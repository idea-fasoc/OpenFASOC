* NGSPICE file created from diff_pair_sample_0810.ext - technology: sky130A

.subckt diff_pair_sample_0810 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t6 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=2.6949 ps=14.6 w=6.91 l=3.91
X1 VTAIL.t3 VN.t0 VDD2.t9 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X2 B.t11 B.t9 B.t10 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=0 ps=0 w=6.91 l=3.91
X3 VDD1.t8 VP.t1 VTAIL.t7 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=1.14015 ps=7.24 w=6.91 l=3.91
X4 VDD2.t8 VN.t1 VTAIL.t16 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X5 VTAIL.t8 VP.t2 VDD1.t7 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X6 VDD1.t6 VP.t3 VTAIL.t9 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=2.6949 ps=14.6 w=6.91 l=3.91
X7 VTAIL.t10 VP.t4 VDD1.t5 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X8 VDD2.t7 VN.t2 VTAIL.t0 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=2.6949 ps=14.6 w=6.91 l=3.91
X9 VTAIL.t2 VN.t3 VDD2.t6 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X10 VDD2.t5 VN.t4 VTAIL.t1 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=1.14015 ps=7.24 w=6.91 l=3.91
X11 VDD2.t4 VN.t5 VTAIL.t5 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=1.14015 ps=7.24 w=6.91 l=3.91
X12 VTAIL.t4 VN.t6 VDD2.t3 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X13 VDD2.t2 VN.t7 VTAIL.t19 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=2.6949 ps=14.6 w=6.91 l=3.91
X14 VTAIL.t11 VP.t5 VDD1.t4 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X15 B.t8 B.t6 B.t7 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=0 ps=0 w=6.91 l=3.91
X16 VDD1.t3 VP.t6 VTAIL.t12 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X17 VTAIL.t13 VP.t7 VDD1.t2 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X18 VDD1.t1 VP.t8 VTAIL.t14 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X19 VDD2.t1 VN.t8 VTAIL.t17 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X20 VTAIL.t18 VN.t9 VDD2.t0 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=1.14015 pd=7.24 as=1.14015 ps=7.24 w=6.91 l=3.91
X21 VDD1.t0 VP.t9 VTAIL.t15 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=1.14015 ps=7.24 w=6.91 l=3.91
X22 B.t5 B.t3 B.t4 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=0 ps=0 w=6.91 l=3.91
X23 B.t2 B.t0 B.t1 w_n6058_n2350# sky130_fd_pr__pfet_01v8 ad=2.6949 pd=14.6 as=0 ps=0 w=6.91 l=3.91
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n25 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n24 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n23 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n53 VP.n22 161.3
R15 VP.n55 VP.n54 161.3
R16 VP.n56 VP.n21 161.3
R17 VP.n59 VP.n58 161.3
R18 VP.n60 VP.n20 161.3
R19 VP.n62 VP.n61 161.3
R20 VP.n63 VP.n19 161.3
R21 VP.n65 VP.n64 161.3
R22 VP.n66 VP.n18 161.3
R23 VP.n68 VP.n67 161.3
R24 VP.n69 VP.n17 161.3
R25 VP.n124 VP.n0 161.3
R26 VP.n123 VP.n122 161.3
R27 VP.n121 VP.n1 161.3
R28 VP.n120 VP.n119 161.3
R29 VP.n118 VP.n2 161.3
R30 VP.n117 VP.n116 161.3
R31 VP.n115 VP.n3 161.3
R32 VP.n114 VP.n113 161.3
R33 VP.n111 VP.n4 161.3
R34 VP.n110 VP.n109 161.3
R35 VP.n108 VP.n5 161.3
R36 VP.n107 VP.n106 161.3
R37 VP.n105 VP.n6 161.3
R38 VP.n104 VP.n103 161.3
R39 VP.n102 VP.n7 161.3
R40 VP.n101 VP.n100 161.3
R41 VP.n99 VP.n8 161.3
R42 VP.n98 VP.n97 161.3
R43 VP.n96 VP.n9 161.3
R44 VP.n95 VP.n94 161.3
R45 VP.n93 VP.n10 161.3
R46 VP.n92 VP.n91 161.3
R47 VP.n90 VP.n11 161.3
R48 VP.n89 VP.n88 161.3
R49 VP.n87 VP.n12 161.3
R50 VP.n85 VP.n84 161.3
R51 VP.n83 VP.n13 161.3
R52 VP.n82 VP.n81 161.3
R53 VP.n80 VP.n14 161.3
R54 VP.n79 VP.n78 161.3
R55 VP.n77 VP.n15 161.3
R56 VP.n76 VP.n75 161.3
R57 VP.n74 VP.n16 161.3
R58 VP.n30 VP.t9 74.666
R59 VP.n31 VP.n30 63.3999
R60 VP.n73 VP.n72 58.6935
R61 VP.n126 VP.n125 58.6935
R62 VP.n71 VP.n70 58.6935
R63 VP.n72 VP.n71 56.6555
R64 VP.n80 VP.n79 54.0911
R65 VP.n119 VP.n118 54.0911
R66 VP.n64 VP.n63 54.0911
R67 VP.n93 VP.n92 52.1486
R68 VP.n106 VP.n105 52.1486
R69 VP.n51 VP.n50 52.1486
R70 VP.n38 VP.n37 52.1486
R71 VP.n99 VP.t8 42.5915
R72 VP.n73 VP.t1 42.5915
R73 VP.n86 VP.t2 42.5915
R74 VP.n112 VP.t5 42.5915
R75 VP.n125 VP.t0 42.5915
R76 VP.n44 VP.t6 42.5915
R77 VP.n70 VP.t3 42.5915
R78 VP.n57 VP.t4 42.5915
R79 VP.n31 VP.t7 42.5915
R80 VP.n94 VP.n93 28.8382
R81 VP.n105 VP.n104 28.8382
R82 VP.n50 VP.n49 28.8382
R83 VP.n39 VP.n38 28.8382
R84 VP.n79 VP.n15 26.8957
R85 VP.n119 VP.n1 26.8957
R86 VP.n64 VP.n18 26.8957
R87 VP.n75 VP.n74 24.4675
R88 VP.n75 VP.n15 24.4675
R89 VP.n81 VP.n80 24.4675
R90 VP.n81 VP.n13 24.4675
R91 VP.n85 VP.n13 24.4675
R92 VP.n88 VP.n87 24.4675
R93 VP.n88 VP.n11 24.4675
R94 VP.n92 VP.n11 24.4675
R95 VP.n94 VP.n9 24.4675
R96 VP.n98 VP.n9 24.4675
R97 VP.n99 VP.n98 24.4675
R98 VP.n100 VP.n99 24.4675
R99 VP.n100 VP.n7 24.4675
R100 VP.n104 VP.n7 24.4675
R101 VP.n106 VP.n5 24.4675
R102 VP.n110 VP.n5 24.4675
R103 VP.n111 VP.n110 24.4675
R104 VP.n113 VP.n3 24.4675
R105 VP.n117 VP.n3 24.4675
R106 VP.n118 VP.n117 24.4675
R107 VP.n123 VP.n1 24.4675
R108 VP.n124 VP.n123 24.4675
R109 VP.n68 VP.n18 24.4675
R110 VP.n69 VP.n68 24.4675
R111 VP.n51 VP.n22 24.4675
R112 VP.n55 VP.n22 24.4675
R113 VP.n56 VP.n55 24.4675
R114 VP.n58 VP.n20 24.4675
R115 VP.n62 VP.n20 24.4675
R116 VP.n63 VP.n62 24.4675
R117 VP.n39 VP.n26 24.4675
R118 VP.n43 VP.n26 24.4675
R119 VP.n44 VP.n43 24.4675
R120 VP.n45 VP.n44 24.4675
R121 VP.n45 VP.n24 24.4675
R122 VP.n49 VP.n24 24.4675
R123 VP.n33 VP.n32 24.4675
R124 VP.n33 VP.n28 24.4675
R125 VP.n37 VP.n28 24.4675
R126 VP.n74 VP.n73 23.4888
R127 VP.n125 VP.n124 23.4888
R128 VP.n70 VP.n69 23.4888
R129 VP.n86 VP.n85 12.7233
R130 VP.n113 VP.n112 12.7233
R131 VP.n58 VP.n57 12.7233
R132 VP.n87 VP.n86 11.7447
R133 VP.n112 VP.n111 11.7447
R134 VP.n57 VP.n56 11.7447
R135 VP.n32 VP.n31 11.7447
R136 VP.n30 VP.n29 2.56981
R137 VP.n71 VP.n17 0.417535
R138 VP.n72 VP.n16 0.417535
R139 VP.n126 VP.n0 0.417535
R140 VP VP.n126 0.394291
R141 VP.n34 VP.n29 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n36 VP.n35 0.189894
R144 VP.n36 VP.n27 0.189894
R145 VP.n40 VP.n27 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n42 VP.n41 0.189894
R148 VP.n42 VP.n25 0.189894
R149 VP.n46 VP.n25 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n48 VP.n47 0.189894
R152 VP.n48 VP.n23 0.189894
R153 VP.n52 VP.n23 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n54 VP.n53 0.189894
R156 VP.n54 VP.n21 0.189894
R157 VP.n59 VP.n21 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n61 VP.n60 0.189894
R160 VP.n61 VP.n19 0.189894
R161 VP.n65 VP.n19 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n67 VP.n66 0.189894
R164 VP.n67 VP.n17 0.189894
R165 VP.n76 VP.n16 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n78 VP.n77 0.189894
R168 VP.n78 VP.n14 0.189894
R169 VP.n82 VP.n14 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n84 VP.n83 0.189894
R172 VP.n84 VP.n12 0.189894
R173 VP.n89 VP.n12 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n91 VP.n90 0.189894
R176 VP.n91 VP.n10 0.189894
R177 VP.n95 VP.n10 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n97 VP.n96 0.189894
R180 VP.n97 VP.n8 0.189894
R181 VP.n101 VP.n8 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n103 VP.n102 0.189894
R184 VP.n103 VP.n6 0.189894
R185 VP.n107 VP.n6 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n109 VP.n108 0.189894
R188 VP.n109 VP.n4 0.189894
R189 VP.n114 VP.n4 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n116 VP.n115 0.189894
R192 VP.n116 VP.n2 0.189894
R193 VP.n120 VP.n2 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n122 VP.n121 0.189894
R196 VP.n122 VP.n0 0.189894
R197 VTAIL.n11 VTAIL.t0 77.9894
R198 VTAIL.n17 VTAIL.t19 77.9893
R199 VTAIL.n2 VTAIL.t6 77.9893
R200 VTAIL.n16 VTAIL.t9 77.9892
R201 VTAIL.n15 VTAIL.n14 73.2853
R202 VTAIL.n13 VTAIL.n12 73.2853
R203 VTAIL.n10 VTAIL.n9 73.2853
R204 VTAIL.n8 VTAIL.n7 73.2853
R205 VTAIL.n19 VTAIL.n18 73.2842
R206 VTAIL.n1 VTAIL.n0 73.2842
R207 VTAIL.n4 VTAIL.n3 73.2842
R208 VTAIL.n6 VTAIL.n5 73.2842
R209 VTAIL.n8 VTAIL.n6 25.6341
R210 VTAIL.n17 VTAIL.n16 21.9789
R211 VTAIL.n18 VTAIL.t16 4.70455
R212 VTAIL.n18 VTAIL.t18 4.70455
R213 VTAIL.n0 VTAIL.t5 4.70455
R214 VTAIL.n0 VTAIL.t3 4.70455
R215 VTAIL.n3 VTAIL.t14 4.70455
R216 VTAIL.n3 VTAIL.t11 4.70455
R217 VTAIL.n5 VTAIL.t7 4.70455
R218 VTAIL.n5 VTAIL.t8 4.70455
R219 VTAIL.n14 VTAIL.t12 4.70455
R220 VTAIL.n14 VTAIL.t10 4.70455
R221 VTAIL.n12 VTAIL.t15 4.70455
R222 VTAIL.n12 VTAIL.t13 4.70455
R223 VTAIL.n9 VTAIL.t17 4.70455
R224 VTAIL.n9 VTAIL.t2 4.70455
R225 VTAIL.n7 VTAIL.t1 4.70455
R226 VTAIL.n7 VTAIL.t4 4.70455
R227 VTAIL.n10 VTAIL.n8 3.65567
R228 VTAIL.n11 VTAIL.n10 3.65567
R229 VTAIL.n15 VTAIL.n13 3.65567
R230 VTAIL.n16 VTAIL.n15 3.65567
R231 VTAIL.n6 VTAIL.n4 3.65567
R232 VTAIL.n4 VTAIL.n2 3.65567
R233 VTAIL.n19 VTAIL.n17 3.65567
R234 VTAIL VTAIL.n1 2.80007
R235 VTAIL.n13 VTAIL.n11 2.29791
R236 VTAIL.n2 VTAIL.n1 2.29791
R237 VTAIL VTAIL.n19 0.856103
R238 VDD1.n1 VDD1.t0 98.3234
R239 VDD1.n3 VDD1.t8 98.3232
R240 VDD1.n5 VDD1.n4 92.649
R241 VDD1.n1 VDD1.n0 89.9641
R242 VDD1.n7 VDD1.n6 89.964
R243 VDD1.n3 VDD1.n2 89.963
R244 VDD1.n7 VDD1.n5 49.4449
R245 VDD1.n6 VDD1.t5 4.70455
R246 VDD1.n6 VDD1.t6 4.70455
R247 VDD1.n0 VDD1.t2 4.70455
R248 VDD1.n0 VDD1.t3 4.70455
R249 VDD1.n4 VDD1.t4 4.70455
R250 VDD1.n4 VDD1.t9 4.70455
R251 VDD1.n2 VDD1.t7 4.70455
R252 VDD1.n2 VDD1.t1 4.70455
R253 VDD1 VDD1.n7 2.68369
R254 VDD1 VDD1.n1 0.972483
R255 VDD1.n5 VDD1.n3 0.858947
R256 VN.n107 VN.n55 161.3
R257 VN.n106 VN.n105 161.3
R258 VN.n104 VN.n56 161.3
R259 VN.n103 VN.n102 161.3
R260 VN.n101 VN.n57 161.3
R261 VN.n100 VN.n99 161.3
R262 VN.n98 VN.n58 161.3
R263 VN.n97 VN.n96 161.3
R264 VN.n94 VN.n59 161.3
R265 VN.n93 VN.n92 161.3
R266 VN.n91 VN.n60 161.3
R267 VN.n90 VN.n89 161.3
R268 VN.n88 VN.n61 161.3
R269 VN.n87 VN.n86 161.3
R270 VN.n85 VN.n62 161.3
R271 VN.n84 VN.n83 161.3
R272 VN.n82 VN.n63 161.3
R273 VN.n81 VN.n80 161.3
R274 VN.n79 VN.n64 161.3
R275 VN.n78 VN.n77 161.3
R276 VN.n76 VN.n65 161.3
R277 VN.n75 VN.n74 161.3
R278 VN.n73 VN.n66 161.3
R279 VN.n72 VN.n71 161.3
R280 VN.n70 VN.n67 161.3
R281 VN.n52 VN.n0 161.3
R282 VN.n51 VN.n50 161.3
R283 VN.n49 VN.n1 161.3
R284 VN.n48 VN.n47 161.3
R285 VN.n46 VN.n2 161.3
R286 VN.n45 VN.n44 161.3
R287 VN.n43 VN.n3 161.3
R288 VN.n42 VN.n41 161.3
R289 VN.n39 VN.n4 161.3
R290 VN.n38 VN.n37 161.3
R291 VN.n36 VN.n5 161.3
R292 VN.n35 VN.n34 161.3
R293 VN.n33 VN.n6 161.3
R294 VN.n32 VN.n31 161.3
R295 VN.n30 VN.n7 161.3
R296 VN.n29 VN.n28 161.3
R297 VN.n27 VN.n8 161.3
R298 VN.n26 VN.n25 161.3
R299 VN.n24 VN.n9 161.3
R300 VN.n23 VN.n22 161.3
R301 VN.n21 VN.n10 161.3
R302 VN.n20 VN.n19 161.3
R303 VN.n18 VN.n11 161.3
R304 VN.n17 VN.n16 161.3
R305 VN.n15 VN.n12 161.3
R306 VN.n13 VN.t5 74.6665
R307 VN.n68 VN.t2 74.6665
R308 VN.n14 VN.n13 63.3999
R309 VN.n69 VN.n68 63.3999
R310 VN.n54 VN.n53 58.6935
R311 VN.n109 VN.n108 58.6935
R312 VN VN.n109 56.6935
R313 VN.n47 VN.n46 54.0911
R314 VN.n102 VN.n101 54.0911
R315 VN.n21 VN.n20 52.1486
R316 VN.n34 VN.n33 52.1486
R317 VN.n76 VN.n75 52.1486
R318 VN.n89 VN.n88 52.1486
R319 VN.n27 VN.t1 42.5915
R320 VN.n14 VN.t0 42.5915
R321 VN.n40 VN.t9 42.5915
R322 VN.n53 VN.t7 42.5915
R323 VN.n82 VN.t8 42.5915
R324 VN.n69 VN.t3 42.5915
R325 VN.n95 VN.t6 42.5915
R326 VN.n108 VN.t4 42.5915
R327 VN.n22 VN.n21 28.8382
R328 VN.n33 VN.n32 28.8382
R329 VN.n77 VN.n76 28.8382
R330 VN.n88 VN.n87 28.8382
R331 VN.n47 VN.n1 26.8957
R332 VN.n102 VN.n56 26.8957
R333 VN.n16 VN.n15 24.4675
R334 VN.n16 VN.n11 24.4675
R335 VN.n20 VN.n11 24.4675
R336 VN.n22 VN.n9 24.4675
R337 VN.n26 VN.n9 24.4675
R338 VN.n27 VN.n26 24.4675
R339 VN.n28 VN.n27 24.4675
R340 VN.n28 VN.n7 24.4675
R341 VN.n32 VN.n7 24.4675
R342 VN.n34 VN.n5 24.4675
R343 VN.n38 VN.n5 24.4675
R344 VN.n39 VN.n38 24.4675
R345 VN.n41 VN.n3 24.4675
R346 VN.n45 VN.n3 24.4675
R347 VN.n46 VN.n45 24.4675
R348 VN.n51 VN.n1 24.4675
R349 VN.n52 VN.n51 24.4675
R350 VN.n75 VN.n66 24.4675
R351 VN.n71 VN.n66 24.4675
R352 VN.n71 VN.n70 24.4675
R353 VN.n87 VN.n62 24.4675
R354 VN.n83 VN.n62 24.4675
R355 VN.n83 VN.n82 24.4675
R356 VN.n82 VN.n81 24.4675
R357 VN.n81 VN.n64 24.4675
R358 VN.n77 VN.n64 24.4675
R359 VN.n101 VN.n100 24.4675
R360 VN.n100 VN.n58 24.4675
R361 VN.n96 VN.n58 24.4675
R362 VN.n94 VN.n93 24.4675
R363 VN.n93 VN.n60 24.4675
R364 VN.n89 VN.n60 24.4675
R365 VN.n107 VN.n106 24.4675
R366 VN.n106 VN.n56 24.4675
R367 VN.n53 VN.n52 23.4888
R368 VN.n108 VN.n107 23.4888
R369 VN.n41 VN.n40 12.7233
R370 VN.n96 VN.n95 12.7233
R371 VN.n15 VN.n14 11.7447
R372 VN.n40 VN.n39 11.7447
R373 VN.n70 VN.n69 11.7447
R374 VN.n95 VN.n94 11.7447
R375 VN.n68 VN.n67 2.56983
R376 VN.n13 VN.n12 2.56983
R377 VN.n109 VN.n55 0.417535
R378 VN.n54 VN.n0 0.417535
R379 VN VN.n54 0.394291
R380 VN.n105 VN.n55 0.189894
R381 VN.n105 VN.n104 0.189894
R382 VN.n104 VN.n103 0.189894
R383 VN.n103 VN.n57 0.189894
R384 VN.n99 VN.n57 0.189894
R385 VN.n99 VN.n98 0.189894
R386 VN.n98 VN.n97 0.189894
R387 VN.n97 VN.n59 0.189894
R388 VN.n92 VN.n59 0.189894
R389 VN.n92 VN.n91 0.189894
R390 VN.n91 VN.n90 0.189894
R391 VN.n90 VN.n61 0.189894
R392 VN.n86 VN.n61 0.189894
R393 VN.n86 VN.n85 0.189894
R394 VN.n85 VN.n84 0.189894
R395 VN.n84 VN.n63 0.189894
R396 VN.n80 VN.n63 0.189894
R397 VN.n80 VN.n79 0.189894
R398 VN.n79 VN.n78 0.189894
R399 VN.n78 VN.n65 0.189894
R400 VN.n74 VN.n65 0.189894
R401 VN.n74 VN.n73 0.189894
R402 VN.n73 VN.n72 0.189894
R403 VN.n72 VN.n67 0.189894
R404 VN.n17 VN.n12 0.189894
R405 VN.n18 VN.n17 0.189894
R406 VN.n19 VN.n18 0.189894
R407 VN.n19 VN.n10 0.189894
R408 VN.n23 VN.n10 0.189894
R409 VN.n24 VN.n23 0.189894
R410 VN.n25 VN.n24 0.189894
R411 VN.n25 VN.n8 0.189894
R412 VN.n29 VN.n8 0.189894
R413 VN.n30 VN.n29 0.189894
R414 VN.n31 VN.n30 0.189894
R415 VN.n31 VN.n6 0.189894
R416 VN.n35 VN.n6 0.189894
R417 VN.n36 VN.n35 0.189894
R418 VN.n37 VN.n36 0.189894
R419 VN.n37 VN.n4 0.189894
R420 VN.n42 VN.n4 0.189894
R421 VN.n43 VN.n42 0.189894
R422 VN.n44 VN.n43 0.189894
R423 VN.n44 VN.n2 0.189894
R424 VN.n48 VN.n2 0.189894
R425 VN.n49 VN.n48 0.189894
R426 VN.n50 VN.n49 0.189894
R427 VN.n50 VN.n0 0.189894
R428 VDD2.n1 VDD2.t4 98.3232
R429 VDD2.n4 VDD2.t5 94.6682
R430 VDD2.n3 VDD2.n2 92.649
R431 VDD2 VDD2.n7 92.6472
R432 VDD2.n6 VDD2.n5 89.9641
R433 VDD2.n1 VDD2.n0 89.963
R434 VDD2.n4 VDD2.n3 47.0343
R435 VDD2.n7 VDD2.t6 4.70455
R436 VDD2.n7 VDD2.t7 4.70455
R437 VDD2.n5 VDD2.t3 4.70455
R438 VDD2.n5 VDD2.t1 4.70455
R439 VDD2.n2 VDD2.t0 4.70455
R440 VDD2.n2 VDD2.t2 4.70455
R441 VDD2.n0 VDD2.t9 4.70455
R442 VDD2.n0 VDD2.t8 4.70455
R443 VDD2.n6 VDD2.n4 3.65567
R444 VDD2 VDD2.n6 0.972483
R445 VDD2.n3 VDD2.n1 0.858947
R446 B.n710 B.n709 585
R447 B.n711 B.n78 585
R448 B.n713 B.n712 585
R449 B.n714 B.n77 585
R450 B.n716 B.n715 585
R451 B.n717 B.n76 585
R452 B.n719 B.n718 585
R453 B.n720 B.n75 585
R454 B.n722 B.n721 585
R455 B.n723 B.n74 585
R456 B.n725 B.n724 585
R457 B.n726 B.n73 585
R458 B.n728 B.n727 585
R459 B.n729 B.n72 585
R460 B.n731 B.n730 585
R461 B.n732 B.n71 585
R462 B.n734 B.n733 585
R463 B.n735 B.n70 585
R464 B.n737 B.n736 585
R465 B.n738 B.n69 585
R466 B.n740 B.n739 585
R467 B.n741 B.n68 585
R468 B.n743 B.n742 585
R469 B.n744 B.n67 585
R470 B.n746 B.n745 585
R471 B.n747 B.n66 585
R472 B.n749 B.n748 585
R473 B.n751 B.n63 585
R474 B.n753 B.n752 585
R475 B.n754 B.n62 585
R476 B.n756 B.n755 585
R477 B.n757 B.n61 585
R478 B.n759 B.n758 585
R479 B.n760 B.n60 585
R480 B.n762 B.n761 585
R481 B.n763 B.n57 585
R482 B.n766 B.n765 585
R483 B.n767 B.n56 585
R484 B.n769 B.n768 585
R485 B.n770 B.n55 585
R486 B.n772 B.n771 585
R487 B.n773 B.n54 585
R488 B.n775 B.n774 585
R489 B.n776 B.n53 585
R490 B.n778 B.n777 585
R491 B.n779 B.n52 585
R492 B.n781 B.n780 585
R493 B.n782 B.n51 585
R494 B.n784 B.n783 585
R495 B.n785 B.n50 585
R496 B.n787 B.n786 585
R497 B.n788 B.n49 585
R498 B.n790 B.n789 585
R499 B.n791 B.n48 585
R500 B.n793 B.n792 585
R501 B.n794 B.n47 585
R502 B.n796 B.n795 585
R503 B.n797 B.n46 585
R504 B.n799 B.n798 585
R505 B.n800 B.n45 585
R506 B.n802 B.n801 585
R507 B.n803 B.n44 585
R508 B.n805 B.n804 585
R509 B.n708 B.n79 585
R510 B.n707 B.n706 585
R511 B.n705 B.n80 585
R512 B.n704 B.n703 585
R513 B.n702 B.n81 585
R514 B.n701 B.n700 585
R515 B.n699 B.n82 585
R516 B.n698 B.n697 585
R517 B.n696 B.n83 585
R518 B.n695 B.n694 585
R519 B.n693 B.n84 585
R520 B.n692 B.n691 585
R521 B.n690 B.n85 585
R522 B.n689 B.n688 585
R523 B.n687 B.n86 585
R524 B.n686 B.n685 585
R525 B.n684 B.n87 585
R526 B.n683 B.n682 585
R527 B.n681 B.n88 585
R528 B.n680 B.n679 585
R529 B.n678 B.n89 585
R530 B.n677 B.n676 585
R531 B.n675 B.n90 585
R532 B.n674 B.n673 585
R533 B.n672 B.n91 585
R534 B.n671 B.n670 585
R535 B.n669 B.n92 585
R536 B.n668 B.n667 585
R537 B.n666 B.n93 585
R538 B.n665 B.n664 585
R539 B.n663 B.n94 585
R540 B.n662 B.n661 585
R541 B.n660 B.n95 585
R542 B.n659 B.n658 585
R543 B.n657 B.n96 585
R544 B.n656 B.n655 585
R545 B.n654 B.n97 585
R546 B.n653 B.n652 585
R547 B.n651 B.n98 585
R548 B.n650 B.n649 585
R549 B.n648 B.n99 585
R550 B.n647 B.n646 585
R551 B.n645 B.n100 585
R552 B.n644 B.n643 585
R553 B.n642 B.n101 585
R554 B.n641 B.n640 585
R555 B.n639 B.n102 585
R556 B.n638 B.n637 585
R557 B.n636 B.n103 585
R558 B.n635 B.n634 585
R559 B.n633 B.n104 585
R560 B.n632 B.n631 585
R561 B.n630 B.n105 585
R562 B.n629 B.n628 585
R563 B.n627 B.n106 585
R564 B.n626 B.n625 585
R565 B.n624 B.n107 585
R566 B.n623 B.n622 585
R567 B.n621 B.n108 585
R568 B.n620 B.n619 585
R569 B.n618 B.n109 585
R570 B.n617 B.n616 585
R571 B.n615 B.n110 585
R572 B.n614 B.n613 585
R573 B.n612 B.n111 585
R574 B.n611 B.n610 585
R575 B.n609 B.n112 585
R576 B.n608 B.n607 585
R577 B.n606 B.n113 585
R578 B.n605 B.n604 585
R579 B.n603 B.n114 585
R580 B.n602 B.n601 585
R581 B.n600 B.n115 585
R582 B.n599 B.n598 585
R583 B.n597 B.n116 585
R584 B.n596 B.n595 585
R585 B.n594 B.n117 585
R586 B.n593 B.n592 585
R587 B.n591 B.n118 585
R588 B.n590 B.n589 585
R589 B.n588 B.n119 585
R590 B.n587 B.n586 585
R591 B.n585 B.n120 585
R592 B.n584 B.n583 585
R593 B.n582 B.n121 585
R594 B.n581 B.n580 585
R595 B.n579 B.n122 585
R596 B.n578 B.n577 585
R597 B.n576 B.n123 585
R598 B.n575 B.n574 585
R599 B.n573 B.n124 585
R600 B.n572 B.n571 585
R601 B.n570 B.n125 585
R602 B.n569 B.n568 585
R603 B.n567 B.n126 585
R604 B.n566 B.n565 585
R605 B.n564 B.n127 585
R606 B.n563 B.n562 585
R607 B.n561 B.n128 585
R608 B.n560 B.n559 585
R609 B.n558 B.n129 585
R610 B.n557 B.n556 585
R611 B.n555 B.n130 585
R612 B.n554 B.n553 585
R613 B.n552 B.n131 585
R614 B.n551 B.n550 585
R615 B.n549 B.n132 585
R616 B.n548 B.n547 585
R617 B.n546 B.n133 585
R618 B.n545 B.n544 585
R619 B.n543 B.n134 585
R620 B.n542 B.n541 585
R621 B.n540 B.n135 585
R622 B.n539 B.n538 585
R623 B.n537 B.n136 585
R624 B.n536 B.n535 585
R625 B.n534 B.n137 585
R626 B.n533 B.n532 585
R627 B.n531 B.n138 585
R628 B.n530 B.n529 585
R629 B.n528 B.n139 585
R630 B.n527 B.n526 585
R631 B.n525 B.n140 585
R632 B.n524 B.n523 585
R633 B.n522 B.n141 585
R634 B.n521 B.n520 585
R635 B.n519 B.n142 585
R636 B.n518 B.n517 585
R637 B.n516 B.n143 585
R638 B.n515 B.n514 585
R639 B.n513 B.n144 585
R640 B.n512 B.n511 585
R641 B.n510 B.n145 585
R642 B.n509 B.n508 585
R643 B.n507 B.n146 585
R644 B.n506 B.n505 585
R645 B.n504 B.n147 585
R646 B.n503 B.n502 585
R647 B.n501 B.n148 585
R648 B.n500 B.n499 585
R649 B.n498 B.n149 585
R650 B.n497 B.n496 585
R651 B.n495 B.n150 585
R652 B.n494 B.n493 585
R653 B.n492 B.n151 585
R654 B.n491 B.n490 585
R655 B.n489 B.n152 585
R656 B.n488 B.n487 585
R657 B.n486 B.n153 585
R658 B.n485 B.n484 585
R659 B.n483 B.n154 585
R660 B.n482 B.n481 585
R661 B.n480 B.n155 585
R662 B.n479 B.n478 585
R663 B.n477 B.n156 585
R664 B.n476 B.n475 585
R665 B.n474 B.n157 585
R666 B.n473 B.n472 585
R667 B.n471 B.n158 585
R668 B.n470 B.n469 585
R669 B.n468 B.n159 585
R670 B.n467 B.n466 585
R671 B.n465 B.n160 585
R672 B.n464 B.n463 585
R673 B.n462 B.n161 585
R674 B.n461 B.n460 585
R675 B.n459 B.n162 585
R676 B.n363 B.n198 585
R677 B.n365 B.n364 585
R678 B.n366 B.n197 585
R679 B.n368 B.n367 585
R680 B.n369 B.n196 585
R681 B.n371 B.n370 585
R682 B.n372 B.n195 585
R683 B.n374 B.n373 585
R684 B.n375 B.n194 585
R685 B.n377 B.n376 585
R686 B.n378 B.n193 585
R687 B.n380 B.n379 585
R688 B.n381 B.n192 585
R689 B.n383 B.n382 585
R690 B.n384 B.n191 585
R691 B.n386 B.n385 585
R692 B.n387 B.n190 585
R693 B.n389 B.n388 585
R694 B.n390 B.n189 585
R695 B.n392 B.n391 585
R696 B.n393 B.n188 585
R697 B.n395 B.n394 585
R698 B.n396 B.n187 585
R699 B.n398 B.n397 585
R700 B.n399 B.n186 585
R701 B.n401 B.n400 585
R702 B.n402 B.n183 585
R703 B.n405 B.n404 585
R704 B.n406 B.n182 585
R705 B.n408 B.n407 585
R706 B.n409 B.n181 585
R707 B.n411 B.n410 585
R708 B.n412 B.n180 585
R709 B.n414 B.n413 585
R710 B.n415 B.n179 585
R711 B.n417 B.n416 585
R712 B.n419 B.n418 585
R713 B.n420 B.n175 585
R714 B.n422 B.n421 585
R715 B.n423 B.n174 585
R716 B.n425 B.n424 585
R717 B.n426 B.n173 585
R718 B.n428 B.n427 585
R719 B.n429 B.n172 585
R720 B.n431 B.n430 585
R721 B.n432 B.n171 585
R722 B.n434 B.n433 585
R723 B.n435 B.n170 585
R724 B.n437 B.n436 585
R725 B.n438 B.n169 585
R726 B.n440 B.n439 585
R727 B.n441 B.n168 585
R728 B.n443 B.n442 585
R729 B.n444 B.n167 585
R730 B.n446 B.n445 585
R731 B.n447 B.n166 585
R732 B.n449 B.n448 585
R733 B.n450 B.n165 585
R734 B.n452 B.n451 585
R735 B.n453 B.n164 585
R736 B.n455 B.n454 585
R737 B.n456 B.n163 585
R738 B.n458 B.n457 585
R739 B.n362 B.n361 585
R740 B.n360 B.n199 585
R741 B.n359 B.n358 585
R742 B.n357 B.n200 585
R743 B.n356 B.n355 585
R744 B.n354 B.n201 585
R745 B.n353 B.n352 585
R746 B.n351 B.n202 585
R747 B.n350 B.n349 585
R748 B.n348 B.n203 585
R749 B.n347 B.n346 585
R750 B.n345 B.n204 585
R751 B.n344 B.n343 585
R752 B.n342 B.n205 585
R753 B.n341 B.n340 585
R754 B.n339 B.n206 585
R755 B.n338 B.n337 585
R756 B.n336 B.n207 585
R757 B.n335 B.n334 585
R758 B.n333 B.n208 585
R759 B.n332 B.n331 585
R760 B.n330 B.n209 585
R761 B.n329 B.n328 585
R762 B.n327 B.n210 585
R763 B.n326 B.n325 585
R764 B.n324 B.n211 585
R765 B.n323 B.n322 585
R766 B.n321 B.n212 585
R767 B.n320 B.n319 585
R768 B.n318 B.n213 585
R769 B.n317 B.n316 585
R770 B.n315 B.n214 585
R771 B.n314 B.n313 585
R772 B.n312 B.n215 585
R773 B.n311 B.n310 585
R774 B.n309 B.n216 585
R775 B.n308 B.n307 585
R776 B.n306 B.n217 585
R777 B.n305 B.n304 585
R778 B.n303 B.n218 585
R779 B.n302 B.n301 585
R780 B.n300 B.n219 585
R781 B.n299 B.n298 585
R782 B.n297 B.n220 585
R783 B.n296 B.n295 585
R784 B.n294 B.n221 585
R785 B.n293 B.n292 585
R786 B.n291 B.n222 585
R787 B.n290 B.n289 585
R788 B.n288 B.n223 585
R789 B.n287 B.n286 585
R790 B.n285 B.n224 585
R791 B.n284 B.n283 585
R792 B.n282 B.n225 585
R793 B.n281 B.n280 585
R794 B.n279 B.n226 585
R795 B.n278 B.n277 585
R796 B.n276 B.n227 585
R797 B.n275 B.n274 585
R798 B.n273 B.n228 585
R799 B.n272 B.n271 585
R800 B.n270 B.n229 585
R801 B.n269 B.n268 585
R802 B.n267 B.n230 585
R803 B.n266 B.n265 585
R804 B.n264 B.n231 585
R805 B.n263 B.n262 585
R806 B.n261 B.n232 585
R807 B.n260 B.n259 585
R808 B.n258 B.n233 585
R809 B.n257 B.n256 585
R810 B.n255 B.n234 585
R811 B.n254 B.n253 585
R812 B.n252 B.n235 585
R813 B.n251 B.n250 585
R814 B.n249 B.n236 585
R815 B.n248 B.n247 585
R816 B.n246 B.n237 585
R817 B.n245 B.n244 585
R818 B.n243 B.n238 585
R819 B.n242 B.n241 585
R820 B.n240 B.n239 585
R821 B.n2 B.n0 585
R822 B.n929 B.n1 585
R823 B.n928 B.n927 585
R824 B.n926 B.n3 585
R825 B.n925 B.n924 585
R826 B.n923 B.n4 585
R827 B.n922 B.n921 585
R828 B.n920 B.n5 585
R829 B.n919 B.n918 585
R830 B.n917 B.n6 585
R831 B.n916 B.n915 585
R832 B.n914 B.n7 585
R833 B.n913 B.n912 585
R834 B.n911 B.n8 585
R835 B.n910 B.n909 585
R836 B.n908 B.n9 585
R837 B.n907 B.n906 585
R838 B.n905 B.n10 585
R839 B.n904 B.n903 585
R840 B.n902 B.n11 585
R841 B.n901 B.n900 585
R842 B.n899 B.n12 585
R843 B.n898 B.n897 585
R844 B.n896 B.n13 585
R845 B.n895 B.n894 585
R846 B.n893 B.n14 585
R847 B.n892 B.n891 585
R848 B.n890 B.n15 585
R849 B.n889 B.n888 585
R850 B.n887 B.n16 585
R851 B.n886 B.n885 585
R852 B.n884 B.n17 585
R853 B.n883 B.n882 585
R854 B.n881 B.n18 585
R855 B.n880 B.n879 585
R856 B.n878 B.n19 585
R857 B.n877 B.n876 585
R858 B.n875 B.n20 585
R859 B.n874 B.n873 585
R860 B.n872 B.n21 585
R861 B.n871 B.n870 585
R862 B.n869 B.n22 585
R863 B.n868 B.n867 585
R864 B.n866 B.n23 585
R865 B.n865 B.n864 585
R866 B.n863 B.n24 585
R867 B.n862 B.n861 585
R868 B.n860 B.n25 585
R869 B.n859 B.n858 585
R870 B.n857 B.n26 585
R871 B.n856 B.n855 585
R872 B.n854 B.n27 585
R873 B.n853 B.n852 585
R874 B.n851 B.n28 585
R875 B.n850 B.n849 585
R876 B.n848 B.n29 585
R877 B.n847 B.n846 585
R878 B.n845 B.n30 585
R879 B.n844 B.n843 585
R880 B.n842 B.n31 585
R881 B.n841 B.n840 585
R882 B.n839 B.n32 585
R883 B.n838 B.n837 585
R884 B.n836 B.n33 585
R885 B.n835 B.n834 585
R886 B.n833 B.n34 585
R887 B.n832 B.n831 585
R888 B.n830 B.n35 585
R889 B.n829 B.n828 585
R890 B.n827 B.n36 585
R891 B.n826 B.n825 585
R892 B.n824 B.n37 585
R893 B.n823 B.n822 585
R894 B.n821 B.n38 585
R895 B.n820 B.n819 585
R896 B.n818 B.n39 585
R897 B.n817 B.n816 585
R898 B.n815 B.n40 585
R899 B.n814 B.n813 585
R900 B.n812 B.n41 585
R901 B.n811 B.n810 585
R902 B.n809 B.n42 585
R903 B.n808 B.n807 585
R904 B.n806 B.n43 585
R905 B.n931 B.n930 585
R906 B.n363 B.n362 478.086
R907 B.n804 B.n43 478.086
R908 B.n459 B.n458 478.086
R909 B.n710 B.n79 478.086
R910 B.n176 B.t3 252.018
R911 B.n184 B.t0 252.018
R912 B.n58 B.t6 252.018
R913 B.n64 B.t9 252.018
R914 B.n176 B.t5 194.042
R915 B.n64 B.t10 194.042
R916 B.n184 B.t2 194.034
R917 B.n58 B.t7 194.034
R918 B.n362 B.n199 163.367
R919 B.n358 B.n199 163.367
R920 B.n358 B.n357 163.367
R921 B.n357 B.n356 163.367
R922 B.n356 B.n201 163.367
R923 B.n352 B.n201 163.367
R924 B.n352 B.n351 163.367
R925 B.n351 B.n350 163.367
R926 B.n350 B.n203 163.367
R927 B.n346 B.n203 163.367
R928 B.n346 B.n345 163.367
R929 B.n345 B.n344 163.367
R930 B.n344 B.n205 163.367
R931 B.n340 B.n205 163.367
R932 B.n340 B.n339 163.367
R933 B.n339 B.n338 163.367
R934 B.n338 B.n207 163.367
R935 B.n334 B.n207 163.367
R936 B.n334 B.n333 163.367
R937 B.n333 B.n332 163.367
R938 B.n332 B.n209 163.367
R939 B.n328 B.n209 163.367
R940 B.n328 B.n327 163.367
R941 B.n327 B.n326 163.367
R942 B.n326 B.n211 163.367
R943 B.n322 B.n211 163.367
R944 B.n322 B.n321 163.367
R945 B.n321 B.n320 163.367
R946 B.n320 B.n213 163.367
R947 B.n316 B.n213 163.367
R948 B.n316 B.n315 163.367
R949 B.n315 B.n314 163.367
R950 B.n314 B.n215 163.367
R951 B.n310 B.n215 163.367
R952 B.n310 B.n309 163.367
R953 B.n309 B.n308 163.367
R954 B.n308 B.n217 163.367
R955 B.n304 B.n217 163.367
R956 B.n304 B.n303 163.367
R957 B.n303 B.n302 163.367
R958 B.n302 B.n219 163.367
R959 B.n298 B.n219 163.367
R960 B.n298 B.n297 163.367
R961 B.n297 B.n296 163.367
R962 B.n296 B.n221 163.367
R963 B.n292 B.n221 163.367
R964 B.n292 B.n291 163.367
R965 B.n291 B.n290 163.367
R966 B.n290 B.n223 163.367
R967 B.n286 B.n223 163.367
R968 B.n286 B.n285 163.367
R969 B.n285 B.n284 163.367
R970 B.n284 B.n225 163.367
R971 B.n280 B.n225 163.367
R972 B.n280 B.n279 163.367
R973 B.n279 B.n278 163.367
R974 B.n278 B.n227 163.367
R975 B.n274 B.n227 163.367
R976 B.n274 B.n273 163.367
R977 B.n273 B.n272 163.367
R978 B.n272 B.n229 163.367
R979 B.n268 B.n229 163.367
R980 B.n268 B.n267 163.367
R981 B.n267 B.n266 163.367
R982 B.n266 B.n231 163.367
R983 B.n262 B.n231 163.367
R984 B.n262 B.n261 163.367
R985 B.n261 B.n260 163.367
R986 B.n260 B.n233 163.367
R987 B.n256 B.n233 163.367
R988 B.n256 B.n255 163.367
R989 B.n255 B.n254 163.367
R990 B.n254 B.n235 163.367
R991 B.n250 B.n235 163.367
R992 B.n250 B.n249 163.367
R993 B.n249 B.n248 163.367
R994 B.n248 B.n237 163.367
R995 B.n244 B.n237 163.367
R996 B.n244 B.n243 163.367
R997 B.n243 B.n242 163.367
R998 B.n242 B.n239 163.367
R999 B.n239 B.n2 163.367
R1000 B.n930 B.n2 163.367
R1001 B.n930 B.n929 163.367
R1002 B.n929 B.n928 163.367
R1003 B.n928 B.n3 163.367
R1004 B.n924 B.n3 163.367
R1005 B.n924 B.n923 163.367
R1006 B.n923 B.n922 163.367
R1007 B.n922 B.n5 163.367
R1008 B.n918 B.n5 163.367
R1009 B.n918 B.n917 163.367
R1010 B.n917 B.n916 163.367
R1011 B.n916 B.n7 163.367
R1012 B.n912 B.n7 163.367
R1013 B.n912 B.n911 163.367
R1014 B.n911 B.n910 163.367
R1015 B.n910 B.n9 163.367
R1016 B.n906 B.n9 163.367
R1017 B.n906 B.n905 163.367
R1018 B.n905 B.n904 163.367
R1019 B.n904 B.n11 163.367
R1020 B.n900 B.n11 163.367
R1021 B.n900 B.n899 163.367
R1022 B.n899 B.n898 163.367
R1023 B.n898 B.n13 163.367
R1024 B.n894 B.n13 163.367
R1025 B.n894 B.n893 163.367
R1026 B.n893 B.n892 163.367
R1027 B.n892 B.n15 163.367
R1028 B.n888 B.n15 163.367
R1029 B.n888 B.n887 163.367
R1030 B.n887 B.n886 163.367
R1031 B.n886 B.n17 163.367
R1032 B.n882 B.n17 163.367
R1033 B.n882 B.n881 163.367
R1034 B.n881 B.n880 163.367
R1035 B.n880 B.n19 163.367
R1036 B.n876 B.n19 163.367
R1037 B.n876 B.n875 163.367
R1038 B.n875 B.n874 163.367
R1039 B.n874 B.n21 163.367
R1040 B.n870 B.n21 163.367
R1041 B.n870 B.n869 163.367
R1042 B.n869 B.n868 163.367
R1043 B.n868 B.n23 163.367
R1044 B.n864 B.n23 163.367
R1045 B.n864 B.n863 163.367
R1046 B.n863 B.n862 163.367
R1047 B.n862 B.n25 163.367
R1048 B.n858 B.n25 163.367
R1049 B.n858 B.n857 163.367
R1050 B.n857 B.n856 163.367
R1051 B.n856 B.n27 163.367
R1052 B.n852 B.n27 163.367
R1053 B.n852 B.n851 163.367
R1054 B.n851 B.n850 163.367
R1055 B.n850 B.n29 163.367
R1056 B.n846 B.n29 163.367
R1057 B.n846 B.n845 163.367
R1058 B.n845 B.n844 163.367
R1059 B.n844 B.n31 163.367
R1060 B.n840 B.n31 163.367
R1061 B.n840 B.n839 163.367
R1062 B.n839 B.n838 163.367
R1063 B.n838 B.n33 163.367
R1064 B.n834 B.n33 163.367
R1065 B.n834 B.n833 163.367
R1066 B.n833 B.n832 163.367
R1067 B.n832 B.n35 163.367
R1068 B.n828 B.n35 163.367
R1069 B.n828 B.n827 163.367
R1070 B.n827 B.n826 163.367
R1071 B.n826 B.n37 163.367
R1072 B.n822 B.n37 163.367
R1073 B.n822 B.n821 163.367
R1074 B.n821 B.n820 163.367
R1075 B.n820 B.n39 163.367
R1076 B.n816 B.n39 163.367
R1077 B.n816 B.n815 163.367
R1078 B.n815 B.n814 163.367
R1079 B.n814 B.n41 163.367
R1080 B.n810 B.n41 163.367
R1081 B.n810 B.n809 163.367
R1082 B.n809 B.n808 163.367
R1083 B.n808 B.n43 163.367
R1084 B.n364 B.n363 163.367
R1085 B.n364 B.n197 163.367
R1086 B.n368 B.n197 163.367
R1087 B.n369 B.n368 163.367
R1088 B.n370 B.n369 163.367
R1089 B.n370 B.n195 163.367
R1090 B.n374 B.n195 163.367
R1091 B.n375 B.n374 163.367
R1092 B.n376 B.n375 163.367
R1093 B.n376 B.n193 163.367
R1094 B.n380 B.n193 163.367
R1095 B.n381 B.n380 163.367
R1096 B.n382 B.n381 163.367
R1097 B.n382 B.n191 163.367
R1098 B.n386 B.n191 163.367
R1099 B.n387 B.n386 163.367
R1100 B.n388 B.n387 163.367
R1101 B.n388 B.n189 163.367
R1102 B.n392 B.n189 163.367
R1103 B.n393 B.n392 163.367
R1104 B.n394 B.n393 163.367
R1105 B.n394 B.n187 163.367
R1106 B.n398 B.n187 163.367
R1107 B.n399 B.n398 163.367
R1108 B.n400 B.n399 163.367
R1109 B.n400 B.n183 163.367
R1110 B.n405 B.n183 163.367
R1111 B.n406 B.n405 163.367
R1112 B.n407 B.n406 163.367
R1113 B.n407 B.n181 163.367
R1114 B.n411 B.n181 163.367
R1115 B.n412 B.n411 163.367
R1116 B.n413 B.n412 163.367
R1117 B.n413 B.n179 163.367
R1118 B.n417 B.n179 163.367
R1119 B.n418 B.n417 163.367
R1120 B.n418 B.n175 163.367
R1121 B.n422 B.n175 163.367
R1122 B.n423 B.n422 163.367
R1123 B.n424 B.n423 163.367
R1124 B.n424 B.n173 163.367
R1125 B.n428 B.n173 163.367
R1126 B.n429 B.n428 163.367
R1127 B.n430 B.n429 163.367
R1128 B.n430 B.n171 163.367
R1129 B.n434 B.n171 163.367
R1130 B.n435 B.n434 163.367
R1131 B.n436 B.n435 163.367
R1132 B.n436 B.n169 163.367
R1133 B.n440 B.n169 163.367
R1134 B.n441 B.n440 163.367
R1135 B.n442 B.n441 163.367
R1136 B.n442 B.n167 163.367
R1137 B.n446 B.n167 163.367
R1138 B.n447 B.n446 163.367
R1139 B.n448 B.n447 163.367
R1140 B.n448 B.n165 163.367
R1141 B.n452 B.n165 163.367
R1142 B.n453 B.n452 163.367
R1143 B.n454 B.n453 163.367
R1144 B.n454 B.n163 163.367
R1145 B.n458 B.n163 163.367
R1146 B.n460 B.n459 163.367
R1147 B.n460 B.n161 163.367
R1148 B.n464 B.n161 163.367
R1149 B.n465 B.n464 163.367
R1150 B.n466 B.n465 163.367
R1151 B.n466 B.n159 163.367
R1152 B.n470 B.n159 163.367
R1153 B.n471 B.n470 163.367
R1154 B.n472 B.n471 163.367
R1155 B.n472 B.n157 163.367
R1156 B.n476 B.n157 163.367
R1157 B.n477 B.n476 163.367
R1158 B.n478 B.n477 163.367
R1159 B.n478 B.n155 163.367
R1160 B.n482 B.n155 163.367
R1161 B.n483 B.n482 163.367
R1162 B.n484 B.n483 163.367
R1163 B.n484 B.n153 163.367
R1164 B.n488 B.n153 163.367
R1165 B.n489 B.n488 163.367
R1166 B.n490 B.n489 163.367
R1167 B.n490 B.n151 163.367
R1168 B.n494 B.n151 163.367
R1169 B.n495 B.n494 163.367
R1170 B.n496 B.n495 163.367
R1171 B.n496 B.n149 163.367
R1172 B.n500 B.n149 163.367
R1173 B.n501 B.n500 163.367
R1174 B.n502 B.n501 163.367
R1175 B.n502 B.n147 163.367
R1176 B.n506 B.n147 163.367
R1177 B.n507 B.n506 163.367
R1178 B.n508 B.n507 163.367
R1179 B.n508 B.n145 163.367
R1180 B.n512 B.n145 163.367
R1181 B.n513 B.n512 163.367
R1182 B.n514 B.n513 163.367
R1183 B.n514 B.n143 163.367
R1184 B.n518 B.n143 163.367
R1185 B.n519 B.n518 163.367
R1186 B.n520 B.n519 163.367
R1187 B.n520 B.n141 163.367
R1188 B.n524 B.n141 163.367
R1189 B.n525 B.n524 163.367
R1190 B.n526 B.n525 163.367
R1191 B.n526 B.n139 163.367
R1192 B.n530 B.n139 163.367
R1193 B.n531 B.n530 163.367
R1194 B.n532 B.n531 163.367
R1195 B.n532 B.n137 163.367
R1196 B.n536 B.n137 163.367
R1197 B.n537 B.n536 163.367
R1198 B.n538 B.n537 163.367
R1199 B.n538 B.n135 163.367
R1200 B.n542 B.n135 163.367
R1201 B.n543 B.n542 163.367
R1202 B.n544 B.n543 163.367
R1203 B.n544 B.n133 163.367
R1204 B.n548 B.n133 163.367
R1205 B.n549 B.n548 163.367
R1206 B.n550 B.n549 163.367
R1207 B.n550 B.n131 163.367
R1208 B.n554 B.n131 163.367
R1209 B.n555 B.n554 163.367
R1210 B.n556 B.n555 163.367
R1211 B.n556 B.n129 163.367
R1212 B.n560 B.n129 163.367
R1213 B.n561 B.n560 163.367
R1214 B.n562 B.n561 163.367
R1215 B.n562 B.n127 163.367
R1216 B.n566 B.n127 163.367
R1217 B.n567 B.n566 163.367
R1218 B.n568 B.n567 163.367
R1219 B.n568 B.n125 163.367
R1220 B.n572 B.n125 163.367
R1221 B.n573 B.n572 163.367
R1222 B.n574 B.n573 163.367
R1223 B.n574 B.n123 163.367
R1224 B.n578 B.n123 163.367
R1225 B.n579 B.n578 163.367
R1226 B.n580 B.n579 163.367
R1227 B.n580 B.n121 163.367
R1228 B.n584 B.n121 163.367
R1229 B.n585 B.n584 163.367
R1230 B.n586 B.n585 163.367
R1231 B.n586 B.n119 163.367
R1232 B.n590 B.n119 163.367
R1233 B.n591 B.n590 163.367
R1234 B.n592 B.n591 163.367
R1235 B.n592 B.n117 163.367
R1236 B.n596 B.n117 163.367
R1237 B.n597 B.n596 163.367
R1238 B.n598 B.n597 163.367
R1239 B.n598 B.n115 163.367
R1240 B.n602 B.n115 163.367
R1241 B.n603 B.n602 163.367
R1242 B.n604 B.n603 163.367
R1243 B.n604 B.n113 163.367
R1244 B.n608 B.n113 163.367
R1245 B.n609 B.n608 163.367
R1246 B.n610 B.n609 163.367
R1247 B.n610 B.n111 163.367
R1248 B.n614 B.n111 163.367
R1249 B.n615 B.n614 163.367
R1250 B.n616 B.n615 163.367
R1251 B.n616 B.n109 163.367
R1252 B.n620 B.n109 163.367
R1253 B.n621 B.n620 163.367
R1254 B.n622 B.n621 163.367
R1255 B.n622 B.n107 163.367
R1256 B.n626 B.n107 163.367
R1257 B.n627 B.n626 163.367
R1258 B.n628 B.n627 163.367
R1259 B.n628 B.n105 163.367
R1260 B.n632 B.n105 163.367
R1261 B.n633 B.n632 163.367
R1262 B.n634 B.n633 163.367
R1263 B.n634 B.n103 163.367
R1264 B.n638 B.n103 163.367
R1265 B.n639 B.n638 163.367
R1266 B.n640 B.n639 163.367
R1267 B.n640 B.n101 163.367
R1268 B.n644 B.n101 163.367
R1269 B.n645 B.n644 163.367
R1270 B.n646 B.n645 163.367
R1271 B.n646 B.n99 163.367
R1272 B.n650 B.n99 163.367
R1273 B.n651 B.n650 163.367
R1274 B.n652 B.n651 163.367
R1275 B.n652 B.n97 163.367
R1276 B.n656 B.n97 163.367
R1277 B.n657 B.n656 163.367
R1278 B.n658 B.n657 163.367
R1279 B.n658 B.n95 163.367
R1280 B.n662 B.n95 163.367
R1281 B.n663 B.n662 163.367
R1282 B.n664 B.n663 163.367
R1283 B.n664 B.n93 163.367
R1284 B.n668 B.n93 163.367
R1285 B.n669 B.n668 163.367
R1286 B.n670 B.n669 163.367
R1287 B.n670 B.n91 163.367
R1288 B.n674 B.n91 163.367
R1289 B.n675 B.n674 163.367
R1290 B.n676 B.n675 163.367
R1291 B.n676 B.n89 163.367
R1292 B.n680 B.n89 163.367
R1293 B.n681 B.n680 163.367
R1294 B.n682 B.n681 163.367
R1295 B.n682 B.n87 163.367
R1296 B.n686 B.n87 163.367
R1297 B.n687 B.n686 163.367
R1298 B.n688 B.n687 163.367
R1299 B.n688 B.n85 163.367
R1300 B.n692 B.n85 163.367
R1301 B.n693 B.n692 163.367
R1302 B.n694 B.n693 163.367
R1303 B.n694 B.n83 163.367
R1304 B.n698 B.n83 163.367
R1305 B.n699 B.n698 163.367
R1306 B.n700 B.n699 163.367
R1307 B.n700 B.n81 163.367
R1308 B.n704 B.n81 163.367
R1309 B.n705 B.n704 163.367
R1310 B.n706 B.n705 163.367
R1311 B.n706 B.n79 163.367
R1312 B.n804 B.n803 163.367
R1313 B.n803 B.n802 163.367
R1314 B.n802 B.n45 163.367
R1315 B.n798 B.n45 163.367
R1316 B.n798 B.n797 163.367
R1317 B.n797 B.n796 163.367
R1318 B.n796 B.n47 163.367
R1319 B.n792 B.n47 163.367
R1320 B.n792 B.n791 163.367
R1321 B.n791 B.n790 163.367
R1322 B.n790 B.n49 163.367
R1323 B.n786 B.n49 163.367
R1324 B.n786 B.n785 163.367
R1325 B.n785 B.n784 163.367
R1326 B.n784 B.n51 163.367
R1327 B.n780 B.n51 163.367
R1328 B.n780 B.n779 163.367
R1329 B.n779 B.n778 163.367
R1330 B.n778 B.n53 163.367
R1331 B.n774 B.n53 163.367
R1332 B.n774 B.n773 163.367
R1333 B.n773 B.n772 163.367
R1334 B.n772 B.n55 163.367
R1335 B.n768 B.n55 163.367
R1336 B.n768 B.n767 163.367
R1337 B.n767 B.n766 163.367
R1338 B.n766 B.n57 163.367
R1339 B.n761 B.n57 163.367
R1340 B.n761 B.n760 163.367
R1341 B.n760 B.n759 163.367
R1342 B.n759 B.n61 163.367
R1343 B.n755 B.n61 163.367
R1344 B.n755 B.n754 163.367
R1345 B.n754 B.n753 163.367
R1346 B.n753 B.n63 163.367
R1347 B.n748 B.n63 163.367
R1348 B.n748 B.n747 163.367
R1349 B.n747 B.n746 163.367
R1350 B.n746 B.n67 163.367
R1351 B.n742 B.n67 163.367
R1352 B.n742 B.n741 163.367
R1353 B.n741 B.n740 163.367
R1354 B.n740 B.n69 163.367
R1355 B.n736 B.n69 163.367
R1356 B.n736 B.n735 163.367
R1357 B.n735 B.n734 163.367
R1358 B.n734 B.n71 163.367
R1359 B.n730 B.n71 163.367
R1360 B.n730 B.n729 163.367
R1361 B.n729 B.n728 163.367
R1362 B.n728 B.n73 163.367
R1363 B.n724 B.n73 163.367
R1364 B.n724 B.n723 163.367
R1365 B.n723 B.n722 163.367
R1366 B.n722 B.n75 163.367
R1367 B.n718 B.n75 163.367
R1368 B.n718 B.n717 163.367
R1369 B.n717 B.n716 163.367
R1370 B.n716 B.n77 163.367
R1371 B.n712 B.n77 163.367
R1372 B.n712 B.n711 163.367
R1373 B.n711 B.n710 163.367
R1374 B.n177 B.t4 111.811
R1375 B.n65 B.t11 111.811
R1376 B.n185 B.t1 111.803
R1377 B.n59 B.t8 111.803
R1378 B.n177 B.n176 82.2308
R1379 B.n185 B.n184 82.2308
R1380 B.n59 B.n58 82.2308
R1381 B.n65 B.n64 82.2308
R1382 B.n178 B.n177 59.5399
R1383 B.n403 B.n185 59.5399
R1384 B.n764 B.n59 59.5399
R1385 B.n750 B.n65 59.5399
R1386 B.n806 B.n805 31.0639
R1387 B.n709 B.n708 31.0639
R1388 B.n457 B.n162 31.0639
R1389 B.n361 B.n198 31.0639
R1390 B B.n931 18.0485
R1391 B.n805 B.n44 10.6151
R1392 B.n801 B.n44 10.6151
R1393 B.n801 B.n800 10.6151
R1394 B.n800 B.n799 10.6151
R1395 B.n799 B.n46 10.6151
R1396 B.n795 B.n46 10.6151
R1397 B.n795 B.n794 10.6151
R1398 B.n794 B.n793 10.6151
R1399 B.n793 B.n48 10.6151
R1400 B.n789 B.n48 10.6151
R1401 B.n789 B.n788 10.6151
R1402 B.n788 B.n787 10.6151
R1403 B.n787 B.n50 10.6151
R1404 B.n783 B.n50 10.6151
R1405 B.n783 B.n782 10.6151
R1406 B.n782 B.n781 10.6151
R1407 B.n781 B.n52 10.6151
R1408 B.n777 B.n52 10.6151
R1409 B.n777 B.n776 10.6151
R1410 B.n776 B.n775 10.6151
R1411 B.n775 B.n54 10.6151
R1412 B.n771 B.n54 10.6151
R1413 B.n771 B.n770 10.6151
R1414 B.n770 B.n769 10.6151
R1415 B.n769 B.n56 10.6151
R1416 B.n765 B.n56 10.6151
R1417 B.n763 B.n762 10.6151
R1418 B.n762 B.n60 10.6151
R1419 B.n758 B.n60 10.6151
R1420 B.n758 B.n757 10.6151
R1421 B.n757 B.n756 10.6151
R1422 B.n756 B.n62 10.6151
R1423 B.n752 B.n62 10.6151
R1424 B.n752 B.n751 10.6151
R1425 B.n749 B.n66 10.6151
R1426 B.n745 B.n66 10.6151
R1427 B.n745 B.n744 10.6151
R1428 B.n744 B.n743 10.6151
R1429 B.n743 B.n68 10.6151
R1430 B.n739 B.n68 10.6151
R1431 B.n739 B.n738 10.6151
R1432 B.n738 B.n737 10.6151
R1433 B.n737 B.n70 10.6151
R1434 B.n733 B.n70 10.6151
R1435 B.n733 B.n732 10.6151
R1436 B.n732 B.n731 10.6151
R1437 B.n731 B.n72 10.6151
R1438 B.n727 B.n72 10.6151
R1439 B.n727 B.n726 10.6151
R1440 B.n726 B.n725 10.6151
R1441 B.n725 B.n74 10.6151
R1442 B.n721 B.n74 10.6151
R1443 B.n721 B.n720 10.6151
R1444 B.n720 B.n719 10.6151
R1445 B.n719 B.n76 10.6151
R1446 B.n715 B.n76 10.6151
R1447 B.n715 B.n714 10.6151
R1448 B.n714 B.n713 10.6151
R1449 B.n713 B.n78 10.6151
R1450 B.n709 B.n78 10.6151
R1451 B.n461 B.n162 10.6151
R1452 B.n462 B.n461 10.6151
R1453 B.n463 B.n462 10.6151
R1454 B.n463 B.n160 10.6151
R1455 B.n467 B.n160 10.6151
R1456 B.n468 B.n467 10.6151
R1457 B.n469 B.n468 10.6151
R1458 B.n469 B.n158 10.6151
R1459 B.n473 B.n158 10.6151
R1460 B.n474 B.n473 10.6151
R1461 B.n475 B.n474 10.6151
R1462 B.n475 B.n156 10.6151
R1463 B.n479 B.n156 10.6151
R1464 B.n480 B.n479 10.6151
R1465 B.n481 B.n480 10.6151
R1466 B.n481 B.n154 10.6151
R1467 B.n485 B.n154 10.6151
R1468 B.n486 B.n485 10.6151
R1469 B.n487 B.n486 10.6151
R1470 B.n487 B.n152 10.6151
R1471 B.n491 B.n152 10.6151
R1472 B.n492 B.n491 10.6151
R1473 B.n493 B.n492 10.6151
R1474 B.n493 B.n150 10.6151
R1475 B.n497 B.n150 10.6151
R1476 B.n498 B.n497 10.6151
R1477 B.n499 B.n498 10.6151
R1478 B.n499 B.n148 10.6151
R1479 B.n503 B.n148 10.6151
R1480 B.n504 B.n503 10.6151
R1481 B.n505 B.n504 10.6151
R1482 B.n505 B.n146 10.6151
R1483 B.n509 B.n146 10.6151
R1484 B.n510 B.n509 10.6151
R1485 B.n511 B.n510 10.6151
R1486 B.n511 B.n144 10.6151
R1487 B.n515 B.n144 10.6151
R1488 B.n516 B.n515 10.6151
R1489 B.n517 B.n516 10.6151
R1490 B.n517 B.n142 10.6151
R1491 B.n521 B.n142 10.6151
R1492 B.n522 B.n521 10.6151
R1493 B.n523 B.n522 10.6151
R1494 B.n523 B.n140 10.6151
R1495 B.n527 B.n140 10.6151
R1496 B.n528 B.n527 10.6151
R1497 B.n529 B.n528 10.6151
R1498 B.n529 B.n138 10.6151
R1499 B.n533 B.n138 10.6151
R1500 B.n534 B.n533 10.6151
R1501 B.n535 B.n534 10.6151
R1502 B.n535 B.n136 10.6151
R1503 B.n539 B.n136 10.6151
R1504 B.n540 B.n539 10.6151
R1505 B.n541 B.n540 10.6151
R1506 B.n541 B.n134 10.6151
R1507 B.n545 B.n134 10.6151
R1508 B.n546 B.n545 10.6151
R1509 B.n547 B.n546 10.6151
R1510 B.n547 B.n132 10.6151
R1511 B.n551 B.n132 10.6151
R1512 B.n552 B.n551 10.6151
R1513 B.n553 B.n552 10.6151
R1514 B.n553 B.n130 10.6151
R1515 B.n557 B.n130 10.6151
R1516 B.n558 B.n557 10.6151
R1517 B.n559 B.n558 10.6151
R1518 B.n559 B.n128 10.6151
R1519 B.n563 B.n128 10.6151
R1520 B.n564 B.n563 10.6151
R1521 B.n565 B.n564 10.6151
R1522 B.n565 B.n126 10.6151
R1523 B.n569 B.n126 10.6151
R1524 B.n570 B.n569 10.6151
R1525 B.n571 B.n570 10.6151
R1526 B.n571 B.n124 10.6151
R1527 B.n575 B.n124 10.6151
R1528 B.n576 B.n575 10.6151
R1529 B.n577 B.n576 10.6151
R1530 B.n577 B.n122 10.6151
R1531 B.n581 B.n122 10.6151
R1532 B.n582 B.n581 10.6151
R1533 B.n583 B.n582 10.6151
R1534 B.n583 B.n120 10.6151
R1535 B.n587 B.n120 10.6151
R1536 B.n588 B.n587 10.6151
R1537 B.n589 B.n588 10.6151
R1538 B.n589 B.n118 10.6151
R1539 B.n593 B.n118 10.6151
R1540 B.n594 B.n593 10.6151
R1541 B.n595 B.n594 10.6151
R1542 B.n595 B.n116 10.6151
R1543 B.n599 B.n116 10.6151
R1544 B.n600 B.n599 10.6151
R1545 B.n601 B.n600 10.6151
R1546 B.n601 B.n114 10.6151
R1547 B.n605 B.n114 10.6151
R1548 B.n606 B.n605 10.6151
R1549 B.n607 B.n606 10.6151
R1550 B.n607 B.n112 10.6151
R1551 B.n611 B.n112 10.6151
R1552 B.n612 B.n611 10.6151
R1553 B.n613 B.n612 10.6151
R1554 B.n613 B.n110 10.6151
R1555 B.n617 B.n110 10.6151
R1556 B.n618 B.n617 10.6151
R1557 B.n619 B.n618 10.6151
R1558 B.n619 B.n108 10.6151
R1559 B.n623 B.n108 10.6151
R1560 B.n624 B.n623 10.6151
R1561 B.n625 B.n624 10.6151
R1562 B.n625 B.n106 10.6151
R1563 B.n629 B.n106 10.6151
R1564 B.n630 B.n629 10.6151
R1565 B.n631 B.n630 10.6151
R1566 B.n631 B.n104 10.6151
R1567 B.n635 B.n104 10.6151
R1568 B.n636 B.n635 10.6151
R1569 B.n637 B.n636 10.6151
R1570 B.n637 B.n102 10.6151
R1571 B.n641 B.n102 10.6151
R1572 B.n642 B.n641 10.6151
R1573 B.n643 B.n642 10.6151
R1574 B.n643 B.n100 10.6151
R1575 B.n647 B.n100 10.6151
R1576 B.n648 B.n647 10.6151
R1577 B.n649 B.n648 10.6151
R1578 B.n649 B.n98 10.6151
R1579 B.n653 B.n98 10.6151
R1580 B.n654 B.n653 10.6151
R1581 B.n655 B.n654 10.6151
R1582 B.n655 B.n96 10.6151
R1583 B.n659 B.n96 10.6151
R1584 B.n660 B.n659 10.6151
R1585 B.n661 B.n660 10.6151
R1586 B.n661 B.n94 10.6151
R1587 B.n665 B.n94 10.6151
R1588 B.n666 B.n665 10.6151
R1589 B.n667 B.n666 10.6151
R1590 B.n667 B.n92 10.6151
R1591 B.n671 B.n92 10.6151
R1592 B.n672 B.n671 10.6151
R1593 B.n673 B.n672 10.6151
R1594 B.n673 B.n90 10.6151
R1595 B.n677 B.n90 10.6151
R1596 B.n678 B.n677 10.6151
R1597 B.n679 B.n678 10.6151
R1598 B.n679 B.n88 10.6151
R1599 B.n683 B.n88 10.6151
R1600 B.n684 B.n683 10.6151
R1601 B.n685 B.n684 10.6151
R1602 B.n685 B.n86 10.6151
R1603 B.n689 B.n86 10.6151
R1604 B.n690 B.n689 10.6151
R1605 B.n691 B.n690 10.6151
R1606 B.n691 B.n84 10.6151
R1607 B.n695 B.n84 10.6151
R1608 B.n696 B.n695 10.6151
R1609 B.n697 B.n696 10.6151
R1610 B.n697 B.n82 10.6151
R1611 B.n701 B.n82 10.6151
R1612 B.n702 B.n701 10.6151
R1613 B.n703 B.n702 10.6151
R1614 B.n703 B.n80 10.6151
R1615 B.n707 B.n80 10.6151
R1616 B.n708 B.n707 10.6151
R1617 B.n365 B.n198 10.6151
R1618 B.n366 B.n365 10.6151
R1619 B.n367 B.n366 10.6151
R1620 B.n367 B.n196 10.6151
R1621 B.n371 B.n196 10.6151
R1622 B.n372 B.n371 10.6151
R1623 B.n373 B.n372 10.6151
R1624 B.n373 B.n194 10.6151
R1625 B.n377 B.n194 10.6151
R1626 B.n378 B.n377 10.6151
R1627 B.n379 B.n378 10.6151
R1628 B.n379 B.n192 10.6151
R1629 B.n383 B.n192 10.6151
R1630 B.n384 B.n383 10.6151
R1631 B.n385 B.n384 10.6151
R1632 B.n385 B.n190 10.6151
R1633 B.n389 B.n190 10.6151
R1634 B.n390 B.n389 10.6151
R1635 B.n391 B.n390 10.6151
R1636 B.n391 B.n188 10.6151
R1637 B.n395 B.n188 10.6151
R1638 B.n396 B.n395 10.6151
R1639 B.n397 B.n396 10.6151
R1640 B.n397 B.n186 10.6151
R1641 B.n401 B.n186 10.6151
R1642 B.n402 B.n401 10.6151
R1643 B.n404 B.n182 10.6151
R1644 B.n408 B.n182 10.6151
R1645 B.n409 B.n408 10.6151
R1646 B.n410 B.n409 10.6151
R1647 B.n410 B.n180 10.6151
R1648 B.n414 B.n180 10.6151
R1649 B.n415 B.n414 10.6151
R1650 B.n416 B.n415 10.6151
R1651 B.n420 B.n419 10.6151
R1652 B.n421 B.n420 10.6151
R1653 B.n421 B.n174 10.6151
R1654 B.n425 B.n174 10.6151
R1655 B.n426 B.n425 10.6151
R1656 B.n427 B.n426 10.6151
R1657 B.n427 B.n172 10.6151
R1658 B.n431 B.n172 10.6151
R1659 B.n432 B.n431 10.6151
R1660 B.n433 B.n432 10.6151
R1661 B.n433 B.n170 10.6151
R1662 B.n437 B.n170 10.6151
R1663 B.n438 B.n437 10.6151
R1664 B.n439 B.n438 10.6151
R1665 B.n439 B.n168 10.6151
R1666 B.n443 B.n168 10.6151
R1667 B.n444 B.n443 10.6151
R1668 B.n445 B.n444 10.6151
R1669 B.n445 B.n166 10.6151
R1670 B.n449 B.n166 10.6151
R1671 B.n450 B.n449 10.6151
R1672 B.n451 B.n450 10.6151
R1673 B.n451 B.n164 10.6151
R1674 B.n455 B.n164 10.6151
R1675 B.n456 B.n455 10.6151
R1676 B.n457 B.n456 10.6151
R1677 B.n361 B.n360 10.6151
R1678 B.n360 B.n359 10.6151
R1679 B.n359 B.n200 10.6151
R1680 B.n355 B.n200 10.6151
R1681 B.n355 B.n354 10.6151
R1682 B.n354 B.n353 10.6151
R1683 B.n353 B.n202 10.6151
R1684 B.n349 B.n202 10.6151
R1685 B.n349 B.n348 10.6151
R1686 B.n348 B.n347 10.6151
R1687 B.n347 B.n204 10.6151
R1688 B.n343 B.n204 10.6151
R1689 B.n343 B.n342 10.6151
R1690 B.n342 B.n341 10.6151
R1691 B.n341 B.n206 10.6151
R1692 B.n337 B.n206 10.6151
R1693 B.n337 B.n336 10.6151
R1694 B.n336 B.n335 10.6151
R1695 B.n335 B.n208 10.6151
R1696 B.n331 B.n208 10.6151
R1697 B.n331 B.n330 10.6151
R1698 B.n330 B.n329 10.6151
R1699 B.n329 B.n210 10.6151
R1700 B.n325 B.n210 10.6151
R1701 B.n325 B.n324 10.6151
R1702 B.n324 B.n323 10.6151
R1703 B.n323 B.n212 10.6151
R1704 B.n319 B.n212 10.6151
R1705 B.n319 B.n318 10.6151
R1706 B.n318 B.n317 10.6151
R1707 B.n317 B.n214 10.6151
R1708 B.n313 B.n214 10.6151
R1709 B.n313 B.n312 10.6151
R1710 B.n312 B.n311 10.6151
R1711 B.n311 B.n216 10.6151
R1712 B.n307 B.n216 10.6151
R1713 B.n307 B.n306 10.6151
R1714 B.n306 B.n305 10.6151
R1715 B.n305 B.n218 10.6151
R1716 B.n301 B.n218 10.6151
R1717 B.n301 B.n300 10.6151
R1718 B.n300 B.n299 10.6151
R1719 B.n299 B.n220 10.6151
R1720 B.n295 B.n220 10.6151
R1721 B.n295 B.n294 10.6151
R1722 B.n294 B.n293 10.6151
R1723 B.n293 B.n222 10.6151
R1724 B.n289 B.n222 10.6151
R1725 B.n289 B.n288 10.6151
R1726 B.n288 B.n287 10.6151
R1727 B.n287 B.n224 10.6151
R1728 B.n283 B.n224 10.6151
R1729 B.n283 B.n282 10.6151
R1730 B.n282 B.n281 10.6151
R1731 B.n281 B.n226 10.6151
R1732 B.n277 B.n226 10.6151
R1733 B.n277 B.n276 10.6151
R1734 B.n276 B.n275 10.6151
R1735 B.n275 B.n228 10.6151
R1736 B.n271 B.n228 10.6151
R1737 B.n271 B.n270 10.6151
R1738 B.n270 B.n269 10.6151
R1739 B.n269 B.n230 10.6151
R1740 B.n265 B.n230 10.6151
R1741 B.n265 B.n264 10.6151
R1742 B.n264 B.n263 10.6151
R1743 B.n263 B.n232 10.6151
R1744 B.n259 B.n232 10.6151
R1745 B.n259 B.n258 10.6151
R1746 B.n258 B.n257 10.6151
R1747 B.n257 B.n234 10.6151
R1748 B.n253 B.n234 10.6151
R1749 B.n253 B.n252 10.6151
R1750 B.n252 B.n251 10.6151
R1751 B.n251 B.n236 10.6151
R1752 B.n247 B.n236 10.6151
R1753 B.n247 B.n246 10.6151
R1754 B.n246 B.n245 10.6151
R1755 B.n245 B.n238 10.6151
R1756 B.n241 B.n238 10.6151
R1757 B.n241 B.n240 10.6151
R1758 B.n240 B.n0 10.6151
R1759 B.n927 B.n1 10.6151
R1760 B.n927 B.n926 10.6151
R1761 B.n926 B.n925 10.6151
R1762 B.n925 B.n4 10.6151
R1763 B.n921 B.n4 10.6151
R1764 B.n921 B.n920 10.6151
R1765 B.n920 B.n919 10.6151
R1766 B.n919 B.n6 10.6151
R1767 B.n915 B.n6 10.6151
R1768 B.n915 B.n914 10.6151
R1769 B.n914 B.n913 10.6151
R1770 B.n913 B.n8 10.6151
R1771 B.n909 B.n8 10.6151
R1772 B.n909 B.n908 10.6151
R1773 B.n908 B.n907 10.6151
R1774 B.n907 B.n10 10.6151
R1775 B.n903 B.n10 10.6151
R1776 B.n903 B.n902 10.6151
R1777 B.n902 B.n901 10.6151
R1778 B.n901 B.n12 10.6151
R1779 B.n897 B.n12 10.6151
R1780 B.n897 B.n896 10.6151
R1781 B.n896 B.n895 10.6151
R1782 B.n895 B.n14 10.6151
R1783 B.n891 B.n14 10.6151
R1784 B.n891 B.n890 10.6151
R1785 B.n890 B.n889 10.6151
R1786 B.n889 B.n16 10.6151
R1787 B.n885 B.n16 10.6151
R1788 B.n885 B.n884 10.6151
R1789 B.n884 B.n883 10.6151
R1790 B.n883 B.n18 10.6151
R1791 B.n879 B.n18 10.6151
R1792 B.n879 B.n878 10.6151
R1793 B.n878 B.n877 10.6151
R1794 B.n877 B.n20 10.6151
R1795 B.n873 B.n20 10.6151
R1796 B.n873 B.n872 10.6151
R1797 B.n872 B.n871 10.6151
R1798 B.n871 B.n22 10.6151
R1799 B.n867 B.n22 10.6151
R1800 B.n867 B.n866 10.6151
R1801 B.n866 B.n865 10.6151
R1802 B.n865 B.n24 10.6151
R1803 B.n861 B.n24 10.6151
R1804 B.n861 B.n860 10.6151
R1805 B.n860 B.n859 10.6151
R1806 B.n859 B.n26 10.6151
R1807 B.n855 B.n26 10.6151
R1808 B.n855 B.n854 10.6151
R1809 B.n854 B.n853 10.6151
R1810 B.n853 B.n28 10.6151
R1811 B.n849 B.n28 10.6151
R1812 B.n849 B.n848 10.6151
R1813 B.n848 B.n847 10.6151
R1814 B.n847 B.n30 10.6151
R1815 B.n843 B.n30 10.6151
R1816 B.n843 B.n842 10.6151
R1817 B.n842 B.n841 10.6151
R1818 B.n841 B.n32 10.6151
R1819 B.n837 B.n32 10.6151
R1820 B.n837 B.n836 10.6151
R1821 B.n836 B.n835 10.6151
R1822 B.n835 B.n34 10.6151
R1823 B.n831 B.n34 10.6151
R1824 B.n831 B.n830 10.6151
R1825 B.n830 B.n829 10.6151
R1826 B.n829 B.n36 10.6151
R1827 B.n825 B.n36 10.6151
R1828 B.n825 B.n824 10.6151
R1829 B.n824 B.n823 10.6151
R1830 B.n823 B.n38 10.6151
R1831 B.n819 B.n38 10.6151
R1832 B.n819 B.n818 10.6151
R1833 B.n818 B.n817 10.6151
R1834 B.n817 B.n40 10.6151
R1835 B.n813 B.n40 10.6151
R1836 B.n813 B.n812 10.6151
R1837 B.n812 B.n811 10.6151
R1838 B.n811 B.n42 10.6151
R1839 B.n807 B.n42 10.6151
R1840 B.n807 B.n806 10.6151
R1841 B.n764 B.n763 6.5566
R1842 B.n751 B.n750 6.5566
R1843 B.n404 B.n403 6.5566
R1844 B.n416 B.n178 6.5566
R1845 B.n765 B.n764 4.05904
R1846 B.n750 B.n749 4.05904
R1847 B.n403 B.n402 4.05904
R1848 B.n419 B.n178 4.05904
R1849 B.n931 B.n0 2.81026
R1850 B.n931 B.n1 2.81026
C0 VDD2 B 2.74558f
C1 VDD2 VN 6.8071f
C2 VTAIL VDD1 9.146541f
C3 VTAIL VP 8.552621f
C4 VN B 1.5554f
C5 VDD1 w_n6058_n2350# 2.93736f
C6 VP w_n6058_n2350# 14.0567f
C7 VDD2 VTAIL 9.20805f
C8 VDD2 w_n6058_n2350# 3.149f
C9 VTAIL B 2.99378f
C10 VTAIL VN 8.53806f
C11 VP VDD1 7.39779f
C12 B w_n6058_n2350# 11.3274f
C13 VN w_n6058_n2350# 13.263901f
C14 VDD2 VDD1 3.02786f
C15 VDD2 VP 0.750115f
C16 B VDD1 2.57665f
C17 VN VDD1 0.156396f
C18 VP B 2.89571f
C19 VTAIL w_n6058_n2350# 2.71789f
C20 VN VP 9.389111f
C21 VDD2 VSUBS 2.615233f
C22 VDD1 VSUBS 2.416192f
C23 VTAIL VSUBS 0.841801f
C24 VN VSUBS 9.65397f
C25 VP VSUBS 5.440804f
C26 B VSUBS 6.561634f
C27 w_n6058_n2350# VSUBS 0.17716p
C28 B.n0 VSUBS 0.006884f
C29 B.n1 VSUBS 0.006884f
C30 B.n2 VSUBS 0.010886f
C31 B.n3 VSUBS 0.010886f
C32 B.n4 VSUBS 0.010886f
C33 B.n5 VSUBS 0.010886f
C34 B.n6 VSUBS 0.010886f
C35 B.n7 VSUBS 0.010886f
C36 B.n8 VSUBS 0.010886f
C37 B.n9 VSUBS 0.010886f
C38 B.n10 VSUBS 0.010886f
C39 B.n11 VSUBS 0.010886f
C40 B.n12 VSUBS 0.010886f
C41 B.n13 VSUBS 0.010886f
C42 B.n14 VSUBS 0.010886f
C43 B.n15 VSUBS 0.010886f
C44 B.n16 VSUBS 0.010886f
C45 B.n17 VSUBS 0.010886f
C46 B.n18 VSUBS 0.010886f
C47 B.n19 VSUBS 0.010886f
C48 B.n20 VSUBS 0.010886f
C49 B.n21 VSUBS 0.010886f
C50 B.n22 VSUBS 0.010886f
C51 B.n23 VSUBS 0.010886f
C52 B.n24 VSUBS 0.010886f
C53 B.n25 VSUBS 0.010886f
C54 B.n26 VSUBS 0.010886f
C55 B.n27 VSUBS 0.010886f
C56 B.n28 VSUBS 0.010886f
C57 B.n29 VSUBS 0.010886f
C58 B.n30 VSUBS 0.010886f
C59 B.n31 VSUBS 0.010886f
C60 B.n32 VSUBS 0.010886f
C61 B.n33 VSUBS 0.010886f
C62 B.n34 VSUBS 0.010886f
C63 B.n35 VSUBS 0.010886f
C64 B.n36 VSUBS 0.010886f
C65 B.n37 VSUBS 0.010886f
C66 B.n38 VSUBS 0.010886f
C67 B.n39 VSUBS 0.010886f
C68 B.n40 VSUBS 0.010886f
C69 B.n41 VSUBS 0.010886f
C70 B.n42 VSUBS 0.010886f
C71 B.n43 VSUBS 0.02401f
C72 B.n44 VSUBS 0.010886f
C73 B.n45 VSUBS 0.010886f
C74 B.n46 VSUBS 0.010886f
C75 B.n47 VSUBS 0.010886f
C76 B.n48 VSUBS 0.010886f
C77 B.n49 VSUBS 0.010886f
C78 B.n50 VSUBS 0.010886f
C79 B.n51 VSUBS 0.010886f
C80 B.n52 VSUBS 0.010886f
C81 B.n53 VSUBS 0.010886f
C82 B.n54 VSUBS 0.010886f
C83 B.n55 VSUBS 0.010886f
C84 B.n56 VSUBS 0.010886f
C85 B.n57 VSUBS 0.010886f
C86 B.t8 VSUBS 0.32299f
C87 B.t7 VSUBS 0.366867f
C88 B.t6 VSUBS 2.01168f
C89 B.n58 VSUBS 0.220952f
C90 B.n59 VSUBS 0.11906f
C91 B.n60 VSUBS 0.010886f
C92 B.n61 VSUBS 0.010886f
C93 B.n62 VSUBS 0.010886f
C94 B.n63 VSUBS 0.010886f
C95 B.t11 VSUBS 0.322988f
C96 B.t10 VSUBS 0.366864f
C97 B.t9 VSUBS 2.01168f
C98 B.n64 VSUBS 0.220954f
C99 B.n65 VSUBS 0.119062f
C100 B.n66 VSUBS 0.010886f
C101 B.n67 VSUBS 0.010886f
C102 B.n68 VSUBS 0.010886f
C103 B.n69 VSUBS 0.010886f
C104 B.n70 VSUBS 0.010886f
C105 B.n71 VSUBS 0.010886f
C106 B.n72 VSUBS 0.010886f
C107 B.n73 VSUBS 0.010886f
C108 B.n74 VSUBS 0.010886f
C109 B.n75 VSUBS 0.010886f
C110 B.n76 VSUBS 0.010886f
C111 B.n77 VSUBS 0.010886f
C112 B.n78 VSUBS 0.010886f
C113 B.n79 VSUBS 0.02401f
C114 B.n80 VSUBS 0.010886f
C115 B.n81 VSUBS 0.010886f
C116 B.n82 VSUBS 0.010886f
C117 B.n83 VSUBS 0.010886f
C118 B.n84 VSUBS 0.010886f
C119 B.n85 VSUBS 0.010886f
C120 B.n86 VSUBS 0.010886f
C121 B.n87 VSUBS 0.010886f
C122 B.n88 VSUBS 0.010886f
C123 B.n89 VSUBS 0.010886f
C124 B.n90 VSUBS 0.010886f
C125 B.n91 VSUBS 0.010886f
C126 B.n92 VSUBS 0.010886f
C127 B.n93 VSUBS 0.010886f
C128 B.n94 VSUBS 0.010886f
C129 B.n95 VSUBS 0.010886f
C130 B.n96 VSUBS 0.010886f
C131 B.n97 VSUBS 0.010886f
C132 B.n98 VSUBS 0.010886f
C133 B.n99 VSUBS 0.010886f
C134 B.n100 VSUBS 0.010886f
C135 B.n101 VSUBS 0.010886f
C136 B.n102 VSUBS 0.010886f
C137 B.n103 VSUBS 0.010886f
C138 B.n104 VSUBS 0.010886f
C139 B.n105 VSUBS 0.010886f
C140 B.n106 VSUBS 0.010886f
C141 B.n107 VSUBS 0.010886f
C142 B.n108 VSUBS 0.010886f
C143 B.n109 VSUBS 0.010886f
C144 B.n110 VSUBS 0.010886f
C145 B.n111 VSUBS 0.010886f
C146 B.n112 VSUBS 0.010886f
C147 B.n113 VSUBS 0.010886f
C148 B.n114 VSUBS 0.010886f
C149 B.n115 VSUBS 0.010886f
C150 B.n116 VSUBS 0.010886f
C151 B.n117 VSUBS 0.010886f
C152 B.n118 VSUBS 0.010886f
C153 B.n119 VSUBS 0.010886f
C154 B.n120 VSUBS 0.010886f
C155 B.n121 VSUBS 0.010886f
C156 B.n122 VSUBS 0.010886f
C157 B.n123 VSUBS 0.010886f
C158 B.n124 VSUBS 0.010886f
C159 B.n125 VSUBS 0.010886f
C160 B.n126 VSUBS 0.010886f
C161 B.n127 VSUBS 0.010886f
C162 B.n128 VSUBS 0.010886f
C163 B.n129 VSUBS 0.010886f
C164 B.n130 VSUBS 0.010886f
C165 B.n131 VSUBS 0.010886f
C166 B.n132 VSUBS 0.010886f
C167 B.n133 VSUBS 0.010886f
C168 B.n134 VSUBS 0.010886f
C169 B.n135 VSUBS 0.010886f
C170 B.n136 VSUBS 0.010886f
C171 B.n137 VSUBS 0.010886f
C172 B.n138 VSUBS 0.010886f
C173 B.n139 VSUBS 0.010886f
C174 B.n140 VSUBS 0.010886f
C175 B.n141 VSUBS 0.010886f
C176 B.n142 VSUBS 0.010886f
C177 B.n143 VSUBS 0.010886f
C178 B.n144 VSUBS 0.010886f
C179 B.n145 VSUBS 0.010886f
C180 B.n146 VSUBS 0.010886f
C181 B.n147 VSUBS 0.010886f
C182 B.n148 VSUBS 0.010886f
C183 B.n149 VSUBS 0.010886f
C184 B.n150 VSUBS 0.010886f
C185 B.n151 VSUBS 0.010886f
C186 B.n152 VSUBS 0.010886f
C187 B.n153 VSUBS 0.010886f
C188 B.n154 VSUBS 0.010886f
C189 B.n155 VSUBS 0.010886f
C190 B.n156 VSUBS 0.010886f
C191 B.n157 VSUBS 0.010886f
C192 B.n158 VSUBS 0.010886f
C193 B.n159 VSUBS 0.010886f
C194 B.n160 VSUBS 0.010886f
C195 B.n161 VSUBS 0.010886f
C196 B.n162 VSUBS 0.02401f
C197 B.n163 VSUBS 0.010886f
C198 B.n164 VSUBS 0.010886f
C199 B.n165 VSUBS 0.010886f
C200 B.n166 VSUBS 0.010886f
C201 B.n167 VSUBS 0.010886f
C202 B.n168 VSUBS 0.010886f
C203 B.n169 VSUBS 0.010886f
C204 B.n170 VSUBS 0.010886f
C205 B.n171 VSUBS 0.010886f
C206 B.n172 VSUBS 0.010886f
C207 B.n173 VSUBS 0.010886f
C208 B.n174 VSUBS 0.010886f
C209 B.n175 VSUBS 0.010886f
C210 B.t4 VSUBS 0.322988f
C211 B.t5 VSUBS 0.366864f
C212 B.t3 VSUBS 2.01168f
C213 B.n176 VSUBS 0.220954f
C214 B.n177 VSUBS 0.119062f
C215 B.n178 VSUBS 0.025221f
C216 B.n179 VSUBS 0.010886f
C217 B.n180 VSUBS 0.010886f
C218 B.n181 VSUBS 0.010886f
C219 B.n182 VSUBS 0.010886f
C220 B.n183 VSUBS 0.010886f
C221 B.t1 VSUBS 0.32299f
C222 B.t2 VSUBS 0.366867f
C223 B.t0 VSUBS 2.01168f
C224 B.n184 VSUBS 0.220952f
C225 B.n185 VSUBS 0.11906f
C226 B.n186 VSUBS 0.010886f
C227 B.n187 VSUBS 0.010886f
C228 B.n188 VSUBS 0.010886f
C229 B.n189 VSUBS 0.010886f
C230 B.n190 VSUBS 0.010886f
C231 B.n191 VSUBS 0.010886f
C232 B.n192 VSUBS 0.010886f
C233 B.n193 VSUBS 0.010886f
C234 B.n194 VSUBS 0.010886f
C235 B.n195 VSUBS 0.010886f
C236 B.n196 VSUBS 0.010886f
C237 B.n197 VSUBS 0.010886f
C238 B.n198 VSUBS 0.025296f
C239 B.n199 VSUBS 0.010886f
C240 B.n200 VSUBS 0.010886f
C241 B.n201 VSUBS 0.010886f
C242 B.n202 VSUBS 0.010886f
C243 B.n203 VSUBS 0.010886f
C244 B.n204 VSUBS 0.010886f
C245 B.n205 VSUBS 0.010886f
C246 B.n206 VSUBS 0.010886f
C247 B.n207 VSUBS 0.010886f
C248 B.n208 VSUBS 0.010886f
C249 B.n209 VSUBS 0.010886f
C250 B.n210 VSUBS 0.010886f
C251 B.n211 VSUBS 0.010886f
C252 B.n212 VSUBS 0.010886f
C253 B.n213 VSUBS 0.010886f
C254 B.n214 VSUBS 0.010886f
C255 B.n215 VSUBS 0.010886f
C256 B.n216 VSUBS 0.010886f
C257 B.n217 VSUBS 0.010886f
C258 B.n218 VSUBS 0.010886f
C259 B.n219 VSUBS 0.010886f
C260 B.n220 VSUBS 0.010886f
C261 B.n221 VSUBS 0.010886f
C262 B.n222 VSUBS 0.010886f
C263 B.n223 VSUBS 0.010886f
C264 B.n224 VSUBS 0.010886f
C265 B.n225 VSUBS 0.010886f
C266 B.n226 VSUBS 0.010886f
C267 B.n227 VSUBS 0.010886f
C268 B.n228 VSUBS 0.010886f
C269 B.n229 VSUBS 0.010886f
C270 B.n230 VSUBS 0.010886f
C271 B.n231 VSUBS 0.010886f
C272 B.n232 VSUBS 0.010886f
C273 B.n233 VSUBS 0.010886f
C274 B.n234 VSUBS 0.010886f
C275 B.n235 VSUBS 0.010886f
C276 B.n236 VSUBS 0.010886f
C277 B.n237 VSUBS 0.010886f
C278 B.n238 VSUBS 0.010886f
C279 B.n239 VSUBS 0.010886f
C280 B.n240 VSUBS 0.010886f
C281 B.n241 VSUBS 0.010886f
C282 B.n242 VSUBS 0.010886f
C283 B.n243 VSUBS 0.010886f
C284 B.n244 VSUBS 0.010886f
C285 B.n245 VSUBS 0.010886f
C286 B.n246 VSUBS 0.010886f
C287 B.n247 VSUBS 0.010886f
C288 B.n248 VSUBS 0.010886f
C289 B.n249 VSUBS 0.010886f
C290 B.n250 VSUBS 0.010886f
C291 B.n251 VSUBS 0.010886f
C292 B.n252 VSUBS 0.010886f
C293 B.n253 VSUBS 0.010886f
C294 B.n254 VSUBS 0.010886f
C295 B.n255 VSUBS 0.010886f
C296 B.n256 VSUBS 0.010886f
C297 B.n257 VSUBS 0.010886f
C298 B.n258 VSUBS 0.010886f
C299 B.n259 VSUBS 0.010886f
C300 B.n260 VSUBS 0.010886f
C301 B.n261 VSUBS 0.010886f
C302 B.n262 VSUBS 0.010886f
C303 B.n263 VSUBS 0.010886f
C304 B.n264 VSUBS 0.010886f
C305 B.n265 VSUBS 0.010886f
C306 B.n266 VSUBS 0.010886f
C307 B.n267 VSUBS 0.010886f
C308 B.n268 VSUBS 0.010886f
C309 B.n269 VSUBS 0.010886f
C310 B.n270 VSUBS 0.010886f
C311 B.n271 VSUBS 0.010886f
C312 B.n272 VSUBS 0.010886f
C313 B.n273 VSUBS 0.010886f
C314 B.n274 VSUBS 0.010886f
C315 B.n275 VSUBS 0.010886f
C316 B.n276 VSUBS 0.010886f
C317 B.n277 VSUBS 0.010886f
C318 B.n278 VSUBS 0.010886f
C319 B.n279 VSUBS 0.010886f
C320 B.n280 VSUBS 0.010886f
C321 B.n281 VSUBS 0.010886f
C322 B.n282 VSUBS 0.010886f
C323 B.n283 VSUBS 0.010886f
C324 B.n284 VSUBS 0.010886f
C325 B.n285 VSUBS 0.010886f
C326 B.n286 VSUBS 0.010886f
C327 B.n287 VSUBS 0.010886f
C328 B.n288 VSUBS 0.010886f
C329 B.n289 VSUBS 0.010886f
C330 B.n290 VSUBS 0.010886f
C331 B.n291 VSUBS 0.010886f
C332 B.n292 VSUBS 0.010886f
C333 B.n293 VSUBS 0.010886f
C334 B.n294 VSUBS 0.010886f
C335 B.n295 VSUBS 0.010886f
C336 B.n296 VSUBS 0.010886f
C337 B.n297 VSUBS 0.010886f
C338 B.n298 VSUBS 0.010886f
C339 B.n299 VSUBS 0.010886f
C340 B.n300 VSUBS 0.010886f
C341 B.n301 VSUBS 0.010886f
C342 B.n302 VSUBS 0.010886f
C343 B.n303 VSUBS 0.010886f
C344 B.n304 VSUBS 0.010886f
C345 B.n305 VSUBS 0.010886f
C346 B.n306 VSUBS 0.010886f
C347 B.n307 VSUBS 0.010886f
C348 B.n308 VSUBS 0.010886f
C349 B.n309 VSUBS 0.010886f
C350 B.n310 VSUBS 0.010886f
C351 B.n311 VSUBS 0.010886f
C352 B.n312 VSUBS 0.010886f
C353 B.n313 VSUBS 0.010886f
C354 B.n314 VSUBS 0.010886f
C355 B.n315 VSUBS 0.010886f
C356 B.n316 VSUBS 0.010886f
C357 B.n317 VSUBS 0.010886f
C358 B.n318 VSUBS 0.010886f
C359 B.n319 VSUBS 0.010886f
C360 B.n320 VSUBS 0.010886f
C361 B.n321 VSUBS 0.010886f
C362 B.n322 VSUBS 0.010886f
C363 B.n323 VSUBS 0.010886f
C364 B.n324 VSUBS 0.010886f
C365 B.n325 VSUBS 0.010886f
C366 B.n326 VSUBS 0.010886f
C367 B.n327 VSUBS 0.010886f
C368 B.n328 VSUBS 0.010886f
C369 B.n329 VSUBS 0.010886f
C370 B.n330 VSUBS 0.010886f
C371 B.n331 VSUBS 0.010886f
C372 B.n332 VSUBS 0.010886f
C373 B.n333 VSUBS 0.010886f
C374 B.n334 VSUBS 0.010886f
C375 B.n335 VSUBS 0.010886f
C376 B.n336 VSUBS 0.010886f
C377 B.n337 VSUBS 0.010886f
C378 B.n338 VSUBS 0.010886f
C379 B.n339 VSUBS 0.010886f
C380 B.n340 VSUBS 0.010886f
C381 B.n341 VSUBS 0.010886f
C382 B.n342 VSUBS 0.010886f
C383 B.n343 VSUBS 0.010886f
C384 B.n344 VSUBS 0.010886f
C385 B.n345 VSUBS 0.010886f
C386 B.n346 VSUBS 0.010886f
C387 B.n347 VSUBS 0.010886f
C388 B.n348 VSUBS 0.010886f
C389 B.n349 VSUBS 0.010886f
C390 B.n350 VSUBS 0.010886f
C391 B.n351 VSUBS 0.010886f
C392 B.n352 VSUBS 0.010886f
C393 B.n353 VSUBS 0.010886f
C394 B.n354 VSUBS 0.010886f
C395 B.n355 VSUBS 0.010886f
C396 B.n356 VSUBS 0.010886f
C397 B.n357 VSUBS 0.010886f
C398 B.n358 VSUBS 0.010886f
C399 B.n359 VSUBS 0.010886f
C400 B.n360 VSUBS 0.010886f
C401 B.n361 VSUBS 0.02401f
C402 B.n362 VSUBS 0.02401f
C403 B.n363 VSUBS 0.025296f
C404 B.n364 VSUBS 0.010886f
C405 B.n365 VSUBS 0.010886f
C406 B.n366 VSUBS 0.010886f
C407 B.n367 VSUBS 0.010886f
C408 B.n368 VSUBS 0.010886f
C409 B.n369 VSUBS 0.010886f
C410 B.n370 VSUBS 0.010886f
C411 B.n371 VSUBS 0.010886f
C412 B.n372 VSUBS 0.010886f
C413 B.n373 VSUBS 0.010886f
C414 B.n374 VSUBS 0.010886f
C415 B.n375 VSUBS 0.010886f
C416 B.n376 VSUBS 0.010886f
C417 B.n377 VSUBS 0.010886f
C418 B.n378 VSUBS 0.010886f
C419 B.n379 VSUBS 0.010886f
C420 B.n380 VSUBS 0.010886f
C421 B.n381 VSUBS 0.010886f
C422 B.n382 VSUBS 0.010886f
C423 B.n383 VSUBS 0.010886f
C424 B.n384 VSUBS 0.010886f
C425 B.n385 VSUBS 0.010886f
C426 B.n386 VSUBS 0.010886f
C427 B.n387 VSUBS 0.010886f
C428 B.n388 VSUBS 0.010886f
C429 B.n389 VSUBS 0.010886f
C430 B.n390 VSUBS 0.010886f
C431 B.n391 VSUBS 0.010886f
C432 B.n392 VSUBS 0.010886f
C433 B.n393 VSUBS 0.010886f
C434 B.n394 VSUBS 0.010886f
C435 B.n395 VSUBS 0.010886f
C436 B.n396 VSUBS 0.010886f
C437 B.n397 VSUBS 0.010886f
C438 B.n398 VSUBS 0.010886f
C439 B.n399 VSUBS 0.010886f
C440 B.n400 VSUBS 0.010886f
C441 B.n401 VSUBS 0.010886f
C442 B.n402 VSUBS 0.007524f
C443 B.n403 VSUBS 0.025221f
C444 B.n404 VSUBS 0.008805f
C445 B.n405 VSUBS 0.010886f
C446 B.n406 VSUBS 0.010886f
C447 B.n407 VSUBS 0.010886f
C448 B.n408 VSUBS 0.010886f
C449 B.n409 VSUBS 0.010886f
C450 B.n410 VSUBS 0.010886f
C451 B.n411 VSUBS 0.010886f
C452 B.n412 VSUBS 0.010886f
C453 B.n413 VSUBS 0.010886f
C454 B.n414 VSUBS 0.010886f
C455 B.n415 VSUBS 0.010886f
C456 B.n416 VSUBS 0.008805f
C457 B.n417 VSUBS 0.010886f
C458 B.n418 VSUBS 0.010886f
C459 B.n419 VSUBS 0.007524f
C460 B.n420 VSUBS 0.010886f
C461 B.n421 VSUBS 0.010886f
C462 B.n422 VSUBS 0.010886f
C463 B.n423 VSUBS 0.010886f
C464 B.n424 VSUBS 0.010886f
C465 B.n425 VSUBS 0.010886f
C466 B.n426 VSUBS 0.010886f
C467 B.n427 VSUBS 0.010886f
C468 B.n428 VSUBS 0.010886f
C469 B.n429 VSUBS 0.010886f
C470 B.n430 VSUBS 0.010886f
C471 B.n431 VSUBS 0.010886f
C472 B.n432 VSUBS 0.010886f
C473 B.n433 VSUBS 0.010886f
C474 B.n434 VSUBS 0.010886f
C475 B.n435 VSUBS 0.010886f
C476 B.n436 VSUBS 0.010886f
C477 B.n437 VSUBS 0.010886f
C478 B.n438 VSUBS 0.010886f
C479 B.n439 VSUBS 0.010886f
C480 B.n440 VSUBS 0.010886f
C481 B.n441 VSUBS 0.010886f
C482 B.n442 VSUBS 0.010886f
C483 B.n443 VSUBS 0.010886f
C484 B.n444 VSUBS 0.010886f
C485 B.n445 VSUBS 0.010886f
C486 B.n446 VSUBS 0.010886f
C487 B.n447 VSUBS 0.010886f
C488 B.n448 VSUBS 0.010886f
C489 B.n449 VSUBS 0.010886f
C490 B.n450 VSUBS 0.010886f
C491 B.n451 VSUBS 0.010886f
C492 B.n452 VSUBS 0.010886f
C493 B.n453 VSUBS 0.010886f
C494 B.n454 VSUBS 0.010886f
C495 B.n455 VSUBS 0.010886f
C496 B.n456 VSUBS 0.010886f
C497 B.n457 VSUBS 0.025296f
C498 B.n458 VSUBS 0.025296f
C499 B.n459 VSUBS 0.02401f
C500 B.n460 VSUBS 0.010886f
C501 B.n461 VSUBS 0.010886f
C502 B.n462 VSUBS 0.010886f
C503 B.n463 VSUBS 0.010886f
C504 B.n464 VSUBS 0.010886f
C505 B.n465 VSUBS 0.010886f
C506 B.n466 VSUBS 0.010886f
C507 B.n467 VSUBS 0.010886f
C508 B.n468 VSUBS 0.010886f
C509 B.n469 VSUBS 0.010886f
C510 B.n470 VSUBS 0.010886f
C511 B.n471 VSUBS 0.010886f
C512 B.n472 VSUBS 0.010886f
C513 B.n473 VSUBS 0.010886f
C514 B.n474 VSUBS 0.010886f
C515 B.n475 VSUBS 0.010886f
C516 B.n476 VSUBS 0.010886f
C517 B.n477 VSUBS 0.010886f
C518 B.n478 VSUBS 0.010886f
C519 B.n479 VSUBS 0.010886f
C520 B.n480 VSUBS 0.010886f
C521 B.n481 VSUBS 0.010886f
C522 B.n482 VSUBS 0.010886f
C523 B.n483 VSUBS 0.010886f
C524 B.n484 VSUBS 0.010886f
C525 B.n485 VSUBS 0.010886f
C526 B.n486 VSUBS 0.010886f
C527 B.n487 VSUBS 0.010886f
C528 B.n488 VSUBS 0.010886f
C529 B.n489 VSUBS 0.010886f
C530 B.n490 VSUBS 0.010886f
C531 B.n491 VSUBS 0.010886f
C532 B.n492 VSUBS 0.010886f
C533 B.n493 VSUBS 0.010886f
C534 B.n494 VSUBS 0.010886f
C535 B.n495 VSUBS 0.010886f
C536 B.n496 VSUBS 0.010886f
C537 B.n497 VSUBS 0.010886f
C538 B.n498 VSUBS 0.010886f
C539 B.n499 VSUBS 0.010886f
C540 B.n500 VSUBS 0.010886f
C541 B.n501 VSUBS 0.010886f
C542 B.n502 VSUBS 0.010886f
C543 B.n503 VSUBS 0.010886f
C544 B.n504 VSUBS 0.010886f
C545 B.n505 VSUBS 0.010886f
C546 B.n506 VSUBS 0.010886f
C547 B.n507 VSUBS 0.010886f
C548 B.n508 VSUBS 0.010886f
C549 B.n509 VSUBS 0.010886f
C550 B.n510 VSUBS 0.010886f
C551 B.n511 VSUBS 0.010886f
C552 B.n512 VSUBS 0.010886f
C553 B.n513 VSUBS 0.010886f
C554 B.n514 VSUBS 0.010886f
C555 B.n515 VSUBS 0.010886f
C556 B.n516 VSUBS 0.010886f
C557 B.n517 VSUBS 0.010886f
C558 B.n518 VSUBS 0.010886f
C559 B.n519 VSUBS 0.010886f
C560 B.n520 VSUBS 0.010886f
C561 B.n521 VSUBS 0.010886f
C562 B.n522 VSUBS 0.010886f
C563 B.n523 VSUBS 0.010886f
C564 B.n524 VSUBS 0.010886f
C565 B.n525 VSUBS 0.010886f
C566 B.n526 VSUBS 0.010886f
C567 B.n527 VSUBS 0.010886f
C568 B.n528 VSUBS 0.010886f
C569 B.n529 VSUBS 0.010886f
C570 B.n530 VSUBS 0.010886f
C571 B.n531 VSUBS 0.010886f
C572 B.n532 VSUBS 0.010886f
C573 B.n533 VSUBS 0.010886f
C574 B.n534 VSUBS 0.010886f
C575 B.n535 VSUBS 0.010886f
C576 B.n536 VSUBS 0.010886f
C577 B.n537 VSUBS 0.010886f
C578 B.n538 VSUBS 0.010886f
C579 B.n539 VSUBS 0.010886f
C580 B.n540 VSUBS 0.010886f
C581 B.n541 VSUBS 0.010886f
C582 B.n542 VSUBS 0.010886f
C583 B.n543 VSUBS 0.010886f
C584 B.n544 VSUBS 0.010886f
C585 B.n545 VSUBS 0.010886f
C586 B.n546 VSUBS 0.010886f
C587 B.n547 VSUBS 0.010886f
C588 B.n548 VSUBS 0.010886f
C589 B.n549 VSUBS 0.010886f
C590 B.n550 VSUBS 0.010886f
C591 B.n551 VSUBS 0.010886f
C592 B.n552 VSUBS 0.010886f
C593 B.n553 VSUBS 0.010886f
C594 B.n554 VSUBS 0.010886f
C595 B.n555 VSUBS 0.010886f
C596 B.n556 VSUBS 0.010886f
C597 B.n557 VSUBS 0.010886f
C598 B.n558 VSUBS 0.010886f
C599 B.n559 VSUBS 0.010886f
C600 B.n560 VSUBS 0.010886f
C601 B.n561 VSUBS 0.010886f
C602 B.n562 VSUBS 0.010886f
C603 B.n563 VSUBS 0.010886f
C604 B.n564 VSUBS 0.010886f
C605 B.n565 VSUBS 0.010886f
C606 B.n566 VSUBS 0.010886f
C607 B.n567 VSUBS 0.010886f
C608 B.n568 VSUBS 0.010886f
C609 B.n569 VSUBS 0.010886f
C610 B.n570 VSUBS 0.010886f
C611 B.n571 VSUBS 0.010886f
C612 B.n572 VSUBS 0.010886f
C613 B.n573 VSUBS 0.010886f
C614 B.n574 VSUBS 0.010886f
C615 B.n575 VSUBS 0.010886f
C616 B.n576 VSUBS 0.010886f
C617 B.n577 VSUBS 0.010886f
C618 B.n578 VSUBS 0.010886f
C619 B.n579 VSUBS 0.010886f
C620 B.n580 VSUBS 0.010886f
C621 B.n581 VSUBS 0.010886f
C622 B.n582 VSUBS 0.010886f
C623 B.n583 VSUBS 0.010886f
C624 B.n584 VSUBS 0.010886f
C625 B.n585 VSUBS 0.010886f
C626 B.n586 VSUBS 0.010886f
C627 B.n587 VSUBS 0.010886f
C628 B.n588 VSUBS 0.010886f
C629 B.n589 VSUBS 0.010886f
C630 B.n590 VSUBS 0.010886f
C631 B.n591 VSUBS 0.010886f
C632 B.n592 VSUBS 0.010886f
C633 B.n593 VSUBS 0.010886f
C634 B.n594 VSUBS 0.010886f
C635 B.n595 VSUBS 0.010886f
C636 B.n596 VSUBS 0.010886f
C637 B.n597 VSUBS 0.010886f
C638 B.n598 VSUBS 0.010886f
C639 B.n599 VSUBS 0.010886f
C640 B.n600 VSUBS 0.010886f
C641 B.n601 VSUBS 0.010886f
C642 B.n602 VSUBS 0.010886f
C643 B.n603 VSUBS 0.010886f
C644 B.n604 VSUBS 0.010886f
C645 B.n605 VSUBS 0.010886f
C646 B.n606 VSUBS 0.010886f
C647 B.n607 VSUBS 0.010886f
C648 B.n608 VSUBS 0.010886f
C649 B.n609 VSUBS 0.010886f
C650 B.n610 VSUBS 0.010886f
C651 B.n611 VSUBS 0.010886f
C652 B.n612 VSUBS 0.010886f
C653 B.n613 VSUBS 0.010886f
C654 B.n614 VSUBS 0.010886f
C655 B.n615 VSUBS 0.010886f
C656 B.n616 VSUBS 0.010886f
C657 B.n617 VSUBS 0.010886f
C658 B.n618 VSUBS 0.010886f
C659 B.n619 VSUBS 0.010886f
C660 B.n620 VSUBS 0.010886f
C661 B.n621 VSUBS 0.010886f
C662 B.n622 VSUBS 0.010886f
C663 B.n623 VSUBS 0.010886f
C664 B.n624 VSUBS 0.010886f
C665 B.n625 VSUBS 0.010886f
C666 B.n626 VSUBS 0.010886f
C667 B.n627 VSUBS 0.010886f
C668 B.n628 VSUBS 0.010886f
C669 B.n629 VSUBS 0.010886f
C670 B.n630 VSUBS 0.010886f
C671 B.n631 VSUBS 0.010886f
C672 B.n632 VSUBS 0.010886f
C673 B.n633 VSUBS 0.010886f
C674 B.n634 VSUBS 0.010886f
C675 B.n635 VSUBS 0.010886f
C676 B.n636 VSUBS 0.010886f
C677 B.n637 VSUBS 0.010886f
C678 B.n638 VSUBS 0.010886f
C679 B.n639 VSUBS 0.010886f
C680 B.n640 VSUBS 0.010886f
C681 B.n641 VSUBS 0.010886f
C682 B.n642 VSUBS 0.010886f
C683 B.n643 VSUBS 0.010886f
C684 B.n644 VSUBS 0.010886f
C685 B.n645 VSUBS 0.010886f
C686 B.n646 VSUBS 0.010886f
C687 B.n647 VSUBS 0.010886f
C688 B.n648 VSUBS 0.010886f
C689 B.n649 VSUBS 0.010886f
C690 B.n650 VSUBS 0.010886f
C691 B.n651 VSUBS 0.010886f
C692 B.n652 VSUBS 0.010886f
C693 B.n653 VSUBS 0.010886f
C694 B.n654 VSUBS 0.010886f
C695 B.n655 VSUBS 0.010886f
C696 B.n656 VSUBS 0.010886f
C697 B.n657 VSUBS 0.010886f
C698 B.n658 VSUBS 0.010886f
C699 B.n659 VSUBS 0.010886f
C700 B.n660 VSUBS 0.010886f
C701 B.n661 VSUBS 0.010886f
C702 B.n662 VSUBS 0.010886f
C703 B.n663 VSUBS 0.010886f
C704 B.n664 VSUBS 0.010886f
C705 B.n665 VSUBS 0.010886f
C706 B.n666 VSUBS 0.010886f
C707 B.n667 VSUBS 0.010886f
C708 B.n668 VSUBS 0.010886f
C709 B.n669 VSUBS 0.010886f
C710 B.n670 VSUBS 0.010886f
C711 B.n671 VSUBS 0.010886f
C712 B.n672 VSUBS 0.010886f
C713 B.n673 VSUBS 0.010886f
C714 B.n674 VSUBS 0.010886f
C715 B.n675 VSUBS 0.010886f
C716 B.n676 VSUBS 0.010886f
C717 B.n677 VSUBS 0.010886f
C718 B.n678 VSUBS 0.010886f
C719 B.n679 VSUBS 0.010886f
C720 B.n680 VSUBS 0.010886f
C721 B.n681 VSUBS 0.010886f
C722 B.n682 VSUBS 0.010886f
C723 B.n683 VSUBS 0.010886f
C724 B.n684 VSUBS 0.010886f
C725 B.n685 VSUBS 0.010886f
C726 B.n686 VSUBS 0.010886f
C727 B.n687 VSUBS 0.010886f
C728 B.n688 VSUBS 0.010886f
C729 B.n689 VSUBS 0.010886f
C730 B.n690 VSUBS 0.010886f
C731 B.n691 VSUBS 0.010886f
C732 B.n692 VSUBS 0.010886f
C733 B.n693 VSUBS 0.010886f
C734 B.n694 VSUBS 0.010886f
C735 B.n695 VSUBS 0.010886f
C736 B.n696 VSUBS 0.010886f
C737 B.n697 VSUBS 0.010886f
C738 B.n698 VSUBS 0.010886f
C739 B.n699 VSUBS 0.010886f
C740 B.n700 VSUBS 0.010886f
C741 B.n701 VSUBS 0.010886f
C742 B.n702 VSUBS 0.010886f
C743 B.n703 VSUBS 0.010886f
C744 B.n704 VSUBS 0.010886f
C745 B.n705 VSUBS 0.010886f
C746 B.n706 VSUBS 0.010886f
C747 B.n707 VSUBS 0.010886f
C748 B.n708 VSUBS 0.025362f
C749 B.n709 VSUBS 0.023944f
C750 B.n710 VSUBS 0.025296f
C751 B.n711 VSUBS 0.010886f
C752 B.n712 VSUBS 0.010886f
C753 B.n713 VSUBS 0.010886f
C754 B.n714 VSUBS 0.010886f
C755 B.n715 VSUBS 0.010886f
C756 B.n716 VSUBS 0.010886f
C757 B.n717 VSUBS 0.010886f
C758 B.n718 VSUBS 0.010886f
C759 B.n719 VSUBS 0.010886f
C760 B.n720 VSUBS 0.010886f
C761 B.n721 VSUBS 0.010886f
C762 B.n722 VSUBS 0.010886f
C763 B.n723 VSUBS 0.010886f
C764 B.n724 VSUBS 0.010886f
C765 B.n725 VSUBS 0.010886f
C766 B.n726 VSUBS 0.010886f
C767 B.n727 VSUBS 0.010886f
C768 B.n728 VSUBS 0.010886f
C769 B.n729 VSUBS 0.010886f
C770 B.n730 VSUBS 0.010886f
C771 B.n731 VSUBS 0.010886f
C772 B.n732 VSUBS 0.010886f
C773 B.n733 VSUBS 0.010886f
C774 B.n734 VSUBS 0.010886f
C775 B.n735 VSUBS 0.010886f
C776 B.n736 VSUBS 0.010886f
C777 B.n737 VSUBS 0.010886f
C778 B.n738 VSUBS 0.010886f
C779 B.n739 VSUBS 0.010886f
C780 B.n740 VSUBS 0.010886f
C781 B.n741 VSUBS 0.010886f
C782 B.n742 VSUBS 0.010886f
C783 B.n743 VSUBS 0.010886f
C784 B.n744 VSUBS 0.010886f
C785 B.n745 VSUBS 0.010886f
C786 B.n746 VSUBS 0.010886f
C787 B.n747 VSUBS 0.010886f
C788 B.n748 VSUBS 0.010886f
C789 B.n749 VSUBS 0.007524f
C790 B.n750 VSUBS 0.025221f
C791 B.n751 VSUBS 0.008805f
C792 B.n752 VSUBS 0.010886f
C793 B.n753 VSUBS 0.010886f
C794 B.n754 VSUBS 0.010886f
C795 B.n755 VSUBS 0.010886f
C796 B.n756 VSUBS 0.010886f
C797 B.n757 VSUBS 0.010886f
C798 B.n758 VSUBS 0.010886f
C799 B.n759 VSUBS 0.010886f
C800 B.n760 VSUBS 0.010886f
C801 B.n761 VSUBS 0.010886f
C802 B.n762 VSUBS 0.010886f
C803 B.n763 VSUBS 0.008805f
C804 B.n764 VSUBS 0.025221f
C805 B.n765 VSUBS 0.007524f
C806 B.n766 VSUBS 0.010886f
C807 B.n767 VSUBS 0.010886f
C808 B.n768 VSUBS 0.010886f
C809 B.n769 VSUBS 0.010886f
C810 B.n770 VSUBS 0.010886f
C811 B.n771 VSUBS 0.010886f
C812 B.n772 VSUBS 0.010886f
C813 B.n773 VSUBS 0.010886f
C814 B.n774 VSUBS 0.010886f
C815 B.n775 VSUBS 0.010886f
C816 B.n776 VSUBS 0.010886f
C817 B.n777 VSUBS 0.010886f
C818 B.n778 VSUBS 0.010886f
C819 B.n779 VSUBS 0.010886f
C820 B.n780 VSUBS 0.010886f
C821 B.n781 VSUBS 0.010886f
C822 B.n782 VSUBS 0.010886f
C823 B.n783 VSUBS 0.010886f
C824 B.n784 VSUBS 0.010886f
C825 B.n785 VSUBS 0.010886f
C826 B.n786 VSUBS 0.010886f
C827 B.n787 VSUBS 0.010886f
C828 B.n788 VSUBS 0.010886f
C829 B.n789 VSUBS 0.010886f
C830 B.n790 VSUBS 0.010886f
C831 B.n791 VSUBS 0.010886f
C832 B.n792 VSUBS 0.010886f
C833 B.n793 VSUBS 0.010886f
C834 B.n794 VSUBS 0.010886f
C835 B.n795 VSUBS 0.010886f
C836 B.n796 VSUBS 0.010886f
C837 B.n797 VSUBS 0.010886f
C838 B.n798 VSUBS 0.010886f
C839 B.n799 VSUBS 0.010886f
C840 B.n800 VSUBS 0.010886f
C841 B.n801 VSUBS 0.010886f
C842 B.n802 VSUBS 0.010886f
C843 B.n803 VSUBS 0.010886f
C844 B.n804 VSUBS 0.025296f
C845 B.n805 VSUBS 0.025296f
C846 B.n806 VSUBS 0.02401f
C847 B.n807 VSUBS 0.010886f
C848 B.n808 VSUBS 0.010886f
C849 B.n809 VSUBS 0.010886f
C850 B.n810 VSUBS 0.010886f
C851 B.n811 VSUBS 0.010886f
C852 B.n812 VSUBS 0.010886f
C853 B.n813 VSUBS 0.010886f
C854 B.n814 VSUBS 0.010886f
C855 B.n815 VSUBS 0.010886f
C856 B.n816 VSUBS 0.010886f
C857 B.n817 VSUBS 0.010886f
C858 B.n818 VSUBS 0.010886f
C859 B.n819 VSUBS 0.010886f
C860 B.n820 VSUBS 0.010886f
C861 B.n821 VSUBS 0.010886f
C862 B.n822 VSUBS 0.010886f
C863 B.n823 VSUBS 0.010886f
C864 B.n824 VSUBS 0.010886f
C865 B.n825 VSUBS 0.010886f
C866 B.n826 VSUBS 0.010886f
C867 B.n827 VSUBS 0.010886f
C868 B.n828 VSUBS 0.010886f
C869 B.n829 VSUBS 0.010886f
C870 B.n830 VSUBS 0.010886f
C871 B.n831 VSUBS 0.010886f
C872 B.n832 VSUBS 0.010886f
C873 B.n833 VSUBS 0.010886f
C874 B.n834 VSUBS 0.010886f
C875 B.n835 VSUBS 0.010886f
C876 B.n836 VSUBS 0.010886f
C877 B.n837 VSUBS 0.010886f
C878 B.n838 VSUBS 0.010886f
C879 B.n839 VSUBS 0.010886f
C880 B.n840 VSUBS 0.010886f
C881 B.n841 VSUBS 0.010886f
C882 B.n842 VSUBS 0.010886f
C883 B.n843 VSUBS 0.010886f
C884 B.n844 VSUBS 0.010886f
C885 B.n845 VSUBS 0.010886f
C886 B.n846 VSUBS 0.010886f
C887 B.n847 VSUBS 0.010886f
C888 B.n848 VSUBS 0.010886f
C889 B.n849 VSUBS 0.010886f
C890 B.n850 VSUBS 0.010886f
C891 B.n851 VSUBS 0.010886f
C892 B.n852 VSUBS 0.010886f
C893 B.n853 VSUBS 0.010886f
C894 B.n854 VSUBS 0.010886f
C895 B.n855 VSUBS 0.010886f
C896 B.n856 VSUBS 0.010886f
C897 B.n857 VSUBS 0.010886f
C898 B.n858 VSUBS 0.010886f
C899 B.n859 VSUBS 0.010886f
C900 B.n860 VSUBS 0.010886f
C901 B.n861 VSUBS 0.010886f
C902 B.n862 VSUBS 0.010886f
C903 B.n863 VSUBS 0.010886f
C904 B.n864 VSUBS 0.010886f
C905 B.n865 VSUBS 0.010886f
C906 B.n866 VSUBS 0.010886f
C907 B.n867 VSUBS 0.010886f
C908 B.n868 VSUBS 0.010886f
C909 B.n869 VSUBS 0.010886f
C910 B.n870 VSUBS 0.010886f
C911 B.n871 VSUBS 0.010886f
C912 B.n872 VSUBS 0.010886f
C913 B.n873 VSUBS 0.010886f
C914 B.n874 VSUBS 0.010886f
C915 B.n875 VSUBS 0.010886f
C916 B.n876 VSUBS 0.010886f
C917 B.n877 VSUBS 0.010886f
C918 B.n878 VSUBS 0.010886f
C919 B.n879 VSUBS 0.010886f
C920 B.n880 VSUBS 0.010886f
C921 B.n881 VSUBS 0.010886f
C922 B.n882 VSUBS 0.010886f
C923 B.n883 VSUBS 0.010886f
C924 B.n884 VSUBS 0.010886f
C925 B.n885 VSUBS 0.010886f
C926 B.n886 VSUBS 0.010886f
C927 B.n887 VSUBS 0.010886f
C928 B.n888 VSUBS 0.010886f
C929 B.n889 VSUBS 0.010886f
C930 B.n890 VSUBS 0.010886f
C931 B.n891 VSUBS 0.010886f
C932 B.n892 VSUBS 0.010886f
C933 B.n893 VSUBS 0.010886f
C934 B.n894 VSUBS 0.010886f
C935 B.n895 VSUBS 0.010886f
C936 B.n896 VSUBS 0.010886f
C937 B.n897 VSUBS 0.010886f
C938 B.n898 VSUBS 0.010886f
C939 B.n899 VSUBS 0.010886f
C940 B.n900 VSUBS 0.010886f
C941 B.n901 VSUBS 0.010886f
C942 B.n902 VSUBS 0.010886f
C943 B.n903 VSUBS 0.010886f
C944 B.n904 VSUBS 0.010886f
C945 B.n905 VSUBS 0.010886f
C946 B.n906 VSUBS 0.010886f
C947 B.n907 VSUBS 0.010886f
C948 B.n908 VSUBS 0.010886f
C949 B.n909 VSUBS 0.010886f
C950 B.n910 VSUBS 0.010886f
C951 B.n911 VSUBS 0.010886f
C952 B.n912 VSUBS 0.010886f
C953 B.n913 VSUBS 0.010886f
C954 B.n914 VSUBS 0.010886f
C955 B.n915 VSUBS 0.010886f
C956 B.n916 VSUBS 0.010886f
C957 B.n917 VSUBS 0.010886f
C958 B.n918 VSUBS 0.010886f
C959 B.n919 VSUBS 0.010886f
C960 B.n920 VSUBS 0.010886f
C961 B.n921 VSUBS 0.010886f
C962 B.n922 VSUBS 0.010886f
C963 B.n923 VSUBS 0.010886f
C964 B.n924 VSUBS 0.010886f
C965 B.n925 VSUBS 0.010886f
C966 B.n926 VSUBS 0.010886f
C967 B.n927 VSUBS 0.010886f
C968 B.n928 VSUBS 0.010886f
C969 B.n929 VSUBS 0.010886f
C970 B.n930 VSUBS 0.010886f
C971 B.n931 VSUBS 0.024649f
C972 VDD2.t4 VSUBS 1.79746f
C973 VDD2.t9 VSUBS 0.188761f
C974 VDD2.t8 VSUBS 0.188761f
C975 VDD2.n0 VSUBS 1.32523f
C976 VDD2.n1 VSUBS 2.08498f
C977 VDD2.t0 VSUBS 0.188761f
C978 VDD2.t2 VSUBS 0.188761f
C979 VDD2.n2 VSUBS 1.36232f
C980 VDD2.n3 VSUBS 4.802259f
C981 VDD2.t5 VSUBS 1.75799f
C982 VDD2.n4 VSUBS 4.74908f
C983 VDD2.t3 VSUBS 0.188761f
C984 VDD2.t1 VSUBS 0.188761f
C985 VDD2.n5 VSUBS 1.32524f
C986 VDD2.n6 VSUBS 1.07422f
C987 VDD2.t6 VSUBS 0.188761f
C988 VDD2.t7 VSUBS 0.188761f
C989 VDD2.n7 VSUBS 1.36226f
C990 VN.n0 VSUBS 0.053627f
C991 VN.t7 VSUBS 2.05455f
C992 VN.n1 VSUBS 0.055265f
C993 VN.n2 VSUBS 0.02851f
C994 VN.n3 VSUBS 0.053135f
C995 VN.n4 VSUBS 0.02851f
C996 VN.t9 VSUBS 2.05455f
C997 VN.n5 VSUBS 0.053135f
C998 VN.n6 VSUBS 0.02851f
C999 VN.n7 VSUBS 0.053135f
C1000 VN.n8 VSUBS 0.02851f
C1001 VN.t1 VSUBS 2.05455f
C1002 VN.n9 VSUBS 0.053135f
C1003 VN.n10 VSUBS 0.02851f
C1004 VN.n11 VSUBS 0.053135f
C1005 VN.n12 VSUBS 0.373751f
C1006 VN.t0 VSUBS 2.05455f
C1007 VN.t5 VSUBS 2.47293f
C1008 VN.n13 VSUBS 0.823005f
C1009 VN.n14 VSUBS 0.848758f
C1010 VN.n15 VSUBS 0.039494f
C1011 VN.n16 VSUBS 0.053135f
C1012 VN.n17 VSUBS 0.02851f
C1013 VN.n18 VSUBS 0.02851f
C1014 VN.n19 VSUBS 0.02851f
C1015 VN.n20 VSUBS 0.051183f
C1016 VN.n21 VSUBS 0.028796f
C1017 VN.n22 VSUBS 0.056394f
C1018 VN.n23 VSUBS 0.02851f
C1019 VN.n24 VSUBS 0.02851f
C1020 VN.n25 VSUBS 0.02851f
C1021 VN.n26 VSUBS 0.053135f
C1022 VN.n27 VSUBS 0.772696f
C1023 VN.n28 VSUBS 0.053135f
C1024 VN.n29 VSUBS 0.02851f
C1025 VN.n30 VSUBS 0.02851f
C1026 VN.n31 VSUBS 0.02851f
C1027 VN.n32 VSUBS 0.056394f
C1028 VN.n33 VSUBS 0.028796f
C1029 VN.n34 VSUBS 0.051183f
C1030 VN.n35 VSUBS 0.02851f
C1031 VN.n36 VSUBS 0.02851f
C1032 VN.n37 VSUBS 0.02851f
C1033 VN.n38 VSUBS 0.053135f
C1034 VN.n39 VSUBS 0.039494f
C1035 VN.n40 VSUBS 0.745794f
C1036 VN.n41 VSUBS 0.040543f
C1037 VN.n42 VSUBS 0.02851f
C1038 VN.n43 VSUBS 0.02851f
C1039 VN.n44 VSUBS 0.02851f
C1040 VN.n45 VSUBS 0.053135f
C1041 VN.n46 VSUBS 0.049972f
C1042 VN.n47 VSUBS 0.031136f
C1043 VN.n48 VSUBS 0.02851f
C1044 VN.n49 VSUBS 0.02851f
C1045 VN.n50 VSUBS 0.02851f
C1046 VN.n51 VSUBS 0.053135f
C1047 VN.n52 VSUBS 0.052086f
C1048 VN.n53 VSUBS 0.876132f
C1049 VN.n54 VSUBS 0.084716f
C1050 VN.n55 VSUBS 0.053627f
C1051 VN.t4 VSUBS 2.05455f
C1052 VN.n56 VSUBS 0.055265f
C1053 VN.n57 VSUBS 0.02851f
C1054 VN.n58 VSUBS 0.053135f
C1055 VN.n59 VSUBS 0.02851f
C1056 VN.t6 VSUBS 2.05455f
C1057 VN.n60 VSUBS 0.053135f
C1058 VN.n61 VSUBS 0.02851f
C1059 VN.n62 VSUBS 0.053135f
C1060 VN.n63 VSUBS 0.02851f
C1061 VN.t8 VSUBS 2.05455f
C1062 VN.n64 VSUBS 0.053135f
C1063 VN.n65 VSUBS 0.02851f
C1064 VN.n66 VSUBS 0.053135f
C1065 VN.n67 VSUBS 0.373751f
C1066 VN.t3 VSUBS 2.05455f
C1067 VN.t2 VSUBS 2.47293f
C1068 VN.n68 VSUBS 0.823005f
C1069 VN.n69 VSUBS 0.848758f
C1070 VN.n70 VSUBS 0.039494f
C1071 VN.n71 VSUBS 0.053135f
C1072 VN.n72 VSUBS 0.02851f
C1073 VN.n73 VSUBS 0.02851f
C1074 VN.n74 VSUBS 0.02851f
C1075 VN.n75 VSUBS 0.051183f
C1076 VN.n76 VSUBS 0.028796f
C1077 VN.n77 VSUBS 0.056394f
C1078 VN.n78 VSUBS 0.02851f
C1079 VN.n79 VSUBS 0.02851f
C1080 VN.n80 VSUBS 0.02851f
C1081 VN.n81 VSUBS 0.053135f
C1082 VN.n82 VSUBS 0.772696f
C1083 VN.n83 VSUBS 0.053135f
C1084 VN.n84 VSUBS 0.02851f
C1085 VN.n85 VSUBS 0.02851f
C1086 VN.n86 VSUBS 0.02851f
C1087 VN.n87 VSUBS 0.056394f
C1088 VN.n88 VSUBS 0.028796f
C1089 VN.n89 VSUBS 0.051183f
C1090 VN.n90 VSUBS 0.02851f
C1091 VN.n91 VSUBS 0.02851f
C1092 VN.n92 VSUBS 0.02851f
C1093 VN.n93 VSUBS 0.053135f
C1094 VN.n94 VSUBS 0.039494f
C1095 VN.n95 VSUBS 0.745794f
C1096 VN.n96 VSUBS 0.040543f
C1097 VN.n97 VSUBS 0.02851f
C1098 VN.n98 VSUBS 0.02851f
C1099 VN.n99 VSUBS 0.02851f
C1100 VN.n100 VSUBS 0.053135f
C1101 VN.n101 VSUBS 0.049972f
C1102 VN.n102 VSUBS 0.031136f
C1103 VN.n103 VSUBS 0.02851f
C1104 VN.n104 VSUBS 0.02851f
C1105 VN.n105 VSUBS 0.02851f
C1106 VN.n106 VSUBS 0.053135f
C1107 VN.n107 VSUBS 0.052086f
C1108 VN.n108 VSUBS 0.876132f
C1109 VN.n109 VSUBS 1.97186f
C1110 VDD1.t0 VSUBS 1.80268f
C1111 VDD1.t2 VSUBS 0.189309f
C1112 VDD1.t3 VSUBS 0.189309f
C1113 VDD1.n0 VSUBS 1.32908f
C1114 VDD1.n1 VSUBS 2.10276f
C1115 VDD1.t8 VSUBS 1.80267f
C1116 VDD1.t7 VSUBS 0.189309f
C1117 VDD1.t1 VSUBS 0.189309f
C1118 VDD1.n2 VSUBS 1.32907f
C1119 VDD1.n3 VSUBS 2.09103f
C1120 VDD1.t4 VSUBS 0.189309f
C1121 VDD1.t9 VSUBS 0.189309f
C1122 VDD1.n4 VSUBS 1.36627f
C1123 VDD1.n5 VSUBS 5.03342f
C1124 VDD1.t5 VSUBS 0.189309f
C1125 VDD1.t6 VSUBS 0.189309f
C1126 VDD1.n6 VSUBS 1.32907f
C1127 VDD1.n7 VSUBS 4.89114f
C1128 VTAIL.t5 VSUBS 0.186325f
C1129 VTAIL.t3 VSUBS 0.186325f
C1130 VTAIL.n0 VSUBS 1.18406f
C1131 VTAIL.n1 VSUBS 1.18971f
C1132 VTAIL.t6 VSUBS 1.60139f
C1133 VTAIL.n2 VSUBS 1.37462f
C1134 VTAIL.t14 VSUBS 0.186325f
C1135 VTAIL.t11 VSUBS 0.186325f
C1136 VTAIL.n3 VSUBS 1.18406f
C1137 VTAIL.n4 VSUBS 1.43307f
C1138 VTAIL.t7 VSUBS 0.186325f
C1139 VTAIL.t8 VSUBS 0.186325f
C1140 VTAIL.n5 VSUBS 1.18406f
C1141 VTAIL.n6 VSUBS 2.95343f
C1142 VTAIL.t1 VSUBS 0.186325f
C1143 VTAIL.t4 VSUBS 0.186325f
C1144 VTAIL.n7 VSUBS 1.18408f
C1145 VTAIL.n8 VSUBS 2.95342f
C1146 VTAIL.t17 VSUBS 0.186325f
C1147 VTAIL.t2 VSUBS 0.186325f
C1148 VTAIL.n9 VSUBS 1.18408f
C1149 VTAIL.n10 VSUBS 1.43306f
C1150 VTAIL.t0 VSUBS 1.6014f
C1151 VTAIL.n11 VSUBS 1.3746f
C1152 VTAIL.t15 VSUBS 0.186325f
C1153 VTAIL.t13 VSUBS 0.186325f
C1154 VTAIL.n12 VSUBS 1.18408f
C1155 VTAIL.n13 VSUBS 1.28377f
C1156 VTAIL.t12 VSUBS 0.186325f
C1157 VTAIL.t10 VSUBS 0.186325f
C1158 VTAIL.n14 VSUBS 1.18408f
C1159 VTAIL.n15 VSUBS 1.43306f
C1160 VTAIL.t9 VSUBS 1.60139f
C1161 VTAIL.n16 VSUBS 2.64238f
C1162 VTAIL.t19 VSUBS 1.60139f
C1163 VTAIL.n17 VSUBS 2.64238f
C1164 VTAIL.t16 VSUBS 0.186325f
C1165 VTAIL.t18 VSUBS 0.186325f
C1166 VTAIL.n18 VSUBS 1.18406f
C1167 VTAIL.n19 VSUBS 1.12526f
C1168 VP.n0 VSUBS 0.059899f
C1169 VP.t0 VSUBS 2.29487f
C1170 VP.n1 VSUBS 0.061729f
C1171 VP.n2 VSUBS 0.031844f
C1172 VP.n3 VSUBS 0.05935f
C1173 VP.n4 VSUBS 0.031844f
C1174 VP.t5 VSUBS 2.29487f
C1175 VP.n5 VSUBS 0.05935f
C1176 VP.n6 VSUBS 0.031844f
C1177 VP.n7 VSUBS 0.05935f
C1178 VP.n8 VSUBS 0.031844f
C1179 VP.t8 VSUBS 2.29487f
C1180 VP.n9 VSUBS 0.05935f
C1181 VP.n10 VSUBS 0.031844f
C1182 VP.n11 VSUBS 0.05935f
C1183 VP.n12 VSUBS 0.031844f
C1184 VP.t2 VSUBS 2.29487f
C1185 VP.n13 VSUBS 0.05935f
C1186 VP.n14 VSUBS 0.031844f
C1187 VP.n15 VSUBS 0.061729f
C1188 VP.n16 VSUBS 0.059899f
C1189 VP.t1 VSUBS 2.29487f
C1190 VP.n17 VSUBS 0.059899f
C1191 VP.t3 VSUBS 2.29487f
C1192 VP.n18 VSUBS 0.061729f
C1193 VP.n19 VSUBS 0.031844f
C1194 VP.n20 VSUBS 0.05935f
C1195 VP.n21 VSUBS 0.031844f
C1196 VP.t4 VSUBS 2.29487f
C1197 VP.n22 VSUBS 0.05935f
C1198 VP.n23 VSUBS 0.031844f
C1199 VP.n24 VSUBS 0.05935f
C1200 VP.n25 VSUBS 0.031844f
C1201 VP.t6 VSUBS 2.29487f
C1202 VP.n26 VSUBS 0.05935f
C1203 VP.n27 VSUBS 0.031844f
C1204 VP.n28 VSUBS 0.05935f
C1205 VP.n29 VSUBS 0.417469f
C1206 VP.t7 VSUBS 2.29487f
C1207 VP.t9 VSUBS 2.76218f
C1208 VP.n30 VSUBS 0.919273f
C1209 VP.n31 VSUBS 0.948035f
C1210 VP.n32 VSUBS 0.044113f
C1211 VP.n33 VSUBS 0.05935f
C1212 VP.n34 VSUBS 0.031844f
C1213 VP.n35 VSUBS 0.031844f
C1214 VP.n36 VSUBS 0.031844f
C1215 VP.n37 VSUBS 0.05717f
C1216 VP.n38 VSUBS 0.032165f
C1217 VP.n39 VSUBS 0.06299f
C1218 VP.n40 VSUBS 0.031844f
C1219 VP.n41 VSUBS 0.031844f
C1220 VP.n42 VSUBS 0.031844f
C1221 VP.n43 VSUBS 0.05935f
C1222 VP.n44 VSUBS 0.863077f
C1223 VP.n45 VSUBS 0.05935f
C1224 VP.n46 VSUBS 0.031844f
C1225 VP.n47 VSUBS 0.031844f
C1226 VP.n48 VSUBS 0.031844f
C1227 VP.n49 VSUBS 0.06299f
C1228 VP.n50 VSUBS 0.032165f
C1229 VP.n51 VSUBS 0.05717f
C1230 VP.n52 VSUBS 0.031844f
C1231 VP.n53 VSUBS 0.031844f
C1232 VP.n54 VSUBS 0.031844f
C1233 VP.n55 VSUBS 0.05935f
C1234 VP.n56 VSUBS 0.044113f
C1235 VP.n57 VSUBS 0.833028f
C1236 VP.n58 VSUBS 0.045285f
C1237 VP.n59 VSUBS 0.031844f
C1238 VP.n60 VSUBS 0.031844f
C1239 VP.n61 VSUBS 0.031844f
C1240 VP.n62 VSUBS 0.05935f
C1241 VP.n63 VSUBS 0.055817f
C1242 VP.n64 VSUBS 0.034778f
C1243 VP.n65 VSUBS 0.031844f
C1244 VP.n66 VSUBS 0.031844f
C1245 VP.n67 VSUBS 0.031844f
C1246 VP.n68 VSUBS 0.05935f
C1247 VP.n69 VSUBS 0.058178f
C1248 VP.n70 VSUBS 0.978611f
C1249 VP.n71 VSUBS 2.19492f
C1250 VP.n72 VSUBS 2.21513f
C1251 VP.n73 VSUBS 0.978611f
C1252 VP.n74 VSUBS 0.058178f
C1253 VP.n75 VSUBS 0.05935f
C1254 VP.n76 VSUBS 0.031844f
C1255 VP.n77 VSUBS 0.031844f
C1256 VP.n78 VSUBS 0.031844f
C1257 VP.n79 VSUBS 0.034778f
C1258 VP.n80 VSUBS 0.055817f
C1259 VP.n81 VSUBS 0.05935f
C1260 VP.n82 VSUBS 0.031844f
C1261 VP.n83 VSUBS 0.031844f
C1262 VP.n84 VSUBS 0.031844f
C1263 VP.n85 VSUBS 0.045285f
C1264 VP.n86 VSUBS 0.833028f
C1265 VP.n87 VSUBS 0.044113f
C1266 VP.n88 VSUBS 0.05935f
C1267 VP.n89 VSUBS 0.031844f
C1268 VP.n90 VSUBS 0.031844f
C1269 VP.n91 VSUBS 0.031844f
C1270 VP.n92 VSUBS 0.05717f
C1271 VP.n93 VSUBS 0.032165f
C1272 VP.n94 VSUBS 0.06299f
C1273 VP.n95 VSUBS 0.031844f
C1274 VP.n96 VSUBS 0.031844f
C1275 VP.n97 VSUBS 0.031844f
C1276 VP.n98 VSUBS 0.05935f
C1277 VP.n99 VSUBS 0.863077f
C1278 VP.n100 VSUBS 0.05935f
C1279 VP.n101 VSUBS 0.031844f
C1280 VP.n102 VSUBS 0.031844f
C1281 VP.n103 VSUBS 0.031844f
C1282 VP.n104 VSUBS 0.06299f
C1283 VP.n105 VSUBS 0.032165f
C1284 VP.n106 VSUBS 0.05717f
C1285 VP.n107 VSUBS 0.031844f
C1286 VP.n108 VSUBS 0.031844f
C1287 VP.n109 VSUBS 0.031844f
C1288 VP.n110 VSUBS 0.05935f
C1289 VP.n111 VSUBS 0.044113f
C1290 VP.n112 VSUBS 0.833028f
C1291 VP.n113 VSUBS 0.045285f
C1292 VP.n114 VSUBS 0.031844f
C1293 VP.n115 VSUBS 0.031844f
C1294 VP.n116 VSUBS 0.031844f
C1295 VP.n117 VSUBS 0.05935f
C1296 VP.n118 VSUBS 0.055817f
C1297 VP.n119 VSUBS 0.034778f
C1298 VP.n120 VSUBS 0.031844f
C1299 VP.n121 VSUBS 0.031844f
C1300 VP.n122 VSUBS 0.031844f
C1301 VP.n123 VSUBS 0.05935f
C1302 VP.n124 VSUBS 0.058178f
C1303 VP.n125 VSUBS 0.978611f
C1304 VP.n126 VSUBS 0.094625f
.ends

