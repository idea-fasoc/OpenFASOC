* NGSPICE file created from diff_pair_sample_1320.ext - technology: sky130A

.subckt diff_pair_sample_1320 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VP.t0 VDD1.t5 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X1 VDD1.t4 VP.t1 VTAIL.t16 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=2.6334 ps=16.29 w=15.96 l=3.61
X2 B.t11 B.t9 B.t10 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=0 ps=0 w=15.96 l=3.61
X3 B.t8 B.t6 B.t7 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=0 ps=0 w=15.96 l=3.61
X4 VDD2.t9 VN.t0 VTAIL.t19 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=6.2244 ps=32.7 w=15.96 l=3.61
X5 VTAIL.t5 VN.t1 VDD2.t8 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X6 VDD2.t7 VN.t2 VTAIL.t2 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X7 VDD1.t3 VP.t2 VTAIL.t15 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=2.6334 ps=16.29 w=15.96 l=3.61
X8 VDD1.t2 VP.t3 VTAIL.t14 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=6.2244 ps=32.7 w=15.96 l=3.61
X9 VDD1.t1 VP.t4 VTAIL.t13 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=6.2244 ps=32.7 w=15.96 l=3.61
X10 VTAIL.t12 VP.t5 VDD1.t0 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X11 VDD2.t6 VN.t3 VTAIL.t1 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=6.2244 ps=32.7 w=15.96 l=3.61
X12 B.t5 B.t3 B.t4 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=0 ps=0 w=15.96 l=3.61
X13 VTAIL.t11 VP.t6 VDD1.t7 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X14 VDD1.t6 VP.t7 VTAIL.t10 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X15 VTAIL.t9 VP.t8 VDD1.t9 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X16 VDD2.t5 VN.t4 VTAIL.t4 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X17 VDD1.t8 VP.t9 VTAIL.t8 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X18 VDD2.t4 VN.t5 VTAIL.t0 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=2.6334 ps=16.29 w=15.96 l=3.61
X19 VTAIL.t6 VN.t6 VDD2.t3 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X20 VDD2.t2 VN.t7 VTAIL.t18 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=2.6334 ps=16.29 w=15.96 l=3.61
X21 B.t2 B.t0 B.t1 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=6.2244 pd=32.7 as=0 ps=0 w=15.96 l=3.61
X22 VTAIL.t3 VN.t8 VDD2.t1 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
X23 VTAIL.t7 VN.t9 VDD2.t0 w_n5698_n4160# sky130_fd_pr__pfet_01v8 ad=2.6334 pd=16.29 as=2.6334 ps=16.29 w=15.96 l=3.61
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n57 VP.n56 161.3
R16 VP.n58 VP.n21 161.3
R17 VP.n60 VP.n59 161.3
R18 VP.n61 VP.n20 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n64 VP.n19 161.3
R21 VP.n66 VP.n65 161.3
R22 VP.n67 VP.n18 161.3
R23 VP.n69 VP.n68 161.3
R24 VP.n123 VP.n122 161.3
R25 VP.n121 VP.n1 161.3
R26 VP.n120 VP.n119 161.3
R27 VP.n118 VP.n2 161.3
R28 VP.n117 VP.n116 161.3
R29 VP.n115 VP.n3 161.3
R30 VP.n114 VP.n113 161.3
R31 VP.n112 VP.n4 161.3
R32 VP.n111 VP.n110 161.3
R33 VP.n108 VP.n5 161.3
R34 VP.n107 VP.n106 161.3
R35 VP.n105 VP.n6 161.3
R36 VP.n104 VP.n103 161.3
R37 VP.n102 VP.n7 161.3
R38 VP.n101 VP.n100 161.3
R39 VP.n99 VP.n8 161.3
R40 VP.n98 VP.n97 161.3
R41 VP.n95 VP.n9 161.3
R42 VP.n94 VP.n93 161.3
R43 VP.n92 VP.n10 161.3
R44 VP.n91 VP.n90 161.3
R45 VP.n89 VP.n11 161.3
R46 VP.n88 VP.n87 161.3
R47 VP.n86 VP.n12 161.3
R48 VP.n85 VP.n84 161.3
R49 VP.n82 VP.n13 161.3
R50 VP.n81 VP.n80 161.3
R51 VP.n79 VP.n14 161.3
R52 VP.n78 VP.n77 161.3
R53 VP.n76 VP.n15 161.3
R54 VP.n75 VP.n74 161.3
R55 VP.n73 VP.n16 161.3
R56 VP.n31 VP.t1 139.361
R57 VP.n71 VP.t2 106.547
R58 VP.n83 VP.t8 106.547
R59 VP.n96 VP.t7 106.547
R60 VP.n109 VP.t5 106.547
R61 VP.n0 VP.t3 106.547
R62 VP.n17 VP.t4 106.547
R63 VP.n55 VP.t0 106.547
R64 VP.n42 VP.t9 106.547
R65 VP.n30 VP.t6 106.547
R66 VP.n72 VP.n71 83.8517
R67 VP.n124 VP.n0 83.8517
R68 VP.n70 VP.n17 83.8517
R69 VP.n31 VP.n30 65.3998
R70 VP.n72 VP.n70 61.6662
R71 VP.n90 VP.n10 56.5617
R72 VP.n103 VP.n6 56.5617
R73 VP.n49 VP.n23 56.5617
R74 VP.n36 VP.n27 56.5617
R75 VP.n77 VP.n14 56.0773
R76 VP.n116 VP.n2 56.0773
R77 VP.n62 VP.n19 56.0773
R78 VP.n81 VP.n14 25.0767
R79 VP.n116 VP.n115 25.0767
R80 VP.n62 VP.n61 25.0767
R81 VP.n75 VP.n16 24.5923
R82 VP.n76 VP.n75 24.5923
R83 VP.n77 VP.n76 24.5923
R84 VP.n82 VP.n81 24.5923
R85 VP.n84 VP.n82 24.5923
R86 VP.n88 VP.n12 24.5923
R87 VP.n89 VP.n88 24.5923
R88 VP.n90 VP.n89 24.5923
R89 VP.n94 VP.n10 24.5923
R90 VP.n95 VP.n94 24.5923
R91 VP.n97 VP.n95 24.5923
R92 VP.n101 VP.n8 24.5923
R93 VP.n102 VP.n101 24.5923
R94 VP.n103 VP.n102 24.5923
R95 VP.n107 VP.n6 24.5923
R96 VP.n108 VP.n107 24.5923
R97 VP.n110 VP.n108 24.5923
R98 VP.n114 VP.n4 24.5923
R99 VP.n115 VP.n114 24.5923
R100 VP.n120 VP.n2 24.5923
R101 VP.n121 VP.n120 24.5923
R102 VP.n122 VP.n121 24.5923
R103 VP.n66 VP.n19 24.5923
R104 VP.n67 VP.n66 24.5923
R105 VP.n68 VP.n67 24.5923
R106 VP.n53 VP.n23 24.5923
R107 VP.n54 VP.n53 24.5923
R108 VP.n56 VP.n54 24.5923
R109 VP.n60 VP.n21 24.5923
R110 VP.n61 VP.n60 24.5923
R111 VP.n40 VP.n27 24.5923
R112 VP.n41 VP.n40 24.5923
R113 VP.n43 VP.n41 24.5923
R114 VP.n47 VP.n25 24.5923
R115 VP.n48 VP.n47 24.5923
R116 VP.n49 VP.n48 24.5923
R117 VP.n34 VP.n29 24.5923
R118 VP.n35 VP.n34 24.5923
R119 VP.n36 VP.n35 24.5923
R120 VP.n84 VP.n83 15.2474
R121 VP.n109 VP.n4 15.2474
R122 VP.n55 VP.n21 15.2474
R123 VP.n97 VP.n96 12.2964
R124 VP.n96 VP.n8 12.2964
R125 VP.n43 VP.n42 12.2964
R126 VP.n42 VP.n25 12.2964
R127 VP.n83 VP.n12 9.3454
R128 VP.n110 VP.n109 9.3454
R129 VP.n56 VP.n55 9.3454
R130 VP.n30 VP.n29 9.3454
R131 VP.n71 VP.n16 6.39438
R132 VP.n122 VP.n0 6.39438
R133 VP.n68 VP.n17 6.39438
R134 VP.n32 VP.n31 3.26188
R135 VP.n70 VP.n69 0.354861
R136 VP.n73 VP.n72 0.354861
R137 VP.n124 VP.n123 0.354861
R138 VP VP.n124 0.267071
R139 VP.n33 VP.n32 0.189894
R140 VP.n33 VP.n28 0.189894
R141 VP.n37 VP.n28 0.189894
R142 VP.n38 VP.n37 0.189894
R143 VP.n39 VP.n38 0.189894
R144 VP.n39 VP.n26 0.189894
R145 VP.n44 VP.n26 0.189894
R146 VP.n45 VP.n44 0.189894
R147 VP.n46 VP.n45 0.189894
R148 VP.n46 VP.n24 0.189894
R149 VP.n50 VP.n24 0.189894
R150 VP.n51 VP.n50 0.189894
R151 VP.n52 VP.n51 0.189894
R152 VP.n52 VP.n22 0.189894
R153 VP.n57 VP.n22 0.189894
R154 VP.n58 VP.n57 0.189894
R155 VP.n59 VP.n58 0.189894
R156 VP.n59 VP.n20 0.189894
R157 VP.n63 VP.n20 0.189894
R158 VP.n64 VP.n63 0.189894
R159 VP.n65 VP.n64 0.189894
R160 VP.n65 VP.n18 0.189894
R161 VP.n69 VP.n18 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n74 VP.n15 0.189894
R164 VP.n78 VP.n15 0.189894
R165 VP.n79 VP.n78 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n80 VP.n13 0.189894
R168 VP.n85 VP.n13 0.189894
R169 VP.n86 VP.n85 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n87 VP.n11 0.189894
R172 VP.n91 VP.n11 0.189894
R173 VP.n92 VP.n91 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n93 VP.n9 0.189894
R176 VP.n98 VP.n9 0.189894
R177 VP.n99 VP.n98 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n100 VP.n7 0.189894
R180 VP.n104 VP.n7 0.189894
R181 VP.n105 VP.n104 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n106 VP.n5 0.189894
R184 VP.n111 VP.n5 0.189894
R185 VP.n112 VP.n111 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n113 VP.n3 0.189894
R188 VP.n117 VP.n3 0.189894
R189 VP.n118 VP.n117 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n119 VP.n1 0.189894
R192 VP.n123 VP.n1 0.189894
R193 VDD1.n1 VDD1.t4 73.4068
R194 VDD1.n3 VDD1.t3 73.4065
R195 VDD1.n5 VDD1.n4 70.4654
R196 VDD1.n7 VDD1.n6 67.9736
R197 VDD1.n1 VDD1.n0 67.9736
R198 VDD1.n3 VDD1.n2 67.9733
R199 VDD1.n7 VDD1.n5 55.8888
R200 VDD1 VDD1.n7 2.48972
R201 VDD1.n6 VDD1.t5 2.03715
R202 VDD1.n6 VDD1.t1 2.03715
R203 VDD1.n0 VDD1.t7 2.03715
R204 VDD1.n0 VDD1.t8 2.03715
R205 VDD1.n4 VDD1.t0 2.03715
R206 VDD1.n4 VDD1.t2 2.03715
R207 VDD1.n2 VDD1.t9 2.03715
R208 VDD1.n2 VDD1.t6 2.03715
R209 VDD1 VDD1.n1 0.907828
R210 VDD1.n5 VDD1.n3 0.794292
R211 VTAIL.n11 VTAIL.t1 53.3314
R212 VTAIL.n16 VTAIL.t13 53.3314
R213 VTAIL.n17 VTAIL.t19 53.3312
R214 VTAIL.n2 VTAIL.t14 53.3312
R215 VTAIL.n15 VTAIL.n14 51.2948
R216 VTAIL.n13 VTAIL.n12 51.2948
R217 VTAIL.n10 VTAIL.n9 51.2948
R218 VTAIL.n8 VTAIL.n7 51.2948
R219 VTAIL.n19 VTAIL.n18 51.2945
R220 VTAIL.n1 VTAIL.n0 51.2945
R221 VTAIL.n4 VTAIL.n3 51.2945
R222 VTAIL.n6 VTAIL.n5 51.2945
R223 VTAIL.n8 VTAIL.n6 32.9186
R224 VTAIL.n17 VTAIL.n16 29.5221
R225 VTAIL.n10 VTAIL.n8 3.39705
R226 VTAIL.n11 VTAIL.n10 3.39705
R227 VTAIL.n15 VTAIL.n13 3.39705
R228 VTAIL.n16 VTAIL.n15 3.39705
R229 VTAIL.n6 VTAIL.n4 3.39705
R230 VTAIL.n4 VTAIL.n2 3.39705
R231 VTAIL.n19 VTAIL.n17 3.39705
R232 VTAIL VTAIL.n1 2.6061
R233 VTAIL.n13 VTAIL.n11 2.1686
R234 VTAIL.n2 VTAIL.n1 2.1686
R235 VTAIL.n18 VTAIL.t2 2.03715
R236 VTAIL.n18 VTAIL.t5 2.03715
R237 VTAIL.n0 VTAIL.t0 2.03715
R238 VTAIL.n0 VTAIL.t3 2.03715
R239 VTAIL.n3 VTAIL.t10 2.03715
R240 VTAIL.n3 VTAIL.t12 2.03715
R241 VTAIL.n5 VTAIL.t15 2.03715
R242 VTAIL.n5 VTAIL.t9 2.03715
R243 VTAIL.n14 VTAIL.t8 2.03715
R244 VTAIL.n14 VTAIL.t17 2.03715
R245 VTAIL.n12 VTAIL.t16 2.03715
R246 VTAIL.n12 VTAIL.t11 2.03715
R247 VTAIL.n9 VTAIL.t4 2.03715
R248 VTAIL.n9 VTAIL.t7 2.03715
R249 VTAIL.n7 VTAIL.t18 2.03715
R250 VTAIL.n7 VTAIL.t6 2.03715
R251 VTAIL VTAIL.n19 0.791448
R252 B.n570 B.n181 585
R253 B.n569 B.n568 585
R254 B.n567 B.n182 585
R255 B.n566 B.n565 585
R256 B.n564 B.n183 585
R257 B.n563 B.n562 585
R258 B.n561 B.n184 585
R259 B.n560 B.n559 585
R260 B.n558 B.n185 585
R261 B.n557 B.n556 585
R262 B.n555 B.n186 585
R263 B.n554 B.n553 585
R264 B.n552 B.n187 585
R265 B.n551 B.n550 585
R266 B.n549 B.n188 585
R267 B.n548 B.n547 585
R268 B.n546 B.n189 585
R269 B.n545 B.n544 585
R270 B.n543 B.n190 585
R271 B.n542 B.n541 585
R272 B.n540 B.n191 585
R273 B.n539 B.n538 585
R274 B.n537 B.n192 585
R275 B.n536 B.n535 585
R276 B.n534 B.n193 585
R277 B.n533 B.n532 585
R278 B.n531 B.n194 585
R279 B.n530 B.n529 585
R280 B.n528 B.n195 585
R281 B.n527 B.n526 585
R282 B.n525 B.n196 585
R283 B.n524 B.n523 585
R284 B.n522 B.n197 585
R285 B.n521 B.n520 585
R286 B.n519 B.n198 585
R287 B.n518 B.n517 585
R288 B.n516 B.n199 585
R289 B.n515 B.n514 585
R290 B.n513 B.n200 585
R291 B.n512 B.n511 585
R292 B.n510 B.n201 585
R293 B.n509 B.n508 585
R294 B.n507 B.n202 585
R295 B.n506 B.n505 585
R296 B.n504 B.n203 585
R297 B.n503 B.n502 585
R298 B.n501 B.n204 585
R299 B.n500 B.n499 585
R300 B.n498 B.n205 585
R301 B.n497 B.n496 585
R302 B.n495 B.n206 585
R303 B.n494 B.n493 585
R304 B.n492 B.n207 585
R305 B.n490 B.n489 585
R306 B.n488 B.n210 585
R307 B.n487 B.n486 585
R308 B.n485 B.n211 585
R309 B.n484 B.n483 585
R310 B.n482 B.n212 585
R311 B.n481 B.n480 585
R312 B.n479 B.n213 585
R313 B.n478 B.n477 585
R314 B.n476 B.n214 585
R315 B.n475 B.n474 585
R316 B.n470 B.n215 585
R317 B.n469 B.n468 585
R318 B.n467 B.n216 585
R319 B.n466 B.n465 585
R320 B.n464 B.n217 585
R321 B.n463 B.n462 585
R322 B.n461 B.n218 585
R323 B.n460 B.n459 585
R324 B.n458 B.n219 585
R325 B.n457 B.n456 585
R326 B.n455 B.n220 585
R327 B.n454 B.n453 585
R328 B.n452 B.n221 585
R329 B.n451 B.n450 585
R330 B.n449 B.n222 585
R331 B.n448 B.n447 585
R332 B.n446 B.n223 585
R333 B.n445 B.n444 585
R334 B.n443 B.n224 585
R335 B.n442 B.n441 585
R336 B.n440 B.n225 585
R337 B.n439 B.n438 585
R338 B.n437 B.n226 585
R339 B.n436 B.n435 585
R340 B.n434 B.n227 585
R341 B.n433 B.n432 585
R342 B.n431 B.n228 585
R343 B.n430 B.n429 585
R344 B.n428 B.n229 585
R345 B.n427 B.n426 585
R346 B.n425 B.n230 585
R347 B.n424 B.n423 585
R348 B.n422 B.n231 585
R349 B.n421 B.n420 585
R350 B.n419 B.n232 585
R351 B.n418 B.n417 585
R352 B.n416 B.n233 585
R353 B.n415 B.n414 585
R354 B.n413 B.n234 585
R355 B.n412 B.n411 585
R356 B.n410 B.n235 585
R357 B.n409 B.n408 585
R358 B.n407 B.n236 585
R359 B.n406 B.n405 585
R360 B.n404 B.n237 585
R361 B.n403 B.n402 585
R362 B.n401 B.n238 585
R363 B.n400 B.n399 585
R364 B.n398 B.n239 585
R365 B.n397 B.n396 585
R366 B.n395 B.n240 585
R367 B.n394 B.n393 585
R368 B.n572 B.n571 585
R369 B.n573 B.n180 585
R370 B.n575 B.n574 585
R371 B.n576 B.n179 585
R372 B.n578 B.n577 585
R373 B.n579 B.n178 585
R374 B.n581 B.n580 585
R375 B.n582 B.n177 585
R376 B.n584 B.n583 585
R377 B.n585 B.n176 585
R378 B.n587 B.n586 585
R379 B.n588 B.n175 585
R380 B.n590 B.n589 585
R381 B.n591 B.n174 585
R382 B.n593 B.n592 585
R383 B.n594 B.n173 585
R384 B.n596 B.n595 585
R385 B.n597 B.n172 585
R386 B.n599 B.n598 585
R387 B.n600 B.n171 585
R388 B.n602 B.n601 585
R389 B.n603 B.n170 585
R390 B.n605 B.n604 585
R391 B.n606 B.n169 585
R392 B.n608 B.n607 585
R393 B.n609 B.n168 585
R394 B.n611 B.n610 585
R395 B.n612 B.n167 585
R396 B.n614 B.n613 585
R397 B.n615 B.n166 585
R398 B.n617 B.n616 585
R399 B.n618 B.n165 585
R400 B.n620 B.n619 585
R401 B.n621 B.n164 585
R402 B.n623 B.n622 585
R403 B.n624 B.n163 585
R404 B.n626 B.n625 585
R405 B.n627 B.n162 585
R406 B.n629 B.n628 585
R407 B.n630 B.n161 585
R408 B.n632 B.n631 585
R409 B.n633 B.n160 585
R410 B.n635 B.n634 585
R411 B.n636 B.n159 585
R412 B.n638 B.n637 585
R413 B.n639 B.n158 585
R414 B.n641 B.n640 585
R415 B.n642 B.n157 585
R416 B.n644 B.n643 585
R417 B.n645 B.n156 585
R418 B.n647 B.n646 585
R419 B.n648 B.n155 585
R420 B.n650 B.n649 585
R421 B.n651 B.n154 585
R422 B.n653 B.n652 585
R423 B.n654 B.n153 585
R424 B.n656 B.n655 585
R425 B.n657 B.n152 585
R426 B.n659 B.n658 585
R427 B.n660 B.n151 585
R428 B.n662 B.n661 585
R429 B.n663 B.n150 585
R430 B.n665 B.n664 585
R431 B.n666 B.n149 585
R432 B.n668 B.n667 585
R433 B.n669 B.n148 585
R434 B.n671 B.n670 585
R435 B.n672 B.n147 585
R436 B.n674 B.n673 585
R437 B.n675 B.n146 585
R438 B.n677 B.n676 585
R439 B.n678 B.n145 585
R440 B.n680 B.n679 585
R441 B.n681 B.n144 585
R442 B.n683 B.n682 585
R443 B.n684 B.n143 585
R444 B.n686 B.n685 585
R445 B.n687 B.n142 585
R446 B.n689 B.n688 585
R447 B.n690 B.n141 585
R448 B.n692 B.n691 585
R449 B.n693 B.n140 585
R450 B.n695 B.n694 585
R451 B.n696 B.n139 585
R452 B.n698 B.n697 585
R453 B.n699 B.n138 585
R454 B.n701 B.n700 585
R455 B.n702 B.n137 585
R456 B.n704 B.n703 585
R457 B.n705 B.n136 585
R458 B.n707 B.n706 585
R459 B.n708 B.n135 585
R460 B.n710 B.n709 585
R461 B.n711 B.n134 585
R462 B.n713 B.n712 585
R463 B.n714 B.n133 585
R464 B.n716 B.n715 585
R465 B.n717 B.n132 585
R466 B.n719 B.n718 585
R467 B.n720 B.n131 585
R468 B.n722 B.n721 585
R469 B.n723 B.n130 585
R470 B.n725 B.n724 585
R471 B.n726 B.n129 585
R472 B.n728 B.n727 585
R473 B.n729 B.n128 585
R474 B.n731 B.n730 585
R475 B.n732 B.n127 585
R476 B.n734 B.n733 585
R477 B.n735 B.n126 585
R478 B.n737 B.n736 585
R479 B.n738 B.n125 585
R480 B.n740 B.n739 585
R481 B.n741 B.n124 585
R482 B.n743 B.n742 585
R483 B.n744 B.n123 585
R484 B.n746 B.n745 585
R485 B.n747 B.n122 585
R486 B.n749 B.n748 585
R487 B.n750 B.n121 585
R488 B.n752 B.n751 585
R489 B.n753 B.n120 585
R490 B.n755 B.n754 585
R491 B.n756 B.n119 585
R492 B.n758 B.n757 585
R493 B.n759 B.n118 585
R494 B.n761 B.n760 585
R495 B.n762 B.n117 585
R496 B.n764 B.n763 585
R497 B.n765 B.n116 585
R498 B.n767 B.n766 585
R499 B.n768 B.n115 585
R500 B.n770 B.n769 585
R501 B.n771 B.n114 585
R502 B.n773 B.n772 585
R503 B.n774 B.n113 585
R504 B.n776 B.n775 585
R505 B.n777 B.n112 585
R506 B.n779 B.n778 585
R507 B.n780 B.n111 585
R508 B.n782 B.n781 585
R509 B.n783 B.n110 585
R510 B.n785 B.n784 585
R511 B.n786 B.n109 585
R512 B.n788 B.n787 585
R513 B.n789 B.n108 585
R514 B.n791 B.n790 585
R515 B.n792 B.n107 585
R516 B.n794 B.n793 585
R517 B.n795 B.n106 585
R518 B.n797 B.n796 585
R519 B.n798 B.n105 585
R520 B.n800 B.n799 585
R521 B.n801 B.n104 585
R522 B.n803 B.n802 585
R523 B.n804 B.n103 585
R524 B.n980 B.n979 585
R525 B.n978 B.n41 585
R526 B.n977 B.n976 585
R527 B.n975 B.n42 585
R528 B.n974 B.n973 585
R529 B.n972 B.n43 585
R530 B.n971 B.n970 585
R531 B.n969 B.n44 585
R532 B.n968 B.n967 585
R533 B.n966 B.n45 585
R534 B.n965 B.n964 585
R535 B.n963 B.n46 585
R536 B.n962 B.n961 585
R537 B.n960 B.n47 585
R538 B.n959 B.n958 585
R539 B.n957 B.n48 585
R540 B.n956 B.n955 585
R541 B.n954 B.n49 585
R542 B.n953 B.n952 585
R543 B.n951 B.n50 585
R544 B.n950 B.n949 585
R545 B.n948 B.n51 585
R546 B.n947 B.n946 585
R547 B.n945 B.n52 585
R548 B.n944 B.n943 585
R549 B.n942 B.n53 585
R550 B.n941 B.n940 585
R551 B.n939 B.n54 585
R552 B.n938 B.n937 585
R553 B.n936 B.n55 585
R554 B.n935 B.n934 585
R555 B.n933 B.n56 585
R556 B.n932 B.n931 585
R557 B.n930 B.n57 585
R558 B.n929 B.n928 585
R559 B.n927 B.n58 585
R560 B.n926 B.n925 585
R561 B.n924 B.n59 585
R562 B.n923 B.n922 585
R563 B.n921 B.n60 585
R564 B.n920 B.n919 585
R565 B.n918 B.n61 585
R566 B.n917 B.n916 585
R567 B.n915 B.n62 585
R568 B.n914 B.n913 585
R569 B.n912 B.n63 585
R570 B.n911 B.n910 585
R571 B.n909 B.n64 585
R572 B.n908 B.n907 585
R573 B.n906 B.n65 585
R574 B.n905 B.n904 585
R575 B.n903 B.n66 585
R576 B.n902 B.n901 585
R577 B.n899 B.n67 585
R578 B.n898 B.n897 585
R579 B.n896 B.n70 585
R580 B.n895 B.n894 585
R581 B.n893 B.n71 585
R582 B.n892 B.n891 585
R583 B.n890 B.n72 585
R584 B.n889 B.n888 585
R585 B.n887 B.n73 585
R586 B.n886 B.n885 585
R587 B.n884 B.n883 585
R588 B.n882 B.n77 585
R589 B.n881 B.n880 585
R590 B.n879 B.n78 585
R591 B.n878 B.n877 585
R592 B.n876 B.n79 585
R593 B.n875 B.n874 585
R594 B.n873 B.n80 585
R595 B.n872 B.n871 585
R596 B.n870 B.n81 585
R597 B.n869 B.n868 585
R598 B.n867 B.n82 585
R599 B.n866 B.n865 585
R600 B.n864 B.n83 585
R601 B.n863 B.n862 585
R602 B.n861 B.n84 585
R603 B.n860 B.n859 585
R604 B.n858 B.n85 585
R605 B.n857 B.n856 585
R606 B.n855 B.n86 585
R607 B.n854 B.n853 585
R608 B.n852 B.n87 585
R609 B.n851 B.n850 585
R610 B.n849 B.n88 585
R611 B.n848 B.n847 585
R612 B.n846 B.n89 585
R613 B.n845 B.n844 585
R614 B.n843 B.n90 585
R615 B.n842 B.n841 585
R616 B.n840 B.n91 585
R617 B.n839 B.n838 585
R618 B.n837 B.n92 585
R619 B.n836 B.n835 585
R620 B.n834 B.n93 585
R621 B.n833 B.n832 585
R622 B.n831 B.n94 585
R623 B.n830 B.n829 585
R624 B.n828 B.n95 585
R625 B.n827 B.n826 585
R626 B.n825 B.n96 585
R627 B.n824 B.n823 585
R628 B.n822 B.n97 585
R629 B.n821 B.n820 585
R630 B.n819 B.n98 585
R631 B.n818 B.n817 585
R632 B.n816 B.n99 585
R633 B.n815 B.n814 585
R634 B.n813 B.n100 585
R635 B.n812 B.n811 585
R636 B.n810 B.n101 585
R637 B.n809 B.n808 585
R638 B.n807 B.n102 585
R639 B.n806 B.n805 585
R640 B.n981 B.n40 585
R641 B.n983 B.n982 585
R642 B.n984 B.n39 585
R643 B.n986 B.n985 585
R644 B.n987 B.n38 585
R645 B.n989 B.n988 585
R646 B.n990 B.n37 585
R647 B.n992 B.n991 585
R648 B.n993 B.n36 585
R649 B.n995 B.n994 585
R650 B.n996 B.n35 585
R651 B.n998 B.n997 585
R652 B.n999 B.n34 585
R653 B.n1001 B.n1000 585
R654 B.n1002 B.n33 585
R655 B.n1004 B.n1003 585
R656 B.n1005 B.n32 585
R657 B.n1007 B.n1006 585
R658 B.n1008 B.n31 585
R659 B.n1010 B.n1009 585
R660 B.n1011 B.n30 585
R661 B.n1013 B.n1012 585
R662 B.n1014 B.n29 585
R663 B.n1016 B.n1015 585
R664 B.n1017 B.n28 585
R665 B.n1019 B.n1018 585
R666 B.n1020 B.n27 585
R667 B.n1022 B.n1021 585
R668 B.n1023 B.n26 585
R669 B.n1025 B.n1024 585
R670 B.n1026 B.n25 585
R671 B.n1028 B.n1027 585
R672 B.n1029 B.n24 585
R673 B.n1031 B.n1030 585
R674 B.n1032 B.n23 585
R675 B.n1034 B.n1033 585
R676 B.n1035 B.n22 585
R677 B.n1037 B.n1036 585
R678 B.n1038 B.n21 585
R679 B.n1040 B.n1039 585
R680 B.n1041 B.n20 585
R681 B.n1043 B.n1042 585
R682 B.n1044 B.n19 585
R683 B.n1046 B.n1045 585
R684 B.n1047 B.n18 585
R685 B.n1049 B.n1048 585
R686 B.n1050 B.n17 585
R687 B.n1052 B.n1051 585
R688 B.n1053 B.n16 585
R689 B.n1055 B.n1054 585
R690 B.n1056 B.n15 585
R691 B.n1058 B.n1057 585
R692 B.n1059 B.n14 585
R693 B.n1061 B.n1060 585
R694 B.n1062 B.n13 585
R695 B.n1064 B.n1063 585
R696 B.n1065 B.n12 585
R697 B.n1067 B.n1066 585
R698 B.n1068 B.n11 585
R699 B.n1070 B.n1069 585
R700 B.n1071 B.n10 585
R701 B.n1073 B.n1072 585
R702 B.n1074 B.n9 585
R703 B.n1076 B.n1075 585
R704 B.n1077 B.n8 585
R705 B.n1079 B.n1078 585
R706 B.n1080 B.n7 585
R707 B.n1082 B.n1081 585
R708 B.n1083 B.n6 585
R709 B.n1085 B.n1084 585
R710 B.n1086 B.n5 585
R711 B.n1088 B.n1087 585
R712 B.n1089 B.n4 585
R713 B.n1091 B.n1090 585
R714 B.n1092 B.n3 585
R715 B.n1094 B.n1093 585
R716 B.n1095 B.n0 585
R717 B.n2 B.n1 585
R718 B.n280 B.n279 585
R719 B.n281 B.n278 585
R720 B.n283 B.n282 585
R721 B.n284 B.n277 585
R722 B.n286 B.n285 585
R723 B.n287 B.n276 585
R724 B.n289 B.n288 585
R725 B.n290 B.n275 585
R726 B.n292 B.n291 585
R727 B.n293 B.n274 585
R728 B.n295 B.n294 585
R729 B.n296 B.n273 585
R730 B.n298 B.n297 585
R731 B.n299 B.n272 585
R732 B.n301 B.n300 585
R733 B.n302 B.n271 585
R734 B.n304 B.n303 585
R735 B.n305 B.n270 585
R736 B.n307 B.n306 585
R737 B.n308 B.n269 585
R738 B.n310 B.n309 585
R739 B.n311 B.n268 585
R740 B.n313 B.n312 585
R741 B.n314 B.n267 585
R742 B.n316 B.n315 585
R743 B.n317 B.n266 585
R744 B.n319 B.n318 585
R745 B.n320 B.n265 585
R746 B.n322 B.n321 585
R747 B.n323 B.n264 585
R748 B.n325 B.n324 585
R749 B.n326 B.n263 585
R750 B.n328 B.n327 585
R751 B.n329 B.n262 585
R752 B.n331 B.n330 585
R753 B.n332 B.n261 585
R754 B.n334 B.n333 585
R755 B.n335 B.n260 585
R756 B.n337 B.n336 585
R757 B.n338 B.n259 585
R758 B.n340 B.n339 585
R759 B.n341 B.n258 585
R760 B.n343 B.n342 585
R761 B.n344 B.n257 585
R762 B.n346 B.n345 585
R763 B.n347 B.n256 585
R764 B.n349 B.n348 585
R765 B.n350 B.n255 585
R766 B.n352 B.n351 585
R767 B.n353 B.n254 585
R768 B.n355 B.n354 585
R769 B.n356 B.n253 585
R770 B.n358 B.n357 585
R771 B.n359 B.n252 585
R772 B.n361 B.n360 585
R773 B.n362 B.n251 585
R774 B.n364 B.n363 585
R775 B.n365 B.n250 585
R776 B.n367 B.n366 585
R777 B.n368 B.n249 585
R778 B.n370 B.n369 585
R779 B.n371 B.n248 585
R780 B.n373 B.n372 585
R781 B.n374 B.n247 585
R782 B.n376 B.n375 585
R783 B.n377 B.n246 585
R784 B.n379 B.n378 585
R785 B.n380 B.n245 585
R786 B.n382 B.n381 585
R787 B.n383 B.n244 585
R788 B.n385 B.n384 585
R789 B.n386 B.n243 585
R790 B.n388 B.n387 585
R791 B.n389 B.n242 585
R792 B.n391 B.n390 585
R793 B.n392 B.n241 585
R794 B.n394 B.n241 530.939
R795 B.n572 B.n181 530.939
R796 B.n806 B.n103 530.939
R797 B.n981 B.n980 530.939
R798 B.n471 B.t6 315.738
R799 B.n208 B.t9 315.738
R800 B.n74 B.t3 315.738
R801 B.n68 B.t0 315.738
R802 B.n1097 B.n1096 256.663
R803 B.n1096 B.n1095 235.042
R804 B.n1096 B.n2 235.042
R805 B.n208 B.t10 189.049
R806 B.n74 B.t5 189.049
R807 B.n471 B.t7 189.03
R808 B.n68 B.t2 189.03
R809 B.n395 B.n394 163.367
R810 B.n396 B.n395 163.367
R811 B.n396 B.n239 163.367
R812 B.n400 B.n239 163.367
R813 B.n401 B.n400 163.367
R814 B.n402 B.n401 163.367
R815 B.n402 B.n237 163.367
R816 B.n406 B.n237 163.367
R817 B.n407 B.n406 163.367
R818 B.n408 B.n407 163.367
R819 B.n408 B.n235 163.367
R820 B.n412 B.n235 163.367
R821 B.n413 B.n412 163.367
R822 B.n414 B.n413 163.367
R823 B.n414 B.n233 163.367
R824 B.n418 B.n233 163.367
R825 B.n419 B.n418 163.367
R826 B.n420 B.n419 163.367
R827 B.n420 B.n231 163.367
R828 B.n424 B.n231 163.367
R829 B.n425 B.n424 163.367
R830 B.n426 B.n425 163.367
R831 B.n426 B.n229 163.367
R832 B.n430 B.n229 163.367
R833 B.n431 B.n430 163.367
R834 B.n432 B.n431 163.367
R835 B.n432 B.n227 163.367
R836 B.n436 B.n227 163.367
R837 B.n437 B.n436 163.367
R838 B.n438 B.n437 163.367
R839 B.n438 B.n225 163.367
R840 B.n442 B.n225 163.367
R841 B.n443 B.n442 163.367
R842 B.n444 B.n443 163.367
R843 B.n444 B.n223 163.367
R844 B.n448 B.n223 163.367
R845 B.n449 B.n448 163.367
R846 B.n450 B.n449 163.367
R847 B.n450 B.n221 163.367
R848 B.n454 B.n221 163.367
R849 B.n455 B.n454 163.367
R850 B.n456 B.n455 163.367
R851 B.n456 B.n219 163.367
R852 B.n460 B.n219 163.367
R853 B.n461 B.n460 163.367
R854 B.n462 B.n461 163.367
R855 B.n462 B.n217 163.367
R856 B.n466 B.n217 163.367
R857 B.n467 B.n466 163.367
R858 B.n468 B.n467 163.367
R859 B.n468 B.n215 163.367
R860 B.n475 B.n215 163.367
R861 B.n476 B.n475 163.367
R862 B.n477 B.n476 163.367
R863 B.n477 B.n213 163.367
R864 B.n481 B.n213 163.367
R865 B.n482 B.n481 163.367
R866 B.n483 B.n482 163.367
R867 B.n483 B.n211 163.367
R868 B.n487 B.n211 163.367
R869 B.n488 B.n487 163.367
R870 B.n489 B.n488 163.367
R871 B.n489 B.n207 163.367
R872 B.n494 B.n207 163.367
R873 B.n495 B.n494 163.367
R874 B.n496 B.n495 163.367
R875 B.n496 B.n205 163.367
R876 B.n500 B.n205 163.367
R877 B.n501 B.n500 163.367
R878 B.n502 B.n501 163.367
R879 B.n502 B.n203 163.367
R880 B.n506 B.n203 163.367
R881 B.n507 B.n506 163.367
R882 B.n508 B.n507 163.367
R883 B.n508 B.n201 163.367
R884 B.n512 B.n201 163.367
R885 B.n513 B.n512 163.367
R886 B.n514 B.n513 163.367
R887 B.n514 B.n199 163.367
R888 B.n518 B.n199 163.367
R889 B.n519 B.n518 163.367
R890 B.n520 B.n519 163.367
R891 B.n520 B.n197 163.367
R892 B.n524 B.n197 163.367
R893 B.n525 B.n524 163.367
R894 B.n526 B.n525 163.367
R895 B.n526 B.n195 163.367
R896 B.n530 B.n195 163.367
R897 B.n531 B.n530 163.367
R898 B.n532 B.n531 163.367
R899 B.n532 B.n193 163.367
R900 B.n536 B.n193 163.367
R901 B.n537 B.n536 163.367
R902 B.n538 B.n537 163.367
R903 B.n538 B.n191 163.367
R904 B.n542 B.n191 163.367
R905 B.n543 B.n542 163.367
R906 B.n544 B.n543 163.367
R907 B.n544 B.n189 163.367
R908 B.n548 B.n189 163.367
R909 B.n549 B.n548 163.367
R910 B.n550 B.n549 163.367
R911 B.n550 B.n187 163.367
R912 B.n554 B.n187 163.367
R913 B.n555 B.n554 163.367
R914 B.n556 B.n555 163.367
R915 B.n556 B.n185 163.367
R916 B.n560 B.n185 163.367
R917 B.n561 B.n560 163.367
R918 B.n562 B.n561 163.367
R919 B.n562 B.n183 163.367
R920 B.n566 B.n183 163.367
R921 B.n567 B.n566 163.367
R922 B.n568 B.n567 163.367
R923 B.n568 B.n181 163.367
R924 B.n802 B.n103 163.367
R925 B.n802 B.n801 163.367
R926 B.n801 B.n800 163.367
R927 B.n800 B.n105 163.367
R928 B.n796 B.n105 163.367
R929 B.n796 B.n795 163.367
R930 B.n795 B.n794 163.367
R931 B.n794 B.n107 163.367
R932 B.n790 B.n107 163.367
R933 B.n790 B.n789 163.367
R934 B.n789 B.n788 163.367
R935 B.n788 B.n109 163.367
R936 B.n784 B.n109 163.367
R937 B.n784 B.n783 163.367
R938 B.n783 B.n782 163.367
R939 B.n782 B.n111 163.367
R940 B.n778 B.n111 163.367
R941 B.n778 B.n777 163.367
R942 B.n777 B.n776 163.367
R943 B.n776 B.n113 163.367
R944 B.n772 B.n113 163.367
R945 B.n772 B.n771 163.367
R946 B.n771 B.n770 163.367
R947 B.n770 B.n115 163.367
R948 B.n766 B.n115 163.367
R949 B.n766 B.n765 163.367
R950 B.n765 B.n764 163.367
R951 B.n764 B.n117 163.367
R952 B.n760 B.n117 163.367
R953 B.n760 B.n759 163.367
R954 B.n759 B.n758 163.367
R955 B.n758 B.n119 163.367
R956 B.n754 B.n119 163.367
R957 B.n754 B.n753 163.367
R958 B.n753 B.n752 163.367
R959 B.n752 B.n121 163.367
R960 B.n748 B.n121 163.367
R961 B.n748 B.n747 163.367
R962 B.n747 B.n746 163.367
R963 B.n746 B.n123 163.367
R964 B.n742 B.n123 163.367
R965 B.n742 B.n741 163.367
R966 B.n741 B.n740 163.367
R967 B.n740 B.n125 163.367
R968 B.n736 B.n125 163.367
R969 B.n736 B.n735 163.367
R970 B.n735 B.n734 163.367
R971 B.n734 B.n127 163.367
R972 B.n730 B.n127 163.367
R973 B.n730 B.n729 163.367
R974 B.n729 B.n728 163.367
R975 B.n728 B.n129 163.367
R976 B.n724 B.n129 163.367
R977 B.n724 B.n723 163.367
R978 B.n723 B.n722 163.367
R979 B.n722 B.n131 163.367
R980 B.n718 B.n131 163.367
R981 B.n718 B.n717 163.367
R982 B.n717 B.n716 163.367
R983 B.n716 B.n133 163.367
R984 B.n712 B.n133 163.367
R985 B.n712 B.n711 163.367
R986 B.n711 B.n710 163.367
R987 B.n710 B.n135 163.367
R988 B.n706 B.n135 163.367
R989 B.n706 B.n705 163.367
R990 B.n705 B.n704 163.367
R991 B.n704 B.n137 163.367
R992 B.n700 B.n137 163.367
R993 B.n700 B.n699 163.367
R994 B.n699 B.n698 163.367
R995 B.n698 B.n139 163.367
R996 B.n694 B.n139 163.367
R997 B.n694 B.n693 163.367
R998 B.n693 B.n692 163.367
R999 B.n692 B.n141 163.367
R1000 B.n688 B.n141 163.367
R1001 B.n688 B.n687 163.367
R1002 B.n687 B.n686 163.367
R1003 B.n686 B.n143 163.367
R1004 B.n682 B.n143 163.367
R1005 B.n682 B.n681 163.367
R1006 B.n681 B.n680 163.367
R1007 B.n680 B.n145 163.367
R1008 B.n676 B.n145 163.367
R1009 B.n676 B.n675 163.367
R1010 B.n675 B.n674 163.367
R1011 B.n674 B.n147 163.367
R1012 B.n670 B.n147 163.367
R1013 B.n670 B.n669 163.367
R1014 B.n669 B.n668 163.367
R1015 B.n668 B.n149 163.367
R1016 B.n664 B.n149 163.367
R1017 B.n664 B.n663 163.367
R1018 B.n663 B.n662 163.367
R1019 B.n662 B.n151 163.367
R1020 B.n658 B.n151 163.367
R1021 B.n658 B.n657 163.367
R1022 B.n657 B.n656 163.367
R1023 B.n656 B.n153 163.367
R1024 B.n652 B.n153 163.367
R1025 B.n652 B.n651 163.367
R1026 B.n651 B.n650 163.367
R1027 B.n650 B.n155 163.367
R1028 B.n646 B.n155 163.367
R1029 B.n646 B.n645 163.367
R1030 B.n645 B.n644 163.367
R1031 B.n644 B.n157 163.367
R1032 B.n640 B.n157 163.367
R1033 B.n640 B.n639 163.367
R1034 B.n639 B.n638 163.367
R1035 B.n638 B.n159 163.367
R1036 B.n634 B.n159 163.367
R1037 B.n634 B.n633 163.367
R1038 B.n633 B.n632 163.367
R1039 B.n632 B.n161 163.367
R1040 B.n628 B.n161 163.367
R1041 B.n628 B.n627 163.367
R1042 B.n627 B.n626 163.367
R1043 B.n626 B.n163 163.367
R1044 B.n622 B.n163 163.367
R1045 B.n622 B.n621 163.367
R1046 B.n621 B.n620 163.367
R1047 B.n620 B.n165 163.367
R1048 B.n616 B.n165 163.367
R1049 B.n616 B.n615 163.367
R1050 B.n615 B.n614 163.367
R1051 B.n614 B.n167 163.367
R1052 B.n610 B.n167 163.367
R1053 B.n610 B.n609 163.367
R1054 B.n609 B.n608 163.367
R1055 B.n608 B.n169 163.367
R1056 B.n604 B.n169 163.367
R1057 B.n604 B.n603 163.367
R1058 B.n603 B.n602 163.367
R1059 B.n602 B.n171 163.367
R1060 B.n598 B.n171 163.367
R1061 B.n598 B.n597 163.367
R1062 B.n597 B.n596 163.367
R1063 B.n596 B.n173 163.367
R1064 B.n592 B.n173 163.367
R1065 B.n592 B.n591 163.367
R1066 B.n591 B.n590 163.367
R1067 B.n590 B.n175 163.367
R1068 B.n586 B.n175 163.367
R1069 B.n586 B.n585 163.367
R1070 B.n585 B.n584 163.367
R1071 B.n584 B.n177 163.367
R1072 B.n580 B.n177 163.367
R1073 B.n580 B.n579 163.367
R1074 B.n579 B.n578 163.367
R1075 B.n578 B.n179 163.367
R1076 B.n574 B.n179 163.367
R1077 B.n574 B.n573 163.367
R1078 B.n573 B.n572 163.367
R1079 B.n980 B.n41 163.367
R1080 B.n976 B.n41 163.367
R1081 B.n976 B.n975 163.367
R1082 B.n975 B.n974 163.367
R1083 B.n974 B.n43 163.367
R1084 B.n970 B.n43 163.367
R1085 B.n970 B.n969 163.367
R1086 B.n969 B.n968 163.367
R1087 B.n968 B.n45 163.367
R1088 B.n964 B.n45 163.367
R1089 B.n964 B.n963 163.367
R1090 B.n963 B.n962 163.367
R1091 B.n962 B.n47 163.367
R1092 B.n958 B.n47 163.367
R1093 B.n958 B.n957 163.367
R1094 B.n957 B.n956 163.367
R1095 B.n956 B.n49 163.367
R1096 B.n952 B.n49 163.367
R1097 B.n952 B.n951 163.367
R1098 B.n951 B.n950 163.367
R1099 B.n950 B.n51 163.367
R1100 B.n946 B.n51 163.367
R1101 B.n946 B.n945 163.367
R1102 B.n945 B.n944 163.367
R1103 B.n944 B.n53 163.367
R1104 B.n940 B.n53 163.367
R1105 B.n940 B.n939 163.367
R1106 B.n939 B.n938 163.367
R1107 B.n938 B.n55 163.367
R1108 B.n934 B.n55 163.367
R1109 B.n934 B.n933 163.367
R1110 B.n933 B.n932 163.367
R1111 B.n932 B.n57 163.367
R1112 B.n928 B.n57 163.367
R1113 B.n928 B.n927 163.367
R1114 B.n927 B.n926 163.367
R1115 B.n926 B.n59 163.367
R1116 B.n922 B.n59 163.367
R1117 B.n922 B.n921 163.367
R1118 B.n921 B.n920 163.367
R1119 B.n920 B.n61 163.367
R1120 B.n916 B.n61 163.367
R1121 B.n916 B.n915 163.367
R1122 B.n915 B.n914 163.367
R1123 B.n914 B.n63 163.367
R1124 B.n910 B.n63 163.367
R1125 B.n910 B.n909 163.367
R1126 B.n909 B.n908 163.367
R1127 B.n908 B.n65 163.367
R1128 B.n904 B.n65 163.367
R1129 B.n904 B.n903 163.367
R1130 B.n903 B.n902 163.367
R1131 B.n902 B.n67 163.367
R1132 B.n897 B.n67 163.367
R1133 B.n897 B.n896 163.367
R1134 B.n896 B.n895 163.367
R1135 B.n895 B.n71 163.367
R1136 B.n891 B.n71 163.367
R1137 B.n891 B.n890 163.367
R1138 B.n890 B.n889 163.367
R1139 B.n889 B.n73 163.367
R1140 B.n885 B.n73 163.367
R1141 B.n885 B.n884 163.367
R1142 B.n884 B.n77 163.367
R1143 B.n880 B.n77 163.367
R1144 B.n880 B.n879 163.367
R1145 B.n879 B.n878 163.367
R1146 B.n878 B.n79 163.367
R1147 B.n874 B.n79 163.367
R1148 B.n874 B.n873 163.367
R1149 B.n873 B.n872 163.367
R1150 B.n872 B.n81 163.367
R1151 B.n868 B.n81 163.367
R1152 B.n868 B.n867 163.367
R1153 B.n867 B.n866 163.367
R1154 B.n866 B.n83 163.367
R1155 B.n862 B.n83 163.367
R1156 B.n862 B.n861 163.367
R1157 B.n861 B.n860 163.367
R1158 B.n860 B.n85 163.367
R1159 B.n856 B.n85 163.367
R1160 B.n856 B.n855 163.367
R1161 B.n855 B.n854 163.367
R1162 B.n854 B.n87 163.367
R1163 B.n850 B.n87 163.367
R1164 B.n850 B.n849 163.367
R1165 B.n849 B.n848 163.367
R1166 B.n848 B.n89 163.367
R1167 B.n844 B.n89 163.367
R1168 B.n844 B.n843 163.367
R1169 B.n843 B.n842 163.367
R1170 B.n842 B.n91 163.367
R1171 B.n838 B.n91 163.367
R1172 B.n838 B.n837 163.367
R1173 B.n837 B.n836 163.367
R1174 B.n836 B.n93 163.367
R1175 B.n832 B.n93 163.367
R1176 B.n832 B.n831 163.367
R1177 B.n831 B.n830 163.367
R1178 B.n830 B.n95 163.367
R1179 B.n826 B.n95 163.367
R1180 B.n826 B.n825 163.367
R1181 B.n825 B.n824 163.367
R1182 B.n824 B.n97 163.367
R1183 B.n820 B.n97 163.367
R1184 B.n820 B.n819 163.367
R1185 B.n819 B.n818 163.367
R1186 B.n818 B.n99 163.367
R1187 B.n814 B.n99 163.367
R1188 B.n814 B.n813 163.367
R1189 B.n813 B.n812 163.367
R1190 B.n812 B.n101 163.367
R1191 B.n808 B.n101 163.367
R1192 B.n808 B.n807 163.367
R1193 B.n807 B.n806 163.367
R1194 B.n982 B.n981 163.367
R1195 B.n982 B.n39 163.367
R1196 B.n986 B.n39 163.367
R1197 B.n987 B.n986 163.367
R1198 B.n988 B.n987 163.367
R1199 B.n988 B.n37 163.367
R1200 B.n992 B.n37 163.367
R1201 B.n993 B.n992 163.367
R1202 B.n994 B.n993 163.367
R1203 B.n994 B.n35 163.367
R1204 B.n998 B.n35 163.367
R1205 B.n999 B.n998 163.367
R1206 B.n1000 B.n999 163.367
R1207 B.n1000 B.n33 163.367
R1208 B.n1004 B.n33 163.367
R1209 B.n1005 B.n1004 163.367
R1210 B.n1006 B.n1005 163.367
R1211 B.n1006 B.n31 163.367
R1212 B.n1010 B.n31 163.367
R1213 B.n1011 B.n1010 163.367
R1214 B.n1012 B.n1011 163.367
R1215 B.n1012 B.n29 163.367
R1216 B.n1016 B.n29 163.367
R1217 B.n1017 B.n1016 163.367
R1218 B.n1018 B.n1017 163.367
R1219 B.n1018 B.n27 163.367
R1220 B.n1022 B.n27 163.367
R1221 B.n1023 B.n1022 163.367
R1222 B.n1024 B.n1023 163.367
R1223 B.n1024 B.n25 163.367
R1224 B.n1028 B.n25 163.367
R1225 B.n1029 B.n1028 163.367
R1226 B.n1030 B.n1029 163.367
R1227 B.n1030 B.n23 163.367
R1228 B.n1034 B.n23 163.367
R1229 B.n1035 B.n1034 163.367
R1230 B.n1036 B.n1035 163.367
R1231 B.n1036 B.n21 163.367
R1232 B.n1040 B.n21 163.367
R1233 B.n1041 B.n1040 163.367
R1234 B.n1042 B.n1041 163.367
R1235 B.n1042 B.n19 163.367
R1236 B.n1046 B.n19 163.367
R1237 B.n1047 B.n1046 163.367
R1238 B.n1048 B.n1047 163.367
R1239 B.n1048 B.n17 163.367
R1240 B.n1052 B.n17 163.367
R1241 B.n1053 B.n1052 163.367
R1242 B.n1054 B.n1053 163.367
R1243 B.n1054 B.n15 163.367
R1244 B.n1058 B.n15 163.367
R1245 B.n1059 B.n1058 163.367
R1246 B.n1060 B.n1059 163.367
R1247 B.n1060 B.n13 163.367
R1248 B.n1064 B.n13 163.367
R1249 B.n1065 B.n1064 163.367
R1250 B.n1066 B.n1065 163.367
R1251 B.n1066 B.n11 163.367
R1252 B.n1070 B.n11 163.367
R1253 B.n1071 B.n1070 163.367
R1254 B.n1072 B.n1071 163.367
R1255 B.n1072 B.n9 163.367
R1256 B.n1076 B.n9 163.367
R1257 B.n1077 B.n1076 163.367
R1258 B.n1078 B.n1077 163.367
R1259 B.n1078 B.n7 163.367
R1260 B.n1082 B.n7 163.367
R1261 B.n1083 B.n1082 163.367
R1262 B.n1084 B.n1083 163.367
R1263 B.n1084 B.n5 163.367
R1264 B.n1088 B.n5 163.367
R1265 B.n1089 B.n1088 163.367
R1266 B.n1090 B.n1089 163.367
R1267 B.n1090 B.n3 163.367
R1268 B.n1094 B.n3 163.367
R1269 B.n1095 B.n1094 163.367
R1270 B.n280 B.n2 163.367
R1271 B.n281 B.n280 163.367
R1272 B.n282 B.n281 163.367
R1273 B.n282 B.n277 163.367
R1274 B.n286 B.n277 163.367
R1275 B.n287 B.n286 163.367
R1276 B.n288 B.n287 163.367
R1277 B.n288 B.n275 163.367
R1278 B.n292 B.n275 163.367
R1279 B.n293 B.n292 163.367
R1280 B.n294 B.n293 163.367
R1281 B.n294 B.n273 163.367
R1282 B.n298 B.n273 163.367
R1283 B.n299 B.n298 163.367
R1284 B.n300 B.n299 163.367
R1285 B.n300 B.n271 163.367
R1286 B.n304 B.n271 163.367
R1287 B.n305 B.n304 163.367
R1288 B.n306 B.n305 163.367
R1289 B.n306 B.n269 163.367
R1290 B.n310 B.n269 163.367
R1291 B.n311 B.n310 163.367
R1292 B.n312 B.n311 163.367
R1293 B.n312 B.n267 163.367
R1294 B.n316 B.n267 163.367
R1295 B.n317 B.n316 163.367
R1296 B.n318 B.n317 163.367
R1297 B.n318 B.n265 163.367
R1298 B.n322 B.n265 163.367
R1299 B.n323 B.n322 163.367
R1300 B.n324 B.n323 163.367
R1301 B.n324 B.n263 163.367
R1302 B.n328 B.n263 163.367
R1303 B.n329 B.n328 163.367
R1304 B.n330 B.n329 163.367
R1305 B.n330 B.n261 163.367
R1306 B.n334 B.n261 163.367
R1307 B.n335 B.n334 163.367
R1308 B.n336 B.n335 163.367
R1309 B.n336 B.n259 163.367
R1310 B.n340 B.n259 163.367
R1311 B.n341 B.n340 163.367
R1312 B.n342 B.n341 163.367
R1313 B.n342 B.n257 163.367
R1314 B.n346 B.n257 163.367
R1315 B.n347 B.n346 163.367
R1316 B.n348 B.n347 163.367
R1317 B.n348 B.n255 163.367
R1318 B.n352 B.n255 163.367
R1319 B.n353 B.n352 163.367
R1320 B.n354 B.n353 163.367
R1321 B.n354 B.n253 163.367
R1322 B.n358 B.n253 163.367
R1323 B.n359 B.n358 163.367
R1324 B.n360 B.n359 163.367
R1325 B.n360 B.n251 163.367
R1326 B.n364 B.n251 163.367
R1327 B.n365 B.n364 163.367
R1328 B.n366 B.n365 163.367
R1329 B.n366 B.n249 163.367
R1330 B.n370 B.n249 163.367
R1331 B.n371 B.n370 163.367
R1332 B.n372 B.n371 163.367
R1333 B.n372 B.n247 163.367
R1334 B.n376 B.n247 163.367
R1335 B.n377 B.n376 163.367
R1336 B.n378 B.n377 163.367
R1337 B.n378 B.n245 163.367
R1338 B.n382 B.n245 163.367
R1339 B.n383 B.n382 163.367
R1340 B.n384 B.n383 163.367
R1341 B.n384 B.n243 163.367
R1342 B.n388 B.n243 163.367
R1343 B.n389 B.n388 163.367
R1344 B.n390 B.n389 163.367
R1345 B.n390 B.n241 163.367
R1346 B.n209 B.t11 112.638
R1347 B.n75 B.t4 112.638
R1348 B.n472 B.t8 112.618
R1349 B.n69 B.t1 112.618
R1350 B.n472 B.n471 76.4126
R1351 B.n209 B.n208 76.4126
R1352 B.n75 B.n74 76.4126
R1353 B.n69 B.n68 76.4126
R1354 B.n473 B.n472 59.5399
R1355 B.n491 B.n209 59.5399
R1356 B.n76 B.n75 59.5399
R1357 B.n900 B.n69 59.5399
R1358 B.n979 B.n40 34.4981
R1359 B.n805 B.n804 34.4981
R1360 B.n571 B.n570 34.4981
R1361 B.n393 B.n392 34.4981
R1362 B B.n1097 18.0485
R1363 B.n983 B.n40 10.6151
R1364 B.n984 B.n983 10.6151
R1365 B.n985 B.n984 10.6151
R1366 B.n985 B.n38 10.6151
R1367 B.n989 B.n38 10.6151
R1368 B.n990 B.n989 10.6151
R1369 B.n991 B.n990 10.6151
R1370 B.n991 B.n36 10.6151
R1371 B.n995 B.n36 10.6151
R1372 B.n996 B.n995 10.6151
R1373 B.n997 B.n996 10.6151
R1374 B.n997 B.n34 10.6151
R1375 B.n1001 B.n34 10.6151
R1376 B.n1002 B.n1001 10.6151
R1377 B.n1003 B.n1002 10.6151
R1378 B.n1003 B.n32 10.6151
R1379 B.n1007 B.n32 10.6151
R1380 B.n1008 B.n1007 10.6151
R1381 B.n1009 B.n1008 10.6151
R1382 B.n1009 B.n30 10.6151
R1383 B.n1013 B.n30 10.6151
R1384 B.n1014 B.n1013 10.6151
R1385 B.n1015 B.n1014 10.6151
R1386 B.n1015 B.n28 10.6151
R1387 B.n1019 B.n28 10.6151
R1388 B.n1020 B.n1019 10.6151
R1389 B.n1021 B.n1020 10.6151
R1390 B.n1021 B.n26 10.6151
R1391 B.n1025 B.n26 10.6151
R1392 B.n1026 B.n1025 10.6151
R1393 B.n1027 B.n1026 10.6151
R1394 B.n1027 B.n24 10.6151
R1395 B.n1031 B.n24 10.6151
R1396 B.n1032 B.n1031 10.6151
R1397 B.n1033 B.n1032 10.6151
R1398 B.n1033 B.n22 10.6151
R1399 B.n1037 B.n22 10.6151
R1400 B.n1038 B.n1037 10.6151
R1401 B.n1039 B.n1038 10.6151
R1402 B.n1039 B.n20 10.6151
R1403 B.n1043 B.n20 10.6151
R1404 B.n1044 B.n1043 10.6151
R1405 B.n1045 B.n1044 10.6151
R1406 B.n1045 B.n18 10.6151
R1407 B.n1049 B.n18 10.6151
R1408 B.n1050 B.n1049 10.6151
R1409 B.n1051 B.n1050 10.6151
R1410 B.n1051 B.n16 10.6151
R1411 B.n1055 B.n16 10.6151
R1412 B.n1056 B.n1055 10.6151
R1413 B.n1057 B.n1056 10.6151
R1414 B.n1057 B.n14 10.6151
R1415 B.n1061 B.n14 10.6151
R1416 B.n1062 B.n1061 10.6151
R1417 B.n1063 B.n1062 10.6151
R1418 B.n1063 B.n12 10.6151
R1419 B.n1067 B.n12 10.6151
R1420 B.n1068 B.n1067 10.6151
R1421 B.n1069 B.n1068 10.6151
R1422 B.n1069 B.n10 10.6151
R1423 B.n1073 B.n10 10.6151
R1424 B.n1074 B.n1073 10.6151
R1425 B.n1075 B.n1074 10.6151
R1426 B.n1075 B.n8 10.6151
R1427 B.n1079 B.n8 10.6151
R1428 B.n1080 B.n1079 10.6151
R1429 B.n1081 B.n1080 10.6151
R1430 B.n1081 B.n6 10.6151
R1431 B.n1085 B.n6 10.6151
R1432 B.n1086 B.n1085 10.6151
R1433 B.n1087 B.n1086 10.6151
R1434 B.n1087 B.n4 10.6151
R1435 B.n1091 B.n4 10.6151
R1436 B.n1092 B.n1091 10.6151
R1437 B.n1093 B.n1092 10.6151
R1438 B.n1093 B.n0 10.6151
R1439 B.n979 B.n978 10.6151
R1440 B.n978 B.n977 10.6151
R1441 B.n977 B.n42 10.6151
R1442 B.n973 B.n42 10.6151
R1443 B.n973 B.n972 10.6151
R1444 B.n972 B.n971 10.6151
R1445 B.n971 B.n44 10.6151
R1446 B.n967 B.n44 10.6151
R1447 B.n967 B.n966 10.6151
R1448 B.n966 B.n965 10.6151
R1449 B.n965 B.n46 10.6151
R1450 B.n961 B.n46 10.6151
R1451 B.n961 B.n960 10.6151
R1452 B.n960 B.n959 10.6151
R1453 B.n959 B.n48 10.6151
R1454 B.n955 B.n48 10.6151
R1455 B.n955 B.n954 10.6151
R1456 B.n954 B.n953 10.6151
R1457 B.n953 B.n50 10.6151
R1458 B.n949 B.n50 10.6151
R1459 B.n949 B.n948 10.6151
R1460 B.n948 B.n947 10.6151
R1461 B.n947 B.n52 10.6151
R1462 B.n943 B.n52 10.6151
R1463 B.n943 B.n942 10.6151
R1464 B.n942 B.n941 10.6151
R1465 B.n941 B.n54 10.6151
R1466 B.n937 B.n54 10.6151
R1467 B.n937 B.n936 10.6151
R1468 B.n936 B.n935 10.6151
R1469 B.n935 B.n56 10.6151
R1470 B.n931 B.n56 10.6151
R1471 B.n931 B.n930 10.6151
R1472 B.n930 B.n929 10.6151
R1473 B.n929 B.n58 10.6151
R1474 B.n925 B.n58 10.6151
R1475 B.n925 B.n924 10.6151
R1476 B.n924 B.n923 10.6151
R1477 B.n923 B.n60 10.6151
R1478 B.n919 B.n60 10.6151
R1479 B.n919 B.n918 10.6151
R1480 B.n918 B.n917 10.6151
R1481 B.n917 B.n62 10.6151
R1482 B.n913 B.n62 10.6151
R1483 B.n913 B.n912 10.6151
R1484 B.n912 B.n911 10.6151
R1485 B.n911 B.n64 10.6151
R1486 B.n907 B.n64 10.6151
R1487 B.n907 B.n906 10.6151
R1488 B.n906 B.n905 10.6151
R1489 B.n905 B.n66 10.6151
R1490 B.n901 B.n66 10.6151
R1491 B.n899 B.n898 10.6151
R1492 B.n898 B.n70 10.6151
R1493 B.n894 B.n70 10.6151
R1494 B.n894 B.n893 10.6151
R1495 B.n893 B.n892 10.6151
R1496 B.n892 B.n72 10.6151
R1497 B.n888 B.n72 10.6151
R1498 B.n888 B.n887 10.6151
R1499 B.n887 B.n886 10.6151
R1500 B.n883 B.n882 10.6151
R1501 B.n882 B.n881 10.6151
R1502 B.n881 B.n78 10.6151
R1503 B.n877 B.n78 10.6151
R1504 B.n877 B.n876 10.6151
R1505 B.n876 B.n875 10.6151
R1506 B.n875 B.n80 10.6151
R1507 B.n871 B.n80 10.6151
R1508 B.n871 B.n870 10.6151
R1509 B.n870 B.n869 10.6151
R1510 B.n869 B.n82 10.6151
R1511 B.n865 B.n82 10.6151
R1512 B.n865 B.n864 10.6151
R1513 B.n864 B.n863 10.6151
R1514 B.n863 B.n84 10.6151
R1515 B.n859 B.n84 10.6151
R1516 B.n859 B.n858 10.6151
R1517 B.n858 B.n857 10.6151
R1518 B.n857 B.n86 10.6151
R1519 B.n853 B.n86 10.6151
R1520 B.n853 B.n852 10.6151
R1521 B.n852 B.n851 10.6151
R1522 B.n851 B.n88 10.6151
R1523 B.n847 B.n88 10.6151
R1524 B.n847 B.n846 10.6151
R1525 B.n846 B.n845 10.6151
R1526 B.n845 B.n90 10.6151
R1527 B.n841 B.n90 10.6151
R1528 B.n841 B.n840 10.6151
R1529 B.n840 B.n839 10.6151
R1530 B.n839 B.n92 10.6151
R1531 B.n835 B.n92 10.6151
R1532 B.n835 B.n834 10.6151
R1533 B.n834 B.n833 10.6151
R1534 B.n833 B.n94 10.6151
R1535 B.n829 B.n94 10.6151
R1536 B.n829 B.n828 10.6151
R1537 B.n828 B.n827 10.6151
R1538 B.n827 B.n96 10.6151
R1539 B.n823 B.n96 10.6151
R1540 B.n823 B.n822 10.6151
R1541 B.n822 B.n821 10.6151
R1542 B.n821 B.n98 10.6151
R1543 B.n817 B.n98 10.6151
R1544 B.n817 B.n816 10.6151
R1545 B.n816 B.n815 10.6151
R1546 B.n815 B.n100 10.6151
R1547 B.n811 B.n100 10.6151
R1548 B.n811 B.n810 10.6151
R1549 B.n810 B.n809 10.6151
R1550 B.n809 B.n102 10.6151
R1551 B.n805 B.n102 10.6151
R1552 B.n804 B.n803 10.6151
R1553 B.n803 B.n104 10.6151
R1554 B.n799 B.n104 10.6151
R1555 B.n799 B.n798 10.6151
R1556 B.n798 B.n797 10.6151
R1557 B.n797 B.n106 10.6151
R1558 B.n793 B.n106 10.6151
R1559 B.n793 B.n792 10.6151
R1560 B.n792 B.n791 10.6151
R1561 B.n791 B.n108 10.6151
R1562 B.n787 B.n108 10.6151
R1563 B.n787 B.n786 10.6151
R1564 B.n786 B.n785 10.6151
R1565 B.n785 B.n110 10.6151
R1566 B.n781 B.n110 10.6151
R1567 B.n781 B.n780 10.6151
R1568 B.n780 B.n779 10.6151
R1569 B.n779 B.n112 10.6151
R1570 B.n775 B.n112 10.6151
R1571 B.n775 B.n774 10.6151
R1572 B.n774 B.n773 10.6151
R1573 B.n773 B.n114 10.6151
R1574 B.n769 B.n114 10.6151
R1575 B.n769 B.n768 10.6151
R1576 B.n768 B.n767 10.6151
R1577 B.n767 B.n116 10.6151
R1578 B.n763 B.n116 10.6151
R1579 B.n763 B.n762 10.6151
R1580 B.n762 B.n761 10.6151
R1581 B.n761 B.n118 10.6151
R1582 B.n757 B.n118 10.6151
R1583 B.n757 B.n756 10.6151
R1584 B.n756 B.n755 10.6151
R1585 B.n755 B.n120 10.6151
R1586 B.n751 B.n120 10.6151
R1587 B.n751 B.n750 10.6151
R1588 B.n750 B.n749 10.6151
R1589 B.n749 B.n122 10.6151
R1590 B.n745 B.n122 10.6151
R1591 B.n745 B.n744 10.6151
R1592 B.n744 B.n743 10.6151
R1593 B.n743 B.n124 10.6151
R1594 B.n739 B.n124 10.6151
R1595 B.n739 B.n738 10.6151
R1596 B.n738 B.n737 10.6151
R1597 B.n737 B.n126 10.6151
R1598 B.n733 B.n126 10.6151
R1599 B.n733 B.n732 10.6151
R1600 B.n732 B.n731 10.6151
R1601 B.n731 B.n128 10.6151
R1602 B.n727 B.n128 10.6151
R1603 B.n727 B.n726 10.6151
R1604 B.n726 B.n725 10.6151
R1605 B.n725 B.n130 10.6151
R1606 B.n721 B.n130 10.6151
R1607 B.n721 B.n720 10.6151
R1608 B.n720 B.n719 10.6151
R1609 B.n719 B.n132 10.6151
R1610 B.n715 B.n132 10.6151
R1611 B.n715 B.n714 10.6151
R1612 B.n714 B.n713 10.6151
R1613 B.n713 B.n134 10.6151
R1614 B.n709 B.n134 10.6151
R1615 B.n709 B.n708 10.6151
R1616 B.n708 B.n707 10.6151
R1617 B.n707 B.n136 10.6151
R1618 B.n703 B.n136 10.6151
R1619 B.n703 B.n702 10.6151
R1620 B.n702 B.n701 10.6151
R1621 B.n701 B.n138 10.6151
R1622 B.n697 B.n138 10.6151
R1623 B.n697 B.n696 10.6151
R1624 B.n696 B.n695 10.6151
R1625 B.n695 B.n140 10.6151
R1626 B.n691 B.n140 10.6151
R1627 B.n691 B.n690 10.6151
R1628 B.n690 B.n689 10.6151
R1629 B.n689 B.n142 10.6151
R1630 B.n685 B.n142 10.6151
R1631 B.n685 B.n684 10.6151
R1632 B.n684 B.n683 10.6151
R1633 B.n683 B.n144 10.6151
R1634 B.n679 B.n144 10.6151
R1635 B.n679 B.n678 10.6151
R1636 B.n678 B.n677 10.6151
R1637 B.n677 B.n146 10.6151
R1638 B.n673 B.n146 10.6151
R1639 B.n673 B.n672 10.6151
R1640 B.n672 B.n671 10.6151
R1641 B.n671 B.n148 10.6151
R1642 B.n667 B.n148 10.6151
R1643 B.n667 B.n666 10.6151
R1644 B.n666 B.n665 10.6151
R1645 B.n665 B.n150 10.6151
R1646 B.n661 B.n150 10.6151
R1647 B.n661 B.n660 10.6151
R1648 B.n660 B.n659 10.6151
R1649 B.n659 B.n152 10.6151
R1650 B.n655 B.n152 10.6151
R1651 B.n655 B.n654 10.6151
R1652 B.n654 B.n653 10.6151
R1653 B.n653 B.n154 10.6151
R1654 B.n649 B.n154 10.6151
R1655 B.n649 B.n648 10.6151
R1656 B.n648 B.n647 10.6151
R1657 B.n647 B.n156 10.6151
R1658 B.n643 B.n156 10.6151
R1659 B.n643 B.n642 10.6151
R1660 B.n642 B.n641 10.6151
R1661 B.n641 B.n158 10.6151
R1662 B.n637 B.n158 10.6151
R1663 B.n637 B.n636 10.6151
R1664 B.n636 B.n635 10.6151
R1665 B.n635 B.n160 10.6151
R1666 B.n631 B.n160 10.6151
R1667 B.n631 B.n630 10.6151
R1668 B.n630 B.n629 10.6151
R1669 B.n629 B.n162 10.6151
R1670 B.n625 B.n162 10.6151
R1671 B.n625 B.n624 10.6151
R1672 B.n624 B.n623 10.6151
R1673 B.n623 B.n164 10.6151
R1674 B.n619 B.n164 10.6151
R1675 B.n619 B.n618 10.6151
R1676 B.n618 B.n617 10.6151
R1677 B.n617 B.n166 10.6151
R1678 B.n613 B.n166 10.6151
R1679 B.n613 B.n612 10.6151
R1680 B.n612 B.n611 10.6151
R1681 B.n611 B.n168 10.6151
R1682 B.n607 B.n168 10.6151
R1683 B.n607 B.n606 10.6151
R1684 B.n606 B.n605 10.6151
R1685 B.n605 B.n170 10.6151
R1686 B.n601 B.n170 10.6151
R1687 B.n601 B.n600 10.6151
R1688 B.n600 B.n599 10.6151
R1689 B.n599 B.n172 10.6151
R1690 B.n595 B.n172 10.6151
R1691 B.n595 B.n594 10.6151
R1692 B.n594 B.n593 10.6151
R1693 B.n593 B.n174 10.6151
R1694 B.n589 B.n174 10.6151
R1695 B.n589 B.n588 10.6151
R1696 B.n588 B.n587 10.6151
R1697 B.n587 B.n176 10.6151
R1698 B.n583 B.n176 10.6151
R1699 B.n583 B.n582 10.6151
R1700 B.n582 B.n581 10.6151
R1701 B.n581 B.n178 10.6151
R1702 B.n577 B.n178 10.6151
R1703 B.n577 B.n576 10.6151
R1704 B.n576 B.n575 10.6151
R1705 B.n575 B.n180 10.6151
R1706 B.n571 B.n180 10.6151
R1707 B.n279 B.n1 10.6151
R1708 B.n279 B.n278 10.6151
R1709 B.n283 B.n278 10.6151
R1710 B.n284 B.n283 10.6151
R1711 B.n285 B.n284 10.6151
R1712 B.n285 B.n276 10.6151
R1713 B.n289 B.n276 10.6151
R1714 B.n290 B.n289 10.6151
R1715 B.n291 B.n290 10.6151
R1716 B.n291 B.n274 10.6151
R1717 B.n295 B.n274 10.6151
R1718 B.n296 B.n295 10.6151
R1719 B.n297 B.n296 10.6151
R1720 B.n297 B.n272 10.6151
R1721 B.n301 B.n272 10.6151
R1722 B.n302 B.n301 10.6151
R1723 B.n303 B.n302 10.6151
R1724 B.n303 B.n270 10.6151
R1725 B.n307 B.n270 10.6151
R1726 B.n308 B.n307 10.6151
R1727 B.n309 B.n308 10.6151
R1728 B.n309 B.n268 10.6151
R1729 B.n313 B.n268 10.6151
R1730 B.n314 B.n313 10.6151
R1731 B.n315 B.n314 10.6151
R1732 B.n315 B.n266 10.6151
R1733 B.n319 B.n266 10.6151
R1734 B.n320 B.n319 10.6151
R1735 B.n321 B.n320 10.6151
R1736 B.n321 B.n264 10.6151
R1737 B.n325 B.n264 10.6151
R1738 B.n326 B.n325 10.6151
R1739 B.n327 B.n326 10.6151
R1740 B.n327 B.n262 10.6151
R1741 B.n331 B.n262 10.6151
R1742 B.n332 B.n331 10.6151
R1743 B.n333 B.n332 10.6151
R1744 B.n333 B.n260 10.6151
R1745 B.n337 B.n260 10.6151
R1746 B.n338 B.n337 10.6151
R1747 B.n339 B.n338 10.6151
R1748 B.n339 B.n258 10.6151
R1749 B.n343 B.n258 10.6151
R1750 B.n344 B.n343 10.6151
R1751 B.n345 B.n344 10.6151
R1752 B.n345 B.n256 10.6151
R1753 B.n349 B.n256 10.6151
R1754 B.n350 B.n349 10.6151
R1755 B.n351 B.n350 10.6151
R1756 B.n351 B.n254 10.6151
R1757 B.n355 B.n254 10.6151
R1758 B.n356 B.n355 10.6151
R1759 B.n357 B.n356 10.6151
R1760 B.n357 B.n252 10.6151
R1761 B.n361 B.n252 10.6151
R1762 B.n362 B.n361 10.6151
R1763 B.n363 B.n362 10.6151
R1764 B.n363 B.n250 10.6151
R1765 B.n367 B.n250 10.6151
R1766 B.n368 B.n367 10.6151
R1767 B.n369 B.n368 10.6151
R1768 B.n369 B.n248 10.6151
R1769 B.n373 B.n248 10.6151
R1770 B.n374 B.n373 10.6151
R1771 B.n375 B.n374 10.6151
R1772 B.n375 B.n246 10.6151
R1773 B.n379 B.n246 10.6151
R1774 B.n380 B.n379 10.6151
R1775 B.n381 B.n380 10.6151
R1776 B.n381 B.n244 10.6151
R1777 B.n385 B.n244 10.6151
R1778 B.n386 B.n385 10.6151
R1779 B.n387 B.n386 10.6151
R1780 B.n387 B.n242 10.6151
R1781 B.n391 B.n242 10.6151
R1782 B.n392 B.n391 10.6151
R1783 B.n393 B.n240 10.6151
R1784 B.n397 B.n240 10.6151
R1785 B.n398 B.n397 10.6151
R1786 B.n399 B.n398 10.6151
R1787 B.n399 B.n238 10.6151
R1788 B.n403 B.n238 10.6151
R1789 B.n404 B.n403 10.6151
R1790 B.n405 B.n404 10.6151
R1791 B.n405 B.n236 10.6151
R1792 B.n409 B.n236 10.6151
R1793 B.n410 B.n409 10.6151
R1794 B.n411 B.n410 10.6151
R1795 B.n411 B.n234 10.6151
R1796 B.n415 B.n234 10.6151
R1797 B.n416 B.n415 10.6151
R1798 B.n417 B.n416 10.6151
R1799 B.n417 B.n232 10.6151
R1800 B.n421 B.n232 10.6151
R1801 B.n422 B.n421 10.6151
R1802 B.n423 B.n422 10.6151
R1803 B.n423 B.n230 10.6151
R1804 B.n427 B.n230 10.6151
R1805 B.n428 B.n427 10.6151
R1806 B.n429 B.n428 10.6151
R1807 B.n429 B.n228 10.6151
R1808 B.n433 B.n228 10.6151
R1809 B.n434 B.n433 10.6151
R1810 B.n435 B.n434 10.6151
R1811 B.n435 B.n226 10.6151
R1812 B.n439 B.n226 10.6151
R1813 B.n440 B.n439 10.6151
R1814 B.n441 B.n440 10.6151
R1815 B.n441 B.n224 10.6151
R1816 B.n445 B.n224 10.6151
R1817 B.n446 B.n445 10.6151
R1818 B.n447 B.n446 10.6151
R1819 B.n447 B.n222 10.6151
R1820 B.n451 B.n222 10.6151
R1821 B.n452 B.n451 10.6151
R1822 B.n453 B.n452 10.6151
R1823 B.n453 B.n220 10.6151
R1824 B.n457 B.n220 10.6151
R1825 B.n458 B.n457 10.6151
R1826 B.n459 B.n458 10.6151
R1827 B.n459 B.n218 10.6151
R1828 B.n463 B.n218 10.6151
R1829 B.n464 B.n463 10.6151
R1830 B.n465 B.n464 10.6151
R1831 B.n465 B.n216 10.6151
R1832 B.n469 B.n216 10.6151
R1833 B.n470 B.n469 10.6151
R1834 B.n474 B.n470 10.6151
R1835 B.n478 B.n214 10.6151
R1836 B.n479 B.n478 10.6151
R1837 B.n480 B.n479 10.6151
R1838 B.n480 B.n212 10.6151
R1839 B.n484 B.n212 10.6151
R1840 B.n485 B.n484 10.6151
R1841 B.n486 B.n485 10.6151
R1842 B.n486 B.n210 10.6151
R1843 B.n490 B.n210 10.6151
R1844 B.n493 B.n492 10.6151
R1845 B.n493 B.n206 10.6151
R1846 B.n497 B.n206 10.6151
R1847 B.n498 B.n497 10.6151
R1848 B.n499 B.n498 10.6151
R1849 B.n499 B.n204 10.6151
R1850 B.n503 B.n204 10.6151
R1851 B.n504 B.n503 10.6151
R1852 B.n505 B.n504 10.6151
R1853 B.n505 B.n202 10.6151
R1854 B.n509 B.n202 10.6151
R1855 B.n510 B.n509 10.6151
R1856 B.n511 B.n510 10.6151
R1857 B.n511 B.n200 10.6151
R1858 B.n515 B.n200 10.6151
R1859 B.n516 B.n515 10.6151
R1860 B.n517 B.n516 10.6151
R1861 B.n517 B.n198 10.6151
R1862 B.n521 B.n198 10.6151
R1863 B.n522 B.n521 10.6151
R1864 B.n523 B.n522 10.6151
R1865 B.n523 B.n196 10.6151
R1866 B.n527 B.n196 10.6151
R1867 B.n528 B.n527 10.6151
R1868 B.n529 B.n528 10.6151
R1869 B.n529 B.n194 10.6151
R1870 B.n533 B.n194 10.6151
R1871 B.n534 B.n533 10.6151
R1872 B.n535 B.n534 10.6151
R1873 B.n535 B.n192 10.6151
R1874 B.n539 B.n192 10.6151
R1875 B.n540 B.n539 10.6151
R1876 B.n541 B.n540 10.6151
R1877 B.n541 B.n190 10.6151
R1878 B.n545 B.n190 10.6151
R1879 B.n546 B.n545 10.6151
R1880 B.n547 B.n546 10.6151
R1881 B.n547 B.n188 10.6151
R1882 B.n551 B.n188 10.6151
R1883 B.n552 B.n551 10.6151
R1884 B.n553 B.n552 10.6151
R1885 B.n553 B.n186 10.6151
R1886 B.n557 B.n186 10.6151
R1887 B.n558 B.n557 10.6151
R1888 B.n559 B.n558 10.6151
R1889 B.n559 B.n184 10.6151
R1890 B.n563 B.n184 10.6151
R1891 B.n564 B.n563 10.6151
R1892 B.n565 B.n564 10.6151
R1893 B.n565 B.n182 10.6151
R1894 B.n569 B.n182 10.6151
R1895 B.n570 B.n569 10.6151
R1896 B.n901 B.n900 9.36635
R1897 B.n883 B.n76 9.36635
R1898 B.n474 B.n473 9.36635
R1899 B.n492 B.n491 9.36635
R1900 B.n1097 B.n0 8.11757
R1901 B.n1097 B.n1 8.11757
R1902 B.n900 B.n899 1.24928
R1903 B.n886 B.n76 1.24928
R1904 B.n473 B.n214 1.24928
R1905 B.n491 B.n490 1.24928
R1906 VN.n106 VN.n105 161.3
R1907 VN.n104 VN.n55 161.3
R1908 VN.n103 VN.n102 161.3
R1909 VN.n101 VN.n56 161.3
R1910 VN.n100 VN.n99 161.3
R1911 VN.n98 VN.n57 161.3
R1912 VN.n97 VN.n96 161.3
R1913 VN.n95 VN.n58 161.3
R1914 VN.n94 VN.n93 161.3
R1915 VN.n92 VN.n59 161.3
R1916 VN.n91 VN.n90 161.3
R1917 VN.n89 VN.n61 161.3
R1918 VN.n88 VN.n87 161.3
R1919 VN.n86 VN.n62 161.3
R1920 VN.n85 VN.n84 161.3
R1921 VN.n83 VN.n63 161.3
R1922 VN.n82 VN.n81 161.3
R1923 VN.n80 VN.n64 161.3
R1924 VN.n79 VN.n78 161.3
R1925 VN.n77 VN.n66 161.3
R1926 VN.n76 VN.n75 161.3
R1927 VN.n74 VN.n67 161.3
R1928 VN.n73 VN.n72 161.3
R1929 VN.n71 VN.n68 161.3
R1930 VN.n52 VN.n51 161.3
R1931 VN.n50 VN.n1 161.3
R1932 VN.n49 VN.n48 161.3
R1933 VN.n47 VN.n2 161.3
R1934 VN.n46 VN.n45 161.3
R1935 VN.n44 VN.n3 161.3
R1936 VN.n43 VN.n42 161.3
R1937 VN.n41 VN.n4 161.3
R1938 VN.n40 VN.n39 161.3
R1939 VN.n37 VN.n5 161.3
R1940 VN.n36 VN.n35 161.3
R1941 VN.n34 VN.n6 161.3
R1942 VN.n33 VN.n32 161.3
R1943 VN.n31 VN.n7 161.3
R1944 VN.n30 VN.n29 161.3
R1945 VN.n28 VN.n8 161.3
R1946 VN.n27 VN.n26 161.3
R1947 VN.n24 VN.n9 161.3
R1948 VN.n23 VN.n22 161.3
R1949 VN.n21 VN.n10 161.3
R1950 VN.n20 VN.n19 161.3
R1951 VN.n18 VN.n11 161.3
R1952 VN.n17 VN.n16 161.3
R1953 VN.n15 VN.n12 161.3
R1954 VN.n70 VN.t3 139.361
R1955 VN.n14 VN.t5 139.361
R1956 VN.n13 VN.t8 106.547
R1957 VN.n25 VN.t2 106.547
R1958 VN.n38 VN.t1 106.547
R1959 VN.n0 VN.t0 106.547
R1960 VN.n69 VN.t9 106.547
R1961 VN.n65 VN.t4 106.547
R1962 VN.n60 VN.t6 106.547
R1963 VN.n54 VN.t7 106.547
R1964 VN.n53 VN.n0 83.8517
R1965 VN.n107 VN.n54 83.8517
R1966 VN.n14 VN.n13 65.3998
R1967 VN.n70 VN.n69 65.3998
R1968 VN VN.n107 61.8315
R1969 VN.n19 VN.n10 56.5617
R1970 VN.n32 VN.n6 56.5617
R1971 VN.n75 VN.n66 56.5617
R1972 VN.n87 VN.n61 56.5617
R1973 VN.n45 VN.n2 56.0773
R1974 VN.n99 VN.n56 56.0773
R1975 VN.n45 VN.n44 25.0767
R1976 VN.n99 VN.n98 25.0767
R1977 VN.n17 VN.n12 24.5923
R1978 VN.n18 VN.n17 24.5923
R1979 VN.n19 VN.n18 24.5923
R1980 VN.n23 VN.n10 24.5923
R1981 VN.n24 VN.n23 24.5923
R1982 VN.n26 VN.n24 24.5923
R1983 VN.n30 VN.n8 24.5923
R1984 VN.n31 VN.n30 24.5923
R1985 VN.n32 VN.n31 24.5923
R1986 VN.n36 VN.n6 24.5923
R1987 VN.n37 VN.n36 24.5923
R1988 VN.n39 VN.n37 24.5923
R1989 VN.n43 VN.n4 24.5923
R1990 VN.n44 VN.n43 24.5923
R1991 VN.n49 VN.n2 24.5923
R1992 VN.n50 VN.n49 24.5923
R1993 VN.n51 VN.n50 24.5923
R1994 VN.n75 VN.n74 24.5923
R1995 VN.n74 VN.n73 24.5923
R1996 VN.n73 VN.n68 24.5923
R1997 VN.n87 VN.n86 24.5923
R1998 VN.n86 VN.n85 24.5923
R1999 VN.n85 VN.n63 24.5923
R2000 VN.n81 VN.n80 24.5923
R2001 VN.n80 VN.n79 24.5923
R2002 VN.n79 VN.n66 24.5923
R2003 VN.n98 VN.n97 24.5923
R2004 VN.n97 VN.n58 24.5923
R2005 VN.n93 VN.n92 24.5923
R2006 VN.n92 VN.n91 24.5923
R2007 VN.n91 VN.n61 24.5923
R2008 VN.n105 VN.n104 24.5923
R2009 VN.n104 VN.n103 24.5923
R2010 VN.n103 VN.n56 24.5923
R2011 VN.n38 VN.n4 15.2474
R2012 VN.n60 VN.n58 15.2474
R2013 VN.n26 VN.n25 12.2964
R2014 VN.n25 VN.n8 12.2964
R2015 VN.n65 VN.n63 12.2964
R2016 VN.n81 VN.n65 12.2964
R2017 VN.n13 VN.n12 9.3454
R2018 VN.n39 VN.n38 9.3454
R2019 VN.n69 VN.n68 9.3454
R2020 VN.n93 VN.n60 9.3454
R2021 VN.n51 VN.n0 6.39438
R2022 VN.n105 VN.n54 6.39438
R2023 VN.n71 VN.n70 3.2619
R2024 VN.n15 VN.n14 3.2619
R2025 VN.n107 VN.n106 0.354861
R2026 VN.n53 VN.n52 0.354861
R2027 VN VN.n53 0.267071
R2028 VN.n106 VN.n55 0.189894
R2029 VN.n102 VN.n55 0.189894
R2030 VN.n102 VN.n101 0.189894
R2031 VN.n101 VN.n100 0.189894
R2032 VN.n100 VN.n57 0.189894
R2033 VN.n96 VN.n57 0.189894
R2034 VN.n96 VN.n95 0.189894
R2035 VN.n95 VN.n94 0.189894
R2036 VN.n94 VN.n59 0.189894
R2037 VN.n90 VN.n59 0.189894
R2038 VN.n90 VN.n89 0.189894
R2039 VN.n89 VN.n88 0.189894
R2040 VN.n88 VN.n62 0.189894
R2041 VN.n84 VN.n62 0.189894
R2042 VN.n84 VN.n83 0.189894
R2043 VN.n83 VN.n82 0.189894
R2044 VN.n82 VN.n64 0.189894
R2045 VN.n78 VN.n64 0.189894
R2046 VN.n78 VN.n77 0.189894
R2047 VN.n77 VN.n76 0.189894
R2048 VN.n76 VN.n67 0.189894
R2049 VN.n72 VN.n67 0.189894
R2050 VN.n72 VN.n71 0.189894
R2051 VN.n16 VN.n15 0.189894
R2052 VN.n16 VN.n11 0.189894
R2053 VN.n20 VN.n11 0.189894
R2054 VN.n21 VN.n20 0.189894
R2055 VN.n22 VN.n21 0.189894
R2056 VN.n22 VN.n9 0.189894
R2057 VN.n27 VN.n9 0.189894
R2058 VN.n28 VN.n27 0.189894
R2059 VN.n29 VN.n28 0.189894
R2060 VN.n29 VN.n7 0.189894
R2061 VN.n33 VN.n7 0.189894
R2062 VN.n34 VN.n33 0.189894
R2063 VN.n35 VN.n34 0.189894
R2064 VN.n35 VN.n5 0.189894
R2065 VN.n40 VN.n5 0.189894
R2066 VN.n41 VN.n40 0.189894
R2067 VN.n42 VN.n41 0.189894
R2068 VN.n42 VN.n3 0.189894
R2069 VN.n46 VN.n3 0.189894
R2070 VN.n47 VN.n46 0.189894
R2071 VN.n48 VN.n47 0.189894
R2072 VN.n48 VN.n1 0.189894
R2073 VN.n52 VN.n1 0.189894
R2074 VDD2.n1 VDD2.t4 73.4065
R2075 VDD2.n3 VDD2.n2 70.4654
R2076 VDD2 VDD2.n7 70.4628
R2077 VDD2.n4 VDD2.t2 70.0102
R2078 VDD2.n6 VDD2.n5 67.9736
R2079 VDD2.n1 VDD2.n0 67.9733
R2080 VDD2.n4 VDD2.n3 53.6075
R2081 VDD2.n6 VDD2.n4 3.39705
R2082 VDD2.n7 VDD2.t0 2.03715
R2083 VDD2.n7 VDD2.t6 2.03715
R2084 VDD2.n5 VDD2.t3 2.03715
R2085 VDD2.n5 VDD2.t5 2.03715
R2086 VDD2.n2 VDD2.t8 2.03715
R2087 VDD2.n2 VDD2.t9 2.03715
R2088 VDD2.n0 VDD2.t1 2.03715
R2089 VDD2.n0 VDD2.t7 2.03715
R2090 VDD2 VDD2.n6 0.907828
R2091 VDD2.n3 VDD2.n1 0.794292
C0 VDD2 VDD1 2.83383f
C1 VN VP 10.6139f
C2 VN w_n5698_n4160# 12.550099f
C3 VN B 1.59143f
C4 VN VDD1 0.156161f
C5 VN VDD2 14.831699f
C6 VTAIL VP 15.7336f
C7 VTAIL w_n5698_n4160# 3.89695f
C8 w_n5698_n4160# VP 13.295f
C9 VTAIL B 5.05414f
C10 VP B 2.8497f
C11 w_n5698_n4160# B 13.355f
C12 VTAIL VDD1 12.4436f
C13 VP VDD1 15.3842f
C14 w_n5698_n4160# VDD1 3.44437f
C15 VDD1 B 3.19197f
C16 VTAIL VDD2 12.5015f
C17 VDD2 VP 0.713045f
C18 VDD2 w_n5698_n4160# 3.64042f
C19 VDD2 B 3.34921f
C20 VN VTAIL 15.7191f
C21 VDD2 VSUBS 2.62159f
C22 VDD1 VSUBS 2.474092f
C23 VTAIL VSUBS 1.674251f
C24 VN VSUBS 9.48722f
C25 VP VSUBS 5.669117f
C26 B VSUBS 6.952431f
C27 w_n5698_n4160# VSUBS 0.290393p
C28 VDD2.t4 VSUBS 3.97035f
C29 VDD2.t1 VSUBS 0.371547f
C30 VDD2.t7 VSUBS 0.371547f
C31 VDD2.n0 VSUBS 3.01553f
C32 VDD2.n1 VSUBS 1.98093f
C33 VDD2.t8 VSUBS 0.371547f
C34 VDD2.t9 VSUBS 0.371547f
C35 VDD2.n2 VSUBS 3.05676f
C36 VDD2.n3 VSUBS 4.678f
C37 VDD2.t2 VSUBS 3.92245f
C38 VDD2.n4 VSUBS 4.88147f
C39 VDD2.t3 VSUBS 0.371547f
C40 VDD2.t5 VSUBS 0.371547f
C41 VDD2.n5 VSUBS 3.01553f
C42 VDD2.n6 VSUBS 1.00331f
C43 VDD2.t0 VSUBS 0.371547f
C44 VDD2.t6 VSUBS 0.371547f
C45 VDD2.n7 VSUBS 3.0567f
C46 VN.t0 VSUBS 3.42561f
C47 VN.n0 VSUBS 1.26698f
C48 VN.n1 VSUBS 0.021668f
C49 VN.n2 VSUBS 0.03684f
C50 VN.n3 VSUBS 0.021668f
C51 VN.n4 VSUBS 0.032644f
C52 VN.n5 VSUBS 0.021668f
C53 VN.n6 VSUBS 0.033297f
C54 VN.n7 VSUBS 0.021668f
C55 VN.n8 VSUBS 0.030263f
C56 VN.n9 VSUBS 0.021668f
C57 VN.n10 VSUBS 0.0297f
C58 VN.n11 VSUBS 0.021668f
C59 VN.n12 VSUBS 0.027883f
C60 VN.t8 VSUBS 3.42561f
C61 VN.n13 VSUBS 1.25857f
C62 VN.t5 VSUBS 3.7432f
C63 VN.n14 VSUBS 1.20121f
C64 VN.n15 VSUBS 0.27167f
C65 VN.n16 VSUBS 0.021668f
C66 VN.n17 VSUBS 0.040182f
C67 VN.n18 VSUBS 0.040182f
C68 VN.n19 VSUBS 0.033297f
C69 VN.n20 VSUBS 0.021668f
C70 VN.n21 VSUBS 0.021668f
C71 VN.n22 VSUBS 0.021668f
C72 VN.n23 VSUBS 0.040182f
C73 VN.n24 VSUBS 0.040182f
C74 VN.t2 VSUBS 3.42561f
C75 VN.n25 VSUBS 1.18607f
C76 VN.n26 VSUBS 0.030263f
C77 VN.n27 VSUBS 0.021668f
C78 VN.n28 VSUBS 0.021668f
C79 VN.n29 VSUBS 0.021668f
C80 VN.n30 VSUBS 0.040182f
C81 VN.n31 VSUBS 0.040182f
C82 VN.n32 VSUBS 0.0297f
C83 VN.n33 VSUBS 0.021668f
C84 VN.n34 VSUBS 0.021668f
C85 VN.n35 VSUBS 0.021668f
C86 VN.n36 VSUBS 0.040182f
C87 VN.n37 VSUBS 0.040182f
C88 VN.t1 VSUBS 3.42561f
C89 VN.n38 VSUBS 1.18607f
C90 VN.n39 VSUBS 0.027883f
C91 VN.n40 VSUBS 0.021668f
C92 VN.n41 VSUBS 0.021668f
C93 VN.n42 VSUBS 0.021668f
C94 VN.n43 VSUBS 0.040182f
C95 VN.n44 VSUBS 0.040557f
C96 VN.n45 VSUBS 0.02578f
C97 VN.n46 VSUBS 0.021668f
C98 VN.n47 VSUBS 0.021668f
C99 VN.n48 VSUBS 0.021668f
C100 VN.n49 VSUBS 0.040182f
C101 VN.n50 VSUBS 0.040182f
C102 VN.n51 VSUBS 0.025503f
C103 VN.n52 VSUBS 0.034967f
C104 VN.n53 VSUBS 0.061957f
C105 VN.t7 VSUBS 3.42561f
C106 VN.n54 VSUBS 1.26698f
C107 VN.n55 VSUBS 0.021668f
C108 VN.n56 VSUBS 0.03684f
C109 VN.n57 VSUBS 0.021668f
C110 VN.n58 VSUBS 0.032644f
C111 VN.n59 VSUBS 0.021668f
C112 VN.t6 VSUBS 3.42561f
C113 VN.n60 VSUBS 1.18607f
C114 VN.n61 VSUBS 0.033297f
C115 VN.n62 VSUBS 0.021668f
C116 VN.n63 VSUBS 0.030263f
C117 VN.n64 VSUBS 0.021668f
C118 VN.t4 VSUBS 3.42561f
C119 VN.n65 VSUBS 1.18607f
C120 VN.n66 VSUBS 0.0297f
C121 VN.n67 VSUBS 0.021668f
C122 VN.n68 VSUBS 0.027883f
C123 VN.t3 VSUBS 3.7432f
C124 VN.t9 VSUBS 3.42561f
C125 VN.n69 VSUBS 1.25857f
C126 VN.n70 VSUBS 1.20121f
C127 VN.n71 VSUBS 0.27167f
C128 VN.n72 VSUBS 0.021668f
C129 VN.n73 VSUBS 0.040182f
C130 VN.n74 VSUBS 0.040182f
C131 VN.n75 VSUBS 0.033297f
C132 VN.n76 VSUBS 0.021668f
C133 VN.n77 VSUBS 0.021668f
C134 VN.n78 VSUBS 0.021668f
C135 VN.n79 VSUBS 0.040182f
C136 VN.n80 VSUBS 0.040182f
C137 VN.n81 VSUBS 0.030263f
C138 VN.n82 VSUBS 0.021668f
C139 VN.n83 VSUBS 0.021668f
C140 VN.n84 VSUBS 0.021668f
C141 VN.n85 VSUBS 0.040182f
C142 VN.n86 VSUBS 0.040182f
C143 VN.n87 VSUBS 0.0297f
C144 VN.n88 VSUBS 0.021668f
C145 VN.n89 VSUBS 0.021668f
C146 VN.n90 VSUBS 0.021668f
C147 VN.n91 VSUBS 0.040182f
C148 VN.n92 VSUBS 0.040182f
C149 VN.n93 VSUBS 0.027883f
C150 VN.n94 VSUBS 0.021668f
C151 VN.n95 VSUBS 0.021668f
C152 VN.n96 VSUBS 0.021668f
C153 VN.n97 VSUBS 0.040182f
C154 VN.n98 VSUBS 0.040557f
C155 VN.n99 VSUBS 0.02578f
C156 VN.n100 VSUBS 0.021668f
C157 VN.n101 VSUBS 0.021668f
C158 VN.n102 VSUBS 0.021668f
C159 VN.n103 VSUBS 0.040182f
C160 VN.n104 VSUBS 0.040182f
C161 VN.n105 VSUBS 0.025503f
C162 VN.n106 VSUBS 0.034967f
C163 VN.n107 VSUBS 1.66322f
C164 B.n0 VSUBS 0.007035f
C165 B.n1 VSUBS 0.007035f
C166 B.n2 VSUBS 0.010405f
C167 B.n3 VSUBS 0.007973f
C168 B.n4 VSUBS 0.007973f
C169 B.n5 VSUBS 0.007973f
C170 B.n6 VSUBS 0.007973f
C171 B.n7 VSUBS 0.007973f
C172 B.n8 VSUBS 0.007973f
C173 B.n9 VSUBS 0.007973f
C174 B.n10 VSUBS 0.007973f
C175 B.n11 VSUBS 0.007973f
C176 B.n12 VSUBS 0.007973f
C177 B.n13 VSUBS 0.007973f
C178 B.n14 VSUBS 0.007973f
C179 B.n15 VSUBS 0.007973f
C180 B.n16 VSUBS 0.007973f
C181 B.n17 VSUBS 0.007973f
C182 B.n18 VSUBS 0.007973f
C183 B.n19 VSUBS 0.007973f
C184 B.n20 VSUBS 0.007973f
C185 B.n21 VSUBS 0.007973f
C186 B.n22 VSUBS 0.007973f
C187 B.n23 VSUBS 0.007973f
C188 B.n24 VSUBS 0.007973f
C189 B.n25 VSUBS 0.007973f
C190 B.n26 VSUBS 0.007973f
C191 B.n27 VSUBS 0.007973f
C192 B.n28 VSUBS 0.007973f
C193 B.n29 VSUBS 0.007973f
C194 B.n30 VSUBS 0.007973f
C195 B.n31 VSUBS 0.007973f
C196 B.n32 VSUBS 0.007973f
C197 B.n33 VSUBS 0.007973f
C198 B.n34 VSUBS 0.007973f
C199 B.n35 VSUBS 0.007973f
C200 B.n36 VSUBS 0.007973f
C201 B.n37 VSUBS 0.007973f
C202 B.n38 VSUBS 0.007973f
C203 B.n39 VSUBS 0.007973f
C204 B.n40 VSUBS 0.018858f
C205 B.n41 VSUBS 0.007973f
C206 B.n42 VSUBS 0.007973f
C207 B.n43 VSUBS 0.007973f
C208 B.n44 VSUBS 0.007973f
C209 B.n45 VSUBS 0.007973f
C210 B.n46 VSUBS 0.007973f
C211 B.n47 VSUBS 0.007973f
C212 B.n48 VSUBS 0.007973f
C213 B.n49 VSUBS 0.007973f
C214 B.n50 VSUBS 0.007973f
C215 B.n51 VSUBS 0.007973f
C216 B.n52 VSUBS 0.007973f
C217 B.n53 VSUBS 0.007973f
C218 B.n54 VSUBS 0.007973f
C219 B.n55 VSUBS 0.007973f
C220 B.n56 VSUBS 0.007973f
C221 B.n57 VSUBS 0.007973f
C222 B.n58 VSUBS 0.007973f
C223 B.n59 VSUBS 0.007973f
C224 B.n60 VSUBS 0.007973f
C225 B.n61 VSUBS 0.007973f
C226 B.n62 VSUBS 0.007973f
C227 B.n63 VSUBS 0.007973f
C228 B.n64 VSUBS 0.007973f
C229 B.n65 VSUBS 0.007973f
C230 B.n66 VSUBS 0.007973f
C231 B.n67 VSUBS 0.007973f
C232 B.t1 VSUBS 0.608284f
C233 B.t2 VSUBS 0.638769f
C234 B.t0 VSUBS 3.00239f
C235 B.n68 VSUBS 0.381452f
C236 B.n69 VSUBS 0.086787f
C237 B.n70 VSUBS 0.007973f
C238 B.n71 VSUBS 0.007973f
C239 B.n72 VSUBS 0.007973f
C240 B.n73 VSUBS 0.007973f
C241 B.t4 VSUBS 0.608266f
C242 B.t5 VSUBS 0.638755f
C243 B.t3 VSUBS 3.00239f
C244 B.n74 VSUBS 0.381466f
C245 B.n75 VSUBS 0.086806f
C246 B.n76 VSUBS 0.018473f
C247 B.n77 VSUBS 0.007973f
C248 B.n78 VSUBS 0.007973f
C249 B.n79 VSUBS 0.007973f
C250 B.n80 VSUBS 0.007973f
C251 B.n81 VSUBS 0.007973f
C252 B.n82 VSUBS 0.007973f
C253 B.n83 VSUBS 0.007973f
C254 B.n84 VSUBS 0.007973f
C255 B.n85 VSUBS 0.007973f
C256 B.n86 VSUBS 0.007973f
C257 B.n87 VSUBS 0.007973f
C258 B.n88 VSUBS 0.007973f
C259 B.n89 VSUBS 0.007973f
C260 B.n90 VSUBS 0.007973f
C261 B.n91 VSUBS 0.007973f
C262 B.n92 VSUBS 0.007973f
C263 B.n93 VSUBS 0.007973f
C264 B.n94 VSUBS 0.007973f
C265 B.n95 VSUBS 0.007973f
C266 B.n96 VSUBS 0.007973f
C267 B.n97 VSUBS 0.007973f
C268 B.n98 VSUBS 0.007973f
C269 B.n99 VSUBS 0.007973f
C270 B.n100 VSUBS 0.007973f
C271 B.n101 VSUBS 0.007973f
C272 B.n102 VSUBS 0.007973f
C273 B.n103 VSUBS 0.018858f
C274 B.n104 VSUBS 0.007973f
C275 B.n105 VSUBS 0.007973f
C276 B.n106 VSUBS 0.007973f
C277 B.n107 VSUBS 0.007973f
C278 B.n108 VSUBS 0.007973f
C279 B.n109 VSUBS 0.007973f
C280 B.n110 VSUBS 0.007973f
C281 B.n111 VSUBS 0.007973f
C282 B.n112 VSUBS 0.007973f
C283 B.n113 VSUBS 0.007973f
C284 B.n114 VSUBS 0.007973f
C285 B.n115 VSUBS 0.007973f
C286 B.n116 VSUBS 0.007973f
C287 B.n117 VSUBS 0.007973f
C288 B.n118 VSUBS 0.007973f
C289 B.n119 VSUBS 0.007973f
C290 B.n120 VSUBS 0.007973f
C291 B.n121 VSUBS 0.007973f
C292 B.n122 VSUBS 0.007973f
C293 B.n123 VSUBS 0.007973f
C294 B.n124 VSUBS 0.007973f
C295 B.n125 VSUBS 0.007973f
C296 B.n126 VSUBS 0.007973f
C297 B.n127 VSUBS 0.007973f
C298 B.n128 VSUBS 0.007973f
C299 B.n129 VSUBS 0.007973f
C300 B.n130 VSUBS 0.007973f
C301 B.n131 VSUBS 0.007973f
C302 B.n132 VSUBS 0.007973f
C303 B.n133 VSUBS 0.007973f
C304 B.n134 VSUBS 0.007973f
C305 B.n135 VSUBS 0.007973f
C306 B.n136 VSUBS 0.007973f
C307 B.n137 VSUBS 0.007973f
C308 B.n138 VSUBS 0.007973f
C309 B.n139 VSUBS 0.007973f
C310 B.n140 VSUBS 0.007973f
C311 B.n141 VSUBS 0.007973f
C312 B.n142 VSUBS 0.007973f
C313 B.n143 VSUBS 0.007973f
C314 B.n144 VSUBS 0.007973f
C315 B.n145 VSUBS 0.007973f
C316 B.n146 VSUBS 0.007973f
C317 B.n147 VSUBS 0.007973f
C318 B.n148 VSUBS 0.007973f
C319 B.n149 VSUBS 0.007973f
C320 B.n150 VSUBS 0.007973f
C321 B.n151 VSUBS 0.007973f
C322 B.n152 VSUBS 0.007973f
C323 B.n153 VSUBS 0.007973f
C324 B.n154 VSUBS 0.007973f
C325 B.n155 VSUBS 0.007973f
C326 B.n156 VSUBS 0.007973f
C327 B.n157 VSUBS 0.007973f
C328 B.n158 VSUBS 0.007973f
C329 B.n159 VSUBS 0.007973f
C330 B.n160 VSUBS 0.007973f
C331 B.n161 VSUBS 0.007973f
C332 B.n162 VSUBS 0.007973f
C333 B.n163 VSUBS 0.007973f
C334 B.n164 VSUBS 0.007973f
C335 B.n165 VSUBS 0.007973f
C336 B.n166 VSUBS 0.007973f
C337 B.n167 VSUBS 0.007973f
C338 B.n168 VSUBS 0.007973f
C339 B.n169 VSUBS 0.007973f
C340 B.n170 VSUBS 0.007973f
C341 B.n171 VSUBS 0.007973f
C342 B.n172 VSUBS 0.007973f
C343 B.n173 VSUBS 0.007973f
C344 B.n174 VSUBS 0.007973f
C345 B.n175 VSUBS 0.007973f
C346 B.n176 VSUBS 0.007973f
C347 B.n177 VSUBS 0.007973f
C348 B.n178 VSUBS 0.007973f
C349 B.n179 VSUBS 0.007973f
C350 B.n180 VSUBS 0.007973f
C351 B.n181 VSUBS 0.019837f
C352 B.n182 VSUBS 0.007973f
C353 B.n183 VSUBS 0.007973f
C354 B.n184 VSUBS 0.007973f
C355 B.n185 VSUBS 0.007973f
C356 B.n186 VSUBS 0.007973f
C357 B.n187 VSUBS 0.007973f
C358 B.n188 VSUBS 0.007973f
C359 B.n189 VSUBS 0.007973f
C360 B.n190 VSUBS 0.007973f
C361 B.n191 VSUBS 0.007973f
C362 B.n192 VSUBS 0.007973f
C363 B.n193 VSUBS 0.007973f
C364 B.n194 VSUBS 0.007973f
C365 B.n195 VSUBS 0.007973f
C366 B.n196 VSUBS 0.007973f
C367 B.n197 VSUBS 0.007973f
C368 B.n198 VSUBS 0.007973f
C369 B.n199 VSUBS 0.007973f
C370 B.n200 VSUBS 0.007973f
C371 B.n201 VSUBS 0.007973f
C372 B.n202 VSUBS 0.007973f
C373 B.n203 VSUBS 0.007973f
C374 B.n204 VSUBS 0.007973f
C375 B.n205 VSUBS 0.007973f
C376 B.n206 VSUBS 0.007973f
C377 B.n207 VSUBS 0.007973f
C378 B.t11 VSUBS 0.608266f
C379 B.t10 VSUBS 0.638755f
C380 B.t9 VSUBS 3.00239f
C381 B.n208 VSUBS 0.381466f
C382 B.n209 VSUBS 0.086806f
C383 B.n210 VSUBS 0.007973f
C384 B.n211 VSUBS 0.007973f
C385 B.n212 VSUBS 0.007973f
C386 B.n213 VSUBS 0.007973f
C387 B.n214 VSUBS 0.004456f
C388 B.n215 VSUBS 0.007973f
C389 B.n216 VSUBS 0.007973f
C390 B.n217 VSUBS 0.007973f
C391 B.n218 VSUBS 0.007973f
C392 B.n219 VSUBS 0.007973f
C393 B.n220 VSUBS 0.007973f
C394 B.n221 VSUBS 0.007973f
C395 B.n222 VSUBS 0.007973f
C396 B.n223 VSUBS 0.007973f
C397 B.n224 VSUBS 0.007973f
C398 B.n225 VSUBS 0.007973f
C399 B.n226 VSUBS 0.007973f
C400 B.n227 VSUBS 0.007973f
C401 B.n228 VSUBS 0.007973f
C402 B.n229 VSUBS 0.007973f
C403 B.n230 VSUBS 0.007973f
C404 B.n231 VSUBS 0.007973f
C405 B.n232 VSUBS 0.007973f
C406 B.n233 VSUBS 0.007973f
C407 B.n234 VSUBS 0.007973f
C408 B.n235 VSUBS 0.007973f
C409 B.n236 VSUBS 0.007973f
C410 B.n237 VSUBS 0.007973f
C411 B.n238 VSUBS 0.007973f
C412 B.n239 VSUBS 0.007973f
C413 B.n240 VSUBS 0.007973f
C414 B.n241 VSUBS 0.018858f
C415 B.n242 VSUBS 0.007973f
C416 B.n243 VSUBS 0.007973f
C417 B.n244 VSUBS 0.007973f
C418 B.n245 VSUBS 0.007973f
C419 B.n246 VSUBS 0.007973f
C420 B.n247 VSUBS 0.007973f
C421 B.n248 VSUBS 0.007973f
C422 B.n249 VSUBS 0.007973f
C423 B.n250 VSUBS 0.007973f
C424 B.n251 VSUBS 0.007973f
C425 B.n252 VSUBS 0.007973f
C426 B.n253 VSUBS 0.007973f
C427 B.n254 VSUBS 0.007973f
C428 B.n255 VSUBS 0.007973f
C429 B.n256 VSUBS 0.007973f
C430 B.n257 VSUBS 0.007973f
C431 B.n258 VSUBS 0.007973f
C432 B.n259 VSUBS 0.007973f
C433 B.n260 VSUBS 0.007973f
C434 B.n261 VSUBS 0.007973f
C435 B.n262 VSUBS 0.007973f
C436 B.n263 VSUBS 0.007973f
C437 B.n264 VSUBS 0.007973f
C438 B.n265 VSUBS 0.007973f
C439 B.n266 VSUBS 0.007973f
C440 B.n267 VSUBS 0.007973f
C441 B.n268 VSUBS 0.007973f
C442 B.n269 VSUBS 0.007973f
C443 B.n270 VSUBS 0.007973f
C444 B.n271 VSUBS 0.007973f
C445 B.n272 VSUBS 0.007973f
C446 B.n273 VSUBS 0.007973f
C447 B.n274 VSUBS 0.007973f
C448 B.n275 VSUBS 0.007973f
C449 B.n276 VSUBS 0.007973f
C450 B.n277 VSUBS 0.007973f
C451 B.n278 VSUBS 0.007973f
C452 B.n279 VSUBS 0.007973f
C453 B.n280 VSUBS 0.007973f
C454 B.n281 VSUBS 0.007973f
C455 B.n282 VSUBS 0.007973f
C456 B.n283 VSUBS 0.007973f
C457 B.n284 VSUBS 0.007973f
C458 B.n285 VSUBS 0.007973f
C459 B.n286 VSUBS 0.007973f
C460 B.n287 VSUBS 0.007973f
C461 B.n288 VSUBS 0.007973f
C462 B.n289 VSUBS 0.007973f
C463 B.n290 VSUBS 0.007973f
C464 B.n291 VSUBS 0.007973f
C465 B.n292 VSUBS 0.007973f
C466 B.n293 VSUBS 0.007973f
C467 B.n294 VSUBS 0.007973f
C468 B.n295 VSUBS 0.007973f
C469 B.n296 VSUBS 0.007973f
C470 B.n297 VSUBS 0.007973f
C471 B.n298 VSUBS 0.007973f
C472 B.n299 VSUBS 0.007973f
C473 B.n300 VSUBS 0.007973f
C474 B.n301 VSUBS 0.007973f
C475 B.n302 VSUBS 0.007973f
C476 B.n303 VSUBS 0.007973f
C477 B.n304 VSUBS 0.007973f
C478 B.n305 VSUBS 0.007973f
C479 B.n306 VSUBS 0.007973f
C480 B.n307 VSUBS 0.007973f
C481 B.n308 VSUBS 0.007973f
C482 B.n309 VSUBS 0.007973f
C483 B.n310 VSUBS 0.007973f
C484 B.n311 VSUBS 0.007973f
C485 B.n312 VSUBS 0.007973f
C486 B.n313 VSUBS 0.007973f
C487 B.n314 VSUBS 0.007973f
C488 B.n315 VSUBS 0.007973f
C489 B.n316 VSUBS 0.007973f
C490 B.n317 VSUBS 0.007973f
C491 B.n318 VSUBS 0.007973f
C492 B.n319 VSUBS 0.007973f
C493 B.n320 VSUBS 0.007973f
C494 B.n321 VSUBS 0.007973f
C495 B.n322 VSUBS 0.007973f
C496 B.n323 VSUBS 0.007973f
C497 B.n324 VSUBS 0.007973f
C498 B.n325 VSUBS 0.007973f
C499 B.n326 VSUBS 0.007973f
C500 B.n327 VSUBS 0.007973f
C501 B.n328 VSUBS 0.007973f
C502 B.n329 VSUBS 0.007973f
C503 B.n330 VSUBS 0.007973f
C504 B.n331 VSUBS 0.007973f
C505 B.n332 VSUBS 0.007973f
C506 B.n333 VSUBS 0.007973f
C507 B.n334 VSUBS 0.007973f
C508 B.n335 VSUBS 0.007973f
C509 B.n336 VSUBS 0.007973f
C510 B.n337 VSUBS 0.007973f
C511 B.n338 VSUBS 0.007973f
C512 B.n339 VSUBS 0.007973f
C513 B.n340 VSUBS 0.007973f
C514 B.n341 VSUBS 0.007973f
C515 B.n342 VSUBS 0.007973f
C516 B.n343 VSUBS 0.007973f
C517 B.n344 VSUBS 0.007973f
C518 B.n345 VSUBS 0.007973f
C519 B.n346 VSUBS 0.007973f
C520 B.n347 VSUBS 0.007973f
C521 B.n348 VSUBS 0.007973f
C522 B.n349 VSUBS 0.007973f
C523 B.n350 VSUBS 0.007973f
C524 B.n351 VSUBS 0.007973f
C525 B.n352 VSUBS 0.007973f
C526 B.n353 VSUBS 0.007973f
C527 B.n354 VSUBS 0.007973f
C528 B.n355 VSUBS 0.007973f
C529 B.n356 VSUBS 0.007973f
C530 B.n357 VSUBS 0.007973f
C531 B.n358 VSUBS 0.007973f
C532 B.n359 VSUBS 0.007973f
C533 B.n360 VSUBS 0.007973f
C534 B.n361 VSUBS 0.007973f
C535 B.n362 VSUBS 0.007973f
C536 B.n363 VSUBS 0.007973f
C537 B.n364 VSUBS 0.007973f
C538 B.n365 VSUBS 0.007973f
C539 B.n366 VSUBS 0.007973f
C540 B.n367 VSUBS 0.007973f
C541 B.n368 VSUBS 0.007973f
C542 B.n369 VSUBS 0.007973f
C543 B.n370 VSUBS 0.007973f
C544 B.n371 VSUBS 0.007973f
C545 B.n372 VSUBS 0.007973f
C546 B.n373 VSUBS 0.007973f
C547 B.n374 VSUBS 0.007973f
C548 B.n375 VSUBS 0.007973f
C549 B.n376 VSUBS 0.007973f
C550 B.n377 VSUBS 0.007973f
C551 B.n378 VSUBS 0.007973f
C552 B.n379 VSUBS 0.007973f
C553 B.n380 VSUBS 0.007973f
C554 B.n381 VSUBS 0.007973f
C555 B.n382 VSUBS 0.007973f
C556 B.n383 VSUBS 0.007973f
C557 B.n384 VSUBS 0.007973f
C558 B.n385 VSUBS 0.007973f
C559 B.n386 VSUBS 0.007973f
C560 B.n387 VSUBS 0.007973f
C561 B.n388 VSUBS 0.007973f
C562 B.n389 VSUBS 0.007973f
C563 B.n390 VSUBS 0.007973f
C564 B.n391 VSUBS 0.007973f
C565 B.n392 VSUBS 0.018858f
C566 B.n393 VSUBS 0.019837f
C567 B.n394 VSUBS 0.019837f
C568 B.n395 VSUBS 0.007973f
C569 B.n396 VSUBS 0.007973f
C570 B.n397 VSUBS 0.007973f
C571 B.n398 VSUBS 0.007973f
C572 B.n399 VSUBS 0.007973f
C573 B.n400 VSUBS 0.007973f
C574 B.n401 VSUBS 0.007973f
C575 B.n402 VSUBS 0.007973f
C576 B.n403 VSUBS 0.007973f
C577 B.n404 VSUBS 0.007973f
C578 B.n405 VSUBS 0.007973f
C579 B.n406 VSUBS 0.007973f
C580 B.n407 VSUBS 0.007973f
C581 B.n408 VSUBS 0.007973f
C582 B.n409 VSUBS 0.007973f
C583 B.n410 VSUBS 0.007973f
C584 B.n411 VSUBS 0.007973f
C585 B.n412 VSUBS 0.007973f
C586 B.n413 VSUBS 0.007973f
C587 B.n414 VSUBS 0.007973f
C588 B.n415 VSUBS 0.007973f
C589 B.n416 VSUBS 0.007973f
C590 B.n417 VSUBS 0.007973f
C591 B.n418 VSUBS 0.007973f
C592 B.n419 VSUBS 0.007973f
C593 B.n420 VSUBS 0.007973f
C594 B.n421 VSUBS 0.007973f
C595 B.n422 VSUBS 0.007973f
C596 B.n423 VSUBS 0.007973f
C597 B.n424 VSUBS 0.007973f
C598 B.n425 VSUBS 0.007973f
C599 B.n426 VSUBS 0.007973f
C600 B.n427 VSUBS 0.007973f
C601 B.n428 VSUBS 0.007973f
C602 B.n429 VSUBS 0.007973f
C603 B.n430 VSUBS 0.007973f
C604 B.n431 VSUBS 0.007973f
C605 B.n432 VSUBS 0.007973f
C606 B.n433 VSUBS 0.007973f
C607 B.n434 VSUBS 0.007973f
C608 B.n435 VSUBS 0.007973f
C609 B.n436 VSUBS 0.007973f
C610 B.n437 VSUBS 0.007973f
C611 B.n438 VSUBS 0.007973f
C612 B.n439 VSUBS 0.007973f
C613 B.n440 VSUBS 0.007973f
C614 B.n441 VSUBS 0.007973f
C615 B.n442 VSUBS 0.007973f
C616 B.n443 VSUBS 0.007973f
C617 B.n444 VSUBS 0.007973f
C618 B.n445 VSUBS 0.007973f
C619 B.n446 VSUBS 0.007973f
C620 B.n447 VSUBS 0.007973f
C621 B.n448 VSUBS 0.007973f
C622 B.n449 VSUBS 0.007973f
C623 B.n450 VSUBS 0.007973f
C624 B.n451 VSUBS 0.007973f
C625 B.n452 VSUBS 0.007973f
C626 B.n453 VSUBS 0.007973f
C627 B.n454 VSUBS 0.007973f
C628 B.n455 VSUBS 0.007973f
C629 B.n456 VSUBS 0.007973f
C630 B.n457 VSUBS 0.007973f
C631 B.n458 VSUBS 0.007973f
C632 B.n459 VSUBS 0.007973f
C633 B.n460 VSUBS 0.007973f
C634 B.n461 VSUBS 0.007973f
C635 B.n462 VSUBS 0.007973f
C636 B.n463 VSUBS 0.007973f
C637 B.n464 VSUBS 0.007973f
C638 B.n465 VSUBS 0.007973f
C639 B.n466 VSUBS 0.007973f
C640 B.n467 VSUBS 0.007973f
C641 B.n468 VSUBS 0.007973f
C642 B.n469 VSUBS 0.007973f
C643 B.n470 VSUBS 0.007973f
C644 B.t8 VSUBS 0.608284f
C645 B.t7 VSUBS 0.638769f
C646 B.t6 VSUBS 3.00239f
C647 B.n471 VSUBS 0.381452f
C648 B.n472 VSUBS 0.086787f
C649 B.n473 VSUBS 0.018473f
C650 B.n474 VSUBS 0.007504f
C651 B.n475 VSUBS 0.007973f
C652 B.n476 VSUBS 0.007973f
C653 B.n477 VSUBS 0.007973f
C654 B.n478 VSUBS 0.007973f
C655 B.n479 VSUBS 0.007973f
C656 B.n480 VSUBS 0.007973f
C657 B.n481 VSUBS 0.007973f
C658 B.n482 VSUBS 0.007973f
C659 B.n483 VSUBS 0.007973f
C660 B.n484 VSUBS 0.007973f
C661 B.n485 VSUBS 0.007973f
C662 B.n486 VSUBS 0.007973f
C663 B.n487 VSUBS 0.007973f
C664 B.n488 VSUBS 0.007973f
C665 B.n489 VSUBS 0.007973f
C666 B.n490 VSUBS 0.004456f
C667 B.n491 VSUBS 0.018473f
C668 B.n492 VSUBS 0.007504f
C669 B.n493 VSUBS 0.007973f
C670 B.n494 VSUBS 0.007973f
C671 B.n495 VSUBS 0.007973f
C672 B.n496 VSUBS 0.007973f
C673 B.n497 VSUBS 0.007973f
C674 B.n498 VSUBS 0.007973f
C675 B.n499 VSUBS 0.007973f
C676 B.n500 VSUBS 0.007973f
C677 B.n501 VSUBS 0.007973f
C678 B.n502 VSUBS 0.007973f
C679 B.n503 VSUBS 0.007973f
C680 B.n504 VSUBS 0.007973f
C681 B.n505 VSUBS 0.007973f
C682 B.n506 VSUBS 0.007973f
C683 B.n507 VSUBS 0.007973f
C684 B.n508 VSUBS 0.007973f
C685 B.n509 VSUBS 0.007973f
C686 B.n510 VSUBS 0.007973f
C687 B.n511 VSUBS 0.007973f
C688 B.n512 VSUBS 0.007973f
C689 B.n513 VSUBS 0.007973f
C690 B.n514 VSUBS 0.007973f
C691 B.n515 VSUBS 0.007973f
C692 B.n516 VSUBS 0.007973f
C693 B.n517 VSUBS 0.007973f
C694 B.n518 VSUBS 0.007973f
C695 B.n519 VSUBS 0.007973f
C696 B.n520 VSUBS 0.007973f
C697 B.n521 VSUBS 0.007973f
C698 B.n522 VSUBS 0.007973f
C699 B.n523 VSUBS 0.007973f
C700 B.n524 VSUBS 0.007973f
C701 B.n525 VSUBS 0.007973f
C702 B.n526 VSUBS 0.007973f
C703 B.n527 VSUBS 0.007973f
C704 B.n528 VSUBS 0.007973f
C705 B.n529 VSUBS 0.007973f
C706 B.n530 VSUBS 0.007973f
C707 B.n531 VSUBS 0.007973f
C708 B.n532 VSUBS 0.007973f
C709 B.n533 VSUBS 0.007973f
C710 B.n534 VSUBS 0.007973f
C711 B.n535 VSUBS 0.007973f
C712 B.n536 VSUBS 0.007973f
C713 B.n537 VSUBS 0.007973f
C714 B.n538 VSUBS 0.007973f
C715 B.n539 VSUBS 0.007973f
C716 B.n540 VSUBS 0.007973f
C717 B.n541 VSUBS 0.007973f
C718 B.n542 VSUBS 0.007973f
C719 B.n543 VSUBS 0.007973f
C720 B.n544 VSUBS 0.007973f
C721 B.n545 VSUBS 0.007973f
C722 B.n546 VSUBS 0.007973f
C723 B.n547 VSUBS 0.007973f
C724 B.n548 VSUBS 0.007973f
C725 B.n549 VSUBS 0.007973f
C726 B.n550 VSUBS 0.007973f
C727 B.n551 VSUBS 0.007973f
C728 B.n552 VSUBS 0.007973f
C729 B.n553 VSUBS 0.007973f
C730 B.n554 VSUBS 0.007973f
C731 B.n555 VSUBS 0.007973f
C732 B.n556 VSUBS 0.007973f
C733 B.n557 VSUBS 0.007973f
C734 B.n558 VSUBS 0.007973f
C735 B.n559 VSUBS 0.007973f
C736 B.n560 VSUBS 0.007973f
C737 B.n561 VSUBS 0.007973f
C738 B.n562 VSUBS 0.007973f
C739 B.n563 VSUBS 0.007973f
C740 B.n564 VSUBS 0.007973f
C741 B.n565 VSUBS 0.007973f
C742 B.n566 VSUBS 0.007973f
C743 B.n567 VSUBS 0.007973f
C744 B.n568 VSUBS 0.007973f
C745 B.n569 VSUBS 0.007973f
C746 B.n570 VSUBS 0.018945f
C747 B.n571 VSUBS 0.01975f
C748 B.n572 VSUBS 0.018858f
C749 B.n573 VSUBS 0.007973f
C750 B.n574 VSUBS 0.007973f
C751 B.n575 VSUBS 0.007973f
C752 B.n576 VSUBS 0.007973f
C753 B.n577 VSUBS 0.007973f
C754 B.n578 VSUBS 0.007973f
C755 B.n579 VSUBS 0.007973f
C756 B.n580 VSUBS 0.007973f
C757 B.n581 VSUBS 0.007973f
C758 B.n582 VSUBS 0.007973f
C759 B.n583 VSUBS 0.007973f
C760 B.n584 VSUBS 0.007973f
C761 B.n585 VSUBS 0.007973f
C762 B.n586 VSUBS 0.007973f
C763 B.n587 VSUBS 0.007973f
C764 B.n588 VSUBS 0.007973f
C765 B.n589 VSUBS 0.007973f
C766 B.n590 VSUBS 0.007973f
C767 B.n591 VSUBS 0.007973f
C768 B.n592 VSUBS 0.007973f
C769 B.n593 VSUBS 0.007973f
C770 B.n594 VSUBS 0.007973f
C771 B.n595 VSUBS 0.007973f
C772 B.n596 VSUBS 0.007973f
C773 B.n597 VSUBS 0.007973f
C774 B.n598 VSUBS 0.007973f
C775 B.n599 VSUBS 0.007973f
C776 B.n600 VSUBS 0.007973f
C777 B.n601 VSUBS 0.007973f
C778 B.n602 VSUBS 0.007973f
C779 B.n603 VSUBS 0.007973f
C780 B.n604 VSUBS 0.007973f
C781 B.n605 VSUBS 0.007973f
C782 B.n606 VSUBS 0.007973f
C783 B.n607 VSUBS 0.007973f
C784 B.n608 VSUBS 0.007973f
C785 B.n609 VSUBS 0.007973f
C786 B.n610 VSUBS 0.007973f
C787 B.n611 VSUBS 0.007973f
C788 B.n612 VSUBS 0.007973f
C789 B.n613 VSUBS 0.007973f
C790 B.n614 VSUBS 0.007973f
C791 B.n615 VSUBS 0.007973f
C792 B.n616 VSUBS 0.007973f
C793 B.n617 VSUBS 0.007973f
C794 B.n618 VSUBS 0.007973f
C795 B.n619 VSUBS 0.007973f
C796 B.n620 VSUBS 0.007973f
C797 B.n621 VSUBS 0.007973f
C798 B.n622 VSUBS 0.007973f
C799 B.n623 VSUBS 0.007973f
C800 B.n624 VSUBS 0.007973f
C801 B.n625 VSUBS 0.007973f
C802 B.n626 VSUBS 0.007973f
C803 B.n627 VSUBS 0.007973f
C804 B.n628 VSUBS 0.007973f
C805 B.n629 VSUBS 0.007973f
C806 B.n630 VSUBS 0.007973f
C807 B.n631 VSUBS 0.007973f
C808 B.n632 VSUBS 0.007973f
C809 B.n633 VSUBS 0.007973f
C810 B.n634 VSUBS 0.007973f
C811 B.n635 VSUBS 0.007973f
C812 B.n636 VSUBS 0.007973f
C813 B.n637 VSUBS 0.007973f
C814 B.n638 VSUBS 0.007973f
C815 B.n639 VSUBS 0.007973f
C816 B.n640 VSUBS 0.007973f
C817 B.n641 VSUBS 0.007973f
C818 B.n642 VSUBS 0.007973f
C819 B.n643 VSUBS 0.007973f
C820 B.n644 VSUBS 0.007973f
C821 B.n645 VSUBS 0.007973f
C822 B.n646 VSUBS 0.007973f
C823 B.n647 VSUBS 0.007973f
C824 B.n648 VSUBS 0.007973f
C825 B.n649 VSUBS 0.007973f
C826 B.n650 VSUBS 0.007973f
C827 B.n651 VSUBS 0.007973f
C828 B.n652 VSUBS 0.007973f
C829 B.n653 VSUBS 0.007973f
C830 B.n654 VSUBS 0.007973f
C831 B.n655 VSUBS 0.007973f
C832 B.n656 VSUBS 0.007973f
C833 B.n657 VSUBS 0.007973f
C834 B.n658 VSUBS 0.007973f
C835 B.n659 VSUBS 0.007973f
C836 B.n660 VSUBS 0.007973f
C837 B.n661 VSUBS 0.007973f
C838 B.n662 VSUBS 0.007973f
C839 B.n663 VSUBS 0.007973f
C840 B.n664 VSUBS 0.007973f
C841 B.n665 VSUBS 0.007973f
C842 B.n666 VSUBS 0.007973f
C843 B.n667 VSUBS 0.007973f
C844 B.n668 VSUBS 0.007973f
C845 B.n669 VSUBS 0.007973f
C846 B.n670 VSUBS 0.007973f
C847 B.n671 VSUBS 0.007973f
C848 B.n672 VSUBS 0.007973f
C849 B.n673 VSUBS 0.007973f
C850 B.n674 VSUBS 0.007973f
C851 B.n675 VSUBS 0.007973f
C852 B.n676 VSUBS 0.007973f
C853 B.n677 VSUBS 0.007973f
C854 B.n678 VSUBS 0.007973f
C855 B.n679 VSUBS 0.007973f
C856 B.n680 VSUBS 0.007973f
C857 B.n681 VSUBS 0.007973f
C858 B.n682 VSUBS 0.007973f
C859 B.n683 VSUBS 0.007973f
C860 B.n684 VSUBS 0.007973f
C861 B.n685 VSUBS 0.007973f
C862 B.n686 VSUBS 0.007973f
C863 B.n687 VSUBS 0.007973f
C864 B.n688 VSUBS 0.007973f
C865 B.n689 VSUBS 0.007973f
C866 B.n690 VSUBS 0.007973f
C867 B.n691 VSUBS 0.007973f
C868 B.n692 VSUBS 0.007973f
C869 B.n693 VSUBS 0.007973f
C870 B.n694 VSUBS 0.007973f
C871 B.n695 VSUBS 0.007973f
C872 B.n696 VSUBS 0.007973f
C873 B.n697 VSUBS 0.007973f
C874 B.n698 VSUBS 0.007973f
C875 B.n699 VSUBS 0.007973f
C876 B.n700 VSUBS 0.007973f
C877 B.n701 VSUBS 0.007973f
C878 B.n702 VSUBS 0.007973f
C879 B.n703 VSUBS 0.007973f
C880 B.n704 VSUBS 0.007973f
C881 B.n705 VSUBS 0.007973f
C882 B.n706 VSUBS 0.007973f
C883 B.n707 VSUBS 0.007973f
C884 B.n708 VSUBS 0.007973f
C885 B.n709 VSUBS 0.007973f
C886 B.n710 VSUBS 0.007973f
C887 B.n711 VSUBS 0.007973f
C888 B.n712 VSUBS 0.007973f
C889 B.n713 VSUBS 0.007973f
C890 B.n714 VSUBS 0.007973f
C891 B.n715 VSUBS 0.007973f
C892 B.n716 VSUBS 0.007973f
C893 B.n717 VSUBS 0.007973f
C894 B.n718 VSUBS 0.007973f
C895 B.n719 VSUBS 0.007973f
C896 B.n720 VSUBS 0.007973f
C897 B.n721 VSUBS 0.007973f
C898 B.n722 VSUBS 0.007973f
C899 B.n723 VSUBS 0.007973f
C900 B.n724 VSUBS 0.007973f
C901 B.n725 VSUBS 0.007973f
C902 B.n726 VSUBS 0.007973f
C903 B.n727 VSUBS 0.007973f
C904 B.n728 VSUBS 0.007973f
C905 B.n729 VSUBS 0.007973f
C906 B.n730 VSUBS 0.007973f
C907 B.n731 VSUBS 0.007973f
C908 B.n732 VSUBS 0.007973f
C909 B.n733 VSUBS 0.007973f
C910 B.n734 VSUBS 0.007973f
C911 B.n735 VSUBS 0.007973f
C912 B.n736 VSUBS 0.007973f
C913 B.n737 VSUBS 0.007973f
C914 B.n738 VSUBS 0.007973f
C915 B.n739 VSUBS 0.007973f
C916 B.n740 VSUBS 0.007973f
C917 B.n741 VSUBS 0.007973f
C918 B.n742 VSUBS 0.007973f
C919 B.n743 VSUBS 0.007973f
C920 B.n744 VSUBS 0.007973f
C921 B.n745 VSUBS 0.007973f
C922 B.n746 VSUBS 0.007973f
C923 B.n747 VSUBS 0.007973f
C924 B.n748 VSUBS 0.007973f
C925 B.n749 VSUBS 0.007973f
C926 B.n750 VSUBS 0.007973f
C927 B.n751 VSUBS 0.007973f
C928 B.n752 VSUBS 0.007973f
C929 B.n753 VSUBS 0.007973f
C930 B.n754 VSUBS 0.007973f
C931 B.n755 VSUBS 0.007973f
C932 B.n756 VSUBS 0.007973f
C933 B.n757 VSUBS 0.007973f
C934 B.n758 VSUBS 0.007973f
C935 B.n759 VSUBS 0.007973f
C936 B.n760 VSUBS 0.007973f
C937 B.n761 VSUBS 0.007973f
C938 B.n762 VSUBS 0.007973f
C939 B.n763 VSUBS 0.007973f
C940 B.n764 VSUBS 0.007973f
C941 B.n765 VSUBS 0.007973f
C942 B.n766 VSUBS 0.007973f
C943 B.n767 VSUBS 0.007973f
C944 B.n768 VSUBS 0.007973f
C945 B.n769 VSUBS 0.007973f
C946 B.n770 VSUBS 0.007973f
C947 B.n771 VSUBS 0.007973f
C948 B.n772 VSUBS 0.007973f
C949 B.n773 VSUBS 0.007973f
C950 B.n774 VSUBS 0.007973f
C951 B.n775 VSUBS 0.007973f
C952 B.n776 VSUBS 0.007973f
C953 B.n777 VSUBS 0.007973f
C954 B.n778 VSUBS 0.007973f
C955 B.n779 VSUBS 0.007973f
C956 B.n780 VSUBS 0.007973f
C957 B.n781 VSUBS 0.007973f
C958 B.n782 VSUBS 0.007973f
C959 B.n783 VSUBS 0.007973f
C960 B.n784 VSUBS 0.007973f
C961 B.n785 VSUBS 0.007973f
C962 B.n786 VSUBS 0.007973f
C963 B.n787 VSUBS 0.007973f
C964 B.n788 VSUBS 0.007973f
C965 B.n789 VSUBS 0.007973f
C966 B.n790 VSUBS 0.007973f
C967 B.n791 VSUBS 0.007973f
C968 B.n792 VSUBS 0.007973f
C969 B.n793 VSUBS 0.007973f
C970 B.n794 VSUBS 0.007973f
C971 B.n795 VSUBS 0.007973f
C972 B.n796 VSUBS 0.007973f
C973 B.n797 VSUBS 0.007973f
C974 B.n798 VSUBS 0.007973f
C975 B.n799 VSUBS 0.007973f
C976 B.n800 VSUBS 0.007973f
C977 B.n801 VSUBS 0.007973f
C978 B.n802 VSUBS 0.007973f
C979 B.n803 VSUBS 0.007973f
C980 B.n804 VSUBS 0.018858f
C981 B.n805 VSUBS 0.019837f
C982 B.n806 VSUBS 0.019837f
C983 B.n807 VSUBS 0.007973f
C984 B.n808 VSUBS 0.007973f
C985 B.n809 VSUBS 0.007973f
C986 B.n810 VSUBS 0.007973f
C987 B.n811 VSUBS 0.007973f
C988 B.n812 VSUBS 0.007973f
C989 B.n813 VSUBS 0.007973f
C990 B.n814 VSUBS 0.007973f
C991 B.n815 VSUBS 0.007973f
C992 B.n816 VSUBS 0.007973f
C993 B.n817 VSUBS 0.007973f
C994 B.n818 VSUBS 0.007973f
C995 B.n819 VSUBS 0.007973f
C996 B.n820 VSUBS 0.007973f
C997 B.n821 VSUBS 0.007973f
C998 B.n822 VSUBS 0.007973f
C999 B.n823 VSUBS 0.007973f
C1000 B.n824 VSUBS 0.007973f
C1001 B.n825 VSUBS 0.007973f
C1002 B.n826 VSUBS 0.007973f
C1003 B.n827 VSUBS 0.007973f
C1004 B.n828 VSUBS 0.007973f
C1005 B.n829 VSUBS 0.007973f
C1006 B.n830 VSUBS 0.007973f
C1007 B.n831 VSUBS 0.007973f
C1008 B.n832 VSUBS 0.007973f
C1009 B.n833 VSUBS 0.007973f
C1010 B.n834 VSUBS 0.007973f
C1011 B.n835 VSUBS 0.007973f
C1012 B.n836 VSUBS 0.007973f
C1013 B.n837 VSUBS 0.007973f
C1014 B.n838 VSUBS 0.007973f
C1015 B.n839 VSUBS 0.007973f
C1016 B.n840 VSUBS 0.007973f
C1017 B.n841 VSUBS 0.007973f
C1018 B.n842 VSUBS 0.007973f
C1019 B.n843 VSUBS 0.007973f
C1020 B.n844 VSUBS 0.007973f
C1021 B.n845 VSUBS 0.007973f
C1022 B.n846 VSUBS 0.007973f
C1023 B.n847 VSUBS 0.007973f
C1024 B.n848 VSUBS 0.007973f
C1025 B.n849 VSUBS 0.007973f
C1026 B.n850 VSUBS 0.007973f
C1027 B.n851 VSUBS 0.007973f
C1028 B.n852 VSUBS 0.007973f
C1029 B.n853 VSUBS 0.007973f
C1030 B.n854 VSUBS 0.007973f
C1031 B.n855 VSUBS 0.007973f
C1032 B.n856 VSUBS 0.007973f
C1033 B.n857 VSUBS 0.007973f
C1034 B.n858 VSUBS 0.007973f
C1035 B.n859 VSUBS 0.007973f
C1036 B.n860 VSUBS 0.007973f
C1037 B.n861 VSUBS 0.007973f
C1038 B.n862 VSUBS 0.007973f
C1039 B.n863 VSUBS 0.007973f
C1040 B.n864 VSUBS 0.007973f
C1041 B.n865 VSUBS 0.007973f
C1042 B.n866 VSUBS 0.007973f
C1043 B.n867 VSUBS 0.007973f
C1044 B.n868 VSUBS 0.007973f
C1045 B.n869 VSUBS 0.007973f
C1046 B.n870 VSUBS 0.007973f
C1047 B.n871 VSUBS 0.007973f
C1048 B.n872 VSUBS 0.007973f
C1049 B.n873 VSUBS 0.007973f
C1050 B.n874 VSUBS 0.007973f
C1051 B.n875 VSUBS 0.007973f
C1052 B.n876 VSUBS 0.007973f
C1053 B.n877 VSUBS 0.007973f
C1054 B.n878 VSUBS 0.007973f
C1055 B.n879 VSUBS 0.007973f
C1056 B.n880 VSUBS 0.007973f
C1057 B.n881 VSUBS 0.007973f
C1058 B.n882 VSUBS 0.007973f
C1059 B.n883 VSUBS 0.007504f
C1060 B.n884 VSUBS 0.007973f
C1061 B.n885 VSUBS 0.007973f
C1062 B.n886 VSUBS 0.004456f
C1063 B.n887 VSUBS 0.007973f
C1064 B.n888 VSUBS 0.007973f
C1065 B.n889 VSUBS 0.007973f
C1066 B.n890 VSUBS 0.007973f
C1067 B.n891 VSUBS 0.007973f
C1068 B.n892 VSUBS 0.007973f
C1069 B.n893 VSUBS 0.007973f
C1070 B.n894 VSUBS 0.007973f
C1071 B.n895 VSUBS 0.007973f
C1072 B.n896 VSUBS 0.007973f
C1073 B.n897 VSUBS 0.007973f
C1074 B.n898 VSUBS 0.007973f
C1075 B.n899 VSUBS 0.004456f
C1076 B.n900 VSUBS 0.018473f
C1077 B.n901 VSUBS 0.007504f
C1078 B.n902 VSUBS 0.007973f
C1079 B.n903 VSUBS 0.007973f
C1080 B.n904 VSUBS 0.007973f
C1081 B.n905 VSUBS 0.007973f
C1082 B.n906 VSUBS 0.007973f
C1083 B.n907 VSUBS 0.007973f
C1084 B.n908 VSUBS 0.007973f
C1085 B.n909 VSUBS 0.007973f
C1086 B.n910 VSUBS 0.007973f
C1087 B.n911 VSUBS 0.007973f
C1088 B.n912 VSUBS 0.007973f
C1089 B.n913 VSUBS 0.007973f
C1090 B.n914 VSUBS 0.007973f
C1091 B.n915 VSUBS 0.007973f
C1092 B.n916 VSUBS 0.007973f
C1093 B.n917 VSUBS 0.007973f
C1094 B.n918 VSUBS 0.007973f
C1095 B.n919 VSUBS 0.007973f
C1096 B.n920 VSUBS 0.007973f
C1097 B.n921 VSUBS 0.007973f
C1098 B.n922 VSUBS 0.007973f
C1099 B.n923 VSUBS 0.007973f
C1100 B.n924 VSUBS 0.007973f
C1101 B.n925 VSUBS 0.007973f
C1102 B.n926 VSUBS 0.007973f
C1103 B.n927 VSUBS 0.007973f
C1104 B.n928 VSUBS 0.007973f
C1105 B.n929 VSUBS 0.007973f
C1106 B.n930 VSUBS 0.007973f
C1107 B.n931 VSUBS 0.007973f
C1108 B.n932 VSUBS 0.007973f
C1109 B.n933 VSUBS 0.007973f
C1110 B.n934 VSUBS 0.007973f
C1111 B.n935 VSUBS 0.007973f
C1112 B.n936 VSUBS 0.007973f
C1113 B.n937 VSUBS 0.007973f
C1114 B.n938 VSUBS 0.007973f
C1115 B.n939 VSUBS 0.007973f
C1116 B.n940 VSUBS 0.007973f
C1117 B.n941 VSUBS 0.007973f
C1118 B.n942 VSUBS 0.007973f
C1119 B.n943 VSUBS 0.007973f
C1120 B.n944 VSUBS 0.007973f
C1121 B.n945 VSUBS 0.007973f
C1122 B.n946 VSUBS 0.007973f
C1123 B.n947 VSUBS 0.007973f
C1124 B.n948 VSUBS 0.007973f
C1125 B.n949 VSUBS 0.007973f
C1126 B.n950 VSUBS 0.007973f
C1127 B.n951 VSUBS 0.007973f
C1128 B.n952 VSUBS 0.007973f
C1129 B.n953 VSUBS 0.007973f
C1130 B.n954 VSUBS 0.007973f
C1131 B.n955 VSUBS 0.007973f
C1132 B.n956 VSUBS 0.007973f
C1133 B.n957 VSUBS 0.007973f
C1134 B.n958 VSUBS 0.007973f
C1135 B.n959 VSUBS 0.007973f
C1136 B.n960 VSUBS 0.007973f
C1137 B.n961 VSUBS 0.007973f
C1138 B.n962 VSUBS 0.007973f
C1139 B.n963 VSUBS 0.007973f
C1140 B.n964 VSUBS 0.007973f
C1141 B.n965 VSUBS 0.007973f
C1142 B.n966 VSUBS 0.007973f
C1143 B.n967 VSUBS 0.007973f
C1144 B.n968 VSUBS 0.007973f
C1145 B.n969 VSUBS 0.007973f
C1146 B.n970 VSUBS 0.007973f
C1147 B.n971 VSUBS 0.007973f
C1148 B.n972 VSUBS 0.007973f
C1149 B.n973 VSUBS 0.007973f
C1150 B.n974 VSUBS 0.007973f
C1151 B.n975 VSUBS 0.007973f
C1152 B.n976 VSUBS 0.007973f
C1153 B.n977 VSUBS 0.007973f
C1154 B.n978 VSUBS 0.007973f
C1155 B.n979 VSUBS 0.019837f
C1156 B.n980 VSUBS 0.019837f
C1157 B.n981 VSUBS 0.018858f
C1158 B.n982 VSUBS 0.007973f
C1159 B.n983 VSUBS 0.007973f
C1160 B.n984 VSUBS 0.007973f
C1161 B.n985 VSUBS 0.007973f
C1162 B.n986 VSUBS 0.007973f
C1163 B.n987 VSUBS 0.007973f
C1164 B.n988 VSUBS 0.007973f
C1165 B.n989 VSUBS 0.007973f
C1166 B.n990 VSUBS 0.007973f
C1167 B.n991 VSUBS 0.007973f
C1168 B.n992 VSUBS 0.007973f
C1169 B.n993 VSUBS 0.007973f
C1170 B.n994 VSUBS 0.007973f
C1171 B.n995 VSUBS 0.007973f
C1172 B.n996 VSUBS 0.007973f
C1173 B.n997 VSUBS 0.007973f
C1174 B.n998 VSUBS 0.007973f
C1175 B.n999 VSUBS 0.007973f
C1176 B.n1000 VSUBS 0.007973f
C1177 B.n1001 VSUBS 0.007973f
C1178 B.n1002 VSUBS 0.007973f
C1179 B.n1003 VSUBS 0.007973f
C1180 B.n1004 VSUBS 0.007973f
C1181 B.n1005 VSUBS 0.007973f
C1182 B.n1006 VSUBS 0.007973f
C1183 B.n1007 VSUBS 0.007973f
C1184 B.n1008 VSUBS 0.007973f
C1185 B.n1009 VSUBS 0.007973f
C1186 B.n1010 VSUBS 0.007973f
C1187 B.n1011 VSUBS 0.007973f
C1188 B.n1012 VSUBS 0.007973f
C1189 B.n1013 VSUBS 0.007973f
C1190 B.n1014 VSUBS 0.007973f
C1191 B.n1015 VSUBS 0.007973f
C1192 B.n1016 VSUBS 0.007973f
C1193 B.n1017 VSUBS 0.007973f
C1194 B.n1018 VSUBS 0.007973f
C1195 B.n1019 VSUBS 0.007973f
C1196 B.n1020 VSUBS 0.007973f
C1197 B.n1021 VSUBS 0.007973f
C1198 B.n1022 VSUBS 0.007973f
C1199 B.n1023 VSUBS 0.007973f
C1200 B.n1024 VSUBS 0.007973f
C1201 B.n1025 VSUBS 0.007973f
C1202 B.n1026 VSUBS 0.007973f
C1203 B.n1027 VSUBS 0.007973f
C1204 B.n1028 VSUBS 0.007973f
C1205 B.n1029 VSUBS 0.007973f
C1206 B.n1030 VSUBS 0.007973f
C1207 B.n1031 VSUBS 0.007973f
C1208 B.n1032 VSUBS 0.007973f
C1209 B.n1033 VSUBS 0.007973f
C1210 B.n1034 VSUBS 0.007973f
C1211 B.n1035 VSUBS 0.007973f
C1212 B.n1036 VSUBS 0.007973f
C1213 B.n1037 VSUBS 0.007973f
C1214 B.n1038 VSUBS 0.007973f
C1215 B.n1039 VSUBS 0.007973f
C1216 B.n1040 VSUBS 0.007973f
C1217 B.n1041 VSUBS 0.007973f
C1218 B.n1042 VSUBS 0.007973f
C1219 B.n1043 VSUBS 0.007973f
C1220 B.n1044 VSUBS 0.007973f
C1221 B.n1045 VSUBS 0.007973f
C1222 B.n1046 VSUBS 0.007973f
C1223 B.n1047 VSUBS 0.007973f
C1224 B.n1048 VSUBS 0.007973f
C1225 B.n1049 VSUBS 0.007973f
C1226 B.n1050 VSUBS 0.007973f
C1227 B.n1051 VSUBS 0.007973f
C1228 B.n1052 VSUBS 0.007973f
C1229 B.n1053 VSUBS 0.007973f
C1230 B.n1054 VSUBS 0.007973f
C1231 B.n1055 VSUBS 0.007973f
C1232 B.n1056 VSUBS 0.007973f
C1233 B.n1057 VSUBS 0.007973f
C1234 B.n1058 VSUBS 0.007973f
C1235 B.n1059 VSUBS 0.007973f
C1236 B.n1060 VSUBS 0.007973f
C1237 B.n1061 VSUBS 0.007973f
C1238 B.n1062 VSUBS 0.007973f
C1239 B.n1063 VSUBS 0.007973f
C1240 B.n1064 VSUBS 0.007973f
C1241 B.n1065 VSUBS 0.007973f
C1242 B.n1066 VSUBS 0.007973f
C1243 B.n1067 VSUBS 0.007973f
C1244 B.n1068 VSUBS 0.007973f
C1245 B.n1069 VSUBS 0.007973f
C1246 B.n1070 VSUBS 0.007973f
C1247 B.n1071 VSUBS 0.007973f
C1248 B.n1072 VSUBS 0.007973f
C1249 B.n1073 VSUBS 0.007973f
C1250 B.n1074 VSUBS 0.007973f
C1251 B.n1075 VSUBS 0.007973f
C1252 B.n1076 VSUBS 0.007973f
C1253 B.n1077 VSUBS 0.007973f
C1254 B.n1078 VSUBS 0.007973f
C1255 B.n1079 VSUBS 0.007973f
C1256 B.n1080 VSUBS 0.007973f
C1257 B.n1081 VSUBS 0.007973f
C1258 B.n1082 VSUBS 0.007973f
C1259 B.n1083 VSUBS 0.007973f
C1260 B.n1084 VSUBS 0.007973f
C1261 B.n1085 VSUBS 0.007973f
C1262 B.n1086 VSUBS 0.007973f
C1263 B.n1087 VSUBS 0.007973f
C1264 B.n1088 VSUBS 0.007973f
C1265 B.n1089 VSUBS 0.007973f
C1266 B.n1090 VSUBS 0.007973f
C1267 B.n1091 VSUBS 0.007973f
C1268 B.n1092 VSUBS 0.007973f
C1269 B.n1093 VSUBS 0.007973f
C1270 B.n1094 VSUBS 0.007973f
C1271 B.n1095 VSUBS 0.010405f
C1272 B.n1096 VSUBS 0.011084f
C1273 B.n1097 VSUBS 0.022041f
C1274 VTAIL.t0 VSUBS 0.359f
C1275 VTAIL.t3 VSUBS 0.359f
C1276 VTAIL.n0 VSUBS 2.72858f
C1277 VTAIL.n1 VSUBS 1.15894f
C1278 VTAIL.t14 VSUBS 3.57979f
C1279 VTAIL.n2 VSUBS 1.35937f
C1280 VTAIL.t10 VSUBS 0.359f
C1281 VTAIL.t12 VSUBS 0.359f
C1282 VTAIL.n3 VSUBS 2.72858f
C1283 VTAIL.n4 VSUBS 1.34416f
C1284 VTAIL.t15 VSUBS 0.359f
C1285 VTAIL.t9 VSUBS 0.359f
C1286 VTAIL.n5 VSUBS 2.72858f
C1287 VTAIL.n6 VSUBS 3.30429f
C1288 VTAIL.t18 VSUBS 0.359f
C1289 VTAIL.t6 VSUBS 0.359f
C1290 VTAIL.n7 VSUBS 2.7286f
C1291 VTAIL.n8 VSUBS 3.30427f
C1292 VTAIL.t4 VSUBS 0.359f
C1293 VTAIL.t7 VSUBS 0.359f
C1294 VTAIL.n9 VSUBS 2.7286f
C1295 VTAIL.n10 VSUBS 1.34414f
C1296 VTAIL.t1 VSUBS 3.5798f
C1297 VTAIL.n11 VSUBS 1.35935f
C1298 VTAIL.t16 VSUBS 0.359f
C1299 VTAIL.t11 VSUBS 0.359f
C1300 VTAIL.n12 VSUBS 2.7286f
C1301 VTAIL.n13 VSUBS 1.23147f
C1302 VTAIL.t8 VSUBS 0.359f
C1303 VTAIL.t17 VSUBS 0.359f
C1304 VTAIL.n14 VSUBS 2.7286f
C1305 VTAIL.n15 VSUBS 1.34414f
C1306 VTAIL.t13 VSUBS 3.57981f
C1307 VTAIL.n16 VSUBS 3.12062f
C1308 VTAIL.t19 VSUBS 3.57979f
C1309 VTAIL.n17 VSUBS 3.12064f
C1310 VTAIL.t2 VSUBS 0.359f
C1311 VTAIL.t5 VSUBS 0.359f
C1312 VTAIL.n18 VSUBS 2.72858f
C1313 VTAIL.n19 VSUBS 1.10517f
C1314 VDD1.t4 VSUBS 3.98012f
C1315 VDD1.t7 VSUBS 0.372461f
C1316 VDD1.t8 VSUBS 0.372461f
C1317 VDD1.n0 VSUBS 3.02294f
C1318 VDD1.n1 VSUBS 1.99573f
C1319 VDD1.t3 VSUBS 3.98011f
C1320 VDD1.t9 VSUBS 0.372461f
C1321 VDD1.t6 VSUBS 0.372461f
C1322 VDD1.n2 VSUBS 3.02294f
C1323 VDD1.n3 VSUBS 1.9858f
C1324 VDD1.t0 VSUBS 0.372461f
C1325 VDD1.t2 VSUBS 0.372461f
C1326 VDD1.n4 VSUBS 3.06427f
C1327 VDD1.n5 VSUBS 4.87344f
C1328 VDD1.t5 VSUBS 0.372461f
C1329 VDD1.t1 VSUBS 0.372461f
C1330 VDD1.n6 VSUBS 3.02294f
C1331 VDD1.n7 VSUBS 4.94881f
C1332 VP.t3 VSUBS 3.68925f
C1333 VP.n0 VSUBS 1.36449f
C1334 VP.n1 VSUBS 0.023336f
C1335 VP.n2 VSUBS 0.039676f
C1336 VP.n3 VSUBS 0.023336f
C1337 VP.n4 VSUBS 0.035156f
C1338 VP.n5 VSUBS 0.023336f
C1339 VP.n6 VSUBS 0.035859f
C1340 VP.n7 VSUBS 0.023336f
C1341 VP.n8 VSUBS 0.032593f
C1342 VP.n9 VSUBS 0.023336f
C1343 VP.n10 VSUBS 0.031985f
C1344 VP.n11 VSUBS 0.023336f
C1345 VP.n12 VSUBS 0.030029f
C1346 VP.n13 VSUBS 0.023336f
C1347 VP.n14 VSUBS 0.027764f
C1348 VP.n15 VSUBS 0.023336f
C1349 VP.n16 VSUBS 0.027465f
C1350 VP.t4 VSUBS 3.68925f
C1351 VP.n17 VSUBS 1.36449f
C1352 VP.n18 VSUBS 0.023336f
C1353 VP.n19 VSUBS 0.039676f
C1354 VP.n20 VSUBS 0.023336f
C1355 VP.n21 VSUBS 0.035156f
C1356 VP.n22 VSUBS 0.023336f
C1357 VP.n23 VSUBS 0.035859f
C1358 VP.n24 VSUBS 0.023336f
C1359 VP.n25 VSUBS 0.032593f
C1360 VP.n26 VSUBS 0.023336f
C1361 VP.n27 VSUBS 0.031985f
C1362 VP.n28 VSUBS 0.023336f
C1363 VP.n29 VSUBS 0.030029f
C1364 VP.t1 VSUBS 4.03128f
C1365 VP.t6 VSUBS 3.68925f
C1366 VP.n30 VSUBS 1.35543f
C1367 VP.n31 VSUBS 1.29365f
C1368 VP.n32 VSUBS 0.292579f
C1369 VP.n33 VSUBS 0.023336f
C1370 VP.n34 VSUBS 0.043274f
C1371 VP.n35 VSUBS 0.043274f
C1372 VP.n36 VSUBS 0.035859f
C1373 VP.n37 VSUBS 0.023336f
C1374 VP.n38 VSUBS 0.023336f
C1375 VP.n39 VSUBS 0.023336f
C1376 VP.n40 VSUBS 0.043274f
C1377 VP.n41 VSUBS 0.043274f
C1378 VP.t9 VSUBS 3.68925f
C1379 VP.n42 VSUBS 1.27735f
C1380 VP.n43 VSUBS 0.032593f
C1381 VP.n44 VSUBS 0.023336f
C1382 VP.n45 VSUBS 0.023336f
C1383 VP.n46 VSUBS 0.023336f
C1384 VP.n47 VSUBS 0.043274f
C1385 VP.n48 VSUBS 0.043274f
C1386 VP.n49 VSUBS 0.031985f
C1387 VP.n50 VSUBS 0.023336f
C1388 VP.n51 VSUBS 0.023336f
C1389 VP.n52 VSUBS 0.023336f
C1390 VP.n53 VSUBS 0.043274f
C1391 VP.n54 VSUBS 0.043274f
C1392 VP.t0 VSUBS 3.68925f
C1393 VP.n55 VSUBS 1.27735f
C1394 VP.n56 VSUBS 0.030029f
C1395 VP.n57 VSUBS 0.023336f
C1396 VP.n58 VSUBS 0.023336f
C1397 VP.n59 VSUBS 0.023336f
C1398 VP.n60 VSUBS 0.043274f
C1399 VP.n61 VSUBS 0.043679f
C1400 VP.n62 VSUBS 0.027764f
C1401 VP.n63 VSUBS 0.023336f
C1402 VP.n64 VSUBS 0.023336f
C1403 VP.n65 VSUBS 0.023336f
C1404 VP.n66 VSUBS 0.043274f
C1405 VP.n67 VSUBS 0.043274f
C1406 VP.n68 VSUBS 0.027465f
C1407 VP.n69 VSUBS 0.037658f
C1408 VP.n70 VSUBS 1.7823f
C1409 VP.t2 VSUBS 3.68925f
C1410 VP.n71 VSUBS 1.36449f
C1411 VP.n72 VSUBS 1.79594f
C1412 VP.n73 VSUBS 0.037658f
C1413 VP.n74 VSUBS 0.023336f
C1414 VP.n75 VSUBS 0.043274f
C1415 VP.n76 VSUBS 0.043274f
C1416 VP.n77 VSUBS 0.039676f
C1417 VP.n78 VSUBS 0.023336f
C1418 VP.n79 VSUBS 0.023336f
C1419 VP.n80 VSUBS 0.023336f
C1420 VP.n81 VSUBS 0.043679f
C1421 VP.n82 VSUBS 0.043274f
C1422 VP.t8 VSUBS 3.68925f
C1423 VP.n83 VSUBS 1.27735f
C1424 VP.n84 VSUBS 0.035156f
C1425 VP.n85 VSUBS 0.023336f
C1426 VP.n86 VSUBS 0.023336f
C1427 VP.n87 VSUBS 0.023336f
C1428 VP.n88 VSUBS 0.043274f
C1429 VP.n89 VSUBS 0.043274f
C1430 VP.n90 VSUBS 0.035859f
C1431 VP.n91 VSUBS 0.023336f
C1432 VP.n92 VSUBS 0.023336f
C1433 VP.n93 VSUBS 0.023336f
C1434 VP.n94 VSUBS 0.043274f
C1435 VP.n95 VSUBS 0.043274f
C1436 VP.t7 VSUBS 3.68925f
C1437 VP.n96 VSUBS 1.27735f
C1438 VP.n97 VSUBS 0.032593f
C1439 VP.n98 VSUBS 0.023336f
C1440 VP.n99 VSUBS 0.023336f
C1441 VP.n100 VSUBS 0.023336f
C1442 VP.n101 VSUBS 0.043274f
C1443 VP.n102 VSUBS 0.043274f
C1444 VP.n103 VSUBS 0.031985f
C1445 VP.n104 VSUBS 0.023336f
C1446 VP.n105 VSUBS 0.023336f
C1447 VP.n106 VSUBS 0.023336f
C1448 VP.n107 VSUBS 0.043274f
C1449 VP.n108 VSUBS 0.043274f
C1450 VP.t5 VSUBS 3.68925f
C1451 VP.n109 VSUBS 1.27735f
C1452 VP.n110 VSUBS 0.030029f
C1453 VP.n111 VSUBS 0.023336f
C1454 VP.n112 VSUBS 0.023336f
C1455 VP.n113 VSUBS 0.023336f
C1456 VP.n114 VSUBS 0.043274f
C1457 VP.n115 VSUBS 0.043679f
C1458 VP.n116 VSUBS 0.027764f
C1459 VP.n117 VSUBS 0.023336f
C1460 VP.n118 VSUBS 0.023336f
C1461 VP.n119 VSUBS 0.023336f
C1462 VP.n120 VSUBS 0.043274f
C1463 VP.n121 VSUBS 0.043274f
C1464 VP.n122 VSUBS 0.027465f
C1465 VP.n123 VSUBS 0.037658f
C1466 VP.n124 VSUBS 0.066726f
.ends

