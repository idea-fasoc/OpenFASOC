* NGSPICE file created from diff_pair_sample_0191.ext - technology: sky130A

.subckt diff_pair_sample_0191 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.1122 pd=1.01 as=0.2652 ps=2.14 w=0.68 l=3.42
X1 VTAIL.t1 VN.t0 VDD2.t3 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0.1122 ps=1.01 w=0.68 l=3.42
X2 B.t11 B.t9 B.t10 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0 ps=0 w=0.68 l=3.42
X3 B.t8 B.t6 B.t7 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0 ps=0 w=0.68 l=3.42
X4 VDD2.t2 VN.t1 VTAIL.t0 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.1122 pd=1.01 as=0.2652 ps=2.14 w=0.68 l=3.42
X5 VTAIL.t7 VP.t1 VDD1.t2 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0.1122 ps=1.01 w=0.68 l=3.42
X6 B.t5 B.t3 B.t4 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0 ps=0 w=0.68 l=3.42
X7 B.t2 B.t0 B.t1 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0 ps=0 w=0.68 l=3.42
X8 VTAIL.t6 VP.t2 VDD1.t1 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0.1122 ps=1.01 w=0.68 l=3.42
X9 VDD2.t1 VN.t2 VTAIL.t2 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.1122 pd=1.01 as=0.2652 ps=2.14 w=0.68 l=3.42
X10 VDD1.t0 VP.t3 VTAIL.t4 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.1122 pd=1.01 as=0.2652 ps=2.14 w=0.68 l=3.42
X11 VTAIL.t3 VN.t3 VDD2.t0 w_n3220_n1104# sky130_fd_pr__pfet_01v8 ad=0.2652 pd=2.14 as=0.1122 ps=1.01 w=0.68 l=3.42
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n7 VP.n6 83.8051
R9 VP.n20 VP.n0 83.8051
R10 VP.n12 VP.n2 56.4773
R11 VP.n7 VP.n5 42.5093
R12 VP.n5 VP.t1 38.7459
R13 VP.n5 VP.t0 37.5466
R14 VP.n10 VP.n4 24.3439
R15 VP.n11 VP.n10 24.3439
R16 VP.n12 VP.n11 24.3439
R17 VP.n16 VP.n2 24.3439
R18 VP.n17 VP.n16 24.3439
R19 VP.n18 VP.n17 24.3439
R20 VP.n6 VP.n4 6.08636
R21 VP.n18 VP.n0 6.08636
R22 VP.n6 VP.t2 4.79231
R23 VP.n0 VP.t3 4.79231
R24 VP.n8 VP.n7 0.355081
R25 VP.n20 VP.n19 0.355081
R26 VP VP.n20 0.26685
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VTAIL.n7 VTAIL.t2 666.538
R35 VTAIL.n0 VTAIL.t3 666.538
R36 VTAIL.n1 VTAIL.t4 666.538
R37 VTAIL.n2 VTAIL.t6 666.538
R38 VTAIL.n6 VTAIL.t5 666.538
R39 VTAIL.n5 VTAIL.t7 666.538
R40 VTAIL.n4 VTAIL.t0 666.538
R41 VTAIL.n3 VTAIL.t1 666.538
R42 VTAIL.n7 VTAIL.n6 16.1858
R43 VTAIL.n3 VTAIL.n2 16.1858
R44 VTAIL.n4 VTAIL.n3 3.23326
R45 VTAIL.n6 VTAIL.n5 3.23326
R46 VTAIL.n2 VTAIL.n1 3.23326
R47 VTAIL VTAIL.n0 1.67507
R48 VTAIL VTAIL.n7 1.55869
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 VDD1 VDD1.n1 669.939
R52 VDD1 VDD1.n0 635.473
R53 VDD1.n0 VDD1.t2 47.802
R54 VDD1.n0 VDD1.t3 47.802
R55 VDD1.n1 VDD1.t1 47.802
R56 VDD1.n1 VDD1.t0 47.802
R57 VN VN.n1 42.6748
R58 VN.n1 VN.t1 38.7461
R59 VN.n0 VN.t3 38.7461
R60 VN.n0 VN.t2 37.5466
R61 VN.n1 VN.t0 37.5466
R62 VN VN.n0 2.2922
R63 VDD2.n2 VDD2.n0 669.414
R64 VDD2.n2 VDD2.n1 635.415
R65 VDD2.n1 VDD2.t3 47.802
R66 VDD2.n1 VDD2.t2 47.802
R67 VDD2.n0 VDD2.t0 47.802
R68 VDD2.n0 VDD2.t1 47.802
R69 VDD2 VDD2.n2 0.0586897
R70 B.n87 B.t2 728.607
R71 B.n93 B.t5 728.607
R72 B.n28 B.t7 728.607
R73 B.n35 B.t10 728.607
R74 B.n88 B.t1 655.88
R75 B.n94 B.t4 655.88
R76 B.n29 B.t8 655.88
R77 B.n36 B.t11 655.88
R78 B.n345 B.n40 585
R79 B.n347 B.n346 585
R80 B.n348 B.n39 585
R81 B.n350 B.n349 585
R82 B.n351 B.n38 585
R83 B.n353 B.n352 585
R84 B.n354 B.n37 585
R85 B.n356 B.n355 585
R86 B.n358 B.n34 585
R87 B.n360 B.n359 585
R88 B.n361 B.n33 585
R89 B.n363 B.n362 585
R90 B.n364 B.n32 585
R91 B.n366 B.n365 585
R92 B.n367 B.n31 585
R93 B.n369 B.n368 585
R94 B.n370 B.n27 585
R95 B.n372 B.n371 585
R96 B.n373 B.n26 585
R97 B.n375 B.n374 585
R98 B.n376 B.n25 585
R99 B.n378 B.n377 585
R100 B.n379 B.n24 585
R101 B.n381 B.n380 585
R102 B.n382 B.n23 585
R103 B.n384 B.n383 585
R104 B.n344 B.n343 585
R105 B.n342 B.n41 585
R106 B.n341 B.n340 585
R107 B.n339 B.n42 585
R108 B.n338 B.n337 585
R109 B.n336 B.n43 585
R110 B.n335 B.n334 585
R111 B.n333 B.n44 585
R112 B.n332 B.n331 585
R113 B.n330 B.n45 585
R114 B.n329 B.n328 585
R115 B.n327 B.n46 585
R116 B.n326 B.n325 585
R117 B.n324 B.n47 585
R118 B.n323 B.n322 585
R119 B.n321 B.n48 585
R120 B.n320 B.n319 585
R121 B.n318 B.n49 585
R122 B.n317 B.n316 585
R123 B.n315 B.n50 585
R124 B.n314 B.n313 585
R125 B.n312 B.n51 585
R126 B.n311 B.n310 585
R127 B.n309 B.n52 585
R128 B.n308 B.n307 585
R129 B.n306 B.n53 585
R130 B.n305 B.n304 585
R131 B.n303 B.n54 585
R132 B.n302 B.n301 585
R133 B.n300 B.n55 585
R134 B.n299 B.n298 585
R135 B.n297 B.n56 585
R136 B.n296 B.n295 585
R137 B.n294 B.n57 585
R138 B.n293 B.n292 585
R139 B.n291 B.n58 585
R140 B.n290 B.n289 585
R141 B.n288 B.n59 585
R142 B.n287 B.n286 585
R143 B.n285 B.n60 585
R144 B.n284 B.n283 585
R145 B.n282 B.n61 585
R146 B.n281 B.n280 585
R147 B.n279 B.n62 585
R148 B.n278 B.n277 585
R149 B.n276 B.n63 585
R150 B.n275 B.n274 585
R151 B.n273 B.n64 585
R152 B.n272 B.n271 585
R153 B.n270 B.n65 585
R154 B.n269 B.n268 585
R155 B.n267 B.n66 585
R156 B.n266 B.n265 585
R157 B.n264 B.n67 585
R158 B.n263 B.n262 585
R159 B.n261 B.n68 585
R160 B.n260 B.n259 585
R161 B.n258 B.n69 585
R162 B.n257 B.n256 585
R163 B.n255 B.n70 585
R164 B.n254 B.n253 585
R165 B.n252 B.n71 585
R166 B.n251 B.n250 585
R167 B.n249 B.n72 585
R168 B.n248 B.n247 585
R169 B.n246 B.n73 585
R170 B.n245 B.n244 585
R171 B.n243 B.n74 585
R172 B.n242 B.n241 585
R173 B.n240 B.n75 585
R174 B.n239 B.n238 585
R175 B.n237 B.n76 585
R176 B.n236 B.n235 585
R177 B.n234 B.n77 585
R178 B.n233 B.n232 585
R179 B.n231 B.n78 585
R180 B.n230 B.n229 585
R181 B.n228 B.n79 585
R182 B.n227 B.n226 585
R183 B.n225 B.n80 585
R184 B.n224 B.n223 585
R185 B.n222 B.n81 585
R186 B.n221 B.n220 585
R187 B.n180 B.n99 585
R188 B.n182 B.n181 585
R189 B.n183 B.n98 585
R190 B.n185 B.n184 585
R191 B.n186 B.n97 585
R192 B.n188 B.n187 585
R193 B.n189 B.n96 585
R194 B.n191 B.n190 585
R195 B.n193 B.n192 585
R196 B.n194 B.n92 585
R197 B.n196 B.n195 585
R198 B.n197 B.n91 585
R199 B.n199 B.n198 585
R200 B.n200 B.n90 585
R201 B.n202 B.n201 585
R202 B.n203 B.n89 585
R203 B.n205 B.n204 585
R204 B.n206 B.n86 585
R205 B.n209 B.n208 585
R206 B.n210 B.n85 585
R207 B.n212 B.n211 585
R208 B.n213 B.n84 585
R209 B.n215 B.n214 585
R210 B.n216 B.n83 585
R211 B.n218 B.n217 585
R212 B.n219 B.n82 585
R213 B.n179 B.n178 585
R214 B.n177 B.n100 585
R215 B.n176 B.n175 585
R216 B.n174 B.n101 585
R217 B.n173 B.n172 585
R218 B.n171 B.n102 585
R219 B.n170 B.n169 585
R220 B.n168 B.n103 585
R221 B.n167 B.n166 585
R222 B.n165 B.n104 585
R223 B.n164 B.n163 585
R224 B.n162 B.n105 585
R225 B.n161 B.n160 585
R226 B.n159 B.n106 585
R227 B.n158 B.n157 585
R228 B.n156 B.n107 585
R229 B.n155 B.n154 585
R230 B.n153 B.n108 585
R231 B.n152 B.n151 585
R232 B.n150 B.n109 585
R233 B.n149 B.n148 585
R234 B.n147 B.n110 585
R235 B.n146 B.n145 585
R236 B.n144 B.n111 585
R237 B.n143 B.n142 585
R238 B.n141 B.n112 585
R239 B.n140 B.n139 585
R240 B.n138 B.n113 585
R241 B.n137 B.n136 585
R242 B.n135 B.n114 585
R243 B.n134 B.n133 585
R244 B.n132 B.n115 585
R245 B.n131 B.n130 585
R246 B.n129 B.n116 585
R247 B.n128 B.n127 585
R248 B.n126 B.n117 585
R249 B.n125 B.n124 585
R250 B.n123 B.n118 585
R251 B.n122 B.n121 585
R252 B.n120 B.n119 585
R253 B.n2 B.n0 585
R254 B.n445 B.n1 585
R255 B.n444 B.n443 585
R256 B.n442 B.n3 585
R257 B.n441 B.n440 585
R258 B.n439 B.n4 585
R259 B.n438 B.n437 585
R260 B.n436 B.n5 585
R261 B.n435 B.n434 585
R262 B.n433 B.n6 585
R263 B.n432 B.n431 585
R264 B.n430 B.n7 585
R265 B.n429 B.n428 585
R266 B.n427 B.n8 585
R267 B.n426 B.n425 585
R268 B.n424 B.n9 585
R269 B.n423 B.n422 585
R270 B.n421 B.n10 585
R271 B.n420 B.n419 585
R272 B.n418 B.n11 585
R273 B.n417 B.n416 585
R274 B.n415 B.n12 585
R275 B.n414 B.n413 585
R276 B.n412 B.n13 585
R277 B.n411 B.n410 585
R278 B.n409 B.n14 585
R279 B.n408 B.n407 585
R280 B.n406 B.n15 585
R281 B.n405 B.n404 585
R282 B.n403 B.n16 585
R283 B.n402 B.n401 585
R284 B.n400 B.n17 585
R285 B.n399 B.n398 585
R286 B.n397 B.n18 585
R287 B.n396 B.n395 585
R288 B.n394 B.n19 585
R289 B.n393 B.n392 585
R290 B.n391 B.n20 585
R291 B.n390 B.n389 585
R292 B.n388 B.n21 585
R293 B.n387 B.n386 585
R294 B.n385 B.n22 585
R295 B.n447 B.n446 585
R296 B.n180 B.n179 550.159
R297 B.n385 B.n384 550.159
R298 B.n221 B.n82 550.159
R299 B.n343 B.n40 550.159
R300 B.n87 B.t0 210.668
R301 B.n35 B.t9 210.668
R302 B.n93 B.t3 210.466
R303 B.n28 B.t6 210.466
R304 B.n179 B.n100 163.367
R305 B.n175 B.n100 163.367
R306 B.n175 B.n174 163.367
R307 B.n174 B.n173 163.367
R308 B.n173 B.n102 163.367
R309 B.n169 B.n102 163.367
R310 B.n169 B.n168 163.367
R311 B.n168 B.n167 163.367
R312 B.n167 B.n104 163.367
R313 B.n163 B.n104 163.367
R314 B.n163 B.n162 163.367
R315 B.n162 B.n161 163.367
R316 B.n161 B.n106 163.367
R317 B.n157 B.n106 163.367
R318 B.n157 B.n156 163.367
R319 B.n156 B.n155 163.367
R320 B.n155 B.n108 163.367
R321 B.n151 B.n108 163.367
R322 B.n151 B.n150 163.367
R323 B.n150 B.n149 163.367
R324 B.n149 B.n110 163.367
R325 B.n145 B.n110 163.367
R326 B.n145 B.n144 163.367
R327 B.n144 B.n143 163.367
R328 B.n143 B.n112 163.367
R329 B.n139 B.n112 163.367
R330 B.n139 B.n138 163.367
R331 B.n138 B.n137 163.367
R332 B.n137 B.n114 163.367
R333 B.n133 B.n114 163.367
R334 B.n133 B.n132 163.367
R335 B.n132 B.n131 163.367
R336 B.n131 B.n116 163.367
R337 B.n127 B.n116 163.367
R338 B.n127 B.n126 163.367
R339 B.n126 B.n125 163.367
R340 B.n125 B.n118 163.367
R341 B.n121 B.n118 163.367
R342 B.n121 B.n120 163.367
R343 B.n120 B.n2 163.367
R344 B.n446 B.n2 163.367
R345 B.n446 B.n445 163.367
R346 B.n445 B.n444 163.367
R347 B.n444 B.n3 163.367
R348 B.n440 B.n3 163.367
R349 B.n440 B.n439 163.367
R350 B.n439 B.n438 163.367
R351 B.n438 B.n5 163.367
R352 B.n434 B.n5 163.367
R353 B.n434 B.n433 163.367
R354 B.n433 B.n432 163.367
R355 B.n432 B.n7 163.367
R356 B.n428 B.n7 163.367
R357 B.n428 B.n427 163.367
R358 B.n427 B.n426 163.367
R359 B.n426 B.n9 163.367
R360 B.n422 B.n9 163.367
R361 B.n422 B.n421 163.367
R362 B.n421 B.n420 163.367
R363 B.n420 B.n11 163.367
R364 B.n416 B.n11 163.367
R365 B.n416 B.n415 163.367
R366 B.n415 B.n414 163.367
R367 B.n414 B.n13 163.367
R368 B.n410 B.n13 163.367
R369 B.n410 B.n409 163.367
R370 B.n409 B.n408 163.367
R371 B.n408 B.n15 163.367
R372 B.n404 B.n15 163.367
R373 B.n404 B.n403 163.367
R374 B.n403 B.n402 163.367
R375 B.n402 B.n17 163.367
R376 B.n398 B.n17 163.367
R377 B.n398 B.n397 163.367
R378 B.n397 B.n396 163.367
R379 B.n396 B.n19 163.367
R380 B.n392 B.n19 163.367
R381 B.n392 B.n391 163.367
R382 B.n391 B.n390 163.367
R383 B.n390 B.n21 163.367
R384 B.n386 B.n21 163.367
R385 B.n386 B.n385 163.367
R386 B.n181 B.n180 163.367
R387 B.n181 B.n98 163.367
R388 B.n185 B.n98 163.367
R389 B.n186 B.n185 163.367
R390 B.n187 B.n186 163.367
R391 B.n187 B.n96 163.367
R392 B.n191 B.n96 163.367
R393 B.n192 B.n191 163.367
R394 B.n192 B.n92 163.367
R395 B.n196 B.n92 163.367
R396 B.n197 B.n196 163.367
R397 B.n198 B.n197 163.367
R398 B.n198 B.n90 163.367
R399 B.n202 B.n90 163.367
R400 B.n203 B.n202 163.367
R401 B.n204 B.n203 163.367
R402 B.n204 B.n86 163.367
R403 B.n209 B.n86 163.367
R404 B.n210 B.n209 163.367
R405 B.n211 B.n210 163.367
R406 B.n211 B.n84 163.367
R407 B.n215 B.n84 163.367
R408 B.n216 B.n215 163.367
R409 B.n217 B.n216 163.367
R410 B.n217 B.n82 163.367
R411 B.n222 B.n221 163.367
R412 B.n223 B.n222 163.367
R413 B.n223 B.n80 163.367
R414 B.n227 B.n80 163.367
R415 B.n228 B.n227 163.367
R416 B.n229 B.n228 163.367
R417 B.n229 B.n78 163.367
R418 B.n233 B.n78 163.367
R419 B.n234 B.n233 163.367
R420 B.n235 B.n234 163.367
R421 B.n235 B.n76 163.367
R422 B.n239 B.n76 163.367
R423 B.n240 B.n239 163.367
R424 B.n241 B.n240 163.367
R425 B.n241 B.n74 163.367
R426 B.n245 B.n74 163.367
R427 B.n246 B.n245 163.367
R428 B.n247 B.n246 163.367
R429 B.n247 B.n72 163.367
R430 B.n251 B.n72 163.367
R431 B.n252 B.n251 163.367
R432 B.n253 B.n252 163.367
R433 B.n253 B.n70 163.367
R434 B.n257 B.n70 163.367
R435 B.n258 B.n257 163.367
R436 B.n259 B.n258 163.367
R437 B.n259 B.n68 163.367
R438 B.n263 B.n68 163.367
R439 B.n264 B.n263 163.367
R440 B.n265 B.n264 163.367
R441 B.n265 B.n66 163.367
R442 B.n269 B.n66 163.367
R443 B.n270 B.n269 163.367
R444 B.n271 B.n270 163.367
R445 B.n271 B.n64 163.367
R446 B.n275 B.n64 163.367
R447 B.n276 B.n275 163.367
R448 B.n277 B.n276 163.367
R449 B.n277 B.n62 163.367
R450 B.n281 B.n62 163.367
R451 B.n282 B.n281 163.367
R452 B.n283 B.n282 163.367
R453 B.n283 B.n60 163.367
R454 B.n287 B.n60 163.367
R455 B.n288 B.n287 163.367
R456 B.n289 B.n288 163.367
R457 B.n289 B.n58 163.367
R458 B.n293 B.n58 163.367
R459 B.n294 B.n293 163.367
R460 B.n295 B.n294 163.367
R461 B.n295 B.n56 163.367
R462 B.n299 B.n56 163.367
R463 B.n300 B.n299 163.367
R464 B.n301 B.n300 163.367
R465 B.n301 B.n54 163.367
R466 B.n305 B.n54 163.367
R467 B.n306 B.n305 163.367
R468 B.n307 B.n306 163.367
R469 B.n307 B.n52 163.367
R470 B.n311 B.n52 163.367
R471 B.n312 B.n311 163.367
R472 B.n313 B.n312 163.367
R473 B.n313 B.n50 163.367
R474 B.n317 B.n50 163.367
R475 B.n318 B.n317 163.367
R476 B.n319 B.n318 163.367
R477 B.n319 B.n48 163.367
R478 B.n323 B.n48 163.367
R479 B.n324 B.n323 163.367
R480 B.n325 B.n324 163.367
R481 B.n325 B.n46 163.367
R482 B.n329 B.n46 163.367
R483 B.n330 B.n329 163.367
R484 B.n331 B.n330 163.367
R485 B.n331 B.n44 163.367
R486 B.n335 B.n44 163.367
R487 B.n336 B.n335 163.367
R488 B.n337 B.n336 163.367
R489 B.n337 B.n42 163.367
R490 B.n341 B.n42 163.367
R491 B.n342 B.n341 163.367
R492 B.n343 B.n342 163.367
R493 B.n384 B.n23 163.367
R494 B.n380 B.n23 163.367
R495 B.n380 B.n379 163.367
R496 B.n379 B.n378 163.367
R497 B.n378 B.n25 163.367
R498 B.n374 B.n25 163.367
R499 B.n374 B.n373 163.367
R500 B.n373 B.n372 163.367
R501 B.n372 B.n27 163.367
R502 B.n368 B.n27 163.367
R503 B.n368 B.n367 163.367
R504 B.n367 B.n366 163.367
R505 B.n366 B.n32 163.367
R506 B.n362 B.n32 163.367
R507 B.n362 B.n361 163.367
R508 B.n361 B.n360 163.367
R509 B.n360 B.n34 163.367
R510 B.n355 B.n34 163.367
R511 B.n355 B.n354 163.367
R512 B.n354 B.n353 163.367
R513 B.n353 B.n38 163.367
R514 B.n349 B.n38 163.367
R515 B.n349 B.n348 163.367
R516 B.n348 B.n347 163.367
R517 B.n347 B.n40 163.367
R518 B.n88 B.n87 72.7278
R519 B.n94 B.n93 72.7278
R520 B.n29 B.n28 72.7278
R521 B.n36 B.n35 72.7278
R522 B.n207 B.n88 59.5399
R523 B.n95 B.n94 59.5399
R524 B.n30 B.n29 59.5399
R525 B.n357 B.n36 59.5399
R526 B.n345 B.n344 35.7468
R527 B.n383 B.n22 35.7468
R528 B.n220 B.n219 35.7468
R529 B.n178 B.n99 35.7468
R530 B B.n447 18.0485
R531 B.n383 B.n382 10.6151
R532 B.n382 B.n381 10.6151
R533 B.n381 B.n24 10.6151
R534 B.n377 B.n24 10.6151
R535 B.n377 B.n376 10.6151
R536 B.n376 B.n375 10.6151
R537 B.n375 B.n26 10.6151
R538 B.n371 B.n370 10.6151
R539 B.n370 B.n369 10.6151
R540 B.n369 B.n31 10.6151
R541 B.n365 B.n31 10.6151
R542 B.n365 B.n364 10.6151
R543 B.n364 B.n363 10.6151
R544 B.n363 B.n33 10.6151
R545 B.n359 B.n33 10.6151
R546 B.n359 B.n358 10.6151
R547 B.n356 B.n37 10.6151
R548 B.n352 B.n37 10.6151
R549 B.n352 B.n351 10.6151
R550 B.n351 B.n350 10.6151
R551 B.n350 B.n39 10.6151
R552 B.n346 B.n39 10.6151
R553 B.n346 B.n345 10.6151
R554 B.n220 B.n81 10.6151
R555 B.n224 B.n81 10.6151
R556 B.n225 B.n224 10.6151
R557 B.n226 B.n225 10.6151
R558 B.n226 B.n79 10.6151
R559 B.n230 B.n79 10.6151
R560 B.n231 B.n230 10.6151
R561 B.n232 B.n231 10.6151
R562 B.n232 B.n77 10.6151
R563 B.n236 B.n77 10.6151
R564 B.n237 B.n236 10.6151
R565 B.n238 B.n237 10.6151
R566 B.n238 B.n75 10.6151
R567 B.n242 B.n75 10.6151
R568 B.n243 B.n242 10.6151
R569 B.n244 B.n243 10.6151
R570 B.n244 B.n73 10.6151
R571 B.n248 B.n73 10.6151
R572 B.n249 B.n248 10.6151
R573 B.n250 B.n249 10.6151
R574 B.n250 B.n71 10.6151
R575 B.n254 B.n71 10.6151
R576 B.n255 B.n254 10.6151
R577 B.n256 B.n255 10.6151
R578 B.n256 B.n69 10.6151
R579 B.n260 B.n69 10.6151
R580 B.n261 B.n260 10.6151
R581 B.n262 B.n261 10.6151
R582 B.n262 B.n67 10.6151
R583 B.n266 B.n67 10.6151
R584 B.n267 B.n266 10.6151
R585 B.n268 B.n267 10.6151
R586 B.n268 B.n65 10.6151
R587 B.n272 B.n65 10.6151
R588 B.n273 B.n272 10.6151
R589 B.n274 B.n273 10.6151
R590 B.n274 B.n63 10.6151
R591 B.n278 B.n63 10.6151
R592 B.n279 B.n278 10.6151
R593 B.n280 B.n279 10.6151
R594 B.n280 B.n61 10.6151
R595 B.n284 B.n61 10.6151
R596 B.n285 B.n284 10.6151
R597 B.n286 B.n285 10.6151
R598 B.n286 B.n59 10.6151
R599 B.n290 B.n59 10.6151
R600 B.n291 B.n290 10.6151
R601 B.n292 B.n291 10.6151
R602 B.n292 B.n57 10.6151
R603 B.n296 B.n57 10.6151
R604 B.n297 B.n296 10.6151
R605 B.n298 B.n297 10.6151
R606 B.n298 B.n55 10.6151
R607 B.n302 B.n55 10.6151
R608 B.n303 B.n302 10.6151
R609 B.n304 B.n303 10.6151
R610 B.n304 B.n53 10.6151
R611 B.n308 B.n53 10.6151
R612 B.n309 B.n308 10.6151
R613 B.n310 B.n309 10.6151
R614 B.n310 B.n51 10.6151
R615 B.n314 B.n51 10.6151
R616 B.n315 B.n314 10.6151
R617 B.n316 B.n315 10.6151
R618 B.n316 B.n49 10.6151
R619 B.n320 B.n49 10.6151
R620 B.n321 B.n320 10.6151
R621 B.n322 B.n321 10.6151
R622 B.n322 B.n47 10.6151
R623 B.n326 B.n47 10.6151
R624 B.n327 B.n326 10.6151
R625 B.n328 B.n327 10.6151
R626 B.n328 B.n45 10.6151
R627 B.n332 B.n45 10.6151
R628 B.n333 B.n332 10.6151
R629 B.n334 B.n333 10.6151
R630 B.n334 B.n43 10.6151
R631 B.n338 B.n43 10.6151
R632 B.n339 B.n338 10.6151
R633 B.n340 B.n339 10.6151
R634 B.n340 B.n41 10.6151
R635 B.n344 B.n41 10.6151
R636 B.n182 B.n99 10.6151
R637 B.n183 B.n182 10.6151
R638 B.n184 B.n183 10.6151
R639 B.n184 B.n97 10.6151
R640 B.n188 B.n97 10.6151
R641 B.n189 B.n188 10.6151
R642 B.n190 B.n189 10.6151
R643 B.n194 B.n193 10.6151
R644 B.n195 B.n194 10.6151
R645 B.n195 B.n91 10.6151
R646 B.n199 B.n91 10.6151
R647 B.n200 B.n199 10.6151
R648 B.n201 B.n200 10.6151
R649 B.n201 B.n89 10.6151
R650 B.n205 B.n89 10.6151
R651 B.n206 B.n205 10.6151
R652 B.n208 B.n85 10.6151
R653 B.n212 B.n85 10.6151
R654 B.n213 B.n212 10.6151
R655 B.n214 B.n213 10.6151
R656 B.n214 B.n83 10.6151
R657 B.n218 B.n83 10.6151
R658 B.n219 B.n218 10.6151
R659 B.n178 B.n177 10.6151
R660 B.n177 B.n176 10.6151
R661 B.n176 B.n101 10.6151
R662 B.n172 B.n101 10.6151
R663 B.n172 B.n171 10.6151
R664 B.n171 B.n170 10.6151
R665 B.n170 B.n103 10.6151
R666 B.n166 B.n103 10.6151
R667 B.n166 B.n165 10.6151
R668 B.n165 B.n164 10.6151
R669 B.n164 B.n105 10.6151
R670 B.n160 B.n105 10.6151
R671 B.n160 B.n159 10.6151
R672 B.n159 B.n158 10.6151
R673 B.n158 B.n107 10.6151
R674 B.n154 B.n107 10.6151
R675 B.n154 B.n153 10.6151
R676 B.n153 B.n152 10.6151
R677 B.n152 B.n109 10.6151
R678 B.n148 B.n109 10.6151
R679 B.n148 B.n147 10.6151
R680 B.n147 B.n146 10.6151
R681 B.n146 B.n111 10.6151
R682 B.n142 B.n111 10.6151
R683 B.n142 B.n141 10.6151
R684 B.n141 B.n140 10.6151
R685 B.n140 B.n113 10.6151
R686 B.n136 B.n113 10.6151
R687 B.n136 B.n135 10.6151
R688 B.n135 B.n134 10.6151
R689 B.n134 B.n115 10.6151
R690 B.n130 B.n115 10.6151
R691 B.n130 B.n129 10.6151
R692 B.n129 B.n128 10.6151
R693 B.n128 B.n117 10.6151
R694 B.n124 B.n117 10.6151
R695 B.n124 B.n123 10.6151
R696 B.n123 B.n122 10.6151
R697 B.n122 B.n119 10.6151
R698 B.n119 B.n0 10.6151
R699 B.n443 B.n1 10.6151
R700 B.n443 B.n442 10.6151
R701 B.n442 B.n441 10.6151
R702 B.n441 B.n4 10.6151
R703 B.n437 B.n4 10.6151
R704 B.n437 B.n436 10.6151
R705 B.n436 B.n435 10.6151
R706 B.n435 B.n6 10.6151
R707 B.n431 B.n6 10.6151
R708 B.n431 B.n430 10.6151
R709 B.n430 B.n429 10.6151
R710 B.n429 B.n8 10.6151
R711 B.n425 B.n8 10.6151
R712 B.n425 B.n424 10.6151
R713 B.n424 B.n423 10.6151
R714 B.n423 B.n10 10.6151
R715 B.n419 B.n10 10.6151
R716 B.n419 B.n418 10.6151
R717 B.n418 B.n417 10.6151
R718 B.n417 B.n12 10.6151
R719 B.n413 B.n12 10.6151
R720 B.n413 B.n412 10.6151
R721 B.n412 B.n411 10.6151
R722 B.n411 B.n14 10.6151
R723 B.n407 B.n14 10.6151
R724 B.n407 B.n406 10.6151
R725 B.n406 B.n405 10.6151
R726 B.n405 B.n16 10.6151
R727 B.n401 B.n16 10.6151
R728 B.n401 B.n400 10.6151
R729 B.n400 B.n399 10.6151
R730 B.n399 B.n18 10.6151
R731 B.n395 B.n18 10.6151
R732 B.n395 B.n394 10.6151
R733 B.n394 B.n393 10.6151
R734 B.n393 B.n20 10.6151
R735 B.n389 B.n20 10.6151
R736 B.n389 B.n388 10.6151
R737 B.n388 B.n387 10.6151
R738 B.n387 B.n22 10.6151
R739 B.n30 B.n26 9.52245
R740 B.n357 B.n356 9.52245
R741 B.n190 B.n95 9.52245
R742 B.n208 B.n207 9.52245
R743 B.n447 B.n0 2.81026
R744 B.n447 B.n1 2.81026
R745 B.n371 B.n30 1.09318
R746 B.n358 B.n357 1.09318
R747 B.n193 B.n95 1.09318
R748 B.n207 B.n206 1.09318
C0 VP VDD2 0.455747f
C1 B VP 1.73481f
C2 VDD1 w_n3220_n1104# 1.29566f
C3 VTAIL VDD2 3.23436f
C4 B VTAIL 1.18534f
C5 VN VDD1 0.157107f
C6 VP VDD1 0.897162f
C7 B VDD2 1.16937f
C8 VN w_n3220_n1104# 5.41523f
C9 VP w_n3220_n1104# 5.82236f
C10 VTAIL VDD1 3.17466f
C11 VN VP 4.70469f
C12 VTAIL w_n3220_n1104# 1.41864f
C13 VDD2 VDD1 1.22119f
C14 B VDD1 1.1027f
C15 VDD2 w_n3220_n1104# 1.3686f
C16 B w_n3220_n1104# 7.21574f
C17 VN VTAIL 1.58666f
C18 VP VTAIL 1.60077f
C19 VN VDD2 0.601756f
C20 B VN 1.04209f
C21 VDD2 VSUBS 0.815797f
C22 VDD1 VSUBS 4.01483f
C23 VTAIL VSUBS 0.498554f
C24 VN VSUBS 6.4488f
C25 VP VSUBS 2.130111f
C26 B VSUBS 3.787019f
C27 w_n3220_n1104# VSUBS 46.0202f
C28 B.n0 VSUBS 0.007392f
C29 B.n1 VSUBS 0.007392f
C30 B.n2 VSUBS 0.011689f
C31 B.n3 VSUBS 0.011689f
C32 B.n4 VSUBS 0.011689f
C33 B.n5 VSUBS 0.011689f
C34 B.n6 VSUBS 0.011689f
C35 B.n7 VSUBS 0.011689f
C36 B.n8 VSUBS 0.011689f
C37 B.n9 VSUBS 0.011689f
C38 B.n10 VSUBS 0.011689f
C39 B.n11 VSUBS 0.011689f
C40 B.n12 VSUBS 0.011689f
C41 B.n13 VSUBS 0.011689f
C42 B.n14 VSUBS 0.011689f
C43 B.n15 VSUBS 0.011689f
C44 B.n16 VSUBS 0.011689f
C45 B.n17 VSUBS 0.011689f
C46 B.n18 VSUBS 0.011689f
C47 B.n19 VSUBS 0.011689f
C48 B.n20 VSUBS 0.011689f
C49 B.n21 VSUBS 0.011689f
C50 B.n22 VSUBS 0.028359f
C51 B.n23 VSUBS 0.011689f
C52 B.n24 VSUBS 0.011689f
C53 B.n25 VSUBS 0.011689f
C54 B.n26 VSUBS 0.011088f
C55 B.n27 VSUBS 0.011689f
C56 B.t8 VSUBS 0.021581f
C57 B.t7 VSUBS 0.027275f
C58 B.t6 VSUBS 0.195475f
C59 B.n28 VSUBS 0.111897f
C60 B.n29 VSUBS 0.073711f
C61 B.n30 VSUBS 0.027083f
C62 B.n31 VSUBS 0.011689f
C63 B.n32 VSUBS 0.011689f
C64 B.n33 VSUBS 0.011689f
C65 B.n34 VSUBS 0.011689f
C66 B.t11 VSUBS 0.021581f
C67 B.t10 VSUBS 0.027275f
C68 B.t9 VSUBS 0.195662f
C69 B.n35 VSUBS 0.11171f
C70 B.n36 VSUBS 0.073711f
C71 B.n37 VSUBS 0.011689f
C72 B.n38 VSUBS 0.011689f
C73 B.n39 VSUBS 0.011689f
C74 B.n40 VSUBS 0.029744f
C75 B.n41 VSUBS 0.011689f
C76 B.n42 VSUBS 0.011689f
C77 B.n43 VSUBS 0.011689f
C78 B.n44 VSUBS 0.011689f
C79 B.n45 VSUBS 0.011689f
C80 B.n46 VSUBS 0.011689f
C81 B.n47 VSUBS 0.011689f
C82 B.n48 VSUBS 0.011689f
C83 B.n49 VSUBS 0.011689f
C84 B.n50 VSUBS 0.011689f
C85 B.n51 VSUBS 0.011689f
C86 B.n52 VSUBS 0.011689f
C87 B.n53 VSUBS 0.011689f
C88 B.n54 VSUBS 0.011689f
C89 B.n55 VSUBS 0.011689f
C90 B.n56 VSUBS 0.011689f
C91 B.n57 VSUBS 0.011689f
C92 B.n58 VSUBS 0.011689f
C93 B.n59 VSUBS 0.011689f
C94 B.n60 VSUBS 0.011689f
C95 B.n61 VSUBS 0.011689f
C96 B.n62 VSUBS 0.011689f
C97 B.n63 VSUBS 0.011689f
C98 B.n64 VSUBS 0.011689f
C99 B.n65 VSUBS 0.011689f
C100 B.n66 VSUBS 0.011689f
C101 B.n67 VSUBS 0.011689f
C102 B.n68 VSUBS 0.011689f
C103 B.n69 VSUBS 0.011689f
C104 B.n70 VSUBS 0.011689f
C105 B.n71 VSUBS 0.011689f
C106 B.n72 VSUBS 0.011689f
C107 B.n73 VSUBS 0.011689f
C108 B.n74 VSUBS 0.011689f
C109 B.n75 VSUBS 0.011689f
C110 B.n76 VSUBS 0.011689f
C111 B.n77 VSUBS 0.011689f
C112 B.n78 VSUBS 0.011689f
C113 B.n79 VSUBS 0.011689f
C114 B.n80 VSUBS 0.011689f
C115 B.n81 VSUBS 0.011689f
C116 B.n82 VSUBS 0.029744f
C117 B.n83 VSUBS 0.011689f
C118 B.n84 VSUBS 0.011689f
C119 B.n85 VSUBS 0.011689f
C120 B.n86 VSUBS 0.011689f
C121 B.t1 VSUBS 0.021581f
C122 B.t2 VSUBS 0.027275f
C123 B.t0 VSUBS 0.195662f
C124 B.n87 VSUBS 0.11171f
C125 B.n88 VSUBS 0.073711f
C126 B.n89 VSUBS 0.011689f
C127 B.n90 VSUBS 0.011689f
C128 B.n91 VSUBS 0.011689f
C129 B.n92 VSUBS 0.011689f
C130 B.t4 VSUBS 0.021581f
C131 B.t5 VSUBS 0.027275f
C132 B.t3 VSUBS 0.195475f
C133 B.n93 VSUBS 0.111897f
C134 B.n94 VSUBS 0.073711f
C135 B.n95 VSUBS 0.027083f
C136 B.n96 VSUBS 0.011689f
C137 B.n97 VSUBS 0.011689f
C138 B.n98 VSUBS 0.011689f
C139 B.n99 VSUBS 0.029744f
C140 B.n100 VSUBS 0.011689f
C141 B.n101 VSUBS 0.011689f
C142 B.n102 VSUBS 0.011689f
C143 B.n103 VSUBS 0.011689f
C144 B.n104 VSUBS 0.011689f
C145 B.n105 VSUBS 0.011689f
C146 B.n106 VSUBS 0.011689f
C147 B.n107 VSUBS 0.011689f
C148 B.n108 VSUBS 0.011689f
C149 B.n109 VSUBS 0.011689f
C150 B.n110 VSUBS 0.011689f
C151 B.n111 VSUBS 0.011689f
C152 B.n112 VSUBS 0.011689f
C153 B.n113 VSUBS 0.011689f
C154 B.n114 VSUBS 0.011689f
C155 B.n115 VSUBS 0.011689f
C156 B.n116 VSUBS 0.011689f
C157 B.n117 VSUBS 0.011689f
C158 B.n118 VSUBS 0.011689f
C159 B.n119 VSUBS 0.011689f
C160 B.n120 VSUBS 0.011689f
C161 B.n121 VSUBS 0.011689f
C162 B.n122 VSUBS 0.011689f
C163 B.n123 VSUBS 0.011689f
C164 B.n124 VSUBS 0.011689f
C165 B.n125 VSUBS 0.011689f
C166 B.n126 VSUBS 0.011689f
C167 B.n127 VSUBS 0.011689f
C168 B.n128 VSUBS 0.011689f
C169 B.n129 VSUBS 0.011689f
C170 B.n130 VSUBS 0.011689f
C171 B.n131 VSUBS 0.011689f
C172 B.n132 VSUBS 0.011689f
C173 B.n133 VSUBS 0.011689f
C174 B.n134 VSUBS 0.011689f
C175 B.n135 VSUBS 0.011689f
C176 B.n136 VSUBS 0.011689f
C177 B.n137 VSUBS 0.011689f
C178 B.n138 VSUBS 0.011689f
C179 B.n139 VSUBS 0.011689f
C180 B.n140 VSUBS 0.011689f
C181 B.n141 VSUBS 0.011689f
C182 B.n142 VSUBS 0.011689f
C183 B.n143 VSUBS 0.011689f
C184 B.n144 VSUBS 0.011689f
C185 B.n145 VSUBS 0.011689f
C186 B.n146 VSUBS 0.011689f
C187 B.n147 VSUBS 0.011689f
C188 B.n148 VSUBS 0.011689f
C189 B.n149 VSUBS 0.011689f
C190 B.n150 VSUBS 0.011689f
C191 B.n151 VSUBS 0.011689f
C192 B.n152 VSUBS 0.011689f
C193 B.n153 VSUBS 0.011689f
C194 B.n154 VSUBS 0.011689f
C195 B.n155 VSUBS 0.011689f
C196 B.n156 VSUBS 0.011689f
C197 B.n157 VSUBS 0.011689f
C198 B.n158 VSUBS 0.011689f
C199 B.n159 VSUBS 0.011689f
C200 B.n160 VSUBS 0.011689f
C201 B.n161 VSUBS 0.011689f
C202 B.n162 VSUBS 0.011689f
C203 B.n163 VSUBS 0.011689f
C204 B.n164 VSUBS 0.011689f
C205 B.n165 VSUBS 0.011689f
C206 B.n166 VSUBS 0.011689f
C207 B.n167 VSUBS 0.011689f
C208 B.n168 VSUBS 0.011689f
C209 B.n169 VSUBS 0.011689f
C210 B.n170 VSUBS 0.011689f
C211 B.n171 VSUBS 0.011689f
C212 B.n172 VSUBS 0.011689f
C213 B.n173 VSUBS 0.011689f
C214 B.n174 VSUBS 0.011689f
C215 B.n175 VSUBS 0.011689f
C216 B.n176 VSUBS 0.011689f
C217 B.n177 VSUBS 0.011689f
C218 B.n178 VSUBS 0.028359f
C219 B.n179 VSUBS 0.028359f
C220 B.n180 VSUBS 0.029744f
C221 B.n181 VSUBS 0.011689f
C222 B.n182 VSUBS 0.011689f
C223 B.n183 VSUBS 0.011689f
C224 B.n184 VSUBS 0.011689f
C225 B.n185 VSUBS 0.011689f
C226 B.n186 VSUBS 0.011689f
C227 B.n187 VSUBS 0.011689f
C228 B.n188 VSUBS 0.011689f
C229 B.n189 VSUBS 0.011689f
C230 B.n190 VSUBS 0.011088f
C231 B.n191 VSUBS 0.011689f
C232 B.n192 VSUBS 0.011689f
C233 B.n193 VSUBS 0.006446f
C234 B.n194 VSUBS 0.011689f
C235 B.n195 VSUBS 0.011689f
C236 B.n196 VSUBS 0.011689f
C237 B.n197 VSUBS 0.011689f
C238 B.n198 VSUBS 0.011689f
C239 B.n199 VSUBS 0.011689f
C240 B.n200 VSUBS 0.011689f
C241 B.n201 VSUBS 0.011689f
C242 B.n202 VSUBS 0.011689f
C243 B.n203 VSUBS 0.011689f
C244 B.n204 VSUBS 0.011689f
C245 B.n205 VSUBS 0.011689f
C246 B.n206 VSUBS 0.006446f
C247 B.n207 VSUBS 0.027083f
C248 B.n208 VSUBS 0.011088f
C249 B.n209 VSUBS 0.011689f
C250 B.n210 VSUBS 0.011689f
C251 B.n211 VSUBS 0.011689f
C252 B.n212 VSUBS 0.011689f
C253 B.n213 VSUBS 0.011689f
C254 B.n214 VSUBS 0.011689f
C255 B.n215 VSUBS 0.011689f
C256 B.n216 VSUBS 0.011689f
C257 B.n217 VSUBS 0.011689f
C258 B.n218 VSUBS 0.011689f
C259 B.n219 VSUBS 0.029744f
C260 B.n220 VSUBS 0.028359f
C261 B.n221 VSUBS 0.028359f
C262 B.n222 VSUBS 0.011689f
C263 B.n223 VSUBS 0.011689f
C264 B.n224 VSUBS 0.011689f
C265 B.n225 VSUBS 0.011689f
C266 B.n226 VSUBS 0.011689f
C267 B.n227 VSUBS 0.011689f
C268 B.n228 VSUBS 0.011689f
C269 B.n229 VSUBS 0.011689f
C270 B.n230 VSUBS 0.011689f
C271 B.n231 VSUBS 0.011689f
C272 B.n232 VSUBS 0.011689f
C273 B.n233 VSUBS 0.011689f
C274 B.n234 VSUBS 0.011689f
C275 B.n235 VSUBS 0.011689f
C276 B.n236 VSUBS 0.011689f
C277 B.n237 VSUBS 0.011689f
C278 B.n238 VSUBS 0.011689f
C279 B.n239 VSUBS 0.011689f
C280 B.n240 VSUBS 0.011689f
C281 B.n241 VSUBS 0.011689f
C282 B.n242 VSUBS 0.011689f
C283 B.n243 VSUBS 0.011689f
C284 B.n244 VSUBS 0.011689f
C285 B.n245 VSUBS 0.011689f
C286 B.n246 VSUBS 0.011689f
C287 B.n247 VSUBS 0.011689f
C288 B.n248 VSUBS 0.011689f
C289 B.n249 VSUBS 0.011689f
C290 B.n250 VSUBS 0.011689f
C291 B.n251 VSUBS 0.011689f
C292 B.n252 VSUBS 0.011689f
C293 B.n253 VSUBS 0.011689f
C294 B.n254 VSUBS 0.011689f
C295 B.n255 VSUBS 0.011689f
C296 B.n256 VSUBS 0.011689f
C297 B.n257 VSUBS 0.011689f
C298 B.n258 VSUBS 0.011689f
C299 B.n259 VSUBS 0.011689f
C300 B.n260 VSUBS 0.011689f
C301 B.n261 VSUBS 0.011689f
C302 B.n262 VSUBS 0.011689f
C303 B.n263 VSUBS 0.011689f
C304 B.n264 VSUBS 0.011689f
C305 B.n265 VSUBS 0.011689f
C306 B.n266 VSUBS 0.011689f
C307 B.n267 VSUBS 0.011689f
C308 B.n268 VSUBS 0.011689f
C309 B.n269 VSUBS 0.011689f
C310 B.n270 VSUBS 0.011689f
C311 B.n271 VSUBS 0.011689f
C312 B.n272 VSUBS 0.011689f
C313 B.n273 VSUBS 0.011689f
C314 B.n274 VSUBS 0.011689f
C315 B.n275 VSUBS 0.011689f
C316 B.n276 VSUBS 0.011689f
C317 B.n277 VSUBS 0.011689f
C318 B.n278 VSUBS 0.011689f
C319 B.n279 VSUBS 0.011689f
C320 B.n280 VSUBS 0.011689f
C321 B.n281 VSUBS 0.011689f
C322 B.n282 VSUBS 0.011689f
C323 B.n283 VSUBS 0.011689f
C324 B.n284 VSUBS 0.011689f
C325 B.n285 VSUBS 0.011689f
C326 B.n286 VSUBS 0.011689f
C327 B.n287 VSUBS 0.011689f
C328 B.n288 VSUBS 0.011689f
C329 B.n289 VSUBS 0.011689f
C330 B.n290 VSUBS 0.011689f
C331 B.n291 VSUBS 0.011689f
C332 B.n292 VSUBS 0.011689f
C333 B.n293 VSUBS 0.011689f
C334 B.n294 VSUBS 0.011689f
C335 B.n295 VSUBS 0.011689f
C336 B.n296 VSUBS 0.011689f
C337 B.n297 VSUBS 0.011689f
C338 B.n298 VSUBS 0.011689f
C339 B.n299 VSUBS 0.011689f
C340 B.n300 VSUBS 0.011689f
C341 B.n301 VSUBS 0.011689f
C342 B.n302 VSUBS 0.011689f
C343 B.n303 VSUBS 0.011689f
C344 B.n304 VSUBS 0.011689f
C345 B.n305 VSUBS 0.011689f
C346 B.n306 VSUBS 0.011689f
C347 B.n307 VSUBS 0.011689f
C348 B.n308 VSUBS 0.011689f
C349 B.n309 VSUBS 0.011689f
C350 B.n310 VSUBS 0.011689f
C351 B.n311 VSUBS 0.011689f
C352 B.n312 VSUBS 0.011689f
C353 B.n313 VSUBS 0.011689f
C354 B.n314 VSUBS 0.011689f
C355 B.n315 VSUBS 0.011689f
C356 B.n316 VSUBS 0.011689f
C357 B.n317 VSUBS 0.011689f
C358 B.n318 VSUBS 0.011689f
C359 B.n319 VSUBS 0.011689f
C360 B.n320 VSUBS 0.011689f
C361 B.n321 VSUBS 0.011689f
C362 B.n322 VSUBS 0.011689f
C363 B.n323 VSUBS 0.011689f
C364 B.n324 VSUBS 0.011689f
C365 B.n325 VSUBS 0.011689f
C366 B.n326 VSUBS 0.011689f
C367 B.n327 VSUBS 0.011689f
C368 B.n328 VSUBS 0.011689f
C369 B.n329 VSUBS 0.011689f
C370 B.n330 VSUBS 0.011689f
C371 B.n331 VSUBS 0.011689f
C372 B.n332 VSUBS 0.011689f
C373 B.n333 VSUBS 0.011689f
C374 B.n334 VSUBS 0.011689f
C375 B.n335 VSUBS 0.011689f
C376 B.n336 VSUBS 0.011689f
C377 B.n337 VSUBS 0.011689f
C378 B.n338 VSUBS 0.011689f
C379 B.n339 VSUBS 0.011689f
C380 B.n340 VSUBS 0.011689f
C381 B.n341 VSUBS 0.011689f
C382 B.n342 VSUBS 0.011689f
C383 B.n343 VSUBS 0.028359f
C384 B.n344 VSUBS 0.029621f
C385 B.n345 VSUBS 0.028482f
C386 B.n346 VSUBS 0.011689f
C387 B.n347 VSUBS 0.011689f
C388 B.n348 VSUBS 0.011689f
C389 B.n349 VSUBS 0.011689f
C390 B.n350 VSUBS 0.011689f
C391 B.n351 VSUBS 0.011689f
C392 B.n352 VSUBS 0.011689f
C393 B.n353 VSUBS 0.011689f
C394 B.n354 VSUBS 0.011689f
C395 B.n355 VSUBS 0.011689f
C396 B.n356 VSUBS 0.011088f
C397 B.n357 VSUBS 0.027083f
C398 B.n358 VSUBS 0.006446f
C399 B.n359 VSUBS 0.011689f
C400 B.n360 VSUBS 0.011689f
C401 B.n361 VSUBS 0.011689f
C402 B.n362 VSUBS 0.011689f
C403 B.n363 VSUBS 0.011689f
C404 B.n364 VSUBS 0.011689f
C405 B.n365 VSUBS 0.011689f
C406 B.n366 VSUBS 0.011689f
C407 B.n367 VSUBS 0.011689f
C408 B.n368 VSUBS 0.011689f
C409 B.n369 VSUBS 0.011689f
C410 B.n370 VSUBS 0.011689f
C411 B.n371 VSUBS 0.006446f
C412 B.n372 VSUBS 0.011689f
C413 B.n373 VSUBS 0.011689f
C414 B.n374 VSUBS 0.011689f
C415 B.n375 VSUBS 0.011689f
C416 B.n376 VSUBS 0.011689f
C417 B.n377 VSUBS 0.011689f
C418 B.n378 VSUBS 0.011689f
C419 B.n379 VSUBS 0.011689f
C420 B.n380 VSUBS 0.011689f
C421 B.n381 VSUBS 0.011689f
C422 B.n382 VSUBS 0.011689f
C423 B.n383 VSUBS 0.029744f
C424 B.n384 VSUBS 0.029744f
C425 B.n385 VSUBS 0.028359f
C426 B.n386 VSUBS 0.011689f
C427 B.n387 VSUBS 0.011689f
C428 B.n388 VSUBS 0.011689f
C429 B.n389 VSUBS 0.011689f
C430 B.n390 VSUBS 0.011689f
C431 B.n391 VSUBS 0.011689f
C432 B.n392 VSUBS 0.011689f
C433 B.n393 VSUBS 0.011689f
C434 B.n394 VSUBS 0.011689f
C435 B.n395 VSUBS 0.011689f
C436 B.n396 VSUBS 0.011689f
C437 B.n397 VSUBS 0.011689f
C438 B.n398 VSUBS 0.011689f
C439 B.n399 VSUBS 0.011689f
C440 B.n400 VSUBS 0.011689f
C441 B.n401 VSUBS 0.011689f
C442 B.n402 VSUBS 0.011689f
C443 B.n403 VSUBS 0.011689f
C444 B.n404 VSUBS 0.011689f
C445 B.n405 VSUBS 0.011689f
C446 B.n406 VSUBS 0.011689f
C447 B.n407 VSUBS 0.011689f
C448 B.n408 VSUBS 0.011689f
C449 B.n409 VSUBS 0.011689f
C450 B.n410 VSUBS 0.011689f
C451 B.n411 VSUBS 0.011689f
C452 B.n412 VSUBS 0.011689f
C453 B.n413 VSUBS 0.011689f
C454 B.n414 VSUBS 0.011689f
C455 B.n415 VSUBS 0.011689f
C456 B.n416 VSUBS 0.011689f
C457 B.n417 VSUBS 0.011689f
C458 B.n418 VSUBS 0.011689f
C459 B.n419 VSUBS 0.011689f
C460 B.n420 VSUBS 0.011689f
C461 B.n421 VSUBS 0.011689f
C462 B.n422 VSUBS 0.011689f
C463 B.n423 VSUBS 0.011689f
C464 B.n424 VSUBS 0.011689f
C465 B.n425 VSUBS 0.011689f
C466 B.n426 VSUBS 0.011689f
C467 B.n427 VSUBS 0.011689f
C468 B.n428 VSUBS 0.011689f
C469 B.n429 VSUBS 0.011689f
C470 B.n430 VSUBS 0.011689f
C471 B.n431 VSUBS 0.011689f
C472 B.n432 VSUBS 0.011689f
C473 B.n433 VSUBS 0.011689f
C474 B.n434 VSUBS 0.011689f
C475 B.n435 VSUBS 0.011689f
C476 B.n436 VSUBS 0.011689f
C477 B.n437 VSUBS 0.011689f
C478 B.n438 VSUBS 0.011689f
C479 B.n439 VSUBS 0.011689f
C480 B.n440 VSUBS 0.011689f
C481 B.n441 VSUBS 0.011689f
C482 B.n442 VSUBS 0.011689f
C483 B.n443 VSUBS 0.011689f
C484 B.n444 VSUBS 0.011689f
C485 B.n445 VSUBS 0.011689f
C486 B.n446 VSUBS 0.011689f
C487 B.n447 VSUBS 0.026469f
C488 VDD2.t0 VSUBS 0.014897f
C489 VDD2.t1 VSUBS 0.014897f
C490 VDD2.n0 VSUBS 0.076463f
C491 VDD2.t3 VSUBS 0.014897f
C492 VDD2.t2 VSUBS 0.014897f
C493 VDD2.n1 VSUBS 0.032477f
C494 VDD2.n2 VSUBS 2.73672f
C495 VN.t2 VSUBS 0.695576f
C496 VN.t3 VSUBS 0.718714f
C497 VN.n0 VSUBS 0.668572f
C498 VN.t1 VSUBS 0.718714f
C499 VN.t0 VSUBS 0.695576f
C500 VN.n1 VSUBS 3.4526f
C501 VDD1.t2 VSUBS 0.014435f
C502 VDD1.t3 VSUBS 0.014435f
C503 VDD1.n0 VSUBS 0.031504f
C504 VDD1.t1 VSUBS 0.014435f
C505 VDD1.t0 VSUBS 0.014435f
C506 VDD1.n1 VSUBS 0.077505f
C507 VTAIL.t3 VSUBS 0.068983f
C508 VTAIL.n0 VSUBS 0.24117f
C509 VTAIL.t4 VSUBS 0.068983f
C510 VTAIL.n1 VSUBS 0.384089f
C511 VTAIL.t6 VSUBS 0.068983f
C512 VTAIL.n2 VSUBS 1.07794f
C513 VTAIL.t1 VSUBS 0.068983f
C514 VTAIL.n3 VSUBS 1.07794f
C515 VTAIL.t0 VSUBS 0.068983f
C516 VTAIL.n4 VSUBS 0.384089f
C517 VTAIL.t7 VSUBS 0.068983f
C518 VTAIL.n5 VSUBS 0.384089f
C519 VTAIL.t5 VSUBS 0.068983f
C520 VTAIL.n6 VSUBS 1.07794f
C521 VTAIL.t2 VSUBS 0.068983f
C522 VTAIL.n7 VSUBS 0.92435f
C523 VP.t3 VSUBS 0.193221f
C524 VP.n0 VSUBS 0.396288f
C525 VP.n1 VSUBS 0.059294f
C526 VP.n2 VSUBS 0.086935f
C527 VP.n3 VSUBS 0.059294f
C528 VP.n4 VSUBS 0.069936f
C529 VP.t1 VSUBS 0.753107f
C530 VP.t0 VSUBS 0.728864f
C531 VP.n5 VSUBS 3.59225f
C532 VP.t2 VSUBS 0.193221f
C533 VP.n6 VSUBS 0.396288f
C534 VP.n7 VSUBS 2.66842f
C535 VP.n8 VSUBS 0.095714f
C536 VP.n9 VSUBS 0.059294f
C537 VP.n10 VSUBS 0.111063f
C538 VP.n11 VSUBS 0.111063f
C539 VP.n12 VSUBS 0.086935f
C540 VP.n13 VSUBS 0.059294f
C541 VP.n14 VSUBS 0.059294f
C542 VP.n15 VSUBS 0.059294f
C543 VP.n16 VSUBS 0.111063f
C544 VP.n17 VSUBS 0.111063f
C545 VP.n18 VSUBS 0.069936f
C546 VP.n19 VSUBS 0.095714f
C547 VP.n20 VSUBS 0.16455f
.ends

