* NGSPICE file created from diff_pair_sample_1718.ext - technology: sky130A

.subckt diff_pair_sample_1718 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=3.67
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=3.67
X2 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=3.67
X3 VTAIL.t5 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=3.67
X4 VTAIL.t7 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=3.67
X5 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=3.67
X6 VDD1.t3 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=3.67
X7 VDD1.t2 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=3.67
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=3.67
X9 VDD2.t3 VN.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=3.67
X10 VDD2.t2 VN.t3 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=3.67
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=3.67
X12 VTAIL.t1 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=3.67
X13 VTAIL.t9 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=3.67
X14 VDD2.t0 VN.t5 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=3.67
X15 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=3.67
R0 VN.n33 VN.n18 161.3
R1 VN.n32 VN.n31 161.3
R2 VN.n30 VN.n19 161.3
R3 VN.n29 VN.n28 161.3
R4 VN.n27 VN.n20 161.3
R5 VN.n26 VN.n25 161.3
R6 VN.n24 VN.n21 161.3
R7 VN.n15 VN.n0 161.3
R8 VN.n14 VN.n13 161.3
R9 VN.n12 VN.n1 161.3
R10 VN.n11 VN.n10 161.3
R11 VN.n9 VN.n2 161.3
R12 VN.n8 VN.n7 161.3
R13 VN.n6 VN.n3 161.3
R14 VN.n5 VN.t3 62.2517
R15 VN.n23 VN.t2 62.2517
R16 VN.n17 VN.n16 57.7148
R17 VN.n35 VN.n34 57.7148
R18 VN.n5 VN.n4 50.4779
R19 VN.n23 VN.n22 50.4779
R20 VN VN.n35 47.5269
R21 VN.n10 VN.n9 40.4934
R22 VN.n10 VN.n1 40.4934
R23 VN.n28 VN.n27 40.4934
R24 VN.n28 VN.n19 40.4934
R25 VN.n16 VN.t0 30.1419
R26 VN.n4 VN.t4 30.1419
R27 VN.n34 VN.t5 30.1419
R28 VN.n22 VN.t1 30.1419
R29 VN.n4 VN.n3 24.4675
R30 VN.n8 VN.n3 24.4675
R31 VN.n9 VN.n8 24.4675
R32 VN.n14 VN.n1 24.4675
R33 VN.n15 VN.n14 24.4675
R34 VN.n16 VN.n15 24.4675
R35 VN.n27 VN.n26 24.4675
R36 VN.n26 VN.n21 24.4675
R37 VN.n22 VN.n21 24.4675
R38 VN.n34 VN.n33 24.4675
R39 VN.n33 VN.n32 24.4675
R40 VN.n32 VN.n19 24.4675
R41 VN.n24 VN.n23 2.5265
R42 VN.n6 VN.n5 2.5265
R43 VN.n35 VN.n18 0.417535
R44 VN.n17 VN.n0 0.417535
R45 VN VN.n17 0.394291
R46 VN.n31 VN.n18 0.189894
R47 VN.n31 VN.n30 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n20 0.189894
R50 VN.n25 VN.n20 0.189894
R51 VN.n25 VN.n24 0.189894
R52 VN.n7 VN.n6 0.189894
R53 VN.n7 VN.n2 0.189894
R54 VN.n11 VN.n2 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n13 VN.n12 0.189894
R57 VN.n13 VN.n0 0.189894
R58 VTAIL.n98 VTAIL.n80 289.615
R59 VTAIL.n20 VTAIL.n2 289.615
R60 VTAIL.n74 VTAIL.n56 289.615
R61 VTAIL.n48 VTAIL.n30 289.615
R62 VTAIL.n89 VTAIL.n88 185
R63 VTAIL.n91 VTAIL.n90 185
R64 VTAIL.n84 VTAIL.n83 185
R65 VTAIL.n97 VTAIL.n96 185
R66 VTAIL.n99 VTAIL.n98 185
R67 VTAIL.n11 VTAIL.n10 185
R68 VTAIL.n13 VTAIL.n12 185
R69 VTAIL.n6 VTAIL.n5 185
R70 VTAIL.n19 VTAIL.n18 185
R71 VTAIL.n21 VTAIL.n20 185
R72 VTAIL.n75 VTAIL.n74 185
R73 VTAIL.n73 VTAIL.n72 185
R74 VTAIL.n60 VTAIL.n59 185
R75 VTAIL.n67 VTAIL.n66 185
R76 VTAIL.n65 VTAIL.n64 185
R77 VTAIL.n49 VTAIL.n48 185
R78 VTAIL.n47 VTAIL.n46 185
R79 VTAIL.n34 VTAIL.n33 185
R80 VTAIL.n41 VTAIL.n40 185
R81 VTAIL.n39 VTAIL.n38 185
R82 VTAIL.n87 VTAIL.t10 147.714
R83 VTAIL.n9 VTAIL.t3 147.714
R84 VTAIL.n63 VTAIL.t2 147.714
R85 VTAIL.n37 VTAIL.t11 147.714
R86 VTAIL.n90 VTAIL.n89 104.615
R87 VTAIL.n90 VTAIL.n83 104.615
R88 VTAIL.n97 VTAIL.n83 104.615
R89 VTAIL.n98 VTAIL.n97 104.615
R90 VTAIL.n12 VTAIL.n11 104.615
R91 VTAIL.n12 VTAIL.n5 104.615
R92 VTAIL.n19 VTAIL.n5 104.615
R93 VTAIL.n20 VTAIL.n19 104.615
R94 VTAIL.n74 VTAIL.n73 104.615
R95 VTAIL.n73 VTAIL.n59 104.615
R96 VTAIL.n66 VTAIL.n59 104.615
R97 VTAIL.n66 VTAIL.n65 104.615
R98 VTAIL.n48 VTAIL.n47 104.615
R99 VTAIL.n47 VTAIL.n33 104.615
R100 VTAIL.n40 VTAIL.n33 104.615
R101 VTAIL.n40 VTAIL.n39 104.615
R102 VTAIL.n55 VTAIL.n54 54.5448
R103 VTAIL.n29 VTAIL.n28 54.5448
R104 VTAIL.n1 VTAIL.n0 54.5447
R105 VTAIL.n27 VTAIL.n26 54.5447
R106 VTAIL.n89 VTAIL.t10 52.3082
R107 VTAIL.n11 VTAIL.t3 52.3082
R108 VTAIL.n65 VTAIL.t2 52.3082
R109 VTAIL.n39 VTAIL.t11 52.3082
R110 VTAIL.n103 VTAIL.n102 32.7672
R111 VTAIL.n25 VTAIL.n24 32.7672
R112 VTAIL.n79 VTAIL.n78 32.7672
R113 VTAIL.n53 VTAIL.n52 32.7672
R114 VTAIL.n29 VTAIL.n27 23.2203
R115 VTAIL.n103 VTAIL.n79 19.7721
R116 VTAIL.n88 VTAIL.n87 15.6631
R117 VTAIL.n10 VTAIL.n9 15.6631
R118 VTAIL.n64 VTAIL.n63 15.6631
R119 VTAIL.n38 VTAIL.n37 15.6631
R120 VTAIL.n91 VTAIL.n86 12.8005
R121 VTAIL.n13 VTAIL.n8 12.8005
R122 VTAIL.n67 VTAIL.n62 12.8005
R123 VTAIL.n41 VTAIL.n36 12.8005
R124 VTAIL.n92 VTAIL.n84 12.0247
R125 VTAIL.n14 VTAIL.n6 12.0247
R126 VTAIL.n68 VTAIL.n60 12.0247
R127 VTAIL.n42 VTAIL.n34 12.0247
R128 VTAIL.n96 VTAIL.n95 11.249
R129 VTAIL.n18 VTAIL.n17 11.249
R130 VTAIL.n72 VTAIL.n71 11.249
R131 VTAIL.n46 VTAIL.n45 11.249
R132 VTAIL.n99 VTAIL.n82 10.4732
R133 VTAIL.n21 VTAIL.n4 10.4732
R134 VTAIL.n75 VTAIL.n58 10.4732
R135 VTAIL.n49 VTAIL.n32 10.4732
R136 VTAIL.n100 VTAIL.n80 9.69747
R137 VTAIL.n22 VTAIL.n2 9.69747
R138 VTAIL.n76 VTAIL.n56 9.69747
R139 VTAIL.n50 VTAIL.n30 9.69747
R140 VTAIL.n102 VTAIL.n101 9.45567
R141 VTAIL.n24 VTAIL.n23 9.45567
R142 VTAIL.n78 VTAIL.n77 9.45567
R143 VTAIL.n52 VTAIL.n51 9.45567
R144 VTAIL.n101 VTAIL.n100 9.3005
R145 VTAIL.n82 VTAIL.n81 9.3005
R146 VTAIL.n95 VTAIL.n94 9.3005
R147 VTAIL.n93 VTAIL.n92 9.3005
R148 VTAIL.n86 VTAIL.n85 9.3005
R149 VTAIL.n23 VTAIL.n22 9.3005
R150 VTAIL.n4 VTAIL.n3 9.3005
R151 VTAIL.n17 VTAIL.n16 9.3005
R152 VTAIL.n15 VTAIL.n14 9.3005
R153 VTAIL.n8 VTAIL.n7 9.3005
R154 VTAIL.n77 VTAIL.n76 9.3005
R155 VTAIL.n58 VTAIL.n57 9.3005
R156 VTAIL.n71 VTAIL.n70 9.3005
R157 VTAIL.n69 VTAIL.n68 9.3005
R158 VTAIL.n62 VTAIL.n61 9.3005
R159 VTAIL.n51 VTAIL.n50 9.3005
R160 VTAIL.n32 VTAIL.n31 9.3005
R161 VTAIL.n45 VTAIL.n44 9.3005
R162 VTAIL.n43 VTAIL.n42 9.3005
R163 VTAIL.n36 VTAIL.n35 9.3005
R164 VTAIL.n87 VTAIL.n85 4.39059
R165 VTAIL.n9 VTAIL.n7 4.39059
R166 VTAIL.n63 VTAIL.n61 4.39059
R167 VTAIL.n37 VTAIL.n35 4.39059
R168 VTAIL.n0 VTAIL.t6 4.31423
R169 VTAIL.n0 VTAIL.t9 4.31423
R170 VTAIL.n26 VTAIL.t4 4.31423
R171 VTAIL.n26 VTAIL.t5 4.31423
R172 VTAIL.n54 VTAIL.t0 4.31423
R173 VTAIL.n54 VTAIL.t1 4.31423
R174 VTAIL.n28 VTAIL.t8 4.31423
R175 VTAIL.n28 VTAIL.t7 4.31423
R176 VTAIL.n102 VTAIL.n80 4.26717
R177 VTAIL.n24 VTAIL.n2 4.26717
R178 VTAIL.n78 VTAIL.n56 4.26717
R179 VTAIL.n52 VTAIL.n30 4.26717
R180 VTAIL.n100 VTAIL.n99 3.49141
R181 VTAIL.n22 VTAIL.n21 3.49141
R182 VTAIL.n76 VTAIL.n75 3.49141
R183 VTAIL.n50 VTAIL.n49 3.49141
R184 VTAIL.n53 VTAIL.n29 3.44878
R185 VTAIL.n79 VTAIL.n55 3.44878
R186 VTAIL.n27 VTAIL.n25 3.44878
R187 VTAIL.n96 VTAIL.n82 2.71565
R188 VTAIL.n18 VTAIL.n4 2.71565
R189 VTAIL.n72 VTAIL.n58 2.71565
R190 VTAIL.n46 VTAIL.n32 2.71565
R191 VTAIL VTAIL.n103 2.52852
R192 VTAIL.n55 VTAIL.n53 2.19447
R193 VTAIL.n25 VTAIL.n1 2.19447
R194 VTAIL.n95 VTAIL.n84 1.93989
R195 VTAIL.n17 VTAIL.n6 1.93989
R196 VTAIL.n71 VTAIL.n60 1.93989
R197 VTAIL.n45 VTAIL.n34 1.93989
R198 VTAIL.n92 VTAIL.n91 1.16414
R199 VTAIL.n14 VTAIL.n13 1.16414
R200 VTAIL.n68 VTAIL.n67 1.16414
R201 VTAIL.n42 VTAIL.n41 1.16414
R202 VTAIL VTAIL.n1 0.920759
R203 VTAIL.n88 VTAIL.n86 0.388379
R204 VTAIL.n10 VTAIL.n8 0.388379
R205 VTAIL.n64 VTAIL.n62 0.388379
R206 VTAIL.n38 VTAIL.n36 0.388379
R207 VTAIL.n93 VTAIL.n85 0.155672
R208 VTAIL.n94 VTAIL.n93 0.155672
R209 VTAIL.n94 VTAIL.n81 0.155672
R210 VTAIL.n101 VTAIL.n81 0.155672
R211 VTAIL.n15 VTAIL.n7 0.155672
R212 VTAIL.n16 VTAIL.n15 0.155672
R213 VTAIL.n16 VTAIL.n3 0.155672
R214 VTAIL.n23 VTAIL.n3 0.155672
R215 VTAIL.n77 VTAIL.n57 0.155672
R216 VTAIL.n70 VTAIL.n57 0.155672
R217 VTAIL.n70 VTAIL.n69 0.155672
R218 VTAIL.n69 VTAIL.n61 0.155672
R219 VTAIL.n51 VTAIL.n31 0.155672
R220 VTAIL.n44 VTAIL.n31 0.155672
R221 VTAIL.n44 VTAIL.n43 0.155672
R222 VTAIL.n43 VTAIL.n35 0.155672
R223 VDD2.n43 VDD2.n25 289.615
R224 VDD2.n18 VDD2.n0 289.615
R225 VDD2.n44 VDD2.n43 185
R226 VDD2.n42 VDD2.n41 185
R227 VDD2.n29 VDD2.n28 185
R228 VDD2.n36 VDD2.n35 185
R229 VDD2.n34 VDD2.n33 185
R230 VDD2.n9 VDD2.n8 185
R231 VDD2.n11 VDD2.n10 185
R232 VDD2.n4 VDD2.n3 185
R233 VDD2.n17 VDD2.n16 185
R234 VDD2.n19 VDD2.n18 185
R235 VDD2.n32 VDD2.t0 147.714
R236 VDD2.n7 VDD2.t2 147.714
R237 VDD2.n43 VDD2.n42 104.615
R238 VDD2.n42 VDD2.n28 104.615
R239 VDD2.n35 VDD2.n28 104.615
R240 VDD2.n35 VDD2.n34 104.615
R241 VDD2.n10 VDD2.n9 104.615
R242 VDD2.n10 VDD2.n3 104.615
R243 VDD2.n17 VDD2.n3 104.615
R244 VDD2.n18 VDD2.n17 104.615
R245 VDD2.n24 VDD2.n23 72.0302
R246 VDD2 VDD2.n49 72.0273
R247 VDD2.n34 VDD2.t0 52.3082
R248 VDD2.n9 VDD2.t2 52.3082
R249 VDD2.n24 VDD2.n22 51.9768
R250 VDD2.n48 VDD2.n47 49.446
R251 VDD2.n48 VDD2.n24 38.8791
R252 VDD2.n33 VDD2.n32 15.6631
R253 VDD2.n8 VDD2.n7 15.6631
R254 VDD2.n36 VDD2.n31 12.8005
R255 VDD2.n11 VDD2.n6 12.8005
R256 VDD2.n37 VDD2.n29 12.0247
R257 VDD2.n12 VDD2.n4 12.0247
R258 VDD2.n41 VDD2.n40 11.249
R259 VDD2.n16 VDD2.n15 11.249
R260 VDD2.n44 VDD2.n27 10.4732
R261 VDD2.n19 VDD2.n2 10.4732
R262 VDD2.n45 VDD2.n25 9.69747
R263 VDD2.n20 VDD2.n0 9.69747
R264 VDD2.n47 VDD2.n46 9.45567
R265 VDD2.n22 VDD2.n21 9.45567
R266 VDD2.n46 VDD2.n45 9.3005
R267 VDD2.n27 VDD2.n26 9.3005
R268 VDD2.n40 VDD2.n39 9.3005
R269 VDD2.n38 VDD2.n37 9.3005
R270 VDD2.n31 VDD2.n30 9.3005
R271 VDD2.n21 VDD2.n20 9.3005
R272 VDD2.n2 VDD2.n1 9.3005
R273 VDD2.n15 VDD2.n14 9.3005
R274 VDD2.n13 VDD2.n12 9.3005
R275 VDD2.n6 VDD2.n5 9.3005
R276 VDD2.n32 VDD2.n30 4.39059
R277 VDD2.n7 VDD2.n5 4.39059
R278 VDD2.n49 VDD2.t4 4.31423
R279 VDD2.n49 VDD2.t3 4.31423
R280 VDD2.n23 VDD2.t1 4.31423
R281 VDD2.n23 VDD2.t5 4.31423
R282 VDD2.n47 VDD2.n25 4.26717
R283 VDD2.n22 VDD2.n0 4.26717
R284 VDD2.n45 VDD2.n44 3.49141
R285 VDD2.n20 VDD2.n19 3.49141
R286 VDD2.n41 VDD2.n27 2.71565
R287 VDD2.n16 VDD2.n2 2.71565
R288 VDD2 VDD2.n48 2.6449
R289 VDD2.n40 VDD2.n29 1.93989
R290 VDD2.n15 VDD2.n4 1.93989
R291 VDD2.n37 VDD2.n36 1.16414
R292 VDD2.n12 VDD2.n11 1.16414
R293 VDD2.n33 VDD2.n31 0.388379
R294 VDD2.n8 VDD2.n6 0.388379
R295 VDD2.n46 VDD2.n26 0.155672
R296 VDD2.n39 VDD2.n26 0.155672
R297 VDD2.n39 VDD2.n38 0.155672
R298 VDD2.n38 VDD2.n30 0.155672
R299 VDD2.n13 VDD2.n5 0.155672
R300 VDD2.n14 VDD2.n13 0.155672
R301 VDD2.n14 VDD2.n1 0.155672
R302 VDD2.n21 VDD2.n1 0.155672
R303 B.n696 B.n695 585
R304 B.n697 B.n696 585
R305 B.n224 B.n126 585
R306 B.n223 B.n222 585
R307 B.n221 B.n220 585
R308 B.n219 B.n218 585
R309 B.n217 B.n216 585
R310 B.n215 B.n214 585
R311 B.n213 B.n212 585
R312 B.n211 B.n210 585
R313 B.n209 B.n208 585
R314 B.n207 B.n206 585
R315 B.n205 B.n204 585
R316 B.n203 B.n202 585
R317 B.n201 B.n200 585
R318 B.n199 B.n198 585
R319 B.n197 B.n196 585
R320 B.n195 B.n194 585
R321 B.n193 B.n192 585
R322 B.n191 B.n190 585
R323 B.n189 B.n188 585
R324 B.n186 B.n185 585
R325 B.n184 B.n183 585
R326 B.n182 B.n181 585
R327 B.n180 B.n179 585
R328 B.n178 B.n177 585
R329 B.n176 B.n175 585
R330 B.n174 B.n173 585
R331 B.n172 B.n171 585
R332 B.n170 B.n169 585
R333 B.n168 B.n167 585
R334 B.n166 B.n165 585
R335 B.n164 B.n163 585
R336 B.n162 B.n161 585
R337 B.n160 B.n159 585
R338 B.n158 B.n157 585
R339 B.n156 B.n155 585
R340 B.n154 B.n153 585
R341 B.n152 B.n151 585
R342 B.n150 B.n149 585
R343 B.n148 B.n147 585
R344 B.n146 B.n145 585
R345 B.n144 B.n143 585
R346 B.n142 B.n141 585
R347 B.n140 B.n139 585
R348 B.n138 B.n137 585
R349 B.n136 B.n135 585
R350 B.n134 B.n133 585
R351 B.n102 B.n101 585
R352 B.n700 B.n699 585
R353 B.n694 B.n127 585
R354 B.n127 B.n99 585
R355 B.n693 B.n98 585
R356 B.n704 B.n98 585
R357 B.n692 B.n97 585
R358 B.n705 B.n97 585
R359 B.n691 B.n96 585
R360 B.n706 B.n96 585
R361 B.n690 B.n689 585
R362 B.n689 B.n92 585
R363 B.n688 B.n91 585
R364 B.n712 B.n91 585
R365 B.n687 B.n90 585
R366 B.n713 B.n90 585
R367 B.n686 B.n89 585
R368 B.n714 B.n89 585
R369 B.n685 B.n684 585
R370 B.n684 B.n85 585
R371 B.n683 B.n84 585
R372 B.n720 B.n84 585
R373 B.n682 B.n83 585
R374 B.n721 B.n83 585
R375 B.n681 B.n82 585
R376 B.n722 B.n82 585
R377 B.n680 B.n679 585
R378 B.n679 B.n78 585
R379 B.n678 B.n77 585
R380 B.n728 B.n77 585
R381 B.n677 B.n76 585
R382 B.n729 B.n76 585
R383 B.n676 B.n75 585
R384 B.n730 B.n75 585
R385 B.n675 B.n674 585
R386 B.n674 B.n71 585
R387 B.n673 B.n70 585
R388 B.n736 B.n70 585
R389 B.n672 B.n69 585
R390 B.n737 B.n69 585
R391 B.n671 B.n68 585
R392 B.n738 B.n68 585
R393 B.n670 B.n669 585
R394 B.n669 B.n64 585
R395 B.n668 B.n63 585
R396 B.n744 B.n63 585
R397 B.n667 B.n62 585
R398 B.n745 B.n62 585
R399 B.n666 B.n61 585
R400 B.n746 B.n61 585
R401 B.n665 B.n664 585
R402 B.n664 B.n57 585
R403 B.n663 B.n56 585
R404 B.n752 B.n56 585
R405 B.n662 B.n55 585
R406 B.n753 B.n55 585
R407 B.n661 B.n54 585
R408 B.n754 B.n54 585
R409 B.n660 B.n659 585
R410 B.n659 B.n50 585
R411 B.n658 B.n49 585
R412 B.n760 B.n49 585
R413 B.n657 B.n48 585
R414 B.n761 B.n48 585
R415 B.n656 B.n47 585
R416 B.n762 B.n47 585
R417 B.n655 B.n654 585
R418 B.n654 B.n43 585
R419 B.n653 B.n42 585
R420 B.n768 B.n42 585
R421 B.n652 B.n41 585
R422 B.n769 B.n41 585
R423 B.n651 B.n40 585
R424 B.n770 B.n40 585
R425 B.n650 B.n649 585
R426 B.n649 B.n36 585
R427 B.n648 B.n35 585
R428 B.n776 B.n35 585
R429 B.n647 B.n34 585
R430 B.n777 B.n34 585
R431 B.n646 B.n33 585
R432 B.n778 B.n33 585
R433 B.n645 B.n644 585
R434 B.n644 B.n29 585
R435 B.n643 B.n28 585
R436 B.n784 B.n28 585
R437 B.n642 B.n27 585
R438 B.n785 B.n27 585
R439 B.n641 B.n26 585
R440 B.n786 B.n26 585
R441 B.n640 B.n639 585
R442 B.n639 B.n22 585
R443 B.n638 B.n21 585
R444 B.n792 B.n21 585
R445 B.n637 B.n20 585
R446 B.n793 B.n20 585
R447 B.n636 B.n19 585
R448 B.n794 B.n19 585
R449 B.n635 B.n634 585
R450 B.n634 B.n15 585
R451 B.n633 B.n14 585
R452 B.n800 B.n14 585
R453 B.n632 B.n13 585
R454 B.n801 B.n13 585
R455 B.n631 B.n12 585
R456 B.n802 B.n12 585
R457 B.n630 B.n629 585
R458 B.n629 B.n8 585
R459 B.n628 B.n7 585
R460 B.n808 B.n7 585
R461 B.n627 B.n6 585
R462 B.n809 B.n6 585
R463 B.n626 B.n5 585
R464 B.n810 B.n5 585
R465 B.n625 B.n624 585
R466 B.n624 B.n4 585
R467 B.n623 B.n225 585
R468 B.n623 B.n622 585
R469 B.n613 B.n226 585
R470 B.n227 B.n226 585
R471 B.n615 B.n614 585
R472 B.n616 B.n615 585
R473 B.n612 B.n232 585
R474 B.n232 B.n231 585
R475 B.n611 B.n610 585
R476 B.n610 B.n609 585
R477 B.n234 B.n233 585
R478 B.n235 B.n234 585
R479 B.n602 B.n601 585
R480 B.n603 B.n602 585
R481 B.n600 B.n240 585
R482 B.n240 B.n239 585
R483 B.n599 B.n598 585
R484 B.n598 B.n597 585
R485 B.n242 B.n241 585
R486 B.n243 B.n242 585
R487 B.n590 B.n589 585
R488 B.n591 B.n590 585
R489 B.n588 B.n248 585
R490 B.n248 B.n247 585
R491 B.n587 B.n586 585
R492 B.n586 B.n585 585
R493 B.n250 B.n249 585
R494 B.n251 B.n250 585
R495 B.n578 B.n577 585
R496 B.n579 B.n578 585
R497 B.n576 B.n256 585
R498 B.n256 B.n255 585
R499 B.n575 B.n574 585
R500 B.n574 B.n573 585
R501 B.n258 B.n257 585
R502 B.n259 B.n258 585
R503 B.n566 B.n565 585
R504 B.n567 B.n566 585
R505 B.n564 B.n264 585
R506 B.n264 B.n263 585
R507 B.n563 B.n562 585
R508 B.n562 B.n561 585
R509 B.n266 B.n265 585
R510 B.n267 B.n266 585
R511 B.n554 B.n553 585
R512 B.n555 B.n554 585
R513 B.n552 B.n272 585
R514 B.n272 B.n271 585
R515 B.n551 B.n550 585
R516 B.n550 B.n549 585
R517 B.n274 B.n273 585
R518 B.n275 B.n274 585
R519 B.n542 B.n541 585
R520 B.n543 B.n542 585
R521 B.n540 B.n280 585
R522 B.n280 B.n279 585
R523 B.n539 B.n538 585
R524 B.n538 B.n537 585
R525 B.n282 B.n281 585
R526 B.n283 B.n282 585
R527 B.n530 B.n529 585
R528 B.n531 B.n530 585
R529 B.n528 B.n288 585
R530 B.n288 B.n287 585
R531 B.n527 B.n526 585
R532 B.n526 B.n525 585
R533 B.n290 B.n289 585
R534 B.n291 B.n290 585
R535 B.n518 B.n517 585
R536 B.n519 B.n518 585
R537 B.n516 B.n296 585
R538 B.n296 B.n295 585
R539 B.n515 B.n514 585
R540 B.n514 B.n513 585
R541 B.n298 B.n297 585
R542 B.n299 B.n298 585
R543 B.n506 B.n505 585
R544 B.n507 B.n506 585
R545 B.n504 B.n304 585
R546 B.n304 B.n303 585
R547 B.n503 B.n502 585
R548 B.n502 B.n501 585
R549 B.n306 B.n305 585
R550 B.n307 B.n306 585
R551 B.n494 B.n493 585
R552 B.n495 B.n494 585
R553 B.n492 B.n312 585
R554 B.n312 B.n311 585
R555 B.n491 B.n490 585
R556 B.n490 B.n489 585
R557 B.n314 B.n313 585
R558 B.n315 B.n314 585
R559 B.n482 B.n481 585
R560 B.n483 B.n482 585
R561 B.n480 B.n320 585
R562 B.n320 B.n319 585
R563 B.n479 B.n478 585
R564 B.n478 B.n477 585
R565 B.n322 B.n321 585
R566 B.n323 B.n322 585
R567 B.n470 B.n469 585
R568 B.n471 B.n470 585
R569 B.n468 B.n328 585
R570 B.n328 B.n327 585
R571 B.n467 B.n466 585
R572 B.n466 B.n465 585
R573 B.n330 B.n329 585
R574 B.n331 B.n330 585
R575 B.n461 B.n460 585
R576 B.n334 B.n333 585
R577 B.n457 B.n456 585
R578 B.n458 B.n457 585
R579 B.n455 B.n358 585
R580 B.n454 B.n453 585
R581 B.n452 B.n451 585
R582 B.n450 B.n449 585
R583 B.n448 B.n447 585
R584 B.n446 B.n445 585
R585 B.n444 B.n443 585
R586 B.n442 B.n441 585
R587 B.n440 B.n439 585
R588 B.n438 B.n437 585
R589 B.n436 B.n435 585
R590 B.n434 B.n433 585
R591 B.n432 B.n431 585
R592 B.n430 B.n429 585
R593 B.n428 B.n427 585
R594 B.n426 B.n425 585
R595 B.n424 B.n423 585
R596 B.n421 B.n420 585
R597 B.n419 B.n418 585
R598 B.n417 B.n416 585
R599 B.n415 B.n414 585
R600 B.n413 B.n412 585
R601 B.n411 B.n410 585
R602 B.n409 B.n408 585
R603 B.n407 B.n406 585
R604 B.n405 B.n404 585
R605 B.n403 B.n402 585
R606 B.n401 B.n400 585
R607 B.n399 B.n398 585
R608 B.n397 B.n396 585
R609 B.n395 B.n394 585
R610 B.n393 B.n392 585
R611 B.n391 B.n390 585
R612 B.n389 B.n388 585
R613 B.n387 B.n386 585
R614 B.n385 B.n384 585
R615 B.n383 B.n382 585
R616 B.n381 B.n380 585
R617 B.n379 B.n378 585
R618 B.n377 B.n376 585
R619 B.n375 B.n374 585
R620 B.n373 B.n372 585
R621 B.n371 B.n370 585
R622 B.n369 B.n368 585
R623 B.n367 B.n366 585
R624 B.n365 B.n364 585
R625 B.n462 B.n332 585
R626 B.n332 B.n331 585
R627 B.n464 B.n463 585
R628 B.n465 B.n464 585
R629 B.n326 B.n325 585
R630 B.n327 B.n326 585
R631 B.n473 B.n472 585
R632 B.n472 B.n471 585
R633 B.n474 B.n324 585
R634 B.n324 B.n323 585
R635 B.n476 B.n475 585
R636 B.n477 B.n476 585
R637 B.n318 B.n317 585
R638 B.n319 B.n318 585
R639 B.n485 B.n484 585
R640 B.n484 B.n483 585
R641 B.n486 B.n316 585
R642 B.n316 B.n315 585
R643 B.n488 B.n487 585
R644 B.n489 B.n488 585
R645 B.n310 B.n309 585
R646 B.n311 B.n310 585
R647 B.n497 B.n496 585
R648 B.n496 B.n495 585
R649 B.n498 B.n308 585
R650 B.n308 B.n307 585
R651 B.n500 B.n499 585
R652 B.n501 B.n500 585
R653 B.n302 B.n301 585
R654 B.n303 B.n302 585
R655 B.n509 B.n508 585
R656 B.n508 B.n507 585
R657 B.n510 B.n300 585
R658 B.n300 B.n299 585
R659 B.n512 B.n511 585
R660 B.n513 B.n512 585
R661 B.n294 B.n293 585
R662 B.n295 B.n294 585
R663 B.n521 B.n520 585
R664 B.n520 B.n519 585
R665 B.n522 B.n292 585
R666 B.n292 B.n291 585
R667 B.n524 B.n523 585
R668 B.n525 B.n524 585
R669 B.n286 B.n285 585
R670 B.n287 B.n286 585
R671 B.n533 B.n532 585
R672 B.n532 B.n531 585
R673 B.n534 B.n284 585
R674 B.n284 B.n283 585
R675 B.n536 B.n535 585
R676 B.n537 B.n536 585
R677 B.n278 B.n277 585
R678 B.n279 B.n278 585
R679 B.n545 B.n544 585
R680 B.n544 B.n543 585
R681 B.n546 B.n276 585
R682 B.n276 B.n275 585
R683 B.n548 B.n547 585
R684 B.n549 B.n548 585
R685 B.n270 B.n269 585
R686 B.n271 B.n270 585
R687 B.n557 B.n556 585
R688 B.n556 B.n555 585
R689 B.n558 B.n268 585
R690 B.n268 B.n267 585
R691 B.n560 B.n559 585
R692 B.n561 B.n560 585
R693 B.n262 B.n261 585
R694 B.n263 B.n262 585
R695 B.n569 B.n568 585
R696 B.n568 B.n567 585
R697 B.n570 B.n260 585
R698 B.n260 B.n259 585
R699 B.n572 B.n571 585
R700 B.n573 B.n572 585
R701 B.n254 B.n253 585
R702 B.n255 B.n254 585
R703 B.n581 B.n580 585
R704 B.n580 B.n579 585
R705 B.n582 B.n252 585
R706 B.n252 B.n251 585
R707 B.n584 B.n583 585
R708 B.n585 B.n584 585
R709 B.n246 B.n245 585
R710 B.n247 B.n246 585
R711 B.n593 B.n592 585
R712 B.n592 B.n591 585
R713 B.n594 B.n244 585
R714 B.n244 B.n243 585
R715 B.n596 B.n595 585
R716 B.n597 B.n596 585
R717 B.n238 B.n237 585
R718 B.n239 B.n238 585
R719 B.n605 B.n604 585
R720 B.n604 B.n603 585
R721 B.n606 B.n236 585
R722 B.n236 B.n235 585
R723 B.n608 B.n607 585
R724 B.n609 B.n608 585
R725 B.n230 B.n229 585
R726 B.n231 B.n230 585
R727 B.n618 B.n617 585
R728 B.n617 B.n616 585
R729 B.n619 B.n228 585
R730 B.n228 B.n227 585
R731 B.n621 B.n620 585
R732 B.n622 B.n621 585
R733 B.n2 B.n0 585
R734 B.n4 B.n2 585
R735 B.n3 B.n1 585
R736 B.n809 B.n3 585
R737 B.n807 B.n806 585
R738 B.n808 B.n807 585
R739 B.n805 B.n9 585
R740 B.n9 B.n8 585
R741 B.n804 B.n803 585
R742 B.n803 B.n802 585
R743 B.n11 B.n10 585
R744 B.n801 B.n11 585
R745 B.n799 B.n798 585
R746 B.n800 B.n799 585
R747 B.n797 B.n16 585
R748 B.n16 B.n15 585
R749 B.n796 B.n795 585
R750 B.n795 B.n794 585
R751 B.n18 B.n17 585
R752 B.n793 B.n18 585
R753 B.n791 B.n790 585
R754 B.n792 B.n791 585
R755 B.n789 B.n23 585
R756 B.n23 B.n22 585
R757 B.n788 B.n787 585
R758 B.n787 B.n786 585
R759 B.n25 B.n24 585
R760 B.n785 B.n25 585
R761 B.n783 B.n782 585
R762 B.n784 B.n783 585
R763 B.n781 B.n30 585
R764 B.n30 B.n29 585
R765 B.n780 B.n779 585
R766 B.n779 B.n778 585
R767 B.n32 B.n31 585
R768 B.n777 B.n32 585
R769 B.n775 B.n774 585
R770 B.n776 B.n775 585
R771 B.n773 B.n37 585
R772 B.n37 B.n36 585
R773 B.n772 B.n771 585
R774 B.n771 B.n770 585
R775 B.n39 B.n38 585
R776 B.n769 B.n39 585
R777 B.n767 B.n766 585
R778 B.n768 B.n767 585
R779 B.n765 B.n44 585
R780 B.n44 B.n43 585
R781 B.n764 B.n763 585
R782 B.n763 B.n762 585
R783 B.n46 B.n45 585
R784 B.n761 B.n46 585
R785 B.n759 B.n758 585
R786 B.n760 B.n759 585
R787 B.n757 B.n51 585
R788 B.n51 B.n50 585
R789 B.n756 B.n755 585
R790 B.n755 B.n754 585
R791 B.n53 B.n52 585
R792 B.n753 B.n53 585
R793 B.n751 B.n750 585
R794 B.n752 B.n751 585
R795 B.n749 B.n58 585
R796 B.n58 B.n57 585
R797 B.n748 B.n747 585
R798 B.n747 B.n746 585
R799 B.n60 B.n59 585
R800 B.n745 B.n60 585
R801 B.n743 B.n742 585
R802 B.n744 B.n743 585
R803 B.n741 B.n65 585
R804 B.n65 B.n64 585
R805 B.n740 B.n739 585
R806 B.n739 B.n738 585
R807 B.n67 B.n66 585
R808 B.n737 B.n67 585
R809 B.n735 B.n734 585
R810 B.n736 B.n735 585
R811 B.n733 B.n72 585
R812 B.n72 B.n71 585
R813 B.n732 B.n731 585
R814 B.n731 B.n730 585
R815 B.n74 B.n73 585
R816 B.n729 B.n74 585
R817 B.n727 B.n726 585
R818 B.n728 B.n727 585
R819 B.n725 B.n79 585
R820 B.n79 B.n78 585
R821 B.n724 B.n723 585
R822 B.n723 B.n722 585
R823 B.n81 B.n80 585
R824 B.n721 B.n81 585
R825 B.n719 B.n718 585
R826 B.n720 B.n719 585
R827 B.n717 B.n86 585
R828 B.n86 B.n85 585
R829 B.n716 B.n715 585
R830 B.n715 B.n714 585
R831 B.n88 B.n87 585
R832 B.n713 B.n88 585
R833 B.n711 B.n710 585
R834 B.n712 B.n711 585
R835 B.n709 B.n93 585
R836 B.n93 B.n92 585
R837 B.n708 B.n707 585
R838 B.n707 B.n706 585
R839 B.n95 B.n94 585
R840 B.n705 B.n95 585
R841 B.n703 B.n702 585
R842 B.n704 B.n703 585
R843 B.n701 B.n100 585
R844 B.n100 B.n99 585
R845 B.n812 B.n811 585
R846 B.n811 B.n810 585
R847 B.n460 B.n332 545.355
R848 B.n699 B.n100 545.355
R849 B.n364 B.n330 545.355
R850 B.n696 B.n127 545.355
R851 B.n697 B.n125 256.663
R852 B.n697 B.n124 256.663
R853 B.n697 B.n123 256.663
R854 B.n697 B.n122 256.663
R855 B.n697 B.n121 256.663
R856 B.n697 B.n120 256.663
R857 B.n697 B.n119 256.663
R858 B.n697 B.n118 256.663
R859 B.n697 B.n117 256.663
R860 B.n697 B.n116 256.663
R861 B.n697 B.n115 256.663
R862 B.n697 B.n114 256.663
R863 B.n697 B.n113 256.663
R864 B.n697 B.n112 256.663
R865 B.n697 B.n111 256.663
R866 B.n697 B.n110 256.663
R867 B.n697 B.n109 256.663
R868 B.n697 B.n108 256.663
R869 B.n697 B.n107 256.663
R870 B.n697 B.n106 256.663
R871 B.n697 B.n105 256.663
R872 B.n697 B.n104 256.663
R873 B.n697 B.n103 256.663
R874 B.n698 B.n697 256.663
R875 B.n459 B.n458 256.663
R876 B.n458 B.n335 256.663
R877 B.n458 B.n336 256.663
R878 B.n458 B.n337 256.663
R879 B.n458 B.n338 256.663
R880 B.n458 B.n339 256.663
R881 B.n458 B.n340 256.663
R882 B.n458 B.n341 256.663
R883 B.n458 B.n342 256.663
R884 B.n458 B.n343 256.663
R885 B.n458 B.n344 256.663
R886 B.n458 B.n345 256.663
R887 B.n458 B.n346 256.663
R888 B.n458 B.n347 256.663
R889 B.n458 B.n348 256.663
R890 B.n458 B.n349 256.663
R891 B.n458 B.n350 256.663
R892 B.n458 B.n351 256.663
R893 B.n458 B.n352 256.663
R894 B.n458 B.n353 256.663
R895 B.n458 B.n354 256.663
R896 B.n458 B.n355 256.663
R897 B.n458 B.n356 256.663
R898 B.n458 B.n357 256.663
R899 B.n361 B.t10 239.381
R900 B.n359 B.t6 239.381
R901 B.n130 B.t17 239.381
R902 B.n128 B.t13 239.381
R903 B.n361 B.t12 232.412
R904 B.n128 B.t15 232.412
R905 B.n359 B.t9 232.412
R906 B.n130 B.t18 232.412
R907 B.n464 B.n332 163.367
R908 B.n464 B.n326 163.367
R909 B.n472 B.n326 163.367
R910 B.n472 B.n324 163.367
R911 B.n476 B.n324 163.367
R912 B.n476 B.n318 163.367
R913 B.n484 B.n318 163.367
R914 B.n484 B.n316 163.367
R915 B.n488 B.n316 163.367
R916 B.n488 B.n310 163.367
R917 B.n496 B.n310 163.367
R918 B.n496 B.n308 163.367
R919 B.n500 B.n308 163.367
R920 B.n500 B.n302 163.367
R921 B.n508 B.n302 163.367
R922 B.n508 B.n300 163.367
R923 B.n512 B.n300 163.367
R924 B.n512 B.n294 163.367
R925 B.n520 B.n294 163.367
R926 B.n520 B.n292 163.367
R927 B.n524 B.n292 163.367
R928 B.n524 B.n286 163.367
R929 B.n532 B.n286 163.367
R930 B.n532 B.n284 163.367
R931 B.n536 B.n284 163.367
R932 B.n536 B.n278 163.367
R933 B.n544 B.n278 163.367
R934 B.n544 B.n276 163.367
R935 B.n548 B.n276 163.367
R936 B.n548 B.n270 163.367
R937 B.n556 B.n270 163.367
R938 B.n556 B.n268 163.367
R939 B.n560 B.n268 163.367
R940 B.n560 B.n262 163.367
R941 B.n568 B.n262 163.367
R942 B.n568 B.n260 163.367
R943 B.n572 B.n260 163.367
R944 B.n572 B.n254 163.367
R945 B.n580 B.n254 163.367
R946 B.n580 B.n252 163.367
R947 B.n584 B.n252 163.367
R948 B.n584 B.n246 163.367
R949 B.n592 B.n246 163.367
R950 B.n592 B.n244 163.367
R951 B.n596 B.n244 163.367
R952 B.n596 B.n238 163.367
R953 B.n604 B.n238 163.367
R954 B.n604 B.n236 163.367
R955 B.n608 B.n236 163.367
R956 B.n608 B.n230 163.367
R957 B.n617 B.n230 163.367
R958 B.n617 B.n228 163.367
R959 B.n621 B.n228 163.367
R960 B.n621 B.n2 163.367
R961 B.n811 B.n2 163.367
R962 B.n811 B.n3 163.367
R963 B.n807 B.n3 163.367
R964 B.n807 B.n9 163.367
R965 B.n803 B.n9 163.367
R966 B.n803 B.n11 163.367
R967 B.n799 B.n11 163.367
R968 B.n799 B.n16 163.367
R969 B.n795 B.n16 163.367
R970 B.n795 B.n18 163.367
R971 B.n791 B.n18 163.367
R972 B.n791 B.n23 163.367
R973 B.n787 B.n23 163.367
R974 B.n787 B.n25 163.367
R975 B.n783 B.n25 163.367
R976 B.n783 B.n30 163.367
R977 B.n779 B.n30 163.367
R978 B.n779 B.n32 163.367
R979 B.n775 B.n32 163.367
R980 B.n775 B.n37 163.367
R981 B.n771 B.n37 163.367
R982 B.n771 B.n39 163.367
R983 B.n767 B.n39 163.367
R984 B.n767 B.n44 163.367
R985 B.n763 B.n44 163.367
R986 B.n763 B.n46 163.367
R987 B.n759 B.n46 163.367
R988 B.n759 B.n51 163.367
R989 B.n755 B.n51 163.367
R990 B.n755 B.n53 163.367
R991 B.n751 B.n53 163.367
R992 B.n751 B.n58 163.367
R993 B.n747 B.n58 163.367
R994 B.n747 B.n60 163.367
R995 B.n743 B.n60 163.367
R996 B.n743 B.n65 163.367
R997 B.n739 B.n65 163.367
R998 B.n739 B.n67 163.367
R999 B.n735 B.n67 163.367
R1000 B.n735 B.n72 163.367
R1001 B.n731 B.n72 163.367
R1002 B.n731 B.n74 163.367
R1003 B.n727 B.n74 163.367
R1004 B.n727 B.n79 163.367
R1005 B.n723 B.n79 163.367
R1006 B.n723 B.n81 163.367
R1007 B.n719 B.n81 163.367
R1008 B.n719 B.n86 163.367
R1009 B.n715 B.n86 163.367
R1010 B.n715 B.n88 163.367
R1011 B.n711 B.n88 163.367
R1012 B.n711 B.n93 163.367
R1013 B.n707 B.n93 163.367
R1014 B.n707 B.n95 163.367
R1015 B.n703 B.n95 163.367
R1016 B.n703 B.n100 163.367
R1017 B.n457 B.n334 163.367
R1018 B.n457 B.n358 163.367
R1019 B.n453 B.n452 163.367
R1020 B.n449 B.n448 163.367
R1021 B.n445 B.n444 163.367
R1022 B.n441 B.n440 163.367
R1023 B.n437 B.n436 163.367
R1024 B.n433 B.n432 163.367
R1025 B.n429 B.n428 163.367
R1026 B.n425 B.n424 163.367
R1027 B.n420 B.n419 163.367
R1028 B.n416 B.n415 163.367
R1029 B.n412 B.n411 163.367
R1030 B.n408 B.n407 163.367
R1031 B.n404 B.n403 163.367
R1032 B.n400 B.n399 163.367
R1033 B.n396 B.n395 163.367
R1034 B.n392 B.n391 163.367
R1035 B.n388 B.n387 163.367
R1036 B.n384 B.n383 163.367
R1037 B.n380 B.n379 163.367
R1038 B.n376 B.n375 163.367
R1039 B.n372 B.n371 163.367
R1040 B.n368 B.n367 163.367
R1041 B.n466 B.n330 163.367
R1042 B.n466 B.n328 163.367
R1043 B.n470 B.n328 163.367
R1044 B.n470 B.n322 163.367
R1045 B.n478 B.n322 163.367
R1046 B.n478 B.n320 163.367
R1047 B.n482 B.n320 163.367
R1048 B.n482 B.n314 163.367
R1049 B.n490 B.n314 163.367
R1050 B.n490 B.n312 163.367
R1051 B.n494 B.n312 163.367
R1052 B.n494 B.n306 163.367
R1053 B.n502 B.n306 163.367
R1054 B.n502 B.n304 163.367
R1055 B.n506 B.n304 163.367
R1056 B.n506 B.n298 163.367
R1057 B.n514 B.n298 163.367
R1058 B.n514 B.n296 163.367
R1059 B.n518 B.n296 163.367
R1060 B.n518 B.n290 163.367
R1061 B.n526 B.n290 163.367
R1062 B.n526 B.n288 163.367
R1063 B.n530 B.n288 163.367
R1064 B.n530 B.n282 163.367
R1065 B.n538 B.n282 163.367
R1066 B.n538 B.n280 163.367
R1067 B.n542 B.n280 163.367
R1068 B.n542 B.n274 163.367
R1069 B.n550 B.n274 163.367
R1070 B.n550 B.n272 163.367
R1071 B.n554 B.n272 163.367
R1072 B.n554 B.n266 163.367
R1073 B.n562 B.n266 163.367
R1074 B.n562 B.n264 163.367
R1075 B.n566 B.n264 163.367
R1076 B.n566 B.n258 163.367
R1077 B.n574 B.n258 163.367
R1078 B.n574 B.n256 163.367
R1079 B.n578 B.n256 163.367
R1080 B.n578 B.n250 163.367
R1081 B.n586 B.n250 163.367
R1082 B.n586 B.n248 163.367
R1083 B.n590 B.n248 163.367
R1084 B.n590 B.n242 163.367
R1085 B.n598 B.n242 163.367
R1086 B.n598 B.n240 163.367
R1087 B.n602 B.n240 163.367
R1088 B.n602 B.n234 163.367
R1089 B.n610 B.n234 163.367
R1090 B.n610 B.n232 163.367
R1091 B.n615 B.n232 163.367
R1092 B.n615 B.n226 163.367
R1093 B.n623 B.n226 163.367
R1094 B.n624 B.n623 163.367
R1095 B.n624 B.n5 163.367
R1096 B.n6 B.n5 163.367
R1097 B.n7 B.n6 163.367
R1098 B.n629 B.n7 163.367
R1099 B.n629 B.n12 163.367
R1100 B.n13 B.n12 163.367
R1101 B.n14 B.n13 163.367
R1102 B.n634 B.n14 163.367
R1103 B.n634 B.n19 163.367
R1104 B.n20 B.n19 163.367
R1105 B.n21 B.n20 163.367
R1106 B.n639 B.n21 163.367
R1107 B.n639 B.n26 163.367
R1108 B.n27 B.n26 163.367
R1109 B.n28 B.n27 163.367
R1110 B.n644 B.n28 163.367
R1111 B.n644 B.n33 163.367
R1112 B.n34 B.n33 163.367
R1113 B.n35 B.n34 163.367
R1114 B.n649 B.n35 163.367
R1115 B.n649 B.n40 163.367
R1116 B.n41 B.n40 163.367
R1117 B.n42 B.n41 163.367
R1118 B.n654 B.n42 163.367
R1119 B.n654 B.n47 163.367
R1120 B.n48 B.n47 163.367
R1121 B.n49 B.n48 163.367
R1122 B.n659 B.n49 163.367
R1123 B.n659 B.n54 163.367
R1124 B.n55 B.n54 163.367
R1125 B.n56 B.n55 163.367
R1126 B.n664 B.n56 163.367
R1127 B.n664 B.n61 163.367
R1128 B.n62 B.n61 163.367
R1129 B.n63 B.n62 163.367
R1130 B.n669 B.n63 163.367
R1131 B.n669 B.n68 163.367
R1132 B.n69 B.n68 163.367
R1133 B.n70 B.n69 163.367
R1134 B.n674 B.n70 163.367
R1135 B.n674 B.n75 163.367
R1136 B.n76 B.n75 163.367
R1137 B.n77 B.n76 163.367
R1138 B.n679 B.n77 163.367
R1139 B.n679 B.n82 163.367
R1140 B.n83 B.n82 163.367
R1141 B.n84 B.n83 163.367
R1142 B.n684 B.n84 163.367
R1143 B.n684 B.n89 163.367
R1144 B.n90 B.n89 163.367
R1145 B.n91 B.n90 163.367
R1146 B.n689 B.n91 163.367
R1147 B.n689 B.n96 163.367
R1148 B.n97 B.n96 163.367
R1149 B.n98 B.n97 163.367
R1150 B.n127 B.n98 163.367
R1151 B.n133 B.n102 163.367
R1152 B.n137 B.n136 163.367
R1153 B.n141 B.n140 163.367
R1154 B.n145 B.n144 163.367
R1155 B.n149 B.n148 163.367
R1156 B.n153 B.n152 163.367
R1157 B.n157 B.n156 163.367
R1158 B.n161 B.n160 163.367
R1159 B.n165 B.n164 163.367
R1160 B.n169 B.n168 163.367
R1161 B.n173 B.n172 163.367
R1162 B.n177 B.n176 163.367
R1163 B.n181 B.n180 163.367
R1164 B.n185 B.n184 163.367
R1165 B.n190 B.n189 163.367
R1166 B.n194 B.n193 163.367
R1167 B.n198 B.n197 163.367
R1168 B.n202 B.n201 163.367
R1169 B.n206 B.n205 163.367
R1170 B.n210 B.n209 163.367
R1171 B.n214 B.n213 163.367
R1172 B.n218 B.n217 163.367
R1173 B.n222 B.n221 163.367
R1174 B.n696 B.n126 163.367
R1175 B.n362 B.t11 154.837
R1176 B.n129 B.t16 154.837
R1177 B.n360 B.t8 154.837
R1178 B.n131 B.t19 154.837
R1179 B.n458 B.n331 150.532
R1180 B.n697 B.n99 150.532
R1181 B.n362 B.n361 77.5763
R1182 B.n360 B.n359 77.5763
R1183 B.n131 B.n130 77.5763
R1184 B.n129 B.n128 77.5763
R1185 B.n465 B.n331 75.8241
R1186 B.n465 B.n327 75.8241
R1187 B.n471 B.n327 75.8241
R1188 B.n471 B.n323 75.8241
R1189 B.n477 B.n323 75.8241
R1190 B.n477 B.n319 75.8241
R1191 B.n483 B.n319 75.8241
R1192 B.n483 B.n315 75.8241
R1193 B.n489 B.n315 75.8241
R1194 B.n495 B.n311 75.8241
R1195 B.n495 B.n307 75.8241
R1196 B.n501 B.n307 75.8241
R1197 B.n501 B.n303 75.8241
R1198 B.n507 B.n303 75.8241
R1199 B.n507 B.n299 75.8241
R1200 B.n513 B.n299 75.8241
R1201 B.n513 B.n295 75.8241
R1202 B.n519 B.n295 75.8241
R1203 B.n519 B.n291 75.8241
R1204 B.n525 B.n291 75.8241
R1205 B.n525 B.n287 75.8241
R1206 B.n531 B.n287 75.8241
R1207 B.n537 B.n283 75.8241
R1208 B.n537 B.n279 75.8241
R1209 B.n543 B.n279 75.8241
R1210 B.n543 B.n275 75.8241
R1211 B.n549 B.n275 75.8241
R1212 B.n549 B.n271 75.8241
R1213 B.n555 B.n271 75.8241
R1214 B.n555 B.n267 75.8241
R1215 B.n561 B.n267 75.8241
R1216 B.n561 B.n263 75.8241
R1217 B.n567 B.n263 75.8241
R1218 B.n573 B.n259 75.8241
R1219 B.n573 B.n255 75.8241
R1220 B.n579 B.n255 75.8241
R1221 B.n579 B.n251 75.8241
R1222 B.n585 B.n251 75.8241
R1223 B.n585 B.n247 75.8241
R1224 B.n591 B.n247 75.8241
R1225 B.n591 B.n243 75.8241
R1226 B.n597 B.n243 75.8241
R1227 B.n597 B.n239 75.8241
R1228 B.n603 B.n239 75.8241
R1229 B.n609 B.n235 75.8241
R1230 B.n609 B.n231 75.8241
R1231 B.n616 B.n231 75.8241
R1232 B.n616 B.n227 75.8241
R1233 B.n622 B.n227 75.8241
R1234 B.n622 B.n4 75.8241
R1235 B.n810 B.n4 75.8241
R1236 B.n810 B.n809 75.8241
R1237 B.n809 B.n808 75.8241
R1238 B.n808 B.n8 75.8241
R1239 B.n802 B.n8 75.8241
R1240 B.n802 B.n801 75.8241
R1241 B.n801 B.n800 75.8241
R1242 B.n800 B.n15 75.8241
R1243 B.n794 B.n793 75.8241
R1244 B.n793 B.n792 75.8241
R1245 B.n792 B.n22 75.8241
R1246 B.n786 B.n22 75.8241
R1247 B.n786 B.n785 75.8241
R1248 B.n785 B.n784 75.8241
R1249 B.n784 B.n29 75.8241
R1250 B.n778 B.n29 75.8241
R1251 B.n778 B.n777 75.8241
R1252 B.n777 B.n776 75.8241
R1253 B.n776 B.n36 75.8241
R1254 B.n770 B.n769 75.8241
R1255 B.n769 B.n768 75.8241
R1256 B.n768 B.n43 75.8241
R1257 B.n762 B.n43 75.8241
R1258 B.n762 B.n761 75.8241
R1259 B.n761 B.n760 75.8241
R1260 B.n760 B.n50 75.8241
R1261 B.n754 B.n50 75.8241
R1262 B.n754 B.n753 75.8241
R1263 B.n753 B.n752 75.8241
R1264 B.n752 B.n57 75.8241
R1265 B.n746 B.n745 75.8241
R1266 B.n745 B.n744 75.8241
R1267 B.n744 B.n64 75.8241
R1268 B.n738 B.n64 75.8241
R1269 B.n738 B.n737 75.8241
R1270 B.n737 B.n736 75.8241
R1271 B.n736 B.n71 75.8241
R1272 B.n730 B.n71 75.8241
R1273 B.n730 B.n729 75.8241
R1274 B.n729 B.n728 75.8241
R1275 B.n728 B.n78 75.8241
R1276 B.n722 B.n78 75.8241
R1277 B.n722 B.n721 75.8241
R1278 B.n720 B.n85 75.8241
R1279 B.n714 B.n85 75.8241
R1280 B.n714 B.n713 75.8241
R1281 B.n713 B.n712 75.8241
R1282 B.n712 B.n92 75.8241
R1283 B.n706 B.n92 75.8241
R1284 B.n706 B.n705 75.8241
R1285 B.n705 B.n704 75.8241
R1286 B.n704 B.n99 75.8241
R1287 B.t7 B.n311 74.7091
R1288 B.n531 B.t4 74.7091
R1289 B.n746 B.t2 74.7091
R1290 B.n721 B.t14 74.7091
R1291 B.n460 B.n459 71.676
R1292 B.n358 B.n335 71.676
R1293 B.n452 B.n336 71.676
R1294 B.n448 B.n337 71.676
R1295 B.n444 B.n338 71.676
R1296 B.n440 B.n339 71.676
R1297 B.n436 B.n340 71.676
R1298 B.n432 B.n341 71.676
R1299 B.n428 B.n342 71.676
R1300 B.n424 B.n343 71.676
R1301 B.n419 B.n344 71.676
R1302 B.n415 B.n345 71.676
R1303 B.n411 B.n346 71.676
R1304 B.n407 B.n347 71.676
R1305 B.n403 B.n348 71.676
R1306 B.n399 B.n349 71.676
R1307 B.n395 B.n350 71.676
R1308 B.n391 B.n351 71.676
R1309 B.n387 B.n352 71.676
R1310 B.n383 B.n353 71.676
R1311 B.n379 B.n354 71.676
R1312 B.n375 B.n355 71.676
R1313 B.n371 B.n356 71.676
R1314 B.n367 B.n357 71.676
R1315 B.n699 B.n698 71.676
R1316 B.n133 B.n103 71.676
R1317 B.n137 B.n104 71.676
R1318 B.n141 B.n105 71.676
R1319 B.n145 B.n106 71.676
R1320 B.n149 B.n107 71.676
R1321 B.n153 B.n108 71.676
R1322 B.n157 B.n109 71.676
R1323 B.n161 B.n110 71.676
R1324 B.n165 B.n111 71.676
R1325 B.n169 B.n112 71.676
R1326 B.n173 B.n113 71.676
R1327 B.n177 B.n114 71.676
R1328 B.n181 B.n115 71.676
R1329 B.n185 B.n116 71.676
R1330 B.n190 B.n117 71.676
R1331 B.n194 B.n118 71.676
R1332 B.n198 B.n119 71.676
R1333 B.n202 B.n120 71.676
R1334 B.n206 B.n121 71.676
R1335 B.n210 B.n122 71.676
R1336 B.n214 B.n123 71.676
R1337 B.n218 B.n124 71.676
R1338 B.n222 B.n125 71.676
R1339 B.n126 B.n125 71.676
R1340 B.n221 B.n124 71.676
R1341 B.n217 B.n123 71.676
R1342 B.n213 B.n122 71.676
R1343 B.n209 B.n121 71.676
R1344 B.n205 B.n120 71.676
R1345 B.n201 B.n119 71.676
R1346 B.n197 B.n118 71.676
R1347 B.n193 B.n117 71.676
R1348 B.n189 B.n116 71.676
R1349 B.n184 B.n115 71.676
R1350 B.n180 B.n114 71.676
R1351 B.n176 B.n113 71.676
R1352 B.n172 B.n112 71.676
R1353 B.n168 B.n111 71.676
R1354 B.n164 B.n110 71.676
R1355 B.n160 B.n109 71.676
R1356 B.n156 B.n108 71.676
R1357 B.n152 B.n107 71.676
R1358 B.n148 B.n106 71.676
R1359 B.n144 B.n105 71.676
R1360 B.n140 B.n104 71.676
R1361 B.n136 B.n103 71.676
R1362 B.n698 B.n102 71.676
R1363 B.n459 B.n334 71.676
R1364 B.n453 B.n335 71.676
R1365 B.n449 B.n336 71.676
R1366 B.n445 B.n337 71.676
R1367 B.n441 B.n338 71.676
R1368 B.n437 B.n339 71.676
R1369 B.n433 B.n340 71.676
R1370 B.n429 B.n341 71.676
R1371 B.n425 B.n342 71.676
R1372 B.n420 B.n343 71.676
R1373 B.n416 B.n344 71.676
R1374 B.n412 B.n345 71.676
R1375 B.n408 B.n346 71.676
R1376 B.n404 B.n347 71.676
R1377 B.n400 B.n348 71.676
R1378 B.n396 B.n349 71.676
R1379 B.n392 B.n350 71.676
R1380 B.n388 B.n351 71.676
R1381 B.n384 B.n352 71.676
R1382 B.n380 B.n353 71.676
R1383 B.n376 B.n354 71.676
R1384 B.n372 B.n355 71.676
R1385 B.n368 B.n356 71.676
R1386 B.n364 B.n357 71.676
R1387 B.n363 B.n362 59.5399
R1388 B.n422 B.n360 59.5399
R1389 B.n132 B.n131 59.5399
R1390 B.n187 B.n129 59.5399
R1391 B.n567 B.t5 56.8682
R1392 B.n770 B.t1 56.8682
R1393 B.n603 B.t3 39.0274
R1394 B.n794 B.t0 39.0274
R1395 B.t3 B.n235 36.7973
R1396 B.t0 B.n15 36.7973
R1397 B.n695 B.n694 35.4346
R1398 B.n701 B.n700 35.4346
R1399 B.n365 B.n329 35.4346
R1400 B.n462 B.n461 35.4346
R1401 B.t5 B.n259 18.9564
R1402 B.t1 B.n36 18.9564
R1403 B B.n812 18.0485
R1404 B.n700 B.n101 10.6151
R1405 B.n134 B.n101 10.6151
R1406 B.n135 B.n134 10.6151
R1407 B.n138 B.n135 10.6151
R1408 B.n139 B.n138 10.6151
R1409 B.n142 B.n139 10.6151
R1410 B.n143 B.n142 10.6151
R1411 B.n146 B.n143 10.6151
R1412 B.n147 B.n146 10.6151
R1413 B.n150 B.n147 10.6151
R1414 B.n151 B.n150 10.6151
R1415 B.n154 B.n151 10.6151
R1416 B.n155 B.n154 10.6151
R1417 B.n158 B.n155 10.6151
R1418 B.n159 B.n158 10.6151
R1419 B.n162 B.n159 10.6151
R1420 B.n163 B.n162 10.6151
R1421 B.n166 B.n163 10.6151
R1422 B.n167 B.n166 10.6151
R1423 B.n171 B.n170 10.6151
R1424 B.n174 B.n171 10.6151
R1425 B.n175 B.n174 10.6151
R1426 B.n178 B.n175 10.6151
R1427 B.n179 B.n178 10.6151
R1428 B.n182 B.n179 10.6151
R1429 B.n183 B.n182 10.6151
R1430 B.n186 B.n183 10.6151
R1431 B.n191 B.n188 10.6151
R1432 B.n192 B.n191 10.6151
R1433 B.n195 B.n192 10.6151
R1434 B.n196 B.n195 10.6151
R1435 B.n199 B.n196 10.6151
R1436 B.n200 B.n199 10.6151
R1437 B.n203 B.n200 10.6151
R1438 B.n204 B.n203 10.6151
R1439 B.n207 B.n204 10.6151
R1440 B.n208 B.n207 10.6151
R1441 B.n211 B.n208 10.6151
R1442 B.n212 B.n211 10.6151
R1443 B.n215 B.n212 10.6151
R1444 B.n216 B.n215 10.6151
R1445 B.n219 B.n216 10.6151
R1446 B.n220 B.n219 10.6151
R1447 B.n223 B.n220 10.6151
R1448 B.n224 B.n223 10.6151
R1449 B.n695 B.n224 10.6151
R1450 B.n467 B.n329 10.6151
R1451 B.n468 B.n467 10.6151
R1452 B.n469 B.n468 10.6151
R1453 B.n469 B.n321 10.6151
R1454 B.n479 B.n321 10.6151
R1455 B.n480 B.n479 10.6151
R1456 B.n481 B.n480 10.6151
R1457 B.n481 B.n313 10.6151
R1458 B.n491 B.n313 10.6151
R1459 B.n492 B.n491 10.6151
R1460 B.n493 B.n492 10.6151
R1461 B.n493 B.n305 10.6151
R1462 B.n503 B.n305 10.6151
R1463 B.n504 B.n503 10.6151
R1464 B.n505 B.n504 10.6151
R1465 B.n505 B.n297 10.6151
R1466 B.n515 B.n297 10.6151
R1467 B.n516 B.n515 10.6151
R1468 B.n517 B.n516 10.6151
R1469 B.n517 B.n289 10.6151
R1470 B.n527 B.n289 10.6151
R1471 B.n528 B.n527 10.6151
R1472 B.n529 B.n528 10.6151
R1473 B.n529 B.n281 10.6151
R1474 B.n539 B.n281 10.6151
R1475 B.n540 B.n539 10.6151
R1476 B.n541 B.n540 10.6151
R1477 B.n541 B.n273 10.6151
R1478 B.n551 B.n273 10.6151
R1479 B.n552 B.n551 10.6151
R1480 B.n553 B.n552 10.6151
R1481 B.n553 B.n265 10.6151
R1482 B.n563 B.n265 10.6151
R1483 B.n564 B.n563 10.6151
R1484 B.n565 B.n564 10.6151
R1485 B.n565 B.n257 10.6151
R1486 B.n575 B.n257 10.6151
R1487 B.n576 B.n575 10.6151
R1488 B.n577 B.n576 10.6151
R1489 B.n577 B.n249 10.6151
R1490 B.n587 B.n249 10.6151
R1491 B.n588 B.n587 10.6151
R1492 B.n589 B.n588 10.6151
R1493 B.n589 B.n241 10.6151
R1494 B.n599 B.n241 10.6151
R1495 B.n600 B.n599 10.6151
R1496 B.n601 B.n600 10.6151
R1497 B.n601 B.n233 10.6151
R1498 B.n611 B.n233 10.6151
R1499 B.n612 B.n611 10.6151
R1500 B.n614 B.n612 10.6151
R1501 B.n614 B.n613 10.6151
R1502 B.n613 B.n225 10.6151
R1503 B.n625 B.n225 10.6151
R1504 B.n626 B.n625 10.6151
R1505 B.n627 B.n626 10.6151
R1506 B.n628 B.n627 10.6151
R1507 B.n630 B.n628 10.6151
R1508 B.n631 B.n630 10.6151
R1509 B.n632 B.n631 10.6151
R1510 B.n633 B.n632 10.6151
R1511 B.n635 B.n633 10.6151
R1512 B.n636 B.n635 10.6151
R1513 B.n637 B.n636 10.6151
R1514 B.n638 B.n637 10.6151
R1515 B.n640 B.n638 10.6151
R1516 B.n641 B.n640 10.6151
R1517 B.n642 B.n641 10.6151
R1518 B.n643 B.n642 10.6151
R1519 B.n645 B.n643 10.6151
R1520 B.n646 B.n645 10.6151
R1521 B.n647 B.n646 10.6151
R1522 B.n648 B.n647 10.6151
R1523 B.n650 B.n648 10.6151
R1524 B.n651 B.n650 10.6151
R1525 B.n652 B.n651 10.6151
R1526 B.n653 B.n652 10.6151
R1527 B.n655 B.n653 10.6151
R1528 B.n656 B.n655 10.6151
R1529 B.n657 B.n656 10.6151
R1530 B.n658 B.n657 10.6151
R1531 B.n660 B.n658 10.6151
R1532 B.n661 B.n660 10.6151
R1533 B.n662 B.n661 10.6151
R1534 B.n663 B.n662 10.6151
R1535 B.n665 B.n663 10.6151
R1536 B.n666 B.n665 10.6151
R1537 B.n667 B.n666 10.6151
R1538 B.n668 B.n667 10.6151
R1539 B.n670 B.n668 10.6151
R1540 B.n671 B.n670 10.6151
R1541 B.n672 B.n671 10.6151
R1542 B.n673 B.n672 10.6151
R1543 B.n675 B.n673 10.6151
R1544 B.n676 B.n675 10.6151
R1545 B.n677 B.n676 10.6151
R1546 B.n678 B.n677 10.6151
R1547 B.n680 B.n678 10.6151
R1548 B.n681 B.n680 10.6151
R1549 B.n682 B.n681 10.6151
R1550 B.n683 B.n682 10.6151
R1551 B.n685 B.n683 10.6151
R1552 B.n686 B.n685 10.6151
R1553 B.n687 B.n686 10.6151
R1554 B.n688 B.n687 10.6151
R1555 B.n690 B.n688 10.6151
R1556 B.n691 B.n690 10.6151
R1557 B.n692 B.n691 10.6151
R1558 B.n693 B.n692 10.6151
R1559 B.n694 B.n693 10.6151
R1560 B.n461 B.n333 10.6151
R1561 B.n456 B.n333 10.6151
R1562 B.n456 B.n455 10.6151
R1563 B.n455 B.n454 10.6151
R1564 B.n454 B.n451 10.6151
R1565 B.n451 B.n450 10.6151
R1566 B.n450 B.n447 10.6151
R1567 B.n447 B.n446 10.6151
R1568 B.n446 B.n443 10.6151
R1569 B.n443 B.n442 10.6151
R1570 B.n442 B.n439 10.6151
R1571 B.n439 B.n438 10.6151
R1572 B.n438 B.n435 10.6151
R1573 B.n435 B.n434 10.6151
R1574 B.n434 B.n431 10.6151
R1575 B.n431 B.n430 10.6151
R1576 B.n430 B.n427 10.6151
R1577 B.n427 B.n426 10.6151
R1578 B.n426 B.n423 10.6151
R1579 B.n421 B.n418 10.6151
R1580 B.n418 B.n417 10.6151
R1581 B.n417 B.n414 10.6151
R1582 B.n414 B.n413 10.6151
R1583 B.n413 B.n410 10.6151
R1584 B.n410 B.n409 10.6151
R1585 B.n409 B.n406 10.6151
R1586 B.n406 B.n405 10.6151
R1587 B.n402 B.n401 10.6151
R1588 B.n401 B.n398 10.6151
R1589 B.n398 B.n397 10.6151
R1590 B.n397 B.n394 10.6151
R1591 B.n394 B.n393 10.6151
R1592 B.n393 B.n390 10.6151
R1593 B.n390 B.n389 10.6151
R1594 B.n389 B.n386 10.6151
R1595 B.n386 B.n385 10.6151
R1596 B.n385 B.n382 10.6151
R1597 B.n382 B.n381 10.6151
R1598 B.n381 B.n378 10.6151
R1599 B.n378 B.n377 10.6151
R1600 B.n377 B.n374 10.6151
R1601 B.n374 B.n373 10.6151
R1602 B.n373 B.n370 10.6151
R1603 B.n370 B.n369 10.6151
R1604 B.n369 B.n366 10.6151
R1605 B.n366 B.n365 10.6151
R1606 B.n463 B.n462 10.6151
R1607 B.n463 B.n325 10.6151
R1608 B.n473 B.n325 10.6151
R1609 B.n474 B.n473 10.6151
R1610 B.n475 B.n474 10.6151
R1611 B.n475 B.n317 10.6151
R1612 B.n485 B.n317 10.6151
R1613 B.n486 B.n485 10.6151
R1614 B.n487 B.n486 10.6151
R1615 B.n487 B.n309 10.6151
R1616 B.n497 B.n309 10.6151
R1617 B.n498 B.n497 10.6151
R1618 B.n499 B.n498 10.6151
R1619 B.n499 B.n301 10.6151
R1620 B.n509 B.n301 10.6151
R1621 B.n510 B.n509 10.6151
R1622 B.n511 B.n510 10.6151
R1623 B.n511 B.n293 10.6151
R1624 B.n521 B.n293 10.6151
R1625 B.n522 B.n521 10.6151
R1626 B.n523 B.n522 10.6151
R1627 B.n523 B.n285 10.6151
R1628 B.n533 B.n285 10.6151
R1629 B.n534 B.n533 10.6151
R1630 B.n535 B.n534 10.6151
R1631 B.n535 B.n277 10.6151
R1632 B.n545 B.n277 10.6151
R1633 B.n546 B.n545 10.6151
R1634 B.n547 B.n546 10.6151
R1635 B.n547 B.n269 10.6151
R1636 B.n557 B.n269 10.6151
R1637 B.n558 B.n557 10.6151
R1638 B.n559 B.n558 10.6151
R1639 B.n559 B.n261 10.6151
R1640 B.n569 B.n261 10.6151
R1641 B.n570 B.n569 10.6151
R1642 B.n571 B.n570 10.6151
R1643 B.n571 B.n253 10.6151
R1644 B.n581 B.n253 10.6151
R1645 B.n582 B.n581 10.6151
R1646 B.n583 B.n582 10.6151
R1647 B.n583 B.n245 10.6151
R1648 B.n593 B.n245 10.6151
R1649 B.n594 B.n593 10.6151
R1650 B.n595 B.n594 10.6151
R1651 B.n595 B.n237 10.6151
R1652 B.n605 B.n237 10.6151
R1653 B.n606 B.n605 10.6151
R1654 B.n607 B.n606 10.6151
R1655 B.n607 B.n229 10.6151
R1656 B.n618 B.n229 10.6151
R1657 B.n619 B.n618 10.6151
R1658 B.n620 B.n619 10.6151
R1659 B.n620 B.n0 10.6151
R1660 B.n806 B.n1 10.6151
R1661 B.n806 B.n805 10.6151
R1662 B.n805 B.n804 10.6151
R1663 B.n804 B.n10 10.6151
R1664 B.n798 B.n10 10.6151
R1665 B.n798 B.n797 10.6151
R1666 B.n797 B.n796 10.6151
R1667 B.n796 B.n17 10.6151
R1668 B.n790 B.n17 10.6151
R1669 B.n790 B.n789 10.6151
R1670 B.n789 B.n788 10.6151
R1671 B.n788 B.n24 10.6151
R1672 B.n782 B.n24 10.6151
R1673 B.n782 B.n781 10.6151
R1674 B.n781 B.n780 10.6151
R1675 B.n780 B.n31 10.6151
R1676 B.n774 B.n31 10.6151
R1677 B.n774 B.n773 10.6151
R1678 B.n773 B.n772 10.6151
R1679 B.n772 B.n38 10.6151
R1680 B.n766 B.n38 10.6151
R1681 B.n766 B.n765 10.6151
R1682 B.n765 B.n764 10.6151
R1683 B.n764 B.n45 10.6151
R1684 B.n758 B.n45 10.6151
R1685 B.n758 B.n757 10.6151
R1686 B.n757 B.n756 10.6151
R1687 B.n756 B.n52 10.6151
R1688 B.n750 B.n52 10.6151
R1689 B.n750 B.n749 10.6151
R1690 B.n749 B.n748 10.6151
R1691 B.n748 B.n59 10.6151
R1692 B.n742 B.n59 10.6151
R1693 B.n742 B.n741 10.6151
R1694 B.n741 B.n740 10.6151
R1695 B.n740 B.n66 10.6151
R1696 B.n734 B.n66 10.6151
R1697 B.n734 B.n733 10.6151
R1698 B.n733 B.n732 10.6151
R1699 B.n732 B.n73 10.6151
R1700 B.n726 B.n73 10.6151
R1701 B.n726 B.n725 10.6151
R1702 B.n725 B.n724 10.6151
R1703 B.n724 B.n80 10.6151
R1704 B.n718 B.n80 10.6151
R1705 B.n718 B.n717 10.6151
R1706 B.n717 B.n716 10.6151
R1707 B.n716 B.n87 10.6151
R1708 B.n710 B.n87 10.6151
R1709 B.n710 B.n709 10.6151
R1710 B.n709 B.n708 10.6151
R1711 B.n708 B.n94 10.6151
R1712 B.n702 B.n94 10.6151
R1713 B.n702 B.n701 10.6151
R1714 B.n170 B.n132 6.5566
R1715 B.n187 B.n186 6.5566
R1716 B.n422 B.n421 6.5566
R1717 B.n405 B.n363 6.5566
R1718 B.n167 B.n132 4.05904
R1719 B.n188 B.n187 4.05904
R1720 B.n423 B.n422 4.05904
R1721 B.n402 B.n363 4.05904
R1722 B.n812 B.n0 2.81026
R1723 B.n812 B.n1 2.81026
R1724 B.n489 B.t7 1.11555
R1725 B.t4 B.n283 1.11555
R1726 B.t2 B.n57 1.11555
R1727 B.t14 B.n720 1.11555
R1728 VP.n14 VP.n11 161.3
R1729 VP.n16 VP.n15 161.3
R1730 VP.n17 VP.n10 161.3
R1731 VP.n19 VP.n18 161.3
R1732 VP.n20 VP.n9 161.3
R1733 VP.n22 VP.n21 161.3
R1734 VP.n23 VP.n8 161.3
R1735 VP.n49 VP.n0 161.3
R1736 VP.n48 VP.n47 161.3
R1737 VP.n46 VP.n1 161.3
R1738 VP.n45 VP.n44 161.3
R1739 VP.n43 VP.n2 161.3
R1740 VP.n42 VP.n41 161.3
R1741 VP.n40 VP.n3 161.3
R1742 VP.n39 VP.n38 161.3
R1743 VP.n37 VP.n4 161.3
R1744 VP.n36 VP.n35 161.3
R1745 VP.n34 VP.n5 161.3
R1746 VP.n33 VP.n32 161.3
R1747 VP.n31 VP.n6 161.3
R1748 VP.n30 VP.n29 161.3
R1749 VP.n28 VP.n7 161.3
R1750 VP.n13 VP.t3 62.2513
R1751 VP.n27 VP.n26 57.7148
R1752 VP.n51 VP.n50 57.7148
R1753 VP.n25 VP.n24 57.7148
R1754 VP.n13 VP.n12 50.4779
R1755 VP.n27 VP.n25 47.4888
R1756 VP.n32 VP.n31 40.4934
R1757 VP.n32 VP.n5 40.4934
R1758 VP.n44 VP.n43 40.4934
R1759 VP.n44 VP.n1 40.4934
R1760 VP.n18 VP.n9 40.4934
R1761 VP.n18 VP.n17 40.4934
R1762 VP.n50 VP.t5 30.1419
R1763 VP.n38 VP.t0 30.1419
R1764 VP.n26 VP.t2 30.1419
R1765 VP.n12 VP.t4 30.1419
R1766 VP.n24 VP.t1 30.1419
R1767 VP.n26 VP.n7 24.4675
R1768 VP.n30 VP.n7 24.4675
R1769 VP.n31 VP.n30 24.4675
R1770 VP.n36 VP.n5 24.4675
R1771 VP.n37 VP.n36 24.4675
R1772 VP.n38 VP.n37 24.4675
R1773 VP.n38 VP.n3 24.4675
R1774 VP.n42 VP.n3 24.4675
R1775 VP.n43 VP.n42 24.4675
R1776 VP.n48 VP.n1 24.4675
R1777 VP.n49 VP.n48 24.4675
R1778 VP.n50 VP.n49 24.4675
R1779 VP.n22 VP.n9 24.4675
R1780 VP.n23 VP.n22 24.4675
R1781 VP.n24 VP.n23 24.4675
R1782 VP.n12 VP.n11 24.4675
R1783 VP.n16 VP.n11 24.4675
R1784 VP.n17 VP.n16 24.4675
R1785 VP.n14 VP.n13 2.52647
R1786 VP.n25 VP.n8 0.417535
R1787 VP.n28 VP.n27 0.417535
R1788 VP.n51 VP.n0 0.417535
R1789 VP VP.n51 0.394291
R1790 VP.n15 VP.n14 0.189894
R1791 VP.n15 VP.n10 0.189894
R1792 VP.n19 VP.n10 0.189894
R1793 VP.n20 VP.n19 0.189894
R1794 VP.n21 VP.n20 0.189894
R1795 VP.n21 VP.n8 0.189894
R1796 VP.n29 VP.n28 0.189894
R1797 VP.n29 VP.n6 0.189894
R1798 VP.n33 VP.n6 0.189894
R1799 VP.n34 VP.n33 0.189894
R1800 VP.n35 VP.n34 0.189894
R1801 VP.n35 VP.n4 0.189894
R1802 VP.n39 VP.n4 0.189894
R1803 VP.n40 VP.n39 0.189894
R1804 VP.n41 VP.n40 0.189894
R1805 VP.n41 VP.n2 0.189894
R1806 VP.n45 VP.n2 0.189894
R1807 VP.n46 VP.n45 0.189894
R1808 VP.n47 VP.n46 0.189894
R1809 VP.n47 VP.n0 0.189894
R1810 VDD1.n18 VDD1.n0 289.615
R1811 VDD1.n41 VDD1.n23 289.615
R1812 VDD1.n19 VDD1.n18 185
R1813 VDD1.n17 VDD1.n16 185
R1814 VDD1.n4 VDD1.n3 185
R1815 VDD1.n11 VDD1.n10 185
R1816 VDD1.n9 VDD1.n8 185
R1817 VDD1.n32 VDD1.n31 185
R1818 VDD1.n34 VDD1.n33 185
R1819 VDD1.n27 VDD1.n26 185
R1820 VDD1.n40 VDD1.n39 185
R1821 VDD1.n42 VDD1.n41 185
R1822 VDD1.n7 VDD1.t2 147.714
R1823 VDD1.n30 VDD1.t3 147.714
R1824 VDD1.n18 VDD1.n17 104.615
R1825 VDD1.n17 VDD1.n3 104.615
R1826 VDD1.n10 VDD1.n3 104.615
R1827 VDD1.n10 VDD1.n9 104.615
R1828 VDD1.n33 VDD1.n32 104.615
R1829 VDD1.n33 VDD1.n26 104.615
R1830 VDD1.n40 VDD1.n26 104.615
R1831 VDD1.n41 VDD1.n40 104.615
R1832 VDD1.n47 VDD1.n46 72.0302
R1833 VDD1.n49 VDD1.n48 71.2235
R1834 VDD1.n9 VDD1.t2 52.3082
R1835 VDD1.n32 VDD1.t3 52.3082
R1836 VDD1 VDD1.n22 52.0904
R1837 VDD1.n47 VDD1.n45 51.9768
R1838 VDD1.n49 VDD1.n47 41.1862
R1839 VDD1.n8 VDD1.n7 15.6631
R1840 VDD1.n31 VDD1.n30 15.6631
R1841 VDD1.n11 VDD1.n6 12.8005
R1842 VDD1.n34 VDD1.n29 12.8005
R1843 VDD1.n12 VDD1.n4 12.0247
R1844 VDD1.n35 VDD1.n27 12.0247
R1845 VDD1.n16 VDD1.n15 11.249
R1846 VDD1.n39 VDD1.n38 11.249
R1847 VDD1.n19 VDD1.n2 10.4732
R1848 VDD1.n42 VDD1.n25 10.4732
R1849 VDD1.n20 VDD1.n0 9.69747
R1850 VDD1.n43 VDD1.n23 9.69747
R1851 VDD1.n22 VDD1.n21 9.45567
R1852 VDD1.n45 VDD1.n44 9.45567
R1853 VDD1.n21 VDD1.n20 9.3005
R1854 VDD1.n2 VDD1.n1 9.3005
R1855 VDD1.n15 VDD1.n14 9.3005
R1856 VDD1.n13 VDD1.n12 9.3005
R1857 VDD1.n6 VDD1.n5 9.3005
R1858 VDD1.n44 VDD1.n43 9.3005
R1859 VDD1.n25 VDD1.n24 9.3005
R1860 VDD1.n38 VDD1.n37 9.3005
R1861 VDD1.n36 VDD1.n35 9.3005
R1862 VDD1.n29 VDD1.n28 9.3005
R1863 VDD1.n7 VDD1.n5 4.39059
R1864 VDD1.n30 VDD1.n28 4.39059
R1865 VDD1.n48 VDD1.t1 4.31423
R1866 VDD1.n48 VDD1.t4 4.31423
R1867 VDD1.n46 VDD1.t5 4.31423
R1868 VDD1.n46 VDD1.t0 4.31423
R1869 VDD1.n22 VDD1.n0 4.26717
R1870 VDD1.n45 VDD1.n23 4.26717
R1871 VDD1.n20 VDD1.n19 3.49141
R1872 VDD1.n43 VDD1.n42 3.49141
R1873 VDD1.n16 VDD1.n2 2.71565
R1874 VDD1.n39 VDD1.n25 2.71565
R1875 VDD1.n15 VDD1.n4 1.93989
R1876 VDD1.n38 VDD1.n27 1.93989
R1877 VDD1.n12 VDD1.n11 1.16414
R1878 VDD1.n35 VDD1.n34 1.16414
R1879 VDD1 VDD1.n49 0.804379
R1880 VDD1.n8 VDD1.n6 0.388379
R1881 VDD1.n31 VDD1.n29 0.388379
R1882 VDD1.n21 VDD1.n1 0.155672
R1883 VDD1.n14 VDD1.n1 0.155672
R1884 VDD1.n14 VDD1.n13 0.155672
R1885 VDD1.n13 VDD1.n5 0.155672
R1886 VDD1.n36 VDD1.n28 0.155672
R1887 VDD1.n37 VDD1.n36 0.155672
R1888 VDD1.n37 VDD1.n24 0.155672
R1889 VDD1.n44 VDD1.n24 0.155672
C0 VTAIL VN 3.96481f
C1 VN VDD1 0.155969f
C2 VDD2 VN 2.97749f
C3 VP VN 6.60451f
C4 VTAIL VDD1 5.71547f
C5 VDD2 VTAIL 5.77556f
C6 VP VTAIL 3.97905f
C7 VDD2 VDD1 1.82247f
C8 VP VDD1 3.37171f
C9 VP VDD2 0.552815f
C10 VDD2 B 5.48705f
C11 VDD1 B 5.667533f
C12 VTAIL B 5.037504f
C13 VN B 15.392489f
C14 VP B 14.035734f
C15 VDD1.n0 B 0.03125f
C16 VDD1.n1 B 0.022779f
C17 VDD1.n2 B 0.012241f
C18 VDD1.n3 B 0.028932f
C19 VDD1.n4 B 0.012961f
C20 VDD1.n5 B 0.393675f
C21 VDD1.n6 B 0.012241f
C22 VDD1.t2 B 0.047452f
C23 VDD1.n7 B 0.090172f
C24 VDD1.n8 B 0.017074f
C25 VDD1.n9 B 0.021699f
C26 VDD1.n10 B 0.028932f
C27 VDD1.n11 B 0.012961f
C28 VDD1.n12 B 0.012241f
C29 VDD1.n13 B 0.022779f
C30 VDD1.n14 B 0.022779f
C31 VDD1.n15 B 0.012241f
C32 VDD1.n16 B 0.012961f
C33 VDD1.n17 B 0.028932f
C34 VDD1.n18 B 0.061275f
C35 VDD1.n19 B 0.012961f
C36 VDD1.n20 B 0.012241f
C37 VDD1.n21 B 0.053587f
C38 VDD1.n22 B 0.062003f
C39 VDD1.n23 B 0.03125f
C40 VDD1.n24 B 0.022779f
C41 VDD1.n25 B 0.012241f
C42 VDD1.n26 B 0.028932f
C43 VDD1.n27 B 0.012961f
C44 VDD1.n28 B 0.393675f
C45 VDD1.n29 B 0.012241f
C46 VDD1.t3 B 0.047452f
C47 VDD1.n30 B 0.090172f
C48 VDD1.n31 B 0.017074f
C49 VDD1.n32 B 0.021699f
C50 VDD1.n33 B 0.028932f
C51 VDD1.n34 B 0.012961f
C52 VDD1.n35 B 0.012241f
C53 VDD1.n36 B 0.022779f
C54 VDD1.n37 B 0.022779f
C55 VDD1.n38 B 0.012241f
C56 VDD1.n39 B 0.012961f
C57 VDD1.n40 B 0.028932f
C58 VDD1.n41 B 0.061275f
C59 VDD1.n42 B 0.012961f
C60 VDD1.n43 B 0.012241f
C61 VDD1.n44 B 0.053587f
C62 VDD1.n45 B 0.061113f
C63 VDD1.t5 B 0.082624f
C64 VDD1.t0 B 0.082624f
C65 VDD1.n46 B 0.67f
C66 VDD1.n47 B 2.57442f
C67 VDD1.t1 B 0.082624f
C68 VDD1.t4 B 0.082624f
C69 VDD1.n48 B 0.664379f
C70 VDD1.n49 B 2.28936f
C71 VP.n0 B 0.045084f
C72 VP.t5 B 1.04933f
C73 VP.n1 B 0.047637f
C74 VP.n2 B 0.023968f
C75 VP.n3 B 0.044671f
C76 VP.n4 B 0.023968f
C77 VP.t0 B 1.04933f
C78 VP.n5 B 0.047637f
C79 VP.n6 B 0.023968f
C80 VP.n7 B 0.044671f
C81 VP.n8 B 0.045084f
C82 VP.t1 B 1.04933f
C83 VP.n9 B 0.047637f
C84 VP.n10 B 0.023968f
C85 VP.n11 B 0.044671f
C86 VP.t3 B 1.35191f
C87 VP.t4 B 1.04933f
C88 VP.n12 B 0.49705f
C89 VP.n13 B 0.487552f
C90 VP.n14 B 0.305437f
C91 VP.n15 B 0.023968f
C92 VP.n16 B 0.044671f
C93 VP.n17 B 0.047637f
C94 VP.n18 B 0.019376f
C95 VP.n19 B 0.023968f
C96 VP.n20 B 0.023968f
C97 VP.n21 B 0.023968f
C98 VP.n22 B 0.044671f
C99 VP.n23 B 0.044671f
C100 VP.n24 B 0.505427f
C101 VP.n25 B 1.28663f
C102 VP.t2 B 1.04933f
C103 VP.n26 B 0.505427f
C104 VP.n27 B 1.30477f
C105 VP.n28 B 0.045084f
C106 VP.n29 B 0.023968f
C107 VP.n30 B 0.044671f
C108 VP.n31 B 0.047637f
C109 VP.n32 B 0.019376f
C110 VP.n33 B 0.023968f
C111 VP.n34 B 0.023968f
C112 VP.n35 B 0.023968f
C113 VP.n36 B 0.044671f
C114 VP.n37 B 0.044671f
C115 VP.n38 B 0.421839f
C116 VP.n39 B 0.023968f
C117 VP.n40 B 0.023968f
C118 VP.n41 B 0.023968f
C119 VP.n42 B 0.044671f
C120 VP.n43 B 0.047637f
C121 VP.n44 B 0.019376f
C122 VP.n45 B 0.023968f
C123 VP.n46 B 0.023968f
C124 VP.n47 B 0.023968f
C125 VP.n48 B 0.044671f
C126 VP.n49 B 0.044671f
C127 VP.n50 B 0.505427f
C128 VP.n51 B 0.067458f
C129 VDD2.n0 B 0.030502f
C130 VDD2.n1 B 0.022234f
C131 VDD2.n2 B 0.011948f
C132 VDD2.n3 B 0.02824f
C133 VDD2.n4 B 0.01265f
C134 VDD2.n5 B 0.38425f
C135 VDD2.n6 B 0.011948f
C136 VDD2.t2 B 0.046316f
C137 VDD2.n7 B 0.088013f
C138 VDD2.n8 B 0.016666f
C139 VDD2.n9 B 0.02118f
C140 VDD2.n10 B 0.02824f
C141 VDD2.n11 B 0.01265f
C142 VDD2.n12 B 0.011948f
C143 VDD2.n13 B 0.022234f
C144 VDD2.n14 B 0.022234f
C145 VDD2.n15 B 0.011948f
C146 VDD2.n16 B 0.01265f
C147 VDD2.n17 B 0.02824f
C148 VDD2.n18 B 0.059808f
C149 VDD2.n19 B 0.01265f
C150 VDD2.n20 B 0.011948f
C151 VDD2.n21 B 0.052304f
C152 VDD2.n22 B 0.05965f
C153 VDD2.t1 B 0.080646f
C154 VDD2.t5 B 0.080646f
C155 VDD2.n23 B 0.653958f
C156 VDD2.n24 B 2.38456f
C157 VDD2.n25 B 0.030502f
C158 VDD2.n26 B 0.022234f
C159 VDD2.n27 B 0.011948f
C160 VDD2.n28 B 0.02824f
C161 VDD2.n29 B 0.01265f
C162 VDD2.n30 B 0.38425f
C163 VDD2.n31 B 0.011948f
C164 VDD2.t0 B 0.046316f
C165 VDD2.n32 B 0.088013f
C166 VDD2.n33 B 0.016666f
C167 VDD2.n34 B 0.02118f
C168 VDD2.n35 B 0.02824f
C169 VDD2.n36 B 0.01265f
C170 VDD2.n37 B 0.011948f
C171 VDD2.n38 B 0.022234f
C172 VDD2.n39 B 0.022234f
C173 VDD2.n40 B 0.011948f
C174 VDD2.n41 B 0.01265f
C175 VDD2.n42 B 0.02824f
C176 VDD2.n43 B 0.059808f
C177 VDD2.n44 B 0.01265f
C178 VDD2.n45 B 0.011948f
C179 VDD2.n46 B 0.052304f
C180 VDD2.n47 B 0.048701f
C181 VDD2.n48 B 2.02438f
C182 VDD2.t4 B 0.080646f
C183 VDD2.t3 B 0.080646f
C184 VDD2.n49 B 0.65393f
C185 VTAIL.t6 B 0.109941f
C186 VTAIL.t9 B 0.109941f
C187 VTAIL.n0 B 0.812653f
C188 VTAIL.n1 B 0.573538f
C189 VTAIL.n2 B 0.041582f
C190 VTAIL.n3 B 0.03031f
C191 VTAIL.n4 B 0.016288f
C192 VTAIL.n5 B 0.038498f
C193 VTAIL.n6 B 0.017246f
C194 VTAIL.n7 B 0.52383f
C195 VTAIL.n8 B 0.016288f
C196 VTAIL.t3 B 0.063141f
C197 VTAIL.n9 B 0.119983f
C198 VTAIL.n10 B 0.022719f
C199 VTAIL.n11 B 0.028873f
C200 VTAIL.n12 B 0.038498f
C201 VTAIL.n13 B 0.017246f
C202 VTAIL.n14 B 0.016288f
C203 VTAIL.n15 B 0.03031f
C204 VTAIL.n16 B 0.03031f
C205 VTAIL.n17 B 0.016288f
C206 VTAIL.n18 B 0.017246f
C207 VTAIL.n19 B 0.038498f
C208 VTAIL.n20 B 0.081533f
C209 VTAIL.n21 B 0.017246f
C210 VTAIL.n22 B 0.016288f
C211 VTAIL.n23 B 0.071304f
C212 VTAIL.n24 B 0.045473f
C213 VTAIL.n25 B 0.577651f
C214 VTAIL.t4 B 0.109941f
C215 VTAIL.t5 B 0.109941f
C216 VTAIL.n26 B 0.812653f
C217 VTAIL.n27 B 2.07792f
C218 VTAIL.t8 B 0.109941f
C219 VTAIL.t7 B 0.109941f
C220 VTAIL.n28 B 0.812658f
C221 VTAIL.n29 B 2.07792f
C222 VTAIL.n30 B 0.041582f
C223 VTAIL.n31 B 0.03031f
C224 VTAIL.n32 B 0.016288f
C225 VTAIL.n33 B 0.038498f
C226 VTAIL.n34 B 0.017246f
C227 VTAIL.n35 B 0.52383f
C228 VTAIL.n36 B 0.016288f
C229 VTAIL.t11 B 0.063141f
C230 VTAIL.n37 B 0.119983f
C231 VTAIL.n38 B 0.022719f
C232 VTAIL.n39 B 0.028873f
C233 VTAIL.n40 B 0.038498f
C234 VTAIL.n41 B 0.017246f
C235 VTAIL.n42 B 0.016288f
C236 VTAIL.n43 B 0.03031f
C237 VTAIL.n44 B 0.03031f
C238 VTAIL.n45 B 0.016288f
C239 VTAIL.n46 B 0.017246f
C240 VTAIL.n47 B 0.038498f
C241 VTAIL.n48 B 0.081533f
C242 VTAIL.n49 B 0.017246f
C243 VTAIL.n50 B 0.016288f
C244 VTAIL.n51 B 0.071304f
C245 VTAIL.n52 B 0.045473f
C246 VTAIL.n53 B 0.577651f
C247 VTAIL.t0 B 0.109941f
C248 VTAIL.t1 B 0.109941f
C249 VTAIL.n54 B 0.812658f
C250 VTAIL.n55 B 0.820437f
C251 VTAIL.n56 B 0.041582f
C252 VTAIL.n57 B 0.03031f
C253 VTAIL.n58 B 0.016288f
C254 VTAIL.n59 B 0.038498f
C255 VTAIL.n60 B 0.017246f
C256 VTAIL.n61 B 0.52383f
C257 VTAIL.n62 B 0.016288f
C258 VTAIL.t2 B 0.063141f
C259 VTAIL.n63 B 0.119983f
C260 VTAIL.n64 B 0.022719f
C261 VTAIL.n65 B 0.028873f
C262 VTAIL.n66 B 0.038498f
C263 VTAIL.n67 B 0.017246f
C264 VTAIL.n68 B 0.016288f
C265 VTAIL.n69 B 0.03031f
C266 VTAIL.n70 B 0.03031f
C267 VTAIL.n71 B 0.016288f
C268 VTAIL.n72 B 0.017246f
C269 VTAIL.n73 B 0.038498f
C270 VTAIL.n74 B 0.081533f
C271 VTAIL.n75 B 0.017246f
C272 VTAIL.n76 B 0.016288f
C273 VTAIL.n77 B 0.071304f
C274 VTAIL.n78 B 0.045473f
C275 VTAIL.n79 B 1.49835f
C276 VTAIL.n80 B 0.041582f
C277 VTAIL.n81 B 0.03031f
C278 VTAIL.n82 B 0.016288f
C279 VTAIL.n83 B 0.038498f
C280 VTAIL.n84 B 0.017246f
C281 VTAIL.n85 B 0.52383f
C282 VTAIL.n86 B 0.016288f
C283 VTAIL.t10 B 0.063141f
C284 VTAIL.n87 B 0.119983f
C285 VTAIL.n88 B 0.022719f
C286 VTAIL.n89 B 0.028873f
C287 VTAIL.n90 B 0.038498f
C288 VTAIL.n91 B 0.017246f
C289 VTAIL.n92 B 0.016288f
C290 VTAIL.n93 B 0.03031f
C291 VTAIL.n94 B 0.03031f
C292 VTAIL.n95 B 0.016288f
C293 VTAIL.n96 B 0.017246f
C294 VTAIL.n97 B 0.038498f
C295 VTAIL.n98 B 0.081533f
C296 VTAIL.n99 B 0.017246f
C297 VTAIL.n100 B 0.016288f
C298 VTAIL.n101 B 0.071304f
C299 VTAIL.n102 B 0.045473f
C300 VTAIL.n103 B 1.40847f
C301 VN.n0 B 0.043691f
C302 VN.t0 B 1.0169f
C303 VN.n1 B 0.046165f
C304 VN.n2 B 0.023228f
C305 VN.n3 B 0.04329f
C306 VN.t3 B 1.31014f
C307 VN.t4 B 1.0169f
C308 VN.n4 B 0.481689f
C309 VN.n5 B 0.472483f
C310 VN.n6 B 0.295997f
C311 VN.n7 B 0.023228f
C312 VN.n8 B 0.04329f
C313 VN.n9 B 0.046165f
C314 VN.n10 B 0.018777f
C315 VN.n11 B 0.023228f
C316 VN.n12 B 0.023228f
C317 VN.n13 B 0.023228f
C318 VN.n14 B 0.04329f
C319 VN.n15 B 0.04329f
C320 VN.n16 B 0.489807f
C321 VN.n17 B 0.065373f
C322 VN.n18 B 0.043691f
C323 VN.t5 B 1.0169f
C324 VN.n19 B 0.046165f
C325 VN.n20 B 0.023228f
C326 VN.n21 B 0.04329f
C327 VN.t2 B 1.31014f
C328 VN.t1 B 1.0169f
C329 VN.n22 B 0.481689f
C330 VN.n23 B 0.472483f
C331 VN.n24 B 0.295997f
C332 VN.n25 B 0.023228f
C333 VN.n26 B 0.04329f
C334 VN.n27 B 0.046165f
C335 VN.n28 B 0.018777f
C336 VN.n29 B 0.023228f
C337 VN.n30 B 0.023228f
C338 VN.n31 B 0.023228f
C339 VN.n32 B 0.04329f
C340 VN.n33 B 0.04329f
C341 VN.n34 B 0.489807f
C342 VN.n35 B 1.2532f
.ends

