* NGSPICE file created from diff_pair_sample_1406.ext - technology: sky130A

.subckt diff_pair_sample_1406 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=0.58
X1 VTAIL.t5 VP.t1 VDD1.t2 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=0.58
X2 B.t11 B.t9 B.t10 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=0.58
X3 VDD2.t3 VN.t0 VTAIL.t1 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=0.58
X4 VDD2.t2 VN.t1 VTAIL.t2 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=0.58
X5 B.t8 B.t6 B.t7 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=0.58
X6 B.t5 B.t3 B.t4 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=0.58
X7 VTAIL.t0 VN.t2 VDD2.t1 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=0.58
X8 VDD1.t1 VP.t2 VTAIL.t4 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=0.58
X9 VTAIL.t7 VP.t3 VDD1.t0 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=0.58
X10 VTAIL.t3 VN.t3 VDD2.t0 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=0.58
X11 B.t2 B.t0 B.t1 w_n1516_n1466# sky130_fd_pr__pfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=0.58
R0 VP.n0 VP.t3 192.59
R1 VP.n0 VP.t0 192.566
R2 VP.n2 VP.t1 171.609
R3 VP.n3 VP.t2 171.609
R4 VP.n4 VP.n3 161.3
R5 VP.n2 VP.n1 161.3
R6 VP.n1 VP.n0 103.153
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n90 VTAIL.n84 756.745
R11 VTAIL.n6 VTAIL.n0 756.745
R12 VTAIL.n18 VTAIL.n12 756.745
R13 VTAIL.n30 VTAIL.n24 756.745
R14 VTAIL.n78 VTAIL.n72 756.745
R15 VTAIL.n66 VTAIL.n60 756.745
R16 VTAIL.n54 VTAIL.n48 756.745
R17 VTAIL.n42 VTAIL.n36 756.745
R18 VTAIL.n89 VTAIL.n88 585
R19 VTAIL.n91 VTAIL.n90 585
R20 VTAIL.n5 VTAIL.n4 585
R21 VTAIL.n7 VTAIL.n6 585
R22 VTAIL.n17 VTAIL.n16 585
R23 VTAIL.n19 VTAIL.n18 585
R24 VTAIL.n29 VTAIL.n28 585
R25 VTAIL.n31 VTAIL.n30 585
R26 VTAIL.n79 VTAIL.n78 585
R27 VTAIL.n77 VTAIL.n76 585
R28 VTAIL.n67 VTAIL.n66 585
R29 VTAIL.n65 VTAIL.n64 585
R30 VTAIL.n55 VTAIL.n54 585
R31 VTAIL.n53 VTAIL.n52 585
R32 VTAIL.n43 VTAIL.n42 585
R33 VTAIL.n41 VTAIL.n40 585
R34 VTAIL.n87 VTAIL.t2 355.474
R35 VTAIL.n3 VTAIL.t3 355.474
R36 VTAIL.n15 VTAIL.t4 355.474
R37 VTAIL.n27 VTAIL.t5 355.474
R38 VTAIL.n75 VTAIL.t6 355.474
R39 VTAIL.n63 VTAIL.t7 355.474
R40 VTAIL.n51 VTAIL.t1 355.474
R41 VTAIL.n39 VTAIL.t0 355.474
R42 VTAIL.n90 VTAIL.n89 171.744
R43 VTAIL.n6 VTAIL.n5 171.744
R44 VTAIL.n18 VTAIL.n17 171.744
R45 VTAIL.n30 VTAIL.n29 171.744
R46 VTAIL.n78 VTAIL.n77 171.744
R47 VTAIL.n66 VTAIL.n65 171.744
R48 VTAIL.n54 VTAIL.n53 171.744
R49 VTAIL.n42 VTAIL.n41 171.744
R50 VTAIL.n89 VTAIL.t2 85.8723
R51 VTAIL.n5 VTAIL.t3 85.8723
R52 VTAIL.n17 VTAIL.t4 85.8723
R53 VTAIL.n29 VTAIL.t5 85.8723
R54 VTAIL.n77 VTAIL.t6 85.8723
R55 VTAIL.n65 VTAIL.t7 85.8723
R56 VTAIL.n53 VTAIL.t1 85.8723
R57 VTAIL.n41 VTAIL.t0 85.8723
R58 VTAIL.n95 VTAIL.n94 33.9308
R59 VTAIL.n11 VTAIL.n10 33.9308
R60 VTAIL.n23 VTAIL.n22 33.9308
R61 VTAIL.n35 VTAIL.n34 33.9308
R62 VTAIL.n83 VTAIL.n82 33.9308
R63 VTAIL.n71 VTAIL.n70 33.9308
R64 VTAIL.n59 VTAIL.n58 33.9308
R65 VTAIL.n47 VTAIL.n46 33.9308
R66 VTAIL.n88 VTAIL.n87 15.8418
R67 VTAIL.n4 VTAIL.n3 15.8418
R68 VTAIL.n16 VTAIL.n15 15.8418
R69 VTAIL.n28 VTAIL.n27 15.8418
R70 VTAIL.n76 VTAIL.n75 15.8418
R71 VTAIL.n64 VTAIL.n63 15.8418
R72 VTAIL.n52 VTAIL.n51 15.8418
R73 VTAIL.n40 VTAIL.n39 15.8418
R74 VTAIL.n95 VTAIL.n83 15.2979
R75 VTAIL.n47 VTAIL.n35 15.2979
R76 VTAIL.n91 VTAIL.n86 12.8005
R77 VTAIL.n7 VTAIL.n2 12.8005
R78 VTAIL.n19 VTAIL.n14 12.8005
R79 VTAIL.n31 VTAIL.n26 12.8005
R80 VTAIL.n79 VTAIL.n74 12.8005
R81 VTAIL.n67 VTAIL.n62 12.8005
R82 VTAIL.n55 VTAIL.n50 12.8005
R83 VTAIL.n43 VTAIL.n38 12.8005
R84 VTAIL.n92 VTAIL.n84 12.0247
R85 VTAIL.n8 VTAIL.n0 12.0247
R86 VTAIL.n20 VTAIL.n12 12.0247
R87 VTAIL.n32 VTAIL.n24 12.0247
R88 VTAIL.n80 VTAIL.n72 12.0247
R89 VTAIL.n68 VTAIL.n60 12.0247
R90 VTAIL.n56 VTAIL.n48 12.0247
R91 VTAIL.n44 VTAIL.n36 12.0247
R92 VTAIL.n94 VTAIL.n93 9.45567
R93 VTAIL.n10 VTAIL.n9 9.45567
R94 VTAIL.n22 VTAIL.n21 9.45567
R95 VTAIL.n34 VTAIL.n33 9.45567
R96 VTAIL.n82 VTAIL.n81 9.45567
R97 VTAIL.n70 VTAIL.n69 9.45567
R98 VTAIL.n58 VTAIL.n57 9.45567
R99 VTAIL.n46 VTAIL.n45 9.45567
R100 VTAIL.n93 VTAIL.n92 9.3005
R101 VTAIL.n86 VTAIL.n85 9.3005
R102 VTAIL.n9 VTAIL.n8 9.3005
R103 VTAIL.n2 VTAIL.n1 9.3005
R104 VTAIL.n21 VTAIL.n20 9.3005
R105 VTAIL.n14 VTAIL.n13 9.3005
R106 VTAIL.n33 VTAIL.n32 9.3005
R107 VTAIL.n26 VTAIL.n25 9.3005
R108 VTAIL.n81 VTAIL.n80 9.3005
R109 VTAIL.n74 VTAIL.n73 9.3005
R110 VTAIL.n69 VTAIL.n68 9.3005
R111 VTAIL.n62 VTAIL.n61 9.3005
R112 VTAIL.n57 VTAIL.n56 9.3005
R113 VTAIL.n50 VTAIL.n49 9.3005
R114 VTAIL.n45 VTAIL.n44 9.3005
R115 VTAIL.n38 VTAIL.n37 9.3005
R116 VTAIL.n75 VTAIL.n73 4.29255
R117 VTAIL.n63 VTAIL.n61 4.29255
R118 VTAIL.n51 VTAIL.n49 4.29255
R119 VTAIL.n39 VTAIL.n37 4.29255
R120 VTAIL.n87 VTAIL.n85 4.29255
R121 VTAIL.n3 VTAIL.n1 4.29255
R122 VTAIL.n15 VTAIL.n13 4.29255
R123 VTAIL.n27 VTAIL.n25 4.29255
R124 VTAIL.n94 VTAIL.n84 1.93989
R125 VTAIL.n10 VTAIL.n0 1.93989
R126 VTAIL.n22 VTAIL.n12 1.93989
R127 VTAIL.n34 VTAIL.n24 1.93989
R128 VTAIL.n82 VTAIL.n72 1.93989
R129 VTAIL.n70 VTAIL.n60 1.93989
R130 VTAIL.n58 VTAIL.n48 1.93989
R131 VTAIL.n46 VTAIL.n36 1.93989
R132 VTAIL.n92 VTAIL.n91 1.16414
R133 VTAIL.n8 VTAIL.n7 1.16414
R134 VTAIL.n20 VTAIL.n19 1.16414
R135 VTAIL.n32 VTAIL.n31 1.16414
R136 VTAIL.n80 VTAIL.n79 1.16414
R137 VTAIL.n68 VTAIL.n67 1.16414
R138 VTAIL.n56 VTAIL.n55 1.16414
R139 VTAIL.n44 VTAIL.n43 1.16414
R140 VTAIL.n59 VTAIL.n47 0.784983
R141 VTAIL.n83 VTAIL.n71 0.784983
R142 VTAIL.n35 VTAIL.n23 0.784983
R143 VTAIL.n71 VTAIL.n59 0.470328
R144 VTAIL.n23 VTAIL.n11 0.470328
R145 VTAIL VTAIL.n11 0.450931
R146 VTAIL.n88 VTAIL.n86 0.388379
R147 VTAIL.n4 VTAIL.n2 0.388379
R148 VTAIL.n16 VTAIL.n14 0.388379
R149 VTAIL.n28 VTAIL.n26 0.388379
R150 VTAIL.n76 VTAIL.n74 0.388379
R151 VTAIL.n64 VTAIL.n62 0.388379
R152 VTAIL.n52 VTAIL.n50 0.388379
R153 VTAIL.n40 VTAIL.n38 0.388379
R154 VTAIL VTAIL.n95 0.334552
R155 VTAIL.n93 VTAIL.n85 0.155672
R156 VTAIL.n9 VTAIL.n1 0.155672
R157 VTAIL.n21 VTAIL.n13 0.155672
R158 VTAIL.n33 VTAIL.n25 0.155672
R159 VTAIL.n81 VTAIL.n73 0.155672
R160 VTAIL.n69 VTAIL.n61 0.155672
R161 VTAIL.n57 VTAIL.n49 0.155672
R162 VTAIL.n45 VTAIL.n37 0.155672
R163 VDD1 VDD1.n1 182.206
R164 VDD1 VDD1.n0 153.524
R165 VDD1.n0 VDD1.t0 13.0547
R166 VDD1.n0 VDD1.t3 13.0547
R167 VDD1.n1 VDD1.t2 13.0547
R168 VDD1.n1 VDD1.t1 13.0547
R169 B.n209 B.n32 585
R170 B.n211 B.n210 585
R171 B.n212 B.n31 585
R172 B.n214 B.n213 585
R173 B.n215 B.n30 585
R174 B.n217 B.n216 585
R175 B.n218 B.n29 585
R176 B.n220 B.n219 585
R177 B.n221 B.n28 585
R178 B.n223 B.n222 585
R179 B.n224 B.n27 585
R180 B.n226 B.n225 585
R181 B.n227 B.n26 585
R182 B.n229 B.n228 585
R183 B.n231 B.n23 585
R184 B.n233 B.n232 585
R185 B.n234 B.n22 585
R186 B.n236 B.n235 585
R187 B.n237 B.n21 585
R188 B.n239 B.n238 585
R189 B.n240 B.n20 585
R190 B.n242 B.n241 585
R191 B.n243 B.n17 585
R192 B.n246 B.n245 585
R193 B.n247 B.n16 585
R194 B.n249 B.n248 585
R195 B.n250 B.n15 585
R196 B.n252 B.n251 585
R197 B.n253 B.n14 585
R198 B.n255 B.n254 585
R199 B.n256 B.n13 585
R200 B.n258 B.n257 585
R201 B.n259 B.n12 585
R202 B.n261 B.n260 585
R203 B.n262 B.n11 585
R204 B.n264 B.n263 585
R205 B.n265 B.n10 585
R206 B.n208 B.n207 585
R207 B.n206 B.n33 585
R208 B.n205 B.n204 585
R209 B.n203 B.n34 585
R210 B.n202 B.n201 585
R211 B.n200 B.n35 585
R212 B.n199 B.n198 585
R213 B.n197 B.n36 585
R214 B.n196 B.n195 585
R215 B.n194 B.n37 585
R216 B.n193 B.n192 585
R217 B.n191 B.n38 585
R218 B.n190 B.n189 585
R219 B.n188 B.n39 585
R220 B.n187 B.n186 585
R221 B.n185 B.n40 585
R222 B.n184 B.n183 585
R223 B.n182 B.n41 585
R224 B.n181 B.n180 585
R225 B.n179 B.n42 585
R226 B.n178 B.n177 585
R227 B.n176 B.n43 585
R228 B.n175 B.n174 585
R229 B.n173 B.n44 585
R230 B.n172 B.n171 585
R231 B.n170 B.n45 585
R232 B.n169 B.n168 585
R233 B.n167 B.n46 585
R234 B.n166 B.n165 585
R235 B.n164 B.n47 585
R236 B.n163 B.n162 585
R237 B.n161 B.n48 585
R238 B.n160 B.n159 585
R239 B.n103 B.n102 585
R240 B.n104 B.n71 585
R241 B.n106 B.n105 585
R242 B.n107 B.n70 585
R243 B.n109 B.n108 585
R244 B.n110 B.n69 585
R245 B.n112 B.n111 585
R246 B.n113 B.n68 585
R247 B.n115 B.n114 585
R248 B.n116 B.n67 585
R249 B.n118 B.n117 585
R250 B.n119 B.n66 585
R251 B.n121 B.n120 585
R252 B.n122 B.n63 585
R253 B.n125 B.n124 585
R254 B.n126 B.n62 585
R255 B.n128 B.n127 585
R256 B.n129 B.n61 585
R257 B.n131 B.n130 585
R258 B.n132 B.n60 585
R259 B.n134 B.n133 585
R260 B.n135 B.n59 585
R261 B.n137 B.n136 585
R262 B.n139 B.n138 585
R263 B.n140 B.n55 585
R264 B.n142 B.n141 585
R265 B.n143 B.n54 585
R266 B.n145 B.n144 585
R267 B.n146 B.n53 585
R268 B.n148 B.n147 585
R269 B.n149 B.n52 585
R270 B.n151 B.n150 585
R271 B.n152 B.n51 585
R272 B.n154 B.n153 585
R273 B.n155 B.n50 585
R274 B.n157 B.n156 585
R275 B.n158 B.n49 585
R276 B.n101 B.n72 585
R277 B.n100 B.n99 585
R278 B.n98 B.n73 585
R279 B.n97 B.n96 585
R280 B.n95 B.n74 585
R281 B.n94 B.n93 585
R282 B.n92 B.n75 585
R283 B.n91 B.n90 585
R284 B.n89 B.n76 585
R285 B.n88 B.n87 585
R286 B.n86 B.n77 585
R287 B.n85 B.n84 585
R288 B.n83 B.n78 585
R289 B.n82 B.n81 585
R290 B.n80 B.n79 585
R291 B.n2 B.n0 585
R292 B.n289 B.n1 585
R293 B.n288 B.n287 585
R294 B.n286 B.n3 585
R295 B.n285 B.n284 585
R296 B.n283 B.n4 585
R297 B.n282 B.n281 585
R298 B.n280 B.n5 585
R299 B.n279 B.n278 585
R300 B.n277 B.n6 585
R301 B.n276 B.n275 585
R302 B.n274 B.n7 585
R303 B.n273 B.n272 585
R304 B.n271 B.n8 585
R305 B.n270 B.n269 585
R306 B.n268 B.n9 585
R307 B.n267 B.n266 585
R308 B.n291 B.n290 585
R309 B.n102 B.n101 511.721
R310 B.n266 B.n265 511.721
R311 B.n160 B.n49 511.721
R312 B.n209 B.n208 511.721
R313 B.n56 B.t9 308.209
R314 B.n64 B.t3 308.209
R315 B.n18 B.t0 308.209
R316 B.n24 B.t6 308.209
R317 B.n56 B.t11 241.706
R318 B.n24 B.t7 241.706
R319 B.n64 B.t5 241.706
R320 B.n18 B.t1 241.706
R321 B.n57 B.t10 224.058
R322 B.n25 B.t8 224.058
R323 B.n65 B.t4 224.058
R324 B.n19 B.t2 224.058
R325 B.n101 B.n100 163.367
R326 B.n100 B.n73 163.367
R327 B.n96 B.n73 163.367
R328 B.n96 B.n95 163.367
R329 B.n95 B.n94 163.367
R330 B.n94 B.n75 163.367
R331 B.n90 B.n75 163.367
R332 B.n90 B.n89 163.367
R333 B.n89 B.n88 163.367
R334 B.n88 B.n77 163.367
R335 B.n84 B.n77 163.367
R336 B.n84 B.n83 163.367
R337 B.n83 B.n82 163.367
R338 B.n82 B.n79 163.367
R339 B.n79 B.n2 163.367
R340 B.n290 B.n2 163.367
R341 B.n290 B.n289 163.367
R342 B.n289 B.n288 163.367
R343 B.n288 B.n3 163.367
R344 B.n284 B.n3 163.367
R345 B.n284 B.n283 163.367
R346 B.n283 B.n282 163.367
R347 B.n282 B.n5 163.367
R348 B.n278 B.n5 163.367
R349 B.n278 B.n277 163.367
R350 B.n277 B.n276 163.367
R351 B.n276 B.n7 163.367
R352 B.n272 B.n7 163.367
R353 B.n272 B.n271 163.367
R354 B.n271 B.n270 163.367
R355 B.n270 B.n9 163.367
R356 B.n266 B.n9 163.367
R357 B.n102 B.n71 163.367
R358 B.n106 B.n71 163.367
R359 B.n107 B.n106 163.367
R360 B.n108 B.n107 163.367
R361 B.n108 B.n69 163.367
R362 B.n112 B.n69 163.367
R363 B.n113 B.n112 163.367
R364 B.n114 B.n113 163.367
R365 B.n114 B.n67 163.367
R366 B.n118 B.n67 163.367
R367 B.n119 B.n118 163.367
R368 B.n120 B.n119 163.367
R369 B.n120 B.n63 163.367
R370 B.n125 B.n63 163.367
R371 B.n126 B.n125 163.367
R372 B.n127 B.n126 163.367
R373 B.n127 B.n61 163.367
R374 B.n131 B.n61 163.367
R375 B.n132 B.n131 163.367
R376 B.n133 B.n132 163.367
R377 B.n133 B.n59 163.367
R378 B.n137 B.n59 163.367
R379 B.n138 B.n137 163.367
R380 B.n138 B.n55 163.367
R381 B.n142 B.n55 163.367
R382 B.n143 B.n142 163.367
R383 B.n144 B.n143 163.367
R384 B.n144 B.n53 163.367
R385 B.n148 B.n53 163.367
R386 B.n149 B.n148 163.367
R387 B.n150 B.n149 163.367
R388 B.n150 B.n51 163.367
R389 B.n154 B.n51 163.367
R390 B.n155 B.n154 163.367
R391 B.n156 B.n155 163.367
R392 B.n156 B.n49 163.367
R393 B.n161 B.n160 163.367
R394 B.n162 B.n161 163.367
R395 B.n162 B.n47 163.367
R396 B.n166 B.n47 163.367
R397 B.n167 B.n166 163.367
R398 B.n168 B.n167 163.367
R399 B.n168 B.n45 163.367
R400 B.n172 B.n45 163.367
R401 B.n173 B.n172 163.367
R402 B.n174 B.n173 163.367
R403 B.n174 B.n43 163.367
R404 B.n178 B.n43 163.367
R405 B.n179 B.n178 163.367
R406 B.n180 B.n179 163.367
R407 B.n180 B.n41 163.367
R408 B.n184 B.n41 163.367
R409 B.n185 B.n184 163.367
R410 B.n186 B.n185 163.367
R411 B.n186 B.n39 163.367
R412 B.n190 B.n39 163.367
R413 B.n191 B.n190 163.367
R414 B.n192 B.n191 163.367
R415 B.n192 B.n37 163.367
R416 B.n196 B.n37 163.367
R417 B.n197 B.n196 163.367
R418 B.n198 B.n197 163.367
R419 B.n198 B.n35 163.367
R420 B.n202 B.n35 163.367
R421 B.n203 B.n202 163.367
R422 B.n204 B.n203 163.367
R423 B.n204 B.n33 163.367
R424 B.n208 B.n33 163.367
R425 B.n265 B.n264 163.367
R426 B.n264 B.n11 163.367
R427 B.n260 B.n11 163.367
R428 B.n260 B.n259 163.367
R429 B.n259 B.n258 163.367
R430 B.n258 B.n13 163.367
R431 B.n254 B.n13 163.367
R432 B.n254 B.n253 163.367
R433 B.n253 B.n252 163.367
R434 B.n252 B.n15 163.367
R435 B.n248 B.n15 163.367
R436 B.n248 B.n247 163.367
R437 B.n247 B.n246 163.367
R438 B.n246 B.n17 163.367
R439 B.n241 B.n17 163.367
R440 B.n241 B.n240 163.367
R441 B.n240 B.n239 163.367
R442 B.n239 B.n21 163.367
R443 B.n235 B.n21 163.367
R444 B.n235 B.n234 163.367
R445 B.n234 B.n233 163.367
R446 B.n233 B.n23 163.367
R447 B.n228 B.n23 163.367
R448 B.n228 B.n227 163.367
R449 B.n227 B.n226 163.367
R450 B.n226 B.n27 163.367
R451 B.n222 B.n27 163.367
R452 B.n222 B.n221 163.367
R453 B.n221 B.n220 163.367
R454 B.n220 B.n29 163.367
R455 B.n216 B.n29 163.367
R456 B.n216 B.n215 163.367
R457 B.n215 B.n214 163.367
R458 B.n214 B.n31 163.367
R459 B.n210 B.n31 163.367
R460 B.n210 B.n209 163.367
R461 B.n58 B.n57 59.5399
R462 B.n123 B.n65 59.5399
R463 B.n244 B.n19 59.5399
R464 B.n230 B.n25 59.5399
R465 B.n267 B.n10 33.2493
R466 B.n207 B.n32 33.2493
R467 B.n159 B.n158 33.2493
R468 B.n103 B.n72 33.2493
R469 B B.n291 18.0485
R470 B.n57 B.n56 17.649
R471 B.n65 B.n64 17.649
R472 B.n19 B.n18 17.649
R473 B.n25 B.n24 17.649
R474 B.n263 B.n10 10.6151
R475 B.n263 B.n262 10.6151
R476 B.n262 B.n261 10.6151
R477 B.n261 B.n12 10.6151
R478 B.n257 B.n12 10.6151
R479 B.n257 B.n256 10.6151
R480 B.n256 B.n255 10.6151
R481 B.n255 B.n14 10.6151
R482 B.n251 B.n14 10.6151
R483 B.n251 B.n250 10.6151
R484 B.n250 B.n249 10.6151
R485 B.n249 B.n16 10.6151
R486 B.n245 B.n16 10.6151
R487 B.n243 B.n242 10.6151
R488 B.n242 B.n20 10.6151
R489 B.n238 B.n20 10.6151
R490 B.n238 B.n237 10.6151
R491 B.n237 B.n236 10.6151
R492 B.n236 B.n22 10.6151
R493 B.n232 B.n22 10.6151
R494 B.n232 B.n231 10.6151
R495 B.n229 B.n26 10.6151
R496 B.n225 B.n26 10.6151
R497 B.n225 B.n224 10.6151
R498 B.n224 B.n223 10.6151
R499 B.n223 B.n28 10.6151
R500 B.n219 B.n28 10.6151
R501 B.n219 B.n218 10.6151
R502 B.n218 B.n217 10.6151
R503 B.n217 B.n30 10.6151
R504 B.n213 B.n30 10.6151
R505 B.n213 B.n212 10.6151
R506 B.n212 B.n211 10.6151
R507 B.n211 B.n32 10.6151
R508 B.n159 B.n48 10.6151
R509 B.n163 B.n48 10.6151
R510 B.n164 B.n163 10.6151
R511 B.n165 B.n164 10.6151
R512 B.n165 B.n46 10.6151
R513 B.n169 B.n46 10.6151
R514 B.n170 B.n169 10.6151
R515 B.n171 B.n170 10.6151
R516 B.n171 B.n44 10.6151
R517 B.n175 B.n44 10.6151
R518 B.n176 B.n175 10.6151
R519 B.n177 B.n176 10.6151
R520 B.n177 B.n42 10.6151
R521 B.n181 B.n42 10.6151
R522 B.n182 B.n181 10.6151
R523 B.n183 B.n182 10.6151
R524 B.n183 B.n40 10.6151
R525 B.n187 B.n40 10.6151
R526 B.n188 B.n187 10.6151
R527 B.n189 B.n188 10.6151
R528 B.n189 B.n38 10.6151
R529 B.n193 B.n38 10.6151
R530 B.n194 B.n193 10.6151
R531 B.n195 B.n194 10.6151
R532 B.n195 B.n36 10.6151
R533 B.n199 B.n36 10.6151
R534 B.n200 B.n199 10.6151
R535 B.n201 B.n200 10.6151
R536 B.n201 B.n34 10.6151
R537 B.n205 B.n34 10.6151
R538 B.n206 B.n205 10.6151
R539 B.n207 B.n206 10.6151
R540 B.n104 B.n103 10.6151
R541 B.n105 B.n104 10.6151
R542 B.n105 B.n70 10.6151
R543 B.n109 B.n70 10.6151
R544 B.n110 B.n109 10.6151
R545 B.n111 B.n110 10.6151
R546 B.n111 B.n68 10.6151
R547 B.n115 B.n68 10.6151
R548 B.n116 B.n115 10.6151
R549 B.n117 B.n116 10.6151
R550 B.n117 B.n66 10.6151
R551 B.n121 B.n66 10.6151
R552 B.n122 B.n121 10.6151
R553 B.n124 B.n62 10.6151
R554 B.n128 B.n62 10.6151
R555 B.n129 B.n128 10.6151
R556 B.n130 B.n129 10.6151
R557 B.n130 B.n60 10.6151
R558 B.n134 B.n60 10.6151
R559 B.n135 B.n134 10.6151
R560 B.n136 B.n135 10.6151
R561 B.n140 B.n139 10.6151
R562 B.n141 B.n140 10.6151
R563 B.n141 B.n54 10.6151
R564 B.n145 B.n54 10.6151
R565 B.n146 B.n145 10.6151
R566 B.n147 B.n146 10.6151
R567 B.n147 B.n52 10.6151
R568 B.n151 B.n52 10.6151
R569 B.n152 B.n151 10.6151
R570 B.n153 B.n152 10.6151
R571 B.n153 B.n50 10.6151
R572 B.n157 B.n50 10.6151
R573 B.n158 B.n157 10.6151
R574 B.n99 B.n72 10.6151
R575 B.n99 B.n98 10.6151
R576 B.n98 B.n97 10.6151
R577 B.n97 B.n74 10.6151
R578 B.n93 B.n74 10.6151
R579 B.n93 B.n92 10.6151
R580 B.n92 B.n91 10.6151
R581 B.n91 B.n76 10.6151
R582 B.n87 B.n76 10.6151
R583 B.n87 B.n86 10.6151
R584 B.n86 B.n85 10.6151
R585 B.n85 B.n78 10.6151
R586 B.n81 B.n78 10.6151
R587 B.n81 B.n80 10.6151
R588 B.n80 B.n0 10.6151
R589 B.n287 B.n1 10.6151
R590 B.n287 B.n286 10.6151
R591 B.n286 B.n285 10.6151
R592 B.n285 B.n4 10.6151
R593 B.n281 B.n4 10.6151
R594 B.n281 B.n280 10.6151
R595 B.n280 B.n279 10.6151
R596 B.n279 B.n6 10.6151
R597 B.n275 B.n6 10.6151
R598 B.n275 B.n274 10.6151
R599 B.n274 B.n273 10.6151
R600 B.n273 B.n8 10.6151
R601 B.n269 B.n8 10.6151
R602 B.n269 B.n268 10.6151
R603 B.n268 B.n267 10.6151
R604 B.n244 B.n243 6.5566
R605 B.n231 B.n230 6.5566
R606 B.n124 B.n123 6.5566
R607 B.n136 B.n58 6.5566
R608 B.n245 B.n244 4.05904
R609 B.n230 B.n229 4.05904
R610 B.n123 B.n122 4.05904
R611 B.n139 B.n58 4.05904
R612 B.n291 B.n0 2.81026
R613 B.n291 B.n1 2.81026
R614 VN.n0 VN.t3 192.59
R615 VN.n1 VN.t0 192.59
R616 VN.n0 VN.t1 192.566
R617 VN.n1 VN.t2 192.566
R618 VN VN.n1 103.534
R619 VN VN.n0 70.265
R620 VDD2.n2 VDD2.n0 181.68
R621 VDD2.n2 VDD2.n1 153.465
R622 VDD2.n1 VDD2.t1 13.0547
R623 VDD2.n1 VDD2.t3 13.0547
R624 VDD2.n0 VDD2.t0 13.0547
R625 VDD2.n0 VDD2.t2 13.0547
R626 VDD2 VDD2.n2 0.0586897
C0 VN VTAIL 0.870484f
C1 VP VDD1 0.941068f
C2 VP VDD2 0.271726f
C3 VTAIL VDD1 2.62202f
C4 w_n1516_n1466# VP 2.16712f
C5 VP B 0.906073f
C6 VTAIL VDD2 2.66269f
C7 VN VDD1 0.152578f
C8 w_n1516_n1466# VTAIL 1.67249f
C9 VTAIL B 1.17712f
C10 VN VDD2 0.822721f
C11 VN w_n1516_n1466# 1.98058f
C12 VN B 0.60112f
C13 VTAIL VP 0.88459f
C14 VDD2 VDD1 0.541442f
C15 w_n1516_n1466# VDD1 0.779539f
C16 B VDD1 0.64719f
C17 VN VP 2.97894f
C18 w_n1516_n1466# VDD2 0.79108f
C19 B VDD2 0.667138f
C20 w_n1516_n1466# B 4.08115f
C21 VDD2 VSUBS 0.40561f
C22 VDD1 VSUBS 2.4611f
C23 VTAIL VSUBS 0.320797f
C24 VN VSUBS 3.06704f
C25 VP VSUBS 0.804339f
C26 B VSUBS 1.636137f
C27 w_n1516_n1466# VSUBS 28.2522f
C28 VDD2.t0 VSUBS 0.041986f
C29 VDD2.t2 VSUBS 0.041986f
C30 VDD2.n0 VSUBS 0.332723f
C31 VDD2.t1 VSUBS 0.041986f
C32 VDD2.t3 VSUBS 0.041986f
C33 VDD2.n1 VSUBS 0.204931f
C34 VDD2.n2 VSUBS 1.93587f
C35 VN.t3 VSUBS 0.162519f
C36 VN.t1 VSUBS 0.162502f
C37 VN.n0 VSUBS 0.173958f
C38 VN.t0 VSUBS 0.162519f
C39 VN.t2 VSUBS 0.162502f
C40 VN.n1 VSUBS 0.489621f
C41 B.n0 VSUBS 0.005395f
C42 B.n1 VSUBS 0.005395f
C43 B.n2 VSUBS 0.008531f
C44 B.n3 VSUBS 0.008531f
C45 B.n4 VSUBS 0.008531f
C46 B.n5 VSUBS 0.008531f
C47 B.n6 VSUBS 0.008531f
C48 B.n7 VSUBS 0.008531f
C49 B.n8 VSUBS 0.008531f
C50 B.n9 VSUBS 0.008531f
C51 B.n10 VSUBS 0.020839f
C52 B.n11 VSUBS 0.008531f
C53 B.n12 VSUBS 0.008531f
C54 B.n13 VSUBS 0.008531f
C55 B.n14 VSUBS 0.008531f
C56 B.n15 VSUBS 0.008531f
C57 B.n16 VSUBS 0.008531f
C58 B.n17 VSUBS 0.008531f
C59 B.t2 VSUBS 0.047014f
C60 B.t1 VSUBS 0.05254f
C61 B.t0 VSUBS 0.081106f
C62 B.n18 VSUBS 0.09329f
C63 B.n19 VSUBS 0.087852f
C64 B.n20 VSUBS 0.008531f
C65 B.n21 VSUBS 0.008531f
C66 B.n22 VSUBS 0.008531f
C67 B.n23 VSUBS 0.008531f
C68 B.t8 VSUBS 0.047014f
C69 B.t7 VSUBS 0.05254f
C70 B.t6 VSUBS 0.081106f
C71 B.n24 VSUBS 0.093289f
C72 B.n25 VSUBS 0.087852f
C73 B.n26 VSUBS 0.008531f
C74 B.n27 VSUBS 0.008531f
C75 B.n28 VSUBS 0.008531f
C76 B.n29 VSUBS 0.008531f
C77 B.n30 VSUBS 0.008531f
C78 B.n31 VSUBS 0.008531f
C79 B.n32 VSUBS 0.019849f
C80 B.n33 VSUBS 0.008531f
C81 B.n34 VSUBS 0.008531f
C82 B.n35 VSUBS 0.008531f
C83 B.n36 VSUBS 0.008531f
C84 B.n37 VSUBS 0.008531f
C85 B.n38 VSUBS 0.008531f
C86 B.n39 VSUBS 0.008531f
C87 B.n40 VSUBS 0.008531f
C88 B.n41 VSUBS 0.008531f
C89 B.n42 VSUBS 0.008531f
C90 B.n43 VSUBS 0.008531f
C91 B.n44 VSUBS 0.008531f
C92 B.n45 VSUBS 0.008531f
C93 B.n46 VSUBS 0.008531f
C94 B.n47 VSUBS 0.008531f
C95 B.n48 VSUBS 0.008531f
C96 B.n49 VSUBS 0.020839f
C97 B.n50 VSUBS 0.008531f
C98 B.n51 VSUBS 0.008531f
C99 B.n52 VSUBS 0.008531f
C100 B.n53 VSUBS 0.008531f
C101 B.n54 VSUBS 0.008531f
C102 B.n55 VSUBS 0.008531f
C103 B.t10 VSUBS 0.047014f
C104 B.t11 VSUBS 0.05254f
C105 B.t9 VSUBS 0.081106f
C106 B.n56 VSUBS 0.093289f
C107 B.n57 VSUBS 0.087852f
C108 B.n58 VSUBS 0.019766f
C109 B.n59 VSUBS 0.008531f
C110 B.n60 VSUBS 0.008531f
C111 B.n61 VSUBS 0.008531f
C112 B.n62 VSUBS 0.008531f
C113 B.n63 VSUBS 0.008531f
C114 B.t4 VSUBS 0.047014f
C115 B.t5 VSUBS 0.05254f
C116 B.t3 VSUBS 0.081106f
C117 B.n64 VSUBS 0.09329f
C118 B.n65 VSUBS 0.087852f
C119 B.n66 VSUBS 0.008531f
C120 B.n67 VSUBS 0.008531f
C121 B.n68 VSUBS 0.008531f
C122 B.n69 VSUBS 0.008531f
C123 B.n70 VSUBS 0.008531f
C124 B.n71 VSUBS 0.008531f
C125 B.n72 VSUBS 0.019559f
C126 B.n73 VSUBS 0.008531f
C127 B.n74 VSUBS 0.008531f
C128 B.n75 VSUBS 0.008531f
C129 B.n76 VSUBS 0.008531f
C130 B.n77 VSUBS 0.008531f
C131 B.n78 VSUBS 0.008531f
C132 B.n79 VSUBS 0.008531f
C133 B.n80 VSUBS 0.008531f
C134 B.n81 VSUBS 0.008531f
C135 B.n82 VSUBS 0.008531f
C136 B.n83 VSUBS 0.008531f
C137 B.n84 VSUBS 0.008531f
C138 B.n85 VSUBS 0.008531f
C139 B.n86 VSUBS 0.008531f
C140 B.n87 VSUBS 0.008531f
C141 B.n88 VSUBS 0.008531f
C142 B.n89 VSUBS 0.008531f
C143 B.n90 VSUBS 0.008531f
C144 B.n91 VSUBS 0.008531f
C145 B.n92 VSUBS 0.008531f
C146 B.n93 VSUBS 0.008531f
C147 B.n94 VSUBS 0.008531f
C148 B.n95 VSUBS 0.008531f
C149 B.n96 VSUBS 0.008531f
C150 B.n97 VSUBS 0.008531f
C151 B.n98 VSUBS 0.008531f
C152 B.n99 VSUBS 0.008531f
C153 B.n100 VSUBS 0.008531f
C154 B.n101 VSUBS 0.019559f
C155 B.n102 VSUBS 0.020839f
C156 B.n103 VSUBS 0.020839f
C157 B.n104 VSUBS 0.008531f
C158 B.n105 VSUBS 0.008531f
C159 B.n106 VSUBS 0.008531f
C160 B.n107 VSUBS 0.008531f
C161 B.n108 VSUBS 0.008531f
C162 B.n109 VSUBS 0.008531f
C163 B.n110 VSUBS 0.008531f
C164 B.n111 VSUBS 0.008531f
C165 B.n112 VSUBS 0.008531f
C166 B.n113 VSUBS 0.008531f
C167 B.n114 VSUBS 0.008531f
C168 B.n115 VSUBS 0.008531f
C169 B.n116 VSUBS 0.008531f
C170 B.n117 VSUBS 0.008531f
C171 B.n118 VSUBS 0.008531f
C172 B.n119 VSUBS 0.008531f
C173 B.n120 VSUBS 0.008531f
C174 B.n121 VSUBS 0.008531f
C175 B.n122 VSUBS 0.005897f
C176 B.n123 VSUBS 0.019766f
C177 B.n124 VSUBS 0.0069f
C178 B.n125 VSUBS 0.008531f
C179 B.n126 VSUBS 0.008531f
C180 B.n127 VSUBS 0.008531f
C181 B.n128 VSUBS 0.008531f
C182 B.n129 VSUBS 0.008531f
C183 B.n130 VSUBS 0.008531f
C184 B.n131 VSUBS 0.008531f
C185 B.n132 VSUBS 0.008531f
C186 B.n133 VSUBS 0.008531f
C187 B.n134 VSUBS 0.008531f
C188 B.n135 VSUBS 0.008531f
C189 B.n136 VSUBS 0.0069f
C190 B.n137 VSUBS 0.008531f
C191 B.n138 VSUBS 0.008531f
C192 B.n139 VSUBS 0.005897f
C193 B.n140 VSUBS 0.008531f
C194 B.n141 VSUBS 0.008531f
C195 B.n142 VSUBS 0.008531f
C196 B.n143 VSUBS 0.008531f
C197 B.n144 VSUBS 0.008531f
C198 B.n145 VSUBS 0.008531f
C199 B.n146 VSUBS 0.008531f
C200 B.n147 VSUBS 0.008531f
C201 B.n148 VSUBS 0.008531f
C202 B.n149 VSUBS 0.008531f
C203 B.n150 VSUBS 0.008531f
C204 B.n151 VSUBS 0.008531f
C205 B.n152 VSUBS 0.008531f
C206 B.n153 VSUBS 0.008531f
C207 B.n154 VSUBS 0.008531f
C208 B.n155 VSUBS 0.008531f
C209 B.n156 VSUBS 0.008531f
C210 B.n157 VSUBS 0.008531f
C211 B.n158 VSUBS 0.020839f
C212 B.n159 VSUBS 0.019559f
C213 B.n160 VSUBS 0.019559f
C214 B.n161 VSUBS 0.008531f
C215 B.n162 VSUBS 0.008531f
C216 B.n163 VSUBS 0.008531f
C217 B.n164 VSUBS 0.008531f
C218 B.n165 VSUBS 0.008531f
C219 B.n166 VSUBS 0.008531f
C220 B.n167 VSUBS 0.008531f
C221 B.n168 VSUBS 0.008531f
C222 B.n169 VSUBS 0.008531f
C223 B.n170 VSUBS 0.008531f
C224 B.n171 VSUBS 0.008531f
C225 B.n172 VSUBS 0.008531f
C226 B.n173 VSUBS 0.008531f
C227 B.n174 VSUBS 0.008531f
C228 B.n175 VSUBS 0.008531f
C229 B.n176 VSUBS 0.008531f
C230 B.n177 VSUBS 0.008531f
C231 B.n178 VSUBS 0.008531f
C232 B.n179 VSUBS 0.008531f
C233 B.n180 VSUBS 0.008531f
C234 B.n181 VSUBS 0.008531f
C235 B.n182 VSUBS 0.008531f
C236 B.n183 VSUBS 0.008531f
C237 B.n184 VSUBS 0.008531f
C238 B.n185 VSUBS 0.008531f
C239 B.n186 VSUBS 0.008531f
C240 B.n187 VSUBS 0.008531f
C241 B.n188 VSUBS 0.008531f
C242 B.n189 VSUBS 0.008531f
C243 B.n190 VSUBS 0.008531f
C244 B.n191 VSUBS 0.008531f
C245 B.n192 VSUBS 0.008531f
C246 B.n193 VSUBS 0.008531f
C247 B.n194 VSUBS 0.008531f
C248 B.n195 VSUBS 0.008531f
C249 B.n196 VSUBS 0.008531f
C250 B.n197 VSUBS 0.008531f
C251 B.n198 VSUBS 0.008531f
C252 B.n199 VSUBS 0.008531f
C253 B.n200 VSUBS 0.008531f
C254 B.n201 VSUBS 0.008531f
C255 B.n202 VSUBS 0.008531f
C256 B.n203 VSUBS 0.008531f
C257 B.n204 VSUBS 0.008531f
C258 B.n205 VSUBS 0.008531f
C259 B.n206 VSUBS 0.008531f
C260 B.n207 VSUBS 0.02055f
C261 B.n208 VSUBS 0.019559f
C262 B.n209 VSUBS 0.020839f
C263 B.n210 VSUBS 0.008531f
C264 B.n211 VSUBS 0.008531f
C265 B.n212 VSUBS 0.008531f
C266 B.n213 VSUBS 0.008531f
C267 B.n214 VSUBS 0.008531f
C268 B.n215 VSUBS 0.008531f
C269 B.n216 VSUBS 0.008531f
C270 B.n217 VSUBS 0.008531f
C271 B.n218 VSUBS 0.008531f
C272 B.n219 VSUBS 0.008531f
C273 B.n220 VSUBS 0.008531f
C274 B.n221 VSUBS 0.008531f
C275 B.n222 VSUBS 0.008531f
C276 B.n223 VSUBS 0.008531f
C277 B.n224 VSUBS 0.008531f
C278 B.n225 VSUBS 0.008531f
C279 B.n226 VSUBS 0.008531f
C280 B.n227 VSUBS 0.008531f
C281 B.n228 VSUBS 0.008531f
C282 B.n229 VSUBS 0.005897f
C283 B.n230 VSUBS 0.019766f
C284 B.n231 VSUBS 0.0069f
C285 B.n232 VSUBS 0.008531f
C286 B.n233 VSUBS 0.008531f
C287 B.n234 VSUBS 0.008531f
C288 B.n235 VSUBS 0.008531f
C289 B.n236 VSUBS 0.008531f
C290 B.n237 VSUBS 0.008531f
C291 B.n238 VSUBS 0.008531f
C292 B.n239 VSUBS 0.008531f
C293 B.n240 VSUBS 0.008531f
C294 B.n241 VSUBS 0.008531f
C295 B.n242 VSUBS 0.008531f
C296 B.n243 VSUBS 0.0069f
C297 B.n244 VSUBS 0.019766f
C298 B.n245 VSUBS 0.005897f
C299 B.n246 VSUBS 0.008531f
C300 B.n247 VSUBS 0.008531f
C301 B.n248 VSUBS 0.008531f
C302 B.n249 VSUBS 0.008531f
C303 B.n250 VSUBS 0.008531f
C304 B.n251 VSUBS 0.008531f
C305 B.n252 VSUBS 0.008531f
C306 B.n253 VSUBS 0.008531f
C307 B.n254 VSUBS 0.008531f
C308 B.n255 VSUBS 0.008531f
C309 B.n256 VSUBS 0.008531f
C310 B.n257 VSUBS 0.008531f
C311 B.n258 VSUBS 0.008531f
C312 B.n259 VSUBS 0.008531f
C313 B.n260 VSUBS 0.008531f
C314 B.n261 VSUBS 0.008531f
C315 B.n262 VSUBS 0.008531f
C316 B.n263 VSUBS 0.008531f
C317 B.n264 VSUBS 0.008531f
C318 B.n265 VSUBS 0.020839f
C319 B.n266 VSUBS 0.019559f
C320 B.n267 VSUBS 0.019559f
C321 B.n268 VSUBS 0.008531f
C322 B.n269 VSUBS 0.008531f
C323 B.n270 VSUBS 0.008531f
C324 B.n271 VSUBS 0.008531f
C325 B.n272 VSUBS 0.008531f
C326 B.n273 VSUBS 0.008531f
C327 B.n274 VSUBS 0.008531f
C328 B.n275 VSUBS 0.008531f
C329 B.n276 VSUBS 0.008531f
C330 B.n277 VSUBS 0.008531f
C331 B.n278 VSUBS 0.008531f
C332 B.n279 VSUBS 0.008531f
C333 B.n280 VSUBS 0.008531f
C334 B.n281 VSUBS 0.008531f
C335 B.n282 VSUBS 0.008531f
C336 B.n283 VSUBS 0.008531f
C337 B.n284 VSUBS 0.008531f
C338 B.n285 VSUBS 0.008531f
C339 B.n286 VSUBS 0.008531f
C340 B.n287 VSUBS 0.008531f
C341 B.n288 VSUBS 0.008531f
C342 B.n289 VSUBS 0.008531f
C343 B.n290 VSUBS 0.008531f
C344 B.n291 VSUBS 0.019318f
C345 VDD1.t0 VSUBS 0.039285f
C346 VDD1.t3 VSUBS 0.039285f
C347 VDD1.n0 VSUBS 0.191856f
C348 VDD1.t2 VSUBS 0.039285f
C349 VDD1.t1 VSUBS 0.039285f
C350 VDD1.n1 VSUBS 0.319706f
C351 VTAIL.n0 VSUBS 0.017325f
C352 VTAIL.n1 VSUBS 0.116217f
C353 VTAIL.n2 VSUBS 0.008884f
C354 VTAIL.t3 VSUBS 0.046685f
C355 VTAIL.n3 VSUBS 0.054767f
C356 VTAIL.n4 VSUBS 0.012381f
C357 VTAIL.n5 VSUBS 0.015748f
C358 VTAIL.n6 VSUBS 0.047972f
C359 VTAIL.n7 VSUBS 0.009406f
C360 VTAIL.n8 VSUBS 0.008884f
C361 VTAIL.n9 VSUBS 0.040246f
C362 VTAIL.n10 VSUBS 0.024059f
C363 VTAIL.n11 VSUBS 0.064291f
C364 VTAIL.n12 VSUBS 0.017325f
C365 VTAIL.n13 VSUBS 0.116217f
C366 VTAIL.n14 VSUBS 0.008884f
C367 VTAIL.t4 VSUBS 0.046685f
C368 VTAIL.n15 VSUBS 0.054767f
C369 VTAIL.n16 VSUBS 0.012381f
C370 VTAIL.n17 VSUBS 0.015748f
C371 VTAIL.n18 VSUBS 0.047972f
C372 VTAIL.n19 VSUBS 0.009406f
C373 VTAIL.n20 VSUBS 0.008884f
C374 VTAIL.n21 VSUBS 0.040246f
C375 VTAIL.n22 VSUBS 0.024059f
C376 VTAIL.n23 VSUBS 0.082086f
C377 VTAIL.n24 VSUBS 0.017325f
C378 VTAIL.n25 VSUBS 0.116217f
C379 VTAIL.n26 VSUBS 0.008884f
C380 VTAIL.t5 VSUBS 0.046685f
C381 VTAIL.n27 VSUBS 0.054767f
C382 VTAIL.n28 VSUBS 0.012381f
C383 VTAIL.n29 VSUBS 0.015748f
C384 VTAIL.n30 VSUBS 0.047972f
C385 VTAIL.n31 VSUBS 0.009406f
C386 VTAIL.n32 VSUBS 0.008884f
C387 VTAIL.n33 VSUBS 0.040246f
C388 VTAIL.n34 VSUBS 0.024059f
C389 VTAIL.n35 VSUBS 0.437766f
C390 VTAIL.n36 VSUBS 0.017325f
C391 VTAIL.n37 VSUBS 0.116217f
C392 VTAIL.n38 VSUBS 0.008884f
C393 VTAIL.t0 VSUBS 0.046685f
C394 VTAIL.n39 VSUBS 0.054767f
C395 VTAIL.n40 VSUBS 0.012381f
C396 VTAIL.n41 VSUBS 0.015748f
C397 VTAIL.n42 VSUBS 0.047972f
C398 VTAIL.n43 VSUBS 0.009406f
C399 VTAIL.n44 VSUBS 0.008884f
C400 VTAIL.n45 VSUBS 0.040246f
C401 VTAIL.n46 VSUBS 0.024059f
C402 VTAIL.n47 VSUBS 0.437766f
C403 VTAIL.n48 VSUBS 0.017325f
C404 VTAIL.n49 VSUBS 0.116217f
C405 VTAIL.n50 VSUBS 0.008884f
C406 VTAIL.t1 VSUBS 0.046685f
C407 VTAIL.n51 VSUBS 0.054767f
C408 VTAIL.n52 VSUBS 0.012381f
C409 VTAIL.n53 VSUBS 0.015748f
C410 VTAIL.n54 VSUBS 0.047972f
C411 VTAIL.n55 VSUBS 0.009406f
C412 VTAIL.n56 VSUBS 0.008884f
C413 VTAIL.n57 VSUBS 0.040246f
C414 VTAIL.n58 VSUBS 0.024059f
C415 VTAIL.n59 VSUBS 0.082086f
C416 VTAIL.n60 VSUBS 0.017325f
C417 VTAIL.n61 VSUBS 0.116217f
C418 VTAIL.n62 VSUBS 0.008884f
C419 VTAIL.t7 VSUBS 0.046685f
C420 VTAIL.n63 VSUBS 0.054767f
C421 VTAIL.n64 VSUBS 0.012381f
C422 VTAIL.n65 VSUBS 0.015748f
C423 VTAIL.n66 VSUBS 0.047972f
C424 VTAIL.n67 VSUBS 0.009406f
C425 VTAIL.n68 VSUBS 0.008884f
C426 VTAIL.n69 VSUBS 0.040246f
C427 VTAIL.n70 VSUBS 0.024059f
C428 VTAIL.n71 VSUBS 0.082086f
C429 VTAIL.n72 VSUBS 0.017325f
C430 VTAIL.n73 VSUBS 0.116217f
C431 VTAIL.n74 VSUBS 0.008884f
C432 VTAIL.t6 VSUBS 0.046685f
C433 VTAIL.n75 VSUBS 0.054767f
C434 VTAIL.n76 VSUBS 0.012381f
C435 VTAIL.n77 VSUBS 0.015748f
C436 VTAIL.n78 VSUBS 0.047972f
C437 VTAIL.n79 VSUBS 0.009406f
C438 VTAIL.n80 VSUBS 0.008884f
C439 VTAIL.n81 VSUBS 0.040246f
C440 VTAIL.n82 VSUBS 0.024059f
C441 VTAIL.n83 VSUBS 0.437766f
C442 VTAIL.n84 VSUBS 0.017325f
C443 VTAIL.n85 VSUBS 0.116217f
C444 VTAIL.n86 VSUBS 0.008884f
C445 VTAIL.t2 VSUBS 0.046685f
C446 VTAIL.n87 VSUBS 0.054767f
C447 VTAIL.n88 VSUBS 0.012381f
C448 VTAIL.n89 VSUBS 0.015748f
C449 VTAIL.n90 VSUBS 0.047972f
C450 VTAIL.n91 VSUBS 0.009406f
C451 VTAIL.n92 VSUBS 0.008884f
C452 VTAIL.n93 VSUBS 0.040246f
C453 VTAIL.n94 VSUBS 0.024059f
C454 VTAIL.n95 VSUBS 0.413772f
C455 VP.t0 VSUBS 0.286307f
C456 VP.t3 VSUBS 0.286336f
C457 VP.n0 VSUBS 0.845335f
C458 VP.n1 VSUBS 2.82377f
C459 VP.t1 VSUBS 0.267602f
C460 VP.n2 VSUBS 0.171873f
C461 VP.t2 VSUBS 0.267602f
C462 VP.n3 VSUBS 0.171873f
C463 VP.n4 VSUBS 0.047195f
.ends

