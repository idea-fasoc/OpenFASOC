* NGSPICE file created from diff_pair_sample_0418.ext - technology: sky130A

.subckt diff_pair_sample_0418 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X1 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=0 ps=0 w=8.23 l=1.68
X2 VDD1.t2 VP.t1 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X3 VTAIL.t17 VP.t2 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X4 VDD1.t7 VP.t3 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=3.2097 ps=17.24 w=8.23 l=1.68
X5 VTAIL.t1 VN.t0 VDD2.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X6 VDD1.t3 VP.t4 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=3.2097 ps=17.24 w=8.23 l=1.68
X7 VTAIL.t14 VP.t5 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X8 VDD1.t0 VP.t6 VTAIL.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X9 VTAIL.t12 VP.t7 VDD1.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X10 VDD2.t8 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=1.35795 ps=8.56 w=8.23 l=1.68
X11 VDD2.t7 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=3.2097 ps=17.24 w=8.23 l=1.68
X12 VDD2.t6 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X13 VTAIL.t0 VN.t4 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X14 VDD2.t4 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=3.2097 ps=17.24 w=8.23 l=1.68
X15 VDD2.t3 VN.t6 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=1.35795 ps=8.56 w=8.23 l=1.68
X16 VTAIL.t3 VN.t7 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X17 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=0 ps=0 w=8.23 l=1.68
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=0 ps=0 w=8.23 l=1.68
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=0 ps=0 w=8.23 l=1.68
X20 VTAIL.t7 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
X21 VDD1.t5 VP.t8 VTAIL.t11 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=1.35795 ps=8.56 w=8.23 l=1.68
X22 VDD1.t8 VP.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2097 pd=17.24 as=1.35795 ps=8.56 w=8.23 l=1.68
X23 VDD2.t0 VN.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.35795 pd=8.56 as=1.35795 ps=8.56 w=8.23 l=1.68
R0 VP.n41 VP.n40 184.788
R1 VP.n70 VP.n69 184.788
R2 VP.n39 VP.n38 184.788
R3 VP.n18 VP.n15 161.3
R4 VP.n20 VP.n19 161.3
R5 VP.n21 VP.n14 161.3
R6 VP.n23 VP.n22 161.3
R7 VP.n24 VP.n13 161.3
R8 VP.n26 VP.n25 161.3
R9 VP.n27 VP.n12 161.3
R10 VP.n29 VP.n28 161.3
R11 VP.n30 VP.n11 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n34 VP.n10 161.3
R14 VP.n36 VP.n35 161.3
R15 VP.n37 VP.n9 161.3
R16 VP.n68 VP.n0 161.3
R17 VP.n67 VP.n66 161.3
R18 VP.n65 VP.n1 161.3
R19 VP.n64 VP.n63 161.3
R20 VP.n61 VP.n2 161.3
R21 VP.n60 VP.n59 161.3
R22 VP.n58 VP.n3 161.3
R23 VP.n57 VP.n56 161.3
R24 VP.n55 VP.n4 161.3
R25 VP.n54 VP.n53 161.3
R26 VP.n52 VP.n5 161.3
R27 VP.n51 VP.n50 161.3
R28 VP.n49 VP.n6 161.3
R29 VP.n47 VP.n46 161.3
R30 VP.n45 VP.n7 161.3
R31 VP.n44 VP.n43 161.3
R32 VP.n42 VP.n8 161.3
R33 VP.n16 VP.t8 145.749
R34 VP.n55 VP.t6 118.061
R35 VP.n41 VP.t9 118.061
R36 VP.n48 VP.t2 118.061
R37 VP.n62 VP.t5 118.061
R38 VP.n69 VP.t4 118.061
R39 VP.n24 VP.t1 118.061
R40 VP.n38 VP.t3 118.061
R41 VP.n31 VP.t7 118.061
R42 VP.n17 VP.t0 118.061
R43 VP.n17 VP.n16 68.3921
R44 VP.n40 VP.n39 45.0876
R45 VP.n43 VP.n7 41.9503
R46 VP.n67 VP.n1 41.9503
R47 VP.n36 VP.n10 41.9503
R48 VP.n50 VP.n5 40.979
R49 VP.n60 VP.n3 40.979
R50 VP.n29 VP.n12 40.979
R51 VP.n19 VP.n14 40.979
R52 VP.n54 VP.n5 40.0078
R53 VP.n56 VP.n3 40.0078
R54 VP.n25 VP.n12 40.0078
R55 VP.n23 VP.n14 40.0078
R56 VP.n47 VP.n7 39.0365
R57 VP.n63 VP.n1 39.0365
R58 VP.n32 VP.n10 39.0365
R59 VP.n43 VP.n42 24.4675
R60 VP.n50 VP.n49 24.4675
R61 VP.n55 VP.n54 24.4675
R62 VP.n56 VP.n55 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n68 VP.n67 24.4675
R65 VP.n37 VP.n36 24.4675
R66 VP.n30 VP.n29 24.4675
R67 VP.n24 VP.n23 24.4675
R68 VP.n25 VP.n24 24.4675
R69 VP.n19 VP.n18 24.4675
R70 VP.n48 VP.n47 23.9782
R71 VP.n63 VP.n62 23.9782
R72 VP.n32 VP.n31 23.9782
R73 VP.n16 VP.n15 18.9635
R74 VP.n42 VP.n41 0.97918
R75 VP.n69 VP.n68 0.97918
R76 VP.n38 VP.n37 0.97918
R77 VP.n49 VP.n48 0.48984
R78 VP.n62 VP.n61 0.48984
R79 VP.n31 VP.n30 0.48984
R80 VP.n18 VP.n17 0.48984
R81 VP.n20 VP.n15 0.189894
R82 VP.n21 VP.n20 0.189894
R83 VP.n22 VP.n21 0.189894
R84 VP.n22 VP.n13 0.189894
R85 VP.n26 VP.n13 0.189894
R86 VP.n27 VP.n26 0.189894
R87 VP.n28 VP.n27 0.189894
R88 VP.n28 VP.n11 0.189894
R89 VP.n33 VP.n11 0.189894
R90 VP.n34 VP.n33 0.189894
R91 VP.n35 VP.n34 0.189894
R92 VP.n35 VP.n9 0.189894
R93 VP.n39 VP.n9 0.189894
R94 VP.n40 VP.n8 0.189894
R95 VP.n44 VP.n8 0.189894
R96 VP.n45 VP.n44 0.189894
R97 VP.n46 VP.n45 0.189894
R98 VP.n46 VP.n6 0.189894
R99 VP.n51 VP.n6 0.189894
R100 VP.n52 VP.n51 0.189894
R101 VP.n53 VP.n52 0.189894
R102 VP.n53 VP.n4 0.189894
R103 VP.n57 VP.n4 0.189894
R104 VP.n58 VP.n57 0.189894
R105 VP.n59 VP.n58 0.189894
R106 VP.n59 VP.n2 0.189894
R107 VP.n64 VP.n2 0.189894
R108 VP.n65 VP.n64 0.189894
R109 VP.n66 VP.n65 0.189894
R110 VP.n66 VP.n0 0.189894
R111 VP.n70 VP.n0 0.189894
R112 VP VP.n70 0.0516364
R113 VDD1.n1 VDD1.t5 69.1918
R114 VDD1.n3 VDD1.t8 69.1917
R115 VDD1.n5 VDD1.n4 66.2973
R116 VDD1.n1 VDD1.n0 65.0533
R117 VDD1.n7 VDD1.n6 65.0531
R118 VDD1.n3 VDD1.n2 65.053
R119 VDD1.n7 VDD1.n5 40.4901
R120 VDD1.n6 VDD1.t9 2.40633
R121 VDD1.n6 VDD1.t7 2.40633
R122 VDD1.n0 VDD1.t1 2.40633
R123 VDD1.n0 VDD1.t2 2.40633
R124 VDD1.n4 VDD1.t6 2.40633
R125 VDD1.n4 VDD1.t3 2.40633
R126 VDD1.n2 VDD1.t4 2.40633
R127 VDD1.n2 VDD1.t0 2.40633
R128 VDD1 VDD1.n7 1.24188
R129 VDD1 VDD1.n1 0.491879
R130 VDD1.n5 VDD1.n3 0.378344
R131 VTAIL.n11 VTAIL.t5 50.7803
R132 VTAIL.n17 VTAIL.t6 50.7802
R133 VTAIL.n2 VTAIL.t15 50.7802
R134 VTAIL.n16 VTAIL.t16 50.7802
R135 VTAIL.n15 VTAIL.n14 48.3745
R136 VTAIL.n13 VTAIL.n12 48.3745
R137 VTAIL.n10 VTAIL.n9 48.3745
R138 VTAIL.n8 VTAIL.n7 48.3745
R139 VTAIL.n19 VTAIL.n18 48.3743
R140 VTAIL.n1 VTAIL.n0 48.3743
R141 VTAIL.n4 VTAIL.n3 48.3743
R142 VTAIL.n6 VTAIL.n5 48.3743
R143 VTAIL.n8 VTAIL.n6 22.9272
R144 VTAIL.n17 VTAIL.n16 21.1945
R145 VTAIL.n18 VTAIL.t4 2.40633
R146 VTAIL.n18 VTAIL.t0 2.40633
R147 VTAIL.n0 VTAIL.t8 2.40633
R148 VTAIL.n0 VTAIL.t3 2.40633
R149 VTAIL.n3 VTAIL.t13 2.40633
R150 VTAIL.n3 VTAIL.t14 2.40633
R151 VTAIL.n5 VTAIL.t10 2.40633
R152 VTAIL.n5 VTAIL.t17 2.40633
R153 VTAIL.n14 VTAIL.t18 2.40633
R154 VTAIL.n14 VTAIL.t12 2.40633
R155 VTAIL.n12 VTAIL.t11 2.40633
R156 VTAIL.n12 VTAIL.t19 2.40633
R157 VTAIL.n9 VTAIL.t9 2.40633
R158 VTAIL.n9 VTAIL.t7 2.40633
R159 VTAIL.n7 VTAIL.t2 2.40633
R160 VTAIL.n7 VTAIL.t1 2.40633
R161 VTAIL.n10 VTAIL.n8 1.73326
R162 VTAIL.n11 VTAIL.n10 1.73326
R163 VTAIL.n15 VTAIL.n13 1.73326
R164 VTAIL.n16 VTAIL.n15 1.73326
R165 VTAIL.n6 VTAIL.n4 1.73326
R166 VTAIL.n4 VTAIL.n2 1.73326
R167 VTAIL.n19 VTAIL.n17 1.73326
R168 VTAIL VTAIL.n1 1.35826
R169 VTAIL.n13 VTAIL.n11 1.33671
R170 VTAIL.n2 VTAIL.n1 1.33671
R171 VTAIL VTAIL.n19 0.3755
R172 B.n713 B.n712 585
R173 B.n714 B.n713 585
R174 B.n259 B.n117 585
R175 B.n258 B.n257 585
R176 B.n256 B.n255 585
R177 B.n254 B.n253 585
R178 B.n252 B.n251 585
R179 B.n250 B.n249 585
R180 B.n248 B.n247 585
R181 B.n246 B.n245 585
R182 B.n244 B.n243 585
R183 B.n242 B.n241 585
R184 B.n240 B.n239 585
R185 B.n238 B.n237 585
R186 B.n236 B.n235 585
R187 B.n234 B.n233 585
R188 B.n232 B.n231 585
R189 B.n230 B.n229 585
R190 B.n228 B.n227 585
R191 B.n226 B.n225 585
R192 B.n224 B.n223 585
R193 B.n222 B.n221 585
R194 B.n220 B.n219 585
R195 B.n218 B.n217 585
R196 B.n216 B.n215 585
R197 B.n214 B.n213 585
R198 B.n212 B.n211 585
R199 B.n210 B.n209 585
R200 B.n208 B.n207 585
R201 B.n206 B.n205 585
R202 B.n204 B.n203 585
R203 B.n202 B.n201 585
R204 B.n200 B.n199 585
R205 B.n198 B.n197 585
R206 B.n196 B.n195 585
R207 B.n194 B.n193 585
R208 B.n192 B.n191 585
R209 B.n190 B.n189 585
R210 B.n188 B.n187 585
R211 B.n186 B.n185 585
R212 B.n184 B.n183 585
R213 B.n181 B.n180 585
R214 B.n179 B.n178 585
R215 B.n177 B.n176 585
R216 B.n175 B.n174 585
R217 B.n173 B.n172 585
R218 B.n171 B.n170 585
R219 B.n169 B.n168 585
R220 B.n167 B.n166 585
R221 B.n165 B.n164 585
R222 B.n163 B.n162 585
R223 B.n161 B.n160 585
R224 B.n159 B.n158 585
R225 B.n157 B.n156 585
R226 B.n155 B.n154 585
R227 B.n153 B.n152 585
R228 B.n151 B.n150 585
R229 B.n149 B.n148 585
R230 B.n147 B.n146 585
R231 B.n145 B.n144 585
R232 B.n143 B.n142 585
R233 B.n141 B.n140 585
R234 B.n139 B.n138 585
R235 B.n137 B.n136 585
R236 B.n135 B.n134 585
R237 B.n133 B.n132 585
R238 B.n131 B.n130 585
R239 B.n129 B.n128 585
R240 B.n127 B.n126 585
R241 B.n125 B.n124 585
R242 B.n82 B.n81 585
R243 B.n717 B.n716 585
R244 B.n711 B.n118 585
R245 B.n118 B.n79 585
R246 B.n710 B.n78 585
R247 B.n721 B.n78 585
R248 B.n709 B.n77 585
R249 B.n722 B.n77 585
R250 B.n708 B.n76 585
R251 B.n723 B.n76 585
R252 B.n707 B.n706 585
R253 B.n706 B.n72 585
R254 B.n705 B.n71 585
R255 B.n729 B.n71 585
R256 B.n704 B.n70 585
R257 B.n730 B.n70 585
R258 B.n703 B.n69 585
R259 B.n731 B.n69 585
R260 B.n702 B.n701 585
R261 B.n701 B.n65 585
R262 B.n700 B.n64 585
R263 B.n737 B.n64 585
R264 B.n699 B.n63 585
R265 B.n738 B.n63 585
R266 B.n698 B.n62 585
R267 B.n739 B.n62 585
R268 B.n697 B.n696 585
R269 B.n696 B.n58 585
R270 B.n695 B.n57 585
R271 B.n745 B.n57 585
R272 B.n694 B.n56 585
R273 B.n746 B.n56 585
R274 B.n693 B.n55 585
R275 B.n747 B.n55 585
R276 B.n692 B.n691 585
R277 B.n691 B.n51 585
R278 B.n690 B.n50 585
R279 B.n753 B.n50 585
R280 B.n689 B.n49 585
R281 B.n754 B.n49 585
R282 B.n688 B.n48 585
R283 B.n755 B.n48 585
R284 B.n687 B.n686 585
R285 B.n686 B.n44 585
R286 B.n685 B.n43 585
R287 B.n761 B.n43 585
R288 B.n684 B.n42 585
R289 B.n762 B.n42 585
R290 B.n683 B.n41 585
R291 B.n763 B.n41 585
R292 B.n682 B.n681 585
R293 B.n681 B.n37 585
R294 B.n680 B.n36 585
R295 B.n769 B.n36 585
R296 B.n679 B.n35 585
R297 B.n770 B.n35 585
R298 B.n678 B.n34 585
R299 B.n771 B.n34 585
R300 B.n677 B.n676 585
R301 B.n676 B.n30 585
R302 B.n675 B.n29 585
R303 B.n777 B.n29 585
R304 B.n674 B.n28 585
R305 B.n778 B.n28 585
R306 B.n673 B.n27 585
R307 B.n779 B.n27 585
R308 B.n672 B.n671 585
R309 B.n671 B.n23 585
R310 B.n670 B.n22 585
R311 B.n785 B.n22 585
R312 B.n669 B.n21 585
R313 B.n786 B.n21 585
R314 B.n668 B.n20 585
R315 B.n787 B.n20 585
R316 B.n667 B.n666 585
R317 B.n666 B.n16 585
R318 B.n665 B.n15 585
R319 B.n793 B.n15 585
R320 B.n664 B.n14 585
R321 B.n794 B.n14 585
R322 B.n663 B.n13 585
R323 B.n795 B.n13 585
R324 B.n662 B.n661 585
R325 B.n661 B.n12 585
R326 B.n660 B.n659 585
R327 B.n660 B.n8 585
R328 B.n658 B.n7 585
R329 B.n802 B.n7 585
R330 B.n657 B.n6 585
R331 B.n803 B.n6 585
R332 B.n656 B.n5 585
R333 B.n804 B.n5 585
R334 B.n655 B.n654 585
R335 B.n654 B.n4 585
R336 B.n653 B.n260 585
R337 B.n653 B.n652 585
R338 B.n643 B.n261 585
R339 B.n262 B.n261 585
R340 B.n645 B.n644 585
R341 B.n646 B.n645 585
R342 B.n642 B.n266 585
R343 B.n270 B.n266 585
R344 B.n641 B.n640 585
R345 B.n640 B.n639 585
R346 B.n268 B.n267 585
R347 B.n269 B.n268 585
R348 B.n632 B.n631 585
R349 B.n633 B.n632 585
R350 B.n630 B.n275 585
R351 B.n275 B.n274 585
R352 B.n629 B.n628 585
R353 B.n628 B.n627 585
R354 B.n277 B.n276 585
R355 B.n278 B.n277 585
R356 B.n620 B.n619 585
R357 B.n621 B.n620 585
R358 B.n618 B.n283 585
R359 B.n283 B.n282 585
R360 B.n617 B.n616 585
R361 B.n616 B.n615 585
R362 B.n285 B.n284 585
R363 B.n286 B.n285 585
R364 B.n608 B.n607 585
R365 B.n609 B.n608 585
R366 B.n606 B.n291 585
R367 B.n291 B.n290 585
R368 B.n605 B.n604 585
R369 B.n604 B.n603 585
R370 B.n293 B.n292 585
R371 B.n294 B.n293 585
R372 B.n596 B.n595 585
R373 B.n597 B.n596 585
R374 B.n594 B.n299 585
R375 B.n299 B.n298 585
R376 B.n593 B.n592 585
R377 B.n592 B.n591 585
R378 B.n301 B.n300 585
R379 B.n302 B.n301 585
R380 B.n584 B.n583 585
R381 B.n585 B.n584 585
R382 B.n582 B.n307 585
R383 B.n307 B.n306 585
R384 B.n581 B.n580 585
R385 B.n580 B.n579 585
R386 B.n309 B.n308 585
R387 B.n310 B.n309 585
R388 B.n572 B.n571 585
R389 B.n573 B.n572 585
R390 B.n570 B.n315 585
R391 B.n315 B.n314 585
R392 B.n569 B.n568 585
R393 B.n568 B.n567 585
R394 B.n317 B.n316 585
R395 B.n318 B.n317 585
R396 B.n560 B.n559 585
R397 B.n561 B.n560 585
R398 B.n558 B.n323 585
R399 B.n323 B.n322 585
R400 B.n557 B.n556 585
R401 B.n556 B.n555 585
R402 B.n325 B.n324 585
R403 B.n326 B.n325 585
R404 B.n548 B.n547 585
R405 B.n549 B.n548 585
R406 B.n546 B.n330 585
R407 B.n334 B.n330 585
R408 B.n545 B.n544 585
R409 B.n544 B.n543 585
R410 B.n332 B.n331 585
R411 B.n333 B.n332 585
R412 B.n536 B.n535 585
R413 B.n537 B.n536 585
R414 B.n534 B.n339 585
R415 B.n339 B.n338 585
R416 B.n533 B.n532 585
R417 B.n532 B.n531 585
R418 B.n341 B.n340 585
R419 B.n342 B.n341 585
R420 B.n527 B.n526 585
R421 B.n345 B.n344 585
R422 B.n523 B.n522 585
R423 B.n524 B.n523 585
R424 B.n521 B.n380 585
R425 B.n520 B.n519 585
R426 B.n518 B.n517 585
R427 B.n516 B.n515 585
R428 B.n514 B.n513 585
R429 B.n512 B.n511 585
R430 B.n510 B.n509 585
R431 B.n508 B.n507 585
R432 B.n506 B.n505 585
R433 B.n504 B.n503 585
R434 B.n502 B.n501 585
R435 B.n500 B.n499 585
R436 B.n498 B.n497 585
R437 B.n496 B.n495 585
R438 B.n494 B.n493 585
R439 B.n492 B.n491 585
R440 B.n490 B.n489 585
R441 B.n488 B.n487 585
R442 B.n486 B.n485 585
R443 B.n484 B.n483 585
R444 B.n482 B.n481 585
R445 B.n480 B.n479 585
R446 B.n478 B.n477 585
R447 B.n476 B.n475 585
R448 B.n474 B.n473 585
R449 B.n472 B.n471 585
R450 B.n470 B.n469 585
R451 B.n468 B.n467 585
R452 B.n466 B.n465 585
R453 B.n464 B.n463 585
R454 B.n462 B.n461 585
R455 B.n460 B.n459 585
R456 B.n458 B.n457 585
R457 B.n456 B.n455 585
R458 B.n454 B.n453 585
R459 B.n452 B.n451 585
R460 B.n450 B.n449 585
R461 B.n447 B.n446 585
R462 B.n445 B.n444 585
R463 B.n443 B.n442 585
R464 B.n441 B.n440 585
R465 B.n439 B.n438 585
R466 B.n437 B.n436 585
R467 B.n435 B.n434 585
R468 B.n433 B.n432 585
R469 B.n431 B.n430 585
R470 B.n429 B.n428 585
R471 B.n427 B.n426 585
R472 B.n425 B.n424 585
R473 B.n423 B.n422 585
R474 B.n421 B.n420 585
R475 B.n419 B.n418 585
R476 B.n417 B.n416 585
R477 B.n415 B.n414 585
R478 B.n413 B.n412 585
R479 B.n411 B.n410 585
R480 B.n409 B.n408 585
R481 B.n407 B.n406 585
R482 B.n405 B.n404 585
R483 B.n403 B.n402 585
R484 B.n401 B.n400 585
R485 B.n399 B.n398 585
R486 B.n397 B.n396 585
R487 B.n395 B.n394 585
R488 B.n393 B.n392 585
R489 B.n391 B.n390 585
R490 B.n389 B.n388 585
R491 B.n387 B.n386 585
R492 B.n528 B.n343 585
R493 B.n343 B.n342 585
R494 B.n530 B.n529 585
R495 B.n531 B.n530 585
R496 B.n337 B.n336 585
R497 B.n338 B.n337 585
R498 B.n539 B.n538 585
R499 B.n538 B.n537 585
R500 B.n540 B.n335 585
R501 B.n335 B.n333 585
R502 B.n542 B.n541 585
R503 B.n543 B.n542 585
R504 B.n329 B.n328 585
R505 B.n334 B.n329 585
R506 B.n551 B.n550 585
R507 B.n550 B.n549 585
R508 B.n552 B.n327 585
R509 B.n327 B.n326 585
R510 B.n554 B.n553 585
R511 B.n555 B.n554 585
R512 B.n321 B.n320 585
R513 B.n322 B.n321 585
R514 B.n563 B.n562 585
R515 B.n562 B.n561 585
R516 B.n564 B.n319 585
R517 B.n319 B.n318 585
R518 B.n566 B.n565 585
R519 B.n567 B.n566 585
R520 B.n313 B.n312 585
R521 B.n314 B.n313 585
R522 B.n575 B.n574 585
R523 B.n574 B.n573 585
R524 B.n576 B.n311 585
R525 B.n311 B.n310 585
R526 B.n578 B.n577 585
R527 B.n579 B.n578 585
R528 B.n305 B.n304 585
R529 B.n306 B.n305 585
R530 B.n587 B.n586 585
R531 B.n586 B.n585 585
R532 B.n588 B.n303 585
R533 B.n303 B.n302 585
R534 B.n590 B.n589 585
R535 B.n591 B.n590 585
R536 B.n297 B.n296 585
R537 B.n298 B.n297 585
R538 B.n599 B.n598 585
R539 B.n598 B.n597 585
R540 B.n600 B.n295 585
R541 B.n295 B.n294 585
R542 B.n602 B.n601 585
R543 B.n603 B.n602 585
R544 B.n289 B.n288 585
R545 B.n290 B.n289 585
R546 B.n611 B.n610 585
R547 B.n610 B.n609 585
R548 B.n612 B.n287 585
R549 B.n287 B.n286 585
R550 B.n614 B.n613 585
R551 B.n615 B.n614 585
R552 B.n281 B.n280 585
R553 B.n282 B.n281 585
R554 B.n623 B.n622 585
R555 B.n622 B.n621 585
R556 B.n624 B.n279 585
R557 B.n279 B.n278 585
R558 B.n626 B.n625 585
R559 B.n627 B.n626 585
R560 B.n273 B.n272 585
R561 B.n274 B.n273 585
R562 B.n635 B.n634 585
R563 B.n634 B.n633 585
R564 B.n636 B.n271 585
R565 B.n271 B.n269 585
R566 B.n638 B.n637 585
R567 B.n639 B.n638 585
R568 B.n265 B.n264 585
R569 B.n270 B.n265 585
R570 B.n648 B.n647 585
R571 B.n647 B.n646 585
R572 B.n649 B.n263 585
R573 B.n263 B.n262 585
R574 B.n651 B.n650 585
R575 B.n652 B.n651 585
R576 B.n3 B.n0 585
R577 B.n4 B.n3 585
R578 B.n801 B.n1 585
R579 B.n802 B.n801 585
R580 B.n800 B.n799 585
R581 B.n800 B.n8 585
R582 B.n798 B.n9 585
R583 B.n12 B.n9 585
R584 B.n797 B.n796 585
R585 B.n796 B.n795 585
R586 B.n11 B.n10 585
R587 B.n794 B.n11 585
R588 B.n792 B.n791 585
R589 B.n793 B.n792 585
R590 B.n790 B.n17 585
R591 B.n17 B.n16 585
R592 B.n789 B.n788 585
R593 B.n788 B.n787 585
R594 B.n19 B.n18 585
R595 B.n786 B.n19 585
R596 B.n784 B.n783 585
R597 B.n785 B.n784 585
R598 B.n782 B.n24 585
R599 B.n24 B.n23 585
R600 B.n781 B.n780 585
R601 B.n780 B.n779 585
R602 B.n26 B.n25 585
R603 B.n778 B.n26 585
R604 B.n776 B.n775 585
R605 B.n777 B.n776 585
R606 B.n774 B.n31 585
R607 B.n31 B.n30 585
R608 B.n773 B.n772 585
R609 B.n772 B.n771 585
R610 B.n33 B.n32 585
R611 B.n770 B.n33 585
R612 B.n768 B.n767 585
R613 B.n769 B.n768 585
R614 B.n766 B.n38 585
R615 B.n38 B.n37 585
R616 B.n765 B.n764 585
R617 B.n764 B.n763 585
R618 B.n40 B.n39 585
R619 B.n762 B.n40 585
R620 B.n760 B.n759 585
R621 B.n761 B.n760 585
R622 B.n758 B.n45 585
R623 B.n45 B.n44 585
R624 B.n757 B.n756 585
R625 B.n756 B.n755 585
R626 B.n47 B.n46 585
R627 B.n754 B.n47 585
R628 B.n752 B.n751 585
R629 B.n753 B.n752 585
R630 B.n750 B.n52 585
R631 B.n52 B.n51 585
R632 B.n749 B.n748 585
R633 B.n748 B.n747 585
R634 B.n54 B.n53 585
R635 B.n746 B.n54 585
R636 B.n744 B.n743 585
R637 B.n745 B.n744 585
R638 B.n742 B.n59 585
R639 B.n59 B.n58 585
R640 B.n741 B.n740 585
R641 B.n740 B.n739 585
R642 B.n61 B.n60 585
R643 B.n738 B.n61 585
R644 B.n736 B.n735 585
R645 B.n737 B.n736 585
R646 B.n734 B.n66 585
R647 B.n66 B.n65 585
R648 B.n733 B.n732 585
R649 B.n732 B.n731 585
R650 B.n68 B.n67 585
R651 B.n730 B.n68 585
R652 B.n728 B.n727 585
R653 B.n729 B.n728 585
R654 B.n726 B.n73 585
R655 B.n73 B.n72 585
R656 B.n725 B.n724 585
R657 B.n724 B.n723 585
R658 B.n75 B.n74 585
R659 B.n722 B.n75 585
R660 B.n720 B.n719 585
R661 B.n721 B.n720 585
R662 B.n718 B.n80 585
R663 B.n80 B.n79 585
R664 B.n805 B.n804 585
R665 B.n803 B.n2 585
R666 B.n716 B.n80 482.89
R667 B.n713 B.n118 482.89
R668 B.n386 B.n341 482.89
R669 B.n526 B.n343 482.89
R670 B.n122 B.t21 324.113
R671 B.n119 B.t14 324.113
R672 B.n384 B.t10 324.113
R673 B.n381 B.t18 324.113
R674 B.n714 B.n116 256.663
R675 B.n714 B.n115 256.663
R676 B.n714 B.n114 256.663
R677 B.n714 B.n113 256.663
R678 B.n714 B.n112 256.663
R679 B.n714 B.n111 256.663
R680 B.n714 B.n110 256.663
R681 B.n714 B.n109 256.663
R682 B.n714 B.n108 256.663
R683 B.n714 B.n107 256.663
R684 B.n714 B.n106 256.663
R685 B.n714 B.n105 256.663
R686 B.n714 B.n104 256.663
R687 B.n714 B.n103 256.663
R688 B.n714 B.n102 256.663
R689 B.n714 B.n101 256.663
R690 B.n714 B.n100 256.663
R691 B.n714 B.n99 256.663
R692 B.n714 B.n98 256.663
R693 B.n714 B.n97 256.663
R694 B.n714 B.n96 256.663
R695 B.n714 B.n95 256.663
R696 B.n714 B.n94 256.663
R697 B.n714 B.n93 256.663
R698 B.n714 B.n92 256.663
R699 B.n714 B.n91 256.663
R700 B.n714 B.n90 256.663
R701 B.n714 B.n89 256.663
R702 B.n714 B.n88 256.663
R703 B.n714 B.n87 256.663
R704 B.n714 B.n86 256.663
R705 B.n714 B.n85 256.663
R706 B.n714 B.n84 256.663
R707 B.n714 B.n83 256.663
R708 B.n715 B.n714 256.663
R709 B.n525 B.n524 256.663
R710 B.n524 B.n346 256.663
R711 B.n524 B.n347 256.663
R712 B.n524 B.n348 256.663
R713 B.n524 B.n349 256.663
R714 B.n524 B.n350 256.663
R715 B.n524 B.n351 256.663
R716 B.n524 B.n352 256.663
R717 B.n524 B.n353 256.663
R718 B.n524 B.n354 256.663
R719 B.n524 B.n355 256.663
R720 B.n524 B.n356 256.663
R721 B.n524 B.n357 256.663
R722 B.n524 B.n358 256.663
R723 B.n524 B.n359 256.663
R724 B.n524 B.n360 256.663
R725 B.n524 B.n361 256.663
R726 B.n524 B.n362 256.663
R727 B.n524 B.n363 256.663
R728 B.n524 B.n364 256.663
R729 B.n524 B.n365 256.663
R730 B.n524 B.n366 256.663
R731 B.n524 B.n367 256.663
R732 B.n524 B.n368 256.663
R733 B.n524 B.n369 256.663
R734 B.n524 B.n370 256.663
R735 B.n524 B.n371 256.663
R736 B.n524 B.n372 256.663
R737 B.n524 B.n373 256.663
R738 B.n524 B.n374 256.663
R739 B.n524 B.n375 256.663
R740 B.n524 B.n376 256.663
R741 B.n524 B.n377 256.663
R742 B.n524 B.n378 256.663
R743 B.n524 B.n379 256.663
R744 B.n807 B.n806 256.663
R745 B.n124 B.n82 163.367
R746 B.n128 B.n127 163.367
R747 B.n132 B.n131 163.367
R748 B.n136 B.n135 163.367
R749 B.n140 B.n139 163.367
R750 B.n144 B.n143 163.367
R751 B.n148 B.n147 163.367
R752 B.n152 B.n151 163.367
R753 B.n156 B.n155 163.367
R754 B.n160 B.n159 163.367
R755 B.n164 B.n163 163.367
R756 B.n168 B.n167 163.367
R757 B.n172 B.n171 163.367
R758 B.n176 B.n175 163.367
R759 B.n180 B.n179 163.367
R760 B.n185 B.n184 163.367
R761 B.n189 B.n188 163.367
R762 B.n193 B.n192 163.367
R763 B.n197 B.n196 163.367
R764 B.n201 B.n200 163.367
R765 B.n205 B.n204 163.367
R766 B.n209 B.n208 163.367
R767 B.n213 B.n212 163.367
R768 B.n217 B.n216 163.367
R769 B.n221 B.n220 163.367
R770 B.n225 B.n224 163.367
R771 B.n229 B.n228 163.367
R772 B.n233 B.n232 163.367
R773 B.n237 B.n236 163.367
R774 B.n241 B.n240 163.367
R775 B.n245 B.n244 163.367
R776 B.n249 B.n248 163.367
R777 B.n253 B.n252 163.367
R778 B.n257 B.n256 163.367
R779 B.n713 B.n117 163.367
R780 B.n532 B.n341 163.367
R781 B.n532 B.n339 163.367
R782 B.n536 B.n339 163.367
R783 B.n536 B.n332 163.367
R784 B.n544 B.n332 163.367
R785 B.n544 B.n330 163.367
R786 B.n548 B.n330 163.367
R787 B.n548 B.n325 163.367
R788 B.n556 B.n325 163.367
R789 B.n556 B.n323 163.367
R790 B.n560 B.n323 163.367
R791 B.n560 B.n317 163.367
R792 B.n568 B.n317 163.367
R793 B.n568 B.n315 163.367
R794 B.n572 B.n315 163.367
R795 B.n572 B.n309 163.367
R796 B.n580 B.n309 163.367
R797 B.n580 B.n307 163.367
R798 B.n584 B.n307 163.367
R799 B.n584 B.n301 163.367
R800 B.n592 B.n301 163.367
R801 B.n592 B.n299 163.367
R802 B.n596 B.n299 163.367
R803 B.n596 B.n293 163.367
R804 B.n604 B.n293 163.367
R805 B.n604 B.n291 163.367
R806 B.n608 B.n291 163.367
R807 B.n608 B.n285 163.367
R808 B.n616 B.n285 163.367
R809 B.n616 B.n283 163.367
R810 B.n620 B.n283 163.367
R811 B.n620 B.n277 163.367
R812 B.n628 B.n277 163.367
R813 B.n628 B.n275 163.367
R814 B.n632 B.n275 163.367
R815 B.n632 B.n268 163.367
R816 B.n640 B.n268 163.367
R817 B.n640 B.n266 163.367
R818 B.n645 B.n266 163.367
R819 B.n645 B.n261 163.367
R820 B.n653 B.n261 163.367
R821 B.n654 B.n653 163.367
R822 B.n654 B.n5 163.367
R823 B.n6 B.n5 163.367
R824 B.n7 B.n6 163.367
R825 B.n660 B.n7 163.367
R826 B.n661 B.n660 163.367
R827 B.n661 B.n13 163.367
R828 B.n14 B.n13 163.367
R829 B.n15 B.n14 163.367
R830 B.n666 B.n15 163.367
R831 B.n666 B.n20 163.367
R832 B.n21 B.n20 163.367
R833 B.n22 B.n21 163.367
R834 B.n671 B.n22 163.367
R835 B.n671 B.n27 163.367
R836 B.n28 B.n27 163.367
R837 B.n29 B.n28 163.367
R838 B.n676 B.n29 163.367
R839 B.n676 B.n34 163.367
R840 B.n35 B.n34 163.367
R841 B.n36 B.n35 163.367
R842 B.n681 B.n36 163.367
R843 B.n681 B.n41 163.367
R844 B.n42 B.n41 163.367
R845 B.n43 B.n42 163.367
R846 B.n686 B.n43 163.367
R847 B.n686 B.n48 163.367
R848 B.n49 B.n48 163.367
R849 B.n50 B.n49 163.367
R850 B.n691 B.n50 163.367
R851 B.n691 B.n55 163.367
R852 B.n56 B.n55 163.367
R853 B.n57 B.n56 163.367
R854 B.n696 B.n57 163.367
R855 B.n696 B.n62 163.367
R856 B.n63 B.n62 163.367
R857 B.n64 B.n63 163.367
R858 B.n701 B.n64 163.367
R859 B.n701 B.n69 163.367
R860 B.n70 B.n69 163.367
R861 B.n71 B.n70 163.367
R862 B.n706 B.n71 163.367
R863 B.n706 B.n76 163.367
R864 B.n77 B.n76 163.367
R865 B.n78 B.n77 163.367
R866 B.n118 B.n78 163.367
R867 B.n523 B.n345 163.367
R868 B.n523 B.n380 163.367
R869 B.n519 B.n518 163.367
R870 B.n515 B.n514 163.367
R871 B.n511 B.n510 163.367
R872 B.n507 B.n506 163.367
R873 B.n503 B.n502 163.367
R874 B.n499 B.n498 163.367
R875 B.n495 B.n494 163.367
R876 B.n491 B.n490 163.367
R877 B.n487 B.n486 163.367
R878 B.n483 B.n482 163.367
R879 B.n479 B.n478 163.367
R880 B.n475 B.n474 163.367
R881 B.n471 B.n470 163.367
R882 B.n467 B.n466 163.367
R883 B.n463 B.n462 163.367
R884 B.n459 B.n458 163.367
R885 B.n455 B.n454 163.367
R886 B.n451 B.n450 163.367
R887 B.n446 B.n445 163.367
R888 B.n442 B.n441 163.367
R889 B.n438 B.n437 163.367
R890 B.n434 B.n433 163.367
R891 B.n430 B.n429 163.367
R892 B.n426 B.n425 163.367
R893 B.n422 B.n421 163.367
R894 B.n418 B.n417 163.367
R895 B.n414 B.n413 163.367
R896 B.n410 B.n409 163.367
R897 B.n406 B.n405 163.367
R898 B.n402 B.n401 163.367
R899 B.n398 B.n397 163.367
R900 B.n394 B.n393 163.367
R901 B.n390 B.n389 163.367
R902 B.n530 B.n343 163.367
R903 B.n530 B.n337 163.367
R904 B.n538 B.n337 163.367
R905 B.n538 B.n335 163.367
R906 B.n542 B.n335 163.367
R907 B.n542 B.n329 163.367
R908 B.n550 B.n329 163.367
R909 B.n550 B.n327 163.367
R910 B.n554 B.n327 163.367
R911 B.n554 B.n321 163.367
R912 B.n562 B.n321 163.367
R913 B.n562 B.n319 163.367
R914 B.n566 B.n319 163.367
R915 B.n566 B.n313 163.367
R916 B.n574 B.n313 163.367
R917 B.n574 B.n311 163.367
R918 B.n578 B.n311 163.367
R919 B.n578 B.n305 163.367
R920 B.n586 B.n305 163.367
R921 B.n586 B.n303 163.367
R922 B.n590 B.n303 163.367
R923 B.n590 B.n297 163.367
R924 B.n598 B.n297 163.367
R925 B.n598 B.n295 163.367
R926 B.n602 B.n295 163.367
R927 B.n602 B.n289 163.367
R928 B.n610 B.n289 163.367
R929 B.n610 B.n287 163.367
R930 B.n614 B.n287 163.367
R931 B.n614 B.n281 163.367
R932 B.n622 B.n281 163.367
R933 B.n622 B.n279 163.367
R934 B.n626 B.n279 163.367
R935 B.n626 B.n273 163.367
R936 B.n634 B.n273 163.367
R937 B.n634 B.n271 163.367
R938 B.n638 B.n271 163.367
R939 B.n638 B.n265 163.367
R940 B.n647 B.n265 163.367
R941 B.n647 B.n263 163.367
R942 B.n651 B.n263 163.367
R943 B.n651 B.n3 163.367
R944 B.n805 B.n3 163.367
R945 B.n801 B.n2 163.367
R946 B.n801 B.n800 163.367
R947 B.n800 B.n9 163.367
R948 B.n796 B.n9 163.367
R949 B.n796 B.n11 163.367
R950 B.n792 B.n11 163.367
R951 B.n792 B.n17 163.367
R952 B.n788 B.n17 163.367
R953 B.n788 B.n19 163.367
R954 B.n784 B.n19 163.367
R955 B.n784 B.n24 163.367
R956 B.n780 B.n24 163.367
R957 B.n780 B.n26 163.367
R958 B.n776 B.n26 163.367
R959 B.n776 B.n31 163.367
R960 B.n772 B.n31 163.367
R961 B.n772 B.n33 163.367
R962 B.n768 B.n33 163.367
R963 B.n768 B.n38 163.367
R964 B.n764 B.n38 163.367
R965 B.n764 B.n40 163.367
R966 B.n760 B.n40 163.367
R967 B.n760 B.n45 163.367
R968 B.n756 B.n45 163.367
R969 B.n756 B.n47 163.367
R970 B.n752 B.n47 163.367
R971 B.n752 B.n52 163.367
R972 B.n748 B.n52 163.367
R973 B.n748 B.n54 163.367
R974 B.n744 B.n54 163.367
R975 B.n744 B.n59 163.367
R976 B.n740 B.n59 163.367
R977 B.n740 B.n61 163.367
R978 B.n736 B.n61 163.367
R979 B.n736 B.n66 163.367
R980 B.n732 B.n66 163.367
R981 B.n732 B.n68 163.367
R982 B.n728 B.n68 163.367
R983 B.n728 B.n73 163.367
R984 B.n724 B.n73 163.367
R985 B.n724 B.n75 163.367
R986 B.n720 B.n75 163.367
R987 B.n720 B.n80 163.367
R988 B.n119 B.t16 108.88
R989 B.n384 B.t13 108.88
R990 B.n122 B.t22 108.871
R991 B.n381 B.t20 108.871
R992 B.n524 B.n342 105.073
R993 B.n714 B.n79 105.073
R994 B.n716 B.n715 71.676
R995 B.n124 B.n83 71.676
R996 B.n128 B.n84 71.676
R997 B.n132 B.n85 71.676
R998 B.n136 B.n86 71.676
R999 B.n140 B.n87 71.676
R1000 B.n144 B.n88 71.676
R1001 B.n148 B.n89 71.676
R1002 B.n152 B.n90 71.676
R1003 B.n156 B.n91 71.676
R1004 B.n160 B.n92 71.676
R1005 B.n164 B.n93 71.676
R1006 B.n168 B.n94 71.676
R1007 B.n172 B.n95 71.676
R1008 B.n176 B.n96 71.676
R1009 B.n180 B.n97 71.676
R1010 B.n185 B.n98 71.676
R1011 B.n189 B.n99 71.676
R1012 B.n193 B.n100 71.676
R1013 B.n197 B.n101 71.676
R1014 B.n201 B.n102 71.676
R1015 B.n205 B.n103 71.676
R1016 B.n209 B.n104 71.676
R1017 B.n213 B.n105 71.676
R1018 B.n217 B.n106 71.676
R1019 B.n221 B.n107 71.676
R1020 B.n225 B.n108 71.676
R1021 B.n229 B.n109 71.676
R1022 B.n233 B.n110 71.676
R1023 B.n237 B.n111 71.676
R1024 B.n241 B.n112 71.676
R1025 B.n245 B.n113 71.676
R1026 B.n249 B.n114 71.676
R1027 B.n253 B.n115 71.676
R1028 B.n257 B.n116 71.676
R1029 B.n117 B.n116 71.676
R1030 B.n256 B.n115 71.676
R1031 B.n252 B.n114 71.676
R1032 B.n248 B.n113 71.676
R1033 B.n244 B.n112 71.676
R1034 B.n240 B.n111 71.676
R1035 B.n236 B.n110 71.676
R1036 B.n232 B.n109 71.676
R1037 B.n228 B.n108 71.676
R1038 B.n224 B.n107 71.676
R1039 B.n220 B.n106 71.676
R1040 B.n216 B.n105 71.676
R1041 B.n212 B.n104 71.676
R1042 B.n208 B.n103 71.676
R1043 B.n204 B.n102 71.676
R1044 B.n200 B.n101 71.676
R1045 B.n196 B.n100 71.676
R1046 B.n192 B.n99 71.676
R1047 B.n188 B.n98 71.676
R1048 B.n184 B.n97 71.676
R1049 B.n179 B.n96 71.676
R1050 B.n175 B.n95 71.676
R1051 B.n171 B.n94 71.676
R1052 B.n167 B.n93 71.676
R1053 B.n163 B.n92 71.676
R1054 B.n159 B.n91 71.676
R1055 B.n155 B.n90 71.676
R1056 B.n151 B.n89 71.676
R1057 B.n147 B.n88 71.676
R1058 B.n143 B.n87 71.676
R1059 B.n139 B.n86 71.676
R1060 B.n135 B.n85 71.676
R1061 B.n131 B.n84 71.676
R1062 B.n127 B.n83 71.676
R1063 B.n715 B.n82 71.676
R1064 B.n526 B.n525 71.676
R1065 B.n380 B.n346 71.676
R1066 B.n518 B.n347 71.676
R1067 B.n514 B.n348 71.676
R1068 B.n510 B.n349 71.676
R1069 B.n506 B.n350 71.676
R1070 B.n502 B.n351 71.676
R1071 B.n498 B.n352 71.676
R1072 B.n494 B.n353 71.676
R1073 B.n490 B.n354 71.676
R1074 B.n486 B.n355 71.676
R1075 B.n482 B.n356 71.676
R1076 B.n478 B.n357 71.676
R1077 B.n474 B.n358 71.676
R1078 B.n470 B.n359 71.676
R1079 B.n466 B.n360 71.676
R1080 B.n462 B.n361 71.676
R1081 B.n458 B.n362 71.676
R1082 B.n454 B.n363 71.676
R1083 B.n450 B.n364 71.676
R1084 B.n445 B.n365 71.676
R1085 B.n441 B.n366 71.676
R1086 B.n437 B.n367 71.676
R1087 B.n433 B.n368 71.676
R1088 B.n429 B.n369 71.676
R1089 B.n425 B.n370 71.676
R1090 B.n421 B.n371 71.676
R1091 B.n417 B.n372 71.676
R1092 B.n413 B.n373 71.676
R1093 B.n409 B.n374 71.676
R1094 B.n405 B.n375 71.676
R1095 B.n401 B.n376 71.676
R1096 B.n397 B.n377 71.676
R1097 B.n393 B.n378 71.676
R1098 B.n389 B.n379 71.676
R1099 B.n525 B.n345 71.676
R1100 B.n519 B.n346 71.676
R1101 B.n515 B.n347 71.676
R1102 B.n511 B.n348 71.676
R1103 B.n507 B.n349 71.676
R1104 B.n503 B.n350 71.676
R1105 B.n499 B.n351 71.676
R1106 B.n495 B.n352 71.676
R1107 B.n491 B.n353 71.676
R1108 B.n487 B.n354 71.676
R1109 B.n483 B.n355 71.676
R1110 B.n479 B.n356 71.676
R1111 B.n475 B.n357 71.676
R1112 B.n471 B.n358 71.676
R1113 B.n467 B.n359 71.676
R1114 B.n463 B.n360 71.676
R1115 B.n459 B.n361 71.676
R1116 B.n455 B.n362 71.676
R1117 B.n451 B.n363 71.676
R1118 B.n446 B.n364 71.676
R1119 B.n442 B.n365 71.676
R1120 B.n438 B.n366 71.676
R1121 B.n434 B.n367 71.676
R1122 B.n430 B.n368 71.676
R1123 B.n426 B.n369 71.676
R1124 B.n422 B.n370 71.676
R1125 B.n418 B.n371 71.676
R1126 B.n414 B.n372 71.676
R1127 B.n410 B.n373 71.676
R1128 B.n406 B.n374 71.676
R1129 B.n402 B.n375 71.676
R1130 B.n398 B.n376 71.676
R1131 B.n394 B.n377 71.676
R1132 B.n390 B.n378 71.676
R1133 B.n386 B.n379 71.676
R1134 B.n806 B.n805 71.676
R1135 B.n806 B.n2 71.676
R1136 B.n120 B.t17 69.8983
R1137 B.n385 B.t12 69.8983
R1138 B.n123 B.t23 69.8885
R1139 B.n382 B.t19 69.8885
R1140 B.n182 B.n123 59.5399
R1141 B.n121 B.n120 59.5399
R1142 B.n448 B.n385 59.5399
R1143 B.n383 B.n382 59.5399
R1144 B.n531 B.n342 55.3874
R1145 B.n531 B.n338 55.3874
R1146 B.n537 B.n338 55.3874
R1147 B.n537 B.n333 55.3874
R1148 B.n543 B.n333 55.3874
R1149 B.n543 B.n334 55.3874
R1150 B.n549 B.n326 55.3874
R1151 B.n555 B.n326 55.3874
R1152 B.n555 B.n322 55.3874
R1153 B.n561 B.n322 55.3874
R1154 B.n561 B.n318 55.3874
R1155 B.n567 B.n318 55.3874
R1156 B.n567 B.n314 55.3874
R1157 B.n573 B.n314 55.3874
R1158 B.n579 B.n310 55.3874
R1159 B.n579 B.n306 55.3874
R1160 B.n585 B.n306 55.3874
R1161 B.n585 B.n302 55.3874
R1162 B.n591 B.n302 55.3874
R1163 B.n597 B.n298 55.3874
R1164 B.n597 B.n294 55.3874
R1165 B.n603 B.n294 55.3874
R1166 B.n603 B.n290 55.3874
R1167 B.n609 B.n290 55.3874
R1168 B.n615 B.n286 55.3874
R1169 B.n615 B.n282 55.3874
R1170 B.n621 B.n282 55.3874
R1171 B.n621 B.n278 55.3874
R1172 B.n627 B.n278 55.3874
R1173 B.n633 B.n274 55.3874
R1174 B.n633 B.n269 55.3874
R1175 B.n639 B.n269 55.3874
R1176 B.n639 B.n270 55.3874
R1177 B.n646 B.n262 55.3874
R1178 B.n652 B.n262 55.3874
R1179 B.n652 B.n4 55.3874
R1180 B.n804 B.n4 55.3874
R1181 B.n804 B.n803 55.3874
R1182 B.n803 B.n802 55.3874
R1183 B.n802 B.n8 55.3874
R1184 B.n12 B.n8 55.3874
R1185 B.n795 B.n12 55.3874
R1186 B.n794 B.n793 55.3874
R1187 B.n793 B.n16 55.3874
R1188 B.n787 B.n16 55.3874
R1189 B.n787 B.n786 55.3874
R1190 B.n785 B.n23 55.3874
R1191 B.n779 B.n23 55.3874
R1192 B.n779 B.n778 55.3874
R1193 B.n778 B.n777 55.3874
R1194 B.n777 B.n30 55.3874
R1195 B.n771 B.n770 55.3874
R1196 B.n770 B.n769 55.3874
R1197 B.n769 B.n37 55.3874
R1198 B.n763 B.n37 55.3874
R1199 B.n763 B.n762 55.3874
R1200 B.n761 B.n44 55.3874
R1201 B.n755 B.n44 55.3874
R1202 B.n755 B.n754 55.3874
R1203 B.n754 B.n753 55.3874
R1204 B.n753 B.n51 55.3874
R1205 B.n747 B.n746 55.3874
R1206 B.n746 B.n745 55.3874
R1207 B.n745 B.n58 55.3874
R1208 B.n739 B.n58 55.3874
R1209 B.n739 B.n738 55.3874
R1210 B.n738 B.n737 55.3874
R1211 B.n737 B.n65 55.3874
R1212 B.n731 B.n65 55.3874
R1213 B.n730 B.n729 55.3874
R1214 B.n729 B.n72 55.3874
R1215 B.n723 B.n72 55.3874
R1216 B.n723 B.n722 55.3874
R1217 B.n722 B.n721 55.3874
R1218 B.n721 B.n79 55.3874
R1219 B.t7 B.n274 53.7584
R1220 B.n786 B.t3 53.7584
R1221 B.n270 B.t5 52.1293
R1222 B.t8 B.n794 52.1293
R1223 B.t9 B.n286 48.8713
R1224 B.t4 B.n30 48.8713
R1225 B.n549 B.t11 45.6132
R1226 B.n731 B.t15 45.6132
R1227 B.t1 B.n298 43.9842
R1228 B.n762 B.t0 43.9842
R1229 B.t2 B.n310 39.0971
R1230 B.t6 B.n51 39.0971
R1231 B.n123 B.n122 38.9823
R1232 B.n120 B.n119 38.9823
R1233 B.n385 B.n384 38.9823
R1234 B.n382 B.n381 38.9823
R1235 B.n528 B.n527 31.3761
R1236 B.n387 B.n340 31.3761
R1237 B.n712 B.n711 31.3761
R1238 B.n718 B.n717 31.3761
R1239 B B.n807 18.0485
R1240 B.n573 B.t2 16.2908
R1241 B.n747 B.t6 16.2908
R1242 B.n591 B.t1 11.4037
R1243 B.t0 B.n761 11.4037
R1244 B.n529 B.n528 10.6151
R1245 B.n529 B.n336 10.6151
R1246 B.n539 B.n336 10.6151
R1247 B.n540 B.n539 10.6151
R1248 B.n541 B.n540 10.6151
R1249 B.n541 B.n328 10.6151
R1250 B.n551 B.n328 10.6151
R1251 B.n552 B.n551 10.6151
R1252 B.n553 B.n552 10.6151
R1253 B.n553 B.n320 10.6151
R1254 B.n563 B.n320 10.6151
R1255 B.n564 B.n563 10.6151
R1256 B.n565 B.n564 10.6151
R1257 B.n565 B.n312 10.6151
R1258 B.n575 B.n312 10.6151
R1259 B.n576 B.n575 10.6151
R1260 B.n577 B.n576 10.6151
R1261 B.n577 B.n304 10.6151
R1262 B.n587 B.n304 10.6151
R1263 B.n588 B.n587 10.6151
R1264 B.n589 B.n588 10.6151
R1265 B.n589 B.n296 10.6151
R1266 B.n599 B.n296 10.6151
R1267 B.n600 B.n599 10.6151
R1268 B.n601 B.n600 10.6151
R1269 B.n601 B.n288 10.6151
R1270 B.n611 B.n288 10.6151
R1271 B.n612 B.n611 10.6151
R1272 B.n613 B.n612 10.6151
R1273 B.n613 B.n280 10.6151
R1274 B.n623 B.n280 10.6151
R1275 B.n624 B.n623 10.6151
R1276 B.n625 B.n624 10.6151
R1277 B.n625 B.n272 10.6151
R1278 B.n635 B.n272 10.6151
R1279 B.n636 B.n635 10.6151
R1280 B.n637 B.n636 10.6151
R1281 B.n637 B.n264 10.6151
R1282 B.n648 B.n264 10.6151
R1283 B.n649 B.n648 10.6151
R1284 B.n650 B.n649 10.6151
R1285 B.n650 B.n0 10.6151
R1286 B.n527 B.n344 10.6151
R1287 B.n522 B.n344 10.6151
R1288 B.n522 B.n521 10.6151
R1289 B.n521 B.n520 10.6151
R1290 B.n520 B.n517 10.6151
R1291 B.n517 B.n516 10.6151
R1292 B.n516 B.n513 10.6151
R1293 B.n513 B.n512 10.6151
R1294 B.n512 B.n509 10.6151
R1295 B.n509 B.n508 10.6151
R1296 B.n508 B.n505 10.6151
R1297 B.n505 B.n504 10.6151
R1298 B.n504 B.n501 10.6151
R1299 B.n501 B.n500 10.6151
R1300 B.n500 B.n497 10.6151
R1301 B.n497 B.n496 10.6151
R1302 B.n496 B.n493 10.6151
R1303 B.n493 B.n492 10.6151
R1304 B.n492 B.n489 10.6151
R1305 B.n489 B.n488 10.6151
R1306 B.n488 B.n485 10.6151
R1307 B.n485 B.n484 10.6151
R1308 B.n484 B.n481 10.6151
R1309 B.n481 B.n480 10.6151
R1310 B.n480 B.n477 10.6151
R1311 B.n477 B.n476 10.6151
R1312 B.n476 B.n473 10.6151
R1313 B.n473 B.n472 10.6151
R1314 B.n472 B.n469 10.6151
R1315 B.n469 B.n468 10.6151
R1316 B.n465 B.n464 10.6151
R1317 B.n464 B.n461 10.6151
R1318 B.n461 B.n460 10.6151
R1319 B.n460 B.n457 10.6151
R1320 B.n457 B.n456 10.6151
R1321 B.n456 B.n453 10.6151
R1322 B.n453 B.n452 10.6151
R1323 B.n452 B.n449 10.6151
R1324 B.n447 B.n444 10.6151
R1325 B.n444 B.n443 10.6151
R1326 B.n443 B.n440 10.6151
R1327 B.n440 B.n439 10.6151
R1328 B.n439 B.n436 10.6151
R1329 B.n436 B.n435 10.6151
R1330 B.n435 B.n432 10.6151
R1331 B.n432 B.n431 10.6151
R1332 B.n431 B.n428 10.6151
R1333 B.n428 B.n427 10.6151
R1334 B.n427 B.n424 10.6151
R1335 B.n424 B.n423 10.6151
R1336 B.n423 B.n420 10.6151
R1337 B.n420 B.n419 10.6151
R1338 B.n419 B.n416 10.6151
R1339 B.n416 B.n415 10.6151
R1340 B.n415 B.n412 10.6151
R1341 B.n412 B.n411 10.6151
R1342 B.n411 B.n408 10.6151
R1343 B.n408 B.n407 10.6151
R1344 B.n407 B.n404 10.6151
R1345 B.n404 B.n403 10.6151
R1346 B.n403 B.n400 10.6151
R1347 B.n400 B.n399 10.6151
R1348 B.n399 B.n396 10.6151
R1349 B.n396 B.n395 10.6151
R1350 B.n395 B.n392 10.6151
R1351 B.n392 B.n391 10.6151
R1352 B.n391 B.n388 10.6151
R1353 B.n388 B.n387 10.6151
R1354 B.n533 B.n340 10.6151
R1355 B.n534 B.n533 10.6151
R1356 B.n535 B.n534 10.6151
R1357 B.n535 B.n331 10.6151
R1358 B.n545 B.n331 10.6151
R1359 B.n546 B.n545 10.6151
R1360 B.n547 B.n546 10.6151
R1361 B.n547 B.n324 10.6151
R1362 B.n557 B.n324 10.6151
R1363 B.n558 B.n557 10.6151
R1364 B.n559 B.n558 10.6151
R1365 B.n559 B.n316 10.6151
R1366 B.n569 B.n316 10.6151
R1367 B.n570 B.n569 10.6151
R1368 B.n571 B.n570 10.6151
R1369 B.n571 B.n308 10.6151
R1370 B.n581 B.n308 10.6151
R1371 B.n582 B.n581 10.6151
R1372 B.n583 B.n582 10.6151
R1373 B.n583 B.n300 10.6151
R1374 B.n593 B.n300 10.6151
R1375 B.n594 B.n593 10.6151
R1376 B.n595 B.n594 10.6151
R1377 B.n595 B.n292 10.6151
R1378 B.n605 B.n292 10.6151
R1379 B.n606 B.n605 10.6151
R1380 B.n607 B.n606 10.6151
R1381 B.n607 B.n284 10.6151
R1382 B.n617 B.n284 10.6151
R1383 B.n618 B.n617 10.6151
R1384 B.n619 B.n618 10.6151
R1385 B.n619 B.n276 10.6151
R1386 B.n629 B.n276 10.6151
R1387 B.n630 B.n629 10.6151
R1388 B.n631 B.n630 10.6151
R1389 B.n631 B.n267 10.6151
R1390 B.n641 B.n267 10.6151
R1391 B.n642 B.n641 10.6151
R1392 B.n644 B.n642 10.6151
R1393 B.n644 B.n643 10.6151
R1394 B.n643 B.n260 10.6151
R1395 B.n655 B.n260 10.6151
R1396 B.n656 B.n655 10.6151
R1397 B.n657 B.n656 10.6151
R1398 B.n658 B.n657 10.6151
R1399 B.n659 B.n658 10.6151
R1400 B.n662 B.n659 10.6151
R1401 B.n663 B.n662 10.6151
R1402 B.n664 B.n663 10.6151
R1403 B.n665 B.n664 10.6151
R1404 B.n667 B.n665 10.6151
R1405 B.n668 B.n667 10.6151
R1406 B.n669 B.n668 10.6151
R1407 B.n670 B.n669 10.6151
R1408 B.n672 B.n670 10.6151
R1409 B.n673 B.n672 10.6151
R1410 B.n674 B.n673 10.6151
R1411 B.n675 B.n674 10.6151
R1412 B.n677 B.n675 10.6151
R1413 B.n678 B.n677 10.6151
R1414 B.n679 B.n678 10.6151
R1415 B.n680 B.n679 10.6151
R1416 B.n682 B.n680 10.6151
R1417 B.n683 B.n682 10.6151
R1418 B.n684 B.n683 10.6151
R1419 B.n685 B.n684 10.6151
R1420 B.n687 B.n685 10.6151
R1421 B.n688 B.n687 10.6151
R1422 B.n689 B.n688 10.6151
R1423 B.n690 B.n689 10.6151
R1424 B.n692 B.n690 10.6151
R1425 B.n693 B.n692 10.6151
R1426 B.n694 B.n693 10.6151
R1427 B.n695 B.n694 10.6151
R1428 B.n697 B.n695 10.6151
R1429 B.n698 B.n697 10.6151
R1430 B.n699 B.n698 10.6151
R1431 B.n700 B.n699 10.6151
R1432 B.n702 B.n700 10.6151
R1433 B.n703 B.n702 10.6151
R1434 B.n704 B.n703 10.6151
R1435 B.n705 B.n704 10.6151
R1436 B.n707 B.n705 10.6151
R1437 B.n708 B.n707 10.6151
R1438 B.n709 B.n708 10.6151
R1439 B.n710 B.n709 10.6151
R1440 B.n711 B.n710 10.6151
R1441 B.n799 B.n1 10.6151
R1442 B.n799 B.n798 10.6151
R1443 B.n798 B.n797 10.6151
R1444 B.n797 B.n10 10.6151
R1445 B.n791 B.n10 10.6151
R1446 B.n791 B.n790 10.6151
R1447 B.n790 B.n789 10.6151
R1448 B.n789 B.n18 10.6151
R1449 B.n783 B.n18 10.6151
R1450 B.n783 B.n782 10.6151
R1451 B.n782 B.n781 10.6151
R1452 B.n781 B.n25 10.6151
R1453 B.n775 B.n25 10.6151
R1454 B.n775 B.n774 10.6151
R1455 B.n774 B.n773 10.6151
R1456 B.n773 B.n32 10.6151
R1457 B.n767 B.n32 10.6151
R1458 B.n767 B.n766 10.6151
R1459 B.n766 B.n765 10.6151
R1460 B.n765 B.n39 10.6151
R1461 B.n759 B.n39 10.6151
R1462 B.n759 B.n758 10.6151
R1463 B.n758 B.n757 10.6151
R1464 B.n757 B.n46 10.6151
R1465 B.n751 B.n46 10.6151
R1466 B.n751 B.n750 10.6151
R1467 B.n750 B.n749 10.6151
R1468 B.n749 B.n53 10.6151
R1469 B.n743 B.n53 10.6151
R1470 B.n743 B.n742 10.6151
R1471 B.n742 B.n741 10.6151
R1472 B.n741 B.n60 10.6151
R1473 B.n735 B.n60 10.6151
R1474 B.n735 B.n734 10.6151
R1475 B.n734 B.n733 10.6151
R1476 B.n733 B.n67 10.6151
R1477 B.n727 B.n67 10.6151
R1478 B.n727 B.n726 10.6151
R1479 B.n726 B.n725 10.6151
R1480 B.n725 B.n74 10.6151
R1481 B.n719 B.n74 10.6151
R1482 B.n719 B.n718 10.6151
R1483 B.n717 B.n81 10.6151
R1484 B.n125 B.n81 10.6151
R1485 B.n126 B.n125 10.6151
R1486 B.n129 B.n126 10.6151
R1487 B.n130 B.n129 10.6151
R1488 B.n133 B.n130 10.6151
R1489 B.n134 B.n133 10.6151
R1490 B.n137 B.n134 10.6151
R1491 B.n138 B.n137 10.6151
R1492 B.n141 B.n138 10.6151
R1493 B.n142 B.n141 10.6151
R1494 B.n145 B.n142 10.6151
R1495 B.n146 B.n145 10.6151
R1496 B.n149 B.n146 10.6151
R1497 B.n150 B.n149 10.6151
R1498 B.n153 B.n150 10.6151
R1499 B.n154 B.n153 10.6151
R1500 B.n157 B.n154 10.6151
R1501 B.n158 B.n157 10.6151
R1502 B.n161 B.n158 10.6151
R1503 B.n162 B.n161 10.6151
R1504 B.n165 B.n162 10.6151
R1505 B.n166 B.n165 10.6151
R1506 B.n169 B.n166 10.6151
R1507 B.n170 B.n169 10.6151
R1508 B.n173 B.n170 10.6151
R1509 B.n174 B.n173 10.6151
R1510 B.n177 B.n174 10.6151
R1511 B.n178 B.n177 10.6151
R1512 B.n181 B.n178 10.6151
R1513 B.n186 B.n183 10.6151
R1514 B.n187 B.n186 10.6151
R1515 B.n190 B.n187 10.6151
R1516 B.n191 B.n190 10.6151
R1517 B.n194 B.n191 10.6151
R1518 B.n195 B.n194 10.6151
R1519 B.n198 B.n195 10.6151
R1520 B.n199 B.n198 10.6151
R1521 B.n203 B.n202 10.6151
R1522 B.n206 B.n203 10.6151
R1523 B.n207 B.n206 10.6151
R1524 B.n210 B.n207 10.6151
R1525 B.n211 B.n210 10.6151
R1526 B.n214 B.n211 10.6151
R1527 B.n215 B.n214 10.6151
R1528 B.n218 B.n215 10.6151
R1529 B.n219 B.n218 10.6151
R1530 B.n222 B.n219 10.6151
R1531 B.n223 B.n222 10.6151
R1532 B.n226 B.n223 10.6151
R1533 B.n227 B.n226 10.6151
R1534 B.n230 B.n227 10.6151
R1535 B.n231 B.n230 10.6151
R1536 B.n234 B.n231 10.6151
R1537 B.n235 B.n234 10.6151
R1538 B.n238 B.n235 10.6151
R1539 B.n239 B.n238 10.6151
R1540 B.n242 B.n239 10.6151
R1541 B.n243 B.n242 10.6151
R1542 B.n246 B.n243 10.6151
R1543 B.n247 B.n246 10.6151
R1544 B.n250 B.n247 10.6151
R1545 B.n251 B.n250 10.6151
R1546 B.n254 B.n251 10.6151
R1547 B.n255 B.n254 10.6151
R1548 B.n258 B.n255 10.6151
R1549 B.n259 B.n258 10.6151
R1550 B.n712 B.n259 10.6151
R1551 B.n334 B.t11 9.77466
R1552 B.t15 B.n730 9.77466
R1553 B.n807 B.n0 8.11757
R1554 B.n807 B.n1 8.11757
R1555 B.n465 B.n383 6.5566
R1556 B.n449 B.n448 6.5566
R1557 B.n183 B.n182 6.5566
R1558 B.n199 B.n121 6.5566
R1559 B.n609 B.t9 6.51661
R1560 B.n771 B.t4 6.51661
R1561 B.n468 B.n383 4.05904
R1562 B.n448 B.n447 4.05904
R1563 B.n182 B.n181 4.05904
R1564 B.n202 B.n121 4.05904
R1565 B.n646 B.t5 3.25855
R1566 B.n795 B.t8 3.25855
R1567 B.n627 B.t7 1.62953
R1568 B.t3 B.n785 1.62953
R1569 VN.n30 VN.n29 184.788
R1570 VN.n61 VN.n60 184.788
R1571 VN.n59 VN.n31 161.3
R1572 VN.n58 VN.n57 161.3
R1573 VN.n56 VN.n32 161.3
R1574 VN.n55 VN.n54 161.3
R1575 VN.n52 VN.n33 161.3
R1576 VN.n51 VN.n50 161.3
R1577 VN.n49 VN.n34 161.3
R1578 VN.n48 VN.n47 161.3
R1579 VN.n46 VN.n35 161.3
R1580 VN.n45 VN.n44 161.3
R1581 VN.n43 VN.n36 161.3
R1582 VN.n42 VN.n41 161.3
R1583 VN.n40 VN.n37 161.3
R1584 VN.n28 VN.n0 161.3
R1585 VN.n27 VN.n26 161.3
R1586 VN.n25 VN.n1 161.3
R1587 VN.n24 VN.n23 161.3
R1588 VN.n21 VN.n2 161.3
R1589 VN.n20 VN.n19 161.3
R1590 VN.n18 VN.n3 161.3
R1591 VN.n17 VN.n16 161.3
R1592 VN.n15 VN.n4 161.3
R1593 VN.n14 VN.n13 161.3
R1594 VN.n12 VN.n5 161.3
R1595 VN.n11 VN.n10 161.3
R1596 VN.n9 VN.n6 161.3
R1597 VN.n7 VN.t6 145.749
R1598 VN.n38 VN.t5 145.749
R1599 VN.n15 VN.t3 118.061
R1600 VN.n8 VN.t7 118.061
R1601 VN.n22 VN.t4 118.061
R1602 VN.n29 VN.t2 118.061
R1603 VN.n46 VN.t9 118.061
R1604 VN.n39 VN.t8 118.061
R1605 VN.n53 VN.t0 118.061
R1606 VN.n60 VN.t1 118.061
R1607 VN.n8 VN.n7 68.3921
R1608 VN.n39 VN.n38 68.3921
R1609 VN VN.n61 45.4683
R1610 VN.n27 VN.n1 41.9503
R1611 VN.n58 VN.n32 41.9503
R1612 VN.n10 VN.n5 40.979
R1613 VN.n20 VN.n3 40.979
R1614 VN.n41 VN.n36 40.979
R1615 VN.n51 VN.n34 40.979
R1616 VN.n14 VN.n5 40.0078
R1617 VN.n16 VN.n3 40.0078
R1618 VN.n45 VN.n36 40.0078
R1619 VN.n47 VN.n34 40.0078
R1620 VN.n23 VN.n1 39.0365
R1621 VN.n54 VN.n32 39.0365
R1622 VN.n10 VN.n9 24.4675
R1623 VN.n15 VN.n14 24.4675
R1624 VN.n16 VN.n15 24.4675
R1625 VN.n21 VN.n20 24.4675
R1626 VN.n28 VN.n27 24.4675
R1627 VN.n41 VN.n40 24.4675
R1628 VN.n47 VN.n46 24.4675
R1629 VN.n46 VN.n45 24.4675
R1630 VN.n52 VN.n51 24.4675
R1631 VN.n59 VN.n58 24.4675
R1632 VN.n23 VN.n22 23.9782
R1633 VN.n54 VN.n53 23.9782
R1634 VN.n38 VN.n37 18.9635
R1635 VN.n7 VN.n6 18.9635
R1636 VN.n29 VN.n28 0.97918
R1637 VN.n60 VN.n59 0.97918
R1638 VN.n9 VN.n8 0.48984
R1639 VN.n22 VN.n21 0.48984
R1640 VN.n40 VN.n39 0.48984
R1641 VN.n53 VN.n52 0.48984
R1642 VN.n61 VN.n31 0.189894
R1643 VN.n57 VN.n31 0.189894
R1644 VN.n57 VN.n56 0.189894
R1645 VN.n56 VN.n55 0.189894
R1646 VN.n55 VN.n33 0.189894
R1647 VN.n50 VN.n33 0.189894
R1648 VN.n50 VN.n49 0.189894
R1649 VN.n49 VN.n48 0.189894
R1650 VN.n48 VN.n35 0.189894
R1651 VN.n44 VN.n35 0.189894
R1652 VN.n44 VN.n43 0.189894
R1653 VN.n43 VN.n42 0.189894
R1654 VN.n42 VN.n37 0.189894
R1655 VN.n11 VN.n6 0.189894
R1656 VN.n12 VN.n11 0.189894
R1657 VN.n13 VN.n12 0.189894
R1658 VN.n13 VN.n4 0.189894
R1659 VN.n17 VN.n4 0.189894
R1660 VN.n18 VN.n17 0.189894
R1661 VN.n19 VN.n18 0.189894
R1662 VN.n19 VN.n2 0.189894
R1663 VN.n24 VN.n2 0.189894
R1664 VN.n25 VN.n24 0.189894
R1665 VN.n26 VN.n25 0.189894
R1666 VN.n26 VN.n0 0.189894
R1667 VN.n30 VN.n0 0.189894
R1668 VN VN.n30 0.0516364
R1669 VDD2.n1 VDD2.t3 69.1917
R1670 VDD2.n4 VDD2.t8 67.459
R1671 VDD2.n3 VDD2.n2 66.2973
R1672 VDD2 VDD2.n7 66.2945
R1673 VDD2.n6 VDD2.n5 65.0533
R1674 VDD2.n1 VDD2.n0 65.053
R1675 VDD2.n4 VDD2.n3 39.0407
R1676 VDD2.n7 VDD2.t1 2.40633
R1677 VDD2.n7 VDD2.t4 2.40633
R1678 VDD2.n5 VDD2.t9 2.40633
R1679 VDD2.n5 VDD2.t0 2.40633
R1680 VDD2.n2 VDD2.t5 2.40633
R1681 VDD2.n2 VDD2.t7 2.40633
R1682 VDD2.n0 VDD2.t2 2.40633
R1683 VDD2.n0 VDD2.t6 2.40633
R1684 VDD2.n6 VDD2.n4 1.73326
R1685 VDD2 VDD2.n6 0.491879
R1686 VDD2.n3 VDD2.n1 0.378344
C0 VDD2 VDD1 1.57251f
C1 VP VDD2 0.465474f
C2 VN VDD1 0.150834f
C3 VDD1 VTAIL 8.494431f
C4 VN VP 6.346971f
C5 VP VTAIL 7.16042f
C6 VN VDD2 6.73484f
C7 VDD2 VTAIL 8.53916f
C8 VN VTAIL 7.146121f
C9 VP VDD1 7.04636f
C10 VDD2 B 5.442591f
C11 VDD1 B 5.424747f
C12 VTAIL B 5.99002f
C13 VN B 13.482271f
C14 VP B 11.975913f
C15 VDD2.t3 B 1.61944f
C16 VDD2.t2 B 0.145902f
C17 VDD2.t6 B 0.145902f
C18 VDD2.n0 B 1.26648f
C19 VDD2.n1 B 0.690953f
C20 VDD2.t5 B 0.145902f
C21 VDD2.t7 B 0.145902f
C22 VDD2.n2 B 1.27406f
C23 VDD2.n3 B 1.9634f
C24 VDD2.t8 B 1.61025f
C25 VDD2.n4 B 2.20743f
C26 VDD2.t9 B 0.145902f
C27 VDD2.t0 B 0.145902f
C28 VDD2.n5 B 1.26649f
C29 VDD2.n6 B 0.339652f
C30 VDD2.t1 B 0.145902f
C31 VDD2.t4 B 0.145902f
C32 VDD2.n7 B 1.27402f
C33 VN.n0 B 0.028794f
C34 VN.t2 B 1.07052f
C35 VN.n1 B 0.023362f
C36 VN.n2 B 0.028794f
C37 VN.t4 B 1.07052f
C38 VN.n3 B 0.023287f
C39 VN.n4 B 0.028794f
C40 VN.t3 B 1.07052f
C41 VN.n5 B 0.023287f
C42 VN.n6 B 0.181956f
C43 VN.t7 B 1.07052f
C44 VN.t6 B 1.16895f
C45 VN.n7 B 0.475741f
C46 VN.n8 B 0.447037f
C47 VN.n9 B 0.0277f
C48 VN.n10 B 0.057081f
C49 VN.n11 B 0.028794f
C50 VN.n12 B 0.028794f
C51 VN.n13 B 0.028794f
C52 VN.n14 B 0.05737f
C53 VN.n15 B 0.425567f
C54 VN.n16 B 0.05737f
C55 VN.n17 B 0.028794f
C56 VN.n18 B 0.028794f
C57 VN.n19 B 0.028794f
C58 VN.n20 B 0.057081f
C59 VN.n21 B 0.0277f
C60 VN.n22 B 0.398397f
C61 VN.n23 B 0.05709f
C62 VN.n24 B 0.028794f
C63 VN.n25 B 0.028794f
C64 VN.n26 B 0.028794f
C65 VN.n27 B 0.056756f
C66 VN.n28 B 0.02823f
C67 VN.n29 B 0.454491f
C68 VN.n30 B 0.030482f
C69 VN.n31 B 0.028794f
C70 VN.t1 B 1.07052f
C71 VN.n32 B 0.023362f
C72 VN.n33 B 0.028794f
C73 VN.t0 B 1.07052f
C74 VN.n34 B 0.023287f
C75 VN.n35 B 0.028794f
C76 VN.t9 B 1.07052f
C77 VN.n36 B 0.023287f
C78 VN.n37 B 0.181956f
C79 VN.t8 B 1.07052f
C80 VN.t5 B 1.16895f
C81 VN.n38 B 0.475741f
C82 VN.n39 B 0.447037f
C83 VN.n40 B 0.0277f
C84 VN.n41 B 0.057081f
C85 VN.n42 B 0.028794f
C86 VN.n43 B 0.028794f
C87 VN.n44 B 0.028794f
C88 VN.n45 B 0.05737f
C89 VN.n46 B 0.425567f
C90 VN.n47 B 0.05737f
C91 VN.n48 B 0.028794f
C92 VN.n49 B 0.028794f
C93 VN.n50 B 0.028794f
C94 VN.n51 B 0.057081f
C95 VN.n52 B 0.0277f
C96 VN.n53 B 0.398397f
C97 VN.n54 B 0.05709f
C98 VN.n55 B 0.028794f
C99 VN.n56 B 0.028794f
C100 VN.n57 B 0.028794f
C101 VN.n58 B 0.056756f
C102 VN.n59 B 0.02823f
C103 VN.n60 B 0.454491f
C104 VN.n61 B 1.36106f
C105 VTAIL.t8 B 0.167175f
C106 VTAIL.t3 B 0.167175f
C107 VTAIL.n0 B 1.38217f
C108 VTAIL.n1 B 0.462136f
C109 VTAIL.t15 B 1.75893f
C110 VTAIL.n2 B 0.572366f
C111 VTAIL.t13 B 0.167175f
C112 VTAIL.t14 B 0.167175f
C113 VTAIL.n3 B 1.38217f
C114 VTAIL.n4 B 0.526042f
C115 VTAIL.t10 B 0.167175f
C116 VTAIL.t17 B 0.167175f
C117 VTAIL.n5 B 1.38217f
C118 VTAIL.n6 B 1.60638f
C119 VTAIL.t2 B 0.167175f
C120 VTAIL.t1 B 0.167175f
C121 VTAIL.n7 B 1.38217f
C122 VTAIL.n8 B 1.60638f
C123 VTAIL.t9 B 0.167175f
C124 VTAIL.t7 B 0.167175f
C125 VTAIL.n9 B 1.38217f
C126 VTAIL.n10 B 0.526038f
C127 VTAIL.t5 B 1.75894f
C128 VTAIL.n11 B 0.572353f
C129 VTAIL.t11 B 0.167175f
C130 VTAIL.t19 B 0.167175f
C131 VTAIL.n12 B 1.38217f
C132 VTAIL.n13 B 0.493193f
C133 VTAIL.t18 B 0.167175f
C134 VTAIL.t12 B 0.167175f
C135 VTAIL.n14 B 1.38217f
C136 VTAIL.n15 B 0.526038f
C137 VTAIL.t16 B 1.75893f
C138 VTAIL.n16 B 1.54203f
C139 VTAIL.t6 B 1.75893f
C140 VTAIL.n17 B 1.54203f
C141 VTAIL.t4 B 0.167175f
C142 VTAIL.t0 B 0.167175f
C143 VTAIL.n18 B 1.38217f
C144 VTAIL.n19 B 0.413582f
C145 VDD1.t5 B 1.64245f
C146 VDD1.t1 B 0.147975f
C147 VDD1.t2 B 0.147975f
C148 VDD1.n0 B 1.28448f
C149 VDD1.n1 B 0.707687f
C150 VDD1.t8 B 1.64245f
C151 VDD1.t4 B 0.147975f
C152 VDD1.t0 B 0.147975f
C153 VDD1.n2 B 1.28448f
C154 VDD1.n3 B 0.70077f
C155 VDD1.t6 B 0.147975f
C156 VDD1.t3 B 0.147975f
C157 VDD1.n4 B 1.29216f
C158 VDD1.n5 B 2.0811f
C159 VDD1.t9 B 0.147975f
C160 VDD1.t7 B 0.147975f
C161 VDD1.n6 B 1.28447f
C162 VDD1.n7 B 2.26912f
C163 VP.n0 B 0.029426f
C164 VP.t4 B 1.09402f
C165 VP.n1 B 0.023875f
C166 VP.n2 B 0.029426f
C167 VP.t5 B 1.09402f
C168 VP.n3 B 0.023799f
C169 VP.n4 B 0.029426f
C170 VP.t6 B 1.09402f
C171 VP.n5 B 0.023799f
C172 VP.n6 B 0.029426f
C173 VP.t2 B 1.09402f
C174 VP.n7 B 0.023875f
C175 VP.n8 B 0.029426f
C176 VP.t9 B 1.09402f
C177 VP.n9 B 0.029426f
C178 VP.t3 B 1.09402f
C179 VP.n10 B 0.023875f
C180 VP.n11 B 0.029426f
C181 VP.t7 B 1.09402f
C182 VP.n12 B 0.023799f
C183 VP.n13 B 0.029426f
C184 VP.t1 B 1.09402f
C185 VP.n14 B 0.023799f
C186 VP.n15 B 0.185951f
C187 VP.t0 B 1.09402f
C188 VP.t8 B 1.19461f
C189 VP.n16 B 0.486187f
C190 VP.n17 B 0.456853f
C191 VP.n18 B 0.028308f
C192 VP.n19 B 0.058334f
C193 VP.n20 B 0.029426f
C194 VP.n21 B 0.029426f
C195 VP.n22 B 0.029426f
C196 VP.n23 B 0.058629f
C197 VP.n24 B 0.434911f
C198 VP.n25 B 0.058629f
C199 VP.n26 B 0.029426f
C200 VP.n27 B 0.029426f
C201 VP.n28 B 0.029426f
C202 VP.n29 B 0.058334f
C203 VP.n30 B 0.028308f
C204 VP.n31 B 0.407145f
C205 VP.n32 B 0.058344f
C206 VP.n33 B 0.029426f
C207 VP.n34 B 0.029426f
C208 VP.n35 B 0.029426f
C209 VP.n36 B 0.058003f
C210 VP.n37 B 0.02885f
C211 VP.n38 B 0.46447f
C212 VP.n39 B 1.37171f
C213 VP.n40 B 1.39518f
C214 VP.n41 B 0.46447f
C215 VP.n42 B 0.02885f
C216 VP.n43 B 0.058003f
C217 VP.n44 B 0.029426f
C218 VP.n45 B 0.029426f
C219 VP.n46 B 0.029426f
C220 VP.n47 B 0.058344f
C221 VP.n48 B 0.407145f
C222 VP.n49 B 0.028308f
C223 VP.n50 B 0.058334f
C224 VP.n51 B 0.029426f
C225 VP.n52 B 0.029426f
C226 VP.n53 B 0.029426f
C227 VP.n54 B 0.058629f
C228 VP.n55 B 0.434911f
C229 VP.n56 B 0.058629f
C230 VP.n57 B 0.029426f
C231 VP.n58 B 0.029426f
C232 VP.n59 B 0.029426f
C233 VP.n60 B 0.058334f
C234 VP.n61 B 0.028308f
C235 VP.n62 B 0.407145f
C236 VP.n63 B 0.058344f
C237 VP.n64 B 0.029426f
C238 VP.n65 B 0.029426f
C239 VP.n66 B 0.029426f
C240 VP.n67 B 0.058003f
C241 VP.n68 B 0.02885f
C242 VP.n69 B 0.46447f
C243 VP.n70 B 0.031152f
.ends

