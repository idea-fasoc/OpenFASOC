* NGSPICE file created from diff_pair_sample_0562.ext - technology: sky130A

.subckt diff_pair_sample_0562 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=2.2803 ps=14.15 w=13.82 l=0.38
X1 VDD1.t9 VP.t0 VTAIL.t3 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X2 VDD1.t8 VP.t1 VTAIL.t2 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=2.2803 ps=14.15 w=13.82 l=0.38
X3 VTAIL.t7 VP.t2 VDD1.t7 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X4 VDD1.t6 VP.t3 VTAIL.t4 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=5.3898 ps=28.42 w=13.82 l=0.38
X5 B.t11 B.t9 B.t10 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=0 ps=0 w=13.82 l=0.38
X6 VDD2.t8 VN.t1 VTAIL.t17 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X7 VDD1.t5 VP.t4 VTAIL.t5 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=5.3898 ps=28.42 w=13.82 l=0.38
X8 VDD1.t4 VP.t5 VTAIL.t0 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X9 VDD2.t7 VN.t2 VTAIL.t19 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=5.3898 ps=28.42 w=13.82 l=0.38
X10 VTAIL.t11 VN.t3 VDD2.t6 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X11 VDD2.t5 VN.t4 VTAIL.t13 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=2.2803 ps=14.15 w=13.82 l=0.38
X12 B.t8 B.t6 B.t7 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=0 ps=0 w=13.82 l=0.38
X13 VTAIL.t15 VN.t5 VDD2.t4 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X14 B.t5 B.t3 B.t4 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=0 ps=0 w=13.82 l=0.38
X15 VTAIL.t8 VP.t6 VDD1.t3 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X16 VTAIL.t6 VP.t7 VDD1.t2 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X17 VDD2.t3 VN.t6 VTAIL.t18 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X18 VTAIL.t12 VN.t7 VDD2.t2 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X19 VTAIL.t14 VN.t8 VDD2.t1 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X20 VDD1.t1 VP.t8 VTAIL.t9 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=2.2803 ps=14.15 w=13.82 l=0.38
X21 VTAIL.t1 VP.t9 VDD1.t0 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=2.2803 ps=14.15 w=13.82 l=0.38
X22 VDD2.t0 VN.t9 VTAIL.t10 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=2.2803 pd=14.15 as=5.3898 ps=28.42 w=13.82 l=0.38
X23 B.t2 B.t0 B.t1 w_n1822_n3732# sky130_fd_pr__pfet_01v8 ad=5.3898 pd=28.42 as=0 ps=0 w=13.82 l=0.38
R0 VN.n2 VN.t4 1002.11
R1 VN.n13 VN.t2 1002.11
R2 VN.n3 VN.t8 981.125
R3 VN.n1 VN.t1 981.125
R4 VN.n8 VN.t5 981.125
R5 VN.n9 VN.t9 981.125
R6 VN.n14 VN.t3 981.125
R7 VN.n12 VN.t6 981.125
R8 VN.n19 VN.t7 981.125
R9 VN.n20 VN.t0 981.125
R10 VN.n10 VN.n9 161.3
R11 VN.n21 VN.n20 161.3
R12 VN.n19 VN.n11 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n8 VN.n0 161.3
R16 VN.n7 VN.n6 161.3
R17 VN.n5 VN.n4 161.3
R18 VN.n16 VN.n13 70.4033
R19 VN.n5 VN.n2 70.4033
R20 VN.n9 VN.n8 48.2005
R21 VN.n20 VN.n19 48.2005
R22 VN VN.n21 42.8092
R23 VN.n4 VN.n3 39.4369
R24 VN.n8 VN.n7 39.4369
R25 VN.n15 VN.n14 39.4369
R26 VN.n19 VN.n18 39.4369
R27 VN.n14 VN.n13 20.9576
R28 VN.n3 VN.n2 20.9576
R29 VN.n4 VN.n1 8.76414
R30 VN.n7 VN.n1 8.76414
R31 VN.n15 VN.n12 8.76414
R32 VN.n18 VN.n12 8.76414
R33 VN.n21 VN.n11 0.189894
R34 VN.n17 VN.n11 0.189894
R35 VN.n17 VN.n16 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n6 VN.n0 0.189894
R38 VN.n10 VN.n0 0.189894
R39 VN VN.n10 0.0516364
R40 VTAIL.n16 VTAIL.t4 55.681
R41 VTAIL.n11 VTAIL.t19 55.681
R42 VTAIL.n17 VTAIL.t10 55.6808
R43 VTAIL.n2 VTAIL.t5 55.6808
R44 VTAIL.n15 VTAIL.n14 53.329
R45 VTAIL.n13 VTAIL.n12 53.329
R46 VTAIL.n10 VTAIL.n9 53.329
R47 VTAIL.n8 VTAIL.n7 53.329
R48 VTAIL.n19 VTAIL.n18 53.3289
R49 VTAIL.n1 VTAIL.n0 53.3289
R50 VTAIL.n4 VTAIL.n3 53.3289
R51 VTAIL.n6 VTAIL.n5 53.3289
R52 VTAIL.n8 VTAIL.n6 25.5048
R53 VTAIL.n17 VTAIL.n16 24.8927
R54 VTAIL.n18 VTAIL.t17 2.35253
R55 VTAIL.n18 VTAIL.t15 2.35253
R56 VTAIL.n0 VTAIL.t13 2.35253
R57 VTAIL.n0 VTAIL.t14 2.35253
R58 VTAIL.n3 VTAIL.t0 2.35253
R59 VTAIL.n3 VTAIL.t8 2.35253
R60 VTAIL.n5 VTAIL.t2 2.35253
R61 VTAIL.n5 VTAIL.t6 2.35253
R62 VTAIL.n14 VTAIL.t3 2.35253
R63 VTAIL.n14 VTAIL.t7 2.35253
R64 VTAIL.n12 VTAIL.t9 2.35253
R65 VTAIL.n12 VTAIL.t1 2.35253
R66 VTAIL.n9 VTAIL.t18 2.35253
R67 VTAIL.n9 VTAIL.t11 2.35253
R68 VTAIL.n7 VTAIL.t16 2.35253
R69 VTAIL.n7 VTAIL.t12 2.35253
R70 VTAIL.n13 VTAIL.n11 0.776362
R71 VTAIL.n2 VTAIL.n1 0.776362
R72 VTAIL.n10 VTAIL.n8 0.612569
R73 VTAIL.n11 VTAIL.n10 0.612569
R74 VTAIL.n15 VTAIL.n13 0.612569
R75 VTAIL.n16 VTAIL.n15 0.612569
R76 VTAIL.n6 VTAIL.n4 0.612569
R77 VTAIL.n4 VTAIL.n2 0.612569
R78 VTAIL.n19 VTAIL.n17 0.612569
R79 VTAIL VTAIL.n1 0.517741
R80 VTAIL VTAIL.n19 0.0953276
R81 VDD2.n1 VDD2.t5 72.9717
R82 VDD2.n4 VDD2.t9 72.3598
R83 VDD2.n3 VDD2.n2 70.4114
R84 VDD2 VDD2.n7 70.4086
R85 VDD2.n6 VDD2.n5 70.0078
R86 VDD2.n1 VDD2.n0 70.0077
R87 VDD2.n4 VDD2.n3 38.5364
R88 VDD2.n7 VDD2.t6 2.35253
R89 VDD2.n7 VDD2.t7 2.35253
R90 VDD2.n5 VDD2.t2 2.35253
R91 VDD2.n5 VDD2.t3 2.35253
R92 VDD2.n2 VDD2.t4 2.35253
R93 VDD2.n2 VDD2.t0 2.35253
R94 VDD2.n0 VDD2.t1 2.35253
R95 VDD2.n0 VDD2.t8 2.35253
R96 VDD2.n6 VDD2.n4 0.612569
R97 VDD2 VDD2.n6 0.211707
R98 VDD2.n3 VDD2.n1 0.0981712
R99 VP.n5 VP.t8 1002.11
R100 VP.n15 VP.t1 981.125
R101 VP.n16 VP.t7 981.125
R102 VP.n1 VP.t5 981.125
R103 VP.n21 VP.t6 981.125
R104 VP.n22 VP.t4 981.125
R105 VP.n12 VP.t3 981.125
R106 VP.n11 VP.t2 981.125
R107 VP.n4 VP.t0 981.125
R108 VP.n6 VP.t9 981.125
R109 VP.n23 VP.n22 161.3
R110 VP.n8 VP.n7 161.3
R111 VP.n10 VP.n9 161.3
R112 VP.n11 VP.n3 161.3
R113 VP.n13 VP.n12 161.3
R114 VP.n21 VP.n0 161.3
R115 VP.n20 VP.n19 161.3
R116 VP.n18 VP.n17 161.3
R117 VP.n16 VP.n2 161.3
R118 VP.n15 VP.n14 161.3
R119 VP.n8 VP.n5 70.4033
R120 VP.n16 VP.n15 48.2005
R121 VP.n22 VP.n21 48.2005
R122 VP.n12 VP.n11 48.2005
R123 VP.n14 VP.n13 42.4285
R124 VP.n17 VP.n16 39.4369
R125 VP.n21 VP.n20 39.4369
R126 VP.n11 VP.n10 39.4369
R127 VP.n7 VP.n6 39.4369
R128 VP.n6 VP.n5 20.9576
R129 VP.n17 VP.n1 8.76414
R130 VP.n20 VP.n1 8.76414
R131 VP.n10 VP.n4 8.76414
R132 VP.n7 VP.n4 8.76414
R133 VP.n9 VP.n8 0.189894
R134 VP.n9 VP.n3 0.189894
R135 VP.n13 VP.n3 0.189894
R136 VP.n14 VP.n2 0.189894
R137 VP.n18 VP.n2 0.189894
R138 VP.n19 VP.n18 0.189894
R139 VP.n19 VP.n0 0.189894
R140 VP.n23 VP.n0 0.189894
R141 VP VP.n23 0.0516364
R142 VDD1.n1 VDD1.t1 72.9718
R143 VDD1.n3 VDD1.t8 72.9717
R144 VDD1.n5 VDD1.n4 70.4114
R145 VDD1.n7 VDD1.n6 70.0078
R146 VDD1.n1 VDD1.n0 70.0078
R147 VDD1.n3 VDD1.n2 70.0077
R148 VDD1.n7 VDD1.n5 39.4255
R149 VDD1.n6 VDD1.t7 2.35253
R150 VDD1.n6 VDD1.t6 2.35253
R151 VDD1.n0 VDD1.t0 2.35253
R152 VDD1.n0 VDD1.t9 2.35253
R153 VDD1.n4 VDD1.t3 2.35253
R154 VDD1.n4 VDD1.t5 2.35253
R155 VDD1.n2 VDD1.t2 2.35253
R156 VDD1.n2 VDD1.t4 2.35253
R157 VDD1 VDD1.n7 0.401362
R158 VDD1 VDD1.n1 0.211707
R159 VDD1.n5 VDD1.n3 0.0981712
R160 B.n119 B.t0 1086.69
R161 B.n267 B.t6 1086.69
R162 B.n44 B.t9 1086.69
R163 B.n36 B.t3 1086.69
R164 B.n341 B.n90 585
R165 B.n340 B.n339 585
R166 B.n338 B.n91 585
R167 B.n337 B.n336 585
R168 B.n335 B.n92 585
R169 B.n334 B.n333 585
R170 B.n332 B.n93 585
R171 B.n331 B.n330 585
R172 B.n329 B.n94 585
R173 B.n328 B.n327 585
R174 B.n326 B.n95 585
R175 B.n325 B.n324 585
R176 B.n323 B.n96 585
R177 B.n322 B.n321 585
R178 B.n320 B.n97 585
R179 B.n319 B.n318 585
R180 B.n317 B.n98 585
R181 B.n316 B.n315 585
R182 B.n314 B.n99 585
R183 B.n313 B.n312 585
R184 B.n311 B.n100 585
R185 B.n310 B.n309 585
R186 B.n308 B.n101 585
R187 B.n307 B.n306 585
R188 B.n305 B.n102 585
R189 B.n304 B.n303 585
R190 B.n302 B.n103 585
R191 B.n301 B.n300 585
R192 B.n299 B.n104 585
R193 B.n298 B.n297 585
R194 B.n296 B.n105 585
R195 B.n295 B.n294 585
R196 B.n293 B.n106 585
R197 B.n292 B.n291 585
R198 B.n290 B.n107 585
R199 B.n289 B.n288 585
R200 B.n287 B.n108 585
R201 B.n286 B.n285 585
R202 B.n284 B.n109 585
R203 B.n283 B.n282 585
R204 B.n281 B.n110 585
R205 B.n280 B.n279 585
R206 B.n278 B.n111 585
R207 B.n277 B.n276 585
R208 B.n275 B.n112 585
R209 B.n274 B.n273 585
R210 B.n272 B.n113 585
R211 B.n271 B.n270 585
R212 B.n266 B.n114 585
R213 B.n265 B.n264 585
R214 B.n263 B.n115 585
R215 B.n262 B.n261 585
R216 B.n260 B.n116 585
R217 B.n259 B.n258 585
R218 B.n257 B.n117 585
R219 B.n256 B.n255 585
R220 B.n254 B.n118 585
R221 B.n252 B.n251 585
R222 B.n250 B.n121 585
R223 B.n249 B.n248 585
R224 B.n247 B.n122 585
R225 B.n246 B.n245 585
R226 B.n244 B.n123 585
R227 B.n243 B.n242 585
R228 B.n241 B.n124 585
R229 B.n240 B.n239 585
R230 B.n238 B.n125 585
R231 B.n237 B.n236 585
R232 B.n235 B.n126 585
R233 B.n234 B.n233 585
R234 B.n232 B.n127 585
R235 B.n231 B.n230 585
R236 B.n229 B.n128 585
R237 B.n228 B.n227 585
R238 B.n226 B.n129 585
R239 B.n225 B.n224 585
R240 B.n223 B.n130 585
R241 B.n222 B.n221 585
R242 B.n220 B.n131 585
R243 B.n219 B.n218 585
R244 B.n217 B.n132 585
R245 B.n216 B.n215 585
R246 B.n214 B.n133 585
R247 B.n213 B.n212 585
R248 B.n211 B.n134 585
R249 B.n210 B.n209 585
R250 B.n208 B.n135 585
R251 B.n207 B.n206 585
R252 B.n205 B.n136 585
R253 B.n204 B.n203 585
R254 B.n202 B.n137 585
R255 B.n201 B.n200 585
R256 B.n199 B.n138 585
R257 B.n198 B.n197 585
R258 B.n196 B.n139 585
R259 B.n195 B.n194 585
R260 B.n193 B.n140 585
R261 B.n192 B.n191 585
R262 B.n190 B.n141 585
R263 B.n189 B.n188 585
R264 B.n187 B.n142 585
R265 B.n186 B.n185 585
R266 B.n184 B.n143 585
R267 B.n183 B.n182 585
R268 B.n343 B.n342 585
R269 B.n344 B.n89 585
R270 B.n346 B.n345 585
R271 B.n347 B.n88 585
R272 B.n349 B.n348 585
R273 B.n350 B.n87 585
R274 B.n352 B.n351 585
R275 B.n353 B.n86 585
R276 B.n355 B.n354 585
R277 B.n356 B.n85 585
R278 B.n358 B.n357 585
R279 B.n359 B.n84 585
R280 B.n361 B.n360 585
R281 B.n362 B.n83 585
R282 B.n364 B.n363 585
R283 B.n365 B.n82 585
R284 B.n367 B.n366 585
R285 B.n368 B.n81 585
R286 B.n370 B.n369 585
R287 B.n371 B.n80 585
R288 B.n373 B.n372 585
R289 B.n374 B.n79 585
R290 B.n376 B.n375 585
R291 B.n377 B.n78 585
R292 B.n379 B.n378 585
R293 B.n380 B.n77 585
R294 B.n382 B.n381 585
R295 B.n383 B.n76 585
R296 B.n385 B.n384 585
R297 B.n386 B.n75 585
R298 B.n388 B.n387 585
R299 B.n389 B.n74 585
R300 B.n391 B.n390 585
R301 B.n392 B.n73 585
R302 B.n394 B.n393 585
R303 B.n395 B.n72 585
R304 B.n397 B.n396 585
R305 B.n398 B.n71 585
R306 B.n400 B.n399 585
R307 B.n401 B.n70 585
R308 B.n403 B.n402 585
R309 B.n404 B.n69 585
R310 B.n561 B.n12 585
R311 B.n560 B.n559 585
R312 B.n558 B.n13 585
R313 B.n557 B.n556 585
R314 B.n555 B.n14 585
R315 B.n554 B.n553 585
R316 B.n552 B.n15 585
R317 B.n551 B.n550 585
R318 B.n549 B.n16 585
R319 B.n548 B.n547 585
R320 B.n546 B.n17 585
R321 B.n545 B.n544 585
R322 B.n543 B.n18 585
R323 B.n542 B.n541 585
R324 B.n540 B.n19 585
R325 B.n539 B.n538 585
R326 B.n537 B.n20 585
R327 B.n536 B.n535 585
R328 B.n534 B.n21 585
R329 B.n533 B.n532 585
R330 B.n531 B.n22 585
R331 B.n530 B.n529 585
R332 B.n528 B.n23 585
R333 B.n527 B.n526 585
R334 B.n525 B.n24 585
R335 B.n524 B.n523 585
R336 B.n522 B.n25 585
R337 B.n521 B.n520 585
R338 B.n519 B.n26 585
R339 B.n518 B.n517 585
R340 B.n516 B.n27 585
R341 B.n515 B.n514 585
R342 B.n513 B.n28 585
R343 B.n512 B.n511 585
R344 B.n510 B.n29 585
R345 B.n509 B.n508 585
R346 B.n507 B.n30 585
R347 B.n506 B.n505 585
R348 B.n504 B.n31 585
R349 B.n503 B.n502 585
R350 B.n501 B.n32 585
R351 B.n500 B.n499 585
R352 B.n498 B.n33 585
R353 B.n497 B.n496 585
R354 B.n495 B.n34 585
R355 B.n494 B.n493 585
R356 B.n492 B.n35 585
R357 B.n490 B.n489 585
R358 B.n488 B.n38 585
R359 B.n487 B.n486 585
R360 B.n485 B.n39 585
R361 B.n484 B.n483 585
R362 B.n482 B.n40 585
R363 B.n481 B.n480 585
R364 B.n479 B.n41 585
R365 B.n478 B.n477 585
R366 B.n476 B.n42 585
R367 B.n475 B.n474 585
R368 B.n473 B.n43 585
R369 B.n472 B.n471 585
R370 B.n470 B.n47 585
R371 B.n469 B.n468 585
R372 B.n467 B.n48 585
R373 B.n466 B.n465 585
R374 B.n464 B.n49 585
R375 B.n463 B.n462 585
R376 B.n461 B.n50 585
R377 B.n460 B.n459 585
R378 B.n458 B.n51 585
R379 B.n457 B.n456 585
R380 B.n455 B.n52 585
R381 B.n454 B.n453 585
R382 B.n452 B.n53 585
R383 B.n451 B.n450 585
R384 B.n449 B.n54 585
R385 B.n448 B.n447 585
R386 B.n446 B.n55 585
R387 B.n445 B.n444 585
R388 B.n443 B.n56 585
R389 B.n442 B.n441 585
R390 B.n440 B.n57 585
R391 B.n439 B.n438 585
R392 B.n437 B.n58 585
R393 B.n436 B.n435 585
R394 B.n434 B.n59 585
R395 B.n433 B.n432 585
R396 B.n431 B.n60 585
R397 B.n430 B.n429 585
R398 B.n428 B.n61 585
R399 B.n427 B.n426 585
R400 B.n425 B.n62 585
R401 B.n424 B.n423 585
R402 B.n422 B.n63 585
R403 B.n421 B.n420 585
R404 B.n419 B.n64 585
R405 B.n418 B.n417 585
R406 B.n416 B.n65 585
R407 B.n415 B.n414 585
R408 B.n413 B.n66 585
R409 B.n412 B.n411 585
R410 B.n410 B.n67 585
R411 B.n409 B.n408 585
R412 B.n407 B.n68 585
R413 B.n406 B.n405 585
R414 B.n563 B.n562 585
R415 B.n564 B.n11 585
R416 B.n566 B.n565 585
R417 B.n567 B.n10 585
R418 B.n569 B.n568 585
R419 B.n570 B.n9 585
R420 B.n572 B.n571 585
R421 B.n573 B.n8 585
R422 B.n575 B.n574 585
R423 B.n576 B.n7 585
R424 B.n578 B.n577 585
R425 B.n579 B.n6 585
R426 B.n581 B.n580 585
R427 B.n582 B.n5 585
R428 B.n584 B.n583 585
R429 B.n585 B.n4 585
R430 B.n587 B.n586 585
R431 B.n588 B.n3 585
R432 B.n590 B.n589 585
R433 B.n591 B.n0 585
R434 B.n2 B.n1 585
R435 B.n154 B.n153 585
R436 B.n156 B.n155 585
R437 B.n157 B.n152 585
R438 B.n159 B.n158 585
R439 B.n160 B.n151 585
R440 B.n162 B.n161 585
R441 B.n163 B.n150 585
R442 B.n165 B.n164 585
R443 B.n166 B.n149 585
R444 B.n168 B.n167 585
R445 B.n169 B.n148 585
R446 B.n171 B.n170 585
R447 B.n172 B.n147 585
R448 B.n174 B.n173 585
R449 B.n175 B.n146 585
R450 B.n177 B.n176 585
R451 B.n178 B.n145 585
R452 B.n180 B.n179 585
R453 B.n181 B.n144 585
R454 B.n183 B.n144 482.89
R455 B.n343 B.n90 482.89
R456 B.n405 B.n404 482.89
R457 B.n562 B.n561 482.89
R458 B.n593 B.n592 256.663
R459 B.n592 B.n591 235.042
R460 B.n592 B.n2 235.042
R461 B.n184 B.n183 163.367
R462 B.n185 B.n184 163.367
R463 B.n185 B.n142 163.367
R464 B.n189 B.n142 163.367
R465 B.n190 B.n189 163.367
R466 B.n191 B.n190 163.367
R467 B.n191 B.n140 163.367
R468 B.n195 B.n140 163.367
R469 B.n196 B.n195 163.367
R470 B.n197 B.n196 163.367
R471 B.n197 B.n138 163.367
R472 B.n201 B.n138 163.367
R473 B.n202 B.n201 163.367
R474 B.n203 B.n202 163.367
R475 B.n203 B.n136 163.367
R476 B.n207 B.n136 163.367
R477 B.n208 B.n207 163.367
R478 B.n209 B.n208 163.367
R479 B.n209 B.n134 163.367
R480 B.n213 B.n134 163.367
R481 B.n214 B.n213 163.367
R482 B.n215 B.n214 163.367
R483 B.n215 B.n132 163.367
R484 B.n219 B.n132 163.367
R485 B.n220 B.n219 163.367
R486 B.n221 B.n220 163.367
R487 B.n221 B.n130 163.367
R488 B.n225 B.n130 163.367
R489 B.n226 B.n225 163.367
R490 B.n227 B.n226 163.367
R491 B.n227 B.n128 163.367
R492 B.n231 B.n128 163.367
R493 B.n232 B.n231 163.367
R494 B.n233 B.n232 163.367
R495 B.n233 B.n126 163.367
R496 B.n237 B.n126 163.367
R497 B.n238 B.n237 163.367
R498 B.n239 B.n238 163.367
R499 B.n239 B.n124 163.367
R500 B.n243 B.n124 163.367
R501 B.n244 B.n243 163.367
R502 B.n245 B.n244 163.367
R503 B.n245 B.n122 163.367
R504 B.n249 B.n122 163.367
R505 B.n250 B.n249 163.367
R506 B.n251 B.n250 163.367
R507 B.n251 B.n118 163.367
R508 B.n256 B.n118 163.367
R509 B.n257 B.n256 163.367
R510 B.n258 B.n257 163.367
R511 B.n258 B.n116 163.367
R512 B.n262 B.n116 163.367
R513 B.n263 B.n262 163.367
R514 B.n264 B.n263 163.367
R515 B.n264 B.n114 163.367
R516 B.n271 B.n114 163.367
R517 B.n272 B.n271 163.367
R518 B.n273 B.n272 163.367
R519 B.n273 B.n112 163.367
R520 B.n277 B.n112 163.367
R521 B.n278 B.n277 163.367
R522 B.n279 B.n278 163.367
R523 B.n279 B.n110 163.367
R524 B.n283 B.n110 163.367
R525 B.n284 B.n283 163.367
R526 B.n285 B.n284 163.367
R527 B.n285 B.n108 163.367
R528 B.n289 B.n108 163.367
R529 B.n290 B.n289 163.367
R530 B.n291 B.n290 163.367
R531 B.n291 B.n106 163.367
R532 B.n295 B.n106 163.367
R533 B.n296 B.n295 163.367
R534 B.n297 B.n296 163.367
R535 B.n297 B.n104 163.367
R536 B.n301 B.n104 163.367
R537 B.n302 B.n301 163.367
R538 B.n303 B.n302 163.367
R539 B.n303 B.n102 163.367
R540 B.n307 B.n102 163.367
R541 B.n308 B.n307 163.367
R542 B.n309 B.n308 163.367
R543 B.n309 B.n100 163.367
R544 B.n313 B.n100 163.367
R545 B.n314 B.n313 163.367
R546 B.n315 B.n314 163.367
R547 B.n315 B.n98 163.367
R548 B.n319 B.n98 163.367
R549 B.n320 B.n319 163.367
R550 B.n321 B.n320 163.367
R551 B.n321 B.n96 163.367
R552 B.n325 B.n96 163.367
R553 B.n326 B.n325 163.367
R554 B.n327 B.n326 163.367
R555 B.n327 B.n94 163.367
R556 B.n331 B.n94 163.367
R557 B.n332 B.n331 163.367
R558 B.n333 B.n332 163.367
R559 B.n333 B.n92 163.367
R560 B.n337 B.n92 163.367
R561 B.n338 B.n337 163.367
R562 B.n339 B.n338 163.367
R563 B.n339 B.n90 163.367
R564 B.n404 B.n403 163.367
R565 B.n403 B.n70 163.367
R566 B.n399 B.n70 163.367
R567 B.n399 B.n398 163.367
R568 B.n398 B.n397 163.367
R569 B.n397 B.n72 163.367
R570 B.n393 B.n72 163.367
R571 B.n393 B.n392 163.367
R572 B.n392 B.n391 163.367
R573 B.n391 B.n74 163.367
R574 B.n387 B.n74 163.367
R575 B.n387 B.n386 163.367
R576 B.n386 B.n385 163.367
R577 B.n385 B.n76 163.367
R578 B.n381 B.n76 163.367
R579 B.n381 B.n380 163.367
R580 B.n380 B.n379 163.367
R581 B.n379 B.n78 163.367
R582 B.n375 B.n78 163.367
R583 B.n375 B.n374 163.367
R584 B.n374 B.n373 163.367
R585 B.n373 B.n80 163.367
R586 B.n369 B.n80 163.367
R587 B.n369 B.n368 163.367
R588 B.n368 B.n367 163.367
R589 B.n367 B.n82 163.367
R590 B.n363 B.n82 163.367
R591 B.n363 B.n362 163.367
R592 B.n362 B.n361 163.367
R593 B.n361 B.n84 163.367
R594 B.n357 B.n84 163.367
R595 B.n357 B.n356 163.367
R596 B.n356 B.n355 163.367
R597 B.n355 B.n86 163.367
R598 B.n351 B.n86 163.367
R599 B.n351 B.n350 163.367
R600 B.n350 B.n349 163.367
R601 B.n349 B.n88 163.367
R602 B.n345 B.n88 163.367
R603 B.n345 B.n344 163.367
R604 B.n344 B.n343 163.367
R605 B.n561 B.n560 163.367
R606 B.n560 B.n13 163.367
R607 B.n556 B.n13 163.367
R608 B.n556 B.n555 163.367
R609 B.n555 B.n554 163.367
R610 B.n554 B.n15 163.367
R611 B.n550 B.n15 163.367
R612 B.n550 B.n549 163.367
R613 B.n549 B.n548 163.367
R614 B.n548 B.n17 163.367
R615 B.n544 B.n17 163.367
R616 B.n544 B.n543 163.367
R617 B.n543 B.n542 163.367
R618 B.n542 B.n19 163.367
R619 B.n538 B.n19 163.367
R620 B.n538 B.n537 163.367
R621 B.n537 B.n536 163.367
R622 B.n536 B.n21 163.367
R623 B.n532 B.n21 163.367
R624 B.n532 B.n531 163.367
R625 B.n531 B.n530 163.367
R626 B.n530 B.n23 163.367
R627 B.n526 B.n23 163.367
R628 B.n526 B.n525 163.367
R629 B.n525 B.n524 163.367
R630 B.n524 B.n25 163.367
R631 B.n520 B.n25 163.367
R632 B.n520 B.n519 163.367
R633 B.n519 B.n518 163.367
R634 B.n518 B.n27 163.367
R635 B.n514 B.n27 163.367
R636 B.n514 B.n513 163.367
R637 B.n513 B.n512 163.367
R638 B.n512 B.n29 163.367
R639 B.n508 B.n29 163.367
R640 B.n508 B.n507 163.367
R641 B.n507 B.n506 163.367
R642 B.n506 B.n31 163.367
R643 B.n502 B.n31 163.367
R644 B.n502 B.n501 163.367
R645 B.n501 B.n500 163.367
R646 B.n500 B.n33 163.367
R647 B.n496 B.n33 163.367
R648 B.n496 B.n495 163.367
R649 B.n495 B.n494 163.367
R650 B.n494 B.n35 163.367
R651 B.n489 B.n35 163.367
R652 B.n489 B.n488 163.367
R653 B.n488 B.n487 163.367
R654 B.n487 B.n39 163.367
R655 B.n483 B.n39 163.367
R656 B.n483 B.n482 163.367
R657 B.n482 B.n481 163.367
R658 B.n481 B.n41 163.367
R659 B.n477 B.n41 163.367
R660 B.n477 B.n476 163.367
R661 B.n476 B.n475 163.367
R662 B.n475 B.n43 163.367
R663 B.n471 B.n43 163.367
R664 B.n471 B.n470 163.367
R665 B.n470 B.n469 163.367
R666 B.n469 B.n48 163.367
R667 B.n465 B.n48 163.367
R668 B.n465 B.n464 163.367
R669 B.n464 B.n463 163.367
R670 B.n463 B.n50 163.367
R671 B.n459 B.n50 163.367
R672 B.n459 B.n458 163.367
R673 B.n458 B.n457 163.367
R674 B.n457 B.n52 163.367
R675 B.n453 B.n52 163.367
R676 B.n453 B.n452 163.367
R677 B.n452 B.n451 163.367
R678 B.n451 B.n54 163.367
R679 B.n447 B.n54 163.367
R680 B.n447 B.n446 163.367
R681 B.n446 B.n445 163.367
R682 B.n445 B.n56 163.367
R683 B.n441 B.n56 163.367
R684 B.n441 B.n440 163.367
R685 B.n440 B.n439 163.367
R686 B.n439 B.n58 163.367
R687 B.n435 B.n58 163.367
R688 B.n435 B.n434 163.367
R689 B.n434 B.n433 163.367
R690 B.n433 B.n60 163.367
R691 B.n429 B.n60 163.367
R692 B.n429 B.n428 163.367
R693 B.n428 B.n427 163.367
R694 B.n427 B.n62 163.367
R695 B.n423 B.n62 163.367
R696 B.n423 B.n422 163.367
R697 B.n422 B.n421 163.367
R698 B.n421 B.n64 163.367
R699 B.n417 B.n64 163.367
R700 B.n417 B.n416 163.367
R701 B.n416 B.n415 163.367
R702 B.n415 B.n66 163.367
R703 B.n411 B.n66 163.367
R704 B.n411 B.n410 163.367
R705 B.n410 B.n409 163.367
R706 B.n409 B.n68 163.367
R707 B.n405 B.n68 163.367
R708 B.n562 B.n11 163.367
R709 B.n566 B.n11 163.367
R710 B.n567 B.n566 163.367
R711 B.n568 B.n567 163.367
R712 B.n568 B.n9 163.367
R713 B.n572 B.n9 163.367
R714 B.n573 B.n572 163.367
R715 B.n574 B.n573 163.367
R716 B.n574 B.n7 163.367
R717 B.n578 B.n7 163.367
R718 B.n579 B.n578 163.367
R719 B.n580 B.n579 163.367
R720 B.n580 B.n5 163.367
R721 B.n584 B.n5 163.367
R722 B.n585 B.n584 163.367
R723 B.n586 B.n585 163.367
R724 B.n586 B.n3 163.367
R725 B.n590 B.n3 163.367
R726 B.n591 B.n590 163.367
R727 B.n154 B.n2 163.367
R728 B.n155 B.n154 163.367
R729 B.n155 B.n152 163.367
R730 B.n159 B.n152 163.367
R731 B.n160 B.n159 163.367
R732 B.n161 B.n160 163.367
R733 B.n161 B.n150 163.367
R734 B.n165 B.n150 163.367
R735 B.n166 B.n165 163.367
R736 B.n167 B.n166 163.367
R737 B.n167 B.n148 163.367
R738 B.n171 B.n148 163.367
R739 B.n172 B.n171 163.367
R740 B.n173 B.n172 163.367
R741 B.n173 B.n146 163.367
R742 B.n177 B.n146 163.367
R743 B.n178 B.n177 163.367
R744 B.n179 B.n178 163.367
R745 B.n179 B.n144 163.367
R746 B.n267 B.t7 124.781
R747 B.n44 B.t11 124.781
R748 B.n119 B.t1 124.764
R749 B.n36 B.t5 124.764
R750 B.n268 B.t8 111.013
R751 B.n45 B.t10 111.013
R752 B.n120 B.t2 110.996
R753 B.n37 B.t4 110.996
R754 B.n253 B.n120 59.5399
R755 B.n269 B.n268 59.5399
R756 B.n46 B.n45 59.5399
R757 B.n491 B.n37 59.5399
R758 B.n563 B.n12 31.3761
R759 B.n406 B.n69 31.3761
R760 B.n342 B.n341 31.3761
R761 B.n182 B.n181 31.3761
R762 B B.n593 18.0485
R763 B.n120 B.n119 13.7702
R764 B.n268 B.n267 13.7702
R765 B.n45 B.n44 13.7702
R766 B.n37 B.n36 13.7702
R767 B.n564 B.n563 10.6151
R768 B.n565 B.n564 10.6151
R769 B.n565 B.n10 10.6151
R770 B.n569 B.n10 10.6151
R771 B.n570 B.n569 10.6151
R772 B.n571 B.n570 10.6151
R773 B.n571 B.n8 10.6151
R774 B.n575 B.n8 10.6151
R775 B.n576 B.n575 10.6151
R776 B.n577 B.n576 10.6151
R777 B.n577 B.n6 10.6151
R778 B.n581 B.n6 10.6151
R779 B.n582 B.n581 10.6151
R780 B.n583 B.n582 10.6151
R781 B.n583 B.n4 10.6151
R782 B.n587 B.n4 10.6151
R783 B.n588 B.n587 10.6151
R784 B.n589 B.n588 10.6151
R785 B.n589 B.n0 10.6151
R786 B.n559 B.n12 10.6151
R787 B.n559 B.n558 10.6151
R788 B.n558 B.n557 10.6151
R789 B.n557 B.n14 10.6151
R790 B.n553 B.n14 10.6151
R791 B.n553 B.n552 10.6151
R792 B.n552 B.n551 10.6151
R793 B.n551 B.n16 10.6151
R794 B.n547 B.n16 10.6151
R795 B.n547 B.n546 10.6151
R796 B.n546 B.n545 10.6151
R797 B.n545 B.n18 10.6151
R798 B.n541 B.n18 10.6151
R799 B.n541 B.n540 10.6151
R800 B.n540 B.n539 10.6151
R801 B.n539 B.n20 10.6151
R802 B.n535 B.n20 10.6151
R803 B.n535 B.n534 10.6151
R804 B.n534 B.n533 10.6151
R805 B.n533 B.n22 10.6151
R806 B.n529 B.n22 10.6151
R807 B.n529 B.n528 10.6151
R808 B.n528 B.n527 10.6151
R809 B.n527 B.n24 10.6151
R810 B.n523 B.n24 10.6151
R811 B.n523 B.n522 10.6151
R812 B.n522 B.n521 10.6151
R813 B.n521 B.n26 10.6151
R814 B.n517 B.n26 10.6151
R815 B.n517 B.n516 10.6151
R816 B.n516 B.n515 10.6151
R817 B.n515 B.n28 10.6151
R818 B.n511 B.n28 10.6151
R819 B.n511 B.n510 10.6151
R820 B.n510 B.n509 10.6151
R821 B.n509 B.n30 10.6151
R822 B.n505 B.n30 10.6151
R823 B.n505 B.n504 10.6151
R824 B.n504 B.n503 10.6151
R825 B.n503 B.n32 10.6151
R826 B.n499 B.n32 10.6151
R827 B.n499 B.n498 10.6151
R828 B.n498 B.n497 10.6151
R829 B.n497 B.n34 10.6151
R830 B.n493 B.n34 10.6151
R831 B.n493 B.n492 10.6151
R832 B.n490 B.n38 10.6151
R833 B.n486 B.n38 10.6151
R834 B.n486 B.n485 10.6151
R835 B.n485 B.n484 10.6151
R836 B.n484 B.n40 10.6151
R837 B.n480 B.n40 10.6151
R838 B.n480 B.n479 10.6151
R839 B.n479 B.n478 10.6151
R840 B.n478 B.n42 10.6151
R841 B.n474 B.n473 10.6151
R842 B.n473 B.n472 10.6151
R843 B.n472 B.n47 10.6151
R844 B.n468 B.n47 10.6151
R845 B.n468 B.n467 10.6151
R846 B.n467 B.n466 10.6151
R847 B.n466 B.n49 10.6151
R848 B.n462 B.n49 10.6151
R849 B.n462 B.n461 10.6151
R850 B.n461 B.n460 10.6151
R851 B.n460 B.n51 10.6151
R852 B.n456 B.n51 10.6151
R853 B.n456 B.n455 10.6151
R854 B.n455 B.n454 10.6151
R855 B.n454 B.n53 10.6151
R856 B.n450 B.n53 10.6151
R857 B.n450 B.n449 10.6151
R858 B.n449 B.n448 10.6151
R859 B.n448 B.n55 10.6151
R860 B.n444 B.n55 10.6151
R861 B.n444 B.n443 10.6151
R862 B.n443 B.n442 10.6151
R863 B.n442 B.n57 10.6151
R864 B.n438 B.n57 10.6151
R865 B.n438 B.n437 10.6151
R866 B.n437 B.n436 10.6151
R867 B.n436 B.n59 10.6151
R868 B.n432 B.n59 10.6151
R869 B.n432 B.n431 10.6151
R870 B.n431 B.n430 10.6151
R871 B.n430 B.n61 10.6151
R872 B.n426 B.n61 10.6151
R873 B.n426 B.n425 10.6151
R874 B.n425 B.n424 10.6151
R875 B.n424 B.n63 10.6151
R876 B.n420 B.n63 10.6151
R877 B.n420 B.n419 10.6151
R878 B.n419 B.n418 10.6151
R879 B.n418 B.n65 10.6151
R880 B.n414 B.n65 10.6151
R881 B.n414 B.n413 10.6151
R882 B.n413 B.n412 10.6151
R883 B.n412 B.n67 10.6151
R884 B.n408 B.n67 10.6151
R885 B.n408 B.n407 10.6151
R886 B.n407 B.n406 10.6151
R887 B.n402 B.n69 10.6151
R888 B.n402 B.n401 10.6151
R889 B.n401 B.n400 10.6151
R890 B.n400 B.n71 10.6151
R891 B.n396 B.n71 10.6151
R892 B.n396 B.n395 10.6151
R893 B.n395 B.n394 10.6151
R894 B.n394 B.n73 10.6151
R895 B.n390 B.n73 10.6151
R896 B.n390 B.n389 10.6151
R897 B.n389 B.n388 10.6151
R898 B.n388 B.n75 10.6151
R899 B.n384 B.n75 10.6151
R900 B.n384 B.n383 10.6151
R901 B.n383 B.n382 10.6151
R902 B.n382 B.n77 10.6151
R903 B.n378 B.n77 10.6151
R904 B.n378 B.n377 10.6151
R905 B.n377 B.n376 10.6151
R906 B.n376 B.n79 10.6151
R907 B.n372 B.n79 10.6151
R908 B.n372 B.n371 10.6151
R909 B.n371 B.n370 10.6151
R910 B.n370 B.n81 10.6151
R911 B.n366 B.n81 10.6151
R912 B.n366 B.n365 10.6151
R913 B.n365 B.n364 10.6151
R914 B.n364 B.n83 10.6151
R915 B.n360 B.n83 10.6151
R916 B.n360 B.n359 10.6151
R917 B.n359 B.n358 10.6151
R918 B.n358 B.n85 10.6151
R919 B.n354 B.n85 10.6151
R920 B.n354 B.n353 10.6151
R921 B.n353 B.n352 10.6151
R922 B.n352 B.n87 10.6151
R923 B.n348 B.n87 10.6151
R924 B.n348 B.n347 10.6151
R925 B.n347 B.n346 10.6151
R926 B.n346 B.n89 10.6151
R927 B.n342 B.n89 10.6151
R928 B.n153 B.n1 10.6151
R929 B.n156 B.n153 10.6151
R930 B.n157 B.n156 10.6151
R931 B.n158 B.n157 10.6151
R932 B.n158 B.n151 10.6151
R933 B.n162 B.n151 10.6151
R934 B.n163 B.n162 10.6151
R935 B.n164 B.n163 10.6151
R936 B.n164 B.n149 10.6151
R937 B.n168 B.n149 10.6151
R938 B.n169 B.n168 10.6151
R939 B.n170 B.n169 10.6151
R940 B.n170 B.n147 10.6151
R941 B.n174 B.n147 10.6151
R942 B.n175 B.n174 10.6151
R943 B.n176 B.n175 10.6151
R944 B.n176 B.n145 10.6151
R945 B.n180 B.n145 10.6151
R946 B.n181 B.n180 10.6151
R947 B.n182 B.n143 10.6151
R948 B.n186 B.n143 10.6151
R949 B.n187 B.n186 10.6151
R950 B.n188 B.n187 10.6151
R951 B.n188 B.n141 10.6151
R952 B.n192 B.n141 10.6151
R953 B.n193 B.n192 10.6151
R954 B.n194 B.n193 10.6151
R955 B.n194 B.n139 10.6151
R956 B.n198 B.n139 10.6151
R957 B.n199 B.n198 10.6151
R958 B.n200 B.n199 10.6151
R959 B.n200 B.n137 10.6151
R960 B.n204 B.n137 10.6151
R961 B.n205 B.n204 10.6151
R962 B.n206 B.n205 10.6151
R963 B.n206 B.n135 10.6151
R964 B.n210 B.n135 10.6151
R965 B.n211 B.n210 10.6151
R966 B.n212 B.n211 10.6151
R967 B.n212 B.n133 10.6151
R968 B.n216 B.n133 10.6151
R969 B.n217 B.n216 10.6151
R970 B.n218 B.n217 10.6151
R971 B.n218 B.n131 10.6151
R972 B.n222 B.n131 10.6151
R973 B.n223 B.n222 10.6151
R974 B.n224 B.n223 10.6151
R975 B.n224 B.n129 10.6151
R976 B.n228 B.n129 10.6151
R977 B.n229 B.n228 10.6151
R978 B.n230 B.n229 10.6151
R979 B.n230 B.n127 10.6151
R980 B.n234 B.n127 10.6151
R981 B.n235 B.n234 10.6151
R982 B.n236 B.n235 10.6151
R983 B.n236 B.n125 10.6151
R984 B.n240 B.n125 10.6151
R985 B.n241 B.n240 10.6151
R986 B.n242 B.n241 10.6151
R987 B.n242 B.n123 10.6151
R988 B.n246 B.n123 10.6151
R989 B.n247 B.n246 10.6151
R990 B.n248 B.n247 10.6151
R991 B.n248 B.n121 10.6151
R992 B.n252 B.n121 10.6151
R993 B.n255 B.n254 10.6151
R994 B.n255 B.n117 10.6151
R995 B.n259 B.n117 10.6151
R996 B.n260 B.n259 10.6151
R997 B.n261 B.n260 10.6151
R998 B.n261 B.n115 10.6151
R999 B.n265 B.n115 10.6151
R1000 B.n266 B.n265 10.6151
R1001 B.n270 B.n266 10.6151
R1002 B.n274 B.n113 10.6151
R1003 B.n275 B.n274 10.6151
R1004 B.n276 B.n275 10.6151
R1005 B.n276 B.n111 10.6151
R1006 B.n280 B.n111 10.6151
R1007 B.n281 B.n280 10.6151
R1008 B.n282 B.n281 10.6151
R1009 B.n282 B.n109 10.6151
R1010 B.n286 B.n109 10.6151
R1011 B.n287 B.n286 10.6151
R1012 B.n288 B.n287 10.6151
R1013 B.n288 B.n107 10.6151
R1014 B.n292 B.n107 10.6151
R1015 B.n293 B.n292 10.6151
R1016 B.n294 B.n293 10.6151
R1017 B.n294 B.n105 10.6151
R1018 B.n298 B.n105 10.6151
R1019 B.n299 B.n298 10.6151
R1020 B.n300 B.n299 10.6151
R1021 B.n300 B.n103 10.6151
R1022 B.n304 B.n103 10.6151
R1023 B.n305 B.n304 10.6151
R1024 B.n306 B.n305 10.6151
R1025 B.n306 B.n101 10.6151
R1026 B.n310 B.n101 10.6151
R1027 B.n311 B.n310 10.6151
R1028 B.n312 B.n311 10.6151
R1029 B.n312 B.n99 10.6151
R1030 B.n316 B.n99 10.6151
R1031 B.n317 B.n316 10.6151
R1032 B.n318 B.n317 10.6151
R1033 B.n318 B.n97 10.6151
R1034 B.n322 B.n97 10.6151
R1035 B.n323 B.n322 10.6151
R1036 B.n324 B.n323 10.6151
R1037 B.n324 B.n95 10.6151
R1038 B.n328 B.n95 10.6151
R1039 B.n329 B.n328 10.6151
R1040 B.n330 B.n329 10.6151
R1041 B.n330 B.n93 10.6151
R1042 B.n334 B.n93 10.6151
R1043 B.n335 B.n334 10.6151
R1044 B.n336 B.n335 10.6151
R1045 B.n336 B.n91 10.6151
R1046 B.n340 B.n91 10.6151
R1047 B.n341 B.n340 10.6151
R1048 B.n492 B.n491 9.36635
R1049 B.n474 B.n46 9.36635
R1050 B.n253 B.n252 9.36635
R1051 B.n269 B.n113 9.36635
R1052 B.n593 B.n0 8.11757
R1053 B.n593 B.n1 8.11757
R1054 B.n491 B.n490 1.24928
R1055 B.n46 B.n42 1.24928
R1056 B.n254 B.n253 1.24928
R1057 B.n270 B.n269 1.24928
C0 VTAIL VDD2 21.3304f
C1 B VDD1 1.69005f
C2 VP w_n1822_n3732# 3.49236f
C3 VN VDD1 0.147962f
C4 VP VTAIL 4.8867f
C5 B VN 0.734536f
C6 w_n1822_n3732# VTAIL 3.3387f
C7 VDD1 VDD2 0.775314f
C8 B VDD2 1.72209f
C9 VP VDD1 5.43767f
C10 VN VDD2 5.29053f
C11 w_n1822_n3732# VDD1 2.03263f
C12 VP B 1.10966f
C13 B w_n1822_n3732# 7.32998f
C14 VDD1 VTAIL 21.301f
C15 VP VN 5.46768f
C16 B VTAIL 2.8065f
C17 w_n1822_n3732# VN 3.26199f
C18 VP VDD2 0.300924f
C19 VN VTAIL 4.87188f
C20 w_n1822_n3732# VDD2 2.0608f
C21 VDD2 VSUBS 1.536721f
C22 VDD1 VSUBS 1.106923f
C23 VTAIL VSUBS 0.658157f
C24 VN VSUBS 4.83061f
C25 VP VSUBS 1.485917f
C26 B VSUBS 2.759749f
C27 w_n1822_n3732# VSUBS 83.498604f
C28 B.n0 VSUBS 0.006559f
C29 B.n1 VSUBS 0.006559f
C30 B.n2 VSUBS 0.009701f
C31 B.n3 VSUBS 0.007434f
C32 B.n4 VSUBS 0.007434f
C33 B.n5 VSUBS 0.007434f
C34 B.n6 VSUBS 0.007434f
C35 B.n7 VSUBS 0.007434f
C36 B.n8 VSUBS 0.007434f
C37 B.n9 VSUBS 0.007434f
C38 B.n10 VSUBS 0.007434f
C39 B.n11 VSUBS 0.007434f
C40 B.n12 VSUBS 0.017669f
C41 B.n13 VSUBS 0.007434f
C42 B.n14 VSUBS 0.007434f
C43 B.n15 VSUBS 0.007434f
C44 B.n16 VSUBS 0.007434f
C45 B.n17 VSUBS 0.007434f
C46 B.n18 VSUBS 0.007434f
C47 B.n19 VSUBS 0.007434f
C48 B.n20 VSUBS 0.007434f
C49 B.n21 VSUBS 0.007434f
C50 B.n22 VSUBS 0.007434f
C51 B.n23 VSUBS 0.007434f
C52 B.n24 VSUBS 0.007434f
C53 B.n25 VSUBS 0.007434f
C54 B.n26 VSUBS 0.007434f
C55 B.n27 VSUBS 0.007434f
C56 B.n28 VSUBS 0.007434f
C57 B.n29 VSUBS 0.007434f
C58 B.n30 VSUBS 0.007434f
C59 B.n31 VSUBS 0.007434f
C60 B.n32 VSUBS 0.007434f
C61 B.n33 VSUBS 0.007434f
C62 B.n34 VSUBS 0.007434f
C63 B.n35 VSUBS 0.007434f
C64 B.t4 VSUBS 0.485058f
C65 B.t5 VSUBS 0.491238f
C66 B.t3 VSUBS 0.220264f
C67 B.n36 VSUBS 0.121645f
C68 B.n37 VSUBS 0.066591f
C69 B.n38 VSUBS 0.007434f
C70 B.n39 VSUBS 0.007434f
C71 B.n40 VSUBS 0.007434f
C72 B.n41 VSUBS 0.007434f
C73 B.n42 VSUBS 0.004154f
C74 B.n43 VSUBS 0.007434f
C75 B.t10 VSUBS 0.485047f
C76 B.t11 VSUBS 0.491226f
C77 B.t9 VSUBS 0.220264f
C78 B.n44 VSUBS 0.121657f
C79 B.n45 VSUBS 0.066602f
C80 B.n46 VSUBS 0.017223f
C81 B.n47 VSUBS 0.007434f
C82 B.n48 VSUBS 0.007434f
C83 B.n49 VSUBS 0.007434f
C84 B.n50 VSUBS 0.007434f
C85 B.n51 VSUBS 0.007434f
C86 B.n52 VSUBS 0.007434f
C87 B.n53 VSUBS 0.007434f
C88 B.n54 VSUBS 0.007434f
C89 B.n55 VSUBS 0.007434f
C90 B.n56 VSUBS 0.007434f
C91 B.n57 VSUBS 0.007434f
C92 B.n58 VSUBS 0.007434f
C93 B.n59 VSUBS 0.007434f
C94 B.n60 VSUBS 0.007434f
C95 B.n61 VSUBS 0.007434f
C96 B.n62 VSUBS 0.007434f
C97 B.n63 VSUBS 0.007434f
C98 B.n64 VSUBS 0.007434f
C99 B.n65 VSUBS 0.007434f
C100 B.n66 VSUBS 0.007434f
C101 B.n67 VSUBS 0.007434f
C102 B.n68 VSUBS 0.007434f
C103 B.n69 VSUBS 0.01622f
C104 B.n70 VSUBS 0.007434f
C105 B.n71 VSUBS 0.007434f
C106 B.n72 VSUBS 0.007434f
C107 B.n73 VSUBS 0.007434f
C108 B.n74 VSUBS 0.007434f
C109 B.n75 VSUBS 0.007434f
C110 B.n76 VSUBS 0.007434f
C111 B.n77 VSUBS 0.007434f
C112 B.n78 VSUBS 0.007434f
C113 B.n79 VSUBS 0.007434f
C114 B.n80 VSUBS 0.007434f
C115 B.n81 VSUBS 0.007434f
C116 B.n82 VSUBS 0.007434f
C117 B.n83 VSUBS 0.007434f
C118 B.n84 VSUBS 0.007434f
C119 B.n85 VSUBS 0.007434f
C120 B.n86 VSUBS 0.007434f
C121 B.n87 VSUBS 0.007434f
C122 B.n88 VSUBS 0.007434f
C123 B.n89 VSUBS 0.007434f
C124 B.n90 VSUBS 0.017669f
C125 B.n91 VSUBS 0.007434f
C126 B.n92 VSUBS 0.007434f
C127 B.n93 VSUBS 0.007434f
C128 B.n94 VSUBS 0.007434f
C129 B.n95 VSUBS 0.007434f
C130 B.n96 VSUBS 0.007434f
C131 B.n97 VSUBS 0.007434f
C132 B.n98 VSUBS 0.007434f
C133 B.n99 VSUBS 0.007434f
C134 B.n100 VSUBS 0.007434f
C135 B.n101 VSUBS 0.007434f
C136 B.n102 VSUBS 0.007434f
C137 B.n103 VSUBS 0.007434f
C138 B.n104 VSUBS 0.007434f
C139 B.n105 VSUBS 0.007434f
C140 B.n106 VSUBS 0.007434f
C141 B.n107 VSUBS 0.007434f
C142 B.n108 VSUBS 0.007434f
C143 B.n109 VSUBS 0.007434f
C144 B.n110 VSUBS 0.007434f
C145 B.n111 VSUBS 0.007434f
C146 B.n112 VSUBS 0.007434f
C147 B.n113 VSUBS 0.006996f
C148 B.n114 VSUBS 0.007434f
C149 B.n115 VSUBS 0.007434f
C150 B.n116 VSUBS 0.007434f
C151 B.n117 VSUBS 0.007434f
C152 B.n118 VSUBS 0.007434f
C153 B.t2 VSUBS 0.485058f
C154 B.t1 VSUBS 0.491238f
C155 B.t0 VSUBS 0.220264f
C156 B.n119 VSUBS 0.121645f
C157 B.n120 VSUBS 0.066591f
C158 B.n121 VSUBS 0.007434f
C159 B.n122 VSUBS 0.007434f
C160 B.n123 VSUBS 0.007434f
C161 B.n124 VSUBS 0.007434f
C162 B.n125 VSUBS 0.007434f
C163 B.n126 VSUBS 0.007434f
C164 B.n127 VSUBS 0.007434f
C165 B.n128 VSUBS 0.007434f
C166 B.n129 VSUBS 0.007434f
C167 B.n130 VSUBS 0.007434f
C168 B.n131 VSUBS 0.007434f
C169 B.n132 VSUBS 0.007434f
C170 B.n133 VSUBS 0.007434f
C171 B.n134 VSUBS 0.007434f
C172 B.n135 VSUBS 0.007434f
C173 B.n136 VSUBS 0.007434f
C174 B.n137 VSUBS 0.007434f
C175 B.n138 VSUBS 0.007434f
C176 B.n139 VSUBS 0.007434f
C177 B.n140 VSUBS 0.007434f
C178 B.n141 VSUBS 0.007434f
C179 B.n142 VSUBS 0.007434f
C180 B.n143 VSUBS 0.007434f
C181 B.n144 VSUBS 0.01622f
C182 B.n145 VSUBS 0.007434f
C183 B.n146 VSUBS 0.007434f
C184 B.n147 VSUBS 0.007434f
C185 B.n148 VSUBS 0.007434f
C186 B.n149 VSUBS 0.007434f
C187 B.n150 VSUBS 0.007434f
C188 B.n151 VSUBS 0.007434f
C189 B.n152 VSUBS 0.007434f
C190 B.n153 VSUBS 0.007434f
C191 B.n154 VSUBS 0.007434f
C192 B.n155 VSUBS 0.007434f
C193 B.n156 VSUBS 0.007434f
C194 B.n157 VSUBS 0.007434f
C195 B.n158 VSUBS 0.007434f
C196 B.n159 VSUBS 0.007434f
C197 B.n160 VSUBS 0.007434f
C198 B.n161 VSUBS 0.007434f
C199 B.n162 VSUBS 0.007434f
C200 B.n163 VSUBS 0.007434f
C201 B.n164 VSUBS 0.007434f
C202 B.n165 VSUBS 0.007434f
C203 B.n166 VSUBS 0.007434f
C204 B.n167 VSUBS 0.007434f
C205 B.n168 VSUBS 0.007434f
C206 B.n169 VSUBS 0.007434f
C207 B.n170 VSUBS 0.007434f
C208 B.n171 VSUBS 0.007434f
C209 B.n172 VSUBS 0.007434f
C210 B.n173 VSUBS 0.007434f
C211 B.n174 VSUBS 0.007434f
C212 B.n175 VSUBS 0.007434f
C213 B.n176 VSUBS 0.007434f
C214 B.n177 VSUBS 0.007434f
C215 B.n178 VSUBS 0.007434f
C216 B.n179 VSUBS 0.007434f
C217 B.n180 VSUBS 0.007434f
C218 B.n181 VSUBS 0.01622f
C219 B.n182 VSUBS 0.017669f
C220 B.n183 VSUBS 0.017669f
C221 B.n184 VSUBS 0.007434f
C222 B.n185 VSUBS 0.007434f
C223 B.n186 VSUBS 0.007434f
C224 B.n187 VSUBS 0.007434f
C225 B.n188 VSUBS 0.007434f
C226 B.n189 VSUBS 0.007434f
C227 B.n190 VSUBS 0.007434f
C228 B.n191 VSUBS 0.007434f
C229 B.n192 VSUBS 0.007434f
C230 B.n193 VSUBS 0.007434f
C231 B.n194 VSUBS 0.007434f
C232 B.n195 VSUBS 0.007434f
C233 B.n196 VSUBS 0.007434f
C234 B.n197 VSUBS 0.007434f
C235 B.n198 VSUBS 0.007434f
C236 B.n199 VSUBS 0.007434f
C237 B.n200 VSUBS 0.007434f
C238 B.n201 VSUBS 0.007434f
C239 B.n202 VSUBS 0.007434f
C240 B.n203 VSUBS 0.007434f
C241 B.n204 VSUBS 0.007434f
C242 B.n205 VSUBS 0.007434f
C243 B.n206 VSUBS 0.007434f
C244 B.n207 VSUBS 0.007434f
C245 B.n208 VSUBS 0.007434f
C246 B.n209 VSUBS 0.007434f
C247 B.n210 VSUBS 0.007434f
C248 B.n211 VSUBS 0.007434f
C249 B.n212 VSUBS 0.007434f
C250 B.n213 VSUBS 0.007434f
C251 B.n214 VSUBS 0.007434f
C252 B.n215 VSUBS 0.007434f
C253 B.n216 VSUBS 0.007434f
C254 B.n217 VSUBS 0.007434f
C255 B.n218 VSUBS 0.007434f
C256 B.n219 VSUBS 0.007434f
C257 B.n220 VSUBS 0.007434f
C258 B.n221 VSUBS 0.007434f
C259 B.n222 VSUBS 0.007434f
C260 B.n223 VSUBS 0.007434f
C261 B.n224 VSUBS 0.007434f
C262 B.n225 VSUBS 0.007434f
C263 B.n226 VSUBS 0.007434f
C264 B.n227 VSUBS 0.007434f
C265 B.n228 VSUBS 0.007434f
C266 B.n229 VSUBS 0.007434f
C267 B.n230 VSUBS 0.007434f
C268 B.n231 VSUBS 0.007434f
C269 B.n232 VSUBS 0.007434f
C270 B.n233 VSUBS 0.007434f
C271 B.n234 VSUBS 0.007434f
C272 B.n235 VSUBS 0.007434f
C273 B.n236 VSUBS 0.007434f
C274 B.n237 VSUBS 0.007434f
C275 B.n238 VSUBS 0.007434f
C276 B.n239 VSUBS 0.007434f
C277 B.n240 VSUBS 0.007434f
C278 B.n241 VSUBS 0.007434f
C279 B.n242 VSUBS 0.007434f
C280 B.n243 VSUBS 0.007434f
C281 B.n244 VSUBS 0.007434f
C282 B.n245 VSUBS 0.007434f
C283 B.n246 VSUBS 0.007434f
C284 B.n247 VSUBS 0.007434f
C285 B.n248 VSUBS 0.007434f
C286 B.n249 VSUBS 0.007434f
C287 B.n250 VSUBS 0.007434f
C288 B.n251 VSUBS 0.007434f
C289 B.n252 VSUBS 0.006996f
C290 B.n253 VSUBS 0.017223f
C291 B.n254 VSUBS 0.004154f
C292 B.n255 VSUBS 0.007434f
C293 B.n256 VSUBS 0.007434f
C294 B.n257 VSUBS 0.007434f
C295 B.n258 VSUBS 0.007434f
C296 B.n259 VSUBS 0.007434f
C297 B.n260 VSUBS 0.007434f
C298 B.n261 VSUBS 0.007434f
C299 B.n262 VSUBS 0.007434f
C300 B.n263 VSUBS 0.007434f
C301 B.n264 VSUBS 0.007434f
C302 B.n265 VSUBS 0.007434f
C303 B.n266 VSUBS 0.007434f
C304 B.t8 VSUBS 0.485047f
C305 B.t7 VSUBS 0.491226f
C306 B.t6 VSUBS 0.220264f
C307 B.n267 VSUBS 0.121657f
C308 B.n268 VSUBS 0.066602f
C309 B.n269 VSUBS 0.017223f
C310 B.n270 VSUBS 0.004154f
C311 B.n271 VSUBS 0.007434f
C312 B.n272 VSUBS 0.007434f
C313 B.n273 VSUBS 0.007434f
C314 B.n274 VSUBS 0.007434f
C315 B.n275 VSUBS 0.007434f
C316 B.n276 VSUBS 0.007434f
C317 B.n277 VSUBS 0.007434f
C318 B.n278 VSUBS 0.007434f
C319 B.n279 VSUBS 0.007434f
C320 B.n280 VSUBS 0.007434f
C321 B.n281 VSUBS 0.007434f
C322 B.n282 VSUBS 0.007434f
C323 B.n283 VSUBS 0.007434f
C324 B.n284 VSUBS 0.007434f
C325 B.n285 VSUBS 0.007434f
C326 B.n286 VSUBS 0.007434f
C327 B.n287 VSUBS 0.007434f
C328 B.n288 VSUBS 0.007434f
C329 B.n289 VSUBS 0.007434f
C330 B.n290 VSUBS 0.007434f
C331 B.n291 VSUBS 0.007434f
C332 B.n292 VSUBS 0.007434f
C333 B.n293 VSUBS 0.007434f
C334 B.n294 VSUBS 0.007434f
C335 B.n295 VSUBS 0.007434f
C336 B.n296 VSUBS 0.007434f
C337 B.n297 VSUBS 0.007434f
C338 B.n298 VSUBS 0.007434f
C339 B.n299 VSUBS 0.007434f
C340 B.n300 VSUBS 0.007434f
C341 B.n301 VSUBS 0.007434f
C342 B.n302 VSUBS 0.007434f
C343 B.n303 VSUBS 0.007434f
C344 B.n304 VSUBS 0.007434f
C345 B.n305 VSUBS 0.007434f
C346 B.n306 VSUBS 0.007434f
C347 B.n307 VSUBS 0.007434f
C348 B.n308 VSUBS 0.007434f
C349 B.n309 VSUBS 0.007434f
C350 B.n310 VSUBS 0.007434f
C351 B.n311 VSUBS 0.007434f
C352 B.n312 VSUBS 0.007434f
C353 B.n313 VSUBS 0.007434f
C354 B.n314 VSUBS 0.007434f
C355 B.n315 VSUBS 0.007434f
C356 B.n316 VSUBS 0.007434f
C357 B.n317 VSUBS 0.007434f
C358 B.n318 VSUBS 0.007434f
C359 B.n319 VSUBS 0.007434f
C360 B.n320 VSUBS 0.007434f
C361 B.n321 VSUBS 0.007434f
C362 B.n322 VSUBS 0.007434f
C363 B.n323 VSUBS 0.007434f
C364 B.n324 VSUBS 0.007434f
C365 B.n325 VSUBS 0.007434f
C366 B.n326 VSUBS 0.007434f
C367 B.n327 VSUBS 0.007434f
C368 B.n328 VSUBS 0.007434f
C369 B.n329 VSUBS 0.007434f
C370 B.n330 VSUBS 0.007434f
C371 B.n331 VSUBS 0.007434f
C372 B.n332 VSUBS 0.007434f
C373 B.n333 VSUBS 0.007434f
C374 B.n334 VSUBS 0.007434f
C375 B.n335 VSUBS 0.007434f
C376 B.n336 VSUBS 0.007434f
C377 B.n337 VSUBS 0.007434f
C378 B.n338 VSUBS 0.007434f
C379 B.n339 VSUBS 0.007434f
C380 B.n340 VSUBS 0.007434f
C381 B.n341 VSUBS 0.016755f
C382 B.n342 VSUBS 0.017134f
C383 B.n343 VSUBS 0.01622f
C384 B.n344 VSUBS 0.007434f
C385 B.n345 VSUBS 0.007434f
C386 B.n346 VSUBS 0.007434f
C387 B.n347 VSUBS 0.007434f
C388 B.n348 VSUBS 0.007434f
C389 B.n349 VSUBS 0.007434f
C390 B.n350 VSUBS 0.007434f
C391 B.n351 VSUBS 0.007434f
C392 B.n352 VSUBS 0.007434f
C393 B.n353 VSUBS 0.007434f
C394 B.n354 VSUBS 0.007434f
C395 B.n355 VSUBS 0.007434f
C396 B.n356 VSUBS 0.007434f
C397 B.n357 VSUBS 0.007434f
C398 B.n358 VSUBS 0.007434f
C399 B.n359 VSUBS 0.007434f
C400 B.n360 VSUBS 0.007434f
C401 B.n361 VSUBS 0.007434f
C402 B.n362 VSUBS 0.007434f
C403 B.n363 VSUBS 0.007434f
C404 B.n364 VSUBS 0.007434f
C405 B.n365 VSUBS 0.007434f
C406 B.n366 VSUBS 0.007434f
C407 B.n367 VSUBS 0.007434f
C408 B.n368 VSUBS 0.007434f
C409 B.n369 VSUBS 0.007434f
C410 B.n370 VSUBS 0.007434f
C411 B.n371 VSUBS 0.007434f
C412 B.n372 VSUBS 0.007434f
C413 B.n373 VSUBS 0.007434f
C414 B.n374 VSUBS 0.007434f
C415 B.n375 VSUBS 0.007434f
C416 B.n376 VSUBS 0.007434f
C417 B.n377 VSUBS 0.007434f
C418 B.n378 VSUBS 0.007434f
C419 B.n379 VSUBS 0.007434f
C420 B.n380 VSUBS 0.007434f
C421 B.n381 VSUBS 0.007434f
C422 B.n382 VSUBS 0.007434f
C423 B.n383 VSUBS 0.007434f
C424 B.n384 VSUBS 0.007434f
C425 B.n385 VSUBS 0.007434f
C426 B.n386 VSUBS 0.007434f
C427 B.n387 VSUBS 0.007434f
C428 B.n388 VSUBS 0.007434f
C429 B.n389 VSUBS 0.007434f
C430 B.n390 VSUBS 0.007434f
C431 B.n391 VSUBS 0.007434f
C432 B.n392 VSUBS 0.007434f
C433 B.n393 VSUBS 0.007434f
C434 B.n394 VSUBS 0.007434f
C435 B.n395 VSUBS 0.007434f
C436 B.n396 VSUBS 0.007434f
C437 B.n397 VSUBS 0.007434f
C438 B.n398 VSUBS 0.007434f
C439 B.n399 VSUBS 0.007434f
C440 B.n400 VSUBS 0.007434f
C441 B.n401 VSUBS 0.007434f
C442 B.n402 VSUBS 0.007434f
C443 B.n403 VSUBS 0.007434f
C444 B.n404 VSUBS 0.01622f
C445 B.n405 VSUBS 0.017669f
C446 B.n406 VSUBS 0.017669f
C447 B.n407 VSUBS 0.007434f
C448 B.n408 VSUBS 0.007434f
C449 B.n409 VSUBS 0.007434f
C450 B.n410 VSUBS 0.007434f
C451 B.n411 VSUBS 0.007434f
C452 B.n412 VSUBS 0.007434f
C453 B.n413 VSUBS 0.007434f
C454 B.n414 VSUBS 0.007434f
C455 B.n415 VSUBS 0.007434f
C456 B.n416 VSUBS 0.007434f
C457 B.n417 VSUBS 0.007434f
C458 B.n418 VSUBS 0.007434f
C459 B.n419 VSUBS 0.007434f
C460 B.n420 VSUBS 0.007434f
C461 B.n421 VSUBS 0.007434f
C462 B.n422 VSUBS 0.007434f
C463 B.n423 VSUBS 0.007434f
C464 B.n424 VSUBS 0.007434f
C465 B.n425 VSUBS 0.007434f
C466 B.n426 VSUBS 0.007434f
C467 B.n427 VSUBS 0.007434f
C468 B.n428 VSUBS 0.007434f
C469 B.n429 VSUBS 0.007434f
C470 B.n430 VSUBS 0.007434f
C471 B.n431 VSUBS 0.007434f
C472 B.n432 VSUBS 0.007434f
C473 B.n433 VSUBS 0.007434f
C474 B.n434 VSUBS 0.007434f
C475 B.n435 VSUBS 0.007434f
C476 B.n436 VSUBS 0.007434f
C477 B.n437 VSUBS 0.007434f
C478 B.n438 VSUBS 0.007434f
C479 B.n439 VSUBS 0.007434f
C480 B.n440 VSUBS 0.007434f
C481 B.n441 VSUBS 0.007434f
C482 B.n442 VSUBS 0.007434f
C483 B.n443 VSUBS 0.007434f
C484 B.n444 VSUBS 0.007434f
C485 B.n445 VSUBS 0.007434f
C486 B.n446 VSUBS 0.007434f
C487 B.n447 VSUBS 0.007434f
C488 B.n448 VSUBS 0.007434f
C489 B.n449 VSUBS 0.007434f
C490 B.n450 VSUBS 0.007434f
C491 B.n451 VSUBS 0.007434f
C492 B.n452 VSUBS 0.007434f
C493 B.n453 VSUBS 0.007434f
C494 B.n454 VSUBS 0.007434f
C495 B.n455 VSUBS 0.007434f
C496 B.n456 VSUBS 0.007434f
C497 B.n457 VSUBS 0.007434f
C498 B.n458 VSUBS 0.007434f
C499 B.n459 VSUBS 0.007434f
C500 B.n460 VSUBS 0.007434f
C501 B.n461 VSUBS 0.007434f
C502 B.n462 VSUBS 0.007434f
C503 B.n463 VSUBS 0.007434f
C504 B.n464 VSUBS 0.007434f
C505 B.n465 VSUBS 0.007434f
C506 B.n466 VSUBS 0.007434f
C507 B.n467 VSUBS 0.007434f
C508 B.n468 VSUBS 0.007434f
C509 B.n469 VSUBS 0.007434f
C510 B.n470 VSUBS 0.007434f
C511 B.n471 VSUBS 0.007434f
C512 B.n472 VSUBS 0.007434f
C513 B.n473 VSUBS 0.007434f
C514 B.n474 VSUBS 0.006996f
C515 B.n475 VSUBS 0.007434f
C516 B.n476 VSUBS 0.007434f
C517 B.n477 VSUBS 0.007434f
C518 B.n478 VSUBS 0.007434f
C519 B.n479 VSUBS 0.007434f
C520 B.n480 VSUBS 0.007434f
C521 B.n481 VSUBS 0.007434f
C522 B.n482 VSUBS 0.007434f
C523 B.n483 VSUBS 0.007434f
C524 B.n484 VSUBS 0.007434f
C525 B.n485 VSUBS 0.007434f
C526 B.n486 VSUBS 0.007434f
C527 B.n487 VSUBS 0.007434f
C528 B.n488 VSUBS 0.007434f
C529 B.n489 VSUBS 0.007434f
C530 B.n490 VSUBS 0.004154f
C531 B.n491 VSUBS 0.017223f
C532 B.n492 VSUBS 0.006996f
C533 B.n493 VSUBS 0.007434f
C534 B.n494 VSUBS 0.007434f
C535 B.n495 VSUBS 0.007434f
C536 B.n496 VSUBS 0.007434f
C537 B.n497 VSUBS 0.007434f
C538 B.n498 VSUBS 0.007434f
C539 B.n499 VSUBS 0.007434f
C540 B.n500 VSUBS 0.007434f
C541 B.n501 VSUBS 0.007434f
C542 B.n502 VSUBS 0.007434f
C543 B.n503 VSUBS 0.007434f
C544 B.n504 VSUBS 0.007434f
C545 B.n505 VSUBS 0.007434f
C546 B.n506 VSUBS 0.007434f
C547 B.n507 VSUBS 0.007434f
C548 B.n508 VSUBS 0.007434f
C549 B.n509 VSUBS 0.007434f
C550 B.n510 VSUBS 0.007434f
C551 B.n511 VSUBS 0.007434f
C552 B.n512 VSUBS 0.007434f
C553 B.n513 VSUBS 0.007434f
C554 B.n514 VSUBS 0.007434f
C555 B.n515 VSUBS 0.007434f
C556 B.n516 VSUBS 0.007434f
C557 B.n517 VSUBS 0.007434f
C558 B.n518 VSUBS 0.007434f
C559 B.n519 VSUBS 0.007434f
C560 B.n520 VSUBS 0.007434f
C561 B.n521 VSUBS 0.007434f
C562 B.n522 VSUBS 0.007434f
C563 B.n523 VSUBS 0.007434f
C564 B.n524 VSUBS 0.007434f
C565 B.n525 VSUBS 0.007434f
C566 B.n526 VSUBS 0.007434f
C567 B.n527 VSUBS 0.007434f
C568 B.n528 VSUBS 0.007434f
C569 B.n529 VSUBS 0.007434f
C570 B.n530 VSUBS 0.007434f
C571 B.n531 VSUBS 0.007434f
C572 B.n532 VSUBS 0.007434f
C573 B.n533 VSUBS 0.007434f
C574 B.n534 VSUBS 0.007434f
C575 B.n535 VSUBS 0.007434f
C576 B.n536 VSUBS 0.007434f
C577 B.n537 VSUBS 0.007434f
C578 B.n538 VSUBS 0.007434f
C579 B.n539 VSUBS 0.007434f
C580 B.n540 VSUBS 0.007434f
C581 B.n541 VSUBS 0.007434f
C582 B.n542 VSUBS 0.007434f
C583 B.n543 VSUBS 0.007434f
C584 B.n544 VSUBS 0.007434f
C585 B.n545 VSUBS 0.007434f
C586 B.n546 VSUBS 0.007434f
C587 B.n547 VSUBS 0.007434f
C588 B.n548 VSUBS 0.007434f
C589 B.n549 VSUBS 0.007434f
C590 B.n550 VSUBS 0.007434f
C591 B.n551 VSUBS 0.007434f
C592 B.n552 VSUBS 0.007434f
C593 B.n553 VSUBS 0.007434f
C594 B.n554 VSUBS 0.007434f
C595 B.n555 VSUBS 0.007434f
C596 B.n556 VSUBS 0.007434f
C597 B.n557 VSUBS 0.007434f
C598 B.n558 VSUBS 0.007434f
C599 B.n559 VSUBS 0.007434f
C600 B.n560 VSUBS 0.007434f
C601 B.n561 VSUBS 0.017669f
C602 B.n562 VSUBS 0.01622f
C603 B.n563 VSUBS 0.01622f
C604 B.n564 VSUBS 0.007434f
C605 B.n565 VSUBS 0.007434f
C606 B.n566 VSUBS 0.007434f
C607 B.n567 VSUBS 0.007434f
C608 B.n568 VSUBS 0.007434f
C609 B.n569 VSUBS 0.007434f
C610 B.n570 VSUBS 0.007434f
C611 B.n571 VSUBS 0.007434f
C612 B.n572 VSUBS 0.007434f
C613 B.n573 VSUBS 0.007434f
C614 B.n574 VSUBS 0.007434f
C615 B.n575 VSUBS 0.007434f
C616 B.n576 VSUBS 0.007434f
C617 B.n577 VSUBS 0.007434f
C618 B.n578 VSUBS 0.007434f
C619 B.n579 VSUBS 0.007434f
C620 B.n580 VSUBS 0.007434f
C621 B.n581 VSUBS 0.007434f
C622 B.n582 VSUBS 0.007434f
C623 B.n583 VSUBS 0.007434f
C624 B.n584 VSUBS 0.007434f
C625 B.n585 VSUBS 0.007434f
C626 B.n586 VSUBS 0.007434f
C627 B.n587 VSUBS 0.007434f
C628 B.n588 VSUBS 0.007434f
C629 B.n589 VSUBS 0.007434f
C630 B.n590 VSUBS 0.007434f
C631 B.n591 VSUBS 0.009701f
C632 B.n592 VSUBS 0.010334f
C633 B.n593 VSUBS 0.020549f
C634 VDD1.t1 VSUBS 3.41337f
C635 VDD1.t0 VSUBS 0.328717f
C636 VDD1.t9 VSUBS 0.328717f
C637 VDD1.n0 VSUBS 2.61387f
C638 VDD1.n1 VSUBS 1.42936f
C639 VDD1.t8 VSUBS 3.41336f
C640 VDD1.t2 VSUBS 0.328717f
C641 VDD1.t4 VSUBS 0.328717f
C642 VDD1.n2 VSUBS 2.61386f
C643 VDD1.n3 VSUBS 1.42551f
C644 VDD1.t3 VSUBS 0.328717f
C645 VDD1.t5 VSUBS 0.328717f
C646 VDD1.n4 VSUBS 2.61789f
C647 VDD1.n5 VSUBS 2.64261f
C648 VDD1.t7 VSUBS 0.328717f
C649 VDD1.t6 VSUBS 0.328717f
C650 VDD1.n6 VSUBS 2.61387f
C651 VDD1.n7 VSUBS 3.22721f
C652 VP.n0 VSUBS 0.063206f
C653 VP.t5 VSUBS 0.944808f
C654 VP.n1 VSUBS 0.36658f
C655 VP.n2 VSUBS 0.063206f
C656 VP.n3 VSUBS 0.063206f
C657 VP.t3 VSUBS 0.944808f
C658 VP.t2 VSUBS 0.944808f
C659 VP.t0 VSUBS 0.944808f
C660 VP.n4 VSUBS 0.36658f
C661 VP.t8 VSUBS 0.952688f
C662 VP.n5 VSUBS 0.368814f
C663 VP.t9 VSUBS 0.944808f
C664 VP.n6 VSUBS 0.386768f
C665 VP.n7 VSUBS 0.014343f
C666 VP.n8 VSUBS 0.197743f
C667 VP.n9 VSUBS 0.063206f
C668 VP.n10 VSUBS 0.014343f
C669 VP.n11 VSUBS 0.386768f
C670 VP.n12 VSUBS 0.376246f
C671 VP.n13 VSUBS 2.65337f
C672 VP.n14 VSUBS 2.70676f
C673 VP.t1 VSUBS 0.944808f
C674 VP.n15 VSUBS 0.376246f
C675 VP.t7 VSUBS 0.944808f
C676 VP.n16 VSUBS 0.386768f
C677 VP.n17 VSUBS 0.014343f
C678 VP.n18 VSUBS 0.063206f
C679 VP.n19 VSUBS 0.063206f
C680 VP.n20 VSUBS 0.014343f
C681 VP.t6 VSUBS 0.944808f
C682 VP.n21 VSUBS 0.386768f
C683 VP.t4 VSUBS 0.944808f
C684 VP.n22 VSUBS 0.376246f
C685 VP.n23 VSUBS 0.048982f
C686 VDD2.t5 VSUBS 3.42663f
C687 VDD2.t1 VSUBS 0.329995f
C688 VDD2.t8 VSUBS 0.329995f
C689 VDD2.n0 VSUBS 2.62403f
C690 VDD2.n1 VSUBS 1.43105f
C691 VDD2.t4 VSUBS 0.329995f
C692 VDD2.t0 VSUBS 0.329995f
C693 VDD2.n2 VSUBS 2.62807f
C694 VDD2.n3 VSUBS 2.56829f
C695 VDD2.t9 VSUBS 3.4202f
C696 VDD2.n4 VSUBS 3.27753f
C697 VDD2.t2 VSUBS 0.329995f
C698 VDD2.t3 VSUBS 0.329995f
C699 VDD2.n5 VSUBS 2.62403f
C700 VDD2.n6 VSUBS 0.672969f
C701 VDD2.t6 VSUBS 0.329995f
C702 VDD2.t7 VSUBS 0.329995f
C703 VDD2.n7 VSUBS 2.62804f
C704 VTAIL.t13 VSUBS 0.351736f
C705 VTAIL.t14 VSUBS 0.351736f
C706 VTAIL.n0 VSUBS 2.6012f
C707 VTAIL.n1 VSUBS 0.917996f
C708 VTAIL.t5 VSUBS 3.42493f
C709 VTAIL.n2 VSUBS 1.06339f
C710 VTAIL.t0 VSUBS 0.351736f
C711 VTAIL.t8 VSUBS 0.351736f
C712 VTAIL.n3 VSUBS 2.6012f
C713 VTAIL.n4 VSUBS 0.910839f
C714 VTAIL.t2 VSUBS 0.351736f
C715 VTAIL.t6 VSUBS 0.351736f
C716 VTAIL.n5 VSUBS 2.6012f
C717 VTAIL.n6 VSUBS 2.64826f
C718 VTAIL.t16 VSUBS 0.351736f
C719 VTAIL.t12 VSUBS 0.351736f
C720 VTAIL.n7 VSUBS 2.60121f
C721 VTAIL.n8 VSUBS 2.64826f
C722 VTAIL.t18 VSUBS 0.351736f
C723 VTAIL.t11 VSUBS 0.351736f
C724 VTAIL.n9 VSUBS 2.60121f
C725 VTAIL.n10 VSUBS 0.910833f
C726 VTAIL.t19 VSUBS 3.42495f
C727 VTAIL.n11 VSUBS 1.06337f
C728 VTAIL.t9 VSUBS 0.351736f
C729 VTAIL.t1 VSUBS 0.351736f
C730 VTAIL.n12 VSUBS 2.60121f
C731 VTAIL.n13 VSUBS 0.927831f
C732 VTAIL.t3 VSUBS 0.351736f
C733 VTAIL.t7 VSUBS 0.351736f
C734 VTAIL.n14 VSUBS 2.60121f
C735 VTAIL.n15 VSUBS 0.910833f
C736 VTAIL.t4 VSUBS 3.42494f
C737 VTAIL.n16 VSUBS 2.72028f
C738 VTAIL.t10 VSUBS 3.42493f
C739 VTAIL.n17 VSUBS 2.7203f
C740 VTAIL.t17 VSUBS 0.351736f
C741 VTAIL.t15 VSUBS 0.351736f
C742 VTAIL.n18 VSUBS 2.6012f
C743 VTAIL.n19 VSUBS 0.85716f
C744 VN.n0 VSUBS 0.061938f
C745 VN.t1 VSUBS 0.92586f
C746 VN.n1 VSUBS 0.359228f
C747 VN.t4 VSUBS 0.933581f
C748 VN.n2 VSUBS 0.361417f
C749 VN.t8 VSUBS 0.92586f
C750 VN.n3 VSUBS 0.379011f
C751 VN.n4 VSUBS 0.014055f
C752 VN.n5 VSUBS 0.193777f
C753 VN.n6 VSUBS 0.061938f
C754 VN.n7 VSUBS 0.014055f
C755 VN.t5 VSUBS 0.92586f
C756 VN.n8 VSUBS 0.379011f
C757 VN.t9 VSUBS 0.92586f
C758 VN.n9 VSUBS 0.3687f
C759 VN.n10 VSUBS 0.048f
C760 VN.n11 VSUBS 0.061938f
C761 VN.t6 VSUBS 0.92586f
C762 VN.n12 VSUBS 0.359228f
C763 VN.t2 VSUBS 0.933581f
C764 VN.n13 VSUBS 0.361417f
C765 VN.t3 VSUBS 0.92586f
C766 VN.n14 VSUBS 0.379011f
C767 VN.n15 VSUBS 0.014055f
C768 VN.n16 VSUBS 0.193777f
C769 VN.n17 VSUBS 0.061938f
C770 VN.n18 VSUBS 0.014055f
C771 VN.t7 VSUBS 0.92586f
C772 VN.n19 VSUBS 0.379011f
C773 VN.t0 VSUBS 0.92586f
C774 VN.n20 VSUBS 0.3687f
C775 VN.n21 VSUBS 2.64079f
.ends

