* NGSPICE file created from diff_pair_sample_0851.ext - technology: sky130A

.subckt diff_pair_sample_0851 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X1 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=0 ps=0 w=14.86 l=1.36
X2 VTAIL.t18 VP.t1 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X3 VDD1.t9 VP.t2 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X4 VTAIL.t16 VP.t3 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X5 VTAIL.t5 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X6 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=0 ps=0 w=14.86 l=1.36
X7 VTAIL.t1 VN.t1 VDD2.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X8 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=0 ps=0 w=14.86 l=1.36
X9 VTAIL.t8 VN.t2 VDD2.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X10 VDD2.t6 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X11 VTAIL.t15 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X12 VTAIL.t3 VN.t4 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X13 VDD1.t2 VP.t5 VTAIL.t14 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=2.4519 ps=15.19 w=14.86 l=1.36
X14 VDD2.t4 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=5.7954 ps=30.5 w=14.86 l=1.36
X15 VDD1.t7 VP.t6 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=5.7954 ps=30.5 w=14.86 l=1.36
X16 VDD1.t6 VP.t7 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=2.4519 ps=15.19 w=14.86 l=1.36
X17 VDD2.t3 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X18 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=5.7954 ps=30.5 w=14.86 l=1.36
X19 VDD2.t1 VN.t8 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=2.4519 ps=15.19 w=14.86 l=1.36
X20 VDD1.t5 VP.t8 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=5.7954 ps=30.5 w=14.86 l=1.36
X21 VDD2.t0 VN.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=2.4519 ps=15.19 w=14.86 l=1.36
X22 VDD1.t4 VP.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4519 pd=15.19 as=2.4519 ps=15.19 w=14.86 l=1.36
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7954 pd=30.5 as=0 ps=0 w=14.86 l=1.36
R0 VP.n13 VP.t7 310.889
R1 VP.n31 VP.t5 292.212
R2 VP.n49 VP.t6 292.212
R3 VP.n28 VP.t8 292.212
R4 VP.n3 VP.t9 263.329
R5 VP.n5 VP.t3 263.329
R6 VP.n1 VP.t0 263.329
R7 VP.n10 VP.t2 263.329
R8 VP.n8 VP.t1 263.329
R9 VP.n12 VP.t4 263.329
R10 VP.n15 VP.n14 161.3
R11 VP.n16 VP.n11 161.3
R12 VP.n18 VP.n17 161.3
R13 VP.n19 VP.n10 161.3
R14 VP.n21 VP.n20 161.3
R15 VP.n22 VP.n9 161.3
R16 VP.n24 VP.n23 161.3
R17 VP.n26 VP.n25 161.3
R18 VP.n27 VP.n7 161.3
R19 VP.n48 VP.n0 161.3
R20 VP.n47 VP.n46 161.3
R21 VP.n45 VP.n44 161.3
R22 VP.n43 VP.n2 161.3
R23 VP.n42 VP.n41 161.3
R24 VP.n40 VP.n3 161.3
R25 VP.n39 VP.n38 161.3
R26 VP.n37 VP.n4 161.3
R27 VP.n36 VP.n35 161.3
R28 VP.n34 VP.n33 161.3
R29 VP.n32 VP.n6 161.3
R30 VP.n29 VP.n28 80.6037
R31 VP.n50 VP.n49 80.6037
R32 VP.n31 VP.n30 80.6037
R33 VP.n38 VP.n37 55.593
R34 VP.n43 VP.n42 55.593
R35 VP.n22 VP.n21 55.593
R36 VP.n17 VP.n16 55.593
R37 VP.n30 VP.n29 48.7552
R38 VP.n13 VP.n12 48.5618
R39 VP.n33 VP.n32 37.1863
R40 VP.n48 VP.n47 37.1863
R41 VP.n27 VP.n26 37.1863
R42 VP.n14 VP.n13 29.6663
R43 VP.n32 VP.n31 29.2126
R44 VP.n49 VP.n48 29.2126
R45 VP.n28 VP.n27 29.2126
R46 VP.n37 VP.n36 25.5611
R47 VP.n44 VP.n43 25.5611
R48 VP.n23 VP.n22 25.5611
R49 VP.n16 VP.n15 25.5611
R50 VP.n38 VP.n3 24.5923
R51 VP.n42 VP.n3 24.5923
R52 VP.n17 VP.n10 24.5923
R53 VP.n21 VP.n10 24.5923
R54 VP.n33 VP.n5 15.2474
R55 VP.n47 VP.n1 15.2474
R56 VP.n26 VP.n8 15.2474
R57 VP.n36 VP.n5 9.3454
R58 VP.n44 VP.n1 9.3454
R59 VP.n23 VP.n8 9.3454
R60 VP.n15 VP.n12 9.3454
R61 VP.n29 VP.n7 0.285035
R62 VP.n30 VP.n6 0.285035
R63 VP.n50 VP.n0 0.285035
R64 VP.n14 VP.n11 0.189894
R65 VP.n18 VP.n11 0.189894
R66 VP.n19 VP.n18 0.189894
R67 VP.n20 VP.n19 0.189894
R68 VP.n20 VP.n9 0.189894
R69 VP.n24 VP.n9 0.189894
R70 VP.n25 VP.n24 0.189894
R71 VP.n25 VP.n7 0.189894
R72 VP.n34 VP.n6 0.189894
R73 VP.n35 VP.n34 0.189894
R74 VP.n35 VP.n4 0.189894
R75 VP.n39 VP.n4 0.189894
R76 VP.n40 VP.n39 0.189894
R77 VP.n41 VP.n40 0.189894
R78 VP.n41 VP.n2 0.189894
R79 VP.n45 VP.n2 0.189894
R80 VP.n46 VP.n45 0.189894
R81 VP.n46 VP.n0 0.189894
R82 VP VP.n50 0.146778
R83 VDD1.n76 VDD1.n0 289.615
R84 VDD1.n159 VDD1.n83 289.615
R85 VDD1.n77 VDD1.n76 185
R86 VDD1.n75 VDD1.n74 185
R87 VDD1.n73 VDD1.n3 185
R88 VDD1.n7 VDD1.n4 185
R89 VDD1.n68 VDD1.n67 185
R90 VDD1.n66 VDD1.n65 185
R91 VDD1.n9 VDD1.n8 185
R92 VDD1.n60 VDD1.n59 185
R93 VDD1.n58 VDD1.n57 185
R94 VDD1.n13 VDD1.n12 185
R95 VDD1.n52 VDD1.n51 185
R96 VDD1.n50 VDD1.n49 185
R97 VDD1.n17 VDD1.n16 185
R98 VDD1.n44 VDD1.n43 185
R99 VDD1.n42 VDD1.n41 185
R100 VDD1.n21 VDD1.n20 185
R101 VDD1.n36 VDD1.n35 185
R102 VDD1.n34 VDD1.n33 185
R103 VDD1.n25 VDD1.n24 185
R104 VDD1.n28 VDD1.n27 185
R105 VDD1.n110 VDD1.n109 185
R106 VDD1.n107 VDD1.n106 185
R107 VDD1.n116 VDD1.n115 185
R108 VDD1.n118 VDD1.n117 185
R109 VDD1.n103 VDD1.n102 185
R110 VDD1.n124 VDD1.n123 185
R111 VDD1.n126 VDD1.n125 185
R112 VDD1.n99 VDD1.n98 185
R113 VDD1.n132 VDD1.n131 185
R114 VDD1.n134 VDD1.n133 185
R115 VDD1.n95 VDD1.n94 185
R116 VDD1.n140 VDD1.n139 185
R117 VDD1.n142 VDD1.n141 185
R118 VDD1.n91 VDD1.n90 185
R119 VDD1.n148 VDD1.n147 185
R120 VDD1.n151 VDD1.n150 185
R121 VDD1.n149 VDD1.n87 185
R122 VDD1.n156 VDD1.n86 185
R123 VDD1.n158 VDD1.n157 185
R124 VDD1.n160 VDD1.n159 185
R125 VDD1.t6 VDD1.n26 147.659
R126 VDD1.t2 VDD1.n108 147.659
R127 VDD1.n76 VDD1.n75 104.615
R128 VDD1.n75 VDD1.n3 104.615
R129 VDD1.n7 VDD1.n3 104.615
R130 VDD1.n67 VDD1.n7 104.615
R131 VDD1.n67 VDD1.n66 104.615
R132 VDD1.n66 VDD1.n8 104.615
R133 VDD1.n59 VDD1.n8 104.615
R134 VDD1.n59 VDD1.n58 104.615
R135 VDD1.n58 VDD1.n12 104.615
R136 VDD1.n51 VDD1.n12 104.615
R137 VDD1.n51 VDD1.n50 104.615
R138 VDD1.n50 VDD1.n16 104.615
R139 VDD1.n43 VDD1.n16 104.615
R140 VDD1.n43 VDD1.n42 104.615
R141 VDD1.n42 VDD1.n20 104.615
R142 VDD1.n35 VDD1.n20 104.615
R143 VDD1.n35 VDD1.n34 104.615
R144 VDD1.n34 VDD1.n24 104.615
R145 VDD1.n27 VDD1.n24 104.615
R146 VDD1.n109 VDD1.n106 104.615
R147 VDD1.n116 VDD1.n106 104.615
R148 VDD1.n117 VDD1.n116 104.615
R149 VDD1.n117 VDD1.n102 104.615
R150 VDD1.n124 VDD1.n102 104.615
R151 VDD1.n125 VDD1.n124 104.615
R152 VDD1.n125 VDD1.n98 104.615
R153 VDD1.n132 VDD1.n98 104.615
R154 VDD1.n133 VDD1.n132 104.615
R155 VDD1.n133 VDD1.n94 104.615
R156 VDD1.n140 VDD1.n94 104.615
R157 VDD1.n141 VDD1.n140 104.615
R158 VDD1.n141 VDD1.n90 104.615
R159 VDD1.n148 VDD1.n90 104.615
R160 VDD1.n150 VDD1.n148 104.615
R161 VDD1.n150 VDD1.n149 104.615
R162 VDD1.n149 VDD1.n86 104.615
R163 VDD1.n158 VDD1.n86 104.615
R164 VDD1.n159 VDD1.n158 104.615
R165 VDD1.n167 VDD1.n166 66.2249
R166 VDD1.n82 VDD1.n81 65.1878
R167 VDD1.n169 VDD1.n168 65.1876
R168 VDD1.n165 VDD1.n164 65.1876
R169 VDD1.n82 VDD1.n80 54.5877
R170 VDD1.n165 VDD1.n163 54.5877
R171 VDD1.n27 VDD1.t6 52.3082
R172 VDD1.n109 VDD1.t2 52.3082
R173 VDD1.n169 VDD1.n167 44.7574
R174 VDD1.n28 VDD1.n26 15.6677
R175 VDD1.n110 VDD1.n108 15.6677
R176 VDD1.n74 VDD1.n73 13.1884
R177 VDD1.n157 VDD1.n156 13.1884
R178 VDD1.n77 VDD1.n2 12.8005
R179 VDD1.n72 VDD1.n4 12.8005
R180 VDD1.n29 VDD1.n25 12.8005
R181 VDD1.n111 VDD1.n107 12.8005
R182 VDD1.n155 VDD1.n87 12.8005
R183 VDD1.n160 VDD1.n85 12.8005
R184 VDD1.n78 VDD1.n0 12.0247
R185 VDD1.n69 VDD1.n68 12.0247
R186 VDD1.n33 VDD1.n32 12.0247
R187 VDD1.n115 VDD1.n114 12.0247
R188 VDD1.n152 VDD1.n151 12.0247
R189 VDD1.n161 VDD1.n83 12.0247
R190 VDD1.n65 VDD1.n6 11.249
R191 VDD1.n36 VDD1.n23 11.249
R192 VDD1.n118 VDD1.n105 11.249
R193 VDD1.n147 VDD1.n89 11.249
R194 VDD1.n64 VDD1.n9 10.4732
R195 VDD1.n37 VDD1.n21 10.4732
R196 VDD1.n119 VDD1.n103 10.4732
R197 VDD1.n146 VDD1.n91 10.4732
R198 VDD1.n61 VDD1.n60 9.69747
R199 VDD1.n41 VDD1.n40 9.69747
R200 VDD1.n123 VDD1.n122 9.69747
R201 VDD1.n143 VDD1.n142 9.69747
R202 VDD1.n80 VDD1.n79 9.45567
R203 VDD1.n163 VDD1.n162 9.45567
R204 VDD1.n54 VDD1.n53 9.3005
R205 VDD1.n56 VDD1.n55 9.3005
R206 VDD1.n11 VDD1.n10 9.3005
R207 VDD1.n62 VDD1.n61 9.3005
R208 VDD1.n64 VDD1.n63 9.3005
R209 VDD1.n6 VDD1.n5 9.3005
R210 VDD1.n70 VDD1.n69 9.3005
R211 VDD1.n72 VDD1.n71 9.3005
R212 VDD1.n79 VDD1.n78 9.3005
R213 VDD1.n2 VDD1.n1 9.3005
R214 VDD1.n15 VDD1.n14 9.3005
R215 VDD1.n48 VDD1.n47 9.3005
R216 VDD1.n46 VDD1.n45 9.3005
R217 VDD1.n19 VDD1.n18 9.3005
R218 VDD1.n40 VDD1.n39 9.3005
R219 VDD1.n38 VDD1.n37 9.3005
R220 VDD1.n23 VDD1.n22 9.3005
R221 VDD1.n32 VDD1.n31 9.3005
R222 VDD1.n30 VDD1.n29 9.3005
R223 VDD1.n162 VDD1.n161 9.3005
R224 VDD1.n85 VDD1.n84 9.3005
R225 VDD1.n130 VDD1.n129 9.3005
R226 VDD1.n128 VDD1.n127 9.3005
R227 VDD1.n101 VDD1.n100 9.3005
R228 VDD1.n122 VDD1.n121 9.3005
R229 VDD1.n120 VDD1.n119 9.3005
R230 VDD1.n105 VDD1.n104 9.3005
R231 VDD1.n114 VDD1.n113 9.3005
R232 VDD1.n112 VDD1.n111 9.3005
R233 VDD1.n97 VDD1.n96 9.3005
R234 VDD1.n136 VDD1.n135 9.3005
R235 VDD1.n138 VDD1.n137 9.3005
R236 VDD1.n93 VDD1.n92 9.3005
R237 VDD1.n144 VDD1.n143 9.3005
R238 VDD1.n146 VDD1.n145 9.3005
R239 VDD1.n89 VDD1.n88 9.3005
R240 VDD1.n153 VDD1.n152 9.3005
R241 VDD1.n155 VDD1.n154 9.3005
R242 VDD1.n57 VDD1.n11 8.92171
R243 VDD1.n44 VDD1.n19 8.92171
R244 VDD1.n126 VDD1.n101 8.92171
R245 VDD1.n139 VDD1.n93 8.92171
R246 VDD1.n56 VDD1.n13 8.14595
R247 VDD1.n45 VDD1.n17 8.14595
R248 VDD1.n127 VDD1.n99 8.14595
R249 VDD1.n138 VDD1.n95 8.14595
R250 VDD1.n53 VDD1.n52 7.3702
R251 VDD1.n49 VDD1.n48 7.3702
R252 VDD1.n131 VDD1.n130 7.3702
R253 VDD1.n135 VDD1.n134 7.3702
R254 VDD1.n52 VDD1.n15 6.59444
R255 VDD1.n49 VDD1.n15 6.59444
R256 VDD1.n131 VDD1.n97 6.59444
R257 VDD1.n134 VDD1.n97 6.59444
R258 VDD1.n53 VDD1.n13 5.81868
R259 VDD1.n48 VDD1.n17 5.81868
R260 VDD1.n130 VDD1.n99 5.81868
R261 VDD1.n135 VDD1.n95 5.81868
R262 VDD1.n57 VDD1.n56 5.04292
R263 VDD1.n45 VDD1.n44 5.04292
R264 VDD1.n127 VDD1.n126 5.04292
R265 VDD1.n139 VDD1.n138 5.04292
R266 VDD1.n30 VDD1.n26 4.38563
R267 VDD1.n112 VDD1.n108 4.38563
R268 VDD1.n60 VDD1.n11 4.26717
R269 VDD1.n41 VDD1.n19 4.26717
R270 VDD1.n123 VDD1.n101 4.26717
R271 VDD1.n142 VDD1.n93 4.26717
R272 VDD1.n61 VDD1.n9 3.49141
R273 VDD1.n40 VDD1.n21 3.49141
R274 VDD1.n122 VDD1.n103 3.49141
R275 VDD1.n143 VDD1.n91 3.49141
R276 VDD1.n65 VDD1.n64 2.71565
R277 VDD1.n37 VDD1.n36 2.71565
R278 VDD1.n119 VDD1.n118 2.71565
R279 VDD1.n147 VDD1.n146 2.71565
R280 VDD1.n80 VDD1.n0 1.93989
R281 VDD1.n68 VDD1.n6 1.93989
R282 VDD1.n33 VDD1.n23 1.93989
R283 VDD1.n115 VDD1.n105 1.93989
R284 VDD1.n151 VDD1.n89 1.93989
R285 VDD1.n163 VDD1.n83 1.93989
R286 VDD1.n168 VDD1.t0 1.33294
R287 VDD1.n168 VDD1.t5 1.33294
R288 VDD1.n81 VDD1.t3 1.33294
R289 VDD1.n81 VDD1.t9 1.33294
R290 VDD1.n166 VDD1.t1 1.33294
R291 VDD1.n166 VDD1.t7 1.33294
R292 VDD1.n164 VDD1.t8 1.33294
R293 VDD1.n164 VDD1.t4 1.33294
R294 VDD1.n78 VDD1.n77 1.16414
R295 VDD1.n69 VDD1.n4 1.16414
R296 VDD1.n32 VDD1.n25 1.16414
R297 VDD1.n114 VDD1.n107 1.16414
R298 VDD1.n152 VDD1.n87 1.16414
R299 VDD1.n161 VDD1.n160 1.16414
R300 VDD1 VDD1.n169 1.03498
R301 VDD1 VDD1.n82 0.422914
R302 VDD1.n74 VDD1.n2 0.388379
R303 VDD1.n73 VDD1.n72 0.388379
R304 VDD1.n29 VDD1.n28 0.388379
R305 VDD1.n111 VDD1.n110 0.388379
R306 VDD1.n156 VDD1.n155 0.388379
R307 VDD1.n157 VDD1.n85 0.388379
R308 VDD1.n167 VDD1.n165 0.309378
R309 VDD1.n79 VDD1.n1 0.155672
R310 VDD1.n71 VDD1.n1 0.155672
R311 VDD1.n71 VDD1.n70 0.155672
R312 VDD1.n70 VDD1.n5 0.155672
R313 VDD1.n63 VDD1.n5 0.155672
R314 VDD1.n63 VDD1.n62 0.155672
R315 VDD1.n62 VDD1.n10 0.155672
R316 VDD1.n55 VDD1.n10 0.155672
R317 VDD1.n55 VDD1.n54 0.155672
R318 VDD1.n54 VDD1.n14 0.155672
R319 VDD1.n47 VDD1.n14 0.155672
R320 VDD1.n47 VDD1.n46 0.155672
R321 VDD1.n46 VDD1.n18 0.155672
R322 VDD1.n39 VDD1.n18 0.155672
R323 VDD1.n39 VDD1.n38 0.155672
R324 VDD1.n38 VDD1.n22 0.155672
R325 VDD1.n31 VDD1.n22 0.155672
R326 VDD1.n31 VDD1.n30 0.155672
R327 VDD1.n113 VDD1.n112 0.155672
R328 VDD1.n113 VDD1.n104 0.155672
R329 VDD1.n120 VDD1.n104 0.155672
R330 VDD1.n121 VDD1.n120 0.155672
R331 VDD1.n121 VDD1.n100 0.155672
R332 VDD1.n128 VDD1.n100 0.155672
R333 VDD1.n129 VDD1.n128 0.155672
R334 VDD1.n129 VDD1.n96 0.155672
R335 VDD1.n136 VDD1.n96 0.155672
R336 VDD1.n137 VDD1.n136 0.155672
R337 VDD1.n137 VDD1.n92 0.155672
R338 VDD1.n144 VDD1.n92 0.155672
R339 VDD1.n145 VDD1.n144 0.155672
R340 VDD1.n145 VDD1.n88 0.155672
R341 VDD1.n153 VDD1.n88 0.155672
R342 VDD1.n154 VDD1.n153 0.155672
R343 VDD1.n154 VDD1.n84 0.155672
R344 VDD1.n162 VDD1.n84 0.155672
R345 VTAIL.n336 VTAIL.n260 289.615
R346 VTAIL.n78 VTAIL.n2 289.615
R347 VTAIL.n254 VTAIL.n178 289.615
R348 VTAIL.n168 VTAIL.n92 289.615
R349 VTAIL.n287 VTAIL.n286 185
R350 VTAIL.n284 VTAIL.n283 185
R351 VTAIL.n293 VTAIL.n292 185
R352 VTAIL.n295 VTAIL.n294 185
R353 VTAIL.n280 VTAIL.n279 185
R354 VTAIL.n301 VTAIL.n300 185
R355 VTAIL.n303 VTAIL.n302 185
R356 VTAIL.n276 VTAIL.n275 185
R357 VTAIL.n309 VTAIL.n308 185
R358 VTAIL.n311 VTAIL.n310 185
R359 VTAIL.n272 VTAIL.n271 185
R360 VTAIL.n317 VTAIL.n316 185
R361 VTAIL.n319 VTAIL.n318 185
R362 VTAIL.n268 VTAIL.n267 185
R363 VTAIL.n325 VTAIL.n324 185
R364 VTAIL.n328 VTAIL.n327 185
R365 VTAIL.n326 VTAIL.n264 185
R366 VTAIL.n333 VTAIL.n263 185
R367 VTAIL.n335 VTAIL.n334 185
R368 VTAIL.n337 VTAIL.n336 185
R369 VTAIL.n29 VTAIL.n28 185
R370 VTAIL.n26 VTAIL.n25 185
R371 VTAIL.n35 VTAIL.n34 185
R372 VTAIL.n37 VTAIL.n36 185
R373 VTAIL.n22 VTAIL.n21 185
R374 VTAIL.n43 VTAIL.n42 185
R375 VTAIL.n45 VTAIL.n44 185
R376 VTAIL.n18 VTAIL.n17 185
R377 VTAIL.n51 VTAIL.n50 185
R378 VTAIL.n53 VTAIL.n52 185
R379 VTAIL.n14 VTAIL.n13 185
R380 VTAIL.n59 VTAIL.n58 185
R381 VTAIL.n61 VTAIL.n60 185
R382 VTAIL.n10 VTAIL.n9 185
R383 VTAIL.n67 VTAIL.n66 185
R384 VTAIL.n70 VTAIL.n69 185
R385 VTAIL.n68 VTAIL.n6 185
R386 VTAIL.n75 VTAIL.n5 185
R387 VTAIL.n77 VTAIL.n76 185
R388 VTAIL.n79 VTAIL.n78 185
R389 VTAIL.n255 VTAIL.n254 185
R390 VTAIL.n253 VTAIL.n252 185
R391 VTAIL.n251 VTAIL.n181 185
R392 VTAIL.n185 VTAIL.n182 185
R393 VTAIL.n246 VTAIL.n245 185
R394 VTAIL.n244 VTAIL.n243 185
R395 VTAIL.n187 VTAIL.n186 185
R396 VTAIL.n238 VTAIL.n237 185
R397 VTAIL.n236 VTAIL.n235 185
R398 VTAIL.n191 VTAIL.n190 185
R399 VTAIL.n230 VTAIL.n229 185
R400 VTAIL.n228 VTAIL.n227 185
R401 VTAIL.n195 VTAIL.n194 185
R402 VTAIL.n222 VTAIL.n221 185
R403 VTAIL.n220 VTAIL.n219 185
R404 VTAIL.n199 VTAIL.n198 185
R405 VTAIL.n214 VTAIL.n213 185
R406 VTAIL.n212 VTAIL.n211 185
R407 VTAIL.n203 VTAIL.n202 185
R408 VTAIL.n206 VTAIL.n205 185
R409 VTAIL.n169 VTAIL.n168 185
R410 VTAIL.n167 VTAIL.n166 185
R411 VTAIL.n165 VTAIL.n95 185
R412 VTAIL.n99 VTAIL.n96 185
R413 VTAIL.n160 VTAIL.n159 185
R414 VTAIL.n158 VTAIL.n157 185
R415 VTAIL.n101 VTAIL.n100 185
R416 VTAIL.n152 VTAIL.n151 185
R417 VTAIL.n150 VTAIL.n149 185
R418 VTAIL.n105 VTAIL.n104 185
R419 VTAIL.n144 VTAIL.n143 185
R420 VTAIL.n142 VTAIL.n141 185
R421 VTAIL.n109 VTAIL.n108 185
R422 VTAIL.n136 VTAIL.n135 185
R423 VTAIL.n134 VTAIL.n133 185
R424 VTAIL.n113 VTAIL.n112 185
R425 VTAIL.n128 VTAIL.n127 185
R426 VTAIL.n126 VTAIL.n125 185
R427 VTAIL.n117 VTAIL.n116 185
R428 VTAIL.n120 VTAIL.n119 185
R429 VTAIL.t11 VTAIL.n204 147.659
R430 VTAIL.t4 VTAIL.n118 147.659
R431 VTAIL.t6 VTAIL.n285 147.659
R432 VTAIL.t13 VTAIL.n27 147.659
R433 VTAIL.n286 VTAIL.n283 104.615
R434 VTAIL.n293 VTAIL.n283 104.615
R435 VTAIL.n294 VTAIL.n293 104.615
R436 VTAIL.n294 VTAIL.n279 104.615
R437 VTAIL.n301 VTAIL.n279 104.615
R438 VTAIL.n302 VTAIL.n301 104.615
R439 VTAIL.n302 VTAIL.n275 104.615
R440 VTAIL.n309 VTAIL.n275 104.615
R441 VTAIL.n310 VTAIL.n309 104.615
R442 VTAIL.n310 VTAIL.n271 104.615
R443 VTAIL.n317 VTAIL.n271 104.615
R444 VTAIL.n318 VTAIL.n317 104.615
R445 VTAIL.n318 VTAIL.n267 104.615
R446 VTAIL.n325 VTAIL.n267 104.615
R447 VTAIL.n327 VTAIL.n325 104.615
R448 VTAIL.n327 VTAIL.n326 104.615
R449 VTAIL.n326 VTAIL.n263 104.615
R450 VTAIL.n335 VTAIL.n263 104.615
R451 VTAIL.n336 VTAIL.n335 104.615
R452 VTAIL.n28 VTAIL.n25 104.615
R453 VTAIL.n35 VTAIL.n25 104.615
R454 VTAIL.n36 VTAIL.n35 104.615
R455 VTAIL.n36 VTAIL.n21 104.615
R456 VTAIL.n43 VTAIL.n21 104.615
R457 VTAIL.n44 VTAIL.n43 104.615
R458 VTAIL.n44 VTAIL.n17 104.615
R459 VTAIL.n51 VTAIL.n17 104.615
R460 VTAIL.n52 VTAIL.n51 104.615
R461 VTAIL.n52 VTAIL.n13 104.615
R462 VTAIL.n59 VTAIL.n13 104.615
R463 VTAIL.n60 VTAIL.n59 104.615
R464 VTAIL.n60 VTAIL.n9 104.615
R465 VTAIL.n67 VTAIL.n9 104.615
R466 VTAIL.n69 VTAIL.n67 104.615
R467 VTAIL.n69 VTAIL.n68 104.615
R468 VTAIL.n68 VTAIL.n5 104.615
R469 VTAIL.n77 VTAIL.n5 104.615
R470 VTAIL.n78 VTAIL.n77 104.615
R471 VTAIL.n254 VTAIL.n253 104.615
R472 VTAIL.n253 VTAIL.n181 104.615
R473 VTAIL.n185 VTAIL.n181 104.615
R474 VTAIL.n245 VTAIL.n185 104.615
R475 VTAIL.n245 VTAIL.n244 104.615
R476 VTAIL.n244 VTAIL.n186 104.615
R477 VTAIL.n237 VTAIL.n186 104.615
R478 VTAIL.n237 VTAIL.n236 104.615
R479 VTAIL.n236 VTAIL.n190 104.615
R480 VTAIL.n229 VTAIL.n190 104.615
R481 VTAIL.n229 VTAIL.n228 104.615
R482 VTAIL.n228 VTAIL.n194 104.615
R483 VTAIL.n221 VTAIL.n194 104.615
R484 VTAIL.n221 VTAIL.n220 104.615
R485 VTAIL.n220 VTAIL.n198 104.615
R486 VTAIL.n213 VTAIL.n198 104.615
R487 VTAIL.n213 VTAIL.n212 104.615
R488 VTAIL.n212 VTAIL.n202 104.615
R489 VTAIL.n205 VTAIL.n202 104.615
R490 VTAIL.n168 VTAIL.n167 104.615
R491 VTAIL.n167 VTAIL.n95 104.615
R492 VTAIL.n99 VTAIL.n95 104.615
R493 VTAIL.n159 VTAIL.n99 104.615
R494 VTAIL.n159 VTAIL.n158 104.615
R495 VTAIL.n158 VTAIL.n100 104.615
R496 VTAIL.n151 VTAIL.n100 104.615
R497 VTAIL.n151 VTAIL.n150 104.615
R498 VTAIL.n150 VTAIL.n104 104.615
R499 VTAIL.n143 VTAIL.n104 104.615
R500 VTAIL.n143 VTAIL.n142 104.615
R501 VTAIL.n142 VTAIL.n108 104.615
R502 VTAIL.n135 VTAIL.n108 104.615
R503 VTAIL.n135 VTAIL.n134 104.615
R504 VTAIL.n134 VTAIL.n112 104.615
R505 VTAIL.n127 VTAIL.n112 104.615
R506 VTAIL.n127 VTAIL.n126 104.615
R507 VTAIL.n126 VTAIL.n116 104.615
R508 VTAIL.n119 VTAIL.n116 104.615
R509 VTAIL.n286 VTAIL.t6 52.3082
R510 VTAIL.n28 VTAIL.t13 52.3082
R511 VTAIL.n205 VTAIL.t11 52.3082
R512 VTAIL.n119 VTAIL.t4 52.3082
R513 VTAIL.n177 VTAIL.n176 48.509
R514 VTAIL.n175 VTAIL.n174 48.509
R515 VTAIL.n91 VTAIL.n90 48.509
R516 VTAIL.n89 VTAIL.n88 48.509
R517 VTAIL.n343 VTAIL.n342 48.5088
R518 VTAIL.n1 VTAIL.n0 48.5088
R519 VTAIL.n85 VTAIL.n84 48.5088
R520 VTAIL.n87 VTAIL.n86 48.5088
R521 VTAIL.n341 VTAIL.n340 36.452
R522 VTAIL.n83 VTAIL.n82 36.452
R523 VTAIL.n259 VTAIL.n258 36.452
R524 VTAIL.n173 VTAIL.n172 36.452
R525 VTAIL.n89 VTAIL.n87 28.091
R526 VTAIL.n341 VTAIL.n259 26.6341
R527 VTAIL.n287 VTAIL.n285 15.6677
R528 VTAIL.n29 VTAIL.n27 15.6677
R529 VTAIL.n206 VTAIL.n204 15.6677
R530 VTAIL.n120 VTAIL.n118 15.6677
R531 VTAIL.n334 VTAIL.n333 13.1884
R532 VTAIL.n76 VTAIL.n75 13.1884
R533 VTAIL.n252 VTAIL.n251 13.1884
R534 VTAIL.n166 VTAIL.n165 13.1884
R535 VTAIL.n288 VTAIL.n284 12.8005
R536 VTAIL.n332 VTAIL.n264 12.8005
R537 VTAIL.n337 VTAIL.n262 12.8005
R538 VTAIL.n30 VTAIL.n26 12.8005
R539 VTAIL.n74 VTAIL.n6 12.8005
R540 VTAIL.n79 VTAIL.n4 12.8005
R541 VTAIL.n255 VTAIL.n180 12.8005
R542 VTAIL.n250 VTAIL.n182 12.8005
R543 VTAIL.n207 VTAIL.n203 12.8005
R544 VTAIL.n169 VTAIL.n94 12.8005
R545 VTAIL.n164 VTAIL.n96 12.8005
R546 VTAIL.n121 VTAIL.n117 12.8005
R547 VTAIL.n292 VTAIL.n291 12.0247
R548 VTAIL.n329 VTAIL.n328 12.0247
R549 VTAIL.n338 VTAIL.n260 12.0247
R550 VTAIL.n34 VTAIL.n33 12.0247
R551 VTAIL.n71 VTAIL.n70 12.0247
R552 VTAIL.n80 VTAIL.n2 12.0247
R553 VTAIL.n256 VTAIL.n178 12.0247
R554 VTAIL.n247 VTAIL.n246 12.0247
R555 VTAIL.n211 VTAIL.n210 12.0247
R556 VTAIL.n170 VTAIL.n92 12.0247
R557 VTAIL.n161 VTAIL.n160 12.0247
R558 VTAIL.n125 VTAIL.n124 12.0247
R559 VTAIL.n295 VTAIL.n282 11.249
R560 VTAIL.n324 VTAIL.n266 11.249
R561 VTAIL.n37 VTAIL.n24 11.249
R562 VTAIL.n66 VTAIL.n8 11.249
R563 VTAIL.n243 VTAIL.n184 11.249
R564 VTAIL.n214 VTAIL.n201 11.249
R565 VTAIL.n157 VTAIL.n98 11.249
R566 VTAIL.n128 VTAIL.n115 11.249
R567 VTAIL.n296 VTAIL.n280 10.4732
R568 VTAIL.n323 VTAIL.n268 10.4732
R569 VTAIL.n38 VTAIL.n22 10.4732
R570 VTAIL.n65 VTAIL.n10 10.4732
R571 VTAIL.n242 VTAIL.n187 10.4732
R572 VTAIL.n215 VTAIL.n199 10.4732
R573 VTAIL.n156 VTAIL.n101 10.4732
R574 VTAIL.n129 VTAIL.n113 10.4732
R575 VTAIL.n300 VTAIL.n299 9.69747
R576 VTAIL.n320 VTAIL.n319 9.69747
R577 VTAIL.n42 VTAIL.n41 9.69747
R578 VTAIL.n62 VTAIL.n61 9.69747
R579 VTAIL.n239 VTAIL.n238 9.69747
R580 VTAIL.n219 VTAIL.n218 9.69747
R581 VTAIL.n153 VTAIL.n152 9.69747
R582 VTAIL.n133 VTAIL.n132 9.69747
R583 VTAIL.n340 VTAIL.n339 9.45567
R584 VTAIL.n82 VTAIL.n81 9.45567
R585 VTAIL.n258 VTAIL.n257 9.45567
R586 VTAIL.n172 VTAIL.n171 9.45567
R587 VTAIL.n339 VTAIL.n338 9.3005
R588 VTAIL.n262 VTAIL.n261 9.3005
R589 VTAIL.n307 VTAIL.n306 9.3005
R590 VTAIL.n305 VTAIL.n304 9.3005
R591 VTAIL.n278 VTAIL.n277 9.3005
R592 VTAIL.n299 VTAIL.n298 9.3005
R593 VTAIL.n297 VTAIL.n296 9.3005
R594 VTAIL.n282 VTAIL.n281 9.3005
R595 VTAIL.n291 VTAIL.n290 9.3005
R596 VTAIL.n289 VTAIL.n288 9.3005
R597 VTAIL.n274 VTAIL.n273 9.3005
R598 VTAIL.n313 VTAIL.n312 9.3005
R599 VTAIL.n315 VTAIL.n314 9.3005
R600 VTAIL.n270 VTAIL.n269 9.3005
R601 VTAIL.n321 VTAIL.n320 9.3005
R602 VTAIL.n323 VTAIL.n322 9.3005
R603 VTAIL.n266 VTAIL.n265 9.3005
R604 VTAIL.n330 VTAIL.n329 9.3005
R605 VTAIL.n332 VTAIL.n331 9.3005
R606 VTAIL.n81 VTAIL.n80 9.3005
R607 VTAIL.n4 VTAIL.n3 9.3005
R608 VTAIL.n49 VTAIL.n48 9.3005
R609 VTAIL.n47 VTAIL.n46 9.3005
R610 VTAIL.n20 VTAIL.n19 9.3005
R611 VTAIL.n41 VTAIL.n40 9.3005
R612 VTAIL.n39 VTAIL.n38 9.3005
R613 VTAIL.n24 VTAIL.n23 9.3005
R614 VTAIL.n33 VTAIL.n32 9.3005
R615 VTAIL.n31 VTAIL.n30 9.3005
R616 VTAIL.n16 VTAIL.n15 9.3005
R617 VTAIL.n55 VTAIL.n54 9.3005
R618 VTAIL.n57 VTAIL.n56 9.3005
R619 VTAIL.n12 VTAIL.n11 9.3005
R620 VTAIL.n63 VTAIL.n62 9.3005
R621 VTAIL.n65 VTAIL.n64 9.3005
R622 VTAIL.n8 VTAIL.n7 9.3005
R623 VTAIL.n72 VTAIL.n71 9.3005
R624 VTAIL.n74 VTAIL.n73 9.3005
R625 VTAIL.n232 VTAIL.n231 9.3005
R626 VTAIL.n234 VTAIL.n233 9.3005
R627 VTAIL.n189 VTAIL.n188 9.3005
R628 VTAIL.n240 VTAIL.n239 9.3005
R629 VTAIL.n242 VTAIL.n241 9.3005
R630 VTAIL.n184 VTAIL.n183 9.3005
R631 VTAIL.n248 VTAIL.n247 9.3005
R632 VTAIL.n250 VTAIL.n249 9.3005
R633 VTAIL.n257 VTAIL.n256 9.3005
R634 VTAIL.n180 VTAIL.n179 9.3005
R635 VTAIL.n193 VTAIL.n192 9.3005
R636 VTAIL.n226 VTAIL.n225 9.3005
R637 VTAIL.n224 VTAIL.n223 9.3005
R638 VTAIL.n197 VTAIL.n196 9.3005
R639 VTAIL.n218 VTAIL.n217 9.3005
R640 VTAIL.n216 VTAIL.n215 9.3005
R641 VTAIL.n201 VTAIL.n200 9.3005
R642 VTAIL.n210 VTAIL.n209 9.3005
R643 VTAIL.n208 VTAIL.n207 9.3005
R644 VTAIL.n146 VTAIL.n145 9.3005
R645 VTAIL.n148 VTAIL.n147 9.3005
R646 VTAIL.n103 VTAIL.n102 9.3005
R647 VTAIL.n154 VTAIL.n153 9.3005
R648 VTAIL.n156 VTAIL.n155 9.3005
R649 VTAIL.n98 VTAIL.n97 9.3005
R650 VTAIL.n162 VTAIL.n161 9.3005
R651 VTAIL.n164 VTAIL.n163 9.3005
R652 VTAIL.n171 VTAIL.n170 9.3005
R653 VTAIL.n94 VTAIL.n93 9.3005
R654 VTAIL.n107 VTAIL.n106 9.3005
R655 VTAIL.n140 VTAIL.n139 9.3005
R656 VTAIL.n138 VTAIL.n137 9.3005
R657 VTAIL.n111 VTAIL.n110 9.3005
R658 VTAIL.n132 VTAIL.n131 9.3005
R659 VTAIL.n130 VTAIL.n129 9.3005
R660 VTAIL.n115 VTAIL.n114 9.3005
R661 VTAIL.n124 VTAIL.n123 9.3005
R662 VTAIL.n122 VTAIL.n121 9.3005
R663 VTAIL.n303 VTAIL.n278 8.92171
R664 VTAIL.n316 VTAIL.n270 8.92171
R665 VTAIL.n45 VTAIL.n20 8.92171
R666 VTAIL.n58 VTAIL.n12 8.92171
R667 VTAIL.n235 VTAIL.n189 8.92171
R668 VTAIL.n222 VTAIL.n197 8.92171
R669 VTAIL.n149 VTAIL.n103 8.92171
R670 VTAIL.n136 VTAIL.n111 8.92171
R671 VTAIL.n304 VTAIL.n276 8.14595
R672 VTAIL.n315 VTAIL.n272 8.14595
R673 VTAIL.n46 VTAIL.n18 8.14595
R674 VTAIL.n57 VTAIL.n14 8.14595
R675 VTAIL.n234 VTAIL.n191 8.14595
R676 VTAIL.n223 VTAIL.n195 8.14595
R677 VTAIL.n148 VTAIL.n105 8.14595
R678 VTAIL.n137 VTAIL.n109 8.14595
R679 VTAIL.n308 VTAIL.n307 7.3702
R680 VTAIL.n312 VTAIL.n311 7.3702
R681 VTAIL.n50 VTAIL.n49 7.3702
R682 VTAIL.n54 VTAIL.n53 7.3702
R683 VTAIL.n231 VTAIL.n230 7.3702
R684 VTAIL.n227 VTAIL.n226 7.3702
R685 VTAIL.n145 VTAIL.n144 7.3702
R686 VTAIL.n141 VTAIL.n140 7.3702
R687 VTAIL.n308 VTAIL.n274 6.59444
R688 VTAIL.n311 VTAIL.n274 6.59444
R689 VTAIL.n50 VTAIL.n16 6.59444
R690 VTAIL.n53 VTAIL.n16 6.59444
R691 VTAIL.n230 VTAIL.n193 6.59444
R692 VTAIL.n227 VTAIL.n193 6.59444
R693 VTAIL.n144 VTAIL.n107 6.59444
R694 VTAIL.n141 VTAIL.n107 6.59444
R695 VTAIL.n307 VTAIL.n276 5.81868
R696 VTAIL.n312 VTAIL.n272 5.81868
R697 VTAIL.n49 VTAIL.n18 5.81868
R698 VTAIL.n54 VTAIL.n14 5.81868
R699 VTAIL.n231 VTAIL.n191 5.81868
R700 VTAIL.n226 VTAIL.n195 5.81868
R701 VTAIL.n145 VTAIL.n105 5.81868
R702 VTAIL.n140 VTAIL.n109 5.81868
R703 VTAIL.n304 VTAIL.n303 5.04292
R704 VTAIL.n316 VTAIL.n315 5.04292
R705 VTAIL.n46 VTAIL.n45 5.04292
R706 VTAIL.n58 VTAIL.n57 5.04292
R707 VTAIL.n235 VTAIL.n234 5.04292
R708 VTAIL.n223 VTAIL.n222 5.04292
R709 VTAIL.n149 VTAIL.n148 5.04292
R710 VTAIL.n137 VTAIL.n136 5.04292
R711 VTAIL.n208 VTAIL.n204 4.38563
R712 VTAIL.n122 VTAIL.n118 4.38563
R713 VTAIL.n289 VTAIL.n285 4.38563
R714 VTAIL.n31 VTAIL.n27 4.38563
R715 VTAIL.n300 VTAIL.n278 4.26717
R716 VTAIL.n319 VTAIL.n270 4.26717
R717 VTAIL.n42 VTAIL.n20 4.26717
R718 VTAIL.n61 VTAIL.n12 4.26717
R719 VTAIL.n238 VTAIL.n189 4.26717
R720 VTAIL.n219 VTAIL.n197 4.26717
R721 VTAIL.n152 VTAIL.n103 4.26717
R722 VTAIL.n133 VTAIL.n111 4.26717
R723 VTAIL.n299 VTAIL.n280 3.49141
R724 VTAIL.n320 VTAIL.n268 3.49141
R725 VTAIL.n41 VTAIL.n22 3.49141
R726 VTAIL.n62 VTAIL.n10 3.49141
R727 VTAIL.n239 VTAIL.n187 3.49141
R728 VTAIL.n218 VTAIL.n199 3.49141
R729 VTAIL.n153 VTAIL.n101 3.49141
R730 VTAIL.n132 VTAIL.n113 3.49141
R731 VTAIL.n296 VTAIL.n295 2.71565
R732 VTAIL.n324 VTAIL.n323 2.71565
R733 VTAIL.n38 VTAIL.n37 2.71565
R734 VTAIL.n66 VTAIL.n65 2.71565
R735 VTAIL.n243 VTAIL.n242 2.71565
R736 VTAIL.n215 VTAIL.n214 2.71565
R737 VTAIL.n157 VTAIL.n156 2.71565
R738 VTAIL.n129 VTAIL.n128 2.71565
R739 VTAIL.n292 VTAIL.n282 1.93989
R740 VTAIL.n328 VTAIL.n266 1.93989
R741 VTAIL.n340 VTAIL.n260 1.93989
R742 VTAIL.n34 VTAIL.n24 1.93989
R743 VTAIL.n70 VTAIL.n8 1.93989
R744 VTAIL.n82 VTAIL.n2 1.93989
R745 VTAIL.n258 VTAIL.n178 1.93989
R746 VTAIL.n246 VTAIL.n184 1.93989
R747 VTAIL.n211 VTAIL.n201 1.93989
R748 VTAIL.n172 VTAIL.n92 1.93989
R749 VTAIL.n160 VTAIL.n98 1.93989
R750 VTAIL.n125 VTAIL.n115 1.93989
R751 VTAIL.n91 VTAIL.n89 1.4574
R752 VTAIL.n173 VTAIL.n91 1.4574
R753 VTAIL.n177 VTAIL.n175 1.4574
R754 VTAIL.n259 VTAIL.n177 1.4574
R755 VTAIL.n87 VTAIL.n85 1.4574
R756 VTAIL.n85 VTAIL.n83 1.4574
R757 VTAIL.n343 VTAIL.n341 1.4574
R758 VTAIL.n342 VTAIL.t0 1.33294
R759 VTAIL.n342 VTAIL.t3 1.33294
R760 VTAIL.n0 VTAIL.t7 1.33294
R761 VTAIL.n0 VTAIL.t1 1.33294
R762 VTAIL.n84 VTAIL.t10 1.33294
R763 VTAIL.n84 VTAIL.t19 1.33294
R764 VTAIL.n86 VTAIL.t14 1.33294
R765 VTAIL.n86 VTAIL.t16 1.33294
R766 VTAIL.n176 VTAIL.t17 1.33294
R767 VTAIL.n176 VTAIL.t18 1.33294
R768 VTAIL.n174 VTAIL.t12 1.33294
R769 VTAIL.n174 VTAIL.t15 1.33294
R770 VTAIL.n90 VTAIL.t2 1.33294
R771 VTAIL.n90 VTAIL.t8 1.33294
R772 VTAIL.n88 VTAIL.t9 1.33294
R773 VTAIL.n88 VTAIL.t5 1.33294
R774 VTAIL.n175 VTAIL.n173 1.19878
R775 VTAIL.n83 VTAIL.n1 1.19878
R776 VTAIL.n291 VTAIL.n284 1.16414
R777 VTAIL.n329 VTAIL.n264 1.16414
R778 VTAIL.n338 VTAIL.n337 1.16414
R779 VTAIL.n33 VTAIL.n26 1.16414
R780 VTAIL.n71 VTAIL.n6 1.16414
R781 VTAIL.n80 VTAIL.n79 1.16414
R782 VTAIL.n256 VTAIL.n255 1.16414
R783 VTAIL.n247 VTAIL.n182 1.16414
R784 VTAIL.n210 VTAIL.n203 1.16414
R785 VTAIL.n170 VTAIL.n169 1.16414
R786 VTAIL.n161 VTAIL.n96 1.16414
R787 VTAIL.n124 VTAIL.n117 1.16414
R788 VTAIL VTAIL.n1 1.15136
R789 VTAIL.n288 VTAIL.n287 0.388379
R790 VTAIL.n333 VTAIL.n332 0.388379
R791 VTAIL.n334 VTAIL.n262 0.388379
R792 VTAIL.n30 VTAIL.n29 0.388379
R793 VTAIL.n75 VTAIL.n74 0.388379
R794 VTAIL.n76 VTAIL.n4 0.388379
R795 VTAIL.n252 VTAIL.n180 0.388379
R796 VTAIL.n251 VTAIL.n250 0.388379
R797 VTAIL.n207 VTAIL.n206 0.388379
R798 VTAIL.n166 VTAIL.n94 0.388379
R799 VTAIL.n165 VTAIL.n164 0.388379
R800 VTAIL.n121 VTAIL.n120 0.388379
R801 VTAIL VTAIL.n343 0.306534
R802 VTAIL.n290 VTAIL.n289 0.155672
R803 VTAIL.n290 VTAIL.n281 0.155672
R804 VTAIL.n297 VTAIL.n281 0.155672
R805 VTAIL.n298 VTAIL.n297 0.155672
R806 VTAIL.n298 VTAIL.n277 0.155672
R807 VTAIL.n305 VTAIL.n277 0.155672
R808 VTAIL.n306 VTAIL.n305 0.155672
R809 VTAIL.n306 VTAIL.n273 0.155672
R810 VTAIL.n313 VTAIL.n273 0.155672
R811 VTAIL.n314 VTAIL.n313 0.155672
R812 VTAIL.n314 VTAIL.n269 0.155672
R813 VTAIL.n321 VTAIL.n269 0.155672
R814 VTAIL.n322 VTAIL.n321 0.155672
R815 VTAIL.n322 VTAIL.n265 0.155672
R816 VTAIL.n330 VTAIL.n265 0.155672
R817 VTAIL.n331 VTAIL.n330 0.155672
R818 VTAIL.n331 VTAIL.n261 0.155672
R819 VTAIL.n339 VTAIL.n261 0.155672
R820 VTAIL.n32 VTAIL.n31 0.155672
R821 VTAIL.n32 VTAIL.n23 0.155672
R822 VTAIL.n39 VTAIL.n23 0.155672
R823 VTAIL.n40 VTAIL.n39 0.155672
R824 VTAIL.n40 VTAIL.n19 0.155672
R825 VTAIL.n47 VTAIL.n19 0.155672
R826 VTAIL.n48 VTAIL.n47 0.155672
R827 VTAIL.n48 VTAIL.n15 0.155672
R828 VTAIL.n55 VTAIL.n15 0.155672
R829 VTAIL.n56 VTAIL.n55 0.155672
R830 VTAIL.n56 VTAIL.n11 0.155672
R831 VTAIL.n63 VTAIL.n11 0.155672
R832 VTAIL.n64 VTAIL.n63 0.155672
R833 VTAIL.n64 VTAIL.n7 0.155672
R834 VTAIL.n72 VTAIL.n7 0.155672
R835 VTAIL.n73 VTAIL.n72 0.155672
R836 VTAIL.n73 VTAIL.n3 0.155672
R837 VTAIL.n81 VTAIL.n3 0.155672
R838 VTAIL.n257 VTAIL.n179 0.155672
R839 VTAIL.n249 VTAIL.n179 0.155672
R840 VTAIL.n249 VTAIL.n248 0.155672
R841 VTAIL.n248 VTAIL.n183 0.155672
R842 VTAIL.n241 VTAIL.n183 0.155672
R843 VTAIL.n241 VTAIL.n240 0.155672
R844 VTAIL.n240 VTAIL.n188 0.155672
R845 VTAIL.n233 VTAIL.n188 0.155672
R846 VTAIL.n233 VTAIL.n232 0.155672
R847 VTAIL.n232 VTAIL.n192 0.155672
R848 VTAIL.n225 VTAIL.n192 0.155672
R849 VTAIL.n225 VTAIL.n224 0.155672
R850 VTAIL.n224 VTAIL.n196 0.155672
R851 VTAIL.n217 VTAIL.n196 0.155672
R852 VTAIL.n217 VTAIL.n216 0.155672
R853 VTAIL.n216 VTAIL.n200 0.155672
R854 VTAIL.n209 VTAIL.n200 0.155672
R855 VTAIL.n209 VTAIL.n208 0.155672
R856 VTAIL.n171 VTAIL.n93 0.155672
R857 VTAIL.n163 VTAIL.n93 0.155672
R858 VTAIL.n163 VTAIL.n162 0.155672
R859 VTAIL.n162 VTAIL.n97 0.155672
R860 VTAIL.n155 VTAIL.n97 0.155672
R861 VTAIL.n155 VTAIL.n154 0.155672
R862 VTAIL.n154 VTAIL.n102 0.155672
R863 VTAIL.n147 VTAIL.n102 0.155672
R864 VTAIL.n147 VTAIL.n146 0.155672
R865 VTAIL.n146 VTAIL.n106 0.155672
R866 VTAIL.n139 VTAIL.n106 0.155672
R867 VTAIL.n139 VTAIL.n138 0.155672
R868 VTAIL.n138 VTAIL.n110 0.155672
R869 VTAIL.n131 VTAIL.n110 0.155672
R870 VTAIL.n131 VTAIL.n130 0.155672
R871 VTAIL.n130 VTAIL.n114 0.155672
R872 VTAIL.n123 VTAIL.n114 0.155672
R873 VTAIL.n123 VTAIL.n122 0.155672
R874 B.n649 B.n648 585
R875 B.n650 B.n131 585
R876 B.n652 B.n651 585
R877 B.n654 B.n130 585
R878 B.n657 B.n656 585
R879 B.n658 B.n129 585
R880 B.n660 B.n659 585
R881 B.n662 B.n128 585
R882 B.n665 B.n664 585
R883 B.n666 B.n127 585
R884 B.n668 B.n667 585
R885 B.n670 B.n126 585
R886 B.n673 B.n672 585
R887 B.n674 B.n125 585
R888 B.n676 B.n675 585
R889 B.n678 B.n124 585
R890 B.n681 B.n680 585
R891 B.n682 B.n123 585
R892 B.n684 B.n683 585
R893 B.n686 B.n122 585
R894 B.n689 B.n688 585
R895 B.n690 B.n121 585
R896 B.n692 B.n691 585
R897 B.n694 B.n120 585
R898 B.n697 B.n696 585
R899 B.n698 B.n119 585
R900 B.n700 B.n699 585
R901 B.n702 B.n118 585
R902 B.n705 B.n704 585
R903 B.n706 B.n117 585
R904 B.n708 B.n707 585
R905 B.n710 B.n116 585
R906 B.n713 B.n712 585
R907 B.n714 B.n115 585
R908 B.n716 B.n715 585
R909 B.n718 B.n114 585
R910 B.n721 B.n720 585
R911 B.n722 B.n113 585
R912 B.n724 B.n723 585
R913 B.n726 B.n112 585
R914 B.n729 B.n728 585
R915 B.n730 B.n111 585
R916 B.n732 B.n731 585
R917 B.n734 B.n110 585
R918 B.n737 B.n736 585
R919 B.n738 B.n109 585
R920 B.n740 B.n739 585
R921 B.n742 B.n108 585
R922 B.n744 B.n743 585
R923 B.n746 B.n745 585
R924 B.n749 B.n748 585
R925 B.n750 B.n103 585
R926 B.n752 B.n751 585
R927 B.n754 B.n102 585
R928 B.n757 B.n756 585
R929 B.n758 B.n101 585
R930 B.n760 B.n759 585
R931 B.n762 B.n100 585
R932 B.n764 B.n763 585
R933 B.n766 B.n765 585
R934 B.n769 B.n768 585
R935 B.n770 B.n95 585
R936 B.n772 B.n771 585
R937 B.n774 B.n94 585
R938 B.n777 B.n776 585
R939 B.n778 B.n93 585
R940 B.n780 B.n779 585
R941 B.n782 B.n92 585
R942 B.n785 B.n784 585
R943 B.n786 B.n91 585
R944 B.n788 B.n787 585
R945 B.n790 B.n90 585
R946 B.n793 B.n792 585
R947 B.n794 B.n89 585
R948 B.n796 B.n795 585
R949 B.n798 B.n88 585
R950 B.n801 B.n800 585
R951 B.n802 B.n87 585
R952 B.n804 B.n803 585
R953 B.n806 B.n86 585
R954 B.n809 B.n808 585
R955 B.n810 B.n85 585
R956 B.n812 B.n811 585
R957 B.n814 B.n84 585
R958 B.n817 B.n816 585
R959 B.n818 B.n83 585
R960 B.n820 B.n819 585
R961 B.n822 B.n82 585
R962 B.n825 B.n824 585
R963 B.n826 B.n81 585
R964 B.n828 B.n827 585
R965 B.n830 B.n80 585
R966 B.n833 B.n832 585
R967 B.n834 B.n79 585
R968 B.n836 B.n835 585
R969 B.n838 B.n78 585
R970 B.n841 B.n840 585
R971 B.n842 B.n77 585
R972 B.n844 B.n843 585
R973 B.n846 B.n76 585
R974 B.n849 B.n848 585
R975 B.n850 B.n75 585
R976 B.n852 B.n851 585
R977 B.n854 B.n74 585
R978 B.n857 B.n856 585
R979 B.n858 B.n73 585
R980 B.n860 B.n859 585
R981 B.n862 B.n72 585
R982 B.n865 B.n864 585
R983 B.n866 B.n71 585
R984 B.n646 B.n69 585
R985 B.n869 B.n69 585
R986 B.n645 B.n68 585
R987 B.n870 B.n68 585
R988 B.n644 B.n67 585
R989 B.n871 B.n67 585
R990 B.n643 B.n642 585
R991 B.n642 B.n63 585
R992 B.n641 B.n62 585
R993 B.n877 B.n62 585
R994 B.n640 B.n61 585
R995 B.n878 B.n61 585
R996 B.n639 B.n60 585
R997 B.n879 B.n60 585
R998 B.n638 B.n637 585
R999 B.n637 B.n56 585
R1000 B.n636 B.n55 585
R1001 B.n885 B.n55 585
R1002 B.n635 B.n54 585
R1003 B.n886 B.n54 585
R1004 B.n634 B.n53 585
R1005 B.n887 B.n53 585
R1006 B.n633 B.n632 585
R1007 B.n632 B.n49 585
R1008 B.n631 B.n48 585
R1009 B.n893 B.n48 585
R1010 B.n630 B.n47 585
R1011 B.n894 B.n47 585
R1012 B.n629 B.n46 585
R1013 B.n895 B.n46 585
R1014 B.n628 B.n627 585
R1015 B.n627 B.n42 585
R1016 B.n626 B.n41 585
R1017 B.n901 B.n41 585
R1018 B.n625 B.n40 585
R1019 B.n902 B.n40 585
R1020 B.n624 B.n39 585
R1021 B.n903 B.n39 585
R1022 B.n623 B.n622 585
R1023 B.n622 B.t3 585
R1024 B.n621 B.n35 585
R1025 B.n909 B.n35 585
R1026 B.n620 B.n34 585
R1027 B.n910 B.n34 585
R1028 B.n619 B.n33 585
R1029 B.n911 B.n33 585
R1030 B.n618 B.n617 585
R1031 B.n617 B.n32 585
R1032 B.n616 B.n28 585
R1033 B.n917 B.n28 585
R1034 B.n615 B.n27 585
R1035 B.n918 B.n27 585
R1036 B.n614 B.n26 585
R1037 B.n919 B.n26 585
R1038 B.n613 B.n612 585
R1039 B.n612 B.n22 585
R1040 B.n611 B.n21 585
R1041 B.n925 B.n21 585
R1042 B.n610 B.n20 585
R1043 B.n926 B.n20 585
R1044 B.n609 B.n19 585
R1045 B.n927 B.n19 585
R1046 B.n608 B.n607 585
R1047 B.n607 B.n15 585
R1048 B.n606 B.n14 585
R1049 B.n933 B.n14 585
R1050 B.n605 B.n13 585
R1051 B.n934 B.n13 585
R1052 B.n604 B.n12 585
R1053 B.n935 B.n12 585
R1054 B.n603 B.n602 585
R1055 B.n602 B.n8 585
R1056 B.n601 B.n7 585
R1057 B.n941 B.n7 585
R1058 B.n600 B.n6 585
R1059 B.n942 B.n6 585
R1060 B.n599 B.n5 585
R1061 B.n943 B.n5 585
R1062 B.n598 B.n597 585
R1063 B.n597 B.n4 585
R1064 B.n596 B.n132 585
R1065 B.n596 B.n595 585
R1066 B.n586 B.n133 585
R1067 B.n134 B.n133 585
R1068 B.n588 B.n587 585
R1069 B.n589 B.n588 585
R1070 B.n585 B.n138 585
R1071 B.n142 B.n138 585
R1072 B.n584 B.n583 585
R1073 B.n583 B.n582 585
R1074 B.n140 B.n139 585
R1075 B.n141 B.n140 585
R1076 B.n575 B.n574 585
R1077 B.n576 B.n575 585
R1078 B.n573 B.n147 585
R1079 B.n147 B.n146 585
R1080 B.n572 B.n571 585
R1081 B.n571 B.n570 585
R1082 B.n149 B.n148 585
R1083 B.n150 B.n149 585
R1084 B.n563 B.n562 585
R1085 B.n564 B.n563 585
R1086 B.n561 B.n155 585
R1087 B.n155 B.n154 585
R1088 B.n560 B.n559 585
R1089 B.n559 B.n558 585
R1090 B.n157 B.n156 585
R1091 B.n551 B.n157 585
R1092 B.n550 B.n549 585
R1093 B.n552 B.n550 585
R1094 B.n548 B.n162 585
R1095 B.n162 B.n161 585
R1096 B.n547 B.n546 585
R1097 B.n546 B.n545 585
R1098 B.n164 B.n163 585
R1099 B.t5 B.n164 585
R1100 B.n538 B.n537 585
R1101 B.n539 B.n538 585
R1102 B.n536 B.n169 585
R1103 B.n169 B.n168 585
R1104 B.n535 B.n534 585
R1105 B.n534 B.n533 585
R1106 B.n171 B.n170 585
R1107 B.n172 B.n171 585
R1108 B.n526 B.n525 585
R1109 B.n527 B.n526 585
R1110 B.n524 B.n177 585
R1111 B.n177 B.n176 585
R1112 B.n523 B.n522 585
R1113 B.n522 B.n521 585
R1114 B.n179 B.n178 585
R1115 B.n180 B.n179 585
R1116 B.n514 B.n513 585
R1117 B.n515 B.n514 585
R1118 B.n512 B.n185 585
R1119 B.n185 B.n184 585
R1120 B.n511 B.n510 585
R1121 B.n510 B.n509 585
R1122 B.n187 B.n186 585
R1123 B.n188 B.n187 585
R1124 B.n502 B.n501 585
R1125 B.n503 B.n502 585
R1126 B.n500 B.n192 585
R1127 B.n196 B.n192 585
R1128 B.n499 B.n498 585
R1129 B.n498 B.n497 585
R1130 B.n194 B.n193 585
R1131 B.n195 B.n194 585
R1132 B.n490 B.n489 585
R1133 B.n491 B.n490 585
R1134 B.n488 B.n201 585
R1135 B.n201 B.n200 585
R1136 B.n487 B.n486 585
R1137 B.n486 B.n485 585
R1138 B.n482 B.n205 585
R1139 B.n481 B.n480 585
R1140 B.n478 B.n206 585
R1141 B.n478 B.n204 585
R1142 B.n477 B.n476 585
R1143 B.n475 B.n474 585
R1144 B.n473 B.n208 585
R1145 B.n471 B.n470 585
R1146 B.n469 B.n209 585
R1147 B.n468 B.n467 585
R1148 B.n465 B.n210 585
R1149 B.n463 B.n462 585
R1150 B.n461 B.n211 585
R1151 B.n460 B.n459 585
R1152 B.n457 B.n212 585
R1153 B.n455 B.n454 585
R1154 B.n453 B.n213 585
R1155 B.n452 B.n451 585
R1156 B.n449 B.n214 585
R1157 B.n447 B.n446 585
R1158 B.n445 B.n215 585
R1159 B.n444 B.n443 585
R1160 B.n441 B.n216 585
R1161 B.n439 B.n438 585
R1162 B.n437 B.n217 585
R1163 B.n436 B.n435 585
R1164 B.n433 B.n218 585
R1165 B.n431 B.n430 585
R1166 B.n429 B.n219 585
R1167 B.n428 B.n427 585
R1168 B.n425 B.n220 585
R1169 B.n423 B.n422 585
R1170 B.n421 B.n221 585
R1171 B.n420 B.n419 585
R1172 B.n417 B.n222 585
R1173 B.n415 B.n414 585
R1174 B.n413 B.n223 585
R1175 B.n412 B.n411 585
R1176 B.n409 B.n224 585
R1177 B.n407 B.n406 585
R1178 B.n405 B.n225 585
R1179 B.n404 B.n403 585
R1180 B.n401 B.n226 585
R1181 B.n399 B.n398 585
R1182 B.n397 B.n227 585
R1183 B.n396 B.n395 585
R1184 B.n393 B.n228 585
R1185 B.n391 B.n390 585
R1186 B.n389 B.n229 585
R1187 B.n388 B.n387 585
R1188 B.n385 B.n230 585
R1189 B.n383 B.n382 585
R1190 B.n381 B.n231 585
R1191 B.n380 B.n379 585
R1192 B.n377 B.n235 585
R1193 B.n375 B.n374 585
R1194 B.n373 B.n236 585
R1195 B.n372 B.n371 585
R1196 B.n369 B.n237 585
R1197 B.n367 B.n366 585
R1198 B.n365 B.n238 585
R1199 B.n363 B.n362 585
R1200 B.n360 B.n241 585
R1201 B.n358 B.n357 585
R1202 B.n356 B.n242 585
R1203 B.n355 B.n354 585
R1204 B.n352 B.n243 585
R1205 B.n350 B.n349 585
R1206 B.n348 B.n244 585
R1207 B.n347 B.n346 585
R1208 B.n344 B.n245 585
R1209 B.n342 B.n341 585
R1210 B.n340 B.n246 585
R1211 B.n339 B.n338 585
R1212 B.n336 B.n247 585
R1213 B.n334 B.n333 585
R1214 B.n332 B.n248 585
R1215 B.n331 B.n330 585
R1216 B.n328 B.n249 585
R1217 B.n326 B.n325 585
R1218 B.n324 B.n250 585
R1219 B.n323 B.n322 585
R1220 B.n320 B.n251 585
R1221 B.n318 B.n317 585
R1222 B.n316 B.n252 585
R1223 B.n315 B.n314 585
R1224 B.n312 B.n253 585
R1225 B.n310 B.n309 585
R1226 B.n308 B.n254 585
R1227 B.n307 B.n306 585
R1228 B.n304 B.n255 585
R1229 B.n302 B.n301 585
R1230 B.n300 B.n256 585
R1231 B.n299 B.n298 585
R1232 B.n296 B.n257 585
R1233 B.n294 B.n293 585
R1234 B.n292 B.n258 585
R1235 B.n291 B.n290 585
R1236 B.n288 B.n259 585
R1237 B.n286 B.n285 585
R1238 B.n284 B.n260 585
R1239 B.n283 B.n282 585
R1240 B.n280 B.n261 585
R1241 B.n278 B.n277 585
R1242 B.n276 B.n262 585
R1243 B.n275 B.n274 585
R1244 B.n272 B.n263 585
R1245 B.n270 B.n269 585
R1246 B.n268 B.n264 585
R1247 B.n267 B.n266 585
R1248 B.n203 B.n202 585
R1249 B.n204 B.n203 585
R1250 B.n484 B.n483 585
R1251 B.n485 B.n484 585
R1252 B.n199 B.n198 585
R1253 B.n200 B.n199 585
R1254 B.n493 B.n492 585
R1255 B.n492 B.n491 585
R1256 B.n494 B.n197 585
R1257 B.n197 B.n195 585
R1258 B.n496 B.n495 585
R1259 B.n497 B.n496 585
R1260 B.n191 B.n190 585
R1261 B.n196 B.n191 585
R1262 B.n505 B.n504 585
R1263 B.n504 B.n503 585
R1264 B.n506 B.n189 585
R1265 B.n189 B.n188 585
R1266 B.n508 B.n507 585
R1267 B.n509 B.n508 585
R1268 B.n183 B.n182 585
R1269 B.n184 B.n183 585
R1270 B.n517 B.n516 585
R1271 B.n516 B.n515 585
R1272 B.n518 B.n181 585
R1273 B.n181 B.n180 585
R1274 B.n520 B.n519 585
R1275 B.n521 B.n520 585
R1276 B.n175 B.n174 585
R1277 B.n176 B.n175 585
R1278 B.n529 B.n528 585
R1279 B.n528 B.n527 585
R1280 B.n530 B.n173 585
R1281 B.n173 B.n172 585
R1282 B.n532 B.n531 585
R1283 B.n533 B.n532 585
R1284 B.n167 B.n166 585
R1285 B.n168 B.n167 585
R1286 B.n541 B.n540 585
R1287 B.n540 B.n539 585
R1288 B.n542 B.n165 585
R1289 B.n165 B.t5 585
R1290 B.n544 B.n543 585
R1291 B.n545 B.n544 585
R1292 B.n160 B.n159 585
R1293 B.n161 B.n160 585
R1294 B.n554 B.n553 585
R1295 B.n553 B.n552 585
R1296 B.n555 B.n158 585
R1297 B.n551 B.n158 585
R1298 B.n557 B.n556 585
R1299 B.n558 B.n557 585
R1300 B.n153 B.n152 585
R1301 B.n154 B.n153 585
R1302 B.n566 B.n565 585
R1303 B.n565 B.n564 585
R1304 B.n567 B.n151 585
R1305 B.n151 B.n150 585
R1306 B.n569 B.n568 585
R1307 B.n570 B.n569 585
R1308 B.n145 B.n144 585
R1309 B.n146 B.n145 585
R1310 B.n578 B.n577 585
R1311 B.n577 B.n576 585
R1312 B.n579 B.n143 585
R1313 B.n143 B.n141 585
R1314 B.n581 B.n580 585
R1315 B.n582 B.n581 585
R1316 B.n137 B.n136 585
R1317 B.n142 B.n137 585
R1318 B.n591 B.n590 585
R1319 B.n590 B.n589 585
R1320 B.n592 B.n135 585
R1321 B.n135 B.n134 585
R1322 B.n594 B.n593 585
R1323 B.n595 B.n594 585
R1324 B.n2 B.n0 585
R1325 B.n4 B.n2 585
R1326 B.n3 B.n1 585
R1327 B.n942 B.n3 585
R1328 B.n940 B.n939 585
R1329 B.n941 B.n940 585
R1330 B.n938 B.n9 585
R1331 B.n9 B.n8 585
R1332 B.n937 B.n936 585
R1333 B.n936 B.n935 585
R1334 B.n11 B.n10 585
R1335 B.n934 B.n11 585
R1336 B.n932 B.n931 585
R1337 B.n933 B.n932 585
R1338 B.n930 B.n16 585
R1339 B.n16 B.n15 585
R1340 B.n929 B.n928 585
R1341 B.n928 B.n927 585
R1342 B.n18 B.n17 585
R1343 B.n926 B.n18 585
R1344 B.n924 B.n923 585
R1345 B.n925 B.n924 585
R1346 B.n922 B.n23 585
R1347 B.n23 B.n22 585
R1348 B.n921 B.n920 585
R1349 B.n920 B.n919 585
R1350 B.n25 B.n24 585
R1351 B.n918 B.n25 585
R1352 B.n916 B.n915 585
R1353 B.n917 B.n916 585
R1354 B.n914 B.n29 585
R1355 B.n32 B.n29 585
R1356 B.n913 B.n912 585
R1357 B.n912 B.n911 585
R1358 B.n31 B.n30 585
R1359 B.n910 B.n31 585
R1360 B.n908 B.n907 585
R1361 B.n909 B.n908 585
R1362 B.n906 B.n36 585
R1363 B.n36 B.t3 585
R1364 B.n905 B.n904 585
R1365 B.n904 B.n903 585
R1366 B.n38 B.n37 585
R1367 B.n902 B.n38 585
R1368 B.n900 B.n899 585
R1369 B.n901 B.n900 585
R1370 B.n898 B.n43 585
R1371 B.n43 B.n42 585
R1372 B.n897 B.n896 585
R1373 B.n896 B.n895 585
R1374 B.n45 B.n44 585
R1375 B.n894 B.n45 585
R1376 B.n892 B.n891 585
R1377 B.n893 B.n892 585
R1378 B.n890 B.n50 585
R1379 B.n50 B.n49 585
R1380 B.n889 B.n888 585
R1381 B.n888 B.n887 585
R1382 B.n52 B.n51 585
R1383 B.n886 B.n52 585
R1384 B.n884 B.n883 585
R1385 B.n885 B.n884 585
R1386 B.n882 B.n57 585
R1387 B.n57 B.n56 585
R1388 B.n881 B.n880 585
R1389 B.n880 B.n879 585
R1390 B.n59 B.n58 585
R1391 B.n878 B.n59 585
R1392 B.n876 B.n875 585
R1393 B.n877 B.n876 585
R1394 B.n874 B.n64 585
R1395 B.n64 B.n63 585
R1396 B.n873 B.n872 585
R1397 B.n872 B.n871 585
R1398 B.n66 B.n65 585
R1399 B.n870 B.n66 585
R1400 B.n868 B.n867 585
R1401 B.n869 B.n868 585
R1402 B.n945 B.n944 585
R1403 B.n944 B.n943 585
R1404 B.n239 B.t10 468.205
R1405 B.n232 B.t18 468.205
R1406 B.n96 B.t21 468.205
R1407 B.n104 B.t14 468.205
R1408 B.n484 B.n205 458.866
R1409 B.n868 B.n71 458.866
R1410 B.n486 B.n203 458.866
R1411 B.n648 B.n69 458.866
R1412 B.n239 B.t13 364.349
R1413 B.n232 B.t20 364.349
R1414 B.n96 B.t22 364.349
R1415 B.n104 B.t16 364.349
R1416 B.n240 B.t12 331.572
R1417 B.n105 B.t17 331.572
R1418 B.n233 B.t19 331.572
R1419 B.n97 B.t23 331.572
R1420 B.n647 B.n70 256.663
R1421 B.n653 B.n70 256.663
R1422 B.n655 B.n70 256.663
R1423 B.n661 B.n70 256.663
R1424 B.n663 B.n70 256.663
R1425 B.n669 B.n70 256.663
R1426 B.n671 B.n70 256.663
R1427 B.n677 B.n70 256.663
R1428 B.n679 B.n70 256.663
R1429 B.n685 B.n70 256.663
R1430 B.n687 B.n70 256.663
R1431 B.n693 B.n70 256.663
R1432 B.n695 B.n70 256.663
R1433 B.n701 B.n70 256.663
R1434 B.n703 B.n70 256.663
R1435 B.n709 B.n70 256.663
R1436 B.n711 B.n70 256.663
R1437 B.n717 B.n70 256.663
R1438 B.n719 B.n70 256.663
R1439 B.n725 B.n70 256.663
R1440 B.n727 B.n70 256.663
R1441 B.n733 B.n70 256.663
R1442 B.n735 B.n70 256.663
R1443 B.n741 B.n70 256.663
R1444 B.n107 B.n70 256.663
R1445 B.n747 B.n70 256.663
R1446 B.n753 B.n70 256.663
R1447 B.n755 B.n70 256.663
R1448 B.n761 B.n70 256.663
R1449 B.n99 B.n70 256.663
R1450 B.n767 B.n70 256.663
R1451 B.n773 B.n70 256.663
R1452 B.n775 B.n70 256.663
R1453 B.n781 B.n70 256.663
R1454 B.n783 B.n70 256.663
R1455 B.n789 B.n70 256.663
R1456 B.n791 B.n70 256.663
R1457 B.n797 B.n70 256.663
R1458 B.n799 B.n70 256.663
R1459 B.n805 B.n70 256.663
R1460 B.n807 B.n70 256.663
R1461 B.n813 B.n70 256.663
R1462 B.n815 B.n70 256.663
R1463 B.n821 B.n70 256.663
R1464 B.n823 B.n70 256.663
R1465 B.n829 B.n70 256.663
R1466 B.n831 B.n70 256.663
R1467 B.n837 B.n70 256.663
R1468 B.n839 B.n70 256.663
R1469 B.n845 B.n70 256.663
R1470 B.n847 B.n70 256.663
R1471 B.n853 B.n70 256.663
R1472 B.n855 B.n70 256.663
R1473 B.n861 B.n70 256.663
R1474 B.n863 B.n70 256.663
R1475 B.n479 B.n204 256.663
R1476 B.n207 B.n204 256.663
R1477 B.n472 B.n204 256.663
R1478 B.n466 B.n204 256.663
R1479 B.n464 B.n204 256.663
R1480 B.n458 B.n204 256.663
R1481 B.n456 B.n204 256.663
R1482 B.n450 B.n204 256.663
R1483 B.n448 B.n204 256.663
R1484 B.n442 B.n204 256.663
R1485 B.n440 B.n204 256.663
R1486 B.n434 B.n204 256.663
R1487 B.n432 B.n204 256.663
R1488 B.n426 B.n204 256.663
R1489 B.n424 B.n204 256.663
R1490 B.n418 B.n204 256.663
R1491 B.n416 B.n204 256.663
R1492 B.n410 B.n204 256.663
R1493 B.n408 B.n204 256.663
R1494 B.n402 B.n204 256.663
R1495 B.n400 B.n204 256.663
R1496 B.n394 B.n204 256.663
R1497 B.n392 B.n204 256.663
R1498 B.n386 B.n204 256.663
R1499 B.n384 B.n204 256.663
R1500 B.n378 B.n204 256.663
R1501 B.n376 B.n204 256.663
R1502 B.n370 B.n204 256.663
R1503 B.n368 B.n204 256.663
R1504 B.n361 B.n204 256.663
R1505 B.n359 B.n204 256.663
R1506 B.n353 B.n204 256.663
R1507 B.n351 B.n204 256.663
R1508 B.n345 B.n204 256.663
R1509 B.n343 B.n204 256.663
R1510 B.n337 B.n204 256.663
R1511 B.n335 B.n204 256.663
R1512 B.n329 B.n204 256.663
R1513 B.n327 B.n204 256.663
R1514 B.n321 B.n204 256.663
R1515 B.n319 B.n204 256.663
R1516 B.n313 B.n204 256.663
R1517 B.n311 B.n204 256.663
R1518 B.n305 B.n204 256.663
R1519 B.n303 B.n204 256.663
R1520 B.n297 B.n204 256.663
R1521 B.n295 B.n204 256.663
R1522 B.n289 B.n204 256.663
R1523 B.n287 B.n204 256.663
R1524 B.n281 B.n204 256.663
R1525 B.n279 B.n204 256.663
R1526 B.n273 B.n204 256.663
R1527 B.n271 B.n204 256.663
R1528 B.n265 B.n204 256.663
R1529 B.n484 B.n199 163.367
R1530 B.n492 B.n199 163.367
R1531 B.n492 B.n197 163.367
R1532 B.n496 B.n197 163.367
R1533 B.n496 B.n191 163.367
R1534 B.n504 B.n191 163.367
R1535 B.n504 B.n189 163.367
R1536 B.n508 B.n189 163.367
R1537 B.n508 B.n183 163.367
R1538 B.n516 B.n183 163.367
R1539 B.n516 B.n181 163.367
R1540 B.n520 B.n181 163.367
R1541 B.n520 B.n175 163.367
R1542 B.n528 B.n175 163.367
R1543 B.n528 B.n173 163.367
R1544 B.n532 B.n173 163.367
R1545 B.n532 B.n167 163.367
R1546 B.n540 B.n167 163.367
R1547 B.n540 B.n165 163.367
R1548 B.n544 B.n165 163.367
R1549 B.n544 B.n160 163.367
R1550 B.n553 B.n160 163.367
R1551 B.n553 B.n158 163.367
R1552 B.n557 B.n158 163.367
R1553 B.n557 B.n153 163.367
R1554 B.n565 B.n153 163.367
R1555 B.n565 B.n151 163.367
R1556 B.n569 B.n151 163.367
R1557 B.n569 B.n145 163.367
R1558 B.n577 B.n145 163.367
R1559 B.n577 B.n143 163.367
R1560 B.n581 B.n143 163.367
R1561 B.n581 B.n137 163.367
R1562 B.n590 B.n137 163.367
R1563 B.n590 B.n135 163.367
R1564 B.n594 B.n135 163.367
R1565 B.n594 B.n2 163.367
R1566 B.n944 B.n2 163.367
R1567 B.n944 B.n3 163.367
R1568 B.n940 B.n3 163.367
R1569 B.n940 B.n9 163.367
R1570 B.n936 B.n9 163.367
R1571 B.n936 B.n11 163.367
R1572 B.n932 B.n11 163.367
R1573 B.n932 B.n16 163.367
R1574 B.n928 B.n16 163.367
R1575 B.n928 B.n18 163.367
R1576 B.n924 B.n18 163.367
R1577 B.n924 B.n23 163.367
R1578 B.n920 B.n23 163.367
R1579 B.n920 B.n25 163.367
R1580 B.n916 B.n25 163.367
R1581 B.n916 B.n29 163.367
R1582 B.n912 B.n29 163.367
R1583 B.n912 B.n31 163.367
R1584 B.n908 B.n31 163.367
R1585 B.n908 B.n36 163.367
R1586 B.n904 B.n36 163.367
R1587 B.n904 B.n38 163.367
R1588 B.n900 B.n38 163.367
R1589 B.n900 B.n43 163.367
R1590 B.n896 B.n43 163.367
R1591 B.n896 B.n45 163.367
R1592 B.n892 B.n45 163.367
R1593 B.n892 B.n50 163.367
R1594 B.n888 B.n50 163.367
R1595 B.n888 B.n52 163.367
R1596 B.n884 B.n52 163.367
R1597 B.n884 B.n57 163.367
R1598 B.n880 B.n57 163.367
R1599 B.n880 B.n59 163.367
R1600 B.n876 B.n59 163.367
R1601 B.n876 B.n64 163.367
R1602 B.n872 B.n64 163.367
R1603 B.n872 B.n66 163.367
R1604 B.n868 B.n66 163.367
R1605 B.n480 B.n478 163.367
R1606 B.n478 B.n477 163.367
R1607 B.n474 B.n473 163.367
R1608 B.n471 B.n209 163.367
R1609 B.n467 B.n465 163.367
R1610 B.n463 B.n211 163.367
R1611 B.n459 B.n457 163.367
R1612 B.n455 B.n213 163.367
R1613 B.n451 B.n449 163.367
R1614 B.n447 B.n215 163.367
R1615 B.n443 B.n441 163.367
R1616 B.n439 B.n217 163.367
R1617 B.n435 B.n433 163.367
R1618 B.n431 B.n219 163.367
R1619 B.n427 B.n425 163.367
R1620 B.n423 B.n221 163.367
R1621 B.n419 B.n417 163.367
R1622 B.n415 B.n223 163.367
R1623 B.n411 B.n409 163.367
R1624 B.n407 B.n225 163.367
R1625 B.n403 B.n401 163.367
R1626 B.n399 B.n227 163.367
R1627 B.n395 B.n393 163.367
R1628 B.n391 B.n229 163.367
R1629 B.n387 B.n385 163.367
R1630 B.n383 B.n231 163.367
R1631 B.n379 B.n377 163.367
R1632 B.n375 B.n236 163.367
R1633 B.n371 B.n369 163.367
R1634 B.n367 B.n238 163.367
R1635 B.n362 B.n360 163.367
R1636 B.n358 B.n242 163.367
R1637 B.n354 B.n352 163.367
R1638 B.n350 B.n244 163.367
R1639 B.n346 B.n344 163.367
R1640 B.n342 B.n246 163.367
R1641 B.n338 B.n336 163.367
R1642 B.n334 B.n248 163.367
R1643 B.n330 B.n328 163.367
R1644 B.n326 B.n250 163.367
R1645 B.n322 B.n320 163.367
R1646 B.n318 B.n252 163.367
R1647 B.n314 B.n312 163.367
R1648 B.n310 B.n254 163.367
R1649 B.n306 B.n304 163.367
R1650 B.n302 B.n256 163.367
R1651 B.n298 B.n296 163.367
R1652 B.n294 B.n258 163.367
R1653 B.n290 B.n288 163.367
R1654 B.n286 B.n260 163.367
R1655 B.n282 B.n280 163.367
R1656 B.n278 B.n262 163.367
R1657 B.n274 B.n272 163.367
R1658 B.n270 B.n264 163.367
R1659 B.n266 B.n203 163.367
R1660 B.n486 B.n201 163.367
R1661 B.n490 B.n201 163.367
R1662 B.n490 B.n194 163.367
R1663 B.n498 B.n194 163.367
R1664 B.n498 B.n192 163.367
R1665 B.n502 B.n192 163.367
R1666 B.n502 B.n187 163.367
R1667 B.n510 B.n187 163.367
R1668 B.n510 B.n185 163.367
R1669 B.n514 B.n185 163.367
R1670 B.n514 B.n179 163.367
R1671 B.n522 B.n179 163.367
R1672 B.n522 B.n177 163.367
R1673 B.n526 B.n177 163.367
R1674 B.n526 B.n171 163.367
R1675 B.n534 B.n171 163.367
R1676 B.n534 B.n169 163.367
R1677 B.n538 B.n169 163.367
R1678 B.n538 B.n164 163.367
R1679 B.n546 B.n164 163.367
R1680 B.n546 B.n162 163.367
R1681 B.n550 B.n162 163.367
R1682 B.n550 B.n157 163.367
R1683 B.n559 B.n157 163.367
R1684 B.n559 B.n155 163.367
R1685 B.n563 B.n155 163.367
R1686 B.n563 B.n149 163.367
R1687 B.n571 B.n149 163.367
R1688 B.n571 B.n147 163.367
R1689 B.n575 B.n147 163.367
R1690 B.n575 B.n140 163.367
R1691 B.n583 B.n140 163.367
R1692 B.n583 B.n138 163.367
R1693 B.n588 B.n138 163.367
R1694 B.n588 B.n133 163.367
R1695 B.n596 B.n133 163.367
R1696 B.n597 B.n596 163.367
R1697 B.n597 B.n5 163.367
R1698 B.n6 B.n5 163.367
R1699 B.n7 B.n6 163.367
R1700 B.n602 B.n7 163.367
R1701 B.n602 B.n12 163.367
R1702 B.n13 B.n12 163.367
R1703 B.n14 B.n13 163.367
R1704 B.n607 B.n14 163.367
R1705 B.n607 B.n19 163.367
R1706 B.n20 B.n19 163.367
R1707 B.n21 B.n20 163.367
R1708 B.n612 B.n21 163.367
R1709 B.n612 B.n26 163.367
R1710 B.n27 B.n26 163.367
R1711 B.n28 B.n27 163.367
R1712 B.n617 B.n28 163.367
R1713 B.n617 B.n33 163.367
R1714 B.n34 B.n33 163.367
R1715 B.n35 B.n34 163.367
R1716 B.n622 B.n35 163.367
R1717 B.n622 B.n39 163.367
R1718 B.n40 B.n39 163.367
R1719 B.n41 B.n40 163.367
R1720 B.n627 B.n41 163.367
R1721 B.n627 B.n46 163.367
R1722 B.n47 B.n46 163.367
R1723 B.n48 B.n47 163.367
R1724 B.n632 B.n48 163.367
R1725 B.n632 B.n53 163.367
R1726 B.n54 B.n53 163.367
R1727 B.n55 B.n54 163.367
R1728 B.n637 B.n55 163.367
R1729 B.n637 B.n60 163.367
R1730 B.n61 B.n60 163.367
R1731 B.n62 B.n61 163.367
R1732 B.n642 B.n62 163.367
R1733 B.n642 B.n67 163.367
R1734 B.n68 B.n67 163.367
R1735 B.n69 B.n68 163.367
R1736 B.n864 B.n862 163.367
R1737 B.n860 B.n73 163.367
R1738 B.n856 B.n854 163.367
R1739 B.n852 B.n75 163.367
R1740 B.n848 B.n846 163.367
R1741 B.n844 B.n77 163.367
R1742 B.n840 B.n838 163.367
R1743 B.n836 B.n79 163.367
R1744 B.n832 B.n830 163.367
R1745 B.n828 B.n81 163.367
R1746 B.n824 B.n822 163.367
R1747 B.n820 B.n83 163.367
R1748 B.n816 B.n814 163.367
R1749 B.n812 B.n85 163.367
R1750 B.n808 B.n806 163.367
R1751 B.n804 B.n87 163.367
R1752 B.n800 B.n798 163.367
R1753 B.n796 B.n89 163.367
R1754 B.n792 B.n790 163.367
R1755 B.n788 B.n91 163.367
R1756 B.n784 B.n782 163.367
R1757 B.n780 B.n93 163.367
R1758 B.n776 B.n774 163.367
R1759 B.n772 B.n95 163.367
R1760 B.n768 B.n766 163.367
R1761 B.n763 B.n762 163.367
R1762 B.n760 B.n101 163.367
R1763 B.n756 B.n754 163.367
R1764 B.n752 B.n103 163.367
R1765 B.n748 B.n746 163.367
R1766 B.n743 B.n742 163.367
R1767 B.n740 B.n109 163.367
R1768 B.n736 B.n734 163.367
R1769 B.n732 B.n111 163.367
R1770 B.n728 B.n726 163.367
R1771 B.n724 B.n113 163.367
R1772 B.n720 B.n718 163.367
R1773 B.n716 B.n115 163.367
R1774 B.n712 B.n710 163.367
R1775 B.n708 B.n117 163.367
R1776 B.n704 B.n702 163.367
R1777 B.n700 B.n119 163.367
R1778 B.n696 B.n694 163.367
R1779 B.n692 B.n121 163.367
R1780 B.n688 B.n686 163.367
R1781 B.n684 B.n123 163.367
R1782 B.n680 B.n678 163.367
R1783 B.n676 B.n125 163.367
R1784 B.n672 B.n670 163.367
R1785 B.n668 B.n127 163.367
R1786 B.n664 B.n662 163.367
R1787 B.n660 B.n129 163.367
R1788 B.n656 B.n654 163.367
R1789 B.n652 B.n131 163.367
R1790 B.n479 B.n205 71.676
R1791 B.n477 B.n207 71.676
R1792 B.n473 B.n472 71.676
R1793 B.n466 B.n209 71.676
R1794 B.n465 B.n464 71.676
R1795 B.n458 B.n211 71.676
R1796 B.n457 B.n456 71.676
R1797 B.n450 B.n213 71.676
R1798 B.n449 B.n448 71.676
R1799 B.n442 B.n215 71.676
R1800 B.n441 B.n440 71.676
R1801 B.n434 B.n217 71.676
R1802 B.n433 B.n432 71.676
R1803 B.n426 B.n219 71.676
R1804 B.n425 B.n424 71.676
R1805 B.n418 B.n221 71.676
R1806 B.n417 B.n416 71.676
R1807 B.n410 B.n223 71.676
R1808 B.n409 B.n408 71.676
R1809 B.n402 B.n225 71.676
R1810 B.n401 B.n400 71.676
R1811 B.n394 B.n227 71.676
R1812 B.n393 B.n392 71.676
R1813 B.n386 B.n229 71.676
R1814 B.n385 B.n384 71.676
R1815 B.n378 B.n231 71.676
R1816 B.n377 B.n376 71.676
R1817 B.n370 B.n236 71.676
R1818 B.n369 B.n368 71.676
R1819 B.n361 B.n238 71.676
R1820 B.n360 B.n359 71.676
R1821 B.n353 B.n242 71.676
R1822 B.n352 B.n351 71.676
R1823 B.n345 B.n244 71.676
R1824 B.n344 B.n343 71.676
R1825 B.n337 B.n246 71.676
R1826 B.n336 B.n335 71.676
R1827 B.n329 B.n248 71.676
R1828 B.n328 B.n327 71.676
R1829 B.n321 B.n250 71.676
R1830 B.n320 B.n319 71.676
R1831 B.n313 B.n252 71.676
R1832 B.n312 B.n311 71.676
R1833 B.n305 B.n254 71.676
R1834 B.n304 B.n303 71.676
R1835 B.n297 B.n256 71.676
R1836 B.n296 B.n295 71.676
R1837 B.n289 B.n258 71.676
R1838 B.n288 B.n287 71.676
R1839 B.n281 B.n260 71.676
R1840 B.n280 B.n279 71.676
R1841 B.n273 B.n262 71.676
R1842 B.n272 B.n271 71.676
R1843 B.n265 B.n264 71.676
R1844 B.n863 B.n71 71.676
R1845 B.n862 B.n861 71.676
R1846 B.n855 B.n73 71.676
R1847 B.n854 B.n853 71.676
R1848 B.n847 B.n75 71.676
R1849 B.n846 B.n845 71.676
R1850 B.n839 B.n77 71.676
R1851 B.n838 B.n837 71.676
R1852 B.n831 B.n79 71.676
R1853 B.n830 B.n829 71.676
R1854 B.n823 B.n81 71.676
R1855 B.n822 B.n821 71.676
R1856 B.n815 B.n83 71.676
R1857 B.n814 B.n813 71.676
R1858 B.n807 B.n85 71.676
R1859 B.n806 B.n805 71.676
R1860 B.n799 B.n87 71.676
R1861 B.n798 B.n797 71.676
R1862 B.n791 B.n89 71.676
R1863 B.n790 B.n789 71.676
R1864 B.n783 B.n91 71.676
R1865 B.n782 B.n781 71.676
R1866 B.n775 B.n93 71.676
R1867 B.n774 B.n773 71.676
R1868 B.n767 B.n95 71.676
R1869 B.n766 B.n99 71.676
R1870 B.n762 B.n761 71.676
R1871 B.n755 B.n101 71.676
R1872 B.n754 B.n753 71.676
R1873 B.n747 B.n103 71.676
R1874 B.n746 B.n107 71.676
R1875 B.n742 B.n741 71.676
R1876 B.n735 B.n109 71.676
R1877 B.n734 B.n733 71.676
R1878 B.n727 B.n111 71.676
R1879 B.n726 B.n725 71.676
R1880 B.n719 B.n113 71.676
R1881 B.n718 B.n717 71.676
R1882 B.n711 B.n115 71.676
R1883 B.n710 B.n709 71.676
R1884 B.n703 B.n117 71.676
R1885 B.n702 B.n701 71.676
R1886 B.n695 B.n119 71.676
R1887 B.n694 B.n693 71.676
R1888 B.n687 B.n121 71.676
R1889 B.n686 B.n685 71.676
R1890 B.n679 B.n123 71.676
R1891 B.n678 B.n677 71.676
R1892 B.n671 B.n125 71.676
R1893 B.n670 B.n669 71.676
R1894 B.n663 B.n127 71.676
R1895 B.n662 B.n661 71.676
R1896 B.n655 B.n129 71.676
R1897 B.n654 B.n653 71.676
R1898 B.n647 B.n131 71.676
R1899 B.n648 B.n647 71.676
R1900 B.n653 B.n652 71.676
R1901 B.n656 B.n655 71.676
R1902 B.n661 B.n660 71.676
R1903 B.n664 B.n663 71.676
R1904 B.n669 B.n668 71.676
R1905 B.n672 B.n671 71.676
R1906 B.n677 B.n676 71.676
R1907 B.n680 B.n679 71.676
R1908 B.n685 B.n684 71.676
R1909 B.n688 B.n687 71.676
R1910 B.n693 B.n692 71.676
R1911 B.n696 B.n695 71.676
R1912 B.n701 B.n700 71.676
R1913 B.n704 B.n703 71.676
R1914 B.n709 B.n708 71.676
R1915 B.n712 B.n711 71.676
R1916 B.n717 B.n716 71.676
R1917 B.n720 B.n719 71.676
R1918 B.n725 B.n724 71.676
R1919 B.n728 B.n727 71.676
R1920 B.n733 B.n732 71.676
R1921 B.n736 B.n735 71.676
R1922 B.n741 B.n740 71.676
R1923 B.n743 B.n107 71.676
R1924 B.n748 B.n747 71.676
R1925 B.n753 B.n752 71.676
R1926 B.n756 B.n755 71.676
R1927 B.n761 B.n760 71.676
R1928 B.n763 B.n99 71.676
R1929 B.n768 B.n767 71.676
R1930 B.n773 B.n772 71.676
R1931 B.n776 B.n775 71.676
R1932 B.n781 B.n780 71.676
R1933 B.n784 B.n783 71.676
R1934 B.n789 B.n788 71.676
R1935 B.n792 B.n791 71.676
R1936 B.n797 B.n796 71.676
R1937 B.n800 B.n799 71.676
R1938 B.n805 B.n804 71.676
R1939 B.n808 B.n807 71.676
R1940 B.n813 B.n812 71.676
R1941 B.n816 B.n815 71.676
R1942 B.n821 B.n820 71.676
R1943 B.n824 B.n823 71.676
R1944 B.n829 B.n828 71.676
R1945 B.n832 B.n831 71.676
R1946 B.n837 B.n836 71.676
R1947 B.n840 B.n839 71.676
R1948 B.n845 B.n844 71.676
R1949 B.n848 B.n847 71.676
R1950 B.n853 B.n852 71.676
R1951 B.n856 B.n855 71.676
R1952 B.n861 B.n860 71.676
R1953 B.n864 B.n863 71.676
R1954 B.n480 B.n479 71.676
R1955 B.n474 B.n207 71.676
R1956 B.n472 B.n471 71.676
R1957 B.n467 B.n466 71.676
R1958 B.n464 B.n463 71.676
R1959 B.n459 B.n458 71.676
R1960 B.n456 B.n455 71.676
R1961 B.n451 B.n450 71.676
R1962 B.n448 B.n447 71.676
R1963 B.n443 B.n442 71.676
R1964 B.n440 B.n439 71.676
R1965 B.n435 B.n434 71.676
R1966 B.n432 B.n431 71.676
R1967 B.n427 B.n426 71.676
R1968 B.n424 B.n423 71.676
R1969 B.n419 B.n418 71.676
R1970 B.n416 B.n415 71.676
R1971 B.n411 B.n410 71.676
R1972 B.n408 B.n407 71.676
R1973 B.n403 B.n402 71.676
R1974 B.n400 B.n399 71.676
R1975 B.n395 B.n394 71.676
R1976 B.n392 B.n391 71.676
R1977 B.n387 B.n386 71.676
R1978 B.n384 B.n383 71.676
R1979 B.n379 B.n378 71.676
R1980 B.n376 B.n375 71.676
R1981 B.n371 B.n370 71.676
R1982 B.n368 B.n367 71.676
R1983 B.n362 B.n361 71.676
R1984 B.n359 B.n358 71.676
R1985 B.n354 B.n353 71.676
R1986 B.n351 B.n350 71.676
R1987 B.n346 B.n345 71.676
R1988 B.n343 B.n342 71.676
R1989 B.n338 B.n337 71.676
R1990 B.n335 B.n334 71.676
R1991 B.n330 B.n329 71.676
R1992 B.n327 B.n326 71.676
R1993 B.n322 B.n321 71.676
R1994 B.n319 B.n318 71.676
R1995 B.n314 B.n313 71.676
R1996 B.n311 B.n310 71.676
R1997 B.n306 B.n305 71.676
R1998 B.n303 B.n302 71.676
R1999 B.n298 B.n297 71.676
R2000 B.n295 B.n294 71.676
R2001 B.n290 B.n289 71.676
R2002 B.n287 B.n286 71.676
R2003 B.n282 B.n281 71.676
R2004 B.n279 B.n278 71.676
R2005 B.n274 B.n273 71.676
R2006 B.n271 B.n270 71.676
R2007 B.n266 B.n265 71.676
R2008 B.n485 B.n204 65.0117
R2009 B.n869 B.n70 65.0117
R2010 B.n364 B.n240 59.5399
R2011 B.n234 B.n233 59.5399
R2012 B.n98 B.n97 59.5399
R2013 B.n106 B.n105 59.5399
R2014 B.n485 B.n200 37.1497
R2015 B.n491 B.n200 37.1497
R2016 B.n491 B.n195 37.1497
R2017 B.n497 B.n195 37.1497
R2018 B.n497 B.n196 37.1497
R2019 B.n503 B.n188 37.1497
R2020 B.n509 B.n188 37.1497
R2021 B.n509 B.n184 37.1497
R2022 B.n515 B.n184 37.1497
R2023 B.n515 B.n180 37.1497
R2024 B.n521 B.n180 37.1497
R2025 B.n521 B.n176 37.1497
R2026 B.n527 B.n176 37.1497
R2027 B.n533 B.n172 37.1497
R2028 B.n533 B.n168 37.1497
R2029 B.n539 B.n168 37.1497
R2030 B.n539 B.t5 37.1497
R2031 B.n545 B.t5 37.1497
R2032 B.n545 B.n161 37.1497
R2033 B.n552 B.n161 37.1497
R2034 B.n552 B.n551 37.1497
R2035 B.n558 B.n154 37.1497
R2036 B.n564 B.n154 37.1497
R2037 B.n564 B.n150 37.1497
R2038 B.n570 B.n150 37.1497
R2039 B.n576 B.n146 37.1497
R2040 B.n576 B.n141 37.1497
R2041 B.n582 B.n141 37.1497
R2042 B.n582 B.n142 37.1497
R2043 B.n589 B.n134 37.1497
R2044 B.n595 B.n134 37.1497
R2045 B.n595 B.n4 37.1497
R2046 B.n943 B.n4 37.1497
R2047 B.n943 B.n942 37.1497
R2048 B.n942 B.n941 37.1497
R2049 B.n941 B.n8 37.1497
R2050 B.n935 B.n8 37.1497
R2051 B.n934 B.n933 37.1497
R2052 B.n933 B.n15 37.1497
R2053 B.n927 B.n15 37.1497
R2054 B.n927 B.n926 37.1497
R2055 B.n925 B.n22 37.1497
R2056 B.n919 B.n22 37.1497
R2057 B.n919 B.n918 37.1497
R2058 B.n918 B.n917 37.1497
R2059 B.n911 B.n32 37.1497
R2060 B.n911 B.n910 37.1497
R2061 B.n910 B.n909 37.1497
R2062 B.n909 B.t3 37.1497
R2063 B.n903 B.t3 37.1497
R2064 B.n903 B.n902 37.1497
R2065 B.n902 B.n901 37.1497
R2066 B.n901 B.n42 37.1497
R2067 B.n895 B.n894 37.1497
R2068 B.n894 B.n893 37.1497
R2069 B.n893 B.n49 37.1497
R2070 B.n887 B.n49 37.1497
R2071 B.n887 B.n886 37.1497
R2072 B.n886 B.n885 37.1497
R2073 B.n885 B.n56 37.1497
R2074 B.n879 B.n56 37.1497
R2075 B.n878 B.n877 37.1497
R2076 B.n877 B.n63 37.1497
R2077 B.n871 B.n63 37.1497
R2078 B.n871 B.n870 37.1497
R2079 B.n870 B.n869 37.1497
R2080 B.t9 B.n172 36.0571
R2081 B.n551 B.t2 36.0571
R2082 B.n32 B.t0 36.0571
R2083 B.t6 B.n42 36.0571
R2084 B.n570 B.t8 34.9645
R2085 B.t1 B.n925 34.9645
R2086 B.n142 B.t4 33.8719
R2087 B.t7 B.n934 33.8719
R2088 B.n240 B.n239 32.7763
R2089 B.n233 B.n232 32.7763
R2090 B.n97 B.n96 32.7763
R2091 B.n105 B.n104 32.7763
R2092 B.n196 B.t11 31.6866
R2093 B.t15 B.n878 31.6866
R2094 B.n867 B.n866 29.8151
R2095 B.n649 B.n646 29.8151
R2096 B.n487 B.n202 29.8151
R2097 B.n483 B.n482 29.8151
R2098 B B.n945 18.0485
R2099 B.n866 B.n865 10.6151
R2100 B.n865 B.n72 10.6151
R2101 B.n859 B.n72 10.6151
R2102 B.n859 B.n858 10.6151
R2103 B.n858 B.n857 10.6151
R2104 B.n857 B.n74 10.6151
R2105 B.n851 B.n74 10.6151
R2106 B.n851 B.n850 10.6151
R2107 B.n850 B.n849 10.6151
R2108 B.n849 B.n76 10.6151
R2109 B.n843 B.n76 10.6151
R2110 B.n843 B.n842 10.6151
R2111 B.n842 B.n841 10.6151
R2112 B.n841 B.n78 10.6151
R2113 B.n835 B.n78 10.6151
R2114 B.n835 B.n834 10.6151
R2115 B.n834 B.n833 10.6151
R2116 B.n833 B.n80 10.6151
R2117 B.n827 B.n80 10.6151
R2118 B.n827 B.n826 10.6151
R2119 B.n826 B.n825 10.6151
R2120 B.n825 B.n82 10.6151
R2121 B.n819 B.n82 10.6151
R2122 B.n819 B.n818 10.6151
R2123 B.n818 B.n817 10.6151
R2124 B.n817 B.n84 10.6151
R2125 B.n811 B.n84 10.6151
R2126 B.n811 B.n810 10.6151
R2127 B.n810 B.n809 10.6151
R2128 B.n809 B.n86 10.6151
R2129 B.n803 B.n86 10.6151
R2130 B.n803 B.n802 10.6151
R2131 B.n802 B.n801 10.6151
R2132 B.n801 B.n88 10.6151
R2133 B.n795 B.n88 10.6151
R2134 B.n795 B.n794 10.6151
R2135 B.n794 B.n793 10.6151
R2136 B.n793 B.n90 10.6151
R2137 B.n787 B.n90 10.6151
R2138 B.n787 B.n786 10.6151
R2139 B.n786 B.n785 10.6151
R2140 B.n785 B.n92 10.6151
R2141 B.n779 B.n92 10.6151
R2142 B.n779 B.n778 10.6151
R2143 B.n778 B.n777 10.6151
R2144 B.n777 B.n94 10.6151
R2145 B.n771 B.n94 10.6151
R2146 B.n771 B.n770 10.6151
R2147 B.n770 B.n769 10.6151
R2148 B.n765 B.n764 10.6151
R2149 B.n764 B.n100 10.6151
R2150 B.n759 B.n100 10.6151
R2151 B.n759 B.n758 10.6151
R2152 B.n758 B.n757 10.6151
R2153 B.n757 B.n102 10.6151
R2154 B.n751 B.n102 10.6151
R2155 B.n751 B.n750 10.6151
R2156 B.n750 B.n749 10.6151
R2157 B.n745 B.n744 10.6151
R2158 B.n744 B.n108 10.6151
R2159 B.n739 B.n108 10.6151
R2160 B.n739 B.n738 10.6151
R2161 B.n738 B.n737 10.6151
R2162 B.n737 B.n110 10.6151
R2163 B.n731 B.n110 10.6151
R2164 B.n731 B.n730 10.6151
R2165 B.n730 B.n729 10.6151
R2166 B.n729 B.n112 10.6151
R2167 B.n723 B.n112 10.6151
R2168 B.n723 B.n722 10.6151
R2169 B.n722 B.n721 10.6151
R2170 B.n721 B.n114 10.6151
R2171 B.n715 B.n114 10.6151
R2172 B.n715 B.n714 10.6151
R2173 B.n714 B.n713 10.6151
R2174 B.n713 B.n116 10.6151
R2175 B.n707 B.n116 10.6151
R2176 B.n707 B.n706 10.6151
R2177 B.n706 B.n705 10.6151
R2178 B.n705 B.n118 10.6151
R2179 B.n699 B.n118 10.6151
R2180 B.n699 B.n698 10.6151
R2181 B.n698 B.n697 10.6151
R2182 B.n697 B.n120 10.6151
R2183 B.n691 B.n120 10.6151
R2184 B.n691 B.n690 10.6151
R2185 B.n690 B.n689 10.6151
R2186 B.n689 B.n122 10.6151
R2187 B.n683 B.n122 10.6151
R2188 B.n683 B.n682 10.6151
R2189 B.n682 B.n681 10.6151
R2190 B.n681 B.n124 10.6151
R2191 B.n675 B.n124 10.6151
R2192 B.n675 B.n674 10.6151
R2193 B.n674 B.n673 10.6151
R2194 B.n673 B.n126 10.6151
R2195 B.n667 B.n126 10.6151
R2196 B.n667 B.n666 10.6151
R2197 B.n666 B.n665 10.6151
R2198 B.n665 B.n128 10.6151
R2199 B.n659 B.n128 10.6151
R2200 B.n659 B.n658 10.6151
R2201 B.n658 B.n657 10.6151
R2202 B.n657 B.n130 10.6151
R2203 B.n651 B.n130 10.6151
R2204 B.n651 B.n650 10.6151
R2205 B.n650 B.n649 10.6151
R2206 B.n488 B.n487 10.6151
R2207 B.n489 B.n488 10.6151
R2208 B.n489 B.n193 10.6151
R2209 B.n499 B.n193 10.6151
R2210 B.n500 B.n499 10.6151
R2211 B.n501 B.n500 10.6151
R2212 B.n501 B.n186 10.6151
R2213 B.n511 B.n186 10.6151
R2214 B.n512 B.n511 10.6151
R2215 B.n513 B.n512 10.6151
R2216 B.n513 B.n178 10.6151
R2217 B.n523 B.n178 10.6151
R2218 B.n524 B.n523 10.6151
R2219 B.n525 B.n524 10.6151
R2220 B.n525 B.n170 10.6151
R2221 B.n535 B.n170 10.6151
R2222 B.n536 B.n535 10.6151
R2223 B.n537 B.n536 10.6151
R2224 B.n537 B.n163 10.6151
R2225 B.n547 B.n163 10.6151
R2226 B.n548 B.n547 10.6151
R2227 B.n549 B.n548 10.6151
R2228 B.n549 B.n156 10.6151
R2229 B.n560 B.n156 10.6151
R2230 B.n561 B.n560 10.6151
R2231 B.n562 B.n561 10.6151
R2232 B.n562 B.n148 10.6151
R2233 B.n572 B.n148 10.6151
R2234 B.n573 B.n572 10.6151
R2235 B.n574 B.n573 10.6151
R2236 B.n574 B.n139 10.6151
R2237 B.n584 B.n139 10.6151
R2238 B.n585 B.n584 10.6151
R2239 B.n587 B.n585 10.6151
R2240 B.n587 B.n586 10.6151
R2241 B.n586 B.n132 10.6151
R2242 B.n598 B.n132 10.6151
R2243 B.n599 B.n598 10.6151
R2244 B.n600 B.n599 10.6151
R2245 B.n601 B.n600 10.6151
R2246 B.n603 B.n601 10.6151
R2247 B.n604 B.n603 10.6151
R2248 B.n605 B.n604 10.6151
R2249 B.n606 B.n605 10.6151
R2250 B.n608 B.n606 10.6151
R2251 B.n609 B.n608 10.6151
R2252 B.n610 B.n609 10.6151
R2253 B.n611 B.n610 10.6151
R2254 B.n613 B.n611 10.6151
R2255 B.n614 B.n613 10.6151
R2256 B.n615 B.n614 10.6151
R2257 B.n616 B.n615 10.6151
R2258 B.n618 B.n616 10.6151
R2259 B.n619 B.n618 10.6151
R2260 B.n620 B.n619 10.6151
R2261 B.n621 B.n620 10.6151
R2262 B.n623 B.n621 10.6151
R2263 B.n624 B.n623 10.6151
R2264 B.n625 B.n624 10.6151
R2265 B.n626 B.n625 10.6151
R2266 B.n628 B.n626 10.6151
R2267 B.n629 B.n628 10.6151
R2268 B.n630 B.n629 10.6151
R2269 B.n631 B.n630 10.6151
R2270 B.n633 B.n631 10.6151
R2271 B.n634 B.n633 10.6151
R2272 B.n635 B.n634 10.6151
R2273 B.n636 B.n635 10.6151
R2274 B.n638 B.n636 10.6151
R2275 B.n639 B.n638 10.6151
R2276 B.n640 B.n639 10.6151
R2277 B.n641 B.n640 10.6151
R2278 B.n643 B.n641 10.6151
R2279 B.n644 B.n643 10.6151
R2280 B.n645 B.n644 10.6151
R2281 B.n646 B.n645 10.6151
R2282 B.n482 B.n481 10.6151
R2283 B.n481 B.n206 10.6151
R2284 B.n476 B.n206 10.6151
R2285 B.n476 B.n475 10.6151
R2286 B.n475 B.n208 10.6151
R2287 B.n470 B.n208 10.6151
R2288 B.n470 B.n469 10.6151
R2289 B.n469 B.n468 10.6151
R2290 B.n468 B.n210 10.6151
R2291 B.n462 B.n210 10.6151
R2292 B.n462 B.n461 10.6151
R2293 B.n461 B.n460 10.6151
R2294 B.n460 B.n212 10.6151
R2295 B.n454 B.n212 10.6151
R2296 B.n454 B.n453 10.6151
R2297 B.n453 B.n452 10.6151
R2298 B.n452 B.n214 10.6151
R2299 B.n446 B.n214 10.6151
R2300 B.n446 B.n445 10.6151
R2301 B.n445 B.n444 10.6151
R2302 B.n444 B.n216 10.6151
R2303 B.n438 B.n216 10.6151
R2304 B.n438 B.n437 10.6151
R2305 B.n437 B.n436 10.6151
R2306 B.n436 B.n218 10.6151
R2307 B.n430 B.n218 10.6151
R2308 B.n430 B.n429 10.6151
R2309 B.n429 B.n428 10.6151
R2310 B.n428 B.n220 10.6151
R2311 B.n422 B.n220 10.6151
R2312 B.n422 B.n421 10.6151
R2313 B.n421 B.n420 10.6151
R2314 B.n420 B.n222 10.6151
R2315 B.n414 B.n222 10.6151
R2316 B.n414 B.n413 10.6151
R2317 B.n413 B.n412 10.6151
R2318 B.n412 B.n224 10.6151
R2319 B.n406 B.n224 10.6151
R2320 B.n406 B.n405 10.6151
R2321 B.n405 B.n404 10.6151
R2322 B.n404 B.n226 10.6151
R2323 B.n398 B.n226 10.6151
R2324 B.n398 B.n397 10.6151
R2325 B.n397 B.n396 10.6151
R2326 B.n396 B.n228 10.6151
R2327 B.n390 B.n228 10.6151
R2328 B.n390 B.n389 10.6151
R2329 B.n389 B.n388 10.6151
R2330 B.n388 B.n230 10.6151
R2331 B.n382 B.n381 10.6151
R2332 B.n381 B.n380 10.6151
R2333 B.n380 B.n235 10.6151
R2334 B.n374 B.n235 10.6151
R2335 B.n374 B.n373 10.6151
R2336 B.n373 B.n372 10.6151
R2337 B.n372 B.n237 10.6151
R2338 B.n366 B.n237 10.6151
R2339 B.n366 B.n365 10.6151
R2340 B.n363 B.n241 10.6151
R2341 B.n357 B.n241 10.6151
R2342 B.n357 B.n356 10.6151
R2343 B.n356 B.n355 10.6151
R2344 B.n355 B.n243 10.6151
R2345 B.n349 B.n243 10.6151
R2346 B.n349 B.n348 10.6151
R2347 B.n348 B.n347 10.6151
R2348 B.n347 B.n245 10.6151
R2349 B.n341 B.n245 10.6151
R2350 B.n341 B.n340 10.6151
R2351 B.n340 B.n339 10.6151
R2352 B.n339 B.n247 10.6151
R2353 B.n333 B.n247 10.6151
R2354 B.n333 B.n332 10.6151
R2355 B.n332 B.n331 10.6151
R2356 B.n331 B.n249 10.6151
R2357 B.n325 B.n249 10.6151
R2358 B.n325 B.n324 10.6151
R2359 B.n324 B.n323 10.6151
R2360 B.n323 B.n251 10.6151
R2361 B.n317 B.n251 10.6151
R2362 B.n317 B.n316 10.6151
R2363 B.n316 B.n315 10.6151
R2364 B.n315 B.n253 10.6151
R2365 B.n309 B.n253 10.6151
R2366 B.n309 B.n308 10.6151
R2367 B.n308 B.n307 10.6151
R2368 B.n307 B.n255 10.6151
R2369 B.n301 B.n255 10.6151
R2370 B.n301 B.n300 10.6151
R2371 B.n300 B.n299 10.6151
R2372 B.n299 B.n257 10.6151
R2373 B.n293 B.n257 10.6151
R2374 B.n293 B.n292 10.6151
R2375 B.n292 B.n291 10.6151
R2376 B.n291 B.n259 10.6151
R2377 B.n285 B.n259 10.6151
R2378 B.n285 B.n284 10.6151
R2379 B.n284 B.n283 10.6151
R2380 B.n283 B.n261 10.6151
R2381 B.n277 B.n261 10.6151
R2382 B.n277 B.n276 10.6151
R2383 B.n276 B.n275 10.6151
R2384 B.n275 B.n263 10.6151
R2385 B.n269 B.n263 10.6151
R2386 B.n269 B.n268 10.6151
R2387 B.n268 B.n267 10.6151
R2388 B.n267 B.n202 10.6151
R2389 B.n483 B.n198 10.6151
R2390 B.n493 B.n198 10.6151
R2391 B.n494 B.n493 10.6151
R2392 B.n495 B.n494 10.6151
R2393 B.n495 B.n190 10.6151
R2394 B.n505 B.n190 10.6151
R2395 B.n506 B.n505 10.6151
R2396 B.n507 B.n506 10.6151
R2397 B.n507 B.n182 10.6151
R2398 B.n517 B.n182 10.6151
R2399 B.n518 B.n517 10.6151
R2400 B.n519 B.n518 10.6151
R2401 B.n519 B.n174 10.6151
R2402 B.n529 B.n174 10.6151
R2403 B.n530 B.n529 10.6151
R2404 B.n531 B.n530 10.6151
R2405 B.n531 B.n166 10.6151
R2406 B.n541 B.n166 10.6151
R2407 B.n542 B.n541 10.6151
R2408 B.n543 B.n542 10.6151
R2409 B.n543 B.n159 10.6151
R2410 B.n554 B.n159 10.6151
R2411 B.n555 B.n554 10.6151
R2412 B.n556 B.n555 10.6151
R2413 B.n556 B.n152 10.6151
R2414 B.n566 B.n152 10.6151
R2415 B.n567 B.n566 10.6151
R2416 B.n568 B.n567 10.6151
R2417 B.n568 B.n144 10.6151
R2418 B.n578 B.n144 10.6151
R2419 B.n579 B.n578 10.6151
R2420 B.n580 B.n579 10.6151
R2421 B.n580 B.n136 10.6151
R2422 B.n591 B.n136 10.6151
R2423 B.n592 B.n591 10.6151
R2424 B.n593 B.n592 10.6151
R2425 B.n593 B.n0 10.6151
R2426 B.n939 B.n1 10.6151
R2427 B.n939 B.n938 10.6151
R2428 B.n938 B.n937 10.6151
R2429 B.n937 B.n10 10.6151
R2430 B.n931 B.n10 10.6151
R2431 B.n931 B.n930 10.6151
R2432 B.n930 B.n929 10.6151
R2433 B.n929 B.n17 10.6151
R2434 B.n923 B.n17 10.6151
R2435 B.n923 B.n922 10.6151
R2436 B.n922 B.n921 10.6151
R2437 B.n921 B.n24 10.6151
R2438 B.n915 B.n24 10.6151
R2439 B.n915 B.n914 10.6151
R2440 B.n914 B.n913 10.6151
R2441 B.n913 B.n30 10.6151
R2442 B.n907 B.n30 10.6151
R2443 B.n907 B.n906 10.6151
R2444 B.n906 B.n905 10.6151
R2445 B.n905 B.n37 10.6151
R2446 B.n899 B.n37 10.6151
R2447 B.n899 B.n898 10.6151
R2448 B.n898 B.n897 10.6151
R2449 B.n897 B.n44 10.6151
R2450 B.n891 B.n44 10.6151
R2451 B.n891 B.n890 10.6151
R2452 B.n890 B.n889 10.6151
R2453 B.n889 B.n51 10.6151
R2454 B.n883 B.n51 10.6151
R2455 B.n883 B.n882 10.6151
R2456 B.n882 B.n881 10.6151
R2457 B.n881 B.n58 10.6151
R2458 B.n875 B.n58 10.6151
R2459 B.n875 B.n874 10.6151
R2460 B.n874 B.n873 10.6151
R2461 B.n873 B.n65 10.6151
R2462 B.n867 B.n65 10.6151
R2463 B.n769 B.n98 9.36635
R2464 B.n745 B.n106 9.36635
R2465 B.n234 B.n230 9.36635
R2466 B.n364 B.n363 9.36635
R2467 B.n503 B.t11 5.46362
R2468 B.n879 B.t15 5.46362
R2469 B.n589 B.t4 3.27837
R2470 B.n935 B.t7 3.27837
R2471 B.n945 B.n0 2.81026
R2472 B.n945 B.n1 2.81026
R2473 B.t8 B.n146 2.18575
R2474 B.n926 B.t1 2.18575
R2475 B.n765 B.n98 1.24928
R2476 B.n749 B.n106 1.24928
R2477 B.n382 B.n234 1.24928
R2478 B.n365 B.n364 1.24928
R2479 B.n527 B.t9 1.09312
R2480 B.n558 B.t2 1.09312
R2481 B.n917 B.t0 1.09312
R2482 B.n895 B.t6 1.09312
R2483 VN.n6 VN.t8 310.889
R2484 VN.n29 VN.t5 310.889
R2485 VN.n21 VN.t7 292.212
R2486 VN.n44 VN.t9 292.212
R2487 VN.n3 VN.t6 263.329
R2488 VN.n5 VN.t1 263.329
R2489 VN.n1 VN.t4 263.329
R2490 VN.n26 VN.t3 263.329
R2491 VN.n28 VN.t2 263.329
R2492 VN.n24 VN.t0 263.329
R2493 VN.n43 VN.n23 161.3
R2494 VN.n42 VN.n41 161.3
R2495 VN.n40 VN.n39 161.3
R2496 VN.n38 VN.n25 161.3
R2497 VN.n37 VN.n36 161.3
R2498 VN.n35 VN.n26 161.3
R2499 VN.n34 VN.n33 161.3
R2500 VN.n32 VN.n27 161.3
R2501 VN.n31 VN.n30 161.3
R2502 VN.n20 VN.n0 161.3
R2503 VN.n19 VN.n18 161.3
R2504 VN.n17 VN.n16 161.3
R2505 VN.n15 VN.n2 161.3
R2506 VN.n14 VN.n13 161.3
R2507 VN.n12 VN.n3 161.3
R2508 VN.n11 VN.n10 161.3
R2509 VN.n9 VN.n4 161.3
R2510 VN.n8 VN.n7 161.3
R2511 VN.n45 VN.n44 80.6037
R2512 VN.n22 VN.n21 80.6037
R2513 VN.n10 VN.n9 55.593
R2514 VN.n15 VN.n14 55.593
R2515 VN.n33 VN.n32 55.593
R2516 VN.n38 VN.n37 55.593
R2517 VN VN.n45 49.0407
R2518 VN.n6 VN.n5 48.5618
R2519 VN.n29 VN.n28 48.5618
R2520 VN.n20 VN.n19 37.1863
R2521 VN.n43 VN.n42 37.1863
R2522 VN.n30 VN.n29 29.6663
R2523 VN.n7 VN.n6 29.6663
R2524 VN.n21 VN.n20 29.2126
R2525 VN.n44 VN.n43 29.2126
R2526 VN.n9 VN.n8 25.5611
R2527 VN.n16 VN.n15 25.5611
R2528 VN.n32 VN.n31 25.5611
R2529 VN.n39 VN.n38 25.5611
R2530 VN.n10 VN.n3 24.5923
R2531 VN.n14 VN.n3 24.5923
R2532 VN.n37 VN.n26 24.5923
R2533 VN.n33 VN.n26 24.5923
R2534 VN.n19 VN.n1 15.2474
R2535 VN.n42 VN.n24 15.2474
R2536 VN.n8 VN.n5 9.3454
R2537 VN.n16 VN.n1 9.3454
R2538 VN.n31 VN.n28 9.3454
R2539 VN.n39 VN.n24 9.3454
R2540 VN.n45 VN.n23 0.285035
R2541 VN.n22 VN.n0 0.285035
R2542 VN.n41 VN.n23 0.189894
R2543 VN.n41 VN.n40 0.189894
R2544 VN.n40 VN.n25 0.189894
R2545 VN.n36 VN.n25 0.189894
R2546 VN.n36 VN.n35 0.189894
R2547 VN.n35 VN.n34 0.189894
R2548 VN.n34 VN.n27 0.189894
R2549 VN.n30 VN.n27 0.189894
R2550 VN.n7 VN.n4 0.189894
R2551 VN.n11 VN.n4 0.189894
R2552 VN.n12 VN.n11 0.189894
R2553 VN.n13 VN.n12 0.189894
R2554 VN.n13 VN.n2 0.189894
R2555 VN.n17 VN.n2 0.189894
R2556 VN.n18 VN.n17 0.189894
R2557 VN.n18 VN.n0 0.189894
R2558 VN VN.n22 0.146778
R2559 VDD2.n161 VDD2.n85 289.615
R2560 VDD2.n76 VDD2.n0 289.615
R2561 VDD2.n162 VDD2.n161 185
R2562 VDD2.n160 VDD2.n159 185
R2563 VDD2.n158 VDD2.n88 185
R2564 VDD2.n92 VDD2.n89 185
R2565 VDD2.n153 VDD2.n152 185
R2566 VDD2.n151 VDD2.n150 185
R2567 VDD2.n94 VDD2.n93 185
R2568 VDD2.n145 VDD2.n144 185
R2569 VDD2.n143 VDD2.n142 185
R2570 VDD2.n98 VDD2.n97 185
R2571 VDD2.n137 VDD2.n136 185
R2572 VDD2.n135 VDD2.n134 185
R2573 VDD2.n102 VDD2.n101 185
R2574 VDD2.n129 VDD2.n128 185
R2575 VDD2.n127 VDD2.n126 185
R2576 VDD2.n106 VDD2.n105 185
R2577 VDD2.n121 VDD2.n120 185
R2578 VDD2.n119 VDD2.n118 185
R2579 VDD2.n110 VDD2.n109 185
R2580 VDD2.n113 VDD2.n112 185
R2581 VDD2.n27 VDD2.n26 185
R2582 VDD2.n24 VDD2.n23 185
R2583 VDD2.n33 VDD2.n32 185
R2584 VDD2.n35 VDD2.n34 185
R2585 VDD2.n20 VDD2.n19 185
R2586 VDD2.n41 VDD2.n40 185
R2587 VDD2.n43 VDD2.n42 185
R2588 VDD2.n16 VDD2.n15 185
R2589 VDD2.n49 VDD2.n48 185
R2590 VDD2.n51 VDD2.n50 185
R2591 VDD2.n12 VDD2.n11 185
R2592 VDD2.n57 VDD2.n56 185
R2593 VDD2.n59 VDD2.n58 185
R2594 VDD2.n8 VDD2.n7 185
R2595 VDD2.n65 VDD2.n64 185
R2596 VDD2.n68 VDD2.n67 185
R2597 VDD2.n66 VDD2.n4 185
R2598 VDD2.n73 VDD2.n3 185
R2599 VDD2.n75 VDD2.n74 185
R2600 VDD2.n77 VDD2.n76 185
R2601 VDD2.t0 VDD2.n111 147.659
R2602 VDD2.t1 VDD2.n25 147.659
R2603 VDD2.n161 VDD2.n160 104.615
R2604 VDD2.n160 VDD2.n88 104.615
R2605 VDD2.n92 VDD2.n88 104.615
R2606 VDD2.n152 VDD2.n92 104.615
R2607 VDD2.n152 VDD2.n151 104.615
R2608 VDD2.n151 VDD2.n93 104.615
R2609 VDD2.n144 VDD2.n93 104.615
R2610 VDD2.n144 VDD2.n143 104.615
R2611 VDD2.n143 VDD2.n97 104.615
R2612 VDD2.n136 VDD2.n97 104.615
R2613 VDD2.n136 VDD2.n135 104.615
R2614 VDD2.n135 VDD2.n101 104.615
R2615 VDD2.n128 VDD2.n101 104.615
R2616 VDD2.n128 VDD2.n127 104.615
R2617 VDD2.n127 VDD2.n105 104.615
R2618 VDD2.n120 VDD2.n105 104.615
R2619 VDD2.n120 VDD2.n119 104.615
R2620 VDD2.n119 VDD2.n109 104.615
R2621 VDD2.n112 VDD2.n109 104.615
R2622 VDD2.n26 VDD2.n23 104.615
R2623 VDD2.n33 VDD2.n23 104.615
R2624 VDD2.n34 VDD2.n33 104.615
R2625 VDD2.n34 VDD2.n19 104.615
R2626 VDD2.n41 VDD2.n19 104.615
R2627 VDD2.n42 VDD2.n41 104.615
R2628 VDD2.n42 VDD2.n15 104.615
R2629 VDD2.n49 VDD2.n15 104.615
R2630 VDD2.n50 VDD2.n49 104.615
R2631 VDD2.n50 VDD2.n11 104.615
R2632 VDD2.n57 VDD2.n11 104.615
R2633 VDD2.n58 VDD2.n57 104.615
R2634 VDD2.n58 VDD2.n7 104.615
R2635 VDD2.n65 VDD2.n7 104.615
R2636 VDD2.n67 VDD2.n65 104.615
R2637 VDD2.n67 VDD2.n66 104.615
R2638 VDD2.n66 VDD2.n3 104.615
R2639 VDD2.n75 VDD2.n3 104.615
R2640 VDD2.n76 VDD2.n75 104.615
R2641 VDD2.n84 VDD2.n83 66.2249
R2642 VDD2 VDD2.n169 66.2221
R2643 VDD2.n168 VDD2.n167 65.1878
R2644 VDD2.n82 VDD2.n81 65.1876
R2645 VDD2.n82 VDD2.n80 54.5877
R2646 VDD2.n166 VDD2.n165 53.1308
R2647 VDD2.n112 VDD2.t0 52.3082
R2648 VDD2.n26 VDD2.t1 52.3082
R2649 VDD2.n166 VDD2.n84 43.4459
R2650 VDD2.n113 VDD2.n111 15.6677
R2651 VDD2.n27 VDD2.n25 15.6677
R2652 VDD2.n159 VDD2.n158 13.1884
R2653 VDD2.n74 VDD2.n73 13.1884
R2654 VDD2.n162 VDD2.n87 12.8005
R2655 VDD2.n157 VDD2.n89 12.8005
R2656 VDD2.n114 VDD2.n110 12.8005
R2657 VDD2.n28 VDD2.n24 12.8005
R2658 VDD2.n72 VDD2.n4 12.8005
R2659 VDD2.n77 VDD2.n2 12.8005
R2660 VDD2.n163 VDD2.n85 12.0247
R2661 VDD2.n154 VDD2.n153 12.0247
R2662 VDD2.n118 VDD2.n117 12.0247
R2663 VDD2.n32 VDD2.n31 12.0247
R2664 VDD2.n69 VDD2.n68 12.0247
R2665 VDD2.n78 VDD2.n0 12.0247
R2666 VDD2.n150 VDD2.n91 11.249
R2667 VDD2.n121 VDD2.n108 11.249
R2668 VDD2.n35 VDD2.n22 11.249
R2669 VDD2.n64 VDD2.n6 11.249
R2670 VDD2.n149 VDD2.n94 10.4732
R2671 VDD2.n122 VDD2.n106 10.4732
R2672 VDD2.n36 VDD2.n20 10.4732
R2673 VDD2.n63 VDD2.n8 10.4732
R2674 VDD2.n146 VDD2.n145 9.69747
R2675 VDD2.n126 VDD2.n125 9.69747
R2676 VDD2.n40 VDD2.n39 9.69747
R2677 VDD2.n60 VDD2.n59 9.69747
R2678 VDD2.n165 VDD2.n164 9.45567
R2679 VDD2.n80 VDD2.n79 9.45567
R2680 VDD2.n139 VDD2.n138 9.3005
R2681 VDD2.n141 VDD2.n140 9.3005
R2682 VDD2.n96 VDD2.n95 9.3005
R2683 VDD2.n147 VDD2.n146 9.3005
R2684 VDD2.n149 VDD2.n148 9.3005
R2685 VDD2.n91 VDD2.n90 9.3005
R2686 VDD2.n155 VDD2.n154 9.3005
R2687 VDD2.n157 VDD2.n156 9.3005
R2688 VDD2.n164 VDD2.n163 9.3005
R2689 VDD2.n87 VDD2.n86 9.3005
R2690 VDD2.n100 VDD2.n99 9.3005
R2691 VDD2.n133 VDD2.n132 9.3005
R2692 VDD2.n131 VDD2.n130 9.3005
R2693 VDD2.n104 VDD2.n103 9.3005
R2694 VDD2.n125 VDD2.n124 9.3005
R2695 VDD2.n123 VDD2.n122 9.3005
R2696 VDD2.n108 VDD2.n107 9.3005
R2697 VDD2.n117 VDD2.n116 9.3005
R2698 VDD2.n115 VDD2.n114 9.3005
R2699 VDD2.n79 VDD2.n78 9.3005
R2700 VDD2.n2 VDD2.n1 9.3005
R2701 VDD2.n47 VDD2.n46 9.3005
R2702 VDD2.n45 VDD2.n44 9.3005
R2703 VDD2.n18 VDD2.n17 9.3005
R2704 VDD2.n39 VDD2.n38 9.3005
R2705 VDD2.n37 VDD2.n36 9.3005
R2706 VDD2.n22 VDD2.n21 9.3005
R2707 VDD2.n31 VDD2.n30 9.3005
R2708 VDD2.n29 VDD2.n28 9.3005
R2709 VDD2.n14 VDD2.n13 9.3005
R2710 VDD2.n53 VDD2.n52 9.3005
R2711 VDD2.n55 VDD2.n54 9.3005
R2712 VDD2.n10 VDD2.n9 9.3005
R2713 VDD2.n61 VDD2.n60 9.3005
R2714 VDD2.n63 VDD2.n62 9.3005
R2715 VDD2.n6 VDD2.n5 9.3005
R2716 VDD2.n70 VDD2.n69 9.3005
R2717 VDD2.n72 VDD2.n71 9.3005
R2718 VDD2.n142 VDD2.n96 8.92171
R2719 VDD2.n129 VDD2.n104 8.92171
R2720 VDD2.n43 VDD2.n18 8.92171
R2721 VDD2.n56 VDD2.n10 8.92171
R2722 VDD2.n141 VDD2.n98 8.14595
R2723 VDD2.n130 VDD2.n102 8.14595
R2724 VDD2.n44 VDD2.n16 8.14595
R2725 VDD2.n55 VDD2.n12 8.14595
R2726 VDD2.n138 VDD2.n137 7.3702
R2727 VDD2.n134 VDD2.n133 7.3702
R2728 VDD2.n48 VDD2.n47 7.3702
R2729 VDD2.n52 VDD2.n51 7.3702
R2730 VDD2.n137 VDD2.n100 6.59444
R2731 VDD2.n134 VDD2.n100 6.59444
R2732 VDD2.n48 VDD2.n14 6.59444
R2733 VDD2.n51 VDD2.n14 6.59444
R2734 VDD2.n138 VDD2.n98 5.81868
R2735 VDD2.n133 VDD2.n102 5.81868
R2736 VDD2.n47 VDD2.n16 5.81868
R2737 VDD2.n52 VDD2.n12 5.81868
R2738 VDD2.n142 VDD2.n141 5.04292
R2739 VDD2.n130 VDD2.n129 5.04292
R2740 VDD2.n44 VDD2.n43 5.04292
R2741 VDD2.n56 VDD2.n55 5.04292
R2742 VDD2.n115 VDD2.n111 4.38563
R2743 VDD2.n29 VDD2.n25 4.38563
R2744 VDD2.n145 VDD2.n96 4.26717
R2745 VDD2.n126 VDD2.n104 4.26717
R2746 VDD2.n40 VDD2.n18 4.26717
R2747 VDD2.n59 VDD2.n10 4.26717
R2748 VDD2.n146 VDD2.n94 3.49141
R2749 VDD2.n125 VDD2.n106 3.49141
R2750 VDD2.n39 VDD2.n20 3.49141
R2751 VDD2.n60 VDD2.n8 3.49141
R2752 VDD2.n150 VDD2.n149 2.71565
R2753 VDD2.n122 VDD2.n121 2.71565
R2754 VDD2.n36 VDD2.n35 2.71565
R2755 VDD2.n64 VDD2.n63 2.71565
R2756 VDD2.n165 VDD2.n85 1.93989
R2757 VDD2.n153 VDD2.n91 1.93989
R2758 VDD2.n118 VDD2.n108 1.93989
R2759 VDD2.n32 VDD2.n22 1.93989
R2760 VDD2.n68 VDD2.n6 1.93989
R2761 VDD2.n80 VDD2.n0 1.93989
R2762 VDD2.n168 VDD2.n166 1.4574
R2763 VDD2.n169 VDD2.t7 1.33294
R2764 VDD2.n169 VDD2.t4 1.33294
R2765 VDD2.n167 VDD2.t9 1.33294
R2766 VDD2.n167 VDD2.t6 1.33294
R2767 VDD2.n83 VDD2.t5 1.33294
R2768 VDD2.n83 VDD2.t2 1.33294
R2769 VDD2.n81 VDD2.t8 1.33294
R2770 VDD2.n81 VDD2.t3 1.33294
R2771 VDD2.n163 VDD2.n162 1.16414
R2772 VDD2.n154 VDD2.n89 1.16414
R2773 VDD2.n117 VDD2.n110 1.16414
R2774 VDD2.n31 VDD2.n24 1.16414
R2775 VDD2.n69 VDD2.n4 1.16414
R2776 VDD2.n78 VDD2.n77 1.16414
R2777 VDD2 VDD2.n168 0.422914
R2778 VDD2.n159 VDD2.n87 0.388379
R2779 VDD2.n158 VDD2.n157 0.388379
R2780 VDD2.n114 VDD2.n113 0.388379
R2781 VDD2.n28 VDD2.n27 0.388379
R2782 VDD2.n73 VDD2.n72 0.388379
R2783 VDD2.n74 VDD2.n2 0.388379
R2784 VDD2.n84 VDD2.n82 0.309378
R2785 VDD2.n164 VDD2.n86 0.155672
R2786 VDD2.n156 VDD2.n86 0.155672
R2787 VDD2.n156 VDD2.n155 0.155672
R2788 VDD2.n155 VDD2.n90 0.155672
R2789 VDD2.n148 VDD2.n90 0.155672
R2790 VDD2.n148 VDD2.n147 0.155672
R2791 VDD2.n147 VDD2.n95 0.155672
R2792 VDD2.n140 VDD2.n95 0.155672
R2793 VDD2.n140 VDD2.n139 0.155672
R2794 VDD2.n139 VDD2.n99 0.155672
R2795 VDD2.n132 VDD2.n99 0.155672
R2796 VDD2.n132 VDD2.n131 0.155672
R2797 VDD2.n131 VDD2.n103 0.155672
R2798 VDD2.n124 VDD2.n103 0.155672
R2799 VDD2.n124 VDD2.n123 0.155672
R2800 VDD2.n123 VDD2.n107 0.155672
R2801 VDD2.n116 VDD2.n107 0.155672
R2802 VDD2.n116 VDD2.n115 0.155672
R2803 VDD2.n30 VDD2.n29 0.155672
R2804 VDD2.n30 VDD2.n21 0.155672
R2805 VDD2.n37 VDD2.n21 0.155672
R2806 VDD2.n38 VDD2.n37 0.155672
R2807 VDD2.n38 VDD2.n17 0.155672
R2808 VDD2.n45 VDD2.n17 0.155672
R2809 VDD2.n46 VDD2.n45 0.155672
R2810 VDD2.n46 VDD2.n13 0.155672
R2811 VDD2.n53 VDD2.n13 0.155672
R2812 VDD2.n54 VDD2.n53 0.155672
R2813 VDD2.n54 VDD2.n9 0.155672
R2814 VDD2.n61 VDD2.n9 0.155672
R2815 VDD2.n62 VDD2.n61 0.155672
R2816 VDD2.n62 VDD2.n5 0.155672
R2817 VDD2.n70 VDD2.n5 0.155672
R2818 VDD2.n71 VDD2.n70 0.155672
R2819 VDD2.n71 VDD2.n1 0.155672
R2820 VDD2.n79 VDD2.n1 0.155672
C0 VDD2 VTAIL 13.098f
C1 VP VDD1 11.2534f
C2 VN VDD1 0.150731f
C3 VP VTAIL 11.010799f
C4 VP VDD2 0.426086f
C5 VN VTAIL 10.9963f
C6 VN VDD2 10.982901f
C7 VP VN 7.09151f
C8 VTAIL VDD1 13.0585f
C9 VDD2 VDD1 1.3681f
C10 VDD2 B 6.263457f
C11 VDD1 B 6.233797f
C12 VTAIL B 8.260687f
C13 VN B 12.657869f
C14 VP B 10.877342f
C15 VDD2.n0 B 0.032063f
C16 VDD2.n1 B 0.022594f
C17 VDD2.n2 B 0.012141f
C18 VDD2.n3 B 0.028697f
C19 VDD2.n4 B 0.012855f
C20 VDD2.n5 B 0.022594f
C21 VDD2.n6 B 0.012141f
C22 VDD2.n7 B 0.028697f
C23 VDD2.n8 B 0.012855f
C24 VDD2.n9 B 0.022594f
C25 VDD2.n10 B 0.012141f
C26 VDD2.n11 B 0.028697f
C27 VDD2.n12 B 0.012855f
C28 VDD2.n13 B 0.022594f
C29 VDD2.n14 B 0.012141f
C30 VDD2.n15 B 0.028697f
C31 VDD2.n16 B 0.012855f
C32 VDD2.n17 B 0.022594f
C33 VDD2.n18 B 0.012141f
C34 VDD2.n19 B 0.028697f
C35 VDD2.n20 B 0.012855f
C36 VDD2.n21 B 0.022594f
C37 VDD2.n22 B 0.012141f
C38 VDD2.n23 B 0.028697f
C39 VDD2.n24 B 0.012855f
C40 VDD2.n25 B 0.146571f
C41 VDD2.t1 B 0.047307f
C42 VDD2.n26 B 0.021523f
C43 VDD2.n27 B 0.016952f
C44 VDD2.n28 B 0.012141f
C45 VDD2.n29 B 1.45551f
C46 VDD2.n30 B 0.022594f
C47 VDD2.n31 B 0.012141f
C48 VDD2.n32 B 0.012855f
C49 VDD2.n33 B 0.028697f
C50 VDD2.n34 B 0.028697f
C51 VDD2.n35 B 0.012855f
C52 VDD2.n36 B 0.012141f
C53 VDD2.n37 B 0.022594f
C54 VDD2.n38 B 0.022594f
C55 VDD2.n39 B 0.012141f
C56 VDD2.n40 B 0.012855f
C57 VDD2.n41 B 0.028697f
C58 VDD2.n42 B 0.028697f
C59 VDD2.n43 B 0.012855f
C60 VDD2.n44 B 0.012141f
C61 VDD2.n45 B 0.022594f
C62 VDD2.n46 B 0.022594f
C63 VDD2.n47 B 0.012141f
C64 VDD2.n48 B 0.012855f
C65 VDD2.n49 B 0.028697f
C66 VDD2.n50 B 0.028697f
C67 VDD2.n51 B 0.012855f
C68 VDD2.n52 B 0.012141f
C69 VDD2.n53 B 0.022594f
C70 VDD2.n54 B 0.022594f
C71 VDD2.n55 B 0.012141f
C72 VDD2.n56 B 0.012855f
C73 VDD2.n57 B 0.028697f
C74 VDD2.n58 B 0.028697f
C75 VDD2.n59 B 0.012855f
C76 VDD2.n60 B 0.012141f
C77 VDD2.n61 B 0.022594f
C78 VDD2.n62 B 0.022594f
C79 VDD2.n63 B 0.012141f
C80 VDD2.n64 B 0.012855f
C81 VDD2.n65 B 0.028697f
C82 VDD2.n66 B 0.028697f
C83 VDD2.n67 B 0.028697f
C84 VDD2.n68 B 0.012855f
C85 VDD2.n69 B 0.012141f
C86 VDD2.n70 B 0.022594f
C87 VDD2.n71 B 0.022594f
C88 VDD2.n72 B 0.012141f
C89 VDD2.n73 B 0.012498f
C90 VDD2.n74 B 0.012498f
C91 VDD2.n75 B 0.028697f
C92 VDD2.n76 B 0.062664f
C93 VDD2.n77 B 0.012855f
C94 VDD2.n78 B 0.012141f
C95 VDD2.n79 B 0.059016f
C96 VDD2.n80 B 0.054966f
C97 VDD2.t8 B 0.265319f
C98 VDD2.t3 B 0.265319f
C99 VDD2.n81 B 2.40111f
C100 VDD2.n82 B 0.460549f
C101 VDD2.t5 B 0.265319f
C102 VDD2.t2 B 0.265319f
C103 VDD2.n83 B 2.40694f
C104 VDD2.n84 B 2.19184f
C105 VDD2.n85 B 0.032063f
C106 VDD2.n86 B 0.022594f
C107 VDD2.n87 B 0.012141f
C108 VDD2.n88 B 0.028697f
C109 VDD2.n89 B 0.012855f
C110 VDD2.n90 B 0.022594f
C111 VDD2.n91 B 0.012141f
C112 VDD2.n92 B 0.028697f
C113 VDD2.n93 B 0.028697f
C114 VDD2.n94 B 0.012855f
C115 VDD2.n95 B 0.022594f
C116 VDD2.n96 B 0.012141f
C117 VDD2.n97 B 0.028697f
C118 VDD2.n98 B 0.012855f
C119 VDD2.n99 B 0.022594f
C120 VDD2.n100 B 0.012141f
C121 VDD2.n101 B 0.028697f
C122 VDD2.n102 B 0.012855f
C123 VDD2.n103 B 0.022594f
C124 VDD2.n104 B 0.012141f
C125 VDD2.n105 B 0.028697f
C126 VDD2.n106 B 0.012855f
C127 VDD2.n107 B 0.022594f
C128 VDD2.n108 B 0.012141f
C129 VDD2.n109 B 0.028697f
C130 VDD2.n110 B 0.012855f
C131 VDD2.n111 B 0.146571f
C132 VDD2.t0 B 0.047307f
C133 VDD2.n112 B 0.021523f
C134 VDD2.n113 B 0.016952f
C135 VDD2.n114 B 0.012141f
C136 VDD2.n115 B 1.45551f
C137 VDD2.n116 B 0.022594f
C138 VDD2.n117 B 0.012141f
C139 VDD2.n118 B 0.012855f
C140 VDD2.n119 B 0.028697f
C141 VDD2.n120 B 0.028697f
C142 VDD2.n121 B 0.012855f
C143 VDD2.n122 B 0.012141f
C144 VDD2.n123 B 0.022594f
C145 VDD2.n124 B 0.022594f
C146 VDD2.n125 B 0.012141f
C147 VDD2.n126 B 0.012855f
C148 VDD2.n127 B 0.028697f
C149 VDD2.n128 B 0.028697f
C150 VDD2.n129 B 0.012855f
C151 VDD2.n130 B 0.012141f
C152 VDD2.n131 B 0.022594f
C153 VDD2.n132 B 0.022594f
C154 VDD2.n133 B 0.012141f
C155 VDD2.n134 B 0.012855f
C156 VDD2.n135 B 0.028697f
C157 VDD2.n136 B 0.028697f
C158 VDD2.n137 B 0.012855f
C159 VDD2.n138 B 0.012141f
C160 VDD2.n139 B 0.022594f
C161 VDD2.n140 B 0.022594f
C162 VDD2.n141 B 0.012141f
C163 VDD2.n142 B 0.012855f
C164 VDD2.n143 B 0.028697f
C165 VDD2.n144 B 0.028697f
C166 VDD2.n145 B 0.012855f
C167 VDD2.n146 B 0.012141f
C168 VDD2.n147 B 0.022594f
C169 VDD2.n148 B 0.022594f
C170 VDD2.n149 B 0.012141f
C171 VDD2.n150 B 0.012855f
C172 VDD2.n151 B 0.028697f
C173 VDD2.n152 B 0.028697f
C174 VDD2.n153 B 0.012855f
C175 VDD2.n154 B 0.012141f
C176 VDD2.n155 B 0.022594f
C177 VDD2.n156 B 0.022594f
C178 VDD2.n157 B 0.012141f
C179 VDD2.n158 B 0.012498f
C180 VDD2.n159 B 0.012498f
C181 VDD2.n160 B 0.028697f
C182 VDD2.n161 B 0.062664f
C183 VDD2.n162 B 0.012855f
C184 VDD2.n163 B 0.012141f
C185 VDD2.n164 B 0.059016f
C186 VDD2.n165 B 0.05087f
C187 VDD2.n166 B 2.38074f
C188 VDD2.t9 B 0.265319f
C189 VDD2.t6 B 0.265319f
C190 VDD2.n167 B 2.40112f
C191 VDD2.n168 B 0.317743f
C192 VDD2.t7 B 0.265319f
C193 VDD2.t4 B 0.265319f
C194 VDD2.n169 B 2.40692f
C195 VN.n0 B 0.041701f
C196 VN.t4 B 1.73026f
C197 VN.n1 B 0.618599f
C198 VN.n2 B 0.031251f
C199 VN.t6 B 1.73026f
C200 VN.n3 B 0.647941f
C201 VN.n4 B 0.031251f
C202 VN.t1 B 1.73026f
C203 VN.n5 B 0.658166f
C204 VN.t8 B 1.83664f
C205 VN.n6 B 0.676923f
C206 VN.n7 B 0.166693f
C207 VN.n8 B 0.041255f
C208 VN.n9 B 0.036331f
C209 VN.n10 B 0.053485f
C210 VN.n11 B 0.031251f
C211 VN.n12 B 0.031251f
C212 VN.n13 B 0.031251f
C213 VN.n14 B 0.053485f
C214 VN.n15 B 0.036331f
C215 VN.n16 B 0.041255f
C216 VN.n17 B 0.031251f
C217 VN.n18 B 0.031251f
C218 VN.n19 B 0.051732f
C219 VN.n20 B 0.018678f
C220 VN.t7 B 1.79498f
C221 VN.n21 B 0.686229f
C222 VN.n22 B 0.029268f
C223 VN.n23 B 0.041701f
C224 VN.t0 B 1.73026f
C225 VN.n24 B 0.618599f
C226 VN.n25 B 0.031251f
C227 VN.t3 B 1.73026f
C228 VN.n26 B 0.647941f
C229 VN.n27 B 0.031251f
C230 VN.t2 B 1.73026f
C231 VN.n28 B 0.658166f
C232 VN.t5 B 1.83664f
C233 VN.n29 B 0.676923f
C234 VN.n30 B 0.166693f
C235 VN.n31 B 0.041255f
C236 VN.n32 B 0.036331f
C237 VN.n33 B 0.053485f
C238 VN.n34 B 0.031251f
C239 VN.n35 B 0.031251f
C240 VN.n36 B 0.031251f
C241 VN.n37 B 0.053485f
C242 VN.n38 B 0.036331f
C243 VN.n39 B 0.041255f
C244 VN.n40 B 0.031251f
C245 VN.n41 B 0.031251f
C246 VN.n42 B 0.051732f
C247 VN.n43 B 0.018678f
C248 VN.t9 B 1.79498f
C249 VN.n44 B 0.686229f
C250 VN.n45 B 1.66362f
C251 VTAIL.t7 B 0.281706f
C252 VTAIL.t1 B 0.281706f
C253 VTAIL.n0 B 2.48493f
C254 VTAIL.n1 B 0.40557f
C255 VTAIL.n2 B 0.034043f
C256 VTAIL.n3 B 0.02399f
C257 VTAIL.n4 B 0.012891f
C258 VTAIL.n5 B 0.03047f
C259 VTAIL.n6 B 0.013649f
C260 VTAIL.n7 B 0.02399f
C261 VTAIL.n8 B 0.012891f
C262 VTAIL.n9 B 0.03047f
C263 VTAIL.n10 B 0.013649f
C264 VTAIL.n11 B 0.02399f
C265 VTAIL.n12 B 0.012891f
C266 VTAIL.n13 B 0.03047f
C267 VTAIL.n14 B 0.013649f
C268 VTAIL.n15 B 0.02399f
C269 VTAIL.n16 B 0.012891f
C270 VTAIL.n17 B 0.03047f
C271 VTAIL.n18 B 0.013649f
C272 VTAIL.n19 B 0.02399f
C273 VTAIL.n20 B 0.012891f
C274 VTAIL.n21 B 0.03047f
C275 VTAIL.n22 B 0.013649f
C276 VTAIL.n23 B 0.02399f
C277 VTAIL.n24 B 0.012891f
C278 VTAIL.n25 B 0.03047f
C279 VTAIL.n26 B 0.013649f
C280 VTAIL.n27 B 0.155624f
C281 VTAIL.t13 B 0.050229f
C282 VTAIL.n28 B 0.022852f
C283 VTAIL.n29 B 0.017999f
C284 VTAIL.n30 B 0.012891f
C285 VTAIL.n31 B 1.54541f
C286 VTAIL.n32 B 0.02399f
C287 VTAIL.n33 B 0.012891f
C288 VTAIL.n34 B 0.013649f
C289 VTAIL.n35 B 0.03047f
C290 VTAIL.n36 B 0.03047f
C291 VTAIL.n37 B 0.013649f
C292 VTAIL.n38 B 0.012891f
C293 VTAIL.n39 B 0.02399f
C294 VTAIL.n40 B 0.02399f
C295 VTAIL.n41 B 0.012891f
C296 VTAIL.n42 B 0.013649f
C297 VTAIL.n43 B 0.03047f
C298 VTAIL.n44 B 0.03047f
C299 VTAIL.n45 B 0.013649f
C300 VTAIL.n46 B 0.012891f
C301 VTAIL.n47 B 0.02399f
C302 VTAIL.n48 B 0.02399f
C303 VTAIL.n49 B 0.012891f
C304 VTAIL.n50 B 0.013649f
C305 VTAIL.n51 B 0.03047f
C306 VTAIL.n52 B 0.03047f
C307 VTAIL.n53 B 0.013649f
C308 VTAIL.n54 B 0.012891f
C309 VTAIL.n55 B 0.02399f
C310 VTAIL.n56 B 0.02399f
C311 VTAIL.n57 B 0.012891f
C312 VTAIL.n58 B 0.013649f
C313 VTAIL.n59 B 0.03047f
C314 VTAIL.n60 B 0.03047f
C315 VTAIL.n61 B 0.013649f
C316 VTAIL.n62 B 0.012891f
C317 VTAIL.n63 B 0.02399f
C318 VTAIL.n64 B 0.02399f
C319 VTAIL.n65 B 0.012891f
C320 VTAIL.n66 B 0.013649f
C321 VTAIL.n67 B 0.03047f
C322 VTAIL.n68 B 0.03047f
C323 VTAIL.n69 B 0.03047f
C324 VTAIL.n70 B 0.013649f
C325 VTAIL.n71 B 0.012891f
C326 VTAIL.n72 B 0.02399f
C327 VTAIL.n73 B 0.02399f
C328 VTAIL.n74 B 0.012891f
C329 VTAIL.n75 B 0.01327f
C330 VTAIL.n76 B 0.01327f
C331 VTAIL.n77 B 0.03047f
C332 VTAIL.n78 B 0.066534f
C333 VTAIL.n79 B 0.013649f
C334 VTAIL.n80 B 0.012891f
C335 VTAIL.n81 B 0.062661f
C336 VTAIL.n82 B 0.037497f
C337 VTAIL.n83 B 0.229815f
C338 VTAIL.t10 B 0.281706f
C339 VTAIL.t19 B 0.281706f
C340 VTAIL.n84 B 2.48493f
C341 VTAIL.n85 B 0.449218f
C342 VTAIL.t14 B 0.281706f
C343 VTAIL.t16 B 0.281706f
C344 VTAIL.n86 B 2.48493f
C345 VTAIL.n87 B 1.87795f
C346 VTAIL.t9 B 0.281706f
C347 VTAIL.t5 B 0.281706f
C348 VTAIL.n88 B 2.48495f
C349 VTAIL.n89 B 1.87794f
C350 VTAIL.t2 B 0.281706f
C351 VTAIL.t8 B 0.281706f
C352 VTAIL.n90 B 2.48495f
C353 VTAIL.n91 B 0.449206f
C354 VTAIL.n92 B 0.034043f
C355 VTAIL.n93 B 0.02399f
C356 VTAIL.n94 B 0.012891f
C357 VTAIL.n95 B 0.03047f
C358 VTAIL.n96 B 0.013649f
C359 VTAIL.n97 B 0.02399f
C360 VTAIL.n98 B 0.012891f
C361 VTAIL.n99 B 0.03047f
C362 VTAIL.n100 B 0.03047f
C363 VTAIL.n101 B 0.013649f
C364 VTAIL.n102 B 0.02399f
C365 VTAIL.n103 B 0.012891f
C366 VTAIL.n104 B 0.03047f
C367 VTAIL.n105 B 0.013649f
C368 VTAIL.n106 B 0.02399f
C369 VTAIL.n107 B 0.012891f
C370 VTAIL.n108 B 0.03047f
C371 VTAIL.n109 B 0.013649f
C372 VTAIL.n110 B 0.02399f
C373 VTAIL.n111 B 0.012891f
C374 VTAIL.n112 B 0.03047f
C375 VTAIL.n113 B 0.013649f
C376 VTAIL.n114 B 0.02399f
C377 VTAIL.n115 B 0.012891f
C378 VTAIL.n116 B 0.03047f
C379 VTAIL.n117 B 0.013649f
C380 VTAIL.n118 B 0.155624f
C381 VTAIL.t4 B 0.050229f
C382 VTAIL.n119 B 0.022852f
C383 VTAIL.n120 B 0.017999f
C384 VTAIL.n121 B 0.012891f
C385 VTAIL.n122 B 1.54541f
C386 VTAIL.n123 B 0.02399f
C387 VTAIL.n124 B 0.012891f
C388 VTAIL.n125 B 0.013649f
C389 VTAIL.n126 B 0.03047f
C390 VTAIL.n127 B 0.03047f
C391 VTAIL.n128 B 0.013649f
C392 VTAIL.n129 B 0.012891f
C393 VTAIL.n130 B 0.02399f
C394 VTAIL.n131 B 0.02399f
C395 VTAIL.n132 B 0.012891f
C396 VTAIL.n133 B 0.013649f
C397 VTAIL.n134 B 0.03047f
C398 VTAIL.n135 B 0.03047f
C399 VTAIL.n136 B 0.013649f
C400 VTAIL.n137 B 0.012891f
C401 VTAIL.n138 B 0.02399f
C402 VTAIL.n139 B 0.02399f
C403 VTAIL.n140 B 0.012891f
C404 VTAIL.n141 B 0.013649f
C405 VTAIL.n142 B 0.03047f
C406 VTAIL.n143 B 0.03047f
C407 VTAIL.n144 B 0.013649f
C408 VTAIL.n145 B 0.012891f
C409 VTAIL.n146 B 0.02399f
C410 VTAIL.n147 B 0.02399f
C411 VTAIL.n148 B 0.012891f
C412 VTAIL.n149 B 0.013649f
C413 VTAIL.n150 B 0.03047f
C414 VTAIL.n151 B 0.03047f
C415 VTAIL.n152 B 0.013649f
C416 VTAIL.n153 B 0.012891f
C417 VTAIL.n154 B 0.02399f
C418 VTAIL.n155 B 0.02399f
C419 VTAIL.n156 B 0.012891f
C420 VTAIL.n157 B 0.013649f
C421 VTAIL.n158 B 0.03047f
C422 VTAIL.n159 B 0.03047f
C423 VTAIL.n160 B 0.013649f
C424 VTAIL.n161 B 0.012891f
C425 VTAIL.n162 B 0.02399f
C426 VTAIL.n163 B 0.02399f
C427 VTAIL.n164 B 0.012891f
C428 VTAIL.n165 B 0.01327f
C429 VTAIL.n166 B 0.01327f
C430 VTAIL.n167 B 0.03047f
C431 VTAIL.n168 B 0.066534f
C432 VTAIL.n169 B 0.013649f
C433 VTAIL.n170 B 0.012891f
C434 VTAIL.n171 B 0.062661f
C435 VTAIL.n172 B 0.037497f
C436 VTAIL.n173 B 0.229815f
C437 VTAIL.t12 B 0.281706f
C438 VTAIL.t15 B 0.281706f
C439 VTAIL.n174 B 2.48495f
C440 VTAIL.n175 B 0.429215f
C441 VTAIL.t17 B 0.281706f
C442 VTAIL.t18 B 0.281706f
C443 VTAIL.n176 B 2.48495f
C444 VTAIL.n177 B 0.449206f
C445 VTAIL.n178 B 0.034043f
C446 VTAIL.n179 B 0.02399f
C447 VTAIL.n180 B 0.012891f
C448 VTAIL.n181 B 0.03047f
C449 VTAIL.n182 B 0.013649f
C450 VTAIL.n183 B 0.02399f
C451 VTAIL.n184 B 0.012891f
C452 VTAIL.n185 B 0.03047f
C453 VTAIL.n186 B 0.03047f
C454 VTAIL.n187 B 0.013649f
C455 VTAIL.n188 B 0.02399f
C456 VTAIL.n189 B 0.012891f
C457 VTAIL.n190 B 0.03047f
C458 VTAIL.n191 B 0.013649f
C459 VTAIL.n192 B 0.02399f
C460 VTAIL.n193 B 0.012891f
C461 VTAIL.n194 B 0.03047f
C462 VTAIL.n195 B 0.013649f
C463 VTAIL.n196 B 0.02399f
C464 VTAIL.n197 B 0.012891f
C465 VTAIL.n198 B 0.03047f
C466 VTAIL.n199 B 0.013649f
C467 VTAIL.n200 B 0.02399f
C468 VTAIL.n201 B 0.012891f
C469 VTAIL.n202 B 0.03047f
C470 VTAIL.n203 B 0.013649f
C471 VTAIL.n204 B 0.155624f
C472 VTAIL.t11 B 0.050229f
C473 VTAIL.n205 B 0.022852f
C474 VTAIL.n206 B 0.017999f
C475 VTAIL.n207 B 0.012891f
C476 VTAIL.n208 B 1.54541f
C477 VTAIL.n209 B 0.02399f
C478 VTAIL.n210 B 0.012891f
C479 VTAIL.n211 B 0.013649f
C480 VTAIL.n212 B 0.03047f
C481 VTAIL.n213 B 0.03047f
C482 VTAIL.n214 B 0.013649f
C483 VTAIL.n215 B 0.012891f
C484 VTAIL.n216 B 0.02399f
C485 VTAIL.n217 B 0.02399f
C486 VTAIL.n218 B 0.012891f
C487 VTAIL.n219 B 0.013649f
C488 VTAIL.n220 B 0.03047f
C489 VTAIL.n221 B 0.03047f
C490 VTAIL.n222 B 0.013649f
C491 VTAIL.n223 B 0.012891f
C492 VTAIL.n224 B 0.02399f
C493 VTAIL.n225 B 0.02399f
C494 VTAIL.n226 B 0.012891f
C495 VTAIL.n227 B 0.013649f
C496 VTAIL.n228 B 0.03047f
C497 VTAIL.n229 B 0.03047f
C498 VTAIL.n230 B 0.013649f
C499 VTAIL.n231 B 0.012891f
C500 VTAIL.n232 B 0.02399f
C501 VTAIL.n233 B 0.02399f
C502 VTAIL.n234 B 0.012891f
C503 VTAIL.n235 B 0.013649f
C504 VTAIL.n236 B 0.03047f
C505 VTAIL.n237 B 0.03047f
C506 VTAIL.n238 B 0.013649f
C507 VTAIL.n239 B 0.012891f
C508 VTAIL.n240 B 0.02399f
C509 VTAIL.n241 B 0.02399f
C510 VTAIL.n242 B 0.012891f
C511 VTAIL.n243 B 0.013649f
C512 VTAIL.n244 B 0.03047f
C513 VTAIL.n245 B 0.03047f
C514 VTAIL.n246 B 0.013649f
C515 VTAIL.n247 B 0.012891f
C516 VTAIL.n248 B 0.02399f
C517 VTAIL.n249 B 0.02399f
C518 VTAIL.n250 B 0.012891f
C519 VTAIL.n251 B 0.01327f
C520 VTAIL.n252 B 0.01327f
C521 VTAIL.n253 B 0.03047f
C522 VTAIL.n254 B 0.066534f
C523 VTAIL.n255 B 0.013649f
C524 VTAIL.n256 B 0.012891f
C525 VTAIL.n257 B 0.062661f
C526 VTAIL.n258 B 0.037497f
C527 VTAIL.n259 B 1.56592f
C528 VTAIL.n260 B 0.034043f
C529 VTAIL.n261 B 0.02399f
C530 VTAIL.n262 B 0.012891f
C531 VTAIL.n263 B 0.03047f
C532 VTAIL.n264 B 0.013649f
C533 VTAIL.n265 B 0.02399f
C534 VTAIL.n266 B 0.012891f
C535 VTAIL.n267 B 0.03047f
C536 VTAIL.n268 B 0.013649f
C537 VTAIL.n269 B 0.02399f
C538 VTAIL.n270 B 0.012891f
C539 VTAIL.n271 B 0.03047f
C540 VTAIL.n272 B 0.013649f
C541 VTAIL.n273 B 0.02399f
C542 VTAIL.n274 B 0.012891f
C543 VTAIL.n275 B 0.03047f
C544 VTAIL.n276 B 0.013649f
C545 VTAIL.n277 B 0.02399f
C546 VTAIL.n278 B 0.012891f
C547 VTAIL.n279 B 0.03047f
C548 VTAIL.n280 B 0.013649f
C549 VTAIL.n281 B 0.02399f
C550 VTAIL.n282 B 0.012891f
C551 VTAIL.n283 B 0.03047f
C552 VTAIL.n284 B 0.013649f
C553 VTAIL.n285 B 0.155624f
C554 VTAIL.t6 B 0.050229f
C555 VTAIL.n286 B 0.022852f
C556 VTAIL.n287 B 0.017999f
C557 VTAIL.n288 B 0.012891f
C558 VTAIL.n289 B 1.54541f
C559 VTAIL.n290 B 0.02399f
C560 VTAIL.n291 B 0.012891f
C561 VTAIL.n292 B 0.013649f
C562 VTAIL.n293 B 0.03047f
C563 VTAIL.n294 B 0.03047f
C564 VTAIL.n295 B 0.013649f
C565 VTAIL.n296 B 0.012891f
C566 VTAIL.n297 B 0.02399f
C567 VTAIL.n298 B 0.02399f
C568 VTAIL.n299 B 0.012891f
C569 VTAIL.n300 B 0.013649f
C570 VTAIL.n301 B 0.03047f
C571 VTAIL.n302 B 0.03047f
C572 VTAIL.n303 B 0.013649f
C573 VTAIL.n304 B 0.012891f
C574 VTAIL.n305 B 0.02399f
C575 VTAIL.n306 B 0.02399f
C576 VTAIL.n307 B 0.012891f
C577 VTAIL.n308 B 0.013649f
C578 VTAIL.n309 B 0.03047f
C579 VTAIL.n310 B 0.03047f
C580 VTAIL.n311 B 0.013649f
C581 VTAIL.n312 B 0.012891f
C582 VTAIL.n313 B 0.02399f
C583 VTAIL.n314 B 0.02399f
C584 VTAIL.n315 B 0.012891f
C585 VTAIL.n316 B 0.013649f
C586 VTAIL.n317 B 0.03047f
C587 VTAIL.n318 B 0.03047f
C588 VTAIL.n319 B 0.013649f
C589 VTAIL.n320 B 0.012891f
C590 VTAIL.n321 B 0.02399f
C591 VTAIL.n322 B 0.02399f
C592 VTAIL.n323 B 0.012891f
C593 VTAIL.n324 B 0.013649f
C594 VTAIL.n325 B 0.03047f
C595 VTAIL.n326 B 0.03047f
C596 VTAIL.n327 B 0.03047f
C597 VTAIL.n328 B 0.013649f
C598 VTAIL.n329 B 0.012891f
C599 VTAIL.n330 B 0.02399f
C600 VTAIL.n331 B 0.02399f
C601 VTAIL.n332 B 0.012891f
C602 VTAIL.n333 B 0.01327f
C603 VTAIL.n334 B 0.01327f
C604 VTAIL.n335 B 0.03047f
C605 VTAIL.n336 B 0.066534f
C606 VTAIL.n337 B 0.013649f
C607 VTAIL.n338 B 0.012891f
C608 VTAIL.n339 B 0.062661f
C609 VTAIL.n340 B 0.037497f
C610 VTAIL.n341 B 1.56592f
C611 VTAIL.t0 B 0.281706f
C612 VTAIL.t3 B 0.281706f
C613 VTAIL.n342 B 2.48493f
C614 VTAIL.n343 B 0.360256f
C615 VDD1.n0 B 0.03235f
C616 VDD1.n1 B 0.022796f
C617 VDD1.n2 B 0.01225f
C618 VDD1.n3 B 0.028954f
C619 VDD1.n4 B 0.01297f
C620 VDD1.n5 B 0.022796f
C621 VDD1.n6 B 0.01225f
C622 VDD1.n7 B 0.028954f
C623 VDD1.n8 B 0.028954f
C624 VDD1.n9 B 0.01297f
C625 VDD1.n10 B 0.022796f
C626 VDD1.n11 B 0.01225f
C627 VDD1.n12 B 0.028954f
C628 VDD1.n13 B 0.01297f
C629 VDD1.n14 B 0.022796f
C630 VDD1.n15 B 0.01225f
C631 VDD1.n16 B 0.028954f
C632 VDD1.n17 B 0.01297f
C633 VDD1.n18 B 0.022796f
C634 VDD1.n19 B 0.01225f
C635 VDD1.n20 B 0.028954f
C636 VDD1.n21 B 0.01297f
C637 VDD1.n22 B 0.022796f
C638 VDD1.n23 B 0.01225f
C639 VDD1.n24 B 0.028954f
C640 VDD1.n25 B 0.01297f
C641 VDD1.n26 B 0.147883f
C642 VDD1.t6 B 0.047731f
C643 VDD1.n27 B 0.021716f
C644 VDD1.n28 B 0.017104f
C645 VDD1.n29 B 0.01225f
C646 VDD1.n30 B 1.46855f
C647 VDD1.n31 B 0.022796f
C648 VDD1.n32 B 0.01225f
C649 VDD1.n33 B 0.01297f
C650 VDD1.n34 B 0.028954f
C651 VDD1.n35 B 0.028954f
C652 VDD1.n36 B 0.01297f
C653 VDD1.n37 B 0.01225f
C654 VDD1.n38 B 0.022796f
C655 VDD1.n39 B 0.022796f
C656 VDD1.n40 B 0.01225f
C657 VDD1.n41 B 0.01297f
C658 VDD1.n42 B 0.028954f
C659 VDD1.n43 B 0.028954f
C660 VDD1.n44 B 0.01297f
C661 VDD1.n45 B 0.01225f
C662 VDD1.n46 B 0.022796f
C663 VDD1.n47 B 0.022796f
C664 VDD1.n48 B 0.01225f
C665 VDD1.n49 B 0.01297f
C666 VDD1.n50 B 0.028954f
C667 VDD1.n51 B 0.028954f
C668 VDD1.n52 B 0.01297f
C669 VDD1.n53 B 0.01225f
C670 VDD1.n54 B 0.022796f
C671 VDD1.n55 B 0.022796f
C672 VDD1.n56 B 0.01225f
C673 VDD1.n57 B 0.01297f
C674 VDD1.n58 B 0.028954f
C675 VDD1.n59 B 0.028954f
C676 VDD1.n60 B 0.01297f
C677 VDD1.n61 B 0.01225f
C678 VDD1.n62 B 0.022796f
C679 VDD1.n63 B 0.022796f
C680 VDD1.n64 B 0.01225f
C681 VDD1.n65 B 0.01297f
C682 VDD1.n66 B 0.028954f
C683 VDD1.n67 B 0.028954f
C684 VDD1.n68 B 0.01297f
C685 VDD1.n69 B 0.01225f
C686 VDD1.n70 B 0.022796f
C687 VDD1.n71 B 0.022796f
C688 VDD1.n72 B 0.01225f
C689 VDD1.n73 B 0.01261f
C690 VDD1.n74 B 0.01261f
C691 VDD1.n75 B 0.028954f
C692 VDD1.n76 B 0.063225f
C693 VDD1.n77 B 0.01297f
C694 VDD1.n78 B 0.01225f
C695 VDD1.n79 B 0.059544f
C696 VDD1.n80 B 0.055458f
C697 VDD1.t3 B 0.267695f
C698 VDD1.t9 B 0.267695f
C699 VDD1.n81 B 2.42262f
C700 VDD1.n82 B 0.471294f
C701 VDD1.n83 B 0.03235f
C702 VDD1.n84 B 0.022796f
C703 VDD1.n85 B 0.01225f
C704 VDD1.n86 B 0.028954f
C705 VDD1.n87 B 0.01297f
C706 VDD1.n88 B 0.022796f
C707 VDD1.n89 B 0.01225f
C708 VDD1.n90 B 0.028954f
C709 VDD1.n91 B 0.01297f
C710 VDD1.n92 B 0.022796f
C711 VDD1.n93 B 0.01225f
C712 VDD1.n94 B 0.028954f
C713 VDD1.n95 B 0.01297f
C714 VDD1.n96 B 0.022796f
C715 VDD1.n97 B 0.01225f
C716 VDD1.n98 B 0.028954f
C717 VDD1.n99 B 0.01297f
C718 VDD1.n100 B 0.022796f
C719 VDD1.n101 B 0.01225f
C720 VDD1.n102 B 0.028954f
C721 VDD1.n103 B 0.01297f
C722 VDD1.n104 B 0.022796f
C723 VDD1.n105 B 0.01225f
C724 VDD1.n106 B 0.028954f
C725 VDD1.n107 B 0.01297f
C726 VDD1.n108 B 0.147883f
C727 VDD1.t2 B 0.047731f
C728 VDD1.n109 B 0.021716f
C729 VDD1.n110 B 0.017104f
C730 VDD1.n111 B 0.01225f
C731 VDD1.n112 B 1.46855f
C732 VDD1.n113 B 0.022796f
C733 VDD1.n114 B 0.01225f
C734 VDD1.n115 B 0.01297f
C735 VDD1.n116 B 0.028954f
C736 VDD1.n117 B 0.028954f
C737 VDD1.n118 B 0.01297f
C738 VDD1.n119 B 0.01225f
C739 VDD1.n120 B 0.022796f
C740 VDD1.n121 B 0.022796f
C741 VDD1.n122 B 0.01225f
C742 VDD1.n123 B 0.01297f
C743 VDD1.n124 B 0.028954f
C744 VDD1.n125 B 0.028954f
C745 VDD1.n126 B 0.01297f
C746 VDD1.n127 B 0.01225f
C747 VDD1.n128 B 0.022796f
C748 VDD1.n129 B 0.022796f
C749 VDD1.n130 B 0.01225f
C750 VDD1.n131 B 0.01297f
C751 VDD1.n132 B 0.028954f
C752 VDD1.n133 B 0.028954f
C753 VDD1.n134 B 0.01297f
C754 VDD1.n135 B 0.01225f
C755 VDD1.n136 B 0.022796f
C756 VDD1.n137 B 0.022796f
C757 VDD1.n138 B 0.01225f
C758 VDD1.n139 B 0.01297f
C759 VDD1.n140 B 0.028954f
C760 VDD1.n141 B 0.028954f
C761 VDD1.n142 B 0.01297f
C762 VDD1.n143 B 0.01225f
C763 VDD1.n144 B 0.022796f
C764 VDD1.n145 B 0.022796f
C765 VDD1.n146 B 0.01225f
C766 VDD1.n147 B 0.01297f
C767 VDD1.n148 B 0.028954f
C768 VDD1.n149 B 0.028954f
C769 VDD1.n150 B 0.028954f
C770 VDD1.n151 B 0.01297f
C771 VDD1.n152 B 0.01225f
C772 VDD1.n153 B 0.022796f
C773 VDD1.n154 B 0.022796f
C774 VDD1.n155 B 0.01225f
C775 VDD1.n156 B 0.01261f
C776 VDD1.n157 B 0.01261f
C777 VDD1.n158 B 0.028954f
C778 VDD1.n159 B 0.063225f
C779 VDD1.n160 B 0.01297f
C780 VDD1.n161 B 0.01225f
C781 VDD1.n162 B 0.059544f
C782 VDD1.n163 B 0.055458f
C783 VDD1.t8 B 0.267695f
C784 VDD1.t4 B 0.267695f
C785 VDD1.n164 B 2.42262f
C786 VDD1.n165 B 0.464673f
C787 VDD1.t1 B 0.267695f
C788 VDD1.t7 B 0.267695f
C789 VDD1.n166 B 2.4285f
C790 VDD1.n167 B 2.29737f
C791 VDD1.t0 B 0.267695f
C792 VDD1.t5 B 0.267695f
C793 VDD1.n168 B 2.42262f
C794 VDD1.n169 B 2.62026f
C795 VP.n0 B 0.042194f
C796 VP.t0 B 1.75074f
C797 VP.n1 B 0.625921f
C798 VP.n2 B 0.031621f
C799 VP.t9 B 1.75074f
C800 VP.n3 B 0.655611f
C801 VP.n4 B 0.031621f
C802 VP.t3 B 1.75074f
C803 VP.n5 B 0.625921f
C804 VP.n6 B 0.042194f
C805 VP.n7 B 0.042194f
C806 VP.t8 B 1.81623f
C807 VP.t1 B 1.75074f
C808 VP.n8 B 0.625921f
C809 VP.n9 B 0.031621f
C810 VP.t2 B 1.75074f
C811 VP.n10 B 0.655611f
C812 VP.n11 B 0.031621f
C813 VP.t4 B 1.75074f
C814 VP.n12 B 0.665957f
C815 VP.t7 B 1.85838f
C816 VP.n13 B 0.684935f
C817 VP.n14 B 0.168666f
C818 VP.n15 B 0.041744f
C819 VP.n16 B 0.036761f
C820 VP.n17 B 0.054118f
C821 VP.n18 B 0.031621f
C822 VP.n19 B 0.031621f
C823 VP.n20 B 0.031621f
C824 VP.n21 B 0.054118f
C825 VP.n22 B 0.036761f
C826 VP.n23 B 0.041744f
C827 VP.n24 B 0.031621f
C828 VP.n25 B 0.031621f
C829 VP.n26 B 0.052344f
C830 VP.n27 B 0.018899f
C831 VP.n28 B 0.694352f
C832 VP.n29 B 1.666f
C833 VP.n30 B 1.68938f
C834 VP.t5 B 1.81623f
C835 VP.n31 B 0.694352f
C836 VP.n32 B 0.018899f
C837 VP.n33 B 0.052344f
C838 VP.n34 B 0.031621f
C839 VP.n35 B 0.031621f
C840 VP.n36 B 0.041744f
C841 VP.n37 B 0.036761f
C842 VP.n38 B 0.054118f
C843 VP.n39 B 0.031621f
C844 VP.n40 B 0.031621f
C845 VP.n41 B 0.031621f
C846 VP.n42 B 0.054118f
C847 VP.n43 B 0.036761f
C848 VP.n44 B 0.041744f
C849 VP.n45 B 0.031621f
C850 VP.n46 B 0.031621f
C851 VP.n47 B 0.052344f
C852 VP.n48 B 0.018899f
C853 VP.t6 B 1.81623f
C854 VP.n49 B 0.694352f
C855 VP.n50 B 0.029614f
.ends

