* NGSPICE file created from diff_pair_sample_1137.ext - technology: sky130A

.subckt diff_pair_sample_1137 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=1.92
X1 VDD2.t4 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=1.92
X2 VTAIL.t5 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=1.92
X3 VTAIL.t10 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=1.92
X4 VDD2.t2 VN.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=1.92
X5 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=1.92
X6 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=1.92
X7 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=1.92
X8 VDD1.t3 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=1.92
X9 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=1.92
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=1.92
X11 VDD2.t1 VN.t4 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=1.92
X12 VTAIL.t7 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=1.92
X13 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=1.92
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=1.92
X15 VTAIL.t0 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=1.92
R0 VN.n21 VN.n12 161.3
R1 VN.n20 VN.n19 161.3
R2 VN.n18 VN.n13 161.3
R3 VN.n17 VN.n16 161.3
R4 VN.n9 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n11 VN.n10 86.3164
R9 VN.n23 VN.n22 86.3164
R10 VN.n3 VN.n2 58.0791
R11 VN.n15 VN.n14 58.0791
R12 VN.n8 VN.n1 52.6866
R13 VN.n20 VN.n13 52.6866
R14 VN.n2 VN.t3 40.2861
R15 VN.n14 VN.t4 40.2861
R16 VN VN.n23 37.805
R17 VN.n9 VN.n8 28.4674
R18 VN.n21 VN.n20 28.4674
R19 VN.n4 VN.n1 24.5923
R20 VN.n10 VN.n9 24.5923
R21 VN.n16 VN.n13 24.5923
R22 VN.n22 VN.n21 24.5923
R23 VN.n17 VN.n14 12.6034
R24 VN.n5 VN.n2 12.6034
R25 VN.n4 VN.n3 12.2964
R26 VN.n16 VN.n15 12.2964
R27 VN.n10 VN.t1 8.78696
R28 VN.n3 VN.t5 8.78696
R29 VN.n22 VN.t0 8.78696
R30 VN.n15 VN.t2 8.78696
R31 VN.n23 VN.n12 0.278335
R32 VN.n11 VN.n0 0.278335
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153485
R40 VTAIL.n11 VTAIL.t6 247.411
R41 VTAIL.n2 VTAIL.t3 247.411
R42 VTAIL.n10 VTAIL.t1 247.411
R43 VTAIL.n7 VTAIL.t9 247.411
R44 VTAIL.n1 VTAIL.n0 219.125
R45 VTAIL.n4 VTAIL.n3 219.125
R46 VTAIL.n9 VTAIL.n8 219.125
R47 VTAIL.n6 VTAIL.n5 219.125
R48 VTAIL.n0 VTAIL.t8 28.2862
R49 VTAIL.n0 VTAIL.t7 28.2862
R50 VTAIL.n3 VTAIL.t2 28.2862
R51 VTAIL.n3 VTAIL.t0 28.2862
R52 VTAIL.n8 VTAIL.t4 28.2862
R53 VTAIL.n8 VTAIL.t5 28.2862
R54 VTAIL.n5 VTAIL.t11 28.2862
R55 VTAIL.n5 VTAIL.t10 28.2862
R56 VTAIL.n6 VTAIL.n4 16.8496
R57 VTAIL.n11 VTAIL.n10 14.91
R58 VTAIL.n7 VTAIL.n6 1.94016
R59 VTAIL.n10 VTAIL.n9 1.94016
R60 VTAIL.n4 VTAIL.n2 1.94016
R61 VTAIL.n9 VTAIL.n7 1.44016
R62 VTAIL.n2 VTAIL.n1 1.44016
R63 VTAIL VTAIL.n11 1.39705
R64 VTAIL VTAIL.n1 0.543603
R65 VDD2.n1 VDD2.t2 265.488
R66 VDD2.n2 VDD2.t5 264.089
R67 VDD2.n1 VDD2.n0 236.233
R68 VDD2 VDD2.n3 236.231
R69 VDD2.n2 VDD2.n1 30.6226
R70 VDD2.n3 VDD2.t3 28.2862
R71 VDD2.n3 VDD2.t1 28.2862
R72 VDD2.n0 VDD2.t0 28.2862
R73 VDD2.n0 VDD2.t4 28.2862
R74 VDD2 VDD2.n2 1.51343
R75 B.n368 B.n367 585
R76 B.n370 B.n83 585
R77 B.n373 B.n372 585
R78 B.n374 B.n82 585
R79 B.n376 B.n375 585
R80 B.n378 B.n81 585
R81 B.n380 B.n379 585
R82 B.n382 B.n381 585
R83 B.n385 B.n384 585
R84 B.n386 B.n76 585
R85 B.n388 B.n387 585
R86 B.n390 B.n75 585
R87 B.n393 B.n392 585
R88 B.n394 B.n74 585
R89 B.n396 B.n395 585
R90 B.n398 B.n73 585
R91 B.n401 B.n400 585
R92 B.n402 B.n70 585
R93 B.n405 B.n404 585
R94 B.n407 B.n69 585
R95 B.n410 B.n409 585
R96 B.n411 B.n68 585
R97 B.n413 B.n412 585
R98 B.n415 B.n67 585
R99 B.n418 B.n417 585
R100 B.n419 B.n66 585
R101 B.n366 B.n64 585
R102 B.n422 B.n64 585
R103 B.n365 B.n63 585
R104 B.n423 B.n63 585
R105 B.n364 B.n62 585
R106 B.n424 B.n62 585
R107 B.n363 B.n362 585
R108 B.n362 B.n58 585
R109 B.n361 B.n57 585
R110 B.n430 B.n57 585
R111 B.n360 B.n56 585
R112 B.n431 B.n56 585
R113 B.n359 B.n55 585
R114 B.n432 B.n55 585
R115 B.n358 B.n357 585
R116 B.n357 B.n51 585
R117 B.n356 B.n50 585
R118 B.n438 B.n50 585
R119 B.n355 B.n49 585
R120 B.n439 B.n49 585
R121 B.n354 B.n48 585
R122 B.n440 B.n48 585
R123 B.n353 B.n352 585
R124 B.n352 B.n44 585
R125 B.n351 B.n43 585
R126 B.n446 B.n43 585
R127 B.n350 B.n42 585
R128 B.n447 B.n42 585
R129 B.n349 B.n41 585
R130 B.n448 B.n41 585
R131 B.n348 B.n347 585
R132 B.n347 B.n37 585
R133 B.n346 B.n36 585
R134 B.n454 B.n36 585
R135 B.n345 B.n35 585
R136 B.n455 B.n35 585
R137 B.n344 B.n34 585
R138 B.n456 B.n34 585
R139 B.n343 B.n342 585
R140 B.n342 B.n30 585
R141 B.n341 B.n29 585
R142 B.n462 B.n29 585
R143 B.n340 B.n28 585
R144 B.n463 B.n28 585
R145 B.n339 B.n27 585
R146 B.n464 B.n27 585
R147 B.n338 B.n337 585
R148 B.n337 B.n23 585
R149 B.n336 B.n22 585
R150 B.n470 B.n22 585
R151 B.n335 B.n21 585
R152 B.n471 B.n21 585
R153 B.n334 B.n20 585
R154 B.n472 B.n20 585
R155 B.n333 B.n332 585
R156 B.n332 B.n16 585
R157 B.n331 B.n15 585
R158 B.n478 B.n15 585
R159 B.n330 B.n14 585
R160 B.n479 B.n14 585
R161 B.n329 B.n13 585
R162 B.n480 B.n13 585
R163 B.n328 B.n327 585
R164 B.n327 B.n12 585
R165 B.n326 B.n325 585
R166 B.n326 B.n8 585
R167 B.n324 B.n7 585
R168 B.n487 B.n7 585
R169 B.n323 B.n6 585
R170 B.n488 B.n6 585
R171 B.n322 B.n5 585
R172 B.n489 B.n5 585
R173 B.n321 B.n320 585
R174 B.n320 B.n4 585
R175 B.n319 B.n84 585
R176 B.n319 B.n318 585
R177 B.n309 B.n85 585
R178 B.n86 B.n85 585
R179 B.n311 B.n310 585
R180 B.n312 B.n311 585
R181 B.n308 B.n90 585
R182 B.n94 B.n90 585
R183 B.n307 B.n306 585
R184 B.n306 B.n305 585
R185 B.n92 B.n91 585
R186 B.n93 B.n92 585
R187 B.n298 B.n297 585
R188 B.n299 B.n298 585
R189 B.n296 B.n99 585
R190 B.n99 B.n98 585
R191 B.n295 B.n294 585
R192 B.n294 B.n293 585
R193 B.n101 B.n100 585
R194 B.n102 B.n101 585
R195 B.n286 B.n285 585
R196 B.n287 B.n286 585
R197 B.n284 B.n107 585
R198 B.n107 B.n106 585
R199 B.n283 B.n282 585
R200 B.n282 B.n281 585
R201 B.n109 B.n108 585
R202 B.n110 B.n109 585
R203 B.n274 B.n273 585
R204 B.n275 B.n274 585
R205 B.n272 B.n115 585
R206 B.n115 B.n114 585
R207 B.n271 B.n270 585
R208 B.n270 B.n269 585
R209 B.n117 B.n116 585
R210 B.n118 B.n117 585
R211 B.n262 B.n261 585
R212 B.n263 B.n262 585
R213 B.n260 B.n123 585
R214 B.n123 B.n122 585
R215 B.n259 B.n258 585
R216 B.n258 B.n257 585
R217 B.n125 B.n124 585
R218 B.n126 B.n125 585
R219 B.n250 B.n249 585
R220 B.n251 B.n250 585
R221 B.n248 B.n131 585
R222 B.n131 B.n130 585
R223 B.n247 B.n246 585
R224 B.n246 B.n245 585
R225 B.n133 B.n132 585
R226 B.n134 B.n133 585
R227 B.n238 B.n237 585
R228 B.n239 B.n238 585
R229 B.n236 B.n139 585
R230 B.n139 B.n138 585
R231 B.n235 B.n234 585
R232 B.n234 B.n233 585
R233 B.n141 B.n140 585
R234 B.n142 B.n141 585
R235 B.n226 B.n225 585
R236 B.n227 B.n226 585
R237 B.n224 B.n147 585
R238 B.n147 B.n146 585
R239 B.n223 B.n222 585
R240 B.n222 B.n221 585
R241 B.n218 B.n151 585
R242 B.n217 B.n216 585
R243 B.n214 B.n152 585
R244 B.n214 B.n150 585
R245 B.n213 B.n212 585
R246 B.n211 B.n210 585
R247 B.n209 B.n154 585
R248 B.n207 B.n206 585
R249 B.n205 B.n155 585
R250 B.n203 B.n202 585
R251 B.n200 B.n158 585
R252 B.n198 B.n197 585
R253 B.n196 B.n159 585
R254 B.n195 B.n194 585
R255 B.n192 B.n160 585
R256 B.n190 B.n189 585
R257 B.n188 B.n161 585
R258 B.n187 B.n186 585
R259 B.n184 B.n162 585
R260 B.n182 B.n181 585
R261 B.n180 B.n163 585
R262 B.n179 B.n178 585
R263 B.n176 B.n167 585
R264 B.n174 B.n173 585
R265 B.n172 B.n168 585
R266 B.n171 B.n170 585
R267 B.n149 B.n148 585
R268 B.n150 B.n149 585
R269 B.n220 B.n219 585
R270 B.n221 B.n220 585
R271 B.n145 B.n144 585
R272 B.n146 B.n145 585
R273 B.n229 B.n228 585
R274 B.n228 B.n227 585
R275 B.n230 B.n143 585
R276 B.n143 B.n142 585
R277 B.n232 B.n231 585
R278 B.n233 B.n232 585
R279 B.n137 B.n136 585
R280 B.n138 B.n137 585
R281 B.n241 B.n240 585
R282 B.n240 B.n239 585
R283 B.n242 B.n135 585
R284 B.n135 B.n134 585
R285 B.n244 B.n243 585
R286 B.n245 B.n244 585
R287 B.n129 B.n128 585
R288 B.n130 B.n129 585
R289 B.n253 B.n252 585
R290 B.n252 B.n251 585
R291 B.n254 B.n127 585
R292 B.n127 B.n126 585
R293 B.n256 B.n255 585
R294 B.n257 B.n256 585
R295 B.n121 B.n120 585
R296 B.n122 B.n121 585
R297 B.n265 B.n264 585
R298 B.n264 B.n263 585
R299 B.n266 B.n119 585
R300 B.n119 B.n118 585
R301 B.n268 B.n267 585
R302 B.n269 B.n268 585
R303 B.n113 B.n112 585
R304 B.n114 B.n113 585
R305 B.n277 B.n276 585
R306 B.n276 B.n275 585
R307 B.n278 B.n111 585
R308 B.n111 B.n110 585
R309 B.n280 B.n279 585
R310 B.n281 B.n280 585
R311 B.n105 B.n104 585
R312 B.n106 B.n105 585
R313 B.n289 B.n288 585
R314 B.n288 B.n287 585
R315 B.n290 B.n103 585
R316 B.n103 B.n102 585
R317 B.n292 B.n291 585
R318 B.n293 B.n292 585
R319 B.n97 B.n96 585
R320 B.n98 B.n97 585
R321 B.n301 B.n300 585
R322 B.n300 B.n299 585
R323 B.n302 B.n95 585
R324 B.n95 B.n93 585
R325 B.n304 B.n303 585
R326 B.n305 B.n304 585
R327 B.n89 B.n88 585
R328 B.n94 B.n89 585
R329 B.n314 B.n313 585
R330 B.n313 B.n312 585
R331 B.n315 B.n87 585
R332 B.n87 B.n86 585
R333 B.n317 B.n316 585
R334 B.n318 B.n317 585
R335 B.n3 B.n0 585
R336 B.n4 B.n3 585
R337 B.n486 B.n1 585
R338 B.n487 B.n486 585
R339 B.n485 B.n484 585
R340 B.n485 B.n8 585
R341 B.n483 B.n9 585
R342 B.n12 B.n9 585
R343 B.n482 B.n481 585
R344 B.n481 B.n480 585
R345 B.n11 B.n10 585
R346 B.n479 B.n11 585
R347 B.n477 B.n476 585
R348 B.n478 B.n477 585
R349 B.n475 B.n17 585
R350 B.n17 B.n16 585
R351 B.n474 B.n473 585
R352 B.n473 B.n472 585
R353 B.n19 B.n18 585
R354 B.n471 B.n19 585
R355 B.n469 B.n468 585
R356 B.n470 B.n469 585
R357 B.n467 B.n24 585
R358 B.n24 B.n23 585
R359 B.n466 B.n465 585
R360 B.n465 B.n464 585
R361 B.n26 B.n25 585
R362 B.n463 B.n26 585
R363 B.n461 B.n460 585
R364 B.n462 B.n461 585
R365 B.n459 B.n31 585
R366 B.n31 B.n30 585
R367 B.n458 B.n457 585
R368 B.n457 B.n456 585
R369 B.n33 B.n32 585
R370 B.n455 B.n33 585
R371 B.n453 B.n452 585
R372 B.n454 B.n453 585
R373 B.n451 B.n38 585
R374 B.n38 B.n37 585
R375 B.n450 B.n449 585
R376 B.n449 B.n448 585
R377 B.n40 B.n39 585
R378 B.n447 B.n40 585
R379 B.n445 B.n444 585
R380 B.n446 B.n445 585
R381 B.n443 B.n45 585
R382 B.n45 B.n44 585
R383 B.n442 B.n441 585
R384 B.n441 B.n440 585
R385 B.n47 B.n46 585
R386 B.n439 B.n47 585
R387 B.n437 B.n436 585
R388 B.n438 B.n437 585
R389 B.n435 B.n52 585
R390 B.n52 B.n51 585
R391 B.n434 B.n433 585
R392 B.n433 B.n432 585
R393 B.n54 B.n53 585
R394 B.n431 B.n54 585
R395 B.n429 B.n428 585
R396 B.n430 B.n429 585
R397 B.n427 B.n59 585
R398 B.n59 B.n58 585
R399 B.n426 B.n425 585
R400 B.n425 B.n424 585
R401 B.n61 B.n60 585
R402 B.n423 B.n61 585
R403 B.n421 B.n420 585
R404 B.n422 B.n421 585
R405 B.n490 B.n489 585
R406 B.n488 B.n2 585
R407 B.n421 B.n66 540.549
R408 B.n368 B.n64 540.549
R409 B.n222 B.n149 540.549
R410 B.n220 B.n151 540.549
R411 B.n71 B.t12 280.195
R412 B.n77 B.t15 280.195
R413 B.n164 B.t9 280.195
R414 B.n156 B.t19 280.195
R415 B.n369 B.n65 256.663
R416 B.n371 B.n65 256.663
R417 B.n377 B.n65 256.663
R418 B.n80 B.n65 256.663
R419 B.n383 B.n65 256.663
R420 B.n389 B.n65 256.663
R421 B.n391 B.n65 256.663
R422 B.n397 B.n65 256.663
R423 B.n399 B.n65 256.663
R424 B.n406 B.n65 256.663
R425 B.n408 B.n65 256.663
R426 B.n414 B.n65 256.663
R427 B.n416 B.n65 256.663
R428 B.n215 B.n150 256.663
R429 B.n153 B.n150 256.663
R430 B.n208 B.n150 256.663
R431 B.n201 B.n150 256.663
R432 B.n199 B.n150 256.663
R433 B.n193 B.n150 256.663
R434 B.n191 B.n150 256.663
R435 B.n185 B.n150 256.663
R436 B.n183 B.n150 256.663
R437 B.n177 B.n150 256.663
R438 B.n175 B.n150 256.663
R439 B.n169 B.n150 256.663
R440 B.n492 B.n491 256.663
R441 B.n221 B.n150 237.49
R442 B.n422 B.n65 237.49
R443 B.n72 B.t13 236.559
R444 B.n78 B.t16 236.559
R445 B.n165 B.t8 236.559
R446 B.n157 B.t18 236.559
R447 B.n71 B.t10 208.226
R448 B.n77 B.t14 208.226
R449 B.n164 B.t6 208.226
R450 B.n156 B.t17 208.226
R451 B.n417 B.n415 163.367
R452 B.n413 B.n68 163.367
R453 B.n409 B.n407 163.367
R454 B.n405 B.n70 163.367
R455 B.n400 B.n398 163.367
R456 B.n396 B.n74 163.367
R457 B.n392 B.n390 163.367
R458 B.n388 B.n76 163.367
R459 B.n384 B.n382 163.367
R460 B.n379 B.n378 163.367
R461 B.n376 B.n82 163.367
R462 B.n372 B.n370 163.367
R463 B.n222 B.n147 163.367
R464 B.n226 B.n147 163.367
R465 B.n226 B.n141 163.367
R466 B.n234 B.n141 163.367
R467 B.n234 B.n139 163.367
R468 B.n238 B.n139 163.367
R469 B.n238 B.n133 163.367
R470 B.n246 B.n133 163.367
R471 B.n246 B.n131 163.367
R472 B.n250 B.n131 163.367
R473 B.n250 B.n125 163.367
R474 B.n258 B.n125 163.367
R475 B.n258 B.n123 163.367
R476 B.n262 B.n123 163.367
R477 B.n262 B.n117 163.367
R478 B.n270 B.n117 163.367
R479 B.n270 B.n115 163.367
R480 B.n274 B.n115 163.367
R481 B.n274 B.n109 163.367
R482 B.n282 B.n109 163.367
R483 B.n282 B.n107 163.367
R484 B.n286 B.n107 163.367
R485 B.n286 B.n101 163.367
R486 B.n294 B.n101 163.367
R487 B.n294 B.n99 163.367
R488 B.n298 B.n99 163.367
R489 B.n298 B.n92 163.367
R490 B.n306 B.n92 163.367
R491 B.n306 B.n90 163.367
R492 B.n311 B.n90 163.367
R493 B.n311 B.n85 163.367
R494 B.n319 B.n85 163.367
R495 B.n320 B.n319 163.367
R496 B.n320 B.n5 163.367
R497 B.n6 B.n5 163.367
R498 B.n7 B.n6 163.367
R499 B.n326 B.n7 163.367
R500 B.n327 B.n326 163.367
R501 B.n327 B.n13 163.367
R502 B.n14 B.n13 163.367
R503 B.n15 B.n14 163.367
R504 B.n332 B.n15 163.367
R505 B.n332 B.n20 163.367
R506 B.n21 B.n20 163.367
R507 B.n22 B.n21 163.367
R508 B.n337 B.n22 163.367
R509 B.n337 B.n27 163.367
R510 B.n28 B.n27 163.367
R511 B.n29 B.n28 163.367
R512 B.n342 B.n29 163.367
R513 B.n342 B.n34 163.367
R514 B.n35 B.n34 163.367
R515 B.n36 B.n35 163.367
R516 B.n347 B.n36 163.367
R517 B.n347 B.n41 163.367
R518 B.n42 B.n41 163.367
R519 B.n43 B.n42 163.367
R520 B.n352 B.n43 163.367
R521 B.n352 B.n48 163.367
R522 B.n49 B.n48 163.367
R523 B.n50 B.n49 163.367
R524 B.n357 B.n50 163.367
R525 B.n357 B.n55 163.367
R526 B.n56 B.n55 163.367
R527 B.n57 B.n56 163.367
R528 B.n362 B.n57 163.367
R529 B.n362 B.n62 163.367
R530 B.n63 B.n62 163.367
R531 B.n64 B.n63 163.367
R532 B.n216 B.n214 163.367
R533 B.n214 B.n213 163.367
R534 B.n210 B.n209 163.367
R535 B.n207 B.n155 163.367
R536 B.n202 B.n200 163.367
R537 B.n198 B.n159 163.367
R538 B.n194 B.n192 163.367
R539 B.n190 B.n161 163.367
R540 B.n186 B.n184 163.367
R541 B.n182 B.n163 163.367
R542 B.n178 B.n176 163.367
R543 B.n174 B.n168 163.367
R544 B.n170 B.n149 163.367
R545 B.n220 B.n145 163.367
R546 B.n228 B.n145 163.367
R547 B.n228 B.n143 163.367
R548 B.n232 B.n143 163.367
R549 B.n232 B.n137 163.367
R550 B.n240 B.n137 163.367
R551 B.n240 B.n135 163.367
R552 B.n244 B.n135 163.367
R553 B.n244 B.n129 163.367
R554 B.n252 B.n129 163.367
R555 B.n252 B.n127 163.367
R556 B.n256 B.n127 163.367
R557 B.n256 B.n121 163.367
R558 B.n264 B.n121 163.367
R559 B.n264 B.n119 163.367
R560 B.n268 B.n119 163.367
R561 B.n268 B.n113 163.367
R562 B.n276 B.n113 163.367
R563 B.n276 B.n111 163.367
R564 B.n280 B.n111 163.367
R565 B.n280 B.n105 163.367
R566 B.n288 B.n105 163.367
R567 B.n288 B.n103 163.367
R568 B.n292 B.n103 163.367
R569 B.n292 B.n97 163.367
R570 B.n300 B.n97 163.367
R571 B.n300 B.n95 163.367
R572 B.n304 B.n95 163.367
R573 B.n304 B.n89 163.367
R574 B.n313 B.n89 163.367
R575 B.n313 B.n87 163.367
R576 B.n317 B.n87 163.367
R577 B.n317 B.n3 163.367
R578 B.n490 B.n3 163.367
R579 B.n486 B.n2 163.367
R580 B.n486 B.n485 163.367
R581 B.n485 B.n9 163.367
R582 B.n481 B.n9 163.367
R583 B.n481 B.n11 163.367
R584 B.n477 B.n11 163.367
R585 B.n477 B.n17 163.367
R586 B.n473 B.n17 163.367
R587 B.n473 B.n19 163.367
R588 B.n469 B.n19 163.367
R589 B.n469 B.n24 163.367
R590 B.n465 B.n24 163.367
R591 B.n465 B.n26 163.367
R592 B.n461 B.n26 163.367
R593 B.n461 B.n31 163.367
R594 B.n457 B.n31 163.367
R595 B.n457 B.n33 163.367
R596 B.n453 B.n33 163.367
R597 B.n453 B.n38 163.367
R598 B.n449 B.n38 163.367
R599 B.n449 B.n40 163.367
R600 B.n445 B.n40 163.367
R601 B.n445 B.n45 163.367
R602 B.n441 B.n45 163.367
R603 B.n441 B.n47 163.367
R604 B.n437 B.n47 163.367
R605 B.n437 B.n52 163.367
R606 B.n433 B.n52 163.367
R607 B.n433 B.n54 163.367
R608 B.n429 B.n54 163.367
R609 B.n429 B.n59 163.367
R610 B.n425 B.n59 163.367
R611 B.n425 B.n61 163.367
R612 B.n421 B.n61 163.367
R613 B.n221 B.n146 125.189
R614 B.n227 B.n146 125.189
R615 B.n227 B.n142 125.189
R616 B.n233 B.n142 125.189
R617 B.n233 B.n138 125.189
R618 B.n239 B.n138 125.189
R619 B.n245 B.n134 125.189
R620 B.n245 B.n130 125.189
R621 B.n251 B.n130 125.189
R622 B.n251 B.n126 125.189
R623 B.n257 B.n126 125.189
R624 B.n257 B.n122 125.189
R625 B.n263 B.n122 125.189
R626 B.n263 B.n118 125.189
R627 B.n269 B.n118 125.189
R628 B.n275 B.n114 125.189
R629 B.n275 B.n110 125.189
R630 B.n281 B.n110 125.189
R631 B.n281 B.n106 125.189
R632 B.n287 B.n106 125.189
R633 B.n293 B.n102 125.189
R634 B.n293 B.n98 125.189
R635 B.n299 B.n98 125.189
R636 B.n299 B.n93 125.189
R637 B.n305 B.n93 125.189
R638 B.n305 B.n94 125.189
R639 B.n312 B.n86 125.189
R640 B.n318 B.n86 125.189
R641 B.n318 B.n4 125.189
R642 B.n489 B.n4 125.189
R643 B.n489 B.n488 125.189
R644 B.n488 B.n487 125.189
R645 B.n487 B.n8 125.189
R646 B.n12 B.n8 125.189
R647 B.n480 B.n12 125.189
R648 B.n479 B.n478 125.189
R649 B.n478 B.n16 125.189
R650 B.n472 B.n16 125.189
R651 B.n472 B.n471 125.189
R652 B.n471 B.n470 125.189
R653 B.n470 B.n23 125.189
R654 B.n464 B.n463 125.189
R655 B.n463 B.n462 125.189
R656 B.n462 B.n30 125.189
R657 B.n456 B.n30 125.189
R658 B.n456 B.n455 125.189
R659 B.n454 B.n37 125.189
R660 B.n448 B.n37 125.189
R661 B.n448 B.n447 125.189
R662 B.n447 B.n446 125.189
R663 B.n446 B.n44 125.189
R664 B.n440 B.n44 125.189
R665 B.n440 B.n439 125.189
R666 B.n439 B.n438 125.189
R667 B.n438 B.n51 125.189
R668 B.n432 B.n431 125.189
R669 B.n431 B.n430 125.189
R670 B.n430 B.n58 125.189
R671 B.n424 B.n58 125.189
R672 B.n424 B.n423 125.189
R673 B.n423 B.n422 125.189
R674 B.n287 B.t0 121.507
R675 B.n464 B.t5 121.507
R676 B.t2 B.n114 81.0047
R677 B.n455 B.t1 81.0047
R678 B.n94 B.t3 73.6407
R679 B.t4 B.n479 73.6407
R680 B.n416 B.n66 71.676
R681 B.n415 B.n414 71.676
R682 B.n408 B.n68 71.676
R683 B.n407 B.n406 71.676
R684 B.n399 B.n70 71.676
R685 B.n398 B.n397 71.676
R686 B.n391 B.n74 71.676
R687 B.n390 B.n389 71.676
R688 B.n383 B.n76 71.676
R689 B.n382 B.n80 71.676
R690 B.n378 B.n377 71.676
R691 B.n371 B.n82 71.676
R692 B.n370 B.n369 71.676
R693 B.n369 B.n368 71.676
R694 B.n372 B.n371 71.676
R695 B.n377 B.n376 71.676
R696 B.n379 B.n80 71.676
R697 B.n384 B.n383 71.676
R698 B.n389 B.n388 71.676
R699 B.n392 B.n391 71.676
R700 B.n397 B.n396 71.676
R701 B.n400 B.n399 71.676
R702 B.n406 B.n405 71.676
R703 B.n409 B.n408 71.676
R704 B.n414 B.n413 71.676
R705 B.n417 B.n416 71.676
R706 B.n215 B.n151 71.676
R707 B.n213 B.n153 71.676
R708 B.n209 B.n208 71.676
R709 B.n201 B.n155 71.676
R710 B.n200 B.n199 71.676
R711 B.n193 B.n159 71.676
R712 B.n192 B.n191 71.676
R713 B.n185 B.n161 71.676
R714 B.n184 B.n183 71.676
R715 B.n177 B.n163 71.676
R716 B.n176 B.n175 71.676
R717 B.n169 B.n168 71.676
R718 B.n216 B.n215 71.676
R719 B.n210 B.n153 71.676
R720 B.n208 B.n207 71.676
R721 B.n202 B.n201 71.676
R722 B.n199 B.n198 71.676
R723 B.n194 B.n193 71.676
R724 B.n191 B.n190 71.676
R725 B.n186 B.n185 71.676
R726 B.n183 B.n182 71.676
R727 B.n178 B.n177 71.676
R728 B.n175 B.n174 71.676
R729 B.n170 B.n169 71.676
R730 B.n491 B.n490 71.676
R731 B.n491 B.n2 71.676
R732 B.n239 B.t7 66.2766
R733 B.n432 B.t11 66.2766
R734 B.n403 B.n72 59.5399
R735 B.n79 B.n78 59.5399
R736 B.n166 B.n165 59.5399
R737 B.n204 B.n157 59.5399
R738 B.t7 B.n134 58.9126
R739 B.t11 B.n51 58.9126
R740 B.n312 B.t3 51.5486
R741 B.n480 B.t4 51.5486
R742 B.n269 B.t2 44.1846
R743 B.t1 B.n454 44.1846
R744 B.n72 B.n71 43.6369
R745 B.n78 B.n77 43.6369
R746 B.n165 B.n164 43.6369
R747 B.n157 B.n156 43.6369
R748 B.n219 B.n218 35.1225
R749 B.n223 B.n148 35.1225
R750 B.n420 B.n419 35.1225
R751 B.n367 B.n366 35.1224
R752 B B.n492 18.0485
R753 B.n219 B.n144 10.6151
R754 B.n229 B.n144 10.6151
R755 B.n230 B.n229 10.6151
R756 B.n231 B.n230 10.6151
R757 B.n231 B.n136 10.6151
R758 B.n241 B.n136 10.6151
R759 B.n242 B.n241 10.6151
R760 B.n243 B.n242 10.6151
R761 B.n243 B.n128 10.6151
R762 B.n253 B.n128 10.6151
R763 B.n254 B.n253 10.6151
R764 B.n255 B.n254 10.6151
R765 B.n255 B.n120 10.6151
R766 B.n265 B.n120 10.6151
R767 B.n266 B.n265 10.6151
R768 B.n267 B.n266 10.6151
R769 B.n267 B.n112 10.6151
R770 B.n277 B.n112 10.6151
R771 B.n278 B.n277 10.6151
R772 B.n279 B.n278 10.6151
R773 B.n279 B.n104 10.6151
R774 B.n289 B.n104 10.6151
R775 B.n290 B.n289 10.6151
R776 B.n291 B.n290 10.6151
R777 B.n291 B.n96 10.6151
R778 B.n301 B.n96 10.6151
R779 B.n302 B.n301 10.6151
R780 B.n303 B.n302 10.6151
R781 B.n303 B.n88 10.6151
R782 B.n314 B.n88 10.6151
R783 B.n315 B.n314 10.6151
R784 B.n316 B.n315 10.6151
R785 B.n316 B.n0 10.6151
R786 B.n218 B.n217 10.6151
R787 B.n217 B.n152 10.6151
R788 B.n212 B.n152 10.6151
R789 B.n212 B.n211 10.6151
R790 B.n211 B.n154 10.6151
R791 B.n206 B.n154 10.6151
R792 B.n206 B.n205 10.6151
R793 B.n203 B.n158 10.6151
R794 B.n197 B.n158 10.6151
R795 B.n197 B.n196 10.6151
R796 B.n196 B.n195 10.6151
R797 B.n195 B.n160 10.6151
R798 B.n189 B.n160 10.6151
R799 B.n189 B.n188 10.6151
R800 B.n188 B.n187 10.6151
R801 B.n187 B.n162 10.6151
R802 B.n181 B.n180 10.6151
R803 B.n180 B.n179 10.6151
R804 B.n179 B.n167 10.6151
R805 B.n173 B.n167 10.6151
R806 B.n173 B.n172 10.6151
R807 B.n172 B.n171 10.6151
R808 B.n171 B.n148 10.6151
R809 B.n224 B.n223 10.6151
R810 B.n225 B.n224 10.6151
R811 B.n225 B.n140 10.6151
R812 B.n235 B.n140 10.6151
R813 B.n236 B.n235 10.6151
R814 B.n237 B.n236 10.6151
R815 B.n237 B.n132 10.6151
R816 B.n247 B.n132 10.6151
R817 B.n248 B.n247 10.6151
R818 B.n249 B.n248 10.6151
R819 B.n249 B.n124 10.6151
R820 B.n259 B.n124 10.6151
R821 B.n260 B.n259 10.6151
R822 B.n261 B.n260 10.6151
R823 B.n261 B.n116 10.6151
R824 B.n271 B.n116 10.6151
R825 B.n272 B.n271 10.6151
R826 B.n273 B.n272 10.6151
R827 B.n273 B.n108 10.6151
R828 B.n283 B.n108 10.6151
R829 B.n284 B.n283 10.6151
R830 B.n285 B.n284 10.6151
R831 B.n285 B.n100 10.6151
R832 B.n295 B.n100 10.6151
R833 B.n296 B.n295 10.6151
R834 B.n297 B.n296 10.6151
R835 B.n297 B.n91 10.6151
R836 B.n307 B.n91 10.6151
R837 B.n308 B.n307 10.6151
R838 B.n310 B.n308 10.6151
R839 B.n310 B.n309 10.6151
R840 B.n309 B.n84 10.6151
R841 B.n321 B.n84 10.6151
R842 B.n322 B.n321 10.6151
R843 B.n323 B.n322 10.6151
R844 B.n324 B.n323 10.6151
R845 B.n325 B.n324 10.6151
R846 B.n328 B.n325 10.6151
R847 B.n329 B.n328 10.6151
R848 B.n330 B.n329 10.6151
R849 B.n331 B.n330 10.6151
R850 B.n333 B.n331 10.6151
R851 B.n334 B.n333 10.6151
R852 B.n335 B.n334 10.6151
R853 B.n336 B.n335 10.6151
R854 B.n338 B.n336 10.6151
R855 B.n339 B.n338 10.6151
R856 B.n340 B.n339 10.6151
R857 B.n341 B.n340 10.6151
R858 B.n343 B.n341 10.6151
R859 B.n344 B.n343 10.6151
R860 B.n345 B.n344 10.6151
R861 B.n346 B.n345 10.6151
R862 B.n348 B.n346 10.6151
R863 B.n349 B.n348 10.6151
R864 B.n350 B.n349 10.6151
R865 B.n351 B.n350 10.6151
R866 B.n353 B.n351 10.6151
R867 B.n354 B.n353 10.6151
R868 B.n355 B.n354 10.6151
R869 B.n356 B.n355 10.6151
R870 B.n358 B.n356 10.6151
R871 B.n359 B.n358 10.6151
R872 B.n360 B.n359 10.6151
R873 B.n361 B.n360 10.6151
R874 B.n363 B.n361 10.6151
R875 B.n364 B.n363 10.6151
R876 B.n365 B.n364 10.6151
R877 B.n366 B.n365 10.6151
R878 B.n484 B.n1 10.6151
R879 B.n484 B.n483 10.6151
R880 B.n483 B.n482 10.6151
R881 B.n482 B.n10 10.6151
R882 B.n476 B.n10 10.6151
R883 B.n476 B.n475 10.6151
R884 B.n475 B.n474 10.6151
R885 B.n474 B.n18 10.6151
R886 B.n468 B.n18 10.6151
R887 B.n468 B.n467 10.6151
R888 B.n467 B.n466 10.6151
R889 B.n466 B.n25 10.6151
R890 B.n460 B.n25 10.6151
R891 B.n460 B.n459 10.6151
R892 B.n459 B.n458 10.6151
R893 B.n458 B.n32 10.6151
R894 B.n452 B.n32 10.6151
R895 B.n452 B.n451 10.6151
R896 B.n451 B.n450 10.6151
R897 B.n450 B.n39 10.6151
R898 B.n444 B.n39 10.6151
R899 B.n444 B.n443 10.6151
R900 B.n443 B.n442 10.6151
R901 B.n442 B.n46 10.6151
R902 B.n436 B.n46 10.6151
R903 B.n436 B.n435 10.6151
R904 B.n435 B.n434 10.6151
R905 B.n434 B.n53 10.6151
R906 B.n428 B.n53 10.6151
R907 B.n428 B.n427 10.6151
R908 B.n427 B.n426 10.6151
R909 B.n426 B.n60 10.6151
R910 B.n420 B.n60 10.6151
R911 B.n419 B.n418 10.6151
R912 B.n418 B.n67 10.6151
R913 B.n412 B.n67 10.6151
R914 B.n412 B.n411 10.6151
R915 B.n411 B.n410 10.6151
R916 B.n410 B.n69 10.6151
R917 B.n404 B.n69 10.6151
R918 B.n402 B.n401 10.6151
R919 B.n401 B.n73 10.6151
R920 B.n395 B.n73 10.6151
R921 B.n395 B.n394 10.6151
R922 B.n394 B.n393 10.6151
R923 B.n393 B.n75 10.6151
R924 B.n387 B.n75 10.6151
R925 B.n387 B.n386 10.6151
R926 B.n386 B.n385 10.6151
R927 B.n381 B.n380 10.6151
R928 B.n380 B.n81 10.6151
R929 B.n375 B.n81 10.6151
R930 B.n375 B.n374 10.6151
R931 B.n374 B.n373 10.6151
R932 B.n373 B.n83 10.6151
R933 B.n367 B.n83 10.6151
R934 B.n205 B.n204 9.36635
R935 B.n181 B.n166 9.36635
R936 B.n404 B.n403 9.36635
R937 B.n381 B.n79 9.36635
R938 B.n492 B.n0 8.11757
R939 B.n492 B.n1 8.11757
R940 B.t0 B.n102 3.68251
R941 B.t5 B.n23 3.68251
R942 B.n204 B.n203 1.24928
R943 B.n166 B.n162 1.24928
R944 B.n403 B.n402 1.24928
R945 B.n385 B.n79 1.24928
R946 VP.n9 VP.n8 161.3
R947 VP.n10 VP.n5 161.3
R948 VP.n12 VP.n11 161.3
R949 VP.n13 VP.n4 161.3
R950 VP.n30 VP.n0 161.3
R951 VP.n29 VP.n28 161.3
R952 VP.n27 VP.n1 161.3
R953 VP.n26 VP.n25 161.3
R954 VP.n23 VP.n2 161.3
R955 VP.n22 VP.n21 161.3
R956 VP.n20 VP.n3 161.3
R957 VP.n19 VP.n18 161.3
R958 VP.n17 VP.n16 86.3164
R959 VP.n32 VP.n31 86.3164
R960 VP.n15 VP.n14 86.3164
R961 VP.n7 VP.n6 58.0791
R962 VP.n22 VP.n3 52.6866
R963 VP.n29 VP.n1 52.6866
R964 VP.n12 VP.n5 52.6866
R965 VP.n6 VP.t3 40.2861
R966 VP.n16 VP.n15 37.5262
R967 VP.n18 VP.n3 28.4674
R968 VP.n30 VP.n29 28.4674
R969 VP.n13 VP.n12 28.4674
R970 VP.n18 VP.n17 24.5923
R971 VP.n23 VP.n22 24.5923
R972 VP.n25 VP.n1 24.5923
R973 VP.n31 VP.n30 24.5923
R974 VP.n14 VP.n13 24.5923
R975 VP.n8 VP.n5 24.5923
R976 VP.n9 VP.n6 12.6034
R977 VP.n24 VP.n23 12.2964
R978 VP.n25 VP.n24 12.2964
R979 VP.n8 VP.n7 12.2964
R980 VP.n31 VP.t2 8.78696
R981 VP.n17 VP.t1 8.78696
R982 VP.n24 VP.t5 8.78696
R983 VP.n14 VP.t4 8.78696
R984 VP.n7 VP.t0 8.78696
R985 VP.n15 VP.n4 0.278335
R986 VP.n19 VP.n16 0.278335
R987 VP.n32 VP.n0 0.278335
R988 VP.n10 VP.n9 0.189894
R989 VP.n11 VP.n10 0.189894
R990 VP.n11 VP.n4 0.189894
R991 VP.n20 VP.n19 0.189894
R992 VP.n21 VP.n20 0.189894
R993 VP.n21 VP.n2 0.189894
R994 VP.n26 VP.n2 0.189894
R995 VP.n27 VP.n26 0.189894
R996 VP.n28 VP.n27 0.189894
R997 VP.n28 VP.n0 0.189894
R998 VP VP.n32 0.153485
R999 VDD1 VDD1.t2 265.603
R1000 VDD1.n1 VDD1.t4 265.488
R1001 VDD1.n1 VDD1.n0 236.233
R1002 VDD1.n3 VDD1.n2 235.804
R1003 VDD1.n3 VDD1.n1 32.1755
R1004 VDD1.n2 VDD1.t5 28.2862
R1005 VDD1.n2 VDD1.t1 28.2862
R1006 VDD1.n0 VDD1.t0 28.2862
R1007 VDD1.n0 VDD1.t3 28.2862
R1008 VDD1 VDD1.n3 0.427224
C0 VDD2 VTAIL 3.16304f
C1 VN VDD2 0.723176f
C2 VP VDD1 0.971668f
C3 VN VTAIL 1.52188f
C4 VP VDD2 0.409984f
C5 VP VTAIL 1.536f
C6 VP VN 4.17864f
C7 VDD2 VDD1 1.1646f
C8 VDD1 VTAIL 3.11421f
C9 VN VDD1 0.158451f
C10 VDD2 B 3.26472f
C11 VDD1 B 3.492629f
C12 VTAIL B 2.462178f
C13 VN B 9.518109f
C14 VP B 8.434814f
C15 VDD1.t2 B 0.053295f
C16 VDD1.t4 B 0.05319f
C17 VDD1.t0 B 0.011028f
C18 VDD1.t3 B 0.011028f
C19 VDD1.n0 B 0.027647f
C20 VDD1.n1 B 1.36439f
C21 VDD1.t5 B 0.011028f
C22 VDD1.t1 B 0.011028f
C23 VDD1.n2 B 0.027261f
C24 VDD1.n3 B 1.24537f
C25 VP.n0 B 0.03585f
C26 VP.t2 B 0.053652f
C27 VP.n1 B 0.048304f
C28 VP.n2 B 0.027194f
C29 VP.t5 B 0.053652f
C30 VP.n3 B 0.02791f
C31 VP.n4 B 0.03585f
C32 VP.t4 B 0.053652f
C33 VP.n5 B 0.048304f
C34 VP.t3 B 0.204054f
C35 VP.n6 B 0.10593f
C36 VP.t0 B 0.053652f
C37 VP.n7 B 0.122064f
C38 VP.n8 B 0.037981f
C39 VP.n9 B 0.20142f
C40 VP.n10 B 0.027194f
C41 VP.n11 B 0.027194f
C42 VP.n12 B 0.02791f
C43 VP.n13 B 0.053275f
C44 VP.n14 B 0.146473f
C45 VP.n15 B 0.941986f
C46 VP.n16 B 0.968111f
C47 VP.t1 B 0.053652f
C48 VP.n17 B 0.146473f
C49 VP.n18 B 0.053275f
C50 VP.n19 B 0.03585f
C51 VP.n20 B 0.027194f
C52 VP.n21 B 0.027194f
C53 VP.n22 B 0.048304f
C54 VP.n23 B 0.037981f
C55 VP.n24 B 0.059037f
C56 VP.n25 B 0.037981f
C57 VP.n26 B 0.027194f
C58 VP.n27 B 0.027194f
C59 VP.n28 B 0.027194f
C60 VP.n29 B 0.02791f
C61 VP.n30 B 0.053275f
C62 VP.n31 B 0.146473f
C63 VP.n32 B 0.028736f
C64 VDD2.t2 B 0.056242f
C65 VDD2.t0 B 0.011661f
C66 VDD2.t4 B 0.011661f
C67 VDD2.n0 B 0.029233f
C68 VDD2.n1 B 1.36189f
C69 VDD2.t5 B 0.055383f
C70 VDD2.n2 B 1.26701f
C71 VDD2.t3 B 0.011661f
C72 VDD2.t1 B 0.011661f
C73 VDD2.n3 B 0.029228f
C74 VTAIL.t8 B 0.017503f
C75 VTAIL.t7 B 0.017503f
C76 VTAIL.n0 B 0.037579f
C77 VTAIL.n1 B 0.245571f
C78 VTAIL.t3 B 0.077561f
C79 VTAIL.n2 B 0.395709f
C80 VTAIL.t2 B 0.017503f
C81 VTAIL.t0 B 0.017503f
C82 VTAIL.n3 B 0.037579f
C83 VTAIL.n4 B 1.12802f
C84 VTAIL.t11 B 0.017503f
C85 VTAIL.t10 B 0.017503f
C86 VTAIL.n5 B 0.037579f
C87 VTAIL.n6 B 1.12802f
C88 VTAIL.t9 B 0.077561f
C89 VTAIL.n7 B 0.395709f
C90 VTAIL.t4 B 0.017503f
C91 VTAIL.t5 B 0.017503f
C92 VTAIL.n8 B 0.037579f
C93 VTAIL.n9 B 0.387956f
C94 VTAIL.t1 B 0.077561f
C95 VTAIL.n10 B 0.93802f
C96 VTAIL.t6 B 0.077561f
C97 VTAIL.n11 B 0.882648f
C98 VN.n0 B 0.035527f
C99 VN.t1 B 0.053168f
C100 VN.n1 B 0.047869f
C101 VN.t3 B 0.202214f
C102 VN.n2 B 0.104974f
C103 VN.t5 B 0.053168f
C104 VN.n3 B 0.120963f
C105 VN.n4 B 0.037638f
C106 VN.n5 B 0.199603f
C107 VN.n6 B 0.026949f
C108 VN.n7 B 0.026949f
C109 VN.n8 B 0.027658f
C110 VN.n9 B 0.052794f
C111 VN.n10 B 0.145152f
C112 VN.n11 B 0.028477f
C113 VN.n12 B 0.035527f
C114 VN.t0 B 0.053168f
C115 VN.n13 B 0.047869f
C116 VN.t4 B 0.202214f
C117 VN.n14 B 0.104974f
C118 VN.t2 B 0.053168f
C119 VN.n15 B 0.120963f
C120 VN.n16 B 0.037638f
C121 VN.n17 B 0.199603f
C122 VN.n18 B 0.026949f
C123 VN.n19 B 0.026949f
C124 VN.n20 B 0.027658f
C125 VN.n21 B 0.052794f
C126 VN.n22 B 0.145152f
C127 VN.n23 B 0.948735f
.ends

