* NGSPICE file created from diff_pair_sample_1347.ext - technology: sky130A

.subckt diff_pair_sample_1347 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X1 VDD1.t1 VP.t1 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X2 VTAIL.t4 VN.t0 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0.29205 ps=2.1 w=1.77 l=1.49
X3 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=1.49
X4 VDD1.t6 VP.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.6903 ps=4.32 w=1.77 l=1.49
X5 VTAIL.t0 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=1.49
X7 VTAIL.t12 VP.t3 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0.29205 ps=2.1 w=1.77 l=1.49
X8 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.6903 ps=4.32 w=1.77 l=1.49
X9 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X10 VTAIL.t11 VP.t4 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0.29205 ps=2.1 w=1.77 l=1.49
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=1.49
X12 VTAIL.t10 VP.t5 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X13 VDD2.t3 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X14 VDD1.t0 VP.t6 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.6903 ps=4.32 w=1.77 l=1.49
X15 VDD2.t2 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.6903 ps=4.32 w=1.77 l=1.49
X16 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X17 VDD1.t2 VP.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.29205 pd=2.1 as=0.29205 ps=2.1 w=1.77 l=1.49
X18 VTAIL.t7 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0.29205 ps=2.1 w=1.77 l=1.49
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=1.49
R0 VP.n26 VP.n25 174.512
R1 VP.n46 VP.n45 174.512
R2 VP.n24 VP.n23 174.512
R3 VP.n12 VP.n9 161.3
R4 VP.n14 VP.n13 161.3
R5 VP.n15 VP.n8 161.3
R6 VP.n18 VP.n17 161.3
R7 VP.n19 VP.n7 161.3
R8 VP.n21 VP.n20 161.3
R9 VP.n22 VP.n6 161.3
R10 VP.n44 VP.n0 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n1 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n37 VP.n2 161.3
R15 VP.n36 VP.n35 161.3
R16 VP.n34 VP.n3 161.3
R17 VP.n33 VP.n32 161.3
R18 VP.n30 VP.n4 161.3
R19 VP.n29 VP.n28 161.3
R20 VP.n27 VP.n5 161.3
R21 VP.n11 VP.t4 63.006
R22 VP.n30 VP.n29 56.5193
R23 VP.n21 VP.n7 56.5193
R24 VP.n43 VP.n1 56.5193
R25 VP.n11 VP.n10 46.4328
R26 VP.n36 VP.n3 40.4934
R27 VP.n37 VP.n36 40.4934
R28 VP.n15 VP.n14 40.4934
R29 VP.n14 VP.n9 40.4934
R30 VP.n26 VP.n24 37.8944
R31 VP.n25 VP.t3 28.6294
R32 VP.n31 VP.t1 28.6294
R33 VP.n38 VP.t5 28.6294
R34 VP.n45 VP.t2 28.6294
R35 VP.n23 VP.t6 28.6294
R36 VP.n16 VP.t0 28.6294
R37 VP.n10 VP.t7 28.6294
R38 VP.n29 VP.n5 24.4675
R39 VP.n32 VP.n30 24.4675
R40 VP.n39 VP.n1 24.4675
R41 VP.n44 VP.n43 24.4675
R42 VP.n22 VP.n21 24.4675
R43 VP.n17 VP.n7 24.4675
R44 VP.n31 VP.n3 20.0634
R45 VP.n38 VP.n37 20.0634
R46 VP.n16 VP.n15 20.0634
R47 VP.n10 VP.n9 20.0634
R48 VP.n12 VP.n11 17.6611
R49 VP.n25 VP.n5 11.2553
R50 VP.n45 VP.n44 11.2553
R51 VP.n23 VP.n22 11.2553
R52 VP.n32 VP.n31 4.40456
R53 VP.n39 VP.n38 4.40456
R54 VP.n17 VP.n16 4.40456
R55 VP.n13 VP.n12 0.189894
R56 VP.n13 VP.n8 0.189894
R57 VP.n18 VP.n8 0.189894
R58 VP.n19 VP.n18 0.189894
R59 VP.n20 VP.n19 0.189894
R60 VP.n20 VP.n6 0.189894
R61 VP.n24 VP.n6 0.189894
R62 VP.n27 VP.n26 0.189894
R63 VP.n28 VP.n27 0.189894
R64 VP.n28 VP.n4 0.189894
R65 VP.n33 VP.n4 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n35 VP.n34 0.189894
R68 VP.n35 VP.n2 0.189894
R69 VP.n40 VP.n2 0.189894
R70 VP.n41 VP.n40 0.189894
R71 VP.n42 VP.n41 0.189894
R72 VP.n42 VP.n0 0.189894
R73 VP.n46 VP.n0 0.189894
R74 VP VP.n46 0.0516364
R75 VDD1 VDD1.n0 102.072
R76 VDD1.n3 VDD1.n2 101.959
R77 VDD1.n3 VDD1.n1 101.959
R78 VDD1.n5 VDD1.n4 101.23
R79 VDD1.n5 VDD1.n3 32.8845
R80 VDD1.n4 VDD1.t4 11.1869
R81 VDD1.n4 VDD1.t0 11.1869
R82 VDD1.n0 VDD1.t7 11.1869
R83 VDD1.n0 VDD1.t2 11.1869
R84 VDD1.n2 VDD1.t3 11.1869
R85 VDD1.n2 VDD1.t6 11.1869
R86 VDD1.n1 VDD1.t5 11.1869
R87 VDD1.n1 VDD1.t1 11.1869
R88 VDD1 VDD1.n5 0.726793
R89 VTAIL.n66 VTAIL.n64 289.615
R90 VTAIL.n4 VTAIL.n2 289.615
R91 VTAIL.n12 VTAIL.n10 289.615
R92 VTAIL.n22 VTAIL.n20 289.615
R93 VTAIL.n58 VTAIL.n56 289.615
R94 VTAIL.n48 VTAIL.n46 289.615
R95 VTAIL.n40 VTAIL.n38 289.615
R96 VTAIL.n30 VTAIL.n28 289.615
R97 VTAIL.n67 VTAIL.n66 185
R98 VTAIL.n5 VTAIL.n4 185
R99 VTAIL.n13 VTAIL.n12 185
R100 VTAIL.n23 VTAIL.n22 185
R101 VTAIL.n59 VTAIL.n58 185
R102 VTAIL.n49 VTAIL.n48 185
R103 VTAIL.n41 VTAIL.n40 185
R104 VTAIL.n31 VTAIL.n30 185
R105 VTAIL.t1 VTAIL.n65 164.876
R106 VTAIL.t7 VTAIL.n3 164.876
R107 VTAIL.t13 VTAIL.n11 164.876
R108 VTAIL.t12 VTAIL.n21 164.876
R109 VTAIL.t9 VTAIL.n57 164.876
R110 VTAIL.t11 VTAIL.n47 164.876
R111 VTAIL.t3 VTAIL.n39 164.876
R112 VTAIL.t4 VTAIL.n29 164.876
R113 VTAIL.n55 VTAIL.n54 84.5504
R114 VTAIL.n37 VTAIL.n36 84.5504
R115 VTAIL.n1 VTAIL.n0 84.5503
R116 VTAIL.n19 VTAIL.n18 84.5503
R117 VTAIL.n66 VTAIL.t1 52.3082
R118 VTAIL.n4 VTAIL.t7 52.3082
R119 VTAIL.n12 VTAIL.t13 52.3082
R120 VTAIL.n22 VTAIL.t12 52.3082
R121 VTAIL.n58 VTAIL.t9 52.3082
R122 VTAIL.n48 VTAIL.t11 52.3082
R123 VTAIL.n40 VTAIL.t3 52.3082
R124 VTAIL.n30 VTAIL.t4 52.3082
R125 VTAIL.n71 VTAIL.n70 33.9308
R126 VTAIL.n9 VTAIL.n8 33.9308
R127 VTAIL.n17 VTAIL.n16 33.9308
R128 VTAIL.n27 VTAIL.n26 33.9308
R129 VTAIL.n63 VTAIL.n62 33.9308
R130 VTAIL.n53 VTAIL.n52 33.9308
R131 VTAIL.n45 VTAIL.n44 33.9308
R132 VTAIL.n35 VTAIL.n34 33.9308
R133 VTAIL.n71 VTAIL.n63 15.4617
R134 VTAIL.n35 VTAIL.n27 15.4617
R135 VTAIL.n67 VTAIL.n65 14.7318
R136 VTAIL.n5 VTAIL.n3 14.7318
R137 VTAIL.n13 VTAIL.n11 14.7318
R138 VTAIL.n23 VTAIL.n21 14.7318
R139 VTAIL.n59 VTAIL.n57 14.7318
R140 VTAIL.n49 VTAIL.n47 14.7318
R141 VTAIL.n41 VTAIL.n39 14.7318
R142 VTAIL.n31 VTAIL.n29 14.7318
R143 VTAIL.n68 VTAIL.n64 12.8005
R144 VTAIL.n6 VTAIL.n2 12.8005
R145 VTAIL.n14 VTAIL.n10 12.8005
R146 VTAIL.n24 VTAIL.n20 12.8005
R147 VTAIL.n60 VTAIL.n56 12.8005
R148 VTAIL.n50 VTAIL.n46 12.8005
R149 VTAIL.n42 VTAIL.n38 12.8005
R150 VTAIL.n32 VTAIL.n28 12.8005
R151 VTAIL.n0 VTAIL.t6 11.1869
R152 VTAIL.n0 VTAIL.t2 11.1869
R153 VTAIL.n18 VTAIL.t14 11.1869
R154 VTAIL.n18 VTAIL.t10 11.1869
R155 VTAIL.n54 VTAIL.t8 11.1869
R156 VTAIL.n54 VTAIL.t15 11.1869
R157 VTAIL.n36 VTAIL.t5 11.1869
R158 VTAIL.n36 VTAIL.t0 11.1869
R159 VTAIL.n70 VTAIL.n69 9.45567
R160 VTAIL.n8 VTAIL.n7 9.45567
R161 VTAIL.n16 VTAIL.n15 9.45567
R162 VTAIL.n26 VTAIL.n25 9.45567
R163 VTAIL.n62 VTAIL.n61 9.45567
R164 VTAIL.n52 VTAIL.n51 9.45567
R165 VTAIL.n44 VTAIL.n43 9.45567
R166 VTAIL.n34 VTAIL.n33 9.45567
R167 VTAIL.n69 VTAIL.n68 9.3005
R168 VTAIL.n7 VTAIL.n6 9.3005
R169 VTAIL.n15 VTAIL.n14 9.3005
R170 VTAIL.n25 VTAIL.n24 9.3005
R171 VTAIL.n61 VTAIL.n60 9.3005
R172 VTAIL.n51 VTAIL.n50 9.3005
R173 VTAIL.n43 VTAIL.n42 9.3005
R174 VTAIL.n33 VTAIL.n32 9.3005
R175 VTAIL.n69 VTAIL.n65 5.62509
R176 VTAIL.n7 VTAIL.n3 5.62509
R177 VTAIL.n15 VTAIL.n11 5.62509
R178 VTAIL.n25 VTAIL.n21 5.62509
R179 VTAIL.n61 VTAIL.n57 5.62509
R180 VTAIL.n51 VTAIL.n47 5.62509
R181 VTAIL.n43 VTAIL.n39 5.62509
R182 VTAIL.n33 VTAIL.n29 5.62509
R183 VTAIL.n37 VTAIL.n35 1.56947
R184 VTAIL.n45 VTAIL.n37 1.56947
R185 VTAIL.n55 VTAIL.n53 1.56947
R186 VTAIL.n63 VTAIL.n55 1.56947
R187 VTAIL.n27 VTAIL.n19 1.56947
R188 VTAIL.n19 VTAIL.n17 1.56947
R189 VTAIL.n9 VTAIL.n1 1.56947
R190 VTAIL VTAIL.n71 1.51128
R191 VTAIL.n70 VTAIL.n64 1.16414
R192 VTAIL.n8 VTAIL.n2 1.16414
R193 VTAIL.n16 VTAIL.n10 1.16414
R194 VTAIL.n26 VTAIL.n20 1.16414
R195 VTAIL.n62 VTAIL.n56 1.16414
R196 VTAIL.n52 VTAIL.n46 1.16414
R197 VTAIL.n44 VTAIL.n38 1.16414
R198 VTAIL.n34 VTAIL.n28 1.16414
R199 VTAIL.n53 VTAIL.n45 0.470328
R200 VTAIL.n17 VTAIL.n9 0.470328
R201 VTAIL.n68 VTAIL.n67 0.388379
R202 VTAIL.n6 VTAIL.n5 0.388379
R203 VTAIL.n14 VTAIL.n13 0.388379
R204 VTAIL.n24 VTAIL.n23 0.388379
R205 VTAIL.n60 VTAIL.n59 0.388379
R206 VTAIL.n50 VTAIL.n49 0.388379
R207 VTAIL.n42 VTAIL.n41 0.388379
R208 VTAIL.n32 VTAIL.n31 0.388379
R209 VTAIL VTAIL.n1 0.0586897
R210 B.n456 B.n455 585
R211 B.n457 B.n456 585
R212 B.n149 B.n83 585
R213 B.n148 B.n147 585
R214 B.n146 B.n145 585
R215 B.n144 B.n143 585
R216 B.n142 B.n141 585
R217 B.n140 B.n139 585
R218 B.n138 B.n137 585
R219 B.n136 B.n135 585
R220 B.n134 B.n133 585
R221 B.n132 B.n131 585
R222 B.n130 B.n129 585
R223 B.n127 B.n126 585
R224 B.n125 B.n124 585
R225 B.n123 B.n122 585
R226 B.n121 B.n120 585
R227 B.n119 B.n118 585
R228 B.n117 B.n116 585
R229 B.n115 B.n114 585
R230 B.n113 B.n112 585
R231 B.n111 B.n110 585
R232 B.n109 B.n108 585
R233 B.n107 B.n106 585
R234 B.n105 B.n104 585
R235 B.n103 B.n102 585
R236 B.n101 B.n100 585
R237 B.n99 B.n98 585
R238 B.n97 B.n96 585
R239 B.n95 B.n94 585
R240 B.n93 B.n92 585
R241 B.n91 B.n90 585
R242 B.n67 B.n66 585
R243 B.n460 B.n459 585
R244 B.n454 B.n84 585
R245 B.n84 B.n64 585
R246 B.n453 B.n63 585
R247 B.n464 B.n63 585
R248 B.n452 B.n62 585
R249 B.n465 B.n62 585
R250 B.n451 B.n61 585
R251 B.n466 B.n61 585
R252 B.n450 B.n449 585
R253 B.n449 B.n57 585
R254 B.n448 B.n56 585
R255 B.n472 B.n56 585
R256 B.n447 B.n55 585
R257 B.n473 B.n55 585
R258 B.n446 B.n54 585
R259 B.n474 B.n54 585
R260 B.n445 B.n444 585
R261 B.n444 B.n50 585
R262 B.n443 B.n49 585
R263 B.n480 B.n49 585
R264 B.n442 B.n48 585
R265 B.n481 B.n48 585
R266 B.n441 B.n47 585
R267 B.n482 B.n47 585
R268 B.n440 B.n439 585
R269 B.n439 B.n43 585
R270 B.n438 B.n42 585
R271 B.n488 B.n42 585
R272 B.n437 B.n41 585
R273 B.n489 B.n41 585
R274 B.n436 B.n40 585
R275 B.n490 B.n40 585
R276 B.n435 B.n434 585
R277 B.n434 B.n36 585
R278 B.n433 B.n35 585
R279 B.n496 B.n35 585
R280 B.n432 B.n34 585
R281 B.n497 B.n34 585
R282 B.n431 B.n33 585
R283 B.n498 B.n33 585
R284 B.n430 B.n429 585
R285 B.n429 B.n32 585
R286 B.n428 B.n28 585
R287 B.n504 B.n28 585
R288 B.n427 B.n27 585
R289 B.n505 B.n27 585
R290 B.n426 B.n26 585
R291 B.n506 B.n26 585
R292 B.n425 B.n424 585
R293 B.n424 B.n22 585
R294 B.n423 B.n21 585
R295 B.n512 B.n21 585
R296 B.n422 B.n20 585
R297 B.n513 B.n20 585
R298 B.n421 B.n19 585
R299 B.n514 B.n19 585
R300 B.n420 B.n419 585
R301 B.n419 B.n15 585
R302 B.n418 B.n14 585
R303 B.n520 B.n14 585
R304 B.n417 B.n13 585
R305 B.n521 B.n13 585
R306 B.n416 B.n12 585
R307 B.n522 B.n12 585
R308 B.n415 B.n414 585
R309 B.n414 B.n8 585
R310 B.n413 B.n7 585
R311 B.n528 B.n7 585
R312 B.n412 B.n6 585
R313 B.n529 B.n6 585
R314 B.n411 B.n5 585
R315 B.n530 B.n5 585
R316 B.n410 B.n409 585
R317 B.n409 B.n4 585
R318 B.n408 B.n150 585
R319 B.n408 B.n407 585
R320 B.n398 B.n151 585
R321 B.n152 B.n151 585
R322 B.n400 B.n399 585
R323 B.n401 B.n400 585
R324 B.n397 B.n156 585
R325 B.n160 B.n156 585
R326 B.n396 B.n395 585
R327 B.n395 B.n394 585
R328 B.n158 B.n157 585
R329 B.n159 B.n158 585
R330 B.n387 B.n386 585
R331 B.n388 B.n387 585
R332 B.n385 B.n165 585
R333 B.n165 B.n164 585
R334 B.n384 B.n383 585
R335 B.n383 B.n382 585
R336 B.n167 B.n166 585
R337 B.n168 B.n167 585
R338 B.n375 B.n374 585
R339 B.n376 B.n375 585
R340 B.n373 B.n173 585
R341 B.n173 B.n172 585
R342 B.n372 B.n371 585
R343 B.n371 B.n370 585
R344 B.n175 B.n174 585
R345 B.n363 B.n175 585
R346 B.n362 B.n361 585
R347 B.n364 B.n362 585
R348 B.n360 B.n180 585
R349 B.n180 B.n179 585
R350 B.n359 B.n358 585
R351 B.n358 B.n357 585
R352 B.n182 B.n181 585
R353 B.n183 B.n182 585
R354 B.n350 B.n349 585
R355 B.n351 B.n350 585
R356 B.n348 B.n187 585
R357 B.n191 B.n187 585
R358 B.n347 B.n346 585
R359 B.n346 B.n345 585
R360 B.n189 B.n188 585
R361 B.n190 B.n189 585
R362 B.n338 B.n337 585
R363 B.n339 B.n338 585
R364 B.n336 B.n196 585
R365 B.n196 B.n195 585
R366 B.n335 B.n334 585
R367 B.n334 B.n333 585
R368 B.n198 B.n197 585
R369 B.n199 B.n198 585
R370 B.n326 B.n325 585
R371 B.n327 B.n326 585
R372 B.n324 B.n203 585
R373 B.n207 B.n203 585
R374 B.n323 B.n322 585
R375 B.n322 B.n321 585
R376 B.n205 B.n204 585
R377 B.n206 B.n205 585
R378 B.n314 B.n313 585
R379 B.n315 B.n314 585
R380 B.n312 B.n212 585
R381 B.n212 B.n211 585
R382 B.n311 B.n310 585
R383 B.n310 B.n309 585
R384 B.n214 B.n213 585
R385 B.n215 B.n214 585
R386 B.n305 B.n304 585
R387 B.n218 B.n217 585
R388 B.n301 B.n300 585
R389 B.n302 B.n301 585
R390 B.n299 B.n234 585
R391 B.n298 B.n297 585
R392 B.n296 B.n295 585
R393 B.n294 B.n293 585
R394 B.n292 B.n291 585
R395 B.n290 B.n289 585
R396 B.n288 B.n287 585
R397 B.n286 B.n285 585
R398 B.n284 B.n283 585
R399 B.n281 B.n280 585
R400 B.n279 B.n278 585
R401 B.n277 B.n276 585
R402 B.n275 B.n274 585
R403 B.n273 B.n272 585
R404 B.n271 B.n270 585
R405 B.n269 B.n268 585
R406 B.n267 B.n266 585
R407 B.n265 B.n264 585
R408 B.n263 B.n262 585
R409 B.n261 B.n260 585
R410 B.n259 B.n258 585
R411 B.n257 B.n256 585
R412 B.n255 B.n254 585
R413 B.n253 B.n252 585
R414 B.n251 B.n250 585
R415 B.n249 B.n248 585
R416 B.n247 B.n246 585
R417 B.n245 B.n244 585
R418 B.n243 B.n242 585
R419 B.n241 B.n240 585
R420 B.n306 B.n216 585
R421 B.n216 B.n215 585
R422 B.n308 B.n307 585
R423 B.n309 B.n308 585
R424 B.n210 B.n209 585
R425 B.n211 B.n210 585
R426 B.n317 B.n316 585
R427 B.n316 B.n315 585
R428 B.n318 B.n208 585
R429 B.n208 B.n206 585
R430 B.n320 B.n319 585
R431 B.n321 B.n320 585
R432 B.n202 B.n201 585
R433 B.n207 B.n202 585
R434 B.n329 B.n328 585
R435 B.n328 B.n327 585
R436 B.n330 B.n200 585
R437 B.n200 B.n199 585
R438 B.n332 B.n331 585
R439 B.n333 B.n332 585
R440 B.n194 B.n193 585
R441 B.n195 B.n194 585
R442 B.n341 B.n340 585
R443 B.n340 B.n339 585
R444 B.n342 B.n192 585
R445 B.n192 B.n190 585
R446 B.n344 B.n343 585
R447 B.n345 B.n344 585
R448 B.n186 B.n185 585
R449 B.n191 B.n186 585
R450 B.n353 B.n352 585
R451 B.n352 B.n351 585
R452 B.n354 B.n184 585
R453 B.n184 B.n183 585
R454 B.n356 B.n355 585
R455 B.n357 B.n356 585
R456 B.n178 B.n177 585
R457 B.n179 B.n178 585
R458 B.n366 B.n365 585
R459 B.n365 B.n364 585
R460 B.n367 B.n176 585
R461 B.n363 B.n176 585
R462 B.n369 B.n368 585
R463 B.n370 B.n369 585
R464 B.n171 B.n170 585
R465 B.n172 B.n171 585
R466 B.n378 B.n377 585
R467 B.n377 B.n376 585
R468 B.n379 B.n169 585
R469 B.n169 B.n168 585
R470 B.n381 B.n380 585
R471 B.n382 B.n381 585
R472 B.n163 B.n162 585
R473 B.n164 B.n163 585
R474 B.n390 B.n389 585
R475 B.n389 B.n388 585
R476 B.n391 B.n161 585
R477 B.n161 B.n159 585
R478 B.n393 B.n392 585
R479 B.n394 B.n393 585
R480 B.n155 B.n154 585
R481 B.n160 B.n155 585
R482 B.n403 B.n402 585
R483 B.n402 B.n401 585
R484 B.n404 B.n153 585
R485 B.n153 B.n152 585
R486 B.n406 B.n405 585
R487 B.n407 B.n406 585
R488 B.n2 B.n0 585
R489 B.n4 B.n2 585
R490 B.n3 B.n1 585
R491 B.n529 B.n3 585
R492 B.n527 B.n526 585
R493 B.n528 B.n527 585
R494 B.n525 B.n9 585
R495 B.n9 B.n8 585
R496 B.n524 B.n523 585
R497 B.n523 B.n522 585
R498 B.n11 B.n10 585
R499 B.n521 B.n11 585
R500 B.n519 B.n518 585
R501 B.n520 B.n519 585
R502 B.n517 B.n16 585
R503 B.n16 B.n15 585
R504 B.n516 B.n515 585
R505 B.n515 B.n514 585
R506 B.n18 B.n17 585
R507 B.n513 B.n18 585
R508 B.n511 B.n510 585
R509 B.n512 B.n511 585
R510 B.n509 B.n23 585
R511 B.n23 B.n22 585
R512 B.n508 B.n507 585
R513 B.n507 B.n506 585
R514 B.n25 B.n24 585
R515 B.n505 B.n25 585
R516 B.n503 B.n502 585
R517 B.n504 B.n503 585
R518 B.n501 B.n29 585
R519 B.n32 B.n29 585
R520 B.n500 B.n499 585
R521 B.n499 B.n498 585
R522 B.n31 B.n30 585
R523 B.n497 B.n31 585
R524 B.n495 B.n494 585
R525 B.n496 B.n495 585
R526 B.n493 B.n37 585
R527 B.n37 B.n36 585
R528 B.n492 B.n491 585
R529 B.n491 B.n490 585
R530 B.n39 B.n38 585
R531 B.n489 B.n39 585
R532 B.n487 B.n486 585
R533 B.n488 B.n487 585
R534 B.n485 B.n44 585
R535 B.n44 B.n43 585
R536 B.n484 B.n483 585
R537 B.n483 B.n482 585
R538 B.n46 B.n45 585
R539 B.n481 B.n46 585
R540 B.n479 B.n478 585
R541 B.n480 B.n479 585
R542 B.n477 B.n51 585
R543 B.n51 B.n50 585
R544 B.n476 B.n475 585
R545 B.n475 B.n474 585
R546 B.n53 B.n52 585
R547 B.n473 B.n53 585
R548 B.n471 B.n470 585
R549 B.n472 B.n471 585
R550 B.n469 B.n58 585
R551 B.n58 B.n57 585
R552 B.n468 B.n467 585
R553 B.n467 B.n466 585
R554 B.n60 B.n59 585
R555 B.n465 B.n60 585
R556 B.n463 B.n462 585
R557 B.n464 B.n463 585
R558 B.n461 B.n65 585
R559 B.n65 B.n64 585
R560 B.n532 B.n531 585
R561 B.n531 B.n530 585
R562 B.n304 B.n216 449.257
R563 B.n459 B.n65 449.257
R564 B.n240 B.n214 449.257
R565 B.n456 B.n84 449.257
R566 B.n457 B.n82 256.663
R567 B.n457 B.n81 256.663
R568 B.n457 B.n80 256.663
R569 B.n457 B.n79 256.663
R570 B.n457 B.n78 256.663
R571 B.n457 B.n77 256.663
R572 B.n457 B.n76 256.663
R573 B.n457 B.n75 256.663
R574 B.n457 B.n74 256.663
R575 B.n457 B.n73 256.663
R576 B.n457 B.n72 256.663
R577 B.n457 B.n71 256.663
R578 B.n457 B.n70 256.663
R579 B.n457 B.n69 256.663
R580 B.n457 B.n68 256.663
R581 B.n458 B.n457 256.663
R582 B.n303 B.n302 256.663
R583 B.n302 B.n219 256.663
R584 B.n302 B.n220 256.663
R585 B.n302 B.n221 256.663
R586 B.n302 B.n222 256.663
R587 B.n302 B.n223 256.663
R588 B.n302 B.n224 256.663
R589 B.n302 B.n225 256.663
R590 B.n302 B.n226 256.663
R591 B.n302 B.n227 256.663
R592 B.n302 B.n228 256.663
R593 B.n302 B.n229 256.663
R594 B.n302 B.n230 256.663
R595 B.n302 B.n231 256.663
R596 B.n302 B.n232 256.663
R597 B.n302 B.n233 256.663
R598 B.n237 B.t8 234.031
R599 B.n235 B.t19 234.031
R600 B.n87 B.t12 234.031
R601 B.n85 B.t16 234.031
R602 B.n302 B.n215 179.56
R603 B.n457 B.n64 179.56
R604 B.n308 B.n216 163.367
R605 B.n308 B.n210 163.367
R606 B.n316 B.n210 163.367
R607 B.n316 B.n208 163.367
R608 B.n320 B.n208 163.367
R609 B.n320 B.n202 163.367
R610 B.n328 B.n202 163.367
R611 B.n328 B.n200 163.367
R612 B.n332 B.n200 163.367
R613 B.n332 B.n194 163.367
R614 B.n340 B.n194 163.367
R615 B.n340 B.n192 163.367
R616 B.n344 B.n192 163.367
R617 B.n344 B.n186 163.367
R618 B.n352 B.n186 163.367
R619 B.n352 B.n184 163.367
R620 B.n356 B.n184 163.367
R621 B.n356 B.n178 163.367
R622 B.n365 B.n178 163.367
R623 B.n365 B.n176 163.367
R624 B.n369 B.n176 163.367
R625 B.n369 B.n171 163.367
R626 B.n377 B.n171 163.367
R627 B.n377 B.n169 163.367
R628 B.n381 B.n169 163.367
R629 B.n381 B.n163 163.367
R630 B.n389 B.n163 163.367
R631 B.n389 B.n161 163.367
R632 B.n393 B.n161 163.367
R633 B.n393 B.n155 163.367
R634 B.n402 B.n155 163.367
R635 B.n402 B.n153 163.367
R636 B.n406 B.n153 163.367
R637 B.n406 B.n2 163.367
R638 B.n531 B.n2 163.367
R639 B.n531 B.n3 163.367
R640 B.n527 B.n3 163.367
R641 B.n527 B.n9 163.367
R642 B.n523 B.n9 163.367
R643 B.n523 B.n11 163.367
R644 B.n519 B.n11 163.367
R645 B.n519 B.n16 163.367
R646 B.n515 B.n16 163.367
R647 B.n515 B.n18 163.367
R648 B.n511 B.n18 163.367
R649 B.n511 B.n23 163.367
R650 B.n507 B.n23 163.367
R651 B.n507 B.n25 163.367
R652 B.n503 B.n25 163.367
R653 B.n503 B.n29 163.367
R654 B.n499 B.n29 163.367
R655 B.n499 B.n31 163.367
R656 B.n495 B.n31 163.367
R657 B.n495 B.n37 163.367
R658 B.n491 B.n37 163.367
R659 B.n491 B.n39 163.367
R660 B.n487 B.n39 163.367
R661 B.n487 B.n44 163.367
R662 B.n483 B.n44 163.367
R663 B.n483 B.n46 163.367
R664 B.n479 B.n46 163.367
R665 B.n479 B.n51 163.367
R666 B.n475 B.n51 163.367
R667 B.n475 B.n53 163.367
R668 B.n471 B.n53 163.367
R669 B.n471 B.n58 163.367
R670 B.n467 B.n58 163.367
R671 B.n467 B.n60 163.367
R672 B.n463 B.n60 163.367
R673 B.n463 B.n65 163.367
R674 B.n301 B.n218 163.367
R675 B.n301 B.n234 163.367
R676 B.n297 B.n296 163.367
R677 B.n293 B.n292 163.367
R678 B.n289 B.n288 163.367
R679 B.n285 B.n284 163.367
R680 B.n280 B.n279 163.367
R681 B.n276 B.n275 163.367
R682 B.n272 B.n271 163.367
R683 B.n268 B.n267 163.367
R684 B.n264 B.n263 163.367
R685 B.n260 B.n259 163.367
R686 B.n256 B.n255 163.367
R687 B.n252 B.n251 163.367
R688 B.n248 B.n247 163.367
R689 B.n244 B.n243 163.367
R690 B.n310 B.n214 163.367
R691 B.n310 B.n212 163.367
R692 B.n314 B.n212 163.367
R693 B.n314 B.n205 163.367
R694 B.n322 B.n205 163.367
R695 B.n322 B.n203 163.367
R696 B.n326 B.n203 163.367
R697 B.n326 B.n198 163.367
R698 B.n334 B.n198 163.367
R699 B.n334 B.n196 163.367
R700 B.n338 B.n196 163.367
R701 B.n338 B.n189 163.367
R702 B.n346 B.n189 163.367
R703 B.n346 B.n187 163.367
R704 B.n350 B.n187 163.367
R705 B.n350 B.n182 163.367
R706 B.n358 B.n182 163.367
R707 B.n358 B.n180 163.367
R708 B.n362 B.n180 163.367
R709 B.n362 B.n175 163.367
R710 B.n371 B.n175 163.367
R711 B.n371 B.n173 163.367
R712 B.n375 B.n173 163.367
R713 B.n375 B.n167 163.367
R714 B.n383 B.n167 163.367
R715 B.n383 B.n165 163.367
R716 B.n387 B.n165 163.367
R717 B.n387 B.n158 163.367
R718 B.n395 B.n158 163.367
R719 B.n395 B.n156 163.367
R720 B.n400 B.n156 163.367
R721 B.n400 B.n151 163.367
R722 B.n408 B.n151 163.367
R723 B.n409 B.n408 163.367
R724 B.n409 B.n5 163.367
R725 B.n6 B.n5 163.367
R726 B.n7 B.n6 163.367
R727 B.n414 B.n7 163.367
R728 B.n414 B.n12 163.367
R729 B.n13 B.n12 163.367
R730 B.n14 B.n13 163.367
R731 B.n419 B.n14 163.367
R732 B.n419 B.n19 163.367
R733 B.n20 B.n19 163.367
R734 B.n21 B.n20 163.367
R735 B.n424 B.n21 163.367
R736 B.n424 B.n26 163.367
R737 B.n27 B.n26 163.367
R738 B.n28 B.n27 163.367
R739 B.n429 B.n28 163.367
R740 B.n429 B.n33 163.367
R741 B.n34 B.n33 163.367
R742 B.n35 B.n34 163.367
R743 B.n434 B.n35 163.367
R744 B.n434 B.n40 163.367
R745 B.n41 B.n40 163.367
R746 B.n42 B.n41 163.367
R747 B.n439 B.n42 163.367
R748 B.n439 B.n47 163.367
R749 B.n48 B.n47 163.367
R750 B.n49 B.n48 163.367
R751 B.n444 B.n49 163.367
R752 B.n444 B.n54 163.367
R753 B.n55 B.n54 163.367
R754 B.n56 B.n55 163.367
R755 B.n449 B.n56 163.367
R756 B.n449 B.n61 163.367
R757 B.n62 B.n61 163.367
R758 B.n63 B.n62 163.367
R759 B.n84 B.n63 163.367
R760 B.n90 B.n67 163.367
R761 B.n94 B.n93 163.367
R762 B.n98 B.n97 163.367
R763 B.n102 B.n101 163.367
R764 B.n106 B.n105 163.367
R765 B.n110 B.n109 163.367
R766 B.n114 B.n113 163.367
R767 B.n118 B.n117 163.367
R768 B.n122 B.n121 163.367
R769 B.n126 B.n125 163.367
R770 B.n131 B.n130 163.367
R771 B.n135 B.n134 163.367
R772 B.n139 B.n138 163.367
R773 B.n143 B.n142 163.367
R774 B.n147 B.n146 163.367
R775 B.n456 B.n83 163.367
R776 B.n237 B.t11 153.855
R777 B.n85 B.t17 153.855
R778 B.n235 B.t21 153.855
R779 B.n87 B.t14 153.855
R780 B.n238 B.t10 118.558
R781 B.n86 B.t18 118.558
R782 B.n236 B.t20 118.558
R783 B.n88 B.t15 118.558
R784 B.n309 B.n215 106.175
R785 B.n309 B.n211 106.175
R786 B.n315 B.n211 106.175
R787 B.n315 B.n206 106.175
R788 B.n321 B.n206 106.175
R789 B.n321 B.n207 106.175
R790 B.n327 B.n199 106.175
R791 B.n333 B.n199 106.175
R792 B.n333 B.n195 106.175
R793 B.n339 B.n195 106.175
R794 B.n339 B.n190 106.175
R795 B.n345 B.n190 106.175
R796 B.n345 B.n191 106.175
R797 B.n351 B.n183 106.175
R798 B.n357 B.n183 106.175
R799 B.n357 B.n179 106.175
R800 B.n364 B.n179 106.175
R801 B.n364 B.n363 106.175
R802 B.n370 B.n172 106.175
R803 B.n376 B.n172 106.175
R804 B.n376 B.n168 106.175
R805 B.n382 B.n168 106.175
R806 B.n388 B.n164 106.175
R807 B.n388 B.n159 106.175
R808 B.n394 B.n159 106.175
R809 B.n394 B.n160 106.175
R810 B.n401 B.n152 106.175
R811 B.n407 B.n152 106.175
R812 B.n407 B.n4 106.175
R813 B.n530 B.n4 106.175
R814 B.n530 B.n529 106.175
R815 B.n529 B.n528 106.175
R816 B.n528 B.n8 106.175
R817 B.n522 B.n8 106.175
R818 B.n521 B.n520 106.175
R819 B.n520 B.n15 106.175
R820 B.n514 B.n15 106.175
R821 B.n514 B.n513 106.175
R822 B.n512 B.n22 106.175
R823 B.n506 B.n22 106.175
R824 B.n506 B.n505 106.175
R825 B.n505 B.n504 106.175
R826 B.n498 B.n32 106.175
R827 B.n498 B.n497 106.175
R828 B.n497 B.n496 106.175
R829 B.n496 B.n36 106.175
R830 B.n490 B.n36 106.175
R831 B.n489 B.n488 106.175
R832 B.n488 B.n43 106.175
R833 B.n482 B.n43 106.175
R834 B.n482 B.n481 106.175
R835 B.n481 B.n480 106.175
R836 B.n480 B.n50 106.175
R837 B.n474 B.n50 106.175
R838 B.n473 B.n472 106.175
R839 B.n472 B.n57 106.175
R840 B.n466 B.n57 106.175
R841 B.n466 B.n465 106.175
R842 B.n465 B.n464 106.175
R843 B.n464 B.n64 106.175
R844 B.n370 B.t5 104.614
R845 B.n504 B.t2 104.614
R846 B.n327 B.t9 95.2454
R847 B.n474 B.t13 95.2454
R848 B.n160 B.t3 76.5087
R849 B.t7 B.n521 76.5087
R850 B.n304 B.n303 71.676
R851 B.n234 B.n219 71.676
R852 B.n296 B.n220 71.676
R853 B.n292 B.n221 71.676
R854 B.n288 B.n222 71.676
R855 B.n284 B.n223 71.676
R856 B.n279 B.n224 71.676
R857 B.n275 B.n225 71.676
R858 B.n271 B.n226 71.676
R859 B.n267 B.n227 71.676
R860 B.n263 B.n228 71.676
R861 B.n259 B.n229 71.676
R862 B.n255 B.n230 71.676
R863 B.n251 B.n231 71.676
R864 B.n247 B.n232 71.676
R865 B.n243 B.n233 71.676
R866 B.n459 B.n458 71.676
R867 B.n90 B.n68 71.676
R868 B.n94 B.n69 71.676
R869 B.n98 B.n70 71.676
R870 B.n102 B.n71 71.676
R871 B.n106 B.n72 71.676
R872 B.n110 B.n73 71.676
R873 B.n114 B.n74 71.676
R874 B.n118 B.n75 71.676
R875 B.n122 B.n76 71.676
R876 B.n126 B.n77 71.676
R877 B.n131 B.n78 71.676
R878 B.n135 B.n79 71.676
R879 B.n139 B.n80 71.676
R880 B.n143 B.n81 71.676
R881 B.n147 B.n82 71.676
R882 B.n83 B.n82 71.676
R883 B.n146 B.n81 71.676
R884 B.n142 B.n80 71.676
R885 B.n138 B.n79 71.676
R886 B.n134 B.n78 71.676
R887 B.n130 B.n77 71.676
R888 B.n125 B.n76 71.676
R889 B.n121 B.n75 71.676
R890 B.n117 B.n74 71.676
R891 B.n113 B.n73 71.676
R892 B.n109 B.n72 71.676
R893 B.n105 B.n71 71.676
R894 B.n101 B.n70 71.676
R895 B.n97 B.n69 71.676
R896 B.n93 B.n68 71.676
R897 B.n458 B.n67 71.676
R898 B.n303 B.n218 71.676
R899 B.n297 B.n219 71.676
R900 B.n293 B.n220 71.676
R901 B.n289 B.n221 71.676
R902 B.n285 B.n222 71.676
R903 B.n280 B.n223 71.676
R904 B.n276 B.n224 71.676
R905 B.n272 B.n225 71.676
R906 B.n268 B.n226 71.676
R907 B.n264 B.n227 71.676
R908 B.n260 B.n228 71.676
R909 B.n256 B.n229 71.676
R910 B.n252 B.n230 71.676
R911 B.n248 B.n231 71.676
R912 B.n244 B.n232 71.676
R913 B.n240 B.n233 71.676
R914 B.n191 B.t4 70.2631
R915 B.t1 B.n489 70.2631
R916 B.t0 B.n164 67.1403
R917 B.n513 B.t6 67.1403
R918 B.n239 B.n238 59.5399
R919 B.n282 B.n236 59.5399
R920 B.n89 B.n88 59.5399
R921 B.n128 B.n86 59.5399
R922 B.n382 B.t0 39.0353
R923 B.t6 B.n512 39.0353
R924 B.n351 B.t4 35.9125
R925 B.n490 B.t1 35.9125
R926 B.n238 B.n237 35.2975
R927 B.n236 B.n235 35.2975
R928 B.n88 B.n87 35.2975
R929 B.n86 B.n85 35.2975
R930 B.n401 B.t3 29.6669
R931 B.n522 B.t7 29.6669
R932 B.n461 B.n460 29.1907
R933 B.n455 B.n454 29.1907
R934 B.n241 B.n213 29.1907
R935 B.n306 B.n305 29.1907
R936 B B.n532 18.0485
R937 B.n207 B.t9 10.9302
R938 B.t13 B.n473 10.9302
R939 B.n460 B.n66 10.6151
R940 B.n91 B.n66 10.6151
R941 B.n92 B.n91 10.6151
R942 B.n95 B.n92 10.6151
R943 B.n96 B.n95 10.6151
R944 B.n99 B.n96 10.6151
R945 B.n100 B.n99 10.6151
R946 B.n103 B.n100 10.6151
R947 B.n104 B.n103 10.6151
R948 B.n107 B.n104 10.6151
R949 B.n108 B.n107 10.6151
R950 B.n112 B.n111 10.6151
R951 B.n115 B.n112 10.6151
R952 B.n116 B.n115 10.6151
R953 B.n119 B.n116 10.6151
R954 B.n120 B.n119 10.6151
R955 B.n123 B.n120 10.6151
R956 B.n124 B.n123 10.6151
R957 B.n127 B.n124 10.6151
R958 B.n132 B.n129 10.6151
R959 B.n133 B.n132 10.6151
R960 B.n136 B.n133 10.6151
R961 B.n137 B.n136 10.6151
R962 B.n140 B.n137 10.6151
R963 B.n141 B.n140 10.6151
R964 B.n144 B.n141 10.6151
R965 B.n145 B.n144 10.6151
R966 B.n148 B.n145 10.6151
R967 B.n149 B.n148 10.6151
R968 B.n455 B.n149 10.6151
R969 B.n311 B.n213 10.6151
R970 B.n312 B.n311 10.6151
R971 B.n313 B.n312 10.6151
R972 B.n313 B.n204 10.6151
R973 B.n323 B.n204 10.6151
R974 B.n324 B.n323 10.6151
R975 B.n325 B.n324 10.6151
R976 B.n325 B.n197 10.6151
R977 B.n335 B.n197 10.6151
R978 B.n336 B.n335 10.6151
R979 B.n337 B.n336 10.6151
R980 B.n337 B.n188 10.6151
R981 B.n347 B.n188 10.6151
R982 B.n348 B.n347 10.6151
R983 B.n349 B.n348 10.6151
R984 B.n349 B.n181 10.6151
R985 B.n359 B.n181 10.6151
R986 B.n360 B.n359 10.6151
R987 B.n361 B.n360 10.6151
R988 B.n361 B.n174 10.6151
R989 B.n372 B.n174 10.6151
R990 B.n373 B.n372 10.6151
R991 B.n374 B.n373 10.6151
R992 B.n374 B.n166 10.6151
R993 B.n384 B.n166 10.6151
R994 B.n385 B.n384 10.6151
R995 B.n386 B.n385 10.6151
R996 B.n386 B.n157 10.6151
R997 B.n396 B.n157 10.6151
R998 B.n397 B.n396 10.6151
R999 B.n399 B.n397 10.6151
R1000 B.n399 B.n398 10.6151
R1001 B.n398 B.n150 10.6151
R1002 B.n410 B.n150 10.6151
R1003 B.n411 B.n410 10.6151
R1004 B.n412 B.n411 10.6151
R1005 B.n413 B.n412 10.6151
R1006 B.n415 B.n413 10.6151
R1007 B.n416 B.n415 10.6151
R1008 B.n417 B.n416 10.6151
R1009 B.n418 B.n417 10.6151
R1010 B.n420 B.n418 10.6151
R1011 B.n421 B.n420 10.6151
R1012 B.n422 B.n421 10.6151
R1013 B.n423 B.n422 10.6151
R1014 B.n425 B.n423 10.6151
R1015 B.n426 B.n425 10.6151
R1016 B.n427 B.n426 10.6151
R1017 B.n428 B.n427 10.6151
R1018 B.n430 B.n428 10.6151
R1019 B.n431 B.n430 10.6151
R1020 B.n432 B.n431 10.6151
R1021 B.n433 B.n432 10.6151
R1022 B.n435 B.n433 10.6151
R1023 B.n436 B.n435 10.6151
R1024 B.n437 B.n436 10.6151
R1025 B.n438 B.n437 10.6151
R1026 B.n440 B.n438 10.6151
R1027 B.n441 B.n440 10.6151
R1028 B.n442 B.n441 10.6151
R1029 B.n443 B.n442 10.6151
R1030 B.n445 B.n443 10.6151
R1031 B.n446 B.n445 10.6151
R1032 B.n447 B.n446 10.6151
R1033 B.n448 B.n447 10.6151
R1034 B.n450 B.n448 10.6151
R1035 B.n451 B.n450 10.6151
R1036 B.n452 B.n451 10.6151
R1037 B.n453 B.n452 10.6151
R1038 B.n454 B.n453 10.6151
R1039 B.n305 B.n217 10.6151
R1040 B.n300 B.n217 10.6151
R1041 B.n300 B.n299 10.6151
R1042 B.n299 B.n298 10.6151
R1043 B.n298 B.n295 10.6151
R1044 B.n295 B.n294 10.6151
R1045 B.n294 B.n291 10.6151
R1046 B.n291 B.n290 10.6151
R1047 B.n290 B.n287 10.6151
R1048 B.n287 B.n286 10.6151
R1049 B.n286 B.n283 10.6151
R1050 B.n281 B.n278 10.6151
R1051 B.n278 B.n277 10.6151
R1052 B.n277 B.n274 10.6151
R1053 B.n274 B.n273 10.6151
R1054 B.n273 B.n270 10.6151
R1055 B.n270 B.n269 10.6151
R1056 B.n269 B.n266 10.6151
R1057 B.n266 B.n265 10.6151
R1058 B.n262 B.n261 10.6151
R1059 B.n261 B.n258 10.6151
R1060 B.n258 B.n257 10.6151
R1061 B.n257 B.n254 10.6151
R1062 B.n254 B.n253 10.6151
R1063 B.n253 B.n250 10.6151
R1064 B.n250 B.n249 10.6151
R1065 B.n249 B.n246 10.6151
R1066 B.n246 B.n245 10.6151
R1067 B.n245 B.n242 10.6151
R1068 B.n242 B.n241 10.6151
R1069 B.n307 B.n306 10.6151
R1070 B.n307 B.n209 10.6151
R1071 B.n317 B.n209 10.6151
R1072 B.n318 B.n317 10.6151
R1073 B.n319 B.n318 10.6151
R1074 B.n319 B.n201 10.6151
R1075 B.n329 B.n201 10.6151
R1076 B.n330 B.n329 10.6151
R1077 B.n331 B.n330 10.6151
R1078 B.n331 B.n193 10.6151
R1079 B.n341 B.n193 10.6151
R1080 B.n342 B.n341 10.6151
R1081 B.n343 B.n342 10.6151
R1082 B.n343 B.n185 10.6151
R1083 B.n353 B.n185 10.6151
R1084 B.n354 B.n353 10.6151
R1085 B.n355 B.n354 10.6151
R1086 B.n355 B.n177 10.6151
R1087 B.n366 B.n177 10.6151
R1088 B.n367 B.n366 10.6151
R1089 B.n368 B.n367 10.6151
R1090 B.n368 B.n170 10.6151
R1091 B.n378 B.n170 10.6151
R1092 B.n379 B.n378 10.6151
R1093 B.n380 B.n379 10.6151
R1094 B.n380 B.n162 10.6151
R1095 B.n390 B.n162 10.6151
R1096 B.n391 B.n390 10.6151
R1097 B.n392 B.n391 10.6151
R1098 B.n392 B.n154 10.6151
R1099 B.n403 B.n154 10.6151
R1100 B.n404 B.n403 10.6151
R1101 B.n405 B.n404 10.6151
R1102 B.n405 B.n0 10.6151
R1103 B.n526 B.n1 10.6151
R1104 B.n526 B.n525 10.6151
R1105 B.n525 B.n524 10.6151
R1106 B.n524 B.n10 10.6151
R1107 B.n518 B.n10 10.6151
R1108 B.n518 B.n517 10.6151
R1109 B.n517 B.n516 10.6151
R1110 B.n516 B.n17 10.6151
R1111 B.n510 B.n17 10.6151
R1112 B.n510 B.n509 10.6151
R1113 B.n509 B.n508 10.6151
R1114 B.n508 B.n24 10.6151
R1115 B.n502 B.n24 10.6151
R1116 B.n502 B.n501 10.6151
R1117 B.n501 B.n500 10.6151
R1118 B.n500 B.n30 10.6151
R1119 B.n494 B.n30 10.6151
R1120 B.n494 B.n493 10.6151
R1121 B.n493 B.n492 10.6151
R1122 B.n492 B.n38 10.6151
R1123 B.n486 B.n38 10.6151
R1124 B.n486 B.n485 10.6151
R1125 B.n485 B.n484 10.6151
R1126 B.n484 B.n45 10.6151
R1127 B.n478 B.n45 10.6151
R1128 B.n478 B.n477 10.6151
R1129 B.n477 B.n476 10.6151
R1130 B.n476 B.n52 10.6151
R1131 B.n470 B.n52 10.6151
R1132 B.n470 B.n469 10.6151
R1133 B.n469 B.n468 10.6151
R1134 B.n468 B.n59 10.6151
R1135 B.n462 B.n59 10.6151
R1136 B.n462 B.n461 10.6151
R1137 B.n111 B.n89 6.5566
R1138 B.n128 B.n127 6.5566
R1139 B.n282 B.n281 6.5566
R1140 B.n265 B.n239 6.5566
R1141 B.n108 B.n89 4.05904
R1142 B.n129 B.n128 4.05904
R1143 B.n283 B.n282 4.05904
R1144 B.n262 B.n239 4.05904
R1145 B.n532 B.n0 2.81026
R1146 B.n532 B.n1 2.81026
R1147 B.n363 B.t5 1.56189
R1148 B.n32 B.t2 1.56189
R1149 VN.n18 VN.n17 174.512
R1150 VN.n37 VN.n36 174.512
R1151 VN.n35 VN.n19 161.3
R1152 VN.n34 VN.n33 161.3
R1153 VN.n32 VN.n20 161.3
R1154 VN.n31 VN.n30 161.3
R1155 VN.n28 VN.n21 161.3
R1156 VN.n27 VN.n26 161.3
R1157 VN.n25 VN.n22 161.3
R1158 VN.n16 VN.n0 161.3
R1159 VN.n15 VN.n14 161.3
R1160 VN.n13 VN.n1 161.3
R1161 VN.n12 VN.n11 161.3
R1162 VN.n9 VN.n2 161.3
R1163 VN.n8 VN.n7 161.3
R1164 VN.n6 VN.n3 161.3
R1165 VN.n5 VN.t7 63.006
R1166 VN.n24 VN.t5 63.006
R1167 VN.n15 VN.n1 56.5193
R1168 VN.n34 VN.n20 56.5193
R1169 VN.n5 VN.n4 46.4328
R1170 VN.n24 VN.n23 46.4328
R1171 VN.n8 VN.n3 40.4934
R1172 VN.n9 VN.n8 40.4934
R1173 VN.n27 VN.n22 40.4934
R1174 VN.n28 VN.n27 40.4934
R1175 VN VN.n37 38.2751
R1176 VN.n4 VN.t3 28.6294
R1177 VN.n10 VN.t6 28.6294
R1178 VN.n17 VN.t2 28.6294
R1179 VN.n23 VN.t1 28.6294
R1180 VN.n29 VN.t4 28.6294
R1181 VN.n36 VN.t0 28.6294
R1182 VN.n11 VN.n1 24.4675
R1183 VN.n16 VN.n15 24.4675
R1184 VN.n30 VN.n20 24.4675
R1185 VN.n35 VN.n34 24.4675
R1186 VN.n4 VN.n3 20.0634
R1187 VN.n10 VN.n9 20.0634
R1188 VN.n23 VN.n22 20.0634
R1189 VN.n29 VN.n28 20.0634
R1190 VN.n25 VN.n24 17.6611
R1191 VN.n6 VN.n5 17.6611
R1192 VN.n17 VN.n16 11.2553
R1193 VN.n36 VN.n35 11.2553
R1194 VN.n11 VN.n10 4.40456
R1195 VN.n30 VN.n29 4.40456
R1196 VN.n37 VN.n19 0.189894
R1197 VN.n33 VN.n19 0.189894
R1198 VN.n33 VN.n32 0.189894
R1199 VN.n32 VN.n31 0.189894
R1200 VN.n31 VN.n21 0.189894
R1201 VN.n26 VN.n21 0.189894
R1202 VN.n26 VN.n25 0.189894
R1203 VN.n7 VN.n6 0.189894
R1204 VN.n7 VN.n2 0.189894
R1205 VN.n12 VN.n2 0.189894
R1206 VN.n13 VN.n12 0.189894
R1207 VN.n14 VN.n13 0.189894
R1208 VN.n14 VN.n0 0.189894
R1209 VN.n18 VN.n0 0.189894
R1210 VN VN.n18 0.0516364
R1211 VDD2.n2 VDD2.n1 101.959
R1212 VDD2.n2 VDD2.n0 101.959
R1213 VDD2 VDD2.n5 101.956
R1214 VDD2.n4 VDD2.n3 101.23
R1215 VDD2.n4 VDD2.n2 32.3015
R1216 VDD2.n5 VDD2.t6 11.1869
R1217 VDD2.n5 VDD2.t2 11.1869
R1218 VDD2.n3 VDD2.t7 11.1869
R1219 VDD2.n3 VDD2.t3 11.1869
R1220 VDD2.n1 VDD2.t1 11.1869
R1221 VDD2.n1 VDD2.t5 11.1869
R1222 VDD2.n0 VDD2.t0 11.1869
R1223 VDD2.n0 VDD2.t4 11.1869
R1224 VDD2 VDD2.n4 0.843172
C0 VP VTAIL 2.14137f
C1 VDD1 VTAIL 3.72735f
C2 VN VTAIL 2.12727f
C3 VTAIL VDD2 3.77433f
C4 VDD1 VP 1.72117f
C5 VN VP 4.41755f
C6 VP VDD2 0.408728f
C7 VDD1 VN 0.155867f
C8 VDD1 VDD2 1.21811f
C9 VN VDD2 1.47032f
C10 VDD2 B 3.285504f
C11 VDD1 B 3.582834f
C12 VTAIL B 3.339865f
C13 VN B 10.06709f
C14 VP B 8.819691f
C15 VDD2.t0 B 0.024813f
C16 VDD2.t4 B 0.024813f
C17 VDD2.n0 B 0.160582f
C18 VDD2.t1 B 0.024813f
C19 VDD2.t5 B 0.024813f
C20 VDD2.n1 B 0.160582f
C21 VDD2.n2 B 1.39081f
C22 VDD2.t7 B 0.024813f
C23 VDD2.t3 B 0.024813f
C24 VDD2.n3 B 0.158712f
C25 VDD2.n4 B 1.22153f
C26 VDD2.t6 B 0.024813f
C27 VDD2.t2 B 0.024813f
C28 VDD2.n5 B 0.16057f
C29 VN.n0 B 0.03086f
C30 VN.t2 B 0.18513f
C31 VN.n1 B 0.051069f
C32 VN.n2 B 0.03086f
C33 VN.t6 B 0.18513f
C34 VN.n3 B 0.056222f
C35 VN.t7 B 0.307366f
C36 VN.t3 B 0.18513f
C37 VN.n4 B 0.170962f
C38 VN.n5 B 0.150231f
C39 VN.n6 B 0.195659f
C40 VN.n7 B 0.03086f
C41 VN.n8 B 0.024947f
C42 VN.n9 B 0.056222f
C43 VN.n10 B 0.104423f
C44 VN.n11 B 0.034231f
C45 VN.n12 B 0.03086f
C46 VN.n13 B 0.03086f
C47 VN.n14 B 0.03086f
C48 VN.n15 B 0.03903f
C49 VN.n16 B 0.042181f
C50 VN.n17 B 0.169132f
C51 VN.n18 B 0.029215f
C52 VN.n19 B 0.03086f
C53 VN.t0 B 0.18513f
C54 VN.n20 B 0.051069f
C55 VN.n21 B 0.03086f
C56 VN.t4 B 0.18513f
C57 VN.n22 B 0.056222f
C58 VN.t5 B 0.307366f
C59 VN.t1 B 0.18513f
C60 VN.n23 B 0.170962f
C61 VN.n24 B 0.150231f
C62 VN.n25 B 0.195659f
C63 VN.n26 B 0.03086f
C64 VN.n27 B 0.024947f
C65 VN.n28 B 0.056222f
C66 VN.n29 B 0.104423f
C67 VN.n30 B 0.034231f
C68 VN.n31 B 0.03086f
C69 VN.n32 B 0.03086f
C70 VN.n33 B 0.03086f
C71 VN.n34 B 0.03903f
C72 VN.n35 B 0.042181f
C73 VN.n36 B 0.169132f
C74 VN.n37 B 1.09184f
C75 VTAIL.t6 B 0.041241f
C76 VTAIL.t2 B 0.041241f
C77 VTAIL.n0 B 0.224724f
C78 VTAIL.n1 B 0.357238f
C79 VTAIL.n2 B 0.03846f
C80 VTAIL.n3 B 0.090116f
C81 VTAIL.t7 B 0.064748f
C82 VTAIL.n4 B 0.066433f
C83 VTAIL.n5 B 0.019519f
C84 VTAIL.n6 B 0.015844f
C85 VTAIL.n7 B 0.175516f
C86 VTAIL.n8 B 0.041977f
C87 VTAIL.n9 B 0.220934f
C88 VTAIL.n10 B 0.03846f
C89 VTAIL.n11 B 0.090116f
C90 VTAIL.t13 B 0.064748f
C91 VTAIL.n12 B 0.066433f
C92 VTAIL.n13 B 0.019519f
C93 VTAIL.n14 B 0.015844f
C94 VTAIL.n15 B 0.175516f
C95 VTAIL.n16 B 0.041977f
C96 VTAIL.n17 B 0.220934f
C97 VTAIL.t14 B 0.041241f
C98 VTAIL.t10 B 0.041241f
C99 VTAIL.n18 B 0.224724f
C100 VTAIL.n19 B 0.500775f
C101 VTAIL.n20 B 0.03846f
C102 VTAIL.n21 B 0.090116f
C103 VTAIL.t12 B 0.064748f
C104 VTAIL.n22 B 0.066433f
C105 VTAIL.n23 B 0.019519f
C106 VTAIL.n24 B 0.015844f
C107 VTAIL.n25 B 0.175516f
C108 VTAIL.n26 B 0.041977f
C109 VTAIL.n27 B 0.870856f
C110 VTAIL.n28 B 0.03846f
C111 VTAIL.n29 B 0.090116f
C112 VTAIL.t4 B 0.064748f
C113 VTAIL.n30 B 0.066433f
C114 VTAIL.n31 B 0.019519f
C115 VTAIL.n32 B 0.015844f
C116 VTAIL.n33 B 0.175516f
C117 VTAIL.n34 B 0.041977f
C118 VTAIL.n35 B 0.870855f
C119 VTAIL.t5 B 0.041241f
C120 VTAIL.t0 B 0.041241f
C121 VTAIL.n36 B 0.224726f
C122 VTAIL.n37 B 0.500773f
C123 VTAIL.n38 B 0.03846f
C124 VTAIL.n39 B 0.090116f
C125 VTAIL.t3 B 0.064748f
C126 VTAIL.n40 B 0.066433f
C127 VTAIL.n41 B 0.019519f
C128 VTAIL.n42 B 0.015844f
C129 VTAIL.n43 B 0.175516f
C130 VTAIL.n44 B 0.041977f
C131 VTAIL.n45 B 0.220934f
C132 VTAIL.n46 B 0.03846f
C133 VTAIL.n47 B 0.090116f
C134 VTAIL.t11 B 0.064748f
C135 VTAIL.n48 B 0.066433f
C136 VTAIL.n49 B 0.019519f
C137 VTAIL.n50 B 0.015844f
C138 VTAIL.n51 B 0.175516f
C139 VTAIL.n52 B 0.041977f
C140 VTAIL.n53 B 0.220934f
C141 VTAIL.t8 B 0.041241f
C142 VTAIL.t15 B 0.041241f
C143 VTAIL.n54 B 0.224726f
C144 VTAIL.n55 B 0.500773f
C145 VTAIL.n56 B 0.03846f
C146 VTAIL.n57 B 0.090116f
C147 VTAIL.t9 B 0.064748f
C148 VTAIL.n58 B 0.066433f
C149 VTAIL.n59 B 0.019519f
C150 VTAIL.n60 B 0.015844f
C151 VTAIL.n61 B 0.175516f
C152 VTAIL.n62 B 0.041977f
C153 VTAIL.n63 B 0.870856f
C154 VTAIL.n64 B 0.03846f
C155 VTAIL.n65 B 0.090116f
C156 VTAIL.t1 B 0.064748f
C157 VTAIL.n66 B 0.066433f
C158 VTAIL.n67 B 0.019519f
C159 VTAIL.n68 B 0.015844f
C160 VTAIL.n69 B 0.175516f
C161 VTAIL.n70 B 0.041977f
C162 VTAIL.n71 B 0.865327f
C163 VDD1.t7 B 0.023751f
C164 VDD1.t2 B 0.023751f
C165 VDD1.n0 B 0.15403f
C166 VDD1.t5 B 0.023751f
C167 VDD1.t1 B 0.023751f
C168 VDD1.n1 B 0.153706f
C169 VDD1.t3 B 0.023751f
C170 VDD1.t6 B 0.023751f
C171 VDD1.n2 B 0.153706f
C172 VDD1.n3 B 1.36724f
C173 VDD1.t4 B 0.023751f
C174 VDD1.t0 B 0.023751f
C175 VDD1.n4 B 0.151916f
C176 VDD1.n5 B 1.18959f
C177 VP.n0 B 0.031067f
C178 VP.t2 B 0.186374f
C179 VP.n1 B 0.051412f
C180 VP.n2 B 0.031067f
C181 VP.t5 B 0.186374f
C182 VP.n3 B 0.0566f
C183 VP.n4 B 0.031067f
C184 VP.n5 B 0.042465f
C185 VP.n6 B 0.031067f
C186 VP.t6 B 0.186374f
C187 VP.n7 B 0.051412f
C188 VP.n8 B 0.031067f
C189 VP.t0 B 0.186374f
C190 VP.n9 B 0.0566f
C191 VP.t4 B 0.309431f
C192 VP.t7 B 0.186374f
C193 VP.n10 B 0.17211f
C194 VP.n11 B 0.151241f
C195 VP.n12 B 0.196974f
C196 VP.n13 B 0.031067f
C197 VP.n14 B 0.025115f
C198 VP.n15 B 0.0566f
C199 VP.n16 B 0.105125f
C200 VP.n17 B 0.034461f
C201 VP.n18 B 0.031067f
C202 VP.n19 B 0.031067f
C203 VP.n20 B 0.031067f
C204 VP.n21 B 0.039292f
C205 VP.n22 B 0.042465f
C206 VP.n23 B 0.170268f
C207 VP.n24 B 1.07865f
C208 VP.t3 B 0.186374f
C209 VP.n25 B 0.170268f
C210 VP.n26 B 1.10812f
C211 VP.n27 B 0.031067f
C212 VP.n28 B 0.031067f
C213 VP.n29 B 0.039292f
C214 VP.n30 B 0.051412f
C215 VP.t1 B 0.186374f
C216 VP.n31 B 0.105125f
C217 VP.n32 B 0.034461f
C218 VP.n33 B 0.031067f
C219 VP.n34 B 0.031067f
C220 VP.n35 B 0.031067f
C221 VP.n36 B 0.025115f
C222 VP.n37 B 0.0566f
C223 VP.n38 B 0.105125f
C224 VP.n39 B 0.034461f
C225 VP.n40 B 0.031067f
C226 VP.n41 B 0.031067f
C227 VP.n42 B 0.031067f
C228 VP.n43 B 0.039292f
C229 VP.n44 B 0.042465f
C230 VP.n45 B 0.170268f
C231 VP.n46 B 0.029412f
.ends

