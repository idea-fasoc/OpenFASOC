* NGSPICE file created from diff_pair_sample_0596.ext - technology: sky130A

.subckt diff_pair_sample_0596 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=0 ps=0 w=7.21 l=3.38
X1 VTAIL.t7 VP.t0 VDD1.t0 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=1.18965 ps=7.54 w=7.21 l=3.38
X2 VDD1.t3 VP.t1 VTAIL.t6 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=1.18965 pd=7.54 as=2.8119 ps=15.2 w=7.21 l=3.38
X3 B.t8 B.t6 B.t7 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=0 ps=0 w=7.21 l=3.38
X4 VDD2.t3 VN.t0 VTAIL.t3 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=1.18965 pd=7.54 as=2.8119 ps=15.2 w=7.21 l=3.38
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=1.18965 pd=7.54 as=2.8119 ps=15.2 w=7.21 l=3.38
X6 VTAIL.t1 VN.t2 VDD2.t1 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=1.18965 ps=7.54 w=7.21 l=3.38
X7 B.t5 B.t3 B.t4 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=0 ps=0 w=7.21 l=3.38
X8 VTAIL.t2 VN.t3 VDD2.t0 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=1.18965 ps=7.54 w=7.21 l=3.38
X9 VTAIL.t5 VP.t2 VDD1.t1 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=1.18965 ps=7.54 w=7.21 l=3.38
X10 B.t2 B.t0 B.t1 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=2.8119 pd=15.2 as=0 ps=0 w=7.21 l=3.38
X11 VDD1.t2 VP.t3 VTAIL.t4 w_n3196_n2410# sky130_fd_pr__pfet_01v8 ad=1.18965 pd=7.54 as=2.8119 ps=15.2 w=7.21 l=3.38
R0 B.n443 B.n442 585
R1 B.n444 B.n59 585
R2 B.n446 B.n445 585
R3 B.n447 B.n58 585
R4 B.n449 B.n448 585
R5 B.n450 B.n57 585
R6 B.n452 B.n451 585
R7 B.n453 B.n56 585
R8 B.n455 B.n454 585
R9 B.n456 B.n55 585
R10 B.n458 B.n457 585
R11 B.n459 B.n54 585
R12 B.n461 B.n460 585
R13 B.n462 B.n53 585
R14 B.n464 B.n463 585
R15 B.n465 B.n52 585
R16 B.n467 B.n466 585
R17 B.n468 B.n51 585
R18 B.n470 B.n469 585
R19 B.n471 B.n50 585
R20 B.n473 B.n472 585
R21 B.n474 B.n49 585
R22 B.n476 B.n475 585
R23 B.n477 B.n48 585
R24 B.n479 B.n478 585
R25 B.n480 B.n47 585
R26 B.n482 B.n481 585
R27 B.n483 B.n44 585
R28 B.n486 B.n485 585
R29 B.n487 B.n43 585
R30 B.n489 B.n488 585
R31 B.n490 B.n42 585
R32 B.n492 B.n491 585
R33 B.n493 B.n41 585
R34 B.n495 B.n494 585
R35 B.n496 B.n37 585
R36 B.n498 B.n497 585
R37 B.n499 B.n36 585
R38 B.n501 B.n500 585
R39 B.n502 B.n35 585
R40 B.n504 B.n503 585
R41 B.n505 B.n34 585
R42 B.n507 B.n506 585
R43 B.n508 B.n33 585
R44 B.n510 B.n509 585
R45 B.n511 B.n32 585
R46 B.n513 B.n512 585
R47 B.n514 B.n31 585
R48 B.n516 B.n515 585
R49 B.n517 B.n30 585
R50 B.n519 B.n518 585
R51 B.n520 B.n29 585
R52 B.n522 B.n521 585
R53 B.n523 B.n28 585
R54 B.n525 B.n524 585
R55 B.n526 B.n27 585
R56 B.n528 B.n527 585
R57 B.n529 B.n26 585
R58 B.n531 B.n530 585
R59 B.n532 B.n25 585
R60 B.n534 B.n533 585
R61 B.n535 B.n24 585
R62 B.n537 B.n536 585
R63 B.n538 B.n23 585
R64 B.n540 B.n539 585
R65 B.n441 B.n60 585
R66 B.n440 B.n439 585
R67 B.n438 B.n61 585
R68 B.n437 B.n436 585
R69 B.n435 B.n62 585
R70 B.n434 B.n433 585
R71 B.n432 B.n63 585
R72 B.n431 B.n430 585
R73 B.n429 B.n64 585
R74 B.n428 B.n427 585
R75 B.n426 B.n65 585
R76 B.n425 B.n424 585
R77 B.n423 B.n66 585
R78 B.n422 B.n421 585
R79 B.n420 B.n67 585
R80 B.n419 B.n418 585
R81 B.n417 B.n68 585
R82 B.n416 B.n415 585
R83 B.n414 B.n69 585
R84 B.n413 B.n412 585
R85 B.n411 B.n70 585
R86 B.n410 B.n409 585
R87 B.n408 B.n71 585
R88 B.n407 B.n406 585
R89 B.n405 B.n72 585
R90 B.n404 B.n403 585
R91 B.n402 B.n73 585
R92 B.n401 B.n400 585
R93 B.n399 B.n74 585
R94 B.n398 B.n397 585
R95 B.n396 B.n75 585
R96 B.n395 B.n394 585
R97 B.n393 B.n76 585
R98 B.n392 B.n391 585
R99 B.n390 B.n77 585
R100 B.n389 B.n388 585
R101 B.n387 B.n78 585
R102 B.n386 B.n385 585
R103 B.n384 B.n79 585
R104 B.n383 B.n382 585
R105 B.n381 B.n80 585
R106 B.n380 B.n379 585
R107 B.n378 B.n81 585
R108 B.n377 B.n376 585
R109 B.n375 B.n82 585
R110 B.n374 B.n373 585
R111 B.n372 B.n83 585
R112 B.n371 B.n370 585
R113 B.n369 B.n84 585
R114 B.n368 B.n367 585
R115 B.n366 B.n85 585
R116 B.n365 B.n364 585
R117 B.n363 B.n86 585
R118 B.n362 B.n361 585
R119 B.n360 B.n87 585
R120 B.n359 B.n358 585
R121 B.n357 B.n88 585
R122 B.n356 B.n355 585
R123 B.n354 B.n89 585
R124 B.n353 B.n352 585
R125 B.n351 B.n90 585
R126 B.n350 B.n349 585
R127 B.n348 B.n91 585
R128 B.n347 B.n346 585
R129 B.n345 B.n92 585
R130 B.n344 B.n343 585
R131 B.n342 B.n93 585
R132 B.n341 B.n340 585
R133 B.n339 B.n94 585
R134 B.n338 B.n337 585
R135 B.n336 B.n95 585
R136 B.n335 B.n334 585
R137 B.n333 B.n96 585
R138 B.n332 B.n331 585
R139 B.n330 B.n97 585
R140 B.n329 B.n328 585
R141 B.n327 B.n98 585
R142 B.n326 B.n325 585
R143 B.n324 B.n99 585
R144 B.n323 B.n322 585
R145 B.n321 B.n100 585
R146 B.n320 B.n319 585
R147 B.n318 B.n101 585
R148 B.n217 B.n216 585
R149 B.n218 B.n135 585
R150 B.n220 B.n219 585
R151 B.n221 B.n134 585
R152 B.n223 B.n222 585
R153 B.n224 B.n133 585
R154 B.n226 B.n225 585
R155 B.n227 B.n132 585
R156 B.n229 B.n228 585
R157 B.n230 B.n131 585
R158 B.n232 B.n231 585
R159 B.n233 B.n130 585
R160 B.n235 B.n234 585
R161 B.n236 B.n129 585
R162 B.n238 B.n237 585
R163 B.n239 B.n128 585
R164 B.n241 B.n240 585
R165 B.n242 B.n127 585
R166 B.n244 B.n243 585
R167 B.n245 B.n126 585
R168 B.n247 B.n246 585
R169 B.n248 B.n125 585
R170 B.n250 B.n249 585
R171 B.n251 B.n124 585
R172 B.n253 B.n252 585
R173 B.n254 B.n123 585
R174 B.n256 B.n255 585
R175 B.n257 B.n120 585
R176 B.n260 B.n259 585
R177 B.n261 B.n119 585
R178 B.n263 B.n262 585
R179 B.n264 B.n118 585
R180 B.n266 B.n265 585
R181 B.n267 B.n117 585
R182 B.n269 B.n268 585
R183 B.n270 B.n116 585
R184 B.n275 B.n274 585
R185 B.n276 B.n115 585
R186 B.n278 B.n277 585
R187 B.n279 B.n114 585
R188 B.n281 B.n280 585
R189 B.n282 B.n113 585
R190 B.n284 B.n283 585
R191 B.n285 B.n112 585
R192 B.n287 B.n286 585
R193 B.n288 B.n111 585
R194 B.n290 B.n289 585
R195 B.n291 B.n110 585
R196 B.n293 B.n292 585
R197 B.n294 B.n109 585
R198 B.n296 B.n295 585
R199 B.n297 B.n108 585
R200 B.n299 B.n298 585
R201 B.n300 B.n107 585
R202 B.n302 B.n301 585
R203 B.n303 B.n106 585
R204 B.n305 B.n304 585
R205 B.n306 B.n105 585
R206 B.n308 B.n307 585
R207 B.n309 B.n104 585
R208 B.n311 B.n310 585
R209 B.n312 B.n103 585
R210 B.n314 B.n313 585
R211 B.n315 B.n102 585
R212 B.n317 B.n316 585
R213 B.n215 B.n136 585
R214 B.n214 B.n213 585
R215 B.n212 B.n137 585
R216 B.n211 B.n210 585
R217 B.n209 B.n138 585
R218 B.n208 B.n207 585
R219 B.n206 B.n139 585
R220 B.n205 B.n204 585
R221 B.n203 B.n140 585
R222 B.n202 B.n201 585
R223 B.n200 B.n141 585
R224 B.n199 B.n198 585
R225 B.n197 B.n142 585
R226 B.n196 B.n195 585
R227 B.n194 B.n143 585
R228 B.n193 B.n192 585
R229 B.n191 B.n144 585
R230 B.n190 B.n189 585
R231 B.n188 B.n145 585
R232 B.n187 B.n186 585
R233 B.n185 B.n146 585
R234 B.n184 B.n183 585
R235 B.n182 B.n147 585
R236 B.n181 B.n180 585
R237 B.n179 B.n148 585
R238 B.n178 B.n177 585
R239 B.n176 B.n149 585
R240 B.n175 B.n174 585
R241 B.n173 B.n150 585
R242 B.n172 B.n171 585
R243 B.n170 B.n151 585
R244 B.n169 B.n168 585
R245 B.n167 B.n152 585
R246 B.n166 B.n165 585
R247 B.n164 B.n153 585
R248 B.n163 B.n162 585
R249 B.n161 B.n154 585
R250 B.n160 B.n159 585
R251 B.n158 B.n155 585
R252 B.n157 B.n156 585
R253 B.n2 B.n0 585
R254 B.n601 B.n1 585
R255 B.n600 B.n599 585
R256 B.n598 B.n3 585
R257 B.n597 B.n596 585
R258 B.n595 B.n4 585
R259 B.n594 B.n593 585
R260 B.n592 B.n5 585
R261 B.n591 B.n590 585
R262 B.n589 B.n6 585
R263 B.n588 B.n587 585
R264 B.n586 B.n7 585
R265 B.n585 B.n584 585
R266 B.n583 B.n8 585
R267 B.n582 B.n581 585
R268 B.n580 B.n9 585
R269 B.n579 B.n578 585
R270 B.n577 B.n10 585
R271 B.n576 B.n575 585
R272 B.n574 B.n11 585
R273 B.n573 B.n572 585
R274 B.n571 B.n12 585
R275 B.n570 B.n569 585
R276 B.n568 B.n13 585
R277 B.n567 B.n566 585
R278 B.n565 B.n14 585
R279 B.n564 B.n563 585
R280 B.n562 B.n15 585
R281 B.n561 B.n560 585
R282 B.n559 B.n16 585
R283 B.n558 B.n557 585
R284 B.n556 B.n17 585
R285 B.n555 B.n554 585
R286 B.n553 B.n18 585
R287 B.n552 B.n551 585
R288 B.n550 B.n19 585
R289 B.n549 B.n548 585
R290 B.n547 B.n20 585
R291 B.n546 B.n545 585
R292 B.n544 B.n21 585
R293 B.n543 B.n542 585
R294 B.n541 B.n22 585
R295 B.n603 B.n602 585
R296 B.n217 B.n136 444.452
R297 B.n541 B.n540 444.452
R298 B.n318 B.n317 444.452
R299 B.n443 B.n60 444.452
R300 B.n271 B.t5 361.337
R301 B.n45 B.t7 361.337
R302 B.n121 B.t2 361.337
R303 B.n38 B.t10 361.337
R304 B.n272 B.t4 289.387
R305 B.n46 B.t8 289.387
R306 B.n122 B.t1 289.387
R307 B.n39 B.t11 289.387
R308 B.n271 B.t3 260.392
R309 B.n121 B.t0 260.392
R310 B.n38 B.t9 260.392
R311 B.n45 B.t6 260.392
R312 B.n213 B.n136 163.367
R313 B.n213 B.n212 163.367
R314 B.n212 B.n211 163.367
R315 B.n211 B.n138 163.367
R316 B.n207 B.n138 163.367
R317 B.n207 B.n206 163.367
R318 B.n206 B.n205 163.367
R319 B.n205 B.n140 163.367
R320 B.n201 B.n140 163.367
R321 B.n201 B.n200 163.367
R322 B.n200 B.n199 163.367
R323 B.n199 B.n142 163.367
R324 B.n195 B.n142 163.367
R325 B.n195 B.n194 163.367
R326 B.n194 B.n193 163.367
R327 B.n193 B.n144 163.367
R328 B.n189 B.n144 163.367
R329 B.n189 B.n188 163.367
R330 B.n188 B.n187 163.367
R331 B.n187 B.n146 163.367
R332 B.n183 B.n146 163.367
R333 B.n183 B.n182 163.367
R334 B.n182 B.n181 163.367
R335 B.n181 B.n148 163.367
R336 B.n177 B.n148 163.367
R337 B.n177 B.n176 163.367
R338 B.n176 B.n175 163.367
R339 B.n175 B.n150 163.367
R340 B.n171 B.n150 163.367
R341 B.n171 B.n170 163.367
R342 B.n170 B.n169 163.367
R343 B.n169 B.n152 163.367
R344 B.n165 B.n152 163.367
R345 B.n165 B.n164 163.367
R346 B.n164 B.n163 163.367
R347 B.n163 B.n154 163.367
R348 B.n159 B.n154 163.367
R349 B.n159 B.n158 163.367
R350 B.n158 B.n157 163.367
R351 B.n157 B.n2 163.367
R352 B.n602 B.n2 163.367
R353 B.n602 B.n601 163.367
R354 B.n601 B.n600 163.367
R355 B.n600 B.n3 163.367
R356 B.n596 B.n3 163.367
R357 B.n596 B.n595 163.367
R358 B.n595 B.n594 163.367
R359 B.n594 B.n5 163.367
R360 B.n590 B.n5 163.367
R361 B.n590 B.n589 163.367
R362 B.n589 B.n588 163.367
R363 B.n588 B.n7 163.367
R364 B.n584 B.n7 163.367
R365 B.n584 B.n583 163.367
R366 B.n583 B.n582 163.367
R367 B.n582 B.n9 163.367
R368 B.n578 B.n9 163.367
R369 B.n578 B.n577 163.367
R370 B.n577 B.n576 163.367
R371 B.n576 B.n11 163.367
R372 B.n572 B.n11 163.367
R373 B.n572 B.n571 163.367
R374 B.n571 B.n570 163.367
R375 B.n570 B.n13 163.367
R376 B.n566 B.n13 163.367
R377 B.n566 B.n565 163.367
R378 B.n565 B.n564 163.367
R379 B.n564 B.n15 163.367
R380 B.n560 B.n15 163.367
R381 B.n560 B.n559 163.367
R382 B.n559 B.n558 163.367
R383 B.n558 B.n17 163.367
R384 B.n554 B.n17 163.367
R385 B.n554 B.n553 163.367
R386 B.n553 B.n552 163.367
R387 B.n552 B.n19 163.367
R388 B.n548 B.n19 163.367
R389 B.n548 B.n547 163.367
R390 B.n547 B.n546 163.367
R391 B.n546 B.n21 163.367
R392 B.n542 B.n21 163.367
R393 B.n542 B.n541 163.367
R394 B.n218 B.n217 163.367
R395 B.n219 B.n218 163.367
R396 B.n219 B.n134 163.367
R397 B.n223 B.n134 163.367
R398 B.n224 B.n223 163.367
R399 B.n225 B.n224 163.367
R400 B.n225 B.n132 163.367
R401 B.n229 B.n132 163.367
R402 B.n230 B.n229 163.367
R403 B.n231 B.n230 163.367
R404 B.n231 B.n130 163.367
R405 B.n235 B.n130 163.367
R406 B.n236 B.n235 163.367
R407 B.n237 B.n236 163.367
R408 B.n237 B.n128 163.367
R409 B.n241 B.n128 163.367
R410 B.n242 B.n241 163.367
R411 B.n243 B.n242 163.367
R412 B.n243 B.n126 163.367
R413 B.n247 B.n126 163.367
R414 B.n248 B.n247 163.367
R415 B.n249 B.n248 163.367
R416 B.n249 B.n124 163.367
R417 B.n253 B.n124 163.367
R418 B.n254 B.n253 163.367
R419 B.n255 B.n254 163.367
R420 B.n255 B.n120 163.367
R421 B.n260 B.n120 163.367
R422 B.n261 B.n260 163.367
R423 B.n262 B.n261 163.367
R424 B.n262 B.n118 163.367
R425 B.n266 B.n118 163.367
R426 B.n267 B.n266 163.367
R427 B.n268 B.n267 163.367
R428 B.n268 B.n116 163.367
R429 B.n275 B.n116 163.367
R430 B.n276 B.n275 163.367
R431 B.n277 B.n276 163.367
R432 B.n277 B.n114 163.367
R433 B.n281 B.n114 163.367
R434 B.n282 B.n281 163.367
R435 B.n283 B.n282 163.367
R436 B.n283 B.n112 163.367
R437 B.n287 B.n112 163.367
R438 B.n288 B.n287 163.367
R439 B.n289 B.n288 163.367
R440 B.n289 B.n110 163.367
R441 B.n293 B.n110 163.367
R442 B.n294 B.n293 163.367
R443 B.n295 B.n294 163.367
R444 B.n295 B.n108 163.367
R445 B.n299 B.n108 163.367
R446 B.n300 B.n299 163.367
R447 B.n301 B.n300 163.367
R448 B.n301 B.n106 163.367
R449 B.n305 B.n106 163.367
R450 B.n306 B.n305 163.367
R451 B.n307 B.n306 163.367
R452 B.n307 B.n104 163.367
R453 B.n311 B.n104 163.367
R454 B.n312 B.n311 163.367
R455 B.n313 B.n312 163.367
R456 B.n313 B.n102 163.367
R457 B.n317 B.n102 163.367
R458 B.n319 B.n318 163.367
R459 B.n319 B.n100 163.367
R460 B.n323 B.n100 163.367
R461 B.n324 B.n323 163.367
R462 B.n325 B.n324 163.367
R463 B.n325 B.n98 163.367
R464 B.n329 B.n98 163.367
R465 B.n330 B.n329 163.367
R466 B.n331 B.n330 163.367
R467 B.n331 B.n96 163.367
R468 B.n335 B.n96 163.367
R469 B.n336 B.n335 163.367
R470 B.n337 B.n336 163.367
R471 B.n337 B.n94 163.367
R472 B.n341 B.n94 163.367
R473 B.n342 B.n341 163.367
R474 B.n343 B.n342 163.367
R475 B.n343 B.n92 163.367
R476 B.n347 B.n92 163.367
R477 B.n348 B.n347 163.367
R478 B.n349 B.n348 163.367
R479 B.n349 B.n90 163.367
R480 B.n353 B.n90 163.367
R481 B.n354 B.n353 163.367
R482 B.n355 B.n354 163.367
R483 B.n355 B.n88 163.367
R484 B.n359 B.n88 163.367
R485 B.n360 B.n359 163.367
R486 B.n361 B.n360 163.367
R487 B.n361 B.n86 163.367
R488 B.n365 B.n86 163.367
R489 B.n366 B.n365 163.367
R490 B.n367 B.n366 163.367
R491 B.n367 B.n84 163.367
R492 B.n371 B.n84 163.367
R493 B.n372 B.n371 163.367
R494 B.n373 B.n372 163.367
R495 B.n373 B.n82 163.367
R496 B.n377 B.n82 163.367
R497 B.n378 B.n377 163.367
R498 B.n379 B.n378 163.367
R499 B.n379 B.n80 163.367
R500 B.n383 B.n80 163.367
R501 B.n384 B.n383 163.367
R502 B.n385 B.n384 163.367
R503 B.n385 B.n78 163.367
R504 B.n389 B.n78 163.367
R505 B.n390 B.n389 163.367
R506 B.n391 B.n390 163.367
R507 B.n391 B.n76 163.367
R508 B.n395 B.n76 163.367
R509 B.n396 B.n395 163.367
R510 B.n397 B.n396 163.367
R511 B.n397 B.n74 163.367
R512 B.n401 B.n74 163.367
R513 B.n402 B.n401 163.367
R514 B.n403 B.n402 163.367
R515 B.n403 B.n72 163.367
R516 B.n407 B.n72 163.367
R517 B.n408 B.n407 163.367
R518 B.n409 B.n408 163.367
R519 B.n409 B.n70 163.367
R520 B.n413 B.n70 163.367
R521 B.n414 B.n413 163.367
R522 B.n415 B.n414 163.367
R523 B.n415 B.n68 163.367
R524 B.n419 B.n68 163.367
R525 B.n420 B.n419 163.367
R526 B.n421 B.n420 163.367
R527 B.n421 B.n66 163.367
R528 B.n425 B.n66 163.367
R529 B.n426 B.n425 163.367
R530 B.n427 B.n426 163.367
R531 B.n427 B.n64 163.367
R532 B.n431 B.n64 163.367
R533 B.n432 B.n431 163.367
R534 B.n433 B.n432 163.367
R535 B.n433 B.n62 163.367
R536 B.n437 B.n62 163.367
R537 B.n438 B.n437 163.367
R538 B.n439 B.n438 163.367
R539 B.n439 B.n60 163.367
R540 B.n540 B.n23 163.367
R541 B.n536 B.n23 163.367
R542 B.n536 B.n535 163.367
R543 B.n535 B.n534 163.367
R544 B.n534 B.n25 163.367
R545 B.n530 B.n25 163.367
R546 B.n530 B.n529 163.367
R547 B.n529 B.n528 163.367
R548 B.n528 B.n27 163.367
R549 B.n524 B.n27 163.367
R550 B.n524 B.n523 163.367
R551 B.n523 B.n522 163.367
R552 B.n522 B.n29 163.367
R553 B.n518 B.n29 163.367
R554 B.n518 B.n517 163.367
R555 B.n517 B.n516 163.367
R556 B.n516 B.n31 163.367
R557 B.n512 B.n31 163.367
R558 B.n512 B.n511 163.367
R559 B.n511 B.n510 163.367
R560 B.n510 B.n33 163.367
R561 B.n506 B.n33 163.367
R562 B.n506 B.n505 163.367
R563 B.n505 B.n504 163.367
R564 B.n504 B.n35 163.367
R565 B.n500 B.n35 163.367
R566 B.n500 B.n499 163.367
R567 B.n499 B.n498 163.367
R568 B.n498 B.n37 163.367
R569 B.n494 B.n37 163.367
R570 B.n494 B.n493 163.367
R571 B.n493 B.n492 163.367
R572 B.n492 B.n42 163.367
R573 B.n488 B.n42 163.367
R574 B.n488 B.n487 163.367
R575 B.n487 B.n486 163.367
R576 B.n486 B.n44 163.367
R577 B.n481 B.n44 163.367
R578 B.n481 B.n480 163.367
R579 B.n480 B.n479 163.367
R580 B.n479 B.n48 163.367
R581 B.n475 B.n48 163.367
R582 B.n475 B.n474 163.367
R583 B.n474 B.n473 163.367
R584 B.n473 B.n50 163.367
R585 B.n469 B.n50 163.367
R586 B.n469 B.n468 163.367
R587 B.n468 B.n467 163.367
R588 B.n467 B.n52 163.367
R589 B.n463 B.n52 163.367
R590 B.n463 B.n462 163.367
R591 B.n462 B.n461 163.367
R592 B.n461 B.n54 163.367
R593 B.n457 B.n54 163.367
R594 B.n457 B.n456 163.367
R595 B.n456 B.n455 163.367
R596 B.n455 B.n56 163.367
R597 B.n451 B.n56 163.367
R598 B.n451 B.n450 163.367
R599 B.n450 B.n449 163.367
R600 B.n449 B.n58 163.367
R601 B.n445 B.n58 163.367
R602 B.n445 B.n444 163.367
R603 B.n444 B.n443 163.367
R604 B.n272 B.n271 71.952
R605 B.n122 B.n121 71.952
R606 B.n39 B.n38 71.952
R607 B.n46 B.n45 71.952
R608 B.n273 B.n272 59.5399
R609 B.n258 B.n122 59.5399
R610 B.n40 B.n39 59.5399
R611 B.n484 B.n46 59.5399
R612 B.n539 B.n22 28.8785
R613 B.n442 B.n441 28.8785
R614 B.n316 B.n101 28.8785
R615 B.n216 B.n215 28.8785
R616 B B.n603 18.0485
R617 B.n539 B.n538 10.6151
R618 B.n538 B.n537 10.6151
R619 B.n537 B.n24 10.6151
R620 B.n533 B.n24 10.6151
R621 B.n533 B.n532 10.6151
R622 B.n532 B.n531 10.6151
R623 B.n531 B.n26 10.6151
R624 B.n527 B.n26 10.6151
R625 B.n527 B.n526 10.6151
R626 B.n526 B.n525 10.6151
R627 B.n525 B.n28 10.6151
R628 B.n521 B.n28 10.6151
R629 B.n521 B.n520 10.6151
R630 B.n520 B.n519 10.6151
R631 B.n519 B.n30 10.6151
R632 B.n515 B.n30 10.6151
R633 B.n515 B.n514 10.6151
R634 B.n514 B.n513 10.6151
R635 B.n513 B.n32 10.6151
R636 B.n509 B.n32 10.6151
R637 B.n509 B.n508 10.6151
R638 B.n508 B.n507 10.6151
R639 B.n507 B.n34 10.6151
R640 B.n503 B.n34 10.6151
R641 B.n503 B.n502 10.6151
R642 B.n502 B.n501 10.6151
R643 B.n501 B.n36 10.6151
R644 B.n497 B.n496 10.6151
R645 B.n496 B.n495 10.6151
R646 B.n495 B.n41 10.6151
R647 B.n491 B.n41 10.6151
R648 B.n491 B.n490 10.6151
R649 B.n490 B.n489 10.6151
R650 B.n489 B.n43 10.6151
R651 B.n485 B.n43 10.6151
R652 B.n483 B.n482 10.6151
R653 B.n482 B.n47 10.6151
R654 B.n478 B.n47 10.6151
R655 B.n478 B.n477 10.6151
R656 B.n477 B.n476 10.6151
R657 B.n476 B.n49 10.6151
R658 B.n472 B.n49 10.6151
R659 B.n472 B.n471 10.6151
R660 B.n471 B.n470 10.6151
R661 B.n470 B.n51 10.6151
R662 B.n466 B.n51 10.6151
R663 B.n466 B.n465 10.6151
R664 B.n465 B.n464 10.6151
R665 B.n464 B.n53 10.6151
R666 B.n460 B.n53 10.6151
R667 B.n460 B.n459 10.6151
R668 B.n459 B.n458 10.6151
R669 B.n458 B.n55 10.6151
R670 B.n454 B.n55 10.6151
R671 B.n454 B.n453 10.6151
R672 B.n453 B.n452 10.6151
R673 B.n452 B.n57 10.6151
R674 B.n448 B.n57 10.6151
R675 B.n448 B.n447 10.6151
R676 B.n447 B.n446 10.6151
R677 B.n446 B.n59 10.6151
R678 B.n442 B.n59 10.6151
R679 B.n320 B.n101 10.6151
R680 B.n321 B.n320 10.6151
R681 B.n322 B.n321 10.6151
R682 B.n322 B.n99 10.6151
R683 B.n326 B.n99 10.6151
R684 B.n327 B.n326 10.6151
R685 B.n328 B.n327 10.6151
R686 B.n328 B.n97 10.6151
R687 B.n332 B.n97 10.6151
R688 B.n333 B.n332 10.6151
R689 B.n334 B.n333 10.6151
R690 B.n334 B.n95 10.6151
R691 B.n338 B.n95 10.6151
R692 B.n339 B.n338 10.6151
R693 B.n340 B.n339 10.6151
R694 B.n340 B.n93 10.6151
R695 B.n344 B.n93 10.6151
R696 B.n345 B.n344 10.6151
R697 B.n346 B.n345 10.6151
R698 B.n346 B.n91 10.6151
R699 B.n350 B.n91 10.6151
R700 B.n351 B.n350 10.6151
R701 B.n352 B.n351 10.6151
R702 B.n352 B.n89 10.6151
R703 B.n356 B.n89 10.6151
R704 B.n357 B.n356 10.6151
R705 B.n358 B.n357 10.6151
R706 B.n358 B.n87 10.6151
R707 B.n362 B.n87 10.6151
R708 B.n363 B.n362 10.6151
R709 B.n364 B.n363 10.6151
R710 B.n364 B.n85 10.6151
R711 B.n368 B.n85 10.6151
R712 B.n369 B.n368 10.6151
R713 B.n370 B.n369 10.6151
R714 B.n370 B.n83 10.6151
R715 B.n374 B.n83 10.6151
R716 B.n375 B.n374 10.6151
R717 B.n376 B.n375 10.6151
R718 B.n376 B.n81 10.6151
R719 B.n380 B.n81 10.6151
R720 B.n381 B.n380 10.6151
R721 B.n382 B.n381 10.6151
R722 B.n382 B.n79 10.6151
R723 B.n386 B.n79 10.6151
R724 B.n387 B.n386 10.6151
R725 B.n388 B.n387 10.6151
R726 B.n388 B.n77 10.6151
R727 B.n392 B.n77 10.6151
R728 B.n393 B.n392 10.6151
R729 B.n394 B.n393 10.6151
R730 B.n394 B.n75 10.6151
R731 B.n398 B.n75 10.6151
R732 B.n399 B.n398 10.6151
R733 B.n400 B.n399 10.6151
R734 B.n400 B.n73 10.6151
R735 B.n404 B.n73 10.6151
R736 B.n405 B.n404 10.6151
R737 B.n406 B.n405 10.6151
R738 B.n406 B.n71 10.6151
R739 B.n410 B.n71 10.6151
R740 B.n411 B.n410 10.6151
R741 B.n412 B.n411 10.6151
R742 B.n412 B.n69 10.6151
R743 B.n416 B.n69 10.6151
R744 B.n417 B.n416 10.6151
R745 B.n418 B.n417 10.6151
R746 B.n418 B.n67 10.6151
R747 B.n422 B.n67 10.6151
R748 B.n423 B.n422 10.6151
R749 B.n424 B.n423 10.6151
R750 B.n424 B.n65 10.6151
R751 B.n428 B.n65 10.6151
R752 B.n429 B.n428 10.6151
R753 B.n430 B.n429 10.6151
R754 B.n430 B.n63 10.6151
R755 B.n434 B.n63 10.6151
R756 B.n435 B.n434 10.6151
R757 B.n436 B.n435 10.6151
R758 B.n436 B.n61 10.6151
R759 B.n440 B.n61 10.6151
R760 B.n441 B.n440 10.6151
R761 B.n216 B.n135 10.6151
R762 B.n220 B.n135 10.6151
R763 B.n221 B.n220 10.6151
R764 B.n222 B.n221 10.6151
R765 B.n222 B.n133 10.6151
R766 B.n226 B.n133 10.6151
R767 B.n227 B.n226 10.6151
R768 B.n228 B.n227 10.6151
R769 B.n228 B.n131 10.6151
R770 B.n232 B.n131 10.6151
R771 B.n233 B.n232 10.6151
R772 B.n234 B.n233 10.6151
R773 B.n234 B.n129 10.6151
R774 B.n238 B.n129 10.6151
R775 B.n239 B.n238 10.6151
R776 B.n240 B.n239 10.6151
R777 B.n240 B.n127 10.6151
R778 B.n244 B.n127 10.6151
R779 B.n245 B.n244 10.6151
R780 B.n246 B.n245 10.6151
R781 B.n246 B.n125 10.6151
R782 B.n250 B.n125 10.6151
R783 B.n251 B.n250 10.6151
R784 B.n252 B.n251 10.6151
R785 B.n252 B.n123 10.6151
R786 B.n256 B.n123 10.6151
R787 B.n257 B.n256 10.6151
R788 B.n259 B.n119 10.6151
R789 B.n263 B.n119 10.6151
R790 B.n264 B.n263 10.6151
R791 B.n265 B.n264 10.6151
R792 B.n265 B.n117 10.6151
R793 B.n269 B.n117 10.6151
R794 B.n270 B.n269 10.6151
R795 B.n274 B.n270 10.6151
R796 B.n278 B.n115 10.6151
R797 B.n279 B.n278 10.6151
R798 B.n280 B.n279 10.6151
R799 B.n280 B.n113 10.6151
R800 B.n284 B.n113 10.6151
R801 B.n285 B.n284 10.6151
R802 B.n286 B.n285 10.6151
R803 B.n286 B.n111 10.6151
R804 B.n290 B.n111 10.6151
R805 B.n291 B.n290 10.6151
R806 B.n292 B.n291 10.6151
R807 B.n292 B.n109 10.6151
R808 B.n296 B.n109 10.6151
R809 B.n297 B.n296 10.6151
R810 B.n298 B.n297 10.6151
R811 B.n298 B.n107 10.6151
R812 B.n302 B.n107 10.6151
R813 B.n303 B.n302 10.6151
R814 B.n304 B.n303 10.6151
R815 B.n304 B.n105 10.6151
R816 B.n308 B.n105 10.6151
R817 B.n309 B.n308 10.6151
R818 B.n310 B.n309 10.6151
R819 B.n310 B.n103 10.6151
R820 B.n314 B.n103 10.6151
R821 B.n315 B.n314 10.6151
R822 B.n316 B.n315 10.6151
R823 B.n215 B.n214 10.6151
R824 B.n214 B.n137 10.6151
R825 B.n210 B.n137 10.6151
R826 B.n210 B.n209 10.6151
R827 B.n209 B.n208 10.6151
R828 B.n208 B.n139 10.6151
R829 B.n204 B.n139 10.6151
R830 B.n204 B.n203 10.6151
R831 B.n203 B.n202 10.6151
R832 B.n202 B.n141 10.6151
R833 B.n198 B.n141 10.6151
R834 B.n198 B.n197 10.6151
R835 B.n197 B.n196 10.6151
R836 B.n196 B.n143 10.6151
R837 B.n192 B.n143 10.6151
R838 B.n192 B.n191 10.6151
R839 B.n191 B.n190 10.6151
R840 B.n190 B.n145 10.6151
R841 B.n186 B.n145 10.6151
R842 B.n186 B.n185 10.6151
R843 B.n185 B.n184 10.6151
R844 B.n184 B.n147 10.6151
R845 B.n180 B.n147 10.6151
R846 B.n180 B.n179 10.6151
R847 B.n179 B.n178 10.6151
R848 B.n178 B.n149 10.6151
R849 B.n174 B.n149 10.6151
R850 B.n174 B.n173 10.6151
R851 B.n173 B.n172 10.6151
R852 B.n172 B.n151 10.6151
R853 B.n168 B.n151 10.6151
R854 B.n168 B.n167 10.6151
R855 B.n167 B.n166 10.6151
R856 B.n166 B.n153 10.6151
R857 B.n162 B.n153 10.6151
R858 B.n162 B.n161 10.6151
R859 B.n161 B.n160 10.6151
R860 B.n160 B.n155 10.6151
R861 B.n156 B.n155 10.6151
R862 B.n156 B.n0 10.6151
R863 B.n599 B.n1 10.6151
R864 B.n599 B.n598 10.6151
R865 B.n598 B.n597 10.6151
R866 B.n597 B.n4 10.6151
R867 B.n593 B.n4 10.6151
R868 B.n593 B.n592 10.6151
R869 B.n592 B.n591 10.6151
R870 B.n591 B.n6 10.6151
R871 B.n587 B.n6 10.6151
R872 B.n587 B.n586 10.6151
R873 B.n586 B.n585 10.6151
R874 B.n585 B.n8 10.6151
R875 B.n581 B.n8 10.6151
R876 B.n581 B.n580 10.6151
R877 B.n580 B.n579 10.6151
R878 B.n579 B.n10 10.6151
R879 B.n575 B.n10 10.6151
R880 B.n575 B.n574 10.6151
R881 B.n574 B.n573 10.6151
R882 B.n573 B.n12 10.6151
R883 B.n569 B.n12 10.6151
R884 B.n569 B.n568 10.6151
R885 B.n568 B.n567 10.6151
R886 B.n567 B.n14 10.6151
R887 B.n563 B.n14 10.6151
R888 B.n563 B.n562 10.6151
R889 B.n562 B.n561 10.6151
R890 B.n561 B.n16 10.6151
R891 B.n557 B.n16 10.6151
R892 B.n557 B.n556 10.6151
R893 B.n556 B.n555 10.6151
R894 B.n555 B.n18 10.6151
R895 B.n551 B.n18 10.6151
R896 B.n551 B.n550 10.6151
R897 B.n550 B.n549 10.6151
R898 B.n549 B.n20 10.6151
R899 B.n545 B.n20 10.6151
R900 B.n545 B.n544 10.6151
R901 B.n544 B.n543 10.6151
R902 B.n543 B.n22 10.6151
R903 B.n497 B.n40 6.5566
R904 B.n485 B.n484 6.5566
R905 B.n259 B.n258 6.5566
R906 B.n274 B.n273 6.5566
R907 B.n40 B.n36 4.05904
R908 B.n484 B.n483 4.05904
R909 B.n258 B.n257 4.05904
R910 B.n273 B.n115 4.05904
R911 B.n603 B.n0 2.81026
R912 B.n603 B.n1 2.81026
R913 VP.n17 VP.n16 161.3
R914 VP.n15 VP.n1 161.3
R915 VP.n14 VP.n13 161.3
R916 VP.n12 VP.n2 161.3
R917 VP.n11 VP.n10 161.3
R918 VP.n9 VP.n3 161.3
R919 VP.n8 VP.n7 161.3
R920 VP.n5 VP.t0 86.5089
R921 VP.n5 VP.t1 85.3711
R922 VP.n6 VP.n4 72.6958
R923 VP.n18 VP.n0 72.6958
R924 VP.n4 VP.t2 51.4091
R925 VP.n0 VP.t3 51.4091
R926 VP.n6 VP.n5 47.5828
R927 VP.n10 VP.n2 40.4934
R928 VP.n14 VP.n2 40.4934
R929 VP.n9 VP.n8 24.4675
R930 VP.n10 VP.n9 24.4675
R931 VP.n15 VP.n14 24.4675
R932 VP.n16 VP.n15 24.4675
R933 VP.n8 VP.n4 17.3721
R934 VP.n16 VP.n0 17.3721
R935 VP.n7 VP.n6 0.354971
R936 VP.n18 VP.n17 0.354971
R937 VP VP.n18 0.26696
R938 VP.n7 VP.n3 0.189894
R939 VP.n11 VP.n3 0.189894
R940 VP.n12 VP.n11 0.189894
R941 VP.n13 VP.n12 0.189894
R942 VP.n13 VP.n1 0.189894
R943 VP.n17 VP.n1 0.189894
R944 VDD1 VDD1.n1 127.409
R945 VDD1 VDD1.n0 87.4181
R946 VDD1.n0 VDD1.t0 4.50882
R947 VDD1.n0 VDD1.t3 4.50882
R948 VDD1.n1 VDD1.t1 4.50882
R949 VDD1.n1 VDD1.t2 4.50882
R950 VTAIL.n265 VTAIL.n264 585
R951 VTAIL.n267 VTAIL.n266 585
R952 VTAIL.n260 VTAIL.n259 585
R953 VTAIL.n273 VTAIL.n272 585
R954 VTAIL.n275 VTAIL.n274 585
R955 VTAIL.n256 VTAIL.n255 585
R956 VTAIL.n281 VTAIL.n280 585
R957 VTAIL.n283 VTAIL.n282 585
R958 VTAIL.n13 VTAIL.n12 585
R959 VTAIL.n15 VTAIL.n14 585
R960 VTAIL.n8 VTAIL.n7 585
R961 VTAIL.n21 VTAIL.n20 585
R962 VTAIL.n23 VTAIL.n22 585
R963 VTAIL.n4 VTAIL.n3 585
R964 VTAIL.n29 VTAIL.n28 585
R965 VTAIL.n31 VTAIL.n30 585
R966 VTAIL.n49 VTAIL.n48 585
R967 VTAIL.n51 VTAIL.n50 585
R968 VTAIL.n44 VTAIL.n43 585
R969 VTAIL.n57 VTAIL.n56 585
R970 VTAIL.n59 VTAIL.n58 585
R971 VTAIL.n40 VTAIL.n39 585
R972 VTAIL.n65 VTAIL.n64 585
R973 VTAIL.n67 VTAIL.n66 585
R974 VTAIL.n85 VTAIL.n84 585
R975 VTAIL.n87 VTAIL.n86 585
R976 VTAIL.n80 VTAIL.n79 585
R977 VTAIL.n93 VTAIL.n92 585
R978 VTAIL.n95 VTAIL.n94 585
R979 VTAIL.n76 VTAIL.n75 585
R980 VTAIL.n101 VTAIL.n100 585
R981 VTAIL.n103 VTAIL.n102 585
R982 VTAIL.n247 VTAIL.n246 585
R983 VTAIL.n245 VTAIL.n244 585
R984 VTAIL.n220 VTAIL.n219 585
R985 VTAIL.n239 VTAIL.n238 585
R986 VTAIL.n237 VTAIL.n236 585
R987 VTAIL.n224 VTAIL.n223 585
R988 VTAIL.n231 VTAIL.n230 585
R989 VTAIL.n229 VTAIL.n228 585
R990 VTAIL.n211 VTAIL.n210 585
R991 VTAIL.n209 VTAIL.n208 585
R992 VTAIL.n184 VTAIL.n183 585
R993 VTAIL.n203 VTAIL.n202 585
R994 VTAIL.n201 VTAIL.n200 585
R995 VTAIL.n188 VTAIL.n187 585
R996 VTAIL.n195 VTAIL.n194 585
R997 VTAIL.n193 VTAIL.n192 585
R998 VTAIL.n175 VTAIL.n174 585
R999 VTAIL.n173 VTAIL.n172 585
R1000 VTAIL.n148 VTAIL.n147 585
R1001 VTAIL.n167 VTAIL.n166 585
R1002 VTAIL.n165 VTAIL.n164 585
R1003 VTAIL.n152 VTAIL.n151 585
R1004 VTAIL.n159 VTAIL.n158 585
R1005 VTAIL.n157 VTAIL.n156 585
R1006 VTAIL.n139 VTAIL.n138 585
R1007 VTAIL.n137 VTAIL.n136 585
R1008 VTAIL.n112 VTAIL.n111 585
R1009 VTAIL.n131 VTAIL.n130 585
R1010 VTAIL.n129 VTAIL.n128 585
R1011 VTAIL.n116 VTAIL.n115 585
R1012 VTAIL.n123 VTAIL.n122 585
R1013 VTAIL.n121 VTAIL.n120 585
R1014 VTAIL.n282 VTAIL.n252 498.474
R1015 VTAIL.n30 VTAIL.n0 498.474
R1016 VTAIL.n66 VTAIL.n36 498.474
R1017 VTAIL.n102 VTAIL.n72 498.474
R1018 VTAIL.n246 VTAIL.n216 498.474
R1019 VTAIL.n210 VTAIL.n180 498.474
R1020 VTAIL.n174 VTAIL.n144 498.474
R1021 VTAIL.n138 VTAIL.n108 498.474
R1022 VTAIL.n263 VTAIL.t3 329.053
R1023 VTAIL.n11 VTAIL.t1 329.053
R1024 VTAIL.n47 VTAIL.t4 329.053
R1025 VTAIL.n83 VTAIL.t5 329.053
R1026 VTAIL.n227 VTAIL.t6 329.053
R1027 VTAIL.n191 VTAIL.t7 329.053
R1028 VTAIL.n155 VTAIL.t0 329.053
R1029 VTAIL.n119 VTAIL.t2 329.053
R1030 VTAIL.n266 VTAIL.n265 171.744
R1031 VTAIL.n266 VTAIL.n259 171.744
R1032 VTAIL.n273 VTAIL.n259 171.744
R1033 VTAIL.n274 VTAIL.n273 171.744
R1034 VTAIL.n274 VTAIL.n255 171.744
R1035 VTAIL.n281 VTAIL.n255 171.744
R1036 VTAIL.n282 VTAIL.n281 171.744
R1037 VTAIL.n14 VTAIL.n13 171.744
R1038 VTAIL.n14 VTAIL.n7 171.744
R1039 VTAIL.n21 VTAIL.n7 171.744
R1040 VTAIL.n22 VTAIL.n21 171.744
R1041 VTAIL.n22 VTAIL.n3 171.744
R1042 VTAIL.n29 VTAIL.n3 171.744
R1043 VTAIL.n30 VTAIL.n29 171.744
R1044 VTAIL.n50 VTAIL.n49 171.744
R1045 VTAIL.n50 VTAIL.n43 171.744
R1046 VTAIL.n57 VTAIL.n43 171.744
R1047 VTAIL.n58 VTAIL.n57 171.744
R1048 VTAIL.n58 VTAIL.n39 171.744
R1049 VTAIL.n65 VTAIL.n39 171.744
R1050 VTAIL.n66 VTAIL.n65 171.744
R1051 VTAIL.n86 VTAIL.n85 171.744
R1052 VTAIL.n86 VTAIL.n79 171.744
R1053 VTAIL.n93 VTAIL.n79 171.744
R1054 VTAIL.n94 VTAIL.n93 171.744
R1055 VTAIL.n94 VTAIL.n75 171.744
R1056 VTAIL.n101 VTAIL.n75 171.744
R1057 VTAIL.n102 VTAIL.n101 171.744
R1058 VTAIL.n246 VTAIL.n245 171.744
R1059 VTAIL.n245 VTAIL.n219 171.744
R1060 VTAIL.n238 VTAIL.n219 171.744
R1061 VTAIL.n238 VTAIL.n237 171.744
R1062 VTAIL.n237 VTAIL.n223 171.744
R1063 VTAIL.n230 VTAIL.n223 171.744
R1064 VTAIL.n230 VTAIL.n229 171.744
R1065 VTAIL.n210 VTAIL.n209 171.744
R1066 VTAIL.n209 VTAIL.n183 171.744
R1067 VTAIL.n202 VTAIL.n183 171.744
R1068 VTAIL.n202 VTAIL.n201 171.744
R1069 VTAIL.n201 VTAIL.n187 171.744
R1070 VTAIL.n194 VTAIL.n187 171.744
R1071 VTAIL.n194 VTAIL.n193 171.744
R1072 VTAIL.n174 VTAIL.n173 171.744
R1073 VTAIL.n173 VTAIL.n147 171.744
R1074 VTAIL.n166 VTAIL.n147 171.744
R1075 VTAIL.n166 VTAIL.n165 171.744
R1076 VTAIL.n165 VTAIL.n151 171.744
R1077 VTAIL.n158 VTAIL.n151 171.744
R1078 VTAIL.n158 VTAIL.n157 171.744
R1079 VTAIL.n138 VTAIL.n137 171.744
R1080 VTAIL.n137 VTAIL.n111 171.744
R1081 VTAIL.n130 VTAIL.n111 171.744
R1082 VTAIL.n130 VTAIL.n129 171.744
R1083 VTAIL.n129 VTAIL.n115 171.744
R1084 VTAIL.n122 VTAIL.n115 171.744
R1085 VTAIL.n122 VTAIL.n121 171.744
R1086 VTAIL.n265 VTAIL.t3 85.8723
R1087 VTAIL.n13 VTAIL.t1 85.8723
R1088 VTAIL.n49 VTAIL.t4 85.8723
R1089 VTAIL.n85 VTAIL.t5 85.8723
R1090 VTAIL.n229 VTAIL.t6 85.8723
R1091 VTAIL.n193 VTAIL.t7 85.8723
R1092 VTAIL.n157 VTAIL.t0 85.8723
R1093 VTAIL.n121 VTAIL.t2 85.8723
R1094 VTAIL.n287 VTAIL.n286 34.7066
R1095 VTAIL.n35 VTAIL.n34 34.7066
R1096 VTAIL.n71 VTAIL.n70 34.7066
R1097 VTAIL.n107 VTAIL.n106 34.7066
R1098 VTAIL.n251 VTAIL.n250 34.7066
R1099 VTAIL.n215 VTAIL.n214 34.7066
R1100 VTAIL.n179 VTAIL.n178 34.7066
R1101 VTAIL.n143 VTAIL.n142 34.7066
R1102 VTAIL.n287 VTAIL.n251 21.7807
R1103 VTAIL.n143 VTAIL.n107 21.7807
R1104 VTAIL.n284 VTAIL.n283 12.8005
R1105 VTAIL.n32 VTAIL.n31 12.8005
R1106 VTAIL.n68 VTAIL.n67 12.8005
R1107 VTAIL.n104 VTAIL.n103 12.8005
R1108 VTAIL.n248 VTAIL.n247 12.8005
R1109 VTAIL.n212 VTAIL.n211 12.8005
R1110 VTAIL.n176 VTAIL.n175 12.8005
R1111 VTAIL.n140 VTAIL.n139 12.8005
R1112 VTAIL.n280 VTAIL.n254 12.0247
R1113 VTAIL.n28 VTAIL.n2 12.0247
R1114 VTAIL.n64 VTAIL.n38 12.0247
R1115 VTAIL.n100 VTAIL.n74 12.0247
R1116 VTAIL.n244 VTAIL.n218 12.0247
R1117 VTAIL.n208 VTAIL.n182 12.0247
R1118 VTAIL.n172 VTAIL.n146 12.0247
R1119 VTAIL.n136 VTAIL.n110 12.0247
R1120 VTAIL.n279 VTAIL.n256 11.249
R1121 VTAIL.n27 VTAIL.n4 11.249
R1122 VTAIL.n63 VTAIL.n40 11.249
R1123 VTAIL.n99 VTAIL.n76 11.249
R1124 VTAIL.n243 VTAIL.n220 11.249
R1125 VTAIL.n207 VTAIL.n184 11.249
R1126 VTAIL.n171 VTAIL.n148 11.249
R1127 VTAIL.n135 VTAIL.n112 11.249
R1128 VTAIL.n264 VTAIL.n263 10.7237
R1129 VTAIL.n12 VTAIL.n11 10.7237
R1130 VTAIL.n48 VTAIL.n47 10.7237
R1131 VTAIL.n84 VTAIL.n83 10.7237
R1132 VTAIL.n228 VTAIL.n227 10.7237
R1133 VTAIL.n192 VTAIL.n191 10.7237
R1134 VTAIL.n156 VTAIL.n155 10.7237
R1135 VTAIL.n120 VTAIL.n119 10.7237
R1136 VTAIL.n276 VTAIL.n275 10.4732
R1137 VTAIL.n24 VTAIL.n23 10.4732
R1138 VTAIL.n60 VTAIL.n59 10.4732
R1139 VTAIL.n96 VTAIL.n95 10.4732
R1140 VTAIL.n240 VTAIL.n239 10.4732
R1141 VTAIL.n204 VTAIL.n203 10.4732
R1142 VTAIL.n168 VTAIL.n167 10.4732
R1143 VTAIL.n132 VTAIL.n131 10.4732
R1144 VTAIL.n272 VTAIL.n258 9.69747
R1145 VTAIL.n20 VTAIL.n6 9.69747
R1146 VTAIL.n56 VTAIL.n42 9.69747
R1147 VTAIL.n92 VTAIL.n78 9.69747
R1148 VTAIL.n236 VTAIL.n222 9.69747
R1149 VTAIL.n200 VTAIL.n186 9.69747
R1150 VTAIL.n164 VTAIL.n150 9.69747
R1151 VTAIL.n128 VTAIL.n114 9.69747
R1152 VTAIL.n286 VTAIL.n285 9.45567
R1153 VTAIL.n34 VTAIL.n33 9.45567
R1154 VTAIL.n70 VTAIL.n69 9.45567
R1155 VTAIL.n106 VTAIL.n105 9.45567
R1156 VTAIL.n250 VTAIL.n249 9.45567
R1157 VTAIL.n214 VTAIL.n213 9.45567
R1158 VTAIL.n178 VTAIL.n177 9.45567
R1159 VTAIL.n142 VTAIL.n141 9.45567
R1160 VTAIL.n262 VTAIL.n261 9.3005
R1161 VTAIL.n269 VTAIL.n268 9.3005
R1162 VTAIL.n271 VTAIL.n270 9.3005
R1163 VTAIL.n258 VTAIL.n257 9.3005
R1164 VTAIL.n277 VTAIL.n276 9.3005
R1165 VTAIL.n279 VTAIL.n278 9.3005
R1166 VTAIL.n254 VTAIL.n253 9.3005
R1167 VTAIL.n285 VTAIL.n284 9.3005
R1168 VTAIL.n10 VTAIL.n9 9.3005
R1169 VTAIL.n17 VTAIL.n16 9.3005
R1170 VTAIL.n19 VTAIL.n18 9.3005
R1171 VTAIL.n6 VTAIL.n5 9.3005
R1172 VTAIL.n25 VTAIL.n24 9.3005
R1173 VTAIL.n27 VTAIL.n26 9.3005
R1174 VTAIL.n2 VTAIL.n1 9.3005
R1175 VTAIL.n33 VTAIL.n32 9.3005
R1176 VTAIL.n46 VTAIL.n45 9.3005
R1177 VTAIL.n53 VTAIL.n52 9.3005
R1178 VTAIL.n55 VTAIL.n54 9.3005
R1179 VTAIL.n42 VTAIL.n41 9.3005
R1180 VTAIL.n61 VTAIL.n60 9.3005
R1181 VTAIL.n63 VTAIL.n62 9.3005
R1182 VTAIL.n38 VTAIL.n37 9.3005
R1183 VTAIL.n69 VTAIL.n68 9.3005
R1184 VTAIL.n82 VTAIL.n81 9.3005
R1185 VTAIL.n89 VTAIL.n88 9.3005
R1186 VTAIL.n91 VTAIL.n90 9.3005
R1187 VTAIL.n78 VTAIL.n77 9.3005
R1188 VTAIL.n97 VTAIL.n96 9.3005
R1189 VTAIL.n99 VTAIL.n98 9.3005
R1190 VTAIL.n74 VTAIL.n73 9.3005
R1191 VTAIL.n105 VTAIL.n104 9.3005
R1192 VTAIL.n226 VTAIL.n225 9.3005
R1193 VTAIL.n233 VTAIL.n232 9.3005
R1194 VTAIL.n235 VTAIL.n234 9.3005
R1195 VTAIL.n222 VTAIL.n221 9.3005
R1196 VTAIL.n241 VTAIL.n240 9.3005
R1197 VTAIL.n243 VTAIL.n242 9.3005
R1198 VTAIL.n218 VTAIL.n217 9.3005
R1199 VTAIL.n249 VTAIL.n248 9.3005
R1200 VTAIL.n190 VTAIL.n189 9.3005
R1201 VTAIL.n197 VTAIL.n196 9.3005
R1202 VTAIL.n199 VTAIL.n198 9.3005
R1203 VTAIL.n186 VTAIL.n185 9.3005
R1204 VTAIL.n205 VTAIL.n204 9.3005
R1205 VTAIL.n207 VTAIL.n206 9.3005
R1206 VTAIL.n182 VTAIL.n181 9.3005
R1207 VTAIL.n213 VTAIL.n212 9.3005
R1208 VTAIL.n154 VTAIL.n153 9.3005
R1209 VTAIL.n161 VTAIL.n160 9.3005
R1210 VTAIL.n163 VTAIL.n162 9.3005
R1211 VTAIL.n150 VTAIL.n149 9.3005
R1212 VTAIL.n169 VTAIL.n168 9.3005
R1213 VTAIL.n171 VTAIL.n170 9.3005
R1214 VTAIL.n146 VTAIL.n145 9.3005
R1215 VTAIL.n177 VTAIL.n176 9.3005
R1216 VTAIL.n118 VTAIL.n117 9.3005
R1217 VTAIL.n125 VTAIL.n124 9.3005
R1218 VTAIL.n127 VTAIL.n126 9.3005
R1219 VTAIL.n114 VTAIL.n113 9.3005
R1220 VTAIL.n133 VTAIL.n132 9.3005
R1221 VTAIL.n135 VTAIL.n134 9.3005
R1222 VTAIL.n110 VTAIL.n109 9.3005
R1223 VTAIL.n141 VTAIL.n140 9.3005
R1224 VTAIL.n271 VTAIL.n260 8.92171
R1225 VTAIL.n19 VTAIL.n8 8.92171
R1226 VTAIL.n55 VTAIL.n44 8.92171
R1227 VTAIL.n91 VTAIL.n80 8.92171
R1228 VTAIL.n235 VTAIL.n224 8.92171
R1229 VTAIL.n199 VTAIL.n188 8.92171
R1230 VTAIL.n163 VTAIL.n152 8.92171
R1231 VTAIL.n127 VTAIL.n116 8.92171
R1232 VTAIL.n268 VTAIL.n267 8.14595
R1233 VTAIL.n16 VTAIL.n15 8.14595
R1234 VTAIL.n52 VTAIL.n51 8.14595
R1235 VTAIL.n88 VTAIL.n87 8.14595
R1236 VTAIL.n232 VTAIL.n231 8.14595
R1237 VTAIL.n196 VTAIL.n195 8.14595
R1238 VTAIL.n160 VTAIL.n159 8.14595
R1239 VTAIL.n124 VTAIL.n123 8.14595
R1240 VTAIL.n286 VTAIL.n252 7.75445
R1241 VTAIL.n34 VTAIL.n0 7.75445
R1242 VTAIL.n70 VTAIL.n36 7.75445
R1243 VTAIL.n106 VTAIL.n72 7.75445
R1244 VTAIL.n250 VTAIL.n216 7.75445
R1245 VTAIL.n214 VTAIL.n180 7.75445
R1246 VTAIL.n178 VTAIL.n144 7.75445
R1247 VTAIL.n142 VTAIL.n108 7.75445
R1248 VTAIL.n264 VTAIL.n262 7.3702
R1249 VTAIL.n12 VTAIL.n10 7.3702
R1250 VTAIL.n48 VTAIL.n46 7.3702
R1251 VTAIL.n84 VTAIL.n82 7.3702
R1252 VTAIL.n228 VTAIL.n226 7.3702
R1253 VTAIL.n192 VTAIL.n190 7.3702
R1254 VTAIL.n156 VTAIL.n154 7.3702
R1255 VTAIL.n120 VTAIL.n118 7.3702
R1256 VTAIL.n284 VTAIL.n252 6.08283
R1257 VTAIL.n32 VTAIL.n0 6.08283
R1258 VTAIL.n68 VTAIL.n36 6.08283
R1259 VTAIL.n104 VTAIL.n72 6.08283
R1260 VTAIL.n248 VTAIL.n216 6.08283
R1261 VTAIL.n212 VTAIL.n180 6.08283
R1262 VTAIL.n176 VTAIL.n144 6.08283
R1263 VTAIL.n140 VTAIL.n108 6.08283
R1264 VTAIL.n267 VTAIL.n262 5.81868
R1265 VTAIL.n15 VTAIL.n10 5.81868
R1266 VTAIL.n51 VTAIL.n46 5.81868
R1267 VTAIL.n87 VTAIL.n82 5.81868
R1268 VTAIL.n231 VTAIL.n226 5.81868
R1269 VTAIL.n195 VTAIL.n190 5.81868
R1270 VTAIL.n159 VTAIL.n154 5.81868
R1271 VTAIL.n123 VTAIL.n118 5.81868
R1272 VTAIL.n268 VTAIL.n260 5.04292
R1273 VTAIL.n16 VTAIL.n8 5.04292
R1274 VTAIL.n52 VTAIL.n44 5.04292
R1275 VTAIL.n88 VTAIL.n80 5.04292
R1276 VTAIL.n232 VTAIL.n224 5.04292
R1277 VTAIL.n196 VTAIL.n188 5.04292
R1278 VTAIL.n160 VTAIL.n152 5.04292
R1279 VTAIL.n124 VTAIL.n116 5.04292
R1280 VTAIL.n272 VTAIL.n271 4.26717
R1281 VTAIL.n20 VTAIL.n19 4.26717
R1282 VTAIL.n56 VTAIL.n55 4.26717
R1283 VTAIL.n92 VTAIL.n91 4.26717
R1284 VTAIL.n236 VTAIL.n235 4.26717
R1285 VTAIL.n200 VTAIL.n199 4.26717
R1286 VTAIL.n164 VTAIL.n163 4.26717
R1287 VTAIL.n128 VTAIL.n127 4.26717
R1288 VTAIL.n275 VTAIL.n258 3.49141
R1289 VTAIL.n23 VTAIL.n6 3.49141
R1290 VTAIL.n59 VTAIL.n42 3.49141
R1291 VTAIL.n95 VTAIL.n78 3.49141
R1292 VTAIL.n239 VTAIL.n222 3.49141
R1293 VTAIL.n203 VTAIL.n186 3.49141
R1294 VTAIL.n167 VTAIL.n150 3.49141
R1295 VTAIL.n131 VTAIL.n114 3.49141
R1296 VTAIL.n179 VTAIL.n143 3.19878
R1297 VTAIL.n251 VTAIL.n215 3.19878
R1298 VTAIL.n107 VTAIL.n71 3.19878
R1299 VTAIL.n276 VTAIL.n256 2.71565
R1300 VTAIL.n24 VTAIL.n4 2.71565
R1301 VTAIL.n60 VTAIL.n40 2.71565
R1302 VTAIL.n96 VTAIL.n76 2.71565
R1303 VTAIL.n240 VTAIL.n220 2.71565
R1304 VTAIL.n204 VTAIL.n184 2.71565
R1305 VTAIL.n168 VTAIL.n148 2.71565
R1306 VTAIL.n132 VTAIL.n112 2.71565
R1307 VTAIL.n263 VTAIL.n261 2.41305
R1308 VTAIL.n11 VTAIL.n9 2.41305
R1309 VTAIL.n47 VTAIL.n45 2.41305
R1310 VTAIL.n83 VTAIL.n81 2.41305
R1311 VTAIL.n227 VTAIL.n225 2.41305
R1312 VTAIL.n191 VTAIL.n189 2.41305
R1313 VTAIL.n155 VTAIL.n153 2.41305
R1314 VTAIL.n119 VTAIL.n117 2.41305
R1315 VTAIL.n280 VTAIL.n279 1.93989
R1316 VTAIL.n28 VTAIL.n27 1.93989
R1317 VTAIL.n64 VTAIL.n63 1.93989
R1318 VTAIL.n100 VTAIL.n99 1.93989
R1319 VTAIL.n244 VTAIL.n243 1.93989
R1320 VTAIL.n208 VTAIL.n207 1.93989
R1321 VTAIL.n172 VTAIL.n171 1.93989
R1322 VTAIL.n136 VTAIL.n135 1.93989
R1323 VTAIL VTAIL.n35 1.65783
R1324 VTAIL VTAIL.n287 1.54145
R1325 VTAIL.n283 VTAIL.n254 1.16414
R1326 VTAIL.n31 VTAIL.n2 1.16414
R1327 VTAIL.n67 VTAIL.n38 1.16414
R1328 VTAIL.n103 VTAIL.n74 1.16414
R1329 VTAIL.n247 VTAIL.n218 1.16414
R1330 VTAIL.n211 VTAIL.n182 1.16414
R1331 VTAIL.n175 VTAIL.n146 1.16414
R1332 VTAIL.n139 VTAIL.n110 1.16414
R1333 VTAIL.n215 VTAIL.n179 0.470328
R1334 VTAIL.n71 VTAIL.n35 0.470328
R1335 VTAIL.n269 VTAIL.n261 0.155672
R1336 VTAIL.n270 VTAIL.n269 0.155672
R1337 VTAIL.n270 VTAIL.n257 0.155672
R1338 VTAIL.n277 VTAIL.n257 0.155672
R1339 VTAIL.n278 VTAIL.n277 0.155672
R1340 VTAIL.n278 VTAIL.n253 0.155672
R1341 VTAIL.n285 VTAIL.n253 0.155672
R1342 VTAIL.n17 VTAIL.n9 0.155672
R1343 VTAIL.n18 VTAIL.n17 0.155672
R1344 VTAIL.n18 VTAIL.n5 0.155672
R1345 VTAIL.n25 VTAIL.n5 0.155672
R1346 VTAIL.n26 VTAIL.n25 0.155672
R1347 VTAIL.n26 VTAIL.n1 0.155672
R1348 VTAIL.n33 VTAIL.n1 0.155672
R1349 VTAIL.n53 VTAIL.n45 0.155672
R1350 VTAIL.n54 VTAIL.n53 0.155672
R1351 VTAIL.n54 VTAIL.n41 0.155672
R1352 VTAIL.n61 VTAIL.n41 0.155672
R1353 VTAIL.n62 VTAIL.n61 0.155672
R1354 VTAIL.n62 VTAIL.n37 0.155672
R1355 VTAIL.n69 VTAIL.n37 0.155672
R1356 VTAIL.n89 VTAIL.n81 0.155672
R1357 VTAIL.n90 VTAIL.n89 0.155672
R1358 VTAIL.n90 VTAIL.n77 0.155672
R1359 VTAIL.n97 VTAIL.n77 0.155672
R1360 VTAIL.n98 VTAIL.n97 0.155672
R1361 VTAIL.n98 VTAIL.n73 0.155672
R1362 VTAIL.n105 VTAIL.n73 0.155672
R1363 VTAIL.n249 VTAIL.n217 0.155672
R1364 VTAIL.n242 VTAIL.n217 0.155672
R1365 VTAIL.n242 VTAIL.n241 0.155672
R1366 VTAIL.n241 VTAIL.n221 0.155672
R1367 VTAIL.n234 VTAIL.n221 0.155672
R1368 VTAIL.n234 VTAIL.n233 0.155672
R1369 VTAIL.n233 VTAIL.n225 0.155672
R1370 VTAIL.n213 VTAIL.n181 0.155672
R1371 VTAIL.n206 VTAIL.n181 0.155672
R1372 VTAIL.n206 VTAIL.n205 0.155672
R1373 VTAIL.n205 VTAIL.n185 0.155672
R1374 VTAIL.n198 VTAIL.n185 0.155672
R1375 VTAIL.n198 VTAIL.n197 0.155672
R1376 VTAIL.n197 VTAIL.n189 0.155672
R1377 VTAIL.n177 VTAIL.n145 0.155672
R1378 VTAIL.n170 VTAIL.n145 0.155672
R1379 VTAIL.n170 VTAIL.n169 0.155672
R1380 VTAIL.n169 VTAIL.n149 0.155672
R1381 VTAIL.n162 VTAIL.n149 0.155672
R1382 VTAIL.n162 VTAIL.n161 0.155672
R1383 VTAIL.n161 VTAIL.n153 0.155672
R1384 VTAIL.n141 VTAIL.n109 0.155672
R1385 VTAIL.n134 VTAIL.n109 0.155672
R1386 VTAIL.n134 VTAIL.n133 0.155672
R1387 VTAIL.n133 VTAIL.n113 0.155672
R1388 VTAIL.n126 VTAIL.n113 0.155672
R1389 VTAIL.n126 VTAIL.n125 0.155672
R1390 VTAIL.n125 VTAIL.n117 0.155672
R1391 VN.n1 VN.t1 86.5092
R1392 VN.n0 VN.t2 86.5092
R1393 VN.n0 VN.t0 85.3711
R1394 VN.n1 VN.t3 85.3711
R1395 VN VN.n1 47.7482
R1396 VN VN.n0 2.38075
R1397 VDD2.n2 VDD2.n0 126.885
R1398 VDD2.n2 VDD2.n1 87.3599
R1399 VDD2.n1 VDD2.t0 4.50882
R1400 VDD2.n1 VDD2.t2 4.50882
R1401 VDD2.n0 VDD2.t1 4.50882
R1402 VDD2.n0 VDD2.t3 4.50882
R1403 VDD2 VDD2.n2 0.0586897
C0 VN VTAIL 3.35941f
C1 VTAIL VDD1 4.56518f
C2 VN w_n3196_n2410# 5.46282f
C3 w_n3196_n2410# VDD1 1.46898f
C4 VN VDD1 0.149552f
C5 VDD2 B 1.33568f
C6 B VP 1.88919f
C7 B VTAIL 3.63613f
C8 VDD2 VP 0.443785f
C9 VDD2 VTAIL 4.62462f
C10 VTAIL VP 3.37351f
C11 B w_n3196_n2410# 8.86386f
C12 VDD2 w_n3196_n2410# 1.54232f
C13 w_n3196_n2410# VP 5.87565f
C14 B VN 1.20048f
C15 VTAIL w_n3196_n2410# 2.94878f
C16 B VDD1 1.2706f
C17 VDD2 VN 3.10948f
C18 VN VP 5.86371f
C19 VDD2 VDD1 1.20819f
C20 VDD1 VP 3.40277f
C21 VDD2 VSUBS 0.969681f
C22 VDD1 VSUBS 5.62981f
C23 VTAIL VSUBS 1.098524f
C24 VN VSUBS 5.88117f
C25 VP VSUBS 2.533082f
C26 B VSUBS 4.543282f
C27 w_n3196_n2410# VSUBS 95.7649f
C28 VDD2.t1 VSUBS 0.158068f
C29 VDD2.t3 VSUBS 0.158068f
C30 VDD2.n0 VSUBS 1.64229f
C31 VDD2.t0 VSUBS 0.158068f
C32 VDD2.t2 VSUBS 0.158068f
C33 VDD2.n1 VSUBS 1.11883f
C34 VDD2.n2 VSUBS 4.01472f
C35 VN.t0 VSUBS 2.65662f
C36 VN.t2 VSUBS 2.67015f
C37 VN.n0 VSUBS 1.56647f
C38 VN.t3 VSUBS 2.65662f
C39 VN.t1 VSUBS 2.67015f
C40 VN.n1 VSUBS 3.5078f
C41 VTAIL.n0 VSUBS 0.028838f
C42 VTAIL.n1 VSUBS 0.027054f
C43 VTAIL.n2 VSUBS 0.014538f
C44 VTAIL.n3 VSUBS 0.034362f
C45 VTAIL.n4 VSUBS 0.015393f
C46 VTAIL.n5 VSUBS 0.027054f
C47 VTAIL.n6 VSUBS 0.014538f
C48 VTAIL.n7 VSUBS 0.034362f
C49 VTAIL.n8 VSUBS 0.015393f
C50 VTAIL.n9 VSUBS 0.761091f
C51 VTAIL.n10 VSUBS 0.014538f
C52 VTAIL.t1 VSUBS 0.073801f
C53 VTAIL.n11 VSUBS 0.154631f
C54 VTAIL.n12 VSUBS 0.025848f
C55 VTAIL.n13 VSUBS 0.025771f
C56 VTAIL.n14 VSUBS 0.034362f
C57 VTAIL.n15 VSUBS 0.015393f
C58 VTAIL.n16 VSUBS 0.014538f
C59 VTAIL.n17 VSUBS 0.027054f
C60 VTAIL.n18 VSUBS 0.027054f
C61 VTAIL.n19 VSUBS 0.014538f
C62 VTAIL.n20 VSUBS 0.015393f
C63 VTAIL.n21 VSUBS 0.034362f
C64 VTAIL.n22 VSUBS 0.034362f
C65 VTAIL.n23 VSUBS 0.015393f
C66 VTAIL.n24 VSUBS 0.014538f
C67 VTAIL.n25 VSUBS 0.027054f
C68 VTAIL.n26 VSUBS 0.027054f
C69 VTAIL.n27 VSUBS 0.014538f
C70 VTAIL.n28 VSUBS 0.015393f
C71 VTAIL.n29 VSUBS 0.034362f
C72 VTAIL.n30 VSUBS 0.084794f
C73 VTAIL.n31 VSUBS 0.015393f
C74 VTAIL.n32 VSUBS 0.028549f
C75 VTAIL.n33 VSUBS 0.067339f
C76 VTAIL.n34 VSUBS 0.06465f
C77 VTAIL.n35 VSUBS 0.211256f
C78 VTAIL.n36 VSUBS 0.028838f
C79 VTAIL.n37 VSUBS 0.027054f
C80 VTAIL.n38 VSUBS 0.014538f
C81 VTAIL.n39 VSUBS 0.034362f
C82 VTAIL.n40 VSUBS 0.015393f
C83 VTAIL.n41 VSUBS 0.027054f
C84 VTAIL.n42 VSUBS 0.014538f
C85 VTAIL.n43 VSUBS 0.034362f
C86 VTAIL.n44 VSUBS 0.015393f
C87 VTAIL.n45 VSUBS 0.761091f
C88 VTAIL.n46 VSUBS 0.014538f
C89 VTAIL.t4 VSUBS 0.073801f
C90 VTAIL.n47 VSUBS 0.154631f
C91 VTAIL.n48 VSUBS 0.025848f
C92 VTAIL.n49 VSUBS 0.025771f
C93 VTAIL.n50 VSUBS 0.034362f
C94 VTAIL.n51 VSUBS 0.015393f
C95 VTAIL.n52 VSUBS 0.014538f
C96 VTAIL.n53 VSUBS 0.027054f
C97 VTAIL.n54 VSUBS 0.027054f
C98 VTAIL.n55 VSUBS 0.014538f
C99 VTAIL.n56 VSUBS 0.015393f
C100 VTAIL.n57 VSUBS 0.034362f
C101 VTAIL.n58 VSUBS 0.034362f
C102 VTAIL.n59 VSUBS 0.015393f
C103 VTAIL.n60 VSUBS 0.014538f
C104 VTAIL.n61 VSUBS 0.027054f
C105 VTAIL.n62 VSUBS 0.027054f
C106 VTAIL.n63 VSUBS 0.014538f
C107 VTAIL.n64 VSUBS 0.015393f
C108 VTAIL.n65 VSUBS 0.034362f
C109 VTAIL.n66 VSUBS 0.084794f
C110 VTAIL.n67 VSUBS 0.015393f
C111 VTAIL.n68 VSUBS 0.028549f
C112 VTAIL.n69 VSUBS 0.067339f
C113 VTAIL.n70 VSUBS 0.06465f
C114 VTAIL.n71 VSUBS 0.345587f
C115 VTAIL.n72 VSUBS 0.028838f
C116 VTAIL.n73 VSUBS 0.027054f
C117 VTAIL.n74 VSUBS 0.014538f
C118 VTAIL.n75 VSUBS 0.034362f
C119 VTAIL.n76 VSUBS 0.015393f
C120 VTAIL.n77 VSUBS 0.027054f
C121 VTAIL.n78 VSUBS 0.014538f
C122 VTAIL.n79 VSUBS 0.034362f
C123 VTAIL.n80 VSUBS 0.015393f
C124 VTAIL.n81 VSUBS 0.761091f
C125 VTAIL.n82 VSUBS 0.014538f
C126 VTAIL.t5 VSUBS 0.073801f
C127 VTAIL.n83 VSUBS 0.154631f
C128 VTAIL.n84 VSUBS 0.025848f
C129 VTAIL.n85 VSUBS 0.025771f
C130 VTAIL.n86 VSUBS 0.034362f
C131 VTAIL.n87 VSUBS 0.015393f
C132 VTAIL.n88 VSUBS 0.014538f
C133 VTAIL.n89 VSUBS 0.027054f
C134 VTAIL.n90 VSUBS 0.027054f
C135 VTAIL.n91 VSUBS 0.014538f
C136 VTAIL.n92 VSUBS 0.015393f
C137 VTAIL.n93 VSUBS 0.034362f
C138 VTAIL.n94 VSUBS 0.034362f
C139 VTAIL.n95 VSUBS 0.015393f
C140 VTAIL.n96 VSUBS 0.014538f
C141 VTAIL.n97 VSUBS 0.027054f
C142 VTAIL.n98 VSUBS 0.027054f
C143 VTAIL.n99 VSUBS 0.014538f
C144 VTAIL.n100 VSUBS 0.015393f
C145 VTAIL.n101 VSUBS 0.034362f
C146 VTAIL.n102 VSUBS 0.084794f
C147 VTAIL.n103 VSUBS 0.015393f
C148 VTAIL.n104 VSUBS 0.028549f
C149 VTAIL.n105 VSUBS 0.067339f
C150 VTAIL.n106 VSUBS 0.06465f
C151 VTAIL.n107 VSUBS 1.49277f
C152 VTAIL.n108 VSUBS 0.028838f
C153 VTAIL.n109 VSUBS 0.027054f
C154 VTAIL.n110 VSUBS 0.014538f
C155 VTAIL.n111 VSUBS 0.034362f
C156 VTAIL.n112 VSUBS 0.015393f
C157 VTAIL.n113 VSUBS 0.027054f
C158 VTAIL.n114 VSUBS 0.014538f
C159 VTAIL.n115 VSUBS 0.034362f
C160 VTAIL.n116 VSUBS 0.015393f
C161 VTAIL.n117 VSUBS 0.761091f
C162 VTAIL.n118 VSUBS 0.014538f
C163 VTAIL.t2 VSUBS 0.073801f
C164 VTAIL.n119 VSUBS 0.154631f
C165 VTAIL.n120 VSUBS 0.025848f
C166 VTAIL.n121 VSUBS 0.025771f
C167 VTAIL.n122 VSUBS 0.034362f
C168 VTAIL.n123 VSUBS 0.015393f
C169 VTAIL.n124 VSUBS 0.014538f
C170 VTAIL.n125 VSUBS 0.027054f
C171 VTAIL.n126 VSUBS 0.027054f
C172 VTAIL.n127 VSUBS 0.014538f
C173 VTAIL.n128 VSUBS 0.015393f
C174 VTAIL.n129 VSUBS 0.034362f
C175 VTAIL.n130 VSUBS 0.034362f
C176 VTAIL.n131 VSUBS 0.015393f
C177 VTAIL.n132 VSUBS 0.014538f
C178 VTAIL.n133 VSUBS 0.027054f
C179 VTAIL.n134 VSUBS 0.027054f
C180 VTAIL.n135 VSUBS 0.014538f
C181 VTAIL.n136 VSUBS 0.015393f
C182 VTAIL.n137 VSUBS 0.034362f
C183 VTAIL.n138 VSUBS 0.084794f
C184 VTAIL.n139 VSUBS 0.015393f
C185 VTAIL.n140 VSUBS 0.028549f
C186 VTAIL.n141 VSUBS 0.067339f
C187 VTAIL.n142 VSUBS 0.06465f
C188 VTAIL.n143 VSUBS 1.49277f
C189 VTAIL.n144 VSUBS 0.028838f
C190 VTAIL.n145 VSUBS 0.027054f
C191 VTAIL.n146 VSUBS 0.014538f
C192 VTAIL.n147 VSUBS 0.034362f
C193 VTAIL.n148 VSUBS 0.015393f
C194 VTAIL.n149 VSUBS 0.027054f
C195 VTAIL.n150 VSUBS 0.014538f
C196 VTAIL.n151 VSUBS 0.034362f
C197 VTAIL.n152 VSUBS 0.015393f
C198 VTAIL.n153 VSUBS 0.761091f
C199 VTAIL.n154 VSUBS 0.014538f
C200 VTAIL.t0 VSUBS 0.073801f
C201 VTAIL.n155 VSUBS 0.154631f
C202 VTAIL.n156 VSUBS 0.025848f
C203 VTAIL.n157 VSUBS 0.025771f
C204 VTAIL.n158 VSUBS 0.034362f
C205 VTAIL.n159 VSUBS 0.015393f
C206 VTAIL.n160 VSUBS 0.014538f
C207 VTAIL.n161 VSUBS 0.027054f
C208 VTAIL.n162 VSUBS 0.027054f
C209 VTAIL.n163 VSUBS 0.014538f
C210 VTAIL.n164 VSUBS 0.015393f
C211 VTAIL.n165 VSUBS 0.034362f
C212 VTAIL.n166 VSUBS 0.034362f
C213 VTAIL.n167 VSUBS 0.015393f
C214 VTAIL.n168 VSUBS 0.014538f
C215 VTAIL.n169 VSUBS 0.027054f
C216 VTAIL.n170 VSUBS 0.027054f
C217 VTAIL.n171 VSUBS 0.014538f
C218 VTAIL.n172 VSUBS 0.015393f
C219 VTAIL.n173 VSUBS 0.034362f
C220 VTAIL.n174 VSUBS 0.084794f
C221 VTAIL.n175 VSUBS 0.015393f
C222 VTAIL.n176 VSUBS 0.028549f
C223 VTAIL.n177 VSUBS 0.067339f
C224 VTAIL.n178 VSUBS 0.06465f
C225 VTAIL.n179 VSUBS 0.345587f
C226 VTAIL.n180 VSUBS 0.028838f
C227 VTAIL.n181 VSUBS 0.027054f
C228 VTAIL.n182 VSUBS 0.014538f
C229 VTAIL.n183 VSUBS 0.034362f
C230 VTAIL.n184 VSUBS 0.015393f
C231 VTAIL.n185 VSUBS 0.027054f
C232 VTAIL.n186 VSUBS 0.014538f
C233 VTAIL.n187 VSUBS 0.034362f
C234 VTAIL.n188 VSUBS 0.015393f
C235 VTAIL.n189 VSUBS 0.761091f
C236 VTAIL.n190 VSUBS 0.014538f
C237 VTAIL.t7 VSUBS 0.073801f
C238 VTAIL.n191 VSUBS 0.154631f
C239 VTAIL.n192 VSUBS 0.025848f
C240 VTAIL.n193 VSUBS 0.025771f
C241 VTAIL.n194 VSUBS 0.034362f
C242 VTAIL.n195 VSUBS 0.015393f
C243 VTAIL.n196 VSUBS 0.014538f
C244 VTAIL.n197 VSUBS 0.027054f
C245 VTAIL.n198 VSUBS 0.027054f
C246 VTAIL.n199 VSUBS 0.014538f
C247 VTAIL.n200 VSUBS 0.015393f
C248 VTAIL.n201 VSUBS 0.034362f
C249 VTAIL.n202 VSUBS 0.034362f
C250 VTAIL.n203 VSUBS 0.015393f
C251 VTAIL.n204 VSUBS 0.014538f
C252 VTAIL.n205 VSUBS 0.027054f
C253 VTAIL.n206 VSUBS 0.027054f
C254 VTAIL.n207 VSUBS 0.014538f
C255 VTAIL.n208 VSUBS 0.015393f
C256 VTAIL.n209 VSUBS 0.034362f
C257 VTAIL.n210 VSUBS 0.084794f
C258 VTAIL.n211 VSUBS 0.015393f
C259 VTAIL.n212 VSUBS 0.028549f
C260 VTAIL.n213 VSUBS 0.067339f
C261 VTAIL.n214 VSUBS 0.06465f
C262 VTAIL.n215 VSUBS 0.345587f
C263 VTAIL.n216 VSUBS 0.028838f
C264 VTAIL.n217 VSUBS 0.027054f
C265 VTAIL.n218 VSUBS 0.014538f
C266 VTAIL.n219 VSUBS 0.034362f
C267 VTAIL.n220 VSUBS 0.015393f
C268 VTAIL.n221 VSUBS 0.027054f
C269 VTAIL.n222 VSUBS 0.014538f
C270 VTAIL.n223 VSUBS 0.034362f
C271 VTAIL.n224 VSUBS 0.015393f
C272 VTAIL.n225 VSUBS 0.761091f
C273 VTAIL.n226 VSUBS 0.014538f
C274 VTAIL.t6 VSUBS 0.073801f
C275 VTAIL.n227 VSUBS 0.154631f
C276 VTAIL.n228 VSUBS 0.025848f
C277 VTAIL.n229 VSUBS 0.025771f
C278 VTAIL.n230 VSUBS 0.034362f
C279 VTAIL.n231 VSUBS 0.015393f
C280 VTAIL.n232 VSUBS 0.014538f
C281 VTAIL.n233 VSUBS 0.027054f
C282 VTAIL.n234 VSUBS 0.027054f
C283 VTAIL.n235 VSUBS 0.014538f
C284 VTAIL.n236 VSUBS 0.015393f
C285 VTAIL.n237 VSUBS 0.034362f
C286 VTAIL.n238 VSUBS 0.034362f
C287 VTAIL.n239 VSUBS 0.015393f
C288 VTAIL.n240 VSUBS 0.014538f
C289 VTAIL.n241 VSUBS 0.027054f
C290 VTAIL.n242 VSUBS 0.027054f
C291 VTAIL.n243 VSUBS 0.014538f
C292 VTAIL.n244 VSUBS 0.015393f
C293 VTAIL.n245 VSUBS 0.034362f
C294 VTAIL.n246 VSUBS 0.084794f
C295 VTAIL.n247 VSUBS 0.015393f
C296 VTAIL.n248 VSUBS 0.028549f
C297 VTAIL.n249 VSUBS 0.067339f
C298 VTAIL.n250 VSUBS 0.06465f
C299 VTAIL.n251 VSUBS 1.49277f
C300 VTAIL.n252 VSUBS 0.028838f
C301 VTAIL.n253 VSUBS 0.027054f
C302 VTAIL.n254 VSUBS 0.014538f
C303 VTAIL.n255 VSUBS 0.034362f
C304 VTAIL.n256 VSUBS 0.015393f
C305 VTAIL.n257 VSUBS 0.027054f
C306 VTAIL.n258 VSUBS 0.014538f
C307 VTAIL.n259 VSUBS 0.034362f
C308 VTAIL.n260 VSUBS 0.015393f
C309 VTAIL.n261 VSUBS 0.761091f
C310 VTAIL.n262 VSUBS 0.014538f
C311 VTAIL.t3 VSUBS 0.073801f
C312 VTAIL.n263 VSUBS 0.154631f
C313 VTAIL.n264 VSUBS 0.025848f
C314 VTAIL.n265 VSUBS 0.025771f
C315 VTAIL.n266 VSUBS 0.034362f
C316 VTAIL.n267 VSUBS 0.015393f
C317 VTAIL.n268 VSUBS 0.014538f
C318 VTAIL.n269 VSUBS 0.027054f
C319 VTAIL.n270 VSUBS 0.027054f
C320 VTAIL.n271 VSUBS 0.014538f
C321 VTAIL.n272 VSUBS 0.015393f
C322 VTAIL.n273 VSUBS 0.034362f
C323 VTAIL.n274 VSUBS 0.034362f
C324 VTAIL.n275 VSUBS 0.015393f
C325 VTAIL.n276 VSUBS 0.014538f
C326 VTAIL.n277 VSUBS 0.027054f
C327 VTAIL.n278 VSUBS 0.027054f
C328 VTAIL.n279 VSUBS 0.014538f
C329 VTAIL.n280 VSUBS 0.015393f
C330 VTAIL.n281 VSUBS 0.034362f
C331 VTAIL.n282 VSUBS 0.084794f
C332 VTAIL.n283 VSUBS 0.015393f
C333 VTAIL.n284 VSUBS 0.028549f
C334 VTAIL.n285 VSUBS 0.067339f
C335 VTAIL.n286 VSUBS 0.06465f
C336 VTAIL.n287 VSUBS 1.34829f
C337 VDD1.t0 VSUBS 0.16207f
C338 VDD1.t3 VSUBS 0.16207f
C339 VDD1.n0 VSUBS 1.14768f
C340 VDD1.t1 VSUBS 0.16207f
C341 VDD1.t2 VSUBS 0.16207f
C342 VDD1.n1 VSUBS 1.70658f
C343 VP.t3 VSUBS 2.32625f
C344 VP.n0 VSUBS 0.995963f
C345 VP.n1 VSUBS 0.035712f
C346 VP.n2 VSUBS 0.02887f
C347 VP.n3 VSUBS 0.035712f
C348 VP.t2 VSUBS 2.32625f
C349 VP.n4 VSUBS 0.995963f
C350 VP.t0 VSUBS 2.78205f
C351 VP.t1 VSUBS 2.76796f
C352 VP.n5 VSUBS 3.64006f
C353 VP.n6 VSUBS 1.89045f
C354 VP.n7 VSUBS 0.057639f
C355 VP.n8 VSUBS 0.057028f
C356 VP.n9 VSUBS 0.066559f
C357 VP.n10 VSUBS 0.070978f
C358 VP.n11 VSUBS 0.035712f
C359 VP.n12 VSUBS 0.035712f
C360 VP.n13 VSUBS 0.035712f
C361 VP.n14 VSUBS 0.070978f
C362 VP.n15 VSUBS 0.066559f
C363 VP.n16 VSUBS 0.057028f
C364 VP.n17 VSUBS 0.057639f
C365 VP.n18 VSUBS 0.083377f
C366 B.n0 VSUBS 0.004737f
C367 B.n1 VSUBS 0.004737f
C368 B.n2 VSUBS 0.007491f
C369 B.n3 VSUBS 0.007491f
C370 B.n4 VSUBS 0.007491f
C371 B.n5 VSUBS 0.007491f
C372 B.n6 VSUBS 0.007491f
C373 B.n7 VSUBS 0.007491f
C374 B.n8 VSUBS 0.007491f
C375 B.n9 VSUBS 0.007491f
C376 B.n10 VSUBS 0.007491f
C377 B.n11 VSUBS 0.007491f
C378 B.n12 VSUBS 0.007491f
C379 B.n13 VSUBS 0.007491f
C380 B.n14 VSUBS 0.007491f
C381 B.n15 VSUBS 0.007491f
C382 B.n16 VSUBS 0.007491f
C383 B.n17 VSUBS 0.007491f
C384 B.n18 VSUBS 0.007491f
C385 B.n19 VSUBS 0.007491f
C386 B.n20 VSUBS 0.007491f
C387 B.n21 VSUBS 0.007491f
C388 B.n22 VSUBS 0.015693f
C389 B.n23 VSUBS 0.007491f
C390 B.n24 VSUBS 0.007491f
C391 B.n25 VSUBS 0.007491f
C392 B.n26 VSUBS 0.007491f
C393 B.n27 VSUBS 0.007491f
C394 B.n28 VSUBS 0.007491f
C395 B.n29 VSUBS 0.007491f
C396 B.n30 VSUBS 0.007491f
C397 B.n31 VSUBS 0.007491f
C398 B.n32 VSUBS 0.007491f
C399 B.n33 VSUBS 0.007491f
C400 B.n34 VSUBS 0.007491f
C401 B.n35 VSUBS 0.007491f
C402 B.n36 VSUBS 0.005178f
C403 B.n37 VSUBS 0.007491f
C404 B.t11 VSUBS 0.119018f
C405 B.t10 VSUBS 0.155608f
C406 B.t9 VSUBS 1.23869f
C407 B.n38 VSUBS 0.2568f
C408 B.n39 VSUBS 0.194436f
C409 B.n40 VSUBS 0.017356f
C410 B.n41 VSUBS 0.007491f
C411 B.n42 VSUBS 0.007491f
C412 B.n43 VSUBS 0.007491f
C413 B.n44 VSUBS 0.007491f
C414 B.t8 VSUBS 0.11902f
C415 B.t7 VSUBS 0.15561f
C416 B.t6 VSUBS 1.23869f
C417 B.n45 VSUBS 0.256798f
C418 B.n46 VSUBS 0.194434f
C419 B.n47 VSUBS 0.007491f
C420 B.n48 VSUBS 0.007491f
C421 B.n49 VSUBS 0.007491f
C422 B.n50 VSUBS 0.007491f
C423 B.n51 VSUBS 0.007491f
C424 B.n52 VSUBS 0.007491f
C425 B.n53 VSUBS 0.007491f
C426 B.n54 VSUBS 0.007491f
C427 B.n55 VSUBS 0.007491f
C428 B.n56 VSUBS 0.007491f
C429 B.n57 VSUBS 0.007491f
C430 B.n58 VSUBS 0.007491f
C431 B.n59 VSUBS 0.007491f
C432 B.n60 VSUBS 0.015693f
C433 B.n61 VSUBS 0.007491f
C434 B.n62 VSUBS 0.007491f
C435 B.n63 VSUBS 0.007491f
C436 B.n64 VSUBS 0.007491f
C437 B.n65 VSUBS 0.007491f
C438 B.n66 VSUBS 0.007491f
C439 B.n67 VSUBS 0.007491f
C440 B.n68 VSUBS 0.007491f
C441 B.n69 VSUBS 0.007491f
C442 B.n70 VSUBS 0.007491f
C443 B.n71 VSUBS 0.007491f
C444 B.n72 VSUBS 0.007491f
C445 B.n73 VSUBS 0.007491f
C446 B.n74 VSUBS 0.007491f
C447 B.n75 VSUBS 0.007491f
C448 B.n76 VSUBS 0.007491f
C449 B.n77 VSUBS 0.007491f
C450 B.n78 VSUBS 0.007491f
C451 B.n79 VSUBS 0.007491f
C452 B.n80 VSUBS 0.007491f
C453 B.n81 VSUBS 0.007491f
C454 B.n82 VSUBS 0.007491f
C455 B.n83 VSUBS 0.007491f
C456 B.n84 VSUBS 0.007491f
C457 B.n85 VSUBS 0.007491f
C458 B.n86 VSUBS 0.007491f
C459 B.n87 VSUBS 0.007491f
C460 B.n88 VSUBS 0.007491f
C461 B.n89 VSUBS 0.007491f
C462 B.n90 VSUBS 0.007491f
C463 B.n91 VSUBS 0.007491f
C464 B.n92 VSUBS 0.007491f
C465 B.n93 VSUBS 0.007491f
C466 B.n94 VSUBS 0.007491f
C467 B.n95 VSUBS 0.007491f
C468 B.n96 VSUBS 0.007491f
C469 B.n97 VSUBS 0.007491f
C470 B.n98 VSUBS 0.007491f
C471 B.n99 VSUBS 0.007491f
C472 B.n100 VSUBS 0.007491f
C473 B.n101 VSUBS 0.015693f
C474 B.n102 VSUBS 0.007491f
C475 B.n103 VSUBS 0.007491f
C476 B.n104 VSUBS 0.007491f
C477 B.n105 VSUBS 0.007491f
C478 B.n106 VSUBS 0.007491f
C479 B.n107 VSUBS 0.007491f
C480 B.n108 VSUBS 0.007491f
C481 B.n109 VSUBS 0.007491f
C482 B.n110 VSUBS 0.007491f
C483 B.n111 VSUBS 0.007491f
C484 B.n112 VSUBS 0.007491f
C485 B.n113 VSUBS 0.007491f
C486 B.n114 VSUBS 0.007491f
C487 B.n115 VSUBS 0.005178f
C488 B.n116 VSUBS 0.007491f
C489 B.n117 VSUBS 0.007491f
C490 B.n118 VSUBS 0.007491f
C491 B.n119 VSUBS 0.007491f
C492 B.n120 VSUBS 0.007491f
C493 B.t1 VSUBS 0.119018f
C494 B.t2 VSUBS 0.155608f
C495 B.t0 VSUBS 1.23869f
C496 B.n121 VSUBS 0.2568f
C497 B.n122 VSUBS 0.194436f
C498 B.n123 VSUBS 0.007491f
C499 B.n124 VSUBS 0.007491f
C500 B.n125 VSUBS 0.007491f
C501 B.n126 VSUBS 0.007491f
C502 B.n127 VSUBS 0.007491f
C503 B.n128 VSUBS 0.007491f
C504 B.n129 VSUBS 0.007491f
C505 B.n130 VSUBS 0.007491f
C506 B.n131 VSUBS 0.007491f
C507 B.n132 VSUBS 0.007491f
C508 B.n133 VSUBS 0.007491f
C509 B.n134 VSUBS 0.007491f
C510 B.n135 VSUBS 0.007491f
C511 B.n136 VSUBS 0.015693f
C512 B.n137 VSUBS 0.007491f
C513 B.n138 VSUBS 0.007491f
C514 B.n139 VSUBS 0.007491f
C515 B.n140 VSUBS 0.007491f
C516 B.n141 VSUBS 0.007491f
C517 B.n142 VSUBS 0.007491f
C518 B.n143 VSUBS 0.007491f
C519 B.n144 VSUBS 0.007491f
C520 B.n145 VSUBS 0.007491f
C521 B.n146 VSUBS 0.007491f
C522 B.n147 VSUBS 0.007491f
C523 B.n148 VSUBS 0.007491f
C524 B.n149 VSUBS 0.007491f
C525 B.n150 VSUBS 0.007491f
C526 B.n151 VSUBS 0.007491f
C527 B.n152 VSUBS 0.007491f
C528 B.n153 VSUBS 0.007491f
C529 B.n154 VSUBS 0.007491f
C530 B.n155 VSUBS 0.007491f
C531 B.n156 VSUBS 0.007491f
C532 B.n157 VSUBS 0.007491f
C533 B.n158 VSUBS 0.007491f
C534 B.n159 VSUBS 0.007491f
C535 B.n160 VSUBS 0.007491f
C536 B.n161 VSUBS 0.007491f
C537 B.n162 VSUBS 0.007491f
C538 B.n163 VSUBS 0.007491f
C539 B.n164 VSUBS 0.007491f
C540 B.n165 VSUBS 0.007491f
C541 B.n166 VSUBS 0.007491f
C542 B.n167 VSUBS 0.007491f
C543 B.n168 VSUBS 0.007491f
C544 B.n169 VSUBS 0.007491f
C545 B.n170 VSUBS 0.007491f
C546 B.n171 VSUBS 0.007491f
C547 B.n172 VSUBS 0.007491f
C548 B.n173 VSUBS 0.007491f
C549 B.n174 VSUBS 0.007491f
C550 B.n175 VSUBS 0.007491f
C551 B.n176 VSUBS 0.007491f
C552 B.n177 VSUBS 0.007491f
C553 B.n178 VSUBS 0.007491f
C554 B.n179 VSUBS 0.007491f
C555 B.n180 VSUBS 0.007491f
C556 B.n181 VSUBS 0.007491f
C557 B.n182 VSUBS 0.007491f
C558 B.n183 VSUBS 0.007491f
C559 B.n184 VSUBS 0.007491f
C560 B.n185 VSUBS 0.007491f
C561 B.n186 VSUBS 0.007491f
C562 B.n187 VSUBS 0.007491f
C563 B.n188 VSUBS 0.007491f
C564 B.n189 VSUBS 0.007491f
C565 B.n190 VSUBS 0.007491f
C566 B.n191 VSUBS 0.007491f
C567 B.n192 VSUBS 0.007491f
C568 B.n193 VSUBS 0.007491f
C569 B.n194 VSUBS 0.007491f
C570 B.n195 VSUBS 0.007491f
C571 B.n196 VSUBS 0.007491f
C572 B.n197 VSUBS 0.007491f
C573 B.n198 VSUBS 0.007491f
C574 B.n199 VSUBS 0.007491f
C575 B.n200 VSUBS 0.007491f
C576 B.n201 VSUBS 0.007491f
C577 B.n202 VSUBS 0.007491f
C578 B.n203 VSUBS 0.007491f
C579 B.n204 VSUBS 0.007491f
C580 B.n205 VSUBS 0.007491f
C581 B.n206 VSUBS 0.007491f
C582 B.n207 VSUBS 0.007491f
C583 B.n208 VSUBS 0.007491f
C584 B.n209 VSUBS 0.007491f
C585 B.n210 VSUBS 0.007491f
C586 B.n211 VSUBS 0.007491f
C587 B.n212 VSUBS 0.007491f
C588 B.n213 VSUBS 0.007491f
C589 B.n214 VSUBS 0.007491f
C590 B.n215 VSUBS 0.015693f
C591 B.n216 VSUBS 0.016694f
C592 B.n217 VSUBS 0.016694f
C593 B.n218 VSUBS 0.007491f
C594 B.n219 VSUBS 0.007491f
C595 B.n220 VSUBS 0.007491f
C596 B.n221 VSUBS 0.007491f
C597 B.n222 VSUBS 0.007491f
C598 B.n223 VSUBS 0.007491f
C599 B.n224 VSUBS 0.007491f
C600 B.n225 VSUBS 0.007491f
C601 B.n226 VSUBS 0.007491f
C602 B.n227 VSUBS 0.007491f
C603 B.n228 VSUBS 0.007491f
C604 B.n229 VSUBS 0.007491f
C605 B.n230 VSUBS 0.007491f
C606 B.n231 VSUBS 0.007491f
C607 B.n232 VSUBS 0.007491f
C608 B.n233 VSUBS 0.007491f
C609 B.n234 VSUBS 0.007491f
C610 B.n235 VSUBS 0.007491f
C611 B.n236 VSUBS 0.007491f
C612 B.n237 VSUBS 0.007491f
C613 B.n238 VSUBS 0.007491f
C614 B.n239 VSUBS 0.007491f
C615 B.n240 VSUBS 0.007491f
C616 B.n241 VSUBS 0.007491f
C617 B.n242 VSUBS 0.007491f
C618 B.n243 VSUBS 0.007491f
C619 B.n244 VSUBS 0.007491f
C620 B.n245 VSUBS 0.007491f
C621 B.n246 VSUBS 0.007491f
C622 B.n247 VSUBS 0.007491f
C623 B.n248 VSUBS 0.007491f
C624 B.n249 VSUBS 0.007491f
C625 B.n250 VSUBS 0.007491f
C626 B.n251 VSUBS 0.007491f
C627 B.n252 VSUBS 0.007491f
C628 B.n253 VSUBS 0.007491f
C629 B.n254 VSUBS 0.007491f
C630 B.n255 VSUBS 0.007491f
C631 B.n256 VSUBS 0.007491f
C632 B.n257 VSUBS 0.005178f
C633 B.n258 VSUBS 0.017356f
C634 B.n259 VSUBS 0.006059f
C635 B.n260 VSUBS 0.007491f
C636 B.n261 VSUBS 0.007491f
C637 B.n262 VSUBS 0.007491f
C638 B.n263 VSUBS 0.007491f
C639 B.n264 VSUBS 0.007491f
C640 B.n265 VSUBS 0.007491f
C641 B.n266 VSUBS 0.007491f
C642 B.n267 VSUBS 0.007491f
C643 B.n268 VSUBS 0.007491f
C644 B.n269 VSUBS 0.007491f
C645 B.n270 VSUBS 0.007491f
C646 B.t4 VSUBS 0.11902f
C647 B.t5 VSUBS 0.15561f
C648 B.t3 VSUBS 1.23869f
C649 B.n271 VSUBS 0.256798f
C650 B.n272 VSUBS 0.194434f
C651 B.n273 VSUBS 0.017356f
C652 B.n274 VSUBS 0.006059f
C653 B.n275 VSUBS 0.007491f
C654 B.n276 VSUBS 0.007491f
C655 B.n277 VSUBS 0.007491f
C656 B.n278 VSUBS 0.007491f
C657 B.n279 VSUBS 0.007491f
C658 B.n280 VSUBS 0.007491f
C659 B.n281 VSUBS 0.007491f
C660 B.n282 VSUBS 0.007491f
C661 B.n283 VSUBS 0.007491f
C662 B.n284 VSUBS 0.007491f
C663 B.n285 VSUBS 0.007491f
C664 B.n286 VSUBS 0.007491f
C665 B.n287 VSUBS 0.007491f
C666 B.n288 VSUBS 0.007491f
C667 B.n289 VSUBS 0.007491f
C668 B.n290 VSUBS 0.007491f
C669 B.n291 VSUBS 0.007491f
C670 B.n292 VSUBS 0.007491f
C671 B.n293 VSUBS 0.007491f
C672 B.n294 VSUBS 0.007491f
C673 B.n295 VSUBS 0.007491f
C674 B.n296 VSUBS 0.007491f
C675 B.n297 VSUBS 0.007491f
C676 B.n298 VSUBS 0.007491f
C677 B.n299 VSUBS 0.007491f
C678 B.n300 VSUBS 0.007491f
C679 B.n301 VSUBS 0.007491f
C680 B.n302 VSUBS 0.007491f
C681 B.n303 VSUBS 0.007491f
C682 B.n304 VSUBS 0.007491f
C683 B.n305 VSUBS 0.007491f
C684 B.n306 VSUBS 0.007491f
C685 B.n307 VSUBS 0.007491f
C686 B.n308 VSUBS 0.007491f
C687 B.n309 VSUBS 0.007491f
C688 B.n310 VSUBS 0.007491f
C689 B.n311 VSUBS 0.007491f
C690 B.n312 VSUBS 0.007491f
C691 B.n313 VSUBS 0.007491f
C692 B.n314 VSUBS 0.007491f
C693 B.n315 VSUBS 0.007491f
C694 B.n316 VSUBS 0.016694f
C695 B.n317 VSUBS 0.016694f
C696 B.n318 VSUBS 0.015693f
C697 B.n319 VSUBS 0.007491f
C698 B.n320 VSUBS 0.007491f
C699 B.n321 VSUBS 0.007491f
C700 B.n322 VSUBS 0.007491f
C701 B.n323 VSUBS 0.007491f
C702 B.n324 VSUBS 0.007491f
C703 B.n325 VSUBS 0.007491f
C704 B.n326 VSUBS 0.007491f
C705 B.n327 VSUBS 0.007491f
C706 B.n328 VSUBS 0.007491f
C707 B.n329 VSUBS 0.007491f
C708 B.n330 VSUBS 0.007491f
C709 B.n331 VSUBS 0.007491f
C710 B.n332 VSUBS 0.007491f
C711 B.n333 VSUBS 0.007491f
C712 B.n334 VSUBS 0.007491f
C713 B.n335 VSUBS 0.007491f
C714 B.n336 VSUBS 0.007491f
C715 B.n337 VSUBS 0.007491f
C716 B.n338 VSUBS 0.007491f
C717 B.n339 VSUBS 0.007491f
C718 B.n340 VSUBS 0.007491f
C719 B.n341 VSUBS 0.007491f
C720 B.n342 VSUBS 0.007491f
C721 B.n343 VSUBS 0.007491f
C722 B.n344 VSUBS 0.007491f
C723 B.n345 VSUBS 0.007491f
C724 B.n346 VSUBS 0.007491f
C725 B.n347 VSUBS 0.007491f
C726 B.n348 VSUBS 0.007491f
C727 B.n349 VSUBS 0.007491f
C728 B.n350 VSUBS 0.007491f
C729 B.n351 VSUBS 0.007491f
C730 B.n352 VSUBS 0.007491f
C731 B.n353 VSUBS 0.007491f
C732 B.n354 VSUBS 0.007491f
C733 B.n355 VSUBS 0.007491f
C734 B.n356 VSUBS 0.007491f
C735 B.n357 VSUBS 0.007491f
C736 B.n358 VSUBS 0.007491f
C737 B.n359 VSUBS 0.007491f
C738 B.n360 VSUBS 0.007491f
C739 B.n361 VSUBS 0.007491f
C740 B.n362 VSUBS 0.007491f
C741 B.n363 VSUBS 0.007491f
C742 B.n364 VSUBS 0.007491f
C743 B.n365 VSUBS 0.007491f
C744 B.n366 VSUBS 0.007491f
C745 B.n367 VSUBS 0.007491f
C746 B.n368 VSUBS 0.007491f
C747 B.n369 VSUBS 0.007491f
C748 B.n370 VSUBS 0.007491f
C749 B.n371 VSUBS 0.007491f
C750 B.n372 VSUBS 0.007491f
C751 B.n373 VSUBS 0.007491f
C752 B.n374 VSUBS 0.007491f
C753 B.n375 VSUBS 0.007491f
C754 B.n376 VSUBS 0.007491f
C755 B.n377 VSUBS 0.007491f
C756 B.n378 VSUBS 0.007491f
C757 B.n379 VSUBS 0.007491f
C758 B.n380 VSUBS 0.007491f
C759 B.n381 VSUBS 0.007491f
C760 B.n382 VSUBS 0.007491f
C761 B.n383 VSUBS 0.007491f
C762 B.n384 VSUBS 0.007491f
C763 B.n385 VSUBS 0.007491f
C764 B.n386 VSUBS 0.007491f
C765 B.n387 VSUBS 0.007491f
C766 B.n388 VSUBS 0.007491f
C767 B.n389 VSUBS 0.007491f
C768 B.n390 VSUBS 0.007491f
C769 B.n391 VSUBS 0.007491f
C770 B.n392 VSUBS 0.007491f
C771 B.n393 VSUBS 0.007491f
C772 B.n394 VSUBS 0.007491f
C773 B.n395 VSUBS 0.007491f
C774 B.n396 VSUBS 0.007491f
C775 B.n397 VSUBS 0.007491f
C776 B.n398 VSUBS 0.007491f
C777 B.n399 VSUBS 0.007491f
C778 B.n400 VSUBS 0.007491f
C779 B.n401 VSUBS 0.007491f
C780 B.n402 VSUBS 0.007491f
C781 B.n403 VSUBS 0.007491f
C782 B.n404 VSUBS 0.007491f
C783 B.n405 VSUBS 0.007491f
C784 B.n406 VSUBS 0.007491f
C785 B.n407 VSUBS 0.007491f
C786 B.n408 VSUBS 0.007491f
C787 B.n409 VSUBS 0.007491f
C788 B.n410 VSUBS 0.007491f
C789 B.n411 VSUBS 0.007491f
C790 B.n412 VSUBS 0.007491f
C791 B.n413 VSUBS 0.007491f
C792 B.n414 VSUBS 0.007491f
C793 B.n415 VSUBS 0.007491f
C794 B.n416 VSUBS 0.007491f
C795 B.n417 VSUBS 0.007491f
C796 B.n418 VSUBS 0.007491f
C797 B.n419 VSUBS 0.007491f
C798 B.n420 VSUBS 0.007491f
C799 B.n421 VSUBS 0.007491f
C800 B.n422 VSUBS 0.007491f
C801 B.n423 VSUBS 0.007491f
C802 B.n424 VSUBS 0.007491f
C803 B.n425 VSUBS 0.007491f
C804 B.n426 VSUBS 0.007491f
C805 B.n427 VSUBS 0.007491f
C806 B.n428 VSUBS 0.007491f
C807 B.n429 VSUBS 0.007491f
C808 B.n430 VSUBS 0.007491f
C809 B.n431 VSUBS 0.007491f
C810 B.n432 VSUBS 0.007491f
C811 B.n433 VSUBS 0.007491f
C812 B.n434 VSUBS 0.007491f
C813 B.n435 VSUBS 0.007491f
C814 B.n436 VSUBS 0.007491f
C815 B.n437 VSUBS 0.007491f
C816 B.n438 VSUBS 0.007491f
C817 B.n439 VSUBS 0.007491f
C818 B.n440 VSUBS 0.007491f
C819 B.n441 VSUBS 0.016694f
C820 B.n442 VSUBS 0.015693f
C821 B.n443 VSUBS 0.016694f
C822 B.n444 VSUBS 0.007491f
C823 B.n445 VSUBS 0.007491f
C824 B.n446 VSUBS 0.007491f
C825 B.n447 VSUBS 0.007491f
C826 B.n448 VSUBS 0.007491f
C827 B.n449 VSUBS 0.007491f
C828 B.n450 VSUBS 0.007491f
C829 B.n451 VSUBS 0.007491f
C830 B.n452 VSUBS 0.007491f
C831 B.n453 VSUBS 0.007491f
C832 B.n454 VSUBS 0.007491f
C833 B.n455 VSUBS 0.007491f
C834 B.n456 VSUBS 0.007491f
C835 B.n457 VSUBS 0.007491f
C836 B.n458 VSUBS 0.007491f
C837 B.n459 VSUBS 0.007491f
C838 B.n460 VSUBS 0.007491f
C839 B.n461 VSUBS 0.007491f
C840 B.n462 VSUBS 0.007491f
C841 B.n463 VSUBS 0.007491f
C842 B.n464 VSUBS 0.007491f
C843 B.n465 VSUBS 0.007491f
C844 B.n466 VSUBS 0.007491f
C845 B.n467 VSUBS 0.007491f
C846 B.n468 VSUBS 0.007491f
C847 B.n469 VSUBS 0.007491f
C848 B.n470 VSUBS 0.007491f
C849 B.n471 VSUBS 0.007491f
C850 B.n472 VSUBS 0.007491f
C851 B.n473 VSUBS 0.007491f
C852 B.n474 VSUBS 0.007491f
C853 B.n475 VSUBS 0.007491f
C854 B.n476 VSUBS 0.007491f
C855 B.n477 VSUBS 0.007491f
C856 B.n478 VSUBS 0.007491f
C857 B.n479 VSUBS 0.007491f
C858 B.n480 VSUBS 0.007491f
C859 B.n481 VSUBS 0.007491f
C860 B.n482 VSUBS 0.007491f
C861 B.n483 VSUBS 0.005178f
C862 B.n484 VSUBS 0.017356f
C863 B.n485 VSUBS 0.006059f
C864 B.n486 VSUBS 0.007491f
C865 B.n487 VSUBS 0.007491f
C866 B.n488 VSUBS 0.007491f
C867 B.n489 VSUBS 0.007491f
C868 B.n490 VSUBS 0.007491f
C869 B.n491 VSUBS 0.007491f
C870 B.n492 VSUBS 0.007491f
C871 B.n493 VSUBS 0.007491f
C872 B.n494 VSUBS 0.007491f
C873 B.n495 VSUBS 0.007491f
C874 B.n496 VSUBS 0.007491f
C875 B.n497 VSUBS 0.006059f
C876 B.n498 VSUBS 0.007491f
C877 B.n499 VSUBS 0.007491f
C878 B.n500 VSUBS 0.007491f
C879 B.n501 VSUBS 0.007491f
C880 B.n502 VSUBS 0.007491f
C881 B.n503 VSUBS 0.007491f
C882 B.n504 VSUBS 0.007491f
C883 B.n505 VSUBS 0.007491f
C884 B.n506 VSUBS 0.007491f
C885 B.n507 VSUBS 0.007491f
C886 B.n508 VSUBS 0.007491f
C887 B.n509 VSUBS 0.007491f
C888 B.n510 VSUBS 0.007491f
C889 B.n511 VSUBS 0.007491f
C890 B.n512 VSUBS 0.007491f
C891 B.n513 VSUBS 0.007491f
C892 B.n514 VSUBS 0.007491f
C893 B.n515 VSUBS 0.007491f
C894 B.n516 VSUBS 0.007491f
C895 B.n517 VSUBS 0.007491f
C896 B.n518 VSUBS 0.007491f
C897 B.n519 VSUBS 0.007491f
C898 B.n520 VSUBS 0.007491f
C899 B.n521 VSUBS 0.007491f
C900 B.n522 VSUBS 0.007491f
C901 B.n523 VSUBS 0.007491f
C902 B.n524 VSUBS 0.007491f
C903 B.n525 VSUBS 0.007491f
C904 B.n526 VSUBS 0.007491f
C905 B.n527 VSUBS 0.007491f
C906 B.n528 VSUBS 0.007491f
C907 B.n529 VSUBS 0.007491f
C908 B.n530 VSUBS 0.007491f
C909 B.n531 VSUBS 0.007491f
C910 B.n532 VSUBS 0.007491f
C911 B.n533 VSUBS 0.007491f
C912 B.n534 VSUBS 0.007491f
C913 B.n535 VSUBS 0.007491f
C914 B.n536 VSUBS 0.007491f
C915 B.n537 VSUBS 0.007491f
C916 B.n538 VSUBS 0.007491f
C917 B.n539 VSUBS 0.016694f
C918 B.n540 VSUBS 0.016694f
C919 B.n541 VSUBS 0.015693f
C920 B.n542 VSUBS 0.007491f
C921 B.n543 VSUBS 0.007491f
C922 B.n544 VSUBS 0.007491f
C923 B.n545 VSUBS 0.007491f
C924 B.n546 VSUBS 0.007491f
C925 B.n547 VSUBS 0.007491f
C926 B.n548 VSUBS 0.007491f
C927 B.n549 VSUBS 0.007491f
C928 B.n550 VSUBS 0.007491f
C929 B.n551 VSUBS 0.007491f
C930 B.n552 VSUBS 0.007491f
C931 B.n553 VSUBS 0.007491f
C932 B.n554 VSUBS 0.007491f
C933 B.n555 VSUBS 0.007491f
C934 B.n556 VSUBS 0.007491f
C935 B.n557 VSUBS 0.007491f
C936 B.n558 VSUBS 0.007491f
C937 B.n559 VSUBS 0.007491f
C938 B.n560 VSUBS 0.007491f
C939 B.n561 VSUBS 0.007491f
C940 B.n562 VSUBS 0.007491f
C941 B.n563 VSUBS 0.007491f
C942 B.n564 VSUBS 0.007491f
C943 B.n565 VSUBS 0.007491f
C944 B.n566 VSUBS 0.007491f
C945 B.n567 VSUBS 0.007491f
C946 B.n568 VSUBS 0.007491f
C947 B.n569 VSUBS 0.007491f
C948 B.n570 VSUBS 0.007491f
C949 B.n571 VSUBS 0.007491f
C950 B.n572 VSUBS 0.007491f
C951 B.n573 VSUBS 0.007491f
C952 B.n574 VSUBS 0.007491f
C953 B.n575 VSUBS 0.007491f
C954 B.n576 VSUBS 0.007491f
C955 B.n577 VSUBS 0.007491f
C956 B.n578 VSUBS 0.007491f
C957 B.n579 VSUBS 0.007491f
C958 B.n580 VSUBS 0.007491f
C959 B.n581 VSUBS 0.007491f
C960 B.n582 VSUBS 0.007491f
C961 B.n583 VSUBS 0.007491f
C962 B.n584 VSUBS 0.007491f
C963 B.n585 VSUBS 0.007491f
C964 B.n586 VSUBS 0.007491f
C965 B.n587 VSUBS 0.007491f
C966 B.n588 VSUBS 0.007491f
C967 B.n589 VSUBS 0.007491f
C968 B.n590 VSUBS 0.007491f
C969 B.n591 VSUBS 0.007491f
C970 B.n592 VSUBS 0.007491f
C971 B.n593 VSUBS 0.007491f
C972 B.n594 VSUBS 0.007491f
C973 B.n595 VSUBS 0.007491f
C974 B.n596 VSUBS 0.007491f
C975 B.n597 VSUBS 0.007491f
C976 B.n598 VSUBS 0.007491f
C977 B.n599 VSUBS 0.007491f
C978 B.n600 VSUBS 0.007491f
C979 B.n601 VSUBS 0.007491f
C980 B.n602 VSUBS 0.007491f
C981 B.n603 VSUBS 0.016962f
.ends

