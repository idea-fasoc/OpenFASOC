* NGSPICE file created from diff_pair_sample_1080.ext - technology: sky130A

.subckt diff_pair_sample_1080 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t0 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=6.3414 ps=33.3 w=16.26 l=2.59
X1 VDD2.t1 VN.t0 VTAIL.t2 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=6.3414 ps=33.3 w=16.26 l=2.59
X2 B.t11 B.t9 B.t10 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=0 ps=0 w=16.26 l=2.59
X3 VDD2.t0 VN.t1 VTAIL.t3 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=6.3414 ps=33.3 w=16.26 l=2.59
X4 B.t8 B.t6 B.t7 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=0 ps=0 w=16.26 l=2.59
X5 B.t5 B.t3 B.t4 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=0 ps=0 w=16.26 l=2.59
X6 B.t2 B.t0 B.t1 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=0 ps=0 w=16.26 l=2.59
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n2138_n4220# sky130_fd_pr__pfet_01v8 ad=6.3414 pd=33.3 as=6.3414 ps=33.3 w=16.26 l=2.59
R0 VP.n0 VP.t1 248.284
R1 VP.n0 VP.t0 200.427
R2 VP VP.n0 0.336784
R3 VTAIL.n354 VTAIL.n270 756.745
R4 VTAIL.n84 VTAIL.n0 756.745
R5 VTAIL.n264 VTAIL.n180 756.745
R6 VTAIL.n174 VTAIL.n90 756.745
R7 VTAIL.n298 VTAIL.n297 585
R8 VTAIL.n303 VTAIL.n302 585
R9 VTAIL.n305 VTAIL.n304 585
R10 VTAIL.n294 VTAIL.n293 585
R11 VTAIL.n311 VTAIL.n310 585
R12 VTAIL.n313 VTAIL.n312 585
R13 VTAIL.n290 VTAIL.n289 585
R14 VTAIL.n319 VTAIL.n318 585
R15 VTAIL.n321 VTAIL.n320 585
R16 VTAIL.n286 VTAIL.n285 585
R17 VTAIL.n327 VTAIL.n326 585
R18 VTAIL.n329 VTAIL.n328 585
R19 VTAIL.n282 VTAIL.n281 585
R20 VTAIL.n335 VTAIL.n334 585
R21 VTAIL.n337 VTAIL.n336 585
R22 VTAIL.n278 VTAIL.n277 585
R23 VTAIL.n344 VTAIL.n343 585
R24 VTAIL.n345 VTAIL.n276 585
R25 VTAIL.n347 VTAIL.n346 585
R26 VTAIL.n274 VTAIL.n273 585
R27 VTAIL.n353 VTAIL.n352 585
R28 VTAIL.n355 VTAIL.n354 585
R29 VTAIL.n28 VTAIL.n27 585
R30 VTAIL.n33 VTAIL.n32 585
R31 VTAIL.n35 VTAIL.n34 585
R32 VTAIL.n24 VTAIL.n23 585
R33 VTAIL.n41 VTAIL.n40 585
R34 VTAIL.n43 VTAIL.n42 585
R35 VTAIL.n20 VTAIL.n19 585
R36 VTAIL.n49 VTAIL.n48 585
R37 VTAIL.n51 VTAIL.n50 585
R38 VTAIL.n16 VTAIL.n15 585
R39 VTAIL.n57 VTAIL.n56 585
R40 VTAIL.n59 VTAIL.n58 585
R41 VTAIL.n12 VTAIL.n11 585
R42 VTAIL.n65 VTAIL.n64 585
R43 VTAIL.n67 VTAIL.n66 585
R44 VTAIL.n8 VTAIL.n7 585
R45 VTAIL.n74 VTAIL.n73 585
R46 VTAIL.n75 VTAIL.n6 585
R47 VTAIL.n77 VTAIL.n76 585
R48 VTAIL.n4 VTAIL.n3 585
R49 VTAIL.n83 VTAIL.n82 585
R50 VTAIL.n85 VTAIL.n84 585
R51 VTAIL.n265 VTAIL.n264 585
R52 VTAIL.n263 VTAIL.n262 585
R53 VTAIL.n184 VTAIL.n183 585
R54 VTAIL.n257 VTAIL.n256 585
R55 VTAIL.n255 VTAIL.n186 585
R56 VTAIL.n254 VTAIL.n253 585
R57 VTAIL.n189 VTAIL.n187 585
R58 VTAIL.n248 VTAIL.n247 585
R59 VTAIL.n246 VTAIL.n245 585
R60 VTAIL.n193 VTAIL.n192 585
R61 VTAIL.n240 VTAIL.n239 585
R62 VTAIL.n238 VTAIL.n237 585
R63 VTAIL.n197 VTAIL.n196 585
R64 VTAIL.n232 VTAIL.n231 585
R65 VTAIL.n230 VTAIL.n229 585
R66 VTAIL.n201 VTAIL.n200 585
R67 VTAIL.n224 VTAIL.n223 585
R68 VTAIL.n222 VTAIL.n221 585
R69 VTAIL.n205 VTAIL.n204 585
R70 VTAIL.n216 VTAIL.n215 585
R71 VTAIL.n214 VTAIL.n213 585
R72 VTAIL.n209 VTAIL.n208 585
R73 VTAIL.n175 VTAIL.n174 585
R74 VTAIL.n173 VTAIL.n172 585
R75 VTAIL.n94 VTAIL.n93 585
R76 VTAIL.n167 VTAIL.n166 585
R77 VTAIL.n165 VTAIL.n96 585
R78 VTAIL.n164 VTAIL.n163 585
R79 VTAIL.n99 VTAIL.n97 585
R80 VTAIL.n158 VTAIL.n157 585
R81 VTAIL.n156 VTAIL.n155 585
R82 VTAIL.n103 VTAIL.n102 585
R83 VTAIL.n150 VTAIL.n149 585
R84 VTAIL.n148 VTAIL.n147 585
R85 VTAIL.n107 VTAIL.n106 585
R86 VTAIL.n142 VTAIL.n141 585
R87 VTAIL.n140 VTAIL.n139 585
R88 VTAIL.n111 VTAIL.n110 585
R89 VTAIL.n134 VTAIL.n133 585
R90 VTAIL.n132 VTAIL.n131 585
R91 VTAIL.n115 VTAIL.n114 585
R92 VTAIL.n126 VTAIL.n125 585
R93 VTAIL.n124 VTAIL.n123 585
R94 VTAIL.n119 VTAIL.n118 585
R95 VTAIL.n299 VTAIL.t2 327.466
R96 VTAIL.n29 VTAIL.t0 327.466
R97 VTAIL.n210 VTAIL.t1 327.466
R98 VTAIL.n120 VTAIL.t3 327.466
R99 VTAIL.n303 VTAIL.n297 171.744
R100 VTAIL.n304 VTAIL.n303 171.744
R101 VTAIL.n304 VTAIL.n293 171.744
R102 VTAIL.n311 VTAIL.n293 171.744
R103 VTAIL.n312 VTAIL.n311 171.744
R104 VTAIL.n312 VTAIL.n289 171.744
R105 VTAIL.n319 VTAIL.n289 171.744
R106 VTAIL.n320 VTAIL.n319 171.744
R107 VTAIL.n320 VTAIL.n285 171.744
R108 VTAIL.n327 VTAIL.n285 171.744
R109 VTAIL.n328 VTAIL.n327 171.744
R110 VTAIL.n328 VTAIL.n281 171.744
R111 VTAIL.n335 VTAIL.n281 171.744
R112 VTAIL.n336 VTAIL.n335 171.744
R113 VTAIL.n336 VTAIL.n277 171.744
R114 VTAIL.n344 VTAIL.n277 171.744
R115 VTAIL.n345 VTAIL.n344 171.744
R116 VTAIL.n346 VTAIL.n345 171.744
R117 VTAIL.n346 VTAIL.n273 171.744
R118 VTAIL.n353 VTAIL.n273 171.744
R119 VTAIL.n354 VTAIL.n353 171.744
R120 VTAIL.n33 VTAIL.n27 171.744
R121 VTAIL.n34 VTAIL.n33 171.744
R122 VTAIL.n34 VTAIL.n23 171.744
R123 VTAIL.n41 VTAIL.n23 171.744
R124 VTAIL.n42 VTAIL.n41 171.744
R125 VTAIL.n42 VTAIL.n19 171.744
R126 VTAIL.n49 VTAIL.n19 171.744
R127 VTAIL.n50 VTAIL.n49 171.744
R128 VTAIL.n50 VTAIL.n15 171.744
R129 VTAIL.n57 VTAIL.n15 171.744
R130 VTAIL.n58 VTAIL.n57 171.744
R131 VTAIL.n58 VTAIL.n11 171.744
R132 VTAIL.n65 VTAIL.n11 171.744
R133 VTAIL.n66 VTAIL.n65 171.744
R134 VTAIL.n66 VTAIL.n7 171.744
R135 VTAIL.n74 VTAIL.n7 171.744
R136 VTAIL.n75 VTAIL.n74 171.744
R137 VTAIL.n76 VTAIL.n75 171.744
R138 VTAIL.n76 VTAIL.n3 171.744
R139 VTAIL.n83 VTAIL.n3 171.744
R140 VTAIL.n84 VTAIL.n83 171.744
R141 VTAIL.n264 VTAIL.n263 171.744
R142 VTAIL.n263 VTAIL.n183 171.744
R143 VTAIL.n256 VTAIL.n183 171.744
R144 VTAIL.n256 VTAIL.n255 171.744
R145 VTAIL.n255 VTAIL.n254 171.744
R146 VTAIL.n254 VTAIL.n187 171.744
R147 VTAIL.n247 VTAIL.n187 171.744
R148 VTAIL.n247 VTAIL.n246 171.744
R149 VTAIL.n246 VTAIL.n192 171.744
R150 VTAIL.n239 VTAIL.n192 171.744
R151 VTAIL.n239 VTAIL.n238 171.744
R152 VTAIL.n238 VTAIL.n196 171.744
R153 VTAIL.n231 VTAIL.n196 171.744
R154 VTAIL.n231 VTAIL.n230 171.744
R155 VTAIL.n230 VTAIL.n200 171.744
R156 VTAIL.n223 VTAIL.n200 171.744
R157 VTAIL.n223 VTAIL.n222 171.744
R158 VTAIL.n222 VTAIL.n204 171.744
R159 VTAIL.n215 VTAIL.n204 171.744
R160 VTAIL.n215 VTAIL.n214 171.744
R161 VTAIL.n214 VTAIL.n208 171.744
R162 VTAIL.n174 VTAIL.n173 171.744
R163 VTAIL.n173 VTAIL.n93 171.744
R164 VTAIL.n166 VTAIL.n93 171.744
R165 VTAIL.n166 VTAIL.n165 171.744
R166 VTAIL.n165 VTAIL.n164 171.744
R167 VTAIL.n164 VTAIL.n97 171.744
R168 VTAIL.n157 VTAIL.n97 171.744
R169 VTAIL.n157 VTAIL.n156 171.744
R170 VTAIL.n156 VTAIL.n102 171.744
R171 VTAIL.n149 VTAIL.n102 171.744
R172 VTAIL.n149 VTAIL.n148 171.744
R173 VTAIL.n148 VTAIL.n106 171.744
R174 VTAIL.n141 VTAIL.n106 171.744
R175 VTAIL.n141 VTAIL.n140 171.744
R176 VTAIL.n140 VTAIL.n110 171.744
R177 VTAIL.n133 VTAIL.n110 171.744
R178 VTAIL.n133 VTAIL.n132 171.744
R179 VTAIL.n132 VTAIL.n114 171.744
R180 VTAIL.n125 VTAIL.n114 171.744
R181 VTAIL.n125 VTAIL.n124 171.744
R182 VTAIL.n124 VTAIL.n118 171.744
R183 VTAIL.t2 VTAIL.n297 85.8723
R184 VTAIL.t0 VTAIL.n27 85.8723
R185 VTAIL.t1 VTAIL.n208 85.8723
R186 VTAIL.t3 VTAIL.n118 85.8723
R187 VTAIL.n359 VTAIL.n358 35.6763
R188 VTAIL.n89 VTAIL.n88 35.6763
R189 VTAIL.n269 VTAIL.n268 35.6763
R190 VTAIL.n179 VTAIL.n178 35.6763
R191 VTAIL.n179 VTAIL.n89 31.4186
R192 VTAIL.n359 VTAIL.n269 28.9014
R193 VTAIL.n299 VTAIL.n298 16.3895
R194 VTAIL.n29 VTAIL.n28 16.3895
R195 VTAIL.n210 VTAIL.n209 16.3895
R196 VTAIL.n120 VTAIL.n119 16.3895
R197 VTAIL.n347 VTAIL.n276 13.1884
R198 VTAIL.n77 VTAIL.n6 13.1884
R199 VTAIL.n257 VTAIL.n186 13.1884
R200 VTAIL.n167 VTAIL.n96 13.1884
R201 VTAIL.n302 VTAIL.n301 12.8005
R202 VTAIL.n343 VTAIL.n342 12.8005
R203 VTAIL.n348 VTAIL.n274 12.8005
R204 VTAIL.n32 VTAIL.n31 12.8005
R205 VTAIL.n73 VTAIL.n72 12.8005
R206 VTAIL.n78 VTAIL.n4 12.8005
R207 VTAIL.n258 VTAIL.n184 12.8005
R208 VTAIL.n253 VTAIL.n188 12.8005
R209 VTAIL.n213 VTAIL.n212 12.8005
R210 VTAIL.n168 VTAIL.n94 12.8005
R211 VTAIL.n163 VTAIL.n98 12.8005
R212 VTAIL.n123 VTAIL.n122 12.8005
R213 VTAIL.n305 VTAIL.n296 12.0247
R214 VTAIL.n341 VTAIL.n278 12.0247
R215 VTAIL.n352 VTAIL.n351 12.0247
R216 VTAIL.n35 VTAIL.n26 12.0247
R217 VTAIL.n71 VTAIL.n8 12.0247
R218 VTAIL.n82 VTAIL.n81 12.0247
R219 VTAIL.n262 VTAIL.n261 12.0247
R220 VTAIL.n252 VTAIL.n189 12.0247
R221 VTAIL.n216 VTAIL.n207 12.0247
R222 VTAIL.n172 VTAIL.n171 12.0247
R223 VTAIL.n162 VTAIL.n99 12.0247
R224 VTAIL.n126 VTAIL.n117 12.0247
R225 VTAIL.n306 VTAIL.n294 11.249
R226 VTAIL.n338 VTAIL.n337 11.249
R227 VTAIL.n355 VTAIL.n272 11.249
R228 VTAIL.n36 VTAIL.n24 11.249
R229 VTAIL.n68 VTAIL.n67 11.249
R230 VTAIL.n85 VTAIL.n2 11.249
R231 VTAIL.n265 VTAIL.n182 11.249
R232 VTAIL.n249 VTAIL.n248 11.249
R233 VTAIL.n217 VTAIL.n205 11.249
R234 VTAIL.n175 VTAIL.n92 11.249
R235 VTAIL.n159 VTAIL.n158 11.249
R236 VTAIL.n127 VTAIL.n115 11.249
R237 VTAIL.n310 VTAIL.n309 10.4732
R238 VTAIL.n334 VTAIL.n280 10.4732
R239 VTAIL.n356 VTAIL.n270 10.4732
R240 VTAIL.n40 VTAIL.n39 10.4732
R241 VTAIL.n64 VTAIL.n10 10.4732
R242 VTAIL.n86 VTAIL.n0 10.4732
R243 VTAIL.n266 VTAIL.n180 10.4732
R244 VTAIL.n245 VTAIL.n191 10.4732
R245 VTAIL.n221 VTAIL.n220 10.4732
R246 VTAIL.n176 VTAIL.n90 10.4732
R247 VTAIL.n155 VTAIL.n101 10.4732
R248 VTAIL.n131 VTAIL.n130 10.4732
R249 VTAIL.n313 VTAIL.n292 9.69747
R250 VTAIL.n333 VTAIL.n282 9.69747
R251 VTAIL.n43 VTAIL.n22 9.69747
R252 VTAIL.n63 VTAIL.n12 9.69747
R253 VTAIL.n244 VTAIL.n193 9.69747
R254 VTAIL.n224 VTAIL.n203 9.69747
R255 VTAIL.n154 VTAIL.n103 9.69747
R256 VTAIL.n134 VTAIL.n113 9.69747
R257 VTAIL.n358 VTAIL.n357 9.45567
R258 VTAIL.n88 VTAIL.n87 9.45567
R259 VTAIL.n268 VTAIL.n267 9.45567
R260 VTAIL.n178 VTAIL.n177 9.45567
R261 VTAIL.n357 VTAIL.n356 9.3005
R262 VTAIL.n272 VTAIL.n271 9.3005
R263 VTAIL.n351 VTAIL.n350 9.3005
R264 VTAIL.n349 VTAIL.n348 9.3005
R265 VTAIL.n288 VTAIL.n287 9.3005
R266 VTAIL.n317 VTAIL.n316 9.3005
R267 VTAIL.n315 VTAIL.n314 9.3005
R268 VTAIL.n292 VTAIL.n291 9.3005
R269 VTAIL.n309 VTAIL.n308 9.3005
R270 VTAIL.n307 VTAIL.n306 9.3005
R271 VTAIL.n296 VTAIL.n295 9.3005
R272 VTAIL.n301 VTAIL.n300 9.3005
R273 VTAIL.n323 VTAIL.n322 9.3005
R274 VTAIL.n325 VTAIL.n324 9.3005
R275 VTAIL.n284 VTAIL.n283 9.3005
R276 VTAIL.n331 VTAIL.n330 9.3005
R277 VTAIL.n333 VTAIL.n332 9.3005
R278 VTAIL.n280 VTAIL.n279 9.3005
R279 VTAIL.n339 VTAIL.n338 9.3005
R280 VTAIL.n341 VTAIL.n340 9.3005
R281 VTAIL.n342 VTAIL.n275 9.3005
R282 VTAIL.n87 VTAIL.n86 9.3005
R283 VTAIL.n2 VTAIL.n1 9.3005
R284 VTAIL.n81 VTAIL.n80 9.3005
R285 VTAIL.n79 VTAIL.n78 9.3005
R286 VTAIL.n18 VTAIL.n17 9.3005
R287 VTAIL.n47 VTAIL.n46 9.3005
R288 VTAIL.n45 VTAIL.n44 9.3005
R289 VTAIL.n22 VTAIL.n21 9.3005
R290 VTAIL.n39 VTAIL.n38 9.3005
R291 VTAIL.n37 VTAIL.n36 9.3005
R292 VTAIL.n26 VTAIL.n25 9.3005
R293 VTAIL.n31 VTAIL.n30 9.3005
R294 VTAIL.n53 VTAIL.n52 9.3005
R295 VTAIL.n55 VTAIL.n54 9.3005
R296 VTAIL.n14 VTAIL.n13 9.3005
R297 VTAIL.n61 VTAIL.n60 9.3005
R298 VTAIL.n63 VTAIL.n62 9.3005
R299 VTAIL.n10 VTAIL.n9 9.3005
R300 VTAIL.n69 VTAIL.n68 9.3005
R301 VTAIL.n71 VTAIL.n70 9.3005
R302 VTAIL.n72 VTAIL.n5 9.3005
R303 VTAIL.n236 VTAIL.n235 9.3005
R304 VTAIL.n195 VTAIL.n194 9.3005
R305 VTAIL.n242 VTAIL.n241 9.3005
R306 VTAIL.n244 VTAIL.n243 9.3005
R307 VTAIL.n191 VTAIL.n190 9.3005
R308 VTAIL.n250 VTAIL.n249 9.3005
R309 VTAIL.n252 VTAIL.n251 9.3005
R310 VTAIL.n188 VTAIL.n185 9.3005
R311 VTAIL.n267 VTAIL.n266 9.3005
R312 VTAIL.n182 VTAIL.n181 9.3005
R313 VTAIL.n261 VTAIL.n260 9.3005
R314 VTAIL.n259 VTAIL.n258 9.3005
R315 VTAIL.n234 VTAIL.n233 9.3005
R316 VTAIL.n199 VTAIL.n198 9.3005
R317 VTAIL.n228 VTAIL.n227 9.3005
R318 VTAIL.n226 VTAIL.n225 9.3005
R319 VTAIL.n203 VTAIL.n202 9.3005
R320 VTAIL.n220 VTAIL.n219 9.3005
R321 VTAIL.n218 VTAIL.n217 9.3005
R322 VTAIL.n207 VTAIL.n206 9.3005
R323 VTAIL.n212 VTAIL.n211 9.3005
R324 VTAIL.n146 VTAIL.n145 9.3005
R325 VTAIL.n105 VTAIL.n104 9.3005
R326 VTAIL.n152 VTAIL.n151 9.3005
R327 VTAIL.n154 VTAIL.n153 9.3005
R328 VTAIL.n101 VTAIL.n100 9.3005
R329 VTAIL.n160 VTAIL.n159 9.3005
R330 VTAIL.n162 VTAIL.n161 9.3005
R331 VTAIL.n98 VTAIL.n95 9.3005
R332 VTAIL.n177 VTAIL.n176 9.3005
R333 VTAIL.n92 VTAIL.n91 9.3005
R334 VTAIL.n171 VTAIL.n170 9.3005
R335 VTAIL.n169 VTAIL.n168 9.3005
R336 VTAIL.n144 VTAIL.n143 9.3005
R337 VTAIL.n109 VTAIL.n108 9.3005
R338 VTAIL.n138 VTAIL.n137 9.3005
R339 VTAIL.n136 VTAIL.n135 9.3005
R340 VTAIL.n113 VTAIL.n112 9.3005
R341 VTAIL.n130 VTAIL.n129 9.3005
R342 VTAIL.n128 VTAIL.n127 9.3005
R343 VTAIL.n117 VTAIL.n116 9.3005
R344 VTAIL.n122 VTAIL.n121 9.3005
R345 VTAIL.n314 VTAIL.n290 8.92171
R346 VTAIL.n330 VTAIL.n329 8.92171
R347 VTAIL.n44 VTAIL.n20 8.92171
R348 VTAIL.n60 VTAIL.n59 8.92171
R349 VTAIL.n241 VTAIL.n240 8.92171
R350 VTAIL.n225 VTAIL.n201 8.92171
R351 VTAIL.n151 VTAIL.n150 8.92171
R352 VTAIL.n135 VTAIL.n111 8.92171
R353 VTAIL.n318 VTAIL.n317 8.14595
R354 VTAIL.n326 VTAIL.n284 8.14595
R355 VTAIL.n48 VTAIL.n47 8.14595
R356 VTAIL.n56 VTAIL.n14 8.14595
R357 VTAIL.n237 VTAIL.n195 8.14595
R358 VTAIL.n229 VTAIL.n228 8.14595
R359 VTAIL.n147 VTAIL.n105 8.14595
R360 VTAIL.n139 VTAIL.n138 8.14595
R361 VTAIL.n321 VTAIL.n288 7.3702
R362 VTAIL.n325 VTAIL.n286 7.3702
R363 VTAIL.n51 VTAIL.n18 7.3702
R364 VTAIL.n55 VTAIL.n16 7.3702
R365 VTAIL.n236 VTAIL.n197 7.3702
R366 VTAIL.n232 VTAIL.n199 7.3702
R367 VTAIL.n146 VTAIL.n107 7.3702
R368 VTAIL.n142 VTAIL.n109 7.3702
R369 VTAIL.n322 VTAIL.n321 6.59444
R370 VTAIL.n322 VTAIL.n286 6.59444
R371 VTAIL.n52 VTAIL.n51 6.59444
R372 VTAIL.n52 VTAIL.n16 6.59444
R373 VTAIL.n233 VTAIL.n197 6.59444
R374 VTAIL.n233 VTAIL.n232 6.59444
R375 VTAIL.n143 VTAIL.n107 6.59444
R376 VTAIL.n143 VTAIL.n142 6.59444
R377 VTAIL.n318 VTAIL.n288 5.81868
R378 VTAIL.n326 VTAIL.n325 5.81868
R379 VTAIL.n48 VTAIL.n18 5.81868
R380 VTAIL.n56 VTAIL.n55 5.81868
R381 VTAIL.n237 VTAIL.n236 5.81868
R382 VTAIL.n229 VTAIL.n199 5.81868
R383 VTAIL.n147 VTAIL.n146 5.81868
R384 VTAIL.n139 VTAIL.n109 5.81868
R385 VTAIL.n317 VTAIL.n290 5.04292
R386 VTAIL.n329 VTAIL.n284 5.04292
R387 VTAIL.n47 VTAIL.n20 5.04292
R388 VTAIL.n59 VTAIL.n14 5.04292
R389 VTAIL.n240 VTAIL.n195 5.04292
R390 VTAIL.n228 VTAIL.n201 5.04292
R391 VTAIL.n150 VTAIL.n105 5.04292
R392 VTAIL.n138 VTAIL.n111 5.04292
R393 VTAIL.n314 VTAIL.n313 4.26717
R394 VTAIL.n330 VTAIL.n282 4.26717
R395 VTAIL.n44 VTAIL.n43 4.26717
R396 VTAIL.n60 VTAIL.n12 4.26717
R397 VTAIL.n241 VTAIL.n193 4.26717
R398 VTAIL.n225 VTAIL.n224 4.26717
R399 VTAIL.n151 VTAIL.n103 4.26717
R400 VTAIL.n135 VTAIL.n134 4.26717
R401 VTAIL.n300 VTAIL.n299 3.70982
R402 VTAIL.n30 VTAIL.n29 3.70982
R403 VTAIL.n211 VTAIL.n210 3.70982
R404 VTAIL.n121 VTAIL.n120 3.70982
R405 VTAIL.n310 VTAIL.n292 3.49141
R406 VTAIL.n334 VTAIL.n333 3.49141
R407 VTAIL.n358 VTAIL.n270 3.49141
R408 VTAIL.n40 VTAIL.n22 3.49141
R409 VTAIL.n64 VTAIL.n63 3.49141
R410 VTAIL.n88 VTAIL.n0 3.49141
R411 VTAIL.n268 VTAIL.n180 3.49141
R412 VTAIL.n245 VTAIL.n244 3.49141
R413 VTAIL.n221 VTAIL.n203 3.49141
R414 VTAIL.n178 VTAIL.n90 3.49141
R415 VTAIL.n155 VTAIL.n154 3.49141
R416 VTAIL.n131 VTAIL.n113 3.49141
R417 VTAIL.n309 VTAIL.n294 2.71565
R418 VTAIL.n337 VTAIL.n280 2.71565
R419 VTAIL.n356 VTAIL.n355 2.71565
R420 VTAIL.n39 VTAIL.n24 2.71565
R421 VTAIL.n67 VTAIL.n10 2.71565
R422 VTAIL.n86 VTAIL.n85 2.71565
R423 VTAIL.n266 VTAIL.n265 2.71565
R424 VTAIL.n248 VTAIL.n191 2.71565
R425 VTAIL.n220 VTAIL.n205 2.71565
R426 VTAIL.n176 VTAIL.n175 2.71565
R427 VTAIL.n158 VTAIL.n101 2.71565
R428 VTAIL.n130 VTAIL.n115 2.71565
R429 VTAIL.n306 VTAIL.n305 1.93989
R430 VTAIL.n338 VTAIL.n278 1.93989
R431 VTAIL.n352 VTAIL.n272 1.93989
R432 VTAIL.n36 VTAIL.n35 1.93989
R433 VTAIL.n68 VTAIL.n8 1.93989
R434 VTAIL.n82 VTAIL.n2 1.93989
R435 VTAIL.n262 VTAIL.n182 1.93989
R436 VTAIL.n249 VTAIL.n189 1.93989
R437 VTAIL.n217 VTAIL.n216 1.93989
R438 VTAIL.n172 VTAIL.n92 1.93989
R439 VTAIL.n159 VTAIL.n99 1.93989
R440 VTAIL.n127 VTAIL.n126 1.93989
R441 VTAIL.n269 VTAIL.n179 1.72895
R442 VTAIL.n302 VTAIL.n296 1.16414
R443 VTAIL.n343 VTAIL.n341 1.16414
R444 VTAIL.n351 VTAIL.n274 1.16414
R445 VTAIL.n32 VTAIL.n26 1.16414
R446 VTAIL.n73 VTAIL.n71 1.16414
R447 VTAIL.n81 VTAIL.n4 1.16414
R448 VTAIL.n261 VTAIL.n184 1.16414
R449 VTAIL.n253 VTAIL.n252 1.16414
R450 VTAIL.n213 VTAIL.n207 1.16414
R451 VTAIL.n171 VTAIL.n94 1.16414
R452 VTAIL.n163 VTAIL.n162 1.16414
R453 VTAIL.n123 VTAIL.n117 1.16414
R454 VTAIL VTAIL.n89 1.15783
R455 VTAIL VTAIL.n359 0.571621
R456 VTAIL.n301 VTAIL.n298 0.388379
R457 VTAIL.n342 VTAIL.n276 0.388379
R458 VTAIL.n348 VTAIL.n347 0.388379
R459 VTAIL.n31 VTAIL.n28 0.388379
R460 VTAIL.n72 VTAIL.n6 0.388379
R461 VTAIL.n78 VTAIL.n77 0.388379
R462 VTAIL.n258 VTAIL.n257 0.388379
R463 VTAIL.n188 VTAIL.n186 0.388379
R464 VTAIL.n212 VTAIL.n209 0.388379
R465 VTAIL.n168 VTAIL.n167 0.388379
R466 VTAIL.n98 VTAIL.n96 0.388379
R467 VTAIL.n122 VTAIL.n119 0.388379
R468 VTAIL.n300 VTAIL.n295 0.155672
R469 VTAIL.n307 VTAIL.n295 0.155672
R470 VTAIL.n308 VTAIL.n307 0.155672
R471 VTAIL.n308 VTAIL.n291 0.155672
R472 VTAIL.n315 VTAIL.n291 0.155672
R473 VTAIL.n316 VTAIL.n315 0.155672
R474 VTAIL.n316 VTAIL.n287 0.155672
R475 VTAIL.n323 VTAIL.n287 0.155672
R476 VTAIL.n324 VTAIL.n323 0.155672
R477 VTAIL.n324 VTAIL.n283 0.155672
R478 VTAIL.n331 VTAIL.n283 0.155672
R479 VTAIL.n332 VTAIL.n331 0.155672
R480 VTAIL.n332 VTAIL.n279 0.155672
R481 VTAIL.n339 VTAIL.n279 0.155672
R482 VTAIL.n340 VTAIL.n339 0.155672
R483 VTAIL.n340 VTAIL.n275 0.155672
R484 VTAIL.n349 VTAIL.n275 0.155672
R485 VTAIL.n350 VTAIL.n349 0.155672
R486 VTAIL.n350 VTAIL.n271 0.155672
R487 VTAIL.n357 VTAIL.n271 0.155672
R488 VTAIL.n30 VTAIL.n25 0.155672
R489 VTAIL.n37 VTAIL.n25 0.155672
R490 VTAIL.n38 VTAIL.n37 0.155672
R491 VTAIL.n38 VTAIL.n21 0.155672
R492 VTAIL.n45 VTAIL.n21 0.155672
R493 VTAIL.n46 VTAIL.n45 0.155672
R494 VTAIL.n46 VTAIL.n17 0.155672
R495 VTAIL.n53 VTAIL.n17 0.155672
R496 VTAIL.n54 VTAIL.n53 0.155672
R497 VTAIL.n54 VTAIL.n13 0.155672
R498 VTAIL.n61 VTAIL.n13 0.155672
R499 VTAIL.n62 VTAIL.n61 0.155672
R500 VTAIL.n62 VTAIL.n9 0.155672
R501 VTAIL.n69 VTAIL.n9 0.155672
R502 VTAIL.n70 VTAIL.n69 0.155672
R503 VTAIL.n70 VTAIL.n5 0.155672
R504 VTAIL.n79 VTAIL.n5 0.155672
R505 VTAIL.n80 VTAIL.n79 0.155672
R506 VTAIL.n80 VTAIL.n1 0.155672
R507 VTAIL.n87 VTAIL.n1 0.155672
R508 VTAIL.n267 VTAIL.n181 0.155672
R509 VTAIL.n260 VTAIL.n181 0.155672
R510 VTAIL.n260 VTAIL.n259 0.155672
R511 VTAIL.n259 VTAIL.n185 0.155672
R512 VTAIL.n251 VTAIL.n185 0.155672
R513 VTAIL.n251 VTAIL.n250 0.155672
R514 VTAIL.n250 VTAIL.n190 0.155672
R515 VTAIL.n243 VTAIL.n190 0.155672
R516 VTAIL.n243 VTAIL.n242 0.155672
R517 VTAIL.n242 VTAIL.n194 0.155672
R518 VTAIL.n235 VTAIL.n194 0.155672
R519 VTAIL.n235 VTAIL.n234 0.155672
R520 VTAIL.n234 VTAIL.n198 0.155672
R521 VTAIL.n227 VTAIL.n198 0.155672
R522 VTAIL.n227 VTAIL.n226 0.155672
R523 VTAIL.n226 VTAIL.n202 0.155672
R524 VTAIL.n219 VTAIL.n202 0.155672
R525 VTAIL.n219 VTAIL.n218 0.155672
R526 VTAIL.n218 VTAIL.n206 0.155672
R527 VTAIL.n211 VTAIL.n206 0.155672
R528 VTAIL.n177 VTAIL.n91 0.155672
R529 VTAIL.n170 VTAIL.n91 0.155672
R530 VTAIL.n170 VTAIL.n169 0.155672
R531 VTAIL.n169 VTAIL.n95 0.155672
R532 VTAIL.n161 VTAIL.n95 0.155672
R533 VTAIL.n161 VTAIL.n160 0.155672
R534 VTAIL.n160 VTAIL.n100 0.155672
R535 VTAIL.n153 VTAIL.n100 0.155672
R536 VTAIL.n153 VTAIL.n152 0.155672
R537 VTAIL.n152 VTAIL.n104 0.155672
R538 VTAIL.n145 VTAIL.n104 0.155672
R539 VTAIL.n145 VTAIL.n144 0.155672
R540 VTAIL.n144 VTAIL.n108 0.155672
R541 VTAIL.n137 VTAIL.n108 0.155672
R542 VTAIL.n137 VTAIL.n136 0.155672
R543 VTAIL.n136 VTAIL.n112 0.155672
R544 VTAIL.n129 VTAIL.n112 0.155672
R545 VTAIL.n129 VTAIL.n128 0.155672
R546 VTAIL.n128 VTAIL.n116 0.155672
R547 VTAIL.n121 VTAIL.n116 0.155672
R548 VDD1.n84 VDD1.n0 756.745
R549 VDD1.n173 VDD1.n89 756.745
R550 VDD1.n85 VDD1.n84 585
R551 VDD1.n83 VDD1.n82 585
R552 VDD1.n4 VDD1.n3 585
R553 VDD1.n77 VDD1.n76 585
R554 VDD1.n75 VDD1.n6 585
R555 VDD1.n74 VDD1.n73 585
R556 VDD1.n9 VDD1.n7 585
R557 VDD1.n68 VDD1.n67 585
R558 VDD1.n66 VDD1.n65 585
R559 VDD1.n13 VDD1.n12 585
R560 VDD1.n60 VDD1.n59 585
R561 VDD1.n58 VDD1.n57 585
R562 VDD1.n17 VDD1.n16 585
R563 VDD1.n52 VDD1.n51 585
R564 VDD1.n50 VDD1.n49 585
R565 VDD1.n21 VDD1.n20 585
R566 VDD1.n44 VDD1.n43 585
R567 VDD1.n42 VDD1.n41 585
R568 VDD1.n25 VDD1.n24 585
R569 VDD1.n36 VDD1.n35 585
R570 VDD1.n34 VDD1.n33 585
R571 VDD1.n29 VDD1.n28 585
R572 VDD1.n117 VDD1.n116 585
R573 VDD1.n122 VDD1.n121 585
R574 VDD1.n124 VDD1.n123 585
R575 VDD1.n113 VDD1.n112 585
R576 VDD1.n130 VDD1.n129 585
R577 VDD1.n132 VDD1.n131 585
R578 VDD1.n109 VDD1.n108 585
R579 VDD1.n138 VDD1.n137 585
R580 VDD1.n140 VDD1.n139 585
R581 VDD1.n105 VDD1.n104 585
R582 VDD1.n146 VDD1.n145 585
R583 VDD1.n148 VDD1.n147 585
R584 VDD1.n101 VDD1.n100 585
R585 VDD1.n154 VDD1.n153 585
R586 VDD1.n156 VDD1.n155 585
R587 VDD1.n97 VDD1.n96 585
R588 VDD1.n163 VDD1.n162 585
R589 VDD1.n164 VDD1.n95 585
R590 VDD1.n166 VDD1.n165 585
R591 VDD1.n93 VDD1.n92 585
R592 VDD1.n172 VDD1.n171 585
R593 VDD1.n174 VDD1.n173 585
R594 VDD1.n30 VDD1.t0 327.466
R595 VDD1.n118 VDD1.t1 327.466
R596 VDD1.n84 VDD1.n83 171.744
R597 VDD1.n83 VDD1.n3 171.744
R598 VDD1.n76 VDD1.n3 171.744
R599 VDD1.n76 VDD1.n75 171.744
R600 VDD1.n75 VDD1.n74 171.744
R601 VDD1.n74 VDD1.n7 171.744
R602 VDD1.n67 VDD1.n7 171.744
R603 VDD1.n67 VDD1.n66 171.744
R604 VDD1.n66 VDD1.n12 171.744
R605 VDD1.n59 VDD1.n12 171.744
R606 VDD1.n59 VDD1.n58 171.744
R607 VDD1.n58 VDD1.n16 171.744
R608 VDD1.n51 VDD1.n16 171.744
R609 VDD1.n51 VDD1.n50 171.744
R610 VDD1.n50 VDD1.n20 171.744
R611 VDD1.n43 VDD1.n20 171.744
R612 VDD1.n43 VDD1.n42 171.744
R613 VDD1.n42 VDD1.n24 171.744
R614 VDD1.n35 VDD1.n24 171.744
R615 VDD1.n35 VDD1.n34 171.744
R616 VDD1.n34 VDD1.n28 171.744
R617 VDD1.n122 VDD1.n116 171.744
R618 VDD1.n123 VDD1.n122 171.744
R619 VDD1.n123 VDD1.n112 171.744
R620 VDD1.n130 VDD1.n112 171.744
R621 VDD1.n131 VDD1.n130 171.744
R622 VDD1.n131 VDD1.n108 171.744
R623 VDD1.n138 VDD1.n108 171.744
R624 VDD1.n139 VDD1.n138 171.744
R625 VDD1.n139 VDD1.n104 171.744
R626 VDD1.n146 VDD1.n104 171.744
R627 VDD1.n147 VDD1.n146 171.744
R628 VDD1.n147 VDD1.n100 171.744
R629 VDD1.n154 VDD1.n100 171.744
R630 VDD1.n155 VDD1.n154 171.744
R631 VDD1.n155 VDD1.n96 171.744
R632 VDD1.n163 VDD1.n96 171.744
R633 VDD1.n164 VDD1.n163 171.744
R634 VDD1.n165 VDD1.n164 171.744
R635 VDD1.n165 VDD1.n92 171.744
R636 VDD1.n172 VDD1.n92 171.744
R637 VDD1.n173 VDD1.n172 171.744
R638 VDD1 VDD1.n177 96.2203
R639 VDD1.t0 VDD1.n28 85.8723
R640 VDD1.t1 VDD1.n116 85.8723
R641 VDD1 VDD1.n88 53.0425
R642 VDD1.n30 VDD1.n29 16.3895
R643 VDD1.n118 VDD1.n117 16.3895
R644 VDD1.n77 VDD1.n6 13.1884
R645 VDD1.n166 VDD1.n95 13.1884
R646 VDD1.n78 VDD1.n4 12.8005
R647 VDD1.n73 VDD1.n8 12.8005
R648 VDD1.n33 VDD1.n32 12.8005
R649 VDD1.n121 VDD1.n120 12.8005
R650 VDD1.n162 VDD1.n161 12.8005
R651 VDD1.n167 VDD1.n93 12.8005
R652 VDD1.n82 VDD1.n81 12.0247
R653 VDD1.n72 VDD1.n9 12.0247
R654 VDD1.n36 VDD1.n27 12.0247
R655 VDD1.n124 VDD1.n115 12.0247
R656 VDD1.n160 VDD1.n97 12.0247
R657 VDD1.n171 VDD1.n170 12.0247
R658 VDD1.n85 VDD1.n2 11.249
R659 VDD1.n69 VDD1.n68 11.249
R660 VDD1.n37 VDD1.n25 11.249
R661 VDD1.n125 VDD1.n113 11.249
R662 VDD1.n157 VDD1.n156 11.249
R663 VDD1.n174 VDD1.n91 11.249
R664 VDD1.n86 VDD1.n0 10.4732
R665 VDD1.n65 VDD1.n11 10.4732
R666 VDD1.n41 VDD1.n40 10.4732
R667 VDD1.n129 VDD1.n128 10.4732
R668 VDD1.n153 VDD1.n99 10.4732
R669 VDD1.n175 VDD1.n89 10.4732
R670 VDD1.n64 VDD1.n13 9.69747
R671 VDD1.n44 VDD1.n23 9.69747
R672 VDD1.n132 VDD1.n111 9.69747
R673 VDD1.n152 VDD1.n101 9.69747
R674 VDD1.n88 VDD1.n87 9.45567
R675 VDD1.n177 VDD1.n176 9.45567
R676 VDD1.n56 VDD1.n55 9.3005
R677 VDD1.n15 VDD1.n14 9.3005
R678 VDD1.n62 VDD1.n61 9.3005
R679 VDD1.n64 VDD1.n63 9.3005
R680 VDD1.n11 VDD1.n10 9.3005
R681 VDD1.n70 VDD1.n69 9.3005
R682 VDD1.n72 VDD1.n71 9.3005
R683 VDD1.n8 VDD1.n5 9.3005
R684 VDD1.n87 VDD1.n86 9.3005
R685 VDD1.n2 VDD1.n1 9.3005
R686 VDD1.n81 VDD1.n80 9.3005
R687 VDD1.n79 VDD1.n78 9.3005
R688 VDD1.n54 VDD1.n53 9.3005
R689 VDD1.n19 VDD1.n18 9.3005
R690 VDD1.n48 VDD1.n47 9.3005
R691 VDD1.n46 VDD1.n45 9.3005
R692 VDD1.n23 VDD1.n22 9.3005
R693 VDD1.n40 VDD1.n39 9.3005
R694 VDD1.n38 VDD1.n37 9.3005
R695 VDD1.n27 VDD1.n26 9.3005
R696 VDD1.n32 VDD1.n31 9.3005
R697 VDD1.n176 VDD1.n175 9.3005
R698 VDD1.n91 VDD1.n90 9.3005
R699 VDD1.n170 VDD1.n169 9.3005
R700 VDD1.n168 VDD1.n167 9.3005
R701 VDD1.n107 VDD1.n106 9.3005
R702 VDD1.n136 VDD1.n135 9.3005
R703 VDD1.n134 VDD1.n133 9.3005
R704 VDD1.n111 VDD1.n110 9.3005
R705 VDD1.n128 VDD1.n127 9.3005
R706 VDD1.n126 VDD1.n125 9.3005
R707 VDD1.n115 VDD1.n114 9.3005
R708 VDD1.n120 VDD1.n119 9.3005
R709 VDD1.n142 VDD1.n141 9.3005
R710 VDD1.n144 VDD1.n143 9.3005
R711 VDD1.n103 VDD1.n102 9.3005
R712 VDD1.n150 VDD1.n149 9.3005
R713 VDD1.n152 VDD1.n151 9.3005
R714 VDD1.n99 VDD1.n98 9.3005
R715 VDD1.n158 VDD1.n157 9.3005
R716 VDD1.n160 VDD1.n159 9.3005
R717 VDD1.n161 VDD1.n94 9.3005
R718 VDD1.n61 VDD1.n60 8.92171
R719 VDD1.n45 VDD1.n21 8.92171
R720 VDD1.n133 VDD1.n109 8.92171
R721 VDD1.n149 VDD1.n148 8.92171
R722 VDD1.n57 VDD1.n15 8.14595
R723 VDD1.n49 VDD1.n48 8.14595
R724 VDD1.n137 VDD1.n136 8.14595
R725 VDD1.n145 VDD1.n103 8.14595
R726 VDD1.n56 VDD1.n17 7.3702
R727 VDD1.n52 VDD1.n19 7.3702
R728 VDD1.n140 VDD1.n107 7.3702
R729 VDD1.n144 VDD1.n105 7.3702
R730 VDD1.n53 VDD1.n17 6.59444
R731 VDD1.n53 VDD1.n52 6.59444
R732 VDD1.n141 VDD1.n140 6.59444
R733 VDD1.n141 VDD1.n105 6.59444
R734 VDD1.n57 VDD1.n56 5.81868
R735 VDD1.n49 VDD1.n19 5.81868
R736 VDD1.n137 VDD1.n107 5.81868
R737 VDD1.n145 VDD1.n144 5.81868
R738 VDD1.n60 VDD1.n15 5.04292
R739 VDD1.n48 VDD1.n21 5.04292
R740 VDD1.n136 VDD1.n109 5.04292
R741 VDD1.n148 VDD1.n103 5.04292
R742 VDD1.n61 VDD1.n13 4.26717
R743 VDD1.n45 VDD1.n44 4.26717
R744 VDD1.n133 VDD1.n132 4.26717
R745 VDD1.n149 VDD1.n101 4.26717
R746 VDD1.n31 VDD1.n30 3.70982
R747 VDD1.n119 VDD1.n118 3.70982
R748 VDD1.n88 VDD1.n0 3.49141
R749 VDD1.n65 VDD1.n64 3.49141
R750 VDD1.n41 VDD1.n23 3.49141
R751 VDD1.n129 VDD1.n111 3.49141
R752 VDD1.n153 VDD1.n152 3.49141
R753 VDD1.n177 VDD1.n89 3.49141
R754 VDD1.n86 VDD1.n85 2.71565
R755 VDD1.n68 VDD1.n11 2.71565
R756 VDD1.n40 VDD1.n25 2.71565
R757 VDD1.n128 VDD1.n113 2.71565
R758 VDD1.n156 VDD1.n99 2.71565
R759 VDD1.n175 VDD1.n174 2.71565
R760 VDD1.n82 VDD1.n2 1.93989
R761 VDD1.n69 VDD1.n9 1.93989
R762 VDD1.n37 VDD1.n36 1.93989
R763 VDD1.n125 VDD1.n124 1.93989
R764 VDD1.n157 VDD1.n97 1.93989
R765 VDD1.n171 VDD1.n91 1.93989
R766 VDD1.n81 VDD1.n4 1.16414
R767 VDD1.n73 VDD1.n72 1.16414
R768 VDD1.n33 VDD1.n27 1.16414
R769 VDD1.n121 VDD1.n115 1.16414
R770 VDD1.n162 VDD1.n160 1.16414
R771 VDD1.n170 VDD1.n93 1.16414
R772 VDD1.n78 VDD1.n77 0.388379
R773 VDD1.n8 VDD1.n6 0.388379
R774 VDD1.n32 VDD1.n29 0.388379
R775 VDD1.n120 VDD1.n117 0.388379
R776 VDD1.n161 VDD1.n95 0.388379
R777 VDD1.n167 VDD1.n166 0.388379
R778 VDD1.n87 VDD1.n1 0.155672
R779 VDD1.n80 VDD1.n1 0.155672
R780 VDD1.n80 VDD1.n79 0.155672
R781 VDD1.n79 VDD1.n5 0.155672
R782 VDD1.n71 VDD1.n5 0.155672
R783 VDD1.n71 VDD1.n70 0.155672
R784 VDD1.n70 VDD1.n10 0.155672
R785 VDD1.n63 VDD1.n10 0.155672
R786 VDD1.n63 VDD1.n62 0.155672
R787 VDD1.n62 VDD1.n14 0.155672
R788 VDD1.n55 VDD1.n14 0.155672
R789 VDD1.n55 VDD1.n54 0.155672
R790 VDD1.n54 VDD1.n18 0.155672
R791 VDD1.n47 VDD1.n18 0.155672
R792 VDD1.n47 VDD1.n46 0.155672
R793 VDD1.n46 VDD1.n22 0.155672
R794 VDD1.n39 VDD1.n22 0.155672
R795 VDD1.n39 VDD1.n38 0.155672
R796 VDD1.n38 VDD1.n26 0.155672
R797 VDD1.n31 VDD1.n26 0.155672
R798 VDD1.n119 VDD1.n114 0.155672
R799 VDD1.n126 VDD1.n114 0.155672
R800 VDD1.n127 VDD1.n126 0.155672
R801 VDD1.n127 VDD1.n110 0.155672
R802 VDD1.n134 VDD1.n110 0.155672
R803 VDD1.n135 VDD1.n134 0.155672
R804 VDD1.n135 VDD1.n106 0.155672
R805 VDD1.n142 VDD1.n106 0.155672
R806 VDD1.n143 VDD1.n142 0.155672
R807 VDD1.n143 VDD1.n102 0.155672
R808 VDD1.n150 VDD1.n102 0.155672
R809 VDD1.n151 VDD1.n150 0.155672
R810 VDD1.n151 VDD1.n98 0.155672
R811 VDD1.n158 VDD1.n98 0.155672
R812 VDD1.n159 VDD1.n158 0.155672
R813 VDD1.n159 VDD1.n94 0.155672
R814 VDD1.n168 VDD1.n94 0.155672
R815 VDD1.n169 VDD1.n168 0.155672
R816 VDD1.n169 VDD1.n90 0.155672
R817 VDD1.n176 VDD1.n90 0.155672
R818 VN VN.t1 248.38
R819 VN VN.t0 200.762
R820 VDD2.n173 VDD2.n89 756.745
R821 VDD2.n84 VDD2.n0 756.745
R822 VDD2.n174 VDD2.n173 585
R823 VDD2.n172 VDD2.n171 585
R824 VDD2.n93 VDD2.n92 585
R825 VDD2.n166 VDD2.n165 585
R826 VDD2.n164 VDD2.n95 585
R827 VDD2.n163 VDD2.n162 585
R828 VDD2.n98 VDD2.n96 585
R829 VDD2.n157 VDD2.n156 585
R830 VDD2.n155 VDD2.n154 585
R831 VDD2.n102 VDD2.n101 585
R832 VDD2.n149 VDD2.n148 585
R833 VDD2.n147 VDD2.n146 585
R834 VDD2.n106 VDD2.n105 585
R835 VDD2.n141 VDD2.n140 585
R836 VDD2.n139 VDD2.n138 585
R837 VDD2.n110 VDD2.n109 585
R838 VDD2.n133 VDD2.n132 585
R839 VDD2.n131 VDD2.n130 585
R840 VDD2.n114 VDD2.n113 585
R841 VDD2.n125 VDD2.n124 585
R842 VDD2.n123 VDD2.n122 585
R843 VDD2.n118 VDD2.n117 585
R844 VDD2.n28 VDD2.n27 585
R845 VDD2.n33 VDD2.n32 585
R846 VDD2.n35 VDD2.n34 585
R847 VDD2.n24 VDD2.n23 585
R848 VDD2.n41 VDD2.n40 585
R849 VDD2.n43 VDD2.n42 585
R850 VDD2.n20 VDD2.n19 585
R851 VDD2.n49 VDD2.n48 585
R852 VDD2.n51 VDD2.n50 585
R853 VDD2.n16 VDD2.n15 585
R854 VDD2.n57 VDD2.n56 585
R855 VDD2.n59 VDD2.n58 585
R856 VDD2.n12 VDD2.n11 585
R857 VDD2.n65 VDD2.n64 585
R858 VDD2.n67 VDD2.n66 585
R859 VDD2.n8 VDD2.n7 585
R860 VDD2.n74 VDD2.n73 585
R861 VDD2.n75 VDD2.n6 585
R862 VDD2.n77 VDD2.n76 585
R863 VDD2.n4 VDD2.n3 585
R864 VDD2.n83 VDD2.n82 585
R865 VDD2.n85 VDD2.n84 585
R866 VDD2.n119 VDD2.t0 327.466
R867 VDD2.n29 VDD2.t1 327.466
R868 VDD2.n173 VDD2.n172 171.744
R869 VDD2.n172 VDD2.n92 171.744
R870 VDD2.n165 VDD2.n92 171.744
R871 VDD2.n165 VDD2.n164 171.744
R872 VDD2.n164 VDD2.n163 171.744
R873 VDD2.n163 VDD2.n96 171.744
R874 VDD2.n156 VDD2.n96 171.744
R875 VDD2.n156 VDD2.n155 171.744
R876 VDD2.n155 VDD2.n101 171.744
R877 VDD2.n148 VDD2.n101 171.744
R878 VDD2.n148 VDD2.n147 171.744
R879 VDD2.n147 VDD2.n105 171.744
R880 VDD2.n140 VDD2.n105 171.744
R881 VDD2.n140 VDD2.n139 171.744
R882 VDD2.n139 VDD2.n109 171.744
R883 VDD2.n132 VDD2.n109 171.744
R884 VDD2.n132 VDD2.n131 171.744
R885 VDD2.n131 VDD2.n113 171.744
R886 VDD2.n124 VDD2.n113 171.744
R887 VDD2.n124 VDD2.n123 171.744
R888 VDD2.n123 VDD2.n117 171.744
R889 VDD2.n33 VDD2.n27 171.744
R890 VDD2.n34 VDD2.n33 171.744
R891 VDD2.n34 VDD2.n23 171.744
R892 VDD2.n41 VDD2.n23 171.744
R893 VDD2.n42 VDD2.n41 171.744
R894 VDD2.n42 VDD2.n19 171.744
R895 VDD2.n49 VDD2.n19 171.744
R896 VDD2.n50 VDD2.n49 171.744
R897 VDD2.n50 VDD2.n15 171.744
R898 VDD2.n57 VDD2.n15 171.744
R899 VDD2.n58 VDD2.n57 171.744
R900 VDD2.n58 VDD2.n11 171.744
R901 VDD2.n65 VDD2.n11 171.744
R902 VDD2.n66 VDD2.n65 171.744
R903 VDD2.n66 VDD2.n7 171.744
R904 VDD2.n74 VDD2.n7 171.744
R905 VDD2.n75 VDD2.n74 171.744
R906 VDD2.n76 VDD2.n75 171.744
R907 VDD2.n76 VDD2.n3 171.744
R908 VDD2.n83 VDD2.n3 171.744
R909 VDD2.n84 VDD2.n83 171.744
R910 VDD2.n178 VDD2.n88 95.0662
R911 VDD2.t0 VDD2.n117 85.8723
R912 VDD2.t1 VDD2.n27 85.8723
R913 VDD2.n178 VDD2.n177 52.355
R914 VDD2.n119 VDD2.n118 16.3895
R915 VDD2.n29 VDD2.n28 16.3895
R916 VDD2.n166 VDD2.n95 13.1884
R917 VDD2.n77 VDD2.n6 13.1884
R918 VDD2.n167 VDD2.n93 12.8005
R919 VDD2.n162 VDD2.n97 12.8005
R920 VDD2.n122 VDD2.n121 12.8005
R921 VDD2.n32 VDD2.n31 12.8005
R922 VDD2.n73 VDD2.n72 12.8005
R923 VDD2.n78 VDD2.n4 12.8005
R924 VDD2.n171 VDD2.n170 12.0247
R925 VDD2.n161 VDD2.n98 12.0247
R926 VDD2.n125 VDD2.n116 12.0247
R927 VDD2.n35 VDD2.n26 12.0247
R928 VDD2.n71 VDD2.n8 12.0247
R929 VDD2.n82 VDD2.n81 12.0247
R930 VDD2.n174 VDD2.n91 11.249
R931 VDD2.n158 VDD2.n157 11.249
R932 VDD2.n126 VDD2.n114 11.249
R933 VDD2.n36 VDD2.n24 11.249
R934 VDD2.n68 VDD2.n67 11.249
R935 VDD2.n85 VDD2.n2 11.249
R936 VDD2.n175 VDD2.n89 10.4732
R937 VDD2.n154 VDD2.n100 10.4732
R938 VDD2.n130 VDD2.n129 10.4732
R939 VDD2.n40 VDD2.n39 10.4732
R940 VDD2.n64 VDD2.n10 10.4732
R941 VDD2.n86 VDD2.n0 10.4732
R942 VDD2.n153 VDD2.n102 9.69747
R943 VDD2.n133 VDD2.n112 9.69747
R944 VDD2.n43 VDD2.n22 9.69747
R945 VDD2.n63 VDD2.n12 9.69747
R946 VDD2.n177 VDD2.n176 9.45567
R947 VDD2.n88 VDD2.n87 9.45567
R948 VDD2.n145 VDD2.n144 9.3005
R949 VDD2.n104 VDD2.n103 9.3005
R950 VDD2.n151 VDD2.n150 9.3005
R951 VDD2.n153 VDD2.n152 9.3005
R952 VDD2.n100 VDD2.n99 9.3005
R953 VDD2.n159 VDD2.n158 9.3005
R954 VDD2.n161 VDD2.n160 9.3005
R955 VDD2.n97 VDD2.n94 9.3005
R956 VDD2.n176 VDD2.n175 9.3005
R957 VDD2.n91 VDD2.n90 9.3005
R958 VDD2.n170 VDD2.n169 9.3005
R959 VDD2.n168 VDD2.n167 9.3005
R960 VDD2.n143 VDD2.n142 9.3005
R961 VDD2.n108 VDD2.n107 9.3005
R962 VDD2.n137 VDD2.n136 9.3005
R963 VDD2.n135 VDD2.n134 9.3005
R964 VDD2.n112 VDD2.n111 9.3005
R965 VDD2.n129 VDD2.n128 9.3005
R966 VDD2.n127 VDD2.n126 9.3005
R967 VDD2.n116 VDD2.n115 9.3005
R968 VDD2.n121 VDD2.n120 9.3005
R969 VDD2.n87 VDD2.n86 9.3005
R970 VDD2.n2 VDD2.n1 9.3005
R971 VDD2.n81 VDD2.n80 9.3005
R972 VDD2.n79 VDD2.n78 9.3005
R973 VDD2.n18 VDD2.n17 9.3005
R974 VDD2.n47 VDD2.n46 9.3005
R975 VDD2.n45 VDD2.n44 9.3005
R976 VDD2.n22 VDD2.n21 9.3005
R977 VDD2.n39 VDD2.n38 9.3005
R978 VDD2.n37 VDD2.n36 9.3005
R979 VDD2.n26 VDD2.n25 9.3005
R980 VDD2.n31 VDD2.n30 9.3005
R981 VDD2.n53 VDD2.n52 9.3005
R982 VDD2.n55 VDD2.n54 9.3005
R983 VDD2.n14 VDD2.n13 9.3005
R984 VDD2.n61 VDD2.n60 9.3005
R985 VDD2.n63 VDD2.n62 9.3005
R986 VDD2.n10 VDD2.n9 9.3005
R987 VDD2.n69 VDD2.n68 9.3005
R988 VDD2.n71 VDD2.n70 9.3005
R989 VDD2.n72 VDD2.n5 9.3005
R990 VDD2.n150 VDD2.n149 8.92171
R991 VDD2.n134 VDD2.n110 8.92171
R992 VDD2.n44 VDD2.n20 8.92171
R993 VDD2.n60 VDD2.n59 8.92171
R994 VDD2.n146 VDD2.n104 8.14595
R995 VDD2.n138 VDD2.n137 8.14595
R996 VDD2.n48 VDD2.n47 8.14595
R997 VDD2.n56 VDD2.n14 8.14595
R998 VDD2.n145 VDD2.n106 7.3702
R999 VDD2.n141 VDD2.n108 7.3702
R1000 VDD2.n51 VDD2.n18 7.3702
R1001 VDD2.n55 VDD2.n16 7.3702
R1002 VDD2.n142 VDD2.n106 6.59444
R1003 VDD2.n142 VDD2.n141 6.59444
R1004 VDD2.n52 VDD2.n51 6.59444
R1005 VDD2.n52 VDD2.n16 6.59444
R1006 VDD2.n146 VDD2.n145 5.81868
R1007 VDD2.n138 VDD2.n108 5.81868
R1008 VDD2.n48 VDD2.n18 5.81868
R1009 VDD2.n56 VDD2.n55 5.81868
R1010 VDD2.n149 VDD2.n104 5.04292
R1011 VDD2.n137 VDD2.n110 5.04292
R1012 VDD2.n47 VDD2.n20 5.04292
R1013 VDD2.n59 VDD2.n14 5.04292
R1014 VDD2.n150 VDD2.n102 4.26717
R1015 VDD2.n134 VDD2.n133 4.26717
R1016 VDD2.n44 VDD2.n43 4.26717
R1017 VDD2.n60 VDD2.n12 4.26717
R1018 VDD2.n120 VDD2.n119 3.70982
R1019 VDD2.n30 VDD2.n29 3.70982
R1020 VDD2.n177 VDD2.n89 3.49141
R1021 VDD2.n154 VDD2.n153 3.49141
R1022 VDD2.n130 VDD2.n112 3.49141
R1023 VDD2.n40 VDD2.n22 3.49141
R1024 VDD2.n64 VDD2.n63 3.49141
R1025 VDD2.n88 VDD2.n0 3.49141
R1026 VDD2.n175 VDD2.n174 2.71565
R1027 VDD2.n157 VDD2.n100 2.71565
R1028 VDD2.n129 VDD2.n114 2.71565
R1029 VDD2.n39 VDD2.n24 2.71565
R1030 VDD2.n67 VDD2.n10 2.71565
R1031 VDD2.n86 VDD2.n85 2.71565
R1032 VDD2.n171 VDD2.n91 1.93989
R1033 VDD2.n158 VDD2.n98 1.93989
R1034 VDD2.n126 VDD2.n125 1.93989
R1035 VDD2.n36 VDD2.n35 1.93989
R1036 VDD2.n68 VDD2.n8 1.93989
R1037 VDD2.n82 VDD2.n2 1.93989
R1038 VDD2.n170 VDD2.n93 1.16414
R1039 VDD2.n162 VDD2.n161 1.16414
R1040 VDD2.n122 VDD2.n116 1.16414
R1041 VDD2.n32 VDD2.n26 1.16414
R1042 VDD2.n73 VDD2.n71 1.16414
R1043 VDD2.n81 VDD2.n4 1.16414
R1044 VDD2 VDD2.n178 0.688
R1045 VDD2.n167 VDD2.n166 0.388379
R1046 VDD2.n97 VDD2.n95 0.388379
R1047 VDD2.n121 VDD2.n118 0.388379
R1048 VDD2.n31 VDD2.n28 0.388379
R1049 VDD2.n72 VDD2.n6 0.388379
R1050 VDD2.n78 VDD2.n77 0.388379
R1051 VDD2.n176 VDD2.n90 0.155672
R1052 VDD2.n169 VDD2.n90 0.155672
R1053 VDD2.n169 VDD2.n168 0.155672
R1054 VDD2.n168 VDD2.n94 0.155672
R1055 VDD2.n160 VDD2.n94 0.155672
R1056 VDD2.n160 VDD2.n159 0.155672
R1057 VDD2.n159 VDD2.n99 0.155672
R1058 VDD2.n152 VDD2.n99 0.155672
R1059 VDD2.n152 VDD2.n151 0.155672
R1060 VDD2.n151 VDD2.n103 0.155672
R1061 VDD2.n144 VDD2.n103 0.155672
R1062 VDD2.n144 VDD2.n143 0.155672
R1063 VDD2.n143 VDD2.n107 0.155672
R1064 VDD2.n136 VDD2.n107 0.155672
R1065 VDD2.n136 VDD2.n135 0.155672
R1066 VDD2.n135 VDD2.n111 0.155672
R1067 VDD2.n128 VDD2.n111 0.155672
R1068 VDD2.n128 VDD2.n127 0.155672
R1069 VDD2.n127 VDD2.n115 0.155672
R1070 VDD2.n120 VDD2.n115 0.155672
R1071 VDD2.n30 VDD2.n25 0.155672
R1072 VDD2.n37 VDD2.n25 0.155672
R1073 VDD2.n38 VDD2.n37 0.155672
R1074 VDD2.n38 VDD2.n21 0.155672
R1075 VDD2.n45 VDD2.n21 0.155672
R1076 VDD2.n46 VDD2.n45 0.155672
R1077 VDD2.n46 VDD2.n17 0.155672
R1078 VDD2.n53 VDD2.n17 0.155672
R1079 VDD2.n54 VDD2.n53 0.155672
R1080 VDD2.n54 VDD2.n13 0.155672
R1081 VDD2.n61 VDD2.n13 0.155672
R1082 VDD2.n62 VDD2.n61 0.155672
R1083 VDD2.n62 VDD2.n9 0.155672
R1084 VDD2.n69 VDD2.n9 0.155672
R1085 VDD2.n70 VDD2.n69 0.155672
R1086 VDD2.n70 VDD2.n5 0.155672
R1087 VDD2.n79 VDD2.n5 0.155672
R1088 VDD2.n80 VDD2.n79 0.155672
R1089 VDD2.n80 VDD2.n1 0.155672
R1090 VDD2.n87 VDD2.n1 0.155672
R1091 B.n471 B.n78 585
R1092 B.n473 B.n472 585
R1093 B.n474 B.n77 585
R1094 B.n476 B.n475 585
R1095 B.n477 B.n76 585
R1096 B.n479 B.n478 585
R1097 B.n480 B.n75 585
R1098 B.n482 B.n481 585
R1099 B.n483 B.n74 585
R1100 B.n485 B.n484 585
R1101 B.n486 B.n73 585
R1102 B.n488 B.n487 585
R1103 B.n489 B.n72 585
R1104 B.n491 B.n490 585
R1105 B.n492 B.n71 585
R1106 B.n494 B.n493 585
R1107 B.n495 B.n70 585
R1108 B.n497 B.n496 585
R1109 B.n498 B.n69 585
R1110 B.n500 B.n499 585
R1111 B.n501 B.n68 585
R1112 B.n503 B.n502 585
R1113 B.n504 B.n67 585
R1114 B.n506 B.n505 585
R1115 B.n507 B.n66 585
R1116 B.n509 B.n508 585
R1117 B.n510 B.n65 585
R1118 B.n512 B.n511 585
R1119 B.n513 B.n64 585
R1120 B.n515 B.n514 585
R1121 B.n516 B.n63 585
R1122 B.n518 B.n517 585
R1123 B.n519 B.n62 585
R1124 B.n521 B.n520 585
R1125 B.n522 B.n61 585
R1126 B.n524 B.n523 585
R1127 B.n525 B.n60 585
R1128 B.n527 B.n526 585
R1129 B.n528 B.n59 585
R1130 B.n530 B.n529 585
R1131 B.n531 B.n58 585
R1132 B.n533 B.n532 585
R1133 B.n534 B.n57 585
R1134 B.n536 B.n535 585
R1135 B.n537 B.n56 585
R1136 B.n539 B.n538 585
R1137 B.n540 B.n55 585
R1138 B.n542 B.n541 585
R1139 B.n543 B.n54 585
R1140 B.n545 B.n544 585
R1141 B.n546 B.n53 585
R1142 B.n548 B.n547 585
R1143 B.n549 B.n49 585
R1144 B.n551 B.n550 585
R1145 B.n552 B.n48 585
R1146 B.n554 B.n553 585
R1147 B.n555 B.n47 585
R1148 B.n557 B.n556 585
R1149 B.n558 B.n46 585
R1150 B.n560 B.n559 585
R1151 B.n561 B.n45 585
R1152 B.n563 B.n562 585
R1153 B.n564 B.n44 585
R1154 B.n566 B.n565 585
R1155 B.n568 B.n41 585
R1156 B.n570 B.n569 585
R1157 B.n571 B.n40 585
R1158 B.n573 B.n572 585
R1159 B.n574 B.n39 585
R1160 B.n576 B.n575 585
R1161 B.n577 B.n38 585
R1162 B.n579 B.n578 585
R1163 B.n580 B.n37 585
R1164 B.n582 B.n581 585
R1165 B.n583 B.n36 585
R1166 B.n585 B.n584 585
R1167 B.n586 B.n35 585
R1168 B.n588 B.n587 585
R1169 B.n589 B.n34 585
R1170 B.n591 B.n590 585
R1171 B.n592 B.n33 585
R1172 B.n594 B.n593 585
R1173 B.n595 B.n32 585
R1174 B.n597 B.n596 585
R1175 B.n598 B.n31 585
R1176 B.n600 B.n599 585
R1177 B.n601 B.n30 585
R1178 B.n603 B.n602 585
R1179 B.n604 B.n29 585
R1180 B.n606 B.n605 585
R1181 B.n607 B.n28 585
R1182 B.n609 B.n608 585
R1183 B.n610 B.n27 585
R1184 B.n612 B.n611 585
R1185 B.n613 B.n26 585
R1186 B.n615 B.n614 585
R1187 B.n616 B.n25 585
R1188 B.n618 B.n617 585
R1189 B.n619 B.n24 585
R1190 B.n621 B.n620 585
R1191 B.n622 B.n23 585
R1192 B.n624 B.n623 585
R1193 B.n625 B.n22 585
R1194 B.n627 B.n626 585
R1195 B.n628 B.n21 585
R1196 B.n630 B.n629 585
R1197 B.n631 B.n20 585
R1198 B.n633 B.n632 585
R1199 B.n634 B.n19 585
R1200 B.n636 B.n635 585
R1201 B.n637 B.n18 585
R1202 B.n639 B.n638 585
R1203 B.n640 B.n17 585
R1204 B.n642 B.n641 585
R1205 B.n643 B.n16 585
R1206 B.n645 B.n644 585
R1207 B.n646 B.n15 585
R1208 B.n648 B.n647 585
R1209 B.n470 B.n469 585
R1210 B.n468 B.n79 585
R1211 B.n467 B.n466 585
R1212 B.n465 B.n80 585
R1213 B.n464 B.n463 585
R1214 B.n462 B.n81 585
R1215 B.n461 B.n460 585
R1216 B.n459 B.n82 585
R1217 B.n458 B.n457 585
R1218 B.n456 B.n83 585
R1219 B.n455 B.n454 585
R1220 B.n453 B.n84 585
R1221 B.n452 B.n451 585
R1222 B.n450 B.n85 585
R1223 B.n449 B.n448 585
R1224 B.n447 B.n86 585
R1225 B.n446 B.n445 585
R1226 B.n444 B.n87 585
R1227 B.n443 B.n442 585
R1228 B.n441 B.n88 585
R1229 B.n440 B.n439 585
R1230 B.n438 B.n89 585
R1231 B.n437 B.n436 585
R1232 B.n435 B.n90 585
R1233 B.n434 B.n433 585
R1234 B.n432 B.n91 585
R1235 B.n431 B.n430 585
R1236 B.n429 B.n92 585
R1237 B.n428 B.n427 585
R1238 B.n426 B.n93 585
R1239 B.n425 B.n424 585
R1240 B.n423 B.n94 585
R1241 B.n422 B.n421 585
R1242 B.n420 B.n95 585
R1243 B.n419 B.n418 585
R1244 B.n417 B.n96 585
R1245 B.n416 B.n415 585
R1246 B.n414 B.n97 585
R1247 B.n413 B.n412 585
R1248 B.n411 B.n98 585
R1249 B.n410 B.n409 585
R1250 B.n408 B.n99 585
R1251 B.n407 B.n406 585
R1252 B.n405 B.n100 585
R1253 B.n404 B.n403 585
R1254 B.n402 B.n101 585
R1255 B.n401 B.n400 585
R1256 B.n399 B.n102 585
R1257 B.n398 B.n397 585
R1258 B.n396 B.n103 585
R1259 B.n395 B.n394 585
R1260 B.n216 B.n167 585
R1261 B.n218 B.n217 585
R1262 B.n219 B.n166 585
R1263 B.n221 B.n220 585
R1264 B.n222 B.n165 585
R1265 B.n224 B.n223 585
R1266 B.n225 B.n164 585
R1267 B.n227 B.n226 585
R1268 B.n228 B.n163 585
R1269 B.n230 B.n229 585
R1270 B.n231 B.n162 585
R1271 B.n233 B.n232 585
R1272 B.n234 B.n161 585
R1273 B.n236 B.n235 585
R1274 B.n237 B.n160 585
R1275 B.n239 B.n238 585
R1276 B.n240 B.n159 585
R1277 B.n242 B.n241 585
R1278 B.n243 B.n158 585
R1279 B.n245 B.n244 585
R1280 B.n246 B.n157 585
R1281 B.n248 B.n247 585
R1282 B.n249 B.n156 585
R1283 B.n251 B.n250 585
R1284 B.n252 B.n155 585
R1285 B.n254 B.n253 585
R1286 B.n255 B.n154 585
R1287 B.n257 B.n256 585
R1288 B.n258 B.n153 585
R1289 B.n260 B.n259 585
R1290 B.n261 B.n152 585
R1291 B.n263 B.n262 585
R1292 B.n264 B.n151 585
R1293 B.n266 B.n265 585
R1294 B.n267 B.n150 585
R1295 B.n269 B.n268 585
R1296 B.n270 B.n149 585
R1297 B.n272 B.n271 585
R1298 B.n273 B.n148 585
R1299 B.n275 B.n274 585
R1300 B.n276 B.n147 585
R1301 B.n278 B.n277 585
R1302 B.n279 B.n146 585
R1303 B.n281 B.n280 585
R1304 B.n282 B.n145 585
R1305 B.n284 B.n283 585
R1306 B.n285 B.n144 585
R1307 B.n287 B.n286 585
R1308 B.n288 B.n143 585
R1309 B.n290 B.n289 585
R1310 B.n291 B.n142 585
R1311 B.n293 B.n292 585
R1312 B.n294 B.n141 585
R1313 B.n296 B.n295 585
R1314 B.n298 B.n138 585
R1315 B.n300 B.n299 585
R1316 B.n301 B.n137 585
R1317 B.n303 B.n302 585
R1318 B.n304 B.n136 585
R1319 B.n306 B.n305 585
R1320 B.n307 B.n135 585
R1321 B.n309 B.n308 585
R1322 B.n310 B.n134 585
R1323 B.n312 B.n311 585
R1324 B.n314 B.n313 585
R1325 B.n315 B.n130 585
R1326 B.n317 B.n316 585
R1327 B.n318 B.n129 585
R1328 B.n320 B.n319 585
R1329 B.n321 B.n128 585
R1330 B.n323 B.n322 585
R1331 B.n324 B.n127 585
R1332 B.n326 B.n325 585
R1333 B.n327 B.n126 585
R1334 B.n329 B.n328 585
R1335 B.n330 B.n125 585
R1336 B.n332 B.n331 585
R1337 B.n333 B.n124 585
R1338 B.n335 B.n334 585
R1339 B.n336 B.n123 585
R1340 B.n338 B.n337 585
R1341 B.n339 B.n122 585
R1342 B.n341 B.n340 585
R1343 B.n342 B.n121 585
R1344 B.n344 B.n343 585
R1345 B.n345 B.n120 585
R1346 B.n347 B.n346 585
R1347 B.n348 B.n119 585
R1348 B.n350 B.n349 585
R1349 B.n351 B.n118 585
R1350 B.n353 B.n352 585
R1351 B.n354 B.n117 585
R1352 B.n356 B.n355 585
R1353 B.n357 B.n116 585
R1354 B.n359 B.n358 585
R1355 B.n360 B.n115 585
R1356 B.n362 B.n361 585
R1357 B.n363 B.n114 585
R1358 B.n365 B.n364 585
R1359 B.n366 B.n113 585
R1360 B.n368 B.n367 585
R1361 B.n369 B.n112 585
R1362 B.n371 B.n370 585
R1363 B.n372 B.n111 585
R1364 B.n374 B.n373 585
R1365 B.n375 B.n110 585
R1366 B.n377 B.n376 585
R1367 B.n378 B.n109 585
R1368 B.n380 B.n379 585
R1369 B.n381 B.n108 585
R1370 B.n383 B.n382 585
R1371 B.n384 B.n107 585
R1372 B.n386 B.n385 585
R1373 B.n387 B.n106 585
R1374 B.n389 B.n388 585
R1375 B.n390 B.n105 585
R1376 B.n392 B.n391 585
R1377 B.n393 B.n104 585
R1378 B.n215 B.n214 585
R1379 B.n213 B.n168 585
R1380 B.n212 B.n211 585
R1381 B.n210 B.n169 585
R1382 B.n209 B.n208 585
R1383 B.n207 B.n170 585
R1384 B.n206 B.n205 585
R1385 B.n204 B.n171 585
R1386 B.n203 B.n202 585
R1387 B.n201 B.n172 585
R1388 B.n200 B.n199 585
R1389 B.n198 B.n173 585
R1390 B.n197 B.n196 585
R1391 B.n195 B.n174 585
R1392 B.n194 B.n193 585
R1393 B.n192 B.n175 585
R1394 B.n191 B.n190 585
R1395 B.n189 B.n176 585
R1396 B.n188 B.n187 585
R1397 B.n186 B.n177 585
R1398 B.n185 B.n184 585
R1399 B.n183 B.n178 585
R1400 B.n182 B.n181 585
R1401 B.n180 B.n179 585
R1402 B.n2 B.n0 585
R1403 B.n685 B.n1 585
R1404 B.n684 B.n683 585
R1405 B.n682 B.n3 585
R1406 B.n681 B.n680 585
R1407 B.n679 B.n4 585
R1408 B.n678 B.n677 585
R1409 B.n676 B.n5 585
R1410 B.n675 B.n674 585
R1411 B.n673 B.n6 585
R1412 B.n672 B.n671 585
R1413 B.n670 B.n7 585
R1414 B.n669 B.n668 585
R1415 B.n667 B.n8 585
R1416 B.n666 B.n665 585
R1417 B.n664 B.n9 585
R1418 B.n663 B.n662 585
R1419 B.n661 B.n10 585
R1420 B.n660 B.n659 585
R1421 B.n658 B.n11 585
R1422 B.n657 B.n656 585
R1423 B.n655 B.n12 585
R1424 B.n654 B.n653 585
R1425 B.n652 B.n13 585
R1426 B.n651 B.n650 585
R1427 B.n649 B.n14 585
R1428 B.n687 B.n686 585
R1429 B.n216 B.n215 535.745
R1430 B.n649 B.n648 535.745
R1431 B.n395 B.n104 535.745
R1432 B.n469 B.n78 535.745
R1433 B.n131 B.t5 509.137
R1434 B.n50 B.t7 509.137
R1435 B.n139 B.t11 509.137
R1436 B.n42 B.t1 509.137
R1437 B.n132 B.t4 452.507
R1438 B.n51 B.t8 452.507
R1439 B.n140 B.t10 452.507
R1440 B.n43 B.t2 452.507
R1441 B.n131 B.t3 359.332
R1442 B.n139 B.t9 359.332
R1443 B.n42 B.t0 359.332
R1444 B.n50 B.t6 359.332
R1445 B.n215 B.n168 163.367
R1446 B.n211 B.n168 163.367
R1447 B.n211 B.n210 163.367
R1448 B.n210 B.n209 163.367
R1449 B.n209 B.n170 163.367
R1450 B.n205 B.n170 163.367
R1451 B.n205 B.n204 163.367
R1452 B.n204 B.n203 163.367
R1453 B.n203 B.n172 163.367
R1454 B.n199 B.n172 163.367
R1455 B.n199 B.n198 163.367
R1456 B.n198 B.n197 163.367
R1457 B.n197 B.n174 163.367
R1458 B.n193 B.n174 163.367
R1459 B.n193 B.n192 163.367
R1460 B.n192 B.n191 163.367
R1461 B.n191 B.n176 163.367
R1462 B.n187 B.n176 163.367
R1463 B.n187 B.n186 163.367
R1464 B.n186 B.n185 163.367
R1465 B.n185 B.n178 163.367
R1466 B.n181 B.n178 163.367
R1467 B.n181 B.n180 163.367
R1468 B.n180 B.n2 163.367
R1469 B.n686 B.n2 163.367
R1470 B.n686 B.n685 163.367
R1471 B.n685 B.n684 163.367
R1472 B.n684 B.n3 163.367
R1473 B.n680 B.n3 163.367
R1474 B.n680 B.n679 163.367
R1475 B.n679 B.n678 163.367
R1476 B.n678 B.n5 163.367
R1477 B.n674 B.n5 163.367
R1478 B.n674 B.n673 163.367
R1479 B.n673 B.n672 163.367
R1480 B.n672 B.n7 163.367
R1481 B.n668 B.n7 163.367
R1482 B.n668 B.n667 163.367
R1483 B.n667 B.n666 163.367
R1484 B.n666 B.n9 163.367
R1485 B.n662 B.n9 163.367
R1486 B.n662 B.n661 163.367
R1487 B.n661 B.n660 163.367
R1488 B.n660 B.n11 163.367
R1489 B.n656 B.n11 163.367
R1490 B.n656 B.n655 163.367
R1491 B.n655 B.n654 163.367
R1492 B.n654 B.n13 163.367
R1493 B.n650 B.n13 163.367
R1494 B.n650 B.n649 163.367
R1495 B.n217 B.n216 163.367
R1496 B.n217 B.n166 163.367
R1497 B.n221 B.n166 163.367
R1498 B.n222 B.n221 163.367
R1499 B.n223 B.n222 163.367
R1500 B.n223 B.n164 163.367
R1501 B.n227 B.n164 163.367
R1502 B.n228 B.n227 163.367
R1503 B.n229 B.n228 163.367
R1504 B.n229 B.n162 163.367
R1505 B.n233 B.n162 163.367
R1506 B.n234 B.n233 163.367
R1507 B.n235 B.n234 163.367
R1508 B.n235 B.n160 163.367
R1509 B.n239 B.n160 163.367
R1510 B.n240 B.n239 163.367
R1511 B.n241 B.n240 163.367
R1512 B.n241 B.n158 163.367
R1513 B.n245 B.n158 163.367
R1514 B.n246 B.n245 163.367
R1515 B.n247 B.n246 163.367
R1516 B.n247 B.n156 163.367
R1517 B.n251 B.n156 163.367
R1518 B.n252 B.n251 163.367
R1519 B.n253 B.n252 163.367
R1520 B.n253 B.n154 163.367
R1521 B.n257 B.n154 163.367
R1522 B.n258 B.n257 163.367
R1523 B.n259 B.n258 163.367
R1524 B.n259 B.n152 163.367
R1525 B.n263 B.n152 163.367
R1526 B.n264 B.n263 163.367
R1527 B.n265 B.n264 163.367
R1528 B.n265 B.n150 163.367
R1529 B.n269 B.n150 163.367
R1530 B.n270 B.n269 163.367
R1531 B.n271 B.n270 163.367
R1532 B.n271 B.n148 163.367
R1533 B.n275 B.n148 163.367
R1534 B.n276 B.n275 163.367
R1535 B.n277 B.n276 163.367
R1536 B.n277 B.n146 163.367
R1537 B.n281 B.n146 163.367
R1538 B.n282 B.n281 163.367
R1539 B.n283 B.n282 163.367
R1540 B.n283 B.n144 163.367
R1541 B.n287 B.n144 163.367
R1542 B.n288 B.n287 163.367
R1543 B.n289 B.n288 163.367
R1544 B.n289 B.n142 163.367
R1545 B.n293 B.n142 163.367
R1546 B.n294 B.n293 163.367
R1547 B.n295 B.n294 163.367
R1548 B.n295 B.n138 163.367
R1549 B.n300 B.n138 163.367
R1550 B.n301 B.n300 163.367
R1551 B.n302 B.n301 163.367
R1552 B.n302 B.n136 163.367
R1553 B.n306 B.n136 163.367
R1554 B.n307 B.n306 163.367
R1555 B.n308 B.n307 163.367
R1556 B.n308 B.n134 163.367
R1557 B.n312 B.n134 163.367
R1558 B.n313 B.n312 163.367
R1559 B.n313 B.n130 163.367
R1560 B.n317 B.n130 163.367
R1561 B.n318 B.n317 163.367
R1562 B.n319 B.n318 163.367
R1563 B.n319 B.n128 163.367
R1564 B.n323 B.n128 163.367
R1565 B.n324 B.n323 163.367
R1566 B.n325 B.n324 163.367
R1567 B.n325 B.n126 163.367
R1568 B.n329 B.n126 163.367
R1569 B.n330 B.n329 163.367
R1570 B.n331 B.n330 163.367
R1571 B.n331 B.n124 163.367
R1572 B.n335 B.n124 163.367
R1573 B.n336 B.n335 163.367
R1574 B.n337 B.n336 163.367
R1575 B.n337 B.n122 163.367
R1576 B.n341 B.n122 163.367
R1577 B.n342 B.n341 163.367
R1578 B.n343 B.n342 163.367
R1579 B.n343 B.n120 163.367
R1580 B.n347 B.n120 163.367
R1581 B.n348 B.n347 163.367
R1582 B.n349 B.n348 163.367
R1583 B.n349 B.n118 163.367
R1584 B.n353 B.n118 163.367
R1585 B.n354 B.n353 163.367
R1586 B.n355 B.n354 163.367
R1587 B.n355 B.n116 163.367
R1588 B.n359 B.n116 163.367
R1589 B.n360 B.n359 163.367
R1590 B.n361 B.n360 163.367
R1591 B.n361 B.n114 163.367
R1592 B.n365 B.n114 163.367
R1593 B.n366 B.n365 163.367
R1594 B.n367 B.n366 163.367
R1595 B.n367 B.n112 163.367
R1596 B.n371 B.n112 163.367
R1597 B.n372 B.n371 163.367
R1598 B.n373 B.n372 163.367
R1599 B.n373 B.n110 163.367
R1600 B.n377 B.n110 163.367
R1601 B.n378 B.n377 163.367
R1602 B.n379 B.n378 163.367
R1603 B.n379 B.n108 163.367
R1604 B.n383 B.n108 163.367
R1605 B.n384 B.n383 163.367
R1606 B.n385 B.n384 163.367
R1607 B.n385 B.n106 163.367
R1608 B.n389 B.n106 163.367
R1609 B.n390 B.n389 163.367
R1610 B.n391 B.n390 163.367
R1611 B.n391 B.n104 163.367
R1612 B.n396 B.n395 163.367
R1613 B.n397 B.n396 163.367
R1614 B.n397 B.n102 163.367
R1615 B.n401 B.n102 163.367
R1616 B.n402 B.n401 163.367
R1617 B.n403 B.n402 163.367
R1618 B.n403 B.n100 163.367
R1619 B.n407 B.n100 163.367
R1620 B.n408 B.n407 163.367
R1621 B.n409 B.n408 163.367
R1622 B.n409 B.n98 163.367
R1623 B.n413 B.n98 163.367
R1624 B.n414 B.n413 163.367
R1625 B.n415 B.n414 163.367
R1626 B.n415 B.n96 163.367
R1627 B.n419 B.n96 163.367
R1628 B.n420 B.n419 163.367
R1629 B.n421 B.n420 163.367
R1630 B.n421 B.n94 163.367
R1631 B.n425 B.n94 163.367
R1632 B.n426 B.n425 163.367
R1633 B.n427 B.n426 163.367
R1634 B.n427 B.n92 163.367
R1635 B.n431 B.n92 163.367
R1636 B.n432 B.n431 163.367
R1637 B.n433 B.n432 163.367
R1638 B.n433 B.n90 163.367
R1639 B.n437 B.n90 163.367
R1640 B.n438 B.n437 163.367
R1641 B.n439 B.n438 163.367
R1642 B.n439 B.n88 163.367
R1643 B.n443 B.n88 163.367
R1644 B.n444 B.n443 163.367
R1645 B.n445 B.n444 163.367
R1646 B.n445 B.n86 163.367
R1647 B.n449 B.n86 163.367
R1648 B.n450 B.n449 163.367
R1649 B.n451 B.n450 163.367
R1650 B.n451 B.n84 163.367
R1651 B.n455 B.n84 163.367
R1652 B.n456 B.n455 163.367
R1653 B.n457 B.n456 163.367
R1654 B.n457 B.n82 163.367
R1655 B.n461 B.n82 163.367
R1656 B.n462 B.n461 163.367
R1657 B.n463 B.n462 163.367
R1658 B.n463 B.n80 163.367
R1659 B.n467 B.n80 163.367
R1660 B.n468 B.n467 163.367
R1661 B.n469 B.n468 163.367
R1662 B.n648 B.n15 163.367
R1663 B.n644 B.n15 163.367
R1664 B.n644 B.n643 163.367
R1665 B.n643 B.n642 163.367
R1666 B.n642 B.n17 163.367
R1667 B.n638 B.n17 163.367
R1668 B.n638 B.n637 163.367
R1669 B.n637 B.n636 163.367
R1670 B.n636 B.n19 163.367
R1671 B.n632 B.n19 163.367
R1672 B.n632 B.n631 163.367
R1673 B.n631 B.n630 163.367
R1674 B.n630 B.n21 163.367
R1675 B.n626 B.n21 163.367
R1676 B.n626 B.n625 163.367
R1677 B.n625 B.n624 163.367
R1678 B.n624 B.n23 163.367
R1679 B.n620 B.n23 163.367
R1680 B.n620 B.n619 163.367
R1681 B.n619 B.n618 163.367
R1682 B.n618 B.n25 163.367
R1683 B.n614 B.n25 163.367
R1684 B.n614 B.n613 163.367
R1685 B.n613 B.n612 163.367
R1686 B.n612 B.n27 163.367
R1687 B.n608 B.n27 163.367
R1688 B.n608 B.n607 163.367
R1689 B.n607 B.n606 163.367
R1690 B.n606 B.n29 163.367
R1691 B.n602 B.n29 163.367
R1692 B.n602 B.n601 163.367
R1693 B.n601 B.n600 163.367
R1694 B.n600 B.n31 163.367
R1695 B.n596 B.n31 163.367
R1696 B.n596 B.n595 163.367
R1697 B.n595 B.n594 163.367
R1698 B.n594 B.n33 163.367
R1699 B.n590 B.n33 163.367
R1700 B.n590 B.n589 163.367
R1701 B.n589 B.n588 163.367
R1702 B.n588 B.n35 163.367
R1703 B.n584 B.n35 163.367
R1704 B.n584 B.n583 163.367
R1705 B.n583 B.n582 163.367
R1706 B.n582 B.n37 163.367
R1707 B.n578 B.n37 163.367
R1708 B.n578 B.n577 163.367
R1709 B.n577 B.n576 163.367
R1710 B.n576 B.n39 163.367
R1711 B.n572 B.n39 163.367
R1712 B.n572 B.n571 163.367
R1713 B.n571 B.n570 163.367
R1714 B.n570 B.n41 163.367
R1715 B.n565 B.n41 163.367
R1716 B.n565 B.n564 163.367
R1717 B.n564 B.n563 163.367
R1718 B.n563 B.n45 163.367
R1719 B.n559 B.n45 163.367
R1720 B.n559 B.n558 163.367
R1721 B.n558 B.n557 163.367
R1722 B.n557 B.n47 163.367
R1723 B.n553 B.n47 163.367
R1724 B.n553 B.n552 163.367
R1725 B.n552 B.n551 163.367
R1726 B.n551 B.n49 163.367
R1727 B.n547 B.n49 163.367
R1728 B.n547 B.n546 163.367
R1729 B.n546 B.n545 163.367
R1730 B.n545 B.n54 163.367
R1731 B.n541 B.n54 163.367
R1732 B.n541 B.n540 163.367
R1733 B.n540 B.n539 163.367
R1734 B.n539 B.n56 163.367
R1735 B.n535 B.n56 163.367
R1736 B.n535 B.n534 163.367
R1737 B.n534 B.n533 163.367
R1738 B.n533 B.n58 163.367
R1739 B.n529 B.n58 163.367
R1740 B.n529 B.n528 163.367
R1741 B.n528 B.n527 163.367
R1742 B.n527 B.n60 163.367
R1743 B.n523 B.n60 163.367
R1744 B.n523 B.n522 163.367
R1745 B.n522 B.n521 163.367
R1746 B.n521 B.n62 163.367
R1747 B.n517 B.n62 163.367
R1748 B.n517 B.n516 163.367
R1749 B.n516 B.n515 163.367
R1750 B.n515 B.n64 163.367
R1751 B.n511 B.n64 163.367
R1752 B.n511 B.n510 163.367
R1753 B.n510 B.n509 163.367
R1754 B.n509 B.n66 163.367
R1755 B.n505 B.n66 163.367
R1756 B.n505 B.n504 163.367
R1757 B.n504 B.n503 163.367
R1758 B.n503 B.n68 163.367
R1759 B.n499 B.n68 163.367
R1760 B.n499 B.n498 163.367
R1761 B.n498 B.n497 163.367
R1762 B.n497 B.n70 163.367
R1763 B.n493 B.n70 163.367
R1764 B.n493 B.n492 163.367
R1765 B.n492 B.n491 163.367
R1766 B.n491 B.n72 163.367
R1767 B.n487 B.n72 163.367
R1768 B.n487 B.n486 163.367
R1769 B.n486 B.n485 163.367
R1770 B.n485 B.n74 163.367
R1771 B.n481 B.n74 163.367
R1772 B.n481 B.n480 163.367
R1773 B.n480 B.n479 163.367
R1774 B.n479 B.n76 163.367
R1775 B.n475 B.n76 163.367
R1776 B.n475 B.n474 163.367
R1777 B.n474 B.n473 163.367
R1778 B.n473 B.n78 163.367
R1779 B.n133 B.n132 59.5399
R1780 B.n297 B.n140 59.5399
R1781 B.n567 B.n43 59.5399
R1782 B.n52 B.n51 59.5399
R1783 B.n132 B.n131 56.6308
R1784 B.n140 B.n139 56.6308
R1785 B.n43 B.n42 56.6308
R1786 B.n51 B.n50 56.6308
R1787 B.n647 B.n14 34.8103
R1788 B.n471 B.n470 34.8103
R1789 B.n394 B.n393 34.8103
R1790 B.n214 B.n167 34.8103
R1791 B B.n687 18.0485
R1792 B.n647 B.n646 10.6151
R1793 B.n646 B.n645 10.6151
R1794 B.n645 B.n16 10.6151
R1795 B.n641 B.n16 10.6151
R1796 B.n641 B.n640 10.6151
R1797 B.n640 B.n639 10.6151
R1798 B.n639 B.n18 10.6151
R1799 B.n635 B.n18 10.6151
R1800 B.n635 B.n634 10.6151
R1801 B.n634 B.n633 10.6151
R1802 B.n633 B.n20 10.6151
R1803 B.n629 B.n20 10.6151
R1804 B.n629 B.n628 10.6151
R1805 B.n628 B.n627 10.6151
R1806 B.n627 B.n22 10.6151
R1807 B.n623 B.n22 10.6151
R1808 B.n623 B.n622 10.6151
R1809 B.n622 B.n621 10.6151
R1810 B.n621 B.n24 10.6151
R1811 B.n617 B.n24 10.6151
R1812 B.n617 B.n616 10.6151
R1813 B.n616 B.n615 10.6151
R1814 B.n615 B.n26 10.6151
R1815 B.n611 B.n26 10.6151
R1816 B.n611 B.n610 10.6151
R1817 B.n610 B.n609 10.6151
R1818 B.n609 B.n28 10.6151
R1819 B.n605 B.n28 10.6151
R1820 B.n605 B.n604 10.6151
R1821 B.n604 B.n603 10.6151
R1822 B.n603 B.n30 10.6151
R1823 B.n599 B.n30 10.6151
R1824 B.n599 B.n598 10.6151
R1825 B.n598 B.n597 10.6151
R1826 B.n597 B.n32 10.6151
R1827 B.n593 B.n32 10.6151
R1828 B.n593 B.n592 10.6151
R1829 B.n592 B.n591 10.6151
R1830 B.n591 B.n34 10.6151
R1831 B.n587 B.n34 10.6151
R1832 B.n587 B.n586 10.6151
R1833 B.n586 B.n585 10.6151
R1834 B.n585 B.n36 10.6151
R1835 B.n581 B.n36 10.6151
R1836 B.n581 B.n580 10.6151
R1837 B.n580 B.n579 10.6151
R1838 B.n579 B.n38 10.6151
R1839 B.n575 B.n38 10.6151
R1840 B.n575 B.n574 10.6151
R1841 B.n574 B.n573 10.6151
R1842 B.n573 B.n40 10.6151
R1843 B.n569 B.n40 10.6151
R1844 B.n569 B.n568 10.6151
R1845 B.n566 B.n44 10.6151
R1846 B.n562 B.n44 10.6151
R1847 B.n562 B.n561 10.6151
R1848 B.n561 B.n560 10.6151
R1849 B.n560 B.n46 10.6151
R1850 B.n556 B.n46 10.6151
R1851 B.n556 B.n555 10.6151
R1852 B.n555 B.n554 10.6151
R1853 B.n554 B.n48 10.6151
R1854 B.n550 B.n549 10.6151
R1855 B.n549 B.n548 10.6151
R1856 B.n548 B.n53 10.6151
R1857 B.n544 B.n53 10.6151
R1858 B.n544 B.n543 10.6151
R1859 B.n543 B.n542 10.6151
R1860 B.n542 B.n55 10.6151
R1861 B.n538 B.n55 10.6151
R1862 B.n538 B.n537 10.6151
R1863 B.n537 B.n536 10.6151
R1864 B.n536 B.n57 10.6151
R1865 B.n532 B.n57 10.6151
R1866 B.n532 B.n531 10.6151
R1867 B.n531 B.n530 10.6151
R1868 B.n530 B.n59 10.6151
R1869 B.n526 B.n59 10.6151
R1870 B.n526 B.n525 10.6151
R1871 B.n525 B.n524 10.6151
R1872 B.n524 B.n61 10.6151
R1873 B.n520 B.n61 10.6151
R1874 B.n520 B.n519 10.6151
R1875 B.n519 B.n518 10.6151
R1876 B.n518 B.n63 10.6151
R1877 B.n514 B.n63 10.6151
R1878 B.n514 B.n513 10.6151
R1879 B.n513 B.n512 10.6151
R1880 B.n512 B.n65 10.6151
R1881 B.n508 B.n65 10.6151
R1882 B.n508 B.n507 10.6151
R1883 B.n507 B.n506 10.6151
R1884 B.n506 B.n67 10.6151
R1885 B.n502 B.n67 10.6151
R1886 B.n502 B.n501 10.6151
R1887 B.n501 B.n500 10.6151
R1888 B.n500 B.n69 10.6151
R1889 B.n496 B.n69 10.6151
R1890 B.n496 B.n495 10.6151
R1891 B.n495 B.n494 10.6151
R1892 B.n494 B.n71 10.6151
R1893 B.n490 B.n71 10.6151
R1894 B.n490 B.n489 10.6151
R1895 B.n489 B.n488 10.6151
R1896 B.n488 B.n73 10.6151
R1897 B.n484 B.n73 10.6151
R1898 B.n484 B.n483 10.6151
R1899 B.n483 B.n482 10.6151
R1900 B.n482 B.n75 10.6151
R1901 B.n478 B.n75 10.6151
R1902 B.n478 B.n477 10.6151
R1903 B.n477 B.n476 10.6151
R1904 B.n476 B.n77 10.6151
R1905 B.n472 B.n77 10.6151
R1906 B.n472 B.n471 10.6151
R1907 B.n394 B.n103 10.6151
R1908 B.n398 B.n103 10.6151
R1909 B.n399 B.n398 10.6151
R1910 B.n400 B.n399 10.6151
R1911 B.n400 B.n101 10.6151
R1912 B.n404 B.n101 10.6151
R1913 B.n405 B.n404 10.6151
R1914 B.n406 B.n405 10.6151
R1915 B.n406 B.n99 10.6151
R1916 B.n410 B.n99 10.6151
R1917 B.n411 B.n410 10.6151
R1918 B.n412 B.n411 10.6151
R1919 B.n412 B.n97 10.6151
R1920 B.n416 B.n97 10.6151
R1921 B.n417 B.n416 10.6151
R1922 B.n418 B.n417 10.6151
R1923 B.n418 B.n95 10.6151
R1924 B.n422 B.n95 10.6151
R1925 B.n423 B.n422 10.6151
R1926 B.n424 B.n423 10.6151
R1927 B.n424 B.n93 10.6151
R1928 B.n428 B.n93 10.6151
R1929 B.n429 B.n428 10.6151
R1930 B.n430 B.n429 10.6151
R1931 B.n430 B.n91 10.6151
R1932 B.n434 B.n91 10.6151
R1933 B.n435 B.n434 10.6151
R1934 B.n436 B.n435 10.6151
R1935 B.n436 B.n89 10.6151
R1936 B.n440 B.n89 10.6151
R1937 B.n441 B.n440 10.6151
R1938 B.n442 B.n441 10.6151
R1939 B.n442 B.n87 10.6151
R1940 B.n446 B.n87 10.6151
R1941 B.n447 B.n446 10.6151
R1942 B.n448 B.n447 10.6151
R1943 B.n448 B.n85 10.6151
R1944 B.n452 B.n85 10.6151
R1945 B.n453 B.n452 10.6151
R1946 B.n454 B.n453 10.6151
R1947 B.n454 B.n83 10.6151
R1948 B.n458 B.n83 10.6151
R1949 B.n459 B.n458 10.6151
R1950 B.n460 B.n459 10.6151
R1951 B.n460 B.n81 10.6151
R1952 B.n464 B.n81 10.6151
R1953 B.n465 B.n464 10.6151
R1954 B.n466 B.n465 10.6151
R1955 B.n466 B.n79 10.6151
R1956 B.n470 B.n79 10.6151
R1957 B.n218 B.n167 10.6151
R1958 B.n219 B.n218 10.6151
R1959 B.n220 B.n219 10.6151
R1960 B.n220 B.n165 10.6151
R1961 B.n224 B.n165 10.6151
R1962 B.n225 B.n224 10.6151
R1963 B.n226 B.n225 10.6151
R1964 B.n226 B.n163 10.6151
R1965 B.n230 B.n163 10.6151
R1966 B.n231 B.n230 10.6151
R1967 B.n232 B.n231 10.6151
R1968 B.n232 B.n161 10.6151
R1969 B.n236 B.n161 10.6151
R1970 B.n237 B.n236 10.6151
R1971 B.n238 B.n237 10.6151
R1972 B.n238 B.n159 10.6151
R1973 B.n242 B.n159 10.6151
R1974 B.n243 B.n242 10.6151
R1975 B.n244 B.n243 10.6151
R1976 B.n244 B.n157 10.6151
R1977 B.n248 B.n157 10.6151
R1978 B.n249 B.n248 10.6151
R1979 B.n250 B.n249 10.6151
R1980 B.n250 B.n155 10.6151
R1981 B.n254 B.n155 10.6151
R1982 B.n255 B.n254 10.6151
R1983 B.n256 B.n255 10.6151
R1984 B.n256 B.n153 10.6151
R1985 B.n260 B.n153 10.6151
R1986 B.n261 B.n260 10.6151
R1987 B.n262 B.n261 10.6151
R1988 B.n262 B.n151 10.6151
R1989 B.n266 B.n151 10.6151
R1990 B.n267 B.n266 10.6151
R1991 B.n268 B.n267 10.6151
R1992 B.n268 B.n149 10.6151
R1993 B.n272 B.n149 10.6151
R1994 B.n273 B.n272 10.6151
R1995 B.n274 B.n273 10.6151
R1996 B.n274 B.n147 10.6151
R1997 B.n278 B.n147 10.6151
R1998 B.n279 B.n278 10.6151
R1999 B.n280 B.n279 10.6151
R2000 B.n280 B.n145 10.6151
R2001 B.n284 B.n145 10.6151
R2002 B.n285 B.n284 10.6151
R2003 B.n286 B.n285 10.6151
R2004 B.n286 B.n143 10.6151
R2005 B.n290 B.n143 10.6151
R2006 B.n291 B.n290 10.6151
R2007 B.n292 B.n291 10.6151
R2008 B.n292 B.n141 10.6151
R2009 B.n296 B.n141 10.6151
R2010 B.n299 B.n298 10.6151
R2011 B.n299 B.n137 10.6151
R2012 B.n303 B.n137 10.6151
R2013 B.n304 B.n303 10.6151
R2014 B.n305 B.n304 10.6151
R2015 B.n305 B.n135 10.6151
R2016 B.n309 B.n135 10.6151
R2017 B.n310 B.n309 10.6151
R2018 B.n311 B.n310 10.6151
R2019 B.n315 B.n314 10.6151
R2020 B.n316 B.n315 10.6151
R2021 B.n316 B.n129 10.6151
R2022 B.n320 B.n129 10.6151
R2023 B.n321 B.n320 10.6151
R2024 B.n322 B.n321 10.6151
R2025 B.n322 B.n127 10.6151
R2026 B.n326 B.n127 10.6151
R2027 B.n327 B.n326 10.6151
R2028 B.n328 B.n327 10.6151
R2029 B.n328 B.n125 10.6151
R2030 B.n332 B.n125 10.6151
R2031 B.n333 B.n332 10.6151
R2032 B.n334 B.n333 10.6151
R2033 B.n334 B.n123 10.6151
R2034 B.n338 B.n123 10.6151
R2035 B.n339 B.n338 10.6151
R2036 B.n340 B.n339 10.6151
R2037 B.n340 B.n121 10.6151
R2038 B.n344 B.n121 10.6151
R2039 B.n345 B.n344 10.6151
R2040 B.n346 B.n345 10.6151
R2041 B.n346 B.n119 10.6151
R2042 B.n350 B.n119 10.6151
R2043 B.n351 B.n350 10.6151
R2044 B.n352 B.n351 10.6151
R2045 B.n352 B.n117 10.6151
R2046 B.n356 B.n117 10.6151
R2047 B.n357 B.n356 10.6151
R2048 B.n358 B.n357 10.6151
R2049 B.n358 B.n115 10.6151
R2050 B.n362 B.n115 10.6151
R2051 B.n363 B.n362 10.6151
R2052 B.n364 B.n363 10.6151
R2053 B.n364 B.n113 10.6151
R2054 B.n368 B.n113 10.6151
R2055 B.n369 B.n368 10.6151
R2056 B.n370 B.n369 10.6151
R2057 B.n370 B.n111 10.6151
R2058 B.n374 B.n111 10.6151
R2059 B.n375 B.n374 10.6151
R2060 B.n376 B.n375 10.6151
R2061 B.n376 B.n109 10.6151
R2062 B.n380 B.n109 10.6151
R2063 B.n381 B.n380 10.6151
R2064 B.n382 B.n381 10.6151
R2065 B.n382 B.n107 10.6151
R2066 B.n386 B.n107 10.6151
R2067 B.n387 B.n386 10.6151
R2068 B.n388 B.n387 10.6151
R2069 B.n388 B.n105 10.6151
R2070 B.n392 B.n105 10.6151
R2071 B.n393 B.n392 10.6151
R2072 B.n214 B.n213 10.6151
R2073 B.n213 B.n212 10.6151
R2074 B.n212 B.n169 10.6151
R2075 B.n208 B.n169 10.6151
R2076 B.n208 B.n207 10.6151
R2077 B.n207 B.n206 10.6151
R2078 B.n206 B.n171 10.6151
R2079 B.n202 B.n171 10.6151
R2080 B.n202 B.n201 10.6151
R2081 B.n201 B.n200 10.6151
R2082 B.n200 B.n173 10.6151
R2083 B.n196 B.n173 10.6151
R2084 B.n196 B.n195 10.6151
R2085 B.n195 B.n194 10.6151
R2086 B.n194 B.n175 10.6151
R2087 B.n190 B.n175 10.6151
R2088 B.n190 B.n189 10.6151
R2089 B.n189 B.n188 10.6151
R2090 B.n188 B.n177 10.6151
R2091 B.n184 B.n177 10.6151
R2092 B.n184 B.n183 10.6151
R2093 B.n183 B.n182 10.6151
R2094 B.n182 B.n179 10.6151
R2095 B.n179 B.n0 10.6151
R2096 B.n683 B.n1 10.6151
R2097 B.n683 B.n682 10.6151
R2098 B.n682 B.n681 10.6151
R2099 B.n681 B.n4 10.6151
R2100 B.n677 B.n4 10.6151
R2101 B.n677 B.n676 10.6151
R2102 B.n676 B.n675 10.6151
R2103 B.n675 B.n6 10.6151
R2104 B.n671 B.n6 10.6151
R2105 B.n671 B.n670 10.6151
R2106 B.n670 B.n669 10.6151
R2107 B.n669 B.n8 10.6151
R2108 B.n665 B.n8 10.6151
R2109 B.n665 B.n664 10.6151
R2110 B.n664 B.n663 10.6151
R2111 B.n663 B.n10 10.6151
R2112 B.n659 B.n10 10.6151
R2113 B.n659 B.n658 10.6151
R2114 B.n658 B.n657 10.6151
R2115 B.n657 B.n12 10.6151
R2116 B.n653 B.n12 10.6151
R2117 B.n653 B.n652 10.6151
R2118 B.n652 B.n651 10.6151
R2119 B.n651 B.n14 10.6151
R2120 B.n568 B.n567 9.36635
R2121 B.n550 B.n52 9.36635
R2122 B.n297 B.n296 9.36635
R2123 B.n314 B.n133 9.36635
R2124 B.n687 B.n0 2.81026
R2125 B.n687 B.n1 2.81026
R2126 B.n567 B.n566 1.24928
R2127 B.n52 B.n48 1.24928
R2128 B.n298 B.n297 1.24928
R2129 B.n311 B.n133 1.24928
C0 VTAIL VP 3.16358f
C1 VTAIL VDD2 6.2413f
C2 w_n2138_n4220# B 9.992531f
C3 VP VN 6.2396f
C4 VTAIL B 4.60726f
C5 VDD2 VN 3.67671f
C6 VDD1 w_n2138_n4220# 2.07587f
C7 VTAIL VDD1 6.19176f
C8 B VN 1.09446f
C9 VP VDD2 0.332653f
C10 VDD1 VN 0.147783f
C11 VTAIL w_n2138_n4220# 3.34984f
C12 VP B 1.54213f
C13 VDD2 B 2.07066f
C14 w_n2138_n4220# VN 3.03001f
C15 VDD1 VP 3.85829f
C16 VDD1 VDD2 0.673901f
C17 VTAIL VN 3.14923f
C18 VP w_n2138_n4220# 3.30233f
C19 VDD1 B 2.04066f
C20 w_n2138_n4220# VDD2 2.10163f
C21 VDD2 VSUBS 1.072472f
C22 VDD1 VSUBS 5.38152f
C23 VTAIL VSUBS 1.167839f
C24 VN VSUBS 8.646471f
C25 VP VSUBS 1.833626f
C26 B VSUBS 4.263251f
C27 w_n2138_n4220# VSUBS 0.1105p
C28 B.n0 VSUBS 0.004492f
C29 B.n1 VSUBS 0.004492f
C30 B.n2 VSUBS 0.007103f
C31 B.n3 VSUBS 0.007103f
C32 B.n4 VSUBS 0.007103f
C33 B.n5 VSUBS 0.007103f
C34 B.n6 VSUBS 0.007103f
C35 B.n7 VSUBS 0.007103f
C36 B.n8 VSUBS 0.007103f
C37 B.n9 VSUBS 0.007103f
C38 B.n10 VSUBS 0.007103f
C39 B.n11 VSUBS 0.007103f
C40 B.n12 VSUBS 0.007103f
C41 B.n13 VSUBS 0.007103f
C42 B.n14 VSUBS 0.016734f
C43 B.n15 VSUBS 0.007103f
C44 B.n16 VSUBS 0.007103f
C45 B.n17 VSUBS 0.007103f
C46 B.n18 VSUBS 0.007103f
C47 B.n19 VSUBS 0.007103f
C48 B.n20 VSUBS 0.007103f
C49 B.n21 VSUBS 0.007103f
C50 B.n22 VSUBS 0.007103f
C51 B.n23 VSUBS 0.007103f
C52 B.n24 VSUBS 0.007103f
C53 B.n25 VSUBS 0.007103f
C54 B.n26 VSUBS 0.007103f
C55 B.n27 VSUBS 0.007103f
C56 B.n28 VSUBS 0.007103f
C57 B.n29 VSUBS 0.007103f
C58 B.n30 VSUBS 0.007103f
C59 B.n31 VSUBS 0.007103f
C60 B.n32 VSUBS 0.007103f
C61 B.n33 VSUBS 0.007103f
C62 B.n34 VSUBS 0.007103f
C63 B.n35 VSUBS 0.007103f
C64 B.n36 VSUBS 0.007103f
C65 B.n37 VSUBS 0.007103f
C66 B.n38 VSUBS 0.007103f
C67 B.n39 VSUBS 0.007103f
C68 B.n40 VSUBS 0.007103f
C69 B.n41 VSUBS 0.007103f
C70 B.t2 VSUBS 0.314055f
C71 B.t1 VSUBS 0.347614f
C72 B.t0 VSUBS 1.90803f
C73 B.n42 VSUBS 0.536032f
C74 B.n43 VSUBS 0.311847f
C75 B.n44 VSUBS 0.007103f
C76 B.n45 VSUBS 0.007103f
C77 B.n46 VSUBS 0.007103f
C78 B.n47 VSUBS 0.007103f
C79 B.n48 VSUBS 0.003969f
C80 B.n49 VSUBS 0.007103f
C81 B.t8 VSUBS 0.314058f
C82 B.t7 VSUBS 0.347617f
C83 B.t6 VSUBS 1.90803f
C84 B.n50 VSUBS 0.536029f
C85 B.n51 VSUBS 0.311843f
C86 B.n52 VSUBS 0.016457f
C87 B.n53 VSUBS 0.007103f
C88 B.n54 VSUBS 0.007103f
C89 B.n55 VSUBS 0.007103f
C90 B.n56 VSUBS 0.007103f
C91 B.n57 VSUBS 0.007103f
C92 B.n58 VSUBS 0.007103f
C93 B.n59 VSUBS 0.007103f
C94 B.n60 VSUBS 0.007103f
C95 B.n61 VSUBS 0.007103f
C96 B.n62 VSUBS 0.007103f
C97 B.n63 VSUBS 0.007103f
C98 B.n64 VSUBS 0.007103f
C99 B.n65 VSUBS 0.007103f
C100 B.n66 VSUBS 0.007103f
C101 B.n67 VSUBS 0.007103f
C102 B.n68 VSUBS 0.007103f
C103 B.n69 VSUBS 0.007103f
C104 B.n70 VSUBS 0.007103f
C105 B.n71 VSUBS 0.007103f
C106 B.n72 VSUBS 0.007103f
C107 B.n73 VSUBS 0.007103f
C108 B.n74 VSUBS 0.007103f
C109 B.n75 VSUBS 0.007103f
C110 B.n76 VSUBS 0.007103f
C111 B.n77 VSUBS 0.007103f
C112 B.n78 VSUBS 0.017944f
C113 B.n79 VSUBS 0.007103f
C114 B.n80 VSUBS 0.007103f
C115 B.n81 VSUBS 0.007103f
C116 B.n82 VSUBS 0.007103f
C117 B.n83 VSUBS 0.007103f
C118 B.n84 VSUBS 0.007103f
C119 B.n85 VSUBS 0.007103f
C120 B.n86 VSUBS 0.007103f
C121 B.n87 VSUBS 0.007103f
C122 B.n88 VSUBS 0.007103f
C123 B.n89 VSUBS 0.007103f
C124 B.n90 VSUBS 0.007103f
C125 B.n91 VSUBS 0.007103f
C126 B.n92 VSUBS 0.007103f
C127 B.n93 VSUBS 0.007103f
C128 B.n94 VSUBS 0.007103f
C129 B.n95 VSUBS 0.007103f
C130 B.n96 VSUBS 0.007103f
C131 B.n97 VSUBS 0.007103f
C132 B.n98 VSUBS 0.007103f
C133 B.n99 VSUBS 0.007103f
C134 B.n100 VSUBS 0.007103f
C135 B.n101 VSUBS 0.007103f
C136 B.n102 VSUBS 0.007103f
C137 B.n103 VSUBS 0.007103f
C138 B.n104 VSUBS 0.017944f
C139 B.n105 VSUBS 0.007103f
C140 B.n106 VSUBS 0.007103f
C141 B.n107 VSUBS 0.007103f
C142 B.n108 VSUBS 0.007103f
C143 B.n109 VSUBS 0.007103f
C144 B.n110 VSUBS 0.007103f
C145 B.n111 VSUBS 0.007103f
C146 B.n112 VSUBS 0.007103f
C147 B.n113 VSUBS 0.007103f
C148 B.n114 VSUBS 0.007103f
C149 B.n115 VSUBS 0.007103f
C150 B.n116 VSUBS 0.007103f
C151 B.n117 VSUBS 0.007103f
C152 B.n118 VSUBS 0.007103f
C153 B.n119 VSUBS 0.007103f
C154 B.n120 VSUBS 0.007103f
C155 B.n121 VSUBS 0.007103f
C156 B.n122 VSUBS 0.007103f
C157 B.n123 VSUBS 0.007103f
C158 B.n124 VSUBS 0.007103f
C159 B.n125 VSUBS 0.007103f
C160 B.n126 VSUBS 0.007103f
C161 B.n127 VSUBS 0.007103f
C162 B.n128 VSUBS 0.007103f
C163 B.n129 VSUBS 0.007103f
C164 B.n130 VSUBS 0.007103f
C165 B.t4 VSUBS 0.314058f
C166 B.t5 VSUBS 0.347617f
C167 B.t3 VSUBS 1.90803f
C168 B.n131 VSUBS 0.536029f
C169 B.n132 VSUBS 0.311843f
C170 B.n133 VSUBS 0.016457f
C171 B.n134 VSUBS 0.007103f
C172 B.n135 VSUBS 0.007103f
C173 B.n136 VSUBS 0.007103f
C174 B.n137 VSUBS 0.007103f
C175 B.n138 VSUBS 0.007103f
C176 B.t10 VSUBS 0.314055f
C177 B.t11 VSUBS 0.347614f
C178 B.t9 VSUBS 1.90803f
C179 B.n139 VSUBS 0.536032f
C180 B.n140 VSUBS 0.311847f
C181 B.n141 VSUBS 0.007103f
C182 B.n142 VSUBS 0.007103f
C183 B.n143 VSUBS 0.007103f
C184 B.n144 VSUBS 0.007103f
C185 B.n145 VSUBS 0.007103f
C186 B.n146 VSUBS 0.007103f
C187 B.n147 VSUBS 0.007103f
C188 B.n148 VSUBS 0.007103f
C189 B.n149 VSUBS 0.007103f
C190 B.n150 VSUBS 0.007103f
C191 B.n151 VSUBS 0.007103f
C192 B.n152 VSUBS 0.007103f
C193 B.n153 VSUBS 0.007103f
C194 B.n154 VSUBS 0.007103f
C195 B.n155 VSUBS 0.007103f
C196 B.n156 VSUBS 0.007103f
C197 B.n157 VSUBS 0.007103f
C198 B.n158 VSUBS 0.007103f
C199 B.n159 VSUBS 0.007103f
C200 B.n160 VSUBS 0.007103f
C201 B.n161 VSUBS 0.007103f
C202 B.n162 VSUBS 0.007103f
C203 B.n163 VSUBS 0.007103f
C204 B.n164 VSUBS 0.007103f
C205 B.n165 VSUBS 0.007103f
C206 B.n166 VSUBS 0.007103f
C207 B.n167 VSUBS 0.017944f
C208 B.n168 VSUBS 0.007103f
C209 B.n169 VSUBS 0.007103f
C210 B.n170 VSUBS 0.007103f
C211 B.n171 VSUBS 0.007103f
C212 B.n172 VSUBS 0.007103f
C213 B.n173 VSUBS 0.007103f
C214 B.n174 VSUBS 0.007103f
C215 B.n175 VSUBS 0.007103f
C216 B.n176 VSUBS 0.007103f
C217 B.n177 VSUBS 0.007103f
C218 B.n178 VSUBS 0.007103f
C219 B.n179 VSUBS 0.007103f
C220 B.n180 VSUBS 0.007103f
C221 B.n181 VSUBS 0.007103f
C222 B.n182 VSUBS 0.007103f
C223 B.n183 VSUBS 0.007103f
C224 B.n184 VSUBS 0.007103f
C225 B.n185 VSUBS 0.007103f
C226 B.n186 VSUBS 0.007103f
C227 B.n187 VSUBS 0.007103f
C228 B.n188 VSUBS 0.007103f
C229 B.n189 VSUBS 0.007103f
C230 B.n190 VSUBS 0.007103f
C231 B.n191 VSUBS 0.007103f
C232 B.n192 VSUBS 0.007103f
C233 B.n193 VSUBS 0.007103f
C234 B.n194 VSUBS 0.007103f
C235 B.n195 VSUBS 0.007103f
C236 B.n196 VSUBS 0.007103f
C237 B.n197 VSUBS 0.007103f
C238 B.n198 VSUBS 0.007103f
C239 B.n199 VSUBS 0.007103f
C240 B.n200 VSUBS 0.007103f
C241 B.n201 VSUBS 0.007103f
C242 B.n202 VSUBS 0.007103f
C243 B.n203 VSUBS 0.007103f
C244 B.n204 VSUBS 0.007103f
C245 B.n205 VSUBS 0.007103f
C246 B.n206 VSUBS 0.007103f
C247 B.n207 VSUBS 0.007103f
C248 B.n208 VSUBS 0.007103f
C249 B.n209 VSUBS 0.007103f
C250 B.n210 VSUBS 0.007103f
C251 B.n211 VSUBS 0.007103f
C252 B.n212 VSUBS 0.007103f
C253 B.n213 VSUBS 0.007103f
C254 B.n214 VSUBS 0.016734f
C255 B.n215 VSUBS 0.016734f
C256 B.n216 VSUBS 0.017944f
C257 B.n217 VSUBS 0.007103f
C258 B.n218 VSUBS 0.007103f
C259 B.n219 VSUBS 0.007103f
C260 B.n220 VSUBS 0.007103f
C261 B.n221 VSUBS 0.007103f
C262 B.n222 VSUBS 0.007103f
C263 B.n223 VSUBS 0.007103f
C264 B.n224 VSUBS 0.007103f
C265 B.n225 VSUBS 0.007103f
C266 B.n226 VSUBS 0.007103f
C267 B.n227 VSUBS 0.007103f
C268 B.n228 VSUBS 0.007103f
C269 B.n229 VSUBS 0.007103f
C270 B.n230 VSUBS 0.007103f
C271 B.n231 VSUBS 0.007103f
C272 B.n232 VSUBS 0.007103f
C273 B.n233 VSUBS 0.007103f
C274 B.n234 VSUBS 0.007103f
C275 B.n235 VSUBS 0.007103f
C276 B.n236 VSUBS 0.007103f
C277 B.n237 VSUBS 0.007103f
C278 B.n238 VSUBS 0.007103f
C279 B.n239 VSUBS 0.007103f
C280 B.n240 VSUBS 0.007103f
C281 B.n241 VSUBS 0.007103f
C282 B.n242 VSUBS 0.007103f
C283 B.n243 VSUBS 0.007103f
C284 B.n244 VSUBS 0.007103f
C285 B.n245 VSUBS 0.007103f
C286 B.n246 VSUBS 0.007103f
C287 B.n247 VSUBS 0.007103f
C288 B.n248 VSUBS 0.007103f
C289 B.n249 VSUBS 0.007103f
C290 B.n250 VSUBS 0.007103f
C291 B.n251 VSUBS 0.007103f
C292 B.n252 VSUBS 0.007103f
C293 B.n253 VSUBS 0.007103f
C294 B.n254 VSUBS 0.007103f
C295 B.n255 VSUBS 0.007103f
C296 B.n256 VSUBS 0.007103f
C297 B.n257 VSUBS 0.007103f
C298 B.n258 VSUBS 0.007103f
C299 B.n259 VSUBS 0.007103f
C300 B.n260 VSUBS 0.007103f
C301 B.n261 VSUBS 0.007103f
C302 B.n262 VSUBS 0.007103f
C303 B.n263 VSUBS 0.007103f
C304 B.n264 VSUBS 0.007103f
C305 B.n265 VSUBS 0.007103f
C306 B.n266 VSUBS 0.007103f
C307 B.n267 VSUBS 0.007103f
C308 B.n268 VSUBS 0.007103f
C309 B.n269 VSUBS 0.007103f
C310 B.n270 VSUBS 0.007103f
C311 B.n271 VSUBS 0.007103f
C312 B.n272 VSUBS 0.007103f
C313 B.n273 VSUBS 0.007103f
C314 B.n274 VSUBS 0.007103f
C315 B.n275 VSUBS 0.007103f
C316 B.n276 VSUBS 0.007103f
C317 B.n277 VSUBS 0.007103f
C318 B.n278 VSUBS 0.007103f
C319 B.n279 VSUBS 0.007103f
C320 B.n280 VSUBS 0.007103f
C321 B.n281 VSUBS 0.007103f
C322 B.n282 VSUBS 0.007103f
C323 B.n283 VSUBS 0.007103f
C324 B.n284 VSUBS 0.007103f
C325 B.n285 VSUBS 0.007103f
C326 B.n286 VSUBS 0.007103f
C327 B.n287 VSUBS 0.007103f
C328 B.n288 VSUBS 0.007103f
C329 B.n289 VSUBS 0.007103f
C330 B.n290 VSUBS 0.007103f
C331 B.n291 VSUBS 0.007103f
C332 B.n292 VSUBS 0.007103f
C333 B.n293 VSUBS 0.007103f
C334 B.n294 VSUBS 0.007103f
C335 B.n295 VSUBS 0.007103f
C336 B.n296 VSUBS 0.006685f
C337 B.n297 VSUBS 0.016457f
C338 B.n298 VSUBS 0.003969f
C339 B.n299 VSUBS 0.007103f
C340 B.n300 VSUBS 0.007103f
C341 B.n301 VSUBS 0.007103f
C342 B.n302 VSUBS 0.007103f
C343 B.n303 VSUBS 0.007103f
C344 B.n304 VSUBS 0.007103f
C345 B.n305 VSUBS 0.007103f
C346 B.n306 VSUBS 0.007103f
C347 B.n307 VSUBS 0.007103f
C348 B.n308 VSUBS 0.007103f
C349 B.n309 VSUBS 0.007103f
C350 B.n310 VSUBS 0.007103f
C351 B.n311 VSUBS 0.003969f
C352 B.n312 VSUBS 0.007103f
C353 B.n313 VSUBS 0.007103f
C354 B.n314 VSUBS 0.006685f
C355 B.n315 VSUBS 0.007103f
C356 B.n316 VSUBS 0.007103f
C357 B.n317 VSUBS 0.007103f
C358 B.n318 VSUBS 0.007103f
C359 B.n319 VSUBS 0.007103f
C360 B.n320 VSUBS 0.007103f
C361 B.n321 VSUBS 0.007103f
C362 B.n322 VSUBS 0.007103f
C363 B.n323 VSUBS 0.007103f
C364 B.n324 VSUBS 0.007103f
C365 B.n325 VSUBS 0.007103f
C366 B.n326 VSUBS 0.007103f
C367 B.n327 VSUBS 0.007103f
C368 B.n328 VSUBS 0.007103f
C369 B.n329 VSUBS 0.007103f
C370 B.n330 VSUBS 0.007103f
C371 B.n331 VSUBS 0.007103f
C372 B.n332 VSUBS 0.007103f
C373 B.n333 VSUBS 0.007103f
C374 B.n334 VSUBS 0.007103f
C375 B.n335 VSUBS 0.007103f
C376 B.n336 VSUBS 0.007103f
C377 B.n337 VSUBS 0.007103f
C378 B.n338 VSUBS 0.007103f
C379 B.n339 VSUBS 0.007103f
C380 B.n340 VSUBS 0.007103f
C381 B.n341 VSUBS 0.007103f
C382 B.n342 VSUBS 0.007103f
C383 B.n343 VSUBS 0.007103f
C384 B.n344 VSUBS 0.007103f
C385 B.n345 VSUBS 0.007103f
C386 B.n346 VSUBS 0.007103f
C387 B.n347 VSUBS 0.007103f
C388 B.n348 VSUBS 0.007103f
C389 B.n349 VSUBS 0.007103f
C390 B.n350 VSUBS 0.007103f
C391 B.n351 VSUBS 0.007103f
C392 B.n352 VSUBS 0.007103f
C393 B.n353 VSUBS 0.007103f
C394 B.n354 VSUBS 0.007103f
C395 B.n355 VSUBS 0.007103f
C396 B.n356 VSUBS 0.007103f
C397 B.n357 VSUBS 0.007103f
C398 B.n358 VSUBS 0.007103f
C399 B.n359 VSUBS 0.007103f
C400 B.n360 VSUBS 0.007103f
C401 B.n361 VSUBS 0.007103f
C402 B.n362 VSUBS 0.007103f
C403 B.n363 VSUBS 0.007103f
C404 B.n364 VSUBS 0.007103f
C405 B.n365 VSUBS 0.007103f
C406 B.n366 VSUBS 0.007103f
C407 B.n367 VSUBS 0.007103f
C408 B.n368 VSUBS 0.007103f
C409 B.n369 VSUBS 0.007103f
C410 B.n370 VSUBS 0.007103f
C411 B.n371 VSUBS 0.007103f
C412 B.n372 VSUBS 0.007103f
C413 B.n373 VSUBS 0.007103f
C414 B.n374 VSUBS 0.007103f
C415 B.n375 VSUBS 0.007103f
C416 B.n376 VSUBS 0.007103f
C417 B.n377 VSUBS 0.007103f
C418 B.n378 VSUBS 0.007103f
C419 B.n379 VSUBS 0.007103f
C420 B.n380 VSUBS 0.007103f
C421 B.n381 VSUBS 0.007103f
C422 B.n382 VSUBS 0.007103f
C423 B.n383 VSUBS 0.007103f
C424 B.n384 VSUBS 0.007103f
C425 B.n385 VSUBS 0.007103f
C426 B.n386 VSUBS 0.007103f
C427 B.n387 VSUBS 0.007103f
C428 B.n388 VSUBS 0.007103f
C429 B.n389 VSUBS 0.007103f
C430 B.n390 VSUBS 0.007103f
C431 B.n391 VSUBS 0.007103f
C432 B.n392 VSUBS 0.007103f
C433 B.n393 VSUBS 0.017944f
C434 B.n394 VSUBS 0.016734f
C435 B.n395 VSUBS 0.016734f
C436 B.n396 VSUBS 0.007103f
C437 B.n397 VSUBS 0.007103f
C438 B.n398 VSUBS 0.007103f
C439 B.n399 VSUBS 0.007103f
C440 B.n400 VSUBS 0.007103f
C441 B.n401 VSUBS 0.007103f
C442 B.n402 VSUBS 0.007103f
C443 B.n403 VSUBS 0.007103f
C444 B.n404 VSUBS 0.007103f
C445 B.n405 VSUBS 0.007103f
C446 B.n406 VSUBS 0.007103f
C447 B.n407 VSUBS 0.007103f
C448 B.n408 VSUBS 0.007103f
C449 B.n409 VSUBS 0.007103f
C450 B.n410 VSUBS 0.007103f
C451 B.n411 VSUBS 0.007103f
C452 B.n412 VSUBS 0.007103f
C453 B.n413 VSUBS 0.007103f
C454 B.n414 VSUBS 0.007103f
C455 B.n415 VSUBS 0.007103f
C456 B.n416 VSUBS 0.007103f
C457 B.n417 VSUBS 0.007103f
C458 B.n418 VSUBS 0.007103f
C459 B.n419 VSUBS 0.007103f
C460 B.n420 VSUBS 0.007103f
C461 B.n421 VSUBS 0.007103f
C462 B.n422 VSUBS 0.007103f
C463 B.n423 VSUBS 0.007103f
C464 B.n424 VSUBS 0.007103f
C465 B.n425 VSUBS 0.007103f
C466 B.n426 VSUBS 0.007103f
C467 B.n427 VSUBS 0.007103f
C468 B.n428 VSUBS 0.007103f
C469 B.n429 VSUBS 0.007103f
C470 B.n430 VSUBS 0.007103f
C471 B.n431 VSUBS 0.007103f
C472 B.n432 VSUBS 0.007103f
C473 B.n433 VSUBS 0.007103f
C474 B.n434 VSUBS 0.007103f
C475 B.n435 VSUBS 0.007103f
C476 B.n436 VSUBS 0.007103f
C477 B.n437 VSUBS 0.007103f
C478 B.n438 VSUBS 0.007103f
C479 B.n439 VSUBS 0.007103f
C480 B.n440 VSUBS 0.007103f
C481 B.n441 VSUBS 0.007103f
C482 B.n442 VSUBS 0.007103f
C483 B.n443 VSUBS 0.007103f
C484 B.n444 VSUBS 0.007103f
C485 B.n445 VSUBS 0.007103f
C486 B.n446 VSUBS 0.007103f
C487 B.n447 VSUBS 0.007103f
C488 B.n448 VSUBS 0.007103f
C489 B.n449 VSUBS 0.007103f
C490 B.n450 VSUBS 0.007103f
C491 B.n451 VSUBS 0.007103f
C492 B.n452 VSUBS 0.007103f
C493 B.n453 VSUBS 0.007103f
C494 B.n454 VSUBS 0.007103f
C495 B.n455 VSUBS 0.007103f
C496 B.n456 VSUBS 0.007103f
C497 B.n457 VSUBS 0.007103f
C498 B.n458 VSUBS 0.007103f
C499 B.n459 VSUBS 0.007103f
C500 B.n460 VSUBS 0.007103f
C501 B.n461 VSUBS 0.007103f
C502 B.n462 VSUBS 0.007103f
C503 B.n463 VSUBS 0.007103f
C504 B.n464 VSUBS 0.007103f
C505 B.n465 VSUBS 0.007103f
C506 B.n466 VSUBS 0.007103f
C507 B.n467 VSUBS 0.007103f
C508 B.n468 VSUBS 0.007103f
C509 B.n469 VSUBS 0.016734f
C510 B.n470 VSUBS 0.017522f
C511 B.n471 VSUBS 0.017157f
C512 B.n472 VSUBS 0.007103f
C513 B.n473 VSUBS 0.007103f
C514 B.n474 VSUBS 0.007103f
C515 B.n475 VSUBS 0.007103f
C516 B.n476 VSUBS 0.007103f
C517 B.n477 VSUBS 0.007103f
C518 B.n478 VSUBS 0.007103f
C519 B.n479 VSUBS 0.007103f
C520 B.n480 VSUBS 0.007103f
C521 B.n481 VSUBS 0.007103f
C522 B.n482 VSUBS 0.007103f
C523 B.n483 VSUBS 0.007103f
C524 B.n484 VSUBS 0.007103f
C525 B.n485 VSUBS 0.007103f
C526 B.n486 VSUBS 0.007103f
C527 B.n487 VSUBS 0.007103f
C528 B.n488 VSUBS 0.007103f
C529 B.n489 VSUBS 0.007103f
C530 B.n490 VSUBS 0.007103f
C531 B.n491 VSUBS 0.007103f
C532 B.n492 VSUBS 0.007103f
C533 B.n493 VSUBS 0.007103f
C534 B.n494 VSUBS 0.007103f
C535 B.n495 VSUBS 0.007103f
C536 B.n496 VSUBS 0.007103f
C537 B.n497 VSUBS 0.007103f
C538 B.n498 VSUBS 0.007103f
C539 B.n499 VSUBS 0.007103f
C540 B.n500 VSUBS 0.007103f
C541 B.n501 VSUBS 0.007103f
C542 B.n502 VSUBS 0.007103f
C543 B.n503 VSUBS 0.007103f
C544 B.n504 VSUBS 0.007103f
C545 B.n505 VSUBS 0.007103f
C546 B.n506 VSUBS 0.007103f
C547 B.n507 VSUBS 0.007103f
C548 B.n508 VSUBS 0.007103f
C549 B.n509 VSUBS 0.007103f
C550 B.n510 VSUBS 0.007103f
C551 B.n511 VSUBS 0.007103f
C552 B.n512 VSUBS 0.007103f
C553 B.n513 VSUBS 0.007103f
C554 B.n514 VSUBS 0.007103f
C555 B.n515 VSUBS 0.007103f
C556 B.n516 VSUBS 0.007103f
C557 B.n517 VSUBS 0.007103f
C558 B.n518 VSUBS 0.007103f
C559 B.n519 VSUBS 0.007103f
C560 B.n520 VSUBS 0.007103f
C561 B.n521 VSUBS 0.007103f
C562 B.n522 VSUBS 0.007103f
C563 B.n523 VSUBS 0.007103f
C564 B.n524 VSUBS 0.007103f
C565 B.n525 VSUBS 0.007103f
C566 B.n526 VSUBS 0.007103f
C567 B.n527 VSUBS 0.007103f
C568 B.n528 VSUBS 0.007103f
C569 B.n529 VSUBS 0.007103f
C570 B.n530 VSUBS 0.007103f
C571 B.n531 VSUBS 0.007103f
C572 B.n532 VSUBS 0.007103f
C573 B.n533 VSUBS 0.007103f
C574 B.n534 VSUBS 0.007103f
C575 B.n535 VSUBS 0.007103f
C576 B.n536 VSUBS 0.007103f
C577 B.n537 VSUBS 0.007103f
C578 B.n538 VSUBS 0.007103f
C579 B.n539 VSUBS 0.007103f
C580 B.n540 VSUBS 0.007103f
C581 B.n541 VSUBS 0.007103f
C582 B.n542 VSUBS 0.007103f
C583 B.n543 VSUBS 0.007103f
C584 B.n544 VSUBS 0.007103f
C585 B.n545 VSUBS 0.007103f
C586 B.n546 VSUBS 0.007103f
C587 B.n547 VSUBS 0.007103f
C588 B.n548 VSUBS 0.007103f
C589 B.n549 VSUBS 0.007103f
C590 B.n550 VSUBS 0.006685f
C591 B.n551 VSUBS 0.007103f
C592 B.n552 VSUBS 0.007103f
C593 B.n553 VSUBS 0.007103f
C594 B.n554 VSUBS 0.007103f
C595 B.n555 VSUBS 0.007103f
C596 B.n556 VSUBS 0.007103f
C597 B.n557 VSUBS 0.007103f
C598 B.n558 VSUBS 0.007103f
C599 B.n559 VSUBS 0.007103f
C600 B.n560 VSUBS 0.007103f
C601 B.n561 VSUBS 0.007103f
C602 B.n562 VSUBS 0.007103f
C603 B.n563 VSUBS 0.007103f
C604 B.n564 VSUBS 0.007103f
C605 B.n565 VSUBS 0.007103f
C606 B.n566 VSUBS 0.003969f
C607 B.n567 VSUBS 0.016457f
C608 B.n568 VSUBS 0.006685f
C609 B.n569 VSUBS 0.007103f
C610 B.n570 VSUBS 0.007103f
C611 B.n571 VSUBS 0.007103f
C612 B.n572 VSUBS 0.007103f
C613 B.n573 VSUBS 0.007103f
C614 B.n574 VSUBS 0.007103f
C615 B.n575 VSUBS 0.007103f
C616 B.n576 VSUBS 0.007103f
C617 B.n577 VSUBS 0.007103f
C618 B.n578 VSUBS 0.007103f
C619 B.n579 VSUBS 0.007103f
C620 B.n580 VSUBS 0.007103f
C621 B.n581 VSUBS 0.007103f
C622 B.n582 VSUBS 0.007103f
C623 B.n583 VSUBS 0.007103f
C624 B.n584 VSUBS 0.007103f
C625 B.n585 VSUBS 0.007103f
C626 B.n586 VSUBS 0.007103f
C627 B.n587 VSUBS 0.007103f
C628 B.n588 VSUBS 0.007103f
C629 B.n589 VSUBS 0.007103f
C630 B.n590 VSUBS 0.007103f
C631 B.n591 VSUBS 0.007103f
C632 B.n592 VSUBS 0.007103f
C633 B.n593 VSUBS 0.007103f
C634 B.n594 VSUBS 0.007103f
C635 B.n595 VSUBS 0.007103f
C636 B.n596 VSUBS 0.007103f
C637 B.n597 VSUBS 0.007103f
C638 B.n598 VSUBS 0.007103f
C639 B.n599 VSUBS 0.007103f
C640 B.n600 VSUBS 0.007103f
C641 B.n601 VSUBS 0.007103f
C642 B.n602 VSUBS 0.007103f
C643 B.n603 VSUBS 0.007103f
C644 B.n604 VSUBS 0.007103f
C645 B.n605 VSUBS 0.007103f
C646 B.n606 VSUBS 0.007103f
C647 B.n607 VSUBS 0.007103f
C648 B.n608 VSUBS 0.007103f
C649 B.n609 VSUBS 0.007103f
C650 B.n610 VSUBS 0.007103f
C651 B.n611 VSUBS 0.007103f
C652 B.n612 VSUBS 0.007103f
C653 B.n613 VSUBS 0.007103f
C654 B.n614 VSUBS 0.007103f
C655 B.n615 VSUBS 0.007103f
C656 B.n616 VSUBS 0.007103f
C657 B.n617 VSUBS 0.007103f
C658 B.n618 VSUBS 0.007103f
C659 B.n619 VSUBS 0.007103f
C660 B.n620 VSUBS 0.007103f
C661 B.n621 VSUBS 0.007103f
C662 B.n622 VSUBS 0.007103f
C663 B.n623 VSUBS 0.007103f
C664 B.n624 VSUBS 0.007103f
C665 B.n625 VSUBS 0.007103f
C666 B.n626 VSUBS 0.007103f
C667 B.n627 VSUBS 0.007103f
C668 B.n628 VSUBS 0.007103f
C669 B.n629 VSUBS 0.007103f
C670 B.n630 VSUBS 0.007103f
C671 B.n631 VSUBS 0.007103f
C672 B.n632 VSUBS 0.007103f
C673 B.n633 VSUBS 0.007103f
C674 B.n634 VSUBS 0.007103f
C675 B.n635 VSUBS 0.007103f
C676 B.n636 VSUBS 0.007103f
C677 B.n637 VSUBS 0.007103f
C678 B.n638 VSUBS 0.007103f
C679 B.n639 VSUBS 0.007103f
C680 B.n640 VSUBS 0.007103f
C681 B.n641 VSUBS 0.007103f
C682 B.n642 VSUBS 0.007103f
C683 B.n643 VSUBS 0.007103f
C684 B.n644 VSUBS 0.007103f
C685 B.n645 VSUBS 0.007103f
C686 B.n646 VSUBS 0.007103f
C687 B.n647 VSUBS 0.017944f
C688 B.n648 VSUBS 0.017944f
C689 B.n649 VSUBS 0.016734f
C690 B.n650 VSUBS 0.007103f
C691 B.n651 VSUBS 0.007103f
C692 B.n652 VSUBS 0.007103f
C693 B.n653 VSUBS 0.007103f
C694 B.n654 VSUBS 0.007103f
C695 B.n655 VSUBS 0.007103f
C696 B.n656 VSUBS 0.007103f
C697 B.n657 VSUBS 0.007103f
C698 B.n658 VSUBS 0.007103f
C699 B.n659 VSUBS 0.007103f
C700 B.n660 VSUBS 0.007103f
C701 B.n661 VSUBS 0.007103f
C702 B.n662 VSUBS 0.007103f
C703 B.n663 VSUBS 0.007103f
C704 B.n664 VSUBS 0.007103f
C705 B.n665 VSUBS 0.007103f
C706 B.n666 VSUBS 0.007103f
C707 B.n667 VSUBS 0.007103f
C708 B.n668 VSUBS 0.007103f
C709 B.n669 VSUBS 0.007103f
C710 B.n670 VSUBS 0.007103f
C711 B.n671 VSUBS 0.007103f
C712 B.n672 VSUBS 0.007103f
C713 B.n673 VSUBS 0.007103f
C714 B.n674 VSUBS 0.007103f
C715 B.n675 VSUBS 0.007103f
C716 B.n676 VSUBS 0.007103f
C717 B.n677 VSUBS 0.007103f
C718 B.n678 VSUBS 0.007103f
C719 B.n679 VSUBS 0.007103f
C720 B.n680 VSUBS 0.007103f
C721 B.n681 VSUBS 0.007103f
C722 B.n682 VSUBS 0.007103f
C723 B.n683 VSUBS 0.007103f
C724 B.n684 VSUBS 0.007103f
C725 B.n685 VSUBS 0.007103f
C726 B.n686 VSUBS 0.007103f
C727 B.n687 VSUBS 0.016083f
C728 VDD2.n0 VSUBS 0.031853f
C729 VDD2.n1 VSUBS 0.028439f
C730 VDD2.n2 VSUBS 0.015282f
C731 VDD2.n3 VSUBS 0.036121f
C732 VDD2.n4 VSUBS 0.016181f
C733 VDD2.n5 VSUBS 0.028439f
C734 VDD2.n6 VSUBS 0.015731f
C735 VDD2.n7 VSUBS 0.036121f
C736 VDD2.n8 VSUBS 0.016181f
C737 VDD2.n9 VSUBS 0.028439f
C738 VDD2.n10 VSUBS 0.015282f
C739 VDD2.n11 VSUBS 0.036121f
C740 VDD2.n12 VSUBS 0.016181f
C741 VDD2.n13 VSUBS 0.028439f
C742 VDD2.n14 VSUBS 0.015282f
C743 VDD2.n15 VSUBS 0.036121f
C744 VDD2.n16 VSUBS 0.016181f
C745 VDD2.n17 VSUBS 0.028439f
C746 VDD2.n18 VSUBS 0.015282f
C747 VDD2.n19 VSUBS 0.036121f
C748 VDD2.n20 VSUBS 0.016181f
C749 VDD2.n21 VSUBS 0.028439f
C750 VDD2.n22 VSUBS 0.015282f
C751 VDD2.n23 VSUBS 0.036121f
C752 VDD2.n24 VSUBS 0.016181f
C753 VDD2.n25 VSUBS 0.028439f
C754 VDD2.n26 VSUBS 0.015282f
C755 VDD2.n27 VSUBS 0.02709f
C756 VDD2.n28 VSUBS 0.022978f
C757 VDD2.t1 VSUBS 0.077416f
C758 VDD2.n29 VSUBS 0.211039f
C759 VDD2.n30 VSUBS 1.97855f
C760 VDD2.n31 VSUBS 0.015282f
C761 VDD2.n32 VSUBS 0.016181f
C762 VDD2.n33 VSUBS 0.036121f
C763 VDD2.n34 VSUBS 0.036121f
C764 VDD2.n35 VSUBS 0.016181f
C765 VDD2.n36 VSUBS 0.015282f
C766 VDD2.n37 VSUBS 0.028439f
C767 VDD2.n38 VSUBS 0.028439f
C768 VDD2.n39 VSUBS 0.015282f
C769 VDD2.n40 VSUBS 0.016181f
C770 VDD2.n41 VSUBS 0.036121f
C771 VDD2.n42 VSUBS 0.036121f
C772 VDD2.n43 VSUBS 0.016181f
C773 VDD2.n44 VSUBS 0.015282f
C774 VDD2.n45 VSUBS 0.028439f
C775 VDD2.n46 VSUBS 0.028439f
C776 VDD2.n47 VSUBS 0.015282f
C777 VDD2.n48 VSUBS 0.016181f
C778 VDD2.n49 VSUBS 0.036121f
C779 VDD2.n50 VSUBS 0.036121f
C780 VDD2.n51 VSUBS 0.016181f
C781 VDD2.n52 VSUBS 0.015282f
C782 VDD2.n53 VSUBS 0.028439f
C783 VDD2.n54 VSUBS 0.028439f
C784 VDD2.n55 VSUBS 0.015282f
C785 VDD2.n56 VSUBS 0.016181f
C786 VDD2.n57 VSUBS 0.036121f
C787 VDD2.n58 VSUBS 0.036121f
C788 VDD2.n59 VSUBS 0.016181f
C789 VDD2.n60 VSUBS 0.015282f
C790 VDD2.n61 VSUBS 0.028439f
C791 VDD2.n62 VSUBS 0.028439f
C792 VDD2.n63 VSUBS 0.015282f
C793 VDD2.n64 VSUBS 0.016181f
C794 VDD2.n65 VSUBS 0.036121f
C795 VDD2.n66 VSUBS 0.036121f
C796 VDD2.n67 VSUBS 0.016181f
C797 VDD2.n68 VSUBS 0.015282f
C798 VDD2.n69 VSUBS 0.028439f
C799 VDD2.n70 VSUBS 0.028439f
C800 VDD2.n71 VSUBS 0.015282f
C801 VDD2.n72 VSUBS 0.015282f
C802 VDD2.n73 VSUBS 0.016181f
C803 VDD2.n74 VSUBS 0.036121f
C804 VDD2.n75 VSUBS 0.036121f
C805 VDD2.n76 VSUBS 0.036121f
C806 VDD2.n77 VSUBS 0.015731f
C807 VDD2.n78 VSUBS 0.015282f
C808 VDD2.n79 VSUBS 0.028439f
C809 VDD2.n80 VSUBS 0.028439f
C810 VDD2.n81 VSUBS 0.015282f
C811 VDD2.n82 VSUBS 0.016181f
C812 VDD2.n83 VSUBS 0.036121f
C813 VDD2.n84 VSUBS 0.089503f
C814 VDD2.n85 VSUBS 0.016181f
C815 VDD2.n86 VSUBS 0.015282f
C816 VDD2.n87 VSUBS 0.072728f
C817 VDD2.n88 VSUBS 0.98218f
C818 VDD2.n89 VSUBS 0.031853f
C819 VDD2.n90 VSUBS 0.028439f
C820 VDD2.n91 VSUBS 0.015282f
C821 VDD2.n92 VSUBS 0.036121f
C822 VDD2.n93 VSUBS 0.016181f
C823 VDD2.n94 VSUBS 0.028439f
C824 VDD2.n95 VSUBS 0.015731f
C825 VDD2.n96 VSUBS 0.036121f
C826 VDD2.n97 VSUBS 0.015282f
C827 VDD2.n98 VSUBS 0.016181f
C828 VDD2.n99 VSUBS 0.028439f
C829 VDD2.n100 VSUBS 0.015282f
C830 VDD2.n101 VSUBS 0.036121f
C831 VDD2.n102 VSUBS 0.016181f
C832 VDD2.n103 VSUBS 0.028439f
C833 VDD2.n104 VSUBS 0.015282f
C834 VDD2.n105 VSUBS 0.036121f
C835 VDD2.n106 VSUBS 0.016181f
C836 VDD2.n107 VSUBS 0.028439f
C837 VDD2.n108 VSUBS 0.015282f
C838 VDD2.n109 VSUBS 0.036121f
C839 VDD2.n110 VSUBS 0.016181f
C840 VDD2.n111 VSUBS 0.028439f
C841 VDD2.n112 VSUBS 0.015282f
C842 VDD2.n113 VSUBS 0.036121f
C843 VDD2.n114 VSUBS 0.016181f
C844 VDD2.n115 VSUBS 0.028439f
C845 VDD2.n116 VSUBS 0.015282f
C846 VDD2.n117 VSUBS 0.02709f
C847 VDD2.n118 VSUBS 0.022978f
C848 VDD2.t0 VSUBS 0.077416f
C849 VDD2.n119 VSUBS 0.211039f
C850 VDD2.n120 VSUBS 1.97855f
C851 VDD2.n121 VSUBS 0.015282f
C852 VDD2.n122 VSUBS 0.016181f
C853 VDD2.n123 VSUBS 0.036121f
C854 VDD2.n124 VSUBS 0.036121f
C855 VDD2.n125 VSUBS 0.016181f
C856 VDD2.n126 VSUBS 0.015282f
C857 VDD2.n127 VSUBS 0.028439f
C858 VDD2.n128 VSUBS 0.028439f
C859 VDD2.n129 VSUBS 0.015282f
C860 VDD2.n130 VSUBS 0.016181f
C861 VDD2.n131 VSUBS 0.036121f
C862 VDD2.n132 VSUBS 0.036121f
C863 VDD2.n133 VSUBS 0.016181f
C864 VDD2.n134 VSUBS 0.015282f
C865 VDD2.n135 VSUBS 0.028439f
C866 VDD2.n136 VSUBS 0.028439f
C867 VDD2.n137 VSUBS 0.015282f
C868 VDD2.n138 VSUBS 0.016181f
C869 VDD2.n139 VSUBS 0.036121f
C870 VDD2.n140 VSUBS 0.036121f
C871 VDD2.n141 VSUBS 0.016181f
C872 VDD2.n142 VSUBS 0.015282f
C873 VDD2.n143 VSUBS 0.028439f
C874 VDD2.n144 VSUBS 0.028439f
C875 VDD2.n145 VSUBS 0.015282f
C876 VDD2.n146 VSUBS 0.016181f
C877 VDD2.n147 VSUBS 0.036121f
C878 VDD2.n148 VSUBS 0.036121f
C879 VDD2.n149 VSUBS 0.016181f
C880 VDD2.n150 VSUBS 0.015282f
C881 VDD2.n151 VSUBS 0.028439f
C882 VDD2.n152 VSUBS 0.028439f
C883 VDD2.n153 VSUBS 0.015282f
C884 VDD2.n154 VSUBS 0.016181f
C885 VDD2.n155 VSUBS 0.036121f
C886 VDD2.n156 VSUBS 0.036121f
C887 VDD2.n157 VSUBS 0.016181f
C888 VDD2.n158 VSUBS 0.015282f
C889 VDD2.n159 VSUBS 0.028439f
C890 VDD2.n160 VSUBS 0.028439f
C891 VDD2.n161 VSUBS 0.015282f
C892 VDD2.n162 VSUBS 0.016181f
C893 VDD2.n163 VSUBS 0.036121f
C894 VDD2.n164 VSUBS 0.036121f
C895 VDD2.n165 VSUBS 0.036121f
C896 VDD2.n166 VSUBS 0.015731f
C897 VDD2.n167 VSUBS 0.015282f
C898 VDD2.n168 VSUBS 0.028439f
C899 VDD2.n169 VSUBS 0.028439f
C900 VDD2.n170 VSUBS 0.015282f
C901 VDD2.n171 VSUBS 0.016181f
C902 VDD2.n172 VSUBS 0.036121f
C903 VDD2.n173 VSUBS 0.089503f
C904 VDD2.n174 VSUBS 0.016181f
C905 VDD2.n175 VSUBS 0.015282f
C906 VDD2.n176 VSUBS 0.072728f
C907 VDD2.n177 VSUBS 0.064894f
C908 VDD2.n178 VSUBS 4.00635f
C909 VN.t0 VSUBS 4.64849f
C910 VN.t1 VSUBS 5.28838f
C911 VDD1.n0 VSUBS 0.031841f
C912 VDD1.n1 VSUBS 0.028429f
C913 VDD1.n2 VSUBS 0.015276f
C914 VDD1.n3 VSUBS 0.036108f
C915 VDD1.n4 VSUBS 0.016175f
C916 VDD1.n5 VSUBS 0.028429f
C917 VDD1.n6 VSUBS 0.015726f
C918 VDD1.n7 VSUBS 0.036108f
C919 VDD1.n8 VSUBS 0.015276f
C920 VDD1.n9 VSUBS 0.016175f
C921 VDD1.n10 VSUBS 0.028429f
C922 VDD1.n11 VSUBS 0.015276f
C923 VDD1.n12 VSUBS 0.036108f
C924 VDD1.n13 VSUBS 0.016175f
C925 VDD1.n14 VSUBS 0.028429f
C926 VDD1.n15 VSUBS 0.015276f
C927 VDD1.n16 VSUBS 0.036108f
C928 VDD1.n17 VSUBS 0.016175f
C929 VDD1.n18 VSUBS 0.028429f
C930 VDD1.n19 VSUBS 0.015276f
C931 VDD1.n20 VSUBS 0.036108f
C932 VDD1.n21 VSUBS 0.016175f
C933 VDD1.n22 VSUBS 0.028429f
C934 VDD1.n23 VSUBS 0.015276f
C935 VDD1.n24 VSUBS 0.036108f
C936 VDD1.n25 VSUBS 0.016175f
C937 VDD1.n26 VSUBS 0.028429f
C938 VDD1.n27 VSUBS 0.015276f
C939 VDD1.n28 VSUBS 0.027081f
C940 VDD1.n29 VSUBS 0.02297f
C941 VDD1.t0 VSUBS 0.077389f
C942 VDD1.n30 VSUBS 0.210964f
C943 VDD1.n31 VSUBS 1.97785f
C944 VDD1.n32 VSUBS 0.015276f
C945 VDD1.n33 VSUBS 0.016175f
C946 VDD1.n34 VSUBS 0.036108f
C947 VDD1.n35 VSUBS 0.036108f
C948 VDD1.n36 VSUBS 0.016175f
C949 VDD1.n37 VSUBS 0.015276f
C950 VDD1.n38 VSUBS 0.028429f
C951 VDD1.n39 VSUBS 0.028429f
C952 VDD1.n40 VSUBS 0.015276f
C953 VDD1.n41 VSUBS 0.016175f
C954 VDD1.n42 VSUBS 0.036108f
C955 VDD1.n43 VSUBS 0.036108f
C956 VDD1.n44 VSUBS 0.016175f
C957 VDD1.n45 VSUBS 0.015276f
C958 VDD1.n46 VSUBS 0.028429f
C959 VDD1.n47 VSUBS 0.028429f
C960 VDD1.n48 VSUBS 0.015276f
C961 VDD1.n49 VSUBS 0.016175f
C962 VDD1.n50 VSUBS 0.036108f
C963 VDD1.n51 VSUBS 0.036108f
C964 VDD1.n52 VSUBS 0.016175f
C965 VDD1.n53 VSUBS 0.015276f
C966 VDD1.n54 VSUBS 0.028429f
C967 VDD1.n55 VSUBS 0.028429f
C968 VDD1.n56 VSUBS 0.015276f
C969 VDD1.n57 VSUBS 0.016175f
C970 VDD1.n58 VSUBS 0.036108f
C971 VDD1.n59 VSUBS 0.036108f
C972 VDD1.n60 VSUBS 0.016175f
C973 VDD1.n61 VSUBS 0.015276f
C974 VDD1.n62 VSUBS 0.028429f
C975 VDD1.n63 VSUBS 0.028429f
C976 VDD1.n64 VSUBS 0.015276f
C977 VDD1.n65 VSUBS 0.016175f
C978 VDD1.n66 VSUBS 0.036108f
C979 VDD1.n67 VSUBS 0.036108f
C980 VDD1.n68 VSUBS 0.016175f
C981 VDD1.n69 VSUBS 0.015276f
C982 VDD1.n70 VSUBS 0.028429f
C983 VDD1.n71 VSUBS 0.028429f
C984 VDD1.n72 VSUBS 0.015276f
C985 VDD1.n73 VSUBS 0.016175f
C986 VDD1.n74 VSUBS 0.036108f
C987 VDD1.n75 VSUBS 0.036108f
C988 VDD1.n76 VSUBS 0.036108f
C989 VDD1.n77 VSUBS 0.015726f
C990 VDD1.n78 VSUBS 0.015276f
C991 VDD1.n79 VSUBS 0.028429f
C992 VDD1.n80 VSUBS 0.028429f
C993 VDD1.n81 VSUBS 0.015276f
C994 VDD1.n82 VSUBS 0.016175f
C995 VDD1.n83 VSUBS 0.036108f
C996 VDD1.n84 VSUBS 0.089471f
C997 VDD1.n85 VSUBS 0.016175f
C998 VDD1.n86 VSUBS 0.015276f
C999 VDD1.n87 VSUBS 0.072702f
C1000 VDD1.n88 VSUBS 0.066449f
C1001 VDD1.n89 VSUBS 0.031841f
C1002 VDD1.n90 VSUBS 0.028429f
C1003 VDD1.n91 VSUBS 0.015276f
C1004 VDD1.n92 VSUBS 0.036108f
C1005 VDD1.n93 VSUBS 0.016175f
C1006 VDD1.n94 VSUBS 0.028429f
C1007 VDD1.n95 VSUBS 0.015726f
C1008 VDD1.n96 VSUBS 0.036108f
C1009 VDD1.n97 VSUBS 0.016175f
C1010 VDD1.n98 VSUBS 0.028429f
C1011 VDD1.n99 VSUBS 0.015276f
C1012 VDD1.n100 VSUBS 0.036108f
C1013 VDD1.n101 VSUBS 0.016175f
C1014 VDD1.n102 VSUBS 0.028429f
C1015 VDD1.n103 VSUBS 0.015276f
C1016 VDD1.n104 VSUBS 0.036108f
C1017 VDD1.n105 VSUBS 0.016175f
C1018 VDD1.n106 VSUBS 0.028429f
C1019 VDD1.n107 VSUBS 0.015276f
C1020 VDD1.n108 VSUBS 0.036108f
C1021 VDD1.n109 VSUBS 0.016175f
C1022 VDD1.n110 VSUBS 0.028429f
C1023 VDD1.n111 VSUBS 0.015276f
C1024 VDD1.n112 VSUBS 0.036108f
C1025 VDD1.n113 VSUBS 0.016175f
C1026 VDD1.n114 VSUBS 0.028429f
C1027 VDD1.n115 VSUBS 0.015276f
C1028 VDD1.n116 VSUBS 0.027081f
C1029 VDD1.n117 VSUBS 0.02297f
C1030 VDD1.t1 VSUBS 0.077389f
C1031 VDD1.n118 VSUBS 0.210964f
C1032 VDD1.n119 VSUBS 1.97785f
C1033 VDD1.n120 VSUBS 0.015276f
C1034 VDD1.n121 VSUBS 0.016175f
C1035 VDD1.n122 VSUBS 0.036108f
C1036 VDD1.n123 VSUBS 0.036108f
C1037 VDD1.n124 VSUBS 0.016175f
C1038 VDD1.n125 VSUBS 0.015276f
C1039 VDD1.n126 VSUBS 0.028429f
C1040 VDD1.n127 VSUBS 0.028429f
C1041 VDD1.n128 VSUBS 0.015276f
C1042 VDD1.n129 VSUBS 0.016175f
C1043 VDD1.n130 VSUBS 0.036108f
C1044 VDD1.n131 VSUBS 0.036108f
C1045 VDD1.n132 VSUBS 0.016175f
C1046 VDD1.n133 VSUBS 0.015276f
C1047 VDD1.n134 VSUBS 0.028429f
C1048 VDD1.n135 VSUBS 0.028429f
C1049 VDD1.n136 VSUBS 0.015276f
C1050 VDD1.n137 VSUBS 0.016175f
C1051 VDD1.n138 VSUBS 0.036108f
C1052 VDD1.n139 VSUBS 0.036108f
C1053 VDD1.n140 VSUBS 0.016175f
C1054 VDD1.n141 VSUBS 0.015276f
C1055 VDD1.n142 VSUBS 0.028429f
C1056 VDD1.n143 VSUBS 0.028429f
C1057 VDD1.n144 VSUBS 0.015276f
C1058 VDD1.n145 VSUBS 0.016175f
C1059 VDD1.n146 VSUBS 0.036108f
C1060 VDD1.n147 VSUBS 0.036108f
C1061 VDD1.n148 VSUBS 0.016175f
C1062 VDD1.n149 VSUBS 0.015276f
C1063 VDD1.n150 VSUBS 0.028429f
C1064 VDD1.n151 VSUBS 0.028429f
C1065 VDD1.n152 VSUBS 0.015276f
C1066 VDD1.n153 VSUBS 0.016175f
C1067 VDD1.n154 VSUBS 0.036108f
C1068 VDD1.n155 VSUBS 0.036108f
C1069 VDD1.n156 VSUBS 0.016175f
C1070 VDD1.n157 VSUBS 0.015276f
C1071 VDD1.n158 VSUBS 0.028429f
C1072 VDD1.n159 VSUBS 0.028429f
C1073 VDD1.n160 VSUBS 0.015276f
C1074 VDD1.n161 VSUBS 0.015276f
C1075 VDD1.n162 VSUBS 0.016175f
C1076 VDD1.n163 VSUBS 0.036108f
C1077 VDD1.n164 VSUBS 0.036108f
C1078 VDD1.n165 VSUBS 0.036108f
C1079 VDD1.n166 VSUBS 0.015726f
C1080 VDD1.n167 VSUBS 0.015276f
C1081 VDD1.n168 VSUBS 0.028429f
C1082 VDD1.n169 VSUBS 0.028429f
C1083 VDD1.n170 VSUBS 0.015276f
C1084 VDD1.n171 VSUBS 0.016175f
C1085 VDD1.n172 VSUBS 0.036108f
C1086 VDD1.n173 VSUBS 0.089471f
C1087 VDD1.n174 VSUBS 0.016175f
C1088 VDD1.n175 VSUBS 0.015276f
C1089 VDD1.n176 VSUBS 0.072702f
C1090 VDD1.n177 VSUBS 1.03968f
C1091 VTAIL.n0 VSUBS 0.031698f
C1092 VTAIL.n1 VSUBS 0.028301f
C1093 VTAIL.n2 VSUBS 0.015208f
C1094 VTAIL.n3 VSUBS 0.035945f
C1095 VTAIL.n4 VSUBS 0.016102f
C1096 VTAIL.n5 VSUBS 0.028301f
C1097 VTAIL.n6 VSUBS 0.015655f
C1098 VTAIL.n7 VSUBS 0.035945f
C1099 VTAIL.n8 VSUBS 0.016102f
C1100 VTAIL.n9 VSUBS 0.028301f
C1101 VTAIL.n10 VSUBS 0.015208f
C1102 VTAIL.n11 VSUBS 0.035945f
C1103 VTAIL.n12 VSUBS 0.016102f
C1104 VTAIL.n13 VSUBS 0.028301f
C1105 VTAIL.n14 VSUBS 0.015208f
C1106 VTAIL.n15 VSUBS 0.035945f
C1107 VTAIL.n16 VSUBS 0.016102f
C1108 VTAIL.n17 VSUBS 0.028301f
C1109 VTAIL.n18 VSUBS 0.015208f
C1110 VTAIL.n19 VSUBS 0.035945f
C1111 VTAIL.n20 VSUBS 0.016102f
C1112 VTAIL.n21 VSUBS 0.028301f
C1113 VTAIL.n22 VSUBS 0.015208f
C1114 VTAIL.n23 VSUBS 0.035945f
C1115 VTAIL.n24 VSUBS 0.016102f
C1116 VTAIL.n25 VSUBS 0.028301f
C1117 VTAIL.n26 VSUBS 0.015208f
C1118 VTAIL.n27 VSUBS 0.026959f
C1119 VTAIL.n28 VSUBS 0.022867f
C1120 VTAIL.t0 VSUBS 0.07704f
C1121 VTAIL.n29 VSUBS 0.210013f
C1122 VTAIL.n30 VSUBS 1.96894f
C1123 VTAIL.n31 VSUBS 0.015208f
C1124 VTAIL.n32 VSUBS 0.016102f
C1125 VTAIL.n33 VSUBS 0.035945f
C1126 VTAIL.n34 VSUBS 0.035945f
C1127 VTAIL.n35 VSUBS 0.016102f
C1128 VTAIL.n36 VSUBS 0.015208f
C1129 VTAIL.n37 VSUBS 0.028301f
C1130 VTAIL.n38 VSUBS 0.028301f
C1131 VTAIL.n39 VSUBS 0.015208f
C1132 VTAIL.n40 VSUBS 0.016102f
C1133 VTAIL.n41 VSUBS 0.035945f
C1134 VTAIL.n42 VSUBS 0.035945f
C1135 VTAIL.n43 VSUBS 0.016102f
C1136 VTAIL.n44 VSUBS 0.015208f
C1137 VTAIL.n45 VSUBS 0.028301f
C1138 VTAIL.n46 VSUBS 0.028301f
C1139 VTAIL.n47 VSUBS 0.015208f
C1140 VTAIL.n48 VSUBS 0.016102f
C1141 VTAIL.n49 VSUBS 0.035945f
C1142 VTAIL.n50 VSUBS 0.035945f
C1143 VTAIL.n51 VSUBS 0.016102f
C1144 VTAIL.n52 VSUBS 0.015208f
C1145 VTAIL.n53 VSUBS 0.028301f
C1146 VTAIL.n54 VSUBS 0.028301f
C1147 VTAIL.n55 VSUBS 0.015208f
C1148 VTAIL.n56 VSUBS 0.016102f
C1149 VTAIL.n57 VSUBS 0.035945f
C1150 VTAIL.n58 VSUBS 0.035945f
C1151 VTAIL.n59 VSUBS 0.016102f
C1152 VTAIL.n60 VSUBS 0.015208f
C1153 VTAIL.n61 VSUBS 0.028301f
C1154 VTAIL.n62 VSUBS 0.028301f
C1155 VTAIL.n63 VSUBS 0.015208f
C1156 VTAIL.n64 VSUBS 0.016102f
C1157 VTAIL.n65 VSUBS 0.035945f
C1158 VTAIL.n66 VSUBS 0.035945f
C1159 VTAIL.n67 VSUBS 0.016102f
C1160 VTAIL.n68 VSUBS 0.015208f
C1161 VTAIL.n69 VSUBS 0.028301f
C1162 VTAIL.n70 VSUBS 0.028301f
C1163 VTAIL.n71 VSUBS 0.015208f
C1164 VTAIL.n72 VSUBS 0.015208f
C1165 VTAIL.n73 VSUBS 0.016102f
C1166 VTAIL.n74 VSUBS 0.035945f
C1167 VTAIL.n75 VSUBS 0.035945f
C1168 VTAIL.n76 VSUBS 0.035945f
C1169 VTAIL.n77 VSUBS 0.015655f
C1170 VTAIL.n78 VSUBS 0.015208f
C1171 VTAIL.n79 VSUBS 0.028301f
C1172 VTAIL.n80 VSUBS 0.028301f
C1173 VTAIL.n81 VSUBS 0.015208f
C1174 VTAIL.n82 VSUBS 0.016102f
C1175 VTAIL.n83 VSUBS 0.035945f
C1176 VTAIL.n84 VSUBS 0.089068f
C1177 VTAIL.n85 VSUBS 0.016102f
C1178 VTAIL.n86 VSUBS 0.015208f
C1179 VTAIL.n87 VSUBS 0.072375f
C1180 VTAIL.n88 VSUBS 0.045087f
C1181 VTAIL.n89 VSUBS 2.25543f
C1182 VTAIL.n90 VSUBS 0.031698f
C1183 VTAIL.n91 VSUBS 0.028301f
C1184 VTAIL.n92 VSUBS 0.015208f
C1185 VTAIL.n93 VSUBS 0.035945f
C1186 VTAIL.n94 VSUBS 0.016102f
C1187 VTAIL.n95 VSUBS 0.028301f
C1188 VTAIL.n96 VSUBS 0.015655f
C1189 VTAIL.n97 VSUBS 0.035945f
C1190 VTAIL.n98 VSUBS 0.015208f
C1191 VTAIL.n99 VSUBS 0.016102f
C1192 VTAIL.n100 VSUBS 0.028301f
C1193 VTAIL.n101 VSUBS 0.015208f
C1194 VTAIL.n102 VSUBS 0.035945f
C1195 VTAIL.n103 VSUBS 0.016102f
C1196 VTAIL.n104 VSUBS 0.028301f
C1197 VTAIL.n105 VSUBS 0.015208f
C1198 VTAIL.n106 VSUBS 0.035945f
C1199 VTAIL.n107 VSUBS 0.016102f
C1200 VTAIL.n108 VSUBS 0.028301f
C1201 VTAIL.n109 VSUBS 0.015208f
C1202 VTAIL.n110 VSUBS 0.035945f
C1203 VTAIL.n111 VSUBS 0.016102f
C1204 VTAIL.n112 VSUBS 0.028301f
C1205 VTAIL.n113 VSUBS 0.015208f
C1206 VTAIL.n114 VSUBS 0.035945f
C1207 VTAIL.n115 VSUBS 0.016102f
C1208 VTAIL.n116 VSUBS 0.028301f
C1209 VTAIL.n117 VSUBS 0.015208f
C1210 VTAIL.n118 VSUBS 0.026959f
C1211 VTAIL.n119 VSUBS 0.022867f
C1212 VTAIL.t3 VSUBS 0.07704f
C1213 VTAIL.n120 VSUBS 0.210013f
C1214 VTAIL.n121 VSUBS 1.96894f
C1215 VTAIL.n122 VSUBS 0.015208f
C1216 VTAIL.n123 VSUBS 0.016102f
C1217 VTAIL.n124 VSUBS 0.035945f
C1218 VTAIL.n125 VSUBS 0.035945f
C1219 VTAIL.n126 VSUBS 0.016102f
C1220 VTAIL.n127 VSUBS 0.015208f
C1221 VTAIL.n128 VSUBS 0.028301f
C1222 VTAIL.n129 VSUBS 0.028301f
C1223 VTAIL.n130 VSUBS 0.015208f
C1224 VTAIL.n131 VSUBS 0.016102f
C1225 VTAIL.n132 VSUBS 0.035945f
C1226 VTAIL.n133 VSUBS 0.035945f
C1227 VTAIL.n134 VSUBS 0.016102f
C1228 VTAIL.n135 VSUBS 0.015208f
C1229 VTAIL.n136 VSUBS 0.028301f
C1230 VTAIL.n137 VSUBS 0.028301f
C1231 VTAIL.n138 VSUBS 0.015208f
C1232 VTAIL.n139 VSUBS 0.016102f
C1233 VTAIL.n140 VSUBS 0.035945f
C1234 VTAIL.n141 VSUBS 0.035945f
C1235 VTAIL.n142 VSUBS 0.016102f
C1236 VTAIL.n143 VSUBS 0.015208f
C1237 VTAIL.n144 VSUBS 0.028301f
C1238 VTAIL.n145 VSUBS 0.028301f
C1239 VTAIL.n146 VSUBS 0.015208f
C1240 VTAIL.n147 VSUBS 0.016102f
C1241 VTAIL.n148 VSUBS 0.035945f
C1242 VTAIL.n149 VSUBS 0.035945f
C1243 VTAIL.n150 VSUBS 0.016102f
C1244 VTAIL.n151 VSUBS 0.015208f
C1245 VTAIL.n152 VSUBS 0.028301f
C1246 VTAIL.n153 VSUBS 0.028301f
C1247 VTAIL.n154 VSUBS 0.015208f
C1248 VTAIL.n155 VSUBS 0.016102f
C1249 VTAIL.n156 VSUBS 0.035945f
C1250 VTAIL.n157 VSUBS 0.035945f
C1251 VTAIL.n158 VSUBS 0.016102f
C1252 VTAIL.n159 VSUBS 0.015208f
C1253 VTAIL.n160 VSUBS 0.028301f
C1254 VTAIL.n161 VSUBS 0.028301f
C1255 VTAIL.n162 VSUBS 0.015208f
C1256 VTAIL.n163 VSUBS 0.016102f
C1257 VTAIL.n164 VSUBS 0.035945f
C1258 VTAIL.n165 VSUBS 0.035945f
C1259 VTAIL.n166 VSUBS 0.035945f
C1260 VTAIL.n167 VSUBS 0.015655f
C1261 VTAIL.n168 VSUBS 0.015208f
C1262 VTAIL.n169 VSUBS 0.028301f
C1263 VTAIL.n170 VSUBS 0.028301f
C1264 VTAIL.n171 VSUBS 0.015208f
C1265 VTAIL.n172 VSUBS 0.016102f
C1266 VTAIL.n173 VSUBS 0.035945f
C1267 VTAIL.n174 VSUBS 0.089068f
C1268 VTAIL.n175 VSUBS 0.016102f
C1269 VTAIL.n176 VSUBS 0.015208f
C1270 VTAIL.n177 VSUBS 0.072375f
C1271 VTAIL.n178 VSUBS 0.045087f
C1272 VTAIL.n179 VSUBS 2.30751f
C1273 VTAIL.n180 VSUBS 0.031698f
C1274 VTAIL.n181 VSUBS 0.028301f
C1275 VTAIL.n182 VSUBS 0.015208f
C1276 VTAIL.n183 VSUBS 0.035945f
C1277 VTAIL.n184 VSUBS 0.016102f
C1278 VTAIL.n185 VSUBS 0.028301f
C1279 VTAIL.n186 VSUBS 0.015655f
C1280 VTAIL.n187 VSUBS 0.035945f
C1281 VTAIL.n188 VSUBS 0.015208f
C1282 VTAIL.n189 VSUBS 0.016102f
C1283 VTAIL.n190 VSUBS 0.028301f
C1284 VTAIL.n191 VSUBS 0.015208f
C1285 VTAIL.n192 VSUBS 0.035945f
C1286 VTAIL.n193 VSUBS 0.016102f
C1287 VTAIL.n194 VSUBS 0.028301f
C1288 VTAIL.n195 VSUBS 0.015208f
C1289 VTAIL.n196 VSUBS 0.035945f
C1290 VTAIL.n197 VSUBS 0.016102f
C1291 VTAIL.n198 VSUBS 0.028301f
C1292 VTAIL.n199 VSUBS 0.015208f
C1293 VTAIL.n200 VSUBS 0.035945f
C1294 VTAIL.n201 VSUBS 0.016102f
C1295 VTAIL.n202 VSUBS 0.028301f
C1296 VTAIL.n203 VSUBS 0.015208f
C1297 VTAIL.n204 VSUBS 0.035945f
C1298 VTAIL.n205 VSUBS 0.016102f
C1299 VTAIL.n206 VSUBS 0.028301f
C1300 VTAIL.n207 VSUBS 0.015208f
C1301 VTAIL.n208 VSUBS 0.026959f
C1302 VTAIL.n209 VSUBS 0.022867f
C1303 VTAIL.t1 VSUBS 0.07704f
C1304 VTAIL.n210 VSUBS 0.210013f
C1305 VTAIL.n211 VSUBS 1.96894f
C1306 VTAIL.n212 VSUBS 0.015208f
C1307 VTAIL.n213 VSUBS 0.016102f
C1308 VTAIL.n214 VSUBS 0.035945f
C1309 VTAIL.n215 VSUBS 0.035945f
C1310 VTAIL.n216 VSUBS 0.016102f
C1311 VTAIL.n217 VSUBS 0.015208f
C1312 VTAIL.n218 VSUBS 0.028301f
C1313 VTAIL.n219 VSUBS 0.028301f
C1314 VTAIL.n220 VSUBS 0.015208f
C1315 VTAIL.n221 VSUBS 0.016102f
C1316 VTAIL.n222 VSUBS 0.035945f
C1317 VTAIL.n223 VSUBS 0.035945f
C1318 VTAIL.n224 VSUBS 0.016102f
C1319 VTAIL.n225 VSUBS 0.015208f
C1320 VTAIL.n226 VSUBS 0.028301f
C1321 VTAIL.n227 VSUBS 0.028301f
C1322 VTAIL.n228 VSUBS 0.015208f
C1323 VTAIL.n229 VSUBS 0.016102f
C1324 VTAIL.n230 VSUBS 0.035945f
C1325 VTAIL.n231 VSUBS 0.035945f
C1326 VTAIL.n232 VSUBS 0.016102f
C1327 VTAIL.n233 VSUBS 0.015208f
C1328 VTAIL.n234 VSUBS 0.028301f
C1329 VTAIL.n235 VSUBS 0.028301f
C1330 VTAIL.n236 VSUBS 0.015208f
C1331 VTAIL.n237 VSUBS 0.016102f
C1332 VTAIL.n238 VSUBS 0.035945f
C1333 VTAIL.n239 VSUBS 0.035945f
C1334 VTAIL.n240 VSUBS 0.016102f
C1335 VTAIL.n241 VSUBS 0.015208f
C1336 VTAIL.n242 VSUBS 0.028301f
C1337 VTAIL.n243 VSUBS 0.028301f
C1338 VTAIL.n244 VSUBS 0.015208f
C1339 VTAIL.n245 VSUBS 0.016102f
C1340 VTAIL.n246 VSUBS 0.035945f
C1341 VTAIL.n247 VSUBS 0.035945f
C1342 VTAIL.n248 VSUBS 0.016102f
C1343 VTAIL.n249 VSUBS 0.015208f
C1344 VTAIL.n250 VSUBS 0.028301f
C1345 VTAIL.n251 VSUBS 0.028301f
C1346 VTAIL.n252 VSUBS 0.015208f
C1347 VTAIL.n253 VSUBS 0.016102f
C1348 VTAIL.n254 VSUBS 0.035945f
C1349 VTAIL.n255 VSUBS 0.035945f
C1350 VTAIL.n256 VSUBS 0.035945f
C1351 VTAIL.n257 VSUBS 0.015655f
C1352 VTAIL.n258 VSUBS 0.015208f
C1353 VTAIL.n259 VSUBS 0.028301f
C1354 VTAIL.n260 VSUBS 0.028301f
C1355 VTAIL.n261 VSUBS 0.015208f
C1356 VTAIL.n262 VSUBS 0.016102f
C1357 VTAIL.n263 VSUBS 0.035945f
C1358 VTAIL.n264 VSUBS 0.089068f
C1359 VTAIL.n265 VSUBS 0.016102f
C1360 VTAIL.n266 VSUBS 0.015208f
C1361 VTAIL.n267 VSUBS 0.072375f
C1362 VTAIL.n268 VSUBS 0.045087f
C1363 VTAIL.n269 VSUBS 2.07796f
C1364 VTAIL.n270 VSUBS 0.031698f
C1365 VTAIL.n271 VSUBS 0.028301f
C1366 VTAIL.n272 VSUBS 0.015208f
C1367 VTAIL.n273 VSUBS 0.035945f
C1368 VTAIL.n274 VSUBS 0.016102f
C1369 VTAIL.n275 VSUBS 0.028301f
C1370 VTAIL.n276 VSUBS 0.015655f
C1371 VTAIL.n277 VSUBS 0.035945f
C1372 VTAIL.n278 VSUBS 0.016102f
C1373 VTAIL.n279 VSUBS 0.028301f
C1374 VTAIL.n280 VSUBS 0.015208f
C1375 VTAIL.n281 VSUBS 0.035945f
C1376 VTAIL.n282 VSUBS 0.016102f
C1377 VTAIL.n283 VSUBS 0.028301f
C1378 VTAIL.n284 VSUBS 0.015208f
C1379 VTAIL.n285 VSUBS 0.035945f
C1380 VTAIL.n286 VSUBS 0.016102f
C1381 VTAIL.n287 VSUBS 0.028301f
C1382 VTAIL.n288 VSUBS 0.015208f
C1383 VTAIL.n289 VSUBS 0.035945f
C1384 VTAIL.n290 VSUBS 0.016102f
C1385 VTAIL.n291 VSUBS 0.028301f
C1386 VTAIL.n292 VSUBS 0.015208f
C1387 VTAIL.n293 VSUBS 0.035945f
C1388 VTAIL.n294 VSUBS 0.016102f
C1389 VTAIL.n295 VSUBS 0.028301f
C1390 VTAIL.n296 VSUBS 0.015208f
C1391 VTAIL.n297 VSUBS 0.026959f
C1392 VTAIL.n298 VSUBS 0.022867f
C1393 VTAIL.t2 VSUBS 0.07704f
C1394 VTAIL.n299 VSUBS 0.210013f
C1395 VTAIL.n300 VSUBS 1.96894f
C1396 VTAIL.n301 VSUBS 0.015208f
C1397 VTAIL.n302 VSUBS 0.016102f
C1398 VTAIL.n303 VSUBS 0.035945f
C1399 VTAIL.n304 VSUBS 0.035945f
C1400 VTAIL.n305 VSUBS 0.016102f
C1401 VTAIL.n306 VSUBS 0.015208f
C1402 VTAIL.n307 VSUBS 0.028301f
C1403 VTAIL.n308 VSUBS 0.028301f
C1404 VTAIL.n309 VSUBS 0.015208f
C1405 VTAIL.n310 VSUBS 0.016102f
C1406 VTAIL.n311 VSUBS 0.035945f
C1407 VTAIL.n312 VSUBS 0.035945f
C1408 VTAIL.n313 VSUBS 0.016102f
C1409 VTAIL.n314 VSUBS 0.015208f
C1410 VTAIL.n315 VSUBS 0.028301f
C1411 VTAIL.n316 VSUBS 0.028301f
C1412 VTAIL.n317 VSUBS 0.015208f
C1413 VTAIL.n318 VSUBS 0.016102f
C1414 VTAIL.n319 VSUBS 0.035945f
C1415 VTAIL.n320 VSUBS 0.035945f
C1416 VTAIL.n321 VSUBS 0.016102f
C1417 VTAIL.n322 VSUBS 0.015208f
C1418 VTAIL.n323 VSUBS 0.028301f
C1419 VTAIL.n324 VSUBS 0.028301f
C1420 VTAIL.n325 VSUBS 0.015208f
C1421 VTAIL.n326 VSUBS 0.016102f
C1422 VTAIL.n327 VSUBS 0.035945f
C1423 VTAIL.n328 VSUBS 0.035945f
C1424 VTAIL.n329 VSUBS 0.016102f
C1425 VTAIL.n330 VSUBS 0.015208f
C1426 VTAIL.n331 VSUBS 0.028301f
C1427 VTAIL.n332 VSUBS 0.028301f
C1428 VTAIL.n333 VSUBS 0.015208f
C1429 VTAIL.n334 VSUBS 0.016102f
C1430 VTAIL.n335 VSUBS 0.035945f
C1431 VTAIL.n336 VSUBS 0.035945f
C1432 VTAIL.n337 VSUBS 0.016102f
C1433 VTAIL.n338 VSUBS 0.015208f
C1434 VTAIL.n339 VSUBS 0.028301f
C1435 VTAIL.n340 VSUBS 0.028301f
C1436 VTAIL.n341 VSUBS 0.015208f
C1437 VTAIL.n342 VSUBS 0.015208f
C1438 VTAIL.n343 VSUBS 0.016102f
C1439 VTAIL.n344 VSUBS 0.035945f
C1440 VTAIL.n345 VSUBS 0.035945f
C1441 VTAIL.n346 VSUBS 0.035945f
C1442 VTAIL.n347 VSUBS 0.015655f
C1443 VTAIL.n348 VSUBS 0.015208f
C1444 VTAIL.n349 VSUBS 0.028301f
C1445 VTAIL.n350 VSUBS 0.028301f
C1446 VTAIL.n351 VSUBS 0.015208f
C1447 VTAIL.n352 VSUBS 0.016102f
C1448 VTAIL.n353 VSUBS 0.035945f
C1449 VTAIL.n354 VSUBS 0.089068f
C1450 VTAIL.n355 VSUBS 0.016102f
C1451 VTAIL.n356 VSUBS 0.015208f
C1452 VTAIL.n357 VSUBS 0.072375f
C1453 VTAIL.n358 VSUBS 0.045087f
C1454 VTAIL.n359 VSUBS 1.97242f
C1455 VP.t1 VSUBS 5.5008f
C1456 VP.t0 VSUBS 4.83581f
C1457 VP.n0 VSUBS 6.17254f
.ends

