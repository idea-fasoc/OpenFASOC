* NGSPICE file created from diff_pair_sample_1760.ext - technology: sky130A

.subckt diff_pair_sample_1760 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=3.2109 ps=19.79 w=19.46 l=3.41
X1 B.t11 B.t9 B.t10 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=0 ps=0 w=19.46 l=3.41
X2 VDD1.t1 VP.t1 VTAIL.t6 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=3.2109 pd=19.79 as=7.5894 ps=39.7 w=19.46 l=3.41
X3 VDD1.t0 VP.t2 VTAIL.t5 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=3.2109 pd=19.79 as=7.5894 ps=39.7 w=19.46 l=3.41
X4 VDD2.t3 VN.t0 VTAIL.t2 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=3.2109 pd=19.79 as=7.5894 ps=39.7 w=19.46 l=3.41
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=3.2109 pd=19.79 as=7.5894 ps=39.7 w=19.46 l=3.41
X6 B.t8 B.t6 B.t7 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=0 ps=0 w=19.46 l=3.41
X7 VTAIL.t1 VN.t2 VDD2.t1 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=3.2109 ps=19.79 w=19.46 l=3.41
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=3.2109 ps=19.79 w=19.46 l=3.41
X9 B.t5 B.t3 B.t4 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=0 ps=0 w=19.46 l=3.41
X10 VTAIL.t4 VP.t3 VDD1.t3 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=3.2109 ps=19.79 w=19.46 l=3.41
X11 B.t2 B.t0 B.t1 w_n3214_n4860# sky130_fd_pr__pfet_01v8 ad=7.5894 pd=39.7 as=0 ps=0 w=19.46 l=3.41
R0 VP.n5 VP.t0 171.585
R1 VP.n5 VP.t2 170.387
R2 VP.n19 VP.n18 161.3
R3 VP.n17 VP.n1 161.3
R4 VP.n16 VP.n15 161.3
R5 VP.n14 VP.n2 161.3
R6 VP.n13 VP.n12 161.3
R7 VP.n11 VP.n3 161.3
R8 VP.n10 VP.n9 161.3
R9 VP.n8 VP.n4 161.3
R10 VP.n6 VP.t3 137.534
R11 VP.n0 VP.t1 137.534
R12 VP.n7 VP.n6 84.3435
R13 VP.n20 VP.n0 84.3435
R14 VP.n7 VP.n5 56.6938
R15 VP.n12 VP.n2 56.5617
R16 VP.n10 VP.n4 24.5923
R17 VP.n11 VP.n10 24.5923
R18 VP.n12 VP.n11 24.5923
R19 VP.n16 VP.n2 24.5923
R20 VP.n17 VP.n16 24.5923
R21 VP.n18 VP.n17 24.5923
R22 VP.n6 VP.n4 5.90254
R23 VP.n18 VP.n0 5.90254
R24 VP.n8 VP.n7 0.354861
R25 VP.n20 VP.n19 0.354861
R26 VP VP.n20 0.267071
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VDD1 VDD1.n1 121.246
R35 VDD1 VDD1.n0 70.6164
R36 VDD1.n0 VDD1.t2 1.67085
R37 VDD1.n0 VDD1.t0 1.67085
R38 VDD1.n1 VDD1.t3 1.67085
R39 VDD1.n1 VDD1.t1 1.67085
R40 VTAIL.n777 VTAIL.n776 585
R41 VTAIL.n774 VTAIL.n773 585
R42 VTAIL.n783 VTAIL.n782 585
R43 VTAIL.n785 VTAIL.n784 585
R44 VTAIL.n770 VTAIL.n769 585
R45 VTAIL.n791 VTAIL.n790 585
R46 VTAIL.n794 VTAIL.n793 585
R47 VTAIL.n792 VTAIL.n766 585
R48 VTAIL.n799 VTAIL.n765 585
R49 VTAIL.n801 VTAIL.n800 585
R50 VTAIL.n803 VTAIL.n802 585
R51 VTAIL.n762 VTAIL.n761 585
R52 VTAIL.n809 VTAIL.n808 585
R53 VTAIL.n811 VTAIL.n810 585
R54 VTAIL.n758 VTAIL.n757 585
R55 VTAIL.n817 VTAIL.n816 585
R56 VTAIL.n819 VTAIL.n818 585
R57 VTAIL.n754 VTAIL.n753 585
R58 VTAIL.n825 VTAIL.n824 585
R59 VTAIL.n827 VTAIL.n826 585
R60 VTAIL.n750 VTAIL.n749 585
R61 VTAIL.n833 VTAIL.n832 585
R62 VTAIL.n835 VTAIL.n834 585
R63 VTAIL.n746 VTAIL.n745 585
R64 VTAIL.n841 VTAIL.n840 585
R65 VTAIL.n843 VTAIL.n842 585
R66 VTAIL.n35 VTAIL.n34 585
R67 VTAIL.n32 VTAIL.n31 585
R68 VTAIL.n41 VTAIL.n40 585
R69 VTAIL.n43 VTAIL.n42 585
R70 VTAIL.n28 VTAIL.n27 585
R71 VTAIL.n49 VTAIL.n48 585
R72 VTAIL.n52 VTAIL.n51 585
R73 VTAIL.n50 VTAIL.n24 585
R74 VTAIL.n57 VTAIL.n23 585
R75 VTAIL.n59 VTAIL.n58 585
R76 VTAIL.n61 VTAIL.n60 585
R77 VTAIL.n20 VTAIL.n19 585
R78 VTAIL.n67 VTAIL.n66 585
R79 VTAIL.n69 VTAIL.n68 585
R80 VTAIL.n16 VTAIL.n15 585
R81 VTAIL.n75 VTAIL.n74 585
R82 VTAIL.n77 VTAIL.n76 585
R83 VTAIL.n12 VTAIL.n11 585
R84 VTAIL.n83 VTAIL.n82 585
R85 VTAIL.n85 VTAIL.n84 585
R86 VTAIL.n8 VTAIL.n7 585
R87 VTAIL.n91 VTAIL.n90 585
R88 VTAIL.n93 VTAIL.n92 585
R89 VTAIL.n4 VTAIL.n3 585
R90 VTAIL.n99 VTAIL.n98 585
R91 VTAIL.n101 VTAIL.n100 585
R92 VTAIL.n141 VTAIL.n140 585
R93 VTAIL.n138 VTAIL.n137 585
R94 VTAIL.n147 VTAIL.n146 585
R95 VTAIL.n149 VTAIL.n148 585
R96 VTAIL.n134 VTAIL.n133 585
R97 VTAIL.n155 VTAIL.n154 585
R98 VTAIL.n158 VTAIL.n157 585
R99 VTAIL.n156 VTAIL.n130 585
R100 VTAIL.n163 VTAIL.n129 585
R101 VTAIL.n165 VTAIL.n164 585
R102 VTAIL.n167 VTAIL.n166 585
R103 VTAIL.n126 VTAIL.n125 585
R104 VTAIL.n173 VTAIL.n172 585
R105 VTAIL.n175 VTAIL.n174 585
R106 VTAIL.n122 VTAIL.n121 585
R107 VTAIL.n181 VTAIL.n180 585
R108 VTAIL.n183 VTAIL.n182 585
R109 VTAIL.n118 VTAIL.n117 585
R110 VTAIL.n189 VTAIL.n188 585
R111 VTAIL.n191 VTAIL.n190 585
R112 VTAIL.n114 VTAIL.n113 585
R113 VTAIL.n197 VTAIL.n196 585
R114 VTAIL.n199 VTAIL.n198 585
R115 VTAIL.n110 VTAIL.n109 585
R116 VTAIL.n205 VTAIL.n204 585
R117 VTAIL.n207 VTAIL.n206 585
R118 VTAIL.n247 VTAIL.n246 585
R119 VTAIL.n244 VTAIL.n243 585
R120 VTAIL.n253 VTAIL.n252 585
R121 VTAIL.n255 VTAIL.n254 585
R122 VTAIL.n240 VTAIL.n239 585
R123 VTAIL.n261 VTAIL.n260 585
R124 VTAIL.n264 VTAIL.n263 585
R125 VTAIL.n262 VTAIL.n236 585
R126 VTAIL.n269 VTAIL.n235 585
R127 VTAIL.n271 VTAIL.n270 585
R128 VTAIL.n273 VTAIL.n272 585
R129 VTAIL.n232 VTAIL.n231 585
R130 VTAIL.n279 VTAIL.n278 585
R131 VTAIL.n281 VTAIL.n280 585
R132 VTAIL.n228 VTAIL.n227 585
R133 VTAIL.n287 VTAIL.n286 585
R134 VTAIL.n289 VTAIL.n288 585
R135 VTAIL.n224 VTAIL.n223 585
R136 VTAIL.n295 VTAIL.n294 585
R137 VTAIL.n297 VTAIL.n296 585
R138 VTAIL.n220 VTAIL.n219 585
R139 VTAIL.n303 VTAIL.n302 585
R140 VTAIL.n305 VTAIL.n304 585
R141 VTAIL.n216 VTAIL.n215 585
R142 VTAIL.n311 VTAIL.n310 585
R143 VTAIL.n313 VTAIL.n312 585
R144 VTAIL.n737 VTAIL.n736 585
R145 VTAIL.n735 VTAIL.n734 585
R146 VTAIL.n640 VTAIL.n639 585
R147 VTAIL.n729 VTAIL.n728 585
R148 VTAIL.n727 VTAIL.n726 585
R149 VTAIL.n644 VTAIL.n643 585
R150 VTAIL.n721 VTAIL.n720 585
R151 VTAIL.n719 VTAIL.n718 585
R152 VTAIL.n648 VTAIL.n647 585
R153 VTAIL.n713 VTAIL.n712 585
R154 VTAIL.n711 VTAIL.n710 585
R155 VTAIL.n652 VTAIL.n651 585
R156 VTAIL.n705 VTAIL.n704 585
R157 VTAIL.n703 VTAIL.n702 585
R158 VTAIL.n656 VTAIL.n655 585
R159 VTAIL.n697 VTAIL.n696 585
R160 VTAIL.n695 VTAIL.n694 585
R161 VTAIL.n693 VTAIL.n659 585
R162 VTAIL.n663 VTAIL.n660 585
R163 VTAIL.n688 VTAIL.n687 585
R164 VTAIL.n686 VTAIL.n685 585
R165 VTAIL.n665 VTAIL.n664 585
R166 VTAIL.n680 VTAIL.n679 585
R167 VTAIL.n678 VTAIL.n677 585
R168 VTAIL.n669 VTAIL.n668 585
R169 VTAIL.n672 VTAIL.n671 585
R170 VTAIL.n631 VTAIL.n630 585
R171 VTAIL.n629 VTAIL.n628 585
R172 VTAIL.n534 VTAIL.n533 585
R173 VTAIL.n623 VTAIL.n622 585
R174 VTAIL.n621 VTAIL.n620 585
R175 VTAIL.n538 VTAIL.n537 585
R176 VTAIL.n615 VTAIL.n614 585
R177 VTAIL.n613 VTAIL.n612 585
R178 VTAIL.n542 VTAIL.n541 585
R179 VTAIL.n607 VTAIL.n606 585
R180 VTAIL.n605 VTAIL.n604 585
R181 VTAIL.n546 VTAIL.n545 585
R182 VTAIL.n599 VTAIL.n598 585
R183 VTAIL.n597 VTAIL.n596 585
R184 VTAIL.n550 VTAIL.n549 585
R185 VTAIL.n591 VTAIL.n590 585
R186 VTAIL.n589 VTAIL.n588 585
R187 VTAIL.n587 VTAIL.n553 585
R188 VTAIL.n557 VTAIL.n554 585
R189 VTAIL.n582 VTAIL.n581 585
R190 VTAIL.n580 VTAIL.n579 585
R191 VTAIL.n559 VTAIL.n558 585
R192 VTAIL.n574 VTAIL.n573 585
R193 VTAIL.n572 VTAIL.n571 585
R194 VTAIL.n563 VTAIL.n562 585
R195 VTAIL.n566 VTAIL.n565 585
R196 VTAIL.n525 VTAIL.n524 585
R197 VTAIL.n523 VTAIL.n522 585
R198 VTAIL.n428 VTAIL.n427 585
R199 VTAIL.n517 VTAIL.n516 585
R200 VTAIL.n515 VTAIL.n514 585
R201 VTAIL.n432 VTAIL.n431 585
R202 VTAIL.n509 VTAIL.n508 585
R203 VTAIL.n507 VTAIL.n506 585
R204 VTAIL.n436 VTAIL.n435 585
R205 VTAIL.n501 VTAIL.n500 585
R206 VTAIL.n499 VTAIL.n498 585
R207 VTAIL.n440 VTAIL.n439 585
R208 VTAIL.n493 VTAIL.n492 585
R209 VTAIL.n491 VTAIL.n490 585
R210 VTAIL.n444 VTAIL.n443 585
R211 VTAIL.n485 VTAIL.n484 585
R212 VTAIL.n483 VTAIL.n482 585
R213 VTAIL.n481 VTAIL.n447 585
R214 VTAIL.n451 VTAIL.n448 585
R215 VTAIL.n476 VTAIL.n475 585
R216 VTAIL.n474 VTAIL.n473 585
R217 VTAIL.n453 VTAIL.n452 585
R218 VTAIL.n468 VTAIL.n467 585
R219 VTAIL.n466 VTAIL.n465 585
R220 VTAIL.n457 VTAIL.n456 585
R221 VTAIL.n460 VTAIL.n459 585
R222 VTAIL.n419 VTAIL.n418 585
R223 VTAIL.n417 VTAIL.n416 585
R224 VTAIL.n322 VTAIL.n321 585
R225 VTAIL.n411 VTAIL.n410 585
R226 VTAIL.n409 VTAIL.n408 585
R227 VTAIL.n326 VTAIL.n325 585
R228 VTAIL.n403 VTAIL.n402 585
R229 VTAIL.n401 VTAIL.n400 585
R230 VTAIL.n330 VTAIL.n329 585
R231 VTAIL.n395 VTAIL.n394 585
R232 VTAIL.n393 VTAIL.n392 585
R233 VTAIL.n334 VTAIL.n333 585
R234 VTAIL.n387 VTAIL.n386 585
R235 VTAIL.n385 VTAIL.n384 585
R236 VTAIL.n338 VTAIL.n337 585
R237 VTAIL.n379 VTAIL.n378 585
R238 VTAIL.n377 VTAIL.n376 585
R239 VTAIL.n375 VTAIL.n341 585
R240 VTAIL.n345 VTAIL.n342 585
R241 VTAIL.n370 VTAIL.n369 585
R242 VTAIL.n368 VTAIL.n367 585
R243 VTAIL.n347 VTAIL.n346 585
R244 VTAIL.n362 VTAIL.n361 585
R245 VTAIL.n360 VTAIL.n359 585
R246 VTAIL.n351 VTAIL.n350 585
R247 VTAIL.n354 VTAIL.n353 585
R248 VTAIL.n842 VTAIL.n742 498.474
R249 VTAIL.n100 VTAIL.n0 498.474
R250 VTAIL.n206 VTAIL.n106 498.474
R251 VTAIL.n312 VTAIL.n212 498.474
R252 VTAIL.n736 VTAIL.n636 498.474
R253 VTAIL.n630 VTAIL.n530 498.474
R254 VTAIL.n524 VTAIL.n424 498.474
R255 VTAIL.n418 VTAIL.n318 498.474
R256 VTAIL.t2 VTAIL.n775 329.036
R257 VTAIL.t1 VTAIL.n33 329.036
R258 VTAIL.t6 VTAIL.n139 329.036
R259 VTAIL.t4 VTAIL.n245 329.036
R260 VTAIL.t5 VTAIL.n670 329.036
R261 VTAIL.t7 VTAIL.n564 329.036
R262 VTAIL.t0 VTAIL.n458 329.036
R263 VTAIL.t3 VTAIL.n352 329.036
R264 VTAIL.n776 VTAIL.n773 171.744
R265 VTAIL.n783 VTAIL.n773 171.744
R266 VTAIL.n784 VTAIL.n783 171.744
R267 VTAIL.n784 VTAIL.n769 171.744
R268 VTAIL.n791 VTAIL.n769 171.744
R269 VTAIL.n793 VTAIL.n791 171.744
R270 VTAIL.n793 VTAIL.n792 171.744
R271 VTAIL.n792 VTAIL.n765 171.744
R272 VTAIL.n801 VTAIL.n765 171.744
R273 VTAIL.n802 VTAIL.n801 171.744
R274 VTAIL.n802 VTAIL.n761 171.744
R275 VTAIL.n809 VTAIL.n761 171.744
R276 VTAIL.n810 VTAIL.n809 171.744
R277 VTAIL.n810 VTAIL.n757 171.744
R278 VTAIL.n817 VTAIL.n757 171.744
R279 VTAIL.n818 VTAIL.n817 171.744
R280 VTAIL.n818 VTAIL.n753 171.744
R281 VTAIL.n825 VTAIL.n753 171.744
R282 VTAIL.n826 VTAIL.n825 171.744
R283 VTAIL.n826 VTAIL.n749 171.744
R284 VTAIL.n833 VTAIL.n749 171.744
R285 VTAIL.n834 VTAIL.n833 171.744
R286 VTAIL.n834 VTAIL.n745 171.744
R287 VTAIL.n841 VTAIL.n745 171.744
R288 VTAIL.n842 VTAIL.n841 171.744
R289 VTAIL.n34 VTAIL.n31 171.744
R290 VTAIL.n41 VTAIL.n31 171.744
R291 VTAIL.n42 VTAIL.n41 171.744
R292 VTAIL.n42 VTAIL.n27 171.744
R293 VTAIL.n49 VTAIL.n27 171.744
R294 VTAIL.n51 VTAIL.n49 171.744
R295 VTAIL.n51 VTAIL.n50 171.744
R296 VTAIL.n50 VTAIL.n23 171.744
R297 VTAIL.n59 VTAIL.n23 171.744
R298 VTAIL.n60 VTAIL.n59 171.744
R299 VTAIL.n60 VTAIL.n19 171.744
R300 VTAIL.n67 VTAIL.n19 171.744
R301 VTAIL.n68 VTAIL.n67 171.744
R302 VTAIL.n68 VTAIL.n15 171.744
R303 VTAIL.n75 VTAIL.n15 171.744
R304 VTAIL.n76 VTAIL.n75 171.744
R305 VTAIL.n76 VTAIL.n11 171.744
R306 VTAIL.n83 VTAIL.n11 171.744
R307 VTAIL.n84 VTAIL.n83 171.744
R308 VTAIL.n84 VTAIL.n7 171.744
R309 VTAIL.n91 VTAIL.n7 171.744
R310 VTAIL.n92 VTAIL.n91 171.744
R311 VTAIL.n92 VTAIL.n3 171.744
R312 VTAIL.n99 VTAIL.n3 171.744
R313 VTAIL.n100 VTAIL.n99 171.744
R314 VTAIL.n140 VTAIL.n137 171.744
R315 VTAIL.n147 VTAIL.n137 171.744
R316 VTAIL.n148 VTAIL.n147 171.744
R317 VTAIL.n148 VTAIL.n133 171.744
R318 VTAIL.n155 VTAIL.n133 171.744
R319 VTAIL.n157 VTAIL.n155 171.744
R320 VTAIL.n157 VTAIL.n156 171.744
R321 VTAIL.n156 VTAIL.n129 171.744
R322 VTAIL.n165 VTAIL.n129 171.744
R323 VTAIL.n166 VTAIL.n165 171.744
R324 VTAIL.n166 VTAIL.n125 171.744
R325 VTAIL.n173 VTAIL.n125 171.744
R326 VTAIL.n174 VTAIL.n173 171.744
R327 VTAIL.n174 VTAIL.n121 171.744
R328 VTAIL.n181 VTAIL.n121 171.744
R329 VTAIL.n182 VTAIL.n181 171.744
R330 VTAIL.n182 VTAIL.n117 171.744
R331 VTAIL.n189 VTAIL.n117 171.744
R332 VTAIL.n190 VTAIL.n189 171.744
R333 VTAIL.n190 VTAIL.n113 171.744
R334 VTAIL.n197 VTAIL.n113 171.744
R335 VTAIL.n198 VTAIL.n197 171.744
R336 VTAIL.n198 VTAIL.n109 171.744
R337 VTAIL.n205 VTAIL.n109 171.744
R338 VTAIL.n206 VTAIL.n205 171.744
R339 VTAIL.n246 VTAIL.n243 171.744
R340 VTAIL.n253 VTAIL.n243 171.744
R341 VTAIL.n254 VTAIL.n253 171.744
R342 VTAIL.n254 VTAIL.n239 171.744
R343 VTAIL.n261 VTAIL.n239 171.744
R344 VTAIL.n263 VTAIL.n261 171.744
R345 VTAIL.n263 VTAIL.n262 171.744
R346 VTAIL.n262 VTAIL.n235 171.744
R347 VTAIL.n271 VTAIL.n235 171.744
R348 VTAIL.n272 VTAIL.n271 171.744
R349 VTAIL.n272 VTAIL.n231 171.744
R350 VTAIL.n279 VTAIL.n231 171.744
R351 VTAIL.n280 VTAIL.n279 171.744
R352 VTAIL.n280 VTAIL.n227 171.744
R353 VTAIL.n287 VTAIL.n227 171.744
R354 VTAIL.n288 VTAIL.n287 171.744
R355 VTAIL.n288 VTAIL.n223 171.744
R356 VTAIL.n295 VTAIL.n223 171.744
R357 VTAIL.n296 VTAIL.n295 171.744
R358 VTAIL.n296 VTAIL.n219 171.744
R359 VTAIL.n303 VTAIL.n219 171.744
R360 VTAIL.n304 VTAIL.n303 171.744
R361 VTAIL.n304 VTAIL.n215 171.744
R362 VTAIL.n311 VTAIL.n215 171.744
R363 VTAIL.n312 VTAIL.n311 171.744
R364 VTAIL.n736 VTAIL.n735 171.744
R365 VTAIL.n735 VTAIL.n639 171.744
R366 VTAIL.n728 VTAIL.n639 171.744
R367 VTAIL.n728 VTAIL.n727 171.744
R368 VTAIL.n727 VTAIL.n643 171.744
R369 VTAIL.n720 VTAIL.n643 171.744
R370 VTAIL.n720 VTAIL.n719 171.744
R371 VTAIL.n719 VTAIL.n647 171.744
R372 VTAIL.n712 VTAIL.n647 171.744
R373 VTAIL.n712 VTAIL.n711 171.744
R374 VTAIL.n711 VTAIL.n651 171.744
R375 VTAIL.n704 VTAIL.n651 171.744
R376 VTAIL.n704 VTAIL.n703 171.744
R377 VTAIL.n703 VTAIL.n655 171.744
R378 VTAIL.n696 VTAIL.n655 171.744
R379 VTAIL.n696 VTAIL.n695 171.744
R380 VTAIL.n695 VTAIL.n659 171.744
R381 VTAIL.n663 VTAIL.n659 171.744
R382 VTAIL.n687 VTAIL.n663 171.744
R383 VTAIL.n687 VTAIL.n686 171.744
R384 VTAIL.n686 VTAIL.n664 171.744
R385 VTAIL.n679 VTAIL.n664 171.744
R386 VTAIL.n679 VTAIL.n678 171.744
R387 VTAIL.n678 VTAIL.n668 171.744
R388 VTAIL.n671 VTAIL.n668 171.744
R389 VTAIL.n630 VTAIL.n629 171.744
R390 VTAIL.n629 VTAIL.n533 171.744
R391 VTAIL.n622 VTAIL.n533 171.744
R392 VTAIL.n622 VTAIL.n621 171.744
R393 VTAIL.n621 VTAIL.n537 171.744
R394 VTAIL.n614 VTAIL.n537 171.744
R395 VTAIL.n614 VTAIL.n613 171.744
R396 VTAIL.n613 VTAIL.n541 171.744
R397 VTAIL.n606 VTAIL.n541 171.744
R398 VTAIL.n606 VTAIL.n605 171.744
R399 VTAIL.n605 VTAIL.n545 171.744
R400 VTAIL.n598 VTAIL.n545 171.744
R401 VTAIL.n598 VTAIL.n597 171.744
R402 VTAIL.n597 VTAIL.n549 171.744
R403 VTAIL.n590 VTAIL.n549 171.744
R404 VTAIL.n590 VTAIL.n589 171.744
R405 VTAIL.n589 VTAIL.n553 171.744
R406 VTAIL.n557 VTAIL.n553 171.744
R407 VTAIL.n581 VTAIL.n557 171.744
R408 VTAIL.n581 VTAIL.n580 171.744
R409 VTAIL.n580 VTAIL.n558 171.744
R410 VTAIL.n573 VTAIL.n558 171.744
R411 VTAIL.n573 VTAIL.n572 171.744
R412 VTAIL.n572 VTAIL.n562 171.744
R413 VTAIL.n565 VTAIL.n562 171.744
R414 VTAIL.n524 VTAIL.n523 171.744
R415 VTAIL.n523 VTAIL.n427 171.744
R416 VTAIL.n516 VTAIL.n427 171.744
R417 VTAIL.n516 VTAIL.n515 171.744
R418 VTAIL.n515 VTAIL.n431 171.744
R419 VTAIL.n508 VTAIL.n431 171.744
R420 VTAIL.n508 VTAIL.n507 171.744
R421 VTAIL.n507 VTAIL.n435 171.744
R422 VTAIL.n500 VTAIL.n435 171.744
R423 VTAIL.n500 VTAIL.n499 171.744
R424 VTAIL.n499 VTAIL.n439 171.744
R425 VTAIL.n492 VTAIL.n439 171.744
R426 VTAIL.n492 VTAIL.n491 171.744
R427 VTAIL.n491 VTAIL.n443 171.744
R428 VTAIL.n484 VTAIL.n443 171.744
R429 VTAIL.n484 VTAIL.n483 171.744
R430 VTAIL.n483 VTAIL.n447 171.744
R431 VTAIL.n451 VTAIL.n447 171.744
R432 VTAIL.n475 VTAIL.n451 171.744
R433 VTAIL.n475 VTAIL.n474 171.744
R434 VTAIL.n474 VTAIL.n452 171.744
R435 VTAIL.n467 VTAIL.n452 171.744
R436 VTAIL.n467 VTAIL.n466 171.744
R437 VTAIL.n466 VTAIL.n456 171.744
R438 VTAIL.n459 VTAIL.n456 171.744
R439 VTAIL.n418 VTAIL.n417 171.744
R440 VTAIL.n417 VTAIL.n321 171.744
R441 VTAIL.n410 VTAIL.n321 171.744
R442 VTAIL.n410 VTAIL.n409 171.744
R443 VTAIL.n409 VTAIL.n325 171.744
R444 VTAIL.n402 VTAIL.n325 171.744
R445 VTAIL.n402 VTAIL.n401 171.744
R446 VTAIL.n401 VTAIL.n329 171.744
R447 VTAIL.n394 VTAIL.n329 171.744
R448 VTAIL.n394 VTAIL.n393 171.744
R449 VTAIL.n393 VTAIL.n333 171.744
R450 VTAIL.n386 VTAIL.n333 171.744
R451 VTAIL.n386 VTAIL.n385 171.744
R452 VTAIL.n385 VTAIL.n337 171.744
R453 VTAIL.n378 VTAIL.n337 171.744
R454 VTAIL.n378 VTAIL.n377 171.744
R455 VTAIL.n377 VTAIL.n341 171.744
R456 VTAIL.n345 VTAIL.n341 171.744
R457 VTAIL.n369 VTAIL.n345 171.744
R458 VTAIL.n369 VTAIL.n368 171.744
R459 VTAIL.n368 VTAIL.n346 171.744
R460 VTAIL.n361 VTAIL.n346 171.744
R461 VTAIL.n361 VTAIL.n360 171.744
R462 VTAIL.n360 VTAIL.n350 171.744
R463 VTAIL.n353 VTAIL.n350 171.744
R464 VTAIL.n776 VTAIL.t2 85.8723
R465 VTAIL.n34 VTAIL.t1 85.8723
R466 VTAIL.n140 VTAIL.t6 85.8723
R467 VTAIL.n246 VTAIL.t4 85.8723
R468 VTAIL.n671 VTAIL.t5 85.8723
R469 VTAIL.n565 VTAIL.t7 85.8723
R470 VTAIL.n459 VTAIL.t0 85.8723
R471 VTAIL.n353 VTAIL.t3 85.8723
R472 VTAIL.n847 VTAIL.n846 34.9005
R473 VTAIL.n105 VTAIL.n104 34.9005
R474 VTAIL.n211 VTAIL.n210 34.9005
R475 VTAIL.n317 VTAIL.n316 34.9005
R476 VTAIL.n741 VTAIL.n740 34.9005
R477 VTAIL.n635 VTAIL.n634 34.9005
R478 VTAIL.n529 VTAIL.n528 34.9005
R479 VTAIL.n423 VTAIL.n422 34.9005
R480 VTAIL.n847 VTAIL.n741 32.3669
R481 VTAIL.n423 VTAIL.n317 32.3669
R482 VTAIL.n800 VTAIL.n799 13.1884
R483 VTAIL.n58 VTAIL.n57 13.1884
R484 VTAIL.n164 VTAIL.n163 13.1884
R485 VTAIL.n270 VTAIL.n269 13.1884
R486 VTAIL.n694 VTAIL.n693 13.1884
R487 VTAIL.n588 VTAIL.n587 13.1884
R488 VTAIL.n482 VTAIL.n481 13.1884
R489 VTAIL.n376 VTAIL.n375 13.1884
R490 VTAIL.n798 VTAIL.n766 12.8005
R491 VTAIL.n803 VTAIL.n764 12.8005
R492 VTAIL.n844 VTAIL.n843 12.8005
R493 VTAIL.n56 VTAIL.n24 12.8005
R494 VTAIL.n61 VTAIL.n22 12.8005
R495 VTAIL.n102 VTAIL.n101 12.8005
R496 VTAIL.n162 VTAIL.n130 12.8005
R497 VTAIL.n167 VTAIL.n128 12.8005
R498 VTAIL.n208 VTAIL.n207 12.8005
R499 VTAIL.n268 VTAIL.n236 12.8005
R500 VTAIL.n273 VTAIL.n234 12.8005
R501 VTAIL.n314 VTAIL.n313 12.8005
R502 VTAIL.n738 VTAIL.n737 12.8005
R503 VTAIL.n697 VTAIL.n658 12.8005
R504 VTAIL.n692 VTAIL.n660 12.8005
R505 VTAIL.n632 VTAIL.n631 12.8005
R506 VTAIL.n591 VTAIL.n552 12.8005
R507 VTAIL.n586 VTAIL.n554 12.8005
R508 VTAIL.n526 VTAIL.n525 12.8005
R509 VTAIL.n485 VTAIL.n446 12.8005
R510 VTAIL.n480 VTAIL.n448 12.8005
R511 VTAIL.n420 VTAIL.n419 12.8005
R512 VTAIL.n379 VTAIL.n340 12.8005
R513 VTAIL.n374 VTAIL.n342 12.8005
R514 VTAIL.n795 VTAIL.n794 12.0247
R515 VTAIL.n804 VTAIL.n762 12.0247
R516 VTAIL.n840 VTAIL.n744 12.0247
R517 VTAIL.n53 VTAIL.n52 12.0247
R518 VTAIL.n62 VTAIL.n20 12.0247
R519 VTAIL.n98 VTAIL.n2 12.0247
R520 VTAIL.n159 VTAIL.n158 12.0247
R521 VTAIL.n168 VTAIL.n126 12.0247
R522 VTAIL.n204 VTAIL.n108 12.0247
R523 VTAIL.n265 VTAIL.n264 12.0247
R524 VTAIL.n274 VTAIL.n232 12.0247
R525 VTAIL.n310 VTAIL.n214 12.0247
R526 VTAIL.n734 VTAIL.n638 12.0247
R527 VTAIL.n698 VTAIL.n656 12.0247
R528 VTAIL.n689 VTAIL.n688 12.0247
R529 VTAIL.n628 VTAIL.n532 12.0247
R530 VTAIL.n592 VTAIL.n550 12.0247
R531 VTAIL.n583 VTAIL.n582 12.0247
R532 VTAIL.n522 VTAIL.n426 12.0247
R533 VTAIL.n486 VTAIL.n444 12.0247
R534 VTAIL.n477 VTAIL.n476 12.0247
R535 VTAIL.n416 VTAIL.n320 12.0247
R536 VTAIL.n380 VTAIL.n338 12.0247
R537 VTAIL.n371 VTAIL.n370 12.0247
R538 VTAIL.n790 VTAIL.n768 11.249
R539 VTAIL.n808 VTAIL.n807 11.249
R540 VTAIL.n839 VTAIL.n746 11.249
R541 VTAIL.n48 VTAIL.n26 11.249
R542 VTAIL.n66 VTAIL.n65 11.249
R543 VTAIL.n97 VTAIL.n4 11.249
R544 VTAIL.n154 VTAIL.n132 11.249
R545 VTAIL.n172 VTAIL.n171 11.249
R546 VTAIL.n203 VTAIL.n110 11.249
R547 VTAIL.n260 VTAIL.n238 11.249
R548 VTAIL.n278 VTAIL.n277 11.249
R549 VTAIL.n309 VTAIL.n216 11.249
R550 VTAIL.n733 VTAIL.n640 11.249
R551 VTAIL.n702 VTAIL.n701 11.249
R552 VTAIL.n685 VTAIL.n662 11.249
R553 VTAIL.n627 VTAIL.n534 11.249
R554 VTAIL.n596 VTAIL.n595 11.249
R555 VTAIL.n579 VTAIL.n556 11.249
R556 VTAIL.n521 VTAIL.n428 11.249
R557 VTAIL.n490 VTAIL.n489 11.249
R558 VTAIL.n473 VTAIL.n450 11.249
R559 VTAIL.n415 VTAIL.n322 11.249
R560 VTAIL.n384 VTAIL.n383 11.249
R561 VTAIL.n367 VTAIL.n344 11.249
R562 VTAIL.n777 VTAIL.n775 10.7239
R563 VTAIL.n35 VTAIL.n33 10.7239
R564 VTAIL.n141 VTAIL.n139 10.7239
R565 VTAIL.n247 VTAIL.n245 10.7239
R566 VTAIL.n672 VTAIL.n670 10.7239
R567 VTAIL.n566 VTAIL.n564 10.7239
R568 VTAIL.n460 VTAIL.n458 10.7239
R569 VTAIL.n354 VTAIL.n352 10.7239
R570 VTAIL.n789 VTAIL.n770 10.4732
R571 VTAIL.n811 VTAIL.n760 10.4732
R572 VTAIL.n836 VTAIL.n835 10.4732
R573 VTAIL.n47 VTAIL.n28 10.4732
R574 VTAIL.n69 VTAIL.n18 10.4732
R575 VTAIL.n94 VTAIL.n93 10.4732
R576 VTAIL.n153 VTAIL.n134 10.4732
R577 VTAIL.n175 VTAIL.n124 10.4732
R578 VTAIL.n200 VTAIL.n199 10.4732
R579 VTAIL.n259 VTAIL.n240 10.4732
R580 VTAIL.n281 VTAIL.n230 10.4732
R581 VTAIL.n306 VTAIL.n305 10.4732
R582 VTAIL.n730 VTAIL.n729 10.4732
R583 VTAIL.n705 VTAIL.n654 10.4732
R584 VTAIL.n684 VTAIL.n665 10.4732
R585 VTAIL.n624 VTAIL.n623 10.4732
R586 VTAIL.n599 VTAIL.n548 10.4732
R587 VTAIL.n578 VTAIL.n559 10.4732
R588 VTAIL.n518 VTAIL.n517 10.4732
R589 VTAIL.n493 VTAIL.n442 10.4732
R590 VTAIL.n472 VTAIL.n453 10.4732
R591 VTAIL.n412 VTAIL.n411 10.4732
R592 VTAIL.n387 VTAIL.n336 10.4732
R593 VTAIL.n366 VTAIL.n347 10.4732
R594 VTAIL.n786 VTAIL.n785 9.69747
R595 VTAIL.n812 VTAIL.n758 9.69747
R596 VTAIL.n832 VTAIL.n748 9.69747
R597 VTAIL.n44 VTAIL.n43 9.69747
R598 VTAIL.n70 VTAIL.n16 9.69747
R599 VTAIL.n90 VTAIL.n6 9.69747
R600 VTAIL.n150 VTAIL.n149 9.69747
R601 VTAIL.n176 VTAIL.n122 9.69747
R602 VTAIL.n196 VTAIL.n112 9.69747
R603 VTAIL.n256 VTAIL.n255 9.69747
R604 VTAIL.n282 VTAIL.n228 9.69747
R605 VTAIL.n302 VTAIL.n218 9.69747
R606 VTAIL.n726 VTAIL.n642 9.69747
R607 VTAIL.n706 VTAIL.n652 9.69747
R608 VTAIL.n681 VTAIL.n680 9.69747
R609 VTAIL.n620 VTAIL.n536 9.69747
R610 VTAIL.n600 VTAIL.n546 9.69747
R611 VTAIL.n575 VTAIL.n574 9.69747
R612 VTAIL.n514 VTAIL.n430 9.69747
R613 VTAIL.n494 VTAIL.n440 9.69747
R614 VTAIL.n469 VTAIL.n468 9.69747
R615 VTAIL.n408 VTAIL.n324 9.69747
R616 VTAIL.n388 VTAIL.n334 9.69747
R617 VTAIL.n363 VTAIL.n362 9.69747
R618 VTAIL.n846 VTAIL.n845 9.45567
R619 VTAIL.n104 VTAIL.n103 9.45567
R620 VTAIL.n210 VTAIL.n209 9.45567
R621 VTAIL.n316 VTAIL.n315 9.45567
R622 VTAIL.n740 VTAIL.n739 9.45567
R623 VTAIL.n634 VTAIL.n633 9.45567
R624 VTAIL.n528 VTAIL.n527 9.45567
R625 VTAIL.n422 VTAIL.n421 9.45567
R626 VTAIL.n821 VTAIL.n820 9.3005
R627 VTAIL.n756 VTAIL.n755 9.3005
R628 VTAIL.n815 VTAIL.n814 9.3005
R629 VTAIL.n813 VTAIL.n812 9.3005
R630 VTAIL.n760 VTAIL.n759 9.3005
R631 VTAIL.n807 VTAIL.n806 9.3005
R632 VTAIL.n805 VTAIL.n804 9.3005
R633 VTAIL.n764 VTAIL.n763 9.3005
R634 VTAIL.n779 VTAIL.n778 9.3005
R635 VTAIL.n781 VTAIL.n780 9.3005
R636 VTAIL.n772 VTAIL.n771 9.3005
R637 VTAIL.n787 VTAIL.n786 9.3005
R638 VTAIL.n789 VTAIL.n788 9.3005
R639 VTAIL.n768 VTAIL.n767 9.3005
R640 VTAIL.n796 VTAIL.n795 9.3005
R641 VTAIL.n798 VTAIL.n797 9.3005
R642 VTAIL.n823 VTAIL.n822 9.3005
R643 VTAIL.n752 VTAIL.n751 9.3005
R644 VTAIL.n829 VTAIL.n828 9.3005
R645 VTAIL.n831 VTAIL.n830 9.3005
R646 VTAIL.n748 VTAIL.n747 9.3005
R647 VTAIL.n837 VTAIL.n836 9.3005
R648 VTAIL.n839 VTAIL.n838 9.3005
R649 VTAIL.n744 VTAIL.n743 9.3005
R650 VTAIL.n845 VTAIL.n844 9.3005
R651 VTAIL.n79 VTAIL.n78 9.3005
R652 VTAIL.n14 VTAIL.n13 9.3005
R653 VTAIL.n73 VTAIL.n72 9.3005
R654 VTAIL.n71 VTAIL.n70 9.3005
R655 VTAIL.n18 VTAIL.n17 9.3005
R656 VTAIL.n65 VTAIL.n64 9.3005
R657 VTAIL.n63 VTAIL.n62 9.3005
R658 VTAIL.n22 VTAIL.n21 9.3005
R659 VTAIL.n37 VTAIL.n36 9.3005
R660 VTAIL.n39 VTAIL.n38 9.3005
R661 VTAIL.n30 VTAIL.n29 9.3005
R662 VTAIL.n45 VTAIL.n44 9.3005
R663 VTAIL.n47 VTAIL.n46 9.3005
R664 VTAIL.n26 VTAIL.n25 9.3005
R665 VTAIL.n54 VTAIL.n53 9.3005
R666 VTAIL.n56 VTAIL.n55 9.3005
R667 VTAIL.n81 VTAIL.n80 9.3005
R668 VTAIL.n10 VTAIL.n9 9.3005
R669 VTAIL.n87 VTAIL.n86 9.3005
R670 VTAIL.n89 VTAIL.n88 9.3005
R671 VTAIL.n6 VTAIL.n5 9.3005
R672 VTAIL.n95 VTAIL.n94 9.3005
R673 VTAIL.n97 VTAIL.n96 9.3005
R674 VTAIL.n2 VTAIL.n1 9.3005
R675 VTAIL.n103 VTAIL.n102 9.3005
R676 VTAIL.n185 VTAIL.n184 9.3005
R677 VTAIL.n120 VTAIL.n119 9.3005
R678 VTAIL.n179 VTAIL.n178 9.3005
R679 VTAIL.n177 VTAIL.n176 9.3005
R680 VTAIL.n124 VTAIL.n123 9.3005
R681 VTAIL.n171 VTAIL.n170 9.3005
R682 VTAIL.n169 VTAIL.n168 9.3005
R683 VTAIL.n128 VTAIL.n127 9.3005
R684 VTAIL.n143 VTAIL.n142 9.3005
R685 VTAIL.n145 VTAIL.n144 9.3005
R686 VTAIL.n136 VTAIL.n135 9.3005
R687 VTAIL.n151 VTAIL.n150 9.3005
R688 VTAIL.n153 VTAIL.n152 9.3005
R689 VTAIL.n132 VTAIL.n131 9.3005
R690 VTAIL.n160 VTAIL.n159 9.3005
R691 VTAIL.n162 VTAIL.n161 9.3005
R692 VTAIL.n187 VTAIL.n186 9.3005
R693 VTAIL.n116 VTAIL.n115 9.3005
R694 VTAIL.n193 VTAIL.n192 9.3005
R695 VTAIL.n195 VTAIL.n194 9.3005
R696 VTAIL.n112 VTAIL.n111 9.3005
R697 VTAIL.n201 VTAIL.n200 9.3005
R698 VTAIL.n203 VTAIL.n202 9.3005
R699 VTAIL.n108 VTAIL.n107 9.3005
R700 VTAIL.n209 VTAIL.n208 9.3005
R701 VTAIL.n291 VTAIL.n290 9.3005
R702 VTAIL.n226 VTAIL.n225 9.3005
R703 VTAIL.n285 VTAIL.n284 9.3005
R704 VTAIL.n283 VTAIL.n282 9.3005
R705 VTAIL.n230 VTAIL.n229 9.3005
R706 VTAIL.n277 VTAIL.n276 9.3005
R707 VTAIL.n275 VTAIL.n274 9.3005
R708 VTAIL.n234 VTAIL.n233 9.3005
R709 VTAIL.n249 VTAIL.n248 9.3005
R710 VTAIL.n251 VTAIL.n250 9.3005
R711 VTAIL.n242 VTAIL.n241 9.3005
R712 VTAIL.n257 VTAIL.n256 9.3005
R713 VTAIL.n259 VTAIL.n258 9.3005
R714 VTAIL.n238 VTAIL.n237 9.3005
R715 VTAIL.n266 VTAIL.n265 9.3005
R716 VTAIL.n268 VTAIL.n267 9.3005
R717 VTAIL.n293 VTAIL.n292 9.3005
R718 VTAIL.n222 VTAIL.n221 9.3005
R719 VTAIL.n299 VTAIL.n298 9.3005
R720 VTAIL.n301 VTAIL.n300 9.3005
R721 VTAIL.n218 VTAIL.n217 9.3005
R722 VTAIL.n307 VTAIL.n306 9.3005
R723 VTAIL.n309 VTAIL.n308 9.3005
R724 VTAIL.n214 VTAIL.n213 9.3005
R725 VTAIL.n315 VTAIL.n314 9.3005
R726 VTAIL.n674 VTAIL.n673 9.3005
R727 VTAIL.n676 VTAIL.n675 9.3005
R728 VTAIL.n667 VTAIL.n666 9.3005
R729 VTAIL.n682 VTAIL.n681 9.3005
R730 VTAIL.n684 VTAIL.n683 9.3005
R731 VTAIL.n662 VTAIL.n661 9.3005
R732 VTAIL.n690 VTAIL.n689 9.3005
R733 VTAIL.n692 VTAIL.n691 9.3005
R734 VTAIL.n646 VTAIL.n645 9.3005
R735 VTAIL.n723 VTAIL.n722 9.3005
R736 VTAIL.n725 VTAIL.n724 9.3005
R737 VTAIL.n642 VTAIL.n641 9.3005
R738 VTAIL.n731 VTAIL.n730 9.3005
R739 VTAIL.n733 VTAIL.n732 9.3005
R740 VTAIL.n638 VTAIL.n637 9.3005
R741 VTAIL.n739 VTAIL.n738 9.3005
R742 VTAIL.n717 VTAIL.n716 9.3005
R743 VTAIL.n715 VTAIL.n714 9.3005
R744 VTAIL.n650 VTAIL.n649 9.3005
R745 VTAIL.n709 VTAIL.n708 9.3005
R746 VTAIL.n707 VTAIL.n706 9.3005
R747 VTAIL.n654 VTAIL.n653 9.3005
R748 VTAIL.n701 VTAIL.n700 9.3005
R749 VTAIL.n699 VTAIL.n698 9.3005
R750 VTAIL.n658 VTAIL.n657 9.3005
R751 VTAIL.n568 VTAIL.n567 9.3005
R752 VTAIL.n570 VTAIL.n569 9.3005
R753 VTAIL.n561 VTAIL.n560 9.3005
R754 VTAIL.n576 VTAIL.n575 9.3005
R755 VTAIL.n578 VTAIL.n577 9.3005
R756 VTAIL.n556 VTAIL.n555 9.3005
R757 VTAIL.n584 VTAIL.n583 9.3005
R758 VTAIL.n586 VTAIL.n585 9.3005
R759 VTAIL.n540 VTAIL.n539 9.3005
R760 VTAIL.n617 VTAIL.n616 9.3005
R761 VTAIL.n619 VTAIL.n618 9.3005
R762 VTAIL.n536 VTAIL.n535 9.3005
R763 VTAIL.n625 VTAIL.n624 9.3005
R764 VTAIL.n627 VTAIL.n626 9.3005
R765 VTAIL.n532 VTAIL.n531 9.3005
R766 VTAIL.n633 VTAIL.n632 9.3005
R767 VTAIL.n611 VTAIL.n610 9.3005
R768 VTAIL.n609 VTAIL.n608 9.3005
R769 VTAIL.n544 VTAIL.n543 9.3005
R770 VTAIL.n603 VTAIL.n602 9.3005
R771 VTAIL.n601 VTAIL.n600 9.3005
R772 VTAIL.n548 VTAIL.n547 9.3005
R773 VTAIL.n595 VTAIL.n594 9.3005
R774 VTAIL.n593 VTAIL.n592 9.3005
R775 VTAIL.n552 VTAIL.n551 9.3005
R776 VTAIL.n462 VTAIL.n461 9.3005
R777 VTAIL.n464 VTAIL.n463 9.3005
R778 VTAIL.n455 VTAIL.n454 9.3005
R779 VTAIL.n470 VTAIL.n469 9.3005
R780 VTAIL.n472 VTAIL.n471 9.3005
R781 VTAIL.n450 VTAIL.n449 9.3005
R782 VTAIL.n478 VTAIL.n477 9.3005
R783 VTAIL.n480 VTAIL.n479 9.3005
R784 VTAIL.n434 VTAIL.n433 9.3005
R785 VTAIL.n511 VTAIL.n510 9.3005
R786 VTAIL.n513 VTAIL.n512 9.3005
R787 VTAIL.n430 VTAIL.n429 9.3005
R788 VTAIL.n519 VTAIL.n518 9.3005
R789 VTAIL.n521 VTAIL.n520 9.3005
R790 VTAIL.n426 VTAIL.n425 9.3005
R791 VTAIL.n527 VTAIL.n526 9.3005
R792 VTAIL.n505 VTAIL.n504 9.3005
R793 VTAIL.n503 VTAIL.n502 9.3005
R794 VTAIL.n438 VTAIL.n437 9.3005
R795 VTAIL.n497 VTAIL.n496 9.3005
R796 VTAIL.n495 VTAIL.n494 9.3005
R797 VTAIL.n442 VTAIL.n441 9.3005
R798 VTAIL.n489 VTAIL.n488 9.3005
R799 VTAIL.n487 VTAIL.n486 9.3005
R800 VTAIL.n446 VTAIL.n445 9.3005
R801 VTAIL.n356 VTAIL.n355 9.3005
R802 VTAIL.n358 VTAIL.n357 9.3005
R803 VTAIL.n349 VTAIL.n348 9.3005
R804 VTAIL.n364 VTAIL.n363 9.3005
R805 VTAIL.n366 VTAIL.n365 9.3005
R806 VTAIL.n344 VTAIL.n343 9.3005
R807 VTAIL.n372 VTAIL.n371 9.3005
R808 VTAIL.n374 VTAIL.n373 9.3005
R809 VTAIL.n328 VTAIL.n327 9.3005
R810 VTAIL.n405 VTAIL.n404 9.3005
R811 VTAIL.n407 VTAIL.n406 9.3005
R812 VTAIL.n324 VTAIL.n323 9.3005
R813 VTAIL.n413 VTAIL.n412 9.3005
R814 VTAIL.n415 VTAIL.n414 9.3005
R815 VTAIL.n320 VTAIL.n319 9.3005
R816 VTAIL.n421 VTAIL.n420 9.3005
R817 VTAIL.n399 VTAIL.n398 9.3005
R818 VTAIL.n397 VTAIL.n396 9.3005
R819 VTAIL.n332 VTAIL.n331 9.3005
R820 VTAIL.n391 VTAIL.n390 9.3005
R821 VTAIL.n389 VTAIL.n388 9.3005
R822 VTAIL.n336 VTAIL.n335 9.3005
R823 VTAIL.n383 VTAIL.n382 9.3005
R824 VTAIL.n381 VTAIL.n380 9.3005
R825 VTAIL.n340 VTAIL.n339 9.3005
R826 VTAIL.n782 VTAIL.n772 8.92171
R827 VTAIL.n816 VTAIL.n815 8.92171
R828 VTAIL.n831 VTAIL.n750 8.92171
R829 VTAIL.n40 VTAIL.n30 8.92171
R830 VTAIL.n74 VTAIL.n73 8.92171
R831 VTAIL.n89 VTAIL.n8 8.92171
R832 VTAIL.n146 VTAIL.n136 8.92171
R833 VTAIL.n180 VTAIL.n179 8.92171
R834 VTAIL.n195 VTAIL.n114 8.92171
R835 VTAIL.n252 VTAIL.n242 8.92171
R836 VTAIL.n286 VTAIL.n285 8.92171
R837 VTAIL.n301 VTAIL.n220 8.92171
R838 VTAIL.n725 VTAIL.n644 8.92171
R839 VTAIL.n710 VTAIL.n709 8.92171
R840 VTAIL.n677 VTAIL.n667 8.92171
R841 VTAIL.n619 VTAIL.n538 8.92171
R842 VTAIL.n604 VTAIL.n603 8.92171
R843 VTAIL.n571 VTAIL.n561 8.92171
R844 VTAIL.n513 VTAIL.n432 8.92171
R845 VTAIL.n498 VTAIL.n497 8.92171
R846 VTAIL.n465 VTAIL.n455 8.92171
R847 VTAIL.n407 VTAIL.n326 8.92171
R848 VTAIL.n392 VTAIL.n391 8.92171
R849 VTAIL.n359 VTAIL.n349 8.92171
R850 VTAIL.n781 VTAIL.n774 8.14595
R851 VTAIL.n819 VTAIL.n756 8.14595
R852 VTAIL.n828 VTAIL.n827 8.14595
R853 VTAIL.n39 VTAIL.n32 8.14595
R854 VTAIL.n77 VTAIL.n14 8.14595
R855 VTAIL.n86 VTAIL.n85 8.14595
R856 VTAIL.n145 VTAIL.n138 8.14595
R857 VTAIL.n183 VTAIL.n120 8.14595
R858 VTAIL.n192 VTAIL.n191 8.14595
R859 VTAIL.n251 VTAIL.n244 8.14595
R860 VTAIL.n289 VTAIL.n226 8.14595
R861 VTAIL.n298 VTAIL.n297 8.14595
R862 VTAIL.n722 VTAIL.n721 8.14595
R863 VTAIL.n713 VTAIL.n650 8.14595
R864 VTAIL.n676 VTAIL.n669 8.14595
R865 VTAIL.n616 VTAIL.n615 8.14595
R866 VTAIL.n607 VTAIL.n544 8.14595
R867 VTAIL.n570 VTAIL.n563 8.14595
R868 VTAIL.n510 VTAIL.n509 8.14595
R869 VTAIL.n501 VTAIL.n438 8.14595
R870 VTAIL.n464 VTAIL.n457 8.14595
R871 VTAIL.n404 VTAIL.n403 8.14595
R872 VTAIL.n395 VTAIL.n332 8.14595
R873 VTAIL.n358 VTAIL.n351 8.14595
R874 VTAIL.n846 VTAIL.n742 7.75445
R875 VTAIL.n104 VTAIL.n0 7.75445
R876 VTAIL.n210 VTAIL.n106 7.75445
R877 VTAIL.n316 VTAIL.n212 7.75445
R878 VTAIL.n740 VTAIL.n636 7.75445
R879 VTAIL.n634 VTAIL.n530 7.75445
R880 VTAIL.n528 VTAIL.n424 7.75445
R881 VTAIL.n422 VTAIL.n318 7.75445
R882 VTAIL.n778 VTAIL.n777 7.3702
R883 VTAIL.n820 VTAIL.n754 7.3702
R884 VTAIL.n824 VTAIL.n752 7.3702
R885 VTAIL.n36 VTAIL.n35 7.3702
R886 VTAIL.n78 VTAIL.n12 7.3702
R887 VTAIL.n82 VTAIL.n10 7.3702
R888 VTAIL.n142 VTAIL.n141 7.3702
R889 VTAIL.n184 VTAIL.n118 7.3702
R890 VTAIL.n188 VTAIL.n116 7.3702
R891 VTAIL.n248 VTAIL.n247 7.3702
R892 VTAIL.n290 VTAIL.n224 7.3702
R893 VTAIL.n294 VTAIL.n222 7.3702
R894 VTAIL.n718 VTAIL.n646 7.3702
R895 VTAIL.n714 VTAIL.n648 7.3702
R896 VTAIL.n673 VTAIL.n672 7.3702
R897 VTAIL.n612 VTAIL.n540 7.3702
R898 VTAIL.n608 VTAIL.n542 7.3702
R899 VTAIL.n567 VTAIL.n566 7.3702
R900 VTAIL.n506 VTAIL.n434 7.3702
R901 VTAIL.n502 VTAIL.n436 7.3702
R902 VTAIL.n461 VTAIL.n460 7.3702
R903 VTAIL.n400 VTAIL.n328 7.3702
R904 VTAIL.n396 VTAIL.n330 7.3702
R905 VTAIL.n355 VTAIL.n354 7.3702
R906 VTAIL.n823 VTAIL.n754 6.59444
R907 VTAIL.n824 VTAIL.n823 6.59444
R908 VTAIL.n81 VTAIL.n12 6.59444
R909 VTAIL.n82 VTAIL.n81 6.59444
R910 VTAIL.n187 VTAIL.n118 6.59444
R911 VTAIL.n188 VTAIL.n187 6.59444
R912 VTAIL.n293 VTAIL.n224 6.59444
R913 VTAIL.n294 VTAIL.n293 6.59444
R914 VTAIL.n718 VTAIL.n717 6.59444
R915 VTAIL.n717 VTAIL.n648 6.59444
R916 VTAIL.n612 VTAIL.n611 6.59444
R917 VTAIL.n611 VTAIL.n542 6.59444
R918 VTAIL.n506 VTAIL.n505 6.59444
R919 VTAIL.n505 VTAIL.n436 6.59444
R920 VTAIL.n400 VTAIL.n399 6.59444
R921 VTAIL.n399 VTAIL.n330 6.59444
R922 VTAIL.n844 VTAIL.n742 6.08283
R923 VTAIL.n102 VTAIL.n0 6.08283
R924 VTAIL.n208 VTAIL.n106 6.08283
R925 VTAIL.n314 VTAIL.n212 6.08283
R926 VTAIL.n738 VTAIL.n636 6.08283
R927 VTAIL.n632 VTAIL.n530 6.08283
R928 VTAIL.n526 VTAIL.n424 6.08283
R929 VTAIL.n420 VTAIL.n318 6.08283
R930 VTAIL.n778 VTAIL.n774 5.81868
R931 VTAIL.n820 VTAIL.n819 5.81868
R932 VTAIL.n827 VTAIL.n752 5.81868
R933 VTAIL.n36 VTAIL.n32 5.81868
R934 VTAIL.n78 VTAIL.n77 5.81868
R935 VTAIL.n85 VTAIL.n10 5.81868
R936 VTAIL.n142 VTAIL.n138 5.81868
R937 VTAIL.n184 VTAIL.n183 5.81868
R938 VTAIL.n191 VTAIL.n116 5.81868
R939 VTAIL.n248 VTAIL.n244 5.81868
R940 VTAIL.n290 VTAIL.n289 5.81868
R941 VTAIL.n297 VTAIL.n222 5.81868
R942 VTAIL.n721 VTAIL.n646 5.81868
R943 VTAIL.n714 VTAIL.n713 5.81868
R944 VTAIL.n673 VTAIL.n669 5.81868
R945 VTAIL.n615 VTAIL.n540 5.81868
R946 VTAIL.n608 VTAIL.n607 5.81868
R947 VTAIL.n567 VTAIL.n563 5.81868
R948 VTAIL.n509 VTAIL.n434 5.81868
R949 VTAIL.n502 VTAIL.n501 5.81868
R950 VTAIL.n461 VTAIL.n457 5.81868
R951 VTAIL.n403 VTAIL.n328 5.81868
R952 VTAIL.n396 VTAIL.n395 5.81868
R953 VTAIL.n355 VTAIL.n351 5.81868
R954 VTAIL.n782 VTAIL.n781 5.04292
R955 VTAIL.n816 VTAIL.n756 5.04292
R956 VTAIL.n828 VTAIL.n750 5.04292
R957 VTAIL.n40 VTAIL.n39 5.04292
R958 VTAIL.n74 VTAIL.n14 5.04292
R959 VTAIL.n86 VTAIL.n8 5.04292
R960 VTAIL.n146 VTAIL.n145 5.04292
R961 VTAIL.n180 VTAIL.n120 5.04292
R962 VTAIL.n192 VTAIL.n114 5.04292
R963 VTAIL.n252 VTAIL.n251 5.04292
R964 VTAIL.n286 VTAIL.n226 5.04292
R965 VTAIL.n298 VTAIL.n220 5.04292
R966 VTAIL.n722 VTAIL.n644 5.04292
R967 VTAIL.n710 VTAIL.n650 5.04292
R968 VTAIL.n677 VTAIL.n676 5.04292
R969 VTAIL.n616 VTAIL.n538 5.04292
R970 VTAIL.n604 VTAIL.n544 5.04292
R971 VTAIL.n571 VTAIL.n570 5.04292
R972 VTAIL.n510 VTAIL.n432 5.04292
R973 VTAIL.n498 VTAIL.n438 5.04292
R974 VTAIL.n465 VTAIL.n464 5.04292
R975 VTAIL.n404 VTAIL.n326 5.04292
R976 VTAIL.n392 VTAIL.n332 5.04292
R977 VTAIL.n359 VTAIL.n358 5.04292
R978 VTAIL.n785 VTAIL.n772 4.26717
R979 VTAIL.n815 VTAIL.n758 4.26717
R980 VTAIL.n832 VTAIL.n831 4.26717
R981 VTAIL.n43 VTAIL.n30 4.26717
R982 VTAIL.n73 VTAIL.n16 4.26717
R983 VTAIL.n90 VTAIL.n89 4.26717
R984 VTAIL.n149 VTAIL.n136 4.26717
R985 VTAIL.n179 VTAIL.n122 4.26717
R986 VTAIL.n196 VTAIL.n195 4.26717
R987 VTAIL.n255 VTAIL.n242 4.26717
R988 VTAIL.n285 VTAIL.n228 4.26717
R989 VTAIL.n302 VTAIL.n301 4.26717
R990 VTAIL.n726 VTAIL.n725 4.26717
R991 VTAIL.n709 VTAIL.n652 4.26717
R992 VTAIL.n680 VTAIL.n667 4.26717
R993 VTAIL.n620 VTAIL.n619 4.26717
R994 VTAIL.n603 VTAIL.n546 4.26717
R995 VTAIL.n574 VTAIL.n561 4.26717
R996 VTAIL.n514 VTAIL.n513 4.26717
R997 VTAIL.n497 VTAIL.n440 4.26717
R998 VTAIL.n468 VTAIL.n455 4.26717
R999 VTAIL.n408 VTAIL.n407 4.26717
R1000 VTAIL.n391 VTAIL.n334 4.26717
R1001 VTAIL.n362 VTAIL.n349 4.26717
R1002 VTAIL.n786 VTAIL.n770 3.49141
R1003 VTAIL.n812 VTAIL.n811 3.49141
R1004 VTAIL.n835 VTAIL.n748 3.49141
R1005 VTAIL.n44 VTAIL.n28 3.49141
R1006 VTAIL.n70 VTAIL.n69 3.49141
R1007 VTAIL.n93 VTAIL.n6 3.49141
R1008 VTAIL.n150 VTAIL.n134 3.49141
R1009 VTAIL.n176 VTAIL.n175 3.49141
R1010 VTAIL.n199 VTAIL.n112 3.49141
R1011 VTAIL.n256 VTAIL.n240 3.49141
R1012 VTAIL.n282 VTAIL.n281 3.49141
R1013 VTAIL.n305 VTAIL.n218 3.49141
R1014 VTAIL.n729 VTAIL.n642 3.49141
R1015 VTAIL.n706 VTAIL.n705 3.49141
R1016 VTAIL.n681 VTAIL.n665 3.49141
R1017 VTAIL.n623 VTAIL.n536 3.49141
R1018 VTAIL.n600 VTAIL.n599 3.49141
R1019 VTAIL.n575 VTAIL.n559 3.49141
R1020 VTAIL.n517 VTAIL.n430 3.49141
R1021 VTAIL.n494 VTAIL.n493 3.49141
R1022 VTAIL.n469 VTAIL.n453 3.49141
R1023 VTAIL.n411 VTAIL.n324 3.49141
R1024 VTAIL.n388 VTAIL.n387 3.49141
R1025 VTAIL.n363 VTAIL.n347 3.49141
R1026 VTAIL.n529 VTAIL.n423 3.22464
R1027 VTAIL.n741 VTAIL.n635 3.22464
R1028 VTAIL.n317 VTAIL.n211 3.22464
R1029 VTAIL.n790 VTAIL.n789 2.71565
R1030 VTAIL.n808 VTAIL.n760 2.71565
R1031 VTAIL.n836 VTAIL.n746 2.71565
R1032 VTAIL.n48 VTAIL.n47 2.71565
R1033 VTAIL.n66 VTAIL.n18 2.71565
R1034 VTAIL.n94 VTAIL.n4 2.71565
R1035 VTAIL.n154 VTAIL.n153 2.71565
R1036 VTAIL.n172 VTAIL.n124 2.71565
R1037 VTAIL.n200 VTAIL.n110 2.71565
R1038 VTAIL.n260 VTAIL.n259 2.71565
R1039 VTAIL.n278 VTAIL.n230 2.71565
R1040 VTAIL.n306 VTAIL.n216 2.71565
R1041 VTAIL.n730 VTAIL.n640 2.71565
R1042 VTAIL.n702 VTAIL.n654 2.71565
R1043 VTAIL.n685 VTAIL.n684 2.71565
R1044 VTAIL.n624 VTAIL.n534 2.71565
R1045 VTAIL.n596 VTAIL.n548 2.71565
R1046 VTAIL.n579 VTAIL.n578 2.71565
R1047 VTAIL.n518 VTAIL.n428 2.71565
R1048 VTAIL.n490 VTAIL.n442 2.71565
R1049 VTAIL.n473 VTAIL.n472 2.71565
R1050 VTAIL.n412 VTAIL.n322 2.71565
R1051 VTAIL.n384 VTAIL.n336 2.71565
R1052 VTAIL.n367 VTAIL.n366 2.71565
R1053 VTAIL.n674 VTAIL.n670 2.41282
R1054 VTAIL.n568 VTAIL.n564 2.41282
R1055 VTAIL.n462 VTAIL.n458 2.41282
R1056 VTAIL.n356 VTAIL.n352 2.41282
R1057 VTAIL.n779 VTAIL.n775 2.41282
R1058 VTAIL.n37 VTAIL.n33 2.41282
R1059 VTAIL.n143 VTAIL.n139 2.41282
R1060 VTAIL.n249 VTAIL.n245 2.41282
R1061 VTAIL.n794 VTAIL.n768 1.93989
R1062 VTAIL.n807 VTAIL.n762 1.93989
R1063 VTAIL.n840 VTAIL.n839 1.93989
R1064 VTAIL.n52 VTAIL.n26 1.93989
R1065 VTAIL.n65 VTAIL.n20 1.93989
R1066 VTAIL.n98 VTAIL.n97 1.93989
R1067 VTAIL.n158 VTAIL.n132 1.93989
R1068 VTAIL.n171 VTAIL.n126 1.93989
R1069 VTAIL.n204 VTAIL.n203 1.93989
R1070 VTAIL.n264 VTAIL.n238 1.93989
R1071 VTAIL.n277 VTAIL.n232 1.93989
R1072 VTAIL.n310 VTAIL.n309 1.93989
R1073 VTAIL.n734 VTAIL.n733 1.93989
R1074 VTAIL.n701 VTAIL.n656 1.93989
R1075 VTAIL.n688 VTAIL.n662 1.93989
R1076 VTAIL.n628 VTAIL.n627 1.93989
R1077 VTAIL.n595 VTAIL.n550 1.93989
R1078 VTAIL.n582 VTAIL.n556 1.93989
R1079 VTAIL.n522 VTAIL.n521 1.93989
R1080 VTAIL.n489 VTAIL.n444 1.93989
R1081 VTAIL.n476 VTAIL.n450 1.93989
R1082 VTAIL.n416 VTAIL.n415 1.93989
R1083 VTAIL.n383 VTAIL.n338 1.93989
R1084 VTAIL.n370 VTAIL.n344 1.93989
R1085 VTAIL VTAIL.n105 1.67076
R1086 VTAIL VTAIL.n847 1.55438
R1087 VTAIL.n795 VTAIL.n766 1.16414
R1088 VTAIL.n804 VTAIL.n803 1.16414
R1089 VTAIL.n843 VTAIL.n744 1.16414
R1090 VTAIL.n53 VTAIL.n24 1.16414
R1091 VTAIL.n62 VTAIL.n61 1.16414
R1092 VTAIL.n101 VTAIL.n2 1.16414
R1093 VTAIL.n159 VTAIL.n130 1.16414
R1094 VTAIL.n168 VTAIL.n167 1.16414
R1095 VTAIL.n207 VTAIL.n108 1.16414
R1096 VTAIL.n265 VTAIL.n236 1.16414
R1097 VTAIL.n274 VTAIL.n273 1.16414
R1098 VTAIL.n313 VTAIL.n214 1.16414
R1099 VTAIL.n737 VTAIL.n638 1.16414
R1100 VTAIL.n698 VTAIL.n697 1.16414
R1101 VTAIL.n689 VTAIL.n660 1.16414
R1102 VTAIL.n631 VTAIL.n532 1.16414
R1103 VTAIL.n592 VTAIL.n591 1.16414
R1104 VTAIL.n583 VTAIL.n554 1.16414
R1105 VTAIL.n525 VTAIL.n426 1.16414
R1106 VTAIL.n486 VTAIL.n485 1.16414
R1107 VTAIL.n477 VTAIL.n448 1.16414
R1108 VTAIL.n419 VTAIL.n320 1.16414
R1109 VTAIL.n380 VTAIL.n379 1.16414
R1110 VTAIL.n371 VTAIL.n342 1.16414
R1111 VTAIL.n635 VTAIL.n529 0.470328
R1112 VTAIL.n211 VTAIL.n105 0.470328
R1113 VTAIL.n799 VTAIL.n798 0.388379
R1114 VTAIL.n800 VTAIL.n764 0.388379
R1115 VTAIL.n57 VTAIL.n56 0.388379
R1116 VTAIL.n58 VTAIL.n22 0.388379
R1117 VTAIL.n163 VTAIL.n162 0.388379
R1118 VTAIL.n164 VTAIL.n128 0.388379
R1119 VTAIL.n269 VTAIL.n268 0.388379
R1120 VTAIL.n270 VTAIL.n234 0.388379
R1121 VTAIL.n694 VTAIL.n658 0.388379
R1122 VTAIL.n693 VTAIL.n692 0.388379
R1123 VTAIL.n588 VTAIL.n552 0.388379
R1124 VTAIL.n587 VTAIL.n586 0.388379
R1125 VTAIL.n482 VTAIL.n446 0.388379
R1126 VTAIL.n481 VTAIL.n480 0.388379
R1127 VTAIL.n376 VTAIL.n340 0.388379
R1128 VTAIL.n375 VTAIL.n374 0.388379
R1129 VTAIL.n780 VTAIL.n779 0.155672
R1130 VTAIL.n780 VTAIL.n771 0.155672
R1131 VTAIL.n787 VTAIL.n771 0.155672
R1132 VTAIL.n788 VTAIL.n787 0.155672
R1133 VTAIL.n788 VTAIL.n767 0.155672
R1134 VTAIL.n796 VTAIL.n767 0.155672
R1135 VTAIL.n797 VTAIL.n796 0.155672
R1136 VTAIL.n797 VTAIL.n763 0.155672
R1137 VTAIL.n805 VTAIL.n763 0.155672
R1138 VTAIL.n806 VTAIL.n805 0.155672
R1139 VTAIL.n806 VTAIL.n759 0.155672
R1140 VTAIL.n813 VTAIL.n759 0.155672
R1141 VTAIL.n814 VTAIL.n813 0.155672
R1142 VTAIL.n814 VTAIL.n755 0.155672
R1143 VTAIL.n821 VTAIL.n755 0.155672
R1144 VTAIL.n822 VTAIL.n821 0.155672
R1145 VTAIL.n822 VTAIL.n751 0.155672
R1146 VTAIL.n829 VTAIL.n751 0.155672
R1147 VTAIL.n830 VTAIL.n829 0.155672
R1148 VTAIL.n830 VTAIL.n747 0.155672
R1149 VTAIL.n837 VTAIL.n747 0.155672
R1150 VTAIL.n838 VTAIL.n837 0.155672
R1151 VTAIL.n838 VTAIL.n743 0.155672
R1152 VTAIL.n845 VTAIL.n743 0.155672
R1153 VTAIL.n38 VTAIL.n37 0.155672
R1154 VTAIL.n38 VTAIL.n29 0.155672
R1155 VTAIL.n45 VTAIL.n29 0.155672
R1156 VTAIL.n46 VTAIL.n45 0.155672
R1157 VTAIL.n46 VTAIL.n25 0.155672
R1158 VTAIL.n54 VTAIL.n25 0.155672
R1159 VTAIL.n55 VTAIL.n54 0.155672
R1160 VTAIL.n55 VTAIL.n21 0.155672
R1161 VTAIL.n63 VTAIL.n21 0.155672
R1162 VTAIL.n64 VTAIL.n63 0.155672
R1163 VTAIL.n64 VTAIL.n17 0.155672
R1164 VTAIL.n71 VTAIL.n17 0.155672
R1165 VTAIL.n72 VTAIL.n71 0.155672
R1166 VTAIL.n72 VTAIL.n13 0.155672
R1167 VTAIL.n79 VTAIL.n13 0.155672
R1168 VTAIL.n80 VTAIL.n79 0.155672
R1169 VTAIL.n80 VTAIL.n9 0.155672
R1170 VTAIL.n87 VTAIL.n9 0.155672
R1171 VTAIL.n88 VTAIL.n87 0.155672
R1172 VTAIL.n88 VTAIL.n5 0.155672
R1173 VTAIL.n95 VTAIL.n5 0.155672
R1174 VTAIL.n96 VTAIL.n95 0.155672
R1175 VTAIL.n96 VTAIL.n1 0.155672
R1176 VTAIL.n103 VTAIL.n1 0.155672
R1177 VTAIL.n144 VTAIL.n143 0.155672
R1178 VTAIL.n144 VTAIL.n135 0.155672
R1179 VTAIL.n151 VTAIL.n135 0.155672
R1180 VTAIL.n152 VTAIL.n151 0.155672
R1181 VTAIL.n152 VTAIL.n131 0.155672
R1182 VTAIL.n160 VTAIL.n131 0.155672
R1183 VTAIL.n161 VTAIL.n160 0.155672
R1184 VTAIL.n161 VTAIL.n127 0.155672
R1185 VTAIL.n169 VTAIL.n127 0.155672
R1186 VTAIL.n170 VTAIL.n169 0.155672
R1187 VTAIL.n170 VTAIL.n123 0.155672
R1188 VTAIL.n177 VTAIL.n123 0.155672
R1189 VTAIL.n178 VTAIL.n177 0.155672
R1190 VTAIL.n178 VTAIL.n119 0.155672
R1191 VTAIL.n185 VTAIL.n119 0.155672
R1192 VTAIL.n186 VTAIL.n185 0.155672
R1193 VTAIL.n186 VTAIL.n115 0.155672
R1194 VTAIL.n193 VTAIL.n115 0.155672
R1195 VTAIL.n194 VTAIL.n193 0.155672
R1196 VTAIL.n194 VTAIL.n111 0.155672
R1197 VTAIL.n201 VTAIL.n111 0.155672
R1198 VTAIL.n202 VTAIL.n201 0.155672
R1199 VTAIL.n202 VTAIL.n107 0.155672
R1200 VTAIL.n209 VTAIL.n107 0.155672
R1201 VTAIL.n250 VTAIL.n249 0.155672
R1202 VTAIL.n250 VTAIL.n241 0.155672
R1203 VTAIL.n257 VTAIL.n241 0.155672
R1204 VTAIL.n258 VTAIL.n257 0.155672
R1205 VTAIL.n258 VTAIL.n237 0.155672
R1206 VTAIL.n266 VTAIL.n237 0.155672
R1207 VTAIL.n267 VTAIL.n266 0.155672
R1208 VTAIL.n267 VTAIL.n233 0.155672
R1209 VTAIL.n275 VTAIL.n233 0.155672
R1210 VTAIL.n276 VTAIL.n275 0.155672
R1211 VTAIL.n276 VTAIL.n229 0.155672
R1212 VTAIL.n283 VTAIL.n229 0.155672
R1213 VTAIL.n284 VTAIL.n283 0.155672
R1214 VTAIL.n284 VTAIL.n225 0.155672
R1215 VTAIL.n291 VTAIL.n225 0.155672
R1216 VTAIL.n292 VTAIL.n291 0.155672
R1217 VTAIL.n292 VTAIL.n221 0.155672
R1218 VTAIL.n299 VTAIL.n221 0.155672
R1219 VTAIL.n300 VTAIL.n299 0.155672
R1220 VTAIL.n300 VTAIL.n217 0.155672
R1221 VTAIL.n307 VTAIL.n217 0.155672
R1222 VTAIL.n308 VTAIL.n307 0.155672
R1223 VTAIL.n308 VTAIL.n213 0.155672
R1224 VTAIL.n315 VTAIL.n213 0.155672
R1225 VTAIL.n739 VTAIL.n637 0.155672
R1226 VTAIL.n732 VTAIL.n637 0.155672
R1227 VTAIL.n732 VTAIL.n731 0.155672
R1228 VTAIL.n731 VTAIL.n641 0.155672
R1229 VTAIL.n724 VTAIL.n641 0.155672
R1230 VTAIL.n724 VTAIL.n723 0.155672
R1231 VTAIL.n723 VTAIL.n645 0.155672
R1232 VTAIL.n716 VTAIL.n645 0.155672
R1233 VTAIL.n716 VTAIL.n715 0.155672
R1234 VTAIL.n715 VTAIL.n649 0.155672
R1235 VTAIL.n708 VTAIL.n649 0.155672
R1236 VTAIL.n708 VTAIL.n707 0.155672
R1237 VTAIL.n707 VTAIL.n653 0.155672
R1238 VTAIL.n700 VTAIL.n653 0.155672
R1239 VTAIL.n700 VTAIL.n699 0.155672
R1240 VTAIL.n699 VTAIL.n657 0.155672
R1241 VTAIL.n691 VTAIL.n657 0.155672
R1242 VTAIL.n691 VTAIL.n690 0.155672
R1243 VTAIL.n690 VTAIL.n661 0.155672
R1244 VTAIL.n683 VTAIL.n661 0.155672
R1245 VTAIL.n683 VTAIL.n682 0.155672
R1246 VTAIL.n682 VTAIL.n666 0.155672
R1247 VTAIL.n675 VTAIL.n666 0.155672
R1248 VTAIL.n675 VTAIL.n674 0.155672
R1249 VTAIL.n633 VTAIL.n531 0.155672
R1250 VTAIL.n626 VTAIL.n531 0.155672
R1251 VTAIL.n626 VTAIL.n625 0.155672
R1252 VTAIL.n625 VTAIL.n535 0.155672
R1253 VTAIL.n618 VTAIL.n535 0.155672
R1254 VTAIL.n618 VTAIL.n617 0.155672
R1255 VTAIL.n617 VTAIL.n539 0.155672
R1256 VTAIL.n610 VTAIL.n539 0.155672
R1257 VTAIL.n610 VTAIL.n609 0.155672
R1258 VTAIL.n609 VTAIL.n543 0.155672
R1259 VTAIL.n602 VTAIL.n543 0.155672
R1260 VTAIL.n602 VTAIL.n601 0.155672
R1261 VTAIL.n601 VTAIL.n547 0.155672
R1262 VTAIL.n594 VTAIL.n547 0.155672
R1263 VTAIL.n594 VTAIL.n593 0.155672
R1264 VTAIL.n593 VTAIL.n551 0.155672
R1265 VTAIL.n585 VTAIL.n551 0.155672
R1266 VTAIL.n585 VTAIL.n584 0.155672
R1267 VTAIL.n584 VTAIL.n555 0.155672
R1268 VTAIL.n577 VTAIL.n555 0.155672
R1269 VTAIL.n577 VTAIL.n576 0.155672
R1270 VTAIL.n576 VTAIL.n560 0.155672
R1271 VTAIL.n569 VTAIL.n560 0.155672
R1272 VTAIL.n569 VTAIL.n568 0.155672
R1273 VTAIL.n527 VTAIL.n425 0.155672
R1274 VTAIL.n520 VTAIL.n425 0.155672
R1275 VTAIL.n520 VTAIL.n519 0.155672
R1276 VTAIL.n519 VTAIL.n429 0.155672
R1277 VTAIL.n512 VTAIL.n429 0.155672
R1278 VTAIL.n512 VTAIL.n511 0.155672
R1279 VTAIL.n511 VTAIL.n433 0.155672
R1280 VTAIL.n504 VTAIL.n433 0.155672
R1281 VTAIL.n504 VTAIL.n503 0.155672
R1282 VTAIL.n503 VTAIL.n437 0.155672
R1283 VTAIL.n496 VTAIL.n437 0.155672
R1284 VTAIL.n496 VTAIL.n495 0.155672
R1285 VTAIL.n495 VTAIL.n441 0.155672
R1286 VTAIL.n488 VTAIL.n441 0.155672
R1287 VTAIL.n488 VTAIL.n487 0.155672
R1288 VTAIL.n487 VTAIL.n445 0.155672
R1289 VTAIL.n479 VTAIL.n445 0.155672
R1290 VTAIL.n479 VTAIL.n478 0.155672
R1291 VTAIL.n478 VTAIL.n449 0.155672
R1292 VTAIL.n471 VTAIL.n449 0.155672
R1293 VTAIL.n471 VTAIL.n470 0.155672
R1294 VTAIL.n470 VTAIL.n454 0.155672
R1295 VTAIL.n463 VTAIL.n454 0.155672
R1296 VTAIL.n463 VTAIL.n462 0.155672
R1297 VTAIL.n421 VTAIL.n319 0.155672
R1298 VTAIL.n414 VTAIL.n319 0.155672
R1299 VTAIL.n414 VTAIL.n413 0.155672
R1300 VTAIL.n413 VTAIL.n323 0.155672
R1301 VTAIL.n406 VTAIL.n323 0.155672
R1302 VTAIL.n406 VTAIL.n405 0.155672
R1303 VTAIL.n405 VTAIL.n327 0.155672
R1304 VTAIL.n398 VTAIL.n327 0.155672
R1305 VTAIL.n398 VTAIL.n397 0.155672
R1306 VTAIL.n397 VTAIL.n331 0.155672
R1307 VTAIL.n390 VTAIL.n331 0.155672
R1308 VTAIL.n390 VTAIL.n389 0.155672
R1309 VTAIL.n389 VTAIL.n335 0.155672
R1310 VTAIL.n382 VTAIL.n335 0.155672
R1311 VTAIL.n382 VTAIL.n381 0.155672
R1312 VTAIL.n381 VTAIL.n339 0.155672
R1313 VTAIL.n373 VTAIL.n339 0.155672
R1314 VTAIL.n373 VTAIL.n372 0.155672
R1315 VTAIL.n372 VTAIL.n343 0.155672
R1316 VTAIL.n365 VTAIL.n343 0.155672
R1317 VTAIL.n365 VTAIL.n364 0.155672
R1318 VTAIL.n364 VTAIL.n348 0.155672
R1319 VTAIL.n357 VTAIL.n348 0.155672
R1320 VTAIL.n357 VTAIL.n356 0.155672
R1321 B.n623 B.n622 585
R1322 B.n624 B.n95 585
R1323 B.n626 B.n625 585
R1324 B.n627 B.n94 585
R1325 B.n629 B.n628 585
R1326 B.n630 B.n93 585
R1327 B.n632 B.n631 585
R1328 B.n633 B.n92 585
R1329 B.n635 B.n634 585
R1330 B.n636 B.n91 585
R1331 B.n638 B.n637 585
R1332 B.n639 B.n90 585
R1333 B.n641 B.n640 585
R1334 B.n642 B.n89 585
R1335 B.n644 B.n643 585
R1336 B.n645 B.n88 585
R1337 B.n647 B.n646 585
R1338 B.n648 B.n87 585
R1339 B.n650 B.n649 585
R1340 B.n651 B.n86 585
R1341 B.n653 B.n652 585
R1342 B.n654 B.n85 585
R1343 B.n656 B.n655 585
R1344 B.n657 B.n84 585
R1345 B.n659 B.n658 585
R1346 B.n660 B.n83 585
R1347 B.n662 B.n661 585
R1348 B.n663 B.n82 585
R1349 B.n665 B.n664 585
R1350 B.n666 B.n81 585
R1351 B.n668 B.n667 585
R1352 B.n669 B.n80 585
R1353 B.n671 B.n670 585
R1354 B.n672 B.n79 585
R1355 B.n674 B.n673 585
R1356 B.n675 B.n78 585
R1357 B.n677 B.n676 585
R1358 B.n678 B.n77 585
R1359 B.n680 B.n679 585
R1360 B.n681 B.n76 585
R1361 B.n683 B.n682 585
R1362 B.n684 B.n75 585
R1363 B.n686 B.n685 585
R1364 B.n687 B.n74 585
R1365 B.n689 B.n688 585
R1366 B.n690 B.n73 585
R1367 B.n692 B.n691 585
R1368 B.n693 B.n72 585
R1369 B.n695 B.n694 585
R1370 B.n696 B.n71 585
R1371 B.n698 B.n697 585
R1372 B.n699 B.n70 585
R1373 B.n701 B.n700 585
R1374 B.n702 B.n69 585
R1375 B.n704 B.n703 585
R1376 B.n705 B.n68 585
R1377 B.n707 B.n706 585
R1378 B.n708 B.n67 585
R1379 B.n710 B.n709 585
R1380 B.n711 B.n66 585
R1381 B.n713 B.n712 585
R1382 B.n714 B.n65 585
R1383 B.n716 B.n715 585
R1384 B.n717 B.n62 585
R1385 B.n720 B.n719 585
R1386 B.n721 B.n61 585
R1387 B.n723 B.n722 585
R1388 B.n724 B.n60 585
R1389 B.n726 B.n725 585
R1390 B.n727 B.n59 585
R1391 B.n729 B.n728 585
R1392 B.n730 B.n55 585
R1393 B.n732 B.n731 585
R1394 B.n733 B.n54 585
R1395 B.n735 B.n734 585
R1396 B.n736 B.n53 585
R1397 B.n738 B.n737 585
R1398 B.n739 B.n52 585
R1399 B.n741 B.n740 585
R1400 B.n742 B.n51 585
R1401 B.n744 B.n743 585
R1402 B.n745 B.n50 585
R1403 B.n747 B.n746 585
R1404 B.n748 B.n49 585
R1405 B.n750 B.n749 585
R1406 B.n751 B.n48 585
R1407 B.n753 B.n752 585
R1408 B.n754 B.n47 585
R1409 B.n756 B.n755 585
R1410 B.n757 B.n46 585
R1411 B.n759 B.n758 585
R1412 B.n760 B.n45 585
R1413 B.n762 B.n761 585
R1414 B.n763 B.n44 585
R1415 B.n765 B.n764 585
R1416 B.n766 B.n43 585
R1417 B.n768 B.n767 585
R1418 B.n769 B.n42 585
R1419 B.n771 B.n770 585
R1420 B.n772 B.n41 585
R1421 B.n774 B.n773 585
R1422 B.n775 B.n40 585
R1423 B.n777 B.n776 585
R1424 B.n778 B.n39 585
R1425 B.n780 B.n779 585
R1426 B.n781 B.n38 585
R1427 B.n783 B.n782 585
R1428 B.n784 B.n37 585
R1429 B.n786 B.n785 585
R1430 B.n787 B.n36 585
R1431 B.n789 B.n788 585
R1432 B.n790 B.n35 585
R1433 B.n792 B.n791 585
R1434 B.n793 B.n34 585
R1435 B.n795 B.n794 585
R1436 B.n796 B.n33 585
R1437 B.n798 B.n797 585
R1438 B.n799 B.n32 585
R1439 B.n801 B.n800 585
R1440 B.n802 B.n31 585
R1441 B.n804 B.n803 585
R1442 B.n805 B.n30 585
R1443 B.n807 B.n806 585
R1444 B.n808 B.n29 585
R1445 B.n810 B.n809 585
R1446 B.n811 B.n28 585
R1447 B.n813 B.n812 585
R1448 B.n814 B.n27 585
R1449 B.n816 B.n815 585
R1450 B.n817 B.n26 585
R1451 B.n819 B.n818 585
R1452 B.n820 B.n25 585
R1453 B.n822 B.n821 585
R1454 B.n823 B.n24 585
R1455 B.n825 B.n824 585
R1456 B.n826 B.n23 585
R1457 B.n828 B.n827 585
R1458 B.n621 B.n96 585
R1459 B.n620 B.n619 585
R1460 B.n618 B.n97 585
R1461 B.n617 B.n616 585
R1462 B.n615 B.n98 585
R1463 B.n614 B.n613 585
R1464 B.n612 B.n99 585
R1465 B.n611 B.n610 585
R1466 B.n609 B.n100 585
R1467 B.n608 B.n607 585
R1468 B.n606 B.n101 585
R1469 B.n605 B.n604 585
R1470 B.n603 B.n102 585
R1471 B.n602 B.n601 585
R1472 B.n600 B.n103 585
R1473 B.n599 B.n598 585
R1474 B.n597 B.n104 585
R1475 B.n596 B.n595 585
R1476 B.n594 B.n105 585
R1477 B.n593 B.n592 585
R1478 B.n591 B.n106 585
R1479 B.n590 B.n589 585
R1480 B.n588 B.n107 585
R1481 B.n587 B.n586 585
R1482 B.n585 B.n108 585
R1483 B.n584 B.n583 585
R1484 B.n582 B.n109 585
R1485 B.n581 B.n580 585
R1486 B.n579 B.n110 585
R1487 B.n578 B.n577 585
R1488 B.n576 B.n111 585
R1489 B.n575 B.n574 585
R1490 B.n573 B.n112 585
R1491 B.n572 B.n571 585
R1492 B.n570 B.n113 585
R1493 B.n569 B.n568 585
R1494 B.n567 B.n114 585
R1495 B.n566 B.n565 585
R1496 B.n564 B.n115 585
R1497 B.n563 B.n562 585
R1498 B.n561 B.n116 585
R1499 B.n560 B.n559 585
R1500 B.n558 B.n117 585
R1501 B.n557 B.n556 585
R1502 B.n555 B.n118 585
R1503 B.n554 B.n553 585
R1504 B.n552 B.n119 585
R1505 B.n551 B.n550 585
R1506 B.n549 B.n120 585
R1507 B.n548 B.n547 585
R1508 B.n546 B.n121 585
R1509 B.n545 B.n544 585
R1510 B.n543 B.n122 585
R1511 B.n542 B.n541 585
R1512 B.n540 B.n123 585
R1513 B.n539 B.n538 585
R1514 B.n537 B.n124 585
R1515 B.n536 B.n535 585
R1516 B.n534 B.n125 585
R1517 B.n533 B.n532 585
R1518 B.n531 B.n126 585
R1519 B.n530 B.n529 585
R1520 B.n528 B.n127 585
R1521 B.n527 B.n526 585
R1522 B.n525 B.n128 585
R1523 B.n524 B.n523 585
R1524 B.n522 B.n129 585
R1525 B.n521 B.n520 585
R1526 B.n519 B.n130 585
R1527 B.n518 B.n517 585
R1528 B.n516 B.n131 585
R1529 B.n515 B.n514 585
R1530 B.n513 B.n132 585
R1531 B.n512 B.n511 585
R1532 B.n510 B.n133 585
R1533 B.n509 B.n508 585
R1534 B.n507 B.n134 585
R1535 B.n506 B.n505 585
R1536 B.n504 B.n135 585
R1537 B.n503 B.n502 585
R1538 B.n501 B.n136 585
R1539 B.n500 B.n499 585
R1540 B.n498 B.n137 585
R1541 B.n289 B.n288 585
R1542 B.n290 B.n207 585
R1543 B.n292 B.n291 585
R1544 B.n293 B.n206 585
R1545 B.n295 B.n294 585
R1546 B.n296 B.n205 585
R1547 B.n298 B.n297 585
R1548 B.n299 B.n204 585
R1549 B.n301 B.n300 585
R1550 B.n302 B.n203 585
R1551 B.n304 B.n303 585
R1552 B.n305 B.n202 585
R1553 B.n307 B.n306 585
R1554 B.n308 B.n201 585
R1555 B.n310 B.n309 585
R1556 B.n311 B.n200 585
R1557 B.n313 B.n312 585
R1558 B.n314 B.n199 585
R1559 B.n316 B.n315 585
R1560 B.n317 B.n198 585
R1561 B.n319 B.n318 585
R1562 B.n320 B.n197 585
R1563 B.n322 B.n321 585
R1564 B.n323 B.n196 585
R1565 B.n325 B.n324 585
R1566 B.n326 B.n195 585
R1567 B.n328 B.n327 585
R1568 B.n329 B.n194 585
R1569 B.n331 B.n330 585
R1570 B.n332 B.n193 585
R1571 B.n334 B.n333 585
R1572 B.n335 B.n192 585
R1573 B.n337 B.n336 585
R1574 B.n338 B.n191 585
R1575 B.n340 B.n339 585
R1576 B.n341 B.n190 585
R1577 B.n343 B.n342 585
R1578 B.n344 B.n189 585
R1579 B.n346 B.n345 585
R1580 B.n347 B.n188 585
R1581 B.n349 B.n348 585
R1582 B.n350 B.n187 585
R1583 B.n352 B.n351 585
R1584 B.n353 B.n186 585
R1585 B.n355 B.n354 585
R1586 B.n356 B.n185 585
R1587 B.n358 B.n357 585
R1588 B.n359 B.n184 585
R1589 B.n361 B.n360 585
R1590 B.n362 B.n183 585
R1591 B.n364 B.n363 585
R1592 B.n365 B.n182 585
R1593 B.n367 B.n366 585
R1594 B.n368 B.n181 585
R1595 B.n370 B.n369 585
R1596 B.n371 B.n180 585
R1597 B.n373 B.n372 585
R1598 B.n374 B.n179 585
R1599 B.n376 B.n375 585
R1600 B.n377 B.n178 585
R1601 B.n379 B.n378 585
R1602 B.n380 B.n177 585
R1603 B.n382 B.n381 585
R1604 B.n383 B.n174 585
R1605 B.n386 B.n385 585
R1606 B.n387 B.n173 585
R1607 B.n389 B.n388 585
R1608 B.n390 B.n172 585
R1609 B.n392 B.n391 585
R1610 B.n393 B.n171 585
R1611 B.n395 B.n394 585
R1612 B.n396 B.n170 585
R1613 B.n401 B.n400 585
R1614 B.n402 B.n169 585
R1615 B.n404 B.n403 585
R1616 B.n405 B.n168 585
R1617 B.n407 B.n406 585
R1618 B.n408 B.n167 585
R1619 B.n410 B.n409 585
R1620 B.n411 B.n166 585
R1621 B.n413 B.n412 585
R1622 B.n414 B.n165 585
R1623 B.n416 B.n415 585
R1624 B.n417 B.n164 585
R1625 B.n419 B.n418 585
R1626 B.n420 B.n163 585
R1627 B.n422 B.n421 585
R1628 B.n423 B.n162 585
R1629 B.n425 B.n424 585
R1630 B.n426 B.n161 585
R1631 B.n428 B.n427 585
R1632 B.n429 B.n160 585
R1633 B.n431 B.n430 585
R1634 B.n432 B.n159 585
R1635 B.n434 B.n433 585
R1636 B.n435 B.n158 585
R1637 B.n437 B.n436 585
R1638 B.n438 B.n157 585
R1639 B.n440 B.n439 585
R1640 B.n441 B.n156 585
R1641 B.n443 B.n442 585
R1642 B.n444 B.n155 585
R1643 B.n446 B.n445 585
R1644 B.n447 B.n154 585
R1645 B.n449 B.n448 585
R1646 B.n450 B.n153 585
R1647 B.n452 B.n451 585
R1648 B.n453 B.n152 585
R1649 B.n455 B.n454 585
R1650 B.n456 B.n151 585
R1651 B.n458 B.n457 585
R1652 B.n459 B.n150 585
R1653 B.n461 B.n460 585
R1654 B.n462 B.n149 585
R1655 B.n464 B.n463 585
R1656 B.n465 B.n148 585
R1657 B.n467 B.n466 585
R1658 B.n468 B.n147 585
R1659 B.n470 B.n469 585
R1660 B.n471 B.n146 585
R1661 B.n473 B.n472 585
R1662 B.n474 B.n145 585
R1663 B.n476 B.n475 585
R1664 B.n477 B.n144 585
R1665 B.n479 B.n478 585
R1666 B.n480 B.n143 585
R1667 B.n482 B.n481 585
R1668 B.n483 B.n142 585
R1669 B.n485 B.n484 585
R1670 B.n486 B.n141 585
R1671 B.n488 B.n487 585
R1672 B.n489 B.n140 585
R1673 B.n491 B.n490 585
R1674 B.n492 B.n139 585
R1675 B.n494 B.n493 585
R1676 B.n495 B.n138 585
R1677 B.n497 B.n496 585
R1678 B.n287 B.n208 585
R1679 B.n286 B.n285 585
R1680 B.n284 B.n209 585
R1681 B.n283 B.n282 585
R1682 B.n281 B.n210 585
R1683 B.n280 B.n279 585
R1684 B.n278 B.n211 585
R1685 B.n277 B.n276 585
R1686 B.n275 B.n212 585
R1687 B.n274 B.n273 585
R1688 B.n272 B.n213 585
R1689 B.n271 B.n270 585
R1690 B.n269 B.n214 585
R1691 B.n268 B.n267 585
R1692 B.n266 B.n215 585
R1693 B.n265 B.n264 585
R1694 B.n263 B.n216 585
R1695 B.n262 B.n261 585
R1696 B.n260 B.n217 585
R1697 B.n259 B.n258 585
R1698 B.n257 B.n218 585
R1699 B.n256 B.n255 585
R1700 B.n254 B.n219 585
R1701 B.n253 B.n252 585
R1702 B.n251 B.n220 585
R1703 B.n250 B.n249 585
R1704 B.n248 B.n221 585
R1705 B.n247 B.n246 585
R1706 B.n245 B.n222 585
R1707 B.n244 B.n243 585
R1708 B.n242 B.n223 585
R1709 B.n241 B.n240 585
R1710 B.n239 B.n224 585
R1711 B.n238 B.n237 585
R1712 B.n236 B.n225 585
R1713 B.n235 B.n234 585
R1714 B.n233 B.n226 585
R1715 B.n232 B.n231 585
R1716 B.n230 B.n227 585
R1717 B.n229 B.n228 585
R1718 B.n2 B.n0 585
R1719 B.n889 B.n1 585
R1720 B.n888 B.n887 585
R1721 B.n886 B.n3 585
R1722 B.n885 B.n884 585
R1723 B.n883 B.n4 585
R1724 B.n882 B.n881 585
R1725 B.n880 B.n5 585
R1726 B.n879 B.n878 585
R1727 B.n877 B.n6 585
R1728 B.n876 B.n875 585
R1729 B.n874 B.n7 585
R1730 B.n873 B.n872 585
R1731 B.n871 B.n8 585
R1732 B.n870 B.n869 585
R1733 B.n868 B.n9 585
R1734 B.n867 B.n866 585
R1735 B.n865 B.n10 585
R1736 B.n864 B.n863 585
R1737 B.n862 B.n11 585
R1738 B.n861 B.n860 585
R1739 B.n859 B.n12 585
R1740 B.n858 B.n857 585
R1741 B.n856 B.n13 585
R1742 B.n855 B.n854 585
R1743 B.n853 B.n14 585
R1744 B.n852 B.n851 585
R1745 B.n850 B.n15 585
R1746 B.n849 B.n848 585
R1747 B.n847 B.n16 585
R1748 B.n846 B.n845 585
R1749 B.n844 B.n17 585
R1750 B.n843 B.n842 585
R1751 B.n841 B.n18 585
R1752 B.n840 B.n839 585
R1753 B.n838 B.n19 585
R1754 B.n837 B.n836 585
R1755 B.n835 B.n20 585
R1756 B.n834 B.n833 585
R1757 B.n832 B.n21 585
R1758 B.n831 B.n830 585
R1759 B.n829 B.n22 585
R1760 B.n891 B.n890 585
R1761 B.n397 B.t2 582.404
R1762 B.n63 B.t7 582.404
R1763 B.n175 B.t5 582.404
R1764 B.n56 B.t10 582.404
R1765 B.n398 B.t1 509.87
R1766 B.n64 B.t8 509.87
R1767 B.n176 B.t4 509.87
R1768 B.n57 B.t11 509.87
R1769 B.n289 B.n208 492.5
R1770 B.n829 B.n828 492.5
R1771 B.n498 B.n497 492.5
R1772 B.n623 B.n96 492.5
R1773 B.n397 B.t0 346.543
R1774 B.n175 B.t3 346.543
R1775 B.n56 B.t9 346.543
R1776 B.n63 B.t6 346.543
R1777 B.n285 B.n208 163.367
R1778 B.n285 B.n284 163.367
R1779 B.n284 B.n283 163.367
R1780 B.n283 B.n210 163.367
R1781 B.n279 B.n210 163.367
R1782 B.n279 B.n278 163.367
R1783 B.n278 B.n277 163.367
R1784 B.n277 B.n212 163.367
R1785 B.n273 B.n212 163.367
R1786 B.n273 B.n272 163.367
R1787 B.n272 B.n271 163.367
R1788 B.n271 B.n214 163.367
R1789 B.n267 B.n214 163.367
R1790 B.n267 B.n266 163.367
R1791 B.n266 B.n265 163.367
R1792 B.n265 B.n216 163.367
R1793 B.n261 B.n216 163.367
R1794 B.n261 B.n260 163.367
R1795 B.n260 B.n259 163.367
R1796 B.n259 B.n218 163.367
R1797 B.n255 B.n218 163.367
R1798 B.n255 B.n254 163.367
R1799 B.n254 B.n253 163.367
R1800 B.n253 B.n220 163.367
R1801 B.n249 B.n220 163.367
R1802 B.n249 B.n248 163.367
R1803 B.n248 B.n247 163.367
R1804 B.n247 B.n222 163.367
R1805 B.n243 B.n222 163.367
R1806 B.n243 B.n242 163.367
R1807 B.n242 B.n241 163.367
R1808 B.n241 B.n224 163.367
R1809 B.n237 B.n224 163.367
R1810 B.n237 B.n236 163.367
R1811 B.n236 B.n235 163.367
R1812 B.n235 B.n226 163.367
R1813 B.n231 B.n226 163.367
R1814 B.n231 B.n230 163.367
R1815 B.n230 B.n229 163.367
R1816 B.n229 B.n2 163.367
R1817 B.n890 B.n2 163.367
R1818 B.n890 B.n889 163.367
R1819 B.n889 B.n888 163.367
R1820 B.n888 B.n3 163.367
R1821 B.n884 B.n3 163.367
R1822 B.n884 B.n883 163.367
R1823 B.n883 B.n882 163.367
R1824 B.n882 B.n5 163.367
R1825 B.n878 B.n5 163.367
R1826 B.n878 B.n877 163.367
R1827 B.n877 B.n876 163.367
R1828 B.n876 B.n7 163.367
R1829 B.n872 B.n7 163.367
R1830 B.n872 B.n871 163.367
R1831 B.n871 B.n870 163.367
R1832 B.n870 B.n9 163.367
R1833 B.n866 B.n9 163.367
R1834 B.n866 B.n865 163.367
R1835 B.n865 B.n864 163.367
R1836 B.n864 B.n11 163.367
R1837 B.n860 B.n11 163.367
R1838 B.n860 B.n859 163.367
R1839 B.n859 B.n858 163.367
R1840 B.n858 B.n13 163.367
R1841 B.n854 B.n13 163.367
R1842 B.n854 B.n853 163.367
R1843 B.n853 B.n852 163.367
R1844 B.n852 B.n15 163.367
R1845 B.n848 B.n15 163.367
R1846 B.n848 B.n847 163.367
R1847 B.n847 B.n846 163.367
R1848 B.n846 B.n17 163.367
R1849 B.n842 B.n17 163.367
R1850 B.n842 B.n841 163.367
R1851 B.n841 B.n840 163.367
R1852 B.n840 B.n19 163.367
R1853 B.n836 B.n19 163.367
R1854 B.n836 B.n835 163.367
R1855 B.n835 B.n834 163.367
R1856 B.n834 B.n21 163.367
R1857 B.n830 B.n21 163.367
R1858 B.n830 B.n829 163.367
R1859 B.n290 B.n289 163.367
R1860 B.n291 B.n290 163.367
R1861 B.n291 B.n206 163.367
R1862 B.n295 B.n206 163.367
R1863 B.n296 B.n295 163.367
R1864 B.n297 B.n296 163.367
R1865 B.n297 B.n204 163.367
R1866 B.n301 B.n204 163.367
R1867 B.n302 B.n301 163.367
R1868 B.n303 B.n302 163.367
R1869 B.n303 B.n202 163.367
R1870 B.n307 B.n202 163.367
R1871 B.n308 B.n307 163.367
R1872 B.n309 B.n308 163.367
R1873 B.n309 B.n200 163.367
R1874 B.n313 B.n200 163.367
R1875 B.n314 B.n313 163.367
R1876 B.n315 B.n314 163.367
R1877 B.n315 B.n198 163.367
R1878 B.n319 B.n198 163.367
R1879 B.n320 B.n319 163.367
R1880 B.n321 B.n320 163.367
R1881 B.n321 B.n196 163.367
R1882 B.n325 B.n196 163.367
R1883 B.n326 B.n325 163.367
R1884 B.n327 B.n326 163.367
R1885 B.n327 B.n194 163.367
R1886 B.n331 B.n194 163.367
R1887 B.n332 B.n331 163.367
R1888 B.n333 B.n332 163.367
R1889 B.n333 B.n192 163.367
R1890 B.n337 B.n192 163.367
R1891 B.n338 B.n337 163.367
R1892 B.n339 B.n338 163.367
R1893 B.n339 B.n190 163.367
R1894 B.n343 B.n190 163.367
R1895 B.n344 B.n343 163.367
R1896 B.n345 B.n344 163.367
R1897 B.n345 B.n188 163.367
R1898 B.n349 B.n188 163.367
R1899 B.n350 B.n349 163.367
R1900 B.n351 B.n350 163.367
R1901 B.n351 B.n186 163.367
R1902 B.n355 B.n186 163.367
R1903 B.n356 B.n355 163.367
R1904 B.n357 B.n356 163.367
R1905 B.n357 B.n184 163.367
R1906 B.n361 B.n184 163.367
R1907 B.n362 B.n361 163.367
R1908 B.n363 B.n362 163.367
R1909 B.n363 B.n182 163.367
R1910 B.n367 B.n182 163.367
R1911 B.n368 B.n367 163.367
R1912 B.n369 B.n368 163.367
R1913 B.n369 B.n180 163.367
R1914 B.n373 B.n180 163.367
R1915 B.n374 B.n373 163.367
R1916 B.n375 B.n374 163.367
R1917 B.n375 B.n178 163.367
R1918 B.n379 B.n178 163.367
R1919 B.n380 B.n379 163.367
R1920 B.n381 B.n380 163.367
R1921 B.n381 B.n174 163.367
R1922 B.n386 B.n174 163.367
R1923 B.n387 B.n386 163.367
R1924 B.n388 B.n387 163.367
R1925 B.n388 B.n172 163.367
R1926 B.n392 B.n172 163.367
R1927 B.n393 B.n392 163.367
R1928 B.n394 B.n393 163.367
R1929 B.n394 B.n170 163.367
R1930 B.n401 B.n170 163.367
R1931 B.n402 B.n401 163.367
R1932 B.n403 B.n402 163.367
R1933 B.n403 B.n168 163.367
R1934 B.n407 B.n168 163.367
R1935 B.n408 B.n407 163.367
R1936 B.n409 B.n408 163.367
R1937 B.n409 B.n166 163.367
R1938 B.n413 B.n166 163.367
R1939 B.n414 B.n413 163.367
R1940 B.n415 B.n414 163.367
R1941 B.n415 B.n164 163.367
R1942 B.n419 B.n164 163.367
R1943 B.n420 B.n419 163.367
R1944 B.n421 B.n420 163.367
R1945 B.n421 B.n162 163.367
R1946 B.n425 B.n162 163.367
R1947 B.n426 B.n425 163.367
R1948 B.n427 B.n426 163.367
R1949 B.n427 B.n160 163.367
R1950 B.n431 B.n160 163.367
R1951 B.n432 B.n431 163.367
R1952 B.n433 B.n432 163.367
R1953 B.n433 B.n158 163.367
R1954 B.n437 B.n158 163.367
R1955 B.n438 B.n437 163.367
R1956 B.n439 B.n438 163.367
R1957 B.n439 B.n156 163.367
R1958 B.n443 B.n156 163.367
R1959 B.n444 B.n443 163.367
R1960 B.n445 B.n444 163.367
R1961 B.n445 B.n154 163.367
R1962 B.n449 B.n154 163.367
R1963 B.n450 B.n449 163.367
R1964 B.n451 B.n450 163.367
R1965 B.n451 B.n152 163.367
R1966 B.n455 B.n152 163.367
R1967 B.n456 B.n455 163.367
R1968 B.n457 B.n456 163.367
R1969 B.n457 B.n150 163.367
R1970 B.n461 B.n150 163.367
R1971 B.n462 B.n461 163.367
R1972 B.n463 B.n462 163.367
R1973 B.n463 B.n148 163.367
R1974 B.n467 B.n148 163.367
R1975 B.n468 B.n467 163.367
R1976 B.n469 B.n468 163.367
R1977 B.n469 B.n146 163.367
R1978 B.n473 B.n146 163.367
R1979 B.n474 B.n473 163.367
R1980 B.n475 B.n474 163.367
R1981 B.n475 B.n144 163.367
R1982 B.n479 B.n144 163.367
R1983 B.n480 B.n479 163.367
R1984 B.n481 B.n480 163.367
R1985 B.n481 B.n142 163.367
R1986 B.n485 B.n142 163.367
R1987 B.n486 B.n485 163.367
R1988 B.n487 B.n486 163.367
R1989 B.n487 B.n140 163.367
R1990 B.n491 B.n140 163.367
R1991 B.n492 B.n491 163.367
R1992 B.n493 B.n492 163.367
R1993 B.n493 B.n138 163.367
R1994 B.n497 B.n138 163.367
R1995 B.n499 B.n498 163.367
R1996 B.n499 B.n136 163.367
R1997 B.n503 B.n136 163.367
R1998 B.n504 B.n503 163.367
R1999 B.n505 B.n504 163.367
R2000 B.n505 B.n134 163.367
R2001 B.n509 B.n134 163.367
R2002 B.n510 B.n509 163.367
R2003 B.n511 B.n510 163.367
R2004 B.n511 B.n132 163.367
R2005 B.n515 B.n132 163.367
R2006 B.n516 B.n515 163.367
R2007 B.n517 B.n516 163.367
R2008 B.n517 B.n130 163.367
R2009 B.n521 B.n130 163.367
R2010 B.n522 B.n521 163.367
R2011 B.n523 B.n522 163.367
R2012 B.n523 B.n128 163.367
R2013 B.n527 B.n128 163.367
R2014 B.n528 B.n527 163.367
R2015 B.n529 B.n528 163.367
R2016 B.n529 B.n126 163.367
R2017 B.n533 B.n126 163.367
R2018 B.n534 B.n533 163.367
R2019 B.n535 B.n534 163.367
R2020 B.n535 B.n124 163.367
R2021 B.n539 B.n124 163.367
R2022 B.n540 B.n539 163.367
R2023 B.n541 B.n540 163.367
R2024 B.n541 B.n122 163.367
R2025 B.n545 B.n122 163.367
R2026 B.n546 B.n545 163.367
R2027 B.n547 B.n546 163.367
R2028 B.n547 B.n120 163.367
R2029 B.n551 B.n120 163.367
R2030 B.n552 B.n551 163.367
R2031 B.n553 B.n552 163.367
R2032 B.n553 B.n118 163.367
R2033 B.n557 B.n118 163.367
R2034 B.n558 B.n557 163.367
R2035 B.n559 B.n558 163.367
R2036 B.n559 B.n116 163.367
R2037 B.n563 B.n116 163.367
R2038 B.n564 B.n563 163.367
R2039 B.n565 B.n564 163.367
R2040 B.n565 B.n114 163.367
R2041 B.n569 B.n114 163.367
R2042 B.n570 B.n569 163.367
R2043 B.n571 B.n570 163.367
R2044 B.n571 B.n112 163.367
R2045 B.n575 B.n112 163.367
R2046 B.n576 B.n575 163.367
R2047 B.n577 B.n576 163.367
R2048 B.n577 B.n110 163.367
R2049 B.n581 B.n110 163.367
R2050 B.n582 B.n581 163.367
R2051 B.n583 B.n582 163.367
R2052 B.n583 B.n108 163.367
R2053 B.n587 B.n108 163.367
R2054 B.n588 B.n587 163.367
R2055 B.n589 B.n588 163.367
R2056 B.n589 B.n106 163.367
R2057 B.n593 B.n106 163.367
R2058 B.n594 B.n593 163.367
R2059 B.n595 B.n594 163.367
R2060 B.n595 B.n104 163.367
R2061 B.n599 B.n104 163.367
R2062 B.n600 B.n599 163.367
R2063 B.n601 B.n600 163.367
R2064 B.n601 B.n102 163.367
R2065 B.n605 B.n102 163.367
R2066 B.n606 B.n605 163.367
R2067 B.n607 B.n606 163.367
R2068 B.n607 B.n100 163.367
R2069 B.n611 B.n100 163.367
R2070 B.n612 B.n611 163.367
R2071 B.n613 B.n612 163.367
R2072 B.n613 B.n98 163.367
R2073 B.n617 B.n98 163.367
R2074 B.n618 B.n617 163.367
R2075 B.n619 B.n618 163.367
R2076 B.n619 B.n96 163.367
R2077 B.n828 B.n23 163.367
R2078 B.n824 B.n23 163.367
R2079 B.n824 B.n823 163.367
R2080 B.n823 B.n822 163.367
R2081 B.n822 B.n25 163.367
R2082 B.n818 B.n25 163.367
R2083 B.n818 B.n817 163.367
R2084 B.n817 B.n816 163.367
R2085 B.n816 B.n27 163.367
R2086 B.n812 B.n27 163.367
R2087 B.n812 B.n811 163.367
R2088 B.n811 B.n810 163.367
R2089 B.n810 B.n29 163.367
R2090 B.n806 B.n29 163.367
R2091 B.n806 B.n805 163.367
R2092 B.n805 B.n804 163.367
R2093 B.n804 B.n31 163.367
R2094 B.n800 B.n31 163.367
R2095 B.n800 B.n799 163.367
R2096 B.n799 B.n798 163.367
R2097 B.n798 B.n33 163.367
R2098 B.n794 B.n33 163.367
R2099 B.n794 B.n793 163.367
R2100 B.n793 B.n792 163.367
R2101 B.n792 B.n35 163.367
R2102 B.n788 B.n35 163.367
R2103 B.n788 B.n787 163.367
R2104 B.n787 B.n786 163.367
R2105 B.n786 B.n37 163.367
R2106 B.n782 B.n37 163.367
R2107 B.n782 B.n781 163.367
R2108 B.n781 B.n780 163.367
R2109 B.n780 B.n39 163.367
R2110 B.n776 B.n39 163.367
R2111 B.n776 B.n775 163.367
R2112 B.n775 B.n774 163.367
R2113 B.n774 B.n41 163.367
R2114 B.n770 B.n41 163.367
R2115 B.n770 B.n769 163.367
R2116 B.n769 B.n768 163.367
R2117 B.n768 B.n43 163.367
R2118 B.n764 B.n43 163.367
R2119 B.n764 B.n763 163.367
R2120 B.n763 B.n762 163.367
R2121 B.n762 B.n45 163.367
R2122 B.n758 B.n45 163.367
R2123 B.n758 B.n757 163.367
R2124 B.n757 B.n756 163.367
R2125 B.n756 B.n47 163.367
R2126 B.n752 B.n47 163.367
R2127 B.n752 B.n751 163.367
R2128 B.n751 B.n750 163.367
R2129 B.n750 B.n49 163.367
R2130 B.n746 B.n49 163.367
R2131 B.n746 B.n745 163.367
R2132 B.n745 B.n744 163.367
R2133 B.n744 B.n51 163.367
R2134 B.n740 B.n51 163.367
R2135 B.n740 B.n739 163.367
R2136 B.n739 B.n738 163.367
R2137 B.n738 B.n53 163.367
R2138 B.n734 B.n53 163.367
R2139 B.n734 B.n733 163.367
R2140 B.n733 B.n732 163.367
R2141 B.n732 B.n55 163.367
R2142 B.n728 B.n55 163.367
R2143 B.n728 B.n727 163.367
R2144 B.n727 B.n726 163.367
R2145 B.n726 B.n60 163.367
R2146 B.n722 B.n60 163.367
R2147 B.n722 B.n721 163.367
R2148 B.n721 B.n720 163.367
R2149 B.n720 B.n62 163.367
R2150 B.n715 B.n62 163.367
R2151 B.n715 B.n714 163.367
R2152 B.n714 B.n713 163.367
R2153 B.n713 B.n66 163.367
R2154 B.n709 B.n66 163.367
R2155 B.n709 B.n708 163.367
R2156 B.n708 B.n707 163.367
R2157 B.n707 B.n68 163.367
R2158 B.n703 B.n68 163.367
R2159 B.n703 B.n702 163.367
R2160 B.n702 B.n701 163.367
R2161 B.n701 B.n70 163.367
R2162 B.n697 B.n70 163.367
R2163 B.n697 B.n696 163.367
R2164 B.n696 B.n695 163.367
R2165 B.n695 B.n72 163.367
R2166 B.n691 B.n72 163.367
R2167 B.n691 B.n690 163.367
R2168 B.n690 B.n689 163.367
R2169 B.n689 B.n74 163.367
R2170 B.n685 B.n74 163.367
R2171 B.n685 B.n684 163.367
R2172 B.n684 B.n683 163.367
R2173 B.n683 B.n76 163.367
R2174 B.n679 B.n76 163.367
R2175 B.n679 B.n678 163.367
R2176 B.n678 B.n677 163.367
R2177 B.n677 B.n78 163.367
R2178 B.n673 B.n78 163.367
R2179 B.n673 B.n672 163.367
R2180 B.n672 B.n671 163.367
R2181 B.n671 B.n80 163.367
R2182 B.n667 B.n80 163.367
R2183 B.n667 B.n666 163.367
R2184 B.n666 B.n665 163.367
R2185 B.n665 B.n82 163.367
R2186 B.n661 B.n82 163.367
R2187 B.n661 B.n660 163.367
R2188 B.n660 B.n659 163.367
R2189 B.n659 B.n84 163.367
R2190 B.n655 B.n84 163.367
R2191 B.n655 B.n654 163.367
R2192 B.n654 B.n653 163.367
R2193 B.n653 B.n86 163.367
R2194 B.n649 B.n86 163.367
R2195 B.n649 B.n648 163.367
R2196 B.n648 B.n647 163.367
R2197 B.n647 B.n88 163.367
R2198 B.n643 B.n88 163.367
R2199 B.n643 B.n642 163.367
R2200 B.n642 B.n641 163.367
R2201 B.n641 B.n90 163.367
R2202 B.n637 B.n90 163.367
R2203 B.n637 B.n636 163.367
R2204 B.n636 B.n635 163.367
R2205 B.n635 B.n92 163.367
R2206 B.n631 B.n92 163.367
R2207 B.n631 B.n630 163.367
R2208 B.n630 B.n629 163.367
R2209 B.n629 B.n94 163.367
R2210 B.n625 B.n94 163.367
R2211 B.n625 B.n624 163.367
R2212 B.n624 B.n623 163.367
R2213 B.n398 B.n397 72.5338
R2214 B.n176 B.n175 72.5338
R2215 B.n57 B.n56 72.5338
R2216 B.n64 B.n63 72.5338
R2217 B.n399 B.n398 59.5399
R2218 B.n384 B.n176 59.5399
R2219 B.n58 B.n57 59.5399
R2220 B.n718 B.n64 59.5399
R2221 B.n827 B.n22 32.0005
R2222 B.n622 B.n621 32.0005
R2223 B.n496 B.n137 32.0005
R2224 B.n288 B.n287 32.0005
R2225 B B.n891 18.0485
R2226 B.n827 B.n826 10.6151
R2227 B.n826 B.n825 10.6151
R2228 B.n825 B.n24 10.6151
R2229 B.n821 B.n24 10.6151
R2230 B.n821 B.n820 10.6151
R2231 B.n820 B.n819 10.6151
R2232 B.n819 B.n26 10.6151
R2233 B.n815 B.n26 10.6151
R2234 B.n815 B.n814 10.6151
R2235 B.n814 B.n813 10.6151
R2236 B.n813 B.n28 10.6151
R2237 B.n809 B.n28 10.6151
R2238 B.n809 B.n808 10.6151
R2239 B.n808 B.n807 10.6151
R2240 B.n807 B.n30 10.6151
R2241 B.n803 B.n30 10.6151
R2242 B.n803 B.n802 10.6151
R2243 B.n802 B.n801 10.6151
R2244 B.n801 B.n32 10.6151
R2245 B.n797 B.n32 10.6151
R2246 B.n797 B.n796 10.6151
R2247 B.n796 B.n795 10.6151
R2248 B.n795 B.n34 10.6151
R2249 B.n791 B.n34 10.6151
R2250 B.n791 B.n790 10.6151
R2251 B.n790 B.n789 10.6151
R2252 B.n789 B.n36 10.6151
R2253 B.n785 B.n36 10.6151
R2254 B.n785 B.n784 10.6151
R2255 B.n784 B.n783 10.6151
R2256 B.n783 B.n38 10.6151
R2257 B.n779 B.n38 10.6151
R2258 B.n779 B.n778 10.6151
R2259 B.n778 B.n777 10.6151
R2260 B.n777 B.n40 10.6151
R2261 B.n773 B.n40 10.6151
R2262 B.n773 B.n772 10.6151
R2263 B.n772 B.n771 10.6151
R2264 B.n771 B.n42 10.6151
R2265 B.n767 B.n42 10.6151
R2266 B.n767 B.n766 10.6151
R2267 B.n766 B.n765 10.6151
R2268 B.n765 B.n44 10.6151
R2269 B.n761 B.n44 10.6151
R2270 B.n761 B.n760 10.6151
R2271 B.n760 B.n759 10.6151
R2272 B.n759 B.n46 10.6151
R2273 B.n755 B.n46 10.6151
R2274 B.n755 B.n754 10.6151
R2275 B.n754 B.n753 10.6151
R2276 B.n753 B.n48 10.6151
R2277 B.n749 B.n48 10.6151
R2278 B.n749 B.n748 10.6151
R2279 B.n748 B.n747 10.6151
R2280 B.n747 B.n50 10.6151
R2281 B.n743 B.n50 10.6151
R2282 B.n743 B.n742 10.6151
R2283 B.n742 B.n741 10.6151
R2284 B.n741 B.n52 10.6151
R2285 B.n737 B.n52 10.6151
R2286 B.n737 B.n736 10.6151
R2287 B.n736 B.n735 10.6151
R2288 B.n735 B.n54 10.6151
R2289 B.n731 B.n730 10.6151
R2290 B.n730 B.n729 10.6151
R2291 B.n729 B.n59 10.6151
R2292 B.n725 B.n59 10.6151
R2293 B.n725 B.n724 10.6151
R2294 B.n724 B.n723 10.6151
R2295 B.n723 B.n61 10.6151
R2296 B.n719 B.n61 10.6151
R2297 B.n717 B.n716 10.6151
R2298 B.n716 B.n65 10.6151
R2299 B.n712 B.n65 10.6151
R2300 B.n712 B.n711 10.6151
R2301 B.n711 B.n710 10.6151
R2302 B.n710 B.n67 10.6151
R2303 B.n706 B.n67 10.6151
R2304 B.n706 B.n705 10.6151
R2305 B.n705 B.n704 10.6151
R2306 B.n704 B.n69 10.6151
R2307 B.n700 B.n69 10.6151
R2308 B.n700 B.n699 10.6151
R2309 B.n699 B.n698 10.6151
R2310 B.n698 B.n71 10.6151
R2311 B.n694 B.n71 10.6151
R2312 B.n694 B.n693 10.6151
R2313 B.n693 B.n692 10.6151
R2314 B.n692 B.n73 10.6151
R2315 B.n688 B.n73 10.6151
R2316 B.n688 B.n687 10.6151
R2317 B.n687 B.n686 10.6151
R2318 B.n686 B.n75 10.6151
R2319 B.n682 B.n75 10.6151
R2320 B.n682 B.n681 10.6151
R2321 B.n681 B.n680 10.6151
R2322 B.n680 B.n77 10.6151
R2323 B.n676 B.n77 10.6151
R2324 B.n676 B.n675 10.6151
R2325 B.n675 B.n674 10.6151
R2326 B.n674 B.n79 10.6151
R2327 B.n670 B.n79 10.6151
R2328 B.n670 B.n669 10.6151
R2329 B.n669 B.n668 10.6151
R2330 B.n668 B.n81 10.6151
R2331 B.n664 B.n81 10.6151
R2332 B.n664 B.n663 10.6151
R2333 B.n663 B.n662 10.6151
R2334 B.n662 B.n83 10.6151
R2335 B.n658 B.n83 10.6151
R2336 B.n658 B.n657 10.6151
R2337 B.n657 B.n656 10.6151
R2338 B.n656 B.n85 10.6151
R2339 B.n652 B.n85 10.6151
R2340 B.n652 B.n651 10.6151
R2341 B.n651 B.n650 10.6151
R2342 B.n650 B.n87 10.6151
R2343 B.n646 B.n87 10.6151
R2344 B.n646 B.n645 10.6151
R2345 B.n645 B.n644 10.6151
R2346 B.n644 B.n89 10.6151
R2347 B.n640 B.n89 10.6151
R2348 B.n640 B.n639 10.6151
R2349 B.n639 B.n638 10.6151
R2350 B.n638 B.n91 10.6151
R2351 B.n634 B.n91 10.6151
R2352 B.n634 B.n633 10.6151
R2353 B.n633 B.n632 10.6151
R2354 B.n632 B.n93 10.6151
R2355 B.n628 B.n93 10.6151
R2356 B.n628 B.n627 10.6151
R2357 B.n627 B.n626 10.6151
R2358 B.n626 B.n95 10.6151
R2359 B.n622 B.n95 10.6151
R2360 B.n500 B.n137 10.6151
R2361 B.n501 B.n500 10.6151
R2362 B.n502 B.n501 10.6151
R2363 B.n502 B.n135 10.6151
R2364 B.n506 B.n135 10.6151
R2365 B.n507 B.n506 10.6151
R2366 B.n508 B.n507 10.6151
R2367 B.n508 B.n133 10.6151
R2368 B.n512 B.n133 10.6151
R2369 B.n513 B.n512 10.6151
R2370 B.n514 B.n513 10.6151
R2371 B.n514 B.n131 10.6151
R2372 B.n518 B.n131 10.6151
R2373 B.n519 B.n518 10.6151
R2374 B.n520 B.n519 10.6151
R2375 B.n520 B.n129 10.6151
R2376 B.n524 B.n129 10.6151
R2377 B.n525 B.n524 10.6151
R2378 B.n526 B.n525 10.6151
R2379 B.n526 B.n127 10.6151
R2380 B.n530 B.n127 10.6151
R2381 B.n531 B.n530 10.6151
R2382 B.n532 B.n531 10.6151
R2383 B.n532 B.n125 10.6151
R2384 B.n536 B.n125 10.6151
R2385 B.n537 B.n536 10.6151
R2386 B.n538 B.n537 10.6151
R2387 B.n538 B.n123 10.6151
R2388 B.n542 B.n123 10.6151
R2389 B.n543 B.n542 10.6151
R2390 B.n544 B.n543 10.6151
R2391 B.n544 B.n121 10.6151
R2392 B.n548 B.n121 10.6151
R2393 B.n549 B.n548 10.6151
R2394 B.n550 B.n549 10.6151
R2395 B.n550 B.n119 10.6151
R2396 B.n554 B.n119 10.6151
R2397 B.n555 B.n554 10.6151
R2398 B.n556 B.n555 10.6151
R2399 B.n556 B.n117 10.6151
R2400 B.n560 B.n117 10.6151
R2401 B.n561 B.n560 10.6151
R2402 B.n562 B.n561 10.6151
R2403 B.n562 B.n115 10.6151
R2404 B.n566 B.n115 10.6151
R2405 B.n567 B.n566 10.6151
R2406 B.n568 B.n567 10.6151
R2407 B.n568 B.n113 10.6151
R2408 B.n572 B.n113 10.6151
R2409 B.n573 B.n572 10.6151
R2410 B.n574 B.n573 10.6151
R2411 B.n574 B.n111 10.6151
R2412 B.n578 B.n111 10.6151
R2413 B.n579 B.n578 10.6151
R2414 B.n580 B.n579 10.6151
R2415 B.n580 B.n109 10.6151
R2416 B.n584 B.n109 10.6151
R2417 B.n585 B.n584 10.6151
R2418 B.n586 B.n585 10.6151
R2419 B.n586 B.n107 10.6151
R2420 B.n590 B.n107 10.6151
R2421 B.n591 B.n590 10.6151
R2422 B.n592 B.n591 10.6151
R2423 B.n592 B.n105 10.6151
R2424 B.n596 B.n105 10.6151
R2425 B.n597 B.n596 10.6151
R2426 B.n598 B.n597 10.6151
R2427 B.n598 B.n103 10.6151
R2428 B.n602 B.n103 10.6151
R2429 B.n603 B.n602 10.6151
R2430 B.n604 B.n603 10.6151
R2431 B.n604 B.n101 10.6151
R2432 B.n608 B.n101 10.6151
R2433 B.n609 B.n608 10.6151
R2434 B.n610 B.n609 10.6151
R2435 B.n610 B.n99 10.6151
R2436 B.n614 B.n99 10.6151
R2437 B.n615 B.n614 10.6151
R2438 B.n616 B.n615 10.6151
R2439 B.n616 B.n97 10.6151
R2440 B.n620 B.n97 10.6151
R2441 B.n621 B.n620 10.6151
R2442 B.n288 B.n207 10.6151
R2443 B.n292 B.n207 10.6151
R2444 B.n293 B.n292 10.6151
R2445 B.n294 B.n293 10.6151
R2446 B.n294 B.n205 10.6151
R2447 B.n298 B.n205 10.6151
R2448 B.n299 B.n298 10.6151
R2449 B.n300 B.n299 10.6151
R2450 B.n300 B.n203 10.6151
R2451 B.n304 B.n203 10.6151
R2452 B.n305 B.n304 10.6151
R2453 B.n306 B.n305 10.6151
R2454 B.n306 B.n201 10.6151
R2455 B.n310 B.n201 10.6151
R2456 B.n311 B.n310 10.6151
R2457 B.n312 B.n311 10.6151
R2458 B.n312 B.n199 10.6151
R2459 B.n316 B.n199 10.6151
R2460 B.n317 B.n316 10.6151
R2461 B.n318 B.n317 10.6151
R2462 B.n318 B.n197 10.6151
R2463 B.n322 B.n197 10.6151
R2464 B.n323 B.n322 10.6151
R2465 B.n324 B.n323 10.6151
R2466 B.n324 B.n195 10.6151
R2467 B.n328 B.n195 10.6151
R2468 B.n329 B.n328 10.6151
R2469 B.n330 B.n329 10.6151
R2470 B.n330 B.n193 10.6151
R2471 B.n334 B.n193 10.6151
R2472 B.n335 B.n334 10.6151
R2473 B.n336 B.n335 10.6151
R2474 B.n336 B.n191 10.6151
R2475 B.n340 B.n191 10.6151
R2476 B.n341 B.n340 10.6151
R2477 B.n342 B.n341 10.6151
R2478 B.n342 B.n189 10.6151
R2479 B.n346 B.n189 10.6151
R2480 B.n347 B.n346 10.6151
R2481 B.n348 B.n347 10.6151
R2482 B.n348 B.n187 10.6151
R2483 B.n352 B.n187 10.6151
R2484 B.n353 B.n352 10.6151
R2485 B.n354 B.n353 10.6151
R2486 B.n354 B.n185 10.6151
R2487 B.n358 B.n185 10.6151
R2488 B.n359 B.n358 10.6151
R2489 B.n360 B.n359 10.6151
R2490 B.n360 B.n183 10.6151
R2491 B.n364 B.n183 10.6151
R2492 B.n365 B.n364 10.6151
R2493 B.n366 B.n365 10.6151
R2494 B.n366 B.n181 10.6151
R2495 B.n370 B.n181 10.6151
R2496 B.n371 B.n370 10.6151
R2497 B.n372 B.n371 10.6151
R2498 B.n372 B.n179 10.6151
R2499 B.n376 B.n179 10.6151
R2500 B.n377 B.n376 10.6151
R2501 B.n378 B.n377 10.6151
R2502 B.n378 B.n177 10.6151
R2503 B.n382 B.n177 10.6151
R2504 B.n383 B.n382 10.6151
R2505 B.n385 B.n173 10.6151
R2506 B.n389 B.n173 10.6151
R2507 B.n390 B.n389 10.6151
R2508 B.n391 B.n390 10.6151
R2509 B.n391 B.n171 10.6151
R2510 B.n395 B.n171 10.6151
R2511 B.n396 B.n395 10.6151
R2512 B.n400 B.n396 10.6151
R2513 B.n404 B.n169 10.6151
R2514 B.n405 B.n404 10.6151
R2515 B.n406 B.n405 10.6151
R2516 B.n406 B.n167 10.6151
R2517 B.n410 B.n167 10.6151
R2518 B.n411 B.n410 10.6151
R2519 B.n412 B.n411 10.6151
R2520 B.n412 B.n165 10.6151
R2521 B.n416 B.n165 10.6151
R2522 B.n417 B.n416 10.6151
R2523 B.n418 B.n417 10.6151
R2524 B.n418 B.n163 10.6151
R2525 B.n422 B.n163 10.6151
R2526 B.n423 B.n422 10.6151
R2527 B.n424 B.n423 10.6151
R2528 B.n424 B.n161 10.6151
R2529 B.n428 B.n161 10.6151
R2530 B.n429 B.n428 10.6151
R2531 B.n430 B.n429 10.6151
R2532 B.n430 B.n159 10.6151
R2533 B.n434 B.n159 10.6151
R2534 B.n435 B.n434 10.6151
R2535 B.n436 B.n435 10.6151
R2536 B.n436 B.n157 10.6151
R2537 B.n440 B.n157 10.6151
R2538 B.n441 B.n440 10.6151
R2539 B.n442 B.n441 10.6151
R2540 B.n442 B.n155 10.6151
R2541 B.n446 B.n155 10.6151
R2542 B.n447 B.n446 10.6151
R2543 B.n448 B.n447 10.6151
R2544 B.n448 B.n153 10.6151
R2545 B.n452 B.n153 10.6151
R2546 B.n453 B.n452 10.6151
R2547 B.n454 B.n453 10.6151
R2548 B.n454 B.n151 10.6151
R2549 B.n458 B.n151 10.6151
R2550 B.n459 B.n458 10.6151
R2551 B.n460 B.n459 10.6151
R2552 B.n460 B.n149 10.6151
R2553 B.n464 B.n149 10.6151
R2554 B.n465 B.n464 10.6151
R2555 B.n466 B.n465 10.6151
R2556 B.n466 B.n147 10.6151
R2557 B.n470 B.n147 10.6151
R2558 B.n471 B.n470 10.6151
R2559 B.n472 B.n471 10.6151
R2560 B.n472 B.n145 10.6151
R2561 B.n476 B.n145 10.6151
R2562 B.n477 B.n476 10.6151
R2563 B.n478 B.n477 10.6151
R2564 B.n478 B.n143 10.6151
R2565 B.n482 B.n143 10.6151
R2566 B.n483 B.n482 10.6151
R2567 B.n484 B.n483 10.6151
R2568 B.n484 B.n141 10.6151
R2569 B.n488 B.n141 10.6151
R2570 B.n489 B.n488 10.6151
R2571 B.n490 B.n489 10.6151
R2572 B.n490 B.n139 10.6151
R2573 B.n494 B.n139 10.6151
R2574 B.n495 B.n494 10.6151
R2575 B.n496 B.n495 10.6151
R2576 B.n287 B.n286 10.6151
R2577 B.n286 B.n209 10.6151
R2578 B.n282 B.n209 10.6151
R2579 B.n282 B.n281 10.6151
R2580 B.n281 B.n280 10.6151
R2581 B.n280 B.n211 10.6151
R2582 B.n276 B.n211 10.6151
R2583 B.n276 B.n275 10.6151
R2584 B.n275 B.n274 10.6151
R2585 B.n274 B.n213 10.6151
R2586 B.n270 B.n213 10.6151
R2587 B.n270 B.n269 10.6151
R2588 B.n269 B.n268 10.6151
R2589 B.n268 B.n215 10.6151
R2590 B.n264 B.n215 10.6151
R2591 B.n264 B.n263 10.6151
R2592 B.n263 B.n262 10.6151
R2593 B.n262 B.n217 10.6151
R2594 B.n258 B.n217 10.6151
R2595 B.n258 B.n257 10.6151
R2596 B.n257 B.n256 10.6151
R2597 B.n256 B.n219 10.6151
R2598 B.n252 B.n219 10.6151
R2599 B.n252 B.n251 10.6151
R2600 B.n251 B.n250 10.6151
R2601 B.n250 B.n221 10.6151
R2602 B.n246 B.n221 10.6151
R2603 B.n246 B.n245 10.6151
R2604 B.n245 B.n244 10.6151
R2605 B.n244 B.n223 10.6151
R2606 B.n240 B.n223 10.6151
R2607 B.n240 B.n239 10.6151
R2608 B.n239 B.n238 10.6151
R2609 B.n238 B.n225 10.6151
R2610 B.n234 B.n225 10.6151
R2611 B.n234 B.n233 10.6151
R2612 B.n233 B.n232 10.6151
R2613 B.n232 B.n227 10.6151
R2614 B.n228 B.n227 10.6151
R2615 B.n228 B.n0 10.6151
R2616 B.n887 B.n1 10.6151
R2617 B.n887 B.n886 10.6151
R2618 B.n886 B.n885 10.6151
R2619 B.n885 B.n4 10.6151
R2620 B.n881 B.n4 10.6151
R2621 B.n881 B.n880 10.6151
R2622 B.n880 B.n879 10.6151
R2623 B.n879 B.n6 10.6151
R2624 B.n875 B.n6 10.6151
R2625 B.n875 B.n874 10.6151
R2626 B.n874 B.n873 10.6151
R2627 B.n873 B.n8 10.6151
R2628 B.n869 B.n8 10.6151
R2629 B.n869 B.n868 10.6151
R2630 B.n868 B.n867 10.6151
R2631 B.n867 B.n10 10.6151
R2632 B.n863 B.n10 10.6151
R2633 B.n863 B.n862 10.6151
R2634 B.n862 B.n861 10.6151
R2635 B.n861 B.n12 10.6151
R2636 B.n857 B.n12 10.6151
R2637 B.n857 B.n856 10.6151
R2638 B.n856 B.n855 10.6151
R2639 B.n855 B.n14 10.6151
R2640 B.n851 B.n14 10.6151
R2641 B.n851 B.n850 10.6151
R2642 B.n850 B.n849 10.6151
R2643 B.n849 B.n16 10.6151
R2644 B.n845 B.n16 10.6151
R2645 B.n845 B.n844 10.6151
R2646 B.n844 B.n843 10.6151
R2647 B.n843 B.n18 10.6151
R2648 B.n839 B.n18 10.6151
R2649 B.n839 B.n838 10.6151
R2650 B.n838 B.n837 10.6151
R2651 B.n837 B.n20 10.6151
R2652 B.n833 B.n20 10.6151
R2653 B.n833 B.n832 10.6151
R2654 B.n832 B.n831 10.6151
R2655 B.n831 B.n22 10.6151
R2656 B.n731 B.n58 6.5566
R2657 B.n719 B.n718 6.5566
R2658 B.n385 B.n384 6.5566
R2659 B.n400 B.n399 6.5566
R2660 B.n58 B.n54 4.05904
R2661 B.n718 B.n717 4.05904
R2662 B.n384 B.n383 4.05904
R2663 B.n399 B.n169 4.05904
R2664 B.n891 B.n0 2.81026
R2665 B.n891 B.n1 2.81026
R2666 VN.n1 VN.t1 171.585
R2667 VN.n0 VN.t2 171.585
R2668 VN.n0 VN.t0 170.387
R2669 VN.n1 VN.t3 170.387
R2670 VN VN.n1 56.859
R2671 VN VN.n0 2.28707
R2672 VDD2.n2 VDD2.n0 120.722
R2673 VDD2.n2 VDD2.n1 70.5582
R2674 VDD2.n1 VDD2.t0 1.67085
R2675 VDD2.n1 VDD2.t2 1.67085
R2676 VDD2.n0 VDD2.t1 1.67085
R2677 VDD2.n0 VDD2.t3 1.67085
R2678 VDD2 VDD2.n2 0.0586897
C0 VDD1 B 1.60598f
C1 VN VP 8.15643f
C2 VDD2 B 1.67155f
C3 VDD1 VN 0.150214f
C4 VDD2 VN 7.83932f
C5 w_n3214_n4860# VP 6.15129f
C6 VTAIL VP 7.53899f
C7 VN B 1.35453f
C8 VDD1 w_n3214_n4860# 1.80799f
C9 VDD1 VTAIL 7.21895f
C10 VDD2 w_n3214_n4860# 1.88199f
C11 VDD2 VTAIL 7.27859f
C12 w_n3214_n4860# B 12.332999f
C13 VTAIL B 7.83024f
C14 VN w_n3214_n4860# 5.73607f
C15 VN VTAIL 7.52488f
C16 VDD1 VP 8.13449f
C17 VTAIL w_n3214_n4860# 5.63935f
C18 VDD2 VP 0.446329f
C19 B VP 2.04734f
C20 VDD1 VDD2 1.21812f
C21 VDD2 VSUBS 1.259394f
C22 VDD1 VSUBS 7.08474f
C23 VTAIL VSUBS 1.654527f
C24 VN VSUBS 6.14702f
C25 VP VSUBS 2.984601f
C26 B VSUBS 5.603952f
C27 w_n3214_n4860# VSUBS 0.190796p
C28 VDD2.t1 VSUBS 0.408124f
C29 VDD2.t3 VSUBS 0.408124f
C30 VDD2.n0 VSUBS 4.48253f
C31 VDD2.t0 VSUBS 0.408124f
C32 VDD2.t2 VSUBS 0.408124f
C33 VDD2.n1 VSUBS 3.44257f
C34 VDD2.n2 VSUBS 5.26097f
C35 VN.t0 VSUBS 4.85174f
C36 VN.t2 VSUBS 4.86355f
C37 VN.n0 VSUBS 3.01883f
C38 VN.t1 VSUBS 4.86355f
C39 VN.t3 VSUBS 4.85174f
C40 VN.n1 VSUBS 4.80184f
C41 B.n0 VSUBS 0.003808f
C42 B.n1 VSUBS 0.003808f
C43 B.n2 VSUBS 0.006021f
C44 B.n3 VSUBS 0.006021f
C45 B.n4 VSUBS 0.006021f
C46 B.n5 VSUBS 0.006021f
C47 B.n6 VSUBS 0.006021f
C48 B.n7 VSUBS 0.006021f
C49 B.n8 VSUBS 0.006021f
C50 B.n9 VSUBS 0.006021f
C51 B.n10 VSUBS 0.006021f
C52 B.n11 VSUBS 0.006021f
C53 B.n12 VSUBS 0.006021f
C54 B.n13 VSUBS 0.006021f
C55 B.n14 VSUBS 0.006021f
C56 B.n15 VSUBS 0.006021f
C57 B.n16 VSUBS 0.006021f
C58 B.n17 VSUBS 0.006021f
C59 B.n18 VSUBS 0.006021f
C60 B.n19 VSUBS 0.006021f
C61 B.n20 VSUBS 0.006021f
C62 B.n21 VSUBS 0.006021f
C63 B.n22 VSUBS 0.013397f
C64 B.n23 VSUBS 0.006021f
C65 B.n24 VSUBS 0.006021f
C66 B.n25 VSUBS 0.006021f
C67 B.n26 VSUBS 0.006021f
C68 B.n27 VSUBS 0.006021f
C69 B.n28 VSUBS 0.006021f
C70 B.n29 VSUBS 0.006021f
C71 B.n30 VSUBS 0.006021f
C72 B.n31 VSUBS 0.006021f
C73 B.n32 VSUBS 0.006021f
C74 B.n33 VSUBS 0.006021f
C75 B.n34 VSUBS 0.006021f
C76 B.n35 VSUBS 0.006021f
C77 B.n36 VSUBS 0.006021f
C78 B.n37 VSUBS 0.006021f
C79 B.n38 VSUBS 0.006021f
C80 B.n39 VSUBS 0.006021f
C81 B.n40 VSUBS 0.006021f
C82 B.n41 VSUBS 0.006021f
C83 B.n42 VSUBS 0.006021f
C84 B.n43 VSUBS 0.006021f
C85 B.n44 VSUBS 0.006021f
C86 B.n45 VSUBS 0.006021f
C87 B.n46 VSUBS 0.006021f
C88 B.n47 VSUBS 0.006021f
C89 B.n48 VSUBS 0.006021f
C90 B.n49 VSUBS 0.006021f
C91 B.n50 VSUBS 0.006021f
C92 B.n51 VSUBS 0.006021f
C93 B.n52 VSUBS 0.006021f
C94 B.n53 VSUBS 0.006021f
C95 B.n54 VSUBS 0.004162f
C96 B.n55 VSUBS 0.006021f
C97 B.t11 VSUBS 0.332439f
C98 B.t10 VSUBS 0.368806f
C99 B.t9 VSUBS 2.56894f
C100 B.n56 VSUBS 0.584369f
C101 B.n57 VSUBS 0.300596f
C102 B.n58 VSUBS 0.013951f
C103 B.n59 VSUBS 0.006021f
C104 B.n60 VSUBS 0.006021f
C105 B.n61 VSUBS 0.006021f
C106 B.n62 VSUBS 0.006021f
C107 B.t8 VSUBS 0.332442f
C108 B.t7 VSUBS 0.368809f
C109 B.t6 VSUBS 2.56894f
C110 B.n63 VSUBS 0.584366f
C111 B.n64 VSUBS 0.300593f
C112 B.n65 VSUBS 0.006021f
C113 B.n66 VSUBS 0.006021f
C114 B.n67 VSUBS 0.006021f
C115 B.n68 VSUBS 0.006021f
C116 B.n69 VSUBS 0.006021f
C117 B.n70 VSUBS 0.006021f
C118 B.n71 VSUBS 0.006021f
C119 B.n72 VSUBS 0.006021f
C120 B.n73 VSUBS 0.006021f
C121 B.n74 VSUBS 0.006021f
C122 B.n75 VSUBS 0.006021f
C123 B.n76 VSUBS 0.006021f
C124 B.n77 VSUBS 0.006021f
C125 B.n78 VSUBS 0.006021f
C126 B.n79 VSUBS 0.006021f
C127 B.n80 VSUBS 0.006021f
C128 B.n81 VSUBS 0.006021f
C129 B.n82 VSUBS 0.006021f
C130 B.n83 VSUBS 0.006021f
C131 B.n84 VSUBS 0.006021f
C132 B.n85 VSUBS 0.006021f
C133 B.n86 VSUBS 0.006021f
C134 B.n87 VSUBS 0.006021f
C135 B.n88 VSUBS 0.006021f
C136 B.n89 VSUBS 0.006021f
C137 B.n90 VSUBS 0.006021f
C138 B.n91 VSUBS 0.006021f
C139 B.n92 VSUBS 0.006021f
C140 B.n93 VSUBS 0.006021f
C141 B.n94 VSUBS 0.006021f
C142 B.n95 VSUBS 0.006021f
C143 B.n96 VSUBS 0.013397f
C144 B.n97 VSUBS 0.006021f
C145 B.n98 VSUBS 0.006021f
C146 B.n99 VSUBS 0.006021f
C147 B.n100 VSUBS 0.006021f
C148 B.n101 VSUBS 0.006021f
C149 B.n102 VSUBS 0.006021f
C150 B.n103 VSUBS 0.006021f
C151 B.n104 VSUBS 0.006021f
C152 B.n105 VSUBS 0.006021f
C153 B.n106 VSUBS 0.006021f
C154 B.n107 VSUBS 0.006021f
C155 B.n108 VSUBS 0.006021f
C156 B.n109 VSUBS 0.006021f
C157 B.n110 VSUBS 0.006021f
C158 B.n111 VSUBS 0.006021f
C159 B.n112 VSUBS 0.006021f
C160 B.n113 VSUBS 0.006021f
C161 B.n114 VSUBS 0.006021f
C162 B.n115 VSUBS 0.006021f
C163 B.n116 VSUBS 0.006021f
C164 B.n117 VSUBS 0.006021f
C165 B.n118 VSUBS 0.006021f
C166 B.n119 VSUBS 0.006021f
C167 B.n120 VSUBS 0.006021f
C168 B.n121 VSUBS 0.006021f
C169 B.n122 VSUBS 0.006021f
C170 B.n123 VSUBS 0.006021f
C171 B.n124 VSUBS 0.006021f
C172 B.n125 VSUBS 0.006021f
C173 B.n126 VSUBS 0.006021f
C174 B.n127 VSUBS 0.006021f
C175 B.n128 VSUBS 0.006021f
C176 B.n129 VSUBS 0.006021f
C177 B.n130 VSUBS 0.006021f
C178 B.n131 VSUBS 0.006021f
C179 B.n132 VSUBS 0.006021f
C180 B.n133 VSUBS 0.006021f
C181 B.n134 VSUBS 0.006021f
C182 B.n135 VSUBS 0.006021f
C183 B.n136 VSUBS 0.006021f
C184 B.n137 VSUBS 0.013397f
C185 B.n138 VSUBS 0.006021f
C186 B.n139 VSUBS 0.006021f
C187 B.n140 VSUBS 0.006021f
C188 B.n141 VSUBS 0.006021f
C189 B.n142 VSUBS 0.006021f
C190 B.n143 VSUBS 0.006021f
C191 B.n144 VSUBS 0.006021f
C192 B.n145 VSUBS 0.006021f
C193 B.n146 VSUBS 0.006021f
C194 B.n147 VSUBS 0.006021f
C195 B.n148 VSUBS 0.006021f
C196 B.n149 VSUBS 0.006021f
C197 B.n150 VSUBS 0.006021f
C198 B.n151 VSUBS 0.006021f
C199 B.n152 VSUBS 0.006021f
C200 B.n153 VSUBS 0.006021f
C201 B.n154 VSUBS 0.006021f
C202 B.n155 VSUBS 0.006021f
C203 B.n156 VSUBS 0.006021f
C204 B.n157 VSUBS 0.006021f
C205 B.n158 VSUBS 0.006021f
C206 B.n159 VSUBS 0.006021f
C207 B.n160 VSUBS 0.006021f
C208 B.n161 VSUBS 0.006021f
C209 B.n162 VSUBS 0.006021f
C210 B.n163 VSUBS 0.006021f
C211 B.n164 VSUBS 0.006021f
C212 B.n165 VSUBS 0.006021f
C213 B.n166 VSUBS 0.006021f
C214 B.n167 VSUBS 0.006021f
C215 B.n168 VSUBS 0.006021f
C216 B.n169 VSUBS 0.004162f
C217 B.n170 VSUBS 0.006021f
C218 B.n171 VSUBS 0.006021f
C219 B.n172 VSUBS 0.006021f
C220 B.n173 VSUBS 0.006021f
C221 B.n174 VSUBS 0.006021f
C222 B.t4 VSUBS 0.332439f
C223 B.t5 VSUBS 0.368806f
C224 B.t3 VSUBS 2.56894f
C225 B.n175 VSUBS 0.584369f
C226 B.n176 VSUBS 0.300596f
C227 B.n177 VSUBS 0.006021f
C228 B.n178 VSUBS 0.006021f
C229 B.n179 VSUBS 0.006021f
C230 B.n180 VSUBS 0.006021f
C231 B.n181 VSUBS 0.006021f
C232 B.n182 VSUBS 0.006021f
C233 B.n183 VSUBS 0.006021f
C234 B.n184 VSUBS 0.006021f
C235 B.n185 VSUBS 0.006021f
C236 B.n186 VSUBS 0.006021f
C237 B.n187 VSUBS 0.006021f
C238 B.n188 VSUBS 0.006021f
C239 B.n189 VSUBS 0.006021f
C240 B.n190 VSUBS 0.006021f
C241 B.n191 VSUBS 0.006021f
C242 B.n192 VSUBS 0.006021f
C243 B.n193 VSUBS 0.006021f
C244 B.n194 VSUBS 0.006021f
C245 B.n195 VSUBS 0.006021f
C246 B.n196 VSUBS 0.006021f
C247 B.n197 VSUBS 0.006021f
C248 B.n198 VSUBS 0.006021f
C249 B.n199 VSUBS 0.006021f
C250 B.n200 VSUBS 0.006021f
C251 B.n201 VSUBS 0.006021f
C252 B.n202 VSUBS 0.006021f
C253 B.n203 VSUBS 0.006021f
C254 B.n204 VSUBS 0.006021f
C255 B.n205 VSUBS 0.006021f
C256 B.n206 VSUBS 0.006021f
C257 B.n207 VSUBS 0.006021f
C258 B.n208 VSUBS 0.013397f
C259 B.n209 VSUBS 0.006021f
C260 B.n210 VSUBS 0.006021f
C261 B.n211 VSUBS 0.006021f
C262 B.n212 VSUBS 0.006021f
C263 B.n213 VSUBS 0.006021f
C264 B.n214 VSUBS 0.006021f
C265 B.n215 VSUBS 0.006021f
C266 B.n216 VSUBS 0.006021f
C267 B.n217 VSUBS 0.006021f
C268 B.n218 VSUBS 0.006021f
C269 B.n219 VSUBS 0.006021f
C270 B.n220 VSUBS 0.006021f
C271 B.n221 VSUBS 0.006021f
C272 B.n222 VSUBS 0.006021f
C273 B.n223 VSUBS 0.006021f
C274 B.n224 VSUBS 0.006021f
C275 B.n225 VSUBS 0.006021f
C276 B.n226 VSUBS 0.006021f
C277 B.n227 VSUBS 0.006021f
C278 B.n228 VSUBS 0.006021f
C279 B.n229 VSUBS 0.006021f
C280 B.n230 VSUBS 0.006021f
C281 B.n231 VSUBS 0.006021f
C282 B.n232 VSUBS 0.006021f
C283 B.n233 VSUBS 0.006021f
C284 B.n234 VSUBS 0.006021f
C285 B.n235 VSUBS 0.006021f
C286 B.n236 VSUBS 0.006021f
C287 B.n237 VSUBS 0.006021f
C288 B.n238 VSUBS 0.006021f
C289 B.n239 VSUBS 0.006021f
C290 B.n240 VSUBS 0.006021f
C291 B.n241 VSUBS 0.006021f
C292 B.n242 VSUBS 0.006021f
C293 B.n243 VSUBS 0.006021f
C294 B.n244 VSUBS 0.006021f
C295 B.n245 VSUBS 0.006021f
C296 B.n246 VSUBS 0.006021f
C297 B.n247 VSUBS 0.006021f
C298 B.n248 VSUBS 0.006021f
C299 B.n249 VSUBS 0.006021f
C300 B.n250 VSUBS 0.006021f
C301 B.n251 VSUBS 0.006021f
C302 B.n252 VSUBS 0.006021f
C303 B.n253 VSUBS 0.006021f
C304 B.n254 VSUBS 0.006021f
C305 B.n255 VSUBS 0.006021f
C306 B.n256 VSUBS 0.006021f
C307 B.n257 VSUBS 0.006021f
C308 B.n258 VSUBS 0.006021f
C309 B.n259 VSUBS 0.006021f
C310 B.n260 VSUBS 0.006021f
C311 B.n261 VSUBS 0.006021f
C312 B.n262 VSUBS 0.006021f
C313 B.n263 VSUBS 0.006021f
C314 B.n264 VSUBS 0.006021f
C315 B.n265 VSUBS 0.006021f
C316 B.n266 VSUBS 0.006021f
C317 B.n267 VSUBS 0.006021f
C318 B.n268 VSUBS 0.006021f
C319 B.n269 VSUBS 0.006021f
C320 B.n270 VSUBS 0.006021f
C321 B.n271 VSUBS 0.006021f
C322 B.n272 VSUBS 0.006021f
C323 B.n273 VSUBS 0.006021f
C324 B.n274 VSUBS 0.006021f
C325 B.n275 VSUBS 0.006021f
C326 B.n276 VSUBS 0.006021f
C327 B.n277 VSUBS 0.006021f
C328 B.n278 VSUBS 0.006021f
C329 B.n279 VSUBS 0.006021f
C330 B.n280 VSUBS 0.006021f
C331 B.n281 VSUBS 0.006021f
C332 B.n282 VSUBS 0.006021f
C333 B.n283 VSUBS 0.006021f
C334 B.n284 VSUBS 0.006021f
C335 B.n285 VSUBS 0.006021f
C336 B.n286 VSUBS 0.006021f
C337 B.n287 VSUBS 0.013397f
C338 B.n288 VSUBS 0.014407f
C339 B.n289 VSUBS 0.014407f
C340 B.n290 VSUBS 0.006021f
C341 B.n291 VSUBS 0.006021f
C342 B.n292 VSUBS 0.006021f
C343 B.n293 VSUBS 0.006021f
C344 B.n294 VSUBS 0.006021f
C345 B.n295 VSUBS 0.006021f
C346 B.n296 VSUBS 0.006021f
C347 B.n297 VSUBS 0.006021f
C348 B.n298 VSUBS 0.006021f
C349 B.n299 VSUBS 0.006021f
C350 B.n300 VSUBS 0.006021f
C351 B.n301 VSUBS 0.006021f
C352 B.n302 VSUBS 0.006021f
C353 B.n303 VSUBS 0.006021f
C354 B.n304 VSUBS 0.006021f
C355 B.n305 VSUBS 0.006021f
C356 B.n306 VSUBS 0.006021f
C357 B.n307 VSUBS 0.006021f
C358 B.n308 VSUBS 0.006021f
C359 B.n309 VSUBS 0.006021f
C360 B.n310 VSUBS 0.006021f
C361 B.n311 VSUBS 0.006021f
C362 B.n312 VSUBS 0.006021f
C363 B.n313 VSUBS 0.006021f
C364 B.n314 VSUBS 0.006021f
C365 B.n315 VSUBS 0.006021f
C366 B.n316 VSUBS 0.006021f
C367 B.n317 VSUBS 0.006021f
C368 B.n318 VSUBS 0.006021f
C369 B.n319 VSUBS 0.006021f
C370 B.n320 VSUBS 0.006021f
C371 B.n321 VSUBS 0.006021f
C372 B.n322 VSUBS 0.006021f
C373 B.n323 VSUBS 0.006021f
C374 B.n324 VSUBS 0.006021f
C375 B.n325 VSUBS 0.006021f
C376 B.n326 VSUBS 0.006021f
C377 B.n327 VSUBS 0.006021f
C378 B.n328 VSUBS 0.006021f
C379 B.n329 VSUBS 0.006021f
C380 B.n330 VSUBS 0.006021f
C381 B.n331 VSUBS 0.006021f
C382 B.n332 VSUBS 0.006021f
C383 B.n333 VSUBS 0.006021f
C384 B.n334 VSUBS 0.006021f
C385 B.n335 VSUBS 0.006021f
C386 B.n336 VSUBS 0.006021f
C387 B.n337 VSUBS 0.006021f
C388 B.n338 VSUBS 0.006021f
C389 B.n339 VSUBS 0.006021f
C390 B.n340 VSUBS 0.006021f
C391 B.n341 VSUBS 0.006021f
C392 B.n342 VSUBS 0.006021f
C393 B.n343 VSUBS 0.006021f
C394 B.n344 VSUBS 0.006021f
C395 B.n345 VSUBS 0.006021f
C396 B.n346 VSUBS 0.006021f
C397 B.n347 VSUBS 0.006021f
C398 B.n348 VSUBS 0.006021f
C399 B.n349 VSUBS 0.006021f
C400 B.n350 VSUBS 0.006021f
C401 B.n351 VSUBS 0.006021f
C402 B.n352 VSUBS 0.006021f
C403 B.n353 VSUBS 0.006021f
C404 B.n354 VSUBS 0.006021f
C405 B.n355 VSUBS 0.006021f
C406 B.n356 VSUBS 0.006021f
C407 B.n357 VSUBS 0.006021f
C408 B.n358 VSUBS 0.006021f
C409 B.n359 VSUBS 0.006021f
C410 B.n360 VSUBS 0.006021f
C411 B.n361 VSUBS 0.006021f
C412 B.n362 VSUBS 0.006021f
C413 B.n363 VSUBS 0.006021f
C414 B.n364 VSUBS 0.006021f
C415 B.n365 VSUBS 0.006021f
C416 B.n366 VSUBS 0.006021f
C417 B.n367 VSUBS 0.006021f
C418 B.n368 VSUBS 0.006021f
C419 B.n369 VSUBS 0.006021f
C420 B.n370 VSUBS 0.006021f
C421 B.n371 VSUBS 0.006021f
C422 B.n372 VSUBS 0.006021f
C423 B.n373 VSUBS 0.006021f
C424 B.n374 VSUBS 0.006021f
C425 B.n375 VSUBS 0.006021f
C426 B.n376 VSUBS 0.006021f
C427 B.n377 VSUBS 0.006021f
C428 B.n378 VSUBS 0.006021f
C429 B.n379 VSUBS 0.006021f
C430 B.n380 VSUBS 0.006021f
C431 B.n381 VSUBS 0.006021f
C432 B.n382 VSUBS 0.006021f
C433 B.n383 VSUBS 0.004162f
C434 B.n384 VSUBS 0.013951f
C435 B.n385 VSUBS 0.00487f
C436 B.n386 VSUBS 0.006021f
C437 B.n387 VSUBS 0.006021f
C438 B.n388 VSUBS 0.006021f
C439 B.n389 VSUBS 0.006021f
C440 B.n390 VSUBS 0.006021f
C441 B.n391 VSUBS 0.006021f
C442 B.n392 VSUBS 0.006021f
C443 B.n393 VSUBS 0.006021f
C444 B.n394 VSUBS 0.006021f
C445 B.n395 VSUBS 0.006021f
C446 B.n396 VSUBS 0.006021f
C447 B.t1 VSUBS 0.332442f
C448 B.t2 VSUBS 0.368809f
C449 B.t0 VSUBS 2.56894f
C450 B.n397 VSUBS 0.584366f
C451 B.n398 VSUBS 0.300593f
C452 B.n399 VSUBS 0.013951f
C453 B.n400 VSUBS 0.00487f
C454 B.n401 VSUBS 0.006021f
C455 B.n402 VSUBS 0.006021f
C456 B.n403 VSUBS 0.006021f
C457 B.n404 VSUBS 0.006021f
C458 B.n405 VSUBS 0.006021f
C459 B.n406 VSUBS 0.006021f
C460 B.n407 VSUBS 0.006021f
C461 B.n408 VSUBS 0.006021f
C462 B.n409 VSUBS 0.006021f
C463 B.n410 VSUBS 0.006021f
C464 B.n411 VSUBS 0.006021f
C465 B.n412 VSUBS 0.006021f
C466 B.n413 VSUBS 0.006021f
C467 B.n414 VSUBS 0.006021f
C468 B.n415 VSUBS 0.006021f
C469 B.n416 VSUBS 0.006021f
C470 B.n417 VSUBS 0.006021f
C471 B.n418 VSUBS 0.006021f
C472 B.n419 VSUBS 0.006021f
C473 B.n420 VSUBS 0.006021f
C474 B.n421 VSUBS 0.006021f
C475 B.n422 VSUBS 0.006021f
C476 B.n423 VSUBS 0.006021f
C477 B.n424 VSUBS 0.006021f
C478 B.n425 VSUBS 0.006021f
C479 B.n426 VSUBS 0.006021f
C480 B.n427 VSUBS 0.006021f
C481 B.n428 VSUBS 0.006021f
C482 B.n429 VSUBS 0.006021f
C483 B.n430 VSUBS 0.006021f
C484 B.n431 VSUBS 0.006021f
C485 B.n432 VSUBS 0.006021f
C486 B.n433 VSUBS 0.006021f
C487 B.n434 VSUBS 0.006021f
C488 B.n435 VSUBS 0.006021f
C489 B.n436 VSUBS 0.006021f
C490 B.n437 VSUBS 0.006021f
C491 B.n438 VSUBS 0.006021f
C492 B.n439 VSUBS 0.006021f
C493 B.n440 VSUBS 0.006021f
C494 B.n441 VSUBS 0.006021f
C495 B.n442 VSUBS 0.006021f
C496 B.n443 VSUBS 0.006021f
C497 B.n444 VSUBS 0.006021f
C498 B.n445 VSUBS 0.006021f
C499 B.n446 VSUBS 0.006021f
C500 B.n447 VSUBS 0.006021f
C501 B.n448 VSUBS 0.006021f
C502 B.n449 VSUBS 0.006021f
C503 B.n450 VSUBS 0.006021f
C504 B.n451 VSUBS 0.006021f
C505 B.n452 VSUBS 0.006021f
C506 B.n453 VSUBS 0.006021f
C507 B.n454 VSUBS 0.006021f
C508 B.n455 VSUBS 0.006021f
C509 B.n456 VSUBS 0.006021f
C510 B.n457 VSUBS 0.006021f
C511 B.n458 VSUBS 0.006021f
C512 B.n459 VSUBS 0.006021f
C513 B.n460 VSUBS 0.006021f
C514 B.n461 VSUBS 0.006021f
C515 B.n462 VSUBS 0.006021f
C516 B.n463 VSUBS 0.006021f
C517 B.n464 VSUBS 0.006021f
C518 B.n465 VSUBS 0.006021f
C519 B.n466 VSUBS 0.006021f
C520 B.n467 VSUBS 0.006021f
C521 B.n468 VSUBS 0.006021f
C522 B.n469 VSUBS 0.006021f
C523 B.n470 VSUBS 0.006021f
C524 B.n471 VSUBS 0.006021f
C525 B.n472 VSUBS 0.006021f
C526 B.n473 VSUBS 0.006021f
C527 B.n474 VSUBS 0.006021f
C528 B.n475 VSUBS 0.006021f
C529 B.n476 VSUBS 0.006021f
C530 B.n477 VSUBS 0.006021f
C531 B.n478 VSUBS 0.006021f
C532 B.n479 VSUBS 0.006021f
C533 B.n480 VSUBS 0.006021f
C534 B.n481 VSUBS 0.006021f
C535 B.n482 VSUBS 0.006021f
C536 B.n483 VSUBS 0.006021f
C537 B.n484 VSUBS 0.006021f
C538 B.n485 VSUBS 0.006021f
C539 B.n486 VSUBS 0.006021f
C540 B.n487 VSUBS 0.006021f
C541 B.n488 VSUBS 0.006021f
C542 B.n489 VSUBS 0.006021f
C543 B.n490 VSUBS 0.006021f
C544 B.n491 VSUBS 0.006021f
C545 B.n492 VSUBS 0.006021f
C546 B.n493 VSUBS 0.006021f
C547 B.n494 VSUBS 0.006021f
C548 B.n495 VSUBS 0.006021f
C549 B.n496 VSUBS 0.014407f
C550 B.n497 VSUBS 0.014407f
C551 B.n498 VSUBS 0.013397f
C552 B.n499 VSUBS 0.006021f
C553 B.n500 VSUBS 0.006021f
C554 B.n501 VSUBS 0.006021f
C555 B.n502 VSUBS 0.006021f
C556 B.n503 VSUBS 0.006021f
C557 B.n504 VSUBS 0.006021f
C558 B.n505 VSUBS 0.006021f
C559 B.n506 VSUBS 0.006021f
C560 B.n507 VSUBS 0.006021f
C561 B.n508 VSUBS 0.006021f
C562 B.n509 VSUBS 0.006021f
C563 B.n510 VSUBS 0.006021f
C564 B.n511 VSUBS 0.006021f
C565 B.n512 VSUBS 0.006021f
C566 B.n513 VSUBS 0.006021f
C567 B.n514 VSUBS 0.006021f
C568 B.n515 VSUBS 0.006021f
C569 B.n516 VSUBS 0.006021f
C570 B.n517 VSUBS 0.006021f
C571 B.n518 VSUBS 0.006021f
C572 B.n519 VSUBS 0.006021f
C573 B.n520 VSUBS 0.006021f
C574 B.n521 VSUBS 0.006021f
C575 B.n522 VSUBS 0.006021f
C576 B.n523 VSUBS 0.006021f
C577 B.n524 VSUBS 0.006021f
C578 B.n525 VSUBS 0.006021f
C579 B.n526 VSUBS 0.006021f
C580 B.n527 VSUBS 0.006021f
C581 B.n528 VSUBS 0.006021f
C582 B.n529 VSUBS 0.006021f
C583 B.n530 VSUBS 0.006021f
C584 B.n531 VSUBS 0.006021f
C585 B.n532 VSUBS 0.006021f
C586 B.n533 VSUBS 0.006021f
C587 B.n534 VSUBS 0.006021f
C588 B.n535 VSUBS 0.006021f
C589 B.n536 VSUBS 0.006021f
C590 B.n537 VSUBS 0.006021f
C591 B.n538 VSUBS 0.006021f
C592 B.n539 VSUBS 0.006021f
C593 B.n540 VSUBS 0.006021f
C594 B.n541 VSUBS 0.006021f
C595 B.n542 VSUBS 0.006021f
C596 B.n543 VSUBS 0.006021f
C597 B.n544 VSUBS 0.006021f
C598 B.n545 VSUBS 0.006021f
C599 B.n546 VSUBS 0.006021f
C600 B.n547 VSUBS 0.006021f
C601 B.n548 VSUBS 0.006021f
C602 B.n549 VSUBS 0.006021f
C603 B.n550 VSUBS 0.006021f
C604 B.n551 VSUBS 0.006021f
C605 B.n552 VSUBS 0.006021f
C606 B.n553 VSUBS 0.006021f
C607 B.n554 VSUBS 0.006021f
C608 B.n555 VSUBS 0.006021f
C609 B.n556 VSUBS 0.006021f
C610 B.n557 VSUBS 0.006021f
C611 B.n558 VSUBS 0.006021f
C612 B.n559 VSUBS 0.006021f
C613 B.n560 VSUBS 0.006021f
C614 B.n561 VSUBS 0.006021f
C615 B.n562 VSUBS 0.006021f
C616 B.n563 VSUBS 0.006021f
C617 B.n564 VSUBS 0.006021f
C618 B.n565 VSUBS 0.006021f
C619 B.n566 VSUBS 0.006021f
C620 B.n567 VSUBS 0.006021f
C621 B.n568 VSUBS 0.006021f
C622 B.n569 VSUBS 0.006021f
C623 B.n570 VSUBS 0.006021f
C624 B.n571 VSUBS 0.006021f
C625 B.n572 VSUBS 0.006021f
C626 B.n573 VSUBS 0.006021f
C627 B.n574 VSUBS 0.006021f
C628 B.n575 VSUBS 0.006021f
C629 B.n576 VSUBS 0.006021f
C630 B.n577 VSUBS 0.006021f
C631 B.n578 VSUBS 0.006021f
C632 B.n579 VSUBS 0.006021f
C633 B.n580 VSUBS 0.006021f
C634 B.n581 VSUBS 0.006021f
C635 B.n582 VSUBS 0.006021f
C636 B.n583 VSUBS 0.006021f
C637 B.n584 VSUBS 0.006021f
C638 B.n585 VSUBS 0.006021f
C639 B.n586 VSUBS 0.006021f
C640 B.n587 VSUBS 0.006021f
C641 B.n588 VSUBS 0.006021f
C642 B.n589 VSUBS 0.006021f
C643 B.n590 VSUBS 0.006021f
C644 B.n591 VSUBS 0.006021f
C645 B.n592 VSUBS 0.006021f
C646 B.n593 VSUBS 0.006021f
C647 B.n594 VSUBS 0.006021f
C648 B.n595 VSUBS 0.006021f
C649 B.n596 VSUBS 0.006021f
C650 B.n597 VSUBS 0.006021f
C651 B.n598 VSUBS 0.006021f
C652 B.n599 VSUBS 0.006021f
C653 B.n600 VSUBS 0.006021f
C654 B.n601 VSUBS 0.006021f
C655 B.n602 VSUBS 0.006021f
C656 B.n603 VSUBS 0.006021f
C657 B.n604 VSUBS 0.006021f
C658 B.n605 VSUBS 0.006021f
C659 B.n606 VSUBS 0.006021f
C660 B.n607 VSUBS 0.006021f
C661 B.n608 VSUBS 0.006021f
C662 B.n609 VSUBS 0.006021f
C663 B.n610 VSUBS 0.006021f
C664 B.n611 VSUBS 0.006021f
C665 B.n612 VSUBS 0.006021f
C666 B.n613 VSUBS 0.006021f
C667 B.n614 VSUBS 0.006021f
C668 B.n615 VSUBS 0.006021f
C669 B.n616 VSUBS 0.006021f
C670 B.n617 VSUBS 0.006021f
C671 B.n618 VSUBS 0.006021f
C672 B.n619 VSUBS 0.006021f
C673 B.n620 VSUBS 0.006021f
C674 B.n621 VSUBS 0.014124f
C675 B.n622 VSUBS 0.013681f
C676 B.n623 VSUBS 0.014407f
C677 B.n624 VSUBS 0.006021f
C678 B.n625 VSUBS 0.006021f
C679 B.n626 VSUBS 0.006021f
C680 B.n627 VSUBS 0.006021f
C681 B.n628 VSUBS 0.006021f
C682 B.n629 VSUBS 0.006021f
C683 B.n630 VSUBS 0.006021f
C684 B.n631 VSUBS 0.006021f
C685 B.n632 VSUBS 0.006021f
C686 B.n633 VSUBS 0.006021f
C687 B.n634 VSUBS 0.006021f
C688 B.n635 VSUBS 0.006021f
C689 B.n636 VSUBS 0.006021f
C690 B.n637 VSUBS 0.006021f
C691 B.n638 VSUBS 0.006021f
C692 B.n639 VSUBS 0.006021f
C693 B.n640 VSUBS 0.006021f
C694 B.n641 VSUBS 0.006021f
C695 B.n642 VSUBS 0.006021f
C696 B.n643 VSUBS 0.006021f
C697 B.n644 VSUBS 0.006021f
C698 B.n645 VSUBS 0.006021f
C699 B.n646 VSUBS 0.006021f
C700 B.n647 VSUBS 0.006021f
C701 B.n648 VSUBS 0.006021f
C702 B.n649 VSUBS 0.006021f
C703 B.n650 VSUBS 0.006021f
C704 B.n651 VSUBS 0.006021f
C705 B.n652 VSUBS 0.006021f
C706 B.n653 VSUBS 0.006021f
C707 B.n654 VSUBS 0.006021f
C708 B.n655 VSUBS 0.006021f
C709 B.n656 VSUBS 0.006021f
C710 B.n657 VSUBS 0.006021f
C711 B.n658 VSUBS 0.006021f
C712 B.n659 VSUBS 0.006021f
C713 B.n660 VSUBS 0.006021f
C714 B.n661 VSUBS 0.006021f
C715 B.n662 VSUBS 0.006021f
C716 B.n663 VSUBS 0.006021f
C717 B.n664 VSUBS 0.006021f
C718 B.n665 VSUBS 0.006021f
C719 B.n666 VSUBS 0.006021f
C720 B.n667 VSUBS 0.006021f
C721 B.n668 VSUBS 0.006021f
C722 B.n669 VSUBS 0.006021f
C723 B.n670 VSUBS 0.006021f
C724 B.n671 VSUBS 0.006021f
C725 B.n672 VSUBS 0.006021f
C726 B.n673 VSUBS 0.006021f
C727 B.n674 VSUBS 0.006021f
C728 B.n675 VSUBS 0.006021f
C729 B.n676 VSUBS 0.006021f
C730 B.n677 VSUBS 0.006021f
C731 B.n678 VSUBS 0.006021f
C732 B.n679 VSUBS 0.006021f
C733 B.n680 VSUBS 0.006021f
C734 B.n681 VSUBS 0.006021f
C735 B.n682 VSUBS 0.006021f
C736 B.n683 VSUBS 0.006021f
C737 B.n684 VSUBS 0.006021f
C738 B.n685 VSUBS 0.006021f
C739 B.n686 VSUBS 0.006021f
C740 B.n687 VSUBS 0.006021f
C741 B.n688 VSUBS 0.006021f
C742 B.n689 VSUBS 0.006021f
C743 B.n690 VSUBS 0.006021f
C744 B.n691 VSUBS 0.006021f
C745 B.n692 VSUBS 0.006021f
C746 B.n693 VSUBS 0.006021f
C747 B.n694 VSUBS 0.006021f
C748 B.n695 VSUBS 0.006021f
C749 B.n696 VSUBS 0.006021f
C750 B.n697 VSUBS 0.006021f
C751 B.n698 VSUBS 0.006021f
C752 B.n699 VSUBS 0.006021f
C753 B.n700 VSUBS 0.006021f
C754 B.n701 VSUBS 0.006021f
C755 B.n702 VSUBS 0.006021f
C756 B.n703 VSUBS 0.006021f
C757 B.n704 VSUBS 0.006021f
C758 B.n705 VSUBS 0.006021f
C759 B.n706 VSUBS 0.006021f
C760 B.n707 VSUBS 0.006021f
C761 B.n708 VSUBS 0.006021f
C762 B.n709 VSUBS 0.006021f
C763 B.n710 VSUBS 0.006021f
C764 B.n711 VSUBS 0.006021f
C765 B.n712 VSUBS 0.006021f
C766 B.n713 VSUBS 0.006021f
C767 B.n714 VSUBS 0.006021f
C768 B.n715 VSUBS 0.006021f
C769 B.n716 VSUBS 0.006021f
C770 B.n717 VSUBS 0.004162f
C771 B.n718 VSUBS 0.013951f
C772 B.n719 VSUBS 0.00487f
C773 B.n720 VSUBS 0.006021f
C774 B.n721 VSUBS 0.006021f
C775 B.n722 VSUBS 0.006021f
C776 B.n723 VSUBS 0.006021f
C777 B.n724 VSUBS 0.006021f
C778 B.n725 VSUBS 0.006021f
C779 B.n726 VSUBS 0.006021f
C780 B.n727 VSUBS 0.006021f
C781 B.n728 VSUBS 0.006021f
C782 B.n729 VSUBS 0.006021f
C783 B.n730 VSUBS 0.006021f
C784 B.n731 VSUBS 0.00487f
C785 B.n732 VSUBS 0.006021f
C786 B.n733 VSUBS 0.006021f
C787 B.n734 VSUBS 0.006021f
C788 B.n735 VSUBS 0.006021f
C789 B.n736 VSUBS 0.006021f
C790 B.n737 VSUBS 0.006021f
C791 B.n738 VSUBS 0.006021f
C792 B.n739 VSUBS 0.006021f
C793 B.n740 VSUBS 0.006021f
C794 B.n741 VSUBS 0.006021f
C795 B.n742 VSUBS 0.006021f
C796 B.n743 VSUBS 0.006021f
C797 B.n744 VSUBS 0.006021f
C798 B.n745 VSUBS 0.006021f
C799 B.n746 VSUBS 0.006021f
C800 B.n747 VSUBS 0.006021f
C801 B.n748 VSUBS 0.006021f
C802 B.n749 VSUBS 0.006021f
C803 B.n750 VSUBS 0.006021f
C804 B.n751 VSUBS 0.006021f
C805 B.n752 VSUBS 0.006021f
C806 B.n753 VSUBS 0.006021f
C807 B.n754 VSUBS 0.006021f
C808 B.n755 VSUBS 0.006021f
C809 B.n756 VSUBS 0.006021f
C810 B.n757 VSUBS 0.006021f
C811 B.n758 VSUBS 0.006021f
C812 B.n759 VSUBS 0.006021f
C813 B.n760 VSUBS 0.006021f
C814 B.n761 VSUBS 0.006021f
C815 B.n762 VSUBS 0.006021f
C816 B.n763 VSUBS 0.006021f
C817 B.n764 VSUBS 0.006021f
C818 B.n765 VSUBS 0.006021f
C819 B.n766 VSUBS 0.006021f
C820 B.n767 VSUBS 0.006021f
C821 B.n768 VSUBS 0.006021f
C822 B.n769 VSUBS 0.006021f
C823 B.n770 VSUBS 0.006021f
C824 B.n771 VSUBS 0.006021f
C825 B.n772 VSUBS 0.006021f
C826 B.n773 VSUBS 0.006021f
C827 B.n774 VSUBS 0.006021f
C828 B.n775 VSUBS 0.006021f
C829 B.n776 VSUBS 0.006021f
C830 B.n777 VSUBS 0.006021f
C831 B.n778 VSUBS 0.006021f
C832 B.n779 VSUBS 0.006021f
C833 B.n780 VSUBS 0.006021f
C834 B.n781 VSUBS 0.006021f
C835 B.n782 VSUBS 0.006021f
C836 B.n783 VSUBS 0.006021f
C837 B.n784 VSUBS 0.006021f
C838 B.n785 VSUBS 0.006021f
C839 B.n786 VSUBS 0.006021f
C840 B.n787 VSUBS 0.006021f
C841 B.n788 VSUBS 0.006021f
C842 B.n789 VSUBS 0.006021f
C843 B.n790 VSUBS 0.006021f
C844 B.n791 VSUBS 0.006021f
C845 B.n792 VSUBS 0.006021f
C846 B.n793 VSUBS 0.006021f
C847 B.n794 VSUBS 0.006021f
C848 B.n795 VSUBS 0.006021f
C849 B.n796 VSUBS 0.006021f
C850 B.n797 VSUBS 0.006021f
C851 B.n798 VSUBS 0.006021f
C852 B.n799 VSUBS 0.006021f
C853 B.n800 VSUBS 0.006021f
C854 B.n801 VSUBS 0.006021f
C855 B.n802 VSUBS 0.006021f
C856 B.n803 VSUBS 0.006021f
C857 B.n804 VSUBS 0.006021f
C858 B.n805 VSUBS 0.006021f
C859 B.n806 VSUBS 0.006021f
C860 B.n807 VSUBS 0.006021f
C861 B.n808 VSUBS 0.006021f
C862 B.n809 VSUBS 0.006021f
C863 B.n810 VSUBS 0.006021f
C864 B.n811 VSUBS 0.006021f
C865 B.n812 VSUBS 0.006021f
C866 B.n813 VSUBS 0.006021f
C867 B.n814 VSUBS 0.006021f
C868 B.n815 VSUBS 0.006021f
C869 B.n816 VSUBS 0.006021f
C870 B.n817 VSUBS 0.006021f
C871 B.n818 VSUBS 0.006021f
C872 B.n819 VSUBS 0.006021f
C873 B.n820 VSUBS 0.006021f
C874 B.n821 VSUBS 0.006021f
C875 B.n822 VSUBS 0.006021f
C876 B.n823 VSUBS 0.006021f
C877 B.n824 VSUBS 0.006021f
C878 B.n825 VSUBS 0.006021f
C879 B.n826 VSUBS 0.006021f
C880 B.n827 VSUBS 0.014407f
C881 B.n828 VSUBS 0.014407f
C882 B.n829 VSUBS 0.013397f
C883 B.n830 VSUBS 0.006021f
C884 B.n831 VSUBS 0.006021f
C885 B.n832 VSUBS 0.006021f
C886 B.n833 VSUBS 0.006021f
C887 B.n834 VSUBS 0.006021f
C888 B.n835 VSUBS 0.006021f
C889 B.n836 VSUBS 0.006021f
C890 B.n837 VSUBS 0.006021f
C891 B.n838 VSUBS 0.006021f
C892 B.n839 VSUBS 0.006021f
C893 B.n840 VSUBS 0.006021f
C894 B.n841 VSUBS 0.006021f
C895 B.n842 VSUBS 0.006021f
C896 B.n843 VSUBS 0.006021f
C897 B.n844 VSUBS 0.006021f
C898 B.n845 VSUBS 0.006021f
C899 B.n846 VSUBS 0.006021f
C900 B.n847 VSUBS 0.006021f
C901 B.n848 VSUBS 0.006021f
C902 B.n849 VSUBS 0.006021f
C903 B.n850 VSUBS 0.006021f
C904 B.n851 VSUBS 0.006021f
C905 B.n852 VSUBS 0.006021f
C906 B.n853 VSUBS 0.006021f
C907 B.n854 VSUBS 0.006021f
C908 B.n855 VSUBS 0.006021f
C909 B.n856 VSUBS 0.006021f
C910 B.n857 VSUBS 0.006021f
C911 B.n858 VSUBS 0.006021f
C912 B.n859 VSUBS 0.006021f
C913 B.n860 VSUBS 0.006021f
C914 B.n861 VSUBS 0.006021f
C915 B.n862 VSUBS 0.006021f
C916 B.n863 VSUBS 0.006021f
C917 B.n864 VSUBS 0.006021f
C918 B.n865 VSUBS 0.006021f
C919 B.n866 VSUBS 0.006021f
C920 B.n867 VSUBS 0.006021f
C921 B.n868 VSUBS 0.006021f
C922 B.n869 VSUBS 0.006021f
C923 B.n870 VSUBS 0.006021f
C924 B.n871 VSUBS 0.006021f
C925 B.n872 VSUBS 0.006021f
C926 B.n873 VSUBS 0.006021f
C927 B.n874 VSUBS 0.006021f
C928 B.n875 VSUBS 0.006021f
C929 B.n876 VSUBS 0.006021f
C930 B.n877 VSUBS 0.006021f
C931 B.n878 VSUBS 0.006021f
C932 B.n879 VSUBS 0.006021f
C933 B.n880 VSUBS 0.006021f
C934 B.n881 VSUBS 0.006021f
C935 B.n882 VSUBS 0.006021f
C936 B.n883 VSUBS 0.006021f
C937 B.n884 VSUBS 0.006021f
C938 B.n885 VSUBS 0.006021f
C939 B.n886 VSUBS 0.006021f
C940 B.n887 VSUBS 0.006021f
C941 B.n888 VSUBS 0.006021f
C942 B.n889 VSUBS 0.006021f
C943 B.n890 VSUBS 0.006021f
C944 B.n891 VSUBS 0.013634f
C945 VTAIL.n0 VSUBS 0.023972f
C946 VTAIL.n1 VSUBS 0.02238f
C947 VTAIL.n2 VSUBS 0.012026f
C948 VTAIL.n3 VSUBS 0.028426f
C949 VTAIL.n4 VSUBS 0.012734f
C950 VTAIL.n5 VSUBS 0.02238f
C951 VTAIL.n6 VSUBS 0.012026f
C952 VTAIL.n7 VSUBS 0.028426f
C953 VTAIL.n8 VSUBS 0.012734f
C954 VTAIL.n9 VSUBS 0.02238f
C955 VTAIL.n10 VSUBS 0.012026f
C956 VTAIL.n11 VSUBS 0.028426f
C957 VTAIL.n12 VSUBS 0.012734f
C958 VTAIL.n13 VSUBS 0.02238f
C959 VTAIL.n14 VSUBS 0.012026f
C960 VTAIL.n15 VSUBS 0.028426f
C961 VTAIL.n16 VSUBS 0.012734f
C962 VTAIL.n17 VSUBS 0.02238f
C963 VTAIL.n18 VSUBS 0.012026f
C964 VTAIL.n19 VSUBS 0.028426f
C965 VTAIL.n20 VSUBS 0.012734f
C966 VTAIL.n21 VSUBS 0.02238f
C967 VTAIL.n22 VSUBS 0.012026f
C968 VTAIL.n23 VSUBS 0.028426f
C969 VTAIL.n24 VSUBS 0.012734f
C970 VTAIL.n25 VSUBS 0.02238f
C971 VTAIL.n26 VSUBS 0.012026f
C972 VTAIL.n27 VSUBS 0.028426f
C973 VTAIL.n28 VSUBS 0.012734f
C974 VTAIL.n29 VSUBS 0.02238f
C975 VTAIL.n30 VSUBS 0.012026f
C976 VTAIL.n31 VSUBS 0.028426f
C977 VTAIL.n32 VSUBS 0.012734f
C978 VTAIL.n33 VSUBS 0.251749f
C979 VTAIL.t1 VSUBS 0.061818f
C980 VTAIL.n34 VSUBS 0.021319f
C981 VTAIL.n35 VSUBS 0.021383f
C982 VTAIL.n36 VSUBS 0.012026f
C983 VTAIL.n37 VSUBS 1.83116f
C984 VTAIL.n38 VSUBS 0.02238f
C985 VTAIL.n39 VSUBS 0.012026f
C986 VTAIL.n40 VSUBS 0.012734f
C987 VTAIL.n41 VSUBS 0.028426f
C988 VTAIL.n42 VSUBS 0.028426f
C989 VTAIL.n43 VSUBS 0.012734f
C990 VTAIL.n44 VSUBS 0.012026f
C991 VTAIL.n45 VSUBS 0.02238f
C992 VTAIL.n46 VSUBS 0.02238f
C993 VTAIL.n47 VSUBS 0.012026f
C994 VTAIL.n48 VSUBS 0.012734f
C995 VTAIL.n49 VSUBS 0.028426f
C996 VTAIL.n50 VSUBS 0.028426f
C997 VTAIL.n51 VSUBS 0.028426f
C998 VTAIL.n52 VSUBS 0.012734f
C999 VTAIL.n53 VSUBS 0.012026f
C1000 VTAIL.n54 VSUBS 0.02238f
C1001 VTAIL.n55 VSUBS 0.02238f
C1002 VTAIL.n56 VSUBS 0.012026f
C1003 VTAIL.n57 VSUBS 0.01238f
C1004 VTAIL.n58 VSUBS 0.01238f
C1005 VTAIL.n59 VSUBS 0.028426f
C1006 VTAIL.n60 VSUBS 0.028426f
C1007 VTAIL.n61 VSUBS 0.012734f
C1008 VTAIL.n62 VSUBS 0.012026f
C1009 VTAIL.n63 VSUBS 0.02238f
C1010 VTAIL.n64 VSUBS 0.02238f
C1011 VTAIL.n65 VSUBS 0.012026f
C1012 VTAIL.n66 VSUBS 0.012734f
C1013 VTAIL.n67 VSUBS 0.028426f
C1014 VTAIL.n68 VSUBS 0.028426f
C1015 VTAIL.n69 VSUBS 0.012734f
C1016 VTAIL.n70 VSUBS 0.012026f
C1017 VTAIL.n71 VSUBS 0.02238f
C1018 VTAIL.n72 VSUBS 0.02238f
C1019 VTAIL.n73 VSUBS 0.012026f
C1020 VTAIL.n74 VSUBS 0.012734f
C1021 VTAIL.n75 VSUBS 0.028426f
C1022 VTAIL.n76 VSUBS 0.028426f
C1023 VTAIL.n77 VSUBS 0.012734f
C1024 VTAIL.n78 VSUBS 0.012026f
C1025 VTAIL.n79 VSUBS 0.02238f
C1026 VTAIL.n80 VSUBS 0.02238f
C1027 VTAIL.n81 VSUBS 0.012026f
C1028 VTAIL.n82 VSUBS 0.012734f
C1029 VTAIL.n83 VSUBS 0.028426f
C1030 VTAIL.n84 VSUBS 0.028426f
C1031 VTAIL.n85 VSUBS 0.012734f
C1032 VTAIL.n86 VSUBS 0.012026f
C1033 VTAIL.n87 VSUBS 0.02238f
C1034 VTAIL.n88 VSUBS 0.02238f
C1035 VTAIL.n89 VSUBS 0.012026f
C1036 VTAIL.n90 VSUBS 0.012734f
C1037 VTAIL.n91 VSUBS 0.028426f
C1038 VTAIL.n92 VSUBS 0.028426f
C1039 VTAIL.n93 VSUBS 0.012734f
C1040 VTAIL.n94 VSUBS 0.012026f
C1041 VTAIL.n95 VSUBS 0.02238f
C1042 VTAIL.n96 VSUBS 0.02238f
C1043 VTAIL.n97 VSUBS 0.012026f
C1044 VTAIL.n98 VSUBS 0.012734f
C1045 VTAIL.n99 VSUBS 0.028426f
C1046 VTAIL.n100 VSUBS 0.070357f
C1047 VTAIL.n101 VSUBS 0.012734f
C1048 VTAIL.n102 VSUBS 0.023617f
C1049 VTAIL.n103 VSUBS 0.056011f
C1050 VTAIL.n104 VSUBS 0.053757f
C1051 VTAIL.n105 VSUBS 0.175866f
C1052 VTAIL.n106 VSUBS 0.023972f
C1053 VTAIL.n107 VSUBS 0.02238f
C1054 VTAIL.n108 VSUBS 0.012026f
C1055 VTAIL.n109 VSUBS 0.028426f
C1056 VTAIL.n110 VSUBS 0.012734f
C1057 VTAIL.n111 VSUBS 0.02238f
C1058 VTAIL.n112 VSUBS 0.012026f
C1059 VTAIL.n113 VSUBS 0.028426f
C1060 VTAIL.n114 VSUBS 0.012734f
C1061 VTAIL.n115 VSUBS 0.02238f
C1062 VTAIL.n116 VSUBS 0.012026f
C1063 VTAIL.n117 VSUBS 0.028426f
C1064 VTAIL.n118 VSUBS 0.012734f
C1065 VTAIL.n119 VSUBS 0.02238f
C1066 VTAIL.n120 VSUBS 0.012026f
C1067 VTAIL.n121 VSUBS 0.028426f
C1068 VTAIL.n122 VSUBS 0.012734f
C1069 VTAIL.n123 VSUBS 0.02238f
C1070 VTAIL.n124 VSUBS 0.012026f
C1071 VTAIL.n125 VSUBS 0.028426f
C1072 VTAIL.n126 VSUBS 0.012734f
C1073 VTAIL.n127 VSUBS 0.02238f
C1074 VTAIL.n128 VSUBS 0.012026f
C1075 VTAIL.n129 VSUBS 0.028426f
C1076 VTAIL.n130 VSUBS 0.012734f
C1077 VTAIL.n131 VSUBS 0.02238f
C1078 VTAIL.n132 VSUBS 0.012026f
C1079 VTAIL.n133 VSUBS 0.028426f
C1080 VTAIL.n134 VSUBS 0.012734f
C1081 VTAIL.n135 VSUBS 0.02238f
C1082 VTAIL.n136 VSUBS 0.012026f
C1083 VTAIL.n137 VSUBS 0.028426f
C1084 VTAIL.n138 VSUBS 0.012734f
C1085 VTAIL.n139 VSUBS 0.251749f
C1086 VTAIL.t6 VSUBS 0.061818f
C1087 VTAIL.n140 VSUBS 0.021319f
C1088 VTAIL.n141 VSUBS 0.021383f
C1089 VTAIL.n142 VSUBS 0.012026f
C1090 VTAIL.n143 VSUBS 1.83116f
C1091 VTAIL.n144 VSUBS 0.02238f
C1092 VTAIL.n145 VSUBS 0.012026f
C1093 VTAIL.n146 VSUBS 0.012734f
C1094 VTAIL.n147 VSUBS 0.028426f
C1095 VTAIL.n148 VSUBS 0.028426f
C1096 VTAIL.n149 VSUBS 0.012734f
C1097 VTAIL.n150 VSUBS 0.012026f
C1098 VTAIL.n151 VSUBS 0.02238f
C1099 VTAIL.n152 VSUBS 0.02238f
C1100 VTAIL.n153 VSUBS 0.012026f
C1101 VTAIL.n154 VSUBS 0.012734f
C1102 VTAIL.n155 VSUBS 0.028426f
C1103 VTAIL.n156 VSUBS 0.028426f
C1104 VTAIL.n157 VSUBS 0.028426f
C1105 VTAIL.n158 VSUBS 0.012734f
C1106 VTAIL.n159 VSUBS 0.012026f
C1107 VTAIL.n160 VSUBS 0.02238f
C1108 VTAIL.n161 VSUBS 0.02238f
C1109 VTAIL.n162 VSUBS 0.012026f
C1110 VTAIL.n163 VSUBS 0.01238f
C1111 VTAIL.n164 VSUBS 0.01238f
C1112 VTAIL.n165 VSUBS 0.028426f
C1113 VTAIL.n166 VSUBS 0.028426f
C1114 VTAIL.n167 VSUBS 0.012734f
C1115 VTAIL.n168 VSUBS 0.012026f
C1116 VTAIL.n169 VSUBS 0.02238f
C1117 VTAIL.n170 VSUBS 0.02238f
C1118 VTAIL.n171 VSUBS 0.012026f
C1119 VTAIL.n172 VSUBS 0.012734f
C1120 VTAIL.n173 VSUBS 0.028426f
C1121 VTAIL.n174 VSUBS 0.028426f
C1122 VTAIL.n175 VSUBS 0.012734f
C1123 VTAIL.n176 VSUBS 0.012026f
C1124 VTAIL.n177 VSUBS 0.02238f
C1125 VTAIL.n178 VSUBS 0.02238f
C1126 VTAIL.n179 VSUBS 0.012026f
C1127 VTAIL.n180 VSUBS 0.012734f
C1128 VTAIL.n181 VSUBS 0.028426f
C1129 VTAIL.n182 VSUBS 0.028426f
C1130 VTAIL.n183 VSUBS 0.012734f
C1131 VTAIL.n184 VSUBS 0.012026f
C1132 VTAIL.n185 VSUBS 0.02238f
C1133 VTAIL.n186 VSUBS 0.02238f
C1134 VTAIL.n187 VSUBS 0.012026f
C1135 VTAIL.n188 VSUBS 0.012734f
C1136 VTAIL.n189 VSUBS 0.028426f
C1137 VTAIL.n190 VSUBS 0.028426f
C1138 VTAIL.n191 VSUBS 0.012734f
C1139 VTAIL.n192 VSUBS 0.012026f
C1140 VTAIL.n193 VSUBS 0.02238f
C1141 VTAIL.n194 VSUBS 0.02238f
C1142 VTAIL.n195 VSUBS 0.012026f
C1143 VTAIL.n196 VSUBS 0.012734f
C1144 VTAIL.n197 VSUBS 0.028426f
C1145 VTAIL.n198 VSUBS 0.028426f
C1146 VTAIL.n199 VSUBS 0.012734f
C1147 VTAIL.n200 VSUBS 0.012026f
C1148 VTAIL.n201 VSUBS 0.02238f
C1149 VTAIL.n202 VSUBS 0.02238f
C1150 VTAIL.n203 VSUBS 0.012026f
C1151 VTAIL.n204 VSUBS 0.012734f
C1152 VTAIL.n205 VSUBS 0.028426f
C1153 VTAIL.n206 VSUBS 0.070357f
C1154 VTAIL.n207 VSUBS 0.012734f
C1155 VTAIL.n208 VSUBS 0.023617f
C1156 VTAIL.n209 VSUBS 0.056011f
C1157 VTAIL.n210 VSUBS 0.053757f
C1158 VTAIL.n211 VSUBS 0.287923f
C1159 VTAIL.n212 VSUBS 0.023972f
C1160 VTAIL.n213 VSUBS 0.02238f
C1161 VTAIL.n214 VSUBS 0.012026f
C1162 VTAIL.n215 VSUBS 0.028426f
C1163 VTAIL.n216 VSUBS 0.012734f
C1164 VTAIL.n217 VSUBS 0.02238f
C1165 VTAIL.n218 VSUBS 0.012026f
C1166 VTAIL.n219 VSUBS 0.028426f
C1167 VTAIL.n220 VSUBS 0.012734f
C1168 VTAIL.n221 VSUBS 0.02238f
C1169 VTAIL.n222 VSUBS 0.012026f
C1170 VTAIL.n223 VSUBS 0.028426f
C1171 VTAIL.n224 VSUBS 0.012734f
C1172 VTAIL.n225 VSUBS 0.02238f
C1173 VTAIL.n226 VSUBS 0.012026f
C1174 VTAIL.n227 VSUBS 0.028426f
C1175 VTAIL.n228 VSUBS 0.012734f
C1176 VTAIL.n229 VSUBS 0.02238f
C1177 VTAIL.n230 VSUBS 0.012026f
C1178 VTAIL.n231 VSUBS 0.028426f
C1179 VTAIL.n232 VSUBS 0.012734f
C1180 VTAIL.n233 VSUBS 0.02238f
C1181 VTAIL.n234 VSUBS 0.012026f
C1182 VTAIL.n235 VSUBS 0.028426f
C1183 VTAIL.n236 VSUBS 0.012734f
C1184 VTAIL.n237 VSUBS 0.02238f
C1185 VTAIL.n238 VSUBS 0.012026f
C1186 VTAIL.n239 VSUBS 0.028426f
C1187 VTAIL.n240 VSUBS 0.012734f
C1188 VTAIL.n241 VSUBS 0.02238f
C1189 VTAIL.n242 VSUBS 0.012026f
C1190 VTAIL.n243 VSUBS 0.028426f
C1191 VTAIL.n244 VSUBS 0.012734f
C1192 VTAIL.n245 VSUBS 0.251749f
C1193 VTAIL.t4 VSUBS 0.061818f
C1194 VTAIL.n246 VSUBS 0.021319f
C1195 VTAIL.n247 VSUBS 0.021383f
C1196 VTAIL.n248 VSUBS 0.012026f
C1197 VTAIL.n249 VSUBS 1.83116f
C1198 VTAIL.n250 VSUBS 0.02238f
C1199 VTAIL.n251 VSUBS 0.012026f
C1200 VTAIL.n252 VSUBS 0.012734f
C1201 VTAIL.n253 VSUBS 0.028426f
C1202 VTAIL.n254 VSUBS 0.028426f
C1203 VTAIL.n255 VSUBS 0.012734f
C1204 VTAIL.n256 VSUBS 0.012026f
C1205 VTAIL.n257 VSUBS 0.02238f
C1206 VTAIL.n258 VSUBS 0.02238f
C1207 VTAIL.n259 VSUBS 0.012026f
C1208 VTAIL.n260 VSUBS 0.012734f
C1209 VTAIL.n261 VSUBS 0.028426f
C1210 VTAIL.n262 VSUBS 0.028426f
C1211 VTAIL.n263 VSUBS 0.028426f
C1212 VTAIL.n264 VSUBS 0.012734f
C1213 VTAIL.n265 VSUBS 0.012026f
C1214 VTAIL.n266 VSUBS 0.02238f
C1215 VTAIL.n267 VSUBS 0.02238f
C1216 VTAIL.n268 VSUBS 0.012026f
C1217 VTAIL.n269 VSUBS 0.01238f
C1218 VTAIL.n270 VSUBS 0.01238f
C1219 VTAIL.n271 VSUBS 0.028426f
C1220 VTAIL.n272 VSUBS 0.028426f
C1221 VTAIL.n273 VSUBS 0.012734f
C1222 VTAIL.n274 VSUBS 0.012026f
C1223 VTAIL.n275 VSUBS 0.02238f
C1224 VTAIL.n276 VSUBS 0.02238f
C1225 VTAIL.n277 VSUBS 0.012026f
C1226 VTAIL.n278 VSUBS 0.012734f
C1227 VTAIL.n279 VSUBS 0.028426f
C1228 VTAIL.n280 VSUBS 0.028426f
C1229 VTAIL.n281 VSUBS 0.012734f
C1230 VTAIL.n282 VSUBS 0.012026f
C1231 VTAIL.n283 VSUBS 0.02238f
C1232 VTAIL.n284 VSUBS 0.02238f
C1233 VTAIL.n285 VSUBS 0.012026f
C1234 VTAIL.n286 VSUBS 0.012734f
C1235 VTAIL.n287 VSUBS 0.028426f
C1236 VTAIL.n288 VSUBS 0.028426f
C1237 VTAIL.n289 VSUBS 0.012734f
C1238 VTAIL.n290 VSUBS 0.012026f
C1239 VTAIL.n291 VSUBS 0.02238f
C1240 VTAIL.n292 VSUBS 0.02238f
C1241 VTAIL.n293 VSUBS 0.012026f
C1242 VTAIL.n294 VSUBS 0.012734f
C1243 VTAIL.n295 VSUBS 0.028426f
C1244 VTAIL.n296 VSUBS 0.028426f
C1245 VTAIL.n297 VSUBS 0.012734f
C1246 VTAIL.n298 VSUBS 0.012026f
C1247 VTAIL.n299 VSUBS 0.02238f
C1248 VTAIL.n300 VSUBS 0.02238f
C1249 VTAIL.n301 VSUBS 0.012026f
C1250 VTAIL.n302 VSUBS 0.012734f
C1251 VTAIL.n303 VSUBS 0.028426f
C1252 VTAIL.n304 VSUBS 0.028426f
C1253 VTAIL.n305 VSUBS 0.012734f
C1254 VTAIL.n306 VSUBS 0.012026f
C1255 VTAIL.n307 VSUBS 0.02238f
C1256 VTAIL.n308 VSUBS 0.02238f
C1257 VTAIL.n309 VSUBS 0.012026f
C1258 VTAIL.n310 VSUBS 0.012734f
C1259 VTAIL.n311 VSUBS 0.028426f
C1260 VTAIL.n312 VSUBS 0.070357f
C1261 VTAIL.n313 VSUBS 0.012734f
C1262 VTAIL.n314 VSUBS 0.023617f
C1263 VTAIL.n315 VSUBS 0.056011f
C1264 VTAIL.n316 VSUBS 0.053757f
C1265 VTAIL.n317 VSUBS 2.00034f
C1266 VTAIL.n318 VSUBS 0.023972f
C1267 VTAIL.n319 VSUBS 0.02238f
C1268 VTAIL.n320 VSUBS 0.012026f
C1269 VTAIL.n321 VSUBS 0.028426f
C1270 VTAIL.n322 VSUBS 0.012734f
C1271 VTAIL.n323 VSUBS 0.02238f
C1272 VTAIL.n324 VSUBS 0.012026f
C1273 VTAIL.n325 VSUBS 0.028426f
C1274 VTAIL.n326 VSUBS 0.012734f
C1275 VTAIL.n327 VSUBS 0.02238f
C1276 VTAIL.n328 VSUBS 0.012026f
C1277 VTAIL.n329 VSUBS 0.028426f
C1278 VTAIL.n330 VSUBS 0.012734f
C1279 VTAIL.n331 VSUBS 0.02238f
C1280 VTAIL.n332 VSUBS 0.012026f
C1281 VTAIL.n333 VSUBS 0.028426f
C1282 VTAIL.n334 VSUBS 0.012734f
C1283 VTAIL.n335 VSUBS 0.02238f
C1284 VTAIL.n336 VSUBS 0.012026f
C1285 VTAIL.n337 VSUBS 0.028426f
C1286 VTAIL.n338 VSUBS 0.012734f
C1287 VTAIL.n339 VSUBS 0.02238f
C1288 VTAIL.n340 VSUBS 0.012026f
C1289 VTAIL.n341 VSUBS 0.028426f
C1290 VTAIL.n342 VSUBS 0.012734f
C1291 VTAIL.n343 VSUBS 0.02238f
C1292 VTAIL.n344 VSUBS 0.012026f
C1293 VTAIL.n345 VSUBS 0.028426f
C1294 VTAIL.n346 VSUBS 0.028426f
C1295 VTAIL.n347 VSUBS 0.012734f
C1296 VTAIL.n348 VSUBS 0.02238f
C1297 VTAIL.n349 VSUBS 0.012026f
C1298 VTAIL.n350 VSUBS 0.028426f
C1299 VTAIL.n351 VSUBS 0.012734f
C1300 VTAIL.n352 VSUBS 0.251749f
C1301 VTAIL.t3 VSUBS 0.061818f
C1302 VTAIL.n353 VSUBS 0.021319f
C1303 VTAIL.n354 VSUBS 0.021383f
C1304 VTAIL.n355 VSUBS 0.012026f
C1305 VTAIL.n356 VSUBS 1.83116f
C1306 VTAIL.n357 VSUBS 0.02238f
C1307 VTAIL.n358 VSUBS 0.012026f
C1308 VTAIL.n359 VSUBS 0.012734f
C1309 VTAIL.n360 VSUBS 0.028426f
C1310 VTAIL.n361 VSUBS 0.028426f
C1311 VTAIL.n362 VSUBS 0.012734f
C1312 VTAIL.n363 VSUBS 0.012026f
C1313 VTAIL.n364 VSUBS 0.02238f
C1314 VTAIL.n365 VSUBS 0.02238f
C1315 VTAIL.n366 VSUBS 0.012026f
C1316 VTAIL.n367 VSUBS 0.012734f
C1317 VTAIL.n368 VSUBS 0.028426f
C1318 VTAIL.n369 VSUBS 0.028426f
C1319 VTAIL.n370 VSUBS 0.012734f
C1320 VTAIL.n371 VSUBS 0.012026f
C1321 VTAIL.n372 VSUBS 0.02238f
C1322 VTAIL.n373 VSUBS 0.02238f
C1323 VTAIL.n374 VSUBS 0.012026f
C1324 VTAIL.n375 VSUBS 0.01238f
C1325 VTAIL.n376 VSUBS 0.01238f
C1326 VTAIL.n377 VSUBS 0.028426f
C1327 VTAIL.n378 VSUBS 0.028426f
C1328 VTAIL.n379 VSUBS 0.012734f
C1329 VTAIL.n380 VSUBS 0.012026f
C1330 VTAIL.n381 VSUBS 0.02238f
C1331 VTAIL.n382 VSUBS 0.02238f
C1332 VTAIL.n383 VSUBS 0.012026f
C1333 VTAIL.n384 VSUBS 0.012734f
C1334 VTAIL.n385 VSUBS 0.028426f
C1335 VTAIL.n386 VSUBS 0.028426f
C1336 VTAIL.n387 VSUBS 0.012734f
C1337 VTAIL.n388 VSUBS 0.012026f
C1338 VTAIL.n389 VSUBS 0.02238f
C1339 VTAIL.n390 VSUBS 0.02238f
C1340 VTAIL.n391 VSUBS 0.012026f
C1341 VTAIL.n392 VSUBS 0.012734f
C1342 VTAIL.n393 VSUBS 0.028426f
C1343 VTAIL.n394 VSUBS 0.028426f
C1344 VTAIL.n395 VSUBS 0.012734f
C1345 VTAIL.n396 VSUBS 0.012026f
C1346 VTAIL.n397 VSUBS 0.02238f
C1347 VTAIL.n398 VSUBS 0.02238f
C1348 VTAIL.n399 VSUBS 0.012026f
C1349 VTAIL.n400 VSUBS 0.012734f
C1350 VTAIL.n401 VSUBS 0.028426f
C1351 VTAIL.n402 VSUBS 0.028426f
C1352 VTAIL.n403 VSUBS 0.012734f
C1353 VTAIL.n404 VSUBS 0.012026f
C1354 VTAIL.n405 VSUBS 0.02238f
C1355 VTAIL.n406 VSUBS 0.02238f
C1356 VTAIL.n407 VSUBS 0.012026f
C1357 VTAIL.n408 VSUBS 0.012734f
C1358 VTAIL.n409 VSUBS 0.028426f
C1359 VTAIL.n410 VSUBS 0.028426f
C1360 VTAIL.n411 VSUBS 0.012734f
C1361 VTAIL.n412 VSUBS 0.012026f
C1362 VTAIL.n413 VSUBS 0.02238f
C1363 VTAIL.n414 VSUBS 0.02238f
C1364 VTAIL.n415 VSUBS 0.012026f
C1365 VTAIL.n416 VSUBS 0.012734f
C1366 VTAIL.n417 VSUBS 0.028426f
C1367 VTAIL.n418 VSUBS 0.070357f
C1368 VTAIL.n419 VSUBS 0.012734f
C1369 VTAIL.n420 VSUBS 0.023617f
C1370 VTAIL.n421 VSUBS 0.056011f
C1371 VTAIL.n422 VSUBS 0.053757f
C1372 VTAIL.n423 VSUBS 2.00034f
C1373 VTAIL.n424 VSUBS 0.023972f
C1374 VTAIL.n425 VSUBS 0.02238f
C1375 VTAIL.n426 VSUBS 0.012026f
C1376 VTAIL.n427 VSUBS 0.028426f
C1377 VTAIL.n428 VSUBS 0.012734f
C1378 VTAIL.n429 VSUBS 0.02238f
C1379 VTAIL.n430 VSUBS 0.012026f
C1380 VTAIL.n431 VSUBS 0.028426f
C1381 VTAIL.n432 VSUBS 0.012734f
C1382 VTAIL.n433 VSUBS 0.02238f
C1383 VTAIL.n434 VSUBS 0.012026f
C1384 VTAIL.n435 VSUBS 0.028426f
C1385 VTAIL.n436 VSUBS 0.012734f
C1386 VTAIL.n437 VSUBS 0.02238f
C1387 VTAIL.n438 VSUBS 0.012026f
C1388 VTAIL.n439 VSUBS 0.028426f
C1389 VTAIL.n440 VSUBS 0.012734f
C1390 VTAIL.n441 VSUBS 0.02238f
C1391 VTAIL.n442 VSUBS 0.012026f
C1392 VTAIL.n443 VSUBS 0.028426f
C1393 VTAIL.n444 VSUBS 0.012734f
C1394 VTAIL.n445 VSUBS 0.02238f
C1395 VTAIL.n446 VSUBS 0.012026f
C1396 VTAIL.n447 VSUBS 0.028426f
C1397 VTAIL.n448 VSUBS 0.012734f
C1398 VTAIL.n449 VSUBS 0.02238f
C1399 VTAIL.n450 VSUBS 0.012026f
C1400 VTAIL.n451 VSUBS 0.028426f
C1401 VTAIL.n452 VSUBS 0.028426f
C1402 VTAIL.n453 VSUBS 0.012734f
C1403 VTAIL.n454 VSUBS 0.02238f
C1404 VTAIL.n455 VSUBS 0.012026f
C1405 VTAIL.n456 VSUBS 0.028426f
C1406 VTAIL.n457 VSUBS 0.012734f
C1407 VTAIL.n458 VSUBS 0.251749f
C1408 VTAIL.t0 VSUBS 0.061818f
C1409 VTAIL.n459 VSUBS 0.021319f
C1410 VTAIL.n460 VSUBS 0.021383f
C1411 VTAIL.n461 VSUBS 0.012026f
C1412 VTAIL.n462 VSUBS 1.83116f
C1413 VTAIL.n463 VSUBS 0.02238f
C1414 VTAIL.n464 VSUBS 0.012026f
C1415 VTAIL.n465 VSUBS 0.012734f
C1416 VTAIL.n466 VSUBS 0.028426f
C1417 VTAIL.n467 VSUBS 0.028426f
C1418 VTAIL.n468 VSUBS 0.012734f
C1419 VTAIL.n469 VSUBS 0.012026f
C1420 VTAIL.n470 VSUBS 0.02238f
C1421 VTAIL.n471 VSUBS 0.02238f
C1422 VTAIL.n472 VSUBS 0.012026f
C1423 VTAIL.n473 VSUBS 0.012734f
C1424 VTAIL.n474 VSUBS 0.028426f
C1425 VTAIL.n475 VSUBS 0.028426f
C1426 VTAIL.n476 VSUBS 0.012734f
C1427 VTAIL.n477 VSUBS 0.012026f
C1428 VTAIL.n478 VSUBS 0.02238f
C1429 VTAIL.n479 VSUBS 0.02238f
C1430 VTAIL.n480 VSUBS 0.012026f
C1431 VTAIL.n481 VSUBS 0.01238f
C1432 VTAIL.n482 VSUBS 0.01238f
C1433 VTAIL.n483 VSUBS 0.028426f
C1434 VTAIL.n484 VSUBS 0.028426f
C1435 VTAIL.n485 VSUBS 0.012734f
C1436 VTAIL.n486 VSUBS 0.012026f
C1437 VTAIL.n487 VSUBS 0.02238f
C1438 VTAIL.n488 VSUBS 0.02238f
C1439 VTAIL.n489 VSUBS 0.012026f
C1440 VTAIL.n490 VSUBS 0.012734f
C1441 VTAIL.n491 VSUBS 0.028426f
C1442 VTAIL.n492 VSUBS 0.028426f
C1443 VTAIL.n493 VSUBS 0.012734f
C1444 VTAIL.n494 VSUBS 0.012026f
C1445 VTAIL.n495 VSUBS 0.02238f
C1446 VTAIL.n496 VSUBS 0.02238f
C1447 VTAIL.n497 VSUBS 0.012026f
C1448 VTAIL.n498 VSUBS 0.012734f
C1449 VTAIL.n499 VSUBS 0.028426f
C1450 VTAIL.n500 VSUBS 0.028426f
C1451 VTAIL.n501 VSUBS 0.012734f
C1452 VTAIL.n502 VSUBS 0.012026f
C1453 VTAIL.n503 VSUBS 0.02238f
C1454 VTAIL.n504 VSUBS 0.02238f
C1455 VTAIL.n505 VSUBS 0.012026f
C1456 VTAIL.n506 VSUBS 0.012734f
C1457 VTAIL.n507 VSUBS 0.028426f
C1458 VTAIL.n508 VSUBS 0.028426f
C1459 VTAIL.n509 VSUBS 0.012734f
C1460 VTAIL.n510 VSUBS 0.012026f
C1461 VTAIL.n511 VSUBS 0.02238f
C1462 VTAIL.n512 VSUBS 0.02238f
C1463 VTAIL.n513 VSUBS 0.012026f
C1464 VTAIL.n514 VSUBS 0.012734f
C1465 VTAIL.n515 VSUBS 0.028426f
C1466 VTAIL.n516 VSUBS 0.028426f
C1467 VTAIL.n517 VSUBS 0.012734f
C1468 VTAIL.n518 VSUBS 0.012026f
C1469 VTAIL.n519 VSUBS 0.02238f
C1470 VTAIL.n520 VSUBS 0.02238f
C1471 VTAIL.n521 VSUBS 0.012026f
C1472 VTAIL.n522 VSUBS 0.012734f
C1473 VTAIL.n523 VSUBS 0.028426f
C1474 VTAIL.n524 VSUBS 0.070357f
C1475 VTAIL.n525 VSUBS 0.012734f
C1476 VTAIL.n526 VSUBS 0.023617f
C1477 VTAIL.n527 VSUBS 0.056011f
C1478 VTAIL.n528 VSUBS 0.053757f
C1479 VTAIL.n529 VSUBS 0.287923f
C1480 VTAIL.n530 VSUBS 0.023972f
C1481 VTAIL.n531 VSUBS 0.02238f
C1482 VTAIL.n532 VSUBS 0.012026f
C1483 VTAIL.n533 VSUBS 0.028426f
C1484 VTAIL.n534 VSUBS 0.012734f
C1485 VTAIL.n535 VSUBS 0.02238f
C1486 VTAIL.n536 VSUBS 0.012026f
C1487 VTAIL.n537 VSUBS 0.028426f
C1488 VTAIL.n538 VSUBS 0.012734f
C1489 VTAIL.n539 VSUBS 0.02238f
C1490 VTAIL.n540 VSUBS 0.012026f
C1491 VTAIL.n541 VSUBS 0.028426f
C1492 VTAIL.n542 VSUBS 0.012734f
C1493 VTAIL.n543 VSUBS 0.02238f
C1494 VTAIL.n544 VSUBS 0.012026f
C1495 VTAIL.n545 VSUBS 0.028426f
C1496 VTAIL.n546 VSUBS 0.012734f
C1497 VTAIL.n547 VSUBS 0.02238f
C1498 VTAIL.n548 VSUBS 0.012026f
C1499 VTAIL.n549 VSUBS 0.028426f
C1500 VTAIL.n550 VSUBS 0.012734f
C1501 VTAIL.n551 VSUBS 0.02238f
C1502 VTAIL.n552 VSUBS 0.012026f
C1503 VTAIL.n553 VSUBS 0.028426f
C1504 VTAIL.n554 VSUBS 0.012734f
C1505 VTAIL.n555 VSUBS 0.02238f
C1506 VTAIL.n556 VSUBS 0.012026f
C1507 VTAIL.n557 VSUBS 0.028426f
C1508 VTAIL.n558 VSUBS 0.028426f
C1509 VTAIL.n559 VSUBS 0.012734f
C1510 VTAIL.n560 VSUBS 0.02238f
C1511 VTAIL.n561 VSUBS 0.012026f
C1512 VTAIL.n562 VSUBS 0.028426f
C1513 VTAIL.n563 VSUBS 0.012734f
C1514 VTAIL.n564 VSUBS 0.251749f
C1515 VTAIL.t7 VSUBS 0.061818f
C1516 VTAIL.n565 VSUBS 0.021319f
C1517 VTAIL.n566 VSUBS 0.021383f
C1518 VTAIL.n567 VSUBS 0.012026f
C1519 VTAIL.n568 VSUBS 1.83116f
C1520 VTAIL.n569 VSUBS 0.02238f
C1521 VTAIL.n570 VSUBS 0.012026f
C1522 VTAIL.n571 VSUBS 0.012734f
C1523 VTAIL.n572 VSUBS 0.028426f
C1524 VTAIL.n573 VSUBS 0.028426f
C1525 VTAIL.n574 VSUBS 0.012734f
C1526 VTAIL.n575 VSUBS 0.012026f
C1527 VTAIL.n576 VSUBS 0.02238f
C1528 VTAIL.n577 VSUBS 0.02238f
C1529 VTAIL.n578 VSUBS 0.012026f
C1530 VTAIL.n579 VSUBS 0.012734f
C1531 VTAIL.n580 VSUBS 0.028426f
C1532 VTAIL.n581 VSUBS 0.028426f
C1533 VTAIL.n582 VSUBS 0.012734f
C1534 VTAIL.n583 VSUBS 0.012026f
C1535 VTAIL.n584 VSUBS 0.02238f
C1536 VTAIL.n585 VSUBS 0.02238f
C1537 VTAIL.n586 VSUBS 0.012026f
C1538 VTAIL.n587 VSUBS 0.01238f
C1539 VTAIL.n588 VSUBS 0.01238f
C1540 VTAIL.n589 VSUBS 0.028426f
C1541 VTAIL.n590 VSUBS 0.028426f
C1542 VTAIL.n591 VSUBS 0.012734f
C1543 VTAIL.n592 VSUBS 0.012026f
C1544 VTAIL.n593 VSUBS 0.02238f
C1545 VTAIL.n594 VSUBS 0.02238f
C1546 VTAIL.n595 VSUBS 0.012026f
C1547 VTAIL.n596 VSUBS 0.012734f
C1548 VTAIL.n597 VSUBS 0.028426f
C1549 VTAIL.n598 VSUBS 0.028426f
C1550 VTAIL.n599 VSUBS 0.012734f
C1551 VTAIL.n600 VSUBS 0.012026f
C1552 VTAIL.n601 VSUBS 0.02238f
C1553 VTAIL.n602 VSUBS 0.02238f
C1554 VTAIL.n603 VSUBS 0.012026f
C1555 VTAIL.n604 VSUBS 0.012734f
C1556 VTAIL.n605 VSUBS 0.028426f
C1557 VTAIL.n606 VSUBS 0.028426f
C1558 VTAIL.n607 VSUBS 0.012734f
C1559 VTAIL.n608 VSUBS 0.012026f
C1560 VTAIL.n609 VSUBS 0.02238f
C1561 VTAIL.n610 VSUBS 0.02238f
C1562 VTAIL.n611 VSUBS 0.012026f
C1563 VTAIL.n612 VSUBS 0.012734f
C1564 VTAIL.n613 VSUBS 0.028426f
C1565 VTAIL.n614 VSUBS 0.028426f
C1566 VTAIL.n615 VSUBS 0.012734f
C1567 VTAIL.n616 VSUBS 0.012026f
C1568 VTAIL.n617 VSUBS 0.02238f
C1569 VTAIL.n618 VSUBS 0.02238f
C1570 VTAIL.n619 VSUBS 0.012026f
C1571 VTAIL.n620 VSUBS 0.012734f
C1572 VTAIL.n621 VSUBS 0.028426f
C1573 VTAIL.n622 VSUBS 0.028426f
C1574 VTAIL.n623 VSUBS 0.012734f
C1575 VTAIL.n624 VSUBS 0.012026f
C1576 VTAIL.n625 VSUBS 0.02238f
C1577 VTAIL.n626 VSUBS 0.02238f
C1578 VTAIL.n627 VSUBS 0.012026f
C1579 VTAIL.n628 VSUBS 0.012734f
C1580 VTAIL.n629 VSUBS 0.028426f
C1581 VTAIL.n630 VSUBS 0.070357f
C1582 VTAIL.n631 VSUBS 0.012734f
C1583 VTAIL.n632 VSUBS 0.023617f
C1584 VTAIL.n633 VSUBS 0.056011f
C1585 VTAIL.n634 VSUBS 0.053757f
C1586 VTAIL.n635 VSUBS 0.287923f
C1587 VTAIL.n636 VSUBS 0.023972f
C1588 VTAIL.n637 VSUBS 0.02238f
C1589 VTAIL.n638 VSUBS 0.012026f
C1590 VTAIL.n639 VSUBS 0.028426f
C1591 VTAIL.n640 VSUBS 0.012734f
C1592 VTAIL.n641 VSUBS 0.02238f
C1593 VTAIL.n642 VSUBS 0.012026f
C1594 VTAIL.n643 VSUBS 0.028426f
C1595 VTAIL.n644 VSUBS 0.012734f
C1596 VTAIL.n645 VSUBS 0.02238f
C1597 VTAIL.n646 VSUBS 0.012026f
C1598 VTAIL.n647 VSUBS 0.028426f
C1599 VTAIL.n648 VSUBS 0.012734f
C1600 VTAIL.n649 VSUBS 0.02238f
C1601 VTAIL.n650 VSUBS 0.012026f
C1602 VTAIL.n651 VSUBS 0.028426f
C1603 VTAIL.n652 VSUBS 0.012734f
C1604 VTAIL.n653 VSUBS 0.02238f
C1605 VTAIL.n654 VSUBS 0.012026f
C1606 VTAIL.n655 VSUBS 0.028426f
C1607 VTAIL.n656 VSUBS 0.012734f
C1608 VTAIL.n657 VSUBS 0.02238f
C1609 VTAIL.n658 VSUBS 0.012026f
C1610 VTAIL.n659 VSUBS 0.028426f
C1611 VTAIL.n660 VSUBS 0.012734f
C1612 VTAIL.n661 VSUBS 0.02238f
C1613 VTAIL.n662 VSUBS 0.012026f
C1614 VTAIL.n663 VSUBS 0.028426f
C1615 VTAIL.n664 VSUBS 0.028426f
C1616 VTAIL.n665 VSUBS 0.012734f
C1617 VTAIL.n666 VSUBS 0.02238f
C1618 VTAIL.n667 VSUBS 0.012026f
C1619 VTAIL.n668 VSUBS 0.028426f
C1620 VTAIL.n669 VSUBS 0.012734f
C1621 VTAIL.n670 VSUBS 0.251749f
C1622 VTAIL.t5 VSUBS 0.061818f
C1623 VTAIL.n671 VSUBS 0.021319f
C1624 VTAIL.n672 VSUBS 0.021383f
C1625 VTAIL.n673 VSUBS 0.012026f
C1626 VTAIL.n674 VSUBS 1.83116f
C1627 VTAIL.n675 VSUBS 0.02238f
C1628 VTAIL.n676 VSUBS 0.012026f
C1629 VTAIL.n677 VSUBS 0.012734f
C1630 VTAIL.n678 VSUBS 0.028426f
C1631 VTAIL.n679 VSUBS 0.028426f
C1632 VTAIL.n680 VSUBS 0.012734f
C1633 VTAIL.n681 VSUBS 0.012026f
C1634 VTAIL.n682 VSUBS 0.02238f
C1635 VTAIL.n683 VSUBS 0.02238f
C1636 VTAIL.n684 VSUBS 0.012026f
C1637 VTAIL.n685 VSUBS 0.012734f
C1638 VTAIL.n686 VSUBS 0.028426f
C1639 VTAIL.n687 VSUBS 0.028426f
C1640 VTAIL.n688 VSUBS 0.012734f
C1641 VTAIL.n689 VSUBS 0.012026f
C1642 VTAIL.n690 VSUBS 0.02238f
C1643 VTAIL.n691 VSUBS 0.02238f
C1644 VTAIL.n692 VSUBS 0.012026f
C1645 VTAIL.n693 VSUBS 0.01238f
C1646 VTAIL.n694 VSUBS 0.01238f
C1647 VTAIL.n695 VSUBS 0.028426f
C1648 VTAIL.n696 VSUBS 0.028426f
C1649 VTAIL.n697 VSUBS 0.012734f
C1650 VTAIL.n698 VSUBS 0.012026f
C1651 VTAIL.n699 VSUBS 0.02238f
C1652 VTAIL.n700 VSUBS 0.02238f
C1653 VTAIL.n701 VSUBS 0.012026f
C1654 VTAIL.n702 VSUBS 0.012734f
C1655 VTAIL.n703 VSUBS 0.028426f
C1656 VTAIL.n704 VSUBS 0.028426f
C1657 VTAIL.n705 VSUBS 0.012734f
C1658 VTAIL.n706 VSUBS 0.012026f
C1659 VTAIL.n707 VSUBS 0.02238f
C1660 VTAIL.n708 VSUBS 0.02238f
C1661 VTAIL.n709 VSUBS 0.012026f
C1662 VTAIL.n710 VSUBS 0.012734f
C1663 VTAIL.n711 VSUBS 0.028426f
C1664 VTAIL.n712 VSUBS 0.028426f
C1665 VTAIL.n713 VSUBS 0.012734f
C1666 VTAIL.n714 VSUBS 0.012026f
C1667 VTAIL.n715 VSUBS 0.02238f
C1668 VTAIL.n716 VSUBS 0.02238f
C1669 VTAIL.n717 VSUBS 0.012026f
C1670 VTAIL.n718 VSUBS 0.012734f
C1671 VTAIL.n719 VSUBS 0.028426f
C1672 VTAIL.n720 VSUBS 0.028426f
C1673 VTAIL.n721 VSUBS 0.012734f
C1674 VTAIL.n722 VSUBS 0.012026f
C1675 VTAIL.n723 VSUBS 0.02238f
C1676 VTAIL.n724 VSUBS 0.02238f
C1677 VTAIL.n725 VSUBS 0.012026f
C1678 VTAIL.n726 VSUBS 0.012734f
C1679 VTAIL.n727 VSUBS 0.028426f
C1680 VTAIL.n728 VSUBS 0.028426f
C1681 VTAIL.n729 VSUBS 0.012734f
C1682 VTAIL.n730 VSUBS 0.012026f
C1683 VTAIL.n731 VSUBS 0.02238f
C1684 VTAIL.n732 VSUBS 0.02238f
C1685 VTAIL.n733 VSUBS 0.012026f
C1686 VTAIL.n734 VSUBS 0.012734f
C1687 VTAIL.n735 VSUBS 0.028426f
C1688 VTAIL.n736 VSUBS 0.070357f
C1689 VTAIL.n737 VSUBS 0.012734f
C1690 VTAIL.n738 VSUBS 0.023617f
C1691 VTAIL.n739 VSUBS 0.056011f
C1692 VTAIL.n740 VSUBS 0.053757f
C1693 VTAIL.n741 VSUBS 2.00034f
C1694 VTAIL.n742 VSUBS 0.023972f
C1695 VTAIL.n743 VSUBS 0.02238f
C1696 VTAIL.n744 VSUBS 0.012026f
C1697 VTAIL.n745 VSUBS 0.028426f
C1698 VTAIL.n746 VSUBS 0.012734f
C1699 VTAIL.n747 VSUBS 0.02238f
C1700 VTAIL.n748 VSUBS 0.012026f
C1701 VTAIL.n749 VSUBS 0.028426f
C1702 VTAIL.n750 VSUBS 0.012734f
C1703 VTAIL.n751 VSUBS 0.02238f
C1704 VTAIL.n752 VSUBS 0.012026f
C1705 VTAIL.n753 VSUBS 0.028426f
C1706 VTAIL.n754 VSUBS 0.012734f
C1707 VTAIL.n755 VSUBS 0.02238f
C1708 VTAIL.n756 VSUBS 0.012026f
C1709 VTAIL.n757 VSUBS 0.028426f
C1710 VTAIL.n758 VSUBS 0.012734f
C1711 VTAIL.n759 VSUBS 0.02238f
C1712 VTAIL.n760 VSUBS 0.012026f
C1713 VTAIL.n761 VSUBS 0.028426f
C1714 VTAIL.n762 VSUBS 0.012734f
C1715 VTAIL.n763 VSUBS 0.02238f
C1716 VTAIL.n764 VSUBS 0.012026f
C1717 VTAIL.n765 VSUBS 0.028426f
C1718 VTAIL.n766 VSUBS 0.012734f
C1719 VTAIL.n767 VSUBS 0.02238f
C1720 VTAIL.n768 VSUBS 0.012026f
C1721 VTAIL.n769 VSUBS 0.028426f
C1722 VTAIL.n770 VSUBS 0.012734f
C1723 VTAIL.n771 VSUBS 0.02238f
C1724 VTAIL.n772 VSUBS 0.012026f
C1725 VTAIL.n773 VSUBS 0.028426f
C1726 VTAIL.n774 VSUBS 0.012734f
C1727 VTAIL.n775 VSUBS 0.251749f
C1728 VTAIL.t2 VSUBS 0.061818f
C1729 VTAIL.n776 VSUBS 0.021319f
C1730 VTAIL.n777 VSUBS 0.021383f
C1731 VTAIL.n778 VSUBS 0.012026f
C1732 VTAIL.n779 VSUBS 1.83116f
C1733 VTAIL.n780 VSUBS 0.02238f
C1734 VTAIL.n781 VSUBS 0.012026f
C1735 VTAIL.n782 VSUBS 0.012734f
C1736 VTAIL.n783 VSUBS 0.028426f
C1737 VTAIL.n784 VSUBS 0.028426f
C1738 VTAIL.n785 VSUBS 0.012734f
C1739 VTAIL.n786 VSUBS 0.012026f
C1740 VTAIL.n787 VSUBS 0.02238f
C1741 VTAIL.n788 VSUBS 0.02238f
C1742 VTAIL.n789 VSUBS 0.012026f
C1743 VTAIL.n790 VSUBS 0.012734f
C1744 VTAIL.n791 VSUBS 0.028426f
C1745 VTAIL.n792 VSUBS 0.028426f
C1746 VTAIL.n793 VSUBS 0.028426f
C1747 VTAIL.n794 VSUBS 0.012734f
C1748 VTAIL.n795 VSUBS 0.012026f
C1749 VTAIL.n796 VSUBS 0.02238f
C1750 VTAIL.n797 VSUBS 0.02238f
C1751 VTAIL.n798 VSUBS 0.012026f
C1752 VTAIL.n799 VSUBS 0.01238f
C1753 VTAIL.n800 VSUBS 0.01238f
C1754 VTAIL.n801 VSUBS 0.028426f
C1755 VTAIL.n802 VSUBS 0.028426f
C1756 VTAIL.n803 VSUBS 0.012734f
C1757 VTAIL.n804 VSUBS 0.012026f
C1758 VTAIL.n805 VSUBS 0.02238f
C1759 VTAIL.n806 VSUBS 0.02238f
C1760 VTAIL.n807 VSUBS 0.012026f
C1761 VTAIL.n808 VSUBS 0.012734f
C1762 VTAIL.n809 VSUBS 0.028426f
C1763 VTAIL.n810 VSUBS 0.028426f
C1764 VTAIL.n811 VSUBS 0.012734f
C1765 VTAIL.n812 VSUBS 0.012026f
C1766 VTAIL.n813 VSUBS 0.02238f
C1767 VTAIL.n814 VSUBS 0.02238f
C1768 VTAIL.n815 VSUBS 0.012026f
C1769 VTAIL.n816 VSUBS 0.012734f
C1770 VTAIL.n817 VSUBS 0.028426f
C1771 VTAIL.n818 VSUBS 0.028426f
C1772 VTAIL.n819 VSUBS 0.012734f
C1773 VTAIL.n820 VSUBS 0.012026f
C1774 VTAIL.n821 VSUBS 0.02238f
C1775 VTAIL.n822 VSUBS 0.02238f
C1776 VTAIL.n823 VSUBS 0.012026f
C1777 VTAIL.n824 VSUBS 0.012734f
C1778 VTAIL.n825 VSUBS 0.028426f
C1779 VTAIL.n826 VSUBS 0.028426f
C1780 VTAIL.n827 VSUBS 0.012734f
C1781 VTAIL.n828 VSUBS 0.012026f
C1782 VTAIL.n829 VSUBS 0.02238f
C1783 VTAIL.n830 VSUBS 0.02238f
C1784 VTAIL.n831 VSUBS 0.012026f
C1785 VTAIL.n832 VSUBS 0.012734f
C1786 VTAIL.n833 VSUBS 0.028426f
C1787 VTAIL.n834 VSUBS 0.028426f
C1788 VTAIL.n835 VSUBS 0.012734f
C1789 VTAIL.n836 VSUBS 0.012026f
C1790 VTAIL.n837 VSUBS 0.02238f
C1791 VTAIL.n838 VSUBS 0.02238f
C1792 VTAIL.n839 VSUBS 0.012026f
C1793 VTAIL.n840 VSUBS 0.012734f
C1794 VTAIL.n841 VSUBS 0.028426f
C1795 VTAIL.n842 VSUBS 0.070357f
C1796 VTAIL.n843 VSUBS 0.012734f
C1797 VTAIL.n844 VSUBS 0.023617f
C1798 VTAIL.n845 VSUBS 0.056011f
C1799 VTAIL.n846 VSUBS 0.053757f
C1800 VTAIL.n847 VSUBS 1.87989f
C1801 VDD1.t2 VSUBS 0.410863f
C1802 VDD1.t0 VSUBS 0.410863f
C1803 VDD1.n0 VSUBS 3.46634f
C1804 VDD1.t3 VSUBS 0.410863f
C1805 VDD1.t1 VSUBS 0.410863f
C1806 VDD1.n1 VSUBS 4.54074f
C1807 VP.t1 VSUBS 4.957f
C1808 VP.n0 VSUBS 1.80128f
C1809 VP.n1 VSUBS 0.02712f
C1810 VP.n2 VSUBS 0.039423f
C1811 VP.n3 VSUBS 0.02712f
C1812 VP.n4 VSUBS 0.031422f
C1813 VP.t0 VSUBS 5.33626f
C1814 VP.t2 VSUBS 5.32331f
C1815 VP.n5 VSUBS 5.25796f
C1816 VP.t3 VSUBS 4.957f
C1817 VP.n6 VSUBS 1.80128f
C1818 VP.n7 VSUBS 1.84855f
C1819 VP.n8 VSUBS 0.043764f
C1820 VP.n9 VSUBS 0.02712f
C1821 VP.n10 VSUBS 0.050291f
C1822 VP.n11 VSUBS 0.050291f
C1823 VP.n12 VSUBS 0.039423f
C1824 VP.n13 VSUBS 0.02712f
C1825 VP.n14 VSUBS 0.02712f
C1826 VP.n15 VSUBS 0.02712f
C1827 VP.n16 VSUBS 0.050291f
C1828 VP.n17 VSUBS 0.050291f
C1829 VP.n18 VSUBS 0.031422f
C1830 VP.n19 VSUBS 0.043764f
C1831 VP.n20 VSUBS 0.075127f
.ends

