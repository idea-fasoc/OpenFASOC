* NGSPICE file created from diff_pair_sample_1374.ext - technology: sky130A

.subckt diff_pair_sample_1374 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=2.07
X1 B.t8 B.t6 B.t7 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=2.07
X2 B.t5 B.t3 B.t4 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=2.07
X3 VDD2.t3 VN.t0 VTAIL.t7 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=2.07
X4 VTAIL.t4 VN.t1 VDD2.t2 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=2.07
X5 VDD2.t1 VN.t2 VTAIL.t6 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=2.07
X6 VTAIL.t5 VN.t3 VDD2.t0 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=2.07
X7 VDD1.t3 VP.t0 VTAIL.t3 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=2.07
X8 VTAIL.t0 VP.t1 VDD1.t2 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=2.07
X9 B.t2 B.t0 B.t1 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=2.07
X10 VDD1.t1 VP.t2 VTAIL.t1 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=2.07
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n2410_n4968# sky130_fd_pr__pfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=2.07
R0 B.n552 B.n551 585
R1 B.n553 B.n90 585
R2 B.n555 B.n554 585
R3 B.n556 B.n89 585
R4 B.n558 B.n557 585
R5 B.n559 B.n88 585
R6 B.n561 B.n560 585
R7 B.n562 B.n87 585
R8 B.n564 B.n563 585
R9 B.n565 B.n86 585
R10 B.n567 B.n566 585
R11 B.n568 B.n85 585
R12 B.n570 B.n569 585
R13 B.n571 B.n84 585
R14 B.n573 B.n572 585
R15 B.n574 B.n83 585
R16 B.n576 B.n575 585
R17 B.n577 B.n82 585
R18 B.n579 B.n578 585
R19 B.n580 B.n81 585
R20 B.n582 B.n581 585
R21 B.n583 B.n80 585
R22 B.n585 B.n584 585
R23 B.n586 B.n79 585
R24 B.n588 B.n587 585
R25 B.n589 B.n78 585
R26 B.n591 B.n590 585
R27 B.n592 B.n77 585
R28 B.n594 B.n593 585
R29 B.n595 B.n76 585
R30 B.n597 B.n596 585
R31 B.n598 B.n75 585
R32 B.n600 B.n599 585
R33 B.n601 B.n74 585
R34 B.n603 B.n602 585
R35 B.n604 B.n73 585
R36 B.n606 B.n605 585
R37 B.n607 B.n72 585
R38 B.n609 B.n608 585
R39 B.n610 B.n71 585
R40 B.n612 B.n611 585
R41 B.n613 B.n70 585
R42 B.n615 B.n614 585
R43 B.n616 B.n69 585
R44 B.n618 B.n617 585
R45 B.n619 B.n68 585
R46 B.n621 B.n620 585
R47 B.n622 B.n67 585
R48 B.n624 B.n623 585
R49 B.n625 B.n66 585
R50 B.n627 B.n626 585
R51 B.n628 B.n65 585
R52 B.n630 B.n629 585
R53 B.n631 B.n64 585
R54 B.n633 B.n632 585
R55 B.n634 B.n63 585
R56 B.n636 B.n635 585
R57 B.n637 B.n62 585
R58 B.n639 B.n638 585
R59 B.n640 B.n61 585
R60 B.n642 B.n641 585
R61 B.n643 B.n60 585
R62 B.n645 B.n644 585
R63 B.n646 B.n59 585
R64 B.n648 B.n647 585
R65 B.n650 B.n649 585
R66 B.n651 B.n55 585
R67 B.n653 B.n652 585
R68 B.n654 B.n54 585
R69 B.n656 B.n655 585
R70 B.n657 B.n53 585
R71 B.n659 B.n658 585
R72 B.n660 B.n52 585
R73 B.n662 B.n661 585
R74 B.n663 B.n49 585
R75 B.n666 B.n665 585
R76 B.n667 B.n48 585
R77 B.n669 B.n668 585
R78 B.n670 B.n47 585
R79 B.n672 B.n671 585
R80 B.n673 B.n46 585
R81 B.n675 B.n674 585
R82 B.n676 B.n45 585
R83 B.n678 B.n677 585
R84 B.n679 B.n44 585
R85 B.n681 B.n680 585
R86 B.n682 B.n43 585
R87 B.n684 B.n683 585
R88 B.n685 B.n42 585
R89 B.n687 B.n686 585
R90 B.n688 B.n41 585
R91 B.n690 B.n689 585
R92 B.n691 B.n40 585
R93 B.n693 B.n692 585
R94 B.n694 B.n39 585
R95 B.n696 B.n695 585
R96 B.n697 B.n38 585
R97 B.n699 B.n698 585
R98 B.n700 B.n37 585
R99 B.n702 B.n701 585
R100 B.n703 B.n36 585
R101 B.n705 B.n704 585
R102 B.n706 B.n35 585
R103 B.n708 B.n707 585
R104 B.n709 B.n34 585
R105 B.n711 B.n710 585
R106 B.n712 B.n33 585
R107 B.n714 B.n713 585
R108 B.n715 B.n32 585
R109 B.n717 B.n716 585
R110 B.n718 B.n31 585
R111 B.n720 B.n719 585
R112 B.n721 B.n30 585
R113 B.n723 B.n722 585
R114 B.n724 B.n29 585
R115 B.n726 B.n725 585
R116 B.n727 B.n28 585
R117 B.n729 B.n728 585
R118 B.n730 B.n27 585
R119 B.n732 B.n731 585
R120 B.n733 B.n26 585
R121 B.n735 B.n734 585
R122 B.n736 B.n25 585
R123 B.n738 B.n737 585
R124 B.n739 B.n24 585
R125 B.n741 B.n740 585
R126 B.n742 B.n23 585
R127 B.n744 B.n743 585
R128 B.n745 B.n22 585
R129 B.n747 B.n746 585
R130 B.n748 B.n21 585
R131 B.n750 B.n749 585
R132 B.n751 B.n20 585
R133 B.n753 B.n752 585
R134 B.n754 B.n19 585
R135 B.n756 B.n755 585
R136 B.n757 B.n18 585
R137 B.n759 B.n758 585
R138 B.n760 B.n17 585
R139 B.n762 B.n761 585
R140 B.n550 B.n91 585
R141 B.n549 B.n548 585
R142 B.n547 B.n92 585
R143 B.n546 B.n545 585
R144 B.n544 B.n93 585
R145 B.n543 B.n542 585
R146 B.n541 B.n94 585
R147 B.n540 B.n539 585
R148 B.n538 B.n95 585
R149 B.n537 B.n536 585
R150 B.n535 B.n96 585
R151 B.n534 B.n533 585
R152 B.n532 B.n97 585
R153 B.n531 B.n530 585
R154 B.n529 B.n98 585
R155 B.n528 B.n527 585
R156 B.n526 B.n99 585
R157 B.n525 B.n524 585
R158 B.n523 B.n100 585
R159 B.n522 B.n521 585
R160 B.n520 B.n101 585
R161 B.n519 B.n518 585
R162 B.n517 B.n102 585
R163 B.n516 B.n515 585
R164 B.n514 B.n103 585
R165 B.n513 B.n512 585
R166 B.n511 B.n104 585
R167 B.n510 B.n509 585
R168 B.n508 B.n105 585
R169 B.n507 B.n506 585
R170 B.n505 B.n106 585
R171 B.n504 B.n503 585
R172 B.n502 B.n107 585
R173 B.n501 B.n500 585
R174 B.n499 B.n108 585
R175 B.n498 B.n497 585
R176 B.n496 B.n109 585
R177 B.n495 B.n494 585
R178 B.n493 B.n110 585
R179 B.n492 B.n491 585
R180 B.n490 B.n111 585
R181 B.n489 B.n488 585
R182 B.n487 B.n112 585
R183 B.n486 B.n485 585
R184 B.n484 B.n113 585
R185 B.n483 B.n482 585
R186 B.n481 B.n114 585
R187 B.n480 B.n479 585
R188 B.n478 B.n115 585
R189 B.n477 B.n476 585
R190 B.n475 B.n116 585
R191 B.n474 B.n473 585
R192 B.n472 B.n117 585
R193 B.n471 B.n470 585
R194 B.n469 B.n118 585
R195 B.n468 B.n467 585
R196 B.n466 B.n119 585
R197 B.n465 B.n464 585
R198 B.n463 B.n120 585
R199 B.n252 B.n251 585
R200 B.n253 B.n194 585
R201 B.n255 B.n254 585
R202 B.n256 B.n193 585
R203 B.n258 B.n257 585
R204 B.n259 B.n192 585
R205 B.n261 B.n260 585
R206 B.n262 B.n191 585
R207 B.n264 B.n263 585
R208 B.n265 B.n190 585
R209 B.n267 B.n266 585
R210 B.n268 B.n189 585
R211 B.n270 B.n269 585
R212 B.n271 B.n188 585
R213 B.n273 B.n272 585
R214 B.n274 B.n187 585
R215 B.n276 B.n275 585
R216 B.n277 B.n186 585
R217 B.n279 B.n278 585
R218 B.n280 B.n185 585
R219 B.n282 B.n281 585
R220 B.n283 B.n184 585
R221 B.n285 B.n284 585
R222 B.n286 B.n183 585
R223 B.n288 B.n287 585
R224 B.n289 B.n182 585
R225 B.n291 B.n290 585
R226 B.n292 B.n181 585
R227 B.n294 B.n293 585
R228 B.n295 B.n180 585
R229 B.n297 B.n296 585
R230 B.n298 B.n179 585
R231 B.n300 B.n299 585
R232 B.n301 B.n178 585
R233 B.n303 B.n302 585
R234 B.n304 B.n177 585
R235 B.n306 B.n305 585
R236 B.n307 B.n176 585
R237 B.n309 B.n308 585
R238 B.n310 B.n175 585
R239 B.n312 B.n311 585
R240 B.n313 B.n174 585
R241 B.n315 B.n314 585
R242 B.n316 B.n173 585
R243 B.n318 B.n317 585
R244 B.n319 B.n172 585
R245 B.n321 B.n320 585
R246 B.n322 B.n171 585
R247 B.n324 B.n323 585
R248 B.n325 B.n170 585
R249 B.n327 B.n326 585
R250 B.n328 B.n169 585
R251 B.n330 B.n329 585
R252 B.n331 B.n168 585
R253 B.n333 B.n332 585
R254 B.n334 B.n167 585
R255 B.n336 B.n335 585
R256 B.n337 B.n166 585
R257 B.n339 B.n338 585
R258 B.n340 B.n165 585
R259 B.n342 B.n341 585
R260 B.n343 B.n164 585
R261 B.n345 B.n344 585
R262 B.n346 B.n163 585
R263 B.n348 B.n347 585
R264 B.n350 B.n349 585
R265 B.n351 B.n159 585
R266 B.n353 B.n352 585
R267 B.n354 B.n158 585
R268 B.n356 B.n355 585
R269 B.n357 B.n157 585
R270 B.n359 B.n358 585
R271 B.n360 B.n156 585
R272 B.n362 B.n361 585
R273 B.n363 B.n153 585
R274 B.n366 B.n365 585
R275 B.n367 B.n152 585
R276 B.n369 B.n368 585
R277 B.n370 B.n151 585
R278 B.n372 B.n371 585
R279 B.n373 B.n150 585
R280 B.n375 B.n374 585
R281 B.n376 B.n149 585
R282 B.n378 B.n377 585
R283 B.n379 B.n148 585
R284 B.n381 B.n380 585
R285 B.n382 B.n147 585
R286 B.n384 B.n383 585
R287 B.n385 B.n146 585
R288 B.n387 B.n386 585
R289 B.n388 B.n145 585
R290 B.n390 B.n389 585
R291 B.n391 B.n144 585
R292 B.n393 B.n392 585
R293 B.n394 B.n143 585
R294 B.n396 B.n395 585
R295 B.n397 B.n142 585
R296 B.n399 B.n398 585
R297 B.n400 B.n141 585
R298 B.n402 B.n401 585
R299 B.n403 B.n140 585
R300 B.n405 B.n404 585
R301 B.n406 B.n139 585
R302 B.n408 B.n407 585
R303 B.n409 B.n138 585
R304 B.n411 B.n410 585
R305 B.n412 B.n137 585
R306 B.n414 B.n413 585
R307 B.n415 B.n136 585
R308 B.n417 B.n416 585
R309 B.n418 B.n135 585
R310 B.n420 B.n419 585
R311 B.n421 B.n134 585
R312 B.n423 B.n422 585
R313 B.n424 B.n133 585
R314 B.n426 B.n425 585
R315 B.n427 B.n132 585
R316 B.n429 B.n428 585
R317 B.n430 B.n131 585
R318 B.n432 B.n431 585
R319 B.n433 B.n130 585
R320 B.n435 B.n434 585
R321 B.n436 B.n129 585
R322 B.n438 B.n437 585
R323 B.n439 B.n128 585
R324 B.n441 B.n440 585
R325 B.n442 B.n127 585
R326 B.n444 B.n443 585
R327 B.n445 B.n126 585
R328 B.n447 B.n446 585
R329 B.n448 B.n125 585
R330 B.n450 B.n449 585
R331 B.n451 B.n124 585
R332 B.n453 B.n452 585
R333 B.n454 B.n123 585
R334 B.n456 B.n455 585
R335 B.n457 B.n122 585
R336 B.n459 B.n458 585
R337 B.n460 B.n121 585
R338 B.n462 B.n461 585
R339 B.n250 B.n195 585
R340 B.n249 B.n248 585
R341 B.n247 B.n196 585
R342 B.n246 B.n245 585
R343 B.n244 B.n197 585
R344 B.n243 B.n242 585
R345 B.n241 B.n198 585
R346 B.n240 B.n239 585
R347 B.n238 B.n199 585
R348 B.n237 B.n236 585
R349 B.n235 B.n200 585
R350 B.n234 B.n233 585
R351 B.n232 B.n201 585
R352 B.n231 B.n230 585
R353 B.n229 B.n202 585
R354 B.n228 B.n227 585
R355 B.n226 B.n203 585
R356 B.n225 B.n224 585
R357 B.n223 B.n204 585
R358 B.n222 B.n221 585
R359 B.n220 B.n205 585
R360 B.n219 B.n218 585
R361 B.n217 B.n206 585
R362 B.n216 B.n215 585
R363 B.n214 B.n207 585
R364 B.n213 B.n212 585
R365 B.n211 B.n208 585
R366 B.n210 B.n209 585
R367 B.n2 B.n0 585
R368 B.n805 B.n1 585
R369 B.n804 B.n803 585
R370 B.n802 B.n3 585
R371 B.n801 B.n800 585
R372 B.n799 B.n4 585
R373 B.n798 B.n797 585
R374 B.n796 B.n5 585
R375 B.n795 B.n794 585
R376 B.n793 B.n6 585
R377 B.n792 B.n791 585
R378 B.n790 B.n7 585
R379 B.n789 B.n788 585
R380 B.n787 B.n8 585
R381 B.n786 B.n785 585
R382 B.n784 B.n9 585
R383 B.n783 B.n782 585
R384 B.n781 B.n10 585
R385 B.n780 B.n779 585
R386 B.n778 B.n11 585
R387 B.n777 B.n776 585
R388 B.n775 B.n12 585
R389 B.n774 B.n773 585
R390 B.n772 B.n13 585
R391 B.n771 B.n770 585
R392 B.n769 B.n14 585
R393 B.n768 B.n767 585
R394 B.n766 B.n15 585
R395 B.n765 B.n764 585
R396 B.n763 B.n16 585
R397 B.n807 B.n806 585
R398 B.n252 B.n195 535.745
R399 B.n763 B.n762 535.745
R400 B.n463 B.n462 535.745
R401 B.n552 B.n91 535.745
R402 B.n154 B.t0 439.928
R403 B.n160 B.t6 439.928
R404 B.n50 B.t9 439.928
R405 B.n56 B.t3 439.928
R406 B.n248 B.n195 163.367
R407 B.n248 B.n247 163.367
R408 B.n247 B.n246 163.367
R409 B.n246 B.n197 163.367
R410 B.n242 B.n197 163.367
R411 B.n242 B.n241 163.367
R412 B.n241 B.n240 163.367
R413 B.n240 B.n199 163.367
R414 B.n236 B.n199 163.367
R415 B.n236 B.n235 163.367
R416 B.n235 B.n234 163.367
R417 B.n234 B.n201 163.367
R418 B.n230 B.n201 163.367
R419 B.n230 B.n229 163.367
R420 B.n229 B.n228 163.367
R421 B.n228 B.n203 163.367
R422 B.n224 B.n203 163.367
R423 B.n224 B.n223 163.367
R424 B.n223 B.n222 163.367
R425 B.n222 B.n205 163.367
R426 B.n218 B.n205 163.367
R427 B.n218 B.n217 163.367
R428 B.n217 B.n216 163.367
R429 B.n216 B.n207 163.367
R430 B.n212 B.n207 163.367
R431 B.n212 B.n211 163.367
R432 B.n211 B.n210 163.367
R433 B.n210 B.n2 163.367
R434 B.n806 B.n2 163.367
R435 B.n806 B.n805 163.367
R436 B.n805 B.n804 163.367
R437 B.n804 B.n3 163.367
R438 B.n800 B.n3 163.367
R439 B.n800 B.n799 163.367
R440 B.n799 B.n798 163.367
R441 B.n798 B.n5 163.367
R442 B.n794 B.n5 163.367
R443 B.n794 B.n793 163.367
R444 B.n793 B.n792 163.367
R445 B.n792 B.n7 163.367
R446 B.n788 B.n7 163.367
R447 B.n788 B.n787 163.367
R448 B.n787 B.n786 163.367
R449 B.n786 B.n9 163.367
R450 B.n782 B.n9 163.367
R451 B.n782 B.n781 163.367
R452 B.n781 B.n780 163.367
R453 B.n780 B.n11 163.367
R454 B.n776 B.n11 163.367
R455 B.n776 B.n775 163.367
R456 B.n775 B.n774 163.367
R457 B.n774 B.n13 163.367
R458 B.n770 B.n13 163.367
R459 B.n770 B.n769 163.367
R460 B.n769 B.n768 163.367
R461 B.n768 B.n15 163.367
R462 B.n764 B.n15 163.367
R463 B.n764 B.n763 163.367
R464 B.n253 B.n252 163.367
R465 B.n254 B.n253 163.367
R466 B.n254 B.n193 163.367
R467 B.n258 B.n193 163.367
R468 B.n259 B.n258 163.367
R469 B.n260 B.n259 163.367
R470 B.n260 B.n191 163.367
R471 B.n264 B.n191 163.367
R472 B.n265 B.n264 163.367
R473 B.n266 B.n265 163.367
R474 B.n266 B.n189 163.367
R475 B.n270 B.n189 163.367
R476 B.n271 B.n270 163.367
R477 B.n272 B.n271 163.367
R478 B.n272 B.n187 163.367
R479 B.n276 B.n187 163.367
R480 B.n277 B.n276 163.367
R481 B.n278 B.n277 163.367
R482 B.n278 B.n185 163.367
R483 B.n282 B.n185 163.367
R484 B.n283 B.n282 163.367
R485 B.n284 B.n283 163.367
R486 B.n284 B.n183 163.367
R487 B.n288 B.n183 163.367
R488 B.n289 B.n288 163.367
R489 B.n290 B.n289 163.367
R490 B.n290 B.n181 163.367
R491 B.n294 B.n181 163.367
R492 B.n295 B.n294 163.367
R493 B.n296 B.n295 163.367
R494 B.n296 B.n179 163.367
R495 B.n300 B.n179 163.367
R496 B.n301 B.n300 163.367
R497 B.n302 B.n301 163.367
R498 B.n302 B.n177 163.367
R499 B.n306 B.n177 163.367
R500 B.n307 B.n306 163.367
R501 B.n308 B.n307 163.367
R502 B.n308 B.n175 163.367
R503 B.n312 B.n175 163.367
R504 B.n313 B.n312 163.367
R505 B.n314 B.n313 163.367
R506 B.n314 B.n173 163.367
R507 B.n318 B.n173 163.367
R508 B.n319 B.n318 163.367
R509 B.n320 B.n319 163.367
R510 B.n320 B.n171 163.367
R511 B.n324 B.n171 163.367
R512 B.n325 B.n324 163.367
R513 B.n326 B.n325 163.367
R514 B.n326 B.n169 163.367
R515 B.n330 B.n169 163.367
R516 B.n331 B.n330 163.367
R517 B.n332 B.n331 163.367
R518 B.n332 B.n167 163.367
R519 B.n336 B.n167 163.367
R520 B.n337 B.n336 163.367
R521 B.n338 B.n337 163.367
R522 B.n338 B.n165 163.367
R523 B.n342 B.n165 163.367
R524 B.n343 B.n342 163.367
R525 B.n344 B.n343 163.367
R526 B.n344 B.n163 163.367
R527 B.n348 B.n163 163.367
R528 B.n349 B.n348 163.367
R529 B.n349 B.n159 163.367
R530 B.n353 B.n159 163.367
R531 B.n354 B.n353 163.367
R532 B.n355 B.n354 163.367
R533 B.n355 B.n157 163.367
R534 B.n359 B.n157 163.367
R535 B.n360 B.n359 163.367
R536 B.n361 B.n360 163.367
R537 B.n361 B.n153 163.367
R538 B.n366 B.n153 163.367
R539 B.n367 B.n366 163.367
R540 B.n368 B.n367 163.367
R541 B.n368 B.n151 163.367
R542 B.n372 B.n151 163.367
R543 B.n373 B.n372 163.367
R544 B.n374 B.n373 163.367
R545 B.n374 B.n149 163.367
R546 B.n378 B.n149 163.367
R547 B.n379 B.n378 163.367
R548 B.n380 B.n379 163.367
R549 B.n380 B.n147 163.367
R550 B.n384 B.n147 163.367
R551 B.n385 B.n384 163.367
R552 B.n386 B.n385 163.367
R553 B.n386 B.n145 163.367
R554 B.n390 B.n145 163.367
R555 B.n391 B.n390 163.367
R556 B.n392 B.n391 163.367
R557 B.n392 B.n143 163.367
R558 B.n396 B.n143 163.367
R559 B.n397 B.n396 163.367
R560 B.n398 B.n397 163.367
R561 B.n398 B.n141 163.367
R562 B.n402 B.n141 163.367
R563 B.n403 B.n402 163.367
R564 B.n404 B.n403 163.367
R565 B.n404 B.n139 163.367
R566 B.n408 B.n139 163.367
R567 B.n409 B.n408 163.367
R568 B.n410 B.n409 163.367
R569 B.n410 B.n137 163.367
R570 B.n414 B.n137 163.367
R571 B.n415 B.n414 163.367
R572 B.n416 B.n415 163.367
R573 B.n416 B.n135 163.367
R574 B.n420 B.n135 163.367
R575 B.n421 B.n420 163.367
R576 B.n422 B.n421 163.367
R577 B.n422 B.n133 163.367
R578 B.n426 B.n133 163.367
R579 B.n427 B.n426 163.367
R580 B.n428 B.n427 163.367
R581 B.n428 B.n131 163.367
R582 B.n432 B.n131 163.367
R583 B.n433 B.n432 163.367
R584 B.n434 B.n433 163.367
R585 B.n434 B.n129 163.367
R586 B.n438 B.n129 163.367
R587 B.n439 B.n438 163.367
R588 B.n440 B.n439 163.367
R589 B.n440 B.n127 163.367
R590 B.n444 B.n127 163.367
R591 B.n445 B.n444 163.367
R592 B.n446 B.n445 163.367
R593 B.n446 B.n125 163.367
R594 B.n450 B.n125 163.367
R595 B.n451 B.n450 163.367
R596 B.n452 B.n451 163.367
R597 B.n452 B.n123 163.367
R598 B.n456 B.n123 163.367
R599 B.n457 B.n456 163.367
R600 B.n458 B.n457 163.367
R601 B.n458 B.n121 163.367
R602 B.n462 B.n121 163.367
R603 B.n464 B.n463 163.367
R604 B.n464 B.n119 163.367
R605 B.n468 B.n119 163.367
R606 B.n469 B.n468 163.367
R607 B.n470 B.n469 163.367
R608 B.n470 B.n117 163.367
R609 B.n474 B.n117 163.367
R610 B.n475 B.n474 163.367
R611 B.n476 B.n475 163.367
R612 B.n476 B.n115 163.367
R613 B.n480 B.n115 163.367
R614 B.n481 B.n480 163.367
R615 B.n482 B.n481 163.367
R616 B.n482 B.n113 163.367
R617 B.n486 B.n113 163.367
R618 B.n487 B.n486 163.367
R619 B.n488 B.n487 163.367
R620 B.n488 B.n111 163.367
R621 B.n492 B.n111 163.367
R622 B.n493 B.n492 163.367
R623 B.n494 B.n493 163.367
R624 B.n494 B.n109 163.367
R625 B.n498 B.n109 163.367
R626 B.n499 B.n498 163.367
R627 B.n500 B.n499 163.367
R628 B.n500 B.n107 163.367
R629 B.n504 B.n107 163.367
R630 B.n505 B.n504 163.367
R631 B.n506 B.n505 163.367
R632 B.n506 B.n105 163.367
R633 B.n510 B.n105 163.367
R634 B.n511 B.n510 163.367
R635 B.n512 B.n511 163.367
R636 B.n512 B.n103 163.367
R637 B.n516 B.n103 163.367
R638 B.n517 B.n516 163.367
R639 B.n518 B.n517 163.367
R640 B.n518 B.n101 163.367
R641 B.n522 B.n101 163.367
R642 B.n523 B.n522 163.367
R643 B.n524 B.n523 163.367
R644 B.n524 B.n99 163.367
R645 B.n528 B.n99 163.367
R646 B.n529 B.n528 163.367
R647 B.n530 B.n529 163.367
R648 B.n530 B.n97 163.367
R649 B.n534 B.n97 163.367
R650 B.n535 B.n534 163.367
R651 B.n536 B.n535 163.367
R652 B.n536 B.n95 163.367
R653 B.n540 B.n95 163.367
R654 B.n541 B.n540 163.367
R655 B.n542 B.n541 163.367
R656 B.n542 B.n93 163.367
R657 B.n546 B.n93 163.367
R658 B.n547 B.n546 163.367
R659 B.n548 B.n547 163.367
R660 B.n548 B.n91 163.367
R661 B.n762 B.n17 163.367
R662 B.n758 B.n17 163.367
R663 B.n758 B.n757 163.367
R664 B.n757 B.n756 163.367
R665 B.n756 B.n19 163.367
R666 B.n752 B.n19 163.367
R667 B.n752 B.n751 163.367
R668 B.n751 B.n750 163.367
R669 B.n750 B.n21 163.367
R670 B.n746 B.n21 163.367
R671 B.n746 B.n745 163.367
R672 B.n745 B.n744 163.367
R673 B.n744 B.n23 163.367
R674 B.n740 B.n23 163.367
R675 B.n740 B.n739 163.367
R676 B.n739 B.n738 163.367
R677 B.n738 B.n25 163.367
R678 B.n734 B.n25 163.367
R679 B.n734 B.n733 163.367
R680 B.n733 B.n732 163.367
R681 B.n732 B.n27 163.367
R682 B.n728 B.n27 163.367
R683 B.n728 B.n727 163.367
R684 B.n727 B.n726 163.367
R685 B.n726 B.n29 163.367
R686 B.n722 B.n29 163.367
R687 B.n722 B.n721 163.367
R688 B.n721 B.n720 163.367
R689 B.n720 B.n31 163.367
R690 B.n716 B.n31 163.367
R691 B.n716 B.n715 163.367
R692 B.n715 B.n714 163.367
R693 B.n714 B.n33 163.367
R694 B.n710 B.n33 163.367
R695 B.n710 B.n709 163.367
R696 B.n709 B.n708 163.367
R697 B.n708 B.n35 163.367
R698 B.n704 B.n35 163.367
R699 B.n704 B.n703 163.367
R700 B.n703 B.n702 163.367
R701 B.n702 B.n37 163.367
R702 B.n698 B.n37 163.367
R703 B.n698 B.n697 163.367
R704 B.n697 B.n696 163.367
R705 B.n696 B.n39 163.367
R706 B.n692 B.n39 163.367
R707 B.n692 B.n691 163.367
R708 B.n691 B.n690 163.367
R709 B.n690 B.n41 163.367
R710 B.n686 B.n41 163.367
R711 B.n686 B.n685 163.367
R712 B.n685 B.n684 163.367
R713 B.n684 B.n43 163.367
R714 B.n680 B.n43 163.367
R715 B.n680 B.n679 163.367
R716 B.n679 B.n678 163.367
R717 B.n678 B.n45 163.367
R718 B.n674 B.n45 163.367
R719 B.n674 B.n673 163.367
R720 B.n673 B.n672 163.367
R721 B.n672 B.n47 163.367
R722 B.n668 B.n47 163.367
R723 B.n668 B.n667 163.367
R724 B.n667 B.n666 163.367
R725 B.n666 B.n49 163.367
R726 B.n661 B.n49 163.367
R727 B.n661 B.n660 163.367
R728 B.n660 B.n659 163.367
R729 B.n659 B.n53 163.367
R730 B.n655 B.n53 163.367
R731 B.n655 B.n654 163.367
R732 B.n654 B.n653 163.367
R733 B.n653 B.n55 163.367
R734 B.n649 B.n55 163.367
R735 B.n649 B.n648 163.367
R736 B.n648 B.n59 163.367
R737 B.n644 B.n59 163.367
R738 B.n644 B.n643 163.367
R739 B.n643 B.n642 163.367
R740 B.n642 B.n61 163.367
R741 B.n638 B.n61 163.367
R742 B.n638 B.n637 163.367
R743 B.n637 B.n636 163.367
R744 B.n636 B.n63 163.367
R745 B.n632 B.n63 163.367
R746 B.n632 B.n631 163.367
R747 B.n631 B.n630 163.367
R748 B.n630 B.n65 163.367
R749 B.n626 B.n65 163.367
R750 B.n626 B.n625 163.367
R751 B.n625 B.n624 163.367
R752 B.n624 B.n67 163.367
R753 B.n620 B.n67 163.367
R754 B.n620 B.n619 163.367
R755 B.n619 B.n618 163.367
R756 B.n618 B.n69 163.367
R757 B.n614 B.n69 163.367
R758 B.n614 B.n613 163.367
R759 B.n613 B.n612 163.367
R760 B.n612 B.n71 163.367
R761 B.n608 B.n71 163.367
R762 B.n608 B.n607 163.367
R763 B.n607 B.n606 163.367
R764 B.n606 B.n73 163.367
R765 B.n602 B.n73 163.367
R766 B.n602 B.n601 163.367
R767 B.n601 B.n600 163.367
R768 B.n600 B.n75 163.367
R769 B.n596 B.n75 163.367
R770 B.n596 B.n595 163.367
R771 B.n595 B.n594 163.367
R772 B.n594 B.n77 163.367
R773 B.n590 B.n77 163.367
R774 B.n590 B.n589 163.367
R775 B.n589 B.n588 163.367
R776 B.n588 B.n79 163.367
R777 B.n584 B.n79 163.367
R778 B.n584 B.n583 163.367
R779 B.n583 B.n582 163.367
R780 B.n582 B.n81 163.367
R781 B.n578 B.n81 163.367
R782 B.n578 B.n577 163.367
R783 B.n577 B.n576 163.367
R784 B.n576 B.n83 163.367
R785 B.n572 B.n83 163.367
R786 B.n572 B.n571 163.367
R787 B.n571 B.n570 163.367
R788 B.n570 B.n85 163.367
R789 B.n566 B.n85 163.367
R790 B.n566 B.n565 163.367
R791 B.n565 B.n564 163.367
R792 B.n564 B.n87 163.367
R793 B.n560 B.n87 163.367
R794 B.n560 B.n559 163.367
R795 B.n559 B.n558 163.367
R796 B.n558 B.n89 163.367
R797 B.n554 B.n89 163.367
R798 B.n554 B.n553 163.367
R799 B.n553 B.n552 163.367
R800 B.n154 B.t2 158.001
R801 B.n56 B.t4 158.001
R802 B.n160 B.t8 157.976
R803 B.n50 B.t10 157.976
R804 B.n155 B.t1 111.457
R805 B.n57 B.t5 111.457
R806 B.n161 B.t7 111.43
R807 B.n51 B.t11 111.43
R808 B.n364 B.n155 59.5399
R809 B.n162 B.n161 59.5399
R810 B.n664 B.n51 59.5399
R811 B.n58 B.n57 59.5399
R812 B.n155 B.n154 46.546
R813 B.n161 B.n160 46.546
R814 B.n51 B.n50 46.546
R815 B.n57 B.n56 46.546
R816 B.n761 B.n16 34.8103
R817 B.n551 B.n550 34.8103
R818 B.n461 B.n120 34.8103
R819 B.n251 B.n250 34.8103
R820 B B.n807 18.0485
R821 B.n761 B.n760 10.6151
R822 B.n760 B.n759 10.6151
R823 B.n759 B.n18 10.6151
R824 B.n755 B.n18 10.6151
R825 B.n755 B.n754 10.6151
R826 B.n754 B.n753 10.6151
R827 B.n753 B.n20 10.6151
R828 B.n749 B.n20 10.6151
R829 B.n749 B.n748 10.6151
R830 B.n748 B.n747 10.6151
R831 B.n747 B.n22 10.6151
R832 B.n743 B.n22 10.6151
R833 B.n743 B.n742 10.6151
R834 B.n742 B.n741 10.6151
R835 B.n741 B.n24 10.6151
R836 B.n737 B.n24 10.6151
R837 B.n737 B.n736 10.6151
R838 B.n736 B.n735 10.6151
R839 B.n735 B.n26 10.6151
R840 B.n731 B.n26 10.6151
R841 B.n731 B.n730 10.6151
R842 B.n730 B.n729 10.6151
R843 B.n729 B.n28 10.6151
R844 B.n725 B.n28 10.6151
R845 B.n725 B.n724 10.6151
R846 B.n724 B.n723 10.6151
R847 B.n723 B.n30 10.6151
R848 B.n719 B.n30 10.6151
R849 B.n719 B.n718 10.6151
R850 B.n718 B.n717 10.6151
R851 B.n717 B.n32 10.6151
R852 B.n713 B.n32 10.6151
R853 B.n713 B.n712 10.6151
R854 B.n712 B.n711 10.6151
R855 B.n711 B.n34 10.6151
R856 B.n707 B.n34 10.6151
R857 B.n707 B.n706 10.6151
R858 B.n706 B.n705 10.6151
R859 B.n705 B.n36 10.6151
R860 B.n701 B.n36 10.6151
R861 B.n701 B.n700 10.6151
R862 B.n700 B.n699 10.6151
R863 B.n699 B.n38 10.6151
R864 B.n695 B.n38 10.6151
R865 B.n695 B.n694 10.6151
R866 B.n694 B.n693 10.6151
R867 B.n693 B.n40 10.6151
R868 B.n689 B.n40 10.6151
R869 B.n689 B.n688 10.6151
R870 B.n688 B.n687 10.6151
R871 B.n687 B.n42 10.6151
R872 B.n683 B.n42 10.6151
R873 B.n683 B.n682 10.6151
R874 B.n682 B.n681 10.6151
R875 B.n681 B.n44 10.6151
R876 B.n677 B.n44 10.6151
R877 B.n677 B.n676 10.6151
R878 B.n676 B.n675 10.6151
R879 B.n675 B.n46 10.6151
R880 B.n671 B.n46 10.6151
R881 B.n671 B.n670 10.6151
R882 B.n670 B.n669 10.6151
R883 B.n669 B.n48 10.6151
R884 B.n665 B.n48 10.6151
R885 B.n663 B.n662 10.6151
R886 B.n662 B.n52 10.6151
R887 B.n658 B.n52 10.6151
R888 B.n658 B.n657 10.6151
R889 B.n657 B.n656 10.6151
R890 B.n656 B.n54 10.6151
R891 B.n652 B.n54 10.6151
R892 B.n652 B.n651 10.6151
R893 B.n651 B.n650 10.6151
R894 B.n647 B.n646 10.6151
R895 B.n646 B.n645 10.6151
R896 B.n645 B.n60 10.6151
R897 B.n641 B.n60 10.6151
R898 B.n641 B.n640 10.6151
R899 B.n640 B.n639 10.6151
R900 B.n639 B.n62 10.6151
R901 B.n635 B.n62 10.6151
R902 B.n635 B.n634 10.6151
R903 B.n634 B.n633 10.6151
R904 B.n633 B.n64 10.6151
R905 B.n629 B.n64 10.6151
R906 B.n629 B.n628 10.6151
R907 B.n628 B.n627 10.6151
R908 B.n627 B.n66 10.6151
R909 B.n623 B.n66 10.6151
R910 B.n623 B.n622 10.6151
R911 B.n622 B.n621 10.6151
R912 B.n621 B.n68 10.6151
R913 B.n617 B.n68 10.6151
R914 B.n617 B.n616 10.6151
R915 B.n616 B.n615 10.6151
R916 B.n615 B.n70 10.6151
R917 B.n611 B.n70 10.6151
R918 B.n611 B.n610 10.6151
R919 B.n610 B.n609 10.6151
R920 B.n609 B.n72 10.6151
R921 B.n605 B.n72 10.6151
R922 B.n605 B.n604 10.6151
R923 B.n604 B.n603 10.6151
R924 B.n603 B.n74 10.6151
R925 B.n599 B.n74 10.6151
R926 B.n599 B.n598 10.6151
R927 B.n598 B.n597 10.6151
R928 B.n597 B.n76 10.6151
R929 B.n593 B.n76 10.6151
R930 B.n593 B.n592 10.6151
R931 B.n592 B.n591 10.6151
R932 B.n591 B.n78 10.6151
R933 B.n587 B.n78 10.6151
R934 B.n587 B.n586 10.6151
R935 B.n586 B.n585 10.6151
R936 B.n585 B.n80 10.6151
R937 B.n581 B.n80 10.6151
R938 B.n581 B.n580 10.6151
R939 B.n580 B.n579 10.6151
R940 B.n579 B.n82 10.6151
R941 B.n575 B.n82 10.6151
R942 B.n575 B.n574 10.6151
R943 B.n574 B.n573 10.6151
R944 B.n573 B.n84 10.6151
R945 B.n569 B.n84 10.6151
R946 B.n569 B.n568 10.6151
R947 B.n568 B.n567 10.6151
R948 B.n567 B.n86 10.6151
R949 B.n563 B.n86 10.6151
R950 B.n563 B.n562 10.6151
R951 B.n562 B.n561 10.6151
R952 B.n561 B.n88 10.6151
R953 B.n557 B.n88 10.6151
R954 B.n557 B.n556 10.6151
R955 B.n556 B.n555 10.6151
R956 B.n555 B.n90 10.6151
R957 B.n551 B.n90 10.6151
R958 B.n465 B.n120 10.6151
R959 B.n466 B.n465 10.6151
R960 B.n467 B.n466 10.6151
R961 B.n467 B.n118 10.6151
R962 B.n471 B.n118 10.6151
R963 B.n472 B.n471 10.6151
R964 B.n473 B.n472 10.6151
R965 B.n473 B.n116 10.6151
R966 B.n477 B.n116 10.6151
R967 B.n478 B.n477 10.6151
R968 B.n479 B.n478 10.6151
R969 B.n479 B.n114 10.6151
R970 B.n483 B.n114 10.6151
R971 B.n484 B.n483 10.6151
R972 B.n485 B.n484 10.6151
R973 B.n485 B.n112 10.6151
R974 B.n489 B.n112 10.6151
R975 B.n490 B.n489 10.6151
R976 B.n491 B.n490 10.6151
R977 B.n491 B.n110 10.6151
R978 B.n495 B.n110 10.6151
R979 B.n496 B.n495 10.6151
R980 B.n497 B.n496 10.6151
R981 B.n497 B.n108 10.6151
R982 B.n501 B.n108 10.6151
R983 B.n502 B.n501 10.6151
R984 B.n503 B.n502 10.6151
R985 B.n503 B.n106 10.6151
R986 B.n507 B.n106 10.6151
R987 B.n508 B.n507 10.6151
R988 B.n509 B.n508 10.6151
R989 B.n509 B.n104 10.6151
R990 B.n513 B.n104 10.6151
R991 B.n514 B.n513 10.6151
R992 B.n515 B.n514 10.6151
R993 B.n515 B.n102 10.6151
R994 B.n519 B.n102 10.6151
R995 B.n520 B.n519 10.6151
R996 B.n521 B.n520 10.6151
R997 B.n521 B.n100 10.6151
R998 B.n525 B.n100 10.6151
R999 B.n526 B.n525 10.6151
R1000 B.n527 B.n526 10.6151
R1001 B.n527 B.n98 10.6151
R1002 B.n531 B.n98 10.6151
R1003 B.n532 B.n531 10.6151
R1004 B.n533 B.n532 10.6151
R1005 B.n533 B.n96 10.6151
R1006 B.n537 B.n96 10.6151
R1007 B.n538 B.n537 10.6151
R1008 B.n539 B.n538 10.6151
R1009 B.n539 B.n94 10.6151
R1010 B.n543 B.n94 10.6151
R1011 B.n544 B.n543 10.6151
R1012 B.n545 B.n544 10.6151
R1013 B.n545 B.n92 10.6151
R1014 B.n549 B.n92 10.6151
R1015 B.n550 B.n549 10.6151
R1016 B.n251 B.n194 10.6151
R1017 B.n255 B.n194 10.6151
R1018 B.n256 B.n255 10.6151
R1019 B.n257 B.n256 10.6151
R1020 B.n257 B.n192 10.6151
R1021 B.n261 B.n192 10.6151
R1022 B.n262 B.n261 10.6151
R1023 B.n263 B.n262 10.6151
R1024 B.n263 B.n190 10.6151
R1025 B.n267 B.n190 10.6151
R1026 B.n268 B.n267 10.6151
R1027 B.n269 B.n268 10.6151
R1028 B.n269 B.n188 10.6151
R1029 B.n273 B.n188 10.6151
R1030 B.n274 B.n273 10.6151
R1031 B.n275 B.n274 10.6151
R1032 B.n275 B.n186 10.6151
R1033 B.n279 B.n186 10.6151
R1034 B.n280 B.n279 10.6151
R1035 B.n281 B.n280 10.6151
R1036 B.n281 B.n184 10.6151
R1037 B.n285 B.n184 10.6151
R1038 B.n286 B.n285 10.6151
R1039 B.n287 B.n286 10.6151
R1040 B.n287 B.n182 10.6151
R1041 B.n291 B.n182 10.6151
R1042 B.n292 B.n291 10.6151
R1043 B.n293 B.n292 10.6151
R1044 B.n293 B.n180 10.6151
R1045 B.n297 B.n180 10.6151
R1046 B.n298 B.n297 10.6151
R1047 B.n299 B.n298 10.6151
R1048 B.n299 B.n178 10.6151
R1049 B.n303 B.n178 10.6151
R1050 B.n304 B.n303 10.6151
R1051 B.n305 B.n304 10.6151
R1052 B.n305 B.n176 10.6151
R1053 B.n309 B.n176 10.6151
R1054 B.n310 B.n309 10.6151
R1055 B.n311 B.n310 10.6151
R1056 B.n311 B.n174 10.6151
R1057 B.n315 B.n174 10.6151
R1058 B.n316 B.n315 10.6151
R1059 B.n317 B.n316 10.6151
R1060 B.n317 B.n172 10.6151
R1061 B.n321 B.n172 10.6151
R1062 B.n322 B.n321 10.6151
R1063 B.n323 B.n322 10.6151
R1064 B.n323 B.n170 10.6151
R1065 B.n327 B.n170 10.6151
R1066 B.n328 B.n327 10.6151
R1067 B.n329 B.n328 10.6151
R1068 B.n329 B.n168 10.6151
R1069 B.n333 B.n168 10.6151
R1070 B.n334 B.n333 10.6151
R1071 B.n335 B.n334 10.6151
R1072 B.n335 B.n166 10.6151
R1073 B.n339 B.n166 10.6151
R1074 B.n340 B.n339 10.6151
R1075 B.n341 B.n340 10.6151
R1076 B.n341 B.n164 10.6151
R1077 B.n345 B.n164 10.6151
R1078 B.n346 B.n345 10.6151
R1079 B.n347 B.n346 10.6151
R1080 B.n351 B.n350 10.6151
R1081 B.n352 B.n351 10.6151
R1082 B.n352 B.n158 10.6151
R1083 B.n356 B.n158 10.6151
R1084 B.n357 B.n356 10.6151
R1085 B.n358 B.n357 10.6151
R1086 B.n358 B.n156 10.6151
R1087 B.n362 B.n156 10.6151
R1088 B.n363 B.n362 10.6151
R1089 B.n365 B.n152 10.6151
R1090 B.n369 B.n152 10.6151
R1091 B.n370 B.n369 10.6151
R1092 B.n371 B.n370 10.6151
R1093 B.n371 B.n150 10.6151
R1094 B.n375 B.n150 10.6151
R1095 B.n376 B.n375 10.6151
R1096 B.n377 B.n376 10.6151
R1097 B.n377 B.n148 10.6151
R1098 B.n381 B.n148 10.6151
R1099 B.n382 B.n381 10.6151
R1100 B.n383 B.n382 10.6151
R1101 B.n383 B.n146 10.6151
R1102 B.n387 B.n146 10.6151
R1103 B.n388 B.n387 10.6151
R1104 B.n389 B.n388 10.6151
R1105 B.n389 B.n144 10.6151
R1106 B.n393 B.n144 10.6151
R1107 B.n394 B.n393 10.6151
R1108 B.n395 B.n394 10.6151
R1109 B.n395 B.n142 10.6151
R1110 B.n399 B.n142 10.6151
R1111 B.n400 B.n399 10.6151
R1112 B.n401 B.n400 10.6151
R1113 B.n401 B.n140 10.6151
R1114 B.n405 B.n140 10.6151
R1115 B.n406 B.n405 10.6151
R1116 B.n407 B.n406 10.6151
R1117 B.n407 B.n138 10.6151
R1118 B.n411 B.n138 10.6151
R1119 B.n412 B.n411 10.6151
R1120 B.n413 B.n412 10.6151
R1121 B.n413 B.n136 10.6151
R1122 B.n417 B.n136 10.6151
R1123 B.n418 B.n417 10.6151
R1124 B.n419 B.n418 10.6151
R1125 B.n419 B.n134 10.6151
R1126 B.n423 B.n134 10.6151
R1127 B.n424 B.n423 10.6151
R1128 B.n425 B.n424 10.6151
R1129 B.n425 B.n132 10.6151
R1130 B.n429 B.n132 10.6151
R1131 B.n430 B.n429 10.6151
R1132 B.n431 B.n430 10.6151
R1133 B.n431 B.n130 10.6151
R1134 B.n435 B.n130 10.6151
R1135 B.n436 B.n435 10.6151
R1136 B.n437 B.n436 10.6151
R1137 B.n437 B.n128 10.6151
R1138 B.n441 B.n128 10.6151
R1139 B.n442 B.n441 10.6151
R1140 B.n443 B.n442 10.6151
R1141 B.n443 B.n126 10.6151
R1142 B.n447 B.n126 10.6151
R1143 B.n448 B.n447 10.6151
R1144 B.n449 B.n448 10.6151
R1145 B.n449 B.n124 10.6151
R1146 B.n453 B.n124 10.6151
R1147 B.n454 B.n453 10.6151
R1148 B.n455 B.n454 10.6151
R1149 B.n455 B.n122 10.6151
R1150 B.n459 B.n122 10.6151
R1151 B.n460 B.n459 10.6151
R1152 B.n461 B.n460 10.6151
R1153 B.n250 B.n249 10.6151
R1154 B.n249 B.n196 10.6151
R1155 B.n245 B.n196 10.6151
R1156 B.n245 B.n244 10.6151
R1157 B.n244 B.n243 10.6151
R1158 B.n243 B.n198 10.6151
R1159 B.n239 B.n198 10.6151
R1160 B.n239 B.n238 10.6151
R1161 B.n238 B.n237 10.6151
R1162 B.n237 B.n200 10.6151
R1163 B.n233 B.n200 10.6151
R1164 B.n233 B.n232 10.6151
R1165 B.n232 B.n231 10.6151
R1166 B.n231 B.n202 10.6151
R1167 B.n227 B.n202 10.6151
R1168 B.n227 B.n226 10.6151
R1169 B.n226 B.n225 10.6151
R1170 B.n225 B.n204 10.6151
R1171 B.n221 B.n204 10.6151
R1172 B.n221 B.n220 10.6151
R1173 B.n220 B.n219 10.6151
R1174 B.n219 B.n206 10.6151
R1175 B.n215 B.n206 10.6151
R1176 B.n215 B.n214 10.6151
R1177 B.n214 B.n213 10.6151
R1178 B.n213 B.n208 10.6151
R1179 B.n209 B.n208 10.6151
R1180 B.n209 B.n0 10.6151
R1181 B.n803 B.n1 10.6151
R1182 B.n803 B.n802 10.6151
R1183 B.n802 B.n801 10.6151
R1184 B.n801 B.n4 10.6151
R1185 B.n797 B.n4 10.6151
R1186 B.n797 B.n796 10.6151
R1187 B.n796 B.n795 10.6151
R1188 B.n795 B.n6 10.6151
R1189 B.n791 B.n6 10.6151
R1190 B.n791 B.n790 10.6151
R1191 B.n790 B.n789 10.6151
R1192 B.n789 B.n8 10.6151
R1193 B.n785 B.n8 10.6151
R1194 B.n785 B.n784 10.6151
R1195 B.n784 B.n783 10.6151
R1196 B.n783 B.n10 10.6151
R1197 B.n779 B.n10 10.6151
R1198 B.n779 B.n778 10.6151
R1199 B.n778 B.n777 10.6151
R1200 B.n777 B.n12 10.6151
R1201 B.n773 B.n12 10.6151
R1202 B.n773 B.n772 10.6151
R1203 B.n772 B.n771 10.6151
R1204 B.n771 B.n14 10.6151
R1205 B.n767 B.n14 10.6151
R1206 B.n767 B.n766 10.6151
R1207 B.n766 B.n765 10.6151
R1208 B.n765 B.n16 10.6151
R1209 B.n665 B.n664 9.36635
R1210 B.n647 B.n58 9.36635
R1211 B.n347 B.n162 9.36635
R1212 B.n365 B.n364 9.36635
R1213 B.n807 B.n0 2.81026
R1214 B.n807 B.n1 2.81026
R1215 B.n664 B.n663 1.24928
R1216 B.n650 B.n58 1.24928
R1217 B.n350 B.n162 1.24928
R1218 B.n364 B.n363 1.24928
R1219 VN.n0 VN.t1 268.887
R1220 VN.n1 VN.t2 268.887
R1221 VN.n0 VN.t0 268.344
R1222 VN.n1 VN.t3 268.344
R1223 VN VN.n1 58.0394
R1224 VN VN.n0 6.99771
R1225 VTAIL.n6 VTAIL.t3 52.1522
R1226 VTAIL.n5 VTAIL.t0 52.1522
R1227 VTAIL.n4 VTAIL.t6 52.1522
R1228 VTAIL.n3 VTAIL.t5 52.1522
R1229 VTAIL.n7 VTAIL.t7 52.152
R1230 VTAIL.n0 VTAIL.t4 52.152
R1231 VTAIL.n1 VTAIL.t1 52.152
R1232 VTAIL.n2 VTAIL.t2 52.152
R1233 VTAIL.n7 VTAIL.n6 31.6772
R1234 VTAIL.n3 VTAIL.n2 31.6772
R1235 VTAIL.n4 VTAIL.n3 2.06947
R1236 VTAIL.n6 VTAIL.n5 2.06947
R1237 VTAIL.n2 VTAIL.n1 2.06947
R1238 VTAIL VTAIL.n0 1.09317
R1239 VTAIL VTAIL.n7 0.976793
R1240 VTAIL.n5 VTAIL.n4 0.470328
R1241 VTAIL.n1 VTAIL.n0 0.470328
R1242 VDD2.n2 VDD2.n0 114.368
R1243 VDD2.n2 VDD2.n1 67.2058
R1244 VDD2.n1 VDD2.t0 1.62575
R1245 VDD2.n1 VDD2.t1 1.62575
R1246 VDD2.n0 VDD2.t2 1.62575
R1247 VDD2.n0 VDD2.t3 1.62575
R1248 VDD2 VDD2.n2 0.0586897
R1249 VP.n2 VP.t1 268.887
R1250 VP.n2 VP.t0 268.344
R1251 VP.n4 VP.t3 232.851
R1252 VP.n11 VP.t2 232.851
R1253 VP.n10 VP.n0 161.3
R1254 VP.n9 VP.n8 161.3
R1255 VP.n7 VP.n1 161.3
R1256 VP.n6 VP.n5 161.3
R1257 VP.n4 VP.n3 88.7756
R1258 VP.n12 VP.n11 88.7756
R1259 VP.n3 VP.n2 57.7605
R1260 VP.n9 VP.n1 56.5617
R1261 VP.n5 VP.n1 24.5923
R1262 VP.n10 VP.n9 24.5923
R1263 VP.n5 VP.n4 22.1332
R1264 VP.n11 VP.n10 22.1332
R1265 VP.n6 VP.n3 0.278335
R1266 VP.n12 VP.n0 0.278335
R1267 VP.n7 VP.n6 0.189894
R1268 VP.n8 VP.n7 0.189894
R1269 VP.n8 VP.n0 0.189894
R1270 VP VP.n12 0.153485
R1271 VDD1 VDD1.n1 114.894
R1272 VDD1 VDD1.n0 67.264
R1273 VDD1.n0 VDD1.t2 1.62575
R1274 VDD1.n0 VDD1.t3 1.62575
R1275 VDD1.n1 VDD1.t0 1.62575
R1276 VDD1.n1 VDD1.t1 1.62575
C0 VN w_n2410_n4968# 4.1246f
C1 VDD2 VTAIL 7.51251f
C2 VDD1 VDD2 0.901321f
C3 VN VTAIL 6.86074f
C4 VN VDD1 0.148981f
C5 w_n2410_n4968# VP 4.43307f
C6 VP VTAIL 6.87484f
C7 VDD1 VP 7.56934f
C8 B VDD2 1.42834f
C9 VN B 1.10543f
C10 VN VDD2 7.35788f
C11 B VP 1.61486f
C12 VDD2 VP 0.361041f
C13 VN VP 7.28595f
C14 w_n2410_n4968# VTAIL 5.80603f
C15 VDD1 w_n2410_n4968# 1.56678f
C16 VDD1 VTAIL 7.46186f
C17 B w_n2410_n4968# 10.836901f
C18 B VTAIL 7.22583f
C19 VDD1 B 1.38488f
C20 VDD2 w_n2410_n4968# 1.61105f
C21 VDD2 VSUBS 1.050461f
C22 VDD1 VSUBS 6.49484f
C23 VTAIL VSUBS 1.54431f
C24 VN VSUBS 5.6311f
C25 VP VSUBS 2.310519f
C26 B VSUBS 4.490677f
C27 w_n2410_n4968# VSUBS 0.146191p
C28 VDD1.t2 VSUBS 0.420996f
C29 VDD1.t3 VSUBS 0.420996f
C30 VDD1.n0 VSUBS 3.53598f
C31 VDD1.t0 VSUBS 0.420996f
C32 VDD1.t1 VSUBS 0.420996f
C33 VDD1.n1 VSUBS 4.58785f
C34 VP.n0 VSUBS 0.044921f
C35 VP.t2 VSUBS 3.88747f
C36 VP.n1 VSUBS 0.049532f
C37 VP.t0 VSUBS 4.09022f
C38 VP.t1 VSUBS 4.09331f
C39 VP.n2 VSUBS 4.64811f
C40 VP.n3 VSUBS 2.2113f
C41 VP.t3 VSUBS 3.88747f
C42 VP.n4 VSUBS 1.46117f
C43 VP.n5 VSUBS 0.060068f
C44 VP.n6 VSUBS 0.044921f
C45 VP.n7 VSUBS 0.034074f
C46 VP.n8 VSUBS 0.034074f
C47 VP.n9 VSUBS 0.049532f
C48 VP.n10 VSUBS 0.060068f
C49 VP.n11 VSUBS 1.46117f
C50 VP.n12 VSUBS 0.039341f
C51 VDD2.t2 VSUBS 0.418144f
C52 VDD2.t3 VSUBS 0.418144f
C53 VDD2.n0 VSUBS 4.52854f
C54 VDD2.t0 VSUBS 0.418144f
C55 VDD2.t1 VSUBS 0.418144f
C56 VDD2.n1 VSUBS 3.5114f
C57 VDD2.n2 VSUBS 5.00541f
C58 VTAIL.t4 VSUBS 3.5799f
C59 VTAIL.n0 VSUBS 0.767909f
C60 VTAIL.t1 VSUBS 3.5799f
C61 VTAIL.n1 VSUBS 0.836397f
C62 VTAIL.t2 VSUBS 3.5799f
C63 VTAIL.n2 VSUBS 2.45381f
C64 VTAIL.t5 VSUBS 3.57992f
C65 VTAIL.n3 VSUBS 2.45378f
C66 VTAIL.t6 VSUBS 3.57992f
C67 VTAIL.n4 VSUBS 0.836371f
C68 VTAIL.t0 VSUBS 3.57992f
C69 VTAIL.n5 VSUBS 0.836371f
C70 VTAIL.t3 VSUBS 3.57991f
C71 VTAIL.n6 VSUBS 2.45379f
C72 VTAIL.t7 VSUBS 3.5799f
C73 VTAIL.n7 VSUBS 2.37716f
C74 VN.t1 VSUBS 4.00786f
C75 VN.t0 VSUBS 4.00484f
C76 VN.n0 VSUBS 2.69f
C77 VN.t2 VSUBS 4.00786f
C78 VN.t3 VSUBS 4.00484f
C79 VN.n1 VSUBS 4.56806f
C80 B.n0 VSUBS 0.00395f
C81 B.n1 VSUBS 0.00395f
C82 B.n2 VSUBS 0.006246f
C83 B.n3 VSUBS 0.006246f
C84 B.n4 VSUBS 0.006246f
C85 B.n5 VSUBS 0.006246f
C86 B.n6 VSUBS 0.006246f
C87 B.n7 VSUBS 0.006246f
C88 B.n8 VSUBS 0.006246f
C89 B.n9 VSUBS 0.006246f
C90 B.n10 VSUBS 0.006246f
C91 B.n11 VSUBS 0.006246f
C92 B.n12 VSUBS 0.006246f
C93 B.n13 VSUBS 0.006246f
C94 B.n14 VSUBS 0.006246f
C95 B.n15 VSUBS 0.006246f
C96 B.n16 VSUBS 0.014715f
C97 B.n17 VSUBS 0.006246f
C98 B.n18 VSUBS 0.006246f
C99 B.n19 VSUBS 0.006246f
C100 B.n20 VSUBS 0.006246f
C101 B.n21 VSUBS 0.006246f
C102 B.n22 VSUBS 0.006246f
C103 B.n23 VSUBS 0.006246f
C104 B.n24 VSUBS 0.006246f
C105 B.n25 VSUBS 0.006246f
C106 B.n26 VSUBS 0.006246f
C107 B.n27 VSUBS 0.006246f
C108 B.n28 VSUBS 0.006246f
C109 B.n29 VSUBS 0.006246f
C110 B.n30 VSUBS 0.006246f
C111 B.n31 VSUBS 0.006246f
C112 B.n32 VSUBS 0.006246f
C113 B.n33 VSUBS 0.006246f
C114 B.n34 VSUBS 0.006246f
C115 B.n35 VSUBS 0.006246f
C116 B.n36 VSUBS 0.006246f
C117 B.n37 VSUBS 0.006246f
C118 B.n38 VSUBS 0.006246f
C119 B.n39 VSUBS 0.006246f
C120 B.n40 VSUBS 0.006246f
C121 B.n41 VSUBS 0.006246f
C122 B.n42 VSUBS 0.006246f
C123 B.n43 VSUBS 0.006246f
C124 B.n44 VSUBS 0.006246f
C125 B.n45 VSUBS 0.006246f
C126 B.n46 VSUBS 0.006246f
C127 B.n47 VSUBS 0.006246f
C128 B.n48 VSUBS 0.006246f
C129 B.n49 VSUBS 0.006246f
C130 B.t11 VSUBS 0.606692f
C131 B.t10 VSUBS 0.62246f
C132 B.t9 VSUBS 1.59872f
C133 B.n50 VSUBS 0.316605f
C134 B.n51 VSUBS 0.062427f
C135 B.n52 VSUBS 0.006246f
C136 B.n53 VSUBS 0.006246f
C137 B.n54 VSUBS 0.006246f
C138 B.n55 VSUBS 0.006246f
C139 B.t5 VSUBS 0.606667f
C140 B.t4 VSUBS 0.62244f
C141 B.t3 VSUBS 1.59872f
C142 B.n56 VSUBS 0.316626f
C143 B.n57 VSUBS 0.062452f
C144 B.n58 VSUBS 0.014471f
C145 B.n59 VSUBS 0.006246f
C146 B.n60 VSUBS 0.006246f
C147 B.n61 VSUBS 0.006246f
C148 B.n62 VSUBS 0.006246f
C149 B.n63 VSUBS 0.006246f
C150 B.n64 VSUBS 0.006246f
C151 B.n65 VSUBS 0.006246f
C152 B.n66 VSUBS 0.006246f
C153 B.n67 VSUBS 0.006246f
C154 B.n68 VSUBS 0.006246f
C155 B.n69 VSUBS 0.006246f
C156 B.n70 VSUBS 0.006246f
C157 B.n71 VSUBS 0.006246f
C158 B.n72 VSUBS 0.006246f
C159 B.n73 VSUBS 0.006246f
C160 B.n74 VSUBS 0.006246f
C161 B.n75 VSUBS 0.006246f
C162 B.n76 VSUBS 0.006246f
C163 B.n77 VSUBS 0.006246f
C164 B.n78 VSUBS 0.006246f
C165 B.n79 VSUBS 0.006246f
C166 B.n80 VSUBS 0.006246f
C167 B.n81 VSUBS 0.006246f
C168 B.n82 VSUBS 0.006246f
C169 B.n83 VSUBS 0.006246f
C170 B.n84 VSUBS 0.006246f
C171 B.n85 VSUBS 0.006246f
C172 B.n86 VSUBS 0.006246f
C173 B.n87 VSUBS 0.006246f
C174 B.n88 VSUBS 0.006246f
C175 B.n89 VSUBS 0.006246f
C176 B.n90 VSUBS 0.006246f
C177 B.n91 VSUBS 0.014715f
C178 B.n92 VSUBS 0.006246f
C179 B.n93 VSUBS 0.006246f
C180 B.n94 VSUBS 0.006246f
C181 B.n95 VSUBS 0.006246f
C182 B.n96 VSUBS 0.006246f
C183 B.n97 VSUBS 0.006246f
C184 B.n98 VSUBS 0.006246f
C185 B.n99 VSUBS 0.006246f
C186 B.n100 VSUBS 0.006246f
C187 B.n101 VSUBS 0.006246f
C188 B.n102 VSUBS 0.006246f
C189 B.n103 VSUBS 0.006246f
C190 B.n104 VSUBS 0.006246f
C191 B.n105 VSUBS 0.006246f
C192 B.n106 VSUBS 0.006246f
C193 B.n107 VSUBS 0.006246f
C194 B.n108 VSUBS 0.006246f
C195 B.n109 VSUBS 0.006246f
C196 B.n110 VSUBS 0.006246f
C197 B.n111 VSUBS 0.006246f
C198 B.n112 VSUBS 0.006246f
C199 B.n113 VSUBS 0.006246f
C200 B.n114 VSUBS 0.006246f
C201 B.n115 VSUBS 0.006246f
C202 B.n116 VSUBS 0.006246f
C203 B.n117 VSUBS 0.006246f
C204 B.n118 VSUBS 0.006246f
C205 B.n119 VSUBS 0.006246f
C206 B.n120 VSUBS 0.014715f
C207 B.n121 VSUBS 0.006246f
C208 B.n122 VSUBS 0.006246f
C209 B.n123 VSUBS 0.006246f
C210 B.n124 VSUBS 0.006246f
C211 B.n125 VSUBS 0.006246f
C212 B.n126 VSUBS 0.006246f
C213 B.n127 VSUBS 0.006246f
C214 B.n128 VSUBS 0.006246f
C215 B.n129 VSUBS 0.006246f
C216 B.n130 VSUBS 0.006246f
C217 B.n131 VSUBS 0.006246f
C218 B.n132 VSUBS 0.006246f
C219 B.n133 VSUBS 0.006246f
C220 B.n134 VSUBS 0.006246f
C221 B.n135 VSUBS 0.006246f
C222 B.n136 VSUBS 0.006246f
C223 B.n137 VSUBS 0.006246f
C224 B.n138 VSUBS 0.006246f
C225 B.n139 VSUBS 0.006246f
C226 B.n140 VSUBS 0.006246f
C227 B.n141 VSUBS 0.006246f
C228 B.n142 VSUBS 0.006246f
C229 B.n143 VSUBS 0.006246f
C230 B.n144 VSUBS 0.006246f
C231 B.n145 VSUBS 0.006246f
C232 B.n146 VSUBS 0.006246f
C233 B.n147 VSUBS 0.006246f
C234 B.n148 VSUBS 0.006246f
C235 B.n149 VSUBS 0.006246f
C236 B.n150 VSUBS 0.006246f
C237 B.n151 VSUBS 0.006246f
C238 B.n152 VSUBS 0.006246f
C239 B.n153 VSUBS 0.006246f
C240 B.t1 VSUBS 0.606667f
C241 B.t2 VSUBS 0.62244f
C242 B.t0 VSUBS 1.59872f
C243 B.n154 VSUBS 0.316626f
C244 B.n155 VSUBS 0.062452f
C245 B.n156 VSUBS 0.006246f
C246 B.n157 VSUBS 0.006246f
C247 B.n158 VSUBS 0.006246f
C248 B.n159 VSUBS 0.006246f
C249 B.t7 VSUBS 0.606692f
C250 B.t8 VSUBS 0.62246f
C251 B.t6 VSUBS 1.59872f
C252 B.n160 VSUBS 0.316605f
C253 B.n161 VSUBS 0.062427f
C254 B.n162 VSUBS 0.014471f
C255 B.n163 VSUBS 0.006246f
C256 B.n164 VSUBS 0.006246f
C257 B.n165 VSUBS 0.006246f
C258 B.n166 VSUBS 0.006246f
C259 B.n167 VSUBS 0.006246f
C260 B.n168 VSUBS 0.006246f
C261 B.n169 VSUBS 0.006246f
C262 B.n170 VSUBS 0.006246f
C263 B.n171 VSUBS 0.006246f
C264 B.n172 VSUBS 0.006246f
C265 B.n173 VSUBS 0.006246f
C266 B.n174 VSUBS 0.006246f
C267 B.n175 VSUBS 0.006246f
C268 B.n176 VSUBS 0.006246f
C269 B.n177 VSUBS 0.006246f
C270 B.n178 VSUBS 0.006246f
C271 B.n179 VSUBS 0.006246f
C272 B.n180 VSUBS 0.006246f
C273 B.n181 VSUBS 0.006246f
C274 B.n182 VSUBS 0.006246f
C275 B.n183 VSUBS 0.006246f
C276 B.n184 VSUBS 0.006246f
C277 B.n185 VSUBS 0.006246f
C278 B.n186 VSUBS 0.006246f
C279 B.n187 VSUBS 0.006246f
C280 B.n188 VSUBS 0.006246f
C281 B.n189 VSUBS 0.006246f
C282 B.n190 VSUBS 0.006246f
C283 B.n191 VSUBS 0.006246f
C284 B.n192 VSUBS 0.006246f
C285 B.n193 VSUBS 0.006246f
C286 B.n194 VSUBS 0.006246f
C287 B.n195 VSUBS 0.014715f
C288 B.n196 VSUBS 0.006246f
C289 B.n197 VSUBS 0.006246f
C290 B.n198 VSUBS 0.006246f
C291 B.n199 VSUBS 0.006246f
C292 B.n200 VSUBS 0.006246f
C293 B.n201 VSUBS 0.006246f
C294 B.n202 VSUBS 0.006246f
C295 B.n203 VSUBS 0.006246f
C296 B.n204 VSUBS 0.006246f
C297 B.n205 VSUBS 0.006246f
C298 B.n206 VSUBS 0.006246f
C299 B.n207 VSUBS 0.006246f
C300 B.n208 VSUBS 0.006246f
C301 B.n209 VSUBS 0.006246f
C302 B.n210 VSUBS 0.006246f
C303 B.n211 VSUBS 0.006246f
C304 B.n212 VSUBS 0.006246f
C305 B.n213 VSUBS 0.006246f
C306 B.n214 VSUBS 0.006246f
C307 B.n215 VSUBS 0.006246f
C308 B.n216 VSUBS 0.006246f
C309 B.n217 VSUBS 0.006246f
C310 B.n218 VSUBS 0.006246f
C311 B.n219 VSUBS 0.006246f
C312 B.n220 VSUBS 0.006246f
C313 B.n221 VSUBS 0.006246f
C314 B.n222 VSUBS 0.006246f
C315 B.n223 VSUBS 0.006246f
C316 B.n224 VSUBS 0.006246f
C317 B.n225 VSUBS 0.006246f
C318 B.n226 VSUBS 0.006246f
C319 B.n227 VSUBS 0.006246f
C320 B.n228 VSUBS 0.006246f
C321 B.n229 VSUBS 0.006246f
C322 B.n230 VSUBS 0.006246f
C323 B.n231 VSUBS 0.006246f
C324 B.n232 VSUBS 0.006246f
C325 B.n233 VSUBS 0.006246f
C326 B.n234 VSUBS 0.006246f
C327 B.n235 VSUBS 0.006246f
C328 B.n236 VSUBS 0.006246f
C329 B.n237 VSUBS 0.006246f
C330 B.n238 VSUBS 0.006246f
C331 B.n239 VSUBS 0.006246f
C332 B.n240 VSUBS 0.006246f
C333 B.n241 VSUBS 0.006246f
C334 B.n242 VSUBS 0.006246f
C335 B.n243 VSUBS 0.006246f
C336 B.n244 VSUBS 0.006246f
C337 B.n245 VSUBS 0.006246f
C338 B.n246 VSUBS 0.006246f
C339 B.n247 VSUBS 0.006246f
C340 B.n248 VSUBS 0.006246f
C341 B.n249 VSUBS 0.006246f
C342 B.n250 VSUBS 0.014715f
C343 B.n251 VSUBS 0.015779f
C344 B.n252 VSUBS 0.015779f
C345 B.n253 VSUBS 0.006246f
C346 B.n254 VSUBS 0.006246f
C347 B.n255 VSUBS 0.006246f
C348 B.n256 VSUBS 0.006246f
C349 B.n257 VSUBS 0.006246f
C350 B.n258 VSUBS 0.006246f
C351 B.n259 VSUBS 0.006246f
C352 B.n260 VSUBS 0.006246f
C353 B.n261 VSUBS 0.006246f
C354 B.n262 VSUBS 0.006246f
C355 B.n263 VSUBS 0.006246f
C356 B.n264 VSUBS 0.006246f
C357 B.n265 VSUBS 0.006246f
C358 B.n266 VSUBS 0.006246f
C359 B.n267 VSUBS 0.006246f
C360 B.n268 VSUBS 0.006246f
C361 B.n269 VSUBS 0.006246f
C362 B.n270 VSUBS 0.006246f
C363 B.n271 VSUBS 0.006246f
C364 B.n272 VSUBS 0.006246f
C365 B.n273 VSUBS 0.006246f
C366 B.n274 VSUBS 0.006246f
C367 B.n275 VSUBS 0.006246f
C368 B.n276 VSUBS 0.006246f
C369 B.n277 VSUBS 0.006246f
C370 B.n278 VSUBS 0.006246f
C371 B.n279 VSUBS 0.006246f
C372 B.n280 VSUBS 0.006246f
C373 B.n281 VSUBS 0.006246f
C374 B.n282 VSUBS 0.006246f
C375 B.n283 VSUBS 0.006246f
C376 B.n284 VSUBS 0.006246f
C377 B.n285 VSUBS 0.006246f
C378 B.n286 VSUBS 0.006246f
C379 B.n287 VSUBS 0.006246f
C380 B.n288 VSUBS 0.006246f
C381 B.n289 VSUBS 0.006246f
C382 B.n290 VSUBS 0.006246f
C383 B.n291 VSUBS 0.006246f
C384 B.n292 VSUBS 0.006246f
C385 B.n293 VSUBS 0.006246f
C386 B.n294 VSUBS 0.006246f
C387 B.n295 VSUBS 0.006246f
C388 B.n296 VSUBS 0.006246f
C389 B.n297 VSUBS 0.006246f
C390 B.n298 VSUBS 0.006246f
C391 B.n299 VSUBS 0.006246f
C392 B.n300 VSUBS 0.006246f
C393 B.n301 VSUBS 0.006246f
C394 B.n302 VSUBS 0.006246f
C395 B.n303 VSUBS 0.006246f
C396 B.n304 VSUBS 0.006246f
C397 B.n305 VSUBS 0.006246f
C398 B.n306 VSUBS 0.006246f
C399 B.n307 VSUBS 0.006246f
C400 B.n308 VSUBS 0.006246f
C401 B.n309 VSUBS 0.006246f
C402 B.n310 VSUBS 0.006246f
C403 B.n311 VSUBS 0.006246f
C404 B.n312 VSUBS 0.006246f
C405 B.n313 VSUBS 0.006246f
C406 B.n314 VSUBS 0.006246f
C407 B.n315 VSUBS 0.006246f
C408 B.n316 VSUBS 0.006246f
C409 B.n317 VSUBS 0.006246f
C410 B.n318 VSUBS 0.006246f
C411 B.n319 VSUBS 0.006246f
C412 B.n320 VSUBS 0.006246f
C413 B.n321 VSUBS 0.006246f
C414 B.n322 VSUBS 0.006246f
C415 B.n323 VSUBS 0.006246f
C416 B.n324 VSUBS 0.006246f
C417 B.n325 VSUBS 0.006246f
C418 B.n326 VSUBS 0.006246f
C419 B.n327 VSUBS 0.006246f
C420 B.n328 VSUBS 0.006246f
C421 B.n329 VSUBS 0.006246f
C422 B.n330 VSUBS 0.006246f
C423 B.n331 VSUBS 0.006246f
C424 B.n332 VSUBS 0.006246f
C425 B.n333 VSUBS 0.006246f
C426 B.n334 VSUBS 0.006246f
C427 B.n335 VSUBS 0.006246f
C428 B.n336 VSUBS 0.006246f
C429 B.n337 VSUBS 0.006246f
C430 B.n338 VSUBS 0.006246f
C431 B.n339 VSUBS 0.006246f
C432 B.n340 VSUBS 0.006246f
C433 B.n341 VSUBS 0.006246f
C434 B.n342 VSUBS 0.006246f
C435 B.n343 VSUBS 0.006246f
C436 B.n344 VSUBS 0.006246f
C437 B.n345 VSUBS 0.006246f
C438 B.n346 VSUBS 0.006246f
C439 B.n347 VSUBS 0.005879f
C440 B.n348 VSUBS 0.006246f
C441 B.n349 VSUBS 0.006246f
C442 B.n350 VSUBS 0.00349f
C443 B.n351 VSUBS 0.006246f
C444 B.n352 VSUBS 0.006246f
C445 B.n353 VSUBS 0.006246f
C446 B.n354 VSUBS 0.006246f
C447 B.n355 VSUBS 0.006246f
C448 B.n356 VSUBS 0.006246f
C449 B.n357 VSUBS 0.006246f
C450 B.n358 VSUBS 0.006246f
C451 B.n359 VSUBS 0.006246f
C452 B.n360 VSUBS 0.006246f
C453 B.n361 VSUBS 0.006246f
C454 B.n362 VSUBS 0.006246f
C455 B.n363 VSUBS 0.00349f
C456 B.n364 VSUBS 0.014471f
C457 B.n365 VSUBS 0.005879f
C458 B.n366 VSUBS 0.006246f
C459 B.n367 VSUBS 0.006246f
C460 B.n368 VSUBS 0.006246f
C461 B.n369 VSUBS 0.006246f
C462 B.n370 VSUBS 0.006246f
C463 B.n371 VSUBS 0.006246f
C464 B.n372 VSUBS 0.006246f
C465 B.n373 VSUBS 0.006246f
C466 B.n374 VSUBS 0.006246f
C467 B.n375 VSUBS 0.006246f
C468 B.n376 VSUBS 0.006246f
C469 B.n377 VSUBS 0.006246f
C470 B.n378 VSUBS 0.006246f
C471 B.n379 VSUBS 0.006246f
C472 B.n380 VSUBS 0.006246f
C473 B.n381 VSUBS 0.006246f
C474 B.n382 VSUBS 0.006246f
C475 B.n383 VSUBS 0.006246f
C476 B.n384 VSUBS 0.006246f
C477 B.n385 VSUBS 0.006246f
C478 B.n386 VSUBS 0.006246f
C479 B.n387 VSUBS 0.006246f
C480 B.n388 VSUBS 0.006246f
C481 B.n389 VSUBS 0.006246f
C482 B.n390 VSUBS 0.006246f
C483 B.n391 VSUBS 0.006246f
C484 B.n392 VSUBS 0.006246f
C485 B.n393 VSUBS 0.006246f
C486 B.n394 VSUBS 0.006246f
C487 B.n395 VSUBS 0.006246f
C488 B.n396 VSUBS 0.006246f
C489 B.n397 VSUBS 0.006246f
C490 B.n398 VSUBS 0.006246f
C491 B.n399 VSUBS 0.006246f
C492 B.n400 VSUBS 0.006246f
C493 B.n401 VSUBS 0.006246f
C494 B.n402 VSUBS 0.006246f
C495 B.n403 VSUBS 0.006246f
C496 B.n404 VSUBS 0.006246f
C497 B.n405 VSUBS 0.006246f
C498 B.n406 VSUBS 0.006246f
C499 B.n407 VSUBS 0.006246f
C500 B.n408 VSUBS 0.006246f
C501 B.n409 VSUBS 0.006246f
C502 B.n410 VSUBS 0.006246f
C503 B.n411 VSUBS 0.006246f
C504 B.n412 VSUBS 0.006246f
C505 B.n413 VSUBS 0.006246f
C506 B.n414 VSUBS 0.006246f
C507 B.n415 VSUBS 0.006246f
C508 B.n416 VSUBS 0.006246f
C509 B.n417 VSUBS 0.006246f
C510 B.n418 VSUBS 0.006246f
C511 B.n419 VSUBS 0.006246f
C512 B.n420 VSUBS 0.006246f
C513 B.n421 VSUBS 0.006246f
C514 B.n422 VSUBS 0.006246f
C515 B.n423 VSUBS 0.006246f
C516 B.n424 VSUBS 0.006246f
C517 B.n425 VSUBS 0.006246f
C518 B.n426 VSUBS 0.006246f
C519 B.n427 VSUBS 0.006246f
C520 B.n428 VSUBS 0.006246f
C521 B.n429 VSUBS 0.006246f
C522 B.n430 VSUBS 0.006246f
C523 B.n431 VSUBS 0.006246f
C524 B.n432 VSUBS 0.006246f
C525 B.n433 VSUBS 0.006246f
C526 B.n434 VSUBS 0.006246f
C527 B.n435 VSUBS 0.006246f
C528 B.n436 VSUBS 0.006246f
C529 B.n437 VSUBS 0.006246f
C530 B.n438 VSUBS 0.006246f
C531 B.n439 VSUBS 0.006246f
C532 B.n440 VSUBS 0.006246f
C533 B.n441 VSUBS 0.006246f
C534 B.n442 VSUBS 0.006246f
C535 B.n443 VSUBS 0.006246f
C536 B.n444 VSUBS 0.006246f
C537 B.n445 VSUBS 0.006246f
C538 B.n446 VSUBS 0.006246f
C539 B.n447 VSUBS 0.006246f
C540 B.n448 VSUBS 0.006246f
C541 B.n449 VSUBS 0.006246f
C542 B.n450 VSUBS 0.006246f
C543 B.n451 VSUBS 0.006246f
C544 B.n452 VSUBS 0.006246f
C545 B.n453 VSUBS 0.006246f
C546 B.n454 VSUBS 0.006246f
C547 B.n455 VSUBS 0.006246f
C548 B.n456 VSUBS 0.006246f
C549 B.n457 VSUBS 0.006246f
C550 B.n458 VSUBS 0.006246f
C551 B.n459 VSUBS 0.006246f
C552 B.n460 VSUBS 0.006246f
C553 B.n461 VSUBS 0.015779f
C554 B.n462 VSUBS 0.015779f
C555 B.n463 VSUBS 0.014715f
C556 B.n464 VSUBS 0.006246f
C557 B.n465 VSUBS 0.006246f
C558 B.n466 VSUBS 0.006246f
C559 B.n467 VSUBS 0.006246f
C560 B.n468 VSUBS 0.006246f
C561 B.n469 VSUBS 0.006246f
C562 B.n470 VSUBS 0.006246f
C563 B.n471 VSUBS 0.006246f
C564 B.n472 VSUBS 0.006246f
C565 B.n473 VSUBS 0.006246f
C566 B.n474 VSUBS 0.006246f
C567 B.n475 VSUBS 0.006246f
C568 B.n476 VSUBS 0.006246f
C569 B.n477 VSUBS 0.006246f
C570 B.n478 VSUBS 0.006246f
C571 B.n479 VSUBS 0.006246f
C572 B.n480 VSUBS 0.006246f
C573 B.n481 VSUBS 0.006246f
C574 B.n482 VSUBS 0.006246f
C575 B.n483 VSUBS 0.006246f
C576 B.n484 VSUBS 0.006246f
C577 B.n485 VSUBS 0.006246f
C578 B.n486 VSUBS 0.006246f
C579 B.n487 VSUBS 0.006246f
C580 B.n488 VSUBS 0.006246f
C581 B.n489 VSUBS 0.006246f
C582 B.n490 VSUBS 0.006246f
C583 B.n491 VSUBS 0.006246f
C584 B.n492 VSUBS 0.006246f
C585 B.n493 VSUBS 0.006246f
C586 B.n494 VSUBS 0.006246f
C587 B.n495 VSUBS 0.006246f
C588 B.n496 VSUBS 0.006246f
C589 B.n497 VSUBS 0.006246f
C590 B.n498 VSUBS 0.006246f
C591 B.n499 VSUBS 0.006246f
C592 B.n500 VSUBS 0.006246f
C593 B.n501 VSUBS 0.006246f
C594 B.n502 VSUBS 0.006246f
C595 B.n503 VSUBS 0.006246f
C596 B.n504 VSUBS 0.006246f
C597 B.n505 VSUBS 0.006246f
C598 B.n506 VSUBS 0.006246f
C599 B.n507 VSUBS 0.006246f
C600 B.n508 VSUBS 0.006246f
C601 B.n509 VSUBS 0.006246f
C602 B.n510 VSUBS 0.006246f
C603 B.n511 VSUBS 0.006246f
C604 B.n512 VSUBS 0.006246f
C605 B.n513 VSUBS 0.006246f
C606 B.n514 VSUBS 0.006246f
C607 B.n515 VSUBS 0.006246f
C608 B.n516 VSUBS 0.006246f
C609 B.n517 VSUBS 0.006246f
C610 B.n518 VSUBS 0.006246f
C611 B.n519 VSUBS 0.006246f
C612 B.n520 VSUBS 0.006246f
C613 B.n521 VSUBS 0.006246f
C614 B.n522 VSUBS 0.006246f
C615 B.n523 VSUBS 0.006246f
C616 B.n524 VSUBS 0.006246f
C617 B.n525 VSUBS 0.006246f
C618 B.n526 VSUBS 0.006246f
C619 B.n527 VSUBS 0.006246f
C620 B.n528 VSUBS 0.006246f
C621 B.n529 VSUBS 0.006246f
C622 B.n530 VSUBS 0.006246f
C623 B.n531 VSUBS 0.006246f
C624 B.n532 VSUBS 0.006246f
C625 B.n533 VSUBS 0.006246f
C626 B.n534 VSUBS 0.006246f
C627 B.n535 VSUBS 0.006246f
C628 B.n536 VSUBS 0.006246f
C629 B.n537 VSUBS 0.006246f
C630 B.n538 VSUBS 0.006246f
C631 B.n539 VSUBS 0.006246f
C632 B.n540 VSUBS 0.006246f
C633 B.n541 VSUBS 0.006246f
C634 B.n542 VSUBS 0.006246f
C635 B.n543 VSUBS 0.006246f
C636 B.n544 VSUBS 0.006246f
C637 B.n545 VSUBS 0.006246f
C638 B.n546 VSUBS 0.006246f
C639 B.n547 VSUBS 0.006246f
C640 B.n548 VSUBS 0.006246f
C641 B.n549 VSUBS 0.006246f
C642 B.n550 VSUBS 0.015408f
C643 B.n551 VSUBS 0.015087f
C644 B.n552 VSUBS 0.015779f
C645 B.n553 VSUBS 0.006246f
C646 B.n554 VSUBS 0.006246f
C647 B.n555 VSUBS 0.006246f
C648 B.n556 VSUBS 0.006246f
C649 B.n557 VSUBS 0.006246f
C650 B.n558 VSUBS 0.006246f
C651 B.n559 VSUBS 0.006246f
C652 B.n560 VSUBS 0.006246f
C653 B.n561 VSUBS 0.006246f
C654 B.n562 VSUBS 0.006246f
C655 B.n563 VSUBS 0.006246f
C656 B.n564 VSUBS 0.006246f
C657 B.n565 VSUBS 0.006246f
C658 B.n566 VSUBS 0.006246f
C659 B.n567 VSUBS 0.006246f
C660 B.n568 VSUBS 0.006246f
C661 B.n569 VSUBS 0.006246f
C662 B.n570 VSUBS 0.006246f
C663 B.n571 VSUBS 0.006246f
C664 B.n572 VSUBS 0.006246f
C665 B.n573 VSUBS 0.006246f
C666 B.n574 VSUBS 0.006246f
C667 B.n575 VSUBS 0.006246f
C668 B.n576 VSUBS 0.006246f
C669 B.n577 VSUBS 0.006246f
C670 B.n578 VSUBS 0.006246f
C671 B.n579 VSUBS 0.006246f
C672 B.n580 VSUBS 0.006246f
C673 B.n581 VSUBS 0.006246f
C674 B.n582 VSUBS 0.006246f
C675 B.n583 VSUBS 0.006246f
C676 B.n584 VSUBS 0.006246f
C677 B.n585 VSUBS 0.006246f
C678 B.n586 VSUBS 0.006246f
C679 B.n587 VSUBS 0.006246f
C680 B.n588 VSUBS 0.006246f
C681 B.n589 VSUBS 0.006246f
C682 B.n590 VSUBS 0.006246f
C683 B.n591 VSUBS 0.006246f
C684 B.n592 VSUBS 0.006246f
C685 B.n593 VSUBS 0.006246f
C686 B.n594 VSUBS 0.006246f
C687 B.n595 VSUBS 0.006246f
C688 B.n596 VSUBS 0.006246f
C689 B.n597 VSUBS 0.006246f
C690 B.n598 VSUBS 0.006246f
C691 B.n599 VSUBS 0.006246f
C692 B.n600 VSUBS 0.006246f
C693 B.n601 VSUBS 0.006246f
C694 B.n602 VSUBS 0.006246f
C695 B.n603 VSUBS 0.006246f
C696 B.n604 VSUBS 0.006246f
C697 B.n605 VSUBS 0.006246f
C698 B.n606 VSUBS 0.006246f
C699 B.n607 VSUBS 0.006246f
C700 B.n608 VSUBS 0.006246f
C701 B.n609 VSUBS 0.006246f
C702 B.n610 VSUBS 0.006246f
C703 B.n611 VSUBS 0.006246f
C704 B.n612 VSUBS 0.006246f
C705 B.n613 VSUBS 0.006246f
C706 B.n614 VSUBS 0.006246f
C707 B.n615 VSUBS 0.006246f
C708 B.n616 VSUBS 0.006246f
C709 B.n617 VSUBS 0.006246f
C710 B.n618 VSUBS 0.006246f
C711 B.n619 VSUBS 0.006246f
C712 B.n620 VSUBS 0.006246f
C713 B.n621 VSUBS 0.006246f
C714 B.n622 VSUBS 0.006246f
C715 B.n623 VSUBS 0.006246f
C716 B.n624 VSUBS 0.006246f
C717 B.n625 VSUBS 0.006246f
C718 B.n626 VSUBS 0.006246f
C719 B.n627 VSUBS 0.006246f
C720 B.n628 VSUBS 0.006246f
C721 B.n629 VSUBS 0.006246f
C722 B.n630 VSUBS 0.006246f
C723 B.n631 VSUBS 0.006246f
C724 B.n632 VSUBS 0.006246f
C725 B.n633 VSUBS 0.006246f
C726 B.n634 VSUBS 0.006246f
C727 B.n635 VSUBS 0.006246f
C728 B.n636 VSUBS 0.006246f
C729 B.n637 VSUBS 0.006246f
C730 B.n638 VSUBS 0.006246f
C731 B.n639 VSUBS 0.006246f
C732 B.n640 VSUBS 0.006246f
C733 B.n641 VSUBS 0.006246f
C734 B.n642 VSUBS 0.006246f
C735 B.n643 VSUBS 0.006246f
C736 B.n644 VSUBS 0.006246f
C737 B.n645 VSUBS 0.006246f
C738 B.n646 VSUBS 0.006246f
C739 B.n647 VSUBS 0.005879f
C740 B.n648 VSUBS 0.006246f
C741 B.n649 VSUBS 0.006246f
C742 B.n650 VSUBS 0.00349f
C743 B.n651 VSUBS 0.006246f
C744 B.n652 VSUBS 0.006246f
C745 B.n653 VSUBS 0.006246f
C746 B.n654 VSUBS 0.006246f
C747 B.n655 VSUBS 0.006246f
C748 B.n656 VSUBS 0.006246f
C749 B.n657 VSUBS 0.006246f
C750 B.n658 VSUBS 0.006246f
C751 B.n659 VSUBS 0.006246f
C752 B.n660 VSUBS 0.006246f
C753 B.n661 VSUBS 0.006246f
C754 B.n662 VSUBS 0.006246f
C755 B.n663 VSUBS 0.00349f
C756 B.n664 VSUBS 0.014471f
C757 B.n665 VSUBS 0.005879f
C758 B.n666 VSUBS 0.006246f
C759 B.n667 VSUBS 0.006246f
C760 B.n668 VSUBS 0.006246f
C761 B.n669 VSUBS 0.006246f
C762 B.n670 VSUBS 0.006246f
C763 B.n671 VSUBS 0.006246f
C764 B.n672 VSUBS 0.006246f
C765 B.n673 VSUBS 0.006246f
C766 B.n674 VSUBS 0.006246f
C767 B.n675 VSUBS 0.006246f
C768 B.n676 VSUBS 0.006246f
C769 B.n677 VSUBS 0.006246f
C770 B.n678 VSUBS 0.006246f
C771 B.n679 VSUBS 0.006246f
C772 B.n680 VSUBS 0.006246f
C773 B.n681 VSUBS 0.006246f
C774 B.n682 VSUBS 0.006246f
C775 B.n683 VSUBS 0.006246f
C776 B.n684 VSUBS 0.006246f
C777 B.n685 VSUBS 0.006246f
C778 B.n686 VSUBS 0.006246f
C779 B.n687 VSUBS 0.006246f
C780 B.n688 VSUBS 0.006246f
C781 B.n689 VSUBS 0.006246f
C782 B.n690 VSUBS 0.006246f
C783 B.n691 VSUBS 0.006246f
C784 B.n692 VSUBS 0.006246f
C785 B.n693 VSUBS 0.006246f
C786 B.n694 VSUBS 0.006246f
C787 B.n695 VSUBS 0.006246f
C788 B.n696 VSUBS 0.006246f
C789 B.n697 VSUBS 0.006246f
C790 B.n698 VSUBS 0.006246f
C791 B.n699 VSUBS 0.006246f
C792 B.n700 VSUBS 0.006246f
C793 B.n701 VSUBS 0.006246f
C794 B.n702 VSUBS 0.006246f
C795 B.n703 VSUBS 0.006246f
C796 B.n704 VSUBS 0.006246f
C797 B.n705 VSUBS 0.006246f
C798 B.n706 VSUBS 0.006246f
C799 B.n707 VSUBS 0.006246f
C800 B.n708 VSUBS 0.006246f
C801 B.n709 VSUBS 0.006246f
C802 B.n710 VSUBS 0.006246f
C803 B.n711 VSUBS 0.006246f
C804 B.n712 VSUBS 0.006246f
C805 B.n713 VSUBS 0.006246f
C806 B.n714 VSUBS 0.006246f
C807 B.n715 VSUBS 0.006246f
C808 B.n716 VSUBS 0.006246f
C809 B.n717 VSUBS 0.006246f
C810 B.n718 VSUBS 0.006246f
C811 B.n719 VSUBS 0.006246f
C812 B.n720 VSUBS 0.006246f
C813 B.n721 VSUBS 0.006246f
C814 B.n722 VSUBS 0.006246f
C815 B.n723 VSUBS 0.006246f
C816 B.n724 VSUBS 0.006246f
C817 B.n725 VSUBS 0.006246f
C818 B.n726 VSUBS 0.006246f
C819 B.n727 VSUBS 0.006246f
C820 B.n728 VSUBS 0.006246f
C821 B.n729 VSUBS 0.006246f
C822 B.n730 VSUBS 0.006246f
C823 B.n731 VSUBS 0.006246f
C824 B.n732 VSUBS 0.006246f
C825 B.n733 VSUBS 0.006246f
C826 B.n734 VSUBS 0.006246f
C827 B.n735 VSUBS 0.006246f
C828 B.n736 VSUBS 0.006246f
C829 B.n737 VSUBS 0.006246f
C830 B.n738 VSUBS 0.006246f
C831 B.n739 VSUBS 0.006246f
C832 B.n740 VSUBS 0.006246f
C833 B.n741 VSUBS 0.006246f
C834 B.n742 VSUBS 0.006246f
C835 B.n743 VSUBS 0.006246f
C836 B.n744 VSUBS 0.006246f
C837 B.n745 VSUBS 0.006246f
C838 B.n746 VSUBS 0.006246f
C839 B.n747 VSUBS 0.006246f
C840 B.n748 VSUBS 0.006246f
C841 B.n749 VSUBS 0.006246f
C842 B.n750 VSUBS 0.006246f
C843 B.n751 VSUBS 0.006246f
C844 B.n752 VSUBS 0.006246f
C845 B.n753 VSUBS 0.006246f
C846 B.n754 VSUBS 0.006246f
C847 B.n755 VSUBS 0.006246f
C848 B.n756 VSUBS 0.006246f
C849 B.n757 VSUBS 0.006246f
C850 B.n758 VSUBS 0.006246f
C851 B.n759 VSUBS 0.006246f
C852 B.n760 VSUBS 0.006246f
C853 B.n761 VSUBS 0.015779f
C854 B.n762 VSUBS 0.015779f
C855 B.n763 VSUBS 0.014715f
C856 B.n764 VSUBS 0.006246f
C857 B.n765 VSUBS 0.006246f
C858 B.n766 VSUBS 0.006246f
C859 B.n767 VSUBS 0.006246f
C860 B.n768 VSUBS 0.006246f
C861 B.n769 VSUBS 0.006246f
C862 B.n770 VSUBS 0.006246f
C863 B.n771 VSUBS 0.006246f
C864 B.n772 VSUBS 0.006246f
C865 B.n773 VSUBS 0.006246f
C866 B.n774 VSUBS 0.006246f
C867 B.n775 VSUBS 0.006246f
C868 B.n776 VSUBS 0.006246f
C869 B.n777 VSUBS 0.006246f
C870 B.n778 VSUBS 0.006246f
C871 B.n779 VSUBS 0.006246f
C872 B.n780 VSUBS 0.006246f
C873 B.n781 VSUBS 0.006246f
C874 B.n782 VSUBS 0.006246f
C875 B.n783 VSUBS 0.006246f
C876 B.n784 VSUBS 0.006246f
C877 B.n785 VSUBS 0.006246f
C878 B.n786 VSUBS 0.006246f
C879 B.n787 VSUBS 0.006246f
C880 B.n788 VSUBS 0.006246f
C881 B.n789 VSUBS 0.006246f
C882 B.n790 VSUBS 0.006246f
C883 B.n791 VSUBS 0.006246f
C884 B.n792 VSUBS 0.006246f
C885 B.n793 VSUBS 0.006246f
C886 B.n794 VSUBS 0.006246f
C887 B.n795 VSUBS 0.006246f
C888 B.n796 VSUBS 0.006246f
C889 B.n797 VSUBS 0.006246f
C890 B.n798 VSUBS 0.006246f
C891 B.n799 VSUBS 0.006246f
C892 B.n800 VSUBS 0.006246f
C893 B.n801 VSUBS 0.006246f
C894 B.n802 VSUBS 0.006246f
C895 B.n803 VSUBS 0.006246f
C896 B.n804 VSUBS 0.006246f
C897 B.n805 VSUBS 0.006246f
C898 B.n806 VSUBS 0.006246f
C899 B.n807 VSUBS 0.014143f
.ends

