* NGSPICE file created from diff_pair_sample_0695.ext - technology: sky130A

.subckt diff_pair_sample_0695 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=1.0527 ps=6.71 w=6.38 l=2
X1 VTAIL.t2 VP.t0 VDD1.t3 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=1.0527 ps=6.71 w=6.38 l=2
X2 VTAIL.t6 VN.t1 VDD2.t0 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=1.0527 ps=6.71 w=6.38 l=2
X3 VDD1.t2 VP.t1 VTAIL.t0 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=1.0527 pd=6.71 as=2.4882 ps=13.54 w=6.38 l=2
X4 VDD2.t3 VN.t2 VTAIL.t5 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=1.0527 pd=6.71 as=2.4882 ps=13.54 w=6.38 l=2
X5 B.t11 B.t9 B.t10 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=0 ps=0 w=6.38 l=2
X6 VDD1.t1 VP.t2 VTAIL.t1 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=1.0527 pd=6.71 as=2.4882 ps=13.54 w=6.38 l=2
X7 B.t8 B.t6 B.t7 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=0 ps=0 w=6.38 l=2
X8 VDD2.t1 VN.t3 VTAIL.t4 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=1.0527 pd=6.71 as=2.4882 ps=13.54 w=6.38 l=2
X9 B.t5 B.t3 B.t4 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=0 ps=0 w=6.38 l=2
X10 B.t2 B.t0 B.t1 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=0 ps=0 w=6.38 l=2
X11 VTAIL.t3 VP.t3 VDD1.t0 w_n2368_n2244# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=13.54 as=1.0527 ps=6.71 w=6.38 l=2
R0 VN.n0 VN.t1 112.546
R1 VN.n1 VN.t2 112.546
R2 VN.n0 VN.t3 112.013
R3 VN.n1 VN.t0 112.013
R4 VN VN.n1 47.7183
R5 VN VN.n0 7.25996
R6 VDD2.n2 VDD2.n0 125.856
R7 VDD2.n2 VDD2.n1 90.6162
R8 VDD2.n1 VDD2.t2 5.09533
R9 VDD2.n1 VDD2.t3 5.09533
R10 VDD2.n0 VDD2.t0 5.09533
R11 VDD2.n0 VDD2.t1 5.09533
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t2 79.0323
R14 VTAIL.n4 VTAIL.t5 79.0323
R15 VTAIL.n3 VTAIL.t7 79.0323
R16 VTAIL.n7 VTAIL.t4 79.0322
R17 VTAIL.n0 VTAIL.t6 79.0322
R18 VTAIL.n1 VTAIL.t0 79.0322
R19 VTAIL.n2 VTAIL.t3 79.0322
R20 VTAIL.n6 VTAIL.t1 79.0322
R21 VTAIL.n7 VTAIL.n6 19.8755
R22 VTAIL.n3 VTAIL.n2 19.8755
R23 VTAIL.n4 VTAIL.n3 2.00912
R24 VTAIL.n6 VTAIL.n5 2.00912
R25 VTAIL.n2 VTAIL.n1 2.00912
R26 VTAIL VTAIL.n0 1.063
R27 VTAIL VTAIL.n7 0.946621
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 VP.n10 VP.n0 161.3
R31 VP.n9 VP.n8 161.3
R32 VP.n7 VP.n1 161.3
R33 VP.n6 VP.n5 161.3
R34 VP.n2 VP.t0 112.546
R35 VP.n2 VP.t2 112.013
R36 VP.n4 VP.n3 90.497
R37 VP.n12 VP.n11 90.497
R38 VP.n4 VP.t3 76.8795
R39 VP.n11 VP.t1 76.8795
R40 VP.n9 VP.n1 56.5617
R41 VP.n3 VP.n2 47.4395
R42 VP.n5 VP.n1 24.5923
R43 VP.n10 VP.n9 24.5923
R44 VP.n5 VP.n4 20.4117
R45 VP.n11 VP.n10 20.4117
R46 VP.n6 VP.n3 0.278335
R47 VP.n12 VP.n0 0.278335
R48 VP.n7 VP.n6 0.189894
R49 VP.n8 VP.n7 0.189894
R50 VP.n8 VP.n0 0.189894
R51 VP VP.n12 0.153485
R52 VDD1 VDD1.n1 126.382
R53 VDD1 VDD1.n0 90.6743
R54 VDD1.n0 VDD1.t3 5.09533
R55 VDD1.n0 VDD1.t1 5.09533
R56 VDD1.n1 VDD1.t0 5.09533
R57 VDD1.n1 VDD1.t2 5.09533
R58 B.n259 B.n80 585
R59 B.n258 B.n257 585
R60 B.n256 B.n81 585
R61 B.n255 B.n254 585
R62 B.n253 B.n82 585
R63 B.n252 B.n251 585
R64 B.n250 B.n83 585
R65 B.n249 B.n248 585
R66 B.n247 B.n84 585
R67 B.n246 B.n245 585
R68 B.n244 B.n85 585
R69 B.n243 B.n242 585
R70 B.n241 B.n86 585
R71 B.n240 B.n239 585
R72 B.n238 B.n87 585
R73 B.n237 B.n236 585
R74 B.n235 B.n88 585
R75 B.n234 B.n233 585
R76 B.n232 B.n89 585
R77 B.n231 B.n230 585
R78 B.n229 B.n90 585
R79 B.n228 B.n227 585
R80 B.n226 B.n91 585
R81 B.n225 B.n224 585
R82 B.n223 B.n92 585
R83 B.n221 B.n220 585
R84 B.n219 B.n95 585
R85 B.n218 B.n217 585
R86 B.n216 B.n96 585
R87 B.n215 B.n214 585
R88 B.n213 B.n97 585
R89 B.n212 B.n211 585
R90 B.n210 B.n98 585
R91 B.n209 B.n208 585
R92 B.n207 B.n99 585
R93 B.n206 B.n205 585
R94 B.n201 B.n100 585
R95 B.n200 B.n199 585
R96 B.n198 B.n101 585
R97 B.n197 B.n196 585
R98 B.n195 B.n102 585
R99 B.n194 B.n193 585
R100 B.n192 B.n103 585
R101 B.n191 B.n190 585
R102 B.n189 B.n104 585
R103 B.n188 B.n187 585
R104 B.n186 B.n105 585
R105 B.n185 B.n184 585
R106 B.n183 B.n106 585
R107 B.n182 B.n181 585
R108 B.n180 B.n107 585
R109 B.n179 B.n178 585
R110 B.n177 B.n108 585
R111 B.n176 B.n175 585
R112 B.n174 B.n109 585
R113 B.n173 B.n172 585
R114 B.n171 B.n110 585
R115 B.n170 B.n169 585
R116 B.n168 B.n111 585
R117 B.n167 B.n166 585
R118 B.n261 B.n260 585
R119 B.n262 B.n79 585
R120 B.n264 B.n263 585
R121 B.n265 B.n78 585
R122 B.n267 B.n266 585
R123 B.n268 B.n77 585
R124 B.n270 B.n269 585
R125 B.n271 B.n76 585
R126 B.n273 B.n272 585
R127 B.n274 B.n75 585
R128 B.n276 B.n275 585
R129 B.n277 B.n74 585
R130 B.n279 B.n278 585
R131 B.n280 B.n73 585
R132 B.n282 B.n281 585
R133 B.n283 B.n72 585
R134 B.n285 B.n284 585
R135 B.n286 B.n71 585
R136 B.n288 B.n287 585
R137 B.n289 B.n70 585
R138 B.n291 B.n290 585
R139 B.n292 B.n69 585
R140 B.n294 B.n293 585
R141 B.n295 B.n68 585
R142 B.n297 B.n296 585
R143 B.n298 B.n67 585
R144 B.n300 B.n299 585
R145 B.n301 B.n66 585
R146 B.n303 B.n302 585
R147 B.n304 B.n65 585
R148 B.n306 B.n305 585
R149 B.n307 B.n64 585
R150 B.n309 B.n308 585
R151 B.n310 B.n63 585
R152 B.n312 B.n311 585
R153 B.n313 B.n62 585
R154 B.n315 B.n314 585
R155 B.n316 B.n61 585
R156 B.n318 B.n317 585
R157 B.n319 B.n60 585
R158 B.n321 B.n320 585
R159 B.n322 B.n59 585
R160 B.n324 B.n323 585
R161 B.n325 B.n58 585
R162 B.n327 B.n326 585
R163 B.n328 B.n57 585
R164 B.n330 B.n329 585
R165 B.n331 B.n56 585
R166 B.n333 B.n332 585
R167 B.n334 B.n55 585
R168 B.n336 B.n335 585
R169 B.n337 B.n54 585
R170 B.n339 B.n338 585
R171 B.n340 B.n53 585
R172 B.n342 B.n341 585
R173 B.n343 B.n52 585
R174 B.n345 B.n344 585
R175 B.n346 B.n51 585
R176 B.n437 B.n16 585
R177 B.n436 B.n435 585
R178 B.n434 B.n17 585
R179 B.n433 B.n432 585
R180 B.n431 B.n18 585
R181 B.n430 B.n429 585
R182 B.n428 B.n19 585
R183 B.n427 B.n426 585
R184 B.n425 B.n20 585
R185 B.n424 B.n423 585
R186 B.n422 B.n21 585
R187 B.n421 B.n420 585
R188 B.n419 B.n22 585
R189 B.n418 B.n417 585
R190 B.n416 B.n23 585
R191 B.n415 B.n414 585
R192 B.n413 B.n24 585
R193 B.n412 B.n411 585
R194 B.n410 B.n25 585
R195 B.n409 B.n408 585
R196 B.n407 B.n26 585
R197 B.n406 B.n405 585
R198 B.n404 B.n27 585
R199 B.n403 B.n402 585
R200 B.n401 B.n28 585
R201 B.n400 B.n399 585
R202 B.n398 B.n29 585
R203 B.n397 B.n396 585
R204 B.n395 B.n33 585
R205 B.n394 B.n393 585
R206 B.n392 B.n34 585
R207 B.n391 B.n390 585
R208 B.n389 B.n35 585
R209 B.n388 B.n387 585
R210 B.n386 B.n36 585
R211 B.n384 B.n383 585
R212 B.n382 B.n39 585
R213 B.n381 B.n380 585
R214 B.n379 B.n40 585
R215 B.n378 B.n377 585
R216 B.n376 B.n41 585
R217 B.n375 B.n374 585
R218 B.n373 B.n42 585
R219 B.n372 B.n371 585
R220 B.n370 B.n43 585
R221 B.n369 B.n368 585
R222 B.n367 B.n44 585
R223 B.n366 B.n365 585
R224 B.n364 B.n45 585
R225 B.n363 B.n362 585
R226 B.n361 B.n46 585
R227 B.n360 B.n359 585
R228 B.n358 B.n47 585
R229 B.n357 B.n356 585
R230 B.n355 B.n48 585
R231 B.n354 B.n353 585
R232 B.n352 B.n49 585
R233 B.n351 B.n350 585
R234 B.n349 B.n50 585
R235 B.n348 B.n347 585
R236 B.n439 B.n438 585
R237 B.n440 B.n15 585
R238 B.n442 B.n441 585
R239 B.n443 B.n14 585
R240 B.n445 B.n444 585
R241 B.n446 B.n13 585
R242 B.n448 B.n447 585
R243 B.n449 B.n12 585
R244 B.n451 B.n450 585
R245 B.n452 B.n11 585
R246 B.n454 B.n453 585
R247 B.n455 B.n10 585
R248 B.n457 B.n456 585
R249 B.n458 B.n9 585
R250 B.n460 B.n459 585
R251 B.n461 B.n8 585
R252 B.n463 B.n462 585
R253 B.n464 B.n7 585
R254 B.n466 B.n465 585
R255 B.n467 B.n6 585
R256 B.n469 B.n468 585
R257 B.n470 B.n5 585
R258 B.n472 B.n471 585
R259 B.n473 B.n4 585
R260 B.n475 B.n474 585
R261 B.n476 B.n3 585
R262 B.n478 B.n477 585
R263 B.n479 B.n0 585
R264 B.n2 B.n1 585
R265 B.n126 B.n125 585
R266 B.n128 B.n127 585
R267 B.n129 B.n124 585
R268 B.n131 B.n130 585
R269 B.n132 B.n123 585
R270 B.n134 B.n133 585
R271 B.n135 B.n122 585
R272 B.n137 B.n136 585
R273 B.n138 B.n121 585
R274 B.n140 B.n139 585
R275 B.n141 B.n120 585
R276 B.n143 B.n142 585
R277 B.n144 B.n119 585
R278 B.n146 B.n145 585
R279 B.n147 B.n118 585
R280 B.n149 B.n148 585
R281 B.n150 B.n117 585
R282 B.n152 B.n151 585
R283 B.n153 B.n116 585
R284 B.n155 B.n154 585
R285 B.n156 B.n115 585
R286 B.n158 B.n157 585
R287 B.n159 B.n114 585
R288 B.n161 B.n160 585
R289 B.n162 B.n113 585
R290 B.n164 B.n163 585
R291 B.n165 B.n112 585
R292 B.n167 B.n112 506.916
R293 B.n261 B.n80 506.916
R294 B.n347 B.n346 506.916
R295 B.n438 B.n437 506.916
R296 B.n202 B.t9 283.796
R297 B.n93 B.t0 283.796
R298 B.n37 B.t6 283.796
R299 B.n30 B.t3 283.796
R300 B.n481 B.n480 256.663
R301 B.n480 B.n479 235.042
R302 B.n480 B.n2 235.042
R303 B.n168 B.n167 163.367
R304 B.n169 B.n168 163.367
R305 B.n169 B.n110 163.367
R306 B.n173 B.n110 163.367
R307 B.n174 B.n173 163.367
R308 B.n175 B.n174 163.367
R309 B.n175 B.n108 163.367
R310 B.n179 B.n108 163.367
R311 B.n180 B.n179 163.367
R312 B.n181 B.n180 163.367
R313 B.n181 B.n106 163.367
R314 B.n185 B.n106 163.367
R315 B.n186 B.n185 163.367
R316 B.n187 B.n186 163.367
R317 B.n187 B.n104 163.367
R318 B.n191 B.n104 163.367
R319 B.n192 B.n191 163.367
R320 B.n193 B.n192 163.367
R321 B.n193 B.n102 163.367
R322 B.n197 B.n102 163.367
R323 B.n198 B.n197 163.367
R324 B.n199 B.n198 163.367
R325 B.n199 B.n100 163.367
R326 B.n206 B.n100 163.367
R327 B.n207 B.n206 163.367
R328 B.n208 B.n207 163.367
R329 B.n208 B.n98 163.367
R330 B.n212 B.n98 163.367
R331 B.n213 B.n212 163.367
R332 B.n214 B.n213 163.367
R333 B.n214 B.n96 163.367
R334 B.n218 B.n96 163.367
R335 B.n219 B.n218 163.367
R336 B.n220 B.n219 163.367
R337 B.n220 B.n92 163.367
R338 B.n225 B.n92 163.367
R339 B.n226 B.n225 163.367
R340 B.n227 B.n226 163.367
R341 B.n227 B.n90 163.367
R342 B.n231 B.n90 163.367
R343 B.n232 B.n231 163.367
R344 B.n233 B.n232 163.367
R345 B.n233 B.n88 163.367
R346 B.n237 B.n88 163.367
R347 B.n238 B.n237 163.367
R348 B.n239 B.n238 163.367
R349 B.n239 B.n86 163.367
R350 B.n243 B.n86 163.367
R351 B.n244 B.n243 163.367
R352 B.n245 B.n244 163.367
R353 B.n245 B.n84 163.367
R354 B.n249 B.n84 163.367
R355 B.n250 B.n249 163.367
R356 B.n251 B.n250 163.367
R357 B.n251 B.n82 163.367
R358 B.n255 B.n82 163.367
R359 B.n256 B.n255 163.367
R360 B.n257 B.n256 163.367
R361 B.n257 B.n80 163.367
R362 B.n346 B.n345 163.367
R363 B.n345 B.n52 163.367
R364 B.n341 B.n52 163.367
R365 B.n341 B.n340 163.367
R366 B.n340 B.n339 163.367
R367 B.n339 B.n54 163.367
R368 B.n335 B.n54 163.367
R369 B.n335 B.n334 163.367
R370 B.n334 B.n333 163.367
R371 B.n333 B.n56 163.367
R372 B.n329 B.n56 163.367
R373 B.n329 B.n328 163.367
R374 B.n328 B.n327 163.367
R375 B.n327 B.n58 163.367
R376 B.n323 B.n58 163.367
R377 B.n323 B.n322 163.367
R378 B.n322 B.n321 163.367
R379 B.n321 B.n60 163.367
R380 B.n317 B.n60 163.367
R381 B.n317 B.n316 163.367
R382 B.n316 B.n315 163.367
R383 B.n315 B.n62 163.367
R384 B.n311 B.n62 163.367
R385 B.n311 B.n310 163.367
R386 B.n310 B.n309 163.367
R387 B.n309 B.n64 163.367
R388 B.n305 B.n64 163.367
R389 B.n305 B.n304 163.367
R390 B.n304 B.n303 163.367
R391 B.n303 B.n66 163.367
R392 B.n299 B.n66 163.367
R393 B.n299 B.n298 163.367
R394 B.n298 B.n297 163.367
R395 B.n297 B.n68 163.367
R396 B.n293 B.n68 163.367
R397 B.n293 B.n292 163.367
R398 B.n292 B.n291 163.367
R399 B.n291 B.n70 163.367
R400 B.n287 B.n70 163.367
R401 B.n287 B.n286 163.367
R402 B.n286 B.n285 163.367
R403 B.n285 B.n72 163.367
R404 B.n281 B.n72 163.367
R405 B.n281 B.n280 163.367
R406 B.n280 B.n279 163.367
R407 B.n279 B.n74 163.367
R408 B.n275 B.n74 163.367
R409 B.n275 B.n274 163.367
R410 B.n274 B.n273 163.367
R411 B.n273 B.n76 163.367
R412 B.n269 B.n76 163.367
R413 B.n269 B.n268 163.367
R414 B.n268 B.n267 163.367
R415 B.n267 B.n78 163.367
R416 B.n263 B.n78 163.367
R417 B.n263 B.n262 163.367
R418 B.n262 B.n261 163.367
R419 B.n437 B.n436 163.367
R420 B.n436 B.n17 163.367
R421 B.n432 B.n17 163.367
R422 B.n432 B.n431 163.367
R423 B.n431 B.n430 163.367
R424 B.n430 B.n19 163.367
R425 B.n426 B.n19 163.367
R426 B.n426 B.n425 163.367
R427 B.n425 B.n424 163.367
R428 B.n424 B.n21 163.367
R429 B.n420 B.n21 163.367
R430 B.n420 B.n419 163.367
R431 B.n419 B.n418 163.367
R432 B.n418 B.n23 163.367
R433 B.n414 B.n23 163.367
R434 B.n414 B.n413 163.367
R435 B.n413 B.n412 163.367
R436 B.n412 B.n25 163.367
R437 B.n408 B.n25 163.367
R438 B.n408 B.n407 163.367
R439 B.n407 B.n406 163.367
R440 B.n406 B.n27 163.367
R441 B.n402 B.n27 163.367
R442 B.n402 B.n401 163.367
R443 B.n401 B.n400 163.367
R444 B.n400 B.n29 163.367
R445 B.n396 B.n29 163.367
R446 B.n396 B.n395 163.367
R447 B.n395 B.n394 163.367
R448 B.n394 B.n34 163.367
R449 B.n390 B.n34 163.367
R450 B.n390 B.n389 163.367
R451 B.n389 B.n388 163.367
R452 B.n388 B.n36 163.367
R453 B.n383 B.n36 163.367
R454 B.n383 B.n382 163.367
R455 B.n382 B.n381 163.367
R456 B.n381 B.n40 163.367
R457 B.n377 B.n40 163.367
R458 B.n377 B.n376 163.367
R459 B.n376 B.n375 163.367
R460 B.n375 B.n42 163.367
R461 B.n371 B.n42 163.367
R462 B.n371 B.n370 163.367
R463 B.n370 B.n369 163.367
R464 B.n369 B.n44 163.367
R465 B.n365 B.n44 163.367
R466 B.n365 B.n364 163.367
R467 B.n364 B.n363 163.367
R468 B.n363 B.n46 163.367
R469 B.n359 B.n46 163.367
R470 B.n359 B.n358 163.367
R471 B.n358 B.n357 163.367
R472 B.n357 B.n48 163.367
R473 B.n353 B.n48 163.367
R474 B.n353 B.n352 163.367
R475 B.n352 B.n351 163.367
R476 B.n351 B.n50 163.367
R477 B.n347 B.n50 163.367
R478 B.n438 B.n15 163.367
R479 B.n442 B.n15 163.367
R480 B.n443 B.n442 163.367
R481 B.n444 B.n443 163.367
R482 B.n444 B.n13 163.367
R483 B.n448 B.n13 163.367
R484 B.n449 B.n448 163.367
R485 B.n450 B.n449 163.367
R486 B.n450 B.n11 163.367
R487 B.n454 B.n11 163.367
R488 B.n455 B.n454 163.367
R489 B.n456 B.n455 163.367
R490 B.n456 B.n9 163.367
R491 B.n460 B.n9 163.367
R492 B.n461 B.n460 163.367
R493 B.n462 B.n461 163.367
R494 B.n462 B.n7 163.367
R495 B.n466 B.n7 163.367
R496 B.n467 B.n466 163.367
R497 B.n468 B.n467 163.367
R498 B.n468 B.n5 163.367
R499 B.n472 B.n5 163.367
R500 B.n473 B.n472 163.367
R501 B.n474 B.n473 163.367
R502 B.n474 B.n3 163.367
R503 B.n478 B.n3 163.367
R504 B.n479 B.n478 163.367
R505 B.n126 B.n2 163.367
R506 B.n127 B.n126 163.367
R507 B.n127 B.n124 163.367
R508 B.n131 B.n124 163.367
R509 B.n132 B.n131 163.367
R510 B.n133 B.n132 163.367
R511 B.n133 B.n122 163.367
R512 B.n137 B.n122 163.367
R513 B.n138 B.n137 163.367
R514 B.n139 B.n138 163.367
R515 B.n139 B.n120 163.367
R516 B.n143 B.n120 163.367
R517 B.n144 B.n143 163.367
R518 B.n145 B.n144 163.367
R519 B.n145 B.n118 163.367
R520 B.n149 B.n118 163.367
R521 B.n150 B.n149 163.367
R522 B.n151 B.n150 163.367
R523 B.n151 B.n116 163.367
R524 B.n155 B.n116 163.367
R525 B.n156 B.n155 163.367
R526 B.n157 B.n156 163.367
R527 B.n157 B.n114 163.367
R528 B.n161 B.n114 163.367
R529 B.n162 B.n161 163.367
R530 B.n163 B.n162 163.367
R531 B.n163 B.n112 163.367
R532 B.n93 B.t1 160.786
R533 B.n37 B.t8 160.786
R534 B.n202 B.t10 160.78
R535 B.n30 B.t5 160.78
R536 B.n94 B.t2 115.599
R537 B.n38 B.t7 115.599
R538 B.n203 B.t11 115.593
R539 B.n31 B.t4 115.593
R540 B.n204 B.n203 59.5399
R541 B.n222 B.n94 59.5399
R542 B.n385 B.n38 59.5399
R543 B.n32 B.n31 59.5399
R544 B.n203 B.n202 45.1884
R545 B.n94 B.n93 45.1884
R546 B.n38 B.n37 45.1884
R547 B.n31 B.n30 45.1884
R548 B.n439 B.n16 32.9371
R549 B.n348 B.n51 32.9371
R550 B.n260 B.n259 32.9371
R551 B.n166 B.n165 32.9371
R552 B B.n481 18.0485
R553 B.n440 B.n439 10.6151
R554 B.n441 B.n440 10.6151
R555 B.n441 B.n14 10.6151
R556 B.n445 B.n14 10.6151
R557 B.n446 B.n445 10.6151
R558 B.n447 B.n446 10.6151
R559 B.n447 B.n12 10.6151
R560 B.n451 B.n12 10.6151
R561 B.n452 B.n451 10.6151
R562 B.n453 B.n452 10.6151
R563 B.n453 B.n10 10.6151
R564 B.n457 B.n10 10.6151
R565 B.n458 B.n457 10.6151
R566 B.n459 B.n458 10.6151
R567 B.n459 B.n8 10.6151
R568 B.n463 B.n8 10.6151
R569 B.n464 B.n463 10.6151
R570 B.n465 B.n464 10.6151
R571 B.n465 B.n6 10.6151
R572 B.n469 B.n6 10.6151
R573 B.n470 B.n469 10.6151
R574 B.n471 B.n470 10.6151
R575 B.n471 B.n4 10.6151
R576 B.n475 B.n4 10.6151
R577 B.n476 B.n475 10.6151
R578 B.n477 B.n476 10.6151
R579 B.n477 B.n0 10.6151
R580 B.n435 B.n16 10.6151
R581 B.n435 B.n434 10.6151
R582 B.n434 B.n433 10.6151
R583 B.n433 B.n18 10.6151
R584 B.n429 B.n18 10.6151
R585 B.n429 B.n428 10.6151
R586 B.n428 B.n427 10.6151
R587 B.n427 B.n20 10.6151
R588 B.n423 B.n20 10.6151
R589 B.n423 B.n422 10.6151
R590 B.n422 B.n421 10.6151
R591 B.n421 B.n22 10.6151
R592 B.n417 B.n22 10.6151
R593 B.n417 B.n416 10.6151
R594 B.n416 B.n415 10.6151
R595 B.n415 B.n24 10.6151
R596 B.n411 B.n24 10.6151
R597 B.n411 B.n410 10.6151
R598 B.n410 B.n409 10.6151
R599 B.n409 B.n26 10.6151
R600 B.n405 B.n26 10.6151
R601 B.n405 B.n404 10.6151
R602 B.n404 B.n403 10.6151
R603 B.n403 B.n28 10.6151
R604 B.n399 B.n398 10.6151
R605 B.n398 B.n397 10.6151
R606 B.n397 B.n33 10.6151
R607 B.n393 B.n33 10.6151
R608 B.n393 B.n392 10.6151
R609 B.n392 B.n391 10.6151
R610 B.n391 B.n35 10.6151
R611 B.n387 B.n35 10.6151
R612 B.n387 B.n386 10.6151
R613 B.n384 B.n39 10.6151
R614 B.n380 B.n39 10.6151
R615 B.n380 B.n379 10.6151
R616 B.n379 B.n378 10.6151
R617 B.n378 B.n41 10.6151
R618 B.n374 B.n41 10.6151
R619 B.n374 B.n373 10.6151
R620 B.n373 B.n372 10.6151
R621 B.n372 B.n43 10.6151
R622 B.n368 B.n43 10.6151
R623 B.n368 B.n367 10.6151
R624 B.n367 B.n366 10.6151
R625 B.n366 B.n45 10.6151
R626 B.n362 B.n45 10.6151
R627 B.n362 B.n361 10.6151
R628 B.n361 B.n360 10.6151
R629 B.n360 B.n47 10.6151
R630 B.n356 B.n47 10.6151
R631 B.n356 B.n355 10.6151
R632 B.n355 B.n354 10.6151
R633 B.n354 B.n49 10.6151
R634 B.n350 B.n49 10.6151
R635 B.n350 B.n349 10.6151
R636 B.n349 B.n348 10.6151
R637 B.n344 B.n51 10.6151
R638 B.n344 B.n343 10.6151
R639 B.n343 B.n342 10.6151
R640 B.n342 B.n53 10.6151
R641 B.n338 B.n53 10.6151
R642 B.n338 B.n337 10.6151
R643 B.n337 B.n336 10.6151
R644 B.n336 B.n55 10.6151
R645 B.n332 B.n55 10.6151
R646 B.n332 B.n331 10.6151
R647 B.n331 B.n330 10.6151
R648 B.n330 B.n57 10.6151
R649 B.n326 B.n57 10.6151
R650 B.n326 B.n325 10.6151
R651 B.n325 B.n324 10.6151
R652 B.n324 B.n59 10.6151
R653 B.n320 B.n59 10.6151
R654 B.n320 B.n319 10.6151
R655 B.n319 B.n318 10.6151
R656 B.n318 B.n61 10.6151
R657 B.n314 B.n61 10.6151
R658 B.n314 B.n313 10.6151
R659 B.n313 B.n312 10.6151
R660 B.n312 B.n63 10.6151
R661 B.n308 B.n63 10.6151
R662 B.n308 B.n307 10.6151
R663 B.n307 B.n306 10.6151
R664 B.n306 B.n65 10.6151
R665 B.n302 B.n65 10.6151
R666 B.n302 B.n301 10.6151
R667 B.n301 B.n300 10.6151
R668 B.n300 B.n67 10.6151
R669 B.n296 B.n67 10.6151
R670 B.n296 B.n295 10.6151
R671 B.n295 B.n294 10.6151
R672 B.n294 B.n69 10.6151
R673 B.n290 B.n69 10.6151
R674 B.n290 B.n289 10.6151
R675 B.n289 B.n288 10.6151
R676 B.n288 B.n71 10.6151
R677 B.n284 B.n71 10.6151
R678 B.n284 B.n283 10.6151
R679 B.n283 B.n282 10.6151
R680 B.n282 B.n73 10.6151
R681 B.n278 B.n73 10.6151
R682 B.n278 B.n277 10.6151
R683 B.n277 B.n276 10.6151
R684 B.n276 B.n75 10.6151
R685 B.n272 B.n75 10.6151
R686 B.n272 B.n271 10.6151
R687 B.n271 B.n270 10.6151
R688 B.n270 B.n77 10.6151
R689 B.n266 B.n77 10.6151
R690 B.n266 B.n265 10.6151
R691 B.n265 B.n264 10.6151
R692 B.n264 B.n79 10.6151
R693 B.n260 B.n79 10.6151
R694 B.n125 B.n1 10.6151
R695 B.n128 B.n125 10.6151
R696 B.n129 B.n128 10.6151
R697 B.n130 B.n129 10.6151
R698 B.n130 B.n123 10.6151
R699 B.n134 B.n123 10.6151
R700 B.n135 B.n134 10.6151
R701 B.n136 B.n135 10.6151
R702 B.n136 B.n121 10.6151
R703 B.n140 B.n121 10.6151
R704 B.n141 B.n140 10.6151
R705 B.n142 B.n141 10.6151
R706 B.n142 B.n119 10.6151
R707 B.n146 B.n119 10.6151
R708 B.n147 B.n146 10.6151
R709 B.n148 B.n147 10.6151
R710 B.n148 B.n117 10.6151
R711 B.n152 B.n117 10.6151
R712 B.n153 B.n152 10.6151
R713 B.n154 B.n153 10.6151
R714 B.n154 B.n115 10.6151
R715 B.n158 B.n115 10.6151
R716 B.n159 B.n158 10.6151
R717 B.n160 B.n159 10.6151
R718 B.n160 B.n113 10.6151
R719 B.n164 B.n113 10.6151
R720 B.n165 B.n164 10.6151
R721 B.n166 B.n111 10.6151
R722 B.n170 B.n111 10.6151
R723 B.n171 B.n170 10.6151
R724 B.n172 B.n171 10.6151
R725 B.n172 B.n109 10.6151
R726 B.n176 B.n109 10.6151
R727 B.n177 B.n176 10.6151
R728 B.n178 B.n177 10.6151
R729 B.n178 B.n107 10.6151
R730 B.n182 B.n107 10.6151
R731 B.n183 B.n182 10.6151
R732 B.n184 B.n183 10.6151
R733 B.n184 B.n105 10.6151
R734 B.n188 B.n105 10.6151
R735 B.n189 B.n188 10.6151
R736 B.n190 B.n189 10.6151
R737 B.n190 B.n103 10.6151
R738 B.n194 B.n103 10.6151
R739 B.n195 B.n194 10.6151
R740 B.n196 B.n195 10.6151
R741 B.n196 B.n101 10.6151
R742 B.n200 B.n101 10.6151
R743 B.n201 B.n200 10.6151
R744 B.n205 B.n201 10.6151
R745 B.n209 B.n99 10.6151
R746 B.n210 B.n209 10.6151
R747 B.n211 B.n210 10.6151
R748 B.n211 B.n97 10.6151
R749 B.n215 B.n97 10.6151
R750 B.n216 B.n215 10.6151
R751 B.n217 B.n216 10.6151
R752 B.n217 B.n95 10.6151
R753 B.n221 B.n95 10.6151
R754 B.n224 B.n223 10.6151
R755 B.n224 B.n91 10.6151
R756 B.n228 B.n91 10.6151
R757 B.n229 B.n228 10.6151
R758 B.n230 B.n229 10.6151
R759 B.n230 B.n89 10.6151
R760 B.n234 B.n89 10.6151
R761 B.n235 B.n234 10.6151
R762 B.n236 B.n235 10.6151
R763 B.n236 B.n87 10.6151
R764 B.n240 B.n87 10.6151
R765 B.n241 B.n240 10.6151
R766 B.n242 B.n241 10.6151
R767 B.n242 B.n85 10.6151
R768 B.n246 B.n85 10.6151
R769 B.n247 B.n246 10.6151
R770 B.n248 B.n247 10.6151
R771 B.n248 B.n83 10.6151
R772 B.n252 B.n83 10.6151
R773 B.n253 B.n252 10.6151
R774 B.n254 B.n253 10.6151
R775 B.n254 B.n81 10.6151
R776 B.n258 B.n81 10.6151
R777 B.n259 B.n258 10.6151
R778 B.n32 B.n28 9.36635
R779 B.n385 B.n384 9.36635
R780 B.n205 B.n204 9.36635
R781 B.n223 B.n222 9.36635
R782 B.n481 B.n0 8.11757
R783 B.n481 B.n1 8.11757
R784 B.n399 B.n32 1.24928
R785 B.n386 B.n385 1.24928
R786 B.n204 B.n99 1.24928
R787 B.n222 B.n221 1.24928
C0 VN B 0.929736f
C1 VTAIL w_n2368_n2244# 2.67683f
C2 VDD2 w_n2368_n2244# 1.23024f
C3 VTAIL VP 2.71205f
C4 VDD2 VP 0.356585f
C5 VTAIL VN 2.69794f
C6 VDD2 VN 2.53907f
C7 VDD1 w_n2368_n2244# 1.18754f
C8 VDD1 VP 2.74615f
C9 VDD1 VN 0.148917f
C10 VP w_n2368_n2244# 4.09519f
C11 VN w_n2368_n2244# 3.79229f
C12 VN VP 4.71561f
C13 VTAIL B 2.88016f
C14 VDD2 B 1.04798f
C15 VTAIL VDD2 3.94441f
C16 VDD1 B 1.00566f
C17 B w_n2368_n2244# 6.93783f
C18 VTAIL VDD1 3.89422f
C19 VDD2 VDD1 0.88379f
C20 VP B 1.42959f
C21 VDD2 VSUBS 0.707636f
C22 VDD1 VSUBS 4.61273f
C23 VTAIL VSUBS 0.67193f
C24 VN VSUBS 4.98799f
C25 VP VSUBS 1.671241f
C26 B VSUBS 3.280509f
C27 w_n2368_n2244# VSUBS 66.23771f
C28 B.n0 VSUBS 0.007383f
C29 B.n1 VSUBS 0.007383f
C30 B.n2 VSUBS 0.010919f
C31 B.n3 VSUBS 0.008367f
C32 B.n4 VSUBS 0.008367f
C33 B.n5 VSUBS 0.008367f
C34 B.n6 VSUBS 0.008367f
C35 B.n7 VSUBS 0.008367f
C36 B.n8 VSUBS 0.008367f
C37 B.n9 VSUBS 0.008367f
C38 B.n10 VSUBS 0.008367f
C39 B.n11 VSUBS 0.008367f
C40 B.n12 VSUBS 0.008367f
C41 B.n13 VSUBS 0.008367f
C42 B.n14 VSUBS 0.008367f
C43 B.n15 VSUBS 0.008367f
C44 B.n16 VSUBS 0.020393f
C45 B.n17 VSUBS 0.008367f
C46 B.n18 VSUBS 0.008367f
C47 B.n19 VSUBS 0.008367f
C48 B.n20 VSUBS 0.008367f
C49 B.n21 VSUBS 0.008367f
C50 B.n22 VSUBS 0.008367f
C51 B.n23 VSUBS 0.008367f
C52 B.n24 VSUBS 0.008367f
C53 B.n25 VSUBS 0.008367f
C54 B.n26 VSUBS 0.008367f
C55 B.n27 VSUBS 0.008367f
C56 B.n28 VSUBS 0.007875f
C57 B.n29 VSUBS 0.008367f
C58 B.t4 VSUBS 0.225399f
C59 B.t5 VSUBS 0.245097f
C60 B.t3 VSUBS 0.709023f
C61 B.n30 VSUBS 0.136882f
C62 B.n31 VSUBS 0.082019f
C63 B.n32 VSUBS 0.019386f
C64 B.n33 VSUBS 0.008367f
C65 B.n34 VSUBS 0.008367f
C66 B.n35 VSUBS 0.008367f
C67 B.n36 VSUBS 0.008367f
C68 B.t7 VSUBS 0.225398f
C69 B.t8 VSUBS 0.245095f
C70 B.t6 VSUBS 0.709023f
C71 B.n37 VSUBS 0.136883f
C72 B.n38 VSUBS 0.08202f
C73 B.n39 VSUBS 0.008367f
C74 B.n40 VSUBS 0.008367f
C75 B.n41 VSUBS 0.008367f
C76 B.n42 VSUBS 0.008367f
C77 B.n43 VSUBS 0.008367f
C78 B.n44 VSUBS 0.008367f
C79 B.n45 VSUBS 0.008367f
C80 B.n46 VSUBS 0.008367f
C81 B.n47 VSUBS 0.008367f
C82 B.n48 VSUBS 0.008367f
C83 B.n49 VSUBS 0.008367f
C84 B.n50 VSUBS 0.008367f
C85 B.n51 VSUBS 0.018982f
C86 B.n52 VSUBS 0.008367f
C87 B.n53 VSUBS 0.008367f
C88 B.n54 VSUBS 0.008367f
C89 B.n55 VSUBS 0.008367f
C90 B.n56 VSUBS 0.008367f
C91 B.n57 VSUBS 0.008367f
C92 B.n58 VSUBS 0.008367f
C93 B.n59 VSUBS 0.008367f
C94 B.n60 VSUBS 0.008367f
C95 B.n61 VSUBS 0.008367f
C96 B.n62 VSUBS 0.008367f
C97 B.n63 VSUBS 0.008367f
C98 B.n64 VSUBS 0.008367f
C99 B.n65 VSUBS 0.008367f
C100 B.n66 VSUBS 0.008367f
C101 B.n67 VSUBS 0.008367f
C102 B.n68 VSUBS 0.008367f
C103 B.n69 VSUBS 0.008367f
C104 B.n70 VSUBS 0.008367f
C105 B.n71 VSUBS 0.008367f
C106 B.n72 VSUBS 0.008367f
C107 B.n73 VSUBS 0.008367f
C108 B.n74 VSUBS 0.008367f
C109 B.n75 VSUBS 0.008367f
C110 B.n76 VSUBS 0.008367f
C111 B.n77 VSUBS 0.008367f
C112 B.n78 VSUBS 0.008367f
C113 B.n79 VSUBS 0.008367f
C114 B.n80 VSUBS 0.020393f
C115 B.n81 VSUBS 0.008367f
C116 B.n82 VSUBS 0.008367f
C117 B.n83 VSUBS 0.008367f
C118 B.n84 VSUBS 0.008367f
C119 B.n85 VSUBS 0.008367f
C120 B.n86 VSUBS 0.008367f
C121 B.n87 VSUBS 0.008367f
C122 B.n88 VSUBS 0.008367f
C123 B.n89 VSUBS 0.008367f
C124 B.n90 VSUBS 0.008367f
C125 B.n91 VSUBS 0.008367f
C126 B.n92 VSUBS 0.008367f
C127 B.t2 VSUBS 0.225398f
C128 B.t1 VSUBS 0.245095f
C129 B.t0 VSUBS 0.709023f
C130 B.n93 VSUBS 0.136883f
C131 B.n94 VSUBS 0.08202f
C132 B.n95 VSUBS 0.008367f
C133 B.n96 VSUBS 0.008367f
C134 B.n97 VSUBS 0.008367f
C135 B.n98 VSUBS 0.008367f
C136 B.n99 VSUBS 0.004676f
C137 B.n100 VSUBS 0.008367f
C138 B.n101 VSUBS 0.008367f
C139 B.n102 VSUBS 0.008367f
C140 B.n103 VSUBS 0.008367f
C141 B.n104 VSUBS 0.008367f
C142 B.n105 VSUBS 0.008367f
C143 B.n106 VSUBS 0.008367f
C144 B.n107 VSUBS 0.008367f
C145 B.n108 VSUBS 0.008367f
C146 B.n109 VSUBS 0.008367f
C147 B.n110 VSUBS 0.008367f
C148 B.n111 VSUBS 0.008367f
C149 B.n112 VSUBS 0.018982f
C150 B.n113 VSUBS 0.008367f
C151 B.n114 VSUBS 0.008367f
C152 B.n115 VSUBS 0.008367f
C153 B.n116 VSUBS 0.008367f
C154 B.n117 VSUBS 0.008367f
C155 B.n118 VSUBS 0.008367f
C156 B.n119 VSUBS 0.008367f
C157 B.n120 VSUBS 0.008367f
C158 B.n121 VSUBS 0.008367f
C159 B.n122 VSUBS 0.008367f
C160 B.n123 VSUBS 0.008367f
C161 B.n124 VSUBS 0.008367f
C162 B.n125 VSUBS 0.008367f
C163 B.n126 VSUBS 0.008367f
C164 B.n127 VSUBS 0.008367f
C165 B.n128 VSUBS 0.008367f
C166 B.n129 VSUBS 0.008367f
C167 B.n130 VSUBS 0.008367f
C168 B.n131 VSUBS 0.008367f
C169 B.n132 VSUBS 0.008367f
C170 B.n133 VSUBS 0.008367f
C171 B.n134 VSUBS 0.008367f
C172 B.n135 VSUBS 0.008367f
C173 B.n136 VSUBS 0.008367f
C174 B.n137 VSUBS 0.008367f
C175 B.n138 VSUBS 0.008367f
C176 B.n139 VSUBS 0.008367f
C177 B.n140 VSUBS 0.008367f
C178 B.n141 VSUBS 0.008367f
C179 B.n142 VSUBS 0.008367f
C180 B.n143 VSUBS 0.008367f
C181 B.n144 VSUBS 0.008367f
C182 B.n145 VSUBS 0.008367f
C183 B.n146 VSUBS 0.008367f
C184 B.n147 VSUBS 0.008367f
C185 B.n148 VSUBS 0.008367f
C186 B.n149 VSUBS 0.008367f
C187 B.n150 VSUBS 0.008367f
C188 B.n151 VSUBS 0.008367f
C189 B.n152 VSUBS 0.008367f
C190 B.n153 VSUBS 0.008367f
C191 B.n154 VSUBS 0.008367f
C192 B.n155 VSUBS 0.008367f
C193 B.n156 VSUBS 0.008367f
C194 B.n157 VSUBS 0.008367f
C195 B.n158 VSUBS 0.008367f
C196 B.n159 VSUBS 0.008367f
C197 B.n160 VSUBS 0.008367f
C198 B.n161 VSUBS 0.008367f
C199 B.n162 VSUBS 0.008367f
C200 B.n163 VSUBS 0.008367f
C201 B.n164 VSUBS 0.008367f
C202 B.n165 VSUBS 0.018982f
C203 B.n166 VSUBS 0.020393f
C204 B.n167 VSUBS 0.020393f
C205 B.n168 VSUBS 0.008367f
C206 B.n169 VSUBS 0.008367f
C207 B.n170 VSUBS 0.008367f
C208 B.n171 VSUBS 0.008367f
C209 B.n172 VSUBS 0.008367f
C210 B.n173 VSUBS 0.008367f
C211 B.n174 VSUBS 0.008367f
C212 B.n175 VSUBS 0.008367f
C213 B.n176 VSUBS 0.008367f
C214 B.n177 VSUBS 0.008367f
C215 B.n178 VSUBS 0.008367f
C216 B.n179 VSUBS 0.008367f
C217 B.n180 VSUBS 0.008367f
C218 B.n181 VSUBS 0.008367f
C219 B.n182 VSUBS 0.008367f
C220 B.n183 VSUBS 0.008367f
C221 B.n184 VSUBS 0.008367f
C222 B.n185 VSUBS 0.008367f
C223 B.n186 VSUBS 0.008367f
C224 B.n187 VSUBS 0.008367f
C225 B.n188 VSUBS 0.008367f
C226 B.n189 VSUBS 0.008367f
C227 B.n190 VSUBS 0.008367f
C228 B.n191 VSUBS 0.008367f
C229 B.n192 VSUBS 0.008367f
C230 B.n193 VSUBS 0.008367f
C231 B.n194 VSUBS 0.008367f
C232 B.n195 VSUBS 0.008367f
C233 B.n196 VSUBS 0.008367f
C234 B.n197 VSUBS 0.008367f
C235 B.n198 VSUBS 0.008367f
C236 B.n199 VSUBS 0.008367f
C237 B.n200 VSUBS 0.008367f
C238 B.n201 VSUBS 0.008367f
C239 B.t11 VSUBS 0.225399f
C240 B.t10 VSUBS 0.245097f
C241 B.t9 VSUBS 0.709023f
C242 B.n202 VSUBS 0.136882f
C243 B.n203 VSUBS 0.082019f
C244 B.n204 VSUBS 0.019386f
C245 B.n205 VSUBS 0.007875f
C246 B.n206 VSUBS 0.008367f
C247 B.n207 VSUBS 0.008367f
C248 B.n208 VSUBS 0.008367f
C249 B.n209 VSUBS 0.008367f
C250 B.n210 VSUBS 0.008367f
C251 B.n211 VSUBS 0.008367f
C252 B.n212 VSUBS 0.008367f
C253 B.n213 VSUBS 0.008367f
C254 B.n214 VSUBS 0.008367f
C255 B.n215 VSUBS 0.008367f
C256 B.n216 VSUBS 0.008367f
C257 B.n217 VSUBS 0.008367f
C258 B.n218 VSUBS 0.008367f
C259 B.n219 VSUBS 0.008367f
C260 B.n220 VSUBS 0.008367f
C261 B.n221 VSUBS 0.004676f
C262 B.n222 VSUBS 0.019386f
C263 B.n223 VSUBS 0.007875f
C264 B.n224 VSUBS 0.008367f
C265 B.n225 VSUBS 0.008367f
C266 B.n226 VSUBS 0.008367f
C267 B.n227 VSUBS 0.008367f
C268 B.n228 VSUBS 0.008367f
C269 B.n229 VSUBS 0.008367f
C270 B.n230 VSUBS 0.008367f
C271 B.n231 VSUBS 0.008367f
C272 B.n232 VSUBS 0.008367f
C273 B.n233 VSUBS 0.008367f
C274 B.n234 VSUBS 0.008367f
C275 B.n235 VSUBS 0.008367f
C276 B.n236 VSUBS 0.008367f
C277 B.n237 VSUBS 0.008367f
C278 B.n238 VSUBS 0.008367f
C279 B.n239 VSUBS 0.008367f
C280 B.n240 VSUBS 0.008367f
C281 B.n241 VSUBS 0.008367f
C282 B.n242 VSUBS 0.008367f
C283 B.n243 VSUBS 0.008367f
C284 B.n244 VSUBS 0.008367f
C285 B.n245 VSUBS 0.008367f
C286 B.n246 VSUBS 0.008367f
C287 B.n247 VSUBS 0.008367f
C288 B.n248 VSUBS 0.008367f
C289 B.n249 VSUBS 0.008367f
C290 B.n250 VSUBS 0.008367f
C291 B.n251 VSUBS 0.008367f
C292 B.n252 VSUBS 0.008367f
C293 B.n253 VSUBS 0.008367f
C294 B.n254 VSUBS 0.008367f
C295 B.n255 VSUBS 0.008367f
C296 B.n256 VSUBS 0.008367f
C297 B.n257 VSUBS 0.008367f
C298 B.n258 VSUBS 0.008367f
C299 B.n259 VSUBS 0.019413f
C300 B.n260 VSUBS 0.019963f
C301 B.n261 VSUBS 0.018982f
C302 B.n262 VSUBS 0.008367f
C303 B.n263 VSUBS 0.008367f
C304 B.n264 VSUBS 0.008367f
C305 B.n265 VSUBS 0.008367f
C306 B.n266 VSUBS 0.008367f
C307 B.n267 VSUBS 0.008367f
C308 B.n268 VSUBS 0.008367f
C309 B.n269 VSUBS 0.008367f
C310 B.n270 VSUBS 0.008367f
C311 B.n271 VSUBS 0.008367f
C312 B.n272 VSUBS 0.008367f
C313 B.n273 VSUBS 0.008367f
C314 B.n274 VSUBS 0.008367f
C315 B.n275 VSUBS 0.008367f
C316 B.n276 VSUBS 0.008367f
C317 B.n277 VSUBS 0.008367f
C318 B.n278 VSUBS 0.008367f
C319 B.n279 VSUBS 0.008367f
C320 B.n280 VSUBS 0.008367f
C321 B.n281 VSUBS 0.008367f
C322 B.n282 VSUBS 0.008367f
C323 B.n283 VSUBS 0.008367f
C324 B.n284 VSUBS 0.008367f
C325 B.n285 VSUBS 0.008367f
C326 B.n286 VSUBS 0.008367f
C327 B.n287 VSUBS 0.008367f
C328 B.n288 VSUBS 0.008367f
C329 B.n289 VSUBS 0.008367f
C330 B.n290 VSUBS 0.008367f
C331 B.n291 VSUBS 0.008367f
C332 B.n292 VSUBS 0.008367f
C333 B.n293 VSUBS 0.008367f
C334 B.n294 VSUBS 0.008367f
C335 B.n295 VSUBS 0.008367f
C336 B.n296 VSUBS 0.008367f
C337 B.n297 VSUBS 0.008367f
C338 B.n298 VSUBS 0.008367f
C339 B.n299 VSUBS 0.008367f
C340 B.n300 VSUBS 0.008367f
C341 B.n301 VSUBS 0.008367f
C342 B.n302 VSUBS 0.008367f
C343 B.n303 VSUBS 0.008367f
C344 B.n304 VSUBS 0.008367f
C345 B.n305 VSUBS 0.008367f
C346 B.n306 VSUBS 0.008367f
C347 B.n307 VSUBS 0.008367f
C348 B.n308 VSUBS 0.008367f
C349 B.n309 VSUBS 0.008367f
C350 B.n310 VSUBS 0.008367f
C351 B.n311 VSUBS 0.008367f
C352 B.n312 VSUBS 0.008367f
C353 B.n313 VSUBS 0.008367f
C354 B.n314 VSUBS 0.008367f
C355 B.n315 VSUBS 0.008367f
C356 B.n316 VSUBS 0.008367f
C357 B.n317 VSUBS 0.008367f
C358 B.n318 VSUBS 0.008367f
C359 B.n319 VSUBS 0.008367f
C360 B.n320 VSUBS 0.008367f
C361 B.n321 VSUBS 0.008367f
C362 B.n322 VSUBS 0.008367f
C363 B.n323 VSUBS 0.008367f
C364 B.n324 VSUBS 0.008367f
C365 B.n325 VSUBS 0.008367f
C366 B.n326 VSUBS 0.008367f
C367 B.n327 VSUBS 0.008367f
C368 B.n328 VSUBS 0.008367f
C369 B.n329 VSUBS 0.008367f
C370 B.n330 VSUBS 0.008367f
C371 B.n331 VSUBS 0.008367f
C372 B.n332 VSUBS 0.008367f
C373 B.n333 VSUBS 0.008367f
C374 B.n334 VSUBS 0.008367f
C375 B.n335 VSUBS 0.008367f
C376 B.n336 VSUBS 0.008367f
C377 B.n337 VSUBS 0.008367f
C378 B.n338 VSUBS 0.008367f
C379 B.n339 VSUBS 0.008367f
C380 B.n340 VSUBS 0.008367f
C381 B.n341 VSUBS 0.008367f
C382 B.n342 VSUBS 0.008367f
C383 B.n343 VSUBS 0.008367f
C384 B.n344 VSUBS 0.008367f
C385 B.n345 VSUBS 0.008367f
C386 B.n346 VSUBS 0.018982f
C387 B.n347 VSUBS 0.020393f
C388 B.n348 VSUBS 0.020393f
C389 B.n349 VSUBS 0.008367f
C390 B.n350 VSUBS 0.008367f
C391 B.n351 VSUBS 0.008367f
C392 B.n352 VSUBS 0.008367f
C393 B.n353 VSUBS 0.008367f
C394 B.n354 VSUBS 0.008367f
C395 B.n355 VSUBS 0.008367f
C396 B.n356 VSUBS 0.008367f
C397 B.n357 VSUBS 0.008367f
C398 B.n358 VSUBS 0.008367f
C399 B.n359 VSUBS 0.008367f
C400 B.n360 VSUBS 0.008367f
C401 B.n361 VSUBS 0.008367f
C402 B.n362 VSUBS 0.008367f
C403 B.n363 VSUBS 0.008367f
C404 B.n364 VSUBS 0.008367f
C405 B.n365 VSUBS 0.008367f
C406 B.n366 VSUBS 0.008367f
C407 B.n367 VSUBS 0.008367f
C408 B.n368 VSUBS 0.008367f
C409 B.n369 VSUBS 0.008367f
C410 B.n370 VSUBS 0.008367f
C411 B.n371 VSUBS 0.008367f
C412 B.n372 VSUBS 0.008367f
C413 B.n373 VSUBS 0.008367f
C414 B.n374 VSUBS 0.008367f
C415 B.n375 VSUBS 0.008367f
C416 B.n376 VSUBS 0.008367f
C417 B.n377 VSUBS 0.008367f
C418 B.n378 VSUBS 0.008367f
C419 B.n379 VSUBS 0.008367f
C420 B.n380 VSUBS 0.008367f
C421 B.n381 VSUBS 0.008367f
C422 B.n382 VSUBS 0.008367f
C423 B.n383 VSUBS 0.008367f
C424 B.n384 VSUBS 0.007875f
C425 B.n385 VSUBS 0.019386f
C426 B.n386 VSUBS 0.004676f
C427 B.n387 VSUBS 0.008367f
C428 B.n388 VSUBS 0.008367f
C429 B.n389 VSUBS 0.008367f
C430 B.n390 VSUBS 0.008367f
C431 B.n391 VSUBS 0.008367f
C432 B.n392 VSUBS 0.008367f
C433 B.n393 VSUBS 0.008367f
C434 B.n394 VSUBS 0.008367f
C435 B.n395 VSUBS 0.008367f
C436 B.n396 VSUBS 0.008367f
C437 B.n397 VSUBS 0.008367f
C438 B.n398 VSUBS 0.008367f
C439 B.n399 VSUBS 0.004676f
C440 B.n400 VSUBS 0.008367f
C441 B.n401 VSUBS 0.008367f
C442 B.n402 VSUBS 0.008367f
C443 B.n403 VSUBS 0.008367f
C444 B.n404 VSUBS 0.008367f
C445 B.n405 VSUBS 0.008367f
C446 B.n406 VSUBS 0.008367f
C447 B.n407 VSUBS 0.008367f
C448 B.n408 VSUBS 0.008367f
C449 B.n409 VSUBS 0.008367f
C450 B.n410 VSUBS 0.008367f
C451 B.n411 VSUBS 0.008367f
C452 B.n412 VSUBS 0.008367f
C453 B.n413 VSUBS 0.008367f
C454 B.n414 VSUBS 0.008367f
C455 B.n415 VSUBS 0.008367f
C456 B.n416 VSUBS 0.008367f
C457 B.n417 VSUBS 0.008367f
C458 B.n418 VSUBS 0.008367f
C459 B.n419 VSUBS 0.008367f
C460 B.n420 VSUBS 0.008367f
C461 B.n421 VSUBS 0.008367f
C462 B.n422 VSUBS 0.008367f
C463 B.n423 VSUBS 0.008367f
C464 B.n424 VSUBS 0.008367f
C465 B.n425 VSUBS 0.008367f
C466 B.n426 VSUBS 0.008367f
C467 B.n427 VSUBS 0.008367f
C468 B.n428 VSUBS 0.008367f
C469 B.n429 VSUBS 0.008367f
C470 B.n430 VSUBS 0.008367f
C471 B.n431 VSUBS 0.008367f
C472 B.n432 VSUBS 0.008367f
C473 B.n433 VSUBS 0.008367f
C474 B.n434 VSUBS 0.008367f
C475 B.n435 VSUBS 0.008367f
C476 B.n436 VSUBS 0.008367f
C477 B.n437 VSUBS 0.020393f
C478 B.n438 VSUBS 0.018982f
C479 B.n439 VSUBS 0.018982f
C480 B.n440 VSUBS 0.008367f
C481 B.n441 VSUBS 0.008367f
C482 B.n442 VSUBS 0.008367f
C483 B.n443 VSUBS 0.008367f
C484 B.n444 VSUBS 0.008367f
C485 B.n445 VSUBS 0.008367f
C486 B.n446 VSUBS 0.008367f
C487 B.n447 VSUBS 0.008367f
C488 B.n448 VSUBS 0.008367f
C489 B.n449 VSUBS 0.008367f
C490 B.n450 VSUBS 0.008367f
C491 B.n451 VSUBS 0.008367f
C492 B.n452 VSUBS 0.008367f
C493 B.n453 VSUBS 0.008367f
C494 B.n454 VSUBS 0.008367f
C495 B.n455 VSUBS 0.008367f
C496 B.n456 VSUBS 0.008367f
C497 B.n457 VSUBS 0.008367f
C498 B.n458 VSUBS 0.008367f
C499 B.n459 VSUBS 0.008367f
C500 B.n460 VSUBS 0.008367f
C501 B.n461 VSUBS 0.008367f
C502 B.n462 VSUBS 0.008367f
C503 B.n463 VSUBS 0.008367f
C504 B.n464 VSUBS 0.008367f
C505 B.n465 VSUBS 0.008367f
C506 B.n466 VSUBS 0.008367f
C507 B.n467 VSUBS 0.008367f
C508 B.n468 VSUBS 0.008367f
C509 B.n469 VSUBS 0.008367f
C510 B.n470 VSUBS 0.008367f
C511 B.n471 VSUBS 0.008367f
C512 B.n472 VSUBS 0.008367f
C513 B.n473 VSUBS 0.008367f
C514 B.n474 VSUBS 0.008367f
C515 B.n475 VSUBS 0.008367f
C516 B.n476 VSUBS 0.008367f
C517 B.n477 VSUBS 0.008367f
C518 B.n478 VSUBS 0.008367f
C519 B.n479 VSUBS 0.010919f
C520 B.n480 VSUBS 0.011631f
C521 B.n481 VSUBS 0.02313f
C522 VDD1.t3 VSUBS 0.137298f
C523 VDD1.t1 VSUBS 0.137298f
C524 VDD1.n0 VSUBS 0.925901f
C525 VDD1.t0 VSUBS 0.137298f
C526 VDD1.t2 VSUBS 0.137298f
C527 VDD1.n1 VSUBS 1.36832f
C528 VP.n0 VSUBS 0.061286f
C529 VP.t1 VSUBS 1.57553f
C530 VP.n1 VSUBS 0.067577f
C531 VP.t2 VSUBS 1.83816f
C532 VP.t0 VSUBS 1.84214f
C533 VP.n2 VSUBS 3.07772f
C534 VP.n3 VSUBS 2.19295f
C535 VP.t3 VSUBS 1.57553f
C536 VP.n4 VSUBS 0.739815f
C537 VP.n5 VSUBS 0.078973f
C538 VP.n6 VSUBS 0.061286f
C539 VP.n7 VSUBS 0.046488f
C540 VP.n8 VSUBS 0.046488f
C541 VP.n9 VSUBS 0.067577f
C542 VP.n10 VSUBS 0.078973f
C543 VP.n11 VSUBS 0.739815f
C544 VP.n12 VSUBS 0.055718f
C545 VTAIL.t6 VSUBS 1.09635f
C546 VTAIL.n0 VSUBS 0.694541f
C547 VTAIL.t0 VSUBS 1.09635f
C548 VTAIL.n1 VSUBS 0.775014f
C549 VTAIL.t3 VSUBS 1.09635f
C550 VTAIL.n2 VSUBS 1.73228f
C551 VTAIL.t7 VSUBS 1.09636f
C552 VTAIL.n3 VSUBS 1.73227f
C553 VTAIL.t5 VSUBS 1.09636f
C554 VTAIL.n4 VSUBS 0.775008f
C555 VTAIL.t2 VSUBS 1.09636f
C556 VTAIL.n5 VSUBS 0.775008f
C557 VTAIL.t1 VSUBS 1.09635f
C558 VTAIL.n6 VSUBS 1.73228f
C559 VTAIL.t4 VSUBS 1.09635f
C560 VTAIL.n7 VSUBS 1.64191f
C561 VDD2.t0 VSUBS 0.135198f
C562 VDD2.t1 VSUBS 0.135198f
C563 VDD2.n0 VSUBS 1.32758f
C564 VDD2.t2 VSUBS 0.135198f
C565 VDD2.t3 VSUBS 0.135198f
C566 VDD2.n1 VSUBS 0.911332f
C567 VDD2.n2 VSUBS 3.44096f
C568 VN.t1 VSUBS 1.76913f
C569 VN.t3 VSUBS 1.76531f
C570 VN.n0 VSUBS 1.21248f
C571 VN.t2 VSUBS 1.76913f
C572 VN.t0 VSUBS 1.76531f
C573 VN.n1 VSUBS 2.97875f
.ends

