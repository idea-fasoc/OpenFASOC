* NGSPICE file created from diff_pair_sample_0008.ext - technology: sky130A

.subckt diff_pair_sample_0008 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t2 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=2.2407 ps=13.91 w=13.58 l=2.95
X1 B.t11 B.t9 B.t10 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=0 ps=0 w=13.58 l=2.95
X2 B.t8 B.t6 B.t7 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=0 ps=0 w=13.58 l=2.95
X3 VDD1.t1 VP.t1 VTAIL.t8 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=2.2407 ps=13.91 w=13.58 l=2.95
X4 VDD2.t5 VN.t0 VTAIL.t11 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=5.2962 ps=27.94 w=13.58 l=2.95
X5 VTAIL.t10 VN.t1 VDD2.t4 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=2.2407 ps=13.91 w=13.58 l=2.95
X6 VDD2.t3 VN.t2 VTAIL.t0 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=5.2962 ps=27.94 w=13.58 l=2.95
X7 B.t5 B.t3 B.t4 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=0 ps=0 w=13.58 l=2.95
X8 VDD2.t2 VN.t3 VTAIL.t3 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=2.2407 ps=13.91 w=13.58 l=2.95
X9 VDD1.t3 VP.t2 VTAIL.t7 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=5.2962 ps=27.94 w=13.58 l=2.95
X10 VDD1.t0 VP.t3 VTAIL.t6 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=5.2962 ps=27.94 w=13.58 l=2.95
X11 VTAIL.t5 VP.t4 VDD1.t4 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=2.2407 ps=13.91 w=13.58 l=2.95
X12 VDD2.t1 VN.t4 VTAIL.t2 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=2.2407 ps=13.91 w=13.58 l=2.95
X13 VDD1.t5 VP.t5 VTAIL.t4 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=2.2407 ps=13.91 w=13.58 l=2.95
X14 VTAIL.t1 VN.t5 VDD2.t0 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=2.2407 pd=13.91 as=2.2407 ps=13.91 w=13.58 l=2.95
X15 B.t2 B.t0 B.t1 w_n3594_n3684# sky130_fd_pr__pfet_01v8 ad=5.2962 pd=27.94 as=0 ps=0 w=13.58 l=2.95
R0 VP.n14 VP.n11 161.3
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n10 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n9 161.3
R5 VP.n22 VP.n21 161.3
R6 VP.n23 VP.n8 161.3
R7 VP.n48 VP.n0 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n45 VP.n1 161.3
R10 VP.n44 VP.n43 161.3
R11 VP.n42 VP.n2 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n39 VP.n3 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n35 VP.n4 161.3
R16 VP.n34 VP.n33 161.3
R17 VP.n32 VP.n5 161.3
R18 VP.n31 VP.n30 161.3
R19 VP.n29 VP.n6 161.3
R20 VP.n28 VP.n27 161.3
R21 VP.n13 VP.t5 143.483
R22 VP.n7 VP.t1 110.942
R23 VP.n36 VP.t0 110.942
R24 VP.n49 VP.t2 110.942
R25 VP.n24 VP.t3 110.942
R26 VP.n12 VP.t4 110.942
R27 VP.n26 VP.n7 109.433
R28 VP.n50 VP.n49 109.433
R29 VP.n25 VP.n24 109.433
R30 VP.n13 VP.n12 61.799
R31 VP.n34 VP.n5 51.2335
R32 VP.n43 VP.n42 51.2335
R33 VP.n18 VP.n17 51.2335
R34 VP.n26 VP.n25 51.2193
R35 VP.n30 VP.n5 29.9206
R36 VP.n43 VP.n1 29.9206
R37 VP.n18 VP.n9 29.9206
R38 VP.n29 VP.n28 24.5923
R39 VP.n30 VP.n29 24.5923
R40 VP.n35 VP.n34 24.5923
R41 VP.n37 VP.n35 24.5923
R42 VP.n41 VP.n3 24.5923
R43 VP.n42 VP.n41 24.5923
R44 VP.n47 VP.n1 24.5923
R45 VP.n48 VP.n47 24.5923
R46 VP.n22 VP.n9 24.5923
R47 VP.n23 VP.n22 24.5923
R48 VP.n16 VP.n11 24.5923
R49 VP.n17 VP.n16 24.5923
R50 VP.n37 VP.n36 12.2964
R51 VP.n36 VP.n3 12.2964
R52 VP.n12 VP.n11 12.2964
R53 VP.n14 VP.n13 5.13236
R54 VP.n28 VP.n7 1.47601
R55 VP.n49 VP.n48 1.47601
R56 VP.n24 VP.n23 1.47601
R57 VP.n25 VP.n8 0.278335
R58 VP.n27 VP.n26 0.278335
R59 VP.n50 VP.n0 0.278335
R60 VP.n15 VP.n14 0.189894
R61 VP.n15 VP.n10 0.189894
R62 VP.n19 VP.n10 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n8 0.189894
R66 VP.n27 VP.n6 0.189894
R67 VP.n31 VP.n6 0.189894
R68 VP.n32 VP.n31 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n33 VP.n4 0.189894
R71 VP.n38 VP.n4 0.189894
R72 VP.n39 VP.n38 0.189894
R73 VP.n40 VP.n39 0.189894
R74 VP.n40 VP.n2 0.189894
R75 VP.n44 VP.n2 0.189894
R76 VP.n45 VP.n44 0.189894
R77 VP.n46 VP.n45 0.189894
R78 VP.n46 VP.n0 0.189894
R79 VP VP.n50 0.153485
R80 VDD1.n68 VDD1.n0 756.745
R81 VDD1.n141 VDD1.n73 756.745
R82 VDD1.n69 VDD1.n68 585
R83 VDD1.n67 VDD1.n66 585
R84 VDD1.n4 VDD1.n3 585
R85 VDD1.n61 VDD1.n60 585
R86 VDD1.n59 VDD1.n58 585
R87 VDD1.n8 VDD1.n7 585
R88 VDD1.n53 VDD1.n52 585
R89 VDD1.n51 VDD1.n50 585
R90 VDD1.n12 VDD1.n11 585
R91 VDD1.n16 VDD1.n14 585
R92 VDD1.n45 VDD1.n44 585
R93 VDD1.n43 VDD1.n42 585
R94 VDD1.n18 VDD1.n17 585
R95 VDD1.n37 VDD1.n36 585
R96 VDD1.n35 VDD1.n34 585
R97 VDD1.n22 VDD1.n21 585
R98 VDD1.n29 VDD1.n28 585
R99 VDD1.n27 VDD1.n26 585
R100 VDD1.n98 VDD1.n97 585
R101 VDD1.n100 VDD1.n99 585
R102 VDD1.n93 VDD1.n92 585
R103 VDD1.n106 VDD1.n105 585
R104 VDD1.n108 VDD1.n107 585
R105 VDD1.n89 VDD1.n88 585
R106 VDD1.n115 VDD1.n114 585
R107 VDD1.n116 VDD1.n87 585
R108 VDD1.n118 VDD1.n117 585
R109 VDD1.n85 VDD1.n84 585
R110 VDD1.n124 VDD1.n123 585
R111 VDD1.n126 VDD1.n125 585
R112 VDD1.n81 VDD1.n80 585
R113 VDD1.n132 VDD1.n131 585
R114 VDD1.n134 VDD1.n133 585
R115 VDD1.n77 VDD1.n76 585
R116 VDD1.n140 VDD1.n139 585
R117 VDD1.n142 VDD1.n141 585
R118 VDD1.n25 VDD1.t5 329.036
R119 VDD1.n96 VDD1.t1 329.036
R120 VDD1.n68 VDD1.n67 171.744
R121 VDD1.n67 VDD1.n3 171.744
R122 VDD1.n60 VDD1.n3 171.744
R123 VDD1.n60 VDD1.n59 171.744
R124 VDD1.n59 VDD1.n7 171.744
R125 VDD1.n52 VDD1.n7 171.744
R126 VDD1.n52 VDD1.n51 171.744
R127 VDD1.n51 VDD1.n11 171.744
R128 VDD1.n16 VDD1.n11 171.744
R129 VDD1.n44 VDD1.n16 171.744
R130 VDD1.n44 VDD1.n43 171.744
R131 VDD1.n43 VDD1.n17 171.744
R132 VDD1.n36 VDD1.n17 171.744
R133 VDD1.n36 VDD1.n35 171.744
R134 VDD1.n35 VDD1.n21 171.744
R135 VDD1.n28 VDD1.n21 171.744
R136 VDD1.n28 VDD1.n27 171.744
R137 VDD1.n99 VDD1.n98 171.744
R138 VDD1.n99 VDD1.n92 171.744
R139 VDD1.n106 VDD1.n92 171.744
R140 VDD1.n107 VDD1.n106 171.744
R141 VDD1.n107 VDD1.n88 171.744
R142 VDD1.n115 VDD1.n88 171.744
R143 VDD1.n116 VDD1.n115 171.744
R144 VDD1.n117 VDD1.n116 171.744
R145 VDD1.n117 VDD1.n84 171.744
R146 VDD1.n124 VDD1.n84 171.744
R147 VDD1.n125 VDD1.n124 171.744
R148 VDD1.n125 VDD1.n80 171.744
R149 VDD1.n132 VDD1.n80 171.744
R150 VDD1.n133 VDD1.n132 171.744
R151 VDD1.n133 VDD1.n76 171.744
R152 VDD1.n140 VDD1.n76 171.744
R153 VDD1.n141 VDD1.n140 171.744
R154 VDD1.n27 VDD1.t5 85.8723
R155 VDD1.n98 VDD1.t1 85.8723
R156 VDD1.n147 VDD1.n146 73.3201
R157 VDD1.n149 VDD1.n148 72.6686
R158 VDD1 VDD1.n72 51.4309
R159 VDD1.n147 VDD1.n145 51.3174
R160 VDD1.n149 VDD1.n147 46.6086
R161 VDD1.n14 VDD1.n12 13.1884
R162 VDD1.n118 VDD1.n85 13.1884
R163 VDD1.n50 VDD1.n49 12.8005
R164 VDD1.n46 VDD1.n45 12.8005
R165 VDD1.n119 VDD1.n87 12.8005
R166 VDD1.n123 VDD1.n122 12.8005
R167 VDD1.n53 VDD1.n10 12.0247
R168 VDD1.n42 VDD1.n15 12.0247
R169 VDD1.n114 VDD1.n113 12.0247
R170 VDD1.n126 VDD1.n83 12.0247
R171 VDD1.n54 VDD1.n8 11.249
R172 VDD1.n41 VDD1.n18 11.249
R173 VDD1.n112 VDD1.n89 11.249
R174 VDD1.n127 VDD1.n81 11.249
R175 VDD1.n26 VDD1.n25 10.7239
R176 VDD1.n97 VDD1.n96 10.7239
R177 VDD1.n58 VDD1.n57 10.4732
R178 VDD1.n38 VDD1.n37 10.4732
R179 VDD1.n109 VDD1.n108 10.4732
R180 VDD1.n131 VDD1.n130 10.4732
R181 VDD1.n61 VDD1.n6 9.69747
R182 VDD1.n34 VDD1.n20 9.69747
R183 VDD1.n105 VDD1.n91 9.69747
R184 VDD1.n134 VDD1.n79 9.69747
R185 VDD1.n72 VDD1.n71 9.45567
R186 VDD1.n145 VDD1.n144 9.45567
R187 VDD1.n24 VDD1.n23 9.3005
R188 VDD1.n31 VDD1.n30 9.3005
R189 VDD1.n33 VDD1.n32 9.3005
R190 VDD1.n20 VDD1.n19 9.3005
R191 VDD1.n39 VDD1.n38 9.3005
R192 VDD1.n41 VDD1.n40 9.3005
R193 VDD1.n15 VDD1.n13 9.3005
R194 VDD1.n47 VDD1.n46 9.3005
R195 VDD1.n71 VDD1.n70 9.3005
R196 VDD1.n2 VDD1.n1 9.3005
R197 VDD1.n65 VDD1.n64 9.3005
R198 VDD1.n63 VDD1.n62 9.3005
R199 VDD1.n6 VDD1.n5 9.3005
R200 VDD1.n57 VDD1.n56 9.3005
R201 VDD1.n55 VDD1.n54 9.3005
R202 VDD1.n10 VDD1.n9 9.3005
R203 VDD1.n49 VDD1.n48 9.3005
R204 VDD1.n144 VDD1.n143 9.3005
R205 VDD1.n138 VDD1.n137 9.3005
R206 VDD1.n136 VDD1.n135 9.3005
R207 VDD1.n79 VDD1.n78 9.3005
R208 VDD1.n130 VDD1.n129 9.3005
R209 VDD1.n128 VDD1.n127 9.3005
R210 VDD1.n83 VDD1.n82 9.3005
R211 VDD1.n122 VDD1.n121 9.3005
R212 VDD1.n95 VDD1.n94 9.3005
R213 VDD1.n102 VDD1.n101 9.3005
R214 VDD1.n104 VDD1.n103 9.3005
R215 VDD1.n91 VDD1.n90 9.3005
R216 VDD1.n110 VDD1.n109 9.3005
R217 VDD1.n112 VDD1.n111 9.3005
R218 VDD1.n113 VDD1.n86 9.3005
R219 VDD1.n120 VDD1.n119 9.3005
R220 VDD1.n75 VDD1.n74 9.3005
R221 VDD1.n62 VDD1.n4 8.92171
R222 VDD1.n33 VDD1.n22 8.92171
R223 VDD1.n104 VDD1.n93 8.92171
R224 VDD1.n135 VDD1.n77 8.92171
R225 VDD1.n66 VDD1.n65 8.14595
R226 VDD1.n30 VDD1.n29 8.14595
R227 VDD1.n101 VDD1.n100 8.14595
R228 VDD1.n139 VDD1.n138 8.14595
R229 VDD1.n72 VDD1.n0 7.3702
R230 VDD1.n69 VDD1.n2 7.3702
R231 VDD1.n26 VDD1.n24 7.3702
R232 VDD1.n97 VDD1.n95 7.3702
R233 VDD1.n142 VDD1.n75 7.3702
R234 VDD1.n145 VDD1.n73 7.3702
R235 VDD1.n70 VDD1.n0 6.59444
R236 VDD1.n70 VDD1.n69 6.59444
R237 VDD1.n143 VDD1.n142 6.59444
R238 VDD1.n143 VDD1.n73 6.59444
R239 VDD1.n66 VDD1.n2 5.81868
R240 VDD1.n29 VDD1.n24 5.81868
R241 VDD1.n100 VDD1.n95 5.81868
R242 VDD1.n139 VDD1.n75 5.81868
R243 VDD1.n65 VDD1.n4 5.04292
R244 VDD1.n30 VDD1.n22 5.04292
R245 VDD1.n101 VDD1.n93 5.04292
R246 VDD1.n138 VDD1.n77 5.04292
R247 VDD1.n62 VDD1.n61 4.26717
R248 VDD1.n34 VDD1.n33 4.26717
R249 VDD1.n105 VDD1.n104 4.26717
R250 VDD1.n135 VDD1.n134 4.26717
R251 VDD1.n58 VDD1.n6 3.49141
R252 VDD1.n37 VDD1.n20 3.49141
R253 VDD1.n108 VDD1.n91 3.49141
R254 VDD1.n131 VDD1.n79 3.49141
R255 VDD1.n57 VDD1.n8 2.71565
R256 VDD1.n38 VDD1.n18 2.71565
R257 VDD1.n109 VDD1.n89 2.71565
R258 VDD1.n130 VDD1.n81 2.71565
R259 VDD1.n25 VDD1.n23 2.41282
R260 VDD1.n96 VDD1.n94 2.41282
R261 VDD1.n148 VDD1.t4 2.39409
R262 VDD1.n148 VDD1.t0 2.39409
R263 VDD1.n146 VDD1.t2 2.39409
R264 VDD1.n146 VDD1.t3 2.39409
R265 VDD1.n54 VDD1.n53 1.93989
R266 VDD1.n42 VDD1.n41 1.93989
R267 VDD1.n114 VDD1.n112 1.93989
R268 VDD1.n127 VDD1.n126 1.93989
R269 VDD1.n50 VDD1.n10 1.16414
R270 VDD1.n45 VDD1.n15 1.16414
R271 VDD1.n113 VDD1.n87 1.16414
R272 VDD1.n123 VDD1.n83 1.16414
R273 VDD1 VDD1.n149 0.649207
R274 VDD1.n49 VDD1.n12 0.388379
R275 VDD1.n46 VDD1.n14 0.388379
R276 VDD1.n119 VDD1.n118 0.388379
R277 VDD1.n122 VDD1.n85 0.388379
R278 VDD1.n71 VDD1.n1 0.155672
R279 VDD1.n64 VDD1.n1 0.155672
R280 VDD1.n64 VDD1.n63 0.155672
R281 VDD1.n63 VDD1.n5 0.155672
R282 VDD1.n56 VDD1.n5 0.155672
R283 VDD1.n56 VDD1.n55 0.155672
R284 VDD1.n55 VDD1.n9 0.155672
R285 VDD1.n48 VDD1.n9 0.155672
R286 VDD1.n48 VDD1.n47 0.155672
R287 VDD1.n47 VDD1.n13 0.155672
R288 VDD1.n40 VDD1.n13 0.155672
R289 VDD1.n40 VDD1.n39 0.155672
R290 VDD1.n39 VDD1.n19 0.155672
R291 VDD1.n32 VDD1.n19 0.155672
R292 VDD1.n32 VDD1.n31 0.155672
R293 VDD1.n31 VDD1.n23 0.155672
R294 VDD1.n102 VDD1.n94 0.155672
R295 VDD1.n103 VDD1.n102 0.155672
R296 VDD1.n103 VDD1.n90 0.155672
R297 VDD1.n110 VDD1.n90 0.155672
R298 VDD1.n111 VDD1.n110 0.155672
R299 VDD1.n111 VDD1.n86 0.155672
R300 VDD1.n120 VDD1.n86 0.155672
R301 VDD1.n121 VDD1.n120 0.155672
R302 VDD1.n121 VDD1.n82 0.155672
R303 VDD1.n128 VDD1.n82 0.155672
R304 VDD1.n129 VDD1.n128 0.155672
R305 VDD1.n129 VDD1.n78 0.155672
R306 VDD1.n136 VDD1.n78 0.155672
R307 VDD1.n137 VDD1.n136 0.155672
R308 VDD1.n137 VDD1.n74 0.155672
R309 VDD1.n144 VDD1.n74 0.155672
R310 VTAIL.n298 VTAIL.n230 756.745
R311 VTAIL.n70 VTAIL.n2 756.745
R312 VTAIL.n224 VTAIL.n156 756.745
R313 VTAIL.n148 VTAIL.n80 756.745
R314 VTAIL.n255 VTAIL.n254 585
R315 VTAIL.n257 VTAIL.n256 585
R316 VTAIL.n250 VTAIL.n249 585
R317 VTAIL.n263 VTAIL.n262 585
R318 VTAIL.n265 VTAIL.n264 585
R319 VTAIL.n246 VTAIL.n245 585
R320 VTAIL.n272 VTAIL.n271 585
R321 VTAIL.n273 VTAIL.n244 585
R322 VTAIL.n275 VTAIL.n274 585
R323 VTAIL.n242 VTAIL.n241 585
R324 VTAIL.n281 VTAIL.n280 585
R325 VTAIL.n283 VTAIL.n282 585
R326 VTAIL.n238 VTAIL.n237 585
R327 VTAIL.n289 VTAIL.n288 585
R328 VTAIL.n291 VTAIL.n290 585
R329 VTAIL.n234 VTAIL.n233 585
R330 VTAIL.n297 VTAIL.n296 585
R331 VTAIL.n299 VTAIL.n298 585
R332 VTAIL.n27 VTAIL.n26 585
R333 VTAIL.n29 VTAIL.n28 585
R334 VTAIL.n22 VTAIL.n21 585
R335 VTAIL.n35 VTAIL.n34 585
R336 VTAIL.n37 VTAIL.n36 585
R337 VTAIL.n18 VTAIL.n17 585
R338 VTAIL.n44 VTAIL.n43 585
R339 VTAIL.n45 VTAIL.n16 585
R340 VTAIL.n47 VTAIL.n46 585
R341 VTAIL.n14 VTAIL.n13 585
R342 VTAIL.n53 VTAIL.n52 585
R343 VTAIL.n55 VTAIL.n54 585
R344 VTAIL.n10 VTAIL.n9 585
R345 VTAIL.n61 VTAIL.n60 585
R346 VTAIL.n63 VTAIL.n62 585
R347 VTAIL.n6 VTAIL.n5 585
R348 VTAIL.n69 VTAIL.n68 585
R349 VTAIL.n71 VTAIL.n70 585
R350 VTAIL.n225 VTAIL.n224 585
R351 VTAIL.n223 VTAIL.n222 585
R352 VTAIL.n160 VTAIL.n159 585
R353 VTAIL.n217 VTAIL.n216 585
R354 VTAIL.n215 VTAIL.n214 585
R355 VTAIL.n164 VTAIL.n163 585
R356 VTAIL.n209 VTAIL.n208 585
R357 VTAIL.n207 VTAIL.n206 585
R358 VTAIL.n168 VTAIL.n167 585
R359 VTAIL.n172 VTAIL.n170 585
R360 VTAIL.n201 VTAIL.n200 585
R361 VTAIL.n199 VTAIL.n198 585
R362 VTAIL.n174 VTAIL.n173 585
R363 VTAIL.n193 VTAIL.n192 585
R364 VTAIL.n191 VTAIL.n190 585
R365 VTAIL.n178 VTAIL.n177 585
R366 VTAIL.n185 VTAIL.n184 585
R367 VTAIL.n183 VTAIL.n182 585
R368 VTAIL.n149 VTAIL.n148 585
R369 VTAIL.n147 VTAIL.n146 585
R370 VTAIL.n84 VTAIL.n83 585
R371 VTAIL.n141 VTAIL.n140 585
R372 VTAIL.n139 VTAIL.n138 585
R373 VTAIL.n88 VTAIL.n87 585
R374 VTAIL.n133 VTAIL.n132 585
R375 VTAIL.n131 VTAIL.n130 585
R376 VTAIL.n92 VTAIL.n91 585
R377 VTAIL.n96 VTAIL.n94 585
R378 VTAIL.n125 VTAIL.n124 585
R379 VTAIL.n123 VTAIL.n122 585
R380 VTAIL.n98 VTAIL.n97 585
R381 VTAIL.n117 VTAIL.n116 585
R382 VTAIL.n115 VTAIL.n114 585
R383 VTAIL.n102 VTAIL.n101 585
R384 VTAIL.n109 VTAIL.n108 585
R385 VTAIL.n107 VTAIL.n106 585
R386 VTAIL.n253 VTAIL.t0 329.036
R387 VTAIL.n25 VTAIL.t7 329.036
R388 VTAIL.n181 VTAIL.t6 329.036
R389 VTAIL.n105 VTAIL.t11 329.036
R390 VTAIL.n256 VTAIL.n255 171.744
R391 VTAIL.n256 VTAIL.n249 171.744
R392 VTAIL.n263 VTAIL.n249 171.744
R393 VTAIL.n264 VTAIL.n263 171.744
R394 VTAIL.n264 VTAIL.n245 171.744
R395 VTAIL.n272 VTAIL.n245 171.744
R396 VTAIL.n273 VTAIL.n272 171.744
R397 VTAIL.n274 VTAIL.n273 171.744
R398 VTAIL.n274 VTAIL.n241 171.744
R399 VTAIL.n281 VTAIL.n241 171.744
R400 VTAIL.n282 VTAIL.n281 171.744
R401 VTAIL.n282 VTAIL.n237 171.744
R402 VTAIL.n289 VTAIL.n237 171.744
R403 VTAIL.n290 VTAIL.n289 171.744
R404 VTAIL.n290 VTAIL.n233 171.744
R405 VTAIL.n297 VTAIL.n233 171.744
R406 VTAIL.n298 VTAIL.n297 171.744
R407 VTAIL.n28 VTAIL.n27 171.744
R408 VTAIL.n28 VTAIL.n21 171.744
R409 VTAIL.n35 VTAIL.n21 171.744
R410 VTAIL.n36 VTAIL.n35 171.744
R411 VTAIL.n36 VTAIL.n17 171.744
R412 VTAIL.n44 VTAIL.n17 171.744
R413 VTAIL.n45 VTAIL.n44 171.744
R414 VTAIL.n46 VTAIL.n45 171.744
R415 VTAIL.n46 VTAIL.n13 171.744
R416 VTAIL.n53 VTAIL.n13 171.744
R417 VTAIL.n54 VTAIL.n53 171.744
R418 VTAIL.n54 VTAIL.n9 171.744
R419 VTAIL.n61 VTAIL.n9 171.744
R420 VTAIL.n62 VTAIL.n61 171.744
R421 VTAIL.n62 VTAIL.n5 171.744
R422 VTAIL.n69 VTAIL.n5 171.744
R423 VTAIL.n70 VTAIL.n69 171.744
R424 VTAIL.n224 VTAIL.n223 171.744
R425 VTAIL.n223 VTAIL.n159 171.744
R426 VTAIL.n216 VTAIL.n159 171.744
R427 VTAIL.n216 VTAIL.n215 171.744
R428 VTAIL.n215 VTAIL.n163 171.744
R429 VTAIL.n208 VTAIL.n163 171.744
R430 VTAIL.n208 VTAIL.n207 171.744
R431 VTAIL.n207 VTAIL.n167 171.744
R432 VTAIL.n172 VTAIL.n167 171.744
R433 VTAIL.n200 VTAIL.n172 171.744
R434 VTAIL.n200 VTAIL.n199 171.744
R435 VTAIL.n199 VTAIL.n173 171.744
R436 VTAIL.n192 VTAIL.n173 171.744
R437 VTAIL.n192 VTAIL.n191 171.744
R438 VTAIL.n191 VTAIL.n177 171.744
R439 VTAIL.n184 VTAIL.n177 171.744
R440 VTAIL.n184 VTAIL.n183 171.744
R441 VTAIL.n148 VTAIL.n147 171.744
R442 VTAIL.n147 VTAIL.n83 171.744
R443 VTAIL.n140 VTAIL.n83 171.744
R444 VTAIL.n140 VTAIL.n139 171.744
R445 VTAIL.n139 VTAIL.n87 171.744
R446 VTAIL.n132 VTAIL.n87 171.744
R447 VTAIL.n132 VTAIL.n131 171.744
R448 VTAIL.n131 VTAIL.n91 171.744
R449 VTAIL.n96 VTAIL.n91 171.744
R450 VTAIL.n124 VTAIL.n96 171.744
R451 VTAIL.n124 VTAIL.n123 171.744
R452 VTAIL.n123 VTAIL.n97 171.744
R453 VTAIL.n116 VTAIL.n97 171.744
R454 VTAIL.n116 VTAIL.n115 171.744
R455 VTAIL.n115 VTAIL.n101 171.744
R456 VTAIL.n108 VTAIL.n101 171.744
R457 VTAIL.n108 VTAIL.n107 171.744
R458 VTAIL.n255 VTAIL.t0 85.8723
R459 VTAIL.n27 VTAIL.t7 85.8723
R460 VTAIL.n183 VTAIL.t6 85.8723
R461 VTAIL.n107 VTAIL.t11 85.8723
R462 VTAIL.n155 VTAIL.n154 55.99
R463 VTAIL.n79 VTAIL.n78 55.99
R464 VTAIL.n1 VTAIL.n0 55.9898
R465 VTAIL.n77 VTAIL.n76 55.9898
R466 VTAIL.n303 VTAIL.n302 32.5732
R467 VTAIL.n75 VTAIL.n74 32.5732
R468 VTAIL.n229 VTAIL.n228 32.5732
R469 VTAIL.n153 VTAIL.n152 32.5732
R470 VTAIL.n79 VTAIL.n77 29.7289
R471 VTAIL.n303 VTAIL.n229 26.9014
R472 VTAIL.n275 VTAIL.n242 13.1884
R473 VTAIL.n47 VTAIL.n14 13.1884
R474 VTAIL.n170 VTAIL.n168 13.1884
R475 VTAIL.n94 VTAIL.n92 13.1884
R476 VTAIL.n276 VTAIL.n244 12.8005
R477 VTAIL.n280 VTAIL.n279 12.8005
R478 VTAIL.n48 VTAIL.n16 12.8005
R479 VTAIL.n52 VTAIL.n51 12.8005
R480 VTAIL.n206 VTAIL.n205 12.8005
R481 VTAIL.n202 VTAIL.n201 12.8005
R482 VTAIL.n130 VTAIL.n129 12.8005
R483 VTAIL.n126 VTAIL.n125 12.8005
R484 VTAIL.n271 VTAIL.n270 12.0247
R485 VTAIL.n283 VTAIL.n240 12.0247
R486 VTAIL.n43 VTAIL.n42 12.0247
R487 VTAIL.n55 VTAIL.n12 12.0247
R488 VTAIL.n209 VTAIL.n166 12.0247
R489 VTAIL.n198 VTAIL.n171 12.0247
R490 VTAIL.n133 VTAIL.n90 12.0247
R491 VTAIL.n122 VTAIL.n95 12.0247
R492 VTAIL.n269 VTAIL.n246 11.249
R493 VTAIL.n284 VTAIL.n238 11.249
R494 VTAIL.n41 VTAIL.n18 11.249
R495 VTAIL.n56 VTAIL.n10 11.249
R496 VTAIL.n210 VTAIL.n164 11.249
R497 VTAIL.n197 VTAIL.n174 11.249
R498 VTAIL.n134 VTAIL.n88 11.249
R499 VTAIL.n121 VTAIL.n98 11.249
R500 VTAIL.n254 VTAIL.n253 10.7239
R501 VTAIL.n26 VTAIL.n25 10.7239
R502 VTAIL.n182 VTAIL.n181 10.7239
R503 VTAIL.n106 VTAIL.n105 10.7239
R504 VTAIL.n266 VTAIL.n265 10.4732
R505 VTAIL.n288 VTAIL.n287 10.4732
R506 VTAIL.n38 VTAIL.n37 10.4732
R507 VTAIL.n60 VTAIL.n59 10.4732
R508 VTAIL.n214 VTAIL.n213 10.4732
R509 VTAIL.n194 VTAIL.n193 10.4732
R510 VTAIL.n138 VTAIL.n137 10.4732
R511 VTAIL.n118 VTAIL.n117 10.4732
R512 VTAIL.n262 VTAIL.n248 9.69747
R513 VTAIL.n291 VTAIL.n236 9.69747
R514 VTAIL.n34 VTAIL.n20 9.69747
R515 VTAIL.n63 VTAIL.n8 9.69747
R516 VTAIL.n217 VTAIL.n162 9.69747
R517 VTAIL.n190 VTAIL.n176 9.69747
R518 VTAIL.n141 VTAIL.n86 9.69747
R519 VTAIL.n114 VTAIL.n100 9.69747
R520 VTAIL.n302 VTAIL.n301 9.45567
R521 VTAIL.n74 VTAIL.n73 9.45567
R522 VTAIL.n228 VTAIL.n227 9.45567
R523 VTAIL.n152 VTAIL.n151 9.45567
R524 VTAIL.n301 VTAIL.n300 9.3005
R525 VTAIL.n295 VTAIL.n294 9.3005
R526 VTAIL.n293 VTAIL.n292 9.3005
R527 VTAIL.n236 VTAIL.n235 9.3005
R528 VTAIL.n287 VTAIL.n286 9.3005
R529 VTAIL.n285 VTAIL.n284 9.3005
R530 VTAIL.n240 VTAIL.n239 9.3005
R531 VTAIL.n279 VTAIL.n278 9.3005
R532 VTAIL.n252 VTAIL.n251 9.3005
R533 VTAIL.n259 VTAIL.n258 9.3005
R534 VTAIL.n261 VTAIL.n260 9.3005
R535 VTAIL.n248 VTAIL.n247 9.3005
R536 VTAIL.n267 VTAIL.n266 9.3005
R537 VTAIL.n269 VTAIL.n268 9.3005
R538 VTAIL.n270 VTAIL.n243 9.3005
R539 VTAIL.n277 VTAIL.n276 9.3005
R540 VTAIL.n232 VTAIL.n231 9.3005
R541 VTAIL.n73 VTAIL.n72 9.3005
R542 VTAIL.n67 VTAIL.n66 9.3005
R543 VTAIL.n65 VTAIL.n64 9.3005
R544 VTAIL.n8 VTAIL.n7 9.3005
R545 VTAIL.n59 VTAIL.n58 9.3005
R546 VTAIL.n57 VTAIL.n56 9.3005
R547 VTAIL.n12 VTAIL.n11 9.3005
R548 VTAIL.n51 VTAIL.n50 9.3005
R549 VTAIL.n24 VTAIL.n23 9.3005
R550 VTAIL.n31 VTAIL.n30 9.3005
R551 VTAIL.n33 VTAIL.n32 9.3005
R552 VTAIL.n20 VTAIL.n19 9.3005
R553 VTAIL.n39 VTAIL.n38 9.3005
R554 VTAIL.n41 VTAIL.n40 9.3005
R555 VTAIL.n42 VTAIL.n15 9.3005
R556 VTAIL.n49 VTAIL.n48 9.3005
R557 VTAIL.n4 VTAIL.n3 9.3005
R558 VTAIL.n180 VTAIL.n179 9.3005
R559 VTAIL.n187 VTAIL.n186 9.3005
R560 VTAIL.n189 VTAIL.n188 9.3005
R561 VTAIL.n176 VTAIL.n175 9.3005
R562 VTAIL.n195 VTAIL.n194 9.3005
R563 VTAIL.n197 VTAIL.n196 9.3005
R564 VTAIL.n171 VTAIL.n169 9.3005
R565 VTAIL.n203 VTAIL.n202 9.3005
R566 VTAIL.n227 VTAIL.n226 9.3005
R567 VTAIL.n158 VTAIL.n157 9.3005
R568 VTAIL.n221 VTAIL.n220 9.3005
R569 VTAIL.n219 VTAIL.n218 9.3005
R570 VTAIL.n162 VTAIL.n161 9.3005
R571 VTAIL.n213 VTAIL.n212 9.3005
R572 VTAIL.n211 VTAIL.n210 9.3005
R573 VTAIL.n166 VTAIL.n165 9.3005
R574 VTAIL.n205 VTAIL.n204 9.3005
R575 VTAIL.n104 VTAIL.n103 9.3005
R576 VTAIL.n111 VTAIL.n110 9.3005
R577 VTAIL.n113 VTAIL.n112 9.3005
R578 VTAIL.n100 VTAIL.n99 9.3005
R579 VTAIL.n119 VTAIL.n118 9.3005
R580 VTAIL.n121 VTAIL.n120 9.3005
R581 VTAIL.n95 VTAIL.n93 9.3005
R582 VTAIL.n127 VTAIL.n126 9.3005
R583 VTAIL.n151 VTAIL.n150 9.3005
R584 VTAIL.n82 VTAIL.n81 9.3005
R585 VTAIL.n145 VTAIL.n144 9.3005
R586 VTAIL.n143 VTAIL.n142 9.3005
R587 VTAIL.n86 VTAIL.n85 9.3005
R588 VTAIL.n137 VTAIL.n136 9.3005
R589 VTAIL.n135 VTAIL.n134 9.3005
R590 VTAIL.n90 VTAIL.n89 9.3005
R591 VTAIL.n129 VTAIL.n128 9.3005
R592 VTAIL.n261 VTAIL.n250 8.92171
R593 VTAIL.n292 VTAIL.n234 8.92171
R594 VTAIL.n33 VTAIL.n22 8.92171
R595 VTAIL.n64 VTAIL.n6 8.92171
R596 VTAIL.n218 VTAIL.n160 8.92171
R597 VTAIL.n189 VTAIL.n178 8.92171
R598 VTAIL.n142 VTAIL.n84 8.92171
R599 VTAIL.n113 VTAIL.n102 8.92171
R600 VTAIL.n258 VTAIL.n257 8.14595
R601 VTAIL.n296 VTAIL.n295 8.14595
R602 VTAIL.n30 VTAIL.n29 8.14595
R603 VTAIL.n68 VTAIL.n67 8.14595
R604 VTAIL.n222 VTAIL.n221 8.14595
R605 VTAIL.n186 VTAIL.n185 8.14595
R606 VTAIL.n146 VTAIL.n145 8.14595
R607 VTAIL.n110 VTAIL.n109 8.14595
R608 VTAIL.n254 VTAIL.n252 7.3702
R609 VTAIL.n299 VTAIL.n232 7.3702
R610 VTAIL.n302 VTAIL.n230 7.3702
R611 VTAIL.n26 VTAIL.n24 7.3702
R612 VTAIL.n71 VTAIL.n4 7.3702
R613 VTAIL.n74 VTAIL.n2 7.3702
R614 VTAIL.n228 VTAIL.n156 7.3702
R615 VTAIL.n225 VTAIL.n158 7.3702
R616 VTAIL.n182 VTAIL.n180 7.3702
R617 VTAIL.n152 VTAIL.n80 7.3702
R618 VTAIL.n149 VTAIL.n82 7.3702
R619 VTAIL.n106 VTAIL.n104 7.3702
R620 VTAIL.n300 VTAIL.n299 6.59444
R621 VTAIL.n300 VTAIL.n230 6.59444
R622 VTAIL.n72 VTAIL.n71 6.59444
R623 VTAIL.n72 VTAIL.n2 6.59444
R624 VTAIL.n226 VTAIL.n156 6.59444
R625 VTAIL.n226 VTAIL.n225 6.59444
R626 VTAIL.n150 VTAIL.n80 6.59444
R627 VTAIL.n150 VTAIL.n149 6.59444
R628 VTAIL.n257 VTAIL.n252 5.81868
R629 VTAIL.n296 VTAIL.n232 5.81868
R630 VTAIL.n29 VTAIL.n24 5.81868
R631 VTAIL.n68 VTAIL.n4 5.81868
R632 VTAIL.n222 VTAIL.n158 5.81868
R633 VTAIL.n185 VTAIL.n180 5.81868
R634 VTAIL.n146 VTAIL.n82 5.81868
R635 VTAIL.n109 VTAIL.n104 5.81868
R636 VTAIL.n258 VTAIL.n250 5.04292
R637 VTAIL.n295 VTAIL.n234 5.04292
R638 VTAIL.n30 VTAIL.n22 5.04292
R639 VTAIL.n67 VTAIL.n6 5.04292
R640 VTAIL.n221 VTAIL.n160 5.04292
R641 VTAIL.n186 VTAIL.n178 5.04292
R642 VTAIL.n145 VTAIL.n84 5.04292
R643 VTAIL.n110 VTAIL.n102 5.04292
R644 VTAIL.n262 VTAIL.n261 4.26717
R645 VTAIL.n292 VTAIL.n291 4.26717
R646 VTAIL.n34 VTAIL.n33 4.26717
R647 VTAIL.n64 VTAIL.n63 4.26717
R648 VTAIL.n218 VTAIL.n217 4.26717
R649 VTAIL.n190 VTAIL.n189 4.26717
R650 VTAIL.n142 VTAIL.n141 4.26717
R651 VTAIL.n114 VTAIL.n113 4.26717
R652 VTAIL.n265 VTAIL.n248 3.49141
R653 VTAIL.n288 VTAIL.n236 3.49141
R654 VTAIL.n37 VTAIL.n20 3.49141
R655 VTAIL.n60 VTAIL.n8 3.49141
R656 VTAIL.n214 VTAIL.n162 3.49141
R657 VTAIL.n193 VTAIL.n176 3.49141
R658 VTAIL.n138 VTAIL.n86 3.49141
R659 VTAIL.n117 VTAIL.n100 3.49141
R660 VTAIL.n153 VTAIL.n79 2.82809
R661 VTAIL.n229 VTAIL.n155 2.82809
R662 VTAIL.n77 VTAIL.n75 2.82809
R663 VTAIL.n266 VTAIL.n246 2.71565
R664 VTAIL.n287 VTAIL.n238 2.71565
R665 VTAIL.n38 VTAIL.n18 2.71565
R666 VTAIL.n59 VTAIL.n10 2.71565
R667 VTAIL.n213 VTAIL.n164 2.71565
R668 VTAIL.n194 VTAIL.n174 2.71565
R669 VTAIL.n137 VTAIL.n88 2.71565
R670 VTAIL.n118 VTAIL.n98 2.71565
R671 VTAIL.n253 VTAIL.n251 2.41282
R672 VTAIL.n25 VTAIL.n23 2.41282
R673 VTAIL.n181 VTAIL.n179 2.41282
R674 VTAIL.n105 VTAIL.n103 2.41282
R675 VTAIL.n0 VTAIL.t3 2.39409
R676 VTAIL.n0 VTAIL.t1 2.39409
R677 VTAIL.n76 VTAIL.t8 2.39409
R678 VTAIL.n76 VTAIL.t9 2.39409
R679 VTAIL.n154 VTAIL.t4 2.39409
R680 VTAIL.n154 VTAIL.t5 2.39409
R681 VTAIL.n78 VTAIL.t2 2.39409
R682 VTAIL.n78 VTAIL.t10 2.39409
R683 VTAIL VTAIL.n303 2.063
R684 VTAIL.n271 VTAIL.n269 1.93989
R685 VTAIL.n284 VTAIL.n283 1.93989
R686 VTAIL.n43 VTAIL.n41 1.93989
R687 VTAIL.n56 VTAIL.n55 1.93989
R688 VTAIL.n210 VTAIL.n209 1.93989
R689 VTAIL.n198 VTAIL.n197 1.93989
R690 VTAIL.n134 VTAIL.n133 1.93989
R691 VTAIL.n122 VTAIL.n121 1.93989
R692 VTAIL.n155 VTAIL.n153 1.88412
R693 VTAIL.n75 VTAIL.n1 1.88412
R694 VTAIL.n270 VTAIL.n244 1.16414
R695 VTAIL.n280 VTAIL.n240 1.16414
R696 VTAIL.n42 VTAIL.n16 1.16414
R697 VTAIL.n52 VTAIL.n12 1.16414
R698 VTAIL.n206 VTAIL.n166 1.16414
R699 VTAIL.n201 VTAIL.n171 1.16414
R700 VTAIL.n130 VTAIL.n90 1.16414
R701 VTAIL.n125 VTAIL.n95 1.16414
R702 VTAIL VTAIL.n1 0.765586
R703 VTAIL.n276 VTAIL.n275 0.388379
R704 VTAIL.n279 VTAIL.n242 0.388379
R705 VTAIL.n48 VTAIL.n47 0.388379
R706 VTAIL.n51 VTAIL.n14 0.388379
R707 VTAIL.n205 VTAIL.n168 0.388379
R708 VTAIL.n202 VTAIL.n170 0.388379
R709 VTAIL.n129 VTAIL.n92 0.388379
R710 VTAIL.n126 VTAIL.n94 0.388379
R711 VTAIL.n259 VTAIL.n251 0.155672
R712 VTAIL.n260 VTAIL.n259 0.155672
R713 VTAIL.n260 VTAIL.n247 0.155672
R714 VTAIL.n267 VTAIL.n247 0.155672
R715 VTAIL.n268 VTAIL.n267 0.155672
R716 VTAIL.n268 VTAIL.n243 0.155672
R717 VTAIL.n277 VTAIL.n243 0.155672
R718 VTAIL.n278 VTAIL.n277 0.155672
R719 VTAIL.n278 VTAIL.n239 0.155672
R720 VTAIL.n285 VTAIL.n239 0.155672
R721 VTAIL.n286 VTAIL.n285 0.155672
R722 VTAIL.n286 VTAIL.n235 0.155672
R723 VTAIL.n293 VTAIL.n235 0.155672
R724 VTAIL.n294 VTAIL.n293 0.155672
R725 VTAIL.n294 VTAIL.n231 0.155672
R726 VTAIL.n301 VTAIL.n231 0.155672
R727 VTAIL.n31 VTAIL.n23 0.155672
R728 VTAIL.n32 VTAIL.n31 0.155672
R729 VTAIL.n32 VTAIL.n19 0.155672
R730 VTAIL.n39 VTAIL.n19 0.155672
R731 VTAIL.n40 VTAIL.n39 0.155672
R732 VTAIL.n40 VTAIL.n15 0.155672
R733 VTAIL.n49 VTAIL.n15 0.155672
R734 VTAIL.n50 VTAIL.n49 0.155672
R735 VTAIL.n50 VTAIL.n11 0.155672
R736 VTAIL.n57 VTAIL.n11 0.155672
R737 VTAIL.n58 VTAIL.n57 0.155672
R738 VTAIL.n58 VTAIL.n7 0.155672
R739 VTAIL.n65 VTAIL.n7 0.155672
R740 VTAIL.n66 VTAIL.n65 0.155672
R741 VTAIL.n66 VTAIL.n3 0.155672
R742 VTAIL.n73 VTAIL.n3 0.155672
R743 VTAIL.n227 VTAIL.n157 0.155672
R744 VTAIL.n220 VTAIL.n157 0.155672
R745 VTAIL.n220 VTAIL.n219 0.155672
R746 VTAIL.n219 VTAIL.n161 0.155672
R747 VTAIL.n212 VTAIL.n161 0.155672
R748 VTAIL.n212 VTAIL.n211 0.155672
R749 VTAIL.n211 VTAIL.n165 0.155672
R750 VTAIL.n204 VTAIL.n165 0.155672
R751 VTAIL.n204 VTAIL.n203 0.155672
R752 VTAIL.n203 VTAIL.n169 0.155672
R753 VTAIL.n196 VTAIL.n169 0.155672
R754 VTAIL.n196 VTAIL.n195 0.155672
R755 VTAIL.n195 VTAIL.n175 0.155672
R756 VTAIL.n188 VTAIL.n175 0.155672
R757 VTAIL.n188 VTAIL.n187 0.155672
R758 VTAIL.n187 VTAIL.n179 0.155672
R759 VTAIL.n151 VTAIL.n81 0.155672
R760 VTAIL.n144 VTAIL.n81 0.155672
R761 VTAIL.n144 VTAIL.n143 0.155672
R762 VTAIL.n143 VTAIL.n85 0.155672
R763 VTAIL.n136 VTAIL.n85 0.155672
R764 VTAIL.n136 VTAIL.n135 0.155672
R765 VTAIL.n135 VTAIL.n89 0.155672
R766 VTAIL.n128 VTAIL.n89 0.155672
R767 VTAIL.n128 VTAIL.n127 0.155672
R768 VTAIL.n127 VTAIL.n93 0.155672
R769 VTAIL.n120 VTAIL.n93 0.155672
R770 VTAIL.n120 VTAIL.n119 0.155672
R771 VTAIL.n119 VTAIL.n99 0.155672
R772 VTAIL.n112 VTAIL.n99 0.155672
R773 VTAIL.n112 VTAIL.n111 0.155672
R774 VTAIL.n111 VTAIL.n103 0.155672
R775 B.n427 B.n426 585
R776 B.n425 B.n128 585
R777 B.n424 B.n423 585
R778 B.n422 B.n129 585
R779 B.n421 B.n420 585
R780 B.n419 B.n130 585
R781 B.n418 B.n417 585
R782 B.n416 B.n131 585
R783 B.n415 B.n414 585
R784 B.n413 B.n132 585
R785 B.n412 B.n411 585
R786 B.n410 B.n133 585
R787 B.n409 B.n408 585
R788 B.n407 B.n134 585
R789 B.n406 B.n405 585
R790 B.n404 B.n135 585
R791 B.n403 B.n402 585
R792 B.n401 B.n136 585
R793 B.n400 B.n399 585
R794 B.n398 B.n137 585
R795 B.n397 B.n396 585
R796 B.n395 B.n138 585
R797 B.n394 B.n393 585
R798 B.n392 B.n139 585
R799 B.n391 B.n390 585
R800 B.n389 B.n140 585
R801 B.n388 B.n387 585
R802 B.n386 B.n141 585
R803 B.n385 B.n384 585
R804 B.n383 B.n142 585
R805 B.n382 B.n381 585
R806 B.n380 B.n143 585
R807 B.n379 B.n378 585
R808 B.n377 B.n144 585
R809 B.n376 B.n375 585
R810 B.n374 B.n145 585
R811 B.n373 B.n372 585
R812 B.n371 B.n146 585
R813 B.n370 B.n369 585
R814 B.n368 B.n147 585
R815 B.n367 B.n366 585
R816 B.n365 B.n148 585
R817 B.n364 B.n363 585
R818 B.n362 B.n149 585
R819 B.n361 B.n360 585
R820 B.n359 B.n150 585
R821 B.n358 B.n357 585
R822 B.n353 B.n151 585
R823 B.n352 B.n351 585
R824 B.n350 B.n152 585
R825 B.n349 B.n348 585
R826 B.n347 B.n153 585
R827 B.n346 B.n345 585
R828 B.n344 B.n154 585
R829 B.n343 B.n342 585
R830 B.n341 B.n155 585
R831 B.n339 B.n338 585
R832 B.n337 B.n158 585
R833 B.n336 B.n335 585
R834 B.n334 B.n159 585
R835 B.n333 B.n332 585
R836 B.n331 B.n160 585
R837 B.n330 B.n329 585
R838 B.n328 B.n161 585
R839 B.n327 B.n326 585
R840 B.n325 B.n162 585
R841 B.n324 B.n323 585
R842 B.n322 B.n163 585
R843 B.n321 B.n320 585
R844 B.n319 B.n164 585
R845 B.n318 B.n317 585
R846 B.n316 B.n165 585
R847 B.n315 B.n314 585
R848 B.n313 B.n166 585
R849 B.n312 B.n311 585
R850 B.n310 B.n167 585
R851 B.n309 B.n308 585
R852 B.n307 B.n168 585
R853 B.n306 B.n305 585
R854 B.n304 B.n169 585
R855 B.n303 B.n302 585
R856 B.n301 B.n170 585
R857 B.n300 B.n299 585
R858 B.n298 B.n171 585
R859 B.n297 B.n296 585
R860 B.n295 B.n172 585
R861 B.n294 B.n293 585
R862 B.n292 B.n173 585
R863 B.n291 B.n290 585
R864 B.n289 B.n174 585
R865 B.n288 B.n287 585
R866 B.n286 B.n175 585
R867 B.n285 B.n284 585
R868 B.n283 B.n176 585
R869 B.n282 B.n281 585
R870 B.n280 B.n177 585
R871 B.n279 B.n278 585
R872 B.n277 B.n178 585
R873 B.n276 B.n275 585
R874 B.n274 B.n179 585
R875 B.n273 B.n272 585
R876 B.n271 B.n180 585
R877 B.n428 B.n127 585
R878 B.n430 B.n429 585
R879 B.n431 B.n126 585
R880 B.n433 B.n432 585
R881 B.n434 B.n125 585
R882 B.n436 B.n435 585
R883 B.n437 B.n124 585
R884 B.n439 B.n438 585
R885 B.n440 B.n123 585
R886 B.n442 B.n441 585
R887 B.n443 B.n122 585
R888 B.n445 B.n444 585
R889 B.n446 B.n121 585
R890 B.n448 B.n447 585
R891 B.n449 B.n120 585
R892 B.n451 B.n450 585
R893 B.n452 B.n119 585
R894 B.n454 B.n453 585
R895 B.n455 B.n118 585
R896 B.n457 B.n456 585
R897 B.n458 B.n117 585
R898 B.n460 B.n459 585
R899 B.n461 B.n116 585
R900 B.n463 B.n462 585
R901 B.n464 B.n115 585
R902 B.n466 B.n465 585
R903 B.n467 B.n114 585
R904 B.n469 B.n468 585
R905 B.n470 B.n113 585
R906 B.n472 B.n471 585
R907 B.n473 B.n112 585
R908 B.n475 B.n474 585
R909 B.n476 B.n111 585
R910 B.n478 B.n477 585
R911 B.n479 B.n110 585
R912 B.n481 B.n480 585
R913 B.n482 B.n109 585
R914 B.n484 B.n483 585
R915 B.n485 B.n108 585
R916 B.n487 B.n486 585
R917 B.n488 B.n107 585
R918 B.n490 B.n489 585
R919 B.n491 B.n106 585
R920 B.n493 B.n492 585
R921 B.n494 B.n105 585
R922 B.n496 B.n495 585
R923 B.n497 B.n104 585
R924 B.n499 B.n498 585
R925 B.n500 B.n103 585
R926 B.n502 B.n501 585
R927 B.n503 B.n102 585
R928 B.n505 B.n504 585
R929 B.n506 B.n101 585
R930 B.n508 B.n507 585
R931 B.n509 B.n100 585
R932 B.n511 B.n510 585
R933 B.n512 B.n99 585
R934 B.n514 B.n513 585
R935 B.n515 B.n98 585
R936 B.n517 B.n516 585
R937 B.n518 B.n97 585
R938 B.n520 B.n519 585
R939 B.n521 B.n96 585
R940 B.n523 B.n522 585
R941 B.n524 B.n95 585
R942 B.n526 B.n525 585
R943 B.n527 B.n94 585
R944 B.n529 B.n528 585
R945 B.n530 B.n93 585
R946 B.n532 B.n531 585
R947 B.n533 B.n92 585
R948 B.n535 B.n534 585
R949 B.n536 B.n91 585
R950 B.n538 B.n537 585
R951 B.n539 B.n90 585
R952 B.n541 B.n540 585
R953 B.n542 B.n89 585
R954 B.n544 B.n543 585
R955 B.n545 B.n88 585
R956 B.n547 B.n546 585
R957 B.n548 B.n87 585
R958 B.n550 B.n549 585
R959 B.n551 B.n86 585
R960 B.n553 B.n552 585
R961 B.n554 B.n85 585
R962 B.n556 B.n555 585
R963 B.n557 B.n84 585
R964 B.n559 B.n558 585
R965 B.n560 B.n83 585
R966 B.n562 B.n561 585
R967 B.n563 B.n82 585
R968 B.n565 B.n564 585
R969 B.n566 B.n81 585
R970 B.n568 B.n567 585
R971 B.n722 B.n25 585
R972 B.n721 B.n720 585
R973 B.n719 B.n26 585
R974 B.n718 B.n717 585
R975 B.n716 B.n27 585
R976 B.n715 B.n714 585
R977 B.n713 B.n28 585
R978 B.n712 B.n711 585
R979 B.n710 B.n29 585
R980 B.n709 B.n708 585
R981 B.n707 B.n30 585
R982 B.n706 B.n705 585
R983 B.n704 B.n31 585
R984 B.n703 B.n702 585
R985 B.n701 B.n32 585
R986 B.n700 B.n699 585
R987 B.n698 B.n33 585
R988 B.n697 B.n696 585
R989 B.n695 B.n34 585
R990 B.n694 B.n693 585
R991 B.n692 B.n35 585
R992 B.n691 B.n690 585
R993 B.n689 B.n36 585
R994 B.n688 B.n687 585
R995 B.n686 B.n37 585
R996 B.n685 B.n684 585
R997 B.n683 B.n38 585
R998 B.n682 B.n681 585
R999 B.n680 B.n39 585
R1000 B.n679 B.n678 585
R1001 B.n677 B.n40 585
R1002 B.n676 B.n675 585
R1003 B.n674 B.n41 585
R1004 B.n673 B.n672 585
R1005 B.n671 B.n42 585
R1006 B.n670 B.n669 585
R1007 B.n668 B.n43 585
R1008 B.n667 B.n666 585
R1009 B.n665 B.n44 585
R1010 B.n664 B.n663 585
R1011 B.n662 B.n45 585
R1012 B.n661 B.n660 585
R1013 B.n659 B.n46 585
R1014 B.n658 B.n657 585
R1015 B.n656 B.n47 585
R1016 B.n655 B.n654 585
R1017 B.n653 B.n652 585
R1018 B.n651 B.n51 585
R1019 B.n650 B.n649 585
R1020 B.n648 B.n52 585
R1021 B.n647 B.n646 585
R1022 B.n645 B.n53 585
R1023 B.n644 B.n643 585
R1024 B.n642 B.n54 585
R1025 B.n641 B.n640 585
R1026 B.n639 B.n55 585
R1027 B.n637 B.n636 585
R1028 B.n635 B.n58 585
R1029 B.n634 B.n633 585
R1030 B.n632 B.n59 585
R1031 B.n631 B.n630 585
R1032 B.n629 B.n60 585
R1033 B.n628 B.n627 585
R1034 B.n626 B.n61 585
R1035 B.n625 B.n624 585
R1036 B.n623 B.n62 585
R1037 B.n622 B.n621 585
R1038 B.n620 B.n63 585
R1039 B.n619 B.n618 585
R1040 B.n617 B.n64 585
R1041 B.n616 B.n615 585
R1042 B.n614 B.n65 585
R1043 B.n613 B.n612 585
R1044 B.n611 B.n66 585
R1045 B.n610 B.n609 585
R1046 B.n608 B.n67 585
R1047 B.n607 B.n606 585
R1048 B.n605 B.n68 585
R1049 B.n604 B.n603 585
R1050 B.n602 B.n69 585
R1051 B.n601 B.n600 585
R1052 B.n599 B.n70 585
R1053 B.n598 B.n597 585
R1054 B.n596 B.n71 585
R1055 B.n595 B.n594 585
R1056 B.n593 B.n72 585
R1057 B.n592 B.n591 585
R1058 B.n590 B.n73 585
R1059 B.n589 B.n588 585
R1060 B.n587 B.n74 585
R1061 B.n586 B.n585 585
R1062 B.n584 B.n75 585
R1063 B.n583 B.n582 585
R1064 B.n581 B.n76 585
R1065 B.n580 B.n579 585
R1066 B.n578 B.n77 585
R1067 B.n577 B.n576 585
R1068 B.n575 B.n78 585
R1069 B.n574 B.n573 585
R1070 B.n572 B.n79 585
R1071 B.n571 B.n570 585
R1072 B.n569 B.n80 585
R1073 B.n724 B.n723 585
R1074 B.n725 B.n24 585
R1075 B.n727 B.n726 585
R1076 B.n728 B.n23 585
R1077 B.n730 B.n729 585
R1078 B.n731 B.n22 585
R1079 B.n733 B.n732 585
R1080 B.n734 B.n21 585
R1081 B.n736 B.n735 585
R1082 B.n737 B.n20 585
R1083 B.n739 B.n738 585
R1084 B.n740 B.n19 585
R1085 B.n742 B.n741 585
R1086 B.n743 B.n18 585
R1087 B.n745 B.n744 585
R1088 B.n746 B.n17 585
R1089 B.n748 B.n747 585
R1090 B.n749 B.n16 585
R1091 B.n751 B.n750 585
R1092 B.n752 B.n15 585
R1093 B.n754 B.n753 585
R1094 B.n755 B.n14 585
R1095 B.n757 B.n756 585
R1096 B.n758 B.n13 585
R1097 B.n760 B.n759 585
R1098 B.n761 B.n12 585
R1099 B.n763 B.n762 585
R1100 B.n764 B.n11 585
R1101 B.n766 B.n765 585
R1102 B.n767 B.n10 585
R1103 B.n769 B.n768 585
R1104 B.n770 B.n9 585
R1105 B.n772 B.n771 585
R1106 B.n773 B.n8 585
R1107 B.n775 B.n774 585
R1108 B.n776 B.n7 585
R1109 B.n778 B.n777 585
R1110 B.n779 B.n6 585
R1111 B.n781 B.n780 585
R1112 B.n782 B.n5 585
R1113 B.n784 B.n783 585
R1114 B.n785 B.n4 585
R1115 B.n787 B.n786 585
R1116 B.n788 B.n3 585
R1117 B.n790 B.n789 585
R1118 B.n791 B.n0 585
R1119 B.n2 B.n1 585
R1120 B.n204 B.n203 585
R1121 B.n205 B.n202 585
R1122 B.n207 B.n206 585
R1123 B.n208 B.n201 585
R1124 B.n210 B.n209 585
R1125 B.n211 B.n200 585
R1126 B.n213 B.n212 585
R1127 B.n214 B.n199 585
R1128 B.n216 B.n215 585
R1129 B.n217 B.n198 585
R1130 B.n219 B.n218 585
R1131 B.n220 B.n197 585
R1132 B.n222 B.n221 585
R1133 B.n223 B.n196 585
R1134 B.n225 B.n224 585
R1135 B.n226 B.n195 585
R1136 B.n228 B.n227 585
R1137 B.n229 B.n194 585
R1138 B.n231 B.n230 585
R1139 B.n232 B.n193 585
R1140 B.n234 B.n233 585
R1141 B.n235 B.n192 585
R1142 B.n237 B.n236 585
R1143 B.n238 B.n191 585
R1144 B.n240 B.n239 585
R1145 B.n241 B.n190 585
R1146 B.n243 B.n242 585
R1147 B.n244 B.n189 585
R1148 B.n246 B.n245 585
R1149 B.n247 B.n188 585
R1150 B.n249 B.n248 585
R1151 B.n250 B.n187 585
R1152 B.n252 B.n251 585
R1153 B.n253 B.n186 585
R1154 B.n255 B.n254 585
R1155 B.n256 B.n185 585
R1156 B.n258 B.n257 585
R1157 B.n259 B.n184 585
R1158 B.n261 B.n260 585
R1159 B.n262 B.n183 585
R1160 B.n264 B.n263 585
R1161 B.n265 B.n182 585
R1162 B.n267 B.n266 585
R1163 B.n268 B.n181 585
R1164 B.n270 B.n269 585
R1165 B.n271 B.n270 540.549
R1166 B.n426 B.n127 540.549
R1167 B.n569 B.n568 540.549
R1168 B.n724 B.n25 540.549
R1169 B.n354 B.t10 467.904
R1170 B.n56 B.t2 467.904
R1171 B.n156 B.t4 467.902
R1172 B.n48 B.t8 467.902
R1173 B.n355 B.t11 404.291
R1174 B.n57 B.t1 404.291
R1175 B.n157 B.t5 404.291
R1176 B.n49 B.t7 404.291
R1177 B.n156 B.t3 319.462
R1178 B.n354 B.t9 319.462
R1179 B.n56 B.t0 319.462
R1180 B.n48 B.t6 319.462
R1181 B.n793 B.n792 256.663
R1182 B.n792 B.n791 235.042
R1183 B.n792 B.n2 235.042
R1184 B.n272 B.n271 163.367
R1185 B.n272 B.n179 163.367
R1186 B.n276 B.n179 163.367
R1187 B.n277 B.n276 163.367
R1188 B.n278 B.n277 163.367
R1189 B.n278 B.n177 163.367
R1190 B.n282 B.n177 163.367
R1191 B.n283 B.n282 163.367
R1192 B.n284 B.n283 163.367
R1193 B.n284 B.n175 163.367
R1194 B.n288 B.n175 163.367
R1195 B.n289 B.n288 163.367
R1196 B.n290 B.n289 163.367
R1197 B.n290 B.n173 163.367
R1198 B.n294 B.n173 163.367
R1199 B.n295 B.n294 163.367
R1200 B.n296 B.n295 163.367
R1201 B.n296 B.n171 163.367
R1202 B.n300 B.n171 163.367
R1203 B.n301 B.n300 163.367
R1204 B.n302 B.n301 163.367
R1205 B.n302 B.n169 163.367
R1206 B.n306 B.n169 163.367
R1207 B.n307 B.n306 163.367
R1208 B.n308 B.n307 163.367
R1209 B.n308 B.n167 163.367
R1210 B.n312 B.n167 163.367
R1211 B.n313 B.n312 163.367
R1212 B.n314 B.n313 163.367
R1213 B.n314 B.n165 163.367
R1214 B.n318 B.n165 163.367
R1215 B.n319 B.n318 163.367
R1216 B.n320 B.n319 163.367
R1217 B.n320 B.n163 163.367
R1218 B.n324 B.n163 163.367
R1219 B.n325 B.n324 163.367
R1220 B.n326 B.n325 163.367
R1221 B.n326 B.n161 163.367
R1222 B.n330 B.n161 163.367
R1223 B.n331 B.n330 163.367
R1224 B.n332 B.n331 163.367
R1225 B.n332 B.n159 163.367
R1226 B.n336 B.n159 163.367
R1227 B.n337 B.n336 163.367
R1228 B.n338 B.n337 163.367
R1229 B.n338 B.n155 163.367
R1230 B.n343 B.n155 163.367
R1231 B.n344 B.n343 163.367
R1232 B.n345 B.n344 163.367
R1233 B.n345 B.n153 163.367
R1234 B.n349 B.n153 163.367
R1235 B.n350 B.n349 163.367
R1236 B.n351 B.n350 163.367
R1237 B.n351 B.n151 163.367
R1238 B.n358 B.n151 163.367
R1239 B.n359 B.n358 163.367
R1240 B.n360 B.n359 163.367
R1241 B.n360 B.n149 163.367
R1242 B.n364 B.n149 163.367
R1243 B.n365 B.n364 163.367
R1244 B.n366 B.n365 163.367
R1245 B.n366 B.n147 163.367
R1246 B.n370 B.n147 163.367
R1247 B.n371 B.n370 163.367
R1248 B.n372 B.n371 163.367
R1249 B.n372 B.n145 163.367
R1250 B.n376 B.n145 163.367
R1251 B.n377 B.n376 163.367
R1252 B.n378 B.n377 163.367
R1253 B.n378 B.n143 163.367
R1254 B.n382 B.n143 163.367
R1255 B.n383 B.n382 163.367
R1256 B.n384 B.n383 163.367
R1257 B.n384 B.n141 163.367
R1258 B.n388 B.n141 163.367
R1259 B.n389 B.n388 163.367
R1260 B.n390 B.n389 163.367
R1261 B.n390 B.n139 163.367
R1262 B.n394 B.n139 163.367
R1263 B.n395 B.n394 163.367
R1264 B.n396 B.n395 163.367
R1265 B.n396 B.n137 163.367
R1266 B.n400 B.n137 163.367
R1267 B.n401 B.n400 163.367
R1268 B.n402 B.n401 163.367
R1269 B.n402 B.n135 163.367
R1270 B.n406 B.n135 163.367
R1271 B.n407 B.n406 163.367
R1272 B.n408 B.n407 163.367
R1273 B.n408 B.n133 163.367
R1274 B.n412 B.n133 163.367
R1275 B.n413 B.n412 163.367
R1276 B.n414 B.n413 163.367
R1277 B.n414 B.n131 163.367
R1278 B.n418 B.n131 163.367
R1279 B.n419 B.n418 163.367
R1280 B.n420 B.n419 163.367
R1281 B.n420 B.n129 163.367
R1282 B.n424 B.n129 163.367
R1283 B.n425 B.n424 163.367
R1284 B.n426 B.n425 163.367
R1285 B.n568 B.n81 163.367
R1286 B.n564 B.n81 163.367
R1287 B.n564 B.n563 163.367
R1288 B.n563 B.n562 163.367
R1289 B.n562 B.n83 163.367
R1290 B.n558 B.n83 163.367
R1291 B.n558 B.n557 163.367
R1292 B.n557 B.n556 163.367
R1293 B.n556 B.n85 163.367
R1294 B.n552 B.n85 163.367
R1295 B.n552 B.n551 163.367
R1296 B.n551 B.n550 163.367
R1297 B.n550 B.n87 163.367
R1298 B.n546 B.n87 163.367
R1299 B.n546 B.n545 163.367
R1300 B.n545 B.n544 163.367
R1301 B.n544 B.n89 163.367
R1302 B.n540 B.n89 163.367
R1303 B.n540 B.n539 163.367
R1304 B.n539 B.n538 163.367
R1305 B.n538 B.n91 163.367
R1306 B.n534 B.n91 163.367
R1307 B.n534 B.n533 163.367
R1308 B.n533 B.n532 163.367
R1309 B.n532 B.n93 163.367
R1310 B.n528 B.n93 163.367
R1311 B.n528 B.n527 163.367
R1312 B.n527 B.n526 163.367
R1313 B.n526 B.n95 163.367
R1314 B.n522 B.n95 163.367
R1315 B.n522 B.n521 163.367
R1316 B.n521 B.n520 163.367
R1317 B.n520 B.n97 163.367
R1318 B.n516 B.n97 163.367
R1319 B.n516 B.n515 163.367
R1320 B.n515 B.n514 163.367
R1321 B.n514 B.n99 163.367
R1322 B.n510 B.n99 163.367
R1323 B.n510 B.n509 163.367
R1324 B.n509 B.n508 163.367
R1325 B.n508 B.n101 163.367
R1326 B.n504 B.n101 163.367
R1327 B.n504 B.n503 163.367
R1328 B.n503 B.n502 163.367
R1329 B.n502 B.n103 163.367
R1330 B.n498 B.n103 163.367
R1331 B.n498 B.n497 163.367
R1332 B.n497 B.n496 163.367
R1333 B.n496 B.n105 163.367
R1334 B.n492 B.n105 163.367
R1335 B.n492 B.n491 163.367
R1336 B.n491 B.n490 163.367
R1337 B.n490 B.n107 163.367
R1338 B.n486 B.n107 163.367
R1339 B.n486 B.n485 163.367
R1340 B.n485 B.n484 163.367
R1341 B.n484 B.n109 163.367
R1342 B.n480 B.n109 163.367
R1343 B.n480 B.n479 163.367
R1344 B.n479 B.n478 163.367
R1345 B.n478 B.n111 163.367
R1346 B.n474 B.n111 163.367
R1347 B.n474 B.n473 163.367
R1348 B.n473 B.n472 163.367
R1349 B.n472 B.n113 163.367
R1350 B.n468 B.n113 163.367
R1351 B.n468 B.n467 163.367
R1352 B.n467 B.n466 163.367
R1353 B.n466 B.n115 163.367
R1354 B.n462 B.n115 163.367
R1355 B.n462 B.n461 163.367
R1356 B.n461 B.n460 163.367
R1357 B.n460 B.n117 163.367
R1358 B.n456 B.n117 163.367
R1359 B.n456 B.n455 163.367
R1360 B.n455 B.n454 163.367
R1361 B.n454 B.n119 163.367
R1362 B.n450 B.n119 163.367
R1363 B.n450 B.n449 163.367
R1364 B.n449 B.n448 163.367
R1365 B.n448 B.n121 163.367
R1366 B.n444 B.n121 163.367
R1367 B.n444 B.n443 163.367
R1368 B.n443 B.n442 163.367
R1369 B.n442 B.n123 163.367
R1370 B.n438 B.n123 163.367
R1371 B.n438 B.n437 163.367
R1372 B.n437 B.n436 163.367
R1373 B.n436 B.n125 163.367
R1374 B.n432 B.n125 163.367
R1375 B.n432 B.n431 163.367
R1376 B.n431 B.n430 163.367
R1377 B.n430 B.n127 163.367
R1378 B.n720 B.n25 163.367
R1379 B.n720 B.n719 163.367
R1380 B.n719 B.n718 163.367
R1381 B.n718 B.n27 163.367
R1382 B.n714 B.n27 163.367
R1383 B.n714 B.n713 163.367
R1384 B.n713 B.n712 163.367
R1385 B.n712 B.n29 163.367
R1386 B.n708 B.n29 163.367
R1387 B.n708 B.n707 163.367
R1388 B.n707 B.n706 163.367
R1389 B.n706 B.n31 163.367
R1390 B.n702 B.n31 163.367
R1391 B.n702 B.n701 163.367
R1392 B.n701 B.n700 163.367
R1393 B.n700 B.n33 163.367
R1394 B.n696 B.n33 163.367
R1395 B.n696 B.n695 163.367
R1396 B.n695 B.n694 163.367
R1397 B.n694 B.n35 163.367
R1398 B.n690 B.n35 163.367
R1399 B.n690 B.n689 163.367
R1400 B.n689 B.n688 163.367
R1401 B.n688 B.n37 163.367
R1402 B.n684 B.n37 163.367
R1403 B.n684 B.n683 163.367
R1404 B.n683 B.n682 163.367
R1405 B.n682 B.n39 163.367
R1406 B.n678 B.n39 163.367
R1407 B.n678 B.n677 163.367
R1408 B.n677 B.n676 163.367
R1409 B.n676 B.n41 163.367
R1410 B.n672 B.n41 163.367
R1411 B.n672 B.n671 163.367
R1412 B.n671 B.n670 163.367
R1413 B.n670 B.n43 163.367
R1414 B.n666 B.n43 163.367
R1415 B.n666 B.n665 163.367
R1416 B.n665 B.n664 163.367
R1417 B.n664 B.n45 163.367
R1418 B.n660 B.n45 163.367
R1419 B.n660 B.n659 163.367
R1420 B.n659 B.n658 163.367
R1421 B.n658 B.n47 163.367
R1422 B.n654 B.n47 163.367
R1423 B.n654 B.n653 163.367
R1424 B.n653 B.n51 163.367
R1425 B.n649 B.n51 163.367
R1426 B.n649 B.n648 163.367
R1427 B.n648 B.n647 163.367
R1428 B.n647 B.n53 163.367
R1429 B.n643 B.n53 163.367
R1430 B.n643 B.n642 163.367
R1431 B.n642 B.n641 163.367
R1432 B.n641 B.n55 163.367
R1433 B.n636 B.n55 163.367
R1434 B.n636 B.n635 163.367
R1435 B.n635 B.n634 163.367
R1436 B.n634 B.n59 163.367
R1437 B.n630 B.n59 163.367
R1438 B.n630 B.n629 163.367
R1439 B.n629 B.n628 163.367
R1440 B.n628 B.n61 163.367
R1441 B.n624 B.n61 163.367
R1442 B.n624 B.n623 163.367
R1443 B.n623 B.n622 163.367
R1444 B.n622 B.n63 163.367
R1445 B.n618 B.n63 163.367
R1446 B.n618 B.n617 163.367
R1447 B.n617 B.n616 163.367
R1448 B.n616 B.n65 163.367
R1449 B.n612 B.n65 163.367
R1450 B.n612 B.n611 163.367
R1451 B.n611 B.n610 163.367
R1452 B.n610 B.n67 163.367
R1453 B.n606 B.n67 163.367
R1454 B.n606 B.n605 163.367
R1455 B.n605 B.n604 163.367
R1456 B.n604 B.n69 163.367
R1457 B.n600 B.n69 163.367
R1458 B.n600 B.n599 163.367
R1459 B.n599 B.n598 163.367
R1460 B.n598 B.n71 163.367
R1461 B.n594 B.n71 163.367
R1462 B.n594 B.n593 163.367
R1463 B.n593 B.n592 163.367
R1464 B.n592 B.n73 163.367
R1465 B.n588 B.n73 163.367
R1466 B.n588 B.n587 163.367
R1467 B.n587 B.n586 163.367
R1468 B.n586 B.n75 163.367
R1469 B.n582 B.n75 163.367
R1470 B.n582 B.n581 163.367
R1471 B.n581 B.n580 163.367
R1472 B.n580 B.n77 163.367
R1473 B.n576 B.n77 163.367
R1474 B.n576 B.n575 163.367
R1475 B.n575 B.n574 163.367
R1476 B.n574 B.n79 163.367
R1477 B.n570 B.n79 163.367
R1478 B.n570 B.n569 163.367
R1479 B.n725 B.n724 163.367
R1480 B.n726 B.n725 163.367
R1481 B.n726 B.n23 163.367
R1482 B.n730 B.n23 163.367
R1483 B.n731 B.n730 163.367
R1484 B.n732 B.n731 163.367
R1485 B.n732 B.n21 163.367
R1486 B.n736 B.n21 163.367
R1487 B.n737 B.n736 163.367
R1488 B.n738 B.n737 163.367
R1489 B.n738 B.n19 163.367
R1490 B.n742 B.n19 163.367
R1491 B.n743 B.n742 163.367
R1492 B.n744 B.n743 163.367
R1493 B.n744 B.n17 163.367
R1494 B.n748 B.n17 163.367
R1495 B.n749 B.n748 163.367
R1496 B.n750 B.n749 163.367
R1497 B.n750 B.n15 163.367
R1498 B.n754 B.n15 163.367
R1499 B.n755 B.n754 163.367
R1500 B.n756 B.n755 163.367
R1501 B.n756 B.n13 163.367
R1502 B.n760 B.n13 163.367
R1503 B.n761 B.n760 163.367
R1504 B.n762 B.n761 163.367
R1505 B.n762 B.n11 163.367
R1506 B.n766 B.n11 163.367
R1507 B.n767 B.n766 163.367
R1508 B.n768 B.n767 163.367
R1509 B.n768 B.n9 163.367
R1510 B.n772 B.n9 163.367
R1511 B.n773 B.n772 163.367
R1512 B.n774 B.n773 163.367
R1513 B.n774 B.n7 163.367
R1514 B.n778 B.n7 163.367
R1515 B.n779 B.n778 163.367
R1516 B.n780 B.n779 163.367
R1517 B.n780 B.n5 163.367
R1518 B.n784 B.n5 163.367
R1519 B.n785 B.n784 163.367
R1520 B.n786 B.n785 163.367
R1521 B.n786 B.n3 163.367
R1522 B.n790 B.n3 163.367
R1523 B.n791 B.n790 163.367
R1524 B.n204 B.n2 163.367
R1525 B.n205 B.n204 163.367
R1526 B.n206 B.n205 163.367
R1527 B.n206 B.n201 163.367
R1528 B.n210 B.n201 163.367
R1529 B.n211 B.n210 163.367
R1530 B.n212 B.n211 163.367
R1531 B.n212 B.n199 163.367
R1532 B.n216 B.n199 163.367
R1533 B.n217 B.n216 163.367
R1534 B.n218 B.n217 163.367
R1535 B.n218 B.n197 163.367
R1536 B.n222 B.n197 163.367
R1537 B.n223 B.n222 163.367
R1538 B.n224 B.n223 163.367
R1539 B.n224 B.n195 163.367
R1540 B.n228 B.n195 163.367
R1541 B.n229 B.n228 163.367
R1542 B.n230 B.n229 163.367
R1543 B.n230 B.n193 163.367
R1544 B.n234 B.n193 163.367
R1545 B.n235 B.n234 163.367
R1546 B.n236 B.n235 163.367
R1547 B.n236 B.n191 163.367
R1548 B.n240 B.n191 163.367
R1549 B.n241 B.n240 163.367
R1550 B.n242 B.n241 163.367
R1551 B.n242 B.n189 163.367
R1552 B.n246 B.n189 163.367
R1553 B.n247 B.n246 163.367
R1554 B.n248 B.n247 163.367
R1555 B.n248 B.n187 163.367
R1556 B.n252 B.n187 163.367
R1557 B.n253 B.n252 163.367
R1558 B.n254 B.n253 163.367
R1559 B.n254 B.n185 163.367
R1560 B.n258 B.n185 163.367
R1561 B.n259 B.n258 163.367
R1562 B.n260 B.n259 163.367
R1563 B.n260 B.n183 163.367
R1564 B.n264 B.n183 163.367
R1565 B.n265 B.n264 163.367
R1566 B.n266 B.n265 163.367
R1567 B.n266 B.n181 163.367
R1568 B.n270 B.n181 163.367
R1569 B.n157 B.n156 63.6126
R1570 B.n355 B.n354 63.6126
R1571 B.n57 B.n56 63.6126
R1572 B.n49 B.n48 63.6126
R1573 B.n340 B.n157 59.5399
R1574 B.n356 B.n355 59.5399
R1575 B.n638 B.n57 59.5399
R1576 B.n50 B.n49 59.5399
R1577 B.n428 B.n427 35.1225
R1578 B.n723 B.n722 35.1224
R1579 B.n567 B.n80 35.1224
R1580 B.n269 B.n180 35.1224
R1581 B B.n793 18.0485
R1582 B.n723 B.n24 10.6151
R1583 B.n727 B.n24 10.6151
R1584 B.n728 B.n727 10.6151
R1585 B.n729 B.n728 10.6151
R1586 B.n729 B.n22 10.6151
R1587 B.n733 B.n22 10.6151
R1588 B.n734 B.n733 10.6151
R1589 B.n735 B.n734 10.6151
R1590 B.n735 B.n20 10.6151
R1591 B.n739 B.n20 10.6151
R1592 B.n740 B.n739 10.6151
R1593 B.n741 B.n740 10.6151
R1594 B.n741 B.n18 10.6151
R1595 B.n745 B.n18 10.6151
R1596 B.n746 B.n745 10.6151
R1597 B.n747 B.n746 10.6151
R1598 B.n747 B.n16 10.6151
R1599 B.n751 B.n16 10.6151
R1600 B.n752 B.n751 10.6151
R1601 B.n753 B.n752 10.6151
R1602 B.n753 B.n14 10.6151
R1603 B.n757 B.n14 10.6151
R1604 B.n758 B.n757 10.6151
R1605 B.n759 B.n758 10.6151
R1606 B.n759 B.n12 10.6151
R1607 B.n763 B.n12 10.6151
R1608 B.n764 B.n763 10.6151
R1609 B.n765 B.n764 10.6151
R1610 B.n765 B.n10 10.6151
R1611 B.n769 B.n10 10.6151
R1612 B.n770 B.n769 10.6151
R1613 B.n771 B.n770 10.6151
R1614 B.n771 B.n8 10.6151
R1615 B.n775 B.n8 10.6151
R1616 B.n776 B.n775 10.6151
R1617 B.n777 B.n776 10.6151
R1618 B.n777 B.n6 10.6151
R1619 B.n781 B.n6 10.6151
R1620 B.n782 B.n781 10.6151
R1621 B.n783 B.n782 10.6151
R1622 B.n783 B.n4 10.6151
R1623 B.n787 B.n4 10.6151
R1624 B.n788 B.n787 10.6151
R1625 B.n789 B.n788 10.6151
R1626 B.n789 B.n0 10.6151
R1627 B.n722 B.n721 10.6151
R1628 B.n721 B.n26 10.6151
R1629 B.n717 B.n26 10.6151
R1630 B.n717 B.n716 10.6151
R1631 B.n716 B.n715 10.6151
R1632 B.n715 B.n28 10.6151
R1633 B.n711 B.n28 10.6151
R1634 B.n711 B.n710 10.6151
R1635 B.n710 B.n709 10.6151
R1636 B.n709 B.n30 10.6151
R1637 B.n705 B.n30 10.6151
R1638 B.n705 B.n704 10.6151
R1639 B.n704 B.n703 10.6151
R1640 B.n703 B.n32 10.6151
R1641 B.n699 B.n32 10.6151
R1642 B.n699 B.n698 10.6151
R1643 B.n698 B.n697 10.6151
R1644 B.n697 B.n34 10.6151
R1645 B.n693 B.n34 10.6151
R1646 B.n693 B.n692 10.6151
R1647 B.n692 B.n691 10.6151
R1648 B.n691 B.n36 10.6151
R1649 B.n687 B.n36 10.6151
R1650 B.n687 B.n686 10.6151
R1651 B.n686 B.n685 10.6151
R1652 B.n685 B.n38 10.6151
R1653 B.n681 B.n38 10.6151
R1654 B.n681 B.n680 10.6151
R1655 B.n680 B.n679 10.6151
R1656 B.n679 B.n40 10.6151
R1657 B.n675 B.n40 10.6151
R1658 B.n675 B.n674 10.6151
R1659 B.n674 B.n673 10.6151
R1660 B.n673 B.n42 10.6151
R1661 B.n669 B.n42 10.6151
R1662 B.n669 B.n668 10.6151
R1663 B.n668 B.n667 10.6151
R1664 B.n667 B.n44 10.6151
R1665 B.n663 B.n44 10.6151
R1666 B.n663 B.n662 10.6151
R1667 B.n662 B.n661 10.6151
R1668 B.n661 B.n46 10.6151
R1669 B.n657 B.n46 10.6151
R1670 B.n657 B.n656 10.6151
R1671 B.n656 B.n655 10.6151
R1672 B.n652 B.n651 10.6151
R1673 B.n651 B.n650 10.6151
R1674 B.n650 B.n52 10.6151
R1675 B.n646 B.n52 10.6151
R1676 B.n646 B.n645 10.6151
R1677 B.n645 B.n644 10.6151
R1678 B.n644 B.n54 10.6151
R1679 B.n640 B.n54 10.6151
R1680 B.n640 B.n639 10.6151
R1681 B.n637 B.n58 10.6151
R1682 B.n633 B.n58 10.6151
R1683 B.n633 B.n632 10.6151
R1684 B.n632 B.n631 10.6151
R1685 B.n631 B.n60 10.6151
R1686 B.n627 B.n60 10.6151
R1687 B.n627 B.n626 10.6151
R1688 B.n626 B.n625 10.6151
R1689 B.n625 B.n62 10.6151
R1690 B.n621 B.n62 10.6151
R1691 B.n621 B.n620 10.6151
R1692 B.n620 B.n619 10.6151
R1693 B.n619 B.n64 10.6151
R1694 B.n615 B.n64 10.6151
R1695 B.n615 B.n614 10.6151
R1696 B.n614 B.n613 10.6151
R1697 B.n613 B.n66 10.6151
R1698 B.n609 B.n66 10.6151
R1699 B.n609 B.n608 10.6151
R1700 B.n608 B.n607 10.6151
R1701 B.n607 B.n68 10.6151
R1702 B.n603 B.n68 10.6151
R1703 B.n603 B.n602 10.6151
R1704 B.n602 B.n601 10.6151
R1705 B.n601 B.n70 10.6151
R1706 B.n597 B.n70 10.6151
R1707 B.n597 B.n596 10.6151
R1708 B.n596 B.n595 10.6151
R1709 B.n595 B.n72 10.6151
R1710 B.n591 B.n72 10.6151
R1711 B.n591 B.n590 10.6151
R1712 B.n590 B.n589 10.6151
R1713 B.n589 B.n74 10.6151
R1714 B.n585 B.n74 10.6151
R1715 B.n585 B.n584 10.6151
R1716 B.n584 B.n583 10.6151
R1717 B.n583 B.n76 10.6151
R1718 B.n579 B.n76 10.6151
R1719 B.n579 B.n578 10.6151
R1720 B.n578 B.n577 10.6151
R1721 B.n577 B.n78 10.6151
R1722 B.n573 B.n78 10.6151
R1723 B.n573 B.n572 10.6151
R1724 B.n572 B.n571 10.6151
R1725 B.n571 B.n80 10.6151
R1726 B.n567 B.n566 10.6151
R1727 B.n566 B.n565 10.6151
R1728 B.n565 B.n82 10.6151
R1729 B.n561 B.n82 10.6151
R1730 B.n561 B.n560 10.6151
R1731 B.n560 B.n559 10.6151
R1732 B.n559 B.n84 10.6151
R1733 B.n555 B.n84 10.6151
R1734 B.n555 B.n554 10.6151
R1735 B.n554 B.n553 10.6151
R1736 B.n553 B.n86 10.6151
R1737 B.n549 B.n86 10.6151
R1738 B.n549 B.n548 10.6151
R1739 B.n548 B.n547 10.6151
R1740 B.n547 B.n88 10.6151
R1741 B.n543 B.n88 10.6151
R1742 B.n543 B.n542 10.6151
R1743 B.n542 B.n541 10.6151
R1744 B.n541 B.n90 10.6151
R1745 B.n537 B.n90 10.6151
R1746 B.n537 B.n536 10.6151
R1747 B.n536 B.n535 10.6151
R1748 B.n535 B.n92 10.6151
R1749 B.n531 B.n92 10.6151
R1750 B.n531 B.n530 10.6151
R1751 B.n530 B.n529 10.6151
R1752 B.n529 B.n94 10.6151
R1753 B.n525 B.n94 10.6151
R1754 B.n525 B.n524 10.6151
R1755 B.n524 B.n523 10.6151
R1756 B.n523 B.n96 10.6151
R1757 B.n519 B.n96 10.6151
R1758 B.n519 B.n518 10.6151
R1759 B.n518 B.n517 10.6151
R1760 B.n517 B.n98 10.6151
R1761 B.n513 B.n98 10.6151
R1762 B.n513 B.n512 10.6151
R1763 B.n512 B.n511 10.6151
R1764 B.n511 B.n100 10.6151
R1765 B.n507 B.n100 10.6151
R1766 B.n507 B.n506 10.6151
R1767 B.n506 B.n505 10.6151
R1768 B.n505 B.n102 10.6151
R1769 B.n501 B.n102 10.6151
R1770 B.n501 B.n500 10.6151
R1771 B.n500 B.n499 10.6151
R1772 B.n499 B.n104 10.6151
R1773 B.n495 B.n104 10.6151
R1774 B.n495 B.n494 10.6151
R1775 B.n494 B.n493 10.6151
R1776 B.n493 B.n106 10.6151
R1777 B.n489 B.n106 10.6151
R1778 B.n489 B.n488 10.6151
R1779 B.n488 B.n487 10.6151
R1780 B.n487 B.n108 10.6151
R1781 B.n483 B.n108 10.6151
R1782 B.n483 B.n482 10.6151
R1783 B.n482 B.n481 10.6151
R1784 B.n481 B.n110 10.6151
R1785 B.n477 B.n110 10.6151
R1786 B.n477 B.n476 10.6151
R1787 B.n476 B.n475 10.6151
R1788 B.n475 B.n112 10.6151
R1789 B.n471 B.n112 10.6151
R1790 B.n471 B.n470 10.6151
R1791 B.n470 B.n469 10.6151
R1792 B.n469 B.n114 10.6151
R1793 B.n465 B.n114 10.6151
R1794 B.n465 B.n464 10.6151
R1795 B.n464 B.n463 10.6151
R1796 B.n463 B.n116 10.6151
R1797 B.n459 B.n116 10.6151
R1798 B.n459 B.n458 10.6151
R1799 B.n458 B.n457 10.6151
R1800 B.n457 B.n118 10.6151
R1801 B.n453 B.n118 10.6151
R1802 B.n453 B.n452 10.6151
R1803 B.n452 B.n451 10.6151
R1804 B.n451 B.n120 10.6151
R1805 B.n447 B.n120 10.6151
R1806 B.n447 B.n446 10.6151
R1807 B.n446 B.n445 10.6151
R1808 B.n445 B.n122 10.6151
R1809 B.n441 B.n122 10.6151
R1810 B.n441 B.n440 10.6151
R1811 B.n440 B.n439 10.6151
R1812 B.n439 B.n124 10.6151
R1813 B.n435 B.n124 10.6151
R1814 B.n435 B.n434 10.6151
R1815 B.n434 B.n433 10.6151
R1816 B.n433 B.n126 10.6151
R1817 B.n429 B.n126 10.6151
R1818 B.n429 B.n428 10.6151
R1819 B.n203 B.n1 10.6151
R1820 B.n203 B.n202 10.6151
R1821 B.n207 B.n202 10.6151
R1822 B.n208 B.n207 10.6151
R1823 B.n209 B.n208 10.6151
R1824 B.n209 B.n200 10.6151
R1825 B.n213 B.n200 10.6151
R1826 B.n214 B.n213 10.6151
R1827 B.n215 B.n214 10.6151
R1828 B.n215 B.n198 10.6151
R1829 B.n219 B.n198 10.6151
R1830 B.n220 B.n219 10.6151
R1831 B.n221 B.n220 10.6151
R1832 B.n221 B.n196 10.6151
R1833 B.n225 B.n196 10.6151
R1834 B.n226 B.n225 10.6151
R1835 B.n227 B.n226 10.6151
R1836 B.n227 B.n194 10.6151
R1837 B.n231 B.n194 10.6151
R1838 B.n232 B.n231 10.6151
R1839 B.n233 B.n232 10.6151
R1840 B.n233 B.n192 10.6151
R1841 B.n237 B.n192 10.6151
R1842 B.n238 B.n237 10.6151
R1843 B.n239 B.n238 10.6151
R1844 B.n239 B.n190 10.6151
R1845 B.n243 B.n190 10.6151
R1846 B.n244 B.n243 10.6151
R1847 B.n245 B.n244 10.6151
R1848 B.n245 B.n188 10.6151
R1849 B.n249 B.n188 10.6151
R1850 B.n250 B.n249 10.6151
R1851 B.n251 B.n250 10.6151
R1852 B.n251 B.n186 10.6151
R1853 B.n255 B.n186 10.6151
R1854 B.n256 B.n255 10.6151
R1855 B.n257 B.n256 10.6151
R1856 B.n257 B.n184 10.6151
R1857 B.n261 B.n184 10.6151
R1858 B.n262 B.n261 10.6151
R1859 B.n263 B.n262 10.6151
R1860 B.n263 B.n182 10.6151
R1861 B.n267 B.n182 10.6151
R1862 B.n268 B.n267 10.6151
R1863 B.n269 B.n268 10.6151
R1864 B.n273 B.n180 10.6151
R1865 B.n274 B.n273 10.6151
R1866 B.n275 B.n274 10.6151
R1867 B.n275 B.n178 10.6151
R1868 B.n279 B.n178 10.6151
R1869 B.n280 B.n279 10.6151
R1870 B.n281 B.n280 10.6151
R1871 B.n281 B.n176 10.6151
R1872 B.n285 B.n176 10.6151
R1873 B.n286 B.n285 10.6151
R1874 B.n287 B.n286 10.6151
R1875 B.n287 B.n174 10.6151
R1876 B.n291 B.n174 10.6151
R1877 B.n292 B.n291 10.6151
R1878 B.n293 B.n292 10.6151
R1879 B.n293 B.n172 10.6151
R1880 B.n297 B.n172 10.6151
R1881 B.n298 B.n297 10.6151
R1882 B.n299 B.n298 10.6151
R1883 B.n299 B.n170 10.6151
R1884 B.n303 B.n170 10.6151
R1885 B.n304 B.n303 10.6151
R1886 B.n305 B.n304 10.6151
R1887 B.n305 B.n168 10.6151
R1888 B.n309 B.n168 10.6151
R1889 B.n310 B.n309 10.6151
R1890 B.n311 B.n310 10.6151
R1891 B.n311 B.n166 10.6151
R1892 B.n315 B.n166 10.6151
R1893 B.n316 B.n315 10.6151
R1894 B.n317 B.n316 10.6151
R1895 B.n317 B.n164 10.6151
R1896 B.n321 B.n164 10.6151
R1897 B.n322 B.n321 10.6151
R1898 B.n323 B.n322 10.6151
R1899 B.n323 B.n162 10.6151
R1900 B.n327 B.n162 10.6151
R1901 B.n328 B.n327 10.6151
R1902 B.n329 B.n328 10.6151
R1903 B.n329 B.n160 10.6151
R1904 B.n333 B.n160 10.6151
R1905 B.n334 B.n333 10.6151
R1906 B.n335 B.n334 10.6151
R1907 B.n335 B.n158 10.6151
R1908 B.n339 B.n158 10.6151
R1909 B.n342 B.n341 10.6151
R1910 B.n342 B.n154 10.6151
R1911 B.n346 B.n154 10.6151
R1912 B.n347 B.n346 10.6151
R1913 B.n348 B.n347 10.6151
R1914 B.n348 B.n152 10.6151
R1915 B.n352 B.n152 10.6151
R1916 B.n353 B.n352 10.6151
R1917 B.n357 B.n353 10.6151
R1918 B.n361 B.n150 10.6151
R1919 B.n362 B.n361 10.6151
R1920 B.n363 B.n362 10.6151
R1921 B.n363 B.n148 10.6151
R1922 B.n367 B.n148 10.6151
R1923 B.n368 B.n367 10.6151
R1924 B.n369 B.n368 10.6151
R1925 B.n369 B.n146 10.6151
R1926 B.n373 B.n146 10.6151
R1927 B.n374 B.n373 10.6151
R1928 B.n375 B.n374 10.6151
R1929 B.n375 B.n144 10.6151
R1930 B.n379 B.n144 10.6151
R1931 B.n380 B.n379 10.6151
R1932 B.n381 B.n380 10.6151
R1933 B.n381 B.n142 10.6151
R1934 B.n385 B.n142 10.6151
R1935 B.n386 B.n385 10.6151
R1936 B.n387 B.n386 10.6151
R1937 B.n387 B.n140 10.6151
R1938 B.n391 B.n140 10.6151
R1939 B.n392 B.n391 10.6151
R1940 B.n393 B.n392 10.6151
R1941 B.n393 B.n138 10.6151
R1942 B.n397 B.n138 10.6151
R1943 B.n398 B.n397 10.6151
R1944 B.n399 B.n398 10.6151
R1945 B.n399 B.n136 10.6151
R1946 B.n403 B.n136 10.6151
R1947 B.n404 B.n403 10.6151
R1948 B.n405 B.n404 10.6151
R1949 B.n405 B.n134 10.6151
R1950 B.n409 B.n134 10.6151
R1951 B.n410 B.n409 10.6151
R1952 B.n411 B.n410 10.6151
R1953 B.n411 B.n132 10.6151
R1954 B.n415 B.n132 10.6151
R1955 B.n416 B.n415 10.6151
R1956 B.n417 B.n416 10.6151
R1957 B.n417 B.n130 10.6151
R1958 B.n421 B.n130 10.6151
R1959 B.n422 B.n421 10.6151
R1960 B.n423 B.n422 10.6151
R1961 B.n423 B.n128 10.6151
R1962 B.n427 B.n128 10.6151
R1963 B.n655 B.n50 9.36635
R1964 B.n638 B.n637 9.36635
R1965 B.n340 B.n339 9.36635
R1966 B.n356 B.n150 9.36635
R1967 B.n793 B.n0 8.11757
R1968 B.n793 B.n1 8.11757
R1969 B.n652 B.n50 1.24928
R1970 B.n639 B.n638 1.24928
R1971 B.n341 B.n340 1.24928
R1972 B.n357 B.n356 1.24928
R1973 VN.n33 VN.n18 161.3
R1974 VN.n32 VN.n31 161.3
R1975 VN.n30 VN.n19 161.3
R1976 VN.n29 VN.n28 161.3
R1977 VN.n27 VN.n20 161.3
R1978 VN.n26 VN.n25 161.3
R1979 VN.n24 VN.n21 161.3
R1980 VN.n15 VN.n0 161.3
R1981 VN.n14 VN.n13 161.3
R1982 VN.n12 VN.n1 161.3
R1983 VN.n11 VN.n10 161.3
R1984 VN.n9 VN.n2 161.3
R1985 VN.n8 VN.n7 161.3
R1986 VN.n6 VN.n3 161.3
R1987 VN.n5 VN.t3 143.483
R1988 VN.n23 VN.t0 143.483
R1989 VN.n4 VN.t5 110.942
R1990 VN.n16 VN.t2 110.942
R1991 VN.n22 VN.t1 110.942
R1992 VN.n34 VN.t4 110.942
R1993 VN.n17 VN.n16 109.433
R1994 VN.n35 VN.n34 109.433
R1995 VN.n5 VN.n4 61.799
R1996 VN.n23 VN.n22 61.799
R1997 VN VN.n35 51.4982
R1998 VN.n10 VN.n9 51.2335
R1999 VN.n28 VN.n27 51.2335
R2000 VN.n10 VN.n1 29.9206
R2001 VN.n28 VN.n19 29.9206
R2002 VN.n8 VN.n3 24.5923
R2003 VN.n9 VN.n8 24.5923
R2004 VN.n14 VN.n1 24.5923
R2005 VN.n15 VN.n14 24.5923
R2006 VN.n27 VN.n26 24.5923
R2007 VN.n26 VN.n21 24.5923
R2008 VN.n33 VN.n32 24.5923
R2009 VN.n32 VN.n19 24.5923
R2010 VN.n4 VN.n3 12.2964
R2011 VN.n22 VN.n21 12.2964
R2012 VN.n24 VN.n23 5.13236
R2013 VN.n6 VN.n5 5.13236
R2014 VN.n16 VN.n15 1.47601
R2015 VN.n34 VN.n33 1.47601
R2016 VN.n35 VN.n18 0.278335
R2017 VN.n17 VN.n0 0.278335
R2018 VN.n31 VN.n18 0.189894
R2019 VN.n31 VN.n30 0.189894
R2020 VN.n30 VN.n29 0.189894
R2021 VN.n29 VN.n20 0.189894
R2022 VN.n25 VN.n20 0.189894
R2023 VN.n25 VN.n24 0.189894
R2024 VN.n7 VN.n6 0.189894
R2025 VN.n7 VN.n2 0.189894
R2026 VN.n11 VN.n2 0.189894
R2027 VN.n12 VN.n11 0.189894
R2028 VN.n13 VN.n12 0.189894
R2029 VN.n13 VN.n0 0.189894
R2030 VN VN.n17 0.153485
R2031 VDD2.n143 VDD2.n75 756.745
R2032 VDD2.n68 VDD2.n0 756.745
R2033 VDD2.n144 VDD2.n143 585
R2034 VDD2.n142 VDD2.n141 585
R2035 VDD2.n79 VDD2.n78 585
R2036 VDD2.n136 VDD2.n135 585
R2037 VDD2.n134 VDD2.n133 585
R2038 VDD2.n83 VDD2.n82 585
R2039 VDD2.n128 VDD2.n127 585
R2040 VDD2.n126 VDD2.n125 585
R2041 VDD2.n87 VDD2.n86 585
R2042 VDD2.n91 VDD2.n89 585
R2043 VDD2.n120 VDD2.n119 585
R2044 VDD2.n118 VDD2.n117 585
R2045 VDD2.n93 VDD2.n92 585
R2046 VDD2.n112 VDD2.n111 585
R2047 VDD2.n110 VDD2.n109 585
R2048 VDD2.n97 VDD2.n96 585
R2049 VDD2.n104 VDD2.n103 585
R2050 VDD2.n102 VDD2.n101 585
R2051 VDD2.n25 VDD2.n24 585
R2052 VDD2.n27 VDD2.n26 585
R2053 VDD2.n20 VDD2.n19 585
R2054 VDD2.n33 VDD2.n32 585
R2055 VDD2.n35 VDD2.n34 585
R2056 VDD2.n16 VDD2.n15 585
R2057 VDD2.n42 VDD2.n41 585
R2058 VDD2.n43 VDD2.n14 585
R2059 VDD2.n45 VDD2.n44 585
R2060 VDD2.n12 VDD2.n11 585
R2061 VDD2.n51 VDD2.n50 585
R2062 VDD2.n53 VDD2.n52 585
R2063 VDD2.n8 VDD2.n7 585
R2064 VDD2.n59 VDD2.n58 585
R2065 VDD2.n61 VDD2.n60 585
R2066 VDD2.n4 VDD2.n3 585
R2067 VDD2.n67 VDD2.n66 585
R2068 VDD2.n69 VDD2.n68 585
R2069 VDD2.n100 VDD2.t1 329.036
R2070 VDD2.n23 VDD2.t2 329.036
R2071 VDD2.n143 VDD2.n142 171.744
R2072 VDD2.n142 VDD2.n78 171.744
R2073 VDD2.n135 VDD2.n78 171.744
R2074 VDD2.n135 VDD2.n134 171.744
R2075 VDD2.n134 VDD2.n82 171.744
R2076 VDD2.n127 VDD2.n82 171.744
R2077 VDD2.n127 VDD2.n126 171.744
R2078 VDD2.n126 VDD2.n86 171.744
R2079 VDD2.n91 VDD2.n86 171.744
R2080 VDD2.n119 VDD2.n91 171.744
R2081 VDD2.n119 VDD2.n118 171.744
R2082 VDD2.n118 VDD2.n92 171.744
R2083 VDD2.n111 VDD2.n92 171.744
R2084 VDD2.n111 VDD2.n110 171.744
R2085 VDD2.n110 VDD2.n96 171.744
R2086 VDD2.n103 VDD2.n96 171.744
R2087 VDD2.n103 VDD2.n102 171.744
R2088 VDD2.n26 VDD2.n25 171.744
R2089 VDD2.n26 VDD2.n19 171.744
R2090 VDD2.n33 VDD2.n19 171.744
R2091 VDD2.n34 VDD2.n33 171.744
R2092 VDD2.n34 VDD2.n15 171.744
R2093 VDD2.n42 VDD2.n15 171.744
R2094 VDD2.n43 VDD2.n42 171.744
R2095 VDD2.n44 VDD2.n43 171.744
R2096 VDD2.n44 VDD2.n11 171.744
R2097 VDD2.n51 VDD2.n11 171.744
R2098 VDD2.n52 VDD2.n51 171.744
R2099 VDD2.n52 VDD2.n7 171.744
R2100 VDD2.n59 VDD2.n7 171.744
R2101 VDD2.n60 VDD2.n59 171.744
R2102 VDD2.n60 VDD2.n3 171.744
R2103 VDD2.n67 VDD2.n3 171.744
R2104 VDD2.n68 VDD2.n67 171.744
R2105 VDD2.n102 VDD2.t1 85.8723
R2106 VDD2.n25 VDD2.t2 85.8723
R2107 VDD2.n74 VDD2.n73 73.3201
R2108 VDD2 VDD2.n149 73.3173
R2109 VDD2.n74 VDD2.n72 51.3174
R2110 VDD2.n148 VDD2.n147 49.252
R2111 VDD2.n148 VDD2.n74 44.6118
R2112 VDD2.n89 VDD2.n87 13.1884
R2113 VDD2.n45 VDD2.n12 13.1884
R2114 VDD2.n125 VDD2.n124 12.8005
R2115 VDD2.n121 VDD2.n120 12.8005
R2116 VDD2.n46 VDD2.n14 12.8005
R2117 VDD2.n50 VDD2.n49 12.8005
R2118 VDD2.n128 VDD2.n85 12.0247
R2119 VDD2.n117 VDD2.n90 12.0247
R2120 VDD2.n41 VDD2.n40 12.0247
R2121 VDD2.n53 VDD2.n10 12.0247
R2122 VDD2.n129 VDD2.n83 11.249
R2123 VDD2.n116 VDD2.n93 11.249
R2124 VDD2.n39 VDD2.n16 11.249
R2125 VDD2.n54 VDD2.n8 11.249
R2126 VDD2.n101 VDD2.n100 10.7239
R2127 VDD2.n24 VDD2.n23 10.7239
R2128 VDD2.n133 VDD2.n132 10.4732
R2129 VDD2.n113 VDD2.n112 10.4732
R2130 VDD2.n36 VDD2.n35 10.4732
R2131 VDD2.n58 VDD2.n57 10.4732
R2132 VDD2.n136 VDD2.n81 9.69747
R2133 VDD2.n109 VDD2.n95 9.69747
R2134 VDD2.n32 VDD2.n18 9.69747
R2135 VDD2.n61 VDD2.n6 9.69747
R2136 VDD2.n147 VDD2.n146 9.45567
R2137 VDD2.n72 VDD2.n71 9.45567
R2138 VDD2.n99 VDD2.n98 9.3005
R2139 VDD2.n106 VDD2.n105 9.3005
R2140 VDD2.n108 VDD2.n107 9.3005
R2141 VDD2.n95 VDD2.n94 9.3005
R2142 VDD2.n114 VDD2.n113 9.3005
R2143 VDD2.n116 VDD2.n115 9.3005
R2144 VDD2.n90 VDD2.n88 9.3005
R2145 VDD2.n122 VDD2.n121 9.3005
R2146 VDD2.n146 VDD2.n145 9.3005
R2147 VDD2.n77 VDD2.n76 9.3005
R2148 VDD2.n140 VDD2.n139 9.3005
R2149 VDD2.n138 VDD2.n137 9.3005
R2150 VDD2.n81 VDD2.n80 9.3005
R2151 VDD2.n132 VDD2.n131 9.3005
R2152 VDD2.n130 VDD2.n129 9.3005
R2153 VDD2.n85 VDD2.n84 9.3005
R2154 VDD2.n124 VDD2.n123 9.3005
R2155 VDD2.n71 VDD2.n70 9.3005
R2156 VDD2.n65 VDD2.n64 9.3005
R2157 VDD2.n63 VDD2.n62 9.3005
R2158 VDD2.n6 VDD2.n5 9.3005
R2159 VDD2.n57 VDD2.n56 9.3005
R2160 VDD2.n55 VDD2.n54 9.3005
R2161 VDD2.n10 VDD2.n9 9.3005
R2162 VDD2.n49 VDD2.n48 9.3005
R2163 VDD2.n22 VDD2.n21 9.3005
R2164 VDD2.n29 VDD2.n28 9.3005
R2165 VDD2.n31 VDD2.n30 9.3005
R2166 VDD2.n18 VDD2.n17 9.3005
R2167 VDD2.n37 VDD2.n36 9.3005
R2168 VDD2.n39 VDD2.n38 9.3005
R2169 VDD2.n40 VDD2.n13 9.3005
R2170 VDD2.n47 VDD2.n46 9.3005
R2171 VDD2.n2 VDD2.n1 9.3005
R2172 VDD2.n137 VDD2.n79 8.92171
R2173 VDD2.n108 VDD2.n97 8.92171
R2174 VDD2.n31 VDD2.n20 8.92171
R2175 VDD2.n62 VDD2.n4 8.92171
R2176 VDD2.n141 VDD2.n140 8.14595
R2177 VDD2.n105 VDD2.n104 8.14595
R2178 VDD2.n28 VDD2.n27 8.14595
R2179 VDD2.n66 VDD2.n65 8.14595
R2180 VDD2.n147 VDD2.n75 7.3702
R2181 VDD2.n144 VDD2.n77 7.3702
R2182 VDD2.n101 VDD2.n99 7.3702
R2183 VDD2.n24 VDD2.n22 7.3702
R2184 VDD2.n69 VDD2.n2 7.3702
R2185 VDD2.n72 VDD2.n0 7.3702
R2186 VDD2.n145 VDD2.n75 6.59444
R2187 VDD2.n145 VDD2.n144 6.59444
R2188 VDD2.n70 VDD2.n69 6.59444
R2189 VDD2.n70 VDD2.n0 6.59444
R2190 VDD2.n141 VDD2.n77 5.81868
R2191 VDD2.n104 VDD2.n99 5.81868
R2192 VDD2.n27 VDD2.n22 5.81868
R2193 VDD2.n66 VDD2.n2 5.81868
R2194 VDD2.n140 VDD2.n79 5.04292
R2195 VDD2.n105 VDD2.n97 5.04292
R2196 VDD2.n28 VDD2.n20 5.04292
R2197 VDD2.n65 VDD2.n4 5.04292
R2198 VDD2.n137 VDD2.n136 4.26717
R2199 VDD2.n109 VDD2.n108 4.26717
R2200 VDD2.n32 VDD2.n31 4.26717
R2201 VDD2.n62 VDD2.n61 4.26717
R2202 VDD2.n133 VDD2.n81 3.49141
R2203 VDD2.n112 VDD2.n95 3.49141
R2204 VDD2.n35 VDD2.n18 3.49141
R2205 VDD2.n58 VDD2.n6 3.49141
R2206 VDD2.n132 VDD2.n83 2.71565
R2207 VDD2.n113 VDD2.n93 2.71565
R2208 VDD2.n36 VDD2.n16 2.71565
R2209 VDD2.n57 VDD2.n8 2.71565
R2210 VDD2.n100 VDD2.n98 2.41282
R2211 VDD2.n23 VDD2.n21 2.41282
R2212 VDD2.n149 VDD2.t4 2.39409
R2213 VDD2.n149 VDD2.t5 2.39409
R2214 VDD2.n73 VDD2.t0 2.39409
R2215 VDD2.n73 VDD2.t3 2.39409
R2216 VDD2 VDD2.n148 2.17938
R2217 VDD2.n129 VDD2.n128 1.93989
R2218 VDD2.n117 VDD2.n116 1.93989
R2219 VDD2.n41 VDD2.n39 1.93989
R2220 VDD2.n54 VDD2.n53 1.93989
R2221 VDD2.n125 VDD2.n85 1.16414
R2222 VDD2.n120 VDD2.n90 1.16414
R2223 VDD2.n40 VDD2.n14 1.16414
R2224 VDD2.n50 VDD2.n10 1.16414
R2225 VDD2.n124 VDD2.n87 0.388379
R2226 VDD2.n121 VDD2.n89 0.388379
R2227 VDD2.n46 VDD2.n45 0.388379
R2228 VDD2.n49 VDD2.n12 0.388379
R2229 VDD2.n146 VDD2.n76 0.155672
R2230 VDD2.n139 VDD2.n76 0.155672
R2231 VDD2.n139 VDD2.n138 0.155672
R2232 VDD2.n138 VDD2.n80 0.155672
R2233 VDD2.n131 VDD2.n80 0.155672
R2234 VDD2.n131 VDD2.n130 0.155672
R2235 VDD2.n130 VDD2.n84 0.155672
R2236 VDD2.n123 VDD2.n84 0.155672
R2237 VDD2.n123 VDD2.n122 0.155672
R2238 VDD2.n122 VDD2.n88 0.155672
R2239 VDD2.n115 VDD2.n88 0.155672
R2240 VDD2.n115 VDD2.n114 0.155672
R2241 VDD2.n114 VDD2.n94 0.155672
R2242 VDD2.n107 VDD2.n94 0.155672
R2243 VDD2.n107 VDD2.n106 0.155672
R2244 VDD2.n106 VDD2.n98 0.155672
R2245 VDD2.n29 VDD2.n21 0.155672
R2246 VDD2.n30 VDD2.n29 0.155672
R2247 VDD2.n30 VDD2.n17 0.155672
R2248 VDD2.n37 VDD2.n17 0.155672
R2249 VDD2.n38 VDD2.n37 0.155672
R2250 VDD2.n38 VDD2.n13 0.155672
R2251 VDD2.n47 VDD2.n13 0.155672
R2252 VDD2.n48 VDD2.n47 0.155672
R2253 VDD2.n48 VDD2.n9 0.155672
R2254 VDD2.n55 VDD2.n9 0.155672
R2255 VDD2.n56 VDD2.n55 0.155672
R2256 VDD2.n56 VDD2.n5 0.155672
R2257 VDD2.n63 VDD2.n5 0.155672
R2258 VDD2.n64 VDD2.n63 0.155672
R2259 VDD2.n64 VDD2.n1 0.155672
R2260 VDD2.n71 VDD2.n1 0.155672
C0 VP w_n3594_n3684# 7.37665f
C1 VDD1 w_n3594_n3684# 2.48492f
C2 VP VN 7.55306f
C3 VDD1 VN 0.151531f
C4 VDD2 w_n3594_n3684# 2.58116f
C5 VDD2 VN 7.7333f
C6 B VP 2.04278f
C7 VDD1 B 2.31061f
C8 VDD1 VP 8.06682f
C9 VDD2 B 2.3931f
C10 VDD2 VP 0.48842f
C11 VDD1 VDD2 1.54348f
C12 VTAIL w_n3594_n3684# 3.22034f
C13 VN VTAIL 7.90661f
C14 VN w_n3594_n3684# 6.91102f
C15 B VTAIL 4.19452f
C16 VP VTAIL 7.92089f
C17 VDD1 VTAIL 8.35978f
C18 B w_n3594_n3684# 10.6027f
C19 B VN 1.2636f
C20 VDD2 VTAIL 8.412991f
C21 VDD2 VSUBS 2.049422f
C22 VDD1 VSUBS 1.995471f
C23 VTAIL VSUBS 1.321212f
C24 VN VSUBS 6.20837f
C25 VP VSUBS 3.256511f
C26 B VSUBS 5.118188f
C27 w_n3594_n3684# VSUBS 0.162636p
C28 VDD2.n0 VSUBS 0.031638f
C29 VDD2.n1 VSUBS 0.027826f
C30 VDD2.n2 VSUBS 0.014952f
C31 VDD2.n3 VSUBS 0.035342f
C32 VDD2.n4 VSUBS 0.015832f
C33 VDD2.n5 VSUBS 0.027826f
C34 VDD2.n6 VSUBS 0.014952f
C35 VDD2.n7 VSUBS 0.035342f
C36 VDD2.n8 VSUBS 0.015832f
C37 VDD2.n9 VSUBS 0.027826f
C38 VDD2.n10 VSUBS 0.014952f
C39 VDD2.n11 VSUBS 0.035342f
C40 VDD2.n12 VSUBS 0.015392f
C41 VDD2.n13 VSUBS 0.027826f
C42 VDD2.n14 VSUBS 0.015832f
C43 VDD2.n15 VSUBS 0.035342f
C44 VDD2.n16 VSUBS 0.015832f
C45 VDD2.n17 VSUBS 0.027826f
C46 VDD2.n18 VSUBS 0.014952f
C47 VDD2.n19 VSUBS 0.035342f
C48 VDD2.n20 VSUBS 0.015832f
C49 VDD2.n21 VSUBS 1.55981f
C50 VDD2.n22 VSUBS 0.014952f
C51 VDD2.t2 VSUBS 0.076304f
C52 VDD2.n23 VSUBS 0.23902f
C53 VDD2.n24 VSUBS 0.026586f
C54 VDD2.n25 VSUBS 0.026506f
C55 VDD2.n26 VSUBS 0.035342f
C56 VDD2.n27 VSUBS 0.015832f
C57 VDD2.n28 VSUBS 0.014952f
C58 VDD2.n29 VSUBS 0.027826f
C59 VDD2.n30 VSUBS 0.027826f
C60 VDD2.n31 VSUBS 0.014952f
C61 VDD2.n32 VSUBS 0.015832f
C62 VDD2.n33 VSUBS 0.035342f
C63 VDD2.n34 VSUBS 0.035342f
C64 VDD2.n35 VSUBS 0.015832f
C65 VDD2.n36 VSUBS 0.014952f
C66 VDD2.n37 VSUBS 0.027826f
C67 VDD2.n38 VSUBS 0.027826f
C68 VDD2.n39 VSUBS 0.014952f
C69 VDD2.n40 VSUBS 0.014952f
C70 VDD2.n41 VSUBS 0.015832f
C71 VDD2.n42 VSUBS 0.035342f
C72 VDD2.n43 VSUBS 0.035342f
C73 VDD2.n44 VSUBS 0.035342f
C74 VDD2.n45 VSUBS 0.015392f
C75 VDD2.n46 VSUBS 0.014952f
C76 VDD2.n47 VSUBS 0.027826f
C77 VDD2.n48 VSUBS 0.027826f
C78 VDD2.n49 VSUBS 0.014952f
C79 VDD2.n50 VSUBS 0.015832f
C80 VDD2.n51 VSUBS 0.035342f
C81 VDD2.n52 VSUBS 0.035342f
C82 VDD2.n53 VSUBS 0.015832f
C83 VDD2.n54 VSUBS 0.014952f
C84 VDD2.n55 VSUBS 0.027826f
C85 VDD2.n56 VSUBS 0.027826f
C86 VDD2.n57 VSUBS 0.014952f
C87 VDD2.n58 VSUBS 0.015832f
C88 VDD2.n59 VSUBS 0.035342f
C89 VDD2.n60 VSUBS 0.035342f
C90 VDD2.n61 VSUBS 0.015832f
C91 VDD2.n62 VSUBS 0.014952f
C92 VDD2.n63 VSUBS 0.027826f
C93 VDD2.n64 VSUBS 0.027826f
C94 VDD2.n65 VSUBS 0.014952f
C95 VDD2.n66 VSUBS 0.015832f
C96 VDD2.n67 VSUBS 0.035342f
C97 VDD2.n68 VSUBS 0.08918f
C98 VDD2.n69 VSUBS 0.015832f
C99 VDD2.n70 VSUBS 0.014952f
C100 VDD2.n71 VSUBS 0.065078f
C101 VDD2.n72 VSUBS 0.073878f
C102 VDD2.t0 VSUBS 0.298607f
C103 VDD2.t3 VSUBS 0.298607f
C104 VDD2.n73 VSUBS 2.38603f
C105 VDD2.n74 VSUBS 3.56115f
C106 VDD2.n75 VSUBS 0.031638f
C107 VDD2.n76 VSUBS 0.027826f
C108 VDD2.n77 VSUBS 0.014952f
C109 VDD2.n78 VSUBS 0.035342f
C110 VDD2.n79 VSUBS 0.015832f
C111 VDD2.n80 VSUBS 0.027826f
C112 VDD2.n81 VSUBS 0.014952f
C113 VDD2.n82 VSUBS 0.035342f
C114 VDD2.n83 VSUBS 0.015832f
C115 VDD2.n84 VSUBS 0.027826f
C116 VDD2.n85 VSUBS 0.014952f
C117 VDD2.n86 VSUBS 0.035342f
C118 VDD2.n87 VSUBS 0.015392f
C119 VDD2.n88 VSUBS 0.027826f
C120 VDD2.n89 VSUBS 0.015392f
C121 VDD2.n90 VSUBS 0.014952f
C122 VDD2.n91 VSUBS 0.035342f
C123 VDD2.n92 VSUBS 0.035342f
C124 VDD2.n93 VSUBS 0.015832f
C125 VDD2.n94 VSUBS 0.027826f
C126 VDD2.n95 VSUBS 0.014952f
C127 VDD2.n96 VSUBS 0.035342f
C128 VDD2.n97 VSUBS 0.015832f
C129 VDD2.n98 VSUBS 1.55981f
C130 VDD2.n99 VSUBS 0.014952f
C131 VDD2.t1 VSUBS 0.076304f
C132 VDD2.n100 VSUBS 0.23902f
C133 VDD2.n101 VSUBS 0.026586f
C134 VDD2.n102 VSUBS 0.026506f
C135 VDD2.n103 VSUBS 0.035342f
C136 VDD2.n104 VSUBS 0.015832f
C137 VDD2.n105 VSUBS 0.014952f
C138 VDD2.n106 VSUBS 0.027826f
C139 VDD2.n107 VSUBS 0.027826f
C140 VDD2.n108 VSUBS 0.014952f
C141 VDD2.n109 VSUBS 0.015832f
C142 VDD2.n110 VSUBS 0.035342f
C143 VDD2.n111 VSUBS 0.035342f
C144 VDD2.n112 VSUBS 0.015832f
C145 VDD2.n113 VSUBS 0.014952f
C146 VDD2.n114 VSUBS 0.027826f
C147 VDD2.n115 VSUBS 0.027826f
C148 VDD2.n116 VSUBS 0.014952f
C149 VDD2.n117 VSUBS 0.015832f
C150 VDD2.n118 VSUBS 0.035342f
C151 VDD2.n119 VSUBS 0.035342f
C152 VDD2.n120 VSUBS 0.015832f
C153 VDD2.n121 VSUBS 0.014952f
C154 VDD2.n122 VSUBS 0.027826f
C155 VDD2.n123 VSUBS 0.027826f
C156 VDD2.n124 VSUBS 0.014952f
C157 VDD2.n125 VSUBS 0.015832f
C158 VDD2.n126 VSUBS 0.035342f
C159 VDD2.n127 VSUBS 0.035342f
C160 VDD2.n128 VSUBS 0.015832f
C161 VDD2.n129 VSUBS 0.014952f
C162 VDD2.n130 VSUBS 0.027826f
C163 VDD2.n131 VSUBS 0.027826f
C164 VDD2.n132 VSUBS 0.014952f
C165 VDD2.n133 VSUBS 0.015832f
C166 VDD2.n134 VSUBS 0.035342f
C167 VDD2.n135 VSUBS 0.035342f
C168 VDD2.n136 VSUBS 0.015832f
C169 VDD2.n137 VSUBS 0.014952f
C170 VDD2.n138 VSUBS 0.027826f
C171 VDD2.n139 VSUBS 0.027826f
C172 VDD2.n140 VSUBS 0.014952f
C173 VDD2.n141 VSUBS 0.015832f
C174 VDD2.n142 VSUBS 0.035342f
C175 VDD2.n143 VSUBS 0.08918f
C176 VDD2.n144 VSUBS 0.015832f
C177 VDD2.n145 VSUBS 0.014952f
C178 VDD2.n146 VSUBS 0.065078f
C179 VDD2.n147 VSUBS 0.064239f
C180 VDD2.n148 VSUBS 3.0929f
C181 VDD2.t4 VSUBS 0.298607f
C182 VDD2.t5 VSUBS 0.298607f
C183 VDD2.n149 VSUBS 2.38599f
C184 VN.n0 VSUBS 0.03615f
C185 VN.t2 VSUBS 3.00297f
C186 VN.n1 VSUBS 0.054336f
C187 VN.n2 VSUBS 0.027421f
C188 VN.n3 VSUBS 0.038298f
C189 VN.t3 VSUBS 3.28382f
C190 VN.t5 VSUBS 3.00297f
C191 VN.n4 VSUBS 1.13715f
C192 VN.n5 VSUBS 1.09869f
C193 VN.n6 VSUBS 0.292313f
C194 VN.n7 VSUBS 0.027421f
C195 VN.n8 VSUBS 0.050849f
C196 VN.n9 VSUBS 0.049544f
C197 VN.n10 VSUBS 0.02669f
C198 VN.n11 VSUBS 0.027421f
C199 VN.n12 VSUBS 0.027421f
C200 VN.n13 VSUBS 0.027421f
C201 VN.n14 VSUBS 0.050849f
C202 VN.n15 VSUBS 0.027253f
C203 VN.n16 VSUBS 1.14253f
C204 VN.n17 VSUBS 0.053613f
C205 VN.n18 VSUBS 0.03615f
C206 VN.t4 VSUBS 3.00297f
C207 VN.n19 VSUBS 0.054336f
C208 VN.n20 VSUBS 0.027421f
C209 VN.n21 VSUBS 0.038298f
C210 VN.t0 VSUBS 3.28382f
C211 VN.t1 VSUBS 3.00297f
C212 VN.n22 VSUBS 1.13715f
C213 VN.n23 VSUBS 1.09869f
C214 VN.n24 VSUBS 0.292313f
C215 VN.n25 VSUBS 0.027421f
C216 VN.n26 VSUBS 0.050849f
C217 VN.n27 VSUBS 0.049544f
C218 VN.n28 VSUBS 0.02669f
C219 VN.n29 VSUBS 0.027421f
C220 VN.n30 VSUBS 0.027421f
C221 VN.n31 VSUBS 0.027421f
C222 VN.n32 VSUBS 0.050849f
C223 VN.n33 VSUBS 0.027253f
C224 VN.n34 VSUBS 1.14253f
C225 VN.n35 VSUBS 1.60424f
C226 B.n0 VSUBS 0.007368f
C227 B.n1 VSUBS 0.007368f
C228 B.n2 VSUBS 0.010897f
C229 B.n3 VSUBS 0.00835f
C230 B.n4 VSUBS 0.00835f
C231 B.n5 VSUBS 0.00835f
C232 B.n6 VSUBS 0.00835f
C233 B.n7 VSUBS 0.00835f
C234 B.n8 VSUBS 0.00835f
C235 B.n9 VSUBS 0.00835f
C236 B.n10 VSUBS 0.00835f
C237 B.n11 VSUBS 0.00835f
C238 B.n12 VSUBS 0.00835f
C239 B.n13 VSUBS 0.00835f
C240 B.n14 VSUBS 0.00835f
C241 B.n15 VSUBS 0.00835f
C242 B.n16 VSUBS 0.00835f
C243 B.n17 VSUBS 0.00835f
C244 B.n18 VSUBS 0.00835f
C245 B.n19 VSUBS 0.00835f
C246 B.n20 VSUBS 0.00835f
C247 B.n21 VSUBS 0.00835f
C248 B.n22 VSUBS 0.00835f
C249 B.n23 VSUBS 0.00835f
C250 B.n24 VSUBS 0.00835f
C251 B.n25 VSUBS 0.021056f
C252 B.n26 VSUBS 0.00835f
C253 B.n27 VSUBS 0.00835f
C254 B.n28 VSUBS 0.00835f
C255 B.n29 VSUBS 0.00835f
C256 B.n30 VSUBS 0.00835f
C257 B.n31 VSUBS 0.00835f
C258 B.n32 VSUBS 0.00835f
C259 B.n33 VSUBS 0.00835f
C260 B.n34 VSUBS 0.00835f
C261 B.n35 VSUBS 0.00835f
C262 B.n36 VSUBS 0.00835f
C263 B.n37 VSUBS 0.00835f
C264 B.n38 VSUBS 0.00835f
C265 B.n39 VSUBS 0.00835f
C266 B.n40 VSUBS 0.00835f
C267 B.n41 VSUBS 0.00835f
C268 B.n42 VSUBS 0.00835f
C269 B.n43 VSUBS 0.00835f
C270 B.n44 VSUBS 0.00835f
C271 B.n45 VSUBS 0.00835f
C272 B.n46 VSUBS 0.00835f
C273 B.n47 VSUBS 0.00835f
C274 B.t7 VSUBS 0.294598f
C275 B.t8 VSUBS 0.337492f
C276 B.t6 VSUBS 2.1786f
C277 B.n48 VSUBS 0.532686f
C278 B.n49 VSUBS 0.32742f
C279 B.n50 VSUBS 0.019347f
C280 B.n51 VSUBS 0.00835f
C281 B.n52 VSUBS 0.00835f
C282 B.n53 VSUBS 0.00835f
C283 B.n54 VSUBS 0.00835f
C284 B.n55 VSUBS 0.00835f
C285 B.t1 VSUBS 0.294602f
C286 B.t2 VSUBS 0.337496f
C287 B.t0 VSUBS 2.1786f
C288 B.n56 VSUBS 0.532682f
C289 B.n57 VSUBS 0.327417f
C290 B.n58 VSUBS 0.00835f
C291 B.n59 VSUBS 0.00835f
C292 B.n60 VSUBS 0.00835f
C293 B.n61 VSUBS 0.00835f
C294 B.n62 VSUBS 0.00835f
C295 B.n63 VSUBS 0.00835f
C296 B.n64 VSUBS 0.00835f
C297 B.n65 VSUBS 0.00835f
C298 B.n66 VSUBS 0.00835f
C299 B.n67 VSUBS 0.00835f
C300 B.n68 VSUBS 0.00835f
C301 B.n69 VSUBS 0.00835f
C302 B.n70 VSUBS 0.00835f
C303 B.n71 VSUBS 0.00835f
C304 B.n72 VSUBS 0.00835f
C305 B.n73 VSUBS 0.00835f
C306 B.n74 VSUBS 0.00835f
C307 B.n75 VSUBS 0.00835f
C308 B.n76 VSUBS 0.00835f
C309 B.n77 VSUBS 0.00835f
C310 B.n78 VSUBS 0.00835f
C311 B.n79 VSUBS 0.00835f
C312 B.n80 VSUBS 0.021056f
C313 B.n81 VSUBS 0.00835f
C314 B.n82 VSUBS 0.00835f
C315 B.n83 VSUBS 0.00835f
C316 B.n84 VSUBS 0.00835f
C317 B.n85 VSUBS 0.00835f
C318 B.n86 VSUBS 0.00835f
C319 B.n87 VSUBS 0.00835f
C320 B.n88 VSUBS 0.00835f
C321 B.n89 VSUBS 0.00835f
C322 B.n90 VSUBS 0.00835f
C323 B.n91 VSUBS 0.00835f
C324 B.n92 VSUBS 0.00835f
C325 B.n93 VSUBS 0.00835f
C326 B.n94 VSUBS 0.00835f
C327 B.n95 VSUBS 0.00835f
C328 B.n96 VSUBS 0.00835f
C329 B.n97 VSUBS 0.00835f
C330 B.n98 VSUBS 0.00835f
C331 B.n99 VSUBS 0.00835f
C332 B.n100 VSUBS 0.00835f
C333 B.n101 VSUBS 0.00835f
C334 B.n102 VSUBS 0.00835f
C335 B.n103 VSUBS 0.00835f
C336 B.n104 VSUBS 0.00835f
C337 B.n105 VSUBS 0.00835f
C338 B.n106 VSUBS 0.00835f
C339 B.n107 VSUBS 0.00835f
C340 B.n108 VSUBS 0.00835f
C341 B.n109 VSUBS 0.00835f
C342 B.n110 VSUBS 0.00835f
C343 B.n111 VSUBS 0.00835f
C344 B.n112 VSUBS 0.00835f
C345 B.n113 VSUBS 0.00835f
C346 B.n114 VSUBS 0.00835f
C347 B.n115 VSUBS 0.00835f
C348 B.n116 VSUBS 0.00835f
C349 B.n117 VSUBS 0.00835f
C350 B.n118 VSUBS 0.00835f
C351 B.n119 VSUBS 0.00835f
C352 B.n120 VSUBS 0.00835f
C353 B.n121 VSUBS 0.00835f
C354 B.n122 VSUBS 0.00835f
C355 B.n123 VSUBS 0.00835f
C356 B.n124 VSUBS 0.00835f
C357 B.n125 VSUBS 0.00835f
C358 B.n126 VSUBS 0.00835f
C359 B.n127 VSUBS 0.019959f
C360 B.n128 VSUBS 0.00835f
C361 B.n129 VSUBS 0.00835f
C362 B.n130 VSUBS 0.00835f
C363 B.n131 VSUBS 0.00835f
C364 B.n132 VSUBS 0.00835f
C365 B.n133 VSUBS 0.00835f
C366 B.n134 VSUBS 0.00835f
C367 B.n135 VSUBS 0.00835f
C368 B.n136 VSUBS 0.00835f
C369 B.n137 VSUBS 0.00835f
C370 B.n138 VSUBS 0.00835f
C371 B.n139 VSUBS 0.00835f
C372 B.n140 VSUBS 0.00835f
C373 B.n141 VSUBS 0.00835f
C374 B.n142 VSUBS 0.00835f
C375 B.n143 VSUBS 0.00835f
C376 B.n144 VSUBS 0.00835f
C377 B.n145 VSUBS 0.00835f
C378 B.n146 VSUBS 0.00835f
C379 B.n147 VSUBS 0.00835f
C380 B.n148 VSUBS 0.00835f
C381 B.n149 VSUBS 0.00835f
C382 B.n150 VSUBS 0.007859f
C383 B.n151 VSUBS 0.00835f
C384 B.n152 VSUBS 0.00835f
C385 B.n153 VSUBS 0.00835f
C386 B.n154 VSUBS 0.00835f
C387 B.n155 VSUBS 0.00835f
C388 B.t5 VSUBS 0.294598f
C389 B.t4 VSUBS 0.337492f
C390 B.t3 VSUBS 2.1786f
C391 B.n156 VSUBS 0.532686f
C392 B.n157 VSUBS 0.32742f
C393 B.n158 VSUBS 0.00835f
C394 B.n159 VSUBS 0.00835f
C395 B.n160 VSUBS 0.00835f
C396 B.n161 VSUBS 0.00835f
C397 B.n162 VSUBS 0.00835f
C398 B.n163 VSUBS 0.00835f
C399 B.n164 VSUBS 0.00835f
C400 B.n165 VSUBS 0.00835f
C401 B.n166 VSUBS 0.00835f
C402 B.n167 VSUBS 0.00835f
C403 B.n168 VSUBS 0.00835f
C404 B.n169 VSUBS 0.00835f
C405 B.n170 VSUBS 0.00835f
C406 B.n171 VSUBS 0.00835f
C407 B.n172 VSUBS 0.00835f
C408 B.n173 VSUBS 0.00835f
C409 B.n174 VSUBS 0.00835f
C410 B.n175 VSUBS 0.00835f
C411 B.n176 VSUBS 0.00835f
C412 B.n177 VSUBS 0.00835f
C413 B.n178 VSUBS 0.00835f
C414 B.n179 VSUBS 0.00835f
C415 B.n180 VSUBS 0.021056f
C416 B.n181 VSUBS 0.00835f
C417 B.n182 VSUBS 0.00835f
C418 B.n183 VSUBS 0.00835f
C419 B.n184 VSUBS 0.00835f
C420 B.n185 VSUBS 0.00835f
C421 B.n186 VSUBS 0.00835f
C422 B.n187 VSUBS 0.00835f
C423 B.n188 VSUBS 0.00835f
C424 B.n189 VSUBS 0.00835f
C425 B.n190 VSUBS 0.00835f
C426 B.n191 VSUBS 0.00835f
C427 B.n192 VSUBS 0.00835f
C428 B.n193 VSUBS 0.00835f
C429 B.n194 VSUBS 0.00835f
C430 B.n195 VSUBS 0.00835f
C431 B.n196 VSUBS 0.00835f
C432 B.n197 VSUBS 0.00835f
C433 B.n198 VSUBS 0.00835f
C434 B.n199 VSUBS 0.00835f
C435 B.n200 VSUBS 0.00835f
C436 B.n201 VSUBS 0.00835f
C437 B.n202 VSUBS 0.00835f
C438 B.n203 VSUBS 0.00835f
C439 B.n204 VSUBS 0.00835f
C440 B.n205 VSUBS 0.00835f
C441 B.n206 VSUBS 0.00835f
C442 B.n207 VSUBS 0.00835f
C443 B.n208 VSUBS 0.00835f
C444 B.n209 VSUBS 0.00835f
C445 B.n210 VSUBS 0.00835f
C446 B.n211 VSUBS 0.00835f
C447 B.n212 VSUBS 0.00835f
C448 B.n213 VSUBS 0.00835f
C449 B.n214 VSUBS 0.00835f
C450 B.n215 VSUBS 0.00835f
C451 B.n216 VSUBS 0.00835f
C452 B.n217 VSUBS 0.00835f
C453 B.n218 VSUBS 0.00835f
C454 B.n219 VSUBS 0.00835f
C455 B.n220 VSUBS 0.00835f
C456 B.n221 VSUBS 0.00835f
C457 B.n222 VSUBS 0.00835f
C458 B.n223 VSUBS 0.00835f
C459 B.n224 VSUBS 0.00835f
C460 B.n225 VSUBS 0.00835f
C461 B.n226 VSUBS 0.00835f
C462 B.n227 VSUBS 0.00835f
C463 B.n228 VSUBS 0.00835f
C464 B.n229 VSUBS 0.00835f
C465 B.n230 VSUBS 0.00835f
C466 B.n231 VSUBS 0.00835f
C467 B.n232 VSUBS 0.00835f
C468 B.n233 VSUBS 0.00835f
C469 B.n234 VSUBS 0.00835f
C470 B.n235 VSUBS 0.00835f
C471 B.n236 VSUBS 0.00835f
C472 B.n237 VSUBS 0.00835f
C473 B.n238 VSUBS 0.00835f
C474 B.n239 VSUBS 0.00835f
C475 B.n240 VSUBS 0.00835f
C476 B.n241 VSUBS 0.00835f
C477 B.n242 VSUBS 0.00835f
C478 B.n243 VSUBS 0.00835f
C479 B.n244 VSUBS 0.00835f
C480 B.n245 VSUBS 0.00835f
C481 B.n246 VSUBS 0.00835f
C482 B.n247 VSUBS 0.00835f
C483 B.n248 VSUBS 0.00835f
C484 B.n249 VSUBS 0.00835f
C485 B.n250 VSUBS 0.00835f
C486 B.n251 VSUBS 0.00835f
C487 B.n252 VSUBS 0.00835f
C488 B.n253 VSUBS 0.00835f
C489 B.n254 VSUBS 0.00835f
C490 B.n255 VSUBS 0.00835f
C491 B.n256 VSUBS 0.00835f
C492 B.n257 VSUBS 0.00835f
C493 B.n258 VSUBS 0.00835f
C494 B.n259 VSUBS 0.00835f
C495 B.n260 VSUBS 0.00835f
C496 B.n261 VSUBS 0.00835f
C497 B.n262 VSUBS 0.00835f
C498 B.n263 VSUBS 0.00835f
C499 B.n264 VSUBS 0.00835f
C500 B.n265 VSUBS 0.00835f
C501 B.n266 VSUBS 0.00835f
C502 B.n267 VSUBS 0.00835f
C503 B.n268 VSUBS 0.00835f
C504 B.n269 VSUBS 0.019959f
C505 B.n270 VSUBS 0.019959f
C506 B.n271 VSUBS 0.021056f
C507 B.n272 VSUBS 0.00835f
C508 B.n273 VSUBS 0.00835f
C509 B.n274 VSUBS 0.00835f
C510 B.n275 VSUBS 0.00835f
C511 B.n276 VSUBS 0.00835f
C512 B.n277 VSUBS 0.00835f
C513 B.n278 VSUBS 0.00835f
C514 B.n279 VSUBS 0.00835f
C515 B.n280 VSUBS 0.00835f
C516 B.n281 VSUBS 0.00835f
C517 B.n282 VSUBS 0.00835f
C518 B.n283 VSUBS 0.00835f
C519 B.n284 VSUBS 0.00835f
C520 B.n285 VSUBS 0.00835f
C521 B.n286 VSUBS 0.00835f
C522 B.n287 VSUBS 0.00835f
C523 B.n288 VSUBS 0.00835f
C524 B.n289 VSUBS 0.00835f
C525 B.n290 VSUBS 0.00835f
C526 B.n291 VSUBS 0.00835f
C527 B.n292 VSUBS 0.00835f
C528 B.n293 VSUBS 0.00835f
C529 B.n294 VSUBS 0.00835f
C530 B.n295 VSUBS 0.00835f
C531 B.n296 VSUBS 0.00835f
C532 B.n297 VSUBS 0.00835f
C533 B.n298 VSUBS 0.00835f
C534 B.n299 VSUBS 0.00835f
C535 B.n300 VSUBS 0.00835f
C536 B.n301 VSUBS 0.00835f
C537 B.n302 VSUBS 0.00835f
C538 B.n303 VSUBS 0.00835f
C539 B.n304 VSUBS 0.00835f
C540 B.n305 VSUBS 0.00835f
C541 B.n306 VSUBS 0.00835f
C542 B.n307 VSUBS 0.00835f
C543 B.n308 VSUBS 0.00835f
C544 B.n309 VSUBS 0.00835f
C545 B.n310 VSUBS 0.00835f
C546 B.n311 VSUBS 0.00835f
C547 B.n312 VSUBS 0.00835f
C548 B.n313 VSUBS 0.00835f
C549 B.n314 VSUBS 0.00835f
C550 B.n315 VSUBS 0.00835f
C551 B.n316 VSUBS 0.00835f
C552 B.n317 VSUBS 0.00835f
C553 B.n318 VSUBS 0.00835f
C554 B.n319 VSUBS 0.00835f
C555 B.n320 VSUBS 0.00835f
C556 B.n321 VSUBS 0.00835f
C557 B.n322 VSUBS 0.00835f
C558 B.n323 VSUBS 0.00835f
C559 B.n324 VSUBS 0.00835f
C560 B.n325 VSUBS 0.00835f
C561 B.n326 VSUBS 0.00835f
C562 B.n327 VSUBS 0.00835f
C563 B.n328 VSUBS 0.00835f
C564 B.n329 VSUBS 0.00835f
C565 B.n330 VSUBS 0.00835f
C566 B.n331 VSUBS 0.00835f
C567 B.n332 VSUBS 0.00835f
C568 B.n333 VSUBS 0.00835f
C569 B.n334 VSUBS 0.00835f
C570 B.n335 VSUBS 0.00835f
C571 B.n336 VSUBS 0.00835f
C572 B.n337 VSUBS 0.00835f
C573 B.n338 VSUBS 0.00835f
C574 B.n339 VSUBS 0.007859f
C575 B.n340 VSUBS 0.019347f
C576 B.n341 VSUBS 0.004666f
C577 B.n342 VSUBS 0.00835f
C578 B.n343 VSUBS 0.00835f
C579 B.n344 VSUBS 0.00835f
C580 B.n345 VSUBS 0.00835f
C581 B.n346 VSUBS 0.00835f
C582 B.n347 VSUBS 0.00835f
C583 B.n348 VSUBS 0.00835f
C584 B.n349 VSUBS 0.00835f
C585 B.n350 VSUBS 0.00835f
C586 B.n351 VSUBS 0.00835f
C587 B.n352 VSUBS 0.00835f
C588 B.n353 VSUBS 0.00835f
C589 B.t11 VSUBS 0.294602f
C590 B.t10 VSUBS 0.337496f
C591 B.t9 VSUBS 2.1786f
C592 B.n354 VSUBS 0.532682f
C593 B.n355 VSUBS 0.327417f
C594 B.n356 VSUBS 0.019347f
C595 B.n357 VSUBS 0.004666f
C596 B.n358 VSUBS 0.00835f
C597 B.n359 VSUBS 0.00835f
C598 B.n360 VSUBS 0.00835f
C599 B.n361 VSUBS 0.00835f
C600 B.n362 VSUBS 0.00835f
C601 B.n363 VSUBS 0.00835f
C602 B.n364 VSUBS 0.00835f
C603 B.n365 VSUBS 0.00835f
C604 B.n366 VSUBS 0.00835f
C605 B.n367 VSUBS 0.00835f
C606 B.n368 VSUBS 0.00835f
C607 B.n369 VSUBS 0.00835f
C608 B.n370 VSUBS 0.00835f
C609 B.n371 VSUBS 0.00835f
C610 B.n372 VSUBS 0.00835f
C611 B.n373 VSUBS 0.00835f
C612 B.n374 VSUBS 0.00835f
C613 B.n375 VSUBS 0.00835f
C614 B.n376 VSUBS 0.00835f
C615 B.n377 VSUBS 0.00835f
C616 B.n378 VSUBS 0.00835f
C617 B.n379 VSUBS 0.00835f
C618 B.n380 VSUBS 0.00835f
C619 B.n381 VSUBS 0.00835f
C620 B.n382 VSUBS 0.00835f
C621 B.n383 VSUBS 0.00835f
C622 B.n384 VSUBS 0.00835f
C623 B.n385 VSUBS 0.00835f
C624 B.n386 VSUBS 0.00835f
C625 B.n387 VSUBS 0.00835f
C626 B.n388 VSUBS 0.00835f
C627 B.n389 VSUBS 0.00835f
C628 B.n390 VSUBS 0.00835f
C629 B.n391 VSUBS 0.00835f
C630 B.n392 VSUBS 0.00835f
C631 B.n393 VSUBS 0.00835f
C632 B.n394 VSUBS 0.00835f
C633 B.n395 VSUBS 0.00835f
C634 B.n396 VSUBS 0.00835f
C635 B.n397 VSUBS 0.00835f
C636 B.n398 VSUBS 0.00835f
C637 B.n399 VSUBS 0.00835f
C638 B.n400 VSUBS 0.00835f
C639 B.n401 VSUBS 0.00835f
C640 B.n402 VSUBS 0.00835f
C641 B.n403 VSUBS 0.00835f
C642 B.n404 VSUBS 0.00835f
C643 B.n405 VSUBS 0.00835f
C644 B.n406 VSUBS 0.00835f
C645 B.n407 VSUBS 0.00835f
C646 B.n408 VSUBS 0.00835f
C647 B.n409 VSUBS 0.00835f
C648 B.n410 VSUBS 0.00835f
C649 B.n411 VSUBS 0.00835f
C650 B.n412 VSUBS 0.00835f
C651 B.n413 VSUBS 0.00835f
C652 B.n414 VSUBS 0.00835f
C653 B.n415 VSUBS 0.00835f
C654 B.n416 VSUBS 0.00835f
C655 B.n417 VSUBS 0.00835f
C656 B.n418 VSUBS 0.00835f
C657 B.n419 VSUBS 0.00835f
C658 B.n420 VSUBS 0.00835f
C659 B.n421 VSUBS 0.00835f
C660 B.n422 VSUBS 0.00835f
C661 B.n423 VSUBS 0.00835f
C662 B.n424 VSUBS 0.00835f
C663 B.n425 VSUBS 0.00835f
C664 B.n426 VSUBS 0.021056f
C665 B.n427 VSUBS 0.020138f
C666 B.n428 VSUBS 0.020877f
C667 B.n429 VSUBS 0.00835f
C668 B.n430 VSUBS 0.00835f
C669 B.n431 VSUBS 0.00835f
C670 B.n432 VSUBS 0.00835f
C671 B.n433 VSUBS 0.00835f
C672 B.n434 VSUBS 0.00835f
C673 B.n435 VSUBS 0.00835f
C674 B.n436 VSUBS 0.00835f
C675 B.n437 VSUBS 0.00835f
C676 B.n438 VSUBS 0.00835f
C677 B.n439 VSUBS 0.00835f
C678 B.n440 VSUBS 0.00835f
C679 B.n441 VSUBS 0.00835f
C680 B.n442 VSUBS 0.00835f
C681 B.n443 VSUBS 0.00835f
C682 B.n444 VSUBS 0.00835f
C683 B.n445 VSUBS 0.00835f
C684 B.n446 VSUBS 0.00835f
C685 B.n447 VSUBS 0.00835f
C686 B.n448 VSUBS 0.00835f
C687 B.n449 VSUBS 0.00835f
C688 B.n450 VSUBS 0.00835f
C689 B.n451 VSUBS 0.00835f
C690 B.n452 VSUBS 0.00835f
C691 B.n453 VSUBS 0.00835f
C692 B.n454 VSUBS 0.00835f
C693 B.n455 VSUBS 0.00835f
C694 B.n456 VSUBS 0.00835f
C695 B.n457 VSUBS 0.00835f
C696 B.n458 VSUBS 0.00835f
C697 B.n459 VSUBS 0.00835f
C698 B.n460 VSUBS 0.00835f
C699 B.n461 VSUBS 0.00835f
C700 B.n462 VSUBS 0.00835f
C701 B.n463 VSUBS 0.00835f
C702 B.n464 VSUBS 0.00835f
C703 B.n465 VSUBS 0.00835f
C704 B.n466 VSUBS 0.00835f
C705 B.n467 VSUBS 0.00835f
C706 B.n468 VSUBS 0.00835f
C707 B.n469 VSUBS 0.00835f
C708 B.n470 VSUBS 0.00835f
C709 B.n471 VSUBS 0.00835f
C710 B.n472 VSUBS 0.00835f
C711 B.n473 VSUBS 0.00835f
C712 B.n474 VSUBS 0.00835f
C713 B.n475 VSUBS 0.00835f
C714 B.n476 VSUBS 0.00835f
C715 B.n477 VSUBS 0.00835f
C716 B.n478 VSUBS 0.00835f
C717 B.n479 VSUBS 0.00835f
C718 B.n480 VSUBS 0.00835f
C719 B.n481 VSUBS 0.00835f
C720 B.n482 VSUBS 0.00835f
C721 B.n483 VSUBS 0.00835f
C722 B.n484 VSUBS 0.00835f
C723 B.n485 VSUBS 0.00835f
C724 B.n486 VSUBS 0.00835f
C725 B.n487 VSUBS 0.00835f
C726 B.n488 VSUBS 0.00835f
C727 B.n489 VSUBS 0.00835f
C728 B.n490 VSUBS 0.00835f
C729 B.n491 VSUBS 0.00835f
C730 B.n492 VSUBS 0.00835f
C731 B.n493 VSUBS 0.00835f
C732 B.n494 VSUBS 0.00835f
C733 B.n495 VSUBS 0.00835f
C734 B.n496 VSUBS 0.00835f
C735 B.n497 VSUBS 0.00835f
C736 B.n498 VSUBS 0.00835f
C737 B.n499 VSUBS 0.00835f
C738 B.n500 VSUBS 0.00835f
C739 B.n501 VSUBS 0.00835f
C740 B.n502 VSUBS 0.00835f
C741 B.n503 VSUBS 0.00835f
C742 B.n504 VSUBS 0.00835f
C743 B.n505 VSUBS 0.00835f
C744 B.n506 VSUBS 0.00835f
C745 B.n507 VSUBS 0.00835f
C746 B.n508 VSUBS 0.00835f
C747 B.n509 VSUBS 0.00835f
C748 B.n510 VSUBS 0.00835f
C749 B.n511 VSUBS 0.00835f
C750 B.n512 VSUBS 0.00835f
C751 B.n513 VSUBS 0.00835f
C752 B.n514 VSUBS 0.00835f
C753 B.n515 VSUBS 0.00835f
C754 B.n516 VSUBS 0.00835f
C755 B.n517 VSUBS 0.00835f
C756 B.n518 VSUBS 0.00835f
C757 B.n519 VSUBS 0.00835f
C758 B.n520 VSUBS 0.00835f
C759 B.n521 VSUBS 0.00835f
C760 B.n522 VSUBS 0.00835f
C761 B.n523 VSUBS 0.00835f
C762 B.n524 VSUBS 0.00835f
C763 B.n525 VSUBS 0.00835f
C764 B.n526 VSUBS 0.00835f
C765 B.n527 VSUBS 0.00835f
C766 B.n528 VSUBS 0.00835f
C767 B.n529 VSUBS 0.00835f
C768 B.n530 VSUBS 0.00835f
C769 B.n531 VSUBS 0.00835f
C770 B.n532 VSUBS 0.00835f
C771 B.n533 VSUBS 0.00835f
C772 B.n534 VSUBS 0.00835f
C773 B.n535 VSUBS 0.00835f
C774 B.n536 VSUBS 0.00835f
C775 B.n537 VSUBS 0.00835f
C776 B.n538 VSUBS 0.00835f
C777 B.n539 VSUBS 0.00835f
C778 B.n540 VSUBS 0.00835f
C779 B.n541 VSUBS 0.00835f
C780 B.n542 VSUBS 0.00835f
C781 B.n543 VSUBS 0.00835f
C782 B.n544 VSUBS 0.00835f
C783 B.n545 VSUBS 0.00835f
C784 B.n546 VSUBS 0.00835f
C785 B.n547 VSUBS 0.00835f
C786 B.n548 VSUBS 0.00835f
C787 B.n549 VSUBS 0.00835f
C788 B.n550 VSUBS 0.00835f
C789 B.n551 VSUBS 0.00835f
C790 B.n552 VSUBS 0.00835f
C791 B.n553 VSUBS 0.00835f
C792 B.n554 VSUBS 0.00835f
C793 B.n555 VSUBS 0.00835f
C794 B.n556 VSUBS 0.00835f
C795 B.n557 VSUBS 0.00835f
C796 B.n558 VSUBS 0.00835f
C797 B.n559 VSUBS 0.00835f
C798 B.n560 VSUBS 0.00835f
C799 B.n561 VSUBS 0.00835f
C800 B.n562 VSUBS 0.00835f
C801 B.n563 VSUBS 0.00835f
C802 B.n564 VSUBS 0.00835f
C803 B.n565 VSUBS 0.00835f
C804 B.n566 VSUBS 0.00835f
C805 B.n567 VSUBS 0.019959f
C806 B.n568 VSUBS 0.019959f
C807 B.n569 VSUBS 0.021056f
C808 B.n570 VSUBS 0.00835f
C809 B.n571 VSUBS 0.00835f
C810 B.n572 VSUBS 0.00835f
C811 B.n573 VSUBS 0.00835f
C812 B.n574 VSUBS 0.00835f
C813 B.n575 VSUBS 0.00835f
C814 B.n576 VSUBS 0.00835f
C815 B.n577 VSUBS 0.00835f
C816 B.n578 VSUBS 0.00835f
C817 B.n579 VSUBS 0.00835f
C818 B.n580 VSUBS 0.00835f
C819 B.n581 VSUBS 0.00835f
C820 B.n582 VSUBS 0.00835f
C821 B.n583 VSUBS 0.00835f
C822 B.n584 VSUBS 0.00835f
C823 B.n585 VSUBS 0.00835f
C824 B.n586 VSUBS 0.00835f
C825 B.n587 VSUBS 0.00835f
C826 B.n588 VSUBS 0.00835f
C827 B.n589 VSUBS 0.00835f
C828 B.n590 VSUBS 0.00835f
C829 B.n591 VSUBS 0.00835f
C830 B.n592 VSUBS 0.00835f
C831 B.n593 VSUBS 0.00835f
C832 B.n594 VSUBS 0.00835f
C833 B.n595 VSUBS 0.00835f
C834 B.n596 VSUBS 0.00835f
C835 B.n597 VSUBS 0.00835f
C836 B.n598 VSUBS 0.00835f
C837 B.n599 VSUBS 0.00835f
C838 B.n600 VSUBS 0.00835f
C839 B.n601 VSUBS 0.00835f
C840 B.n602 VSUBS 0.00835f
C841 B.n603 VSUBS 0.00835f
C842 B.n604 VSUBS 0.00835f
C843 B.n605 VSUBS 0.00835f
C844 B.n606 VSUBS 0.00835f
C845 B.n607 VSUBS 0.00835f
C846 B.n608 VSUBS 0.00835f
C847 B.n609 VSUBS 0.00835f
C848 B.n610 VSUBS 0.00835f
C849 B.n611 VSUBS 0.00835f
C850 B.n612 VSUBS 0.00835f
C851 B.n613 VSUBS 0.00835f
C852 B.n614 VSUBS 0.00835f
C853 B.n615 VSUBS 0.00835f
C854 B.n616 VSUBS 0.00835f
C855 B.n617 VSUBS 0.00835f
C856 B.n618 VSUBS 0.00835f
C857 B.n619 VSUBS 0.00835f
C858 B.n620 VSUBS 0.00835f
C859 B.n621 VSUBS 0.00835f
C860 B.n622 VSUBS 0.00835f
C861 B.n623 VSUBS 0.00835f
C862 B.n624 VSUBS 0.00835f
C863 B.n625 VSUBS 0.00835f
C864 B.n626 VSUBS 0.00835f
C865 B.n627 VSUBS 0.00835f
C866 B.n628 VSUBS 0.00835f
C867 B.n629 VSUBS 0.00835f
C868 B.n630 VSUBS 0.00835f
C869 B.n631 VSUBS 0.00835f
C870 B.n632 VSUBS 0.00835f
C871 B.n633 VSUBS 0.00835f
C872 B.n634 VSUBS 0.00835f
C873 B.n635 VSUBS 0.00835f
C874 B.n636 VSUBS 0.00835f
C875 B.n637 VSUBS 0.007859f
C876 B.n638 VSUBS 0.019347f
C877 B.n639 VSUBS 0.004666f
C878 B.n640 VSUBS 0.00835f
C879 B.n641 VSUBS 0.00835f
C880 B.n642 VSUBS 0.00835f
C881 B.n643 VSUBS 0.00835f
C882 B.n644 VSUBS 0.00835f
C883 B.n645 VSUBS 0.00835f
C884 B.n646 VSUBS 0.00835f
C885 B.n647 VSUBS 0.00835f
C886 B.n648 VSUBS 0.00835f
C887 B.n649 VSUBS 0.00835f
C888 B.n650 VSUBS 0.00835f
C889 B.n651 VSUBS 0.00835f
C890 B.n652 VSUBS 0.004666f
C891 B.n653 VSUBS 0.00835f
C892 B.n654 VSUBS 0.00835f
C893 B.n655 VSUBS 0.007859f
C894 B.n656 VSUBS 0.00835f
C895 B.n657 VSUBS 0.00835f
C896 B.n658 VSUBS 0.00835f
C897 B.n659 VSUBS 0.00835f
C898 B.n660 VSUBS 0.00835f
C899 B.n661 VSUBS 0.00835f
C900 B.n662 VSUBS 0.00835f
C901 B.n663 VSUBS 0.00835f
C902 B.n664 VSUBS 0.00835f
C903 B.n665 VSUBS 0.00835f
C904 B.n666 VSUBS 0.00835f
C905 B.n667 VSUBS 0.00835f
C906 B.n668 VSUBS 0.00835f
C907 B.n669 VSUBS 0.00835f
C908 B.n670 VSUBS 0.00835f
C909 B.n671 VSUBS 0.00835f
C910 B.n672 VSUBS 0.00835f
C911 B.n673 VSUBS 0.00835f
C912 B.n674 VSUBS 0.00835f
C913 B.n675 VSUBS 0.00835f
C914 B.n676 VSUBS 0.00835f
C915 B.n677 VSUBS 0.00835f
C916 B.n678 VSUBS 0.00835f
C917 B.n679 VSUBS 0.00835f
C918 B.n680 VSUBS 0.00835f
C919 B.n681 VSUBS 0.00835f
C920 B.n682 VSUBS 0.00835f
C921 B.n683 VSUBS 0.00835f
C922 B.n684 VSUBS 0.00835f
C923 B.n685 VSUBS 0.00835f
C924 B.n686 VSUBS 0.00835f
C925 B.n687 VSUBS 0.00835f
C926 B.n688 VSUBS 0.00835f
C927 B.n689 VSUBS 0.00835f
C928 B.n690 VSUBS 0.00835f
C929 B.n691 VSUBS 0.00835f
C930 B.n692 VSUBS 0.00835f
C931 B.n693 VSUBS 0.00835f
C932 B.n694 VSUBS 0.00835f
C933 B.n695 VSUBS 0.00835f
C934 B.n696 VSUBS 0.00835f
C935 B.n697 VSUBS 0.00835f
C936 B.n698 VSUBS 0.00835f
C937 B.n699 VSUBS 0.00835f
C938 B.n700 VSUBS 0.00835f
C939 B.n701 VSUBS 0.00835f
C940 B.n702 VSUBS 0.00835f
C941 B.n703 VSUBS 0.00835f
C942 B.n704 VSUBS 0.00835f
C943 B.n705 VSUBS 0.00835f
C944 B.n706 VSUBS 0.00835f
C945 B.n707 VSUBS 0.00835f
C946 B.n708 VSUBS 0.00835f
C947 B.n709 VSUBS 0.00835f
C948 B.n710 VSUBS 0.00835f
C949 B.n711 VSUBS 0.00835f
C950 B.n712 VSUBS 0.00835f
C951 B.n713 VSUBS 0.00835f
C952 B.n714 VSUBS 0.00835f
C953 B.n715 VSUBS 0.00835f
C954 B.n716 VSUBS 0.00835f
C955 B.n717 VSUBS 0.00835f
C956 B.n718 VSUBS 0.00835f
C957 B.n719 VSUBS 0.00835f
C958 B.n720 VSUBS 0.00835f
C959 B.n721 VSUBS 0.00835f
C960 B.n722 VSUBS 0.021056f
C961 B.n723 VSUBS 0.019959f
C962 B.n724 VSUBS 0.019959f
C963 B.n725 VSUBS 0.00835f
C964 B.n726 VSUBS 0.00835f
C965 B.n727 VSUBS 0.00835f
C966 B.n728 VSUBS 0.00835f
C967 B.n729 VSUBS 0.00835f
C968 B.n730 VSUBS 0.00835f
C969 B.n731 VSUBS 0.00835f
C970 B.n732 VSUBS 0.00835f
C971 B.n733 VSUBS 0.00835f
C972 B.n734 VSUBS 0.00835f
C973 B.n735 VSUBS 0.00835f
C974 B.n736 VSUBS 0.00835f
C975 B.n737 VSUBS 0.00835f
C976 B.n738 VSUBS 0.00835f
C977 B.n739 VSUBS 0.00835f
C978 B.n740 VSUBS 0.00835f
C979 B.n741 VSUBS 0.00835f
C980 B.n742 VSUBS 0.00835f
C981 B.n743 VSUBS 0.00835f
C982 B.n744 VSUBS 0.00835f
C983 B.n745 VSUBS 0.00835f
C984 B.n746 VSUBS 0.00835f
C985 B.n747 VSUBS 0.00835f
C986 B.n748 VSUBS 0.00835f
C987 B.n749 VSUBS 0.00835f
C988 B.n750 VSUBS 0.00835f
C989 B.n751 VSUBS 0.00835f
C990 B.n752 VSUBS 0.00835f
C991 B.n753 VSUBS 0.00835f
C992 B.n754 VSUBS 0.00835f
C993 B.n755 VSUBS 0.00835f
C994 B.n756 VSUBS 0.00835f
C995 B.n757 VSUBS 0.00835f
C996 B.n758 VSUBS 0.00835f
C997 B.n759 VSUBS 0.00835f
C998 B.n760 VSUBS 0.00835f
C999 B.n761 VSUBS 0.00835f
C1000 B.n762 VSUBS 0.00835f
C1001 B.n763 VSUBS 0.00835f
C1002 B.n764 VSUBS 0.00835f
C1003 B.n765 VSUBS 0.00835f
C1004 B.n766 VSUBS 0.00835f
C1005 B.n767 VSUBS 0.00835f
C1006 B.n768 VSUBS 0.00835f
C1007 B.n769 VSUBS 0.00835f
C1008 B.n770 VSUBS 0.00835f
C1009 B.n771 VSUBS 0.00835f
C1010 B.n772 VSUBS 0.00835f
C1011 B.n773 VSUBS 0.00835f
C1012 B.n774 VSUBS 0.00835f
C1013 B.n775 VSUBS 0.00835f
C1014 B.n776 VSUBS 0.00835f
C1015 B.n777 VSUBS 0.00835f
C1016 B.n778 VSUBS 0.00835f
C1017 B.n779 VSUBS 0.00835f
C1018 B.n780 VSUBS 0.00835f
C1019 B.n781 VSUBS 0.00835f
C1020 B.n782 VSUBS 0.00835f
C1021 B.n783 VSUBS 0.00835f
C1022 B.n784 VSUBS 0.00835f
C1023 B.n785 VSUBS 0.00835f
C1024 B.n786 VSUBS 0.00835f
C1025 B.n787 VSUBS 0.00835f
C1026 B.n788 VSUBS 0.00835f
C1027 B.n789 VSUBS 0.00835f
C1028 B.n790 VSUBS 0.00835f
C1029 B.n791 VSUBS 0.010897f
C1030 B.n792 VSUBS 0.011608f
C1031 B.n793 VSUBS 0.023083f
C1032 VTAIL.t3 VSUBS 0.30963f
C1033 VTAIL.t1 VSUBS 0.30963f
C1034 VTAIL.n0 VSUBS 2.30299f
C1035 VTAIL.n1 VSUBS 0.923635f
C1036 VTAIL.n2 VSUBS 0.032806f
C1037 VTAIL.n3 VSUBS 0.028853f
C1038 VTAIL.n4 VSUBS 0.015504f
C1039 VTAIL.n5 VSUBS 0.036647f
C1040 VTAIL.n6 VSUBS 0.016416f
C1041 VTAIL.n7 VSUBS 0.028853f
C1042 VTAIL.n8 VSUBS 0.015504f
C1043 VTAIL.n9 VSUBS 0.036647f
C1044 VTAIL.n10 VSUBS 0.016416f
C1045 VTAIL.n11 VSUBS 0.028853f
C1046 VTAIL.n12 VSUBS 0.015504f
C1047 VTAIL.n13 VSUBS 0.036647f
C1048 VTAIL.n14 VSUBS 0.01596f
C1049 VTAIL.n15 VSUBS 0.028853f
C1050 VTAIL.n16 VSUBS 0.016416f
C1051 VTAIL.n17 VSUBS 0.036647f
C1052 VTAIL.n18 VSUBS 0.016416f
C1053 VTAIL.n19 VSUBS 0.028853f
C1054 VTAIL.n20 VSUBS 0.015504f
C1055 VTAIL.n21 VSUBS 0.036647f
C1056 VTAIL.n22 VSUBS 0.016416f
C1057 VTAIL.n23 VSUBS 1.61739f
C1058 VTAIL.n24 VSUBS 0.015504f
C1059 VTAIL.t7 VSUBS 0.079121f
C1060 VTAIL.n25 VSUBS 0.247844f
C1061 VTAIL.n26 VSUBS 0.027568f
C1062 VTAIL.n27 VSUBS 0.027485f
C1063 VTAIL.n28 VSUBS 0.036647f
C1064 VTAIL.n29 VSUBS 0.016416f
C1065 VTAIL.n30 VSUBS 0.015504f
C1066 VTAIL.n31 VSUBS 0.028853f
C1067 VTAIL.n32 VSUBS 0.028853f
C1068 VTAIL.n33 VSUBS 0.015504f
C1069 VTAIL.n34 VSUBS 0.016416f
C1070 VTAIL.n35 VSUBS 0.036647f
C1071 VTAIL.n36 VSUBS 0.036647f
C1072 VTAIL.n37 VSUBS 0.016416f
C1073 VTAIL.n38 VSUBS 0.015504f
C1074 VTAIL.n39 VSUBS 0.028853f
C1075 VTAIL.n40 VSUBS 0.028853f
C1076 VTAIL.n41 VSUBS 0.015504f
C1077 VTAIL.n42 VSUBS 0.015504f
C1078 VTAIL.n43 VSUBS 0.016416f
C1079 VTAIL.n44 VSUBS 0.036647f
C1080 VTAIL.n45 VSUBS 0.036647f
C1081 VTAIL.n46 VSUBS 0.036647f
C1082 VTAIL.n47 VSUBS 0.01596f
C1083 VTAIL.n48 VSUBS 0.015504f
C1084 VTAIL.n49 VSUBS 0.028853f
C1085 VTAIL.n50 VSUBS 0.028853f
C1086 VTAIL.n51 VSUBS 0.015504f
C1087 VTAIL.n52 VSUBS 0.016416f
C1088 VTAIL.n53 VSUBS 0.036647f
C1089 VTAIL.n54 VSUBS 0.036647f
C1090 VTAIL.n55 VSUBS 0.016416f
C1091 VTAIL.n56 VSUBS 0.015504f
C1092 VTAIL.n57 VSUBS 0.028853f
C1093 VTAIL.n58 VSUBS 0.028853f
C1094 VTAIL.n59 VSUBS 0.015504f
C1095 VTAIL.n60 VSUBS 0.016416f
C1096 VTAIL.n61 VSUBS 0.036647f
C1097 VTAIL.n62 VSUBS 0.036647f
C1098 VTAIL.n63 VSUBS 0.016416f
C1099 VTAIL.n64 VSUBS 0.015504f
C1100 VTAIL.n65 VSUBS 0.028853f
C1101 VTAIL.n66 VSUBS 0.028853f
C1102 VTAIL.n67 VSUBS 0.015504f
C1103 VTAIL.n68 VSUBS 0.016416f
C1104 VTAIL.n69 VSUBS 0.036647f
C1105 VTAIL.n70 VSUBS 0.092473f
C1106 VTAIL.n71 VSUBS 0.016416f
C1107 VTAIL.n72 VSUBS 0.015504f
C1108 VTAIL.n73 VSUBS 0.067481f
C1109 VTAIL.n74 VSUBS 0.046694f
C1110 VTAIL.n75 VSUBS 0.463091f
C1111 VTAIL.t8 VSUBS 0.30963f
C1112 VTAIL.t9 VSUBS 0.30963f
C1113 VTAIL.n76 VSUBS 2.30299f
C1114 VTAIL.n77 VSUBS 2.94636f
C1115 VTAIL.t2 VSUBS 0.30963f
C1116 VTAIL.t10 VSUBS 0.30963f
C1117 VTAIL.n78 VSUBS 2.30301f
C1118 VTAIL.n79 VSUBS 2.94634f
C1119 VTAIL.n80 VSUBS 0.032806f
C1120 VTAIL.n81 VSUBS 0.028853f
C1121 VTAIL.n82 VSUBS 0.015504f
C1122 VTAIL.n83 VSUBS 0.036647f
C1123 VTAIL.n84 VSUBS 0.016416f
C1124 VTAIL.n85 VSUBS 0.028853f
C1125 VTAIL.n86 VSUBS 0.015504f
C1126 VTAIL.n87 VSUBS 0.036647f
C1127 VTAIL.n88 VSUBS 0.016416f
C1128 VTAIL.n89 VSUBS 0.028853f
C1129 VTAIL.n90 VSUBS 0.015504f
C1130 VTAIL.n91 VSUBS 0.036647f
C1131 VTAIL.n92 VSUBS 0.01596f
C1132 VTAIL.n93 VSUBS 0.028853f
C1133 VTAIL.n94 VSUBS 0.01596f
C1134 VTAIL.n95 VSUBS 0.015504f
C1135 VTAIL.n96 VSUBS 0.036647f
C1136 VTAIL.n97 VSUBS 0.036647f
C1137 VTAIL.n98 VSUBS 0.016416f
C1138 VTAIL.n99 VSUBS 0.028853f
C1139 VTAIL.n100 VSUBS 0.015504f
C1140 VTAIL.n101 VSUBS 0.036647f
C1141 VTAIL.n102 VSUBS 0.016416f
C1142 VTAIL.n103 VSUBS 1.61739f
C1143 VTAIL.n104 VSUBS 0.015504f
C1144 VTAIL.t11 VSUBS 0.079121f
C1145 VTAIL.n105 VSUBS 0.247844f
C1146 VTAIL.n106 VSUBS 0.027568f
C1147 VTAIL.n107 VSUBS 0.027485f
C1148 VTAIL.n108 VSUBS 0.036647f
C1149 VTAIL.n109 VSUBS 0.016416f
C1150 VTAIL.n110 VSUBS 0.015504f
C1151 VTAIL.n111 VSUBS 0.028853f
C1152 VTAIL.n112 VSUBS 0.028853f
C1153 VTAIL.n113 VSUBS 0.015504f
C1154 VTAIL.n114 VSUBS 0.016416f
C1155 VTAIL.n115 VSUBS 0.036647f
C1156 VTAIL.n116 VSUBS 0.036647f
C1157 VTAIL.n117 VSUBS 0.016416f
C1158 VTAIL.n118 VSUBS 0.015504f
C1159 VTAIL.n119 VSUBS 0.028853f
C1160 VTAIL.n120 VSUBS 0.028853f
C1161 VTAIL.n121 VSUBS 0.015504f
C1162 VTAIL.n122 VSUBS 0.016416f
C1163 VTAIL.n123 VSUBS 0.036647f
C1164 VTAIL.n124 VSUBS 0.036647f
C1165 VTAIL.n125 VSUBS 0.016416f
C1166 VTAIL.n126 VSUBS 0.015504f
C1167 VTAIL.n127 VSUBS 0.028853f
C1168 VTAIL.n128 VSUBS 0.028853f
C1169 VTAIL.n129 VSUBS 0.015504f
C1170 VTAIL.n130 VSUBS 0.016416f
C1171 VTAIL.n131 VSUBS 0.036647f
C1172 VTAIL.n132 VSUBS 0.036647f
C1173 VTAIL.n133 VSUBS 0.016416f
C1174 VTAIL.n134 VSUBS 0.015504f
C1175 VTAIL.n135 VSUBS 0.028853f
C1176 VTAIL.n136 VSUBS 0.028853f
C1177 VTAIL.n137 VSUBS 0.015504f
C1178 VTAIL.n138 VSUBS 0.016416f
C1179 VTAIL.n139 VSUBS 0.036647f
C1180 VTAIL.n140 VSUBS 0.036647f
C1181 VTAIL.n141 VSUBS 0.016416f
C1182 VTAIL.n142 VSUBS 0.015504f
C1183 VTAIL.n143 VSUBS 0.028853f
C1184 VTAIL.n144 VSUBS 0.028853f
C1185 VTAIL.n145 VSUBS 0.015504f
C1186 VTAIL.n146 VSUBS 0.016416f
C1187 VTAIL.n147 VSUBS 0.036647f
C1188 VTAIL.n148 VSUBS 0.092473f
C1189 VTAIL.n149 VSUBS 0.016416f
C1190 VTAIL.n150 VSUBS 0.015504f
C1191 VTAIL.n151 VSUBS 0.067481f
C1192 VTAIL.n152 VSUBS 0.046694f
C1193 VTAIL.n153 VSUBS 0.463091f
C1194 VTAIL.t4 VSUBS 0.30963f
C1195 VTAIL.t5 VSUBS 0.30963f
C1196 VTAIL.n154 VSUBS 2.30301f
C1197 VTAIL.n155 VSUBS 1.11537f
C1198 VTAIL.n156 VSUBS 0.032806f
C1199 VTAIL.n157 VSUBS 0.028853f
C1200 VTAIL.n158 VSUBS 0.015504f
C1201 VTAIL.n159 VSUBS 0.036647f
C1202 VTAIL.n160 VSUBS 0.016416f
C1203 VTAIL.n161 VSUBS 0.028853f
C1204 VTAIL.n162 VSUBS 0.015504f
C1205 VTAIL.n163 VSUBS 0.036647f
C1206 VTAIL.n164 VSUBS 0.016416f
C1207 VTAIL.n165 VSUBS 0.028853f
C1208 VTAIL.n166 VSUBS 0.015504f
C1209 VTAIL.n167 VSUBS 0.036647f
C1210 VTAIL.n168 VSUBS 0.01596f
C1211 VTAIL.n169 VSUBS 0.028853f
C1212 VTAIL.n170 VSUBS 0.01596f
C1213 VTAIL.n171 VSUBS 0.015504f
C1214 VTAIL.n172 VSUBS 0.036647f
C1215 VTAIL.n173 VSUBS 0.036647f
C1216 VTAIL.n174 VSUBS 0.016416f
C1217 VTAIL.n175 VSUBS 0.028853f
C1218 VTAIL.n176 VSUBS 0.015504f
C1219 VTAIL.n177 VSUBS 0.036647f
C1220 VTAIL.n178 VSUBS 0.016416f
C1221 VTAIL.n179 VSUBS 1.61739f
C1222 VTAIL.n180 VSUBS 0.015504f
C1223 VTAIL.t6 VSUBS 0.079121f
C1224 VTAIL.n181 VSUBS 0.247844f
C1225 VTAIL.n182 VSUBS 0.027568f
C1226 VTAIL.n183 VSUBS 0.027485f
C1227 VTAIL.n184 VSUBS 0.036647f
C1228 VTAIL.n185 VSUBS 0.016416f
C1229 VTAIL.n186 VSUBS 0.015504f
C1230 VTAIL.n187 VSUBS 0.028853f
C1231 VTAIL.n188 VSUBS 0.028853f
C1232 VTAIL.n189 VSUBS 0.015504f
C1233 VTAIL.n190 VSUBS 0.016416f
C1234 VTAIL.n191 VSUBS 0.036647f
C1235 VTAIL.n192 VSUBS 0.036647f
C1236 VTAIL.n193 VSUBS 0.016416f
C1237 VTAIL.n194 VSUBS 0.015504f
C1238 VTAIL.n195 VSUBS 0.028853f
C1239 VTAIL.n196 VSUBS 0.028853f
C1240 VTAIL.n197 VSUBS 0.015504f
C1241 VTAIL.n198 VSUBS 0.016416f
C1242 VTAIL.n199 VSUBS 0.036647f
C1243 VTAIL.n200 VSUBS 0.036647f
C1244 VTAIL.n201 VSUBS 0.016416f
C1245 VTAIL.n202 VSUBS 0.015504f
C1246 VTAIL.n203 VSUBS 0.028853f
C1247 VTAIL.n204 VSUBS 0.028853f
C1248 VTAIL.n205 VSUBS 0.015504f
C1249 VTAIL.n206 VSUBS 0.016416f
C1250 VTAIL.n207 VSUBS 0.036647f
C1251 VTAIL.n208 VSUBS 0.036647f
C1252 VTAIL.n209 VSUBS 0.016416f
C1253 VTAIL.n210 VSUBS 0.015504f
C1254 VTAIL.n211 VSUBS 0.028853f
C1255 VTAIL.n212 VSUBS 0.028853f
C1256 VTAIL.n213 VSUBS 0.015504f
C1257 VTAIL.n214 VSUBS 0.016416f
C1258 VTAIL.n215 VSUBS 0.036647f
C1259 VTAIL.n216 VSUBS 0.036647f
C1260 VTAIL.n217 VSUBS 0.016416f
C1261 VTAIL.n218 VSUBS 0.015504f
C1262 VTAIL.n219 VSUBS 0.028853f
C1263 VTAIL.n220 VSUBS 0.028853f
C1264 VTAIL.n221 VSUBS 0.015504f
C1265 VTAIL.n222 VSUBS 0.016416f
C1266 VTAIL.n223 VSUBS 0.036647f
C1267 VTAIL.n224 VSUBS 0.092473f
C1268 VTAIL.n225 VSUBS 0.016416f
C1269 VTAIL.n226 VSUBS 0.015504f
C1270 VTAIL.n227 VSUBS 0.067481f
C1271 VTAIL.n228 VSUBS 0.046694f
C1272 VTAIL.n229 VSUBS 2.03118f
C1273 VTAIL.n230 VSUBS 0.032806f
C1274 VTAIL.n231 VSUBS 0.028853f
C1275 VTAIL.n232 VSUBS 0.015504f
C1276 VTAIL.n233 VSUBS 0.036647f
C1277 VTAIL.n234 VSUBS 0.016416f
C1278 VTAIL.n235 VSUBS 0.028853f
C1279 VTAIL.n236 VSUBS 0.015504f
C1280 VTAIL.n237 VSUBS 0.036647f
C1281 VTAIL.n238 VSUBS 0.016416f
C1282 VTAIL.n239 VSUBS 0.028853f
C1283 VTAIL.n240 VSUBS 0.015504f
C1284 VTAIL.n241 VSUBS 0.036647f
C1285 VTAIL.n242 VSUBS 0.01596f
C1286 VTAIL.n243 VSUBS 0.028853f
C1287 VTAIL.n244 VSUBS 0.016416f
C1288 VTAIL.n245 VSUBS 0.036647f
C1289 VTAIL.n246 VSUBS 0.016416f
C1290 VTAIL.n247 VSUBS 0.028853f
C1291 VTAIL.n248 VSUBS 0.015504f
C1292 VTAIL.n249 VSUBS 0.036647f
C1293 VTAIL.n250 VSUBS 0.016416f
C1294 VTAIL.n251 VSUBS 1.61739f
C1295 VTAIL.n252 VSUBS 0.015504f
C1296 VTAIL.t0 VSUBS 0.079121f
C1297 VTAIL.n253 VSUBS 0.247844f
C1298 VTAIL.n254 VSUBS 0.027568f
C1299 VTAIL.n255 VSUBS 0.027485f
C1300 VTAIL.n256 VSUBS 0.036647f
C1301 VTAIL.n257 VSUBS 0.016416f
C1302 VTAIL.n258 VSUBS 0.015504f
C1303 VTAIL.n259 VSUBS 0.028853f
C1304 VTAIL.n260 VSUBS 0.028853f
C1305 VTAIL.n261 VSUBS 0.015504f
C1306 VTAIL.n262 VSUBS 0.016416f
C1307 VTAIL.n263 VSUBS 0.036647f
C1308 VTAIL.n264 VSUBS 0.036647f
C1309 VTAIL.n265 VSUBS 0.016416f
C1310 VTAIL.n266 VSUBS 0.015504f
C1311 VTAIL.n267 VSUBS 0.028853f
C1312 VTAIL.n268 VSUBS 0.028853f
C1313 VTAIL.n269 VSUBS 0.015504f
C1314 VTAIL.n270 VSUBS 0.015504f
C1315 VTAIL.n271 VSUBS 0.016416f
C1316 VTAIL.n272 VSUBS 0.036647f
C1317 VTAIL.n273 VSUBS 0.036647f
C1318 VTAIL.n274 VSUBS 0.036647f
C1319 VTAIL.n275 VSUBS 0.01596f
C1320 VTAIL.n276 VSUBS 0.015504f
C1321 VTAIL.n277 VSUBS 0.028853f
C1322 VTAIL.n278 VSUBS 0.028853f
C1323 VTAIL.n279 VSUBS 0.015504f
C1324 VTAIL.n280 VSUBS 0.016416f
C1325 VTAIL.n281 VSUBS 0.036647f
C1326 VTAIL.n282 VSUBS 0.036647f
C1327 VTAIL.n283 VSUBS 0.016416f
C1328 VTAIL.n284 VSUBS 0.015504f
C1329 VTAIL.n285 VSUBS 0.028853f
C1330 VTAIL.n286 VSUBS 0.028853f
C1331 VTAIL.n287 VSUBS 0.015504f
C1332 VTAIL.n288 VSUBS 0.016416f
C1333 VTAIL.n289 VSUBS 0.036647f
C1334 VTAIL.n290 VSUBS 0.036647f
C1335 VTAIL.n291 VSUBS 0.016416f
C1336 VTAIL.n292 VSUBS 0.015504f
C1337 VTAIL.n293 VSUBS 0.028853f
C1338 VTAIL.n294 VSUBS 0.028853f
C1339 VTAIL.n295 VSUBS 0.015504f
C1340 VTAIL.n296 VSUBS 0.016416f
C1341 VTAIL.n297 VSUBS 0.036647f
C1342 VTAIL.n298 VSUBS 0.092473f
C1343 VTAIL.n299 VSUBS 0.016416f
C1344 VTAIL.n300 VSUBS 0.015504f
C1345 VTAIL.n301 VSUBS 0.067481f
C1346 VTAIL.n302 VSUBS 0.046694f
C1347 VTAIL.n303 VSUBS 1.96005f
C1348 VDD1.n0 VSUBS 0.031783f
C1349 VDD1.n1 VSUBS 0.027953f
C1350 VDD1.n2 VSUBS 0.015021f
C1351 VDD1.n3 VSUBS 0.035504f
C1352 VDD1.n4 VSUBS 0.015904f
C1353 VDD1.n5 VSUBS 0.027953f
C1354 VDD1.n6 VSUBS 0.015021f
C1355 VDD1.n7 VSUBS 0.035504f
C1356 VDD1.n8 VSUBS 0.015904f
C1357 VDD1.n9 VSUBS 0.027953f
C1358 VDD1.n10 VSUBS 0.015021f
C1359 VDD1.n11 VSUBS 0.035504f
C1360 VDD1.n12 VSUBS 0.015463f
C1361 VDD1.n13 VSUBS 0.027953f
C1362 VDD1.n14 VSUBS 0.015463f
C1363 VDD1.n15 VSUBS 0.015021f
C1364 VDD1.n16 VSUBS 0.035504f
C1365 VDD1.n17 VSUBS 0.035504f
C1366 VDD1.n18 VSUBS 0.015904f
C1367 VDD1.n19 VSUBS 0.027953f
C1368 VDD1.n20 VSUBS 0.015021f
C1369 VDD1.n21 VSUBS 0.035504f
C1370 VDD1.n22 VSUBS 0.015904f
C1371 VDD1.n23 VSUBS 1.56696f
C1372 VDD1.n24 VSUBS 0.015021f
C1373 VDD1.t5 VSUBS 0.076654f
C1374 VDD1.n25 VSUBS 0.240117f
C1375 VDD1.n26 VSUBS 0.026708f
C1376 VDD1.n27 VSUBS 0.026628f
C1377 VDD1.n28 VSUBS 0.035504f
C1378 VDD1.n29 VSUBS 0.015904f
C1379 VDD1.n30 VSUBS 0.015021f
C1380 VDD1.n31 VSUBS 0.027953f
C1381 VDD1.n32 VSUBS 0.027953f
C1382 VDD1.n33 VSUBS 0.015021f
C1383 VDD1.n34 VSUBS 0.015904f
C1384 VDD1.n35 VSUBS 0.035504f
C1385 VDD1.n36 VSUBS 0.035504f
C1386 VDD1.n37 VSUBS 0.015904f
C1387 VDD1.n38 VSUBS 0.015021f
C1388 VDD1.n39 VSUBS 0.027953f
C1389 VDD1.n40 VSUBS 0.027953f
C1390 VDD1.n41 VSUBS 0.015021f
C1391 VDD1.n42 VSUBS 0.015904f
C1392 VDD1.n43 VSUBS 0.035504f
C1393 VDD1.n44 VSUBS 0.035504f
C1394 VDD1.n45 VSUBS 0.015904f
C1395 VDD1.n46 VSUBS 0.015021f
C1396 VDD1.n47 VSUBS 0.027953f
C1397 VDD1.n48 VSUBS 0.027953f
C1398 VDD1.n49 VSUBS 0.015021f
C1399 VDD1.n50 VSUBS 0.015904f
C1400 VDD1.n51 VSUBS 0.035504f
C1401 VDD1.n52 VSUBS 0.035504f
C1402 VDD1.n53 VSUBS 0.015904f
C1403 VDD1.n54 VSUBS 0.015021f
C1404 VDD1.n55 VSUBS 0.027953f
C1405 VDD1.n56 VSUBS 0.027953f
C1406 VDD1.n57 VSUBS 0.015021f
C1407 VDD1.n58 VSUBS 0.015904f
C1408 VDD1.n59 VSUBS 0.035504f
C1409 VDD1.n60 VSUBS 0.035504f
C1410 VDD1.n61 VSUBS 0.015904f
C1411 VDD1.n62 VSUBS 0.015021f
C1412 VDD1.n63 VSUBS 0.027953f
C1413 VDD1.n64 VSUBS 0.027953f
C1414 VDD1.n65 VSUBS 0.015021f
C1415 VDD1.n66 VSUBS 0.015904f
C1416 VDD1.n67 VSUBS 0.035504f
C1417 VDD1.n68 VSUBS 0.089589f
C1418 VDD1.n69 VSUBS 0.015904f
C1419 VDD1.n70 VSUBS 0.015021f
C1420 VDD1.n71 VSUBS 0.065377f
C1421 VDD1.n72 VSUBS 0.075147f
C1422 VDD1.n73 VSUBS 0.031783f
C1423 VDD1.n74 VSUBS 0.027953f
C1424 VDD1.n75 VSUBS 0.015021f
C1425 VDD1.n76 VSUBS 0.035504f
C1426 VDD1.n77 VSUBS 0.015904f
C1427 VDD1.n78 VSUBS 0.027953f
C1428 VDD1.n79 VSUBS 0.015021f
C1429 VDD1.n80 VSUBS 0.035504f
C1430 VDD1.n81 VSUBS 0.015904f
C1431 VDD1.n82 VSUBS 0.027953f
C1432 VDD1.n83 VSUBS 0.015021f
C1433 VDD1.n84 VSUBS 0.035504f
C1434 VDD1.n85 VSUBS 0.015463f
C1435 VDD1.n86 VSUBS 0.027953f
C1436 VDD1.n87 VSUBS 0.015904f
C1437 VDD1.n88 VSUBS 0.035504f
C1438 VDD1.n89 VSUBS 0.015904f
C1439 VDD1.n90 VSUBS 0.027953f
C1440 VDD1.n91 VSUBS 0.015021f
C1441 VDD1.n92 VSUBS 0.035504f
C1442 VDD1.n93 VSUBS 0.015904f
C1443 VDD1.n94 VSUBS 1.56696f
C1444 VDD1.n95 VSUBS 0.015021f
C1445 VDD1.t1 VSUBS 0.076654f
C1446 VDD1.n96 VSUBS 0.240117f
C1447 VDD1.n97 VSUBS 0.026708f
C1448 VDD1.n98 VSUBS 0.026628f
C1449 VDD1.n99 VSUBS 0.035504f
C1450 VDD1.n100 VSUBS 0.015904f
C1451 VDD1.n101 VSUBS 0.015021f
C1452 VDD1.n102 VSUBS 0.027953f
C1453 VDD1.n103 VSUBS 0.027953f
C1454 VDD1.n104 VSUBS 0.015021f
C1455 VDD1.n105 VSUBS 0.015904f
C1456 VDD1.n106 VSUBS 0.035504f
C1457 VDD1.n107 VSUBS 0.035504f
C1458 VDD1.n108 VSUBS 0.015904f
C1459 VDD1.n109 VSUBS 0.015021f
C1460 VDD1.n110 VSUBS 0.027953f
C1461 VDD1.n111 VSUBS 0.027953f
C1462 VDD1.n112 VSUBS 0.015021f
C1463 VDD1.n113 VSUBS 0.015021f
C1464 VDD1.n114 VSUBS 0.015904f
C1465 VDD1.n115 VSUBS 0.035504f
C1466 VDD1.n116 VSUBS 0.035504f
C1467 VDD1.n117 VSUBS 0.035504f
C1468 VDD1.n118 VSUBS 0.015463f
C1469 VDD1.n119 VSUBS 0.015021f
C1470 VDD1.n120 VSUBS 0.027953f
C1471 VDD1.n121 VSUBS 0.027953f
C1472 VDD1.n122 VSUBS 0.015021f
C1473 VDD1.n123 VSUBS 0.015904f
C1474 VDD1.n124 VSUBS 0.035504f
C1475 VDD1.n125 VSUBS 0.035504f
C1476 VDD1.n126 VSUBS 0.015904f
C1477 VDD1.n127 VSUBS 0.015021f
C1478 VDD1.n128 VSUBS 0.027953f
C1479 VDD1.n129 VSUBS 0.027953f
C1480 VDD1.n130 VSUBS 0.015021f
C1481 VDD1.n131 VSUBS 0.015904f
C1482 VDD1.n132 VSUBS 0.035504f
C1483 VDD1.n133 VSUBS 0.035504f
C1484 VDD1.n134 VSUBS 0.015904f
C1485 VDD1.n135 VSUBS 0.015021f
C1486 VDD1.n136 VSUBS 0.027953f
C1487 VDD1.n137 VSUBS 0.027953f
C1488 VDD1.n138 VSUBS 0.015021f
C1489 VDD1.n139 VSUBS 0.015904f
C1490 VDD1.n140 VSUBS 0.035504f
C1491 VDD1.n141 VSUBS 0.089589f
C1492 VDD1.n142 VSUBS 0.015904f
C1493 VDD1.n143 VSUBS 0.015021f
C1494 VDD1.n144 VSUBS 0.065377f
C1495 VDD1.n145 VSUBS 0.074217f
C1496 VDD1.t2 VSUBS 0.299976f
C1497 VDD1.t3 VSUBS 0.299976f
C1498 VDD1.n146 VSUBS 2.39697f
C1499 VDD1.n147 VSUBS 3.72795f
C1500 VDD1.t4 VSUBS 0.299976f
C1501 VDD1.t0 VSUBS 0.299976f
C1502 VDD1.n148 VSUBS 2.38931f
C1503 VDD1.n149 VSUBS 3.66985f
C1504 VP.n0 VSUBS 0.039683f
C1505 VP.t2 VSUBS 3.29651f
C1506 VP.n1 VSUBS 0.059648f
C1507 VP.n2 VSUBS 0.030101f
C1508 VP.n3 VSUBS 0.042042f
C1509 VP.n4 VSUBS 0.030101f
C1510 VP.n5 VSUBS 0.029299f
C1511 VP.n6 VSUBS 0.030101f
C1512 VP.t1 VSUBS 3.29651f
C1513 VP.n7 VSUBS 1.25421f
C1514 VP.n8 VSUBS 0.039683f
C1515 VP.t3 VSUBS 3.29651f
C1516 VP.n9 VSUBS 0.059648f
C1517 VP.n10 VSUBS 0.030101f
C1518 VP.n11 VSUBS 0.042042f
C1519 VP.t5 VSUBS 3.60482f
C1520 VP.t4 VSUBS 3.29651f
C1521 VP.n12 VSUBS 1.2483f
C1522 VP.n13 VSUBS 1.20609f
C1523 VP.n14 VSUBS 0.320887f
C1524 VP.n15 VSUBS 0.030101f
C1525 VP.n16 VSUBS 0.05582f
C1526 VP.n17 VSUBS 0.054387f
C1527 VP.n18 VSUBS 0.029299f
C1528 VP.n19 VSUBS 0.030101f
C1529 VP.n20 VSUBS 0.030101f
C1530 VP.n21 VSUBS 0.030101f
C1531 VP.n22 VSUBS 0.05582f
C1532 VP.n23 VSUBS 0.029917f
C1533 VP.n24 VSUBS 1.25421f
C1534 VP.n25 VSUBS 1.74495f
C1535 VP.n26 VSUBS 1.76613f
C1536 VP.n27 VSUBS 0.039683f
C1537 VP.n28 VSUBS 0.029917f
C1538 VP.n29 VSUBS 0.05582f
C1539 VP.n30 VSUBS 0.059648f
C1540 VP.n31 VSUBS 0.030101f
C1541 VP.n32 VSUBS 0.030101f
C1542 VP.n33 VSUBS 0.030101f
C1543 VP.n34 VSUBS 0.054387f
C1544 VP.n35 VSUBS 0.05582f
C1545 VP.t0 VSUBS 3.29651f
C1546 VP.n36 VSUBS 1.15404f
C1547 VP.n37 VSUBS 0.042042f
C1548 VP.n38 VSUBS 0.030101f
C1549 VP.n39 VSUBS 0.030101f
C1550 VP.n40 VSUBS 0.030101f
C1551 VP.n41 VSUBS 0.05582f
C1552 VP.n42 VSUBS 0.054387f
C1553 VP.n43 VSUBS 0.029299f
C1554 VP.n44 VSUBS 0.030101f
C1555 VP.n45 VSUBS 0.030101f
C1556 VP.n46 VSUBS 0.030101f
C1557 VP.n47 VSUBS 0.05582f
C1558 VP.n48 VSUBS 0.029917f
C1559 VP.n49 VSUBS 1.25421f
C1560 VP.n50 VSUBS 0.058854f
.ends

