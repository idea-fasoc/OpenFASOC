* NGSPICE file created from diff_pair_sample_1229.ext - technology: sky130A

.subckt diff_pair_sample_1229 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.87265 pd=17.74 as=6.7899 ps=35.6 w=17.41 l=0.55
X1 VDD2.t3 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.87265 pd=17.74 as=6.7899 ps=35.6 w=17.41 l=0.55
X2 VTAIL.t6 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=2.87265 ps=17.74 w=17.41 l=0.55
X3 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=0 ps=0 w=17.41 l=0.55
X4 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.87265 pd=17.74 as=6.7899 ps=35.6 w=17.41 l=0.55
X5 VTAIL.t1 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=2.87265 ps=17.74 w=17.41 l=0.55
X6 VDD1.t1 VP.t2 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.87265 pd=17.74 as=6.7899 ps=35.6 w=17.41 l=0.55
X7 VTAIL.t7 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=2.87265 ps=17.74 w=17.41 l=0.55
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=0 ps=0 w=17.41 l=0.55
X9 VTAIL.t4 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=2.87265 ps=17.74 w=17.41 l=0.55
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=0 ps=0 w=17.41 l=0.55
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.7899 pd=35.6 as=0 ps=0 w=17.41 l=0.55
R0 VP.n0 VP.t3 855.718
R1 VP.n0 VP.t0 855.693
R2 VP.n2 VP.t1 834.736
R3 VP.n3 VP.t2 834.736
R4 VP.n4 VP.n3 161.3
R5 VP.n2 VP.n1 161.3
R6 VP.n1 VP.n0 114.343
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n778 VTAIL.n686 289.615
R11 VTAIL.n92 VTAIL.n0 289.615
R12 VTAIL.n190 VTAIL.n98 289.615
R13 VTAIL.n288 VTAIL.n196 289.615
R14 VTAIL.n680 VTAIL.n588 289.615
R15 VTAIL.n582 VTAIL.n490 289.615
R16 VTAIL.n484 VTAIL.n392 289.615
R17 VTAIL.n386 VTAIL.n294 289.615
R18 VTAIL.n719 VTAIL.n718 185
R19 VTAIL.n721 VTAIL.n720 185
R20 VTAIL.n714 VTAIL.n713 185
R21 VTAIL.n727 VTAIL.n726 185
R22 VTAIL.n729 VTAIL.n728 185
R23 VTAIL.n710 VTAIL.n709 185
R24 VTAIL.n735 VTAIL.n734 185
R25 VTAIL.n737 VTAIL.n736 185
R26 VTAIL.n706 VTAIL.n705 185
R27 VTAIL.n743 VTAIL.n742 185
R28 VTAIL.n745 VTAIL.n744 185
R29 VTAIL.n702 VTAIL.n701 185
R30 VTAIL.n751 VTAIL.n750 185
R31 VTAIL.n753 VTAIL.n752 185
R32 VTAIL.n698 VTAIL.n697 185
R33 VTAIL.n760 VTAIL.n759 185
R34 VTAIL.n761 VTAIL.n696 185
R35 VTAIL.n763 VTAIL.n762 185
R36 VTAIL.n694 VTAIL.n693 185
R37 VTAIL.n769 VTAIL.n768 185
R38 VTAIL.n771 VTAIL.n770 185
R39 VTAIL.n690 VTAIL.n689 185
R40 VTAIL.n777 VTAIL.n776 185
R41 VTAIL.n779 VTAIL.n778 185
R42 VTAIL.n33 VTAIL.n32 185
R43 VTAIL.n35 VTAIL.n34 185
R44 VTAIL.n28 VTAIL.n27 185
R45 VTAIL.n41 VTAIL.n40 185
R46 VTAIL.n43 VTAIL.n42 185
R47 VTAIL.n24 VTAIL.n23 185
R48 VTAIL.n49 VTAIL.n48 185
R49 VTAIL.n51 VTAIL.n50 185
R50 VTAIL.n20 VTAIL.n19 185
R51 VTAIL.n57 VTAIL.n56 185
R52 VTAIL.n59 VTAIL.n58 185
R53 VTAIL.n16 VTAIL.n15 185
R54 VTAIL.n65 VTAIL.n64 185
R55 VTAIL.n67 VTAIL.n66 185
R56 VTAIL.n12 VTAIL.n11 185
R57 VTAIL.n74 VTAIL.n73 185
R58 VTAIL.n75 VTAIL.n10 185
R59 VTAIL.n77 VTAIL.n76 185
R60 VTAIL.n8 VTAIL.n7 185
R61 VTAIL.n83 VTAIL.n82 185
R62 VTAIL.n85 VTAIL.n84 185
R63 VTAIL.n4 VTAIL.n3 185
R64 VTAIL.n91 VTAIL.n90 185
R65 VTAIL.n93 VTAIL.n92 185
R66 VTAIL.n131 VTAIL.n130 185
R67 VTAIL.n133 VTAIL.n132 185
R68 VTAIL.n126 VTAIL.n125 185
R69 VTAIL.n139 VTAIL.n138 185
R70 VTAIL.n141 VTAIL.n140 185
R71 VTAIL.n122 VTAIL.n121 185
R72 VTAIL.n147 VTAIL.n146 185
R73 VTAIL.n149 VTAIL.n148 185
R74 VTAIL.n118 VTAIL.n117 185
R75 VTAIL.n155 VTAIL.n154 185
R76 VTAIL.n157 VTAIL.n156 185
R77 VTAIL.n114 VTAIL.n113 185
R78 VTAIL.n163 VTAIL.n162 185
R79 VTAIL.n165 VTAIL.n164 185
R80 VTAIL.n110 VTAIL.n109 185
R81 VTAIL.n172 VTAIL.n171 185
R82 VTAIL.n173 VTAIL.n108 185
R83 VTAIL.n175 VTAIL.n174 185
R84 VTAIL.n106 VTAIL.n105 185
R85 VTAIL.n181 VTAIL.n180 185
R86 VTAIL.n183 VTAIL.n182 185
R87 VTAIL.n102 VTAIL.n101 185
R88 VTAIL.n189 VTAIL.n188 185
R89 VTAIL.n191 VTAIL.n190 185
R90 VTAIL.n229 VTAIL.n228 185
R91 VTAIL.n231 VTAIL.n230 185
R92 VTAIL.n224 VTAIL.n223 185
R93 VTAIL.n237 VTAIL.n236 185
R94 VTAIL.n239 VTAIL.n238 185
R95 VTAIL.n220 VTAIL.n219 185
R96 VTAIL.n245 VTAIL.n244 185
R97 VTAIL.n247 VTAIL.n246 185
R98 VTAIL.n216 VTAIL.n215 185
R99 VTAIL.n253 VTAIL.n252 185
R100 VTAIL.n255 VTAIL.n254 185
R101 VTAIL.n212 VTAIL.n211 185
R102 VTAIL.n261 VTAIL.n260 185
R103 VTAIL.n263 VTAIL.n262 185
R104 VTAIL.n208 VTAIL.n207 185
R105 VTAIL.n270 VTAIL.n269 185
R106 VTAIL.n271 VTAIL.n206 185
R107 VTAIL.n273 VTAIL.n272 185
R108 VTAIL.n204 VTAIL.n203 185
R109 VTAIL.n279 VTAIL.n278 185
R110 VTAIL.n281 VTAIL.n280 185
R111 VTAIL.n200 VTAIL.n199 185
R112 VTAIL.n287 VTAIL.n286 185
R113 VTAIL.n289 VTAIL.n288 185
R114 VTAIL.n681 VTAIL.n680 185
R115 VTAIL.n679 VTAIL.n678 185
R116 VTAIL.n592 VTAIL.n591 185
R117 VTAIL.n673 VTAIL.n672 185
R118 VTAIL.n671 VTAIL.n670 185
R119 VTAIL.n596 VTAIL.n595 185
R120 VTAIL.n600 VTAIL.n598 185
R121 VTAIL.n665 VTAIL.n664 185
R122 VTAIL.n663 VTAIL.n662 185
R123 VTAIL.n602 VTAIL.n601 185
R124 VTAIL.n657 VTAIL.n656 185
R125 VTAIL.n655 VTAIL.n654 185
R126 VTAIL.n606 VTAIL.n605 185
R127 VTAIL.n649 VTAIL.n648 185
R128 VTAIL.n647 VTAIL.n646 185
R129 VTAIL.n610 VTAIL.n609 185
R130 VTAIL.n641 VTAIL.n640 185
R131 VTAIL.n639 VTAIL.n638 185
R132 VTAIL.n614 VTAIL.n613 185
R133 VTAIL.n633 VTAIL.n632 185
R134 VTAIL.n631 VTAIL.n630 185
R135 VTAIL.n618 VTAIL.n617 185
R136 VTAIL.n625 VTAIL.n624 185
R137 VTAIL.n623 VTAIL.n622 185
R138 VTAIL.n583 VTAIL.n582 185
R139 VTAIL.n581 VTAIL.n580 185
R140 VTAIL.n494 VTAIL.n493 185
R141 VTAIL.n575 VTAIL.n574 185
R142 VTAIL.n573 VTAIL.n572 185
R143 VTAIL.n498 VTAIL.n497 185
R144 VTAIL.n502 VTAIL.n500 185
R145 VTAIL.n567 VTAIL.n566 185
R146 VTAIL.n565 VTAIL.n564 185
R147 VTAIL.n504 VTAIL.n503 185
R148 VTAIL.n559 VTAIL.n558 185
R149 VTAIL.n557 VTAIL.n556 185
R150 VTAIL.n508 VTAIL.n507 185
R151 VTAIL.n551 VTAIL.n550 185
R152 VTAIL.n549 VTAIL.n548 185
R153 VTAIL.n512 VTAIL.n511 185
R154 VTAIL.n543 VTAIL.n542 185
R155 VTAIL.n541 VTAIL.n540 185
R156 VTAIL.n516 VTAIL.n515 185
R157 VTAIL.n535 VTAIL.n534 185
R158 VTAIL.n533 VTAIL.n532 185
R159 VTAIL.n520 VTAIL.n519 185
R160 VTAIL.n527 VTAIL.n526 185
R161 VTAIL.n525 VTAIL.n524 185
R162 VTAIL.n485 VTAIL.n484 185
R163 VTAIL.n483 VTAIL.n482 185
R164 VTAIL.n396 VTAIL.n395 185
R165 VTAIL.n477 VTAIL.n476 185
R166 VTAIL.n475 VTAIL.n474 185
R167 VTAIL.n400 VTAIL.n399 185
R168 VTAIL.n404 VTAIL.n402 185
R169 VTAIL.n469 VTAIL.n468 185
R170 VTAIL.n467 VTAIL.n466 185
R171 VTAIL.n406 VTAIL.n405 185
R172 VTAIL.n461 VTAIL.n460 185
R173 VTAIL.n459 VTAIL.n458 185
R174 VTAIL.n410 VTAIL.n409 185
R175 VTAIL.n453 VTAIL.n452 185
R176 VTAIL.n451 VTAIL.n450 185
R177 VTAIL.n414 VTAIL.n413 185
R178 VTAIL.n445 VTAIL.n444 185
R179 VTAIL.n443 VTAIL.n442 185
R180 VTAIL.n418 VTAIL.n417 185
R181 VTAIL.n437 VTAIL.n436 185
R182 VTAIL.n435 VTAIL.n434 185
R183 VTAIL.n422 VTAIL.n421 185
R184 VTAIL.n429 VTAIL.n428 185
R185 VTAIL.n427 VTAIL.n426 185
R186 VTAIL.n387 VTAIL.n386 185
R187 VTAIL.n385 VTAIL.n384 185
R188 VTAIL.n298 VTAIL.n297 185
R189 VTAIL.n379 VTAIL.n378 185
R190 VTAIL.n377 VTAIL.n376 185
R191 VTAIL.n302 VTAIL.n301 185
R192 VTAIL.n306 VTAIL.n304 185
R193 VTAIL.n371 VTAIL.n370 185
R194 VTAIL.n369 VTAIL.n368 185
R195 VTAIL.n308 VTAIL.n307 185
R196 VTAIL.n363 VTAIL.n362 185
R197 VTAIL.n361 VTAIL.n360 185
R198 VTAIL.n312 VTAIL.n311 185
R199 VTAIL.n355 VTAIL.n354 185
R200 VTAIL.n353 VTAIL.n352 185
R201 VTAIL.n316 VTAIL.n315 185
R202 VTAIL.n347 VTAIL.n346 185
R203 VTAIL.n345 VTAIL.n344 185
R204 VTAIL.n320 VTAIL.n319 185
R205 VTAIL.n339 VTAIL.n338 185
R206 VTAIL.n337 VTAIL.n336 185
R207 VTAIL.n324 VTAIL.n323 185
R208 VTAIL.n331 VTAIL.n330 185
R209 VTAIL.n329 VTAIL.n328 185
R210 VTAIL.n717 VTAIL.t2 147.659
R211 VTAIL.n31 VTAIL.t1 147.659
R212 VTAIL.n129 VTAIL.t3 147.659
R213 VTAIL.n227 VTAIL.t6 147.659
R214 VTAIL.n621 VTAIL.t5 147.659
R215 VTAIL.n523 VTAIL.t4 147.659
R216 VTAIL.n425 VTAIL.t0 147.659
R217 VTAIL.n327 VTAIL.t7 147.659
R218 VTAIL.n720 VTAIL.n719 104.615
R219 VTAIL.n720 VTAIL.n713 104.615
R220 VTAIL.n727 VTAIL.n713 104.615
R221 VTAIL.n728 VTAIL.n727 104.615
R222 VTAIL.n728 VTAIL.n709 104.615
R223 VTAIL.n735 VTAIL.n709 104.615
R224 VTAIL.n736 VTAIL.n735 104.615
R225 VTAIL.n736 VTAIL.n705 104.615
R226 VTAIL.n743 VTAIL.n705 104.615
R227 VTAIL.n744 VTAIL.n743 104.615
R228 VTAIL.n744 VTAIL.n701 104.615
R229 VTAIL.n751 VTAIL.n701 104.615
R230 VTAIL.n752 VTAIL.n751 104.615
R231 VTAIL.n752 VTAIL.n697 104.615
R232 VTAIL.n760 VTAIL.n697 104.615
R233 VTAIL.n761 VTAIL.n760 104.615
R234 VTAIL.n762 VTAIL.n761 104.615
R235 VTAIL.n762 VTAIL.n693 104.615
R236 VTAIL.n769 VTAIL.n693 104.615
R237 VTAIL.n770 VTAIL.n769 104.615
R238 VTAIL.n770 VTAIL.n689 104.615
R239 VTAIL.n777 VTAIL.n689 104.615
R240 VTAIL.n778 VTAIL.n777 104.615
R241 VTAIL.n34 VTAIL.n33 104.615
R242 VTAIL.n34 VTAIL.n27 104.615
R243 VTAIL.n41 VTAIL.n27 104.615
R244 VTAIL.n42 VTAIL.n41 104.615
R245 VTAIL.n42 VTAIL.n23 104.615
R246 VTAIL.n49 VTAIL.n23 104.615
R247 VTAIL.n50 VTAIL.n49 104.615
R248 VTAIL.n50 VTAIL.n19 104.615
R249 VTAIL.n57 VTAIL.n19 104.615
R250 VTAIL.n58 VTAIL.n57 104.615
R251 VTAIL.n58 VTAIL.n15 104.615
R252 VTAIL.n65 VTAIL.n15 104.615
R253 VTAIL.n66 VTAIL.n65 104.615
R254 VTAIL.n66 VTAIL.n11 104.615
R255 VTAIL.n74 VTAIL.n11 104.615
R256 VTAIL.n75 VTAIL.n74 104.615
R257 VTAIL.n76 VTAIL.n75 104.615
R258 VTAIL.n76 VTAIL.n7 104.615
R259 VTAIL.n83 VTAIL.n7 104.615
R260 VTAIL.n84 VTAIL.n83 104.615
R261 VTAIL.n84 VTAIL.n3 104.615
R262 VTAIL.n91 VTAIL.n3 104.615
R263 VTAIL.n92 VTAIL.n91 104.615
R264 VTAIL.n132 VTAIL.n131 104.615
R265 VTAIL.n132 VTAIL.n125 104.615
R266 VTAIL.n139 VTAIL.n125 104.615
R267 VTAIL.n140 VTAIL.n139 104.615
R268 VTAIL.n140 VTAIL.n121 104.615
R269 VTAIL.n147 VTAIL.n121 104.615
R270 VTAIL.n148 VTAIL.n147 104.615
R271 VTAIL.n148 VTAIL.n117 104.615
R272 VTAIL.n155 VTAIL.n117 104.615
R273 VTAIL.n156 VTAIL.n155 104.615
R274 VTAIL.n156 VTAIL.n113 104.615
R275 VTAIL.n163 VTAIL.n113 104.615
R276 VTAIL.n164 VTAIL.n163 104.615
R277 VTAIL.n164 VTAIL.n109 104.615
R278 VTAIL.n172 VTAIL.n109 104.615
R279 VTAIL.n173 VTAIL.n172 104.615
R280 VTAIL.n174 VTAIL.n173 104.615
R281 VTAIL.n174 VTAIL.n105 104.615
R282 VTAIL.n181 VTAIL.n105 104.615
R283 VTAIL.n182 VTAIL.n181 104.615
R284 VTAIL.n182 VTAIL.n101 104.615
R285 VTAIL.n189 VTAIL.n101 104.615
R286 VTAIL.n190 VTAIL.n189 104.615
R287 VTAIL.n230 VTAIL.n229 104.615
R288 VTAIL.n230 VTAIL.n223 104.615
R289 VTAIL.n237 VTAIL.n223 104.615
R290 VTAIL.n238 VTAIL.n237 104.615
R291 VTAIL.n238 VTAIL.n219 104.615
R292 VTAIL.n245 VTAIL.n219 104.615
R293 VTAIL.n246 VTAIL.n245 104.615
R294 VTAIL.n246 VTAIL.n215 104.615
R295 VTAIL.n253 VTAIL.n215 104.615
R296 VTAIL.n254 VTAIL.n253 104.615
R297 VTAIL.n254 VTAIL.n211 104.615
R298 VTAIL.n261 VTAIL.n211 104.615
R299 VTAIL.n262 VTAIL.n261 104.615
R300 VTAIL.n262 VTAIL.n207 104.615
R301 VTAIL.n270 VTAIL.n207 104.615
R302 VTAIL.n271 VTAIL.n270 104.615
R303 VTAIL.n272 VTAIL.n271 104.615
R304 VTAIL.n272 VTAIL.n203 104.615
R305 VTAIL.n279 VTAIL.n203 104.615
R306 VTAIL.n280 VTAIL.n279 104.615
R307 VTAIL.n280 VTAIL.n199 104.615
R308 VTAIL.n287 VTAIL.n199 104.615
R309 VTAIL.n288 VTAIL.n287 104.615
R310 VTAIL.n680 VTAIL.n679 104.615
R311 VTAIL.n679 VTAIL.n591 104.615
R312 VTAIL.n672 VTAIL.n591 104.615
R313 VTAIL.n672 VTAIL.n671 104.615
R314 VTAIL.n671 VTAIL.n595 104.615
R315 VTAIL.n600 VTAIL.n595 104.615
R316 VTAIL.n664 VTAIL.n600 104.615
R317 VTAIL.n664 VTAIL.n663 104.615
R318 VTAIL.n663 VTAIL.n601 104.615
R319 VTAIL.n656 VTAIL.n601 104.615
R320 VTAIL.n656 VTAIL.n655 104.615
R321 VTAIL.n655 VTAIL.n605 104.615
R322 VTAIL.n648 VTAIL.n605 104.615
R323 VTAIL.n648 VTAIL.n647 104.615
R324 VTAIL.n647 VTAIL.n609 104.615
R325 VTAIL.n640 VTAIL.n609 104.615
R326 VTAIL.n640 VTAIL.n639 104.615
R327 VTAIL.n639 VTAIL.n613 104.615
R328 VTAIL.n632 VTAIL.n613 104.615
R329 VTAIL.n632 VTAIL.n631 104.615
R330 VTAIL.n631 VTAIL.n617 104.615
R331 VTAIL.n624 VTAIL.n617 104.615
R332 VTAIL.n624 VTAIL.n623 104.615
R333 VTAIL.n582 VTAIL.n581 104.615
R334 VTAIL.n581 VTAIL.n493 104.615
R335 VTAIL.n574 VTAIL.n493 104.615
R336 VTAIL.n574 VTAIL.n573 104.615
R337 VTAIL.n573 VTAIL.n497 104.615
R338 VTAIL.n502 VTAIL.n497 104.615
R339 VTAIL.n566 VTAIL.n502 104.615
R340 VTAIL.n566 VTAIL.n565 104.615
R341 VTAIL.n565 VTAIL.n503 104.615
R342 VTAIL.n558 VTAIL.n503 104.615
R343 VTAIL.n558 VTAIL.n557 104.615
R344 VTAIL.n557 VTAIL.n507 104.615
R345 VTAIL.n550 VTAIL.n507 104.615
R346 VTAIL.n550 VTAIL.n549 104.615
R347 VTAIL.n549 VTAIL.n511 104.615
R348 VTAIL.n542 VTAIL.n511 104.615
R349 VTAIL.n542 VTAIL.n541 104.615
R350 VTAIL.n541 VTAIL.n515 104.615
R351 VTAIL.n534 VTAIL.n515 104.615
R352 VTAIL.n534 VTAIL.n533 104.615
R353 VTAIL.n533 VTAIL.n519 104.615
R354 VTAIL.n526 VTAIL.n519 104.615
R355 VTAIL.n526 VTAIL.n525 104.615
R356 VTAIL.n484 VTAIL.n483 104.615
R357 VTAIL.n483 VTAIL.n395 104.615
R358 VTAIL.n476 VTAIL.n395 104.615
R359 VTAIL.n476 VTAIL.n475 104.615
R360 VTAIL.n475 VTAIL.n399 104.615
R361 VTAIL.n404 VTAIL.n399 104.615
R362 VTAIL.n468 VTAIL.n404 104.615
R363 VTAIL.n468 VTAIL.n467 104.615
R364 VTAIL.n467 VTAIL.n405 104.615
R365 VTAIL.n460 VTAIL.n405 104.615
R366 VTAIL.n460 VTAIL.n459 104.615
R367 VTAIL.n459 VTAIL.n409 104.615
R368 VTAIL.n452 VTAIL.n409 104.615
R369 VTAIL.n452 VTAIL.n451 104.615
R370 VTAIL.n451 VTAIL.n413 104.615
R371 VTAIL.n444 VTAIL.n413 104.615
R372 VTAIL.n444 VTAIL.n443 104.615
R373 VTAIL.n443 VTAIL.n417 104.615
R374 VTAIL.n436 VTAIL.n417 104.615
R375 VTAIL.n436 VTAIL.n435 104.615
R376 VTAIL.n435 VTAIL.n421 104.615
R377 VTAIL.n428 VTAIL.n421 104.615
R378 VTAIL.n428 VTAIL.n427 104.615
R379 VTAIL.n386 VTAIL.n385 104.615
R380 VTAIL.n385 VTAIL.n297 104.615
R381 VTAIL.n378 VTAIL.n297 104.615
R382 VTAIL.n378 VTAIL.n377 104.615
R383 VTAIL.n377 VTAIL.n301 104.615
R384 VTAIL.n306 VTAIL.n301 104.615
R385 VTAIL.n370 VTAIL.n306 104.615
R386 VTAIL.n370 VTAIL.n369 104.615
R387 VTAIL.n369 VTAIL.n307 104.615
R388 VTAIL.n362 VTAIL.n307 104.615
R389 VTAIL.n362 VTAIL.n361 104.615
R390 VTAIL.n361 VTAIL.n311 104.615
R391 VTAIL.n354 VTAIL.n311 104.615
R392 VTAIL.n354 VTAIL.n353 104.615
R393 VTAIL.n353 VTAIL.n315 104.615
R394 VTAIL.n346 VTAIL.n315 104.615
R395 VTAIL.n346 VTAIL.n345 104.615
R396 VTAIL.n345 VTAIL.n319 104.615
R397 VTAIL.n338 VTAIL.n319 104.615
R398 VTAIL.n338 VTAIL.n337 104.615
R399 VTAIL.n337 VTAIL.n323 104.615
R400 VTAIL.n330 VTAIL.n323 104.615
R401 VTAIL.n330 VTAIL.n329 104.615
R402 VTAIL.n719 VTAIL.t2 52.3082
R403 VTAIL.n33 VTAIL.t1 52.3082
R404 VTAIL.n131 VTAIL.t3 52.3082
R405 VTAIL.n229 VTAIL.t6 52.3082
R406 VTAIL.n623 VTAIL.t5 52.3082
R407 VTAIL.n525 VTAIL.t4 52.3082
R408 VTAIL.n427 VTAIL.t0 52.3082
R409 VTAIL.n329 VTAIL.t7 52.3082
R410 VTAIL.n783 VTAIL.n782 30.052
R411 VTAIL.n97 VTAIL.n96 30.052
R412 VTAIL.n195 VTAIL.n194 30.052
R413 VTAIL.n293 VTAIL.n292 30.052
R414 VTAIL.n685 VTAIL.n684 30.052
R415 VTAIL.n587 VTAIL.n586 30.052
R416 VTAIL.n489 VTAIL.n488 30.052
R417 VTAIL.n391 VTAIL.n390 30.052
R418 VTAIL.n783 VTAIL.n685 28.1341
R419 VTAIL.n391 VTAIL.n293 28.1341
R420 VTAIL.n718 VTAIL.n717 15.6677
R421 VTAIL.n32 VTAIL.n31 15.6677
R422 VTAIL.n130 VTAIL.n129 15.6677
R423 VTAIL.n228 VTAIL.n227 15.6677
R424 VTAIL.n622 VTAIL.n621 15.6677
R425 VTAIL.n524 VTAIL.n523 15.6677
R426 VTAIL.n426 VTAIL.n425 15.6677
R427 VTAIL.n328 VTAIL.n327 15.6677
R428 VTAIL.n763 VTAIL.n694 13.1884
R429 VTAIL.n77 VTAIL.n8 13.1884
R430 VTAIL.n175 VTAIL.n106 13.1884
R431 VTAIL.n273 VTAIL.n204 13.1884
R432 VTAIL.n598 VTAIL.n596 13.1884
R433 VTAIL.n500 VTAIL.n498 13.1884
R434 VTAIL.n402 VTAIL.n400 13.1884
R435 VTAIL.n304 VTAIL.n302 13.1884
R436 VTAIL.n721 VTAIL.n716 12.8005
R437 VTAIL.n764 VTAIL.n696 12.8005
R438 VTAIL.n768 VTAIL.n767 12.8005
R439 VTAIL.n35 VTAIL.n30 12.8005
R440 VTAIL.n78 VTAIL.n10 12.8005
R441 VTAIL.n82 VTAIL.n81 12.8005
R442 VTAIL.n133 VTAIL.n128 12.8005
R443 VTAIL.n176 VTAIL.n108 12.8005
R444 VTAIL.n180 VTAIL.n179 12.8005
R445 VTAIL.n231 VTAIL.n226 12.8005
R446 VTAIL.n274 VTAIL.n206 12.8005
R447 VTAIL.n278 VTAIL.n277 12.8005
R448 VTAIL.n670 VTAIL.n669 12.8005
R449 VTAIL.n666 VTAIL.n665 12.8005
R450 VTAIL.n625 VTAIL.n620 12.8005
R451 VTAIL.n572 VTAIL.n571 12.8005
R452 VTAIL.n568 VTAIL.n567 12.8005
R453 VTAIL.n527 VTAIL.n522 12.8005
R454 VTAIL.n474 VTAIL.n473 12.8005
R455 VTAIL.n470 VTAIL.n469 12.8005
R456 VTAIL.n429 VTAIL.n424 12.8005
R457 VTAIL.n376 VTAIL.n375 12.8005
R458 VTAIL.n372 VTAIL.n371 12.8005
R459 VTAIL.n331 VTAIL.n326 12.8005
R460 VTAIL.n722 VTAIL.n714 12.0247
R461 VTAIL.n759 VTAIL.n758 12.0247
R462 VTAIL.n771 VTAIL.n692 12.0247
R463 VTAIL.n36 VTAIL.n28 12.0247
R464 VTAIL.n73 VTAIL.n72 12.0247
R465 VTAIL.n85 VTAIL.n6 12.0247
R466 VTAIL.n134 VTAIL.n126 12.0247
R467 VTAIL.n171 VTAIL.n170 12.0247
R468 VTAIL.n183 VTAIL.n104 12.0247
R469 VTAIL.n232 VTAIL.n224 12.0247
R470 VTAIL.n269 VTAIL.n268 12.0247
R471 VTAIL.n281 VTAIL.n202 12.0247
R472 VTAIL.n673 VTAIL.n594 12.0247
R473 VTAIL.n662 VTAIL.n599 12.0247
R474 VTAIL.n626 VTAIL.n618 12.0247
R475 VTAIL.n575 VTAIL.n496 12.0247
R476 VTAIL.n564 VTAIL.n501 12.0247
R477 VTAIL.n528 VTAIL.n520 12.0247
R478 VTAIL.n477 VTAIL.n398 12.0247
R479 VTAIL.n466 VTAIL.n403 12.0247
R480 VTAIL.n430 VTAIL.n422 12.0247
R481 VTAIL.n379 VTAIL.n300 12.0247
R482 VTAIL.n368 VTAIL.n305 12.0247
R483 VTAIL.n332 VTAIL.n324 12.0247
R484 VTAIL.n726 VTAIL.n725 11.249
R485 VTAIL.n757 VTAIL.n698 11.249
R486 VTAIL.n772 VTAIL.n690 11.249
R487 VTAIL.n40 VTAIL.n39 11.249
R488 VTAIL.n71 VTAIL.n12 11.249
R489 VTAIL.n86 VTAIL.n4 11.249
R490 VTAIL.n138 VTAIL.n137 11.249
R491 VTAIL.n169 VTAIL.n110 11.249
R492 VTAIL.n184 VTAIL.n102 11.249
R493 VTAIL.n236 VTAIL.n235 11.249
R494 VTAIL.n267 VTAIL.n208 11.249
R495 VTAIL.n282 VTAIL.n200 11.249
R496 VTAIL.n674 VTAIL.n592 11.249
R497 VTAIL.n661 VTAIL.n602 11.249
R498 VTAIL.n630 VTAIL.n629 11.249
R499 VTAIL.n576 VTAIL.n494 11.249
R500 VTAIL.n563 VTAIL.n504 11.249
R501 VTAIL.n532 VTAIL.n531 11.249
R502 VTAIL.n478 VTAIL.n396 11.249
R503 VTAIL.n465 VTAIL.n406 11.249
R504 VTAIL.n434 VTAIL.n433 11.249
R505 VTAIL.n380 VTAIL.n298 11.249
R506 VTAIL.n367 VTAIL.n308 11.249
R507 VTAIL.n336 VTAIL.n335 11.249
R508 VTAIL.n729 VTAIL.n712 10.4732
R509 VTAIL.n754 VTAIL.n753 10.4732
R510 VTAIL.n776 VTAIL.n775 10.4732
R511 VTAIL.n43 VTAIL.n26 10.4732
R512 VTAIL.n68 VTAIL.n67 10.4732
R513 VTAIL.n90 VTAIL.n89 10.4732
R514 VTAIL.n141 VTAIL.n124 10.4732
R515 VTAIL.n166 VTAIL.n165 10.4732
R516 VTAIL.n188 VTAIL.n187 10.4732
R517 VTAIL.n239 VTAIL.n222 10.4732
R518 VTAIL.n264 VTAIL.n263 10.4732
R519 VTAIL.n286 VTAIL.n285 10.4732
R520 VTAIL.n678 VTAIL.n677 10.4732
R521 VTAIL.n658 VTAIL.n657 10.4732
R522 VTAIL.n633 VTAIL.n616 10.4732
R523 VTAIL.n580 VTAIL.n579 10.4732
R524 VTAIL.n560 VTAIL.n559 10.4732
R525 VTAIL.n535 VTAIL.n518 10.4732
R526 VTAIL.n482 VTAIL.n481 10.4732
R527 VTAIL.n462 VTAIL.n461 10.4732
R528 VTAIL.n437 VTAIL.n420 10.4732
R529 VTAIL.n384 VTAIL.n383 10.4732
R530 VTAIL.n364 VTAIL.n363 10.4732
R531 VTAIL.n339 VTAIL.n322 10.4732
R532 VTAIL.n730 VTAIL.n710 9.69747
R533 VTAIL.n750 VTAIL.n700 9.69747
R534 VTAIL.n779 VTAIL.n688 9.69747
R535 VTAIL.n44 VTAIL.n24 9.69747
R536 VTAIL.n64 VTAIL.n14 9.69747
R537 VTAIL.n93 VTAIL.n2 9.69747
R538 VTAIL.n142 VTAIL.n122 9.69747
R539 VTAIL.n162 VTAIL.n112 9.69747
R540 VTAIL.n191 VTAIL.n100 9.69747
R541 VTAIL.n240 VTAIL.n220 9.69747
R542 VTAIL.n260 VTAIL.n210 9.69747
R543 VTAIL.n289 VTAIL.n198 9.69747
R544 VTAIL.n681 VTAIL.n590 9.69747
R545 VTAIL.n654 VTAIL.n604 9.69747
R546 VTAIL.n634 VTAIL.n614 9.69747
R547 VTAIL.n583 VTAIL.n492 9.69747
R548 VTAIL.n556 VTAIL.n506 9.69747
R549 VTAIL.n536 VTAIL.n516 9.69747
R550 VTAIL.n485 VTAIL.n394 9.69747
R551 VTAIL.n458 VTAIL.n408 9.69747
R552 VTAIL.n438 VTAIL.n418 9.69747
R553 VTAIL.n387 VTAIL.n296 9.69747
R554 VTAIL.n360 VTAIL.n310 9.69747
R555 VTAIL.n340 VTAIL.n320 9.69747
R556 VTAIL.n782 VTAIL.n781 9.45567
R557 VTAIL.n96 VTAIL.n95 9.45567
R558 VTAIL.n194 VTAIL.n193 9.45567
R559 VTAIL.n292 VTAIL.n291 9.45567
R560 VTAIL.n684 VTAIL.n683 9.45567
R561 VTAIL.n586 VTAIL.n585 9.45567
R562 VTAIL.n488 VTAIL.n487 9.45567
R563 VTAIL.n390 VTAIL.n389 9.45567
R564 VTAIL.n781 VTAIL.n780 9.3005
R565 VTAIL.n688 VTAIL.n687 9.3005
R566 VTAIL.n775 VTAIL.n774 9.3005
R567 VTAIL.n773 VTAIL.n772 9.3005
R568 VTAIL.n692 VTAIL.n691 9.3005
R569 VTAIL.n767 VTAIL.n766 9.3005
R570 VTAIL.n739 VTAIL.n738 9.3005
R571 VTAIL.n708 VTAIL.n707 9.3005
R572 VTAIL.n733 VTAIL.n732 9.3005
R573 VTAIL.n731 VTAIL.n730 9.3005
R574 VTAIL.n712 VTAIL.n711 9.3005
R575 VTAIL.n725 VTAIL.n724 9.3005
R576 VTAIL.n723 VTAIL.n722 9.3005
R577 VTAIL.n716 VTAIL.n715 9.3005
R578 VTAIL.n741 VTAIL.n740 9.3005
R579 VTAIL.n704 VTAIL.n703 9.3005
R580 VTAIL.n747 VTAIL.n746 9.3005
R581 VTAIL.n749 VTAIL.n748 9.3005
R582 VTAIL.n700 VTAIL.n699 9.3005
R583 VTAIL.n755 VTAIL.n754 9.3005
R584 VTAIL.n757 VTAIL.n756 9.3005
R585 VTAIL.n758 VTAIL.n695 9.3005
R586 VTAIL.n765 VTAIL.n764 9.3005
R587 VTAIL.n95 VTAIL.n94 9.3005
R588 VTAIL.n2 VTAIL.n1 9.3005
R589 VTAIL.n89 VTAIL.n88 9.3005
R590 VTAIL.n87 VTAIL.n86 9.3005
R591 VTAIL.n6 VTAIL.n5 9.3005
R592 VTAIL.n81 VTAIL.n80 9.3005
R593 VTAIL.n53 VTAIL.n52 9.3005
R594 VTAIL.n22 VTAIL.n21 9.3005
R595 VTAIL.n47 VTAIL.n46 9.3005
R596 VTAIL.n45 VTAIL.n44 9.3005
R597 VTAIL.n26 VTAIL.n25 9.3005
R598 VTAIL.n39 VTAIL.n38 9.3005
R599 VTAIL.n37 VTAIL.n36 9.3005
R600 VTAIL.n30 VTAIL.n29 9.3005
R601 VTAIL.n55 VTAIL.n54 9.3005
R602 VTAIL.n18 VTAIL.n17 9.3005
R603 VTAIL.n61 VTAIL.n60 9.3005
R604 VTAIL.n63 VTAIL.n62 9.3005
R605 VTAIL.n14 VTAIL.n13 9.3005
R606 VTAIL.n69 VTAIL.n68 9.3005
R607 VTAIL.n71 VTAIL.n70 9.3005
R608 VTAIL.n72 VTAIL.n9 9.3005
R609 VTAIL.n79 VTAIL.n78 9.3005
R610 VTAIL.n193 VTAIL.n192 9.3005
R611 VTAIL.n100 VTAIL.n99 9.3005
R612 VTAIL.n187 VTAIL.n186 9.3005
R613 VTAIL.n185 VTAIL.n184 9.3005
R614 VTAIL.n104 VTAIL.n103 9.3005
R615 VTAIL.n179 VTAIL.n178 9.3005
R616 VTAIL.n151 VTAIL.n150 9.3005
R617 VTAIL.n120 VTAIL.n119 9.3005
R618 VTAIL.n145 VTAIL.n144 9.3005
R619 VTAIL.n143 VTAIL.n142 9.3005
R620 VTAIL.n124 VTAIL.n123 9.3005
R621 VTAIL.n137 VTAIL.n136 9.3005
R622 VTAIL.n135 VTAIL.n134 9.3005
R623 VTAIL.n128 VTAIL.n127 9.3005
R624 VTAIL.n153 VTAIL.n152 9.3005
R625 VTAIL.n116 VTAIL.n115 9.3005
R626 VTAIL.n159 VTAIL.n158 9.3005
R627 VTAIL.n161 VTAIL.n160 9.3005
R628 VTAIL.n112 VTAIL.n111 9.3005
R629 VTAIL.n167 VTAIL.n166 9.3005
R630 VTAIL.n169 VTAIL.n168 9.3005
R631 VTAIL.n170 VTAIL.n107 9.3005
R632 VTAIL.n177 VTAIL.n176 9.3005
R633 VTAIL.n291 VTAIL.n290 9.3005
R634 VTAIL.n198 VTAIL.n197 9.3005
R635 VTAIL.n285 VTAIL.n284 9.3005
R636 VTAIL.n283 VTAIL.n282 9.3005
R637 VTAIL.n202 VTAIL.n201 9.3005
R638 VTAIL.n277 VTAIL.n276 9.3005
R639 VTAIL.n249 VTAIL.n248 9.3005
R640 VTAIL.n218 VTAIL.n217 9.3005
R641 VTAIL.n243 VTAIL.n242 9.3005
R642 VTAIL.n241 VTAIL.n240 9.3005
R643 VTAIL.n222 VTAIL.n221 9.3005
R644 VTAIL.n235 VTAIL.n234 9.3005
R645 VTAIL.n233 VTAIL.n232 9.3005
R646 VTAIL.n226 VTAIL.n225 9.3005
R647 VTAIL.n251 VTAIL.n250 9.3005
R648 VTAIL.n214 VTAIL.n213 9.3005
R649 VTAIL.n257 VTAIL.n256 9.3005
R650 VTAIL.n259 VTAIL.n258 9.3005
R651 VTAIL.n210 VTAIL.n209 9.3005
R652 VTAIL.n265 VTAIL.n264 9.3005
R653 VTAIL.n267 VTAIL.n266 9.3005
R654 VTAIL.n268 VTAIL.n205 9.3005
R655 VTAIL.n275 VTAIL.n274 9.3005
R656 VTAIL.n608 VTAIL.n607 9.3005
R657 VTAIL.n651 VTAIL.n650 9.3005
R658 VTAIL.n653 VTAIL.n652 9.3005
R659 VTAIL.n604 VTAIL.n603 9.3005
R660 VTAIL.n659 VTAIL.n658 9.3005
R661 VTAIL.n661 VTAIL.n660 9.3005
R662 VTAIL.n599 VTAIL.n597 9.3005
R663 VTAIL.n667 VTAIL.n666 9.3005
R664 VTAIL.n683 VTAIL.n682 9.3005
R665 VTAIL.n590 VTAIL.n589 9.3005
R666 VTAIL.n677 VTAIL.n676 9.3005
R667 VTAIL.n675 VTAIL.n674 9.3005
R668 VTAIL.n594 VTAIL.n593 9.3005
R669 VTAIL.n669 VTAIL.n668 9.3005
R670 VTAIL.n645 VTAIL.n644 9.3005
R671 VTAIL.n643 VTAIL.n642 9.3005
R672 VTAIL.n612 VTAIL.n611 9.3005
R673 VTAIL.n637 VTAIL.n636 9.3005
R674 VTAIL.n635 VTAIL.n634 9.3005
R675 VTAIL.n616 VTAIL.n615 9.3005
R676 VTAIL.n629 VTAIL.n628 9.3005
R677 VTAIL.n627 VTAIL.n626 9.3005
R678 VTAIL.n620 VTAIL.n619 9.3005
R679 VTAIL.n510 VTAIL.n509 9.3005
R680 VTAIL.n553 VTAIL.n552 9.3005
R681 VTAIL.n555 VTAIL.n554 9.3005
R682 VTAIL.n506 VTAIL.n505 9.3005
R683 VTAIL.n561 VTAIL.n560 9.3005
R684 VTAIL.n563 VTAIL.n562 9.3005
R685 VTAIL.n501 VTAIL.n499 9.3005
R686 VTAIL.n569 VTAIL.n568 9.3005
R687 VTAIL.n585 VTAIL.n584 9.3005
R688 VTAIL.n492 VTAIL.n491 9.3005
R689 VTAIL.n579 VTAIL.n578 9.3005
R690 VTAIL.n577 VTAIL.n576 9.3005
R691 VTAIL.n496 VTAIL.n495 9.3005
R692 VTAIL.n571 VTAIL.n570 9.3005
R693 VTAIL.n547 VTAIL.n546 9.3005
R694 VTAIL.n545 VTAIL.n544 9.3005
R695 VTAIL.n514 VTAIL.n513 9.3005
R696 VTAIL.n539 VTAIL.n538 9.3005
R697 VTAIL.n537 VTAIL.n536 9.3005
R698 VTAIL.n518 VTAIL.n517 9.3005
R699 VTAIL.n531 VTAIL.n530 9.3005
R700 VTAIL.n529 VTAIL.n528 9.3005
R701 VTAIL.n522 VTAIL.n521 9.3005
R702 VTAIL.n412 VTAIL.n411 9.3005
R703 VTAIL.n455 VTAIL.n454 9.3005
R704 VTAIL.n457 VTAIL.n456 9.3005
R705 VTAIL.n408 VTAIL.n407 9.3005
R706 VTAIL.n463 VTAIL.n462 9.3005
R707 VTAIL.n465 VTAIL.n464 9.3005
R708 VTAIL.n403 VTAIL.n401 9.3005
R709 VTAIL.n471 VTAIL.n470 9.3005
R710 VTAIL.n487 VTAIL.n486 9.3005
R711 VTAIL.n394 VTAIL.n393 9.3005
R712 VTAIL.n481 VTAIL.n480 9.3005
R713 VTAIL.n479 VTAIL.n478 9.3005
R714 VTAIL.n398 VTAIL.n397 9.3005
R715 VTAIL.n473 VTAIL.n472 9.3005
R716 VTAIL.n449 VTAIL.n448 9.3005
R717 VTAIL.n447 VTAIL.n446 9.3005
R718 VTAIL.n416 VTAIL.n415 9.3005
R719 VTAIL.n441 VTAIL.n440 9.3005
R720 VTAIL.n439 VTAIL.n438 9.3005
R721 VTAIL.n420 VTAIL.n419 9.3005
R722 VTAIL.n433 VTAIL.n432 9.3005
R723 VTAIL.n431 VTAIL.n430 9.3005
R724 VTAIL.n424 VTAIL.n423 9.3005
R725 VTAIL.n314 VTAIL.n313 9.3005
R726 VTAIL.n357 VTAIL.n356 9.3005
R727 VTAIL.n359 VTAIL.n358 9.3005
R728 VTAIL.n310 VTAIL.n309 9.3005
R729 VTAIL.n365 VTAIL.n364 9.3005
R730 VTAIL.n367 VTAIL.n366 9.3005
R731 VTAIL.n305 VTAIL.n303 9.3005
R732 VTAIL.n373 VTAIL.n372 9.3005
R733 VTAIL.n389 VTAIL.n388 9.3005
R734 VTAIL.n296 VTAIL.n295 9.3005
R735 VTAIL.n383 VTAIL.n382 9.3005
R736 VTAIL.n381 VTAIL.n380 9.3005
R737 VTAIL.n300 VTAIL.n299 9.3005
R738 VTAIL.n375 VTAIL.n374 9.3005
R739 VTAIL.n351 VTAIL.n350 9.3005
R740 VTAIL.n349 VTAIL.n348 9.3005
R741 VTAIL.n318 VTAIL.n317 9.3005
R742 VTAIL.n343 VTAIL.n342 9.3005
R743 VTAIL.n341 VTAIL.n340 9.3005
R744 VTAIL.n322 VTAIL.n321 9.3005
R745 VTAIL.n335 VTAIL.n334 9.3005
R746 VTAIL.n333 VTAIL.n332 9.3005
R747 VTAIL.n326 VTAIL.n325 9.3005
R748 VTAIL.n734 VTAIL.n733 8.92171
R749 VTAIL.n749 VTAIL.n702 8.92171
R750 VTAIL.n780 VTAIL.n686 8.92171
R751 VTAIL.n48 VTAIL.n47 8.92171
R752 VTAIL.n63 VTAIL.n16 8.92171
R753 VTAIL.n94 VTAIL.n0 8.92171
R754 VTAIL.n146 VTAIL.n145 8.92171
R755 VTAIL.n161 VTAIL.n114 8.92171
R756 VTAIL.n192 VTAIL.n98 8.92171
R757 VTAIL.n244 VTAIL.n243 8.92171
R758 VTAIL.n259 VTAIL.n212 8.92171
R759 VTAIL.n290 VTAIL.n196 8.92171
R760 VTAIL.n682 VTAIL.n588 8.92171
R761 VTAIL.n653 VTAIL.n606 8.92171
R762 VTAIL.n638 VTAIL.n637 8.92171
R763 VTAIL.n584 VTAIL.n490 8.92171
R764 VTAIL.n555 VTAIL.n508 8.92171
R765 VTAIL.n540 VTAIL.n539 8.92171
R766 VTAIL.n486 VTAIL.n392 8.92171
R767 VTAIL.n457 VTAIL.n410 8.92171
R768 VTAIL.n442 VTAIL.n441 8.92171
R769 VTAIL.n388 VTAIL.n294 8.92171
R770 VTAIL.n359 VTAIL.n312 8.92171
R771 VTAIL.n344 VTAIL.n343 8.92171
R772 VTAIL.n737 VTAIL.n708 8.14595
R773 VTAIL.n746 VTAIL.n745 8.14595
R774 VTAIL.n51 VTAIL.n22 8.14595
R775 VTAIL.n60 VTAIL.n59 8.14595
R776 VTAIL.n149 VTAIL.n120 8.14595
R777 VTAIL.n158 VTAIL.n157 8.14595
R778 VTAIL.n247 VTAIL.n218 8.14595
R779 VTAIL.n256 VTAIL.n255 8.14595
R780 VTAIL.n650 VTAIL.n649 8.14595
R781 VTAIL.n641 VTAIL.n612 8.14595
R782 VTAIL.n552 VTAIL.n551 8.14595
R783 VTAIL.n543 VTAIL.n514 8.14595
R784 VTAIL.n454 VTAIL.n453 8.14595
R785 VTAIL.n445 VTAIL.n416 8.14595
R786 VTAIL.n356 VTAIL.n355 8.14595
R787 VTAIL.n347 VTAIL.n318 8.14595
R788 VTAIL.n738 VTAIL.n706 7.3702
R789 VTAIL.n742 VTAIL.n704 7.3702
R790 VTAIL.n52 VTAIL.n20 7.3702
R791 VTAIL.n56 VTAIL.n18 7.3702
R792 VTAIL.n150 VTAIL.n118 7.3702
R793 VTAIL.n154 VTAIL.n116 7.3702
R794 VTAIL.n248 VTAIL.n216 7.3702
R795 VTAIL.n252 VTAIL.n214 7.3702
R796 VTAIL.n646 VTAIL.n608 7.3702
R797 VTAIL.n642 VTAIL.n610 7.3702
R798 VTAIL.n548 VTAIL.n510 7.3702
R799 VTAIL.n544 VTAIL.n512 7.3702
R800 VTAIL.n450 VTAIL.n412 7.3702
R801 VTAIL.n446 VTAIL.n414 7.3702
R802 VTAIL.n352 VTAIL.n314 7.3702
R803 VTAIL.n348 VTAIL.n316 7.3702
R804 VTAIL.n741 VTAIL.n706 6.59444
R805 VTAIL.n742 VTAIL.n741 6.59444
R806 VTAIL.n55 VTAIL.n20 6.59444
R807 VTAIL.n56 VTAIL.n55 6.59444
R808 VTAIL.n153 VTAIL.n118 6.59444
R809 VTAIL.n154 VTAIL.n153 6.59444
R810 VTAIL.n251 VTAIL.n216 6.59444
R811 VTAIL.n252 VTAIL.n251 6.59444
R812 VTAIL.n646 VTAIL.n645 6.59444
R813 VTAIL.n645 VTAIL.n610 6.59444
R814 VTAIL.n548 VTAIL.n547 6.59444
R815 VTAIL.n547 VTAIL.n512 6.59444
R816 VTAIL.n450 VTAIL.n449 6.59444
R817 VTAIL.n449 VTAIL.n414 6.59444
R818 VTAIL.n352 VTAIL.n351 6.59444
R819 VTAIL.n351 VTAIL.n316 6.59444
R820 VTAIL.n738 VTAIL.n737 5.81868
R821 VTAIL.n745 VTAIL.n704 5.81868
R822 VTAIL.n52 VTAIL.n51 5.81868
R823 VTAIL.n59 VTAIL.n18 5.81868
R824 VTAIL.n150 VTAIL.n149 5.81868
R825 VTAIL.n157 VTAIL.n116 5.81868
R826 VTAIL.n248 VTAIL.n247 5.81868
R827 VTAIL.n255 VTAIL.n214 5.81868
R828 VTAIL.n649 VTAIL.n608 5.81868
R829 VTAIL.n642 VTAIL.n641 5.81868
R830 VTAIL.n551 VTAIL.n510 5.81868
R831 VTAIL.n544 VTAIL.n543 5.81868
R832 VTAIL.n453 VTAIL.n412 5.81868
R833 VTAIL.n446 VTAIL.n445 5.81868
R834 VTAIL.n355 VTAIL.n314 5.81868
R835 VTAIL.n348 VTAIL.n347 5.81868
R836 VTAIL.n734 VTAIL.n708 5.04292
R837 VTAIL.n746 VTAIL.n702 5.04292
R838 VTAIL.n782 VTAIL.n686 5.04292
R839 VTAIL.n48 VTAIL.n22 5.04292
R840 VTAIL.n60 VTAIL.n16 5.04292
R841 VTAIL.n96 VTAIL.n0 5.04292
R842 VTAIL.n146 VTAIL.n120 5.04292
R843 VTAIL.n158 VTAIL.n114 5.04292
R844 VTAIL.n194 VTAIL.n98 5.04292
R845 VTAIL.n244 VTAIL.n218 5.04292
R846 VTAIL.n256 VTAIL.n212 5.04292
R847 VTAIL.n292 VTAIL.n196 5.04292
R848 VTAIL.n684 VTAIL.n588 5.04292
R849 VTAIL.n650 VTAIL.n606 5.04292
R850 VTAIL.n638 VTAIL.n612 5.04292
R851 VTAIL.n586 VTAIL.n490 5.04292
R852 VTAIL.n552 VTAIL.n508 5.04292
R853 VTAIL.n540 VTAIL.n514 5.04292
R854 VTAIL.n488 VTAIL.n392 5.04292
R855 VTAIL.n454 VTAIL.n410 5.04292
R856 VTAIL.n442 VTAIL.n416 5.04292
R857 VTAIL.n390 VTAIL.n294 5.04292
R858 VTAIL.n356 VTAIL.n312 5.04292
R859 VTAIL.n344 VTAIL.n318 5.04292
R860 VTAIL.n717 VTAIL.n715 4.38563
R861 VTAIL.n31 VTAIL.n29 4.38563
R862 VTAIL.n129 VTAIL.n127 4.38563
R863 VTAIL.n227 VTAIL.n225 4.38563
R864 VTAIL.n621 VTAIL.n619 4.38563
R865 VTAIL.n523 VTAIL.n521 4.38563
R866 VTAIL.n425 VTAIL.n423 4.38563
R867 VTAIL.n327 VTAIL.n325 4.38563
R868 VTAIL.n733 VTAIL.n710 4.26717
R869 VTAIL.n750 VTAIL.n749 4.26717
R870 VTAIL.n780 VTAIL.n779 4.26717
R871 VTAIL.n47 VTAIL.n24 4.26717
R872 VTAIL.n64 VTAIL.n63 4.26717
R873 VTAIL.n94 VTAIL.n93 4.26717
R874 VTAIL.n145 VTAIL.n122 4.26717
R875 VTAIL.n162 VTAIL.n161 4.26717
R876 VTAIL.n192 VTAIL.n191 4.26717
R877 VTAIL.n243 VTAIL.n220 4.26717
R878 VTAIL.n260 VTAIL.n259 4.26717
R879 VTAIL.n290 VTAIL.n289 4.26717
R880 VTAIL.n682 VTAIL.n681 4.26717
R881 VTAIL.n654 VTAIL.n653 4.26717
R882 VTAIL.n637 VTAIL.n614 4.26717
R883 VTAIL.n584 VTAIL.n583 4.26717
R884 VTAIL.n556 VTAIL.n555 4.26717
R885 VTAIL.n539 VTAIL.n516 4.26717
R886 VTAIL.n486 VTAIL.n485 4.26717
R887 VTAIL.n458 VTAIL.n457 4.26717
R888 VTAIL.n441 VTAIL.n418 4.26717
R889 VTAIL.n388 VTAIL.n387 4.26717
R890 VTAIL.n360 VTAIL.n359 4.26717
R891 VTAIL.n343 VTAIL.n320 4.26717
R892 VTAIL.n730 VTAIL.n729 3.49141
R893 VTAIL.n753 VTAIL.n700 3.49141
R894 VTAIL.n776 VTAIL.n688 3.49141
R895 VTAIL.n44 VTAIL.n43 3.49141
R896 VTAIL.n67 VTAIL.n14 3.49141
R897 VTAIL.n90 VTAIL.n2 3.49141
R898 VTAIL.n142 VTAIL.n141 3.49141
R899 VTAIL.n165 VTAIL.n112 3.49141
R900 VTAIL.n188 VTAIL.n100 3.49141
R901 VTAIL.n240 VTAIL.n239 3.49141
R902 VTAIL.n263 VTAIL.n210 3.49141
R903 VTAIL.n286 VTAIL.n198 3.49141
R904 VTAIL.n678 VTAIL.n590 3.49141
R905 VTAIL.n657 VTAIL.n604 3.49141
R906 VTAIL.n634 VTAIL.n633 3.49141
R907 VTAIL.n580 VTAIL.n492 3.49141
R908 VTAIL.n559 VTAIL.n506 3.49141
R909 VTAIL.n536 VTAIL.n535 3.49141
R910 VTAIL.n482 VTAIL.n394 3.49141
R911 VTAIL.n461 VTAIL.n408 3.49141
R912 VTAIL.n438 VTAIL.n437 3.49141
R913 VTAIL.n384 VTAIL.n296 3.49141
R914 VTAIL.n363 VTAIL.n310 3.49141
R915 VTAIL.n340 VTAIL.n339 3.49141
R916 VTAIL.n726 VTAIL.n712 2.71565
R917 VTAIL.n754 VTAIL.n698 2.71565
R918 VTAIL.n775 VTAIL.n690 2.71565
R919 VTAIL.n40 VTAIL.n26 2.71565
R920 VTAIL.n68 VTAIL.n12 2.71565
R921 VTAIL.n89 VTAIL.n4 2.71565
R922 VTAIL.n138 VTAIL.n124 2.71565
R923 VTAIL.n166 VTAIL.n110 2.71565
R924 VTAIL.n187 VTAIL.n102 2.71565
R925 VTAIL.n236 VTAIL.n222 2.71565
R926 VTAIL.n264 VTAIL.n208 2.71565
R927 VTAIL.n285 VTAIL.n200 2.71565
R928 VTAIL.n677 VTAIL.n592 2.71565
R929 VTAIL.n658 VTAIL.n602 2.71565
R930 VTAIL.n630 VTAIL.n616 2.71565
R931 VTAIL.n579 VTAIL.n494 2.71565
R932 VTAIL.n560 VTAIL.n504 2.71565
R933 VTAIL.n532 VTAIL.n518 2.71565
R934 VTAIL.n481 VTAIL.n396 2.71565
R935 VTAIL.n462 VTAIL.n406 2.71565
R936 VTAIL.n434 VTAIL.n420 2.71565
R937 VTAIL.n383 VTAIL.n298 2.71565
R938 VTAIL.n364 VTAIL.n308 2.71565
R939 VTAIL.n336 VTAIL.n322 2.71565
R940 VTAIL.n725 VTAIL.n714 1.93989
R941 VTAIL.n759 VTAIL.n757 1.93989
R942 VTAIL.n772 VTAIL.n771 1.93989
R943 VTAIL.n39 VTAIL.n28 1.93989
R944 VTAIL.n73 VTAIL.n71 1.93989
R945 VTAIL.n86 VTAIL.n85 1.93989
R946 VTAIL.n137 VTAIL.n126 1.93989
R947 VTAIL.n171 VTAIL.n169 1.93989
R948 VTAIL.n184 VTAIL.n183 1.93989
R949 VTAIL.n235 VTAIL.n224 1.93989
R950 VTAIL.n269 VTAIL.n267 1.93989
R951 VTAIL.n282 VTAIL.n281 1.93989
R952 VTAIL.n674 VTAIL.n673 1.93989
R953 VTAIL.n662 VTAIL.n661 1.93989
R954 VTAIL.n629 VTAIL.n618 1.93989
R955 VTAIL.n576 VTAIL.n575 1.93989
R956 VTAIL.n564 VTAIL.n563 1.93989
R957 VTAIL.n531 VTAIL.n520 1.93989
R958 VTAIL.n478 VTAIL.n477 1.93989
R959 VTAIL.n466 VTAIL.n465 1.93989
R960 VTAIL.n433 VTAIL.n422 1.93989
R961 VTAIL.n380 VTAIL.n379 1.93989
R962 VTAIL.n368 VTAIL.n367 1.93989
R963 VTAIL.n335 VTAIL.n324 1.93989
R964 VTAIL.n722 VTAIL.n721 1.16414
R965 VTAIL.n758 VTAIL.n696 1.16414
R966 VTAIL.n768 VTAIL.n692 1.16414
R967 VTAIL.n36 VTAIL.n35 1.16414
R968 VTAIL.n72 VTAIL.n10 1.16414
R969 VTAIL.n82 VTAIL.n6 1.16414
R970 VTAIL.n134 VTAIL.n133 1.16414
R971 VTAIL.n170 VTAIL.n108 1.16414
R972 VTAIL.n180 VTAIL.n104 1.16414
R973 VTAIL.n232 VTAIL.n231 1.16414
R974 VTAIL.n268 VTAIL.n206 1.16414
R975 VTAIL.n278 VTAIL.n202 1.16414
R976 VTAIL.n670 VTAIL.n594 1.16414
R977 VTAIL.n665 VTAIL.n599 1.16414
R978 VTAIL.n626 VTAIL.n625 1.16414
R979 VTAIL.n572 VTAIL.n496 1.16414
R980 VTAIL.n567 VTAIL.n501 1.16414
R981 VTAIL.n528 VTAIL.n527 1.16414
R982 VTAIL.n474 VTAIL.n398 1.16414
R983 VTAIL.n469 VTAIL.n403 1.16414
R984 VTAIL.n430 VTAIL.n429 1.16414
R985 VTAIL.n376 VTAIL.n300 1.16414
R986 VTAIL.n371 VTAIL.n305 1.16414
R987 VTAIL.n332 VTAIL.n331 1.16414
R988 VTAIL.n489 VTAIL.n391 0.759121
R989 VTAIL.n685 VTAIL.n587 0.759121
R990 VTAIL.n293 VTAIL.n195 0.759121
R991 VTAIL.n587 VTAIL.n489 0.470328
R992 VTAIL.n195 VTAIL.n97 0.470328
R993 VTAIL VTAIL.n97 0.438
R994 VTAIL.n718 VTAIL.n716 0.388379
R995 VTAIL.n764 VTAIL.n763 0.388379
R996 VTAIL.n767 VTAIL.n694 0.388379
R997 VTAIL.n32 VTAIL.n30 0.388379
R998 VTAIL.n78 VTAIL.n77 0.388379
R999 VTAIL.n81 VTAIL.n8 0.388379
R1000 VTAIL.n130 VTAIL.n128 0.388379
R1001 VTAIL.n176 VTAIL.n175 0.388379
R1002 VTAIL.n179 VTAIL.n106 0.388379
R1003 VTAIL.n228 VTAIL.n226 0.388379
R1004 VTAIL.n274 VTAIL.n273 0.388379
R1005 VTAIL.n277 VTAIL.n204 0.388379
R1006 VTAIL.n669 VTAIL.n596 0.388379
R1007 VTAIL.n666 VTAIL.n598 0.388379
R1008 VTAIL.n622 VTAIL.n620 0.388379
R1009 VTAIL.n571 VTAIL.n498 0.388379
R1010 VTAIL.n568 VTAIL.n500 0.388379
R1011 VTAIL.n524 VTAIL.n522 0.388379
R1012 VTAIL.n473 VTAIL.n400 0.388379
R1013 VTAIL.n470 VTAIL.n402 0.388379
R1014 VTAIL.n426 VTAIL.n424 0.388379
R1015 VTAIL.n375 VTAIL.n302 0.388379
R1016 VTAIL.n372 VTAIL.n304 0.388379
R1017 VTAIL.n328 VTAIL.n326 0.388379
R1018 VTAIL VTAIL.n783 0.321621
R1019 VTAIL.n723 VTAIL.n715 0.155672
R1020 VTAIL.n724 VTAIL.n723 0.155672
R1021 VTAIL.n724 VTAIL.n711 0.155672
R1022 VTAIL.n731 VTAIL.n711 0.155672
R1023 VTAIL.n732 VTAIL.n731 0.155672
R1024 VTAIL.n732 VTAIL.n707 0.155672
R1025 VTAIL.n739 VTAIL.n707 0.155672
R1026 VTAIL.n740 VTAIL.n739 0.155672
R1027 VTAIL.n740 VTAIL.n703 0.155672
R1028 VTAIL.n747 VTAIL.n703 0.155672
R1029 VTAIL.n748 VTAIL.n747 0.155672
R1030 VTAIL.n748 VTAIL.n699 0.155672
R1031 VTAIL.n755 VTAIL.n699 0.155672
R1032 VTAIL.n756 VTAIL.n755 0.155672
R1033 VTAIL.n756 VTAIL.n695 0.155672
R1034 VTAIL.n765 VTAIL.n695 0.155672
R1035 VTAIL.n766 VTAIL.n765 0.155672
R1036 VTAIL.n766 VTAIL.n691 0.155672
R1037 VTAIL.n773 VTAIL.n691 0.155672
R1038 VTAIL.n774 VTAIL.n773 0.155672
R1039 VTAIL.n774 VTAIL.n687 0.155672
R1040 VTAIL.n781 VTAIL.n687 0.155672
R1041 VTAIL.n37 VTAIL.n29 0.155672
R1042 VTAIL.n38 VTAIL.n37 0.155672
R1043 VTAIL.n38 VTAIL.n25 0.155672
R1044 VTAIL.n45 VTAIL.n25 0.155672
R1045 VTAIL.n46 VTAIL.n45 0.155672
R1046 VTAIL.n46 VTAIL.n21 0.155672
R1047 VTAIL.n53 VTAIL.n21 0.155672
R1048 VTAIL.n54 VTAIL.n53 0.155672
R1049 VTAIL.n54 VTAIL.n17 0.155672
R1050 VTAIL.n61 VTAIL.n17 0.155672
R1051 VTAIL.n62 VTAIL.n61 0.155672
R1052 VTAIL.n62 VTAIL.n13 0.155672
R1053 VTAIL.n69 VTAIL.n13 0.155672
R1054 VTAIL.n70 VTAIL.n69 0.155672
R1055 VTAIL.n70 VTAIL.n9 0.155672
R1056 VTAIL.n79 VTAIL.n9 0.155672
R1057 VTAIL.n80 VTAIL.n79 0.155672
R1058 VTAIL.n80 VTAIL.n5 0.155672
R1059 VTAIL.n87 VTAIL.n5 0.155672
R1060 VTAIL.n88 VTAIL.n87 0.155672
R1061 VTAIL.n88 VTAIL.n1 0.155672
R1062 VTAIL.n95 VTAIL.n1 0.155672
R1063 VTAIL.n135 VTAIL.n127 0.155672
R1064 VTAIL.n136 VTAIL.n135 0.155672
R1065 VTAIL.n136 VTAIL.n123 0.155672
R1066 VTAIL.n143 VTAIL.n123 0.155672
R1067 VTAIL.n144 VTAIL.n143 0.155672
R1068 VTAIL.n144 VTAIL.n119 0.155672
R1069 VTAIL.n151 VTAIL.n119 0.155672
R1070 VTAIL.n152 VTAIL.n151 0.155672
R1071 VTAIL.n152 VTAIL.n115 0.155672
R1072 VTAIL.n159 VTAIL.n115 0.155672
R1073 VTAIL.n160 VTAIL.n159 0.155672
R1074 VTAIL.n160 VTAIL.n111 0.155672
R1075 VTAIL.n167 VTAIL.n111 0.155672
R1076 VTAIL.n168 VTAIL.n167 0.155672
R1077 VTAIL.n168 VTAIL.n107 0.155672
R1078 VTAIL.n177 VTAIL.n107 0.155672
R1079 VTAIL.n178 VTAIL.n177 0.155672
R1080 VTAIL.n178 VTAIL.n103 0.155672
R1081 VTAIL.n185 VTAIL.n103 0.155672
R1082 VTAIL.n186 VTAIL.n185 0.155672
R1083 VTAIL.n186 VTAIL.n99 0.155672
R1084 VTAIL.n193 VTAIL.n99 0.155672
R1085 VTAIL.n233 VTAIL.n225 0.155672
R1086 VTAIL.n234 VTAIL.n233 0.155672
R1087 VTAIL.n234 VTAIL.n221 0.155672
R1088 VTAIL.n241 VTAIL.n221 0.155672
R1089 VTAIL.n242 VTAIL.n241 0.155672
R1090 VTAIL.n242 VTAIL.n217 0.155672
R1091 VTAIL.n249 VTAIL.n217 0.155672
R1092 VTAIL.n250 VTAIL.n249 0.155672
R1093 VTAIL.n250 VTAIL.n213 0.155672
R1094 VTAIL.n257 VTAIL.n213 0.155672
R1095 VTAIL.n258 VTAIL.n257 0.155672
R1096 VTAIL.n258 VTAIL.n209 0.155672
R1097 VTAIL.n265 VTAIL.n209 0.155672
R1098 VTAIL.n266 VTAIL.n265 0.155672
R1099 VTAIL.n266 VTAIL.n205 0.155672
R1100 VTAIL.n275 VTAIL.n205 0.155672
R1101 VTAIL.n276 VTAIL.n275 0.155672
R1102 VTAIL.n276 VTAIL.n201 0.155672
R1103 VTAIL.n283 VTAIL.n201 0.155672
R1104 VTAIL.n284 VTAIL.n283 0.155672
R1105 VTAIL.n284 VTAIL.n197 0.155672
R1106 VTAIL.n291 VTAIL.n197 0.155672
R1107 VTAIL.n683 VTAIL.n589 0.155672
R1108 VTAIL.n676 VTAIL.n589 0.155672
R1109 VTAIL.n676 VTAIL.n675 0.155672
R1110 VTAIL.n675 VTAIL.n593 0.155672
R1111 VTAIL.n668 VTAIL.n593 0.155672
R1112 VTAIL.n668 VTAIL.n667 0.155672
R1113 VTAIL.n667 VTAIL.n597 0.155672
R1114 VTAIL.n660 VTAIL.n597 0.155672
R1115 VTAIL.n660 VTAIL.n659 0.155672
R1116 VTAIL.n659 VTAIL.n603 0.155672
R1117 VTAIL.n652 VTAIL.n603 0.155672
R1118 VTAIL.n652 VTAIL.n651 0.155672
R1119 VTAIL.n651 VTAIL.n607 0.155672
R1120 VTAIL.n644 VTAIL.n607 0.155672
R1121 VTAIL.n644 VTAIL.n643 0.155672
R1122 VTAIL.n643 VTAIL.n611 0.155672
R1123 VTAIL.n636 VTAIL.n611 0.155672
R1124 VTAIL.n636 VTAIL.n635 0.155672
R1125 VTAIL.n635 VTAIL.n615 0.155672
R1126 VTAIL.n628 VTAIL.n615 0.155672
R1127 VTAIL.n628 VTAIL.n627 0.155672
R1128 VTAIL.n627 VTAIL.n619 0.155672
R1129 VTAIL.n585 VTAIL.n491 0.155672
R1130 VTAIL.n578 VTAIL.n491 0.155672
R1131 VTAIL.n578 VTAIL.n577 0.155672
R1132 VTAIL.n577 VTAIL.n495 0.155672
R1133 VTAIL.n570 VTAIL.n495 0.155672
R1134 VTAIL.n570 VTAIL.n569 0.155672
R1135 VTAIL.n569 VTAIL.n499 0.155672
R1136 VTAIL.n562 VTAIL.n499 0.155672
R1137 VTAIL.n562 VTAIL.n561 0.155672
R1138 VTAIL.n561 VTAIL.n505 0.155672
R1139 VTAIL.n554 VTAIL.n505 0.155672
R1140 VTAIL.n554 VTAIL.n553 0.155672
R1141 VTAIL.n553 VTAIL.n509 0.155672
R1142 VTAIL.n546 VTAIL.n509 0.155672
R1143 VTAIL.n546 VTAIL.n545 0.155672
R1144 VTAIL.n545 VTAIL.n513 0.155672
R1145 VTAIL.n538 VTAIL.n513 0.155672
R1146 VTAIL.n538 VTAIL.n537 0.155672
R1147 VTAIL.n537 VTAIL.n517 0.155672
R1148 VTAIL.n530 VTAIL.n517 0.155672
R1149 VTAIL.n530 VTAIL.n529 0.155672
R1150 VTAIL.n529 VTAIL.n521 0.155672
R1151 VTAIL.n487 VTAIL.n393 0.155672
R1152 VTAIL.n480 VTAIL.n393 0.155672
R1153 VTAIL.n480 VTAIL.n479 0.155672
R1154 VTAIL.n479 VTAIL.n397 0.155672
R1155 VTAIL.n472 VTAIL.n397 0.155672
R1156 VTAIL.n472 VTAIL.n471 0.155672
R1157 VTAIL.n471 VTAIL.n401 0.155672
R1158 VTAIL.n464 VTAIL.n401 0.155672
R1159 VTAIL.n464 VTAIL.n463 0.155672
R1160 VTAIL.n463 VTAIL.n407 0.155672
R1161 VTAIL.n456 VTAIL.n407 0.155672
R1162 VTAIL.n456 VTAIL.n455 0.155672
R1163 VTAIL.n455 VTAIL.n411 0.155672
R1164 VTAIL.n448 VTAIL.n411 0.155672
R1165 VTAIL.n448 VTAIL.n447 0.155672
R1166 VTAIL.n447 VTAIL.n415 0.155672
R1167 VTAIL.n440 VTAIL.n415 0.155672
R1168 VTAIL.n440 VTAIL.n439 0.155672
R1169 VTAIL.n439 VTAIL.n419 0.155672
R1170 VTAIL.n432 VTAIL.n419 0.155672
R1171 VTAIL.n432 VTAIL.n431 0.155672
R1172 VTAIL.n431 VTAIL.n423 0.155672
R1173 VTAIL.n389 VTAIL.n295 0.155672
R1174 VTAIL.n382 VTAIL.n295 0.155672
R1175 VTAIL.n382 VTAIL.n381 0.155672
R1176 VTAIL.n381 VTAIL.n299 0.155672
R1177 VTAIL.n374 VTAIL.n299 0.155672
R1178 VTAIL.n374 VTAIL.n373 0.155672
R1179 VTAIL.n373 VTAIL.n303 0.155672
R1180 VTAIL.n366 VTAIL.n303 0.155672
R1181 VTAIL.n366 VTAIL.n365 0.155672
R1182 VTAIL.n365 VTAIL.n309 0.155672
R1183 VTAIL.n358 VTAIL.n309 0.155672
R1184 VTAIL.n358 VTAIL.n357 0.155672
R1185 VTAIL.n357 VTAIL.n313 0.155672
R1186 VTAIL.n350 VTAIL.n313 0.155672
R1187 VTAIL.n350 VTAIL.n349 0.155672
R1188 VTAIL.n349 VTAIL.n317 0.155672
R1189 VTAIL.n342 VTAIL.n317 0.155672
R1190 VTAIL.n342 VTAIL.n341 0.155672
R1191 VTAIL.n341 VTAIL.n321 0.155672
R1192 VTAIL.n334 VTAIL.n321 0.155672
R1193 VTAIL.n334 VTAIL.n333 0.155672
R1194 VTAIL.n333 VTAIL.n325 0.155672
R1195 VDD1 VDD1.n1 100.073
R1196 VDD1 VDD1.n0 58.6068
R1197 VDD1.n0 VDD1.t0 1.13778
R1198 VDD1.n0 VDD1.t3 1.13778
R1199 VDD1.n1 VDD1.t2 1.13778
R1200 VDD1.n1 VDD1.t1 1.13778
R1201 B.n407 B.t4 968.188
R1202 B.n555 B.t15 968.188
R1203 B.n99 B.t12 968.188
R1204 B.n97 B.t8 968.188
R1205 B.n766 B.n765 585
R1206 B.n767 B.n766 585
R1207 B.n347 B.n96 585
R1208 B.n346 B.n345 585
R1209 B.n344 B.n343 585
R1210 B.n342 B.n341 585
R1211 B.n340 B.n339 585
R1212 B.n338 B.n337 585
R1213 B.n336 B.n335 585
R1214 B.n334 B.n333 585
R1215 B.n332 B.n331 585
R1216 B.n330 B.n329 585
R1217 B.n328 B.n327 585
R1218 B.n326 B.n325 585
R1219 B.n324 B.n323 585
R1220 B.n322 B.n321 585
R1221 B.n320 B.n319 585
R1222 B.n318 B.n317 585
R1223 B.n316 B.n315 585
R1224 B.n314 B.n313 585
R1225 B.n312 B.n311 585
R1226 B.n310 B.n309 585
R1227 B.n308 B.n307 585
R1228 B.n306 B.n305 585
R1229 B.n304 B.n303 585
R1230 B.n302 B.n301 585
R1231 B.n300 B.n299 585
R1232 B.n298 B.n297 585
R1233 B.n296 B.n295 585
R1234 B.n294 B.n293 585
R1235 B.n292 B.n291 585
R1236 B.n290 B.n289 585
R1237 B.n288 B.n287 585
R1238 B.n286 B.n285 585
R1239 B.n284 B.n283 585
R1240 B.n282 B.n281 585
R1241 B.n280 B.n279 585
R1242 B.n278 B.n277 585
R1243 B.n276 B.n275 585
R1244 B.n274 B.n273 585
R1245 B.n272 B.n271 585
R1246 B.n270 B.n269 585
R1247 B.n268 B.n267 585
R1248 B.n266 B.n265 585
R1249 B.n264 B.n263 585
R1250 B.n262 B.n261 585
R1251 B.n260 B.n259 585
R1252 B.n258 B.n257 585
R1253 B.n256 B.n255 585
R1254 B.n254 B.n253 585
R1255 B.n252 B.n251 585
R1256 B.n250 B.n249 585
R1257 B.n248 B.n247 585
R1258 B.n246 B.n245 585
R1259 B.n244 B.n243 585
R1260 B.n242 B.n241 585
R1261 B.n240 B.n239 585
R1262 B.n238 B.n237 585
R1263 B.n236 B.n235 585
R1264 B.n233 B.n232 585
R1265 B.n231 B.n230 585
R1266 B.n229 B.n228 585
R1267 B.n227 B.n226 585
R1268 B.n225 B.n224 585
R1269 B.n223 B.n222 585
R1270 B.n221 B.n220 585
R1271 B.n219 B.n218 585
R1272 B.n217 B.n216 585
R1273 B.n215 B.n214 585
R1274 B.n213 B.n212 585
R1275 B.n211 B.n210 585
R1276 B.n209 B.n208 585
R1277 B.n207 B.n206 585
R1278 B.n205 B.n204 585
R1279 B.n203 B.n202 585
R1280 B.n201 B.n200 585
R1281 B.n199 B.n198 585
R1282 B.n197 B.n196 585
R1283 B.n195 B.n194 585
R1284 B.n193 B.n192 585
R1285 B.n191 B.n190 585
R1286 B.n189 B.n188 585
R1287 B.n187 B.n186 585
R1288 B.n185 B.n184 585
R1289 B.n183 B.n182 585
R1290 B.n181 B.n180 585
R1291 B.n179 B.n178 585
R1292 B.n177 B.n176 585
R1293 B.n175 B.n174 585
R1294 B.n173 B.n172 585
R1295 B.n171 B.n170 585
R1296 B.n169 B.n168 585
R1297 B.n167 B.n166 585
R1298 B.n165 B.n164 585
R1299 B.n163 B.n162 585
R1300 B.n161 B.n160 585
R1301 B.n159 B.n158 585
R1302 B.n157 B.n156 585
R1303 B.n155 B.n154 585
R1304 B.n153 B.n152 585
R1305 B.n151 B.n150 585
R1306 B.n149 B.n148 585
R1307 B.n147 B.n146 585
R1308 B.n145 B.n144 585
R1309 B.n143 B.n142 585
R1310 B.n141 B.n140 585
R1311 B.n139 B.n138 585
R1312 B.n137 B.n136 585
R1313 B.n135 B.n134 585
R1314 B.n133 B.n132 585
R1315 B.n131 B.n130 585
R1316 B.n129 B.n128 585
R1317 B.n127 B.n126 585
R1318 B.n125 B.n124 585
R1319 B.n123 B.n122 585
R1320 B.n121 B.n120 585
R1321 B.n119 B.n118 585
R1322 B.n117 B.n116 585
R1323 B.n115 B.n114 585
R1324 B.n113 B.n112 585
R1325 B.n111 B.n110 585
R1326 B.n109 B.n108 585
R1327 B.n107 B.n106 585
R1328 B.n105 B.n104 585
R1329 B.n103 B.n102 585
R1330 B.n32 B.n31 585
R1331 B.n764 B.n33 585
R1332 B.n768 B.n33 585
R1333 B.n763 B.n762 585
R1334 B.n762 B.n29 585
R1335 B.n761 B.n28 585
R1336 B.n774 B.n28 585
R1337 B.n760 B.n27 585
R1338 B.n775 B.n27 585
R1339 B.n759 B.n26 585
R1340 B.n776 B.n26 585
R1341 B.n758 B.n757 585
R1342 B.n757 B.n22 585
R1343 B.n756 B.n21 585
R1344 B.n782 B.n21 585
R1345 B.n755 B.n20 585
R1346 B.n783 B.n20 585
R1347 B.n754 B.n19 585
R1348 B.n784 B.n19 585
R1349 B.n753 B.n752 585
R1350 B.n752 B.n15 585
R1351 B.n751 B.n14 585
R1352 B.n790 B.n14 585
R1353 B.n750 B.n13 585
R1354 B.n791 B.n13 585
R1355 B.n749 B.n12 585
R1356 B.n792 B.n12 585
R1357 B.n748 B.n747 585
R1358 B.n747 B.n11 585
R1359 B.n746 B.n7 585
R1360 B.n798 B.n7 585
R1361 B.n745 B.n6 585
R1362 B.n799 B.n6 585
R1363 B.n744 B.n5 585
R1364 B.n800 B.n5 585
R1365 B.n743 B.n742 585
R1366 B.n742 B.n4 585
R1367 B.n741 B.n348 585
R1368 B.n741 B.n740 585
R1369 B.n730 B.n349 585
R1370 B.n733 B.n349 585
R1371 B.n732 B.n731 585
R1372 B.n734 B.n732 585
R1373 B.n729 B.n354 585
R1374 B.n354 B.n353 585
R1375 B.n728 B.n727 585
R1376 B.n727 B.n726 585
R1377 B.n356 B.n355 585
R1378 B.n357 B.n356 585
R1379 B.n719 B.n718 585
R1380 B.n720 B.n719 585
R1381 B.n717 B.n362 585
R1382 B.n362 B.n361 585
R1383 B.n716 B.n715 585
R1384 B.n715 B.n714 585
R1385 B.n364 B.n363 585
R1386 B.n365 B.n364 585
R1387 B.n707 B.n706 585
R1388 B.n708 B.n707 585
R1389 B.n705 B.n370 585
R1390 B.n370 B.n369 585
R1391 B.n704 B.n703 585
R1392 B.n703 B.n702 585
R1393 B.n372 B.n371 585
R1394 B.n373 B.n372 585
R1395 B.n695 B.n694 585
R1396 B.n696 B.n695 585
R1397 B.n376 B.n375 585
R1398 B.n445 B.n443 585
R1399 B.n446 B.n442 585
R1400 B.n446 B.n377 585
R1401 B.n449 B.n448 585
R1402 B.n450 B.n441 585
R1403 B.n452 B.n451 585
R1404 B.n454 B.n440 585
R1405 B.n457 B.n456 585
R1406 B.n458 B.n439 585
R1407 B.n460 B.n459 585
R1408 B.n462 B.n438 585
R1409 B.n465 B.n464 585
R1410 B.n466 B.n437 585
R1411 B.n468 B.n467 585
R1412 B.n470 B.n436 585
R1413 B.n473 B.n472 585
R1414 B.n474 B.n435 585
R1415 B.n476 B.n475 585
R1416 B.n478 B.n434 585
R1417 B.n481 B.n480 585
R1418 B.n482 B.n433 585
R1419 B.n484 B.n483 585
R1420 B.n486 B.n432 585
R1421 B.n489 B.n488 585
R1422 B.n490 B.n431 585
R1423 B.n492 B.n491 585
R1424 B.n494 B.n430 585
R1425 B.n497 B.n496 585
R1426 B.n498 B.n429 585
R1427 B.n500 B.n499 585
R1428 B.n502 B.n428 585
R1429 B.n505 B.n504 585
R1430 B.n506 B.n427 585
R1431 B.n508 B.n507 585
R1432 B.n510 B.n426 585
R1433 B.n513 B.n512 585
R1434 B.n514 B.n425 585
R1435 B.n516 B.n515 585
R1436 B.n518 B.n424 585
R1437 B.n521 B.n520 585
R1438 B.n522 B.n423 585
R1439 B.n524 B.n523 585
R1440 B.n526 B.n422 585
R1441 B.n529 B.n528 585
R1442 B.n530 B.n421 585
R1443 B.n532 B.n531 585
R1444 B.n534 B.n420 585
R1445 B.n537 B.n536 585
R1446 B.n538 B.n419 585
R1447 B.n540 B.n539 585
R1448 B.n542 B.n418 585
R1449 B.n545 B.n544 585
R1450 B.n546 B.n417 585
R1451 B.n548 B.n547 585
R1452 B.n550 B.n416 585
R1453 B.n553 B.n552 585
R1454 B.n554 B.n415 585
R1455 B.n559 B.n558 585
R1456 B.n561 B.n414 585
R1457 B.n564 B.n563 585
R1458 B.n565 B.n413 585
R1459 B.n567 B.n566 585
R1460 B.n569 B.n412 585
R1461 B.n572 B.n571 585
R1462 B.n573 B.n411 585
R1463 B.n575 B.n574 585
R1464 B.n577 B.n410 585
R1465 B.n580 B.n579 585
R1466 B.n581 B.n406 585
R1467 B.n583 B.n582 585
R1468 B.n585 B.n405 585
R1469 B.n588 B.n587 585
R1470 B.n589 B.n404 585
R1471 B.n591 B.n590 585
R1472 B.n593 B.n403 585
R1473 B.n596 B.n595 585
R1474 B.n597 B.n402 585
R1475 B.n599 B.n598 585
R1476 B.n601 B.n401 585
R1477 B.n604 B.n603 585
R1478 B.n605 B.n400 585
R1479 B.n607 B.n606 585
R1480 B.n609 B.n399 585
R1481 B.n612 B.n611 585
R1482 B.n613 B.n398 585
R1483 B.n615 B.n614 585
R1484 B.n617 B.n397 585
R1485 B.n620 B.n619 585
R1486 B.n621 B.n396 585
R1487 B.n623 B.n622 585
R1488 B.n625 B.n395 585
R1489 B.n628 B.n627 585
R1490 B.n629 B.n394 585
R1491 B.n631 B.n630 585
R1492 B.n633 B.n393 585
R1493 B.n636 B.n635 585
R1494 B.n637 B.n392 585
R1495 B.n639 B.n638 585
R1496 B.n641 B.n391 585
R1497 B.n644 B.n643 585
R1498 B.n645 B.n390 585
R1499 B.n647 B.n646 585
R1500 B.n649 B.n389 585
R1501 B.n652 B.n651 585
R1502 B.n653 B.n388 585
R1503 B.n655 B.n654 585
R1504 B.n657 B.n387 585
R1505 B.n660 B.n659 585
R1506 B.n661 B.n386 585
R1507 B.n663 B.n662 585
R1508 B.n665 B.n385 585
R1509 B.n668 B.n667 585
R1510 B.n669 B.n384 585
R1511 B.n671 B.n670 585
R1512 B.n673 B.n383 585
R1513 B.n676 B.n675 585
R1514 B.n677 B.n382 585
R1515 B.n679 B.n678 585
R1516 B.n681 B.n381 585
R1517 B.n684 B.n683 585
R1518 B.n685 B.n380 585
R1519 B.n687 B.n686 585
R1520 B.n689 B.n379 585
R1521 B.n692 B.n691 585
R1522 B.n693 B.n378 585
R1523 B.n698 B.n697 585
R1524 B.n697 B.n696 585
R1525 B.n699 B.n374 585
R1526 B.n374 B.n373 585
R1527 B.n701 B.n700 585
R1528 B.n702 B.n701 585
R1529 B.n368 B.n367 585
R1530 B.n369 B.n368 585
R1531 B.n710 B.n709 585
R1532 B.n709 B.n708 585
R1533 B.n711 B.n366 585
R1534 B.n366 B.n365 585
R1535 B.n713 B.n712 585
R1536 B.n714 B.n713 585
R1537 B.n360 B.n359 585
R1538 B.n361 B.n360 585
R1539 B.n722 B.n721 585
R1540 B.n721 B.n720 585
R1541 B.n723 B.n358 585
R1542 B.n358 B.n357 585
R1543 B.n725 B.n724 585
R1544 B.n726 B.n725 585
R1545 B.n352 B.n351 585
R1546 B.n353 B.n352 585
R1547 B.n736 B.n735 585
R1548 B.n735 B.n734 585
R1549 B.n737 B.n350 585
R1550 B.n733 B.n350 585
R1551 B.n739 B.n738 585
R1552 B.n740 B.n739 585
R1553 B.n2 B.n0 585
R1554 B.n4 B.n2 585
R1555 B.n3 B.n1 585
R1556 B.n799 B.n3 585
R1557 B.n797 B.n796 585
R1558 B.n798 B.n797 585
R1559 B.n795 B.n8 585
R1560 B.n11 B.n8 585
R1561 B.n794 B.n793 585
R1562 B.n793 B.n792 585
R1563 B.n10 B.n9 585
R1564 B.n791 B.n10 585
R1565 B.n789 B.n788 585
R1566 B.n790 B.n789 585
R1567 B.n787 B.n16 585
R1568 B.n16 B.n15 585
R1569 B.n786 B.n785 585
R1570 B.n785 B.n784 585
R1571 B.n18 B.n17 585
R1572 B.n783 B.n18 585
R1573 B.n781 B.n780 585
R1574 B.n782 B.n781 585
R1575 B.n779 B.n23 585
R1576 B.n23 B.n22 585
R1577 B.n778 B.n777 585
R1578 B.n777 B.n776 585
R1579 B.n25 B.n24 585
R1580 B.n775 B.n25 585
R1581 B.n773 B.n772 585
R1582 B.n774 B.n773 585
R1583 B.n771 B.n30 585
R1584 B.n30 B.n29 585
R1585 B.n770 B.n769 585
R1586 B.n769 B.n768 585
R1587 B.n802 B.n801 585
R1588 B.n801 B.n800 585
R1589 B.n697 B.n376 449.257
R1590 B.n769 B.n32 449.257
R1591 B.n695 B.n378 449.257
R1592 B.n766 B.n33 449.257
R1593 B.n407 B.t7 392.192
R1594 B.n97 B.t10 392.192
R1595 B.n555 B.t17 392.192
R1596 B.n99 B.t13 392.192
R1597 B.n408 B.t6 375.125
R1598 B.n98 B.t11 375.125
R1599 B.n556 B.t16 375.125
R1600 B.n100 B.t14 375.125
R1601 B.n767 B.n95 256.663
R1602 B.n767 B.n94 256.663
R1603 B.n767 B.n93 256.663
R1604 B.n767 B.n92 256.663
R1605 B.n767 B.n91 256.663
R1606 B.n767 B.n90 256.663
R1607 B.n767 B.n89 256.663
R1608 B.n767 B.n88 256.663
R1609 B.n767 B.n87 256.663
R1610 B.n767 B.n86 256.663
R1611 B.n767 B.n85 256.663
R1612 B.n767 B.n84 256.663
R1613 B.n767 B.n83 256.663
R1614 B.n767 B.n82 256.663
R1615 B.n767 B.n81 256.663
R1616 B.n767 B.n80 256.663
R1617 B.n767 B.n79 256.663
R1618 B.n767 B.n78 256.663
R1619 B.n767 B.n77 256.663
R1620 B.n767 B.n76 256.663
R1621 B.n767 B.n75 256.663
R1622 B.n767 B.n74 256.663
R1623 B.n767 B.n73 256.663
R1624 B.n767 B.n72 256.663
R1625 B.n767 B.n71 256.663
R1626 B.n767 B.n70 256.663
R1627 B.n767 B.n69 256.663
R1628 B.n767 B.n68 256.663
R1629 B.n767 B.n67 256.663
R1630 B.n767 B.n66 256.663
R1631 B.n767 B.n65 256.663
R1632 B.n767 B.n64 256.663
R1633 B.n767 B.n63 256.663
R1634 B.n767 B.n62 256.663
R1635 B.n767 B.n61 256.663
R1636 B.n767 B.n60 256.663
R1637 B.n767 B.n59 256.663
R1638 B.n767 B.n58 256.663
R1639 B.n767 B.n57 256.663
R1640 B.n767 B.n56 256.663
R1641 B.n767 B.n55 256.663
R1642 B.n767 B.n54 256.663
R1643 B.n767 B.n53 256.663
R1644 B.n767 B.n52 256.663
R1645 B.n767 B.n51 256.663
R1646 B.n767 B.n50 256.663
R1647 B.n767 B.n49 256.663
R1648 B.n767 B.n48 256.663
R1649 B.n767 B.n47 256.663
R1650 B.n767 B.n46 256.663
R1651 B.n767 B.n45 256.663
R1652 B.n767 B.n44 256.663
R1653 B.n767 B.n43 256.663
R1654 B.n767 B.n42 256.663
R1655 B.n767 B.n41 256.663
R1656 B.n767 B.n40 256.663
R1657 B.n767 B.n39 256.663
R1658 B.n767 B.n38 256.663
R1659 B.n767 B.n37 256.663
R1660 B.n767 B.n36 256.663
R1661 B.n767 B.n35 256.663
R1662 B.n767 B.n34 256.663
R1663 B.n444 B.n377 256.663
R1664 B.n447 B.n377 256.663
R1665 B.n453 B.n377 256.663
R1666 B.n455 B.n377 256.663
R1667 B.n461 B.n377 256.663
R1668 B.n463 B.n377 256.663
R1669 B.n469 B.n377 256.663
R1670 B.n471 B.n377 256.663
R1671 B.n477 B.n377 256.663
R1672 B.n479 B.n377 256.663
R1673 B.n485 B.n377 256.663
R1674 B.n487 B.n377 256.663
R1675 B.n493 B.n377 256.663
R1676 B.n495 B.n377 256.663
R1677 B.n501 B.n377 256.663
R1678 B.n503 B.n377 256.663
R1679 B.n509 B.n377 256.663
R1680 B.n511 B.n377 256.663
R1681 B.n517 B.n377 256.663
R1682 B.n519 B.n377 256.663
R1683 B.n525 B.n377 256.663
R1684 B.n527 B.n377 256.663
R1685 B.n533 B.n377 256.663
R1686 B.n535 B.n377 256.663
R1687 B.n541 B.n377 256.663
R1688 B.n543 B.n377 256.663
R1689 B.n549 B.n377 256.663
R1690 B.n551 B.n377 256.663
R1691 B.n560 B.n377 256.663
R1692 B.n562 B.n377 256.663
R1693 B.n568 B.n377 256.663
R1694 B.n570 B.n377 256.663
R1695 B.n576 B.n377 256.663
R1696 B.n578 B.n377 256.663
R1697 B.n584 B.n377 256.663
R1698 B.n586 B.n377 256.663
R1699 B.n592 B.n377 256.663
R1700 B.n594 B.n377 256.663
R1701 B.n600 B.n377 256.663
R1702 B.n602 B.n377 256.663
R1703 B.n608 B.n377 256.663
R1704 B.n610 B.n377 256.663
R1705 B.n616 B.n377 256.663
R1706 B.n618 B.n377 256.663
R1707 B.n624 B.n377 256.663
R1708 B.n626 B.n377 256.663
R1709 B.n632 B.n377 256.663
R1710 B.n634 B.n377 256.663
R1711 B.n640 B.n377 256.663
R1712 B.n642 B.n377 256.663
R1713 B.n648 B.n377 256.663
R1714 B.n650 B.n377 256.663
R1715 B.n656 B.n377 256.663
R1716 B.n658 B.n377 256.663
R1717 B.n664 B.n377 256.663
R1718 B.n666 B.n377 256.663
R1719 B.n672 B.n377 256.663
R1720 B.n674 B.n377 256.663
R1721 B.n680 B.n377 256.663
R1722 B.n682 B.n377 256.663
R1723 B.n688 B.n377 256.663
R1724 B.n690 B.n377 256.663
R1725 B.n697 B.n374 163.367
R1726 B.n701 B.n374 163.367
R1727 B.n701 B.n368 163.367
R1728 B.n709 B.n368 163.367
R1729 B.n709 B.n366 163.367
R1730 B.n713 B.n366 163.367
R1731 B.n713 B.n360 163.367
R1732 B.n721 B.n360 163.367
R1733 B.n721 B.n358 163.367
R1734 B.n725 B.n358 163.367
R1735 B.n725 B.n352 163.367
R1736 B.n735 B.n352 163.367
R1737 B.n735 B.n350 163.367
R1738 B.n739 B.n350 163.367
R1739 B.n739 B.n2 163.367
R1740 B.n801 B.n2 163.367
R1741 B.n801 B.n3 163.367
R1742 B.n797 B.n3 163.367
R1743 B.n797 B.n8 163.367
R1744 B.n793 B.n8 163.367
R1745 B.n793 B.n10 163.367
R1746 B.n789 B.n10 163.367
R1747 B.n789 B.n16 163.367
R1748 B.n785 B.n16 163.367
R1749 B.n785 B.n18 163.367
R1750 B.n781 B.n18 163.367
R1751 B.n781 B.n23 163.367
R1752 B.n777 B.n23 163.367
R1753 B.n777 B.n25 163.367
R1754 B.n773 B.n25 163.367
R1755 B.n773 B.n30 163.367
R1756 B.n769 B.n30 163.367
R1757 B.n446 B.n445 163.367
R1758 B.n448 B.n446 163.367
R1759 B.n452 B.n441 163.367
R1760 B.n456 B.n454 163.367
R1761 B.n460 B.n439 163.367
R1762 B.n464 B.n462 163.367
R1763 B.n468 B.n437 163.367
R1764 B.n472 B.n470 163.367
R1765 B.n476 B.n435 163.367
R1766 B.n480 B.n478 163.367
R1767 B.n484 B.n433 163.367
R1768 B.n488 B.n486 163.367
R1769 B.n492 B.n431 163.367
R1770 B.n496 B.n494 163.367
R1771 B.n500 B.n429 163.367
R1772 B.n504 B.n502 163.367
R1773 B.n508 B.n427 163.367
R1774 B.n512 B.n510 163.367
R1775 B.n516 B.n425 163.367
R1776 B.n520 B.n518 163.367
R1777 B.n524 B.n423 163.367
R1778 B.n528 B.n526 163.367
R1779 B.n532 B.n421 163.367
R1780 B.n536 B.n534 163.367
R1781 B.n540 B.n419 163.367
R1782 B.n544 B.n542 163.367
R1783 B.n548 B.n417 163.367
R1784 B.n552 B.n550 163.367
R1785 B.n559 B.n415 163.367
R1786 B.n563 B.n561 163.367
R1787 B.n567 B.n413 163.367
R1788 B.n571 B.n569 163.367
R1789 B.n575 B.n411 163.367
R1790 B.n579 B.n577 163.367
R1791 B.n583 B.n406 163.367
R1792 B.n587 B.n585 163.367
R1793 B.n591 B.n404 163.367
R1794 B.n595 B.n593 163.367
R1795 B.n599 B.n402 163.367
R1796 B.n603 B.n601 163.367
R1797 B.n607 B.n400 163.367
R1798 B.n611 B.n609 163.367
R1799 B.n615 B.n398 163.367
R1800 B.n619 B.n617 163.367
R1801 B.n623 B.n396 163.367
R1802 B.n627 B.n625 163.367
R1803 B.n631 B.n394 163.367
R1804 B.n635 B.n633 163.367
R1805 B.n639 B.n392 163.367
R1806 B.n643 B.n641 163.367
R1807 B.n647 B.n390 163.367
R1808 B.n651 B.n649 163.367
R1809 B.n655 B.n388 163.367
R1810 B.n659 B.n657 163.367
R1811 B.n663 B.n386 163.367
R1812 B.n667 B.n665 163.367
R1813 B.n671 B.n384 163.367
R1814 B.n675 B.n673 163.367
R1815 B.n679 B.n382 163.367
R1816 B.n683 B.n681 163.367
R1817 B.n687 B.n380 163.367
R1818 B.n691 B.n689 163.367
R1819 B.n695 B.n372 163.367
R1820 B.n703 B.n372 163.367
R1821 B.n703 B.n370 163.367
R1822 B.n707 B.n370 163.367
R1823 B.n707 B.n364 163.367
R1824 B.n715 B.n364 163.367
R1825 B.n715 B.n362 163.367
R1826 B.n719 B.n362 163.367
R1827 B.n719 B.n356 163.367
R1828 B.n727 B.n356 163.367
R1829 B.n727 B.n354 163.367
R1830 B.n732 B.n354 163.367
R1831 B.n732 B.n349 163.367
R1832 B.n741 B.n349 163.367
R1833 B.n742 B.n741 163.367
R1834 B.n742 B.n5 163.367
R1835 B.n6 B.n5 163.367
R1836 B.n7 B.n6 163.367
R1837 B.n747 B.n7 163.367
R1838 B.n747 B.n12 163.367
R1839 B.n13 B.n12 163.367
R1840 B.n14 B.n13 163.367
R1841 B.n752 B.n14 163.367
R1842 B.n752 B.n19 163.367
R1843 B.n20 B.n19 163.367
R1844 B.n21 B.n20 163.367
R1845 B.n757 B.n21 163.367
R1846 B.n757 B.n26 163.367
R1847 B.n27 B.n26 163.367
R1848 B.n28 B.n27 163.367
R1849 B.n762 B.n28 163.367
R1850 B.n762 B.n33 163.367
R1851 B.n104 B.n103 163.367
R1852 B.n108 B.n107 163.367
R1853 B.n112 B.n111 163.367
R1854 B.n116 B.n115 163.367
R1855 B.n120 B.n119 163.367
R1856 B.n124 B.n123 163.367
R1857 B.n128 B.n127 163.367
R1858 B.n132 B.n131 163.367
R1859 B.n136 B.n135 163.367
R1860 B.n140 B.n139 163.367
R1861 B.n144 B.n143 163.367
R1862 B.n148 B.n147 163.367
R1863 B.n152 B.n151 163.367
R1864 B.n156 B.n155 163.367
R1865 B.n160 B.n159 163.367
R1866 B.n164 B.n163 163.367
R1867 B.n168 B.n167 163.367
R1868 B.n172 B.n171 163.367
R1869 B.n176 B.n175 163.367
R1870 B.n180 B.n179 163.367
R1871 B.n184 B.n183 163.367
R1872 B.n188 B.n187 163.367
R1873 B.n192 B.n191 163.367
R1874 B.n196 B.n195 163.367
R1875 B.n200 B.n199 163.367
R1876 B.n204 B.n203 163.367
R1877 B.n208 B.n207 163.367
R1878 B.n212 B.n211 163.367
R1879 B.n216 B.n215 163.367
R1880 B.n220 B.n219 163.367
R1881 B.n224 B.n223 163.367
R1882 B.n228 B.n227 163.367
R1883 B.n232 B.n231 163.367
R1884 B.n237 B.n236 163.367
R1885 B.n241 B.n240 163.367
R1886 B.n245 B.n244 163.367
R1887 B.n249 B.n248 163.367
R1888 B.n253 B.n252 163.367
R1889 B.n257 B.n256 163.367
R1890 B.n261 B.n260 163.367
R1891 B.n265 B.n264 163.367
R1892 B.n269 B.n268 163.367
R1893 B.n273 B.n272 163.367
R1894 B.n277 B.n276 163.367
R1895 B.n281 B.n280 163.367
R1896 B.n285 B.n284 163.367
R1897 B.n289 B.n288 163.367
R1898 B.n293 B.n292 163.367
R1899 B.n297 B.n296 163.367
R1900 B.n301 B.n300 163.367
R1901 B.n305 B.n304 163.367
R1902 B.n309 B.n308 163.367
R1903 B.n313 B.n312 163.367
R1904 B.n317 B.n316 163.367
R1905 B.n321 B.n320 163.367
R1906 B.n325 B.n324 163.367
R1907 B.n329 B.n328 163.367
R1908 B.n333 B.n332 163.367
R1909 B.n337 B.n336 163.367
R1910 B.n341 B.n340 163.367
R1911 B.n345 B.n344 163.367
R1912 B.n766 B.n96 163.367
R1913 B.n444 B.n376 71.676
R1914 B.n448 B.n447 71.676
R1915 B.n453 B.n452 71.676
R1916 B.n456 B.n455 71.676
R1917 B.n461 B.n460 71.676
R1918 B.n464 B.n463 71.676
R1919 B.n469 B.n468 71.676
R1920 B.n472 B.n471 71.676
R1921 B.n477 B.n476 71.676
R1922 B.n480 B.n479 71.676
R1923 B.n485 B.n484 71.676
R1924 B.n488 B.n487 71.676
R1925 B.n493 B.n492 71.676
R1926 B.n496 B.n495 71.676
R1927 B.n501 B.n500 71.676
R1928 B.n504 B.n503 71.676
R1929 B.n509 B.n508 71.676
R1930 B.n512 B.n511 71.676
R1931 B.n517 B.n516 71.676
R1932 B.n520 B.n519 71.676
R1933 B.n525 B.n524 71.676
R1934 B.n528 B.n527 71.676
R1935 B.n533 B.n532 71.676
R1936 B.n536 B.n535 71.676
R1937 B.n541 B.n540 71.676
R1938 B.n544 B.n543 71.676
R1939 B.n549 B.n548 71.676
R1940 B.n552 B.n551 71.676
R1941 B.n560 B.n559 71.676
R1942 B.n563 B.n562 71.676
R1943 B.n568 B.n567 71.676
R1944 B.n571 B.n570 71.676
R1945 B.n576 B.n575 71.676
R1946 B.n579 B.n578 71.676
R1947 B.n584 B.n583 71.676
R1948 B.n587 B.n586 71.676
R1949 B.n592 B.n591 71.676
R1950 B.n595 B.n594 71.676
R1951 B.n600 B.n599 71.676
R1952 B.n603 B.n602 71.676
R1953 B.n608 B.n607 71.676
R1954 B.n611 B.n610 71.676
R1955 B.n616 B.n615 71.676
R1956 B.n619 B.n618 71.676
R1957 B.n624 B.n623 71.676
R1958 B.n627 B.n626 71.676
R1959 B.n632 B.n631 71.676
R1960 B.n635 B.n634 71.676
R1961 B.n640 B.n639 71.676
R1962 B.n643 B.n642 71.676
R1963 B.n648 B.n647 71.676
R1964 B.n651 B.n650 71.676
R1965 B.n656 B.n655 71.676
R1966 B.n659 B.n658 71.676
R1967 B.n664 B.n663 71.676
R1968 B.n667 B.n666 71.676
R1969 B.n672 B.n671 71.676
R1970 B.n675 B.n674 71.676
R1971 B.n680 B.n679 71.676
R1972 B.n683 B.n682 71.676
R1973 B.n688 B.n687 71.676
R1974 B.n691 B.n690 71.676
R1975 B.n34 B.n32 71.676
R1976 B.n104 B.n35 71.676
R1977 B.n108 B.n36 71.676
R1978 B.n112 B.n37 71.676
R1979 B.n116 B.n38 71.676
R1980 B.n120 B.n39 71.676
R1981 B.n124 B.n40 71.676
R1982 B.n128 B.n41 71.676
R1983 B.n132 B.n42 71.676
R1984 B.n136 B.n43 71.676
R1985 B.n140 B.n44 71.676
R1986 B.n144 B.n45 71.676
R1987 B.n148 B.n46 71.676
R1988 B.n152 B.n47 71.676
R1989 B.n156 B.n48 71.676
R1990 B.n160 B.n49 71.676
R1991 B.n164 B.n50 71.676
R1992 B.n168 B.n51 71.676
R1993 B.n172 B.n52 71.676
R1994 B.n176 B.n53 71.676
R1995 B.n180 B.n54 71.676
R1996 B.n184 B.n55 71.676
R1997 B.n188 B.n56 71.676
R1998 B.n192 B.n57 71.676
R1999 B.n196 B.n58 71.676
R2000 B.n200 B.n59 71.676
R2001 B.n204 B.n60 71.676
R2002 B.n208 B.n61 71.676
R2003 B.n212 B.n62 71.676
R2004 B.n216 B.n63 71.676
R2005 B.n220 B.n64 71.676
R2006 B.n224 B.n65 71.676
R2007 B.n228 B.n66 71.676
R2008 B.n232 B.n67 71.676
R2009 B.n237 B.n68 71.676
R2010 B.n241 B.n69 71.676
R2011 B.n245 B.n70 71.676
R2012 B.n249 B.n71 71.676
R2013 B.n253 B.n72 71.676
R2014 B.n257 B.n73 71.676
R2015 B.n261 B.n74 71.676
R2016 B.n265 B.n75 71.676
R2017 B.n269 B.n76 71.676
R2018 B.n273 B.n77 71.676
R2019 B.n277 B.n78 71.676
R2020 B.n281 B.n79 71.676
R2021 B.n285 B.n80 71.676
R2022 B.n289 B.n81 71.676
R2023 B.n293 B.n82 71.676
R2024 B.n297 B.n83 71.676
R2025 B.n301 B.n84 71.676
R2026 B.n305 B.n85 71.676
R2027 B.n309 B.n86 71.676
R2028 B.n313 B.n87 71.676
R2029 B.n317 B.n88 71.676
R2030 B.n321 B.n89 71.676
R2031 B.n325 B.n90 71.676
R2032 B.n329 B.n91 71.676
R2033 B.n333 B.n92 71.676
R2034 B.n337 B.n93 71.676
R2035 B.n341 B.n94 71.676
R2036 B.n345 B.n95 71.676
R2037 B.n96 B.n95 71.676
R2038 B.n344 B.n94 71.676
R2039 B.n340 B.n93 71.676
R2040 B.n336 B.n92 71.676
R2041 B.n332 B.n91 71.676
R2042 B.n328 B.n90 71.676
R2043 B.n324 B.n89 71.676
R2044 B.n320 B.n88 71.676
R2045 B.n316 B.n87 71.676
R2046 B.n312 B.n86 71.676
R2047 B.n308 B.n85 71.676
R2048 B.n304 B.n84 71.676
R2049 B.n300 B.n83 71.676
R2050 B.n296 B.n82 71.676
R2051 B.n292 B.n81 71.676
R2052 B.n288 B.n80 71.676
R2053 B.n284 B.n79 71.676
R2054 B.n280 B.n78 71.676
R2055 B.n276 B.n77 71.676
R2056 B.n272 B.n76 71.676
R2057 B.n268 B.n75 71.676
R2058 B.n264 B.n74 71.676
R2059 B.n260 B.n73 71.676
R2060 B.n256 B.n72 71.676
R2061 B.n252 B.n71 71.676
R2062 B.n248 B.n70 71.676
R2063 B.n244 B.n69 71.676
R2064 B.n240 B.n68 71.676
R2065 B.n236 B.n67 71.676
R2066 B.n231 B.n66 71.676
R2067 B.n227 B.n65 71.676
R2068 B.n223 B.n64 71.676
R2069 B.n219 B.n63 71.676
R2070 B.n215 B.n62 71.676
R2071 B.n211 B.n61 71.676
R2072 B.n207 B.n60 71.676
R2073 B.n203 B.n59 71.676
R2074 B.n199 B.n58 71.676
R2075 B.n195 B.n57 71.676
R2076 B.n191 B.n56 71.676
R2077 B.n187 B.n55 71.676
R2078 B.n183 B.n54 71.676
R2079 B.n179 B.n53 71.676
R2080 B.n175 B.n52 71.676
R2081 B.n171 B.n51 71.676
R2082 B.n167 B.n50 71.676
R2083 B.n163 B.n49 71.676
R2084 B.n159 B.n48 71.676
R2085 B.n155 B.n47 71.676
R2086 B.n151 B.n46 71.676
R2087 B.n147 B.n45 71.676
R2088 B.n143 B.n44 71.676
R2089 B.n139 B.n43 71.676
R2090 B.n135 B.n42 71.676
R2091 B.n131 B.n41 71.676
R2092 B.n127 B.n40 71.676
R2093 B.n123 B.n39 71.676
R2094 B.n119 B.n38 71.676
R2095 B.n115 B.n37 71.676
R2096 B.n111 B.n36 71.676
R2097 B.n107 B.n35 71.676
R2098 B.n103 B.n34 71.676
R2099 B.n445 B.n444 71.676
R2100 B.n447 B.n441 71.676
R2101 B.n454 B.n453 71.676
R2102 B.n455 B.n439 71.676
R2103 B.n462 B.n461 71.676
R2104 B.n463 B.n437 71.676
R2105 B.n470 B.n469 71.676
R2106 B.n471 B.n435 71.676
R2107 B.n478 B.n477 71.676
R2108 B.n479 B.n433 71.676
R2109 B.n486 B.n485 71.676
R2110 B.n487 B.n431 71.676
R2111 B.n494 B.n493 71.676
R2112 B.n495 B.n429 71.676
R2113 B.n502 B.n501 71.676
R2114 B.n503 B.n427 71.676
R2115 B.n510 B.n509 71.676
R2116 B.n511 B.n425 71.676
R2117 B.n518 B.n517 71.676
R2118 B.n519 B.n423 71.676
R2119 B.n526 B.n525 71.676
R2120 B.n527 B.n421 71.676
R2121 B.n534 B.n533 71.676
R2122 B.n535 B.n419 71.676
R2123 B.n542 B.n541 71.676
R2124 B.n543 B.n417 71.676
R2125 B.n550 B.n549 71.676
R2126 B.n551 B.n415 71.676
R2127 B.n561 B.n560 71.676
R2128 B.n562 B.n413 71.676
R2129 B.n569 B.n568 71.676
R2130 B.n570 B.n411 71.676
R2131 B.n577 B.n576 71.676
R2132 B.n578 B.n406 71.676
R2133 B.n585 B.n584 71.676
R2134 B.n586 B.n404 71.676
R2135 B.n593 B.n592 71.676
R2136 B.n594 B.n402 71.676
R2137 B.n601 B.n600 71.676
R2138 B.n602 B.n400 71.676
R2139 B.n609 B.n608 71.676
R2140 B.n610 B.n398 71.676
R2141 B.n617 B.n616 71.676
R2142 B.n618 B.n396 71.676
R2143 B.n625 B.n624 71.676
R2144 B.n626 B.n394 71.676
R2145 B.n633 B.n632 71.676
R2146 B.n634 B.n392 71.676
R2147 B.n641 B.n640 71.676
R2148 B.n642 B.n390 71.676
R2149 B.n649 B.n648 71.676
R2150 B.n650 B.n388 71.676
R2151 B.n657 B.n656 71.676
R2152 B.n658 B.n386 71.676
R2153 B.n665 B.n664 71.676
R2154 B.n666 B.n384 71.676
R2155 B.n673 B.n672 71.676
R2156 B.n674 B.n382 71.676
R2157 B.n681 B.n680 71.676
R2158 B.n682 B.n380 71.676
R2159 B.n689 B.n688 71.676
R2160 B.n690 B.n378 71.676
R2161 B.n409 B.n408 59.5399
R2162 B.n557 B.n556 59.5399
R2163 B.n101 B.n100 59.5399
R2164 B.n234 B.n98 59.5399
R2165 B.n696 B.n377 55.7642
R2166 B.n768 B.n767 55.7642
R2167 B.n696 B.n373 32.9738
R2168 B.n702 B.n373 32.9738
R2169 B.n702 B.n369 32.9738
R2170 B.n708 B.n369 32.9738
R2171 B.n714 B.n365 32.9738
R2172 B.n714 B.n361 32.9738
R2173 B.n720 B.n361 32.9738
R2174 B.n720 B.n357 32.9738
R2175 B.n726 B.n357 32.9738
R2176 B.n734 B.n353 32.9738
R2177 B.n734 B.n733 32.9738
R2178 B.n740 B.n4 32.9738
R2179 B.n800 B.n4 32.9738
R2180 B.n800 B.n799 32.9738
R2181 B.n799 B.n798 32.9738
R2182 B.n792 B.n11 32.9738
R2183 B.n792 B.n791 32.9738
R2184 B.n790 B.n15 32.9738
R2185 B.n784 B.n15 32.9738
R2186 B.n784 B.n783 32.9738
R2187 B.n783 B.n782 32.9738
R2188 B.n782 B.n22 32.9738
R2189 B.n776 B.n775 32.9738
R2190 B.n775 B.n774 32.9738
R2191 B.n774 B.n29 32.9738
R2192 B.n768 B.n29 32.9738
R2193 B.n740 B.t0 29.5795
R2194 B.n798 B.t1 29.5795
R2195 B.n770 B.n31 29.1907
R2196 B.n765 B.n764 29.1907
R2197 B.n694 B.n693 29.1907
R2198 B.n698 B.n375 29.1907
R2199 B.n708 B.t5 23.7607
R2200 B.n776 B.t9 23.7607
R2201 B B.n802 18.0485
R2202 B.n408 B.n407 17.0672
R2203 B.n556 B.n555 17.0672
R2204 B.n100 B.n99 17.0672
R2205 B.n98 B.n97 17.0672
R2206 B.n726 B.t3 16.9721
R2207 B.t2 B.n790 16.9721
R2208 B.t3 B.n353 16.0023
R2209 B.n791 B.t2 16.0023
R2210 B.n102 B.n31 10.6151
R2211 B.n105 B.n102 10.6151
R2212 B.n106 B.n105 10.6151
R2213 B.n109 B.n106 10.6151
R2214 B.n110 B.n109 10.6151
R2215 B.n113 B.n110 10.6151
R2216 B.n114 B.n113 10.6151
R2217 B.n117 B.n114 10.6151
R2218 B.n118 B.n117 10.6151
R2219 B.n121 B.n118 10.6151
R2220 B.n122 B.n121 10.6151
R2221 B.n125 B.n122 10.6151
R2222 B.n126 B.n125 10.6151
R2223 B.n129 B.n126 10.6151
R2224 B.n130 B.n129 10.6151
R2225 B.n133 B.n130 10.6151
R2226 B.n134 B.n133 10.6151
R2227 B.n137 B.n134 10.6151
R2228 B.n138 B.n137 10.6151
R2229 B.n141 B.n138 10.6151
R2230 B.n142 B.n141 10.6151
R2231 B.n145 B.n142 10.6151
R2232 B.n146 B.n145 10.6151
R2233 B.n149 B.n146 10.6151
R2234 B.n150 B.n149 10.6151
R2235 B.n153 B.n150 10.6151
R2236 B.n154 B.n153 10.6151
R2237 B.n157 B.n154 10.6151
R2238 B.n158 B.n157 10.6151
R2239 B.n161 B.n158 10.6151
R2240 B.n162 B.n161 10.6151
R2241 B.n165 B.n162 10.6151
R2242 B.n166 B.n165 10.6151
R2243 B.n169 B.n166 10.6151
R2244 B.n170 B.n169 10.6151
R2245 B.n173 B.n170 10.6151
R2246 B.n174 B.n173 10.6151
R2247 B.n177 B.n174 10.6151
R2248 B.n178 B.n177 10.6151
R2249 B.n181 B.n178 10.6151
R2250 B.n182 B.n181 10.6151
R2251 B.n185 B.n182 10.6151
R2252 B.n186 B.n185 10.6151
R2253 B.n189 B.n186 10.6151
R2254 B.n190 B.n189 10.6151
R2255 B.n193 B.n190 10.6151
R2256 B.n194 B.n193 10.6151
R2257 B.n197 B.n194 10.6151
R2258 B.n198 B.n197 10.6151
R2259 B.n201 B.n198 10.6151
R2260 B.n202 B.n201 10.6151
R2261 B.n205 B.n202 10.6151
R2262 B.n206 B.n205 10.6151
R2263 B.n209 B.n206 10.6151
R2264 B.n210 B.n209 10.6151
R2265 B.n213 B.n210 10.6151
R2266 B.n214 B.n213 10.6151
R2267 B.n218 B.n217 10.6151
R2268 B.n221 B.n218 10.6151
R2269 B.n222 B.n221 10.6151
R2270 B.n225 B.n222 10.6151
R2271 B.n226 B.n225 10.6151
R2272 B.n229 B.n226 10.6151
R2273 B.n230 B.n229 10.6151
R2274 B.n233 B.n230 10.6151
R2275 B.n238 B.n235 10.6151
R2276 B.n239 B.n238 10.6151
R2277 B.n242 B.n239 10.6151
R2278 B.n243 B.n242 10.6151
R2279 B.n246 B.n243 10.6151
R2280 B.n247 B.n246 10.6151
R2281 B.n250 B.n247 10.6151
R2282 B.n251 B.n250 10.6151
R2283 B.n254 B.n251 10.6151
R2284 B.n255 B.n254 10.6151
R2285 B.n258 B.n255 10.6151
R2286 B.n259 B.n258 10.6151
R2287 B.n262 B.n259 10.6151
R2288 B.n263 B.n262 10.6151
R2289 B.n266 B.n263 10.6151
R2290 B.n267 B.n266 10.6151
R2291 B.n270 B.n267 10.6151
R2292 B.n271 B.n270 10.6151
R2293 B.n274 B.n271 10.6151
R2294 B.n275 B.n274 10.6151
R2295 B.n278 B.n275 10.6151
R2296 B.n279 B.n278 10.6151
R2297 B.n282 B.n279 10.6151
R2298 B.n283 B.n282 10.6151
R2299 B.n286 B.n283 10.6151
R2300 B.n287 B.n286 10.6151
R2301 B.n290 B.n287 10.6151
R2302 B.n291 B.n290 10.6151
R2303 B.n294 B.n291 10.6151
R2304 B.n295 B.n294 10.6151
R2305 B.n298 B.n295 10.6151
R2306 B.n299 B.n298 10.6151
R2307 B.n302 B.n299 10.6151
R2308 B.n303 B.n302 10.6151
R2309 B.n306 B.n303 10.6151
R2310 B.n307 B.n306 10.6151
R2311 B.n310 B.n307 10.6151
R2312 B.n311 B.n310 10.6151
R2313 B.n314 B.n311 10.6151
R2314 B.n315 B.n314 10.6151
R2315 B.n318 B.n315 10.6151
R2316 B.n319 B.n318 10.6151
R2317 B.n322 B.n319 10.6151
R2318 B.n323 B.n322 10.6151
R2319 B.n326 B.n323 10.6151
R2320 B.n327 B.n326 10.6151
R2321 B.n330 B.n327 10.6151
R2322 B.n331 B.n330 10.6151
R2323 B.n334 B.n331 10.6151
R2324 B.n335 B.n334 10.6151
R2325 B.n338 B.n335 10.6151
R2326 B.n339 B.n338 10.6151
R2327 B.n342 B.n339 10.6151
R2328 B.n343 B.n342 10.6151
R2329 B.n346 B.n343 10.6151
R2330 B.n347 B.n346 10.6151
R2331 B.n765 B.n347 10.6151
R2332 B.n694 B.n371 10.6151
R2333 B.n704 B.n371 10.6151
R2334 B.n705 B.n704 10.6151
R2335 B.n706 B.n705 10.6151
R2336 B.n706 B.n363 10.6151
R2337 B.n716 B.n363 10.6151
R2338 B.n717 B.n716 10.6151
R2339 B.n718 B.n717 10.6151
R2340 B.n718 B.n355 10.6151
R2341 B.n728 B.n355 10.6151
R2342 B.n729 B.n728 10.6151
R2343 B.n731 B.n729 10.6151
R2344 B.n731 B.n730 10.6151
R2345 B.n730 B.n348 10.6151
R2346 B.n743 B.n348 10.6151
R2347 B.n744 B.n743 10.6151
R2348 B.n745 B.n744 10.6151
R2349 B.n746 B.n745 10.6151
R2350 B.n748 B.n746 10.6151
R2351 B.n749 B.n748 10.6151
R2352 B.n750 B.n749 10.6151
R2353 B.n751 B.n750 10.6151
R2354 B.n753 B.n751 10.6151
R2355 B.n754 B.n753 10.6151
R2356 B.n755 B.n754 10.6151
R2357 B.n756 B.n755 10.6151
R2358 B.n758 B.n756 10.6151
R2359 B.n759 B.n758 10.6151
R2360 B.n760 B.n759 10.6151
R2361 B.n761 B.n760 10.6151
R2362 B.n763 B.n761 10.6151
R2363 B.n764 B.n763 10.6151
R2364 B.n443 B.n375 10.6151
R2365 B.n443 B.n442 10.6151
R2366 B.n449 B.n442 10.6151
R2367 B.n450 B.n449 10.6151
R2368 B.n451 B.n450 10.6151
R2369 B.n451 B.n440 10.6151
R2370 B.n457 B.n440 10.6151
R2371 B.n458 B.n457 10.6151
R2372 B.n459 B.n458 10.6151
R2373 B.n459 B.n438 10.6151
R2374 B.n465 B.n438 10.6151
R2375 B.n466 B.n465 10.6151
R2376 B.n467 B.n466 10.6151
R2377 B.n467 B.n436 10.6151
R2378 B.n473 B.n436 10.6151
R2379 B.n474 B.n473 10.6151
R2380 B.n475 B.n474 10.6151
R2381 B.n475 B.n434 10.6151
R2382 B.n481 B.n434 10.6151
R2383 B.n482 B.n481 10.6151
R2384 B.n483 B.n482 10.6151
R2385 B.n483 B.n432 10.6151
R2386 B.n489 B.n432 10.6151
R2387 B.n490 B.n489 10.6151
R2388 B.n491 B.n490 10.6151
R2389 B.n491 B.n430 10.6151
R2390 B.n497 B.n430 10.6151
R2391 B.n498 B.n497 10.6151
R2392 B.n499 B.n498 10.6151
R2393 B.n499 B.n428 10.6151
R2394 B.n505 B.n428 10.6151
R2395 B.n506 B.n505 10.6151
R2396 B.n507 B.n506 10.6151
R2397 B.n507 B.n426 10.6151
R2398 B.n513 B.n426 10.6151
R2399 B.n514 B.n513 10.6151
R2400 B.n515 B.n514 10.6151
R2401 B.n515 B.n424 10.6151
R2402 B.n521 B.n424 10.6151
R2403 B.n522 B.n521 10.6151
R2404 B.n523 B.n522 10.6151
R2405 B.n523 B.n422 10.6151
R2406 B.n529 B.n422 10.6151
R2407 B.n530 B.n529 10.6151
R2408 B.n531 B.n530 10.6151
R2409 B.n531 B.n420 10.6151
R2410 B.n537 B.n420 10.6151
R2411 B.n538 B.n537 10.6151
R2412 B.n539 B.n538 10.6151
R2413 B.n539 B.n418 10.6151
R2414 B.n545 B.n418 10.6151
R2415 B.n546 B.n545 10.6151
R2416 B.n547 B.n546 10.6151
R2417 B.n547 B.n416 10.6151
R2418 B.n553 B.n416 10.6151
R2419 B.n554 B.n553 10.6151
R2420 B.n558 B.n554 10.6151
R2421 B.n564 B.n414 10.6151
R2422 B.n565 B.n564 10.6151
R2423 B.n566 B.n565 10.6151
R2424 B.n566 B.n412 10.6151
R2425 B.n572 B.n412 10.6151
R2426 B.n573 B.n572 10.6151
R2427 B.n574 B.n573 10.6151
R2428 B.n574 B.n410 10.6151
R2429 B.n581 B.n580 10.6151
R2430 B.n582 B.n581 10.6151
R2431 B.n582 B.n405 10.6151
R2432 B.n588 B.n405 10.6151
R2433 B.n589 B.n588 10.6151
R2434 B.n590 B.n589 10.6151
R2435 B.n590 B.n403 10.6151
R2436 B.n596 B.n403 10.6151
R2437 B.n597 B.n596 10.6151
R2438 B.n598 B.n597 10.6151
R2439 B.n598 B.n401 10.6151
R2440 B.n604 B.n401 10.6151
R2441 B.n605 B.n604 10.6151
R2442 B.n606 B.n605 10.6151
R2443 B.n606 B.n399 10.6151
R2444 B.n612 B.n399 10.6151
R2445 B.n613 B.n612 10.6151
R2446 B.n614 B.n613 10.6151
R2447 B.n614 B.n397 10.6151
R2448 B.n620 B.n397 10.6151
R2449 B.n621 B.n620 10.6151
R2450 B.n622 B.n621 10.6151
R2451 B.n622 B.n395 10.6151
R2452 B.n628 B.n395 10.6151
R2453 B.n629 B.n628 10.6151
R2454 B.n630 B.n629 10.6151
R2455 B.n630 B.n393 10.6151
R2456 B.n636 B.n393 10.6151
R2457 B.n637 B.n636 10.6151
R2458 B.n638 B.n637 10.6151
R2459 B.n638 B.n391 10.6151
R2460 B.n644 B.n391 10.6151
R2461 B.n645 B.n644 10.6151
R2462 B.n646 B.n645 10.6151
R2463 B.n646 B.n389 10.6151
R2464 B.n652 B.n389 10.6151
R2465 B.n653 B.n652 10.6151
R2466 B.n654 B.n653 10.6151
R2467 B.n654 B.n387 10.6151
R2468 B.n660 B.n387 10.6151
R2469 B.n661 B.n660 10.6151
R2470 B.n662 B.n661 10.6151
R2471 B.n662 B.n385 10.6151
R2472 B.n668 B.n385 10.6151
R2473 B.n669 B.n668 10.6151
R2474 B.n670 B.n669 10.6151
R2475 B.n670 B.n383 10.6151
R2476 B.n676 B.n383 10.6151
R2477 B.n677 B.n676 10.6151
R2478 B.n678 B.n677 10.6151
R2479 B.n678 B.n381 10.6151
R2480 B.n684 B.n381 10.6151
R2481 B.n685 B.n684 10.6151
R2482 B.n686 B.n685 10.6151
R2483 B.n686 B.n379 10.6151
R2484 B.n692 B.n379 10.6151
R2485 B.n693 B.n692 10.6151
R2486 B.n699 B.n698 10.6151
R2487 B.n700 B.n699 10.6151
R2488 B.n700 B.n367 10.6151
R2489 B.n710 B.n367 10.6151
R2490 B.n711 B.n710 10.6151
R2491 B.n712 B.n711 10.6151
R2492 B.n712 B.n359 10.6151
R2493 B.n722 B.n359 10.6151
R2494 B.n723 B.n722 10.6151
R2495 B.n724 B.n723 10.6151
R2496 B.n724 B.n351 10.6151
R2497 B.n736 B.n351 10.6151
R2498 B.n737 B.n736 10.6151
R2499 B.n738 B.n737 10.6151
R2500 B.n738 B.n0 10.6151
R2501 B.n796 B.n1 10.6151
R2502 B.n796 B.n795 10.6151
R2503 B.n795 B.n794 10.6151
R2504 B.n794 B.n9 10.6151
R2505 B.n788 B.n9 10.6151
R2506 B.n788 B.n787 10.6151
R2507 B.n787 B.n786 10.6151
R2508 B.n786 B.n17 10.6151
R2509 B.n780 B.n17 10.6151
R2510 B.n780 B.n779 10.6151
R2511 B.n779 B.n778 10.6151
R2512 B.n778 B.n24 10.6151
R2513 B.n772 B.n24 10.6151
R2514 B.n772 B.n771 10.6151
R2515 B.n771 B.n770 10.6151
R2516 B.t5 B.n365 9.21364
R2517 B.t9 B.n22 9.21364
R2518 B.n217 B.n101 6.5566
R2519 B.n234 B.n233 6.5566
R2520 B.n557 B.n414 6.5566
R2521 B.n410 B.n409 6.5566
R2522 B.n214 B.n101 4.05904
R2523 B.n235 B.n234 4.05904
R2524 B.n558 B.n557 4.05904
R2525 B.n580 B.n409 4.05904
R2526 B.n733 B.t0 3.39481
R2527 B.n11 B.t1 3.39481
R2528 B.n802 B.n0 2.81026
R2529 B.n802 B.n1 2.81026
R2530 VN.n0 VN.t2 855.718
R2531 VN.n1 VN.t1 855.718
R2532 VN.n0 VN.t0 855.693
R2533 VN.n1 VN.t3 855.693
R2534 VN VN.n1 114.724
R2535 VN VN.n0 70.265
R2536 VDD2.n2 VDD2.n0 99.5479
R2537 VDD2.n2 VDD2.n1 58.5486
R2538 VDD2.n1 VDD2.t0 1.13778
R2539 VDD2.n1 VDD2.t2 1.13778
R2540 VDD2.n0 VDD2.t1 1.13778
R2541 VDD2.n0 VDD2.t3 1.13778
R2542 VDD2 VDD2.n2 0.0586897
C0 VDD2 VP 0.263965f
C1 VN VDD1 0.147252f
C2 VN VTAIL 3.3083f
C3 VN VP 5.7144f
C4 VTAIL VDD1 10.1483f
C5 VDD1 VP 4.08131f
C6 VTAIL VP 3.3224f
C7 VN VDD2 3.96482f
C8 VDD1 VDD2 0.534602f
C9 VTAIL VDD2 10.1888f
C10 VDD2 B 3.043485f
C11 VDD1 B 7.47869f
C12 VTAIL B 11.715693f
C13 VN B 9.06813f
C14 VP B 4.94191f
C15 VDD2.t1 B 0.406548f
C16 VDD2.t3 B 0.406548f
C17 VDD2.n0 B 4.55825f
C18 VDD2.t0 B 0.406548f
C19 VDD2.t2 B 0.406548f
C20 VDD2.n1 B 3.69493f
C21 VDD2.n2 B 4.24203f
C22 VN.t2 B 1.45871f
C23 VN.t0 B 1.45869f
C24 VN.n0 B 1.07485f
C25 VN.t1 B 1.45871f
C26 VN.t3 B 1.45869f
C27 VN.n1 B 2.03834f
C28 VDD1.t0 B 0.403447f
C29 VDD1.t3 B 0.403447f
C30 VDD1.n0 B 3.66708f
C31 VDD1.t2 B 0.403447f
C32 VDD1.t1 B 0.403447f
C33 VDD1.n1 B 4.55432f
C34 VTAIL.n0 B 0.021394f
C35 VTAIL.n1 B 0.016402f
C36 VTAIL.n2 B 0.008813f
C37 VTAIL.n3 B 0.020832f
C38 VTAIL.n4 B 0.009332f
C39 VTAIL.n5 B 0.016402f
C40 VTAIL.n6 B 0.008813f
C41 VTAIL.n7 B 0.020832f
C42 VTAIL.n8 B 0.009073f
C43 VTAIL.n9 B 0.016402f
C44 VTAIL.n10 B 0.009332f
C45 VTAIL.n11 B 0.020832f
C46 VTAIL.n12 B 0.009332f
C47 VTAIL.n13 B 0.016402f
C48 VTAIL.n14 B 0.008813f
C49 VTAIL.n15 B 0.020832f
C50 VTAIL.n16 B 0.009332f
C51 VTAIL.n17 B 0.016402f
C52 VTAIL.n18 B 0.008813f
C53 VTAIL.n19 B 0.020832f
C54 VTAIL.n20 B 0.009332f
C55 VTAIL.n21 B 0.016402f
C56 VTAIL.n22 B 0.008813f
C57 VTAIL.n23 B 0.020832f
C58 VTAIL.n24 B 0.009332f
C59 VTAIL.n25 B 0.016402f
C60 VTAIL.n26 B 0.008813f
C61 VTAIL.n27 B 0.020832f
C62 VTAIL.n28 B 0.009332f
C63 VTAIL.n29 B 1.24826f
C64 VTAIL.n30 B 0.008813f
C65 VTAIL.t1 B 0.034485f
C66 VTAIL.n31 B 0.116885f
C67 VTAIL.n32 B 0.012306f
C68 VTAIL.n33 B 0.015624f
C69 VTAIL.n34 B 0.020832f
C70 VTAIL.n35 B 0.009332f
C71 VTAIL.n36 B 0.008813f
C72 VTAIL.n37 B 0.016402f
C73 VTAIL.n38 B 0.016402f
C74 VTAIL.n39 B 0.008813f
C75 VTAIL.n40 B 0.009332f
C76 VTAIL.n41 B 0.020832f
C77 VTAIL.n42 B 0.020832f
C78 VTAIL.n43 B 0.009332f
C79 VTAIL.n44 B 0.008813f
C80 VTAIL.n45 B 0.016402f
C81 VTAIL.n46 B 0.016402f
C82 VTAIL.n47 B 0.008813f
C83 VTAIL.n48 B 0.009332f
C84 VTAIL.n49 B 0.020832f
C85 VTAIL.n50 B 0.020832f
C86 VTAIL.n51 B 0.009332f
C87 VTAIL.n52 B 0.008813f
C88 VTAIL.n53 B 0.016402f
C89 VTAIL.n54 B 0.016402f
C90 VTAIL.n55 B 0.008813f
C91 VTAIL.n56 B 0.009332f
C92 VTAIL.n57 B 0.020832f
C93 VTAIL.n58 B 0.020832f
C94 VTAIL.n59 B 0.009332f
C95 VTAIL.n60 B 0.008813f
C96 VTAIL.n61 B 0.016402f
C97 VTAIL.n62 B 0.016402f
C98 VTAIL.n63 B 0.008813f
C99 VTAIL.n64 B 0.009332f
C100 VTAIL.n65 B 0.020832f
C101 VTAIL.n66 B 0.020832f
C102 VTAIL.n67 B 0.009332f
C103 VTAIL.n68 B 0.008813f
C104 VTAIL.n69 B 0.016402f
C105 VTAIL.n70 B 0.016402f
C106 VTAIL.n71 B 0.008813f
C107 VTAIL.n72 B 0.008813f
C108 VTAIL.n73 B 0.009332f
C109 VTAIL.n74 B 0.020832f
C110 VTAIL.n75 B 0.020832f
C111 VTAIL.n76 B 0.020832f
C112 VTAIL.n77 B 0.009073f
C113 VTAIL.n78 B 0.008813f
C114 VTAIL.n79 B 0.016402f
C115 VTAIL.n80 B 0.016402f
C116 VTAIL.n81 B 0.008813f
C117 VTAIL.n82 B 0.009332f
C118 VTAIL.n83 B 0.020832f
C119 VTAIL.n84 B 0.020832f
C120 VTAIL.n85 B 0.009332f
C121 VTAIL.n86 B 0.008813f
C122 VTAIL.n87 B 0.016402f
C123 VTAIL.n88 B 0.016402f
C124 VTAIL.n89 B 0.008813f
C125 VTAIL.n90 B 0.009332f
C126 VTAIL.n91 B 0.020832f
C127 VTAIL.n92 B 0.042162f
C128 VTAIL.n93 B 0.009332f
C129 VTAIL.n94 B 0.008813f
C130 VTAIL.n95 B 0.035447f
C131 VTAIL.n96 B 0.023211f
C132 VTAIL.n97 B 0.060571f
C133 VTAIL.n98 B 0.021394f
C134 VTAIL.n99 B 0.016402f
C135 VTAIL.n100 B 0.008813f
C136 VTAIL.n101 B 0.020832f
C137 VTAIL.n102 B 0.009332f
C138 VTAIL.n103 B 0.016402f
C139 VTAIL.n104 B 0.008813f
C140 VTAIL.n105 B 0.020832f
C141 VTAIL.n106 B 0.009073f
C142 VTAIL.n107 B 0.016402f
C143 VTAIL.n108 B 0.009332f
C144 VTAIL.n109 B 0.020832f
C145 VTAIL.n110 B 0.009332f
C146 VTAIL.n111 B 0.016402f
C147 VTAIL.n112 B 0.008813f
C148 VTAIL.n113 B 0.020832f
C149 VTAIL.n114 B 0.009332f
C150 VTAIL.n115 B 0.016402f
C151 VTAIL.n116 B 0.008813f
C152 VTAIL.n117 B 0.020832f
C153 VTAIL.n118 B 0.009332f
C154 VTAIL.n119 B 0.016402f
C155 VTAIL.n120 B 0.008813f
C156 VTAIL.n121 B 0.020832f
C157 VTAIL.n122 B 0.009332f
C158 VTAIL.n123 B 0.016402f
C159 VTAIL.n124 B 0.008813f
C160 VTAIL.n125 B 0.020832f
C161 VTAIL.n126 B 0.009332f
C162 VTAIL.n127 B 1.24826f
C163 VTAIL.n128 B 0.008813f
C164 VTAIL.t3 B 0.034485f
C165 VTAIL.n129 B 0.116885f
C166 VTAIL.n130 B 0.012306f
C167 VTAIL.n131 B 0.015624f
C168 VTAIL.n132 B 0.020832f
C169 VTAIL.n133 B 0.009332f
C170 VTAIL.n134 B 0.008813f
C171 VTAIL.n135 B 0.016402f
C172 VTAIL.n136 B 0.016402f
C173 VTAIL.n137 B 0.008813f
C174 VTAIL.n138 B 0.009332f
C175 VTAIL.n139 B 0.020832f
C176 VTAIL.n140 B 0.020832f
C177 VTAIL.n141 B 0.009332f
C178 VTAIL.n142 B 0.008813f
C179 VTAIL.n143 B 0.016402f
C180 VTAIL.n144 B 0.016402f
C181 VTAIL.n145 B 0.008813f
C182 VTAIL.n146 B 0.009332f
C183 VTAIL.n147 B 0.020832f
C184 VTAIL.n148 B 0.020832f
C185 VTAIL.n149 B 0.009332f
C186 VTAIL.n150 B 0.008813f
C187 VTAIL.n151 B 0.016402f
C188 VTAIL.n152 B 0.016402f
C189 VTAIL.n153 B 0.008813f
C190 VTAIL.n154 B 0.009332f
C191 VTAIL.n155 B 0.020832f
C192 VTAIL.n156 B 0.020832f
C193 VTAIL.n157 B 0.009332f
C194 VTAIL.n158 B 0.008813f
C195 VTAIL.n159 B 0.016402f
C196 VTAIL.n160 B 0.016402f
C197 VTAIL.n161 B 0.008813f
C198 VTAIL.n162 B 0.009332f
C199 VTAIL.n163 B 0.020832f
C200 VTAIL.n164 B 0.020832f
C201 VTAIL.n165 B 0.009332f
C202 VTAIL.n166 B 0.008813f
C203 VTAIL.n167 B 0.016402f
C204 VTAIL.n168 B 0.016402f
C205 VTAIL.n169 B 0.008813f
C206 VTAIL.n170 B 0.008813f
C207 VTAIL.n171 B 0.009332f
C208 VTAIL.n172 B 0.020832f
C209 VTAIL.n173 B 0.020832f
C210 VTAIL.n174 B 0.020832f
C211 VTAIL.n175 B 0.009073f
C212 VTAIL.n176 B 0.008813f
C213 VTAIL.n177 B 0.016402f
C214 VTAIL.n178 B 0.016402f
C215 VTAIL.n179 B 0.008813f
C216 VTAIL.n180 B 0.009332f
C217 VTAIL.n181 B 0.020832f
C218 VTAIL.n182 B 0.020832f
C219 VTAIL.n183 B 0.009332f
C220 VTAIL.n184 B 0.008813f
C221 VTAIL.n185 B 0.016402f
C222 VTAIL.n186 B 0.016402f
C223 VTAIL.n187 B 0.008813f
C224 VTAIL.n188 B 0.009332f
C225 VTAIL.n189 B 0.020832f
C226 VTAIL.n190 B 0.042162f
C227 VTAIL.n191 B 0.009332f
C228 VTAIL.n192 B 0.008813f
C229 VTAIL.n193 B 0.035447f
C230 VTAIL.n194 B 0.023211f
C231 VTAIL.n195 B 0.077542f
C232 VTAIL.n196 B 0.021394f
C233 VTAIL.n197 B 0.016402f
C234 VTAIL.n198 B 0.008813f
C235 VTAIL.n199 B 0.020832f
C236 VTAIL.n200 B 0.009332f
C237 VTAIL.n201 B 0.016402f
C238 VTAIL.n202 B 0.008813f
C239 VTAIL.n203 B 0.020832f
C240 VTAIL.n204 B 0.009073f
C241 VTAIL.n205 B 0.016402f
C242 VTAIL.n206 B 0.009332f
C243 VTAIL.n207 B 0.020832f
C244 VTAIL.n208 B 0.009332f
C245 VTAIL.n209 B 0.016402f
C246 VTAIL.n210 B 0.008813f
C247 VTAIL.n211 B 0.020832f
C248 VTAIL.n212 B 0.009332f
C249 VTAIL.n213 B 0.016402f
C250 VTAIL.n214 B 0.008813f
C251 VTAIL.n215 B 0.020832f
C252 VTAIL.n216 B 0.009332f
C253 VTAIL.n217 B 0.016402f
C254 VTAIL.n218 B 0.008813f
C255 VTAIL.n219 B 0.020832f
C256 VTAIL.n220 B 0.009332f
C257 VTAIL.n221 B 0.016402f
C258 VTAIL.n222 B 0.008813f
C259 VTAIL.n223 B 0.020832f
C260 VTAIL.n224 B 0.009332f
C261 VTAIL.n225 B 1.24826f
C262 VTAIL.n226 B 0.008813f
C263 VTAIL.t6 B 0.034485f
C264 VTAIL.n227 B 0.116885f
C265 VTAIL.n228 B 0.012306f
C266 VTAIL.n229 B 0.015624f
C267 VTAIL.n230 B 0.020832f
C268 VTAIL.n231 B 0.009332f
C269 VTAIL.n232 B 0.008813f
C270 VTAIL.n233 B 0.016402f
C271 VTAIL.n234 B 0.016402f
C272 VTAIL.n235 B 0.008813f
C273 VTAIL.n236 B 0.009332f
C274 VTAIL.n237 B 0.020832f
C275 VTAIL.n238 B 0.020832f
C276 VTAIL.n239 B 0.009332f
C277 VTAIL.n240 B 0.008813f
C278 VTAIL.n241 B 0.016402f
C279 VTAIL.n242 B 0.016402f
C280 VTAIL.n243 B 0.008813f
C281 VTAIL.n244 B 0.009332f
C282 VTAIL.n245 B 0.020832f
C283 VTAIL.n246 B 0.020832f
C284 VTAIL.n247 B 0.009332f
C285 VTAIL.n248 B 0.008813f
C286 VTAIL.n249 B 0.016402f
C287 VTAIL.n250 B 0.016402f
C288 VTAIL.n251 B 0.008813f
C289 VTAIL.n252 B 0.009332f
C290 VTAIL.n253 B 0.020832f
C291 VTAIL.n254 B 0.020832f
C292 VTAIL.n255 B 0.009332f
C293 VTAIL.n256 B 0.008813f
C294 VTAIL.n257 B 0.016402f
C295 VTAIL.n258 B 0.016402f
C296 VTAIL.n259 B 0.008813f
C297 VTAIL.n260 B 0.009332f
C298 VTAIL.n261 B 0.020832f
C299 VTAIL.n262 B 0.020832f
C300 VTAIL.n263 B 0.009332f
C301 VTAIL.n264 B 0.008813f
C302 VTAIL.n265 B 0.016402f
C303 VTAIL.n266 B 0.016402f
C304 VTAIL.n267 B 0.008813f
C305 VTAIL.n268 B 0.008813f
C306 VTAIL.n269 B 0.009332f
C307 VTAIL.n270 B 0.020832f
C308 VTAIL.n271 B 0.020832f
C309 VTAIL.n272 B 0.020832f
C310 VTAIL.n273 B 0.009073f
C311 VTAIL.n274 B 0.008813f
C312 VTAIL.n275 B 0.016402f
C313 VTAIL.n276 B 0.016402f
C314 VTAIL.n277 B 0.008813f
C315 VTAIL.n278 B 0.009332f
C316 VTAIL.n279 B 0.020832f
C317 VTAIL.n280 B 0.020832f
C318 VTAIL.n281 B 0.009332f
C319 VTAIL.n282 B 0.008813f
C320 VTAIL.n283 B 0.016402f
C321 VTAIL.n284 B 0.016402f
C322 VTAIL.n285 B 0.008813f
C323 VTAIL.n286 B 0.009332f
C324 VTAIL.n287 B 0.020832f
C325 VTAIL.n288 B 0.042162f
C326 VTAIL.n289 B 0.009332f
C327 VTAIL.n290 B 0.008813f
C328 VTAIL.n291 B 0.035447f
C329 VTAIL.n292 B 0.023211f
C330 VTAIL.n293 B 1.1088f
C331 VTAIL.n294 B 0.021394f
C332 VTAIL.n295 B 0.016402f
C333 VTAIL.n296 B 0.008813f
C334 VTAIL.n297 B 0.020832f
C335 VTAIL.n298 B 0.009332f
C336 VTAIL.n299 B 0.016402f
C337 VTAIL.n300 B 0.008813f
C338 VTAIL.n301 B 0.020832f
C339 VTAIL.n302 B 0.009073f
C340 VTAIL.n303 B 0.016402f
C341 VTAIL.n304 B 0.009073f
C342 VTAIL.n305 B 0.008813f
C343 VTAIL.n306 B 0.020832f
C344 VTAIL.n307 B 0.020832f
C345 VTAIL.n308 B 0.009332f
C346 VTAIL.n309 B 0.016402f
C347 VTAIL.n310 B 0.008813f
C348 VTAIL.n311 B 0.020832f
C349 VTAIL.n312 B 0.009332f
C350 VTAIL.n313 B 0.016402f
C351 VTAIL.n314 B 0.008813f
C352 VTAIL.n315 B 0.020832f
C353 VTAIL.n316 B 0.009332f
C354 VTAIL.n317 B 0.016402f
C355 VTAIL.n318 B 0.008813f
C356 VTAIL.n319 B 0.020832f
C357 VTAIL.n320 B 0.009332f
C358 VTAIL.n321 B 0.016402f
C359 VTAIL.n322 B 0.008813f
C360 VTAIL.n323 B 0.020832f
C361 VTAIL.n324 B 0.009332f
C362 VTAIL.n325 B 1.24826f
C363 VTAIL.n326 B 0.008813f
C364 VTAIL.t7 B 0.034485f
C365 VTAIL.n327 B 0.116885f
C366 VTAIL.n328 B 0.012306f
C367 VTAIL.n329 B 0.015624f
C368 VTAIL.n330 B 0.020832f
C369 VTAIL.n331 B 0.009332f
C370 VTAIL.n332 B 0.008813f
C371 VTAIL.n333 B 0.016402f
C372 VTAIL.n334 B 0.016402f
C373 VTAIL.n335 B 0.008813f
C374 VTAIL.n336 B 0.009332f
C375 VTAIL.n337 B 0.020832f
C376 VTAIL.n338 B 0.020832f
C377 VTAIL.n339 B 0.009332f
C378 VTAIL.n340 B 0.008813f
C379 VTAIL.n341 B 0.016402f
C380 VTAIL.n342 B 0.016402f
C381 VTAIL.n343 B 0.008813f
C382 VTAIL.n344 B 0.009332f
C383 VTAIL.n345 B 0.020832f
C384 VTAIL.n346 B 0.020832f
C385 VTAIL.n347 B 0.009332f
C386 VTAIL.n348 B 0.008813f
C387 VTAIL.n349 B 0.016402f
C388 VTAIL.n350 B 0.016402f
C389 VTAIL.n351 B 0.008813f
C390 VTAIL.n352 B 0.009332f
C391 VTAIL.n353 B 0.020832f
C392 VTAIL.n354 B 0.020832f
C393 VTAIL.n355 B 0.009332f
C394 VTAIL.n356 B 0.008813f
C395 VTAIL.n357 B 0.016402f
C396 VTAIL.n358 B 0.016402f
C397 VTAIL.n359 B 0.008813f
C398 VTAIL.n360 B 0.009332f
C399 VTAIL.n361 B 0.020832f
C400 VTAIL.n362 B 0.020832f
C401 VTAIL.n363 B 0.009332f
C402 VTAIL.n364 B 0.008813f
C403 VTAIL.n365 B 0.016402f
C404 VTAIL.n366 B 0.016402f
C405 VTAIL.n367 B 0.008813f
C406 VTAIL.n368 B 0.009332f
C407 VTAIL.n369 B 0.020832f
C408 VTAIL.n370 B 0.020832f
C409 VTAIL.n371 B 0.009332f
C410 VTAIL.n372 B 0.008813f
C411 VTAIL.n373 B 0.016402f
C412 VTAIL.n374 B 0.016402f
C413 VTAIL.n375 B 0.008813f
C414 VTAIL.n376 B 0.009332f
C415 VTAIL.n377 B 0.020832f
C416 VTAIL.n378 B 0.020832f
C417 VTAIL.n379 B 0.009332f
C418 VTAIL.n380 B 0.008813f
C419 VTAIL.n381 B 0.016402f
C420 VTAIL.n382 B 0.016402f
C421 VTAIL.n383 B 0.008813f
C422 VTAIL.n384 B 0.009332f
C423 VTAIL.n385 B 0.020832f
C424 VTAIL.n386 B 0.042162f
C425 VTAIL.n387 B 0.009332f
C426 VTAIL.n388 B 0.008813f
C427 VTAIL.n389 B 0.035447f
C428 VTAIL.n390 B 0.023211f
C429 VTAIL.n391 B 1.1088f
C430 VTAIL.n392 B 0.021394f
C431 VTAIL.n393 B 0.016402f
C432 VTAIL.n394 B 0.008813f
C433 VTAIL.n395 B 0.020832f
C434 VTAIL.n396 B 0.009332f
C435 VTAIL.n397 B 0.016402f
C436 VTAIL.n398 B 0.008813f
C437 VTAIL.n399 B 0.020832f
C438 VTAIL.n400 B 0.009073f
C439 VTAIL.n401 B 0.016402f
C440 VTAIL.n402 B 0.009073f
C441 VTAIL.n403 B 0.008813f
C442 VTAIL.n404 B 0.020832f
C443 VTAIL.n405 B 0.020832f
C444 VTAIL.n406 B 0.009332f
C445 VTAIL.n407 B 0.016402f
C446 VTAIL.n408 B 0.008813f
C447 VTAIL.n409 B 0.020832f
C448 VTAIL.n410 B 0.009332f
C449 VTAIL.n411 B 0.016402f
C450 VTAIL.n412 B 0.008813f
C451 VTAIL.n413 B 0.020832f
C452 VTAIL.n414 B 0.009332f
C453 VTAIL.n415 B 0.016402f
C454 VTAIL.n416 B 0.008813f
C455 VTAIL.n417 B 0.020832f
C456 VTAIL.n418 B 0.009332f
C457 VTAIL.n419 B 0.016402f
C458 VTAIL.n420 B 0.008813f
C459 VTAIL.n421 B 0.020832f
C460 VTAIL.n422 B 0.009332f
C461 VTAIL.n423 B 1.24826f
C462 VTAIL.n424 B 0.008813f
C463 VTAIL.t0 B 0.034485f
C464 VTAIL.n425 B 0.116885f
C465 VTAIL.n426 B 0.012306f
C466 VTAIL.n427 B 0.015624f
C467 VTAIL.n428 B 0.020832f
C468 VTAIL.n429 B 0.009332f
C469 VTAIL.n430 B 0.008813f
C470 VTAIL.n431 B 0.016402f
C471 VTAIL.n432 B 0.016402f
C472 VTAIL.n433 B 0.008813f
C473 VTAIL.n434 B 0.009332f
C474 VTAIL.n435 B 0.020832f
C475 VTAIL.n436 B 0.020832f
C476 VTAIL.n437 B 0.009332f
C477 VTAIL.n438 B 0.008813f
C478 VTAIL.n439 B 0.016402f
C479 VTAIL.n440 B 0.016402f
C480 VTAIL.n441 B 0.008813f
C481 VTAIL.n442 B 0.009332f
C482 VTAIL.n443 B 0.020832f
C483 VTAIL.n444 B 0.020832f
C484 VTAIL.n445 B 0.009332f
C485 VTAIL.n446 B 0.008813f
C486 VTAIL.n447 B 0.016402f
C487 VTAIL.n448 B 0.016402f
C488 VTAIL.n449 B 0.008813f
C489 VTAIL.n450 B 0.009332f
C490 VTAIL.n451 B 0.020832f
C491 VTAIL.n452 B 0.020832f
C492 VTAIL.n453 B 0.009332f
C493 VTAIL.n454 B 0.008813f
C494 VTAIL.n455 B 0.016402f
C495 VTAIL.n456 B 0.016402f
C496 VTAIL.n457 B 0.008813f
C497 VTAIL.n458 B 0.009332f
C498 VTAIL.n459 B 0.020832f
C499 VTAIL.n460 B 0.020832f
C500 VTAIL.n461 B 0.009332f
C501 VTAIL.n462 B 0.008813f
C502 VTAIL.n463 B 0.016402f
C503 VTAIL.n464 B 0.016402f
C504 VTAIL.n465 B 0.008813f
C505 VTAIL.n466 B 0.009332f
C506 VTAIL.n467 B 0.020832f
C507 VTAIL.n468 B 0.020832f
C508 VTAIL.n469 B 0.009332f
C509 VTAIL.n470 B 0.008813f
C510 VTAIL.n471 B 0.016402f
C511 VTAIL.n472 B 0.016402f
C512 VTAIL.n473 B 0.008813f
C513 VTAIL.n474 B 0.009332f
C514 VTAIL.n475 B 0.020832f
C515 VTAIL.n476 B 0.020832f
C516 VTAIL.n477 B 0.009332f
C517 VTAIL.n478 B 0.008813f
C518 VTAIL.n479 B 0.016402f
C519 VTAIL.n480 B 0.016402f
C520 VTAIL.n481 B 0.008813f
C521 VTAIL.n482 B 0.009332f
C522 VTAIL.n483 B 0.020832f
C523 VTAIL.n484 B 0.042162f
C524 VTAIL.n485 B 0.009332f
C525 VTAIL.n486 B 0.008813f
C526 VTAIL.n487 B 0.035447f
C527 VTAIL.n488 B 0.023211f
C528 VTAIL.n489 B 0.077542f
C529 VTAIL.n490 B 0.021394f
C530 VTAIL.n491 B 0.016402f
C531 VTAIL.n492 B 0.008813f
C532 VTAIL.n493 B 0.020832f
C533 VTAIL.n494 B 0.009332f
C534 VTAIL.n495 B 0.016402f
C535 VTAIL.n496 B 0.008813f
C536 VTAIL.n497 B 0.020832f
C537 VTAIL.n498 B 0.009073f
C538 VTAIL.n499 B 0.016402f
C539 VTAIL.n500 B 0.009073f
C540 VTAIL.n501 B 0.008813f
C541 VTAIL.n502 B 0.020832f
C542 VTAIL.n503 B 0.020832f
C543 VTAIL.n504 B 0.009332f
C544 VTAIL.n505 B 0.016402f
C545 VTAIL.n506 B 0.008813f
C546 VTAIL.n507 B 0.020832f
C547 VTAIL.n508 B 0.009332f
C548 VTAIL.n509 B 0.016402f
C549 VTAIL.n510 B 0.008813f
C550 VTAIL.n511 B 0.020832f
C551 VTAIL.n512 B 0.009332f
C552 VTAIL.n513 B 0.016402f
C553 VTAIL.n514 B 0.008813f
C554 VTAIL.n515 B 0.020832f
C555 VTAIL.n516 B 0.009332f
C556 VTAIL.n517 B 0.016402f
C557 VTAIL.n518 B 0.008813f
C558 VTAIL.n519 B 0.020832f
C559 VTAIL.n520 B 0.009332f
C560 VTAIL.n521 B 1.24826f
C561 VTAIL.n522 B 0.008813f
C562 VTAIL.t4 B 0.034485f
C563 VTAIL.n523 B 0.116885f
C564 VTAIL.n524 B 0.012306f
C565 VTAIL.n525 B 0.015624f
C566 VTAIL.n526 B 0.020832f
C567 VTAIL.n527 B 0.009332f
C568 VTAIL.n528 B 0.008813f
C569 VTAIL.n529 B 0.016402f
C570 VTAIL.n530 B 0.016402f
C571 VTAIL.n531 B 0.008813f
C572 VTAIL.n532 B 0.009332f
C573 VTAIL.n533 B 0.020832f
C574 VTAIL.n534 B 0.020832f
C575 VTAIL.n535 B 0.009332f
C576 VTAIL.n536 B 0.008813f
C577 VTAIL.n537 B 0.016402f
C578 VTAIL.n538 B 0.016402f
C579 VTAIL.n539 B 0.008813f
C580 VTAIL.n540 B 0.009332f
C581 VTAIL.n541 B 0.020832f
C582 VTAIL.n542 B 0.020832f
C583 VTAIL.n543 B 0.009332f
C584 VTAIL.n544 B 0.008813f
C585 VTAIL.n545 B 0.016402f
C586 VTAIL.n546 B 0.016402f
C587 VTAIL.n547 B 0.008813f
C588 VTAIL.n548 B 0.009332f
C589 VTAIL.n549 B 0.020832f
C590 VTAIL.n550 B 0.020832f
C591 VTAIL.n551 B 0.009332f
C592 VTAIL.n552 B 0.008813f
C593 VTAIL.n553 B 0.016402f
C594 VTAIL.n554 B 0.016402f
C595 VTAIL.n555 B 0.008813f
C596 VTAIL.n556 B 0.009332f
C597 VTAIL.n557 B 0.020832f
C598 VTAIL.n558 B 0.020832f
C599 VTAIL.n559 B 0.009332f
C600 VTAIL.n560 B 0.008813f
C601 VTAIL.n561 B 0.016402f
C602 VTAIL.n562 B 0.016402f
C603 VTAIL.n563 B 0.008813f
C604 VTAIL.n564 B 0.009332f
C605 VTAIL.n565 B 0.020832f
C606 VTAIL.n566 B 0.020832f
C607 VTAIL.n567 B 0.009332f
C608 VTAIL.n568 B 0.008813f
C609 VTAIL.n569 B 0.016402f
C610 VTAIL.n570 B 0.016402f
C611 VTAIL.n571 B 0.008813f
C612 VTAIL.n572 B 0.009332f
C613 VTAIL.n573 B 0.020832f
C614 VTAIL.n574 B 0.020832f
C615 VTAIL.n575 B 0.009332f
C616 VTAIL.n576 B 0.008813f
C617 VTAIL.n577 B 0.016402f
C618 VTAIL.n578 B 0.016402f
C619 VTAIL.n579 B 0.008813f
C620 VTAIL.n580 B 0.009332f
C621 VTAIL.n581 B 0.020832f
C622 VTAIL.n582 B 0.042162f
C623 VTAIL.n583 B 0.009332f
C624 VTAIL.n584 B 0.008813f
C625 VTAIL.n585 B 0.035447f
C626 VTAIL.n586 B 0.023211f
C627 VTAIL.n587 B 0.077542f
C628 VTAIL.n588 B 0.021394f
C629 VTAIL.n589 B 0.016402f
C630 VTAIL.n590 B 0.008813f
C631 VTAIL.n591 B 0.020832f
C632 VTAIL.n592 B 0.009332f
C633 VTAIL.n593 B 0.016402f
C634 VTAIL.n594 B 0.008813f
C635 VTAIL.n595 B 0.020832f
C636 VTAIL.n596 B 0.009073f
C637 VTAIL.n597 B 0.016402f
C638 VTAIL.n598 B 0.009073f
C639 VTAIL.n599 B 0.008813f
C640 VTAIL.n600 B 0.020832f
C641 VTAIL.n601 B 0.020832f
C642 VTAIL.n602 B 0.009332f
C643 VTAIL.n603 B 0.016402f
C644 VTAIL.n604 B 0.008813f
C645 VTAIL.n605 B 0.020832f
C646 VTAIL.n606 B 0.009332f
C647 VTAIL.n607 B 0.016402f
C648 VTAIL.n608 B 0.008813f
C649 VTAIL.n609 B 0.020832f
C650 VTAIL.n610 B 0.009332f
C651 VTAIL.n611 B 0.016402f
C652 VTAIL.n612 B 0.008813f
C653 VTAIL.n613 B 0.020832f
C654 VTAIL.n614 B 0.009332f
C655 VTAIL.n615 B 0.016402f
C656 VTAIL.n616 B 0.008813f
C657 VTAIL.n617 B 0.020832f
C658 VTAIL.n618 B 0.009332f
C659 VTAIL.n619 B 1.24826f
C660 VTAIL.n620 B 0.008813f
C661 VTAIL.t5 B 0.034485f
C662 VTAIL.n621 B 0.116885f
C663 VTAIL.n622 B 0.012306f
C664 VTAIL.n623 B 0.015624f
C665 VTAIL.n624 B 0.020832f
C666 VTAIL.n625 B 0.009332f
C667 VTAIL.n626 B 0.008813f
C668 VTAIL.n627 B 0.016402f
C669 VTAIL.n628 B 0.016402f
C670 VTAIL.n629 B 0.008813f
C671 VTAIL.n630 B 0.009332f
C672 VTAIL.n631 B 0.020832f
C673 VTAIL.n632 B 0.020832f
C674 VTAIL.n633 B 0.009332f
C675 VTAIL.n634 B 0.008813f
C676 VTAIL.n635 B 0.016402f
C677 VTAIL.n636 B 0.016402f
C678 VTAIL.n637 B 0.008813f
C679 VTAIL.n638 B 0.009332f
C680 VTAIL.n639 B 0.020832f
C681 VTAIL.n640 B 0.020832f
C682 VTAIL.n641 B 0.009332f
C683 VTAIL.n642 B 0.008813f
C684 VTAIL.n643 B 0.016402f
C685 VTAIL.n644 B 0.016402f
C686 VTAIL.n645 B 0.008813f
C687 VTAIL.n646 B 0.009332f
C688 VTAIL.n647 B 0.020832f
C689 VTAIL.n648 B 0.020832f
C690 VTAIL.n649 B 0.009332f
C691 VTAIL.n650 B 0.008813f
C692 VTAIL.n651 B 0.016402f
C693 VTAIL.n652 B 0.016402f
C694 VTAIL.n653 B 0.008813f
C695 VTAIL.n654 B 0.009332f
C696 VTAIL.n655 B 0.020832f
C697 VTAIL.n656 B 0.020832f
C698 VTAIL.n657 B 0.009332f
C699 VTAIL.n658 B 0.008813f
C700 VTAIL.n659 B 0.016402f
C701 VTAIL.n660 B 0.016402f
C702 VTAIL.n661 B 0.008813f
C703 VTAIL.n662 B 0.009332f
C704 VTAIL.n663 B 0.020832f
C705 VTAIL.n664 B 0.020832f
C706 VTAIL.n665 B 0.009332f
C707 VTAIL.n666 B 0.008813f
C708 VTAIL.n667 B 0.016402f
C709 VTAIL.n668 B 0.016402f
C710 VTAIL.n669 B 0.008813f
C711 VTAIL.n670 B 0.009332f
C712 VTAIL.n671 B 0.020832f
C713 VTAIL.n672 B 0.020832f
C714 VTAIL.n673 B 0.009332f
C715 VTAIL.n674 B 0.008813f
C716 VTAIL.n675 B 0.016402f
C717 VTAIL.n676 B 0.016402f
C718 VTAIL.n677 B 0.008813f
C719 VTAIL.n678 B 0.009332f
C720 VTAIL.n679 B 0.020832f
C721 VTAIL.n680 B 0.042162f
C722 VTAIL.n681 B 0.009332f
C723 VTAIL.n682 B 0.008813f
C724 VTAIL.n683 B 0.035447f
C725 VTAIL.n684 B 0.023211f
C726 VTAIL.n685 B 1.1088f
C727 VTAIL.n686 B 0.021394f
C728 VTAIL.n687 B 0.016402f
C729 VTAIL.n688 B 0.008813f
C730 VTAIL.n689 B 0.020832f
C731 VTAIL.n690 B 0.009332f
C732 VTAIL.n691 B 0.016402f
C733 VTAIL.n692 B 0.008813f
C734 VTAIL.n693 B 0.020832f
C735 VTAIL.n694 B 0.009073f
C736 VTAIL.n695 B 0.016402f
C737 VTAIL.n696 B 0.009332f
C738 VTAIL.n697 B 0.020832f
C739 VTAIL.n698 B 0.009332f
C740 VTAIL.n699 B 0.016402f
C741 VTAIL.n700 B 0.008813f
C742 VTAIL.n701 B 0.020832f
C743 VTAIL.n702 B 0.009332f
C744 VTAIL.n703 B 0.016402f
C745 VTAIL.n704 B 0.008813f
C746 VTAIL.n705 B 0.020832f
C747 VTAIL.n706 B 0.009332f
C748 VTAIL.n707 B 0.016402f
C749 VTAIL.n708 B 0.008813f
C750 VTAIL.n709 B 0.020832f
C751 VTAIL.n710 B 0.009332f
C752 VTAIL.n711 B 0.016402f
C753 VTAIL.n712 B 0.008813f
C754 VTAIL.n713 B 0.020832f
C755 VTAIL.n714 B 0.009332f
C756 VTAIL.n715 B 1.24826f
C757 VTAIL.n716 B 0.008813f
C758 VTAIL.t2 B 0.034485f
C759 VTAIL.n717 B 0.116885f
C760 VTAIL.n718 B 0.012306f
C761 VTAIL.n719 B 0.015624f
C762 VTAIL.n720 B 0.020832f
C763 VTAIL.n721 B 0.009332f
C764 VTAIL.n722 B 0.008813f
C765 VTAIL.n723 B 0.016402f
C766 VTAIL.n724 B 0.016402f
C767 VTAIL.n725 B 0.008813f
C768 VTAIL.n726 B 0.009332f
C769 VTAIL.n727 B 0.020832f
C770 VTAIL.n728 B 0.020832f
C771 VTAIL.n729 B 0.009332f
C772 VTAIL.n730 B 0.008813f
C773 VTAIL.n731 B 0.016402f
C774 VTAIL.n732 B 0.016402f
C775 VTAIL.n733 B 0.008813f
C776 VTAIL.n734 B 0.009332f
C777 VTAIL.n735 B 0.020832f
C778 VTAIL.n736 B 0.020832f
C779 VTAIL.n737 B 0.009332f
C780 VTAIL.n738 B 0.008813f
C781 VTAIL.n739 B 0.016402f
C782 VTAIL.n740 B 0.016402f
C783 VTAIL.n741 B 0.008813f
C784 VTAIL.n742 B 0.009332f
C785 VTAIL.n743 B 0.020832f
C786 VTAIL.n744 B 0.020832f
C787 VTAIL.n745 B 0.009332f
C788 VTAIL.n746 B 0.008813f
C789 VTAIL.n747 B 0.016402f
C790 VTAIL.n748 B 0.016402f
C791 VTAIL.n749 B 0.008813f
C792 VTAIL.n750 B 0.009332f
C793 VTAIL.n751 B 0.020832f
C794 VTAIL.n752 B 0.020832f
C795 VTAIL.n753 B 0.009332f
C796 VTAIL.n754 B 0.008813f
C797 VTAIL.n755 B 0.016402f
C798 VTAIL.n756 B 0.016402f
C799 VTAIL.n757 B 0.008813f
C800 VTAIL.n758 B 0.008813f
C801 VTAIL.n759 B 0.009332f
C802 VTAIL.n760 B 0.020832f
C803 VTAIL.n761 B 0.020832f
C804 VTAIL.n762 B 0.020832f
C805 VTAIL.n763 B 0.009073f
C806 VTAIL.n764 B 0.008813f
C807 VTAIL.n765 B 0.016402f
C808 VTAIL.n766 B 0.016402f
C809 VTAIL.n767 B 0.008813f
C810 VTAIL.n768 B 0.009332f
C811 VTAIL.n769 B 0.020832f
C812 VTAIL.n770 B 0.020832f
C813 VTAIL.n771 B 0.009332f
C814 VTAIL.n772 B 0.008813f
C815 VTAIL.n773 B 0.016402f
C816 VTAIL.n774 B 0.016402f
C817 VTAIL.n775 B 0.008813f
C818 VTAIL.n776 B 0.009332f
C819 VTAIL.n777 B 0.020832f
C820 VTAIL.n778 B 0.042162f
C821 VTAIL.n779 B 0.009332f
C822 VTAIL.n780 B 0.008813f
C823 VTAIL.n781 B 0.035447f
C824 VTAIL.n782 B 0.023211f
C825 VTAIL.n783 B 1.08567f
C826 VP.t0 B 1.47841f
C827 VP.t3 B 1.47843f
C828 VP.n0 B 2.04715f
C829 VP.n1 B 3.98171f
C830 VP.t1 B 1.46474f
C831 VP.n2 B 0.558294f
C832 VP.t2 B 1.46474f
C833 VP.n3 B 0.558294f
C834 VP.n4 B 0.041788f
.ends

