* NGSPICE file created from diff_pair_sample_1233.ext - technology: sky130A

.subckt diff_pair_sample_1233 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.61
X1 VDD2.t9 VN.t0 VTAIL.t0 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X2 VTAIL.t5 VN.t1 VDD2.t8 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X3 VTAIL.t7 VP.t1 VDD1.t8 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X4 VDD2.t7 VN.t2 VTAIL.t1 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X5 VDD1.t7 VP.t2 VTAIL.t15 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.61
X6 VTAIL.t8 VP.t3 VDD1.t6 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X7 VTAIL.t4 VN.t3 VDD2.t6 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X8 VDD1.t5 VP.t4 VTAIL.t12 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X9 VDD2.t5 VN.t4 VTAIL.t3 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.61
X10 VDD2.t4 VN.t5 VTAIL.t16 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.61
X11 VDD1.t4 VP.t5 VTAIL.t10 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X12 VTAIL.t17 VN.t6 VDD2.t3 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X13 B.t11 B.t9 B.t10 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.61
X14 B.t8 B.t6 B.t7 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.61
X15 VTAIL.t9 VP.t6 VDD1.t3 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X16 VTAIL.t18 VN.t7 VDD2.t2 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X17 B.t5 B.t3 B.t4 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.61
X18 VTAIL.t13 VP.t7 VDD1.t2 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.39105 ps=2.7 w=2.37 l=0.61
X19 VDD2.t1 VN.t8 VTAIL.t19 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.61
X20 B.t2 B.t0 B.t1 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0 ps=0 w=2.37 l=0.61
X21 VDD1.t1 VP.t8 VTAIL.t6 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.9243 pd=5.52 as=0.39105 ps=2.7 w=2.37 l=0.61
X22 VDD2.t0 VN.t9 VTAIL.t2 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.61
X23 VDD1.t0 VP.t9 VTAIL.t14 w_n2098_n1442# sky130_fd_pr__pfet_01v8 ad=0.39105 pd=2.7 as=0.9243 ps=5.52 w=2.37 l=0.61
R0 VP.n6 VP.t8 185.097
R1 VP.n23 VP.n22 161.3
R2 VP.n9 VP.n4 161.3
R3 VP.n10 VP.n3 161.3
R4 VP.n12 VP.n11 161.3
R5 VP.n21 VP.n0 161.3
R6 VP.n20 VP.n19 161.3
R7 VP.n17 VP.n16 161.3
R8 VP.n15 VP.n2 161.3
R9 VP.n14 VP.n13 161.3
R10 VP.n14 VP.t2 158.429
R11 VP.n16 VP.t6 158.429
R12 VP.n1 VP.t4 158.429
R13 VP.n20 VP.t3 158.429
R14 VP.n22 VP.t9 158.429
R15 VP.n11 VP.t0 158.429
R16 VP.n9 VP.t7 158.429
R17 VP.n8 VP.t5 158.429
R18 VP.n7 VP.t1 158.429
R19 VP.n8 VP.n5 80.6037
R20 VP.n18 VP.n1 80.6037
R21 VP.n16 VP.n1 48.2005
R22 VP.n20 VP.n1 48.2005
R23 VP.n9 VP.n8 48.2005
R24 VP.n8 VP.n7 48.2005
R25 VP.n15 VP.n14 47.4702
R26 VP.n22 VP.n21 47.4702
R27 VP.n11 VP.n10 47.4702
R28 VP.n6 VP.n5 45.2144
R29 VP.n13 VP.n12 35.0308
R30 VP.n7 VP.n6 13.6377
R31 VP.n16 VP.n15 0.730803
R32 VP.n21 VP.n20 0.730803
R33 VP.n10 VP.n9 0.730803
R34 VP.n5 VP.n4 0.285035
R35 VP.n18 VP.n17 0.285035
R36 VP.n19 VP.n18 0.285035
R37 VP.n4 VP.n3 0.189894
R38 VP.n12 VP.n3 0.189894
R39 VP.n13 VP.n2 0.189894
R40 VP.n17 VP.n2 0.189894
R41 VP.n19 VP.n0 0.189894
R42 VP.n23 VP.n0 0.189894
R43 VP VP.n23 0.0516364
R44 VTAIL.n16 VTAIL.t11 168.97
R45 VTAIL.n11 VTAIL.t3 168.97
R46 VTAIL.n17 VTAIL.t2 168.97
R47 VTAIL.n2 VTAIL.t14 168.97
R48 VTAIL.n15 VTAIL.n14 155.256
R49 VTAIL.n13 VTAIL.n12 155.256
R50 VTAIL.n10 VTAIL.n9 155.256
R51 VTAIL.n8 VTAIL.n7 155.256
R52 VTAIL.n19 VTAIL.n18 155.255
R53 VTAIL.n1 VTAIL.n0 155.255
R54 VTAIL.n4 VTAIL.n3 155.255
R55 VTAIL.n6 VTAIL.n5 155.255
R56 VTAIL.n8 VTAIL.n6 16.0307
R57 VTAIL.n17 VTAIL.n16 15.2203
R58 VTAIL.n18 VTAIL.t1 13.7157
R59 VTAIL.n18 VTAIL.t17 13.7157
R60 VTAIL.n0 VTAIL.t19 13.7157
R61 VTAIL.n0 VTAIL.t5 13.7157
R62 VTAIL.n3 VTAIL.t12 13.7157
R63 VTAIL.n3 VTAIL.t8 13.7157
R64 VTAIL.n5 VTAIL.t15 13.7157
R65 VTAIL.n5 VTAIL.t9 13.7157
R66 VTAIL.n14 VTAIL.t10 13.7157
R67 VTAIL.n14 VTAIL.t13 13.7157
R68 VTAIL.n12 VTAIL.t6 13.7157
R69 VTAIL.n12 VTAIL.t7 13.7157
R70 VTAIL.n9 VTAIL.t0 13.7157
R71 VTAIL.n9 VTAIL.t18 13.7157
R72 VTAIL.n7 VTAIL.t16 13.7157
R73 VTAIL.n7 VTAIL.t4 13.7157
R74 VTAIL.n13 VTAIL.n11 0.8755
R75 VTAIL.n2 VTAIL.n1 0.8755
R76 VTAIL.n10 VTAIL.n8 0.810845
R77 VTAIL.n11 VTAIL.n10 0.810845
R78 VTAIL.n15 VTAIL.n13 0.810845
R79 VTAIL.n16 VTAIL.n15 0.810845
R80 VTAIL.n6 VTAIL.n4 0.810845
R81 VTAIL.n4 VTAIL.n2 0.810845
R82 VTAIL.n19 VTAIL.n17 0.810845
R83 VTAIL VTAIL.n1 0.666448
R84 VTAIL VTAIL.n19 0.144897
R85 VDD1.n1 VDD1.t1 186.459
R86 VDD1.n3 VDD1.t7 186.459
R87 VDD1.n5 VDD1.n4 172.487
R88 VDD1.n7 VDD1.n6 171.934
R89 VDD1.n1 VDD1.n0 171.934
R90 VDD1.n3 VDD1.n2 171.934
R91 VDD1.n7 VDD1.n5 30.5957
R92 VDD1.n6 VDD1.t2 13.7157
R93 VDD1.n6 VDD1.t9 13.7157
R94 VDD1.n0 VDD1.t8 13.7157
R95 VDD1.n0 VDD1.t4 13.7157
R96 VDD1.n4 VDD1.t6 13.7157
R97 VDD1.n4 VDD1.t0 13.7157
R98 VDD1.n2 VDD1.t3 13.7157
R99 VDD1.n2 VDD1.t5 13.7157
R100 VDD1 VDD1.n7 0.550069
R101 VDD1 VDD1.n1 0.261276
R102 VDD1.n5 VDD1.n3 0.14774
R103 VN.n3 VN.t8 185.097
R104 VN.n13 VN.t4 185.097
R105 VN.n9 VN.n8 161.3
R106 VN.n19 VN.n18 161.3
R107 VN.n17 VN.n10 161.3
R108 VN.n16 VN.n15 161.3
R109 VN.n7 VN.n0 161.3
R110 VN.n6 VN.n5 161.3
R111 VN.n2 VN.t1 158.429
R112 VN.n1 VN.t2 158.429
R113 VN.n6 VN.t6 158.429
R114 VN.n8 VN.t9 158.429
R115 VN.n12 VN.t7 158.429
R116 VN.n11 VN.t0 158.429
R117 VN.n16 VN.t3 158.429
R118 VN.n18 VN.t5 158.429
R119 VN.n14 VN.n11 80.6037
R120 VN.n4 VN.n1 80.6037
R121 VN.n2 VN.n1 48.2005
R122 VN.n6 VN.n1 48.2005
R123 VN.n12 VN.n11 48.2005
R124 VN.n16 VN.n11 48.2005
R125 VN.n8 VN.n7 47.4702
R126 VN.n18 VN.n17 47.4702
R127 VN.n14 VN.n13 45.2144
R128 VN.n4 VN.n3 45.2144
R129 VN VN.n19 35.4115
R130 VN.n3 VN.n2 13.6377
R131 VN.n13 VN.n12 13.6377
R132 VN.n7 VN.n6 0.730803
R133 VN.n17 VN.n16 0.730803
R134 VN.n15 VN.n14 0.285035
R135 VN.n5 VN.n4 0.285035
R136 VN.n19 VN.n10 0.189894
R137 VN.n15 VN.n10 0.189894
R138 VN.n5 VN.n0 0.189894
R139 VN.n9 VN.n0 0.189894
R140 VN VN.n9 0.0516364
R141 VDD2.n1 VDD2.t1 186.459
R142 VDD2.n4 VDD2.t4 185.649
R143 VDD2.n3 VDD2.n2 172.487
R144 VDD2 VDD2.n7 172.483
R145 VDD2.n6 VDD2.n5 171.934
R146 VDD2.n1 VDD2.n0 171.934
R147 VDD2.n4 VDD2.n3 29.6075
R148 VDD2.n7 VDD2.t2 13.7157
R149 VDD2.n7 VDD2.t5 13.7157
R150 VDD2.n5 VDD2.t6 13.7157
R151 VDD2.n5 VDD2.t9 13.7157
R152 VDD2.n2 VDD2.t3 13.7157
R153 VDD2.n2 VDD2.t0 13.7157
R154 VDD2.n0 VDD2.t8 13.7157
R155 VDD2.n0 VDD2.t7 13.7157
R156 VDD2.n6 VDD2.n4 0.810845
R157 VDD2 VDD2.n6 0.261276
R158 VDD2.n3 VDD2.n1 0.14774
R159 B.n185 B.n62 585
R160 B.n184 B.n183 585
R161 B.n182 B.n63 585
R162 B.n181 B.n180 585
R163 B.n179 B.n64 585
R164 B.n178 B.n177 585
R165 B.n176 B.n65 585
R166 B.n175 B.n174 585
R167 B.n173 B.n66 585
R168 B.n172 B.n171 585
R169 B.n170 B.n67 585
R170 B.n169 B.n168 585
R171 B.n167 B.n68 585
R172 B.n165 B.n164 585
R173 B.n163 B.n71 585
R174 B.n162 B.n161 585
R175 B.n160 B.n72 585
R176 B.n159 B.n158 585
R177 B.n157 B.n73 585
R178 B.n156 B.n155 585
R179 B.n154 B.n74 585
R180 B.n153 B.n152 585
R181 B.n151 B.n75 585
R182 B.n150 B.n149 585
R183 B.n145 B.n76 585
R184 B.n144 B.n143 585
R185 B.n142 B.n77 585
R186 B.n141 B.n140 585
R187 B.n139 B.n78 585
R188 B.n138 B.n137 585
R189 B.n136 B.n79 585
R190 B.n135 B.n134 585
R191 B.n133 B.n80 585
R192 B.n132 B.n131 585
R193 B.n130 B.n81 585
R194 B.n129 B.n128 585
R195 B.n187 B.n186 585
R196 B.n188 B.n61 585
R197 B.n190 B.n189 585
R198 B.n191 B.n60 585
R199 B.n193 B.n192 585
R200 B.n194 B.n59 585
R201 B.n196 B.n195 585
R202 B.n197 B.n58 585
R203 B.n199 B.n198 585
R204 B.n200 B.n57 585
R205 B.n202 B.n201 585
R206 B.n203 B.n56 585
R207 B.n205 B.n204 585
R208 B.n206 B.n55 585
R209 B.n208 B.n207 585
R210 B.n209 B.n54 585
R211 B.n211 B.n210 585
R212 B.n212 B.n53 585
R213 B.n214 B.n213 585
R214 B.n215 B.n52 585
R215 B.n217 B.n216 585
R216 B.n218 B.n51 585
R217 B.n220 B.n219 585
R218 B.n221 B.n50 585
R219 B.n223 B.n222 585
R220 B.n224 B.n49 585
R221 B.n226 B.n225 585
R222 B.n227 B.n48 585
R223 B.n229 B.n228 585
R224 B.n230 B.n47 585
R225 B.n232 B.n231 585
R226 B.n233 B.n46 585
R227 B.n235 B.n234 585
R228 B.n236 B.n45 585
R229 B.n238 B.n237 585
R230 B.n239 B.n44 585
R231 B.n241 B.n240 585
R232 B.n242 B.n43 585
R233 B.n244 B.n243 585
R234 B.n245 B.n42 585
R235 B.n247 B.n246 585
R236 B.n248 B.n41 585
R237 B.n250 B.n249 585
R238 B.n251 B.n40 585
R239 B.n253 B.n252 585
R240 B.n254 B.n39 585
R241 B.n256 B.n255 585
R242 B.n257 B.n38 585
R243 B.n259 B.n258 585
R244 B.n260 B.n37 585
R245 B.n315 B.n14 585
R246 B.n314 B.n313 585
R247 B.n312 B.n15 585
R248 B.n311 B.n310 585
R249 B.n309 B.n16 585
R250 B.n308 B.n307 585
R251 B.n306 B.n17 585
R252 B.n305 B.n304 585
R253 B.n303 B.n18 585
R254 B.n302 B.n301 585
R255 B.n300 B.n19 585
R256 B.n299 B.n298 585
R257 B.n297 B.n20 585
R258 B.n296 B.n295 585
R259 B.n294 B.n21 585
R260 B.n293 B.n292 585
R261 B.n291 B.n25 585
R262 B.n290 B.n289 585
R263 B.n288 B.n26 585
R264 B.n287 B.n286 585
R265 B.n285 B.n27 585
R266 B.n284 B.n283 585
R267 B.n282 B.n28 585
R268 B.n280 B.n279 585
R269 B.n278 B.n31 585
R270 B.n277 B.n276 585
R271 B.n275 B.n32 585
R272 B.n274 B.n273 585
R273 B.n272 B.n33 585
R274 B.n271 B.n270 585
R275 B.n269 B.n34 585
R276 B.n268 B.n267 585
R277 B.n266 B.n35 585
R278 B.n265 B.n264 585
R279 B.n263 B.n36 585
R280 B.n262 B.n261 585
R281 B.n317 B.n316 585
R282 B.n318 B.n13 585
R283 B.n320 B.n319 585
R284 B.n321 B.n12 585
R285 B.n323 B.n322 585
R286 B.n324 B.n11 585
R287 B.n326 B.n325 585
R288 B.n327 B.n10 585
R289 B.n329 B.n328 585
R290 B.n330 B.n9 585
R291 B.n332 B.n331 585
R292 B.n333 B.n8 585
R293 B.n335 B.n334 585
R294 B.n336 B.n7 585
R295 B.n338 B.n337 585
R296 B.n339 B.n6 585
R297 B.n341 B.n340 585
R298 B.n342 B.n5 585
R299 B.n344 B.n343 585
R300 B.n345 B.n4 585
R301 B.n347 B.n346 585
R302 B.n348 B.n3 585
R303 B.n350 B.n349 585
R304 B.n351 B.n0 585
R305 B.n2 B.n1 585
R306 B.n94 B.n93 585
R307 B.n96 B.n95 585
R308 B.n97 B.n92 585
R309 B.n99 B.n98 585
R310 B.n100 B.n91 585
R311 B.n102 B.n101 585
R312 B.n103 B.n90 585
R313 B.n105 B.n104 585
R314 B.n106 B.n89 585
R315 B.n108 B.n107 585
R316 B.n109 B.n88 585
R317 B.n111 B.n110 585
R318 B.n112 B.n87 585
R319 B.n114 B.n113 585
R320 B.n115 B.n86 585
R321 B.n117 B.n116 585
R322 B.n118 B.n85 585
R323 B.n120 B.n119 585
R324 B.n121 B.n84 585
R325 B.n123 B.n122 585
R326 B.n124 B.n83 585
R327 B.n126 B.n125 585
R328 B.n127 B.n82 585
R329 B.n129 B.n82 545.355
R330 B.n187 B.n62 545.355
R331 B.n261 B.n260 545.355
R332 B.n316 B.n315 545.355
R333 B.n146 B.t0 297.87
R334 B.n69 B.t6 297.87
R335 B.n29 B.t3 297.87
R336 B.n22 B.t9 297.87
R337 B.n353 B.n352 256.663
R338 B.n352 B.n351 235.042
R339 B.n352 B.n2 235.042
R340 B.n69 B.t7 193.315
R341 B.n29 B.t5 193.315
R342 B.n146 B.t1 193.315
R343 B.n22 B.t11 193.315
R344 B.n70 B.t8 175.085
R345 B.n30 B.t4 175.085
R346 B.n147 B.t2 175.085
R347 B.n23 B.t10 175.085
R348 B.n130 B.n129 163.367
R349 B.n131 B.n130 163.367
R350 B.n131 B.n80 163.367
R351 B.n135 B.n80 163.367
R352 B.n136 B.n135 163.367
R353 B.n137 B.n136 163.367
R354 B.n137 B.n78 163.367
R355 B.n141 B.n78 163.367
R356 B.n142 B.n141 163.367
R357 B.n143 B.n142 163.367
R358 B.n143 B.n76 163.367
R359 B.n150 B.n76 163.367
R360 B.n151 B.n150 163.367
R361 B.n152 B.n151 163.367
R362 B.n152 B.n74 163.367
R363 B.n156 B.n74 163.367
R364 B.n157 B.n156 163.367
R365 B.n158 B.n157 163.367
R366 B.n158 B.n72 163.367
R367 B.n162 B.n72 163.367
R368 B.n163 B.n162 163.367
R369 B.n164 B.n163 163.367
R370 B.n164 B.n68 163.367
R371 B.n169 B.n68 163.367
R372 B.n170 B.n169 163.367
R373 B.n171 B.n170 163.367
R374 B.n171 B.n66 163.367
R375 B.n175 B.n66 163.367
R376 B.n176 B.n175 163.367
R377 B.n177 B.n176 163.367
R378 B.n177 B.n64 163.367
R379 B.n181 B.n64 163.367
R380 B.n182 B.n181 163.367
R381 B.n183 B.n182 163.367
R382 B.n183 B.n62 163.367
R383 B.n260 B.n259 163.367
R384 B.n259 B.n38 163.367
R385 B.n255 B.n38 163.367
R386 B.n255 B.n254 163.367
R387 B.n254 B.n253 163.367
R388 B.n253 B.n40 163.367
R389 B.n249 B.n40 163.367
R390 B.n249 B.n248 163.367
R391 B.n248 B.n247 163.367
R392 B.n247 B.n42 163.367
R393 B.n243 B.n42 163.367
R394 B.n243 B.n242 163.367
R395 B.n242 B.n241 163.367
R396 B.n241 B.n44 163.367
R397 B.n237 B.n44 163.367
R398 B.n237 B.n236 163.367
R399 B.n236 B.n235 163.367
R400 B.n235 B.n46 163.367
R401 B.n231 B.n46 163.367
R402 B.n231 B.n230 163.367
R403 B.n230 B.n229 163.367
R404 B.n229 B.n48 163.367
R405 B.n225 B.n48 163.367
R406 B.n225 B.n224 163.367
R407 B.n224 B.n223 163.367
R408 B.n223 B.n50 163.367
R409 B.n219 B.n50 163.367
R410 B.n219 B.n218 163.367
R411 B.n218 B.n217 163.367
R412 B.n217 B.n52 163.367
R413 B.n213 B.n52 163.367
R414 B.n213 B.n212 163.367
R415 B.n212 B.n211 163.367
R416 B.n211 B.n54 163.367
R417 B.n207 B.n54 163.367
R418 B.n207 B.n206 163.367
R419 B.n206 B.n205 163.367
R420 B.n205 B.n56 163.367
R421 B.n201 B.n56 163.367
R422 B.n201 B.n200 163.367
R423 B.n200 B.n199 163.367
R424 B.n199 B.n58 163.367
R425 B.n195 B.n58 163.367
R426 B.n195 B.n194 163.367
R427 B.n194 B.n193 163.367
R428 B.n193 B.n60 163.367
R429 B.n189 B.n60 163.367
R430 B.n189 B.n188 163.367
R431 B.n188 B.n187 163.367
R432 B.n315 B.n314 163.367
R433 B.n314 B.n15 163.367
R434 B.n310 B.n15 163.367
R435 B.n310 B.n309 163.367
R436 B.n309 B.n308 163.367
R437 B.n308 B.n17 163.367
R438 B.n304 B.n17 163.367
R439 B.n304 B.n303 163.367
R440 B.n303 B.n302 163.367
R441 B.n302 B.n19 163.367
R442 B.n298 B.n19 163.367
R443 B.n298 B.n297 163.367
R444 B.n297 B.n296 163.367
R445 B.n296 B.n21 163.367
R446 B.n292 B.n21 163.367
R447 B.n292 B.n291 163.367
R448 B.n291 B.n290 163.367
R449 B.n290 B.n26 163.367
R450 B.n286 B.n26 163.367
R451 B.n286 B.n285 163.367
R452 B.n285 B.n284 163.367
R453 B.n284 B.n28 163.367
R454 B.n279 B.n28 163.367
R455 B.n279 B.n278 163.367
R456 B.n278 B.n277 163.367
R457 B.n277 B.n32 163.367
R458 B.n273 B.n32 163.367
R459 B.n273 B.n272 163.367
R460 B.n272 B.n271 163.367
R461 B.n271 B.n34 163.367
R462 B.n267 B.n34 163.367
R463 B.n267 B.n266 163.367
R464 B.n266 B.n265 163.367
R465 B.n265 B.n36 163.367
R466 B.n261 B.n36 163.367
R467 B.n316 B.n13 163.367
R468 B.n320 B.n13 163.367
R469 B.n321 B.n320 163.367
R470 B.n322 B.n321 163.367
R471 B.n322 B.n11 163.367
R472 B.n326 B.n11 163.367
R473 B.n327 B.n326 163.367
R474 B.n328 B.n327 163.367
R475 B.n328 B.n9 163.367
R476 B.n332 B.n9 163.367
R477 B.n333 B.n332 163.367
R478 B.n334 B.n333 163.367
R479 B.n334 B.n7 163.367
R480 B.n338 B.n7 163.367
R481 B.n339 B.n338 163.367
R482 B.n340 B.n339 163.367
R483 B.n340 B.n5 163.367
R484 B.n344 B.n5 163.367
R485 B.n345 B.n344 163.367
R486 B.n346 B.n345 163.367
R487 B.n346 B.n3 163.367
R488 B.n350 B.n3 163.367
R489 B.n351 B.n350 163.367
R490 B.n94 B.n2 163.367
R491 B.n95 B.n94 163.367
R492 B.n95 B.n92 163.367
R493 B.n99 B.n92 163.367
R494 B.n100 B.n99 163.367
R495 B.n101 B.n100 163.367
R496 B.n101 B.n90 163.367
R497 B.n105 B.n90 163.367
R498 B.n106 B.n105 163.367
R499 B.n107 B.n106 163.367
R500 B.n107 B.n88 163.367
R501 B.n111 B.n88 163.367
R502 B.n112 B.n111 163.367
R503 B.n113 B.n112 163.367
R504 B.n113 B.n86 163.367
R505 B.n117 B.n86 163.367
R506 B.n118 B.n117 163.367
R507 B.n119 B.n118 163.367
R508 B.n119 B.n84 163.367
R509 B.n123 B.n84 163.367
R510 B.n124 B.n123 163.367
R511 B.n125 B.n124 163.367
R512 B.n125 B.n82 163.367
R513 B.n148 B.n147 59.5399
R514 B.n166 B.n70 59.5399
R515 B.n281 B.n30 59.5399
R516 B.n24 B.n23 59.5399
R517 B.n186 B.n185 35.4346
R518 B.n317 B.n14 35.4346
R519 B.n262 B.n37 35.4346
R520 B.n128 B.n127 35.4346
R521 B.n147 B.n146 18.2308
R522 B.n70 B.n69 18.2308
R523 B.n30 B.n29 18.2308
R524 B.n23 B.n22 18.2308
R525 B B.n353 18.0485
R526 B.n318 B.n317 10.6151
R527 B.n319 B.n318 10.6151
R528 B.n319 B.n12 10.6151
R529 B.n323 B.n12 10.6151
R530 B.n324 B.n323 10.6151
R531 B.n325 B.n324 10.6151
R532 B.n325 B.n10 10.6151
R533 B.n329 B.n10 10.6151
R534 B.n330 B.n329 10.6151
R535 B.n331 B.n330 10.6151
R536 B.n331 B.n8 10.6151
R537 B.n335 B.n8 10.6151
R538 B.n336 B.n335 10.6151
R539 B.n337 B.n336 10.6151
R540 B.n337 B.n6 10.6151
R541 B.n341 B.n6 10.6151
R542 B.n342 B.n341 10.6151
R543 B.n343 B.n342 10.6151
R544 B.n343 B.n4 10.6151
R545 B.n347 B.n4 10.6151
R546 B.n348 B.n347 10.6151
R547 B.n349 B.n348 10.6151
R548 B.n349 B.n0 10.6151
R549 B.n313 B.n14 10.6151
R550 B.n313 B.n312 10.6151
R551 B.n312 B.n311 10.6151
R552 B.n311 B.n16 10.6151
R553 B.n307 B.n16 10.6151
R554 B.n307 B.n306 10.6151
R555 B.n306 B.n305 10.6151
R556 B.n305 B.n18 10.6151
R557 B.n301 B.n18 10.6151
R558 B.n301 B.n300 10.6151
R559 B.n300 B.n299 10.6151
R560 B.n299 B.n20 10.6151
R561 B.n295 B.n294 10.6151
R562 B.n294 B.n293 10.6151
R563 B.n293 B.n25 10.6151
R564 B.n289 B.n25 10.6151
R565 B.n289 B.n288 10.6151
R566 B.n288 B.n287 10.6151
R567 B.n287 B.n27 10.6151
R568 B.n283 B.n27 10.6151
R569 B.n283 B.n282 10.6151
R570 B.n280 B.n31 10.6151
R571 B.n276 B.n31 10.6151
R572 B.n276 B.n275 10.6151
R573 B.n275 B.n274 10.6151
R574 B.n274 B.n33 10.6151
R575 B.n270 B.n33 10.6151
R576 B.n270 B.n269 10.6151
R577 B.n269 B.n268 10.6151
R578 B.n268 B.n35 10.6151
R579 B.n264 B.n35 10.6151
R580 B.n264 B.n263 10.6151
R581 B.n263 B.n262 10.6151
R582 B.n258 B.n37 10.6151
R583 B.n258 B.n257 10.6151
R584 B.n257 B.n256 10.6151
R585 B.n256 B.n39 10.6151
R586 B.n252 B.n39 10.6151
R587 B.n252 B.n251 10.6151
R588 B.n251 B.n250 10.6151
R589 B.n250 B.n41 10.6151
R590 B.n246 B.n41 10.6151
R591 B.n246 B.n245 10.6151
R592 B.n245 B.n244 10.6151
R593 B.n244 B.n43 10.6151
R594 B.n240 B.n43 10.6151
R595 B.n240 B.n239 10.6151
R596 B.n239 B.n238 10.6151
R597 B.n238 B.n45 10.6151
R598 B.n234 B.n45 10.6151
R599 B.n234 B.n233 10.6151
R600 B.n233 B.n232 10.6151
R601 B.n232 B.n47 10.6151
R602 B.n228 B.n47 10.6151
R603 B.n228 B.n227 10.6151
R604 B.n227 B.n226 10.6151
R605 B.n226 B.n49 10.6151
R606 B.n222 B.n49 10.6151
R607 B.n222 B.n221 10.6151
R608 B.n221 B.n220 10.6151
R609 B.n220 B.n51 10.6151
R610 B.n216 B.n51 10.6151
R611 B.n216 B.n215 10.6151
R612 B.n215 B.n214 10.6151
R613 B.n214 B.n53 10.6151
R614 B.n210 B.n53 10.6151
R615 B.n210 B.n209 10.6151
R616 B.n209 B.n208 10.6151
R617 B.n208 B.n55 10.6151
R618 B.n204 B.n55 10.6151
R619 B.n204 B.n203 10.6151
R620 B.n203 B.n202 10.6151
R621 B.n202 B.n57 10.6151
R622 B.n198 B.n57 10.6151
R623 B.n198 B.n197 10.6151
R624 B.n197 B.n196 10.6151
R625 B.n196 B.n59 10.6151
R626 B.n192 B.n59 10.6151
R627 B.n192 B.n191 10.6151
R628 B.n191 B.n190 10.6151
R629 B.n190 B.n61 10.6151
R630 B.n186 B.n61 10.6151
R631 B.n93 B.n1 10.6151
R632 B.n96 B.n93 10.6151
R633 B.n97 B.n96 10.6151
R634 B.n98 B.n97 10.6151
R635 B.n98 B.n91 10.6151
R636 B.n102 B.n91 10.6151
R637 B.n103 B.n102 10.6151
R638 B.n104 B.n103 10.6151
R639 B.n104 B.n89 10.6151
R640 B.n108 B.n89 10.6151
R641 B.n109 B.n108 10.6151
R642 B.n110 B.n109 10.6151
R643 B.n110 B.n87 10.6151
R644 B.n114 B.n87 10.6151
R645 B.n115 B.n114 10.6151
R646 B.n116 B.n115 10.6151
R647 B.n116 B.n85 10.6151
R648 B.n120 B.n85 10.6151
R649 B.n121 B.n120 10.6151
R650 B.n122 B.n121 10.6151
R651 B.n122 B.n83 10.6151
R652 B.n126 B.n83 10.6151
R653 B.n127 B.n126 10.6151
R654 B.n128 B.n81 10.6151
R655 B.n132 B.n81 10.6151
R656 B.n133 B.n132 10.6151
R657 B.n134 B.n133 10.6151
R658 B.n134 B.n79 10.6151
R659 B.n138 B.n79 10.6151
R660 B.n139 B.n138 10.6151
R661 B.n140 B.n139 10.6151
R662 B.n140 B.n77 10.6151
R663 B.n144 B.n77 10.6151
R664 B.n145 B.n144 10.6151
R665 B.n149 B.n145 10.6151
R666 B.n153 B.n75 10.6151
R667 B.n154 B.n153 10.6151
R668 B.n155 B.n154 10.6151
R669 B.n155 B.n73 10.6151
R670 B.n159 B.n73 10.6151
R671 B.n160 B.n159 10.6151
R672 B.n161 B.n160 10.6151
R673 B.n161 B.n71 10.6151
R674 B.n165 B.n71 10.6151
R675 B.n168 B.n167 10.6151
R676 B.n168 B.n67 10.6151
R677 B.n172 B.n67 10.6151
R678 B.n173 B.n172 10.6151
R679 B.n174 B.n173 10.6151
R680 B.n174 B.n65 10.6151
R681 B.n178 B.n65 10.6151
R682 B.n179 B.n178 10.6151
R683 B.n180 B.n179 10.6151
R684 B.n180 B.n63 10.6151
R685 B.n184 B.n63 10.6151
R686 B.n185 B.n184 10.6151
R687 B.n24 B.n20 9.36635
R688 B.n281 B.n280 9.36635
R689 B.n149 B.n148 9.36635
R690 B.n167 B.n166 9.36635
R691 B.n353 B.n0 8.11757
R692 B.n353 B.n1 8.11757
R693 B.n295 B.n24 1.24928
R694 B.n282 B.n281 1.24928
R695 B.n148 B.n75 1.24928
R696 B.n166 B.n165 1.24928
C0 VN w_n2098_n1442# 3.67533f
C1 VP VN 3.68837f
C2 B VDD1 0.966619f
C3 VDD2 VDD1 0.914318f
C4 VTAIL w_n2098_n1442# 1.47508f
C5 VP VTAIL 1.85287f
C6 B VDD2 1.00758f
C7 w_n2098_n1442# VDD1 1.28451f
C8 VTAIL VN 1.83866f
C9 VP VDD1 1.74133f
C10 B w_n2098_n1442# 4.49363f
C11 w_n2098_n1442# VDD2 1.32387f
C12 VP B 1.09859f
C13 VP VDD2 0.335341f
C14 VN VDD1 0.154851f
C15 B VN 0.661189f
C16 VTAIL VDD1 4.92196f
C17 VN VDD2 1.56295f
C18 VP w_n2098_n1442# 3.93886f
C19 B VTAIL 0.953933f
C20 VTAIL VDD2 4.96082f
C21 VDD2 VSUBS 0.795829f
C22 VDD1 VSUBS 0.794107f
C23 VTAIL VSUBS 0.312651f
C24 VN VSUBS 3.56032f
C25 VP VSUBS 1.235044f
C26 B VSUBS 1.982085f
C27 w_n2098_n1442# VSUBS 38.4941f
C28 B.n0 VSUBS 0.007331f
C29 B.n1 VSUBS 0.007331f
C30 B.n2 VSUBS 0.010843f
C31 B.n3 VSUBS 0.008309f
C32 B.n4 VSUBS 0.008309f
C33 B.n5 VSUBS 0.008309f
C34 B.n6 VSUBS 0.008309f
C35 B.n7 VSUBS 0.008309f
C36 B.n8 VSUBS 0.008309f
C37 B.n9 VSUBS 0.008309f
C38 B.n10 VSUBS 0.008309f
C39 B.n11 VSUBS 0.008309f
C40 B.n12 VSUBS 0.008309f
C41 B.n13 VSUBS 0.008309f
C42 B.n14 VSUBS 0.021046f
C43 B.n15 VSUBS 0.008309f
C44 B.n16 VSUBS 0.008309f
C45 B.n17 VSUBS 0.008309f
C46 B.n18 VSUBS 0.008309f
C47 B.n19 VSUBS 0.008309f
C48 B.n20 VSUBS 0.00782f
C49 B.n21 VSUBS 0.008309f
C50 B.t10 VSUBS 0.062888f
C51 B.t11 VSUBS 0.067754f
C52 B.t9 VSUBS 0.079683f
C53 B.n22 VSUBS 0.068962f
C54 B.n23 VSUBS 0.063457f
C55 B.n24 VSUBS 0.019251f
C56 B.n25 VSUBS 0.008309f
C57 B.n26 VSUBS 0.008309f
C58 B.n27 VSUBS 0.008309f
C59 B.n28 VSUBS 0.008309f
C60 B.t4 VSUBS 0.062888f
C61 B.t5 VSUBS 0.067754f
C62 B.t3 VSUBS 0.079683f
C63 B.n29 VSUBS 0.068962f
C64 B.n30 VSUBS 0.063457f
C65 B.n31 VSUBS 0.008309f
C66 B.n32 VSUBS 0.008309f
C67 B.n33 VSUBS 0.008309f
C68 B.n34 VSUBS 0.008309f
C69 B.n35 VSUBS 0.008309f
C70 B.n36 VSUBS 0.008309f
C71 B.n37 VSUBS 0.020009f
C72 B.n38 VSUBS 0.008309f
C73 B.n39 VSUBS 0.008309f
C74 B.n40 VSUBS 0.008309f
C75 B.n41 VSUBS 0.008309f
C76 B.n42 VSUBS 0.008309f
C77 B.n43 VSUBS 0.008309f
C78 B.n44 VSUBS 0.008309f
C79 B.n45 VSUBS 0.008309f
C80 B.n46 VSUBS 0.008309f
C81 B.n47 VSUBS 0.008309f
C82 B.n48 VSUBS 0.008309f
C83 B.n49 VSUBS 0.008309f
C84 B.n50 VSUBS 0.008309f
C85 B.n51 VSUBS 0.008309f
C86 B.n52 VSUBS 0.008309f
C87 B.n53 VSUBS 0.008309f
C88 B.n54 VSUBS 0.008309f
C89 B.n55 VSUBS 0.008309f
C90 B.n56 VSUBS 0.008309f
C91 B.n57 VSUBS 0.008309f
C92 B.n58 VSUBS 0.008309f
C93 B.n59 VSUBS 0.008309f
C94 B.n60 VSUBS 0.008309f
C95 B.n61 VSUBS 0.008309f
C96 B.n62 VSUBS 0.021046f
C97 B.n63 VSUBS 0.008309f
C98 B.n64 VSUBS 0.008309f
C99 B.n65 VSUBS 0.008309f
C100 B.n66 VSUBS 0.008309f
C101 B.n67 VSUBS 0.008309f
C102 B.n68 VSUBS 0.008309f
C103 B.t8 VSUBS 0.062888f
C104 B.t7 VSUBS 0.067754f
C105 B.t6 VSUBS 0.079683f
C106 B.n69 VSUBS 0.068962f
C107 B.n70 VSUBS 0.063457f
C108 B.n71 VSUBS 0.008309f
C109 B.n72 VSUBS 0.008309f
C110 B.n73 VSUBS 0.008309f
C111 B.n74 VSUBS 0.008309f
C112 B.n75 VSUBS 0.004643f
C113 B.n76 VSUBS 0.008309f
C114 B.n77 VSUBS 0.008309f
C115 B.n78 VSUBS 0.008309f
C116 B.n79 VSUBS 0.008309f
C117 B.n80 VSUBS 0.008309f
C118 B.n81 VSUBS 0.008309f
C119 B.n82 VSUBS 0.020009f
C120 B.n83 VSUBS 0.008309f
C121 B.n84 VSUBS 0.008309f
C122 B.n85 VSUBS 0.008309f
C123 B.n86 VSUBS 0.008309f
C124 B.n87 VSUBS 0.008309f
C125 B.n88 VSUBS 0.008309f
C126 B.n89 VSUBS 0.008309f
C127 B.n90 VSUBS 0.008309f
C128 B.n91 VSUBS 0.008309f
C129 B.n92 VSUBS 0.008309f
C130 B.n93 VSUBS 0.008309f
C131 B.n94 VSUBS 0.008309f
C132 B.n95 VSUBS 0.008309f
C133 B.n96 VSUBS 0.008309f
C134 B.n97 VSUBS 0.008309f
C135 B.n98 VSUBS 0.008309f
C136 B.n99 VSUBS 0.008309f
C137 B.n100 VSUBS 0.008309f
C138 B.n101 VSUBS 0.008309f
C139 B.n102 VSUBS 0.008309f
C140 B.n103 VSUBS 0.008309f
C141 B.n104 VSUBS 0.008309f
C142 B.n105 VSUBS 0.008309f
C143 B.n106 VSUBS 0.008309f
C144 B.n107 VSUBS 0.008309f
C145 B.n108 VSUBS 0.008309f
C146 B.n109 VSUBS 0.008309f
C147 B.n110 VSUBS 0.008309f
C148 B.n111 VSUBS 0.008309f
C149 B.n112 VSUBS 0.008309f
C150 B.n113 VSUBS 0.008309f
C151 B.n114 VSUBS 0.008309f
C152 B.n115 VSUBS 0.008309f
C153 B.n116 VSUBS 0.008309f
C154 B.n117 VSUBS 0.008309f
C155 B.n118 VSUBS 0.008309f
C156 B.n119 VSUBS 0.008309f
C157 B.n120 VSUBS 0.008309f
C158 B.n121 VSUBS 0.008309f
C159 B.n122 VSUBS 0.008309f
C160 B.n123 VSUBS 0.008309f
C161 B.n124 VSUBS 0.008309f
C162 B.n125 VSUBS 0.008309f
C163 B.n126 VSUBS 0.008309f
C164 B.n127 VSUBS 0.020009f
C165 B.n128 VSUBS 0.021046f
C166 B.n129 VSUBS 0.021046f
C167 B.n130 VSUBS 0.008309f
C168 B.n131 VSUBS 0.008309f
C169 B.n132 VSUBS 0.008309f
C170 B.n133 VSUBS 0.008309f
C171 B.n134 VSUBS 0.008309f
C172 B.n135 VSUBS 0.008309f
C173 B.n136 VSUBS 0.008309f
C174 B.n137 VSUBS 0.008309f
C175 B.n138 VSUBS 0.008309f
C176 B.n139 VSUBS 0.008309f
C177 B.n140 VSUBS 0.008309f
C178 B.n141 VSUBS 0.008309f
C179 B.n142 VSUBS 0.008309f
C180 B.n143 VSUBS 0.008309f
C181 B.n144 VSUBS 0.008309f
C182 B.n145 VSUBS 0.008309f
C183 B.t2 VSUBS 0.062888f
C184 B.t1 VSUBS 0.067754f
C185 B.t0 VSUBS 0.079683f
C186 B.n146 VSUBS 0.068962f
C187 B.n147 VSUBS 0.063457f
C188 B.n148 VSUBS 0.019251f
C189 B.n149 VSUBS 0.00782f
C190 B.n150 VSUBS 0.008309f
C191 B.n151 VSUBS 0.008309f
C192 B.n152 VSUBS 0.008309f
C193 B.n153 VSUBS 0.008309f
C194 B.n154 VSUBS 0.008309f
C195 B.n155 VSUBS 0.008309f
C196 B.n156 VSUBS 0.008309f
C197 B.n157 VSUBS 0.008309f
C198 B.n158 VSUBS 0.008309f
C199 B.n159 VSUBS 0.008309f
C200 B.n160 VSUBS 0.008309f
C201 B.n161 VSUBS 0.008309f
C202 B.n162 VSUBS 0.008309f
C203 B.n163 VSUBS 0.008309f
C204 B.n164 VSUBS 0.008309f
C205 B.n165 VSUBS 0.004643f
C206 B.n166 VSUBS 0.019251f
C207 B.n167 VSUBS 0.00782f
C208 B.n168 VSUBS 0.008309f
C209 B.n169 VSUBS 0.008309f
C210 B.n170 VSUBS 0.008309f
C211 B.n171 VSUBS 0.008309f
C212 B.n172 VSUBS 0.008309f
C213 B.n173 VSUBS 0.008309f
C214 B.n174 VSUBS 0.008309f
C215 B.n175 VSUBS 0.008309f
C216 B.n176 VSUBS 0.008309f
C217 B.n177 VSUBS 0.008309f
C218 B.n178 VSUBS 0.008309f
C219 B.n179 VSUBS 0.008309f
C220 B.n180 VSUBS 0.008309f
C221 B.n181 VSUBS 0.008309f
C222 B.n182 VSUBS 0.008309f
C223 B.n183 VSUBS 0.008309f
C224 B.n184 VSUBS 0.008309f
C225 B.n185 VSUBS 0.020142f
C226 B.n186 VSUBS 0.020914f
C227 B.n187 VSUBS 0.020009f
C228 B.n188 VSUBS 0.008309f
C229 B.n189 VSUBS 0.008309f
C230 B.n190 VSUBS 0.008309f
C231 B.n191 VSUBS 0.008309f
C232 B.n192 VSUBS 0.008309f
C233 B.n193 VSUBS 0.008309f
C234 B.n194 VSUBS 0.008309f
C235 B.n195 VSUBS 0.008309f
C236 B.n196 VSUBS 0.008309f
C237 B.n197 VSUBS 0.008309f
C238 B.n198 VSUBS 0.008309f
C239 B.n199 VSUBS 0.008309f
C240 B.n200 VSUBS 0.008309f
C241 B.n201 VSUBS 0.008309f
C242 B.n202 VSUBS 0.008309f
C243 B.n203 VSUBS 0.008309f
C244 B.n204 VSUBS 0.008309f
C245 B.n205 VSUBS 0.008309f
C246 B.n206 VSUBS 0.008309f
C247 B.n207 VSUBS 0.008309f
C248 B.n208 VSUBS 0.008309f
C249 B.n209 VSUBS 0.008309f
C250 B.n210 VSUBS 0.008309f
C251 B.n211 VSUBS 0.008309f
C252 B.n212 VSUBS 0.008309f
C253 B.n213 VSUBS 0.008309f
C254 B.n214 VSUBS 0.008309f
C255 B.n215 VSUBS 0.008309f
C256 B.n216 VSUBS 0.008309f
C257 B.n217 VSUBS 0.008309f
C258 B.n218 VSUBS 0.008309f
C259 B.n219 VSUBS 0.008309f
C260 B.n220 VSUBS 0.008309f
C261 B.n221 VSUBS 0.008309f
C262 B.n222 VSUBS 0.008309f
C263 B.n223 VSUBS 0.008309f
C264 B.n224 VSUBS 0.008309f
C265 B.n225 VSUBS 0.008309f
C266 B.n226 VSUBS 0.008309f
C267 B.n227 VSUBS 0.008309f
C268 B.n228 VSUBS 0.008309f
C269 B.n229 VSUBS 0.008309f
C270 B.n230 VSUBS 0.008309f
C271 B.n231 VSUBS 0.008309f
C272 B.n232 VSUBS 0.008309f
C273 B.n233 VSUBS 0.008309f
C274 B.n234 VSUBS 0.008309f
C275 B.n235 VSUBS 0.008309f
C276 B.n236 VSUBS 0.008309f
C277 B.n237 VSUBS 0.008309f
C278 B.n238 VSUBS 0.008309f
C279 B.n239 VSUBS 0.008309f
C280 B.n240 VSUBS 0.008309f
C281 B.n241 VSUBS 0.008309f
C282 B.n242 VSUBS 0.008309f
C283 B.n243 VSUBS 0.008309f
C284 B.n244 VSUBS 0.008309f
C285 B.n245 VSUBS 0.008309f
C286 B.n246 VSUBS 0.008309f
C287 B.n247 VSUBS 0.008309f
C288 B.n248 VSUBS 0.008309f
C289 B.n249 VSUBS 0.008309f
C290 B.n250 VSUBS 0.008309f
C291 B.n251 VSUBS 0.008309f
C292 B.n252 VSUBS 0.008309f
C293 B.n253 VSUBS 0.008309f
C294 B.n254 VSUBS 0.008309f
C295 B.n255 VSUBS 0.008309f
C296 B.n256 VSUBS 0.008309f
C297 B.n257 VSUBS 0.008309f
C298 B.n258 VSUBS 0.008309f
C299 B.n259 VSUBS 0.008309f
C300 B.n260 VSUBS 0.020009f
C301 B.n261 VSUBS 0.021046f
C302 B.n262 VSUBS 0.021046f
C303 B.n263 VSUBS 0.008309f
C304 B.n264 VSUBS 0.008309f
C305 B.n265 VSUBS 0.008309f
C306 B.n266 VSUBS 0.008309f
C307 B.n267 VSUBS 0.008309f
C308 B.n268 VSUBS 0.008309f
C309 B.n269 VSUBS 0.008309f
C310 B.n270 VSUBS 0.008309f
C311 B.n271 VSUBS 0.008309f
C312 B.n272 VSUBS 0.008309f
C313 B.n273 VSUBS 0.008309f
C314 B.n274 VSUBS 0.008309f
C315 B.n275 VSUBS 0.008309f
C316 B.n276 VSUBS 0.008309f
C317 B.n277 VSUBS 0.008309f
C318 B.n278 VSUBS 0.008309f
C319 B.n279 VSUBS 0.008309f
C320 B.n280 VSUBS 0.00782f
C321 B.n281 VSUBS 0.019251f
C322 B.n282 VSUBS 0.004643f
C323 B.n283 VSUBS 0.008309f
C324 B.n284 VSUBS 0.008309f
C325 B.n285 VSUBS 0.008309f
C326 B.n286 VSUBS 0.008309f
C327 B.n287 VSUBS 0.008309f
C328 B.n288 VSUBS 0.008309f
C329 B.n289 VSUBS 0.008309f
C330 B.n290 VSUBS 0.008309f
C331 B.n291 VSUBS 0.008309f
C332 B.n292 VSUBS 0.008309f
C333 B.n293 VSUBS 0.008309f
C334 B.n294 VSUBS 0.008309f
C335 B.n295 VSUBS 0.004643f
C336 B.n296 VSUBS 0.008309f
C337 B.n297 VSUBS 0.008309f
C338 B.n298 VSUBS 0.008309f
C339 B.n299 VSUBS 0.008309f
C340 B.n300 VSUBS 0.008309f
C341 B.n301 VSUBS 0.008309f
C342 B.n302 VSUBS 0.008309f
C343 B.n303 VSUBS 0.008309f
C344 B.n304 VSUBS 0.008309f
C345 B.n305 VSUBS 0.008309f
C346 B.n306 VSUBS 0.008309f
C347 B.n307 VSUBS 0.008309f
C348 B.n308 VSUBS 0.008309f
C349 B.n309 VSUBS 0.008309f
C350 B.n310 VSUBS 0.008309f
C351 B.n311 VSUBS 0.008309f
C352 B.n312 VSUBS 0.008309f
C353 B.n313 VSUBS 0.008309f
C354 B.n314 VSUBS 0.008309f
C355 B.n315 VSUBS 0.021046f
C356 B.n316 VSUBS 0.020009f
C357 B.n317 VSUBS 0.020009f
C358 B.n318 VSUBS 0.008309f
C359 B.n319 VSUBS 0.008309f
C360 B.n320 VSUBS 0.008309f
C361 B.n321 VSUBS 0.008309f
C362 B.n322 VSUBS 0.008309f
C363 B.n323 VSUBS 0.008309f
C364 B.n324 VSUBS 0.008309f
C365 B.n325 VSUBS 0.008309f
C366 B.n326 VSUBS 0.008309f
C367 B.n327 VSUBS 0.008309f
C368 B.n328 VSUBS 0.008309f
C369 B.n329 VSUBS 0.008309f
C370 B.n330 VSUBS 0.008309f
C371 B.n331 VSUBS 0.008309f
C372 B.n332 VSUBS 0.008309f
C373 B.n333 VSUBS 0.008309f
C374 B.n334 VSUBS 0.008309f
C375 B.n335 VSUBS 0.008309f
C376 B.n336 VSUBS 0.008309f
C377 B.n337 VSUBS 0.008309f
C378 B.n338 VSUBS 0.008309f
C379 B.n339 VSUBS 0.008309f
C380 B.n340 VSUBS 0.008309f
C381 B.n341 VSUBS 0.008309f
C382 B.n342 VSUBS 0.008309f
C383 B.n343 VSUBS 0.008309f
C384 B.n344 VSUBS 0.008309f
C385 B.n345 VSUBS 0.008309f
C386 B.n346 VSUBS 0.008309f
C387 B.n347 VSUBS 0.008309f
C388 B.n348 VSUBS 0.008309f
C389 B.n349 VSUBS 0.008309f
C390 B.n350 VSUBS 0.008309f
C391 B.n351 VSUBS 0.010843f
C392 B.n352 VSUBS 0.01155f
C393 B.n353 VSUBS 0.022968f
C394 VDD2.t1 VSUBS 0.244886f
C395 VDD2.t8 VSUBS 0.035968f
C396 VDD2.t7 VSUBS 0.035968f
C397 VDD2.n0 VSUBS 0.162034f
C398 VDD2.n1 VSUBS 0.593549f
C399 VDD2.t3 VSUBS 0.035968f
C400 VDD2.t0 VSUBS 0.035968f
C401 VDD2.n2 VSUBS 0.163065f
C402 VDD2.n3 VSUBS 1.06537f
C403 VDD2.t4 VSUBS 0.243568f
C404 VDD2.n4 VSUBS 1.24926f
C405 VDD2.t6 VSUBS 0.035968f
C406 VDD2.t9 VSUBS 0.035968f
C407 VDD2.n5 VSUBS 0.162034f
C408 VDD2.n6 VSUBS 0.295355f
C409 VDD2.t2 VSUBS 0.035968f
C410 VDD2.t5 VSUBS 0.035968f
C411 VDD2.n7 VSUBS 0.163057f
C412 VN.n0 VSUBS 0.04901f
C413 VN.t2 VSUBS 0.21644f
C414 VN.n1 VSUBS 0.152666f
C415 VN.t8 VSUBS 0.236844f
C416 VN.t1 VSUBS 0.21644f
C417 VN.n2 VSUBS 0.152437f
C418 VN.n3 VSUBS 0.122829f
C419 VN.n4 VSUBS 0.238384f
C420 VN.n5 VSUBS 0.065398f
C421 VN.t6 VSUBS 0.21644f
C422 VN.n6 VSUBS 0.141695f
C423 VN.n7 VSUBS 0.011121f
C424 VN.t9 VSUBS 0.21644f
C425 VN.n8 VSUBS 0.141393f
C426 VN.n9 VSUBS 0.037981f
C427 VN.n10 VSUBS 0.04901f
C428 VN.t0 VSUBS 0.21644f
C429 VN.n11 VSUBS 0.152666f
C430 VN.t3 VSUBS 0.21644f
C431 VN.t4 VSUBS 0.236844f
C432 VN.t7 VSUBS 0.21644f
C433 VN.n12 VSUBS 0.152437f
C434 VN.n13 VSUBS 0.122829f
C435 VN.n14 VSUBS 0.238384f
C436 VN.n15 VSUBS 0.065398f
C437 VN.n16 VSUBS 0.141695f
C438 VN.n17 VSUBS 0.011121f
C439 VN.t5 VSUBS 0.21644f
C440 VN.n18 VSUBS 0.141393f
C441 VN.n19 VSUBS 1.49544f
C442 VDD1.t1 VSUBS 0.236632f
C443 VDD1.t8 VSUBS 0.034755f
C444 VDD1.t4 VSUBS 0.034755f
C445 VDD1.n0 VSUBS 0.156573f
C446 VDD1.n1 VSUBS 0.577407f
C447 VDD1.t7 VSUBS 0.236632f
C448 VDD1.t3 VSUBS 0.034755f
C449 VDD1.t5 VSUBS 0.034755f
C450 VDD1.n2 VSUBS 0.156572f
C451 VDD1.n3 VSUBS 0.573541f
C452 VDD1.t6 VSUBS 0.034755f
C453 VDD1.t0 VSUBS 0.034755f
C454 VDD1.n4 VSUBS 0.157568f
C455 VDD1.n5 VSUBS 1.08187f
C456 VDD1.t2 VSUBS 0.034755f
C457 VDD1.t9 VSUBS 0.034755f
C458 VDD1.n6 VSUBS 0.156573f
C459 VDD1.n7 VSUBS 1.24014f
C460 VTAIL.t19 VSUBS 0.043335f
C461 VTAIL.t5 VSUBS 0.043335f
C462 VTAIL.n0 VSUBS 0.166047f
C463 VTAIL.n1 VSUBS 0.388609f
C464 VTAIL.t14 VSUBS 0.26468f
C465 VTAIL.n2 VSUBS 0.418929f
C466 VTAIL.t12 VSUBS 0.043335f
C467 VTAIL.t8 VSUBS 0.043335f
C468 VTAIL.n3 VSUBS 0.166047f
C469 VTAIL.n4 VSUBS 0.394555f
C470 VTAIL.t15 VSUBS 0.043335f
C471 VTAIL.t9 VSUBS 0.043335f
C472 VTAIL.n5 VSUBS 0.166047f
C473 VTAIL.n6 VSUBS 0.921612f
C474 VTAIL.t16 VSUBS 0.043335f
C475 VTAIL.t4 VSUBS 0.043335f
C476 VTAIL.n7 VSUBS 0.166048f
C477 VTAIL.n8 VSUBS 0.921611f
C478 VTAIL.t0 VSUBS 0.043335f
C479 VTAIL.t18 VSUBS 0.043335f
C480 VTAIL.n9 VSUBS 0.166048f
C481 VTAIL.n10 VSUBS 0.394554f
C482 VTAIL.t3 VSUBS 0.264681f
C483 VTAIL.n11 VSUBS 0.418928f
C484 VTAIL.t6 VSUBS 0.043335f
C485 VTAIL.t7 VSUBS 0.043335f
C486 VTAIL.n12 VSUBS 0.166048f
C487 VTAIL.n13 VSUBS 0.399374f
C488 VTAIL.t10 VSUBS 0.043335f
C489 VTAIL.t13 VSUBS 0.043335f
C490 VTAIL.n14 VSUBS 0.166048f
C491 VTAIL.n15 VSUBS 0.394554f
C492 VTAIL.t11 VSUBS 0.264681f
C493 VTAIL.n16 VSUBS 0.880747f
C494 VTAIL.t2 VSUBS 0.26468f
C495 VTAIL.n17 VSUBS 0.880748f
C496 VTAIL.t1 VSUBS 0.043335f
C497 VTAIL.t17 VSUBS 0.043335f
C498 VTAIL.n18 VSUBS 0.166047f
C499 VTAIL.n19 VSUBS 0.344903f
C500 VP.n0 VSUBS 0.050808f
C501 VP.t4 VSUBS 0.224379f
C502 VP.n1 VSUBS 0.158265f
C503 VP.n2 VSUBS 0.050808f
C504 VP.n3 VSUBS 0.050808f
C505 VP.t0 VSUBS 0.224379f
C506 VP.t7 VSUBS 0.224379f
C507 VP.n4 VSUBS 0.067797f
C508 VP.t5 VSUBS 0.224379f
C509 VP.n5 VSUBS 0.247127f
C510 VP.t1 VSUBS 0.224379f
C511 VP.t8 VSUBS 0.245531f
C512 VP.n6 VSUBS 0.127334f
C513 VP.n7 VSUBS 0.158029f
C514 VP.n8 VSUBS 0.158265f
C515 VP.n9 VSUBS 0.146892f
C516 VP.n10 VSUBS 0.011529f
C517 VP.n11 VSUBS 0.146579f
C518 VP.n12 VSUBS 1.51652f
C519 VP.n13 VSUBS 1.56866f
C520 VP.t2 VSUBS 0.224379f
C521 VP.n14 VSUBS 0.146579f
C522 VP.n15 VSUBS 0.011529f
C523 VP.t6 VSUBS 0.224379f
C524 VP.n16 VSUBS 0.146892f
C525 VP.n17 VSUBS 0.067797f
C526 VP.n18 VSUBS 0.067638f
C527 VP.n19 VSUBS 0.067797f
C528 VP.t3 VSUBS 0.224379f
C529 VP.n20 VSUBS 0.146892f
C530 VP.n21 VSUBS 0.011529f
C531 VP.t9 VSUBS 0.224379f
C532 VP.n22 VSUBS 0.146579f
C533 VP.n23 VSUBS 0.039374f
.ends

