* NGSPICE file created from diff_pair_sample_1645.ext - technology: sky130A

.subckt diff_pair_sample_1645 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.47
X1 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.47
X2 VDD2.t2 VN.t1 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.47
X3 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.47
X4 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.47
X5 VDD1.t1 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.47
X6 VDD1.t0 VP.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.47
X7 VDD2.t1 VN.t2 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3365 pd=8.43 as=3.159 ps=16.98 w=8.1 l=0.47
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.47
X9 VTAIL.t3 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=1.3365 ps=8.43 w=8.1 l=0.47
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.47
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.159 pd=16.98 as=0 ps=0 w=8.1 l=0.47
R0 VN.n0 VN.t3 519.904
R1 VN.n1 VN.t2 519.904
R2 VN.n0 VN.t1 519.879
R3 VN.n1 VN.t0 519.879
R4 VN VN.n1 107.368
R5 VN VN.n0 70.265
R6 VDD2.n2 VDD2.n0 96.106
R7 VDD2.n2 VDD2.n1 63.3397
R8 VDD2.n1 VDD2.t3 2.44494
R9 VDD2.n1 VDD2.t1 2.44494
R10 VDD2.n0 VDD2.t0 2.44494
R11 VDD2.n0 VDD2.t2 2.44494
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n346 VTAIL.n308 289.615
R14 VTAIL.n38 VTAIL.n0 289.615
R15 VTAIL.n82 VTAIL.n44 289.615
R16 VTAIL.n126 VTAIL.n88 289.615
R17 VTAIL.n302 VTAIL.n264 289.615
R18 VTAIL.n258 VTAIL.n220 289.615
R19 VTAIL.n214 VTAIL.n176 289.615
R20 VTAIL.n170 VTAIL.n132 289.615
R21 VTAIL.n323 VTAIL.n322 185
R22 VTAIL.n320 VTAIL.n319 185
R23 VTAIL.n329 VTAIL.n328 185
R24 VTAIL.n331 VTAIL.n330 185
R25 VTAIL.n316 VTAIL.n315 185
R26 VTAIL.n337 VTAIL.n336 185
R27 VTAIL.n339 VTAIL.n338 185
R28 VTAIL.n312 VTAIL.n311 185
R29 VTAIL.n345 VTAIL.n344 185
R30 VTAIL.n347 VTAIL.n346 185
R31 VTAIL.n15 VTAIL.n14 185
R32 VTAIL.n12 VTAIL.n11 185
R33 VTAIL.n21 VTAIL.n20 185
R34 VTAIL.n23 VTAIL.n22 185
R35 VTAIL.n8 VTAIL.n7 185
R36 VTAIL.n29 VTAIL.n28 185
R37 VTAIL.n31 VTAIL.n30 185
R38 VTAIL.n4 VTAIL.n3 185
R39 VTAIL.n37 VTAIL.n36 185
R40 VTAIL.n39 VTAIL.n38 185
R41 VTAIL.n59 VTAIL.n58 185
R42 VTAIL.n56 VTAIL.n55 185
R43 VTAIL.n65 VTAIL.n64 185
R44 VTAIL.n67 VTAIL.n66 185
R45 VTAIL.n52 VTAIL.n51 185
R46 VTAIL.n73 VTAIL.n72 185
R47 VTAIL.n75 VTAIL.n74 185
R48 VTAIL.n48 VTAIL.n47 185
R49 VTAIL.n81 VTAIL.n80 185
R50 VTAIL.n83 VTAIL.n82 185
R51 VTAIL.n103 VTAIL.n102 185
R52 VTAIL.n100 VTAIL.n99 185
R53 VTAIL.n109 VTAIL.n108 185
R54 VTAIL.n111 VTAIL.n110 185
R55 VTAIL.n96 VTAIL.n95 185
R56 VTAIL.n117 VTAIL.n116 185
R57 VTAIL.n119 VTAIL.n118 185
R58 VTAIL.n92 VTAIL.n91 185
R59 VTAIL.n125 VTAIL.n124 185
R60 VTAIL.n127 VTAIL.n126 185
R61 VTAIL.n303 VTAIL.n302 185
R62 VTAIL.n301 VTAIL.n300 185
R63 VTAIL.n268 VTAIL.n267 185
R64 VTAIL.n295 VTAIL.n294 185
R65 VTAIL.n293 VTAIL.n292 185
R66 VTAIL.n272 VTAIL.n271 185
R67 VTAIL.n287 VTAIL.n286 185
R68 VTAIL.n285 VTAIL.n284 185
R69 VTAIL.n276 VTAIL.n275 185
R70 VTAIL.n279 VTAIL.n278 185
R71 VTAIL.n259 VTAIL.n258 185
R72 VTAIL.n257 VTAIL.n256 185
R73 VTAIL.n224 VTAIL.n223 185
R74 VTAIL.n251 VTAIL.n250 185
R75 VTAIL.n249 VTAIL.n248 185
R76 VTAIL.n228 VTAIL.n227 185
R77 VTAIL.n243 VTAIL.n242 185
R78 VTAIL.n241 VTAIL.n240 185
R79 VTAIL.n232 VTAIL.n231 185
R80 VTAIL.n235 VTAIL.n234 185
R81 VTAIL.n215 VTAIL.n214 185
R82 VTAIL.n213 VTAIL.n212 185
R83 VTAIL.n180 VTAIL.n179 185
R84 VTAIL.n207 VTAIL.n206 185
R85 VTAIL.n205 VTAIL.n204 185
R86 VTAIL.n184 VTAIL.n183 185
R87 VTAIL.n199 VTAIL.n198 185
R88 VTAIL.n197 VTAIL.n196 185
R89 VTAIL.n188 VTAIL.n187 185
R90 VTAIL.n191 VTAIL.n190 185
R91 VTAIL.n171 VTAIL.n170 185
R92 VTAIL.n169 VTAIL.n168 185
R93 VTAIL.n136 VTAIL.n135 185
R94 VTAIL.n163 VTAIL.n162 185
R95 VTAIL.n161 VTAIL.n160 185
R96 VTAIL.n140 VTAIL.n139 185
R97 VTAIL.n155 VTAIL.n154 185
R98 VTAIL.n153 VTAIL.n152 185
R99 VTAIL.n144 VTAIL.n143 185
R100 VTAIL.n147 VTAIL.n146 185
R101 VTAIL.t5 VTAIL.n321 147.659
R102 VTAIL.t3 VTAIL.n13 147.659
R103 VTAIL.t7 VTAIL.n57 147.659
R104 VTAIL.t2 VTAIL.n101 147.659
R105 VTAIL.t0 VTAIL.n277 147.659
R106 VTAIL.t1 VTAIL.n233 147.659
R107 VTAIL.t4 VTAIL.n189 147.659
R108 VTAIL.t6 VTAIL.n145 147.659
R109 VTAIL.n322 VTAIL.n319 104.615
R110 VTAIL.n329 VTAIL.n319 104.615
R111 VTAIL.n330 VTAIL.n329 104.615
R112 VTAIL.n330 VTAIL.n315 104.615
R113 VTAIL.n337 VTAIL.n315 104.615
R114 VTAIL.n338 VTAIL.n337 104.615
R115 VTAIL.n338 VTAIL.n311 104.615
R116 VTAIL.n345 VTAIL.n311 104.615
R117 VTAIL.n346 VTAIL.n345 104.615
R118 VTAIL.n14 VTAIL.n11 104.615
R119 VTAIL.n21 VTAIL.n11 104.615
R120 VTAIL.n22 VTAIL.n21 104.615
R121 VTAIL.n22 VTAIL.n7 104.615
R122 VTAIL.n29 VTAIL.n7 104.615
R123 VTAIL.n30 VTAIL.n29 104.615
R124 VTAIL.n30 VTAIL.n3 104.615
R125 VTAIL.n37 VTAIL.n3 104.615
R126 VTAIL.n38 VTAIL.n37 104.615
R127 VTAIL.n58 VTAIL.n55 104.615
R128 VTAIL.n65 VTAIL.n55 104.615
R129 VTAIL.n66 VTAIL.n65 104.615
R130 VTAIL.n66 VTAIL.n51 104.615
R131 VTAIL.n73 VTAIL.n51 104.615
R132 VTAIL.n74 VTAIL.n73 104.615
R133 VTAIL.n74 VTAIL.n47 104.615
R134 VTAIL.n81 VTAIL.n47 104.615
R135 VTAIL.n82 VTAIL.n81 104.615
R136 VTAIL.n102 VTAIL.n99 104.615
R137 VTAIL.n109 VTAIL.n99 104.615
R138 VTAIL.n110 VTAIL.n109 104.615
R139 VTAIL.n110 VTAIL.n95 104.615
R140 VTAIL.n117 VTAIL.n95 104.615
R141 VTAIL.n118 VTAIL.n117 104.615
R142 VTAIL.n118 VTAIL.n91 104.615
R143 VTAIL.n125 VTAIL.n91 104.615
R144 VTAIL.n126 VTAIL.n125 104.615
R145 VTAIL.n302 VTAIL.n301 104.615
R146 VTAIL.n301 VTAIL.n267 104.615
R147 VTAIL.n294 VTAIL.n267 104.615
R148 VTAIL.n294 VTAIL.n293 104.615
R149 VTAIL.n293 VTAIL.n271 104.615
R150 VTAIL.n286 VTAIL.n271 104.615
R151 VTAIL.n286 VTAIL.n285 104.615
R152 VTAIL.n285 VTAIL.n275 104.615
R153 VTAIL.n278 VTAIL.n275 104.615
R154 VTAIL.n258 VTAIL.n257 104.615
R155 VTAIL.n257 VTAIL.n223 104.615
R156 VTAIL.n250 VTAIL.n223 104.615
R157 VTAIL.n250 VTAIL.n249 104.615
R158 VTAIL.n249 VTAIL.n227 104.615
R159 VTAIL.n242 VTAIL.n227 104.615
R160 VTAIL.n242 VTAIL.n241 104.615
R161 VTAIL.n241 VTAIL.n231 104.615
R162 VTAIL.n234 VTAIL.n231 104.615
R163 VTAIL.n214 VTAIL.n213 104.615
R164 VTAIL.n213 VTAIL.n179 104.615
R165 VTAIL.n206 VTAIL.n179 104.615
R166 VTAIL.n206 VTAIL.n205 104.615
R167 VTAIL.n205 VTAIL.n183 104.615
R168 VTAIL.n198 VTAIL.n183 104.615
R169 VTAIL.n198 VTAIL.n197 104.615
R170 VTAIL.n197 VTAIL.n187 104.615
R171 VTAIL.n190 VTAIL.n187 104.615
R172 VTAIL.n170 VTAIL.n169 104.615
R173 VTAIL.n169 VTAIL.n135 104.615
R174 VTAIL.n162 VTAIL.n135 104.615
R175 VTAIL.n162 VTAIL.n161 104.615
R176 VTAIL.n161 VTAIL.n139 104.615
R177 VTAIL.n154 VTAIL.n139 104.615
R178 VTAIL.n154 VTAIL.n153 104.615
R179 VTAIL.n153 VTAIL.n143 104.615
R180 VTAIL.n146 VTAIL.n143 104.615
R181 VTAIL.n322 VTAIL.t5 52.3082
R182 VTAIL.n14 VTAIL.t3 52.3082
R183 VTAIL.n58 VTAIL.t7 52.3082
R184 VTAIL.n102 VTAIL.t2 52.3082
R185 VTAIL.n278 VTAIL.t0 52.3082
R186 VTAIL.n234 VTAIL.t1 52.3082
R187 VTAIL.n190 VTAIL.t4 52.3082
R188 VTAIL.n146 VTAIL.t6 52.3082
R189 VTAIL.n351 VTAIL.n350 31.0217
R190 VTAIL.n43 VTAIL.n42 31.0217
R191 VTAIL.n87 VTAIL.n86 31.0217
R192 VTAIL.n131 VTAIL.n130 31.0217
R193 VTAIL.n307 VTAIL.n306 31.0217
R194 VTAIL.n263 VTAIL.n262 31.0217
R195 VTAIL.n219 VTAIL.n218 31.0217
R196 VTAIL.n175 VTAIL.n174 31.0217
R197 VTAIL.n351 VTAIL.n307 20.0393
R198 VTAIL.n175 VTAIL.n131 20.0393
R199 VTAIL.n323 VTAIL.n321 15.6677
R200 VTAIL.n15 VTAIL.n13 15.6677
R201 VTAIL.n59 VTAIL.n57 15.6677
R202 VTAIL.n103 VTAIL.n101 15.6677
R203 VTAIL.n279 VTAIL.n277 15.6677
R204 VTAIL.n235 VTAIL.n233 15.6677
R205 VTAIL.n191 VTAIL.n189 15.6677
R206 VTAIL.n147 VTAIL.n145 15.6677
R207 VTAIL.n324 VTAIL.n320 12.8005
R208 VTAIL.n16 VTAIL.n12 12.8005
R209 VTAIL.n60 VTAIL.n56 12.8005
R210 VTAIL.n104 VTAIL.n100 12.8005
R211 VTAIL.n280 VTAIL.n276 12.8005
R212 VTAIL.n236 VTAIL.n232 12.8005
R213 VTAIL.n192 VTAIL.n188 12.8005
R214 VTAIL.n148 VTAIL.n144 12.8005
R215 VTAIL.n328 VTAIL.n327 12.0247
R216 VTAIL.n20 VTAIL.n19 12.0247
R217 VTAIL.n64 VTAIL.n63 12.0247
R218 VTAIL.n108 VTAIL.n107 12.0247
R219 VTAIL.n284 VTAIL.n283 12.0247
R220 VTAIL.n240 VTAIL.n239 12.0247
R221 VTAIL.n196 VTAIL.n195 12.0247
R222 VTAIL.n152 VTAIL.n151 12.0247
R223 VTAIL.n331 VTAIL.n318 11.249
R224 VTAIL.n23 VTAIL.n10 11.249
R225 VTAIL.n67 VTAIL.n54 11.249
R226 VTAIL.n111 VTAIL.n98 11.249
R227 VTAIL.n287 VTAIL.n274 11.249
R228 VTAIL.n243 VTAIL.n230 11.249
R229 VTAIL.n199 VTAIL.n186 11.249
R230 VTAIL.n155 VTAIL.n142 11.249
R231 VTAIL.n332 VTAIL.n316 10.4732
R232 VTAIL.n24 VTAIL.n8 10.4732
R233 VTAIL.n68 VTAIL.n52 10.4732
R234 VTAIL.n112 VTAIL.n96 10.4732
R235 VTAIL.n288 VTAIL.n272 10.4732
R236 VTAIL.n244 VTAIL.n228 10.4732
R237 VTAIL.n200 VTAIL.n184 10.4732
R238 VTAIL.n156 VTAIL.n140 10.4732
R239 VTAIL.n336 VTAIL.n335 9.69747
R240 VTAIL.n28 VTAIL.n27 9.69747
R241 VTAIL.n72 VTAIL.n71 9.69747
R242 VTAIL.n116 VTAIL.n115 9.69747
R243 VTAIL.n292 VTAIL.n291 9.69747
R244 VTAIL.n248 VTAIL.n247 9.69747
R245 VTAIL.n204 VTAIL.n203 9.69747
R246 VTAIL.n160 VTAIL.n159 9.69747
R247 VTAIL.n350 VTAIL.n349 9.45567
R248 VTAIL.n42 VTAIL.n41 9.45567
R249 VTAIL.n86 VTAIL.n85 9.45567
R250 VTAIL.n130 VTAIL.n129 9.45567
R251 VTAIL.n306 VTAIL.n305 9.45567
R252 VTAIL.n262 VTAIL.n261 9.45567
R253 VTAIL.n218 VTAIL.n217 9.45567
R254 VTAIL.n174 VTAIL.n173 9.45567
R255 VTAIL.n310 VTAIL.n309 9.3005
R256 VTAIL.n349 VTAIL.n348 9.3005
R257 VTAIL.n341 VTAIL.n340 9.3005
R258 VTAIL.n314 VTAIL.n313 9.3005
R259 VTAIL.n335 VTAIL.n334 9.3005
R260 VTAIL.n333 VTAIL.n332 9.3005
R261 VTAIL.n318 VTAIL.n317 9.3005
R262 VTAIL.n327 VTAIL.n326 9.3005
R263 VTAIL.n325 VTAIL.n324 9.3005
R264 VTAIL.n343 VTAIL.n342 9.3005
R265 VTAIL.n2 VTAIL.n1 9.3005
R266 VTAIL.n41 VTAIL.n40 9.3005
R267 VTAIL.n33 VTAIL.n32 9.3005
R268 VTAIL.n6 VTAIL.n5 9.3005
R269 VTAIL.n27 VTAIL.n26 9.3005
R270 VTAIL.n25 VTAIL.n24 9.3005
R271 VTAIL.n10 VTAIL.n9 9.3005
R272 VTAIL.n19 VTAIL.n18 9.3005
R273 VTAIL.n17 VTAIL.n16 9.3005
R274 VTAIL.n35 VTAIL.n34 9.3005
R275 VTAIL.n46 VTAIL.n45 9.3005
R276 VTAIL.n85 VTAIL.n84 9.3005
R277 VTAIL.n77 VTAIL.n76 9.3005
R278 VTAIL.n50 VTAIL.n49 9.3005
R279 VTAIL.n71 VTAIL.n70 9.3005
R280 VTAIL.n69 VTAIL.n68 9.3005
R281 VTAIL.n54 VTAIL.n53 9.3005
R282 VTAIL.n63 VTAIL.n62 9.3005
R283 VTAIL.n61 VTAIL.n60 9.3005
R284 VTAIL.n79 VTAIL.n78 9.3005
R285 VTAIL.n90 VTAIL.n89 9.3005
R286 VTAIL.n129 VTAIL.n128 9.3005
R287 VTAIL.n121 VTAIL.n120 9.3005
R288 VTAIL.n94 VTAIL.n93 9.3005
R289 VTAIL.n115 VTAIL.n114 9.3005
R290 VTAIL.n113 VTAIL.n112 9.3005
R291 VTAIL.n98 VTAIL.n97 9.3005
R292 VTAIL.n107 VTAIL.n106 9.3005
R293 VTAIL.n105 VTAIL.n104 9.3005
R294 VTAIL.n123 VTAIL.n122 9.3005
R295 VTAIL.n266 VTAIL.n265 9.3005
R296 VTAIL.n299 VTAIL.n298 9.3005
R297 VTAIL.n297 VTAIL.n296 9.3005
R298 VTAIL.n270 VTAIL.n269 9.3005
R299 VTAIL.n291 VTAIL.n290 9.3005
R300 VTAIL.n289 VTAIL.n288 9.3005
R301 VTAIL.n274 VTAIL.n273 9.3005
R302 VTAIL.n283 VTAIL.n282 9.3005
R303 VTAIL.n281 VTAIL.n280 9.3005
R304 VTAIL.n305 VTAIL.n304 9.3005
R305 VTAIL.n261 VTAIL.n260 9.3005
R306 VTAIL.n222 VTAIL.n221 9.3005
R307 VTAIL.n255 VTAIL.n254 9.3005
R308 VTAIL.n253 VTAIL.n252 9.3005
R309 VTAIL.n226 VTAIL.n225 9.3005
R310 VTAIL.n247 VTAIL.n246 9.3005
R311 VTAIL.n245 VTAIL.n244 9.3005
R312 VTAIL.n230 VTAIL.n229 9.3005
R313 VTAIL.n239 VTAIL.n238 9.3005
R314 VTAIL.n237 VTAIL.n236 9.3005
R315 VTAIL.n217 VTAIL.n216 9.3005
R316 VTAIL.n178 VTAIL.n177 9.3005
R317 VTAIL.n211 VTAIL.n210 9.3005
R318 VTAIL.n209 VTAIL.n208 9.3005
R319 VTAIL.n182 VTAIL.n181 9.3005
R320 VTAIL.n203 VTAIL.n202 9.3005
R321 VTAIL.n201 VTAIL.n200 9.3005
R322 VTAIL.n186 VTAIL.n185 9.3005
R323 VTAIL.n195 VTAIL.n194 9.3005
R324 VTAIL.n193 VTAIL.n192 9.3005
R325 VTAIL.n173 VTAIL.n172 9.3005
R326 VTAIL.n134 VTAIL.n133 9.3005
R327 VTAIL.n167 VTAIL.n166 9.3005
R328 VTAIL.n165 VTAIL.n164 9.3005
R329 VTAIL.n138 VTAIL.n137 9.3005
R330 VTAIL.n159 VTAIL.n158 9.3005
R331 VTAIL.n157 VTAIL.n156 9.3005
R332 VTAIL.n142 VTAIL.n141 9.3005
R333 VTAIL.n151 VTAIL.n150 9.3005
R334 VTAIL.n149 VTAIL.n148 9.3005
R335 VTAIL.n339 VTAIL.n314 8.92171
R336 VTAIL.n31 VTAIL.n6 8.92171
R337 VTAIL.n75 VTAIL.n50 8.92171
R338 VTAIL.n119 VTAIL.n94 8.92171
R339 VTAIL.n295 VTAIL.n270 8.92171
R340 VTAIL.n251 VTAIL.n226 8.92171
R341 VTAIL.n207 VTAIL.n182 8.92171
R342 VTAIL.n163 VTAIL.n138 8.92171
R343 VTAIL.n340 VTAIL.n312 8.14595
R344 VTAIL.n350 VTAIL.n308 8.14595
R345 VTAIL.n32 VTAIL.n4 8.14595
R346 VTAIL.n42 VTAIL.n0 8.14595
R347 VTAIL.n76 VTAIL.n48 8.14595
R348 VTAIL.n86 VTAIL.n44 8.14595
R349 VTAIL.n120 VTAIL.n92 8.14595
R350 VTAIL.n130 VTAIL.n88 8.14595
R351 VTAIL.n306 VTAIL.n264 8.14595
R352 VTAIL.n296 VTAIL.n268 8.14595
R353 VTAIL.n262 VTAIL.n220 8.14595
R354 VTAIL.n252 VTAIL.n224 8.14595
R355 VTAIL.n218 VTAIL.n176 8.14595
R356 VTAIL.n208 VTAIL.n180 8.14595
R357 VTAIL.n174 VTAIL.n132 8.14595
R358 VTAIL.n164 VTAIL.n136 8.14595
R359 VTAIL.n344 VTAIL.n343 7.3702
R360 VTAIL.n348 VTAIL.n347 7.3702
R361 VTAIL.n36 VTAIL.n35 7.3702
R362 VTAIL.n40 VTAIL.n39 7.3702
R363 VTAIL.n80 VTAIL.n79 7.3702
R364 VTAIL.n84 VTAIL.n83 7.3702
R365 VTAIL.n124 VTAIL.n123 7.3702
R366 VTAIL.n128 VTAIL.n127 7.3702
R367 VTAIL.n304 VTAIL.n303 7.3702
R368 VTAIL.n300 VTAIL.n299 7.3702
R369 VTAIL.n260 VTAIL.n259 7.3702
R370 VTAIL.n256 VTAIL.n255 7.3702
R371 VTAIL.n216 VTAIL.n215 7.3702
R372 VTAIL.n212 VTAIL.n211 7.3702
R373 VTAIL.n172 VTAIL.n171 7.3702
R374 VTAIL.n168 VTAIL.n167 7.3702
R375 VTAIL.n344 VTAIL.n310 6.59444
R376 VTAIL.n347 VTAIL.n310 6.59444
R377 VTAIL.n36 VTAIL.n2 6.59444
R378 VTAIL.n39 VTAIL.n2 6.59444
R379 VTAIL.n80 VTAIL.n46 6.59444
R380 VTAIL.n83 VTAIL.n46 6.59444
R381 VTAIL.n124 VTAIL.n90 6.59444
R382 VTAIL.n127 VTAIL.n90 6.59444
R383 VTAIL.n303 VTAIL.n266 6.59444
R384 VTAIL.n300 VTAIL.n266 6.59444
R385 VTAIL.n259 VTAIL.n222 6.59444
R386 VTAIL.n256 VTAIL.n222 6.59444
R387 VTAIL.n215 VTAIL.n178 6.59444
R388 VTAIL.n212 VTAIL.n178 6.59444
R389 VTAIL.n171 VTAIL.n134 6.59444
R390 VTAIL.n168 VTAIL.n134 6.59444
R391 VTAIL.n343 VTAIL.n312 5.81868
R392 VTAIL.n348 VTAIL.n308 5.81868
R393 VTAIL.n35 VTAIL.n4 5.81868
R394 VTAIL.n40 VTAIL.n0 5.81868
R395 VTAIL.n79 VTAIL.n48 5.81868
R396 VTAIL.n84 VTAIL.n44 5.81868
R397 VTAIL.n123 VTAIL.n92 5.81868
R398 VTAIL.n128 VTAIL.n88 5.81868
R399 VTAIL.n304 VTAIL.n264 5.81868
R400 VTAIL.n299 VTAIL.n268 5.81868
R401 VTAIL.n260 VTAIL.n220 5.81868
R402 VTAIL.n255 VTAIL.n224 5.81868
R403 VTAIL.n216 VTAIL.n176 5.81868
R404 VTAIL.n211 VTAIL.n180 5.81868
R405 VTAIL.n172 VTAIL.n132 5.81868
R406 VTAIL.n167 VTAIL.n136 5.81868
R407 VTAIL.n340 VTAIL.n339 5.04292
R408 VTAIL.n32 VTAIL.n31 5.04292
R409 VTAIL.n76 VTAIL.n75 5.04292
R410 VTAIL.n120 VTAIL.n119 5.04292
R411 VTAIL.n296 VTAIL.n295 5.04292
R412 VTAIL.n252 VTAIL.n251 5.04292
R413 VTAIL.n208 VTAIL.n207 5.04292
R414 VTAIL.n164 VTAIL.n163 5.04292
R415 VTAIL.n325 VTAIL.n321 4.38564
R416 VTAIL.n17 VTAIL.n13 4.38564
R417 VTAIL.n61 VTAIL.n57 4.38564
R418 VTAIL.n105 VTAIL.n101 4.38564
R419 VTAIL.n237 VTAIL.n233 4.38564
R420 VTAIL.n193 VTAIL.n189 4.38564
R421 VTAIL.n149 VTAIL.n145 4.38564
R422 VTAIL.n281 VTAIL.n277 4.38564
R423 VTAIL.n336 VTAIL.n314 4.26717
R424 VTAIL.n28 VTAIL.n6 4.26717
R425 VTAIL.n72 VTAIL.n50 4.26717
R426 VTAIL.n116 VTAIL.n94 4.26717
R427 VTAIL.n292 VTAIL.n270 4.26717
R428 VTAIL.n248 VTAIL.n226 4.26717
R429 VTAIL.n204 VTAIL.n182 4.26717
R430 VTAIL.n160 VTAIL.n138 4.26717
R431 VTAIL.n335 VTAIL.n316 3.49141
R432 VTAIL.n27 VTAIL.n8 3.49141
R433 VTAIL.n71 VTAIL.n52 3.49141
R434 VTAIL.n115 VTAIL.n96 3.49141
R435 VTAIL.n291 VTAIL.n272 3.49141
R436 VTAIL.n247 VTAIL.n228 3.49141
R437 VTAIL.n203 VTAIL.n184 3.49141
R438 VTAIL.n159 VTAIL.n140 3.49141
R439 VTAIL.n332 VTAIL.n331 2.71565
R440 VTAIL.n24 VTAIL.n23 2.71565
R441 VTAIL.n68 VTAIL.n67 2.71565
R442 VTAIL.n112 VTAIL.n111 2.71565
R443 VTAIL.n288 VTAIL.n287 2.71565
R444 VTAIL.n244 VTAIL.n243 2.71565
R445 VTAIL.n200 VTAIL.n199 2.71565
R446 VTAIL.n156 VTAIL.n155 2.71565
R447 VTAIL.n328 VTAIL.n318 1.93989
R448 VTAIL.n20 VTAIL.n10 1.93989
R449 VTAIL.n64 VTAIL.n54 1.93989
R450 VTAIL.n108 VTAIL.n98 1.93989
R451 VTAIL.n284 VTAIL.n274 1.93989
R452 VTAIL.n240 VTAIL.n230 1.93989
R453 VTAIL.n196 VTAIL.n186 1.93989
R454 VTAIL.n152 VTAIL.n142 1.93989
R455 VTAIL.n327 VTAIL.n320 1.16414
R456 VTAIL.n19 VTAIL.n12 1.16414
R457 VTAIL.n63 VTAIL.n56 1.16414
R458 VTAIL.n107 VTAIL.n100 1.16414
R459 VTAIL.n283 VTAIL.n276 1.16414
R460 VTAIL.n239 VTAIL.n232 1.16414
R461 VTAIL.n195 VTAIL.n188 1.16414
R462 VTAIL.n151 VTAIL.n144 1.16414
R463 VTAIL.n219 VTAIL.n175 0.690155
R464 VTAIL.n307 VTAIL.n263 0.690155
R465 VTAIL.n131 VTAIL.n87 0.690155
R466 VTAIL.n263 VTAIL.n219 0.470328
R467 VTAIL.n87 VTAIL.n43 0.470328
R468 VTAIL VTAIL.n43 0.403517
R469 VTAIL.n324 VTAIL.n323 0.388379
R470 VTAIL.n16 VTAIL.n15 0.388379
R471 VTAIL.n60 VTAIL.n59 0.388379
R472 VTAIL.n104 VTAIL.n103 0.388379
R473 VTAIL.n280 VTAIL.n279 0.388379
R474 VTAIL.n236 VTAIL.n235 0.388379
R475 VTAIL.n192 VTAIL.n191 0.388379
R476 VTAIL.n148 VTAIL.n147 0.388379
R477 VTAIL VTAIL.n351 0.287138
R478 VTAIL.n326 VTAIL.n325 0.155672
R479 VTAIL.n326 VTAIL.n317 0.155672
R480 VTAIL.n333 VTAIL.n317 0.155672
R481 VTAIL.n334 VTAIL.n333 0.155672
R482 VTAIL.n334 VTAIL.n313 0.155672
R483 VTAIL.n341 VTAIL.n313 0.155672
R484 VTAIL.n342 VTAIL.n341 0.155672
R485 VTAIL.n342 VTAIL.n309 0.155672
R486 VTAIL.n349 VTAIL.n309 0.155672
R487 VTAIL.n18 VTAIL.n17 0.155672
R488 VTAIL.n18 VTAIL.n9 0.155672
R489 VTAIL.n25 VTAIL.n9 0.155672
R490 VTAIL.n26 VTAIL.n25 0.155672
R491 VTAIL.n26 VTAIL.n5 0.155672
R492 VTAIL.n33 VTAIL.n5 0.155672
R493 VTAIL.n34 VTAIL.n33 0.155672
R494 VTAIL.n34 VTAIL.n1 0.155672
R495 VTAIL.n41 VTAIL.n1 0.155672
R496 VTAIL.n62 VTAIL.n61 0.155672
R497 VTAIL.n62 VTAIL.n53 0.155672
R498 VTAIL.n69 VTAIL.n53 0.155672
R499 VTAIL.n70 VTAIL.n69 0.155672
R500 VTAIL.n70 VTAIL.n49 0.155672
R501 VTAIL.n77 VTAIL.n49 0.155672
R502 VTAIL.n78 VTAIL.n77 0.155672
R503 VTAIL.n78 VTAIL.n45 0.155672
R504 VTAIL.n85 VTAIL.n45 0.155672
R505 VTAIL.n106 VTAIL.n105 0.155672
R506 VTAIL.n106 VTAIL.n97 0.155672
R507 VTAIL.n113 VTAIL.n97 0.155672
R508 VTAIL.n114 VTAIL.n113 0.155672
R509 VTAIL.n114 VTAIL.n93 0.155672
R510 VTAIL.n121 VTAIL.n93 0.155672
R511 VTAIL.n122 VTAIL.n121 0.155672
R512 VTAIL.n122 VTAIL.n89 0.155672
R513 VTAIL.n129 VTAIL.n89 0.155672
R514 VTAIL.n305 VTAIL.n265 0.155672
R515 VTAIL.n298 VTAIL.n265 0.155672
R516 VTAIL.n298 VTAIL.n297 0.155672
R517 VTAIL.n297 VTAIL.n269 0.155672
R518 VTAIL.n290 VTAIL.n269 0.155672
R519 VTAIL.n290 VTAIL.n289 0.155672
R520 VTAIL.n289 VTAIL.n273 0.155672
R521 VTAIL.n282 VTAIL.n273 0.155672
R522 VTAIL.n282 VTAIL.n281 0.155672
R523 VTAIL.n261 VTAIL.n221 0.155672
R524 VTAIL.n254 VTAIL.n221 0.155672
R525 VTAIL.n254 VTAIL.n253 0.155672
R526 VTAIL.n253 VTAIL.n225 0.155672
R527 VTAIL.n246 VTAIL.n225 0.155672
R528 VTAIL.n246 VTAIL.n245 0.155672
R529 VTAIL.n245 VTAIL.n229 0.155672
R530 VTAIL.n238 VTAIL.n229 0.155672
R531 VTAIL.n238 VTAIL.n237 0.155672
R532 VTAIL.n217 VTAIL.n177 0.155672
R533 VTAIL.n210 VTAIL.n177 0.155672
R534 VTAIL.n210 VTAIL.n209 0.155672
R535 VTAIL.n209 VTAIL.n181 0.155672
R536 VTAIL.n202 VTAIL.n181 0.155672
R537 VTAIL.n202 VTAIL.n201 0.155672
R538 VTAIL.n201 VTAIL.n185 0.155672
R539 VTAIL.n194 VTAIL.n185 0.155672
R540 VTAIL.n194 VTAIL.n193 0.155672
R541 VTAIL.n173 VTAIL.n133 0.155672
R542 VTAIL.n166 VTAIL.n133 0.155672
R543 VTAIL.n166 VTAIL.n165 0.155672
R544 VTAIL.n165 VTAIL.n137 0.155672
R545 VTAIL.n158 VTAIL.n137 0.155672
R546 VTAIL.n158 VTAIL.n157 0.155672
R547 VTAIL.n157 VTAIL.n141 0.155672
R548 VTAIL.n150 VTAIL.n141 0.155672
R549 VTAIL.n150 VTAIL.n149 0.155672
R550 B.n272 B.t12 622.518
R551 B.n270 B.t8 622.518
R552 B.n71 B.t15 622.518
R553 B.n68 B.t4 622.518
R554 B.n480 B.n479 585
R555 B.n206 B.n66 585
R556 B.n205 B.n204 585
R557 B.n203 B.n202 585
R558 B.n201 B.n200 585
R559 B.n199 B.n198 585
R560 B.n197 B.n196 585
R561 B.n195 B.n194 585
R562 B.n193 B.n192 585
R563 B.n191 B.n190 585
R564 B.n189 B.n188 585
R565 B.n187 B.n186 585
R566 B.n185 B.n184 585
R567 B.n183 B.n182 585
R568 B.n181 B.n180 585
R569 B.n179 B.n178 585
R570 B.n177 B.n176 585
R571 B.n175 B.n174 585
R572 B.n173 B.n172 585
R573 B.n171 B.n170 585
R574 B.n169 B.n168 585
R575 B.n167 B.n166 585
R576 B.n165 B.n164 585
R577 B.n163 B.n162 585
R578 B.n161 B.n160 585
R579 B.n159 B.n158 585
R580 B.n157 B.n156 585
R581 B.n155 B.n154 585
R582 B.n153 B.n152 585
R583 B.n151 B.n150 585
R584 B.n149 B.n148 585
R585 B.n147 B.n146 585
R586 B.n145 B.n144 585
R587 B.n143 B.n142 585
R588 B.n141 B.n140 585
R589 B.n139 B.n138 585
R590 B.n137 B.n136 585
R591 B.n135 B.n134 585
R592 B.n133 B.n132 585
R593 B.n131 B.n130 585
R594 B.n129 B.n128 585
R595 B.n127 B.n126 585
R596 B.n125 B.n124 585
R597 B.n123 B.n122 585
R598 B.n121 B.n120 585
R599 B.n119 B.n118 585
R600 B.n117 B.n116 585
R601 B.n115 B.n114 585
R602 B.n113 B.n112 585
R603 B.n111 B.n110 585
R604 B.n109 B.n108 585
R605 B.n107 B.n106 585
R606 B.n105 B.n104 585
R607 B.n103 B.n102 585
R608 B.n101 B.n100 585
R609 B.n99 B.n98 585
R610 B.n97 B.n96 585
R611 B.n95 B.n94 585
R612 B.n93 B.n92 585
R613 B.n91 B.n90 585
R614 B.n89 B.n88 585
R615 B.n87 B.n86 585
R616 B.n85 B.n84 585
R617 B.n83 B.n82 585
R618 B.n81 B.n80 585
R619 B.n79 B.n78 585
R620 B.n77 B.n76 585
R621 B.n75 B.n74 585
R622 B.n32 B.n31 585
R623 B.n485 B.n484 585
R624 B.n478 B.n67 585
R625 B.n67 B.n29 585
R626 B.n477 B.n28 585
R627 B.n489 B.n28 585
R628 B.n476 B.n27 585
R629 B.n490 B.n27 585
R630 B.n475 B.n26 585
R631 B.n491 B.n26 585
R632 B.n474 B.n473 585
R633 B.n473 B.n25 585
R634 B.n472 B.n21 585
R635 B.n497 B.n21 585
R636 B.n471 B.n20 585
R637 B.n498 B.n20 585
R638 B.n470 B.n19 585
R639 B.n499 B.n19 585
R640 B.n469 B.n468 585
R641 B.n468 B.n15 585
R642 B.n467 B.n14 585
R643 B.n505 B.n14 585
R644 B.n466 B.n13 585
R645 B.n506 B.n13 585
R646 B.n465 B.n12 585
R647 B.n507 B.n12 585
R648 B.n464 B.n463 585
R649 B.n463 B.n11 585
R650 B.n462 B.n7 585
R651 B.n513 B.n7 585
R652 B.n461 B.n6 585
R653 B.n514 B.n6 585
R654 B.n460 B.n5 585
R655 B.n515 B.n5 585
R656 B.n459 B.n458 585
R657 B.n458 B.n4 585
R658 B.n457 B.n207 585
R659 B.n457 B.n456 585
R660 B.n446 B.n208 585
R661 B.n449 B.n208 585
R662 B.n448 B.n447 585
R663 B.n450 B.n448 585
R664 B.n445 B.n213 585
R665 B.n213 B.n212 585
R666 B.n444 B.n443 585
R667 B.n443 B.n442 585
R668 B.n215 B.n214 585
R669 B.n216 B.n215 585
R670 B.n435 B.n434 585
R671 B.n436 B.n435 585
R672 B.n433 B.n221 585
R673 B.n221 B.n220 585
R674 B.n432 B.n431 585
R675 B.n431 B.n430 585
R676 B.n223 B.n222 585
R677 B.n423 B.n223 585
R678 B.n422 B.n421 585
R679 B.n424 B.n422 585
R680 B.n420 B.n228 585
R681 B.n228 B.n227 585
R682 B.n419 B.n418 585
R683 B.n418 B.n417 585
R684 B.n230 B.n229 585
R685 B.n231 B.n230 585
R686 B.n413 B.n412 585
R687 B.n234 B.n233 585
R688 B.n409 B.n408 585
R689 B.n410 B.n409 585
R690 B.n407 B.n269 585
R691 B.n406 B.n405 585
R692 B.n404 B.n403 585
R693 B.n402 B.n401 585
R694 B.n400 B.n399 585
R695 B.n398 B.n397 585
R696 B.n396 B.n395 585
R697 B.n394 B.n393 585
R698 B.n392 B.n391 585
R699 B.n390 B.n389 585
R700 B.n388 B.n387 585
R701 B.n386 B.n385 585
R702 B.n384 B.n383 585
R703 B.n382 B.n381 585
R704 B.n380 B.n379 585
R705 B.n378 B.n377 585
R706 B.n376 B.n375 585
R707 B.n374 B.n373 585
R708 B.n372 B.n371 585
R709 B.n370 B.n369 585
R710 B.n368 B.n367 585
R711 B.n366 B.n365 585
R712 B.n364 B.n363 585
R713 B.n362 B.n361 585
R714 B.n360 B.n359 585
R715 B.n358 B.n357 585
R716 B.n356 B.n355 585
R717 B.n353 B.n352 585
R718 B.n351 B.n350 585
R719 B.n349 B.n348 585
R720 B.n347 B.n346 585
R721 B.n345 B.n344 585
R722 B.n343 B.n342 585
R723 B.n341 B.n340 585
R724 B.n339 B.n338 585
R725 B.n337 B.n336 585
R726 B.n335 B.n334 585
R727 B.n332 B.n331 585
R728 B.n330 B.n329 585
R729 B.n328 B.n327 585
R730 B.n326 B.n325 585
R731 B.n324 B.n323 585
R732 B.n322 B.n321 585
R733 B.n320 B.n319 585
R734 B.n318 B.n317 585
R735 B.n316 B.n315 585
R736 B.n314 B.n313 585
R737 B.n312 B.n311 585
R738 B.n310 B.n309 585
R739 B.n308 B.n307 585
R740 B.n306 B.n305 585
R741 B.n304 B.n303 585
R742 B.n302 B.n301 585
R743 B.n300 B.n299 585
R744 B.n298 B.n297 585
R745 B.n296 B.n295 585
R746 B.n294 B.n293 585
R747 B.n292 B.n291 585
R748 B.n290 B.n289 585
R749 B.n288 B.n287 585
R750 B.n286 B.n285 585
R751 B.n284 B.n283 585
R752 B.n282 B.n281 585
R753 B.n280 B.n279 585
R754 B.n278 B.n277 585
R755 B.n276 B.n275 585
R756 B.n274 B.n268 585
R757 B.n410 B.n268 585
R758 B.n414 B.n232 585
R759 B.n232 B.n231 585
R760 B.n416 B.n415 585
R761 B.n417 B.n416 585
R762 B.n226 B.n225 585
R763 B.n227 B.n226 585
R764 B.n426 B.n425 585
R765 B.n425 B.n424 585
R766 B.n427 B.n224 585
R767 B.n423 B.n224 585
R768 B.n429 B.n428 585
R769 B.n430 B.n429 585
R770 B.n219 B.n218 585
R771 B.n220 B.n219 585
R772 B.n438 B.n437 585
R773 B.n437 B.n436 585
R774 B.n439 B.n217 585
R775 B.n217 B.n216 585
R776 B.n441 B.n440 585
R777 B.n442 B.n441 585
R778 B.n211 B.n210 585
R779 B.n212 B.n211 585
R780 B.n452 B.n451 585
R781 B.n451 B.n450 585
R782 B.n453 B.n209 585
R783 B.n449 B.n209 585
R784 B.n455 B.n454 585
R785 B.n456 B.n455 585
R786 B.n2 B.n0 585
R787 B.n4 B.n2 585
R788 B.n3 B.n1 585
R789 B.n514 B.n3 585
R790 B.n512 B.n511 585
R791 B.n513 B.n512 585
R792 B.n510 B.n8 585
R793 B.n11 B.n8 585
R794 B.n509 B.n508 585
R795 B.n508 B.n507 585
R796 B.n10 B.n9 585
R797 B.n506 B.n10 585
R798 B.n504 B.n503 585
R799 B.n505 B.n504 585
R800 B.n502 B.n16 585
R801 B.n16 B.n15 585
R802 B.n501 B.n500 585
R803 B.n500 B.n499 585
R804 B.n18 B.n17 585
R805 B.n498 B.n18 585
R806 B.n496 B.n495 585
R807 B.n497 B.n496 585
R808 B.n494 B.n22 585
R809 B.n25 B.n22 585
R810 B.n493 B.n492 585
R811 B.n492 B.n491 585
R812 B.n24 B.n23 585
R813 B.n490 B.n24 585
R814 B.n488 B.n487 585
R815 B.n489 B.n488 585
R816 B.n486 B.n30 585
R817 B.n30 B.n29 585
R818 B.n517 B.n516 585
R819 B.n516 B.n515 585
R820 B.n412 B.n232 516.524
R821 B.n484 B.n30 516.524
R822 B.n268 B.n230 516.524
R823 B.n480 B.n67 516.524
R824 B.n482 B.n481 256.663
R825 B.n482 B.n65 256.663
R826 B.n482 B.n64 256.663
R827 B.n482 B.n63 256.663
R828 B.n482 B.n62 256.663
R829 B.n482 B.n61 256.663
R830 B.n482 B.n60 256.663
R831 B.n482 B.n59 256.663
R832 B.n482 B.n58 256.663
R833 B.n482 B.n57 256.663
R834 B.n482 B.n56 256.663
R835 B.n482 B.n55 256.663
R836 B.n482 B.n54 256.663
R837 B.n482 B.n53 256.663
R838 B.n482 B.n52 256.663
R839 B.n482 B.n51 256.663
R840 B.n482 B.n50 256.663
R841 B.n482 B.n49 256.663
R842 B.n482 B.n48 256.663
R843 B.n482 B.n47 256.663
R844 B.n482 B.n46 256.663
R845 B.n482 B.n45 256.663
R846 B.n482 B.n44 256.663
R847 B.n482 B.n43 256.663
R848 B.n482 B.n42 256.663
R849 B.n482 B.n41 256.663
R850 B.n482 B.n40 256.663
R851 B.n482 B.n39 256.663
R852 B.n482 B.n38 256.663
R853 B.n482 B.n37 256.663
R854 B.n482 B.n36 256.663
R855 B.n482 B.n35 256.663
R856 B.n482 B.n34 256.663
R857 B.n482 B.n33 256.663
R858 B.n483 B.n482 256.663
R859 B.n411 B.n410 256.663
R860 B.n410 B.n235 256.663
R861 B.n410 B.n236 256.663
R862 B.n410 B.n237 256.663
R863 B.n410 B.n238 256.663
R864 B.n410 B.n239 256.663
R865 B.n410 B.n240 256.663
R866 B.n410 B.n241 256.663
R867 B.n410 B.n242 256.663
R868 B.n410 B.n243 256.663
R869 B.n410 B.n244 256.663
R870 B.n410 B.n245 256.663
R871 B.n410 B.n246 256.663
R872 B.n410 B.n247 256.663
R873 B.n410 B.n248 256.663
R874 B.n410 B.n249 256.663
R875 B.n410 B.n250 256.663
R876 B.n410 B.n251 256.663
R877 B.n410 B.n252 256.663
R878 B.n410 B.n253 256.663
R879 B.n410 B.n254 256.663
R880 B.n410 B.n255 256.663
R881 B.n410 B.n256 256.663
R882 B.n410 B.n257 256.663
R883 B.n410 B.n258 256.663
R884 B.n410 B.n259 256.663
R885 B.n410 B.n260 256.663
R886 B.n410 B.n261 256.663
R887 B.n410 B.n262 256.663
R888 B.n410 B.n263 256.663
R889 B.n410 B.n264 256.663
R890 B.n410 B.n265 256.663
R891 B.n410 B.n266 256.663
R892 B.n410 B.n267 256.663
R893 B.n272 B.t14 230.745
R894 B.n68 B.t6 230.745
R895 B.n270 B.t11 230.745
R896 B.n71 B.t16 230.745
R897 B.n273 B.t13 215.231
R898 B.n69 B.t7 215.231
R899 B.n271 B.t10 215.231
R900 B.n72 B.t17 215.231
R901 B.n416 B.n232 163.367
R902 B.n416 B.n226 163.367
R903 B.n425 B.n226 163.367
R904 B.n425 B.n224 163.367
R905 B.n429 B.n224 163.367
R906 B.n429 B.n219 163.367
R907 B.n437 B.n219 163.367
R908 B.n437 B.n217 163.367
R909 B.n441 B.n217 163.367
R910 B.n441 B.n211 163.367
R911 B.n451 B.n211 163.367
R912 B.n451 B.n209 163.367
R913 B.n455 B.n209 163.367
R914 B.n455 B.n2 163.367
R915 B.n516 B.n2 163.367
R916 B.n516 B.n3 163.367
R917 B.n512 B.n3 163.367
R918 B.n512 B.n8 163.367
R919 B.n508 B.n8 163.367
R920 B.n508 B.n10 163.367
R921 B.n504 B.n10 163.367
R922 B.n504 B.n16 163.367
R923 B.n500 B.n16 163.367
R924 B.n500 B.n18 163.367
R925 B.n496 B.n18 163.367
R926 B.n496 B.n22 163.367
R927 B.n492 B.n22 163.367
R928 B.n492 B.n24 163.367
R929 B.n488 B.n24 163.367
R930 B.n488 B.n30 163.367
R931 B.n409 B.n234 163.367
R932 B.n409 B.n269 163.367
R933 B.n405 B.n404 163.367
R934 B.n401 B.n400 163.367
R935 B.n397 B.n396 163.367
R936 B.n393 B.n392 163.367
R937 B.n389 B.n388 163.367
R938 B.n385 B.n384 163.367
R939 B.n381 B.n380 163.367
R940 B.n377 B.n376 163.367
R941 B.n373 B.n372 163.367
R942 B.n369 B.n368 163.367
R943 B.n365 B.n364 163.367
R944 B.n361 B.n360 163.367
R945 B.n357 B.n356 163.367
R946 B.n352 B.n351 163.367
R947 B.n348 B.n347 163.367
R948 B.n344 B.n343 163.367
R949 B.n340 B.n339 163.367
R950 B.n336 B.n335 163.367
R951 B.n331 B.n330 163.367
R952 B.n327 B.n326 163.367
R953 B.n323 B.n322 163.367
R954 B.n319 B.n318 163.367
R955 B.n315 B.n314 163.367
R956 B.n311 B.n310 163.367
R957 B.n307 B.n306 163.367
R958 B.n303 B.n302 163.367
R959 B.n299 B.n298 163.367
R960 B.n295 B.n294 163.367
R961 B.n291 B.n290 163.367
R962 B.n287 B.n286 163.367
R963 B.n283 B.n282 163.367
R964 B.n279 B.n278 163.367
R965 B.n275 B.n268 163.367
R966 B.n418 B.n230 163.367
R967 B.n418 B.n228 163.367
R968 B.n422 B.n228 163.367
R969 B.n422 B.n223 163.367
R970 B.n431 B.n223 163.367
R971 B.n431 B.n221 163.367
R972 B.n435 B.n221 163.367
R973 B.n435 B.n215 163.367
R974 B.n443 B.n215 163.367
R975 B.n443 B.n213 163.367
R976 B.n448 B.n213 163.367
R977 B.n448 B.n208 163.367
R978 B.n457 B.n208 163.367
R979 B.n458 B.n457 163.367
R980 B.n458 B.n5 163.367
R981 B.n6 B.n5 163.367
R982 B.n7 B.n6 163.367
R983 B.n463 B.n7 163.367
R984 B.n463 B.n12 163.367
R985 B.n13 B.n12 163.367
R986 B.n14 B.n13 163.367
R987 B.n468 B.n14 163.367
R988 B.n468 B.n19 163.367
R989 B.n20 B.n19 163.367
R990 B.n21 B.n20 163.367
R991 B.n473 B.n21 163.367
R992 B.n473 B.n26 163.367
R993 B.n27 B.n26 163.367
R994 B.n28 B.n27 163.367
R995 B.n67 B.n28 163.367
R996 B.n74 B.n32 163.367
R997 B.n78 B.n77 163.367
R998 B.n82 B.n81 163.367
R999 B.n86 B.n85 163.367
R1000 B.n90 B.n89 163.367
R1001 B.n94 B.n93 163.367
R1002 B.n98 B.n97 163.367
R1003 B.n102 B.n101 163.367
R1004 B.n106 B.n105 163.367
R1005 B.n110 B.n109 163.367
R1006 B.n114 B.n113 163.367
R1007 B.n118 B.n117 163.367
R1008 B.n122 B.n121 163.367
R1009 B.n126 B.n125 163.367
R1010 B.n130 B.n129 163.367
R1011 B.n134 B.n133 163.367
R1012 B.n138 B.n137 163.367
R1013 B.n142 B.n141 163.367
R1014 B.n146 B.n145 163.367
R1015 B.n150 B.n149 163.367
R1016 B.n154 B.n153 163.367
R1017 B.n158 B.n157 163.367
R1018 B.n162 B.n161 163.367
R1019 B.n166 B.n165 163.367
R1020 B.n170 B.n169 163.367
R1021 B.n174 B.n173 163.367
R1022 B.n178 B.n177 163.367
R1023 B.n182 B.n181 163.367
R1024 B.n186 B.n185 163.367
R1025 B.n190 B.n189 163.367
R1026 B.n194 B.n193 163.367
R1027 B.n198 B.n197 163.367
R1028 B.n202 B.n201 163.367
R1029 B.n204 B.n66 163.367
R1030 B.n410 B.n231 111.028
R1031 B.n482 B.n29 111.028
R1032 B.n412 B.n411 71.676
R1033 B.n269 B.n235 71.676
R1034 B.n404 B.n236 71.676
R1035 B.n400 B.n237 71.676
R1036 B.n396 B.n238 71.676
R1037 B.n392 B.n239 71.676
R1038 B.n388 B.n240 71.676
R1039 B.n384 B.n241 71.676
R1040 B.n380 B.n242 71.676
R1041 B.n376 B.n243 71.676
R1042 B.n372 B.n244 71.676
R1043 B.n368 B.n245 71.676
R1044 B.n364 B.n246 71.676
R1045 B.n360 B.n247 71.676
R1046 B.n356 B.n248 71.676
R1047 B.n351 B.n249 71.676
R1048 B.n347 B.n250 71.676
R1049 B.n343 B.n251 71.676
R1050 B.n339 B.n252 71.676
R1051 B.n335 B.n253 71.676
R1052 B.n330 B.n254 71.676
R1053 B.n326 B.n255 71.676
R1054 B.n322 B.n256 71.676
R1055 B.n318 B.n257 71.676
R1056 B.n314 B.n258 71.676
R1057 B.n310 B.n259 71.676
R1058 B.n306 B.n260 71.676
R1059 B.n302 B.n261 71.676
R1060 B.n298 B.n262 71.676
R1061 B.n294 B.n263 71.676
R1062 B.n290 B.n264 71.676
R1063 B.n286 B.n265 71.676
R1064 B.n282 B.n266 71.676
R1065 B.n278 B.n267 71.676
R1066 B.n484 B.n483 71.676
R1067 B.n74 B.n33 71.676
R1068 B.n78 B.n34 71.676
R1069 B.n82 B.n35 71.676
R1070 B.n86 B.n36 71.676
R1071 B.n90 B.n37 71.676
R1072 B.n94 B.n38 71.676
R1073 B.n98 B.n39 71.676
R1074 B.n102 B.n40 71.676
R1075 B.n106 B.n41 71.676
R1076 B.n110 B.n42 71.676
R1077 B.n114 B.n43 71.676
R1078 B.n118 B.n44 71.676
R1079 B.n122 B.n45 71.676
R1080 B.n126 B.n46 71.676
R1081 B.n130 B.n47 71.676
R1082 B.n134 B.n48 71.676
R1083 B.n138 B.n49 71.676
R1084 B.n142 B.n50 71.676
R1085 B.n146 B.n51 71.676
R1086 B.n150 B.n52 71.676
R1087 B.n154 B.n53 71.676
R1088 B.n158 B.n54 71.676
R1089 B.n162 B.n55 71.676
R1090 B.n166 B.n56 71.676
R1091 B.n170 B.n57 71.676
R1092 B.n174 B.n58 71.676
R1093 B.n178 B.n59 71.676
R1094 B.n182 B.n60 71.676
R1095 B.n186 B.n61 71.676
R1096 B.n190 B.n62 71.676
R1097 B.n194 B.n63 71.676
R1098 B.n198 B.n64 71.676
R1099 B.n202 B.n65 71.676
R1100 B.n481 B.n66 71.676
R1101 B.n481 B.n480 71.676
R1102 B.n204 B.n65 71.676
R1103 B.n201 B.n64 71.676
R1104 B.n197 B.n63 71.676
R1105 B.n193 B.n62 71.676
R1106 B.n189 B.n61 71.676
R1107 B.n185 B.n60 71.676
R1108 B.n181 B.n59 71.676
R1109 B.n177 B.n58 71.676
R1110 B.n173 B.n57 71.676
R1111 B.n169 B.n56 71.676
R1112 B.n165 B.n55 71.676
R1113 B.n161 B.n54 71.676
R1114 B.n157 B.n53 71.676
R1115 B.n153 B.n52 71.676
R1116 B.n149 B.n51 71.676
R1117 B.n145 B.n50 71.676
R1118 B.n141 B.n49 71.676
R1119 B.n137 B.n48 71.676
R1120 B.n133 B.n47 71.676
R1121 B.n129 B.n46 71.676
R1122 B.n125 B.n45 71.676
R1123 B.n121 B.n44 71.676
R1124 B.n117 B.n43 71.676
R1125 B.n113 B.n42 71.676
R1126 B.n109 B.n41 71.676
R1127 B.n105 B.n40 71.676
R1128 B.n101 B.n39 71.676
R1129 B.n97 B.n38 71.676
R1130 B.n93 B.n37 71.676
R1131 B.n89 B.n36 71.676
R1132 B.n85 B.n35 71.676
R1133 B.n81 B.n34 71.676
R1134 B.n77 B.n33 71.676
R1135 B.n483 B.n32 71.676
R1136 B.n411 B.n234 71.676
R1137 B.n405 B.n235 71.676
R1138 B.n401 B.n236 71.676
R1139 B.n397 B.n237 71.676
R1140 B.n393 B.n238 71.676
R1141 B.n389 B.n239 71.676
R1142 B.n385 B.n240 71.676
R1143 B.n381 B.n241 71.676
R1144 B.n377 B.n242 71.676
R1145 B.n373 B.n243 71.676
R1146 B.n369 B.n244 71.676
R1147 B.n365 B.n245 71.676
R1148 B.n361 B.n246 71.676
R1149 B.n357 B.n247 71.676
R1150 B.n352 B.n248 71.676
R1151 B.n348 B.n249 71.676
R1152 B.n344 B.n250 71.676
R1153 B.n340 B.n251 71.676
R1154 B.n336 B.n252 71.676
R1155 B.n331 B.n253 71.676
R1156 B.n327 B.n254 71.676
R1157 B.n323 B.n255 71.676
R1158 B.n319 B.n256 71.676
R1159 B.n315 B.n257 71.676
R1160 B.n311 B.n258 71.676
R1161 B.n307 B.n259 71.676
R1162 B.n303 B.n260 71.676
R1163 B.n299 B.n261 71.676
R1164 B.n295 B.n262 71.676
R1165 B.n291 B.n263 71.676
R1166 B.n287 B.n264 71.676
R1167 B.n283 B.n265 71.676
R1168 B.n279 B.n266 71.676
R1169 B.n275 B.n267 71.676
R1170 B.n333 B.n273 59.5399
R1171 B.n354 B.n271 59.5399
R1172 B.n73 B.n72 59.5399
R1173 B.n70 B.n69 59.5399
R1174 B.n417 B.n231 55.9257
R1175 B.n417 B.n227 55.9257
R1176 B.n424 B.n227 55.9257
R1177 B.n424 B.n423 55.9257
R1178 B.n430 B.n220 55.9257
R1179 B.n436 B.n220 55.9257
R1180 B.n436 B.n216 55.9257
R1181 B.n442 B.n216 55.9257
R1182 B.n450 B.n212 55.9257
R1183 B.n450 B.n449 55.9257
R1184 B.n456 B.n4 55.9257
R1185 B.n515 B.n4 55.9257
R1186 B.n515 B.n514 55.9257
R1187 B.n514 B.n513 55.9257
R1188 B.n507 B.n11 55.9257
R1189 B.n507 B.n506 55.9257
R1190 B.n505 B.n15 55.9257
R1191 B.n499 B.n15 55.9257
R1192 B.n499 B.n498 55.9257
R1193 B.n498 B.n497 55.9257
R1194 B.n491 B.n25 55.9257
R1195 B.n491 B.n490 55.9257
R1196 B.n490 B.n489 55.9257
R1197 B.n489 B.n29 55.9257
R1198 B.n442 B.t2 48.5239
R1199 B.t0 B.n505 48.5239
R1200 B.n456 B.t3 43.5893
R1201 B.n513 B.t1 43.5893
R1202 B.n430 B.t9 38.6547
R1203 B.n497 B.t5 38.6547
R1204 B.n486 B.n485 33.5615
R1205 B.n479 B.n478 33.5615
R1206 B.n274 B.n229 33.5615
R1207 B.n414 B.n413 33.5615
R1208 B B.n517 18.0485
R1209 B.n423 B.t9 17.2715
R1210 B.n25 B.t5 17.2715
R1211 B.n273 B.n272 15.5157
R1212 B.n271 B.n270 15.5157
R1213 B.n72 B.n71 15.5157
R1214 B.n69 B.n68 15.5157
R1215 B.n449 B.t3 12.3369
R1216 B.n11 B.t1 12.3369
R1217 B.n485 B.n31 10.6151
R1218 B.n75 B.n31 10.6151
R1219 B.n76 B.n75 10.6151
R1220 B.n79 B.n76 10.6151
R1221 B.n80 B.n79 10.6151
R1222 B.n83 B.n80 10.6151
R1223 B.n84 B.n83 10.6151
R1224 B.n87 B.n84 10.6151
R1225 B.n88 B.n87 10.6151
R1226 B.n91 B.n88 10.6151
R1227 B.n92 B.n91 10.6151
R1228 B.n95 B.n92 10.6151
R1229 B.n96 B.n95 10.6151
R1230 B.n99 B.n96 10.6151
R1231 B.n100 B.n99 10.6151
R1232 B.n103 B.n100 10.6151
R1233 B.n104 B.n103 10.6151
R1234 B.n107 B.n104 10.6151
R1235 B.n108 B.n107 10.6151
R1236 B.n111 B.n108 10.6151
R1237 B.n112 B.n111 10.6151
R1238 B.n115 B.n112 10.6151
R1239 B.n116 B.n115 10.6151
R1240 B.n119 B.n116 10.6151
R1241 B.n120 B.n119 10.6151
R1242 B.n123 B.n120 10.6151
R1243 B.n124 B.n123 10.6151
R1244 B.n127 B.n124 10.6151
R1245 B.n128 B.n127 10.6151
R1246 B.n132 B.n131 10.6151
R1247 B.n135 B.n132 10.6151
R1248 B.n136 B.n135 10.6151
R1249 B.n139 B.n136 10.6151
R1250 B.n140 B.n139 10.6151
R1251 B.n143 B.n140 10.6151
R1252 B.n144 B.n143 10.6151
R1253 B.n147 B.n144 10.6151
R1254 B.n148 B.n147 10.6151
R1255 B.n152 B.n151 10.6151
R1256 B.n155 B.n152 10.6151
R1257 B.n156 B.n155 10.6151
R1258 B.n159 B.n156 10.6151
R1259 B.n160 B.n159 10.6151
R1260 B.n163 B.n160 10.6151
R1261 B.n164 B.n163 10.6151
R1262 B.n167 B.n164 10.6151
R1263 B.n168 B.n167 10.6151
R1264 B.n171 B.n168 10.6151
R1265 B.n172 B.n171 10.6151
R1266 B.n175 B.n172 10.6151
R1267 B.n176 B.n175 10.6151
R1268 B.n179 B.n176 10.6151
R1269 B.n180 B.n179 10.6151
R1270 B.n183 B.n180 10.6151
R1271 B.n184 B.n183 10.6151
R1272 B.n187 B.n184 10.6151
R1273 B.n188 B.n187 10.6151
R1274 B.n191 B.n188 10.6151
R1275 B.n192 B.n191 10.6151
R1276 B.n195 B.n192 10.6151
R1277 B.n196 B.n195 10.6151
R1278 B.n199 B.n196 10.6151
R1279 B.n200 B.n199 10.6151
R1280 B.n203 B.n200 10.6151
R1281 B.n205 B.n203 10.6151
R1282 B.n206 B.n205 10.6151
R1283 B.n479 B.n206 10.6151
R1284 B.n419 B.n229 10.6151
R1285 B.n420 B.n419 10.6151
R1286 B.n421 B.n420 10.6151
R1287 B.n421 B.n222 10.6151
R1288 B.n432 B.n222 10.6151
R1289 B.n433 B.n432 10.6151
R1290 B.n434 B.n433 10.6151
R1291 B.n434 B.n214 10.6151
R1292 B.n444 B.n214 10.6151
R1293 B.n445 B.n444 10.6151
R1294 B.n447 B.n445 10.6151
R1295 B.n447 B.n446 10.6151
R1296 B.n446 B.n207 10.6151
R1297 B.n459 B.n207 10.6151
R1298 B.n460 B.n459 10.6151
R1299 B.n461 B.n460 10.6151
R1300 B.n462 B.n461 10.6151
R1301 B.n464 B.n462 10.6151
R1302 B.n465 B.n464 10.6151
R1303 B.n466 B.n465 10.6151
R1304 B.n467 B.n466 10.6151
R1305 B.n469 B.n467 10.6151
R1306 B.n470 B.n469 10.6151
R1307 B.n471 B.n470 10.6151
R1308 B.n472 B.n471 10.6151
R1309 B.n474 B.n472 10.6151
R1310 B.n475 B.n474 10.6151
R1311 B.n476 B.n475 10.6151
R1312 B.n477 B.n476 10.6151
R1313 B.n478 B.n477 10.6151
R1314 B.n413 B.n233 10.6151
R1315 B.n408 B.n233 10.6151
R1316 B.n408 B.n407 10.6151
R1317 B.n407 B.n406 10.6151
R1318 B.n406 B.n403 10.6151
R1319 B.n403 B.n402 10.6151
R1320 B.n402 B.n399 10.6151
R1321 B.n399 B.n398 10.6151
R1322 B.n398 B.n395 10.6151
R1323 B.n395 B.n394 10.6151
R1324 B.n394 B.n391 10.6151
R1325 B.n391 B.n390 10.6151
R1326 B.n390 B.n387 10.6151
R1327 B.n387 B.n386 10.6151
R1328 B.n386 B.n383 10.6151
R1329 B.n383 B.n382 10.6151
R1330 B.n382 B.n379 10.6151
R1331 B.n379 B.n378 10.6151
R1332 B.n378 B.n375 10.6151
R1333 B.n375 B.n374 10.6151
R1334 B.n374 B.n371 10.6151
R1335 B.n371 B.n370 10.6151
R1336 B.n370 B.n367 10.6151
R1337 B.n367 B.n366 10.6151
R1338 B.n366 B.n363 10.6151
R1339 B.n363 B.n362 10.6151
R1340 B.n362 B.n359 10.6151
R1341 B.n359 B.n358 10.6151
R1342 B.n358 B.n355 10.6151
R1343 B.n353 B.n350 10.6151
R1344 B.n350 B.n349 10.6151
R1345 B.n349 B.n346 10.6151
R1346 B.n346 B.n345 10.6151
R1347 B.n345 B.n342 10.6151
R1348 B.n342 B.n341 10.6151
R1349 B.n341 B.n338 10.6151
R1350 B.n338 B.n337 10.6151
R1351 B.n337 B.n334 10.6151
R1352 B.n332 B.n329 10.6151
R1353 B.n329 B.n328 10.6151
R1354 B.n328 B.n325 10.6151
R1355 B.n325 B.n324 10.6151
R1356 B.n324 B.n321 10.6151
R1357 B.n321 B.n320 10.6151
R1358 B.n320 B.n317 10.6151
R1359 B.n317 B.n316 10.6151
R1360 B.n316 B.n313 10.6151
R1361 B.n313 B.n312 10.6151
R1362 B.n312 B.n309 10.6151
R1363 B.n309 B.n308 10.6151
R1364 B.n308 B.n305 10.6151
R1365 B.n305 B.n304 10.6151
R1366 B.n304 B.n301 10.6151
R1367 B.n301 B.n300 10.6151
R1368 B.n300 B.n297 10.6151
R1369 B.n297 B.n296 10.6151
R1370 B.n296 B.n293 10.6151
R1371 B.n293 B.n292 10.6151
R1372 B.n292 B.n289 10.6151
R1373 B.n289 B.n288 10.6151
R1374 B.n288 B.n285 10.6151
R1375 B.n285 B.n284 10.6151
R1376 B.n284 B.n281 10.6151
R1377 B.n281 B.n280 10.6151
R1378 B.n280 B.n277 10.6151
R1379 B.n277 B.n276 10.6151
R1380 B.n276 B.n274 10.6151
R1381 B.n415 B.n414 10.6151
R1382 B.n415 B.n225 10.6151
R1383 B.n426 B.n225 10.6151
R1384 B.n427 B.n426 10.6151
R1385 B.n428 B.n427 10.6151
R1386 B.n428 B.n218 10.6151
R1387 B.n438 B.n218 10.6151
R1388 B.n439 B.n438 10.6151
R1389 B.n440 B.n439 10.6151
R1390 B.n440 B.n210 10.6151
R1391 B.n452 B.n210 10.6151
R1392 B.n453 B.n452 10.6151
R1393 B.n454 B.n453 10.6151
R1394 B.n454 B.n0 10.6151
R1395 B.n511 B.n1 10.6151
R1396 B.n511 B.n510 10.6151
R1397 B.n510 B.n509 10.6151
R1398 B.n509 B.n9 10.6151
R1399 B.n503 B.n9 10.6151
R1400 B.n503 B.n502 10.6151
R1401 B.n502 B.n501 10.6151
R1402 B.n501 B.n17 10.6151
R1403 B.n495 B.n17 10.6151
R1404 B.n495 B.n494 10.6151
R1405 B.n494 B.n493 10.6151
R1406 B.n493 B.n23 10.6151
R1407 B.n487 B.n23 10.6151
R1408 B.n487 B.n486 10.6151
R1409 B.n128 B.n73 9.36635
R1410 B.n151 B.n70 9.36635
R1411 B.n355 B.n354 9.36635
R1412 B.n333 B.n332 9.36635
R1413 B.t2 B.n212 7.40237
R1414 B.n506 B.t0 7.40237
R1415 B.n517 B.n0 2.81026
R1416 B.n517 B.n1 2.81026
R1417 B.n131 B.n73 1.24928
R1418 B.n148 B.n70 1.24928
R1419 B.n354 B.n353 1.24928
R1420 B.n334 B.n333 1.24928
R1421 VP.n0 VP.t0 519.904
R1422 VP.n0 VP.t2 519.879
R1423 VP.n2 VP.t1 498.921
R1424 VP.n3 VP.t3 498.921
R1425 VP.n4 VP.n3 161.3
R1426 VP.n2 VP.n1 161.3
R1427 VP.n1 VP.n0 106.987
R1428 VP.n3 VP.n2 48.2005
R1429 VP.n4 VP.n1 0.189894
R1430 VP VP.n4 0.0516364
R1431 VDD1 VDD1.n1 96.6309
R1432 VDD1 VDD1.n0 63.3979
R1433 VDD1.n0 VDD1.t3 2.44494
R1434 VDD1.n0 VDD1.t1 2.44494
R1435 VDD1.n1 VDD1.t2 2.44494
R1436 VDD1.n1 VDD1.t0 2.44494
C0 VN VP 3.93304f
C1 VDD1 VP 1.95759f
C2 VDD2 VP 0.259207f
C3 VN VTAIL 1.55355f
C4 VTAIL VDD1 5.76766f
C5 VTAIL VDD2 5.80759f
C6 VTAIL VP 1.56766f
C7 VN VDD1 0.147512f
C8 VN VDD2 1.8461f
C9 VDD2 VDD1 0.516926f
C10 VDD2 B 2.251829f
C11 VDD1 B 4.75409f
C12 VTAIL B 6.42629f
C13 VN B 5.92647f
C14 VP B 4.133857f
C15 VDD1.t3 B 0.141718f
C16 VDD1.t1 B 0.141718f
C17 VDD1.n0 B 1.21979f
C18 VDD1.t2 B 0.141718f
C19 VDD1.t0 B 0.141718f
C20 VDD1.n1 B 1.60073f
C21 VP.t2 B 0.329934f
C22 VP.t0 B 0.329942f
C23 VP.n0 B 0.617141f
C24 VP.n1 B 1.65631f
C25 VP.t1 B 0.324216f
C26 VP.n2 B 0.141844f
C27 VP.t3 B 0.324216f
C28 VP.n3 B 0.141844f
C29 VP.n4 B 0.022955f
C30 VTAIL.n0 B 0.020622f
C31 VTAIL.n1 B 0.01426f
C32 VTAIL.n2 B 0.007663f
C33 VTAIL.n3 B 0.018112f
C34 VTAIL.n4 B 0.008114f
C35 VTAIL.n5 B 0.01426f
C36 VTAIL.n6 B 0.007663f
C37 VTAIL.n7 B 0.018112f
C38 VTAIL.n8 B 0.008114f
C39 VTAIL.n9 B 0.01426f
C40 VTAIL.n10 B 0.007663f
C41 VTAIL.n11 B 0.018112f
C42 VTAIL.n12 B 0.008114f
C43 VTAIL.n13 B 0.068367f
C44 VTAIL.t3 B 0.029541f
C45 VTAIL.n14 B 0.013584f
C46 VTAIL.n15 B 0.0107f
C47 VTAIL.n16 B 0.007663f
C48 VTAIL.n17 B 0.476811f
C49 VTAIL.n18 B 0.01426f
C50 VTAIL.n19 B 0.007663f
C51 VTAIL.n20 B 0.008114f
C52 VTAIL.n21 B 0.018112f
C53 VTAIL.n22 B 0.018112f
C54 VTAIL.n23 B 0.008114f
C55 VTAIL.n24 B 0.007663f
C56 VTAIL.n25 B 0.01426f
C57 VTAIL.n26 B 0.01426f
C58 VTAIL.n27 B 0.007663f
C59 VTAIL.n28 B 0.008114f
C60 VTAIL.n29 B 0.018112f
C61 VTAIL.n30 B 0.018112f
C62 VTAIL.n31 B 0.008114f
C63 VTAIL.n32 B 0.007663f
C64 VTAIL.n33 B 0.01426f
C65 VTAIL.n34 B 0.01426f
C66 VTAIL.n35 B 0.007663f
C67 VTAIL.n36 B 0.008114f
C68 VTAIL.n37 B 0.018112f
C69 VTAIL.n38 B 0.040231f
C70 VTAIL.n39 B 0.008114f
C71 VTAIL.n40 B 0.007663f
C72 VTAIL.n41 B 0.031794f
C73 VTAIL.n42 B 0.022579f
C74 VTAIL.n43 B 0.051628f
C75 VTAIL.n44 B 0.020622f
C76 VTAIL.n45 B 0.01426f
C77 VTAIL.n46 B 0.007663f
C78 VTAIL.n47 B 0.018112f
C79 VTAIL.n48 B 0.008114f
C80 VTAIL.n49 B 0.01426f
C81 VTAIL.n50 B 0.007663f
C82 VTAIL.n51 B 0.018112f
C83 VTAIL.n52 B 0.008114f
C84 VTAIL.n53 B 0.01426f
C85 VTAIL.n54 B 0.007663f
C86 VTAIL.n55 B 0.018112f
C87 VTAIL.n56 B 0.008114f
C88 VTAIL.n57 B 0.068367f
C89 VTAIL.t7 B 0.029541f
C90 VTAIL.n58 B 0.013584f
C91 VTAIL.n59 B 0.0107f
C92 VTAIL.n60 B 0.007663f
C93 VTAIL.n61 B 0.476811f
C94 VTAIL.n62 B 0.01426f
C95 VTAIL.n63 B 0.007663f
C96 VTAIL.n64 B 0.008114f
C97 VTAIL.n65 B 0.018112f
C98 VTAIL.n66 B 0.018112f
C99 VTAIL.n67 B 0.008114f
C100 VTAIL.n68 B 0.007663f
C101 VTAIL.n69 B 0.01426f
C102 VTAIL.n70 B 0.01426f
C103 VTAIL.n71 B 0.007663f
C104 VTAIL.n72 B 0.008114f
C105 VTAIL.n73 B 0.018112f
C106 VTAIL.n74 B 0.018112f
C107 VTAIL.n75 B 0.008114f
C108 VTAIL.n76 B 0.007663f
C109 VTAIL.n77 B 0.01426f
C110 VTAIL.n78 B 0.01426f
C111 VTAIL.n79 B 0.007663f
C112 VTAIL.n80 B 0.008114f
C113 VTAIL.n81 B 0.018112f
C114 VTAIL.n82 B 0.040231f
C115 VTAIL.n83 B 0.008114f
C116 VTAIL.n84 B 0.007663f
C117 VTAIL.n85 B 0.031794f
C118 VTAIL.n86 B 0.022579f
C119 VTAIL.n87 B 0.064799f
C120 VTAIL.n88 B 0.020622f
C121 VTAIL.n89 B 0.01426f
C122 VTAIL.n90 B 0.007663f
C123 VTAIL.n91 B 0.018112f
C124 VTAIL.n92 B 0.008114f
C125 VTAIL.n93 B 0.01426f
C126 VTAIL.n94 B 0.007663f
C127 VTAIL.n95 B 0.018112f
C128 VTAIL.n96 B 0.008114f
C129 VTAIL.n97 B 0.01426f
C130 VTAIL.n98 B 0.007663f
C131 VTAIL.n99 B 0.018112f
C132 VTAIL.n100 B 0.008114f
C133 VTAIL.n101 B 0.068367f
C134 VTAIL.t2 B 0.029541f
C135 VTAIL.n102 B 0.013584f
C136 VTAIL.n103 B 0.0107f
C137 VTAIL.n104 B 0.007663f
C138 VTAIL.n105 B 0.476811f
C139 VTAIL.n106 B 0.01426f
C140 VTAIL.n107 B 0.007663f
C141 VTAIL.n108 B 0.008114f
C142 VTAIL.n109 B 0.018112f
C143 VTAIL.n110 B 0.018112f
C144 VTAIL.n111 B 0.008114f
C145 VTAIL.n112 B 0.007663f
C146 VTAIL.n113 B 0.01426f
C147 VTAIL.n114 B 0.01426f
C148 VTAIL.n115 B 0.007663f
C149 VTAIL.n116 B 0.008114f
C150 VTAIL.n117 B 0.018112f
C151 VTAIL.n118 B 0.018112f
C152 VTAIL.n119 B 0.008114f
C153 VTAIL.n120 B 0.007663f
C154 VTAIL.n121 B 0.01426f
C155 VTAIL.n122 B 0.01426f
C156 VTAIL.n123 B 0.007663f
C157 VTAIL.n124 B 0.008114f
C158 VTAIL.n125 B 0.018112f
C159 VTAIL.n126 B 0.040231f
C160 VTAIL.n127 B 0.008114f
C161 VTAIL.n128 B 0.007663f
C162 VTAIL.n129 B 0.031794f
C163 VTAIL.n130 B 0.022579f
C164 VTAIL.n131 B 0.589473f
C165 VTAIL.n132 B 0.020622f
C166 VTAIL.n133 B 0.01426f
C167 VTAIL.n134 B 0.007663f
C168 VTAIL.n135 B 0.018112f
C169 VTAIL.n136 B 0.008114f
C170 VTAIL.n137 B 0.01426f
C171 VTAIL.n138 B 0.007663f
C172 VTAIL.n139 B 0.018112f
C173 VTAIL.n140 B 0.008114f
C174 VTAIL.n141 B 0.01426f
C175 VTAIL.n142 B 0.007663f
C176 VTAIL.n143 B 0.018112f
C177 VTAIL.n144 B 0.008114f
C178 VTAIL.n145 B 0.068367f
C179 VTAIL.t6 B 0.029541f
C180 VTAIL.n146 B 0.013584f
C181 VTAIL.n147 B 0.0107f
C182 VTAIL.n148 B 0.007663f
C183 VTAIL.n149 B 0.476811f
C184 VTAIL.n150 B 0.01426f
C185 VTAIL.n151 B 0.007663f
C186 VTAIL.n152 B 0.008114f
C187 VTAIL.n153 B 0.018112f
C188 VTAIL.n154 B 0.018112f
C189 VTAIL.n155 B 0.008114f
C190 VTAIL.n156 B 0.007663f
C191 VTAIL.n157 B 0.01426f
C192 VTAIL.n158 B 0.01426f
C193 VTAIL.n159 B 0.007663f
C194 VTAIL.n160 B 0.008114f
C195 VTAIL.n161 B 0.018112f
C196 VTAIL.n162 B 0.018112f
C197 VTAIL.n163 B 0.008114f
C198 VTAIL.n164 B 0.007663f
C199 VTAIL.n165 B 0.01426f
C200 VTAIL.n166 B 0.01426f
C201 VTAIL.n167 B 0.007663f
C202 VTAIL.n168 B 0.008114f
C203 VTAIL.n169 B 0.018112f
C204 VTAIL.n170 B 0.040231f
C205 VTAIL.n171 B 0.008114f
C206 VTAIL.n172 B 0.007663f
C207 VTAIL.n173 B 0.031794f
C208 VTAIL.n174 B 0.022579f
C209 VTAIL.n175 B 0.589473f
C210 VTAIL.n176 B 0.020622f
C211 VTAIL.n177 B 0.01426f
C212 VTAIL.n178 B 0.007663f
C213 VTAIL.n179 B 0.018112f
C214 VTAIL.n180 B 0.008114f
C215 VTAIL.n181 B 0.01426f
C216 VTAIL.n182 B 0.007663f
C217 VTAIL.n183 B 0.018112f
C218 VTAIL.n184 B 0.008114f
C219 VTAIL.n185 B 0.01426f
C220 VTAIL.n186 B 0.007663f
C221 VTAIL.n187 B 0.018112f
C222 VTAIL.n188 B 0.008114f
C223 VTAIL.n189 B 0.068367f
C224 VTAIL.t4 B 0.029541f
C225 VTAIL.n190 B 0.013584f
C226 VTAIL.n191 B 0.0107f
C227 VTAIL.n192 B 0.007663f
C228 VTAIL.n193 B 0.476811f
C229 VTAIL.n194 B 0.01426f
C230 VTAIL.n195 B 0.007663f
C231 VTAIL.n196 B 0.008114f
C232 VTAIL.n197 B 0.018112f
C233 VTAIL.n198 B 0.018112f
C234 VTAIL.n199 B 0.008114f
C235 VTAIL.n200 B 0.007663f
C236 VTAIL.n201 B 0.01426f
C237 VTAIL.n202 B 0.01426f
C238 VTAIL.n203 B 0.007663f
C239 VTAIL.n204 B 0.008114f
C240 VTAIL.n205 B 0.018112f
C241 VTAIL.n206 B 0.018112f
C242 VTAIL.n207 B 0.008114f
C243 VTAIL.n208 B 0.007663f
C244 VTAIL.n209 B 0.01426f
C245 VTAIL.n210 B 0.01426f
C246 VTAIL.n211 B 0.007663f
C247 VTAIL.n212 B 0.008114f
C248 VTAIL.n213 B 0.018112f
C249 VTAIL.n214 B 0.040231f
C250 VTAIL.n215 B 0.008114f
C251 VTAIL.n216 B 0.007663f
C252 VTAIL.n217 B 0.031794f
C253 VTAIL.n218 B 0.022579f
C254 VTAIL.n219 B 0.064799f
C255 VTAIL.n220 B 0.020622f
C256 VTAIL.n221 B 0.01426f
C257 VTAIL.n222 B 0.007663f
C258 VTAIL.n223 B 0.018112f
C259 VTAIL.n224 B 0.008114f
C260 VTAIL.n225 B 0.01426f
C261 VTAIL.n226 B 0.007663f
C262 VTAIL.n227 B 0.018112f
C263 VTAIL.n228 B 0.008114f
C264 VTAIL.n229 B 0.01426f
C265 VTAIL.n230 B 0.007663f
C266 VTAIL.n231 B 0.018112f
C267 VTAIL.n232 B 0.008114f
C268 VTAIL.n233 B 0.068367f
C269 VTAIL.t1 B 0.029541f
C270 VTAIL.n234 B 0.013584f
C271 VTAIL.n235 B 0.0107f
C272 VTAIL.n236 B 0.007663f
C273 VTAIL.n237 B 0.476811f
C274 VTAIL.n238 B 0.01426f
C275 VTAIL.n239 B 0.007663f
C276 VTAIL.n240 B 0.008114f
C277 VTAIL.n241 B 0.018112f
C278 VTAIL.n242 B 0.018112f
C279 VTAIL.n243 B 0.008114f
C280 VTAIL.n244 B 0.007663f
C281 VTAIL.n245 B 0.01426f
C282 VTAIL.n246 B 0.01426f
C283 VTAIL.n247 B 0.007663f
C284 VTAIL.n248 B 0.008114f
C285 VTAIL.n249 B 0.018112f
C286 VTAIL.n250 B 0.018112f
C287 VTAIL.n251 B 0.008114f
C288 VTAIL.n252 B 0.007663f
C289 VTAIL.n253 B 0.01426f
C290 VTAIL.n254 B 0.01426f
C291 VTAIL.n255 B 0.007663f
C292 VTAIL.n256 B 0.008114f
C293 VTAIL.n257 B 0.018112f
C294 VTAIL.n258 B 0.040231f
C295 VTAIL.n259 B 0.008114f
C296 VTAIL.n260 B 0.007663f
C297 VTAIL.n261 B 0.031794f
C298 VTAIL.n262 B 0.022579f
C299 VTAIL.n263 B 0.064799f
C300 VTAIL.n264 B 0.020622f
C301 VTAIL.n265 B 0.01426f
C302 VTAIL.n266 B 0.007663f
C303 VTAIL.n267 B 0.018112f
C304 VTAIL.n268 B 0.008114f
C305 VTAIL.n269 B 0.01426f
C306 VTAIL.n270 B 0.007663f
C307 VTAIL.n271 B 0.018112f
C308 VTAIL.n272 B 0.008114f
C309 VTAIL.n273 B 0.01426f
C310 VTAIL.n274 B 0.007663f
C311 VTAIL.n275 B 0.018112f
C312 VTAIL.n276 B 0.008114f
C313 VTAIL.n277 B 0.068367f
C314 VTAIL.t0 B 0.029541f
C315 VTAIL.n278 B 0.013584f
C316 VTAIL.n279 B 0.0107f
C317 VTAIL.n280 B 0.007663f
C318 VTAIL.n281 B 0.476811f
C319 VTAIL.n282 B 0.01426f
C320 VTAIL.n283 B 0.007663f
C321 VTAIL.n284 B 0.008114f
C322 VTAIL.n285 B 0.018112f
C323 VTAIL.n286 B 0.018112f
C324 VTAIL.n287 B 0.008114f
C325 VTAIL.n288 B 0.007663f
C326 VTAIL.n289 B 0.01426f
C327 VTAIL.n290 B 0.01426f
C328 VTAIL.n291 B 0.007663f
C329 VTAIL.n292 B 0.008114f
C330 VTAIL.n293 B 0.018112f
C331 VTAIL.n294 B 0.018112f
C332 VTAIL.n295 B 0.008114f
C333 VTAIL.n296 B 0.007663f
C334 VTAIL.n297 B 0.01426f
C335 VTAIL.n298 B 0.01426f
C336 VTAIL.n299 B 0.007663f
C337 VTAIL.n300 B 0.008114f
C338 VTAIL.n301 B 0.018112f
C339 VTAIL.n302 B 0.040231f
C340 VTAIL.n303 B 0.008114f
C341 VTAIL.n304 B 0.007663f
C342 VTAIL.n305 B 0.031794f
C343 VTAIL.n306 B 0.022579f
C344 VTAIL.n307 B 0.589473f
C345 VTAIL.n308 B 0.020622f
C346 VTAIL.n309 B 0.01426f
C347 VTAIL.n310 B 0.007663f
C348 VTAIL.n311 B 0.018112f
C349 VTAIL.n312 B 0.008114f
C350 VTAIL.n313 B 0.01426f
C351 VTAIL.n314 B 0.007663f
C352 VTAIL.n315 B 0.018112f
C353 VTAIL.n316 B 0.008114f
C354 VTAIL.n317 B 0.01426f
C355 VTAIL.n318 B 0.007663f
C356 VTAIL.n319 B 0.018112f
C357 VTAIL.n320 B 0.008114f
C358 VTAIL.n321 B 0.068367f
C359 VTAIL.t5 B 0.029541f
C360 VTAIL.n322 B 0.013584f
C361 VTAIL.n323 B 0.0107f
C362 VTAIL.n324 B 0.007663f
C363 VTAIL.n325 B 0.476811f
C364 VTAIL.n326 B 0.01426f
C365 VTAIL.n327 B 0.007663f
C366 VTAIL.n328 B 0.008114f
C367 VTAIL.n329 B 0.018112f
C368 VTAIL.n330 B 0.018112f
C369 VTAIL.n331 B 0.008114f
C370 VTAIL.n332 B 0.007663f
C371 VTAIL.n333 B 0.01426f
C372 VTAIL.n334 B 0.01426f
C373 VTAIL.n335 B 0.007663f
C374 VTAIL.n336 B 0.008114f
C375 VTAIL.n337 B 0.018112f
C376 VTAIL.n338 B 0.018112f
C377 VTAIL.n339 B 0.008114f
C378 VTAIL.n340 B 0.007663f
C379 VTAIL.n341 B 0.01426f
C380 VTAIL.n342 B 0.01426f
C381 VTAIL.n343 B 0.007663f
C382 VTAIL.n344 B 0.008114f
C383 VTAIL.n345 B 0.018112f
C384 VTAIL.n346 B 0.040231f
C385 VTAIL.n347 B 0.008114f
C386 VTAIL.n348 B 0.007663f
C387 VTAIL.n349 B 0.031794f
C388 VTAIL.n350 B 0.022579f
C389 VTAIL.n351 B 0.570954f
C390 VDD2.t0 B 0.143744f
C391 VDD2.t2 B 0.143744f
C392 VDD2.n0 B 1.6039f
C393 VDD2.t3 B 0.143744f
C394 VDD2.t1 B 0.143744f
C395 VDD2.n1 B 1.237f
C396 VDD2.n2 B 2.32938f
C397 VN.t3 B 0.326457f
C398 VN.t1 B 0.326449f
C399 VN.n0 B 0.26945f
C400 VN.t2 B 0.326457f
C401 VN.t0 B 0.326449f
C402 VN.n1 B 0.619648f
.ends

