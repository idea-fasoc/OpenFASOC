* NGSPICE file created from diff_pair_sample_0968.ext - technology: sky130A

.subckt diff_pair_sample_0968 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=3.1746 ps=19.57 w=19.24 l=0.78
X1 VDD1.t8 VP.t1 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=3.1746 ps=19.57 w=19.24 l=0.78
X2 VDD2.t9 VN.t0 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X3 VDD1.t7 VP.t2 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=7.5036 ps=39.26 w=19.24 l=0.78
X4 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=0 ps=0 w=19.24 l=0.78
X5 VDD1.t6 VP.t3 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=7.5036 ps=39.26 w=19.24 l=0.78
X6 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=0 ps=0 w=19.24 l=0.78
X7 VDD2.t8 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=7.5036 ps=39.26 w=19.24 l=0.78
X8 VDD2.t7 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=3.1746 ps=19.57 w=19.24 l=0.78
X9 VTAIL.t8 VN.t3 VDD2.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X10 VTAIL.t16 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X11 VDD2.t5 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=7.5036 ps=39.26 w=19.24 l=0.78
X12 VTAIL.t5 VN.t5 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X13 VTAIL.t6 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X14 VDD1.t4 VP.t5 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=0 ps=0 w=19.24 l=0.78
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=0 ps=0 w=19.24 l=0.78
X17 VDD1.t3 VP.t6 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X18 VTAIL.t14 VP.t7 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X19 VTAIL.t2 VN.t7 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X20 VDD2.t1 VN.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5036 pd=39.26 as=3.1746 ps=19.57 w=19.24 l=0.78
X21 VDD2.t0 VN.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X22 VTAIL.t17 VP.t8 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
X23 VTAIL.t13 VP.t9 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1746 pd=19.57 as=3.1746 ps=19.57 w=19.24 l=0.78
R0 VP.n6 VP.t0 666.87
R1 VP.n14 VP.t1 644.831
R2 VP.n16 VP.t7 644.831
R3 VP.n1 VP.t5 644.831
R4 VP.n20 VP.t8 644.831
R5 VP.n22 VP.t3 644.831
R6 VP.n11 VP.t2 644.831
R7 VP.n9 VP.t9 644.831
R8 VP.n8 VP.t6 644.831
R9 VP.n7 VP.t4 644.831
R10 VP.n23 VP.n22 161.3
R11 VP.n10 VP.n3 161.3
R12 VP.n12 VP.n11 161.3
R13 VP.n21 VP.n0 161.3
R14 VP.n15 VP.n2 161.3
R15 VP.n14 VP.n13 161.3
R16 VP.n8 VP.n5 80.6037
R17 VP.n9 VP.n4 80.6037
R18 VP.n20 VP.n19 80.6037
R19 VP.n18 VP.n1 80.6037
R20 VP.n17 VP.n16 80.6037
R21 VP.n13 VP.n12 48.6558
R22 VP.n16 VP.n1 48.2005
R23 VP.n20 VP.n1 48.2005
R24 VP.n9 VP.n8 48.2005
R25 VP.n8 VP.n7 48.2005
R26 VP.n16 VP.n15 36.5157
R27 VP.n21 VP.n20 36.5157
R28 VP.n10 VP.n9 36.5157
R29 VP.n6 VP.n5 31.7379
R30 VP.n7 VP.n6 16.9109
R31 VP.n15 VP.n14 11.6853
R32 VP.n22 VP.n21 11.6853
R33 VP.n11 VP.n10 11.6853
R34 VP.n5 VP.n4 0.380177
R35 VP.n18 VP.n17 0.380177
R36 VP.n19 VP.n18 0.380177
R37 VP.n4 VP.n3 0.285035
R38 VP.n17 VP.n2 0.285035
R39 VP.n19 VP.n0 0.285035
R40 VP.n12 VP.n3 0.189894
R41 VP.n13 VP.n2 0.189894
R42 VP.n23 VP.n0 0.189894
R43 VP VP.n23 0.0516364
R44 VTAIL.n11 VTAIL.t7 43.4099
R45 VTAIL.n16 VTAIL.t18 43.4097
R46 VTAIL.n17 VTAIL.t1 43.4097
R47 VTAIL.n2 VTAIL.t10 43.4097
R48 VTAIL.n15 VTAIL.n14 42.3808
R49 VTAIL.n13 VTAIL.n12 42.3808
R50 VTAIL.n10 VTAIL.n9 42.3808
R51 VTAIL.n8 VTAIL.n7 42.3808
R52 VTAIL.n19 VTAIL.n18 42.3808
R53 VTAIL.n1 VTAIL.n0 42.3808
R54 VTAIL.n4 VTAIL.n3 42.3808
R55 VTAIL.n6 VTAIL.n5 42.3808
R56 VTAIL.n8 VTAIL.n6 30.8669
R57 VTAIL.n17 VTAIL.n16 29.91
R58 VTAIL.n18 VTAIL.t0 1.02961
R59 VTAIL.n18 VTAIL.t6 1.02961
R60 VTAIL.n0 VTAIL.t4 1.02961
R61 VTAIL.n0 VTAIL.t8 1.02961
R62 VTAIL.n3 VTAIL.t12 1.02961
R63 VTAIL.n3 VTAIL.t17 1.02961
R64 VTAIL.n5 VTAIL.t15 1.02961
R65 VTAIL.n5 VTAIL.t14 1.02961
R66 VTAIL.n14 VTAIL.t11 1.02961
R67 VTAIL.n14 VTAIL.t13 1.02961
R68 VTAIL.n12 VTAIL.t9 1.02961
R69 VTAIL.n12 VTAIL.t16 1.02961
R70 VTAIL.n9 VTAIL.t19 1.02961
R71 VTAIL.n9 VTAIL.t2 1.02961
R72 VTAIL.n7 VTAIL.t3 1.02961
R73 VTAIL.n7 VTAIL.t5 1.02961
R74 VTAIL.n10 VTAIL.n8 0.957397
R75 VTAIL.n11 VTAIL.n10 0.957397
R76 VTAIL.n15 VTAIL.n13 0.957397
R77 VTAIL.n16 VTAIL.n15 0.957397
R78 VTAIL.n6 VTAIL.n4 0.957397
R79 VTAIL.n4 VTAIL.n2 0.957397
R80 VTAIL.n19 VTAIL.n17 0.957397
R81 VTAIL.n13 VTAIL.n11 0.948776
R82 VTAIL.n2 VTAIL.n1 0.948776
R83 VTAIL VTAIL.n1 0.776362
R84 VTAIL VTAIL.n19 0.181534
R85 VDD1.n1 VDD1.t9 61.0456
R86 VDD1.n3 VDD1.t8 61.0454
R87 VDD1.n5 VDD1.n4 59.7219
R88 VDD1.n1 VDD1.n0 59.0596
R89 VDD1.n3 VDD1.n2 59.0596
R90 VDD1.n7 VDD1.n6 59.0594
R91 VDD1.n7 VDD1.n5 45.9082
R92 VDD1.n6 VDD1.t0 1.02961
R93 VDD1.n6 VDD1.t7 1.02961
R94 VDD1.n0 VDD1.t5 1.02961
R95 VDD1.n0 VDD1.t3 1.02961
R96 VDD1.n4 VDD1.t1 1.02961
R97 VDD1.n4 VDD1.t6 1.02961
R98 VDD1.n2 VDD1.t2 1.02961
R99 VDD1.n2 VDD1.t4 1.02961
R100 VDD1 VDD1.n7 0.659983
R101 VDD1 VDD1.n1 0.297914
R102 VDD1.n5 VDD1.n3 0.184378
R103 B.n126 B.t21 796.549
R104 B.n123 B.t17 796.549
R105 B.n514 B.t10 796.549
R106 B.n511 B.t14 796.549
R107 B.n904 B.n903 585
R108 B.n905 B.n904 585
R109 B.n391 B.n121 585
R110 B.n390 B.n389 585
R111 B.n388 B.n387 585
R112 B.n386 B.n385 585
R113 B.n384 B.n383 585
R114 B.n382 B.n381 585
R115 B.n380 B.n379 585
R116 B.n378 B.n377 585
R117 B.n376 B.n375 585
R118 B.n374 B.n373 585
R119 B.n372 B.n371 585
R120 B.n370 B.n369 585
R121 B.n368 B.n367 585
R122 B.n366 B.n365 585
R123 B.n364 B.n363 585
R124 B.n362 B.n361 585
R125 B.n360 B.n359 585
R126 B.n358 B.n357 585
R127 B.n356 B.n355 585
R128 B.n354 B.n353 585
R129 B.n352 B.n351 585
R130 B.n350 B.n349 585
R131 B.n348 B.n347 585
R132 B.n346 B.n345 585
R133 B.n344 B.n343 585
R134 B.n342 B.n341 585
R135 B.n340 B.n339 585
R136 B.n338 B.n337 585
R137 B.n336 B.n335 585
R138 B.n334 B.n333 585
R139 B.n332 B.n331 585
R140 B.n330 B.n329 585
R141 B.n328 B.n327 585
R142 B.n326 B.n325 585
R143 B.n324 B.n323 585
R144 B.n322 B.n321 585
R145 B.n320 B.n319 585
R146 B.n318 B.n317 585
R147 B.n316 B.n315 585
R148 B.n314 B.n313 585
R149 B.n312 B.n311 585
R150 B.n310 B.n309 585
R151 B.n308 B.n307 585
R152 B.n306 B.n305 585
R153 B.n304 B.n303 585
R154 B.n302 B.n301 585
R155 B.n300 B.n299 585
R156 B.n298 B.n297 585
R157 B.n296 B.n295 585
R158 B.n294 B.n293 585
R159 B.n292 B.n291 585
R160 B.n290 B.n289 585
R161 B.n288 B.n287 585
R162 B.n286 B.n285 585
R163 B.n284 B.n283 585
R164 B.n282 B.n281 585
R165 B.n280 B.n279 585
R166 B.n278 B.n277 585
R167 B.n276 B.n275 585
R168 B.n274 B.n273 585
R169 B.n272 B.n271 585
R170 B.n270 B.n269 585
R171 B.n268 B.n267 585
R172 B.n266 B.n265 585
R173 B.n264 B.n263 585
R174 B.n262 B.n261 585
R175 B.n260 B.n259 585
R176 B.n258 B.n257 585
R177 B.n256 B.n255 585
R178 B.n254 B.n253 585
R179 B.n252 B.n251 585
R180 B.n249 B.n248 585
R181 B.n247 B.n246 585
R182 B.n245 B.n244 585
R183 B.n243 B.n242 585
R184 B.n241 B.n240 585
R185 B.n239 B.n238 585
R186 B.n237 B.n236 585
R187 B.n235 B.n234 585
R188 B.n233 B.n232 585
R189 B.n231 B.n230 585
R190 B.n229 B.n228 585
R191 B.n227 B.n226 585
R192 B.n225 B.n224 585
R193 B.n223 B.n222 585
R194 B.n221 B.n220 585
R195 B.n219 B.n218 585
R196 B.n217 B.n216 585
R197 B.n215 B.n214 585
R198 B.n213 B.n212 585
R199 B.n211 B.n210 585
R200 B.n209 B.n208 585
R201 B.n207 B.n206 585
R202 B.n205 B.n204 585
R203 B.n203 B.n202 585
R204 B.n201 B.n200 585
R205 B.n199 B.n198 585
R206 B.n197 B.n196 585
R207 B.n195 B.n194 585
R208 B.n193 B.n192 585
R209 B.n191 B.n190 585
R210 B.n189 B.n188 585
R211 B.n187 B.n186 585
R212 B.n185 B.n184 585
R213 B.n183 B.n182 585
R214 B.n181 B.n180 585
R215 B.n179 B.n178 585
R216 B.n177 B.n176 585
R217 B.n175 B.n174 585
R218 B.n173 B.n172 585
R219 B.n171 B.n170 585
R220 B.n169 B.n168 585
R221 B.n167 B.n166 585
R222 B.n165 B.n164 585
R223 B.n163 B.n162 585
R224 B.n161 B.n160 585
R225 B.n159 B.n158 585
R226 B.n157 B.n156 585
R227 B.n155 B.n154 585
R228 B.n153 B.n152 585
R229 B.n151 B.n150 585
R230 B.n149 B.n148 585
R231 B.n147 B.n146 585
R232 B.n145 B.n144 585
R233 B.n143 B.n142 585
R234 B.n141 B.n140 585
R235 B.n139 B.n138 585
R236 B.n137 B.n136 585
R237 B.n135 B.n134 585
R238 B.n133 B.n132 585
R239 B.n131 B.n130 585
R240 B.n129 B.n128 585
R241 B.n54 B.n53 585
R242 B.n908 B.n907 585
R243 B.n902 B.n122 585
R244 B.n122 B.n51 585
R245 B.n901 B.n50 585
R246 B.n912 B.n50 585
R247 B.n900 B.n49 585
R248 B.n913 B.n49 585
R249 B.n899 B.n48 585
R250 B.n914 B.n48 585
R251 B.n898 B.n897 585
R252 B.n897 B.n47 585
R253 B.n896 B.n43 585
R254 B.n920 B.n43 585
R255 B.n895 B.n42 585
R256 B.n921 B.n42 585
R257 B.n894 B.n41 585
R258 B.n922 B.n41 585
R259 B.n893 B.n892 585
R260 B.n892 B.n37 585
R261 B.n891 B.n36 585
R262 B.n928 B.n36 585
R263 B.n890 B.n35 585
R264 B.n929 B.n35 585
R265 B.n889 B.n34 585
R266 B.n930 B.n34 585
R267 B.n888 B.n887 585
R268 B.n887 B.n30 585
R269 B.n886 B.n29 585
R270 B.n936 B.n29 585
R271 B.n885 B.n28 585
R272 B.n937 B.n28 585
R273 B.n884 B.n27 585
R274 B.n938 B.n27 585
R275 B.n883 B.n882 585
R276 B.n882 B.n23 585
R277 B.n881 B.n22 585
R278 B.n944 B.n22 585
R279 B.n880 B.n21 585
R280 B.n945 B.n21 585
R281 B.n879 B.n20 585
R282 B.n946 B.n20 585
R283 B.n878 B.n877 585
R284 B.n877 B.n16 585
R285 B.n876 B.n15 585
R286 B.t8 B.n15 585
R287 B.n875 B.n14 585
R288 B.n952 B.n14 585
R289 B.n874 B.n13 585
R290 B.n953 B.n13 585
R291 B.n873 B.n872 585
R292 B.n872 B.n12 585
R293 B.n871 B.n870 585
R294 B.n871 B.n8 585
R295 B.n869 B.n7 585
R296 B.n960 B.n7 585
R297 B.n868 B.n6 585
R298 B.n961 B.n6 585
R299 B.n867 B.n5 585
R300 B.n962 B.n5 585
R301 B.n866 B.n865 585
R302 B.n865 B.n4 585
R303 B.n864 B.n392 585
R304 B.n864 B.n863 585
R305 B.n853 B.n393 585
R306 B.n856 B.n393 585
R307 B.n855 B.n854 585
R308 B.n857 B.n855 585
R309 B.n852 B.n398 585
R310 B.n398 B.n397 585
R311 B.n851 B.n850 585
R312 B.n850 B.t2 585
R313 B.n400 B.n399 585
R314 B.n401 B.n400 585
R315 B.n843 B.n842 585
R316 B.n844 B.n843 585
R317 B.n841 B.n406 585
R318 B.n406 B.n405 585
R319 B.n840 B.n839 585
R320 B.n839 B.n838 585
R321 B.n408 B.n407 585
R322 B.n409 B.n408 585
R323 B.n831 B.n830 585
R324 B.n832 B.n831 585
R325 B.n829 B.n413 585
R326 B.n417 B.n413 585
R327 B.n828 B.n827 585
R328 B.n827 B.n826 585
R329 B.n415 B.n414 585
R330 B.n416 B.n415 585
R331 B.n819 B.n818 585
R332 B.n820 B.n819 585
R333 B.n817 B.n422 585
R334 B.n422 B.n421 585
R335 B.n816 B.n815 585
R336 B.n815 B.n814 585
R337 B.n424 B.n423 585
R338 B.n425 B.n424 585
R339 B.n807 B.n806 585
R340 B.n808 B.n807 585
R341 B.n805 B.n430 585
R342 B.n430 B.n429 585
R343 B.n804 B.n803 585
R344 B.n803 B.n802 585
R345 B.n432 B.n431 585
R346 B.n795 B.n432 585
R347 B.n794 B.n793 585
R348 B.n796 B.n794 585
R349 B.n792 B.n437 585
R350 B.n437 B.n436 585
R351 B.n791 B.n790 585
R352 B.n790 B.n789 585
R353 B.n439 B.n438 585
R354 B.n440 B.n439 585
R355 B.n785 B.n784 585
R356 B.n443 B.n442 585
R357 B.n781 B.n780 585
R358 B.n782 B.n781 585
R359 B.n779 B.n510 585
R360 B.n778 B.n777 585
R361 B.n776 B.n775 585
R362 B.n774 B.n773 585
R363 B.n772 B.n771 585
R364 B.n770 B.n769 585
R365 B.n768 B.n767 585
R366 B.n766 B.n765 585
R367 B.n764 B.n763 585
R368 B.n762 B.n761 585
R369 B.n760 B.n759 585
R370 B.n758 B.n757 585
R371 B.n756 B.n755 585
R372 B.n754 B.n753 585
R373 B.n752 B.n751 585
R374 B.n750 B.n749 585
R375 B.n748 B.n747 585
R376 B.n746 B.n745 585
R377 B.n744 B.n743 585
R378 B.n742 B.n741 585
R379 B.n740 B.n739 585
R380 B.n738 B.n737 585
R381 B.n736 B.n735 585
R382 B.n734 B.n733 585
R383 B.n732 B.n731 585
R384 B.n730 B.n729 585
R385 B.n728 B.n727 585
R386 B.n726 B.n725 585
R387 B.n724 B.n723 585
R388 B.n722 B.n721 585
R389 B.n720 B.n719 585
R390 B.n718 B.n717 585
R391 B.n716 B.n715 585
R392 B.n714 B.n713 585
R393 B.n712 B.n711 585
R394 B.n710 B.n709 585
R395 B.n708 B.n707 585
R396 B.n706 B.n705 585
R397 B.n704 B.n703 585
R398 B.n702 B.n701 585
R399 B.n700 B.n699 585
R400 B.n698 B.n697 585
R401 B.n696 B.n695 585
R402 B.n694 B.n693 585
R403 B.n692 B.n691 585
R404 B.n690 B.n689 585
R405 B.n688 B.n687 585
R406 B.n686 B.n685 585
R407 B.n684 B.n683 585
R408 B.n682 B.n681 585
R409 B.n680 B.n679 585
R410 B.n678 B.n677 585
R411 B.n676 B.n675 585
R412 B.n674 B.n673 585
R413 B.n672 B.n671 585
R414 B.n670 B.n669 585
R415 B.n668 B.n667 585
R416 B.n666 B.n665 585
R417 B.n664 B.n663 585
R418 B.n662 B.n661 585
R419 B.n660 B.n659 585
R420 B.n658 B.n657 585
R421 B.n656 B.n655 585
R422 B.n654 B.n653 585
R423 B.n652 B.n651 585
R424 B.n650 B.n649 585
R425 B.n648 B.n647 585
R426 B.n646 B.n645 585
R427 B.n644 B.n643 585
R428 B.n641 B.n640 585
R429 B.n639 B.n638 585
R430 B.n637 B.n636 585
R431 B.n635 B.n634 585
R432 B.n633 B.n632 585
R433 B.n631 B.n630 585
R434 B.n629 B.n628 585
R435 B.n627 B.n626 585
R436 B.n625 B.n624 585
R437 B.n623 B.n622 585
R438 B.n621 B.n620 585
R439 B.n619 B.n618 585
R440 B.n617 B.n616 585
R441 B.n615 B.n614 585
R442 B.n613 B.n612 585
R443 B.n611 B.n610 585
R444 B.n609 B.n608 585
R445 B.n607 B.n606 585
R446 B.n605 B.n604 585
R447 B.n603 B.n602 585
R448 B.n601 B.n600 585
R449 B.n599 B.n598 585
R450 B.n597 B.n596 585
R451 B.n595 B.n594 585
R452 B.n593 B.n592 585
R453 B.n591 B.n590 585
R454 B.n589 B.n588 585
R455 B.n587 B.n586 585
R456 B.n585 B.n584 585
R457 B.n583 B.n582 585
R458 B.n581 B.n580 585
R459 B.n579 B.n578 585
R460 B.n577 B.n576 585
R461 B.n575 B.n574 585
R462 B.n573 B.n572 585
R463 B.n571 B.n570 585
R464 B.n569 B.n568 585
R465 B.n567 B.n566 585
R466 B.n565 B.n564 585
R467 B.n563 B.n562 585
R468 B.n561 B.n560 585
R469 B.n559 B.n558 585
R470 B.n557 B.n556 585
R471 B.n555 B.n554 585
R472 B.n553 B.n552 585
R473 B.n551 B.n550 585
R474 B.n549 B.n548 585
R475 B.n547 B.n546 585
R476 B.n545 B.n544 585
R477 B.n543 B.n542 585
R478 B.n541 B.n540 585
R479 B.n539 B.n538 585
R480 B.n537 B.n536 585
R481 B.n535 B.n534 585
R482 B.n533 B.n532 585
R483 B.n531 B.n530 585
R484 B.n529 B.n528 585
R485 B.n527 B.n526 585
R486 B.n525 B.n524 585
R487 B.n523 B.n522 585
R488 B.n521 B.n520 585
R489 B.n519 B.n518 585
R490 B.n517 B.n516 585
R491 B.n786 B.n441 585
R492 B.n441 B.n440 585
R493 B.n788 B.n787 585
R494 B.n789 B.n788 585
R495 B.n435 B.n434 585
R496 B.n436 B.n435 585
R497 B.n798 B.n797 585
R498 B.n797 B.n796 585
R499 B.n799 B.n433 585
R500 B.n795 B.n433 585
R501 B.n801 B.n800 585
R502 B.n802 B.n801 585
R503 B.n428 B.n427 585
R504 B.n429 B.n428 585
R505 B.n810 B.n809 585
R506 B.n809 B.n808 585
R507 B.n811 B.n426 585
R508 B.n426 B.n425 585
R509 B.n813 B.n812 585
R510 B.n814 B.n813 585
R511 B.n420 B.n419 585
R512 B.n421 B.n420 585
R513 B.n822 B.n821 585
R514 B.n821 B.n820 585
R515 B.n823 B.n418 585
R516 B.n418 B.n416 585
R517 B.n825 B.n824 585
R518 B.n826 B.n825 585
R519 B.n412 B.n411 585
R520 B.n417 B.n412 585
R521 B.n834 B.n833 585
R522 B.n833 B.n832 585
R523 B.n835 B.n410 585
R524 B.n410 B.n409 585
R525 B.n837 B.n836 585
R526 B.n838 B.n837 585
R527 B.n404 B.n403 585
R528 B.n405 B.n404 585
R529 B.n846 B.n845 585
R530 B.n845 B.n844 585
R531 B.n847 B.n402 585
R532 B.n402 B.n401 585
R533 B.n849 B.n848 585
R534 B.t2 B.n849 585
R535 B.n396 B.n395 585
R536 B.n397 B.n396 585
R537 B.n859 B.n858 585
R538 B.n858 B.n857 585
R539 B.n860 B.n394 585
R540 B.n856 B.n394 585
R541 B.n862 B.n861 585
R542 B.n863 B.n862 585
R543 B.n3 B.n0 585
R544 B.n4 B.n3 585
R545 B.n959 B.n1 585
R546 B.n960 B.n959 585
R547 B.n958 B.n957 585
R548 B.n958 B.n8 585
R549 B.n956 B.n9 585
R550 B.n12 B.n9 585
R551 B.n955 B.n954 585
R552 B.n954 B.n953 585
R553 B.n11 B.n10 585
R554 B.n952 B.n11 585
R555 B.n951 B.n950 585
R556 B.t8 B.n951 585
R557 B.n949 B.n17 585
R558 B.n17 B.n16 585
R559 B.n948 B.n947 585
R560 B.n947 B.n946 585
R561 B.n19 B.n18 585
R562 B.n945 B.n19 585
R563 B.n943 B.n942 585
R564 B.n944 B.n943 585
R565 B.n941 B.n24 585
R566 B.n24 B.n23 585
R567 B.n940 B.n939 585
R568 B.n939 B.n938 585
R569 B.n26 B.n25 585
R570 B.n937 B.n26 585
R571 B.n935 B.n934 585
R572 B.n936 B.n935 585
R573 B.n933 B.n31 585
R574 B.n31 B.n30 585
R575 B.n932 B.n931 585
R576 B.n931 B.n930 585
R577 B.n33 B.n32 585
R578 B.n929 B.n33 585
R579 B.n927 B.n926 585
R580 B.n928 B.n927 585
R581 B.n925 B.n38 585
R582 B.n38 B.n37 585
R583 B.n924 B.n923 585
R584 B.n923 B.n922 585
R585 B.n40 B.n39 585
R586 B.n921 B.n40 585
R587 B.n919 B.n918 585
R588 B.n920 B.n919 585
R589 B.n917 B.n44 585
R590 B.n47 B.n44 585
R591 B.n916 B.n915 585
R592 B.n915 B.n914 585
R593 B.n46 B.n45 585
R594 B.n913 B.n46 585
R595 B.n911 B.n910 585
R596 B.n912 B.n911 585
R597 B.n909 B.n52 585
R598 B.n52 B.n51 585
R599 B.n963 B.n962 585
R600 B.n961 B.n2 585
R601 B.n907 B.n52 564.573
R602 B.n904 B.n122 564.573
R603 B.n516 B.n439 564.573
R604 B.n784 B.n441 564.573
R605 B.n905 B.n120 256.663
R606 B.n905 B.n119 256.663
R607 B.n905 B.n118 256.663
R608 B.n905 B.n117 256.663
R609 B.n905 B.n116 256.663
R610 B.n905 B.n115 256.663
R611 B.n905 B.n114 256.663
R612 B.n905 B.n113 256.663
R613 B.n905 B.n112 256.663
R614 B.n905 B.n111 256.663
R615 B.n905 B.n110 256.663
R616 B.n905 B.n109 256.663
R617 B.n905 B.n108 256.663
R618 B.n905 B.n107 256.663
R619 B.n905 B.n106 256.663
R620 B.n905 B.n105 256.663
R621 B.n905 B.n104 256.663
R622 B.n905 B.n103 256.663
R623 B.n905 B.n102 256.663
R624 B.n905 B.n101 256.663
R625 B.n905 B.n100 256.663
R626 B.n905 B.n99 256.663
R627 B.n905 B.n98 256.663
R628 B.n905 B.n97 256.663
R629 B.n905 B.n96 256.663
R630 B.n905 B.n95 256.663
R631 B.n905 B.n94 256.663
R632 B.n905 B.n93 256.663
R633 B.n905 B.n92 256.663
R634 B.n905 B.n91 256.663
R635 B.n905 B.n90 256.663
R636 B.n905 B.n89 256.663
R637 B.n905 B.n88 256.663
R638 B.n905 B.n87 256.663
R639 B.n905 B.n86 256.663
R640 B.n905 B.n85 256.663
R641 B.n905 B.n84 256.663
R642 B.n905 B.n83 256.663
R643 B.n905 B.n82 256.663
R644 B.n905 B.n81 256.663
R645 B.n905 B.n80 256.663
R646 B.n905 B.n79 256.663
R647 B.n905 B.n78 256.663
R648 B.n905 B.n77 256.663
R649 B.n905 B.n76 256.663
R650 B.n905 B.n75 256.663
R651 B.n905 B.n74 256.663
R652 B.n905 B.n73 256.663
R653 B.n905 B.n72 256.663
R654 B.n905 B.n71 256.663
R655 B.n905 B.n70 256.663
R656 B.n905 B.n69 256.663
R657 B.n905 B.n68 256.663
R658 B.n905 B.n67 256.663
R659 B.n905 B.n66 256.663
R660 B.n905 B.n65 256.663
R661 B.n905 B.n64 256.663
R662 B.n905 B.n63 256.663
R663 B.n905 B.n62 256.663
R664 B.n905 B.n61 256.663
R665 B.n905 B.n60 256.663
R666 B.n905 B.n59 256.663
R667 B.n905 B.n58 256.663
R668 B.n905 B.n57 256.663
R669 B.n905 B.n56 256.663
R670 B.n905 B.n55 256.663
R671 B.n906 B.n905 256.663
R672 B.n783 B.n782 256.663
R673 B.n782 B.n444 256.663
R674 B.n782 B.n445 256.663
R675 B.n782 B.n446 256.663
R676 B.n782 B.n447 256.663
R677 B.n782 B.n448 256.663
R678 B.n782 B.n449 256.663
R679 B.n782 B.n450 256.663
R680 B.n782 B.n451 256.663
R681 B.n782 B.n452 256.663
R682 B.n782 B.n453 256.663
R683 B.n782 B.n454 256.663
R684 B.n782 B.n455 256.663
R685 B.n782 B.n456 256.663
R686 B.n782 B.n457 256.663
R687 B.n782 B.n458 256.663
R688 B.n782 B.n459 256.663
R689 B.n782 B.n460 256.663
R690 B.n782 B.n461 256.663
R691 B.n782 B.n462 256.663
R692 B.n782 B.n463 256.663
R693 B.n782 B.n464 256.663
R694 B.n782 B.n465 256.663
R695 B.n782 B.n466 256.663
R696 B.n782 B.n467 256.663
R697 B.n782 B.n468 256.663
R698 B.n782 B.n469 256.663
R699 B.n782 B.n470 256.663
R700 B.n782 B.n471 256.663
R701 B.n782 B.n472 256.663
R702 B.n782 B.n473 256.663
R703 B.n782 B.n474 256.663
R704 B.n782 B.n475 256.663
R705 B.n782 B.n476 256.663
R706 B.n782 B.n477 256.663
R707 B.n782 B.n478 256.663
R708 B.n782 B.n479 256.663
R709 B.n782 B.n480 256.663
R710 B.n782 B.n481 256.663
R711 B.n782 B.n482 256.663
R712 B.n782 B.n483 256.663
R713 B.n782 B.n484 256.663
R714 B.n782 B.n485 256.663
R715 B.n782 B.n486 256.663
R716 B.n782 B.n487 256.663
R717 B.n782 B.n488 256.663
R718 B.n782 B.n489 256.663
R719 B.n782 B.n490 256.663
R720 B.n782 B.n491 256.663
R721 B.n782 B.n492 256.663
R722 B.n782 B.n493 256.663
R723 B.n782 B.n494 256.663
R724 B.n782 B.n495 256.663
R725 B.n782 B.n496 256.663
R726 B.n782 B.n497 256.663
R727 B.n782 B.n498 256.663
R728 B.n782 B.n499 256.663
R729 B.n782 B.n500 256.663
R730 B.n782 B.n501 256.663
R731 B.n782 B.n502 256.663
R732 B.n782 B.n503 256.663
R733 B.n782 B.n504 256.663
R734 B.n782 B.n505 256.663
R735 B.n782 B.n506 256.663
R736 B.n782 B.n507 256.663
R737 B.n782 B.n508 256.663
R738 B.n782 B.n509 256.663
R739 B.n965 B.n964 256.663
R740 B.n128 B.n54 163.367
R741 B.n132 B.n131 163.367
R742 B.n136 B.n135 163.367
R743 B.n140 B.n139 163.367
R744 B.n144 B.n143 163.367
R745 B.n148 B.n147 163.367
R746 B.n152 B.n151 163.367
R747 B.n156 B.n155 163.367
R748 B.n160 B.n159 163.367
R749 B.n164 B.n163 163.367
R750 B.n168 B.n167 163.367
R751 B.n172 B.n171 163.367
R752 B.n176 B.n175 163.367
R753 B.n180 B.n179 163.367
R754 B.n184 B.n183 163.367
R755 B.n188 B.n187 163.367
R756 B.n192 B.n191 163.367
R757 B.n196 B.n195 163.367
R758 B.n200 B.n199 163.367
R759 B.n204 B.n203 163.367
R760 B.n208 B.n207 163.367
R761 B.n212 B.n211 163.367
R762 B.n216 B.n215 163.367
R763 B.n220 B.n219 163.367
R764 B.n224 B.n223 163.367
R765 B.n228 B.n227 163.367
R766 B.n232 B.n231 163.367
R767 B.n236 B.n235 163.367
R768 B.n240 B.n239 163.367
R769 B.n244 B.n243 163.367
R770 B.n248 B.n247 163.367
R771 B.n253 B.n252 163.367
R772 B.n257 B.n256 163.367
R773 B.n261 B.n260 163.367
R774 B.n265 B.n264 163.367
R775 B.n269 B.n268 163.367
R776 B.n273 B.n272 163.367
R777 B.n277 B.n276 163.367
R778 B.n281 B.n280 163.367
R779 B.n285 B.n284 163.367
R780 B.n289 B.n288 163.367
R781 B.n293 B.n292 163.367
R782 B.n297 B.n296 163.367
R783 B.n301 B.n300 163.367
R784 B.n305 B.n304 163.367
R785 B.n309 B.n308 163.367
R786 B.n313 B.n312 163.367
R787 B.n317 B.n316 163.367
R788 B.n321 B.n320 163.367
R789 B.n325 B.n324 163.367
R790 B.n329 B.n328 163.367
R791 B.n333 B.n332 163.367
R792 B.n337 B.n336 163.367
R793 B.n341 B.n340 163.367
R794 B.n345 B.n344 163.367
R795 B.n349 B.n348 163.367
R796 B.n353 B.n352 163.367
R797 B.n357 B.n356 163.367
R798 B.n361 B.n360 163.367
R799 B.n365 B.n364 163.367
R800 B.n369 B.n368 163.367
R801 B.n373 B.n372 163.367
R802 B.n377 B.n376 163.367
R803 B.n381 B.n380 163.367
R804 B.n385 B.n384 163.367
R805 B.n389 B.n388 163.367
R806 B.n904 B.n121 163.367
R807 B.n790 B.n439 163.367
R808 B.n790 B.n437 163.367
R809 B.n794 B.n437 163.367
R810 B.n794 B.n432 163.367
R811 B.n803 B.n432 163.367
R812 B.n803 B.n430 163.367
R813 B.n807 B.n430 163.367
R814 B.n807 B.n424 163.367
R815 B.n815 B.n424 163.367
R816 B.n815 B.n422 163.367
R817 B.n819 B.n422 163.367
R818 B.n819 B.n415 163.367
R819 B.n827 B.n415 163.367
R820 B.n827 B.n413 163.367
R821 B.n831 B.n413 163.367
R822 B.n831 B.n408 163.367
R823 B.n839 B.n408 163.367
R824 B.n839 B.n406 163.367
R825 B.n843 B.n406 163.367
R826 B.n843 B.n400 163.367
R827 B.n850 B.n400 163.367
R828 B.n850 B.n398 163.367
R829 B.n855 B.n398 163.367
R830 B.n855 B.n393 163.367
R831 B.n864 B.n393 163.367
R832 B.n865 B.n864 163.367
R833 B.n865 B.n5 163.367
R834 B.n6 B.n5 163.367
R835 B.n7 B.n6 163.367
R836 B.n871 B.n7 163.367
R837 B.n872 B.n871 163.367
R838 B.n872 B.n13 163.367
R839 B.n14 B.n13 163.367
R840 B.n15 B.n14 163.367
R841 B.n877 B.n15 163.367
R842 B.n877 B.n20 163.367
R843 B.n21 B.n20 163.367
R844 B.n22 B.n21 163.367
R845 B.n882 B.n22 163.367
R846 B.n882 B.n27 163.367
R847 B.n28 B.n27 163.367
R848 B.n29 B.n28 163.367
R849 B.n887 B.n29 163.367
R850 B.n887 B.n34 163.367
R851 B.n35 B.n34 163.367
R852 B.n36 B.n35 163.367
R853 B.n892 B.n36 163.367
R854 B.n892 B.n41 163.367
R855 B.n42 B.n41 163.367
R856 B.n43 B.n42 163.367
R857 B.n897 B.n43 163.367
R858 B.n897 B.n48 163.367
R859 B.n49 B.n48 163.367
R860 B.n50 B.n49 163.367
R861 B.n122 B.n50 163.367
R862 B.n781 B.n443 163.367
R863 B.n781 B.n510 163.367
R864 B.n777 B.n776 163.367
R865 B.n773 B.n772 163.367
R866 B.n769 B.n768 163.367
R867 B.n765 B.n764 163.367
R868 B.n761 B.n760 163.367
R869 B.n757 B.n756 163.367
R870 B.n753 B.n752 163.367
R871 B.n749 B.n748 163.367
R872 B.n745 B.n744 163.367
R873 B.n741 B.n740 163.367
R874 B.n737 B.n736 163.367
R875 B.n733 B.n732 163.367
R876 B.n729 B.n728 163.367
R877 B.n725 B.n724 163.367
R878 B.n721 B.n720 163.367
R879 B.n717 B.n716 163.367
R880 B.n713 B.n712 163.367
R881 B.n709 B.n708 163.367
R882 B.n705 B.n704 163.367
R883 B.n701 B.n700 163.367
R884 B.n697 B.n696 163.367
R885 B.n693 B.n692 163.367
R886 B.n689 B.n688 163.367
R887 B.n685 B.n684 163.367
R888 B.n681 B.n680 163.367
R889 B.n677 B.n676 163.367
R890 B.n673 B.n672 163.367
R891 B.n669 B.n668 163.367
R892 B.n665 B.n664 163.367
R893 B.n661 B.n660 163.367
R894 B.n657 B.n656 163.367
R895 B.n653 B.n652 163.367
R896 B.n649 B.n648 163.367
R897 B.n645 B.n644 163.367
R898 B.n640 B.n639 163.367
R899 B.n636 B.n635 163.367
R900 B.n632 B.n631 163.367
R901 B.n628 B.n627 163.367
R902 B.n624 B.n623 163.367
R903 B.n620 B.n619 163.367
R904 B.n616 B.n615 163.367
R905 B.n612 B.n611 163.367
R906 B.n608 B.n607 163.367
R907 B.n604 B.n603 163.367
R908 B.n600 B.n599 163.367
R909 B.n596 B.n595 163.367
R910 B.n592 B.n591 163.367
R911 B.n588 B.n587 163.367
R912 B.n584 B.n583 163.367
R913 B.n580 B.n579 163.367
R914 B.n576 B.n575 163.367
R915 B.n572 B.n571 163.367
R916 B.n568 B.n567 163.367
R917 B.n564 B.n563 163.367
R918 B.n560 B.n559 163.367
R919 B.n556 B.n555 163.367
R920 B.n552 B.n551 163.367
R921 B.n548 B.n547 163.367
R922 B.n544 B.n543 163.367
R923 B.n540 B.n539 163.367
R924 B.n536 B.n535 163.367
R925 B.n532 B.n531 163.367
R926 B.n528 B.n527 163.367
R927 B.n524 B.n523 163.367
R928 B.n520 B.n519 163.367
R929 B.n788 B.n441 163.367
R930 B.n788 B.n435 163.367
R931 B.n797 B.n435 163.367
R932 B.n797 B.n433 163.367
R933 B.n801 B.n433 163.367
R934 B.n801 B.n428 163.367
R935 B.n809 B.n428 163.367
R936 B.n809 B.n426 163.367
R937 B.n813 B.n426 163.367
R938 B.n813 B.n420 163.367
R939 B.n821 B.n420 163.367
R940 B.n821 B.n418 163.367
R941 B.n825 B.n418 163.367
R942 B.n825 B.n412 163.367
R943 B.n833 B.n412 163.367
R944 B.n833 B.n410 163.367
R945 B.n837 B.n410 163.367
R946 B.n837 B.n404 163.367
R947 B.n845 B.n404 163.367
R948 B.n845 B.n402 163.367
R949 B.n849 B.n402 163.367
R950 B.n849 B.n396 163.367
R951 B.n858 B.n396 163.367
R952 B.n858 B.n394 163.367
R953 B.n862 B.n394 163.367
R954 B.n862 B.n3 163.367
R955 B.n963 B.n3 163.367
R956 B.n959 B.n2 163.367
R957 B.n959 B.n958 163.367
R958 B.n958 B.n9 163.367
R959 B.n954 B.n9 163.367
R960 B.n954 B.n11 163.367
R961 B.n951 B.n11 163.367
R962 B.n951 B.n17 163.367
R963 B.n947 B.n17 163.367
R964 B.n947 B.n19 163.367
R965 B.n943 B.n19 163.367
R966 B.n943 B.n24 163.367
R967 B.n939 B.n24 163.367
R968 B.n939 B.n26 163.367
R969 B.n935 B.n26 163.367
R970 B.n935 B.n31 163.367
R971 B.n931 B.n31 163.367
R972 B.n931 B.n33 163.367
R973 B.n927 B.n33 163.367
R974 B.n927 B.n38 163.367
R975 B.n923 B.n38 163.367
R976 B.n923 B.n40 163.367
R977 B.n919 B.n40 163.367
R978 B.n919 B.n44 163.367
R979 B.n915 B.n44 163.367
R980 B.n915 B.n46 163.367
R981 B.n911 B.n46 163.367
R982 B.n911 B.n52 163.367
R983 B.n123 B.t19 92.5856
R984 B.n514 B.t13 92.5856
R985 B.n126 B.t22 92.5598
R986 B.n511 B.t16 92.5598
R987 B.n907 B.n906 71.676
R988 B.n128 B.n55 71.676
R989 B.n132 B.n56 71.676
R990 B.n136 B.n57 71.676
R991 B.n140 B.n58 71.676
R992 B.n144 B.n59 71.676
R993 B.n148 B.n60 71.676
R994 B.n152 B.n61 71.676
R995 B.n156 B.n62 71.676
R996 B.n160 B.n63 71.676
R997 B.n164 B.n64 71.676
R998 B.n168 B.n65 71.676
R999 B.n172 B.n66 71.676
R1000 B.n176 B.n67 71.676
R1001 B.n180 B.n68 71.676
R1002 B.n184 B.n69 71.676
R1003 B.n188 B.n70 71.676
R1004 B.n192 B.n71 71.676
R1005 B.n196 B.n72 71.676
R1006 B.n200 B.n73 71.676
R1007 B.n204 B.n74 71.676
R1008 B.n208 B.n75 71.676
R1009 B.n212 B.n76 71.676
R1010 B.n216 B.n77 71.676
R1011 B.n220 B.n78 71.676
R1012 B.n224 B.n79 71.676
R1013 B.n228 B.n80 71.676
R1014 B.n232 B.n81 71.676
R1015 B.n236 B.n82 71.676
R1016 B.n240 B.n83 71.676
R1017 B.n244 B.n84 71.676
R1018 B.n248 B.n85 71.676
R1019 B.n253 B.n86 71.676
R1020 B.n257 B.n87 71.676
R1021 B.n261 B.n88 71.676
R1022 B.n265 B.n89 71.676
R1023 B.n269 B.n90 71.676
R1024 B.n273 B.n91 71.676
R1025 B.n277 B.n92 71.676
R1026 B.n281 B.n93 71.676
R1027 B.n285 B.n94 71.676
R1028 B.n289 B.n95 71.676
R1029 B.n293 B.n96 71.676
R1030 B.n297 B.n97 71.676
R1031 B.n301 B.n98 71.676
R1032 B.n305 B.n99 71.676
R1033 B.n309 B.n100 71.676
R1034 B.n313 B.n101 71.676
R1035 B.n317 B.n102 71.676
R1036 B.n321 B.n103 71.676
R1037 B.n325 B.n104 71.676
R1038 B.n329 B.n105 71.676
R1039 B.n333 B.n106 71.676
R1040 B.n337 B.n107 71.676
R1041 B.n341 B.n108 71.676
R1042 B.n345 B.n109 71.676
R1043 B.n349 B.n110 71.676
R1044 B.n353 B.n111 71.676
R1045 B.n357 B.n112 71.676
R1046 B.n361 B.n113 71.676
R1047 B.n365 B.n114 71.676
R1048 B.n369 B.n115 71.676
R1049 B.n373 B.n116 71.676
R1050 B.n377 B.n117 71.676
R1051 B.n381 B.n118 71.676
R1052 B.n385 B.n119 71.676
R1053 B.n389 B.n120 71.676
R1054 B.n121 B.n120 71.676
R1055 B.n388 B.n119 71.676
R1056 B.n384 B.n118 71.676
R1057 B.n380 B.n117 71.676
R1058 B.n376 B.n116 71.676
R1059 B.n372 B.n115 71.676
R1060 B.n368 B.n114 71.676
R1061 B.n364 B.n113 71.676
R1062 B.n360 B.n112 71.676
R1063 B.n356 B.n111 71.676
R1064 B.n352 B.n110 71.676
R1065 B.n348 B.n109 71.676
R1066 B.n344 B.n108 71.676
R1067 B.n340 B.n107 71.676
R1068 B.n336 B.n106 71.676
R1069 B.n332 B.n105 71.676
R1070 B.n328 B.n104 71.676
R1071 B.n324 B.n103 71.676
R1072 B.n320 B.n102 71.676
R1073 B.n316 B.n101 71.676
R1074 B.n312 B.n100 71.676
R1075 B.n308 B.n99 71.676
R1076 B.n304 B.n98 71.676
R1077 B.n300 B.n97 71.676
R1078 B.n296 B.n96 71.676
R1079 B.n292 B.n95 71.676
R1080 B.n288 B.n94 71.676
R1081 B.n284 B.n93 71.676
R1082 B.n280 B.n92 71.676
R1083 B.n276 B.n91 71.676
R1084 B.n272 B.n90 71.676
R1085 B.n268 B.n89 71.676
R1086 B.n264 B.n88 71.676
R1087 B.n260 B.n87 71.676
R1088 B.n256 B.n86 71.676
R1089 B.n252 B.n85 71.676
R1090 B.n247 B.n84 71.676
R1091 B.n243 B.n83 71.676
R1092 B.n239 B.n82 71.676
R1093 B.n235 B.n81 71.676
R1094 B.n231 B.n80 71.676
R1095 B.n227 B.n79 71.676
R1096 B.n223 B.n78 71.676
R1097 B.n219 B.n77 71.676
R1098 B.n215 B.n76 71.676
R1099 B.n211 B.n75 71.676
R1100 B.n207 B.n74 71.676
R1101 B.n203 B.n73 71.676
R1102 B.n199 B.n72 71.676
R1103 B.n195 B.n71 71.676
R1104 B.n191 B.n70 71.676
R1105 B.n187 B.n69 71.676
R1106 B.n183 B.n68 71.676
R1107 B.n179 B.n67 71.676
R1108 B.n175 B.n66 71.676
R1109 B.n171 B.n65 71.676
R1110 B.n167 B.n64 71.676
R1111 B.n163 B.n63 71.676
R1112 B.n159 B.n62 71.676
R1113 B.n155 B.n61 71.676
R1114 B.n151 B.n60 71.676
R1115 B.n147 B.n59 71.676
R1116 B.n143 B.n58 71.676
R1117 B.n139 B.n57 71.676
R1118 B.n135 B.n56 71.676
R1119 B.n131 B.n55 71.676
R1120 B.n906 B.n54 71.676
R1121 B.n784 B.n783 71.676
R1122 B.n510 B.n444 71.676
R1123 B.n776 B.n445 71.676
R1124 B.n772 B.n446 71.676
R1125 B.n768 B.n447 71.676
R1126 B.n764 B.n448 71.676
R1127 B.n760 B.n449 71.676
R1128 B.n756 B.n450 71.676
R1129 B.n752 B.n451 71.676
R1130 B.n748 B.n452 71.676
R1131 B.n744 B.n453 71.676
R1132 B.n740 B.n454 71.676
R1133 B.n736 B.n455 71.676
R1134 B.n732 B.n456 71.676
R1135 B.n728 B.n457 71.676
R1136 B.n724 B.n458 71.676
R1137 B.n720 B.n459 71.676
R1138 B.n716 B.n460 71.676
R1139 B.n712 B.n461 71.676
R1140 B.n708 B.n462 71.676
R1141 B.n704 B.n463 71.676
R1142 B.n700 B.n464 71.676
R1143 B.n696 B.n465 71.676
R1144 B.n692 B.n466 71.676
R1145 B.n688 B.n467 71.676
R1146 B.n684 B.n468 71.676
R1147 B.n680 B.n469 71.676
R1148 B.n676 B.n470 71.676
R1149 B.n672 B.n471 71.676
R1150 B.n668 B.n472 71.676
R1151 B.n664 B.n473 71.676
R1152 B.n660 B.n474 71.676
R1153 B.n656 B.n475 71.676
R1154 B.n652 B.n476 71.676
R1155 B.n648 B.n477 71.676
R1156 B.n644 B.n478 71.676
R1157 B.n639 B.n479 71.676
R1158 B.n635 B.n480 71.676
R1159 B.n631 B.n481 71.676
R1160 B.n627 B.n482 71.676
R1161 B.n623 B.n483 71.676
R1162 B.n619 B.n484 71.676
R1163 B.n615 B.n485 71.676
R1164 B.n611 B.n486 71.676
R1165 B.n607 B.n487 71.676
R1166 B.n603 B.n488 71.676
R1167 B.n599 B.n489 71.676
R1168 B.n595 B.n490 71.676
R1169 B.n591 B.n491 71.676
R1170 B.n587 B.n492 71.676
R1171 B.n583 B.n493 71.676
R1172 B.n579 B.n494 71.676
R1173 B.n575 B.n495 71.676
R1174 B.n571 B.n496 71.676
R1175 B.n567 B.n497 71.676
R1176 B.n563 B.n498 71.676
R1177 B.n559 B.n499 71.676
R1178 B.n555 B.n500 71.676
R1179 B.n551 B.n501 71.676
R1180 B.n547 B.n502 71.676
R1181 B.n543 B.n503 71.676
R1182 B.n539 B.n504 71.676
R1183 B.n535 B.n505 71.676
R1184 B.n531 B.n506 71.676
R1185 B.n527 B.n507 71.676
R1186 B.n523 B.n508 71.676
R1187 B.n519 B.n509 71.676
R1188 B.n783 B.n443 71.676
R1189 B.n777 B.n444 71.676
R1190 B.n773 B.n445 71.676
R1191 B.n769 B.n446 71.676
R1192 B.n765 B.n447 71.676
R1193 B.n761 B.n448 71.676
R1194 B.n757 B.n449 71.676
R1195 B.n753 B.n450 71.676
R1196 B.n749 B.n451 71.676
R1197 B.n745 B.n452 71.676
R1198 B.n741 B.n453 71.676
R1199 B.n737 B.n454 71.676
R1200 B.n733 B.n455 71.676
R1201 B.n729 B.n456 71.676
R1202 B.n725 B.n457 71.676
R1203 B.n721 B.n458 71.676
R1204 B.n717 B.n459 71.676
R1205 B.n713 B.n460 71.676
R1206 B.n709 B.n461 71.676
R1207 B.n705 B.n462 71.676
R1208 B.n701 B.n463 71.676
R1209 B.n697 B.n464 71.676
R1210 B.n693 B.n465 71.676
R1211 B.n689 B.n466 71.676
R1212 B.n685 B.n467 71.676
R1213 B.n681 B.n468 71.676
R1214 B.n677 B.n469 71.676
R1215 B.n673 B.n470 71.676
R1216 B.n669 B.n471 71.676
R1217 B.n665 B.n472 71.676
R1218 B.n661 B.n473 71.676
R1219 B.n657 B.n474 71.676
R1220 B.n653 B.n475 71.676
R1221 B.n649 B.n476 71.676
R1222 B.n645 B.n477 71.676
R1223 B.n640 B.n478 71.676
R1224 B.n636 B.n479 71.676
R1225 B.n632 B.n480 71.676
R1226 B.n628 B.n481 71.676
R1227 B.n624 B.n482 71.676
R1228 B.n620 B.n483 71.676
R1229 B.n616 B.n484 71.676
R1230 B.n612 B.n485 71.676
R1231 B.n608 B.n486 71.676
R1232 B.n604 B.n487 71.676
R1233 B.n600 B.n488 71.676
R1234 B.n596 B.n489 71.676
R1235 B.n592 B.n490 71.676
R1236 B.n588 B.n491 71.676
R1237 B.n584 B.n492 71.676
R1238 B.n580 B.n493 71.676
R1239 B.n576 B.n494 71.676
R1240 B.n572 B.n495 71.676
R1241 B.n568 B.n496 71.676
R1242 B.n564 B.n497 71.676
R1243 B.n560 B.n498 71.676
R1244 B.n556 B.n499 71.676
R1245 B.n552 B.n500 71.676
R1246 B.n548 B.n501 71.676
R1247 B.n544 B.n502 71.676
R1248 B.n540 B.n503 71.676
R1249 B.n536 B.n504 71.676
R1250 B.n532 B.n505 71.676
R1251 B.n528 B.n506 71.676
R1252 B.n524 B.n507 71.676
R1253 B.n520 B.n508 71.676
R1254 B.n516 B.n509 71.676
R1255 B.n964 B.n963 71.676
R1256 B.n964 B.n2 71.676
R1257 B.n124 B.t20 71.0583
R1258 B.n515 B.t12 71.0583
R1259 B.n127 B.t23 71.0326
R1260 B.n512 B.t15 71.0326
R1261 B.n782 B.n440 61.4731
R1262 B.n905 B.n51 61.4731
R1263 B.n250 B.n127 59.5399
R1264 B.n125 B.n124 59.5399
R1265 B.n642 B.n515 59.5399
R1266 B.n513 B.n512 59.5399
R1267 B.n786 B.n785 36.6834
R1268 B.n517 B.n438 36.6834
R1269 B.n903 B.n902 36.6834
R1270 B.n909 B.n908 36.6834
R1271 B.n789 B.n440 30.5124
R1272 B.n789 B.n436 30.5124
R1273 B.n796 B.n436 30.5124
R1274 B.n796 B.n795 30.5124
R1275 B.n802 B.n429 30.5124
R1276 B.n808 B.n429 30.5124
R1277 B.n808 B.n425 30.5124
R1278 B.n814 B.n425 30.5124
R1279 B.n814 B.n421 30.5124
R1280 B.n820 B.n421 30.5124
R1281 B.n826 B.n416 30.5124
R1282 B.n826 B.n417 30.5124
R1283 B.n832 B.n409 30.5124
R1284 B.n838 B.n409 30.5124
R1285 B.n844 B.n405 30.5124
R1286 B.n844 B.n401 30.5124
R1287 B.t2 B.n401 30.5124
R1288 B.t2 B.n397 30.5124
R1289 B.n857 B.n397 30.5124
R1290 B.n857 B.n856 30.5124
R1291 B.n863 B.n4 30.5124
R1292 B.n962 B.n4 30.5124
R1293 B.n962 B.n961 30.5124
R1294 B.n961 B.n960 30.5124
R1295 B.n960 B.n8 30.5124
R1296 B.n953 B.n12 30.5124
R1297 B.n953 B.n952 30.5124
R1298 B.n952 B.t8 30.5124
R1299 B.t8 B.n16 30.5124
R1300 B.n946 B.n16 30.5124
R1301 B.n946 B.n945 30.5124
R1302 B.n944 B.n23 30.5124
R1303 B.n938 B.n23 30.5124
R1304 B.n937 B.n936 30.5124
R1305 B.n936 B.n30 30.5124
R1306 B.n930 B.n929 30.5124
R1307 B.n929 B.n928 30.5124
R1308 B.n928 B.n37 30.5124
R1309 B.n922 B.n37 30.5124
R1310 B.n922 B.n921 30.5124
R1311 B.n921 B.n920 30.5124
R1312 B.n914 B.n47 30.5124
R1313 B.n914 B.n913 30.5124
R1314 B.n913 B.n912 30.5124
R1315 B.n912 B.n51 30.5124
R1316 B.t3 B.n416 24.2306
R1317 B.t1 B.n30 24.2306
R1318 B.n795 B.t11 22.4357
R1319 B.n838 B.t9 22.4357
R1320 B.n863 B.t7 22.4357
R1321 B.t4 B.n8 22.4357
R1322 B.t0 B.n944 22.4357
R1323 B.n47 B.t18 22.4357
R1324 B.n127 B.n126 21.5278
R1325 B.n124 B.n123 21.5278
R1326 B.n515 B.n514 21.5278
R1327 B.n512 B.n511 21.5278
R1328 B B.n965 18.0485
R1329 B.n832 B.t5 16.1539
R1330 B.n938 B.t6 16.1539
R1331 B.n417 B.t5 14.3591
R1332 B.t6 B.n937 14.3591
R1333 B.n787 B.n786 10.6151
R1334 B.n787 B.n434 10.6151
R1335 B.n798 B.n434 10.6151
R1336 B.n799 B.n798 10.6151
R1337 B.n800 B.n799 10.6151
R1338 B.n800 B.n427 10.6151
R1339 B.n810 B.n427 10.6151
R1340 B.n811 B.n810 10.6151
R1341 B.n812 B.n811 10.6151
R1342 B.n812 B.n419 10.6151
R1343 B.n822 B.n419 10.6151
R1344 B.n823 B.n822 10.6151
R1345 B.n824 B.n823 10.6151
R1346 B.n824 B.n411 10.6151
R1347 B.n834 B.n411 10.6151
R1348 B.n835 B.n834 10.6151
R1349 B.n836 B.n835 10.6151
R1350 B.n836 B.n403 10.6151
R1351 B.n846 B.n403 10.6151
R1352 B.n847 B.n846 10.6151
R1353 B.n848 B.n847 10.6151
R1354 B.n848 B.n395 10.6151
R1355 B.n859 B.n395 10.6151
R1356 B.n860 B.n859 10.6151
R1357 B.n861 B.n860 10.6151
R1358 B.n861 B.n0 10.6151
R1359 B.n785 B.n442 10.6151
R1360 B.n780 B.n442 10.6151
R1361 B.n780 B.n779 10.6151
R1362 B.n779 B.n778 10.6151
R1363 B.n778 B.n775 10.6151
R1364 B.n775 B.n774 10.6151
R1365 B.n774 B.n771 10.6151
R1366 B.n771 B.n770 10.6151
R1367 B.n770 B.n767 10.6151
R1368 B.n767 B.n766 10.6151
R1369 B.n766 B.n763 10.6151
R1370 B.n763 B.n762 10.6151
R1371 B.n762 B.n759 10.6151
R1372 B.n759 B.n758 10.6151
R1373 B.n758 B.n755 10.6151
R1374 B.n755 B.n754 10.6151
R1375 B.n754 B.n751 10.6151
R1376 B.n751 B.n750 10.6151
R1377 B.n750 B.n747 10.6151
R1378 B.n747 B.n746 10.6151
R1379 B.n746 B.n743 10.6151
R1380 B.n743 B.n742 10.6151
R1381 B.n742 B.n739 10.6151
R1382 B.n739 B.n738 10.6151
R1383 B.n738 B.n735 10.6151
R1384 B.n735 B.n734 10.6151
R1385 B.n734 B.n731 10.6151
R1386 B.n731 B.n730 10.6151
R1387 B.n730 B.n727 10.6151
R1388 B.n727 B.n726 10.6151
R1389 B.n726 B.n723 10.6151
R1390 B.n723 B.n722 10.6151
R1391 B.n722 B.n719 10.6151
R1392 B.n719 B.n718 10.6151
R1393 B.n718 B.n715 10.6151
R1394 B.n715 B.n714 10.6151
R1395 B.n714 B.n711 10.6151
R1396 B.n711 B.n710 10.6151
R1397 B.n710 B.n707 10.6151
R1398 B.n707 B.n706 10.6151
R1399 B.n706 B.n703 10.6151
R1400 B.n703 B.n702 10.6151
R1401 B.n702 B.n699 10.6151
R1402 B.n699 B.n698 10.6151
R1403 B.n698 B.n695 10.6151
R1404 B.n695 B.n694 10.6151
R1405 B.n694 B.n691 10.6151
R1406 B.n691 B.n690 10.6151
R1407 B.n690 B.n687 10.6151
R1408 B.n687 B.n686 10.6151
R1409 B.n686 B.n683 10.6151
R1410 B.n683 B.n682 10.6151
R1411 B.n682 B.n679 10.6151
R1412 B.n679 B.n678 10.6151
R1413 B.n678 B.n675 10.6151
R1414 B.n675 B.n674 10.6151
R1415 B.n674 B.n671 10.6151
R1416 B.n671 B.n670 10.6151
R1417 B.n670 B.n667 10.6151
R1418 B.n667 B.n666 10.6151
R1419 B.n666 B.n663 10.6151
R1420 B.n663 B.n662 10.6151
R1421 B.n659 B.n658 10.6151
R1422 B.n658 B.n655 10.6151
R1423 B.n655 B.n654 10.6151
R1424 B.n654 B.n651 10.6151
R1425 B.n651 B.n650 10.6151
R1426 B.n650 B.n647 10.6151
R1427 B.n647 B.n646 10.6151
R1428 B.n646 B.n643 10.6151
R1429 B.n641 B.n638 10.6151
R1430 B.n638 B.n637 10.6151
R1431 B.n637 B.n634 10.6151
R1432 B.n634 B.n633 10.6151
R1433 B.n633 B.n630 10.6151
R1434 B.n630 B.n629 10.6151
R1435 B.n629 B.n626 10.6151
R1436 B.n626 B.n625 10.6151
R1437 B.n625 B.n622 10.6151
R1438 B.n622 B.n621 10.6151
R1439 B.n621 B.n618 10.6151
R1440 B.n618 B.n617 10.6151
R1441 B.n617 B.n614 10.6151
R1442 B.n614 B.n613 10.6151
R1443 B.n613 B.n610 10.6151
R1444 B.n610 B.n609 10.6151
R1445 B.n609 B.n606 10.6151
R1446 B.n606 B.n605 10.6151
R1447 B.n605 B.n602 10.6151
R1448 B.n602 B.n601 10.6151
R1449 B.n601 B.n598 10.6151
R1450 B.n598 B.n597 10.6151
R1451 B.n597 B.n594 10.6151
R1452 B.n594 B.n593 10.6151
R1453 B.n593 B.n590 10.6151
R1454 B.n590 B.n589 10.6151
R1455 B.n589 B.n586 10.6151
R1456 B.n586 B.n585 10.6151
R1457 B.n585 B.n582 10.6151
R1458 B.n582 B.n581 10.6151
R1459 B.n581 B.n578 10.6151
R1460 B.n578 B.n577 10.6151
R1461 B.n577 B.n574 10.6151
R1462 B.n574 B.n573 10.6151
R1463 B.n573 B.n570 10.6151
R1464 B.n570 B.n569 10.6151
R1465 B.n569 B.n566 10.6151
R1466 B.n566 B.n565 10.6151
R1467 B.n565 B.n562 10.6151
R1468 B.n562 B.n561 10.6151
R1469 B.n561 B.n558 10.6151
R1470 B.n558 B.n557 10.6151
R1471 B.n557 B.n554 10.6151
R1472 B.n554 B.n553 10.6151
R1473 B.n553 B.n550 10.6151
R1474 B.n550 B.n549 10.6151
R1475 B.n549 B.n546 10.6151
R1476 B.n546 B.n545 10.6151
R1477 B.n545 B.n542 10.6151
R1478 B.n542 B.n541 10.6151
R1479 B.n541 B.n538 10.6151
R1480 B.n538 B.n537 10.6151
R1481 B.n537 B.n534 10.6151
R1482 B.n534 B.n533 10.6151
R1483 B.n533 B.n530 10.6151
R1484 B.n530 B.n529 10.6151
R1485 B.n529 B.n526 10.6151
R1486 B.n526 B.n525 10.6151
R1487 B.n525 B.n522 10.6151
R1488 B.n522 B.n521 10.6151
R1489 B.n521 B.n518 10.6151
R1490 B.n518 B.n517 10.6151
R1491 B.n791 B.n438 10.6151
R1492 B.n792 B.n791 10.6151
R1493 B.n793 B.n792 10.6151
R1494 B.n793 B.n431 10.6151
R1495 B.n804 B.n431 10.6151
R1496 B.n805 B.n804 10.6151
R1497 B.n806 B.n805 10.6151
R1498 B.n806 B.n423 10.6151
R1499 B.n816 B.n423 10.6151
R1500 B.n817 B.n816 10.6151
R1501 B.n818 B.n817 10.6151
R1502 B.n818 B.n414 10.6151
R1503 B.n828 B.n414 10.6151
R1504 B.n829 B.n828 10.6151
R1505 B.n830 B.n829 10.6151
R1506 B.n830 B.n407 10.6151
R1507 B.n840 B.n407 10.6151
R1508 B.n841 B.n840 10.6151
R1509 B.n842 B.n841 10.6151
R1510 B.n842 B.n399 10.6151
R1511 B.n851 B.n399 10.6151
R1512 B.n852 B.n851 10.6151
R1513 B.n854 B.n852 10.6151
R1514 B.n854 B.n853 10.6151
R1515 B.n853 B.n392 10.6151
R1516 B.n866 B.n392 10.6151
R1517 B.n867 B.n866 10.6151
R1518 B.n868 B.n867 10.6151
R1519 B.n869 B.n868 10.6151
R1520 B.n870 B.n869 10.6151
R1521 B.n873 B.n870 10.6151
R1522 B.n874 B.n873 10.6151
R1523 B.n875 B.n874 10.6151
R1524 B.n876 B.n875 10.6151
R1525 B.n878 B.n876 10.6151
R1526 B.n879 B.n878 10.6151
R1527 B.n880 B.n879 10.6151
R1528 B.n881 B.n880 10.6151
R1529 B.n883 B.n881 10.6151
R1530 B.n884 B.n883 10.6151
R1531 B.n885 B.n884 10.6151
R1532 B.n886 B.n885 10.6151
R1533 B.n888 B.n886 10.6151
R1534 B.n889 B.n888 10.6151
R1535 B.n890 B.n889 10.6151
R1536 B.n891 B.n890 10.6151
R1537 B.n893 B.n891 10.6151
R1538 B.n894 B.n893 10.6151
R1539 B.n895 B.n894 10.6151
R1540 B.n896 B.n895 10.6151
R1541 B.n898 B.n896 10.6151
R1542 B.n899 B.n898 10.6151
R1543 B.n900 B.n899 10.6151
R1544 B.n901 B.n900 10.6151
R1545 B.n902 B.n901 10.6151
R1546 B.n957 B.n1 10.6151
R1547 B.n957 B.n956 10.6151
R1548 B.n956 B.n955 10.6151
R1549 B.n955 B.n10 10.6151
R1550 B.n950 B.n10 10.6151
R1551 B.n950 B.n949 10.6151
R1552 B.n949 B.n948 10.6151
R1553 B.n948 B.n18 10.6151
R1554 B.n942 B.n18 10.6151
R1555 B.n942 B.n941 10.6151
R1556 B.n941 B.n940 10.6151
R1557 B.n940 B.n25 10.6151
R1558 B.n934 B.n25 10.6151
R1559 B.n934 B.n933 10.6151
R1560 B.n933 B.n932 10.6151
R1561 B.n932 B.n32 10.6151
R1562 B.n926 B.n32 10.6151
R1563 B.n926 B.n925 10.6151
R1564 B.n925 B.n924 10.6151
R1565 B.n924 B.n39 10.6151
R1566 B.n918 B.n39 10.6151
R1567 B.n918 B.n917 10.6151
R1568 B.n917 B.n916 10.6151
R1569 B.n916 B.n45 10.6151
R1570 B.n910 B.n45 10.6151
R1571 B.n910 B.n909 10.6151
R1572 B.n908 B.n53 10.6151
R1573 B.n129 B.n53 10.6151
R1574 B.n130 B.n129 10.6151
R1575 B.n133 B.n130 10.6151
R1576 B.n134 B.n133 10.6151
R1577 B.n137 B.n134 10.6151
R1578 B.n138 B.n137 10.6151
R1579 B.n141 B.n138 10.6151
R1580 B.n142 B.n141 10.6151
R1581 B.n145 B.n142 10.6151
R1582 B.n146 B.n145 10.6151
R1583 B.n149 B.n146 10.6151
R1584 B.n150 B.n149 10.6151
R1585 B.n153 B.n150 10.6151
R1586 B.n154 B.n153 10.6151
R1587 B.n157 B.n154 10.6151
R1588 B.n158 B.n157 10.6151
R1589 B.n161 B.n158 10.6151
R1590 B.n162 B.n161 10.6151
R1591 B.n165 B.n162 10.6151
R1592 B.n166 B.n165 10.6151
R1593 B.n169 B.n166 10.6151
R1594 B.n170 B.n169 10.6151
R1595 B.n173 B.n170 10.6151
R1596 B.n174 B.n173 10.6151
R1597 B.n177 B.n174 10.6151
R1598 B.n178 B.n177 10.6151
R1599 B.n181 B.n178 10.6151
R1600 B.n182 B.n181 10.6151
R1601 B.n185 B.n182 10.6151
R1602 B.n186 B.n185 10.6151
R1603 B.n189 B.n186 10.6151
R1604 B.n190 B.n189 10.6151
R1605 B.n193 B.n190 10.6151
R1606 B.n194 B.n193 10.6151
R1607 B.n197 B.n194 10.6151
R1608 B.n198 B.n197 10.6151
R1609 B.n201 B.n198 10.6151
R1610 B.n202 B.n201 10.6151
R1611 B.n205 B.n202 10.6151
R1612 B.n206 B.n205 10.6151
R1613 B.n209 B.n206 10.6151
R1614 B.n210 B.n209 10.6151
R1615 B.n213 B.n210 10.6151
R1616 B.n214 B.n213 10.6151
R1617 B.n217 B.n214 10.6151
R1618 B.n218 B.n217 10.6151
R1619 B.n221 B.n218 10.6151
R1620 B.n222 B.n221 10.6151
R1621 B.n225 B.n222 10.6151
R1622 B.n226 B.n225 10.6151
R1623 B.n229 B.n226 10.6151
R1624 B.n230 B.n229 10.6151
R1625 B.n233 B.n230 10.6151
R1626 B.n234 B.n233 10.6151
R1627 B.n237 B.n234 10.6151
R1628 B.n238 B.n237 10.6151
R1629 B.n241 B.n238 10.6151
R1630 B.n242 B.n241 10.6151
R1631 B.n245 B.n242 10.6151
R1632 B.n246 B.n245 10.6151
R1633 B.n249 B.n246 10.6151
R1634 B.n254 B.n251 10.6151
R1635 B.n255 B.n254 10.6151
R1636 B.n258 B.n255 10.6151
R1637 B.n259 B.n258 10.6151
R1638 B.n262 B.n259 10.6151
R1639 B.n263 B.n262 10.6151
R1640 B.n266 B.n263 10.6151
R1641 B.n267 B.n266 10.6151
R1642 B.n271 B.n270 10.6151
R1643 B.n274 B.n271 10.6151
R1644 B.n275 B.n274 10.6151
R1645 B.n278 B.n275 10.6151
R1646 B.n279 B.n278 10.6151
R1647 B.n282 B.n279 10.6151
R1648 B.n283 B.n282 10.6151
R1649 B.n286 B.n283 10.6151
R1650 B.n287 B.n286 10.6151
R1651 B.n290 B.n287 10.6151
R1652 B.n291 B.n290 10.6151
R1653 B.n294 B.n291 10.6151
R1654 B.n295 B.n294 10.6151
R1655 B.n298 B.n295 10.6151
R1656 B.n299 B.n298 10.6151
R1657 B.n302 B.n299 10.6151
R1658 B.n303 B.n302 10.6151
R1659 B.n306 B.n303 10.6151
R1660 B.n307 B.n306 10.6151
R1661 B.n310 B.n307 10.6151
R1662 B.n311 B.n310 10.6151
R1663 B.n314 B.n311 10.6151
R1664 B.n315 B.n314 10.6151
R1665 B.n318 B.n315 10.6151
R1666 B.n319 B.n318 10.6151
R1667 B.n322 B.n319 10.6151
R1668 B.n323 B.n322 10.6151
R1669 B.n326 B.n323 10.6151
R1670 B.n327 B.n326 10.6151
R1671 B.n330 B.n327 10.6151
R1672 B.n331 B.n330 10.6151
R1673 B.n334 B.n331 10.6151
R1674 B.n335 B.n334 10.6151
R1675 B.n338 B.n335 10.6151
R1676 B.n339 B.n338 10.6151
R1677 B.n342 B.n339 10.6151
R1678 B.n343 B.n342 10.6151
R1679 B.n346 B.n343 10.6151
R1680 B.n347 B.n346 10.6151
R1681 B.n350 B.n347 10.6151
R1682 B.n351 B.n350 10.6151
R1683 B.n354 B.n351 10.6151
R1684 B.n355 B.n354 10.6151
R1685 B.n358 B.n355 10.6151
R1686 B.n359 B.n358 10.6151
R1687 B.n362 B.n359 10.6151
R1688 B.n363 B.n362 10.6151
R1689 B.n366 B.n363 10.6151
R1690 B.n367 B.n366 10.6151
R1691 B.n370 B.n367 10.6151
R1692 B.n371 B.n370 10.6151
R1693 B.n374 B.n371 10.6151
R1694 B.n375 B.n374 10.6151
R1695 B.n378 B.n375 10.6151
R1696 B.n379 B.n378 10.6151
R1697 B.n382 B.n379 10.6151
R1698 B.n383 B.n382 10.6151
R1699 B.n386 B.n383 10.6151
R1700 B.n387 B.n386 10.6151
R1701 B.n390 B.n387 10.6151
R1702 B.n391 B.n390 10.6151
R1703 B.n903 B.n391 10.6151
R1704 B.n965 B.n0 8.11757
R1705 B.n965 B.n1 8.11757
R1706 B.n802 B.t11 8.07719
R1707 B.t9 B.n405 8.07719
R1708 B.n856 B.t7 8.07719
R1709 B.n12 B.t4 8.07719
R1710 B.n945 B.t0 8.07719
R1711 B.n920 B.t18 8.07719
R1712 B.n659 B.n513 6.5566
R1713 B.n643 B.n642 6.5566
R1714 B.n251 B.n250 6.5566
R1715 B.n267 B.n125 6.5566
R1716 B.n820 B.t3 6.28237
R1717 B.n930 B.t1 6.28237
R1718 B.n662 B.n513 4.05904
R1719 B.n642 B.n641 4.05904
R1720 B.n250 B.n249 4.05904
R1721 B.n270 B.n125 4.05904
R1722 VN.n3 VN.t2 666.87
R1723 VN.n13 VN.t4 666.87
R1724 VN.n2 VN.t3 644.831
R1725 VN.n1 VN.t9 644.831
R1726 VN.n6 VN.t6 644.831
R1727 VN.n8 VN.t1 644.831
R1728 VN.n12 VN.t7 644.831
R1729 VN.n11 VN.t0 644.831
R1730 VN.n16 VN.t5 644.831
R1731 VN.n18 VN.t8 644.831
R1732 VN.n9 VN.n8 161.3
R1733 VN.n19 VN.n18 161.3
R1734 VN.n17 VN.n10 161.3
R1735 VN.n7 VN.n0 161.3
R1736 VN.n16 VN.n15 80.6037
R1737 VN.n14 VN.n11 80.6037
R1738 VN.n6 VN.n5 80.6037
R1739 VN.n4 VN.n1 80.6037
R1740 VN VN.n19 49.0365
R1741 VN.n2 VN.n1 48.2005
R1742 VN.n6 VN.n1 48.2005
R1743 VN.n12 VN.n11 48.2005
R1744 VN.n16 VN.n11 48.2005
R1745 VN.n7 VN.n6 36.5157
R1746 VN.n17 VN.n16 36.5157
R1747 VN.n14 VN.n13 31.7379
R1748 VN.n4 VN.n3 31.7379
R1749 VN.n3 VN.n2 16.9109
R1750 VN.n13 VN.n12 16.9109
R1751 VN.n8 VN.n7 11.6853
R1752 VN.n18 VN.n17 11.6853
R1753 VN.n15 VN.n14 0.380177
R1754 VN.n5 VN.n4 0.380177
R1755 VN.n15 VN.n10 0.285035
R1756 VN.n5 VN.n0 0.285035
R1757 VN.n19 VN.n10 0.189894
R1758 VN.n9 VN.n0 0.189894
R1759 VN VN.n9 0.0516364
R1760 VDD2.n1 VDD2.t7 61.0454
R1761 VDD2.n4 VDD2.t1 60.0887
R1762 VDD2.n3 VDD2.n2 59.7219
R1763 VDD2 VDD2.n7 59.7189
R1764 VDD2.n6 VDD2.n5 59.0596
R1765 VDD2.n1 VDD2.n0 59.0596
R1766 VDD2.n4 VDD2.n3 44.8468
R1767 VDD2.n7 VDD2.t2 1.02961
R1768 VDD2.n7 VDD2.t5 1.02961
R1769 VDD2.n5 VDD2.t4 1.02961
R1770 VDD2.n5 VDD2.t9 1.02961
R1771 VDD2.n2 VDD2.t3 1.02961
R1772 VDD2.n2 VDD2.t8 1.02961
R1773 VDD2.n0 VDD2.t6 1.02961
R1774 VDD2.n0 VDD2.t0 1.02961
R1775 VDD2.n6 VDD2.n4 0.957397
R1776 VDD2 VDD2.n6 0.297914
R1777 VDD2.n3 VDD2.n1 0.184378
C0 VN VP 7.05483f
C1 VDD2 VN 11.0763f
C2 VTAIL VDD1 20.182499f
C3 VP VDD1 11.272901f
C4 VDD2 VDD1 1.02438f
C5 VN VDD1 0.149511f
C6 VTAIL VP 10.693f
C7 VDD2 VTAIL 20.2136f
C8 VDD2 VP 0.353124f
C9 VTAIL VN 10.6781f
C10 VDD2 B 6.360659f
C11 VDD1 B 6.287717f
C12 VTAIL B 9.23552f
C13 VN B 10.637541f
C14 VP B 8.37477f
C15 VDD2.t7 B 4.26451f
C16 VDD2.t6 B 0.365017f
C17 VDD2.t0 B 0.365017f
C18 VDD2.n0 B 3.33131f
C19 VDD2.n1 B 0.643228f
C20 VDD2.t3 B 0.365017f
C21 VDD2.t8 B 0.365017f
C22 VDD2.n2 B 3.33506f
C23 VDD2.n3 B 2.30551f
C24 VDD2.t1 B 4.25895f
C25 VDD2.n4 B 2.86696f
C26 VDD2.t4 B 0.365017f
C27 VDD2.t9 B 0.365017f
C28 VDD2.n5 B 3.3313f
C29 VDD2.n6 B 0.300015f
C30 VDD2.t2 B 0.365017f
C31 VDD2.t5 B 0.365017f
C32 VDD2.n7 B 3.33502f
C33 VN.n0 B 0.054275f
C34 VN.t9 B 1.72933f
C35 VN.n1 B 0.656549f
C36 VN.t2 B 1.75073f
C37 VN.t3 B 1.72933f
C38 VN.n2 B 0.655777f
C39 VN.n3 B 0.630078f
C40 VN.n4 B 0.247138f
C41 VN.n5 B 0.067749f
C42 VN.t6 B 1.72933f
C43 VN.n6 B 0.654543f
C44 VN.n7 B 0.00923f
C45 VN.t1 B 1.72933f
C46 VN.n8 B 0.64105f
C47 VN.n9 B 0.031521f
C48 VN.n10 B 0.054275f
C49 VN.t0 B 1.72933f
C50 VN.n11 B 0.656549f
C51 VN.t5 B 1.72933f
C52 VN.t4 B 1.75073f
C53 VN.t7 B 1.72933f
C54 VN.n12 B 0.655777f
C55 VN.n13 B 0.630078f
C56 VN.n14 B 0.247138f
C57 VN.n15 B 0.067749f
C58 VN.n16 B 0.654543f
C59 VN.n17 B 0.00923f
C60 VN.t8 B 1.72933f
C61 VN.n18 B 0.64105f
C62 VN.n19 B 2.14839f
C63 VDD1.t9 B 4.27963f
C64 VDD1.t5 B 0.366312f
C65 VDD1.t3 B 0.366312f
C66 VDD1.n0 B 3.34312f
C67 VDD1.n1 B 0.651288f
C68 VDD1.t8 B 4.27963f
C69 VDD1.t2 B 0.366312f
C70 VDD1.t4 B 0.366312f
C71 VDD1.n2 B 3.34312f
C72 VDD1.n3 B 0.645509f
C73 VDD1.t1 B 0.366312f
C74 VDD1.t6 B 0.366312f
C75 VDD1.n4 B 3.34689f
C76 VDD1.n5 B 2.39155f
C77 VDD1.t0 B 0.366312f
C78 VDD1.t7 B 0.366312f
C79 VDD1.n6 B 3.34311f
C80 VDD1.n7 B 2.87137f
C81 VTAIL.t4 B 0.374713f
C82 VTAIL.t8 B 0.374713f
C83 VTAIL.n0 B 3.33964f
C84 VTAIL.n1 B 0.391948f
C85 VTAIL.t10 B 4.26705f
C86 VTAIL.n2 B 0.500853f
C87 VTAIL.t12 B 0.374713f
C88 VTAIL.t17 B 0.374713f
C89 VTAIL.n3 B 3.33964f
C90 VTAIL.n4 B 0.407009f
C91 VTAIL.t15 B 0.374713f
C92 VTAIL.t14 B 0.374713f
C93 VTAIL.n5 B 3.33964f
C94 VTAIL.n6 B 2.13495f
C95 VTAIL.t3 B 0.374713f
C96 VTAIL.t5 B 0.374713f
C97 VTAIL.n7 B 3.33963f
C98 VTAIL.n8 B 2.13496f
C99 VTAIL.t19 B 0.374713f
C100 VTAIL.t2 B 0.374713f
C101 VTAIL.n9 B 3.33963f
C102 VTAIL.n10 B 0.407016f
C103 VTAIL.t7 B 4.26706f
C104 VTAIL.n11 B 0.500848f
C105 VTAIL.t9 B 0.374713f
C106 VTAIL.t16 B 0.374713f
C107 VTAIL.n12 B 3.33963f
C108 VTAIL.n13 B 0.406332f
C109 VTAIL.t11 B 0.374713f
C110 VTAIL.t13 B 0.374713f
C111 VTAIL.n14 B 3.33963f
C112 VTAIL.n15 B 0.407016f
C113 VTAIL.t18 B 4.26705f
C114 VTAIL.n16 B 2.15349f
C115 VTAIL.t1 B 4.26705f
C116 VTAIL.n17 B 2.15349f
C117 VTAIL.t0 B 0.374713f
C118 VTAIL.t6 B 0.374713f
C119 VTAIL.n18 B 3.33964f
C120 VTAIL.n19 B 0.345395f
C121 VP.n0 B 0.054759f
C122 VP.t5 B 1.74475f
C123 VP.n1 B 0.662403f
C124 VP.n2 B 0.054759f
C125 VP.n3 B 0.054759f
C126 VP.t2 B 1.74475f
C127 VP.t9 B 1.74475f
C128 VP.n4 B 0.068353f
C129 VP.t6 B 1.74475f
C130 VP.n5 B 0.249341f
C131 VP.t4 B 1.74475f
C132 VP.t0 B 1.76634f
C133 VP.n6 B 0.635696f
C134 VP.n7 B 0.661624f
C135 VP.n8 B 0.662403f
C136 VP.n9 B 0.660379f
C137 VP.n10 B 0.009312f
C138 VP.n11 B 0.646765f
C139 VP.n12 B 2.14083f
C140 VP.n13 B 2.17123f
C141 VP.t1 B 1.74475f
C142 VP.n14 B 0.646765f
C143 VP.n15 B 0.009312f
C144 VP.t7 B 1.74475f
C145 VP.n16 B 0.660379f
C146 VP.n17 B 0.068353f
C147 VP.n18 B 0.082075f
C148 VP.n19 B 0.068353f
C149 VP.t8 B 1.74475f
C150 VP.n20 B 0.660379f
C151 VP.n21 B 0.009312f
C152 VP.t3 B 1.74475f
C153 VP.n22 B 0.646765f
C154 VP.n23 B 0.031802f
.ends

