* NGSPICE file created from diff_pair_sample_1661.ext - technology: sky130A

.subckt diff_pair_sample_1661 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X1 VTAIL.t18 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X2 VDD1.t9 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.22
X3 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.22
X4 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.22
X5 VDD1.t8 VP.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.22
X6 VTAIL.t2 VP.t2 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X7 VDD1.t6 VP.t3 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.22
X8 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.22
X9 VDD1.t5 VP.t4 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X10 VDD2.t3 VN.t2 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X11 VTAIL.t16 VN.t3 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X12 VDD2.t7 VN.t4 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.22
X13 VDD2.t8 VN.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X14 VDD1.t4 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.22
X15 VTAIL.t5 VP.t6 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X16 VTAIL.t7 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X17 VDD2.t0 VN.t6 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.22
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.22
X19 VDD2.t1 VN.t7 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.22
X20 VDD2.t4 VN.t8 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.22
X21 VTAIL.t0 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X22 VTAIL.t10 VN.t9 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
X23 VDD1.t0 VP.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.22
R0 VN.n8 VN.t7 1863
R1 VN.n2 VN.t8 1863
R2 VN.n18 VN.t4 1863
R3 VN.n12 VN.t6 1863
R4 VN.n7 VN.t1 1811.88
R5 VN.n5 VN.t2 1811.88
R6 VN.n1 VN.t3 1811.88
R7 VN.n17 VN.t9 1811.88
R8 VN.n15 VN.t5 1811.88
R9 VN.n11 VN.t0 1811.88
R10 VN.n13 VN.n12 161.489
R11 VN.n3 VN.n2 161.489
R12 VN.n9 VN.n8 161.3
R13 VN.n19 VN.n18 161.3
R14 VN.n16 VN.n10 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n6 VN.n0 161.3
R17 VN.n4 VN.n3 161.3
R18 VN.n4 VN.n1 43.8187
R19 VN.n7 VN.n6 43.8187
R20 VN.n17 VN.n16 43.8187
R21 VN.n14 VN.n11 43.8187
R22 VN VN.n19 43.1122
R23 VN.n5 VN.n4 36.5157
R24 VN.n6 VN.n5 36.5157
R25 VN.n16 VN.n15 36.5157
R26 VN.n15 VN.n14 36.5157
R27 VN.n2 VN.n1 29.2126
R28 VN.n8 VN.n7 29.2126
R29 VN.n18 VN.n17 29.2126
R30 VN.n12 VN.n11 29.2126
R31 VN.n19 VN.n10 0.189894
R32 VN.n13 VN.n10 0.189894
R33 VN.n3 VN.n0 0.189894
R34 VN.n9 VN.n0 0.189894
R35 VN VN.n9 0.0516364
R36 VDD2.n1 VDD2.t4 60.7204
R37 VDD2.n4 VDD2.t7 60.2464
R38 VDD2.n3 VDD2.n2 59.2473
R39 VDD2 VDD2.n7 59.2447
R40 VDD2.n6 VDD2.n5 58.9473
R41 VDD2.n1 VDD2.n0 58.9471
R42 VDD2.n4 VDD2.n3 39.1054
R43 VDD2.n7 VDD2.t9 1.29971
R44 VDD2.n7 VDD2.t0 1.29971
R45 VDD2.n5 VDD2.t6 1.29971
R46 VDD2.n5 VDD2.t8 1.29971
R47 VDD2.n2 VDD2.t2 1.29971
R48 VDD2.n2 VDD2.t1 1.29971
R49 VDD2.n0 VDD2.t5 1.29971
R50 VDD2.n0 VDD2.t3 1.29971
R51 VDD2.n6 VDD2.n4 0.474638
R52 VDD2 VDD2.n6 0.177224
R53 VDD2.n3 VDD2.n1 0.0636885
R54 VTAIL.n16 VTAIL.t6 43.5677
R55 VTAIL.n11 VTAIL.t13 43.5677
R56 VTAIL.n17 VTAIL.t12 43.5675
R57 VTAIL.n2 VTAIL.t3 43.5675
R58 VTAIL.n15 VTAIL.n14 42.2685
R59 VTAIL.n13 VTAIL.n12 42.2685
R60 VTAIL.n10 VTAIL.n9 42.2685
R61 VTAIL.n8 VTAIL.n7 42.2685
R62 VTAIL.n19 VTAIL.n18 42.2683
R63 VTAIL.n1 VTAIL.n0 42.2683
R64 VTAIL.n4 VTAIL.n3 42.2683
R65 VTAIL.n6 VTAIL.n5 42.2683
R66 VTAIL.n8 VTAIL.n6 26.4531
R67 VTAIL.n17 VTAIL.n16 25.9789
R68 VTAIL.n18 VTAIL.t17 1.29971
R69 VTAIL.n18 VTAIL.t18 1.29971
R70 VTAIL.n0 VTAIL.t11 1.29971
R71 VTAIL.n0 VTAIL.t16 1.29971
R72 VTAIL.n3 VTAIL.t1 1.29971
R73 VTAIL.n3 VTAIL.t2 1.29971
R74 VTAIL.n5 VTAIL.t9 1.29971
R75 VTAIL.n5 VTAIL.t5 1.29971
R76 VTAIL.n14 VTAIL.t8 1.29971
R77 VTAIL.n14 VTAIL.t0 1.29971
R78 VTAIL.n12 VTAIL.t4 1.29971
R79 VTAIL.n12 VTAIL.t7 1.29971
R80 VTAIL.n9 VTAIL.t14 1.29971
R81 VTAIL.n9 VTAIL.t19 1.29971
R82 VTAIL.n7 VTAIL.t15 1.29971
R83 VTAIL.n7 VTAIL.t10 1.29971
R84 VTAIL.n13 VTAIL.n11 0.707397
R85 VTAIL.n2 VTAIL.n1 0.707397
R86 VTAIL.n10 VTAIL.n8 0.474638
R87 VTAIL.n11 VTAIL.n10 0.474638
R88 VTAIL.n15 VTAIL.n13 0.474638
R89 VTAIL.n16 VTAIL.n15 0.474638
R90 VTAIL.n6 VTAIL.n4 0.474638
R91 VTAIL.n4 VTAIL.n2 0.474638
R92 VTAIL.n19 VTAIL.n17 0.474638
R93 VTAIL VTAIL.n1 0.414293
R94 VTAIL VTAIL.n19 0.0608448
R95 B.n165 B.t21 1900.35
R96 B.n159 B.t10 1900.35
R97 B.n64 B.t18 1900.35
R98 B.n71 B.t14 1900.35
R99 B.n495 B.n494 585
R100 B.n497 B.n97 585
R101 B.n500 B.n499 585
R102 B.n501 B.n96 585
R103 B.n503 B.n502 585
R104 B.n505 B.n95 585
R105 B.n508 B.n507 585
R106 B.n509 B.n94 585
R107 B.n511 B.n510 585
R108 B.n513 B.n93 585
R109 B.n516 B.n515 585
R110 B.n517 B.n92 585
R111 B.n519 B.n518 585
R112 B.n521 B.n91 585
R113 B.n524 B.n523 585
R114 B.n525 B.n90 585
R115 B.n527 B.n526 585
R116 B.n529 B.n89 585
R117 B.n532 B.n531 585
R118 B.n533 B.n88 585
R119 B.n535 B.n534 585
R120 B.n537 B.n87 585
R121 B.n540 B.n539 585
R122 B.n541 B.n86 585
R123 B.n543 B.n542 585
R124 B.n545 B.n85 585
R125 B.n548 B.n547 585
R126 B.n549 B.n84 585
R127 B.n551 B.n550 585
R128 B.n553 B.n83 585
R129 B.n556 B.n555 585
R130 B.n557 B.n82 585
R131 B.n559 B.n558 585
R132 B.n561 B.n81 585
R133 B.n564 B.n563 585
R134 B.n565 B.n80 585
R135 B.n567 B.n566 585
R136 B.n569 B.n79 585
R137 B.n572 B.n571 585
R138 B.n573 B.n78 585
R139 B.n575 B.n574 585
R140 B.n577 B.n77 585
R141 B.n580 B.n579 585
R142 B.n581 B.n76 585
R143 B.n583 B.n582 585
R144 B.n585 B.n75 585
R145 B.n588 B.n587 585
R146 B.n589 B.n74 585
R147 B.n591 B.n590 585
R148 B.n593 B.n73 585
R149 B.n596 B.n595 585
R150 B.n598 B.n70 585
R151 B.n600 B.n599 585
R152 B.n602 B.n69 585
R153 B.n605 B.n604 585
R154 B.n606 B.n68 585
R155 B.n608 B.n607 585
R156 B.n610 B.n67 585
R157 B.n613 B.n612 585
R158 B.n614 B.n63 585
R159 B.n616 B.n615 585
R160 B.n618 B.n62 585
R161 B.n621 B.n620 585
R162 B.n622 B.n61 585
R163 B.n624 B.n623 585
R164 B.n626 B.n60 585
R165 B.n629 B.n628 585
R166 B.n630 B.n59 585
R167 B.n632 B.n631 585
R168 B.n634 B.n58 585
R169 B.n637 B.n636 585
R170 B.n638 B.n57 585
R171 B.n640 B.n639 585
R172 B.n642 B.n56 585
R173 B.n645 B.n644 585
R174 B.n646 B.n55 585
R175 B.n648 B.n647 585
R176 B.n650 B.n54 585
R177 B.n653 B.n652 585
R178 B.n654 B.n53 585
R179 B.n656 B.n655 585
R180 B.n658 B.n52 585
R181 B.n661 B.n660 585
R182 B.n662 B.n51 585
R183 B.n664 B.n663 585
R184 B.n666 B.n50 585
R185 B.n669 B.n668 585
R186 B.n670 B.n49 585
R187 B.n672 B.n671 585
R188 B.n674 B.n48 585
R189 B.n677 B.n676 585
R190 B.n678 B.n47 585
R191 B.n680 B.n679 585
R192 B.n682 B.n46 585
R193 B.n685 B.n684 585
R194 B.n686 B.n45 585
R195 B.n688 B.n687 585
R196 B.n690 B.n44 585
R197 B.n693 B.n692 585
R198 B.n694 B.n43 585
R199 B.n696 B.n695 585
R200 B.n698 B.n42 585
R201 B.n701 B.n700 585
R202 B.n702 B.n41 585
R203 B.n704 B.n703 585
R204 B.n706 B.n40 585
R205 B.n709 B.n708 585
R206 B.n710 B.n39 585
R207 B.n712 B.n711 585
R208 B.n714 B.n38 585
R209 B.n717 B.n716 585
R210 B.n718 B.n37 585
R211 B.n493 B.n35 585
R212 B.n721 B.n35 585
R213 B.n492 B.n34 585
R214 B.n722 B.n34 585
R215 B.n491 B.n33 585
R216 B.n723 B.n33 585
R217 B.n490 B.n489 585
R218 B.n489 B.n29 585
R219 B.n488 B.n28 585
R220 B.n729 B.n28 585
R221 B.n487 B.n27 585
R222 B.n730 B.n27 585
R223 B.n486 B.n26 585
R224 B.n731 B.n26 585
R225 B.n485 B.n484 585
R226 B.n484 B.n22 585
R227 B.n483 B.n21 585
R228 B.n737 B.n21 585
R229 B.n482 B.n20 585
R230 B.n738 B.n20 585
R231 B.n481 B.n19 585
R232 B.n739 B.n19 585
R233 B.n480 B.n479 585
R234 B.n479 B.n15 585
R235 B.n478 B.n14 585
R236 B.n745 B.n14 585
R237 B.n477 B.n13 585
R238 B.n746 B.n13 585
R239 B.n476 B.n12 585
R240 B.n747 B.n12 585
R241 B.n475 B.n474 585
R242 B.n474 B.n11 585
R243 B.n473 B.n7 585
R244 B.n753 B.n7 585
R245 B.n472 B.n6 585
R246 B.n754 B.n6 585
R247 B.n471 B.n5 585
R248 B.n755 B.n5 585
R249 B.n470 B.n469 585
R250 B.n469 B.n4 585
R251 B.n468 B.n98 585
R252 B.n468 B.n467 585
R253 B.n457 B.n99 585
R254 B.n460 B.n99 585
R255 B.n459 B.n458 585
R256 B.n461 B.n459 585
R257 B.n456 B.n103 585
R258 B.n107 B.n103 585
R259 B.n455 B.n454 585
R260 B.n454 B.n453 585
R261 B.n105 B.n104 585
R262 B.n106 B.n105 585
R263 B.n446 B.n445 585
R264 B.n447 B.n446 585
R265 B.n444 B.n111 585
R266 B.n115 B.n111 585
R267 B.n443 B.n442 585
R268 B.n442 B.n441 585
R269 B.n113 B.n112 585
R270 B.n114 B.n113 585
R271 B.n434 B.n433 585
R272 B.n435 B.n434 585
R273 B.n432 B.n120 585
R274 B.n120 B.n119 585
R275 B.n431 B.n430 585
R276 B.n430 B.n429 585
R277 B.n122 B.n121 585
R278 B.n123 B.n122 585
R279 B.n422 B.n421 585
R280 B.n423 B.n422 585
R281 B.n420 B.n128 585
R282 B.n128 B.n127 585
R283 B.n419 B.n418 585
R284 B.n418 B.n417 585
R285 B.n414 B.n132 585
R286 B.n413 B.n412 585
R287 B.n410 B.n133 585
R288 B.n410 B.n131 585
R289 B.n409 B.n408 585
R290 B.n407 B.n406 585
R291 B.n405 B.n135 585
R292 B.n403 B.n402 585
R293 B.n401 B.n136 585
R294 B.n400 B.n399 585
R295 B.n397 B.n137 585
R296 B.n395 B.n394 585
R297 B.n393 B.n138 585
R298 B.n392 B.n391 585
R299 B.n389 B.n139 585
R300 B.n387 B.n386 585
R301 B.n385 B.n140 585
R302 B.n384 B.n383 585
R303 B.n381 B.n141 585
R304 B.n379 B.n378 585
R305 B.n377 B.n142 585
R306 B.n376 B.n375 585
R307 B.n373 B.n143 585
R308 B.n371 B.n370 585
R309 B.n369 B.n144 585
R310 B.n368 B.n367 585
R311 B.n365 B.n145 585
R312 B.n363 B.n362 585
R313 B.n361 B.n146 585
R314 B.n360 B.n359 585
R315 B.n357 B.n147 585
R316 B.n355 B.n354 585
R317 B.n353 B.n148 585
R318 B.n352 B.n351 585
R319 B.n349 B.n149 585
R320 B.n347 B.n346 585
R321 B.n345 B.n150 585
R322 B.n344 B.n343 585
R323 B.n341 B.n151 585
R324 B.n339 B.n338 585
R325 B.n337 B.n152 585
R326 B.n336 B.n335 585
R327 B.n333 B.n153 585
R328 B.n331 B.n330 585
R329 B.n329 B.n154 585
R330 B.n328 B.n327 585
R331 B.n325 B.n155 585
R332 B.n323 B.n322 585
R333 B.n321 B.n156 585
R334 B.n320 B.n319 585
R335 B.n317 B.n157 585
R336 B.n315 B.n314 585
R337 B.n312 B.n158 585
R338 B.n311 B.n310 585
R339 B.n308 B.n161 585
R340 B.n306 B.n305 585
R341 B.n304 B.n162 585
R342 B.n303 B.n302 585
R343 B.n300 B.n163 585
R344 B.n298 B.n297 585
R345 B.n296 B.n164 585
R346 B.n295 B.n294 585
R347 B.n292 B.n291 585
R348 B.n290 B.n289 585
R349 B.n288 B.n169 585
R350 B.n286 B.n285 585
R351 B.n284 B.n170 585
R352 B.n283 B.n282 585
R353 B.n280 B.n171 585
R354 B.n278 B.n277 585
R355 B.n276 B.n172 585
R356 B.n275 B.n274 585
R357 B.n272 B.n173 585
R358 B.n270 B.n269 585
R359 B.n268 B.n174 585
R360 B.n267 B.n266 585
R361 B.n264 B.n175 585
R362 B.n262 B.n261 585
R363 B.n260 B.n176 585
R364 B.n259 B.n258 585
R365 B.n256 B.n177 585
R366 B.n254 B.n253 585
R367 B.n252 B.n178 585
R368 B.n251 B.n250 585
R369 B.n248 B.n179 585
R370 B.n246 B.n245 585
R371 B.n244 B.n180 585
R372 B.n243 B.n242 585
R373 B.n240 B.n181 585
R374 B.n238 B.n237 585
R375 B.n236 B.n182 585
R376 B.n235 B.n234 585
R377 B.n232 B.n183 585
R378 B.n230 B.n229 585
R379 B.n228 B.n184 585
R380 B.n227 B.n226 585
R381 B.n224 B.n185 585
R382 B.n222 B.n221 585
R383 B.n220 B.n186 585
R384 B.n219 B.n218 585
R385 B.n216 B.n187 585
R386 B.n214 B.n213 585
R387 B.n212 B.n188 585
R388 B.n211 B.n210 585
R389 B.n208 B.n189 585
R390 B.n206 B.n205 585
R391 B.n204 B.n190 585
R392 B.n203 B.n202 585
R393 B.n200 B.n191 585
R394 B.n198 B.n197 585
R395 B.n196 B.n192 585
R396 B.n195 B.n194 585
R397 B.n130 B.n129 585
R398 B.n131 B.n130 585
R399 B.n416 B.n415 585
R400 B.n417 B.n416 585
R401 B.n126 B.n125 585
R402 B.n127 B.n126 585
R403 B.n425 B.n424 585
R404 B.n424 B.n423 585
R405 B.n426 B.n124 585
R406 B.n124 B.n123 585
R407 B.n428 B.n427 585
R408 B.n429 B.n428 585
R409 B.n118 B.n117 585
R410 B.n119 B.n118 585
R411 B.n437 B.n436 585
R412 B.n436 B.n435 585
R413 B.n438 B.n116 585
R414 B.n116 B.n114 585
R415 B.n440 B.n439 585
R416 B.n441 B.n440 585
R417 B.n110 B.n109 585
R418 B.n115 B.n110 585
R419 B.n449 B.n448 585
R420 B.n448 B.n447 585
R421 B.n450 B.n108 585
R422 B.n108 B.n106 585
R423 B.n452 B.n451 585
R424 B.n453 B.n452 585
R425 B.n102 B.n101 585
R426 B.n107 B.n102 585
R427 B.n463 B.n462 585
R428 B.n462 B.n461 585
R429 B.n464 B.n100 585
R430 B.n460 B.n100 585
R431 B.n466 B.n465 585
R432 B.n467 B.n466 585
R433 B.n2 B.n0 585
R434 B.n4 B.n2 585
R435 B.n3 B.n1 585
R436 B.n754 B.n3 585
R437 B.n752 B.n751 585
R438 B.n753 B.n752 585
R439 B.n750 B.n8 585
R440 B.n11 B.n8 585
R441 B.n749 B.n748 585
R442 B.n748 B.n747 585
R443 B.n10 B.n9 585
R444 B.n746 B.n10 585
R445 B.n744 B.n743 585
R446 B.n745 B.n744 585
R447 B.n742 B.n16 585
R448 B.n16 B.n15 585
R449 B.n741 B.n740 585
R450 B.n740 B.n739 585
R451 B.n18 B.n17 585
R452 B.n738 B.n18 585
R453 B.n736 B.n735 585
R454 B.n737 B.n736 585
R455 B.n734 B.n23 585
R456 B.n23 B.n22 585
R457 B.n733 B.n732 585
R458 B.n732 B.n731 585
R459 B.n25 B.n24 585
R460 B.n730 B.n25 585
R461 B.n728 B.n727 585
R462 B.n729 B.n728 585
R463 B.n726 B.n30 585
R464 B.n30 B.n29 585
R465 B.n725 B.n724 585
R466 B.n724 B.n723 585
R467 B.n32 B.n31 585
R468 B.n722 B.n32 585
R469 B.n720 B.n719 585
R470 B.n721 B.n720 585
R471 B.n757 B.n756 585
R472 B.n756 B.n755 585
R473 B.n416 B.n132 458.866
R474 B.n720 B.n37 458.866
R475 B.n418 B.n130 458.866
R476 B.n495 B.n35 458.866
R477 B.n496 B.n36 256.663
R478 B.n498 B.n36 256.663
R479 B.n504 B.n36 256.663
R480 B.n506 B.n36 256.663
R481 B.n512 B.n36 256.663
R482 B.n514 B.n36 256.663
R483 B.n520 B.n36 256.663
R484 B.n522 B.n36 256.663
R485 B.n528 B.n36 256.663
R486 B.n530 B.n36 256.663
R487 B.n536 B.n36 256.663
R488 B.n538 B.n36 256.663
R489 B.n544 B.n36 256.663
R490 B.n546 B.n36 256.663
R491 B.n552 B.n36 256.663
R492 B.n554 B.n36 256.663
R493 B.n560 B.n36 256.663
R494 B.n562 B.n36 256.663
R495 B.n568 B.n36 256.663
R496 B.n570 B.n36 256.663
R497 B.n576 B.n36 256.663
R498 B.n578 B.n36 256.663
R499 B.n584 B.n36 256.663
R500 B.n586 B.n36 256.663
R501 B.n592 B.n36 256.663
R502 B.n594 B.n36 256.663
R503 B.n601 B.n36 256.663
R504 B.n603 B.n36 256.663
R505 B.n609 B.n36 256.663
R506 B.n611 B.n36 256.663
R507 B.n617 B.n36 256.663
R508 B.n619 B.n36 256.663
R509 B.n625 B.n36 256.663
R510 B.n627 B.n36 256.663
R511 B.n633 B.n36 256.663
R512 B.n635 B.n36 256.663
R513 B.n641 B.n36 256.663
R514 B.n643 B.n36 256.663
R515 B.n649 B.n36 256.663
R516 B.n651 B.n36 256.663
R517 B.n657 B.n36 256.663
R518 B.n659 B.n36 256.663
R519 B.n665 B.n36 256.663
R520 B.n667 B.n36 256.663
R521 B.n673 B.n36 256.663
R522 B.n675 B.n36 256.663
R523 B.n681 B.n36 256.663
R524 B.n683 B.n36 256.663
R525 B.n689 B.n36 256.663
R526 B.n691 B.n36 256.663
R527 B.n697 B.n36 256.663
R528 B.n699 B.n36 256.663
R529 B.n705 B.n36 256.663
R530 B.n707 B.n36 256.663
R531 B.n713 B.n36 256.663
R532 B.n715 B.n36 256.663
R533 B.n411 B.n131 256.663
R534 B.n134 B.n131 256.663
R535 B.n404 B.n131 256.663
R536 B.n398 B.n131 256.663
R537 B.n396 B.n131 256.663
R538 B.n390 B.n131 256.663
R539 B.n388 B.n131 256.663
R540 B.n382 B.n131 256.663
R541 B.n380 B.n131 256.663
R542 B.n374 B.n131 256.663
R543 B.n372 B.n131 256.663
R544 B.n366 B.n131 256.663
R545 B.n364 B.n131 256.663
R546 B.n358 B.n131 256.663
R547 B.n356 B.n131 256.663
R548 B.n350 B.n131 256.663
R549 B.n348 B.n131 256.663
R550 B.n342 B.n131 256.663
R551 B.n340 B.n131 256.663
R552 B.n334 B.n131 256.663
R553 B.n332 B.n131 256.663
R554 B.n326 B.n131 256.663
R555 B.n324 B.n131 256.663
R556 B.n318 B.n131 256.663
R557 B.n316 B.n131 256.663
R558 B.n309 B.n131 256.663
R559 B.n307 B.n131 256.663
R560 B.n301 B.n131 256.663
R561 B.n299 B.n131 256.663
R562 B.n293 B.n131 256.663
R563 B.n168 B.n131 256.663
R564 B.n287 B.n131 256.663
R565 B.n281 B.n131 256.663
R566 B.n279 B.n131 256.663
R567 B.n273 B.n131 256.663
R568 B.n271 B.n131 256.663
R569 B.n265 B.n131 256.663
R570 B.n263 B.n131 256.663
R571 B.n257 B.n131 256.663
R572 B.n255 B.n131 256.663
R573 B.n249 B.n131 256.663
R574 B.n247 B.n131 256.663
R575 B.n241 B.n131 256.663
R576 B.n239 B.n131 256.663
R577 B.n233 B.n131 256.663
R578 B.n231 B.n131 256.663
R579 B.n225 B.n131 256.663
R580 B.n223 B.n131 256.663
R581 B.n217 B.n131 256.663
R582 B.n215 B.n131 256.663
R583 B.n209 B.n131 256.663
R584 B.n207 B.n131 256.663
R585 B.n201 B.n131 256.663
R586 B.n199 B.n131 256.663
R587 B.n193 B.n131 256.663
R588 B.n416 B.n126 163.367
R589 B.n424 B.n126 163.367
R590 B.n424 B.n124 163.367
R591 B.n428 B.n124 163.367
R592 B.n428 B.n118 163.367
R593 B.n436 B.n118 163.367
R594 B.n436 B.n116 163.367
R595 B.n440 B.n116 163.367
R596 B.n440 B.n110 163.367
R597 B.n448 B.n110 163.367
R598 B.n448 B.n108 163.367
R599 B.n452 B.n108 163.367
R600 B.n452 B.n102 163.367
R601 B.n462 B.n102 163.367
R602 B.n462 B.n100 163.367
R603 B.n466 B.n100 163.367
R604 B.n466 B.n2 163.367
R605 B.n756 B.n2 163.367
R606 B.n756 B.n3 163.367
R607 B.n752 B.n3 163.367
R608 B.n752 B.n8 163.367
R609 B.n748 B.n8 163.367
R610 B.n748 B.n10 163.367
R611 B.n744 B.n10 163.367
R612 B.n744 B.n16 163.367
R613 B.n740 B.n16 163.367
R614 B.n740 B.n18 163.367
R615 B.n736 B.n18 163.367
R616 B.n736 B.n23 163.367
R617 B.n732 B.n23 163.367
R618 B.n732 B.n25 163.367
R619 B.n728 B.n25 163.367
R620 B.n728 B.n30 163.367
R621 B.n724 B.n30 163.367
R622 B.n724 B.n32 163.367
R623 B.n720 B.n32 163.367
R624 B.n412 B.n410 163.367
R625 B.n410 B.n409 163.367
R626 B.n406 B.n405 163.367
R627 B.n403 B.n136 163.367
R628 B.n399 B.n397 163.367
R629 B.n395 B.n138 163.367
R630 B.n391 B.n389 163.367
R631 B.n387 B.n140 163.367
R632 B.n383 B.n381 163.367
R633 B.n379 B.n142 163.367
R634 B.n375 B.n373 163.367
R635 B.n371 B.n144 163.367
R636 B.n367 B.n365 163.367
R637 B.n363 B.n146 163.367
R638 B.n359 B.n357 163.367
R639 B.n355 B.n148 163.367
R640 B.n351 B.n349 163.367
R641 B.n347 B.n150 163.367
R642 B.n343 B.n341 163.367
R643 B.n339 B.n152 163.367
R644 B.n335 B.n333 163.367
R645 B.n331 B.n154 163.367
R646 B.n327 B.n325 163.367
R647 B.n323 B.n156 163.367
R648 B.n319 B.n317 163.367
R649 B.n315 B.n158 163.367
R650 B.n310 B.n308 163.367
R651 B.n306 B.n162 163.367
R652 B.n302 B.n300 163.367
R653 B.n298 B.n164 163.367
R654 B.n294 B.n292 163.367
R655 B.n289 B.n288 163.367
R656 B.n286 B.n170 163.367
R657 B.n282 B.n280 163.367
R658 B.n278 B.n172 163.367
R659 B.n274 B.n272 163.367
R660 B.n270 B.n174 163.367
R661 B.n266 B.n264 163.367
R662 B.n262 B.n176 163.367
R663 B.n258 B.n256 163.367
R664 B.n254 B.n178 163.367
R665 B.n250 B.n248 163.367
R666 B.n246 B.n180 163.367
R667 B.n242 B.n240 163.367
R668 B.n238 B.n182 163.367
R669 B.n234 B.n232 163.367
R670 B.n230 B.n184 163.367
R671 B.n226 B.n224 163.367
R672 B.n222 B.n186 163.367
R673 B.n218 B.n216 163.367
R674 B.n214 B.n188 163.367
R675 B.n210 B.n208 163.367
R676 B.n206 B.n190 163.367
R677 B.n202 B.n200 163.367
R678 B.n198 B.n192 163.367
R679 B.n194 B.n130 163.367
R680 B.n418 B.n128 163.367
R681 B.n422 B.n128 163.367
R682 B.n422 B.n122 163.367
R683 B.n430 B.n122 163.367
R684 B.n430 B.n120 163.367
R685 B.n434 B.n120 163.367
R686 B.n434 B.n113 163.367
R687 B.n442 B.n113 163.367
R688 B.n442 B.n111 163.367
R689 B.n446 B.n111 163.367
R690 B.n446 B.n105 163.367
R691 B.n454 B.n105 163.367
R692 B.n454 B.n103 163.367
R693 B.n459 B.n103 163.367
R694 B.n459 B.n99 163.367
R695 B.n468 B.n99 163.367
R696 B.n469 B.n468 163.367
R697 B.n469 B.n5 163.367
R698 B.n6 B.n5 163.367
R699 B.n7 B.n6 163.367
R700 B.n474 B.n7 163.367
R701 B.n474 B.n12 163.367
R702 B.n13 B.n12 163.367
R703 B.n14 B.n13 163.367
R704 B.n479 B.n14 163.367
R705 B.n479 B.n19 163.367
R706 B.n20 B.n19 163.367
R707 B.n21 B.n20 163.367
R708 B.n484 B.n21 163.367
R709 B.n484 B.n26 163.367
R710 B.n27 B.n26 163.367
R711 B.n28 B.n27 163.367
R712 B.n489 B.n28 163.367
R713 B.n489 B.n33 163.367
R714 B.n34 B.n33 163.367
R715 B.n35 B.n34 163.367
R716 B.n716 B.n714 163.367
R717 B.n712 B.n39 163.367
R718 B.n708 B.n706 163.367
R719 B.n704 B.n41 163.367
R720 B.n700 B.n698 163.367
R721 B.n696 B.n43 163.367
R722 B.n692 B.n690 163.367
R723 B.n688 B.n45 163.367
R724 B.n684 B.n682 163.367
R725 B.n680 B.n47 163.367
R726 B.n676 B.n674 163.367
R727 B.n672 B.n49 163.367
R728 B.n668 B.n666 163.367
R729 B.n664 B.n51 163.367
R730 B.n660 B.n658 163.367
R731 B.n656 B.n53 163.367
R732 B.n652 B.n650 163.367
R733 B.n648 B.n55 163.367
R734 B.n644 B.n642 163.367
R735 B.n640 B.n57 163.367
R736 B.n636 B.n634 163.367
R737 B.n632 B.n59 163.367
R738 B.n628 B.n626 163.367
R739 B.n624 B.n61 163.367
R740 B.n620 B.n618 163.367
R741 B.n616 B.n63 163.367
R742 B.n612 B.n610 163.367
R743 B.n608 B.n68 163.367
R744 B.n604 B.n602 163.367
R745 B.n600 B.n70 163.367
R746 B.n595 B.n593 163.367
R747 B.n591 B.n74 163.367
R748 B.n587 B.n585 163.367
R749 B.n583 B.n76 163.367
R750 B.n579 B.n577 163.367
R751 B.n575 B.n78 163.367
R752 B.n571 B.n569 163.367
R753 B.n567 B.n80 163.367
R754 B.n563 B.n561 163.367
R755 B.n559 B.n82 163.367
R756 B.n555 B.n553 163.367
R757 B.n551 B.n84 163.367
R758 B.n547 B.n545 163.367
R759 B.n543 B.n86 163.367
R760 B.n539 B.n537 163.367
R761 B.n535 B.n88 163.367
R762 B.n531 B.n529 163.367
R763 B.n527 B.n90 163.367
R764 B.n523 B.n521 163.367
R765 B.n519 B.n92 163.367
R766 B.n515 B.n513 163.367
R767 B.n511 B.n94 163.367
R768 B.n507 B.n505 163.367
R769 B.n503 B.n96 163.367
R770 B.n499 B.n497 163.367
R771 B.n165 B.t23 83.5406
R772 B.n71 B.t16 83.5406
R773 B.n159 B.t13 83.5208
R774 B.n64 B.t19 83.5208
R775 B.n166 B.t22 72.8739
R776 B.n72 B.t17 72.8739
R777 B.n160 B.t12 72.8542
R778 B.n65 B.t20 72.8542
R779 B.n411 B.n132 71.676
R780 B.n409 B.n134 71.676
R781 B.n405 B.n404 71.676
R782 B.n398 B.n136 71.676
R783 B.n397 B.n396 71.676
R784 B.n390 B.n138 71.676
R785 B.n389 B.n388 71.676
R786 B.n382 B.n140 71.676
R787 B.n381 B.n380 71.676
R788 B.n374 B.n142 71.676
R789 B.n373 B.n372 71.676
R790 B.n366 B.n144 71.676
R791 B.n365 B.n364 71.676
R792 B.n358 B.n146 71.676
R793 B.n357 B.n356 71.676
R794 B.n350 B.n148 71.676
R795 B.n349 B.n348 71.676
R796 B.n342 B.n150 71.676
R797 B.n341 B.n340 71.676
R798 B.n334 B.n152 71.676
R799 B.n333 B.n332 71.676
R800 B.n326 B.n154 71.676
R801 B.n325 B.n324 71.676
R802 B.n318 B.n156 71.676
R803 B.n317 B.n316 71.676
R804 B.n309 B.n158 71.676
R805 B.n308 B.n307 71.676
R806 B.n301 B.n162 71.676
R807 B.n300 B.n299 71.676
R808 B.n293 B.n164 71.676
R809 B.n292 B.n168 71.676
R810 B.n288 B.n287 71.676
R811 B.n281 B.n170 71.676
R812 B.n280 B.n279 71.676
R813 B.n273 B.n172 71.676
R814 B.n272 B.n271 71.676
R815 B.n265 B.n174 71.676
R816 B.n264 B.n263 71.676
R817 B.n257 B.n176 71.676
R818 B.n256 B.n255 71.676
R819 B.n249 B.n178 71.676
R820 B.n248 B.n247 71.676
R821 B.n241 B.n180 71.676
R822 B.n240 B.n239 71.676
R823 B.n233 B.n182 71.676
R824 B.n232 B.n231 71.676
R825 B.n225 B.n184 71.676
R826 B.n224 B.n223 71.676
R827 B.n217 B.n186 71.676
R828 B.n216 B.n215 71.676
R829 B.n209 B.n188 71.676
R830 B.n208 B.n207 71.676
R831 B.n201 B.n190 71.676
R832 B.n200 B.n199 71.676
R833 B.n193 B.n192 71.676
R834 B.n715 B.n37 71.676
R835 B.n714 B.n713 71.676
R836 B.n707 B.n39 71.676
R837 B.n706 B.n705 71.676
R838 B.n699 B.n41 71.676
R839 B.n698 B.n697 71.676
R840 B.n691 B.n43 71.676
R841 B.n690 B.n689 71.676
R842 B.n683 B.n45 71.676
R843 B.n682 B.n681 71.676
R844 B.n675 B.n47 71.676
R845 B.n674 B.n673 71.676
R846 B.n667 B.n49 71.676
R847 B.n666 B.n665 71.676
R848 B.n659 B.n51 71.676
R849 B.n658 B.n657 71.676
R850 B.n651 B.n53 71.676
R851 B.n650 B.n649 71.676
R852 B.n643 B.n55 71.676
R853 B.n642 B.n641 71.676
R854 B.n635 B.n57 71.676
R855 B.n634 B.n633 71.676
R856 B.n627 B.n59 71.676
R857 B.n626 B.n625 71.676
R858 B.n619 B.n61 71.676
R859 B.n618 B.n617 71.676
R860 B.n611 B.n63 71.676
R861 B.n610 B.n609 71.676
R862 B.n603 B.n68 71.676
R863 B.n602 B.n601 71.676
R864 B.n594 B.n70 71.676
R865 B.n593 B.n592 71.676
R866 B.n586 B.n74 71.676
R867 B.n585 B.n584 71.676
R868 B.n578 B.n76 71.676
R869 B.n577 B.n576 71.676
R870 B.n570 B.n78 71.676
R871 B.n569 B.n568 71.676
R872 B.n562 B.n80 71.676
R873 B.n561 B.n560 71.676
R874 B.n554 B.n82 71.676
R875 B.n553 B.n552 71.676
R876 B.n546 B.n84 71.676
R877 B.n545 B.n544 71.676
R878 B.n538 B.n86 71.676
R879 B.n537 B.n536 71.676
R880 B.n530 B.n88 71.676
R881 B.n529 B.n528 71.676
R882 B.n522 B.n90 71.676
R883 B.n521 B.n520 71.676
R884 B.n514 B.n92 71.676
R885 B.n513 B.n512 71.676
R886 B.n506 B.n94 71.676
R887 B.n505 B.n504 71.676
R888 B.n498 B.n96 71.676
R889 B.n497 B.n496 71.676
R890 B.n496 B.n495 71.676
R891 B.n499 B.n498 71.676
R892 B.n504 B.n503 71.676
R893 B.n507 B.n506 71.676
R894 B.n512 B.n511 71.676
R895 B.n515 B.n514 71.676
R896 B.n520 B.n519 71.676
R897 B.n523 B.n522 71.676
R898 B.n528 B.n527 71.676
R899 B.n531 B.n530 71.676
R900 B.n536 B.n535 71.676
R901 B.n539 B.n538 71.676
R902 B.n544 B.n543 71.676
R903 B.n547 B.n546 71.676
R904 B.n552 B.n551 71.676
R905 B.n555 B.n554 71.676
R906 B.n560 B.n559 71.676
R907 B.n563 B.n562 71.676
R908 B.n568 B.n567 71.676
R909 B.n571 B.n570 71.676
R910 B.n576 B.n575 71.676
R911 B.n579 B.n578 71.676
R912 B.n584 B.n583 71.676
R913 B.n587 B.n586 71.676
R914 B.n592 B.n591 71.676
R915 B.n595 B.n594 71.676
R916 B.n601 B.n600 71.676
R917 B.n604 B.n603 71.676
R918 B.n609 B.n608 71.676
R919 B.n612 B.n611 71.676
R920 B.n617 B.n616 71.676
R921 B.n620 B.n619 71.676
R922 B.n625 B.n624 71.676
R923 B.n628 B.n627 71.676
R924 B.n633 B.n632 71.676
R925 B.n636 B.n635 71.676
R926 B.n641 B.n640 71.676
R927 B.n644 B.n643 71.676
R928 B.n649 B.n648 71.676
R929 B.n652 B.n651 71.676
R930 B.n657 B.n656 71.676
R931 B.n660 B.n659 71.676
R932 B.n665 B.n664 71.676
R933 B.n668 B.n667 71.676
R934 B.n673 B.n672 71.676
R935 B.n676 B.n675 71.676
R936 B.n681 B.n680 71.676
R937 B.n684 B.n683 71.676
R938 B.n689 B.n688 71.676
R939 B.n692 B.n691 71.676
R940 B.n697 B.n696 71.676
R941 B.n700 B.n699 71.676
R942 B.n705 B.n704 71.676
R943 B.n708 B.n707 71.676
R944 B.n713 B.n712 71.676
R945 B.n716 B.n715 71.676
R946 B.n412 B.n411 71.676
R947 B.n406 B.n134 71.676
R948 B.n404 B.n403 71.676
R949 B.n399 B.n398 71.676
R950 B.n396 B.n395 71.676
R951 B.n391 B.n390 71.676
R952 B.n388 B.n387 71.676
R953 B.n383 B.n382 71.676
R954 B.n380 B.n379 71.676
R955 B.n375 B.n374 71.676
R956 B.n372 B.n371 71.676
R957 B.n367 B.n366 71.676
R958 B.n364 B.n363 71.676
R959 B.n359 B.n358 71.676
R960 B.n356 B.n355 71.676
R961 B.n351 B.n350 71.676
R962 B.n348 B.n347 71.676
R963 B.n343 B.n342 71.676
R964 B.n340 B.n339 71.676
R965 B.n335 B.n334 71.676
R966 B.n332 B.n331 71.676
R967 B.n327 B.n326 71.676
R968 B.n324 B.n323 71.676
R969 B.n319 B.n318 71.676
R970 B.n316 B.n315 71.676
R971 B.n310 B.n309 71.676
R972 B.n307 B.n306 71.676
R973 B.n302 B.n301 71.676
R974 B.n299 B.n298 71.676
R975 B.n294 B.n293 71.676
R976 B.n289 B.n168 71.676
R977 B.n287 B.n286 71.676
R978 B.n282 B.n281 71.676
R979 B.n279 B.n278 71.676
R980 B.n274 B.n273 71.676
R981 B.n271 B.n270 71.676
R982 B.n266 B.n265 71.676
R983 B.n263 B.n262 71.676
R984 B.n258 B.n257 71.676
R985 B.n255 B.n254 71.676
R986 B.n250 B.n249 71.676
R987 B.n247 B.n246 71.676
R988 B.n242 B.n241 71.676
R989 B.n239 B.n238 71.676
R990 B.n234 B.n233 71.676
R991 B.n231 B.n230 71.676
R992 B.n226 B.n225 71.676
R993 B.n223 B.n222 71.676
R994 B.n218 B.n217 71.676
R995 B.n215 B.n214 71.676
R996 B.n210 B.n209 71.676
R997 B.n207 B.n206 71.676
R998 B.n202 B.n201 71.676
R999 B.n199 B.n198 71.676
R1000 B.n194 B.n193 71.676
R1001 B.n167 B.n166 59.5399
R1002 B.n313 B.n160 59.5399
R1003 B.n66 B.n65 59.5399
R1004 B.n597 B.n72 59.5399
R1005 B.n417 B.n131 59.5179
R1006 B.n721 B.n36 59.5179
R1007 B.n417 B.n127 36.4616
R1008 B.n423 B.n127 36.4616
R1009 B.n423 B.n123 36.4616
R1010 B.n429 B.n123 36.4616
R1011 B.n435 B.n119 36.4616
R1012 B.n435 B.n114 36.4616
R1013 B.n441 B.n114 36.4616
R1014 B.n441 B.n115 36.4616
R1015 B.n453 B.n106 36.4616
R1016 B.n461 B.n460 36.4616
R1017 B.n467 B.n4 36.4616
R1018 B.n755 B.n4 36.4616
R1019 B.n755 B.n754 36.4616
R1020 B.n754 B.n753 36.4616
R1021 B.n747 B.n11 36.4616
R1022 B.n745 B.n15 36.4616
R1023 B.n738 B.n737 36.4616
R1024 B.n737 B.n22 36.4616
R1025 B.n731 B.n22 36.4616
R1026 B.n731 B.n730 36.4616
R1027 B.n729 B.n29 36.4616
R1028 B.n723 B.n29 36.4616
R1029 B.n723 B.n722 36.4616
R1030 B.n722 B.n721 36.4616
R1031 B.n107 B.t2 35.3892
R1032 B.t7 B.n746 35.3892
R1033 B.n447 B.t9 32.1721
R1034 B.n739 B.t6 32.1721
R1035 B.n719 B.n718 29.8151
R1036 B.n419 B.n129 29.8151
R1037 B.n415 B.n414 29.8151
R1038 B.n494 B.n493 29.8151
R1039 B.n447 B.t5 26.8102
R1040 B.n739 B.t0 26.8102
R1041 B.t11 B.n119 25.7378
R1042 B.n730 B.t15 25.7378
R1043 B.t1 B.n107 23.593
R1044 B.n746 B.t8 23.593
R1045 B.n460 B.t3 21.4482
R1046 B.n11 B.t4 21.4482
R1047 B B.n757 18.0485
R1048 B.n467 B.t3 15.0139
R1049 B.n753 B.t4 15.0139
R1050 B.n453 B.t1 12.8691
R1051 B.t8 B.n745 12.8691
R1052 B.n429 B.t11 10.7244
R1053 B.t15 B.n729 10.7244
R1054 B.n166 B.n165 10.6672
R1055 B.n160 B.n159 10.6672
R1056 B.n65 B.n64 10.6672
R1057 B.n72 B.n71 10.6672
R1058 B.n718 B.n717 10.6151
R1059 B.n717 B.n38 10.6151
R1060 B.n711 B.n38 10.6151
R1061 B.n711 B.n710 10.6151
R1062 B.n710 B.n709 10.6151
R1063 B.n709 B.n40 10.6151
R1064 B.n703 B.n40 10.6151
R1065 B.n703 B.n702 10.6151
R1066 B.n702 B.n701 10.6151
R1067 B.n701 B.n42 10.6151
R1068 B.n695 B.n42 10.6151
R1069 B.n695 B.n694 10.6151
R1070 B.n694 B.n693 10.6151
R1071 B.n693 B.n44 10.6151
R1072 B.n687 B.n44 10.6151
R1073 B.n687 B.n686 10.6151
R1074 B.n686 B.n685 10.6151
R1075 B.n685 B.n46 10.6151
R1076 B.n679 B.n46 10.6151
R1077 B.n679 B.n678 10.6151
R1078 B.n678 B.n677 10.6151
R1079 B.n677 B.n48 10.6151
R1080 B.n671 B.n48 10.6151
R1081 B.n671 B.n670 10.6151
R1082 B.n670 B.n669 10.6151
R1083 B.n669 B.n50 10.6151
R1084 B.n663 B.n50 10.6151
R1085 B.n663 B.n662 10.6151
R1086 B.n662 B.n661 10.6151
R1087 B.n661 B.n52 10.6151
R1088 B.n655 B.n52 10.6151
R1089 B.n655 B.n654 10.6151
R1090 B.n654 B.n653 10.6151
R1091 B.n653 B.n54 10.6151
R1092 B.n647 B.n54 10.6151
R1093 B.n647 B.n646 10.6151
R1094 B.n646 B.n645 10.6151
R1095 B.n645 B.n56 10.6151
R1096 B.n639 B.n56 10.6151
R1097 B.n639 B.n638 10.6151
R1098 B.n638 B.n637 10.6151
R1099 B.n637 B.n58 10.6151
R1100 B.n631 B.n58 10.6151
R1101 B.n631 B.n630 10.6151
R1102 B.n630 B.n629 10.6151
R1103 B.n629 B.n60 10.6151
R1104 B.n623 B.n60 10.6151
R1105 B.n623 B.n622 10.6151
R1106 B.n622 B.n621 10.6151
R1107 B.n621 B.n62 10.6151
R1108 B.n615 B.n614 10.6151
R1109 B.n614 B.n613 10.6151
R1110 B.n613 B.n67 10.6151
R1111 B.n607 B.n67 10.6151
R1112 B.n607 B.n606 10.6151
R1113 B.n606 B.n605 10.6151
R1114 B.n605 B.n69 10.6151
R1115 B.n599 B.n69 10.6151
R1116 B.n599 B.n598 10.6151
R1117 B.n596 B.n73 10.6151
R1118 B.n590 B.n73 10.6151
R1119 B.n590 B.n589 10.6151
R1120 B.n589 B.n588 10.6151
R1121 B.n588 B.n75 10.6151
R1122 B.n582 B.n75 10.6151
R1123 B.n582 B.n581 10.6151
R1124 B.n581 B.n580 10.6151
R1125 B.n580 B.n77 10.6151
R1126 B.n574 B.n77 10.6151
R1127 B.n574 B.n573 10.6151
R1128 B.n573 B.n572 10.6151
R1129 B.n572 B.n79 10.6151
R1130 B.n566 B.n79 10.6151
R1131 B.n566 B.n565 10.6151
R1132 B.n565 B.n564 10.6151
R1133 B.n564 B.n81 10.6151
R1134 B.n558 B.n81 10.6151
R1135 B.n558 B.n557 10.6151
R1136 B.n557 B.n556 10.6151
R1137 B.n556 B.n83 10.6151
R1138 B.n550 B.n83 10.6151
R1139 B.n550 B.n549 10.6151
R1140 B.n549 B.n548 10.6151
R1141 B.n548 B.n85 10.6151
R1142 B.n542 B.n85 10.6151
R1143 B.n542 B.n541 10.6151
R1144 B.n541 B.n540 10.6151
R1145 B.n540 B.n87 10.6151
R1146 B.n534 B.n87 10.6151
R1147 B.n534 B.n533 10.6151
R1148 B.n533 B.n532 10.6151
R1149 B.n532 B.n89 10.6151
R1150 B.n526 B.n89 10.6151
R1151 B.n526 B.n525 10.6151
R1152 B.n525 B.n524 10.6151
R1153 B.n524 B.n91 10.6151
R1154 B.n518 B.n91 10.6151
R1155 B.n518 B.n517 10.6151
R1156 B.n517 B.n516 10.6151
R1157 B.n516 B.n93 10.6151
R1158 B.n510 B.n93 10.6151
R1159 B.n510 B.n509 10.6151
R1160 B.n509 B.n508 10.6151
R1161 B.n508 B.n95 10.6151
R1162 B.n502 B.n95 10.6151
R1163 B.n502 B.n501 10.6151
R1164 B.n501 B.n500 10.6151
R1165 B.n500 B.n97 10.6151
R1166 B.n494 B.n97 10.6151
R1167 B.n420 B.n419 10.6151
R1168 B.n421 B.n420 10.6151
R1169 B.n421 B.n121 10.6151
R1170 B.n431 B.n121 10.6151
R1171 B.n432 B.n431 10.6151
R1172 B.n433 B.n432 10.6151
R1173 B.n433 B.n112 10.6151
R1174 B.n443 B.n112 10.6151
R1175 B.n444 B.n443 10.6151
R1176 B.n445 B.n444 10.6151
R1177 B.n445 B.n104 10.6151
R1178 B.n455 B.n104 10.6151
R1179 B.n456 B.n455 10.6151
R1180 B.n458 B.n456 10.6151
R1181 B.n458 B.n457 10.6151
R1182 B.n457 B.n98 10.6151
R1183 B.n470 B.n98 10.6151
R1184 B.n471 B.n470 10.6151
R1185 B.n472 B.n471 10.6151
R1186 B.n473 B.n472 10.6151
R1187 B.n475 B.n473 10.6151
R1188 B.n476 B.n475 10.6151
R1189 B.n477 B.n476 10.6151
R1190 B.n478 B.n477 10.6151
R1191 B.n480 B.n478 10.6151
R1192 B.n481 B.n480 10.6151
R1193 B.n482 B.n481 10.6151
R1194 B.n483 B.n482 10.6151
R1195 B.n485 B.n483 10.6151
R1196 B.n486 B.n485 10.6151
R1197 B.n487 B.n486 10.6151
R1198 B.n488 B.n487 10.6151
R1199 B.n490 B.n488 10.6151
R1200 B.n491 B.n490 10.6151
R1201 B.n492 B.n491 10.6151
R1202 B.n493 B.n492 10.6151
R1203 B.n414 B.n413 10.6151
R1204 B.n413 B.n133 10.6151
R1205 B.n408 B.n133 10.6151
R1206 B.n408 B.n407 10.6151
R1207 B.n407 B.n135 10.6151
R1208 B.n402 B.n135 10.6151
R1209 B.n402 B.n401 10.6151
R1210 B.n401 B.n400 10.6151
R1211 B.n400 B.n137 10.6151
R1212 B.n394 B.n137 10.6151
R1213 B.n394 B.n393 10.6151
R1214 B.n393 B.n392 10.6151
R1215 B.n392 B.n139 10.6151
R1216 B.n386 B.n139 10.6151
R1217 B.n386 B.n385 10.6151
R1218 B.n385 B.n384 10.6151
R1219 B.n384 B.n141 10.6151
R1220 B.n378 B.n141 10.6151
R1221 B.n378 B.n377 10.6151
R1222 B.n377 B.n376 10.6151
R1223 B.n376 B.n143 10.6151
R1224 B.n370 B.n143 10.6151
R1225 B.n370 B.n369 10.6151
R1226 B.n369 B.n368 10.6151
R1227 B.n368 B.n145 10.6151
R1228 B.n362 B.n145 10.6151
R1229 B.n362 B.n361 10.6151
R1230 B.n361 B.n360 10.6151
R1231 B.n360 B.n147 10.6151
R1232 B.n354 B.n147 10.6151
R1233 B.n354 B.n353 10.6151
R1234 B.n353 B.n352 10.6151
R1235 B.n352 B.n149 10.6151
R1236 B.n346 B.n149 10.6151
R1237 B.n346 B.n345 10.6151
R1238 B.n345 B.n344 10.6151
R1239 B.n344 B.n151 10.6151
R1240 B.n338 B.n151 10.6151
R1241 B.n338 B.n337 10.6151
R1242 B.n337 B.n336 10.6151
R1243 B.n336 B.n153 10.6151
R1244 B.n330 B.n153 10.6151
R1245 B.n330 B.n329 10.6151
R1246 B.n329 B.n328 10.6151
R1247 B.n328 B.n155 10.6151
R1248 B.n322 B.n155 10.6151
R1249 B.n322 B.n321 10.6151
R1250 B.n321 B.n320 10.6151
R1251 B.n320 B.n157 10.6151
R1252 B.n314 B.n157 10.6151
R1253 B.n312 B.n311 10.6151
R1254 B.n311 B.n161 10.6151
R1255 B.n305 B.n161 10.6151
R1256 B.n305 B.n304 10.6151
R1257 B.n304 B.n303 10.6151
R1258 B.n303 B.n163 10.6151
R1259 B.n297 B.n163 10.6151
R1260 B.n297 B.n296 10.6151
R1261 B.n296 B.n295 10.6151
R1262 B.n291 B.n290 10.6151
R1263 B.n290 B.n169 10.6151
R1264 B.n285 B.n169 10.6151
R1265 B.n285 B.n284 10.6151
R1266 B.n284 B.n283 10.6151
R1267 B.n283 B.n171 10.6151
R1268 B.n277 B.n171 10.6151
R1269 B.n277 B.n276 10.6151
R1270 B.n276 B.n275 10.6151
R1271 B.n275 B.n173 10.6151
R1272 B.n269 B.n173 10.6151
R1273 B.n269 B.n268 10.6151
R1274 B.n268 B.n267 10.6151
R1275 B.n267 B.n175 10.6151
R1276 B.n261 B.n175 10.6151
R1277 B.n261 B.n260 10.6151
R1278 B.n260 B.n259 10.6151
R1279 B.n259 B.n177 10.6151
R1280 B.n253 B.n177 10.6151
R1281 B.n253 B.n252 10.6151
R1282 B.n252 B.n251 10.6151
R1283 B.n251 B.n179 10.6151
R1284 B.n245 B.n179 10.6151
R1285 B.n245 B.n244 10.6151
R1286 B.n244 B.n243 10.6151
R1287 B.n243 B.n181 10.6151
R1288 B.n237 B.n181 10.6151
R1289 B.n237 B.n236 10.6151
R1290 B.n236 B.n235 10.6151
R1291 B.n235 B.n183 10.6151
R1292 B.n229 B.n183 10.6151
R1293 B.n229 B.n228 10.6151
R1294 B.n228 B.n227 10.6151
R1295 B.n227 B.n185 10.6151
R1296 B.n221 B.n185 10.6151
R1297 B.n221 B.n220 10.6151
R1298 B.n220 B.n219 10.6151
R1299 B.n219 B.n187 10.6151
R1300 B.n213 B.n187 10.6151
R1301 B.n213 B.n212 10.6151
R1302 B.n212 B.n211 10.6151
R1303 B.n211 B.n189 10.6151
R1304 B.n205 B.n189 10.6151
R1305 B.n205 B.n204 10.6151
R1306 B.n204 B.n203 10.6151
R1307 B.n203 B.n191 10.6151
R1308 B.n197 B.n191 10.6151
R1309 B.n197 B.n196 10.6151
R1310 B.n196 B.n195 10.6151
R1311 B.n195 B.n129 10.6151
R1312 B.n415 B.n125 10.6151
R1313 B.n425 B.n125 10.6151
R1314 B.n426 B.n425 10.6151
R1315 B.n427 B.n426 10.6151
R1316 B.n427 B.n117 10.6151
R1317 B.n437 B.n117 10.6151
R1318 B.n438 B.n437 10.6151
R1319 B.n439 B.n438 10.6151
R1320 B.n439 B.n109 10.6151
R1321 B.n449 B.n109 10.6151
R1322 B.n450 B.n449 10.6151
R1323 B.n451 B.n450 10.6151
R1324 B.n451 B.n101 10.6151
R1325 B.n463 B.n101 10.6151
R1326 B.n464 B.n463 10.6151
R1327 B.n465 B.n464 10.6151
R1328 B.n465 B.n0 10.6151
R1329 B.n751 B.n1 10.6151
R1330 B.n751 B.n750 10.6151
R1331 B.n750 B.n749 10.6151
R1332 B.n749 B.n9 10.6151
R1333 B.n743 B.n9 10.6151
R1334 B.n743 B.n742 10.6151
R1335 B.n742 B.n741 10.6151
R1336 B.n741 B.n17 10.6151
R1337 B.n735 B.n17 10.6151
R1338 B.n735 B.n734 10.6151
R1339 B.n734 B.n733 10.6151
R1340 B.n733 B.n24 10.6151
R1341 B.n727 B.n24 10.6151
R1342 B.n727 B.n726 10.6151
R1343 B.n726 B.n725 10.6151
R1344 B.n725 B.n31 10.6151
R1345 B.n719 B.n31 10.6151
R1346 B.t5 B.n106 9.65197
R1347 B.t0 B.n15 9.65197
R1348 B.n66 B.n62 9.36635
R1349 B.n597 B.n596 9.36635
R1350 B.n314 B.n313 9.36635
R1351 B.n291 B.n167 9.36635
R1352 B.n115 B.t9 4.29004
R1353 B.t6 B.n738 4.29004
R1354 B.n757 B.n0 2.81026
R1355 B.n757 B.n1 2.81026
R1356 B.n615 B.n66 1.24928
R1357 B.n598 B.n597 1.24928
R1358 B.n313 B.n312 1.24928
R1359 B.n295 B.n167 1.24928
R1360 B.n461 B.t2 1.07289
R1361 B.n747 B.t7 1.07289
R1362 VP.n19 VP.t5 1863
R1363 VP.n12 VP.t3 1863
R1364 VP.n4 VP.t0 1863
R1365 VP.n10 VP.t1 1863
R1366 VP.n18 VP.t2 1811.88
R1367 VP.n16 VP.t9 1811.88
R1368 VP.n1 VP.t6 1811.88
R1369 VP.n3 VP.t7 1811.88
R1370 VP.n7 VP.t4 1811.88
R1371 VP.n9 VP.t8 1811.88
R1372 VP.n5 VP.n4 161.489
R1373 VP.n20 VP.n19 161.3
R1374 VP.n6 VP.n5 161.3
R1375 VP.n8 VP.n2 161.3
R1376 VP.n11 VP.n10 161.3
R1377 VP.n17 VP.n0 161.3
R1378 VP.n15 VP.n14 161.3
R1379 VP.n13 VP.n12 161.3
R1380 VP.n15 VP.n1 43.8187
R1381 VP.n18 VP.n17 43.8187
R1382 VP.n6 VP.n3 43.8187
R1383 VP.n9 VP.n8 43.8187
R1384 VP.n13 VP.n11 42.7316
R1385 VP.n16 VP.n15 36.5157
R1386 VP.n17 VP.n16 36.5157
R1387 VP.n7 VP.n6 36.5157
R1388 VP.n8 VP.n7 36.5157
R1389 VP.n12 VP.n1 29.2126
R1390 VP.n19 VP.n18 29.2126
R1391 VP.n4 VP.n3 29.2126
R1392 VP.n10 VP.n9 29.2126
R1393 VP.n5 VP.n2 0.189894
R1394 VP.n11 VP.n2 0.189894
R1395 VP.n14 VP.n13 0.189894
R1396 VP.n14 VP.n0 0.189894
R1397 VP.n20 VP.n0 0.189894
R1398 VP VP.n20 0.0516364
R1399 VDD1.n1 VDD1.t9 60.7206
R1400 VDD1.n3 VDD1.t6 60.7204
R1401 VDD1.n5 VDD1.n4 59.2473
R1402 VDD1.n7 VDD1.n6 58.9473
R1403 VDD1.n1 VDD1.n0 58.9473
R1404 VDD1.n3 VDD1.n2 58.9471
R1405 VDD1.n7 VDD1.n5 39.9255
R1406 VDD1.n6 VDD1.t1 1.29971
R1407 VDD1.n6 VDD1.t8 1.29971
R1408 VDD1.n0 VDD1.t2 1.29971
R1409 VDD1.n0 VDD1.t5 1.29971
R1410 VDD1.n4 VDD1.t7 1.29971
R1411 VDD1.n4 VDD1.t4 1.29971
R1412 VDD1.n2 VDD1.t3 1.29971
R1413 VDD1.n2 VDD1.t0 1.29971
R1414 VDD1 VDD1.n7 0.297914
R1415 VDD1 VDD1.n1 0.177224
R1416 VDD1.n5 VDD1.n3 0.0636885
C0 VDD1 VDD2 0.677382f
C1 VTAIL VN 3.4411f
C2 VP VN 5.48587f
C3 VTAIL VDD2 29.756699f
C4 VDD2 VP 0.281262f
C5 VDD1 VTAIL 29.730501f
C6 VDD2 VN 4.02785f
C7 VDD1 VP 4.15447f
C8 VTAIL VP 3.45609f
C9 VDD1 VN 0.14795f
C10 VDD2 B 5.050187f
C11 VDD1 B 4.856892f
C12 VTAIL B 7.03112f
C13 VN B 7.9304f
C14 VP B 5.408829f
C15 VDD1.t9 B 4.55761f
C16 VDD1.t2 B 0.395646f
C17 VDD1.t5 B 0.395646f
C18 VDD1.n0 B 3.56682f
C19 VDD1.n1 B 0.783384f
C20 VDD1.t6 B 4.55759f
C21 VDD1.t3 B 0.395646f
C22 VDD1.t0 B 0.395646f
C23 VDD1.n2 B 3.56681f
C24 VDD1.n3 B 0.783444f
C25 VDD1.t7 B 0.395646f
C26 VDD1.t4 B 0.395646f
C27 VDD1.n4 B 3.56873f
C28 VDD1.n5 B 2.51655f
C29 VDD1.t1 B 0.395646f
C30 VDD1.t8 B 0.395646f
C31 VDD1.n6 B 3.56682f
C32 VDD1.n7 B 3.21687f
C33 VP.n0 B 0.058141f
C34 VP.t2 B 0.549883f
C35 VP.t9 B 0.549883f
C36 VP.t6 B 0.549883f
C37 VP.n1 B 0.215556f
C38 VP.n2 B 0.058141f
C39 VP.t8 B 0.549883f
C40 VP.t4 B 0.549883f
C41 VP.t7 B 0.549883f
C42 VP.n3 B 0.215556f
C43 VP.t0 B 0.555867f
C44 VP.n4 B 0.233247f
C45 VP.n5 B 0.131251f
C46 VP.n6 B 0.02108f
C47 VP.n7 B 0.215556f
C48 VP.n8 B 0.02108f
C49 VP.n9 B 0.215556f
C50 VP.t1 B 0.555867f
C51 VP.n10 B 0.233161f
C52 VP.n11 B 2.46946f
C53 VP.t3 B 0.555867f
C54 VP.n12 B 0.233161f
C55 VP.n13 B 2.51851f
C56 VP.n14 B 0.058141f
C57 VP.n15 B 0.02108f
C58 VP.n16 B 0.215556f
C59 VP.n17 B 0.02108f
C60 VP.n18 B 0.215556f
C61 VP.t5 B 0.555867f
C62 VP.n19 B 0.233161f
C63 VP.n20 B 0.045057f
C64 VTAIL.t11 B 0.403913f
C65 VTAIL.t16 B 0.403913f
C66 VTAIL.n0 B 3.53049f
C67 VTAIL.n1 B 0.47367f
C68 VTAIL.t3 B 4.50598f
C69 VTAIL.n2 B 0.606288f
C70 VTAIL.t1 B 0.403913f
C71 VTAIL.t2 B 0.403913f
C72 VTAIL.n3 B 3.53049f
C73 VTAIL.n4 B 0.455038f
C74 VTAIL.t9 B 0.403913f
C75 VTAIL.t5 B 0.403913f
C76 VTAIL.n5 B 3.53049f
C77 VTAIL.n6 B 2.38168f
C78 VTAIL.t15 B 0.403913f
C79 VTAIL.t10 B 0.403913f
C80 VTAIL.n7 B 3.5305f
C81 VTAIL.n8 B 2.38167f
C82 VTAIL.t14 B 0.403913f
C83 VTAIL.t19 B 0.403913f
C84 VTAIL.n9 B 3.5305f
C85 VTAIL.n10 B 0.455027f
C86 VTAIL.t13 B 4.506f
C87 VTAIL.n11 B 0.606261f
C88 VTAIL.t4 B 0.403913f
C89 VTAIL.t7 B 0.403913f
C90 VTAIL.n12 B 3.5305f
C91 VTAIL.n13 B 0.480181f
C92 VTAIL.t8 B 0.403913f
C93 VTAIL.t0 B 0.403913f
C94 VTAIL.n14 B 3.5305f
C95 VTAIL.n15 B 0.455027f
C96 VTAIL.t6 B 4.506f
C97 VTAIL.n16 B 2.45652f
C98 VTAIL.t12 B 4.50598f
C99 VTAIL.n17 B 2.45654f
C100 VTAIL.t17 B 0.403913f
C101 VTAIL.t18 B 0.403913f
C102 VTAIL.n18 B 3.53049f
C103 VTAIL.n19 B 0.410319f
C104 VDD2.t4 B 4.56047f
C105 VDD2.t5 B 0.395896f
C106 VDD2.t3 B 0.395896f
C107 VDD2.n0 B 3.56906f
C108 VDD2.n1 B 0.783939f
C109 VDD2.t2 B 0.395896f
C110 VDD2.t1 B 0.395896f
C111 VDD2.n2 B 3.57099f
C112 VDD2.n3 B 2.43073f
C113 VDD2.t7 B 4.55708f
C114 VDD2.n4 B 3.24511f
C115 VDD2.t6 B 0.395896f
C116 VDD2.t8 B 0.395896f
C117 VDD2.n5 B 3.56907f
C118 VDD2.n6 B 0.35053f
C119 VDD2.t9 B 0.395896f
C120 VDD2.t0 B 0.395896f
C121 VDD2.n7 B 3.57096f
C122 VN.n0 B 0.05647f
C123 VN.t1 B 0.534079f
C124 VN.t2 B 0.534079f
C125 VN.t3 B 0.534079f
C126 VN.n1 B 0.209361f
C127 VN.t8 B 0.539891f
C128 VN.n2 B 0.226543f
C129 VN.n3 B 0.127479f
C130 VN.n4 B 0.020474f
C131 VN.n5 B 0.209361f
C132 VN.n6 B 0.020474f
C133 VN.n7 B 0.209361f
C134 VN.t7 B 0.539891f
C135 VN.n8 B 0.22646f
C136 VN.n9 B 0.043762f
C137 VN.n10 B 0.05647f
C138 VN.t4 B 0.539891f
C139 VN.t9 B 0.534079f
C140 VN.t5 B 0.534079f
C141 VN.t0 B 0.534079f
C142 VN.n11 B 0.209361f
C143 VN.t6 B 0.539891f
C144 VN.n12 B 0.226543f
C145 VN.n13 B 0.127479f
C146 VN.n14 B 0.020474f
C147 VN.n15 B 0.209361f
C148 VN.n16 B 0.020474f
C149 VN.n17 B 0.209361f
C150 VN.n18 B 0.22646f
C151 VN.n19 B 2.43552f
.ends

