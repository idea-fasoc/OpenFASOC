* NGSPICE file created from diff_pair_sample_0134.ext - technology: sky130A

.subckt diff_pair_sample_0134 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X1 VTAIL.t6 VP.t0 VDD1.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X2 VDD2.t4 VN.t1 VTAIL.t18 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=1.28865 ps=8.14 w=7.81 l=2.81
X3 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=0 ps=0 w=7.81 l=2.81
X4 VTAIL.t2 VP.t1 VDD1.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X5 VDD1.t7 VP.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=1.28865 ps=8.14 w=7.81 l=2.81
X6 VDD1.t6 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=3.0459 ps=16.4 w=7.81 l=2.81
X7 VDD2.t3 VN.t2 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X8 VDD1.t5 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=3.0459 ps=16.4 w=7.81 l=2.81
X9 VDD1.t4 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X10 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=0 ps=0 w=7.81 l=2.81
X11 VDD2.t1 VN.t3 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=1.28865 ps=8.14 w=7.81 l=2.81
X12 VTAIL.t15 VN.t4 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X13 VTAIL.t7 VP.t6 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=0 ps=0 w=7.81 l=2.81
X15 VTAIL.t0 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X16 VTAIL.t14 VN.t5 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X17 VDD2.t5 VN.t6 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=3.0459 ps=16.4 w=7.81 l=2.81
X18 VTAIL.t12 VN.t7 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=0 ps=0 w=7.81 l=2.81
X20 VDD1.t1 VP.t8 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0459 pd=16.4 as=1.28865 ps=8.14 w=7.81 l=2.81
X21 VDD1.t0 VP.t9 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X22 VDD2.t7 VN.t8 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=1.28865 ps=8.14 w=7.81 l=2.81
X23 VDD2.t9 VN.t9 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.28865 pd=8.14 as=3.0459 ps=16.4 w=7.81 l=2.81
R0 VN.n85 VN.n44 161.3
R1 VN.n84 VN.n83 161.3
R2 VN.n82 VN.n45 161.3
R3 VN.n81 VN.n80 161.3
R4 VN.n79 VN.n46 161.3
R5 VN.n78 VN.n77 161.3
R6 VN.n76 VN.n47 161.3
R7 VN.n75 VN.n74 161.3
R8 VN.n73 VN.n48 161.3
R9 VN.n72 VN.n71 161.3
R10 VN.n70 VN.n50 161.3
R11 VN.n69 VN.n68 161.3
R12 VN.n67 VN.n51 161.3
R13 VN.n65 VN.n64 161.3
R14 VN.n63 VN.n52 161.3
R15 VN.n62 VN.n61 161.3
R16 VN.n60 VN.n53 161.3
R17 VN.n59 VN.n58 161.3
R18 VN.n57 VN.n54 161.3
R19 VN.n41 VN.n0 161.3
R20 VN.n40 VN.n39 161.3
R21 VN.n38 VN.n1 161.3
R22 VN.n37 VN.n36 161.3
R23 VN.n35 VN.n2 161.3
R24 VN.n34 VN.n33 161.3
R25 VN.n32 VN.n3 161.3
R26 VN.n31 VN.n30 161.3
R27 VN.n28 VN.n4 161.3
R28 VN.n27 VN.n26 161.3
R29 VN.n25 VN.n5 161.3
R30 VN.n24 VN.n23 161.3
R31 VN.n22 VN.n6 161.3
R32 VN.n20 VN.n19 161.3
R33 VN.n18 VN.n7 161.3
R34 VN.n17 VN.n16 161.3
R35 VN.n15 VN.n8 161.3
R36 VN.n14 VN.n13 161.3
R37 VN.n12 VN.n9 161.3
R38 VN.n43 VN.n42 109.288
R39 VN.n87 VN.n86 109.288
R40 VN.n11 VN.t3 99.6097
R41 VN.n56 VN.t6 99.6097
R42 VN.n10 VN.t5 66.9831
R43 VN.n21 VN.t2 66.9831
R44 VN.n29 VN.t4 66.9831
R45 VN.n42 VN.t9 66.9831
R46 VN.n55 VN.t7 66.9831
R47 VN.n66 VN.t8 66.9831
R48 VN.n49 VN.t0 66.9831
R49 VN.n86 VN.t1 66.9831
R50 VN.n16 VN.n15 56.5193
R51 VN.n61 VN.n60 56.5193
R52 VN.n27 VN.n5 56.5193
R53 VN.n72 VN.n50 56.5193
R54 VN.n11 VN.n10 54.5315
R55 VN.n56 VN.n55 54.5315
R56 VN VN.n87 51.3012
R57 VN.n36 VN.n35 44.3785
R58 VN.n80 VN.n79 44.3785
R59 VN.n36 VN.n1 36.6083
R60 VN.n80 VN.n45 36.6083
R61 VN.n14 VN.n9 24.4675
R62 VN.n15 VN.n14 24.4675
R63 VN.n16 VN.n7 24.4675
R64 VN.n20 VN.n7 24.4675
R65 VN.n23 VN.n22 24.4675
R66 VN.n23 VN.n5 24.4675
R67 VN.n28 VN.n27 24.4675
R68 VN.n30 VN.n28 24.4675
R69 VN.n34 VN.n3 24.4675
R70 VN.n35 VN.n34 24.4675
R71 VN.n40 VN.n1 24.4675
R72 VN.n41 VN.n40 24.4675
R73 VN.n60 VN.n59 24.4675
R74 VN.n59 VN.n54 24.4675
R75 VN.n68 VN.n50 24.4675
R76 VN.n68 VN.n67 24.4675
R77 VN.n65 VN.n52 24.4675
R78 VN.n61 VN.n52 24.4675
R79 VN.n79 VN.n78 24.4675
R80 VN.n78 VN.n47 24.4675
R81 VN.n74 VN.n73 24.4675
R82 VN.n73 VN.n72 24.4675
R83 VN.n85 VN.n84 24.4675
R84 VN.n84 VN.n45 24.4675
R85 VN.n10 VN.n9 19.0848
R86 VN.n30 VN.n29 19.0848
R87 VN.n55 VN.n54 19.0848
R88 VN.n74 VN.n49 19.0848
R89 VN.n21 VN.n20 12.234
R90 VN.n22 VN.n21 12.234
R91 VN.n67 VN.n66 12.234
R92 VN.n66 VN.n65 12.234
R93 VN.n29 VN.n3 5.38324
R94 VN.n49 VN.n47 5.38324
R95 VN.n57 VN.n56 5.13245
R96 VN.n12 VN.n11 5.13245
R97 VN.n42 VN.n41 1.46852
R98 VN.n86 VN.n85 1.46852
R99 VN.n87 VN.n44 0.278367
R100 VN.n43 VN.n0 0.278367
R101 VN.n83 VN.n44 0.189894
R102 VN.n83 VN.n82 0.189894
R103 VN.n82 VN.n81 0.189894
R104 VN.n81 VN.n46 0.189894
R105 VN.n77 VN.n46 0.189894
R106 VN.n77 VN.n76 0.189894
R107 VN.n76 VN.n75 0.189894
R108 VN.n75 VN.n48 0.189894
R109 VN.n71 VN.n48 0.189894
R110 VN.n71 VN.n70 0.189894
R111 VN.n70 VN.n69 0.189894
R112 VN.n69 VN.n51 0.189894
R113 VN.n64 VN.n51 0.189894
R114 VN.n64 VN.n63 0.189894
R115 VN.n63 VN.n62 0.189894
R116 VN.n62 VN.n53 0.189894
R117 VN.n58 VN.n53 0.189894
R118 VN.n58 VN.n57 0.189894
R119 VN.n13 VN.n12 0.189894
R120 VN.n13 VN.n8 0.189894
R121 VN.n17 VN.n8 0.189894
R122 VN.n18 VN.n17 0.189894
R123 VN.n19 VN.n18 0.189894
R124 VN.n19 VN.n6 0.189894
R125 VN.n24 VN.n6 0.189894
R126 VN.n25 VN.n24 0.189894
R127 VN.n26 VN.n25 0.189894
R128 VN.n26 VN.n4 0.189894
R129 VN.n31 VN.n4 0.189894
R130 VN.n32 VN.n31 0.189894
R131 VN.n33 VN.n32 0.189894
R132 VN.n33 VN.n2 0.189894
R133 VN.n37 VN.n2 0.189894
R134 VN.n38 VN.n37 0.189894
R135 VN.n39 VN.n38 0.189894
R136 VN.n39 VN.n0 0.189894
R137 VN VN.n43 0.153454
R138 VDD2.n1 VDD2.t1 70.2685
R139 VDD2.n4 VDD2.t4 67.5617
R140 VDD2.n3 VDD2.n2 67.0013
R141 VDD2 VDD2.n7 66.9985
R142 VDD2.n6 VDD2.n5 65.0266
R143 VDD2.n1 VDD2.n0 65.0265
R144 VDD2.n4 VDD2.n3 43.3058
R145 VDD2.n6 VDD2.n4 2.7074
R146 VDD2.n7 VDD2.t8 2.53571
R147 VDD2.n7 VDD2.t5 2.53571
R148 VDD2.n5 VDD2.t2 2.53571
R149 VDD2.n5 VDD2.t7 2.53571
R150 VDD2.n2 VDD2.t0 2.53571
R151 VDD2.n2 VDD2.t9 2.53571
R152 VDD2.n0 VDD2.t6 2.53571
R153 VDD2.n0 VDD2.t3 2.53571
R154 VDD2 VDD2.n6 0.735414
R155 VDD2.n3 VDD2.n1 0.621878
R156 VTAIL.n16 VTAIL.t4 50.883
R157 VTAIL.n11 VTAIL.t13 50.8829
R158 VTAIL.n17 VTAIL.t10 50.8828
R159 VTAIL.n2 VTAIL.t1 50.8828
R160 VTAIL.n15 VTAIL.n14 48.3478
R161 VTAIL.n13 VTAIL.n12 48.3478
R162 VTAIL.n10 VTAIL.n9 48.3478
R163 VTAIL.n8 VTAIL.n7 48.3478
R164 VTAIL.n19 VTAIL.n18 48.3477
R165 VTAIL.n1 VTAIL.n0 48.3477
R166 VTAIL.n4 VTAIL.n3 48.3477
R167 VTAIL.n6 VTAIL.n5 48.3477
R168 VTAIL.n8 VTAIL.n6 24.5134
R169 VTAIL.n17 VTAIL.n16 21.8065
R170 VTAIL.n10 VTAIL.n8 2.7074
R171 VTAIL.n11 VTAIL.n10 2.7074
R172 VTAIL.n15 VTAIL.n13 2.7074
R173 VTAIL.n16 VTAIL.n15 2.7074
R174 VTAIL.n6 VTAIL.n4 2.7074
R175 VTAIL.n4 VTAIL.n2 2.7074
R176 VTAIL.n19 VTAIL.n17 2.7074
R177 VTAIL.n18 VTAIL.t17 2.53571
R178 VTAIL.n18 VTAIL.t15 2.53571
R179 VTAIL.n0 VTAIL.t16 2.53571
R180 VTAIL.n0 VTAIL.t14 2.53571
R181 VTAIL.n3 VTAIL.t3 2.53571
R182 VTAIL.n3 VTAIL.t0 2.53571
R183 VTAIL.n5 VTAIL.t9 2.53571
R184 VTAIL.n5 VTAIL.t7 2.53571
R185 VTAIL.n14 VTAIL.t5 2.53571
R186 VTAIL.n14 VTAIL.t6 2.53571
R187 VTAIL.n12 VTAIL.t8 2.53571
R188 VTAIL.n12 VTAIL.t2 2.53571
R189 VTAIL.n9 VTAIL.t11 2.53571
R190 VTAIL.n9 VTAIL.t12 2.53571
R191 VTAIL.n7 VTAIL.t18 2.53571
R192 VTAIL.n7 VTAIL.t19 2.53571
R193 VTAIL VTAIL.n1 2.08886
R194 VTAIL.n13 VTAIL.n11 1.82378
R195 VTAIL.n2 VTAIL.n1 1.82378
R196 VTAIL VTAIL.n19 0.619035
R197 B.n857 B.n856 585
R198 B.n286 B.n150 585
R199 B.n285 B.n284 585
R200 B.n283 B.n282 585
R201 B.n281 B.n280 585
R202 B.n279 B.n278 585
R203 B.n277 B.n276 585
R204 B.n275 B.n274 585
R205 B.n273 B.n272 585
R206 B.n271 B.n270 585
R207 B.n269 B.n268 585
R208 B.n267 B.n266 585
R209 B.n265 B.n264 585
R210 B.n263 B.n262 585
R211 B.n261 B.n260 585
R212 B.n259 B.n258 585
R213 B.n257 B.n256 585
R214 B.n255 B.n254 585
R215 B.n253 B.n252 585
R216 B.n251 B.n250 585
R217 B.n249 B.n248 585
R218 B.n247 B.n246 585
R219 B.n245 B.n244 585
R220 B.n243 B.n242 585
R221 B.n241 B.n240 585
R222 B.n239 B.n238 585
R223 B.n237 B.n236 585
R224 B.n235 B.n234 585
R225 B.n233 B.n232 585
R226 B.n230 B.n229 585
R227 B.n228 B.n227 585
R228 B.n226 B.n225 585
R229 B.n224 B.n223 585
R230 B.n222 B.n221 585
R231 B.n220 B.n219 585
R232 B.n218 B.n217 585
R233 B.n216 B.n215 585
R234 B.n214 B.n213 585
R235 B.n212 B.n211 585
R236 B.n209 B.n208 585
R237 B.n207 B.n206 585
R238 B.n205 B.n204 585
R239 B.n203 B.n202 585
R240 B.n201 B.n200 585
R241 B.n199 B.n198 585
R242 B.n197 B.n196 585
R243 B.n195 B.n194 585
R244 B.n193 B.n192 585
R245 B.n191 B.n190 585
R246 B.n189 B.n188 585
R247 B.n187 B.n186 585
R248 B.n185 B.n184 585
R249 B.n183 B.n182 585
R250 B.n181 B.n180 585
R251 B.n179 B.n178 585
R252 B.n177 B.n176 585
R253 B.n175 B.n174 585
R254 B.n173 B.n172 585
R255 B.n171 B.n170 585
R256 B.n169 B.n168 585
R257 B.n167 B.n166 585
R258 B.n165 B.n164 585
R259 B.n163 B.n162 585
R260 B.n161 B.n160 585
R261 B.n159 B.n158 585
R262 B.n157 B.n156 585
R263 B.n117 B.n116 585
R264 B.n862 B.n861 585
R265 B.n855 B.n151 585
R266 B.n151 B.n114 585
R267 B.n854 B.n113 585
R268 B.n866 B.n113 585
R269 B.n853 B.n112 585
R270 B.n867 B.n112 585
R271 B.n852 B.n111 585
R272 B.n868 B.n111 585
R273 B.n851 B.n850 585
R274 B.n850 B.n107 585
R275 B.n849 B.n106 585
R276 B.n874 B.n106 585
R277 B.n848 B.n105 585
R278 B.n875 B.n105 585
R279 B.n847 B.n104 585
R280 B.n876 B.n104 585
R281 B.n846 B.n845 585
R282 B.n845 B.n100 585
R283 B.n844 B.n99 585
R284 B.n882 B.n99 585
R285 B.n843 B.n98 585
R286 B.n883 B.n98 585
R287 B.n842 B.n97 585
R288 B.n884 B.n97 585
R289 B.n841 B.n840 585
R290 B.n840 B.n93 585
R291 B.n839 B.n92 585
R292 B.n890 B.n92 585
R293 B.n838 B.n91 585
R294 B.n891 B.n91 585
R295 B.n837 B.n90 585
R296 B.n892 B.n90 585
R297 B.n836 B.n835 585
R298 B.n835 B.n86 585
R299 B.n834 B.n85 585
R300 B.n898 B.n85 585
R301 B.n833 B.n84 585
R302 B.n899 B.n84 585
R303 B.n832 B.n83 585
R304 B.n900 B.n83 585
R305 B.n831 B.n830 585
R306 B.n830 B.n82 585
R307 B.n829 B.n78 585
R308 B.n906 B.n78 585
R309 B.n828 B.n77 585
R310 B.n907 B.n77 585
R311 B.n827 B.n76 585
R312 B.n908 B.n76 585
R313 B.n826 B.n825 585
R314 B.n825 B.n72 585
R315 B.n824 B.n71 585
R316 B.n914 B.n71 585
R317 B.n823 B.n70 585
R318 B.n915 B.n70 585
R319 B.n822 B.n69 585
R320 B.n916 B.n69 585
R321 B.n821 B.n820 585
R322 B.n820 B.n65 585
R323 B.n819 B.n64 585
R324 B.n922 B.n64 585
R325 B.n818 B.n63 585
R326 B.n923 B.n63 585
R327 B.n817 B.n62 585
R328 B.n924 B.n62 585
R329 B.n816 B.n815 585
R330 B.n815 B.n58 585
R331 B.n814 B.n57 585
R332 B.n930 B.n57 585
R333 B.n813 B.n56 585
R334 B.n931 B.n56 585
R335 B.n812 B.n55 585
R336 B.n932 B.n55 585
R337 B.n811 B.n810 585
R338 B.n810 B.n51 585
R339 B.n809 B.n50 585
R340 B.n938 B.n50 585
R341 B.n808 B.n49 585
R342 B.n939 B.n49 585
R343 B.n807 B.n48 585
R344 B.n940 B.n48 585
R345 B.n806 B.n805 585
R346 B.n805 B.n44 585
R347 B.n804 B.n43 585
R348 B.n946 B.n43 585
R349 B.n803 B.n42 585
R350 B.n947 B.n42 585
R351 B.n802 B.n41 585
R352 B.n948 B.n41 585
R353 B.n801 B.n800 585
R354 B.n800 B.n37 585
R355 B.n799 B.n36 585
R356 B.n954 B.n36 585
R357 B.n798 B.n35 585
R358 B.n955 B.n35 585
R359 B.n797 B.n34 585
R360 B.n956 B.n34 585
R361 B.n796 B.n795 585
R362 B.n795 B.n33 585
R363 B.n794 B.n29 585
R364 B.n962 B.n29 585
R365 B.n793 B.n28 585
R366 B.n963 B.n28 585
R367 B.n792 B.n27 585
R368 B.n964 B.n27 585
R369 B.n791 B.n790 585
R370 B.n790 B.n23 585
R371 B.n789 B.n22 585
R372 B.n970 B.n22 585
R373 B.n788 B.n21 585
R374 B.n971 B.n21 585
R375 B.n787 B.n20 585
R376 B.n972 B.n20 585
R377 B.n786 B.n785 585
R378 B.n785 B.n16 585
R379 B.n784 B.n15 585
R380 B.n978 B.n15 585
R381 B.n783 B.n14 585
R382 B.n979 B.n14 585
R383 B.n782 B.n13 585
R384 B.n980 B.n13 585
R385 B.n781 B.n780 585
R386 B.n780 B.n12 585
R387 B.n779 B.n778 585
R388 B.n779 B.n8 585
R389 B.n777 B.n7 585
R390 B.n987 B.n7 585
R391 B.n776 B.n6 585
R392 B.n988 B.n6 585
R393 B.n775 B.n5 585
R394 B.n989 B.n5 585
R395 B.n774 B.n773 585
R396 B.n773 B.n4 585
R397 B.n772 B.n287 585
R398 B.n772 B.n771 585
R399 B.n762 B.n288 585
R400 B.n289 B.n288 585
R401 B.n764 B.n763 585
R402 B.n765 B.n764 585
R403 B.n761 B.n294 585
R404 B.n294 B.n293 585
R405 B.n760 B.n759 585
R406 B.n759 B.n758 585
R407 B.n296 B.n295 585
R408 B.n297 B.n296 585
R409 B.n751 B.n750 585
R410 B.n752 B.n751 585
R411 B.n749 B.n302 585
R412 B.n302 B.n301 585
R413 B.n748 B.n747 585
R414 B.n747 B.n746 585
R415 B.n304 B.n303 585
R416 B.n305 B.n304 585
R417 B.n739 B.n738 585
R418 B.n740 B.n739 585
R419 B.n737 B.n310 585
R420 B.n310 B.n309 585
R421 B.n736 B.n735 585
R422 B.n735 B.n734 585
R423 B.n312 B.n311 585
R424 B.n727 B.n312 585
R425 B.n726 B.n725 585
R426 B.n728 B.n726 585
R427 B.n724 B.n317 585
R428 B.n317 B.n316 585
R429 B.n723 B.n722 585
R430 B.n722 B.n721 585
R431 B.n319 B.n318 585
R432 B.n320 B.n319 585
R433 B.n714 B.n713 585
R434 B.n715 B.n714 585
R435 B.n712 B.n325 585
R436 B.n325 B.n324 585
R437 B.n711 B.n710 585
R438 B.n710 B.n709 585
R439 B.n327 B.n326 585
R440 B.n328 B.n327 585
R441 B.n702 B.n701 585
R442 B.n703 B.n702 585
R443 B.n700 B.n332 585
R444 B.n336 B.n332 585
R445 B.n699 B.n698 585
R446 B.n698 B.n697 585
R447 B.n334 B.n333 585
R448 B.n335 B.n334 585
R449 B.n690 B.n689 585
R450 B.n691 B.n690 585
R451 B.n688 B.n341 585
R452 B.n341 B.n340 585
R453 B.n687 B.n686 585
R454 B.n686 B.n685 585
R455 B.n343 B.n342 585
R456 B.n344 B.n343 585
R457 B.n678 B.n677 585
R458 B.n679 B.n678 585
R459 B.n676 B.n349 585
R460 B.n349 B.n348 585
R461 B.n675 B.n674 585
R462 B.n674 B.n673 585
R463 B.n351 B.n350 585
R464 B.n352 B.n351 585
R465 B.n666 B.n665 585
R466 B.n667 B.n666 585
R467 B.n664 B.n357 585
R468 B.n357 B.n356 585
R469 B.n663 B.n662 585
R470 B.n662 B.n661 585
R471 B.n359 B.n358 585
R472 B.n360 B.n359 585
R473 B.n654 B.n653 585
R474 B.n655 B.n654 585
R475 B.n652 B.n365 585
R476 B.n365 B.n364 585
R477 B.n651 B.n650 585
R478 B.n650 B.n649 585
R479 B.n367 B.n366 585
R480 B.n642 B.n367 585
R481 B.n641 B.n640 585
R482 B.n643 B.n641 585
R483 B.n639 B.n372 585
R484 B.n372 B.n371 585
R485 B.n638 B.n637 585
R486 B.n637 B.n636 585
R487 B.n374 B.n373 585
R488 B.n375 B.n374 585
R489 B.n629 B.n628 585
R490 B.n630 B.n629 585
R491 B.n627 B.n380 585
R492 B.n380 B.n379 585
R493 B.n626 B.n625 585
R494 B.n625 B.n624 585
R495 B.n382 B.n381 585
R496 B.n383 B.n382 585
R497 B.n617 B.n616 585
R498 B.n618 B.n617 585
R499 B.n615 B.n388 585
R500 B.n388 B.n387 585
R501 B.n614 B.n613 585
R502 B.n613 B.n612 585
R503 B.n390 B.n389 585
R504 B.n391 B.n390 585
R505 B.n605 B.n604 585
R506 B.n606 B.n605 585
R507 B.n603 B.n396 585
R508 B.n396 B.n395 585
R509 B.n602 B.n601 585
R510 B.n601 B.n600 585
R511 B.n398 B.n397 585
R512 B.n399 B.n398 585
R513 B.n593 B.n592 585
R514 B.n594 B.n593 585
R515 B.n591 B.n404 585
R516 B.n404 B.n403 585
R517 B.n590 B.n589 585
R518 B.n589 B.n588 585
R519 B.n406 B.n405 585
R520 B.n407 B.n406 585
R521 B.n584 B.n583 585
R522 B.n410 B.n409 585
R523 B.n580 B.n579 585
R524 B.n581 B.n580 585
R525 B.n578 B.n444 585
R526 B.n577 B.n576 585
R527 B.n575 B.n574 585
R528 B.n573 B.n572 585
R529 B.n571 B.n570 585
R530 B.n569 B.n568 585
R531 B.n567 B.n566 585
R532 B.n565 B.n564 585
R533 B.n563 B.n562 585
R534 B.n561 B.n560 585
R535 B.n559 B.n558 585
R536 B.n557 B.n556 585
R537 B.n555 B.n554 585
R538 B.n553 B.n552 585
R539 B.n551 B.n550 585
R540 B.n549 B.n548 585
R541 B.n547 B.n546 585
R542 B.n545 B.n544 585
R543 B.n543 B.n542 585
R544 B.n541 B.n540 585
R545 B.n539 B.n538 585
R546 B.n537 B.n536 585
R547 B.n535 B.n534 585
R548 B.n533 B.n532 585
R549 B.n531 B.n530 585
R550 B.n529 B.n528 585
R551 B.n527 B.n526 585
R552 B.n525 B.n524 585
R553 B.n523 B.n522 585
R554 B.n521 B.n520 585
R555 B.n519 B.n518 585
R556 B.n517 B.n516 585
R557 B.n515 B.n514 585
R558 B.n513 B.n512 585
R559 B.n511 B.n510 585
R560 B.n509 B.n508 585
R561 B.n507 B.n506 585
R562 B.n505 B.n504 585
R563 B.n503 B.n502 585
R564 B.n501 B.n500 585
R565 B.n499 B.n498 585
R566 B.n497 B.n496 585
R567 B.n495 B.n494 585
R568 B.n493 B.n492 585
R569 B.n491 B.n490 585
R570 B.n489 B.n488 585
R571 B.n487 B.n486 585
R572 B.n485 B.n484 585
R573 B.n483 B.n482 585
R574 B.n481 B.n480 585
R575 B.n479 B.n478 585
R576 B.n477 B.n476 585
R577 B.n475 B.n474 585
R578 B.n473 B.n472 585
R579 B.n471 B.n470 585
R580 B.n469 B.n468 585
R581 B.n467 B.n466 585
R582 B.n465 B.n464 585
R583 B.n463 B.n462 585
R584 B.n461 B.n460 585
R585 B.n459 B.n458 585
R586 B.n457 B.n456 585
R587 B.n455 B.n454 585
R588 B.n453 B.n452 585
R589 B.n451 B.n443 585
R590 B.n581 B.n443 585
R591 B.n585 B.n408 585
R592 B.n408 B.n407 585
R593 B.n587 B.n586 585
R594 B.n588 B.n587 585
R595 B.n402 B.n401 585
R596 B.n403 B.n402 585
R597 B.n596 B.n595 585
R598 B.n595 B.n594 585
R599 B.n597 B.n400 585
R600 B.n400 B.n399 585
R601 B.n599 B.n598 585
R602 B.n600 B.n599 585
R603 B.n394 B.n393 585
R604 B.n395 B.n394 585
R605 B.n608 B.n607 585
R606 B.n607 B.n606 585
R607 B.n609 B.n392 585
R608 B.n392 B.n391 585
R609 B.n611 B.n610 585
R610 B.n612 B.n611 585
R611 B.n386 B.n385 585
R612 B.n387 B.n386 585
R613 B.n620 B.n619 585
R614 B.n619 B.n618 585
R615 B.n621 B.n384 585
R616 B.n384 B.n383 585
R617 B.n623 B.n622 585
R618 B.n624 B.n623 585
R619 B.n378 B.n377 585
R620 B.n379 B.n378 585
R621 B.n632 B.n631 585
R622 B.n631 B.n630 585
R623 B.n633 B.n376 585
R624 B.n376 B.n375 585
R625 B.n635 B.n634 585
R626 B.n636 B.n635 585
R627 B.n370 B.n369 585
R628 B.n371 B.n370 585
R629 B.n645 B.n644 585
R630 B.n644 B.n643 585
R631 B.n646 B.n368 585
R632 B.n642 B.n368 585
R633 B.n648 B.n647 585
R634 B.n649 B.n648 585
R635 B.n363 B.n362 585
R636 B.n364 B.n363 585
R637 B.n657 B.n656 585
R638 B.n656 B.n655 585
R639 B.n658 B.n361 585
R640 B.n361 B.n360 585
R641 B.n660 B.n659 585
R642 B.n661 B.n660 585
R643 B.n355 B.n354 585
R644 B.n356 B.n355 585
R645 B.n669 B.n668 585
R646 B.n668 B.n667 585
R647 B.n670 B.n353 585
R648 B.n353 B.n352 585
R649 B.n672 B.n671 585
R650 B.n673 B.n672 585
R651 B.n347 B.n346 585
R652 B.n348 B.n347 585
R653 B.n681 B.n680 585
R654 B.n680 B.n679 585
R655 B.n682 B.n345 585
R656 B.n345 B.n344 585
R657 B.n684 B.n683 585
R658 B.n685 B.n684 585
R659 B.n339 B.n338 585
R660 B.n340 B.n339 585
R661 B.n693 B.n692 585
R662 B.n692 B.n691 585
R663 B.n694 B.n337 585
R664 B.n337 B.n335 585
R665 B.n696 B.n695 585
R666 B.n697 B.n696 585
R667 B.n331 B.n330 585
R668 B.n336 B.n331 585
R669 B.n705 B.n704 585
R670 B.n704 B.n703 585
R671 B.n706 B.n329 585
R672 B.n329 B.n328 585
R673 B.n708 B.n707 585
R674 B.n709 B.n708 585
R675 B.n323 B.n322 585
R676 B.n324 B.n323 585
R677 B.n717 B.n716 585
R678 B.n716 B.n715 585
R679 B.n718 B.n321 585
R680 B.n321 B.n320 585
R681 B.n720 B.n719 585
R682 B.n721 B.n720 585
R683 B.n315 B.n314 585
R684 B.n316 B.n315 585
R685 B.n730 B.n729 585
R686 B.n729 B.n728 585
R687 B.n731 B.n313 585
R688 B.n727 B.n313 585
R689 B.n733 B.n732 585
R690 B.n734 B.n733 585
R691 B.n308 B.n307 585
R692 B.n309 B.n308 585
R693 B.n742 B.n741 585
R694 B.n741 B.n740 585
R695 B.n743 B.n306 585
R696 B.n306 B.n305 585
R697 B.n745 B.n744 585
R698 B.n746 B.n745 585
R699 B.n300 B.n299 585
R700 B.n301 B.n300 585
R701 B.n754 B.n753 585
R702 B.n753 B.n752 585
R703 B.n755 B.n298 585
R704 B.n298 B.n297 585
R705 B.n757 B.n756 585
R706 B.n758 B.n757 585
R707 B.n292 B.n291 585
R708 B.n293 B.n292 585
R709 B.n767 B.n766 585
R710 B.n766 B.n765 585
R711 B.n768 B.n290 585
R712 B.n290 B.n289 585
R713 B.n770 B.n769 585
R714 B.n771 B.n770 585
R715 B.n3 B.n0 585
R716 B.n4 B.n3 585
R717 B.n986 B.n1 585
R718 B.n987 B.n986 585
R719 B.n985 B.n984 585
R720 B.n985 B.n8 585
R721 B.n983 B.n9 585
R722 B.n12 B.n9 585
R723 B.n982 B.n981 585
R724 B.n981 B.n980 585
R725 B.n11 B.n10 585
R726 B.n979 B.n11 585
R727 B.n977 B.n976 585
R728 B.n978 B.n977 585
R729 B.n975 B.n17 585
R730 B.n17 B.n16 585
R731 B.n974 B.n973 585
R732 B.n973 B.n972 585
R733 B.n19 B.n18 585
R734 B.n971 B.n19 585
R735 B.n969 B.n968 585
R736 B.n970 B.n969 585
R737 B.n967 B.n24 585
R738 B.n24 B.n23 585
R739 B.n966 B.n965 585
R740 B.n965 B.n964 585
R741 B.n26 B.n25 585
R742 B.n963 B.n26 585
R743 B.n961 B.n960 585
R744 B.n962 B.n961 585
R745 B.n959 B.n30 585
R746 B.n33 B.n30 585
R747 B.n958 B.n957 585
R748 B.n957 B.n956 585
R749 B.n32 B.n31 585
R750 B.n955 B.n32 585
R751 B.n953 B.n952 585
R752 B.n954 B.n953 585
R753 B.n951 B.n38 585
R754 B.n38 B.n37 585
R755 B.n950 B.n949 585
R756 B.n949 B.n948 585
R757 B.n40 B.n39 585
R758 B.n947 B.n40 585
R759 B.n945 B.n944 585
R760 B.n946 B.n945 585
R761 B.n943 B.n45 585
R762 B.n45 B.n44 585
R763 B.n942 B.n941 585
R764 B.n941 B.n940 585
R765 B.n47 B.n46 585
R766 B.n939 B.n47 585
R767 B.n937 B.n936 585
R768 B.n938 B.n937 585
R769 B.n935 B.n52 585
R770 B.n52 B.n51 585
R771 B.n934 B.n933 585
R772 B.n933 B.n932 585
R773 B.n54 B.n53 585
R774 B.n931 B.n54 585
R775 B.n929 B.n928 585
R776 B.n930 B.n929 585
R777 B.n927 B.n59 585
R778 B.n59 B.n58 585
R779 B.n926 B.n925 585
R780 B.n925 B.n924 585
R781 B.n61 B.n60 585
R782 B.n923 B.n61 585
R783 B.n921 B.n920 585
R784 B.n922 B.n921 585
R785 B.n919 B.n66 585
R786 B.n66 B.n65 585
R787 B.n918 B.n917 585
R788 B.n917 B.n916 585
R789 B.n68 B.n67 585
R790 B.n915 B.n68 585
R791 B.n913 B.n912 585
R792 B.n914 B.n913 585
R793 B.n911 B.n73 585
R794 B.n73 B.n72 585
R795 B.n910 B.n909 585
R796 B.n909 B.n908 585
R797 B.n75 B.n74 585
R798 B.n907 B.n75 585
R799 B.n905 B.n904 585
R800 B.n906 B.n905 585
R801 B.n903 B.n79 585
R802 B.n82 B.n79 585
R803 B.n902 B.n901 585
R804 B.n901 B.n900 585
R805 B.n81 B.n80 585
R806 B.n899 B.n81 585
R807 B.n897 B.n896 585
R808 B.n898 B.n897 585
R809 B.n895 B.n87 585
R810 B.n87 B.n86 585
R811 B.n894 B.n893 585
R812 B.n893 B.n892 585
R813 B.n89 B.n88 585
R814 B.n891 B.n89 585
R815 B.n889 B.n888 585
R816 B.n890 B.n889 585
R817 B.n887 B.n94 585
R818 B.n94 B.n93 585
R819 B.n886 B.n885 585
R820 B.n885 B.n884 585
R821 B.n96 B.n95 585
R822 B.n883 B.n96 585
R823 B.n881 B.n880 585
R824 B.n882 B.n881 585
R825 B.n879 B.n101 585
R826 B.n101 B.n100 585
R827 B.n878 B.n877 585
R828 B.n877 B.n876 585
R829 B.n103 B.n102 585
R830 B.n875 B.n103 585
R831 B.n873 B.n872 585
R832 B.n874 B.n873 585
R833 B.n871 B.n108 585
R834 B.n108 B.n107 585
R835 B.n870 B.n869 585
R836 B.n869 B.n868 585
R837 B.n110 B.n109 585
R838 B.n867 B.n110 585
R839 B.n865 B.n864 585
R840 B.n866 B.n865 585
R841 B.n863 B.n115 585
R842 B.n115 B.n114 585
R843 B.n990 B.n989 585
R844 B.n988 B.n2 585
R845 B.n861 B.n115 516.524
R846 B.n857 B.n151 516.524
R847 B.n443 B.n406 516.524
R848 B.n583 B.n408 516.524
R849 B.n154 B.t14 275.327
R850 B.n152 B.t21 275.327
R851 B.n448 B.t18 275.327
R852 B.n445 B.t10 275.327
R853 B.n859 B.n858 256.663
R854 B.n859 B.n149 256.663
R855 B.n859 B.n148 256.663
R856 B.n859 B.n147 256.663
R857 B.n859 B.n146 256.663
R858 B.n859 B.n145 256.663
R859 B.n859 B.n144 256.663
R860 B.n859 B.n143 256.663
R861 B.n859 B.n142 256.663
R862 B.n859 B.n141 256.663
R863 B.n859 B.n140 256.663
R864 B.n859 B.n139 256.663
R865 B.n859 B.n138 256.663
R866 B.n859 B.n137 256.663
R867 B.n859 B.n136 256.663
R868 B.n859 B.n135 256.663
R869 B.n859 B.n134 256.663
R870 B.n859 B.n133 256.663
R871 B.n859 B.n132 256.663
R872 B.n859 B.n131 256.663
R873 B.n859 B.n130 256.663
R874 B.n859 B.n129 256.663
R875 B.n859 B.n128 256.663
R876 B.n859 B.n127 256.663
R877 B.n859 B.n126 256.663
R878 B.n859 B.n125 256.663
R879 B.n859 B.n124 256.663
R880 B.n859 B.n123 256.663
R881 B.n859 B.n122 256.663
R882 B.n859 B.n121 256.663
R883 B.n859 B.n120 256.663
R884 B.n859 B.n119 256.663
R885 B.n859 B.n118 256.663
R886 B.n860 B.n859 256.663
R887 B.n582 B.n581 256.663
R888 B.n581 B.n411 256.663
R889 B.n581 B.n412 256.663
R890 B.n581 B.n413 256.663
R891 B.n581 B.n414 256.663
R892 B.n581 B.n415 256.663
R893 B.n581 B.n416 256.663
R894 B.n581 B.n417 256.663
R895 B.n581 B.n418 256.663
R896 B.n581 B.n419 256.663
R897 B.n581 B.n420 256.663
R898 B.n581 B.n421 256.663
R899 B.n581 B.n422 256.663
R900 B.n581 B.n423 256.663
R901 B.n581 B.n424 256.663
R902 B.n581 B.n425 256.663
R903 B.n581 B.n426 256.663
R904 B.n581 B.n427 256.663
R905 B.n581 B.n428 256.663
R906 B.n581 B.n429 256.663
R907 B.n581 B.n430 256.663
R908 B.n581 B.n431 256.663
R909 B.n581 B.n432 256.663
R910 B.n581 B.n433 256.663
R911 B.n581 B.n434 256.663
R912 B.n581 B.n435 256.663
R913 B.n581 B.n436 256.663
R914 B.n581 B.n437 256.663
R915 B.n581 B.n438 256.663
R916 B.n581 B.n439 256.663
R917 B.n581 B.n440 256.663
R918 B.n581 B.n441 256.663
R919 B.n581 B.n442 256.663
R920 B.n992 B.n991 256.663
R921 B.n156 B.n117 163.367
R922 B.n160 B.n159 163.367
R923 B.n164 B.n163 163.367
R924 B.n168 B.n167 163.367
R925 B.n172 B.n171 163.367
R926 B.n176 B.n175 163.367
R927 B.n180 B.n179 163.367
R928 B.n184 B.n183 163.367
R929 B.n188 B.n187 163.367
R930 B.n192 B.n191 163.367
R931 B.n196 B.n195 163.367
R932 B.n200 B.n199 163.367
R933 B.n204 B.n203 163.367
R934 B.n208 B.n207 163.367
R935 B.n213 B.n212 163.367
R936 B.n217 B.n216 163.367
R937 B.n221 B.n220 163.367
R938 B.n225 B.n224 163.367
R939 B.n229 B.n228 163.367
R940 B.n234 B.n233 163.367
R941 B.n238 B.n237 163.367
R942 B.n242 B.n241 163.367
R943 B.n246 B.n245 163.367
R944 B.n250 B.n249 163.367
R945 B.n254 B.n253 163.367
R946 B.n258 B.n257 163.367
R947 B.n262 B.n261 163.367
R948 B.n266 B.n265 163.367
R949 B.n270 B.n269 163.367
R950 B.n274 B.n273 163.367
R951 B.n278 B.n277 163.367
R952 B.n282 B.n281 163.367
R953 B.n284 B.n150 163.367
R954 B.n589 B.n406 163.367
R955 B.n589 B.n404 163.367
R956 B.n593 B.n404 163.367
R957 B.n593 B.n398 163.367
R958 B.n601 B.n398 163.367
R959 B.n601 B.n396 163.367
R960 B.n605 B.n396 163.367
R961 B.n605 B.n390 163.367
R962 B.n613 B.n390 163.367
R963 B.n613 B.n388 163.367
R964 B.n617 B.n388 163.367
R965 B.n617 B.n382 163.367
R966 B.n625 B.n382 163.367
R967 B.n625 B.n380 163.367
R968 B.n629 B.n380 163.367
R969 B.n629 B.n374 163.367
R970 B.n637 B.n374 163.367
R971 B.n637 B.n372 163.367
R972 B.n641 B.n372 163.367
R973 B.n641 B.n367 163.367
R974 B.n650 B.n367 163.367
R975 B.n650 B.n365 163.367
R976 B.n654 B.n365 163.367
R977 B.n654 B.n359 163.367
R978 B.n662 B.n359 163.367
R979 B.n662 B.n357 163.367
R980 B.n666 B.n357 163.367
R981 B.n666 B.n351 163.367
R982 B.n674 B.n351 163.367
R983 B.n674 B.n349 163.367
R984 B.n678 B.n349 163.367
R985 B.n678 B.n343 163.367
R986 B.n686 B.n343 163.367
R987 B.n686 B.n341 163.367
R988 B.n690 B.n341 163.367
R989 B.n690 B.n334 163.367
R990 B.n698 B.n334 163.367
R991 B.n698 B.n332 163.367
R992 B.n702 B.n332 163.367
R993 B.n702 B.n327 163.367
R994 B.n710 B.n327 163.367
R995 B.n710 B.n325 163.367
R996 B.n714 B.n325 163.367
R997 B.n714 B.n319 163.367
R998 B.n722 B.n319 163.367
R999 B.n722 B.n317 163.367
R1000 B.n726 B.n317 163.367
R1001 B.n726 B.n312 163.367
R1002 B.n735 B.n312 163.367
R1003 B.n735 B.n310 163.367
R1004 B.n739 B.n310 163.367
R1005 B.n739 B.n304 163.367
R1006 B.n747 B.n304 163.367
R1007 B.n747 B.n302 163.367
R1008 B.n751 B.n302 163.367
R1009 B.n751 B.n296 163.367
R1010 B.n759 B.n296 163.367
R1011 B.n759 B.n294 163.367
R1012 B.n764 B.n294 163.367
R1013 B.n764 B.n288 163.367
R1014 B.n772 B.n288 163.367
R1015 B.n773 B.n772 163.367
R1016 B.n773 B.n5 163.367
R1017 B.n6 B.n5 163.367
R1018 B.n7 B.n6 163.367
R1019 B.n779 B.n7 163.367
R1020 B.n780 B.n779 163.367
R1021 B.n780 B.n13 163.367
R1022 B.n14 B.n13 163.367
R1023 B.n15 B.n14 163.367
R1024 B.n785 B.n15 163.367
R1025 B.n785 B.n20 163.367
R1026 B.n21 B.n20 163.367
R1027 B.n22 B.n21 163.367
R1028 B.n790 B.n22 163.367
R1029 B.n790 B.n27 163.367
R1030 B.n28 B.n27 163.367
R1031 B.n29 B.n28 163.367
R1032 B.n795 B.n29 163.367
R1033 B.n795 B.n34 163.367
R1034 B.n35 B.n34 163.367
R1035 B.n36 B.n35 163.367
R1036 B.n800 B.n36 163.367
R1037 B.n800 B.n41 163.367
R1038 B.n42 B.n41 163.367
R1039 B.n43 B.n42 163.367
R1040 B.n805 B.n43 163.367
R1041 B.n805 B.n48 163.367
R1042 B.n49 B.n48 163.367
R1043 B.n50 B.n49 163.367
R1044 B.n810 B.n50 163.367
R1045 B.n810 B.n55 163.367
R1046 B.n56 B.n55 163.367
R1047 B.n57 B.n56 163.367
R1048 B.n815 B.n57 163.367
R1049 B.n815 B.n62 163.367
R1050 B.n63 B.n62 163.367
R1051 B.n64 B.n63 163.367
R1052 B.n820 B.n64 163.367
R1053 B.n820 B.n69 163.367
R1054 B.n70 B.n69 163.367
R1055 B.n71 B.n70 163.367
R1056 B.n825 B.n71 163.367
R1057 B.n825 B.n76 163.367
R1058 B.n77 B.n76 163.367
R1059 B.n78 B.n77 163.367
R1060 B.n830 B.n78 163.367
R1061 B.n830 B.n83 163.367
R1062 B.n84 B.n83 163.367
R1063 B.n85 B.n84 163.367
R1064 B.n835 B.n85 163.367
R1065 B.n835 B.n90 163.367
R1066 B.n91 B.n90 163.367
R1067 B.n92 B.n91 163.367
R1068 B.n840 B.n92 163.367
R1069 B.n840 B.n97 163.367
R1070 B.n98 B.n97 163.367
R1071 B.n99 B.n98 163.367
R1072 B.n845 B.n99 163.367
R1073 B.n845 B.n104 163.367
R1074 B.n105 B.n104 163.367
R1075 B.n106 B.n105 163.367
R1076 B.n850 B.n106 163.367
R1077 B.n850 B.n111 163.367
R1078 B.n112 B.n111 163.367
R1079 B.n113 B.n112 163.367
R1080 B.n151 B.n113 163.367
R1081 B.n580 B.n410 163.367
R1082 B.n580 B.n444 163.367
R1083 B.n576 B.n575 163.367
R1084 B.n572 B.n571 163.367
R1085 B.n568 B.n567 163.367
R1086 B.n564 B.n563 163.367
R1087 B.n560 B.n559 163.367
R1088 B.n556 B.n555 163.367
R1089 B.n552 B.n551 163.367
R1090 B.n548 B.n547 163.367
R1091 B.n544 B.n543 163.367
R1092 B.n540 B.n539 163.367
R1093 B.n536 B.n535 163.367
R1094 B.n532 B.n531 163.367
R1095 B.n528 B.n527 163.367
R1096 B.n524 B.n523 163.367
R1097 B.n520 B.n519 163.367
R1098 B.n516 B.n515 163.367
R1099 B.n512 B.n511 163.367
R1100 B.n508 B.n507 163.367
R1101 B.n504 B.n503 163.367
R1102 B.n500 B.n499 163.367
R1103 B.n496 B.n495 163.367
R1104 B.n492 B.n491 163.367
R1105 B.n488 B.n487 163.367
R1106 B.n484 B.n483 163.367
R1107 B.n480 B.n479 163.367
R1108 B.n476 B.n475 163.367
R1109 B.n472 B.n471 163.367
R1110 B.n468 B.n467 163.367
R1111 B.n464 B.n463 163.367
R1112 B.n460 B.n459 163.367
R1113 B.n456 B.n455 163.367
R1114 B.n452 B.n443 163.367
R1115 B.n587 B.n408 163.367
R1116 B.n587 B.n402 163.367
R1117 B.n595 B.n402 163.367
R1118 B.n595 B.n400 163.367
R1119 B.n599 B.n400 163.367
R1120 B.n599 B.n394 163.367
R1121 B.n607 B.n394 163.367
R1122 B.n607 B.n392 163.367
R1123 B.n611 B.n392 163.367
R1124 B.n611 B.n386 163.367
R1125 B.n619 B.n386 163.367
R1126 B.n619 B.n384 163.367
R1127 B.n623 B.n384 163.367
R1128 B.n623 B.n378 163.367
R1129 B.n631 B.n378 163.367
R1130 B.n631 B.n376 163.367
R1131 B.n635 B.n376 163.367
R1132 B.n635 B.n370 163.367
R1133 B.n644 B.n370 163.367
R1134 B.n644 B.n368 163.367
R1135 B.n648 B.n368 163.367
R1136 B.n648 B.n363 163.367
R1137 B.n656 B.n363 163.367
R1138 B.n656 B.n361 163.367
R1139 B.n660 B.n361 163.367
R1140 B.n660 B.n355 163.367
R1141 B.n668 B.n355 163.367
R1142 B.n668 B.n353 163.367
R1143 B.n672 B.n353 163.367
R1144 B.n672 B.n347 163.367
R1145 B.n680 B.n347 163.367
R1146 B.n680 B.n345 163.367
R1147 B.n684 B.n345 163.367
R1148 B.n684 B.n339 163.367
R1149 B.n692 B.n339 163.367
R1150 B.n692 B.n337 163.367
R1151 B.n696 B.n337 163.367
R1152 B.n696 B.n331 163.367
R1153 B.n704 B.n331 163.367
R1154 B.n704 B.n329 163.367
R1155 B.n708 B.n329 163.367
R1156 B.n708 B.n323 163.367
R1157 B.n716 B.n323 163.367
R1158 B.n716 B.n321 163.367
R1159 B.n720 B.n321 163.367
R1160 B.n720 B.n315 163.367
R1161 B.n729 B.n315 163.367
R1162 B.n729 B.n313 163.367
R1163 B.n733 B.n313 163.367
R1164 B.n733 B.n308 163.367
R1165 B.n741 B.n308 163.367
R1166 B.n741 B.n306 163.367
R1167 B.n745 B.n306 163.367
R1168 B.n745 B.n300 163.367
R1169 B.n753 B.n300 163.367
R1170 B.n753 B.n298 163.367
R1171 B.n757 B.n298 163.367
R1172 B.n757 B.n292 163.367
R1173 B.n766 B.n292 163.367
R1174 B.n766 B.n290 163.367
R1175 B.n770 B.n290 163.367
R1176 B.n770 B.n3 163.367
R1177 B.n990 B.n3 163.367
R1178 B.n986 B.n2 163.367
R1179 B.n986 B.n985 163.367
R1180 B.n985 B.n9 163.367
R1181 B.n981 B.n9 163.367
R1182 B.n981 B.n11 163.367
R1183 B.n977 B.n11 163.367
R1184 B.n977 B.n17 163.367
R1185 B.n973 B.n17 163.367
R1186 B.n973 B.n19 163.367
R1187 B.n969 B.n19 163.367
R1188 B.n969 B.n24 163.367
R1189 B.n965 B.n24 163.367
R1190 B.n965 B.n26 163.367
R1191 B.n961 B.n26 163.367
R1192 B.n961 B.n30 163.367
R1193 B.n957 B.n30 163.367
R1194 B.n957 B.n32 163.367
R1195 B.n953 B.n32 163.367
R1196 B.n953 B.n38 163.367
R1197 B.n949 B.n38 163.367
R1198 B.n949 B.n40 163.367
R1199 B.n945 B.n40 163.367
R1200 B.n945 B.n45 163.367
R1201 B.n941 B.n45 163.367
R1202 B.n941 B.n47 163.367
R1203 B.n937 B.n47 163.367
R1204 B.n937 B.n52 163.367
R1205 B.n933 B.n52 163.367
R1206 B.n933 B.n54 163.367
R1207 B.n929 B.n54 163.367
R1208 B.n929 B.n59 163.367
R1209 B.n925 B.n59 163.367
R1210 B.n925 B.n61 163.367
R1211 B.n921 B.n61 163.367
R1212 B.n921 B.n66 163.367
R1213 B.n917 B.n66 163.367
R1214 B.n917 B.n68 163.367
R1215 B.n913 B.n68 163.367
R1216 B.n913 B.n73 163.367
R1217 B.n909 B.n73 163.367
R1218 B.n909 B.n75 163.367
R1219 B.n905 B.n75 163.367
R1220 B.n905 B.n79 163.367
R1221 B.n901 B.n79 163.367
R1222 B.n901 B.n81 163.367
R1223 B.n897 B.n81 163.367
R1224 B.n897 B.n87 163.367
R1225 B.n893 B.n87 163.367
R1226 B.n893 B.n89 163.367
R1227 B.n889 B.n89 163.367
R1228 B.n889 B.n94 163.367
R1229 B.n885 B.n94 163.367
R1230 B.n885 B.n96 163.367
R1231 B.n881 B.n96 163.367
R1232 B.n881 B.n101 163.367
R1233 B.n877 B.n101 163.367
R1234 B.n877 B.n103 163.367
R1235 B.n873 B.n103 163.367
R1236 B.n873 B.n108 163.367
R1237 B.n869 B.n108 163.367
R1238 B.n869 B.n110 163.367
R1239 B.n865 B.n110 163.367
R1240 B.n865 B.n115 163.367
R1241 B.n152 B.t22 135.968
R1242 B.n448 B.t20 135.968
R1243 B.n154 B.t16 135.958
R1244 B.n445 B.t13 135.958
R1245 B.n581 B.n407 105.082
R1246 B.n859 B.n114 105.082
R1247 B.n153 B.t23 75.07
R1248 B.n449 B.t19 75.07
R1249 B.n155 B.t17 75.0613
R1250 B.n446 B.t12 75.0613
R1251 B.n861 B.n860 71.676
R1252 B.n156 B.n118 71.676
R1253 B.n160 B.n119 71.676
R1254 B.n164 B.n120 71.676
R1255 B.n168 B.n121 71.676
R1256 B.n172 B.n122 71.676
R1257 B.n176 B.n123 71.676
R1258 B.n180 B.n124 71.676
R1259 B.n184 B.n125 71.676
R1260 B.n188 B.n126 71.676
R1261 B.n192 B.n127 71.676
R1262 B.n196 B.n128 71.676
R1263 B.n200 B.n129 71.676
R1264 B.n204 B.n130 71.676
R1265 B.n208 B.n131 71.676
R1266 B.n213 B.n132 71.676
R1267 B.n217 B.n133 71.676
R1268 B.n221 B.n134 71.676
R1269 B.n225 B.n135 71.676
R1270 B.n229 B.n136 71.676
R1271 B.n234 B.n137 71.676
R1272 B.n238 B.n138 71.676
R1273 B.n242 B.n139 71.676
R1274 B.n246 B.n140 71.676
R1275 B.n250 B.n141 71.676
R1276 B.n254 B.n142 71.676
R1277 B.n258 B.n143 71.676
R1278 B.n262 B.n144 71.676
R1279 B.n266 B.n145 71.676
R1280 B.n270 B.n146 71.676
R1281 B.n274 B.n147 71.676
R1282 B.n278 B.n148 71.676
R1283 B.n282 B.n149 71.676
R1284 B.n858 B.n150 71.676
R1285 B.n858 B.n857 71.676
R1286 B.n284 B.n149 71.676
R1287 B.n281 B.n148 71.676
R1288 B.n277 B.n147 71.676
R1289 B.n273 B.n146 71.676
R1290 B.n269 B.n145 71.676
R1291 B.n265 B.n144 71.676
R1292 B.n261 B.n143 71.676
R1293 B.n257 B.n142 71.676
R1294 B.n253 B.n141 71.676
R1295 B.n249 B.n140 71.676
R1296 B.n245 B.n139 71.676
R1297 B.n241 B.n138 71.676
R1298 B.n237 B.n137 71.676
R1299 B.n233 B.n136 71.676
R1300 B.n228 B.n135 71.676
R1301 B.n224 B.n134 71.676
R1302 B.n220 B.n133 71.676
R1303 B.n216 B.n132 71.676
R1304 B.n212 B.n131 71.676
R1305 B.n207 B.n130 71.676
R1306 B.n203 B.n129 71.676
R1307 B.n199 B.n128 71.676
R1308 B.n195 B.n127 71.676
R1309 B.n191 B.n126 71.676
R1310 B.n187 B.n125 71.676
R1311 B.n183 B.n124 71.676
R1312 B.n179 B.n123 71.676
R1313 B.n175 B.n122 71.676
R1314 B.n171 B.n121 71.676
R1315 B.n167 B.n120 71.676
R1316 B.n163 B.n119 71.676
R1317 B.n159 B.n118 71.676
R1318 B.n860 B.n117 71.676
R1319 B.n583 B.n582 71.676
R1320 B.n444 B.n411 71.676
R1321 B.n575 B.n412 71.676
R1322 B.n571 B.n413 71.676
R1323 B.n567 B.n414 71.676
R1324 B.n563 B.n415 71.676
R1325 B.n559 B.n416 71.676
R1326 B.n555 B.n417 71.676
R1327 B.n551 B.n418 71.676
R1328 B.n547 B.n419 71.676
R1329 B.n543 B.n420 71.676
R1330 B.n539 B.n421 71.676
R1331 B.n535 B.n422 71.676
R1332 B.n531 B.n423 71.676
R1333 B.n527 B.n424 71.676
R1334 B.n523 B.n425 71.676
R1335 B.n519 B.n426 71.676
R1336 B.n515 B.n427 71.676
R1337 B.n511 B.n428 71.676
R1338 B.n507 B.n429 71.676
R1339 B.n503 B.n430 71.676
R1340 B.n499 B.n431 71.676
R1341 B.n495 B.n432 71.676
R1342 B.n491 B.n433 71.676
R1343 B.n487 B.n434 71.676
R1344 B.n483 B.n435 71.676
R1345 B.n479 B.n436 71.676
R1346 B.n475 B.n437 71.676
R1347 B.n471 B.n438 71.676
R1348 B.n467 B.n439 71.676
R1349 B.n463 B.n440 71.676
R1350 B.n459 B.n441 71.676
R1351 B.n455 B.n442 71.676
R1352 B.n582 B.n410 71.676
R1353 B.n576 B.n411 71.676
R1354 B.n572 B.n412 71.676
R1355 B.n568 B.n413 71.676
R1356 B.n564 B.n414 71.676
R1357 B.n560 B.n415 71.676
R1358 B.n556 B.n416 71.676
R1359 B.n552 B.n417 71.676
R1360 B.n548 B.n418 71.676
R1361 B.n544 B.n419 71.676
R1362 B.n540 B.n420 71.676
R1363 B.n536 B.n421 71.676
R1364 B.n532 B.n422 71.676
R1365 B.n528 B.n423 71.676
R1366 B.n524 B.n424 71.676
R1367 B.n520 B.n425 71.676
R1368 B.n516 B.n426 71.676
R1369 B.n512 B.n427 71.676
R1370 B.n508 B.n428 71.676
R1371 B.n504 B.n429 71.676
R1372 B.n500 B.n430 71.676
R1373 B.n496 B.n431 71.676
R1374 B.n492 B.n432 71.676
R1375 B.n488 B.n433 71.676
R1376 B.n484 B.n434 71.676
R1377 B.n480 B.n435 71.676
R1378 B.n476 B.n436 71.676
R1379 B.n472 B.n437 71.676
R1380 B.n468 B.n438 71.676
R1381 B.n464 B.n439 71.676
R1382 B.n460 B.n440 71.676
R1383 B.n456 B.n441 71.676
R1384 B.n452 B.n442 71.676
R1385 B.n991 B.n990 71.676
R1386 B.n991 B.n2 71.676
R1387 B.n155 B.n154 60.8975
R1388 B.n153 B.n152 60.8975
R1389 B.n449 B.n448 60.8975
R1390 B.n446 B.n445 60.8975
R1391 B.n210 B.n155 59.5399
R1392 B.n231 B.n153 59.5399
R1393 B.n450 B.n449 59.5399
R1394 B.n447 B.n446 59.5399
R1395 B.n588 B.n407 57.1652
R1396 B.n588 B.n403 57.1652
R1397 B.n594 B.n403 57.1652
R1398 B.n594 B.n399 57.1652
R1399 B.n600 B.n399 57.1652
R1400 B.n600 B.n395 57.1652
R1401 B.n606 B.n395 57.1652
R1402 B.n612 B.n391 57.1652
R1403 B.n612 B.n387 57.1652
R1404 B.n618 B.n387 57.1652
R1405 B.n618 B.n383 57.1652
R1406 B.n624 B.n383 57.1652
R1407 B.n624 B.n379 57.1652
R1408 B.n630 B.n379 57.1652
R1409 B.n630 B.n375 57.1652
R1410 B.n636 B.n375 57.1652
R1411 B.n636 B.n371 57.1652
R1412 B.n643 B.n371 57.1652
R1413 B.n643 B.n642 57.1652
R1414 B.n649 B.n364 57.1652
R1415 B.n655 B.n364 57.1652
R1416 B.n655 B.n360 57.1652
R1417 B.n661 B.n360 57.1652
R1418 B.n661 B.n356 57.1652
R1419 B.n667 B.n356 57.1652
R1420 B.n667 B.n352 57.1652
R1421 B.n673 B.n352 57.1652
R1422 B.n679 B.n348 57.1652
R1423 B.n679 B.n344 57.1652
R1424 B.n685 B.n344 57.1652
R1425 B.n685 B.n340 57.1652
R1426 B.n691 B.n340 57.1652
R1427 B.n691 B.n335 57.1652
R1428 B.n697 B.n335 57.1652
R1429 B.n697 B.n336 57.1652
R1430 B.n703 B.n328 57.1652
R1431 B.n709 B.n328 57.1652
R1432 B.n709 B.n324 57.1652
R1433 B.n715 B.n324 57.1652
R1434 B.n715 B.n320 57.1652
R1435 B.n721 B.n320 57.1652
R1436 B.n721 B.n316 57.1652
R1437 B.n728 B.n316 57.1652
R1438 B.n728 B.n727 57.1652
R1439 B.n734 B.n309 57.1652
R1440 B.n740 B.n309 57.1652
R1441 B.n740 B.n305 57.1652
R1442 B.n746 B.n305 57.1652
R1443 B.n746 B.n301 57.1652
R1444 B.n752 B.n301 57.1652
R1445 B.n752 B.n297 57.1652
R1446 B.n758 B.n297 57.1652
R1447 B.n765 B.n293 57.1652
R1448 B.n765 B.n289 57.1652
R1449 B.n771 B.n289 57.1652
R1450 B.n771 B.n4 57.1652
R1451 B.n989 B.n4 57.1652
R1452 B.n989 B.n988 57.1652
R1453 B.n988 B.n987 57.1652
R1454 B.n987 B.n8 57.1652
R1455 B.n12 B.n8 57.1652
R1456 B.n980 B.n12 57.1652
R1457 B.n980 B.n979 57.1652
R1458 B.n978 B.n16 57.1652
R1459 B.n972 B.n16 57.1652
R1460 B.n972 B.n971 57.1652
R1461 B.n971 B.n970 57.1652
R1462 B.n970 B.n23 57.1652
R1463 B.n964 B.n23 57.1652
R1464 B.n964 B.n963 57.1652
R1465 B.n963 B.n962 57.1652
R1466 B.n956 B.n33 57.1652
R1467 B.n956 B.n955 57.1652
R1468 B.n955 B.n954 57.1652
R1469 B.n954 B.n37 57.1652
R1470 B.n948 B.n37 57.1652
R1471 B.n948 B.n947 57.1652
R1472 B.n947 B.n946 57.1652
R1473 B.n946 B.n44 57.1652
R1474 B.n940 B.n44 57.1652
R1475 B.n939 B.n938 57.1652
R1476 B.n938 B.n51 57.1652
R1477 B.n932 B.n51 57.1652
R1478 B.n932 B.n931 57.1652
R1479 B.n931 B.n930 57.1652
R1480 B.n930 B.n58 57.1652
R1481 B.n924 B.n58 57.1652
R1482 B.n924 B.n923 57.1652
R1483 B.n922 B.n65 57.1652
R1484 B.n916 B.n65 57.1652
R1485 B.n916 B.n915 57.1652
R1486 B.n915 B.n914 57.1652
R1487 B.n914 B.n72 57.1652
R1488 B.n908 B.n72 57.1652
R1489 B.n908 B.n907 57.1652
R1490 B.n907 B.n906 57.1652
R1491 B.n900 B.n82 57.1652
R1492 B.n900 B.n899 57.1652
R1493 B.n899 B.n898 57.1652
R1494 B.n898 B.n86 57.1652
R1495 B.n892 B.n86 57.1652
R1496 B.n892 B.n891 57.1652
R1497 B.n891 B.n890 57.1652
R1498 B.n890 B.n93 57.1652
R1499 B.n884 B.n93 57.1652
R1500 B.n884 B.n883 57.1652
R1501 B.n883 B.n882 57.1652
R1502 B.n882 B.n100 57.1652
R1503 B.n876 B.n875 57.1652
R1504 B.n875 B.n874 57.1652
R1505 B.n874 B.n107 57.1652
R1506 B.n868 B.n107 57.1652
R1507 B.n868 B.n867 57.1652
R1508 B.n867 B.n866 57.1652
R1509 B.n866 B.n114 57.1652
R1510 B.n734 B.t0 54.6432
R1511 B.n962 B.t2 54.6432
R1512 B.n606 B.t11 51.2806
R1513 B.n876 B.t15 51.2806
R1514 B.n336 B.t3 46.2366
R1515 B.t5 B.n939 46.2366
R1516 B.t1 B.n293 41.1927
R1517 B.n979 B.t8 41.1927
R1518 B.n649 B.t9 37.8301
R1519 B.n906 B.t4 37.8301
R1520 B.n585 B.n584 33.5615
R1521 B.n451 B.n405 33.5615
R1522 B.n856 B.n855 33.5615
R1523 B.n863 B.n862 33.5615
R1524 B.n673 B.t7 32.7861
R1525 B.t6 B.n922 32.7861
R1526 B.t7 B.n348 24.3796
R1527 B.n923 B.t6 24.3796
R1528 B.n642 B.t9 19.3356
R1529 B.n82 B.t4 19.3356
R1530 B B.n992 18.0485
R1531 B.n758 B.t1 15.973
R1532 B.t8 B.n978 15.973
R1533 B.n703 B.t3 10.929
R1534 B.n940 B.t5 10.929
R1535 B.n586 B.n585 10.6151
R1536 B.n586 B.n401 10.6151
R1537 B.n596 B.n401 10.6151
R1538 B.n597 B.n596 10.6151
R1539 B.n598 B.n597 10.6151
R1540 B.n598 B.n393 10.6151
R1541 B.n608 B.n393 10.6151
R1542 B.n609 B.n608 10.6151
R1543 B.n610 B.n609 10.6151
R1544 B.n610 B.n385 10.6151
R1545 B.n620 B.n385 10.6151
R1546 B.n621 B.n620 10.6151
R1547 B.n622 B.n621 10.6151
R1548 B.n622 B.n377 10.6151
R1549 B.n632 B.n377 10.6151
R1550 B.n633 B.n632 10.6151
R1551 B.n634 B.n633 10.6151
R1552 B.n634 B.n369 10.6151
R1553 B.n645 B.n369 10.6151
R1554 B.n646 B.n645 10.6151
R1555 B.n647 B.n646 10.6151
R1556 B.n647 B.n362 10.6151
R1557 B.n657 B.n362 10.6151
R1558 B.n658 B.n657 10.6151
R1559 B.n659 B.n658 10.6151
R1560 B.n659 B.n354 10.6151
R1561 B.n669 B.n354 10.6151
R1562 B.n670 B.n669 10.6151
R1563 B.n671 B.n670 10.6151
R1564 B.n671 B.n346 10.6151
R1565 B.n681 B.n346 10.6151
R1566 B.n682 B.n681 10.6151
R1567 B.n683 B.n682 10.6151
R1568 B.n683 B.n338 10.6151
R1569 B.n693 B.n338 10.6151
R1570 B.n694 B.n693 10.6151
R1571 B.n695 B.n694 10.6151
R1572 B.n695 B.n330 10.6151
R1573 B.n705 B.n330 10.6151
R1574 B.n706 B.n705 10.6151
R1575 B.n707 B.n706 10.6151
R1576 B.n707 B.n322 10.6151
R1577 B.n717 B.n322 10.6151
R1578 B.n718 B.n717 10.6151
R1579 B.n719 B.n718 10.6151
R1580 B.n719 B.n314 10.6151
R1581 B.n730 B.n314 10.6151
R1582 B.n731 B.n730 10.6151
R1583 B.n732 B.n731 10.6151
R1584 B.n732 B.n307 10.6151
R1585 B.n742 B.n307 10.6151
R1586 B.n743 B.n742 10.6151
R1587 B.n744 B.n743 10.6151
R1588 B.n744 B.n299 10.6151
R1589 B.n754 B.n299 10.6151
R1590 B.n755 B.n754 10.6151
R1591 B.n756 B.n755 10.6151
R1592 B.n756 B.n291 10.6151
R1593 B.n767 B.n291 10.6151
R1594 B.n768 B.n767 10.6151
R1595 B.n769 B.n768 10.6151
R1596 B.n769 B.n0 10.6151
R1597 B.n584 B.n409 10.6151
R1598 B.n579 B.n409 10.6151
R1599 B.n579 B.n578 10.6151
R1600 B.n578 B.n577 10.6151
R1601 B.n577 B.n574 10.6151
R1602 B.n574 B.n573 10.6151
R1603 B.n573 B.n570 10.6151
R1604 B.n570 B.n569 10.6151
R1605 B.n569 B.n566 10.6151
R1606 B.n566 B.n565 10.6151
R1607 B.n565 B.n562 10.6151
R1608 B.n562 B.n561 10.6151
R1609 B.n561 B.n558 10.6151
R1610 B.n558 B.n557 10.6151
R1611 B.n557 B.n554 10.6151
R1612 B.n554 B.n553 10.6151
R1613 B.n553 B.n550 10.6151
R1614 B.n550 B.n549 10.6151
R1615 B.n549 B.n546 10.6151
R1616 B.n546 B.n545 10.6151
R1617 B.n545 B.n542 10.6151
R1618 B.n542 B.n541 10.6151
R1619 B.n541 B.n538 10.6151
R1620 B.n538 B.n537 10.6151
R1621 B.n537 B.n534 10.6151
R1622 B.n534 B.n533 10.6151
R1623 B.n533 B.n530 10.6151
R1624 B.n530 B.n529 10.6151
R1625 B.n526 B.n525 10.6151
R1626 B.n525 B.n522 10.6151
R1627 B.n522 B.n521 10.6151
R1628 B.n521 B.n518 10.6151
R1629 B.n518 B.n517 10.6151
R1630 B.n517 B.n514 10.6151
R1631 B.n514 B.n513 10.6151
R1632 B.n513 B.n510 10.6151
R1633 B.n510 B.n509 10.6151
R1634 B.n506 B.n505 10.6151
R1635 B.n505 B.n502 10.6151
R1636 B.n502 B.n501 10.6151
R1637 B.n501 B.n498 10.6151
R1638 B.n498 B.n497 10.6151
R1639 B.n497 B.n494 10.6151
R1640 B.n494 B.n493 10.6151
R1641 B.n493 B.n490 10.6151
R1642 B.n490 B.n489 10.6151
R1643 B.n489 B.n486 10.6151
R1644 B.n486 B.n485 10.6151
R1645 B.n485 B.n482 10.6151
R1646 B.n482 B.n481 10.6151
R1647 B.n481 B.n478 10.6151
R1648 B.n478 B.n477 10.6151
R1649 B.n477 B.n474 10.6151
R1650 B.n474 B.n473 10.6151
R1651 B.n473 B.n470 10.6151
R1652 B.n470 B.n469 10.6151
R1653 B.n469 B.n466 10.6151
R1654 B.n466 B.n465 10.6151
R1655 B.n465 B.n462 10.6151
R1656 B.n462 B.n461 10.6151
R1657 B.n461 B.n458 10.6151
R1658 B.n458 B.n457 10.6151
R1659 B.n457 B.n454 10.6151
R1660 B.n454 B.n453 10.6151
R1661 B.n453 B.n451 10.6151
R1662 B.n590 B.n405 10.6151
R1663 B.n591 B.n590 10.6151
R1664 B.n592 B.n591 10.6151
R1665 B.n592 B.n397 10.6151
R1666 B.n602 B.n397 10.6151
R1667 B.n603 B.n602 10.6151
R1668 B.n604 B.n603 10.6151
R1669 B.n604 B.n389 10.6151
R1670 B.n614 B.n389 10.6151
R1671 B.n615 B.n614 10.6151
R1672 B.n616 B.n615 10.6151
R1673 B.n616 B.n381 10.6151
R1674 B.n626 B.n381 10.6151
R1675 B.n627 B.n626 10.6151
R1676 B.n628 B.n627 10.6151
R1677 B.n628 B.n373 10.6151
R1678 B.n638 B.n373 10.6151
R1679 B.n639 B.n638 10.6151
R1680 B.n640 B.n639 10.6151
R1681 B.n640 B.n366 10.6151
R1682 B.n651 B.n366 10.6151
R1683 B.n652 B.n651 10.6151
R1684 B.n653 B.n652 10.6151
R1685 B.n653 B.n358 10.6151
R1686 B.n663 B.n358 10.6151
R1687 B.n664 B.n663 10.6151
R1688 B.n665 B.n664 10.6151
R1689 B.n665 B.n350 10.6151
R1690 B.n675 B.n350 10.6151
R1691 B.n676 B.n675 10.6151
R1692 B.n677 B.n676 10.6151
R1693 B.n677 B.n342 10.6151
R1694 B.n687 B.n342 10.6151
R1695 B.n688 B.n687 10.6151
R1696 B.n689 B.n688 10.6151
R1697 B.n689 B.n333 10.6151
R1698 B.n699 B.n333 10.6151
R1699 B.n700 B.n699 10.6151
R1700 B.n701 B.n700 10.6151
R1701 B.n701 B.n326 10.6151
R1702 B.n711 B.n326 10.6151
R1703 B.n712 B.n711 10.6151
R1704 B.n713 B.n712 10.6151
R1705 B.n713 B.n318 10.6151
R1706 B.n723 B.n318 10.6151
R1707 B.n724 B.n723 10.6151
R1708 B.n725 B.n724 10.6151
R1709 B.n725 B.n311 10.6151
R1710 B.n736 B.n311 10.6151
R1711 B.n737 B.n736 10.6151
R1712 B.n738 B.n737 10.6151
R1713 B.n738 B.n303 10.6151
R1714 B.n748 B.n303 10.6151
R1715 B.n749 B.n748 10.6151
R1716 B.n750 B.n749 10.6151
R1717 B.n750 B.n295 10.6151
R1718 B.n760 B.n295 10.6151
R1719 B.n761 B.n760 10.6151
R1720 B.n763 B.n761 10.6151
R1721 B.n763 B.n762 10.6151
R1722 B.n762 B.n287 10.6151
R1723 B.n774 B.n287 10.6151
R1724 B.n775 B.n774 10.6151
R1725 B.n776 B.n775 10.6151
R1726 B.n777 B.n776 10.6151
R1727 B.n778 B.n777 10.6151
R1728 B.n781 B.n778 10.6151
R1729 B.n782 B.n781 10.6151
R1730 B.n783 B.n782 10.6151
R1731 B.n784 B.n783 10.6151
R1732 B.n786 B.n784 10.6151
R1733 B.n787 B.n786 10.6151
R1734 B.n788 B.n787 10.6151
R1735 B.n789 B.n788 10.6151
R1736 B.n791 B.n789 10.6151
R1737 B.n792 B.n791 10.6151
R1738 B.n793 B.n792 10.6151
R1739 B.n794 B.n793 10.6151
R1740 B.n796 B.n794 10.6151
R1741 B.n797 B.n796 10.6151
R1742 B.n798 B.n797 10.6151
R1743 B.n799 B.n798 10.6151
R1744 B.n801 B.n799 10.6151
R1745 B.n802 B.n801 10.6151
R1746 B.n803 B.n802 10.6151
R1747 B.n804 B.n803 10.6151
R1748 B.n806 B.n804 10.6151
R1749 B.n807 B.n806 10.6151
R1750 B.n808 B.n807 10.6151
R1751 B.n809 B.n808 10.6151
R1752 B.n811 B.n809 10.6151
R1753 B.n812 B.n811 10.6151
R1754 B.n813 B.n812 10.6151
R1755 B.n814 B.n813 10.6151
R1756 B.n816 B.n814 10.6151
R1757 B.n817 B.n816 10.6151
R1758 B.n818 B.n817 10.6151
R1759 B.n819 B.n818 10.6151
R1760 B.n821 B.n819 10.6151
R1761 B.n822 B.n821 10.6151
R1762 B.n823 B.n822 10.6151
R1763 B.n824 B.n823 10.6151
R1764 B.n826 B.n824 10.6151
R1765 B.n827 B.n826 10.6151
R1766 B.n828 B.n827 10.6151
R1767 B.n829 B.n828 10.6151
R1768 B.n831 B.n829 10.6151
R1769 B.n832 B.n831 10.6151
R1770 B.n833 B.n832 10.6151
R1771 B.n834 B.n833 10.6151
R1772 B.n836 B.n834 10.6151
R1773 B.n837 B.n836 10.6151
R1774 B.n838 B.n837 10.6151
R1775 B.n839 B.n838 10.6151
R1776 B.n841 B.n839 10.6151
R1777 B.n842 B.n841 10.6151
R1778 B.n843 B.n842 10.6151
R1779 B.n844 B.n843 10.6151
R1780 B.n846 B.n844 10.6151
R1781 B.n847 B.n846 10.6151
R1782 B.n848 B.n847 10.6151
R1783 B.n849 B.n848 10.6151
R1784 B.n851 B.n849 10.6151
R1785 B.n852 B.n851 10.6151
R1786 B.n853 B.n852 10.6151
R1787 B.n854 B.n853 10.6151
R1788 B.n855 B.n854 10.6151
R1789 B.n984 B.n1 10.6151
R1790 B.n984 B.n983 10.6151
R1791 B.n983 B.n982 10.6151
R1792 B.n982 B.n10 10.6151
R1793 B.n976 B.n10 10.6151
R1794 B.n976 B.n975 10.6151
R1795 B.n975 B.n974 10.6151
R1796 B.n974 B.n18 10.6151
R1797 B.n968 B.n18 10.6151
R1798 B.n968 B.n967 10.6151
R1799 B.n967 B.n966 10.6151
R1800 B.n966 B.n25 10.6151
R1801 B.n960 B.n25 10.6151
R1802 B.n960 B.n959 10.6151
R1803 B.n959 B.n958 10.6151
R1804 B.n958 B.n31 10.6151
R1805 B.n952 B.n31 10.6151
R1806 B.n952 B.n951 10.6151
R1807 B.n951 B.n950 10.6151
R1808 B.n950 B.n39 10.6151
R1809 B.n944 B.n39 10.6151
R1810 B.n944 B.n943 10.6151
R1811 B.n943 B.n942 10.6151
R1812 B.n942 B.n46 10.6151
R1813 B.n936 B.n46 10.6151
R1814 B.n936 B.n935 10.6151
R1815 B.n935 B.n934 10.6151
R1816 B.n934 B.n53 10.6151
R1817 B.n928 B.n53 10.6151
R1818 B.n928 B.n927 10.6151
R1819 B.n927 B.n926 10.6151
R1820 B.n926 B.n60 10.6151
R1821 B.n920 B.n60 10.6151
R1822 B.n920 B.n919 10.6151
R1823 B.n919 B.n918 10.6151
R1824 B.n918 B.n67 10.6151
R1825 B.n912 B.n67 10.6151
R1826 B.n912 B.n911 10.6151
R1827 B.n911 B.n910 10.6151
R1828 B.n910 B.n74 10.6151
R1829 B.n904 B.n74 10.6151
R1830 B.n904 B.n903 10.6151
R1831 B.n903 B.n902 10.6151
R1832 B.n902 B.n80 10.6151
R1833 B.n896 B.n80 10.6151
R1834 B.n896 B.n895 10.6151
R1835 B.n895 B.n894 10.6151
R1836 B.n894 B.n88 10.6151
R1837 B.n888 B.n88 10.6151
R1838 B.n888 B.n887 10.6151
R1839 B.n887 B.n886 10.6151
R1840 B.n886 B.n95 10.6151
R1841 B.n880 B.n95 10.6151
R1842 B.n880 B.n879 10.6151
R1843 B.n879 B.n878 10.6151
R1844 B.n878 B.n102 10.6151
R1845 B.n872 B.n102 10.6151
R1846 B.n872 B.n871 10.6151
R1847 B.n871 B.n870 10.6151
R1848 B.n870 B.n109 10.6151
R1849 B.n864 B.n109 10.6151
R1850 B.n864 B.n863 10.6151
R1851 B.n862 B.n116 10.6151
R1852 B.n157 B.n116 10.6151
R1853 B.n158 B.n157 10.6151
R1854 B.n161 B.n158 10.6151
R1855 B.n162 B.n161 10.6151
R1856 B.n165 B.n162 10.6151
R1857 B.n166 B.n165 10.6151
R1858 B.n169 B.n166 10.6151
R1859 B.n170 B.n169 10.6151
R1860 B.n173 B.n170 10.6151
R1861 B.n174 B.n173 10.6151
R1862 B.n177 B.n174 10.6151
R1863 B.n178 B.n177 10.6151
R1864 B.n181 B.n178 10.6151
R1865 B.n182 B.n181 10.6151
R1866 B.n185 B.n182 10.6151
R1867 B.n186 B.n185 10.6151
R1868 B.n189 B.n186 10.6151
R1869 B.n190 B.n189 10.6151
R1870 B.n193 B.n190 10.6151
R1871 B.n194 B.n193 10.6151
R1872 B.n197 B.n194 10.6151
R1873 B.n198 B.n197 10.6151
R1874 B.n201 B.n198 10.6151
R1875 B.n202 B.n201 10.6151
R1876 B.n205 B.n202 10.6151
R1877 B.n206 B.n205 10.6151
R1878 B.n209 B.n206 10.6151
R1879 B.n214 B.n211 10.6151
R1880 B.n215 B.n214 10.6151
R1881 B.n218 B.n215 10.6151
R1882 B.n219 B.n218 10.6151
R1883 B.n222 B.n219 10.6151
R1884 B.n223 B.n222 10.6151
R1885 B.n226 B.n223 10.6151
R1886 B.n227 B.n226 10.6151
R1887 B.n230 B.n227 10.6151
R1888 B.n235 B.n232 10.6151
R1889 B.n236 B.n235 10.6151
R1890 B.n239 B.n236 10.6151
R1891 B.n240 B.n239 10.6151
R1892 B.n243 B.n240 10.6151
R1893 B.n244 B.n243 10.6151
R1894 B.n247 B.n244 10.6151
R1895 B.n248 B.n247 10.6151
R1896 B.n251 B.n248 10.6151
R1897 B.n252 B.n251 10.6151
R1898 B.n255 B.n252 10.6151
R1899 B.n256 B.n255 10.6151
R1900 B.n259 B.n256 10.6151
R1901 B.n260 B.n259 10.6151
R1902 B.n263 B.n260 10.6151
R1903 B.n264 B.n263 10.6151
R1904 B.n267 B.n264 10.6151
R1905 B.n268 B.n267 10.6151
R1906 B.n271 B.n268 10.6151
R1907 B.n272 B.n271 10.6151
R1908 B.n275 B.n272 10.6151
R1909 B.n276 B.n275 10.6151
R1910 B.n279 B.n276 10.6151
R1911 B.n280 B.n279 10.6151
R1912 B.n283 B.n280 10.6151
R1913 B.n285 B.n283 10.6151
R1914 B.n286 B.n285 10.6151
R1915 B.n856 B.n286 10.6151
R1916 B.n529 B.n447 9.36635
R1917 B.n506 B.n450 9.36635
R1918 B.n210 B.n209 9.36635
R1919 B.n232 B.n231 9.36635
R1920 B.n992 B.n0 8.11757
R1921 B.n992 B.n1 8.11757
R1922 B.t11 B.n391 5.8851
R1923 B.t15 B.n100 5.8851
R1924 B.n727 B.t0 2.52247
R1925 B.n33 B.t2 2.52247
R1926 B.n526 B.n447 1.24928
R1927 B.n509 B.n450 1.24928
R1928 B.n211 B.n210 1.24928
R1929 B.n231 B.n230 1.24928
R1930 VP.n26 VP.n23 161.3
R1931 VP.n28 VP.n27 161.3
R1932 VP.n29 VP.n22 161.3
R1933 VP.n31 VP.n30 161.3
R1934 VP.n32 VP.n21 161.3
R1935 VP.n34 VP.n33 161.3
R1936 VP.n36 VP.n20 161.3
R1937 VP.n38 VP.n37 161.3
R1938 VP.n39 VP.n19 161.3
R1939 VP.n41 VP.n40 161.3
R1940 VP.n42 VP.n18 161.3
R1941 VP.n45 VP.n44 161.3
R1942 VP.n46 VP.n17 161.3
R1943 VP.n48 VP.n47 161.3
R1944 VP.n49 VP.n16 161.3
R1945 VP.n51 VP.n50 161.3
R1946 VP.n52 VP.n15 161.3
R1947 VP.n54 VP.n53 161.3
R1948 VP.n55 VP.n14 161.3
R1949 VP.n100 VP.n0 161.3
R1950 VP.n99 VP.n98 161.3
R1951 VP.n97 VP.n1 161.3
R1952 VP.n96 VP.n95 161.3
R1953 VP.n94 VP.n2 161.3
R1954 VP.n93 VP.n92 161.3
R1955 VP.n91 VP.n3 161.3
R1956 VP.n90 VP.n89 161.3
R1957 VP.n87 VP.n4 161.3
R1958 VP.n86 VP.n85 161.3
R1959 VP.n84 VP.n5 161.3
R1960 VP.n83 VP.n82 161.3
R1961 VP.n81 VP.n6 161.3
R1962 VP.n79 VP.n78 161.3
R1963 VP.n77 VP.n7 161.3
R1964 VP.n76 VP.n75 161.3
R1965 VP.n74 VP.n8 161.3
R1966 VP.n73 VP.n72 161.3
R1967 VP.n71 VP.n9 161.3
R1968 VP.n70 VP.n69 161.3
R1969 VP.n67 VP.n10 161.3
R1970 VP.n66 VP.n65 161.3
R1971 VP.n64 VP.n11 161.3
R1972 VP.n63 VP.n62 161.3
R1973 VP.n61 VP.n12 161.3
R1974 VP.n60 VP.n59 161.3
R1975 VP.n58 VP.n13 109.288
R1976 VP.n102 VP.n101 109.288
R1977 VP.n57 VP.n56 109.288
R1978 VP.n25 VP.t2 99.6097
R1979 VP.n13 VP.t8 66.9831
R1980 VP.n68 VP.t6 66.9831
R1981 VP.n80 VP.t9 66.9831
R1982 VP.n88 VP.t7 66.9831
R1983 VP.n101 VP.t4 66.9831
R1984 VP.n56 VP.t3 66.9831
R1985 VP.n43 VP.t0 66.9831
R1986 VP.n35 VP.t5 66.9831
R1987 VP.n24 VP.t1 66.9831
R1988 VP.n75 VP.n74 56.5193
R1989 VP.n41 VP.n19 56.5193
R1990 VP.n86 VP.n5 56.5193
R1991 VP.n30 VP.n29 56.5193
R1992 VP.n25 VP.n24 54.5315
R1993 VP.n58 VP.n57 51.0223
R1994 VP.n66 VP.n11 44.3785
R1995 VP.n95 VP.n94 44.3785
R1996 VP.n50 VP.n49 44.3785
R1997 VP.n62 VP.n11 36.6083
R1998 VP.n95 VP.n1 36.6083
R1999 VP.n50 VP.n15 36.6083
R2000 VP.n61 VP.n60 24.4675
R2001 VP.n62 VP.n61 24.4675
R2002 VP.n67 VP.n66 24.4675
R2003 VP.n69 VP.n67 24.4675
R2004 VP.n73 VP.n9 24.4675
R2005 VP.n74 VP.n73 24.4675
R2006 VP.n75 VP.n7 24.4675
R2007 VP.n79 VP.n7 24.4675
R2008 VP.n82 VP.n81 24.4675
R2009 VP.n82 VP.n5 24.4675
R2010 VP.n87 VP.n86 24.4675
R2011 VP.n89 VP.n87 24.4675
R2012 VP.n93 VP.n3 24.4675
R2013 VP.n94 VP.n93 24.4675
R2014 VP.n99 VP.n1 24.4675
R2015 VP.n100 VP.n99 24.4675
R2016 VP.n54 VP.n15 24.4675
R2017 VP.n55 VP.n54 24.4675
R2018 VP.n42 VP.n41 24.4675
R2019 VP.n44 VP.n42 24.4675
R2020 VP.n48 VP.n17 24.4675
R2021 VP.n49 VP.n48 24.4675
R2022 VP.n30 VP.n21 24.4675
R2023 VP.n34 VP.n21 24.4675
R2024 VP.n37 VP.n36 24.4675
R2025 VP.n37 VP.n19 24.4675
R2026 VP.n28 VP.n23 24.4675
R2027 VP.n29 VP.n28 24.4675
R2028 VP.n68 VP.n9 19.0848
R2029 VP.n89 VP.n88 19.0848
R2030 VP.n44 VP.n43 19.0848
R2031 VP.n24 VP.n23 19.0848
R2032 VP.n80 VP.n79 12.234
R2033 VP.n81 VP.n80 12.234
R2034 VP.n35 VP.n34 12.234
R2035 VP.n36 VP.n35 12.234
R2036 VP.n69 VP.n68 5.38324
R2037 VP.n88 VP.n3 5.38324
R2038 VP.n43 VP.n17 5.38324
R2039 VP.n26 VP.n25 5.13245
R2040 VP.n60 VP.n13 1.46852
R2041 VP.n101 VP.n100 1.46852
R2042 VP.n56 VP.n55 1.46852
R2043 VP.n57 VP.n14 0.278367
R2044 VP.n59 VP.n58 0.278367
R2045 VP.n102 VP.n0 0.278367
R2046 VP.n27 VP.n26 0.189894
R2047 VP.n27 VP.n22 0.189894
R2048 VP.n31 VP.n22 0.189894
R2049 VP.n32 VP.n31 0.189894
R2050 VP.n33 VP.n32 0.189894
R2051 VP.n33 VP.n20 0.189894
R2052 VP.n38 VP.n20 0.189894
R2053 VP.n39 VP.n38 0.189894
R2054 VP.n40 VP.n39 0.189894
R2055 VP.n40 VP.n18 0.189894
R2056 VP.n45 VP.n18 0.189894
R2057 VP.n46 VP.n45 0.189894
R2058 VP.n47 VP.n46 0.189894
R2059 VP.n47 VP.n16 0.189894
R2060 VP.n51 VP.n16 0.189894
R2061 VP.n52 VP.n51 0.189894
R2062 VP.n53 VP.n52 0.189894
R2063 VP.n53 VP.n14 0.189894
R2064 VP.n59 VP.n12 0.189894
R2065 VP.n63 VP.n12 0.189894
R2066 VP.n64 VP.n63 0.189894
R2067 VP.n65 VP.n64 0.189894
R2068 VP.n65 VP.n10 0.189894
R2069 VP.n70 VP.n10 0.189894
R2070 VP.n71 VP.n70 0.189894
R2071 VP.n72 VP.n71 0.189894
R2072 VP.n72 VP.n8 0.189894
R2073 VP.n76 VP.n8 0.189894
R2074 VP.n77 VP.n76 0.189894
R2075 VP.n78 VP.n77 0.189894
R2076 VP.n78 VP.n6 0.189894
R2077 VP.n83 VP.n6 0.189894
R2078 VP.n84 VP.n83 0.189894
R2079 VP.n85 VP.n84 0.189894
R2080 VP.n85 VP.n4 0.189894
R2081 VP.n90 VP.n4 0.189894
R2082 VP.n91 VP.n90 0.189894
R2083 VP.n92 VP.n91 0.189894
R2084 VP.n92 VP.n2 0.189894
R2085 VP.n96 VP.n2 0.189894
R2086 VP.n97 VP.n96 0.189894
R2087 VP.n98 VP.n97 0.189894
R2088 VP.n98 VP.n0 0.189894
R2089 VP VP.n102 0.153454
R2090 VDD1.n1 VDD1.t7 70.2686
R2091 VDD1.n3 VDD1.t1 70.2685
R2092 VDD1.n5 VDD1.n4 67.0013
R2093 VDD1.n7 VDD1.n6 65.0266
R2094 VDD1.n1 VDD1.n0 65.0266
R2095 VDD1.n3 VDD1.n2 65.0265
R2096 VDD1.n7 VDD1.n5 45.2423
R2097 VDD1.n6 VDD1.t9 2.53571
R2098 VDD1.n6 VDD1.t6 2.53571
R2099 VDD1.n0 VDD1.t8 2.53571
R2100 VDD1.n0 VDD1.t4 2.53571
R2101 VDD1.n4 VDD1.t2 2.53571
R2102 VDD1.n4 VDD1.t5 2.53571
R2103 VDD1.n2 VDD1.t3 2.53571
R2104 VDD1.n2 VDD1.t0 2.53571
R2105 VDD1 VDD1.n7 1.97248
R2106 VDD1 VDD1.n1 0.735414
R2107 VDD1.n5 VDD1.n3 0.621878
C0 VDD1 VP 7.68285f
C1 VN VP 7.9334f
C2 VTAIL VP 8.16507f
C3 VDD2 VP 0.609985f
C4 VDD1 VN 0.153773f
C5 VDD1 VTAIL 8.589621f
C6 VTAIL VN 8.15086f
C7 VDD2 VDD1 2.31022f
C8 VDD2 VN 7.22981f
C9 VDD2 VTAIL 8.643089f
C10 VDD2 B 6.755968f
C11 VDD1 B 6.695352f
C12 VTAIL B 6.702909f
C13 VN B 18.81827f
C14 VP B 17.398855f
C15 VDD1.t7 B 1.76932f
C16 VDD1.t8 B 0.16017f
C17 VDD1.t4 B 0.16017f
C18 VDD1.n0 B 1.37464f
C19 VDD1.n1 B 0.99766f
C20 VDD1.t1 B 1.76931f
C21 VDD1.t3 B 0.16017f
C22 VDD1.t0 B 0.16017f
C23 VDD1.n2 B 1.37464f
C24 VDD1.n3 B 0.989143f
C25 VDD1.t2 B 0.16017f
C26 VDD1.t5 B 0.16017f
C27 VDD1.n4 B 1.39285f
C28 VDD1.n5 B 2.99772f
C29 VDD1.t9 B 0.16017f
C30 VDD1.t6 B 0.16017f
C31 VDD1.n6 B 1.37464f
C32 VDD1.n7 B 3.05235f
C33 VP.n0 B 0.029258f
C34 VP.t4 B 1.30663f
C35 VP.n1 B 0.044745f
C36 VP.n2 B 0.022192f
C37 VP.n3 B 0.025433f
C38 VP.n4 B 0.022192f
C39 VP.n5 B 0.036725f
C40 VP.n6 B 0.022192f
C41 VP.t9 B 1.30663f
C42 VP.n7 B 0.041361f
C43 VP.n8 B 0.022192f
C44 VP.n9 B 0.036868f
C45 VP.n10 B 0.022192f
C46 VP.n11 B 0.0184f
C47 VP.n12 B 0.022192f
C48 VP.t8 B 1.30663f
C49 VP.n13 B 0.545786f
C50 VP.n14 B 0.029258f
C51 VP.t3 B 1.30663f
C52 VP.n15 B 0.044745f
C53 VP.n16 B 0.022192f
C54 VP.n17 B 0.025433f
C55 VP.n18 B 0.022192f
C56 VP.n19 B 0.036725f
C57 VP.n20 B 0.022192f
C58 VP.t5 B 1.30663f
C59 VP.n21 B 0.041361f
C60 VP.n22 B 0.022192f
C61 VP.n23 B 0.036868f
C62 VP.t2 B 1.5108f
C63 VP.t1 B 1.30663f
C64 VP.n24 B 0.54957f
C65 VP.n25 B 0.523903f
C66 VP.n26 B 0.233187f
C67 VP.n27 B 0.022192f
C68 VP.n28 B 0.041361f
C69 VP.n29 B 0.028068f
C70 VP.n30 B 0.036725f
C71 VP.n31 B 0.022192f
C72 VP.n32 B 0.022192f
C73 VP.n33 B 0.022192f
C74 VP.n34 B 0.031151f
C75 VP.n35 B 0.475382f
C76 VP.n36 B 0.031151f
C77 VP.n37 B 0.041361f
C78 VP.n38 B 0.022192f
C79 VP.n39 B 0.022192f
C80 VP.n40 B 0.022192f
C81 VP.n41 B 0.028068f
C82 VP.n42 B 0.041361f
C83 VP.t0 B 1.30663f
C84 VP.n43 B 0.475382f
C85 VP.n44 B 0.036868f
C86 VP.n45 B 0.022192f
C87 VP.n46 B 0.022192f
C88 VP.n47 B 0.022192f
C89 VP.n48 B 0.041361f
C90 VP.n49 B 0.043008f
C91 VP.n50 B 0.0184f
C92 VP.n51 B 0.022192f
C93 VP.n52 B 0.022192f
C94 VP.n53 B 0.022192f
C95 VP.n54 B 0.041361f
C96 VP.n55 B 0.022166f
C97 VP.n56 B 0.545786f
C98 VP.n57 B 1.27757f
C99 VP.n58 B 1.29321f
C100 VP.n59 B 0.029258f
C101 VP.n60 B 0.022166f
C102 VP.n61 B 0.041361f
C103 VP.n62 B 0.044745f
C104 VP.n63 B 0.022192f
C105 VP.n64 B 0.022192f
C106 VP.n65 B 0.022192f
C107 VP.n66 B 0.043008f
C108 VP.n67 B 0.041361f
C109 VP.t6 B 1.30663f
C110 VP.n68 B 0.475382f
C111 VP.n69 B 0.025433f
C112 VP.n70 B 0.022192f
C113 VP.n71 B 0.022192f
C114 VP.n72 B 0.022192f
C115 VP.n73 B 0.041361f
C116 VP.n74 B 0.028068f
C117 VP.n75 B 0.036725f
C118 VP.n76 B 0.022192f
C119 VP.n77 B 0.022192f
C120 VP.n78 B 0.022192f
C121 VP.n79 B 0.031151f
C122 VP.n80 B 0.475382f
C123 VP.n81 B 0.031151f
C124 VP.n82 B 0.041361f
C125 VP.n83 B 0.022192f
C126 VP.n84 B 0.022192f
C127 VP.n85 B 0.022192f
C128 VP.n86 B 0.028068f
C129 VP.n87 B 0.041361f
C130 VP.t7 B 1.30663f
C131 VP.n88 B 0.475382f
C132 VP.n89 B 0.036868f
C133 VP.n90 B 0.022192f
C134 VP.n91 B 0.022192f
C135 VP.n92 B 0.022192f
C136 VP.n93 B 0.041361f
C137 VP.n94 B 0.043008f
C138 VP.n95 B 0.0184f
C139 VP.n96 B 0.022192f
C140 VP.n97 B 0.022192f
C141 VP.n98 B 0.022192f
C142 VP.n99 B 0.041361f
C143 VP.n100 B 0.022166f
C144 VP.n101 B 0.545786f
C145 VP.n102 B 0.042127f
C146 VTAIL.t16 B 0.167032f
C147 VTAIL.t14 B 0.167032f
C148 VTAIL.n0 B 1.3578f
C149 VTAIL.n1 B 0.604729f
C150 VTAIL.t1 B 1.73131f
C151 VTAIL.n2 B 0.740703f
C152 VTAIL.t3 B 0.167032f
C153 VTAIL.t0 B 0.167032f
C154 VTAIL.n3 B 1.3578f
C155 VTAIL.n4 B 0.735727f
C156 VTAIL.t9 B 0.167032f
C157 VTAIL.t7 B 0.167032f
C158 VTAIL.n5 B 1.3578f
C159 VTAIL.n6 B 1.92656f
C160 VTAIL.t18 B 0.167032f
C161 VTAIL.t19 B 0.167032f
C162 VTAIL.n7 B 1.3578f
C163 VTAIL.n8 B 1.92656f
C164 VTAIL.t11 B 0.167032f
C165 VTAIL.t12 B 0.167032f
C166 VTAIL.n9 B 1.3578f
C167 VTAIL.n10 B 0.735724f
C168 VTAIL.t13 B 1.73132f
C169 VTAIL.n11 B 0.740692f
C170 VTAIL.t8 B 0.167032f
C171 VTAIL.t2 B 0.167032f
C172 VTAIL.n12 B 1.3578f
C173 VTAIL.n13 B 0.658667f
C174 VTAIL.t5 B 0.167032f
C175 VTAIL.t6 B 0.167032f
C176 VTAIL.n14 B 1.3578f
C177 VTAIL.n15 B 0.735724f
C178 VTAIL.t4 B 1.73132f
C179 VTAIL.n16 B 1.77253f
C180 VTAIL.t10 B 1.73131f
C181 VTAIL.n17 B 1.77254f
C182 VTAIL.t17 B 0.167032f
C183 VTAIL.t15 B 0.167032f
C184 VTAIL.n18 B 1.3578f
C185 VTAIL.n19 B 0.553608f
C186 VDD2.t1 B 1.73067f
C187 VDD2.t6 B 0.156672f
C188 VDD2.t3 B 0.156672f
C189 VDD2.n0 B 1.34462f
C190 VDD2.n1 B 0.967539f
C191 VDD2.t0 B 0.156672f
C192 VDD2.t9 B 0.156672f
C193 VDD2.n2 B 1.36243f
C194 VDD2.n3 B 2.80288f
C195 VDD2.t4 B 1.7113f
C196 VDD2.n4 B 2.92059f
C197 VDD2.t2 B 0.156672f
C198 VDD2.t7 B 0.156672f
C199 VDD2.n5 B 1.34462f
C200 VDD2.n6 B 0.492263f
C201 VDD2.t8 B 0.156672f
C202 VDD2.t5 B 0.156672f
C203 VDD2.n7 B 1.36239f
C204 VN.n0 B 0.028606f
C205 VN.t9 B 1.27751f
C206 VN.n1 B 0.043748f
C207 VN.n2 B 0.021697f
C208 VN.n3 B 0.024866f
C209 VN.n4 B 0.021697f
C210 VN.n5 B 0.035907f
C211 VN.n6 B 0.021697f
C212 VN.t2 B 1.27751f
C213 VN.n7 B 0.040439f
C214 VN.n8 B 0.021697f
C215 VN.n9 B 0.036046f
C216 VN.t3 B 1.47713f
C217 VN.t5 B 1.27751f
C218 VN.n10 B 0.53732f
C219 VN.n11 B 0.512225f
C220 VN.n12 B 0.22799f
C221 VN.n13 B 0.021697f
C222 VN.n14 B 0.040439f
C223 VN.n15 B 0.027442f
C224 VN.n16 B 0.035907f
C225 VN.n17 B 0.021697f
C226 VN.n18 B 0.021697f
C227 VN.n19 B 0.021697f
C228 VN.n20 B 0.030456f
C229 VN.n21 B 0.464786f
C230 VN.n22 B 0.030456f
C231 VN.n23 B 0.040439f
C232 VN.n24 B 0.021697f
C233 VN.n25 B 0.021697f
C234 VN.n26 B 0.021697f
C235 VN.n27 B 0.027442f
C236 VN.n28 B 0.040439f
C237 VN.t4 B 1.27751f
C238 VN.n29 B 0.464786f
C239 VN.n30 B 0.036046f
C240 VN.n31 B 0.021697f
C241 VN.n32 B 0.021697f
C242 VN.n33 B 0.021697f
C243 VN.n34 B 0.040439f
C244 VN.n35 B 0.042049f
C245 VN.n36 B 0.01799f
C246 VN.n37 B 0.021697f
C247 VN.n38 B 0.021697f
C248 VN.n39 B 0.021697f
C249 VN.n40 B 0.040439f
C250 VN.n41 B 0.021672f
C251 VN.n42 B 0.53362f
C252 VN.n43 B 0.041189f
C253 VN.n44 B 0.028606f
C254 VN.t1 B 1.27751f
C255 VN.n45 B 0.043748f
C256 VN.n46 B 0.021697f
C257 VN.n47 B 0.024866f
C258 VN.n48 B 0.021697f
C259 VN.t0 B 1.27751f
C260 VN.n49 B 0.464786f
C261 VN.n50 B 0.035907f
C262 VN.n51 B 0.021697f
C263 VN.t8 B 1.27751f
C264 VN.n52 B 0.040439f
C265 VN.n53 B 0.021697f
C266 VN.n54 B 0.036046f
C267 VN.t6 B 1.47713f
C268 VN.t7 B 1.27751f
C269 VN.n55 B 0.53732f
C270 VN.n56 B 0.512225f
C271 VN.n57 B 0.22799f
C272 VN.n58 B 0.021697f
C273 VN.n59 B 0.040439f
C274 VN.n60 B 0.027442f
C275 VN.n61 B 0.035907f
C276 VN.n62 B 0.021697f
C277 VN.n63 B 0.021697f
C278 VN.n64 B 0.021697f
C279 VN.n65 B 0.030456f
C280 VN.n66 B 0.464786f
C281 VN.n67 B 0.030456f
C282 VN.n68 B 0.040439f
C283 VN.n69 B 0.021697f
C284 VN.n70 B 0.021697f
C285 VN.n71 B 0.021697f
C286 VN.n72 B 0.027442f
C287 VN.n73 B 0.040439f
C288 VN.n74 B 0.036046f
C289 VN.n75 B 0.021697f
C290 VN.n76 B 0.021697f
C291 VN.n77 B 0.021697f
C292 VN.n78 B 0.040439f
C293 VN.n79 B 0.042049f
C294 VN.n80 B 0.01799f
C295 VN.n81 B 0.021697f
C296 VN.n82 B 0.021697f
C297 VN.n83 B 0.021697f
C298 VN.n84 B 0.040439f
C299 VN.n85 B 0.021672f
C300 VN.n86 B 0.53362f
C301 VN.n87 B 1.26072f
.ends

