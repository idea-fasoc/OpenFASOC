* NGSPICE file created from diff_pair_sample_1622.ext - technology: sky130A

.subckt diff_pair_sample_1622 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=2.9733 ps=18.35 w=18.02 l=1.79
X1 B.t11 B.t9 B.t10 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=0 ps=0 w=18.02 l=1.79
X2 B.t8 B.t6 B.t7 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=0 ps=0 w=18.02 l=1.79
X3 B.t5 B.t3 B.t4 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=0 ps=0 w=18.02 l=1.79
X4 VDD2.t5 VN.t0 VTAIL.t2 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=7.0278 ps=36.82 w=18.02 l=1.79
X5 VDD2.t4 VN.t1 VTAIL.t1 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=2.9733 ps=18.35 w=18.02 l=1.79
X6 VTAIL.t4 VN.t2 VDD2.t3 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=2.9733 ps=18.35 w=18.02 l=1.79
X7 VTAIL.t7 VP.t1 VDD1.t4 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=2.9733 ps=18.35 w=18.02 l=1.79
X8 VDD1.t3 VP.t2 VTAIL.t11 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=7.0278 ps=36.82 w=18.02 l=1.79
X9 VDD1.t2 VP.t3 VTAIL.t8 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=2.9733 ps=18.35 w=18.02 l=1.79
X10 VDD1.t1 VP.t4 VTAIL.t10 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=7.0278 ps=36.82 w=18.02 l=1.79
X11 B.t2 B.t0 B.t1 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=0 ps=0 w=18.02 l=1.79
X12 VTAIL.t9 VP.t5 VDD1.t0 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=2.9733 ps=18.35 w=18.02 l=1.79
X13 VDD2.t2 VN.t3 VTAIL.t0 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=7.0278 ps=36.82 w=18.02 l=1.79
X14 VDD2.t1 VN.t4 VTAIL.t3 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=7.0278 pd=36.82 as=2.9733 ps=18.35 w=18.02 l=1.79
X15 VTAIL.t5 VN.t5 VDD2.t0 w_n2666_n4572# sky130_fd_pr__pfet_01v8 ad=2.9733 pd=18.35 as=2.9733 ps=18.35 w=18.02 l=1.79
R0 VP.n7 VP.t3 278.62
R1 VP.n25 VP.t1 242.617
R2 VP.n18 VP.t0 242.617
R3 VP.n32 VP.t2 242.617
R4 VP.n8 VP.t5 242.617
R5 VP.n15 VP.t4 242.617
R6 VP.n18 VP.n17 179.99
R7 VP.n33 VP.n32 179.99
R8 VP.n16 VP.n15 179.99
R9 VP.n10 VP.n9 161.3
R10 VP.n11 VP.n6 161.3
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n5 161.3
R13 VP.n31 VP.n0 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n1 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n2 161.3
R18 VP.n24 VP.n23 161.3
R19 VP.n22 VP.n3 161.3
R20 VP.n21 VP.n20 161.3
R21 VP.n19 VP.n4 161.3
R22 VP.n17 VP.n16 49.9929
R23 VP.n20 VP.n3 46.3896
R24 VP.n30 VP.n1 46.3896
R25 VP.n13 VP.n6 46.3896
R26 VP.n8 VP.n7 44.58
R27 VP.n24 VP.n3 34.7644
R28 VP.n26 VP.n1 34.7644
R29 VP.n9 VP.n6 34.7644
R30 VP.n20 VP.n19 24.5923
R31 VP.n25 VP.n24 24.5923
R32 VP.n26 VP.n25 24.5923
R33 VP.n31 VP.n30 24.5923
R34 VP.n14 VP.n13 24.5923
R35 VP.n9 VP.n8 24.5923
R36 VP.n10 VP.n7 12.1133
R37 VP.n19 VP.n18 5.90254
R38 VP.n32 VP.n31 5.90254
R39 VP.n15 VP.n14 5.90254
R40 VP.n11 VP.n10 0.189894
R41 VP.n12 VP.n11 0.189894
R42 VP.n12 VP.n5 0.189894
R43 VP.n16 VP.n5 0.189894
R44 VP.n17 VP.n4 0.189894
R45 VP.n21 VP.n4 0.189894
R46 VP.n22 VP.n21 0.189894
R47 VP.n23 VP.n22 0.189894
R48 VP.n23 VP.n2 0.189894
R49 VP.n27 VP.n2 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n29 VP.n28 0.189894
R52 VP.n29 VP.n0 0.189894
R53 VP.n33 VP.n0 0.189894
R54 VP VP.n33 0.0516364
R55 VTAIL.n7 VTAIL.t2 56.6909
R56 VTAIL.n11 VTAIL.t0 56.6906
R57 VTAIL.n2 VTAIL.t11 56.6906
R58 VTAIL.n10 VTAIL.t10 56.6906
R59 VTAIL.n9 VTAIL.n8 54.8871
R60 VTAIL.n6 VTAIL.n5 54.8871
R61 VTAIL.n1 VTAIL.n0 54.8868
R62 VTAIL.n4 VTAIL.n3 54.8868
R63 VTAIL.n6 VTAIL.n4 31.5565
R64 VTAIL.n11 VTAIL.n10 29.7289
R65 VTAIL.n7 VTAIL.n6 1.82809
R66 VTAIL.n10 VTAIL.n9 1.82809
R67 VTAIL.n4 VTAIL.n2 1.82809
R68 VTAIL.n0 VTAIL.t3 1.80433
R69 VTAIL.n0 VTAIL.t5 1.80433
R70 VTAIL.n3 VTAIL.t6 1.80433
R71 VTAIL.n3 VTAIL.t7 1.80433
R72 VTAIL.n8 VTAIL.t8 1.80433
R73 VTAIL.n8 VTAIL.t9 1.80433
R74 VTAIL.n5 VTAIL.t1 1.80433
R75 VTAIL.n5 VTAIL.t4 1.80433
R76 VTAIL.n9 VTAIL.n7 1.38412
R77 VTAIL.n2 VTAIL.n1 1.38412
R78 VTAIL VTAIL.n11 1.313
R79 VTAIL VTAIL.n1 0.515586
R80 VDD1 VDD1.t2 74.7986
R81 VDD1.n1 VDD1.t5 74.6848
R82 VDD1.n1 VDD1.n0 71.9671
R83 VDD1.n3 VDD1.n2 71.5656
R84 VDD1.n3 VDD1.n1 46.6862
R85 VDD1.n2 VDD1.t0 1.80433
R86 VDD1.n2 VDD1.t1 1.80433
R87 VDD1.n0 VDD1.t4 1.80433
R88 VDD1.n0 VDD1.t3 1.80433
R89 VDD1 VDD1.n3 0.399207
R90 B.n548 B.n547 585
R91 B.n549 B.n86 585
R92 B.n551 B.n550 585
R93 B.n552 B.n85 585
R94 B.n554 B.n553 585
R95 B.n555 B.n84 585
R96 B.n557 B.n556 585
R97 B.n558 B.n83 585
R98 B.n560 B.n559 585
R99 B.n561 B.n82 585
R100 B.n563 B.n562 585
R101 B.n564 B.n81 585
R102 B.n566 B.n565 585
R103 B.n567 B.n80 585
R104 B.n569 B.n568 585
R105 B.n570 B.n79 585
R106 B.n572 B.n571 585
R107 B.n573 B.n78 585
R108 B.n575 B.n574 585
R109 B.n576 B.n77 585
R110 B.n578 B.n577 585
R111 B.n579 B.n76 585
R112 B.n581 B.n580 585
R113 B.n582 B.n75 585
R114 B.n584 B.n583 585
R115 B.n585 B.n74 585
R116 B.n587 B.n586 585
R117 B.n588 B.n73 585
R118 B.n590 B.n589 585
R119 B.n591 B.n72 585
R120 B.n593 B.n592 585
R121 B.n594 B.n71 585
R122 B.n596 B.n595 585
R123 B.n597 B.n70 585
R124 B.n599 B.n598 585
R125 B.n600 B.n69 585
R126 B.n602 B.n601 585
R127 B.n603 B.n68 585
R128 B.n605 B.n604 585
R129 B.n606 B.n67 585
R130 B.n608 B.n607 585
R131 B.n609 B.n66 585
R132 B.n611 B.n610 585
R133 B.n612 B.n65 585
R134 B.n614 B.n613 585
R135 B.n615 B.n64 585
R136 B.n617 B.n616 585
R137 B.n618 B.n63 585
R138 B.n620 B.n619 585
R139 B.n621 B.n62 585
R140 B.n623 B.n622 585
R141 B.n624 B.n61 585
R142 B.n626 B.n625 585
R143 B.n627 B.n60 585
R144 B.n629 B.n628 585
R145 B.n630 B.n59 585
R146 B.n632 B.n631 585
R147 B.n633 B.n58 585
R148 B.n635 B.n634 585
R149 B.n637 B.n55 585
R150 B.n639 B.n638 585
R151 B.n640 B.n54 585
R152 B.n642 B.n641 585
R153 B.n643 B.n53 585
R154 B.n645 B.n644 585
R155 B.n646 B.n52 585
R156 B.n648 B.n647 585
R157 B.n649 B.n51 585
R158 B.n651 B.n650 585
R159 B.n653 B.n652 585
R160 B.n654 B.n47 585
R161 B.n656 B.n655 585
R162 B.n657 B.n46 585
R163 B.n659 B.n658 585
R164 B.n660 B.n45 585
R165 B.n662 B.n661 585
R166 B.n663 B.n44 585
R167 B.n665 B.n664 585
R168 B.n666 B.n43 585
R169 B.n668 B.n667 585
R170 B.n669 B.n42 585
R171 B.n671 B.n670 585
R172 B.n672 B.n41 585
R173 B.n674 B.n673 585
R174 B.n675 B.n40 585
R175 B.n677 B.n676 585
R176 B.n678 B.n39 585
R177 B.n680 B.n679 585
R178 B.n681 B.n38 585
R179 B.n683 B.n682 585
R180 B.n684 B.n37 585
R181 B.n686 B.n685 585
R182 B.n687 B.n36 585
R183 B.n689 B.n688 585
R184 B.n690 B.n35 585
R185 B.n692 B.n691 585
R186 B.n693 B.n34 585
R187 B.n695 B.n694 585
R188 B.n696 B.n33 585
R189 B.n698 B.n697 585
R190 B.n699 B.n32 585
R191 B.n701 B.n700 585
R192 B.n702 B.n31 585
R193 B.n704 B.n703 585
R194 B.n705 B.n30 585
R195 B.n707 B.n706 585
R196 B.n708 B.n29 585
R197 B.n710 B.n709 585
R198 B.n711 B.n28 585
R199 B.n713 B.n712 585
R200 B.n714 B.n27 585
R201 B.n716 B.n715 585
R202 B.n717 B.n26 585
R203 B.n719 B.n718 585
R204 B.n720 B.n25 585
R205 B.n722 B.n721 585
R206 B.n723 B.n24 585
R207 B.n725 B.n724 585
R208 B.n726 B.n23 585
R209 B.n728 B.n727 585
R210 B.n729 B.n22 585
R211 B.n731 B.n730 585
R212 B.n732 B.n21 585
R213 B.n734 B.n733 585
R214 B.n735 B.n20 585
R215 B.n737 B.n736 585
R216 B.n738 B.n19 585
R217 B.n740 B.n739 585
R218 B.n546 B.n87 585
R219 B.n545 B.n544 585
R220 B.n543 B.n88 585
R221 B.n542 B.n541 585
R222 B.n540 B.n89 585
R223 B.n539 B.n538 585
R224 B.n537 B.n90 585
R225 B.n536 B.n535 585
R226 B.n534 B.n91 585
R227 B.n533 B.n532 585
R228 B.n531 B.n92 585
R229 B.n530 B.n529 585
R230 B.n528 B.n93 585
R231 B.n527 B.n526 585
R232 B.n525 B.n94 585
R233 B.n524 B.n523 585
R234 B.n522 B.n95 585
R235 B.n521 B.n520 585
R236 B.n519 B.n96 585
R237 B.n518 B.n517 585
R238 B.n516 B.n97 585
R239 B.n515 B.n514 585
R240 B.n513 B.n98 585
R241 B.n512 B.n511 585
R242 B.n510 B.n99 585
R243 B.n509 B.n508 585
R244 B.n507 B.n100 585
R245 B.n506 B.n505 585
R246 B.n504 B.n101 585
R247 B.n503 B.n502 585
R248 B.n501 B.n102 585
R249 B.n500 B.n499 585
R250 B.n498 B.n103 585
R251 B.n497 B.n496 585
R252 B.n495 B.n104 585
R253 B.n494 B.n493 585
R254 B.n492 B.n105 585
R255 B.n491 B.n490 585
R256 B.n489 B.n106 585
R257 B.n488 B.n487 585
R258 B.n486 B.n107 585
R259 B.n485 B.n484 585
R260 B.n483 B.n108 585
R261 B.n482 B.n481 585
R262 B.n480 B.n109 585
R263 B.n479 B.n478 585
R264 B.n477 B.n110 585
R265 B.n476 B.n475 585
R266 B.n474 B.n111 585
R267 B.n473 B.n472 585
R268 B.n471 B.n112 585
R269 B.n470 B.n469 585
R270 B.n468 B.n113 585
R271 B.n467 B.n466 585
R272 B.n465 B.n114 585
R273 B.n464 B.n463 585
R274 B.n462 B.n115 585
R275 B.n461 B.n460 585
R276 B.n459 B.n116 585
R277 B.n458 B.n457 585
R278 B.n456 B.n117 585
R279 B.n455 B.n454 585
R280 B.n453 B.n118 585
R281 B.n452 B.n451 585
R282 B.n450 B.n119 585
R283 B.n449 B.n448 585
R284 B.n447 B.n120 585
R285 B.n254 B.n253 585
R286 B.n255 B.n188 585
R287 B.n257 B.n256 585
R288 B.n258 B.n187 585
R289 B.n260 B.n259 585
R290 B.n261 B.n186 585
R291 B.n263 B.n262 585
R292 B.n264 B.n185 585
R293 B.n266 B.n265 585
R294 B.n267 B.n184 585
R295 B.n269 B.n268 585
R296 B.n270 B.n183 585
R297 B.n272 B.n271 585
R298 B.n273 B.n182 585
R299 B.n275 B.n274 585
R300 B.n276 B.n181 585
R301 B.n278 B.n277 585
R302 B.n279 B.n180 585
R303 B.n281 B.n280 585
R304 B.n282 B.n179 585
R305 B.n284 B.n283 585
R306 B.n285 B.n178 585
R307 B.n287 B.n286 585
R308 B.n288 B.n177 585
R309 B.n290 B.n289 585
R310 B.n291 B.n176 585
R311 B.n293 B.n292 585
R312 B.n294 B.n175 585
R313 B.n296 B.n295 585
R314 B.n297 B.n174 585
R315 B.n299 B.n298 585
R316 B.n300 B.n173 585
R317 B.n302 B.n301 585
R318 B.n303 B.n172 585
R319 B.n305 B.n304 585
R320 B.n306 B.n171 585
R321 B.n308 B.n307 585
R322 B.n309 B.n170 585
R323 B.n311 B.n310 585
R324 B.n312 B.n169 585
R325 B.n314 B.n313 585
R326 B.n315 B.n168 585
R327 B.n317 B.n316 585
R328 B.n318 B.n167 585
R329 B.n320 B.n319 585
R330 B.n321 B.n166 585
R331 B.n323 B.n322 585
R332 B.n324 B.n165 585
R333 B.n326 B.n325 585
R334 B.n327 B.n164 585
R335 B.n329 B.n328 585
R336 B.n330 B.n163 585
R337 B.n332 B.n331 585
R338 B.n333 B.n162 585
R339 B.n335 B.n334 585
R340 B.n336 B.n161 585
R341 B.n338 B.n337 585
R342 B.n339 B.n160 585
R343 B.n341 B.n340 585
R344 B.n343 B.n157 585
R345 B.n345 B.n344 585
R346 B.n346 B.n156 585
R347 B.n348 B.n347 585
R348 B.n349 B.n155 585
R349 B.n351 B.n350 585
R350 B.n352 B.n154 585
R351 B.n354 B.n353 585
R352 B.n355 B.n153 585
R353 B.n357 B.n356 585
R354 B.n359 B.n358 585
R355 B.n360 B.n149 585
R356 B.n362 B.n361 585
R357 B.n363 B.n148 585
R358 B.n365 B.n364 585
R359 B.n366 B.n147 585
R360 B.n368 B.n367 585
R361 B.n369 B.n146 585
R362 B.n371 B.n370 585
R363 B.n372 B.n145 585
R364 B.n374 B.n373 585
R365 B.n375 B.n144 585
R366 B.n377 B.n376 585
R367 B.n378 B.n143 585
R368 B.n380 B.n379 585
R369 B.n381 B.n142 585
R370 B.n383 B.n382 585
R371 B.n384 B.n141 585
R372 B.n386 B.n385 585
R373 B.n387 B.n140 585
R374 B.n389 B.n388 585
R375 B.n390 B.n139 585
R376 B.n392 B.n391 585
R377 B.n393 B.n138 585
R378 B.n395 B.n394 585
R379 B.n396 B.n137 585
R380 B.n398 B.n397 585
R381 B.n399 B.n136 585
R382 B.n401 B.n400 585
R383 B.n402 B.n135 585
R384 B.n404 B.n403 585
R385 B.n405 B.n134 585
R386 B.n407 B.n406 585
R387 B.n408 B.n133 585
R388 B.n410 B.n409 585
R389 B.n411 B.n132 585
R390 B.n413 B.n412 585
R391 B.n414 B.n131 585
R392 B.n416 B.n415 585
R393 B.n417 B.n130 585
R394 B.n419 B.n418 585
R395 B.n420 B.n129 585
R396 B.n422 B.n421 585
R397 B.n423 B.n128 585
R398 B.n425 B.n424 585
R399 B.n426 B.n127 585
R400 B.n428 B.n427 585
R401 B.n429 B.n126 585
R402 B.n431 B.n430 585
R403 B.n432 B.n125 585
R404 B.n434 B.n433 585
R405 B.n435 B.n124 585
R406 B.n437 B.n436 585
R407 B.n438 B.n123 585
R408 B.n440 B.n439 585
R409 B.n441 B.n122 585
R410 B.n443 B.n442 585
R411 B.n444 B.n121 585
R412 B.n446 B.n445 585
R413 B.n252 B.n189 585
R414 B.n251 B.n250 585
R415 B.n249 B.n190 585
R416 B.n248 B.n247 585
R417 B.n246 B.n191 585
R418 B.n245 B.n244 585
R419 B.n243 B.n192 585
R420 B.n242 B.n241 585
R421 B.n240 B.n193 585
R422 B.n239 B.n238 585
R423 B.n237 B.n194 585
R424 B.n236 B.n235 585
R425 B.n234 B.n195 585
R426 B.n233 B.n232 585
R427 B.n231 B.n196 585
R428 B.n230 B.n229 585
R429 B.n228 B.n197 585
R430 B.n227 B.n226 585
R431 B.n225 B.n198 585
R432 B.n224 B.n223 585
R433 B.n222 B.n199 585
R434 B.n221 B.n220 585
R435 B.n219 B.n200 585
R436 B.n218 B.n217 585
R437 B.n216 B.n201 585
R438 B.n215 B.n214 585
R439 B.n213 B.n202 585
R440 B.n212 B.n211 585
R441 B.n210 B.n203 585
R442 B.n209 B.n208 585
R443 B.n207 B.n204 585
R444 B.n206 B.n205 585
R445 B.n2 B.n0 585
R446 B.n789 B.n1 585
R447 B.n788 B.n787 585
R448 B.n786 B.n3 585
R449 B.n785 B.n784 585
R450 B.n783 B.n4 585
R451 B.n782 B.n781 585
R452 B.n780 B.n5 585
R453 B.n779 B.n778 585
R454 B.n777 B.n6 585
R455 B.n776 B.n775 585
R456 B.n774 B.n7 585
R457 B.n773 B.n772 585
R458 B.n771 B.n8 585
R459 B.n770 B.n769 585
R460 B.n768 B.n9 585
R461 B.n767 B.n766 585
R462 B.n765 B.n10 585
R463 B.n764 B.n763 585
R464 B.n762 B.n11 585
R465 B.n761 B.n760 585
R466 B.n759 B.n12 585
R467 B.n758 B.n757 585
R468 B.n756 B.n13 585
R469 B.n755 B.n754 585
R470 B.n753 B.n14 585
R471 B.n752 B.n751 585
R472 B.n750 B.n15 585
R473 B.n749 B.n748 585
R474 B.n747 B.n16 585
R475 B.n746 B.n745 585
R476 B.n744 B.n17 585
R477 B.n743 B.n742 585
R478 B.n741 B.n18 585
R479 B.n791 B.n790 585
R480 B.n254 B.n189 526.135
R481 B.n741 B.n740 526.135
R482 B.n447 B.n446 526.135
R483 B.n548 B.n87 526.135
R484 B.n150 B.t9 448.995
R485 B.n158 B.t3 448.995
R486 B.n48 B.t6 448.995
R487 B.n56 B.t0 448.995
R488 B.n250 B.n189 163.367
R489 B.n250 B.n249 163.367
R490 B.n249 B.n248 163.367
R491 B.n248 B.n191 163.367
R492 B.n244 B.n191 163.367
R493 B.n244 B.n243 163.367
R494 B.n243 B.n242 163.367
R495 B.n242 B.n193 163.367
R496 B.n238 B.n193 163.367
R497 B.n238 B.n237 163.367
R498 B.n237 B.n236 163.367
R499 B.n236 B.n195 163.367
R500 B.n232 B.n195 163.367
R501 B.n232 B.n231 163.367
R502 B.n231 B.n230 163.367
R503 B.n230 B.n197 163.367
R504 B.n226 B.n197 163.367
R505 B.n226 B.n225 163.367
R506 B.n225 B.n224 163.367
R507 B.n224 B.n199 163.367
R508 B.n220 B.n199 163.367
R509 B.n220 B.n219 163.367
R510 B.n219 B.n218 163.367
R511 B.n218 B.n201 163.367
R512 B.n214 B.n201 163.367
R513 B.n214 B.n213 163.367
R514 B.n213 B.n212 163.367
R515 B.n212 B.n203 163.367
R516 B.n208 B.n203 163.367
R517 B.n208 B.n207 163.367
R518 B.n207 B.n206 163.367
R519 B.n206 B.n2 163.367
R520 B.n790 B.n2 163.367
R521 B.n790 B.n789 163.367
R522 B.n789 B.n788 163.367
R523 B.n788 B.n3 163.367
R524 B.n784 B.n3 163.367
R525 B.n784 B.n783 163.367
R526 B.n783 B.n782 163.367
R527 B.n782 B.n5 163.367
R528 B.n778 B.n5 163.367
R529 B.n778 B.n777 163.367
R530 B.n777 B.n776 163.367
R531 B.n776 B.n7 163.367
R532 B.n772 B.n7 163.367
R533 B.n772 B.n771 163.367
R534 B.n771 B.n770 163.367
R535 B.n770 B.n9 163.367
R536 B.n766 B.n9 163.367
R537 B.n766 B.n765 163.367
R538 B.n765 B.n764 163.367
R539 B.n764 B.n11 163.367
R540 B.n760 B.n11 163.367
R541 B.n760 B.n759 163.367
R542 B.n759 B.n758 163.367
R543 B.n758 B.n13 163.367
R544 B.n754 B.n13 163.367
R545 B.n754 B.n753 163.367
R546 B.n753 B.n752 163.367
R547 B.n752 B.n15 163.367
R548 B.n748 B.n15 163.367
R549 B.n748 B.n747 163.367
R550 B.n747 B.n746 163.367
R551 B.n746 B.n17 163.367
R552 B.n742 B.n17 163.367
R553 B.n742 B.n741 163.367
R554 B.n255 B.n254 163.367
R555 B.n256 B.n255 163.367
R556 B.n256 B.n187 163.367
R557 B.n260 B.n187 163.367
R558 B.n261 B.n260 163.367
R559 B.n262 B.n261 163.367
R560 B.n262 B.n185 163.367
R561 B.n266 B.n185 163.367
R562 B.n267 B.n266 163.367
R563 B.n268 B.n267 163.367
R564 B.n268 B.n183 163.367
R565 B.n272 B.n183 163.367
R566 B.n273 B.n272 163.367
R567 B.n274 B.n273 163.367
R568 B.n274 B.n181 163.367
R569 B.n278 B.n181 163.367
R570 B.n279 B.n278 163.367
R571 B.n280 B.n279 163.367
R572 B.n280 B.n179 163.367
R573 B.n284 B.n179 163.367
R574 B.n285 B.n284 163.367
R575 B.n286 B.n285 163.367
R576 B.n286 B.n177 163.367
R577 B.n290 B.n177 163.367
R578 B.n291 B.n290 163.367
R579 B.n292 B.n291 163.367
R580 B.n292 B.n175 163.367
R581 B.n296 B.n175 163.367
R582 B.n297 B.n296 163.367
R583 B.n298 B.n297 163.367
R584 B.n298 B.n173 163.367
R585 B.n302 B.n173 163.367
R586 B.n303 B.n302 163.367
R587 B.n304 B.n303 163.367
R588 B.n304 B.n171 163.367
R589 B.n308 B.n171 163.367
R590 B.n309 B.n308 163.367
R591 B.n310 B.n309 163.367
R592 B.n310 B.n169 163.367
R593 B.n314 B.n169 163.367
R594 B.n315 B.n314 163.367
R595 B.n316 B.n315 163.367
R596 B.n316 B.n167 163.367
R597 B.n320 B.n167 163.367
R598 B.n321 B.n320 163.367
R599 B.n322 B.n321 163.367
R600 B.n322 B.n165 163.367
R601 B.n326 B.n165 163.367
R602 B.n327 B.n326 163.367
R603 B.n328 B.n327 163.367
R604 B.n328 B.n163 163.367
R605 B.n332 B.n163 163.367
R606 B.n333 B.n332 163.367
R607 B.n334 B.n333 163.367
R608 B.n334 B.n161 163.367
R609 B.n338 B.n161 163.367
R610 B.n339 B.n338 163.367
R611 B.n340 B.n339 163.367
R612 B.n340 B.n157 163.367
R613 B.n345 B.n157 163.367
R614 B.n346 B.n345 163.367
R615 B.n347 B.n346 163.367
R616 B.n347 B.n155 163.367
R617 B.n351 B.n155 163.367
R618 B.n352 B.n351 163.367
R619 B.n353 B.n352 163.367
R620 B.n353 B.n153 163.367
R621 B.n357 B.n153 163.367
R622 B.n358 B.n357 163.367
R623 B.n358 B.n149 163.367
R624 B.n362 B.n149 163.367
R625 B.n363 B.n362 163.367
R626 B.n364 B.n363 163.367
R627 B.n364 B.n147 163.367
R628 B.n368 B.n147 163.367
R629 B.n369 B.n368 163.367
R630 B.n370 B.n369 163.367
R631 B.n370 B.n145 163.367
R632 B.n374 B.n145 163.367
R633 B.n375 B.n374 163.367
R634 B.n376 B.n375 163.367
R635 B.n376 B.n143 163.367
R636 B.n380 B.n143 163.367
R637 B.n381 B.n380 163.367
R638 B.n382 B.n381 163.367
R639 B.n382 B.n141 163.367
R640 B.n386 B.n141 163.367
R641 B.n387 B.n386 163.367
R642 B.n388 B.n387 163.367
R643 B.n388 B.n139 163.367
R644 B.n392 B.n139 163.367
R645 B.n393 B.n392 163.367
R646 B.n394 B.n393 163.367
R647 B.n394 B.n137 163.367
R648 B.n398 B.n137 163.367
R649 B.n399 B.n398 163.367
R650 B.n400 B.n399 163.367
R651 B.n400 B.n135 163.367
R652 B.n404 B.n135 163.367
R653 B.n405 B.n404 163.367
R654 B.n406 B.n405 163.367
R655 B.n406 B.n133 163.367
R656 B.n410 B.n133 163.367
R657 B.n411 B.n410 163.367
R658 B.n412 B.n411 163.367
R659 B.n412 B.n131 163.367
R660 B.n416 B.n131 163.367
R661 B.n417 B.n416 163.367
R662 B.n418 B.n417 163.367
R663 B.n418 B.n129 163.367
R664 B.n422 B.n129 163.367
R665 B.n423 B.n422 163.367
R666 B.n424 B.n423 163.367
R667 B.n424 B.n127 163.367
R668 B.n428 B.n127 163.367
R669 B.n429 B.n428 163.367
R670 B.n430 B.n429 163.367
R671 B.n430 B.n125 163.367
R672 B.n434 B.n125 163.367
R673 B.n435 B.n434 163.367
R674 B.n436 B.n435 163.367
R675 B.n436 B.n123 163.367
R676 B.n440 B.n123 163.367
R677 B.n441 B.n440 163.367
R678 B.n442 B.n441 163.367
R679 B.n442 B.n121 163.367
R680 B.n446 B.n121 163.367
R681 B.n448 B.n447 163.367
R682 B.n448 B.n119 163.367
R683 B.n452 B.n119 163.367
R684 B.n453 B.n452 163.367
R685 B.n454 B.n453 163.367
R686 B.n454 B.n117 163.367
R687 B.n458 B.n117 163.367
R688 B.n459 B.n458 163.367
R689 B.n460 B.n459 163.367
R690 B.n460 B.n115 163.367
R691 B.n464 B.n115 163.367
R692 B.n465 B.n464 163.367
R693 B.n466 B.n465 163.367
R694 B.n466 B.n113 163.367
R695 B.n470 B.n113 163.367
R696 B.n471 B.n470 163.367
R697 B.n472 B.n471 163.367
R698 B.n472 B.n111 163.367
R699 B.n476 B.n111 163.367
R700 B.n477 B.n476 163.367
R701 B.n478 B.n477 163.367
R702 B.n478 B.n109 163.367
R703 B.n482 B.n109 163.367
R704 B.n483 B.n482 163.367
R705 B.n484 B.n483 163.367
R706 B.n484 B.n107 163.367
R707 B.n488 B.n107 163.367
R708 B.n489 B.n488 163.367
R709 B.n490 B.n489 163.367
R710 B.n490 B.n105 163.367
R711 B.n494 B.n105 163.367
R712 B.n495 B.n494 163.367
R713 B.n496 B.n495 163.367
R714 B.n496 B.n103 163.367
R715 B.n500 B.n103 163.367
R716 B.n501 B.n500 163.367
R717 B.n502 B.n501 163.367
R718 B.n502 B.n101 163.367
R719 B.n506 B.n101 163.367
R720 B.n507 B.n506 163.367
R721 B.n508 B.n507 163.367
R722 B.n508 B.n99 163.367
R723 B.n512 B.n99 163.367
R724 B.n513 B.n512 163.367
R725 B.n514 B.n513 163.367
R726 B.n514 B.n97 163.367
R727 B.n518 B.n97 163.367
R728 B.n519 B.n518 163.367
R729 B.n520 B.n519 163.367
R730 B.n520 B.n95 163.367
R731 B.n524 B.n95 163.367
R732 B.n525 B.n524 163.367
R733 B.n526 B.n525 163.367
R734 B.n526 B.n93 163.367
R735 B.n530 B.n93 163.367
R736 B.n531 B.n530 163.367
R737 B.n532 B.n531 163.367
R738 B.n532 B.n91 163.367
R739 B.n536 B.n91 163.367
R740 B.n537 B.n536 163.367
R741 B.n538 B.n537 163.367
R742 B.n538 B.n89 163.367
R743 B.n542 B.n89 163.367
R744 B.n543 B.n542 163.367
R745 B.n544 B.n543 163.367
R746 B.n544 B.n87 163.367
R747 B.n740 B.n19 163.367
R748 B.n736 B.n19 163.367
R749 B.n736 B.n735 163.367
R750 B.n735 B.n734 163.367
R751 B.n734 B.n21 163.367
R752 B.n730 B.n21 163.367
R753 B.n730 B.n729 163.367
R754 B.n729 B.n728 163.367
R755 B.n728 B.n23 163.367
R756 B.n724 B.n23 163.367
R757 B.n724 B.n723 163.367
R758 B.n723 B.n722 163.367
R759 B.n722 B.n25 163.367
R760 B.n718 B.n25 163.367
R761 B.n718 B.n717 163.367
R762 B.n717 B.n716 163.367
R763 B.n716 B.n27 163.367
R764 B.n712 B.n27 163.367
R765 B.n712 B.n711 163.367
R766 B.n711 B.n710 163.367
R767 B.n710 B.n29 163.367
R768 B.n706 B.n29 163.367
R769 B.n706 B.n705 163.367
R770 B.n705 B.n704 163.367
R771 B.n704 B.n31 163.367
R772 B.n700 B.n31 163.367
R773 B.n700 B.n699 163.367
R774 B.n699 B.n698 163.367
R775 B.n698 B.n33 163.367
R776 B.n694 B.n33 163.367
R777 B.n694 B.n693 163.367
R778 B.n693 B.n692 163.367
R779 B.n692 B.n35 163.367
R780 B.n688 B.n35 163.367
R781 B.n688 B.n687 163.367
R782 B.n687 B.n686 163.367
R783 B.n686 B.n37 163.367
R784 B.n682 B.n37 163.367
R785 B.n682 B.n681 163.367
R786 B.n681 B.n680 163.367
R787 B.n680 B.n39 163.367
R788 B.n676 B.n39 163.367
R789 B.n676 B.n675 163.367
R790 B.n675 B.n674 163.367
R791 B.n674 B.n41 163.367
R792 B.n670 B.n41 163.367
R793 B.n670 B.n669 163.367
R794 B.n669 B.n668 163.367
R795 B.n668 B.n43 163.367
R796 B.n664 B.n43 163.367
R797 B.n664 B.n663 163.367
R798 B.n663 B.n662 163.367
R799 B.n662 B.n45 163.367
R800 B.n658 B.n45 163.367
R801 B.n658 B.n657 163.367
R802 B.n657 B.n656 163.367
R803 B.n656 B.n47 163.367
R804 B.n652 B.n47 163.367
R805 B.n652 B.n651 163.367
R806 B.n651 B.n51 163.367
R807 B.n647 B.n51 163.367
R808 B.n647 B.n646 163.367
R809 B.n646 B.n645 163.367
R810 B.n645 B.n53 163.367
R811 B.n641 B.n53 163.367
R812 B.n641 B.n640 163.367
R813 B.n640 B.n639 163.367
R814 B.n639 B.n55 163.367
R815 B.n634 B.n55 163.367
R816 B.n634 B.n633 163.367
R817 B.n633 B.n632 163.367
R818 B.n632 B.n59 163.367
R819 B.n628 B.n59 163.367
R820 B.n628 B.n627 163.367
R821 B.n627 B.n626 163.367
R822 B.n626 B.n61 163.367
R823 B.n622 B.n61 163.367
R824 B.n622 B.n621 163.367
R825 B.n621 B.n620 163.367
R826 B.n620 B.n63 163.367
R827 B.n616 B.n63 163.367
R828 B.n616 B.n615 163.367
R829 B.n615 B.n614 163.367
R830 B.n614 B.n65 163.367
R831 B.n610 B.n65 163.367
R832 B.n610 B.n609 163.367
R833 B.n609 B.n608 163.367
R834 B.n608 B.n67 163.367
R835 B.n604 B.n67 163.367
R836 B.n604 B.n603 163.367
R837 B.n603 B.n602 163.367
R838 B.n602 B.n69 163.367
R839 B.n598 B.n69 163.367
R840 B.n598 B.n597 163.367
R841 B.n597 B.n596 163.367
R842 B.n596 B.n71 163.367
R843 B.n592 B.n71 163.367
R844 B.n592 B.n591 163.367
R845 B.n591 B.n590 163.367
R846 B.n590 B.n73 163.367
R847 B.n586 B.n73 163.367
R848 B.n586 B.n585 163.367
R849 B.n585 B.n584 163.367
R850 B.n584 B.n75 163.367
R851 B.n580 B.n75 163.367
R852 B.n580 B.n579 163.367
R853 B.n579 B.n578 163.367
R854 B.n578 B.n77 163.367
R855 B.n574 B.n77 163.367
R856 B.n574 B.n573 163.367
R857 B.n573 B.n572 163.367
R858 B.n572 B.n79 163.367
R859 B.n568 B.n79 163.367
R860 B.n568 B.n567 163.367
R861 B.n567 B.n566 163.367
R862 B.n566 B.n81 163.367
R863 B.n562 B.n81 163.367
R864 B.n562 B.n561 163.367
R865 B.n561 B.n560 163.367
R866 B.n560 B.n83 163.367
R867 B.n556 B.n83 163.367
R868 B.n556 B.n555 163.367
R869 B.n555 B.n554 163.367
R870 B.n554 B.n85 163.367
R871 B.n550 B.n85 163.367
R872 B.n550 B.n549 163.367
R873 B.n549 B.n548 163.367
R874 B.n150 B.t11 153.911
R875 B.n56 B.t1 153.911
R876 B.n158 B.t5 153.887
R877 B.n48 B.t7 153.887
R878 B.n151 B.t10 112.796
R879 B.n57 B.t2 112.796
R880 B.n159 B.t4 112.772
R881 B.n49 B.t8 112.772
R882 B.n152 B.n151 59.5399
R883 B.n342 B.n159 59.5399
R884 B.n50 B.n49 59.5399
R885 B.n636 B.n57 59.5399
R886 B.n151 B.n150 41.1157
R887 B.n159 B.n158 41.1157
R888 B.n49 B.n48 41.1157
R889 B.n57 B.n56 41.1157
R890 B.n739 B.n18 34.1859
R891 B.n547 B.n546 34.1859
R892 B.n445 B.n120 34.1859
R893 B.n253 B.n252 34.1859
R894 B B.n791 18.0485
R895 B.n739 B.n738 10.6151
R896 B.n738 B.n737 10.6151
R897 B.n737 B.n20 10.6151
R898 B.n733 B.n20 10.6151
R899 B.n733 B.n732 10.6151
R900 B.n732 B.n731 10.6151
R901 B.n731 B.n22 10.6151
R902 B.n727 B.n22 10.6151
R903 B.n727 B.n726 10.6151
R904 B.n726 B.n725 10.6151
R905 B.n725 B.n24 10.6151
R906 B.n721 B.n24 10.6151
R907 B.n721 B.n720 10.6151
R908 B.n720 B.n719 10.6151
R909 B.n719 B.n26 10.6151
R910 B.n715 B.n26 10.6151
R911 B.n715 B.n714 10.6151
R912 B.n714 B.n713 10.6151
R913 B.n713 B.n28 10.6151
R914 B.n709 B.n28 10.6151
R915 B.n709 B.n708 10.6151
R916 B.n708 B.n707 10.6151
R917 B.n707 B.n30 10.6151
R918 B.n703 B.n30 10.6151
R919 B.n703 B.n702 10.6151
R920 B.n702 B.n701 10.6151
R921 B.n701 B.n32 10.6151
R922 B.n697 B.n32 10.6151
R923 B.n697 B.n696 10.6151
R924 B.n696 B.n695 10.6151
R925 B.n695 B.n34 10.6151
R926 B.n691 B.n34 10.6151
R927 B.n691 B.n690 10.6151
R928 B.n690 B.n689 10.6151
R929 B.n689 B.n36 10.6151
R930 B.n685 B.n36 10.6151
R931 B.n685 B.n684 10.6151
R932 B.n684 B.n683 10.6151
R933 B.n683 B.n38 10.6151
R934 B.n679 B.n38 10.6151
R935 B.n679 B.n678 10.6151
R936 B.n678 B.n677 10.6151
R937 B.n677 B.n40 10.6151
R938 B.n673 B.n40 10.6151
R939 B.n673 B.n672 10.6151
R940 B.n672 B.n671 10.6151
R941 B.n671 B.n42 10.6151
R942 B.n667 B.n42 10.6151
R943 B.n667 B.n666 10.6151
R944 B.n666 B.n665 10.6151
R945 B.n665 B.n44 10.6151
R946 B.n661 B.n44 10.6151
R947 B.n661 B.n660 10.6151
R948 B.n660 B.n659 10.6151
R949 B.n659 B.n46 10.6151
R950 B.n655 B.n46 10.6151
R951 B.n655 B.n654 10.6151
R952 B.n654 B.n653 10.6151
R953 B.n650 B.n649 10.6151
R954 B.n649 B.n648 10.6151
R955 B.n648 B.n52 10.6151
R956 B.n644 B.n52 10.6151
R957 B.n644 B.n643 10.6151
R958 B.n643 B.n642 10.6151
R959 B.n642 B.n54 10.6151
R960 B.n638 B.n54 10.6151
R961 B.n638 B.n637 10.6151
R962 B.n635 B.n58 10.6151
R963 B.n631 B.n58 10.6151
R964 B.n631 B.n630 10.6151
R965 B.n630 B.n629 10.6151
R966 B.n629 B.n60 10.6151
R967 B.n625 B.n60 10.6151
R968 B.n625 B.n624 10.6151
R969 B.n624 B.n623 10.6151
R970 B.n623 B.n62 10.6151
R971 B.n619 B.n62 10.6151
R972 B.n619 B.n618 10.6151
R973 B.n618 B.n617 10.6151
R974 B.n617 B.n64 10.6151
R975 B.n613 B.n64 10.6151
R976 B.n613 B.n612 10.6151
R977 B.n612 B.n611 10.6151
R978 B.n611 B.n66 10.6151
R979 B.n607 B.n66 10.6151
R980 B.n607 B.n606 10.6151
R981 B.n606 B.n605 10.6151
R982 B.n605 B.n68 10.6151
R983 B.n601 B.n68 10.6151
R984 B.n601 B.n600 10.6151
R985 B.n600 B.n599 10.6151
R986 B.n599 B.n70 10.6151
R987 B.n595 B.n70 10.6151
R988 B.n595 B.n594 10.6151
R989 B.n594 B.n593 10.6151
R990 B.n593 B.n72 10.6151
R991 B.n589 B.n72 10.6151
R992 B.n589 B.n588 10.6151
R993 B.n588 B.n587 10.6151
R994 B.n587 B.n74 10.6151
R995 B.n583 B.n74 10.6151
R996 B.n583 B.n582 10.6151
R997 B.n582 B.n581 10.6151
R998 B.n581 B.n76 10.6151
R999 B.n577 B.n76 10.6151
R1000 B.n577 B.n576 10.6151
R1001 B.n576 B.n575 10.6151
R1002 B.n575 B.n78 10.6151
R1003 B.n571 B.n78 10.6151
R1004 B.n571 B.n570 10.6151
R1005 B.n570 B.n569 10.6151
R1006 B.n569 B.n80 10.6151
R1007 B.n565 B.n80 10.6151
R1008 B.n565 B.n564 10.6151
R1009 B.n564 B.n563 10.6151
R1010 B.n563 B.n82 10.6151
R1011 B.n559 B.n82 10.6151
R1012 B.n559 B.n558 10.6151
R1013 B.n558 B.n557 10.6151
R1014 B.n557 B.n84 10.6151
R1015 B.n553 B.n84 10.6151
R1016 B.n553 B.n552 10.6151
R1017 B.n552 B.n551 10.6151
R1018 B.n551 B.n86 10.6151
R1019 B.n547 B.n86 10.6151
R1020 B.n449 B.n120 10.6151
R1021 B.n450 B.n449 10.6151
R1022 B.n451 B.n450 10.6151
R1023 B.n451 B.n118 10.6151
R1024 B.n455 B.n118 10.6151
R1025 B.n456 B.n455 10.6151
R1026 B.n457 B.n456 10.6151
R1027 B.n457 B.n116 10.6151
R1028 B.n461 B.n116 10.6151
R1029 B.n462 B.n461 10.6151
R1030 B.n463 B.n462 10.6151
R1031 B.n463 B.n114 10.6151
R1032 B.n467 B.n114 10.6151
R1033 B.n468 B.n467 10.6151
R1034 B.n469 B.n468 10.6151
R1035 B.n469 B.n112 10.6151
R1036 B.n473 B.n112 10.6151
R1037 B.n474 B.n473 10.6151
R1038 B.n475 B.n474 10.6151
R1039 B.n475 B.n110 10.6151
R1040 B.n479 B.n110 10.6151
R1041 B.n480 B.n479 10.6151
R1042 B.n481 B.n480 10.6151
R1043 B.n481 B.n108 10.6151
R1044 B.n485 B.n108 10.6151
R1045 B.n486 B.n485 10.6151
R1046 B.n487 B.n486 10.6151
R1047 B.n487 B.n106 10.6151
R1048 B.n491 B.n106 10.6151
R1049 B.n492 B.n491 10.6151
R1050 B.n493 B.n492 10.6151
R1051 B.n493 B.n104 10.6151
R1052 B.n497 B.n104 10.6151
R1053 B.n498 B.n497 10.6151
R1054 B.n499 B.n498 10.6151
R1055 B.n499 B.n102 10.6151
R1056 B.n503 B.n102 10.6151
R1057 B.n504 B.n503 10.6151
R1058 B.n505 B.n504 10.6151
R1059 B.n505 B.n100 10.6151
R1060 B.n509 B.n100 10.6151
R1061 B.n510 B.n509 10.6151
R1062 B.n511 B.n510 10.6151
R1063 B.n511 B.n98 10.6151
R1064 B.n515 B.n98 10.6151
R1065 B.n516 B.n515 10.6151
R1066 B.n517 B.n516 10.6151
R1067 B.n517 B.n96 10.6151
R1068 B.n521 B.n96 10.6151
R1069 B.n522 B.n521 10.6151
R1070 B.n523 B.n522 10.6151
R1071 B.n523 B.n94 10.6151
R1072 B.n527 B.n94 10.6151
R1073 B.n528 B.n527 10.6151
R1074 B.n529 B.n528 10.6151
R1075 B.n529 B.n92 10.6151
R1076 B.n533 B.n92 10.6151
R1077 B.n534 B.n533 10.6151
R1078 B.n535 B.n534 10.6151
R1079 B.n535 B.n90 10.6151
R1080 B.n539 B.n90 10.6151
R1081 B.n540 B.n539 10.6151
R1082 B.n541 B.n540 10.6151
R1083 B.n541 B.n88 10.6151
R1084 B.n545 B.n88 10.6151
R1085 B.n546 B.n545 10.6151
R1086 B.n253 B.n188 10.6151
R1087 B.n257 B.n188 10.6151
R1088 B.n258 B.n257 10.6151
R1089 B.n259 B.n258 10.6151
R1090 B.n259 B.n186 10.6151
R1091 B.n263 B.n186 10.6151
R1092 B.n264 B.n263 10.6151
R1093 B.n265 B.n264 10.6151
R1094 B.n265 B.n184 10.6151
R1095 B.n269 B.n184 10.6151
R1096 B.n270 B.n269 10.6151
R1097 B.n271 B.n270 10.6151
R1098 B.n271 B.n182 10.6151
R1099 B.n275 B.n182 10.6151
R1100 B.n276 B.n275 10.6151
R1101 B.n277 B.n276 10.6151
R1102 B.n277 B.n180 10.6151
R1103 B.n281 B.n180 10.6151
R1104 B.n282 B.n281 10.6151
R1105 B.n283 B.n282 10.6151
R1106 B.n283 B.n178 10.6151
R1107 B.n287 B.n178 10.6151
R1108 B.n288 B.n287 10.6151
R1109 B.n289 B.n288 10.6151
R1110 B.n289 B.n176 10.6151
R1111 B.n293 B.n176 10.6151
R1112 B.n294 B.n293 10.6151
R1113 B.n295 B.n294 10.6151
R1114 B.n295 B.n174 10.6151
R1115 B.n299 B.n174 10.6151
R1116 B.n300 B.n299 10.6151
R1117 B.n301 B.n300 10.6151
R1118 B.n301 B.n172 10.6151
R1119 B.n305 B.n172 10.6151
R1120 B.n306 B.n305 10.6151
R1121 B.n307 B.n306 10.6151
R1122 B.n307 B.n170 10.6151
R1123 B.n311 B.n170 10.6151
R1124 B.n312 B.n311 10.6151
R1125 B.n313 B.n312 10.6151
R1126 B.n313 B.n168 10.6151
R1127 B.n317 B.n168 10.6151
R1128 B.n318 B.n317 10.6151
R1129 B.n319 B.n318 10.6151
R1130 B.n319 B.n166 10.6151
R1131 B.n323 B.n166 10.6151
R1132 B.n324 B.n323 10.6151
R1133 B.n325 B.n324 10.6151
R1134 B.n325 B.n164 10.6151
R1135 B.n329 B.n164 10.6151
R1136 B.n330 B.n329 10.6151
R1137 B.n331 B.n330 10.6151
R1138 B.n331 B.n162 10.6151
R1139 B.n335 B.n162 10.6151
R1140 B.n336 B.n335 10.6151
R1141 B.n337 B.n336 10.6151
R1142 B.n337 B.n160 10.6151
R1143 B.n341 B.n160 10.6151
R1144 B.n344 B.n343 10.6151
R1145 B.n344 B.n156 10.6151
R1146 B.n348 B.n156 10.6151
R1147 B.n349 B.n348 10.6151
R1148 B.n350 B.n349 10.6151
R1149 B.n350 B.n154 10.6151
R1150 B.n354 B.n154 10.6151
R1151 B.n355 B.n354 10.6151
R1152 B.n356 B.n355 10.6151
R1153 B.n360 B.n359 10.6151
R1154 B.n361 B.n360 10.6151
R1155 B.n361 B.n148 10.6151
R1156 B.n365 B.n148 10.6151
R1157 B.n366 B.n365 10.6151
R1158 B.n367 B.n366 10.6151
R1159 B.n367 B.n146 10.6151
R1160 B.n371 B.n146 10.6151
R1161 B.n372 B.n371 10.6151
R1162 B.n373 B.n372 10.6151
R1163 B.n373 B.n144 10.6151
R1164 B.n377 B.n144 10.6151
R1165 B.n378 B.n377 10.6151
R1166 B.n379 B.n378 10.6151
R1167 B.n379 B.n142 10.6151
R1168 B.n383 B.n142 10.6151
R1169 B.n384 B.n383 10.6151
R1170 B.n385 B.n384 10.6151
R1171 B.n385 B.n140 10.6151
R1172 B.n389 B.n140 10.6151
R1173 B.n390 B.n389 10.6151
R1174 B.n391 B.n390 10.6151
R1175 B.n391 B.n138 10.6151
R1176 B.n395 B.n138 10.6151
R1177 B.n396 B.n395 10.6151
R1178 B.n397 B.n396 10.6151
R1179 B.n397 B.n136 10.6151
R1180 B.n401 B.n136 10.6151
R1181 B.n402 B.n401 10.6151
R1182 B.n403 B.n402 10.6151
R1183 B.n403 B.n134 10.6151
R1184 B.n407 B.n134 10.6151
R1185 B.n408 B.n407 10.6151
R1186 B.n409 B.n408 10.6151
R1187 B.n409 B.n132 10.6151
R1188 B.n413 B.n132 10.6151
R1189 B.n414 B.n413 10.6151
R1190 B.n415 B.n414 10.6151
R1191 B.n415 B.n130 10.6151
R1192 B.n419 B.n130 10.6151
R1193 B.n420 B.n419 10.6151
R1194 B.n421 B.n420 10.6151
R1195 B.n421 B.n128 10.6151
R1196 B.n425 B.n128 10.6151
R1197 B.n426 B.n425 10.6151
R1198 B.n427 B.n426 10.6151
R1199 B.n427 B.n126 10.6151
R1200 B.n431 B.n126 10.6151
R1201 B.n432 B.n431 10.6151
R1202 B.n433 B.n432 10.6151
R1203 B.n433 B.n124 10.6151
R1204 B.n437 B.n124 10.6151
R1205 B.n438 B.n437 10.6151
R1206 B.n439 B.n438 10.6151
R1207 B.n439 B.n122 10.6151
R1208 B.n443 B.n122 10.6151
R1209 B.n444 B.n443 10.6151
R1210 B.n445 B.n444 10.6151
R1211 B.n252 B.n251 10.6151
R1212 B.n251 B.n190 10.6151
R1213 B.n247 B.n190 10.6151
R1214 B.n247 B.n246 10.6151
R1215 B.n246 B.n245 10.6151
R1216 B.n245 B.n192 10.6151
R1217 B.n241 B.n192 10.6151
R1218 B.n241 B.n240 10.6151
R1219 B.n240 B.n239 10.6151
R1220 B.n239 B.n194 10.6151
R1221 B.n235 B.n194 10.6151
R1222 B.n235 B.n234 10.6151
R1223 B.n234 B.n233 10.6151
R1224 B.n233 B.n196 10.6151
R1225 B.n229 B.n196 10.6151
R1226 B.n229 B.n228 10.6151
R1227 B.n228 B.n227 10.6151
R1228 B.n227 B.n198 10.6151
R1229 B.n223 B.n198 10.6151
R1230 B.n223 B.n222 10.6151
R1231 B.n222 B.n221 10.6151
R1232 B.n221 B.n200 10.6151
R1233 B.n217 B.n200 10.6151
R1234 B.n217 B.n216 10.6151
R1235 B.n216 B.n215 10.6151
R1236 B.n215 B.n202 10.6151
R1237 B.n211 B.n202 10.6151
R1238 B.n211 B.n210 10.6151
R1239 B.n210 B.n209 10.6151
R1240 B.n209 B.n204 10.6151
R1241 B.n205 B.n204 10.6151
R1242 B.n205 B.n0 10.6151
R1243 B.n787 B.n1 10.6151
R1244 B.n787 B.n786 10.6151
R1245 B.n786 B.n785 10.6151
R1246 B.n785 B.n4 10.6151
R1247 B.n781 B.n4 10.6151
R1248 B.n781 B.n780 10.6151
R1249 B.n780 B.n779 10.6151
R1250 B.n779 B.n6 10.6151
R1251 B.n775 B.n6 10.6151
R1252 B.n775 B.n774 10.6151
R1253 B.n774 B.n773 10.6151
R1254 B.n773 B.n8 10.6151
R1255 B.n769 B.n8 10.6151
R1256 B.n769 B.n768 10.6151
R1257 B.n768 B.n767 10.6151
R1258 B.n767 B.n10 10.6151
R1259 B.n763 B.n10 10.6151
R1260 B.n763 B.n762 10.6151
R1261 B.n762 B.n761 10.6151
R1262 B.n761 B.n12 10.6151
R1263 B.n757 B.n12 10.6151
R1264 B.n757 B.n756 10.6151
R1265 B.n756 B.n755 10.6151
R1266 B.n755 B.n14 10.6151
R1267 B.n751 B.n14 10.6151
R1268 B.n751 B.n750 10.6151
R1269 B.n750 B.n749 10.6151
R1270 B.n749 B.n16 10.6151
R1271 B.n745 B.n16 10.6151
R1272 B.n745 B.n744 10.6151
R1273 B.n744 B.n743 10.6151
R1274 B.n743 B.n18 10.6151
R1275 B.n653 B.n50 9.36635
R1276 B.n636 B.n635 9.36635
R1277 B.n342 B.n341 9.36635
R1278 B.n359 B.n152 9.36635
R1279 B.n791 B.n0 2.81026
R1280 B.n791 B.n1 2.81026
R1281 B.n650 B.n50 1.24928
R1282 B.n637 B.n636 1.24928
R1283 B.n343 B.n342 1.24928
R1284 B.n356 B.n152 1.24928
R1285 VN.n2 VN.t4 278.62
R1286 VN.n14 VN.t0 278.62
R1287 VN.n3 VN.t5 242.617
R1288 VN.n10 VN.t3 242.617
R1289 VN.n15 VN.t2 242.617
R1290 VN.n22 VN.t1 242.617
R1291 VN.n11 VN.n10 179.99
R1292 VN.n23 VN.n22 179.99
R1293 VN.n21 VN.n12 161.3
R1294 VN.n20 VN.n19 161.3
R1295 VN.n18 VN.n13 161.3
R1296 VN.n17 VN.n16 161.3
R1297 VN.n9 VN.n0 161.3
R1298 VN.n8 VN.n7 161.3
R1299 VN.n6 VN.n1 161.3
R1300 VN.n5 VN.n4 161.3
R1301 VN VN.n23 50.3736
R1302 VN.n8 VN.n1 46.3896
R1303 VN.n20 VN.n13 46.3896
R1304 VN.n15 VN.n14 44.58
R1305 VN.n3 VN.n2 44.58
R1306 VN.n4 VN.n1 34.7644
R1307 VN.n16 VN.n13 34.7644
R1308 VN.n4 VN.n3 24.5923
R1309 VN.n9 VN.n8 24.5923
R1310 VN.n16 VN.n15 24.5923
R1311 VN.n21 VN.n20 24.5923
R1312 VN.n17 VN.n14 12.1133
R1313 VN.n5 VN.n2 12.1133
R1314 VN.n10 VN.n9 5.90254
R1315 VN.n22 VN.n21 5.90254
R1316 VN.n23 VN.n12 0.189894
R1317 VN.n19 VN.n12 0.189894
R1318 VN.n19 VN.n18 0.189894
R1319 VN.n18 VN.n17 0.189894
R1320 VN.n6 VN.n5 0.189894
R1321 VN.n7 VN.n6 0.189894
R1322 VN.n7 VN.n0 0.189894
R1323 VN.n11 VN.n0 0.189894
R1324 VN VN.n11 0.0516364
R1325 VDD2.n1 VDD2.t1 74.6848
R1326 VDD2.n2 VDD2.t4 73.3697
R1327 VDD2.n1 VDD2.n0 71.9671
R1328 VDD2 VDD2.n3 71.9644
R1329 VDD2.n2 VDD2.n1 45.1894
R1330 VDD2.n3 VDD2.t3 1.80433
R1331 VDD2.n3 VDD2.t5 1.80433
R1332 VDD2.n0 VDD2.t0 1.80433
R1333 VDD2.n0 VDD2.t2 1.80433
R1334 VDD2 VDD2.n2 1.42938
C0 B VN 1.06972f
C1 VTAIL w_n2666_n4572# 3.78524f
C2 VN VDD2 9.101f
C3 VTAIL VDD1 10.345099f
C4 VTAIL VP 8.83786f
C5 w_n2666_n4572# B 10.2451f
C6 B VDD1 2.34007f
C7 w_n2666_n4572# VDD2 2.5765f
C8 B VP 1.63735f
C9 VDD1 VDD2 1.117f
C10 w_n2666_n4572# VN 4.95845f
C11 VP VDD2 0.390543f
C12 VDD1 VN 0.149841f
C13 VTAIL B 4.59138f
C14 VP VN 7.24827f
C15 VTAIL VDD2 10.3875f
C16 w_n2666_n4572# VDD1 2.51735f
C17 VTAIL VN 8.82335f
C18 w_n2666_n4572# VP 5.30087f
C19 B VDD2 2.39477f
C20 VP VDD1 9.336821f
C21 VDD2 VSUBS 1.854546f
C22 VDD1 VSUBS 2.261043f
C23 VTAIL VSUBS 1.256679f
C24 VN VSUBS 5.4157f
C25 VP VSUBS 2.516816f
C26 B VSUBS 4.346079f
C27 w_n2666_n4572# VSUBS 0.149051p
C28 VDD2.t1 VSUBS 4.16378f
C29 VDD2.t0 VSUBS 0.383639f
C30 VDD2.t2 VSUBS 0.383639f
C31 VDD2.n0 VSUBS 3.20346f
C32 VDD2.n1 VSUBS 3.77276f
C33 VDD2.t4 VSUBS 4.15075f
C34 VDD2.n2 VSUBS 3.59299f
C35 VDD2.t3 VSUBS 0.383639f
C36 VDD2.t5 VSUBS 0.383639f
C37 VDD2.n3 VSUBS 3.20341f
C38 VN.n0 VSUBS 0.033969f
C39 VN.t3 VSUBS 3.01388f
C40 VN.n1 VSUBS 0.029027f
C41 VN.t4 VSUBS 3.17089f
C42 VN.n2 VSUBS 1.12594f
C43 VN.t5 VSUBS 3.01388f
C44 VN.n3 VSUBS 1.14578f
C45 VN.n4 VSUBS 0.06827f
C46 VN.n5 VSUBS 0.250967f
C47 VN.n6 VSUBS 0.033969f
C48 VN.n7 VSUBS 0.033969f
C49 VN.n8 VSUBS 0.064454f
C50 VN.n9 VSUBS 0.039358f
C51 VN.n10 VSUBS 1.13396f
C52 VN.n11 VSUBS 0.035514f
C53 VN.n12 VSUBS 0.033969f
C54 VN.t1 VSUBS 3.01388f
C55 VN.n13 VSUBS 0.029027f
C56 VN.t0 VSUBS 3.17089f
C57 VN.n14 VSUBS 1.12594f
C58 VN.t2 VSUBS 3.01388f
C59 VN.n15 VSUBS 1.14578f
C60 VN.n16 VSUBS 0.06827f
C61 VN.n17 VSUBS 0.250967f
C62 VN.n18 VSUBS 0.033969f
C63 VN.n19 VSUBS 0.033969f
C64 VN.n20 VSUBS 0.064454f
C65 VN.n21 VSUBS 0.039358f
C66 VN.n22 VSUBS 1.13396f
C67 VN.n23 VSUBS 1.87764f
C68 B.n0 VSUBS 0.004896f
C69 B.n1 VSUBS 0.004896f
C70 B.n2 VSUBS 0.007743f
C71 B.n3 VSUBS 0.007743f
C72 B.n4 VSUBS 0.007743f
C73 B.n5 VSUBS 0.007743f
C74 B.n6 VSUBS 0.007743f
C75 B.n7 VSUBS 0.007743f
C76 B.n8 VSUBS 0.007743f
C77 B.n9 VSUBS 0.007743f
C78 B.n10 VSUBS 0.007743f
C79 B.n11 VSUBS 0.007743f
C80 B.n12 VSUBS 0.007743f
C81 B.n13 VSUBS 0.007743f
C82 B.n14 VSUBS 0.007743f
C83 B.n15 VSUBS 0.007743f
C84 B.n16 VSUBS 0.007743f
C85 B.n17 VSUBS 0.007743f
C86 B.n18 VSUBS 0.0183f
C87 B.n19 VSUBS 0.007743f
C88 B.n20 VSUBS 0.007743f
C89 B.n21 VSUBS 0.007743f
C90 B.n22 VSUBS 0.007743f
C91 B.n23 VSUBS 0.007743f
C92 B.n24 VSUBS 0.007743f
C93 B.n25 VSUBS 0.007743f
C94 B.n26 VSUBS 0.007743f
C95 B.n27 VSUBS 0.007743f
C96 B.n28 VSUBS 0.007743f
C97 B.n29 VSUBS 0.007743f
C98 B.n30 VSUBS 0.007743f
C99 B.n31 VSUBS 0.007743f
C100 B.n32 VSUBS 0.007743f
C101 B.n33 VSUBS 0.007743f
C102 B.n34 VSUBS 0.007743f
C103 B.n35 VSUBS 0.007743f
C104 B.n36 VSUBS 0.007743f
C105 B.n37 VSUBS 0.007743f
C106 B.n38 VSUBS 0.007743f
C107 B.n39 VSUBS 0.007743f
C108 B.n40 VSUBS 0.007743f
C109 B.n41 VSUBS 0.007743f
C110 B.n42 VSUBS 0.007743f
C111 B.n43 VSUBS 0.007743f
C112 B.n44 VSUBS 0.007743f
C113 B.n45 VSUBS 0.007743f
C114 B.n46 VSUBS 0.007743f
C115 B.n47 VSUBS 0.007743f
C116 B.t8 VSUBS 0.672957f
C117 B.t7 VSUBS 0.69032f
C118 B.t6 VSUBS 1.53795f
C119 B.n48 VSUBS 0.326692f
C120 B.n49 VSUBS 0.076027f
C121 B.n50 VSUBS 0.017939f
C122 B.n51 VSUBS 0.007743f
C123 B.n52 VSUBS 0.007743f
C124 B.n53 VSUBS 0.007743f
C125 B.n54 VSUBS 0.007743f
C126 B.n55 VSUBS 0.007743f
C127 B.t2 VSUBS 0.672933f
C128 B.t1 VSUBS 0.690299f
C129 B.t0 VSUBS 1.53795f
C130 B.n56 VSUBS 0.326712f
C131 B.n57 VSUBS 0.076051f
C132 B.n58 VSUBS 0.007743f
C133 B.n59 VSUBS 0.007743f
C134 B.n60 VSUBS 0.007743f
C135 B.n61 VSUBS 0.007743f
C136 B.n62 VSUBS 0.007743f
C137 B.n63 VSUBS 0.007743f
C138 B.n64 VSUBS 0.007743f
C139 B.n65 VSUBS 0.007743f
C140 B.n66 VSUBS 0.007743f
C141 B.n67 VSUBS 0.007743f
C142 B.n68 VSUBS 0.007743f
C143 B.n69 VSUBS 0.007743f
C144 B.n70 VSUBS 0.007743f
C145 B.n71 VSUBS 0.007743f
C146 B.n72 VSUBS 0.007743f
C147 B.n73 VSUBS 0.007743f
C148 B.n74 VSUBS 0.007743f
C149 B.n75 VSUBS 0.007743f
C150 B.n76 VSUBS 0.007743f
C151 B.n77 VSUBS 0.007743f
C152 B.n78 VSUBS 0.007743f
C153 B.n79 VSUBS 0.007743f
C154 B.n80 VSUBS 0.007743f
C155 B.n81 VSUBS 0.007743f
C156 B.n82 VSUBS 0.007743f
C157 B.n83 VSUBS 0.007743f
C158 B.n84 VSUBS 0.007743f
C159 B.n85 VSUBS 0.007743f
C160 B.n86 VSUBS 0.007743f
C161 B.n87 VSUBS 0.0183f
C162 B.n88 VSUBS 0.007743f
C163 B.n89 VSUBS 0.007743f
C164 B.n90 VSUBS 0.007743f
C165 B.n91 VSUBS 0.007743f
C166 B.n92 VSUBS 0.007743f
C167 B.n93 VSUBS 0.007743f
C168 B.n94 VSUBS 0.007743f
C169 B.n95 VSUBS 0.007743f
C170 B.n96 VSUBS 0.007743f
C171 B.n97 VSUBS 0.007743f
C172 B.n98 VSUBS 0.007743f
C173 B.n99 VSUBS 0.007743f
C174 B.n100 VSUBS 0.007743f
C175 B.n101 VSUBS 0.007743f
C176 B.n102 VSUBS 0.007743f
C177 B.n103 VSUBS 0.007743f
C178 B.n104 VSUBS 0.007743f
C179 B.n105 VSUBS 0.007743f
C180 B.n106 VSUBS 0.007743f
C181 B.n107 VSUBS 0.007743f
C182 B.n108 VSUBS 0.007743f
C183 B.n109 VSUBS 0.007743f
C184 B.n110 VSUBS 0.007743f
C185 B.n111 VSUBS 0.007743f
C186 B.n112 VSUBS 0.007743f
C187 B.n113 VSUBS 0.007743f
C188 B.n114 VSUBS 0.007743f
C189 B.n115 VSUBS 0.007743f
C190 B.n116 VSUBS 0.007743f
C191 B.n117 VSUBS 0.007743f
C192 B.n118 VSUBS 0.007743f
C193 B.n119 VSUBS 0.007743f
C194 B.n120 VSUBS 0.0183f
C195 B.n121 VSUBS 0.007743f
C196 B.n122 VSUBS 0.007743f
C197 B.n123 VSUBS 0.007743f
C198 B.n124 VSUBS 0.007743f
C199 B.n125 VSUBS 0.007743f
C200 B.n126 VSUBS 0.007743f
C201 B.n127 VSUBS 0.007743f
C202 B.n128 VSUBS 0.007743f
C203 B.n129 VSUBS 0.007743f
C204 B.n130 VSUBS 0.007743f
C205 B.n131 VSUBS 0.007743f
C206 B.n132 VSUBS 0.007743f
C207 B.n133 VSUBS 0.007743f
C208 B.n134 VSUBS 0.007743f
C209 B.n135 VSUBS 0.007743f
C210 B.n136 VSUBS 0.007743f
C211 B.n137 VSUBS 0.007743f
C212 B.n138 VSUBS 0.007743f
C213 B.n139 VSUBS 0.007743f
C214 B.n140 VSUBS 0.007743f
C215 B.n141 VSUBS 0.007743f
C216 B.n142 VSUBS 0.007743f
C217 B.n143 VSUBS 0.007743f
C218 B.n144 VSUBS 0.007743f
C219 B.n145 VSUBS 0.007743f
C220 B.n146 VSUBS 0.007743f
C221 B.n147 VSUBS 0.007743f
C222 B.n148 VSUBS 0.007743f
C223 B.n149 VSUBS 0.007743f
C224 B.t10 VSUBS 0.672933f
C225 B.t11 VSUBS 0.690299f
C226 B.t9 VSUBS 1.53795f
C227 B.n150 VSUBS 0.326712f
C228 B.n151 VSUBS 0.076051f
C229 B.n152 VSUBS 0.017939f
C230 B.n153 VSUBS 0.007743f
C231 B.n154 VSUBS 0.007743f
C232 B.n155 VSUBS 0.007743f
C233 B.n156 VSUBS 0.007743f
C234 B.n157 VSUBS 0.007743f
C235 B.t4 VSUBS 0.672957f
C236 B.t5 VSUBS 0.69032f
C237 B.t3 VSUBS 1.53795f
C238 B.n158 VSUBS 0.326692f
C239 B.n159 VSUBS 0.076027f
C240 B.n160 VSUBS 0.007743f
C241 B.n161 VSUBS 0.007743f
C242 B.n162 VSUBS 0.007743f
C243 B.n163 VSUBS 0.007743f
C244 B.n164 VSUBS 0.007743f
C245 B.n165 VSUBS 0.007743f
C246 B.n166 VSUBS 0.007743f
C247 B.n167 VSUBS 0.007743f
C248 B.n168 VSUBS 0.007743f
C249 B.n169 VSUBS 0.007743f
C250 B.n170 VSUBS 0.007743f
C251 B.n171 VSUBS 0.007743f
C252 B.n172 VSUBS 0.007743f
C253 B.n173 VSUBS 0.007743f
C254 B.n174 VSUBS 0.007743f
C255 B.n175 VSUBS 0.007743f
C256 B.n176 VSUBS 0.007743f
C257 B.n177 VSUBS 0.007743f
C258 B.n178 VSUBS 0.007743f
C259 B.n179 VSUBS 0.007743f
C260 B.n180 VSUBS 0.007743f
C261 B.n181 VSUBS 0.007743f
C262 B.n182 VSUBS 0.007743f
C263 B.n183 VSUBS 0.007743f
C264 B.n184 VSUBS 0.007743f
C265 B.n185 VSUBS 0.007743f
C266 B.n186 VSUBS 0.007743f
C267 B.n187 VSUBS 0.007743f
C268 B.n188 VSUBS 0.007743f
C269 B.n189 VSUBS 0.0183f
C270 B.n190 VSUBS 0.007743f
C271 B.n191 VSUBS 0.007743f
C272 B.n192 VSUBS 0.007743f
C273 B.n193 VSUBS 0.007743f
C274 B.n194 VSUBS 0.007743f
C275 B.n195 VSUBS 0.007743f
C276 B.n196 VSUBS 0.007743f
C277 B.n197 VSUBS 0.007743f
C278 B.n198 VSUBS 0.007743f
C279 B.n199 VSUBS 0.007743f
C280 B.n200 VSUBS 0.007743f
C281 B.n201 VSUBS 0.007743f
C282 B.n202 VSUBS 0.007743f
C283 B.n203 VSUBS 0.007743f
C284 B.n204 VSUBS 0.007743f
C285 B.n205 VSUBS 0.007743f
C286 B.n206 VSUBS 0.007743f
C287 B.n207 VSUBS 0.007743f
C288 B.n208 VSUBS 0.007743f
C289 B.n209 VSUBS 0.007743f
C290 B.n210 VSUBS 0.007743f
C291 B.n211 VSUBS 0.007743f
C292 B.n212 VSUBS 0.007743f
C293 B.n213 VSUBS 0.007743f
C294 B.n214 VSUBS 0.007743f
C295 B.n215 VSUBS 0.007743f
C296 B.n216 VSUBS 0.007743f
C297 B.n217 VSUBS 0.007743f
C298 B.n218 VSUBS 0.007743f
C299 B.n219 VSUBS 0.007743f
C300 B.n220 VSUBS 0.007743f
C301 B.n221 VSUBS 0.007743f
C302 B.n222 VSUBS 0.007743f
C303 B.n223 VSUBS 0.007743f
C304 B.n224 VSUBS 0.007743f
C305 B.n225 VSUBS 0.007743f
C306 B.n226 VSUBS 0.007743f
C307 B.n227 VSUBS 0.007743f
C308 B.n228 VSUBS 0.007743f
C309 B.n229 VSUBS 0.007743f
C310 B.n230 VSUBS 0.007743f
C311 B.n231 VSUBS 0.007743f
C312 B.n232 VSUBS 0.007743f
C313 B.n233 VSUBS 0.007743f
C314 B.n234 VSUBS 0.007743f
C315 B.n235 VSUBS 0.007743f
C316 B.n236 VSUBS 0.007743f
C317 B.n237 VSUBS 0.007743f
C318 B.n238 VSUBS 0.007743f
C319 B.n239 VSUBS 0.007743f
C320 B.n240 VSUBS 0.007743f
C321 B.n241 VSUBS 0.007743f
C322 B.n242 VSUBS 0.007743f
C323 B.n243 VSUBS 0.007743f
C324 B.n244 VSUBS 0.007743f
C325 B.n245 VSUBS 0.007743f
C326 B.n246 VSUBS 0.007743f
C327 B.n247 VSUBS 0.007743f
C328 B.n248 VSUBS 0.007743f
C329 B.n249 VSUBS 0.007743f
C330 B.n250 VSUBS 0.007743f
C331 B.n251 VSUBS 0.007743f
C332 B.n252 VSUBS 0.0183f
C333 B.n253 VSUBS 0.019046f
C334 B.n254 VSUBS 0.019046f
C335 B.n255 VSUBS 0.007743f
C336 B.n256 VSUBS 0.007743f
C337 B.n257 VSUBS 0.007743f
C338 B.n258 VSUBS 0.007743f
C339 B.n259 VSUBS 0.007743f
C340 B.n260 VSUBS 0.007743f
C341 B.n261 VSUBS 0.007743f
C342 B.n262 VSUBS 0.007743f
C343 B.n263 VSUBS 0.007743f
C344 B.n264 VSUBS 0.007743f
C345 B.n265 VSUBS 0.007743f
C346 B.n266 VSUBS 0.007743f
C347 B.n267 VSUBS 0.007743f
C348 B.n268 VSUBS 0.007743f
C349 B.n269 VSUBS 0.007743f
C350 B.n270 VSUBS 0.007743f
C351 B.n271 VSUBS 0.007743f
C352 B.n272 VSUBS 0.007743f
C353 B.n273 VSUBS 0.007743f
C354 B.n274 VSUBS 0.007743f
C355 B.n275 VSUBS 0.007743f
C356 B.n276 VSUBS 0.007743f
C357 B.n277 VSUBS 0.007743f
C358 B.n278 VSUBS 0.007743f
C359 B.n279 VSUBS 0.007743f
C360 B.n280 VSUBS 0.007743f
C361 B.n281 VSUBS 0.007743f
C362 B.n282 VSUBS 0.007743f
C363 B.n283 VSUBS 0.007743f
C364 B.n284 VSUBS 0.007743f
C365 B.n285 VSUBS 0.007743f
C366 B.n286 VSUBS 0.007743f
C367 B.n287 VSUBS 0.007743f
C368 B.n288 VSUBS 0.007743f
C369 B.n289 VSUBS 0.007743f
C370 B.n290 VSUBS 0.007743f
C371 B.n291 VSUBS 0.007743f
C372 B.n292 VSUBS 0.007743f
C373 B.n293 VSUBS 0.007743f
C374 B.n294 VSUBS 0.007743f
C375 B.n295 VSUBS 0.007743f
C376 B.n296 VSUBS 0.007743f
C377 B.n297 VSUBS 0.007743f
C378 B.n298 VSUBS 0.007743f
C379 B.n299 VSUBS 0.007743f
C380 B.n300 VSUBS 0.007743f
C381 B.n301 VSUBS 0.007743f
C382 B.n302 VSUBS 0.007743f
C383 B.n303 VSUBS 0.007743f
C384 B.n304 VSUBS 0.007743f
C385 B.n305 VSUBS 0.007743f
C386 B.n306 VSUBS 0.007743f
C387 B.n307 VSUBS 0.007743f
C388 B.n308 VSUBS 0.007743f
C389 B.n309 VSUBS 0.007743f
C390 B.n310 VSUBS 0.007743f
C391 B.n311 VSUBS 0.007743f
C392 B.n312 VSUBS 0.007743f
C393 B.n313 VSUBS 0.007743f
C394 B.n314 VSUBS 0.007743f
C395 B.n315 VSUBS 0.007743f
C396 B.n316 VSUBS 0.007743f
C397 B.n317 VSUBS 0.007743f
C398 B.n318 VSUBS 0.007743f
C399 B.n319 VSUBS 0.007743f
C400 B.n320 VSUBS 0.007743f
C401 B.n321 VSUBS 0.007743f
C402 B.n322 VSUBS 0.007743f
C403 B.n323 VSUBS 0.007743f
C404 B.n324 VSUBS 0.007743f
C405 B.n325 VSUBS 0.007743f
C406 B.n326 VSUBS 0.007743f
C407 B.n327 VSUBS 0.007743f
C408 B.n328 VSUBS 0.007743f
C409 B.n329 VSUBS 0.007743f
C410 B.n330 VSUBS 0.007743f
C411 B.n331 VSUBS 0.007743f
C412 B.n332 VSUBS 0.007743f
C413 B.n333 VSUBS 0.007743f
C414 B.n334 VSUBS 0.007743f
C415 B.n335 VSUBS 0.007743f
C416 B.n336 VSUBS 0.007743f
C417 B.n337 VSUBS 0.007743f
C418 B.n338 VSUBS 0.007743f
C419 B.n339 VSUBS 0.007743f
C420 B.n340 VSUBS 0.007743f
C421 B.n341 VSUBS 0.007287f
C422 B.n342 VSUBS 0.017939f
C423 B.n343 VSUBS 0.004327f
C424 B.n344 VSUBS 0.007743f
C425 B.n345 VSUBS 0.007743f
C426 B.n346 VSUBS 0.007743f
C427 B.n347 VSUBS 0.007743f
C428 B.n348 VSUBS 0.007743f
C429 B.n349 VSUBS 0.007743f
C430 B.n350 VSUBS 0.007743f
C431 B.n351 VSUBS 0.007743f
C432 B.n352 VSUBS 0.007743f
C433 B.n353 VSUBS 0.007743f
C434 B.n354 VSUBS 0.007743f
C435 B.n355 VSUBS 0.007743f
C436 B.n356 VSUBS 0.004327f
C437 B.n357 VSUBS 0.007743f
C438 B.n358 VSUBS 0.007743f
C439 B.n359 VSUBS 0.007287f
C440 B.n360 VSUBS 0.007743f
C441 B.n361 VSUBS 0.007743f
C442 B.n362 VSUBS 0.007743f
C443 B.n363 VSUBS 0.007743f
C444 B.n364 VSUBS 0.007743f
C445 B.n365 VSUBS 0.007743f
C446 B.n366 VSUBS 0.007743f
C447 B.n367 VSUBS 0.007743f
C448 B.n368 VSUBS 0.007743f
C449 B.n369 VSUBS 0.007743f
C450 B.n370 VSUBS 0.007743f
C451 B.n371 VSUBS 0.007743f
C452 B.n372 VSUBS 0.007743f
C453 B.n373 VSUBS 0.007743f
C454 B.n374 VSUBS 0.007743f
C455 B.n375 VSUBS 0.007743f
C456 B.n376 VSUBS 0.007743f
C457 B.n377 VSUBS 0.007743f
C458 B.n378 VSUBS 0.007743f
C459 B.n379 VSUBS 0.007743f
C460 B.n380 VSUBS 0.007743f
C461 B.n381 VSUBS 0.007743f
C462 B.n382 VSUBS 0.007743f
C463 B.n383 VSUBS 0.007743f
C464 B.n384 VSUBS 0.007743f
C465 B.n385 VSUBS 0.007743f
C466 B.n386 VSUBS 0.007743f
C467 B.n387 VSUBS 0.007743f
C468 B.n388 VSUBS 0.007743f
C469 B.n389 VSUBS 0.007743f
C470 B.n390 VSUBS 0.007743f
C471 B.n391 VSUBS 0.007743f
C472 B.n392 VSUBS 0.007743f
C473 B.n393 VSUBS 0.007743f
C474 B.n394 VSUBS 0.007743f
C475 B.n395 VSUBS 0.007743f
C476 B.n396 VSUBS 0.007743f
C477 B.n397 VSUBS 0.007743f
C478 B.n398 VSUBS 0.007743f
C479 B.n399 VSUBS 0.007743f
C480 B.n400 VSUBS 0.007743f
C481 B.n401 VSUBS 0.007743f
C482 B.n402 VSUBS 0.007743f
C483 B.n403 VSUBS 0.007743f
C484 B.n404 VSUBS 0.007743f
C485 B.n405 VSUBS 0.007743f
C486 B.n406 VSUBS 0.007743f
C487 B.n407 VSUBS 0.007743f
C488 B.n408 VSUBS 0.007743f
C489 B.n409 VSUBS 0.007743f
C490 B.n410 VSUBS 0.007743f
C491 B.n411 VSUBS 0.007743f
C492 B.n412 VSUBS 0.007743f
C493 B.n413 VSUBS 0.007743f
C494 B.n414 VSUBS 0.007743f
C495 B.n415 VSUBS 0.007743f
C496 B.n416 VSUBS 0.007743f
C497 B.n417 VSUBS 0.007743f
C498 B.n418 VSUBS 0.007743f
C499 B.n419 VSUBS 0.007743f
C500 B.n420 VSUBS 0.007743f
C501 B.n421 VSUBS 0.007743f
C502 B.n422 VSUBS 0.007743f
C503 B.n423 VSUBS 0.007743f
C504 B.n424 VSUBS 0.007743f
C505 B.n425 VSUBS 0.007743f
C506 B.n426 VSUBS 0.007743f
C507 B.n427 VSUBS 0.007743f
C508 B.n428 VSUBS 0.007743f
C509 B.n429 VSUBS 0.007743f
C510 B.n430 VSUBS 0.007743f
C511 B.n431 VSUBS 0.007743f
C512 B.n432 VSUBS 0.007743f
C513 B.n433 VSUBS 0.007743f
C514 B.n434 VSUBS 0.007743f
C515 B.n435 VSUBS 0.007743f
C516 B.n436 VSUBS 0.007743f
C517 B.n437 VSUBS 0.007743f
C518 B.n438 VSUBS 0.007743f
C519 B.n439 VSUBS 0.007743f
C520 B.n440 VSUBS 0.007743f
C521 B.n441 VSUBS 0.007743f
C522 B.n442 VSUBS 0.007743f
C523 B.n443 VSUBS 0.007743f
C524 B.n444 VSUBS 0.007743f
C525 B.n445 VSUBS 0.019046f
C526 B.n446 VSUBS 0.019046f
C527 B.n447 VSUBS 0.0183f
C528 B.n448 VSUBS 0.007743f
C529 B.n449 VSUBS 0.007743f
C530 B.n450 VSUBS 0.007743f
C531 B.n451 VSUBS 0.007743f
C532 B.n452 VSUBS 0.007743f
C533 B.n453 VSUBS 0.007743f
C534 B.n454 VSUBS 0.007743f
C535 B.n455 VSUBS 0.007743f
C536 B.n456 VSUBS 0.007743f
C537 B.n457 VSUBS 0.007743f
C538 B.n458 VSUBS 0.007743f
C539 B.n459 VSUBS 0.007743f
C540 B.n460 VSUBS 0.007743f
C541 B.n461 VSUBS 0.007743f
C542 B.n462 VSUBS 0.007743f
C543 B.n463 VSUBS 0.007743f
C544 B.n464 VSUBS 0.007743f
C545 B.n465 VSUBS 0.007743f
C546 B.n466 VSUBS 0.007743f
C547 B.n467 VSUBS 0.007743f
C548 B.n468 VSUBS 0.007743f
C549 B.n469 VSUBS 0.007743f
C550 B.n470 VSUBS 0.007743f
C551 B.n471 VSUBS 0.007743f
C552 B.n472 VSUBS 0.007743f
C553 B.n473 VSUBS 0.007743f
C554 B.n474 VSUBS 0.007743f
C555 B.n475 VSUBS 0.007743f
C556 B.n476 VSUBS 0.007743f
C557 B.n477 VSUBS 0.007743f
C558 B.n478 VSUBS 0.007743f
C559 B.n479 VSUBS 0.007743f
C560 B.n480 VSUBS 0.007743f
C561 B.n481 VSUBS 0.007743f
C562 B.n482 VSUBS 0.007743f
C563 B.n483 VSUBS 0.007743f
C564 B.n484 VSUBS 0.007743f
C565 B.n485 VSUBS 0.007743f
C566 B.n486 VSUBS 0.007743f
C567 B.n487 VSUBS 0.007743f
C568 B.n488 VSUBS 0.007743f
C569 B.n489 VSUBS 0.007743f
C570 B.n490 VSUBS 0.007743f
C571 B.n491 VSUBS 0.007743f
C572 B.n492 VSUBS 0.007743f
C573 B.n493 VSUBS 0.007743f
C574 B.n494 VSUBS 0.007743f
C575 B.n495 VSUBS 0.007743f
C576 B.n496 VSUBS 0.007743f
C577 B.n497 VSUBS 0.007743f
C578 B.n498 VSUBS 0.007743f
C579 B.n499 VSUBS 0.007743f
C580 B.n500 VSUBS 0.007743f
C581 B.n501 VSUBS 0.007743f
C582 B.n502 VSUBS 0.007743f
C583 B.n503 VSUBS 0.007743f
C584 B.n504 VSUBS 0.007743f
C585 B.n505 VSUBS 0.007743f
C586 B.n506 VSUBS 0.007743f
C587 B.n507 VSUBS 0.007743f
C588 B.n508 VSUBS 0.007743f
C589 B.n509 VSUBS 0.007743f
C590 B.n510 VSUBS 0.007743f
C591 B.n511 VSUBS 0.007743f
C592 B.n512 VSUBS 0.007743f
C593 B.n513 VSUBS 0.007743f
C594 B.n514 VSUBS 0.007743f
C595 B.n515 VSUBS 0.007743f
C596 B.n516 VSUBS 0.007743f
C597 B.n517 VSUBS 0.007743f
C598 B.n518 VSUBS 0.007743f
C599 B.n519 VSUBS 0.007743f
C600 B.n520 VSUBS 0.007743f
C601 B.n521 VSUBS 0.007743f
C602 B.n522 VSUBS 0.007743f
C603 B.n523 VSUBS 0.007743f
C604 B.n524 VSUBS 0.007743f
C605 B.n525 VSUBS 0.007743f
C606 B.n526 VSUBS 0.007743f
C607 B.n527 VSUBS 0.007743f
C608 B.n528 VSUBS 0.007743f
C609 B.n529 VSUBS 0.007743f
C610 B.n530 VSUBS 0.007743f
C611 B.n531 VSUBS 0.007743f
C612 B.n532 VSUBS 0.007743f
C613 B.n533 VSUBS 0.007743f
C614 B.n534 VSUBS 0.007743f
C615 B.n535 VSUBS 0.007743f
C616 B.n536 VSUBS 0.007743f
C617 B.n537 VSUBS 0.007743f
C618 B.n538 VSUBS 0.007743f
C619 B.n539 VSUBS 0.007743f
C620 B.n540 VSUBS 0.007743f
C621 B.n541 VSUBS 0.007743f
C622 B.n542 VSUBS 0.007743f
C623 B.n543 VSUBS 0.007743f
C624 B.n544 VSUBS 0.007743f
C625 B.n545 VSUBS 0.007743f
C626 B.n546 VSUBS 0.019174f
C627 B.n547 VSUBS 0.018172f
C628 B.n548 VSUBS 0.019046f
C629 B.n549 VSUBS 0.007743f
C630 B.n550 VSUBS 0.007743f
C631 B.n551 VSUBS 0.007743f
C632 B.n552 VSUBS 0.007743f
C633 B.n553 VSUBS 0.007743f
C634 B.n554 VSUBS 0.007743f
C635 B.n555 VSUBS 0.007743f
C636 B.n556 VSUBS 0.007743f
C637 B.n557 VSUBS 0.007743f
C638 B.n558 VSUBS 0.007743f
C639 B.n559 VSUBS 0.007743f
C640 B.n560 VSUBS 0.007743f
C641 B.n561 VSUBS 0.007743f
C642 B.n562 VSUBS 0.007743f
C643 B.n563 VSUBS 0.007743f
C644 B.n564 VSUBS 0.007743f
C645 B.n565 VSUBS 0.007743f
C646 B.n566 VSUBS 0.007743f
C647 B.n567 VSUBS 0.007743f
C648 B.n568 VSUBS 0.007743f
C649 B.n569 VSUBS 0.007743f
C650 B.n570 VSUBS 0.007743f
C651 B.n571 VSUBS 0.007743f
C652 B.n572 VSUBS 0.007743f
C653 B.n573 VSUBS 0.007743f
C654 B.n574 VSUBS 0.007743f
C655 B.n575 VSUBS 0.007743f
C656 B.n576 VSUBS 0.007743f
C657 B.n577 VSUBS 0.007743f
C658 B.n578 VSUBS 0.007743f
C659 B.n579 VSUBS 0.007743f
C660 B.n580 VSUBS 0.007743f
C661 B.n581 VSUBS 0.007743f
C662 B.n582 VSUBS 0.007743f
C663 B.n583 VSUBS 0.007743f
C664 B.n584 VSUBS 0.007743f
C665 B.n585 VSUBS 0.007743f
C666 B.n586 VSUBS 0.007743f
C667 B.n587 VSUBS 0.007743f
C668 B.n588 VSUBS 0.007743f
C669 B.n589 VSUBS 0.007743f
C670 B.n590 VSUBS 0.007743f
C671 B.n591 VSUBS 0.007743f
C672 B.n592 VSUBS 0.007743f
C673 B.n593 VSUBS 0.007743f
C674 B.n594 VSUBS 0.007743f
C675 B.n595 VSUBS 0.007743f
C676 B.n596 VSUBS 0.007743f
C677 B.n597 VSUBS 0.007743f
C678 B.n598 VSUBS 0.007743f
C679 B.n599 VSUBS 0.007743f
C680 B.n600 VSUBS 0.007743f
C681 B.n601 VSUBS 0.007743f
C682 B.n602 VSUBS 0.007743f
C683 B.n603 VSUBS 0.007743f
C684 B.n604 VSUBS 0.007743f
C685 B.n605 VSUBS 0.007743f
C686 B.n606 VSUBS 0.007743f
C687 B.n607 VSUBS 0.007743f
C688 B.n608 VSUBS 0.007743f
C689 B.n609 VSUBS 0.007743f
C690 B.n610 VSUBS 0.007743f
C691 B.n611 VSUBS 0.007743f
C692 B.n612 VSUBS 0.007743f
C693 B.n613 VSUBS 0.007743f
C694 B.n614 VSUBS 0.007743f
C695 B.n615 VSUBS 0.007743f
C696 B.n616 VSUBS 0.007743f
C697 B.n617 VSUBS 0.007743f
C698 B.n618 VSUBS 0.007743f
C699 B.n619 VSUBS 0.007743f
C700 B.n620 VSUBS 0.007743f
C701 B.n621 VSUBS 0.007743f
C702 B.n622 VSUBS 0.007743f
C703 B.n623 VSUBS 0.007743f
C704 B.n624 VSUBS 0.007743f
C705 B.n625 VSUBS 0.007743f
C706 B.n626 VSUBS 0.007743f
C707 B.n627 VSUBS 0.007743f
C708 B.n628 VSUBS 0.007743f
C709 B.n629 VSUBS 0.007743f
C710 B.n630 VSUBS 0.007743f
C711 B.n631 VSUBS 0.007743f
C712 B.n632 VSUBS 0.007743f
C713 B.n633 VSUBS 0.007743f
C714 B.n634 VSUBS 0.007743f
C715 B.n635 VSUBS 0.007287f
C716 B.n636 VSUBS 0.017939f
C717 B.n637 VSUBS 0.004327f
C718 B.n638 VSUBS 0.007743f
C719 B.n639 VSUBS 0.007743f
C720 B.n640 VSUBS 0.007743f
C721 B.n641 VSUBS 0.007743f
C722 B.n642 VSUBS 0.007743f
C723 B.n643 VSUBS 0.007743f
C724 B.n644 VSUBS 0.007743f
C725 B.n645 VSUBS 0.007743f
C726 B.n646 VSUBS 0.007743f
C727 B.n647 VSUBS 0.007743f
C728 B.n648 VSUBS 0.007743f
C729 B.n649 VSUBS 0.007743f
C730 B.n650 VSUBS 0.004327f
C731 B.n651 VSUBS 0.007743f
C732 B.n652 VSUBS 0.007743f
C733 B.n653 VSUBS 0.007287f
C734 B.n654 VSUBS 0.007743f
C735 B.n655 VSUBS 0.007743f
C736 B.n656 VSUBS 0.007743f
C737 B.n657 VSUBS 0.007743f
C738 B.n658 VSUBS 0.007743f
C739 B.n659 VSUBS 0.007743f
C740 B.n660 VSUBS 0.007743f
C741 B.n661 VSUBS 0.007743f
C742 B.n662 VSUBS 0.007743f
C743 B.n663 VSUBS 0.007743f
C744 B.n664 VSUBS 0.007743f
C745 B.n665 VSUBS 0.007743f
C746 B.n666 VSUBS 0.007743f
C747 B.n667 VSUBS 0.007743f
C748 B.n668 VSUBS 0.007743f
C749 B.n669 VSUBS 0.007743f
C750 B.n670 VSUBS 0.007743f
C751 B.n671 VSUBS 0.007743f
C752 B.n672 VSUBS 0.007743f
C753 B.n673 VSUBS 0.007743f
C754 B.n674 VSUBS 0.007743f
C755 B.n675 VSUBS 0.007743f
C756 B.n676 VSUBS 0.007743f
C757 B.n677 VSUBS 0.007743f
C758 B.n678 VSUBS 0.007743f
C759 B.n679 VSUBS 0.007743f
C760 B.n680 VSUBS 0.007743f
C761 B.n681 VSUBS 0.007743f
C762 B.n682 VSUBS 0.007743f
C763 B.n683 VSUBS 0.007743f
C764 B.n684 VSUBS 0.007743f
C765 B.n685 VSUBS 0.007743f
C766 B.n686 VSUBS 0.007743f
C767 B.n687 VSUBS 0.007743f
C768 B.n688 VSUBS 0.007743f
C769 B.n689 VSUBS 0.007743f
C770 B.n690 VSUBS 0.007743f
C771 B.n691 VSUBS 0.007743f
C772 B.n692 VSUBS 0.007743f
C773 B.n693 VSUBS 0.007743f
C774 B.n694 VSUBS 0.007743f
C775 B.n695 VSUBS 0.007743f
C776 B.n696 VSUBS 0.007743f
C777 B.n697 VSUBS 0.007743f
C778 B.n698 VSUBS 0.007743f
C779 B.n699 VSUBS 0.007743f
C780 B.n700 VSUBS 0.007743f
C781 B.n701 VSUBS 0.007743f
C782 B.n702 VSUBS 0.007743f
C783 B.n703 VSUBS 0.007743f
C784 B.n704 VSUBS 0.007743f
C785 B.n705 VSUBS 0.007743f
C786 B.n706 VSUBS 0.007743f
C787 B.n707 VSUBS 0.007743f
C788 B.n708 VSUBS 0.007743f
C789 B.n709 VSUBS 0.007743f
C790 B.n710 VSUBS 0.007743f
C791 B.n711 VSUBS 0.007743f
C792 B.n712 VSUBS 0.007743f
C793 B.n713 VSUBS 0.007743f
C794 B.n714 VSUBS 0.007743f
C795 B.n715 VSUBS 0.007743f
C796 B.n716 VSUBS 0.007743f
C797 B.n717 VSUBS 0.007743f
C798 B.n718 VSUBS 0.007743f
C799 B.n719 VSUBS 0.007743f
C800 B.n720 VSUBS 0.007743f
C801 B.n721 VSUBS 0.007743f
C802 B.n722 VSUBS 0.007743f
C803 B.n723 VSUBS 0.007743f
C804 B.n724 VSUBS 0.007743f
C805 B.n725 VSUBS 0.007743f
C806 B.n726 VSUBS 0.007743f
C807 B.n727 VSUBS 0.007743f
C808 B.n728 VSUBS 0.007743f
C809 B.n729 VSUBS 0.007743f
C810 B.n730 VSUBS 0.007743f
C811 B.n731 VSUBS 0.007743f
C812 B.n732 VSUBS 0.007743f
C813 B.n733 VSUBS 0.007743f
C814 B.n734 VSUBS 0.007743f
C815 B.n735 VSUBS 0.007743f
C816 B.n736 VSUBS 0.007743f
C817 B.n737 VSUBS 0.007743f
C818 B.n738 VSUBS 0.007743f
C819 B.n739 VSUBS 0.019046f
C820 B.n740 VSUBS 0.019046f
C821 B.n741 VSUBS 0.0183f
C822 B.n742 VSUBS 0.007743f
C823 B.n743 VSUBS 0.007743f
C824 B.n744 VSUBS 0.007743f
C825 B.n745 VSUBS 0.007743f
C826 B.n746 VSUBS 0.007743f
C827 B.n747 VSUBS 0.007743f
C828 B.n748 VSUBS 0.007743f
C829 B.n749 VSUBS 0.007743f
C830 B.n750 VSUBS 0.007743f
C831 B.n751 VSUBS 0.007743f
C832 B.n752 VSUBS 0.007743f
C833 B.n753 VSUBS 0.007743f
C834 B.n754 VSUBS 0.007743f
C835 B.n755 VSUBS 0.007743f
C836 B.n756 VSUBS 0.007743f
C837 B.n757 VSUBS 0.007743f
C838 B.n758 VSUBS 0.007743f
C839 B.n759 VSUBS 0.007743f
C840 B.n760 VSUBS 0.007743f
C841 B.n761 VSUBS 0.007743f
C842 B.n762 VSUBS 0.007743f
C843 B.n763 VSUBS 0.007743f
C844 B.n764 VSUBS 0.007743f
C845 B.n765 VSUBS 0.007743f
C846 B.n766 VSUBS 0.007743f
C847 B.n767 VSUBS 0.007743f
C848 B.n768 VSUBS 0.007743f
C849 B.n769 VSUBS 0.007743f
C850 B.n770 VSUBS 0.007743f
C851 B.n771 VSUBS 0.007743f
C852 B.n772 VSUBS 0.007743f
C853 B.n773 VSUBS 0.007743f
C854 B.n774 VSUBS 0.007743f
C855 B.n775 VSUBS 0.007743f
C856 B.n776 VSUBS 0.007743f
C857 B.n777 VSUBS 0.007743f
C858 B.n778 VSUBS 0.007743f
C859 B.n779 VSUBS 0.007743f
C860 B.n780 VSUBS 0.007743f
C861 B.n781 VSUBS 0.007743f
C862 B.n782 VSUBS 0.007743f
C863 B.n783 VSUBS 0.007743f
C864 B.n784 VSUBS 0.007743f
C865 B.n785 VSUBS 0.007743f
C866 B.n786 VSUBS 0.007743f
C867 B.n787 VSUBS 0.007743f
C868 B.n788 VSUBS 0.007743f
C869 B.n789 VSUBS 0.007743f
C870 B.n790 VSUBS 0.007743f
C871 B.n791 VSUBS 0.017532f
C872 VDD1.t2 VSUBS 4.13129f
C873 VDD1.t5 VSUBS 4.13001f
C874 VDD1.t4 VSUBS 0.380528f
C875 VDD1.t3 VSUBS 0.380528f
C876 VDD1.n0 VSUBS 3.17748f
C877 VDD1.n1 VSUBS 3.85606f
C878 VDD1.t0 VSUBS 0.380528f
C879 VDD1.t1 VSUBS 0.380528f
C880 VDD1.n2 VSUBS 3.17346f
C881 VDD1.n3 VSUBS 3.52314f
C882 VTAIL.t3 VSUBS 0.387184f
C883 VTAIL.t5 VSUBS 0.387184f
C884 VTAIL.n0 VSUBS 3.07122f
C885 VTAIL.n1 VSUBS 0.811476f
C886 VTAIL.t11 VSUBS 4.00817f
C887 VTAIL.n2 VSUBS 1.04547f
C888 VTAIL.t6 VSUBS 0.387184f
C889 VTAIL.t7 VSUBS 0.387184f
C890 VTAIL.n3 VSUBS 3.07122f
C891 VTAIL.n4 VSUBS 2.85584f
C892 VTAIL.t1 VSUBS 0.387184f
C893 VTAIL.t4 VSUBS 0.387184f
C894 VTAIL.n5 VSUBS 3.07122f
C895 VTAIL.n6 VSUBS 2.85583f
C896 VTAIL.t2 VSUBS 4.00818f
C897 VTAIL.n7 VSUBS 1.04546f
C898 VTAIL.t8 VSUBS 0.387184f
C899 VTAIL.t9 VSUBS 0.387184f
C900 VTAIL.n8 VSUBS 3.07122f
C901 VTAIL.n9 VSUBS 0.926461f
C902 VTAIL.t10 VSUBS 4.00817f
C903 VTAIL.n10 VSUBS 2.81472f
C904 VTAIL.t0 VSUBS 4.00817f
C905 VTAIL.n11 VSUBS 2.76959f
C906 VP.n0 VSUBS 0.034588f
C907 VP.t2 VSUBS 3.06881f
C908 VP.n1 VSUBS 0.029556f
C909 VP.n2 VSUBS 0.034588f
C910 VP.t1 VSUBS 3.06881f
C911 VP.n3 VSUBS 0.029556f
C912 VP.n4 VSUBS 0.034588f
C913 VP.t0 VSUBS 3.06881f
C914 VP.n5 VSUBS 0.034588f
C915 VP.t4 VSUBS 3.06881f
C916 VP.n6 VSUBS 0.029556f
C917 VP.t3 VSUBS 3.22868f
C918 VP.n7 VSUBS 1.14646f
C919 VP.t5 VSUBS 3.06881f
C920 VP.n8 VSUBS 1.16667f
C921 VP.n9 VSUBS 0.069515f
C922 VP.n10 VSUBS 0.255541f
C923 VP.n11 VSUBS 0.034588f
C924 VP.n12 VSUBS 0.034588f
C925 VP.n13 VSUBS 0.065629f
C926 VP.n14 VSUBS 0.040076f
C927 VP.n15 VSUBS 1.15463f
C928 VP.n16 VSUBS 1.88938f
C929 VP.n17 VSUBS 1.91432f
C930 VP.n18 VSUBS 1.15463f
C931 VP.n19 VSUBS 0.040076f
C932 VP.n20 VSUBS 0.065629f
C933 VP.n21 VSUBS 0.034588f
C934 VP.n22 VSUBS 0.034588f
C935 VP.n23 VSUBS 0.034588f
C936 VP.n24 VSUBS 0.069515f
C937 VP.n25 VSUBS 1.10636f
C938 VP.n26 VSUBS 0.069515f
C939 VP.n27 VSUBS 0.034588f
C940 VP.n28 VSUBS 0.034588f
C941 VP.n29 VSUBS 0.034588f
C942 VP.n30 VSUBS 0.065629f
C943 VP.n31 VSUBS 0.040076f
C944 VP.n32 VSUBS 1.15463f
C945 VP.n33 VSUBS 0.036161f
.ends

