* NGSPICE file created from diff_pair_sample_0019.ext - technology: sky130A

.subckt diff_pair_sample_0019 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.1
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.1
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.1
X3 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.1
X4 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.1
X5 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.1
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.1
X7 VTAIL.t6 VN.t1 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.1
X8 VDD2.t2 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.1
X9 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.1
X10 VDD2.t0 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.1
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.1
R0 VN.n1 VN.t3 113.725
R1 VN.n0 VN.t1 113.725
R2 VN.n0 VN.t2 112.71
R3 VN.n1 VN.t0 112.71
R4 VN VN.n1 49.5666
R5 VN VN.n0 2.82039
R6 VDD2.n2 VDD2.n0 108.269
R7 VDD2.n2 VDD2.n1 66.9068
R8 VDD2.n1 VDD2.t1 1.94549
R9 VDD2.n1 VDD2.t0 1.94549
R10 VDD2.n0 VDD2.t3 1.94549
R11 VDD2.n0 VDD2.t2 1.94549
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n426 VTAIL.n378 289.615
R14 VTAIL.n48 VTAIL.n0 289.615
R15 VTAIL.n102 VTAIL.n54 289.615
R16 VTAIL.n156 VTAIL.n108 289.615
R17 VTAIL.n372 VTAIL.n324 289.615
R18 VTAIL.n318 VTAIL.n270 289.615
R19 VTAIL.n264 VTAIL.n216 289.615
R20 VTAIL.n210 VTAIL.n162 289.615
R21 VTAIL.n394 VTAIL.n393 185
R22 VTAIL.n399 VTAIL.n398 185
R23 VTAIL.n401 VTAIL.n400 185
R24 VTAIL.n390 VTAIL.n389 185
R25 VTAIL.n407 VTAIL.n406 185
R26 VTAIL.n409 VTAIL.n408 185
R27 VTAIL.n386 VTAIL.n385 185
R28 VTAIL.n416 VTAIL.n415 185
R29 VTAIL.n417 VTAIL.n384 185
R30 VTAIL.n419 VTAIL.n418 185
R31 VTAIL.n382 VTAIL.n381 185
R32 VTAIL.n425 VTAIL.n424 185
R33 VTAIL.n427 VTAIL.n426 185
R34 VTAIL.n16 VTAIL.n15 185
R35 VTAIL.n21 VTAIL.n20 185
R36 VTAIL.n23 VTAIL.n22 185
R37 VTAIL.n12 VTAIL.n11 185
R38 VTAIL.n29 VTAIL.n28 185
R39 VTAIL.n31 VTAIL.n30 185
R40 VTAIL.n8 VTAIL.n7 185
R41 VTAIL.n38 VTAIL.n37 185
R42 VTAIL.n39 VTAIL.n6 185
R43 VTAIL.n41 VTAIL.n40 185
R44 VTAIL.n4 VTAIL.n3 185
R45 VTAIL.n47 VTAIL.n46 185
R46 VTAIL.n49 VTAIL.n48 185
R47 VTAIL.n70 VTAIL.n69 185
R48 VTAIL.n75 VTAIL.n74 185
R49 VTAIL.n77 VTAIL.n76 185
R50 VTAIL.n66 VTAIL.n65 185
R51 VTAIL.n83 VTAIL.n82 185
R52 VTAIL.n85 VTAIL.n84 185
R53 VTAIL.n62 VTAIL.n61 185
R54 VTAIL.n92 VTAIL.n91 185
R55 VTAIL.n93 VTAIL.n60 185
R56 VTAIL.n95 VTAIL.n94 185
R57 VTAIL.n58 VTAIL.n57 185
R58 VTAIL.n101 VTAIL.n100 185
R59 VTAIL.n103 VTAIL.n102 185
R60 VTAIL.n124 VTAIL.n123 185
R61 VTAIL.n129 VTAIL.n128 185
R62 VTAIL.n131 VTAIL.n130 185
R63 VTAIL.n120 VTAIL.n119 185
R64 VTAIL.n137 VTAIL.n136 185
R65 VTAIL.n139 VTAIL.n138 185
R66 VTAIL.n116 VTAIL.n115 185
R67 VTAIL.n146 VTAIL.n145 185
R68 VTAIL.n147 VTAIL.n114 185
R69 VTAIL.n149 VTAIL.n148 185
R70 VTAIL.n112 VTAIL.n111 185
R71 VTAIL.n155 VTAIL.n154 185
R72 VTAIL.n157 VTAIL.n156 185
R73 VTAIL.n373 VTAIL.n372 185
R74 VTAIL.n371 VTAIL.n370 185
R75 VTAIL.n328 VTAIL.n327 185
R76 VTAIL.n365 VTAIL.n364 185
R77 VTAIL.n363 VTAIL.n330 185
R78 VTAIL.n362 VTAIL.n361 185
R79 VTAIL.n333 VTAIL.n331 185
R80 VTAIL.n356 VTAIL.n355 185
R81 VTAIL.n354 VTAIL.n353 185
R82 VTAIL.n337 VTAIL.n336 185
R83 VTAIL.n348 VTAIL.n347 185
R84 VTAIL.n346 VTAIL.n345 185
R85 VTAIL.n341 VTAIL.n340 185
R86 VTAIL.n319 VTAIL.n318 185
R87 VTAIL.n317 VTAIL.n316 185
R88 VTAIL.n274 VTAIL.n273 185
R89 VTAIL.n311 VTAIL.n310 185
R90 VTAIL.n309 VTAIL.n276 185
R91 VTAIL.n308 VTAIL.n307 185
R92 VTAIL.n279 VTAIL.n277 185
R93 VTAIL.n302 VTAIL.n301 185
R94 VTAIL.n300 VTAIL.n299 185
R95 VTAIL.n283 VTAIL.n282 185
R96 VTAIL.n294 VTAIL.n293 185
R97 VTAIL.n292 VTAIL.n291 185
R98 VTAIL.n287 VTAIL.n286 185
R99 VTAIL.n265 VTAIL.n264 185
R100 VTAIL.n263 VTAIL.n262 185
R101 VTAIL.n220 VTAIL.n219 185
R102 VTAIL.n257 VTAIL.n256 185
R103 VTAIL.n255 VTAIL.n222 185
R104 VTAIL.n254 VTAIL.n253 185
R105 VTAIL.n225 VTAIL.n223 185
R106 VTAIL.n248 VTAIL.n247 185
R107 VTAIL.n246 VTAIL.n245 185
R108 VTAIL.n229 VTAIL.n228 185
R109 VTAIL.n240 VTAIL.n239 185
R110 VTAIL.n238 VTAIL.n237 185
R111 VTAIL.n233 VTAIL.n232 185
R112 VTAIL.n211 VTAIL.n210 185
R113 VTAIL.n209 VTAIL.n208 185
R114 VTAIL.n166 VTAIL.n165 185
R115 VTAIL.n203 VTAIL.n202 185
R116 VTAIL.n201 VTAIL.n168 185
R117 VTAIL.n200 VTAIL.n199 185
R118 VTAIL.n171 VTAIL.n169 185
R119 VTAIL.n194 VTAIL.n193 185
R120 VTAIL.n192 VTAIL.n191 185
R121 VTAIL.n175 VTAIL.n174 185
R122 VTAIL.n186 VTAIL.n185 185
R123 VTAIL.n184 VTAIL.n183 185
R124 VTAIL.n179 VTAIL.n178 185
R125 VTAIL.n395 VTAIL.t5 149.524
R126 VTAIL.n17 VTAIL.t6 149.524
R127 VTAIL.n71 VTAIL.t2 149.524
R128 VTAIL.n125 VTAIL.t1 149.524
R129 VTAIL.n342 VTAIL.t0 149.524
R130 VTAIL.n288 VTAIL.t3 149.524
R131 VTAIL.n234 VTAIL.t4 149.524
R132 VTAIL.n180 VTAIL.t7 149.524
R133 VTAIL.n399 VTAIL.n393 104.615
R134 VTAIL.n400 VTAIL.n399 104.615
R135 VTAIL.n400 VTAIL.n389 104.615
R136 VTAIL.n407 VTAIL.n389 104.615
R137 VTAIL.n408 VTAIL.n407 104.615
R138 VTAIL.n408 VTAIL.n385 104.615
R139 VTAIL.n416 VTAIL.n385 104.615
R140 VTAIL.n417 VTAIL.n416 104.615
R141 VTAIL.n418 VTAIL.n417 104.615
R142 VTAIL.n418 VTAIL.n381 104.615
R143 VTAIL.n425 VTAIL.n381 104.615
R144 VTAIL.n426 VTAIL.n425 104.615
R145 VTAIL.n21 VTAIL.n15 104.615
R146 VTAIL.n22 VTAIL.n21 104.615
R147 VTAIL.n22 VTAIL.n11 104.615
R148 VTAIL.n29 VTAIL.n11 104.615
R149 VTAIL.n30 VTAIL.n29 104.615
R150 VTAIL.n30 VTAIL.n7 104.615
R151 VTAIL.n38 VTAIL.n7 104.615
R152 VTAIL.n39 VTAIL.n38 104.615
R153 VTAIL.n40 VTAIL.n39 104.615
R154 VTAIL.n40 VTAIL.n3 104.615
R155 VTAIL.n47 VTAIL.n3 104.615
R156 VTAIL.n48 VTAIL.n47 104.615
R157 VTAIL.n75 VTAIL.n69 104.615
R158 VTAIL.n76 VTAIL.n75 104.615
R159 VTAIL.n76 VTAIL.n65 104.615
R160 VTAIL.n83 VTAIL.n65 104.615
R161 VTAIL.n84 VTAIL.n83 104.615
R162 VTAIL.n84 VTAIL.n61 104.615
R163 VTAIL.n92 VTAIL.n61 104.615
R164 VTAIL.n93 VTAIL.n92 104.615
R165 VTAIL.n94 VTAIL.n93 104.615
R166 VTAIL.n94 VTAIL.n57 104.615
R167 VTAIL.n101 VTAIL.n57 104.615
R168 VTAIL.n102 VTAIL.n101 104.615
R169 VTAIL.n129 VTAIL.n123 104.615
R170 VTAIL.n130 VTAIL.n129 104.615
R171 VTAIL.n130 VTAIL.n119 104.615
R172 VTAIL.n137 VTAIL.n119 104.615
R173 VTAIL.n138 VTAIL.n137 104.615
R174 VTAIL.n138 VTAIL.n115 104.615
R175 VTAIL.n146 VTAIL.n115 104.615
R176 VTAIL.n147 VTAIL.n146 104.615
R177 VTAIL.n148 VTAIL.n147 104.615
R178 VTAIL.n148 VTAIL.n111 104.615
R179 VTAIL.n155 VTAIL.n111 104.615
R180 VTAIL.n156 VTAIL.n155 104.615
R181 VTAIL.n372 VTAIL.n371 104.615
R182 VTAIL.n371 VTAIL.n327 104.615
R183 VTAIL.n364 VTAIL.n327 104.615
R184 VTAIL.n364 VTAIL.n363 104.615
R185 VTAIL.n363 VTAIL.n362 104.615
R186 VTAIL.n362 VTAIL.n331 104.615
R187 VTAIL.n355 VTAIL.n331 104.615
R188 VTAIL.n355 VTAIL.n354 104.615
R189 VTAIL.n354 VTAIL.n336 104.615
R190 VTAIL.n347 VTAIL.n336 104.615
R191 VTAIL.n347 VTAIL.n346 104.615
R192 VTAIL.n346 VTAIL.n340 104.615
R193 VTAIL.n318 VTAIL.n317 104.615
R194 VTAIL.n317 VTAIL.n273 104.615
R195 VTAIL.n310 VTAIL.n273 104.615
R196 VTAIL.n310 VTAIL.n309 104.615
R197 VTAIL.n309 VTAIL.n308 104.615
R198 VTAIL.n308 VTAIL.n277 104.615
R199 VTAIL.n301 VTAIL.n277 104.615
R200 VTAIL.n301 VTAIL.n300 104.615
R201 VTAIL.n300 VTAIL.n282 104.615
R202 VTAIL.n293 VTAIL.n282 104.615
R203 VTAIL.n293 VTAIL.n292 104.615
R204 VTAIL.n292 VTAIL.n286 104.615
R205 VTAIL.n264 VTAIL.n263 104.615
R206 VTAIL.n263 VTAIL.n219 104.615
R207 VTAIL.n256 VTAIL.n219 104.615
R208 VTAIL.n256 VTAIL.n255 104.615
R209 VTAIL.n255 VTAIL.n254 104.615
R210 VTAIL.n254 VTAIL.n223 104.615
R211 VTAIL.n247 VTAIL.n223 104.615
R212 VTAIL.n247 VTAIL.n246 104.615
R213 VTAIL.n246 VTAIL.n228 104.615
R214 VTAIL.n239 VTAIL.n228 104.615
R215 VTAIL.n239 VTAIL.n238 104.615
R216 VTAIL.n238 VTAIL.n232 104.615
R217 VTAIL.n210 VTAIL.n209 104.615
R218 VTAIL.n209 VTAIL.n165 104.615
R219 VTAIL.n202 VTAIL.n165 104.615
R220 VTAIL.n202 VTAIL.n201 104.615
R221 VTAIL.n201 VTAIL.n200 104.615
R222 VTAIL.n200 VTAIL.n169 104.615
R223 VTAIL.n193 VTAIL.n169 104.615
R224 VTAIL.n193 VTAIL.n192 104.615
R225 VTAIL.n192 VTAIL.n174 104.615
R226 VTAIL.n185 VTAIL.n174 104.615
R227 VTAIL.n185 VTAIL.n184 104.615
R228 VTAIL.n184 VTAIL.n178 104.615
R229 VTAIL.t5 VTAIL.n393 52.3082
R230 VTAIL.t6 VTAIL.n15 52.3082
R231 VTAIL.t2 VTAIL.n69 52.3082
R232 VTAIL.t1 VTAIL.n123 52.3082
R233 VTAIL.t0 VTAIL.n340 52.3082
R234 VTAIL.t3 VTAIL.n286 52.3082
R235 VTAIL.t4 VTAIL.n232 52.3082
R236 VTAIL.t7 VTAIL.n178 52.3082
R237 VTAIL.n431 VTAIL.n430 36.452
R238 VTAIL.n53 VTAIL.n52 36.452
R239 VTAIL.n107 VTAIL.n106 36.452
R240 VTAIL.n161 VTAIL.n160 36.452
R241 VTAIL.n377 VTAIL.n376 36.452
R242 VTAIL.n323 VTAIL.n322 36.452
R243 VTAIL.n269 VTAIL.n268 36.452
R244 VTAIL.n215 VTAIL.n214 36.452
R245 VTAIL.n431 VTAIL.n377 24.0996
R246 VTAIL.n215 VTAIL.n161 24.0996
R247 VTAIL.n419 VTAIL.n384 13.1884
R248 VTAIL.n41 VTAIL.n6 13.1884
R249 VTAIL.n95 VTAIL.n60 13.1884
R250 VTAIL.n149 VTAIL.n114 13.1884
R251 VTAIL.n365 VTAIL.n330 13.1884
R252 VTAIL.n311 VTAIL.n276 13.1884
R253 VTAIL.n257 VTAIL.n222 13.1884
R254 VTAIL.n203 VTAIL.n168 13.1884
R255 VTAIL.n415 VTAIL.n414 12.8005
R256 VTAIL.n420 VTAIL.n382 12.8005
R257 VTAIL.n37 VTAIL.n36 12.8005
R258 VTAIL.n42 VTAIL.n4 12.8005
R259 VTAIL.n91 VTAIL.n90 12.8005
R260 VTAIL.n96 VTAIL.n58 12.8005
R261 VTAIL.n145 VTAIL.n144 12.8005
R262 VTAIL.n150 VTAIL.n112 12.8005
R263 VTAIL.n366 VTAIL.n328 12.8005
R264 VTAIL.n361 VTAIL.n332 12.8005
R265 VTAIL.n312 VTAIL.n274 12.8005
R266 VTAIL.n307 VTAIL.n278 12.8005
R267 VTAIL.n258 VTAIL.n220 12.8005
R268 VTAIL.n253 VTAIL.n224 12.8005
R269 VTAIL.n204 VTAIL.n166 12.8005
R270 VTAIL.n199 VTAIL.n170 12.8005
R271 VTAIL.n413 VTAIL.n386 12.0247
R272 VTAIL.n424 VTAIL.n423 12.0247
R273 VTAIL.n35 VTAIL.n8 12.0247
R274 VTAIL.n46 VTAIL.n45 12.0247
R275 VTAIL.n89 VTAIL.n62 12.0247
R276 VTAIL.n100 VTAIL.n99 12.0247
R277 VTAIL.n143 VTAIL.n116 12.0247
R278 VTAIL.n154 VTAIL.n153 12.0247
R279 VTAIL.n370 VTAIL.n369 12.0247
R280 VTAIL.n360 VTAIL.n333 12.0247
R281 VTAIL.n316 VTAIL.n315 12.0247
R282 VTAIL.n306 VTAIL.n279 12.0247
R283 VTAIL.n262 VTAIL.n261 12.0247
R284 VTAIL.n252 VTAIL.n225 12.0247
R285 VTAIL.n208 VTAIL.n207 12.0247
R286 VTAIL.n198 VTAIL.n171 12.0247
R287 VTAIL.n410 VTAIL.n409 11.249
R288 VTAIL.n427 VTAIL.n380 11.249
R289 VTAIL.n32 VTAIL.n31 11.249
R290 VTAIL.n49 VTAIL.n2 11.249
R291 VTAIL.n86 VTAIL.n85 11.249
R292 VTAIL.n103 VTAIL.n56 11.249
R293 VTAIL.n140 VTAIL.n139 11.249
R294 VTAIL.n157 VTAIL.n110 11.249
R295 VTAIL.n373 VTAIL.n326 11.249
R296 VTAIL.n357 VTAIL.n356 11.249
R297 VTAIL.n319 VTAIL.n272 11.249
R298 VTAIL.n303 VTAIL.n302 11.249
R299 VTAIL.n265 VTAIL.n218 11.249
R300 VTAIL.n249 VTAIL.n248 11.249
R301 VTAIL.n211 VTAIL.n164 11.249
R302 VTAIL.n195 VTAIL.n194 11.249
R303 VTAIL.n406 VTAIL.n388 10.4732
R304 VTAIL.n428 VTAIL.n378 10.4732
R305 VTAIL.n28 VTAIL.n10 10.4732
R306 VTAIL.n50 VTAIL.n0 10.4732
R307 VTAIL.n82 VTAIL.n64 10.4732
R308 VTAIL.n104 VTAIL.n54 10.4732
R309 VTAIL.n136 VTAIL.n118 10.4732
R310 VTAIL.n158 VTAIL.n108 10.4732
R311 VTAIL.n374 VTAIL.n324 10.4732
R312 VTAIL.n353 VTAIL.n335 10.4732
R313 VTAIL.n320 VTAIL.n270 10.4732
R314 VTAIL.n299 VTAIL.n281 10.4732
R315 VTAIL.n266 VTAIL.n216 10.4732
R316 VTAIL.n245 VTAIL.n227 10.4732
R317 VTAIL.n212 VTAIL.n162 10.4732
R318 VTAIL.n191 VTAIL.n173 10.4732
R319 VTAIL.n395 VTAIL.n394 10.2747
R320 VTAIL.n17 VTAIL.n16 10.2747
R321 VTAIL.n71 VTAIL.n70 10.2747
R322 VTAIL.n125 VTAIL.n124 10.2747
R323 VTAIL.n342 VTAIL.n341 10.2747
R324 VTAIL.n288 VTAIL.n287 10.2747
R325 VTAIL.n234 VTAIL.n233 10.2747
R326 VTAIL.n180 VTAIL.n179 10.2747
R327 VTAIL.n405 VTAIL.n390 9.69747
R328 VTAIL.n27 VTAIL.n12 9.69747
R329 VTAIL.n81 VTAIL.n66 9.69747
R330 VTAIL.n135 VTAIL.n120 9.69747
R331 VTAIL.n352 VTAIL.n337 9.69747
R332 VTAIL.n298 VTAIL.n283 9.69747
R333 VTAIL.n244 VTAIL.n229 9.69747
R334 VTAIL.n190 VTAIL.n175 9.69747
R335 VTAIL.n430 VTAIL.n429 9.45567
R336 VTAIL.n52 VTAIL.n51 9.45567
R337 VTAIL.n106 VTAIL.n105 9.45567
R338 VTAIL.n160 VTAIL.n159 9.45567
R339 VTAIL.n376 VTAIL.n375 9.45567
R340 VTAIL.n322 VTAIL.n321 9.45567
R341 VTAIL.n268 VTAIL.n267 9.45567
R342 VTAIL.n214 VTAIL.n213 9.45567
R343 VTAIL.n429 VTAIL.n428 9.3005
R344 VTAIL.n380 VTAIL.n379 9.3005
R345 VTAIL.n423 VTAIL.n422 9.3005
R346 VTAIL.n421 VTAIL.n420 9.3005
R347 VTAIL.n397 VTAIL.n396 9.3005
R348 VTAIL.n392 VTAIL.n391 9.3005
R349 VTAIL.n403 VTAIL.n402 9.3005
R350 VTAIL.n405 VTAIL.n404 9.3005
R351 VTAIL.n388 VTAIL.n387 9.3005
R352 VTAIL.n411 VTAIL.n410 9.3005
R353 VTAIL.n413 VTAIL.n412 9.3005
R354 VTAIL.n414 VTAIL.n383 9.3005
R355 VTAIL.n51 VTAIL.n50 9.3005
R356 VTAIL.n2 VTAIL.n1 9.3005
R357 VTAIL.n45 VTAIL.n44 9.3005
R358 VTAIL.n43 VTAIL.n42 9.3005
R359 VTAIL.n19 VTAIL.n18 9.3005
R360 VTAIL.n14 VTAIL.n13 9.3005
R361 VTAIL.n25 VTAIL.n24 9.3005
R362 VTAIL.n27 VTAIL.n26 9.3005
R363 VTAIL.n10 VTAIL.n9 9.3005
R364 VTAIL.n33 VTAIL.n32 9.3005
R365 VTAIL.n35 VTAIL.n34 9.3005
R366 VTAIL.n36 VTAIL.n5 9.3005
R367 VTAIL.n105 VTAIL.n104 9.3005
R368 VTAIL.n56 VTAIL.n55 9.3005
R369 VTAIL.n99 VTAIL.n98 9.3005
R370 VTAIL.n97 VTAIL.n96 9.3005
R371 VTAIL.n73 VTAIL.n72 9.3005
R372 VTAIL.n68 VTAIL.n67 9.3005
R373 VTAIL.n79 VTAIL.n78 9.3005
R374 VTAIL.n81 VTAIL.n80 9.3005
R375 VTAIL.n64 VTAIL.n63 9.3005
R376 VTAIL.n87 VTAIL.n86 9.3005
R377 VTAIL.n89 VTAIL.n88 9.3005
R378 VTAIL.n90 VTAIL.n59 9.3005
R379 VTAIL.n159 VTAIL.n158 9.3005
R380 VTAIL.n110 VTAIL.n109 9.3005
R381 VTAIL.n153 VTAIL.n152 9.3005
R382 VTAIL.n151 VTAIL.n150 9.3005
R383 VTAIL.n127 VTAIL.n126 9.3005
R384 VTAIL.n122 VTAIL.n121 9.3005
R385 VTAIL.n133 VTAIL.n132 9.3005
R386 VTAIL.n135 VTAIL.n134 9.3005
R387 VTAIL.n118 VTAIL.n117 9.3005
R388 VTAIL.n141 VTAIL.n140 9.3005
R389 VTAIL.n143 VTAIL.n142 9.3005
R390 VTAIL.n144 VTAIL.n113 9.3005
R391 VTAIL.n344 VTAIL.n343 9.3005
R392 VTAIL.n339 VTAIL.n338 9.3005
R393 VTAIL.n350 VTAIL.n349 9.3005
R394 VTAIL.n352 VTAIL.n351 9.3005
R395 VTAIL.n335 VTAIL.n334 9.3005
R396 VTAIL.n358 VTAIL.n357 9.3005
R397 VTAIL.n360 VTAIL.n359 9.3005
R398 VTAIL.n332 VTAIL.n329 9.3005
R399 VTAIL.n375 VTAIL.n374 9.3005
R400 VTAIL.n326 VTAIL.n325 9.3005
R401 VTAIL.n369 VTAIL.n368 9.3005
R402 VTAIL.n367 VTAIL.n366 9.3005
R403 VTAIL.n290 VTAIL.n289 9.3005
R404 VTAIL.n285 VTAIL.n284 9.3005
R405 VTAIL.n296 VTAIL.n295 9.3005
R406 VTAIL.n298 VTAIL.n297 9.3005
R407 VTAIL.n281 VTAIL.n280 9.3005
R408 VTAIL.n304 VTAIL.n303 9.3005
R409 VTAIL.n306 VTAIL.n305 9.3005
R410 VTAIL.n278 VTAIL.n275 9.3005
R411 VTAIL.n321 VTAIL.n320 9.3005
R412 VTAIL.n272 VTAIL.n271 9.3005
R413 VTAIL.n315 VTAIL.n314 9.3005
R414 VTAIL.n313 VTAIL.n312 9.3005
R415 VTAIL.n236 VTAIL.n235 9.3005
R416 VTAIL.n231 VTAIL.n230 9.3005
R417 VTAIL.n242 VTAIL.n241 9.3005
R418 VTAIL.n244 VTAIL.n243 9.3005
R419 VTAIL.n227 VTAIL.n226 9.3005
R420 VTAIL.n250 VTAIL.n249 9.3005
R421 VTAIL.n252 VTAIL.n251 9.3005
R422 VTAIL.n224 VTAIL.n221 9.3005
R423 VTAIL.n267 VTAIL.n266 9.3005
R424 VTAIL.n218 VTAIL.n217 9.3005
R425 VTAIL.n261 VTAIL.n260 9.3005
R426 VTAIL.n259 VTAIL.n258 9.3005
R427 VTAIL.n182 VTAIL.n181 9.3005
R428 VTAIL.n177 VTAIL.n176 9.3005
R429 VTAIL.n188 VTAIL.n187 9.3005
R430 VTAIL.n190 VTAIL.n189 9.3005
R431 VTAIL.n173 VTAIL.n172 9.3005
R432 VTAIL.n196 VTAIL.n195 9.3005
R433 VTAIL.n198 VTAIL.n197 9.3005
R434 VTAIL.n170 VTAIL.n167 9.3005
R435 VTAIL.n213 VTAIL.n212 9.3005
R436 VTAIL.n164 VTAIL.n163 9.3005
R437 VTAIL.n207 VTAIL.n206 9.3005
R438 VTAIL.n205 VTAIL.n204 9.3005
R439 VTAIL.n402 VTAIL.n401 8.92171
R440 VTAIL.n24 VTAIL.n23 8.92171
R441 VTAIL.n78 VTAIL.n77 8.92171
R442 VTAIL.n132 VTAIL.n131 8.92171
R443 VTAIL.n349 VTAIL.n348 8.92171
R444 VTAIL.n295 VTAIL.n294 8.92171
R445 VTAIL.n241 VTAIL.n240 8.92171
R446 VTAIL.n187 VTAIL.n186 8.92171
R447 VTAIL.n398 VTAIL.n392 8.14595
R448 VTAIL.n20 VTAIL.n14 8.14595
R449 VTAIL.n74 VTAIL.n68 8.14595
R450 VTAIL.n128 VTAIL.n122 8.14595
R451 VTAIL.n345 VTAIL.n339 8.14595
R452 VTAIL.n291 VTAIL.n285 8.14595
R453 VTAIL.n237 VTAIL.n231 8.14595
R454 VTAIL.n183 VTAIL.n177 8.14595
R455 VTAIL.n397 VTAIL.n394 7.3702
R456 VTAIL.n19 VTAIL.n16 7.3702
R457 VTAIL.n73 VTAIL.n70 7.3702
R458 VTAIL.n127 VTAIL.n124 7.3702
R459 VTAIL.n344 VTAIL.n341 7.3702
R460 VTAIL.n290 VTAIL.n287 7.3702
R461 VTAIL.n236 VTAIL.n233 7.3702
R462 VTAIL.n182 VTAIL.n179 7.3702
R463 VTAIL.n398 VTAIL.n397 5.81868
R464 VTAIL.n20 VTAIL.n19 5.81868
R465 VTAIL.n74 VTAIL.n73 5.81868
R466 VTAIL.n128 VTAIL.n127 5.81868
R467 VTAIL.n345 VTAIL.n344 5.81868
R468 VTAIL.n291 VTAIL.n290 5.81868
R469 VTAIL.n237 VTAIL.n236 5.81868
R470 VTAIL.n183 VTAIL.n182 5.81868
R471 VTAIL.n401 VTAIL.n392 5.04292
R472 VTAIL.n23 VTAIL.n14 5.04292
R473 VTAIL.n77 VTAIL.n68 5.04292
R474 VTAIL.n131 VTAIL.n122 5.04292
R475 VTAIL.n348 VTAIL.n339 5.04292
R476 VTAIL.n294 VTAIL.n285 5.04292
R477 VTAIL.n240 VTAIL.n231 5.04292
R478 VTAIL.n186 VTAIL.n177 5.04292
R479 VTAIL.n402 VTAIL.n390 4.26717
R480 VTAIL.n24 VTAIL.n12 4.26717
R481 VTAIL.n78 VTAIL.n66 4.26717
R482 VTAIL.n132 VTAIL.n120 4.26717
R483 VTAIL.n349 VTAIL.n337 4.26717
R484 VTAIL.n295 VTAIL.n283 4.26717
R485 VTAIL.n241 VTAIL.n229 4.26717
R486 VTAIL.n187 VTAIL.n175 4.26717
R487 VTAIL.n406 VTAIL.n405 3.49141
R488 VTAIL.n430 VTAIL.n378 3.49141
R489 VTAIL.n28 VTAIL.n27 3.49141
R490 VTAIL.n52 VTAIL.n0 3.49141
R491 VTAIL.n82 VTAIL.n81 3.49141
R492 VTAIL.n106 VTAIL.n54 3.49141
R493 VTAIL.n136 VTAIL.n135 3.49141
R494 VTAIL.n160 VTAIL.n108 3.49141
R495 VTAIL.n376 VTAIL.n324 3.49141
R496 VTAIL.n353 VTAIL.n352 3.49141
R497 VTAIL.n322 VTAIL.n270 3.49141
R498 VTAIL.n299 VTAIL.n298 3.49141
R499 VTAIL.n268 VTAIL.n216 3.49141
R500 VTAIL.n245 VTAIL.n244 3.49141
R501 VTAIL.n214 VTAIL.n162 3.49141
R502 VTAIL.n191 VTAIL.n190 3.49141
R503 VTAIL.n269 VTAIL.n215 2.9574
R504 VTAIL.n377 VTAIL.n323 2.9574
R505 VTAIL.n161 VTAIL.n107 2.9574
R506 VTAIL.n396 VTAIL.n395 2.84303
R507 VTAIL.n18 VTAIL.n17 2.84303
R508 VTAIL.n72 VTAIL.n71 2.84303
R509 VTAIL.n126 VTAIL.n125 2.84303
R510 VTAIL.n343 VTAIL.n342 2.84303
R511 VTAIL.n289 VTAIL.n288 2.84303
R512 VTAIL.n235 VTAIL.n234 2.84303
R513 VTAIL.n181 VTAIL.n180 2.84303
R514 VTAIL.n409 VTAIL.n388 2.71565
R515 VTAIL.n428 VTAIL.n427 2.71565
R516 VTAIL.n31 VTAIL.n10 2.71565
R517 VTAIL.n50 VTAIL.n49 2.71565
R518 VTAIL.n85 VTAIL.n64 2.71565
R519 VTAIL.n104 VTAIL.n103 2.71565
R520 VTAIL.n139 VTAIL.n118 2.71565
R521 VTAIL.n158 VTAIL.n157 2.71565
R522 VTAIL.n374 VTAIL.n373 2.71565
R523 VTAIL.n356 VTAIL.n335 2.71565
R524 VTAIL.n320 VTAIL.n319 2.71565
R525 VTAIL.n302 VTAIL.n281 2.71565
R526 VTAIL.n266 VTAIL.n265 2.71565
R527 VTAIL.n248 VTAIL.n227 2.71565
R528 VTAIL.n212 VTAIL.n211 2.71565
R529 VTAIL.n194 VTAIL.n173 2.71565
R530 VTAIL.n410 VTAIL.n386 1.93989
R531 VTAIL.n424 VTAIL.n380 1.93989
R532 VTAIL.n32 VTAIL.n8 1.93989
R533 VTAIL.n46 VTAIL.n2 1.93989
R534 VTAIL.n86 VTAIL.n62 1.93989
R535 VTAIL.n100 VTAIL.n56 1.93989
R536 VTAIL.n140 VTAIL.n116 1.93989
R537 VTAIL.n154 VTAIL.n110 1.93989
R538 VTAIL.n370 VTAIL.n326 1.93989
R539 VTAIL.n357 VTAIL.n333 1.93989
R540 VTAIL.n316 VTAIL.n272 1.93989
R541 VTAIL.n303 VTAIL.n279 1.93989
R542 VTAIL.n262 VTAIL.n218 1.93989
R543 VTAIL.n249 VTAIL.n225 1.93989
R544 VTAIL.n208 VTAIL.n164 1.93989
R545 VTAIL.n195 VTAIL.n171 1.93989
R546 VTAIL VTAIL.n53 1.53714
R547 VTAIL VTAIL.n431 1.42076
R548 VTAIL.n415 VTAIL.n413 1.16414
R549 VTAIL.n423 VTAIL.n382 1.16414
R550 VTAIL.n37 VTAIL.n35 1.16414
R551 VTAIL.n45 VTAIL.n4 1.16414
R552 VTAIL.n91 VTAIL.n89 1.16414
R553 VTAIL.n99 VTAIL.n58 1.16414
R554 VTAIL.n145 VTAIL.n143 1.16414
R555 VTAIL.n153 VTAIL.n112 1.16414
R556 VTAIL.n369 VTAIL.n328 1.16414
R557 VTAIL.n361 VTAIL.n360 1.16414
R558 VTAIL.n315 VTAIL.n274 1.16414
R559 VTAIL.n307 VTAIL.n306 1.16414
R560 VTAIL.n261 VTAIL.n220 1.16414
R561 VTAIL.n253 VTAIL.n252 1.16414
R562 VTAIL.n207 VTAIL.n166 1.16414
R563 VTAIL.n199 VTAIL.n198 1.16414
R564 VTAIL.n323 VTAIL.n269 0.470328
R565 VTAIL.n107 VTAIL.n53 0.470328
R566 VTAIL.n414 VTAIL.n384 0.388379
R567 VTAIL.n420 VTAIL.n419 0.388379
R568 VTAIL.n36 VTAIL.n6 0.388379
R569 VTAIL.n42 VTAIL.n41 0.388379
R570 VTAIL.n90 VTAIL.n60 0.388379
R571 VTAIL.n96 VTAIL.n95 0.388379
R572 VTAIL.n144 VTAIL.n114 0.388379
R573 VTAIL.n150 VTAIL.n149 0.388379
R574 VTAIL.n366 VTAIL.n365 0.388379
R575 VTAIL.n332 VTAIL.n330 0.388379
R576 VTAIL.n312 VTAIL.n311 0.388379
R577 VTAIL.n278 VTAIL.n276 0.388379
R578 VTAIL.n258 VTAIL.n257 0.388379
R579 VTAIL.n224 VTAIL.n222 0.388379
R580 VTAIL.n204 VTAIL.n203 0.388379
R581 VTAIL.n170 VTAIL.n168 0.388379
R582 VTAIL.n396 VTAIL.n391 0.155672
R583 VTAIL.n403 VTAIL.n391 0.155672
R584 VTAIL.n404 VTAIL.n403 0.155672
R585 VTAIL.n404 VTAIL.n387 0.155672
R586 VTAIL.n411 VTAIL.n387 0.155672
R587 VTAIL.n412 VTAIL.n411 0.155672
R588 VTAIL.n412 VTAIL.n383 0.155672
R589 VTAIL.n421 VTAIL.n383 0.155672
R590 VTAIL.n422 VTAIL.n421 0.155672
R591 VTAIL.n422 VTAIL.n379 0.155672
R592 VTAIL.n429 VTAIL.n379 0.155672
R593 VTAIL.n18 VTAIL.n13 0.155672
R594 VTAIL.n25 VTAIL.n13 0.155672
R595 VTAIL.n26 VTAIL.n25 0.155672
R596 VTAIL.n26 VTAIL.n9 0.155672
R597 VTAIL.n33 VTAIL.n9 0.155672
R598 VTAIL.n34 VTAIL.n33 0.155672
R599 VTAIL.n34 VTAIL.n5 0.155672
R600 VTAIL.n43 VTAIL.n5 0.155672
R601 VTAIL.n44 VTAIL.n43 0.155672
R602 VTAIL.n44 VTAIL.n1 0.155672
R603 VTAIL.n51 VTAIL.n1 0.155672
R604 VTAIL.n72 VTAIL.n67 0.155672
R605 VTAIL.n79 VTAIL.n67 0.155672
R606 VTAIL.n80 VTAIL.n79 0.155672
R607 VTAIL.n80 VTAIL.n63 0.155672
R608 VTAIL.n87 VTAIL.n63 0.155672
R609 VTAIL.n88 VTAIL.n87 0.155672
R610 VTAIL.n88 VTAIL.n59 0.155672
R611 VTAIL.n97 VTAIL.n59 0.155672
R612 VTAIL.n98 VTAIL.n97 0.155672
R613 VTAIL.n98 VTAIL.n55 0.155672
R614 VTAIL.n105 VTAIL.n55 0.155672
R615 VTAIL.n126 VTAIL.n121 0.155672
R616 VTAIL.n133 VTAIL.n121 0.155672
R617 VTAIL.n134 VTAIL.n133 0.155672
R618 VTAIL.n134 VTAIL.n117 0.155672
R619 VTAIL.n141 VTAIL.n117 0.155672
R620 VTAIL.n142 VTAIL.n141 0.155672
R621 VTAIL.n142 VTAIL.n113 0.155672
R622 VTAIL.n151 VTAIL.n113 0.155672
R623 VTAIL.n152 VTAIL.n151 0.155672
R624 VTAIL.n152 VTAIL.n109 0.155672
R625 VTAIL.n159 VTAIL.n109 0.155672
R626 VTAIL.n375 VTAIL.n325 0.155672
R627 VTAIL.n368 VTAIL.n325 0.155672
R628 VTAIL.n368 VTAIL.n367 0.155672
R629 VTAIL.n367 VTAIL.n329 0.155672
R630 VTAIL.n359 VTAIL.n329 0.155672
R631 VTAIL.n359 VTAIL.n358 0.155672
R632 VTAIL.n358 VTAIL.n334 0.155672
R633 VTAIL.n351 VTAIL.n334 0.155672
R634 VTAIL.n351 VTAIL.n350 0.155672
R635 VTAIL.n350 VTAIL.n338 0.155672
R636 VTAIL.n343 VTAIL.n338 0.155672
R637 VTAIL.n321 VTAIL.n271 0.155672
R638 VTAIL.n314 VTAIL.n271 0.155672
R639 VTAIL.n314 VTAIL.n313 0.155672
R640 VTAIL.n313 VTAIL.n275 0.155672
R641 VTAIL.n305 VTAIL.n275 0.155672
R642 VTAIL.n305 VTAIL.n304 0.155672
R643 VTAIL.n304 VTAIL.n280 0.155672
R644 VTAIL.n297 VTAIL.n280 0.155672
R645 VTAIL.n297 VTAIL.n296 0.155672
R646 VTAIL.n296 VTAIL.n284 0.155672
R647 VTAIL.n289 VTAIL.n284 0.155672
R648 VTAIL.n267 VTAIL.n217 0.155672
R649 VTAIL.n260 VTAIL.n217 0.155672
R650 VTAIL.n260 VTAIL.n259 0.155672
R651 VTAIL.n259 VTAIL.n221 0.155672
R652 VTAIL.n251 VTAIL.n221 0.155672
R653 VTAIL.n251 VTAIL.n250 0.155672
R654 VTAIL.n250 VTAIL.n226 0.155672
R655 VTAIL.n243 VTAIL.n226 0.155672
R656 VTAIL.n243 VTAIL.n242 0.155672
R657 VTAIL.n242 VTAIL.n230 0.155672
R658 VTAIL.n235 VTAIL.n230 0.155672
R659 VTAIL.n213 VTAIL.n163 0.155672
R660 VTAIL.n206 VTAIL.n163 0.155672
R661 VTAIL.n206 VTAIL.n205 0.155672
R662 VTAIL.n205 VTAIL.n167 0.155672
R663 VTAIL.n197 VTAIL.n167 0.155672
R664 VTAIL.n197 VTAIL.n196 0.155672
R665 VTAIL.n196 VTAIL.n172 0.155672
R666 VTAIL.n189 VTAIL.n172 0.155672
R667 VTAIL.n189 VTAIL.n188 0.155672
R668 VTAIL.n188 VTAIL.n176 0.155672
R669 VTAIL.n181 VTAIL.n176 0.155672
R670 B.n568 B.n567 585
R671 B.n570 B.n118 585
R672 B.n573 B.n572 585
R673 B.n574 B.n117 585
R674 B.n576 B.n575 585
R675 B.n578 B.n116 585
R676 B.n581 B.n580 585
R677 B.n582 B.n115 585
R678 B.n584 B.n583 585
R679 B.n586 B.n114 585
R680 B.n589 B.n588 585
R681 B.n590 B.n113 585
R682 B.n592 B.n591 585
R683 B.n594 B.n112 585
R684 B.n597 B.n596 585
R685 B.n598 B.n111 585
R686 B.n600 B.n599 585
R687 B.n602 B.n110 585
R688 B.n605 B.n604 585
R689 B.n606 B.n109 585
R690 B.n608 B.n607 585
R691 B.n610 B.n108 585
R692 B.n613 B.n612 585
R693 B.n614 B.n107 585
R694 B.n616 B.n615 585
R695 B.n618 B.n106 585
R696 B.n621 B.n620 585
R697 B.n622 B.n105 585
R698 B.n624 B.n623 585
R699 B.n626 B.n104 585
R700 B.n629 B.n628 585
R701 B.n630 B.n103 585
R702 B.n632 B.n631 585
R703 B.n634 B.n102 585
R704 B.n636 B.n635 585
R705 B.n638 B.n637 585
R706 B.n641 B.n640 585
R707 B.n642 B.n97 585
R708 B.n644 B.n643 585
R709 B.n646 B.n96 585
R710 B.n649 B.n648 585
R711 B.n650 B.n95 585
R712 B.n652 B.n651 585
R713 B.n654 B.n94 585
R714 B.n657 B.n656 585
R715 B.n658 B.n91 585
R716 B.n661 B.n660 585
R717 B.n663 B.n90 585
R718 B.n666 B.n665 585
R719 B.n667 B.n89 585
R720 B.n669 B.n668 585
R721 B.n671 B.n88 585
R722 B.n674 B.n673 585
R723 B.n675 B.n87 585
R724 B.n677 B.n676 585
R725 B.n679 B.n86 585
R726 B.n682 B.n681 585
R727 B.n683 B.n85 585
R728 B.n685 B.n684 585
R729 B.n687 B.n84 585
R730 B.n690 B.n689 585
R731 B.n691 B.n83 585
R732 B.n693 B.n692 585
R733 B.n695 B.n82 585
R734 B.n698 B.n697 585
R735 B.n699 B.n81 585
R736 B.n701 B.n700 585
R737 B.n703 B.n80 585
R738 B.n706 B.n705 585
R739 B.n707 B.n79 585
R740 B.n709 B.n708 585
R741 B.n711 B.n78 585
R742 B.n714 B.n713 585
R743 B.n715 B.n77 585
R744 B.n717 B.n716 585
R745 B.n719 B.n76 585
R746 B.n722 B.n721 585
R747 B.n723 B.n75 585
R748 B.n725 B.n724 585
R749 B.n727 B.n74 585
R750 B.n730 B.n729 585
R751 B.n731 B.n73 585
R752 B.n566 B.n71 585
R753 B.n734 B.n71 585
R754 B.n565 B.n70 585
R755 B.n735 B.n70 585
R756 B.n564 B.n69 585
R757 B.n736 B.n69 585
R758 B.n563 B.n562 585
R759 B.n562 B.n65 585
R760 B.n561 B.n64 585
R761 B.n742 B.n64 585
R762 B.n560 B.n63 585
R763 B.n743 B.n63 585
R764 B.n559 B.n62 585
R765 B.n744 B.n62 585
R766 B.n558 B.n557 585
R767 B.n557 B.n58 585
R768 B.n556 B.n57 585
R769 B.n750 B.n57 585
R770 B.n555 B.n56 585
R771 B.n751 B.n56 585
R772 B.n554 B.n55 585
R773 B.n752 B.n55 585
R774 B.n553 B.n552 585
R775 B.n552 B.n51 585
R776 B.n551 B.n50 585
R777 B.n758 B.n50 585
R778 B.n550 B.n49 585
R779 B.n759 B.n49 585
R780 B.n549 B.n48 585
R781 B.n760 B.n48 585
R782 B.n548 B.n547 585
R783 B.n547 B.n44 585
R784 B.n546 B.n43 585
R785 B.n766 B.n43 585
R786 B.n545 B.n42 585
R787 B.n767 B.n42 585
R788 B.n544 B.n41 585
R789 B.n768 B.n41 585
R790 B.n543 B.n542 585
R791 B.n542 B.n37 585
R792 B.n541 B.n36 585
R793 B.n774 B.n36 585
R794 B.n540 B.n35 585
R795 B.n775 B.n35 585
R796 B.n539 B.n34 585
R797 B.n776 B.n34 585
R798 B.n538 B.n537 585
R799 B.n537 B.n30 585
R800 B.n536 B.n29 585
R801 B.n782 B.n29 585
R802 B.n535 B.n28 585
R803 B.n783 B.n28 585
R804 B.n534 B.n27 585
R805 B.n784 B.n27 585
R806 B.n533 B.n532 585
R807 B.n532 B.n23 585
R808 B.n531 B.n22 585
R809 B.n790 B.n22 585
R810 B.n530 B.n21 585
R811 B.n791 B.n21 585
R812 B.n529 B.n20 585
R813 B.n792 B.n20 585
R814 B.n528 B.n527 585
R815 B.n527 B.n19 585
R816 B.n526 B.n15 585
R817 B.n798 B.n15 585
R818 B.n525 B.n14 585
R819 B.n799 B.n14 585
R820 B.n524 B.n13 585
R821 B.n800 B.n13 585
R822 B.n523 B.n522 585
R823 B.n522 B.n12 585
R824 B.n521 B.n520 585
R825 B.n521 B.n8 585
R826 B.n519 B.n7 585
R827 B.n807 B.n7 585
R828 B.n518 B.n6 585
R829 B.n808 B.n6 585
R830 B.n517 B.n5 585
R831 B.n809 B.n5 585
R832 B.n516 B.n515 585
R833 B.n515 B.n4 585
R834 B.n514 B.n119 585
R835 B.n514 B.n513 585
R836 B.n504 B.n120 585
R837 B.n121 B.n120 585
R838 B.n506 B.n505 585
R839 B.n507 B.n506 585
R840 B.n503 B.n126 585
R841 B.n126 B.n125 585
R842 B.n502 B.n501 585
R843 B.n501 B.n500 585
R844 B.n128 B.n127 585
R845 B.n493 B.n128 585
R846 B.n492 B.n491 585
R847 B.n494 B.n492 585
R848 B.n490 B.n133 585
R849 B.n133 B.n132 585
R850 B.n489 B.n488 585
R851 B.n488 B.n487 585
R852 B.n135 B.n134 585
R853 B.n136 B.n135 585
R854 B.n480 B.n479 585
R855 B.n481 B.n480 585
R856 B.n478 B.n141 585
R857 B.n141 B.n140 585
R858 B.n477 B.n476 585
R859 B.n476 B.n475 585
R860 B.n143 B.n142 585
R861 B.n144 B.n143 585
R862 B.n468 B.n467 585
R863 B.n469 B.n468 585
R864 B.n466 B.n148 585
R865 B.n152 B.n148 585
R866 B.n465 B.n464 585
R867 B.n464 B.n463 585
R868 B.n150 B.n149 585
R869 B.n151 B.n150 585
R870 B.n456 B.n455 585
R871 B.n457 B.n456 585
R872 B.n454 B.n157 585
R873 B.n157 B.n156 585
R874 B.n453 B.n452 585
R875 B.n452 B.n451 585
R876 B.n159 B.n158 585
R877 B.n160 B.n159 585
R878 B.n444 B.n443 585
R879 B.n445 B.n444 585
R880 B.n442 B.n165 585
R881 B.n165 B.n164 585
R882 B.n441 B.n440 585
R883 B.n440 B.n439 585
R884 B.n167 B.n166 585
R885 B.n168 B.n167 585
R886 B.n432 B.n431 585
R887 B.n433 B.n432 585
R888 B.n430 B.n173 585
R889 B.n173 B.n172 585
R890 B.n429 B.n428 585
R891 B.n428 B.n427 585
R892 B.n175 B.n174 585
R893 B.n176 B.n175 585
R894 B.n420 B.n419 585
R895 B.n421 B.n420 585
R896 B.n418 B.n181 585
R897 B.n181 B.n180 585
R898 B.n417 B.n416 585
R899 B.n416 B.n415 585
R900 B.n183 B.n182 585
R901 B.n184 B.n183 585
R902 B.n408 B.n407 585
R903 B.n409 B.n408 585
R904 B.n406 B.n189 585
R905 B.n189 B.n188 585
R906 B.n405 B.n404 585
R907 B.n404 B.n403 585
R908 B.n400 B.n193 585
R909 B.n399 B.n398 585
R910 B.n396 B.n194 585
R911 B.n396 B.n192 585
R912 B.n395 B.n394 585
R913 B.n393 B.n392 585
R914 B.n391 B.n196 585
R915 B.n389 B.n388 585
R916 B.n387 B.n197 585
R917 B.n386 B.n385 585
R918 B.n383 B.n198 585
R919 B.n381 B.n380 585
R920 B.n379 B.n199 585
R921 B.n378 B.n377 585
R922 B.n375 B.n200 585
R923 B.n373 B.n372 585
R924 B.n371 B.n201 585
R925 B.n370 B.n369 585
R926 B.n367 B.n202 585
R927 B.n365 B.n364 585
R928 B.n363 B.n203 585
R929 B.n362 B.n361 585
R930 B.n359 B.n204 585
R931 B.n357 B.n356 585
R932 B.n355 B.n205 585
R933 B.n354 B.n353 585
R934 B.n351 B.n206 585
R935 B.n349 B.n348 585
R936 B.n347 B.n207 585
R937 B.n346 B.n345 585
R938 B.n343 B.n208 585
R939 B.n341 B.n340 585
R940 B.n339 B.n209 585
R941 B.n338 B.n337 585
R942 B.n335 B.n210 585
R943 B.n333 B.n332 585
R944 B.n331 B.n211 585
R945 B.n329 B.n328 585
R946 B.n326 B.n214 585
R947 B.n324 B.n323 585
R948 B.n322 B.n215 585
R949 B.n321 B.n320 585
R950 B.n318 B.n216 585
R951 B.n316 B.n315 585
R952 B.n314 B.n217 585
R953 B.n313 B.n312 585
R954 B.n310 B.n218 585
R955 B.n308 B.n307 585
R956 B.n306 B.n219 585
R957 B.n305 B.n304 585
R958 B.n302 B.n223 585
R959 B.n300 B.n299 585
R960 B.n298 B.n224 585
R961 B.n297 B.n296 585
R962 B.n294 B.n225 585
R963 B.n292 B.n291 585
R964 B.n290 B.n226 585
R965 B.n289 B.n288 585
R966 B.n286 B.n227 585
R967 B.n284 B.n283 585
R968 B.n282 B.n228 585
R969 B.n281 B.n280 585
R970 B.n278 B.n229 585
R971 B.n276 B.n275 585
R972 B.n274 B.n230 585
R973 B.n273 B.n272 585
R974 B.n270 B.n231 585
R975 B.n268 B.n267 585
R976 B.n266 B.n232 585
R977 B.n265 B.n264 585
R978 B.n262 B.n233 585
R979 B.n260 B.n259 585
R980 B.n258 B.n234 585
R981 B.n257 B.n256 585
R982 B.n254 B.n235 585
R983 B.n252 B.n251 585
R984 B.n250 B.n236 585
R985 B.n249 B.n248 585
R986 B.n246 B.n237 585
R987 B.n244 B.n243 585
R988 B.n242 B.n238 585
R989 B.n241 B.n240 585
R990 B.n191 B.n190 585
R991 B.n192 B.n191 585
R992 B.n402 B.n401 585
R993 B.n403 B.n402 585
R994 B.n187 B.n186 585
R995 B.n188 B.n187 585
R996 B.n411 B.n410 585
R997 B.n410 B.n409 585
R998 B.n412 B.n185 585
R999 B.n185 B.n184 585
R1000 B.n414 B.n413 585
R1001 B.n415 B.n414 585
R1002 B.n179 B.n178 585
R1003 B.n180 B.n179 585
R1004 B.n423 B.n422 585
R1005 B.n422 B.n421 585
R1006 B.n424 B.n177 585
R1007 B.n177 B.n176 585
R1008 B.n426 B.n425 585
R1009 B.n427 B.n426 585
R1010 B.n171 B.n170 585
R1011 B.n172 B.n171 585
R1012 B.n435 B.n434 585
R1013 B.n434 B.n433 585
R1014 B.n436 B.n169 585
R1015 B.n169 B.n168 585
R1016 B.n438 B.n437 585
R1017 B.n439 B.n438 585
R1018 B.n163 B.n162 585
R1019 B.n164 B.n163 585
R1020 B.n447 B.n446 585
R1021 B.n446 B.n445 585
R1022 B.n448 B.n161 585
R1023 B.n161 B.n160 585
R1024 B.n450 B.n449 585
R1025 B.n451 B.n450 585
R1026 B.n155 B.n154 585
R1027 B.n156 B.n155 585
R1028 B.n459 B.n458 585
R1029 B.n458 B.n457 585
R1030 B.n460 B.n153 585
R1031 B.n153 B.n151 585
R1032 B.n462 B.n461 585
R1033 B.n463 B.n462 585
R1034 B.n147 B.n146 585
R1035 B.n152 B.n147 585
R1036 B.n471 B.n470 585
R1037 B.n470 B.n469 585
R1038 B.n472 B.n145 585
R1039 B.n145 B.n144 585
R1040 B.n474 B.n473 585
R1041 B.n475 B.n474 585
R1042 B.n139 B.n138 585
R1043 B.n140 B.n139 585
R1044 B.n483 B.n482 585
R1045 B.n482 B.n481 585
R1046 B.n484 B.n137 585
R1047 B.n137 B.n136 585
R1048 B.n486 B.n485 585
R1049 B.n487 B.n486 585
R1050 B.n131 B.n130 585
R1051 B.n132 B.n131 585
R1052 B.n496 B.n495 585
R1053 B.n495 B.n494 585
R1054 B.n497 B.n129 585
R1055 B.n493 B.n129 585
R1056 B.n499 B.n498 585
R1057 B.n500 B.n499 585
R1058 B.n124 B.n123 585
R1059 B.n125 B.n124 585
R1060 B.n509 B.n508 585
R1061 B.n508 B.n507 585
R1062 B.n510 B.n122 585
R1063 B.n122 B.n121 585
R1064 B.n512 B.n511 585
R1065 B.n513 B.n512 585
R1066 B.n3 B.n0 585
R1067 B.n4 B.n3 585
R1068 B.n806 B.n1 585
R1069 B.n807 B.n806 585
R1070 B.n805 B.n804 585
R1071 B.n805 B.n8 585
R1072 B.n803 B.n9 585
R1073 B.n12 B.n9 585
R1074 B.n802 B.n801 585
R1075 B.n801 B.n800 585
R1076 B.n11 B.n10 585
R1077 B.n799 B.n11 585
R1078 B.n797 B.n796 585
R1079 B.n798 B.n797 585
R1080 B.n795 B.n16 585
R1081 B.n19 B.n16 585
R1082 B.n794 B.n793 585
R1083 B.n793 B.n792 585
R1084 B.n18 B.n17 585
R1085 B.n791 B.n18 585
R1086 B.n789 B.n788 585
R1087 B.n790 B.n789 585
R1088 B.n787 B.n24 585
R1089 B.n24 B.n23 585
R1090 B.n786 B.n785 585
R1091 B.n785 B.n784 585
R1092 B.n26 B.n25 585
R1093 B.n783 B.n26 585
R1094 B.n781 B.n780 585
R1095 B.n782 B.n781 585
R1096 B.n779 B.n31 585
R1097 B.n31 B.n30 585
R1098 B.n778 B.n777 585
R1099 B.n777 B.n776 585
R1100 B.n33 B.n32 585
R1101 B.n775 B.n33 585
R1102 B.n773 B.n772 585
R1103 B.n774 B.n773 585
R1104 B.n771 B.n38 585
R1105 B.n38 B.n37 585
R1106 B.n770 B.n769 585
R1107 B.n769 B.n768 585
R1108 B.n40 B.n39 585
R1109 B.n767 B.n40 585
R1110 B.n765 B.n764 585
R1111 B.n766 B.n765 585
R1112 B.n763 B.n45 585
R1113 B.n45 B.n44 585
R1114 B.n762 B.n761 585
R1115 B.n761 B.n760 585
R1116 B.n47 B.n46 585
R1117 B.n759 B.n47 585
R1118 B.n757 B.n756 585
R1119 B.n758 B.n757 585
R1120 B.n755 B.n52 585
R1121 B.n52 B.n51 585
R1122 B.n754 B.n753 585
R1123 B.n753 B.n752 585
R1124 B.n54 B.n53 585
R1125 B.n751 B.n54 585
R1126 B.n749 B.n748 585
R1127 B.n750 B.n749 585
R1128 B.n747 B.n59 585
R1129 B.n59 B.n58 585
R1130 B.n746 B.n745 585
R1131 B.n745 B.n744 585
R1132 B.n61 B.n60 585
R1133 B.n743 B.n61 585
R1134 B.n741 B.n740 585
R1135 B.n742 B.n741 585
R1136 B.n739 B.n66 585
R1137 B.n66 B.n65 585
R1138 B.n738 B.n737 585
R1139 B.n737 B.n736 585
R1140 B.n68 B.n67 585
R1141 B.n735 B.n68 585
R1142 B.n733 B.n732 585
R1143 B.n734 B.n733 585
R1144 B.n810 B.n809 585
R1145 B.n808 B.n2 585
R1146 B.n733 B.n73 487.695
R1147 B.n568 B.n71 487.695
R1148 B.n404 B.n191 487.695
R1149 B.n402 B.n193 487.695
R1150 B.n98 B.t13 317.659
R1151 B.n220 B.t7 317.659
R1152 B.n92 B.t10 317.659
R1153 B.n212 B.t17 317.659
R1154 B.n92 B.t8 287.836
R1155 B.n98 B.t12 287.836
R1156 B.n220 B.t4 287.836
R1157 B.n212 B.t15 287.836
R1158 B.n569 B.n72 256.663
R1159 B.n571 B.n72 256.663
R1160 B.n577 B.n72 256.663
R1161 B.n579 B.n72 256.663
R1162 B.n585 B.n72 256.663
R1163 B.n587 B.n72 256.663
R1164 B.n593 B.n72 256.663
R1165 B.n595 B.n72 256.663
R1166 B.n601 B.n72 256.663
R1167 B.n603 B.n72 256.663
R1168 B.n609 B.n72 256.663
R1169 B.n611 B.n72 256.663
R1170 B.n617 B.n72 256.663
R1171 B.n619 B.n72 256.663
R1172 B.n625 B.n72 256.663
R1173 B.n627 B.n72 256.663
R1174 B.n633 B.n72 256.663
R1175 B.n101 B.n72 256.663
R1176 B.n639 B.n72 256.663
R1177 B.n645 B.n72 256.663
R1178 B.n647 B.n72 256.663
R1179 B.n653 B.n72 256.663
R1180 B.n655 B.n72 256.663
R1181 B.n662 B.n72 256.663
R1182 B.n664 B.n72 256.663
R1183 B.n670 B.n72 256.663
R1184 B.n672 B.n72 256.663
R1185 B.n678 B.n72 256.663
R1186 B.n680 B.n72 256.663
R1187 B.n686 B.n72 256.663
R1188 B.n688 B.n72 256.663
R1189 B.n694 B.n72 256.663
R1190 B.n696 B.n72 256.663
R1191 B.n702 B.n72 256.663
R1192 B.n704 B.n72 256.663
R1193 B.n710 B.n72 256.663
R1194 B.n712 B.n72 256.663
R1195 B.n718 B.n72 256.663
R1196 B.n720 B.n72 256.663
R1197 B.n726 B.n72 256.663
R1198 B.n728 B.n72 256.663
R1199 B.n397 B.n192 256.663
R1200 B.n195 B.n192 256.663
R1201 B.n390 B.n192 256.663
R1202 B.n384 B.n192 256.663
R1203 B.n382 B.n192 256.663
R1204 B.n376 B.n192 256.663
R1205 B.n374 B.n192 256.663
R1206 B.n368 B.n192 256.663
R1207 B.n366 B.n192 256.663
R1208 B.n360 B.n192 256.663
R1209 B.n358 B.n192 256.663
R1210 B.n352 B.n192 256.663
R1211 B.n350 B.n192 256.663
R1212 B.n344 B.n192 256.663
R1213 B.n342 B.n192 256.663
R1214 B.n336 B.n192 256.663
R1215 B.n334 B.n192 256.663
R1216 B.n327 B.n192 256.663
R1217 B.n325 B.n192 256.663
R1218 B.n319 B.n192 256.663
R1219 B.n317 B.n192 256.663
R1220 B.n311 B.n192 256.663
R1221 B.n309 B.n192 256.663
R1222 B.n303 B.n192 256.663
R1223 B.n301 B.n192 256.663
R1224 B.n295 B.n192 256.663
R1225 B.n293 B.n192 256.663
R1226 B.n287 B.n192 256.663
R1227 B.n285 B.n192 256.663
R1228 B.n279 B.n192 256.663
R1229 B.n277 B.n192 256.663
R1230 B.n271 B.n192 256.663
R1231 B.n269 B.n192 256.663
R1232 B.n263 B.n192 256.663
R1233 B.n261 B.n192 256.663
R1234 B.n255 B.n192 256.663
R1235 B.n253 B.n192 256.663
R1236 B.n247 B.n192 256.663
R1237 B.n245 B.n192 256.663
R1238 B.n239 B.n192 256.663
R1239 B.n812 B.n811 256.663
R1240 B.n99 B.t14 251.138
R1241 B.n221 B.t6 251.138
R1242 B.n93 B.t11 251.138
R1243 B.n213 B.t16 251.138
R1244 B.n729 B.n727 163.367
R1245 B.n725 B.n75 163.367
R1246 B.n721 B.n719 163.367
R1247 B.n717 B.n77 163.367
R1248 B.n713 B.n711 163.367
R1249 B.n709 B.n79 163.367
R1250 B.n705 B.n703 163.367
R1251 B.n701 B.n81 163.367
R1252 B.n697 B.n695 163.367
R1253 B.n693 B.n83 163.367
R1254 B.n689 B.n687 163.367
R1255 B.n685 B.n85 163.367
R1256 B.n681 B.n679 163.367
R1257 B.n677 B.n87 163.367
R1258 B.n673 B.n671 163.367
R1259 B.n669 B.n89 163.367
R1260 B.n665 B.n663 163.367
R1261 B.n661 B.n91 163.367
R1262 B.n656 B.n654 163.367
R1263 B.n652 B.n95 163.367
R1264 B.n648 B.n646 163.367
R1265 B.n644 B.n97 163.367
R1266 B.n640 B.n638 163.367
R1267 B.n635 B.n634 163.367
R1268 B.n632 B.n103 163.367
R1269 B.n628 B.n626 163.367
R1270 B.n624 B.n105 163.367
R1271 B.n620 B.n618 163.367
R1272 B.n616 B.n107 163.367
R1273 B.n612 B.n610 163.367
R1274 B.n608 B.n109 163.367
R1275 B.n604 B.n602 163.367
R1276 B.n600 B.n111 163.367
R1277 B.n596 B.n594 163.367
R1278 B.n592 B.n113 163.367
R1279 B.n588 B.n586 163.367
R1280 B.n584 B.n115 163.367
R1281 B.n580 B.n578 163.367
R1282 B.n576 B.n117 163.367
R1283 B.n572 B.n570 163.367
R1284 B.n404 B.n189 163.367
R1285 B.n408 B.n189 163.367
R1286 B.n408 B.n183 163.367
R1287 B.n416 B.n183 163.367
R1288 B.n416 B.n181 163.367
R1289 B.n420 B.n181 163.367
R1290 B.n420 B.n175 163.367
R1291 B.n428 B.n175 163.367
R1292 B.n428 B.n173 163.367
R1293 B.n432 B.n173 163.367
R1294 B.n432 B.n167 163.367
R1295 B.n440 B.n167 163.367
R1296 B.n440 B.n165 163.367
R1297 B.n444 B.n165 163.367
R1298 B.n444 B.n159 163.367
R1299 B.n452 B.n159 163.367
R1300 B.n452 B.n157 163.367
R1301 B.n456 B.n157 163.367
R1302 B.n456 B.n150 163.367
R1303 B.n464 B.n150 163.367
R1304 B.n464 B.n148 163.367
R1305 B.n468 B.n148 163.367
R1306 B.n468 B.n143 163.367
R1307 B.n476 B.n143 163.367
R1308 B.n476 B.n141 163.367
R1309 B.n480 B.n141 163.367
R1310 B.n480 B.n135 163.367
R1311 B.n488 B.n135 163.367
R1312 B.n488 B.n133 163.367
R1313 B.n492 B.n133 163.367
R1314 B.n492 B.n128 163.367
R1315 B.n501 B.n128 163.367
R1316 B.n501 B.n126 163.367
R1317 B.n506 B.n126 163.367
R1318 B.n506 B.n120 163.367
R1319 B.n514 B.n120 163.367
R1320 B.n515 B.n514 163.367
R1321 B.n515 B.n5 163.367
R1322 B.n6 B.n5 163.367
R1323 B.n7 B.n6 163.367
R1324 B.n521 B.n7 163.367
R1325 B.n522 B.n521 163.367
R1326 B.n522 B.n13 163.367
R1327 B.n14 B.n13 163.367
R1328 B.n15 B.n14 163.367
R1329 B.n527 B.n15 163.367
R1330 B.n527 B.n20 163.367
R1331 B.n21 B.n20 163.367
R1332 B.n22 B.n21 163.367
R1333 B.n532 B.n22 163.367
R1334 B.n532 B.n27 163.367
R1335 B.n28 B.n27 163.367
R1336 B.n29 B.n28 163.367
R1337 B.n537 B.n29 163.367
R1338 B.n537 B.n34 163.367
R1339 B.n35 B.n34 163.367
R1340 B.n36 B.n35 163.367
R1341 B.n542 B.n36 163.367
R1342 B.n542 B.n41 163.367
R1343 B.n42 B.n41 163.367
R1344 B.n43 B.n42 163.367
R1345 B.n547 B.n43 163.367
R1346 B.n547 B.n48 163.367
R1347 B.n49 B.n48 163.367
R1348 B.n50 B.n49 163.367
R1349 B.n552 B.n50 163.367
R1350 B.n552 B.n55 163.367
R1351 B.n56 B.n55 163.367
R1352 B.n57 B.n56 163.367
R1353 B.n557 B.n57 163.367
R1354 B.n557 B.n62 163.367
R1355 B.n63 B.n62 163.367
R1356 B.n64 B.n63 163.367
R1357 B.n562 B.n64 163.367
R1358 B.n562 B.n69 163.367
R1359 B.n70 B.n69 163.367
R1360 B.n71 B.n70 163.367
R1361 B.n398 B.n396 163.367
R1362 B.n396 B.n395 163.367
R1363 B.n392 B.n391 163.367
R1364 B.n389 B.n197 163.367
R1365 B.n385 B.n383 163.367
R1366 B.n381 B.n199 163.367
R1367 B.n377 B.n375 163.367
R1368 B.n373 B.n201 163.367
R1369 B.n369 B.n367 163.367
R1370 B.n365 B.n203 163.367
R1371 B.n361 B.n359 163.367
R1372 B.n357 B.n205 163.367
R1373 B.n353 B.n351 163.367
R1374 B.n349 B.n207 163.367
R1375 B.n345 B.n343 163.367
R1376 B.n341 B.n209 163.367
R1377 B.n337 B.n335 163.367
R1378 B.n333 B.n211 163.367
R1379 B.n328 B.n326 163.367
R1380 B.n324 B.n215 163.367
R1381 B.n320 B.n318 163.367
R1382 B.n316 B.n217 163.367
R1383 B.n312 B.n310 163.367
R1384 B.n308 B.n219 163.367
R1385 B.n304 B.n302 163.367
R1386 B.n300 B.n224 163.367
R1387 B.n296 B.n294 163.367
R1388 B.n292 B.n226 163.367
R1389 B.n288 B.n286 163.367
R1390 B.n284 B.n228 163.367
R1391 B.n280 B.n278 163.367
R1392 B.n276 B.n230 163.367
R1393 B.n272 B.n270 163.367
R1394 B.n268 B.n232 163.367
R1395 B.n264 B.n262 163.367
R1396 B.n260 B.n234 163.367
R1397 B.n256 B.n254 163.367
R1398 B.n252 B.n236 163.367
R1399 B.n248 B.n246 163.367
R1400 B.n244 B.n238 163.367
R1401 B.n240 B.n191 163.367
R1402 B.n402 B.n187 163.367
R1403 B.n410 B.n187 163.367
R1404 B.n410 B.n185 163.367
R1405 B.n414 B.n185 163.367
R1406 B.n414 B.n179 163.367
R1407 B.n422 B.n179 163.367
R1408 B.n422 B.n177 163.367
R1409 B.n426 B.n177 163.367
R1410 B.n426 B.n171 163.367
R1411 B.n434 B.n171 163.367
R1412 B.n434 B.n169 163.367
R1413 B.n438 B.n169 163.367
R1414 B.n438 B.n163 163.367
R1415 B.n446 B.n163 163.367
R1416 B.n446 B.n161 163.367
R1417 B.n450 B.n161 163.367
R1418 B.n450 B.n155 163.367
R1419 B.n458 B.n155 163.367
R1420 B.n458 B.n153 163.367
R1421 B.n462 B.n153 163.367
R1422 B.n462 B.n147 163.367
R1423 B.n470 B.n147 163.367
R1424 B.n470 B.n145 163.367
R1425 B.n474 B.n145 163.367
R1426 B.n474 B.n139 163.367
R1427 B.n482 B.n139 163.367
R1428 B.n482 B.n137 163.367
R1429 B.n486 B.n137 163.367
R1430 B.n486 B.n131 163.367
R1431 B.n495 B.n131 163.367
R1432 B.n495 B.n129 163.367
R1433 B.n499 B.n129 163.367
R1434 B.n499 B.n124 163.367
R1435 B.n508 B.n124 163.367
R1436 B.n508 B.n122 163.367
R1437 B.n512 B.n122 163.367
R1438 B.n512 B.n3 163.367
R1439 B.n810 B.n3 163.367
R1440 B.n806 B.n2 163.367
R1441 B.n806 B.n805 163.367
R1442 B.n805 B.n9 163.367
R1443 B.n801 B.n9 163.367
R1444 B.n801 B.n11 163.367
R1445 B.n797 B.n11 163.367
R1446 B.n797 B.n16 163.367
R1447 B.n793 B.n16 163.367
R1448 B.n793 B.n18 163.367
R1449 B.n789 B.n18 163.367
R1450 B.n789 B.n24 163.367
R1451 B.n785 B.n24 163.367
R1452 B.n785 B.n26 163.367
R1453 B.n781 B.n26 163.367
R1454 B.n781 B.n31 163.367
R1455 B.n777 B.n31 163.367
R1456 B.n777 B.n33 163.367
R1457 B.n773 B.n33 163.367
R1458 B.n773 B.n38 163.367
R1459 B.n769 B.n38 163.367
R1460 B.n769 B.n40 163.367
R1461 B.n765 B.n40 163.367
R1462 B.n765 B.n45 163.367
R1463 B.n761 B.n45 163.367
R1464 B.n761 B.n47 163.367
R1465 B.n757 B.n47 163.367
R1466 B.n757 B.n52 163.367
R1467 B.n753 B.n52 163.367
R1468 B.n753 B.n54 163.367
R1469 B.n749 B.n54 163.367
R1470 B.n749 B.n59 163.367
R1471 B.n745 B.n59 163.367
R1472 B.n745 B.n61 163.367
R1473 B.n741 B.n61 163.367
R1474 B.n741 B.n66 163.367
R1475 B.n737 B.n66 163.367
R1476 B.n737 B.n68 163.367
R1477 B.n733 B.n68 163.367
R1478 B.n403 B.n192 81.851
R1479 B.n734 B.n72 81.851
R1480 B.n728 B.n73 71.676
R1481 B.n727 B.n726 71.676
R1482 B.n720 B.n75 71.676
R1483 B.n719 B.n718 71.676
R1484 B.n712 B.n77 71.676
R1485 B.n711 B.n710 71.676
R1486 B.n704 B.n79 71.676
R1487 B.n703 B.n702 71.676
R1488 B.n696 B.n81 71.676
R1489 B.n695 B.n694 71.676
R1490 B.n688 B.n83 71.676
R1491 B.n687 B.n686 71.676
R1492 B.n680 B.n85 71.676
R1493 B.n679 B.n678 71.676
R1494 B.n672 B.n87 71.676
R1495 B.n671 B.n670 71.676
R1496 B.n664 B.n89 71.676
R1497 B.n663 B.n662 71.676
R1498 B.n655 B.n91 71.676
R1499 B.n654 B.n653 71.676
R1500 B.n647 B.n95 71.676
R1501 B.n646 B.n645 71.676
R1502 B.n639 B.n97 71.676
R1503 B.n638 B.n101 71.676
R1504 B.n634 B.n633 71.676
R1505 B.n627 B.n103 71.676
R1506 B.n626 B.n625 71.676
R1507 B.n619 B.n105 71.676
R1508 B.n618 B.n617 71.676
R1509 B.n611 B.n107 71.676
R1510 B.n610 B.n609 71.676
R1511 B.n603 B.n109 71.676
R1512 B.n602 B.n601 71.676
R1513 B.n595 B.n111 71.676
R1514 B.n594 B.n593 71.676
R1515 B.n587 B.n113 71.676
R1516 B.n586 B.n585 71.676
R1517 B.n579 B.n115 71.676
R1518 B.n578 B.n577 71.676
R1519 B.n571 B.n117 71.676
R1520 B.n570 B.n569 71.676
R1521 B.n569 B.n568 71.676
R1522 B.n572 B.n571 71.676
R1523 B.n577 B.n576 71.676
R1524 B.n580 B.n579 71.676
R1525 B.n585 B.n584 71.676
R1526 B.n588 B.n587 71.676
R1527 B.n593 B.n592 71.676
R1528 B.n596 B.n595 71.676
R1529 B.n601 B.n600 71.676
R1530 B.n604 B.n603 71.676
R1531 B.n609 B.n608 71.676
R1532 B.n612 B.n611 71.676
R1533 B.n617 B.n616 71.676
R1534 B.n620 B.n619 71.676
R1535 B.n625 B.n624 71.676
R1536 B.n628 B.n627 71.676
R1537 B.n633 B.n632 71.676
R1538 B.n635 B.n101 71.676
R1539 B.n640 B.n639 71.676
R1540 B.n645 B.n644 71.676
R1541 B.n648 B.n647 71.676
R1542 B.n653 B.n652 71.676
R1543 B.n656 B.n655 71.676
R1544 B.n662 B.n661 71.676
R1545 B.n665 B.n664 71.676
R1546 B.n670 B.n669 71.676
R1547 B.n673 B.n672 71.676
R1548 B.n678 B.n677 71.676
R1549 B.n681 B.n680 71.676
R1550 B.n686 B.n685 71.676
R1551 B.n689 B.n688 71.676
R1552 B.n694 B.n693 71.676
R1553 B.n697 B.n696 71.676
R1554 B.n702 B.n701 71.676
R1555 B.n705 B.n704 71.676
R1556 B.n710 B.n709 71.676
R1557 B.n713 B.n712 71.676
R1558 B.n718 B.n717 71.676
R1559 B.n721 B.n720 71.676
R1560 B.n726 B.n725 71.676
R1561 B.n729 B.n728 71.676
R1562 B.n397 B.n193 71.676
R1563 B.n395 B.n195 71.676
R1564 B.n391 B.n390 71.676
R1565 B.n384 B.n197 71.676
R1566 B.n383 B.n382 71.676
R1567 B.n376 B.n199 71.676
R1568 B.n375 B.n374 71.676
R1569 B.n368 B.n201 71.676
R1570 B.n367 B.n366 71.676
R1571 B.n360 B.n203 71.676
R1572 B.n359 B.n358 71.676
R1573 B.n352 B.n205 71.676
R1574 B.n351 B.n350 71.676
R1575 B.n344 B.n207 71.676
R1576 B.n343 B.n342 71.676
R1577 B.n336 B.n209 71.676
R1578 B.n335 B.n334 71.676
R1579 B.n327 B.n211 71.676
R1580 B.n326 B.n325 71.676
R1581 B.n319 B.n215 71.676
R1582 B.n318 B.n317 71.676
R1583 B.n311 B.n217 71.676
R1584 B.n310 B.n309 71.676
R1585 B.n303 B.n219 71.676
R1586 B.n302 B.n301 71.676
R1587 B.n295 B.n224 71.676
R1588 B.n294 B.n293 71.676
R1589 B.n287 B.n226 71.676
R1590 B.n286 B.n285 71.676
R1591 B.n279 B.n228 71.676
R1592 B.n278 B.n277 71.676
R1593 B.n271 B.n230 71.676
R1594 B.n270 B.n269 71.676
R1595 B.n263 B.n232 71.676
R1596 B.n262 B.n261 71.676
R1597 B.n255 B.n234 71.676
R1598 B.n254 B.n253 71.676
R1599 B.n247 B.n236 71.676
R1600 B.n246 B.n245 71.676
R1601 B.n239 B.n238 71.676
R1602 B.n398 B.n397 71.676
R1603 B.n392 B.n195 71.676
R1604 B.n390 B.n389 71.676
R1605 B.n385 B.n384 71.676
R1606 B.n382 B.n381 71.676
R1607 B.n377 B.n376 71.676
R1608 B.n374 B.n373 71.676
R1609 B.n369 B.n368 71.676
R1610 B.n366 B.n365 71.676
R1611 B.n361 B.n360 71.676
R1612 B.n358 B.n357 71.676
R1613 B.n353 B.n352 71.676
R1614 B.n350 B.n349 71.676
R1615 B.n345 B.n344 71.676
R1616 B.n342 B.n341 71.676
R1617 B.n337 B.n336 71.676
R1618 B.n334 B.n333 71.676
R1619 B.n328 B.n327 71.676
R1620 B.n325 B.n324 71.676
R1621 B.n320 B.n319 71.676
R1622 B.n317 B.n316 71.676
R1623 B.n312 B.n311 71.676
R1624 B.n309 B.n308 71.676
R1625 B.n304 B.n303 71.676
R1626 B.n301 B.n300 71.676
R1627 B.n296 B.n295 71.676
R1628 B.n293 B.n292 71.676
R1629 B.n288 B.n287 71.676
R1630 B.n285 B.n284 71.676
R1631 B.n280 B.n279 71.676
R1632 B.n277 B.n276 71.676
R1633 B.n272 B.n271 71.676
R1634 B.n269 B.n268 71.676
R1635 B.n264 B.n263 71.676
R1636 B.n261 B.n260 71.676
R1637 B.n256 B.n255 71.676
R1638 B.n253 B.n252 71.676
R1639 B.n248 B.n247 71.676
R1640 B.n245 B.n244 71.676
R1641 B.n240 B.n239 71.676
R1642 B.n811 B.n810 71.676
R1643 B.n811 B.n2 71.676
R1644 B.n93 B.n92 66.5217
R1645 B.n99 B.n98 66.5217
R1646 B.n221 B.n220 66.5217
R1647 B.n213 B.n212 66.5217
R1648 B.n659 B.n93 59.5399
R1649 B.n100 B.n99 59.5399
R1650 B.n222 B.n221 59.5399
R1651 B.n330 B.n213 59.5399
R1652 B.n403 B.n188 48.3991
R1653 B.n409 B.n188 48.3991
R1654 B.n409 B.n184 48.3991
R1655 B.n415 B.n184 48.3991
R1656 B.n415 B.n180 48.3991
R1657 B.n421 B.n180 48.3991
R1658 B.n421 B.n176 48.3991
R1659 B.n427 B.n176 48.3991
R1660 B.n433 B.n172 48.3991
R1661 B.n433 B.n168 48.3991
R1662 B.n439 B.n168 48.3991
R1663 B.n439 B.n164 48.3991
R1664 B.n445 B.n164 48.3991
R1665 B.n445 B.n160 48.3991
R1666 B.n451 B.n160 48.3991
R1667 B.n451 B.n156 48.3991
R1668 B.n457 B.n156 48.3991
R1669 B.n457 B.n151 48.3991
R1670 B.n463 B.n151 48.3991
R1671 B.n463 B.n152 48.3991
R1672 B.n469 B.n144 48.3991
R1673 B.n475 B.n144 48.3991
R1674 B.n475 B.n140 48.3991
R1675 B.n481 B.n140 48.3991
R1676 B.n481 B.n136 48.3991
R1677 B.n487 B.n136 48.3991
R1678 B.n487 B.n132 48.3991
R1679 B.n494 B.n132 48.3991
R1680 B.n494 B.n493 48.3991
R1681 B.n500 B.n125 48.3991
R1682 B.n507 B.n125 48.3991
R1683 B.n507 B.n121 48.3991
R1684 B.n513 B.n121 48.3991
R1685 B.n513 B.n4 48.3991
R1686 B.n809 B.n4 48.3991
R1687 B.n809 B.n808 48.3991
R1688 B.n808 B.n807 48.3991
R1689 B.n807 B.n8 48.3991
R1690 B.n12 B.n8 48.3991
R1691 B.n800 B.n12 48.3991
R1692 B.n800 B.n799 48.3991
R1693 B.n799 B.n798 48.3991
R1694 B.n792 B.n19 48.3991
R1695 B.n792 B.n791 48.3991
R1696 B.n791 B.n790 48.3991
R1697 B.n790 B.n23 48.3991
R1698 B.n784 B.n23 48.3991
R1699 B.n784 B.n783 48.3991
R1700 B.n783 B.n782 48.3991
R1701 B.n782 B.n30 48.3991
R1702 B.n776 B.n30 48.3991
R1703 B.n775 B.n774 48.3991
R1704 B.n774 B.n37 48.3991
R1705 B.n768 B.n37 48.3991
R1706 B.n768 B.n767 48.3991
R1707 B.n767 B.n766 48.3991
R1708 B.n766 B.n44 48.3991
R1709 B.n760 B.n44 48.3991
R1710 B.n760 B.n759 48.3991
R1711 B.n759 B.n758 48.3991
R1712 B.n758 B.n51 48.3991
R1713 B.n752 B.n51 48.3991
R1714 B.n752 B.n751 48.3991
R1715 B.n750 B.n58 48.3991
R1716 B.n744 B.n58 48.3991
R1717 B.n744 B.n743 48.3991
R1718 B.n743 B.n742 48.3991
R1719 B.n742 B.n65 48.3991
R1720 B.n736 B.n65 48.3991
R1721 B.n736 B.n735 48.3991
R1722 B.n735 B.n734 48.3991
R1723 B.n493 B.t2 41.2816
R1724 B.n19 B.t3 41.2816
R1725 B.n152 B.t1 37.0112
R1726 B.t0 B.n775 37.0112
R1727 B.n401 B.n400 31.6883
R1728 B.n405 B.n190 31.6883
R1729 B.n567 B.n566 31.6883
R1730 B.n732 B.n731 31.6883
R1731 B.t5 B.n172 25.6233
R1732 B.n751 B.t9 25.6233
R1733 B.n427 B.t5 22.7763
R1734 B.t9 B.n750 22.7763
R1735 B B.n812 18.0485
R1736 B.n469 B.t1 11.3884
R1737 B.n776 B.t0 11.3884
R1738 B.n401 B.n186 10.6151
R1739 B.n411 B.n186 10.6151
R1740 B.n412 B.n411 10.6151
R1741 B.n413 B.n412 10.6151
R1742 B.n413 B.n178 10.6151
R1743 B.n423 B.n178 10.6151
R1744 B.n424 B.n423 10.6151
R1745 B.n425 B.n424 10.6151
R1746 B.n425 B.n170 10.6151
R1747 B.n435 B.n170 10.6151
R1748 B.n436 B.n435 10.6151
R1749 B.n437 B.n436 10.6151
R1750 B.n437 B.n162 10.6151
R1751 B.n447 B.n162 10.6151
R1752 B.n448 B.n447 10.6151
R1753 B.n449 B.n448 10.6151
R1754 B.n449 B.n154 10.6151
R1755 B.n459 B.n154 10.6151
R1756 B.n460 B.n459 10.6151
R1757 B.n461 B.n460 10.6151
R1758 B.n461 B.n146 10.6151
R1759 B.n471 B.n146 10.6151
R1760 B.n472 B.n471 10.6151
R1761 B.n473 B.n472 10.6151
R1762 B.n473 B.n138 10.6151
R1763 B.n483 B.n138 10.6151
R1764 B.n484 B.n483 10.6151
R1765 B.n485 B.n484 10.6151
R1766 B.n485 B.n130 10.6151
R1767 B.n496 B.n130 10.6151
R1768 B.n497 B.n496 10.6151
R1769 B.n498 B.n497 10.6151
R1770 B.n498 B.n123 10.6151
R1771 B.n509 B.n123 10.6151
R1772 B.n510 B.n509 10.6151
R1773 B.n511 B.n510 10.6151
R1774 B.n511 B.n0 10.6151
R1775 B.n400 B.n399 10.6151
R1776 B.n399 B.n194 10.6151
R1777 B.n394 B.n194 10.6151
R1778 B.n394 B.n393 10.6151
R1779 B.n393 B.n196 10.6151
R1780 B.n388 B.n196 10.6151
R1781 B.n388 B.n387 10.6151
R1782 B.n387 B.n386 10.6151
R1783 B.n386 B.n198 10.6151
R1784 B.n380 B.n198 10.6151
R1785 B.n380 B.n379 10.6151
R1786 B.n379 B.n378 10.6151
R1787 B.n378 B.n200 10.6151
R1788 B.n372 B.n200 10.6151
R1789 B.n372 B.n371 10.6151
R1790 B.n371 B.n370 10.6151
R1791 B.n370 B.n202 10.6151
R1792 B.n364 B.n202 10.6151
R1793 B.n364 B.n363 10.6151
R1794 B.n363 B.n362 10.6151
R1795 B.n362 B.n204 10.6151
R1796 B.n356 B.n204 10.6151
R1797 B.n356 B.n355 10.6151
R1798 B.n355 B.n354 10.6151
R1799 B.n354 B.n206 10.6151
R1800 B.n348 B.n206 10.6151
R1801 B.n348 B.n347 10.6151
R1802 B.n347 B.n346 10.6151
R1803 B.n346 B.n208 10.6151
R1804 B.n340 B.n208 10.6151
R1805 B.n340 B.n339 10.6151
R1806 B.n339 B.n338 10.6151
R1807 B.n338 B.n210 10.6151
R1808 B.n332 B.n210 10.6151
R1809 B.n332 B.n331 10.6151
R1810 B.n329 B.n214 10.6151
R1811 B.n323 B.n214 10.6151
R1812 B.n323 B.n322 10.6151
R1813 B.n322 B.n321 10.6151
R1814 B.n321 B.n216 10.6151
R1815 B.n315 B.n216 10.6151
R1816 B.n315 B.n314 10.6151
R1817 B.n314 B.n313 10.6151
R1818 B.n313 B.n218 10.6151
R1819 B.n307 B.n306 10.6151
R1820 B.n306 B.n305 10.6151
R1821 B.n305 B.n223 10.6151
R1822 B.n299 B.n223 10.6151
R1823 B.n299 B.n298 10.6151
R1824 B.n298 B.n297 10.6151
R1825 B.n297 B.n225 10.6151
R1826 B.n291 B.n225 10.6151
R1827 B.n291 B.n290 10.6151
R1828 B.n290 B.n289 10.6151
R1829 B.n289 B.n227 10.6151
R1830 B.n283 B.n227 10.6151
R1831 B.n283 B.n282 10.6151
R1832 B.n282 B.n281 10.6151
R1833 B.n281 B.n229 10.6151
R1834 B.n275 B.n229 10.6151
R1835 B.n275 B.n274 10.6151
R1836 B.n274 B.n273 10.6151
R1837 B.n273 B.n231 10.6151
R1838 B.n267 B.n231 10.6151
R1839 B.n267 B.n266 10.6151
R1840 B.n266 B.n265 10.6151
R1841 B.n265 B.n233 10.6151
R1842 B.n259 B.n233 10.6151
R1843 B.n259 B.n258 10.6151
R1844 B.n258 B.n257 10.6151
R1845 B.n257 B.n235 10.6151
R1846 B.n251 B.n235 10.6151
R1847 B.n251 B.n250 10.6151
R1848 B.n250 B.n249 10.6151
R1849 B.n249 B.n237 10.6151
R1850 B.n243 B.n237 10.6151
R1851 B.n243 B.n242 10.6151
R1852 B.n242 B.n241 10.6151
R1853 B.n241 B.n190 10.6151
R1854 B.n406 B.n405 10.6151
R1855 B.n407 B.n406 10.6151
R1856 B.n407 B.n182 10.6151
R1857 B.n417 B.n182 10.6151
R1858 B.n418 B.n417 10.6151
R1859 B.n419 B.n418 10.6151
R1860 B.n419 B.n174 10.6151
R1861 B.n429 B.n174 10.6151
R1862 B.n430 B.n429 10.6151
R1863 B.n431 B.n430 10.6151
R1864 B.n431 B.n166 10.6151
R1865 B.n441 B.n166 10.6151
R1866 B.n442 B.n441 10.6151
R1867 B.n443 B.n442 10.6151
R1868 B.n443 B.n158 10.6151
R1869 B.n453 B.n158 10.6151
R1870 B.n454 B.n453 10.6151
R1871 B.n455 B.n454 10.6151
R1872 B.n455 B.n149 10.6151
R1873 B.n465 B.n149 10.6151
R1874 B.n466 B.n465 10.6151
R1875 B.n467 B.n466 10.6151
R1876 B.n467 B.n142 10.6151
R1877 B.n477 B.n142 10.6151
R1878 B.n478 B.n477 10.6151
R1879 B.n479 B.n478 10.6151
R1880 B.n479 B.n134 10.6151
R1881 B.n489 B.n134 10.6151
R1882 B.n490 B.n489 10.6151
R1883 B.n491 B.n490 10.6151
R1884 B.n491 B.n127 10.6151
R1885 B.n502 B.n127 10.6151
R1886 B.n503 B.n502 10.6151
R1887 B.n505 B.n503 10.6151
R1888 B.n505 B.n504 10.6151
R1889 B.n504 B.n119 10.6151
R1890 B.n516 B.n119 10.6151
R1891 B.n517 B.n516 10.6151
R1892 B.n518 B.n517 10.6151
R1893 B.n519 B.n518 10.6151
R1894 B.n520 B.n519 10.6151
R1895 B.n523 B.n520 10.6151
R1896 B.n524 B.n523 10.6151
R1897 B.n525 B.n524 10.6151
R1898 B.n526 B.n525 10.6151
R1899 B.n528 B.n526 10.6151
R1900 B.n529 B.n528 10.6151
R1901 B.n530 B.n529 10.6151
R1902 B.n531 B.n530 10.6151
R1903 B.n533 B.n531 10.6151
R1904 B.n534 B.n533 10.6151
R1905 B.n535 B.n534 10.6151
R1906 B.n536 B.n535 10.6151
R1907 B.n538 B.n536 10.6151
R1908 B.n539 B.n538 10.6151
R1909 B.n540 B.n539 10.6151
R1910 B.n541 B.n540 10.6151
R1911 B.n543 B.n541 10.6151
R1912 B.n544 B.n543 10.6151
R1913 B.n545 B.n544 10.6151
R1914 B.n546 B.n545 10.6151
R1915 B.n548 B.n546 10.6151
R1916 B.n549 B.n548 10.6151
R1917 B.n550 B.n549 10.6151
R1918 B.n551 B.n550 10.6151
R1919 B.n553 B.n551 10.6151
R1920 B.n554 B.n553 10.6151
R1921 B.n555 B.n554 10.6151
R1922 B.n556 B.n555 10.6151
R1923 B.n558 B.n556 10.6151
R1924 B.n559 B.n558 10.6151
R1925 B.n560 B.n559 10.6151
R1926 B.n561 B.n560 10.6151
R1927 B.n563 B.n561 10.6151
R1928 B.n564 B.n563 10.6151
R1929 B.n565 B.n564 10.6151
R1930 B.n566 B.n565 10.6151
R1931 B.n804 B.n1 10.6151
R1932 B.n804 B.n803 10.6151
R1933 B.n803 B.n802 10.6151
R1934 B.n802 B.n10 10.6151
R1935 B.n796 B.n10 10.6151
R1936 B.n796 B.n795 10.6151
R1937 B.n795 B.n794 10.6151
R1938 B.n794 B.n17 10.6151
R1939 B.n788 B.n17 10.6151
R1940 B.n788 B.n787 10.6151
R1941 B.n787 B.n786 10.6151
R1942 B.n786 B.n25 10.6151
R1943 B.n780 B.n25 10.6151
R1944 B.n780 B.n779 10.6151
R1945 B.n779 B.n778 10.6151
R1946 B.n778 B.n32 10.6151
R1947 B.n772 B.n32 10.6151
R1948 B.n772 B.n771 10.6151
R1949 B.n771 B.n770 10.6151
R1950 B.n770 B.n39 10.6151
R1951 B.n764 B.n39 10.6151
R1952 B.n764 B.n763 10.6151
R1953 B.n763 B.n762 10.6151
R1954 B.n762 B.n46 10.6151
R1955 B.n756 B.n46 10.6151
R1956 B.n756 B.n755 10.6151
R1957 B.n755 B.n754 10.6151
R1958 B.n754 B.n53 10.6151
R1959 B.n748 B.n53 10.6151
R1960 B.n748 B.n747 10.6151
R1961 B.n747 B.n746 10.6151
R1962 B.n746 B.n60 10.6151
R1963 B.n740 B.n60 10.6151
R1964 B.n740 B.n739 10.6151
R1965 B.n739 B.n738 10.6151
R1966 B.n738 B.n67 10.6151
R1967 B.n732 B.n67 10.6151
R1968 B.n731 B.n730 10.6151
R1969 B.n730 B.n74 10.6151
R1970 B.n724 B.n74 10.6151
R1971 B.n724 B.n723 10.6151
R1972 B.n723 B.n722 10.6151
R1973 B.n722 B.n76 10.6151
R1974 B.n716 B.n76 10.6151
R1975 B.n716 B.n715 10.6151
R1976 B.n715 B.n714 10.6151
R1977 B.n714 B.n78 10.6151
R1978 B.n708 B.n78 10.6151
R1979 B.n708 B.n707 10.6151
R1980 B.n707 B.n706 10.6151
R1981 B.n706 B.n80 10.6151
R1982 B.n700 B.n80 10.6151
R1983 B.n700 B.n699 10.6151
R1984 B.n699 B.n698 10.6151
R1985 B.n698 B.n82 10.6151
R1986 B.n692 B.n82 10.6151
R1987 B.n692 B.n691 10.6151
R1988 B.n691 B.n690 10.6151
R1989 B.n690 B.n84 10.6151
R1990 B.n684 B.n84 10.6151
R1991 B.n684 B.n683 10.6151
R1992 B.n683 B.n682 10.6151
R1993 B.n682 B.n86 10.6151
R1994 B.n676 B.n86 10.6151
R1995 B.n676 B.n675 10.6151
R1996 B.n675 B.n674 10.6151
R1997 B.n674 B.n88 10.6151
R1998 B.n668 B.n88 10.6151
R1999 B.n668 B.n667 10.6151
R2000 B.n667 B.n666 10.6151
R2001 B.n666 B.n90 10.6151
R2002 B.n660 B.n90 10.6151
R2003 B.n658 B.n657 10.6151
R2004 B.n657 B.n94 10.6151
R2005 B.n651 B.n94 10.6151
R2006 B.n651 B.n650 10.6151
R2007 B.n650 B.n649 10.6151
R2008 B.n649 B.n96 10.6151
R2009 B.n643 B.n96 10.6151
R2010 B.n643 B.n642 10.6151
R2011 B.n642 B.n641 10.6151
R2012 B.n637 B.n636 10.6151
R2013 B.n636 B.n102 10.6151
R2014 B.n631 B.n102 10.6151
R2015 B.n631 B.n630 10.6151
R2016 B.n630 B.n629 10.6151
R2017 B.n629 B.n104 10.6151
R2018 B.n623 B.n104 10.6151
R2019 B.n623 B.n622 10.6151
R2020 B.n622 B.n621 10.6151
R2021 B.n621 B.n106 10.6151
R2022 B.n615 B.n106 10.6151
R2023 B.n615 B.n614 10.6151
R2024 B.n614 B.n613 10.6151
R2025 B.n613 B.n108 10.6151
R2026 B.n607 B.n108 10.6151
R2027 B.n607 B.n606 10.6151
R2028 B.n606 B.n605 10.6151
R2029 B.n605 B.n110 10.6151
R2030 B.n599 B.n110 10.6151
R2031 B.n599 B.n598 10.6151
R2032 B.n598 B.n597 10.6151
R2033 B.n597 B.n112 10.6151
R2034 B.n591 B.n112 10.6151
R2035 B.n591 B.n590 10.6151
R2036 B.n590 B.n589 10.6151
R2037 B.n589 B.n114 10.6151
R2038 B.n583 B.n114 10.6151
R2039 B.n583 B.n582 10.6151
R2040 B.n582 B.n581 10.6151
R2041 B.n581 B.n116 10.6151
R2042 B.n575 B.n116 10.6151
R2043 B.n575 B.n574 10.6151
R2044 B.n574 B.n573 10.6151
R2045 B.n573 B.n118 10.6151
R2046 B.n567 B.n118 10.6151
R2047 B.n331 B.n330 9.36635
R2048 B.n307 B.n222 9.36635
R2049 B.n660 B.n659 9.36635
R2050 B.n637 B.n100 9.36635
R2051 B.n812 B.n0 8.11757
R2052 B.n812 B.n1 8.11757
R2053 B.n500 B.t2 7.11794
R2054 B.n798 B.t3 7.11794
R2055 B.n330 B.n329 1.24928
R2056 B.n222 B.n218 1.24928
R2057 B.n659 B.n658 1.24928
R2058 B.n641 B.n100 1.24928
R2059 VP.n15 VP.n14 161.3
R2060 VP.n13 VP.n1 161.3
R2061 VP.n12 VP.n11 161.3
R2062 VP.n10 VP.n2 161.3
R2063 VP.n9 VP.n8 161.3
R2064 VP.n7 VP.n3 161.3
R2065 VP.n4 VP.t0 113.725
R2066 VP.n4 VP.t3 112.71
R2067 VP.n6 VP.t2 79.1418
R2068 VP.n0 VP.t1 79.1418
R2069 VP.n6 VP.n5 67.3751
R2070 VP.n16 VP.n0 67.3751
R2071 VP.n12 VP.n2 56.5617
R2072 VP.n5 VP.n4 49.4013
R2073 VP.n8 VP.n7 24.5923
R2074 VP.n8 VP.n2 24.5923
R2075 VP.n13 VP.n12 24.5923
R2076 VP.n14 VP.n13 24.5923
R2077 VP.n7 VP.n6 22.8709
R2078 VP.n14 VP.n0 22.8709
R2079 VP.n5 VP.n3 0.354861
R2080 VP.n16 VP.n15 0.354861
R2081 VP VP.n16 0.267071
R2082 VP.n9 VP.n3 0.189894
R2083 VP.n10 VP.n9 0.189894
R2084 VP.n11 VP.n10 0.189894
R2085 VP.n11 VP.n1 0.189894
R2086 VP.n15 VP.n1 0.189894
R2087 VDD1 VDD1.n1 108.793
R2088 VDD1 VDD1.n0 66.965
R2089 VDD1.n0 VDD1.t3 1.94549
R2090 VDD1.n0 VDD1.t0 1.94549
R2091 VDD1.n1 VDD1.t1 1.94549
R2092 VDD1.n1 VDD1.t2 1.94549
C0 VP VTAIL 4.28089f
C1 VDD1 VDD2 1.14914f
C2 VDD1 VN 0.149929f
C3 VN VDD2 4.19446f
C4 VDD1 VTAIL 5.11105f
C5 VDD1 VP 4.47027f
C6 VTAIL VDD2 5.16861f
C7 VP VDD2 0.426598f
C8 VTAIL VN 4.26678f
C9 VP VN 6.2084f
C10 VDD2 B 3.913343f
C11 VDD1 B 8.09246f
C12 VTAIL B 9.256787f
C13 VN B 11.50516f
C14 VP B 9.881944f
C15 VDD1.t3 B 0.221981f
C16 VDD1.t0 B 0.221981f
C17 VDD1.n0 B 1.96113f
C18 VDD1.t1 B 0.221981f
C19 VDD1.t2 B 0.221981f
C20 VDD1.n1 B 2.60694f
C21 VP.t1 B 2.04546f
C22 VP.n0 B 0.828236f
C23 VP.n1 B 0.023911f
C24 VP.n2 B 0.034758f
C25 VP.n3 B 0.038586f
C26 VP.t2 B 2.04546f
C27 VP.t0 B 2.32023f
C28 VP.t3 B 2.31248f
C29 VP.n4 B 2.7821f
C30 VP.n5 B 1.32188f
C31 VP.n6 B 0.828236f
C32 VP.n7 B 0.042808f
C33 VP.n8 B 0.044341f
C34 VP.n9 B 0.023911f
C35 VP.n10 B 0.023911f
C36 VP.n11 B 0.023911f
C37 VP.n12 B 0.034758f
C38 VP.n13 B 0.044341f
C39 VP.n14 B 0.042808f
C40 VP.n15 B 0.038586f
C41 VP.n16 B 0.047231f
C42 VTAIL.n0 B 0.025655f
C43 VTAIL.n1 B 0.017416f
C44 VTAIL.n2 B 0.009359f
C45 VTAIL.n3 B 0.022121f
C46 VTAIL.n4 B 0.009909f
C47 VTAIL.n5 B 0.017416f
C48 VTAIL.n6 B 0.009634f
C49 VTAIL.n7 B 0.022121f
C50 VTAIL.n8 B 0.009909f
C51 VTAIL.n9 B 0.017416f
C52 VTAIL.n10 B 0.009359f
C53 VTAIL.n11 B 0.022121f
C54 VTAIL.n12 B 0.009909f
C55 VTAIL.n13 B 0.017416f
C56 VTAIL.n14 B 0.009359f
C57 VTAIL.n15 B 0.016591f
C58 VTAIL.n16 B 0.015638f
C59 VTAIL.t6 B 0.037191f
C60 VTAIL.n17 B 0.113403f
C61 VTAIL.n18 B 0.737626f
C62 VTAIL.n19 B 0.009359f
C63 VTAIL.n20 B 0.009909f
C64 VTAIL.n21 B 0.022121f
C65 VTAIL.n22 B 0.022121f
C66 VTAIL.n23 B 0.009909f
C67 VTAIL.n24 B 0.009359f
C68 VTAIL.n25 B 0.017416f
C69 VTAIL.n26 B 0.017416f
C70 VTAIL.n27 B 0.009359f
C71 VTAIL.n28 B 0.009909f
C72 VTAIL.n29 B 0.022121f
C73 VTAIL.n30 B 0.022121f
C74 VTAIL.n31 B 0.009909f
C75 VTAIL.n32 B 0.009359f
C76 VTAIL.n33 B 0.017416f
C77 VTAIL.n34 B 0.017416f
C78 VTAIL.n35 B 0.009359f
C79 VTAIL.n36 B 0.009359f
C80 VTAIL.n37 B 0.009909f
C81 VTAIL.n38 B 0.022121f
C82 VTAIL.n39 B 0.022121f
C83 VTAIL.n40 B 0.022121f
C84 VTAIL.n41 B 0.009634f
C85 VTAIL.n42 B 0.009359f
C86 VTAIL.n43 B 0.017416f
C87 VTAIL.n44 B 0.017416f
C88 VTAIL.n45 B 0.009359f
C89 VTAIL.n46 B 0.009909f
C90 VTAIL.n47 B 0.022121f
C91 VTAIL.n48 B 0.049965f
C92 VTAIL.n49 B 0.009909f
C93 VTAIL.n50 B 0.009359f
C94 VTAIL.n51 B 0.045491f
C95 VTAIL.n52 B 0.028323f
C96 VTAIL.n53 B 0.130438f
C97 VTAIL.n54 B 0.025655f
C98 VTAIL.n55 B 0.017416f
C99 VTAIL.n56 B 0.009359f
C100 VTAIL.n57 B 0.022121f
C101 VTAIL.n58 B 0.009909f
C102 VTAIL.n59 B 0.017416f
C103 VTAIL.n60 B 0.009634f
C104 VTAIL.n61 B 0.022121f
C105 VTAIL.n62 B 0.009909f
C106 VTAIL.n63 B 0.017416f
C107 VTAIL.n64 B 0.009359f
C108 VTAIL.n65 B 0.022121f
C109 VTAIL.n66 B 0.009909f
C110 VTAIL.n67 B 0.017416f
C111 VTAIL.n68 B 0.009359f
C112 VTAIL.n69 B 0.016591f
C113 VTAIL.n70 B 0.015638f
C114 VTAIL.t2 B 0.037191f
C115 VTAIL.n71 B 0.113403f
C116 VTAIL.n72 B 0.737626f
C117 VTAIL.n73 B 0.009359f
C118 VTAIL.n74 B 0.009909f
C119 VTAIL.n75 B 0.022121f
C120 VTAIL.n76 B 0.022121f
C121 VTAIL.n77 B 0.009909f
C122 VTAIL.n78 B 0.009359f
C123 VTAIL.n79 B 0.017416f
C124 VTAIL.n80 B 0.017416f
C125 VTAIL.n81 B 0.009359f
C126 VTAIL.n82 B 0.009909f
C127 VTAIL.n83 B 0.022121f
C128 VTAIL.n84 B 0.022121f
C129 VTAIL.n85 B 0.009909f
C130 VTAIL.n86 B 0.009359f
C131 VTAIL.n87 B 0.017416f
C132 VTAIL.n88 B 0.017416f
C133 VTAIL.n89 B 0.009359f
C134 VTAIL.n90 B 0.009359f
C135 VTAIL.n91 B 0.009909f
C136 VTAIL.n92 B 0.022121f
C137 VTAIL.n93 B 0.022121f
C138 VTAIL.n94 B 0.022121f
C139 VTAIL.n95 B 0.009634f
C140 VTAIL.n96 B 0.009359f
C141 VTAIL.n97 B 0.017416f
C142 VTAIL.n98 B 0.017416f
C143 VTAIL.n99 B 0.009359f
C144 VTAIL.n100 B 0.009909f
C145 VTAIL.n101 B 0.022121f
C146 VTAIL.n102 B 0.049965f
C147 VTAIL.n103 B 0.009909f
C148 VTAIL.n104 B 0.009359f
C149 VTAIL.n105 B 0.045491f
C150 VTAIL.n106 B 0.028323f
C151 VTAIL.n107 B 0.210142f
C152 VTAIL.n108 B 0.025655f
C153 VTAIL.n109 B 0.017416f
C154 VTAIL.n110 B 0.009359f
C155 VTAIL.n111 B 0.022121f
C156 VTAIL.n112 B 0.009909f
C157 VTAIL.n113 B 0.017416f
C158 VTAIL.n114 B 0.009634f
C159 VTAIL.n115 B 0.022121f
C160 VTAIL.n116 B 0.009909f
C161 VTAIL.n117 B 0.017416f
C162 VTAIL.n118 B 0.009359f
C163 VTAIL.n119 B 0.022121f
C164 VTAIL.n120 B 0.009909f
C165 VTAIL.n121 B 0.017416f
C166 VTAIL.n122 B 0.009359f
C167 VTAIL.n123 B 0.016591f
C168 VTAIL.n124 B 0.015638f
C169 VTAIL.t1 B 0.037191f
C170 VTAIL.n125 B 0.113403f
C171 VTAIL.n126 B 0.737626f
C172 VTAIL.n127 B 0.009359f
C173 VTAIL.n128 B 0.009909f
C174 VTAIL.n129 B 0.022121f
C175 VTAIL.n130 B 0.022121f
C176 VTAIL.n131 B 0.009909f
C177 VTAIL.n132 B 0.009359f
C178 VTAIL.n133 B 0.017416f
C179 VTAIL.n134 B 0.017416f
C180 VTAIL.n135 B 0.009359f
C181 VTAIL.n136 B 0.009909f
C182 VTAIL.n137 B 0.022121f
C183 VTAIL.n138 B 0.022121f
C184 VTAIL.n139 B 0.009909f
C185 VTAIL.n140 B 0.009359f
C186 VTAIL.n141 B 0.017416f
C187 VTAIL.n142 B 0.017416f
C188 VTAIL.n143 B 0.009359f
C189 VTAIL.n144 B 0.009359f
C190 VTAIL.n145 B 0.009909f
C191 VTAIL.n146 B 0.022121f
C192 VTAIL.n147 B 0.022121f
C193 VTAIL.n148 B 0.022121f
C194 VTAIL.n149 B 0.009634f
C195 VTAIL.n150 B 0.009359f
C196 VTAIL.n151 B 0.017416f
C197 VTAIL.n152 B 0.017416f
C198 VTAIL.n153 B 0.009359f
C199 VTAIL.n154 B 0.009909f
C200 VTAIL.n155 B 0.022121f
C201 VTAIL.n156 B 0.049965f
C202 VTAIL.n157 B 0.009909f
C203 VTAIL.n158 B 0.009359f
C204 VTAIL.n159 B 0.045491f
C205 VTAIL.n160 B 0.028323f
C206 VTAIL.n161 B 1.07878f
C207 VTAIL.n162 B 0.025655f
C208 VTAIL.n163 B 0.017416f
C209 VTAIL.n164 B 0.009359f
C210 VTAIL.n165 B 0.022121f
C211 VTAIL.n166 B 0.009909f
C212 VTAIL.n167 B 0.017416f
C213 VTAIL.n168 B 0.009634f
C214 VTAIL.n169 B 0.022121f
C215 VTAIL.n170 B 0.009359f
C216 VTAIL.n171 B 0.009909f
C217 VTAIL.n172 B 0.017416f
C218 VTAIL.n173 B 0.009359f
C219 VTAIL.n174 B 0.022121f
C220 VTAIL.n175 B 0.009909f
C221 VTAIL.n176 B 0.017416f
C222 VTAIL.n177 B 0.009359f
C223 VTAIL.n178 B 0.016591f
C224 VTAIL.n179 B 0.015638f
C225 VTAIL.t7 B 0.037191f
C226 VTAIL.n180 B 0.113403f
C227 VTAIL.n181 B 0.737626f
C228 VTAIL.n182 B 0.009359f
C229 VTAIL.n183 B 0.009909f
C230 VTAIL.n184 B 0.022121f
C231 VTAIL.n185 B 0.022121f
C232 VTAIL.n186 B 0.009909f
C233 VTAIL.n187 B 0.009359f
C234 VTAIL.n188 B 0.017416f
C235 VTAIL.n189 B 0.017416f
C236 VTAIL.n190 B 0.009359f
C237 VTAIL.n191 B 0.009909f
C238 VTAIL.n192 B 0.022121f
C239 VTAIL.n193 B 0.022121f
C240 VTAIL.n194 B 0.009909f
C241 VTAIL.n195 B 0.009359f
C242 VTAIL.n196 B 0.017416f
C243 VTAIL.n197 B 0.017416f
C244 VTAIL.n198 B 0.009359f
C245 VTAIL.n199 B 0.009909f
C246 VTAIL.n200 B 0.022121f
C247 VTAIL.n201 B 0.022121f
C248 VTAIL.n202 B 0.022121f
C249 VTAIL.n203 B 0.009634f
C250 VTAIL.n204 B 0.009359f
C251 VTAIL.n205 B 0.017416f
C252 VTAIL.n206 B 0.017416f
C253 VTAIL.n207 B 0.009359f
C254 VTAIL.n208 B 0.009909f
C255 VTAIL.n209 B 0.022121f
C256 VTAIL.n210 B 0.049965f
C257 VTAIL.n211 B 0.009909f
C258 VTAIL.n212 B 0.009359f
C259 VTAIL.n213 B 0.045491f
C260 VTAIL.n214 B 0.028323f
C261 VTAIL.n215 B 1.07878f
C262 VTAIL.n216 B 0.025655f
C263 VTAIL.n217 B 0.017416f
C264 VTAIL.n218 B 0.009359f
C265 VTAIL.n219 B 0.022121f
C266 VTAIL.n220 B 0.009909f
C267 VTAIL.n221 B 0.017416f
C268 VTAIL.n222 B 0.009634f
C269 VTAIL.n223 B 0.022121f
C270 VTAIL.n224 B 0.009359f
C271 VTAIL.n225 B 0.009909f
C272 VTAIL.n226 B 0.017416f
C273 VTAIL.n227 B 0.009359f
C274 VTAIL.n228 B 0.022121f
C275 VTAIL.n229 B 0.009909f
C276 VTAIL.n230 B 0.017416f
C277 VTAIL.n231 B 0.009359f
C278 VTAIL.n232 B 0.016591f
C279 VTAIL.n233 B 0.015638f
C280 VTAIL.t4 B 0.037191f
C281 VTAIL.n234 B 0.113403f
C282 VTAIL.n235 B 0.737626f
C283 VTAIL.n236 B 0.009359f
C284 VTAIL.n237 B 0.009909f
C285 VTAIL.n238 B 0.022121f
C286 VTAIL.n239 B 0.022121f
C287 VTAIL.n240 B 0.009909f
C288 VTAIL.n241 B 0.009359f
C289 VTAIL.n242 B 0.017416f
C290 VTAIL.n243 B 0.017416f
C291 VTAIL.n244 B 0.009359f
C292 VTAIL.n245 B 0.009909f
C293 VTAIL.n246 B 0.022121f
C294 VTAIL.n247 B 0.022121f
C295 VTAIL.n248 B 0.009909f
C296 VTAIL.n249 B 0.009359f
C297 VTAIL.n250 B 0.017416f
C298 VTAIL.n251 B 0.017416f
C299 VTAIL.n252 B 0.009359f
C300 VTAIL.n253 B 0.009909f
C301 VTAIL.n254 B 0.022121f
C302 VTAIL.n255 B 0.022121f
C303 VTAIL.n256 B 0.022121f
C304 VTAIL.n257 B 0.009634f
C305 VTAIL.n258 B 0.009359f
C306 VTAIL.n259 B 0.017416f
C307 VTAIL.n260 B 0.017416f
C308 VTAIL.n261 B 0.009359f
C309 VTAIL.n262 B 0.009909f
C310 VTAIL.n263 B 0.022121f
C311 VTAIL.n264 B 0.049965f
C312 VTAIL.n265 B 0.009909f
C313 VTAIL.n266 B 0.009359f
C314 VTAIL.n267 B 0.045491f
C315 VTAIL.n268 B 0.028323f
C316 VTAIL.n269 B 0.210142f
C317 VTAIL.n270 B 0.025655f
C318 VTAIL.n271 B 0.017416f
C319 VTAIL.n272 B 0.009359f
C320 VTAIL.n273 B 0.022121f
C321 VTAIL.n274 B 0.009909f
C322 VTAIL.n275 B 0.017416f
C323 VTAIL.n276 B 0.009634f
C324 VTAIL.n277 B 0.022121f
C325 VTAIL.n278 B 0.009359f
C326 VTAIL.n279 B 0.009909f
C327 VTAIL.n280 B 0.017416f
C328 VTAIL.n281 B 0.009359f
C329 VTAIL.n282 B 0.022121f
C330 VTAIL.n283 B 0.009909f
C331 VTAIL.n284 B 0.017416f
C332 VTAIL.n285 B 0.009359f
C333 VTAIL.n286 B 0.016591f
C334 VTAIL.n287 B 0.015638f
C335 VTAIL.t3 B 0.037191f
C336 VTAIL.n288 B 0.113403f
C337 VTAIL.n289 B 0.737626f
C338 VTAIL.n290 B 0.009359f
C339 VTAIL.n291 B 0.009909f
C340 VTAIL.n292 B 0.022121f
C341 VTAIL.n293 B 0.022121f
C342 VTAIL.n294 B 0.009909f
C343 VTAIL.n295 B 0.009359f
C344 VTAIL.n296 B 0.017416f
C345 VTAIL.n297 B 0.017416f
C346 VTAIL.n298 B 0.009359f
C347 VTAIL.n299 B 0.009909f
C348 VTAIL.n300 B 0.022121f
C349 VTAIL.n301 B 0.022121f
C350 VTAIL.n302 B 0.009909f
C351 VTAIL.n303 B 0.009359f
C352 VTAIL.n304 B 0.017416f
C353 VTAIL.n305 B 0.017416f
C354 VTAIL.n306 B 0.009359f
C355 VTAIL.n307 B 0.009909f
C356 VTAIL.n308 B 0.022121f
C357 VTAIL.n309 B 0.022121f
C358 VTAIL.n310 B 0.022121f
C359 VTAIL.n311 B 0.009634f
C360 VTAIL.n312 B 0.009359f
C361 VTAIL.n313 B 0.017416f
C362 VTAIL.n314 B 0.017416f
C363 VTAIL.n315 B 0.009359f
C364 VTAIL.n316 B 0.009909f
C365 VTAIL.n317 B 0.022121f
C366 VTAIL.n318 B 0.049965f
C367 VTAIL.n319 B 0.009909f
C368 VTAIL.n320 B 0.009359f
C369 VTAIL.n321 B 0.045491f
C370 VTAIL.n322 B 0.028323f
C371 VTAIL.n323 B 0.210142f
C372 VTAIL.n324 B 0.025655f
C373 VTAIL.n325 B 0.017416f
C374 VTAIL.n326 B 0.009359f
C375 VTAIL.n327 B 0.022121f
C376 VTAIL.n328 B 0.009909f
C377 VTAIL.n329 B 0.017416f
C378 VTAIL.n330 B 0.009634f
C379 VTAIL.n331 B 0.022121f
C380 VTAIL.n332 B 0.009359f
C381 VTAIL.n333 B 0.009909f
C382 VTAIL.n334 B 0.017416f
C383 VTAIL.n335 B 0.009359f
C384 VTAIL.n336 B 0.022121f
C385 VTAIL.n337 B 0.009909f
C386 VTAIL.n338 B 0.017416f
C387 VTAIL.n339 B 0.009359f
C388 VTAIL.n340 B 0.016591f
C389 VTAIL.n341 B 0.015638f
C390 VTAIL.t0 B 0.037191f
C391 VTAIL.n342 B 0.113403f
C392 VTAIL.n343 B 0.737626f
C393 VTAIL.n344 B 0.009359f
C394 VTAIL.n345 B 0.009909f
C395 VTAIL.n346 B 0.022121f
C396 VTAIL.n347 B 0.022121f
C397 VTAIL.n348 B 0.009909f
C398 VTAIL.n349 B 0.009359f
C399 VTAIL.n350 B 0.017416f
C400 VTAIL.n351 B 0.017416f
C401 VTAIL.n352 B 0.009359f
C402 VTAIL.n353 B 0.009909f
C403 VTAIL.n354 B 0.022121f
C404 VTAIL.n355 B 0.022121f
C405 VTAIL.n356 B 0.009909f
C406 VTAIL.n357 B 0.009359f
C407 VTAIL.n358 B 0.017416f
C408 VTAIL.n359 B 0.017416f
C409 VTAIL.n360 B 0.009359f
C410 VTAIL.n361 B 0.009909f
C411 VTAIL.n362 B 0.022121f
C412 VTAIL.n363 B 0.022121f
C413 VTAIL.n364 B 0.022121f
C414 VTAIL.n365 B 0.009634f
C415 VTAIL.n366 B 0.009359f
C416 VTAIL.n367 B 0.017416f
C417 VTAIL.n368 B 0.017416f
C418 VTAIL.n369 B 0.009359f
C419 VTAIL.n370 B 0.009909f
C420 VTAIL.n371 B 0.022121f
C421 VTAIL.n372 B 0.049965f
C422 VTAIL.n373 B 0.009909f
C423 VTAIL.n374 B 0.009359f
C424 VTAIL.n375 B 0.045491f
C425 VTAIL.n376 B 0.028323f
C426 VTAIL.n377 B 1.07878f
C427 VTAIL.n378 B 0.025655f
C428 VTAIL.n379 B 0.017416f
C429 VTAIL.n380 B 0.009359f
C430 VTAIL.n381 B 0.022121f
C431 VTAIL.n382 B 0.009909f
C432 VTAIL.n383 B 0.017416f
C433 VTAIL.n384 B 0.009634f
C434 VTAIL.n385 B 0.022121f
C435 VTAIL.n386 B 0.009909f
C436 VTAIL.n387 B 0.017416f
C437 VTAIL.n388 B 0.009359f
C438 VTAIL.n389 B 0.022121f
C439 VTAIL.n390 B 0.009909f
C440 VTAIL.n391 B 0.017416f
C441 VTAIL.n392 B 0.009359f
C442 VTAIL.n393 B 0.016591f
C443 VTAIL.n394 B 0.015638f
C444 VTAIL.t5 B 0.037191f
C445 VTAIL.n395 B 0.113403f
C446 VTAIL.n396 B 0.737626f
C447 VTAIL.n397 B 0.009359f
C448 VTAIL.n398 B 0.009909f
C449 VTAIL.n399 B 0.022121f
C450 VTAIL.n400 B 0.022121f
C451 VTAIL.n401 B 0.009909f
C452 VTAIL.n402 B 0.009359f
C453 VTAIL.n403 B 0.017416f
C454 VTAIL.n404 B 0.017416f
C455 VTAIL.n405 B 0.009359f
C456 VTAIL.n406 B 0.009909f
C457 VTAIL.n407 B 0.022121f
C458 VTAIL.n408 B 0.022121f
C459 VTAIL.n409 B 0.009909f
C460 VTAIL.n410 B 0.009359f
C461 VTAIL.n411 B 0.017416f
C462 VTAIL.n412 B 0.017416f
C463 VTAIL.n413 B 0.009359f
C464 VTAIL.n414 B 0.009359f
C465 VTAIL.n415 B 0.009909f
C466 VTAIL.n416 B 0.022121f
C467 VTAIL.n417 B 0.022121f
C468 VTAIL.n418 B 0.022121f
C469 VTAIL.n419 B 0.009634f
C470 VTAIL.n420 B 0.009359f
C471 VTAIL.n421 B 0.017416f
C472 VTAIL.n422 B 0.017416f
C473 VTAIL.n423 B 0.009359f
C474 VTAIL.n424 B 0.009909f
C475 VTAIL.n425 B 0.022121f
C476 VTAIL.n426 B 0.049965f
C477 VTAIL.n427 B 0.009909f
C478 VTAIL.n428 B 0.009359f
C479 VTAIL.n429 B 0.045491f
C480 VTAIL.n430 B 0.028323f
C481 VTAIL.n431 B 0.99255f
C482 VDD2.t3 B 0.219688f
C483 VDD2.t2 B 0.219688f
C484 VDD2.n0 B 2.55434f
C485 VDD2.t1 B 0.219688f
C486 VDD2.t0 B 0.219688f
C487 VDD2.n1 B 1.94045f
C488 VDD2.n2 B 3.76039f
C489 VN.t2 B 2.26116f
C490 VN.t1 B 2.26874f
C491 VN.n0 B 1.38392f
C492 VN.t3 B 2.26874f
C493 VN.t0 B 2.26116f
C494 VN.n1 B 2.72988f
.ends

