* NGSPICE file created from diff_pair_sample_0842.ext - technology: sky130A

.subckt diff_pair_sample_0842 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.4056 ps=2.86 w=1.04 l=2.89
X1 B.t11 B.t9 B.t10 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0 ps=0 w=1.04 l=2.89
X2 VTAIL.t0 VN.t0 VDD2.t7 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0.1716 ps=1.37 w=1.04 l=2.89
X3 VDD1.t6 VP.t1 VTAIL.t9 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.4056 ps=2.86 w=1.04 l=2.89
X4 VDD2.t6 VN.t1 VTAIL.t1 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.4056 ps=2.86 w=1.04 l=2.89
X5 VDD2.t5 VN.t2 VTAIL.t7 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X6 VTAIL.t6 VN.t3 VDD2.t4 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X7 VTAIL.t8 VP.t2 VDD1.t5 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0.1716 ps=1.37 w=1.04 l=2.89
X8 VTAIL.t14 VP.t3 VDD1.t4 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X9 VDD2.t3 VN.t4 VTAIL.t3 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.4056 ps=2.86 w=1.04 l=2.89
X10 VTAIL.t10 VP.t4 VDD1.t3 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X11 VDD1.t2 VP.t5 VTAIL.t12 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X12 VDD2.t2 VN.t5 VTAIL.t2 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X13 VTAIL.t5 VN.t6 VDD2.t1 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0.1716 ps=1.37 w=1.04 l=2.89
X14 B.t8 B.t6 B.t7 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0 ps=0 w=1.04 l=2.89
X15 VTAIL.t15 VP.t6 VDD1.t1 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0.1716 ps=1.37 w=1.04 l=2.89
X16 VTAIL.t4 VN.t7 VDD2.t0 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X17 VDD1.t0 VP.t7 VTAIL.t13 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.1716 pd=1.37 as=0.1716 ps=1.37 w=1.04 l=2.89
X18 B.t5 B.t3 B.t4 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0 ps=0 w=1.04 l=2.89
X19 B.t2 B.t0 B.t1 w_n4190_n1176# sky130_fd_pr__pfet_01v8 ad=0.4056 pd=2.86 as=0 ps=0 w=1.04 l=2.89
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n28 VP.n27 161.3
R6 VP.n29 VP.n13 161.3
R7 VP.n31 VP.n30 161.3
R8 VP.n32 VP.n12 161.3
R9 VP.n34 VP.n33 161.3
R10 VP.n35 VP.n11 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n38 VP.n10 161.3
R13 VP.n74 VP.n0 161.3
R14 VP.n73 VP.n72 161.3
R15 VP.n71 VP.n1 161.3
R16 VP.n70 VP.n69 161.3
R17 VP.n68 VP.n2 161.3
R18 VP.n67 VP.n66 161.3
R19 VP.n65 VP.n3 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n53 VP.n52 161.3
R27 VP.n51 VP.n7 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n8 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n45 VP.n9 161.3
R32 VP.n44 VP.n43 161.3
R33 VP.n42 VP.n41 106.974
R34 VP.n76 VP.n75 106.974
R35 VP.n40 VP.n39 106.974
R36 VP.n60 VP.n5 56.5617
R37 VP.n24 VP.n15 56.5617
R38 VP.n18 VP.n17 56.2048
R39 VP.n41 VP.n40 43.9466
R40 VP.n49 VP.n48 43.4833
R41 VP.n69 VP.n68 43.4833
R42 VP.n33 VP.n32 43.4833
R43 VP.n17 VP.t6 42.2769
R44 VP.n48 VP.n47 37.6707
R45 VP.n69 VP.n1 37.6707
R46 VP.n33 VP.n11 37.6707
R47 VP.n43 VP.n9 24.5923
R48 VP.n47 VP.n9 24.5923
R49 VP.n49 VP.n7 24.5923
R50 VP.n53 VP.n7 24.5923
R51 VP.n56 VP.n55 24.5923
R52 VP.n56 VP.n5 24.5923
R53 VP.n61 VP.n60 24.5923
R54 VP.n63 VP.n61 24.5923
R55 VP.n67 VP.n3 24.5923
R56 VP.n68 VP.n67 24.5923
R57 VP.n73 VP.n1 24.5923
R58 VP.n74 VP.n73 24.5923
R59 VP.n37 VP.n11 24.5923
R60 VP.n38 VP.n37 24.5923
R61 VP.n25 VP.n24 24.5923
R62 VP.n27 VP.n25 24.5923
R63 VP.n31 VP.n13 24.5923
R64 VP.n32 VP.n31 24.5923
R65 VP.n20 VP.n19 24.5923
R66 VP.n20 VP.n15 24.5923
R67 VP.n55 VP.n54 17.7066
R68 VP.n63 VP.n62 17.7066
R69 VP.n27 VP.n26 17.7066
R70 VP.n19 VP.n18 17.7066
R71 VP.n42 VP.t2 8.67316
R72 VP.n54 VP.t7 8.67316
R73 VP.n62 VP.t4 8.67316
R74 VP.n75 VP.t0 8.67316
R75 VP.n39 VP.t1 8.67316
R76 VP.n26 VP.t3 8.67316
R77 VP.n18 VP.t5 8.67316
R78 VP.n54 VP.n53 6.88621
R79 VP.n62 VP.n3 6.88621
R80 VP.n26 VP.n13 6.88621
R81 VP.n17 VP.n16 5.01074
R82 VP.n43 VP.n42 3.93519
R83 VP.n75 VP.n74 3.93519
R84 VP.n39 VP.n38 3.93519
R85 VP.n40 VP.n10 0.278335
R86 VP.n44 VP.n41 0.278335
R87 VP.n76 VP.n0 0.278335
R88 VP.n21 VP.n16 0.189894
R89 VP.n22 VP.n21 0.189894
R90 VP.n23 VP.n22 0.189894
R91 VP.n23 VP.n14 0.189894
R92 VP.n28 VP.n14 0.189894
R93 VP.n29 VP.n28 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n12 0.189894
R96 VP.n34 VP.n12 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n10 0.189894
R100 VP.n45 VP.n44 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n46 VP.n8 0.189894
R103 VP.n50 VP.n8 0.189894
R104 VP.n51 VP.n50 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n52 VP.n6 0.189894
R107 VP.n57 VP.n6 0.189894
R108 VP.n58 VP.n57 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n59 VP.n4 0.189894
R111 VP.n64 VP.n4 0.189894
R112 VP.n65 VP.n64 0.189894
R113 VP.n66 VP.n65 0.189894
R114 VP.n66 VP.n2 0.189894
R115 VP.n70 VP.n2 0.189894
R116 VP.n71 VP.n70 0.189894
R117 VP.n72 VP.n71 0.189894
R118 VP.n72 VP.n0 0.189894
R119 VP VP.n76 0.153485
R120 VTAIL.n15 VTAIL.t1 371.358
R121 VTAIL.n2 VTAIL.t5 371.358
R122 VTAIL.n3 VTAIL.t11 371.358
R123 VTAIL.n6 VTAIL.t8 371.358
R124 VTAIL.n14 VTAIL.t9 371.358
R125 VTAIL.n11 VTAIL.t15 371.358
R126 VTAIL.n10 VTAIL.t3 371.358
R127 VTAIL.n7 VTAIL.t0 371.358
R128 VTAIL.n1 VTAIL.n0 328.421
R129 VTAIL.n5 VTAIL.n4 328.421
R130 VTAIL.n13 VTAIL.n12 328.421
R131 VTAIL.n9 VTAIL.n8 328.421
R132 VTAIL.n0 VTAIL.t7 31.2553
R133 VTAIL.n0 VTAIL.t4 31.2553
R134 VTAIL.n4 VTAIL.t13 31.2553
R135 VTAIL.n4 VTAIL.t10 31.2553
R136 VTAIL.n12 VTAIL.t12 31.2553
R137 VTAIL.n12 VTAIL.t14 31.2553
R138 VTAIL.n8 VTAIL.t2 31.2553
R139 VTAIL.n8 VTAIL.t6 31.2553
R140 VTAIL.n15 VTAIL.n14 16.0393
R141 VTAIL.n7 VTAIL.n6 16.0393
R142 VTAIL.n9 VTAIL.n7 2.77636
R143 VTAIL.n10 VTAIL.n9 2.77636
R144 VTAIL.n13 VTAIL.n11 2.77636
R145 VTAIL.n14 VTAIL.n13 2.77636
R146 VTAIL.n6 VTAIL.n5 2.77636
R147 VTAIL.n5 VTAIL.n3 2.77636
R148 VTAIL.n2 VTAIL.n1 2.77636
R149 VTAIL VTAIL.n15 2.71817
R150 VTAIL.n11 VTAIL.n10 0.470328
R151 VTAIL.n3 VTAIL.n2 0.470328
R152 VTAIL VTAIL.n1 0.0586897
R153 VDD1 VDD1.n0 346.546
R154 VDD1.n3 VDD1.n2 346.433
R155 VDD1.n3 VDD1.n1 346.433
R156 VDD1.n5 VDD1.n4 345.101
R157 VDD1.n5 VDD1.n3 37.6862
R158 VDD1.n4 VDD1.t4 31.2553
R159 VDD1.n4 VDD1.t6 31.2553
R160 VDD1.n0 VDD1.t1 31.2553
R161 VDD1.n0 VDD1.t2 31.2553
R162 VDD1.n2 VDD1.t3 31.2553
R163 VDD1.n2 VDD1.t7 31.2553
R164 VDD1.n1 VDD1.t5 31.2553
R165 VDD1.n1 VDD1.t0 31.2553
R166 VDD1 VDD1.n5 1.33024
R167 B.n273 B.n104 585
R168 B.n272 B.n271 585
R169 B.n270 B.n105 585
R170 B.n269 B.n268 585
R171 B.n267 B.n106 585
R172 B.n266 B.n265 585
R173 B.n264 B.n107 585
R174 B.n263 B.n262 585
R175 B.n261 B.n108 585
R176 B.n260 B.n259 585
R177 B.n255 B.n109 585
R178 B.n254 B.n253 585
R179 B.n252 B.n110 585
R180 B.n251 B.n250 585
R181 B.n249 B.n111 585
R182 B.n248 B.n247 585
R183 B.n246 B.n112 585
R184 B.n245 B.n244 585
R185 B.n243 B.n113 585
R186 B.n241 B.n240 585
R187 B.n239 B.n116 585
R188 B.n238 B.n237 585
R189 B.n236 B.n117 585
R190 B.n235 B.n234 585
R191 B.n233 B.n118 585
R192 B.n232 B.n231 585
R193 B.n230 B.n119 585
R194 B.n229 B.n228 585
R195 B.n275 B.n274 585
R196 B.n276 B.n103 585
R197 B.n278 B.n277 585
R198 B.n279 B.n102 585
R199 B.n281 B.n280 585
R200 B.n282 B.n101 585
R201 B.n284 B.n283 585
R202 B.n285 B.n100 585
R203 B.n287 B.n286 585
R204 B.n288 B.n99 585
R205 B.n290 B.n289 585
R206 B.n291 B.n98 585
R207 B.n293 B.n292 585
R208 B.n294 B.n97 585
R209 B.n296 B.n295 585
R210 B.n297 B.n96 585
R211 B.n299 B.n298 585
R212 B.n300 B.n95 585
R213 B.n302 B.n301 585
R214 B.n303 B.n94 585
R215 B.n305 B.n304 585
R216 B.n306 B.n93 585
R217 B.n308 B.n307 585
R218 B.n309 B.n92 585
R219 B.n311 B.n310 585
R220 B.n312 B.n91 585
R221 B.n314 B.n313 585
R222 B.n315 B.n90 585
R223 B.n317 B.n316 585
R224 B.n318 B.n89 585
R225 B.n320 B.n319 585
R226 B.n321 B.n88 585
R227 B.n323 B.n322 585
R228 B.n324 B.n87 585
R229 B.n326 B.n325 585
R230 B.n327 B.n86 585
R231 B.n329 B.n328 585
R232 B.n330 B.n85 585
R233 B.n332 B.n331 585
R234 B.n333 B.n84 585
R235 B.n335 B.n334 585
R236 B.n336 B.n83 585
R237 B.n338 B.n337 585
R238 B.n339 B.n82 585
R239 B.n341 B.n340 585
R240 B.n342 B.n81 585
R241 B.n344 B.n343 585
R242 B.n345 B.n80 585
R243 B.n347 B.n346 585
R244 B.n348 B.n79 585
R245 B.n350 B.n349 585
R246 B.n351 B.n78 585
R247 B.n353 B.n352 585
R248 B.n354 B.n77 585
R249 B.n356 B.n355 585
R250 B.n357 B.n76 585
R251 B.n359 B.n358 585
R252 B.n360 B.n75 585
R253 B.n362 B.n361 585
R254 B.n363 B.n74 585
R255 B.n365 B.n364 585
R256 B.n366 B.n73 585
R257 B.n368 B.n367 585
R258 B.n369 B.n72 585
R259 B.n371 B.n370 585
R260 B.n372 B.n71 585
R261 B.n374 B.n373 585
R262 B.n375 B.n70 585
R263 B.n377 B.n376 585
R264 B.n378 B.n69 585
R265 B.n380 B.n379 585
R266 B.n381 B.n68 585
R267 B.n383 B.n382 585
R268 B.n384 B.n67 585
R269 B.n386 B.n385 585
R270 B.n387 B.n66 585
R271 B.n389 B.n388 585
R272 B.n390 B.n65 585
R273 B.n392 B.n391 585
R274 B.n393 B.n64 585
R275 B.n395 B.n394 585
R276 B.n396 B.n63 585
R277 B.n398 B.n397 585
R278 B.n399 B.n62 585
R279 B.n401 B.n400 585
R280 B.n402 B.n61 585
R281 B.n404 B.n403 585
R282 B.n405 B.n60 585
R283 B.n407 B.n406 585
R284 B.n408 B.n59 585
R285 B.n410 B.n409 585
R286 B.n411 B.n58 585
R287 B.n413 B.n412 585
R288 B.n414 B.n57 585
R289 B.n416 B.n415 585
R290 B.n417 B.n56 585
R291 B.n419 B.n418 585
R292 B.n420 B.n55 585
R293 B.n422 B.n421 585
R294 B.n423 B.n54 585
R295 B.n425 B.n424 585
R296 B.n426 B.n53 585
R297 B.n428 B.n427 585
R298 B.n429 B.n52 585
R299 B.n431 B.n430 585
R300 B.n432 B.n51 585
R301 B.n434 B.n433 585
R302 B.n435 B.n50 585
R303 B.n437 B.n436 585
R304 B.n438 B.n49 585
R305 B.n440 B.n439 585
R306 B.n441 B.n48 585
R307 B.n485 B.n484 585
R308 B.n483 B.n30 585
R309 B.n482 B.n481 585
R310 B.n480 B.n31 585
R311 B.n479 B.n478 585
R312 B.n477 B.n32 585
R313 B.n476 B.n475 585
R314 B.n474 B.n33 585
R315 B.n473 B.n472 585
R316 B.n471 B.n470 585
R317 B.n469 B.n37 585
R318 B.n468 B.n467 585
R319 B.n466 B.n38 585
R320 B.n465 B.n464 585
R321 B.n463 B.n39 585
R322 B.n462 B.n461 585
R323 B.n460 B.n40 585
R324 B.n459 B.n458 585
R325 B.n457 B.n41 585
R326 B.n455 B.n454 585
R327 B.n453 B.n44 585
R328 B.n452 B.n451 585
R329 B.n450 B.n45 585
R330 B.n449 B.n448 585
R331 B.n447 B.n46 585
R332 B.n446 B.n445 585
R333 B.n444 B.n47 585
R334 B.n443 B.n442 585
R335 B.n486 B.n29 585
R336 B.n488 B.n487 585
R337 B.n489 B.n28 585
R338 B.n491 B.n490 585
R339 B.n492 B.n27 585
R340 B.n494 B.n493 585
R341 B.n495 B.n26 585
R342 B.n497 B.n496 585
R343 B.n498 B.n25 585
R344 B.n500 B.n499 585
R345 B.n501 B.n24 585
R346 B.n503 B.n502 585
R347 B.n504 B.n23 585
R348 B.n506 B.n505 585
R349 B.n507 B.n22 585
R350 B.n509 B.n508 585
R351 B.n510 B.n21 585
R352 B.n512 B.n511 585
R353 B.n513 B.n20 585
R354 B.n515 B.n514 585
R355 B.n516 B.n19 585
R356 B.n518 B.n517 585
R357 B.n519 B.n18 585
R358 B.n521 B.n520 585
R359 B.n522 B.n17 585
R360 B.n524 B.n523 585
R361 B.n525 B.n16 585
R362 B.n527 B.n526 585
R363 B.n528 B.n15 585
R364 B.n530 B.n529 585
R365 B.n531 B.n14 585
R366 B.n533 B.n532 585
R367 B.n534 B.n13 585
R368 B.n536 B.n535 585
R369 B.n537 B.n12 585
R370 B.n539 B.n538 585
R371 B.n540 B.n11 585
R372 B.n542 B.n541 585
R373 B.n543 B.n10 585
R374 B.n545 B.n544 585
R375 B.n546 B.n9 585
R376 B.n548 B.n547 585
R377 B.n549 B.n8 585
R378 B.n551 B.n550 585
R379 B.n552 B.n7 585
R380 B.n554 B.n553 585
R381 B.n555 B.n6 585
R382 B.n557 B.n556 585
R383 B.n558 B.n5 585
R384 B.n560 B.n559 585
R385 B.n561 B.n4 585
R386 B.n563 B.n562 585
R387 B.n564 B.n3 585
R388 B.n566 B.n565 585
R389 B.n567 B.n0 585
R390 B.n2 B.n1 585
R391 B.n148 B.n147 585
R392 B.n149 B.n146 585
R393 B.n151 B.n150 585
R394 B.n152 B.n145 585
R395 B.n154 B.n153 585
R396 B.n155 B.n144 585
R397 B.n157 B.n156 585
R398 B.n158 B.n143 585
R399 B.n160 B.n159 585
R400 B.n161 B.n142 585
R401 B.n163 B.n162 585
R402 B.n164 B.n141 585
R403 B.n166 B.n165 585
R404 B.n167 B.n140 585
R405 B.n169 B.n168 585
R406 B.n170 B.n139 585
R407 B.n172 B.n171 585
R408 B.n173 B.n138 585
R409 B.n175 B.n174 585
R410 B.n176 B.n137 585
R411 B.n178 B.n177 585
R412 B.n179 B.n136 585
R413 B.n181 B.n180 585
R414 B.n182 B.n135 585
R415 B.n184 B.n183 585
R416 B.n185 B.n134 585
R417 B.n187 B.n186 585
R418 B.n188 B.n133 585
R419 B.n190 B.n189 585
R420 B.n191 B.n132 585
R421 B.n193 B.n192 585
R422 B.n194 B.n131 585
R423 B.n196 B.n195 585
R424 B.n197 B.n130 585
R425 B.n199 B.n198 585
R426 B.n200 B.n129 585
R427 B.n202 B.n201 585
R428 B.n203 B.n128 585
R429 B.n205 B.n204 585
R430 B.n206 B.n127 585
R431 B.n208 B.n207 585
R432 B.n209 B.n126 585
R433 B.n211 B.n210 585
R434 B.n212 B.n125 585
R435 B.n214 B.n213 585
R436 B.n215 B.n124 585
R437 B.n217 B.n216 585
R438 B.n218 B.n123 585
R439 B.n220 B.n219 585
R440 B.n221 B.n122 585
R441 B.n223 B.n222 585
R442 B.n224 B.n121 585
R443 B.n226 B.n225 585
R444 B.n227 B.n120 585
R445 B.n228 B.n227 521.33
R446 B.n274 B.n273 521.33
R447 B.n442 B.n441 521.33
R448 B.n484 B.n29 521.33
R449 B.n114 B.t7 424.423
R450 B.n256 B.t10 424.423
R451 B.n42 B.t2 424.423
R452 B.n34 B.t5 424.423
R453 B.n115 B.t8 361.974
R454 B.n257 B.t11 361.974
R455 B.n43 B.t1 361.974
R456 B.n35 B.t4 361.974
R457 B.n569 B.n568 256.663
R458 B.n568 B.n567 235.042
R459 B.n568 B.n2 235.042
R460 B.n114 B.t6 209.236
R461 B.n256 B.t9 209.236
R462 B.n42 B.t0 209.236
R463 B.n34 B.t3 209.236
R464 B.n228 B.n119 163.367
R465 B.n232 B.n119 163.367
R466 B.n233 B.n232 163.367
R467 B.n234 B.n233 163.367
R468 B.n234 B.n117 163.367
R469 B.n238 B.n117 163.367
R470 B.n239 B.n238 163.367
R471 B.n240 B.n239 163.367
R472 B.n240 B.n113 163.367
R473 B.n245 B.n113 163.367
R474 B.n246 B.n245 163.367
R475 B.n247 B.n246 163.367
R476 B.n247 B.n111 163.367
R477 B.n251 B.n111 163.367
R478 B.n252 B.n251 163.367
R479 B.n253 B.n252 163.367
R480 B.n253 B.n109 163.367
R481 B.n260 B.n109 163.367
R482 B.n261 B.n260 163.367
R483 B.n262 B.n261 163.367
R484 B.n262 B.n107 163.367
R485 B.n266 B.n107 163.367
R486 B.n267 B.n266 163.367
R487 B.n268 B.n267 163.367
R488 B.n268 B.n105 163.367
R489 B.n272 B.n105 163.367
R490 B.n273 B.n272 163.367
R491 B.n441 B.n440 163.367
R492 B.n440 B.n49 163.367
R493 B.n436 B.n49 163.367
R494 B.n436 B.n435 163.367
R495 B.n435 B.n434 163.367
R496 B.n434 B.n51 163.367
R497 B.n430 B.n51 163.367
R498 B.n430 B.n429 163.367
R499 B.n429 B.n428 163.367
R500 B.n428 B.n53 163.367
R501 B.n424 B.n53 163.367
R502 B.n424 B.n423 163.367
R503 B.n423 B.n422 163.367
R504 B.n422 B.n55 163.367
R505 B.n418 B.n55 163.367
R506 B.n418 B.n417 163.367
R507 B.n417 B.n416 163.367
R508 B.n416 B.n57 163.367
R509 B.n412 B.n57 163.367
R510 B.n412 B.n411 163.367
R511 B.n411 B.n410 163.367
R512 B.n410 B.n59 163.367
R513 B.n406 B.n59 163.367
R514 B.n406 B.n405 163.367
R515 B.n405 B.n404 163.367
R516 B.n404 B.n61 163.367
R517 B.n400 B.n61 163.367
R518 B.n400 B.n399 163.367
R519 B.n399 B.n398 163.367
R520 B.n398 B.n63 163.367
R521 B.n394 B.n63 163.367
R522 B.n394 B.n393 163.367
R523 B.n393 B.n392 163.367
R524 B.n392 B.n65 163.367
R525 B.n388 B.n65 163.367
R526 B.n388 B.n387 163.367
R527 B.n387 B.n386 163.367
R528 B.n386 B.n67 163.367
R529 B.n382 B.n67 163.367
R530 B.n382 B.n381 163.367
R531 B.n381 B.n380 163.367
R532 B.n380 B.n69 163.367
R533 B.n376 B.n69 163.367
R534 B.n376 B.n375 163.367
R535 B.n375 B.n374 163.367
R536 B.n374 B.n71 163.367
R537 B.n370 B.n71 163.367
R538 B.n370 B.n369 163.367
R539 B.n369 B.n368 163.367
R540 B.n368 B.n73 163.367
R541 B.n364 B.n73 163.367
R542 B.n364 B.n363 163.367
R543 B.n363 B.n362 163.367
R544 B.n362 B.n75 163.367
R545 B.n358 B.n75 163.367
R546 B.n358 B.n357 163.367
R547 B.n357 B.n356 163.367
R548 B.n356 B.n77 163.367
R549 B.n352 B.n77 163.367
R550 B.n352 B.n351 163.367
R551 B.n351 B.n350 163.367
R552 B.n350 B.n79 163.367
R553 B.n346 B.n79 163.367
R554 B.n346 B.n345 163.367
R555 B.n345 B.n344 163.367
R556 B.n344 B.n81 163.367
R557 B.n340 B.n81 163.367
R558 B.n340 B.n339 163.367
R559 B.n339 B.n338 163.367
R560 B.n338 B.n83 163.367
R561 B.n334 B.n83 163.367
R562 B.n334 B.n333 163.367
R563 B.n333 B.n332 163.367
R564 B.n332 B.n85 163.367
R565 B.n328 B.n85 163.367
R566 B.n328 B.n327 163.367
R567 B.n327 B.n326 163.367
R568 B.n326 B.n87 163.367
R569 B.n322 B.n87 163.367
R570 B.n322 B.n321 163.367
R571 B.n321 B.n320 163.367
R572 B.n320 B.n89 163.367
R573 B.n316 B.n89 163.367
R574 B.n316 B.n315 163.367
R575 B.n315 B.n314 163.367
R576 B.n314 B.n91 163.367
R577 B.n310 B.n91 163.367
R578 B.n310 B.n309 163.367
R579 B.n309 B.n308 163.367
R580 B.n308 B.n93 163.367
R581 B.n304 B.n93 163.367
R582 B.n304 B.n303 163.367
R583 B.n303 B.n302 163.367
R584 B.n302 B.n95 163.367
R585 B.n298 B.n95 163.367
R586 B.n298 B.n297 163.367
R587 B.n297 B.n296 163.367
R588 B.n296 B.n97 163.367
R589 B.n292 B.n97 163.367
R590 B.n292 B.n291 163.367
R591 B.n291 B.n290 163.367
R592 B.n290 B.n99 163.367
R593 B.n286 B.n99 163.367
R594 B.n286 B.n285 163.367
R595 B.n285 B.n284 163.367
R596 B.n284 B.n101 163.367
R597 B.n280 B.n101 163.367
R598 B.n280 B.n279 163.367
R599 B.n279 B.n278 163.367
R600 B.n278 B.n103 163.367
R601 B.n274 B.n103 163.367
R602 B.n484 B.n483 163.367
R603 B.n483 B.n482 163.367
R604 B.n482 B.n31 163.367
R605 B.n478 B.n31 163.367
R606 B.n478 B.n477 163.367
R607 B.n477 B.n476 163.367
R608 B.n476 B.n33 163.367
R609 B.n472 B.n33 163.367
R610 B.n472 B.n471 163.367
R611 B.n471 B.n37 163.367
R612 B.n467 B.n37 163.367
R613 B.n467 B.n466 163.367
R614 B.n466 B.n465 163.367
R615 B.n465 B.n39 163.367
R616 B.n461 B.n39 163.367
R617 B.n461 B.n460 163.367
R618 B.n460 B.n459 163.367
R619 B.n459 B.n41 163.367
R620 B.n454 B.n41 163.367
R621 B.n454 B.n453 163.367
R622 B.n453 B.n452 163.367
R623 B.n452 B.n45 163.367
R624 B.n448 B.n45 163.367
R625 B.n448 B.n447 163.367
R626 B.n447 B.n446 163.367
R627 B.n446 B.n47 163.367
R628 B.n442 B.n47 163.367
R629 B.n488 B.n29 163.367
R630 B.n489 B.n488 163.367
R631 B.n490 B.n489 163.367
R632 B.n490 B.n27 163.367
R633 B.n494 B.n27 163.367
R634 B.n495 B.n494 163.367
R635 B.n496 B.n495 163.367
R636 B.n496 B.n25 163.367
R637 B.n500 B.n25 163.367
R638 B.n501 B.n500 163.367
R639 B.n502 B.n501 163.367
R640 B.n502 B.n23 163.367
R641 B.n506 B.n23 163.367
R642 B.n507 B.n506 163.367
R643 B.n508 B.n507 163.367
R644 B.n508 B.n21 163.367
R645 B.n512 B.n21 163.367
R646 B.n513 B.n512 163.367
R647 B.n514 B.n513 163.367
R648 B.n514 B.n19 163.367
R649 B.n518 B.n19 163.367
R650 B.n519 B.n518 163.367
R651 B.n520 B.n519 163.367
R652 B.n520 B.n17 163.367
R653 B.n524 B.n17 163.367
R654 B.n525 B.n524 163.367
R655 B.n526 B.n525 163.367
R656 B.n526 B.n15 163.367
R657 B.n530 B.n15 163.367
R658 B.n531 B.n530 163.367
R659 B.n532 B.n531 163.367
R660 B.n532 B.n13 163.367
R661 B.n536 B.n13 163.367
R662 B.n537 B.n536 163.367
R663 B.n538 B.n537 163.367
R664 B.n538 B.n11 163.367
R665 B.n542 B.n11 163.367
R666 B.n543 B.n542 163.367
R667 B.n544 B.n543 163.367
R668 B.n544 B.n9 163.367
R669 B.n548 B.n9 163.367
R670 B.n549 B.n548 163.367
R671 B.n550 B.n549 163.367
R672 B.n550 B.n7 163.367
R673 B.n554 B.n7 163.367
R674 B.n555 B.n554 163.367
R675 B.n556 B.n555 163.367
R676 B.n556 B.n5 163.367
R677 B.n560 B.n5 163.367
R678 B.n561 B.n560 163.367
R679 B.n562 B.n561 163.367
R680 B.n562 B.n3 163.367
R681 B.n566 B.n3 163.367
R682 B.n567 B.n566 163.367
R683 B.n148 B.n2 163.367
R684 B.n149 B.n148 163.367
R685 B.n150 B.n149 163.367
R686 B.n150 B.n145 163.367
R687 B.n154 B.n145 163.367
R688 B.n155 B.n154 163.367
R689 B.n156 B.n155 163.367
R690 B.n156 B.n143 163.367
R691 B.n160 B.n143 163.367
R692 B.n161 B.n160 163.367
R693 B.n162 B.n161 163.367
R694 B.n162 B.n141 163.367
R695 B.n166 B.n141 163.367
R696 B.n167 B.n166 163.367
R697 B.n168 B.n167 163.367
R698 B.n168 B.n139 163.367
R699 B.n172 B.n139 163.367
R700 B.n173 B.n172 163.367
R701 B.n174 B.n173 163.367
R702 B.n174 B.n137 163.367
R703 B.n178 B.n137 163.367
R704 B.n179 B.n178 163.367
R705 B.n180 B.n179 163.367
R706 B.n180 B.n135 163.367
R707 B.n184 B.n135 163.367
R708 B.n185 B.n184 163.367
R709 B.n186 B.n185 163.367
R710 B.n186 B.n133 163.367
R711 B.n190 B.n133 163.367
R712 B.n191 B.n190 163.367
R713 B.n192 B.n191 163.367
R714 B.n192 B.n131 163.367
R715 B.n196 B.n131 163.367
R716 B.n197 B.n196 163.367
R717 B.n198 B.n197 163.367
R718 B.n198 B.n129 163.367
R719 B.n202 B.n129 163.367
R720 B.n203 B.n202 163.367
R721 B.n204 B.n203 163.367
R722 B.n204 B.n127 163.367
R723 B.n208 B.n127 163.367
R724 B.n209 B.n208 163.367
R725 B.n210 B.n209 163.367
R726 B.n210 B.n125 163.367
R727 B.n214 B.n125 163.367
R728 B.n215 B.n214 163.367
R729 B.n216 B.n215 163.367
R730 B.n216 B.n123 163.367
R731 B.n220 B.n123 163.367
R732 B.n221 B.n220 163.367
R733 B.n222 B.n221 163.367
R734 B.n222 B.n121 163.367
R735 B.n226 B.n121 163.367
R736 B.n227 B.n226 163.367
R737 B.n115 B.n114 62.449
R738 B.n257 B.n256 62.449
R739 B.n43 B.n42 62.449
R740 B.n35 B.n34 62.449
R741 B.n242 B.n115 59.5399
R742 B.n258 B.n257 59.5399
R743 B.n456 B.n43 59.5399
R744 B.n36 B.n35 59.5399
R745 B.n486 B.n485 33.8737
R746 B.n443 B.n48 33.8737
R747 B.n275 B.n104 33.8737
R748 B.n229 B.n120 33.8737
R749 B B.n569 18.0485
R750 B.n487 B.n486 10.6151
R751 B.n487 B.n28 10.6151
R752 B.n491 B.n28 10.6151
R753 B.n492 B.n491 10.6151
R754 B.n493 B.n492 10.6151
R755 B.n493 B.n26 10.6151
R756 B.n497 B.n26 10.6151
R757 B.n498 B.n497 10.6151
R758 B.n499 B.n498 10.6151
R759 B.n499 B.n24 10.6151
R760 B.n503 B.n24 10.6151
R761 B.n504 B.n503 10.6151
R762 B.n505 B.n504 10.6151
R763 B.n505 B.n22 10.6151
R764 B.n509 B.n22 10.6151
R765 B.n510 B.n509 10.6151
R766 B.n511 B.n510 10.6151
R767 B.n511 B.n20 10.6151
R768 B.n515 B.n20 10.6151
R769 B.n516 B.n515 10.6151
R770 B.n517 B.n516 10.6151
R771 B.n517 B.n18 10.6151
R772 B.n521 B.n18 10.6151
R773 B.n522 B.n521 10.6151
R774 B.n523 B.n522 10.6151
R775 B.n523 B.n16 10.6151
R776 B.n527 B.n16 10.6151
R777 B.n528 B.n527 10.6151
R778 B.n529 B.n528 10.6151
R779 B.n529 B.n14 10.6151
R780 B.n533 B.n14 10.6151
R781 B.n534 B.n533 10.6151
R782 B.n535 B.n534 10.6151
R783 B.n535 B.n12 10.6151
R784 B.n539 B.n12 10.6151
R785 B.n540 B.n539 10.6151
R786 B.n541 B.n540 10.6151
R787 B.n541 B.n10 10.6151
R788 B.n545 B.n10 10.6151
R789 B.n546 B.n545 10.6151
R790 B.n547 B.n546 10.6151
R791 B.n547 B.n8 10.6151
R792 B.n551 B.n8 10.6151
R793 B.n552 B.n551 10.6151
R794 B.n553 B.n552 10.6151
R795 B.n553 B.n6 10.6151
R796 B.n557 B.n6 10.6151
R797 B.n558 B.n557 10.6151
R798 B.n559 B.n558 10.6151
R799 B.n559 B.n4 10.6151
R800 B.n563 B.n4 10.6151
R801 B.n564 B.n563 10.6151
R802 B.n565 B.n564 10.6151
R803 B.n565 B.n0 10.6151
R804 B.n485 B.n30 10.6151
R805 B.n481 B.n30 10.6151
R806 B.n481 B.n480 10.6151
R807 B.n480 B.n479 10.6151
R808 B.n479 B.n32 10.6151
R809 B.n475 B.n32 10.6151
R810 B.n475 B.n474 10.6151
R811 B.n474 B.n473 10.6151
R812 B.n470 B.n469 10.6151
R813 B.n469 B.n468 10.6151
R814 B.n468 B.n38 10.6151
R815 B.n464 B.n38 10.6151
R816 B.n464 B.n463 10.6151
R817 B.n463 B.n462 10.6151
R818 B.n462 B.n40 10.6151
R819 B.n458 B.n40 10.6151
R820 B.n458 B.n457 10.6151
R821 B.n455 B.n44 10.6151
R822 B.n451 B.n44 10.6151
R823 B.n451 B.n450 10.6151
R824 B.n450 B.n449 10.6151
R825 B.n449 B.n46 10.6151
R826 B.n445 B.n46 10.6151
R827 B.n445 B.n444 10.6151
R828 B.n444 B.n443 10.6151
R829 B.n439 B.n48 10.6151
R830 B.n439 B.n438 10.6151
R831 B.n438 B.n437 10.6151
R832 B.n437 B.n50 10.6151
R833 B.n433 B.n50 10.6151
R834 B.n433 B.n432 10.6151
R835 B.n432 B.n431 10.6151
R836 B.n431 B.n52 10.6151
R837 B.n427 B.n52 10.6151
R838 B.n427 B.n426 10.6151
R839 B.n426 B.n425 10.6151
R840 B.n425 B.n54 10.6151
R841 B.n421 B.n54 10.6151
R842 B.n421 B.n420 10.6151
R843 B.n420 B.n419 10.6151
R844 B.n419 B.n56 10.6151
R845 B.n415 B.n56 10.6151
R846 B.n415 B.n414 10.6151
R847 B.n414 B.n413 10.6151
R848 B.n413 B.n58 10.6151
R849 B.n409 B.n58 10.6151
R850 B.n409 B.n408 10.6151
R851 B.n408 B.n407 10.6151
R852 B.n407 B.n60 10.6151
R853 B.n403 B.n60 10.6151
R854 B.n403 B.n402 10.6151
R855 B.n402 B.n401 10.6151
R856 B.n401 B.n62 10.6151
R857 B.n397 B.n62 10.6151
R858 B.n397 B.n396 10.6151
R859 B.n396 B.n395 10.6151
R860 B.n395 B.n64 10.6151
R861 B.n391 B.n64 10.6151
R862 B.n391 B.n390 10.6151
R863 B.n390 B.n389 10.6151
R864 B.n389 B.n66 10.6151
R865 B.n385 B.n66 10.6151
R866 B.n385 B.n384 10.6151
R867 B.n384 B.n383 10.6151
R868 B.n383 B.n68 10.6151
R869 B.n379 B.n68 10.6151
R870 B.n379 B.n378 10.6151
R871 B.n378 B.n377 10.6151
R872 B.n377 B.n70 10.6151
R873 B.n373 B.n70 10.6151
R874 B.n373 B.n372 10.6151
R875 B.n372 B.n371 10.6151
R876 B.n371 B.n72 10.6151
R877 B.n367 B.n72 10.6151
R878 B.n367 B.n366 10.6151
R879 B.n366 B.n365 10.6151
R880 B.n365 B.n74 10.6151
R881 B.n361 B.n74 10.6151
R882 B.n361 B.n360 10.6151
R883 B.n360 B.n359 10.6151
R884 B.n359 B.n76 10.6151
R885 B.n355 B.n76 10.6151
R886 B.n355 B.n354 10.6151
R887 B.n354 B.n353 10.6151
R888 B.n353 B.n78 10.6151
R889 B.n349 B.n78 10.6151
R890 B.n349 B.n348 10.6151
R891 B.n348 B.n347 10.6151
R892 B.n347 B.n80 10.6151
R893 B.n343 B.n80 10.6151
R894 B.n343 B.n342 10.6151
R895 B.n342 B.n341 10.6151
R896 B.n341 B.n82 10.6151
R897 B.n337 B.n82 10.6151
R898 B.n337 B.n336 10.6151
R899 B.n336 B.n335 10.6151
R900 B.n335 B.n84 10.6151
R901 B.n331 B.n84 10.6151
R902 B.n331 B.n330 10.6151
R903 B.n330 B.n329 10.6151
R904 B.n329 B.n86 10.6151
R905 B.n325 B.n86 10.6151
R906 B.n325 B.n324 10.6151
R907 B.n324 B.n323 10.6151
R908 B.n323 B.n88 10.6151
R909 B.n319 B.n88 10.6151
R910 B.n319 B.n318 10.6151
R911 B.n318 B.n317 10.6151
R912 B.n317 B.n90 10.6151
R913 B.n313 B.n90 10.6151
R914 B.n313 B.n312 10.6151
R915 B.n312 B.n311 10.6151
R916 B.n311 B.n92 10.6151
R917 B.n307 B.n92 10.6151
R918 B.n307 B.n306 10.6151
R919 B.n306 B.n305 10.6151
R920 B.n305 B.n94 10.6151
R921 B.n301 B.n94 10.6151
R922 B.n301 B.n300 10.6151
R923 B.n300 B.n299 10.6151
R924 B.n299 B.n96 10.6151
R925 B.n295 B.n96 10.6151
R926 B.n295 B.n294 10.6151
R927 B.n294 B.n293 10.6151
R928 B.n293 B.n98 10.6151
R929 B.n289 B.n98 10.6151
R930 B.n289 B.n288 10.6151
R931 B.n288 B.n287 10.6151
R932 B.n287 B.n100 10.6151
R933 B.n283 B.n100 10.6151
R934 B.n283 B.n282 10.6151
R935 B.n282 B.n281 10.6151
R936 B.n281 B.n102 10.6151
R937 B.n277 B.n102 10.6151
R938 B.n277 B.n276 10.6151
R939 B.n276 B.n275 10.6151
R940 B.n147 B.n1 10.6151
R941 B.n147 B.n146 10.6151
R942 B.n151 B.n146 10.6151
R943 B.n152 B.n151 10.6151
R944 B.n153 B.n152 10.6151
R945 B.n153 B.n144 10.6151
R946 B.n157 B.n144 10.6151
R947 B.n158 B.n157 10.6151
R948 B.n159 B.n158 10.6151
R949 B.n159 B.n142 10.6151
R950 B.n163 B.n142 10.6151
R951 B.n164 B.n163 10.6151
R952 B.n165 B.n164 10.6151
R953 B.n165 B.n140 10.6151
R954 B.n169 B.n140 10.6151
R955 B.n170 B.n169 10.6151
R956 B.n171 B.n170 10.6151
R957 B.n171 B.n138 10.6151
R958 B.n175 B.n138 10.6151
R959 B.n176 B.n175 10.6151
R960 B.n177 B.n176 10.6151
R961 B.n177 B.n136 10.6151
R962 B.n181 B.n136 10.6151
R963 B.n182 B.n181 10.6151
R964 B.n183 B.n182 10.6151
R965 B.n183 B.n134 10.6151
R966 B.n187 B.n134 10.6151
R967 B.n188 B.n187 10.6151
R968 B.n189 B.n188 10.6151
R969 B.n189 B.n132 10.6151
R970 B.n193 B.n132 10.6151
R971 B.n194 B.n193 10.6151
R972 B.n195 B.n194 10.6151
R973 B.n195 B.n130 10.6151
R974 B.n199 B.n130 10.6151
R975 B.n200 B.n199 10.6151
R976 B.n201 B.n200 10.6151
R977 B.n201 B.n128 10.6151
R978 B.n205 B.n128 10.6151
R979 B.n206 B.n205 10.6151
R980 B.n207 B.n206 10.6151
R981 B.n207 B.n126 10.6151
R982 B.n211 B.n126 10.6151
R983 B.n212 B.n211 10.6151
R984 B.n213 B.n212 10.6151
R985 B.n213 B.n124 10.6151
R986 B.n217 B.n124 10.6151
R987 B.n218 B.n217 10.6151
R988 B.n219 B.n218 10.6151
R989 B.n219 B.n122 10.6151
R990 B.n223 B.n122 10.6151
R991 B.n224 B.n223 10.6151
R992 B.n225 B.n224 10.6151
R993 B.n225 B.n120 10.6151
R994 B.n230 B.n229 10.6151
R995 B.n231 B.n230 10.6151
R996 B.n231 B.n118 10.6151
R997 B.n235 B.n118 10.6151
R998 B.n236 B.n235 10.6151
R999 B.n237 B.n236 10.6151
R1000 B.n237 B.n116 10.6151
R1001 B.n241 B.n116 10.6151
R1002 B.n244 B.n243 10.6151
R1003 B.n244 B.n112 10.6151
R1004 B.n248 B.n112 10.6151
R1005 B.n249 B.n248 10.6151
R1006 B.n250 B.n249 10.6151
R1007 B.n250 B.n110 10.6151
R1008 B.n254 B.n110 10.6151
R1009 B.n255 B.n254 10.6151
R1010 B.n259 B.n255 10.6151
R1011 B.n263 B.n108 10.6151
R1012 B.n264 B.n263 10.6151
R1013 B.n265 B.n264 10.6151
R1014 B.n265 B.n106 10.6151
R1015 B.n269 B.n106 10.6151
R1016 B.n270 B.n269 10.6151
R1017 B.n271 B.n270 10.6151
R1018 B.n271 B.n104 10.6151
R1019 B.n473 B.n36 9.36635
R1020 B.n456 B.n455 9.36635
R1021 B.n242 B.n241 9.36635
R1022 B.n258 B.n108 9.36635
R1023 B.n569 B.n0 8.11757
R1024 B.n569 B.n1 8.11757
R1025 B.n470 B.n36 1.24928
R1026 B.n457 B.n456 1.24928
R1027 B.n243 B.n242 1.24928
R1028 B.n259 B.n258 1.24928
R1029 VN.n59 VN.n31 161.3
R1030 VN.n58 VN.n57 161.3
R1031 VN.n56 VN.n32 161.3
R1032 VN.n55 VN.n54 161.3
R1033 VN.n53 VN.n33 161.3
R1034 VN.n52 VN.n51 161.3
R1035 VN.n50 VN.n34 161.3
R1036 VN.n49 VN.n48 161.3
R1037 VN.n47 VN.n35 161.3
R1038 VN.n46 VN.n45 161.3
R1039 VN.n44 VN.n37 161.3
R1040 VN.n43 VN.n42 161.3
R1041 VN.n41 VN.n38 161.3
R1042 VN.n28 VN.n0 161.3
R1043 VN.n27 VN.n26 161.3
R1044 VN.n25 VN.n1 161.3
R1045 VN.n24 VN.n23 161.3
R1046 VN.n22 VN.n2 161.3
R1047 VN.n21 VN.n20 161.3
R1048 VN.n19 VN.n3 161.3
R1049 VN.n18 VN.n17 161.3
R1050 VN.n15 VN.n4 161.3
R1051 VN.n14 VN.n13 161.3
R1052 VN.n12 VN.n5 161.3
R1053 VN.n11 VN.n10 161.3
R1054 VN.n9 VN.n6 161.3
R1055 VN.n30 VN.n29 106.974
R1056 VN.n61 VN.n60 106.974
R1057 VN.n14 VN.n5 56.5617
R1058 VN.n46 VN.n37 56.5617
R1059 VN.n8 VN.n7 56.2048
R1060 VN.n40 VN.n39 56.2048
R1061 VN VN.n61 44.2255
R1062 VN.n23 VN.n22 43.4833
R1063 VN.n54 VN.n53 43.4833
R1064 VN.n7 VN.t6 42.2769
R1065 VN.n39 VN.t4 42.2769
R1066 VN.n23 VN.n1 37.6707
R1067 VN.n54 VN.n32 37.6707
R1068 VN.n10 VN.n9 24.5923
R1069 VN.n10 VN.n5 24.5923
R1070 VN.n15 VN.n14 24.5923
R1071 VN.n17 VN.n15 24.5923
R1072 VN.n21 VN.n3 24.5923
R1073 VN.n22 VN.n21 24.5923
R1074 VN.n27 VN.n1 24.5923
R1075 VN.n28 VN.n27 24.5923
R1076 VN.n42 VN.n37 24.5923
R1077 VN.n42 VN.n41 24.5923
R1078 VN.n53 VN.n52 24.5923
R1079 VN.n52 VN.n34 24.5923
R1080 VN.n48 VN.n47 24.5923
R1081 VN.n47 VN.n46 24.5923
R1082 VN.n59 VN.n58 24.5923
R1083 VN.n58 VN.n32 24.5923
R1084 VN.n9 VN.n8 17.7066
R1085 VN.n17 VN.n16 17.7066
R1086 VN.n41 VN.n40 17.7066
R1087 VN.n48 VN.n36 17.7066
R1088 VN.n8 VN.t2 8.67316
R1089 VN.n16 VN.t7 8.67316
R1090 VN.n29 VN.t1 8.67316
R1091 VN.n40 VN.t3 8.67316
R1092 VN.n36 VN.t5 8.67316
R1093 VN.n60 VN.t0 8.67316
R1094 VN.n16 VN.n3 6.88621
R1095 VN.n36 VN.n34 6.88621
R1096 VN.n39 VN.n38 5.01074
R1097 VN.n7 VN.n6 5.01074
R1098 VN.n29 VN.n28 3.93519
R1099 VN.n60 VN.n59 3.93519
R1100 VN.n61 VN.n31 0.278335
R1101 VN.n30 VN.n0 0.278335
R1102 VN.n57 VN.n31 0.189894
R1103 VN.n57 VN.n56 0.189894
R1104 VN.n56 VN.n55 0.189894
R1105 VN.n55 VN.n33 0.189894
R1106 VN.n51 VN.n33 0.189894
R1107 VN.n51 VN.n50 0.189894
R1108 VN.n50 VN.n49 0.189894
R1109 VN.n49 VN.n35 0.189894
R1110 VN.n45 VN.n35 0.189894
R1111 VN.n45 VN.n44 0.189894
R1112 VN.n44 VN.n43 0.189894
R1113 VN.n43 VN.n38 0.189894
R1114 VN.n11 VN.n6 0.189894
R1115 VN.n12 VN.n11 0.189894
R1116 VN.n13 VN.n12 0.189894
R1117 VN.n13 VN.n4 0.189894
R1118 VN.n18 VN.n4 0.189894
R1119 VN.n19 VN.n18 0.189894
R1120 VN.n20 VN.n19 0.189894
R1121 VN.n20 VN.n2 0.189894
R1122 VN.n24 VN.n2 0.189894
R1123 VN.n25 VN.n24 0.189894
R1124 VN.n26 VN.n25 0.189894
R1125 VN.n26 VN.n0 0.189894
R1126 VN VN.n30 0.153485
R1127 VDD2.n2 VDD2.n1 346.433
R1128 VDD2.n2 VDD2.n0 346.433
R1129 VDD2 VDD2.n5 346.43
R1130 VDD2.n4 VDD2.n3 345.099
R1131 VDD2.n4 VDD2.n2 37.1032
R1132 VDD2.n5 VDD2.t4 31.2553
R1133 VDD2.n5 VDD2.t3 31.2553
R1134 VDD2.n3 VDD2.t7 31.2553
R1135 VDD2.n3 VDD2.t2 31.2553
R1136 VDD2.n1 VDD2.t0 31.2553
R1137 VDD2.n1 VDD2.t6 31.2553
R1138 VDD2.n0 VDD2.t1 31.2553
R1139 VDD2.n0 VDD2.t5 31.2553
R1140 VDD2 VDD2.n4 1.44662
C0 VDD1 w_n4190_n1176# 1.74018f
C1 VTAIL VDD1 4.66689f
C2 VN w_n4190_n1176# 8.42027f
C3 VN VTAIL 2.60157f
C4 VDD2 VDD1 1.92583f
C5 VN VDD2 1.20506f
C6 B VP 2.04608f
C7 VTAIL w_n4190_n1176# 1.72011f
C8 VDD2 w_n4190_n1176# 1.86599f
C9 VDD2 VTAIL 4.72325f
C10 B VDD1 1.44137f
C11 B VN 1.13248f
C12 VP VDD1 1.6013f
C13 VN VP 5.98871f
C14 B w_n4190_n1176# 7.58188f
C15 B VTAIL 1.2826f
C16 VN VDD1 0.159268f
C17 B VDD2 1.54718f
C18 VP w_n4190_n1176# 8.957459f
C19 VP VTAIL 2.61568f
C20 VP VDD2 0.559482f
C21 VDD2 VSUBS 1.180874f
C22 VDD1 VSUBS 1.861283f
C23 VTAIL VSUBS 0.568003f
C24 VN VSUBS 7.44256f
C25 VP VSUBS 3.22262f
C26 B VSUBS 4.135168f
C27 w_n4190_n1176# VSUBS 63.503597f
C28 VDD2.t1 VSUBS 0.015715f
C29 VDD2.t5 VSUBS 0.015715f
C30 VDD2.n0 VSUBS 0.05362f
C31 VDD2.t0 VSUBS 0.015715f
C32 VDD2.t6 VSUBS 0.015715f
C33 VDD2.n1 VSUBS 0.05362f
C34 VDD2.n2 VSUBS 2.11625f
C35 VDD2.t7 VSUBS 0.015715f
C36 VDD2.t2 VSUBS 0.015715f
C37 VDD2.n3 VSUBS 0.052054f
C38 VDD2.n4 VSUBS 1.66887f
C39 VDD2.t4 VSUBS 0.015715f
C40 VDD2.t3 VSUBS 0.015715f
C41 VDD2.n5 VSUBS 0.053615f
C42 VN.n0 VSUBS 0.076321f
C43 VN.t1 VSUBS 0.331342f
C44 VN.n1 VSUBS 0.115821f
C45 VN.n2 VSUBS 0.057893f
C46 VN.n3 VSUBS 0.069197f
C47 VN.n4 VSUBS 0.057893f
C48 VN.n5 VSUBS 0.084156f
C49 VN.n6 VSUBS 0.61319f
C50 VN.t2 VSUBS 0.331342f
C51 VN.t6 VSUBS 0.814595f
C52 VN.n7 VSUBS 0.413529f
C53 VN.n8 VSUBS 0.406623f
C54 VN.n9 VSUBS 0.092517f
C55 VN.n10 VSUBS 0.107357f
C56 VN.n11 VSUBS 0.057893f
C57 VN.n12 VSUBS 0.057893f
C58 VN.n13 VSUBS 0.057893f
C59 VN.n14 VSUBS 0.084156f
C60 VN.n15 VSUBS 0.107357f
C61 VN.t7 VSUBS 0.331342f
C62 VN.n16 VSUBS 0.215544f
C63 VN.n17 VSUBS 0.092517f
C64 VN.n18 VSUBS 0.057893f
C65 VN.n19 VSUBS 0.057893f
C66 VN.n20 VSUBS 0.057893f
C67 VN.n21 VSUBS 0.107357f
C68 VN.n22 VSUBS 0.112422f
C69 VN.n23 VSUBS 0.047426f
C70 VN.n24 VSUBS 0.057893f
C71 VN.n25 VSUBS 0.057893f
C72 VN.n26 VSUBS 0.057893f
C73 VN.n27 VSUBS 0.107357f
C74 VN.n28 VSUBS 0.062837f
C75 VN.n29 VSUBS 0.411311f
C76 VN.n30 VSUBS 0.108636f
C77 VN.n31 VSUBS 0.076321f
C78 VN.t0 VSUBS 0.331342f
C79 VN.n32 VSUBS 0.115821f
C80 VN.n33 VSUBS 0.057893f
C81 VN.n34 VSUBS 0.069197f
C82 VN.n35 VSUBS 0.057893f
C83 VN.t5 VSUBS 0.331342f
C84 VN.n36 VSUBS 0.215544f
C85 VN.n37 VSUBS 0.084156f
C86 VN.n38 VSUBS 0.61319f
C87 VN.t3 VSUBS 0.331342f
C88 VN.t4 VSUBS 0.814595f
C89 VN.n39 VSUBS 0.413529f
C90 VN.n40 VSUBS 0.406623f
C91 VN.n41 VSUBS 0.092517f
C92 VN.n42 VSUBS 0.107357f
C93 VN.n43 VSUBS 0.057893f
C94 VN.n44 VSUBS 0.057893f
C95 VN.n45 VSUBS 0.057893f
C96 VN.n46 VSUBS 0.084156f
C97 VN.n47 VSUBS 0.107357f
C98 VN.n48 VSUBS 0.092517f
C99 VN.n49 VSUBS 0.057893f
C100 VN.n50 VSUBS 0.057893f
C101 VN.n51 VSUBS 0.057893f
C102 VN.n52 VSUBS 0.107357f
C103 VN.n53 VSUBS 0.112422f
C104 VN.n54 VSUBS 0.047426f
C105 VN.n55 VSUBS 0.057893f
C106 VN.n56 VSUBS 0.057893f
C107 VN.n57 VSUBS 0.057893f
C108 VN.n58 VSUBS 0.107357f
C109 VN.n59 VSUBS 0.062837f
C110 VN.n60 VSUBS 0.411311f
C111 VN.n61 VSUBS 2.69491f
C112 B.n0 VSUBS 0.011032f
C113 B.n1 VSUBS 0.011032f
C114 B.n2 VSUBS 0.016316f
C115 B.n3 VSUBS 0.012503f
C116 B.n4 VSUBS 0.012503f
C117 B.n5 VSUBS 0.012503f
C118 B.n6 VSUBS 0.012503f
C119 B.n7 VSUBS 0.012503f
C120 B.n8 VSUBS 0.012503f
C121 B.n9 VSUBS 0.012503f
C122 B.n10 VSUBS 0.012503f
C123 B.n11 VSUBS 0.012503f
C124 B.n12 VSUBS 0.012503f
C125 B.n13 VSUBS 0.012503f
C126 B.n14 VSUBS 0.012503f
C127 B.n15 VSUBS 0.012503f
C128 B.n16 VSUBS 0.012503f
C129 B.n17 VSUBS 0.012503f
C130 B.n18 VSUBS 0.012503f
C131 B.n19 VSUBS 0.012503f
C132 B.n20 VSUBS 0.012503f
C133 B.n21 VSUBS 0.012503f
C134 B.n22 VSUBS 0.012503f
C135 B.n23 VSUBS 0.012503f
C136 B.n24 VSUBS 0.012503f
C137 B.n25 VSUBS 0.012503f
C138 B.n26 VSUBS 0.012503f
C139 B.n27 VSUBS 0.012503f
C140 B.n28 VSUBS 0.012503f
C141 B.n29 VSUBS 0.029536f
C142 B.n30 VSUBS 0.012503f
C143 B.n31 VSUBS 0.012503f
C144 B.n32 VSUBS 0.012503f
C145 B.n33 VSUBS 0.012503f
C146 B.t4 VSUBS 0.034931f
C147 B.t5 VSUBS 0.044986f
C148 B.t3 VSUBS 0.271458f
C149 B.n34 VSUBS 0.113827f
C150 B.n35 VSUBS 0.086174f
C151 B.n36 VSUBS 0.028968f
C152 B.n37 VSUBS 0.012503f
C153 B.n38 VSUBS 0.012503f
C154 B.n39 VSUBS 0.012503f
C155 B.n40 VSUBS 0.012503f
C156 B.n41 VSUBS 0.012503f
C157 B.t1 VSUBS 0.034931f
C158 B.t2 VSUBS 0.044986f
C159 B.t0 VSUBS 0.271458f
C160 B.n42 VSUBS 0.113827f
C161 B.n43 VSUBS 0.086174f
C162 B.n44 VSUBS 0.012503f
C163 B.n45 VSUBS 0.012503f
C164 B.n46 VSUBS 0.012503f
C165 B.n47 VSUBS 0.012503f
C166 B.n48 VSUBS 0.029536f
C167 B.n49 VSUBS 0.012503f
C168 B.n50 VSUBS 0.012503f
C169 B.n51 VSUBS 0.012503f
C170 B.n52 VSUBS 0.012503f
C171 B.n53 VSUBS 0.012503f
C172 B.n54 VSUBS 0.012503f
C173 B.n55 VSUBS 0.012503f
C174 B.n56 VSUBS 0.012503f
C175 B.n57 VSUBS 0.012503f
C176 B.n58 VSUBS 0.012503f
C177 B.n59 VSUBS 0.012503f
C178 B.n60 VSUBS 0.012503f
C179 B.n61 VSUBS 0.012503f
C180 B.n62 VSUBS 0.012503f
C181 B.n63 VSUBS 0.012503f
C182 B.n64 VSUBS 0.012503f
C183 B.n65 VSUBS 0.012503f
C184 B.n66 VSUBS 0.012503f
C185 B.n67 VSUBS 0.012503f
C186 B.n68 VSUBS 0.012503f
C187 B.n69 VSUBS 0.012503f
C188 B.n70 VSUBS 0.012503f
C189 B.n71 VSUBS 0.012503f
C190 B.n72 VSUBS 0.012503f
C191 B.n73 VSUBS 0.012503f
C192 B.n74 VSUBS 0.012503f
C193 B.n75 VSUBS 0.012503f
C194 B.n76 VSUBS 0.012503f
C195 B.n77 VSUBS 0.012503f
C196 B.n78 VSUBS 0.012503f
C197 B.n79 VSUBS 0.012503f
C198 B.n80 VSUBS 0.012503f
C199 B.n81 VSUBS 0.012503f
C200 B.n82 VSUBS 0.012503f
C201 B.n83 VSUBS 0.012503f
C202 B.n84 VSUBS 0.012503f
C203 B.n85 VSUBS 0.012503f
C204 B.n86 VSUBS 0.012503f
C205 B.n87 VSUBS 0.012503f
C206 B.n88 VSUBS 0.012503f
C207 B.n89 VSUBS 0.012503f
C208 B.n90 VSUBS 0.012503f
C209 B.n91 VSUBS 0.012503f
C210 B.n92 VSUBS 0.012503f
C211 B.n93 VSUBS 0.012503f
C212 B.n94 VSUBS 0.012503f
C213 B.n95 VSUBS 0.012503f
C214 B.n96 VSUBS 0.012503f
C215 B.n97 VSUBS 0.012503f
C216 B.n98 VSUBS 0.012503f
C217 B.n99 VSUBS 0.012503f
C218 B.n100 VSUBS 0.012503f
C219 B.n101 VSUBS 0.012503f
C220 B.n102 VSUBS 0.012503f
C221 B.n103 VSUBS 0.012503f
C222 B.n104 VSUBS 0.02898f
C223 B.n105 VSUBS 0.012503f
C224 B.n106 VSUBS 0.012503f
C225 B.n107 VSUBS 0.012503f
C226 B.n108 VSUBS 0.011768f
C227 B.n109 VSUBS 0.012503f
C228 B.n110 VSUBS 0.012503f
C229 B.n111 VSUBS 0.012503f
C230 B.n112 VSUBS 0.012503f
C231 B.n113 VSUBS 0.012503f
C232 B.t8 VSUBS 0.034931f
C233 B.t7 VSUBS 0.044986f
C234 B.t6 VSUBS 0.271458f
C235 B.n114 VSUBS 0.113827f
C236 B.n115 VSUBS 0.086174f
C237 B.n116 VSUBS 0.012503f
C238 B.n117 VSUBS 0.012503f
C239 B.n118 VSUBS 0.012503f
C240 B.n119 VSUBS 0.012503f
C241 B.n120 VSUBS 0.029536f
C242 B.n121 VSUBS 0.012503f
C243 B.n122 VSUBS 0.012503f
C244 B.n123 VSUBS 0.012503f
C245 B.n124 VSUBS 0.012503f
C246 B.n125 VSUBS 0.012503f
C247 B.n126 VSUBS 0.012503f
C248 B.n127 VSUBS 0.012503f
C249 B.n128 VSUBS 0.012503f
C250 B.n129 VSUBS 0.012503f
C251 B.n130 VSUBS 0.012503f
C252 B.n131 VSUBS 0.012503f
C253 B.n132 VSUBS 0.012503f
C254 B.n133 VSUBS 0.012503f
C255 B.n134 VSUBS 0.012503f
C256 B.n135 VSUBS 0.012503f
C257 B.n136 VSUBS 0.012503f
C258 B.n137 VSUBS 0.012503f
C259 B.n138 VSUBS 0.012503f
C260 B.n139 VSUBS 0.012503f
C261 B.n140 VSUBS 0.012503f
C262 B.n141 VSUBS 0.012503f
C263 B.n142 VSUBS 0.012503f
C264 B.n143 VSUBS 0.012503f
C265 B.n144 VSUBS 0.012503f
C266 B.n145 VSUBS 0.012503f
C267 B.n146 VSUBS 0.012503f
C268 B.n147 VSUBS 0.012503f
C269 B.n148 VSUBS 0.012503f
C270 B.n149 VSUBS 0.012503f
C271 B.n150 VSUBS 0.012503f
C272 B.n151 VSUBS 0.012503f
C273 B.n152 VSUBS 0.012503f
C274 B.n153 VSUBS 0.012503f
C275 B.n154 VSUBS 0.012503f
C276 B.n155 VSUBS 0.012503f
C277 B.n156 VSUBS 0.012503f
C278 B.n157 VSUBS 0.012503f
C279 B.n158 VSUBS 0.012503f
C280 B.n159 VSUBS 0.012503f
C281 B.n160 VSUBS 0.012503f
C282 B.n161 VSUBS 0.012503f
C283 B.n162 VSUBS 0.012503f
C284 B.n163 VSUBS 0.012503f
C285 B.n164 VSUBS 0.012503f
C286 B.n165 VSUBS 0.012503f
C287 B.n166 VSUBS 0.012503f
C288 B.n167 VSUBS 0.012503f
C289 B.n168 VSUBS 0.012503f
C290 B.n169 VSUBS 0.012503f
C291 B.n170 VSUBS 0.012503f
C292 B.n171 VSUBS 0.012503f
C293 B.n172 VSUBS 0.012503f
C294 B.n173 VSUBS 0.012503f
C295 B.n174 VSUBS 0.012503f
C296 B.n175 VSUBS 0.012503f
C297 B.n176 VSUBS 0.012503f
C298 B.n177 VSUBS 0.012503f
C299 B.n178 VSUBS 0.012503f
C300 B.n179 VSUBS 0.012503f
C301 B.n180 VSUBS 0.012503f
C302 B.n181 VSUBS 0.012503f
C303 B.n182 VSUBS 0.012503f
C304 B.n183 VSUBS 0.012503f
C305 B.n184 VSUBS 0.012503f
C306 B.n185 VSUBS 0.012503f
C307 B.n186 VSUBS 0.012503f
C308 B.n187 VSUBS 0.012503f
C309 B.n188 VSUBS 0.012503f
C310 B.n189 VSUBS 0.012503f
C311 B.n190 VSUBS 0.012503f
C312 B.n191 VSUBS 0.012503f
C313 B.n192 VSUBS 0.012503f
C314 B.n193 VSUBS 0.012503f
C315 B.n194 VSUBS 0.012503f
C316 B.n195 VSUBS 0.012503f
C317 B.n196 VSUBS 0.012503f
C318 B.n197 VSUBS 0.012503f
C319 B.n198 VSUBS 0.012503f
C320 B.n199 VSUBS 0.012503f
C321 B.n200 VSUBS 0.012503f
C322 B.n201 VSUBS 0.012503f
C323 B.n202 VSUBS 0.012503f
C324 B.n203 VSUBS 0.012503f
C325 B.n204 VSUBS 0.012503f
C326 B.n205 VSUBS 0.012503f
C327 B.n206 VSUBS 0.012503f
C328 B.n207 VSUBS 0.012503f
C329 B.n208 VSUBS 0.012503f
C330 B.n209 VSUBS 0.012503f
C331 B.n210 VSUBS 0.012503f
C332 B.n211 VSUBS 0.012503f
C333 B.n212 VSUBS 0.012503f
C334 B.n213 VSUBS 0.012503f
C335 B.n214 VSUBS 0.012503f
C336 B.n215 VSUBS 0.012503f
C337 B.n216 VSUBS 0.012503f
C338 B.n217 VSUBS 0.012503f
C339 B.n218 VSUBS 0.012503f
C340 B.n219 VSUBS 0.012503f
C341 B.n220 VSUBS 0.012503f
C342 B.n221 VSUBS 0.012503f
C343 B.n222 VSUBS 0.012503f
C344 B.n223 VSUBS 0.012503f
C345 B.n224 VSUBS 0.012503f
C346 B.n225 VSUBS 0.012503f
C347 B.n226 VSUBS 0.012503f
C348 B.n227 VSUBS 0.029536f
C349 B.n228 VSUBS 0.030405f
C350 B.n229 VSUBS 0.030405f
C351 B.n230 VSUBS 0.012503f
C352 B.n231 VSUBS 0.012503f
C353 B.n232 VSUBS 0.012503f
C354 B.n233 VSUBS 0.012503f
C355 B.n234 VSUBS 0.012503f
C356 B.n235 VSUBS 0.012503f
C357 B.n236 VSUBS 0.012503f
C358 B.n237 VSUBS 0.012503f
C359 B.n238 VSUBS 0.012503f
C360 B.n239 VSUBS 0.012503f
C361 B.n240 VSUBS 0.012503f
C362 B.n241 VSUBS 0.011768f
C363 B.n242 VSUBS 0.028968f
C364 B.n243 VSUBS 0.006987f
C365 B.n244 VSUBS 0.012503f
C366 B.n245 VSUBS 0.012503f
C367 B.n246 VSUBS 0.012503f
C368 B.n247 VSUBS 0.012503f
C369 B.n248 VSUBS 0.012503f
C370 B.n249 VSUBS 0.012503f
C371 B.n250 VSUBS 0.012503f
C372 B.n251 VSUBS 0.012503f
C373 B.n252 VSUBS 0.012503f
C374 B.n253 VSUBS 0.012503f
C375 B.n254 VSUBS 0.012503f
C376 B.n255 VSUBS 0.012503f
C377 B.t11 VSUBS 0.034931f
C378 B.t10 VSUBS 0.044986f
C379 B.t9 VSUBS 0.271458f
C380 B.n256 VSUBS 0.113827f
C381 B.n257 VSUBS 0.086174f
C382 B.n258 VSUBS 0.028968f
C383 B.n259 VSUBS 0.006987f
C384 B.n260 VSUBS 0.012503f
C385 B.n261 VSUBS 0.012503f
C386 B.n262 VSUBS 0.012503f
C387 B.n263 VSUBS 0.012503f
C388 B.n264 VSUBS 0.012503f
C389 B.n265 VSUBS 0.012503f
C390 B.n266 VSUBS 0.012503f
C391 B.n267 VSUBS 0.012503f
C392 B.n268 VSUBS 0.012503f
C393 B.n269 VSUBS 0.012503f
C394 B.n270 VSUBS 0.012503f
C395 B.n271 VSUBS 0.012503f
C396 B.n272 VSUBS 0.012503f
C397 B.n273 VSUBS 0.030405f
C398 B.n274 VSUBS 0.029536f
C399 B.n275 VSUBS 0.030961f
C400 B.n276 VSUBS 0.012503f
C401 B.n277 VSUBS 0.012503f
C402 B.n278 VSUBS 0.012503f
C403 B.n279 VSUBS 0.012503f
C404 B.n280 VSUBS 0.012503f
C405 B.n281 VSUBS 0.012503f
C406 B.n282 VSUBS 0.012503f
C407 B.n283 VSUBS 0.012503f
C408 B.n284 VSUBS 0.012503f
C409 B.n285 VSUBS 0.012503f
C410 B.n286 VSUBS 0.012503f
C411 B.n287 VSUBS 0.012503f
C412 B.n288 VSUBS 0.012503f
C413 B.n289 VSUBS 0.012503f
C414 B.n290 VSUBS 0.012503f
C415 B.n291 VSUBS 0.012503f
C416 B.n292 VSUBS 0.012503f
C417 B.n293 VSUBS 0.012503f
C418 B.n294 VSUBS 0.012503f
C419 B.n295 VSUBS 0.012503f
C420 B.n296 VSUBS 0.012503f
C421 B.n297 VSUBS 0.012503f
C422 B.n298 VSUBS 0.012503f
C423 B.n299 VSUBS 0.012503f
C424 B.n300 VSUBS 0.012503f
C425 B.n301 VSUBS 0.012503f
C426 B.n302 VSUBS 0.012503f
C427 B.n303 VSUBS 0.012503f
C428 B.n304 VSUBS 0.012503f
C429 B.n305 VSUBS 0.012503f
C430 B.n306 VSUBS 0.012503f
C431 B.n307 VSUBS 0.012503f
C432 B.n308 VSUBS 0.012503f
C433 B.n309 VSUBS 0.012503f
C434 B.n310 VSUBS 0.012503f
C435 B.n311 VSUBS 0.012503f
C436 B.n312 VSUBS 0.012503f
C437 B.n313 VSUBS 0.012503f
C438 B.n314 VSUBS 0.012503f
C439 B.n315 VSUBS 0.012503f
C440 B.n316 VSUBS 0.012503f
C441 B.n317 VSUBS 0.012503f
C442 B.n318 VSUBS 0.012503f
C443 B.n319 VSUBS 0.012503f
C444 B.n320 VSUBS 0.012503f
C445 B.n321 VSUBS 0.012503f
C446 B.n322 VSUBS 0.012503f
C447 B.n323 VSUBS 0.012503f
C448 B.n324 VSUBS 0.012503f
C449 B.n325 VSUBS 0.012503f
C450 B.n326 VSUBS 0.012503f
C451 B.n327 VSUBS 0.012503f
C452 B.n328 VSUBS 0.012503f
C453 B.n329 VSUBS 0.012503f
C454 B.n330 VSUBS 0.012503f
C455 B.n331 VSUBS 0.012503f
C456 B.n332 VSUBS 0.012503f
C457 B.n333 VSUBS 0.012503f
C458 B.n334 VSUBS 0.012503f
C459 B.n335 VSUBS 0.012503f
C460 B.n336 VSUBS 0.012503f
C461 B.n337 VSUBS 0.012503f
C462 B.n338 VSUBS 0.012503f
C463 B.n339 VSUBS 0.012503f
C464 B.n340 VSUBS 0.012503f
C465 B.n341 VSUBS 0.012503f
C466 B.n342 VSUBS 0.012503f
C467 B.n343 VSUBS 0.012503f
C468 B.n344 VSUBS 0.012503f
C469 B.n345 VSUBS 0.012503f
C470 B.n346 VSUBS 0.012503f
C471 B.n347 VSUBS 0.012503f
C472 B.n348 VSUBS 0.012503f
C473 B.n349 VSUBS 0.012503f
C474 B.n350 VSUBS 0.012503f
C475 B.n351 VSUBS 0.012503f
C476 B.n352 VSUBS 0.012503f
C477 B.n353 VSUBS 0.012503f
C478 B.n354 VSUBS 0.012503f
C479 B.n355 VSUBS 0.012503f
C480 B.n356 VSUBS 0.012503f
C481 B.n357 VSUBS 0.012503f
C482 B.n358 VSUBS 0.012503f
C483 B.n359 VSUBS 0.012503f
C484 B.n360 VSUBS 0.012503f
C485 B.n361 VSUBS 0.012503f
C486 B.n362 VSUBS 0.012503f
C487 B.n363 VSUBS 0.012503f
C488 B.n364 VSUBS 0.012503f
C489 B.n365 VSUBS 0.012503f
C490 B.n366 VSUBS 0.012503f
C491 B.n367 VSUBS 0.012503f
C492 B.n368 VSUBS 0.012503f
C493 B.n369 VSUBS 0.012503f
C494 B.n370 VSUBS 0.012503f
C495 B.n371 VSUBS 0.012503f
C496 B.n372 VSUBS 0.012503f
C497 B.n373 VSUBS 0.012503f
C498 B.n374 VSUBS 0.012503f
C499 B.n375 VSUBS 0.012503f
C500 B.n376 VSUBS 0.012503f
C501 B.n377 VSUBS 0.012503f
C502 B.n378 VSUBS 0.012503f
C503 B.n379 VSUBS 0.012503f
C504 B.n380 VSUBS 0.012503f
C505 B.n381 VSUBS 0.012503f
C506 B.n382 VSUBS 0.012503f
C507 B.n383 VSUBS 0.012503f
C508 B.n384 VSUBS 0.012503f
C509 B.n385 VSUBS 0.012503f
C510 B.n386 VSUBS 0.012503f
C511 B.n387 VSUBS 0.012503f
C512 B.n388 VSUBS 0.012503f
C513 B.n389 VSUBS 0.012503f
C514 B.n390 VSUBS 0.012503f
C515 B.n391 VSUBS 0.012503f
C516 B.n392 VSUBS 0.012503f
C517 B.n393 VSUBS 0.012503f
C518 B.n394 VSUBS 0.012503f
C519 B.n395 VSUBS 0.012503f
C520 B.n396 VSUBS 0.012503f
C521 B.n397 VSUBS 0.012503f
C522 B.n398 VSUBS 0.012503f
C523 B.n399 VSUBS 0.012503f
C524 B.n400 VSUBS 0.012503f
C525 B.n401 VSUBS 0.012503f
C526 B.n402 VSUBS 0.012503f
C527 B.n403 VSUBS 0.012503f
C528 B.n404 VSUBS 0.012503f
C529 B.n405 VSUBS 0.012503f
C530 B.n406 VSUBS 0.012503f
C531 B.n407 VSUBS 0.012503f
C532 B.n408 VSUBS 0.012503f
C533 B.n409 VSUBS 0.012503f
C534 B.n410 VSUBS 0.012503f
C535 B.n411 VSUBS 0.012503f
C536 B.n412 VSUBS 0.012503f
C537 B.n413 VSUBS 0.012503f
C538 B.n414 VSUBS 0.012503f
C539 B.n415 VSUBS 0.012503f
C540 B.n416 VSUBS 0.012503f
C541 B.n417 VSUBS 0.012503f
C542 B.n418 VSUBS 0.012503f
C543 B.n419 VSUBS 0.012503f
C544 B.n420 VSUBS 0.012503f
C545 B.n421 VSUBS 0.012503f
C546 B.n422 VSUBS 0.012503f
C547 B.n423 VSUBS 0.012503f
C548 B.n424 VSUBS 0.012503f
C549 B.n425 VSUBS 0.012503f
C550 B.n426 VSUBS 0.012503f
C551 B.n427 VSUBS 0.012503f
C552 B.n428 VSUBS 0.012503f
C553 B.n429 VSUBS 0.012503f
C554 B.n430 VSUBS 0.012503f
C555 B.n431 VSUBS 0.012503f
C556 B.n432 VSUBS 0.012503f
C557 B.n433 VSUBS 0.012503f
C558 B.n434 VSUBS 0.012503f
C559 B.n435 VSUBS 0.012503f
C560 B.n436 VSUBS 0.012503f
C561 B.n437 VSUBS 0.012503f
C562 B.n438 VSUBS 0.012503f
C563 B.n439 VSUBS 0.012503f
C564 B.n440 VSUBS 0.012503f
C565 B.n441 VSUBS 0.029536f
C566 B.n442 VSUBS 0.030405f
C567 B.n443 VSUBS 0.030405f
C568 B.n444 VSUBS 0.012503f
C569 B.n445 VSUBS 0.012503f
C570 B.n446 VSUBS 0.012503f
C571 B.n447 VSUBS 0.012503f
C572 B.n448 VSUBS 0.012503f
C573 B.n449 VSUBS 0.012503f
C574 B.n450 VSUBS 0.012503f
C575 B.n451 VSUBS 0.012503f
C576 B.n452 VSUBS 0.012503f
C577 B.n453 VSUBS 0.012503f
C578 B.n454 VSUBS 0.012503f
C579 B.n455 VSUBS 0.011768f
C580 B.n456 VSUBS 0.028968f
C581 B.n457 VSUBS 0.006987f
C582 B.n458 VSUBS 0.012503f
C583 B.n459 VSUBS 0.012503f
C584 B.n460 VSUBS 0.012503f
C585 B.n461 VSUBS 0.012503f
C586 B.n462 VSUBS 0.012503f
C587 B.n463 VSUBS 0.012503f
C588 B.n464 VSUBS 0.012503f
C589 B.n465 VSUBS 0.012503f
C590 B.n466 VSUBS 0.012503f
C591 B.n467 VSUBS 0.012503f
C592 B.n468 VSUBS 0.012503f
C593 B.n469 VSUBS 0.012503f
C594 B.n470 VSUBS 0.006987f
C595 B.n471 VSUBS 0.012503f
C596 B.n472 VSUBS 0.012503f
C597 B.n473 VSUBS 0.011768f
C598 B.n474 VSUBS 0.012503f
C599 B.n475 VSUBS 0.012503f
C600 B.n476 VSUBS 0.012503f
C601 B.n477 VSUBS 0.012503f
C602 B.n478 VSUBS 0.012503f
C603 B.n479 VSUBS 0.012503f
C604 B.n480 VSUBS 0.012503f
C605 B.n481 VSUBS 0.012503f
C606 B.n482 VSUBS 0.012503f
C607 B.n483 VSUBS 0.012503f
C608 B.n484 VSUBS 0.030405f
C609 B.n485 VSUBS 0.030405f
C610 B.n486 VSUBS 0.029536f
C611 B.n487 VSUBS 0.012503f
C612 B.n488 VSUBS 0.012503f
C613 B.n489 VSUBS 0.012503f
C614 B.n490 VSUBS 0.012503f
C615 B.n491 VSUBS 0.012503f
C616 B.n492 VSUBS 0.012503f
C617 B.n493 VSUBS 0.012503f
C618 B.n494 VSUBS 0.012503f
C619 B.n495 VSUBS 0.012503f
C620 B.n496 VSUBS 0.012503f
C621 B.n497 VSUBS 0.012503f
C622 B.n498 VSUBS 0.012503f
C623 B.n499 VSUBS 0.012503f
C624 B.n500 VSUBS 0.012503f
C625 B.n501 VSUBS 0.012503f
C626 B.n502 VSUBS 0.012503f
C627 B.n503 VSUBS 0.012503f
C628 B.n504 VSUBS 0.012503f
C629 B.n505 VSUBS 0.012503f
C630 B.n506 VSUBS 0.012503f
C631 B.n507 VSUBS 0.012503f
C632 B.n508 VSUBS 0.012503f
C633 B.n509 VSUBS 0.012503f
C634 B.n510 VSUBS 0.012503f
C635 B.n511 VSUBS 0.012503f
C636 B.n512 VSUBS 0.012503f
C637 B.n513 VSUBS 0.012503f
C638 B.n514 VSUBS 0.012503f
C639 B.n515 VSUBS 0.012503f
C640 B.n516 VSUBS 0.012503f
C641 B.n517 VSUBS 0.012503f
C642 B.n518 VSUBS 0.012503f
C643 B.n519 VSUBS 0.012503f
C644 B.n520 VSUBS 0.012503f
C645 B.n521 VSUBS 0.012503f
C646 B.n522 VSUBS 0.012503f
C647 B.n523 VSUBS 0.012503f
C648 B.n524 VSUBS 0.012503f
C649 B.n525 VSUBS 0.012503f
C650 B.n526 VSUBS 0.012503f
C651 B.n527 VSUBS 0.012503f
C652 B.n528 VSUBS 0.012503f
C653 B.n529 VSUBS 0.012503f
C654 B.n530 VSUBS 0.012503f
C655 B.n531 VSUBS 0.012503f
C656 B.n532 VSUBS 0.012503f
C657 B.n533 VSUBS 0.012503f
C658 B.n534 VSUBS 0.012503f
C659 B.n535 VSUBS 0.012503f
C660 B.n536 VSUBS 0.012503f
C661 B.n537 VSUBS 0.012503f
C662 B.n538 VSUBS 0.012503f
C663 B.n539 VSUBS 0.012503f
C664 B.n540 VSUBS 0.012503f
C665 B.n541 VSUBS 0.012503f
C666 B.n542 VSUBS 0.012503f
C667 B.n543 VSUBS 0.012503f
C668 B.n544 VSUBS 0.012503f
C669 B.n545 VSUBS 0.012503f
C670 B.n546 VSUBS 0.012503f
C671 B.n547 VSUBS 0.012503f
C672 B.n548 VSUBS 0.012503f
C673 B.n549 VSUBS 0.012503f
C674 B.n550 VSUBS 0.012503f
C675 B.n551 VSUBS 0.012503f
C676 B.n552 VSUBS 0.012503f
C677 B.n553 VSUBS 0.012503f
C678 B.n554 VSUBS 0.012503f
C679 B.n555 VSUBS 0.012503f
C680 B.n556 VSUBS 0.012503f
C681 B.n557 VSUBS 0.012503f
C682 B.n558 VSUBS 0.012503f
C683 B.n559 VSUBS 0.012503f
C684 B.n560 VSUBS 0.012503f
C685 B.n561 VSUBS 0.012503f
C686 B.n562 VSUBS 0.012503f
C687 B.n563 VSUBS 0.012503f
C688 B.n564 VSUBS 0.012503f
C689 B.n565 VSUBS 0.012503f
C690 B.n566 VSUBS 0.012503f
C691 B.n567 VSUBS 0.016316f
C692 B.n568 VSUBS 0.017381f
C693 B.n569 VSUBS 0.034563f
C694 VDD1.t1 VSUBS 0.015482f
C695 VDD1.t2 VSUBS 0.015482f
C696 VDD1.n0 VSUBS 0.052985f
C697 VDD1.t5 VSUBS 0.015482f
C698 VDD1.t0 VSUBS 0.015482f
C699 VDD1.n1 VSUBS 0.052827f
C700 VDD1.t3 VSUBS 0.015482f
C701 VDD1.t7 VSUBS 0.015482f
C702 VDD1.n2 VSUBS 0.052827f
C703 VDD1.n3 VSUBS 2.12419f
C704 VDD1.t4 VSUBS 0.015482f
C705 VDD1.t6 VSUBS 0.015482f
C706 VDD1.n4 VSUBS 0.051283f
C707 VDD1.n5 VSUBS 1.66741f
C708 VTAIL.t7 VSUBS 0.031296f
C709 VTAIL.t4 VSUBS 0.031296f
C710 VTAIL.n0 VSUBS 0.089254f
C711 VTAIL.n1 VSUBS 0.601409f
C712 VTAIL.t5 VSUBS 0.157215f
C713 VTAIL.n2 VSUBS 0.669309f
C714 VTAIL.t11 VSUBS 0.157215f
C715 VTAIL.n3 VSUBS 0.669309f
C716 VTAIL.t13 VSUBS 0.031296f
C717 VTAIL.t10 VSUBS 0.031296f
C718 VTAIL.n4 VSUBS 0.089254f
C719 VTAIL.n5 VSUBS 0.934873f
C720 VTAIL.t8 VSUBS 0.157215f
C721 VTAIL.n6 VSUBS 1.57954f
C722 VTAIL.t0 VSUBS 0.157215f
C723 VTAIL.n7 VSUBS 1.57954f
C724 VTAIL.t2 VSUBS 0.031296f
C725 VTAIL.t6 VSUBS 0.031296f
C726 VTAIL.n8 VSUBS 0.089254f
C727 VTAIL.n9 VSUBS 0.934873f
C728 VTAIL.t3 VSUBS 0.157215f
C729 VTAIL.n10 VSUBS 0.669309f
C730 VTAIL.t15 VSUBS 0.157215f
C731 VTAIL.n11 VSUBS 0.669309f
C732 VTAIL.t12 VSUBS 0.031296f
C733 VTAIL.t14 VSUBS 0.031296f
C734 VTAIL.n12 VSUBS 0.089254f
C735 VTAIL.n13 VSUBS 0.934873f
C736 VTAIL.t9 VSUBS 0.157215f
C737 VTAIL.n14 VSUBS 1.57954f
C738 VTAIL.t1 VSUBS 0.157215f
C739 VTAIL.n15 VSUBS 1.5724f
C740 VP.n0 VSUBS 0.088417f
C741 VP.t0 VSUBS 0.383856f
C742 VP.n1 VSUBS 0.134177f
C743 VP.n2 VSUBS 0.067068f
C744 VP.n3 VSUBS 0.080164f
C745 VP.n4 VSUBS 0.067068f
C746 VP.n5 VSUBS 0.097494f
C747 VP.n6 VSUBS 0.067068f
C748 VP.t7 VSUBS 0.383856f
C749 VP.n7 VSUBS 0.124371f
C750 VP.n8 VSUBS 0.067068f
C751 VP.n9 VSUBS 0.124371f
C752 VP.n10 VSUBS 0.088417f
C753 VP.t1 VSUBS 0.383856f
C754 VP.n11 VSUBS 0.134177f
C755 VP.n12 VSUBS 0.067068f
C756 VP.n13 VSUBS 0.080164f
C757 VP.n14 VSUBS 0.067068f
C758 VP.n15 VSUBS 0.097494f
C759 VP.n16 VSUBS 0.710374f
C760 VP.t5 VSUBS 0.383856f
C761 VP.t6 VSUBS 0.943698f
C762 VP.n17 VSUBS 0.479068f
C763 VP.n18 VSUBS 0.471068f
C764 VP.n19 VSUBS 0.10718f
C765 VP.n20 VSUBS 0.124371f
C766 VP.n21 VSUBS 0.067068f
C767 VP.n22 VSUBS 0.067068f
C768 VP.n23 VSUBS 0.067068f
C769 VP.n24 VSUBS 0.097494f
C770 VP.n25 VSUBS 0.124371f
C771 VP.t3 VSUBS 0.383856f
C772 VP.n26 VSUBS 0.249705f
C773 VP.n27 VSUBS 0.10718f
C774 VP.n28 VSUBS 0.067068f
C775 VP.n29 VSUBS 0.067068f
C776 VP.n30 VSUBS 0.067068f
C777 VP.n31 VSUBS 0.124371f
C778 VP.n32 VSUBS 0.13024f
C779 VP.n33 VSUBS 0.054942f
C780 VP.n34 VSUBS 0.067068f
C781 VP.n35 VSUBS 0.067068f
C782 VP.n36 VSUBS 0.067068f
C783 VP.n37 VSUBS 0.124371f
C784 VP.n38 VSUBS 0.072796f
C785 VP.n39 VSUBS 0.476499f
C786 VP.n40 VSUBS 3.0852f
C787 VP.n41 VSUBS 3.14021f
C788 VP.t2 VSUBS 0.383856f
C789 VP.n42 VSUBS 0.476499f
C790 VP.n43 VSUBS 0.072796f
C791 VP.n44 VSUBS 0.088417f
C792 VP.n45 VSUBS 0.067068f
C793 VP.n46 VSUBS 0.067068f
C794 VP.n47 VSUBS 0.134177f
C795 VP.n48 VSUBS 0.054942f
C796 VP.n49 VSUBS 0.13024f
C797 VP.n50 VSUBS 0.067068f
C798 VP.n51 VSUBS 0.067068f
C799 VP.n52 VSUBS 0.067068f
C800 VP.n53 VSUBS 0.080164f
C801 VP.n54 VSUBS 0.249705f
C802 VP.n55 VSUBS 0.10718f
C803 VP.n56 VSUBS 0.124371f
C804 VP.n57 VSUBS 0.067068f
C805 VP.n58 VSUBS 0.067068f
C806 VP.n59 VSUBS 0.067068f
C807 VP.n60 VSUBS 0.097494f
C808 VP.n61 VSUBS 0.124371f
C809 VP.t4 VSUBS 0.383856f
C810 VP.n62 VSUBS 0.249705f
C811 VP.n63 VSUBS 0.10718f
C812 VP.n64 VSUBS 0.067068f
C813 VP.n65 VSUBS 0.067068f
C814 VP.n66 VSUBS 0.067068f
C815 VP.n67 VSUBS 0.124371f
C816 VP.n68 VSUBS 0.13024f
C817 VP.n69 VSUBS 0.054942f
C818 VP.n70 VSUBS 0.067068f
C819 VP.n71 VSUBS 0.067068f
C820 VP.n72 VSUBS 0.067068f
C821 VP.n73 VSUBS 0.124371f
C822 VP.n74 VSUBS 0.072796f
C823 VP.n75 VSUBS 0.476499f
C824 VP.n76 VSUBS 0.125854f
.ends

