* NGSPICE file created from diff_pair_sample_1670.ext - technology: sky130A

.subckt diff_pair_sample_1670 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=0 ps=0 w=11.48 l=1.91
X1 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=0 ps=0 w=11.48 l=1.91
X2 VDD1.t5 VP.t0 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=1.8942 ps=11.81 w=11.48 l=1.91
X3 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=4.4772 ps=23.74 w=11.48 l=1.91
X4 VDD1.t4 VP.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=1.8942 ps=11.81 w=11.48 l=1.91
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=0 ps=0 w=11.48 l=1.91
X6 VTAIL.t5 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=1.8942 ps=11.81 w=11.48 l=1.91
X7 VDD2.t4 VN.t1 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=1.8942 ps=11.81 w=11.48 l=1.91
X8 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=0 ps=0 w=11.48 l=1.91
X9 VDD2.t3 VN.t2 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=4.4772 ps=23.74 w=11.48 l=1.91
X10 VTAIL.t2 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=1.8942 ps=11.81 w=11.48 l=1.91
X11 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4772 pd=23.74 as=1.8942 ps=11.81 w=11.48 l=1.91
X12 VDD1.t2 VP.t3 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=4.4772 ps=23.74 w=11.48 l=1.91
X13 VTAIL.t4 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=1.8942 ps=11.81 w=11.48 l=1.91
X14 VDD1.t1 VP.t4 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=4.4772 ps=23.74 w=11.48 l=1.91
X15 VTAIL.t8 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8942 pd=11.81 as=1.8942 ps=11.81 w=11.48 l=1.91
R0 B.n560 B.n559 585
R1 B.n562 B.n115 585
R2 B.n565 B.n564 585
R3 B.n566 B.n114 585
R4 B.n568 B.n567 585
R5 B.n570 B.n113 585
R6 B.n573 B.n572 585
R7 B.n574 B.n112 585
R8 B.n576 B.n575 585
R9 B.n578 B.n111 585
R10 B.n581 B.n580 585
R11 B.n582 B.n110 585
R12 B.n584 B.n583 585
R13 B.n586 B.n109 585
R14 B.n589 B.n588 585
R15 B.n590 B.n108 585
R16 B.n592 B.n591 585
R17 B.n594 B.n107 585
R18 B.n597 B.n596 585
R19 B.n598 B.n106 585
R20 B.n600 B.n599 585
R21 B.n602 B.n105 585
R22 B.n605 B.n604 585
R23 B.n606 B.n104 585
R24 B.n608 B.n607 585
R25 B.n610 B.n103 585
R26 B.n613 B.n612 585
R27 B.n614 B.n102 585
R28 B.n616 B.n615 585
R29 B.n618 B.n101 585
R30 B.n621 B.n620 585
R31 B.n622 B.n100 585
R32 B.n624 B.n623 585
R33 B.n626 B.n99 585
R34 B.n629 B.n628 585
R35 B.n630 B.n98 585
R36 B.n632 B.n631 585
R37 B.n634 B.n97 585
R38 B.n636 B.n635 585
R39 B.n638 B.n637 585
R40 B.n641 B.n640 585
R41 B.n642 B.n92 585
R42 B.n644 B.n643 585
R43 B.n646 B.n91 585
R44 B.n649 B.n648 585
R45 B.n650 B.n90 585
R46 B.n652 B.n651 585
R47 B.n654 B.n89 585
R48 B.n657 B.n656 585
R49 B.n658 B.n86 585
R50 B.n661 B.n660 585
R51 B.n663 B.n85 585
R52 B.n666 B.n665 585
R53 B.n667 B.n84 585
R54 B.n669 B.n668 585
R55 B.n671 B.n83 585
R56 B.n674 B.n673 585
R57 B.n675 B.n82 585
R58 B.n677 B.n676 585
R59 B.n679 B.n81 585
R60 B.n682 B.n681 585
R61 B.n683 B.n80 585
R62 B.n685 B.n684 585
R63 B.n687 B.n79 585
R64 B.n690 B.n689 585
R65 B.n691 B.n78 585
R66 B.n693 B.n692 585
R67 B.n695 B.n77 585
R68 B.n698 B.n697 585
R69 B.n699 B.n76 585
R70 B.n701 B.n700 585
R71 B.n703 B.n75 585
R72 B.n706 B.n705 585
R73 B.n707 B.n74 585
R74 B.n709 B.n708 585
R75 B.n711 B.n73 585
R76 B.n714 B.n713 585
R77 B.n715 B.n72 585
R78 B.n717 B.n716 585
R79 B.n719 B.n71 585
R80 B.n722 B.n721 585
R81 B.n723 B.n70 585
R82 B.n725 B.n724 585
R83 B.n727 B.n69 585
R84 B.n730 B.n729 585
R85 B.n731 B.n68 585
R86 B.n733 B.n732 585
R87 B.n735 B.n67 585
R88 B.n738 B.n737 585
R89 B.n739 B.n66 585
R90 B.n558 B.n64 585
R91 B.n742 B.n64 585
R92 B.n557 B.n63 585
R93 B.n743 B.n63 585
R94 B.n556 B.n62 585
R95 B.n744 B.n62 585
R96 B.n555 B.n554 585
R97 B.n554 B.n58 585
R98 B.n553 B.n57 585
R99 B.n750 B.n57 585
R100 B.n552 B.n56 585
R101 B.n751 B.n56 585
R102 B.n551 B.n55 585
R103 B.n752 B.n55 585
R104 B.n550 B.n549 585
R105 B.n549 B.n51 585
R106 B.n548 B.n50 585
R107 B.n758 B.n50 585
R108 B.n547 B.n49 585
R109 B.n759 B.n49 585
R110 B.n546 B.n48 585
R111 B.n760 B.n48 585
R112 B.n545 B.n544 585
R113 B.n544 B.n44 585
R114 B.n543 B.n43 585
R115 B.n766 B.n43 585
R116 B.n542 B.n42 585
R117 B.n767 B.n42 585
R118 B.n541 B.n41 585
R119 B.n768 B.n41 585
R120 B.n540 B.n539 585
R121 B.n539 B.n37 585
R122 B.n538 B.n36 585
R123 B.n774 B.n36 585
R124 B.n537 B.n35 585
R125 B.n775 B.n35 585
R126 B.n536 B.n34 585
R127 B.n776 B.n34 585
R128 B.n535 B.n534 585
R129 B.n534 B.n30 585
R130 B.n533 B.n29 585
R131 B.n782 B.n29 585
R132 B.n532 B.n28 585
R133 B.n783 B.n28 585
R134 B.n531 B.n27 585
R135 B.n784 B.n27 585
R136 B.n530 B.n529 585
R137 B.n529 B.n26 585
R138 B.n528 B.n22 585
R139 B.n790 B.n22 585
R140 B.n527 B.n21 585
R141 B.n791 B.n21 585
R142 B.n526 B.n20 585
R143 B.n792 B.n20 585
R144 B.n525 B.n524 585
R145 B.n524 B.n16 585
R146 B.n523 B.n15 585
R147 B.n798 B.n15 585
R148 B.n522 B.n14 585
R149 B.n799 B.n14 585
R150 B.n521 B.n13 585
R151 B.n800 B.n13 585
R152 B.n520 B.n519 585
R153 B.n519 B.n12 585
R154 B.n518 B.n517 585
R155 B.n518 B.n8 585
R156 B.n516 B.n7 585
R157 B.n807 B.n7 585
R158 B.n515 B.n6 585
R159 B.n808 B.n6 585
R160 B.n514 B.n5 585
R161 B.n809 B.n5 585
R162 B.n513 B.n512 585
R163 B.n512 B.n4 585
R164 B.n511 B.n116 585
R165 B.n511 B.n510 585
R166 B.n501 B.n117 585
R167 B.n118 B.n117 585
R168 B.n503 B.n502 585
R169 B.n504 B.n503 585
R170 B.n500 B.n122 585
R171 B.n126 B.n122 585
R172 B.n499 B.n498 585
R173 B.n498 B.n497 585
R174 B.n124 B.n123 585
R175 B.n125 B.n124 585
R176 B.n490 B.n489 585
R177 B.n491 B.n490 585
R178 B.n488 B.n131 585
R179 B.n131 B.n130 585
R180 B.n487 B.n486 585
R181 B.n486 B.n485 585
R182 B.n133 B.n132 585
R183 B.n478 B.n133 585
R184 B.n477 B.n476 585
R185 B.n479 B.n477 585
R186 B.n475 B.n138 585
R187 B.n138 B.n137 585
R188 B.n474 B.n473 585
R189 B.n473 B.n472 585
R190 B.n140 B.n139 585
R191 B.n141 B.n140 585
R192 B.n465 B.n464 585
R193 B.n466 B.n465 585
R194 B.n463 B.n146 585
R195 B.n146 B.n145 585
R196 B.n462 B.n461 585
R197 B.n461 B.n460 585
R198 B.n148 B.n147 585
R199 B.n149 B.n148 585
R200 B.n453 B.n452 585
R201 B.n454 B.n453 585
R202 B.n451 B.n154 585
R203 B.n154 B.n153 585
R204 B.n450 B.n449 585
R205 B.n449 B.n448 585
R206 B.n156 B.n155 585
R207 B.n157 B.n156 585
R208 B.n441 B.n440 585
R209 B.n442 B.n441 585
R210 B.n439 B.n162 585
R211 B.n162 B.n161 585
R212 B.n438 B.n437 585
R213 B.n437 B.n436 585
R214 B.n164 B.n163 585
R215 B.n165 B.n164 585
R216 B.n429 B.n428 585
R217 B.n430 B.n429 585
R218 B.n427 B.n170 585
R219 B.n170 B.n169 585
R220 B.n426 B.n425 585
R221 B.n425 B.n424 585
R222 B.n172 B.n171 585
R223 B.n173 B.n172 585
R224 B.n417 B.n416 585
R225 B.n418 B.n417 585
R226 B.n415 B.n178 585
R227 B.n178 B.n177 585
R228 B.n414 B.n413 585
R229 B.n413 B.n412 585
R230 B.n409 B.n182 585
R231 B.n408 B.n407 585
R232 B.n405 B.n183 585
R233 B.n405 B.n181 585
R234 B.n404 B.n403 585
R235 B.n402 B.n401 585
R236 B.n400 B.n185 585
R237 B.n398 B.n397 585
R238 B.n396 B.n186 585
R239 B.n395 B.n394 585
R240 B.n392 B.n187 585
R241 B.n390 B.n389 585
R242 B.n388 B.n188 585
R243 B.n387 B.n386 585
R244 B.n384 B.n189 585
R245 B.n382 B.n381 585
R246 B.n380 B.n190 585
R247 B.n379 B.n378 585
R248 B.n376 B.n191 585
R249 B.n374 B.n373 585
R250 B.n372 B.n192 585
R251 B.n371 B.n370 585
R252 B.n368 B.n193 585
R253 B.n366 B.n365 585
R254 B.n364 B.n194 585
R255 B.n363 B.n362 585
R256 B.n360 B.n195 585
R257 B.n358 B.n357 585
R258 B.n356 B.n196 585
R259 B.n355 B.n354 585
R260 B.n352 B.n197 585
R261 B.n350 B.n349 585
R262 B.n348 B.n198 585
R263 B.n347 B.n346 585
R264 B.n344 B.n199 585
R265 B.n342 B.n341 585
R266 B.n340 B.n200 585
R267 B.n339 B.n338 585
R268 B.n336 B.n201 585
R269 B.n334 B.n333 585
R270 B.n332 B.n202 585
R271 B.n330 B.n329 585
R272 B.n327 B.n205 585
R273 B.n325 B.n324 585
R274 B.n323 B.n206 585
R275 B.n322 B.n321 585
R276 B.n319 B.n207 585
R277 B.n317 B.n316 585
R278 B.n315 B.n208 585
R279 B.n314 B.n313 585
R280 B.n311 B.n209 585
R281 B.n309 B.n308 585
R282 B.n307 B.n210 585
R283 B.n306 B.n305 585
R284 B.n303 B.n214 585
R285 B.n301 B.n300 585
R286 B.n299 B.n215 585
R287 B.n298 B.n297 585
R288 B.n295 B.n216 585
R289 B.n293 B.n292 585
R290 B.n291 B.n217 585
R291 B.n290 B.n289 585
R292 B.n287 B.n218 585
R293 B.n285 B.n284 585
R294 B.n283 B.n219 585
R295 B.n282 B.n281 585
R296 B.n279 B.n220 585
R297 B.n277 B.n276 585
R298 B.n275 B.n221 585
R299 B.n274 B.n273 585
R300 B.n271 B.n222 585
R301 B.n269 B.n268 585
R302 B.n267 B.n223 585
R303 B.n266 B.n265 585
R304 B.n263 B.n224 585
R305 B.n261 B.n260 585
R306 B.n259 B.n225 585
R307 B.n258 B.n257 585
R308 B.n255 B.n226 585
R309 B.n253 B.n252 585
R310 B.n251 B.n227 585
R311 B.n250 B.n249 585
R312 B.n247 B.n228 585
R313 B.n245 B.n244 585
R314 B.n243 B.n229 585
R315 B.n242 B.n241 585
R316 B.n239 B.n230 585
R317 B.n237 B.n236 585
R318 B.n235 B.n231 585
R319 B.n234 B.n233 585
R320 B.n180 B.n179 585
R321 B.n181 B.n180 585
R322 B.n411 B.n410 585
R323 B.n412 B.n411 585
R324 B.n176 B.n175 585
R325 B.n177 B.n176 585
R326 B.n420 B.n419 585
R327 B.n419 B.n418 585
R328 B.n421 B.n174 585
R329 B.n174 B.n173 585
R330 B.n423 B.n422 585
R331 B.n424 B.n423 585
R332 B.n168 B.n167 585
R333 B.n169 B.n168 585
R334 B.n432 B.n431 585
R335 B.n431 B.n430 585
R336 B.n433 B.n166 585
R337 B.n166 B.n165 585
R338 B.n435 B.n434 585
R339 B.n436 B.n435 585
R340 B.n160 B.n159 585
R341 B.n161 B.n160 585
R342 B.n444 B.n443 585
R343 B.n443 B.n442 585
R344 B.n445 B.n158 585
R345 B.n158 B.n157 585
R346 B.n447 B.n446 585
R347 B.n448 B.n447 585
R348 B.n152 B.n151 585
R349 B.n153 B.n152 585
R350 B.n456 B.n455 585
R351 B.n455 B.n454 585
R352 B.n457 B.n150 585
R353 B.n150 B.n149 585
R354 B.n459 B.n458 585
R355 B.n460 B.n459 585
R356 B.n144 B.n143 585
R357 B.n145 B.n144 585
R358 B.n468 B.n467 585
R359 B.n467 B.n466 585
R360 B.n469 B.n142 585
R361 B.n142 B.n141 585
R362 B.n471 B.n470 585
R363 B.n472 B.n471 585
R364 B.n136 B.n135 585
R365 B.n137 B.n136 585
R366 B.n481 B.n480 585
R367 B.n480 B.n479 585
R368 B.n482 B.n134 585
R369 B.n478 B.n134 585
R370 B.n484 B.n483 585
R371 B.n485 B.n484 585
R372 B.n129 B.n128 585
R373 B.n130 B.n129 585
R374 B.n493 B.n492 585
R375 B.n492 B.n491 585
R376 B.n494 B.n127 585
R377 B.n127 B.n125 585
R378 B.n496 B.n495 585
R379 B.n497 B.n496 585
R380 B.n121 B.n120 585
R381 B.n126 B.n121 585
R382 B.n506 B.n505 585
R383 B.n505 B.n504 585
R384 B.n507 B.n119 585
R385 B.n119 B.n118 585
R386 B.n509 B.n508 585
R387 B.n510 B.n509 585
R388 B.n3 B.n0 585
R389 B.n4 B.n3 585
R390 B.n806 B.n1 585
R391 B.n807 B.n806 585
R392 B.n805 B.n804 585
R393 B.n805 B.n8 585
R394 B.n803 B.n9 585
R395 B.n12 B.n9 585
R396 B.n802 B.n801 585
R397 B.n801 B.n800 585
R398 B.n11 B.n10 585
R399 B.n799 B.n11 585
R400 B.n797 B.n796 585
R401 B.n798 B.n797 585
R402 B.n795 B.n17 585
R403 B.n17 B.n16 585
R404 B.n794 B.n793 585
R405 B.n793 B.n792 585
R406 B.n19 B.n18 585
R407 B.n791 B.n19 585
R408 B.n789 B.n788 585
R409 B.n790 B.n789 585
R410 B.n787 B.n23 585
R411 B.n26 B.n23 585
R412 B.n786 B.n785 585
R413 B.n785 B.n784 585
R414 B.n25 B.n24 585
R415 B.n783 B.n25 585
R416 B.n781 B.n780 585
R417 B.n782 B.n781 585
R418 B.n779 B.n31 585
R419 B.n31 B.n30 585
R420 B.n778 B.n777 585
R421 B.n777 B.n776 585
R422 B.n33 B.n32 585
R423 B.n775 B.n33 585
R424 B.n773 B.n772 585
R425 B.n774 B.n773 585
R426 B.n771 B.n38 585
R427 B.n38 B.n37 585
R428 B.n770 B.n769 585
R429 B.n769 B.n768 585
R430 B.n40 B.n39 585
R431 B.n767 B.n40 585
R432 B.n765 B.n764 585
R433 B.n766 B.n765 585
R434 B.n763 B.n45 585
R435 B.n45 B.n44 585
R436 B.n762 B.n761 585
R437 B.n761 B.n760 585
R438 B.n47 B.n46 585
R439 B.n759 B.n47 585
R440 B.n757 B.n756 585
R441 B.n758 B.n757 585
R442 B.n755 B.n52 585
R443 B.n52 B.n51 585
R444 B.n754 B.n753 585
R445 B.n753 B.n752 585
R446 B.n54 B.n53 585
R447 B.n751 B.n54 585
R448 B.n749 B.n748 585
R449 B.n750 B.n749 585
R450 B.n747 B.n59 585
R451 B.n59 B.n58 585
R452 B.n746 B.n745 585
R453 B.n745 B.n744 585
R454 B.n61 B.n60 585
R455 B.n743 B.n61 585
R456 B.n741 B.n740 585
R457 B.n742 B.n741 585
R458 B.n810 B.n809 585
R459 B.n808 B.n2 585
R460 B.n741 B.n66 473.281
R461 B.n560 B.n64 473.281
R462 B.n413 B.n180 473.281
R463 B.n411 B.n182 473.281
R464 B.n87 B.t13 351.551
R465 B.n93 B.t17 351.551
R466 B.n211 B.t6 351.551
R467 B.n203 B.t10 351.551
R468 B.n93 B.t18 316.841
R469 B.n211 B.t9 316.841
R470 B.n87 B.t15 316.841
R471 B.n203 B.t12 316.841
R472 B.n94 B.t19 273.399
R473 B.n212 B.t8 273.399
R474 B.n88 B.t16 273.399
R475 B.n204 B.t11 273.399
R476 B.n561 B.n65 256.663
R477 B.n563 B.n65 256.663
R478 B.n569 B.n65 256.663
R479 B.n571 B.n65 256.663
R480 B.n577 B.n65 256.663
R481 B.n579 B.n65 256.663
R482 B.n585 B.n65 256.663
R483 B.n587 B.n65 256.663
R484 B.n593 B.n65 256.663
R485 B.n595 B.n65 256.663
R486 B.n601 B.n65 256.663
R487 B.n603 B.n65 256.663
R488 B.n609 B.n65 256.663
R489 B.n611 B.n65 256.663
R490 B.n617 B.n65 256.663
R491 B.n619 B.n65 256.663
R492 B.n625 B.n65 256.663
R493 B.n627 B.n65 256.663
R494 B.n633 B.n65 256.663
R495 B.n96 B.n65 256.663
R496 B.n639 B.n65 256.663
R497 B.n645 B.n65 256.663
R498 B.n647 B.n65 256.663
R499 B.n653 B.n65 256.663
R500 B.n655 B.n65 256.663
R501 B.n662 B.n65 256.663
R502 B.n664 B.n65 256.663
R503 B.n670 B.n65 256.663
R504 B.n672 B.n65 256.663
R505 B.n678 B.n65 256.663
R506 B.n680 B.n65 256.663
R507 B.n686 B.n65 256.663
R508 B.n688 B.n65 256.663
R509 B.n694 B.n65 256.663
R510 B.n696 B.n65 256.663
R511 B.n702 B.n65 256.663
R512 B.n704 B.n65 256.663
R513 B.n710 B.n65 256.663
R514 B.n712 B.n65 256.663
R515 B.n718 B.n65 256.663
R516 B.n720 B.n65 256.663
R517 B.n726 B.n65 256.663
R518 B.n728 B.n65 256.663
R519 B.n734 B.n65 256.663
R520 B.n736 B.n65 256.663
R521 B.n406 B.n181 256.663
R522 B.n184 B.n181 256.663
R523 B.n399 B.n181 256.663
R524 B.n393 B.n181 256.663
R525 B.n391 B.n181 256.663
R526 B.n385 B.n181 256.663
R527 B.n383 B.n181 256.663
R528 B.n377 B.n181 256.663
R529 B.n375 B.n181 256.663
R530 B.n369 B.n181 256.663
R531 B.n367 B.n181 256.663
R532 B.n361 B.n181 256.663
R533 B.n359 B.n181 256.663
R534 B.n353 B.n181 256.663
R535 B.n351 B.n181 256.663
R536 B.n345 B.n181 256.663
R537 B.n343 B.n181 256.663
R538 B.n337 B.n181 256.663
R539 B.n335 B.n181 256.663
R540 B.n328 B.n181 256.663
R541 B.n326 B.n181 256.663
R542 B.n320 B.n181 256.663
R543 B.n318 B.n181 256.663
R544 B.n312 B.n181 256.663
R545 B.n310 B.n181 256.663
R546 B.n304 B.n181 256.663
R547 B.n302 B.n181 256.663
R548 B.n296 B.n181 256.663
R549 B.n294 B.n181 256.663
R550 B.n288 B.n181 256.663
R551 B.n286 B.n181 256.663
R552 B.n280 B.n181 256.663
R553 B.n278 B.n181 256.663
R554 B.n272 B.n181 256.663
R555 B.n270 B.n181 256.663
R556 B.n264 B.n181 256.663
R557 B.n262 B.n181 256.663
R558 B.n256 B.n181 256.663
R559 B.n254 B.n181 256.663
R560 B.n248 B.n181 256.663
R561 B.n246 B.n181 256.663
R562 B.n240 B.n181 256.663
R563 B.n238 B.n181 256.663
R564 B.n232 B.n181 256.663
R565 B.n812 B.n811 256.663
R566 B.n737 B.n735 163.367
R567 B.n733 B.n68 163.367
R568 B.n729 B.n727 163.367
R569 B.n725 B.n70 163.367
R570 B.n721 B.n719 163.367
R571 B.n717 B.n72 163.367
R572 B.n713 B.n711 163.367
R573 B.n709 B.n74 163.367
R574 B.n705 B.n703 163.367
R575 B.n701 B.n76 163.367
R576 B.n697 B.n695 163.367
R577 B.n693 B.n78 163.367
R578 B.n689 B.n687 163.367
R579 B.n685 B.n80 163.367
R580 B.n681 B.n679 163.367
R581 B.n677 B.n82 163.367
R582 B.n673 B.n671 163.367
R583 B.n669 B.n84 163.367
R584 B.n665 B.n663 163.367
R585 B.n661 B.n86 163.367
R586 B.n656 B.n654 163.367
R587 B.n652 B.n90 163.367
R588 B.n648 B.n646 163.367
R589 B.n644 B.n92 163.367
R590 B.n640 B.n638 163.367
R591 B.n635 B.n634 163.367
R592 B.n632 B.n98 163.367
R593 B.n628 B.n626 163.367
R594 B.n624 B.n100 163.367
R595 B.n620 B.n618 163.367
R596 B.n616 B.n102 163.367
R597 B.n612 B.n610 163.367
R598 B.n608 B.n104 163.367
R599 B.n604 B.n602 163.367
R600 B.n600 B.n106 163.367
R601 B.n596 B.n594 163.367
R602 B.n592 B.n108 163.367
R603 B.n588 B.n586 163.367
R604 B.n584 B.n110 163.367
R605 B.n580 B.n578 163.367
R606 B.n576 B.n112 163.367
R607 B.n572 B.n570 163.367
R608 B.n568 B.n114 163.367
R609 B.n564 B.n562 163.367
R610 B.n413 B.n178 163.367
R611 B.n417 B.n178 163.367
R612 B.n417 B.n172 163.367
R613 B.n425 B.n172 163.367
R614 B.n425 B.n170 163.367
R615 B.n429 B.n170 163.367
R616 B.n429 B.n164 163.367
R617 B.n437 B.n164 163.367
R618 B.n437 B.n162 163.367
R619 B.n441 B.n162 163.367
R620 B.n441 B.n156 163.367
R621 B.n449 B.n156 163.367
R622 B.n449 B.n154 163.367
R623 B.n453 B.n154 163.367
R624 B.n453 B.n148 163.367
R625 B.n461 B.n148 163.367
R626 B.n461 B.n146 163.367
R627 B.n465 B.n146 163.367
R628 B.n465 B.n140 163.367
R629 B.n473 B.n140 163.367
R630 B.n473 B.n138 163.367
R631 B.n477 B.n138 163.367
R632 B.n477 B.n133 163.367
R633 B.n486 B.n133 163.367
R634 B.n486 B.n131 163.367
R635 B.n490 B.n131 163.367
R636 B.n490 B.n124 163.367
R637 B.n498 B.n124 163.367
R638 B.n498 B.n122 163.367
R639 B.n503 B.n122 163.367
R640 B.n503 B.n117 163.367
R641 B.n511 B.n117 163.367
R642 B.n512 B.n511 163.367
R643 B.n512 B.n5 163.367
R644 B.n6 B.n5 163.367
R645 B.n7 B.n6 163.367
R646 B.n518 B.n7 163.367
R647 B.n519 B.n518 163.367
R648 B.n519 B.n13 163.367
R649 B.n14 B.n13 163.367
R650 B.n15 B.n14 163.367
R651 B.n524 B.n15 163.367
R652 B.n524 B.n20 163.367
R653 B.n21 B.n20 163.367
R654 B.n22 B.n21 163.367
R655 B.n529 B.n22 163.367
R656 B.n529 B.n27 163.367
R657 B.n28 B.n27 163.367
R658 B.n29 B.n28 163.367
R659 B.n534 B.n29 163.367
R660 B.n534 B.n34 163.367
R661 B.n35 B.n34 163.367
R662 B.n36 B.n35 163.367
R663 B.n539 B.n36 163.367
R664 B.n539 B.n41 163.367
R665 B.n42 B.n41 163.367
R666 B.n43 B.n42 163.367
R667 B.n544 B.n43 163.367
R668 B.n544 B.n48 163.367
R669 B.n49 B.n48 163.367
R670 B.n50 B.n49 163.367
R671 B.n549 B.n50 163.367
R672 B.n549 B.n55 163.367
R673 B.n56 B.n55 163.367
R674 B.n57 B.n56 163.367
R675 B.n554 B.n57 163.367
R676 B.n554 B.n62 163.367
R677 B.n63 B.n62 163.367
R678 B.n64 B.n63 163.367
R679 B.n407 B.n405 163.367
R680 B.n405 B.n404 163.367
R681 B.n401 B.n400 163.367
R682 B.n398 B.n186 163.367
R683 B.n394 B.n392 163.367
R684 B.n390 B.n188 163.367
R685 B.n386 B.n384 163.367
R686 B.n382 B.n190 163.367
R687 B.n378 B.n376 163.367
R688 B.n374 B.n192 163.367
R689 B.n370 B.n368 163.367
R690 B.n366 B.n194 163.367
R691 B.n362 B.n360 163.367
R692 B.n358 B.n196 163.367
R693 B.n354 B.n352 163.367
R694 B.n350 B.n198 163.367
R695 B.n346 B.n344 163.367
R696 B.n342 B.n200 163.367
R697 B.n338 B.n336 163.367
R698 B.n334 B.n202 163.367
R699 B.n329 B.n327 163.367
R700 B.n325 B.n206 163.367
R701 B.n321 B.n319 163.367
R702 B.n317 B.n208 163.367
R703 B.n313 B.n311 163.367
R704 B.n309 B.n210 163.367
R705 B.n305 B.n303 163.367
R706 B.n301 B.n215 163.367
R707 B.n297 B.n295 163.367
R708 B.n293 B.n217 163.367
R709 B.n289 B.n287 163.367
R710 B.n285 B.n219 163.367
R711 B.n281 B.n279 163.367
R712 B.n277 B.n221 163.367
R713 B.n273 B.n271 163.367
R714 B.n269 B.n223 163.367
R715 B.n265 B.n263 163.367
R716 B.n261 B.n225 163.367
R717 B.n257 B.n255 163.367
R718 B.n253 B.n227 163.367
R719 B.n249 B.n247 163.367
R720 B.n245 B.n229 163.367
R721 B.n241 B.n239 163.367
R722 B.n237 B.n231 163.367
R723 B.n233 B.n180 163.367
R724 B.n411 B.n176 163.367
R725 B.n419 B.n176 163.367
R726 B.n419 B.n174 163.367
R727 B.n423 B.n174 163.367
R728 B.n423 B.n168 163.367
R729 B.n431 B.n168 163.367
R730 B.n431 B.n166 163.367
R731 B.n435 B.n166 163.367
R732 B.n435 B.n160 163.367
R733 B.n443 B.n160 163.367
R734 B.n443 B.n158 163.367
R735 B.n447 B.n158 163.367
R736 B.n447 B.n152 163.367
R737 B.n455 B.n152 163.367
R738 B.n455 B.n150 163.367
R739 B.n459 B.n150 163.367
R740 B.n459 B.n144 163.367
R741 B.n467 B.n144 163.367
R742 B.n467 B.n142 163.367
R743 B.n471 B.n142 163.367
R744 B.n471 B.n136 163.367
R745 B.n480 B.n136 163.367
R746 B.n480 B.n134 163.367
R747 B.n484 B.n134 163.367
R748 B.n484 B.n129 163.367
R749 B.n492 B.n129 163.367
R750 B.n492 B.n127 163.367
R751 B.n496 B.n127 163.367
R752 B.n496 B.n121 163.367
R753 B.n505 B.n121 163.367
R754 B.n505 B.n119 163.367
R755 B.n509 B.n119 163.367
R756 B.n509 B.n3 163.367
R757 B.n810 B.n3 163.367
R758 B.n806 B.n2 163.367
R759 B.n806 B.n805 163.367
R760 B.n805 B.n9 163.367
R761 B.n801 B.n9 163.367
R762 B.n801 B.n11 163.367
R763 B.n797 B.n11 163.367
R764 B.n797 B.n17 163.367
R765 B.n793 B.n17 163.367
R766 B.n793 B.n19 163.367
R767 B.n789 B.n19 163.367
R768 B.n789 B.n23 163.367
R769 B.n785 B.n23 163.367
R770 B.n785 B.n25 163.367
R771 B.n781 B.n25 163.367
R772 B.n781 B.n31 163.367
R773 B.n777 B.n31 163.367
R774 B.n777 B.n33 163.367
R775 B.n773 B.n33 163.367
R776 B.n773 B.n38 163.367
R777 B.n769 B.n38 163.367
R778 B.n769 B.n40 163.367
R779 B.n765 B.n40 163.367
R780 B.n765 B.n45 163.367
R781 B.n761 B.n45 163.367
R782 B.n761 B.n47 163.367
R783 B.n757 B.n47 163.367
R784 B.n757 B.n52 163.367
R785 B.n753 B.n52 163.367
R786 B.n753 B.n54 163.367
R787 B.n749 B.n54 163.367
R788 B.n749 B.n59 163.367
R789 B.n745 B.n59 163.367
R790 B.n745 B.n61 163.367
R791 B.n741 B.n61 163.367
R792 B.n412 B.n181 79.4395
R793 B.n742 B.n65 79.4395
R794 B.n736 B.n66 71.676
R795 B.n735 B.n734 71.676
R796 B.n728 B.n68 71.676
R797 B.n727 B.n726 71.676
R798 B.n720 B.n70 71.676
R799 B.n719 B.n718 71.676
R800 B.n712 B.n72 71.676
R801 B.n711 B.n710 71.676
R802 B.n704 B.n74 71.676
R803 B.n703 B.n702 71.676
R804 B.n696 B.n76 71.676
R805 B.n695 B.n694 71.676
R806 B.n688 B.n78 71.676
R807 B.n687 B.n686 71.676
R808 B.n680 B.n80 71.676
R809 B.n679 B.n678 71.676
R810 B.n672 B.n82 71.676
R811 B.n671 B.n670 71.676
R812 B.n664 B.n84 71.676
R813 B.n663 B.n662 71.676
R814 B.n655 B.n86 71.676
R815 B.n654 B.n653 71.676
R816 B.n647 B.n90 71.676
R817 B.n646 B.n645 71.676
R818 B.n639 B.n92 71.676
R819 B.n638 B.n96 71.676
R820 B.n634 B.n633 71.676
R821 B.n627 B.n98 71.676
R822 B.n626 B.n625 71.676
R823 B.n619 B.n100 71.676
R824 B.n618 B.n617 71.676
R825 B.n611 B.n102 71.676
R826 B.n610 B.n609 71.676
R827 B.n603 B.n104 71.676
R828 B.n602 B.n601 71.676
R829 B.n595 B.n106 71.676
R830 B.n594 B.n593 71.676
R831 B.n587 B.n108 71.676
R832 B.n586 B.n585 71.676
R833 B.n579 B.n110 71.676
R834 B.n578 B.n577 71.676
R835 B.n571 B.n112 71.676
R836 B.n570 B.n569 71.676
R837 B.n563 B.n114 71.676
R838 B.n562 B.n561 71.676
R839 B.n561 B.n560 71.676
R840 B.n564 B.n563 71.676
R841 B.n569 B.n568 71.676
R842 B.n572 B.n571 71.676
R843 B.n577 B.n576 71.676
R844 B.n580 B.n579 71.676
R845 B.n585 B.n584 71.676
R846 B.n588 B.n587 71.676
R847 B.n593 B.n592 71.676
R848 B.n596 B.n595 71.676
R849 B.n601 B.n600 71.676
R850 B.n604 B.n603 71.676
R851 B.n609 B.n608 71.676
R852 B.n612 B.n611 71.676
R853 B.n617 B.n616 71.676
R854 B.n620 B.n619 71.676
R855 B.n625 B.n624 71.676
R856 B.n628 B.n627 71.676
R857 B.n633 B.n632 71.676
R858 B.n635 B.n96 71.676
R859 B.n640 B.n639 71.676
R860 B.n645 B.n644 71.676
R861 B.n648 B.n647 71.676
R862 B.n653 B.n652 71.676
R863 B.n656 B.n655 71.676
R864 B.n662 B.n661 71.676
R865 B.n665 B.n664 71.676
R866 B.n670 B.n669 71.676
R867 B.n673 B.n672 71.676
R868 B.n678 B.n677 71.676
R869 B.n681 B.n680 71.676
R870 B.n686 B.n685 71.676
R871 B.n689 B.n688 71.676
R872 B.n694 B.n693 71.676
R873 B.n697 B.n696 71.676
R874 B.n702 B.n701 71.676
R875 B.n705 B.n704 71.676
R876 B.n710 B.n709 71.676
R877 B.n713 B.n712 71.676
R878 B.n718 B.n717 71.676
R879 B.n721 B.n720 71.676
R880 B.n726 B.n725 71.676
R881 B.n729 B.n728 71.676
R882 B.n734 B.n733 71.676
R883 B.n737 B.n736 71.676
R884 B.n406 B.n182 71.676
R885 B.n404 B.n184 71.676
R886 B.n400 B.n399 71.676
R887 B.n393 B.n186 71.676
R888 B.n392 B.n391 71.676
R889 B.n385 B.n188 71.676
R890 B.n384 B.n383 71.676
R891 B.n377 B.n190 71.676
R892 B.n376 B.n375 71.676
R893 B.n369 B.n192 71.676
R894 B.n368 B.n367 71.676
R895 B.n361 B.n194 71.676
R896 B.n360 B.n359 71.676
R897 B.n353 B.n196 71.676
R898 B.n352 B.n351 71.676
R899 B.n345 B.n198 71.676
R900 B.n344 B.n343 71.676
R901 B.n337 B.n200 71.676
R902 B.n336 B.n335 71.676
R903 B.n328 B.n202 71.676
R904 B.n327 B.n326 71.676
R905 B.n320 B.n206 71.676
R906 B.n319 B.n318 71.676
R907 B.n312 B.n208 71.676
R908 B.n311 B.n310 71.676
R909 B.n304 B.n210 71.676
R910 B.n303 B.n302 71.676
R911 B.n296 B.n215 71.676
R912 B.n295 B.n294 71.676
R913 B.n288 B.n217 71.676
R914 B.n287 B.n286 71.676
R915 B.n280 B.n219 71.676
R916 B.n279 B.n278 71.676
R917 B.n272 B.n221 71.676
R918 B.n271 B.n270 71.676
R919 B.n264 B.n223 71.676
R920 B.n263 B.n262 71.676
R921 B.n256 B.n225 71.676
R922 B.n255 B.n254 71.676
R923 B.n248 B.n227 71.676
R924 B.n247 B.n246 71.676
R925 B.n240 B.n229 71.676
R926 B.n239 B.n238 71.676
R927 B.n232 B.n231 71.676
R928 B.n407 B.n406 71.676
R929 B.n401 B.n184 71.676
R930 B.n399 B.n398 71.676
R931 B.n394 B.n393 71.676
R932 B.n391 B.n390 71.676
R933 B.n386 B.n385 71.676
R934 B.n383 B.n382 71.676
R935 B.n378 B.n377 71.676
R936 B.n375 B.n374 71.676
R937 B.n370 B.n369 71.676
R938 B.n367 B.n366 71.676
R939 B.n362 B.n361 71.676
R940 B.n359 B.n358 71.676
R941 B.n354 B.n353 71.676
R942 B.n351 B.n350 71.676
R943 B.n346 B.n345 71.676
R944 B.n343 B.n342 71.676
R945 B.n338 B.n337 71.676
R946 B.n335 B.n334 71.676
R947 B.n329 B.n328 71.676
R948 B.n326 B.n325 71.676
R949 B.n321 B.n320 71.676
R950 B.n318 B.n317 71.676
R951 B.n313 B.n312 71.676
R952 B.n310 B.n309 71.676
R953 B.n305 B.n304 71.676
R954 B.n302 B.n301 71.676
R955 B.n297 B.n296 71.676
R956 B.n294 B.n293 71.676
R957 B.n289 B.n288 71.676
R958 B.n286 B.n285 71.676
R959 B.n281 B.n280 71.676
R960 B.n278 B.n277 71.676
R961 B.n273 B.n272 71.676
R962 B.n270 B.n269 71.676
R963 B.n265 B.n264 71.676
R964 B.n262 B.n261 71.676
R965 B.n257 B.n256 71.676
R966 B.n254 B.n253 71.676
R967 B.n249 B.n248 71.676
R968 B.n246 B.n245 71.676
R969 B.n241 B.n240 71.676
R970 B.n238 B.n237 71.676
R971 B.n233 B.n232 71.676
R972 B.n811 B.n810 71.676
R973 B.n811 B.n2 71.676
R974 B.n659 B.n88 59.5399
R975 B.n95 B.n94 59.5399
R976 B.n213 B.n212 59.5399
R977 B.n331 B.n204 59.5399
R978 B.n412 B.n177 44.6439
R979 B.n418 B.n177 44.6439
R980 B.n418 B.n173 44.6439
R981 B.n424 B.n173 44.6439
R982 B.n424 B.n169 44.6439
R983 B.n430 B.n169 44.6439
R984 B.n436 B.n165 44.6439
R985 B.n436 B.n161 44.6439
R986 B.n442 B.n161 44.6439
R987 B.n442 B.n157 44.6439
R988 B.n448 B.n157 44.6439
R989 B.n448 B.n153 44.6439
R990 B.n454 B.n153 44.6439
R991 B.n454 B.n149 44.6439
R992 B.n460 B.n149 44.6439
R993 B.n466 B.n145 44.6439
R994 B.n466 B.n141 44.6439
R995 B.n472 B.n141 44.6439
R996 B.n472 B.n137 44.6439
R997 B.n479 B.n137 44.6439
R998 B.n479 B.n478 44.6439
R999 B.n485 B.n130 44.6439
R1000 B.n491 B.n130 44.6439
R1001 B.n491 B.n125 44.6439
R1002 B.n497 B.n125 44.6439
R1003 B.n497 B.n126 44.6439
R1004 B.n504 B.n118 44.6439
R1005 B.n510 B.n118 44.6439
R1006 B.n510 B.n4 44.6439
R1007 B.n809 B.n4 44.6439
R1008 B.n809 B.n808 44.6439
R1009 B.n808 B.n807 44.6439
R1010 B.n807 B.n8 44.6439
R1011 B.n12 B.n8 44.6439
R1012 B.n800 B.n12 44.6439
R1013 B.n799 B.n798 44.6439
R1014 B.n798 B.n16 44.6439
R1015 B.n792 B.n16 44.6439
R1016 B.n792 B.n791 44.6439
R1017 B.n791 B.n790 44.6439
R1018 B.n784 B.n26 44.6439
R1019 B.n784 B.n783 44.6439
R1020 B.n783 B.n782 44.6439
R1021 B.n782 B.n30 44.6439
R1022 B.n776 B.n30 44.6439
R1023 B.n776 B.n775 44.6439
R1024 B.n774 B.n37 44.6439
R1025 B.n768 B.n37 44.6439
R1026 B.n768 B.n767 44.6439
R1027 B.n767 B.n766 44.6439
R1028 B.n766 B.n44 44.6439
R1029 B.n760 B.n44 44.6439
R1030 B.n760 B.n759 44.6439
R1031 B.n759 B.n758 44.6439
R1032 B.n758 B.n51 44.6439
R1033 B.n752 B.n751 44.6439
R1034 B.n751 B.n750 44.6439
R1035 B.n750 B.n58 44.6439
R1036 B.n744 B.n58 44.6439
R1037 B.n744 B.n743 44.6439
R1038 B.n743 B.n742 44.6439
R1039 B.n485 B.t2 43.9874
R1040 B.n790 B.t3 43.9874
R1041 B.n88 B.n87 43.4429
R1042 B.n94 B.n93 43.4429
R1043 B.n212 B.n211 43.4429
R1044 B.n204 B.n203 43.4429
R1045 B.n410 B.n409 30.7517
R1046 B.n414 B.n179 30.7517
R1047 B.n559 B.n558 30.7517
R1048 B.n740 B.n739 30.7517
R1049 B.n430 B.t7 28.2309
R1050 B.n752 B.t14 28.2309
R1051 B.n126 B.t5 26.9178
R1052 B.t0 B.n799 26.9178
R1053 B.t4 B.n145 25.6048
R1054 B.n775 B.t1 25.6048
R1055 B.n460 B.t4 19.0396
R1056 B.t1 B.n774 19.0396
R1057 B B.n812 18.0485
R1058 B.n504 B.t5 17.7266
R1059 B.n800 B.t0 17.7266
R1060 B.t7 B.n165 16.4135
R1061 B.t14 B.n51 16.4135
R1062 B.n410 B.n175 10.6151
R1063 B.n420 B.n175 10.6151
R1064 B.n421 B.n420 10.6151
R1065 B.n422 B.n421 10.6151
R1066 B.n422 B.n167 10.6151
R1067 B.n432 B.n167 10.6151
R1068 B.n433 B.n432 10.6151
R1069 B.n434 B.n433 10.6151
R1070 B.n434 B.n159 10.6151
R1071 B.n444 B.n159 10.6151
R1072 B.n445 B.n444 10.6151
R1073 B.n446 B.n445 10.6151
R1074 B.n446 B.n151 10.6151
R1075 B.n456 B.n151 10.6151
R1076 B.n457 B.n456 10.6151
R1077 B.n458 B.n457 10.6151
R1078 B.n458 B.n143 10.6151
R1079 B.n468 B.n143 10.6151
R1080 B.n469 B.n468 10.6151
R1081 B.n470 B.n469 10.6151
R1082 B.n470 B.n135 10.6151
R1083 B.n481 B.n135 10.6151
R1084 B.n482 B.n481 10.6151
R1085 B.n483 B.n482 10.6151
R1086 B.n483 B.n128 10.6151
R1087 B.n493 B.n128 10.6151
R1088 B.n494 B.n493 10.6151
R1089 B.n495 B.n494 10.6151
R1090 B.n495 B.n120 10.6151
R1091 B.n506 B.n120 10.6151
R1092 B.n507 B.n506 10.6151
R1093 B.n508 B.n507 10.6151
R1094 B.n508 B.n0 10.6151
R1095 B.n409 B.n408 10.6151
R1096 B.n408 B.n183 10.6151
R1097 B.n403 B.n183 10.6151
R1098 B.n403 B.n402 10.6151
R1099 B.n402 B.n185 10.6151
R1100 B.n397 B.n185 10.6151
R1101 B.n397 B.n396 10.6151
R1102 B.n396 B.n395 10.6151
R1103 B.n395 B.n187 10.6151
R1104 B.n389 B.n187 10.6151
R1105 B.n389 B.n388 10.6151
R1106 B.n388 B.n387 10.6151
R1107 B.n387 B.n189 10.6151
R1108 B.n381 B.n189 10.6151
R1109 B.n381 B.n380 10.6151
R1110 B.n380 B.n379 10.6151
R1111 B.n379 B.n191 10.6151
R1112 B.n373 B.n191 10.6151
R1113 B.n373 B.n372 10.6151
R1114 B.n372 B.n371 10.6151
R1115 B.n371 B.n193 10.6151
R1116 B.n365 B.n193 10.6151
R1117 B.n365 B.n364 10.6151
R1118 B.n364 B.n363 10.6151
R1119 B.n363 B.n195 10.6151
R1120 B.n357 B.n195 10.6151
R1121 B.n357 B.n356 10.6151
R1122 B.n356 B.n355 10.6151
R1123 B.n355 B.n197 10.6151
R1124 B.n349 B.n197 10.6151
R1125 B.n349 B.n348 10.6151
R1126 B.n348 B.n347 10.6151
R1127 B.n347 B.n199 10.6151
R1128 B.n341 B.n199 10.6151
R1129 B.n341 B.n340 10.6151
R1130 B.n340 B.n339 10.6151
R1131 B.n339 B.n201 10.6151
R1132 B.n333 B.n201 10.6151
R1133 B.n333 B.n332 10.6151
R1134 B.n330 B.n205 10.6151
R1135 B.n324 B.n205 10.6151
R1136 B.n324 B.n323 10.6151
R1137 B.n323 B.n322 10.6151
R1138 B.n322 B.n207 10.6151
R1139 B.n316 B.n207 10.6151
R1140 B.n316 B.n315 10.6151
R1141 B.n315 B.n314 10.6151
R1142 B.n314 B.n209 10.6151
R1143 B.n308 B.n307 10.6151
R1144 B.n307 B.n306 10.6151
R1145 B.n306 B.n214 10.6151
R1146 B.n300 B.n214 10.6151
R1147 B.n300 B.n299 10.6151
R1148 B.n299 B.n298 10.6151
R1149 B.n298 B.n216 10.6151
R1150 B.n292 B.n216 10.6151
R1151 B.n292 B.n291 10.6151
R1152 B.n291 B.n290 10.6151
R1153 B.n290 B.n218 10.6151
R1154 B.n284 B.n218 10.6151
R1155 B.n284 B.n283 10.6151
R1156 B.n283 B.n282 10.6151
R1157 B.n282 B.n220 10.6151
R1158 B.n276 B.n220 10.6151
R1159 B.n276 B.n275 10.6151
R1160 B.n275 B.n274 10.6151
R1161 B.n274 B.n222 10.6151
R1162 B.n268 B.n222 10.6151
R1163 B.n268 B.n267 10.6151
R1164 B.n267 B.n266 10.6151
R1165 B.n266 B.n224 10.6151
R1166 B.n260 B.n224 10.6151
R1167 B.n260 B.n259 10.6151
R1168 B.n259 B.n258 10.6151
R1169 B.n258 B.n226 10.6151
R1170 B.n252 B.n226 10.6151
R1171 B.n252 B.n251 10.6151
R1172 B.n251 B.n250 10.6151
R1173 B.n250 B.n228 10.6151
R1174 B.n244 B.n228 10.6151
R1175 B.n244 B.n243 10.6151
R1176 B.n243 B.n242 10.6151
R1177 B.n242 B.n230 10.6151
R1178 B.n236 B.n230 10.6151
R1179 B.n236 B.n235 10.6151
R1180 B.n235 B.n234 10.6151
R1181 B.n234 B.n179 10.6151
R1182 B.n415 B.n414 10.6151
R1183 B.n416 B.n415 10.6151
R1184 B.n416 B.n171 10.6151
R1185 B.n426 B.n171 10.6151
R1186 B.n427 B.n426 10.6151
R1187 B.n428 B.n427 10.6151
R1188 B.n428 B.n163 10.6151
R1189 B.n438 B.n163 10.6151
R1190 B.n439 B.n438 10.6151
R1191 B.n440 B.n439 10.6151
R1192 B.n440 B.n155 10.6151
R1193 B.n450 B.n155 10.6151
R1194 B.n451 B.n450 10.6151
R1195 B.n452 B.n451 10.6151
R1196 B.n452 B.n147 10.6151
R1197 B.n462 B.n147 10.6151
R1198 B.n463 B.n462 10.6151
R1199 B.n464 B.n463 10.6151
R1200 B.n464 B.n139 10.6151
R1201 B.n474 B.n139 10.6151
R1202 B.n475 B.n474 10.6151
R1203 B.n476 B.n475 10.6151
R1204 B.n476 B.n132 10.6151
R1205 B.n487 B.n132 10.6151
R1206 B.n488 B.n487 10.6151
R1207 B.n489 B.n488 10.6151
R1208 B.n489 B.n123 10.6151
R1209 B.n499 B.n123 10.6151
R1210 B.n500 B.n499 10.6151
R1211 B.n502 B.n500 10.6151
R1212 B.n502 B.n501 10.6151
R1213 B.n501 B.n116 10.6151
R1214 B.n513 B.n116 10.6151
R1215 B.n514 B.n513 10.6151
R1216 B.n515 B.n514 10.6151
R1217 B.n516 B.n515 10.6151
R1218 B.n517 B.n516 10.6151
R1219 B.n520 B.n517 10.6151
R1220 B.n521 B.n520 10.6151
R1221 B.n522 B.n521 10.6151
R1222 B.n523 B.n522 10.6151
R1223 B.n525 B.n523 10.6151
R1224 B.n526 B.n525 10.6151
R1225 B.n527 B.n526 10.6151
R1226 B.n528 B.n527 10.6151
R1227 B.n530 B.n528 10.6151
R1228 B.n531 B.n530 10.6151
R1229 B.n532 B.n531 10.6151
R1230 B.n533 B.n532 10.6151
R1231 B.n535 B.n533 10.6151
R1232 B.n536 B.n535 10.6151
R1233 B.n537 B.n536 10.6151
R1234 B.n538 B.n537 10.6151
R1235 B.n540 B.n538 10.6151
R1236 B.n541 B.n540 10.6151
R1237 B.n542 B.n541 10.6151
R1238 B.n543 B.n542 10.6151
R1239 B.n545 B.n543 10.6151
R1240 B.n546 B.n545 10.6151
R1241 B.n547 B.n546 10.6151
R1242 B.n548 B.n547 10.6151
R1243 B.n550 B.n548 10.6151
R1244 B.n551 B.n550 10.6151
R1245 B.n552 B.n551 10.6151
R1246 B.n553 B.n552 10.6151
R1247 B.n555 B.n553 10.6151
R1248 B.n556 B.n555 10.6151
R1249 B.n557 B.n556 10.6151
R1250 B.n558 B.n557 10.6151
R1251 B.n804 B.n1 10.6151
R1252 B.n804 B.n803 10.6151
R1253 B.n803 B.n802 10.6151
R1254 B.n802 B.n10 10.6151
R1255 B.n796 B.n10 10.6151
R1256 B.n796 B.n795 10.6151
R1257 B.n795 B.n794 10.6151
R1258 B.n794 B.n18 10.6151
R1259 B.n788 B.n18 10.6151
R1260 B.n788 B.n787 10.6151
R1261 B.n787 B.n786 10.6151
R1262 B.n786 B.n24 10.6151
R1263 B.n780 B.n24 10.6151
R1264 B.n780 B.n779 10.6151
R1265 B.n779 B.n778 10.6151
R1266 B.n778 B.n32 10.6151
R1267 B.n772 B.n32 10.6151
R1268 B.n772 B.n771 10.6151
R1269 B.n771 B.n770 10.6151
R1270 B.n770 B.n39 10.6151
R1271 B.n764 B.n39 10.6151
R1272 B.n764 B.n763 10.6151
R1273 B.n763 B.n762 10.6151
R1274 B.n762 B.n46 10.6151
R1275 B.n756 B.n46 10.6151
R1276 B.n756 B.n755 10.6151
R1277 B.n755 B.n754 10.6151
R1278 B.n754 B.n53 10.6151
R1279 B.n748 B.n53 10.6151
R1280 B.n748 B.n747 10.6151
R1281 B.n747 B.n746 10.6151
R1282 B.n746 B.n60 10.6151
R1283 B.n740 B.n60 10.6151
R1284 B.n739 B.n738 10.6151
R1285 B.n738 B.n67 10.6151
R1286 B.n732 B.n67 10.6151
R1287 B.n732 B.n731 10.6151
R1288 B.n731 B.n730 10.6151
R1289 B.n730 B.n69 10.6151
R1290 B.n724 B.n69 10.6151
R1291 B.n724 B.n723 10.6151
R1292 B.n723 B.n722 10.6151
R1293 B.n722 B.n71 10.6151
R1294 B.n716 B.n71 10.6151
R1295 B.n716 B.n715 10.6151
R1296 B.n715 B.n714 10.6151
R1297 B.n714 B.n73 10.6151
R1298 B.n708 B.n73 10.6151
R1299 B.n708 B.n707 10.6151
R1300 B.n707 B.n706 10.6151
R1301 B.n706 B.n75 10.6151
R1302 B.n700 B.n75 10.6151
R1303 B.n700 B.n699 10.6151
R1304 B.n699 B.n698 10.6151
R1305 B.n698 B.n77 10.6151
R1306 B.n692 B.n77 10.6151
R1307 B.n692 B.n691 10.6151
R1308 B.n691 B.n690 10.6151
R1309 B.n690 B.n79 10.6151
R1310 B.n684 B.n79 10.6151
R1311 B.n684 B.n683 10.6151
R1312 B.n683 B.n682 10.6151
R1313 B.n682 B.n81 10.6151
R1314 B.n676 B.n81 10.6151
R1315 B.n676 B.n675 10.6151
R1316 B.n675 B.n674 10.6151
R1317 B.n674 B.n83 10.6151
R1318 B.n668 B.n83 10.6151
R1319 B.n668 B.n667 10.6151
R1320 B.n667 B.n666 10.6151
R1321 B.n666 B.n85 10.6151
R1322 B.n660 B.n85 10.6151
R1323 B.n658 B.n657 10.6151
R1324 B.n657 B.n89 10.6151
R1325 B.n651 B.n89 10.6151
R1326 B.n651 B.n650 10.6151
R1327 B.n650 B.n649 10.6151
R1328 B.n649 B.n91 10.6151
R1329 B.n643 B.n91 10.6151
R1330 B.n643 B.n642 10.6151
R1331 B.n642 B.n641 10.6151
R1332 B.n637 B.n636 10.6151
R1333 B.n636 B.n97 10.6151
R1334 B.n631 B.n97 10.6151
R1335 B.n631 B.n630 10.6151
R1336 B.n630 B.n629 10.6151
R1337 B.n629 B.n99 10.6151
R1338 B.n623 B.n99 10.6151
R1339 B.n623 B.n622 10.6151
R1340 B.n622 B.n621 10.6151
R1341 B.n621 B.n101 10.6151
R1342 B.n615 B.n101 10.6151
R1343 B.n615 B.n614 10.6151
R1344 B.n614 B.n613 10.6151
R1345 B.n613 B.n103 10.6151
R1346 B.n607 B.n103 10.6151
R1347 B.n607 B.n606 10.6151
R1348 B.n606 B.n605 10.6151
R1349 B.n605 B.n105 10.6151
R1350 B.n599 B.n105 10.6151
R1351 B.n599 B.n598 10.6151
R1352 B.n598 B.n597 10.6151
R1353 B.n597 B.n107 10.6151
R1354 B.n591 B.n107 10.6151
R1355 B.n591 B.n590 10.6151
R1356 B.n590 B.n589 10.6151
R1357 B.n589 B.n109 10.6151
R1358 B.n583 B.n109 10.6151
R1359 B.n583 B.n582 10.6151
R1360 B.n582 B.n581 10.6151
R1361 B.n581 B.n111 10.6151
R1362 B.n575 B.n111 10.6151
R1363 B.n575 B.n574 10.6151
R1364 B.n574 B.n573 10.6151
R1365 B.n573 B.n113 10.6151
R1366 B.n567 B.n113 10.6151
R1367 B.n567 B.n566 10.6151
R1368 B.n566 B.n565 10.6151
R1369 B.n565 B.n115 10.6151
R1370 B.n559 B.n115 10.6151
R1371 B.n332 B.n331 9.36635
R1372 B.n308 B.n213 9.36635
R1373 B.n660 B.n659 9.36635
R1374 B.n637 B.n95 9.36635
R1375 B.n812 B.n0 8.11757
R1376 B.n812 B.n1 8.11757
R1377 B.n331 B.n330 1.24928
R1378 B.n213 B.n209 1.24928
R1379 B.n659 B.n658 1.24928
R1380 B.n641 B.n95 1.24928
R1381 B.n478 B.t2 0.65702
R1382 B.n26 B.t3 0.65702
R1383 VP.n6 VP.t0 176.095
R1384 VP.n9 VP.n8 161.3
R1385 VP.n10 VP.n5 161.3
R1386 VP.n12 VP.n11 161.3
R1387 VP.n13 VP.n4 161.3
R1388 VP.n30 VP.n0 161.3
R1389 VP.n29 VP.n28 161.3
R1390 VP.n27 VP.n1 161.3
R1391 VP.n26 VP.n25 161.3
R1392 VP.n23 VP.n2 161.3
R1393 VP.n22 VP.n21 161.3
R1394 VP.n20 VP.n3 161.3
R1395 VP.n19 VP.n18 161.3
R1396 VP.n17 VP.t1 144.852
R1397 VP.n24 VP.t5 144.852
R1398 VP.n31 VP.t4 144.852
R1399 VP.n14 VP.t3 144.852
R1400 VP.n7 VP.t2 144.852
R1401 VP.n17 VP.n16 86.7496
R1402 VP.n32 VP.n31 86.7496
R1403 VP.n15 VP.n14 86.7496
R1404 VP.n7 VP.n6 57.7381
R1405 VP.n22 VP.n3 53.0692
R1406 VP.n29 VP.n1 53.0692
R1407 VP.n12 VP.n5 53.0692
R1408 VP.n16 VP.n15 45.6435
R1409 VP.n18 VP.n3 27.752
R1410 VP.n30 VP.n29 27.752
R1411 VP.n13 VP.n12 27.752
R1412 VP.n23 VP.n22 24.3439
R1413 VP.n25 VP.n1 24.3439
R1414 VP.n8 VP.n5 24.3439
R1415 VP.n18 VP.n17 23.8571
R1416 VP.n31 VP.n30 23.8571
R1417 VP.n14 VP.n13 23.8571
R1418 VP.n9 VP.n6 12.7265
R1419 VP.n24 VP.n23 12.1722
R1420 VP.n25 VP.n24 12.1722
R1421 VP.n8 VP.n7 12.1722
R1422 VP.n15 VP.n4 0.278398
R1423 VP.n19 VP.n16 0.278398
R1424 VP.n32 VP.n0 0.278398
R1425 VP.n10 VP.n9 0.189894
R1426 VP.n11 VP.n10 0.189894
R1427 VP.n11 VP.n4 0.189894
R1428 VP.n20 VP.n19 0.189894
R1429 VP.n21 VP.n20 0.189894
R1430 VP.n21 VP.n2 0.189894
R1431 VP.n26 VP.n2 0.189894
R1432 VP.n27 VP.n26 0.189894
R1433 VP.n28 VP.n27 0.189894
R1434 VP.n28 VP.n0 0.189894
R1435 VP VP.n32 0.153422
R1436 VTAIL.n250 VTAIL.n194 289.615
R1437 VTAIL.n58 VTAIL.n2 289.615
R1438 VTAIL.n188 VTAIL.n132 289.615
R1439 VTAIL.n124 VTAIL.n68 289.615
R1440 VTAIL.n215 VTAIL.n214 185
R1441 VTAIL.n217 VTAIL.n216 185
R1442 VTAIL.n210 VTAIL.n209 185
R1443 VTAIL.n223 VTAIL.n222 185
R1444 VTAIL.n225 VTAIL.n224 185
R1445 VTAIL.n206 VTAIL.n205 185
R1446 VTAIL.n232 VTAIL.n231 185
R1447 VTAIL.n233 VTAIL.n204 185
R1448 VTAIL.n235 VTAIL.n234 185
R1449 VTAIL.n202 VTAIL.n201 185
R1450 VTAIL.n241 VTAIL.n240 185
R1451 VTAIL.n243 VTAIL.n242 185
R1452 VTAIL.n198 VTAIL.n197 185
R1453 VTAIL.n249 VTAIL.n248 185
R1454 VTAIL.n251 VTAIL.n250 185
R1455 VTAIL.n23 VTAIL.n22 185
R1456 VTAIL.n25 VTAIL.n24 185
R1457 VTAIL.n18 VTAIL.n17 185
R1458 VTAIL.n31 VTAIL.n30 185
R1459 VTAIL.n33 VTAIL.n32 185
R1460 VTAIL.n14 VTAIL.n13 185
R1461 VTAIL.n40 VTAIL.n39 185
R1462 VTAIL.n41 VTAIL.n12 185
R1463 VTAIL.n43 VTAIL.n42 185
R1464 VTAIL.n10 VTAIL.n9 185
R1465 VTAIL.n49 VTAIL.n48 185
R1466 VTAIL.n51 VTAIL.n50 185
R1467 VTAIL.n6 VTAIL.n5 185
R1468 VTAIL.n57 VTAIL.n56 185
R1469 VTAIL.n59 VTAIL.n58 185
R1470 VTAIL.n189 VTAIL.n188 185
R1471 VTAIL.n187 VTAIL.n186 185
R1472 VTAIL.n136 VTAIL.n135 185
R1473 VTAIL.n181 VTAIL.n180 185
R1474 VTAIL.n179 VTAIL.n178 185
R1475 VTAIL.n140 VTAIL.n139 185
R1476 VTAIL.n144 VTAIL.n142 185
R1477 VTAIL.n173 VTAIL.n172 185
R1478 VTAIL.n171 VTAIL.n170 185
R1479 VTAIL.n146 VTAIL.n145 185
R1480 VTAIL.n165 VTAIL.n164 185
R1481 VTAIL.n163 VTAIL.n162 185
R1482 VTAIL.n150 VTAIL.n149 185
R1483 VTAIL.n157 VTAIL.n156 185
R1484 VTAIL.n155 VTAIL.n154 185
R1485 VTAIL.n125 VTAIL.n124 185
R1486 VTAIL.n123 VTAIL.n122 185
R1487 VTAIL.n72 VTAIL.n71 185
R1488 VTAIL.n117 VTAIL.n116 185
R1489 VTAIL.n115 VTAIL.n114 185
R1490 VTAIL.n76 VTAIL.n75 185
R1491 VTAIL.n80 VTAIL.n78 185
R1492 VTAIL.n109 VTAIL.n108 185
R1493 VTAIL.n107 VTAIL.n106 185
R1494 VTAIL.n82 VTAIL.n81 185
R1495 VTAIL.n101 VTAIL.n100 185
R1496 VTAIL.n99 VTAIL.n98 185
R1497 VTAIL.n86 VTAIL.n85 185
R1498 VTAIL.n93 VTAIL.n92 185
R1499 VTAIL.n91 VTAIL.n90 185
R1500 VTAIL.n213 VTAIL.t1 149.524
R1501 VTAIL.n21 VTAIL.t6 149.524
R1502 VTAIL.n153 VTAIL.t7 149.524
R1503 VTAIL.n89 VTAIL.t11 149.524
R1504 VTAIL.n216 VTAIL.n215 104.615
R1505 VTAIL.n216 VTAIL.n209 104.615
R1506 VTAIL.n223 VTAIL.n209 104.615
R1507 VTAIL.n224 VTAIL.n223 104.615
R1508 VTAIL.n224 VTAIL.n205 104.615
R1509 VTAIL.n232 VTAIL.n205 104.615
R1510 VTAIL.n233 VTAIL.n232 104.615
R1511 VTAIL.n234 VTAIL.n233 104.615
R1512 VTAIL.n234 VTAIL.n201 104.615
R1513 VTAIL.n241 VTAIL.n201 104.615
R1514 VTAIL.n242 VTAIL.n241 104.615
R1515 VTAIL.n242 VTAIL.n197 104.615
R1516 VTAIL.n249 VTAIL.n197 104.615
R1517 VTAIL.n250 VTAIL.n249 104.615
R1518 VTAIL.n24 VTAIL.n23 104.615
R1519 VTAIL.n24 VTAIL.n17 104.615
R1520 VTAIL.n31 VTAIL.n17 104.615
R1521 VTAIL.n32 VTAIL.n31 104.615
R1522 VTAIL.n32 VTAIL.n13 104.615
R1523 VTAIL.n40 VTAIL.n13 104.615
R1524 VTAIL.n41 VTAIL.n40 104.615
R1525 VTAIL.n42 VTAIL.n41 104.615
R1526 VTAIL.n42 VTAIL.n9 104.615
R1527 VTAIL.n49 VTAIL.n9 104.615
R1528 VTAIL.n50 VTAIL.n49 104.615
R1529 VTAIL.n50 VTAIL.n5 104.615
R1530 VTAIL.n57 VTAIL.n5 104.615
R1531 VTAIL.n58 VTAIL.n57 104.615
R1532 VTAIL.n188 VTAIL.n187 104.615
R1533 VTAIL.n187 VTAIL.n135 104.615
R1534 VTAIL.n180 VTAIL.n135 104.615
R1535 VTAIL.n180 VTAIL.n179 104.615
R1536 VTAIL.n179 VTAIL.n139 104.615
R1537 VTAIL.n144 VTAIL.n139 104.615
R1538 VTAIL.n172 VTAIL.n144 104.615
R1539 VTAIL.n172 VTAIL.n171 104.615
R1540 VTAIL.n171 VTAIL.n145 104.615
R1541 VTAIL.n164 VTAIL.n145 104.615
R1542 VTAIL.n164 VTAIL.n163 104.615
R1543 VTAIL.n163 VTAIL.n149 104.615
R1544 VTAIL.n156 VTAIL.n149 104.615
R1545 VTAIL.n156 VTAIL.n155 104.615
R1546 VTAIL.n124 VTAIL.n123 104.615
R1547 VTAIL.n123 VTAIL.n71 104.615
R1548 VTAIL.n116 VTAIL.n71 104.615
R1549 VTAIL.n116 VTAIL.n115 104.615
R1550 VTAIL.n115 VTAIL.n75 104.615
R1551 VTAIL.n80 VTAIL.n75 104.615
R1552 VTAIL.n108 VTAIL.n80 104.615
R1553 VTAIL.n108 VTAIL.n107 104.615
R1554 VTAIL.n107 VTAIL.n81 104.615
R1555 VTAIL.n100 VTAIL.n81 104.615
R1556 VTAIL.n100 VTAIL.n99 104.615
R1557 VTAIL.n99 VTAIL.n85 104.615
R1558 VTAIL.n92 VTAIL.n85 104.615
R1559 VTAIL.n92 VTAIL.n91 104.615
R1560 VTAIL.n215 VTAIL.t1 52.3082
R1561 VTAIL.n23 VTAIL.t6 52.3082
R1562 VTAIL.n155 VTAIL.t7 52.3082
R1563 VTAIL.n91 VTAIL.t11 52.3082
R1564 VTAIL.n131 VTAIL.n130 46.9626
R1565 VTAIL.n67 VTAIL.n66 46.9626
R1566 VTAIL.n1 VTAIL.n0 46.9625
R1567 VTAIL.n65 VTAIL.n64 46.9625
R1568 VTAIL.n255 VTAIL.n254 33.7369
R1569 VTAIL.n63 VTAIL.n62 33.7369
R1570 VTAIL.n193 VTAIL.n192 33.7369
R1571 VTAIL.n129 VTAIL.n128 33.7369
R1572 VTAIL.n67 VTAIL.n65 26.1255
R1573 VTAIL.n255 VTAIL.n193 24.1945
R1574 VTAIL.n235 VTAIL.n202 13.1884
R1575 VTAIL.n43 VTAIL.n10 13.1884
R1576 VTAIL.n142 VTAIL.n140 13.1884
R1577 VTAIL.n78 VTAIL.n76 13.1884
R1578 VTAIL.n236 VTAIL.n204 12.8005
R1579 VTAIL.n240 VTAIL.n239 12.8005
R1580 VTAIL.n44 VTAIL.n12 12.8005
R1581 VTAIL.n48 VTAIL.n47 12.8005
R1582 VTAIL.n178 VTAIL.n177 12.8005
R1583 VTAIL.n174 VTAIL.n173 12.8005
R1584 VTAIL.n114 VTAIL.n113 12.8005
R1585 VTAIL.n110 VTAIL.n109 12.8005
R1586 VTAIL.n231 VTAIL.n230 12.0247
R1587 VTAIL.n243 VTAIL.n200 12.0247
R1588 VTAIL.n39 VTAIL.n38 12.0247
R1589 VTAIL.n51 VTAIL.n8 12.0247
R1590 VTAIL.n181 VTAIL.n138 12.0247
R1591 VTAIL.n170 VTAIL.n143 12.0247
R1592 VTAIL.n117 VTAIL.n74 12.0247
R1593 VTAIL.n106 VTAIL.n79 12.0247
R1594 VTAIL.n229 VTAIL.n206 11.249
R1595 VTAIL.n244 VTAIL.n198 11.249
R1596 VTAIL.n37 VTAIL.n14 11.249
R1597 VTAIL.n52 VTAIL.n6 11.249
R1598 VTAIL.n182 VTAIL.n136 11.249
R1599 VTAIL.n169 VTAIL.n146 11.249
R1600 VTAIL.n118 VTAIL.n72 11.249
R1601 VTAIL.n105 VTAIL.n82 11.249
R1602 VTAIL.n226 VTAIL.n225 10.4732
R1603 VTAIL.n248 VTAIL.n247 10.4732
R1604 VTAIL.n34 VTAIL.n33 10.4732
R1605 VTAIL.n56 VTAIL.n55 10.4732
R1606 VTAIL.n186 VTAIL.n185 10.4732
R1607 VTAIL.n166 VTAIL.n165 10.4732
R1608 VTAIL.n122 VTAIL.n121 10.4732
R1609 VTAIL.n102 VTAIL.n101 10.4732
R1610 VTAIL.n214 VTAIL.n213 10.2747
R1611 VTAIL.n22 VTAIL.n21 10.2747
R1612 VTAIL.n154 VTAIL.n153 10.2747
R1613 VTAIL.n90 VTAIL.n89 10.2747
R1614 VTAIL.n222 VTAIL.n208 9.69747
R1615 VTAIL.n251 VTAIL.n196 9.69747
R1616 VTAIL.n30 VTAIL.n16 9.69747
R1617 VTAIL.n59 VTAIL.n4 9.69747
R1618 VTAIL.n189 VTAIL.n134 9.69747
R1619 VTAIL.n162 VTAIL.n148 9.69747
R1620 VTAIL.n125 VTAIL.n70 9.69747
R1621 VTAIL.n98 VTAIL.n84 9.69747
R1622 VTAIL.n254 VTAIL.n253 9.45567
R1623 VTAIL.n62 VTAIL.n61 9.45567
R1624 VTAIL.n192 VTAIL.n191 9.45567
R1625 VTAIL.n128 VTAIL.n127 9.45567
R1626 VTAIL.n253 VTAIL.n252 9.3005
R1627 VTAIL.n196 VTAIL.n195 9.3005
R1628 VTAIL.n247 VTAIL.n246 9.3005
R1629 VTAIL.n245 VTAIL.n244 9.3005
R1630 VTAIL.n200 VTAIL.n199 9.3005
R1631 VTAIL.n239 VTAIL.n238 9.3005
R1632 VTAIL.n212 VTAIL.n211 9.3005
R1633 VTAIL.n219 VTAIL.n218 9.3005
R1634 VTAIL.n221 VTAIL.n220 9.3005
R1635 VTAIL.n208 VTAIL.n207 9.3005
R1636 VTAIL.n227 VTAIL.n226 9.3005
R1637 VTAIL.n229 VTAIL.n228 9.3005
R1638 VTAIL.n230 VTAIL.n203 9.3005
R1639 VTAIL.n237 VTAIL.n236 9.3005
R1640 VTAIL.n61 VTAIL.n60 9.3005
R1641 VTAIL.n4 VTAIL.n3 9.3005
R1642 VTAIL.n55 VTAIL.n54 9.3005
R1643 VTAIL.n53 VTAIL.n52 9.3005
R1644 VTAIL.n8 VTAIL.n7 9.3005
R1645 VTAIL.n47 VTAIL.n46 9.3005
R1646 VTAIL.n20 VTAIL.n19 9.3005
R1647 VTAIL.n27 VTAIL.n26 9.3005
R1648 VTAIL.n29 VTAIL.n28 9.3005
R1649 VTAIL.n16 VTAIL.n15 9.3005
R1650 VTAIL.n35 VTAIL.n34 9.3005
R1651 VTAIL.n37 VTAIL.n36 9.3005
R1652 VTAIL.n38 VTAIL.n11 9.3005
R1653 VTAIL.n45 VTAIL.n44 9.3005
R1654 VTAIL.n152 VTAIL.n151 9.3005
R1655 VTAIL.n159 VTAIL.n158 9.3005
R1656 VTAIL.n161 VTAIL.n160 9.3005
R1657 VTAIL.n148 VTAIL.n147 9.3005
R1658 VTAIL.n167 VTAIL.n166 9.3005
R1659 VTAIL.n169 VTAIL.n168 9.3005
R1660 VTAIL.n143 VTAIL.n141 9.3005
R1661 VTAIL.n175 VTAIL.n174 9.3005
R1662 VTAIL.n191 VTAIL.n190 9.3005
R1663 VTAIL.n134 VTAIL.n133 9.3005
R1664 VTAIL.n185 VTAIL.n184 9.3005
R1665 VTAIL.n183 VTAIL.n182 9.3005
R1666 VTAIL.n138 VTAIL.n137 9.3005
R1667 VTAIL.n177 VTAIL.n176 9.3005
R1668 VTAIL.n88 VTAIL.n87 9.3005
R1669 VTAIL.n95 VTAIL.n94 9.3005
R1670 VTAIL.n97 VTAIL.n96 9.3005
R1671 VTAIL.n84 VTAIL.n83 9.3005
R1672 VTAIL.n103 VTAIL.n102 9.3005
R1673 VTAIL.n105 VTAIL.n104 9.3005
R1674 VTAIL.n79 VTAIL.n77 9.3005
R1675 VTAIL.n111 VTAIL.n110 9.3005
R1676 VTAIL.n127 VTAIL.n126 9.3005
R1677 VTAIL.n70 VTAIL.n69 9.3005
R1678 VTAIL.n121 VTAIL.n120 9.3005
R1679 VTAIL.n119 VTAIL.n118 9.3005
R1680 VTAIL.n74 VTAIL.n73 9.3005
R1681 VTAIL.n113 VTAIL.n112 9.3005
R1682 VTAIL.n221 VTAIL.n210 8.92171
R1683 VTAIL.n252 VTAIL.n194 8.92171
R1684 VTAIL.n29 VTAIL.n18 8.92171
R1685 VTAIL.n60 VTAIL.n2 8.92171
R1686 VTAIL.n190 VTAIL.n132 8.92171
R1687 VTAIL.n161 VTAIL.n150 8.92171
R1688 VTAIL.n126 VTAIL.n68 8.92171
R1689 VTAIL.n97 VTAIL.n86 8.92171
R1690 VTAIL.n218 VTAIL.n217 8.14595
R1691 VTAIL.n26 VTAIL.n25 8.14595
R1692 VTAIL.n158 VTAIL.n157 8.14595
R1693 VTAIL.n94 VTAIL.n93 8.14595
R1694 VTAIL.n214 VTAIL.n212 7.3702
R1695 VTAIL.n22 VTAIL.n20 7.3702
R1696 VTAIL.n154 VTAIL.n152 7.3702
R1697 VTAIL.n90 VTAIL.n88 7.3702
R1698 VTAIL.n217 VTAIL.n212 5.81868
R1699 VTAIL.n25 VTAIL.n20 5.81868
R1700 VTAIL.n157 VTAIL.n152 5.81868
R1701 VTAIL.n93 VTAIL.n88 5.81868
R1702 VTAIL.n218 VTAIL.n210 5.04292
R1703 VTAIL.n254 VTAIL.n194 5.04292
R1704 VTAIL.n26 VTAIL.n18 5.04292
R1705 VTAIL.n62 VTAIL.n2 5.04292
R1706 VTAIL.n192 VTAIL.n132 5.04292
R1707 VTAIL.n158 VTAIL.n150 5.04292
R1708 VTAIL.n128 VTAIL.n68 5.04292
R1709 VTAIL.n94 VTAIL.n86 5.04292
R1710 VTAIL.n222 VTAIL.n221 4.26717
R1711 VTAIL.n252 VTAIL.n251 4.26717
R1712 VTAIL.n30 VTAIL.n29 4.26717
R1713 VTAIL.n60 VTAIL.n59 4.26717
R1714 VTAIL.n190 VTAIL.n189 4.26717
R1715 VTAIL.n162 VTAIL.n161 4.26717
R1716 VTAIL.n126 VTAIL.n125 4.26717
R1717 VTAIL.n98 VTAIL.n97 4.26717
R1718 VTAIL.n225 VTAIL.n208 3.49141
R1719 VTAIL.n248 VTAIL.n196 3.49141
R1720 VTAIL.n33 VTAIL.n16 3.49141
R1721 VTAIL.n56 VTAIL.n4 3.49141
R1722 VTAIL.n186 VTAIL.n134 3.49141
R1723 VTAIL.n165 VTAIL.n148 3.49141
R1724 VTAIL.n122 VTAIL.n70 3.49141
R1725 VTAIL.n101 VTAIL.n84 3.49141
R1726 VTAIL.n213 VTAIL.n211 2.84303
R1727 VTAIL.n21 VTAIL.n19 2.84303
R1728 VTAIL.n153 VTAIL.n151 2.84303
R1729 VTAIL.n89 VTAIL.n87 2.84303
R1730 VTAIL.n226 VTAIL.n206 2.71565
R1731 VTAIL.n247 VTAIL.n198 2.71565
R1732 VTAIL.n34 VTAIL.n14 2.71565
R1733 VTAIL.n55 VTAIL.n6 2.71565
R1734 VTAIL.n185 VTAIL.n136 2.71565
R1735 VTAIL.n166 VTAIL.n146 2.71565
R1736 VTAIL.n121 VTAIL.n72 2.71565
R1737 VTAIL.n102 VTAIL.n82 2.71565
R1738 VTAIL.n231 VTAIL.n229 1.93989
R1739 VTAIL.n244 VTAIL.n243 1.93989
R1740 VTAIL.n39 VTAIL.n37 1.93989
R1741 VTAIL.n52 VTAIL.n51 1.93989
R1742 VTAIL.n182 VTAIL.n181 1.93989
R1743 VTAIL.n170 VTAIL.n169 1.93989
R1744 VTAIL.n118 VTAIL.n117 1.93989
R1745 VTAIL.n106 VTAIL.n105 1.93989
R1746 VTAIL.n129 VTAIL.n67 1.93153
R1747 VTAIL.n193 VTAIL.n131 1.93153
R1748 VTAIL.n65 VTAIL.n63 1.93153
R1749 VTAIL.n0 VTAIL.t0 1.72524
R1750 VTAIL.n0 VTAIL.t2 1.72524
R1751 VTAIL.n64 VTAIL.t10 1.72524
R1752 VTAIL.n64 VTAIL.t8 1.72524
R1753 VTAIL.n130 VTAIL.t9 1.72524
R1754 VTAIL.n130 VTAIL.t5 1.72524
R1755 VTAIL.n66 VTAIL.t3 1.72524
R1756 VTAIL.n66 VTAIL.t4 1.72524
R1757 VTAIL.n131 VTAIL.n129 1.43584
R1758 VTAIL.n63 VTAIL.n1 1.43584
R1759 VTAIL VTAIL.n255 1.39059
R1760 VTAIL.n230 VTAIL.n204 1.16414
R1761 VTAIL.n240 VTAIL.n200 1.16414
R1762 VTAIL.n38 VTAIL.n12 1.16414
R1763 VTAIL.n48 VTAIL.n8 1.16414
R1764 VTAIL.n178 VTAIL.n138 1.16414
R1765 VTAIL.n173 VTAIL.n143 1.16414
R1766 VTAIL.n114 VTAIL.n74 1.16414
R1767 VTAIL.n109 VTAIL.n79 1.16414
R1768 VTAIL VTAIL.n1 0.541448
R1769 VTAIL.n236 VTAIL.n235 0.388379
R1770 VTAIL.n239 VTAIL.n202 0.388379
R1771 VTAIL.n44 VTAIL.n43 0.388379
R1772 VTAIL.n47 VTAIL.n10 0.388379
R1773 VTAIL.n177 VTAIL.n140 0.388379
R1774 VTAIL.n174 VTAIL.n142 0.388379
R1775 VTAIL.n113 VTAIL.n76 0.388379
R1776 VTAIL.n110 VTAIL.n78 0.388379
R1777 VTAIL.n219 VTAIL.n211 0.155672
R1778 VTAIL.n220 VTAIL.n219 0.155672
R1779 VTAIL.n220 VTAIL.n207 0.155672
R1780 VTAIL.n227 VTAIL.n207 0.155672
R1781 VTAIL.n228 VTAIL.n227 0.155672
R1782 VTAIL.n228 VTAIL.n203 0.155672
R1783 VTAIL.n237 VTAIL.n203 0.155672
R1784 VTAIL.n238 VTAIL.n237 0.155672
R1785 VTAIL.n238 VTAIL.n199 0.155672
R1786 VTAIL.n245 VTAIL.n199 0.155672
R1787 VTAIL.n246 VTAIL.n245 0.155672
R1788 VTAIL.n246 VTAIL.n195 0.155672
R1789 VTAIL.n253 VTAIL.n195 0.155672
R1790 VTAIL.n27 VTAIL.n19 0.155672
R1791 VTAIL.n28 VTAIL.n27 0.155672
R1792 VTAIL.n28 VTAIL.n15 0.155672
R1793 VTAIL.n35 VTAIL.n15 0.155672
R1794 VTAIL.n36 VTAIL.n35 0.155672
R1795 VTAIL.n36 VTAIL.n11 0.155672
R1796 VTAIL.n45 VTAIL.n11 0.155672
R1797 VTAIL.n46 VTAIL.n45 0.155672
R1798 VTAIL.n46 VTAIL.n7 0.155672
R1799 VTAIL.n53 VTAIL.n7 0.155672
R1800 VTAIL.n54 VTAIL.n53 0.155672
R1801 VTAIL.n54 VTAIL.n3 0.155672
R1802 VTAIL.n61 VTAIL.n3 0.155672
R1803 VTAIL.n191 VTAIL.n133 0.155672
R1804 VTAIL.n184 VTAIL.n133 0.155672
R1805 VTAIL.n184 VTAIL.n183 0.155672
R1806 VTAIL.n183 VTAIL.n137 0.155672
R1807 VTAIL.n176 VTAIL.n137 0.155672
R1808 VTAIL.n176 VTAIL.n175 0.155672
R1809 VTAIL.n175 VTAIL.n141 0.155672
R1810 VTAIL.n168 VTAIL.n141 0.155672
R1811 VTAIL.n168 VTAIL.n167 0.155672
R1812 VTAIL.n167 VTAIL.n147 0.155672
R1813 VTAIL.n160 VTAIL.n147 0.155672
R1814 VTAIL.n160 VTAIL.n159 0.155672
R1815 VTAIL.n159 VTAIL.n151 0.155672
R1816 VTAIL.n127 VTAIL.n69 0.155672
R1817 VTAIL.n120 VTAIL.n69 0.155672
R1818 VTAIL.n120 VTAIL.n119 0.155672
R1819 VTAIL.n119 VTAIL.n73 0.155672
R1820 VTAIL.n112 VTAIL.n73 0.155672
R1821 VTAIL.n112 VTAIL.n111 0.155672
R1822 VTAIL.n111 VTAIL.n77 0.155672
R1823 VTAIL.n104 VTAIL.n77 0.155672
R1824 VTAIL.n104 VTAIL.n103 0.155672
R1825 VTAIL.n103 VTAIL.n83 0.155672
R1826 VTAIL.n96 VTAIL.n83 0.155672
R1827 VTAIL.n96 VTAIL.n95 0.155672
R1828 VTAIL.n95 VTAIL.n87 0.155672
R1829 VDD1.n56 VDD1.n0 289.615
R1830 VDD1.n117 VDD1.n61 289.615
R1831 VDD1.n57 VDD1.n56 185
R1832 VDD1.n55 VDD1.n54 185
R1833 VDD1.n4 VDD1.n3 185
R1834 VDD1.n49 VDD1.n48 185
R1835 VDD1.n47 VDD1.n46 185
R1836 VDD1.n8 VDD1.n7 185
R1837 VDD1.n12 VDD1.n10 185
R1838 VDD1.n41 VDD1.n40 185
R1839 VDD1.n39 VDD1.n38 185
R1840 VDD1.n14 VDD1.n13 185
R1841 VDD1.n33 VDD1.n32 185
R1842 VDD1.n31 VDD1.n30 185
R1843 VDD1.n18 VDD1.n17 185
R1844 VDD1.n25 VDD1.n24 185
R1845 VDD1.n23 VDD1.n22 185
R1846 VDD1.n82 VDD1.n81 185
R1847 VDD1.n84 VDD1.n83 185
R1848 VDD1.n77 VDD1.n76 185
R1849 VDD1.n90 VDD1.n89 185
R1850 VDD1.n92 VDD1.n91 185
R1851 VDD1.n73 VDD1.n72 185
R1852 VDD1.n99 VDD1.n98 185
R1853 VDD1.n100 VDD1.n71 185
R1854 VDD1.n102 VDD1.n101 185
R1855 VDD1.n69 VDD1.n68 185
R1856 VDD1.n108 VDD1.n107 185
R1857 VDD1.n110 VDD1.n109 185
R1858 VDD1.n65 VDD1.n64 185
R1859 VDD1.n116 VDD1.n115 185
R1860 VDD1.n118 VDD1.n117 185
R1861 VDD1.n21 VDD1.t5 149.524
R1862 VDD1.n80 VDD1.t4 149.524
R1863 VDD1.n56 VDD1.n55 104.615
R1864 VDD1.n55 VDD1.n3 104.615
R1865 VDD1.n48 VDD1.n3 104.615
R1866 VDD1.n48 VDD1.n47 104.615
R1867 VDD1.n47 VDD1.n7 104.615
R1868 VDD1.n12 VDD1.n7 104.615
R1869 VDD1.n40 VDD1.n12 104.615
R1870 VDD1.n40 VDD1.n39 104.615
R1871 VDD1.n39 VDD1.n13 104.615
R1872 VDD1.n32 VDD1.n13 104.615
R1873 VDD1.n32 VDD1.n31 104.615
R1874 VDD1.n31 VDD1.n17 104.615
R1875 VDD1.n24 VDD1.n17 104.615
R1876 VDD1.n24 VDD1.n23 104.615
R1877 VDD1.n83 VDD1.n82 104.615
R1878 VDD1.n83 VDD1.n76 104.615
R1879 VDD1.n90 VDD1.n76 104.615
R1880 VDD1.n91 VDD1.n90 104.615
R1881 VDD1.n91 VDD1.n72 104.615
R1882 VDD1.n99 VDD1.n72 104.615
R1883 VDD1.n100 VDD1.n99 104.615
R1884 VDD1.n101 VDD1.n100 104.615
R1885 VDD1.n101 VDD1.n68 104.615
R1886 VDD1.n108 VDD1.n68 104.615
R1887 VDD1.n109 VDD1.n108 104.615
R1888 VDD1.n109 VDD1.n64 104.615
R1889 VDD1.n116 VDD1.n64 104.615
R1890 VDD1.n117 VDD1.n116 104.615
R1891 VDD1.n123 VDD1.n122 64.0687
R1892 VDD1.n125 VDD1.n124 63.6413
R1893 VDD1.n23 VDD1.t5 52.3082
R1894 VDD1.n82 VDD1.t4 52.3082
R1895 VDD1 VDD1.n60 51.9221
R1896 VDD1.n123 VDD1.n121 51.8086
R1897 VDD1.n125 VDD1.n123 41.4362
R1898 VDD1.n10 VDD1.n8 13.1884
R1899 VDD1.n102 VDD1.n69 13.1884
R1900 VDD1.n46 VDD1.n45 12.8005
R1901 VDD1.n42 VDD1.n41 12.8005
R1902 VDD1.n103 VDD1.n71 12.8005
R1903 VDD1.n107 VDD1.n106 12.8005
R1904 VDD1.n49 VDD1.n6 12.0247
R1905 VDD1.n38 VDD1.n11 12.0247
R1906 VDD1.n98 VDD1.n97 12.0247
R1907 VDD1.n110 VDD1.n67 12.0247
R1908 VDD1.n50 VDD1.n4 11.249
R1909 VDD1.n37 VDD1.n14 11.249
R1910 VDD1.n96 VDD1.n73 11.249
R1911 VDD1.n111 VDD1.n65 11.249
R1912 VDD1.n54 VDD1.n53 10.4732
R1913 VDD1.n34 VDD1.n33 10.4732
R1914 VDD1.n93 VDD1.n92 10.4732
R1915 VDD1.n115 VDD1.n114 10.4732
R1916 VDD1.n22 VDD1.n21 10.2747
R1917 VDD1.n81 VDD1.n80 10.2747
R1918 VDD1.n57 VDD1.n2 9.69747
R1919 VDD1.n30 VDD1.n16 9.69747
R1920 VDD1.n89 VDD1.n75 9.69747
R1921 VDD1.n118 VDD1.n63 9.69747
R1922 VDD1.n60 VDD1.n59 9.45567
R1923 VDD1.n121 VDD1.n120 9.45567
R1924 VDD1.n20 VDD1.n19 9.3005
R1925 VDD1.n27 VDD1.n26 9.3005
R1926 VDD1.n29 VDD1.n28 9.3005
R1927 VDD1.n16 VDD1.n15 9.3005
R1928 VDD1.n35 VDD1.n34 9.3005
R1929 VDD1.n37 VDD1.n36 9.3005
R1930 VDD1.n11 VDD1.n9 9.3005
R1931 VDD1.n43 VDD1.n42 9.3005
R1932 VDD1.n59 VDD1.n58 9.3005
R1933 VDD1.n2 VDD1.n1 9.3005
R1934 VDD1.n53 VDD1.n52 9.3005
R1935 VDD1.n51 VDD1.n50 9.3005
R1936 VDD1.n6 VDD1.n5 9.3005
R1937 VDD1.n45 VDD1.n44 9.3005
R1938 VDD1.n120 VDD1.n119 9.3005
R1939 VDD1.n63 VDD1.n62 9.3005
R1940 VDD1.n114 VDD1.n113 9.3005
R1941 VDD1.n112 VDD1.n111 9.3005
R1942 VDD1.n67 VDD1.n66 9.3005
R1943 VDD1.n106 VDD1.n105 9.3005
R1944 VDD1.n79 VDD1.n78 9.3005
R1945 VDD1.n86 VDD1.n85 9.3005
R1946 VDD1.n88 VDD1.n87 9.3005
R1947 VDD1.n75 VDD1.n74 9.3005
R1948 VDD1.n94 VDD1.n93 9.3005
R1949 VDD1.n96 VDD1.n95 9.3005
R1950 VDD1.n97 VDD1.n70 9.3005
R1951 VDD1.n104 VDD1.n103 9.3005
R1952 VDD1.n58 VDD1.n0 8.92171
R1953 VDD1.n29 VDD1.n18 8.92171
R1954 VDD1.n88 VDD1.n77 8.92171
R1955 VDD1.n119 VDD1.n61 8.92171
R1956 VDD1.n26 VDD1.n25 8.14595
R1957 VDD1.n85 VDD1.n84 8.14595
R1958 VDD1.n22 VDD1.n20 7.3702
R1959 VDD1.n81 VDD1.n79 7.3702
R1960 VDD1.n25 VDD1.n20 5.81868
R1961 VDD1.n84 VDD1.n79 5.81868
R1962 VDD1.n60 VDD1.n0 5.04292
R1963 VDD1.n26 VDD1.n18 5.04292
R1964 VDD1.n85 VDD1.n77 5.04292
R1965 VDD1.n121 VDD1.n61 5.04292
R1966 VDD1.n58 VDD1.n57 4.26717
R1967 VDD1.n30 VDD1.n29 4.26717
R1968 VDD1.n89 VDD1.n88 4.26717
R1969 VDD1.n119 VDD1.n118 4.26717
R1970 VDD1.n54 VDD1.n2 3.49141
R1971 VDD1.n33 VDD1.n16 3.49141
R1972 VDD1.n92 VDD1.n75 3.49141
R1973 VDD1.n115 VDD1.n63 3.49141
R1974 VDD1.n21 VDD1.n19 2.84303
R1975 VDD1.n80 VDD1.n78 2.84303
R1976 VDD1.n53 VDD1.n4 2.71565
R1977 VDD1.n34 VDD1.n14 2.71565
R1978 VDD1.n93 VDD1.n73 2.71565
R1979 VDD1.n114 VDD1.n65 2.71565
R1980 VDD1.n50 VDD1.n49 1.93989
R1981 VDD1.n38 VDD1.n37 1.93989
R1982 VDD1.n98 VDD1.n96 1.93989
R1983 VDD1.n111 VDD1.n110 1.93989
R1984 VDD1.n124 VDD1.t3 1.72524
R1985 VDD1.n124 VDD1.t2 1.72524
R1986 VDD1.n122 VDD1.t0 1.72524
R1987 VDD1.n122 VDD1.t1 1.72524
R1988 VDD1.n46 VDD1.n6 1.16414
R1989 VDD1.n41 VDD1.n11 1.16414
R1990 VDD1.n97 VDD1.n71 1.16414
R1991 VDD1.n107 VDD1.n67 1.16414
R1992 VDD1 VDD1.n125 0.425069
R1993 VDD1.n45 VDD1.n8 0.388379
R1994 VDD1.n42 VDD1.n10 0.388379
R1995 VDD1.n103 VDD1.n102 0.388379
R1996 VDD1.n106 VDD1.n69 0.388379
R1997 VDD1.n59 VDD1.n1 0.155672
R1998 VDD1.n52 VDD1.n1 0.155672
R1999 VDD1.n52 VDD1.n51 0.155672
R2000 VDD1.n51 VDD1.n5 0.155672
R2001 VDD1.n44 VDD1.n5 0.155672
R2002 VDD1.n44 VDD1.n43 0.155672
R2003 VDD1.n43 VDD1.n9 0.155672
R2004 VDD1.n36 VDD1.n9 0.155672
R2005 VDD1.n36 VDD1.n35 0.155672
R2006 VDD1.n35 VDD1.n15 0.155672
R2007 VDD1.n28 VDD1.n15 0.155672
R2008 VDD1.n28 VDD1.n27 0.155672
R2009 VDD1.n27 VDD1.n19 0.155672
R2010 VDD1.n86 VDD1.n78 0.155672
R2011 VDD1.n87 VDD1.n86 0.155672
R2012 VDD1.n87 VDD1.n74 0.155672
R2013 VDD1.n94 VDD1.n74 0.155672
R2014 VDD1.n95 VDD1.n94 0.155672
R2015 VDD1.n95 VDD1.n70 0.155672
R2016 VDD1.n104 VDD1.n70 0.155672
R2017 VDD1.n105 VDD1.n104 0.155672
R2018 VDD1.n105 VDD1.n66 0.155672
R2019 VDD1.n112 VDD1.n66 0.155672
R2020 VDD1.n113 VDD1.n112 0.155672
R2021 VDD1.n113 VDD1.n62 0.155672
R2022 VDD1.n120 VDD1.n62 0.155672
R2023 VN.n2 VN.t4 176.095
R2024 VN.n14 VN.t2 176.095
R2025 VN.n21 VN.n12 161.3
R2026 VN.n20 VN.n19 161.3
R2027 VN.n18 VN.n13 161.3
R2028 VN.n17 VN.n16 161.3
R2029 VN.n9 VN.n0 161.3
R2030 VN.n8 VN.n7 161.3
R2031 VN.n6 VN.n1 161.3
R2032 VN.n5 VN.n4 161.3
R2033 VN.n3 VN.t3 144.852
R2034 VN.n10 VN.t0 144.852
R2035 VN.n15 VN.t5 144.852
R2036 VN.n22 VN.t1 144.852
R2037 VN.n11 VN.n10 86.7496
R2038 VN.n23 VN.n22 86.7496
R2039 VN.n3 VN.n2 57.7381
R2040 VN.n15 VN.n14 57.7381
R2041 VN.n8 VN.n1 53.0692
R2042 VN.n20 VN.n13 53.0692
R2043 VN VN.n23 45.9224
R2044 VN.n9 VN.n8 27.752
R2045 VN.n21 VN.n20 27.752
R2046 VN.n4 VN.n1 24.3439
R2047 VN.n16 VN.n13 24.3439
R2048 VN.n10 VN.n9 23.8571
R2049 VN.n22 VN.n21 23.8571
R2050 VN.n17 VN.n14 12.7265
R2051 VN.n5 VN.n2 12.7265
R2052 VN.n4 VN.n3 12.1722
R2053 VN.n16 VN.n15 12.1722
R2054 VN.n23 VN.n12 0.278398
R2055 VN.n11 VN.n0 0.278398
R2056 VN.n19 VN.n12 0.189894
R2057 VN.n19 VN.n18 0.189894
R2058 VN.n18 VN.n17 0.189894
R2059 VN.n6 VN.n5 0.189894
R2060 VN.n7 VN.n6 0.189894
R2061 VN.n7 VN.n0 0.189894
R2062 VN VN.n11 0.153422
R2063 VDD2.n119 VDD2.n63 289.615
R2064 VDD2.n56 VDD2.n0 289.615
R2065 VDD2.n120 VDD2.n119 185
R2066 VDD2.n118 VDD2.n117 185
R2067 VDD2.n67 VDD2.n66 185
R2068 VDD2.n112 VDD2.n111 185
R2069 VDD2.n110 VDD2.n109 185
R2070 VDD2.n71 VDD2.n70 185
R2071 VDD2.n75 VDD2.n73 185
R2072 VDD2.n104 VDD2.n103 185
R2073 VDD2.n102 VDD2.n101 185
R2074 VDD2.n77 VDD2.n76 185
R2075 VDD2.n96 VDD2.n95 185
R2076 VDD2.n94 VDD2.n93 185
R2077 VDD2.n81 VDD2.n80 185
R2078 VDD2.n88 VDD2.n87 185
R2079 VDD2.n86 VDD2.n85 185
R2080 VDD2.n21 VDD2.n20 185
R2081 VDD2.n23 VDD2.n22 185
R2082 VDD2.n16 VDD2.n15 185
R2083 VDD2.n29 VDD2.n28 185
R2084 VDD2.n31 VDD2.n30 185
R2085 VDD2.n12 VDD2.n11 185
R2086 VDD2.n38 VDD2.n37 185
R2087 VDD2.n39 VDD2.n10 185
R2088 VDD2.n41 VDD2.n40 185
R2089 VDD2.n8 VDD2.n7 185
R2090 VDD2.n47 VDD2.n46 185
R2091 VDD2.n49 VDD2.n48 185
R2092 VDD2.n4 VDD2.n3 185
R2093 VDD2.n55 VDD2.n54 185
R2094 VDD2.n57 VDD2.n56 185
R2095 VDD2.n84 VDD2.t4 149.524
R2096 VDD2.n19 VDD2.t1 149.524
R2097 VDD2.n119 VDD2.n118 104.615
R2098 VDD2.n118 VDD2.n66 104.615
R2099 VDD2.n111 VDD2.n66 104.615
R2100 VDD2.n111 VDD2.n110 104.615
R2101 VDD2.n110 VDD2.n70 104.615
R2102 VDD2.n75 VDD2.n70 104.615
R2103 VDD2.n103 VDD2.n75 104.615
R2104 VDD2.n103 VDD2.n102 104.615
R2105 VDD2.n102 VDD2.n76 104.615
R2106 VDD2.n95 VDD2.n76 104.615
R2107 VDD2.n95 VDD2.n94 104.615
R2108 VDD2.n94 VDD2.n80 104.615
R2109 VDD2.n87 VDD2.n80 104.615
R2110 VDD2.n87 VDD2.n86 104.615
R2111 VDD2.n22 VDD2.n21 104.615
R2112 VDD2.n22 VDD2.n15 104.615
R2113 VDD2.n29 VDD2.n15 104.615
R2114 VDD2.n30 VDD2.n29 104.615
R2115 VDD2.n30 VDD2.n11 104.615
R2116 VDD2.n38 VDD2.n11 104.615
R2117 VDD2.n39 VDD2.n38 104.615
R2118 VDD2.n40 VDD2.n39 104.615
R2119 VDD2.n40 VDD2.n7 104.615
R2120 VDD2.n47 VDD2.n7 104.615
R2121 VDD2.n48 VDD2.n47 104.615
R2122 VDD2.n48 VDD2.n3 104.615
R2123 VDD2.n55 VDD2.n3 104.615
R2124 VDD2.n56 VDD2.n55 104.615
R2125 VDD2.n62 VDD2.n61 64.0687
R2126 VDD2 VDD2.n125 64.0658
R2127 VDD2.n86 VDD2.t4 52.3082
R2128 VDD2.n21 VDD2.t1 52.3082
R2129 VDD2.n62 VDD2.n60 51.8086
R2130 VDD2.n124 VDD2.n123 50.4157
R2131 VDD2.n124 VDD2.n62 39.8877
R2132 VDD2.n73 VDD2.n71 13.1884
R2133 VDD2.n41 VDD2.n8 13.1884
R2134 VDD2.n109 VDD2.n108 12.8005
R2135 VDD2.n105 VDD2.n104 12.8005
R2136 VDD2.n42 VDD2.n10 12.8005
R2137 VDD2.n46 VDD2.n45 12.8005
R2138 VDD2.n112 VDD2.n69 12.0247
R2139 VDD2.n101 VDD2.n74 12.0247
R2140 VDD2.n37 VDD2.n36 12.0247
R2141 VDD2.n49 VDD2.n6 12.0247
R2142 VDD2.n113 VDD2.n67 11.249
R2143 VDD2.n100 VDD2.n77 11.249
R2144 VDD2.n35 VDD2.n12 11.249
R2145 VDD2.n50 VDD2.n4 11.249
R2146 VDD2.n117 VDD2.n116 10.4732
R2147 VDD2.n97 VDD2.n96 10.4732
R2148 VDD2.n32 VDD2.n31 10.4732
R2149 VDD2.n54 VDD2.n53 10.4732
R2150 VDD2.n85 VDD2.n84 10.2747
R2151 VDD2.n20 VDD2.n19 10.2747
R2152 VDD2.n120 VDD2.n65 9.69747
R2153 VDD2.n93 VDD2.n79 9.69747
R2154 VDD2.n28 VDD2.n14 9.69747
R2155 VDD2.n57 VDD2.n2 9.69747
R2156 VDD2.n123 VDD2.n122 9.45567
R2157 VDD2.n60 VDD2.n59 9.45567
R2158 VDD2.n83 VDD2.n82 9.3005
R2159 VDD2.n90 VDD2.n89 9.3005
R2160 VDD2.n92 VDD2.n91 9.3005
R2161 VDD2.n79 VDD2.n78 9.3005
R2162 VDD2.n98 VDD2.n97 9.3005
R2163 VDD2.n100 VDD2.n99 9.3005
R2164 VDD2.n74 VDD2.n72 9.3005
R2165 VDD2.n106 VDD2.n105 9.3005
R2166 VDD2.n122 VDD2.n121 9.3005
R2167 VDD2.n65 VDD2.n64 9.3005
R2168 VDD2.n116 VDD2.n115 9.3005
R2169 VDD2.n114 VDD2.n113 9.3005
R2170 VDD2.n69 VDD2.n68 9.3005
R2171 VDD2.n108 VDD2.n107 9.3005
R2172 VDD2.n59 VDD2.n58 9.3005
R2173 VDD2.n2 VDD2.n1 9.3005
R2174 VDD2.n53 VDD2.n52 9.3005
R2175 VDD2.n51 VDD2.n50 9.3005
R2176 VDD2.n6 VDD2.n5 9.3005
R2177 VDD2.n45 VDD2.n44 9.3005
R2178 VDD2.n18 VDD2.n17 9.3005
R2179 VDD2.n25 VDD2.n24 9.3005
R2180 VDD2.n27 VDD2.n26 9.3005
R2181 VDD2.n14 VDD2.n13 9.3005
R2182 VDD2.n33 VDD2.n32 9.3005
R2183 VDD2.n35 VDD2.n34 9.3005
R2184 VDD2.n36 VDD2.n9 9.3005
R2185 VDD2.n43 VDD2.n42 9.3005
R2186 VDD2.n121 VDD2.n63 8.92171
R2187 VDD2.n92 VDD2.n81 8.92171
R2188 VDD2.n27 VDD2.n16 8.92171
R2189 VDD2.n58 VDD2.n0 8.92171
R2190 VDD2.n89 VDD2.n88 8.14595
R2191 VDD2.n24 VDD2.n23 8.14595
R2192 VDD2.n85 VDD2.n83 7.3702
R2193 VDD2.n20 VDD2.n18 7.3702
R2194 VDD2.n88 VDD2.n83 5.81868
R2195 VDD2.n23 VDD2.n18 5.81868
R2196 VDD2.n123 VDD2.n63 5.04292
R2197 VDD2.n89 VDD2.n81 5.04292
R2198 VDD2.n24 VDD2.n16 5.04292
R2199 VDD2.n60 VDD2.n0 5.04292
R2200 VDD2.n121 VDD2.n120 4.26717
R2201 VDD2.n93 VDD2.n92 4.26717
R2202 VDD2.n28 VDD2.n27 4.26717
R2203 VDD2.n58 VDD2.n57 4.26717
R2204 VDD2.n117 VDD2.n65 3.49141
R2205 VDD2.n96 VDD2.n79 3.49141
R2206 VDD2.n31 VDD2.n14 3.49141
R2207 VDD2.n54 VDD2.n2 3.49141
R2208 VDD2.n84 VDD2.n82 2.84303
R2209 VDD2.n19 VDD2.n17 2.84303
R2210 VDD2.n116 VDD2.n67 2.71565
R2211 VDD2.n97 VDD2.n77 2.71565
R2212 VDD2.n32 VDD2.n12 2.71565
R2213 VDD2.n53 VDD2.n4 2.71565
R2214 VDD2.n113 VDD2.n112 1.93989
R2215 VDD2.n101 VDD2.n100 1.93989
R2216 VDD2.n37 VDD2.n35 1.93989
R2217 VDD2.n50 VDD2.n49 1.93989
R2218 VDD2.n125 VDD2.t0 1.72524
R2219 VDD2.n125 VDD2.t3 1.72524
R2220 VDD2.n61 VDD2.t2 1.72524
R2221 VDD2.n61 VDD2.t5 1.72524
R2222 VDD2 VDD2.n124 1.50697
R2223 VDD2.n109 VDD2.n69 1.16414
R2224 VDD2.n104 VDD2.n74 1.16414
R2225 VDD2.n36 VDD2.n10 1.16414
R2226 VDD2.n46 VDD2.n6 1.16414
R2227 VDD2.n108 VDD2.n71 0.388379
R2228 VDD2.n105 VDD2.n73 0.388379
R2229 VDD2.n42 VDD2.n41 0.388379
R2230 VDD2.n45 VDD2.n8 0.388379
R2231 VDD2.n122 VDD2.n64 0.155672
R2232 VDD2.n115 VDD2.n64 0.155672
R2233 VDD2.n115 VDD2.n114 0.155672
R2234 VDD2.n114 VDD2.n68 0.155672
R2235 VDD2.n107 VDD2.n68 0.155672
R2236 VDD2.n107 VDD2.n106 0.155672
R2237 VDD2.n106 VDD2.n72 0.155672
R2238 VDD2.n99 VDD2.n72 0.155672
R2239 VDD2.n99 VDD2.n98 0.155672
R2240 VDD2.n98 VDD2.n78 0.155672
R2241 VDD2.n91 VDD2.n78 0.155672
R2242 VDD2.n91 VDD2.n90 0.155672
R2243 VDD2.n90 VDD2.n82 0.155672
R2244 VDD2.n25 VDD2.n17 0.155672
R2245 VDD2.n26 VDD2.n25 0.155672
R2246 VDD2.n26 VDD2.n13 0.155672
R2247 VDD2.n33 VDD2.n13 0.155672
R2248 VDD2.n34 VDD2.n33 0.155672
R2249 VDD2.n34 VDD2.n9 0.155672
R2250 VDD2.n43 VDD2.n9 0.155672
R2251 VDD2.n44 VDD2.n43 0.155672
R2252 VDD2.n44 VDD2.n5 0.155672
R2253 VDD2.n51 VDD2.n5 0.155672
R2254 VDD2.n52 VDD2.n51 0.155672
R2255 VDD2.n52 VDD2.n1 0.155672
R2256 VDD2.n59 VDD2.n1 0.155672
C0 VDD2 VTAIL 7.58671f
C1 VDD1 VN 0.149464f
C2 VDD1 VP 6.27383f
C3 VDD2 VN 6.02714f
C4 VN VTAIL 6.04881f
C5 VDD2 VP 0.39949f
C6 VP VTAIL 6.06316f
C7 VDD2 VDD1 1.16244f
C8 VDD1 VTAIL 7.54125f
C9 VP VN 6.16441f
C10 VDD2 B 5.337653f
C11 VDD1 B 5.430751f
C12 VTAIL B 7.143257f
C13 VN B 10.8773f
C14 VP B 9.400101f
C15 VDD2.n0 B 0.030844f
C16 VDD2.n1 B 0.02153f
C17 VDD2.n2 B 0.011569f
C18 VDD2.n3 B 0.027346f
C19 VDD2.n4 B 0.01225f
C20 VDD2.n5 B 0.02153f
C21 VDD2.n6 B 0.011569f
C22 VDD2.n7 B 0.027346f
C23 VDD2.n8 B 0.01191f
C24 VDD2.n9 B 0.02153f
C25 VDD2.n10 B 0.01225f
C26 VDD2.n11 B 0.027346f
C27 VDD2.n12 B 0.01225f
C28 VDD2.n13 B 0.02153f
C29 VDD2.n14 B 0.011569f
C30 VDD2.n15 B 0.027346f
C31 VDD2.n16 B 0.01225f
C32 VDD2.n17 B 1.03638f
C33 VDD2.n18 B 0.011569f
C34 VDD2.t1 B 0.046126f
C35 VDD2.n19 B 0.150934f
C36 VDD2.n20 B 0.019332f
C37 VDD2.n21 B 0.02051f
C38 VDD2.n22 B 0.027346f
C39 VDD2.n23 B 0.01225f
C40 VDD2.n24 B 0.011569f
C41 VDD2.n25 B 0.02153f
C42 VDD2.n26 B 0.02153f
C43 VDD2.n27 B 0.011569f
C44 VDD2.n28 B 0.01225f
C45 VDD2.n29 B 0.027346f
C46 VDD2.n30 B 0.027346f
C47 VDD2.n31 B 0.01225f
C48 VDD2.n32 B 0.011569f
C49 VDD2.n33 B 0.02153f
C50 VDD2.n34 B 0.02153f
C51 VDD2.n35 B 0.011569f
C52 VDD2.n36 B 0.011569f
C53 VDD2.n37 B 0.01225f
C54 VDD2.n38 B 0.027346f
C55 VDD2.n39 B 0.027346f
C56 VDD2.n40 B 0.027346f
C57 VDD2.n41 B 0.01191f
C58 VDD2.n42 B 0.011569f
C59 VDD2.n43 B 0.02153f
C60 VDD2.n44 B 0.02153f
C61 VDD2.n45 B 0.011569f
C62 VDD2.n46 B 0.01225f
C63 VDD2.n47 B 0.027346f
C64 VDD2.n48 B 0.027346f
C65 VDD2.n49 B 0.01225f
C66 VDD2.n50 B 0.011569f
C67 VDD2.n51 B 0.02153f
C68 VDD2.n52 B 0.02153f
C69 VDD2.n53 B 0.011569f
C70 VDD2.n54 B 0.01225f
C71 VDD2.n55 B 0.027346f
C72 VDD2.n56 B 0.060227f
C73 VDD2.n57 B 0.01225f
C74 VDD2.n58 B 0.011569f
C75 VDD2.n59 B 0.05212f
C76 VDD2.n60 B 0.052483f
C77 VDD2.t2 B 0.195321f
C78 VDD2.t5 B 0.195321f
C79 VDD2.n61 B 1.73923f
C80 VDD2.n62 B 2.02225f
C81 VDD2.n63 B 0.030844f
C82 VDD2.n64 B 0.02153f
C83 VDD2.n65 B 0.011569f
C84 VDD2.n66 B 0.027346f
C85 VDD2.n67 B 0.01225f
C86 VDD2.n68 B 0.02153f
C87 VDD2.n69 B 0.011569f
C88 VDD2.n70 B 0.027346f
C89 VDD2.n71 B 0.01191f
C90 VDD2.n72 B 0.02153f
C91 VDD2.n73 B 0.01191f
C92 VDD2.n74 B 0.011569f
C93 VDD2.n75 B 0.027346f
C94 VDD2.n76 B 0.027346f
C95 VDD2.n77 B 0.01225f
C96 VDD2.n78 B 0.02153f
C97 VDD2.n79 B 0.011569f
C98 VDD2.n80 B 0.027346f
C99 VDD2.n81 B 0.01225f
C100 VDD2.n82 B 1.03638f
C101 VDD2.n83 B 0.011569f
C102 VDD2.t4 B 0.046126f
C103 VDD2.n84 B 0.150934f
C104 VDD2.n85 B 0.019332f
C105 VDD2.n86 B 0.02051f
C106 VDD2.n87 B 0.027346f
C107 VDD2.n88 B 0.01225f
C108 VDD2.n89 B 0.011569f
C109 VDD2.n90 B 0.02153f
C110 VDD2.n91 B 0.02153f
C111 VDD2.n92 B 0.011569f
C112 VDD2.n93 B 0.01225f
C113 VDD2.n94 B 0.027346f
C114 VDD2.n95 B 0.027346f
C115 VDD2.n96 B 0.01225f
C116 VDD2.n97 B 0.011569f
C117 VDD2.n98 B 0.02153f
C118 VDD2.n99 B 0.02153f
C119 VDD2.n100 B 0.011569f
C120 VDD2.n101 B 0.01225f
C121 VDD2.n102 B 0.027346f
C122 VDD2.n103 B 0.027346f
C123 VDD2.n104 B 0.01225f
C124 VDD2.n105 B 0.011569f
C125 VDD2.n106 B 0.02153f
C126 VDD2.n107 B 0.02153f
C127 VDD2.n108 B 0.011569f
C128 VDD2.n109 B 0.01225f
C129 VDD2.n110 B 0.027346f
C130 VDD2.n111 B 0.027346f
C131 VDD2.n112 B 0.01225f
C132 VDD2.n113 B 0.011569f
C133 VDD2.n114 B 0.02153f
C134 VDD2.n115 B 0.02153f
C135 VDD2.n116 B 0.011569f
C136 VDD2.n117 B 0.01225f
C137 VDD2.n118 B 0.027346f
C138 VDD2.n119 B 0.060227f
C139 VDD2.n120 B 0.01225f
C140 VDD2.n121 B 0.011569f
C141 VDD2.n122 B 0.05212f
C142 VDD2.n123 B 0.048725f
C143 VDD2.n124 B 2.01042f
C144 VDD2.t0 B 0.195321f
C145 VDD2.t3 B 0.195321f
C146 VDD2.n125 B 1.7392f
C147 VN.n0 B 0.037263f
C148 VN.t0 B 1.68627f
C149 VN.n1 B 0.050391f
C150 VN.t4 B 1.81825f
C151 VN.n2 B 0.678302f
C152 VN.t3 B 1.68627f
C153 VN.n3 B 0.67104f
C154 VN.n4 B 0.039869f
C155 VN.n5 B 0.209187f
C156 VN.n6 B 0.028262f
C157 VN.n7 B 0.028262f
C158 VN.n8 B 0.029723f
C159 VN.n9 B 0.055176f
C160 VN.n10 B 0.695559f
C161 VN.n11 B 0.030312f
C162 VN.n12 B 0.037263f
C163 VN.t1 B 1.68627f
C164 VN.n13 B 0.050391f
C165 VN.t2 B 1.81825f
C166 VN.n14 B 0.678302f
C167 VN.t5 B 1.68627f
C168 VN.n15 B 0.67104f
C169 VN.n16 B 0.039869f
C170 VN.n17 B 0.209187f
C171 VN.n18 B 0.028262f
C172 VN.n19 B 0.028262f
C173 VN.n20 B 0.029723f
C174 VN.n21 B 0.055176f
C175 VN.n22 B 0.695559f
C176 VN.n23 B 1.37063f
C177 VDD1.n0 B 0.031116f
C178 VDD1.n1 B 0.02172f
C179 VDD1.n2 B 0.011671f
C180 VDD1.n3 B 0.027587f
C181 VDD1.n4 B 0.012358f
C182 VDD1.n5 B 0.02172f
C183 VDD1.n6 B 0.011671f
C184 VDD1.n7 B 0.027587f
C185 VDD1.n8 B 0.012015f
C186 VDD1.n9 B 0.02172f
C187 VDD1.n10 B 0.012015f
C188 VDD1.n11 B 0.011671f
C189 VDD1.n12 B 0.027587f
C190 VDD1.n13 B 0.027587f
C191 VDD1.n14 B 0.012358f
C192 VDD1.n15 B 0.02172f
C193 VDD1.n16 B 0.011671f
C194 VDD1.n17 B 0.027587f
C195 VDD1.n18 B 0.012358f
C196 VDD1.n19 B 1.0455f
C197 VDD1.n20 B 0.011671f
C198 VDD1.t5 B 0.046532f
C199 VDD1.n21 B 0.152264f
C200 VDD1.n22 B 0.019502f
C201 VDD1.n23 B 0.02069f
C202 VDD1.n24 B 0.027587f
C203 VDD1.n25 B 0.012358f
C204 VDD1.n26 B 0.011671f
C205 VDD1.n27 B 0.02172f
C206 VDD1.n28 B 0.02172f
C207 VDD1.n29 B 0.011671f
C208 VDD1.n30 B 0.012358f
C209 VDD1.n31 B 0.027587f
C210 VDD1.n32 B 0.027587f
C211 VDD1.n33 B 0.012358f
C212 VDD1.n34 B 0.011671f
C213 VDD1.n35 B 0.02172f
C214 VDD1.n36 B 0.02172f
C215 VDD1.n37 B 0.011671f
C216 VDD1.n38 B 0.012358f
C217 VDD1.n39 B 0.027587f
C218 VDD1.n40 B 0.027587f
C219 VDD1.n41 B 0.012358f
C220 VDD1.n42 B 0.011671f
C221 VDD1.n43 B 0.02172f
C222 VDD1.n44 B 0.02172f
C223 VDD1.n45 B 0.011671f
C224 VDD1.n46 B 0.012358f
C225 VDD1.n47 B 0.027587f
C226 VDD1.n48 B 0.027587f
C227 VDD1.n49 B 0.012358f
C228 VDD1.n50 B 0.011671f
C229 VDD1.n51 B 0.02172f
C230 VDD1.n52 B 0.02172f
C231 VDD1.n53 B 0.011671f
C232 VDD1.n54 B 0.012358f
C233 VDD1.n55 B 0.027587f
C234 VDD1.n56 B 0.060758f
C235 VDD1.n57 B 0.012358f
C236 VDD1.n58 B 0.011671f
C237 VDD1.n59 B 0.052579f
C238 VDD1.n60 B 0.053466f
C239 VDD1.n61 B 0.031116f
C240 VDD1.n62 B 0.02172f
C241 VDD1.n63 B 0.011671f
C242 VDD1.n64 B 0.027587f
C243 VDD1.n65 B 0.012358f
C244 VDD1.n66 B 0.02172f
C245 VDD1.n67 B 0.011671f
C246 VDD1.n68 B 0.027587f
C247 VDD1.n69 B 0.012015f
C248 VDD1.n70 B 0.02172f
C249 VDD1.n71 B 0.012358f
C250 VDD1.n72 B 0.027587f
C251 VDD1.n73 B 0.012358f
C252 VDD1.n74 B 0.02172f
C253 VDD1.n75 B 0.011671f
C254 VDD1.n76 B 0.027587f
C255 VDD1.n77 B 0.012358f
C256 VDD1.n78 B 1.0455f
C257 VDD1.n79 B 0.011671f
C258 VDD1.t4 B 0.046532f
C259 VDD1.n80 B 0.152264f
C260 VDD1.n81 B 0.019502f
C261 VDD1.n82 B 0.02069f
C262 VDD1.n83 B 0.027587f
C263 VDD1.n84 B 0.012358f
C264 VDD1.n85 B 0.011671f
C265 VDD1.n86 B 0.02172f
C266 VDD1.n87 B 0.02172f
C267 VDD1.n88 B 0.011671f
C268 VDD1.n89 B 0.012358f
C269 VDD1.n90 B 0.027587f
C270 VDD1.n91 B 0.027587f
C271 VDD1.n92 B 0.012358f
C272 VDD1.n93 B 0.011671f
C273 VDD1.n94 B 0.02172f
C274 VDD1.n95 B 0.02172f
C275 VDD1.n96 B 0.011671f
C276 VDD1.n97 B 0.011671f
C277 VDD1.n98 B 0.012358f
C278 VDD1.n99 B 0.027587f
C279 VDD1.n100 B 0.027587f
C280 VDD1.n101 B 0.027587f
C281 VDD1.n102 B 0.012015f
C282 VDD1.n103 B 0.011671f
C283 VDD1.n104 B 0.02172f
C284 VDD1.n105 B 0.02172f
C285 VDD1.n106 B 0.011671f
C286 VDD1.n107 B 0.012358f
C287 VDD1.n108 B 0.027587f
C288 VDD1.n109 B 0.027587f
C289 VDD1.n110 B 0.012358f
C290 VDD1.n111 B 0.011671f
C291 VDD1.n112 B 0.02172f
C292 VDD1.n113 B 0.02172f
C293 VDD1.n114 B 0.011671f
C294 VDD1.n115 B 0.012358f
C295 VDD1.n116 B 0.027587f
C296 VDD1.n117 B 0.060758f
C297 VDD1.n118 B 0.012358f
C298 VDD1.n119 B 0.011671f
C299 VDD1.n120 B 0.052579f
C300 VDD1.n121 B 0.052945f
C301 VDD1.t0 B 0.197041f
C302 VDD1.t1 B 0.197041f
C303 VDD1.n122 B 1.75455f
C304 VDD1.n123 B 2.13224f
C305 VDD1.t3 B 0.197041f
C306 VDD1.t2 B 0.197041f
C307 VDD1.n124 B 1.75219f
C308 VDD1.n125 B 2.21911f
C309 VTAIL.t0 B 0.212887f
C310 VTAIL.t2 B 0.212887f
C311 VTAIL.n0 B 1.8264f
C312 VTAIL.n1 B 0.376504f
C313 VTAIL.n2 B 0.033618f
C314 VTAIL.n3 B 0.023467f
C315 VTAIL.n4 B 0.01261f
C316 VTAIL.n5 B 0.029806f
C317 VTAIL.n6 B 0.013352f
C318 VTAIL.n7 B 0.023467f
C319 VTAIL.n8 B 0.01261f
C320 VTAIL.n9 B 0.029806f
C321 VTAIL.n10 B 0.012981f
C322 VTAIL.n11 B 0.023467f
C323 VTAIL.n12 B 0.013352f
C324 VTAIL.n13 B 0.029806f
C325 VTAIL.n14 B 0.013352f
C326 VTAIL.n15 B 0.023467f
C327 VTAIL.n16 B 0.01261f
C328 VTAIL.n17 B 0.029806f
C329 VTAIL.n18 B 0.013352f
C330 VTAIL.n19 B 1.12958f
C331 VTAIL.n20 B 0.01261f
C332 VTAIL.t6 B 0.050274f
C333 VTAIL.n21 B 0.164509f
C334 VTAIL.n22 B 0.02107f
C335 VTAIL.n23 B 0.022354f
C336 VTAIL.n24 B 0.029806f
C337 VTAIL.n25 B 0.013352f
C338 VTAIL.n26 B 0.01261f
C339 VTAIL.n27 B 0.023467f
C340 VTAIL.n28 B 0.023467f
C341 VTAIL.n29 B 0.01261f
C342 VTAIL.n30 B 0.013352f
C343 VTAIL.n31 B 0.029806f
C344 VTAIL.n32 B 0.029806f
C345 VTAIL.n33 B 0.013352f
C346 VTAIL.n34 B 0.01261f
C347 VTAIL.n35 B 0.023467f
C348 VTAIL.n36 B 0.023467f
C349 VTAIL.n37 B 0.01261f
C350 VTAIL.n38 B 0.01261f
C351 VTAIL.n39 B 0.013352f
C352 VTAIL.n40 B 0.029806f
C353 VTAIL.n41 B 0.029806f
C354 VTAIL.n42 B 0.029806f
C355 VTAIL.n43 B 0.012981f
C356 VTAIL.n44 B 0.01261f
C357 VTAIL.n45 B 0.023467f
C358 VTAIL.n46 B 0.023467f
C359 VTAIL.n47 B 0.01261f
C360 VTAIL.n48 B 0.013352f
C361 VTAIL.n49 B 0.029806f
C362 VTAIL.n50 B 0.029806f
C363 VTAIL.n51 B 0.013352f
C364 VTAIL.n52 B 0.01261f
C365 VTAIL.n53 B 0.023467f
C366 VTAIL.n54 B 0.023467f
C367 VTAIL.n55 B 0.01261f
C368 VTAIL.n56 B 0.013352f
C369 VTAIL.n57 B 0.029806f
C370 VTAIL.n58 B 0.065644f
C371 VTAIL.n59 B 0.013352f
C372 VTAIL.n60 B 0.01261f
C373 VTAIL.n61 B 0.056807f
C374 VTAIL.n62 B 0.036923f
C375 VTAIL.n63 B 0.276041f
C376 VTAIL.t10 B 0.212887f
C377 VTAIL.t8 B 0.212887f
C378 VTAIL.n64 B 1.8264f
C379 VTAIL.n65 B 1.73221f
C380 VTAIL.t3 B 0.212887f
C381 VTAIL.t4 B 0.212887f
C382 VTAIL.n66 B 1.82641f
C383 VTAIL.n67 B 1.7322f
C384 VTAIL.n68 B 0.033618f
C385 VTAIL.n69 B 0.023467f
C386 VTAIL.n70 B 0.01261f
C387 VTAIL.n71 B 0.029806f
C388 VTAIL.n72 B 0.013352f
C389 VTAIL.n73 B 0.023467f
C390 VTAIL.n74 B 0.01261f
C391 VTAIL.n75 B 0.029806f
C392 VTAIL.n76 B 0.012981f
C393 VTAIL.n77 B 0.023467f
C394 VTAIL.n78 B 0.012981f
C395 VTAIL.n79 B 0.01261f
C396 VTAIL.n80 B 0.029806f
C397 VTAIL.n81 B 0.029806f
C398 VTAIL.n82 B 0.013352f
C399 VTAIL.n83 B 0.023467f
C400 VTAIL.n84 B 0.01261f
C401 VTAIL.n85 B 0.029806f
C402 VTAIL.n86 B 0.013352f
C403 VTAIL.n87 B 1.12958f
C404 VTAIL.n88 B 0.01261f
C405 VTAIL.t11 B 0.050274f
C406 VTAIL.n89 B 0.164509f
C407 VTAIL.n90 B 0.02107f
C408 VTAIL.n91 B 0.022354f
C409 VTAIL.n92 B 0.029806f
C410 VTAIL.n93 B 0.013352f
C411 VTAIL.n94 B 0.01261f
C412 VTAIL.n95 B 0.023467f
C413 VTAIL.n96 B 0.023467f
C414 VTAIL.n97 B 0.01261f
C415 VTAIL.n98 B 0.013352f
C416 VTAIL.n99 B 0.029806f
C417 VTAIL.n100 B 0.029806f
C418 VTAIL.n101 B 0.013352f
C419 VTAIL.n102 B 0.01261f
C420 VTAIL.n103 B 0.023467f
C421 VTAIL.n104 B 0.023467f
C422 VTAIL.n105 B 0.01261f
C423 VTAIL.n106 B 0.013352f
C424 VTAIL.n107 B 0.029806f
C425 VTAIL.n108 B 0.029806f
C426 VTAIL.n109 B 0.013352f
C427 VTAIL.n110 B 0.01261f
C428 VTAIL.n111 B 0.023467f
C429 VTAIL.n112 B 0.023467f
C430 VTAIL.n113 B 0.01261f
C431 VTAIL.n114 B 0.013352f
C432 VTAIL.n115 B 0.029806f
C433 VTAIL.n116 B 0.029806f
C434 VTAIL.n117 B 0.013352f
C435 VTAIL.n118 B 0.01261f
C436 VTAIL.n119 B 0.023467f
C437 VTAIL.n120 B 0.023467f
C438 VTAIL.n121 B 0.01261f
C439 VTAIL.n122 B 0.013352f
C440 VTAIL.n123 B 0.029806f
C441 VTAIL.n124 B 0.065644f
C442 VTAIL.n125 B 0.013352f
C443 VTAIL.n126 B 0.01261f
C444 VTAIL.n127 B 0.056807f
C445 VTAIL.n128 B 0.036923f
C446 VTAIL.n129 B 0.276041f
C447 VTAIL.t9 B 0.212887f
C448 VTAIL.t5 B 0.212887f
C449 VTAIL.n130 B 1.82641f
C450 VTAIL.n131 B 0.481606f
C451 VTAIL.n132 B 0.033618f
C452 VTAIL.n133 B 0.023467f
C453 VTAIL.n134 B 0.01261f
C454 VTAIL.n135 B 0.029806f
C455 VTAIL.n136 B 0.013352f
C456 VTAIL.n137 B 0.023467f
C457 VTAIL.n138 B 0.01261f
C458 VTAIL.n139 B 0.029806f
C459 VTAIL.n140 B 0.012981f
C460 VTAIL.n141 B 0.023467f
C461 VTAIL.n142 B 0.012981f
C462 VTAIL.n143 B 0.01261f
C463 VTAIL.n144 B 0.029806f
C464 VTAIL.n145 B 0.029806f
C465 VTAIL.n146 B 0.013352f
C466 VTAIL.n147 B 0.023467f
C467 VTAIL.n148 B 0.01261f
C468 VTAIL.n149 B 0.029806f
C469 VTAIL.n150 B 0.013352f
C470 VTAIL.n151 B 1.12958f
C471 VTAIL.n152 B 0.01261f
C472 VTAIL.t7 B 0.050274f
C473 VTAIL.n153 B 0.164509f
C474 VTAIL.n154 B 0.02107f
C475 VTAIL.n155 B 0.022354f
C476 VTAIL.n156 B 0.029806f
C477 VTAIL.n157 B 0.013352f
C478 VTAIL.n158 B 0.01261f
C479 VTAIL.n159 B 0.023467f
C480 VTAIL.n160 B 0.023467f
C481 VTAIL.n161 B 0.01261f
C482 VTAIL.n162 B 0.013352f
C483 VTAIL.n163 B 0.029806f
C484 VTAIL.n164 B 0.029806f
C485 VTAIL.n165 B 0.013352f
C486 VTAIL.n166 B 0.01261f
C487 VTAIL.n167 B 0.023467f
C488 VTAIL.n168 B 0.023467f
C489 VTAIL.n169 B 0.01261f
C490 VTAIL.n170 B 0.013352f
C491 VTAIL.n171 B 0.029806f
C492 VTAIL.n172 B 0.029806f
C493 VTAIL.n173 B 0.013352f
C494 VTAIL.n174 B 0.01261f
C495 VTAIL.n175 B 0.023467f
C496 VTAIL.n176 B 0.023467f
C497 VTAIL.n177 B 0.01261f
C498 VTAIL.n178 B 0.013352f
C499 VTAIL.n179 B 0.029806f
C500 VTAIL.n180 B 0.029806f
C501 VTAIL.n181 B 0.013352f
C502 VTAIL.n182 B 0.01261f
C503 VTAIL.n183 B 0.023467f
C504 VTAIL.n184 B 0.023467f
C505 VTAIL.n185 B 0.01261f
C506 VTAIL.n186 B 0.013352f
C507 VTAIL.n187 B 0.029806f
C508 VTAIL.n188 B 0.065644f
C509 VTAIL.n189 B 0.013352f
C510 VTAIL.n190 B 0.01261f
C511 VTAIL.n191 B 0.056807f
C512 VTAIL.n192 B 0.036923f
C513 VTAIL.n193 B 1.38062f
C514 VTAIL.n194 B 0.033618f
C515 VTAIL.n195 B 0.023467f
C516 VTAIL.n196 B 0.01261f
C517 VTAIL.n197 B 0.029806f
C518 VTAIL.n198 B 0.013352f
C519 VTAIL.n199 B 0.023467f
C520 VTAIL.n200 B 0.01261f
C521 VTAIL.n201 B 0.029806f
C522 VTAIL.n202 B 0.012981f
C523 VTAIL.n203 B 0.023467f
C524 VTAIL.n204 B 0.013352f
C525 VTAIL.n205 B 0.029806f
C526 VTAIL.n206 B 0.013352f
C527 VTAIL.n207 B 0.023467f
C528 VTAIL.n208 B 0.01261f
C529 VTAIL.n209 B 0.029806f
C530 VTAIL.n210 B 0.013352f
C531 VTAIL.n211 B 1.12958f
C532 VTAIL.n212 B 0.01261f
C533 VTAIL.t1 B 0.050274f
C534 VTAIL.n213 B 0.164509f
C535 VTAIL.n214 B 0.02107f
C536 VTAIL.n215 B 0.022354f
C537 VTAIL.n216 B 0.029806f
C538 VTAIL.n217 B 0.013352f
C539 VTAIL.n218 B 0.01261f
C540 VTAIL.n219 B 0.023467f
C541 VTAIL.n220 B 0.023467f
C542 VTAIL.n221 B 0.01261f
C543 VTAIL.n222 B 0.013352f
C544 VTAIL.n223 B 0.029806f
C545 VTAIL.n224 B 0.029806f
C546 VTAIL.n225 B 0.013352f
C547 VTAIL.n226 B 0.01261f
C548 VTAIL.n227 B 0.023467f
C549 VTAIL.n228 B 0.023467f
C550 VTAIL.n229 B 0.01261f
C551 VTAIL.n230 B 0.01261f
C552 VTAIL.n231 B 0.013352f
C553 VTAIL.n232 B 0.029806f
C554 VTAIL.n233 B 0.029806f
C555 VTAIL.n234 B 0.029806f
C556 VTAIL.n235 B 0.012981f
C557 VTAIL.n236 B 0.01261f
C558 VTAIL.n237 B 0.023467f
C559 VTAIL.n238 B 0.023467f
C560 VTAIL.n239 B 0.01261f
C561 VTAIL.n240 B 0.013352f
C562 VTAIL.n241 B 0.029806f
C563 VTAIL.n242 B 0.029806f
C564 VTAIL.n243 B 0.013352f
C565 VTAIL.n244 B 0.01261f
C566 VTAIL.n245 B 0.023467f
C567 VTAIL.n246 B 0.023467f
C568 VTAIL.n247 B 0.01261f
C569 VTAIL.n248 B 0.013352f
C570 VTAIL.n249 B 0.029806f
C571 VTAIL.n250 B 0.065644f
C572 VTAIL.n251 B 0.013352f
C573 VTAIL.n252 B 0.01261f
C574 VTAIL.n253 B 0.056807f
C575 VTAIL.n254 B 0.036923f
C576 VTAIL.n255 B 1.33972f
C577 VP.n0 B 0.038166f
C578 VP.t4 B 1.7271f
C579 VP.n1 B 0.051612f
C580 VP.n2 B 0.028947f
C581 VP.t5 B 1.7271f
C582 VP.n3 B 0.030443f
C583 VP.n4 B 0.038166f
C584 VP.t3 B 1.7271f
C585 VP.n5 B 0.051612f
C586 VP.t0 B 1.86228f
C587 VP.n6 B 0.694726f
C588 VP.t2 B 1.7271f
C589 VP.n7 B 0.687288f
C590 VP.n8 B 0.040835f
C591 VP.n9 B 0.214252f
C592 VP.n10 B 0.028947f
C593 VP.n11 B 0.028947f
C594 VP.n12 B 0.030443f
C595 VP.n13 B 0.056512f
C596 VP.n14 B 0.712401f
C597 VP.n15 B 1.38802f
C598 VP.n16 B 1.41075f
C599 VP.t1 B 1.7271f
C600 VP.n17 B 0.712401f
C601 VP.n18 B 0.056512f
C602 VP.n19 B 0.038166f
C603 VP.n20 B 0.028947f
C604 VP.n21 B 0.028947f
C605 VP.n22 B 0.051612f
C606 VP.n23 B 0.040835f
C607 VP.n24 B 0.619687f
C608 VP.n25 B 0.040835f
C609 VP.n26 B 0.028947f
C610 VP.n27 B 0.028947f
C611 VP.n28 B 0.028947f
C612 VP.n29 B 0.030443f
C613 VP.n30 B 0.056512f
C614 VP.n31 B 0.712401f
C615 VP.n32 B 0.031046f
.ends

