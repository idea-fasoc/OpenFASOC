* NGSPICE file created from diff_pair_sample_0746.ext - technology: sky130A

.subckt diff_pair_sample_0746 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X1 VTAIL.t18 VN.t0 VDD2.t9 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X2 VDD1.t8 VP.t1 VTAIL.t10 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X3 B.t11 B.t9 B.t10 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=3.98
X4 VTAIL.t2 VN.t1 VDD2.t8 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X5 VDD2.t7 VN.t2 VTAIL.t4 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.27885 ps=2.02 w=1.69 l=3.98
X6 VDD1.t7 VP.t2 VTAIL.t17 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.27885 ps=2.02 w=1.69 l=3.98
X7 VDD1.t6 VP.t3 VTAIL.t11 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.27885 ps=2.02 w=1.69 l=3.98
X8 VTAIL.t8 VP.t4 VDD1.t5 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X9 VDD2.t6 VN.t3 VTAIL.t1 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.6591 ps=4.16 w=1.69 l=3.98
X10 VTAIL.t14 VP.t5 VDD1.t4 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X11 B.t8 B.t6 B.t7 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=3.98
X12 B.t5 B.t3 B.t4 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=3.98
X13 VDD1.t3 VP.t6 VTAIL.t13 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.6591 ps=4.16 w=1.69 l=3.98
X14 VTAIL.t16 VP.t7 VDD1.t2 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X15 VTAIL.t0 VN.t4 VDD2.t5 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X16 VDD2.t4 VN.t5 VTAIL.t5 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X17 VTAIL.t19 VN.t6 VDD2.t3 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X18 VDD2.t2 VN.t7 VTAIL.t3 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.6591 ps=4.16 w=1.69 l=3.98
X19 VDD2.t1 VN.t8 VTAIL.t7 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
X20 VDD2.t0 VN.t9 VTAIL.t6 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.27885 ps=2.02 w=1.69 l=3.98
X21 VDD1.t1 VP.t8 VTAIL.t9 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.6591 ps=4.16 w=1.69 l=3.98
X22 B.t2 B.t0 B.t1 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=3.98
X23 VTAIL.t15 VP.t9 VDD1.t0 w_n6142_n1306# sky130_fd_pr__pfet_01v8 ad=0.27885 pd=2.02 as=0.27885 ps=2.02 w=1.69 l=3.98
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n46 VP.n45 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n59 VP.n58 161.3
R17 VP.n60 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n73 VP.n18 161.3
R26 VP.n130 VP.n0 161.3
R27 VP.n129 VP.n128 161.3
R28 VP.n127 VP.n1 161.3
R29 VP.n126 VP.n125 161.3
R30 VP.n124 VP.n2 161.3
R31 VP.n123 VP.n122 161.3
R32 VP.n121 VP.n3 161.3
R33 VP.n120 VP.n119 161.3
R34 VP.n117 VP.n4 161.3
R35 VP.n116 VP.n115 161.3
R36 VP.n114 VP.n5 161.3
R37 VP.n113 VP.n112 161.3
R38 VP.n111 VP.n6 161.3
R39 VP.n110 VP.n109 161.3
R40 VP.n108 VP.n7 161.3
R41 VP.n107 VP.n106 161.3
R42 VP.n105 VP.n8 161.3
R43 VP.n103 VP.n102 161.3
R44 VP.n101 VP.n9 161.3
R45 VP.n100 VP.n99 161.3
R46 VP.n98 VP.n10 161.3
R47 VP.n97 VP.n96 161.3
R48 VP.n95 VP.n11 161.3
R49 VP.n94 VP.n93 161.3
R50 VP.n92 VP.n12 161.3
R51 VP.n91 VP.n90 161.3
R52 VP.n89 VP.n88 161.3
R53 VP.n87 VP.n14 161.3
R54 VP.n86 VP.n85 161.3
R55 VP.n84 VP.n15 161.3
R56 VP.n83 VP.n82 161.3
R57 VP.n81 VP.n16 161.3
R58 VP.n80 VP.n79 161.3
R59 VP.n78 VP.n17 161.3
R60 VP.n32 VP.n31 72.0574
R61 VP.n77 VP.n76 64.0762
R62 VP.n132 VP.n131 64.0762
R63 VP.n75 VP.n74 64.0762
R64 VP.n82 VP.n15 56.5193
R65 VP.n125 VP.n124 56.5193
R66 VP.n68 VP.n67 56.5193
R67 VP.n77 VP.n75 53.0154
R68 VP.n98 VP.n97 49.7204
R69 VP.n111 VP.n110 49.7204
R70 VP.n54 VP.n53 49.7204
R71 VP.n41 VP.n40 49.7204
R72 VP.n32 VP.t2 42.5531
R73 VP.n97 VP.n11 31.2664
R74 VP.n112 VP.n111 31.2664
R75 VP.n55 VP.n54 31.2664
R76 VP.n40 VP.n29 31.2664
R77 VP.n80 VP.n17 24.4675
R78 VP.n81 VP.n80 24.4675
R79 VP.n82 VP.n81 24.4675
R80 VP.n86 VP.n15 24.4675
R81 VP.n87 VP.n86 24.4675
R82 VP.n88 VP.n87 24.4675
R83 VP.n92 VP.n91 24.4675
R84 VP.n93 VP.n92 24.4675
R85 VP.n93 VP.n11 24.4675
R86 VP.n99 VP.n98 24.4675
R87 VP.n99 VP.n9 24.4675
R88 VP.n103 VP.n9 24.4675
R89 VP.n106 VP.n105 24.4675
R90 VP.n106 VP.n7 24.4675
R91 VP.n110 VP.n7 24.4675
R92 VP.n112 VP.n5 24.4675
R93 VP.n116 VP.n5 24.4675
R94 VP.n117 VP.n116 24.4675
R95 VP.n119 VP.n3 24.4675
R96 VP.n123 VP.n3 24.4675
R97 VP.n124 VP.n123 24.4675
R98 VP.n125 VP.n1 24.4675
R99 VP.n129 VP.n1 24.4675
R100 VP.n130 VP.n129 24.4675
R101 VP.n68 VP.n19 24.4675
R102 VP.n72 VP.n19 24.4675
R103 VP.n73 VP.n72 24.4675
R104 VP.n55 VP.n23 24.4675
R105 VP.n59 VP.n23 24.4675
R106 VP.n60 VP.n59 24.4675
R107 VP.n62 VP.n21 24.4675
R108 VP.n66 VP.n21 24.4675
R109 VP.n67 VP.n66 24.4675
R110 VP.n42 VP.n41 24.4675
R111 VP.n42 VP.n27 24.4675
R112 VP.n46 VP.n27 24.4675
R113 VP.n49 VP.n48 24.4675
R114 VP.n49 VP.n25 24.4675
R115 VP.n53 VP.n25 24.4675
R116 VP.n35 VP.n34 24.4675
R117 VP.n36 VP.n35 24.4675
R118 VP.n36 VP.n29 24.4675
R119 VP.n88 VP.n13 21.5315
R120 VP.n119 VP.n118 21.5315
R121 VP.n62 VP.n61 21.5315
R122 VP.n76 VP.n17 18.1061
R123 VP.n131 VP.n130 18.1061
R124 VP.n74 VP.n73 18.1061
R125 VP.n104 VP.n103 12.234
R126 VP.n105 VP.n104 12.234
R127 VP.n47 VP.n46 12.234
R128 VP.n48 VP.n47 12.234
R129 VP.n76 VP.t3 10.2339
R130 VP.n13 VP.t9 10.2339
R131 VP.n104 VP.t1 10.2339
R132 VP.n118 VP.t4 10.2339
R133 VP.n131 VP.t8 10.2339
R134 VP.n74 VP.t6 10.2339
R135 VP.n61 VP.t5 10.2339
R136 VP.n47 VP.t0 10.2339
R137 VP.n31 VP.t7 10.2339
R138 VP.n91 VP.n13 2.93654
R139 VP.n118 VP.n117 2.93654
R140 VP.n61 VP.n60 2.93654
R141 VP.n34 VP.n31 2.93654
R142 VP.n33 VP.n32 2.75932
R143 VP.n75 VP.n18 0.417535
R144 VP.n78 VP.n77 0.417535
R145 VP.n132 VP.n0 0.417535
R146 VP VP.n132 0.394291
R147 VP.n33 VP.n30 0.189894
R148 VP.n37 VP.n30 0.189894
R149 VP.n38 VP.n37 0.189894
R150 VP.n39 VP.n38 0.189894
R151 VP.n39 VP.n28 0.189894
R152 VP.n43 VP.n28 0.189894
R153 VP.n44 VP.n43 0.189894
R154 VP.n45 VP.n44 0.189894
R155 VP.n45 VP.n26 0.189894
R156 VP.n50 VP.n26 0.189894
R157 VP.n51 VP.n50 0.189894
R158 VP.n52 VP.n51 0.189894
R159 VP.n52 VP.n24 0.189894
R160 VP.n56 VP.n24 0.189894
R161 VP.n57 VP.n56 0.189894
R162 VP.n58 VP.n57 0.189894
R163 VP.n58 VP.n22 0.189894
R164 VP.n63 VP.n22 0.189894
R165 VP.n64 VP.n63 0.189894
R166 VP.n65 VP.n64 0.189894
R167 VP.n65 VP.n20 0.189894
R168 VP.n69 VP.n20 0.189894
R169 VP.n70 VP.n69 0.189894
R170 VP.n71 VP.n70 0.189894
R171 VP.n71 VP.n18 0.189894
R172 VP.n79 VP.n78 0.189894
R173 VP.n79 VP.n16 0.189894
R174 VP.n83 VP.n16 0.189894
R175 VP.n84 VP.n83 0.189894
R176 VP.n85 VP.n84 0.189894
R177 VP.n85 VP.n14 0.189894
R178 VP.n89 VP.n14 0.189894
R179 VP.n90 VP.n89 0.189894
R180 VP.n90 VP.n12 0.189894
R181 VP.n94 VP.n12 0.189894
R182 VP.n95 VP.n94 0.189894
R183 VP.n96 VP.n95 0.189894
R184 VP.n96 VP.n10 0.189894
R185 VP.n100 VP.n10 0.189894
R186 VP.n101 VP.n100 0.189894
R187 VP.n102 VP.n101 0.189894
R188 VP.n102 VP.n8 0.189894
R189 VP.n107 VP.n8 0.189894
R190 VP.n108 VP.n107 0.189894
R191 VP.n109 VP.n108 0.189894
R192 VP.n109 VP.n6 0.189894
R193 VP.n113 VP.n6 0.189894
R194 VP.n114 VP.n113 0.189894
R195 VP.n115 VP.n114 0.189894
R196 VP.n115 VP.n4 0.189894
R197 VP.n120 VP.n4 0.189894
R198 VP.n121 VP.n120 0.189894
R199 VP.n122 VP.n121 0.189894
R200 VP.n122 VP.n2 0.189894
R201 VP.n126 VP.n2 0.189894
R202 VP.n127 VP.n126 0.189894
R203 VP.n128 VP.n127 0.189894
R204 VP.n128 VP.n0 0.189894
R205 VTAIL.n17 VTAIL.t3 252.861
R206 VTAIL.n2 VTAIL.t9 252.861
R207 VTAIL.n16 VTAIL.t13 252.861
R208 VTAIL.n11 VTAIL.t1 252.861
R209 VTAIL.n19 VTAIL.n18 233.626
R210 VTAIL.n1 VTAIL.n0 233.626
R211 VTAIL.n4 VTAIL.n3 233.626
R212 VTAIL.n6 VTAIL.n5 233.626
R213 VTAIL.n15 VTAIL.n14 233.626
R214 VTAIL.n13 VTAIL.n12 233.626
R215 VTAIL.n10 VTAIL.n9 233.626
R216 VTAIL.n8 VTAIL.n7 233.626
R217 VTAIL.n8 VTAIL.n6 21.2548
R218 VTAIL.n18 VTAIL.t7 19.2342
R219 VTAIL.n18 VTAIL.t0 19.2342
R220 VTAIL.n0 VTAIL.t6 19.2342
R221 VTAIL.n0 VTAIL.t19 19.2342
R222 VTAIL.n3 VTAIL.t10 19.2342
R223 VTAIL.n3 VTAIL.t8 19.2342
R224 VTAIL.n5 VTAIL.t11 19.2342
R225 VTAIL.n5 VTAIL.t15 19.2342
R226 VTAIL.n14 VTAIL.t12 19.2342
R227 VTAIL.n14 VTAIL.t14 19.2342
R228 VTAIL.n12 VTAIL.t17 19.2342
R229 VTAIL.n12 VTAIL.t16 19.2342
R230 VTAIL.n9 VTAIL.t5 19.2342
R231 VTAIL.n9 VTAIL.t2 19.2342
R232 VTAIL.n7 VTAIL.t4 19.2342
R233 VTAIL.n7 VTAIL.t18 19.2342
R234 VTAIL.n17 VTAIL.n16 17.5393
R235 VTAIL.n10 VTAIL.n8 3.71602
R236 VTAIL.n11 VTAIL.n10 3.71602
R237 VTAIL.n15 VTAIL.n13 3.71602
R238 VTAIL.n16 VTAIL.n15 3.71602
R239 VTAIL.n6 VTAIL.n4 3.71602
R240 VTAIL.n4 VTAIL.n2 3.71602
R241 VTAIL.n19 VTAIL.n17 3.71602
R242 VTAIL VTAIL.n1 2.84533
R243 VTAIL.n13 VTAIL.n11 2.32809
R244 VTAIL.n2 VTAIL.n1 2.32809
R245 VTAIL VTAIL.n19 0.87119
R246 VDD1.n3 VDD1.t6 273.255
R247 VDD1.n1 VDD1.t7 273.255
R248 VDD1.n5 VDD1.n4 253.036
R249 VDD1.n3 VDD1.n2 250.305
R250 VDD1.n7 VDD1.n6 250.305
R251 VDD1.n1 VDD1.n0 250.305
R252 VDD1.n7 VDD1.n5 45.2617
R253 VDD1.n6 VDD1.t4 19.2342
R254 VDD1.n6 VDD1.t3 19.2342
R255 VDD1.n0 VDD1.t2 19.2342
R256 VDD1.n0 VDD1.t9 19.2342
R257 VDD1.n4 VDD1.t5 19.2342
R258 VDD1.n4 VDD1.t1 19.2342
R259 VDD1.n2 VDD1.t0 19.2342
R260 VDD1.n2 VDD1.t8 19.2342
R261 VDD1 VDD1.n7 2.72895
R262 VDD1 VDD1.n1 0.987569
R263 VDD1.n5 VDD1.n3 0.874033
R264 VN.n113 VN.n58 161.3
R265 VN.n112 VN.n111 161.3
R266 VN.n110 VN.n59 161.3
R267 VN.n109 VN.n108 161.3
R268 VN.n107 VN.n60 161.3
R269 VN.n106 VN.n105 161.3
R270 VN.n104 VN.n61 161.3
R271 VN.n103 VN.n102 161.3
R272 VN.n100 VN.n62 161.3
R273 VN.n99 VN.n98 161.3
R274 VN.n97 VN.n63 161.3
R275 VN.n96 VN.n95 161.3
R276 VN.n94 VN.n64 161.3
R277 VN.n93 VN.n92 161.3
R278 VN.n91 VN.n65 161.3
R279 VN.n90 VN.n89 161.3
R280 VN.n88 VN.n66 161.3
R281 VN.n86 VN.n85 161.3
R282 VN.n84 VN.n67 161.3
R283 VN.n83 VN.n82 161.3
R284 VN.n81 VN.n68 161.3
R285 VN.n80 VN.n79 161.3
R286 VN.n78 VN.n69 161.3
R287 VN.n77 VN.n76 161.3
R288 VN.n75 VN.n70 161.3
R289 VN.n74 VN.n73 161.3
R290 VN.n55 VN.n0 161.3
R291 VN.n54 VN.n53 161.3
R292 VN.n52 VN.n1 161.3
R293 VN.n51 VN.n50 161.3
R294 VN.n49 VN.n2 161.3
R295 VN.n48 VN.n47 161.3
R296 VN.n46 VN.n3 161.3
R297 VN.n45 VN.n44 161.3
R298 VN.n42 VN.n4 161.3
R299 VN.n41 VN.n40 161.3
R300 VN.n39 VN.n5 161.3
R301 VN.n38 VN.n37 161.3
R302 VN.n36 VN.n6 161.3
R303 VN.n35 VN.n34 161.3
R304 VN.n33 VN.n7 161.3
R305 VN.n32 VN.n31 161.3
R306 VN.n30 VN.n8 161.3
R307 VN.n28 VN.n27 161.3
R308 VN.n26 VN.n9 161.3
R309 VN.n25 VN.n24 161.3
R310 VN.n23 VN.n10 161.3
R311 VN.n22 VN.n21 161.3
R312 VN.n20 VN.n11 161.3
R313 VN.n19 VN.n18 161.3
R314 VN.n17 VN.n12 161.3
R315 VN.n16 VN.n15 161.3
R316 VN.n14 VN.n13 72.0574
R317 VN.n72 VN.n71 72.0574
R318 VN.n57 VN.n56 64.0762
R319 VN.n115 VN.n114 64.0762
R320 VN.n50 VN.n49 56.5193
R321 VN.n108 VN.n107 56.5193
R322 VN VN.n115 53.0534
R323 VN.n23 VN.n22 49.7204
R324 VN.n36 VN.n35 49.7204
R325 VN.n81 VN.n80 49.7204
R326 VN.n94 VN.n93 49.7204
R327 VN.n14 VN.t9 42.5534
R328 VN.n72 VN.t3 42.5534
R329 VN.n22 VN.n11 31.2664
R330 VN.n37 VN.n36 31.2664
R331 VN.n80 VN.n69 31.2664
R332 VN.n95 VN.n94 31.2664
R333 VN.n17 VN.n16 24.4675
R334 VN.n18 VN.n17 24.4675
R335 VN.n18 VN.n11 24.4675
R336 VN.n24 VN.n23 24.4675
R337 VN.n24 VN.n9 24.4675
R338 VN.n28 VN.n9 24.4675
R339 VN.n31 VN.n30 24.4675
R340 VN.n31 VN.n7 24.4675
R341 VN.n35 VN.n7 24.4675
R342 VN.n37 VN.n5 24.4675
R343 VN.n41 VN.n5 24.4675
R344 VN.n42 VN.n41 24.4675
R345 VN.n44 VN.n3 24.4675
R346 VN.n48 VN.n3 24.4675
R347 VN.n49 VN.n48 24.4675
R348 VN.n50 VN.n1 24.4675
R349 VN.n54 VN.n1 24.4675
R350 VN.n55 VN.n54 24.4675
R351 VN.n76 VN.n69 24.4675
R352 VN.n76 VN.n75 24.4675
R353 VN.n75 VN.n74 24.4675
R354 VN.n93 VN.n65 24.4675
R355 VN.n89 VN.n65 24.4675
R356 VN.n89 VN.n88 24.4675
R357 VN.n86 VN.n67 24.4675
R358 VN.n82 VN.n67 24.4675
R359 VN.n82 VN.n81 24.4675
R360 VN.n107 VN.n106 24.4675
R361 VN.n106 VN.n61 24.4675
R362 VN.n102 VN.n61 24.4675
R363 VN.n100 VN.n99 24.4675
R364 VN.n99 VN.n63 24.4675
R365 VN.n95 VN.n63 24.4675
R366 VN.n113 VN.n112 24.4675
R367 VN.n112 VN.n59 24.4675
R368 VN.n108 VN.n59 24.4675
R369 VN.n44 VN.n43 21.5315
R370 VN.n102 VN.n101 21.5315
R371 VN.n56 VN.n55 18.1061
R372 VN.n114 VN.n113 18.1061
R373 VN.n29 VN.n28 12.234
R374 VN.n30 VN.n29 12.234
R375 VN.n88 VN.n87 12.234
R376 VN.n87 VN.n86 12.234
R377 VN.n13 VN.t6 10.2339
R378 VN.n29 VN.t8 10.2339
R379 VN.n43 VN.t4 10.2339
R380 VN.n56 VN.t7 10.2339
R381 VN.n71 VN.t1 10.2339
R382 VN.n87 VN.t5 10.2339
R383 VN.n101 VN.t0 10.2339
R384 VN.n114 VN.t2 10.2339
R385 VN.n16 VN.n13 2.93654
R386 VN.n43 VN.n42 2.93654
R387 VN.n74 VN.n71 2.93654
R388 VN.n101 VN.n100 2.93654
R389 VN.n73 VN.n72 2.75934
R390 VN.n15 VN.n14 2.75934
R391 VN.n115 VN.n58 0.417535
R392 VN.n57 VN.n0 0.417535
R393 VN VN.n57 0.394291
R394 VN.n111 VN.n58 0.189894
R395 VN.n111 VN.n110 0.189894
R396 VN.n110 VN.n109 0.189894
R397 VN.n109 VN.n60 0.189894
R398 VN.n105 VN.n60 0.189894
R399 VN.n105 VN.n104 0.189894
R400 VN.n104 VN.n103 0.189894
R401 VN.n103 VN.n62 0.189894
R402 VN.n98 VN.n62 0.189894
R403 VN.n98 VN.n97 0.189894
R404 VN.n97 VN.n96 0.189894
R405 VN.n96 VN.n64 0.189894
R406 VN.n92 VN.n64 0.189894
R407 VN.n92 VN.n91 0.189894
R408 VN.n91 VN.n90 0.189894
R409 VN.n90 VN.n66 0.189894
R410 VN.n85 VN.n66 0.189894
R411 VN.n85 VN.n84 0.189894
R412 VN.n84 VN.n83 0.189894
R413 VN.n83 VN.n68 0.189894
R414 VN.n79 VN.n68 0.189894
R415 VN.n79 VN.n78 0.189894
R416 VN.n78 VN.n77 0.189894
R417 VN.n77 VN.n70 0.189894
R418 VN.n73 VN.n70 0.189894
R419 VN.n15 VN.n12 0.189894
R420 VN.n19 VN.n12 0.189894
R421 VN.n20 VN.n19 0.189894
R422 VN.n21 VN.n20 0.189894
R423 VN.n21 VN.n10 0.189894
R424 VN.n25 VN.n10 0.189894
R425 VN.n26 VN.n25 0.189894
R426 VN.n27 VN.n26 0.189894
R427 VN.n27 VN.n8 0.189894
R428 VN.n32 VN.n8 0.189894
R429 VN.n33 VN.n32 0.189894
R430 VN.n34 VN.n33 0.189894
R431 VN.n34 VN.n6 0.189894
R432 VN.n38 VN.n6 0.189894
R433 VN.n39 VN.n38 0.189894
R434 VN.n40 VN.n39 0.189894
R435 VN.n40 VN.n4 0.189894
R436 VN.n45 VN.n4 0.189894
R437 VN.n46 VN.n45 0.189894
R438 VN.n47 VN.n46 0.189894
R439 VN.n47 VN.n2 0.189894
R440 VN.n51 VN.n2 0.189894
R441 VN.n52 VN.n51 0.189894
R442 VN.n53 VN.n52 0.189894
R443 VN.n53 VN.n0 0.189894
R444 VDD2.n1 VDD2.t0 273.255
R445 VDD2.n4 VDD2.t7 269.539
R446 VDD2.n3 VDD2.n2 253.036
R447 VDD2 VDD2.n7 253.034
R448 VDD2.n1 VDD2.n0 250.305
R449 VDD2.n6 VDD2.n5 250.305
R450 VDD2.n4 VDD2.n3 42.8209
R451 VDD2.n7 VDD2.t8 19.2342
R452 VDD2.n7 VDD2.t6 19.2342
R453 VDD2.n5 VDD2.t9 19.2342
R454 VDD2.n5 VDD2.t4 19.2342
R455 VDD2.n2 VDD2.t5 19.2342
R456 VDD2.n2 VDD2.t2 19.2342
R457 VDD2.n0 VDD2.t3 19.2342
R458 VDD2.n0 VDD2.t1 19.2342
R459 VDD2.n6 VDD2.n4 3.71602
R460 VDD2 VDD2.n6 0.987569
R461 VDD2.n3 VDD2.n1 0.874033
R462 B.n640 B.n639 585
R463 B.n641 B.n64 585
R464 B.n643 B.n642 585
R465 B.n644 B.n63 585
R466 B.n646 B.n645 585
R467 B.n647 B.n62 585
R468 B.n649 B.n648 585
R469 B.n650 B.n61 585
R470 B.n652 B.n651 585
R471 B.n653 B.n57 585
R472 B.n655 B.n654 585
R473 B.n656 B.n56 585
R474 B.n658 B.n657 585
R475 B.n659 B.n55 585
R476 B.n661 B.n660 585
R477 B.n662 B.n54 585
R478 B.n664 B.n663 585
R479 B.n665 B.n53 585
R480 B.n667 B.n666 585
R481 B.n668 B.n52 585
R482 B.n670 B.n669 585
R483 B.n672 B.n49 585
R484 B.n674 B.n673 585
R485 B.n675 B.n48 585
R486 B.n677 B.n676 585
R487 B.n678 B.n47 585
R488 B.n680 B.n679 585
R489 B.n681 B.n46 585
R490 B.n683 B.n682 585
R491 B.n684 B.n45 585
R492 B.n686 B.n685 585
R493 B.n687 B.n44 585
R494 B.n638 B.n65 585
R495 B.n637 B.n636 585
R496 B.n635 B.n66 585
R497 B.n634 B.n633 585
R498 B.n632 B.n67 585
R499 B.n631 B.n630 585
R500 B.n629 B.n68 585
R501 B.n628 B.n627 585
R502 B.n626 B.n69 585
R503 B.n625 B.n624 585
R504 B.n623 B.n70 585
R505 B.n622 B.n621 585
R506 B.n620 B.n71 585
R507 B.n619 B.n618 585
R508 B.n617 B.n72 585
R509 B.n616 B.n615 585
R510 B.n614 B.n73 585
R511 B.n613 B.n612 585
R512 B.n611 B.n74 585
R513 B.n610 B.n609 585
R514 B.n608 B.n75 585
R515 B.n607 B.n606 585
R516 B.n605 B.n76 585
R517 B.n604 B.n603 585
R518 B.n602 B.n77 585
R519 B.n601 B.n600 585
R520 B.n599 B.n78 585
R521 B.n598 B.n597 585
R522 B.n596 B.n79 585
R523 B.n595 B.n594 585
R524 B.n593 B.n80 585
R525 B.n592 B.n591 585
R526 B.n590 B.n81 585
R527 B.n589 B.n588 585
R528 B.n587 B.n82 585
R529 B.n586 B.n585 585
R530 B.n584 B.n83 585
R531 B.n583 B.n582 585
R532 B.n581 B.n84 585
R533 B.n580 B.n579 585
R534 B.n578 B.n85 585
R535 B.n577 B.n576 585
R536 B.n575 B.n86 585
R537 B.n574 B.n573 585
R538 B.n572 B.n87 585
R539 B.n571 B.n570 585
R540 B.n569 B.n88 585
R541 B.n568 B.n567 585
R542 B.n566 B.n89 585
R543 B.n565 B.n564 585
R544 B.n563 B.n90 585
R545 B.n562 B.n561 585
R546 B.n560 B.n91 585
R547 B.n559 B.n558 585
R548 B.n557 B.n92 585
R549 B.n556 B.n555 585
R550 B.n554 B.n93 585
R551 B.n553 B.n552 585
R552 B.n551 B.n94 585
R553 B.n550 B.n549 585
R554 B.n548 B.n95 585
R555 B.n547 B.n546 585
R556 B.n545 B.n96 585
R557 B.n544 B.n543 585
R558 B.n542 B.n97 585
R559 B.n541 B.n540 585
R560 B.n539 B.n98 585
R561 B.n538 B.n537 585
R562 B.n536 B.n99 585
R563 B.n535 B.n534 585
R564 B.n533 B.n100 585
R565 B.n532 B.n531 585
R566 B.n530 B.n101 585
R567 B.n529 B.n528 585
R568 B.n527 B.n102 585
R569 B.n526 B.n525 585
R570 B.n524 B.n103 585
R571 B.n523 B.n522 585
R572 B.n521 B.n104 585
R573 B.n520 B.n519 585
R574 B.n518 B.n105 585
R575 B.n517 B.n516 585
R576 B.n515 B.n106 585
R577 B.n514 B.n513 585
R578 B.n512 B.n107 585
R579 B.n511 B.n510 585
R580 B.n509 B.n108 585
R581 B.n508 B.n507 585
R582 B.n506 B.n109 585
R583 B.n505 B.n504 585
R584 B.n503 B.n110 585
R585 B.n502 B.n501 585
R586 B.n500 B.n111 585
R587 B.n499 B.n498 585
R588 B.n497 B.n112 585
R589 B.n496 B.n495 585
R590 B.n494 B.n113 585
R591 B.n493 B.n492 585
R592 B.n491 B.n114 585
R593 B.n490 B.n489 585
R594 B.n488 B.n115 585
R595 B.n487 B.n486 585
R596 B.n485 B.n116 585
R597 B.n484 B.n483 585
R598 B.n482 B.n117 585
R599 B.n481 B.n480 585
R600 B.n479 B.n118 585
R601 B.n478 B.n477 585
R602 B.n476 B.n119 585
R603 B.n475 B.n474 585
R604 B.n473 B.n120 585
R605 B.n472 B.n471 585
R606 B.n470 B.n121 585
R607 B.n469 B.n468 585
R608 B.n467 B.n122 585
R609 B.n466 B.n465 585
R610 B.n464 B.n123 585
R611 B.n463 B.n462 585
R612 B.n461 B.n124 585
R613 B.n460 B.n459 585
R614 B.n458 B.n125 585
R615 B.n457 B.n456 585
R616 B.n455 B.n126 585
R617 B.n454 B.n453 585
R618 B.n452 B.n127 585
R619 B.n451 B.n450 585
R620 B.n449 B.n128 585
R621 B.n448 B.n447 585
R622 B.n446 B.n129 585
R623 B.n445 B.n444 585
R624 B.n443 B.n130 585
R625 B.n442 B.n441 585
R626 B.n440 B.n131 585
R627 B.n439 B.n438 585
R628 B.n437 B.n132 585
R629 B.n436 B.n435 585
R630 B.n434 B.n133 585
R631 B.n433 B.n432 585
R632 B.n431 B.n134 585
R633 B.n430 B.n429 585
R634 B.n428 B.n135 585
R635 B.n427 B.n426 585
R636 B.n425 B.n136 585
R637 B.n424 B.n423 585
R638 B.n422 B.n137 585
R639 B.n421 B.n420 585
R640 B.n419 B.n138 585
R641 B.n418 B.n417 585
R642 B.n416 B.n139 585
R643 B.n415 B.n414 585
R644 B.n413 B.n140 585
R645 B.n412 B.n411 585
R646 B.n410 B.n141 585
R647 B.n409 B.n408 585
R648 B.n407 B.n142 585
R649 B.n406 B.n405 585
R650 B.n404 B.n143 585
R651 B.n403 B.n402 585
R652 B.n401 B.n144 585
R653 B.n400 B.n399 585
R654 B.n398 B.n145 585
R655 B.n397 B.n396 585
R656 B.n395 B.n146 585
R657 B.n394 B.n393 585
R658 B.n392 B.n147 585
R659 B.n391 B.n390 585
R660 B.n389 B.n148 585
R661 B.n388 B.n387 585
R662 B.n386 B.n149 585
R663 B.n337 B.n336 585
R664 B.n338 B.n169 585
R665 B.n340 B.n339 585
R666 B.n341 B.n168 585
R667 B.n343 B.n342 585
R668 B.n344 B.n167 585
R669 B.n346 B.n345 585
R670 B.n347 B.n166 585
R671 B.n349 B.n348 585
R672 B.n350 B.n165 585
R673 B.n352 B.n351 585
R674 B.n354 B.n162 585
R675 B.n356 B.n355 585
R676 B.n357 B.n161 585
R677 B.n359 B.n358 585
R678 B.n360 B.n160 585
R679 B.n362 B.n361 585
R680 B.n363 B.n159 585
R681 B.n365 B.n364 585
R682 B.n366 B.n158 585
R683 B.n368 B.n367 585
R684 B.n370 B.n369 585
R685 B.n371 B.n154 585
R686 B.n373 B.n372 585
R687 B.n374 B.n153 585
R688 B.n376 B.n375 585
R689 B.n377 B.n152 585
R690 B.n379 B.n378 585
R691 B.n380 B.n151 585
R692 B.n382 B.n381 585
R693 B.n383 B.n150 585
R694 B.n385 B.n384 585
R695 B.n335 B.n170 585
R696 B.n334 B.n333 585
R697 B.n332 B.n171 585
R698 B.n331 B.n330 585
R699 B.n329 B.n172 585
R700 B.n328 B.n327 585
R701 B.n326 B.n173 585
R702 B.n325 B.n324 585
R703 B.n323 B.n174 585
R704 B.n322 B.n321 585
R705 B.n320 B.n175 585
R706 B.n319 B.n318 585
R707 B.n317 B.n176 585
R708 B.n316 B.n315 585
R709 B.n314 B.n177 585
R710 B.n313 B.n312 585
R711 B.n311 B.n178 585
R712 B.n310 B.n309 585
R713 B.n308 B.n179 585
R714 B.n307 B.n306 585
R715 B.n305 B.n180 585
R716 B.n304 B.n303 585
R717 B.n302 B.n181 585
R718 B.n301 B.n300 585
R719 B.n299 B.n182 585
R720 B.n298 B.n297 585
R721 B.n296 B.n183 585
R722 B.n295 B.n294 585
R723 B.n293 B.n184 585
R724 B.n292 B.n291 585
R725 B.n290 B.n185 585
R726 B.n289 B.n288 585
R727 B.n287 B.n186 585
R728 B.n286 B.n285 585
R729 B.n284 B.n187 585
R730 B.n283 B.n282 585
R731 B.n281 B.n188 585
R732 B.n280 B.n279 585
R733 B.n278 B.n189 585
R734 B.n277 B.n276 585
R735 B.n275 B.n190 585
R736 B.n274 B.n273 585
R737 B.n272 B.n191 585
R738 B.n271 B.n270 585
R739 B.n269 B.n192 585
R740 B.n268 B.n267 585
R741 B.n266 B.n193 585
R742 B.n265 B.n264 585
R743 B.n263 B.n194 585
R744 B.n262 B.n261 585
R745 B.n260 B.n195 585
R746 B.n259 B.n258 585
R747 B.n257 B.n196 585
R748 B.n256 B.n255 585
R749 B.n254 B.n197 585
R750 B.n253 B.n252 585
R751 B.n251 B.n198 585
R752 B.n250 B.n249 585
R753 B.n248 B.n199 585
R754 B.n247 B.n246 585
R755 B.n245 B.n200 585
R756 B.n244 B.n243 585
R757 B.n242 B.n201 585
R758 B.n241 B.n240 585
R759 B.n239 B.n202 585
R760 B.n238 B.n237 585
R761 B.n236 B.n203 585
R762 B.n235 B.n234 585
R763 B.n233 B.n204 585
R764 B.n232 B.n231 585
R765 B.n230 B.n205 585
R766 B.n229 B.n228 585
R767 B.n227 B.n206 585
R768 B.n226 B.n225 585
R769 B.n224 B.n207 585
R770 B.n223 B.n222 585
R771 B.n221 B.n208 585
R772 B.n220 B.n219 585
R773 B.n218 B.n209 585
R774 B.n217 B.n216 585
R775 B.n215 B.n210 585
R776 B.n214 B.n213 585
R777 B.n212 B.n211 585
R778 B.n2 B.n0 585
R779 B.n813 B.n1 585
R780 B.n812 B.n811 585
R781 B.n810 B.n3 585
R782 B.n809 B.n808 585
R783 B.n807 B.n4 585
R784 B.n806 B.n805 585
R785 B.n804 B.n5 585
R786 B.n803 B.n802 585
R787 B.n801 B.n6 585
R788 B.n800 B.n799 585
R789 B.n798 B.n7 585
R790 B.n797 B.n796 585
R791 B.n795 B.n8 585
R792 B.n794 B.n793 585
R793 B.n792 B.n9 585
R794 B.n791 B.n790 585
R795 B.n789 B.n10 585
R796 B.n788 B.n787 585
R797 B.n786 B.n11 585
R798 B.n785 B.n784 585
R799 B.n783 B.n12 585
R800 B.n782 B.n781 585
R801 B.n780 B.n13 585
R802 B.n779 B.n778 585
R803 B.n777 B.n14 585
R804 B.n776 B.n775 585
R805 B.n774 B.n15 585
R806 B.n773 B.n772 585
R807 B.n771 B.n16 585
R808 B.n770 B.n769 585
R809 B.n768 B.n17 585
R810 B.n767 B.n766 585
R811 B.n765 B.n18 585
R812 B.n764 B.n763 585
R813 B.n762 B.n19 585
R814 B.n761 B.n760 585
R815 B.n759 B.n20 585
R816 B.n758 B.n757 585
R817 B.n756 B.n21 585
R818 B.n755 B.n754 585
R819 B.n753 B.n22 585
R820 B.n752 B.n751 585
R821 B.n750 B.n23 585
R822 B.n749 B.n748 585
R823 B.n747 B.n24 585
R824 B.n746 B.n745 585
R825 B.n744 B.n25 585
R826 B.n743 B.n742 585
R827 B.n741 B.n26 585
R828 B.n740 B.n739 585
R829 B.n738 B.n27 585
R830 B.n737 B.n736 585
R831 B.n735 B.n28 585
R832 B.n734 B.n733 585
R833 B.n732 B.n29 585
R834 B.n731 B.n730 585
R835 B.n729 B.n30 585
R836 B.n728 B.n727 585
R837 B.n726 B.n31 585
R838 B.n725 B.n724 585
R839 B.n723 B.n32 585
R840 B.n722 B.n721 585
R841 B.n720 B.n33 585
R842 B.n719 B.n718 585
R843 B.n717 B.n34 585
R844 B.n716 B.n715 585
R845 B.n714 B.n35 585
R846 B.n713 B.n712 585
R847 B.n711 B.n36 585
R848 B.n710 B.n709 585
R849 B.n708 B.n37 585
R850 B.n707 B.n706 585
R851 B.n705 B.n38 585
R852 B.n704 B.n703 585
R853 B.n702 B.n39 585
R854 B.n701 B.n700 585
R855 B.n699 B.n40 585
R856 B.n698 B.n697 585
R857 B.n696 B.n41 585
R858 B.n695 B.n694 585
R859 B.n693 B.n42 585
R860 B.n692 B.n691 585
R861 B.n690 B.n43 585
R862 B.n689 B.n688 585
R863 B.n815 B.n814 585
R864 B.n337 B.n170 540.549
R865 B.n688 B.n687 540.549
R866 B.n386 B.n385 540.549
R867 B.n639 B.n638 540.549
R868 B.n155 B.t8 334.284
R869 B.n58 B.t1 334.284
R870 B.n163 B.t11 334.284
R871 B.n50 B.t4 334.284
R872 B.n156 B.t7 250.696
R873 B.n59 B.t2 250.696
R874 B.n164 B.t10 250.696
R875 B.n51 B.t5 250.696
R876 B.n155 B.t6 209.875
R877 B.n163 B.t9 209.875
R878 B.n50 B.t3 209.875
R879 B.n58 B.t0 209.875
R880 B.n333 B.n170 163.367
R881 B.n333 B.n332 163.367
R882 B.n332 B.n331 163.367
R883 B.n331 B.n172 163.367
R884 B.n327 B.n172 163.367
R885 B.n327 B.n326 163.367
R886 B.n326 B.n325 163.367
R887 B.n325 B.n174 163.367
R888 B.n321 B.n174 163.367
R889 B.n321 B.n320 163.367
R890 B.n320 B.n319 163.367
R891 B.n319 B.n176 163.367
R892 B.n315 B.n176 163.367
R893 B.n315 B.n314 163.367
R894 B.n314 B.n313 163.367
R895 B.n313 B.n178 163.367
R896 B.n309 B.n178 163.367
R897 B.n309 B.n308 163.367
R898 B.n308 B.n307 163.367
R899 B.n307 B.n180 163.367
R900 B.n303 B.n180 163.367
R901 B.n303 B.n302 163.367
R902 B.n302 B.n301 163.367
R903 B.n301 B.n182 163.367
R904 B.n297 B.n182 163.367
R905 B.n297 B.n296 163.367
R906 B.n296 B.n295 163.367
R907 B.n295 B.n184 163.367
R908 B.n291 B.n184 163.367
R909 B.n291 B.n290 163.367
R910 B.n290 B.n289 163.367
R911 B.n289 B.n186 163.367
R912 B.n285 B.n186 163.367
R913 B.n285 B.n284 163.367
R914 B.n284 B.n283 163.367
R915 B.n283 B.n188 163.367
R916 B.n279 B.n188 163.367
R917 B.n279 B.n278 163.367
R918 B.n278 B.n277 163.367
R919 B.n277 B.n190 163.367
R920 B.n273 B.n190 163.367
R921 B.n273 B.n272 163.367
R922 B.n272 B.n271 163.367
R923 B.n271 B.n192 163.367
R924 B.n267 B.n192 163.367
R925 B.n267 B.n266 163.367
R926 B.n266 B.n265 163.367
R927 B.n265 B.n194 163.367
R928 B.n261 B.n194 163.367
R929 B.n261 B.n260 163.367
R930 B.n260 B.n259 163.367
R931 B.n259 B.n196 163.367
R932 B.n255 B.n196 163.367
R933 B.n255 B.n254 163.367
R934 B.n254 B.n253 163.367
R935 B.n253 B.n198 163.367
R936 B.n249 B.n198 163.367
R937 B.n249 B.n248 163.367
R938 B.n248 B.n247 163.367
R939 B.n247 B.n200 163.367
R940 B.n243 B.n200 163.367
R941 B.n243 B.n242 163.367
R942 B.n242 B.n241 163.367
R943 B.n241 B.n202 163.367
R944 B.n237 B.n202 163.367
R945 B.n237 B.n236 163.367
R946 B.n236 B.n235 163.367
R947 B.n235 B.n204 163.367
R948 B.n231 B.n204 163.367
R949 B.n231 B.n230 163.367
R950 B.n230 B.n229 163.367
R951 B.n229 B.n206 163.367
R952 B.n225 B.n206 163.367
R953 B.n225 B.n224 163.367
R954 B.n224 B.n223 163.367
R955 B.n223 B.n208 163.367
R956 B.n219 B.n208 163.367
R957 B.n219 B.n218 163.367
R958 B.n218 B.n217 163.367
R959 B.n217 B.n210 163.367
R960 B.n213 B.n210 163.367
R961 B.n213 B.n212 163.367
R962 B.n212 B.n2 163.367
R963 B.n814 B.n2 163.367
R964 B.n814 B.n813 163.367
R965 B.n813 B.n812 163.367
R966 B.n812 B.n3 163.367
R967 B.n808 B.n3 163.367
R968 B.n808 B.n807 163.367
R969 B.n807 B.n806 163.367
R970 B.n806 B.n5 163.367
R971 B.n802 B.n5 163.367
R972 B.n802 B.n801 163.367
R973 B.n801 B.n800 163.367
R974 B.n800 B.n7 163.367
R975 B.n796 B.n7 163.367
R976 B.n796 B.n795 163.367
R977 B.n795 B.n794 163.367
R978 B.n794 B.n9 163.367
R979 B.n790 B.n9 163.367
R980 B.n790 B.n789 163.367
R981 B.n789 B.n788 163.367
R982 B.n788 B.n11 163.367
R983 B.n784 B.n11 163.367
R984 B.n784 B.n783 163.367
R985 B.n783 B.n782 163.367
R986 B.n782 B.n13 163.367
R987 B.n778 B.n13 163.367
R988 B.n778 B.n777 163.367
R989 B.n777 B.n776 163.367
R990 B.n776 B.n15 163.367
R991 B.n772 B.n15 163.367
R992 B.n772 B.n771 163.367
R993 B.n771 B.n770 163.367
R994 B.n770 B.n17 163.367
R995 B.n766 B.n17 163.367
R996 B.n766 B.n765 163.367
R997 B.n765 B.n764 163.367
R998 B.n764 B.n19 163.367
R999 B.n760 B.n19 163.367
R1000 B.n760 B.n759 163.367
R1001 B.n759 B.n758 163.367
R1002 B.n758 B.n21 163.367
R1003 B.n754 B.n21 163.367
R1004 B.n754 B.n753 163.367
R1005 B.n753 B.n752 163.367
R1006 B.n752 B.n23 163.367
R1007 B.n748 B.n23 163.367
R1008 B.n748 B.n747 163.367
R1009 B.n747 B.n746 163.367
R1010 B.n746 B.n25 163.367
R1011 B.n742 B.n25 163.367
R1012 B.n742 B.n741 163.367
R1013 B.n741 B.n740 163.367
R1014 B.n740 B.n27 163.367
R1015 B.n736 B.n27 163.367
R1016 B.n736 B.n735 163.367
R1017 B.n735 B.n734 163.367
R1018 B.n734 B.n29 163.367
R1019 B.n730 B.n29 163.367
R1020 B.n730 B.n729 163.367
R1021 B.n729 B.n728 163.367
R1022 B.n728 B.n31 163.367
R1023 B.n724 B.n31 163.367
R1024 B.n724 B.n723 163.367
R1025 B.n723 B.n722 163.367
R1026 B.n722 B.n33 163.367
R1027 B.n718 B.n33 163.367
R1028 B.n718 B.n717 163.367
R1029 B.n717 B.n716 163.367
R1030 B.n716 B.n35 163.367
R1031 B.n712 B.n35 163.367
R1032 B.n712 B.n711 163.367
R1033 B.n711 B.n710 163.367
R1034 B.n710 B.n37 163.367
R1035 B.n706 B.n37 163.367
R1036 B.n706 B.n705 163.367
R1037 B.n705 B.n704 163.367
R1038 B.n704 B.n39 163.367
R1039 B.n700 B.n39 163.367
R1040 B.n700 B.n699 163.367
R1041 B.n699 B.n698 163.367
R1042 B.n698 B.n41 163.367
R1043 B.n694 B.n41 163.367
R1044 B.n694 B.n693 163.367
R1045 B.n693 B.n692 163.367
R1046 B.n692 B.n43 163.367
R1047 B.n688 B.n43 163.367
R1048 B.n338 B.n337 163.367
R1049 B.n339 B.n338 163.367
R1050 B.n339 B.n168 163.367
R1051 B.n343 B.n168 163.367
R1052 B.n344 B.n343 163.367
R1053 B.n345 B.n344 163.367
R1054 B.n345 B.n166 163.367
R1055 B.n349 B.n166 163.367
R1056 B.n350 B.n349 163.367
R1057 B.n351 B.n350 163.367
R1058 B.n351 B.n162 163.367
R1059 B.n356 B.n162 163.367
R1060 B.n357 B.n356 163.367
R1061 B.n358 B.n357 163.367
R1062 B.n358 B.n160 163.367
R1063 B.n362 B.n160 163.367
R1064 B.n363 B.n362 163.367
R1065 B.n364 B.n363 163.367
R1066 B.n364 B.n158 163.367
R1067 B.n368 B.n158 163.367
R1068 B.n369 B.n368 163.367
R1069 B.n369 B.n154 163.367
R1070 B.n373 B.n154 163.367
R1071 B.n374 B.n373 163.367
R1072 B.n375 B.n374 163.367
R1073 B.n375 B.n152 163.367
R1074 B.n379 B.n152 163.367
R1075 B.n380 B.n379 163.367
R1076 B.n381 B.n380 163.367
R1077 B.n381 B.n150 163.367
R1078 B.n385 B.n150 163.367
R1079 B.n387 B.n386 163.367
R1080 B.n387 B.n148 163.367
R1081 B.n391 B.n148 163.367
R1082 B.n392 B.n391 163.367
R1083 B.n393 B.n392 163.367
R1084 B.n393 B.n146 163.367
R1085 B.n397 B.n146 163.367
R1086 B.n398 B.n397 163.367
R1087 B.n399 B.n398 163.367
R1088 B.n399 B.n144 163.367
R1089 B.n403 B.n144 163.367
R1090 B.n404 B.n403 163.367
R1091 B.n405 B.n404 163.367
R1092 B.n405 B.n142 163.367
R1093 B.n409 B.n142 163.367
R1094 B.n410 B.n409 163.367
R1095 B.n411 B.n410 163.367
R1096 B.n411 B.n140 163.367
R1097 B.n415 B.n140 163.367
R1098 B.n416 B.n415 163.367
R1099 B.n417 B.n416 163.367
R1100 B.n417 B.n138 163.367
R1101 B.n421 B.n138 163.367
R1102 B.n422 B.n421 163.367
R1103 B.n423 B.n422 163.367
R1104 B.n423 B.n136 163.367
R1105 B.n427 B.n136 163.367
R1106 B.n428 B.n427 163.367
R1107 B.n429 B.n428 163.367
R1108 B.n429 B.n134 163.367
R1109 B.n433 B.n134 163.367
R1110 B.n434 B.n433 163.367
R1111 B.n435 B.n434 163.367
R1112 B.n435 B.n132 163.367
R1113 B.n439 B.n132 163.367
R1114 B.n440 B.n439 163.367
R1115 B.n441 B.n440 163.367
R1116 B.n441 B.n130 163.367
R1117 B.n445 B.n130 163.367
R1118 B.n446 B.n445 163.367
R1119 B.n447 B.n446 163.367
R1120 B.n447 B.n128 163.367
R1121 B.n451 B.n128 163.367
R1122 B.n452 B.n451 163.367
R1123 B.n453 B.n452 163.367
R1124 B.n453 B.n126 163.367
R1125 B.n457 B.n126 163.367
R1126 B.n458 B.n457 163.367
R1127 B.n459 B.n458 163.367
R1128 B.n459 B.n124 163.367
R1129 B.n463 B.n124 163.367
R1130 B.n464 B.n463 163.367
R1131 B.n465 B.n464 163.367
R1132 B.n465 B.n122 163.367
R1133 B.n469 B.n122 163.367
R1134 B.n470 B.n469 163.367
R1135 B.n471 B.n470 163.367
R1136 B.n471 B.n120 163.367
R1137 B.n475 B.n120 163.367
R1138 B.n476 B.n475 163.367
R1139 B.n477 B.n476 163.367
R1140 B.n477 B.n118 163.367
R1141 B.n481 B.n118 163.367
R1142 B.n482 B.n481 163.367
R1143 B.n483 B.n482 163.367
R1144 B.n483 B.n116 163.367
R1145 B.n487 B.n116 163.367
R1146 B.n488 B.n487 163.367
R1147 B.n489 B.n488 163.367
R1148 B.n489 B.n114 163.367
R1149 B.n493 B.n114 163.367
R1150 B.n494 B.n493 163.367
R1151 B.n495 B.n494 163.367
R1152 B.n495 B.n112 163.367
R1153 B.n499 B.n112 163.367
R1154 B.n500 B.n499 163.367
R1155 B.n501 B.n500 163.367
R1156 B.n501 B.n110 163.367
R1157 B.n505 B.n110 163.367
R1158 B.n506 B.n505 163.367
R1159 B.n507 B.n506 163.367
R1160 B.n507 B.n108 163.367
R1161 B.n511 B.n108 163.367
R1162 B.n512 B.n511 163.367
R1163 B.n513 B.n512 163.367
R1164 B.n513 B.n106 163.367
R1165 B.n517 B.n106 163.367
R1166 B.n518 B.n517 163.367
R1167 B.n519 B.n518 163.367
R1168 B.n519 B.n104 163.367
R1169 B.n523 B.n104 163.367
R1170 B.n524 B.n523 163.367
R1171 B.n525 B.n524 163.367
R1172 B.n525 B.n102 163.367
R1173 B.n529 B.n102 163.367
R1174 B.n530 B.n529 163.367
R1175 B.n531 B.n530 163.367
R1176 B.n531 B.n100 163.367
R1177 B.n535 B.n100 163.367
R1178 B.n536 B.n535 163.367
R1179 B.n537 B.n536 163.367
R1180 B.n537 B.n98 163.367
R1181 B.n541 B.n98 163.367
R1182 B.n542 B.n541 163.367
R1183 B.n543 B.n542 163.367
R1184 B.n543 B.n96 163.367
R1185 B.n547 B.n96 163.367
R1186 B.n548 B.n547 163.367
R1187 B.n549 B.n548 163.367
R1188 B.n549 B.n94 163.367
R1189 B.n553 B.n94 163.367
R1190 B.n554 B.n553 163.367
R1191 B.n555 B.n554 163.367
R1192 B.n555 B.n92 163.367
R1193 B.n559 B.n92 163.367
R1194 B.n560 B.n559 163.367
R1195 B.n561 B.n560 163.367
R1196 B.n561 B.n90 163.367
R1197 B.n565 B.n90 163.367
R1198 B.n566 B.n565 163.367
R1199 B.n567 B.n566 163.367
R1200 B.n567 B.n88 163.367
R1201 B.n571 B.n88 163.367
R1202 B.n572 B.n571 163.367
R1203 B.n573 B.n572 163.367
R1204 B.n573 B.n86 163.367
R1205 B.n577 B.n86 163.367
R1206 B.n578 B.n577 163.367
R1207 B.n579 B.n578 163.367
R1208 B.n579 B.n84 163.367
R1209 B.n583 B.n84 163.367
R1210 B.n584 B.n583 163.367
R1211 B.n585 B.n584 163.367
R1212 B.n585 B.n82 163.367
R1213 B.n589 B.n82 163.367
R1214 B.n590 B.n589 163.367
R1215 B.n591 B.n590 163.367
R1216 B.n591 B.n80 163.367
R1217 B.n595 B.n80 163.367
R1218 B.n596 B.n595 163.367
R1219 B.n597 B.n596 163.367
R1220 B.n597 B.n78 163.367
R1221 B.n601 B.n78 163.367
R1222 B.n602 B.n601 163.367
R1223 B.n603 B.n602 163.367
R1224 B.n603 B.n76 163.367
R1225 B.n607 B.n76 163.367
R1226 B.n608 B.n607 163.367
R1227 B.n609 B.n608 163.367
R1228 B.n609 B.n74 163.367
R1229 B.n613 B.n74 163.367
R1230 B.n614 B.n613 163.367
R1231 B.n615 B.n614 163.367
R1232 B.n615 B.n72 163.367
R1233 B.n619 B.n72 163.367
R1234 B.n620 B.n619 163.367
R1235 B.n621 B.n620 163.367
R1236 B.n621 B.n70 163.367
R1237 B.n625 B.n70 163.367
R1238 B.n626 B.n625 163.367
R1239 B.n627 B.n626 163.367
R1240 B.n627 B.n68 163.367
R1241 B.n631 B.n68 163.367
R1242 B.n632 B.n631 163.367
R1243 B.n633 B.n632 163.367
R1244 B.n633 B.n66 163.367
R1245 B.n637 B.n66 163.367
R1246 B.n638 B.n637 163.367
R1247 B.n687 B.n686 163.367
R1248 B.n686 B.n45 163.367
R1249 B.n682 B.n45 163.367
R1250 B.n682 B.n681 163.367
R1251 B.n681 B.n680 163.367
R1252 B.n680 B.n47 163.367
R1253 B.n676 B.n47 163.367
R1254 B.n676 B.n675 163.367
R1255 B.n675 B.n674 163.367
R1256 B.n674 B.n49 163.367
R1257 B.n669 B.n49 163.367
R1258 B.n669 B.n668 163.367
R1259 B.n668 B.n667 163.367
R1260 B.n667 B.n53 163.367
R1261 B.n663 B.n53 163.367
R1262 B.n663 B.n662 163.367
R1263 B.n662 B.n661 163.367
R1264 B.n661 B.n55 163.367
R1265 B.n657 B.n55 163.367
R1266 B.n657 B.n656 163.367
R1267 B.n656 B.n655 163.367
R1268 B.n655 B.n57 163.367
R1269 B.n651 B.n57 163.367
R1270 B.n651 B.n650 163.367
R1271 B.n650 B.n649 163.367
R1272 B.n649 B.n62 163.367
R1273 B.n645 B.n62 163.367
R1274 B.n645 B.n644 163.367
R1275 B.n644 B.n643 163.367
R1276 B.n643 B.n64 163.367
R1277 B.n639 B.n64 163.367
R1278 B.n156 B.n155 83.5884
R1279 B.n164 B.n163 83.5884
R1280 B.n51 B.n50 83.5884
R1281 B.n59 B.n58 83.5884
R1282 B.n157 B.n156 59.5399
R1283 B.n353 B.n164 59.5399
R1284 B.n671 B.n51 59.5399
R1285 B.n60 B.n59 59.5399
R1286 B.n640 B.n65 35.1225
R1287 B.n689 B.n44 35.1224
R1288 B.n384 B.n149 35.1224
R1289 B.n336 B.n335 35.1224
R1290 B B.n815 18.0485
R1291 B.n685 B.n44 10.6151
R1292 B.n685 B.n684 10.6151
R1293 B.n684 B.n683 10.6151
R1294 B.n683 B.n46 10.6151
R1295 B.n679 B.n46 10.6151
R1296 B.n679 B.n678 10.6151
R1297 B.n678 B.n677 10.6151
R1298 B.n677 B.n48 10.6151
R1299 B.n673 B.n48 10.6151
R1300 B.n673 B.n672 10.6151
R1301 B.n670 B.n52 10.6151
R1302 B.n666 B.n52 10.6151
R1303 B.n666 B.n665 10.6151
R1304 B.n665 B.n664 10.6151
R1305 B.n664 B.n54 10.6151
R1306 B.n660 B.n54 10.6151
R1307 B.n660 B.n659 10.6151
R1308 B.n659 B.n658 10.6151
R1309 B.n658 B.n56 10.6151
R1310 B.n654 B.n653 10.6151
R1311 B.n653 B.n652 10.6151
R1312 B.n652 B.n61 10.6151
R1313 B.n648 B.n61 10.6151
R1314 B.n648 B.n647 10.6151
R1315 B.n647 B.n646 10.6151
R1316 B.n646 B.n63 10.6151
R1317 B.n642 B.n63 10.6151
R1318 B.n642 B.n641 10.6151
R1319 B.n641 B.n640 10.6151
R1320 B.n388 B.n149 10.6151
R1321 B.n389 B.n388 10.6151
R1322 B.n390 B.n389 10.6151
R1323 B.n390 B.n147 10.6151
R1324 B.n394 B.n147 10.6151
R1325 B.n395 B.n394 10.6151
R1326 B.n396 B.n395 10.6151
R1327 B.n396 B.n145 10.6151
R1328 B.n400 B.n145 10.6151
R1329 B.n401 B.n400 10.6151
R1330 B.n402 B.n401 10.6151
R1331 B.n402 B.n143 10.6151
R1332 B.n406 B.n143 10.6151
R1333 B.n407 B.n406 10.6151
R1334 B.n408 B.n407 10.6151
R1335 B.n408 B.n141 10.6151
R1336 B.n412 B.n141 10.6151
R1337 B.n413 B.n412 10.6151
R1338 B.n414 B.n413 10.6151
R1339 B.n414 B.n139 10.6151
R1340 B.n418 B.n139 10.6151
R1341 B.n419 B.n418 10.6151
R1342 B.n420 B.n419 10.6151
R1343 B.n420 B.n137 10.6151
R1344 B.n424 B.n137 10.6151
R1345 B.n425 B.n424 10.6151
R1346 B.n426 B.n425 10.6151
R1347 B.n426 B.n135 10.6151
R1348 B.n430 B.n135 10.6151
R1349 B.n431 B.n430 10.6151
R1350 B.n432 B.n431 10.6151
R1351 B.n432 B.n133 10.6151
R1352 B.n436 B.n133 10.6151
R1353 B.n437 B.n436 10.6151
R1354 B.n438 B.n437 10.6151
R1355 B.n438 B.n131 10.6151
R1356 B.n442 B.n131 10.6151
R1357 B.n443 B.n442 10.6151
R1358 B.n444 B.n443 10.6151
R1359 B.n444 B.n129 10.6151
R1360 B.n448 B.n129 10.6151
R1361 B.n449 B.n448 10.6151
R1362 B.n450 B.n449 10.6151
R1363 B.n450 B.n127 10.6151
R1364 B.n454 B.n127 10.6151
R1365 B.n455 B.n454 10.6151
R1366 B.n456 B.n455 10.6151
R1367 B.n456 B.n125 10.6151
R1368 B.n460 B.n125 10.6151
R1369 B.n461 B.n460 10.6151
R1370 B.n462 B.n461 10.6151
R1371 B.n462 B.n123 10.6151
R1372 B.n466 B.n123 10.6151
R1373 B.n467 B.n466 10.6151
R1374 B.n468 B.n467 10.6151
R1375 B.n468 B.n121 10.6151
R1376 B.n472 B.n121 10.6151
R1377 B.n473 B.n472 10.6151
R1378 B.n474 B.n473 10.6151
R1379 B.n474 B.n119 10.6151
R1380 B.n478 B.n119 10.6151
R1381 B.n479 B.n478 10.6151
R1382 B.n480 B.n479 10.6151
R1383 B.n480 B.n117 10.6151
R1384 B.n484 B.n117 10.6151
R1385 B.n485 B.n484 10.6151
R1386 B.n486 B.n485 10.6151
R1387 B.n486 B.n115 10.6151
R1388 B.n490 B.n115 10.6151
R1389 B.n491 B.n490 10.6151
R1390 B.n492 B.n491 10.6151
R1391 B.n492 B.n113 10.6151
R1392 B.n496 B.n113 10.6151
R1393 B.n497 B.n496 10.6151
R1394 B.n498 B.n497 10.6151
R1395 B.n498 B.n111 10.6151
R1396 B.n502 B.n111 10.6151
R1397 B.n503 B.n502 10.6151
R1398 B.n504 B.n503 10.6151
R1399 B.n504 B.n109 10.6151
R1400 B.n508 B.n109 10.6151
R1401 B.n509 B.n508 10.6151
R1402 B.n510 B.n509 10.6151
R1403 B.n510 B.n107 10.6151
R1404 B.n514 B.n107 10.6151
R1405 B.n515 B.n514 10.6151
R1406 B.n516 B.n515 10.6151
R1407 B.n516 B.n105 10.6151
R1408 B.n520 B.n105 10.6151
R1409 B.n521 B.n520 10.6151
R1410 B.n522 B.n521 10.6151
R1411 B.n522 B.n103 10.6151
R1412 B.n526 B.n103 10.6151
R1413 B.n527 B.n526 10.6151
R1414 B.n528 B.n527 10.6151
R1415 B.n528 B.n101 10.6151
R1416 B.n532 B.n101 10.6151
R1417 B.n533 B.n532 10.6151
R1418 B.n534 B.n533 10.6151
R1419 B.n534 B.n99 10.6151
R1420 B.n538 B.n99 10.6151
R1421 B.n539 B.n538 10.6151
R1422 B.n540 B.n539 10.6151
R1423 B.n540 B.n97 10.6151
R1424 B.n544 B.n97 10.6151
R1425 B.n545 B.n544 10.6151
R1426 B.n546 B.n545 10.6151
R1427 B.n546 B.n95 10.6151
R1428 B.n550 B.n95 10.6151
R1429 B.n551 B.n550 10.6151
R1430 B.n552 B.n551 10.6151
R1431 B.n552 B.n93 10.6151
R1432 B.n556 B.n93 10.6151
R1433 B.n557 B.n556 10.6151
R1434 B.n558 B.n557 10.6151
R1435 B.n558 B.n91 10.6151
R1436 B.n562 B.n91 10.6151
R1437 B.n563 B.n562 10.6151
R1438 B.n564 B.n563 10.6151
R1439 B.n564 B.n89 10.6151
R1440 B.n568 B.n89 10.6151
R1441 B.n569 B.n568 10.6151
R1442 B.n570 B.n569 10.6151
R1443 B.n570 B.n87 10.6151
R1444 B.n574 B.n87 10.6151
R1445 B.n575 B.n574 10.6151
R1446 B.n576 B.n575 10.6151
R1447 B.n576 B.n85 10.6151
R1448 B.n580 B.n85 10.6151
R1449 B.n581 B.n580 10.6151
R1450 B.n582 B.n581 10.6151
R1451 B.n582 B.n83 10.6151
R1452 B.n586 B.n83 10.6151
R1453 B.n587 B.n586 10.6151
R1454 B.n588 B.n587 10.6151
R1455 B.n588 B.n81 10.6151
R1456 B.n592 B.n81 10.6151
R1457 B.n593 B.n592 10.6151
R1458 B.n594 B.n593 10.6151
R1459 B.n594 B.n79 10.6151
R1460 B.n598 B.n79 10.6151
R1461 B.n599 B.n598 10.6151
R1462 B.n600 B.n599 10.6151
R1463 B.n600 B.n77 10.6151
R1464 B.n604 B.n77 10.6151
R1465 B.n605 B.n604 10.6151
R1466 B.n606 B.n605 10.6151
R1467 B.n606 B.n75 10.6151
R1468 B.n610 B.n75 10.6151
R1469 B.n611 B.n610 10.6151
R1470 B.n612 B.n611 10.6151
R1471 B.n612 B.n73 10.6151
R1472 B.n616 B.n73 10.6151
R1473 B.n617 B.n616 10.6151
R1474 B.n618 B.n617 10.6151
R1475 B.n618 B.n71 10.6151
R1476 B.n622 B.n71 10.6151
R1477 B.n623 B.n622 10.6151
R1478 B.n624 B.n623 10.6151
R1479 B.n624 B.n69 10.6151
R1480 B.n628 B.n69 10.6151
R1481 B.n629 B.n628 10.6151
R1482 B.n630 B.n629 10.6151
R1483 B.n630 B.n67 10.6151
R1484 B.n634 B.n67 10.6151
R1485 B.n635 B.n634 10.6151
R1486 B.n636 B.n635 10.6151
R1487 B.n636 B.n65 10.6151
R1488 B.n336 B.n169 10.6151
R1489 B.n340 B.n169 10.6151
R1490 B.n341 B.n340 10.6151
R1491 B.n342 B.n341 10.6151
R1492 B.n342 B.n167 10.6151
R1493 B.n346 B.n167 10.6151
R1494 B.n347 B.n346 10.6151
R1495 B.n348 B.n347 10.6151
R1496 B.n348 B.n165 10.6151
R1497 B.n352 B.n165 10.6151
R1498 B.n355 B.n354 10.6151
R1499 B.n355 B.n161 10.6151
R1500 B.n359 B.n161 10.6151
R1501 B.n360 B.n359 10.6151
R1502 B.n361 B.n360 10.6151
R1503 B.n361 B.n159 10.6151
R1504 B.n365 B.n159 10.6151
R1505 B.n366 B.n365 10.6151
R1506 B.n367 B.n366 10.6151
R1507 B.n371 B.n370 10.6151
R1508 B.n372 B.n371 10.6151
R1509 B.n372 B.n153 10.6151
R1510 B.n376 B.n153 10.6151
R1511 B.n377 B.n376 10.6151
R1512 B.n378 B.n377 10.6151
R1513 B.n378 B.n151 10.6151
R1514 B.n382 B.n151 10.6151
R1515 B.n383 B.n382 10.6151
R1516 B.n384 B.n383 10.6151
R1517 B.n335 B.n334 10.6151
R1518 B.n334 B.n171 10.6151
R1519 B.n330 B.n171 10.6151
R1520 B.n330 B.n329 10.6151
R1521 B.n329 B.n328 10.6151
R1522 B.n328 B.n173 10.6151
R1523 B.n324 B.n173 10.6151
R1524 B.n324 B.n323 10.6151
R1525 B.n323 B.n322 10.6151
R1526 B.n322 B.n175 10.6151
R1527 B.n318 B.n175 10.6151
R1528 B.n318 B.n317 10.6151
R1529 B.n317 B.n316 10.6151
R1530 B.n316 B.n177 10.6151
R1531 B.n312 B.n177 10.6151
R1532 B.n312 B.n311 10.6151
R1533 B.n311 B.n310 10.6151
R1534 B.n310 B.n179 10.6151
R1535 B.n306 B.n179 10.6151
R1536 B.n306 B.n305 10.6151
R1537 B.n305 B.n304 10.6151
R1538 B.n304 B.n181 10.6151
R1539 B.n300 B.n181 10.6151
R1540 B.n300 B.n299 10.6151
R1541 B.n299 B.n298 10.6151
R1542 B.n298 B.n183 10.6151
R1543 B.n294 B.n183 10.6151
R1544 B.n294 B.n293 10.6151
R1545 B.n293 B.n292 10.6151
R1546 B.n292 B.n185 10.6151
R1547 B.n288 B.n185 10.6151
R1548 B.n288 B.n287 10.6151
R1549 B.n287 B.n286 10.6151
R1550 B.n286 B.n187 10.6151
R1551 B.n282 B.n187 10.6151
R1552 B.n282 B.n281 10.6151
R1553 B.n281 B.n280 10.6151
R1554 B.n280 B.n189 10.6151
R1555 B.n276 B.n189 10.6151
R1556 B.n276 B.n275 10.6151
R1557 B.n275 B.n274 10.6151
R1558 B.n274 B.n191 10.6151
R1559 B.n270 B.n191 10.6151
R1560 B.n270 B.n269 10.6151
R1561 B.n269 B.n268 10.6151
R1562 B.n268 B.n193 10.6151
R1563 B.n264 B.n193 10.6151
R1564 B.n264 B.n263 10.6151
R1565 B.n263 B.n262 10.6151
R1566 B.n262 B.n195 10.6151
R1567 B.n258 B.n195 10.6151
R1568 B.n258 B.n257 10.6151
R1569 B.n257 B.n256 10.6151
R1570 B.n256 B.n197 10.6151
R1571 B.n252 B.n197 10.6151
R1572 B.n252 B.n251 10.6151
R1573 B.n251 B.n250 10.6151
R1574 B.n250 B.n199 10.6151
R1575 B.n246 B.n199 10.6151
R1576 B.n246 B.n245 10.6151
R1577 B.n245 B.n244 10.6151
R1578 B.n244 B.n201 10.6151
R1579 B.n240 B.n201 10.6151
R1580 B.n240 B.n239 10.6151
R1581 B.n239 B.n238 10.6151
R1582 B.n238 B.n203 10.6151
R1583 B.n234 B.n203 10.6151
R1584 B.n234 B.n233 10.6151
R1585 B.n233 B.n232 10.6151
R1586 B.n232 B.n205 10.6151
R1587 B.n228 B.n205 10.6151
R1588 B.n228 B.n227 10.6151
R1589 B.n227 B.n226 10.6151
R1590 B.n226 B.n207 10.6151
R1591 B.n222 B.n207 10.6151
R1592 B.n222 B.n221 10.6151
R1593 B.n221 B.n220 10.6151
R1594 B.n220 B.n209 10.6151
R1595 B.n216 B.n209 10.6151
R1596 B.n216 B.n215 10.6151
R1597 B.n215 B.n214 10.6151
R1598 B.n214 B.n211 10.6151
R1599 B.n211 B.n0 10.6151
R1600 B.n811 B.n1 10.6151
R1601 B.n811 B.n810 10.6151
R1602 B.n810 B.n809 10.6151
R1603 B.n809 B.n4 10.6151
R1604 B.n805 B.n4 10.6151
R1605 B.n805 B.n804 10.6151
R1606 B.n804 B.n803 10.6151
R1607 B.n803 B.n6 10.6151
R1608 B.n799 B.n6 10.6151
R1609 B.n799 B.n798 10.6151
R1610 B.n798 B.n797 10.6151
R1611 B.n797 B.n8 10.6151
R1612 B.n793 B.n8 10.6151
R1613 B.n793 B.n792 10.6151
R1614 B.n792 B.n791 10.6151
R1615 B.n791 B.n10 10.6151
R1616 B.n787 B.n10 10.6151
R1617 B.n787 B.n786 10.6151
R1618 B.n786 B.n785 10.6151
R1619 B.n785 B.n12 10.6151
R1620 B.n781 B.n12 10.6151
R1621 B.n781 B.n780 10.6151
R1622 B.n780 B.n779 10.6151
R1623 B.n779 B.n14 10.6151
R1624 B.n775 B.n14 10.6151
R1625 B.n775 B.n774 10.6151
R1626 B.n774 B.n773 10.6151
R1627 B.n773 B.n16 10.6151
R1628 B.n769 B.n16 10.6151
R1629 B.n769 B.n768 10.6151
R1630 B.n768 B.n767 10.6151
R1631 B.n767 B.n18 10.6151
R1632 B.n763 B.n18 10.6151
R1633 B.n763 B.n762 10.6151
R1634 B.n762 B.n761 10.6151
R1635 B.n761 B.n20 10.6151
R1636 B.n757 B.n20 10.6151
R1637 B.n757 B.n756 10.6151
R1638 B.n756 B.n755 10.6151
R1639 B.n755 B.n22 10.6151
R1640 B.n751 B.n22 10.6151
R1641 B.n751 B.n750 10.6151
R1642 B.n750 B.n749 10.6151
R1643 B.n749 B.n24 10.6151
R1644 B.n745 B.n24 10.6151
R1645 B.n745 B.n744 10.6151
R1646 B.n744 B.n743 10.6151
R1647 B.n743 B.n26 10.6151
R1648 B.n739 B.n26 10.6151
R1649 B.n739 B.n738 10.6151
R1650 B.n738 B.n737 10.6151
R1651 B.n737 B.n28 10.6151
R1652 B.n733 B.n28 10.6151
R1653 B.n733 B.n732 10.6151
R1654 B.n732 B.n731 10.6151
R1655 B.n731 B.n30 10.6151
R1656 B.n727 B.n30 10.6151
R1657 B.n727 B.n726 10.6151
R1658 B.n726 B.n725 10.6151
R1659 B.n725 B.n32 10.6151
R1660 B.n721 B.n32 10.6151
R1661 B.n721 B.n720 10.6151
R1662 B.n720 B.n719 10.6151
R1663 B.n719 B.n34 10.6151
R1664 B.n715 B.n34 10.6151
R1665 B.n715 B.n714 10.6151
R1666 B.n714 B.n713 10.6151
R1667 B.n713 B.n36 10.6151
R1668 B.n709 B.n36 10.6151
R1669 B.n709 B.n708 10.6151
R1670 B.n708 B.n707 10.6151
R1671 B.n707 B.n38 10.6151
R1672 B.n703 B.n38 10.6151
R1673 B.n703 B.n702 10.6151
R1674 B.n702 B.n701 10.6151
R1675 B.n701 B.n40 10.6151
R1676 B.n697 B.n40 10.6151
R1677 B.n697 B.n696 10.6151
R1678 B.n696 B.n695 10.6151
R1679 B.n695 B.n42 10.6151
R1680 B.n691 B.n42 10.6151
R1681 B.n691 B.n690 10.6151
R1682 B.n690 B.n689 10.6151
R1683 B.n672 B.n671 9.36635
R1684 B.n654 B.n60 9.36635
R1685 B.n353 B.n352 9.36635
R1686 B.n370 B.n157 9.36635
R1687 B.n815 B.n0 2.81026
R1688 B.n815 B.n1 2.81026
R1689 B.n671 B.n670 1.24928
R1690 B.n60 B.n56 1.24928
R1691 B.n354 B.n353 1.24928
R1692 B.n367 B.n157 1.24928
C0 VP VDD1 2.6962f
C1 VP VDD2 0.767987f
C2 VN w_n6142_n1306# 13.4461f
C3 VTAIL w_n6142_n1306# 1.97974f
C4 B w_n6142_n1306# 10.087999f
C5 VDD1 w_n6142_n1306# 2.60276f
C6 VDD2 w_n6142_n1306# 2.81722f
C7 VTAIL VN 4.33419f
C8 B VN 1.52541f
C9 VP w_n6142_n1306# 14.244401f
C10 VDD1 VN 0.163488f
C11 B VTAIL 1.59809f
C12 VDD2 VN 2.09708f
C13 VDD1 VTAIL 7.22941f
C14 B VDD1 2.17925f
C15 VP VN 8.53625f
C16 VDD2 VTAIL 7.29219f
C17 B VDD2 2.35148f
C18 VP VTAIL 4.3484f
C19 B VP 2.88397f
C20 VDD2 VDD1 3.0732f
C21 VDD2 VSUBS 2.715641f
C22 VDD1 VSUBS 2.400377f
C23 VTAIL VSUBS 0.724842f
C24 VN VSUBS 10.60009f
C25 VP VSUBS 5.257891f
C26 B VSUBS 5.799528f
C27 w_n6142_n1306# VSUBS 0.10267p
C28 B.n0 VSUBS 0.009622f
C29 B.n1 VSUBS 0.009622f
C30 B.n2 VSUBS 0.015216f
C31 B.n3 VSUBS 0.015216f
C32 B.n4 VSUBS 0.015216f
C33 B.n5 VSUBS 0.015216f
C34 B.n6 VSUBS 0.015216f
C35 B.n7 VSUBS 0.015216f
C36 B.n8 VSUBS 0.015216f
C37 B.n9 VSUBS 0.015216f
C38 B.n10 VSUBS 0.015216f
C39 B.n11 VSUBS 0.015216f
C40 B.n12 VSUBS 0.015216f
C41 B.n13 VSUBS 0.015216f
C42 B.n14 VSUBS 0.015216f
C43 B.n15 VSUBS 0.015216f
C44 B.n16 VSUBS 0.015216f
C45 B.n17 VSUBS 0.015216f
C46 B.n18 VSUBS 0.015216f
C47 B.n19 VSUBS 0.015216f
C48 B.n20 VSUBS 0.015216f
C49 B.n21 VSUBS 0.015216f
C50 B.n22 VSUBS 0.015216f
C51 B.n23 VSUBS 0.015216f
C52 B.n24 VSUBS 0.015216f
C53 B.n25 VSUBS 0.015216f
C54 B.n26 VSUBS 0.015216f
C55 B.n27 VSUBS 0.015216f
C56 B.n28 VSUBS 0.015216f
C57 B.n29 VSUBS 0.015216f
C58 B.n30 VSUBS 0.015216f
C59 B.n31 VSUBS 0.015216f
C60 B.n32 VSUBS 0.015216f
C61 B.n33 VSUBS 0.015216f
C62 B.n34 VSUBS 0.015216f
C63 B.n35 VSUBS 0.015216f
C64 B.n36 VSUBS 0.015216f
C65 B.n37 VSUBS 0.015216f
C66 B.n38 VSUBS 0.015216f
C67 B.n39 VSUBS 0.015216f
C68 B.n40 VSUBS 0.015216f
C69 B.n41 VSUBS 0.015216f
C70 B.n42 VSUBS 0.015216f
C71 B.n43 VSUBS 0.015216f
C72 B.n44 VSUBS 0.038286f
C73 B.n45 VSUBS 0.015216f
C74 B.n46 VSUBS 0.015216f
C75 B.n47 VSUBS 0.015216f
C76 B.n48 VSUBS 0.015216f
C77 B.n49 VSUBS 0.015216f
C78 B.t5 VSUBS 0.075837f
C79 B.t4 VSUBS 0.103528f
C80 B.t3 VSUBS 0.733886f
C81 B.n50 VSUBS 0.172852f
C82 B.n51 VSUBS 0.132441f
C83 B.n52 VSUBS 0.015216f
C84 B.n53 VSUBS 0.015216f
C85 B.n54 VSUBS 0.015216f
C86 B.n55 VSUBS 0.015216f
C87 B.n56 VSUBS 0.008503f
C88 B.n57 VSUBS 0.015216f
C89 B.t2 VSUBS 0.075837f
C90 B.t1 VSUBS 0.103528f
C91 B.t0 VSUBS 0.733886f
C92 B.n58 VSUBS 0.172852f
C93 B.n59 VSUBS 0.132441f
C94 B.n60 VSUBS 0.035253f
C95 B.n61 VSUBS 0.015216f
C96 B.n62 VSUBS 0.015216f
C97 B.n63 VSUBS 0.015216f
C98 B.n64 VSUBS 0.015216f
C99 B.n65 VSUBS 0.038123f
C100 B.n66 VSUBS 0.015216f
C101 B.n67 VSUBS 0.015216f
C102 B.n68 VSUBS 0.015216f
C103 B.n69 VSUBS 0.015216f
C104 B.n70 VSUBS 0.015216f
C105 B.n71 VSUBS 0.015216f
C106 B.n72 VSUBS 0.015216f
C107 B.n73 VSUBS 0.015216f
C108 B.n74 VSUBS 0.015216f
C109 B.n75 VSUBS 0.015216f
C110 B.n76 VSUBS 0.015216f
C111 B.n77 VSUBS 0.015216f
C112 B.n78 VSUBS 0.015216f
C113 B.n79 VSUBS 0.015216f
C114 B.n80 VSUBS 0.015216f
C115 B.n81 VSUBS 0.015216f
C116 B.n82 VSUBS 0.015216f
C117 B.n83 VSUBS 0.015216f
C118 B.n84 VSUBS 0.015216f
C119 B.n85 VSUBS 0.015216f
C120 B.n86 VSUBS 0.015216f
C121 B.n87 VSUBS 0.015216f
C122 B.n88 VSUBS 0.015216f
C123 B.n89 VSUBS 0.015216f
C124 B.n90 VSUBS 0.015216f
C125 B.n91 VSUBS 0.015216f
C126 B.n92 VSUBS 0.015216f
C127 B.n93 VSUBS 0.015216f
C128 B.n94 VSUBS 0.015216f
C129 B.n95 VSUBS 0.015216f
C130 B.n96 VSUBS 0.015216f
C131 B.n97 VSUBS 0.015216f
C132 B.n98 VSUBS 0.015216f
C133 B.n99 VSUBS 0.015216f
C134 B.n100 VSUBS 0.015216f
C135 B.n101 VSUBS 0.015216f
C136 B.n102 VSUBS 0.015216f
C137 B.n103 VSUBS 0.015216f
C138 B.n104 VSUBS 0.015216f
C139 B.n105 VSUBS 0.015216f
C140 B.n106 VSUBS 0.015216f
C141 B.n107 VSUBS 0.015216f
C142 B.n108 VSUBS 0.015216f
C143 B.n109 VSUBS 0.015216f
C144 B.n110 VSUBS 0.015216f
C145 B.n111 VSUBS 0.015216f
C146 B.n112 VSUBS 0.015216f
C147 B.n113 VSUBS 0.015216f
C148 B.n114 VSUBS 0.015216f
C149 B.n115 VSUBS 0.015216f
C150 B.n116 VSUBS 0.015216f
C151 B.n117 VSUBS 0.015216f
C152 B.n118 VSUBS 0.015216f
C153 B.n119 VSUBS 0.015216f
C154 B.n120 VSUBS 0.015216f
C155 B.n121 VSUBS 0.015216f
C156 B.n122 VSUBS 0.015216f
C157 B.n123 VSUBS 0.015216f
C158 B.n124 VSUBS 0.015216f
C159 B.n125 VSUBS 0.015216f
C160 B.n126 VSUBS 0.015216f
C161 B.n127 VSUBS 0.015216f
C162 B.n128 VSUBS 0.015216f
C163 B.n129 VSUBS 0.015216f
C164 B.n130 VSUBS 0.015216f
C165 B.n131 VSUBS 0.015216f
C166 B.n132 VSUBS 0.015216f
C167 B.n133 VSUBS 0.015216f
C168 B.n134 VSUBS 0.015216f
C169 B.n135 VSUBS 0.015216f
C170 B.n136 VSUBS 0.015216f
C171 B.n137 VSUBS 0.015216f
C172 B.n138 VSUBS 0.015216f
C173 B.n139 VSUBS 0.015216f
C174 B.n140 VSUBS 0.015216f
C175 B.n141 VSUBS 0.015216f
C176 B.n142 VSUBS 0.015216f
C177 B.n143 VSUBS 0.015216f
C178 B.n144 VSUBS 0.015216f
C179 B.n145 VSUBS 0.015216f
C180 B.n146 VSUBS 0.015216f
C181 B.n147 VSUBS 0.015216f
C182 B.n148 VSUBS 0.015216f
C183 B.n149 VSUBS 0.036451f
C184 B.n150 VSUBS 0.015216f
C185 B.n151 VSUBS 0.015216f
C186 B.n152 VSUBS 0.015216f
C187 B.n153 VSUBS 0.015216f
C188 B.n154 VSUBS 0.015216f
C189 B.t7 VSUBS 0.075837f
C190 B.t8 VSUBS 0.103528f
C191 B.t6 VSUBS 0.733886f
C192 B.n155 VSUBS 0.172852f
C193 B.n156 VSUBS 0.132441f
C194 B.n157 VSUBS 0.035253f
C195 B.n158 VSUBS 0.015216f
C196 B.n159 VSUBS 0.015216f
C197 B.n160 VSUBS 0.015216f
C198 B.n161 VSUBS 0.015216f
C199 B.n162 VSUBS 0.015216f
C200 B.t10 VSUBS 0.075837f
C201 B.t11 VSUBS 0.103528f
C202 B.t9 VSUBS 0.733886f
C203 B.n163 VSUBS 0.172852f
C204 B.n164 VSUBS 0.132441f
C205 B.n165 VSUBS 0.015216f
C206 B.n166 VSUBS 0.015216f
C207 B.n167 VSUBS 0.015216f
C208 B.n168 VSUBS 0.015216f
C209 B.n169 VSUBS 0.015216f
C210 B.n170 VSUBS 0.036451f
C211 B.n171 VSUBS 0.015216f
C212 B.n172 VSUBS 0.015216f
C213 B.n173 VSUBS 0.015216f
C214 B.n174 VSUBS 0.015216f
C215 B.n175 VSUBS 0.015216f
C216 B.n176 VSUBS 0.015216f
C217 B.n177 VSUBS 0.015216f
C218 B.n178 VSUBS 0.015216f
C219 B.n179 VSUBS 0.015216f
C220 B.n180 VSUBS 0.015216f
C221 B.n181 VSUBS 0.015216f
C222 B.n182 VSUBS 0.015216f
C223 B.n183 VSUBS 0.015216f
C224 B.n184 VSUBS 0.015216f
C225 B.n185 VSUBS 0.015216f
C226 B.n186 VSUBS 0.015216f
C227 B.n187 VSUBS 0.015216f
C228 B.n188 VSUBS 0.015216f
C229 B.n189 VSUBS 0.015216f
C230 B.n190 VSUBS 0.015216f
C231 B.n191 VSUBS 0.015216f
C232 B.n192 VSUBS 0.015216f
C233 B.n193 VSUBS 0.015216f
C234 B.n194 VSUBS 0.015216f
C235 B.n195 VSUBS 0.015216f
C236 B.n196 VSUBS 0.015216f
C237 B.n197 VSUBS 0.015216f
C238 B.n198 VSUBS 0.015216f
C239 B.n199 VSUBS 0.015216f
C240 B.n200 VSUBS 0.015216f
C241 B.n201 VSUBS 0.015216f
C242 B.n202 VSUBS 0.015216f
C243 B.n203 VSUBS 0.015216f
C244 B.n204 VSUBS 0.015216f
C245 B.n205 VSUBS 0.015216f
C246 B.n206 VSUBS 0.015216f
C247 B.n207 VSUBS 0.015216f
C248 B.n208 VSUBS 0.015216f
C249 B.n209 VSUBS 0.015216f
C250 B.n210 VSUBS 0.015216f
C251 B.n211 VSUBS 0.015216f
C252 B.n212 VSUBS 0.015216f
C253 B.n213 VSUBS 0.015216f
C254 B.n214 VSUBS 0.015216f
C255 B.n215 VSUBS 0.015216f
C256 B.n216 VSUBS 0.015216f
C257 B.n217 VSUBS 0.015216f
C258 B.n218 VSUBS 0.015216f
C259 B.n219 VSUBS 0.015216f
C260 B.n220 VSUBS 0.015216f
C261 B.n221 VSUBS 0.015216f
C262 B.n222 VSUBS 0.015216f
C263 B.n223 VSUBS 0.015216f
C264 B.n224 VSUBS 0.015216f
C265 B.n225 VSUBS 0.015216f
C266 B.n226 VSUBS 0.015216f
C267 B.n227 VSUBS 0.015216f
C268 B.n228 VSUBS 0.015216f
C269 B.n229 VSUBS 0.015216f
C270 B.n230 VSUBS 0.015216f
C271 B.n231 VSUBS 0.015216f
C272 B.n232 VSUBS 0.015216f
C273 B.n233 VSUBS 0.015216f
C274 B.n234 VSUBS 0.015216f
C275 B.n235 VSUBS 0.015216f
C276 B.n236 VSUBS 0.015216f
C277 B.n237 VSUBS 0.015216f
C278 B.n238 VSUBS 0.015216f
C279 B.n239 VSUBS 0.015216f
C280 B.n240 VSUBS 0.015216f
C281 B.n241 VSUBS 0.015216f
C282 B.n242 VSUBS 0.015216f
C283 B.n243 VSUBS 0.015216f
C284 B.n244 VSUBS 0.015216f
C285 B.n245 VSUBS 0.015216f
C286 B.n246 VSUBS 0.015216f
C287 B.n247 VSUBS 0.015216f
C288 B.n248 VSUBS 0.015216f
C289 B.n249 VSUBS 0.015216f
C290 B.n250 VSUBS 0.015216f
C291 B.n251 VSUBS 0.015216f
C292 B.n252 VSUBS 0.015216f
C293 B.n253 VSUBS 0.015216f
C294 B.n254 VSUBS 0.015216f
C295 B.n255 VSUBS 0.015216f
C296 B.n256 VSUBS 0.015216f
C297 B.n257 VSUBS 0.015216f
C298 B.n258 VSUBS 0.015216f
C299 B.n259 VSUBS 0.015216f
C300 B.n260 VSUBS 0.015216f
C301 B.n261 VSUBS 0.015216f
C302 B.n262 VSUBS 0.015216f
C303 B.n263 VSUBS 0.015216f
C304 B.n264 VSUBS 0.015216f
C305 B.n265 VSUBS 0.015216f
C306 B.n266 VSUBS 0.015216f
C307 B.n267 VSUBS 0.015216f
C308 B.n268 VSUBS 0.015216f
C309 B.n269 VSUBS 0.015216f
C310 B.n270 VSUBS 0.015216f
C311 B.n271 VSUBS 0.015216f
C312 B.n272 VSUBS 0.015216f
C313 B.n273 VSUBS 0.015216f
C314 B.n274 VSUBS 0.015216f
C315 B.n275 VSUBS 0.015216f
C316 B.n276 VSUBS 0.015216f
C317 B.n277 VSUBS 0.015216f
C318 B.n278 VSUBS 0.015216f
C319 B.n279 VSUBS 0.015216f
C320 B.n280 VSUBS 0.015216f
C321 B.n281 VSUBS 0.015216f
C322 B.n282 VSUBS 0.015216f
C323 B.n283 VSUBS 0.015216f
C324 B.n284 VSUBS 0.015216f
C325 B.n285 VSUBS 0.015216f
C326 B.n286 VSUBS 0.015216f
C327 B.n287 VSUBS 0.015216f
C328 B.n288 VSUBS 0.015216f
C329 B.n289 VSUBS 0.015216f
C330 B.n290 VSUBS 0.015216f
C331 B.n291 VSUBS 0.015216f
C332 B.n292 VSUBS 0.015216f
C333 B.n293 VSUBS 0.015216f
C334 B.n294 VSUBS 0.015216f
C335 B.n295 VSUBS 0.015216f
C336 B.n296 VSUBS 0.015216f
C337 B.n297 VSUBS 0.015216f
C338 B.n298 VSUBS 0.015216f
C339 B.n299 VSUBS 0.015216f
C340 B.n300 VSUBS 0.015216f
C341 B.n301 VSUBS 0.015216f
C342 B.n302 VSUBS 0.015216f
C343 B.n303 VSUBS 0.015216f
C344 B.n304 VSUBS 0.015216f
C345 B.n305 VSUBS 0.015216f
C346 B.n306 VSUBS 0.015216f
C347 B.n307 VSUBS 0.015216f
C348 B.n308 VSUBS 0.015216f
C349 B.n309 VSUBS 0.015216f
C350 B.n310 VSUBS 0.015216f
C351 B.n311 VSUBS 0.015216f
C352 B.n312 VSUBS 0.015216f
C353 B.n313 VSUBS 0.015216f
C354 B.n314 VSUBS 0.015216f
C355 B.n315 VSUBS 0.015216f
C356 B.n316 VSUBS 0.015216f
C357 B.n317 VSUBS 0.015216f
C358 B.n318 VSUBS 0.015216f
C359 B.n319 VSUBS 0.015216f
C360 B.n320 VSUBS 0.015216f
C361 B.n321 VSUBS 0.015216f
C362 B.n322 VSUBS 0.015216f
C363 B.n323 VSUBS 0.015216f
C364 B.n324 VSUBS 0.015216f
C365 B.n325 VSUBS 0.015216f
C366 B.n326 VSUBS 0.015216f
C367 B.n327 VSUBS 0.015216f
C368 B.n328 VSUBS 0.015216f
C369 B.n329 VSUBS 0.015216f
C370 B.n330 VSUBS 0.015216f
C371 B.n331 VSUBS 0.015216f
C372 B.n332 VSUBS 0.015216f
C373 B.n333 VSUBS 0.015216f
C374 B.n334 VSUBS 0.015216f
C375 B.n335 VSUBS 0.036451f
C376 B.n336 VSUBS 0.038286f
C377 B.n337 VSUBS 0.038286f
C378 B.n338 VSUBS 0.015216f
C379 B.n339 VSUBS 0.015216f
C380 B.n340 VSUBS 0.015216f
C381 B.n341 VSUBS 0.015216f
C382 B.n342 VSUBS 0.015216f
C383 B.n343 VSUBS 0.015216f
C384 B.n344 VSUBS 0.015216f
C385 B.n345 VSUBS 0.015216f
C386 B.n346 VSUBS 0.015216f
C387 B.n347 VSUBS 0.015216f
C388 B.n348 VSUBS 0.015216f
C389 B.n349 VSUBS 0.015216f
C390 B.n350 VSUBS 0.015216f
C391 B.n351 VSUBS 0.015216f
C392 B.n352 VSUBS 0.014321f
C393 B.n353 VSUBS 0.035253f
C394 B.n354 VSUBS 0.008503f
C395 B.n355 VSUBS 0.015216f
C396 B.n356 VSUBS 0.015216f
C397 B.n357 VSUBS 0.015216f
C398 B.n358 VSUBS 0.015216f
C399 B.n359 VSUBS 0.015216f
C400 B.n360 VSUBS 0.015216f
C401 B.n361 VSUBS 0.015216f
C402 B.n362 VSUBS 0.015216f
C403 B.n363 VSUBS 0.015216f
C404 B.n364 VSUBS 0.015216f
C405 B.n365 VSUBS 0.015216f
C406 B.n366 VSUBS 0.015216f
C407 B.n367 VSUBS 0.008503f
C408 B.n368 VSUBS 0.015216f
C409 B.n369 VSUBS 0.015216f
C410 B.n370 VSUBS 0.014321f
C411 B.n371 VSUBS 0.015216f
C412 B.n372 VSUBS 0.015216f
C413 B.n373 VSUBS 0.015216f
C414 B.n374 VSUBS 0.015216f
C415 B.n375 VSUBS 0.015216f
C416 B.n376 VSUBS 0.015216f
C417 B.n377 VSUBS 0.015216f
C418 B.n378 VSUBS 0.015216f
C419 B.n379 VSUBS 0.015216f
C420 B.n380 VSUBS 0.015216f
C421 B.n381 VSUBS 0.015216f
C422 B.n382 VSUBS 0.015216f
C423 B.n383 VSUBS 0.015216f
C424 B.n384 VSUBS 0.038286f
C425 B.n385 VSUBS 0.038286f
C426 B.n386 VSUBS 0.036451f
C427 B.n387 VSUBS 0.015216f
C428 B.n388 VSUBS 0.015216f
C429 B.n389 VSUBS 0.015216f
C430 B.n390 VSUBS 0.015216f
C431 B.n391 VSUBS 0.015216f
C432 B.n392 VSUBS 0.015216f
C433 B.n393 VSUBS 0.015216f
C434 B.n394 VSUBS 0.015216f
C435 B.n395 VSUBS 0.015216f
C436 B.n396 VSUBS 0.015216f
C437 B.n397 VSUBS 0.015216f
C438 B.n398 VSUBS 0.015216f
C439 B.n399 VSUBS 0.015216f
C440 B.n400 VSUBS 0.015216f
C441 B.n401 VSUBS 0.015216f
C442 B.n402 VSUBS 0.015216f
C443 B.n403 VSUBS 0.015216f
C444 B.n404 VSUBS 0.015216f
C445 B.n405 VSUBS 0.015216f
C446 B.n406 VSUBS 0.015216f
C447 B.n407 VSUBS 0.015216f
C448 B.n408 VSUBS 0.015216f
C449 B.n409 VSUBS 0.015216f
C450 B.n410 VSUBS 0.015216f
C451 B.n411 VSUBS 0.015216f
C452 B.n412 VSUBS 0.015216f
C453 B.n413 VSUBS 0.015216f
C454 B.n414 VSUBS 0.015216f
C455 B.n415 VSUBS 0.015216f
C456 B.n416 VSUBS 0.015216f
C457 B.n417 VSUBS 0.015216f
C458 B.n418 VSUBS 0.015216f
C459 B.n419 VSUBS 0.015216f
C460 B.n420 VSUBS 0.015216f
C461 B.n421 VSUBS 0.015216f
C462 B.n422 VSUBS 0.015216f
C463 B.n423 VSUBS 0.015216f
C464 B.n424 VSUBS 0.015216f
C465 B.n425 VSUBS 0.015216f
C466 B.n426 VSUBS 0.015216f
C467 B.n427 VSUBS 0.015216f
C468 B.n428 VSUBS 0.015216f
C469 B.n429 VSUBS 0.015216f
C470 B.n430 VSUBS 0.015216f
C471 B.n431 VSUBS 0.015216f
C472 B.n432 VSUBS 0.015216f
C473 B.n433 VSUBS 0.015216f
C474 B.n434 VSUBS 0.015216f
C475 B.n435 VSUBS 0.015216f
C476 B.n436 VSUBS 0.015216f
C477 B.n437 VSUBS 0.015216f
C478 B.n438 VSUBS 0.015216f
C479 B.n439 VSUBS 0.015216f
C480 B.n440 VSUBS 0.015216f
C481 B.n441 VSUBS 0.015216f
C482 B.n442 VSUBS 0.015216f
C483 B.n443 VSUBS 0.015216f
C484 B.n444 VSUBS 0.015216f
C485 B.n445 VSUBS 0.015216f
C486 B.n446 VSUBS 0.015216f
C487 B.n447 VSUBS 0.015216f
C488 B.n448 VSUBS 0.015216f
C489 B.n449 VSUBS 0.015216f
C490 B.n450 VSUBS 0.015216f
C491 B.n451 VSUBS 0.015216f
C492 B.n452 VSUBS 0.015216f
C493 B.n453 VSUBS 0.015216f
C494 B.n454 VSUBS 0.015216f
C495 B.n455 VSUBS 0.015216f
C496 B.n456 VSUBS 0.015216f
C497 B.n457 VSUBS 0.015216f
C498 B.n458 VSUBS 0.015216f
C499 B.n459 VSUBS 0.015216f
C500 B.n460 VSUBS 0.015216f
C501 B.n461 VSUBS 0.015216f
C502 B.n462 VSUBS 0.015216f
C503 B.n463 VSUBS 0.015216f
C504 B.n464 VSUBS 0.015216f
C505 B.n465 VSUBS 0.015216f
C506 B.n466 VSUBS 0.015216f
C507 B.n467 VSUBS 0.015216f
C508 B.n468 VSUBS 0.015216f
C509 B.n469 VSUBS 0.015216f
C510 B.n470 VSUBS 0.015216f
C511 B.n471 VSUBS 0.015216f
C512 B.n472 VSUBS 0.015216f
C513 B.n473 VSUBS 0.015216f
C514 B.n474 VSUBS 0.015216f
C515 B.n475 VSUBS 0.015216f
C516 B.n476 VSUBS 0.015216f
C517 B.n477 VSUBS 0.015216f
C518 B.n478 VSUBS 0.015216f
C519 B.n479 VSUBS 0.015216f
C520 B.n480 VSUBS 0.015216f
C521 B.n481 VSUBS 0.015216f
C522 B.n482 VSUBS 0.015216f
C523 B.n483 VSUBS 0.015216f
C524 B.n484 VSUBS 0.015216f
C525 B.n485 VSUBS 0.015216f
C526 B.n486 VSUBS 0.015216f
C527 B.n487 VSUBS 0.015216f
C528 B.n488 VSUBS 0.015216f
C529 B.n489 VSUBS 0.015216f
C530 B.n490 VSUBS 0.015216f
C531 B.n491 VSUBS 0.015216f
C532 B.n492 VSUBS 0.015216f
C533 B.n493 VSUBS 0.015216f
C534 B.n494 VSUBS 0.015216f
C535 B.n495 VSUBS 0.015216f
C536 B.n496 VSUBS 0.015216f
C537 B.n497 VSUBS 0.015216f
C538 B.n498 VSUBS 0.015216f
C539 B.n499 VSUBS 0.015216f
C540 B.n500 VSUBS 0.015216f
C541 B.n501 VSUBS 0.015216f
C542 B.n502 VSUBS 0.015216f
C543 B.n503 VSUBS 0.015216f
C544 B.n504 VSUBS 0.015216f
C545 B.n505 VSUBS 0.015216f
C546 B.n506 VSUBS 0.015216f
C547 B.n507 VSUBS 0.015216f
C548 B.n508 VSUBS 0.015216f
C549 B.n509 VSUBS 0.015216f
C550 B.n510 VSUBS 0.015216f
C551 B.n511 VSUBS 0.015216f
C552 B.n512 VSUBS 0.015216f
C553 B.n513 VSUBS 0.015216f
C554 B.n514 VSUBS 0.015216f
C555 B.n515 VSUBS 0.015216f
C556 B.n516 VSUBS 0.015216f
C557 B.n517 VSUBS 0.015216f
C558 B.n518 VSUBS 0.015216f
C559 B.n519 VSUBS 0.015216f
C560 B.n520 VSUBS 0.015216f
C561 B.n521 VSUBS 0.015216f
C562 B.n522 VSUBS 0.015216f
C563 B.n523 VSUBS 0.015216f
C564 B.n524 VSUBS 0.015216f
C565 B.n525 VSUBS 0.015216f
C566 B.n526 VSUBS 0.015216f
C567 B.n527 VSUBS 0.015216f
C568 B.n528 VSUBS 0.015216f
C569 B.n529 VSUBS 0.015216f
C570 B.n530 VSUBS 0.015216f
C571 B.n531 VSUBS 0.015216f
C572 B.n532 VSUBS 0.015216f
C573 B.n533 VSUBS 0.015216f
C574 B.n534 VSUBS 0.015216f
C575 B.n535 VSUBS 0.015216f
C576 B.n536 VSUBS 0.015216f
C577 B.n537 VSUBS 0.015216f
C578 B.n538 VSUBS 0.015216f
C579 B.n539 VSUBS 0.015216f
C580 B.n540 VSUBS 0.015216f
C581 B.n541 VSUBS 0.015216f
C582 B.n542 VSUBS 0.015216f
C583 B.n543 VSUBS 0.015216f
C584 B.n544 VSUBS 0.015216f
C585 B.n545 VSUBS 0.015216f
C586 B.n546 VSUBS 0.015216f
C587 B.n547 VSUBS 0.015216f
C588 B.n548 VSUBS 0.015216f
C589 B.n549 VSUBS 0.015216f
C590 B.n550 VSUBS 0.015216f
C591 B.n551 VSUBS 0.015216f
C592 B.n552 VSUBS 0.015216f
C593 B.n553 VSUBS 0.015216f
C594 B.n554 VSUBS 0.015216f
C595 B.n555 VSUBS 0.015216f
C596 B.n556 VSUBS 0.015216f
C597 B.n557 VSUBS 0.015216f
C598 B.n558 VSUBS 0.015216f
C599 B.n559 VSUBS 0.015216f
C600 B.n560 VSUBS 0.015216f
C601 B.n561 VSUBS 0.015216f
C602 B.n562 VSUBS 0.015216f
C603 B.n563 VSUBS 0.015216f
C604 B.n564 VSUBS 0.015216f
C605 B.n565 VSUBS 0.015216f
C606 B.n566 VSUBS 0.015216f
C607 B.n567 VSUBS 0.015216f
C608 B.n568 VSUBS 0.015216f
C609 B.n569 VSUBS 0.015216f
C610 B.n570 VSUBS 0.015216f
C611 B.n571 VSUBS 0.015216f
C612 B.n572 VSUBS 0.015216f
C613 B.n573 VSUBS 0.015216f
C614 B.n574 VSUBS 0.015216f
C615 B.n575 VSUBS 0.015216f
C616 B.n576 VSUBS 0.015216f
C617 B.n577 VSUBS 0.015216f
C618 B.n578 VSUBS 0.015216f
C619 B.n579 VSUBS 0.015216f
C620 B.n580 VSUBS 0.015216f
C621 B.n581 VSUBS 0.015216f
C622 B.n582 VSUBS 0.015216f
C623 B.n583 VSUBS 0.015216f
C624 B.n584 VSUBS 0.015216f
C625 B.n585 VSUBS 0.015216f
C626 B.n586 VSUBS 0.015216f
C627 B.n587 VSUBS 0.015216f
C628 B.n588 VSUBS 0.015216f
C629 B.n589 VSUBS 0.015216f
C630 B.n590 VSUBS 0.015216f
C631 B.n591 VSUBS 0.015216f
C632 B.n592 VSUBS 0.015216f
C633 B.n593 VSUBS 0.015216f
C634 B.n594 VSUBS 0.015216f
C635 B.n595 VSUBS 0.015216f
C636 B.n596 VSUBS 0.015216f
C637 B.n597 VSUBS 0.015216f
C638 B.n598 VSUBS 0.015216f
C639 B.n599 VSUBS 0.015216f
C640 B.n600 VSUBS 0.015216f
C641 B.n601 VSUBS 0.015216f
C642 B.n602 VSUBS 0.015216f
C643 B.n603 VSUBS 0.015216f
C644 B.n604 VSUBS 0.015216f
C645 B.n605 VSUBS 0.015216f
C646 B.n606 VSUBS 0.015216f
C647 B.n607 VSUBS 0.015216f
C648 B.n608 VSUBS 0.015216f
C649 B.n609 VSUBS 0.015216f
C650 B.n610 VSUBS 0.015216f
C651 B.n611 VSUBS 0.015216f
C652 B.n612 VSUBS 0.015216f
C653 B.n613 VSUBS 0.015216f
C654 B.n614 VSUBS 0.015216f
C655 B.n615 VSUBS 0.015216f
C656 B.n616 VSUBS 0.015216f
C657 B.n617 VSUBS 0.015216f
C658 B.n618 VSUBS 0.015216f
C659 B.n619 VSUBS 0.015216f
C660 B.n620 VSUBS 0.015216f
C661 B.n621 VSUBS 0.015216f
C662 B.n622 VSUBS 0.015216f
C663 B.n623 VSUBS 0.015216f
C664 B.n624 VSUBS 0.015216f
C665 B.n625 VSUBS 0.015216f
C666 B.n626 VSUBS 0.015216f
C667 B.n627 VSUBS 0.015216f
C668 B.n628 VSUBS 0.015216f
C669 B.n629 VSUBS 0.015216f
C670 B.n630 VSUBS 0.015216f
C671 B.n631 VSUBS 0.015216f
C672 B.n632 VSUBS 0.015216f
C673 B.n633 VSUBS 0.015216f
C674 B.n634 VSUBS 0.015216f
C675 B.n635 VSUBS 0.015216f
C676 B.n636 VSUBS 0.015216f
C677 B.n637 VSUBS 0.015216f
C678 B.n638 VSUBS 0.036451f
C679 B.n639 VSUBS 0.038286f
C680 B.n640 VSUBS 0.036614f
C681 B.n641 VSUBS 0.015216f
C682 B.n642 VSUBS 0.015216f
C683 B.n643 VSUBS 0.015216f
C684 B.n644 VSUBS 0.015216f
C685 B.n645 VSUBS 0.015216f
C686 B.n646 VSUBS 0.015216f
C687 B.n647 VSUBS 0.015216f
C688 B.n648 VSUBS 0.015216f
C689 B.n649 VSUBS 0.015216f
C690 B.n650 VSUBS 0.015216f
C691 B.n651 VSUBS 0.015216f
C692 B.n652 VSUBS 0.015216f
C693 B.n653 VSUBS 0.015216f
C694 B.n654 VSUBS 0.014321f
C695 B.n655 VSUBS 0.015216f
C696 B.n656 VSUBS 0.015216f
C697 B.n657 VSUBS 0.015216f
C698 B.n658 VSUBS 0.015216f
C699 B.n659 VSUBS 0.015216f
C700 B.n660 VSUBS 0.015216f
C701 B.n661 VSUBS 0.015216f
C702 B.n662 VSUBS 0.015216f
C703 B.n663 VSUBS 0.015216f
C704 B.n664 VSUBS 0.015216f
C705 B.n665 VSUBS 0.015216f
C706 B.n666 VSUBS 0.015216f
C707 B.n667 VSUBS 0.015216f
C708 B.n668 VSUBS 0.015216f
C709 B.n669 VSUBS 0.015216f
C710 B.n670 VSUBS 0.008503f
C711 B.n671 VSUBS 0.035253f
C712 B.n672 VSUBS 0.014321f
C713 B.n673 VSUBS 0.015216f
C714 B.n674 VSUBS 0.015216f
C715 B.n675 VSUBS 0.015216f
C716 B.n676 VSUBS 0.015216f
C717 B.n677 VSUBS 0.015216f
C718 B.n678 VSUBS 0.015216f
C719 B.n679 VSUBS 0.015216f
C720 B.n680 VSUBS 0.015216f
C721 B.n681 VSUBS 0.015216f
C722 B.n682 VSUBS 0.015216f
C723 B.n683 VSUBS 0.015216f
C724 B.n684 VSUBS 0.015216f
C725 B.n685 VSUBS 0.015216f
C726 B.n686 VSUBS 0.015216f
C727 B.n687 VSUBS 0.038286f
C728 B.n688 VSUBS 0.036451f
C729 B.n689 VSUBS 0.036451f
C730 B.n690 VSUBS 0.015216f
C731 B.n691 VSUBS 0.015216f
C732 B.n692 VSUBS 0.015216f
C733 B.n693 VSUBS 0.015216f
C734 B.n694 VSUBS 0.015216f
C735 B.n695 VSUBS 0.015216f
C736 B.n696 VSUBS 0.015216f
C737 B.n697 VSUBS 0.015216f
C738 B.n698 VSUBS 0.015216f
C739 B.n699 VSUBS 0.015216f
C740 B.n700 VSUBS 0.015216f
C741 B.n701 VSUBS 0.015216f
C742 B.n702 VSUBS 0.015216f
C743 B.n703 VSUBS 0.015216f
C744 B.n704 VSUBS 0.015216f
C745 B.n705 VSUBS 0.015216f
C746 B.n706 VSUBS 0.015216f
C747 B.n707 VSUBS 0.015216f
C748 B.n708 VSUBS 0.015216f
C749 B.n709 VSUBS 0.015216f
C750 B.n710 VSUBS 0.015216f
C751 B.n711 VSUBS 0.015216f
C752 B.n712 VSUBS 0.015216f
C753 B.n713 VSUBS 0.015216f
C754 B.n714 VSUBS 0.015216f
C755 B.n715 VSUBS 0.015216f
C756 B.n716 VSUBS 0.015216f
C757 B.n717 VSUBS 0.015216f
C758 B.n718 VSUBS 0.015216f
C759 B.n719 VSUBS 0.015216f
C760 B.n720 VSUBS 0.015216f
C761 B.n721 VSUBS 0.015216f
C762 B.n722 VSUBS 0.015216f
C763 B.n723 VSUBS 0.015216f
C764 B.n724 VSUBS 0.015216f
C765 B.n725 VSUBS 0.015216f
C766 B.n726 VSUBS 0.015216f
C767 B.n727 VSUBS 0.015216f
C768 B.n728 VSUBS 0.015216f
C769 B.n729 VSUBS 0.015216f
C770 B.n730 VSUBS 0.015216f
C771 B.n731 VSUBS 0.015216f
C772 B.n732 VSUBS 0.015216f
C773 B.n733 VSUBS 0.015216f
C774 B.n734 VSUBS 0.015216f
C775 B.n735 VSUBS 0.015216f
C776 B.n736 VSUBS 0.015216f
C777 B.n737 VSUBS 0.015216f
C778 B.n738 VSUBS 0.015216f
C779 B.n739 VSUBS 0.015216f
C780 B.n740 VSUBS 0.015216f
C781 B.n741 VSUBS 0.015216f
C782 B.n742 VSUBS 0.015216f
C783 B.n743 VSUBS 0.015216f
C784 B.n744 VSUBS 0.015216f
C785 B.n745 VSUBS 0.015216f
C786 B.n746 VSUBS 0.015216f
C787 B.n747 VSUBS 0.015216f
C788 B.n748 VSUBS 0.015216f
C789 B.n749 VSUBS 0.015216f
C790 B.n750 VSUBS 0.015216f
C791 B.n751 VSUBS 0.015216f
C792 B.n752 VSUBS 0.015216f
C793 B.n753 VSUBS 0.015216f
C794 B.n754 VSUBS 0.015216f
C795 B.n755 VSUBS 0.015216f
C796 B.n756 VSUBS 0.015216f
C797 B.n757 VSUBS 0.015216f
C798 B.n758 VSUBS 0.015216f
C799 B.n759 VSUBS 0.015216f
C800 B.n760 VSUBS 0.015216f
C801 B.n761 VSUBS 0.015216f
C802 B.n762 VSUBS 0.015216f
C803 B.n763 VSUBS 0.015216f
C804 B.n764 VSUBS 0.015216f
C805 B.n765 VSUBS 0.015216f
C806 B.n766 VSUBS 0.015216f
C807 B.n767 VSUBS 0.015216f
C808 B.n768 VSUBS 0.015216f
C809 B.n769 VSUBS 0.015216f
C810 B.n770 VSUBS 0.015216f
C811 B.n771 VSUBS 0.015216f
C812 B.n772 VSUBS 0.015216f
C813 B.n773 VSUBS 0.015216f
C814 B.n774 VSUBS 0.015216f
C815 B.n775 VSUBS 0.015216f
C816 B.n776 VSUBS 0.015216f
C817 B.n777 VSUBS 0.015216f
C818 B.n778 VSUBS 0.015216f
C819 B.n779 VSUBS 0.015216f
C820 B.n780 VSUBS 0.015216f
C821 B.n781 VSUBS 0.015216f
C822 B.n782 VSUBS 0.015216f
C823 B.n783 VSUBS 0.015216f
C824 B.n784 VSUBS 0.015216f
C825 B.n785 VSUBS 0.015216f
C826 B.n786 VSUBS 0.015216f
C827 B.n787 VSUBS 0.015216f
C828 B.n788 VSUBS 0.015216f
C829 B.n789 VSUBS 0.015216f
C830 B.n790 VSUBS 0.015216f
C831 B.n791 VSUBS 0.015216f
C832 B.n792 VSUBS 0.015216f
C833 B.n793 VSUBS 0.015216f
C834 B.n794 VSUBS 0.015216f
C835 B.n795 VSUBS 0.015216f
C836 B.n796 VSUBS 0.015216f
C837 B.n797 VSUBS 0.015216f
C838 B.n798 VSUBS 0.015216f
C839 B.n799 VSUBS 0.015216f
C840 B.n800 VSUBS 0.015216f
C841 B.n801 VSUBS 0.015216f
C842 B.n802 VSUBS 0.015216f
C843 B.n803 VSUBS 0.015216f
C844 B.n804 VSUBS 0.015216f
C845 B.n805 VSUBS 0.015216f
C846 B.n806 VSUBS 0.015216f
C847 B.n807 VSUBS 0.015216f
C848 B.n808 VSUBS 0.015216f
C849 B.n809 VSUBS 0.015216f
C850 B.n810 VSUBS 0.015216f
C851 B.n811 VSUBS 0.015216f
C852 B.n812 VSUBS 0.015216f
C853 B.n813 VSUBS 0.015216f
C854 B.n814 VSUBS 0.015216f
C855 B.n815 VSUBS 0.034454f
C856 VDD2.t0 VSUBS 0.373014f
C857 VDD2.t3 VSUBS 0.058918f
C858 VDD2.t1 VSUBS 0.058918f
C859 VDD2.n0 VSUBS 0.221525f
C860 VDD2.n1 VSUBS 2.11135f
C861 VDD2.t5 VSUBS 0.058918f
C862 VDD2.t2 VSUBS 0.058918f
C863 VDD2.n2 VSUBS 0.236485f
C864 VDD2.n3 VSUBS 5.40916f
C865 VDD2.t7 VSUBS 0.35914f
C866 VDD2.n4 VSUBS 5.04177f
C867 VDD2.t9 VSUBS 0.058918f
C868 VDD2.t4 VSUBS 0.058918f
C869 VDD2.n5 VSUBS 0.221525f
C870 VDD2.n6 VSUBS 1.11984f
C871 VDD2.t8 VSUBS 0.058918f
C872 VDD2.t6 VSUBS 0.058918f
C873 VDD2.n7 VSUBS 0.236461f
C874 VN.n0 VSUBS 0.093954f
C875 VN.t7 VSUBS 0.755826f
C876 VN.n1 VSUBS 0.093092f
C877 VN.n2 VSUBS 0.049949f
C878 VN.n3 VSUBS 0.093092f
C879 VN.n4 VSUBS 0.049949f
C880 VN.t4 VSUBS 0.755826f
C881 VN.n5 VSUBS 0.093092f
C882 VN.n6 VSUBS 0.049949f
C883 VN.n7 VSUBS 0.093092f
C884 VN.n8 VSUBS 0.049949f
C885 VN.t8 VSUBS 0.755826f
C886 VN.n9 VSUBS 0.093092f
C887 VN.n10 VSUBS 0.049949f
C888 VN.n11 VSUBS 0.100288f
C889 VN.n12 VSUBS 0.049949f
C890 VN.t6 VSUBS 0.755826f
C891 VN.n13 VSUBS 0.52589f
C892 VN.t9 VSUBS 1.32554f
C893 VN.n14 VSUBS 0.654773f
C894 VN.n15 VSUBS 0.670847f
C895 VN.n16 VSUBS 0.052647f
C896 VN.n17 VSUBS 0.093092f
C897 VN.n18 VSUBS 0.093092f
C898 VN.n19 VSUBS 0.049949f
C899 VN.n20 VSUBS 0.049949f
C900 VN.n21 VSUBS 0.049949f
C901 VN.n22 VSUBS 0.046488f
C902 VN.n23 VSUBS 0.092158f
C903 VN.n24 VSUBS 0.093092f
C904 VN.n25 VSUBS 0.049949f
C905 VN.n26 VSUBS 0.049949f
C906 VN.n27 VSUBS 0.049949f
C907 VN.n28 VSUBS 0.070112f
C908 VN.n29 VSUBS 0.359804f
C909 VN.n30 VSUBS 0.070112f
C910 VN.n31 VSUBS 0.093092f
C911 VN.n32 VSUBS 0.049949f
C912 VN.n33 VSUBS 0.049949f
C913 VN.n34 VSUBS 0.049949f
C914 VN.n35 VSUBS 0.092158f
C915 VN.n36 VSUBS 0.046488f
C916 VN.n37 VSUBS 0.100288f
C917 VN.n38 VSUBS 0.049949f
C918 VN.n39 VSUBS 0.049949f
C919 VN.n40 VSUBS 0.049949f
C920 VN.n41 VSUBS 0.093092f
C921 VN.n42 VSUBS 0.052647f
C922 VN.n43 VSUBS 0.359804f
C923 VN.n44 VSUBS 0.087577f
C924 VN.n45 VSUBS 0.049949f
C925 VN.n46 VSUBS 0.049949f
C926 VN.n47 VSUBS 0.049949f
C927 VN.n48 VSUBS 0.093092f
C928 VN.n49 VSUBS 0.068049f
C929 VN.n50 VSUBS 0.077792f
C930 VN.n51 VSUBS 0.049949f
C931 VN.n52 VSUBS 0.049949f
C932 VN.n53 VSUBS 0.049949f
C933 VN.n54 VSUBS 0.093092f
C934 VN.n55 VSUBS 0.081142f
C935 VN.n56 VSUBS 0.571961f
C936 VN.n57 VSUBS 0.164956f
C937 VN.n58 VSUBS 0.093954f
C938 VN.t2 VSUBS 0.755826f
C939 VN.n59 VSUBS 0.093092f
C940 VN.n60 VSUBS 0.049949f
C941 VN.n61 VSUBS 0.093092f
C942 VN.n62 VSUBS 0.049949f
C943 VN.t0 VSUBS 0.755826f
C944 VN.n63 VSUBS 0.093092f
C945 VN.n64 VSUBS 0.049949f
C946 VN.n65 VSUBS 0.093092f
C947 VN.n66 VSUBS 0.049949f
C948 VN.t5 VSUBS 0.755826f
C949 VN.n67 VSUBS 0.093092f
C950 VN.n68 VSUBS 0.049949f
C951 VN.n69 VSUBS 0.100288f
C952 VN.n70 VSUBS 0.049949f
C953 VN.t1 VSUBS 0.755826f
C954 VN.n71 VSUBS 0.52589f
C955 VN.t3 VSUBS 1.32554f
C956 VN.n72 VSUBS 0.654773f
C957 VN.n73 VSUBS 0.670847f
C958 VN.n74 VSUBS 0.052647f
C959 VN.n75 VSUBS 0.093092f
C960 VN.n76 VSUBS 0.093092f
C961 VN.n77 VSUBS 0.049949f
C962 VN.n78 VSUBS 0.049949f
C963 VN.n79 VSUBS 0.049949f
C964 VN.n80 VSUBS 0.046488f
C965 VN.n81 VSUBS 0.092158f
C966 VN.n82 VSUBS 0.093092f
C967 VN.n83 VSUBS 0.049949f
C968 VN.n84 VSUBS 0.049949f
C969 VN.n85 VSUBS 0.049949f
C970 VN.n86 VSUBS 0.070112f
C971 VN.n87 VSUBS 0.359804f
C972 VN.n88 VSUBS 0.070112f
C973 VN.n89 VSUBS 0.093092f
C974 VN.n90 VSUBS 0.049949f
C975 VN.n91 VSUBS 0.049949f
C976 VN.n92 VSUBS 0.049949f
C977 VN.n93 VSUBS 0.092158f
C978 VN.n94 VSUBS 0.046488f
C979 VN.n95 VSUBS 0.100288f
C980 VN.n96 VSUBS 0.049949f
C981 VN.n97 VSUBS 0.049949f
C982 VN.n98 VSUBS 0.049949f
C983 VN.n99 VSUBS 0.093092f
C984 VN.n100 VSUBS 0.052647f
C985 VN.n101 VSUBS 0.359804f
C986 VN.n102 VSUBS 0.087577f
C987 VN.n103 VSUBS 0.049949f
C988 VN.n104 VSUBS 0.049949f
C989 VN.n105 VSUBS 0.049949f
C990 VN.n106 VSUBS 0.093092f
C991 VN.n107 VSUBS 0.068049f
C992 VN.n108 VSUBS 0.077792f
C993 VN.n109 VSUBS 0.049949f
C994 VN.n110 VSUBS 0.049949f
C995 VN.n111 VSUBS 0.049949f
C996 VN.n112 VSUBS 0.093092f
C997 VN.n113 VSUBS 0.081142f
C998 VN.n114 VSUBS 0.571961f
C999 VN.n115 VSUBS 3.17079f
C1000 VDD1.t7 VSUBS 0.3717f
C1001 VDD1.t2 VSUBS 0.05871f
C1002 VDD1.t9 VSUBS 0.05871f
C1003 VDD1.n0 VSUBS 0.220745f
C1004 VDD1.n1 VSUBS 2.11883f
C1005 VDD1.t6 VSUBS 0.3717f
C1006 VDD1.t0 VSUBS 0.05871f
C1007 VDD1.t8 VSUBS 0.05871f
C1008 VDD1.n2 VSUBS 0.220744f
C1009 VDD1.n3 VSUBS 2.10391f
C1010 VDD1.t5 VSUBS 0.05871f
C1011 VDD1.t1 VSUBS 0.05871f
C1012 VDD1.n4 VSUBS 0.235651f
C1013 VDD1.n5 VSUBS 5.6581f
C1014 VDD1.t4 VSUBS 0.05871f
C1015 VDD1.t3 VSUBS 0.05871f
C1016 VDD1.n6 VSUBS 0.220745f
C1017 VDD1.n7 VSUBS 5.28187f
C1018 VTAIL.t6 VSUBS 0.054203f
C1019 VTAIL.t19 VSUBS 0.054203f
C1020 VTAIL.n0 VSUBS 0.174707f
C1021 VTAIL.n1 VSUBS 1.0656f
C1022 VTAIL.t9 VSUBS 0.302123f
C1023 VTAIL.n2 VSUBS 1.19988f
C1024 VTAIL.t10 VSUBS 0.054203f
C1025 VTAIL.t8 VSUBS 0.054203f
C1026 VTAIL.n3 VSUBS 0.174707f
C1027 VTAIL.n4 VSUBS 1.36098f
C1028 VTAIL.t11 VSUBS 0.054203f
C1029 VTAIL.t15 VSUBS 0.054203f
C1030 VTAIL.n5 VSUBS 0.174707f
C1031 VTAIL.n6 VSUBS 2.58875f
C1032 VTAIL.t4 VSUBS 0.054203f
C1033 VTAIL.t18 VSUBS 0.054203f
C1034 VTAIL.n7 VSUBS 0.174707f
C1035 VTAIL.n8 VSUBS 2.58875f
C1036 VTAIL.t5 VSUBS 0.054203f
C1037 VTAIL.t2 VSUBS 0.054203f
C1038 VTAIL.n9 VSUBS 0.174707f
C1039 VTAIL.n10 VSUBS 1.36098f
C1040 VTAIL.t1 VSUBS 0.302124f
C1041 VTAIL.n11 VSUBS 1.19988f
C1042 VTAIL.t17 VSUBS 0.054203f
C1043 VTAIL.t16 VSUBS 0.054203f
C1044 VTAIL.n12 VSUBS 0.174707f
C1045 VTAIL.n13 VSUBS 1.17947f
C1046 VTAIL.t12 VSUBS 0.054203f
C1047 VTAIL.t14 VSUBS 0.054203f
C1048 VTAIL.n14 VSUBS 0.174707f
C1049 VTAIL.n15 VSUBS 1.36098f
C1050 VTAIL.t13 VSUBS 0.302124f
C1051 VTAIL.n16 VSUBS 2.12324f
C1052 VTAIL.t3 VSUBS 0.302123f
C1053 VTAIL.n17 VSUBS 2.12325f
C1054 VTAIL.t7 VSUBS 0.054203f
C1055 VTAIL.t0 VSUBS 0.054203f
C1056 VTAIL.n18 VSUBS 0.174707f
C1057 VTAIL.n19 VSUBS 0.988935f
C1058 VP.n0 VSUBS 0.108498f
C1059 VP.t8 VSUBS 0.872834f
C1060 VP.n1 VSUBS 0.107503f
C1061 VP.n2 VSUBS 0.057681f
C1062 VP.n3 VSUBS 0.107503f
C1063 VP.n4 VSUBS 0.057681f
C1064 VP.t4 VSUBS 0.872834f
C1065 VP.n5 VSUBS 0.107503f
C1066 VP.n6 VSUBS 0.057681f
C1067 VP.n7 VSUBS 0.107503f
C1068 VP.n8 VSUBS 0.057681f
C1069 VP.t1 VSUBS 0.872834f
C1070 VP.n9 VSUBS 0.107503f
C1071 VP.n10 VSUBS 0.057681f
C1072 VP.n11 VSUBS 0.115813f
C1073 VP.n12 VSUBS 0.057681f
C1074 VP.t9 VSUBS 0.872834f
C1075 VP.n13 VSUBS 0.415505f
C1076 VP.n14 VSUBS 0.057681f
C1077 VP.n15 VSUBS 0.078584f
C1078 VP.n16 VSUBS 0.057681f
C1079 VP.n17 VSUBS 0.093704f
C1080 VP.n18 VSUBS 0.108498f
C1081 VP.t6 VSUBS 0.872834f
C1082 VP.n19 VSUBS 0.107503f
C1083 VP.n20 VSUBS 0.057681f
C1084 VP.n21 VSUBS 0.107503f
C1085 VP.n22 VSUBS 0.057681f
C1086 VP.t5 VSUBS 0.872834f
C1087 VP.n23 VSUBS 0.107503f
C1088 VP.n24 VSUBS 0.057681f
C1089 VP.n25 VSUBS 0.107503f
C1090 VP.n26 VSUBS 0.057681f
C1091 VP.t0 VSUBS 0.872834f
C1092 VP.n27 VSUBS 0.107503f
C1093 VP.n28 VSUBS 0.057681f
C1094 VP.n29 VSUBS 0.115813f
C1095 VP.n30 VSUBS 0.057681f
C1096 VP.t7 VSUBS 0.872834f
C1097 VP.n31 VSUBS 0.607302f
C1098 VP.t2 VSUBS 1.53074f
C1099 VP.n32 VSUBS 0.756141f
C1100 VP.n33 VSUBS 0.774702f
C1101 VP.n34 VSUBS 0.060797f
C1102 VP.n35 VSUBS 0.107503f
C1103 VP.n36 VSUBS 0.107503f
C1104 VP.n37 VSUBS 0.057681f
C1105 VP.n38 VSUBS 0.057681f
C1106 VP.n39 VSUBS 0.057681f
C1107 VP.n40 VSUBS 0.053684f
C1108 VP.n41 VSUBS 0.106425f
C1109 VP.n42 VSUBS 0.107503f
C1110 VP.n43 VSUBS 0.057681f
C1111 VP.n44 VSUBS 0.057681f
C1112 VP.n45 VSUBS 0.057681f
C1113 VP.n46 VSUBS 0.080966f
C1114 VP.n47 VSUBS 0.415505f
C1115 VP.n48 VSUBS 0.080966f
C1116 VP.n49 VSUBS 0.107503f
C1117 VP.n50 VSUBS 0.057681f
C1118 VP.n51 VSUBS 0.057681f
C1119 VP.n52 VSUBS 0.057681f
C1120 VP.n53 VSUBS 0.106425f
C1121 VP.n54 VSUBS 0.053684f
C1122 VP.n55 VSUBS 0.115813f
C1123 VP.n56 VSUBS 0.057681f
C1124 VP.n57 VSUBS 0.057681f
C1125 VP.n58 VSUBS 0.057681f
C1126 VP.n59 VSUBS 0.107503f
C1127 VP.n60 VSUBS 0.060797f
C1128 VP.n61 VSUBS 0.415505f
C1129 VP.n62 VSUBS 0.101134f
C1130 VP.n63 VSUBS 0.057681f
C1131 VP.n64 VSUBS 0.057681f
C1132 VP.n65 VSUBS 0.057681f
C1133 VP.n66 VSUBS 0.107503f
C1134 VP.n67 VSUBS 0.078584f
C1135 VP.n68 VSUBS 0.089835f
C1136 VP.n69 VSUBS 0.057681f
C1137 VP.n70 VSUBS 0.057681f
C1138 VP.n71 VSUBS 0.057681f
C1139 VP.n72 VSUBS 0.107503f
C1140 VP.n73 VSUBS 0.093704f
C1141 VP.n74 VSUBS 0.660505f
C1142 VP.n75 VSUBS 3.6472f
C1143 VP.t3 VSUBS 0.872834f
C1144 VP.n76 VSUBS 0.660505f
C1145 VP.n77 VSUBS 3.68631f
C1146 VP.n78 VSUBS 0.108498f
C1147 VP.n79 VSUBS 0.057681f
C1148 VP.n80 VSUBS 0.107503f
C1149 VP.n81 VSUBS 0.107503f
C1150 VP.n82 VSUBS 0.089835f
C1151 VP.n83 VSUBS 0.057681f
C1152 VP.n84 VSUBS 0.057681f
C1153 VP.n85 VSUBS 0.057681f
C1154 VP.n86 VSUBS 0.107503f
C1155 VP.n87 VSUBS 0.107503f
C1156 VP.n88 VSUBS 0.101134f
C1157 VP.n89 VSUBS 0.057681f
C1158 VP.n90 VSUBS 0.057681f
C1159 VP.n91 VSUBS 0.060797f
C1160 VP.n92 VSUBS 0.107503f
C1161 VP.n93 VSUBS 0.107503f
C1162 VP.n94 VSUBS 0.057681f
C1163 VP.n95 VSUBS 0.057681f
C1164 VP.n96 VSUBS 0.057681f
C1165 VP.n97 VSUBS 0.053684f
C1166 VP.n98 VSUBS 0.106425f
C1167 VP.n99 VSUBS 0.107503f
C1168 VP.n100 VSUBS 0.057681f
C1169 VP.n101 VSUBS 0.057681f
C1170 VP.n102 VSUBS 0.057681f
C1171 VP.n103 VSUBS 0.080966f
C1172 VP.n104 VSUBS 0.415505f
C1173 VP.n105 VSUBS 0.080966f
C1174 VP.n106 VSUBS 0.107503f
C1175 VP.n107 VSUBS 0.057681f
C1176 VP.n108 VSUBS 0.057681f
C1177 VP.n109 VSUBS 0.057681f
C1178 VP.n110 VSUBS 0.106425f
C1179 VP.n111 VSUBS 0.053684f
C1180 VP.n112 VSUBS 0.115813f
C1181 VP.n113 VSUBS 0.057681f
C1182 VP.n114 VSUBS 0.057681f
C1183 VP.n115 VSUBS 0.057681f
C1184 VP.n116 VSUBS 0.107503f
C1185 VP.n117 VSUBS 0.060797f
C1186 VP.n118 VSUBS 0.415505f
C1187 VP.n119 VSUBS 0.101134f
C1188 VP.n120 VSUBS 0.057681f
C1189 VP.n121 VSUBS 0.057681f
C1190 VP.n122 VSUBS 0.057681f
C1191 VP.n123 VSUBS 0.107503f
C1192 VP.n124 VSUBS 0.078584f
C1193 VP.n125 VSUBS 0.089835f
C1194 VP.n126 VSUBS 0.057681f
C1195 VP.n127 VSUBS 0.057681f
C1196 VP.n128 VSUBS 0.057681f
C1197 VP.n129 VSUBS 0.107503f
C1198 VP.n130 VSUBS 0.093704f
C1199 VP.n131 VSUBS 0.660505f
C1200 VP.n132 VSUBS 0.190492f
.ends

