* NGSPICE file created from diff_pair_sample_1635.ext - technology: sky130A

.subckt diff_pair_sample_1635 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0.37785 ps=2.62 w=2.29 l=1.68
X1 VDD1.t7 VP.t0 VTAIL.t7 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.8931 ps=5.36 w=2.29 l=1.68
X2 VTAIL.t14 VN.t1 VDD2.t0 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
X3 VDD2.t5 VN.t2 VTAIL.t13 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.8931 ps=5.36 w=2.29 l=1.68
X4 B.t11 B.t9 B.t10 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0 ps=0 w=2.29 l=1.68
X5 VDD2.t6 VN.t3 VTAIL.t12 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
X6 VTAIL.t6 VP.t1 VDD1.t6 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
X7 VTAIL.t5 VP.t2 VDD1.t5 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0.37785 ps=2.62 w=2.29 l=1.68
X8 VTAIL.t11 VN.t4 VDD2.t2 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
X9 B.t8 B.t6 B.t7 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0 ps=0 w=2.29 l=1.68
X10 VTAIL.t4 VP.t3 VDD1.t4 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0.37785 ps=2.62 w=2.29 l=1.68
X11 VDD2.t1 VN.t5 VTAIL.t10 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
X12 B.t5 B.t3 B.t4 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0 ps=0 w=2.29 l=1.68
X13 VDD2.t7 VN.t6 VTAIL.t9 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.8931 ps=5.36 w=2.29 l=1.68
X14 B.t2 B.t0 B.t1 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0 ps=0 w=2.29 l=1.68
X15 VDD1.t3 VP.t4 VTAIL.t3 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
X16 VTAIL.t2 VP.t5 VDD1.t2 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
X17 VTAIL.t8 VN.t7 VDD2.t3 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.8931 pd=5.36 as=0.37785 ps=2.62 w=2.29 l=1.68
X18 VDD1.t1 VP.t6 VTAIL.t1 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.8931 ps=5.36 w=2.29 l=1.68
X19 VDD1.t0 VP.t7 VTAIL.t0 w_n2980_n1426# sky130_fd_pr__pfet_01v8 ad=0.37785 pd=2.62 as=0.37785 ps=2.62 w=2.29 l=1.68
R0 VN.n22 VN.n21 185.034
R1 VN.n45 VN.n44 185.034
R2 VN.n43 VN.n23 161.3
R3 VN.n42 VN.n41 161.3
R4 VN.n40 VN.n24 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n36 VN.n25 161.3
R7 VN.n35 VN.n34 161.3
R8 VN.n33 VN.n26 161.3
R9 VN.n32 VN.n31 161.3
R10 VN.n30 VN.n27 161.3
R11 VN.n20 VN.n0 161.3
R12 VN.n19 VN.n18 161.3
R13 VN.n17 VN.n1 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n13 VN.n2 161.3
R16 VN.n12 VN.n11 161.3
R17 VN.n10 VN.n3 161.3
R18 VN.n9 VN.n8 161.3
R19 VN.n7 VN.n4 161.3
R20 VN.n6 VN.n5 68.7155
R21 VN.n29 VN.n28 68.7155
R22 VN.n5 VN.t7 60.3516
R23 VN.n28 VN.t2 60.3516
R24 VN.n19 VN.n1 41.4647
R25 VN.n42 VN.n24 41.4647
R26 VN.n8 VN.n3 40.4934
R27 VN.n12 VN.n3 40.4934
R28 VN.n31 VN.n26 40.4934
R29 VN.n35 VN.n26 40.4934
R30 VN.n15 VN.n1 39.5221
R31 VN.n38 VN.n24 39.5221
R32 VN VN.n45 39.4418
R33 VN.n6 VN.t3 32.8511
R34 VN.n14 VN.t1 32.8511
R35 VN.n21 VN.t6 32.8511
R36 VN.n29 VN.t4 32.8511
R37 VN.n37 VN.t5 32.8511
R38 VN.n44 VN.t0 32.8511
R39 VN.n8 VN.n7 24.4675
R40 VN.n13 VN.n12 24.4675
R41 VN.n20 VN.n19 24.4675
R42 VN.n31 VN.n30 24.4675
R43 VN.n36 VN.n35 24.4675
R44 VN.n43 VN.n42 24.4675
R45 VN.n15 VN.n14 24.2228
R46 VN.n38 VN.n37 24.2228
R47 VN.n28 VN.n27 18.9997
R48 VN.n5 VN.n4 18.9997
R49 VN.n21 VN.n20 0.73451
R50 VN.n44 VN.n43 0.73451
R51 VN.n7 VN.n6 0.24517
R52 VN.n14 VN.n13 0.24517
R53 VN.n30 VN.n29 0.24517
R54 VN.n37 VN.n36 0.24517
R55 VN.n45 VN.n23 0.189894
R56 VN.n41 VN.n23 0.189894
R57 VN.n41 VN.n40 0.189894
R58 VN.n40 VN.n39 0.189894
R59 VN.n39 VN.n25 0.189894
R60 VN.n34 VN.n25 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n32 0.189894
R63 VN.n32 VN.n27 0.189894
R64 VN.n9 VN.n4 0.189894
R65 VN.n10 VN.n9 0.189894
R66 VN.n11 VN.n10 0.189894
R67 VN.n11 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n18 VN.n17 0.189894
R71 VN.n18 VN.n0 0.189894
R72 VN.n22 VN.n0 0.189894
R73 VN VN.n22 0.0516364
R74 VDD2.n2 VDD2.n1 171.194
R75 VDD2.n2 VDD2.n0 171.194
R76 VDD2 VDD2.n5 171.19
R77 VDD2.n4 VDD2.n3 170.382
R78 VDD2.n4 VDD2.n2 33.4868
R79 VDD2.n5 VDD2.t2 14.1948
R80 VDD2.n5 VDD2.t5 14.1948
R81 VDD2.n3 VDD2.t4 14.1948
R82 VDD2.n3 VDD2.t1 14.1948
R83 VDD2.n1 VDD2.t0 14.1948
R84 VDD2.n1 VDD2.t7 14.1948
R85 VDD2.n0 VDD2.t3 14.1948
R86 VDD2.n0 VDD2.t6 14.1948
R87 VDD2 VDD2.n4 0.925069
R88 VTAIL.n11 VTAIL.t4 167.898
R89 VTAIL.n10 VTAIL.t13 167.898
R90 VTAIL.n7 VTAIL.t15 167.898
R91 VTAIL.n14 VTAIL.t7 167.898
R92 VTAIL.n15 VTAIL.t9 167.898
R93 VTAIL.n2 VTAIL.t8 167.898
R94 VTAIL.n3 VTAIL.t1 167.898
R95 VTAIL.n6 VTAIL.t5 167.898
R96 VTAIL.n13 VTAIL.n12 153.703
R97 VTAIL.n9 VTAIL.n8 153.703
R98 VTAIL.n1 VTAIL.n0 153.703
R99 VTAIL.n5 VTAIL.n4 153.703
R100 VTAIL.n15 VTAIL.n14 16.0738
R101 VTAIL.n7 VTAIL.n6 16.0738
R102 VTAIL.n0 VTAIL.t12 14.1948
R103 VTAIL.n0 VTAIL.t14 14.1948
R104 VTAIL.n4 VTAIL.t0 14.1948
R105 VTAIL.n4 VTAIL.t6 14.1948
R106 VTAIL.n12 VTAIL.t3 14.1948
R107 VTAIL.n12 VTAIL.t2 14.1948
R108 VTAIL.n8 VTAIL.t10 14.1948
R109 VTAIL.n8 VTAIL.t11 14.1948
R110 VTAIL.n9 VTAIL.n7 1.73326
R111 VTAIL.n10 VTAIL.n9 1.73326
R112 VTAIL.n13 VTAIL.n11 1.73326
R113 VTAIL.n14 VTAIL.n13 1.73326
R114 VTAIL.n6 VTAIL.n5 1.73326
R115 VTAIL.n5 VTAIL.n3 1.73326
R116 VTAIL.n2 VTAIL.n1 1.73326
R117 VTAIL VTAIL.n15 1.67507
R118 VTAIL.n11 VTAIL.n10 0.470328
R119 VTAIL.n3 VTAIL.n2 0.470328
R120 VTAIL VTAIL.n1 0.0586897
R121 VP.n31 VP.n30 185.034
R122 VP.n54 VP.n53 185.034
R123 VP.n29 VP.n28 185.034
R124 VP.n14 VP.n11 161.3
R125 VP.n16 VP.n15 161.3
R126 VP.n17 VP.n10 161.3
R127 VP.n19 VP.n18 161.3
R128 VP.n20 VP.n9 161.3
R129 VP.n23 VP.n22 161.3
R130 VP.n24 VP.n8 161.3
R131 VP.n26 VP.n25 161.3
R132 VP.n27 VP.n7 161.3
R133 VP.n52 VP.n0 161.3
R134 VP.n51 VP.n50 161.3
R135 VP.n49 VP.n1 161.3
R136 VP.n48 VP.n47 161.3
R137 VP.n45 VP.n2 161.3
R138 VP.n44 VP.n43 161.3
R139 VP.n42 VP.n3 161.3
R140 VP.n41 VP.n40 161.3
R141 VP.n39 VP.n4 161.3
R142 VP.n37 VP.n36 161.3
R143 VP.n35 VP.n5 161.3
R144 VP.n34 VP.n33 161.3
R145 VP.n32 VP.n6 161.3
R146 VP.n13 VP.n12 68.7155
R147 VP.n12 VP.t3 60.3516
R148 VP.n33 VP.n5 41.4647
R149 VP.n51 VP.n1 41.4647
R150 VP.n26 VP.n8 41.4647
R151 VP.n40 VP.n3 40.4934
R152 VP.n44 VP.n3 40.4934
R153 VP.n19 VP.n10 40.4934
R154 VP.n15 VP.n10 40.4934
R155 VP.n37 VP.n5 39.5221
R156 VP.n47 VP.n1 39.5221
R157 VP.n22 VP.n8 39.5221
R158 VP.n30 VP.n29 39.0611
R159 VP.n31 VP.t2 32.8511
R160 VP.n38 VP.t7 32.8511
R161 VP.n46 VP.t1 32.8511
R162 VP.n53 VP.t6 32.8511
R163 VP.n28 VP.t0 32.8511
R164 VP.n21 VP.t5 32.8511
R165 VP.n13 VP.t4 32.8511
R166 VP.n33 VP.n32 24.4675
R167 VP.n40 VP.n39 24.4675
R168 VP.n45 VP.n44 24.4675
R169 VP.n52 VP.n51 24.4675
R170 VP.n27 VP.n26 24.4675
R171 VP.n20 VP.n19 24.4675
R172 VP.n15 VP.n14 24.4675
R173 VP.n38 VP.n37 24.2228
R174 VP.n47 VP.n46 24.2228
R175 VP.n22 VP.n21 24.2228
R176 VP.n12 VP.n11 18.9997
R177 VP.n32 VP.n31 0.73451
R178 VP.n53 VP.n52 0.73451
R179 VP.n28 VP.n27 0.73451
R180 VP.n39 VP.n38 0.24517
R181 VP.n46 VP.n45 0.24517
R182 VP.n21 VP.n20 0.24517
R183 VP.n14 VP.n13 0.24517
R184 VP.n16 VP.n11 0.189894
R185 VP.n17 VP.n16 0.189894
R186 VP.n18 VP.n17 0.189894
R187 VP.n18 VP.n9 0.189894
R188 VP.n23 VP.n9 0.189894
R189 VP.n24 VP.n23 0.189894
R190 VP.n25 VP.n24 0.189894
R191 VP.n25 VP.n7 0.189894
R192 VP.n29 VP.n7 0.189894
R193 VP.n30 VP.n6 0.189894
R194 VP.n34 VP.n6 0.189894
R195 VP.n35 VP.n34 0.189894
R196 VP.n36 VP.n35 0.189894
R197 VP.n36 VP.n4 0.189894
R198 VP.n41 VP.n4 0.189894
R199 VP.n42 VP.n41 0.189894
R200 VP.n43 VP.n42 0.189894
R201 VP.n43 VP.n2 0.189894
R202 VP.n48 VP.n2 0.189894
R203 VP.n49 VP.n48 0.189894
R204 VP.n50 VP.n49 0.189894
R205 VP.n50 VP.n0 0.189894
R206 VP.n54 VP.n0 0.189894
R207 VP VP.n54 0.0516364
R208 VDD1 VDD1.n0 171.306
R209 VDD1.n3 VDD1.n2 171.194
R210 VDD1.n3 VDD1.n1 171.194
R211 VDD1.n5 VDD1.n4 170.382
R212 VDD1.n5 VDD1.n3 34.0699
R213 VDD1.n4 VDD1.t2 14.1948
R214 VDD1.n4 VDD1.t7 14.1948
R215 VDD1.n0 VDD1.t4 14.1948
R216 VDD1.n0 VDD1.t3 14.1948
R217 VDD1.n2 VDD1.t6 14.1948
R218 VDD1.n2 VDD1.t1 14.1948
R219 VDD1.n1 VDD1.t5 14.1948
R220 VDD1.n1 VDD1.t0 14.1948
R221 VDD1 VDD1.n5 0.80869
R222 B.n230 B.n81 585
R223 B.n229 B.n228 585
R224 B.n227 B.n82 585
R225 B.n226 B.n225 585
R226 B.n224 B.n83 585
R227 B.n223 B.n222 585
R228 B.n221 B.n84 585
R229 B.n220 B.n219 585
R230 B.n218 B.n85 585
R231 B.n217 B.n216 585
R232 B.n215 B.n86 585
R233 B.n214 B.n213 585
R234 B.n212 B.n87 585
R235 B.n210 B.n209 585
R236 B.n208 B.n90 585
R237 B.n207 B.n206 585
R238 B.n205 B.n91 585
R239 B.n204 B.n203 585
R240 B.n202 B.n92 585
R241 B.n201 B.n200 585
R242 B.n199 B.n93 585
R243 B.n198 B.n197 585
R244 B.n196 B.n94 585
R245 B.n195 B.n194 585
R246 B.n190 B.n95 585
R247 B.n189 B.n188 585
R248 B.n187 B.n96 585
R249 B.n186 B.n185 585
R250 B.n184 B.n97 585
R251 B.n183 B.n182 585
R252 B.n181 B.n98 585
R253 B.n180 B.n179 585
R254 B.n178 B.n99 585
R255 B.n177 B.n176 585
R256 B.n175 B.n100 585
R257 B.n174 B.n173 585
R258 B.n232 B.n231 585
R259 B.n233 B.n80 585
R260 B.n235 B.n234 585
R261 B.n236 B.n79 585
R262 B.n238 B.n237 585
R263 B.n239 B.n78 585
R264 B.n241 B.n240 585
R265 B.n242 B.n77 585
R266 B.n244 B.n243 585
R267 B.n245 B.n76 585
R268 B.n247 B.n246 585
R269 B.n248 B.n75 585
R270 B.n250 B.n249 585
R271 B.n251 B.n74 585
R272 B.n253 B.n252 585
R273 B.n254 B.n73 585
R274 B.n256 B.n255 585
R275 B.n257 B.n72 585
R276 B.n259 B.n258 585
R277 B.n260 B.n71 585
R278 B.n262 B.n261 585
R279 B.n263 B.n70 585
R280 B.n265 B.n264 585
R281 B.n266 B.n69 585
R282 B.n268 B.n267 585
R283 B.n269 B.n68 585
R284 B.n271 B.n270 585
R285 B.n272 B.n67 585
R286 B.n274 B.n273 585
R287 B.n275 B.n66 585
R288 B.n277 B.n276 585
R289 B.n278 B.n65 585
R290 B.n280 B.n279 585
R291 B.n281 B.n64 585
R292 B.n283 B.n282 585
R293 B.n284 B.n63 585
R294 B.n286 B.n285 585
R295 B.n287 B.n62 585
R296 B.n289 B.n288 585
R297 B.n290 B.n61 585
R298 B.n292 B.n291 585
R299 B.n293 B.n60 585
R300 B.n295 B.n294 585
R301 B.n296 B.n59 585
R302 B.n298 B.n297 585
R303 B.n299 B.n58 585
R304 B.n301 B.n300 585
R305 B.n302 B.n57 585
R306 B.n304 B.n303 585
R307 B.n305 B.n56 585
R308 B.n307 B.n306 585
R309 B.n308 B.n55 585
R310 B.n310 B.n309 585
R311 B.n311 B.n54 585
R312 B.n313 B.n312 585
R313 B.n314 B.n53 585
R314 B.n316 B.n315 585
R315 B.n317 B.n52 585
R316 B.n319 B.n318 585
R317 B.n320 B.n51 585
R318 B.n322 B.n321 585
R319 B.n323 B.n50 585
R320 B.n325 B.n324 585
R321 B.n326 B.n49 585
R322 B.n328 B.n327 585
R323 B.n329 B.n48 585
R324 B.n331 B.n330 585
R325 B.n332 B.n47 585
R326 B.n334 B.n333 585
R327 B.n335 B.n46 585
R328 B.n337 B.n336 585
R329 B.n338 B.n45 585
R330 B.n340 B.n339 585
R331 B.n341 B.n44 585
R332 B.n343 B.n342 585
R333 B.n344 B.n43 585
R334 B.n400 B.n399 585
R335 B.n398 B.n21 585
R336 B.n397 B.n396 585
R337 B.n395 B.n22 585
R338 B.n394 B.n393 585
R339 B.n392 B.n23 585
R340 B.n391 B.n390 585
R341 B.n389 B.n24 585
R342 B.n388 B.n387 585
R343 B.n386 B.n25 585
R344 B.n385 B.n384 585
R345 B.n383 B.n26 585
R346 B.n382 B.n381 585
R347 B.n379 B.n27 585
R348 B.n378 B.n377 585
R349 B.n376 B.n30 585
R350 B.n375 B.n374 585
R351 B.n373 B.n31 585
R352 B.n372 B.n371 585
R353 B.n370 B.n32 585
R354 B.n369 B.n368 585
R355 B.n367 B.n33 585
R356 B.n366 B.n365 585
R357 B.n364 B.n363 585
R358 B.n362 B.n37 585
R359 B.n361 B.n360 585
R360 B.n359 B.n38 585
R361 B.n358 B.n357 585
R362 B.n356 B.n39 585
R363 B.n355 B.n354 585
R364 B.n353 B.n40 585
R365 B.n352 B.n351 585
R366 B.n350 B.n41 585
R367 B.n349 B.n348 585
R368 B.n347 B.n42 585
R369 B.n346 B.n345 585
R370 B.n401 B.n20 585
R371 B.n403 B.n402 585
R372 B.n404 B.n19 585
R373 B.n406 B.n405 585
R374 B.n407 B.n18 585
R375 B.n409 B.n408 585
R376 B.n410 B.n17 585
R377 B.n412 B.n411 585
R378 B.n413 B.n16 585
R379 B.n415 B.n414 585
R380 B.n416 B.n15 585
R381 B.n418 B.n417 585
R382 B.n419 B.n14 585
R383 B.n421 B.n420 585
R384 B.n422 B.n13 585
R385 B.n424 B.n423 585
R386 B.n425 B.n12 585
R387 B.n427 B.n426 585
R388 B.n428 B.n11 585
R389 B.n430 B.n429 585
R390 B.n431 B.n10 585
R391 B.n433 B.n432 585
R392 B.n434 B.n9 585
R393 B.n436 B.n435 585
R394 B.n437 B.n8 585
R395 B.n439 B.n438 585
R396 B.n440 B.n7 585
R397 B.n442 B.n441 585
R398 B.n443 B.n6 585
R399 B.n445 B.n444 585
R400 B.n446 B.n5 585
R401 B.n448 B.n447 585
R402 B.n449 B.n4 585
R403 B.n451 B.n450 585
R404 B.n452 B.n3 585
R405 B.n454 B.n453 585
R406 B.n455 B.n0 585
R407 B.n2 B.n1 585
R408 B.n120 B.n119 585
R409 B.n121 B.n118 585
R410 B.n123 B.n122 585
R411 B.n124 B.n117 585
R412 B.n126 B.n125 585
R413 B.n127 B.n116 585
R414 B.n129 B.n128 585
R415 B.n130 B.n115 585
R416 B.n132 B.n131 585
R417 B.n133 B.n114 585
R418 B.n135 B.n134 585
R419 B.n136 B.n113 585
R420 B.n138 B.n137 585
R421 B.n139 B.n112 585
R422 B.n141 B.n140 585
R423 B.n142 B.n111 585
R424 B.n144 B.n143 585
R425 B.n145 B.n110 585
R426 B.n147 B.n146 585
R427 B.n148 B.n109 585
R428 B.n150 B.n149 585
R429 B.n151 B.n108 585
R430 B.n153 B.n152 585
R431 B.n154 B.n107 585
R432 B.n156 B.n155 585
R433 B.n157 B.n106 585
R434 B.n159 B.n158 585
R435 B.n160 B.n105 585
R436 B.n162 B.n161 585
R437 B.n163 B.n104 585
R438 B.n165 B.n164 585
R439 B.n166 B.n103 585
R440 B.n168 B.n167 585
R441 B.n169 B.n102 585
R442 B.n171 B.n170 585
R443 B.n172 B.n101 585
R444 B.n174 B.n101 502.111
R445 B.n232 B.n81 502.111
R446 B.n346 B.n43 502.111
R447 B.n401 B.n400 502.111
R448 B.n457 B.n456 256.663
R449 B.n191 B.t3 238.904
R450 B.n88 B.t0 238.904
R451 B.n34 B.t9 238.904
R452 B.n28 B.t6 238.904
R453 B.n456 B.n455 235.042
R454 B.n456 B.n2 235.042
R455 B.n88 B.t1 212.994
R456 B.n34 B.t11 212.994
R457 B.n191 B.t4 212.994
R458 B.n28 B.t8 212.994
R459 B.n89 B.t2 174.012
R460 B.n35 B.t10 174.012
R461 B.n192 B.t5 174.012
R462 B.n29 B.t7 174.012
R463 B.n175 B.n174 163.367
R464 B.n176 B.n175 163.367
R465 B.n176 B.n99 163.367
R466 B.n180 B.n99 163.367
R467 B.n181 B.n180 163.367
R468 B.n182 B.n181 163.367
R469 B.n182 B.n97 163.367
R470 B.n186 B.n97 163.367
R471 B.n187 B.n186 163.367
R472 B.n188 B.n187 163.367
R473 B.n188 B.n95 163.367
R474 B.n195 B.n95 163.367
R475 B.n196 B.n195 163.367
R476 B.n197 B.n196 163.367
R477 B.n197 B.n93 163.367
R478 B.n201 B.n93 163.367
R479 B.n202 B.n201 163.367
R480 B.n203 B.n202 163.367
R481 B.n203 B.n91 163.367
R482 B.n207 B.n91 163.367
R483 B.n208 B.n207 163.367
R484 B.n209 B.n208 163.367
R485 B.n209 B.n87 163.367
R486 B.n214 B.n87 163.367
R487 B.n215 B.n214 163.367
R488 B.n216 B.n215 163.367
R489 B.n216 B.n85 163.367
R490 B.n220 B.n85 163.367
R491 B.n221 B.n220 163.367
R492 B.n222 B.n221 163.367
R493 B.n222 B.n83 163.367
R494 B.n226 B.n83 163.367
R495 B.n227 B.n226 163.367
R496 B.n228 B.n227 163.367
R497 B.n228 B.n81 163.367
R498 B.n342 B.n43 163.367
R499 B.n342 B.n341 163.367
R500 B.n341 B.n340 163.367
R501 B.n340 B.n45 163.367
R502 B.n336 B.n45 163.367
R503 B.n336 B.n335 163.367
R504 B.n335 B.n334 163.367
R505 B.n334 B.n47 163.367
R506 B.n330 B.n47 163.367
R507 B.n330 B.n329 163.367
R508 B.n329 B.n328 163.367
R509 B.n328 B.n49 163.367
R510 B.n324 B.n49 163.367
R511 B.n324 B.n323 163.367
R512 B.n323 B.n322 163.367
R513 B.n322 B.n51 163.367
R514 B.n318 B.n51 163.367
R515 B.n318 B.n317 163.367
R516 B.n317 B.n316 163.367
R517 B.n316 B.n53 163.367
R518 B.n312 B.n53 163.367
R519 B.n312 B.n311 163.367
R520 B.n311 B.n310 163.367
R521 B.n310 B.n55 163.367
R522 B.n306 B.n55 163.367
R523 B.n306 B.n305 163.367
R524 B.n305 B.n304 163.367
R525 B.n304 B.n57 163.367
R526 B.n300 B.n57 163.367
R527 B.n300 B.n299 163.367
R528 B.n299 B.n298 163.367
R529 B.n298 B.n59 163.367
R530 B.n294 B.n59 163.367
R531 B.n294 B.n293 163.367
R532 B.n293 B.n292 163.367
R533 B.n292 B.n61 163.367
R534 B.n288 B.n61 163.367
R535 B.n288 B.n287 163.367
R536 B.n287 B.n286 163.367
R537 B.n286 B.n63 163.367
R538 B.n282 B.n63 163.367
R539 B.n282 B.n281 163.367
R540 B.n281 B.n280 163.367
R541 B.n280 B.n65 163.367
R542 B.n276 B.n65 163.367
R543 B.n276 B.n275 163.367
R544 B.n275 B.n274 163.367
R545 B.n274 B.n67 163.367
R546 B.n270 B.n67 163.367
R547 B.n270 B.n269 163.367
R548 B.n269 B.n268 163.367
R549 B.n268 B.n69 163.367
R550 B.n264 B.n69 163.367
R551 B.n264 B.n263 163.367
R552 B.n263 B.n262 163.367
R553 B.n262 B.n71 163.367
R554 B.n258 B.n71 163.367
R555 B.n258 B.n257 163.367
R556 B.n257 B.n256 163.367
R557 B.n256 B.n73 163.367
R558 B.n252 B.n73 163.367
R559 B.n252 B.n251 163.367
R560 B.n251 B.n250 163.367
R561 B.n250 B.n75 163.367
R562 B.n246 B.n75 163.367
R563 B.n246 B.n245 163.367
R564 B.n245 B.n244 163.367
R565 B.n244 B.n77 163.367
R566 B.n240 B.n77 163.367
R567 B.n240 B.n239 163.367
R568 B.n239 B.n238 163.367
R569 B.n238 B.n79 163.367
R570 B.n234 B.n79 163.367
R571 B.n234 B.n233 163.367
R572 B.n233 B.n232 163.367
R573 B.n400 B.n21 163.367
R574 B.n396 B.n21 163.367
R575 B.n396 B.n395 163.367
R576 B.n395 B.n394 163.367
R577 B.n394 B.n23 163.367
R578 B.n390 B.n23 163.367
R579 B.n390 B.n389 163.367
R580 B.n389 B.n388 163.367
R581 B.n388 B.n25 163.367
R582 B.n384 B.n25 163.367
R583 B.n384 B.n383 163.367
R584 B.n383 B.n382 163.367
R585 B.n382 B.n27 163.367
R586 B.n377 B.n27 163.367
R587 B.n377 B.n376 163.367
R588 B.n376 B.n375 163.367
R589 B.n375 B.n31 163.367
R590 B.n371 B.n31 163.367
R591 B.n371 B.n370 163.367
R592 B.n370 B.n369 163.367
R593 B.n369 B.n33 163.367
R594 B.n365 B.n33 163.367
R595 B.n365 B.n364 163.367
R596 B.n364 B.n37 163.367
R597 B.n360 B.n37 163.367
R598 B.n360 B.n359 163.367
R599 B.n359 B.n358 163.367
R600 B.n358 B.n39 163.367
R601 B.n354 B.n39 163.367
R602 B.n354 B.n353 163.367
R603 B.n353 B.n352 163.367
R604 B.n352 B.n41 163.367
R605 B.n348 B.n41 163.367
R606 B.n348 B.n347 163.367
R607 B.n347 B.n346 163.367
R608 B.n402 B.n401 163.367
R609 B.n402 B.n19 163.367
R610 B.n406 B.n19 163.367
R611 B.n407 B.n406 163.367
R612 B.n408 B.n407 163.367
R613 B.n408 B.n17 163.367
R614 B.n412 B.n17 163.367
R615 B.n413 B.n412 163.367
R616 B.n414 B.n413 163.367
R617 B.n414 B.n15 163.367
R618 B.n418 B.n15 163.367
R619 B.n419 B.n418 163.367
R620 B.n420 B.n419 163.367
R621 B.n420 B.n13 163.367
R622 B.n424 B.n13 163.367
R623 B.n425 B.n424 163.367
R624 B.n426 B.n425 163.367
R625 B.n426 B.n11 163.367
R626 B.n430 B.n11 163.367
R627 B.n431 B.n430 163.367
R628 B.n432 B.n431 163.367
R629 B.n432 B.n9 163.367
R630 B.n436 B.n9 163.367
R631 B.n437 B.n436 163.367
R632 B.n438 B.n437 163.367
R633 B.n438 B.n7 163.367
R634 B.n442 B.n7 163.367
R635 B.n443 B.n442 163.367
R636 B.n444 B.n443 163.367
R637 B.n444 B.n5 163.367
R638 B.n448 B.n5 163.367
R639 B.n449 B.n448 163.367
R640 B.n450 B.n449 163.367
R641 B.n450 B.n3 163.367
R642 B.n454 B.n3 163.367
R643 B.n455 B.n454 163.367
R644 B.n120 B.n2 163.367
R645 B.n121 B.n120 163.367
R646 B.n122 B.n121 163.367
R647 B.n122 B.n117 163.367
R648 B.n126 B.n117 163.367
R649 B.n127 B.n126 163.367
R650 B.n128 B.n127 163.367
R651 B.n128 B.n115 163.367
R652 B.n132 B.n115 163.367
R653 B.n133 B.n132 163.367
R654 B.n134 B.n133 163.367
R655 B.n134 B.n113 163.367
R656 B.n138 B.n113 163.367
R657 B.n139 B.n138 163.367
R658 B.n140 B.n139 163.367
R659 B.n140 B.n111 163.367
R660 B.n144 B.n111 163.367
R661 B.n145 B.n144 163.367
R662 B.n146 B.n145 163.367
R663 B.n146 B.n109 163.367
R664 B.n150 B.n109 163.367
R665 B.n151 B.n150 163.367
R666 B.n152 B.n151 163.367
R667 B.n152 B.n107 163.367
R668 B.n156 B.n107 163.367
R669 B.n157 B.n156 163.367
R670 B.n158 B.n157 163.367
R671 B.n158 B.n105 163.367
R672 B.n162 B.n105 163.367
R673 B.n163 B.n162 163.367
R674 B.n164 B.n163 163.367
R675 B.n164 B.n103 163.367
R676 B.n168 B.n103 163.367
R677 B.n169 B.n168 163.367
R678 B.n170 B.n169 163.367
R679 B.n170 B.n101 163.367
R680 B.n193 B.n192 59.5399
R681 B.n211 B.n89 59.5399
R682 B.n36 B.n35 59.5399
R683 B.n380 B.n29 59.5399
R684 B.n192 B.n191 38.9823
R685 B.n89 B.n88 38.9823
R686 B.n35 B.n34 38.9823
R687 B.n29 B.n28 38.9823
R688 B.n399 B.n20 32.6249
R689 B.n345 B.n344 32.6249
R690 B.n231 B.n230 32.6249
R691 B.n173 B.n172 32.6249
R692 B B.n457 18.0485
R693 B.n403 B.n20 10.6151
R694 B.n404 B.n403 10.6151
R695 B.n405 B.n404 10.6151
R696 B.n405 B.n18 10.6151
R697 B.n409 B.n18 10.6151
R698 B.n410 B.n409 10.6151
R699 B.n411 B.n410 10.6151
R700 B.n411 B.n16 10.6151
R701 B.n415 B.n16 10.6151
R702 B.n416 B.n415 10.6151
R703 B.n417 B.n416 10.6151
R704 B.n417 B.n14 10.6151
R705 B.n421 B.n14 10.6151
R706 B.n422 B.n421 10.6151
R707 B.n423 B.n422 10.6151
R708 B.n423 B.n12 10.6151
R709 B.n427 B.n12 10.6151
R710 B.n428 B.n427 10.6151
R711 B.n429 B.n428 10.6151
R712 B.n429 B.n10 10.6151
R713 B.n433 B.n10 10.6151
R714 B.n434 B.n433 10.6151
R715 B.n435 B.n434 10.6151
R716 B.n435 B.n8 10.6151
R717 B.n439 B.n8 10.6151
R718 B.n440 B.n439 10.6151
R719 B.n441 B.n440 10.6151
R720 B.n441 B.n6 10.6151
R721 B.n445 B.n6 10.6151
R722 B.n446 B.n445 10.6151
R723 B.n447 B.n446 10.6151
R724 B.n447 B.n4 10.6151
R725 B.n451 B.n4 10.6151
R726 B.n452 B.n451 10.6151
R727 B.n453 B.n452 10.6151
R728 B.n453 B.n0 10.6151
R729 B.n399 B.n398 10.6151
R730 B.n398 B.n397 10.6151
R731 B.n397 B.n22 10.6151
R732 B.n393 B.n22 10.6151
R733 B.n393 B.n392 10.6151
R734 B.n392 B.n391 10.6151
R735 B.n391 B.n24 10.6151
R736 B.n387 B.n24 10.6151
R737 B.n387 B.n386 10.6151
R738 B.n386 B.n385 10.6151
R739 B.n385 B.n26 10.6151
R740 B.n381 B.n26 10.6151
R741 B.n379 B.n378 10.6151
R742 B.n378 B.n30 10.6151
R743 B.n374 B.n30 10.6151
R744 B.n374 B.n373 10.6151
R745 B.n373 B.n372 10.6151
R746 B.n372 B.n32 10.6151
R747 B.n368 B.n32 10.6151
R748 B.n368 B.n367 10.6151
R749 B.n367 B.n366 10.6151
R750 B.n363 B.n362 10.6151
R751 B.n362 B.n361 10.6151
R752 B.n361 B.n38 10.6151
R753 B.n357 B.n38 10.6151
R754 B.n357 B.n356 10.6151
R755 B.n356 B.n355 10.6151
R756 B.n355 B.n40 10.6151
R757 B.n351 B.n40 10.6151
R758 B.n351 B.n350 10.6151
R759 B.n350 B.n349 10.6151
R760 B.n349 B.n42 10.6151
R761 B.n345 B.n42 10.6151
R762 B.n344 B.n343 10.6151
R763 B.n343 B.n44 10.6151
R764 B.n339 B.n44 10.6151
R765 B.n339 B.n338 10.6151
R766 B.n338 B.n337 10.6151
R767 B.n337 B.n46 10.6151
R768 B.n333 B.n46 10.6151
R769 B.n333 B.n332 10.6151
R770 B.n332 B.n331 10.6151
R771 B.n331 B.n48 10.6151
R772 B.n327 B.n48 10.6151
R773 B.n327 B.n326 10.6151
R774 B.n326 B.n325 10.6151
R775 B.n325 B.n50 10.6151
R776 B.n321 B.n50 10.6151
R777 B.n321 B.n320 10.6151
R778 B.n320 B.n319 10.6151
R779 B.n319 B.n52 10.6151
R780 B.n315 B.n52 10.6151
R781 B.n315 B.n314 10.6151
R782 B.n314 B.n313 10.6151
R783 B.n313 B.n54 10.6151
R784 B.n309 B.n54 10.6151
R785 B.n309 B.n308 10.6151
R786 B.n308 B.n307 10.6151
R787 B.n307 B.n56 10.6151
R788 B.n303 B.n56 10.6151
R789 B.n303 B.n302 10.6151
R790 B.n302 B.n301 10.6151
R791 B.n301 B.n58 10.6151
R792 B.n297 B.n58 10.6151
R793 B.n297 B.n296 10.6151
R794 B.n296 B.n295 10.6151
R795 B.n295 B.n60 10.6151
R796 B.n291 B.n60 10.6151
R797 B.n291 B.n290 10.6151
R798 B.n290 B.n289 10.6151
R799 B.n289 B.n62 10.6151
R800 B.n285 B.n62 10.6151
R801 B.n285 B.n284 10.6151
R802 B.n284 B.n283 10.6151
R803 B.n283 B.n64 10.6151
R804 B.n279 B.n64 10.6151
R805 B.n279 B.n278 10.6151
R806 B.n278 B.n277 10.6151
R807 B.n277 B.n66 10.6151
R808 B.n273 B.n66 10.6151
R809 B.n273 B.n272 10.6151
R810 B.n272 B.n271 10.6151
R811 B.n271 B.n68 10.6151
R812 B.n267 B.n68 10.6151
R813 B.n267 B.n266 10.6151
R814 B.n266 B.n265 10.6151
R815 B.n265 B.n70 10.6151
R816 B.n261 B.n70 10.6151
R817 B.n261 B.n260 10.6151
R818 B.n260 B.n259 10.6151
R819 B.n259 B.n72 10.6151
R820 B.n255 B.n72 10.6151
R821 B.n255 B.n254 10.6151
R822 B.n254 B.n253 10.6151
R823 B.n253 B.n74 10.6151
R824 B.n249 B.n74 10.6151
R825 B.n249 B.n248 10.6151
R826 B.n248 B.n247 10.6151
R827 B.n247 B.n76 10.6151
R828 B.n243 B.n76 10.6151
R829 B.n243 B.n242 10.6151
R830 B.n242 B.n241 10.6151
R831 B.n241 B.n78 10.6151
R832 B.n237 B.n78 10.6151
R833 B.n237 B.n236 10.6151
R834 B.n236 B.n235 10.6151
R835 B.n235 B.n80 10.6151
R836 B.n231 B.n80 10.6151
R837 B.n119 B.n1 10.6151
R838 B.n119 B.n118 10.6151
R839 B.n123 B.n118 10.6151
R840 B.n124 B.n123 10.6151
R841 B.n125 B.n124 10.6151
R842 B.n125 B.n116 10.6151
R843 B.n129 B.n116 10.6151
R844 B.n130 B.n129 10.6151
R845 B.n131 B.n130 10.6151
R846 B.n131 B.n114 10.6151
R847 B.n135 B.n114 10.6151
R848 B.n136 B.n135 10.6151
R849 B.n137 B.n136 10.6151
R850 B.n137 B.n112 10.6151
R851 B.n141 B.n112 10.6151
R852 B.n142 B.n141 10.6151
R853 B.n143 B.n142 10.6151
R854 B.n143 B.n110 10.6151
R855 B.n147 B.n110 10.6151
R856 B.n148 B.n147 10.6151
R857 B.n149 B.n148 10.6151
R858 B.n149 B.n108 10.6151
R859 B.n153 B.n108 10.6151
R860 B.n154 B.n153 10.6151
R861 B.n155 B.n154 10.6151
R862 B.n155 B.n106 10.6151
R863 B.n159 B.n106 10.6151
R864 B.n160 B.n159 10.6151
R865 B.n161 B.n160 10.6151
R866 B.n161 B.n104 10.6151
R867 B.n165 B.n104 10.6151
R868 B.n166 B.n165 10.6151
R869 B.n167 B.n166 10.6151
R870 B.n167 B.n102 10.6151
R871 B.n171 B.n102 10.6151
R872 B.n172 B.n171 10.6151
R873 B.n173 B.n100 10.6151
R874 B.n177 B.n100 10.6151
R875 B.n178 B.n177 10.6151
R876 B.n179 B.n178 10.6151
R877 B.n179 B.n98 10.6151
R878 B.n183 B.n98 10.6151
R879 B.n184 B.n183 10.6151
R880 B.n185 B.n184 10.6151
R881 B.n185 B.n96 10.6151
R882 B.n189 B.n96 10.6151
R883 B.n190 B.n189 10.6151
R884 B.n194 B.n190 10.6151
R885 B.n198 B.n94 10.6151
R886 B.n199 B.n198 10.6151
R887 B.n200 B.n199 10.6151
R888 B.n200 B.n92 10.6151
R889 B.n204 B.n92 10.6151
R890 B.n205 B.n204 10.6151
R891 B.n206 B.n205 10.6151
R892 B.n206 B.n90 10.6151
R893 B.n210 B.n90 10.6151
R894 B.n213 B.n212 10.6151
R895 B.n213 B.n86 10.6151
R896 B.n217 B.n86 10.6151
R897 B.n218 B.n217 10.6151
R898 B.n219 B.n218 10.6151
R899 B.n219 B.n84 10.6151
R900 B.n223 B.n84 10.6151
R901 B.n224 B.n223 10.6151
R902 B.n225 B.n224 10.6151
R903 B.n225 B.n82 10.6151
R904 B.n229 B.n82 10.6151
R905 B.n230 B.n229 10.6151
R906 B.n381 B.n380 9.36635
R907 B.n363 B.n36 9.36635
R908 B.n194 B.n193 9.36635
R909 B.n212 B.n211 9.36635
R910 B.n457 B.n0 8.11757
R911 B.n457 B.n1 8.11757
R912 B.n380 B.n379 1.24928
R913 B.n366 B.n36 1.24928
R914 B.n193 B.n94 1.24928
R915 B.n211 B.n210 1.24928
C0 w_n2980_n1426# VP 6.01475f
C1 VTAIL VDD2 4.13616f
C2 B VDD2 1.17415f
C3 VN VDD2 1.85084f
C4 VTAIL VP 2.54643f
C5 VTAIL w_n2980_n1426# 1.84512f
C6 B VP 1.53299f
C7 B w_n2980_n1426# 6.00306f
C8 VDD1 VDD2 1.29537f
C9 VN VP 4.749629f
C10 VN w_n2980_n1426# 5.63423f
C11 VDD1 VP 2.12149f
C12 VDD1 w_n2980_n1426# 1.38048f
C13 VTAIL B 1.47484f
C14 VTAIL VN 2.53232f
C15 VN B 0.89456f
C16 VDD1 VTAIL 4.08791f
C17 VDD2 VP 0.427676f
C18 w_n2980_n1426# VDD2 1.45593f
C19 VDD1 B 1.10683f
C20 VDD1 VN 0.155112f
C21 VDD2 VSUBS 0.947887f
C22 VDD1 VSUBS 1.636885f
C23 VTAIL VSUBS 0.451869f
C24 VN VSUBS 5.09105f
C25 VP VSUBS 2.080152f
C26 B VSUBS 2.980108f
C27 w_n2980_n1426# VSUBS 54.104897f
C28 B.n0 VSUBS 0.007361f
C29 B.n1 VSUBS 0.007361f
C30 B.n2 VSUBS 0.010886f
C31 B.n3 VSUBS 0.008342f
C32 B.n4 VSUBS 0.008342f
C33 B.n5 VSUBS 0.008342f
C34 B.n6 VSUBS 0.008342f
C35 B.n7 VSUBS 0.008342f
C36 B.n8 VSUBS 0.008342f
C37 B.n9 VSUBS 0.008342f
C38 B.n10 VSUBS 0.008342f
C39 B.n11 VSUBS 0.008342f
C40 B.n12 VSUBS 0.008342f
C41 B.n13 VSUBS 0.008342f
C42 B.n14 VSUBS 0.008342f
C43 B.n15 VSUBS 0.008342f
C44 B.n16 VSUBS 0.008342f
C45 B.n17 VSUBS 0.008342f
C46 B.n18 VSUBS 0.008342f
C47 B.n19 VSUBS 0.008342f
C48 B.n20 VSUBS 0.018773f
C49 B.n21 VSUBS 0.008342f
C50 B.n22 VSUBS 0.008342f
C51 B.n23 VSUBS 0.008342f
C52 B.n24 VSUBS 0.008342f
C53 B.n25 VSUBS 0.008342f
C54 B.n26 VSUBS 0.008342f
C55 B.n27 VSUBS 0.008342f
C56 B.t7 VSUBS 0.060626f
C57 B.t8 VSUBS 0.070906f
C58 B.t6 VSUBS 0.222655f
C59 B.n28 VSUBS 0.079835f
C60 B.n29 VSUBS 0.068066f
C61 B.n30 VSUBS 0.008342f
C62 B.n31 VSUBS 0.008342f
C63 B.n32 VSUBS 0.008342f
C64 B.n33 VSUBS 0.008342f
C65 B.t10 VSUBS 0.060626f
C66 B.t11 VSUBS 0.070906f
C67 B.t9 VSUBS 0.222655f
C68 B.n34 VSUBS 0.079835f
C69 B.n35 VSUBS 0.068066f
C70 B.n36 VSUBS 0.019329f
C71 B.n37 VSUBS 0.008342f
C72 B.n38 VSUBS 0.008342f
C73 B.n39 VSUBS 0.008342f
C74 B.n40 VSUBS 0.008342f
C75 B.n41 VSUBS 0.008342f
C76 B.n42 VSUBS 0.008342f
C77 B.n43 VSUBS 0.018773f
C78 B.n44 VSUBS 0.008342f
C79 B.n45 VSUBS 0.008342f
C80 B.n46 VSUBS 0.008342f
C81 B.n47 VSUBS 0.008342f
C82 B.n48 VSUBS 0.008342f
C83 B.n49 VSUBS 0.008342f
C84 B.n50 VSUBS 0.008342f
C85 B.n51 VSUBS 0.008342f
C86 B.n52 VSUBS 0.008342f
C87 B.n53 VSUBS 0.008342f
C88 B.n54 VSUBS 0.008342f
C89 B.n55 VSUBS 0.008342f
C90 B.n56 VSUBS 0.008342f
C91 B.n57 VSUBS 0.008342f
C92 B.n58 VSUBS 0.008342f
C93 B.n59 VSUBS 0.008342f
C94 B.n60 VSUBS 0.008342f
C95 B.n61 VSUBS 0.008342f
C96 B.n62 VSUBS 0.008342f
C97 B.n63 VSUBS 0.008342f
C98 B.n64 VSUBS 0.008342f
C99 B.n65 VSUBS 0.008342f
C100 B.n66 VSUBS 0.008342f
C101 B.n67 VSUBS 0.008342f
C102 B.n68 VSUBS 0.008342f
C103 B.n69 VSUBS 0.008342f
C104 B.n70 VSUBS 0.008342f
C105 B.n71 VSUBS 0.008342f
C106 B.n72 VSUBS 0.008342f
C107 B.n73 VSUBS 0.008342f
C108 B.n74 VSUBS 0.008342f
C109 B.n75 VSUBS 0.008342f
C110 B.n76 VSUBS 0.008342f
C111 B.n77 VSUBS 0.008342f
C112 B.n78 VSUBS 0.008342f
C113 B.n79 VSUBS 0.008342f
C114 B.n80 VSUBS 0.008342f
C115 B.n81 VSUBS 0.020241f
C116 B.n82 VSUBS 0.008342f
C117 B.n83 VSUBS 0.008342f
C118 B.n84 VSUBS 0.008342f
C119 B.n85 VSUBS 0.008342f
C120 B.n86 VSUBS 0.008342f
C121 B.n87 VSUBS 0.008342f
C122 B.t2 VSUBS 0.060626f
C123 B.t1 VSUBS 0.070906f
C124 B.t0 VSUBS 0.222655f
C125 B.n88 VSUBS 0.079835f
C126 B.n89 VSUBS 0.068066f
C127 B.n90 VSUBS 0.008342f
C128 B.n91 VSUBS 0.008342f
C129 B.n92 VSUBS 0.008342f
C130 B.n93 VSUBS 0.008342f
C131 B.n94 VSUBS 0.004662f
C132 B.n95 VSUBS 0.008342f
C133 B.n96 VSUBS 0.008342f
C134 B.n97 VSUBS 0.008342f
C135 B.n98 VSUBS 0.008342f
C136 B.n99 VSUBS 0.008342f
C137 B.n100 VSUBS 0.008342f
C138 B.n101 VSUBS 0.018773f
C139 B.n102 VSUBS 0.008342f
C140 B.n103 VSUBS 0.008342f
C141 B.n104 VSUBS 0.008342f
C142 B.n105 VSUBS 0.008342f
C143 B.n106 VSUBS 0.008342f
C144 B.n107 VSUBS 0.008342f
C145 B.n108 VSUBS 0.008342f
C146 B.n109 VSUBS 0.008342f
C147 B.n110 VSUBS 0.008342f
C148 B.n111 VSUBS 0.008342f
C149 B.n112 VSUBS 0.008342f
C150 B.n113 VSUBS 0.008342f
C151 B.n114 VSUBS 0.008342f
C152 B.n115 VSUBS 0.008342f
C153 B.n116 VSUBS 0.008342f
C154 B.n117 VSUBS 0.008342f
C155 B.n118 VSUBS 0.008342f
C156 B.n119 VSUBS 0.008342f
C157 B.n120 VSUBS 0.008342f
C158 B.n121 VSUBS 0.008342f
C159 B.n122 VSUBS 0.008342f
C160 B.n123 VSUBS 0.008342f
C161 B.n124 VSUBS 0.008342f
C162 B.n125 VSUBS 0.008342f
C163 B.n126 VSUBS 0.008342f
C164 B.n127 VSUBS 0.008342f
C165 B.n128 VSUBS 0.008342f
C166 B.n129 VSUBS 0.008342f
C167 B.n130 VSUBS 0.008342f
C168 B.n131 VSUBS 0.008342f
C169 B.n132 VSUBS 0.008342f
C170 B.n133 VSUBS 0.008342f
C171 B.n134 VSUBS 0.008342f
C172 B.n135 VSUBS 0.008342f
C173 B.n136 VSUBS 0.008342f
C174 B.n137 VSUBS 0.008342f
C175 B.n138 VSUBS 0.008342f
C176 B.n139 VSUBS 0.008342f
C177 B.n140 VSUBS 0.008342f
C178 B.n141 VSUBS 0.008342f
C179 B.n142 VSUBS 0.008342f
C180 B.n143 VSUBS 0.008342f
C181 B.n144 VSUBS 0.008342f
C182 B.n145 VSUBS 0.008342f
C183 B.n146 VSUBS 0.008342f
C184 B.n147 VSUBS 0.008342f
C185 B.n148 VSUBS 0.008342f
C186 B.n149 VSUBS 0.008342f
C187 B.n150 VSUBS 0.008342f
C188 B.n151 VSUBS 0.008342f
C189 B.n152 VSUBS 0.008342f
C190 B.n153 VSUBS 0.008342f
C191 B.n154 VSUBS 0.008342f
C192 B.n155 VSUBS 0.008342f
C193 B.n156 VSUBS 0.008342f
C194 B.n157 VSUBS 0.008342f
C195 B.n158 VSUBS 0.008342f
C196 B.n159 VSUBS 0.008342f
C197 B.n160 VSUBS 0.008342f
C198 B.n161 VSUBS 0.008342f
C199 B.n162 VSUBS 0.008342f
C200 B.n163 VSUBS 0.008342f
C201 B.n164 VSUBS 0.008342f
C202 B.n165 VSUBS 0.008342f
C203 B.n166 VSUBS 0.008342f
C204 B.n167 VSUBS 0.008342f
C205 B.n168 VSUBS 0.008342f
C206 B.n169 VSUBS 0.008342f
C207 B.n170 VSUBS 0.008342f
C208 B.n171 VSUBS 0.008342f
C209 B.n172 VSUBS 0.018773f
C210 B.n173 VSUBS 0.020241f
C211 B.n174 VSUBS 0.020241f
C212 B.n175 VSUBS 0.008342f
C213 B.n176 VSUBS 0.008342f
C214 B.n177 VSUBS 0.008342f
C215 B.n178 VSUBS 0.008342f
C216 B.n179 VSUBS 0.008342f
C217 B.n180 VSUBS 0.008342f
C218 B.n181 VSUBS 0.008342f
C219 B.n182 VSUBS 0.008342f
C220 B.n183 VSUBS 0.008342f
C221 B.n184 VSUBS 0.008342f
C222 B.n185 VSUBS 0.008342f
C223 B.n186 VSUBS 0.008342f
C224 B.n187 VSUBS 0.008342f
C225 B.n188 VSUBS 0.008342f
C226 B.n189 VSUBS 0.008342f
C227 B.n190 VSUBS 0.008342f
C228 B.t5 VSUBS 0.060626f
C229 B.t4 VSUBS 0.070906f
C230 B.t3 VSUBS 0.222655f
C231 B.n191 VSUBS 0.079835f
C232 B.n192 VSUBS 0.068066f
C233 B.n193 VSUBS 0.019329f
C234 B.n194 VSUBS 0.007852f
C235 B.n195 VSUBS 0.008342f
C236 B.n196 VSUBS 0.008342f
C237 B.n197 VSUBS 0.008342f
C238 B.n198 VSUBS 0.008342f
C239 B.n199 VSUBS 0.008342f
C240 B.n200 VSUBS 0.008342f
C241 B.n201 VSUBS 0.008342f
C242 B.n202 VSUBS 0.008342f
C243 B.n203 VSUBS 0.008342f
C244 B.n204 VSUBS 0.008342f
C245 B.n205 VSUBS 0.008342f
C246 B.n206 VSUBS 0.008342f
C247 B.n207 VSUBS 0.008342f
C248 B.n208 VSUBS 0.008342f
C249 B.n209 VSUBS 0.008342f
C250 B.n210 VSUBS 0.004662f
C251 B.n211 VSUBS 0.019329f
C252 B.n212 VSUBS 0.007852f
C253 B.n213 VSUBS 0.008342f
C254 B.n214 VSUBS 0.008342f
C255 B.n215 VSUBS 0.008342f
C256 B.n216 VSUBS 0.008342f
C257 B.n217 VSUBS 0.008342f
C258 B.n218 VSUBS 0.008342f
C259 B.n219 VSUBS 0.008342f
C260 B.n220 VSUBS 0.008342f
C261 B.n221 VSUBS 0.008342f
C262 B.n222 VSUBS 0.008342f
C263 B.n223 VSUBS 0.008342f
C264 B.n224 VSUBS 0.008342f
C265 B.n225 VSUBS 0.008342f
C266 B.n226 VSUBS 0.008342f
C267 B.n227 VSUBS 0.008342f
C268 B.n228 VSUBS 0.008342f
C269 B.n229 VSUBS 0.008342f
C270 B.n230 VSUBS 0.019254f
C271 B.n231 VSUBS 0.019759f
C272 B.n232 VSUBS 0.018773f
C273 B.n233 VSUBS 0.008342f
C274 B.n234 VSUBS 0.008342f
C275 B.n235 VSUBS 0.008342f
C276 B.n236 VSUBS 0.008342f
C277 B.n237 VSUBS 0.008342f
C278 B.n238 VSUBS 0.008342f
C279 B.n239 VSUBS 0.008342f
C280 B.n240 VSUBS 0.008342f
C281 B.n241 VSUBS 0.008342f
C282 B.n242 VSUBS 0.008342f
C283 B.n243 VSUBS 0.008342f
C284 B.n244 VSUBS 0.008342f
C285 B.n245 VSUBS 0.008342f
C286 B.n246 VSUBS 0.008342f
C287 B.n247 VSUBS 0.008342f
C288 B.n248 VSUBS 0.008342f
C289 B.n249 VSUBS 0.008342f
C290 B.n250 VSUBS 0.008342f
C291 B.n251 VSUBS 0.008342f
C292 B.n252 VSUBS 0.008342f
C293 B.n253 VSUBS 0.008342f
C294 B.n254 VSUBS 0.008342f
C295 B.n255 VSUBS 0.008342f
C296 B.n256 VSUBS 0.008342f
C297 B.n257 VSUBS 0.008342f
C298 B.n258 VSUBS 0.008342f
C299 B.n259 VSUBS 0.008342f
C300 B.n260 VSUBS 0.008342f
C301 B.n261 VSUBS 0.008342f
C302 B.n262 VSUBS 0.008342f
C303 B.n263 VSUBS 0.008342f
C304 B.n264 VSUBS 0.008342f
C305 B.n265 VSUBS 0.008342f
C306 B.n266 VSUBS 0.008342f
C307 B.n267 VSUBS 0.008342f
C308 B.n268 VSUBS 0.008342f
C309 B.n269 VSUBS 0.008342f
C310 B.n270 VSUBS 0.008342f
C311 B.n271 VSUBS 0.008342f
C312 B.n272 VSUBS 0.008342f
C313 B.n273 VSUBS 0.008342f
C314 B.n274 VSUBS 0.008342f
C315 B.n275 VSUBS 0.008342f
C316 B.n276 VSUBS 0.008342f
C317 B.n277 VSUBS 0.008342f
C318 B.n278 VSUBS 0.008342f
C319 B.n279 VSUBS 0.008342f
C320 B.n280 VSUBS 0.008342f
C321 B.n281 VSUBS 0.008342f
C322 B.n282 VSUBS 0.008342f
C323 B.n283 VSUBS 0.008342f
C324 B.n284 VSUBS 0.008342f
C325 B.n285 VSUBS 0.008342f
C326 B.n286 VSUBS 0.008342f
C327 B.n287 VSUBS 0.008342f
C328 B.n288 VSUBS 0.008342f
C329 B.n289 VSUBS 0.008342f
C330 B.n290 VSUBS 0.008342f
C331 B.n291 VSUBS 0.008342f
C332 B.n292 VSUBS 0.008342f
C333 B.n293 VSUBS 0.008342f
C334 B.n294 VSUBS 0.008342f
C335 B.n295 VSUBS 0.008342f
C336 B.n296 VSUBS 0.008342f
C337 B.n297 VSUBS 0.008342f
C338 B.n298 VSUBS 0.008342f
C339 B.n299 VSUBS 0.008342f
C340 B.n300 VSUBS 0.008342f
C341 B.n301 VSUBS 0.008342f
C342 B.n302 VSUBS 0.008342f
C343 B.n303 VSUBS 0.008342f
C344 B.n304 VSUBS 0.008342f
C345 B.n305 VSUBS 0.008342f
C346 B.n306 VSUBS 0.008342f
C347 B.n307 VSUBS 0.008342f
C348 B.n308 VSUBS 0.008342f
C349 B.n309 VSUBS 0.008342f
C350 B.n310 VSUBS 0.008342f
C351 B.n311 VSUBS 0.008342f
C352 B.n312 VSUBS 0.008342f
C353 B.n313 VSUBS 0.008342f
C354 B.n314 VSUBS 0.008342f
C355 B.n315 VSUBS 0.008342f
C356 B.n316 VSUBS 0.008342f
C357 B.n317 VSUBS 0.008342f
C358 B.n318 VSUBS 0.008342f
C359 B.n319 VSUBS 0.008342f
C360 B.n320 VSUBS 0.008342f
C361 B.n321 VSUBS 0.008342f
C362 B.n322 VSUBS 0.008342f
C363 B.n323 VSUBS 0.008342f
C364 B.n324 VSUBS 0.008342f
C365 B.n325 VSUBS 0.008342f
C366 B.n326 VSUBS 0.008342f
C367 B.n327 VSUBS 0.008342f
C368 B.n328 VSUBS 0.008342f
C369 B.n329 VSUBS 0.008342f
C370 B.n330 VSUBS 0.008342f
C371 B.n331 VSUBS 0.008342f
C372 B.n332 VSUBS 0.008342f
C373 B.n333 VSUBS 0.008342f
C374 B.n334 VSUBS 0.008342f
C375 B.n335 VSUBS 0.008342f
C376 B.n336 VSUBS 0.008342f
C377 B.n337 VSUBS 0.008342f
C378 B.n338 VSUBS 0.008342f
C379 B.n339 VSUBS 0.008342f
C380 B.n340 VSUBS 0.008342f
C381 B.n341 VSUBS 0.008342f
C382 B.n342 VSUBS 0.008342f
C383 B.n343 VSUBS 0.008342f
C384 B.n344 VSUBS 0.018773f
C385 B.n345 VSUBS 0.020241f
C386 B.n346 VSUBS 0.020241f
C387 B.n347 VSUBS 0.008342f
C388 B.n348 VSUBS 0.008342f
C389 B.n349 VSUBS 0.008342f
C390 B.n350 VSUBS 0.008342f
C391 B.n351 VSUBS 0.008342f
C392 B.n352 VSUBS 0.008342f
C393 B.n353 VSUBS 0.008342f
C394 B.n354 VSUBS 0.008342f
C395 B.n355 VSUBS 0.008342f
C396 B.n356 VSUBS 0.008342f
C397 B.n357 VSUBS 0.008342f
C398 B.n358 VSUBS 0.008342f
C399 B.n359 VSUBS 0.008342f
C400 B.n360 VSUBS 0.008342f
C401 B.n361 VSUBS 0.008342f
C402 B.n362 VSUBS 0.008342f
C403 B.n363 VSUBS 0.007852f
C404 B.n364 VSUBS 0.008342f
C405 B.n365 VSUBS 0.008342f
C406 B.n366 VSUBS 0.004662f
C407 B.n367 VSUBS 0.008342f
C408 B.n368 VSUBS 0.008342f
C409 B.n369 VSUBS 0.008342f
C410 B.n370 VSUBS 0.008342f
C411 B.n371 VSUBS 0.008342f
C412 B.n372 VSUBS 0.008342f
C413 B.n373 VSUBS 0.008342f
C414 B.n374 VSUBS 0.008342f
C415 B.n375 VSUBS 0.008342f
C416 B.n376 VSUBS 0.008342f
C417 B.n377 VSUBS 0.008342f
C418 B.n378 VSUBS 0.008342f
C419 B.n379 VSUBS 0.004662f
C420 B.n380 VSUBS 0.019329f
C421 B.n381 VSUBS 0.007852f
C422 B.n382 VSUBS 0.008342f
C423 B.n383 VSUBS 0.008342f
C424 B.n384 VSUBS 0.008342f
C425 B.n385 VSUBS 0.008342f
C426 B.n386 VSUBS 0.008342f
C427 B.n387 VSUBS 0.008342f
C428 B.n388 VSUBS 0.008342f
C429 B.n389 VSUBS 0.008342f
C430 B.n390 VSUBS 0.008342f
C431 B.n391 VSUBS 0.008342f
C432 B.n392 VSUBS 0.008342f
C433 B.n393 VSUBS 0.008342f
C434 B.n394 VSUBS 0.008342f
C435 B.n395 VSUBS 0.008342f
C436 B.n396 VSUBS 0.008342f
C437 B.n397 VSUBS 0.008342f
C438 B.n398 VSUBS 0.008342f
C439 B.n399 VSUBS 0.020241f
C440 B.n400 VSUBS 0.020241f
C441 B.n401 VSUBS 0.018773f
C442 B.n402 VSUBS 0.008342f
C443 B.n403 VSUBS 0.008342f
C444 B.n404 VSUBS 0.008342f
C445 B.n405 VSUBS 0.008342f
C446 B.n406 VSUBS 0.008342f
C447 B.n407 VSUBS 0.008342f
C448 B.n408 VSUBS 0.008342f
C449 B.n409 VSUBS 0.008342f
C450 B.n410 VSUBS 0.008342f
C451 B.n411 VSUBS 0.008342f
C452 B.n412 VSUBS 0.008342f
C453 B.n413 VSUBS 0.008342f
C454 B.n414 VSUBS 0.008342f
C455 B.n415 VSUBS 0.008342f
C456 B.n416 VSUBS 0.008342f
C457 B.n417 VSUBS 0.008342f
C458 B.n418 VSUBS 0.008342f
C459 B.n419 VSUBS 0.008342f
C460 B.n420 VSUBS 0.008342f
C461 B.n421 VSUBS 0.008342f
C462 B.n422 VSUBS 0.008342f
C463 B.n423 VSUBS 0.008342f
C464 B.n424 VSUBS 0.008342f
C465 B.n425 VSUBS 0.008342f
C466 B.n426 VSUBS 0.008342f
C467 B.n427 VSUBS 0.008342f
C468 B.n428 VSUBS 0.008342f
C469 B.n429 VSUBS 0.008342f
C470 B.n430 VSUBS 0.008342f
C471 B.n431 VSUBS 0.008342f
C472 B.n432 VSUBS 0.008342f
C473 B.n433 VSUBS 0.008342f
C474 B.n434 VSUBS 0.008342f
C475 B.n435 VSUBS 0.008342f
C476 B.n436 VSUBS 0.008342f
C477 B.n437 VSUBS 0.008342f
C478 B.n438 VSUBS 0.008342f
C479 B.n439 VSUBS 0.008342f
C480 B.n440 VSUBS 0.008342f
C481 B.n441 VSUBS 0.008342f
C482 B.n442 VSUBS 0.008342f
C483 B.n443 VSUBS 0.008342f
C484 B.n444 VSUBS 0.008342f
C485 B.n445 VSUBS 0.008342f
C486 B.n446 VSUBS 0.008342f
C487 B.n447 VSUBS 0.008342f
C488 B.n448 VSUBS 0.008342f
C489 B.n449 VSUBS 0.008342f
C490 B.n450 VSUBS 0.008342f
C491 B.n451 VSUBS 0.008342f
C492 B.n452 VSUBS 0.008342f
C493 B.n453 VSUBS 0.008342f
C494 B.n454 VSUBS 0.008342f
C495 B.n455 VSUBS 0.010886f
C496 B.n456 VSUBS 0.011597f
C497 B.n457 VSUBS 0.023062f
C498 VDD1.t4 VSUBS 0.045212f
C499 VDD1.t3 VSUBS 0.045212f
C500 VDD1.n0 VSUBS 0.204921f
C501 VDD1.t5 VSUBS 0.045212f
C502 VDD1.t0 VSUBS 0.045212f
C503 VDD1.n1 VSUBS 0.20454f
C504 VDD1.t6 VSUBS 0.045212f
C505 VDD1.t1 VSUBS 0.045212f
C506 VDD1.n2 VSUBS 0.20454f
C507 VDD1.n3 VSUBS 2.38992f
C508 VDD1.t2 VSUBS 0.045212f
C509 VDD1.t7 VSUBS 0.045212f
C510 VDD1.n4 VSUBS 0.202138f
C511 VDD1.n5 VSUBS 1.97992f
C512 VP.n0 VSUBS 0.059496f
C513 VP.t6 VSUBS 0.548093f
C514 VP.n1 VSUBS 0.048173f
C515 VP.n2 VSUBS 0.059496f
C516 VP.t1 VSUBS 0.548093f
C517 VP.n3 VSUBS 0.048097f
C518 VP.n4 VSUBS 0.059496f
C519 VP.t7 VSUBS 0.548093f
C520 VP.n5 VSUBS 0.048173f
C521 VP.n6 VSUBS 0.059496f
C522 VP.t2 VSUBS 0.548093f
C523 VP.n7 VSUBS 0.059496f
C524 VP.t0 VSUBS 0.548093f
C525 VP.n8 VSUBS 0.048173f
C526 VP.n9 VSUBS 0.059496f
C527 VP.t5 VSUBS 0.548093f
C528 VP.n10 VSUBS 0.048097f
C529 VP.n11 VSUBS 0.375705f
C530 VP.t4 VSUBS 0.548093f
C531 VP.t3 VSUBS 0.783175f
C532 VP.n12 VSUBS 0.396345f
C533 VP.n13 VSUBS 0.368723f
C534 VP.n14 VSUBS 0.056685f
C535 VP.n15 VSUBS 0.118248f
C536 VP.n16 VSUBS 0.059496f
C537 VP.n17 VSUBS 0.059496f
C538 VP.n18 VSUBS 0.059496f
C539 VP.n19 VSUBS 0.118248f
C540 VP.n20 VSUBS 0.056685f
C541 VP.n21 VSUBS 0.268561f
C542 VP.n22 VSUBS 0.118255f
C543 VP.n23 VSUBS 0.059496f
C544 VP.n24 VSUBS 0.059496f
C545 VP.n25 VSUBS 0.059496f
C546 VP.n26 VSUBS 0.117613f
C547 VP.n27 VSUBS 0.05778f
C548 VP.n28 VSUBS 0.383833f
C549 VP.n29 VSUBS 2.18625f
C550 VP.n30 VSUBS 2.241f
C551 VP.n31 VSUBS 0.383833f
C552 VP.n32 VSUBS 0.05778f
C553 VP.n33 VSUBS 0.117613f
C554 VP.n34 VSUBS 0.059496f
C555 VP.n35 VSUBS 0.059496f
C556 VP.n36 VSUBS 0.059496f
C557 VP.n37 VSUBS 0.118255f
C558 VP.n38 VSUBS 0.268561f
C559 VP.n39 VSUBS 0.056685f
C560 VP.n40 VSUBS 0.118248f
C561 VP.n41 VSUBS 0.059496f
C562 VP.n42 VSUBS 0.059496f
C563 VP.n43 VSUBS 0.059496f
C564 VP.n44 VSUBS 0.118248f
C565 VP.n45 VSUBS 0.056685f
C566 VP.n46 VSUBS 0.268561f
C567 VP.n47 VSUBS 0.118255f
C568 VP.n48 VSUBS 0.059496f
C569 VP.n49 VSUBS 0.059496f
C570 VP.n50 VSUBS 0.059496f
C571 VP.n51 VSUBS 0.117613f
C572 VP.n52 VSUBS 0.05778f
C573 VP.n53 VSUBS 0.383833f
C574 VP.n54 VSUBS 0.063068f
C575 VTAIL.t12 VSUBS 0.050575f
C576 VTAIL.t14 VSUBS 0.050575f
C577 VTAIL.n0 VSUBS 0.191292f
C578 VTAIL.n1 VSUBS 0.484342f
C579 VTAIL.t8 VSUBS 0.305666f
C580 VTAIL.n2 VSUBS 0.544969f
C581 VTAIL.t1 VSUBS 0.305666f
C582 VTAIL.n3 VSUBS 0.544969f
C583 VTAIL.t0 VSUBS 0.050575f
C584 VTAIL.t6 VSUBS 0.050575f
C585 VTAIL.n4 VSUBS 0.191292f
C586 VTAIL.n5 VSUBS 0.635143f
C587 VTAIL.t5 VSUBS 0.305666f
C588 VTAIL.n6 VSUBS 1.21611f
C589 VTAIL.t15 VSUBS 0.305667f
C590 VTAIL.n7 VSUBS 1.21611f
C591 VTAIL.t10 VSUBS 0.050575f
C592 VTAIL.t11 VSUBS 0.050575f
C593 VTAIL.n8 VSUBS 0.191293f
C594 VTAIL.n9 VSUBS 0.635142f
C595 VTAIL.t13 VSUBS 0.305667f
C596 VTAIL.n10 VSUBS 0.544968f
C597 VTAIL.t4 VSUBS 0.305667f
C598 VTAIL.n11 VSUBS 0.544968f
C599 VTAIL.t3 VSUBS 0.050575f
C600 VTAIL.t2 VSUBS 0.050575f
C601 VTAIL.n12 VSUBS 0.191293f
C602 VTAIL.n13 VSUBS 0.635142f
C603 VTAIL.t7 VSUBS 0.305667f
C604 VTAIL.n14 VSUBS 1.21611f
C605 VTAIL.t9 VSUBS 0.305666f
C606 VTAIL.n15 VSUBS 1.21087f
C607 VDD2.t3 VSUBS 0.03035f
C608 VDD2.t6 VSUBS 0.03035f
C609 VDD2.n0 VSUBS 0.137304f
C610 VDD2.t0 VSUBS 0.03035f
C611 VDD2.t7 VSUBS 0.03035f
C612 VDD2.n1 VSUBS 0.137304f
C613 VDD2.n2 VSUBS 1.56885f
C614 VDD2.t4 VSUBS 0.03035f
C615 VDD2.t1 VSUBS 0.03035f
C616 VDD2.n3 VSUBS 0.135691f
C617 VDD2.n4 VSUBS 1.30889f
C618 VDD2.t2 VSUBS 0.03035f
C619 VDD2.t5 VSUBS 0.03035f
C620 VDD2.n5 VSUBS 0.137296f
C621 VN.n0 VSUBS 0.049504f
C622 VN.t6 VSUBS 0.456042f
C623 VN.n1 VSUBS 0.040083f
C624 VN.n2 VSUBS 0.049504f
C625 VN.t1 VSUBS 0.456042f
C626 VN.n3 VSUBS 0.040019f
C627 VN.n4 VSUBS 0.312607f
C628 VN.t3 VSUBS 0.456042f
C629 VN.t7 VSUBS 0.651643f
C630 VN.n5 VSUBS 0.32978f
C631 VN.n6 VSUBS 0.306797f
C632 VN.n7 VSUBS 0.047165f
C633 VN.n8 VSUBS 0.098388f
C634 VN.n9 VSUBS 0.049504f
C635 VN.n10 VSUBS 0.049504f
C636 VN.n11 VSUBS 0.049504f
C637 VN.n12 VSUBS 0.098388f
C638 VN.n13 VSUBS 0.047165f
C639 VN.n14 VSUBS 0.223457f
C640 VN.n15 VSUBS 0.098395f
C641 VN.n16 VSUBS 0.049504f
C642 VN.n17 VSUBS 0.049504f
C643 VN.n18 VSUBS 0.049504f
C644 VN.n19 VSUBS 0.09786f
C645 VN.n20 VSUBS 0.048076f
C646 VN.n21 VSUBS 0.31937f
C647 VN.n22 VSUBS 0.052476f
C648 VN.n23 VSUBS 0.049504f
C649 VN.t0 VSUBS 0.456042f
C650 VN.n24 VSUBS 0.040083f
C651 VN.n25 VSUBS 0.049504f
C652 VN.t5 VSUBS 0.456042f
C653 VN.n26 VSUBS 0.040019f
C654 VN.n27 VSUBS 0.312607f
C655 VN.t4 VSUBS 0.456042f
C656 VN.t2 VSUBS 0.651643f
C657 VN.n28 VSUBS 0.32978f
C658 VN.n29 VSUBS 0.306797f
C659 VN.n30 VSUBS 0.047165f
C660 VN.n31 VSUBS 0.098388f
C661 VN.n32 VSUBS 0.049504f
C662 VN.n33 VSUBS 0.049504f
C663 VN.n34 VSUBS 0.049504f
C664 VN.n35 VSUBS 0.098388f
C665 VN.n36 VSUBS 0.047165f
C666 VN.n37 VSUBS 0.223457f
C667 VN.n38 VSUBS 0.098395f
C668 VN.n39 VSUBS 0.049504f
C669 VN.n40 VSUBS 0.049504f
C670 VN.n41 VSUBS 0.049504f
C671 VN.n42 VSUBS 0.09786f
C672 VN.n43 VSUBS 0.048076f
C673 VN.n44 VSUBS 0.31937f
C674 VN.n45 VSUBS 1.85173f
.ends

