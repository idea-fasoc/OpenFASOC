* NGSPICE file created from diff_pair_sample_0734.ext - technology: sky130A

.subckt diff_pair_sample_0734 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=2.87
X1 B.t11 B.t9 B.t10 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=2.87
X2 VTAIL.t4 VN.t0 VDD2.t7 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X3 B.t8 B.t6 B.t7 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=2.87
X4 B.t5 B.t3 B.t4 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=2.87
X5 VTAIL.t5 VN.t1 VDD2.t6 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=2.87
X6 VTAIL.t7 VN.t2 VDD2.t5 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=2.87
X7 VDD1.t1 VP.t1 VTAIL.t14 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X8 VDD2.t4 VN.t3 VTAIL.t6 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X9 VTAIL.t13 VP.t2 VDD1.t2 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X10 VTAIL.t12 VP.t3 VDD1.t3 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0.627 ps=4.13 w=3.8 l=2.87
X11 VTAIL.t11 VP.t4 VDD1.t0 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X12 VDD2.t3 VN.t4 VTAIL.t3 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=2.87
X13 VDD1.t4 VP.t5 VTAIL.t10 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=2.87
X14 VDD2.t2 VN.t5 VTAIL.t1 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X15 VTAIL.t2 VN.t6 VDD2.t1 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X16 VDD2.t0 VN.t7 VTAIL.t0 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=2.87
X17 VDD1.t5 VP.t6 VTAIL.t9 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=1.482 ps=8.38 w=3.8 l=2.87
X18 VDD1.t6 VP.t7 VTAIL.t8 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=0.627 pd=4.13 as=0.627 ps=4.13 w=3.8 l=2.87
X19 B.t2 B.t0 B.t1 w_n4170_n1728# sky130_fd_pr__pfet_01v8 ad=1.482 pd=8.38 as=0 ps=0 w=3.8 l=2.87
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n28 VP.n27 161.3
R6 VP.n29 VP.n13 161.3
R7 VP.n31 VP.n30 161.3
R8 VP.n32 VP.n12 161.3
R9 VP.n34 VP.n33 161.3
R10 VP.n35 VP.n11 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n38 VP.n10 161.3
R13 VP.n74 VP.n0 161.3
R14 VP.n73 VP.n72 161.3
R15 VP.n71 VP.n1 161.3
R16 VP.n70 VP.n69 161.3
R17 VP.n68 VP.n2 161.3
R18 VP.n67 VP.n66 161.3
R19 VP.n65 VP.n3 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n53 VP.n52 161.3
R27 VP.n51 VP.n7 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n8 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n45 VP.n9 161.3
R32 VP.n44 VP.n43 161.3
R33 VP.n42 VP.n41 108.45
R34 VP.n76 VP.n75 108.45
R35 VP.n40 VP.n39 108.45
R36 VP.n17 VP.t0 64.9524
R37 VP.n18 VP.n17 56.7106
R38 VP.n60 VP.n5 56.5617
R39 VP.n24 VP.n15 56.5617
R40 VP.n41 VP.n40 45.9163
R41 VP.n49 VP.n48 45.4209
R42 VP.n69 VP.n68 45.4209
R43 VP.n33 VP.n32 45.4209
R44 VP.n48 VP.n47 35.7332
R45 VP.n69 VP.n1 35.7332
R46 VP.n33 VP.n11 35.7332
R47 VP.n42 VP.t3 31.9099
R48 VP.n54 VP.t7 31.9099
R49 VP.n62 VP.t2 31.9099
R50 VP.n75 VP.t6 31.9099
R51 VP.n39 VP.t5 31.9099
R52 VP.n26 VP.t4 31.9099
R53 VP.n18 VP.t1 31.9099
R54 VP.n43 VP.n9 24.5923
R55 VP.n47 VP.n9 24.5923
R56 VP.n49 VP.n7 24.5923
R57 VP.n53 VP.n7 24.5923
R58 VP.n56 VP.n55 24.5923
R59 VP.n56 VP.n5 24.5923
R60 VP.n61 VP.n60 24.5923
R61 VP.n63 VP.n61 24.5923
R62 VP.n67 VP.n3 24.5923
R63 VP.n68 VP.n67 24.5923
R64 VP.n73 VP.n1 24.5923
R65 VP.n74 VP.n73 24.5923
R66 VP.n37 VP.n11 24.5923
R67 VP.n38 VP.n37 24.5923
R68 VP.n25 VP.n24 24.5923
R69 VP.n27 VP.n25 24.5923
R70 VP.n31 VP.n13 24.5923
R71 VP.n32 VP.n31 24.5923
R72 VP.n20 VP.n19 24.5923
R73 VP.n20 VP.n15 24.5923
R74 VP.n55 VP.n54 17.2148
R75 VP.n63 VP.n62 17.2148
R76 VP.n27 VP.n26 17.2148
R77 VP.n19 VP.n18 17.2148
R78 VP.n54 VP.n53 7.37805
R79 VP.n62 VP.n3 7.37805
R80 VP.n26 VP.n13 7.37805
R81 VP.n17 VP.n16 5.07592
R82 VP.n43 VP.n42 2.45968
R83 VP.n75 VP.n74 2.45968
R84 VP.n39 VP.n38 2.45968
R85 VP.n40 VP.n10 0.278335
R86 VP.n44 VP.n41 0.278335
R87 VP.n76 VP.n0 0.278335
R88 VP.n21 VP.n16 0.189894
R89 VP.n22 VP.n21 0.189894
R90 VP.n23 VP.n22 0.189894
R91 VP.n23 VP.n14 0.189894
R92 VP.n28 VP.n14 0.189894
R93 VP.n29 VP.n28 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n12 0.189894
R96 VP.n34 VP.n12 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n10 0.189894
R100 VP.n45 VP.n44 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n46 VP.n8 0.189894
R103 VP.n50 VP.n8 0.189894
R104 VP.n51 VP.n50 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n52 VP.n6 0.189894
R107 VP.n57 VP.n6 0.189894
R108 VP.n58 VP.n57 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n59 VP.n4 0.189894
R111 VP.n64 VP.n4 0.189894
R112 VP.n65 VP.n64 0.189894
R113 VP.n66 VP.n65 0.189894
R114 VP.n66 VP.n2 0.189894
R115 VP.n70 VP.n2 0.189894
R116 VP.n71 VP.n70 0.189894
R117 VP.n72 VP.n71 0.189894
R118 VP.n72 VP.n0 0.189894
R119 VP VP.n76 0.153485
R120 VDD1 VDD1.n0 114.231
R121 VDD1.n3 VDD1.n2 114.117
R122 VDD1.n3 VDD1.n1 114.117
R123 VDD1.n5 VDD1.n4 112.793
R124 VDD1.n5 VDD1.n3 39.988
R125 VDD1.n4 VDD1.t0 8.55445
R126 VDD1.n4 VDD1.t4 8.55445
R127 VDD1.n0 VDD1.t7 8.55445
R128 VDD1.n0 VDD1.t1 8.55445
R129 VDD1.n2 VDD1.t2 8.55445
R130 VDD1.n2 VDD1.t5 8.55445
R131 VDD1.n1 VDD1.t3 8.55445
R132 VDD1.n1 VDD1.t6 8.55445
R133 VDD1 VDD1.n5 1.32162
R134 VTAIL.n162 VTAIL.n148 756.745
R135 VTAIL.n16 VTAIL.n2 756.745
R136 VTAIL.n36 VTAIL.n22 756.745
R137 VTAIL.n58 VTAIL.n44 756.745
R138 VTAIL.n142 VTAIL.n128 756.745
R139 VTAIL.n120 VTAIL.n106 756.745
R140 VTAIL.n100 VTAIL.n86 756.745
R141 VTAIL.n78 VTAIL.n64 756.745
R142 VTAIL.n155 VTAIL.n154 585
R143 VTAIL.n152 VTAIL.n151 585
R144 VTAIL.n161 VTAIL.n160 585
R145 VTAIL.n163 VTAIL.n162 585
R146 VTAIL.n9 VTAIL.n8 585
R147 VTAIL.n6 VTAIL.n5 585
R148 VTAIL.n15 VTAIL.n14 585
R149 VTAIL.n17 VTAIL.n16 585
R150 VTAIL.n29 VTAIL.n28 585
R151 VTAIL.n26 VTAIL.n25 585
R152 VTAIL.n35 VTAIL.n34 585
R153 VTAIL.n37 VTAIL.n36 585
R154 VTAIL.n51 VTAIL.n50 585
R155 VTAIL.n48 VTAIL.n47 585
R156 VTAIL.n57 VTAIL.n56 585
R157 VTAIL.n59 VTAIL.n58 585
R158 VTAIL.n143 VTAIL.n142 585
R159 VTAIL.n141 VTAIL.n140 585
R160 VTAIL.n132 VTAIL.n131 585
R161 VTAIL.n135 VTAIL.n134 585
R162 VTAIL.n121 VTAIL.n120 585
R163 VTAIL.n119 VTAIL.n118 585
R164 VTAIL.n110 VTAIL.n109 585
R165 VTAIL.n113 VTAIL.n112 585
R166 VTAIL.n101 VTAIL.n100 585
R167 VTAIL.n99 VTAIL.n98 585
R168 VTAIL.n90 VTAIL.n89 585
R169 VTAIL.n93 VTAIL.n92 585
R170 VTAIL.n79 VTAIL.n78 585
R171 VTAIL.n77 VTAIL.n76 585
R172 VTAIL.n68 VTAIL.n67 585
R173 VTAIL.n71 VTAIL.n70 585
R174 VTAIL.t0 VTAIL.n153 330.707
R175 VTAIL.t7 VTAIL.n7 330.707
R176 VTAIL.t9 VTAIL.n27 330.707
R177 VTAIL.t12 VTAIL.n49 330.707
R178 VTAIL.t10 VTAIL.n133 330.707
R179 VTAIL.t15 VTAIL.n111 330.707
R180 VTAIL.t3 VTAIL.n91 330.707
R181 VTAIL.t5 VTAIL.n69 330.707
R182 VTAIL.n154 VTAIL.n151 171.744
R183 VTAIL.n161 VTAIL.n151 171.744
R184 VTAIL.n162 VTAIL.n161 171.744
R185 VTAIL.n8 VTAIL.n5 171.744
R186 VTAIL.n15 VTAIL.n5 171.744
R187 VTAIL.n16 VTAIL.n15 171.744
R188 VTAIL.n28 VTAIL.n25 171.744
R189 VTAIL.n35 VTAIL.n25 171.744
R190 VTAIL.n36 VTAIL.n35 171.744
R191 VTAIL.n50 VTAIL.n47 171.744
R192 VTAIL.n57 VTAIL.n47 171.744
R193 VTAIL.n58 VTAIL.n57 171.744
R194 VTAIL.n142 VTAIL.n141 171.744
R195 VTAIL.n141 VTAIL.n131 171.744
R196 VTAIL.n134 VTAIL.n131 171.744
R197 VTAIL.n120 VTAIL.n119 171.744
R198 VTAIL.n119 VTAIL.n109 171.744
R199 VTAIL.n112 VTAIL.n109 171.744
R200 VTAIL.n100 VTAIL.n99 171.744
R201 VTAIL.n99 VTAIL.n89 171.744
R202 VTAIL.n92 VTAIL.n89 171.744
R203 VTAIL.n78 VTAIL.n77 171.744
R204 VTAIL.n77 VTAIL.n67 171.744
R205 VTAIL.n70 VTAIL.n67 171.744
R206 VTAIL.n127 VTAIL.n126 96.1138
R207 VTAIL.n85 VTAIL.n84 96.1138
R208 VTAIL.n1 VTAIL.n0 96.1136
R209 VTAIL.n43 VTAIL.n42 96.1136
R210 VTAIL.n154 VTAIL.t0 85.8723
R211 VTAIL.n8 VTAIL.t7 85.8723
R212 VTAIL.n28 VTAIL.t9 85.8723
R213 VTAIL.n50 VTAIL.t12 85.8723
R214 VTAIL.n134 VTAIL.t10 85.8723
R215 VTAIL.n112 VTAIL.t15 85.8723
R216 VTAIL.n92 VTAIL.t3 85.8723
R217 VTAIL.n70 VTAIL.t5 85.8723
R218 VTAIL.n167 VTAIL.n166 31.4096
R219 VTAIL.n21 VTAIL.n20 31.4096
R220 VTAIL.n41 VTAIL.n40 31.4096
R221 VTAIL.n63 VTAIL.n62 31.4096
R222 VTAIL.n147 VTAIL.n146 31.4096
R223 VTAIL.n125 VTAIL.n124 31.4096
R224 VTAIL.n105 VTAIL.n104 31.4096
R225 VTAIL.n83 VTAIL.n82 31.4096
R226 VTAIL.n167 VTAIL.n147 18.4014
R227 VTAIL.n83 VTAIL.n63 18.4014
R228 VTAIL.n155 VTAIL.n153 16.3201
R229 VTAIL.n9 VTAIL.n7 16.3201
R230 VTAIL.n29 VTAIL.n27 16.3201
R231 VTAIL.n51 VTAIL.n49 16.3201
R232 VTAIL.n135 VTAIL.n133 16.3201
R233 VTAIL.n113 VTAIL.n111 16.3201
R234 VTAIL.n93 VTAIL.n91 16.3201
R235 VTAIL.n71 VTAIL.n69 16.3201
R236 VTAIL.n156 VTAIL.n152 12.8005
R237 VTAIL.n10 VTAIL.n6 12.8005
R238 VTAIL.n30 VTAIL.n26 12.8005
R239 VTAIL.n52 VTAIL.n48 12.8005
R240 VTAIL.n136 VTAIL.n132 12.8005
R241 VTAIL.n114 VTAIL.n110 12.8005
R242 VTAIL.n94 VTAIL.n90 12.8005
R243 VTAIL.n72 VTAIL.n68 12.8005
R244 VTAIL.n160 VTAIL.n159 12.0247
R245 VTAIL.n14 VTAIL.n13 12.0247
R246 VTAIL.n34 VTAIL.n33 12.0247
R247 VTAIL.n56 VTAIL.n55 12.0247
R248 VTAIL.n140 VTAIL.n139 12.0247
R249 VTAIL.n118 VTAIL.n117 12.0247
R250 VTAIL.n98 VTAIL.n97 12.0247
R251 VTAIL.n76 VTAIL.n75 12.0247
R252 VTAIL.n163 VTAIL.n150 11.249
R253 VTAIL.n17 VTAIL.n4 11.249
R254 VTAIL.n37 VTAIL.n24 11.249
R255 VTAIL.n59 VTAIL.n46 11.249
R256 VTAIL.n143 VTAIL.n130 11.249
R257 VTAIL.n121 VTAIL.n108 11.249
R258 VTAIL.n101 VTAIL.n88 11.249
R259 VTAIL.n79 VTAIL.n66 11.249
R260 VTAIL.n164 VTAIL.n148 10.4732
R261 VTAIL.n18 VTAIL.n2 10.4732
R262 VTAIL.n38 VTAIL.n22 10.4732
R263 VTAIL.n60 VTAIL.n44 10.4732
R264 VTAIL.n144 VTAIL.n128 10.4732
R265 VTAIL.n122 VTAIL.n106 10.4732
R266 VTAIL.n102 VTAIL.n86 10.4732
R267 VTAIL.n80 VTAIL.n64 10.4732
R268 VTAIL.n166 VTAIL.n165 9.45567
R269 VTAIL.n20 VTAIL.n19 9.45567
R270 VTAIL.n40 VTAIL.n39 9.45567
R271 VTAIL.n62 VTAIL.n61 9.45567
R272 VTAIL.n146 VTAIL.n145 9.45567
R273 VTAIL.n124 VTAIL.n123 9.45567
R274 VTAIL.n104 VTAIL.n103 9.45567
R275 VTAIL.n82 VTAIL.n81 9.45567
R276 VTAIL.n165 VTAIL.n164 9.3005
R277 VTAIL.n150 VTAIL.n149 9.3005
R278 VTAIL.n159 VTAIL.n158 9.3005
R279 VTAIL.n157 VTAIL.n156 9.3005
R280 VTAIL.n19 VTAIL.n18 9.3005
R281 VTAIL.n4 VTAIL.n3 9.3005
R282 VTAIL.n13 VTAIL.n12 9.3005
R283 VTAIL.n11 VTAIL.n10 9.3005
R284 VTAIL.n39 VTAIL.n38 9.3005
R285 VTAIL.n24 VTAIL.n23 9.3005
R286 VTAIL.n33 VTAIL.n32 9.3005
R287 VTAIL.n31 VTAIL.n30 9.3005
R288 VTAIL.n61 VTAIL.n60 9.3005
R289 VTAIL.n46 VTAIL.n45 9.3005
R290 VTAIL.n55 VTAIL.n54 9.3005
R291 VTAIL.n53 VTAIL.n52 9.3005
R292 VTAIL.n145 VTAIL.n144 9.3005
R293 VTAIL.n130 VTAIL.n129 9.3005
R294 VTAIL.n139 VTAIL.n138 9.3005
R295 VTAIL.n137 VTAIL.n136 9.3005
R296 VTAIL.n123 VTAIL.n122 9.3005
R297 VTAIL.n108 VTAIL.n107 9.3005
R298 VTAIL.n117 VTAIL.n116 9.3005
R299 VTAIL.n115 VTAIL.n114 9.3005
R300 VTAIL.n103 VTAIL.n102 9.3005
R301 VTAIL.n88 VTAIL.n87 9.3005
R302 VTAIL.n97 VTAIL.n96 9.3005
R303 VTAIL.n95 VTAIL.n94 9.3005
R304 VTAIL.n81 VTAIL.n80 9.3005
R305 VTAIL.n66 VTAIL.n65 9.3005
R306 VTAIL.n75 VTAIL.n74 9.3005
R307 VTAIL.n73 VTAIL.n72 9.3005
R308 VTAIL.n0 VTAIL.t1 8.55445
R309 VTAIL.n0 VTAIL.t4 8.55445
R310 VTAIL.n42 VTAIL.t8 8.55445
R311 VTAIL.n42 VTAIL.t13 8.55445
R312 VTAIL.n126 VTAIL.t14 8.55445
R313 VTAIL.n126 VTAIL.t11 8.55445
R314 VTAIL.n84 VTAIL.t6 8.55445
R315 VTAIL.n84 VTAIL.t2 8.55445
R316 VTAIL.n157 VTAIL.n153 3.78097
R317 VTAIL.n11 VTAIL.n7 3.78097
R318 VTAIL.n31 VTAIL.n27 3.78097
R319 VTAIL.n53 VTAIL.n49 3.78097
R320 VTAIL.n137 VTAIL.n133 3.78097
R321 VTAIL.n115 VTAIL.n111 3.78097
R322 VTAIL.n95 VTAIL.n91 3.78097
R323 VTAIL.n73 VTAIL.n69 3.78097
R324 VTAIL.n166 VTAIL.n148 3.49141
R325 VTAIL.n20 VTAIL.n2 3.49141
R326 VTAIL.n40 VTAIL.n22 3.49141
R327 VTAIL.n62 VTAIL.n44 3.49141
R328 VTAIL.n146 VTAIL.n128 3.49141
R329 VTAIL.n124 VTAIL.n106 3.49141
R330 VTAIL.n104 VTAIL.n86 3.49141
R331 VTAIL.n82 VTAIL.n64 3.49141
R332 VTAIL.n85 VTAIL.n83 2.75912
R333 VTAIL.n105 VTAIL.n85 2.75912
R334 VTAIL.n127 VTAIL.n125 2.75912
R335 VTAIL.n147 VTAIL.n127 2.75912
R336 VTAIL.n63 VTAIL.n43 2.75912
R337 VTAIL.n43 VTAIL.n41 2.75912
R338 VTAIL.n21 VTAIL.n1 2.75912
R339 VTAIL.n164 VTAIL.n163 2.71565
R340 VTAIL.n18 VTAIL.n17 2.71565
R341 VTAIL.n38 VTAIL.n37 2.71565
R342 VTAIL.n60 VTAIL.n59 2.71565
R343 VTAIL.n144 VTAIL.n143 2.71565
R344 VTAIL.n122 VTAIL.n121 2.71565
R345 VTAIL.n102 VTAIL.n101 2.71565
R346 VTAIL.n80 VTAIL.n79 2.71565
R347 VTAIL VTAIL.n167 2.70093
R348 VTAIL.n160 VTAIL.n150 1.93989
R349 VTAIL.n14 VTAIL.n4 1.93989
R350 VTAIL.n34 VTAIL.n24 1.93989
R351 VTAIL.n56 VTAIL.n46 1.93989
R352 VTAIL.n140 VTAIL.n130 1.93989
R353 VTAIL.n118 VTAIL.n108 1.93989
R354 VTAIL.n98 VTAIL.n88 1.93989
R355 VTAIL.n76 VTAIL.n66 1.93989
R356 VTAIL.n159 VTAIL.n152 1.16414
R357 VTAIL.n13 VTAIL.n6 1.16414
R358 VTAIL.n33 VTAIL.n26 1.16414
R359 VTAIL.n55 VTAIL.n48 1.16414
R360 VTAIL.n139 VTAIL.n132 1.16414
R361 VTAIL.n117 VTAIL.n110 1.16414
R362 VTAIL.n97 VTAIL.n90 1.16414
R363 VTAIL.n75 VTAIL.n68 1.16414
R364 VTAIL.n125 VTAIL.n105 0.470328
R365 VTAIL.n41 VTAIL.n21 0.470328
R366 VTAIL.n156 VTAIL.n155 0.388379
R367 VTAIL.n10 VTAIL.n9 0.388379
R368 VTAIL.n30 VTAIL.n29 0.388379
R369 VTAIL.n52 VTAIL.n51 0.388379
R370 VTAIL.n136 VTAIL.n135 0.388379
R371 VTAIL.n114 VTAIL.n113 0.388379
R372 VTAIL.n94 VTAIL.n93 0.388379
R373 VTAIL.n72 VTAIL.n71 0.388379
R374 VTAIL.n158 VTAIL.n157 0.155672
R375 VTAIL.n158 VTAIL.n149 0.155672
R376 VTAIL.n165 VTAIL.n149 0.155672
R377 VTAIL.n12 VTAIL.n11 0.155672
R378 VTAIL.n12 VTAIL.n3 0.155672
R379 VTAIL.n19 VTAIL.n3 0.155672
R380 VTAIL.n32 VTAIL.n31 0.155672
R381 VTAIL.n32 VTAIL.n23 0.155672
R382 VTAIL.n39 VTAIL.n23 0.155672
R383 VTAIL.n54 VTAIL.n53 0.155672
R384 VTAIL.n54 VTAIL.n45 0.155672
R385 VTAIL.n61 VTAIL.n45 0.155672
R386 VTAIL.n145 VTAIL.n129 0.155672
R387 VTAIL.n138 VTAIL.n129 0.155672
R388 VTAIL.n138 VTAIL.n137 0.155672
R389 VTAIL.n123 VTAIL.n107 0.155672
R390 VTAIL.n116 VTAIL.n107 0.155672
R391 VTAIL.n116 VTAIL.n115 0.155672
R392 VTAIL.n103 VTAIL.n87 0.155672
R393 VTAIL.n96 VTAIL.n87 0.155672
R394 VTAIL.n96 VTAIL.n95 0.155672
R395 VTAIL.n81 VTAIL.n65 0.155672
R396 VTAIL.n74 VTAIL.n65 0.155672
R397 VTAIL.n74 VTAIL.n73 0.155672
R398 VTAIL VTAIL.n1 0.0586897
R399 B.n484 B.n483 585
R400 B.n485 B.n56 585
R401 B.n487 B.n486 585
R402 B.n488 B.n55 585
R403 B.n490 B.n489 585
R404 B.n491 B.n54 585
R405 B.n493 B.n492 585
R406 B.n494 B.n53 585
R407 B.n496 B.n495 585
R408 B.n497 B.n52 585
R409 B.n499 B.n498 585
R410 B.n500 B.n51 585
R411 B.n502 B.n501 585
R412 B.n503 B.n50 585
R413 B.n505 B.n504 585
R414 B.n506 B.n49 585
R415 B.n508 B.n507 585
R416 B.n509 B.n46 585
R417 B.n512 B.n511 585
R418 B.n513 B.n45 585
R419 B.n515 B.n514 585
R420 B.n516 B.n44 585
R421 B.n518 B.n517 585
R422 B.n519 B.n43 585
R423 B.n521 B.n520 585
R424 B.n522 B.n39 585
R425 B.n524 B.n523 585
R426 B.n525 B.n38 585
R427 B.n527 B.n526 585
R428 B.n528 B.n37 585
R429 B.n530 B.n529 585
R430 B.n531 B.n36 585
R431 B.n533 B.n532 585
R432 B.n534 B.n35 585
R433 B.n536 B.n535 585
R434 B.n537 B.n34 585
R435 B.n539 B.n538 585
R436 B.n540 B.n33 585
R437 B.n542 B.n541 585
R438 B.n543 B.n32 585
R439 B.n545 B.n544 585
R440 B.n546 B.n31 585
R441 B.n548 B.n547 585
R442 B.n549 B.n30 585
R443 B.n551 B.n550 585
R444 B.n482 B.n57 585
R445 B.n481 B.n480 585
R446 B.n479 B.n58 585
R447 B.n478 B.n477 585
R448 B.n476 B.n59 585
R449 B.n475 B.n474 585
R450 B.n473 B.n60 585
R451 B.n472 B.n471 585
R452 B.n470 B.n61 585
R453 B.n469 B.n468 585
R454 B.n467 B.n62 585
R455 B.n466 B.n465 585
R456 B.n464 B.n63 585
R457 B.n463 B.n462 585
R458 B.n461 B.n64 585
R459 B.n460 B.n459 585
R460 B.n458 B.n65 585
R461 B.n457 B.n456 585
R462 B.n455 B.n66 585
R463 B.n454 B.n453 585
R464 B.n452 B.n67 585
R465 B.n451 B.n450 585
R466 B.n449 B.n68 585
R467 B.n448 B.n447 585
R468 B.n446 B.n69 585
R469 B.n445 B.n444 585
R470 B.n443 B.n70 585
R471 B.n442 B.n441 585
R472 B.n440 B.n71 585
R473 B.n439 B.n438 585
R474 B.n437 B.n72 585
R475 B.n436 B.n435 585
R476 B.n434 B.n73 585
R477 B.n433 B.n432 585
R478 B.n431 B.n74 585
R479 B.n430 B.n429 585
R480 B.n428 B.n75 585
R481 B.n427 B.n426 585
R482 B.n425 B.n76 585
R483 B.n424 B.n423 585
R484 B.n422 B.n77 585
R485 B.n421 B.n420 585
R486 B.n419 B.n78 585
R487 B.n418 B.n417 585
R488 B.n416 B.n79 585
R489 B.n415 B.n414 585
R490 B.n413 B.n80 585
R491 B.n412 B.n411 585
R492 B.n410 B.n81 585
R493 B.n409 B.n408 585
R494 B.n407 B.n82 585
R495 B.n406 B.n405 585
R496 B.n404 B.n83 585
R497 B.n403 B.n402 585
R498 B.n401 B.n84 585
R499 B.n400 B.n399 585
R500 B.n398 B.n85 585
R501 B.n397 B.n396 585
R502 B.n395 B.n86 585
R503 B.n394 B.n393 585
R504 B.n392 B.n87 585
R505 B.n391 B.n390 585
R506 B.n389 B.n88 585
R507 B.n388 B.n387 585
R508 B.n386 B.n89 585
R509 B.n385 B.n384 585
R510 B.n383 B.n90 585
R511 B.n382 B.n381 585
R512 B.n380 B.n91 585
R513 B.n379 B.n378 585
R514 B.n377 B.n92 585
R515 B.n376 B.n375 585
R516 B.n374 B.n93 585
R517 B.n373 B.n372 585
R518 B.n371 B.n94 585
R519 B.n370 B.n369 585
R520 B.n368 B.n95 585
R521 B.n367 B.n366 585
R522 B.n365 B.n96 585
R523 B.n364 B.n363 585
R524 B.n362 B.n97 585
R525 B.n361 B.n360 585
R526 B.n359 B.n98 585
R527 B.n358 B.n357 585
R528 B.n356 B.n99 585
R529 B.n355 B.n354 585
R530 B.n353 B.n100 585
R531 B.n352 B.n351 585
R532 B.n350 B.n101 585
R533 B.n349 B.n348 585
R534 B.n347 B.n102 585
R535 B.n346 B.n345 585
R536 B.n344 B.n103 585
R537 B.n343 B.n342 585
R538 B.n341 B.n104 585
R539 B.n340 B.n339 585
R540 B.n338 B.n105 585
R541 B.n337 B.n336 585
R542 B.n335 B.n106 585
R543 B.n334 B.n333 585
R544 B.n332 B.n107 585
R545 B.n331 B.n330 585
R546 B.n329 B.n108 585
R547 B.n328 B.n327 585
R548 B.n326 B.n109 585
R549 B.n325 B.n324 585
R550 B.n323 B.n110 585
R551 B.n322 B.n321 585
R552 B.n320 B.n111 585
R553 B.n319 B.n318 585
R554 B.n317 B.n112 585
R555 B.n246 B.n245 585
R556 B.n247 B.n136 585
R557 B.n249 B.n248 585
R558 B.n250 B.n135 585
R559 B.n252 B.n251 585
R560 B.n253 B.n134 585
R561 B.n255 B.n254 585
R562 B.n256 B.n133 585
R563 B.n258 B.n257 585
R564 B.n259 B.n132 585
R565 B.n261 B.n260 585
R566 B.n262 B.n131 585
R567 B.n264 B.n263 585
R568 B.n265 B.n130 585
R569 B.n267 B.n266 585
R570 B.n268 B.n129 585
R571 B.n270 B.n269 585
R572 B.n271 B.n126 585
R573 B.n274 B.n273 585
R574 B.n275 B.n125 585
R575 B.n277 B.n276 585
R576 B.n278 B.n124 585
R577 B.n280 B.n279 585
R578 B.n281 B.n123 585
R579 B.n283 B.n282 585
R580 B.n284 B.n122 585
R581 B.n289 B.n288 585
R582 B.n290 B.n121 585
R583 B.n292 B.n291 585
R584 B.n293 B.n120 585
R585 B.n295 B.n294 585
R586 B.n296 B.n119 585
R587 B.n298 B.n297 585
R588 B.n299 B.n118 585
R589 B.n301 B.n300 585
R590 B.n302 B.n117 585
R591 B.n304 B.n303 585
R592 B.n305 B.n116 585
R593 B.n307 B.n306 585
R594 B.n308 B.n115 585
R595 B.n310 B.n309 585
R596 B.n311 B.n114 585
R597 B.n313 B.n312 585
R598 B.n314 B.n113 585
R599 B.n316 B.n315 585
R600 B.n244 B.n137 585
R601 B.n243 B.n242 585
R602 B.n241 B.n138 585
R603 B.n240 B.n239 585
R604 B.n238 B.n139 585
R605 B.n237 B.n236 585
R606 B.n235 B.n140 585
R607 B.n234 B.n233 585
R608 B.n232 B.n141 585
R609 B.n231 B.n230 585
R610 B.n229 B.n142 585
R611 B.n228 B.n227 585
R612 B.n226 B.n143 585
R613 B.n225 B.n224 585
R614 B.n223 B.n144 585
R615 B.n222 B.n221 585
R616 B.n220 B.n145 585
R617 B.n219 B.n218 585
R618 B.n217 B.n146 585
R619 B.n216 B.n215 585
R620 B.n214 B.n147 585
R621 B.n213 B.n212 585
R622 B.n211 B.n148 585
R623 B.n210 B.n209 585
R624 B.n208 B.n149 585
R625 B.n207 B.n206 585
R626 B.n205 B.n150 585
R627 B.n204 B.n203 585
R628 B.n202 B.n151 585
R629 B.n201 B.n200 585
R630 B.n199 B.n152 585
R631 B.n198 B.n197 585
R632 B.n196 B.n153 585
R633 B.n195 B.n194 585
R634 B.n193 B.n154 585
R635 B.n192 B.n191 585
R636 B.n190 B.n155 585
R637 B.n189 B.n188 585
R638 B.n187 B.n156 585
R639 B.n186 B.n185 585
R640 B.n184 B.n157 585
R641 B.n183 B.n182 585
R642 B.n181 B.n158 585
R643 B.n180 B.n179 585
R644 B.n178 B.n159 585
R645 B.n177 B.n176 585
R646 B.n175 B.n160 585
R647 B.n174 B.n173 585
R648 B.n172 B.n161 585
R649 B.n171 B.n170 585
R650 B.n169 B.n162 585
R651 B.n168 B.n167 585
R652 B.n166 B.n163 585
R653 B.n165 B.n164 585
R654 B.n2 B.n0 585
R655 B.n633 B.n1 585
R656 B.n632 B.n631 585
R657 B.n630 B.n3 585
R658 B.n629 B.n628 585
R659 B.n627 B.n4 585
R660 B.n626 B.n625 585
R661 B.n624 B.n5 585
R662 B.n623 B.n622 585
R663 B.n621 B.n6 585
R664 B.n620 B.n619 585
R665 B.n618 B.n7 585
R666 B.n617 B.n616 585
R667 B.n615 B.n8 585
R668 B.n614 B.n613 585
R669 B.n612 B.n9 585
R670 B.n611 B.n610 585
R671 B.n609 B.n10 585
R672 B.n608 B.n607 585
R673 B.n606 B.n11 585
R674 B.n605 B.n604 585
R675 B.n603 B.n12 585
R676 B.n602 B.n601 585
R677 B.n600 B.n13 585
R678 B.n599 B.n598 585
R679 B.n597 B.n14 585
R680 B.n596 B.n595 585
R681 B.n594 B.n15 585
R682 B.n593 B.n592 585
R683 B.n591 B.n16 585
R684 B.n590 B.n589 585
R685 B.n588 B.n17 585
R686 B.n587 B.n586 585
R687 B.n585 B.n18 585
R688 B.n584 B.n583 585
R689 B.n582 B.n19 585
R690 B.n581 B.n580 585
R691 B.n579 B.n20 585
R692 B.n578 B.n577 585
R693 B.n576 B.n21 585
R694 B.n575 B.n574 585
R695 B.n573 B.n22 585
R696 B.n572 B.n571 585
R697 B.n570 B.n23 585
R698 B.n569 B.n568 585
R699 B.n567 B.n24 585
R700 B.n566 B.n565 585
R701 B.n564 B.n25 585
R702 B.n563 B.n562 585
R703 B.n561 B.n26 585
R704 B.n560 B.n559 585
R705 B.n558 B.n27 585
R706 B.n557 B.n556 585
R707 B.n555 B.n28 585
R708 B.n554 B.n553 585
R709 B.n552 B.n29 585
R710 B.n635 B.n634 585
R711 B.n245 B.n244 492.5
R712 B.n550 B.n29 492.5
R713 B.n315 B.n112 492.5
R714 B.n483 B.n482 492.5
R715 B.n285 B.t8 293.812
R716 B.n47 B.t10 293.812
R717 B.n127 B.t5 293.812
R718 B.n40 B.t1 293.812
R719 B.n285 B.t6 240.331
R720 B.n127 B.t3 240.331
R721 B.n40 B.t0 240.331
R722 B.n47 B.t9 240.331
R723 B.n286 B.t7 231.75
R724 B.n48 B.t11 231.75
R725 B.n128 B.t4 231.75
R726 B.n41 B.t2 231.75
R727 B.n244 B.n243 163.367
R728 B.n243 B.n138 163.367
R729 B.n239 B.n138 163.367
R730 B.n239 B.n238 163.367
R731 B.n238 B.n237 163.367
R732 B.n237 B.n140 163.367
R733 B.n233 B.n140 163.367
R734 B.n233 B.n232 163.367
R735 B.n232 B.n231 163.367
R736 B.n231 B.n142 163.367
R737 B.n227 B.n142 163.367
R738 B.n227 B.n226 163.367
R739 B.n226 B.n225 163.367
R740 B.n225 B.n144 163.367
R741 B.n221 B.n144 163.367
R742 B.n221 B.n220 163.367
R743 B.n220 B.n219 163.367
R744 B.n219 B.n146 163.367
R745 B.n215 B.n146 163.367
R746 B.n215 B.n214 163.367
R747 B.n214 B.n213 163.367
R748 B.n213 B.n148 163.367
R749 B.n209 B.n148 163.367
R750 B.n209 B.n208 163.367
R751 B.n208 B.n207 163.367
R752 B.n207 B.n150 163.367
R753 B.n203 B.n150 163.367
R754 B.n203 B.n202 163.367
R755 B.n202 B.n201 163.367
R756 B.n201 B.n152 163.367
R757 B.n197 B.n152 163.367
R758 B.n197 B.n196 163.367
R759 B.n196 B.n195 163.367
R760 B.n195 B.n154 163.367
R761 B.n191 B.n154 163.367
R762 B.n191 B.n190 163.367
R763 B.n190 B.n189 163.367
R764 B.n189 B.n156 163.367
R765 B.n185 B.n156 163.367
R766 B.n185 B.n184 163.367
R767 B.n184 B.n183 163.367
R768 B.n183 B.n158 163.367
R769 B.n179 B.n158 163.367
R770 B.n179 B.n178 163.367
R771 B.n178 B.n177 163.367
R772 B.n177 B.n160 163.367
R773 B.n173 B.n160 163.367
R774 B.n173 B.n172 163.367
R775 B.n172 B.n171 163.367
R776 B.n171 B.n162 163.367
R777 B.n167 B.n162 163.367
R778 B.n167 B.n166 163.367
R779 B.n166 B.n165 163.367
R780 B.n165 B.n2 163.367
R781 B.n634 B.n2 163.367
R782 B.n634 B.n633 163.367
R783 B.n633 B.n632 163.367
R784 B.n632 B.n3 163.367
R785 B.n628 B.n3 163.367
R786 B.n628 B.n627 163.367
R787 B.n627 B.n626 163.367
R788 B.n626 B.n5 163.367
R789 B.n622 B.n5 163.367
R790 B.n622 B.n621 163.367
R791 B.n621 B.n620 163.367
R792 B.n620 B.n7 163.367
R793 B.n616 B.n7 163.367
R794 B.n616 B.n615 163.367
R795 B.n615 B.n614 163.367
R796 B.n614 B.n9 163.367
R797 B.n610 B.n9 163.367
R798 B.n610 B.n609 163.367
R799 B.n609 B.n608 163.367
R800 B.n608 B.n11 163.367
R801 B.n604 B.n11 163.367
R802 B.n604 B.n603 163.367
R803 B.n603 B.n602 163.367
R804 B.n602 B.n13 163.367
R805 B.n598 B.n13 163.367
R806 B.n598 B.n597 163.367
R807 B.n597 B.n596 163.367
R808 B.n596 B.n15 163.367
R809 B.n592 B.n15 163.367
R810 B.n592 B.n591 163.367
R811 B.n591 B.n590 163.367
R812 B.n590 B.n17 163.367
R813 B.n586 B.n17 163.367
R814 B.n586 B.n585 163.367
R815 B.n585 B.n584 163.367
R816 B.n584 B.n19 163.367
R817 B.n580 B.n19 163.367
R818 B.n580 B.n579 163.367
R819 B.n579 B.n578 163.367
R820 B.n578 B.n21 163.367
R821 B.n574 B.n21 163.367
R822 B.n574 B.n573 163.367
R823 B.n573 B.n572 163.367
R824 B.n572 B.n23 163.367
R825 B.n568 B.n23 163.367
R826 B.n568 B.n567 163.367
R827 B.n567 B.n566 163.367
R828 B.n566 B.n25 163.367
R829 B.n562 B.n25 163.367
R830 B.n562 B.n561 163.367
R831 B.n561 B.n560 163.367
R832 B.n560 B.n27 163.367
R833 B.n556 B.n27 163.367
R834 B.n556 B.n555 163.367
R835 B.n555 B.n554 163.367
R836 B.n554 B.n29 163.367
R837 B.n245 B.n136 163.367
R838 B.n249 B.n136 163.367
R839 B.n250 B.n249 163.367
R840 B.n251 B.n250 163.367
R841 B.n251 B.n134 163.367
R842 B.n255 B.n134 163.367
R843 B.n256 B.n255 163.367
R844 B.n257 B.n256 163.367
R845 B.n257 B.n132 163.367
R846 B.n261 B.n132 163.367
R847 B.n262 B.n261 163.367
R848 B.n263 B.n262 163.367
R849 B.n263 B.n130 163.367
R850 B.n267 B.n130 163.367
R851 B.n268 B.n267 163.367
R852 B.n269 B.n268 163.367
R853 B.n269 B.n126 163.367
R854 B.n274 B.n126 163.367
R855 B.n275 B.n274 163.367
R856 B.n276 B.n275 163.367
R857 B.n276 B.n124 163.367
R858 B.n280 B.n124 163.367
R859 B.n281 B.n280 163.367
R860 B.n282 B.n281 163.367
R861 B.n282 B.n122 163.367
R862 B.n289 B.n122 163.367
R863 B.n290 B.n289 163.367
R864 B.n291 B.n290 163.367
R865 B.n291 B.n120 163.367
R866 B.n295 B.n120 163.367
R867 B.n296 B.n295 163.367
R868 B.n297 B.n296 163.367
R869 B.n297 B.n118 163.367
R870 B.n301 B.n118 163.367
R871 B.n302 B.n301 163.367
R872 B.n303 B.n302 163.367
R873 B.n303 B.n116 163.367
R874 B.n307 B.n116 163.367
R875 B.n308 B.n307 163.367
R876 B.n309 B.n308 163.367
R877 B.n309 B.n114 163.367
R878 B.n313 B.n114 163.367
R879 B.n314 B.n313 163.367
R880 B.n315 B.n314 163.367
R881 B.n319 B.n112 163.367
R882 B.n320 B.n319 163.367
R883 B.n321 B.n320 163.367
R884 B.n321 B.n110 163.367
R885 B.n325 B.n110 163.367
R886 B.n326 B.n325 163.367
R887 B.n327 B.n326 163.367
R888 B.n327 B.n108 163.367
R889 B.n331 B.n108 163.367
R890 B.n332 B.n331 163.367
R891 B.n333 B.n332 163.367
R892 B.n333 B.n106 163.367
R893 B.n337 B.n106 163.367
R894 B.n338 B.n337 163.367
R895 B.n339 B.n338 163.367
R896 B.n339 B.n104 163.367
R897 B.n343 B.n104 163.367
R898 B.n344 B.n343 163.367
R899 B.n345 B.n344 163.367
R900 B.n345 B.n102 163.367
R901 B.n349 B.n102 163.367
R902 B.n350 B.n349 163.367
R903 B.n351 B.n350 163.367
R904 B.n351 B.n100 163.367
R905 B.n355 B.n100 163.367
R906 B.n356 B.n355 163.367
R907 B.n357 B.n356 163.367
R908 B.n357 B.n98 163.367
R909 B.n361 B.n98 163.367
R910 B.n362 B.n361 163.367
R911 B.n363 B.n362 163.367
R912 B.n363 B.n96 163.367
R913 B.n367 B.n96 163.367
R914 B.n368 B.n367 163.367
R915 B.n369 B.n368 163.367
R916 B.n369 B.n94 163.367
R917 B.n373 B.n94 163.367
R918 B.n374 B.n373 163.367
R919 B.n375 B.n374 163.367
R920 B.n375 B.n92 163.367
R921 B.n379 B.n92 163.367
R922 B.n380 B.n379 163.367
R923 B.n381 B.n380 163.367
R924 B.n381 B.n90 163.367
R925 B.n385 B.n90 163.367
R926 B.n386 B.n385 163.367
R927 B.n387 B.n386 163.367
R928 B.n387 B.n88 163.367
R929 B.n391 B.n88 163.367
R930 B.n392 B.n391 163.367
R931 B.n393 B.n392 163.367
R932 B.n393 B.n86 163.367
R933 B.n397 B.n86 163.367
R934 B.n398 B.n397 163.367
R935 B.n399 B.n398 163.367
R936 B.n399 B.n84 163.367
R937 B.n403 B.n84 163.367
R938 B.n404 B.n403 163.367
R939 B.n405 B.n404 163.367
R940 B.n405 B.n82 163.367
R941 B.n409 B.n82 163.367
R942 B.n410 B.n409 163.367
R943 B.n411 B.n410 163.367
R944 B.n411 B.n80 163.367
R945 B.n415 B.n80 163.367
R946 B.n416 B.n415 163.367
R947 B.n417 B.n416 163.367
R948 B.n417 B.n78 163.367
R949 B.n421 B.n78 163.367
R950 B.n422 B.n421 163.367
R951 B.n423 B.n422 163.367
R952 B.n423 B.n76 163.367
R953 B.n427 B.n76 163.367
R954 B.n428 B.n427 163.367
R955 B.n429 B.n428 163.367
R956 B.n429 B.n74 163.367
R957 B.n433 B.n74 163.367
R958 B.n434 B.n433 163.367
R959 B.n435 B.n434 163.367
R960 B.n435 B.n72 163.367
R961 B.n439 B.n72 163.367
R962 B.n440 B.n439 163.367
R963 B.n441 B.n440 163.367
R964 B.n441 B.n70 163.367
R965 B.n445 B.n70 163.367
R966 B.n446 B.n445 163.367
R967 B.n447 B.n446 163.367
R968 B.n447 B.n68 163.367
R969 B.n451 B.n68 163.367
R970 B.n452 B.n451 163.367
R971 B.n453 B.n452 163.367
R972 B.n453 B.n66 163.367
R973 B.n457 B.n66 163.367
R974 B.n458 B.n457 163.367
R975 B.n459 B.n458 163.367
R976 B.n459 B.n64 163.367
R977 B.n463 B.n64 163.367
R978 B.n464 B.n463 163.367
R979 B.n465 B.n464 163.367
R980 B.n465 B.n62 163.367
R981 B.n469 B.n62 163.367
R982 B.n470 B.n469 163.367
R983 B.n471 B.n470 163.367
R984 B.n471 B.n60 163.367
R985 B.n475 B.n60 163.367
R986 B.n476 B.n475 163.367
R987 B.n477 B.n476 163.367
R988 B.n477 B.n58 163.367
R989 B.n481 B.n58 163.367
R990 B.n482 B.n481 163.367
R991 B.n550 B.n549 163.367
R992 B.n549 B.n548 163.367
R993 B.n548 B.n31 163.367
R994 B.n544 B.n31 163.367
R995 B.n544 B.n543 163.367
R996 B.n543 B.n542 163.367
R997 B.n542 B.n33 163.367
R998 B.n538 B.n33 163.367
R999 B.n538 B.n537 163.367
R1000 B.n537 B.n536 163.367
R1001 B.n536 B.n35 163.367
R1002 B.n532 B.n35 163.367
R1003 B.n532 B.n531 163.367
R1004 B.n531 B.n530 163.367
R1005 B.n530 B.n37 163.367
R1006 B.n526 B.n37 163.367
R1007 B.n526 B.n525 163.367
R1008 B.n525 B.n524 163.367
R1009 B.n524 B.n39 163.367
R1010 B.n520 B.n39 163.367
R1011 B.n520 B.n519 163.367
R1012 B.n519 B.n518 163.367
R1013 B.n518 B.n44 163.367
R1014 B.n514 B.n44 163.367
R1015 B.n514 B.n513 163.367
R1016 B.n513 B.n512 163.367
R1017 B.n512 B.n46 163.367
R1018 B.n507 B.n46 163.367
R1019 B.n507 B.n506 163.367
R1020 B.n506 B.n505 163.367
R1021 B.n505 B.n50 163.367
R1022 B.n501 B.n50 163.367
R1023 B.n501 B.n500 163.367
R1024 B.n500 B.n499 163.367
R1025 B.n499 B.n52 163.367
R1026 B.n495 B.n52 163.367
R1027 B.n495 B.n494 163.367
R1028 B.n494 B.n493 163.367
R1029 B.n493 B.n54 163.367
R1030 B.n489 B.n54 163.367
R1031 B.n489 B.n488 163.367
R1032 B.n488 B.n487 163.367
R1033 B.n487 B.n56 163.367
R1034 B.n483 B.n56 163.367
R1035 B.n286 B.n285 62.0611
R1036 B.n128 B.n127 62.0611
R1037 B.n41 B.n40 62.0611
R1038 B.n48 B.n47 62.0611
R1039 B.n287 B.n286 59.5399
R1040 B.n272 B.n128 59.5399
R1041 B.n42 B.n41 59.5399
R1042 B.n510 B.n48 59.5399
R1043 B.n552 B.n551 32.0005
R1044 B.n484 B.n57 32.0005
R1045 B.n317 B.n316 32.0005
R1046 B.n246 B.n137 32.0005
R1047 B B.n635 18.0485
R1048 B.n551 B.n30 10.6151
R1049 B.n547 B.n30 10.6151
R1050 B.n547 B.n546 10.6151
R1051 B.n546 B.n545 10.6151
R1052 B.n545 B.n32 10.6151
R1053 B.n541 B.n32 10.6151
R1054 B.n541 B.n540 10.6151
R1055 B.n540 B.n539 10.6151
R1056 B.n539 B.n34 10.6151
R1057 B.n535 B.n34 10.6151
R1058 B.n535 B.n534 10.6151
R1059 B.n534 B.n533 10.6151
R1060 B.n533 B.n36 10.6151
R1061 B.n529 B.n36 10.6151
R1062 B.n529 B.n528 10.6151
R1063 B.n528 B.n527 10.6151
R1064 B.n527 B.n38 10.6151
R1065 B.n523 B.n522 10.6151
R1066 B.n522 B.n521 10.6151
R1067 B.n521 B.n43 10.6151
R1068 B.n517 B.n43 10.6151
R1069 B.n517 B.n516 10.6151
R1070 B.n516 B.n515 10.6151
R1071 B.n515 B.n45 10.6151
R1072 B.n511 B.n45 10.6151
R1073 B.n509 B.n508 10.6151
R1074 B.n508 B.n49 10.6151
R1075 B.n504 B.n49 10.6151
R1076 B.n504 B.n503 10.6151
R1077 B.n503 B.n502 10.6151
R1078 B.n502 B.n51 10.6151
R1079 B.n498 B.n51 10.6151
R1080 B.n498 B.n497 10.6151
R1081 B.n497 B.n496 10.6151
R1082 B.n496 B.n53 10.6151
R1083 B.n492 B.n53 10.6151
R1084 B.n492 B.n491 10.6151
R1085 B.n491 B.n490 10.6151
R1086 B.n490 B.n55 10.6151
R1087 B.n486 B.n55 10.6151
R1088 B.n486 B.n485 10.6151
R1089 B.n485 B.n484 10.6151
R1090 B.n318 B.n317 10.6151
R1091 B.n318 B.n111 10.6151
R1092 B.n322 B.n111 10.6151
R1093 B.n323 B.n322 10.6151
R1094 B.n324 B.n323 10.6151
R1095 B.n324 B.n109 10.6151
R1096 B.n328 B.n109 10.6151
R1097 B.n329 B.n328 10.6151
R1098 B.n330 B.n329 10.6151
R1099 B.n330 B.n107 10.6151
R1100 B.n334 B.n107 10.6151
R1101 B.n335 B.n334 10.6151
R1102 B.n336 B.n335 10.6151
R1103 B.n336 B.n105 10.6151
R1104 B.n340 B.n105 10.6151
R1105 B.n341 B.n340 10.6151
R1106 B.n342 B.n341 10.6151
R1107 B.n342 B.n103 10.6151
R1108 B.n346 B.n103 10.6151
R1109 B.n347 B.n346 10.6151
R1110 B.n348 B.n347 10.6151
R1111 B.n348 B.n101 10.6151
R1112 B.n352 B.n101 10.6151
R1113 B.n353 B.n352 10.6151
R1114 B.n354 B.n353 10.6151
R1115 B.n354 B.n99 10.6151
R1116 B.n358 B.n99 10.6151
R1117 B.n359 B.n358 10.6151
R1118 B.n360 B.n359 10.6151
R1119 B.n360 B.n97 10.6151
R1120 B.n364 B.n97 10.6151
R1121 B.n365 B.n364 10.6151
R1122 B.n366 B.n365 10.6151
R1123 B.n366 B.n95 10.6151
R1124 B.n370 B.n95 10.6151
R1125 B.n371 B.n370 10.6151
R1126 B.n372 B.n371 10.6151
R1127 B.n372 B.n93 10.6151
R1128 B.n376 B.n93 10.6151
R1129 B.n377 B.n376 10.6151
R1130 B.n378 B.n377 10.6151
R1131 B.n378 B.n91 10.6151
R1132 B.n382 B.n91 10.6151
R1133 B.n383 B.n382 10.6151
R1134 B.n384 B.n383 10.6151
R1135 B.n384 B.n89 10.6151
R1136 B.n388 B.n89 10.6151
R1137 B.n389 B.n388 10.6151
R1138 B.n390 B.n389 10.6151
R1139 B.n390 B.n87 10.6151
R1140 B.n394 B.n87 10.6151
R1141 B.n395 B.n394 10.6151
R1142 B.n396 B.n395 10.6151
R1143 B.n396 B.n85 10.6151
R1144 B.n400 B.n85 10.6151
R1145 B.n401 B.n400 10.6151
R1146 B.n402 B.n401 10.6151
R1147 B.n402 B.n83 10.6151
R1148 B.n406 B.n83 10.6151
R1149 B.n407 B.n406 10.6151
R1150 B.n408 B.n407 10.6151
R1151 B.n408 B.n81 10.6151
R1152 B.n412 B.n81 10.6151
R1153 B.n413 B.n412 10.6151
R1154 B.n414 B.n413 10.6151
R1155 B.n414 B.n79 10.6151
R1156 B.n418 B.n79 10.6151
R1157 B.n419 B.n418 10.6151
R1158 B.n420 B.n419 10.6151
R1159 B.n420 B.n77 10.6151
R1160 B.n424 B.n77 10.6151
R1161 B.n425 B.n424 10.6151
R1162 B.n426 B.n425 10.6151
R1163 B.n426 B.n75 10.6151
R1164 B.n430 B.n75 10.6151
R1165 B.n431 B.n430 10.6151
R1166 B.n432 B.n431 10.6151
R1167 B.n432 B.n73 10.6151
R1168 B.n436 B.n73 10.6151
R1169 B.n437 B.n436 10.6151
R1170 B.n438 B.n437 10.6151
R1171 B.n438 B.n71 10.6151
R1172 B.n442 B.n71 10.6151
R1173 B.n443 B.n442 10.6151
R1174 B.n444 B.n443 10.6151
R1175 B.n444 B.n69 10.6151
R1176 B.n448 B.n69 10.6151
R1177 B.n449 B.n448 10.6151
R1178 B.n450 B.n449 10.6151
R1179 B.n450 B.n67 10.6151
R1180 B.n454 B.n67 10.6151
R1181 B.n455 B.n454 10.6151
R1182 B.n456 B.n455 10.6151
R1183 B.n456 B.n65 10.6151
R1184 B.n460 B.n65 10.6151
R1185 B.n461 B.n460 10.6151
R1186 B.n462 B.n461 10.6151
R1187 B.n462 B.n63 10.6151
R1188 B.n466 B.n63 10.6151
R1189 B.n467 B.n466 10.6151
R1190 B.n468 B.n467 10.6151
R1191 B.n468 B.n61 10.6151
R1192 B.n472 B.n61 10.6151
R1193 B.n473 B.n472 10.6151
R1194 B.n474 B.n473 10.6151
R1195 B.n474 B.n59 10.6151
R1196 B.n478 B.n59 10.6151
R1197 B.n479 B.n478 10.6151
R1198 B.n480 B.n479 10.6151
R1199 B.n480 B.n57 10.6151
R1200 B.n247 B.n246 10.6151
R1201 B.n248 B.n247 10.6151
R1202 B.n248 B.n135 10.6151
R1203 B.n252 B.n135 10.6151
R1204 B.n253 B.n252 10.6151
R1205 B.n254 B.n253 10.6151
R1206 B.n254 B.n133 10.6151
R1207 B.n258 B.n133 10.6151
R1208 B.n259 B.n258 10.6151
R1209 B.n260 B.n259 10.6151
R1210 B.n260 B.n131 10.6151
R1211 B.n264 B.n131 10.6151
R1212 B.n265 B.n264 10.6151
R1213 B.n266 B.n265 10.6151
R1214 B.n266 B.n129 10.6151
R1215 B.n270 B.n129 10.6151
R1216 B.n271 B.n270 10.6151
R1217 B.n273 B.n125 10.6151
R1218 B.n277 B.n125 10.6151
R1219 B.n278 B.n277 10.6151
R1220 B.n279 B.n278 10.6151
R1221 B.n279 B.n123 10.6151
R1222 B.n283 B.n123 10.6151
R1223 B.n284 B.n283 10.6151
R1224 B.n288 B.n284 10.6151
R1225 B.n292 B.n121 10.6151
R1226 B.n293 B.n292 10.6151
R1227 B.n294 B.n293 10.6151
R1228 B.n294 B.n119 10.6151
R1229 B.n298 B.n119 10.6151
R1230 B.n299 B.n298 10.6151
R1231 B.n300 B.n299 10.6151
R1232 B.n300 B.n117 10.6151
R1233 B.n304 B.n117 10.6151
R1234 B.n305 B.n304 10.6151
R1235 B.n306 B.n305 10.6151
R1236 B.n306 B.n115 10.6151
R1237 B.n310 B.n115 10.6151
R1238 B.n311 B.n310 10.6151
R1239 B.n312 B.n311 10.6151
R1240 B.n312 B.n113 10.6151
R1241 B.n316 B.n113 10.6151
R1242 B.n242 B.n137 10.6151
R1243 B.n242 B.n241 10.6151
R1244 B.n241 B.n240 10.6151
R1245 B.n240 B.n139 10.6151
R1246 B.n236 B.n139 10.6151
R1247 B.n236 B.n235 10.6151
R1248 B.n235 B.n234 10.6151
R1249 B.n234 B.n141 10.6151
R1250 B.n230 B.n141 10.6151
R1251 B.n230 B.n229 10.6151
R1252 B.n229 B.n228 10.6151
R1253 B.n228 B.n143 10.6151
R1254 B.n224 B.n143 10.6151
R1255 B.n224 B.n223 10.6151
R1256 B.n223 B.n222 10.6151
R1257 B.n222 B.n145 10.6151
R1258 B.n218 B.n145 10.6151
R1259 B.n218 B.n217 10.6151
R1260 B.n217 B.n216 10.6151
R1261 B.n216 B.n147 10.6151
R1262 B.n212 B.n147 10.6151
R1263 B.n212 B.n211 10.6151
R1264 B.n211 B.n210 10.6151
R1265 B.n210 B.n149 10.6151
R1266 B.n206 B.n149 10.6151
R1267 B.n206 B.n205 10.6151
R1268 B.n205 B.n204 10.6151
R1269 B.n204 B.n151 10.6151
R1270 B.n200 B.n151 10.6151
R1271 B.n200 B.n199 10.6151
R1272 B.n199 B.n198 10.6151
R1273 B.n198 B.n153 10.6151
R1274 B.n194 B.n153 10.6151
R1275 B.n194 B.n193 10.6151
R1276 B.n193 B.n192 10.6151
R1277 B.n192 B.n155 10.6151
R1278 B.n188 B.n155 10.6151
R1279 B.n188 B.n187 10.6151
R1280 B.n187 B.n186 10.6151
R1281 B.n186 B.n157 10.6151
R1282 B.n182 B.n157 10.6151
R1283 B.n182 B.n181 10.6151
R1284 B.n181 B.n180 10.6151
R1285 B.n180 B.n159 10.6151
R1286 B.n176 B.n159 10.6151
R1287 B.n176 B.n175 10.6151
R1288 B.n175 B.n174 10.6151
R1289 B.n174 B.n161 10.6151
R1290 B.n170 B.n161 10.6151
R1291 B.n170 B.n169 10.6151
R1292 B.n169 B.n168 10.6151
R1293 B.n168 B.n163 10.6151
R1294 B.n164 B.n163 10.6151
R1295 B.n164 B.n0 10.6151
R1296 B.n631 B.n1 10.6151
R1297 B.n631 B.n630 10.6151
R1298 B.n630 B.n629 10.6151
R1299 B.n629 B.n4 10.6151
R1300 B.n625 B.n4 10.6151
R1301 B.n625 B.n624 10.6151
R1302 B.n624 B.n623 10.6151
R1303 B.n623 B.n6 10.6151
R1304 B.n619 B.n6 10.6151
R1305 B.n619 B.n618 10.6151
R1306 B.n618 B.n617 10.6151
R1307 B.n617 B.n8 10.6151
R1308 B.n613 B.n8 10.6151
R1309 B.n613 B.n612 10.6151
R1310 B.n612 B.n611 10.6151
R1311 B.n611 B.n10 10.6151
R1312 B.n607 B.n10 10.6151
R1313 B.n607 B.n606 10.6151
R1314 B.n606 B.n605 10.6151
R1315 B.n605 B.n12 10.6151
R1316 B.n601 B.n12 10.6151
R1317 B.n601 B.n600 10.6151
R1318 B.n600 B.n599 10.6151
R1319 B.n599 B.n14 10.6151
R1320 B.n595 B.n14 10.6151
R1321 B.n595 B.n594 10.6151
R1322 B.n594 B.n593 10.6151
R1323 B.n593 B.n16 10.6151
R1324 B.n589 B.n16 10.6151
R1325 B.n589 B.n588 10.6151
R1326 B.n588 B.n587 10.6151
R1327 B.n587 B.n18 10.6151
R1328 B.n583 B.n18 10.6151
R1329 B.n583 B.n582 10.6151
R1330 B.n582 B.n581 10.6151
R1331 B.n581 B.n20 10.6151
R1332 B.n577 B.n20 10.6151
R1333 B.n577 B.n576 10.6151
R1334 B.n576 B.n575 10.6151
R1335 B.n575 B.n22 10.6151
R1336 B.n571 B.n22 10.6151
R1337 B.n571 B.n570 10.6151
R1338 B.n570 B.n569 10.6151
R1339 B.n569 B.n24 10.6151
R1340 B.n565 B.n24 10.6151
R1341 B.n565 B.n564 10.6151
R1342 B.n564 B.n563 10.6151
R1343 B.n563 B.n26 10.6151
R1344 B.n559 B.n26 10.6151
R1345 B.n559 B.n558 10.6151
R1346 B.n558 B.n557 10.6151
R1347 B.n557 B.n28 10.6151
R1348 B.n553 B.n28 10.6151
R1349 B.n553 B.n552 10.6151
R1350 B.n523 B.n42 6.5566
R1351 B.n511 B.n510 6.5566
R1352 B.n273 B.n272 6.5566
R1353 B.n288 B.n287 6.5566
R1354 B.n42 B.n38 4.05904
R1355 B.n510 B.n509 4.05904
R1356 B.n272 B.n271 4.05904
R1357 B.n287 B.n121 4.05904
R1358 B.n635 B.n0 2.81026
R1359 B.n635 B.n1 2.81026
R1360 VN.n59 VN.n31 161.3
R1361 VN.n58 VN.n57 161.3
R1362 VN.n56 VN.n32 161.3
R1363 VN.n55 VN.n54 161.3
R1364 VN.n53 VN.n33 161.3
R1365 VN.n52 VN.n51 161.3
R1366 VN.n50 VN.n34 161.3
R1367 VN.n49 VN.n48 161.3
R1368 VN.n47 VN.n35 161.3
R1369 VN.n46 VN.n45 161.3
R1370 VN.n44 VN.n37 161.3
R1371 VN.n43 VN.n42 161.3
R1372 VN.n41 VN.n38 161.3
R1373 VN.n28 VN.n0 161.3
R1374 VN.n27 VN.n26 161.3
R1375 VN.n25 VN.n1 161.3
R1376 VN.n24 VN.n23 161.3
R1377 VN.n22 VN.n2 161.3
R1378 VN.n21 VN.n20 161.3
R1379 VN.n19 VN.n3 161.3
R1380 VN.n18 VN.n17 161.3
R1381 VN.n15 VN.n4 161.3
R1382 VN.n14 VN.n13 161.3
R1383 VN.n12 VN.n5 161.3
R1384 VN.n11 VN.n10 161.3
R1385 VN.n9 VN.n6 161.3
R1386 VN.n30 VN.n29 108.45
R1387 VN.n61 VN.n60 108.45
R1388 VN.n7 VN.t2 64.9524
R1389 VN.n39 VN.t4 64.9524
R1390 VN.n8 VN.n7 56.7106
R1391 VN.n40 VN.n39 56.7106
R1392 VN.n14 VN.n5 56.5617
R1393 VN.n46 VN.n37 56.5617
R1394 VN VN.n61 46.1952
R1395 VN.n23 VN.n22 45.4209
R1396 VN.n54 VN.n53 45.4209
R1397 VN.n23 VN.n1 35.7332
R1398 VN.n54 VN.n32 35.7332
R1399 VN.n8 VN.t5 31.9099
R1400 VN.n16 VN.t0 31.9099
R1401 VN.n29 VN.t7 31.9099
R1402 VN.n40 VN.t6 31.9099
R1403 VN.n36 VN.t3 31.9099
R1404 VN.n60 VN.t1 31.9099
R1405 VN.n10 VN.n9 24.5923
R1406 VN.n10 VN.n5 24.5923
R1407 VN.n15 VN.n14 24.5923
R1408 VN.n17 VN.n15 24.5923
R1409 VN.n21 VN.n3 24.5923
R1410 VN.n22 VN.n21 24.5923
R1411 VN.n27 VN.n1 24.5923
R1412 VN.n28 VN.n27 24.5923
R1413 VN.n42 VN.n37 24.5923
R1414 VN.n42 VN.n41 24.5923
R1415 VN.n53 VN.n52 24.5923
R1416 VN.n52 VN.n34 24.5923
R1417 VN.n48 VN.n47 24.5923
R1418 VN.n47 VN.n46 24.5923
R1419 VN.n59 VN.n58 24.5923
R1420 VN.n58 VN.n32 24.5923
R1421 VN.n9 VN.n8 17.2148
R1422 VN.n17 VN.n16 17.2148
R1423 VN.n41 VN.n40 17.2148
R1424 VN.n48 VN.n36 17.2148
R1425 VN.n16 VN.n3 7.37805
R1426 VN.n36 VN.n34 7.37805
R1427 VN.n39 VN.n38 5.07592
R1428 VN.n7 VN.n6 5.07592
R1429 VN.n29 VN.n28 2.45968
R1430 VN.n60 VN.n59 2.45968
R1431 VN.n61 VN.n31 0.278335
R1432 VN.n30 VN.n0 0.278335
R1433 VN.n57 VN.n31 0.189894
R1434 VN.n57 VN.n56 0.189894
R1435 VN.n56 VN.n55 0.189894
R1436 VN.n55 VN.n33 0.189894
R1437 VN.n51 VN.n33 0.189894
R1438 VN.n51 VN.n50 0.189894
R1439 VN.n50 VN.n49 0.189894
R1440 VN.n49 VN.n35 0.189894
R1441 VN.n45 VN.n35 0.189894
R1442 VN.n45 VN.n44 0.189894
R1443 VN.n44 VN.n43 0.189894
R1444 VN.n43 VN.n38 0.189894
R1445 VN.n11 VN.n6 0.189894
R1446 VN.n12 VN.n11 0.189894
R1447 VN.n13 VN.n12 0.189894
R1448 VN.n13 VN.n4 0.189894
R1449 VN.n18 VN.n4 0.189894
R1450 VN.n19 VN.n18 0.189894
R1451 VN.n20 VN.n19 0.189894
R1452 VN.n20 VN.n2 0.189894
R1453 VN.n24 VN.n2 0.189894
R1454 VN.n25 VN.n24 0.189894
R1455 VN.n26 VN.n25 0.189894
R1456 VN.n26 VN.n0 0.189894
R1457 VN VN.n30 0.153485
R1458 VDD2.n2 VDD2.n1 114.117
R1459 VDD2.n2 VDD2.n0 114.117
R1460 VDD2 VDD2.n5 114.114
R1461 VDD2.n4 VDD2.n3 112.793
R1462 VDD2.n4 VDD2.n2 39.4049
R1463 VDD2.n5 VDD2.t1 8.55445
R1464 VDD2.n5 VDD2.t3 8.55445
R1465 VDD2.n3 VDD2.t6 8.55445
R1466 VDD2.n3 VDD2.t4 8.55445
R1467 VDD2.n1 VDD2.t7 8.55445
R1468 VDD2.n1 VDD2.t0 8.55445
R1469 VDD2.n0 VDD2.t5 8.55445
R1470 VDD2.n0 VDD2.t2 8.55445
R1471 VDD2 VDD2.n4 1.438
C0 B VN 1.22109f
C1 VDD2 B 1.61447f
C2 B VP 2.13112f
C3 VDD1 VN 0.15667f
C4 VTAIL VN 4.20386f
C5 VDD2 VDD1 1.91584f
C6 VDD1 VP 3.52032f
C7 VDD2 VTAIL 5.58702f
C8 VTAIL VP 4.21797f
C9 w_n4170_n1728# VN 8.40944f
C10 VDD2 w_n4170_n1728# 1.94126f
C11 w_n4170_n1728# VP 8.95043f
C12 VDD2 VN 3.12582f
C13 VP VN 6.47342f
C14 VDD1 B 1.50977f
C15 VTAIL B 2.32696f
C16 VDD2 VP 0.553511f
C17 w_n4170_n1728# B 8.25639f
C18 VDD1 VTAIL 5.53079f
C19 VDD1 w_n4170_n1728# 1.81562f
C20 w_n4170_n1728# VTAIL 2.38835f
C21 VDD2 VSUBS 1.535089f
C22 VDD1 VSUBS 2.242884f
C23 VTAIL VSUBS 0.661185f
C24 VN VSUBS 6.89548f
C25 VP VSUBS 3.275881f
C26 B VSUBS 4.344413f
C27 w_n4170_n1728# VSUBS 90.8226f
C28 VDD2.t5 VSUBS 0.072428f
C29 VDD2.t2 VSUBS 0.072428f
C30 VDD2.n0 VSUBS 0.423675f
C31 VDD2.t7 VSUBS 0.072428f
C32 VDD2.t0 VSUBS 0.072428f
C33 VDD2.n1 VSUBS 0.423675f
C34 VDD2.n2 VSUBS 3.10549f
C35 VDD2.t6 VSUBS 0.072428f
C36 VDD2.t4 VSUBS 0.072428f
C37 VDD2.n3 VSUBS 0.415997f
C38 VDD2.n4 VSUBS 2.46003f
C39 VDD2.t1 VSUBS 0.072428f
C40 VDD2.t3 VSUBS 0.072428f
C41 VDD2.n5 VSUBS 0.423651f
C42 VN.n0 VSUBS 0.054634f
C43 VN.t7 VSUBS 1.15551f
C44 VN.n1 VSUBS 0.083238f
C45 VN.n2 VSUBS 0.041442f
C46 VN.n3 VSUBS 0.050293f
C47 VN.n4 VSUBS 0.041442f
C48 VN.n5 VSUBS 0.060242f
C49 VN.n6 VSUBS 0.438092f
C50 VN.t5 VSUBS 1.15551f
C51 VN.t2 VSUBS 1.53138f
C52 VN.n7 VSUBS 0.5666f
C53 VN.n8 VSUBS 0.595759f
C54 VN.n9 VSUBS 0.065468f
C55 VN.n10 VSUBS 0.07685f
C56 VN.n11 VSUBS 0.041442f
C57 VN.n12 VSUBS 0.041442f
C58 VN.n13 VSUBS 0.041442f
C59 VN.n14 VSUBS 0.060242f
C60 VN.n15 VSUBS 0.07685f
C61 VN.t0 VSUBS 1.15551f
C62 VN.n16 VSUBS 0.460145f
C63 VN.n17 VSUBS 0.065468f
C64 VN.n18 VSUBS 0.041442f
C65 VN.n19 VSUBS 0.041442f
C66 VN.n20 VSUBS 0.041442f
C67 VN.n21 VSUBS 0.07685f
C68 VN.n22 VSUBS 0.079286f
C69 VN.n23 VSUBS 0.034811f
C70 VN.n24 VSUBS 0.041442f
C71 VN.n25 VSUBS 0.041442f
C72 VN.n26 VSUBS 0.041442f
C73 VN.n27 VSUBS 0.07685f
C74 VN.n28 VSUBS 0.042705f
C75 VN.n29 VSUBS 0.595995f
C76 VN.n30 VSUBS 0.078794f
C77 VN.n31 VSUBS 0.054634f
C78 VN.t1 VSUBS 1.15551f
C79 VN.n32 VSUBS 0.083238f
C80 VN.n33 VSUBS 0.041442f
C81 VN.n34 VSUBS 0.050293f
C82 VN.n35 VSUBS 0.041442f
C83 VN.t3 VSUBS 1.15551f
C84 VN.n36 VSUBS 0.460145f
C85 VN.n37 VSUBS 0.060242f
C86 VN.n38 VSUBS 0.438092f
C87 VN.t6 VSUBS 1.15551f
C88 VN.t4 VSUBS 1.53138f
C89 VN.n39 VSUBS 0.5666f
C90 VN.n40 VSUBS 0.595759f
C91 VN.n41 VSUBS 0.065468f
C92 VN.n42 VSUBS 0.07685f
C93 VN.n43 VSUBS 0.041442f
C94 VN.n44 VSUBS 0.041442f
C95 VN.n45 VSUBS 0.041442f
C96 VN.n46 VSUBS 0.060242f
C97 VN.n47 VSUBS 0.07685f
C98 VN.n48 VSUBS 0.065468f
C99 VN.n49 VSUBS 0.041442f
C100 VN.n50 VSUBS 0.041442f
C101 VN.n51 VSUBS 0.041442f
C102 VN.n52 VSUBS 0.07685f
C103 VN.n53 VSUBS 0.079286f
C104 VN.n54 VSUBS 0.034811f
C105 VN.n55 VSUBS 0.041442f
C106 VN.n56 VSUBS 0.041442f
C107 VN.n57 VSUBS 0.041442f
C108 VN.n58 VSUBS 0.07685f
C109 VN.n59 VSUBS 0.042705f
C110 VN.n60 VSUBS 0.595995f
C111 VN.n61 VSUBS 2.06304f
C112 B.n0 VSUBS 0.006858f
C113 B.n1 VSUBS 0.006858f
C114 B.n2 VSUBS 0.010846f
C115 B.n3 VSUBS 0.010846f
C116 B.n4 VSUBS 0.010846f
C117 B.n5 VSUBS 0.010846f
C118 B.n6 VSUBS 0.010846f
C119 B.n7 VSUBS 0.010846f
C120 B.n8 VSUBS 0.010846f
C121 B.n9 VSUBS 0.010846f
C122 B.n10 VSUBS 0.010846f
C123 B.n11 VSUBS 0.010846f
C124 B.n12 VSUBS 0.010846f
C125 B.n13 VSUBS 0.010846f
C126 B.n14 VSUBS 0.010846f
C127 B.n15 VSUBS 0.010846f
C128 B.n16 VSUBS 0.010846f
C129 B.n17 VSUBS 0.010846f
C130 B.n18 VSUBS 0.010846f
C131 B.n19 VSUBS 0.010846f
C132 B.n20 VSUBS 0.010846f
C133 B.n21 VSUBS 0.010846f
C134 B.n22 VSUBS 0.010846f
C135 B.n23 VSUBS 0.010846f
C136 B.n24 VSUBS 0.010846f
C137 B.n25 VSUBS 0.010846f
C138 B.n26 VSUBS 0.010846f
C139 B.n27 VSUBS 0.010846f
C140 B.n28 VSUBS 0.010846f
C141 B.n29 VSUBS 0.024005f
C142 B.n30 VSUBS 0.010846f
C143 B.n31 VSUBS 0.010846f
C144 B.n32 VSUBS 0.010846f
C145 B.n33 VSUBS 0.010846f
C146 B.n34 VSUBS 0.010846f
C147 B.n35 VSUBS 0.010846f
C148 B.n36 VSUBS 0.010846f
C149 B.n37 VSUBS 0.010846f
C150 B.n38 VSUBS 0.007496f
C151 B.n39 VSUBS 0.010846f
C152 B.t2 VSUBS 0.084654f
C153 B.t1 VSUBS 0.118326f
C154 B.t0 VSUBS 0.817399f
C155 B.n40 VSUBS 0.206428f
C156 B.n41 VSUBS 0.174883f
C157 B.n42 VSUBS 0.025129f
C158 B.n43 VSUBS 0.010846f
C159 B.n44 VSUBS 0.010846f
C160 B.n45 VSUBS 0.010846f
C161 B.n46 VSUBS 0.010846f
C162 B.t11 VSUBS 0.084655f
C163 B.t10 VSUBS 0.118327f
C164 B.t9 VSUBS 0.817399f
C165 B.n47 VSUBS 0.206427f
C166 B.n48 VSUBS 0.174882f
C167 B.n49 VSUBS 0.010846f
C168 B.n50 VSUBS 0.010846f
C169 B.n51 VSUBS 0.010846f
C170 B.n52 VSUBS 0.010846f
C171 B.n53 VSUBS 0.010846f
C172 B.n54 VSUBS 0.010846f
C173 B.n55 VSUBS 0.010846f
C174 B.n56 VSUBS 0.010846f
C175 B.n57 VSUBS 0.025312f
C176 B.n58 VSUBS 0.010846f
C177 B.n59 VSUBS 0.010846f
C178 B.n60 VSUBS 0.010846f
C179 B.n61 VSUBS 0.010846f
C180 B.n62 VSUBS 0.010846f
C181 B.n63 VSUBS 0.010846f
C182 B.n64 VSUBS 0.010846f
C183 B.n65 VSUBS 0.010846f
C184 B.n66 VSUBS 0.010846f
C185 B.n67 VSUBS 0.010846f
C186 B.n68 VSUBS 0.010846f
C187 B.n69 VSUBS 0.010846f
C188 B.n70 VSUBS 0.010846f
C189 B.n71 VSUBS 0.010846f
C190 B.n72 VSUBS 0.010846f
C191 B.n73 VSUBS 0.010846f
C192 B.n74 VSUBS 0.010846f
C193 B.n75 VSUBS 0.010846f
C194 B.n76 VSUBS 0.010846f
C195 B.n77 VSUBS 0.010846f
C196 B.n78 VSUBS 0.010846f
C197 B.n79 VSUBS 0.010846f
C198 B.n80 VSUBS 0.010846f
C199 B.n81 VSUBS 0.010846f
C200 B.n82 VSUBS 0.010846f
C201 B.n83 VSUBS 0.010846f
C202 B.n84 VSUBS 0.010846f
C203 B.n85 VSUBS 0.010846f
C204 B.n86 VSUBS 0.010846f
C205 B.n87 VSUBS 0.010846f
C206 B.n88 VSUBS 0.010846f
C207 B.n89 VSUBS 0.010846f
C208 B.n90 VSUBS 0.010846f
C209 B.n91 VSUBS 0.010846f
C210 B.n92 VSUBS 0.010846f
C211 B.n93 VSUBS 0.010846f
C212 B.n94 VSUBS 0.010846f
C213 B.n95 VSUBS 0.010846f
C214 B.n96 VSUBS 0.010846f
C215 B.n97 VSUBS 0.010846f
C216 B.n98 VSUBS 0.010846f
C217 B.n99 VSUBS 0.010846f
C218 B.n100 VSUBS 0.010846f
C219 B.n101 VSUBS 0.010846f
C220 B.n102 VSUBS 0.010846f
C221 B.n103 VSUBS 0.010846f
C222 B.n104 VSUBS 0.010846f
C223 B.n105 VSUBS 0.010846f
C224 B.n106 VSUBS 0.010846f
C225 B.n107 VSUBS 0.010846f
C226 B.n108 VSUBS 0.010846f
C227 B.n109 VSUBS 0.010846f
C228 B.n110 VSUBS 0.010846f
C229 B.n111 VSUBS 0.010846f
C230 B.n112 VSUBS 0.024005f
C231 B.n113 VSUBS 0.010846f
C232 B.n114 VSUBS 0.010846f
C233 B.n115 VSUBS 0.010846f
C234 B.n116 VSUBS 0.010846f
C235 B.n117 VSUBS 0.010846f
C236 B.n118 VSUBS 0.010846f
C237 B.n119 VSUBS 0.010846f
C238 B.n120 VSUBS 0.010846f
C239 B.n121 VSUBS 0.007496f
C240 B.n122 VSUBS 0.010846f
C241 B.n123 VSUBS 0.010846f
C242 B.n124 VSUBS 0.010846f
C243 B.n125 VSUBS 0.010846f
C244 B.n126 VSUBS 0.010846f
C245 B.t4 VSUBS 0.084654f
C246 B.t5 VSUBS 0.118326f
C247 B.t3 VSUBS 0.817399f
C248 B.n127 VSUBS 0.206428f
C249 B.n128 VSUBS 0.174883f
C250 B.n129 VSUBS 0.010846f
C251 B.n130 VSUBS 0.010846f
C252 B.n131 VSUBS 0.010846f
C253 B.n132 VSUBS 0.010846f
C254 B.n133 VSUBS 0.010846f
C255 B.n134 VSUBS 0.010846f
C256 B.n135 VSUBS 0.010846f
C257 B.n136 VSUBS 0.010846f
C258 B.n137 VSUBS 0.024005f
C259 B.n138 VSUBS 0.010846f
C260 B.n139 VSUBS 0.010846f
C261 B.n140 VSUBS 0.010846f
C262 B.n141 VSUBS 0.010846f
C263 B.n142 VSUBS 0.010846f
C264 B.n143 VSUBS 0.010846f
C265 B.n144 VSUBS 0.010846f
C266 B.n145 VSUBS 0.010846f
C267 B.n146 VSUBS 0.010846f
C268 B.n147 VSUBS 0.010846f
C269 B.n148 VSUBS 0.010846f
C270 B.n149 VSUBS 0.010846f
C271 B.n150 VSUBS 0.010846f
C272 B.n151 VSUBS 0.010846f
C273 B.n152 VSUBS 0.010846f
C274 B.n153 VSUBS 0.010846f
C275 B.n154 VSUBS 0.010846f
C276 B.n155 VSUBS 0.010846f
C277 B.n156 VSUBS 0.010846f
C278 B.n157 VSUBS 0.010846f
C279 B.n158 VSUBS 0.010846f
C280 B.n159 VSUBS 0.010846f
C281 B.n160 VSUBS 0.010846f
C282 B.n161 VSUBS 0.010846f
C283 B.n162 VSUBS 0.010846f
C284 B.n163 VSUBS 0.010846f
C285 B.n164 VSUBS 0.010846f
C286 B.n165 VSUBS 0.010846f
C287 B.n166 VSUBS 0.010846f
C288 B.n167 VSUBS 0.010846f
C289 B.n168 VSUBS 0.010846f
C290 B.n169 VSUBS 0.010846f
C291 B.n170 VSUBS 0.010846f
C292 B.n171 VSUBS 0.010846f
C293 B.n172 VSUBS 0.010846f
C294 B.n173 VSUBS 0.010846f
C295 B.n174 VSUBS 0.010846f
C296 B.n175 VSUBS 0.010846f
C297 B.n176 VSUBS 0.010846f
C298 B.n177 VSUBS 0.010846f
C299 B.n178 VSUBS 0.010846f
C300 B.n179 VSUBS 0.010846f
C301 B.n180 VSUBS 0.010846f
C302 B.n181 VSUBS 0.010846f
C303 B.n182 VSUBS 0.010846f
C304 B.n183 VSUBS 0.010846f
C305 B.n184 VSUBS 0.010846f
C306 B.n185 VSUBS 0.010846f
C307 B.n186 VSUBS 0.010846f
C308 B.n187 VSUBS 0.010846f
C309 B.n188 VSUBS 0.010846f
C310 B.n189 VSUBS 0.010846f
C311 B.n190 VSUBS 0.010846f
C312 B.n191 VSUBS 0.010846f
C313 B.n192 VSUBS 0.010846f
C314 B.n193 VSUBS 0.010846f
C315 B.n194 VSUBS 0.010846f
C316 B.n195 VSUBS 0.010846f
C317 B.n196 VSUBS 0.010846f
C318 B.n197 VSUBS 0.010846f
C319 B.n198 VSUBS 0.010846f
C320 B.n199 VSUBS 0.010846f
C321 B.n200 VSUBS 0.010846f
C322 B.n201 VSUBS 0.010846f
C323 B.n202 VSUBS 0.010846f
C324 B.n203 VSUBS 0.010846f
C325 B.n204 VSUBS 0.010846f
C326 B.n205 VSUBS 0.010846f
C327 B.n206 VSUBS 0.010846f
C328 B.n207 VSUBS 0.010846f
C329 B.n208 VSUBS 0.010846f
C330 B.n209 VSUBS 0.010846f
C331 B.n210 VSUBS 0.010846f
C332 B.n211 VSUBS 0.010846f
C333 B.n212 VSUBS 0.010846f
C334 B.n213 VSUBS 0.010846f
C335 B.n214 VSUBS 0.010846f
C336 B.n215 VSUBS 0.010846f
C337 B.n216 VSUBS 0.010846f
C338 B.n217 VSUBS 0.010846f
C339 B.n218 VSUBS 0.010846f
C340 B.n219 VSUBS 0.010846f
C341 B.n220 VSUBS 0.010846f
C342 B.n221 VSUBS 0.010846f
C343 B.n222 VSUBS 0.010846f
C344 B.n223 VSUBS 0.010846f
C345 B.n224 VSUBS 0.010846f
C346 B.n225 VSUBS 0.010846f
C347 B.n226 VSUBS 0.010846f
C348 B.n227 VSUBS 0.010846f
C349 B.n228 VSUBS 0.010846f
C350 B.n229 VSUBS 0.010846f
C351 B.n230 VSUBS 0.010846f
C352 B.n231 VSUBS 0.010846f
C353 B.n232 VSUBS 0.010846f
C354 B.n233 VSUBS 0.010846f
C355 B.n234 VSUBS 0.010846f
C356 B.n235 VSUBS 0.010846f
C357 B.n236 VSUBS 0.010846f
C358 B.n237 VSUBS 0.010846f
C359 B.n238 VSUBS 0.010846f
C360 B.n239 VSUBS 0.010846f
C361 B.n240 VSUBS 0.010846f
C362 B.n241 VSUBS 0.010846f
C363 B.n242 VSUBS 0.010846f
C364 B.n243 VSUBS 0.010846f
C365 B.n244 VSUBS 0.024005f
C366 B.n245 VSUBS 0.026078f
C367 B.n246 VSUBS 0.026078f
C368 B.n247 VSUBS 0.010846f
C369 B.n248 VSUBS 0.010846f
C370 B.n249 VSUBS 0.010846f
C371 B.n250 VSUBS 0.010846f
C372 B.n251 VSUBS 0.010846f
C373 B.n252 VSUBS 0.010846f
C374 B.n253 VSUBS 0.010846f
C375 B.n254 VSUBS 0.010846f
C376 B.n255 VSUBS 0.010846f
C377 B.n256 VSUBS 0.010846f
C378 B.n257 VSUBS 0.010846f
C379 B.n258 VSUBS 0.010846f
C380 B.n259 VSUBS 0.010846f
C381 B.n260 VSUBS 0.010846f
C382 B.n261 VSUBS 0.010846f
C383 B.n262 VSUBS 0.010846f
C384 B.n263 VSUBS 0.010846f
C385 B.n264 VSUBS 0.010846f
C386 B.n265 VSUBS 0.010846f
C387 B.n266 VSUBS 0.010846f
C388 B.n267 VSUBS 0.010846f
C389 B.n268 VSUBS 0.010846f
C390 B.n269 VSUBS 0.010846f
C391 B.n270 VSUBS 0.010846f
C392 B.n271 VSUBS 0.007496f
C393 B.n272 VSUBS 0.025129f
C394 B.n273 VSUBS 0.008772f
C395 B.n274 VSUBS 0.010846f
C396 B.n275 VSUBS 0.010846f
C397 B.n276 VSUBS 0.010846f
C398 B.n277 VSUBS 0.010846f
C399 B.n278 VSUBS 0.010846f
C400 B.n279 VSUBS 0.010846f
C401 B.n280 VSUBS 0.010846f
C402 B.n281 VSUBS 0.010846f
C403 B.n282 VSUBS 0.010846f
C404 B.n283 VSUBS 0.010846f
C405 B.n284 VSUBS 0.010846f
C406 B.t7 VSUBS 0.084655f
C407 B.t8 VSUBS 0.118327f
C408 B.t6 VSUBS 0.817399f
C409 B.n285 VSUBS 0.206427f
C410 B.n286 VSUBS 0.174882f
C411 B.n287 VSUBS 0.025129f
C412 B.n288 VSUBS 0.008772f
C413 B.n289 VSUBS 0.010846f
C414 B.n290 VSUBS 0.010846f
C415 B.n291 VSUBS 0.010846f
C416 B.n292 VSUBS 0.010846f
C417 B.n293 VSUBS 0.010846f
C418 B.n294 VSUBS 0.010846f
C419 B.n295 VSUBS 0.010846f
C420 B.n296 VSUBS 0.010846f
C421 B.n297 VSUBS 0.010846f
C422 B.n298 VSUBS 0.010846f
C423 B.n299 VSUBS 0.010846f
C424 B.n300 VSUBS 0.010846f
C425 B.n301 VSUBS 0.010846f
C426 B.n302 VSUBS 0.010846f
C427 B.n303 VSUBS 0.010846f
C428 B.n304 VSUBS 0.010846f
C429 B.n305 VSUBS 0.010846f
C430 B.n306 VSUBS 0.010846f
C431 B.n307 VSUBS 0.010846f
C432 B.n308 VSUBS 0.010846f
C433 B.n309 VSUBS 0.010846f
C434 B.n310 VSUBS 0.010846f
C435 B.n311 VSUBS 0.010846f
C436 B.n312 VSUBS 0.010846f
C437 B.n313 VSUBS 0.010846f
C438 B.n314 VSUBS 0.010846f
C439 B.n315 VSUBS 0.026078f
C440 B.n316 VSUBS 0.026078f
C441 B.n317 VSUBS 0.024005f
C442 B.n318 VSUBS 0.010846f
C443 B.n319 VSUBS 0.010846f
C444 B.n320 VSUBS 0.010846f
C445 B.n321 VSUBS 0.010846f
C446 B.n322 VSUBS 0.010846f
C447 B.n323 VSUBS 0.010846f
C448 B.n324 VSUBS 0.010846f
C449 B.n325 VSUBS 0.010846f
C450 B.n326 VSUBS 0.010846f
C451 B.n327 VSUBS 0.010846f
C452 B.n328 VSUBS 0.010846f
C453 B.n329 VSUBS 0.010846f
C454 B.n330 VSUBS 0.010846f
C455 B.n331 VSUBS 0.010846f
C456 B.n332 VSUBS 0.010846f
C457 B.n333 VSUBS 0.010846f
C458 B.n334 VSUBS 0.010846f
C459 B.n335 VSUBS 0.010846f
C460 B.n336 VSUBS 0.010846f
C461 B.n337 VSUBS 0.010846f
C462 B.n338 VSUBS 0.010846f
C463 B.n339 VSUBS 0.010846f
C464 B.n340 VSUBS 0.010846f
C465 B.n341 VSUBS 0.010846f
C466 B.n342 VSUBS 0.010846f
C467 B.n343 VSUBS 0.010846f
C468 B.n344 VSUBS 0.010846f
C469 B.n345 VSUBS 0.010846f
C470 B.n346 VSUBS 0.010846f
C471 B.n347 VSUBS 0.010846f
C472 B.n348 VSUBS 0.010846f
C473 B.n349 VSUBS 0.010846f
C474 B.n350 VSUBS 0.010846f
C475 B.n351 VSUBS 0.010846f
C476 B.n352 VSUBS 0.010846f
C477 B.n353 VSUBS 0.010846f
C478 B.n354 VSUBS 0.010846f
C479 B.n355 VSUBS 0.010846f
C480 B.n356 VSUBS 0.010846f
C481 B.n357 VSUBS 0.010846f
C482 B.n358 VSUBS 0.010846f
C483 B.n359 VSUBS 0.010846f
C484 B.n360 VSUBS 0.010846f
C485 B.n361 VSUBS 0.010846f
C486 B.n362 VSUBS 0.010846f
C487 B.n363 VSUBS 0.010846f
C488 B.n364 VSUBS 0.010846f
C489 B.n365 VSUBS 0.010846f
C490 B.n366 VSUBS 0.010846f
C491 B.n367 VSUBS 0.010846f
C492 B.n368 VSUBS 0.010846f
C493 B.n369 VSUBS 0.010846f
C494 B.n370 VSUBS 0.010846f
C495 B.n371 VSUBS 0.010846f
C496 B.n372 VSUBS 0.010846f
C497 B.n373 VSUBS 0.010846f
C498 B.n374 VSUBS 0.010846f
C499 B.n375 VSUBS 0.010846f
C500 B.n376 VSUBS 0.010846f
C501 B.n377 VSUBS 0.010846f
C502 B.n378 VSUBS 0.010846f
C503 B.n379 VSUBS 0.010846f
C504 B.n380 VSUBS 0.010846f
C505 B.n381 VSUBS 0.010846f
C506 B.n382 VSUBS 0.010846f
C507 B.n383 VSUBS 0.010846f
C508 B.n384 VSUBS 0.010846f
C509 B.n385 VSUBS 0.010846f
C510 B.n386 VSUBS 0.010846f
C511 B.n387 VSUBS 0.010846f
C512 B.n388 VSUBS 0.010846f
C513 B.n389 VSUBS 0.010846f
C514 B.n390 VSUBS 0.010846f
C515 B.n391 VSUBS 0.010846f
C516 B.n392 VSUBS 0.010846f
C517 B.n393 VSUBS 0.010846f
C518 B.n394 VSUBS 0.010846f
C519 B.n395 VSUBS 0.010846f
C520 B.n396 VSUBS 0.010846f
C521 B.n397 VSUBS 0.010846f
C522 B.n398 VSUBS 0.010846f
C523 B.n399 VSUBS 0.010846f
C524 B.n400 VSUBS 0.010846f
C525 B.n401 VSUBS 0.010846f
C526 B.n402 VSUBS 0.010846f
C527 B.n403 VSUBS 0.010846f
C528 B.n404 VSUBS 0.010846f
C529 B.n405 VSUBS 0.010846f
C530 B.n406 VSUBS 0.010846f
C531 B.n407 VSUBS 0.010846f
C532 B.n408 VSUBS 0.010846f
C533 B.n409 VSUBS 0.010846f
C534 B.n410 VSUBS 0.010846f
C535 B.n411 VSUBS 0.010846f
C536 B.n412 VSUBS 0.010846f
C537 B.n413 VSUBS 0.010846f
C538 B.n414 VSUBS 0.010846f
C539 B.n415 VSUBS 0.010846f
C540 B.n416 VSUBS 0.010846f
C541 B.n417 VSUBS 0.010846f
C542 B.n418 VSUBS 0.010846f
C543 B.n419 VSUBS 0.010846f
C544 B.n420 VSUBS 0.010846f
C545 B.n421 VSUBS 0.010846f
C546 B.n422 VSUBS 0.010846f
C547 B.n423 VSUBS 0.010846f
C548 B.n424 VSUBS 0.010846f
C549 B.n425 VSUBS 0.010846f
C550 B.n426 VSUBS 0.010846f
C551 B.n427 VSUBS 0.010846f
C552 B.n428 VSUBS 0.010846f
C553 B.n429 VSUBS 0.010846f
C554 B.n430 VSUBS 0.010846f
C555 B.n431 VSUBS 0.010846f
C556 B.n432 VSUBS 0.010846f
C557 B.n433 VSUBS 0.010846f
C558 B.n434 VSUBS 0.010846f
C559 B.n435 VSUBS 0.010846f
C560 B.n436 VSUBS 0.010846f
C561 B.n437 VSUBS 0.010846f
C562 B.n438 VSUBS 0.010846f
C563 B.n439 VSUBS 0.010846f
C564 B.n440 VSUBS 0.010846f
C565 B.n441 VSUBS 0.010846f
C566 B.n442 VSUBS 0.010846f
C567 B.n443 VSUBS 0.010846f
C568 B.n444 VSUBS 0.010846f
C569 B.n445 VSUBS 0.010846f
C570 B.n446 VSUBS 0.010846f
C571 B.n447 VSUBS 0.010846f
C572 B.n448 VSUBS 0.010846f
C573 B.n449 VSUBS 0.010846f
C574 B.n450 VSUBS 0.010846f
C575 B.n451 VSUBS 0.010846f
C576 B.n452 VSUBS 0.010846f
C577 B.n453 VSUBS 0.010846f
C578 B.n454 VSUBS 0.010846f
C579 B.n455 VSUBS 0.010846f
C580 B.n456 VSUBS 0.010846f
C581 B.n457 VSUBS 0.010846f
C582 B.n458 VSUBS 0.010846f
C583 B.n459 VSUBS 0.010846f
C584 B.n460 VSUBS 0.010846f
C585 B.n461 VSUBS 0.010846f
C586 B.n462 VSUBS 0.010846f
C587 B.n463 VSUBS 0.010846f
C588 B.n464 VSUBS 0.010846f
C589 B.n465 VSUBS 0.010846f
C590 B.n466 VSUBS 0.010846f
C591 B.n467 VSUBS 0.010846f
C592 B.n468 VSUBS 0.010846f
C593 B.n469 VSUBS 0.010846f
C594 B.n470 VSUBS 0.010846f
C595 B.n471 VSUBS 0.010846f
C596 B.n472 VSUBS 0.010846f
C597 B.n473 VSUBS 0.010846f
C598 B.n474 VSUBS 0.010846f
C599 B.n475 VSUBS 0.010846f
C600 B.n476 VSUBS 0.010846f
C601 B.n477 VSUBS 0.010846f
C602 B.n478 VSUBS 0.010846f
C603 B.n479 VSUBS 0.010846f
C604 B.n480 VSUBS 0.010846f
C605 B.n481 VSUBS 0.010846f
C606 B.n482 VSUBS 0.024005f
C607 B.n483 VSUBS 0.026078f
C608 B.n484 VSUBS 0.02477f
C609 B.n485 VSUBS 0.010846f
C610 B.n486 VSUBS 0.010846f
C611 B.n487 VSUBS 0.010846f
C612 B.n488 VSUBS 0.010846f
C613 B.n489 VSUBS 0.010846f
C614 B.n490 VSUBS 0.010846f
C615 B.n491 VSUBS 0.010846f
C616 B.n492 VSUBS 0.010846f
C617 B.n493 VSUBS 0.010846f
C618 B.n494 VSUBS 0.010846f
C619 B.n495 VSUBS 0.010846f
C620 B.n496 VSUBS 0.010846f
C621 B.n497 VSUBS 0.010846f
C622 B.n498 VSUBS 0.010846f
C623 B.n499 VSUBS 0.010846f
C624 B.n500 VSUBS 0.010846f
C625 B.n501 VSUBS 0.010846f
C626 B.n502 VSUBS 0.010846f
C627 B.n503 VSUBS 0.010846f
C628 B.n504 VSUBS 0.010846f
C629 B.n505 VSUBS 0.010846f
C630 B.n506 VSUBS 0.010846f
C631 B.n507 VSUBS 0.010846f
C632 B.n508 VSUBS 0.010846f
C633 B.n509 VSUBS 0.007496f
C634 B.n510 VSUBS 0.025129f
C635 B.n511 VSUBS 0.008772f
C636 B.n512 VSUBS 0.010846f
C637 B.n513 VSUBS 0.010846f
C638 B.n514 VSUBS 0.010846f
C639 B.n515 VSUBS 0.010846f
C640 B.n516 VSUBS 0.010846f
C641 B.n517 VSUBS 0.010846f
C642 B.n518 VSUBS 0.010846f
C643 B.n519 VSUBS 0.010846f
C644 B.n520 VSUBS 0.010846f
C645 B.n521 VSUBS 0.010846f
C646 B.n522 VSUBS 0.010846f
C647 B.n523 VSUBS 0.008772f
C648 B.n524 VSUBS 0.010846f
C649 B.n525 VSUBS 0.010846f
C650 B.n526 VSUBS 0.010846f
C651 B.n527 VSUBS 0.010846f
C652 B.n528 VSUBS 0.010846f
C653 B.n529 VSUBS 0.010846f
C654 B.n530 VSUBS 0.010846f
C655 B.n531 VSUBS 0.010846f
C656 B.n532 VSUBS 0.010846f
C657 B.n533 VSUBS 0.010846f
C658 B.n534 VSUBS 0.010846f
C659 B.n535 VSUBS 0.010846f
C660 B.n536 VSUBS 0.010846f
C661 B.n537 VSUBS 0.010846f
C662 B.n538 VSUBS 0.010846f
C663 B.n539 VSUBS 0.010846f
C664 B.n540 VSUBS 0.010846f
C665 B.n541 VSUBS 0.010846f
C666 B.n542 VSUBS 0.010846f
C667 B.n543 VSUBS 0.010846f
C668 B.n544 VSUBS 0.010846f
C669 B.n545 VSUBS 0.010846f
C670 B.n546 VSUBS 0.010846f
C671 B.n547 VSUBS 0.010846f
C672 B.n548 VSUBS 0.010846f
C673 B.n549 VSUBS 0.010846f
C674 B.n550 VSUBS 0.026078f
C675 B.n551 VSUBS 0.026078f
C676 B.n552 VSUBS 0.024005f
C677 B.n553 VSUBS 0.010846f
C678 B.n554 VSUBS 0.010846f
C679 B.n555 VSUBS 0.010846f
C680 B.n556 VSUBS 0.010846f
C681 B.n557 VSUBS 0.010846f
C682 B.n558 VSUBS 0.010846f
C683 B.n559 VSUBS 0.010846f
C684 B.n560 VSUBS 0.010846f
C685 B.n561 VSUBS 0.010846f
C686 B.n562 VSUBS 0.010846f
C687 B.n563 VSUBS 0.010846f
C688 B.n564 VSUBS 0.010846f
C689 B.n565 VSUBS 0.010846f
C690 B.n566 VSUBS 0.010846f
C691 B.n567 VSUBS 0.010846f
C692 B.n568 VSUBS 0.010846f
C693 B.n569 VSUBS 0.010846f
C694 B.n570 VSUBS 0.010846f
C695 B.n571 VSUBS 0.010846f
C696 B.n572 VSUBS 0.010846f
C697 B.n573 VSUBS 0.010846f
C698 B.n574 VSUBS 0.010846f
C699 B.n575 VSUBS 0.010846f
C700 B.n576 VSUBS 0.010846f
C701 B.n577 VSUBS 0.010846f
C702 B.n578 VSUBS 0.010846f
C703 B.n579 VSUBS 0.010846f
C704 B.n580 VSUBS 0.010846f
C705 B.n581 VSUBS 0.010846f
C706 B.n582 VSUBS 0.010846f
C707 B.n583 VSUBS 0.010846f
C708 B.n584 VSUBS 0.010846f
C709 B.n585 VSUBS 0.010846f
C710 B.n586 VSUBS 0.010846f
C711 B.n587 VSUBS 0.010846f
C712 B.n588 VSUBS 0.010846f
C713 B.n589 VSUBS 0.010846f
C714 B.n590 VSUBS 0.010846f
C715 B.n591 VSUBS 0.010846f
C716 B.n592 VSUBS 0.010846f
C717 B.n593 VSUBS 0.010846f
C718 B.n594 VSUBS 0.010846f
C719 B.n595 VSUBS 0.010846f
C720 B.n596 VSUBS 0.010846f
C721 B.n597 VSUBS 0.010846f
C722 B.n598 VSUBS 0.010846f
C723 B.n599 VSUBS 0.010846f
C724 B.n600 VSUBS 0.010846f
C725 B.n601 VSUBS 0.010846f
C726 B.n602 VSUBS 0.010846f
C727 B.n603 VSUBS 0.010846f
C728 B.n604 VSUBS 0.010846f
C729 B.n605 VSUBS 0.010846f
C730 B.n606 VSUBS 0.010846f
C731 B.n607 VSUBS 0.010846f
C732 B.n608 VSUBS 0.010846f
C733 B.n609 VSUBS 0.010846f
C734 B.n610 VSUBS 0.010846f
C735 B.n611 VSUBS 0.010846f
C736 B.n612 VSUBS 0.010846f
C737 B.n613 VSUBS 0.010846f
C738 B.n614 VSUBS 0.010846f
C739 B.n615 VSUBS 0.010846f
C740 B.n616 VSUBS 0.010846f
C741 B.n617 VSUBS 0.010846f
C742 B.n618 VSUBS 0.010846f
C743 B.n619 VSUBS 0.010846f
C744 B.n620 VSUBS 0.010846f
C745 B.n621 VSUBS 0.010846f
C746 B.n622 VSUBS 0.010846f
C747 B.n623 VSUBS 0.010846f
C748 B.n624 VSUBS 0.010846f
C749 B.n625 VSUBS 0.010846f
C750 B.n626 VSUBS 0.010846f
C751 B.n627 VSUBS 0.010846f
C752 B.n628 VSUBS 0.010846f
C753 B.n629 VSUBS 0.010846f
C754 B.n630 VSUBS 0.010846f
C755 B.n631 VSUBS 0.010846f
C756 B.n632 VSUBS 0.010846f
C757 B.n633 VSUBS 0.010846f
C758 B.n634 VSUBS 0.010846f
C759 B.n635 VSUBS 0.024559f
C760 VTAIL.t1 VSUBS 0.099954f
C761 VTAIL.t4 VSUBS 0.099954f
C762 VTAIL.n0 VSUBS 0.495079f
C763 VTAIL.n1 VSUBS 0.797574f
C764 VTAIL.n2 VSUBS 0.034178f
C765 VTAIL.n3 VSUBS 0.033286f
C766 VTAIL.n4 VSUBS 0.017886f
C767 VTAIL.n5 VSUBS 0.042277f
C768 VTAIL.n6 VSUBS 0.018939f
C769 VTAIL.n7 VSUBS 0.126308f
C770 VTAIL.t7 VSUBS 0.092224f
C771 VTAIL.n8 VSUBS 0.031708f
C772 VTAIL.n9 VSUBS 0.026592f
C773 VTAIL.n10 VSUBS 0.017886f
C774 VTAIL.n11 VSUBS 0.428985f
C775 VTAIL.n12 VSUBS 0.033286f
C776 VTAIL.n13 VSUBS 0.017886f
C777 VTAIL.n14 VSUBS 0.018939f
C778 VTAIL.n15 VSUBS 0.042277f
C779 VTAIL.n16 VSUBS 0.094185f
C780 VTAIL.n17 VSUBS 0.018939f
C781 VTAIL.n18 VSUBS 0.017886f
C782 VTAIL.n19 VSUBS 0.075121f
C783 VTAIL.n20 VSUBS 0.046946f
C784 VTAIL.n21 VSUBS 0.373671f
C785 VTAIL.n22 VSUBS 0.034178f
C786 VTAIL.n23 VSUBS 0.033286f
C787 VTAIL.n24 VSUBS 0.017886f
C788 VTAIL.n25 VSUBS 0.042277f
C789 VTAIL.n26 VSUBS 0.018939f
C790 VTAIL.n27 VSUBS 0.126308f
C791 VTAIL.t9 VSUBS 0.092224f
C792 VTAIL.n28 VSUBS 0.031708f
C793 VTAIL.n29 VSUBS 0.026592f
C794 VTAIL.n30 VSUBS 0.017886f
C795 VTAIL.n31 VSUBS 0.428985f
C796 VTAIL.n32 VSUBS 0.033286f
C797 VTAIL.n33 VSUBS 0.017886f
C798 VTAIL.n34 VSUBS 0.018939f
C799 VTAIL.n35 VSUBS 0.042277f
C800 VTAIL.n36 VSUBS 0.094185f
C801 VTAIL.n37 VSUBS 0.018939f
C802 VTAIL.n38 VSUBS 0.017886f
C803 VTAIL.n39 VSUBS 0.075121f
C804 VTAIL.n40 VSUBS 0.046946f
C805 VTAIL.n41 VSUBS 0.373671f
C806 VTAIL.t8 VSUBS 0.099954f
C807 VTAIL.t13 VSUBS 0.099954f
C808 VTAIL.n42 VSUBS 0.495079f
C809 VTAIL.n43 VSUBS 1.08721f
C810 VTAIL.n44 VSUBS 0.034178f
C811 VTAIL.n45 VSUBS 0.033286f
C812 VTAIL.n46 VSUBS 0.017886f
C813 VTAIL.n47 VSUBS 0.042277f
C814 VTAIL.n48 VSUBS 0.018939f
C815 VTAIL.n49 VSUBS 0.126308f
C816 VTAIL.t12 VSUBS 0.092224f
C817 VTAIL.n50 VSUBS 0.031708f
C818 VTAIL.n51 VSUBS 0.026592f
C819 VTAIL.n52 VSUBS 0.017886f
C820 VTAIL.n53 VSUBS 0.428985f
C821 VTAIL.n54 VSUBS 0.033286f
C822 VTAIL.n55 VSUBS 0.017886f
C823 VTAIL.n56 VSUBS 0.018939f
C824 VTAIL.n57 VSUBS 0.042277f
C825 VTAIL.n58 VSUBS 0.094185f
C826 VTAIL.n59 VSUBS 0.018939f
C827 VTAIL.n60 VSUBS 0.017886f
C828 VTAIL.n61 VSUBS 0.075121f
C829 VTAIL.n62 VSUBS 0.046946f
C830 VTAIL.n63 VSUBS 1.42266f
C831 VTAIL.n64 VSUBS 0.034178f
C832 VTAIL.n65 VSUBS 0.033286f
C833 VTAIL.n66 VSUBS 0.017886f
C834 VTAIL.n67 VSUBS 0.042277f
C835 VTAIL.n68 VSUBS 0.018939f
C836 VTAIL.n69 VSUBS 0.126308f
C837 VTAIL.t5 VSUBS 0.092224f
C838 VTAIL.n70 VSUBS 0.031708f
C839 VTAIL.n71 VSUBS 0.026592f
C840 VTAIL.n72 VSUBS 0.017886f
C841 VTAIL.n73 VSUBS 0.428985f
C842 VTAIL.n74 VSUBS 0.033286f
C843 VTAIL.n75 VSUBS 0.017886f
C844 VTAIL.n76 VSUBS 0.018939f
C845 VTAIL.n77 VSUBS 0.042277f
C846 VTAIL.n78 VSUBS 0.094185f
C847 VTAIL.n79 VSUBS 0.018939f
C848 VTAIL.n80 VSUBS 0.017886f
C849 VTAIL.n81 VSUBS 0.075121f
C850 VTAIL.n82 VSUBS 0.046946f
C851 VTAIL.n83 VSUBS 1.42266f
C852 VTAIL.t6 VSUBS 0.099954f
C853 VTAIL.t2 VSUBS 0.099954f
C854 VTAIL.n84 VSUBS 0.495082f
C855 VTAIL.n85 VSUBS 1.08721f
C856 VTAIL.n86 VSUBS 0.034178f
C857 VTAIL.n87 VSUBS 0.033286f
C858 VTAIL.n88 VSUBS 0.017886f
C859 VTAIL.n89 VSUBS 0.042277f
C860 VTAIL.n90 VSUBS 0.018939f
C861 VTAIL.n91 VSUBS 0.126308f
C862 VTAIL.t3 VSUBS 0.092224f
C863 VTAIL.n92 VSUBS 0.031708f
C864 VTAIL.n93 VSUBS 0.026592f
C865 VTAIL.n94 VSUBS 0.017886f
C866 VTAIL.n95 VSUBS 0.428985f
C867 VTAIL.n96 VSUBS 0.033286f
C868 VTAIL.n97 VSUBS 0.017886f
C869 VTAIL.n98 VSUBS 0.018939f
C870 VTAIL.n99 VSUBS 0.042277f
C871 VTAIL.n100 VSUBS 0.094185f
C872 VTAIL.n101 VSUBS 0.018939f
C873 VTAIL.n102 VSUBS 0.017886f
C874 VTAIL.n103 VSUBS 0.075121f
C875 VTAIL.n104 VSUBS 0.046946f
C876 VTAIL.n105 VSUBS 0.373671f
C877 VTAIL.n106 VSUBS 0.034178f
C878 VTAIL.n107 VSUBS 0.033286f
C879 VTAIL.n108 VSUBS 0.017886f
C880 VTAIL.n109 VSUBS 0.042277f
C881 VTAIL.n110 VSUBS 0.018939f
C882 VTAIL.n111 VSUBS 0.126308f
C883 VTAIL.t15 VSUBS 0.092224f
C884 VTAIL.n112 VSUBS 0.031708f
C885 VTAIL.n113 VSUBS 0.026592f
C886 VTAIL.n114 VSUBS 0.017886f
C887 VTAIL.n115 VSUBS 0.428985f
C888 VTAIL.n116 VSUBS 0.033286f
C889 VTAIL.n117 VSUBS 0.017886f
C890 VTAIL.n118 VSUBS 0.018939f
C891 VTAIL.n119 VSUBS 0.042277f
C892 VTAIL.n120 VSUBS 0.094185f
C893 VTAIL.n121 VSUBS 0.018939f
C894 VTAIL.n122 VSUBS 0.017886f
C895 VTAIL.n123 VSUBS 0.075121f
C896 VTAIL.n124 VSUBS 0.046946f
C897 VTAIL.n125 VSUBS 0.373671f
C898 VTAIL.t14 VSUBS 0.099954f
C899 VTAIL.t11 VSUBS 0.099954f
C900 VTAIL.n126 VSUBS 0.495082f
C901 VTAIL.n127 VSUBS 1.08721f
C902 VTAIL.n128 VSUBS 0.034178f
C903 VTAIL.n129 VSUBS 0.033286f
C904 VTAIL.n130 VSUBS 0.017886f
C905 VTAIL.n131 VSUBS 0.042277f
C906 VTAIL.n132 VSUBS 0.018939f
C907 VTAIL.n133 VSUBS 0.126308f
C908 VTAIL.t10 VSUBS 0.092224f
C909 VTAIL.n134 VSUBS 0.031708f
C910 VTAIL.n135 VSUBS 0.026592f
C911 VTAIL.n136 VSUBS 0.017886f
C912 VTAIL.n137 VSUBS 0.428985f
C913 VTAIL.n138 VSUBS 0.033286f
C914 VTAIL.n139 VSUBS 0.017886f
C915 VTAIL.n140 VSUBS 0.018939f
C916 VTAIL.n141 VSUBS 0.042277f
C917 VTAIL.n142 VSUBS 0.094185f
C918 VTAIL.n143 VSUBS 0.018939f
C919 VTAIL.n144 VSUBS 0.017886f
C920 VTAIL.n145 VSUBS 0.075121f
C921 VTAIL.n146 VSUBS 0.046946f
C922 VTAIL.n147 VSUBS 1.42266f
C923 VTAIL.n148 VSUBS 0.034178f
C924 VTAIL.n149 VSUBS 0.033286f
C925 VTAIL.n150 VSUBS 0.017886f
C926 VTAIL.n151 VSUBS 0.042277f
C927 VTAIL.n152 VSUBS 0.018939f
C928 VTAIL.n153 VSUBS 0.126308f
C929 VTAIL.t0 VSUBS 0.092224f
C930 VTAIL.n154 VSUBS 0.031708f
C931 VTAIL.n155 VSUBS 0.026592f
C932 VTAIL.n156 VSUBS 0.017886f
C933 VTAIL.n157 VSUBS 0.428985f
C934 VTAIL.n158 VSUBS 0.033286f
C935 VTAIL.n159 VSUBS 0.017886f
C936 VTAIL.n160 VSUBS 0.018939f
C937 VTAIL.n161 VSUBS 0.042277f
C938 VTAIL.n162 VSUBS 0.094185f
C939 VTAIL.n163 VSUBS 0.018939f
C940 VTAIL.n164 VSUBS 0.017886f
C941 VTAIL.n165 VSUBS 0.075121f
C942 VTAIL.n166 VSUBS 0.046946f
C943 VTAIL.n167 VSUBS 1.41642f
C944 VDD1.t7 VSUBS 0.074166f
C945 VDD1.t1 VSUBS 0.074166f
C946 VDD1.n0 VSUBS 0.434618f
C947 VDD1.t3 VSUBS 0.074166f
C948 VDD1.t6 VSUBS 0.074166f
C949 VDD1.n1 VSUBS 0.433842f
C950 VDD1.t2 VSUBS 0.074166f
C951 VDD1.t5 VSUBS 0.074166f
C952 VDD1.n2 VSUBS 0.433842f
C953 VDD1.n3 VSUBS 3.23151f
C954 VDD1.t0 VSUBS 0.074166f
C955 VDD1.t4 VSUBS 0.074166f
C956 VDD1.n4 VSUBS 0.425977f
C957 VDD1.n5 VSUBS 2.54953f
C958 VP.n0 VSUBS 0.062427f
C959 VP.t6 VSUBS 1.32033f
C960 VP.n1 VSUBS 0.09511f
C961 VP.n2 VSUBS 0.047353f
C962 VP.n3 VSUBS 0.057466f
C963 VP.n4 VSUBS 0.047353f
C964 VP.n5 VSUBS 0.068835f
C965 VP.n6 VSUBS 0.047353f
C966 VP.t7 VSUBS 1.32033f
C967 VP.n7 VSUBS 0.087812f
C968 VP.n8 VSUBS 0.047353f
C969 VP.n9 VSUBS 0.087812f
C970 VP.n10 VSUBS 0.062427f
C971 VP.t5 VSUBS 1.32033f
C972 VP.n11 VSUBS 0.09511f
C973 VP.n12 VSUBS 0.047353f
C974 VP.n13 VSUBS 0.057466f
C975 VP.n14 VSUBS 0.047353f
C976 VP.n15 VSUBS 0.068835f
C977 VP.n16 VSUBS 0.500581f
C978 VP.t1 VSUBS 1.32033f
C979 VP.t0 VSUBS 1.74981f
C980 VP.n17 VSUBS 0.647419f
C981 VP.n18 VSUBS 0.680736f
C982 VP.n19 VSUBS 0.074807f
C983 VP.n20 VSUBS 0.087812f
C984 VP.n21 VSUBS 0.047353f
C985 VP.n22 VSUBS 0.047353f
C986 VP.n23 VSUBS 0.047353f
C987 VP.n24 VSUBS 0.068835f
C988 VP.n25 VSUBS 0.087812f
C989 VP.t4 VSUBS 1.32033f
C990 VP.n26 VSUBS 0.525779f
C991 VP.n27 VSUBS 0.074807f
C992 VP.n28 VSUBS 0.047353f
C993 VP.n29 VSUBS 0.047353f
C994 VP.n30 VSUBS 0.047353f
C995 VP.n31 VSUBS 0.087812f
C996 VP.n32 VSUBS 0.090595f
C997 VP.n33 VSUBS 0.039776f
C998 VP.n34 VSUBS 0.047353f
C999 VP.n35 VSUBS 0.047353f
C1000 VP.n36 VSUBS 0.047353f
C1001 VP.n37 VSUBS 0.087812f
C1002 VP.n38 VSUBS 0.048797f
C1003 VP.n39 VSUBS 0.681007f
C1004 VP.n40 VSUBS 2.3315f
C1005 VP.n41 VSUBS 2.36868f
C1006 VP.t3 VSUBS 1.32033f
C1007 VP.n42 VSUBS 0.681007f
C1008 VP.n43 VSUBS 0.048797f
C1009 VP.n44 VSUBS 0.062427f
C1010 VP.n45 VSUBS 0.047353f
C1011 VP.n46 VSUBS 0.047353f
C1012 VP.n47 VSUBS 0.09511f
C1013 VP.n48 VSUBS 0.039776f
C1014 VP.n49 VSUBS 0.090595f
C1015 VP.n50 VSUBS 0.047353f
C1016 VP.n51 VSUBS 0.047353f
C1017 VP.n52 VSUBS 0.047353f
C1018 VP.n53 VSUBS 0.057466f
C1019 VP.n54 VSUBS 0.525779f
C1020 VP.n55 VSUBS 0.074807f
C1021 VP.n56 VSUBS 0.087812f
C1022 VP.n57 VSUBS 0.047353f
C1023 VP.n58 VSUBS 0.047353f
C1024 VP.n59 VSUBS 0.047353f
C1025 VP.n60 VSUBS 0.068835f
C1026 VP.n61 VSUBS 0.087812f
C1027 VP.t2 VSUBS 1.32033f
C1028 VP.n62 VSUBS 0.525779f
C1029 VP.n63 VSUBS 0.074807f
C1030 VP.n64 VSUBS 0.047353f
C1031 VP.n65 VSUBS 0.047353f
C1032 VP.n66 VSUBS 0.047353f
C1033 VP.n67 VSUBS 0.087812f
C1034 VP.n68 VSUBS 0.090595f
C1035 VP.n69 VSUBS 0.039776f
C1036 VP.n70 VSUBS 0.047353f
C1037 VP.n71 VSUBS 0.047353f
C1038 VP.n72 VSUBS 0.047353f
C1039 VP.n73 VSUBS 0.087812f
C1040 VP.n74 VSUBS 0.048797f
C1041 VP.n75 VSUBS 0.681007f
C1042 VP.n76 VSUBS 0.090033f
.ends

