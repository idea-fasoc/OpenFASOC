* NGSPICE file created from diff_pair_sample_0406.ext - technology: sky130A

.subckt diff_pair_sample_0406 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=3.10365 ps=19.14 w=18.81 l=1.55
X1 VTAIL.t10 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=3.10365 ps=19.14 w=18.81 l=1.55
X2 VDD1.t1 VP.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=3.10365 ps=19.14 w=18.81 l=1.55
X3 VDD2.t5 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=7.3359 ps=38.4 w=18.81 l=1.55
X4 VTAIL.t3 VN.t1 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=3.10365 ps=19.14 w=18.81 l=1.55
X5 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=3.10365 ps=19.14 w=18.81 l=1.55
X6 VDD1.t0 VP.t3 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=3.10365 ps=19.14 w=18.81 l=1.55
X7 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=0 ps=0 w=18.81 l=1.55
X8 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=0 ps=0 w=18.81 l=1.55
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=0 ps=0 w=18.81 l=1.55
X10 VDD1.t5 VP.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=7.3359 ps=38.4 w=18.81 l=1.55
X11 VDD1.t4 VP.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=7.3359 ps=38.4 w=18.81 l=1.55
X12 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=3.10365 ps=19.14 w=18.81 l=1.55
X13 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=7.3359 ps=38.4 w=18.81 l=1.55
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3359 pd=38.4 as=0 ps=0 w=18.81 l=1.55
X15 VTAIL.t4 VN.t5 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=3.10365 pd=19.14 as=3.10365 ps=19.14 w=18.81 l=1.55
R0 VP.n6 VP.t3 324.25
R1 VP.n17 VP.t2 292.466
R2 VP.n24 VP.t1 292.466
R3 VP.n31 VP.t5 292.466
R4 VP.n14 VP.t4 292.466
R5 VP.n7 VP.t0 292.466
R6 VP.n17 VP.n16 179.406
R7 VP.n32 VP.n31 179.406
R8 VP.n15 VP.n14 179.406
R9 VP.n9 VP.n8 161.3
R10 VP.n10 VP.n5 161.3
R11 VP.n12 VP.n11 161.3
R12 VP.n13 VP.n4 161.3
R13 VP.n30 VP.n0 161.3
R14 VP.n29 VP.n28 161.3
R15 VP.n27 VP.n1 161.3
R16 VP.n26 VP.n25 161.3
R17 VP.n23 VP.n2 161.3
R18 VP.n22 VP.n21 161.3
R19 VP.n20 VP.n3 161.3
R20 VP.n19 VP.n18 161.3
R21 VP.n22 VP.n3 56.5193
R22 VP.n29 VP.n1 56.5193
R23 VP.n12 VP.n5 56.5193
R24 VP.n7 VP.n6 53.7793
R25 VP.n16 VP.n15 49.599
R26 VP.n18 VP.n3 24.4675
R27 VP.n23 VP.n22 24.4675
R28 VP.n25 VP.n1 24.4675
R29 VP.n30 VP.n29 24.4675
R30 VP.n13 VP.n12 24.4675
R31 VP.n8 VP.n5 24.4675
R32 VP.n9 VP.n6 18.144
R33 VP.n24 VP.n23 12.234
R34 VP.n25 VP.n24 12.234
R35 VP.n8 VP.n7 12.234
R36 VP.n18 VP.n17 6.36192
R37 VP.n31 VP.n30 6.36192
R38 VP.n14 VP.n13 6.36192
R39 VP.n10 VP.n9 0.189894
R40 VP.n11 VP.n10 0.189894
R41 VP.n11 VP.n4 0.189894
R42 VP.n15 VP.n4 0.189894
R43 VP.n19 VP.n16 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n21 VP.n20 0.189894
R46 VP.n21 VP.n2 0.189894
R47 VP.n26 VP.n2 0.189894
R48 VP.n27 VP.n26 0.189894
R49 VP.n28 VP.n27 0.189894
R50 VP.n28 VP.n0 0.189894
R51 VP.n32 VP.n0 0.189894
R52 VP VP.n32 0.0516364
R53 VDD1.n102 VDD1.n101 289.615
R54 VDD1.n205 VDD1.n204 289.615
R55 VDD1.n101 VDD1.n100 185
R56 VDD1.n2 VDD1.n1 185
R57 VDD1.n95 VDD1.n94 185
R58 VDD1.n93 VDD1.n92 185
R59 VDD1.n6 VDD1.n5 185
R60 VDD1.n87 VDD1.n86 185
R61 VDD1.n85 VDD1.n84 185
R62 VDD1.n10 VDD1.n9 185
R63 VDD1.n79 VDD1.n78 185
R64 VDD1.n77 VDD1.n76 185
R65 VDD1.n14 VDD1.n13 185
R66 VDD1.n71 VDD1.n70 185
R67 VDD1.n69 VDD1.n68 185
R68 VDD1.n18 VDD1.n17 185
R69 VDD1.n63 VDD1.n62 185
R70 VDD1.n61 VDD1.n60 185
R71 VDD1.n22 VDD1.n21 185
R72 VDD1.n26 VDD1.n24 185
R73 VDD1.n55 VDD1.n54 185
R74 VDD1.n53 VDD1.n52 185
R75 VDD1.n28 VDD1.n27 185
R76 VDD1.n47 VDD1.n46 185
R77 VDD1.n45 VDD1.n44 185
R78 VDD1.n32 VDD1.n31 185
R79 VDD1.n39 VDD1.n38 185
R80 VDD1.n37 VDD1.n36 185
R81 VDD1.n138 VDD1.n137 185
R82 VDD1.n140 VDD1.n139 185
R83 VDD1.n133 VDD1.n132 185
R84 VDD1.n146 VDD1.n145 185
R85 VDD1.n148 VDD1.n147 185
R86 VDD1.n129 VDD1.n128 185
R87 VDD1.n155 VDD1.n154 185
R88 VDD1.n156 VDD1.n127 185
R89 VDD1.n158 VDD1.n157 185
R90 VDD1.n125 VDD1.n124 185
R91 VDD1.n164 VDD1.n163 185
R92 VDD1.n166 VDD1.n165 185
R93 VDD1.n121 VDD1.n120 185
R94 VDD1.n172 VDD1.n171 185
R95 VDD1.n174 VDD1.n173 185
R96 VDD1.n117 VDD1.n116 185
R97 VDD1.n180 VDD1.n179 185
R98 VDD1.n182 VDD1.n181 185
R99 VDD1.n113 VDD1.n112 185
R100 VDD1.n188 VDD1.n187 185
R101 VDD1.n190 VDD1.n189 185
R102 VDD1.n109 VDD1.n108 185
R103 VDD1.n196 VDD1.n195 185
R104 VDD1.n198 VDD1.n197 185
R105 VDD1.n105 VDD1.n104 185
R106 VDD1.n204 VDD1.n203 185
R107 VDD1.n35 VDD1.t0 149.524
R108 VDD1.n136 VDD1.t1 149.524
R109 VDD1.n101 VDD1.n1 104.615
R110 VDD1.n94 VDD1.n1 104.615
R111 VDD1.n94 VDD1.n93 104.615
R112 VDD1.n93 VDD1.n5 104.615
R113 VDD1.n86 VDD1.n5 104.615
R114 VDD1.n86 VDD1.n85 104.615
R115 VDD1.n85 VDD1.n9 104.615
R116 VDD1.n78 VDD1.n9 104.615
R117 VDD1.n78 VDD1.n77 104.615
R118 VDD1.n77 VDD1.n13 104.615
R119 VDD1.n70 VDD1.n13 104.615
R120 VDD1.n70 VDD1.n69 104.615
R121 VDD1.n69 VDD1.n17 104.615
R122 VDD1.n62 VDD1.n17 104.615
R123 VDD1.n62 VDD1.n61 104.615
R124 VDD1.n61 VDD1.n21 104.615
R125 VDD1.n26 VDD1.n21 104.615
R126 VDD1.n54 VDD1.n26 104.615
R127 VDD1.n54 VDD1.n53 104.615
R128 VDD1.n53 VDD1.n27 104.615
R129 VDD1.n46 VDD1.n27 104.615
R130 VDD1.n46 VDD1.n45 104.615
R131 VDD1.n45 VDD1.n31 104.615
R132 VDD1.n38 VDD1.n31 104.615
R133 VDD1.n38 VDD1.n37 104.615
R134 VDD1.n139 VDD1.n138 104.615
R135 VDD1.n139 VDD1.n132 104.615
R136 VDD1.n146 VDD1.n132 104.615
R137 VDD1.n147 VDD1.n146 104.615
R138 VDD1.n147 VDD1.n128 104.615
R139 VDD1.n155 VDD1.n128 104.615
R140 VDD1.n156 VDD1.n155 104.615
R141 VDD1.n157 VDD1.n156 104.615
R142 VDD1.n157 VDD1.n124 104.615
R143 VDD1.n164 VDD1.n124 104.615
R144 VDD1.n165 VDD1.n164 104.615
R145 VDD1.n165 VDD1.n120 104.615
R146 VDD1.n172 VDD1.n120 104.615
R147 VDD1.n173 VDD1.n172 104.615
R148 VDD1.n173 VDD1.n116 104.615
R149 VDD1.n180 VDD1.n116 104.615
R150 VDD1.n181 VDD1.n180 104.615
R151 VDD1.n181 VDD1.n112 104.615
R152 VDD1.n188 VDD1.n112 104.615
R153 VDD1.n189 VDD1.n188 104.615
R154 VDD1.n189 VDD1.n108 104.615
R155 VDD1.n196 VDD1.n108 104.615
R156 VDD1.n197 VDD1.n196 104.615
R157 VDD1.n197 VDD1.n104 104.615
R158 VDD1.n204 VDD1.n104 104.615
R159 VDD1.n207 VDD1.n206 64.5906
R160 VDD1.n209 VDD1.n208 64.2406
R161 VDD1 VDD1.n102 53.8227
R162 VDD1.n207 VDD1.n205 53.7092
R163 VDD1.n37 VDD1.t0 52.3082
R164 VDD1.n138 VDD1.t1 52.3082
R165 VDD1.n209 VDD1.n207 46.5914
R166 VDD1.n24 VDD1.n22 13.1884
R167 VDD1.n158 VDD1.n125 13.1884
R168 VDD1.n100 VDD1.n0 12.8005
R169 VDD1.n60 VDD1.n59 12.8005
R170 VDD1.n56 VDD1.n55 12.8005
R171 VDD1.n159 VDD1.n127 12.8005
R172 VDD1.n163 VDD1.n162 12.8005
R173 VDD1.n203 VDD1.n103 12.8005
R174 VDD1.n99 VDD1.n2 12.0247
R175 VDD1.n63 VDD1.n20 12.0247
R176 VDD1.n52 VDD1.n25 12.0247
R177 VDD1.n154 VDD1.n153 12.0247
R178 VDD1.n166 VDD1.n123 12.0247
R179 VDD1.n202 VDD1.n105 12.0247
R180 VDD1.n96 VDD1.n95 11.249
R181 VDD1.n64 VDD1.n18 11.249
R182 VDD1.n51 VDD1.n28 11.249
R183 VDD1.n152 VDD1.n129 11.249
R184 VDD1.n167 VDD1.n121 11.249
R185 VDD1.n199 VDD1.n198 11.249
R186 VDD1.n92 VDD1.n4 10.4732
R187 VDD1.n68 VDD1.n67 10.4732
R188 VDD1.n48 VDD1.n47 10.4732
R189 VDD1.n149 VDD1.n148 10.4732
R190 VDD1.n171 VDD1.n170 10.4732
R191 VDD1.n195 VDD1.n107 10.4732
R192 VDD1.n36 VDD1.n35 10.2747
R193 VDD1.n137 VDD1.n136 10.2747
R194 VDD1.n91 VDD1.n6 9.69747
R195 VDD1.n71 VDD1.n16 9.69747
R196 VDD1.n44 VDD1.n30 9.69747
R197 VDD1.n145 VDD1.n131 9.69747
R198 VDD1.n174 VDD1.n119 9.69747
R199 VDD1.n194 VDD1.n109 9.69747
R200 VDD1.n98 VDD1.n0 9.45567
R201 VDD1.n201 VDD1.n103 9.45567
R202 VDD1.n34 VDD1.n33 9.3005
R203 VDD1.n41 VDD1.n40 9.3005
R204 VDD1.n43 VDD1.n42 9.3005
R205 VDD1.n30 VDD1.n29 9.3005
R206 VDD1.n49 VDD1.n48 9.3005
R207 VDD1.n51 VDD1.n50 9.3005
R208 VDD1.n25 VDD1.n23 9.3005
R209 VDD1.n57 VDD1.n56 9.3005
R210 VDD1.n83 VDD1.n82 9.3005
R211 VDD1.n8 VDD1.n7 9.3005
R212 VDD1.n89 VDD1.n88 9.3005
R213 VDD1.n91 VDD1.n90 9.3005
R214 VDD1.n4 VDD1.n3 9.3005
R215 VDD1.n97 VDD1.n96 9.3005
R216 VDD1.n99 VDD1.n98 9.3005
R217 VDD1.n81 VDD1.n80 9.3005
R218 VDD1.n12 VDD1.n11 9.3005
R219 VDD1.n75 VDD1.n74 9.3005
R220 VDD1.n73 VDD1.n72 9.3005
R221 VDD1.n16 VDD1.n15 9.3005
R222 VDD1.n67 VDD1.n66 9.3005
R223 VDD1.n65 VDD1.n64 9.3005
R224 VDD1.n20 VDD1.n19 9.3005
R225 VDD1.n59 VDD1.n58 9.3005
R226 VDD1.n184 VDD1.n183 9.3005
R227 VDD1.n186 VDD1.n185 9.3005
R228 VDD1.n111 VDD1.n110 9.3005
R229 VDD1.n192 VDD1.n191 9.3005
R230 VDD1.n194 VDD1.n193 9.3005
R231 VDD1.n107 VDD1.n106 9.3005
R232 VDD1.n200 VDD1.n199 9.3005
R233 VDD1.n202 VDD1.n201 9.3005
R234 VDD1.n178 VDD1.n177 9.3005
R235 VDD1.n176 VDD1.n175 9.3005
R236 VDD1.n119 VDD1.n118 9.3005
R237 VDD1.n170 VDD1.n169 9.3005
R238 VDD1.n168 VDD1.n167 9.3005
R239 VDD1.n123 VDD1.n122 9.3005
R240 VDD1.n162 VDD1.n161 9.3005
R241 VDD1.n135 VDD1.n134 9.3005
R242 VDD1.n142 VDD1.n141 9.3005
R243 VDD1.n144 VDD1.n143 9.3005
R244 VDD1.n131 VDD1.n130 9.3005
R245 VDD1.n150 VDD1.n149 9.3005
R246 VDD1.n152 VDD1.n151 9.3005
R247 VDD1.n153 VDD1.n126 9.3005
R248 VDD1.n160 VDD1.n159 9.3005
R249 VDD1.n115 VDD1.n114 9.3005
R250 VDD1.n88 VDD1.n87 8.92171
R251 VDD1.n72 VDD1.n14 8.92171
R252 VDD1.n43 VDD1.n32 8.92171
R253 VDD1.n144 VDD1.n133 8.92171
R254 VDD1.n175 VDD1.n117 8.92171
R255 VDD1.n191 VDD1.n190 8.92171
R256 VDD1.n84 VDD1.n8 8.14595
R257 VDD1.n76 VDD1.n75 8.14595
R258 VDD1.n40 VDD1.n39 8.14595
R259 VDD1.n141 VDD1.n140 8.14595
R260 VDD1.n179 VDD1.n178 8.14595
R261 VDD1.n187 VDD1.n111 8.14595
R262 VDD1.n83 VDD1.n10 7.3702
R263 VDD1.n79 VDD1.n12 7.3702
R264 VDD1.n36 VDD1.n34 7.3702
R265 VDD1.n137 VDD1.n135 7.3702
R266 VDD1.n182 VDD1.n115 7.3702
R267 VDD1.n186 VDD1.n113 7.3702
R268 VDD1.n80 VDD1.n10 6.59444
R269 VDD1.n80 VDD1.n79 6.59444
R270 VDD1.n183 VDD1.n182 6.59444
R271 VDD1.n183 VDD1.n113 6.59444
R272 VDD1.n84 VDD1.n83 5.81868
R273 VDD1.n76 VDD1.n12 5.81868
R274 VDD1.n39 VDD1.n34 5.81868
R275 VDD1.n140 VDD1.n135 5.81868
R276 VDD1.n179 VDD1.n115 5.81868
R277 VDD1.n187 VDD1.n186 5.81868
R278 VDD1.n87 VDD1.n8 5.04292
R279 VDD1.n75 VDD1.n14 5.04292
R280 VDD1.n40 VDD1.n32 5.04292
R281 VDD1.n141 VDD1.n133 5.04292
R282 VDD1.n178 VDD1.n117 5.04292
R283 VDD1.n190 VDD1.n111 5.04292
R284 VDD1.n88 VDD1.n6 4.26717
R285 VDD1.n72 VDD1.n71 4.26717
R286 VDD1.n44 VDD1.n43 4.26717
R287 VDD1.n145 VDD1.n144 4.26717
R288 VDD1.n175 VDD1.n174 4.26717
R289 VDD1.n191 VDD1.n109 4.26717
R290 VDD1.n92 VDD1.n91 3.49141
R291 VDD1.n68 VDD1.n16 3.49141
R292 VDD1.n47 VDD1.n30 3.49141
R293 VDD1.n148 VDD1.n131 3.49141
R294 VDD1.n171 VDD1.n119 3.49141
R295 VDD1.n195 VDD1.n194 3.49141
R296 VDD1.n136 VDD1.n134 2.84303
R297 VDD1.n35 VDD1.n33 2.84303
R298 VDD1.n95 VDD1.n4 2.71565
R299 VDD1.n67 VDD1.n18 2.71565
R300 VDD1.n48 VDD1.n28 2.71565
R301 VDD1.n149 VDD1.n129 2.71565
R302 VDD1.n170 VDD1.n121 2.71565
R303 VDD1.n198 VDD1.n107 2.71565
R304 VDD1.n96 VDD1.n2 1.93989
R305 VDD1.n64 VDD1.n63 1.93989
R306 VDD1.n52 VDD1.n51 1.93989
R307 VDD1.n154 VDD1.n152 1.93989
R308 VDD1.n167 VDD1.n166 1.93989
R309 VDD1.n199 VDD1.n105 1.93989
R310 VDD1.n100 VDD1.n99 1.16414
R311 VDD1.n60 VDD1.n20 1.16414
R312 VDD1.n55 VDD1.n25 1.16414
R313 VDD1.n153 VDD1.n127 1.16414
R314 VDD1.n163 VDD1.n123 1.16414
R315 VDD1.n203 VDD1.n202 1.16414
R316 VDD1.n208 VDD1.t3 1.05313
R317 VDD1.n208 VDD1.t5 1.05313
R318 VDD1.n206 VDD1.t2 1.05313
R319 VDD1.n206 VDD1.t4 1.05313
R320 VDD1.n102 VDD1.n0 0.388379
R321 VDD1.n59 VDD1.n22 0.388379
R322 VDD1.n56 VDD1.n24 0.388379
R323 VDD1.n159 VDD1.n158 0.388379
R324 VDD1.n162 VDD1.n125 0.388379
R325 VDD1.n205 VDD1.n103 0.388379
R326 VDD1 VDD1.n209 0.347483
R327 VDD1.n98 VDD1.n97 0.155672
R328 VDD1.n97 VDD1.n3 0.155672
R329 VDD1.n90 VDD1.n3 0.155672
R330 VDD1.n90 VDD1.n89 0.155672
R331 VDD1.n89 VDD1.n7 0.155672
R332 VDD1.n82 VDD1.n7 0.155672
R333 VDD1.n82 VDD1.n81 0.155672
R334 VDD1.n81 VDD1.n11 0.155672
R335 VDD1.n74 VDD1.n11 0.155672
R336 VDD1.n74 VDD1.n73 0.155672
R337 VDD1.n73 VDD1.n15 0.155672
R338 VDD1.n66 VDD1.n15 0.155672
R339 VDD1.n66 VDD1.n65 0.155672
R340 VDD1.n65 VDD1.n19 0.155672
R341 VDD1.n58 VDD1.n19 0.155672
R342 VDD1.n58 VDD1.n57 0.155672
R343 VDD1.n57 VDD1.n23 0.155672
R344 VDD1.n50 VDD1.n23 0.155672
R345 VDD1.n50 VDD1.n49 0.155672
R346 VDD1.n49 VDD1.n29 0.155672
R347 VDD1.n42 VDD1.n29 0.155672
R348 VDD1.n42 VDD1.n41 0.155672
R349 VDD1.n41 VDD1.n33 0.155672
R350 VDD1.n142 VDD1.n134 0.155672
R351 VDD1.n143 VDD1.n142 0.155672
R352 VDD1.n143 VDD1.n130 0.155672
R353 VDD1.n150 VDD1.n130 0.155672
R354 VDD1.n151 VDD1.n150 0.155672
R355 VDD1.n151 VDD1.n126 0.155672
R356 VDD1.n160 VDD1.n126 0.155672
R357 VDD1.n161 VDD1.n160 0.155672
R358 VDD1.n161 VDD1.n122 0.155672
R359 VDD1.n168 VDD1.n122 0.155672
R360 VDD1.n169 VDD1.n168 0.155672
R361 VDD1.n169 VDD1.n118 0.155672
R362 VDD1.n176 VDD1.n118 0.155672
R363 VDD1.n177 VDD1.n176 0.155672
R364 VDD1.n177 VDD1.n114 0.155672
R365 VDD1.n184 VDD1.n114 0.155672
R366 VDD1.n185 VDD1.n184 0.155672
R367 VDD1.n185 VDD1.n110 0.155672
R368 VDD1.n192 VDD1.n110 0.155672
R369 VDD1.n193 VDD1.n192 0.155672
R370 VDD1.n193 VDD1.n106 0.155672
R371 VDD1.n200 VDD1.n106 0.155672
R372 VDD1.n201 VDD1.n200 0.155672
R373 VTAIL.n422 VTAIL.n421 289.615
R374 VTAIL.n104 VTAIL.n103 289.615
R375 VTAIL.n318 VTAIL.n317 289.615
R376 VTAIL.n212 VTAIL.n211 289.615
R377 VTAIL.n355 VTAIL.n354 185
R378 VTAIL.n357 VTAIL.n356 185
R379 VTAIL.n350 VTAIL.n349 185
R380 VTAIL.n363 VTAIL.n362 185
R381 VTAIL.n365 VTAIL.n364 185
R382 VTAIL.n346 VTAIL.n345 185
R383 VTAIL.n372 VTAIL.n371 185
R384 VTAIL.n373 VTAIL.n344 185
R385 VTAIL.n375 VTAIL.n374 185
R386 VTAIL.n342 VTAIL.n341 185
R387 VTAIL.n381 VTAIL.n380 185
R388 VTAIL.n383 VTAIL.n382 185
R389 VTAIL.n338 VTAIL.n337 185
R390 VTAIL.n389 VTAIL.n388 185
R391 VTAIL.n391 VTAIL.n390 185
R392 VTAIL.n334 VTAIL.n333 185
R393 VTAIL.n397 VTAIL.n396 185
R394 VTAIL.n399 VTAIL.n398 185
R395 VTAIL.n330 VTAIL.n329 185
R396 VTAIL.n405 VTAIL.n404 185
R397 VTAIL.n407 VTAIL.n406 185
R398 VTAIL.n326 VTAIL.n325 185
R399 VTAIL.n413 VTAIL.n412 185
R400 VTAIL.n415 VTAIL.n414 185
R401 VTAIL.n322 VTAIL.n321 185
R402 VTAIL.n421 VTAIL.n420 185
R403 VTAIL.n37 VTAIL.n36 185
R404 VTAIL.n39 VTAIL.n38 185
R405 VTAIL.n32 VTAIL.n31 185
R406 VTAIL.n45 VTAIL.n44 185
R407 VTAIL.n47 VTAIL.n46 185
R408 VTAIL.n28 VTAIL.n27 185
R409 VTAIL.n54 VTAIL.n53 185
R410 VTAIL.n55 VTAIL.n26 185
R411 VTAIL.n57 VTAIL.n56 185
R412 VTAIL.n24 VTAIL.n23 185
R413 VTAIL.n63 VTAIL.n62 185
R414 VTAIL.n65 VTAIL.n64 185
R415 VTAIL.n20 VTAIL.n19 185
R416 VTAIL.n71 VTAIL.n70 185
R417 VTAIL.n73 VTAIL.n72 185
R418 VTAIL.n16 VTAIL.n15 185
R419 VTAIL.n79 VTAIL.n78 185
R420 VTAIL.n81 VTAIL.n80 185
R421 VTAIL.n12 VTAIL.n11 185
R422 VTAIL.n87 VTAIL.n86 185
R423 VTAIL.n89 VTAIL.n88 185
R424 VTAIL.n8 VTAIL.n7 185
R425 VTAIL.n95 VTAIL.n94 185
R426 VTAIL.n97 VTAIL.n96 185
R427 VTAIL.n4 VTAIL.n3 185
R428 VTAIL.n103 VTAIL.n102 185
R429 VTAIL.n317 VTAIL.n316 185
R430 VTAIL.n218 VTAIL.n217 185
R431 VTAIL.n311 VTAIL.n310 185
R432 VTAIL.n309 VTAIL.n308 185
R433 VTAIL.n222 VTAIL.n221 185
R434 VTAIL.n303 VTAIL.n302 185
R435 VTAIL.n301 VTAIL.n300 185
R436 VTAIL.n226 VTAIL.n225 185
R437 VTAIL.n295 VTAIL.n294 185
R438 VTAIL.n293 VTAIL.n292 185
R439 VTAIL.n230 VTAIL.n229 185
R440 VTAIL.n287 VTAIL.n286 185
R441 VTAIL.n285 VTAIL.n284 185
R442 VTAIL.n234 VTAIL.n233 185
R443 VTAIL.n279 VTAIL.n278 185
R444 VTAIL.n277 VTAIL.n276 185
R445 VTAIL.n238 VTAIL.n237 185
R446 VTAIL.n242 VTAIL.n240 185
R447 VTAIL.n271 VTAIL.n270 185
R448 VTAIL.n269 VTAIL.n268 185
R449 VTAIL.n244 VTAIL.n243 185
R450 VTAIL.n263 VTAIL.n262 185
R451 VTAIL.n261 VTAIL.n260 185
R452 VTAIL.n248 VTAIL.n247 185
R453 VTAIL.n255 VTAIL.n254 185
R454 VTAIL.n253 VTAIL.n252 185
R455 VTAIL.n211 VTAIL.n210 185
R456 VTAIL.n112 VTAIL.n111 185
R457 VTAIL.n205 VTAIL.n204 185
R458 VTAIL.n203 VTAIL.n202 185
R459 VTAIL.n116 VTAIL.n115 185
R460 VTAIL.n197 VTAIL.n196 185
R461 VTAIL.n195 VTAIL.n194 185
R462 VTAIL.n120 VTAIL.n119 185
R463 VTAIL.n189 VTAIL.n188 185
R464 VTAIL.n187 VTAIL.n186 185
R465 VTAIL.n124 VTAIL.n123 185
R466 VTAIL.n181 VTAIL.n180 185
R467 VTAIL.n179 VTAIL.n178 185
R468 VTAIL.n128 VTAIL.n127 185
R469 VTAIL.n173 VTAIL.n172 185
R470 VTAIL.n171 VTAIL.n170 185
R471 VTAIL.n132 VTAIL.n131 185
R472 VTAIL.n136 VTAIL.n134 185
R473 VTAIL.n165 VTAIL.n164 185
R474 VTAIL.n163 VTAIL.n162 185
R475 VTAIL.n138 VTAIL.n137 185
R476 VTAIL.n157 VTAIL.n156 185
R477 VTAIL.n155 VTAIL.n154 185
R478 VTAIL.n142 VTAIL.n141 185
R479 VTAIL.n149 VTAIL.n148 185
R480 VTAIL.n147 VTAIL.n146 185
R481 VTAIL.n353 VTAIL.t5 149.524
R482 VTAIL.n35 VTAIL.t6 149.524
R483 VTAIL.n251 VTAIL.t7 149.524
R484 VTAIL.n145 VTAIL.t0 149.524
R485 VTAIL.n356 VTAIL.n355 104.615
R486 VTAIL.n356 VTAIL.n349 104.615
R487 VTAIL.n363 VTAIL.n349 104.615
R488 VTAIL.n364 VTAIL.n363 104.615
R489 VTAIL.n364 VTAIL.n345 104.615
R490 VTAIL.n372 VTAIL.n345 104.615
R491 VTAIL.n373 VTAIL.n372 104.615
R492 VTAIL.n374 VTAIL.n373 104.615
R493 VTAIL.n374 VTAIL.n341 104.615
R494 VTAIL.n381 VTAIL.n341 104.615
R495 VTAIL.n382 VTAIL.n381 104.615
R496 VTAIL.n382 VTAIL.n337 104.615
R497 VTAIL.n389 VTAIL.n337 104.615
R498 VTAIL.n390 VTAIL.n389 104.615
R499 VTAIL.n390 VTAIL.n333 104.615
R500 VTAIL.n397 VTAIL.n333 104.615
R501 VTAIL.n398 VTAIL.n397 104.615
R502 VTAIL.n398 VTAIL.n329 104.615
R503 VTAIL.n405 VTAIL.n329 104.615
R504 VTAIL.n406 VTAIL.n405 104.615
R505 VTAIL.n406 VTAIL.n325 104.615
R506 VTAIL.n413 VTAIL.n325 104.615
R507 VTAIL.n414 VTAIL.n413 104.615
R508 VTAIL.n414 VTAIL.n321 104.615
R509 VTAIL.n421 VTAIL.n321 104.615
R510 VTAIL.n38 VTAIL.n37 104.615
R511 VTAIL.n38 VTAIL.n31 104.615
R512 VTAIL.n45 VTAIL.n31 104.615
R513 VTAIL.n46 VTAIL.n45 104.615
R514 VTAIL.n46 VTAIL.n27 104.615
R515 VTAIL.n54 VTAIL.n27 104.615
R516 VTAIL.n55 VTAIL.n54 104.615
R517 VTAIL.n56 VTAIL.n55 104.615
R518 VTAIL.n56 VTAIL.n23 104.615
R519 VTAIL.n63 VTAIL.n23 104.615
R520 VTAIL.n64 VTAIL.n63 104.615
R521 VTAIL.n64 VTAIL.n19 104.615
R522 VTAIL.n71 VTAIL.n19 104.615
R523 VTAIL.n72 VTAIL.n71 104.615
R524 VTAIL.n72 VTAIL.n15 104.615
R525 VTAIL.n79 VTAIL.n15 104.615
R526 VTAIL.n80 VTAIL.n79 104.615
R527 VTAIL.n80 VTAIL.n11 104.615
R528 VTAIL.n87 VTAIL.n11 104.615
R529 VTAIL.n88 VTAIL.n87 104.615
R530 VTAIL.n88 VTAIL.n7 104.615
R531 VTAIL.n95 VTAIL.n7 104.615
R532 VTAIL.n96 VTAIL.n95 104.615
R533 VTAIL.n96 VTAIL.n3 104.615
R534 VTAIL.n103 VTAIL.n3 104.615
R535 VTAIL.n317 VTAIL.n217 104.615
R536 VTAIL.n310 VTAIL.n217 104.615
R537 VTAIL.n310 VTAIL.n309 104.615
R538 VTAIL.n309 VTAIL.n221 104.615
R539 VTAIL.n302 VTAIL.n221 104.615
R540 VTAIL.n302 VTAIL.n301 104.615
R541 VTAIL.n301 VTAIL.n225 104.615
R542 VTAIL.n294 VTAIL.n225 104.615
R543 VTAIL.n294 VTAIL.n293 104.615
R544 VTAIL.n293 VTAIL.n229 104.615
R545 VTAIL.n286 VTAIL.n229 104.615
R546 VTAIL.n286 VTAIL.n285 104.615
R547 VTAIL.n285 VTAIL.n233 104.615
R548 VTAIL.n278 VTAIL.n233 104.615
R549 VTAIL.n278 VTAIL.n277 104.615
R550 VTAIL.n277 VTAIL.n237 104.615
R551 VTAIL.n242 VTAIL.n237 104.615
R552 VTAIL.n270 VTAIL.n242 104.615
R553 VTAIL.n270 VTAIL.n269 104.615
R554 VTAIL.n269 VTAIL.n243 104.615
R555 VTAIL.n262 VTAIL.n243 104.615
R556 VTAIL.n262 VTAIL.n261 104.615
R557 VTAIL.n261 VTAIL.n247 104.615
R558 VTAIL.n254 VTAIL.n247 104.615
R559 VTAIL.n254 VTAIL.n253 104.615
R560 VTAIL.n211 VTAIL.n111 104.615
R561 VTAIL.n204 VTAIL.n111 104.615
R562 VTAIL.n204 VTAIL.n203 104.615
R563 VTAIL.n203 VTAIL.n115 104.615
R564 VTAIL.n196 VTAIL.n115 104.615
R565 VTAIL.n196 VTAIL.n195 104.615
R566 VTAIL.n195 VTAIL.n119 104.615
R567 VTAIL.n188 VTAIL.n119 104.615
R568 VTAIL.n188 VTAIL.n187 104.615
R569 VTAIL.n187 VTAIL.n123 104.615
R570 VTAIL.n180 VTAIL.n123 104.615
R571 VTAIL.n180 VTAIL.n179 104.615
R572 VTAIL.n179 VTAIL.n127 104.615
R573 VTAIL.n172 VTAIL.n127 104.615
R574 VTAIL.n172 VTAIL.n171 104.615
R575 VTAIL.n171 VTAIL.n131 104.615
R576 VTAIL.n136 VTAIL.n131 104.615
R577 VTAIL.n164 VTAIL.n136 104.615
R578 VTAIL.n164 VTAIL.n163 104.615
R579 VTAIL.n163 VTAIL.n137 104.615
R580 VTAIL.n156 VTAIL.n137 104.615
R581 VTAIL.n156 VTAIL.n155 104.615
R582 VTAIL.n155 VTAIL.n141 104.615
R583 VTAIL.n148 VTAIL.n141 104.615
R584 VTAIL.n148 VTAIL.n147 104.615
R585 VTAIL.n355 VTAIL.t5 52.3082
R586 VTAIL.n37 VTAIL.t6 52.3082
R587 VTAIL.n253 VTAIL.t7 52.3082
R588 VTAIL.n147 VTAIL.t0 52.3082
R589 VTAIL.n215 VTAIL.n214 47.563
R590 VTAIL.n109 VTAIL.n108 47.563
R591 VTAIL.n1 VTAIL.n0 47.562
R592 VTAIL.n107 VTAIL.n106 47.562
R593 VTAIL.n423 VTAIL.n422 35.8702
R594 VTAIL.n105 VTAIL.n104 35.8702
R595 VTAIL.n319 VTAIL.n318 35.8702
R596 VTAIL.n213 VTAIL.n212 35.8702
R597 VTAIL.n109 VTAIL.n107 31.8238
R598 VTAIL.n423 VTAIL.n319 30.2031
R599 VTAIL.n375 VTAIL.n342 13.1884
R600 VTAIL.n57 VTAIL.n24 13.1884
R601 VTAIL.n240 VTAIL.n238 13.1884
R602 VTAIL.n134 VTAIL.n132 13.1884
R603 VTAIL.n376 VTAIL.n344 12.8005
R604 VTAIL.n380 VTAIL.n379 12.8005
R605 VTAIL.n420 VTAIL.n320 12.8005
R606 VTAIL.n58 VTAIL.n26 12.8005
R607 VTAIL.n62 VTAIL.n61 12.8005
R608 VTAIL.n102 VTAIL.n2 12.8005
R609 VTAIL.n316 VTAIL.n216 12.8005
R610 VTAIL.n276 VTAIL.n275 12.8005
R611 VTAIL.n272 VTAIL.n271 12.8005
R612 VTAIL.n210 VTAIL.n110 12.8005
R613 VTAIL.n170 VTAIL.n169 12.8005
R614 VTAIL.n166 VTAIL.n165 12.8005
R615 VTAIL.n371 VTAIL.n370 12.0247
R616 VTAIL.n383 VTAIL.n340 12.0247
R617 VTAIL.n419 VTAIL.n322 12.0247
R618 VTAIL.n53 VTAIL.n52 12.0247
R619 VTAIL.n65 VTAIL.n22 12.0247
R620 VTAIL.n101 VTAIL.n4 12.0247
R621 VTAIL.n315 VTAIL.n218 12.0247
R622 VTAIL.n279 VTAIL.n236 12.0247
R623 VTAIL.n268 VTAIL.n241 12.0247
R624 VTAIL.n209 VTAIL.n112 12.0247
R625 VTAIL.n173 VTAIL.n130 12.0247
R626 VTAIL.n162 VTAIL.n135 12.0247
R627 VTAIL.n369 VTAIL.n346 11.249
R628 VTAIL.n384 VTAIL.n338 11.249
R629 VTAIL.n416 VTAIL.n415 11.249
R630 VTAIL.n51 VTAIL.n28 11.249
R631 VTAIL.n66 VTAIL.n20 11.249
R632 VTAIL.n98 VTAIL.n97 11.249
R633 VTAIL.n312 VTAIL.n311 11.249
R634 VTAIL.n280 VTAIL.n234 11.249
R635 VTAIL.n267 VTAIL.n244 11.249
R636 VTAIL.n206 VTAIL.n205 11.249
R637 VTAIL.n174 VTAIL.n128 11.249
R638 VTAIL.n161 VTAIL.n138 11.249
R639 VTAIL.n366 VTAIL.n365 10.4732
R640 VTAIL.n388 VTAIL.n387 10.4732
R641 VTAIL.n412 VTAIL.n324 10.4732
R642 VTAIL.n48 VTAIL.n47 10.4732
R643 VTAIL.n70 VTAIL.n69 10.4732
R644 VTAIL.n94 VTAIL.n6 10.4732
R645 VTAIL.n308 VTAIL.n220 10.4732
R646 VTAIL.n284 VTAIL.n283 10.4732
R647 VTAIL.n264 VTAIL.n263 10.4732
R648 VTAIL.n202 VTAIL.n114 10.4732
R649 VTAIL.n178 VTAIL.n177 10.4732
R650 VTAIL.n158 VTAIL.n157 10.4732
R651 VTAIL.n354 VTAIL.n353 10.2747
R652 VTAIL.n36 VTAIL.n35 10.2747
R653 VTAIL.n252 VTAIL.n251 10.2747
R654 VTAIL.n146 VTAIL.n145 10.2747
R655 VTAIL.n362 VTAIL.n348 9.69747
R656 VTAIL.n391 VTAIL.n336 9.69747
R657 VTAIL.n411 VTAIL.n326 9.69747
R658 VTAIL.n44 VTAIL.n30 9.69747
R659 VTAIL.n73 VTAIL.n18 9.69747
R660 VTAIL.n93 VTAIL.n8 9.69747
R661 VTAIL.n307 VTAIL.n222 9.69747
R662 VTAIL.n287 VTAIL.n232 9.69747
R663 VTAIL.n260 VTAIL.n246 9.69747
R664 VTAIL.n201 VTAIL.n116 9.69747
R665 VTAIL.n181 VTAIL.n126 9.69747
R666 VTAIL.n154 VTAIL.n140 9.69747
R667 VTAIL.n418 VTAIL.n320 9.45567
R668 VTAIL.n100 VTAIL.n2 9.45567
R669 VTAIL.n314 VTAIL.n216 9.45567
R670 VTAIL.n208 VTAIL.n110 9.45567
R671 VTAIL.n401 VTAIL.n400 9.3005
R672 VTAIL.n403 VTAIL.n402 9.3005
R673 VTAIL.n328 VTAIL.n327 9.3005
R674 VTAIL.n409 VTAIL.n408 9.3005
R675 VTAIL.n411 VTAIL.n410 9.3005
R676 VTAIL.n324 VTAIL.n323 9.3005
R677 VTAIL.n417 VTAIL.n416 9.3005
R678 VTAIL.n419 VTAIL.n418 9.3005
R679 VTAIL.n395 VTAIL.n394 9.3005
R680 VTAIL.n393 VTAIL.n392 9.3005
R681 VTAIL.n336 VTAIL.n335 9.3005
R682 VTAIL.n387 VTAIL.n386 9.3005
R683 VTAIL.n385 VTAIL.n384 9.3005
R684 VTAIL.n340 VTAIL.n339 9.3005
R685 VTAIL.n379 VTAIL.n378 9.3005
R686 VTAIL.n352 VTAIL.n351 9.3005
R687 VTAIL.n359 VTAIL.n358 9.3005
R688 VTAIL.n361 VTAIL.n360 9.3005
R689 VTAIL.n348 VTAIL.n347 9.3005
R690 VTAIL.n367 VTAIL.n366 9.3005
R691 VTAIL.n369 VTAIL.n368 9.3005
R692 VTAIL.n370 VTAIL.n343 9.3005
R693 VTAIL.n377 VTAIL.n376 9.3005
R694 VTAIL.n332 VTAIL.n331 9.3005
R695 VTAIL.n83 VTAIL.n82 9.3005
R696 VTAIL.n85 VTAIL.n84 9.3005
R697 VTAIL.n10 VTAIL.n9 9.3005
R698 VTAIL.n91 VTAIL.n90 9.3005
R699 VTAIL.n93 VTAIL.n92 9.3005
R700 VTAIL.n6 VTAIL.n5 9.3005
R701 VTAIL.n99 VTAIL.n98 9.3005
R702 VTAIL.n101 VTAIL.n100 9.3005
R703 VTAIL.n77 VTAIL.n76 9.3005
R704 VTAIL.n75 VTAIL.n74 9.3005
R705 VTAIL.n18 VTAIL.n17 9.3005
R706 VTAIL.n69 VTAIL.n68 9.3005
R707 VTAIL.n67 VTAIL.n66 9.3005
R708 VTAIL.n22 VTAIL.n21 9.3005
R709 VTAIL.n61 VTAIL.n60 9.3005
R710 VTAIL.n34 VTAIL.n33 9.3005
R711 VTAIL.n41 VTAIL.n40 9.3005
R712 VTAIL.n43 VTAIL.n42 9.3005
R713 VTAIL.n30 VTAIL.n29 9.3005
R714 VTAIL.n49 VTAIL.n48 9.3005
R715 VTAIL.n51 VTAIL.n50 9.3005
R716 VTAIL.n52 VTAIL.n25 9.3005
R717 VTAIL.n59 VTAIL.n58 9.3005
R718 VTAIL.n14 VTAIL.n13 9.3005
R719 VTAIL.n315 VTAIL.n314 9.3005
R720 VTAIL.n313 VTAIL.n312 9.3005
R721 VTAIL.n220 VTAIL.n219 9.3005
R722 VTAIL.n307 VTAIL.n306 9.3005
R723 VTAIL.n305 VTAIL.n304 9.3005
R724 VTAIL.n224 VTAIL.n223 9.3005
R725 VTAIL.n299 VTAIL.n298 9.3005
R726 VTAIL.n297 VTAIL.n296 9.3005
R727 VTAIL.n228 VTAIL.n227 9.3005
R728 VTAIL.n291 VTAIL.n290 9.3005
R729 VTAIL.n289 VTAIL.n288 9.3005
R730 VTAIL.n232 VTAIL.n231 9.3005
R731 VTAIL.n283 VTAIL.n282 9.3005
R732 VTAIL.n281 VTAIL.n280 9.3005
R733 VTAIL.n236 VTAIL.n235 9.3005
R734 VTAIL.n275 VTAIL.n274 9.3005
R735 VTAIL.n273 VTAIL.n272 9.3005
R736 VTAIL.n241 VTAIL.n239 9.3005
R737 VTAIL.n267 VTAIL.n266 9.3005
R738 VTAIL.n265 VTAIL.n264 9.3005
R739 VTAIL.n246 VTAIL.n245 9.3005
R740 VTAIL.n259 VTAIL.n258 9.3005
R741 VTAIL.n257 VTAIL.n256 9.3005
R742 VTAIL.n250 VTAIL.n249 9.3005
R743 VTAIL.n144 VTAIL.n143 9.3005
R744 VTAIL.n151 VTAIL.n150 9.3005
R745 VTAIL.n153 VTAIL.n152 9.3005
R746 VTAIL.n140 VTAIL.n139 9.3005
R747 VTAIL.n159 VTAIL.n158 9.3005
R748 VTAIL.n161 VTAIL.n160 9.3005
R749 VTAIL.n135 VTAIL.n133 9.3005
R750 VTAIL.n167 VTAIL.n166 9.3005
R751 VTAIL.n193 VTAIL.n192 9.3005
R752 VTAIL.n118 VTAIL.n117 9.3005
R753 VTAIL.n199 VTAIL.n198 9.3005
R754 VTAIL.n201 VTAIL.n200 9.3005
R755 VTAIL.n114 VTAIL.n113 9.3005
R756 VTAIL.n207 VTAIL.n206 9.3005
R757 VTAIL.n209 VTAIL.n208 9.3005
R758 VTAIL.n191 VTAIL.n190 9.3005
R759 VTAIL.n122 VTAIL.n121 9.3005
R760 VTAIL.n185 VTAIL.n184 9.3005
R761 VTAIL.n183 VTAIL.n182 9.3005
R762 VTAIL.n126 VTAIL.n125 9.3005
R763 VTAIL.n177 VTAIL.n176 9.3005
R764 VTAIL.n175 VTAIL.n174 9.3005
R765 VTAIL.n130 VTAIL.n129 9.3005
R766 VTAIL.n169 VTAIL.n168 9.3005
R767 VTAIL.n361 VTAIL.n350 8.92171
R768 VTAIL.n392 VTAIL.n334 8.92171
R769 VTAIL.n408 VTAIL.n407 8.92171
R770 VTAIL.n43 VTAIL.n32 8.92171
R771 VTAIL.n74 VTAIL.n16 8.92171
R772 VTAIL.n90 VTAIL.n89 8.92171
R773 VTAIL.n304 VTAIL.n303 8.92171
R774 VTAIL.n288 VTAIL.n230 8.92171
R775 VTAIL.n259 VTAIL.n248 8.92171
R776 VTAIL.n198 VTAIL.n197 8.92171
R777 VTAIL.n182 VTAIL.n124 8.92171
R778 VTAIL.n153 VTAIL.n142 8.92171
R779 VTAIL.n358 VTAIL.n357 8.14595
R780 VTAIL.n396 VTAIL.n395 8.14595
R781 VTAIL.n404 VTAIL.n328 8.14595
R782 VTAIL.n40 VTAIL.n39 8.14595
R783 VTAIL.n78 VTAIL.n77 8.14595
R784 VTAIL.n86 VTAIL.n10 8.14595
R785 VTAIL.n300 VTAIL.n224 8.14595
R786 VTAIL.n292 VTAIL.n291 8.14595
R787 VTAIL.n256 VTAIL.n255 8.14595
R788 VTAIL.n194 VTAIL.n118 8.14595
R789 VTAIL.n186 VTAIL.n185 8.14595
R790 VTAIL.n150 VTAIL.n149 8.14595
R791 VTAIL.n354 VTAIL.n352 7.3702
R792 VTAIL.n399 VTAIL.n332 7.3702
R793 VTAIL.n403 VTAIL.n330 7.3702
R794 VTAIL.n36 VTAIL.n34 7.3702
R795 VTAIL.n81 VTAIL.n14 7.3702
R796 VTAIL.n85 VTAIL.n12 7.3702
R797 VTAIL.n299 VTAIL.n226 7.3702
R798 VTAIL.n295 VTAIL.n228 7.3702
R799 VTAIL.n252 VTAIL.n250 7.3702
R800 VTAIL.n193 VTAIL.n120 7.3702
R801 VTAIL.n189 VTAIL.n122 7.3702
R802 VTAIL.n146 VTAIL.n144 7.3702
R803 VTAIL.n400 VTAIL.n399 6.59444
R804 VTAIL.n400 VTAIL.n330 6.59444
R805 VTAIL.n82 VTAIL.n81 6.59444
R806 VTAIL.n82 VTAIL.n12 6.59444
R807 VTAIL.n296 VTAIL.n226 6.59444
R808 VTAIL.n296 VTAIL.n295 6.59444
R809 VTAIL.n190 VTAIL.n120 6.59444
R810 VTAIL.n190 VTAIL.n189 6.59444
R811 VTAIL.n357 VTAIL.n352 5.81868
R812 VTAIL.n396 VTAIL.n332 5.81868
R813 VTAIL.n404 VTAIL.n403 5.81868
R814 VTAIL.n39 VTAIL.n34 5.81868
R815 VTAIL.n78 VTAIL.n14 5.81868
R816 VTAIL.n86 VTAIL.n85 5.81868
R817 VTAIL.n300 VTAIL.n299 5.81868
R818 VTAIL.n292 VTAIL.n228 5.81868
R819 VTAIL.n255 VTAIL.n250 5.81868
R820 VTAIL.n194 VTAIL.n193 5.81868
R821 VTAIL.n186 VTAIL.n122 5.81868
R822 VTAIL.n149 VTAIL.n144 5.81868
R823 VTAIL.n358 VTAIL.n350 5.04292
R824 VTAIL.n395 VTAIL.n334 5.04292
R825 VTAIL.n407 VTAIL.n328 5.04292
R826 VTAIL.n40 VTAIL.n32 5.04292
R827 VTAIL.n77 VTAIL.n16 5.04292
R828 VTAIL.n89 VTAIL.n10 5.04292
R829 VTAIL.n303 VTAIL.n224 5.04292
R830 VTAIL.n291 VTAIL.n230 5.04292
R831 VTAIL.n256 VTAIL.n248 5.04292
R832 VTAIL.n197 VTAIL.n118 5.04292
R833 VTAIL.n185 VTAIL.n124 5.04292
R834 VTAIL.n150 VTAIL.n142 5.04292
R835 VTAIL.n362 VTAIL.n361 4.26717
R836 VTAIL.n392 VTAIL.n391 4.26717
R837 VTAIL.n408 VTAIL.n326 4.26717
R838 VTAIL.n44 VTAIL.n43 4.26717
R839 VTAIL.n74 VTAIL.n73 4.26717
R840 VTAIL.n90 VTAIL.n8 4.26717
R841 VTAIL.n304 VTAIL.n222 4.26717
R842 VTAIL.n288 VTAIL.n287 4.26717
R843 VTAIL.n260 VTAIL.n259 4.26717
R844 VTAIL.n198 VTAIL.n116 4.26717
R845 VTAIL.n182 VTAIL.n181 4.26717
R846 VTAIL.n154 VTAIL.n153 4.26717
R847 VTAIL.n365 VTAIL.n348 3.49141
R848 VTAIL.n388 VTAIL.n336 3.49141
R849 VTAIL.n412 VTAIL.n411 3.49141
R850 VTAIL.n47 VTAIL.n30 3.49141
R851 VTAIL.n70 VTAIL.n18 3.49141
R852 VTAIL.n94 VTAIL.n93 3.49141
R853 VTAIL.n308 VTAIL.n307 3.49141
R854 VTAIL.n284 VTAIL.n232 3.49141
R855 VTAIL.n263 VTAIL.n246 3.49141
R856 VTAIL.n202 VTAIL.n201 3.49141
R857 VTAIL.n178 VTAIL.n126 3.49141
R858 VTAIL.n157 VTAIL.n140 3.49141
R859 VTAIL.n353 VTAIL.n351 2.84303
R860 VTAIL.n35 VTAIL.n33 2.84303
R861 VTAIL.n251 VTAIL.n249 2.84303
R862 VTAIL.n145 VTAIL.n143 2.84303
R863 VTAIL.n366 VTAIL.n346 2.71565
R864 VTAIL.n387 VTAIL.n338 2.71565
R865 VTAIL.n415 VTAIL.n324 2.71565
R866 VTAIL.n48 VTAIL.n28 2.71565
R867 VTAIL.n69 VTAIL.n20 2.71565
R868 VTAIL.n97 VTAIL.n6 2.71565
R869 VTAIL.n311 VTAIL.n220 2.71565
R870 VTAIL.n283 VTAIL.n234 2.71565
R871 VTAIL.n264 VTAIL.n244 2.71565
R872 VTAIL.n205 VTAIL.n114 2.71565
R873 VTAIL.n177 VTAIL.n128 2.71565
R874 VTAIL.n158 VTAIL.n138 2.71565
R875 VTAIL.n371 VTAIL.n369 1.93989
R876 VTAIL.n384 VTAIL.n383 1.93989
R877 VTAIL.n416 VTAIL.n322 1.93989
R878 VTAIL.n53 VTAIL.n51 1.93989
R879 VTAIL.n66 VTAIL.n65 1.93989
R880 VTAIL.n98 VTAIL.n4 1.93989
R881 VTAIL.n312 VTAIL.n218 1.93989
R882 VTAIL.n280 VTAIL.n279 1.93989
R883 VTAIL.n268 VTAIL.n267 1.93989
R884 VTAIL.n206 VTAIL.n112 1.93989
R885 VTAIL.n174 VTAIL.n173 1.93989
R886 VTAIL.n162 VTAIL.n161 1.93989
R887 VTAIL.n213 VTAIL.n109 1.62119
R888 VTAIL.n319 VTAIL.n215 1.62119
R889 VTAIL.n107 VTAIL.n105 1.62119
R890 VTAIL.n215 VTAIL.n213 1.28067
R891 VTAIL.n105 VTAIL.n1 1.28067
R892 VTAIL.n370 VTAIL.n344 1.16414
R893 VTAIL.n380 VTAIL.n340 1.16414
R894 VTAIL.n420 VTAIL.n419 1.16414
R895 VTAIL.n52 VTAIL.n26 1.16414
R896 VTAIL.n62 VTAIL.n22 1.16414
R897 VTAIL.n102 VTAIL.n101 1.16414
R898 VTAIL.n316 VTAIL.n315 1.16414
R899 VTAIL.n276 VTAIL.n236 1.16414
R900 VTAIL.n271 VTAIL.n241 1.16414
R901 VTAIL.n210 VTAIL.n209 1.16414
R902 VTAIL.n170 VTAIL.n130 1.16414
R903 VTAIL.n165 VTAIL.n135 1.16414
R904 VTAIL VTAIL.n423 1.15783
R905 VTAIL.n0 VTAIL.t1 1.05313
R906 VTAIL.n0 VTAIL.t4 1.05313
R907 VTAIL.n106 VTAIL.t9 1.05313
R908 VTAIL.n106 VTAIL.t10 1.05313
R909 VTAIL.n214 VTAIL.t8 1.05313
R910 VTAIL.n214 VTAIL.t11 1.05313
R911 VTAIL.n108 VTAIL.t2 1.05313
R912 VTAIL.n108 VTAIL.t3 1.05313
R913 VTAIL VTAIL.n1 0.463862
R914 VTAIL.n376 VTAIL.n375 0.388379
R915 VTAIL.n379 VTAIL.n342 0.388379
R916 VTAIL.n422 VTAIL.n320 0.388379
R917 VTAIL.n58 VTAIL.n57 0.388379
R918 VTAIL.n61 VTAIL.n24 0.388379
R919 VTAIL.n104 VTAIL.n2 0.388379
R920 VTAIL.n318 VTAIL.n216 0.388379
R921 VTAIL.n275 VTAIL.n238 0.388379
R922 VTAIL.n272 VTAIL.n240 0.388379
R923 VTAIL.n212 VTAIL.n110 0.388379
R924 VTAIL.n169 VTAIL.n132 0.388379
R925 VTAIL.n166 VTAIL.n134 0.388379
R926 VTAIL.n359 VTAIL.n351 0.155672
R927 VTAIL.n360 VTAIL.n359 0.155672
R928 VTAIL.n360 VTAIL.n347 0.155672
R929 VTAIL.n367 VTAIL.n347 0.155672
R930 VTAIL.n368 VTAIL.n367 0.155672
R931 VTAIL.n368 VTAIL.n343 0.155672
R932 VTAIL.n377 VTAIL.n343 0.155672
R933 VTAIL.n378 VTAIL.n377 0.155672
R934 VTAIL.n378 VTAIL.n339 0.155672
R935 VTAIL.n385 VTAIL.n339 0.155672
R936 VTAIL.n386 VTAIL.n385 0.155672
R937 VTAIL.n386 VTAIL.n335 0.155672
R938 VTAIL.n393 VTAIL.n335 0.155672
R939 VTAIL.n394 VTAIL.n393 0.155672
R940 VTAIL.n394 VTAIL.n331 0.155672
R941 VTAIL.n401 VTAIL.n331 0.155672
R942 VTAIL.n402 VTAIL.n401 0.155672
R943 VTAIL.n402 VTAIL.n327 0.155672
R944 VTAIL.n409 VTAIL.n327 0.155672
R945 VTAIL.n410 VTAIL.n409 0.155672
R946 VTAIL.n410 VTAIL.n323 0.155672
R947 VTAIL.n417 VTAIL.n323 0.155672
R948 VTAIL.n418 VTAIL.n417 0.155672
R949 VTAIL.n41 VTAIL.n33 0.155672
R950 VTAIL.n42 VTAIL.n41 0.155672
R951 VTAIL.n42 VTAIL.n29 0.155672
R952 VTAIL.n49 VTAIL.n29 0.155672
R953 VTAIL.n50 VTAIL.n49 0.155672
R954 VTAIL.n50 VTAIL.n25 0.155672
R955 VTAIL.n59 VTAIL.n25 0.155672
R956 VTAIL.n60 VTAIL.n59 0.155672
R957 VTAIL.n60 VTAIL.n21 0.155672
R958 VTAIL.n67 VTAIL.n21 0.155672
R959 VTAIL.n68 VTAIL.n67 0.155672
R960 VTAIL.n68 VTAIL.n17 0.155672
R961 VTAIL.n75 VTAIL.n17 0.155672
R962 VTAIL.n76 VTAIL.n75 0.155672
R963 VTAIL.n76 VTAIL.n13 0.155672
R964 VTAIL.n83 VTAIL.n13 0.155672
R965 VTAIL.n84 VTAIL.n83 0.155672
R966 VTAIL.n84 VTAIL.n9 0.155672
R967 VTAIL.n91 VTAIL.n9 0.155672
R968 VTAIL.n92 VTAIL.n91 0.155672
R969 VTAIL.n92 VTAIL.n5 0.155672
R970 VTAIL.n99 VTAIL.n5 0.155672
R971 VTAIL.n100 VTAIL.n99 0.155672
R972 VTAIL.n314 VTAIL.n313 0.155672
R973 VTAIL.n313 VTAIL.n219 0.155672
R974 VTAIL.n306 VTAIL.n219 0.155672
R975 VTAIL.n306 VTAIL.n305 0.155672
R976 VTAIL.n305 VTAIL.n223 0.155672
R977 VTAIL.n298 VTAIL.n223 0.155672
R978 VTAIL.n298 VTAIL.n297 0.155672
R979 VTAIL.n297 VTAIL.n227 0.155672
R980 VTAIL.n290 VTAIL.n227 0.155672
R981 VTAIL.n290 VTAIL.n289 0.155672
R982 VTAIL.n289 VTAIL.n231 0.155672
R983 VTAIL.n282 VTAIL.n231 0.155672
R984 VTAIL.n282 VTAIL.n281 0.155672
R985 VTAIL.n281 VTAIL.n235 0.155672
R986 VTAIL.n274 VTAIL.n235 0.155672
R987 VTAIL.n274 VTAIL.n273 0.155672
R988 VTAIL.n273 VTAIL.n239 0.155672
R989 VTAIL.n266 VTAIL.n239 0.155672
R990 VTAIL.n266 VTAIL.n265 0.155672
R991 VTAIL.n265 VTAIL.n245 0.155672
R992 VTAIL.n258 VTAIL.n245 0.155672
R993 VTAIL.n258 VTAIL.n257 0.155672
R994 VTAIL.n257 VTAIL.n249 0.155672
R995 VTAIL.n208 VTAIL.n207 0.155672
R996 VTAIL.n207 VTAIL.n113 0.155672
R997 VTAIL.n200 VTAIL.n113 0.155672
R998 VTAIL.n200 VTAIL.n199 0.155672
R999 VTAIL.n199 VTAIL.n117 0.155672
R1000 VTAIL.n192 VTAIL.n117 0.155672
R1001 VTAIL.n192 VTAIL.n191 0.155672
R1002 VTAIL.n191 VTAIL.n121 0.155672
R1003 VTAIL.n184 VTAIL.n121 0.155672
R1004 VTAIL.n184 VTAIL.n183 0.155672
R1005 VTAIL.n183 VTAIL.n125 0.155672
R1006 VTAIL.n176 VTAIL.n125 0.155672
R1007 VTAIL.n176 VTAIL.n175 0.155672
R1008 VTAIL.n175 VTAIL.n129 0.155672
R1009 VTAIL.n168 VTAIL.n129 0.155672
R1010 VTAIL.n168 VTAIL.n167 0.155672
R1011 VTAIL.n167 VTAIL.n133 0.155672
R1012 VTAIL.n160 VTAIL.n133 0.155672
R1013 VTAIL.n160 VTAIL.n159 0.155672
R1014 VTAIL.n159 VTAIL.n139 0.155672
R1015 VTAIL.n152 VTAIL.n139 0.155672
R1016 VTAIL.n152 VTAIL.n151 0.155672
R1017 VTAIL.n151 VTAIL.n143 0.155672
R1018 B.n654 B.n653 585
R1019 B.n654 B.n57 585
R1020 B.n657 B.n656 585
R1021 B.n658 B.n128 585
R1022 B.n660 B.n659 585
R1023 B.n662 B.n127 585
R1024 B.n665 B.n664 585
R1025 B.n666 B.n126 585
R1026 B.n668 B.n667 585
R1027 B.n670 B.n125 585
R1028 B.n673 B.n672 585
R1029 B.n674 B.n124 585
R1030 B.n676 B.n675 585
R1031 B.n678 B.n123 585
R1032 B.n681 B.n680 585
R1033 B.n682 B.n122 585
R1034 B.n684 B.n683 585
R1035 B.n686 B.n121 585
R1036 B.n689 B.n688 585
R1037 B.n690 B.n120 585
R1038 B.n692 B.n691 585
R1039 B.n694 B.n119 585
R1040 B.n697 B.n696 585
R1041 B.n698 B.n118 585
R1042 B.n700 B.n699 585
R1043 B.n702 B.n117 585
R1044 B.n705 B.n704 585
R1045 B.n706 B.n116 585
R1046 B.n708 B.n707 585
R1047 B.n710 B.n115 585
R1048 B.n713 B.n712 585
R1049 B.n714 B.n114 585
R1050 B.n716 B.n715 585
R1051 B.n718 B.n113 585
R1052 B.n721 B.n720 585
R1053 B.n722 B.n112 585
R1054 B.n724 B.n723 585
R1055 B.n726 B.n111 585
R1056 B.n729 B.n728 585
R1057 B.n730 B.n110 585
R1058 B.n732 B.n731 585
R1059 B.n734 B.n109 585
R1060 B.n737 B.n736 585
R1061 B.n738 B.n108 585
R1062 B.n740 B.n739 585
R1063 B.n742 B.n107 585
R1064 B.n745 B.n744 585
R1065 B.n746 B.n106 585
R1066 B.n748 B.n747 585
R1067 B.n750 B.n105 585
R1068 B.n753 B.n752 585
R1069 B.n754 B.n104 585
R1070 B.n756 B.n755 585
R1071 B.n758 B.n103 585
R1072 B.n761 B.n760 585
R1073 B.n762 B.n102 585
R1074 B.n764 B.n763 585
R1075 B.n766 B.n101 585
R1076 B.n769 B.n768 585
R1077 B.n770 B.n100 585
R1078 B.n772 B.n771 585
R1079 B.n774 B.n99 585
R1080 B.n777 B.n776 585
R1081 B.n779 B.n96 585
R1082 B.n781 B.n780 585
R1083 B.n783 B.n95 585
R1084 B.n786 B.n785 585
R1085 B.n787 B.n94 585
R1086 B.n789 B.n788 585
R1087 B.n791 B.n93 585
R1088 B.n793 B.n792 585
R1089 B.n795 B.n794 585
R1090 B.n798 B.n797 585
R1091 B.n799 B.n88 585
R1092 B.n801 B.n800 585
R1093 B.n803 B.n87 585
R1094 B.n806 B.n805 585
R1095 B.n807 B.n86 585
R1096 B.n809 B.n808 585
R1097 B.n811 B.n85 585
R1098 B.n814 B.n813 585
R1099 B.n815 B.n84 585
R1100 B.n817 B.n816 585
R1101 B.n819 B.n83 585
R1102 B.n822 B.n821 585
R1103 B.n823 B.n82 585
R1104 B.n825 B.n824 585
R1105 B.n827 B.n81 585
R1106 B.n830 B.n829 585
R1107 B.n831 B.n80 585
R1108 B.n833 B.n832 585
R1109 B.n835 B.n79 585
R1110 B.n838 B.n837 585
R1111 B.n839 B.n78 585
R1112 B.n841 B.n840 585
R1113 B.n843 B.n77 585
R1114 B.n846 B.n845 585
R1115 B.n847 B.n76 585
R1116 B.n849 B.n848 585
R1117 B.n851 B.n75 585
R1118 B.n854 B.n853 585
R1119 B.n855 B.n74 585
R1120 B.n857 B.n856 585
R1121 B.n859 B.n73 585
R1122 B.n862 B.n861 585
R1123 B.n863 B.n72 585
R1124 B.n865 B.n864 585
R1125 B.n867 B.n71 585
R1126 B.n870 B.n869 585
R1127 B.n871 B.n70 585
R1128 B.n873 B.n872 585
R1129 B.n875 B.n69 585
R1130 B.n878 B.n877 585
R1131 B.n879 B.n68 585
R1132 B.n881 B.n880 585
R1133 B.n883 B.n67 585
R1134 B.n886 B.n885 585
R1135 B.n887 B.n66 585
R1136 B.n889 B.n888 585
R1137 B.n891 B.n65 585
R1138 B.n894 B.n893 585
R1139 B.n895 B.n64 585
R1140 B.n897 B.n896 585
R1141 B.n899 B.n63 585
R1142 B.n902 B.n901 585
R1143 B.n903 B.n62 585
R1144 B.n905 B.n904 585
R1145 B.n907 B.n61 585
R1146 B.n910 B.n909 585
R1147 B.n911 B.n60 585
R1148 B.n913 B.n912 585
R1149 B.n915 B.n59 585
R1150 B.n918 B.n917 585
R1151 B.n919 B.n58 585
R1152 B.n652 B.n56 585
R1153 B.n922 B.n56 585
R1154 B.n651 B.n55 585
R1155 B.n923 B.n55 585
R1156 B.n650 B.n54 585
R1157 B.n924 B.n54 585
R1158 B.n649 B.n648 585
R1159 B.n648 B.n50 585
R1160 B.n647 B.n49 585
R1161 B.n930 B.n49 585
R1162 B.n646 B.n48 585
R1163 B.n931 B.n48 585
R1164 B.n645 B.n47 585
R1165 B.n932 B.n47 585
R1166 B.n644 B.n643 585
R1167 B.n643 B.n43 585
R1168 B.n642 B.n42 585
R1169 B.n938 B.n42 585
R1170 B.n641 B.n41 585
R1171 B.n939 B.n41 585
R1172 B.n640 B.n40 585
R1173 B.n940 B.n40 585
R1174 B.n639 B.n638 585
R1175 B.n638 B.n36 585
R1176 B.n637 B.n35 585
R1177 B.n946 B.n35 585
R1178 B.n636 B.n34 585
R1179 B.n947 B.n34 585
R1180 B.n635 B.n33 585
R1181 B.n948 B.n33 585
R1182 B.n634 B.n633 585
R1183 B.n633 B.n29 585
R1184 B.n632 B.n28 585
R1185 B.n954 B.n28 585
R1186 B.n631 B.n27 585
R1187 B.n955 B.n27 585
R1188 B.n630 B.n26 585
R1189 B.n956 B.n26 585
R1190 B.n629 B.n628 585
R1191 B.n628 B.n22 585
R1192 B.n627 B.n21 585
R1193 B.n962 B.n21 585
R1194 B.n626 B.n20 585
R1195 B.n963 B.n20 585
R1196 B.n625 B.n19 585
R1197 B.n964 B.n19 585
R1198 B.n624 B.n623 585
R1199 B.n623 B.n15 585
R1200 B.n622 B.n14 585
R1201 B.n970 B.n14 585
R1202 B.n621 B.n13 585
R1203 B.n971 B.n13 585
R1204 B.n620 B.n12 585
R1205 B.n972 B.n12 585
R1206 B.n619 B.n618 585
R1207 B.n618 B.n8 585
R1208 B.n617 B.n7 585
R1209 B.n978 B.n7 585
R1210 B.n616 B.n6 585
R1211 B.n979 B.n6 585
R1212 B.n615 B.n5 585
R1213 B.n980 B.n5 585
R1214 B.n614 B.n613 585
R1215 B.n613 B.n4 585
R1216 B.n612 B.n129 585
R1217 B.n612 B.n611 585
R1218 B.n602 B.n130 585
R1219 B.n131 B.n130 585
R1220 B.n604 B.n603 585
R1221 B.n605 B.n604 585
R1222 B.n601 B.n135 585
R1223 B.n139 B.n135 585
R1224 B.n600 B.n599 585
R1225 B.n599 B.n598 585
R1226 B.n137 B.n136 585
R1227 B.n138 B.n137 585
R1228 B.n591 B.n590 585
R1229 B.n592 B.n591 585
R1230 B.n589 B.n144 585
R1231 B.n144 B.n143 585
R1232 B.n588 B.n587 585
R1233 B.n587 B.n586 585
R1234 B.n146 B.n145 585
R1235 B.n147 B.n146 585
R1236 B.n579 B.n578 585
R1237 B.n580 B.n579 585
R1238 B.n577 B.n152 585
R1239 B.n152 B.n151 585
R1240 B.n576 B.n575 585
R1241 B.n575 B.n574 585
R1242 B.n154 B.n153 585
R1243 B.n155 B.n154 585
R1244 B.n567 B.n566 585
R1245 B.n568 B.n567 585
R1246 B.n565 B.n160 585
R1247 B.n160 B.n159 585
R1248 B.n564 B.n563 585
R1249 B.n563 B.n562 585
R1250 B.n162 B.n161 585
R1251 B.n163 B.n162 585
R1252 B.n555 B.n554 585
R1253 B.n556 B.n555 585
R1254 B.n553 B.n168 585
R1255 B.n168 B.n167 585
R1256 B.n552 B.n551 585
R1257 B.n551 B.n550 585
R1258 B.n170 B.n169 585
R1259 B.n171 B.n170 585
R1260 B.n543 B.n542 585
R1261 B.n544 B.n543 585
R1262 B.n541 B.n175 585
R1263 B.n179 B.n175 585
R1264 B.n540 B.n539 585
R1265 B.n539 B.n538 585
R1266 B.n177 B.n176 585
R1267 B.n178 B.n177 585
R1268 B.n531 B.n530 585
R1269 B.n532 B.n531 585
R1270 B.n529 B.n184 585
R1271 B.n184 B.n183 585
R1272 B.n528 B.n527 585
R1273 B.n527 B.n526 585
R1274 B.n523 B.n188 585
R1275 B.n522 B.n521 585
R1276 B.n519 B.n189 585
R1277 B.n519 B.n187 585
R1278 B.n518 B.n517 585
R1279 B.n516 B.n515 585
R1280 B.n514 B.n191 585
R1281 B.n512 B.n511 585
R1282 B.n510 B.n192 585
R1283 B.n509 B.n508 585
R1284 B.n506 B.n193 585
R1285 B.n504 B.n503 585
R1286 B.n502 B.n194 585
R1287 B.n501 B.n500 585
R1288 B.n498 B.n195 585
R1289 B.n496 B.n495 585
R1290 B.n494 B.n196 585
R1291 B.n493 B.n492 585
R1292 B.n490 B.n197 585
R1293 B.n488 B.n487 585
R1294 B.n486 B.n198 585
R1295 B.n485 B.n484 585
R1296 B.n482 B.n199 585
R1297 B.n480 B.n479 585
R1298 B.n478 B.n200 585
R1299 B.n477 B.n476 585
R1300 B.n474 B.n201 585
R1301 B.n472 B.n471 585
R1302 B.n470 B.n202 585
R1303 B.n469 B.n468 585
R1304 B.n466 B.n203 585
R1305 B.n464 B.n463 585
R1306 B.n462 B.n204 585
R1307 B.n461 B.n460 585
R1308 B.n458 B.n205 585
R1309 B.n456 B.n455 585
R1310 B.n454 B.n206 585
R1311 B.n453 B.n452 585
R1312 B.n450 B.n207 585
R1313 B.n448 B.n447 585
R1314 B.n446 B.n208 585
R1315 B.n445 B.n444 585
R1316 B.n442 B.n209 585
R1317 B.n440 B.n439 585
R1318 B.n438 B.n210 585
R1319 B.n437 B.n436 585
R1320 B.n434 B.n211 585
R1321 B.n432 B.n431 585
R1322 B.n430 B.n212 585
R1323 B.n429 B.n428 585
R1324 B.n426 B.n213 585
R1325 B.n424 B.n423 585
R1326 B.n422 B.n214 585
R1327 B.n421 B.n420 585
R1328 B.n418 B.n215 585
R1329 B.n416 B.n415 585
R1330 B.n414 B.n216 585
R1331 B.n413 B.n412 585
R1332 B.n410 B.n217 585
R1333 B.n408 B.n407 585
R1334 B.n406 B.n218 585
R1335 B.n405 B.n404 585
R1336 B.n402 B.n219 585
R1337 B.n400 B.n399 585
R1338 B.n398 B.n220 585
R1339 B.n397 B.n396 585
R1340 B.n394 B.n224 585
R1341 B.n392 B.n391 585
R1342 B.n390 B.n225 585
R1343 B.n389 B.n388 585
R1344 B.n386 B.n226 585
R1345 B.n384 B.n383 585
R1346 B.n381 B.n227 585
R1347 B.n380 B.n379 585
R1348 B.n377 B.n230 585
R1349 B.n375 B.n374 585
R1350 B.n373 B.n231 585
R1351 B.n372 B.n371 585
R1352 B.n369 B.n232 585
R1353 B.n367 B.n366 585
R1354 B.n365 B.n233 585
R1355 B.n364 B.n363 585
R1356 B.n361 B.n234 585
R1357 B.n359 B.n358 585
R1358 B.n357 B.n235 585
R1359 B.n356 B.n355 585
R1360 B.n353 B.n236 585
R1361 B.n351 B.n350 585
R1362 B.n349 B.n237 585
R1363 B.n348 B.n347 585
R1364 B.n345 B.n238 585
R1365 B.n343 B.n342 585
R1366 B.n341 B.n239 585
R1367 B.n340 B.n339 585
R1368 B.n337 B.n240 585
R1369 B.n335 B.n334 585
R1370 B.n333 B.n241 585
R1371 B.n332 B.n331 585
R1372 B.n329 B.n242 585
R1373 B.n327 B.n326 585
R1374 B.n325 B.n243 585
R1375 B.n324 B.n323 585
R1376 B.n321 B.n244 585
R1377 B.n319 B.n318 585
R1378 B.n317 B.n245 585
R1379 B.n316 B.n315 585
R1380 B.n313 B.n246 585
R1381 B.n311 B.n310 585
R1382 B.n309 B.n247 585
R1383 B.n308 B.n307 585
R1384 B.n305 B.n248 585
R1385 B.n303 B.n302 585
R1386 B.n301 B.n249 585
R1387 B.n300 B.n299 585
R1388 B.n297 B.n250 585
R1389 B.n295 B.n294 585
R1390 B.n293 B.n251 585
R1391 B.n292 B.n291 585
R1392 B.n289 B.n252 585
R1393 B.n287 B.n286 585
R1394 B.n285 B.n253 585
R1395 B.n284 B.n283 585
R1396 B.n281 B.n254 585
R1397 B.n279 B.n278 585
R1398 B.n277 B.n255 585
R1399 B.n276 B.n275 585
R1400 B.n273 B.n256 585
R1401 B.n271 B.n270 585
R1402 B.n269 B.n257 585
R1403 B.n268 B.n267 585
R1404 B.n265 B.n258 585
R1405 B.n263 B.n262 585
R1406 B.n261 B.n260 585
R1407 B.n186 B.n185 585
R1408 B.n525 B.n524 585
R1409 B.n526 B.n525 585
R1410 B.n182 B.n181 585
R1411 B.n183 B.n182 585
R1412 B.n534 B.n533 585
R1413 B.n533 B.n532 585
R1414 B.n535 B.n180 585
R1415 B.n180 B.n178 585
R1416 B.n537 B.n536 585
R1417 B.n538 B.n537 585
R1418 B.n174 B.n173 585
R1419 B.n179 B.n174 585
R1420 B.n546 B.n545 585
R1421 B.n545 B.n544 585
R1422 B.n547 B.n172 585
R1423 B.n172 B.n171 585
R1424 B.n549 B.n548 585
R1425 B.n550 B.n549 585
R1426 B.n166 B.n165 585
R1427 B.n167 B.n166 585
R1428 B.n558 B.n557 585
R1429 B.n557 B.n556 585
R1430 B.n559 B.n164 585
R1431 B.n164 B.n163 585
R1432 B.n561 B.n560 585
R1433 B.n562 B.n561 585
R1434 B.n158 B.n157 585
R1435 B.n159 B.n158 585
R1436 B.n570 B.n569 585
R1437 B.n569 B.n568 585
R1438 B.n571 B.n156 585
R1439 B.n156 B.n155 585
R1440 B.n573 B.n572 585
R1441 B.n574 B.n573 585
R1442 B.n150 B.n149 585
R1443 B.n151 B.n150 585
R1444 B.n582 B.n581 585
R1445 B.n581 B.n580 585
R1446 B.n583 B.n148 585
R1447 B.n148 B.n147 585
R1448 B.n585 B.n584 585
R1449 B.n586 B.n585 585
R1450 B.n142 B.n141 585
R1451 B.n143 B.n142 585
R1452 B.n594 B.n593 585
R1453 B.n593 B.n592 585
R1454 B.n595 B.n140 585
R1455 B.n140 B.n138 585
R1456 B.n597 B.n596 585
R1457 B.n598 B.n597 585
R1458 B.n134 B.n133 585
R1459 B.n139 B.n134 585
R1460 B.n607 B.n606 585
R1461 B.n606 B.n605 585
R1462 B.n608 B.n132 585
R1463 B.n132 B.n131 585
R1464 B.n610 B.n609 585
R1465 B.n611 B.n610 585
R1466 B.n2 B.n0 585
R1467 B.n4 B.n2 585
R1468 B.n3 B.n1 585
R1469 B.n979 B.n3 585
R1470 B.n977 B.n976 585
R1471 B.n978 B.n977 585
R1472 B.n975 B.n9 585
R1473 B.n9 B.n8 585
R1474 B.n974 B.n973 585
R1475 B.n973 B.n972 585
R1476 B.n11 B.n10 585
R1477 B.n971 B.n11 585
R1478 B.n969 B.n968 585
R1479 B.n970 B.n969 585
R1480 B.n967 B.n16 585
R1481 B.n16 B.n15 585
R1482 B.n966 B.n965 585
R1483 B.n965 B.n964 585
R1484 B.n18 B.n17 585
R1485 B.n963 B.n18 585
R1486 B.n961 B.n960 585
R1487 B.n962 B.n961 585
R1488 B.n959 B.n23 585
R1489 B.n23 B.n22 585
R1490 B.n958 B.n957 585
R1491 B.n957 B.n956 585
R1492 B.n25 B.n24 585
R1493 B.n955 B.n25 585
R1494 B.n953 B.n952 585
R1495 B.n954 B.n953 585
R1496 B.n951 B.n30 585
R1497 B.n30 B.n29 585
R1498 B.n950 B.n949 585
R1499 B.n949 B.n948 585
R1500 B.n32 B.n31 585
R1501 B.n947 B.n32 585
R1502 B.n945 B.n944 585
R1503 B.n946 B.n945 585
R1504 B.n943 B.n37 585
R1505 B.n37 B.n36 585
R1506 B.n942 B.n941 585
R1507 B.n941 B.n940 585
R1508 B.n39 B.n38 585
R1509 B.n939 B.n39 585
R1510 B.n937 B.n936 585
R1511 B.n938 B.n937 585
R1512 B.n935 B.n44 585
R1513 B.n44 B.n43 585
R1514 B.n934 B.n933 585
R1515 B.n933 B.n932 585
R1516 B.n46 B.n45 585
R1517 B.n931 B.n46 585
R1518 B.n929 B.n928 585
R1519 B.n930 B.n929 585
R1520 B.n927 B.n51 585
R1521 B.n51 B.n50 585
R1522 B.n926 B.n925 585
R1523 B.n925 B.n924 585
R1524 B.n53 B.n52 585
R1525 B.n923 B.n53 585
R1526 B.n921 B.n920 585
R1527 B.n922 B.n921 585
R1528 B.n982 B.n981 585
R1529 B.n981 B.n980 585
R1530 B.n525 B.n188 526.135
R1531 B.n921 B.n58 526.135
R1532 B.n527 B.n186 526.135
R1533 B.n654 B.n56 526.135
R1534 B.n228 B.t14 498.087
R1535 B.n221 B.t6 498.087
R1536 B.n89 B.t10 498.087
R1537 B.n97 B.t17 498.087
R1538 B.n228 B.t16 435.786
R1539 B.n221 B.t9 435.786
R1540 B.n89 B.t12 435.786
R1541 B.n97 B.t18 435.786
R1542 B.n229 B.t15 399.327
R1543 B.n98 B.t19 399.327
R1544 B.n222 B.t8 399.327
R1545 B.n90 B.t13 399.327
R1546 B.n655 B.n57 256.663
R1547 B.n661 B.n57 256.663
R1548 B.n663 B.n57 256.663
R1549 B.n669 B.n57 256.663
R1550 B.n671 B.n57 256.663
R1551 B.n677 B.n57 256.663
R1552 B.n679 B.n57 256.663
R1553 B.n685 B.n57 256.663
R1554 B.n687 B.n57 256.663
R1555 B.n693 B.n57 256.663
R1556 B.n695 B.n57 256.663
R1557 B.n701 B.n57 256.663
R1558 B.n703 B.n57 256.663
R1559 B.n709 B.n57 256.663
R1560 B.n711 B.n57 256.663
R1561 B.n717 B.n57 256.663
R1562 B.n719 B.n57 256.663
R1563 B.n725 B.n57 256.663
R1564 B.n727 B.n57 256.663
R1565 B.n733 B.n57 256.663
R1566 B.n735 B.n57 256.663
R1567 B.n741 B.n57 256.663
R1568 B.n743 B.n57 256.663
R1569 B.n749 B.n57 256.663
R1570 B.n751 B.n57 256.663
R1571 B.n757 B.n57 256.663
R1572 B.n759 B.n57 256.663
R1573 B.n765 B.n57 256.663
R1574 B.n767 B.n57 256.663
R1575 B.n773 B.n57 256.663
R1576 B.n775 B.n57 256.663
R1577 B.n782 B.n57 256.663
R1578 B.n784 B.n57 256.663
R1579 B.n790 B.n57 256.663
R1580 B.n92 B.n57 256.663
R1581 B.n796 B.n57 256.663
R1582 B.n802 B.n57 256.663
R1583 B.n804 B.n57 256.663
R1584 B.n810 B.n57 256.663
R1585 B.n812 B.n57 256.663
R1586 B.n818 B.n57 256.663
R1587 B.n820 B.n57 256.663
R1588 B.n826 B.n57 256.663
R1589 B.n828 B.n57 256.663
R1590 B.n834 B.n57 256.663
R1591 B.n836 B.n57 256.663
R1592 B.n842 B.n57 256.663
R1593 B.n844 B.n57 256.663
R1594 B.n850 B.n57 256.663
R1595 B.n852 B.n57 256.663
R1596 B.n858 B.n57 256.663
R1597 B.n860 B.n57 256.663
R1598 B.n866 B.n57 256.663
R1599 B.n868 B.n57 256.663
R1600 B.n874 B.n57 256.663
R1601 B.n876 B.n57 256.663
R1602 B.n882 B.n57 256.663
R1603 B.n884 B.n57 256.663
R1604 B.n890 B.n57 256.663
R1605 B.n892 B.n57 256.663
R1606 B.n898 B.n57 256.663
R1607 B.n900 B.n57 256.663
R1608 B.n906 B.n57 256.663
R1609 B.n908 B.n57 256.663
R1610 B.n914 B.n57 256.663
R1611 B.n916 B.n57 256.663
R1612 B.n520 B.n187 256.663
R1613 B.n190 B.n187 256.663
R1614 B.n513 B.n187 256.663
R1615 B.n507 B.n187 256.663
R1616 B.n505 B.n187 256.663
R1617 B.n499 B.n187 256.663
R1618 B.n497 B.n187 256.663
R1619 B.n491 B.n187 256.663
R1620 B.n489 B.n187 256.663
R1621 B.n483 B.n187 256.663
R1622 B.n481 B.n187 256.663
R1623 B.n475 B.n187 256.663
R1624 B.n473 B.n187 256.663
R1625 B.n467 B.n187 256.663
R1626 B.n465 B.n187 256.663
R1627 B.n459 B.n187 256.663
R1628 B.n457 B.n187 256.663
R1629 B.n451 B.n187 256.663
R1630 B.n449 B.n187 256.663
R1631 B.n443 B.n187 256.663
R1632 B.n441 B.n187 256.663
R1633 B.n435 B.n187 256.663
R1634 B.n433 B.n187 256.663
R1635 B.n427 B.n187 256.663
R1636 B.n425 B.n187 256.663
R1637 B.n419 B.n187 256.663
R1638 B.n417 B.n187 256.663
R1639 B.n411 B.n187 256.663
R1640 B.n409 B.n187 256.663
R1641 B.n403 B.n187 256.663
R1642 B.n401 B.n187 256.663
R1643 B.n395 B.n187 256.663
R1644 B.n393 B.n187 256.663
R1645 B.n387 B.n187 256.663
R1646 B.n385 B.n187 256.663
R1647 B.n378 B.n187 256.663
R1648 B.n376 B.n187 256.663
R1649 B.n370 B.n187 256.663
R1650 B.n368 B.n187 256.663
R1651 B.n362 B.n187 256.663
R1652 B.n360 B.n187 256.663
R1653 B.n354 B.n187 256.663
R1654 B.n352 B.n187 256.663
R1655 B.n346 B.n187 256.663
R1656 B.n344 B.n187 256.663
R1657 B.n338 B.n187 256.663
R1658 B.n336 B.n187 256.663
R1659 B.n330 B.n187 256.663
R1660 B.n328 B.n187 256.663
R1661 B.n322 B.n187 256.663
R1662 B.n320 B.n187 256.663
R1663 B.n314 B.n187 256.663
R1664 B.n312 B.n187 256.663
R1665 B.n306 B.n187 256.663
R1666 B.n304 B.n187 256.663
R1667 B.n298 B.n187 256.663
R1668 B.n296 B.n187 256.663
R1669 B.n290 B.n187 256.663
R1670 B.n288 B.n187 256.663
R1671 B.n282 B.n187 256.663
R1672 B.n280 B.n187 256.663
R1673 B.n274 B.n187 256.663
R1674 B.n272 B.n187 256.663
R1675 B.n266 B.n187 256.663
R1676 B.n264 B.n187 256.663
R1677 B.n259 B.n187 256.663
R1678 B.n525 B.n182 163.367
R1679 B.n533 B.n182 163.367
R1680 B.n533 B.n180 163.367
R1681 B.n537 B.n180 163.367
R1682 B.n537 B.n174 163.367
R1683 B.n545 B.n174 163.367
R1684 B.n545 B.n172 163.367
R1685 B.n549 B.n172 163.367
R1686 B.n549 B.n166 163.367
R1687 B.n557 B.n166 163.367
R1688 B.n557 B.n164 163.367
R1689 B.n561 B.n164 163.367
R1690 B.n561 B.n158 163.367
R1691 B.n569 B.n158 163.367
R1692 B.n569 B.n156 163.367
R1693 B.n573 B.n156 163.367
R1694 B.n573 B.n150 163.367
R1695 B.n581 B.n150 163.367
R1696 B.n581 B.n148 163.367
R1697 B.n585 B.n148 163.367
R1698 B.n585 B.n142 163.367
R1699 B.n593 B.n142 163.367
R1700 B.n593 B.n140 163.367
R1701 B.n597 B.n140 163.367
R1702 B.n597 B.n134 163.367
R1703 B.n606 B.n134 163.367
R1704 B.n606 B.n132 163.367
R1705 B.n610 B.n132 163.367
R1706 B.n610 B.n2 163.367
R1707 B.n981 B.n2 163.367
R1708 B.n981 B.n3 163.367
R1709 B.n977 B.n3 163.367
R1710 B.n977 B.n9 163.367
R1711 B.n973 B.n9 163.367
R1712 B.n973 B.n11 163.367
R1713 B.n969 B.n11 163.367
R1714 B.n969 B.n16 163.367
R1715 B.n965 B.n16 163.367
R1716 B.n965 B.n18 163.367
R1717 B.n961 B.n18 163.367
R1718 B.n961 B.n23 163.367
R1719 B.n957 B.n23 163.367
R1720 B.n957 B.n25 163.367
R1721 B.n953 B.n25 163.367
R1722 B.n953 B.n30 163.367
R1723 B.n949 B.n30 163.367
R1724 B.n949 B.n32 163.367
R1725 B.n945 B.n32 163.367
R1726 B.n945 B.n37 163.367
R1727 B.n941 B.n37 163.367
R1728 B.n941 B.n39 163.367
R1729 B.n937 B.n39 163.367
R1730 B.n937 B.n44 163.367
R1731 B.n933 B.n44 163.367
R1732 B.n933 B.n46 163.367
R1733 B.n929 B.n46 163.367
R1734 B.n929 B.n51 163.367
R1735 B.n925 B.n51 163.367
R1736 B.n925 B.n53 163.367
R1737 B.n921 B.n53 163.367
R1738 B.n521 B.n519 163.367
R1739 B.n519 B.n518 163.367
R1740 B.n515 B.n514 163.367
R1741 B.n512 B.n192 163.367
R1742 B.n508 B.n506 163.367
R1743 B.n504 B.n194 163.367
R1744 B.n500 B.n498 163.367
R1745 B.n496 B.n196 163.367
R1746 B.n492 B.n490 163.367
R1747 B.n488 B.n198 163.367
R1748 B.n484 B.n482 163.367
R1749 B.n480 B.n200 163.367
R1750 B.n476 B.n474 163.367
R1751 B.n472 B.n202 163.367
R1752 B.n468 B.n466 163.367
R1753 B.n464 B.n204 163.367
R1754 B.n460 B.n458 163.367
R1755 B.n456 B.n206 163.367
R1756 B.n452 B.n450 163.367
R1757 B.n448 B.n208 163.367
R1758 B.n444 B.n442 163.367
R1759 B.n440 B.n210 163.367
R1760 B.n436 B.n434 163.367
R1761 B.n432 B.n212 163.367
R1762 B.n428 B.n426 163.367
R1763 B.n424 B.n214 163.367
R1764 B.n420 B.n418 163.367
R1765 B.n416 B.n216 163.367
R1766 B.n412 B.n410 163.367
R1767 B.n408 B.n218 163.367
R1768 B.n404 B.n402 163.367
R1769 B.n400 B.n220 163.367
R1770 B.n396 B.n394 163.367
R1771 B.n392 B.n225 163.367
R1772 B.n388 B.n386 163.367
R1773 B.n384 B.n227 163.367
R1774 B.n379 B.n377 163.367
R1775 B.n375 B.n231 163.367
R1776 B.n371 B.n369 163.367
R1777 B.n367 B.n233 163.367
R1778 B.n363 B.n361 163.367
R1779 B.n359 B.n235 163.367
R1780 B.n355 B.n353 163.367
R1781 B.n351 B.n237 163.367
R1782 B.n347 B.n345 163.367
R1783 B.n343 B.n239 163.367
R1784 B.n339 B.n337 163.367
R1785 B.n335 B.n241 163.367
R1786 B.n331 B.n329 163.367
R1787 B.n327 B.n243 163.367
R1788 B.n323 B.n321 163.367
R1789 B.n319 B.n245 163.367
R1790 B.n315 B.n313 163.367
R1791 B.n311 B.n247 163.367
R1792 B.n307 B.n305 163.367
R1793 B.n303 B.n249 163.367
R1794 B.n299 B.n297 163.367
R1795 B.n295 B.n251 163.367
R1796 B.n291 B.n289 163.367
R1797 B.n287 B.n253 163.367
R1798 B.n283 B.n281 163.367
R1799 B.n279 B.n255 163.367
R1800 B.n275 B.n273 163.367
R1801 B.n271 B.n257 163.367
R1802 B.n267 B.n265 163.367
R1803 B.n263 B.n260 163.367
R1804 B.n527 B.n184 163.367
R1805 B.n531 B.n184 163.367
R1806 B.n531 B.n177 163.367
R1807 B.n539 B.n177 163.367
R1808 B.n539 B.n175 163.367
R1809 B.n543 B.n175 163.367
R1810 B.n543 B.n170 163.367
R1811 B.n551 B.n170 163.367
R1812 B.n551 B.n168 163.367
R1813 B.n555 B.n168 163.367
R1814 B.n555 B.n162 163.367
R1815 B.n563 B.n162 163.367
R1816 B.n563 B.n160 163.367
R1817 B.n567 B.n160 163.367
R1818 B.n567 B.n154 163.367
R1819 B.n575 B.n154 163.367
R1820 B.n575 B.n152 163.367
R1821 B.n579 B.n152 163.367
R1822 B.n579 B.n146 163.367
R1823 B.n587 B.n146 163.367
R1824 B.n587 B.n144 163.367
R1825 B.n591 B.n144 163.367
R1826 B.n591 B.n137 163.367
R1827 B.n599 B.n137 163.367
R1828 B.n599 B.n135 163.367
R1829 B.n604 B.n135 163.367
R1830 B.n604 B.n130 163.367
R1831 B.n612 B.n130 163.367
R1832 B.n613 B.n612 163.367
R1833 B.n613 B.n5 163.367
R1834 B.n6 B.n5 163.367
R1835 B.n7 B.n6 163.367
R1836 B.n618 B.n7 163.367
R1837 B.n618 B.n12 163.367
R1838 B.n13 B.n12 163.367
R1839 B.n14 B.n13 163.367
R1840 B.n623 B.n14 163.367
R1841 B.n623 B.n19 163.367
R1842 B.n20 B.n19 163.367
R1843 B.n21 B.n20 163.367
R1844 B.n628 B.n21 163.367
R1845 B.n628 B.n26 163.367
R1846 B.n27 B.n26 163.367
R1847 B.n28 B.n27 163.367
R1848 B.n633 B.n28 163.367
R1849 B.n633 B.n33 163.367
R1850 B.n34 B.n33 163.367
R1851 B.n35 B.n34 163.367
R1852 B.n638 B.n35 163.367
R1853 B.n638 B.n40 163.367
R1854 B.n41 B.n40 163.367
R1855 B.n42 B.n41 163.367
R1856 B.n643 B.n42 163.367
R1857 B.n643 B.n47 163.367
R1858 B.n48 B.n47 163.367
R1859 B.n49 B.n48 163.367
R1860 B.n648 B.n49 163.367
R1861 B.n648 B.n54 163.367
R1862 B.n55 B.n54 163.367
R1863 B.n56 B.n55 163.367
R1864 B.n917 B.n915 163.367
R1865 B.n913 B.n60 163.367
R1866 B.n909 B.n907 163.367
R1867 B.n905 B.n62 163.367
R1868 B.n901 B.n899 163.367
R1869 B.n897 B.n64 163.367
R1870 B.n893 B.n891 163.367
R1871 B.n889 B.n66 163.367
R1872 B.n885 B.n883 163.367
R1873 B.n881 B.n68 163.367
R1874 B.n877 B.n875 163.367
R1875 B.n873 B.n70 163.367
R1876 B.n869 B.n867 163.367
R1877 B.n865 B.n72 163.367
R1878 B.n861 B.n859 163.367
R1879 B.n857 B.n74 163.367
R1880 B.n853 B.n851 163.367
R1881 B.n849 B.n76 163.367
R1882 B.n845 B.n843 163.367
R1883 B.n841 B.n78 163.367
R1884 B.n837 B.n835 163.367
R1885 B.n833 B.n80 163.367
R1886 B.n829 B.n827 163.367
R1887 B.n825 B.n82 163.367
R1888 B.n821 B.n819 163.367
R1889 B.n817 B.n84 163.367
R1890 B.n813 B.n811 163.367
R1891 B.n809 B.n86 163.367
R1892 B.n805 B.n803 163.367
R1893 B.n801 B.n88 163.367
R1894 B.n797 B.n795 163.367
R1895 B.n792 B.n791 163.367
R1896 B.n789 B.n94 163.367
R1897 B.n785 B.n783 163.367
R1898 B.n781 B.n96 163.367
R1899 B.n776 B.n774 163.367
R1900 B.n772 B.n100 163.367
R1901 B.n768 B.n766 163.367
R1902 B.n764 B.n102 163.367
R1903 B.n760 B.n758 163.367
R1904 B.n756 B.n104 163.367
R1905 B.n752 B.n750 163.367
R1906 B.n748 B.n106 163.367
R1907 B.n744 B.n742 163.367
R1908 B.n740 B.n108 163.367
R1909 B.n736 B.n734 163.367
R1910 B.n732 B.n110 163.367
R1911 B.n728 B.n726 163.367
R1912 B.n724 B.n112 163.367
R1913 B.n720 B.n718 163.367
R1914 B.n716 B.n114 163.367
R1915 B.n712 B.n710 163.367
R1916 B.n708 B.n116 163.367
R1917 B.n704 B.n702 163.367
R1918 B.n700 B.n118 163.367
R1919 B.n696 B.n694 163.367
R1920 B.n692 B.n120 163.367
R1921 B.n688 B.n686 163.367
R1922 B.n684 B.n122 163.367
R1923 B.n680 B.n678 163.367
R1924 B.n676 B.n124 163.367
R1925 B.n672 B.n670 163.367
R1926 B.n668 B.n126 163.367
R1927 B.n664 B.n662 163.367
R1928 B.n660 B.n128 163.367
R1929 B.n656 B.n654 163.367
R1930 B.n520 B.n188 71.676
R1931 B.n518 B.n190 71.676
R1932 B.n514 B.n513 71.676
R1933 B.n507 B.n192 71.676
R1934 B.n506 B.n505 71.676
R1935 B.n499 B.n194 71.676
R1936 B.n498 B.n497 71.676
R1937 B.n491 B.n196 71.676
R1938 B.n490 B.n489 71.676
R1939 B.n483 B.n198 71.676
R1940 B.n482 B.n481 71.676
R1941 B.n475 B.n200 71.676
R1942 B.n474 B.n473 71.676
R1943 B.n467 B.n202 71.676
R1944 B.n466 B.n465 71.676
R1945 B.n459 B.n204 71.676
R1946 B.n458 B.n457 71.676
R1947 B.n451 B.n206 71.676
R1948 B.n450 B.n449 71.676
R1949 B.n443 B.n208 71.676
R1950 B.n442 B.n441 71.676
R1951 B.n435 B.n210 71.676
R1952 B.n434 B.n433 71.676
R1953 B.n427 B.n212 71.676
R1954 B.n426 B.n425 71.676
R1955 B.n419 B.n214 71.676
R1956 B.n418 B.n417 71.676
R1957 B.n411 B.n216 71.676
R1958 B.n410 B.n409 71.676
R1959 B.n403 B.n218 71.676
R1960 B.n402 B.n401 71.676
R1961 B.n395 B.n220 71.676
R1962 B.n394 B.n393 71.676
R1963 B.n387 B.n225 71.676
R1964 B.n386 B.n385 71.676
R1965 B.n378 B.n227 71.676
R1966 B.n377 B.n376 71.676
R1967 B.n370 B.n231 71.676
R1968 B.n369 B.n368 71.676
R1969 B.n362 B.n233 71.676
R1970 B.n361 B.n360 71.676
R1971 B.n354 B.n235 71.676
R1972 B.n353 B.n352 71.676
R1973 B.n346 B.n237 71.676
R1974 B.n345 B.n344 71.676
R1975 B.n338 B.n239 71.676
R1976 B.n337 B.n336 71.676
R1977 B.n330 B.n241 71.676
R1978 B.n329 B.n328 71.676
R1979 B.n322 B.n243 71.676
R1980 B.n321 B.n320 71.676
R1981 B.n314 B.n245 71.676
R1982 B.n313 B.n312 71.676
R1983 B.n306 B.n247 71.676
R1984 B.n305 B.n304 71.676
R1985 B.n298 B.n249 71.676
R1986 B.n297 B.n296 71.676
R1987 B.n290 B.n251 71.676
R1988 B.n289 B.n288 71.676
R1989 B.n282 B.n253 71.676
R1990 B.n281 B.n280 71.676
R1991 B.n274 B.n255 71.676
R1992 B.n273 B.n272 71.676
R1993 B.n266 B.n257 71.676
R1994 B.n265 B.n264 71.676
R1995 B.n260 B.n259 71.676
R1996 B.n916 B.n58 71.676
R1997 B.n915 B.n914 71.676
R1998 B.n908 B.n60 71.676
R1999 B.n907 B.n906 71.676
R2000 B.n900 B.n62 71.676
R2001 B.n899 B.n898 71.676
R2002 B.n892 B.n64 71.676
R2003 B.n891 B.n890 71.676
R2004 B.n884 B.n66 71.676
R2005 B.n883 B.n882 71.676
R2006 B.n876 B.n68 71.676
R2007 B.n875 B.n874 71.676
R2008 B.n868 B.n70 71.676
R2009 B.n867 B.n866 71.676
R2010 B.n860 B.n72 71.676
R2011 B.n859 B.n858 71.676
R2012 B.n852 B.n74 71.676
R2013 B.n851 B.n850 71.676
R2014 B.n844 B.n76 71.676
R2015 B.n843 B.n842 71.676
R2016 B.n836 B.n78 71.676
R2017 B.n835 B.n834 71.676
R2018 B.n828 B.n80 71.676
R2019 B.n827 B.n826 71.676
R2020 B.n820 B.n82 71.676
R2021 B.n819 B.n818 71.676
R2022 B.n812 B.n84 71.676
R2023 B.n811 B.n810 71.676
R2024 B.n804 B.n86 71.676
R2025 B.n803 B.n802 71.676
R2026 B.n796 B.n88 71.676
R2027 B.n795 B.n92 71.676
R2028 B.n791 B.n790 71.676
R2029 B.n784 B.n94 71.676
R2030 B.n783 B.n782 71.676
R2031 B.n775 B.n96 71.676
R2032 B.n774 B.n773 71.676
R2033 B.n767 B.n100 71.676
R2034 B.n766 B.n765 71.676
R2035 B.n759 B.n102 71.676
R2036 B.n758 B.n757 71.676
R2037 B.n751 B.n104 71.676
R2038 B.n750 B.n749 71.676
R2039 B.n743 B.n106 71.676
R2040 B.n742 B.n741 71.676
R2041 B.n735 B.n108 71.676
R2042 B.n734 B.n733 71.676
R2043 B.n727 B.n110 71.676
R2044 B.n726 B.n725 71.676
R2045 B.n719 B.n112 71.676
R2046 B.n718 B.n717 71.676
R2047 B.n711 B.n114 71.676
R2048 B.n710 B.n709 71.676
R2049 B.n703 B.n116 71.676
R2050 B.n702 B.n701 71.676
R2051 B.n695 B.n118 71.676
R2052 B.n694 B.n693 71.676
R2053 B.n687 B.n120 71.676
R2054 B.n686 B.n685 71.676
R2055 B.n679 B.n122 71.676
R2056 B.n678 B.n677 71.676
R2057 B.n671 B.n124 71.676
R2058 B.n670 B.n669 71.676
R2059 B.n663 B.n126 71.676
R2060 B.n662 B.n661 71.676
R2061 B.n655 B.n128 71.676
R2062 B.n656 B.n655 71.676
R2063 B.n661 B.n660 71.676
R2064 B.n664 B.n663 71.676
R2065 B.n669 B.n668 71.676
R2066 B.n672 B.n671 71.676
R2067 B.n677 B.n676 71.676
R2068 B.n680 B.n679 71.676
R2069 B.n685 B.n684 71.676
R2070 B.n688 B.n687 71.676
R2071 B.n693 B.n692 71.676
R2072 B.n696 B.n695 71.676
R2073 B.n701 B.n700 71.676
R2074 B.n704 B.n703 71.676
R2075 B.n709 B.n708 71.676
R2076 B.n712 B.n711 71.676
R2077 B.n717 B.n716 71.676
R2078 B.n720 B.n719 71.676
R2079 B.n725 B.n724 71.676
R2080 B.n728 B.n727 71.676
R2081 B.n733 B.n732 71.676
R2082 B.n736 B.n735 71.676
R2083 B.n741 B.n740 71.676
R2084 B.n744 B.n743 71.676
R2085 B.n749 B.n748 71.676
R2086 B.n752 B.n751 71.676
R2087 B.n757 B.n756 71.676
R2088 B.n760 B.n759 71.676
R2089 B.n765 B.n764 71.676
R2090 B.n768 B.n767 71.676
R2091 B.n773 B.n772 71.676
R2092 B.n776 B.n775 71.676
R2093 B.n782 B.n781 71.676
R2094 B.n785 B.n784 71.676
R2095 B.n790 B.n789 71.676
R2096 B.n792 B.n92 71.676
R2097 B.n797 B.n796 71.676
R2098 B.n802 B.n801 71.676
R2099 B.n805 B.n804 71.676
R2100 B.n810 B.n809 71.676
R2101 B.n813 B.n812 71.676
R2102 B.n818 B.n817 71.676
R2103 B.n821 B.n820 71.676
R2104 B.n826 B.n825 71.676
R2105 B.n829 B.n828 71.676
R2106 B.n834 B.n833 71.676
R2107 B.n837 B.n836 71.676
R2108 B.n842 B.n841 71.676
R2109 B.n845 B.n844 71.676
R2110 B.n850 B.n849 71.676
R2111 B.n853 B.n852 71.676
R2112 B.n858 B.n857 71.676
R2113 B.n861 B.n860 71.676
R2114 B.n866 B.n865 71.676
R2115 B.n869 B.n868 71.676
R2116 B.n874 B.n873 71.676
R2117 B.n877 B.n876 71.676
R2118 B.n882 B.n881 71.676
R2119 B.n885 B.n884 71.676
R2120 B.n890 B.n889 71.676
R2121 B.n893 B.n892 71.676
R2122 B.n898 B.n897 71.676
R2123 B.n901 B.n900 71.676
R2124 B.n906 B.n905 71.676
R2125 B.n909 B.n908 71.676
R2126 B.n914 B.n913 71.676
R2127 B.n917 B.n916 71.676
R2128 B.n521 B.n520 71.676
R2129 B.n515 B.n190 71.676
R2130 B.n513 B.n512 71.676
R2131 B.n508 B.n507 71.676
R2132 B.n505 B.n504 71.676
R2133 B.n500 B.n499 71.676
R2134 B.n497 B.n496 71.676
R2135 B.n492 B.n491 71.676
R2136 B.n489 B.n488 71.676
R2137 B.n484 B.n483 71.676
R2138 B.n481 B.n480 71.676
R2139 B.n476 B.n475 71.676
R2140 B.n473 B.n472 71.676
R2141 B.n468 B.n467 71.676
R2142 B.n465 B.n464 71.676
R2143 B.n460 B.n459 71.676
R2144 B.n457 B.n456 71.676
R2145 B.n452 B.n451 71.676
R2146 B.n449 B.n448 71.676
R2147 B.n444 B.n443 71.676
R2148 B.n441 B.n440 71.676
R2149 B.n436 B.n435 71.676
R2150 B.n433 B.n432 71.676
R2151 B.n428 B.n427 71.676
R2152 B.n425 B.n424 71.676
R2153 B.n420 B.n419 71.676
R2154 B.n417 B.n416 71.676
R2155 B.n412 B.n411 71.676
R2156 B.n409 B.n408 71.676
R2157 B.n404 B.n403 71.676
R2158 B.n401 B.n400 71.676
R2159 B.n396 B.n395 71.676
R2160 B.n393 B.n392 71.676
R2161 B.n388 B.n387 71.676
R2162 B.n385 B.n384 71.676
R2163 B.n379 B.n378 71.676
R2164 B.n376 B.n375 71.676
R2165 B.n371 B.n370 71.676
R2166 B.n368 B.n367 71.676
R2167 B.n363 B.n362 71.676
R2168 B.n360 B.n359 71.676
R2169 B.n355 B.n354 71.676
R2170 B.n352 B.n351 71.676
R2171 B.n347 B.n346 71.676
R2172 B.n344 B.n343 71.676
R2173 B.n339 B.n338 71.676
R2174 B.n336 B.n335 71.676
R2175 B.n331 B.n330 71.676
R2176 B.n328 B.n327 71.676
R2177 B.n323 B.n322 71.676
R2178 B.n320 B.n319 71.676
R2179 B.n315 B.n314 71.676
R2180 B.n312 B.n311 71.676
R2181 B.n307 B.n306 71.676
R2182 B.n304 B.n303 71.676
R2183 B.n299 B.n298 71.676
R2184 B.n296 B.n295 71.676
R2185 B.n291 B.n290 71.676
R2186 B.n288 B.n287 71.676
R2187 B.n283 B.n282 71.676
R2188 B.n280 B.n279 71.676
R2189 B.n275 B.n274 71.676
R2190 B.n272 B.n271 71.676
R2191 B.n267 B.n266 71.676
R2192 B.n264 B.n263 71.676
R2193 B.n259 B.n186 71.676
R2194 B.n526 B.n187 63.484
R2195 B.n922 B.n57 63.484
R2196 B.n382 B.n229 59.5399
R2197 B.n223 B.n222 59.5399
R2198 B.n91 B.n90 59.5399
R2199 B.n778 B.n98 59.5399
R2200 B.n229 B.n228 36.4611
R2201 B.n222 B.n221 36.4611
R2202 B.n90 B.n89 36.4611
R2203 B.n98 B.n97 36.4611
R2204 B.n920 B.n919 34.1859
R2205 B.n653 B.n652 34.1859
R2206 B.n528 B.n185 34.1859
R2207 B.n524 B.n523 34.1859
R2208 B.n526 B.n183 31.0572
R2209 B.n532 B.n183 31.0572
R2210 B.n532 B.n178 31.0572
R2211 B.n538 B.n178 31.0572
R2212 B.n538 B.n179 31.0572
R2213 B.n544 B.n171 31.0572
R2214 B.n550 B.n171 31.0572
R2215 B.n550 B.n167 31.0572
R2216 B.n556 B.n167 31.0572
R2217 B.n556 B.n163 31.0572
R2218 B.n562 B.n163 31.0572
R2219 B.n562 B.n159 31.0572
R2220 B.n568 B.n159 31.0572
R2221 B.n574 B.n155 31.0572
R2222 B.n574 B.n151 31.0572
R2223 B.n580 B.n151 31.0572
R2224 B.n580 B.n147 31.0572
R2225 B.n586 B.n147 31.0572
R2226 B.n592 B.n143 31.0572
R2227 B.n592 B.n138 31.0572
R2228 B.n598 B.n138 31.0572
R2229 B.n598 B.n139 31.0572
R2230 B.n605 B.n131 31.0572
R2231 B.n611 B.n131 31.0572
R2232 B.n611 B.n4 31.0572
R2233 B.n980 B.n4 31.0572
R2234 B.n980 B.n979 31.0572
R2235 B.n979 B.n978 31.0572
R2236 B.n978 B.n8 31.0572
R2237 B.n972 B.n8 31.0572
R2238 B.n971 B.n970 31.0572
R2239 B.n970 B.n15 31.0572
R2240 B.n964 B.n15 31.0572
R2241 B.n964 B.n963 31.0572
R2242 B.n962 B.n22 31.0572
R2243 B.n956 B.n22 31.0572
R2244 B.n956 B.n955 31.0572
R2245 B.n955 B.n954 31.0572
R2246 B.n954 B.n29 31.0572
R2247 B.n948 B.n947 31.0572
R2248 B.n947 B.n946 31.0572
R2249 B.n946 B.n36 31.0572
R2250 B.n940 B.n36 31.0572
R2251 B.n940 B.n939 31.0572
R2252 B.n939 B.n938 31.0572
R2253 B.n938 B.n43 31.0572
R2254 B.n932 B.n43 31.0572
R2255 B.n931 B.n930 31.0572
R2256 B.n930 B.n50 31.0572
R2257 B.n924 B.n50 31.0572
R2258 B.n924 B.n923 31.0572
R2259 B.n923 B.n922 31.0572
R2260 B.t3 B.n143 27.8602
R2261 B.n963 B.t4 27.8602
R2262 B.n179 B.t7 26.0333
R2263 B.t11 B.n931 26.0333
R2264 B.n139 B.t0 19.6393
R2265 B.t1 B.n971 19.6393
R2266 B B.n982 18.0485
R2267 B.n568 B.t2 17.8124
R2268 B.n948 B.t5 17.8124
R2269 B.t2 B.n155 13.2453
R2270 B.t5 B.n29 13.2453
R2271 B.n605 B.t0 11.4184
R2272 B.n972 B.t1 11.4184
R2273 B.n919 B.n918 10.6151
R2274 B.n918 B.n59 10.6151
R2275 B.n912 B.n59 10.6151
R2276 B.n912 B.n911 10.6151
R2277 B.n911 B.n910 10.6151
R2278 B.n910 B.n61 10.6151
R2279 B.n904 B.n61 10.6151
R2280 B.n904 B.n903 10.6151
R2281 B.n903 B.n902 10.6151
R2282 B.n902 B.n63 10.6151
R2283 B.n896 B.n63 10.6151
R2284 B.n896 B.n895 10.6151
R2285 B.n895 B.n894 10.6151
R2286 B.n894 B.n65 10.6151
R2287 B.n888 B.n65 10.6151
R2288 B.n888 B.n887 10.6151
R2289 B.n887 B.n886 10.6151
R2290 B.n886 B.n67 10.6151
R2291 B.n880 B.n67 10.6151
R2292 B.n880 B.n879 10.6151
R2293 B.n879 B.n878 10.6151
R2294 B.n878 B.n69 10.6151
R2295 B.n872 B.n69 10.6151
R2296 B.n872 B.n871 10.6151
R2297 B.n871 B.n870 10.6151
R2298 B.n870 B.n71 10.6151
R2299 B.n864 B.n71 10.6151
R2300 B.n864 B.n863 10.6151
R2301 B.n863 B.n862 10.6151
R2302 B.n862 B.n73 10.6151
R2303 B.n856 B.n73 10.6151
R2304 B.n856 B.n855 10.6151
R2305 B.n855 B.n854 10.6151
R2306 B.n854 B.n75 10.6151
R2307 B.n848 B.n75 10.6151
R2308 B.n848 B.n847 10.6151
R2309 B.n847 B.n846 10.6151
R2310 B.n846 B.n77 10.6151
R2311 B.n840 B.n77 10.6151
R2312 B.n840 B.n839 10.6151
R2313 B.n839 B.n838 10.6151
R2314 B.n838 B.n79 10.6151
R2315 B.n832 B.n79 10.6151
R2316 B.n832 B.n831 10.6151
R2317 B.n831 B.n830 10.6151
R2318 B.n830 B.n81 10.6151
R2319 B.n824 B.n81 10.6151
R2320 B.n824 B.n823 10.6151
R2321 B.n823 B.n822 10.6151
R2322 B.n822 B.n83 10.6151
R2323 B.n816 B.n83 10.6151
R2324 B.n816 B.n815 10.6151
R2325 B.n815 B.n814 10.6151
R2326 B.n814 B.n85 10.6151
R2327 B.n808 B.n85 10.6151
R2328 B.n808 B.n807 10.6151
R2329 B.n807 B.n806 10.6151
R2330 B.n806 B.n87 10.6151
R2331 B.n800 B.n87 10.6151
R2332 B.n800 B.n799 10.6151
R2333 B.n799 B.n798 10.6151
R2334 B.n794 B.n793 10.6151
R2335 B.n793 B.n93 10.6151
R2336 B.n788 B.n93 10.6151
R2337 B.n788 B.n787 10.6151
R2338 B.n787 B.n786 10.6151
R2339 B.n786 B.n95 10.6151
R2340 B.n780 B.n95 10.6151
R2341 B.n780 B.n779 10.6151
R2342 B.n777 B.n99 10.6151
R2343 B.n771 B.n99 10.6151
R2344 B.n771 B.n770 10.6151
R2345 B.n770 B.n769 10.6151
R2346 B.n769 B.n101 10.6151
R2347 B.n763 B.n101 10.6151
R2348 B.n763 B.n762 10.6151
R2349 B.n762 B.n761 10.6151
R2350 B.n761 B.n103 10.6151
R2351 B.n755 B.n103 10.6151
R2352 B.n755 B.n754 10.6151
R2353 B.n754 B.n753 10.6151
R2354 B.n753 B.n105 10.6151
R2355 B.n747 B.n105 10.6151
R2356 B.n747 B.n746 10.6151
R2357 B.n746 B.n745 10.6151
R2358 B.n745 B.n107 10.6151
R2359 B.n739 B.n107 10.6151
R2360 B.n739 B.n738 10.6151
R2361 B.n738 B.n737 10.6151
R2362 B.n737 B.n109 10.6151
R2363 B.n731 B.n109 10.6151
R2364 B.n731 B.n730 10.6151
R2365 B.n730 B.n729 10.6151
R2366 B.n729 B.n111 10.6151
R2367 B.n723 B.n111 10.6151
R2368 B.n723 B.n722 10.6151
R2369 B.n722 B.n721 10.6151
R2370 B.n721 B.n113 10.6151
R2371 B.n715 B.n113 10.6151
R2372 B.n715 B.n714 10.6151
R2373 B.n714 B.n713 10.6151
R2374 B.n713 B.n115 10.6151
R2375 B.n707 B.n115 10.6151
R2376 B.n707 B.n706 10.6151
R2377 B.n706 B.n705 10.6151
R2378 B.n705 B.n117 10.6151
R2379 B.n699 B.n117 10.6151
R2380 B.n699 B.n698 10.6151
R2381 B.n698 B.n697 10.6151
R2382 B.n697 B.n119 10.6151
R2383 B.n691 B.n119 10.6151
R2384 B.n691 B.n690 10.6151
R2385 B.n690 B.n689 10.6151
R2386 B.n689 B.n121 10.6151
R2387 B.n683 B.n121 10.6151
R2388 B.n683 B.n682 10.6151
R2389 B.n682 B.n681 10.6151
R2390 B.n681 B.n123 10.6151
R2391 B.n675 B.n123 10.6151
R2392 B.n675 B.n674 10.6151
R2393 B.n674 B.n673 10.6151
R2394 B.n673 B.n125 10.6151
R2395 B.n667 B.n125 10.6151
R2396 B.n667 B.n666 10.6151
R2397 B.n666 B.n665 10.6151
R2398 B.n665 B.n127 10.6151
R2399 B.n659 B.n127 10.6151
R2400 B.n659 B.n658 10.6151
R2401 B.n658 B.n657 10.6151
R2402 B.n657 B.n653 10.6151
R2403 B.n529 B.n528 10.6151
R2404 B.n530 B.n529 10.6151
R2405 B.n530 B.n176 10.6151
R2406 B.n540 B.n176 10.6151
R2407 B.n541 B.n540 10.6151
R2408 B.n542 B.n541 10.6151
R2409 B.n542 B.n169 10.6151
R2410 B.n552 B.n169 10.6151
R2411 B.n553 B.n552 10.6151
R2412 B.n554 B.n553 10.6151
R2413 B.n554 B.n161 10.6151
R2414 B.n564 B.n161 10.6151
R2415 B.n565 B.n564 10.6151
R2416 B.n566 B.n565 10.6151
R2417 B.n566 B.n153 10.6151
R2418 B.n576 B.n153 10.6151
R2419 B.n577 B.n576 10.6151
R2420 B.n578 B.n577 10.6151
R2421 B.n578 B.n145 10.6151
R2422 B.n588 B.n145 10.6151
R2423 B.n589 B.n588 10.6151
R2424 B.n590 B.n589 10.6151
R2425 B.n590 B.n136 10.6151
R2426 B.n600 B.n136 10.6151
R2427 B.n601 B.n600 10.6151
R2428 B.n603 B.n601 10.6151
R2429 B.n603 B.n602 10.6151
R2430 B.n602 B.n129 10.6151
R2431 B.n614 B.n129 10.6151
R2432 B.n615 B.n614 10.6151
R2433 B.n616 B.n615 10.6151
R2434 B.n617 B.n616 10.6151
R2435 B.n619 B.n617 10.6151
R2436 B.n620 B.n619 10.6151
R2437 B.n621 B.n620 10.6151
R2438 B.n622 B.n621 10.6151
R2439 B.n624 B.n622 10.6151
R2440 B.n625 B.n624 10.6151
R2441 B.n626 B.n625 10.6151
R2442 B.n627 B.n626 10.6151
R2443 B.n629 B.n627 10.6151
R2444 B.n630 B.n629 10.6151
R2445 B.n631 B.n630 10.6151
R2446 B.n632 B.n631 10.6151
R2447 B.n634 B.n632 10.6151
R2448 B.n635 B.n634 10.6151
R2449 B.n636 B.n635 10.6151
R2450 B.n637 B.n636 10.6151
R2451 B.n639 B.n637 10.6151
R2452 B.n640 B.n639 10.6151
R2453 B.n641 B.n640 10.6151
R2454 B.n642 B.n641 10.6151
R2455 B.n644 B.n642 10.6151
R2456 B.n645 B.n644 10.6151
R2457 B.n646 B.n645 10.6151
R2458 B.n647 B.n646 10.6151
R2459 B.n649 B.n647 10.6151
R2460 B.n650 B.n649 10.6151
R2461 B.n651 B.n650 10.6151
R2462 B.n652 B.n651 10.6151
R2463 B.n523 B.n522 10.6151
R2464 B.n522 B.n189 10.6151
R2465 B.n517 B.n189 10.6151
R2466 B.n517 B.n516 10.6151
R2467 B.n516 B.n191 10.6151
R2468 B.n511 B.n191 10.6151
R2469 B.n511 B.n510 10.6151
R2470 B.n510 B.n509 10.6151
R2471 B.n509 B.n193 10.6151
R2472 B.n503 B.n193 10.6151
R2473 B.n503 B.n502 10.6151
R2474 B.n502 B.n501 10.6151
R2475 B.n501 B.n195 10.6151
R2476 B.n495 B.n195 10.6151
R2477 B.n495 B.n494 10.6151
R2478 B.n494 B.n493 10.6151
R2479 B.n493 B.n197 10.6151
R2480 B.n487 B.n197 10.6151
R2481 B.n487 B.n486 10.6151
R2482 B.n486 B.n485 10.6151
R2483 B.n485 B.n199 10.6151
R2484 B.n479 B.n199 10.6151
R2485 B.n479 B.n478 10.6151
R2486 B.n478 B.n477 10.6151
R2487 B.n477 B.n201 10.6151
R2488 B.n471 B.n201 10.6151
R2489 B.n471 B.n470 10.6151
R2490 B.n470 B.n469 10.6151
R2491 B.n469 B.n203 10.6151
R2492 B.n463 B.n203 10.6151
R2493 B.n463 B.n462 10.6151
R2494 B.n462 B.n461 10.6151
R2495 B.n461 B.n205 10.6151
R2496 B.n455 B.n205 10.6151
R2497 B.n455 B.n454 10.6151
R2498 B.n454 B.n453 10.6151
R2499 B.n453 B.n207 10.6151
R2500 B.n447 B.n207 10.6151
R2501 B.n447 B.n446 10.6151
R2502 B.n446 B.n445 10.6151
R2503 B.n445 B.n209 10.6151
R2504 B.n439 B.n209 10.6151
R2505 B.n439 B.n438 10.6151
R2506 B.n438 B.n437 10.6151
R2507 B.n437 B.n211 10.6151
R2508 B.n431 B.n211 10.6151
R2509 B.n431 B.n430 10.6151
R2510 B.n430 B.n429 10.6151
R2511 B.n429 B.n213 10.6151
R2512 B.n423 B.n213 10.6151
R2513 B.n423 B.n422 10.6151
R2514 B.n422 B.n421 10.6151
R2515 B.n421 B.n215 10.6151
R2516 B.n415 B.n215 10.6151
R2517 B.n415 B.n414 10.6151
R2518 B.n414 B.n413 10.6151
R2519 B.n413 B.n217 10.6151
R2520 B.n407 B.n217 10.6151
R2521 B.n407 B.n406 10.6151
R2522 B.n406 B.n405 10.6151
R2523 B.n405 B.n219 10.6151
R2524 B.n399 B.n398 10.6151
R2525 B.n398 B.n397 10.6151
R2526 B.n397 B.n224 10.6151
R2527 B.n391 B.n224 10.6151
R2528 B.n391 B.n390 10.6151
R2529 B.n390 B.n389 10.6151
R2530 B.n389 B.n226 10.6151
R2531 B.n383 B.n226 10.6151
R2532 B.n381 B.n380 10.6151
R2533 B.n380 B.n230 10.6151
R2534 B.n374 B.n230 10.6151
R2535 B.n374 B.n373 10.6151
R2536 B.n373 B.n372 10.6151
R2537 B.n372 B.n232 10.6151
R2538 B.n366 B.n232 10.6151
R2539 B.n366 B.n365 10.6151
R2540 B.n365 B.n364 10.6151
R2541 B.n364 B.n234 10.6151
R2542 B.n358 B.n234 10.6151
R2543 B.n358 B.n357 10.6151
R2544 B.n357 B.n356 10.6151
R2545 B.n356 B.n236 10.6151
R2546 B.n350 B.n236 10.6151
R2547 B.n350 B.n349 10.6151
R2548 B.n349 B.n348 10.6151
R2549 B.n348 B.n238 10.6151
R2550 B.n342 B.n238 10.6151
R2551 B.n342 B.n341 10.6151
R2552 B.n341 B.n340 10.6151
R2553 B.n340 B.n240 10.6151
R2554 B.n334 B.n240 10.6151
R2555 B.n334 B.n333 10.6151
R2556 B.n333 B.n332 10.6151
R2557 B.n332 B.n242 10.6151
R2558 B.n326 B.n242 10.6151
R2559 B.n326 B.n325 10.6151
R2560 B.n325 B.n324 10.6151
R2561 B.n324 B.n244 10.6151
R2562 B.n318 B.n244 10.6151
R2563 B.n318 B.n317 10.6151
R2564 B.n317 B.n316 10.6151
R2565 B.n316 B.n246 10.6151
R2566 B.n310 B.n246 10.6151
R2567 B.n310 B.n309 10.6151
R2568 B.n309 B.n308 10.6151
R2569 B.n308 B.n248 10.6151
R2570 B.n302 B.n248 10.6151
R2571 B.n302 B.n301 10.6151
R2572 B.n301 B.n300 10.6151
R2573 B.n300 B.n250 10.6151
R2574 B.n294 B.n250 10.6151
R2575 B.n294 B.n293 10.6151
R2576 B.n293 B.n292 10.6151
R2577 B.n292 B.n252 10.6151
R2578 B.n286 B.n252 10.6151
R2579 B.n286 B.n285 10.6151
R2580 B.n285 B.n284 10.6151
R2581 B.n284 B.n254 10.6151
R2582 B.n278 B.n254 10.6151
R2583 B.n278 B.n277 10.6151
R2584 B.n277 B.n276 10.6151
R2585 B.n276 B.n256 10.6151
R2586 B.n270 B.n256 10.6151
R2587 B.n270 B.n269 10.6151
R2588 B.n269 B.n268 10.6151
R2589 B.n268 B.n258 10.6151
R2590 B.n262 B.n258 10.6151
R2591 B.n262 B.n261 10.6151
R2592 B.n261 B.n185 10.6151
R2593 B.n524 B.n181 10.6151
R2594 B.n534 B.n181 10.6151
R2595 B.n535 B.n534 10.6151
R2596 B.n536 B.n535 10.6151
R2597 B.n536 B.n173 10.6151
R2598 B.n546 B.n173 10.6151
R2599 B.n547 B.n546 10.6151
R2600 B.n548 B.n547 10.6151
R2601 B.n548 B.n165 10.6151
R2602 B.n558 B.n165 10.6151
R2603 B.n559 B.n558 10.6151
R2604 B.n560 B.n559 10.6151
R2605 B.n560 B.n157 10.6151
R2606 B.n570 B.n157 10.6151
R2607 B.n571 B.n570 10.6151
R2608 B.n572 B.n571 10.6151
R2609 B.n572 B.n149 10.6151
R2610 B.n582 B.n149 10.6151
R2611 B.n583 B.n582 10.6151
R2612 B.n584 B.n583 10.6151
R2613 B.n584 B.n141 10.6151
R2614 B.n594 B.n141 10.6151
R2615 B.n595 B.n594 10.6151
R2616 B.n596 B.n595 10.6151
R2617 B.n596 B.n133 10.6151
R2618 B.n607 B.n133 10.6151
R2619 B.n608 B.n607 10.6151
R2620 B.n609 B.n608 10.6151
R2621 B.n609 B.n0 10.6151
R2622 B.n976 B.n1 10.6151
R2623 B.n976 B.n975 10.6151
R2624 B.n975 B.n974 10.6151
R2625 B.n974 B.n10 10.6151
R2626 B.n968 B.n10 10.6151
R2627 B.n968 B.n967 10.6151
R2628 B.n967 B.n966 10.6151
R2629 B.n966 B.n17 10.6151
R2630 B.n960 B.n17 10.6151
R2631 B.n960 B.n959 10.6151
R2632 B.n959 B.n958 10.6151
R2633 B.n958 B.n24 10.6151
R2634 B.n952 B.n24 10.6151
R2635 B.n952 B.n951 10.6151
R2636 B.n951 B.n950 10.6151
R2637 B.n950 B.n31 10.6151
R2638 B.n944 B.n31 10.6151
R2639 B.n944 B.n943 10.6151
R2640 B.n943 B.n942 10.6151
R2641 B.n942 B.n38 10.6151
R2642 B.n936 B.n38 10.6151
R2643 B.n936 B.n935 10.6151
R2644 B.n935 B.n934 10.6151
R2645 B.n934 B.n45 10.6151
R2646 B.n928 B.n45 10.6151
R2647 B.n928 B.n927 10.6151
R2648 B.n927 B.n926 10.6151
R2649 B.n926 B.n52 10.6151
R2650 B.n920 B.n52 10.6151
R2651 B.n794 B.n91 6.5566
R2652 B.n779 B.n778 6.5566
R2653 B.n399 B.n223 6.5566
R2654 B.n383 B.n382 6.5566
R2655 B.n544 B.t7 5.02437
R2656 B.n932 B.t11 5.02437
R2657 B.n798 B.n91 4.05904
R2658 B.n778 B.n777 4.05904
R2659 B.n223 B.n219 4.05904
R2660 B.n382 B.n381 4.05904
R2661 B.n586 B.t3 3.19751
R2662 B.t4 B.n962 3.19751
R2663 B.n982 B.n0 2.81026
R2664 B.n982 B.n1 2.81026
R2665 VN.n2 VN.t2 324.25
R2666 VN.n14 VN.t4 324.25
R2667 VN.n3 VN.t5 292.466
R2668 VN.n10 VN.t0 292.466
R2669 VN.n15 VN.t1 292.466
R2670 VN.n22 VN.t3 292.466
R2671 VN.n11 VN.n10 179.406
R2672 VN.n23 VN.n22 179.406
R2673 VN.n21 VN.n12 161.3
R2674 VN.n20 VN.n19 161.3
R2675 VN.n18 VN.n13 161.3
R2676 VN.n17 VN.n16 161.3
R2677 VN.n9 VN.n0 161.3
R2678 VN.n8 VN.n7 161.3
R2679 VN.n6 VN.n1 161.3
R2680 VN.n5 VN.n4 161.3
R2681 VN.n8 VN.n1 56.5193
R2682 VN.n20 VN.n13 56.5193
R2683 VN.n3 VN.n2 53.7793
R2684 VN.n15 VN.n14 53.7793
R2685 VN VN.n23 49.9797
R2686 VN.n4 VN.n1 24.4675
R2687 VN.n9 VN.n8 24.4675
R2688 VN.n16 VN.n13 24.4675
R2689 VN.n21 VN.n20 24.4675
R2690 VN.n17 VN.n14 18.144
R2691 VN.n5 VN.n2 18.144
R2692 VN.n4 VN.n3 12.234
R2693 VN.n16 VN.n15 12.234
R2694 VN.n10 VN.n9 6.36192
R2695 VN.n22 VN.n21 6.36192
R2696 VN.n23 VN.n12 0.189894
R2697 VN.n19 VN.n12 0.189894
R2698 VN.n19 VN.n18 0.189894
R2699 VN.n18 VN.n17 0.189894
R2700 VN.n6 VN.n5 0.189894
R2701 VN.n7 VN.n6 0.189894
R2702 VN.n7 VN.n0 0.189894
R2703 VN.n11 VN.n0 0.189894
R2704 VN VN.n11 0.0516364
R2705 VDD2.n207 VDD2.n206 289.615
R2706 VDD2.n102 VDD2.n101 289.615
R2707 VDD2.n206 VDD2.n205 185
R2708 VDD2.n107 VDD2.n106 185
R2709 VDD2.n200 VDD2.n199 185
R2710 VDD2.n198 VDD2.n197 185
R2711 VDD2.n111 VDD2.n110 185
R2712 VDD2.n192 VDD2.n191 185
R2713 VDD2.n190 VDD2.n189 185
R2714 VDD2.n115 VDD2.n114 185
R2715 VDD2.n184 VDD2.n183 185
R2716 VDD2.n182 VDD2.n181 185
R2717 VDD2.n119 VDD2.n118 185
R2718 VDD2.n176 VDD2.n175 185
R2719 VDD2.n174 VDD2.n173 185
R2720 VDD2.n123 VDD2.n122 185
R2721 VDD2.n168 VDD2.n167 185
R2722 VDD2.n166 VDD2.n165 185
R2723 VDD2.n127 VDD2.n126 185
R2724 VDD2.n131 VDD2.n129 185
R2725 VDD2.n160 VDD2.n159 185
R2726 VDD2.n158 VDD2.n157 185
R2727 VDD2.n133 VDD2.n132 185
R2728 VDD2.n152 VDD2.n151 185
R2729 VDD2.n150 VDD2.n149 185
R2730 VDD2.n137 VDD2.n136 185
R2731 VDD2.n144 VDD2.n143 185
R2732 VDD2.n142 VDD2.n141 185
R2733 VDD2.n35 VDD2.n34 185
R2734 VDD2.n37 VDD2.n36 185
R2735 VDD2.n30 VDD2.n29 185
R2736 VDD2.n43 VDD2.n42 185
R2737 VDD2.n45 VDD2.n44 185
R2738 VDD2.n26 VDD2.n25 185
R2739 VDD2.n52 VDD2.n51 185
R2740 VDD2.n53 VDD2.n24 185
R2741 VDD2.n55 VDD2.n54 185
R2742 VDD2.n22 VDD2.n21 185
R2743 VDD2.n61 VDD2.n60 185
R2744 VDD2.n63 VDD2.n62 185
R2745 VDD2.n18 VDD2.n17 185
R2746 VDD2.n69 VDD2.n68 185
R2747 VDD2.n71 VDD2.n70 185
R2748 VDD2.n14 VDD2.n13 185
R2749 VDD2.n77 VDD2.n76 185
R2750 VDD2.n79 VDD2.n78 185
R2751 VDD2.n10 VDD2.n9 185
R2752 VDD2.n85 VDD2.n84 185
R2753 VDD2.n87 VDD2.n86 185
R2754 VDD2.n6 VDD2.n5 185
R2755 VDD2.n93 VDD2.n92 185
R2756 VDD2.n95 VDD2.n94 185
R2757 VDD2.n2 VDD2.n1 185
R2758 VDD2.n101 VDD2.n100 185
R2759 VDD2.n140 VDD2.t2 149.524
R2760 VDD2.n33 VDD2.t3 149.524
R2761 VDD2.n206 VDD2.n106 104.615
R2762 VDD2.n199 VDD2.n106 104.615
R2763 VDD2.n199 VDD2.n198 104.615
R2764 VDD2.n198 VDD2.n110 104.615
R2765 VDD2.n191 VDD2.n110 104.615
R2766 VDD2.n191 VDD2.n190 104.615
R2767 VDD2.n190 VDD2.n114 104.615
R2768 VDD2.n183 VDD2.n114 104.615
R2769 VDD2.n183 VDD2.n182 104.615
R2770 VDD2.n182 VDD2.n118 104.615
R2771 VDD2.n175 VDD2.n118 104.615
R2772 VDD2.n175 VDD2.n174 104.615
R2773 VDD2.n174 VDD2.n122 104.615
R2774 VDD2.n167 VDD2.n122 104.615
R2775 VDD2.n167 VDD2.n166 104.615
R2776 VDD2.n166 VDD2.n126 104.615
R2777 VDD2.n131 VDD2.n126 104.615
R2778 VDD2.n159 VDD2.n131 104.615
R2779 VDD2.n159 VDD2.n158 104.615
R2780 VDD2.n158 VDD2.n132 104.615
R2781 VDD2.n151 VDD2.n132 104.615
R2782 VDD2.n151 VDD2.n150 104.615
R2783 VDD2.n150 VDD2.n136 104.615
R2784 VDD2.n143 VDD2.n136 104.615
R2785 VDD2.n143 VDD2.n142 104.615
R2786 VDD2.n36 VDD2.n35 104.615
R2787 VDD2.n36 VDD2.n29 104.615
R2788 VDD2.n43 VDD2.n29 104.615
R2789 VDD2.n44 VDD2.n43 104.615
R2790 VDD2.n44 VDD2.n25 104.615
R2791 VDD2.n52 VDD2.n25 104.615
R2792 VDD2.n53 VDD2.n52 104.615
R2793 VDD2.n54 VDD2.n53 104.615
R2794 VDD2.n54 VDD2.n21 104.615
R2795 VDD2.n61 VDD2.n21 104.615
R2796 VDD2.n62 VDD2.n61 104.615
R2797 VDD2.n62 VDD2.n17 104.615
R2798 VDD2.n69 VDD2.n17 104.615
R2799 VDD2.n70 VDD2.n69 104.615
R2800 VDD2.n70 VDD2.n13 104.615
R2801 VDD2.n77 VDD2.n13 104.615
R2802 VDD2.n78 VDD2.n77 104.615
R2803 VDD2.n78 VDD2.n9 104.615
R2804 VDD2.n85 VDD2.n9 104.615
R2805 VDD2.n86 VDD2.n85 104.615
R2806 VDD2.n86 VDD2.n5 104.615
R2807 VDD2.n93 VDD2.n5 104.615
R2808 VDD2.n94 VDD2.n93 104.615
R2809 VDD2.n94 VDD2.n1 104.615
R2810 VDD2.n101 VDD2.n1 104.615
R2811 VDD2.n104 VDD2.n103 64.5906
R2812 VDD2 VDD2.n209 64.5876
R2813 VDD2.n104 VDD2.n102 53.7092
R2814 VDD2.n208 VDD2.n207 52.549
R2815 VDD2.n142 VDD2.t2 52.3082
R2816 VDD2.n35 VDD2.t3 52.3082
R2817 VDD2.n208 VDD2.n104 45.1981
R2818 VDD2.n129 VDD2.n127 13.1884
R2819 VDD2.n55 VDD2.n22 13.1884
R2820 VDD2.n205 VDD2.n105 12.8005
R2821 VDD2.n165 VDD2.n164 12.8005
R2822 VDD2.n161 VDD2.n160 12.8005
R2823 VDD2.n56 VDD2.n24 12.8005
R2824 VDD2.n60 VDD2.n59 12.8005
R2825 VDD2.n100 VDD2.n0 12.8005
R2826 VDD2.n204 VDD2.n107 12.0247
R2827 VDD2.n168 VDD2.n125 12.0247
R2828 VDD2.n157 VDD2.n130 12.0247
R2829 VDD2.n51 VDD2.n50 12.0247
R2830 VDD2.n63 VDD2.n20 12.0247
R2831 VDD2.n99 VDD2.n2 12.0247
R2832 VDD2.n201 VDD2.n200 11.249
R2833 VDD2.n169 VDD2.n123 11.249
R2834 VDD2.n156 VDD2.n133 11.249
R2835 VDD2.n49 VDD2.n26 11.249
R2836 VDD2.n64 VDD2.n18 11.249
R2837 VDD2.n96 VDD2.n95 11.249
R2838 VDD2.n197 VDD2.n109 10.4732
R2839 VDD2.n173 VDD2.n172 10.4732
R2840 VDD2.n153 VDD2.n152 10.4732
R2841 VDD2.n46 VDD2.n45 10.4732
R2842 VDD2.n68 VDD2.n67 10.4732
R2843 VDD2.n92 VDD2.n4 10.4732
R2844 VDD2.n141 VDD2.n140 10.2747
R2845 VDD2.n34 VDD2.n33 10.2747
R2846 VDD2.n196 VDD2.n111 9.69747
R2847 VDD2.n176 VDD2.n121 9.69747
R2848 VDD2.n149 VDD2.n135 9.69747
R2849 VDD2.n42 VDD2.n28 9.69747
R2850 VDD2.n71 VDD2.n16 9.69747
R2851 VDD2.n91 VDD2.n6 9.69747
R2852 VDD2.n203 VDD2.n105 9.45567
R2853 VDD2.n98 VDD2.n0 9.45567
R2854 VDD2.n139 VDD2.n138 9.3005
R2855 VDD2.n146 VDD2.n145 9.3005
R2856 VDD2.n148 VDD2.n147 9.3005
R2857 VDD2.n135 VDD2.n134 9.3005
R2858 VDD2.n154 VDD2.n153 9.3005
R2859 VDD2.n156 VDD2.n155 9.3005
R2860 VDD2.n130 VDD2.n128 9.3005
R2861 VDD2.n162 VDD2.n161 9.3005
R2862 VDD2.n188 VDD2.n187 9.3005
R2863 VDD2.n113 VDD2.n112 9.3005
R2864 VDD2.n194 VDD2.n193 9.3005
R2865 VDD2.n196 VDD2.n195 9.3005
R2866 VDD2.n109 VDD2.n108 9.3005
R2867 VDD2.n202 VDD2.n201 9.3005
R2868 VDD2.n204 VDD2.n203 9.3005
R2869 VDD2.n186 VDD2.n185 9.3005
R2870 VDD2.n117 VDD2.n116 9.3005
R2871 VDD2.n180 VDD2.n179 9.3005
R2872 VDD2.n178 VDD2.n177 9.3005
R2873 VDD2.n121 VDD2.n120 9.3005
R2874 VDD2.n172 VDD2.n171 9.3005
R2875 VDD2.n170 VDD2.n169 9.3005
R2876 VDD2.n125 VDD2.n124 9.3005
R2877 VDD2.n164 VDD2.n163 9.3005
R2878 VDD2.n81 VDD2.n80 9.3005
R2879 VDD2.n83 VDD2.n82 9.3005
R2880 VDD2.n8 VDD2.n7 9.3005
R2881 VDD2.n89 VDD2.n88 9.3005
R2882 VDD2.n91 VDD2.n90 9.3005
R2883 VDD2.n4 VDD2.n3 9.3005
R2884 VDD2.n97 VDD2.n96 9.3005
R2885 VDD2.n99 VDD2.n98 9.3005
R2886 VDD2.n75 VDD2.n74 9.3005
R2887 VDD2.n73 VDD2.n72 9.3005
R2888 VDD2.n16 VDD2.n15 9.3005
R2889 VDD2.n67 VDD2.n66 9.3005
R2890 VDD2.n65 VDD2.n64 9.3005
R2891 VDD2.n20 VDD2.n19 9.3005
R2892 VDD2.n59 VDD2.n58 9.3005
R2893 VDD2.n32 VDD2.n31 9.3005
R2894 VDD2.n39 VDD2.n38 9.3005
R2895 VDD2.n41 VDD2.n40 9.3005
R2896 VDD2.n28 VDD2.n27 9.3005
R2897 VDD2.n47 VDD2.n46 9.3005
R2898 VDD2.n49 VDD2.n48 9.3005
R2899 VDD2.n50 VDD2.n23 9.3005
R2900 VDD2.n57 VDD2.n56 9.3005
R2901 VDD2.n12 VDD2.n11 9.3005
R2902 VDD2.n193 VDD2.n192 8.92171
R2903 VDD2.n177 VDD2.n119 8.92171
R2904 VDD2.n148 VDD2.n137 8.92171
R2905 VDD2.n41 VDD2.n30 8.92171
R2906 VDD2.n72 VDD2.n14 8.92171
R2907 VDD2.n88 VDD2.n87 8.92171
R2908 VDD2.n189 VDD2.n113 8.14595
R2909 VDD2.n181 VDD2.n180 8.14595
R2910 VDD2.n145 VDD2.n144 8.14595
R2911 VDD2.n38 VDD2.n37 8.14595
R2912 VDD2.n76 VDD2.n75 8.14595
R2913 VDD2.n84 VDD2.n8 8.14595
R2914 VDD2.n188 VDD2.n115 7.3702
R2915 VDD2.n184 VDD2.n117 7.3702
R2916 VDD2.n141 VDD2.n139 7.3702
R2917 VDD2.n34 VDD2.n32 7.3702
R2918 VDD2.n79 VDD2.n12 7.3702
R2919 VDD2.n83 VDD2.n10 7.3702
R2920 VDD2.n185 VDD2.n115 6.59444
R2921 VDD2.n185 VDD2.n184 6.59444
R2922 VDD2.n80 VDD2.n79 6.59444
R2923 VDD2.n80 VDD2.n10 6.59444
R2924 VDD2.n189 VDD2.n188 5.81868
R2925 VDD2.n181 VDD2.n117 5.81868
R2926 VDD2.n144 VDD2.n139 5.81868
R2927 VDD2.n37 VDD2.n32 5.81868
R2928 VDD2.n76 VDD2.n12 5.81868
R2929 VDD2.n84 VDD2.n83 5.81868
R2930 VDD2.n192 VDD2.n113 5.04292
R2931 VDD2.n180 VDD2.n119 5.04292
R2932 VDD2.n145 VDD2.n137 5.04292
R2933 VDD2.n38 VDD2.n30 5.04292
R2934 VDD2.n75 VDD2.n14 5.04292
R2935 VDD2.n87 VDD2.n8 5.04292
R2936 VDD2.n193 VDD2.n111 4.26717
R2937 VDD2.n177 VDD2.n176 4.26717
R2938 VDD2.n149 VDD2.n148 4.26717
R2939 VDD2.n42 VDD2.n41 4.26717
R2940 VDD2.n72 VDD2.n71 4.26717
R2941 VDD2.n88 VDD2.n6 4.26717
R2942 VDD2.n197 VDD2.n196 3.49141
R2943 VDD2.n173 VDD2.n121 3.49141
R2944 VDD2.n152 VDD2.n135 3.49141
R2945 VDD2.n45 VDD2.n28 3.49141
R2946 VDD2.n68 VDD2.n16 3.49141
R2947 VDD2.n92 VDD2.n91 3.49141
R2948 VDD2.n33 VDD2.n31 2.84303
R2949 VDD2.n140 VDD2.n138 2.84303
R2950 VDD2.n200 VDD2.n109 2.71565
R2951 VDD2.n172 VDD2.n123 2.71565
R2952 VDD2.n153 VDD2.n133 2.71565
R2953 VDD2.n46 VDD2.n26 2.71565
R2954 VDD2.n67 VDD2.n18 2.71565
R2955 VDD2.n95 VDD2.n4 2.71565
R2956 VDD2.n201 VDD2.n107 1.93989
R2957 VDD2.n169 VDD2.n168 1.93989
R2958 VDD2.n157 VDD2.n156 1.93989
R2959 VDD2.n51 VDD2.n49 1.93989
R2960 VDD2.n64 VDD2.n63 1.93989
R2961 VDD2.n96 VDD2.n2 1.93989
R2962 VDD2 VDD2.n208 1.27421
R2963 VDD2.n205 VDD2.n204 1.16414
R2964 VDD2.n165 VDD2.n125 1.16414
R2965 VDD2.n160 VDD2.n130 1.16414
R2966 VDD2.n50 VDD2.n24 1.16414
R2967 VDD2.n60 VDD2.n20 1.16414
R2968 VDD2.n100 VDD2.n99 1.16414
R2969 VDD2.n209 VDD2.t4 1.05313
R2970 VDD2.n209 VDD2.t1 1.05313
R2971 VDD2.n103 VDD2.t0 1.05313
R2972 VDD2.n103 VDD2.t5 1.05313
R2973 VDD2.n207 VDD2.n105 0.388379
R2974 VDD2.n164 VDD2.n127 0.388379
R2975 VDD2.n161 VDD2.n129 0.388379
R2976 VDD2.n56 VDD2.n55 0.388379
R2977 VDD2.n59 VDD2.n22 0.388379
R2978 VDD2.n102 VDD2.n0 0.388379
R2979 VDD2.n203 VDD2.n202 0.155672
R2980 VDD2.n202 VDD2.n108 0.155672
R2981 VDD2.n195 VDD2.n108 0.155672
R2982 VDD2.n195 VDD2.n194 0.155672
R2983 VDD2.n194 VDD2.n112 0.155672
R2984 VDD2.n187 VDD2.n112 0.155672
R2985 VDD2.n187 VDD2.n186 0.155672
R2986 VDD2.n186 VDD2.n116 0.155672
R2987 VDD2.n179 VDD2.n116 0.155672
R2988 VDD2.n179 VDD2.n178 0.155672
R2989 VDD2.n178 VDD2.n120 0.155672
R2990 VDD2.n171 VDD2.n120 0.155672
R2991 VDD2.n171 VDD2.n170 0.155672
R2992 VDD2.n170 VDD2.n124 0.155672
R2993 VDD2.n163 VDD2.n124 0.155672
R2994 VDD2.n163 VDD2.n162 0.155672
R2995 VDD2.n162 VDD2.n128 0.155672
R2996 VDD2.n155 VDD2.n128 0.155672
R2997 VDD2.n155 VDD2.n154 0.155672
R2998 VDD2.n154 VDD2.n134 0.155672
R2999 VDD2.n147 VDD2.n134 0.155672
R3000 VDD2.n147 VDD2.n146 0.155672
R3001 VDD2.n146 VDD2.n138 0.155672
R3002 VDD2.n39 VDD2.n31 0.155672
R3003 VDD2.n40 VDD2.n39 0.155672
R3004 VDD2.n40 VDD2.n27 0.155672
R3005 VDD2.n47 VDD2.n27 0.155672
R3006 VDD2.n48 VDD2.n47 0.155672
R3007 VDD2.n48 VDD2.n23 0.155672
R3008 VDD2.n57 VDD2.n23 0.155672
R3009 VDD2.n58 VDD2.n57 0.155672
R3010 VDD2.n58 VDD2.n19 0.155672
R3011 VDD2.n65 VDD2.n19 0.155672
R3012 VDD2.n66 VDD2.n65 0.155672
R3013 VDD2.n66 VDD2.n15 0.155672
R3014 VDD2.n73 VDD2.n15 0.155672
R3015 VDD2.n74 VDD2.n73 0.155672
R3016 VDD2.n74 VDD2.n11 0.155672
R3017 VDD2.n81 VDD2.n11 0.155672
R3018 VDD2.n82 VDD2.n81 0.155672
R3019 VDD2.n82 VDD2.n7 0.155672
R3020 VDD2.n89 VDD2.n7 0.155672
R3021 VDD2.n90 VDD2.n89 0.155672
R3022 VDD2.n90 VDD2.n3 0.155672
R3023 VDD2.n97 VDD2.n3 0.155672
R3024 VDD2.n98 VDD2.n97 0.155672
C0 VN VP 7.16886f
C1 VTAIL VP 8.75087f
C2 VDD1 VP 9.314099f
C3 VN VTAIL 8.73629f
C4 VDD2 VP 0.370236f
C5 VDD1 VN 0.149371f
C6 VDD1 VTAIL 11.0222f
C7 VDD2 VN 9.09859f
C8 VDD2 VTAIL 11.062f
C9 VDD1 VDD2 1.02769f
C10 VDD2 B 6.365029f
C11 VDD1 B 6.445857f
C12 VTAIL B 9.704607f
C13 VN B 10.586842f
C14 VP B 8.787124f
C15 VDD2.n0 B 0.012184f
C16 VDD2.n1 B 0.027437f
C17 VDD2.n2 B 0.012291f
C18 VDD2.n3 B 0.021602f
C19 VDD2.n4 B 0.011608f
C20 VDD2.n5 B 0.027437f
C21 VDD2.n6 B 0.012291f
C22 VDD2.n7 B 0.021602f
C23 VDD2.n8 B 0.011608f
C24 VDD2.n9 B 0.027437f
C25 VDD2.n10 B 0.012291f
C26 VDD2.n11 B 0.021602f
C27 VDD2.n12 B 0.011608f
C28 VDD2.n13 B 0.027437f
C29 VDD2.n14 B 0.012291f
C30 VDD2.n15 B 0.021602f
C31 VDD2.n16 B 0.011608f
C32 VDD2.n17 B 0.027437f
C33 VDD2.n18 B 0.012291f
C34 VDD2.n19 B 0.021602f
C35 VDD2.n20 B 0.011608f
C36 VDD2.n21 B 0.027437f
C37 VDD2.n22 B 0.011949f
C38 VDD2.n23 B 0.021602f
C39 VDD2.n24 B 0.012291f
C40 VDD2.n25 B 0.027437f
C41 VDD2.n26 B 0.012291f
C42 VDD2.n27 B 0.021602f
C43 VDD2.n28 B 0.011608f
C44 VDD2.n29 B 0.027437f
C45 VDD2.n30 B 0.012291f
C46 VDD2.n31 B 1.74408f
C47 VDD2.n32 B 0.011608f
C48 VDD2.t3 B 0.047131f
C49 VDD2.n33 B 0.212223f
C50 VDD2.n34 B 0.019396f
C51 VDD2.n35 B 0.020577f
C52 VDD2.n36 B 0.027437f
C53 VDD2.n37 B 0.012291f
C54 VDD2.n38 B 0.011608f
C55 VDD2.n39 B 0.021602f
C56 VDD2.n40 B 0.021602f
C57 VDD2.n41 B 0.011608f
C58 VDD2.n42 B 0.012291f
C59 VDD2.n43 B 0.027437f
C60 VDD2.n44 B 0.027437f
C61 VDD2.n45 B 0.012291f
C62 VDD2.n46 B 0.011608f
C63 VDD2.n47 B 0.021602f
C64 VDD2.n48 B 0.021602f
C65 VDD2.n49 B 0.011608f
C66 VDD2.n50 B 0.011608f
C67 VDD2.n51 B 0.012291f
C68 VDD2.n52 B 0.027437f
C69 VDD2.n53 B 0.027437f
C70 VDD2.n54 B 0.027437f
C71 VDD2.n55 B 0.011949f
C72 VDD2.n56 B 0.011608f
C73 VDD2.n57 B 0.021602f
C74 VDD2.n58 B 0.021602f
C75 VDD2.n59 B 0.011608f
C76 VDD2.n60 B 0.012291f
C77 VDD2.n61 B 0.027437f
C78 VDD2.n62 B 0.027437f
C79 VDD2.n63 B 0.012291f
C80 VDD2.n64 B 0.011608f
C81 VDD2.n65 B 0.021602f
C82 VDD2.n66 B 0.021602f
C83 VDD2.n67 B 0.011608f
C84 VDD2.n68 B 0.012291f
C85 VDD2.n69 B 0.027437f
C86 VDD2.n70 B 0.027437f
C87 VDD2.n71 B 0.012291f
C88 VDD2.n72 B 0.011608f
C89 VDD2.n73 B 0.021602f
C90 VDD2.n74 B 0.021602f
C91 VDD2.n75 B 0.011608f
C92 VDD2.n76 B 0.012291f
C93 VDD2.n77 B 0.027437f
C94 VDD2.n78 B 0.027437f
C95 VDD2.n79 B 0.012291f
C96 VDD2.n80 B 0.011608f
C97 VDD2.n81 B 0.021602f
C98 VDD2.n82 B 0.021602f
C99 VDD2.n83 B 0.011608f
C100 VDD2.n84 B 0.012291f
C101 VDD2.n85 B 0.027437f
C102 VDD2.n86 B 0.027437f
C103 VDD2.n87 B 0.012291f
C104 VDD2.n88 B 0.011608f
C105 VDD2.n89 B 0.021602f
C106 VDD2.n90 B 0.021602f
C107 VDD2.n91 B 0.011608f
C108 VDD2.n92 B 0.012291f
C109 VDD2.n93 B 0.027437f
C110 VDD2.n94 B 0.027437f
C111 VDD2.n95 B 0.012291f
C112 VDD2.n96 B 0.011608f
C113 VDD2.n97 B 0.021602f
C114 VDD2.n98 B 0.056128f
C115 VDD2.n99 B 0.011608f
C116 VDD2.n100 B 0.012291f
C117 VDD2.n101 B 0.056561f
C118 VDD2.n102 B 0.065363f
C119 VDD2.t0 B 0.321093f
C120 VDD2.t5 B 0.321093f
C121 VDD2.n103 B 2.94033f
C122 VDD2.n104 B 2.28425f
C123 VDD2.n105 B 0.012184f
C124 VDD2.n106 B 0.027437f
C125 VDD2.n107 B 0.012291f
C126 VDD2.n108 B 0.021602f
C127 VDD2.n109 B 0.011608f
C128 VDD2.n110 B 0.027437f
C129 VDD2.n111 B 0.012291f
C130 VDD2.n112 B 0.021602f
C131 VDD2.n113 B 0.011608f
C132 VDD2.n114 B 0.027437f
C133 VDD2.n115 B 0.012291f
C134 VDD2.n116 B 0.021602f
C135 VDD2.n117 B 0.011608f
C136 VDD2.n118 B 0.027437f
C137 VDD2.n119 B 0.012291f
C138 VDD2.n120 B 0.021602f
C139 VDD2.n121 B 0.011608f
C140 VDD2.n122 B 0.027437f
C141 VDD2.n123 B 0.012291f
C142 VDD2.n124 B 0.021602f
C143 VDD2.n125 B 0.011608f
C144 VDD2.n126 B 0.027437f
C145 VDD2.n127 B 0.011949f
C146 VDD2.n128 B 0.021602f
C147 VDD2.n129 B 0.011949f
C148 VDD2.n130 B 0.011608f
C149 VDD2.n131 B 0.027437f
C150 VDD2.n132 B 0.027437f
C151 VDD2.n133 B 0.012291f
C152 VDD2.n134 B 0.021602f
C153 VDD2.n135 B 0.011608f
C154 VDD2.n136 B 0.027437f
C155 VDD2.n137 B 0.012291f
C156 VDD2.n138 B 1.74408f
C157 VDD2.n139 B 0.011608f
C158 VDD2.t2 B 0.047131f
C159 VDD2.n140 B 0.212223f
C160 VDD2.n141 B 0.019396f
C161 VDD2.n142 B 0.020577f
C162 VDD2.n143 B 0.027437f
C163 VDD2.n144 B 0.012291f
C164 VDD2.n145 B 0.011608f
C165 VDD2.n146 B 0.021602f
C166 VDD2.n147 B 0.021602f
C167 VDD2.n148 B 0.011608f
C168 VDD2.n149 B 0.012291f
C169 VDD2.n150 B 0.027437f
C170 VDD2.n151 B 0.027437f
C171 VDD2.n152 B 0.012291f
C172 VDD2.n153 B 0.011608f
C173 VDD2.n154 B 0.021602f
C174 VDD2.n155 B 0.021602f
C175 VDD2.n156 B 0.011608f
C176 VDD2.n157 B 0.012291f
C177 VDD2.n158 B 0.027437f
C178 VDD2.n159 B 0.027437f
C179 VDD2.n160 B 0.012291f
C180 VDD2.n161 B 0.011608f
C181 VDD2.n162 B 0.021602f
C182 VDD2.n163 B 0.021602f
C183 VDD2.n164 B 0.011608f
C184 VDD2.n165 B 0.012291f
C185 VDD2.n166 B 0.027437f
C186 VDD2.n167 B 0.027437f
C187 VDD2.n168 B 0.012291f
C188 VDD2.n169 B 0.011608f
C189 VDD2.n170 B 0.021602f
C190 VDD2.n171 B 0.021602f
C191 VDD2.n172 B 0.011608f
C192 VDD2.n173 B 0.012291f
C193 VDD2.n174 B 0.027437f
C194 VDD2.n175 B 0.027437f
C195 VDD2.n176 B 0.012291f
C196 VDD2.n177 B 0.011608f
C197 VDD2.n178 B 0.021602f
C198 VDD2.n179 B 0.021602f
C199 VDD2.n180 B 0.011608f
C200 VDD2.n181 B 0.012291f
C201 VDD2.n182 B 0.027437f
C202 VDD2.n183 B 0.027437f
C203 VDD2.n184 B 0.012291f
C204 VDD2.n185 B 0.011608f
C205 VDD2.n186 B 0.021602f
C206 VDD2.n187 B 0.021602f
C207 VDD2.n188 B 0.011608f
C208 VDD2.n189 B 0.012291f
C209 VDD2.n190 B 0.027437f
C210 VDD2.n191 B 0.027437f
C211 VDD2.n192 B 0.012291f
C212 VDD2.n193 B 0.011608f
C213 VDD2.n194 B 0.021602f
C214 VDD2.n195 B 0.021602f
C215 VDD2.n196 B 0.011608f
C216 VDD2.n197 B 0.012291f
C217 VDD2.n198 B 0.027437f
C218 VDD2.n199 B 0.027437f
C219 VDD2.n200 B 0.012291f
C220 VDD2.n201 B 0.011608f
C221 VDD2.n202 B 0.021602f
C222 VDD2.n203 B 0.056128f
C223 VDD2.n204 B 0.011608f
C224 VDD2.n205 B 0.012291f
C225 VDD2.n206 B 0.056561f
C226 VDD2.n207 B 0.062642f
C227 VDD2.n208 B 2.42002f
C228 VDD2.t4 B 0.321093f
C229 VDD2.t1 B 0.321093f
C230 VDD2.n209 B 2.9403f
C231 VN.n0 B 0.030893f
C232 VN.t0 B 2.47949f
C233 VN.n1 B 0.039934f
C234 VN.t2 B 2.57671f
C235 VN.n2 B 0.948185f
C236 VN.t5 B 2.47949f
C237 VN.n3 B 0.928591f
C238 VN.n4 B 0.043364f
C239 VN.n5 B 0.19486f
C240 VN.n6 B 0.030893f
C241 VN.n7 B 0.030893f
C242 VN.n8 B 0.050264f
C243 VN.n9 B 0.036542f
C244 VN.n10 B 0.930803f
C245 VN.n11 B 0.030785f
C246 VN.n12 B 0.030893f
C247 VN.t3 B 2.47949f
C248 VN.n13 B 0.039934f
C249 VN.t4 B 2.57671f
C250 VN.n14 B 0.948185f
C251 VN.t1 B 2.47949f
C252 VN.n15 B 0.928591f
C253 VN.n16 B 0.043364f
C254 VN.n17 B 0.19486f
C255 VN.n18 B 0.030893f
C256 VN.n19 B 0.030893f
C257 VN.n20 B 0.050264f
C258 VN.n21 B 0.036542f
C259 VN.n22 B 0.930803f
C260 VN.n23 B 1.68626f
C261 VTAIL.t1 B 0.331622f
C262 VTAIL.t4 B 0.331622f
C263 VTAIL.n0 B 2.97431f
C264 VTAIL.n1 B 0.332909f
C265 VTAIL.n2 B 0.012583f
C266 VTAIL.n3 B 0.028336f
C267 VTAIL.n4 B 0.012694f
C268 VTAIL.n5 B 0.02231f
C269 VTAIL.n6 B 0.011989f
C270 VTAIL.n7 B 0.028336f
C271 VTAIL.n8 B 0.012694f
C272 VTAIL.n9 B 0.02231f
C273 VTAIL.n10 B 0.011989f
C274 VTAIL.n11 B 0.028336f
C275 VTAIL.n12 B 0.012694f
C276 VTAIL.n13 B 0.02231f
C277 VTAIL.n14 B 0.011989f
C278 VTAIL.n15 B 0.028336f
C279 VTAIL.n16 B 0.012694f
C280 VTAIL.n17 B 0.02231f
C281 VTAIL.n18 B 0.011989f
C282 VTAIL.n19 B 0.028336f
C283 VTAIL.n20 B 0.012694f
C284 VTAIL.n21 B 0.02231f
C285 VTAIL.n22 B 0.011989f
C286 VTAIL.n23 B 0.028336f
C287 VTAIL.n24 B 0.012341f
C288 VTAIL.n25 B 0.02231f
C289 VTAIL.n26 B 0.012694f
C290 VTAIL.n27 B 0.028336f
C291 VTAIL.n28 B 0.012694f
C292 VTAIL.n29 B 0.02231f
C293 VTAIL.n30 B 0.011989f
C294 VTAIL.n31 B 0.028336f
C295 VTAIL.n32 B 0.012694f
C296 VTAIL.n33 B 1.80128f
C297 VTAIL.n34 B 0.011989f
C298 VTAIL.t6 B 0.048676f
C299 VTAIL.n35 B 0.219182f
C300 VTAIL.n36 B 0.020032f
C301 VTAIL.n37 B 0.021252f
C302 VTAIL.n38 B 0.028336f
C303 VTAIL.n39 B 0.012694f
C304 VTAIL.n40 B 0.011989f
C305 VTAIL.n41 B 0.02231f
C306 VTAIL.n42 B 0.02231f
C307 VTAIL.n43 B 0.011989f
C308 VTAIL.n44 B 0.012694f
C309 VTAIL.n45 B 0.028336f
C310 VTAIL.n46 B 0.028336f
C311 VTAIL.n47 B 0.012694f
C312 VTAIL.n48 B 0.011989f
C313 VTAIL.n49 B 0.02231f
C314 VTAIL.n50 B 0.02231f
C315 VTAIL.n51 B 0.011989f
C316 VTAIL.n52 B 0.011989f
C317 VTAIL.n53 B 0.012694f
C318 VTAIL.n54 B 0.028336f
C319 VTAIL.n55 B 0.028336f
C320 VTAIL.n56 B 0.028336f
C321 VTAIL.n57 B 0.012341f
C322 VTAIL.n58 B 0.011989f
C323 VTAIL.n59 B 0.02231f
C324 VTAIL.n60 B 0.02231f
C325 VTAIL.n61 B 0.011989f
C326 VTAIL.n62 B 0.012694f
C327 VTAIL.n63 B 0.028336f
C328 VTAIL.n64 B 0.028336f
C329 VTAIL.n65 B 0.012694f
C330 VTAIL.n66 B 0.011989f
C331 VTAIL.n67 B 0.02231f
C332 VTAIL.n68 B 0.02231f
C333 VTAIL.n69 B 0.011989f
C334 VTAIL.n70 B 0.012694f
C335 VTAIL.n71 B 0.028336f
C336 VTAIL.n72 B 0.028336f
C337 VTAIL.n73 B 0.012694f
C338 VTAIL.n74 B 0.011989f
C339 VTAIL.n75 B 0.02231f
C340 VTAIL.n76 B 0.02231f
C341 VTAIL.n77 B 0.011989f
C342 VTAIL.n78 B 0.012694f
C343 VTAIL.n79 B 0.028336f
C344 VTAIL.n80 B 0.028336f
C345 VTAIL.n81 B 0.012694f
C346 VTAIL.n82 B 0.011989f
C347 VTAIL.n83 B 0.02231f
C348 VTAIL.n84 B 0.02231f
C349 VTAIL.n85 B 0.011989f
C350 VTAIL.n86 B 0.012694f
C351 VTAIL.n87 B 0.028336f
C352 VTAIL.n88 B 0.028336f
C353 VTAIL.n89 B 0.012694f
C354 VTAIL.n90 B 0.011989f
C355 VTAIL.n91 B 0.02231f
C356 VTAIL.n92 B 0.02231f
C357 VTAIL.n93 B 0.011989f
C358 VTAIL.n94 B 0.012694f
C359 VTAIL.n95 B 0.028336f
C360 VTAIL.n96 B 0.028336f
C361 VTAIL.n97 B 0.012694f
C362 VTAIL.n98 B 0.011989f
C363 VTAIL.n99 B 0.02231f
C364 VTAIL.n100 B 0.057969f
C365 VTAIL.n101 B 0.011989f
C366 VTAIL.n102 B 0.012694f
C367 VTAIL.n103 B 0.058415f
C368 VTAIL.n104 B 0.049332f
C369 VTAIL.n105 B 0.230869f
C370 VTAIL.t9 B 0.331622f
C371 VTAIL.t10 B 0.331622f
C372 VTAIL.n106 B 2.97431f
C373 VTAIL.n107 B 2.02585f
C374 VTAIL.t2 B 0.331622f
C375 VTAIL.t3 B 0.331622f
C376 VTAIL.n108 B 2.9743f
C377 VTAIL.n109 B 2.02586f
C378 VTAIL.n110 B 0.012583f
C379 VTAIL.n111 B 0.028336f
C380 VTAIL.n112 B 0.012694f
C381 VTAIL.n113 B 0.02231f
C382 VTAIL.n114 B 0.011989f
C383 VTAIL.n115 B 0.028336f
C384 VTAIL.n116 B 0.012694f
C385 VTAIL.n117 B 0.02231f
C386 VTAIL.n118 B 0.011989f
C387 VTAIL.n119 B 0.028336f
C388 VTAIL.n120 B 0.012694f
C389 VTAIL.n121 B 0.02231f
C390 VTAIL.n122 B 0.011989f
C391 VTAIL.n123 B 0.028336f
C392 VTAIL.n124 B 0.012694f
C393 VTAIL.n125 B 0.02231f
C394 VTAIL.n126 B 0.011989f
C395 VTAIL.n127 B 0.028336f
C396 VTAIL.n128 B 0.012694f
C397 VTAIL.n129 B 0.02231f
C398 VTAIL.n130 B 0.011989f
C399 VTAIL.n131 B 0.028336f
C400 VTAIL.n132 B 0.012341f
C401 VTAIL.n133 B 0.02231f
C402 VTAIL.n134 B 0.012341f
C403 VTAIL.n135 B 0.011989f
C404 VTAIL.n136 B 0.028336f
C405 VTAIL.n137 B 0.028336f
C406 VTAIL.n138 B 0.012694f
C407 VTAIL.n139 B 0.02231f
C408 VTAIL.n140 B 0.011989f
C409 VTAIL.n141 B 0.028336f
C410 VTAIL.n142 B 0.012694f
C411 VTAIL.n143 B 1.80128f
C412 VTAIL.n144 B 0.011989f
C413 VTAIL.t0 B 0.048676f
C414 VTAIL.n145 B 0.219182f
C415 VTAIL.n146 B 0.020032f
C416 VTAIL.n147 B 0.021252f
C417 VTAIL.n148 B 0.028336f
C418 VTAIL.n149 B 0.012694f
C419 VTAIL.n150 B 0.011989f
C420 VTAIL.n151 B 0.02231f
C421 VTAIL.n152 B 0.02231f
C422 VTAIL.n153 B 0.011989f
C423 VTAIL.n154 B 0.012694f
C424 VTAIL.n155 B 0.028336f
C425 VTAIL.n156 B 0.028336f
C426 VTAIL.n157 B 0.012694f
C427 VTAIL.n158 B 0.011989f
C428 VTAIL.n159 B 0.02231f
C429 VTAIL.n160 B 0.02231f
C430 VTAIL.n161 B 0.011989f
C431 VTAIL.n162 B 0.012694f
C432 VTAIL.n163 B 0.028336f
C433 VTAIL.n164 B 0.028336f
C434 VTAIL.n165 B 0.012694f
C435 VTAIL.n166 B 0.011989f
C436 VTAIL.n167 B 0.02231f
C437 VTAIL.n168 B 0.02231f
C438 VTAIL.n169 B 0.011989f
C439 VTAIL.n170 B 0.012694f
C440 VTAIL.n171 B 0.028336f
C441 VTAIL.n172 B 0.028336f
C442 VTAIL.n173 B 0.012694f
C443 VTAIL.n174 B 0.011989f
C444 VTAIL.n175 B 0.02231f
C445 VTAIL.n176 B 0.02231f
C446 VTAIL.n177 B 0.011989f
C447 VTAIL.n178 B 0.012694f
C448 VTAIL.n179 B 0.028336f
C449 VTAIL.n180 B 0.028336f
C450 VTAIL.n181 B 0.012694f
C451 VTAIL.n182 B 0.011989f
C452 VTAIL.n183 B 0.02231f
C453 VTAIL.n184 B 0.02231f
C454 VTAIL.n185 B 0.011989f
C455 VTAIL.n186 B 0.012694f
C456 VTAIL.n187 B 0.028336f
C457 VTAIL.n188 B 0.028336f
C458 VTAIL.n189 B 0.012694f
C459 VTAIL.n190 B 0.011989f
C460 VTAIL.n191 B 0.02231f
C461 VTAIL.n192 B 0.02231f
C462 VTAIL.n193 B 0.011989f
C463 VTAIL.n194 B 0.012694f
C464 VTAIL.n195 B 0.028336f
C465 VTAIL.n196 B 0.028336f
C466 VTAIL.n197 B 0.012694f
C467 VTAIL.n198 B 0.011989f
C468 VTAIL.n199 B 0.02231f
C469 VTAIL.n200 B 0.02231f
C470 VTAIL.n201 B 0.011989f
C471 VTAIL.n202 B 0.012694f
C472 VTAIL.n203 B 0.028336f
C473 VTAIL.n204 B 0.028336f
C474 VTAIL.n205 B 0.012694f
C475 VTAIL.n206 B 0.011989f
C476 VTAIL.n207 B 0.02231f
C477 VTAIL.n208 B 0.057969f
C478 VTAIL.n209 B 0.011989f
C479 VTAIL.n210 B 0.012694f
C480 VTAIL.n211 B 0.058415f
C481 VTAIL.n212 B 0.049332f
C482 VTAIL.n213 B 0.230869f
C483 VTAIL.t8 B 0.331622f
C484 VTAIL.t11 B 0.331622f
C485 VTAIL.n214 B 2.9743f
C486 VTAIL.n215 B 0.416115f
C487 VTAIL.n216 B 0.012583f
C488 VTAIL.n217 B 0.028336f
C489 VTAIL.n218 B 0.012694f
C490 VTAIL.n219 B 0.02231f
C491 VTAIL.n220 B 0.011989f
C492 VTAIL.n221 B 0.028336f
C493 VTAIL.n222 B 0.012694f
C494 VTAIL.n223 B 0.02231f
C495 VTAIL.n224 B 0.011989f
C496 VTAIL.n225 B 0.028336f
C497 VTAIL.n226 B 0.012694f
C498 VTAIL.n227 B 0.02231f
C499 VTAIL.n228 B 0.011989f
C500 VTAIL.n229 B 0.028336f
C501 VTAIL.n230 B 0.012694f
C502 VTAIL.n231 B 0.02231f
C503 VTAIL.n232 B 0.011989f
C504 VTAIL.n233 B 0.028336f
C505 VTAIL.n234 B 0.012694f
C506 VTAIL.n235 B 0.02231f
C507 VTAIL.n236 B 0.011989f
C508 VTAIL.n237 B 0.028336f
C509 VTAIL.n238 B 0.012341f
C510 VTAIL.n239 B 0.02231f
C511 VTAIL.n240 B 0.012341f
C512 VTAIL.n241 B 0.011989f
C513 VTAIL.n242 B 0.028336f
C514 VTAIL.n243 B 0.028336f
C515 VTAIL.n244 B 0.012694f
C516 VTAIL.n245 B 0.02231f
C517 VTAIL.n246 B 0.011989f
C518 VTAIL.n247 B 0.028336f
C519 VTAIL.n248 B 0.012694f
C520 VTAIL.n249 B 1.80128f
C521 VTAIL.n250 B 0.011989f
C522 VTAIL.t7 B 0.048676f
C523 VTAIL.n251 B 0.219183f
C524 VTAIL.n252 B 0.020032f
C525 VTAIL.n253 B 0.021252f
C526 VTAIL.n254 B 0.028336f
C527 VTAIL.n255 B 0.012694f
C528 VTAIL.n256 B 0.011989f
C529 VTAIL.n257 B 0.02231f
C530 VTAIL.n258 B 0.02231f
C531 VTAIL.n259 B 0.011989f
C532 VTAIL.n260 B 0.012694f
C533 VTAIL.n261 B 0.028336f
C534 VTAIL.n262 B 0.028336f
C535 VTAIL.n263 B 0.012694f
C536 VTAIL.n264 B 0.011989f
C537 VTAIL.n265 B 0.02231f
C538 VTAIL.n266 B 0.02231f
C539 VTAIL.n267 B 0.011989f
C540 VTAIL.n268 B 0.012694f
C541 VTAIL.n269 B 0.028336f
C542 VTAIL.n270 B 0.028336f
C543 VTAIL.n271 B 0.012694f
C544 VTAIL.n272 B 0.011989f
C545 VTAIL.n273 B 0.02231f
C546 VTAIL.n274 B 0.02231f
C547 VTAIL.n275 B 0.011989f
C548 VTAIL.n276 B 0.012694f
C549 VTAIL.n277 B 0.028336f
C550 VTAIL.n278 B 0.028336f
C551 VTAIL.n279 B 0.012694f
C552 VTAIL.n280 B 0.011989f
C553 VTAIL.n281 B 0.02231f
C554 VTAIL.n282 B 0.02231f
C555 VTAIL.n283 B 0.011989f
C556 VTAIL.n284 B 0.012694f
C557 VTAIL.n285 B 0.028336f
C558 VTAIL.n286 B 0.028336f
C559 VTAIL.n287 B 0.012694f
C560 VTAIL.n288 B 0.011989f
C561 VTAIL.n289 B 0.02231f
C562 VTAIL.n290 B 0.02231f
C563 VTAIL.n291 B 0.011989f
C564 VTAIL.n292 B 0.012694f
C565 VTAIL.n293 B 0.028336f
C566 VTAIL.n294 B 0.028336f
C567 VTAIL.n295 B 0.012694f
C568 VTAIL.n296 B 0.011989f
C569 VTAIL.n297 B 0.02231f
C570 VTAIL.n298 B 0.02231f
C571 VTAIL.n299 B 0.011989f
C572 VTAIL.n300 B 0.012694f
C573 VTAIL.n301 B 0.028336f
C574 VTAIL.n302 B 0.028336f
C575 VTAIL.n303 B 0.012694f
C576 VTAIL.n304 B 0.011989f
C577 VTAIL.n305 B 0.02231f
C578 VTAIL.n306 B 0.02231f
C579 VTAIL.n307 B 0.011989f
C580 VTAIL.n308 B 0.012694f
C581 VTAIL.n309 B 0.028336f
C582 VTAIL.n310 B 0.028336f
C583 VTAIL.n311 B 0.012694f
C584 VTAIL.n312 B 0.011989f
C585 VTAIL.n313 B 0.02231f
C586 VTAIL.n314 B 0.057969f
C587 VTAIL.n315 B 0.011989f
C588 VTAIL.n316 B 0.012694f
C589 VTAIL.n317 B 0.058415f
C590 VTAIL.n318 B 0.049332f
C591 VTAIL.n319 B 1.72411f
C592 VTAIL.n320 B 0.012583f
C593 VTAIL.n321 B 0.028336f
C594 VTAIL.n322 B 0.012694f
C595 VTAIL.n323 B 0.02231f
C596 VTAIL.n324 B 0.011989f
C597 VTAIL.n325 B 0.028336f
C598 VTAIL.n326 B 0.012694f
C599 VTAIL.n327 B 0.02231f
C600 VTAIL.n328 B 0.011989f
C601 VTAIL.n329 B 0.028336f
C602 VTAIL.n330 B 0.012694f
C603 VTAIL.n331 B 0.02231f
C604 VTAIL.n332 B 0.011989f
C605 VTAIL.n333 B 0.028336f
C606 VTAIL.n334 B 0.012694f
C607 VTAIL.n335 B 0.02231f
C608 VTAIL.n336 B 0.011989f
C609 VTAIL.n337 B 0.028336f
C610 VTAIL.n338 B 0.012694f
C611 VTAIL.n339 B 0.02231f
C612 VTAIL.n340 B 0.011989f
C613 VTAIL.n341 B 0.028336f
C614 VTAIL.n342 B 0.012341f
C615 VTAIL.n343 B 0.02231f
C616 VTAIL.n344 B 0.012694f
C617 VTAIL.n345 B 0.028336f
C618 VTAIL.n346 B 0.012694f
C619 VTAIL.n347 B 0.02231f
C620 VTAIL.n348 B 0.011989f
C621 VTAIL.n349 B 0.028336f
C622 VTAIL.n350 B 0.012694f
C623 VTAIL.n351 B 1.80128f
C624 VTAIL.n352 B 0.011989f
C625 VTAIL.t5 B 0.048676f
C626 VTAIL.n353 B 0.219182f
C627 VTAIL.n354 B 0.020032f
C628 VTAIL.n355 B 0.021252f
C629 VTAIL.n356 B 0.028336f
C630 VTAIL.n357 B 0.012694f
C631 VTAIL.n358 B 0.011989f
C632 VTAIL.n359 B 0.02231f
C633 VTAIL.n360 B 0.02231f
C634 VTAIL.n361 B 0.011989f
C635 VTAIL.n362 B 0.012694f
C636 VTAIL.n363 B 0.028336f
C637 VTAIL.n364 B 0.028336f
C638 VTAIL.n365 B 0.012694f
C639 VTAIL.n366 B 0.011989f
C640 VTAIL.n367 B 0.02231f
C641 VTAIL.n368 B 0.02231f
C642 VTAIL.n369 B 0.011989f
C643 VTAIL.n370 B 0.011989f
C644 VTAIL.n371 B 0.012694f
C645 VTAIL.n372 B 0.028336f
C646 VTAIL.n373 B 0.028336f
C647 VTAIL.n374 B 0.028336f
C648 VTAIL.n375 B 0.012341f
C649 VTAIL.n376 B 0.011989f
C650 VTAIL.n377 B 0.02231f
C651 VTAIL.n378 B 0.02231f
C652 VTAIL.n379 B 0.011989f
C653 VTAIL.n380 B 0.012694f
C654 VTAIL.n381 B 0.028336f
C655 VTAIL.n382 B 0.028336f
C656 VTAIL.n383 B 0.012694f
C657 VTAIL.n384 B 0.011989f
C658 VTAIL.n385 B 0.02231f
C659 VTAIL.n386 B 0.02231f
C660 VTAIL.n387 B 0.011989f
C661 VTAIL.n388 B 0.012694f
C662 VTAIL.n389 B 0.028336f
C663 VTAIL.n390 B 0.028336f
C664 VTAIL.n391 B 0.012694f
C665 VTAIL.n392 B 0.011989f
C666 VTAIL.n393 B 0.02231f
C667 VTAIL.n394 B 0.02231f
C668 VTAIL.n395 B 0.011989f
C669 VTAIL.n396 B 0.012694f
C670 VTAIL.n397 B 0.028336f
C671 VTAIL.n398 B 0.028336f
C672 VTAIL.n399 B 0.012694f
C673 VTAIL.n400 B 0.011989f
C674 VTAIL.n401 B 0.02231f
C675 VTAIL.n402 B 0.02231f
C676 VTAIL.n403 B 0.011989f
C677 VTAIL.n404 B 0.012694f
C678 VTAIL.n405 B 0.028336f
C679 VTAIL.n406 B 0.028336f
C680 VTAIL.n407 B 0.012694f
C681 VTAIL.n408 B 0.011989f
C682 VTAIL.n409 B 0.02231f
C683 VTAIL.n410 B 0.02231f
C684 VTAIL.n411 B 0.011989f
C685 VTAIL.n412 B 0.012694f
C686 VTAIL.n413 B 0.028336f
C687 VTAIL.n414 B 0.028336f
C688 VTAIL.n415 B 0.012694f
C689 VTAIL.n416 B 0.011989f
C690 VTAIL.n417 B 0.02231f
C691 VTAIL.n418 B 0.057969f
C692 VTAIL.n419 B 0.011989f
C693 VTAIL.n420 B 0.012694f
C694 VTAIL.n421 B 0.058415f
C695 VTAIL.n422 B 0.049332f
C696 VTAIL.n423 B 1.6908f
C697 VDD1.n0 B 0.012196f
C698 VDD1.n1 B 0.027464f
C699 VDD1.n2 B 0.012303f
C700 VDD1.n3 B 0.021623f
C701 VDD1.n4 B 0.011619f
C702 VDD1.n5 B 0.027464f
C703 VDD1.n6 B 0.012303f
C704 VDD1.n7 B 0.021623f
C705 VDD1.n8 B 0.011619f
C706 VDD1.n9 B 0.027464f
C707 VDD1.n10 B 0.012303f
C708 VDD1.n11 B 0.021623f
C709 VDD1.n12 B 0.011619f
C710 VDD1.n13 B 0.027464f
C711 VDD1.n14 B 0.012303f
C712 VDD1.n15 B 0.021623f
C713 VDD1.n16 B 0.011619f
C714 VDD1.n17 B 0.027464f
C715 VDD1.n18 B 0.012303f
C716 VDD1.n19 B 0.021623f
C717 VDD1.n20 B 0.011619f
C718 VDD1.n21 B 0.027464f
C719 VDD1.n22 B 0.011961f
C720 VDD1.n23 B 0.021623f
C721 VDD1.n24 B 0.011961f
C722 VDD1.n25 B 0.011619f
C723 VDD1.n26 B 0.027464f
C724 VDD1.n27 B 0.027464f
C725 VDD1.n28 B 0.012303f
C726 VDD1.n29 B 0.021623f
C727 VDD1.n30 B 0.011619f
C728 VDD1.n31 B 0.027464f
C729 VDD1.n32 B 0.012303f
C730 VDD1.n33 B 1.74582f
C731 VDD1.n34 B 0.011619f
C732 VDD1.t0 B 0.047178f
C733 VDD1.n35 B 0.212435f
C734 VDD1.n36 B 0.019415f
C735 VDD1.n37 B 0.020598f
C736 VDD1.n38 B 0.027464f
C737 VDD1.n39 B 0.012303f
C738 VDD1.n40 B 0.011619f
C739 VDD1.n41 B 0.021623f
C740 VDD1.n42 B 0.021623f
C741 VDD1.n43 B 0.011619f
C742 VDD1.n44 B 0.012303f
C743 VDD1.n45 B 0.027464f
C744 VDD1.n46 B 0.027464f
C745 VDD1.n47 B 0.012303f
C746 VDD1.n48 B 0.011619f
C747 VDD1.n49 B 0.021623f
C748 VDD1.n50 B 0.021623f
C749 VDD1.n51 B 0.011619f
C750 VDD1.n52 B 0.012303f
C751 VDD1.n53 B 0.027464f
C752 VDD1.n54 B 0.027464f
C753 VDD1.n55 B 0.012303f
C754 VDD1.n56 B 0.011619f
C755 VDD1.n57 B 0.021623f
C756 VDD1.n58 B 0.021623f
C757 VDD1.n59 B 0.011619f
C758 VDD1.n60 B 0.012303f
C759 VDD1.n61 B 0.027464f
C760 VDD1.n62 B 0.027464f
C761 VDD1.n63 B 0.012303f
C762 VDD1.n64 B 0.011619f
C763 VDD1.n65 B 0.021623f
C764 VDD1.n66 B 0.021623f
C765 VDD1.n67 B 0.011619f
C766 VDD1.n68 B 0.012303f
C767 VDD1.n69 B 0.027464f
C768 VDD1.n70 B 0.027464f
C769 VDD1.n71 B 0.012303f
C770 VDD1.n72 B 0.011619f
C771 VDD1.n73 B 0.021623f
C772 VDD1.n74 B 0.021623f
C773 VDD1.n75 B 0.011619f
C774 VDD1.n76 B 0.012303f
C775 VDD1.n77 B 0.027464f
C776 VDD1.n78 B 0.027464f
C777 VDD1.n79 B 0.012303f
C778 VDD1.n80 B 0.011619f
C779 VDD1.n81 B 0.021623f
C780 VDD1.n82 B 0.021623f
C781 VDD1.n83 B 0.011619f
C782 VDD1.n84 B 0.012303f
C783 VDD1.n85 B 0.027464f
C784 VDD1.n86 B 0.027464f
C785 VDD1.n87 B 0.012303f
C786 VDD1.n88 B 0.011619f
C787 VDD1.n89 B 0.021623f
C788 VDD1.n90 B 0.021623f
C789 VDD1.n91 B 0.011619f
C790 VDD1.n92 B 0.012303f
C791 VDD1.n93 B 0.027464f
C792 VDD1.n94 B 0.027464f
C793 VDD1.n95 B 0.012303f
C794 VDD1.n96 B 0.011619f
C795 VDD1.n97 B 0.021623f
C796 VDD1.n98 B 0.056184f
C797 VDD1.n99 B 0.011619f
C798 VDD1.n100 B 0.012303f
C799 VDD1.n101 B 0.056617f
C800 VDD1.n102 B 0.065866f
C801 VDD1.n103 B 0.012196f
C802 VDD1.n104 B 0.027464f
C803 VDD1.n105 B 0.012303f
C804 VDD1.n106 B 0.021623f
C805 VDD1.n107 B 0.011619f
C806 VDD1.n108 B 0.027464f
C807 VDD1.n109 B 0.012303f
C808 VDD1.n110 B 0.021623f
C809 VDD1.n111 B 0.011619f
C810 VDD1.n112 B 0.027464f
C811 VDD1.n113 B 0.012303f
C812 VDD1.n114 B 0.021623f
C813 VDD1.n115 B 0.011619f
C814 VDD1.n116 B 0.027464f
C815 VDD1.n117 B 0.012303f
C816 VDD1.n118 B 0.021623f
C817 VDD1.n119 B 0.011619f
C818 VDD1.n120 B 0.027464f
C819 VDD1.n121 B 0.012303f
C820 VDD1.n122 B 0.021623f
C821 VDD1.n123 B 0.011619f
C822 VDD1.n124 B 0.027464f
C823 VDD1.n125 B 0.011961f
C824 VDD1.n126 B 0.021623f
C825 VDD1.n127 B 0.012303f
C826 VDD1.n128 B 0.027464f
C827 VDD1.n129 B 0.012303f
C828 VDD1.n130 B 0.021623f
C829 VDD1.n131 B 0.011619f
C830 VDD1.n132 B 0.027464f
C831 VDD1.n133 B 0.012303f
C832 VDD1.n134 B 1.74582f
C833 VDD1.n135 B 0.011619f
C834 VDD1.t1 B 0.047178f
C835 VDD1.n136 B 0.212435f
C836 VDD1.n137 B 0.019415f
C837 VDD1.n138 B 0.020598f
C838 VDD1.n139 B 0.027464f
C839 VDD1.n140 B 0.012303f
C840 VDD1.n141 B 0.011619f
C841 VDD1.n142 B 0.021623f
C842 VDD1.n143 B 0.021623f
C843 VDD1.n144 B 0.011619f
C844 VDD1.n145 B 0.012303f
C845 VDD1.n146 B 0.027464f
C846 VDD1.n147 B 0.027464f
C847 VDD1.n148 B 0.012303f
C848 VDD1.n149 B 0.011619f
C849 VDD1.n150 B 0.021623f
C850 VDD1.n151 B 0.021623f
C851 VDD1.n152 B 0.011619f
C852 VDD1.n153 B 0.011619f
C853 VDD1.n154 B 0.012303f
C854 VDD1.n155 B 0.027464f
C855 VDD1.n156 B 0.027464f
C856 VDD1.n157 B 0.027464f
C857 VDD1.n158 B 0.011961f
C858 VDD1.n159 B 0.011619f
C859 VDD1.n160 B 0.021623f
C860 VDD1.n161 B 0.021623f
C861 VDD1.n162 B 0.011619f
C862 VDD1.n163 B 0.012303f
C863 VDD1.n164 B 0.027464f
C864 VDD1.n165 B 0.027464f
C865 VDD1.n166 B 0.012303f
C866 VDD1.n167 B 0.011619f
C867 VDD1.n168 B 0.021623f
C868 VDD1.n169 B 0.021623f
C869 VDD1.n170 B 0.011619f
C870 VDD1.n171 B 0.012303f
C871 VDD1.n172 B 0.027464f
C872 VDD1.n173 B 0.027464f
C873 VDD1.n174 B 0.012303f
C874 VDD1.n175 B 0.011619f
C875 VDD1.n176 B 0.021623f
C876 VDD1.n177 B 0.021623f
C877 VDD1.n178 B 0.011619f
C878 VDD1.n179 B 0.012303f
C879 VDD1.n180 B 0.027464f
C880 VDD1.n181 B 0.027464f
C881 VDD1.n182 B 0.012303f
C882 VDD1.n183 B 0.011619f
C883 VDD1.n184 B 0.021623f
C884 VDD1.n185 B 0.021623f
C885 VDD1.n186 B 0.011619f
C886 VDD1.n187 B 0.012303f
C887 VDD1.n188 B 0.027464f
C888 VDD1.n189 B 0.027464f
C889 VDD1.n190 B 0.012303f
C890 VDD1.n191 B 0.011619f
C891 VDD1.n192 B 0.021623f
C892 VDD1.n193 B 0.021623f
C893 VDD1.n194 B 0.011619f
C894 VDD1.n195 B 0.012303f
C895 VDD1.n196 B 0.027464f
C896 VDD1.n197 B 0.027464f
C897 VDD1.n198 B 0.012303f
C898 VDD1.n199 B 0.011619f
C899 VDD1.n200 B 0.021623f
C900 VDD1.n201 B 0.056184f
C901 VDD1.n202 B 0.011619f
C902 VDD1.n203 B 0.012303f
C903 VDD1.n204 B 0.056617f
C904 VDD1.n205 B 0.065428f
C905 VDD1.t2 B 0.321413f
C906 VDD1.t4 B 0.321413f
C907 VDD1.n206 B 2.94327f
C908 VDD1.n207 B 2.37354f
C909 VDD1.t3 B 0.321413f
C910 VDD1.t5 B 0.321413f
C911 VDD1.n208 B 2.94153f
C912 VDD1.n209 B 2.59928f
C913 VP.n0 B 0.031319f
C914 VP.t5 B 2.51361f
C915 VP.n1 B 0.040483f
C916 VP.n2 B 0.031319f
C917 VP.t1 B 2.51361f
C918 VP.n3 B 0.050956f
C919 VP.n4 B 0.031319f
C920 VP.t4 B 2.51361f
C921 VP.n5 B 0.040483f
C922 VP.t3 B 2.61217f
C923 VP.n6 B 0.961233f
C924 VP.t0 B 2.51361f
C925 VP.n7 B 0.94137f
C926 VP.n8 B 0.043961f
C927 VP.n9 B 0.197542f
C928 VP.n10 B 0.031319f
C929 VP.n11 B 0.031319f
C930 VP.n12 B 0.050956f
C931 VP.n13 B 0.037045f
C932 VP.n14 B 0.943612f
C933 VP.n15 B 1.6891f
C934 VP.n16 B 1.7118f
C935 VP.t2 B 2.51361f
C936 VP.n17 B 0.943612f
C937 VP.n18 B 0.037045f
C938 VP.n19 B 0.031319f
C939 VP.n20 B 0.031319f
C940 VP.n21 B 0.031319f
C941 VP.n22 B 0.040483f
C942 VP.n23 B 0.043961f
C943 VP.n24 B 0.881805f
C944 VP.n25 B 0.043961f
C945 VP.n26 B 0.031319f
C946 VP.n27 B 0.031319f
C947 VP.n28 B 0.031319f
C948 VP.n29 B 0.050956f
C949 VP.n30 B 0.037045f
C950 VP.n31 B 0.943612f
C951 VP.n32 B 0.031208f
.ends

