* NGSPICE file created from diff_pair_sample_0824.ext - technology: sky130A

.subckt diff_pair_sample_0824 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=0 ps=0 w=12.57 l=2.34
X1 VTAIL.t15 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X2 VTAIL.t14 VN.t1 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X3 VTAIL.t13 VN.t2 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=2.07405 ps=12.9 w=12.57 l=2.34
X4 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=0 ps=0 w=12.57 l=2.34
X5 VTAIL.t0 VP.t0 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X6 VTAIL.t12 VN.t3 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=2.07405 ps=12.9 w=12.57 l=2.34
X7 VTAIL.t1 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X8 VDD2.t7 VN.t4 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X9 VTAIL.t2 VP.t2 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=2.07405 ps=12.9 w=12.57 l=2.34
X10 VTAIL.t5 VP.t3 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=2.07405 ps=12.9 w=12.57 l=2.34
X11 VDD2.t6 VN.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=4.9023 ps=25.92 w=12.57 l=2.34
X12 VDD2.t5 VN.t6 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=4.9023 ps=25.92 w=12.57 l=2.34
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=0 ps=0 w=12.57 l=2.34
X14 VDD1.t3 VP.t4 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=4.9023 ps=25.92 w=12.57 l=2.34
X15 VDD1.t2 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=4.9023 ps=25.92 w=12.57 l=2.34
X16 VDD1.t1 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X17 VDD1.t0 VP.t7 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X18 VDD2.t2 VN.t7 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.07405 pd=12.9 as=2.07405 ps=12.9 w=12.57 l=2.34
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.9023 pd=25.92 as=0 ps=0 w=12.57 l=2.34
R0 B.n869 B.n868 585
R1 B.n328 B.n136 585
R2 B.n327 B.n326 585
R3 B.n325 B.n324 585
R4 B.n323 B.n322 585
R5 B.n321 B.n320 585
R6 B.n319 B.n318 585
R7 B.n317 B.n316 585
R8 B.n315 B.n314 585
R9 B.n313 B.n312 585
R10 B.n311 B.n310 585
R11 B.n309 B.n308 585
R12 B.n307 B.n306 585
R13 B.n305 B.n304 585
R14 B.n303 B.n302 585
R15 B.n301 B.n300 585
R16 B.n299 B.n298 585
R17 B.n297 B.n296 585
R18 B.n295 B.n294 585
R19 B.n293 B.n292 585
R20 B.n291 B.n290 585
R21 B.n289 B.n288 585
R22 B.n287 B.n286 585
R23 B.n285 B.n284 585
R24 B.n283 B.n282 585
R25 B.n281 B.n280 585
R26 B.n279 B.n278 585
R27 B.n277 B.n276 585
R28 B.n275 B.n274 585
R29 B.n273 B.n272 585
R30 B.n271 B.n270 585
R31 B.n269 B.n268 585
R32 B.n267 B.n266 585
R33 B.n265 B.n264 585
R34 B.n263 B.n262 585
R35 B.n261 B.n260 585
R36 B.n259 B.n258 585
R37 B.n257 B.n256 585
R38 B.n255 B.n254 585
R39 B.n253 B.n252 585
R40 B.n251 B.n250 585
R41 B.n249 B.n248 585
R42 B.n247 B.n246 585
R43 B.n244 B.n243 585
R44 B.n242 B.n241 585
R45 B.n240 B.n239 585
R46 B.n238 B.n237 585
R47 B.n236 B.n235 585
R48 B.n234 B.n233 585
R49 B.n232 B.n231 585
R50 B.n230 B.n229 585
R51 B.n228 B.n227 585
R52 B.n226 B.n225 585
R53 B.n223 B.n222 585
R54 B.n221 B.n220 585
R55 B.n219 B.n218 585
R56 B.n217 B.n216 585
R57 B.n215 B.n214 585
R58 B.n213 B.n212 585
R59 B.n211 B.n210 585
R60 B.n209 B.n208 585
R61 B.n207 B.n206 585
R62 B.n205 B.n204 585
R63 B.n203 B.n202 585
R64 B.n201 B.n200 585
R65 B.n199 B.n198 585
R66 B.n197 B.n196 585
R67 B.n195 B.n194 585
R68 B.n193 B.n192 585
R69 B.n191 B.n190 585
R70 B.n189 B.n188 585
R71 B.n187 B.n186 585
R72 B.n185 B.n184 585
R73 B.n183 B.n182 585
R74 B.n181 B.n180 585
R75 B.n179 B.n178 585
R76 B.n177 B.n176 585
R77 B.n175 B.n174 585
R78 B.n173 B.n172 585
R79 B.n171 B.n170 585
R80 B.n169 B.n168 585
R81 B.n167 B.n166 585
R82 B.n165 B.n164 585
R83 B.n163 B.n162 585
R84 B.n161 B.n160 585
R85 B.n159 B.n158 585
R86 B.n157 B.n156 585
R87 B.n155 B.n154 585
R88 B.n153 B.n152 585
R89 B.n151 B.n150 585
R90 B.n149 B.n148 585
R91 B.n147 B.n146 585
R92 B.n145 B.n144 585
R93 B.n143 B.n142 585
R94 B.n89 B.n88 585
R95 B.n874 B.n873 585
R96 B.n867 B.n137 585
R97 B.n137 B.n86 585
R98 B.n866 B.n85 585
R99 B.n878 B.n85 585
R100 B.n865 B.n84 585
R101 B.n879 B.n84 585
R102 B.n864 B.n83 585
R103 B.n880 B.n83 585
R104 B.n863 B.n862 585
R105 B.n862 B.n79 585
R106 B.n861 B.n78 585
R107 B.n886 B.n78 585
R108 B.n860 B.n77 585
R109 B.n887 B.n77 585
R110 B.n859 B.n76 585
R111 B.n888 B.n76 585
R112 B.n858 B.n857 585
R113 B.n857 B.n72 585
R114 B.n856 B.n71 585
R115 B.n894 B.n71 585
R116 B.n855 B.n70 585
R117 B.n895 B.n70 585
R118 B.n854 B.n69 585
R119 B.n896 B.n69 585
R120 B.n853 B.n852 585
R121 B.n852 B.n65 585
R122 B.n851 B.n64 585
R123 B.n902 B.n64 585
R124 B.n850 B.n63 585
R125 B.n903 B.n63 585
R126 B.n849 B.n62 585
R127 B.n904 B.n62 585
R128 B.n848 B.n847 585
R129 B.n847 B.n58 585
R130 B.n846 B.n57 585
R131 B.n910 B.n57 585
R132 B.n845 B.n56 585
R133 B.n911 B.n56 585
R134 B.n844 B.n55 585
R135 B.n912 B.n55 585
R136 B.n843 B.n842 585
R137 B.n842 B.n51 585
R138 B.n841 B.n50 585
R139 B.n918 B.n50 585
R140 B.n840 B.n49 585
R141 B.n919 B.n49 585
R142 B.n839 B.n48 585
R143 B.n920 B.n48 585
R144 B.n838 B.n837 585
R145 B.n837 B.n44 585
R146 B.n836 B.n43 585
R147 B.n926 B.n43 585
R148 B.n835 B.n42 585
R149 B.n927 B.n42 585
R150 B.n834 B.n41 585
R151 B.n928 B.n41 585
R152 B.n833 B.n832 585
R153 B.n832 B.n37 585
R154 B.n831 B.n36 585
R155 B.n934 B.n36 585
R156 B.n830 B.n35 585
R157 B.n935 B.n35 585
R158 B.n829 B.n34 585
R159 B.n936 B.n34 585
R160 B.n828 B.n827 585
R161 B.n827 B.n30 585
R162 B.n826 B.n29 585
R163 B.n942 B.n29 585
R164 B.n825 B.n28 585
R165 B.n943 B.n28 585
R166 B.n824 B.n27 585
R167 B.n944 B.n27 585
R168 B.n823 B.n822 585
R169 B.n822 B.n23 585
R170 B.n821 B.n22 585
R171 B.n950 B.n22 585
R172 B.n820 B.n21 585
R173 B.n951 B.n21 585
R174 B.n819 B.n20 585
R175 B.n952 B.n20 585
R176 B.n818 B.n817 585
R177 B.n817 B.n16 585
R178 B.n816 B.n15 585
R179 B.n958 B.n15 585
R180 B.n815 B.n14 585
R181 B.n959 B.n14 585
R182 B.n814 B.n13 585
R183 B.n960 B.n13 585
R184 B.n813 B.n812 585
R185 B.n812 B.n12 585
R186 B.n811 B.n810 585
R187 B.n811 B.n8 585
R188 B.n809 B.n7 585
R189 B.n967 B.n7 585
R190 B.n808 B.n6 585
R191 B.n968 B.n6 585
R192 B.n807 B.n5 585
R193 B.n969 B.n5 585
R194 B.n806 B.n805 585
R195 B.n805 B.n4 585
R196 B.n804 B.n329 585
R197 B.n804 B.n803 585
R198 B.n794 B.n330 585
R199 B.n331 B.n330 585
R200 B.n796 B.n795 585
R201 B.n797 B.n796 585
R202 B.n793 B.n336 585
R203 B.n336 B.n335 585
R204 B.n792 B.n791 585
R205 B.n791 B.n790 585
R206 B.n338 B.n337 585
R207 B.n339 B.n338 585
R208 B.n783 B.n782 585
R209 B.n784 B.n783 585
R210 B.n781 B.n344 585
R211 B.n344 B.n343 585
R212 B.n780 B.n779 585
R213 B.n779 B.n778 585
R214 B.n346 B.n345 585
R215 B.n347 B.n346 585
R216 B.n771 B.n770 585
R217 B.n772 B.n771 585
R218 B.n769 B.n351 585
R219 B.n355 B.n351 585
R220 B.n768 B.n767 585
R221 B.n767 B.n766 585
R222 B.n353 B.n352 585
R223 B.n354 B.n353 585
R224 B.n759 B.n758 585
R225 B.n760 B.n759 585
R226 B.n757 B.n360 585
R227 B.n360 B.n359 585
R228 B.n756 B.n755 585
R229 B.n755 B.n754 585
R230 B.n362 B.n361 585
R231 B.n363 B.n362 585
R232 B.n747 B.n746 585
R233 B.n748 B.n747 585
R234 B.n745 B.n367 585
R235 B.n371 B.n367 585
R236 B.n744 B.n743 585
R237 B.n743 B.n742 585
R238 B.n369 B.n368 585
R239 B.n370 B.n369 585
R240 B.n735 B.n734 585
R241 B.n736 B.n735 585
R242 B.n733 B.n376 585
R243 B.n376 B.n375 585
R244 B.n732 B.n731 585
R245 B.n731 B.n730 585
R246 B.n378 B.n377 585
R247 B.n379 B.n378 585
R248 B.n723 B.n722 585
R249 B.n724 B.n723 585
R250 B.n721 B.n383 585
R251 B.n387 B.n383 585
R252 B.n720 B.n719 585
R253 B.n719 B.n718 585
R254 B.n385 B.n384 585
R255 B.n386 B.n385 585
R256 B.n711 B.n710 585
R257 B.n712 B.n711 585
R258 B.n709 B.n392 585
R259 B.n392 B.n391 585
R260 B.n708 B.n707 585
R261 B.n707 B.n706 585
R262 B.n394 B.n393 585
R263 B.n395 B.n394 585
R264 B.n699 B.n698 585
R265 B.n700 B.n699 585
R266 B.n697 B.n400 585
R267 B.n400 B.n399 585
R268 B.n696 B.n695 585
R269 B.n695 B.n694 585
R270 B.n402 B.n401 585
R271 B.n403 B.n402 585
R272 B.n687 B.n686 585
R273 B.n688 B.n687 585
R274 B.n685 B.n408 585
R275 B.n408 B.n407 585
R276 B.n684 B.n683 585
R277 B.n683 B.n682 585
R278 B.n410 B.n409 585
R279 B.n411 B.n410 585
R280 B.n675 B.n674 585
R281 B.n676 B.n675 585
R282 B.n673 B.n416 585
R283 B.n416 B.n415 585
R284 B.n672 B.n671 585
R285 B.n671 B.n670 585
R286 B.n418 B.n417 585
R287 B.n419 B.n418 585
R288 B.n666 B.n665 585
R289 B.n422 B.n421 585
R290 B.n662 B.n661 585
R291 B.n663 B.n662 585
R292 B.n660 B.n470 585
R293 B.n659 B.n658 585
R294 B.n657 B.n656 585
R295 B.n655 B.n654 585
R296 B.n653 B.n652 585
R297 B.n651 B.n650 585
R298 B.n649 B.n648 585
R299 B.n647 B.n646 585
R300 B.n645 B.n644 585
R301 B.n643 B.n642 585
R302 B.n641 B.n640 585
R303 B.n639 B.n638 585
R304 B.n637 B.n636 585
R305 B.n635 B.n634 585
R306 B.n633 B.n632 585
R307 B.n631 B.n630 585
R308 B.n629 B.n628 585
R309 B.n627 B.n626 585
R310 B.n625 B.n624 585
R311 B.n623 B.n622 585
R312 B.n621 B.n620 585
R313 B.n619 B.n618 585
R314 B.n617 B.n616 585
R315 B.n615 B.n614 585
R316 B.n613 B.n612 585
R317 B.n611 B.n610 585
R318 B.n609 B.n608 585
R319 B.n607 B.n606 585
R320 B.n605 B.n604 585
R321 B.n603 B.n602 585
R322 B.n601 B.n600 585
R323 B.n599 B.n598 585
R324 B.n597 B.n596 585
R325 B.n595 B.n594 585
R326 B.n593 B.n592 585
R327 B.n591 B.n590 585
R328 B.n589 B.n588 585
R329 B.n587 B.n586 585
R330 B.n585 B.n584 585
R331 B.n583 B.n582 585
R332 B.n581 B.n580 585
R333 B.n579 B.n578 585
R334 B.n577 B.n576 585
R335 B.n575 B.n574 585
R336 B.n573 B.n572 585
R337 B.n571 B.n570 585
R338 B.n569 B.n568 585
R339 B.n567 B.n566 585
R340 B.n565 B.n564 585
R341 B.n563 B.n562 585
R342 B.n561 B.n560 585
R343 B.n559 B.n558 585
R344 B.n557 B.n556 585
R345 B.n555 B.n554 585
R346 B.n553 B.n552 585
R347 B.n551 B.n550 585
R348 B.n549 B.n548 585
R349 B.n547 B.n546 585
R350 B.n545 B.n544 585
R351 B.n543 B.n542 585
R352 B.n541 B.n540 585
R353 B.n539 B.n538 585
R354 B.n537 B.n536 585
R355 B.n535 B.n534 585
R356 B.n533 B.n532 585
R357 B.n531 B.n530 585
R358 B.n529 B.n528 585
R359 B.n527 B.n526 585
R360 B.n525 B.n524 585
R361 B.n523 B.n522 585
R362 B.n521 B.n520 585
R363 B.n519 B.n518 585
R364 B.n517 B.n516 585
R365 B.n515 B.n514 585
R366 B.n513 B.n512 585
R367 B.n511 B.n510 585
R368 B.n509 B.n508 585
R369 B.n507 B.n506 585
R370 B.n505 B.n504 585
R371 B.n503 B.n502 585
R372 B.n501 B.n500 585
R373 B.n499 B.n498 585
R374 B.n497 B.n496 585
R375 B.n495 B.n494 585
R376 B.n493 B.n492 585
R377 B.n491 B.n490 585
R378 B.n489 B.n488 585
R379 B.n487 B.n486 585
R380 B.n485 B.n484 585
R381 B.n483 B.n482 585
R382 B.n481 B.n480 585
R383 B.n479 B.n478 585
R384 B.n477 B.n469 585
R385 B.n663 B.n469 585
R386 B.n667 B.n420 585
R387 B.n420 B.n419 585
R388 B.n669 B.n668 585
R389 B.n670 B.n669 585
R390 B.n414 B.n413 585
R391 B.n415 B.n414 585
R392 B.n678 B.n677 585
R393 B.n677 B.n676 585
R394 B.n679 B.n412 585
R395 B.n412 B.n411 585
R396 B.n681 B.n680 585
R397 B.n682 B.n681 585
R398 B.n406 B.n405 585
R399 B.n407 B.n406 585
R400 B.n690 B.n689 585
R401 B.n689 B.n688 585
R402 B.n691 B.n404 585
R403 B.n404 B.n403 585
R404 B.n693 B.n692 585
R405 B.n694 B.n693 585
R406 B.n398 B.n397 585
R407 B.n399 B.n398 585
R408 B.n702 B.n701 585
R409 B.n701 B.n700 585
R410 B.n703 B.n396 585
R411 B.n396 B.n395 585
R412 B.n705 B.n704 585
R413 B.n706 B.n705 585
R414 B.n390 B.n389 585
R415 B.n391 B.n390 585
R416 B.n714 B.n713 585
R417 B.n713 B.n712 585
R418 B.n715 B.n388 585
R419 B.n388 B.n386 585
R420 B.n717 B.n716 585
R421 B.n718 B.n717 585
R422 B.n382 B.n381 585
R423 B.n387 B.n382 585
R424 B.n726 B.n725 585
R425 B.n725 B.n724 585
R426 B.n727 B.n380 585
R427 B.n380 B.n379 585
R428 B.n729 B.n728 585
R429 B.n730 B.n729 585
R430 B.n374 B.n373 585
R431 B.n375 B.n374 585
R432 B.n738 B.n737 585
R433 B.n737 B.n736 585
R434 B.n739 B.n372 585
R435 B.n372 B.n370 585
R436 B.n741 B.n740 585
R437 B.n742 B.n741 585
R438 B.n366 B.n365 585
R439 B.n371 B.n366 585
R440 B.n750 B.n749 585
R441 B.n749 B.n748 585
R442 B.n751 B.n364 585
R443 B.n364 B.n363 585
R444 B.n753 B.n752 585
R445 B.n754 B.n753 585
R446 B.n358 B.n357 585
R447 B.n359 B.n358 585
R448 B.n762 B.n761 585
R449 B.n761 B.n760 585
R450 B.n763 B.n356 585
R451 B.n356 B.n354 585
R452 B.n765 B.n764 585
R453 B.n766 B.n765 585
R454 B.n350 B.n349 585
R455 B.n355 B.n350 585
R456 B.n774 B.n773 585
R457 B.n773 B.n772 585
R458 B.n775 B.n348 585
R459 B.n348 B.n347 585
R460 B.n777 B.n776 585
R461 B.n778 B.n777 585
R462 B.n342 B.n341 585
R463 B.n343 B.n342 585
R464 B.n786 B.n785 585
R465 B.n785 B.n784 585
R466 B.n787 B.n340 585
R467 B.n340 B.n339 585
R468 B.n789 B.n788 585
R469 B.n790 B.n789 585
R470 B.n334 B.n333 585
R471 B.n335 B.n334 585
R472 B.n799 B.n798 585
R473 B.n798 B.n797 585
R474 B.n800 B.n332 585
R475 B.n332 B.n331 585
R476 B.n802 B.n801 585
R477 B.n803 B.n802 585
R478 B.n3 B.n0 585
R479 B.n4 B.n3 585
R480 B.n966 B.n1 585
R481 B.n967 B.n966 585
R482 B.n965 B.n964 585
R483 B.n965 B.n8 585
R484 B.n963 B.n9 585
R485 B.n12 B.n9 585
R486 B.n962 B.n961 585
R487 B.n961 B.n960 585
R488 B.n11 B.n10 585
R489 B.n959 B.n11 585
R490 B.n957 B.n956 585
R491 B.n958 B.n957 585
R492 B.n955 B.n17 585
R493 B.n17 B.n16 585
R494 B.n954 B.n953 585
R495 B.n953 B.n952 585
R496 B.n19 B.n18 585
R497 B.n951 B.n19 585
R498 B.n949 B.n948 585
R499 B.n950 B.n949 585
R500 B.n947 B.n24 585
R501 B.n24 B.n23 585
R502 B.n946 B.n945 585
R503 B.n945 B.n944 585
R504 B.n26 B.n25 585
R505 B.n943 B.n26 585
R506 B.n941 B.n940 585
R507 B.n942 B.n941 585
R508 B.n939 B.n31 585
R509 B.n31 B.n30 585
R510 B.n938 B.n937 585
R511 B.n937 B.n936 585
R512 B.n33 B.n32 585
R513 B.n935 B.n33 585
R514 B.n933 B.n932 585
R515 B.n934 B.n933 585
R516 B.n931 B.n38 585
R517 B.n38 B.n37 585
R518 B.n930 B.n929 585
R519 B.n929 B.n928 585
R520 B.n40 B.n39 585
R521 B.n927 B.n40 585
R522 B.n925 B.n924 585
R523 B.n926 B.n925 585
R524 B.n923 B.n45 585
R525 B.n45 B.n44 585
R526 B.n922 B.n921 585
R527 B.n921 B.n920 585
R528 B.n47 B.n46 585
R529 B.n919 B.n47 585
R530 B.n917 B.n916 585
R531 B.n918 B.n917 585
R532 B.n915 B.n52 585
R533 B.n52 B.n51 585
R534 B.n914 B.n913 585
R535 B.n913 B.n912 585
R536 B.n54 B.n53 585
R537 B.n911 B.n54 585
R538 B.n909 B.n908 585
R539 B.n910 B.n909 585
R540 B.n907 B.n59 585
R541 B.n59 B.n58 585
R542 B.n906 B.n905 585
R543 B.n905 B.n904 585
R544 B.n61 B.n60 585
R545 B.n903 B.n61 585
R546 B.n901 B.n900 585
R547 B.n902 B.n901 585
R548 B.n899 B.n66 585
R549 B.n66 B.n65 585
R550 B.n898 B.n897 585
R551 B.n897 B.n896 585
R552 B.n68 B.n67 585
R553 B.n895 B.n68 585
R554 B.n893 B.n892 585
R555 B.n894 B.n893 585
R556 B.n891 B.n73 585
R557 B.n73 B.n72 585
R558 B.n890 B.n889 585
R559 B.n889 B.n888 585
R560 B.n75 B.n74 585
R561 B.n887 B.n75 585
R562 B.n885 B.n884 585
R563 B.n886 B.n885 585
R564 B.n883 B.n80 585
R565 B.n80 B.n79 585
R566 B.n882 B.n881 585
R567 B.n881 B.n880 585
R568 B.n82 B.n81 585
R569 B.n879 B.n82 585
R570 B.n877 B.n876 585
R571 B.n878 B.n877 585
R572 B.n875 B.n87 585
R573 B.n87 B.n86 585
R574 B.n970 B.n969 585
R575 B.n968 B.n2 585
R576 B.n873 B.n87 492.5
R577 B.n869 B.n137 492.5
R578 B.n469 B.n418 492.5
R579 B.n665 B.n420 492.5
R580 B.n140 B.t12 337.079
R581 B.n138 B.t16 337.079
R582 B.n474 B.t8 337.079
R583 B.n471 B.t19 337.079
R584 B.n871 B.n870 256.663
R585 B.n871 B.n135 256.663
R586 B.n871 B.n134 256.663
R587 B.n871 B.n133 256.663
R588 B.n871 B.n132 256.663
R589 B.n871 B.n131 256.663
R590 B.n871 B.n130 256.663
R591 B.n871 B.n129 256.663
R592 B.n871 B.n128 256.663
R593 B.n871 B.n127 256.663
R594 B.n871 B.n126 256.663
R595 B.n871 B.n125 256.663
R596 B.n871 B.n124 256.663
R597 B.n871 B.n123 256.663
R598 B.n871 B.n122 256.663
R599 B.n871 B.n121 256.663
R600 B.n871 B.n120 256.663
R601 B.n871 B.n119 256.663
R602 B.n871 B.n118 256.663
R603 B.n871 B.n117 256.663
R604 B.n871 B.n116 256.663
R605 B.n871 B.n115 256.663
R606 B.n871 B.n114 256.663
R607 B.n871 B.n113 256.663
R608 B.n871 B.n112 256.663
R609 B.n871 B.n111 256.663
R610 B.n871 B.n110 256.663
R611 B.n871 B.n109 256.663
R612 B.n871 B.n108 256.663
R613 B.n871 B.n107 256.663
R614 B.n871 B.n106 256.663
R615 B.n871 B.n105 256.663
R616 B.n871 B.n104 256.663
R617 B.n871 B.n103 256.663
R618 B.n871 B.n102 256.663
R619 B.n871 B.n101 256.663
R620 B.n871 B.n100 256.663
R621 B.n871 B.n99 256.663
R622 B.n871 B.n98 256.663
R623 B.n871 B.n97 256.663
R624 B.n871 B.n96 256.663
R625 B.n871 B.n95 256.663
R626 B.n871 B.n94 256.663
R627 B.n871 B.n93 256.663
R628 B.n871 B.n92 256.663
R629 B.n871 B.n91 256.663
R630 B.n871 B.n90 256.663
R631 B.n872 B.n871 256.663
R632 B.n664 B.n663 256.663
R633 B.n663 B.n423 256.663
R634 B.n663 B.n424 256.663
R635 B.n663 B.n425 256.663
R636 B.n663 B.n426 256.663
R637 B.n663 B.n427 256.663
R638 B.n663 B.n428 256.663
R639 B.n663 B.n429 256.663
R640 B.n663 B.n430 256.663
R641 B.n663 B.n431 256.663
R642 B.n663 B.n432 256.663
R643 B.n663 B.n433 256.663
R644 B.n663 B.n434 256.663
R645 B.n663 B.n435 256.663
R646 B.n663 B.n436 256.663
R647 B.n663 B.n437 256.663
R648 B.n663 B.n438 256.663
R649 B.n663 B.n439 256.663
R650 B.n663 B.n440 256.663
R651 B.n663 B.n441 256.663
R652 B.n663 B.n442 256.663
R653 B.n663 B.n443 256.663
R654 B.n663 B.n444 256.663
R655 B.n663 B.n445 256.663
R656 B.n663 B.n446 256.663
R657 B.n663 B.n447 256.663
R658 B.n663 B.n448 256.663
R659 B.n663 B.n449 256.663
R660 B.n663 B.n450 256.663
R661 B.n663 B.n451 256.663
R662 B.n663 B.n452 256.663
R663 B.n663 B.n453 256.663
R664 B.n663 B.n454 256.663
R665 B.n663 B.n455 256.663
R666 B.n663 B.n456 256.663
R667 B.n663 B.n457 256.663
R668 B.n663 B.n458 256.663
R669 B.n663 B.n459 256.663
R670 B.n663 B.n460 256.663
R671 B.n663 B.n461 256.663
R672 B.n663 B.n462 256.663
R673 B.n663 B.n463 256.663
R674 B.n663 B.n464 256.663
R675 B.n663 B.n465 256.663
R676 B.n663 B.n466 256.663
R677 B.n663 B.n467 256.663
R678 B.n663 B.n468 256.663
R679 B.n972 B.n971 256.663
R680 B.n142 B.n89 163.367
R681 B.n146 B.n145 163.367
R682 B.n150 B.n149 163.367
R683 B.n154 B.n153 163.367
R684 B.n158 B.n157 163.367
R685 B.n162 B.n161 163.367
R686 B.n166 B.n165 163.367
R687 B.n170 B.n169 163.367
R688 B.n174 B.n173 163.367
R689 B.n178 B.n177 163.367
R690 B.n182 B.n181 163.367
R691 B.n186 B.n185 163.367
R692 B.n190 B.n189 163.367
R693 B.n194 B.n193 163.367
R694 B.n198 B.n197 163.367
R695 B.n202 B.n201 163.367
R696 B.n206 B.n205 163.367
R697 B.n210 B.n209 163.367
R698 B.n214 B.n213 163.367
R699 B.n218 B.n217 163.367
R700 B.n222 B.n221 163.367
R701 B.n227 B.n226 163.367
R702 B.n231 B.n230 163.367
R703 B.n235 B.n234 163.367
R704 B.n239 B.n238 163.367
R705 B.n243 B.n242 163.367
R706 B.n248 B.n247 163.367
R707 B.n252 B.n251 163.367
R708 B.n256 B.n255 163.367
R709 B.n260 B.n259 163.367
R710 B.n264 B.n263 163.367
R711 B.n268 B.n267 163.367
R712 B.n272 B.n271 163.367
R713 B.n276 B.n275 163.367
R714 B.n280 B.n279 163.367
R715 B.n284 B.n283 163.367
R716 B.n288 B.n287 163.367
R717 B.n292 B.n291 163.367
R718 B.n296 B.n295 163.367
R719 B.n300 B.n299 163.367
R720 B.n304 B.n303 163.367
R721 B.n308 B.n307 163.367
R722 B.n312 B.n311 163.367
R723 B.n316 B.n315 163.367
R724 B.n320 B.n319 163.367
R725 B.n324 B.n323 163.367
R726 B.n326 B.n136 163.367
R727 B.n671 B.n418 163.367
R728 B.n671 B.n416 163.367
R729 B.n675 B.n416 163.367
R730 B.n675 B.n410 163.367
R731 B.n683 B.n410 163.367
R732 B.n683 B.n408 163.367
R733 B.n687 B.n408 163.367
R734 B.n687 B.n402 163.367
R735 B.n695 B.n402 163.367
R736 B.n695 B.n400 163.367
R737 B.n699 B.n400 163.367
R738 B.n699 B.n394 163.367
R739 B.n707 B.n394 163.367
R740 B.n707 B.n392 163.367
R741 B.n711 B.n392 163.367
R742 B.n711 B.n385 163.367
R743 B.n719 B.n385 163.367
R744 B.n719 B.n383 163.367
R745 B.n723 B.n383 163.367
R746 B.n723 B.n378 163.367
R747 B.n731 B.n378 163.367
R748 B.n731 B.n376 163.367
R749 B.n735 B.n376 163.367
R750 B.n735 B.n369 163.367
R751 B.n743 B.n369 163.367
R752 B.n743 B.n367 163.367
R753 B.n747 B.n367 163.367
R754 B.n747 B.n362 163.367
R755 B.n755 B.n362 163.367
R756 B.n755 B.n360 163.367
R757 B.n759 B.n360 163.367
R758 B.n759 B.n353 163.367
R759 B.n767 B.n353 163.367
R760 B.n767 B.n351 163.367
R761 B.n771 B.n351 163.367
R762 B.n771 B.n346 163.367
R763 B.n779 B.n346 163.367
R764 B.n779 B.n344 163.367
R765 B.n783 B.n344 163.367
R766 B.n783 B.n338 163.367
R767 B.n791 B.n338 163.367
R768 B.n791 B.n336 163.367
R769 B.n796 B.n336 163.367
R770 B.n796 B.n330 163.367
R771 B.n804 B.n330 163.367
R772 B.n805 B.n804 163.367
R773 B.n805 B.n5 163.367
R774 B.n6 B.n5 163.367
R775 B.n7 B.n6 163.367
R776 B.n811 B.n7 163.367
R777 B.n812 B.n811 163.367
R778 B.n812 B.n13 163.367
R779 B.n14 B.n13 163.367
R780 B.n15 B.n14 163.367
R781 B.n817 B.n15 163.367
R782 B.n817 B.n20 163.367
R783 B.n21 B.n20 163.367
R784 B.n22 B.n21 163.367
R785 B.n822 B.n22 163.367
R786 B.n822 B.n27 163.367
R787 B.n28 B.n27 163.367
R788 B.n29 B.n28 163.367
R789 B.n827 B.n29 163.367
R790 B.n827 B.n34 163.367
R791 B.n35 B.n34 163.367
R792 B.n36 B.n35 163.367
R793 B.n832 B.n36 163.367
R794 B.n832 B.n41 163.367
R795 B.n42 B.n41 163.367
R796 B.n43 B.n42 163.367
R797 B.n837 B.n43 163.367
R798 B.n837 B.n48 163.367
R799 B.n49 B.n48 163.367
R800 B.n50 B.n49 163.367
R801 B.n842 B.n50 163.367
R802 B.n842 B.n55 163.367
R803 B.n56 B.n55 163.367
R804 B.n57 B.n56 163.367
R805 B.n847 B.n57 163.367
R806 B.n847 B.n62 163.367
R807 B.n63 B.n62 163.367
R808 B.n64 B.n63 163.367
R809 B.n852 B.n64 163.367
R810 B.n852 B.n69 163.367
R811 B.n70 B.n69 163.367
R812 B.n71 B.n70 163.367
R813 B.n857 B.n71 163.367
R814 B.n857 B.n76 163.367
R815 B.n77 B.n76 163.367
R816 B.n78 B.n77 163.367
R817 B.n862 B.n78 163.367
R818 B.n862 B.n83 163.367
R819 B.n84 B.n83 163.367
R820 B.n85 B.n84 163.367
R821 B.n137 B.n85 163.367
R822 B.n662 B.n422 163.367
R823 B.n662 B.n470 163.367
R824 B.n658 B.n657 163.367
R825 B.n654 B.n653 163.367
R826 B.n650 B.n649 163.367
R827 B.n646 B.n645 163.367
R828 B.n642 B.n641 163.367
R829 B.n638 B.n637 163.367
R830 B.n634 B.n633 163.367
R831 B.n630 B.n629 163.367
R832 B.n626 B.n625 163.367
R833 B.n622 B.n621 163.367
R834 B.n618 B.n617 163.367
R835 B.n614 B.n613 163.367
R836 B.n610 B.n609 163.367
R837 B.n606 B.n605 163.367
R838 B.n602 B.n601 163.367
R839 B.n598 B.n597 163.367
R840 B.n594 B.n593 163.367
R841 B.n590 B.n589 163.367
R842 B.n586 B.n585 163.367
R843 B.n582 B.n581 163.367
R844 B.n578 B.n577 163.367
R845 B.n574 B.n573 163.367
R846 B.n570 B.n569 163.367
R847 B.n566 B.n565 163.367
R848 B.n562 B.n561 163.367
R849 B.n558 B.n557 163.367
R850 B.n554 B.n553 163.367
R851 B.n550 B.n549 163.367
R852 B.n546 B.n545 163.367
R853 B.n542 B.n541 163.367
R854 B.n538 B.n537 163.367
R855 B.n534 B.n533 163.367
R856 B.n530 B.n529 163.367
R857 B.n526 B.n525 163.367
R858 B.n522 B.n521 163.367
R859 B.n518 B.n517 163.367
R860 B.n514 B.n513 163.367
R861 B.n510 B.n509 163.367
R862 B.n506 B.n505 163.367
R863 B.n502 B.n501 163.367
R864 B.n498 B.n497 163.367
R865 B.n494 B.n493 163.367
R866 B.n490 B.n489 163.367
R867 B.n486 B.n485 163.367
R868 B.n482 B.n481 163.367
R869 B.n478 B.n469 163.367
R870 B.n669 B.n420 163.367
R871 B.n669 B.n414 163.367
R872 B.n677 B.n414 163.367
R873 B.n677 B.n412 163.367
R874 B.n681 B.n412 163.367
R875 B.n681 B.n406 163.367
R876 B.n689 B.n406 163.367
R877 B.n689 B.n404 163.367
R878 B.n693 B.n404 163.367
R879 B.n693 B.n398 163.367
R880 B.n701 B.n398 163.367
R881 B.n701 B.n396 163.367
R882 B.n705 B.n396 163.367
R883 B.n705 B.n390 163.367
R884 B.n713 B.n390 163.367
R885 B.n713 B.n388 163.367
R886 B.n717 B.n388 163.367
R887 B.n717 B.n382 163.367
R888 B.n725 B.n382 163.367
R889 B.n725 B.n380 163.367
R890 B.n729 B.n380 163.367
R891 B.n729 B.n374 163.367
R892 B.n737 B.n374 163.367
R893 B.n737 B.n372 163.367
R894 B.n741 B.n372 163.367
R895 B.n741 B.n366 163.367
R896 B.n749 B.n366 163.367
R897 B.n749 B.n364 163.367
R898 B.n753 B.n364 163.367
R899 B.n753 B.n358 163.367
R900 B.n761 B.n358 163.367
R901 B.n761 B.n356 163.367
R902 B.n765 B.n356 163.367
R903 B.n765 B.n350 163.367
R904 B.n773 B.n350 163.367
R905 B.n773 B.n348 163.367
R906 B.n777 B.n348 163.367
R907 B.n777 B.n342 163.367
R908 B.n785 B.n342 163.367
R909 B.n785 B.n340 163.367
R910 B.n789 B.n340 163.367
R911 B.n789 B.n334 163.367
R912 B.n798 B.n334 163.367
R913 B.n798 B.n332 163.367
R914 B.n802 B.n332 163.367
R915 B.n802 B.n3 163.367
R916 B.n970 B.n3 163.367
R917 B.n966 B.n2 163.367
R918 B.n966 B.n965 163.367
R919 B.n965 B.n9 163.367
R920 B.n961 B.n9 163.367
R921 B.n961 B.n11 163.367
R922 B.n957 B.n11 163.367
R923 B.n957 B.n17 163.367
R924 B.n953 B.n17 163.367
R925 B.n953 B.n19 163.367
R926 B.n949 B.n19 163.367
R927 B.n949 B.n24 163.367
R928 B.n945 B.n24 163.367
R929 B.n945 B.n26 163.367
R930 B.n941 B.n26 163.367
R931 B.n941 B.n31 163.367
R932 B.n937 B.n31 163.367
R933 B.n937 B.n33 163.367
R934 B.n933 B.n33 163.367
R935 B.n933 B.n38 163.367
R936 B.n929 B.n38 163.367
R937 B.n929 B.n40 163.367
R938 B.n925 B.n40 163.367
R939 B.n925 B.n45 163.367
R940 B.n921 B.n45 163.367
R941 B.n921 B.n47 163.367
R942 B.n917 B.n47 163.367
R943 B.n917 B.n52 163.367
R944 B.n913 B.n52 163.367
R945 B.n913 B.n54 163.367
R946 B.n909 B.n54 163.367
R947 B.n909 B.n59 163.367
R948 B.n905 B.n59 163.367
R949 B.n905 B.n61 163.367
R950 B.n901 B.n61 163.367
R951 B.n901 B.n66 163.367
R952 B.n897 B.n66 163.367
R953 B.n897 B.n68 163.367
R954 B.n893 B.n68 163.367
R955 B.n893 B.n73 163.367
R956 B.n889 B.n73 163.367
R957 B.n889 B.n75 163.367
R958 B.n885 B.n75 163.367
R959 B.n885 B.n80 163.367
R960 B.n881 B.n80 163.367
R961 B.n881 B.n82 163.367
R962 B.n877 B.n82 163.367
R963 B.n877 B.n87 163.367
R964 B.n138 B.t17 125.897
R965 B.n474 B.t11 125.897
R966 B.n140 B.t14 125.882
R967 B.n471 B.t21 125.882
R968 B.n139 B.t18 74.1156
R969 B.n475 B.t10 74.1156
R970 B.n141 B.t15 74.0998
R971 B.n472 B.t20 74.0998
R972 B.n873 B.n872 71.676
R973 B.n142 B.n90 71.676
R974 B.n146 B.n91 71.676
R975 B.n150 B.n92 71.676
R976 B.n154 B.n93 71.676
R977 B.n158 B.n94 71.676
R978 B.n162 B.n95 71.676
R979 B.n166 B.n96 71.676
R980 B.n170 B.n97 71.676
R981 B.n174 B.n98 71.676
R982 B.n178 B.n99 71.676
R983 B.n182 B.n100 71.676
R984 B.n186 B.n101 71.676
R985 B.n190 B.n102 71.676
R986 B.n194 B.n103 71.676
R987 B.n198 B.n104 71.676
R988 B.n202 B.n105 71.676
R989 B.n206 B.n106 71.676
R990 B.n210 B.n107 71.676
R991 B.n214 B.n108 71.676
R992 B.n218 B.n109 71.676
R993 B.n222 B.n110 71.676
R994 B.n227 B.n111 71.676
R995 B.n231 B.n112 71.676
R996 B.n235 B.n113 71.676
R997 B.n239 B.n114 71.676
R998 B.n243 B.n115 71.676
R999 B.n248 B.n116 71.676
R1000 B.n252 B.n117 71.676
R1001 B.n256 B.n118 71.676
R1002 B.n260 B.n119 71.676
R1003 B.n264 B.n120 71.676
R1004 B.n268 B.n121 71.676
R1005 B.n272 B.n122 71.676
R1006 B.n276 B.n123 71.676
R1007 B.n280 B.n124 71.676
R1008 B.n284 B.n125 71.676
R1009 B.n288 B.n126 71.676
R1010 B.n292 B.n127 71.676
R1011 B.n296 B.n128 71.676
R1012 B.n300 B.n129 71.676
R1013 B.n304 B.n130 71.676
R1014 B.n308 B.n131 71.676
R1015 B.n312 B.n132 71.676
R1016 B.n316 B.n133 71.676
R1017 B.n320 B.n134 71.676
R1018 B.n324 B.n135 71.676
R1019 B.n870 B.n136 71.676
R1020 B.n870 B.n869 71.676
R1021 B.n326 B.n135 71.676
R1022 B.n323 B.n134 71.676
R1023 B.n319 B.n133 71.676
R1024 B.n315 B.n132 71.676
R1025 B.n311 B.n131 71.676
R1026 B.n307 B.n130 71.676
R1027 B.n303 B.n129 71.676
R1028 B.n299 B.n128 71.676
R1029 B.n295 B.n127 71.676
R1030 B.n291 B.n126 71.676
R1031 B.n287 B.n125 71.676
R1032 B.n283 B.n124 71.676
R1033 B.n279 B.n123 71.676
R1034 B.n275 B.n122 71.676
R1035 B.n271 B.n121 71.676
R1036 B.n267 B.n120 71.676
R1037 B.n263 B.n119 71.676
R1038 B.n259 B.n118 71.676
R1039 B.n255 B.n117 71.676
R1040 B.n251 B.n116 71.676
R1041 B.n247 B.n115 71.676
R1042 B.n242 B.n114 71.676
R1043 B.n238 B.n113 71.676
R1044 B.n234 B.n112 71.676
R1045 B.n230 B.n111 71.676
R1046 B.n226 B.n110 71.676
R1047 B.n221 B.n109 71.676
R1048 B.n217 B.n108 71.676
R1049 B.n213 B.n107 71.676
R1050 B.n209 B.n106 71.676
R1051 B.n205 B.n105 71.676
R1052 B.n201 B.n104 71.676
R1053 B.n197 B.n103 71.676
R1054 B.n193 B.n102 71.676
R1055 B.n189 B.n101 71.676
R1056 B.n185 B.n100 71.676
R1057 B.n181 B.n99 71.676
R1058 B.n177 B.n98 71.676
R1059 B.n173 B.n97 71.676
R1060 B.n169 B.n96 71.676
R1061 B.n165 B.n95 71.676
R1062 B.n161 B.n94 71.676
R1063 B.n157 B.n93 71.676
R1064 B.n153 B.n92 71.676
R1065 B.n149 B.n91 71.676
R1066 B.n145 B.n90 71.676
R1067 B.n872 B.n89 71.676
R1068 B.n665 B.n664 71.676
R1069 B.n470 B.n423 71.676
R1070 B.n657 B.n424 71.676
R1071 B.n653 B.n425 71.676
R1072 B.n649 B.n426 71.676
R1073 B.n645 B.n427 71.676
R1074 B.n641 B.n428 71.676
R1075 B.n637 B.n429 71.676
R1076 B.n633 B.n430 71.676
R1077 B.n629 B.n431 71.676
R1078 B.n625 B.n432 71.676
R1079 B.n621 B.n433 71.676
R1080 B.n617 B.n434 71.676
R1081 B.n613 B.n435 71.676
R1082 B.n609 B.n436 71.676
R1083 B.n605 B.n437 71.676
R1084 B.n601 B.n438 71.676
R1085 B.n597 B.n439 71.676
R1086 B.n593 B.n440 71.676
R1087 B.n589 B.n441 71.676
R1088 B.n585 B.n442 71.676
R1089 B.n581 B.n443 71.676
R1090 B.n577 B.n444 71.676
R1091 B.n573 B.n445 71.676
R1092 B.n569 B.n446 71.676
R1093 B.n565 B.n447 71.676
R1094 B.n561 B.n448 71.676
R1095 B.n557 B.n449 71.676
R1096 B.n553 B.n450 71.676
R1097 B.n549 B.n451 71.676
R1098 B.n545 B.n452 71.676
R1099 B.n541 B.n453 71.676
R1100 B.n537 B.n454 71.676
R1101 B.n533 B.n455 71.676
R1102 B.n529 B.n456 71.676
R1103 B.n525 B.n457 71.676
R1104 B.n521 B.n458 71.676
R1105 B.n517 B.n459 71.676
R1106 B.n513 B.n460 71.676
R1107 B.n509 B.n461 71.676
R1108 B.n505 B.n462 71.676
R1109 B.n501 B.n463 71.676
R1110 B.n497 B.n464 71.676
R1111 B.n493 B.n465 71.676
R1112 B.n489 B.n466 71.676
R1113 B.n485 B.n467 71.676
R1114 B.n481 B.n468 71.676
R1115 B.n664 B.n422 71.676
R1116 B.n658 B.n423 71.676
R1117 B.n654 B.n424 71.676
R1118 B.n650 B.n425 71.676
R1119 B.n646 B.n426 71.676
R1120 B.n642 B.n427 71.676
R1121 B.n638 B.n428 71.676
R1122 B.n634 B.n429 71.676
R1123 B.n630 B.n430 71.676
R1124 B.n626 B.n431 71.676
R1125 B.n622 B.n432 71.676
R1126 B.n618 B.n433 71.676
R1127 B.n614 B.n434 71.676
R1128 B.n610 B.n435 71.676
R1129 B.n606 B.n436 71.676
R1130 B.n602 B.n437 71.676
R1131 B.n598 B.n438 71.676
R1132 B.n594 B.n439 71.676
R1133 B.n590 B.n440 71.676
R1134 B.n586 B.n441 71.676
R1135 B.n582 B.n442 71.676
R1136 B.n578 B.n443 71.676
R1137 B.n574 B.n444 71.676
R1138 B.n570 B.n445 71.676
R1139 B.n566 B.n446 71.676
R1140 B.n562 B.n447 71.676
R1141 B.n558 B.n448 71.676
R1142 B.n554 B.n449 71.676
R1143 B.n550 B.n450 71.676
R1144 B.n546 B.n451 71.676
R1145 B.n542 B.n452 71.676
R1146 B.n538 B.n453 71.676
R1147 B.n534 B.n454 71.676
R1148 B.n530 B.n455 71.676
R1149 B.n526 B.n456 71.676
R1150 B.n522 B.n457 71.676
R1151 B.n518 B.n458 71.676
R1152 B.n514 B.n459 71.676
R1153 B.n510 B.n460 71.676
R1154 B.n506 B.n461 71.676
R1155 B.n502 B.n462 71.676
R1156 B.n498 B.n463 71.676
R1157 B.n494 B.n464 71.676
R1158 B.n490 B.n465 71.676
R1159 B.n486 B.n466 71.676
R1160 B.n482 B.n467 71.676
R1161 B.n478 B.n468 71.676
R1162 B.n971 B.n970 71.676
R1163 B.n971 B.n2 71.676
R1164 B.n663 B.n419 70.8887
R1165 B.n871 B.n86 70.8887
R1166 B.n224 B.n141 59.5399
R1167 B.n245 B.n139 59.5399
R1168 B.n476 B.n475 59.5399
R1169 B.n473 B.n472 59.5399
R1170 B.n141 B.n140 51.7823
R1171 B.n139 B.n138 51.7823
R1172 B.n475 B.n474 51.7823
R1173 B.n472 B.n471 51.7823
R1174 B.n670 B.n419 41.917
R1175 B.n670 B.n415 41.917
R1176 B.n676 B.n415 41.917
R1177 B.n676 B.n411 41.917
R1178 B.n682 B.n411 41.917
R1179 B.n682 B.n407 41.917
R1180 B.n688 B.n407 41.917
R1181 B.n694 B.n403 41.917
R1182 B.n694 B.n399 41.917
R1183 B.n700 B.n399 41.917
R1184 B.n700 B.n395 41.917
R1185 B.n706 B.n395 41.917
R1186 B.n706 B.n391 41.917
R1187 B.n712 B.n391 41.917
R1188 B.n712 B.n386 41.917
R1189 B.n718 B.n386 41.917
R1190 B.n718 B.n387 41.917
R1191 B.n724 B.n379 41.917
R1192 B.n730 B.n379 41.917
R1193 B.n730 B.n375 41.917
R1194 B.n736 B.n375 41.917
R1195 B.n736 B.n370 41.917
R1196 B.n742 B.n370 41.917
R1197 B.n742 B.n371 41.917
R1198 B.n748 B.n363 41.917
R1199 B.n754 B.n363 41.917
R1200 B.n754 B.n359 41.917
R1201 B.n760 B.n359 41.917
R1202 B.n760 B.n354 41.917
R1203 B.n766 B.n354 41.917
R1204 B.n766 B.n355 41.917
R1205 B.n772 B.n347 41.917
R1206 B.n778 B.n347 41.917
R1207 B.n778 B.n343 41.917
R1208 B.n784 B.n343 41.917
R1209 B.n784 B.n339 41.917
R1210 B.n790 B.n339 41.917
R1211 B.n797 B.n335 41.917
R1212 B.n797 B.n331 41.917
R1213 B.n803 B.n331 41.917
R1214 B.n803 B.n4 41.917
R1215 B.n969 B.n4 41.917
R1216 B.n969 B.n968 41.917
R1217 B.n968 B.n967 41.917
R1218 B.n967 B.n8 41.917
R1219 B.n12 B.n8 41.917
R1220 B.n960 B.n12 41.917
R1221 B.n960 B.n959 41.917
R1222 B.n958 B.n16 41.917
R1223 B.n952 B.n16 41.917
R1224 B.n952 B.n951 41.917
R1225 B.n951 B.n950 41.917
R1226 B.n950 B.n23 41.917
R1227 B.n944 B.n23 41.917
R1228 B.n943 B.n942 41.917
R1229 B.n942 B.n30 41.917
R1230 B.n936 B.n30 41.917
R1231 B.n936 B.n935 41.917
R1232 B.n935 B.n934 41.917
R1233 B.n934 B.n37 41.917
R1234 B.n928 B.n37 41.917
R1235 B.n927 B.n926 41.917
R1236 B.n926 B.n44 41.917
R1237 B.n920 B.n44 41.917
R1238 B.n920 B.n919 41.917
R1239 B.n919 B.n918 41.917
R1240 B.n918 B.n51 41.917
R1241 B.n912 B.n51 41.917
R1242 B.n911 B.n910 41.917
R1243 B.n910 B.n58 41.917
R1244 B.n904 B.n58 41.917
R1245 B.n904 B.n903 41.917
R1246 B.n903 B.n902 41.917
R1247 B.n902 B.n65 41.917
R1248 B.n896 B.n65 41.917
R1249 B.n896 B.n895 41.917
R1250 B.n895 B.n894 41.917
R1251 B.n894 B.n72 41.917
R1252 B.n888 B.n887 41.917
R1253 B.n887 B.n886 41.917
R1254 B.n886 B.n79 41.917
R1255 B.n880 B.n79 41.917
R1256 B.n880 B.n879 41.917
R1257 B.n879 B.n878 41.917
R1258 B.n878 B.n86 41.917
R1259 B.n790 B.t6 40.6842
R1260 B.t3 B.n958 40.6842
R1261 B.n772 B.t1 36.9856
R1262 B.n944 B.t7 36.9856
R1263 B.n667 B.n666 32.0005
R1264 B.n477 B.n417 32.0005
R1265 B.n868 B.n867 32.0005
R1266 B.n875 B.n874 32.0005
R1267 B.n748 B.t5 30.8215
R1268 B.n928 B.t0 30.8215
R1269 B.t9 B.n403 27.1229
R1270 B.t13 B.n72 27.1229
R1271 B.n724 B.t2 24.6573
R1272 B.n912 B.t4 24.6573
R1273 B B.n972 18.0485
R1274 B.n387 B.t2 17.2602
R1275 B.t4 B.n911 17.2602
R1276 B.n688 B.t9 14.7946
R1277 B.n888 B.t13 14.7946
R1278 B.n371 B.t5 11.096
R1279 B.t0 B.n927 11.096
R1280 B.n668 B.n667 10.6151
R1281 B.n668 B.n413 10.6151
R1282 B.n678 B.n413 10.6151
R1283 B.n679 B.n678 10.6151
R1284 B.n680 B.n679 10.6151
R1285 B.n680 B.n405 10.6151
R1286 B.n690 B.n405 10.6151
R1287 B.n691 B.n690 10.6151
R1288 B.n692 B.n691 10.6151
R1289 B.n692 B.n397 10.6151
R1290 B.n702 B.n397 10.6151
R1291 B.n703 B.n702 10.6151
R1292 B.n704 B.n703 10.6151
R1293 B.n704 B.n389 10.6151
R1294 B.n714 B.n389 10.6151
R1295 B.n715 B.n714 10.6151
R1296 B.n716 B.n715 10.6151
R1297 B.n716 B.n381 10.6151
R1298 B.n726 B.n381 10.6151
R1299 B.n727 B.n726 10.6151
R1300 B.n728 B.n727 10.6151
R1301 B.n728 B.n373 10.6151
R1302 B.n738 B.n373 10.6151
R1303 B.n739 B.n738 10.6151
R1304 B.n740 B.n739 10.6151
R1305 B.n740 B.n365 10.6151
R1306 B.n750 B.n365 10.6151
R1307 B.n751 B.n750 10.6151
R1308 B.n752 B.n751 10.6151
R1309 B.n752 B.n357 10.6151
R1310 B.n762 B.n357 10.6151
R1311 B.n763 B.n762 10.6151
R1312 B.n764 B.n763 10.6151
R1313 B.n764 B.n349 10.6151
R1314 B.n774 B.n349 10.6151
R1315 B.n775 B.n774 10.6151
R1316 B.n776 B.n775 10.6151
R1317 B.n776 B.n341 10.6151
R1318 B.n786 B.n341 10.6151
R1319 B.n787 B.n786 10.6151
R1320 B.n788 B.n787 10.6151
R1321 B.n788 B.n333 10.6151
R1322 B.n799 B.n333 10.6151
R1323 B.n800 B.n799 10.6151
R1324 B.n801 B.n800 10.6151
R1325 B.n801 B.n0 10.6151
R1326 B.n666 B.n421 10.6151
R1327 B.n661 B.n421 10.6151
R1328 B.n661 B.n660 10.6151
R1329 B.n660 B.n659 10.6151
R1330 B.n659 B.n656 10.6151
R1331 B.n656 B.n655 10.6151
R1332 B.n655 B.n652 10.6151
R1333 B.n652 B.n651 10.6151
R1334 B.n651 B.n648 10.6151
R1335 B.n648 B.n647 10.6151
R1336 B.n647 B.n644 10.6151
R1337 B.n644 B.n643 10.6151
R1338 B.n643 B.n640 10.6151
R1339 B.n640 B.n639 10.6151
R1340 B.n639 B.n636 10.6151
R1341 B.n636 B.n635 10.6151
R1342 B.n635 B.n632 10.6151
R1343 B.n632 B.n631 10.6151
R1344 B.n631 B.n628 10.6151
R1345 B.n628 B.n627 10.6151
R1346 B.n627 B.n624 10.6151
R1347 B.n624 B.n623 10.6151
R1348 B.n623 B.n620 10.6151
R1349 B.n620 B.n619 10.6151
R1350 B.n619 B.n616 10.6151
R1351 B.n616 B.n615 10.6151
R1352 B.n615 B.n612 10.6151
R1353 B.n612 B.n611 10.6151
R1354 B.n611 B.n608 10.6151
R1355 B.n608 B.n607 10.6151
R1356 B.n607 B.n604 10.6151
R1357 B.n604 B.n603 10.6151
R1358 B.n603 B.n600 10.6151
R1359 B.n600 B.n599 10.6151
R1360 B.n599 B.n596 10.6151
R1361 B.n596 B.n595 10.6151
R1362 B.n595 B.n592 10.6151
R1363 B.n592 B.n591 10.6151
R1364 B.n591 B.n588 10.6151
R1365 B.n588 B.n587 10.6151
R1366 B.n587 B.n584 10.6151
R1367 B.n584 B.n583 10.6151
R1368 B.n580 B.n579 10.6151
R1369 B.n579 B.n576 10.6151
R1370 B.n576 B.n575 10.6151
R1371 B.n575 B.n572 10.6151
R1372 B.n572 B.n571 10.6151
R1373 B.n571 B.n568 10.6151
R1374 B.n568 B.n567 10.6151
R1375 B.n567 B.n564 10.6151
R1376 B.n564 B.n563 10.6151
R1377 B.n560 B.n559 10.6151
R1378 B.n559 B.n556 10.6151
R1379 B.n556 B.n555 10.6151
R1380 B.n555 B.n552 10.6151
R1381 B.n552 B.n551 10.6151
R1382 B.n551 B.n548 10.6151
R1383 B.n548 B.n547 10.6151
R1384 B.n547 B.n544 10.6151
R1385 B.n544 B.n543 10.6151
R1386 B.n543 B.n540 10.6151
R1387 B.n540 B.n539 10.6151
R1388 B.n539 B.n536 10.6151
R1389 B.n536 B.n535 10.6151
R1390 B.n535 B.n532 10.6151
R1391 B.n532 B.n531 10.6151
R1392 B.n531 B.n528 10.6151
R1393 B.n528 B.n527 10.6151
R1394 B.n527 B.n524 10.6151
R1395 B.n524 B.n523 10.6151
R1396 B.n523 B.n520 10.6151
R1397 B.n520 B.n519 10.6151
R1398 B.n519 B.n516 10.6151
R1399 B.n516 B.n515 10.6151
R1400 B.n515 B.n512 10.6151
R1401 B.n512 B.n511 10.6151
R1402 B.n511 B.n508 10.6151
R1403 B.n508 B.n507 10.6151
R1404 B.n507 B.n504 10.6151
R1405 B.n504 B.n503 10.6151
R1406 B.n503 B.n500 10.6151
R1407 B.n500 B.n499 10.6151
R1408 B.n499 B.n496 10.6151
R1409 B.n496 B.n495 10.6151
R1410 B.n495 B.n492 10.6151
R1411 B.n492 B.n491 10.6151
R1412 B.n491 B.n488 10.6151
R1413 B.n488 B.n487 10.6151
R1414 B.n487 B.n484 10.6151
R1415 B.n484 B.n483 10.6151
R1416 B.n483 B.n480 10.6151
R1417 B.n480 B.n479 10.6151
R1418 B.n479 B.n477 10.6151
R1419 B.n672 B.n417 10.6151
R1420 B.n673 B.n672 10.6151
R1421 B.n674 B.n673 10.6151
R1422 B.n674 B.n409 10.6151
R1423 B.n684 B.n409 10.6151
R1424 B.n685 B.n684 10.6151
R1425 B.n686 B.n685 10.6151
R1426 B.n686 B.n401 10.6151
R1427 B.n696 B.n401 10.6151
R1428 B.n697 B.n696 10.6151
R1429 B.n698 B.n697 10.6151
R1430 B.n698 B.n393 10.6151
R1431 B.n708 B.n393 10.6151
R1432 B.n709 B.n708 10.6151
R1433 B.n710 B.n709 10.6151
R1434 B.n710 B.n384 10.6151
R1435 B.n720 B.n384 10.6151
R1436 B.n721 B.n720 10.6151
R1437 B.n722 B.n721 10.6151
R1438 B.n722 B.n377 10.6151
R1439 B.n732 B.n377 10.6151
R1440 B.n733 B.n732 10.6151
R1441 B.n734 B.n733 10.6151
R1442 B.n734 B.n368 10.6151
R1443 B.n744 B.n368 10.6151
R1444 B.n745 B.n744 10.6151
R1445 B.n746 B.n745 10.6151
R1446 B.n746 B.n361 10.6151
R1447 B.n756 B.n361 10.6151
R1448 B.n757 B.n756 10.6151
R1449 B.n758 B.n757 10.6151
R1450 B.n758 B.n352 10.6151
R1451 B.n768 B.n352 10.6151
R1452 B.n769 B.n768 10.6151
R1453 B.n770 B.n769 10.6151
R1454 B.n770 B.n345 10.6151
R1455 B.n780 B.n345 10.6151
R1456 B.n781 B.n780 10.6151
R1457 B.n782 B.n781 10.6151
R1458 B.n782 B.n337 10.6151
R1459 B.n792 B.n337 10.6151
R1460 B.n793 B.n792 10.6151
R1461 B.n795 B.n793 10.6151
R1462 B.n795 B.n794 10.6151
R1463 B.n794 B.n329 10.6151
R1464 B.n806 B.n329 10.6151
R1465 B.n807 B.n806 10.6151
R1466 B.n808 B.n807 10.6151
R1467 B.n809 B.n808 10.6151
R1468 B.n810 B.n809 10.6151
R1469 B.n813 B.n810 10.6151
R1470 B.n814 B.n813 10.6151
R1471 B.n815 B.n814 10.6151
R1472 B.n816 B.n815 10.6151
R1473 B.n818 B.n816 10.6151
R1474 B.n819 B.n818 10.6151
R1475 B.n820 B.n819 10.6151
R1476 B.n821 B.n820 10.6151
R1477 B.n823 B.n821 10.6151
R1478 B.n824 B.n823 10.6151
R1479 B.n825 B.n824 10.6151
R1480 B.n826 B.n825 10.6151
R1481 B.n828 B.n826 10.6151
R1482 B.n829 B.n828 10.6151
R1483 B.n830 B.n829 10.6151
R1484 B.n831 B.n830 10.6151
R1485 B.n833 B.n831 10.6151
R1486 B.n834 B.n833 10.6151
R1487 B.n835 B.n834 10.6151
R1488 B.n836 B.n835 10.6151
R1489 B.n838 B.n836 10.6151
R1490 B.n839 B.n838 10.6151
R1491 B.n840 B.n839 10.6151
R1492 B.n841 B.n840 10.6151
R1493 B.n843 B.n841 10.6151
R1494 B.n844 B.n843 10.6151
R1495 B.n845 B.n844 10.6151
R1496 B.n846 B.n845 10.6151
R1497 B.n848 B.n846 10.6151
R1498 B.n849 B.n848 10.6151
R1499 B.n850 B.n849 10.6151
R1500 B.n851 B.n850 10.6151
R1501 B.n853 B.n851 10.6151
R1502 B.n854 B.n853 10.6151
R1503 B.n855 B.n854 10.6151
R1504 B.n856 B.n855 10.6151
R1505 B.n858 B.n856 10.6151
R1506 B.n859 B.n858 10.6151
R1507 B.n860 B.n859 10.6151
R1508 B.n861 B.n860 10.6151
R1509 B.n863 B.n861 10.6151
R1510 B.n864 B.n863 10.6151
R1511 B.n865 B.n864 10.6151
R1512 B.n866 B.n865 10.6151
R1513 B.n867 B.n866 10.6151
R1514 B.n964 B.n1 10.6151
R1515 B.n964 B.n963 10.6151
R1516 B.n963 B.n962 10.6151
R1517 B.n962 B.n10 10.6151
R1518 B.n956 B.n10 10.6151
R1519 B.n956 B.n955 10.6151
R1520 B.n955 B.n954 10.6151
R1521 B.n954 B.n18 10.6151
R1522 B.n948 B.n18 10.6151
R1523 B.n948 B.n947 10.6151
R1524 B.n947 B.n946 10.6151
R1525 B.n946 B.n25 10.6151
R1526 B.n940 B.n25 10.6151
R1527 B.n940 B.n939 10.6151
R1528 B.n939 B.n938 10.6151
R1529 B.n938 B.n32 10.6151
R1530 B.n932 B.n32 10.6151
R1531 B.n932 B.n931 10.6151
R1532 B.n931 B.n930 10.6151
R1533 B.n930 B.n39 10.6151
R1534 B.n924 B.n39 10.6151
R1535 B.n924 B.n923 10.6151
R1536 B.n923 B.n922 10.6151
R1537 B.n922 B.n46 10.6151
R1538 B.n916 B.n46 10.6151
R1539 B.n916 B.n915 10.6151
R1540 B.n915 B.n914 10.6151
R1541 B.n914 B.n53 10.6151
R1542 B.n908 B.n53 10.6151
R1543 B.n908 B.n907 10.6151
R1544 B.n907 B.n906 10.6151
R1545 B.n906 B.n60 10.6151
R1546 B.n900 B.n60 10.6151
R1547 B.n900 B.n899 10.6151
R1548 B.n899 B.n898 10.6151
R1549 B.n898 B.n67 10.6151
R1550 B.n892 B.n67 10.6151
R1551 B.n892 B.n891 10.6151
R1552 B.n891 B.n890 10.6151
R1553 B.n890 B.n74 10.6151
R1554 B.n884 B.n74 10.6151
R1555 B.n884 B.n883 10.6151
R1556 B.n883 B.n882 10.6151
R1557 B.n882 B.n81 10.6151
R1558 B.n876 B.n81 10.6151
R1559 B.n876 B.n875 10.6151
R1560 B.n874 B.n88 10.6151
R1561 B.n143 B.n88 10.6151
R1562 B.n144 B.n143 10.6151
R1563 B.n147 B.n144 10.6151
R1564 B.n148 B.n147 10.6151
R1565 B.n151 B.n148 10.6151
R1566 B.n152 B.n151 10.6151
R1567 B.n155 B.n152 10.6151
R1568 B.n156 B.n155 10.6151
R1569 B.n159 B.n156 10.6151
R1570 B.n160 B.n159 10.6151
R1571 B.n163 B.n160 10.6151
R1572 B.n164 B.n163 10.6151
R1573 B.n167 B.n164 10.6151
R1574 B.n168 B.n167 10.6151
R1575 B.n171 B.n168 10.6151
R1576 B.n172 B.n171 10.6151
R1577 B.n175 B.n172 10.6151
R1578 B.n176 B.n175 10.6151
R1579 B.n179 B.n176 10.6151
R1580 B.n180 B.n179 10.6151
R1581 B.n183 B.n180 10.6151
R1582 B.n184 B.n183 10.6151
R1583 B.n187 B.n184 10.6151
R1584 B.n188 B.n187 10.6151
R1585 B.n191 B.n188 10.6151
R1586 B.n192 B.n191 10.6151
R1587 B.n195 B.n192 10.6151
R1588 B.n196 B.n195 10.6151
R1589 B.n199 B.n196 10.6151
R1590 B.n200 B.n199 10.6151
R1591 B.n203 B.n200 10.6151
R1592 B.n204 B.n203 10.6151
R1593 B.n207 B.n204 10.6151
R1594 B.n208 B.n207 10.6151
R1595 B.n211 B.n208 10.6151
R1596 B.n212 B.n211 10.6151
R1597 B.n215 B.n212 10.6151
R1598 B.n216 B.n215 10.6151
R1599 B.n219 B.n216 10.6151
R1600 B.n220 B.n219 10.6151
R1601 B.n223 B.n220 10.6151
R1602 B.n228 B.n225 10.6151
R1603 B.n229 B.n228 10.6151
R1604 B.n232 B.n229 10.6151
R1605 B.n233 B.n232 10.6151
R1606 B.n236 B.n233 10.6151
R1607 B.n237 B.n236 10.6151
R1608 B.n240 B.n237 10.6151
R1609 B.n241 B.n240 10.6151
R1610 B.n244 B.n241 10.6151
R1611 B.n249 B.n246 10.6151
R1612 B.n250 B.n249 10.6151
R1613 B.n253 B.n250 10.6151
R1614 B.n254 B.n253 10.6151
R1615 B.n257 B.n254 10.6151
R1616 B.n258 B.n257 10.6151
R1617 B.n261 B.n258 10.6151
R1618 B.n262 B.n261 10.6151
R1619 B.n265 B.n262 10.6151
R1620 B.n266 B.n265 10.6151
R1621 B.n269 B.n266 10.6151
R1622 B.n270 B.n269 10.6151
R1623 B.n273 B.n270 10.6151
R1624 B.n274 B.n273 10.6151
R1625 B.n277 B.n274 10.6151
R1626 B.n278 B.n277 10.6151
R1627 B.n281 B.n278 10.6151
R1628 B.n282 B.n281 10.6151
R1629 B.n285 B.n282 10.6151
R1630 B.n286 B.n285 10.6151
R1631 B.n289 B.n286 10.6151
R1632 B.n290 B.n289 10.6151
R1633 B.n293 B.n290 10.6151
R1634 B.n294 B.n293 10.6151
R1635 B.n297 B.n294 10.6151
R1636 B.n298 B.n297 10.6151
R1637 B.n301 B.n298 10.6151
R1638 B.n302 B.n301 10.6151
R1639 B.n305 B.n302 10.6151
R1640 B.n306 B.n305 10.6151
R1641 B.n309 B.n306 10.6151
R1642 B.n310 B.n309 10.6151
R1643 B.n313 B.n310 10.6151
R1644 B.n314 B.n313 10.6151
R1645 B.n317 B.n314 10.6151
R1646 B.n318 B.n317 10.6151
R1647 B.n321 B.n318 10.6151
R1648 B.n322 B.n321 10.6151
R1649 B.n325 B.n322 10.6151
R1650 B.n327 B.n325 10.6151
R1651 B.n328 B.n327 10.6151
R1652 B.n868 B.n328 10.6151
R1653 B.n583 B.n473 9.36635
R1654 B.n560 B.n476 9.36635
R1655 B.n224 B.n223 9.36635
R1656 B.n246 B.n245 9.36635
R1657 B.n972 B.n0 8.11757
R1658 B.n972 B.n1 8.11757
R1659 B.n355 B.t1 4.93185
R1660 B.t7 B.n943 4.93185
R1661 B.n580 B.n473 1.24928
R1662 B.n563 B.n476 1.24928
R1663 B.n225 B.n224 1.24928
R1664 B.n245 B.n244 1.24928
R1665 B.t6 B.n335 1.23334
R1666 B.n959 B.t3 1.23334
R1667 VN.n51 VN.n27 161.3
R1668 VN.n50 VN.n49 161.3
R1669 VN.n48 VN.n28 161.3
R1670 VN.n47 VN.n46 161.3
R1671 VN.n45 VN.n29 161.3
R1672 VN.n43 VN.n42 161.3
R1673 VN.n41 VN.n30 161.3
R1674 VN.n40 VN.n39 161.3
R1675 VN.n38 VN.n31 161.3
R1676 VN.n37 VN.n36 161.3
R1677 VN.n35 VN.n32 161.3
R1678 VN.n24 VN.n0 161.3
R1679 VN.n23 VN.n22 161.3
R1680 VN.n21 VN.n1 161.3
R1681 VN.n20 VN.n19 161.3
R1682 VN.n18 VN.n2 161.3
R1683 VN.n16 VN.n15 161.3
R1684 VN.n14 VN.n3 161.3
R1685 VN.n13 VN.n12 161.3
R1686 VN.n11 VN.n4 161.3
R1687 VN.n10 VN.n9 161.3
R1688 VN.n8 VN.n5 161.3
R1689 VN.n7 VN.t2 161.194
R1690 VN.n34 VN.t5 161.194
R1691 VN.n6 VN.t4 129.46
R1692 VN.n17 VN.t0 129.46
R1693 VN.n25 VN.t6 129.46
R1694 VN.n33 VN.t1 129.46
R1695 VN.n44 VN.t7 129.46
R1696 VN.n52 VN.t3 129.46
R1697 VN.n26 VN.n25 98.2783
R1698 VN.n53 VN.n52 98.2783
R1699 VN.n7 VN.n6 68.0271
R1700 VN.n34 VN.n33 68.0271
R1701 VN.n12 VN.n11 56.5193
R1702 VN.n39 VN.n38 56.5193
R1703 VN VN.n53 50.3845
R1704 VN.n19 VN.n1 48.2635
R1705 VN.n46 VN.n28 48.2635
R1706 VN.n23 VN.n1 32.7233
R1707 VN.n50 VN.n28 32.7233
R1708 VN.n10 VN.n5 24.4675
R1709 VN.n11 VN.n10 24.4675
R1710 VN.n12 VN.n3 24.4675
R1711 VN.n16 VN.n3 24.4675
R1712 VN.n19 VN.n18 24.4675
R1713 VN.n24 VN.n23 24.4675
R1714 VN.n38 VN.n37 24.4675
R1715 VN.n37 VN.n32 24.4675
R1716 VN.n46 VN.n45 24.4675
R1717 VN.n43 VN.n30 24.4675
R1718 VN.n39 VN.n30 24.4675
R1719 VN.n51 VN.n50 24.4675
R1720 VN.n18 VN.n17 20.3081
R1721 VN.n45 VN.n44 20.3081
R1722 VN.n25 VN.n24 12.4787
R1723 VN.n52 VN.n51 12.4787
R1724 VN.n35 VN.n34 9.75521
R1725 VN.n8 VN.n7 9.75521
R1726 VN.n6 VN.n5 4.15989
R1727 VN.n17 VN.n16 4.15989
R1728 VN.n33 VN.n32 4.15989
R1729 VN.n44 VN.n43 4.15989
R1730 VN.n53 VN.n27 0.278367
R1731 VN.n26 VN.n0 0.278367
R1732 VN.n49 VN.n27 0.189894
R1733 VN.n49 VN.n48 0.189894
R1734 VN.n48 VN.n47 0.189894
R1735 VN.n47 VN.n29 0.189894
R1736 VN.n42 VN.n29 0.189894
R1737 VN.n42 VN.n41 0.189894
R1738 VN.n41 VN.n40 0.189894
R1739 VN.n40 VN.n31 0.189894
R1740 VN.n36 VN.n31 0.189894
R1741 VN.n36 VN.n35 0.189894
R1742 VN.n9 VN.n8 0.189894
R1743 VN.n9 VN.n4 0.189894
R1744 VN.n13 VN.n4 0.189894
R1745 VN.n14 VN.n13 0.189894
R1746 VN.n15 VN.n14 0.189894
R1747 VN.n15 VN.n2 0.189894
R1748 VN.n20 VN.n2 0.189894
R1749 VN.n21 VN.n20 0.189894
R1750 VN.n22 VN.n21 0.189894
R1751 VN.n22 VN.n0 0.189894
R1752 VN VN.n26 0.153454
R1753 VDD2.n2 VDD2.n1 64.6283
R1754 VDD2.n2 VDD2.n0 64.6283
R1755 VDD2 VDD2.n5 64.6255
R1756 VDD2.n4 VDD2.n3 63.533
R1757 VDD2.n4 VDD2.n2 44.9093
R1758 VDD2.n5 VDD2.t3 1.57568
R1759 VDD2.n5 VDD2.t6 1.57568
R1760 VDD2.n3 VDD2.t1 1.57568
R1761 VDD2.n3 VDD2.t2 1.57568
R1762 VDD2.n1 VDD2.t0 1.57568
R1763 VDD2.n1 VDD2.t5 1.57568
R1764 VDD2.n0 VDD2.t4 1.57568
R1765 VDD2.n0 VDD2.t7 1.57568
R1766 VDD2 VDD2.n4 1.20955
R1767 VTAIL.n11 VTAIL.t5 48.4293
R1768 VTAIL.n10 VTAIL.t10 48.4293
R1769 VTAIL.n7 VTAIL.t12 48.4293
R1770 VTAIL.n15 VTAIL.t9 48.4292
R1771 VTAIL.n2 VTAIL.t13 48.4292
R1772 VTAIL.n3 VTAIL.t6 48.4292
R1773 VTAIL.n6 VTAIL.t2 48.4292
R1774 VTAIL.n14 VTAIL.t3 48.4292
R1775 VTAIL.n13 VTAIL.n12 46.8542
R1776 VTAIL.n9 VTAIL.n8 46.8542
R1777 VTAIL.n1 VTAIL.n0 46.854
R1778 VTAIL.n5 VTAIL.n4 46.854
R1779 VTAIL.n15 VTAIL.n14 25.5048
R1780 VTAIL.n7 VTAIL.n6 25.5048
R1781 VTAIL.n9 VTAIL.n7 2.30222
R1782 VTAIL.n10 VTAIL.n9 2.30222
R1783 VTAIL.n13 VTAIL.n11 2.30222
R1784 VTAIL.n14 VTAIL.n13 2.30222
R1785 VTAIL.n6 VTAIL.n5 2.30222
R1786 VTAIL.n5 VTAIL.n3 2.30222
R1787 VTAIL.n2 VTAIL.n1 2.30222
R1788 VTAIL VTAIL.n15 2.24403
R1789 VTAIL.n0 VTAIL.t11 1.57568
R1790 VTAIL.n0 VTAIL.t15 1.57568
R1791 VTAIL.n4 VTAIL.t4 1.57568
R1792 VTAIL.n4 VTAIL.t1 1.57568
R1793 VTAIL.n12 VTAIL.t7 1.57568
R1794 VTAIL.n12 VTAIL.t0 1.57568
R1795 VTAIL.n8 VTAIL.t8 1.57568
R1796 VTAIL.n8 VTAIL.t14 1.57568
R1797 VTAIL.n11 VTAIL.n10 0.470328
R1798 VTAIL.n3 VTAIL.n2 0.470328
R1799 VTAIL VTAIL.n1 0.0586897
R1800 VP.n16 VP.n13 161.3
R1801 VP.n18 VP.n17 161.3
R1802 VP.n19 VP.n12 161.3
R1803 VP.n21 VP.n20 161.3
R1804 VP.n22 VP.n11 161.3
R1805 VP.n24 VP.n23 161.3
R1806 VP.n26 VP.n10 161.3
R1807 VP.n28 VP.n27 161.3
R1808 VP.n29 VP.n9 161.3
R1809 VP.n31 VP.n30 161.3
R1810 VP.n32 VP.n8 161.3
R1811 VP.n62 VP.n0 161.3
R1812 VP.n61 VP.n60 161.3
R1813 VP.n59 VP.n1 161.3
R1814 VP.n58 VP.n57 161.3
R1815 VP.n56 VP.n2 161.3
R1816 VP.n54 VP.n53 161.3
R1817 VP.n52 VP.n3 161.3
R1818 VP.n51 VP.n50 161.3
R1819 VP.n49 VP.n4 161.3
R1820 VP.n48 VP.n47 161.3
R1821 VP.n46 VP.n5 161.3
R1822 VP.n45 VP.n44 161.3
R1823 VP.n42 VP.n6 161.3
R1824 VP.n41 VP.n40 161.3
R1825 VP.n39 VP.n7 161.3
R1826 VP.n38 VP.n37 161.3
R1827 VP.n15 VP.t3 161.194
R1828 VP.n36 VP.t2 129.46
R1829 VP.n43 VP.t7 129.46
R1830 VP.n55 VP.t1 129.46
R1831 VP.n63 VP.t5 129.46
R1832 VP.n33 VP.t4 129.46
R1833 VP.n25 VP.t0 129.46
R1834 VP.n14 VP.t6 129.46
R1835 VP.n36 VP.n35 98.2783
R1836 VP.n64 VP.n63 98.2783
R1837 VP.n34 VP.n33 98.2783
R1838 VP.n15 VP.n14 68.0271
R1839 VP.n50 VP.n49 56.5193
R1840 VP.n20 VP.n19 56.5193
R1841 VP.n35 VP.n34 50.1056
R1842 VP.n42 VP.n41 48.2635
R1843 VP.n57 VP.n1 48.2635
R1844 VP.n27 VP.n9 48.2635
R1845 VP.n41 VP.n7 32.7233
R1846 VP.n61 VP.n1 32.7233
R1847 VP.n31 VP.n9 32.7233
R1848 VP.n37 VP.n7 24.4675
R1849 VP.n44 VP.n42 24.4675
R1850 VP.n48 VP.n5 24.4675
R1851 VP.n49 VP.n48 24.4675
R1852 VP.n50 VP.n3 24.4675
R1853 VP.n54 VP.n3 24.4675
R1854 VP.n57 VP.n56 24.4675
R1855 VP.n62 VP.n61 24.4675
R1856 VP.n32 VP.n31 24.4675
R1857 VP.n20 VP.n11 24.4675
R1858 VP.n24 VP.n11 24.4675
R1859 VP.n27 VP.n26 24.4675
R1860 VP.n18 VP.n13 24.4675
R1861 VP.n19 VP.n18 24.4675
R1862 VP.n44 VP.n43 20.3081
R1863 VP.n56 VP.n55 20.3081
R1864 VP.n26 VP.n25 20.3081
R1865 VP.n37 VP.n36 12.4787
R1866 VP.n63 VP.n62 12.4787
R1867 VP.n33 VP.n32 12.4787
R1868 VP.n16 VP.n15 9.75521
R1869 VP.n43 VP.n5 4.15989
R1870 VP.n55 VP.n54 4.15989
R1871 VP.n25 VP.n24 4.15989
R1872 VP.n14 VP.n13 4.15989
R1873 VP.n34 VP.n8 0.278367
R1874 VP.n38 VP.n35 0.278367
R1875 VP.n64 VP.n0 0.278367
R1876 VP.n17 VP.n16 0.189894
R1877 VP.n17 VP.n12 0.189894
R1878 VP.n21 VP.n12 0.189894
R1879 VP.n22 VP.n21 0.189894
R1880 VP.n23 VP.n22 0.189894
R1881 VP.n23 VP.n10 0.189894
R1882 VP.n28 VP.n10 0.189894
R1883 VP.n29 VP.n28 0.189894
R1884 VP.n30 VP.n29 0.189894
R1885 VP.n30 VP.n8 0.189894
R1886 VP.n39 VP.n38 0.189894
R1887 VP.n40 VP.n39 0.189894
R1888 VP.n40 VP.n6 0.189894
R1889 VP.n45 VP.n6 0.189894
R1890 VP.n46 VP.n45 0.189894
R1891 VP.n47 VP.n46 0.189894
R1892 VP.n47 VP.n4 0.189894
R1893 VP.n51 VP.n4 0.189894
R1894 VP.n52 VP.n51 0.189894
R1895 VP.n53 VP.n52 0.189894
R1896 VP.n53 VP.n2 0.189894
R1897 VP.n58 VP.n2 0.189894
R1898 VP.n59 VP.n58 0.189894
R1899 VP.n60 VP.n59 0.189894
R1900 VP.n60 VP.n0 0.189894
R1901 VP VP.n64 0.153454
R1902 VDD1 VDD1.n0 64.742
R1903 VDD1.n3 VDD1.n2 64.6283
R1904 VDD1.n3 VDD1.n1 64.6283
R1905 VDD1.n5 VDD1.n4 63.5328
R1906 VDD1.n5 VDD1.n3 45.4923
R1907 VDD1.n4 VDD1.t7 1.57568
R1908 VDD1.n4 VDD1.t3 1.57568
R1909 VDD1.n0 VDD1.t4 1.57568
R1910 VDD1.n0 VDD1.t1 1.57568
R1911 VDD1.n2 VDD1.t6 1.57568
R1912 VDD1.n2 VDD1.t2 1.57568
R1913 VDD1.n1 VDD1.t5 1.57568
R1914 VDD1.n1 VDD1.t0 1.57568
R1915 VDD1 VDD1.n5 1.09317
C0 VP VDD2 0.491783f
C1 VN VDD1 0.151036f
C2 VTAIL VDD1 8.25521f
C3 VP VDD1 9.23229f
C4 VDD2 VDD1 1.64054f
C5 VTAIL VN 9.17295f
C6 VP VN 7.45143f
C7 VDD2 VN 8.8928f
C8 VP VTAIL 9.18705f
C9 VDD2 VTAIL 8.307879f
C10 VDD2 B 5.137979f
C11 VDD1 B 5.54745f
C12 VTAIL B 10.648677f
C13 VN B 14.5704f
C14 VP B 13.111974f
C15 VDD1.t4 B 0.245254f
C16 VDD1.t1 B 0.245254f
C17 VDD1.n0 B 2.20216f
C18 VDD1.t5 B 0.245254f
C19 VDD1.t0 B 0.245254f
C20 VDD1.n1 B 2.20116f
C21 VDD1.t6 B 0.245254f
C22 VDD1.t2 B 0.245254f
C23 VDD1.n2 B 2.20116f
C24 VDD1.n3 B 3.17587f
C25 VDD1.t7 B 0.245254f
C26 VDD1.t3 B 0.245254f
C27 VDD1.n4 B 2.19294f
C28 VDD1.n5 B 2.89802f
C29 VP.n0 B 0.03157f
C30 VP.t5 B 1.92152f
C31 VP.n1 B 0.021401f
C32 VP.n2 B 0.023945f
C33 VP.t1 B 1.92152f
C34 VP.n3 B 0.044628f
C35 VP.n4 B 0.023945f
C36 VP.n5 B 0.02634f
C37 VP.n6 B 0.023945f
C38 VP.n7 B 0.048296f
C39 VP.n8 B 0.03157f
C40 VP.t4 B 1.92152f
C41 VP.n9 B 0.021401f
C42 VP.n10 B 0.023945f
C43 VP.t0 B 1.92152f
C44 VP.n11 B 0.044628f
C45 VP.n12 B 0.023945f
C46 VP.n13 B 0.02634f
C47 VP.t3 B 2.08152f
C48 VP.t6 B 1.92152f
C49 VP.n14 B 0.738055f
C50 VP.n15 B 0.73419f
C51 VP.n16 B 0.207149f
C52 VP.n17 B 0.023945f
C53 VP.n18 B 0.044628f
C54 VP.n19 B 0.034956f
C55 VP.n20 B 0.034956f
C56 VP.n21 B 0.023945f
C57 VP.n22 B 0.023945f
C58 VP.n23 B 0.023945f
C59 VP.n24 B 0.02634f
C60 VP.n25 B 0.679984f
C61 VP.n26 B 0.040882f
C62 VP.n27 B 0.044844f
C63 VP.n28 B 0.023945f
C64 VP.n29 B 0.023945f
C65 VP.n30 B 0.023945f
C66 VP.n31 B 0.048296f
C67 VP.n32 B 0.033831f
C68 VP.n33 B 0.755083f
C69 VP.n34 B 1.3327f
C70 VP.n35 B 1.34988f
C71 VP.t2 B 1.92152f
C72 VP.n36 B 0.755083f
C73 VP.n37 B 0.033831f
C74 VP.n38 B 0.03157f
C75 VP.n39 B 0.023945f
C76 VP.n40 B 0.023945f
C77 VP.n41 B 0.021401f
C78 VP.n42 B 0.044844f
C79 VP.t7 B 1.92152f
C80 VP.n43 B 0.679984f
C81 VP.n44 B 0.040882f
C82 VP.n45 B 0.023945f
C83 VP.n46 B 0.023945f
C84 VP.n47 B 0.023945f
C85 VP.n48 B 0.044628f
C86 VP.n49 B 0.034956f
C87 VP.n50 B 0.034956f
C88 VP.n51 B 0.023945f
C89 VP.n52 B 0.023945f
C90 VP.n53 B 0.023945f
C91 VP.n54 B 0.02634f
C92 VP.n55 B 0.679984f
C93 VP.n56 B 0.040882f
C94 VP.n57 B 0.044844f
C95 VP.n58 B 0.023945f
C96 VP.n59 B 0.023945f
C97 VP.n60 B 0.023945f
C98 VP.n61 B 0.048296f
C99 VP.n62 B 0.033831f
C100 VP.n63 B 0.755083f
C101 VP.n64 B 0.035604f
C102 VTAIL.t11 B 0.1939f
C103 VTAIL.t15 B 0.1939f
C104 VTAIL.n0 B 1.67782f
C105 VTAIL.n1 B 0.338747f
C106 VTAIL.t13 B 2.14117f
C107 VTAIL.n2 B 0.430108f
C108 VTAIL.t6 B 2.14117f
C109 VTAIL.n3 B 0.430108f
C110 VTAIL.t4 B 0.1939f
C111 VTAIL.t1 B 0.1939f
C112 VTAIL.n4 B 1.67782f
C113 VTAIL.n5 B 0.479863f
C114 VTAIL.t2 B 2.14117f
C115 VTAIL.n6 B 1.49208f
C116 VTAIL.t12 B 2.14118f
C117 VTAIL.n7 B 1.49207f
C118 VTAIL.t8 B 0.1939f
C119 VTAIL.t14 B 0.1939f
C120 VTAIL.n8 B 1.67782f
C121 VTAIL.n9 B 0.479858f
C122 VTAIL.t10 B 2.14118f
C123 VTAIL.n10 B 0.430095f
C124 VTAIL.t5 B 2.14118f
C125 VTAIL.n11 B 0.430095f
C126 VTAIL.t7 B 0.1939f
C127 VTAIL.t0 B 0.1939f
C128 VTAIL.n12 B 1.67782f
C129 VTAIL.n13 B 0.479858f
C130 VTAIL.t3 B 2.14117f
C131 VTAIL.n14 B 1.49208f
C132 VTAIL.t9 B 2.14117f
C133 VTAIL.n15 B 1.48842f
C134 VDD2.t4 B 0.242312f
C135 VDD2.t7 B 0.242312f
C136 VDD2.n0 B 2.17476f
C137 VDD2.t0 B 0.242312f
C138 VDD2.t5 B 0.242312f
C139 VDD2.n1 B 2.17476f
C140 VDD2.n2 B 3.08684f
C141 VDD2.t1 B 0.242312f
C142 VDD2.t2 B 0.242312f
C143 VDD2.n3 B 2.16665f
C144 VDD2.n4 B 2.83323f
C145 VDD2.t3 B 0.242312f
C146 VDD2.t6 B 0.242312f
C147 VDD2.n5 B 2.17472f
C148 VN.n0 B 0.031164f
C149 VN.t6 B 1.89679f
C150 VN.n1 B 0.021126f
C151 VN.n2 B 0.023637f
C152 VN.t0 B 1.89679f
C153 VN.n3 B 0.044054f
C154 VN.n4 B 0.023637f
C155 VN.n5 B 0.026001f
C156 VN.t2 B 2.05474f
C157 VN.t4 B 1.89679f
C158 VN.n6 B 0.72856f
C159 VN.n7 B 0.724744f
C160 VN.n8 B 0.204484f
C161 VN.n9 B 0.023637f
C162 VN.n10 B 0.044054f
C163 VN.n11 B 0.034506f
C164 VN.n12 B 0.034506f
C165 VN.n13 B 0.023637f
C166 VN.n14 B 0.023637f
C167 VN.n15 B 0.023637f
C168 VN.n16 B 0.026001f
C169 VN.n17 B 0.671235f
C170 VN.n18 B 0.040356f
C171 VN.n19 B 0.044267f
C172 VN.n20 B 0.023637f
C173 VN.n21 B 0.023637f
C174 VN.n22 B 0.023637f
C175 VN.n23 B 0.047674f
C176 VN.n24 B 0.033396f
C177 VN.n25 B 0.745368f
C178 VN.n26 B 0.035146f
C179 VN.n27 B 0.031164f
C180 VN.t3 B 1.89679f
C181 VN.n28 B 0.021126f
C182 VN.n29 B 0.023637f
C183 VN.t7 B 1.89679f
C184 VN.n30 B 0.044054f
C185 VN.n31 B 0.023637f
C186 VN.n32 B 0.026001f
C187 VN.t5 B 2.05474f
C188 VN.t1 B 1.89679f
C189 VN.n33 B 0.72856f
C190 VN.n34 B 0.724744f
C191 VN.n35 B 0.204484f
C192 VN.n36 B 0.023637f
C193 VN.n37 B 0.044054f
C194 VN.n38 B 0.034506f
C195 VN.n39 B 0.034506f
C196 VN.n40 B 0.023637f
C197 VN.n41 B 0.023637f
C198 VN.n42 B 0.023637f
C199 VN.n43 B 0.026001f
C200 VN.n44 B 0.671235f
C201 VN.n45 B 0.040356f
C202 VN.n46 B 0.044267f
C203 VN.n47 B 0.023637f
C204 VN.n48 B 0.023637f
C205 VN.n49 B 0.023637f
C206 VN.n50 B 0.047674f
C207 VN.n51 B 0.033396f
C208 VN.n52 B 0.745368f
C209 VN.n53 B 1.32826f
.ends

