* NGSPICE file created from diff_pair_sample_1788.ext - technology: sky130A

.subckt diff_pair_sample_1788 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X1 VDD1.t6 VP.t1 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=1.32
X2 VTAIL.t8 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=1.32
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=1.32
X4 VDD2.t7 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X5 VDD2.t6 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=1.32
X6 VTAIL.t7 VN.t2 VDD2.t5 B.t21 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X7 VDD2.t4 VN.t3 VTAIL.t6 B.t20 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X8 VTAIL.t5 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=1.32
X9 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=1.32
X10 VDD1.t4 VP.t3 VTAIL.t13 B.t20 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X11 VDD1.t3 VP.t4 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=1.32
X12 VTAIL.t15 VP.t5 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X13 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=1.32
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=1.32
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=1.32
X16 VTAIL.t9 VP.t6 VDD1.t1 B.t21 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X17 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=1.32
X18 VTAIL.t4 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=1.32
X19 VTAIL.t10 VP.t7 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=1.32
R0 VP.n25 VP.n5 174.827
R1 VP.n44 VP.n43 174.827
R2 VP.n24 VP.n23 174.827
R3 VP.n12 VP.n9 161.3
R4 VP.n14 VP.n13 161.3
R5 VP.n15 VP.n8 161.3
R6 VP.n18 VP.n17 161.3
R7 VP.n19 VP.n7 161.3
R8 VP.n21 VP.n20 161.3
R9 VP.n22 VP.n6 161.3
R10 VP.n42 VP.n0 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n39 VP.n1 161.3
R13 VP.n38 VP.n37 161.3
R14 VP.n35 VP.n2 161.3
R15 VP.n34 VP.n33 161.3
R16 VP.n32 VP.n3 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n28 VP.n4 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n11 VP.t2 128.549
R21 VP.n5 VP.t7 100.418
R22 VP.n29 VP.t0 100.418
R23 VP.n36 VP.t5 100.418
R24 VP.n43 VP.t4 100.418
R25 VP.n23 VP.t1 100.418
R26 VP.n16 VP.t6 100.418
R27 VP.n10 VP.t3 100.418
R28 VP.n11 VP.n10 61.9082
R29 VP.n35 VP.n34 56.5617
R30 VP.n15 VP.n14 56.5617
R31 VP.n30 VP.n28 50.2647
R32 VP.n41 VP.n1 50.2647
R33 VP.n21 VP.n7 50.2647
R34 VP.n25 VP.n24 39.8793
R35 VP.n28 VP.n27 30.8893
R36 VP.n42 VP.n41 30.8893
R37 VP.n22 VP.n21 30.8893
R38 VP.n12 VP.n11 27.4757
R39 VP.n34 VP.n3 24.5923
R40 VP.n37 VP.n35 24.5923
R41 VP.n17 VP.n15 24.5923
R42 VP.n14 VP.n9 24.5923
R43 VP.n30 VP.n29 20.9036
R44 VP.n36 VP.n1 20.9036
R45 VP.n16 VP.n7 20.9036
R46 VP.n27 VP.n5 11.0668
R47 VP.n43 VP.n42 11.0668
R48 VP.n23 VP.n22 11.0668
R49 VP.n29 VP.n3 3.68928
R50 VP.n37 VP.n36 3.68928
R51 VP.n17 VP.n16 3.68928
R52 VP.n10 VP.n9 3.68928
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VTAIL.n11 VTAIL.t8 58.1546
R73 VTAIL.n10 VTAIL.t0 58.1546
R74 VTAIL.n7 VTAIL.t4 58.1546
R75 VTAIL.n14 VTAIL.t12 58.1537
R76 VTAIL.n15 VTAIL.t2 58.1536
R77 VTAIL.n2 VTAIL.t5 58.1536
R78 VTAIL.n3 VTAIL.t14 58.1536
R79 VTAIL.n6 VTAIL.t10 58.1536
R80 VTAIL.n13 VTAIL.n12 54.5546
R81 VTAIL.n9 VTAIL.n8 54.5546
R82 VTAIL.n1 VTAIL.n0 54.5545
R83 VTAIL.n5 VTAIL.n4 54.5545
R84 VTAIL.n15 VTAIL.n14 18.5307
R85 VTAIL.n7 VTAIL.n6 18.5307
R86 VTAIL.n0 VTAIL.t6 3.6005
R87 VTAIL.n0 VTAIL.t7 3.6005
R88 VTAIL.n4 VTAIL.t11 3.6005
R89 VTAIL.n4 VTAIL.t15 3.6005
R90 VTAIL.n12 VTAIL.t13 3.6005
R91 VTAIL.n12 VTAIL.t9 3.6005
R92 VTAIL.n8 VTAIL.t3 3.6005
R93 VTAIL.n8 VTAIL.t1 3.6005
R94 VTAIL.n9 VTAIL.n7 1.42291
R95 VTAIL.n10 VTAIL.n9 1.42291
R96 VTAIL.n13 VTAIL.n11 1.42291
R97 VTAIL.n14 VTAIL.n13 1.42291
R98 VTAIL.n6 VTAIL.n5 1.42291
R99 VTAIL.n5 VTAIL.n3 1.42291
R100 VTAIL.n2 VTAIL.n1 1.42291
R101 VTAIL VTAIL.n15 1.36472
R102 VTAIL.n11 VTAIL.n10 0.470328
R103 VTAIL.n3 VTAIL.n2 0.470328
R104 VTAIL VTAIL.n1 0.0586897
R105 VDD1 VDD1.n0 72.0028
R106 VDD1.n3 VDD1.n2 71.8892
R107 VDD1.n3 VDD1.n1 71.8892
R108 VDD1.n5 VDD1.n4 71.2325
R109 VDD1.n5 VDD1.n3 35.4405
R110 VDD1.n4 VDD1.t1 3.6005
R111 VDD1.n4 VDD1.t6 3.6005
R112 VDD1.n0 VDD1.t5 3.6005
R113 VDD1.n0 VDD1.t4 3.6005
R114 VDD1.n2 VDD1.t2 3.6005
R115 VDD1.n2 VDD1.t3 3.6005
R116 VDD1.n1 VDD1.t0 3.6005
R117 VDD1.n1 VDD1.t7 3.6005
R118 VDD1 VDD1.n5 0.653517
R119 B.n547 B.n546 585
R120 B.n548 B.n547 585
R121 B.n200 B.n89 585
R122 B.n199 B.n198 585
R123 B.n197 B.n196 585
R124 B.n195 B.n194 585
R125 B.n193 B.n192 585
R126 B.n191 B.n190 585
R127 B.n189 B.n188 585
R128 B.n187 B.n186 585
R129 B.n185 B.n184 585
R130 B.n183 B.n182 585
R131 B.n181 B.n180 585
R132 B.n179 B.n178 585
R133 B.n177 B.n176 585
R134 B.n175 B.n174 585
R135 B.n173 B.n172 585
R136 B.n171 B.n170 585
R137 B.n169 B.n168 585
R138 B.n167 B.n166 585
R139 B.n165 B.n164 585
R140 B.n163 B.n162 585
R141 B.n161 B.n160 585
R142 B.n159 B.n158 585
R143 B.n157 B.n156 585
R144 B.n155 B.n154 585
R145 B.n153 B.n152 585
R146 B.n151 B.n150 585
R147 B.n149 B.n148 585
R148 B.n147 B.n146 585
R149 B.n145 B.n144 585
R150 B.n143 B.n142 585
R151 B.n141 B.n140 585
R152 B.n138 B.n137 585
R153 B.n136 B.n135 585
R154 B.n134 B.n133 585
R155 B.n132 B.n131 585
R156 B.n130 B.n129 585
R157 B.n128 B.n127 585
R158 B.n126 B.n125 585
R159 B.n124 B.n123 585
R160 B.n122 B.n121 585
R161 B.n120 B.n119 585
R162 B.n118 B.n117 585
R163 B.n116 B.n115 585
R164 B.n114 B.n113 585
R165 B.n112 B.n111 585
R166 B.n110 B.n109 585
R167 B.n108 B.n107 585
R168 B.n106 B.n105 585
R169 B.n104 B.n103 585
R170 B.n102 B.n101 585
R171 B.n100 B.n99 585
R172 B.n98 B.n97 585
R173 B.n96 B.n95 585
R174 B.n60 B.n59 585
R175 B.n545 B.n61 585
R176 B.n549 B.n61 585
R177 B.n544 B.n543 585
R178 B.n543 B.n57 585
R179 B.n542 B.n56 585
R180 B.n555 B.n56 585
R181 B.n541 B.n55 585
R182 B.n556 B.n55 585
R183 B.n540 B.n54 585
R184 B.n557 B.n54 585
R185 B.n539 B.n538 585
R186 B.n538 B.n53 585
R187 B.n537 B.n49 585
R188 B.n563 B.n49 585
R189 B.n536 B.n48 585
R190 B.n564 B.n48 585
R191 B.n535 B.n47 585
R192 B.n565 B.n47 585
R193 B.n534 B.n533 585
R194 B.n533 B.n43 585
R195 B.n532 B.n42 585
R196 B.n571 B.n42 585
R197 B.n531 B.n41 585
R198 B.n572 B.n41 585
R199 B.n530 B.n40 585
R200 B.n573 B.n40 585
R201 B.n529 B.n528 585
R202 B.n528 B.n39 585
R203 B.n527 B.n35 585
R204 B.n579 B.n35 585
R205 B.n526 B.n34 585
R206 B.n580 B.n34 585
R207 B.n525 B.n33 585
R208 B.n581 B.n33 585
R209 B.n524 B.n523 585
R210 B.n523 B.n29 585
R211 B.n522 B.n28 585
R212 B.n587 B.n28 585
R213 B.n521 B.n27 585
R214 B.n588 B.n27 585
R215 B.n520 B.n26 585
R216 B.n589 B.n26 585
R217 B.n519 B.n518 585
R218 B.n518 B.n22 585
R219 B.n517 B.n21 585
R220 B.n595 B.n21 585
R221 B.n516 B.n20 585
R222 B.n596 B.n20 585
R223 B.n515 B.n19 585
R224 B.n597 B.n19 585
R225 B.n514 B.n513 585
R226 B.n513 B.n15 585
R227 B.n512 B.n14 585
R228 B.n603 B.n14 585
R229 B.n511 B.n13 585
R230 B.n604 B.n13 585
R231 B.n510 B.n12 585
R232 B.n605 B.n12 585
R233 B.n509 B.n508 585
R234 B.n508 B.n507 585
R235 B.n506 B.n505 585
R236 B.n506 B.n8 585
R237 B.n504 B.n7 585
R238 B.n612 B.n7 585
R239 B.n503 B.n6 585
R240 B.n613 B.n6 585
R241 B.n502 B.n5 585
R242 B.n614 B.n5 585
R243 B.n501 B.n500 585
R244 B.n500 B.n4 585
R245 B.n499 B.n201 585
R246 B.n499 B.n498 585
R247 B.n489 B.n202 585
R248 B.n203 B.n202 585
R249 B.n491 B.n490 585
R250 B.n492 B.n491 585
R251 B.n488 B.n208 585
R252 B.n208 B.n207 585
R253 B.n487 B.n486 585
R254 B.n486 B.n485 585
R255 B.n210 B.n209 585
R256 B.n211 B.n210 585
R257 B.n478 B.n477 585
R258 B.n479 B.n478 585
R259 B.n476 B.n215 585
R260 B.n219 B.n215 585
R261 B.n475 B.n474 585
R262 B.n474 B.n473 585
R263 B.n217 B.n216 585
R264 B.n218 B.n217 585
R265 B.n466 B.n465 585
R266 B.n467 B.n466 585
R267 B.n464 B.n224 585
R268 B.n224 B.n223 585
R269 B.n463 B.n462 585
R270 B.n462 B.n461 585
R271 B.n226 B.n225 585
R272 B.n227 B.n226 585
R273 B.n454 B.n453 585
R274 B.n455 B.n454 585
R275 B.n452 B.n232 585
R276 B.n232 B.n231 585
R277 B.n451 B.n450 585
R278 B.n450 B.n449 585
R279 B.n234 B.n233 585
R280 B.n442 B.n234 585
R281 B.n441 B.n440 585
R282 B.n443 B.n441 585
R283 B.n439 B.n239 585
R284 B.n239 B.n238 585
R285 B.n438 B.n437 585
R286 B.n437 B.n436 585
R287 B.n241 B.n240 585
R288 B.n242 B.n241 585
R289 B.n429 B.n428 585
R290 B.n430 B.n429 585
R291 B.n427 B.n247 585
R292 B.n247 B.n246 585
R293 B.n426 B.n425 585
R294 B.n425 B.n424 585
R295 B.n249 B.n248 585
R296 B.n417 B.n249 585
R297 B.n416 B.n415 585
R298 B.n418 B.n416 585
R299 B.n414 B.n254 585
R300 B.n254 B.n253 585
R301 B.n413 B.n412 585
R302 B.n412 B.n411 585
R303 B.n256 B.n255 585
R304 B.n257 B.n256 585
R305 B.n404 B.n403 585
R306 B.n405 B.n404 585
R307 B.n260 B.n259 585
R308 B.n293 B.n292 585
R309 B.n294 B.n290 585
R310 B.n290 B.n261 585
R311 B.n296 B.n295 585
R312 B.n298 B.n289 585
R313 B.n301 B.n300 585
R314 B.n302 B.n288 585
R315 B.n304 B.n303 585
R316 B.n306 B.n287 585
R317 B.n309 B.n308 585
R318 B.n310 B.n286 585
R319 B.n312 B.n311 585
R320 B.n314 B.n285 585
R321 B.n317 B.n316 585
R322 B.n318 B.n284 585
R323 B.n320 B.n319 585
R324 B.n322 B.n283 585
R325 B.n325 B.n324 585
R326 B.n326 B.n282 585
R327 B.n328 B.n327 585
R328 B.n330 B.n281 585
R329 B.n333 B.n332 585
R330 B.n334 B.n278 585
R331 B.n337 B.n336 585
R332 B.n339 B.n277 585
R333 B.n342 B.n341 585
R334 B.n343 B.n276 585
R335 B.n345 B.n344 585
R336 B.n347 B.n275 585
R337 B.n350 B.n349 585
R338 B.n351 B.n274 585
R339 B.n356 B.n355 585
R340 B.n358 B.n273 585
R341 B.n361 B.n360 585
R342 B.n362 B.n272 585
R343 B.n364 B.n363 585
R344 B.n366 B.n271 585
R345 B.n369 B.n368 585
R346 B.n370 B.n270 585
R347 B.n372 B.n371 585
R348 B.n374 B.n269 585
R349 B.n377 B.n376 585
R350 B.n378 B.n268 585
R351 B.n380 B.n379 585
R352 B.n382 B.n267 585
R353 B.n385 B.n384 585
R354 B.n386 B.n266 585
R355 B.n388 B.n387 585
R356 B.n390 B.n265 585
R357 B.n393 B.n392 585
R358 B.n394 B.n264 585
R359 B.n396 B.n395 585
R360 B.n398 B.n263 585
R361 B.n401 B.n400 585
R362 B.n402 B.n262 585
R363 B.n407 B.n406 585
R364 B.n406 B.n405 585
R365 B.n408 B.n258 585
R366 B.n258 B.n257 585
R367 B.n410 B.n409 585
R368 B.n411 B.n410 585
R369 B.n252 B.n251 585
R370 B.n253 B.n252 585
R371 B.n420 B.n419 585
R372 B.n419 B.n418 585
R373 B.n421 B.n250 585
R374 B.n417 B.n250 585
R375 B.n423 B.n422 585
R376 B.n424 B.n423 585
R377 B.n245 B.n244 585
R378 B.n246 B.n245 585
R379 B.n432 B.n431 585
R380 B.n431 B.n430 585
R381 B.n433 B.n243 585
R382 B.n243 B.n242 585
R383 B.n435 B.n434 585
R384 B.n436 B.n435 585
R385 B.n237 B.n236 585
R386 B.n238 B.n237 585
R387 B.n445 B.n444 585
R388 B.n444 B.n443 585
R389 B.n446 B.n235 585
R390 B.n442 B.n235 585
R391 B.n448 B.n447 585
R392 B.n449 B.n448 585
R393 B.n230 B.n229 585
R394 B.n231 B.n230 585
R395 B.n457 B.n456 585
R396 B.n456 B.n455 585
R397 B.n458 B.n228 585
R398 B.n228 B.n227 585
R399 B.n460 B.n459 585
R400 B.n461 B.n460 585
R401 B.n222 B.n221 585
R402 B.n223 B.n222 585
R403 B.n469 B.n468 585
R404 B.n468 B.n467 585
R405 B.n470 B.n220 585
R406 B.n220 B.n218 585
R407 B.n472 B.n471 585
R408 B.n473 B.n472 585
R409 B.n214 B.n213 585
R410 B.n219 B.n214 585
R411 B.n481 B.n480 585
R412 B.n480 B.n479 585
R413 B.n482 B.n212 585
R414 B.n212 B.n211 585
R415 B.n484 B.n483 585
R416 B.n485 B.n484 585
R417 B.n206 B.n205 585
R418 B.n207 B.n206 585
R419 B.n494 B.n493 585
R420 B.n493 B.n492 585
R421 B.n495 B.n204 585
R422 B.n204 B.n203 585
R423 B.n497 B.n496 585
R424 B.n498 B.n497 585
R425 B.n3 B.n0 585
R426 B.n4 B.n3 585
R427 B.n611 B.n1 585
R428 B.n612 B.n611 585
R429 B.n610 B.n609 585
R430 B.n610 B.n8 585
R431 B.n608 B.n9 585
R432 B.n507 B.n9 585
R433 B.n607 B.n606 585
R434 B.n606 B.n605 585
R435 B.n11 B.n10 585
R436 B.n604 B.n11 585
R437 B.n602 B.n601 585
R438 B.n603 B.n602 585
R439 B.n600 B.n16 585
R440 B.n16 B.n15 585
R441 B.n599 B.n598 585
R442 B.n598 B.n597 585
R443 B.n18 B.n17 585
R444 B.n596 B.n18 585
R445 B.n594 B.n593 585
R446 B.n595 B.n594 585
R447 B.n592 B.n23 585
R448 B.n23 B.n22 585
R449 B.n591 B.n590 585
R450 B.n590 B.n589 585
R451 B.n25 B.n24 585
R452 B.n588 B.n25 585
R453 B.n586 B.n585 585
R454 B.n587 B.n586 585
R455 B.n584 B.n30 585
R456 B.n30 B.n29 585
R457 B.n583 B.n582 585
R458 B.n582 B.n581 585
R459 B.n32 B.n31 585
R460 B.n580 B.n32 585
R461 B.n578 B.n577 585
R462 B.n579 B.n578 585
R463 B.n576 B.n36 585
R464 B.n39 B.n36 585
R465 B.n575 B.n574 585
R466 B.n574 B.n573 585
R467 B.n38 B.n37 585
R468 B.n572 B.n38 585
R469 B.n570 B.n569 585
R470 B.n571 B.n570 585
R471 B.n568 B.n44 585
R472 B.n44 B.n43 585
R473 B.n567 B.n566 585
R474 B.n566 B.n565 585
R475 B.n46 B.n45 585
R476 B.n564 B.n46 585
R477 B.n562 B.n561 585
R478 B.n563 B.n562 585
R479 B.n560 B.n50 585
R480 B.n53 B.n50 585
R481 B.n559 B.n558 585
R482 B.n558 B.n557 585
R483 B.n52 B.n51 585
R484 B.n556 B.n52 585
R485 B.n554 B.n553 585
R486 B.n555 B.n554 585
R487 B.n552 B.n58 585
R488 B.n58 B.n57 585
R489 B.n551 B.n550 585
R490 B.n550 B.n549 585
R491 B.n615 B.n614 585
R492 B.n613 B.n2 585
R493 B.n550 B.n60 444.452
R494 B.n547 B.n61 444.452
R495 B.n404 B.n262 444.452
R496 B.n406 B.n260 444.452
R497 B.n93 B.t17 305.118
R498 B.n90 B.t10 305.118
R499 B.n352 B.t6 305.118
R500 B.n279 B.t14 305.118
R501 B.n548 B.n88 256.663
R502 B.n548 B.n87 256.663
R503 B.n548 B.n86 256.663
R504 B.n548 B.n85 256.663
R505 B.n548 B.n84 256.663
R506 B.n548 B.n83 256.663
R507 B.n548 B.n82 256.663
R508 B.n548 B.n81 256.663
R509 B.n548 B.n80 256.663
R510 B.n548 B.n79 256.663
R511 B.n548 B.n78 256.663
R512 B.n548 B.n77 256.663
R513 B.n548 B.n76 256.663
R514 B.n548 B.n75 256.663
R515 B.n548 B.n74 256.663
R516 B.n548 B.n73 256.663
R517 B.n548 B.n72 256.663
R518 B.n548 B.n71 256.663
R519 B.n548 B.n70 256.663
R520 B.n548 B.n69 256.663
R521 B.n548 B.n68 256.663
R522 B.n548 B.n67 256.663
R523 B.n548 B.n66 256.663
R524 B.n548 B.n65 256.663
R525 B.n548 B.n64 256.663
R526 B.n548 B.n63 256.663
R527 B.n548 B.n62 256.663
R528 B.n291 B.n261 256.663
R529 B.n297 B.n261 256.663
R530 B.n299 B.n261 256.663
R531 B.n305 B.n261 256.663
R532 B.n307 B.n261 256.663
R533 B.n313 B.n261 256.663
R534 B.n315 B.n261 256.663
R535 B.n321 B.n261 256.663
R536 B.n323 B.n261 256.663
R537 B.n329 B.n261 256.663
R538 B.n331 B.n261 256.663
R539 B.n338 B.n261 256.663
R540 B.n340 B.n261 256.663
R541 B.n346 B.n261 256.663
R542 B.n348 B.n261 256.663
R543 B.n357 B.n261 256.663
R544 B.n359 B.n261 256.663
R545 B.n365 B.n261 256.663
R546 B.n367 B.n261 256.663
R547 B.n373 B.n261 256.663
R548 B.n375 B.n261 256.663
R549 B.n381 B.n261 256.663
R550 B.n383 B.n261 256.663
R551 B.n389 B.n261 256.663
R552 B.n391 B.n261 256.663
R553 B.n397 B.n261 256.663
R554 B.n399 B.n261 256.663
R555 B.n617 B.n616 256.663
R556 B.n97 B.n96 163.367
R557 B.n101 B.n100 163.367
R558 B.n105 B.n104 163.367
R559 B.n109 B.n108 163.367
R560 B.n113 B.n112 163.367
R561 B.n117 B.n116 163.367
R562 B.n121 B.n120 163.367
R563 B.n125 B.n124 163.367
R564 B.n129 B.n128 163.367
R565 B.n133 B.n132 163.367
R566 B.n137 B.n136 163.367
R567 B.n142 B.n141 163.367
R568 B.n146 B.n145 163.367
R569 B.n150 B.n149 163.367
R570 B.n154 B.n153 163.367
R571 B.n158 B.n157 163.367
R572 B.n162 B.n161 163.367
R573 B.n166 B.n165 163.367
R574 B.n170 B.n169 163.367
R575 B.n174 B.n173 163.367
R576 B.n178 B.n177 163.367
R577 B.n182 B.n181 163.367
R578 B.n186 B.n185 163.367
R579 B.n190 B.n189 163.367
R580 B.n194 B.n193 163.367
R581 B.n198 B.n197 163.367
R582 B.n547 B.n89 163.367
R583 B.n404 B.n256 163.367
R584 B.n412 B.n256 163.367
R585 B.n412 B.n254 163.367
R586 B.n416 B.n254 163.367
R587 B.n416 B.n249 163.367
R588 B.n425 B.n249 163.367
R589 B.n425 B.n247 163.367
R590 B.n429 B.n247 163.367
R591 B.n429 B.n241 163.367
R592 B.n437 B.n241 163.367
R593 B.n437 B.n239 163.367
R594 B.n441 B.n239 163.367
R595 B.n441 B.n234 163.367
R596 B.n450 B.n234 163.367
R597 B.n450 B.n232 163.367
R598 B.n454 B.n232 163.367
R599 B.n454 B.n226 163.367
R600 B.n462 B.n226 163.367
R601 B.n462 B.n224 163.367
R602 B.n466 B.n224 163.367
R603 B.n466 B.n217 163.367
R604 B.n474 B.n217 163.367
R605 B.n474 B.n215 163.367
R606 B.n478 B.n215 163.367
R607 B.n478 B.n210 163.367
R608 B.n486 B.n210 163.367
R609 B.n486 B.n208 163.367
R610 B.n491 B.n208 163.367
R611 B.n491 B.n202 163.367
R612 B.n499 B.n202 163.367
R613 B.n500 B.n499 163.367
R614 B.n500 B.n5 163.367
R615 B.n6 B.n5 163.367
R616 B.n7 B.n6 163.367
R617 B.n506 B.n7 163.367
R618 B.n508 B.n506 163.367
R619 B.n508 B.n12 163.367
R620 B.n13 B.n12 163.367
R621 B.n14 B.n13 163.367
R622 B.n513 B.n14 163.367
R623 B.n513 B.n19 163.367
R624 B.n20 B.n19 163.367
R625 B.n21 B.n20 163.367
R626 B.n518 B.n21 163.367
R627 B.n518 B.n26 163.367
R628 B.n27 B.n26 163.367
R629 B.n28 B.n27 163.367
R630 B.n523 B.n28 163.367
R631 B.n523 B.n33 163.367
R632 B.n34 B.n33 163.367
R633 B.n35 B.n34 163.367
R634 B.n528 B.n35 163.367
R635 B.n528 B.n40 163.367
R636 B.n41 B.n40 163.367
R637 B.n42 B.n41 163.367
R638 B.n533 B.n42 163.367
R639 B.n533 B.n47 163.367
R640 B.n48 B.n47 163.367
R641 B.n49 B.n48 163.367
R642 B.n538 B.n49 163.367
R643 B.n538 B.n54 163.367
R644 B.n55 B.n54 163.367
R645 B.n56 B.n55 163.367
R646 B.n543 B.n56 163.367
R647 B.n543 B.n61 163.367
R648 B.n292 B.n290 163.367
R649 B.n296 B.n290 163.367
R650 B.n300 B.n298 163.367
R651 B.n304 B.n288 163.367
R652 B.n308 B.n306 163.367
R653 B.n312 B.n286 163.367
R654 B.n316 B.n314 163.367
R655 B.n320 B.n284 163.367
R656 B.n324 B.n322 163.367
R657 B.n328 B.n282 163.367
R658 B.n332 B.n330 163.367
R659 B.n337 B.n278 163.367
R660 B.n341 B.n339 163.367
R661 B.n345 B.n276 163.367
R662 B.n349 B.n347 163.367
R663 B.n356 B.n274 163.367
R664 B.n360 B.n358 163.367
R665 B.n364 B.n272 163.367
R666 B.n368 B.n366 163.367
R667 B.n372 B.n270 163.367
R668 B.n376 B.n374 163.367
R669 B.n380 B.n268 163.367
R670 B.n384 B.n382 163.367
R671 B.n388 B.n266 163.367
R672 B.n392 B.n390 163.367
R673 B.n396 B.n264 163.367
R674 B.n400 B.n398 163.367
R675 B.n406 B.n258 163.367
R676 B.n410 B.n258 163.367
R677 B.n410 B.n252 163.367
R678 B.n419 B.n252 163.367
R679 B.n419 B.n250 163.367
R680 B.n423 B.n250 163.367
R681 B.n423 B.n245 163.367
R682 B.n431 B.n245 163.367
R683 B.n431 B.n243 163.367
R684 B.n435 B.n243 163.367
R685 B.n435 B.n237 163.367
R686 B.n444 B.n237 163.367
R687 B.n444 B.n235 163.367
R688 B.n448 B.n235 163.367
R689 B.n448 B.n230 163.367
R690 B.n456 B.n230 163.367
R691 B.n456 B.n228 163.367
R692 B.n460 B.n228 163.367
R693 B.n460 B.n222 163.367
R694 B.n468 B.n222 163.367
R695 B.n468 B.n220 163.367
R696 B.n472 B.n220 163.367
R697 B.n472 B.n214 163.367
R698 B.n480 B.n214 163.367
R699 B.n480 B.n212 163.367
R700 B.n484 B.n212 163.367
R701 B.n484 B.n206 163.367
R702 B.n493 B.n206 163.367
R703 B.n493 B.n204 163.367
R704 B.n497 B.n204 163.367
R705 B.n497 B.n3 163.367
R706 B.n615 B.n3 163.367
R707 B.n611 B.n2 163.367
R708 B.n611 B.n610 163.367
R709 B.n610 B.n9 163.367
R710 B.n606 B.n9 163.367
R711 B.n606 B.n11 163.367
R712 B.n602 B.n11 163.367
R713 B.n602 B.n16 163.367
R714 B.n598 B.n16 163.367
R715 B.n598 B.n18 163.367
R716 B.n594 B.n18 163.367
R717 B.n594 B.n23 163.367
R718 B.n590 B.n23 163.367
R719 B.n590 B.n25 163.367
R720 B.n586 B.n25 163.367
R721 B.n586 B.n30 163.367
R722 B.n582 B.n30 163.367
R723 B.n582 B.n32 163.367
R724 B.n578 B.n32 163.367
R725 B.n578 B.n36 163.367
R726 B.n574 B.n36 163.367
R727 B.n574 B.n38 163.367
R728 B.n570 B.n38 163.367
R729 B.n570 B.n44 163.367
R730 B.n566 B.n44 163.367
R731 B.n566 B.n46 163.367
R732 B.n562 B.n46 163.367
R733 B.n562 B.n50 163.367
R734 B.n558 B.n50 163.367
R735 B.n558 B.n52 163.367
R736 B.n554 B.n52 163.367
R737 B.n554 B.n58 163.367
R738 B.n550 B.n58 163.367
R739 B.n405 B.n261 117.401
R740 B.n549 B.n548 117.401
R741 B.n90 B.t12 102.928
R742 B.n352 B.t9 102.928
R743 B.n93 B.t18 102.922
R744 B.n279 B.t16 102.922
R745 B.n62 B.n60 71.676
R746 B.n97 B.n63 71.676
R747 B.n101 B.n64 71.676
R748 B.n105 B.n65 71.676
R749 B.n109 B.n66 71.676
R750 B.n113 B.n67 71.676
R751 B.n117 B.n68 71.676
R752 B.n121 B.n69 71.676
R753 B.n125 B.n70 71.676
R754 B.n129 B.n71 71.676
R755 B.n133 B.n72 71.676
R756 B.n137 B.n73 71.676
R757 B.n142 B.n74 71.676
R758 B.n146 B.n75 71.676
R759 B.n150 B.n76 71.676
R760 B.n154 B.n77 71.676
R761 B.n158 B.n78 71.676
R762 B.n162 B.n79 71.676
R763 B.n166 B.n80 71.676
R764 B.n170 B.n81 71.676
R765 B.n174 B.n82 71.676
R766 B.n178 B.n83 71.676
R767 B.n182 B.n84 71.676
R768 B.n186 B.n85 71.676
R769 B.n190 B.n86 71.676
R770 B.n194 B.n87 71.676
R771 B.n198 B.n88 71.676
R772 B.n89 B.n88 71.676
R773 B.n197 B.n87 71.676
R774 B.n193 B.n86 71.676
R775 B.n189 B.n85 71.676
R776 B.n185 B.n84 71.676
R777 B.n181 B.n83 71.676
R778 B.n177 B.n82 71.676
R779 B.n173 B.n81 71.676
R780 B.n169 B.n80 71.676
R781 B.n165 B.n79 71.676
R782 B.n161 B.n78 71.676
R783 B.n157 B.n77 71.676
R784 B.n153 B.n76 71.676
R785 B.n149 B.n75 71.676
R786 B.n145 B.n74 71.676
R787 B.n141 B.n73 71.676
R788 B.n136 B.n72 71.676
R789 B.n132 B.n71 71.676
R790 B.n128 B.n70 71.676
R791 B.n124 B.n69 71.676
R792 B.n120 B.n68 71.676
R793 B.n116 B.n67 71.676
R794 B.n112 B.n66 71.676
R795 B.n108 B.n65 71.676
R796 B.n104 B.n64 71.676
R797 B.n100 B.n63 71.676
R798 B.n96 B.n62 71.676
R799 B.n291 B.n260 71.676
R800 B.n297 B.n296 71.676
R801 B.n300 B.n299 71.676
R802 B.n305 B.n304 71.676
R803 B.n308 B.n307 71.676
R804 B.n313 B.n312 71.676
R805 B.n316 B.n315 71.676
R806 B.n321 B.n320 71.676
R807 B.n324 B.n323 71.676
R808 B.n329 B.n328 71.676
R809 B.n332 B.n331 71.676
R810 B.n338 B.n337 71.676
R811 B.n341 B.n340 71.676
R812 B.n346 B.n345 71.676
R813 B.n349 B.n348 71.676
R814 B.n357 B.n356 71.676
R815 B.n360 B.n359 71.676
R816 B.n365 B.n364 71.676
R817 B.n368 B.n367 71.676
R818 B.n373 B.n372 71.676
R819 B.n376 B.n375 71.676
R820 B.n381 B.n380 71.676
R821 B.n384 B.n383 71.676
R822 B.n389 B.n388 71.676
R823 B.n392 B.n391 71.676
R824 B.n397 B.n396 71.676
R825 B.n400 B.n399 71.676
R826 B.n292 B.n291 71.676
R827 B.n298 B.n297 71.676
R828 B.n299 B.n288 71.676
R829 B.n306 B.n305 71.676
R830 B.n307 B.n286 71.676
R831 B.n314 B.n313 71.676
R832 B.n315 B.n284 71.676
R833 B.n322 B.n321 71.676
R834 B.n323 B.n282 71.676
R835 B.n330 B.n329 71.676
R836 B.n331 B.n278 71.676
R837 B.n339 B.n338 71.676
R838 B.n340 B.n276 71.676
R839 B.n347 B.n346 71.676
R840 B.n348 B.n274 71.676
R841 B.n358 B.n357 71.676
R842 B.n359 B.n272 71.676
R843 B.n366 B.n365 71.676
R844 B.n367 B.n270 71.676
R845 B.n374 B.n373 71.676
R846 B.n375 B.n268 71.676
R847 B.n382 B.n381 71.676
R848 B.n383 B.n266 71.676
R849 B.n390 B.n389 71.676
R850 B.n391 B.n264 71.676
R851 B.n398 B.n397 71.676
R852 B.n399 B.n262 71.676
R853 B.n616 B.n615 71.676
R854 B.n616 B.n2 71.676
R855 B.n91 B.t13 70.928
R856 B.n353 B.t8 70.928
R857 B.n94 B.t19 70.9222
R858 B.n280 B.t15 70.9222
R859 B.n405 B.n257 69.4205
R860 B.n411 B.n257 69.4205
R861 B.n411 B.n253 69.4205
R862 B.n418 B.n253 69.4205
R863 B.n418 B.n417 69.4205
R864 B.n424 B.n246 69.4205
R865 B.n430 B.n246 69.4205
R866 B.n430 B.n242 69.4205
R867 B.n436 B.n242 69.4205
R868 B.n436 B.n238 69.4205
R869 B.n443 B.n238 69.4205
R870 B.n443 B.n442 69.4205
R871 B.n449 B.n231 69.4205
R872 B.n455 B.n231 69.4205
R873 B.n455 B.n227 69.4205
R874 B.n461 B.n227 69.4205
R875 B.n467 B.n223 69.4205
R876 B.n467 B.n218 69.4205
R877 B.n473 B.n218 69.4205
R878 B.n473 B.n219 69.4205
R879 B.n479 B.n211 69.4205
R880 B.n485 B.n211 69.4205
R881 B.n485 B.n207 69.4205
R882 B.n492 B.n207 69.4205
R883 B.n498 B.n203 69.4205
R884 B.n498 B.n4 69.4205
R885 B.n614 B.n4 69.4205
R886 B.n614 B.n613 69.4205
R887 B.n613 B.n612 69.4205
R888 B.n612 B.n8 69.4205
R889 B.n507 B.n8 69.4205
R890 B.n605 B.n604 69.4205
R891 B.n604 B.n603 69.4205
R892 B.n603 B.n15 69.4205
R893 B.n597 B.n15 69.4205
R894 B.n596 B.n595 69.4205
R895 B.n595 B.n22 69.4205
R896 B.n589 B.n22 69.4205
R897 B.n589 B.n588 69.4205
R898 B.n587 B.n29 69.4205
R899 B.n581 B.n29 69.4205
R900 B.n581 B.n580 69.4205
R901 B.n580 B.n579 69.4205
R902 B.n573 B.n39 69.4205
R903 B.n573 B.n572 69.4205
R904 B.n572 B.n571 69.4205
R905 B.n571 B.n43 69.4205
R906 B.n565 B.n43 69.4205
R907 B.n565 B.n564 69.4205
R908 B.n564 B.n563 69.4205
R909 B.n557 B.n53 69.4205
R910 B.n557 B.n556 69.4205
R911 B.n556 B.n555 69.4205
R912 B.n555 B.n57 69.4205
R913 B.n549 B.n57 69.4205
R914 B.n442 B.t4 63.2952
R915 B.n39 B.t2 63.2952
R916 B.n139 B.n94 59.5399
R917 B.n92 B.n91 59.5399
R918 B.n354 B.n353 59.5399
R919 B.n335 B.n280 59.5399
R920 B.n417 B.t7 59.2116
R921 B.n53 B.t11 59.2116
R922 B.n461 B.t3 53.0863
R923 B.t21 B.n587 53.0863
R924 B.n219 B.t1 42.8775
R925 B.t20 B.n596 42.8775
R926 B.t0 B.n203 36.7522
R927 B.n507 B.t5 36.7522
R928 B.n492 B.t0 32.6687
R929 B.n605 B.t5 32.6687
R930 B.n94 B.n93 32.0005
R931 B.n91 B.n90 32.0005
R932 B.n353 B.n352 32.0005
R933 B.n280 B.n279 32.0005
R934 B.n546 B.n545 28.8785
R935 B.n407 B.n259 28.8785
R936 B.n403 B.n402 28.8785
R937 B.n551 B.n59 28.8785
R938 B.n479 B.t1 26.5434
R939 B.n597 B.t20 26.5434
R940 B B.n617 18.0485
R941 B.t3 B.n223 16.3346
R942 B.n588 B.t21 16.3346
R943 B.n408 B.n407 10.6151
R944 B.n409 B.n408 10.6151
R945 B.n409 B.n251 10.6151
R946 B.n420 B.n251 10.6151
R947 B.n421 B.n420 10.6151
R948 B.n422 B.n421 10.6151
R949 B.n422 B.n244 10.6151
R950 B.n432 B.n244 10.6151
R951 B.n433 B.n432 10.6151
R952 B.n434 B.n433 10.6151
R953 B.n434 B.n236 10.6151
R954 B.n445 B.n236 10.6151
R955 B.n446 B.n445 10.6151
R956 B.n447 B.n446 10.6151
R957 B.n447 B.n229 10.6151
R958 B.n457 B.n229 10.6151
R959 B.n458 B.n457 10.6151
R960 B.n459 B.n458 10.6151
R961 B.n459 B.n221 10.6151
R962 B.n469 B.n221 10.6151
R963 B.n470 B.n469 10.6151
R964 B.n471 B.n470 10.6151
R965 B.n471 B.n213 10.6151
R966 B.n481 B.n213 10.6151
R967 B.n482 B.n481 10.6151
R968 B.n483 B.n482 10.6151
R969 B.n483 B.n205 10.6151
R970 B.n494 B.n205 10.6151
R971 B.n495 B.n494 10.6151
R972 B.n496 B.n495 10.6151
R973 B.n496 B.n0 10.6151
R974 B.n293 B.n259 10.6151
R975 B.n294 B.n293 10.6151
R976 B.n295 B.n294 10.6151
R977 B.n295 B.n289 10.6151
R978 B.n301 B.n289 10.6151
R979 B.n302 B.n301 10.6151
R980 B.n303 B.n302 10.6151
R981 B.n303 B.n287 10.6151
R982 B.n309 B.n287 10.6151
R983 B.n310 B.n309 10.6151
R984 B.n311 B.n310 10.6151
R985 B.n311 B.n285 10.6151
R986 B.n317 B.n285 10.6151
R987 B.n318 B.n317 10.6151
R988 B.n319 B.n318 10.6151
R989 B.n319 B.n283 10.6151
R990 B.n325 B.n283 10.6151
R991 B.n326 B.n325 10.6151
R992 B.n327 B.n326 10.6151
R993 B.n327 B.n281 10.6151
R994 B.n333 B.n281 10.6151
R995 B.n334 B.n333 10.6151
R996 B.n336 B.n277 10.6151
R997 B.n342 B.n277 10.6151
R998 B.n343 B.n342 10.6151
R999 B.n344 B.n343 10.6151
R1000 B.n344 B.n275 10.6151
R1001 B.n350 B.n275 10.6151
R1002 B.n351 B.n350 10.6151
R1003 B.n355 B.n351 10.6151
R1004 B.n361 B.n273 10.6151
R1005 B.n362 B.n361 10.6151
R1006 B.n363 B.n362 10.6151
R1007 B.n363 B.n271 10.6151
R1008 B.n369 B.n271 10.6151
R1009 B.n370 B.n369 10.6151
R1010 B.n371 B.n370 10.6151
R1011 B.n371 B.n269 10.6151
R1012 B.n377 B.n269 10.6151
R1013 B.n378 B.n377 10.6151
R1014 B.n379 B.n378 10.6151
R1015 B.n379 B.n267 10.6151
R1016 B.n385 B.n267 10.6151
R1017 B.n386 B.n385 10.6151
R1018 B.n387 B.n386 10.6151
R1019 B.n387 B.n265 10.6151
R1020 B.n393 B.n265 10.6151
R1021 B.n394 B.n393 10.6151
R1022 B.n395 B.n394 10.6151
R1023 B.n395 B.n263 10.6151
R1024 B.n401 B.n263 10.6151
R1025 B.n402 B.n401 10.6151
R1026 B.n403 B.n255 10.6151
R1027 B.n413 B.n255 10.6151
R1028 B.n414 B.n413 10.6151
R1029 B.n415 B.n414 10.6151
R1030 B.n415 B.n248 10.6151
R1031 B.n426 B.n248 10.6151
R1032 B.n427 B.n426 10.6151
R1033 B.n428 B.n427 10.6151
R1034 B.n428 B.n240 10.6151
R1035 B.n438 B.n240 10.6151
R1036 B.n439 B.n438 10.6151
R1037 B.n440 B.n439 10.6151
R1038 B.n440 B.n233 10.6151
R1039 B.n451 B.n233 10.6151
R1040 B.n452 B.n451 10.6151
R1041 B.n453 B.n452 10.6151
R1042 B.n453 B.n225 10.6151
R1043 B.n463 B.n225 10.6151
R1044 B.n464 B.n463 10.6151
R1045 B.n465 B.n464 10.6151
R1046 B.n465 B.n216 10.6151
R1047 B.n475 B.n216 10.6151
R1048 B.n476 B.n475 10.6151
R1049 B.n477 B.n476 10.6151
R1050 B.n477 B.n209 10.6151
R1051 B.n487 B.n209 10.6151
R1052 B.n488 B.n487 10.6151
R1053 B.n490 B.n488 10.6151
R1054 B.n490 B.n489 10.6151
R1055 B.n489 B.n201 10.6151
R1056 B.n501 B.n201 10.6151
R1057 B.n502 B.n501 10.6151
R1058 B.n503 B.n502 10.6151
R1059 B.n504 B.n503 10.6151
R1060 B.n505 B.n504 10.6151
R1061 B.n509 B.n505 10.6151
R1062 B.n510 B.n509 10.6151
R1063 B.n511 B.n510 10.6151
R1064 B.n512 B.n511 10.6151
R1065 B.n514 B.n512 10.6151
R1066 B.n515 B.n514 10.6151
R1067 B.n516 B.n515 10.6151
R1068 B.n517 B.n516 10.6151
R1069 B.n519 B.n517 10.6151
R1070 B.n520 B.n519 10.6151
R1071 B.n521 B.n520 10.6151
R1072 B.n522 B.n521 10.6151
R1073 B.n524 B.n522 10.6151
R1074 B.n525 B.n524 10.6151
R1075 B.n526 B.n525 10.6151
R1076 B.n527 B.n526 10.6151
R1077 B.n529 B.n527 10.6151
R1078 B.n530 B.n529 10.6151
R1079 B.n531 B.n530 10.6151
R1080 B.n532 B.n531 10.6151
R1081 B.n534 B.n532 10.6151
R1082 B.n535 B.n534 10.6151
R1083 B.n536 B.n535 10.6151
R1084 B.n537 B.n536 10.6151
R1085 B.n539 B.n537 10.6151
R1086 B.n540 B.n539 10.6151
R1087 B.n541 B.n540 10.6151
R1088 B.n542 B.n541 10.6151
R1089 B.n544 B.n542 10.6151
R1090 B.n545 B.n544 10.6151
R1091 B.n609 B.n1 10.6151
R1092 B.n609 B.n608 10.6151
R1093 B.n608 B.n607 10.6151
R1094 B.n607 B.n10 10.6151
R1095 B.n601 B.n10 10.6151
R1096 B.n601 B.n600 10.6151
R1097 B.n600 B.n599 10.6151
R1098 B.n599 B.n17 10.6151
R1099 B.n593 B.n17 10.6151
R1100 B.n593 B.n592 10.6151
R1101 B.n592 B.n591 10.6151
R1102 B.n591 B.n24 10.6151
R1103 B.n585 B.n24 10.6151
R1104 B.n585 B.n584 10.6151
R1105 B.n584 B.n583 10.6151
R1106 B.n583 B.n31 10.6151
R1107 B.n577 B.n31 10.6151
R1108 B.n577 B.n576 10.6151
R1109 B.n576 B.n575 10.6151
R1110 B.n575 B.n37 10.6151
R1111 B.n569 B.n37 10.6151
R1112 B.n569 B.n568 10.6151
R1113 B.n568 B.n567 10.6151
R1114 B.n567 B.n45 10.6151
R1115 B.n561 B.n45 10.6151
R1116 B.n561 B.n560 10.6151
R1117 B.n560 B.n559 10.6151
R1118 B.n559 B.n51 10.6151
R1119 B.n553 B.n51 10.6151
R1120 B.n553 B.n552 10.6151
R1121 B.n552 B.n551 10.6151
R1122 B.n95 B.n59 10.6151
R1123 B.n98 B.n95 10.6151
R1124 B.n99 B.n98 10.6151
R1125 B.n102 B.n99 10.6151
R1126 B.n103 B.n102 10.6151
R1127 B.n106 B.n103 10.6151
R1128 B.n107 B.n106 10.6151
R1129 B.n110 B.n107 10.6151
R1130 B.n111 B.n110 10.6151
R1131 B.n114 B.n111 10.6151
R1132 B.n115 B.n114 10.6151
R1133 B.n118 B.n115 10.6151
R1134 B.n119 B.n118 10.6151
R1135 B.n122 B.n119 10.6151
R1136 B.n123 B.n122 10.6151
R1137 B.n126 B.n123 10.6151
R1138 B.n127 B.n126 10.6151
R1139 B.n130 B.n127 10.6151
R1140 B.n131 B.n130 10.6151
R1141 B.n134 B.n131 10.6151
R1142 B.n135 B.n134 10.6151
R1143 B.n138 B.n135 10.6151
R1144 B.n143 B.n140 10.6151
R1145 B.n144 B.n143 10.6151
R1146 B.n147 B.n144 10.6151
R1147 B.n148 B.n147 10.6151
R1148 B.n151 B.n148 10.6151
R1149 B.n152 B.n151 10.6151
R1150 B.n155 B.n152 10.6151
R1151 B.n156 B.n155 10.6151
R1152 B.n160 B.n159 10.6151
R1153 B.n163 B.n160 10.6151
R1154 B.n164 B.n163 10.6151
R1155 B.n167 B.n164 10.6151
R1156 B.n168 B.n167 10.6151
R1157 B.n171 B.n168 10.6151
R1158 B.n172 B.n171 10.6151
R1159 B.n175 B.n172 10.6151
R1160 B.n176 B.n175 10.6151
R1161 B.n179 B.n176 10.6151
R1162 B.n180 B.n179 10.6151
R1163 B.n183 B.n180 10.6151
R1164 B.n184 B.n183 10.6151
R1165 B.n187 B.n184 10.6151
R1166 B.n188 B.n187 10.6151
R1167 B.n191 B.n188 10.6151
R1168 B.n192 B.n191 10.6151
R1169 B.n195 B.n192 10.6151
R1170 B.n196 B.n195 10.6151
R1171 B.n199 B.n196 10.6151
R1172 B.n200 B.n199 10.6151
R1173 B.n546 B.n200 10.6151
R1174 B.n424 B.t7 10.2093
R1175 B.n563 B.t11 10.2093
R1176 B.n617 B.n0 8.11757
R1177 B.n617 B.n1 8.11757
R1178 B.n336 B.n335 6.5566
R1179 B.n355 B.n354 6.5566
R1180 B.n140 B.n139 6.5566
R1181 B.n156 B.n92 6.5566
R1182 B.n449 B.t4 6.12579
R1183 B.n579 B.t2 6.12579
R1184 B.n335 B.n334 4.05904
R1185 B.n354 B.n273 4.05904
R1186 B.n139 B.n138 4.05904
R1187 B.n159 B.n92 4.05904
R1188 VN.n18 VN.n17 174.827
R1189 VN.n37 VN.n36 174.827
R1190 VN.n35 VN.n19 161.3
R1191 VN.n34 VN.n33 161.3
R1192 VN.n32 VN.n20 161.3
R1193 VN.n31 VN.n30 161.3
R1194 VN.n29 VN.n21 161.3
R1195 VN.n28 VN.n27 161.3
R1196 VN.n26 VN.n23 161.3
R1197 VN.n16 VN.n0 161.3
R1198 VN.n15 VN.n14 161.3
R1199 VN.n13 VN.n1 161.3
R1200 VN.n12 VN.n11 161.3
R1201 VN.n9 VN.n2 161.3
R1202 VN.n8 VN.n7 161.3
R1203 VN.n6 VN.n3 161.3
R1204 VN.n5 VN.t4 128.549
R1205 VN.n25 VN.t5 128.549
R1206 VN.n4 VN.t3 100.418
R1207 VN.n10 VN.t2 100.418
R1208 VN.n17 VN.t1 100.418
R1209 VN.n24 VN.t6 100.418
R1210 VN.n22 VN.t0 100.418
R1211 VN.n36 VN.t7 100.418
R1212 VN.n5 VN.n4 61.9082
R1213 VN.n25 VN.n24 61.9082
R1214 VN.n9 VN.n8 56.5617
R1215 VN.n29 VN.n28 56.5617
R1216 VN.n15 VN.n1 50.2647
R1217 VN.n34 VN.n20 50.2647
R1218 VN VN.n37 40.26
R1219 VN.n16 VN.n15 30.8893
R1220 VN.n35 VN.n34 30.8893
R1221 VN.n26 VN.n25 27.4757
R1222 VN.n6 VN.n5 27.4757
R1223 VN.n8 VN.n3 24.5923
R1224 VN.n11 VN.n9 24.5923
R1225 VN.n28 VN.n23 24.5923
R1226 VN.n30 VN.n29 24.5923
R1227 VN.n10 VN.n1 20.9036
R1228 VN.n22 VN.n20 20.9036
R1229 VN.n17 VN.n16 11.0668
R1230 VN.n36 VN.n35 11.0668
R1231 VN.n4 VN.n3 3.68928
R1232 VN.n11 VN.n10 3.68928
R1233 VN.n24 VN.n23 3.68928
R1234 VN.n30 VN.n22 3.68928
R1235 VN.n37 VN.n19 0.189894
R1236 VN.n33 VN.n19 0.189894
R1237 VN.n33 VN.n32 0.189894
R1238 VN.n32 VN.n31 0.189894
R1239 VN.n31 VN.n21 0.189894
R1240 VN.n27 VN.n21 0.189894
R1241 VN.n27 VN.n26 0.189894
R1242 VN.n7 VN.n6 0.189894
R1243 VN.n7 VN.n2 0.189894
R1244 VN.n12 VN.n2 0.189894
R1245 VN.n13 VN.n12 0.189894
R1246 VN.n14 VN.n13 0.189894
R1247 VN.n14 VN.n0 0.189894
R1248 VN.n18 VN.n0 0.189894
R1249 VN VN.n18 0.0516364
R1250 VDD2.n2 VDD2.n1 71.8892
R1251 VDD2.n2 VDD2.n0 71.8892
R1252 VDD2 VDD2.n5 71.8855
R1253 VDD2.n4 VDD2.n3 71.2334
R1254 VDD2.n4 VDD2.n2 34.8575
R1255 VDD2.n5 VDD2.t1 3.6005
R1256 VDD2.n5 VDD2.t2 3.6005
R1257 VDD2.n3 VDD2.t0 3.6005
R1258 VDD2.n3 VDD2.t7 3.6005
R1259 VDD2.n1 VDD2.t5 3.6005
R1260 VDD2.n1 VDD2.t6 3.6005
R1261 VDD2.n0 VDD2.t3 3.6005
R1262 VDD2.n0 VDD2.t4 3.6005
R1263 VDD2 VDD2.n4 0.769897
C0 VDD2 VP 0.383613f
C1 VDD2 VTAIL 5.53495f
C2 VN VP 4.8913f
C3 VN VTAIL 3.89035f
C4 VDD2 VDD1 1.13614f
C5 VTAIL VP 3.90446f
C6 VN VDD1 0.149562f
C7 VDD1 VP 3.78312f
C8 VTAIL VDD1 5.48911f
C9 VN VDD2 3.54982f
C10 VDD2 B 3.557438f
C11 VDD1 B 3.865369f
C12 VTAIL B 5.510256f
C13 VN B 9.987261f
C14 VP B 8.502308f
C15 VDD2.t3 B 0.107718f
C16 VDD2.t4 B 0.107718f
C17 VDD2.n0 B 0.902628f
C18 VDD2.t5 B 0.107718f
C19 VDD2.t6 B 0.107718f
C20 VDD2.n1 B 0.902628f
C21 VDD2.n2 B 2.09339f
C22 VDD2.t0 B 0.107718f
C23 VDD2.t7 B 0.107718f
C24 VDD2.n3 B 0.899296f
C25 VDD2.n4 B 1.96299f
C26 VDD2.t1 B 0.107718f
C27 VDD2.t2 B 0.107718f
C28 VDD2.n5 B 0.902604f
C29 VN.n0 B 0.035236f
C30 VN.t1 B 0.673455f
C31 VN.n1 B 0.059514f
C32 VN.n2 B 0.035236f
C33 VN.n3 B 0.037923f
C34 VN.t4 B 0.757264f
C35 VN.t3 B 0.673455f
C36 VN.n4 B 0.318548f
C37 VN.n5 B 0.35001f
C38 VN.n6 B 0.185574f
C39 VN.n7 B 0.035236f
C40 VN.n8 B 0.051221f
C41 VN.n9 B 0.051221f
C42 VN.t2 B 0.673455f
C43 VN.n10 B 0.271225f
C44 VN.n11 B 0.037923f
C45 VN.n12 B 0.035236f
C46 VN.n13 B 0.035236f
C47 VN.n14 B 0.035236f
C48 VN.n15 B 0.033222f
C49 VN.n16 B 0.052466f
C50 VN.n17 B 0.33419f
C51 VN.n18 B 0.032586f
C52 VN.n19 B 0.035236f
C53 VN.t7 B 0.673455f
C54 VN.n20 B 0.059514f
C55 VN.n21 B 0.035236f
C56 VN.t0 B 0.673455f
C57 VN.n22 B 0.271225f
C58 VN.n23 B 0.037923f
C59 VN.t5 B 0.757264f
C60 VN.t6 B 0.673455f
C61 VN.n24 B 0.318548f
C62 VN.n25 B 0.35001f
C63 VN.n26 B 0.185574f
C64 VN.n27 B 0.035236f
C65 VN.n28 B 0.051221f
C66 VN.n29 B 0.051221f
C67 VN.n30 B 0.037923f
C68 VN.n31 B 0.035236f
C69 VN.n32 B 0.035236f
C70 VN.n33 B 0.035236f
C71 VN.n34 B 0.033222f
C72 VN.n35 B 0.052466f
C73 VN.n36 B 0.33419f
C74 VN.n37 B 1.36043f
C75 VDD1.t5 B 0.110188f
C76 VDD1.t4 B 0.110188f
C77 VDD1.n0 B 0.924001f
C78 VDD1.t0 B 0.110188f
C79 VDD1.t7 B 0.110188f
C80 VDD1.n1 B 0.923324f
C81 VDD1.t2 B 0.110188f
C82 VDD1.t3 B 0.110188f
C83 VDD1.n2 B 0.923324f
C84 VDD1.n3 B 2.19524f
C85 VDD1.t1 B 0.110188f
C86 VDD1.t6 B 0.110188f
C87 VDD1.n4 B 0.919913f
C88 VDD1.n5 B 2.03828f
C89 VTAIL.t6 B 0.095762f
C90 VTAIL.t7 B 0.095762f
C91 VTAIL.n0 B 0.749472f
C92 VTAIL.n1 B 0.292957f
C93 VTAIL.t5 B 0.95401f
C94 VTAIL.n2 B 0.378813f
C95 VTAIL.t14 B 0.95401f
C96 VTAIL.n3 B 0.378813f
C97 VTAIL.t11 B 0.095762f
C98 VTAIL.t15 B 0.095762f
C99 VTAIL.n4 B 0.749472f
C100 VTAIL.n5 B 0.389811f
C101 VTAIL.t10 B 0.95401f
C102 VTAIL.n6 B 1.08236f
C103 VTAIL.t4 B 0.95401f
C104 VTAIL.n7 B 1.08236f
C105 VTAIL.t3 B 0.095762f
C106 VTAIL.t1 B 0.095762f
C107 VTAIL.n8 B 0.749475f
C108 VTAIL.n9 B 0.389808f
C109 VTAIL.t0 B 0.95401f
C110 VTAIL.n10 B 0.378813f
C111 VTAIL.t8 B 0.95401f
C112 VTAIL.n11 B 0.378813f
C113 VTAIL.t13 B 0.095762f
C114 VTAIL.t9 B 0.095762f
C115 VTAIL.n12 B 0.749475f
C116 VTAIL.n13 B 0.389808f
C117 VTAIL.t12 B 0.954006f
C118 VTAIL.n14 B 1.08236f
C119 VTAIL.t2 B 0.95401f
C120 VTAIL.n15 B 1.07823f
C121 VP.n0 B 0.036241f
C122 VP.t4 B 0.69267f
C123 VP.n1 B 0.061212f
C124 VP.n2 B 0.036241f
C125 VP.n3 B 0.039005f
C126 VP.n4 B 0.036241f
C127 VP.t7 B 0.69267f
C128 VP.n5 B 0.343725f
C129 VP.n6 B 0.036241f
C130 VP.t1 B 0.69267f
C131 VP.n7 B 0.061212f
C132 VP.n8 B 0.036241f
C133 VP.n9 B 0.039005f
C134 VP.t2 B 0.778871f
C135 VP.t3 B 0.69267f
C136 VP.n10 B 0.327637f
C137 VP.n11 B 0.359997f
C138 VP.n12 B 0.190869f
C139 VP.n13 B 0.036241f
C140 VP.n14 B 0.052682f
C141 VP.n15 B 0.052682f
C142 VP.t6 B 0.69267f
C143 VP.n16 B 0.278964f
C144 VP.n17 B 0.039005f
C145 VP.n18 B 0.036241f
C146 VP.n19 B 0.036241f
C147 VP.n20 B 0.036241f
C148 VP.n21 B 0.03417f
C149 VP.n22 B 0.053963f
C150 VP.n23 B 0.343725f
C151 VP.n24 B 1.37538f
C152 VP.n25 B 1.40814f
C153 VP.n26 B 0.036241f
C154 VP.n27 B 0.053963f
C155 VP.n28 B 0.03417f
C156 VP.t0 B 0.69267f
C157 VP.n29 B 0.278964f
C158 VP.n30 B 0.061212f
C159 VP.n31 B 0.036241f
C160 VP.n32 B 0.036241f
C161 VP.n33 B 0.036241f
C162 VP.n34 B 0.052682f
C163 VP.n35 B 0.052682f
C164 VP.t5 B 0.69267f
C165 VP.n36 B 0.278964f
C166 VP.n37 B 0.039005f
C167 VP.n38 B 0.036241f
C168 VP.n39 B 0.036241f
C169 VP.n40 B 0.036241f
C170 VP.n41 B 0.03417f
C171 VP.n42 B 0.053963f
C172 VP.n43 B 0.343725f
C173 VP.n44 B 0.033516f
.ends

