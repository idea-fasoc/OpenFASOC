* NGSPICE file created from diff_pair_sample_0444.ext - technology: sky130A

.subckt diff_pair_sample_0444 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X1 VDD2.t6 VN.t1 VTAIL.t8 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X2 VTAIL.t14 VN.t2 VDD2.t5 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X3 VTAIL.t2 VP.t0 VDD1.t7 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X4 VDD1.t6 VP.t1 VTAIL.t7 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X5 VDD1.t5 VP.t2 VTAIL.t4 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=5.5068 ps=29.02 w=14.12 l=0.4
X6 VTAIL.t11 VN.t3 VDD2.t4 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X7 B.t11 B.t9 B.t10 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=0 ps=0 w=14.12 l=0.4
X8 B.t8 B.t6 B.t7 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=0 ps=0 w=14.12 l=0.4
X9 VDD2.t3 VN.t4 VTAIL.t13 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=5.5068 ps=29.02 w=14.12 l=0.4
X10 VTAIL.t0 VP.t3 VDD1.t4 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X11 VDD2.t2 VN.t5 VTAIL.t9 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=5.5068 ps=29.02 w=14.12 l=0.4
X12 VTAIL.t6 VP.t4 VDD1.t3 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=2.3298 ps=14.45 w=14.12 l=0.4
X13 VTAIL.t1 VP.t5 VDD1.t2 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=2.3298 ps=14.45 w=14.12 l=0.4
X14 B.t5 B.t3 B.t4 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=0 ps=0 w=14.12 l=0.4
X15 VDD1.t1 VP.t6 VTAIL.t3 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=2.3298 ps=14.45 w=14.12 l=0.4
X16 VTAIL.t10 VN.t6 VDD2.t1 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=2.3298 ps=14.45 w=14.12 l=0.4
X17 B.t2 B.t0 B.t1 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=0 ps=0 w=14.12 l=0.4
X18 VDD1.t0 VP.t7 VTAIL.t5 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=2.3298 pd=14.45 as=5.5068 ps=29.02 w=14.12 l=0.4
X19 VTAIL.t15 VN.t7 VDD2.t0 w_n1700_n3792# sky130_fd_pr__pfet_01v8 ad=5.5068 pd=29.02 as=2.3298 ps=14.45 w=14.12 l=0.4
R0 VN.n1 VN.t7 982.591
R1 VN.n7 VN.t4 982.591
R2 VN.n4 VN.t5 970.116
R3 VN.n10 VN.t6 970.116
R4 VN.n2 VN.t0 948.938
R5 VN.n3 VN.t3 948.938
R6 VN.n8 VN.t2 948.938
R7 VN.n9 VN.t1 948.938
R8 VN.n5 VN.n4 161.3
R9 VN.n11 VN.n10 161.3
R10 VN.n9 VN.n6 161.3
R11 VN.n3 VN.n0 161.3
R12 VN.n7 VN.n6 74.6542
R13 VN.n1 VN.n0 74.6542
R14 VN.n3 VN.n2 48.2005
R15 VN.n9 VN.n8 48.2005
R16 VN VN.n11 42.7297
R17 VN.n4 VN.n3 27.0217
R18 VN.n10 VN.n9 27.0217
R19 VN.n8 VN.n7 12.4607
R20 VN.n2 VN.n1 12.4607
R21 VN.n11 VN.n6 0.189894
R22 VN.n5 VN.n0 0.189894
R23 VN VN.n5 0.0516364
R24 VTAIL.n626 VTAIL.n554 756.745
R25 VTAIL.n74 VTAIL.n2 756.745
R26 VTAIL.n152 VTAIL.n80 756.745
R27 VTAIL.n232 VTAIL.n160 756.745
R28 VTAIL.n548 VTAIL.n476 756.745
R29 VTAIL.n468 VTAIL.n396 756.745
R30 VTAIL.n390 VTAIL.n318 756.745
R31 VTAIL.n310 VTAIL.n238 756.745
R32 VTAIL.n578 VTAIL.n577 585
R33 VTAIL.n583 VTAIL.n582 585
R34 VTAIL.n585 VTAIL.n584 585
R35 VTAIL.n574 VTAIL.n573 585
R36 VTAIL.n591 VTAIL.n590 585
R37 VTAIL.n593 VTAIL.n592 585
R38 VTAIL.n570 VTAIL.n569 585
R39 VTAIL.n599 VTAIL.n598 585
R40 VTAIL.n601 VTAIL.n600 585
R41 VTAIL.n566 VTAIL.n565 585
R42 VTAIL.n607 VTAIL.n606 585
R43 VTAIL.n609 VTAIL.n608 585
R44 VTAIL.n562 VTAIL.n561 585
R45 VTAIL.n615 VTAIL.n614 585
R46 VTAIL.n617 VTAIL.n616 585
R47 VTAIL.n558 VTAIL.n557 585
R48 VTAIL.n624 VTAIL.n623 585
R49 VTAIL.n625 VTAIL.n556 585
R50 VTAIL.n627 VTAIL.n626 585
R51 VTAIL.n26 VTAIL.n25 585
R52 VTAIL.n31 VTAIL.n30 585
R53 VTAIL.n33 VTAIL.n32 585
R54 VTAIL.n22 VTAIL.n21 585
R55 VTAIL.n39 VTAIL.n38 585
R56 VTAIL.n41 VTAIL.n40 585
R57 VTAIL.n18 VTAIL.n17 585
R58 VTAIL.n47 VTAIL.n46 585
R59 VTAIL.n49 VTAIL.n48 585
R60 VTAIL.n14 VTAIL.n13 585
R61 VTAIL.n55 VTAIL.n54 585
R62 VTAIL.n57 VTAIL.n56 585
R63 VTAIL.n10 VTAIL.n9 585
R64 VTAIL.n63 VTAIL.n62 585
R65 VTAIL.n65 VTAIL.n64 585
R66 VTAIL.n6 VTAIL.n5 585
R67 VTAIL.n72 VTAIL.n71 585
R68 VTAIL.n73 VTAIL.n4 585
R69 VTAIL.n75 VTAIL.n74 585
R70 VTAIL.n104 VTAIL.n103 585
R71 VTAIL.n109 VTAIL.n108 585
R72 VTAIL.n111 VTAIL.n110 585
R73 VTAIL.n100 VTAIL.n99 585
R74 VTAIL.n117 VTAIL.n116 585
R75 VTAIL.n119 VTAIL.n118 585
R76 VTAIL.n96 VTAIL.n95 585
R77 VTAIL.n125 VTAIL.n124 585
R78 VTAIL.n127 VTAIL.n126 585
R79 VTAIL.n92 VTAIL.n91 585
R80 VTAIL.n133 VTAIL.n132 585
R81 VTAIL.n135 VTAIL.n134 585
R82 VTAIL.n88 VTAIL.n87 585
R83 VTAIL.n141 VTAIL.n140 585
R84 VTAIL.n143 VTAIL.n142 585
R85 VTAIL.n84 VTAIL.n83 585
R86 VTAIL.n150 VTAIL.n149 585
R87 VTAIL.n151 VTAIL.n82 585
R88 VTAIL.n153 VTAIL.n152 585
R89 VTAIL.n184 VTAIL.n183 585
R90 VTAIL.n189 VTAIL.n188 585
R91 VTAIL.n191 VTAIL.n190 585
R92 VTAIL.n180 VTAIL.n179 585
R93 VTAIL.n197 VTAIL.n196 585
R94 VTAIL.n199 VTAIL.n198 585
R95 VTAIL.n176 VTAIL.n175 585
R96 VTAIL.n205 VTAIL.n204 585
R97 VTAIL.n207 VTAIL.n206 585
R98 VTAIL.n172 VTAIL.n171 585
R99 VTAIL.n213 VTAIL.n212 585
R100 VTAIL.n215 VTAIL.n214 585
R101 VTAIL.n168 VTAIL.n167 585
R102 VTAIL.n221 VTAIL.n220 585
R103 VTAIL.n223 VTAIL.n222 585
R104 VTAIL.n164 VTAIL.n163 585
R105 VTAIL.n230 VTAIL.n229 585
R106 VTAIL.n231 VTAIL.n162 585
R107 VTAIL.n233 VTAIL.n232 585
R108 VTAIL.n549 VTAIL.n548 585
R109 VTAIL.n547 VTAIL.n478 585
R110 VTAIL.n546 VTAIL.n545 585
R111 VTAIL.n481 VTAIL.n479 585
R112 VTAIL.n540 VTAIL.n539 585
R113 VTAIL.n538 VTAIL.n537 585
R114 VTAIL.n485 VTAIL.n484 585
R115 VTAIL.n532 VTAIL.n531 585
R116 VTAIL.n530 VTAIL.n529 585
R117 VTAIL.n489 VTAIL.n488 585
R118 VTAIL.n524 VTAIL.n523 585
R119 VTAIL.n522 VTAIL.n521 585
R120 VTAIL.n493 VTAIL.n492 585
R121 VTAIL.n516 VTAIL.n515 585
R122 VTAIL.n514 VTAIL.n513 585
R123 VTAIL.n497 VTAIL.n496 585
R124 VTAIL.n508 VTAIL.n507 585
R125 VTAIL.n506 VTAIL.n505 585
R126 VTAIL.n501 VTAIL.n500 585
R127 VTAIL.n469 VTAIL.n468 585
R128 VTAIL.n467 VTAIL.n398 585
R129 VTAIL.n466 VTAIL.n465 585
R130 VTAIL.n401 VTAIL.n399 585
R131 VTAIL.n460 VTAIL.n459 585
R132 VTAIL.n458 VTAIL.n457 585
R133 VTAIL.n405 VTAIL.n404 585
R134 VTAIL.n452 VTAIL.n451 585
R135 VTAIL.n450 VTAIL.n449 585
R136 VTAIL.n409 VTAIL.n408 585
R137 VTAIL.n444 VTAIL.n443 585
R138 VTAIL.n442 VTAIL.n441 585
R139 VTAIL.n413 VTAIL.n412 585
R140 VTAIL.n436 VTAIL.n435 585
R141 VTAIL.n434 VTAIL.n433 585
R142 VTAIL.n417 VTAIL.n416 585
R143 VTAIL.n428 VTAIL.n427 585
R144 VTAIL.n426 VTAIL.n425 585
R145 VTAIL.n421 VTAIL.n420 585
R146 VTAIL.n391 VTAIL.n390 585
R147 VTAIL.n389 VTAIL.n320 585
R148 VTAIL.n388 VTAIL.n387 585
R149 VTAIL.n323 VTAIL.n321 585
R150 VTAIL.n382 VTAIL.n381 585
R151 VTAIL.n380 VTAIL.n379 585
R152 VTAIL.n327 VTAIL.n326 585
R153 VTAIL.n374 VTAIL.n373 585
R154 VTAIL.n372 VTAIL.n371 585
R155 VTAIL.n331 VTAIL.n330 585
R156 VTAIL.n366 VTAIL.n365 585
R157 VTAIL.n364 VTAIL.n363 585
R158 VTAIL.n335 VTAIL.n334 585
R159 VTAIL.n358 VTAIL.n357 585
R160 VTAIL.n356 VTAIL.n355 585
R161 VTAIL.n339 VTAIL.n338 585
R162 VTAIL.n350 VTAIL.n349 585
R163 VTAIL.n348 VTAIL.n347 585
R164 VTAIL.n343 VTAIL.n342 585
R165 VTAIL.n311 VTAIL.n310 585
R166 VTAIL.n309 VTAIL.n240 585
R167 VTAIL.n308 VTAIL.n307 585
R168 VTAIL.n243 VTAIL.n241 585
R169 VTAIL.n302 VTAIL.n301 585
R170 VTAIL.n300 VTAIL.n299 585
R171 VTAIL.n247 VTAIL.n246 585
R172 VTAIL.n294 VTAIL.n293 585
R173 VTAIL.n292 VTAIL.n291 585
R174 VTAIL.n251 VTAIL.n250 585
R175 VTAIL.n286 VTAIL.n285 585
R176 VTAIL.n284 VTAIL.n283 585
R177 VTAIL.n255 VTAIL.n254 585
R178 VTAIL.n278 VTAIL.n277 585
R179 VTAIL.n276 VTAIL.n275 585
R180 VTAIL.n259 VTAIL.n258 585
R181 VTAIL.n270 VTAIL.n269 585
R182 VTAIL.n268 VTAIL.n267 585
R183 VTAIL.n263 VTAIL.n262 585
R184 VTAIL.n579 VTAIL.t9 327.466
R185 VTAIL.n27 VTAIL.t15 327.466
R186 VTAIL.n105 VTAIL.t4 327.466
R187 VTAIL.n185 VTAIL.t1 327.466
R188 VTAIL.n502 VTAIL.t5 327.466
R189 VTAIL.n422 VTAIL.t6 327.466
R190 VTAIL.n344 VTAIL.t13 327.466
R191 VTAIL.n264 VTAIL.t10 327.466
R192 VTAIL.n583 VTAIL.n577 171.744
R193 VTAIL.n584 VTAIL.n583 171.744
R194 VTAIL.n584 VTAIL.n573 171.744
R195 VTAIL.n591 VTAIL.n573 171.744
R196 VTAIL.n592 VTAIL.n591 171.744
R197 VTAIL.n592 VTAIL.n569 171.744
R198 VTAIL.n599 VTAIL.n569 171.744
R199 VTAIL.n600 VTAIL.n599 171.744
R200 VTAIL.n600 VTAIL.n565 171.744
R201 VTAIL.n607 VTAIL.n565 171.744
R202 VTAIL.n608 VTAIL.n607 171.744
R203 VTAIL.n608 VTAIL.n561 171.744
R204 VTAIL.n615 VTAIL.n561 171.744
R205 VTAIL.n616 VTAIL.n615 171.744
R206 VTAIL.n616 VTAIL.n557 171.744
R207 VTAIL.n624 VTAIL.n557 171.744
R208 VTAIL.n625 VTAIL.n624 171.744
R209 VTAIL.n626 VTAIL.n625 171.744
R210 VTAIL.n31 VTAIL.n25 171.744
R211 VTAIL.n32 VTAIL.n31 171.744
R212 VTAIL.n32 VTAIL.n21 171.744
R213 VTAIL.n39 VTAIL.n21 171.744
R214 VTAIL.n40 VTAIL.n39 171.744
R215 VTAIL.n40 VTAIL.n17 171.744
R216 VTAIL.n47 VTAIL.n17 171.744
R217 VTAIL.n48 VTAIL.n47 171.744
R218 VTAIL.n48 VTAIL.n13 171.744
R219 VTAIL.n55 VTAIL.n13 171.744
R220 VTAIL.n56 VTAIL.n55 171.744
R221 VTAIL.n56 VTAIL.n9 171.744
R222 VTAIL.n63 VTAIL.n9 171.744
R223 VTAIL.n64 VTAIL.n63 171.744
R224 VTAIL.n64 VTAIL.n5 171.744
R225 VTAIL.n72 VTAIL.n5 171.744
R226 VTAIL.n73 VTAIL.n72 171.744
R227 VTAIL.n74 VTAIL.n73 171.744
R228 VTAIL.n109 VTAIL.n103 171.744
R229 VTAIL.n110 VTAIL.n109 171.744
R230 VTAIL.n110 VTAIL.n99 171.744
R231 VTAIL.n117 VTAIL.n99 171.744
R232 VTAIL.n118 VTAIL.n117 171.744
R233 VTAIL.n118 VTAIL.n95 171.744
R234 VTAIL.n125 VTAIL.n95 171.744
R235 VTAIL.n126 VTAIL.n125 171.744
R236 VTAIL.n126 VTAIL.n91 171.744
R237 VTAIL.n133 VTAIL.n91 171.744
R238 VTAIL.n134 VTAIL.n133 171.744
R239 VTAIL.n134 VTAIL.n87 171.744
R240 VTAIL.n141 VTAIL.n87 171.744
R241 VTAIL.n142 VTAIL.n141 171.744
R242 VTAIL.n142 VTAIL.n83 171.744
R243 VTAIL.n150 VTAIL.n83 171.744
R244 VTAIL.n151 VTAIL.n150 171.744
R245 VTAIL.n152 VTAIL.n151 171.744
R246 VTAIL.n189 VTAIL.n183 171.744
R247 VTAIL.n190 VTAIL.n189 171.744
R248 VTAIL.n190 VTAIL.n179 171.744
R249 VTAIL.n197 VTAIL.n179 171.744
R250 VTAIL.n198 VTAIL.n197 171.744
R251 VTAIL.n198 VTAIL.n175 171.744
R252 VTAIL.n205 VTAIL.n175 171.744
R253 VTAIL.n206 VTAIL.n205 171.744
R254 VTAIL.n206 VTAIL.n171 171.744
R255 VTAIL.n213 VTAIL.n171 171.744
R256 VTAIL.n214 VTAIL.n213 171.744
R257 VTAIL.n214 VTAIL.n167 171.744
R258 VTAIL.n221 VTAIL.n167 171.744
R259 VTAIL.n222 VTAIL.n221 171.744
R260 VTAIL.n222 VTAIL.n163 171.744
R261 VTAIL.n230 VTAIL.n163 171.744
R262 VTAIL.n231 VTAIL.n230 171.744
R263 VTAIL.n232 VTAIL.n231 171.744
R264 VTAIL.n548 VTAIL.n547 171.744
R265 VTAIL.n547 VTAIL.n546 171.744
R266 VTAIL.n546 VTAIL.n479 171.744
R267 VTAIL.n539 VTAIL.n479 171.744
R268 VTAIL.n539 VTAIL.n538 171.744
R269 VTAIL.n538 VTAIL.n484 171.744
R270 VTAIL.n531 VTAIL.n484 171.744
R271 VTAIL.n531 VTAIL.n530 171.744
R272 VTAIL.n530 VTAIL.n488 171.744
R273 VTAIL.n523 VTAIL.n488 171.744
R274 VTAIL.n523 VTAIL.n522 171.744
R275 VTAIL.n522 VTAIL.n492 171.744
R276 VTAIL.n515 VTAIL.n492 171.744
R277 VTAIL.n515 VTAIL.n514 171.744
R278 VTAIL.n514 VTAIL.n496 171.744
R279 VTAIL.n507 VTAIL.n496 171.744
R280 VTAIL.n507 VTAIL.n506 171.744
R281 VTAIL.n506 VTAIL.n500 171.744
R282 VTAIL.n468 VTAIL.n467 171.744
R283 VTAIL.n467 VTAIL.n466 171.744
R284 VTAIL.n466 VTAIL.n399 171.744
R285 VTAIL.n459 VTAIL.n399 171.744
R286 VTAIL.n459 VTAIL.n458 171.744
R287 VTAIL.n458 VTAIL.n404 171.744
R288 VTAIL.n451 VTAIL.n404 171.744
R289 VTAIL.n451 VTAIL.n450 171.744
R290 VTAIL.n450 VTAIL.n408 171.744
R291 VTAIL.n443 VTAIL.n408 171.744
R292 VTAIL.n443 VTAIL.n442 171.744
R293 VTAIL.n442 VTAIL.n412 171.744
R294 VTAIL.n435 VTAIL.n412 171.744
R295 VTAIL.n435 VTAIL.n434 171.744
R296 VTAIL.n434 VTAIL.n416 171.744
R297 VTAIL.n427 VTAIL.n416 171.744
R298 VTAIL.n427 VTAIL.n426 171.744
R299 VTAIL.n426 VTAIL.n420 171.744
R300 VTAIL.n390 VTAIL.n389 171.744
R301 VTAIL.n389 VTAIL.n388 171.744
R302 VTAIL.n388 VTAIL.n321 171.744
R303 VTAIL.n381 VTAIL.n321 171.744
R304 VTAIL.n381 VTAIL.n380 171.744
R305 VTAIL.n380 VTAIL.n326 171.744
R306 VTAIL.n373 VTAIL.n326 171.744
R307 VTAIL.n373 VTAIL.n372 171.744
R308 VTAIL.n372 VTAIL.n330 171.744
R309 VTAIL.n365 VTAIL.n330 171.744
R310 VTAIL.n365 VTAIL.n364 171.744
R311 VTAIL.n364 VTAIL.n334 171.744
R312 VTAIL.n357 VTAIL.n334 171.744
R313 VTAIL.n357 VTAIL.n356 171.744
R314 VTAIL.n356 VTAIL.n338 171.744
R315 VTAIL.n349 VTAIL.n338 171.744
R316 VTAIL.n349 VTAIL.n348 171.744
R317 VTAIL.n348 VTAIL.n342 171.744
R318 VTAIL.n310 VTAIL.n309 171.744
R319 VTAIL.n309 VTAIL.n308 171.744
R320 VTAIL.n308 VTAIL.n241 171.744
R321 VTAIL.n301 VTAIL.n241 171.744
R322 VTAIL.n301 VTAIL.n300 171.744
R323 VTAIL.n300 VTAIL.n246 171.744
R324 VTAIL.n293 VTAIL.n246 171.744
R325 VTAIL.n293 VTAIL.n292 171.744
R326 VTAIL.n292 VTAIL.n250 171.744
R327 VTAIL.n285 VTAIL.n250 171.744
R328 VTAIL.n285 VTAIL.n284 171.744
R329 VTAIL.n284 VTAIL.n254 171.744
R330 VTAIL.n277 VTAIL.n254 171.744
R331 VTAIL.n277 VTAIL.n276 171.744
R332 VTAIL.n276 VTAIL.n258 171.744
R333 VTAIL.n269 VTAIL.n258 171.744
R334 VTAIL.n269 VTAIL.n268 171.744
R335 VTAIL.n268 VTAIL.n262 171.744
R336 VTAIL.t9 VTAIL.n577 85.8723
R337 VTAIL.t15 VTAIL.n25 85.8723
R338 VTAIL.t4 VTAIL.n103 85.8723
R339 VTAIL.t1 VTAIL.n183 85.8723
R340 VTAIL.t5 VTAIL.n500 85.8723
R341 VTAIL.t6 VTAIL.n420 85.8723
R342 VTAIL.t13 VTAIL.n342 85.8723
R343 VTAIL.t10 VTAIL.n262 85.8723
R344 VTAIL.n475 VTAIL.n474 58.5343
R345 VTAIL.n317 VTAIL.n316 58.5343
R346 VTAIL.n1 VTAIL.n0 58.5341
R347 VTAIL.n159 VTAIL.n158 58.5341
R348 VTAIL.n631 VTAIL.n630 36.0641
R349 VTAIL.n79 VTAIL.n78 36.0641
R350 VTAIL.n157 VTAIL.n156 36.0641
R351 VTAIL.n237 VTAIL.n236 36.0641
R352 VTAIL.n553 VTAIL.n552 36.0641
R353 VTAIL.n473 VTAIL.n472 36.0641
R354 VTAIL.n395 VTAIL.n394 36.0641
R355 VTAIL.n315 VTAIL.n314 36.0641
R356 VTAIL.n631 VTAIL.n553 25.1686
R357 VTAIL.n315 VTAIL.n237 25.1686
R358 VTAIL.n579 VTAIL.n578 16.3895
R359 VTAIL.n27 VTAIL.n26 16.3895
R360 VTAIL.n105 VTAIL.n104 16.3895
R361 VTAIL.n185 VTAIL.n184 16.3895
R362 VTAIL.n502 VTAIL.n501 16.3895
R363 VTAIL.n422 VTAIL.n421 16.3895
R364 VTAIL.n344 VTAIL.n343 16.3895
R365 VTAIL.n264 VTAIL.n263 16.3895
R366 VTAIL.n627 VTAIL.n556 13.1884
R367 VTAIL.n75 VTAIL.n4 13.1884
R368 VTAIL.n153 VTAIL.n82 13.1884
R369 VTAIL.n233 VTAIL.n162 13.1884
R370 VTAIL.n549 VTAIL.n478 13.1884
R371 VTAIL.n469 VTAIL.n398 13.1884
R372 VTAIL.n391 VTAIL.n320 13.1884
R373 VTAIL.n311 VTAIL.n240 13.1884
R374 VTAIL.n582 VTAIL.n581 12.8005
R375 VTAIL.n623 VTAIL.n622 12.8005
R376 VTAIL.n628 VTAIL.n554 12.8005
R377 VTAIL.n30 VTAIL.n29 12.8005
R378 VTAIL.n71 VTAIL.n70 12.8005
R379 VTAIL.n76 VTAIL.n2 12.8005
R380 VTAIL.n108 VTAIL.n107 12.8005
R381 VTAIL.n149 VTAIL.n148 12.8005
R382 VTAIL.n154 VTAIL.n80 12.8005
R383 VTAIL.n188 VTAIL.n187 12.8005
R384 VTAIL.n229 VTAIL.n228 12.8005
R385 VTAIL.n234 VTAIL.n160 12.8005
R386 VTAIL.n550 VTAIL.n476 12.8005
R387 VTAIL.n545 VTAIL.n480 12.8005
R388 VTAIL.n505 VTAIL.n504 12.8005
R389 VTAIL.n470 VTAIL.n396 12.8005
R390 VTAIL.n465 VTAIL.n400 12.8005
R391 VTAIL.n425 VTAIL.n424 12.8005
R392 VTAIL.n392 VTAIL.n318 12.8005
R393 VTAIL.n387 VTAIL.n322 12.8005
R394 VTAIL.n347 VTAIL.n346 12.8005
R395 VTAIL.n312 VTAIL.n238 12.8005
R396 VTAIL.n307 VTAIL.n242 12.8005
R397 VTAIL.n267 VTAIL.n266 12.8005
R398 VTAIL.n585 VTAIL.n576 12.0247
R399 VTAIL.n621 VTAIL.n558 12.0247
R400 VTAIL.n33 VTAIL.n24 12.0247
R401 VTAIL.n69 VTAIL.n6 12.0247
R402 VTAIL.n111 VTAIL.n102 12.0247
R403 VTAIL.n147 VTAIL.n84 12.0247
R404 VTAIL.n191 VTAIL.n182 12.0247
R405 VTAIL.n227 VTAIL.n164 12.0247
R406 VTAIL.n544 VTAIL.n481 12.0247
R407 VTAIL.n508 VTAIL.n499 12.0247
R408 VTAIL.n464 VTAIL.n401 12.0247
R409 VTAIL.n428 VTAIL.n419 12.0247
R410 VTAIL.n386 VTAIL.n323 12.0247
R411 VTAIL.n350 VTAIL.n341 12.0247
R412 VTAIL.n306 VTAIL.n243 12.0247
R413 VTAIL.n270 VTAIL.n261 12.0247
R414 VTAIL.n586 VTAIL.n574 11.249
R415 VTAIL.n618 VTAIL.n617 11.249
R416 VTAIL.n34 VTAIL.n22 11.249
R417 VTAIL.n66 VTAIL.n65 11.249
R418 VTAIL.n112 VTAIL.n100 11.249
R419 VTAIL.n144 VTAIL.n143 11.249
R420 VTAIL.n192 VTAIL.n180 11.249
R421 VTAIL.n224 VTAIL.n223 11.249
R422 VTAIL.n541 VTAIL.n540 11.249
R423 VTAIL.n509 VTAIL.n497 11.249
R424 VTAIL.n461 VTAIL.n460 11.249
R425 VTAIL.n429 VTAIL.n417 11.249
R426 VTAIL.n383 VTAIL.n382 11.249
R427 VTAIL.n351 VTAIL.n339 11.249
R428 VTAIL.n303 VTAIL.n302 11.249
R429 VTAIL.n271 VTAIL.n259 11.249
R430 VTAIL.n590 VTAIL.n589 10.4732
R431 VTAIL.n614 VTAIL.n560 10.4732
R432 VTAIL.n38 VTAIL.n37 10.4732
R433 VTAIL.n62 VTAIL.n8 10.4732
R434 VTAIL.n116 VTAIL.n115 10.4732
R435 VTAIL.n140 VTAIL.n86 10.4732
R436 VTAIL.n196 VTAIL.n195 10.4732
R437 VTAIL.n220 VTAIL.n166 10.4732
R438 VTAIL.n537 VTAIL.n483 10.4732
R439 VTAIL.n513 VTAIL.n512 10.4732
R440 VTAIL.n457 VTAIL.n403 10.4732
R441 VTAIL.n433 VTAIL.n432 10.4732
R442 VTAIL.n379 VTAIL.n325 10.4732
R443 VTAIL.n355 VTAIL.n354 10.4732
R444 VTAIL.n299 VTAIL.n245 10.4732
R445 VTAIL.n275 VTAIL.n274 10.4732
R446 VTAIL.n593 VTAIL.n572 9.69747
R447 VTAIL.n613 VTAIL.n562 9.69747
R448 VTAIL.n41 VTAIL.n20 9.69747
R449 VTAIL.n61 VTAIL.n10 9.69747
R450 VTAIL.n119 VTAIL.n98 9.69747
R451 VTAIL.n139 VTAIL.n88 9.69747
R452 VTAIL.n199 VTAIL.n178 9.69747
R453 VTAIL.n219 VTAIL.n168 9.69747
R454 VTAIL.n536 VTAIL.n485 9.69747
R455 VTAIL.n516 VTAIL.n495 9.69747
R456 VTAIL.n456 VTAIL.n405 9.69747
R457 VTAIL.n436 VTAIL.n415 9.69747
R458 VTAIL.n378 VTAIL.n327 9.69747
R459 VTAIL.n358 VTAIL.n337 9.69747
R460 VTAIL.n298 VTAIL.n247 9.69747
R461 VTAIL.n278 VTAIL.n257 9.69747
R462 VTAIL.n630 VTAIL.n629 9.45567
R463 VTAIL.n78 VTAIL.n77 9.45567
R464 VTAIL.n156 VTAIL.n155 9.45567
R465 VTAIL.n236 VTAIL.n235 9.45567
R466 VTAIL.n552 VTAIL.n551 9.45567
R467 VTAIL.n472 VTAIL.n471 9.45567
R468 VTAIL.n394 VTAIL.n393 9.45567
R469 VTAIL.n314 VTAIL.n313 9.45567
R470 VTAIL.n629 VTAIL.n628 9.3005
R471 VTAIL.n568 VTAIL.n567 9.3005
R472 VTAIL.n597 VTAIL.n596 9.3005
R473 VTAIL.n595 VTAIL.n594 9.3005
R474 VTAIL.n572 VTAIL.n571 9.3005
R475 VTAIL.n589 VTAIL.n588 9.3005
R476 VTAIL.n587 VTAIL.n586 9.3005
R477 VTAIL.n576 VTAIL.n575 9.3005
R478 VTAIL.n581 VTAIL.n580 9.3005
R479 VTAIL.n603 VTAIL.n602 9.3005
R480 VTAIL.n605 VTAIL.n604 9.3005
R481 VTAIL.n564 VTAIL.n563 9.3005
R482 VTAIL.n611 VTAIL.n610 9.3005
R483 VTAIL.n613 VTAIL.n612 9.3005
R484 VTAIL.n560 VTAIL.n559 9.3005
R485 VTAIL.n619 VTAIL.n618 9.3005
R486 VTAIL.n621 VTAIL.n620 9.3005
R487 VTAIL.n622 VTAIL.n555 9.3005
R488 VTAIL.n77 VTAIL.n76 9.3005
R489 VTAIL.n16 VTAIL.n15 9.3005
R490 VTAIL.n45 VTAIL.n44 9.3005
R491 VTAIL.n43 VTAIL.n42 9.3005
R492 VTAIL.n20 VTAIL.n19 9.3005
R493 VTAIL.n37 VTAIL.n36 9.3005
R494 VTAIL.n35 VTAIL.n34 9.3005
R495 VTAIL.n24 VTAIL.n23 9.3005
R496 VTAIL.n29 VTAIL.n28 9.3005
R497 VTAIL.n51 VTAIL.n50 9.3005
R498 VTAIL.n53 VTAIL.n52 9.3005
R499 VTAIL.n12 VTAIL.n11 9.3005
R500 VTAIL.n59 VTAIL.n58 9.3005
R501 VTAIL.n61 VTAIL.n60 9.3005
R502 VTAIL.n8 VTAIL.n7 9.3005
R503 VTAIL.n67 VTAIL.n66 9.3005
R504 VTAIL.n69 VTAIL.n68 9.3005
R505 VTAIL.n70 VTAIL.n3 9.3005
R506 VTAIL.n155 VTAIL.n154 9.3005
R507 VTAIL.n94 VTAIL.n93 9.3005
R508 VTAIL.n123 VTAIL.n122 9.3005
R509 VTAIL.n121 VTAIL.n120 9.3005
R510 VTAIL.n98 VTAIL.n97 9.3005
R511 VTAIL.n115 VTAIL.n114 9.3005
R512 VTAIL.n113 VTAIL.n112 9.3005
R513 VTAIL.n102 VTAIL.n101 9.3005
R514 VTAIL.n107 VTAIL.n106 9.3005
R515 VTAIL.n129 VTAIL.n128 9.3005
R516 VTAIL.n131 VTAIL.n130 9.3005
R517 VTAIL.n90 VTAIL.n89 9.3005
R518 VTAIL.n137 VTAIL.n136 9.3005
R519 VTAIL.n139 VTAIL.n138 9.3005
R520 VTAIL.n86 VTAIL.n85 9.3005
R521 VTAIL.n145 VTAIL.n144 9.3005
R522 VTAIL.n147 VTAIL.n146 9.3005
R523 VTAIL.n148 VTAIL.n81 9.3005
R524 VTAIL.n235 VTAIL.n234 9.3005
R525 VTAIL.n174 VTAIL.n173 9.3005
R526 VTAIL.n203 VTAIL.n202 9.3005
R527 VTAIL.n201 VTAIL.n200 9.3005
R528 VTAIL.n178 VTAIL.n177 9.3005
R529 VTAIL.n195 VTAIL.n194 9.3005
R530 VTAIL.n193 VTAIL.n192 9.3005
R531 VTAIL.n182 VTAIL.n181 9.3005
R532 VTAIL.n187 VTAIL.n186 9.3005
R533 VTAIL.n209 VTAIL.n208 9.3005
R534 VTAIL.n211 VTAIL.n210 9.3005
R535 VTAIL.n170 VTAIL.n169 9.3005
R536 VTAIL.n217 VTAIL.n216 9.3005
R537 VTAIL.n219 VTAIL.n218 9.3005
R538 VTAIL.n166 VTAIL.n165 9.3005
R539 VTAIL.n225 VTAIL.n224 9.3005
R540 VTAIL.n227 VTAIL.n226 9.3005
R541 VTAIL.n228 VTAIL.n161 9.3005
R542 VTAIL.n528 VTAIL.n527 9.3005
R543 VTAIL.n487 VTAIL.n486 9.3005
R544 VTAIL.n534 VTAIL.n533 9.3005
R545 VTAIL.n536 VTAIL.n535 9.3005
R546 VTAIL.n483 VTAIL.n482 9.3005
R547 VTAIL.n542 VTAIL.n541 9.3005
R548 VTAIL.n544 VTAIL.n543 9.3005
R549 VTAIL.n480 VTAIL.n477 9.3005
R550 VTAIL.n551 VTAIL.n550 9.3005
R551 VTAIL.n526 VTAIL.n525 9.3005
R552 VTAIL.n491 VTAIL.n490 9.3005
R553 VTAIL.n520 VTAIL.n519 9.3005
R554 VTAIL.n518 VTAIL.n517 9.3005
R555 VTAIL.n495 VTAIL.n494 9.3005
R556 VTAIL.n512 VTAIL.n511 9.3005
R557 VTAIL.n510 VTAIL.n509 9.3005
R558 VTAIL.n499 VTAIL.n498 9.3005
R559 VTAIL.n504 VTAIL.n503 9.3005
R560 VTAIL.n448 VTAIL.n447 9.3005
R561 VTAIL.n407 VTAIL.n406 9.3005
R562 VTAIL.n454 VTAIL.n453 9.3005
R563 VTAIL.n456 VTAIL.n455 9.3005
R564 VTAIL.n403 VTAIL.n402 9.3005
R565 VTAIL.n462 VTAIL.n461 9.3005
R566 VTAIL.n464 VTAIL.n463 9.3005
R567 VTAIL.n400 VTAIL.n397 9.3005
R568 VTAIL.n471 VTAIL.n470 9.3005
R569 VTAIL.n446 VTAIL.n445 9.3005
R570 VTAIL.n411 VTAIL.n410 9.3005
R571 VTAIL.n440 VTAIL.n439 9.3005
R572 VTAIL.n438 VTAIL.n437 9.3005
R573 VTAIL.n415 VTAIL.n414 9.3005
R574 VTAIL.n432 VTAIL.n431 9.3005
R575 VTAIL.n430 VTAIL.n429 9.3005
R576 VTAIL.n419 VTAIL.n418 9.3005
R577 VTAIL.n424 VTAIL.n423 9.3005
R578 VTAIL.n370 VTAIL.n369 9.3005
R579 VTAIL.n329 VTAIL.n328 9.3005
R580 VTAIL.n376 VTAIL.n375 9.3005
R581 VTAIL.n378 VTAIL.n377 9.3005
R582 VTAIL.n325 VTAIL.n324 9.3005
R583 VTAIL.n384 VTAIL.n383 9.3005
R584 VTAIL.n386 VTAIL.n385 9.3005
R585 VTAIL.n322 VTAIL.n319 9.3005
R586 VTAIL.n393 VTAIL.n392 9.3005
R587 VTAIL.n368 VTAIL.n367 9.3005
R588 VTAIL.n333 VTAIL.n332 9.3005
R589 VTAIL.n362 VTAIL.n361 9.3005
R590 VTAIL.n360 VTAIL.n359 9.3005
R591 VTAIL.n337 VTAIL.n336 9.3005
R592 VTAIL.n354 VTAIL.n353 9.3005
R593 VTAIL.n352 VTAIL.n351 9.3005
R594 VTAIL.n341 VTAIL.n340 9.3005
R595 VTAIL.n346 VTAIL.n345 9.3005
R596 VTAIL.n290 VTAIL.n289 9.3005
R597 VTAIL.n249 VTAIL.n248 9.3005
R598 VTAIL.n296 VTAIL.n295 9.3005
R599 VTAIL.n298 VTAIL.n297 9.3005
R600 VTAIL.n245 VTAIL.n244 9.3005
R601 VTAIL.n304 VTAIL.n303 9.3005
R602 VTAIL.n306 VTAIL.n305 9.3005
R603 VTAIL.n242 VTAIL.n239 9.3005
R604 VTAIL.n313 VTAIL.n312 9.3005
R605 VTAIL.n288 VTAIL.n287 9.3005
R606 VTAIL.n253 VTAIL.n252 9.3005
R607 VTAIL.n282 VTAIL.n281 9.3005
R608 VTAIL.n280 VTAIL.n279 9.3005
R609 VTAIL.n257 VTAIL.n256 9.3005
R610 VTAIL.n274 VTAIL.n273 9.3005
R611 VTAIL.n272 VTAIL.n271 9.3005
R612 VTAIL.n261 VTAIL.n260 9.3005
R613 VTAIL.n266 VTAIL.n265 9.3005
R614 VTAIL.n594 VTAIL.n570 8.92171
R615 VTAIL.n610 VTAIL.n609 8.92171
R616 VTAIL.n42 VTAIL.n18 8.92171
R617 VTAIL.n58 VTAIL.n57 8.92171
R618 VTAIL.n120 VTAIL.n96 8.92171
R619 VTAIL.n136 VTAIL.n135 8.92171
R620 VTAIL.n200 VTAIL.n176 8.92171
R621 VTAIL.n216 VTAIL.n215 8.92171
R622 VTAIL.n533 VTAIL.n532 8.92171
R623 VTAIL.n517 VTAIL.n493 8.92171
R624 VTAIL.n453 VTAIL.n452 8.92171
R625 VTAIL.n437 VTAIL.n413 8.92171
R626 VTAIL.n375 VTAIL.n374 8.92171
R627 VTAIL.n359 VTAIL.n335 8.92171
R628 VTAIL.n295 VTAIL.n294 8.92171
R629 VTAIL.n279 VTAIL.n255 8.92171
R630 VTAIL.n598 VTAIL.n597 8.14595
R631 VTAIL.n606 VTAIL.n564 8.14595
R632 VTAIL.n46 VTAIL.n45 8.14595
R633 VTAIL.n54 VTAIL.n12 8.14595
R634 VTAIL.n124 VTAIL.n123 8.14595
R635 VTAIL.n132 VTAIL.n90 8.14595
R636 VTAIL.n204 VTAIL.n203 8.14595
R637 VTAIL.n212 VTAIL.n170 8.14595
R638 VTAIL.n529 VTAIL.n487 8.14595
R639 VTAIL.n521 VTAIL.n520 8.14595
R640 VTAIL.n449 VTAIL.n407 8.14595
R641 VTAIL.n441 VTAIL.n440 8.14595
R642 VTAIL.n371 VTAIL.n329 8.14595
R643 VTAIL.n363 VTAIL.n362 8.14595
R644 VTAIL.n291 VTAIL.n249 8.14595
R645 VTAIL.n283 VTAIL.n282 8.14595
R646 VTAIL.n601 VTAIL.n568 7.3702
R647 VTAIL.n605 VTAIL.n566 7.3702
R648 VTAIL.n49 VTAIL.n16 7.3702
R649 VTAIL.n53 VTAIL.n14 7.3702
R650 VTAIL.n127 VTAIL.n94 7.3702
R651 VTAIL.n131 VTAIL.n92 7.3702
R652 VTAIL.n207 VTAIL.n174 7.3702
R653 VTAIL.n211 VTAIL.n172 7.3702
R654 VTAIL.n528 VTAIL.n489 7.3702
R655 VTAIL.n524 VTAIL.n491 7.3702
R656 VTAIL.n448 VTAIL.n409 7.3702
R657 VTAIL.n444 VTAIL.n411 7.3702
R658 VTAIL.n370 VTAIL.n331 7.3702
R659 VTAIL.n366 VTAIL.n333 7.3702
R660 VTAIL.n290 VTAIL.n251 7.3702
R661 VTAIL.n286 VTAIL.n253 7.3702
R662 VTAIL.n602 VTAIL.n601 6.59444
R663 VTAIL.n602 VTAIL.n566 6.59444
R664 VTAIL.n50 VTAIL.n49 6.59444
R665 VTAIL.n50 VTAIL.n14 6.59444
R666 VTAIL.n128 VTAIL.n127 6.59444
R667 VTAIL.n128 VTAIL.n92 6.59444
R668 VTAIL.n208 VTAIL.n207 6.59444
R669 VTAIL.n208 VTAIL.n172 6.59444
R670 VTAIL.n525 VTAIL.n489 6.59444
R671 VTAIL.n525 VTAIL.n524 6.59444
R672 VTAIL.n445 VTAIL.n409 6.59444
R673 VTAIL.n445 VTAIL.n444 6.59444
R674 VTAIL.n367 VTAIL.n331 6.59444
R675 VTAIL.n367 VTAIL.n366 6.59444
R676 VTAIL.n287 VTAIL.n251 6.59444
R677 VTAIL.n287 VTAIL.n286 6.59444
R678 VTAIL.n598 VTAIL.n568 5.81868
R679 VTAIL.n606 VTAIL.n605 5.81868
R680 VTAIL.n46 VTAIL.n16 5.81868
R681 VTAIL.n54 VTAIL.n53 5.81868
R682 VTAIL.n124 VTAIL.n94 5.81868
R683 VTAIL.n132 VTAIL.n131 5.81868
R684 VTAIL.n204 VTAIL.n174 5.81868
R685 VTAIL.n212 VTAIL.n211 5.81868
R686 VTAIL.n529 VTAIL.n528 5.81868
R687 VTAIL.n521 VTAIL.n491 5.81868
R688 VTAIL.n449 VTAIL.n448 5.81868
R689 VTAIL.n441 VTAIL.n411 5.81868
R690 VTAIL.n371 VTAIL.n370 5.81868
R691 VTAIL.n363 VTAIL.n333 5.81868
R692 VTAIL.n291 VTAIL.n290 5.81868
R693 VTAIL.n283 VTAIL.n253 5.81868
R694 VTAIL.n597 VTAIL.n570 5.04292
R695 VTAIL.n609 VTAIL.n564 5.04292
R696 VTAIL.n45 VTAIL.n18 5.04292
R697 VTAIL.n57 VTAIL.n12 5.04292
R698 VTAIL.n123 VTAIL.n96 5.04292
R699 VTAIL.n135 VTAIL.n90 5.04292
R700 VTAIL.n203 VTAIL.n176 5.04292
R701 VTAIL.n215 VTAIL.n170 5.04292
R702 VTAIL.n532 VTAIL.n487 5.04292
R703 VTAIL.n520 VTAIL.n493 5.04292
R704 VTAIL.n452 VTAIL.n407 5.04292
R705 VTAIL.n440 VTAIL.n413 5.04292
R706 VTAIL.n374 VTAIL.n329 5.04292
R707 VTAIL.n362 VTAIL.n335 5.04292
R708 VTAIL.n294 VTAIL.n249 5.04292
R709 VTAIL.n282 VTAIL.n255 5.04292
R710 VTAIL.n594 VTAIL.n593 4.26717
R711 VTAIL.n610 VTAIL.n562 4.26717
R712 VTAIL.n42 VTAIL.n41 4.26717
R713 VTAIL.n58 VTAIL.n10 4.26717
R714 VTAIL.n120 VTAIL.n119 4.26717
R715 VTAIL.n136 VTAIL.n88 4.26717
R716 VTAIL.n200 VTAIL.n199 4.26717
R717 VTAIL.n216 VTAIL.n168 4.26717
R718 VTAIL.n533 VTAIL.n485 4.26717
R719 VTAIL.n517 VTAIL.n516 4.26717
R720 VTAIL.n453 VTAIL.n405 4.26717
R721 VTAIL.n437 VTAIL.n436 4.26717
R722 VTAIL.n375 VTAIL.n327 4.26717
R723 VTAIL.n359 VTAIL.n358 4.26717
R724 VTAIL.n295 VTAIL.n247 4.26717
R725 VTAIL.n279 VTAIL.n278 4.26717
R726 VTAIL.n580 VTAIL.n579 3.70982
R727 VTAIL.n28 VTAIL.n27 3.70982
R728 VTAIL.n106 VTAIL.n105 3.70982
R729 VTAIL.n186 VTAIL.n185 3.70982
R730 VTAIL.n503 VTAIL.n502 3.70982
R731 VTAIL.n423 VTAIL.n422 3.70982
R732 VTAIL.n345 VTAIL.n344 3.70982
R733 VTAIL.n265 VTAIL.n264 3.70982
R734 VTAIL.n590 VTAIL.n572 3.49141
R735 VTAIL.n614 VTAIL.n613 3.49141
R736 VTAIL.n38 VTAIL.n20 3.49141
R737 VTAIL.n62 VTAIL.n61 3.49141
R738 VTAIL.n116 VTAIL.n98 3.49141
R739 VTAIL.n140 VTAIL.n139 3.49141
R740 VTAIL.n196 VTAIL.n178 3.49141
R741 VTAIL.n220 VTAIL.n219 3.49141
R742 VTAIL.n537 VTAIL.n536 3.49141
R743 VTAIL.n513 VTAIL.n495 3.49141
R744 VTAIL.n457 VTAIL.n456 3.49141
R745 VTAIL.n433 VTAIL.n415 3.49141
R746 VTAIL.n379 VTAIL.n378 3.49141
R747 VTAIL.n355 VTAIL.n337 3.49141
R748 VTAIL.n299 VTAIL.n298 3.49141
R749 VTAIL.n275 VTAIL.n257 3.49141
R750 VTAIL.n589 VTAIL.n574 2.71565
R751 VTAIL.n617 VTAIL.n560 2.71565
R752 VTAIL.n37 VTAIL.n22 2.71565
R753 VTAIL.n65 VTAIL.n8 2.71565
R754 VTAIL.n115 VTAIL.n100 2.71565
R755 VTAIL.n143 VTAIL.n86 2.71565
R756 VTAIL.n195 VTAIL.n180 2.71565
R757 VTAIL.n223 VTAIL.n166 2.71565
R758 VTAIL.n540 VTAIL.n483 2.71565
R759 VTAIL.n512 VTAIL.n497 2.71565
R760 VTAIL.n460 VTAIL.n403 2.71565
R761 VTAIL.n432 VTAIL.n417 2.71565
R762 VTAIL.n382 VTAIL.n325 2.71565
R763 VTAIL.n354 VTAIL.n339 2.71565
R764 VTAIL.n302 VTAIL.n245 2.71565
R765 VTAIL.n274 VTAIL.n259 2.71565
R766 VTAIL.n0 VTAIL.t12 2.30255
R767 VTAIL.n0 VTAIL.t11 2.30255
R768 VTAIL.n158 VTAIL.t3 2.30255
R769 VTAIL.n158 VTAIL.t0 2.30255
R770 VTAIL.n474 VTAIL.t7 2.30255
R771 VTAIL.n474 VTAIL.t2 2.30255
R772 VTAIL.n316 VTAIL.t8 2.30255
R773 VTAIL.n316 VTAIL.t14 2.30255
R774 VTAIL.n586 VTAIL.n585 1.93989
R775 VTAIL.n618 VTAIL.n558 1.93989
R776 VTAIL.n34 VTAIL.n33 1.93989
R777 VTAIL.n66 VTAIL.n6 1.93989
R778 VTAIL.n112 VTAIL.n111 1.93989
R779 VTAIL.n144 VTAIL.n84 1.93989
R780 VTAIL.n192 VTAIL.n191 1.93989
R781 VTAIL.n224 VTAIL.n164 1.93989
R782 VTAIL.n541 VTAIL.n481 1.93989
R783 VTAIL.n509 VTAIL.n508 1.93989
R784 VTAIL.n461 VTAIL.n401 1.93989
R785 VTAIL.n429 VTAIL.n428 1.93989
R786 VTAIL.n383 VTAIL.n323 1.93989
R787 VTAIL.n351 VTAIL.n350 1.93989
R788 VTAIL.n303 VTAIL.n243 1.93989
R789 VTAIL.n271 VTAIL.n270 1.93989
R790 VTAIL.n582 VTAIL.n576 1.16414
R791 VTAIL.n623 VTAIL.n621 1.16414
R792 VTAIL.n630 VTAIL.n554 1.16414
R793 VTAIL.n30 VTAIL.n24 1.16414
R794 VTAIL.n71 VTAIL.n69 1.16414
R795 VTAIL.n78 VTAIL.n2 1.16414
R796 VTAIL.n108 VTAIL.n102 1.16414
R797 VTAIL.n149 VTAIL.n147 1.16414
R798 VTAIL.n156 VTAIL.n80 1.16414
R799 VTAIL.n188 VTAIL.n182 1.16414
R800 VTAIL.n229 VTAIL.n227 1.16414
R801 VTAIL.n236 VTAIL.n160 1.16414
R802 VTAIL.n552 VTAIL.n476 1.16414
R803 VTAIL.n545 VTAIL.n544 1.16414
R804 VTAIL.n505 VTAIL.n499 1.16414
R805 VTAIL.n472 VTAIL.n396 1.16414
R806 VTAIL.n465 VTAIL.n464 1.16414
R807 VTAIL.n425 VTAIL.n419 1.16414
R808 VTAIL.n394 VTAIL.n318 1.16414
R809 VTAIL.n387 VTAIL.n386 1.16414
R810 VTAIL.n347 VTAIL.n341 1.16414
R811 VTAIL.n314 VTAIL.n238 1.16414
R812 VTAIL.n307 VTAIL.n306 1.16414
R813 VTAIL.n267 VTAIL.n261 1.16414
R814 VTAIL.n317 VTAIL.n315 0.62981
R815 VTAIL.n395 VTAIL.n317 0.62981
R816 VTAIL.n475 VTAIL.n473 0.62981
R817 VTAIL.n553 VTAIL.n475 0.62981
R818 VTAIL.n237 VTAIL.n159 0.62981
R819 VTAIL.n159 VTAIL.n157 0.62981
R820 VTAIL.n79 VTAIL.n1 0.62981
R821 VTAIL VTAIL.n631 0.571621
R822 VTAIL.n473 VTAIL.n395 0.470328
R823 VTAIL.n157 VTAIL.n79 0.470328
R824 VTAIL.n581 VTAIL.n578 0.388379
R825 VTAIL.n622 VTAIL.n556 0.388379
R826 VTAIL.n628 VTAIL.n627 0.388379
R827 VTAIL.n29 VTAIL.n26 0.388379
R828 VTAIL.n70 VTAIL.n4 0.388379
R829 VTAIL.n76 VTAIL.n75 0.388379
R830 VTAIL.n107 VTAIL.n104 0.388379
R831 VTAIL.n148 VTAIL.n82 0.388379
R832 VTAIL.n154 VTAIL.n153 0.388379
R833 VTAIL.n187 VTAIL.n184 0.388379
R834 VTAIL.n228 VTAIL.n162 0.388379
R835 VTAIL.n234 VTAIL.n233 0.388379
R836 VTAIL.n550 VTAIL.n549 0.388379
R837 VTAIL.n480 VTAIL.n478 0.388379
R838 VTAIL.n504 VTAIL.n501 0.388379
R839 VTAIL.n470 VTAIL.n469 0.388379
R840 VTAIL.n400 VTAIL.n398 0.388379
R841 VTAIL.n424 VTAIL.n421 0.388379
R842 VTAIL.n392 VTAIL.n391 0.388379
R843 VTAIL.n322 VTAIL.n320 0.388379
R844 VTAIL.n346 VTAIL.n343 0.388379
R845 VTAIL.n312 VTAIL.n311 0.388379
R846 VTAIL.n242 VTAIL.n240 0.388379
R847 VTAIL.n266 VTAIL.n263 0.388379
R848 VTAIL.n580 VTAIL.n575 0.155672
R849 VTAIL.n587 VTAIL.n575 0.155672
R850 VTAIL.n588 VTAIL.n587 0.155672
R851 VTAIL.n588 VTAIL.n571 0.155672
R852 VTAIL.n595 VTAIL.n571 0.155672
R853 VTAIL.n596 VTAIL.n595 0.155672
R854 VTAIL.n596 VTAIL.n567 0.155672
R855 VTAIL.n603 VTAIL.n567 0.155672
R856 VTAIL.n604 VTAIL.n603 0.155672
R857 VTAIL.n604 VTAIL.n563 0.155672
R858 VTAIL.n611 VTAIL.n563 0.155672
R859 VTAIL.n612 VTAIL.n611 0.155672
R860 VTAIL.n612 VTAIL.n559 0.155672
R861 VTAIL.n619 VTAIL.n559 0.155672
R862 VTAIL.n620 VTAIL.n619 0.155672
R863 VTAIL.n620 VTAIL.n555 0.155672
R864 VTAIL.n629 VTAIL.n555 0.155672
R865 VTAIL.n28 VTAIL.n23 0.155672
R866 VTAIL.n35 VTAIL.n23 0.155672
R867 VTAIL.n36 VTAIL.n35 0.155672
R868 VTAIL.n36 VTAIL.n19 0.155672
R869 VTAIL.n43 VTAIL.n19 0.155672
R870 VTAIL.n44 VTAIL.n43 0.155672
R871 VTAIL.n44 VTAIL.n15 0.155672
R872 VTAIL.n51 VTAIL.n15 0.155672
R873 VTAIL.n52 VTAIL.n51 0.155672
R874 VTAIL.n52 VTAIL.n11 0.155672
R875 VTAIL.n59 VTAIL.n11 0.155672
R876 VTAIL.n60 VTAIL.n59 0.155672
R877 VTAIL.n60 VTAIL.n7 0.155672
R878 VTAIL.n67 VTAIL.n7 0.155672
R879 VTAIL.n68 VTAIL.n67 0.155672
R880 VTAIL.n68 VTAIL.n3 0.155672
R881 VTAIL.n77 VTAIL.n3 0.155672
R882 VTAIL.n106 VTAIL.n101 0.155672
R883 VTAIL.n113 VTAIL.n101 0.155672
R884 VTAIL.n114 VTAIL.n113 0.155672
R885 VTAIL.n114 VTAIL.n97 0.155672
R886 VTAIL.n121 VTAIL.n97 0.155672
R887 VTAIL.n122 VTAIL.n121 0.155672
R888 VTAIL.n122 VTAIL.n93 0.155672
R889 VTAIL.n129 VTAIL.n93 0.155672
R890 VTAIL.n130 VTAIL.n129 0.155672
R891 VTAIL.n130 VTAIL.n89 0.155672
R892 VTAIL.n137 VTAIL.n89 0.155672
R893 VTAIL.n138 VTAIL.n137 0.155672
R894 VTAIL.n138 VTAIL.n85 0.155672
R895 VTAIL.n145 VTAIL.n85 0.155672
R896 VTAIL.n146 VTAIL.n145 0.155672
R897 VTAIL.n146 VTAIL.n81 0.155672
R898 VTAIL.n155 VTAIL.n81 0.155672
R899 VTAIL.n186 VTAIL.n181 0.155672
R900 VTAIL.n193 VTAIL.n181 0.155672
R901 VTAIL.n194 VTAIL.n193 0.155672
R902 VTAIL.n194 VTAIL.n177 0.155672
R903 VTAIL.n201 VTAIL.n177 0.155672
R904 VTAIL.n202 VTAIL.n201 0.155672
R905 VTAIL.n202 VTAIL.n173 0.155672
R906 VTAIL.n209 VTAIL.n173 0.155672
R907 VTAIL.n210 VTAIL.n209 0.155672
R908 VTAIL.n210 VTAIL.n169 0.155672
R909 VTAIL.n217 VTAIL.n169 0.155672
R910 VTAIL.n218 VTAIL.n217 0.155672
R911 VTAIL.n218 VTAIL.n165 0.155672
R912 VTAIL.n225 VTAIL.n165 0.155672
R913 VTAIL.n226 VTAIL.n225 0.155672
R914 VTAIL.n226 VTAIL.n161 0.155672
R915 VTAIL.n235 VTAIL.n161 0.155672
R916 VTAIL.n551 VTAIL.n477 0.155672
R917 VTAIL.n543 VTAIL.n477 0.155672
R918 VTAIL.n543 VTAIL.n542 0.155672
R919 VTAIL.n542 VTAIL.n482 0.155672
R920 VTAIL.n535 VTAIL.n482 0.155672
R921 VTAIL.n535 VTAIL.n534 0.155672
R922 VTAIL.n534 VTAIL.n486 0.155672
R923 VTAIL.n527 VTAIL.n486 0.155672
R924 VTAIL.n527 VTAIL.n526 0.155672
R925 VTAIL.n526 VTAIL.n490 0.155672
R926 VTAIL.n519 VTAIL.n490 0.155672
R927 VTAIL.n519 VTAIL.n518 0.155672
R928 VTAIL.n518 VTAIL.n494 0.155672
R929 VTAIL.n511 VTAIL.n494 0.155672
R930 VTAIL.n511 VTAIL.n510 0.155672
R931 VTAIL.n510 VTAIL.n498 0.155672
R932 VTAIL.n503 VTAIL.n498 0.155672
R933 VTAIL.n471 VTAIL.n397 0.155672
R934 VTAIL.n463 VTAIL.n397 0.155672
R935 VTAIL.n463 VTAIL.n462 0.155672
R936 VTAIL.n462 VTAIL.n402 0.155672
R937 VTAIL.n455 VTAIL.n402 0.155672
R938 VTAIL.n455 VTAIL.n454 0.155672
R939 VTAIL.n454 VTAIL.n406 0.155672
R940 VTAIL.n447 VTAIL.n406 0.155672
R941 VTAIL.n447 VTAIL.n446 0.155672
R942 VTAIL.n446 VTAIL.n410 0.155672
R943 VTAIL.n439 VTAIL.n410 0.155672
R944 VTAIL.n439 VTAIL.n438 0.155672
R945 VTAIL.n438 VTAIL.n414 0.155672
R946 VTAIL.n431 VTAIL.n414 0.155672
R947 VTAIL.n431 VTAIL.n430 0.155672
R948 VTAIL.n430 VTAIL.n418 0.155672
R949 VTAIL.n423 VTAIL.n418 0.155672
R950 VTAIL.n393 VTAIL.n319 0.155672
R951 VTAIL.n385 VTAIL.n319 0.155672
R952 VTAIL.n385 VTAIL.n384 0.155672
R953 VTAIL.n384 VTAIL.n324 0.155672
R954 VTAIL.n377 VTAIL.n324 0.155672
R955 VTAIL.n377 VTAIL.n376 0.155672
R956 VTAIL.n376 VTAIL.n328 0.155672
R957 VTAIL.n369 VTAIL.n328 0.155672
R958 VTAIL.n369 VTAIL.n368 0.155672
R959 VTAIL.n368 VTAIL.n332 0.155672
R960 VTAIL.n361 VTAIL.n332 0.155672
R961 VTAIL.n361 VTAIL.n360 0.155672
R962 VTAIL.n360 VTAIL.n336 0.155672
R963 VTAIL.n353 VTAIL.n336 0.155672
R964 VTAIL.n353 VTAIL.n352 0.155672
R965 VTAIL.n352 VTAIL.n340 0.155672
R966 VTAIL.n345 VTAIL.n340 0.155672
R967 VTAIL.n313 VTAIL.n239 0.155672
R968 VTAIL.n305 VTAIL.n239 0.155672
R969 VTAIL.n305 VTAIL.n304 0.155672
R970 VTAIL.n304 VTAIL.n244 0.155672
R971 VTAIL.n297 VTAIL.n244 0.155672
R972 VTAIL.n297 VTAIL.n296 0.155672
R973 VTAIL.n296 VTAIL.n248 0.155672
R974 VTAIL.n289 VTAIL.n248 0.155672
R975 VTAIL.n289 VTAIL.n288 0.155672
R976 VTAIL.n288 VTAIL.n252 0.155672
R977 VTAIL.n281 VTAIL.n252 0.155672
R978 VTAIL.n281 VTAIL.n280 0.155672
R979 VTAIL.n280 VTAIL.n256 0.155672
R980 VTAIL.n273 VTAIL.n256 0.155672
R981 VTAIL.n273 VTAIL.n272 0.155672
R982 VTAIL.n272 VTAIL.n260 0.155672
R983 VTAIL.n265 VTAIL.n260 0.155672
R984 VTAIL VTAIL.n1 0.0586897
R985 VDD2.n2 VDD2.n1 75.4722
R986 VDD2.n2 VDD2.n0 75.4722
R987 VDD2 VDD2.n5 75.4694
R988 VDD2.n4 VDD2.n3 75.2131
R989 VDD2.n4 VDD2.n2 38.7196
R990 VDD2.n5 VDD2.t5 2.30255
R991 VDD2.n5 VDD2.t3 2.30255
R992 VDD2.n3 VDD2.t1 2.30255
R993 VDD2.n3 VDD2.t6 2.30255
R994 VDD2.n1 VDD2.t4 2.30255
R995 VDD2.n1 VDD2.t2 2.30255
R996 VDD2.n0 VDD2.t0 2.30255
R997 VDD2.n0 VDD2.t7 2.30255
R998 VDD2 VDD2.n4 0.373345
R999 VP.n3 VP.t4 982.591
R1000 VP.n12 VP.t2 970.116
R1001 VP.n1 VP.t5 970.116
R1002 VP.n6 VP.t7 970.116
R1003 VP.n10 VP.t6 948.938
R1004 VP.n11 VP.t3 948.938
R1005 VP.n5 VP.t0 948.938
R1006 VP.n4 VP.t1 948.938
R1007 VP.n13 VP.n12 161.3
R1008 VP.n5 VP.n2 161.3
R1009 VP.n7 VP.n6 161.3
R1010 VP.n11 VP.n0 161.3
R1011 VP.n10 VP.n9 161.3
R1012 VP.n8 VP.n1 161.3
R1013 VP.n3 VP.n2 74.6542
R1014 VP.n11 VP.n10 48.2005
R1015 VP.n5 VP.n4 48.2005
R1016 VP.n8 VP.n7 42.349
R1017 VP.n10 VP.n1 27.0217
R1018 VP.n12 VP.n11 27.0217
R1019 VP.n6 VP.n5 27.0217
R1020 VP.n4 VP.n3 12.4607
R1021 VP.n7 VP.n2 0.189894
R1022 VP.n9 VP.n8 0.189894
R1023 VP.n9 VP.n0 0.189894
R1024 VP.n13 VP.n0 0.189894
R1025 VP VP.n13 0.0516364
R1026 VDD1 VDD1.n0 75.586
R1027 VDD1.n3 VDD1.n2 75.4722
R1028 VDD1.n3 VDD1.n1 75.4722
R1029 VDD1.n5 VDD1.n4 75.2129
R1030 VDD1.n5 VDD1.n3 39.3026
R1031 VDD1.n4 VDD1.t7 2.30255
R1032 VDD1.n4 VDD1.t0 2.30255
R1033 VDD1.n0 VDD1.t3 2.30255
R1034 VDD1.n0 VDD1.t6 2.30255
R1035 VDD1.n2 VDD1.t4 2.30255
R1036 VDD1.n2 VDD1.t5 2.30255
R1037 VDD1.n1 VDD1.t2 2.30255
R1038 VDD1.n1 VDD1.t1 2.30255
R1039 VDD1 VDD1.n5 0.256966
R1040 B.n112 B.t0 1060.15
R1041 B.n120 B.t9 1060.15
R1042 B.n36 B.t6 1060.15
R1043 B.n42 B.t3 1060.15
R1044 B.n399 B.n68 585
R1045 B.n401 B.n400 585
R1046 B.n402 B.n67 585
R1047 B.n404 B.n403 585
R1048 B.n405 B.n66 585
R1049 B.n407 B.n406 585
R1050 B.n408 B.n65 585
R1051 B.n410 B.n409 585
R1052 B.n411 B.n64 585
R1053 B.n413 B.n412 585
R1054 B.n414 B.n63 585
R1055 B.n416 B.n415 585
R1056 B.n417 B.n62 585
R1057 B.n419 B.n418 585
R1058 B.n420 B.n61 585
R1059 B.n422 B.n421 585
R1060 B.n423 B.n60 585
R1061 B.n425 B.n424 585
R1062 B.n426 B.n59 585
R1063 B.n428 B.n427 585
R1064 B.n429 B.n58 585
R1065 B.n431 B.n430 585
R1066 B.n432 B.n57 585
R1067 B.n434 B.n433 585
R1068 B.n435 B.n56 585
R1069 B.n437 B.n436 585
R1070 B.n438 B.n55 585
R1071 B.n440 B.n439 585
R1072 B.n441 B.n54 585
R1073 B.n443 B.n442 585
R1074 B.n444 B.n53 585
R1075 B.n446 B.n445 585
R1076 B.n447 B.n52 585
R1077 B.n449 B.n448 585
R1078 B.n450 B.n51 585
R1079 B.n452 B.n451 585
R1080 B.n453 B.n50 585
R1081 B.n455 B.n454 585
R1082 B.n456 B.n49 585
R1083 B.n458 B.n457 585
R1084 B.n459 B.n48 585
R1085 B.n461 B.n460 585
R1086 B.n462 B.n47 585
R1087 B.n464 B.n463 585
R1088 B.n465 B.n46 585
R1089 B.n467 B.n466 585
R1090 B.n468 B.n45 585
R1091 B.n470 B.n469 585
R1092 B.n472 B.n471 585
R1093 B.n473 B.n41 585
R1094 B.n475 B.n474 585
R1095 B.n476 B.n40 585
R1096 B.n478 B.n477 585
R1097 B.n479 B.n39 585
R1098 B.n481 B.n480 585
R1099 B.n482 B.n38 585
R1100 B.n484 B.n483 585
R1101 B.n486 B.n35 585
R1102 B.n488 B.n487 585
R1103 B.n489 B.n34 585
R1104 B.n491 B.n490 585
R1105 B.n492 B.n33 585
R1106 B.n494 B.n493 585
R1107 B.n495 B.n32 585
R1108 B.n497 B.n496 585
R1109 B.n498 B.n31 585
R1110 B.n500 B.n499 585
R1111 B.n501 B.n30 585
R1112 B.n503 B.n502 585
R1113 B.n504 B.n29 585
R1114 B.n506 B.n505 585
R1115 B.n507 B.n28 585
R1116 B.n509 B.n508 585
R1117 B.n510 B.n27 585
R1118 B.n512 B.n511 585
R1119 B.n513 B.n26 585
R1120 B.n515 B.n514 585
R1121 B.n516 B.n25 585
R1122 B.n518 B.n517 585
R1123 B.n519 B.n24 585
R1124 B.n521 B.n520 585
R1125 B.n522 B.n23 585
R1126 B.n524 B.n523 585
R1127 B.n525 B.n22 585
R1128 B.n527 B.n526 585
R1129 B.n528 B.n21 585
R1130 B.n530 B.n529 585
R1131 B.n531 B.n20 585
R1132 B.n533 B.n532 585
R1133 B.n534 B.n19 585
R1134 B.n536 B.n535 585
R1135 B.n537 B.n18 585
R1136 B.n539 B.n538 585
R1137 B.n540 B.n17 585
R1138 B.n542 B.n541 585
R1139 B.n543 B.n16 585
R1140 B.n545 B.n544 585
R1141 B.n546 B.n15 585
R1142 B.n548 B.n547 585
R1143 B.n549 B.n14 585
R1144 B.n551 B.n550 585
R1145 B.n552 B.n13 585
R1146 B.n554 B.n553 585
R1147 B.n555 B.n12 585
R1148 B.n557 B.n556 585
R1149 B.n398 B.n397 585
R1150 B.n396 B.n69 585
R1151 B.n395 B.n394 585
R1152 B.n393 B.n70 585
R1153 B.n392 B.n391 585
R1154 B.n390 B.n71 585
R1155 B.n389 B.n388 585
R1156 B.n387 B.n72 585
R1157 B.n386 B.n385 585
R1158 B.n384 B.n73 585
R1159 B.n383 B.n382 585
R1160 B.n381 B.n74 585
R1161 B.n380 B.n379 585
R1162 B.n378 B.n75 585
R1163 B.n377 B.n376 585
R1164 B.n375 B.n76 585
R1165 B.n374 B.n373 585
R1166 B.n372 B.n77 585
R1167 B.n371 B.n370 585
R1168 B.n369 B.n78 585
R1169 B.n368 B.n367 585
R1170 B.n366 B.n79 585
R1171 B.n365 B.n364 585
R1172 B.n363 B.n80 585
R1173 B.n362 B.n361 585
R1174 B.n360 B.n81 585
R1175 B.n359 B.n358 585
R1176 B.n357 B.n82 585
R1177 B.n356 B.n355 585
R1178 B.n354 B.n83 585
R1179 B.n353 B.n352 585
R1180 B.n351 B.n84 585
R1181 B.n350 B.n349 585
R1182 B.n348 B.n85 585
R1183 B.n347 B.n346 585
R1184 B.n345 B.n86 585
R1185 B.n344 B.n343 585
R1186 B.n342 B.n87 585
R1187 B.n341 B.n340 585
R1188 B.n182 B.n181 585
R1189 B.n183 B.n144 585
R1190 B.n185 B.n184 585
R1191 B.n186 B.n143 585
R1192 B.n188 B.n187 585
R1193 B.n189 B.n142 585
R1194 B.n191 B.n190 585
R1195 B.n192 B.n141 585
R1196 B.n194 B.n193 585
R1197 B.n195 B.n140 585
R1198 B.n197 B.n196 585
R1199 B.n198 B.n139 585
R1200 B.n200 B.n199 585
R1201 B.n201 B.n138 585
R1202 B.n203 B.n202 585
R1203 B.n204 B.n137 585
R1204 B.n206 B.n205 585
R1205 B.n207 B.n136 585
R1206 B.n209 B.n208 585
R1207 B.n210 B.n135 585
R1208 B.n212 B.n211 585
R1209 B.n213 B.n134 585
R1210 B.n215 B.n214 585
R1211 B.n216 B.n133 585
R1212 B.n218 B.n217 585
R1213 B.n219 B.n132 585
R1214 B.n221 B.n220 585
R1215 B.n222 B.n131 585
R1216 B.n224 B.n223 585
R1217 B.n225 B.n130 585
R1218 B.n227 B.n226 585
R1219 B.n228 B.n129 585
R1220 B.n230 B.n229 585
R1221 B.n231 B.n128 585
R1222 B.n233 B.n232 585
R1223 B.n234 B.n127 585
R1224 B.n236 B.n235 585
R1225 B.n237 B.n126 585
R1226 B.n239 B.n238 585
R1227 B.n240 B.n125 585
R1228 B.n242 B.n241 585
R1229 B.n243 B.n124 585
R1230 B.n245 B.n244 585
R1231 B.n246 B.n123 585
R1232 B.n248 B.n247 585
R1233 B.n249 B.n122 585
R1234 B.n251 B.n250 585
R1235 B.n252 B.n119 585
R1236 B.n255 B.n254 585
R1237 B.n256 B.n118 585
R1238 B.n258 B.n257 585
R1239 B.n259 B.n117 585
R1240 B.n261 B.n260 585
R1241 B.n262 B.n116 585
R1242 B.n264 B.n263 585
R1243 B.n265 B.n115 585
R1244 B.n267 B.n266 585
R1245 B.n269 B.n268 585
R1246 B.n270 B.n111 585
R1247 B.n272 B.n271 585
R1248 B.n273 B.n110 585
R1249 B.n275 B.n274 585
R1250 B.n276 B.n109 585
R1251 B.n278 B.n277 585
R1252 B.n279 B.n108 585
R1253 B.n281 B.n280 585
R1254 B.n282 B.n107 585
R1255 B.n284 B.n283 585
R1256 B.n285 B.n106 585
R1257 B.n287 B.n286 585
R1258 B.n288 B.n105 585
R1259 B.n290 B.n289 585
R1260 B.n291 B.n104 585
R1261 B.n293 B.n292 585
R1262 B.n294 B.n103 585
R1263 B.n296 B.n295 585
R1264 B.n297 B.n102 585
R1265 B.n299 B.n298 585
R1266 B.n300 B.n101 585
R1267 B.n302 B.n301 585
R1268 B.n303 B.n100 585
R1269 B.n305 B.n304 585
R1270 B.n306 B.n99 585
R1271 B.n308 B.n307 585
R1272 B.n309 B.n98 585
R1273 B.n311 B.n310 585
R1274 B.n312 B.n97 585
R1275 B.n314 B.n313 585
R1276 B.n315 B.n96 585
R1277 B.n317 B.n316 585
R1278 B.n318 B.n95 585
R1279 B.n320 B.n319 585
R1280 B.n321 B.n94 585
R1281 B.n323 B.n322 585
R1282 B.n324 B.n93 585
R1283 B.n326 B.n325 585
R1284 B.n327 B.n92 585
R1285 B.n329 B.n328 585
R1286 B.n330 B.n91 585
R1287 B.n332 B.n331 585
R1288 B.n333 B.n90 585
R1289 B.n335 B.n334 585
R1290 B.n336 B.n89 585
R1291 B.n338 B.n337 585
R1292 B.n339 B.n88 585
R1293 B.n180 B.n145 585
R1294 B.n179 B.n178 585
R1295 B.n177 B.n146 585
R1296 B.n176 B.n175 585
R1297 B.n174 B.n147 585
R1298 B.n173 B.n172 585
R1299 B.n171 B.n148 585
R1300 B.n170 B.n169 585
R1301 B.n168 B.n149 585
R1302 B.n167 B.n166 585
R1303 B.n165 B.n150 585
R1304 B.n164 B.n163 585
R1305 B.n162 B.n151 585
R1306 B.n161 B.n160 585
R1307 B.n159 B.n152 585
R1308 B.n158 B.n157 585
R1309 B.n156 B.n153 585
R1310 B.n155 B.n154 585
R1311 B.n2 B.n0 585
R1312 B.n585 B.n1 585
R1313 B.n584 B.n583 585
R1314 B.n582 B.n3 585
R1315 B.n581 B.n580 585
R1316 B.n579 B.n4 585
R1317 B.n578 B.n577 585
R1318 B.n576 B.n5 585
R1319 B.n575 B.n574 585
R1320 B.n573 B.n6 585
R1321 B.n572 B.n571 585
R1322 B.n570 B.n7 585
R1323 B.n569 B.n568 585
R1324 B.n567 B.n8 585
R1325 B.n566 B.n565 585
R1326 B.n564 B.n9 585
R1327 B.n563 B.n562 585
R1328 B.n561 B.n10 585
R1329 B.n560 B.n559 585
R1330 B.n558 B.n11 585
R1331 B.n587 B.n586 585
R1332 B.n182 B.n145 497.305
R1333 B.n556 B.n11 497.305
R1334 B.n340 B.n339 497.305
R1335 B.n399 B.n398 497.305
R1336 B.n112 B.t2 427.981
R1337 B.n42 B.t4 427.981
R1338 B.n120 B.t11 427.981
R1339 B.n36 B.t7 427.981
R1340 B.n113 B.t1 413.824
R1341 B.n43 B.t5 413.824
R1342 B.n121 B.t10 413.824
R1343 B.n37 B.t8 413.824
R1344 B.n178 B.n145 163.367
R1345 B.n178 B.n177 163.367
R1346 B.n177 B.n176 163.367
R1347 B.n176 B.n147 163.367
R1348 B.n172 B.n147 163.367
R1349 B.n172 B.n171 163.367
R1350 B.n171 B.n170 163.367
R1351 B.n170 B.n149 163.367
R1352 B.n166 B.n149 163.367
R1353 B.n166 B.n165 163.367
R1354 B.n165 B.n164 163.367
R1355 B.n164 B.n151 163.367
R1356 B.n160 B.n151 163.367
R1357 B.n160 B.n159 163.367
R1358 B.n159 B.n158 163.367
R1359 B.n158 B.n153 163.367
R1360 B.n154 B.n153 163.367
R1361 B.n154 B.n2 163.367
R1362 B.n586 B.n2 163.367
R1363 B.n586 B.n585 163.367
R1364 B.n585 B.n584 163.367
R1365 B.n584 B.n3 163.367
R1366 B.n580 B.n3 163.367
R1367 B.n580 B.n579 163.367
R1368 B.n579 B.n578 163.367
R1369 B.n578 B.n5 163.367
R1370 B.n574 B.n5 163.367
R1371 B.n574 B.n573 163.367
R1372 B.n573 B.n572 163.367
R1373 B.n572 B.n7 163.367
R1374 B.n568 B.n7 163.367
R1375 B.n568 B.n567 163.367
R1376 B.n567 B.n566 163.367
R1377 B.n566 B.n9 163.367
R1378 B.n562 B.n9 163.367
R1379 B.n562 B.n561 163.367
R1380 B.n561 B.n560 163.367
R1381 B.n560 B.n11 163.367
R1382 B.n183 B.n182 163.367
R1383 B.n184 B.n183 163.367
R1384 B.n184 B.n143 163.367
R1385 B.n188 B.n143 163.367
R1386 B.n189 B.n188 163.367
R1387 B.n190 B.n189 163.367
R1388 B.n190 B.n141 163.367
R1389 B.n194 B.n141 163.367
R1390 B.n195 B.n194 163.367
R1391 B.n196 B.n195 163.367
R1392 B.n196 B.n139 163.367
R1393 B.n200 B.n139 163.367
R1394 B.n201 B.n200 163.367
R1395 B.n202 B.n201 163.367
R1396 B.n202 B.n137 163.367
R1397 B.n206 B.n137 163.367
R1398 B.n207 B.n206 163.367
R1399 B.n208 B.n207 163.367
R1400 B.n208 B.n135 163.367
R1401 B.n212 B.n135 163.367
R1402 B.n213 B.n212 163.367
R1403 B.n214 B.n213 163.367
R1404 B.n214 B.n133 163.367
R1405 B.n218 B.n133 163.367
R1406 B.n219 B.n218 163.367
R1407 B.n220 B.n219 163.367
R1408 B.n220 B.n131 163.367
R1409 B.n224 B.n131 163.367
R1410 B.n225 B.n224 163.367
R1411 B.n226 B.n225 163.367
R1412 B.n226 B.n129 163.367
R1413 B.n230 B.n129 163.367
R1414 B.n231 B.n230 163.367
R1415 B.n232 B.n231 163.367
R1416 B.n232 B.n127 163.367
R1417 B.n236 B.n127 163.367
R1418 B.n237 B.n236 163.367
R1419 B.n238 B.n237 163.367
R1420 B.n238 B.n125 163.367
R1421 B.n242 B.n125 163.367
R1422 B.n243 B.n242 163.367
R1423 B.n244 B.n243 163.367
R1424 B.n244 B.n123 163.367
R1425 B.n248 B.n123 163.367
R1426 B.n249 B.n248 163.367
R1427 B.n250 B.n249 163.367
R1428 B.n250 B.n119 163.367
R1429 B.n255 B.n119 163.367
R1430 B.n256 B.n255 163.367
R1431 B.n257 B.n256 163.367
R1432 B.n257 B.n117 163.367
R1433 B.n261 B.n117 163.367
R1434 B.n262 B.n261 163.367
R1435 B.n263 B.n262 163.367
R1436 B.n263 B.n115 163.367
R1437 B.n267 B.n115 163.367
R1438 B.n268 B.n267 163.367
R1439 B.n268 B.n111 163.367
R1440 B.n272 B.n111 163.367
R1441 B.n273 B.n272 163.367
R1442 B.n274 B.n273 163.367
R1443 B.n274 B.n109 163.367
R1444 B.n278 B.n109 163.367
R1445 B.n279 B.n278 163.367
R1446 B.n280 B.n279 163.367
R1447 B.n280 B.n107 163.367
R1448 B.n284 B.n107 163.367
R1449 B.n285 B.n284 163.367
R1450 B.n286 B.n285 163.367
R1451 B.n286 B.n105 163.367
R1452 B.n290 B.n105 163.367
R1453 B.n291 B.n290 163.367
R1454 B.n292 B.n291 163.367
R1455 B.n292 B.n103 163.367
R1456 B.n296 B.n103 163.367
R1457 B.n297 B.n296 163.367
R1458 B.n298 B.n297 163.367
R1459 B.n298 B.n101 163.367
R1460 B.n302 B.n101 163.367
R1461 B.n303 B.n302 163.367
R1462 B.n304 B.n303 163.367
R1463 B.n304 B.n99 163.367
R1464 B.n308 B.n99 163.367
R1465 B.n309 B.n308 163.367
R1466 B.n310 B.n309 163.367
R1467 B.n310 B.n97 163.367
R1468 B.n314 B.n97 163.367
R1469 B.n315 B.n314 163.367
R1470 B.n316 B.n315 163.367
R1471 B.n316 B.n95 163.367
R1472 B.n320 B.n95 163.367
R1473 B.n321 B.n320 163.367
R1474 B.n322 B.n321 163.367
R1475 B.n322 B.n93 163.367
R1476 B.n326 B.n93 163.367
R1477 B.n327 B.n326 163.367
R1478 B.n328 B.n327 163.367
R1479 B.n328 B.n91 163.367
R1480 B.n332 B.n91 163.367
R1481 B.n333 B.n332 163.367
R1482 B.n334 B.n333 163.367
R1483 B.n334 B.n89 163.367
R1484 B.n338 B.n89 163.367
R1485 B.n339 B.n338 163.367
R1486 B.n340 B.n87 163.367
R1487 B.n344 B.n87 163.367
R1488 B.n345 B.n344 163.367
R1489 B.n346 B.n345 163.367
R1490 B.n346 B.n85 163.367
R1491 B.n350 B.n85 163.367
R1492 B.n351 B.n350 163.367
R1493 B.n352 B.n351 163.367
R1494 B.n352 B.n83 163.367
R1495 B.n356 B.n83 163.367
R1496 B.n357 B.n356 163.367
R1497 B.n358 B.n357 163.367
R1498 B.n358 B.n81 163.367
R1499 B.n362 B.n81 163.367
R1500 B.n363 B.n362 163.367
R1501 B.n364 B.n363 163.367
R1502 B.n364 B.n79 163.367
R1503 B.n368 B.n79 163.367
R1504 B.n369 B.n368 163.367
R1505 B.n370 B.n369 163.367
R1506 B.n370 B.n77 163.367
R1507 B.n374 B.n77 163.367
R1508 B.n375 B.n374 163.367
R1509 B.n376 B.n375 163.367
R1510 B.n376 B.n75 163.367
R1511 B.n380 B.n75 163.367
R1512 B.n381 B.n380 163.367
R1513 B.n382 B.n381 163.367
R1514 B.n382 B.n73 163.367
R1515 B.n386 B.n73 163.367
R1516 B.n387 B.n386 163.367
R1517 B.n388 B.n387 163.367
R1518 B.n388 B.n71 163.367
R1519 B.n392 B.n71 163.367
R1520 B.n393 B.n392 163.367
R1521 B.n394 B.n393 163.367
R1522 B.n394 B.n69 163.367
R1523 B.n398 B.n69 163.367
R1524 B.n556 B.n555 163.367
R1525 B.n555 B.n554 163.367
R1526 B.n554 B.n13 163.367
R1527 B.n550 B.n13 163.367
R1528 B.n550 B.n549 163.367
R1529 B.n549 B.n548 163.367
R1530 B.n548 B.n15 163.367
R1531 B.n544 B.n15 163.367
R1532 B.n544 B.n543 163.367
R1533 B.n543 B.n542 163.367
R1534 B.n542 B.n17 163.367
R1535 B.n538 B.n17 163.367
R1536 B.n538 B.n537 163.367
R1537 B.n537 B.n536 163.367
R1538 B.n536 B.n19 163.367
R1539 B.n532 B.n19 163.367
R1540 B.n532 B.n531 163.367
R1541 B.n531 B.n530 163.367
R1542 B.n530 B.n21 163.367
R1543 B.n526 B.n21 163.367
R1544 B.n526 B.n525 163.367
R1545 B.n525 B.n524 163.367
R1546 B.n524 B.n23 163.367
R1547 B.n520 B.n23 163.367
R1548 B.n520 B.n519 163.367
R1549 B.n519 B.n518 163.367
R1550 B.n518 B.n25 163.367
R1551 B.n514 B.n25 163.367
R1552 B.n514 B.n513 163.367
R1553 B.n513 B.n512 163.367
R1554 B.n512 B.n27 163.367
R1555 B.n508 B.n27 163.367
R1556 B.n508 B.n507 163.367
R1557 B.n507 B.n506 163.367
R1558 B.n506 B.n29 163.367
R1559 B.n502 B.n29 163.367
R1560 B.n502 B.n501 163.367
R1561 B.n501 B.n500 163.367
R1562 B.n500 B.n31 163.367
R1563 B.n496 B.n31 163.367
R1564 B.n496 B.n495 163.367
R1565 B.n495 B.n494 163.367
R1566 B.n494 B.n33 163.367
R1567 B.n490 B.n33 163.367
R1568 B.n490 B.n489 163.367
R1569 B.n489 B.n488 163.367
R1570 B.n488 B.n35 163.367
R1571 B.n483 B.n35 163.367
R1572 B.n483 B.n482 163.367
R1573 B.n482 B.n481 163.367
R1574 B.n481 B.n39 163.367
R1575 B.n477 B.n39 163.367
R1576 B.n477 B.n476 163.367
R1577 B.n476 B.n475 163.367
R1578 B.n475 B.n41 163.367
R1579 B.n471 B.n41 163.367
R1580 B.n471 B.n470 163.367
R1581 B.n470 B.n45 163.367
R1582 B.n466 B.n45 163.367
R1583 B.n466 B.n465 163.367
R1584 B.n465 B.n464 163.367
R1585 B.n464 B.n47 163.367
R1586 B.n460 B.n47 163.367
R1587 B.n460 B.n459 163.367
R1588 B.n459 B.n458 163.367
R1589 B.n458 B.n49 163.367
R1590 B.n454 B.n49 163.367
R1591 B.n454 B.n453 163.367
R1592 B.n453 B.n452 163.367
R1593 B.n452 B.n51 163.367
R1594 B.n448 B.n51 163.367
R1595 B.n448 B.n447 163.367
R1596 B.n447 B.n446 163.367
R1597 B.n446 B.n53 163.367
R1598 B.n442 B.n53 163.367
R1599 B.n442 B.n441 163.367
R1600 B.n441 B.n440 163.367
R1601 B.n440 B.n55 163.367
R1602 B.n436 B.n55 163.367
R1603 B.n436 B.n435 163.367
R1604 B.n435 B.n434 163.367
R1605 B.n434 B.n57 163.367
R1606 B.n430 B.n57 163.367
R1607 B.n430 B.n429 163.367
R1608 B.n429 B.n428 163.367
R1609 B.n428 B.n59 163.367
R1610 B.n424 B.n59 163.367
R1611 B.n424 B.n423 163.367
R1612 B.n423 B.n422 163.367
R1613 B.n422 B.n61 163.367
R1614 B.n418 B.n61 163.367
R1615 B.n418 B.n417 163.367
R1616 B.n417 B.n416 163.367
R1617 B.n416 B.n63 163.367
R1618 B.n412 B.n63 163.367
R1619 B.n412 B.n411 163.367
R1620 B.n411 B.n410 163.367
R1621 B.n410 B.n65 163.367
R1622 B.n406 B.n65 163.367
R1623 B.n406 B.n405 163.367
R1624 B.n405 B.n404 163.367
R1625 B.n404 B.n67 163.367
R1626 B.n400 B.n67 163.367
R1627 B.n400 B.n399 163.367
R1628 B.n114 B.n113 59.5399
R1629 B.n253 B.n121 59.5399
R1630 B.n485 B.n37 59.5399
R1631 B.n44 B.n43 59.5399
R1632 B.n558 B.n557 32.3127
R1633 B.n397 B.n68 32.3127
R1634 B.n341 B.n88 32.3127
R1635 B.n181 B.n180 32.3127
R1636 B B.n587 18.0485
R1637 B.n113 B.n112 14.1581
R1638 B.n121 B.n120 14.1581
R1639 B.n37 B.n36 14.1581
R1640 B.n43 B.n42 14.1581
R1641 B.n557 B.n12 10.6151
R1642 B.n553 B.n12 10.6151
R1643 B.n553 B.n552 10.6151
R1644 B.n552 B.n551 10.6151
R1645 B.n551 B.n14 10.6151
R1646 B.n547 B.n14 10.6151
R1647 B.n547 B.n546 10.6151
R1648 B.n546 B.n545 10.6151
R1649 B.n545 B.n16 10.6151
R1650 B.n541 B.n16 10.6151
R1651 B.n541 B.n540 10.6151
R1652 B.n540 B.n539 10.6151
R1653 B.n539 B.n18 10.6151
R1654 B.n535 B.n18 10.6151
R1655 B.n535 B.n534 10.6151
R1656 B.n534 B.n533 10.6151
R1657 B.n533 B.n20 10.6151
R1658 B.n529 B.n20 10.6151
R1659 B.n529 B.n528 10.6151
R1660 B.n528 B.n527 10.6151
R1661 B.n527 B.n22 10.6151
R1662 B.n523 B.n22 10.6151
R1663 B.n523 B.n522 10.6151
R1664 B.n522 B.n521 10.6151
R1665 B.n521 B.n24 10.6151
R1666 B.n517 B.n24 10.6151
R1667 B.n517 B.n516 10.6151
R1668 B.n516 B.n515 10.6151
R1669 B.n515 B.n26 10.6151
R1670 B.n511 B.n26 10.6151
R1671 B.n511 B.n510 10.6151
R1672 B.n510 B.n509 10.6151
R1673 B.n509 B.n28 10.6151
R1674 B.n505 B.n28 10.6151
R1675 B.n505 B.n504 10.6151
R1676 B.n504 B.n503 10.6151
R1677 B.n503 B.n30 10.6151
R1678 B.n499 B.n30 10.6151
R1679 B.n499 B.n498 10.6151
R1680 B.n498 B.n497 10.6151
R1681 B.n497 B.n32 10.6151
R1682 B.n493 B.n32 10.6151
R1683 B.n493 B.n492 10.6151
R1684 B.n492 B.n491 10.6151
R1685 B.n491 B.n34 10.6151
R1686 B.n487 B.n34 10.6151
R1687 B.n487 B.n486 10.6151
R1688 B.n484 B.n38 10.6151
R1689 B.n480 B.n38 10.6151
R1690 B.n480 B.n479 10.6151
R1691 B.n479 B.n478 10.6151
R1692 B.n478 B.n40 10.6151
R1693 B.n474 B.n40 10.6151
R1694 B.n474 B.n473 10.6151
R1695 B.n473 B.n472 10.6151
R1696 B.n469 B.n468 10.6151
R1697 B.n468 B.n467 10.6151
R1698 B.n467 B.n46 10.6151
R1699 B.n463 B.n46 10.6151
R1700 B.n463 B.n462 10.6151
R1701 B.n462 B.n461 10.6151
R1702 B.n461 B.n48 10.6151
R1703 B.n457 B.n48 10.6151
R1704 B.n457 B.n456 10.6151
R1705 B.n456 B.n455 10.6151
R1706 B.n455 B.n50 10.6151
R1707 B.n451 B.n50 10.6151
R1708 B.n451 B.n450 10.6151
R1709 B.n450 B.n449 10.6151
R1710 B.n449 B.n52 10.6151
R1711 B.n445 B.n52 10.6151
R1712 B.n445 B.n444 10.6151
R1713 B.n444 B.n443 10.6151
R1714 B.n443 B.n54 10.6151
R1715 B.n439 B.n54 10.6151
R1716 B.n439 B.n438 10.6151
R1717 B.n438 B.n437 10.6151
R1718 B.n437 B.n56 10.6151
R1719 B.n433 B.n56 10.6151
R1720 B.n433 B.n432 10.6151
R1721 B.n432 B.n431 10.6151
R1722 B.n431 B.n58 10.6151
R1723 B.n427 B.n58 10.6151
R1724 B.n427 B.n426 10.6151
R1725 B.n426 B.n425 10.6151
R1726 B.n425 B.n60 10.6151
R1727 B.n421 B.n60 10.6151
R1728 B.n421 B.n420 10.6151
R1729 B.n420 B.n419 10.6151
R1730 B.n419 B.n62 10.6151
R1731 B.n415 B.n62 10.6151
R1732 B.n415 B.n414 10.6151
R1733 B.n414 B.n413 10.6151
R1734 B.n413 B.n64 10.6151
R1735 B.n409 B.n64 10.6151
R1736 B.n409 B.n408 10.6151
R1737 B.n408 B.n407 10.6151
R1738 B.n407 B.n66 10.6151
R1739 B.n403 B.n66 10.6151
R1740 B.n403 B.n402 10.6151
R1741 B.n402 B.n401 10.6151
R1742 B.n401 B.n68 10.6151
R1743 B.n342 B.n341 10.6151
R1744 B.n343 B.n342 10.6151
R1745 B.n343 B.n86 10.6151
R1746 B.n347 B.n86 10.6151
R1747 B.n348 B.n347 10.6151
R1748 B.n349 B.n348 10.6151
R1749 B.n349 B.n84 10.6151
R1750 B.n353 B.n84 10.6151
R1751 B.n354 B.n353 10.6151
R1752 B.n355 B.n354 10.6151
R1753 B.n355 B.n82 10.6151
R1754 B.n359 B.n82 10.6151
R1755 B.n360 B.n359 10.6151
R1756 B.n361 B.n360 10.6151
R1757 B.n361 B.n80 10.6151
R1758 B.n365 B.n80 10.6151
R1759 B.n366 B.n365 10.6151
R1760 B.n367 B.n366 10.6151
R1761 B.n367 B.n78 10.6151
R1762 B.n371 B.n78 10.6151
R1763 B.n372 B.n371 10.6151
R1764 B.n373 B.n372 10.6151
R1765 B.n373 B.n76 10.6151
R1766 B.n377 B.n76 10.6151
R1767 B.n378 B.n377 10.6151
R1768 B.n379 B.n378 10.6151
R1769 B.n379 B.n74 10.6151
R1770 B.n383 B.n74 10.6151
R1771 B.n384 B.n383 10.6151
R1772 B.n385 B.n384 10.6151
R1773 B.n385 B.n72 10.6151
R1774 B.n389 B.n72 10.6151
R1775 B.n390 B.n389 10.6151
R1776 B.n391 B.n390 10.6151
R1777 B.n391 B.n70 10.6151
R1778 B.n395 B.n70 10.6151
R1779 B.n396 B.n395 10.6151
R1780 B.n397 B.n396 10.6151
R1781 B.n181 B.n144 10.6151
R1782 B.n185 B.n144 10.6151
R1783 B.n186 B.n185 10.6151
R1784 B.n187 B.n186 10.6151
R1785 B.n187 B.n142 10.6151
R1786 B.n191 B.n142 10.6151
R1787 B.n192 B.n191 10.6151
R1788 B.n193 B.n192 10.6151
R1789 B.n193 B.n140 10.6151
R1790 B.n197 B.n140 10.6151
R1791 B.n198 B.n197 10.6151
R1792 B.n199 B.n198 10.6151
R1793 B.n199 B.n138 10.6151
R1794 B.n203 B.n138 10.6151
R1795 B.n204 B.n203 10.6151
R1796 B.n205 B.n204 10.6151
R1797 B.n205 B.n136 10.6151
R1798 B.n209 B.n136 10.6151
R1799 B.n210 B.n209 10.6151
R1800 B.n211 B.n210 10.6151
R1801 B.n211 B.n134 10.6151
R1802 B.n215 B.n134 10.6151
R1803 B.n216 B.n215 10.6151
R1804 B.n217 B.n216 10.6151
R1805 B.n217 B.n132 10.6151
R1806 B.n221 B.n132 10.6151
R1807 B.n222 B.n221 10.6151
R1808 B.n223 B.n222 10.6151
R1809 B.n223 B.n130 10.6151
R1810 B.n227 B.n130 10.6151
R1811 B.n228 B.n227 10.6151
R1812 B.n229 B.n228 10.6151
R1813 B.n229 B.n128 10.6151
R1814 B.n233 B.n128 10.6151
R1815 B.n234 B.n233 10.6151
R1816 B.n235 B.n234 10.6151
R1817 B.n235 B.n126 10.6151
R1818 B.n239 B.n126 10.6151
R1819 B.n240 B.n239 10.6151
R1820 B.n241 B.n240 10.6151
R1821 B.n241 B.n124 10.6151
R1822 B.n245 B.n124 10.6151
R1823 B.n246 B.n245 10.6151
R1824 B.n247 B.n246 10.6151
R1825 B.n247 B.n122 10.6151
R1826 B.n251 B.n122 10.6151
R1827 B.n252 B.n251 10.6151
R1828 B.n254 B.n118 10.6151
R1829 B.n258 B.n118 10.6151
R1830 B.n259 B.n258 10.6151
R1831 B.n260 B.n259 10.6151
R1832 B.n260 B.n116 10.6151
R1833 B.n264 B.n116 10.6151
R1834 B.n265 B.n264 10.6151
R1835 B.n266 B.n265 10.6151
R1836 B.n270 B.n269 10.6151
R1837 B.n271 B.n270 10.6151
R1838 B.n271 B.n110 10.6151
R1839 B.n275 B.n110 10.6151
R1840 B.n276 B.n275 10.6151
R1841 B.n277 B.n276 10.6151
R1842 B.n277 B.n108 10.6151
R1843 B.n281 B.n108 10.6151
R1844 B.n282 B.n281 10.6151
R1845 B.n283 B.n282 10.6151
R1846 B.n283 B.n106 10.6151
R1847 B.n287 B.n106 10.6151
R1848 B.n288 B.n287 10.6151
R1849 B.n289 B.n288 10.6151
R1850 B.n289 B.n104 10.6151
R1851 B.n293 B.n104 10.6151
R1852 B.n294 B.n293 10.6151
R1853 B.n295 B.n294 10.6151
R1854 B.n295 B.n102 10.6151
R1855 B.n299 B.n102 10.6151
R1856 B.n300 B.n299 10.6151
R1857 B.n301 B.n300 10.6151
R1858 B.n301 B.n100 10.6151
R1859 B.n305 B.n100 10.6151
R1860 B.n306 B.n305 10.6151
R1861 B.n307 B.n306 10.6151
R1862 B.n307 B.n98 10.6151
R1863 B.n311 B.n98 10.6151
R1864 B.n312 B.n311 10.6151
R1865 B.n313 B.n312 10.6151
R1866 B.n313 B.n96 10.6151
R1867 B.n317 B.n96 10.6151
R1868 B.n318 B.n317 10.6151
R1869 B.n319 B.n318 10.6151
R1870 B.n319 B.n94 10.6151
R1871 B.n323 B.n94 10.6151
R1872 B.n324 B.n323 10.6151
R1873 B.n325 B.n324 10.6151
R1874 B.n325 B.n92 10.6151
R1875 B.n329 B.n92 10.6151
R1876 B.n330 B.n329 10.6151
R1877 B.n331 B.n330 10.6151
R1878 B.n331 B.n90 10.6151
R1879 B.n335 B.n90 10.6151
R1880 B.n336 B.n335 10.6151
R1881 B.n337 B.n336 10.6151
R1882 B.n337 B.n88 10.6151
R1883 B.n180 B.n179 10.6151
R1884 B.n179 B.n146 10.6151
R1885 B.n175 B.n146 10.6151
R1886 B.n175 B.n174 10.6151
R1887 B.n174 B.n173 10.6151
R1888 B.n173 B.n148 10.6151
R1889 B.n169 B.n148 10.6151
R1890 B.n169 B.n168 10.6151
R1891 B.n168 B.n167 10.6151
R1892 B.n167 B.n150 10.6151
R1893 B.n163 B.n150 10.6151
R1894 B.n163 B.n162 10.6151
R1895 B.n162 B.n161 10.6151
R1896 B.n161 B.n152 10.6151
R1897 B.n157 B.n152 10.6151
R1898 B.n157 B.n156 10.6151
R1899 B.n156 B.n155 10.6151
R1900 B.n155 B.n0 10.6151
R1901 B.n583 B.n1 10.6151
R1902 B.n583 B.n582 10.6151
R1903 B.n582 B.n581 10.6151
R1904 B.n581 B.n4 10.6151
R1905 B.n577 B.n4 10.6151
R1906 B.n577 B.n576 10.6151
R1907 B.n576 B.n575 10.6151
R1908 B.n575 B.n6 10.6151
R1909 B.n571 B.n6 10.6151
R1910 B.n571 B.n570 10.6151
R1911 B.n570 B.n569 10.6151
R1912 B.n569 B.n8 10.6151
R1913 B.n565 B.n8 10.6151
R1914 B.n565 B.n564 10.6151
R1915 B.n564 B.n563 10.6151
R1916 B.n563 B.n10 10.6151
R1917 B.n559 B.n10 10.6151
R1918 B.n559 B.n558 10.6151
R1919 B.n485 B.n484 6.5566
R1920 B.n472 B.n44 6.5566
R1921 B.n254 B.n253 6.5566
R1922 B.n266 B.n114 6.5566
R1923 B.n486 B.n485 4.05904
R1924 B.n469 B.n44 4.05904
R1925 B.n253 B.n252 4.05904
R1926 B.n269 B.n114 4.05904
R1927 B.n587 B.n0 2.81026
R1928 B.n587 B.n1 2.81026
C0 B w_n1700_n3792# 7.34554f
C1 VN w_n1700_n3792# 2.87388f
C2 VDD2 VP 0.285404f
C3 B VP 1.08405f
C4 VP VN 5.35789f
C5 VDD2 B 1.06295f
C6 VDD2 VN 4.65422f
C7 VDD1 VTAIL 16.585901f
C8 B VN 0.736688f
C9 VDD1 w_n1700_n3792# 1.22812f
C10 VTAIL w_n1700_n3792# 4.80617f
C11 VP VDD1 4.79175f
C12 VDD2 VDD1 0.676501f
C13 VP VTAIL 4.19628f
C14 B VDD1 1.03554f
C15 VN VDD1 0.147587f
C16 VDD2 VTAIL 16.6255f
C17 B VTAIL 4.12392f
C18 VN VTAIL 4.18217f
C19 VP w_n1700_n3792# 3.08809f
C20 VDD2 w_n1700_n3792# 1.25053f
C21 VDD2 VSUBS 1.38527f
C22 VDD1 VSUBS 1.638804f
C23 VTAIL VSUBS 0.838951f
C24 VN VSUBS 4.7524f
C25 VP VSUBS 1.431837f
C26 B VSUBS 2.72461f
C27 w_n1700_n3792# VSUBS 79.1316f
C28 B.n0 VSUBS 0.005241f
C29 B.n1 VSUBS 0.005241f
C30 B.n2 VSUBS 0.008289f
C31 B.n3 VSUBS 0.008289f
C32 B.n4 VSUBS 0.008289f
C33 B.n5 VSUBS 0.008289f
C34 B.n6 VSUBS 0.008289f
C35 B.n7 VSUBS 0.008289f
C36 B.n8 VSUBS 0.008289f
C37 B.n9 VSUBS 0.008289f
C38 B.n10 VSUBS 0.008289f
C39 B.n11 VSUBS 0.01903f
C40 B.n12 VSUBS 0.008289f
C41 B.n13 VSUBS 0.008289f
C42 B.n14 VSUBS 0.008289f
C43 B.n15 VSUBS 0.008289f
C44 B.n16 VSUBS 0.008289f
C45 B.n17 VSUBS 0.008289f
C46 B.n18 VSUBS 0.008289f
C47 B.n19 VSUBS 0.008289f
C48 B.n20 VSUBS 0.008289f
C49 B.n21 VSUBS 0.008289f
C50 B.n22 VSUBS 0.008289f
C51 B.n23 VSUBS 0.008289f
C52 B.n24 VSUBS 0.008289f
C53 B.n25 VSUBS 0.008289f
C54 B.n26 VSUBS 0.008289f
C55 B.n27 VSUBS 0.008289f
C56 B.n28 VSUBS 0.008289f
C57 B.n29 VSUBS 0.008289f
C58 B.n30 VSUBS 0.008289f
C59 B.n31 VSUBS 0.008289f
C60 B.n32 VSUBS 0.008289f
C61 B.n33 VSUBS 0.008289f
C62 B.n34 VSUBS 0.008289f
C63 B.n35 VSUBS 0.008289f
C64 B.t8 VSUBS 0.306883f
C65 B.t7 VSUBS 0.317116f
C66 B.t6 VSUBS 0.26457f
C67 B.n36 VSUBS 0.384011f
C68 B.n37 VSUBS 0.321167f
C69 B.n38 VSUBS 0.008289f
C70 B.n39 VSUBS 0.008289f
C71 B.n40 VSUBS 0.008289f
C72 B.n41 VSUBS 0.008289f
C73 B.t5 VSUBS 0.306887f
C74 B.t4 VSUBS 0.31712f
C75 B.t3 VSUBS 0.26457f
C76 B.n42 VSUBS 0.384007f
C77 B.n43 VSUBS 0.321163f
C78 B.n44 VSUBS 0.019204f
C79 B.n45 VSUBS 0.008289f
C80 B.n46 VSUBS 0.008289f
C81 B.n47 VSUBS 0.008289f
C82 B.n48 VSUBS 0.008289f
C83 B.n49 VSUBS 0.008289f
C84 B.n50 VSUBS 0.008289f
C85 B.n51 VSUBS 0.008289f
C86 B.n52 VSUBS 0.008289f
C87 B.n53 VSUBS 0.008289f
C88 B.n54 VSUBS 0.008289f
C89 B.n55 VSUBS 0.008289f
C90 B.n56 VSUBS 0.008289f
C91 B.n57 VSUBS 0.008289f
C92 B.n58 VSUBS 0.008289f
C93 B.n59 VSUBS 0.008289f
C94 B.n60 VSUBS 0.008289f
C95 B.n61 VSUBS 0.008289f
C96 B.n62 VSUBS 0.008289f
C97 B.n63 VSUBS 0.008289f
C98 B.n64 VSUBS 0.008289f
C99 B.n65 VSUBS 0.008289f
C100 B.n66 VSUBS 0.008289f
C101 B.n67 VSUBS 0.008289f
C102 B.n68 VSUBS 0.018499f
C103 B.n69 VSUBS 0.008289f
C104 B.n70 VSUBS 0.008289f
C105 B.n71 VSUBS 0.008289f
C106 B.n72 VSUBS 0.008289f
C107 B.n73 VSUBS 0.008289f
C108 B.n74 VSUBS 0.008289f
C109 B.n75 VSUBS 0.008289f
C110 B.n76 VSUBS 0.008289f
C111 B.n77 VSUBS 0.008289f
C112 B.n78 VSUBS 0.008289f
C113 B.n79 VSUBS 0.008289f
C114 B.n80 VSUBS 0.008289f
C115 B.n81 VSUBS 0.008289f
C116 B.n82 VSUBS 0.008289f
C117 B.n83 VSUBS 0.008289f
C118 B.n84 VSUBS 0.008289f
C119 B.n85 VSUBS 0.008289f
C120 B.n86 VSUBS 0.008289f
C121 B.n87 VSUBS 0.008289f
C122 B.n88 VSUBS 0.019489f
C123 B.n89 VSUBS 0.008289f
C124 B.n90 VSUBS 0.008289f
C125 B.n91 VSUBS 0.008289f
C126 B.n92 VSUBS 0.008289f
C127 B.n93 VSUBS 0.008289f
C128 B.n94 VSUBS 0.008289f
C129 B.n95 VSUBS 0.008289f
C130 B.n96 VSUBS 0.008289f
C131 B.n97 VSUBS 0.008289f
C132 B.n98 VSUBS 0.008289f
C133 B.n99 VSUBS 0.008289f
C134 B.n100 VSUBS 0.008289f
C135 B.n101 VSUBS 0.008289f
C136 B.n102 VSUBS 0.008289f
C137 B.n103 VSUBS 0.008289f
C138 B.n104 VSUBS 0.008289f
C139 B.n105 VSUBS 0.008289f
C140 B.n106 VSUBS 0.008289f
C141 B.n107 VSUBS 0.008289f
C142 B.n108 VSUBS 0.008289f
C143 B.n109 VSUBS 0.008289f
C144 B.n110 VSUBS 0.008289f
C145 B.n111 VSUBS 0.008289f
C146 B.t1 VSUBS 0.306887f
C147 B.t2 VSUBS 0.31712f
C148 B.t0 VSUBS 0.26457f
C149 B.n112 VSUBS 0.384007f
C150 B.n113 VSUBS 0.321163f
C151 B.n114 VSUBS 0.019204f
C152 B.n115 VSUBS 0.008289f
C153 B.n116 VSUBS 0.008289f
C154 B.n117 VSUBS 0.008289f
C155 B.n118 VSUBS 0.008289f
C156 B.n119 VSUBS 0.008289f
C157 B.t10 VSUBS 0.306883f
C158 B.t11 VSUBS 0.317116f
C159 B.t9 VSUBS 0.26457f
C160 B.n120 VSUBS 0.384011f
C161 B.n121 VSUBS 0.321167f
C162 B.n122 VSUBS 0.008289f
C163 B.n123 VSUBS 0.008289f
C164 B.n124 VSUBS 0.008289f
C165 B.n125 VSUBS 0.008289f
C166 B.n126 VSUBS 0.008289f
C167 B.n127 VSUBS 0.008289f
C168 B.n128 VSUBS 0.008289f
C169 B.n129 VSUBS 0.008289f
C170 B.n130 VSUBS 0.008289f
C171 B.n131 VSUBS 0.008289f
C172 B.n132 VSUBS 0.008289f
C173 B.n133 VSUBS 0.008289f
C174 B.n134 VSUBS 0.008289f
C175 B.n135 VSUBS 0.008289f
C176 B.n136 VSUBS 0.008289f
C177 B.n137 VSUBS 0.008289f
C178 B.n138 VSUBS 0.008289f
C179 B.n139 VSUBS 0.008289f
C180 B.n140 VSUBS 0.008289f
C181 B.n141 VSUBS 0.008289f
C182 B.n142 VSUBS 0.008289f
C183 B.n143 VSUBS 0.008289f
C184 B.n144 VSUBS 0.008289f
C185 B.n145 VSUBS 0.01903f
C186 B.n146 VSUBS 0.008289f
C187 B.n147 VSUBS 0.008289f
C188 B.n148 VSUBS 0.008289f
C189 B.n149 VSUBS 0.008289f
C190 B.n150 VSUBS 0.008289f
C191 B.n151 VSUBS 0.008289f
C192 B.n152 VSUBS 0.008289f
C193 B.n153 VSUBS 0.008289f
C194 B.n154 VSUBS 0.008289f
C195 B.n155 VSUBS 0.008289f
C196 B.n156 VSUBS 0.008289f
C197 B.n157 VSUBS 0.008289f
C198 B.n158 VSUBS 0.008289f
C199 B.n159 VSUBS 0.008289f
C200 B.n160 VSUBS 0.008289f
C201 B.n161 VSUBS 0.008289f
C202 B.n162 VSUBS 0.008289f
C203 B.n163 VSUBS 0.008289f
C204 B.n164 VSUBS 0.008289f
C205 B.n165 VSUBS 0.008289f
C206 B.n166 VSUBS 0.008289f
C207 B.n167 VSUBS 0.008289f
C208 B.n168 VSUBS 0.008289f
C209 B.n169 VSUBS 0.008289f
C210 B.n170 VSUBS 0.008289f
C211 B.n171 VSUBS 0.008289f
C212 B.n172 VSUBS 0.008289f
C213 B.n173 VSUBS 0.008289f
C214 B.n174 VSUBS 0.008289f
C215 B.n175 VSUBS 0.008289f
C216 B.n176 VSUBS 0.008289f
C217 B.n177 VSUBS 0.008289f
C218 B.n178 VSUBS 0.008289f
C219 B.n179 VSUBS 0.008289f
C220 B.n180 VSUBS 0.01903f
C221 B.n181 VSUBS 0.019489f
C222 B.n182 VSUBS 0.019489f
C223 B.n183 VSUBS 0.008289f
C224 B.n184 VSUBS 0.008289f
C225 B.n185 VSUBS 0.008289f
C226 B.n186 VSUBS 0.008289f
C227 B.n187 VSUBS 0.008289f
C228 B.n188 VSUBS 0.008289f
C229 B.n189 VSUBS 0.008289f
C230 B.n190 VSUBS 0.008289f
C231 B.n191 VSUBS 0.008289f
C232 B.n192 VSUBS 0.008289f
C233 B.n193 VSUBS 0.008289f
C234 B.n194 VSUBS 0.008289f
C235 B.n195 VSUBS 0.008289f
C236 B.n196 VSUBS 0.008289f
C237 B.n197 VSUBS 0.008289f
C238 B.n198 VSUBS 0.008289f
C239 B.n199 VSUBS 0.008289f
C240 B.n200 VSUBS 0.008289f
C241 B.n201 VSUBS 0.008289f
C242 B.n202 VSUBS 0.008289f
C243 B.n203 VSUBS 0.008289f
C244 B.n204 VSUBS 0.008289f
C245 B.n205 VSUBS 0.008289f
C246 B.n206 VSUBS 0.008289f
C247 B.n207 VSUBS 0.008289f
C248 B.n208 VSUBS 0.008289f
C249 B.n209 VSUBS 0.008289f
C250 B.n210 VSUBS 0.008289f
C251 B.n211 VSUBS 0.008289f
C252 B.n212 VSUBS 0.008289f
C253 B.n213 VSUBS 0.008289f
C254 B.n214 VSUBS 0.008289f
C255 B.n215 VSUBS 0.008289f
C256 B.n216 VSUBS 0.008289f
C257 B.n217 VSUBS 0.008289f
C258 B.n218 VSUBS 0.008289f
C259 B.n219 VSUBS 0.008289f
C260 B.n220 VSUBS 0.008289f
C261 B.n221 VSUBS 0.008289f
C262 B.n222 VSUBS 0.008289f
C263 B.n223 VSUBS 0.008289f
C264 B.n224 VSUBS 0.008289f
C265 B.n225 VSUBS 0.008289f
C266 B.n226 VSUBS 0.008289f
C267 B.n227 VSUBS 0.008289f
C268 B.n228 VSUBS 0.008289f
C269 B.n229 VSUBS 0.008289f
C270 B.n230 VSUBS 0.008289f
C271 B.n231 VSUBS 0.008289f
C272 B.n232 VSUBS 0.008289f
C273 B.n233 VSUBS 0.008289f
C274 B.n234 VSUBS 0.008289f
C275 B.n235 VSUBS 0.008289f
C276 B.n236 VSUBS 0.008289f
C277 B.n237 VSUBS 0.008289f
C278 B.n238 VSUBS 0.008289f
C279 B.n239 VSUBS 0.008289f
C280 B.n240 VSUBS 0.008289f
C281 B.n241 VSUBS 0.008289f
C282 B.n242 VSUBS 0.008289f
C283 B.n243 VSUBS 0.008289f
C284 B.n244 VSUBS 0.008289f
C285 B.n245 VSUBS 0.008289f
C286 B.n246 VSUBS 0.008289f
C287 B.n247 VSUBS 0.008289f
C288 B.n248 VSUBS 0.008289f
C289 B.n249 VSUBS 0.008289f
C290 B.n250 VSUBS 0.008289f
C291 B.n251 VSUBS 0.008289f
C292 B.n252 VSUBS 0.005729f
C293 B.n253 VSUBS 0.019204f
C294 B.n254 VSUBS 0.006704f
C295 B.n255 VSUBS 0.008289f
C296 B.n256 VSUBS 0.008289f
C297 B.n257 VSUBS 0.008289f
C298 B.n258 VSUBS 0.008289f
C299 B.n259 VSUBS 0.008289f
C300 B.n260 VSUBS 0.008289f
C301 B.n261 VSUBS 0.008289f
C302 B.n262 VSUBS 0.008289f
C303 B.n263 VSUBS 0.008289f
C304 B.n264 VSUBS 0.008289f
C305 B.n265 VSUBS 0.008289f
C306 B.n266 VSUBS 0.006704f
C307 B.n267 VSUBS 0.008289f
C308 B.n268 VSUBS 0.008289f
C309 B.n269 VSUBS 0.005729f
C310 B.n270 VSUBS 0.008289f
C311 B.n271 VSUBS 0.008289f
C312 B.n272 VSUBS 0.008289f
C313 B.n273 VSUBS 0.008289f
C314 B.n274 VSUBS 0.008289f
C315 B.n275 VSUBS 0.008289f
C316 B.n276 VSUBS 0.008289f
C317 B.n277 VSUBS 0.008289f
C318 B.n278 VSUBS 0.008289f
C319 B.n279 VSUBS 0.008289f
C320 B.n280 VSUBS 0.008289f
C321 B.n281 VSUBS 0.008289f
C322 B.n282 VSUBS 0.008289f
C323 B.n283 VSUBS 0.008289f
C324 B.n284 VSUBS 0.008289f
C325 B.n285 VSUBS 0.008289f
C326 B.n286 VSUBS 0.008289f
C327 B.n287 VSUBS 0.008289f
C328 B.n288 VSUBS 0.008289f
C329 B.n289 VSUBS 0.008289f
C330 B.n290 VSUBS 0.008289f
C331 B.n291 VSUBS 0.008289f
C332 B.n292 VSUBS 0.008289f
C333 B.n293 VSUBS 0.008289f
C334 B.n294 VSUBS 0.008289f
C335 B.n295 VSUBS 0.008289f
C336 B.n296 VSUBS 0.008289f
C337 B.n297 VSUBS 0.008289f
C338 B.n298 VSUBS 0.008289f
C339 B.n299 VSUBS 0.008289f
C340 B.n300 VSUBS 0.008289f
C341 B.n301 VSUBS 0.008289f
C342 B.n302 VSUBS 0.008289f
C343 B.n303 VSUBS 0.008289f
C344 B.n304 VSUBS 0.008289f
C345 B.n305 VSUBS 0.008289f
C346 B.n306 VSUBS 0.008289f
C347 B.n307 VSUBS 0.008289f
C348 B.n308 VSUBS 0.008289f
C349 B.n309 VSUBS 0.008289f
C350 B.n310 VSUBS 0.008289f
C351 B.n311 VSUBS 0.008289f
C352 B.n312 VSUBS 0.008289f
C353 B.n313 VSUBS 0.008289f
C354 B.n314 VSUBS 0.008289f
C355 B.n315 VSUBS 0.008289f
C356 B.n316 VSUBS 0.008289f
C357 B.n317 VSUBS 0.008289f
C358 B.n318 VSUBS 0.008289f
C359 B.n319 VSUBS 0.008289f
C360 B.n320 VSUBS 0.008289f
C361 B.n321 VSUBS 0.008289f
C362 B.n322 VSUBS 0.008289f
C363 B.n323 VSUBS 0.008289f
C364 B.n324 VSUBS 0.008289f
C365 B.n325 VSUBS 0.008289f
C366 B.n326 VSUBS 0.008289f
C367 B.n327 VSUBS 0.008289f
C368 B.n328 VSUBS 0.008289f
C369 B.n329 VSUBS 0.008289f
C370 B.n330 VSUBS 0.008289f
C371 B.n331 VSUBS 0.008289f
C372 B.n332 VSUBS 0.008289f
C373 B.n333 VSUBS 0.008289f
C374 B.n334 VSUBS 0.008289f
C375 B.n335 VSUBS 0.008289f
C376 B.n336 VSUBS 0.008289f
C377 B.n337 VSUBS 0.008289f
C378 B.n338 VSUBS 0.008289f
C379 B.n339 VSUBS 0.019489f
C380 B.n340 VSUBS 0.01903f
C381 B.n341 VSUBS 0.01903f
C382 B.n342 VSUBS 0.008289f
C383 B.n343 VSUBS 0.008289f
C384 B.n344 VSUBS 0.008289f
C385 B.n345 VSUBS 0.008289f
C386 B.n346 VSUBS 0.008289f
C387 B.n347 VSUBS 0.008289f
C388 B.n348 VSUBS 0.008289f
C389 B.n349 VSUBS 0.008289f
C390 B.n350 VSUBS 0.008289f
C391 B.n351 VSUBS 0.008289f
C392 B.n352 VSUBS 0.008289f
C393 B.n353 VSUBS 0.008289f
C394 B.n354 VSUBS 0.008289f
C395 B.n355 VSUBS 0.008289f
C396 B.n356 VSUBS 0.008289f
C397 B.n357 VSUBS 0.008289f
C398 B.n358 VSUBS 0.008289f
C399 B.n359 VSUBS 0.008289f
C400 B.n360 VSUBS 0.008289f
C401 B.n361 VSUBS 0.008289f
C402 B.n362 VSUBS 0.008289f
C403 B.n363 VSUBS 0.008289f
C404 B.n364 VSUBS 0.008289f
C405 B.n365 VSUBS 0.008289f
C406 B.n366 VSUBS 0.008289f
C407 B.n367 VSUBS 0.008289f
C408 B.n368 VSUBS 0.008289f
C409 B.n369 VSUBS 0.008289f
C410 B.n370 VSUBS 0.008289f
C411 B.n371 VSUBS 0.008289f
C412 B.n372 VSUBS 0.008289f
C413 B.n373 VSUBS 0.008289f
C414 B.n374 VSUBS 0.008289f
C415 B.n375 VSUBS 0.008289f
C416 B.n376 VSUBS 0.008289f
C417 B.n377 VSUBS 0.008289f
C418 B.n378 VSUBS 0.008289f
C419 B.n379 VSUBS 0.008289f
C420 B.n380 VSUBS 0.008289f
C421 B.n381 VSUBS 0.008289f
C422 B.n382 VSUBS 0.008289f
C423 B.n383 VSUBS 0.008289f
C424 B.n384 VSUBS 0.008289f
C425 B.n385 VSUBS 0.008289f
C426 B.n386 VSUBS 0.008289f
C427 B.n387 VSUBS 0.008289f
C428 B.n388 VSUBS 0.008289f
C429 B.n389 VSUBS 0.008289f
C430 B.n390 VSUBS 0.008289f
C431 B.n391 VSUBS 0.008289f
C432 B.n392 VSUBS 0.008289f
C433 B.n393 VSUBS 0.008289f
C434 B.n394 VSUBS 0.008289f
C435 B.n395 VSUBS 0.008289f
C436 B.n396 VSUBS 0.008289f
C437 B.n397 VSUBS 0.02002f
C438 B.n398 VSUBS 0.01903f
C439 B.n399 VSUBS 0.019489f
C440 B.n400 VSUBS 0.008289f
C441 B.n401 VSUBS 0.008289f
C442 B.n402 VSUBS 0.008289f
C443 B.n403 VSUBS 0.008289f
C444 B.n404 VSUBS 0.008289f
C445 B.n405 VSUBS 0.008289f
C446 B.n406 VSUBS 0.008289f
C447 B.n407 VSUBS 0.008289f
C448 B.n408 VSUBS 0.008289f
C449 B.n409 VSUBS 0.008289f
C450 B.n410 VSUBS 0.008289f
C451 B.n411 VSUBS 0.008289f
C452 B.n412 VSUBS 0.008289f
C453 B.n413 VSUBS 0.008289f
C454 B.n414 VSUBS 0.008289f
C455 B.n415 VSUBS 0.008289f
C456 B.n416 VSUBS 0.008289f
C457 B.n417 VSUBS 0.008289f
C458 B.n418 VSUBS 0.008289f
C459 B.n419 VSUBS 0.008289f
C460 B.n420 VSUBS 0.008289f
C461 B.n421 VSUBS 0.008289f
C462 B.n422 VSUBS 0.008289f
C463 B.n423 VSUBS 0.008289f
C464 B.n424 VSUBS 0.008289f
C465 B.n425 VSUBS 0.008289f
C466 B.n426 VSUBS 0.008289f
C467 B.n427 VSUBS 0.008289f
C468 B.n428 VSUBS 0.008289f
C469 B.n429 VSUBS 0.008289f
C470 B.n430 VSUBS 0.008289f
C471 B.n431 VSUBS 0.008289f
C472 B.n432 VSUBS 0.008289f
C473 B.n433 VSUBS 0.008289f
C474 B.n434 VSUBS 0.008289f
C475 B.n435 VSUBS 0.008289f
C476 B.n436 VSUBS 0.008289f
C477 B.n437 VSUBS 0.008289f
C478 B.n438 VSUBS 0.008289f
C479 B.n439 VSUBS 0.008289f
C480 B.n440 VSUBS 0.008289f
C481 B.n441 VSUBS 0.008289f
C482 B.n442 VSUBS 0.008289f
C483 B.n443 VSUBS 0.008289f
C484 B.n444 VSUBS 0.008289f
C485 B.n445 VSUBS 0.008289f
C486 B.n446 VSUBS 0.008289f
C487 B.n447 VSUBS 0.008289f
C488 B.n448 VSUBS 0.008289f
C489 B.n449 VSUBS 0.008289f
C490 B.n450 VSUBS 0.008289f
C491 B.n451 VSUBS 0.008289f
C492 B.n452 VSUBS 0.008289f
C493 B.n453 VSUBS 0.008289f
C494 B.n454 VSUBS 0.008289f
C495 B.n455 VSUBS 0.008289f
C496 B.n456 VSUBS 0.008289f
C497 B.n457 VSUBS 0.008289f
C498 B.n458 VSUBS 0.008289f
C499 B.n459 VSUBS 0.008289f
C500 B.n460 VSUBS 0.008289f
C501 B.n461 VSUBS 0.008289f
C502 B.n462 VSUBS 0.008289f
C503 B.n463 VSUBS 0.008289f
C504 B.n464 VSUBS 0.008289f
C505 B.n465 VSUBS 0.008289f
C506 B.n466 VSUBS 0.008289f
C507 B.n467 VSUBS 0.008289f
C508 B.n468 VSUBS 0.008289f
C509 B.n469 VSUBS 0.005729f
C510 B.n470 VSUBS 0.008289f
C511 B.n471 VSUBS 0.008289f
C512 B.n472 VSUBS 0.006704f
C513 B.n473 VSUBS 0.008289f
C514 B.n474 VSUBS 0.008289f
C515 B.n475 VSUBS 0.008289f
C516 B.n476 VSUBS 0.008289f
C517 B.n477 VSUBS 0.008289f
C518 B.n478 VSUBS 0.008289f
C519 B.n479 VSUBS 0.008289f
C520 B.n480 VSUBS 0.008289f
C521 B.n481 VSUBS 0.008289f
C522 B.n482 VSUBS 0.008289f
C523 B.n483 VSUBS 0.008289f
C524 B.n484 VSUBS 0.006704f
C525 B.n485 VSUBS 0.019204f
C526 B.n486 VSUBS 0.005729f
C527 B.n487 VSUBS 0.008289f
C528 B.n488 VSUBS 0.008289f
C529 B.n489 VSUBS 0.008289f
C530 B.n490 VSUBS 0.008289f
C531 B.n491 VSUBS 0.008289f
C532 B.n492 VSUBS 0.008289f
C533 B.n493 VSUBS 0.008289f
C534 B.n494 VSUBS 0.008289f
C535 B.n495 VSUBS 0.008289f
C536 B.n496 VSUBS 0.008289f
C537 B.n497 VSUBS 0.008289f
C538 B.n498 VSUBS 0.008289f
C539 B.n499 VSUBS 0.008289f
C540 B.n500 VSUBS 0.008289f
C541 B.n501 VSUBS 0.008289f
C542 B.n502 VSUBS 0.008289f
C543 B.n503 VSUBS 0.008289f
C544 B.n504 VSUBS 0.008289f
C545 B.n505 VSUBS 0.008289f
C546 B.n506 VSUBS 0.008289f
C547 B.n507 VSUBS 0.008289f
C548 B.n508 VSUBS 0.008289f
C549 B.n509 VSUBS 0.008289f
C550 B.n510 VSUBS 0.008289f
C551 B.n511 VSUBS 0.008289f
C552 B.n512 VSUBS 0.008289f
C553 B.n513 VSUBS 0.008289f
C554 B.n514 VSUBS 0.008289f
C555 B.n515 VSUBS 0.008289f
C556 B.n516 VSUBS 0.008289f
C557 B.n517 VSUBS 0.008289f
C558 B.n518 VSUBS 0.008289f
C559 B.n519 VSUBS 0.008289f
C560 B.n520 VSUBS 0.008289f
C561 B.n521 VSUBS 0.008289f
C562 B.n522 VSUBS 0.008289f
C563 B.n523 VSUBS 0.008289f
C564 B.n524 VSUBS 0.008289f
C565 B.n525 VSUBS 0.008289f
C566 B.n526 VSUBS 0.008289f
C567 B.n527 VSUBS 0.008289f
C568 B.n528 VSUBS 0.008289f
C569 B.n529 VSUBS 0.008289f
C570 B.n530 VSUBS 0.008289f
C571 B.n531 VSUBS 0.008289f
C572 B.n532 VSUBS 0.008289f
C573 B.n533 VSUBS 0.008289f
C574 B.n534 VSUBS 0.008289f
C575 B.n535 VSUBS 0.008289f
C576 B.n536 VSUBS 0.008289f
C577 B.n537 VSUBS 0.008289f
C578 B.n538 VSUBS 0.008289f
C579 B.n539 VSUBS 0.008289f
C580 B.n540 VSUBS 0.008289f
C581 B.n541 VSUBS 0.008289f
C582 B.n542 VSUBS 0.008289f
C583 B.n543 VSUBS 0.008289f
C584 B.n544 VSUBS 0.008289f
C585 B.n545 VSUBS 0.008289f
C586 B.n546 VSUBS 0.008289f
C587 B.n547 VSUBS 0.008289f
C588 B.n548 VSUBS 0.008289f
C589 B.n549 VSUBS 0.008289f
C590 B.n550 VSUBS 0.008289f
C591 B.n551 VSUBS 0.008289f
C592 B.n552 VSUBS 0.008289f
C593 B.n553 VSUBS 0.008289f
C594 B.n554 VSUBS 0.008289f
C595 B.n555 VSUBS 0.008289f
C596 B.n556 VSUBS 0.019489f
C597 B.n557 VSUBS 0.019489f
C598 B.n558 VSUBS 0.01903f
C599 B.n559 VSUBS 0.008289f
C600 B.n560 VSUBS 0.008289f
C601 B.n561 VSUBS 0.008289f
C602 B.n562 VSUBS 0.008289f
C603 B.n563 VSUBS 0.008289f
C604 B.n564 VSUBS 0.008289f
C605 B.n565 VSUBS 0.008289f
C606 B.n566 VSUBS 0.008289f
C607 B.n567 VSUBS 0.008289f
C608 B.n568 VSUBS 0.008289f
C609 B.n569 VSUBS 0.008289f
C610 B.n570 VSUBS 0.008289f
C611 B.n571 VSUBS 0.008289f
C612 B.n572 VSUBS 0.008289f
C613 B.n573 VSUBS 0.008289f
C614 B.n574 VSUBS 0.008289f
C615 B.n575 VSUBS 0.008289f
C616 B.n576 VSUBS 0.008289f
C617 B.n577 VSUBS 0.008289f
C618 B.n578 VSUBS 0.008289f
C619 B.n579 VSUBS 0.008289f
C620 B.n580 VSUBS 0.008289f
C621 B.n581 VSUBS 0.008289f
C622 B.n582 VSUBS 0.008289f
C623 B.n583 VSUBS 0.008289f
C624 B.n584 VSUBS 0.008289f
C625 B.n585 VSUBS 0.008289f
C626 B.n586 VSUBS 0.008289f
C627 B.n587 VSUBS 0.018769f
C628 VDD1.t3 VSUBS 0.347276f
C629 VDD1.t6 VSUBS 0.347276f
C630 VDD1.n0 VSUBS 2.81432f
C631 VDD1.t2 VSUBS 0.347276f
C632 VDD1.t1 VSUBS 0.347276f
C633 VDD1.n1 VSUBS 2.81325f
C634 VDD1.t4 VSUBS 0.347276f
C635 VDD1.t5 VSUBS 0.347276f
C636 VDD1.n2 VSUBS 2.81325f
C637 VDD1.n3 VSUBS 3.34517f
C638 VDD1.t7 VSUBS 0.347276f
C639 VDD1.t0 VSUBS 0.347276f
C640 VDD1.n4 VSUBS 2.81092f
C641 VDD1.n5 VSUBS 3.27947f
C642 VP.n0 VSUBS 0.064465f
C643 VP.t5 VSUBS 1.0443f
C644 VP.n1 VSUBS 0.40692f
C645 VP.n2 VSUBS 0.216354f
C646 VP.t0 VSUBS 1.03554f
C647 VP.t1 VSUBS 1.03554f
C648 VP.t4 VSUBS 1.04947f
C649 VP.n3 VSUBS 0.402242f
C650 VP.n4 VSUBS 0.417265f
C651 VP.n5 VSUBS 0.417265f
C652 VP.t7 VSUBS 1.0443f
C653 VP.n6 VSUBS 0.40692f
C654 VP.n7 VSUBS 2.69767f
C655 VP.n8 VSUBS 2.75254f
C656 VP.n9 VSUBS 0.064465f
C657 VP.t6 VSUBS 1.03554f
C658 VP.n10 VSUBS 0.417265f
C659 VP.t3 VSUBS 1.03554f
C660 VP.n11 VSUBS 0.417265f
C661 VP.t2 VSUBS 1.0443f
C662 VP.n12 VSUBS 0.40692f
C663 VP.n13 VSUBS 0.049958f
C664 VDD2.t0 VSUBS 0.34752f
C665 VDD2.t7 VSUBS 0.34752f
C666 VDD2.n0 VSUBS 2.81523f
C667 VDD2.t4 VSUBS 0.34752f
C668 VDD2.t2 VSUBS 0.34752f
C669 VDD2.n1 VSUBS 2.81523f
C670 VDD2.n2 VSUBS 3.2809f
C671 VDD2.t1 VSUBS 0.34752f
C672 VDD2.t6 VSUBS 0.34752f
C673 VDD2.n3 VSUBS 2.81291f
C674 VDD2.n4 VSUBS 3.24502f
C675 VDD2.t5 VSUBS 0.34752f
C676 VDD2.t3 VSUBS 0.34752f
C677 VDD2.n5 VSUBS 2.81519f
C678 VTAIL.t12 VSUBS 0.299913f
C679 VTAIL.t11 VSUBS 0.299913f
C680 VTAIL.n0 VSUBS 2.28809f
C681 VTAIL.n1 VSUBS 0.657025f
C682 VTAIL.n2 VSUBS 0.028966f
C683 VTAIL.n3 VSUBS 0.026879f
C684 VTAIL.n4 VSUBS 0.014868f
C685 VTAIL.n5 VSUBS 0.034139f
C686 VTAIL.n6 VSUBS 0.015293f
C687 VTAIL.n7 VSUBS 0.026879f
C688 VTAIL.n8 VSUBS 0.014443f
C689 VTAIL.n9 VSUBS 0.034139f
C690 VTAIL.n10 VSUBS 0.015293f
C691 VTAIL.n11 VSUBS 0.026879f
C692 VTAIL.n12 VSUBS 0.014443f
C693 VTAIL.n13 VSUBS 0.034139f
C694 VTAIL.n14 VSUBS 0.015293f
C695 VTAIL.n15 VSUBS 0.026879f
C696 VTAIL.n16 VSUBS 0.014443f
C697 VTAIL.n17 VSUBS 0.034139f
C698 VTAIL.n18 VSUBS 0.015293f
C699 VTAIL.n19 VSUBS 0.026879f
C700 VTAIL.n20 VSUBS 0.014443f
C701 VTAIL.n21 VSUBS 0.034139f
C702 VTAIL.n22 VSUBS 0.015293f
C703 VTAIL.n23 VSUBS 0.026879f
C704 VTAIL.n24 VSUBS 0.014443f
C705 VTAIL.n25 VSUBS 0.025604f
C706 VTAIL.n26 VSUBS 0.021718f
C707 VTAIL.t15 VSUBS 0.073026f
C708 VTAIL.n27 VSUBS 0.182495f
C709 VTAIL.n28 VSUBS 1.60887f
C710 VTAIL.n29 VSUBS 0.014443f
C711 VTAIL.n30 VSUBS 0.015293f
C712 VTAIL.n31 VSUBS 0.034139f
C713 VTAIL.n32 VSUBS 0.034139f
C714 VTAIL.n33 VSUBS 0.015293f
C715 VTAIL.n34 VSUBS 0.014443f
C716 VTAIL.n35 VSUBS 0.026879f
C717 VTAIL.n36 VSUBS 0.026879f
C718 VTAIL.n37 VSUBS 0.014443f
C719 VTAIL.n38 VSUBS 0.015293f
C720 VTAIL.n39 VSUBS 0.034139f
C721 VTAIL.n40 VSUBS 0.034139f
C722 VTAIL.n41 VSUBS 0.015293f
C723 VTAIL.n42 VSUBS 0.014443f
C724 VTAIL.n43 VSUBS 0.026879f
C725 VTAIL.n44 VSUBS 0.026879f
C726 VTAIL.n45 VSUBS 0.014443f
C727 VTAIL.n46 VSUBS 0.015293f
C728 VTAIL.n47 VSUBS 0.034139f
C729 VTAIL.n48 VSUBS 0.034139f
C730 VTAIL.n49 VSUBS 0.015293f
C731 VTAIL.n50 VSUBS 0.014443f
C732 VTAIL.n51 VSUBS 0.026879f
C733 VTAIL.n52 VSUBS 0.026879f
C734 VTAIL.n53 VSUBS 0.014443f
C735 VTAIL.n54 VSUBS 0.015293f
C736 VTAIL.n55 VSUBS 0.034139f
C737 VTAIL.n56 VSUBS 0.034139f
C738 VTAIL.n57 VSUBS 0.015293f
C739 VTAIL.n58 VSUBS 0.014443f
C740 VTAIL.n59 VSUBS 0.026879f
C741 VTAIL.n60 VSUBS 0.026879f
C742 VTAIL.n61 VSUBS 0.014443f
C743 VTAIL.n62 VSUBS 0.015293f
C744 VTAIL.n63 VSUBS 0.034139f
C745 VTAIL.n64 VSUBS 0.034139f
C746 VTAIL.n65 VSUBS 0.015293f
C747 VTAIL.n66 VSUBS 0.014443f
C748 VTAIL.n67 VSUBS 0.026879f
C749 VTAIL.n68 VSUBS 0.026879f
C750 VTAIL.n69 VSUBS 0.014443f
C751 VTAIL.n70 VSUBS 0.014443f
C752 VTAIL.n71 VSUBS 0.015293f
C753 VTAIL.n72 VSUBS 0.034139f
C754 VTAIL.n73 VSUBS 0.034139f
C755 VTAIL.n74 VSUBS 0.080711f
C756 VTAIL.n75 VSUBS 0.014868f
C757 VTAIL.n76 VSUBS 0.014443f
C758 VTAIL.n77 VSUBS 0.069472f
C759 VTAIL.n78 VSUBS 0.040718f
C760 VTAIL.n79 VSUBS 0.122307f
C761 VTAIL.n80 VSUBS 0.028966f
C762 VTAIL.n81 VSUBS 0.026879f
C763 VTAIL.n82 VSUBS 0.014868f
C764 VTAIL.n83 VSUBS 0.034139f
C765 VTAIL.n84 VSUBS 0.015293f
C766 VTAIL.n85 VSUBS 0.026879f
C767 VTAIL.n86 VSUBS 0.014443f
C768 VTAIL.n87 VSUBS 0.034139f
C769 VTAIL.n88 VSUBS 0.015293f
C770 VTAIL.n89 VSUBS 0.026879f
C771 VTAIL.n90 VSUBS 0.014443f
C772 VTAIL.n91 VSUBS 0.034139f
C773 VTAIL.n92 VSUBS 0.015293f
C774 VTAIL.n93 VSUBS 0.026879f
C775 VTAIL.n94 VSUBS 0.014443f
C776 VTAIL.n95 VSUBS 0.034139f
C777 VTAIL.n96 VSUBS 0.015293f
C778 VTAIL.n97 VSUBS 0.026879f
C779 VTAIL.n98 VSUBS 0.014443f
C780 VTAIL.n99 VSUBS 0.034139f
C781 VTAIL.n100 VSUBS 0.015293f
C782 VTAIL.n101 VSUBS 0.026879f
C783 VTAIL.n102 VSUBS 0.014443f
C784 VTAIL.n103 VSUBS 0.025604f
C785 VTAIL.n104 VSUBS 0.021718f
C786 VTAIL.t4 VSUBS 0.073026f
C787 VTAIL.n105 VSUBS 0.182495f
C788 VTAIL.n106 VSUBS 1.60887f
C789 VTAIL.n107 VSUBS 0.014443f
C790 VTAIL.n108 VSUBS 0.015293f
C791 VTAIL.n109 VSUBS 0.034139f
C792 VTAIL.n110 VSUBS 0.034139f
C793 VTAIL.n111 VSUBS 0.015293f
C794 VTAIL.n112 VSUBS 0.014443f
C795 VTAIL.n113 VSUBS 0.026879f
C796 VTAIL.n114 VSUBS 0.026879f
C797 VTAIL.n115 VSUBS 0.014443f
C798 VTAIL.n116 VSUBS 0.015293f
C799 VTAIL.n117 VSUBS 0.034139f
C800 VTAIL.n118 VSUBS 0.034139f
C801 VTAIL.n119 VSUBS 0.015293f
C802 VTAIL.n120 VSUBS 0.014443f
C803 VTAIL.n121 VSUBS 0.026879f
C804 VTAIL.n122 VSUBS 0.026879f
C805 VTAIL.n123 VSUBS 0.014443f
C806 VTAIL.n124 VSUBS 0.015293f
C807 VTAIL.n125 VSUBS 0.034139f
C808 VTAIL.n126 VSUBS 0.034139f
C809 VTAIL.n127 VSUBS 0.015293f
C810 VTAIL.n128 VSUBS 0.014443f
C811 VTAIL.n129 VSUBS 0.026879f
C812 VTAIL.n130 VSUBS 0.026879f
C813 VTAIL.n131 VSUBS 0.014443f
C814 VTAIL.n132 VSUBS 0.015293f
C815 VTAIL.n133 VSUBS 0.034139f
C816 VTAIL.n134 VSUBS 0.034139f
C817 VTAIL.n135 VSUBS 0.015293f
C818 VTAIL.n136 VSUBS 0.014443f
C819 VTAIL.n137 VSUBS 0.026879f
C820 VTAIL.n138 VSUBS 0.026879f
C821 VTAIL.n139 VSUBS 0.014443f
C822 VTAIL.n140 VSUBS 0.015293f
C823 VTAIL.n141 VSUBS 0.034139f
C824 VTAIL.n142 VSUBS 0.034139f
C825 VTAIL.n143 VSUBS 0.015293f
C826 VTAIL.n144 VSUBS 0.014443f
C827 VTAIL.n145 VSUBS 0.026879f
C828 VTAIL.n146 VSUBS 0.026879f
C829 VTAIL.n147 VSUBS 0.014443f
C830 VTAIL.n148 VSUBS 0.014443f
C831 VTAIL.n149 VSUBS 0.015293f
C832 VTAIL.n150 VSUBS 0.034139f
C833 VTAIL.n151 VSUBS 0.034139f
C834 VTAIL.n152 VSUBS 0.080711f
C835 VTAIL.n153 VSUBS 0.014868f
C836 VTAIL.n154 VSUBS 0.014443f
C837 VTAIL.n155 VSUBS 0.069472f
C838 VTAIL.n156 VSUBS 0.040718f
C839 VTAIL.n157 VSUBS 0.122307f
C840 VTAIL.t3 VSUBS 0.299913f
C841 VTAIL.t0 VSUBS 0.299913f
C842 VTAIL.n158 VSUBS 2.28809f
C843 VTAIL.n159 VSUBS 0.706489f
C844 VTAIL.n160 VSUBS 0.028966f
C845 VTAIL.n161 VSUBS 0.026879f
C846 VTAIL.n162 VSUBS 0.014868f
C847 VTAIL.n163 VSUBS 0.034139f
C848 VTAIL.n164 VSUBS 0.015293f
C849 VTAIL.n165 VSUBS 0.026879f
C850 VTAIL.n166 VSUBS 0.014443f
C851 VTAIL.n167 VSUBS 0.034139f
C852 VTAIL.n168 VSUBS 0.015293f
C853 VTAIL.n169 VSUBS 0.026879f
C854 VTAIL.n170 VSUBS 0.014443f
C855 VTAIL.n171 VSUBS 0.034139f
C856 VTAIL.n172 VSUBS 0.015293f
C857 VTAIL.n173 VSUBS 0.026879f
C858 VTAIL.n174 VSUBS 0.014443f
C859 VTAIL.n175 VSUBS 0.034139f
C860 VTAIL.n176 VSUBS 0.015293f
C861 VTAIL.n177 VSUBS 0.026879f
C862 VTAIL.n178 VSUBS 0.014443f
C863 VTAIL.n179 VSUBS 0.034139f
C864 VTAIL.n180 VSUBS 0.015293f
C865 VTAIL.n181 VSUBS 0.026879f
C866 VTAIL.n182 VSUBS 0.014443f
C867 VTAIL.n183 VSUBS 0.025604f
C868 VTAIL.n184 VSUBS 0.021718f
C869 VTAIL.t1 VSUBS 0.073026f
C870 VTAIL.n185 VSUBS 0.182495f
C871 VTAIL.n186 VSUBS 1.60887f
C872 VTAIL.n187 VSUBS 0.014443f
C873 VTAIL.n188 VSUBS 0.015293f
C874 VTAIL.n189 VSUBS 0.034139f
C875 VTAIL.n190 VSUBS 0.034139f
C876 VTAIL.n191 VSUBS 0.015293f
C877 VTAIL.n192 VSUBS 0.014443f
C878 VTAIL.n193 VSUBS 0.026879f
C879 VTAIL.n194 VSUBS 0.026879f
C880 VTAIL.n195 VSUBS 0.014443f
C881 VTAIL.n196 VSUBS 0.015293f
C882 VTAIL.n197 VSUBS 0.034139f
C883 VTAIL.n198 VSUBS 0.034139f
C884 VTAIL.n199 VSUBS 0.015293f
C885 VTAIL.n200 VSUBS 0.014443f
C886 VTAIL.n201 VSUBS 0.026879f
C887 VTAIL.n202 VSUBS 0.026879f
C888 VTAIL.n203 VSUBS 0.014443f
C889 VTAIL.n204 VSUBS 0.015293f
C890 VTAIL.n205 VSUBS 0.034139f
C891 VTAIL.n206 VSUBS 0.034139f
C892 VTAIL.n207 VSUBS 0.015293f
C893 VTAIL.n208 VSUBS 0.014443f
C894 VTAIL.n209 VSUBS 0.026879f
C895 VTAIL.n210 VSUBS 0.026879f
C896 VTAIL.n211 VSUBS 0.014443f
C897 VTAIL.n212 VSUBS 0.015293f
C898 VTAIL.n213 VSUBS 0.034139f
C899 VTAIL.n214 VSUBS 0.034139f
C900 VTAIL.n215 VSUBS 0.015293f
C901 VTAIL.n216 VSUBS 0.014443f
C902 VTAIL.n217 VSUBS 0.026879f
C903 VTAIL.n218 VSUBS 0.026879f
C904 VTAIL.n219 VSUBS 0.014443f
C905 VTAIL.n220 VSUBS 0.015293f
C906 VTAIL.n221 VSUBS 0.034139f
C907 VTAIL.n222 VSUBS 0.034139f
C908 VTAIL.n223 VSUBS 0.015293f
C909 VTAIL.n224 VSUBS 0.014443f
C910 VTAIL.n225 VSUBS 0.026879f
C911 VTAIL.n226 VSUBS 0.026879f
C912 VTAIL.n227 VSUBS 0.014443f
C913 VTAIL.n228 VSUBS 0.014443f
C914 VTAIL.n229 VSUBS 0.015293f
C915 VTAIL.n230 VSUBS 0.034139f
C916 VTAIL.n231 VSUBS 0.034139f
C917 VTAIL.n232 VSUBS 0.080711f
C918 VTAIL.n233 VSUBS 0.014868f
C919 VTAIL.n234 VSUBS 0.014443f
C920 VTAIL.n235 VSUBS 0.069472f
C921 VTAIL.n236 VSUBS 0.040718f
C922 VTAIL.n237 VSUBS 1.55547f
C923 VTAIL.n238 VSUBS 0.028966f
C924 VTAIL.n239 VSUBS 0.026879f
C925 VTAIL.n240 VSUBS 0.014868f
C926 VTAIL.n241 VSUBS 0.034139f
C927 VTAIL.n242 VSUBS 0.014443f
C928 VTAIL.n243 VSUBS 0.015293f
C929 VTAIL.n244 VSUBS 0.026879f
C930 VTAIL.n245 VSUBS 0.014443f
C931 VTAIL.n246 VSUBS 0.034139f
C932 VTAIL.n247 VSUBS 0.015293f
C933 VTAIL.n248 VSUBS 0.026879f
C934 VTAIL.n249 VSUBS 0.014443f
C935 VTAIL.n250 VSUBS 0.034139f
C936 VTAIL.n251 VSUBS 0.015293f
C937 VTAIL.n252 VSUBS 0.026879f
C938 VTAIL.n253 VSUBS 0.014443f
C939 VTAIL.n254 VSUBS 0.034139f
C940 VTAIL.n255 VSUBS 0.015293f
C941 VTAIL.n256 VSUBS 0.026879f
C942 VTAIL.n257 VSUBS 0.014443f
C943 VTAIL.n258 VSUBS 0.034139f
C944 VTAIL.n259 VSUBS 0.015293f
C945 VTAIL.n260 VSUBS 0.026879f
C946 VTAIL.n261 VSUBS 0.014443f
C947 VTAIL.n262 VSUBS 0.025604f
C948 VTAIL.n263 VSUBS 0.021718f
C949 VTAIL.t10 VSUBS 0.073026f
C950 VTAIL.n264 VSUBS 0.182495f
C951 VTAIL.n265 VSUBS 1.60887f
C952 VTAIL.n266 VSUBS 0.014443f
C953 VTAIL.n267 VSUBS 0.015293f
C954 VTAIL.n268 VSUBS 0.034139f
C955 VTAIL.n269 VSUBS 0.034139f
C956 VTAIL.n270 VSUBS 0.015293f
C957 VTAIL.n271 VSUBS 0.014443f
C958 VTAIL.n272 VSUBS 0.026879f
C959 VTAIL.n273 VSUBS 0.026879f
C960 VTAIL.n274 VSUBS 0.014443f
C961 VTAIL.n275 VSUBS 0.015293f
C962 VTAIL.n276 VSUBS 0.034139f
C963 VTAIL.n277 VSUBS 0.034139f
C964 VTAIL.n278 VSUBS 0.015293f
C965 VTAIL.n279 VSUBS 0.014443f
C966 VTAIL.n280 VSUBS 0.026879f
C967 VTAIL.n281 VSUBS 0.026879f
C968 VTAIL.n282 VSUBS 0.014443f
C969 VTAIL.n283 VSUBS 0.015293f
C970 VTAIL.n284 VSUBS 0.034139f
C971 VTAIL.n285 VSUBS 0.034139f
C972 VTAIL.n286 VSUBS 0.015293f
C973 VTAIL.n287 VSUBS 0.014443f
C974 VTAIL.n288 VSUBS 0.026879f
C975 VTAIL.n289 VSUBS 0.026879f
C976 VTAIL.n290 VSUBS 0.014443f
C977 VTAIL.n291 VSUBS 0.015293f
C978 VTAIL.n292 VSUBS 0.034139f
C979 VTAIL.n293 VSUBS 0.034139f
C980 VTAIL.n294 VSUBS 0.015293f
C981 VTAIL.n295 VSUBS 0.014443f
C982 VTAIL.n296 VSUBS 0.026879f
C983 VTAIL.n297 VSUBS 0.026879f
C984 VTAIL.n298 VSUBS 0.014443f
C985 VTAIL.n299 VSUBS 0.015293f
C986 VTAIL.n300 VSUBS 0.034139f
C987 VTAIL.n301 VSUBS 0.034139f
C988 VTAIL.n302 VSUBS 0.015293f
C989 VTAIL.n303 VSUBS 0.014443f
C990 VTAIL.n304 VSUBS 0.026879f
C991 VTAIL.n305 VSUBS 0.026879f
C992 VTAIL.n306 VSUBS 0.014443f
C993 VTAIL.n307 VSUBS 0.015293f
C994 VTAIL.n308 VSUBS 0.034139f
C995 VTAIL.n309 VSUBS 0.034139f
C996 VTAIL.n310 VSUBS 0.080711f
C997 VTAIL.n311 VSUBS 0.014868f
C998 VTAIL.n312 VSUBS 0.014443f
C999 VTAIL.n313 VSUBS 0.069472f
C1000 VTAIL.n314 VSUBS 0.040718f
C1001 VTAIL.n315 VSUBS 1.55547f
C1002 VTAIL.t8 VSUBS 0.299913f
C1003 VTAIL.t14 VSUBS 0.299913f
C1004 VTAIL.n316 VSUBS 2.28811f
C1005 VTAIL.n317 VSUBS 0.706475f
C1006 VTAIL.n318 VSUBS 0.028966f
C1007 VTAIL.n319 VSUBS 0.026879f
C1008 VTAIL.n320 VSUBS 0.014868f
C1009 VTAIL.n321 VSUBS 0.034139f
C1010 VTAIL.n322 VSUBS 0.014443f
C1011 VTAIL.n323 VSUBS 0.015293f
C1012 VTAIL.n324 VSUBS 0.026879f
C1013 VTAIL.n325 VSUBS 0.014443f
C1014 VTAIL.n326 VSUBS 0.034139f
C1015 VTAIL.n327 VSUBS 0.015293f
C1016 VTAIL.n328 VSUBS 0.026879f
C1017 VTAIL.n329 VSUBS 0.014443f
C1018 VTAIL.n330 VSUBS 0.034139f
C1019 VTAIL.n331 VSUBS 0.015293f
C1020 VTAIL.n332 VSUBS 0.026879f
C1021 VTAIL.n333 VSUBS 0.014443f
C1022 VTAIL.n334 VSUBS 0.034139f
C1023 VTAIL.n335 VSUBS 0.015293f
C1024 VTAIL.n336 VSUBS 0.026879f
C1025 VTAIL.n337 VSUBS 0.014443f
C1026 VTAIL.n338 VSUBS 0.034139f
C1027 VTAIL.n339 VSUBS 0.015293f
C1028 VTAIL.n340 VSUBS 0.026879f
C1029 VTAIL.n341 VSUBS 0.014443f
C1030 VTAIL.n342 VSUBS 0.025604f
C1031 VTAIL.n343 VSUBS 0.021718f
C1032 VTAIL.t13 VSUBS 0.073026f
C1033 VTAIL.n344 VSUBS 0.182495f
C1034 VTAIL.n345 VSUBS 1.60887f
C1035 VTAIL.n346 VSUBS 0.014443f
C1036 VTAIL.n347 VSUBS 0.015293f
C1037 VTAIL.n348 VSUBS 0.034139f
C1038 VTAIL.n349 VSUBS 0.034139f
C1039 VTAIL.n350 VSUBS 0.015293f
C1040 VTAIL.n351 VSUBS 0.014443f
C1041 VTAIL.n352 VSUBS 0.026879f
C1042 VTAIL.n353 VSUBS 0.026879f
C1043 VTAIL.n354 VSUBS 0.014443f
C1044 VTAIL.n355 VSUBS 0.015293f
C1045 VTAIL.n356 VSUBS 0.034139f
C1046 VTAIL.n357 VSUBS 0.034139f
C1047 VTAIL.n358 VSUBS 0.015293f
C1048 VTAIL.n359 VSUBS 0.014443f
C1049 VTAIL.n360 VSUBS 0.026879f
C1050 VTAIL.n361 VSUBS 0.026879f
C1051 VTAIL.n362 VSUBS 0.014443f
C1052 VTAIL.n363 VSUBS 0.015293f
C1053 VTAIL.n364 VSUBS 0.034139f
C1054 VTAIL.n365 VSUBS 0.034139f
C1055 VTAIL.n366 VSUBS 0.015293f
C1056 VTAIL.n367 VSUBS 0.014443f
C1057 VTAIL.n368 VSUBS 0.026879f
C1058 VTAIL.n369 VSUBS 0.026879f
C1059 VTAIL.n370 VSUBS 0.014443f
C1060 VTAIL.n371 VSUBS 0.015293f
C1061 VTAIL.n372 VSUBS 0.034139f
C1062 VTAIL.n373 VSUBS 0.034139f
C1063 VTAIL.n374 VSUBS 0.015293f
C1064 VTAIL.n375 VSUBS 0.014443f
C1065 VTAIL.n376 VSUBS 0.026879f
C1066 VTAIL.n377 VSUBS 0.026879f
C1067 VTAIL.n378 VSUBS 0.014443f
C1068 VTAIL.n379 VSUBS 0.015293f
C1069 VTAIL.n380 VSUBS 0.034139f
C1070 VTAIL.n381 VSUBS 0.034139f
C1071 VTAIL.n382 VSUBS 0.015293f
C1072 VTAIL.n383 VSUBS 0.014443f
C1073 VTAIL.n384 VSUBS 0.026879f
C1074 VTAIL.n385 VSUBS 0.026879f
C1075 VTAIL.n386 VSUBS 0.014443f
C1076 VTAIL.n387 VSUBS 0.015293f
C1077 VTAIL.n388 VSUBS 0.034139f
C1078 VTAIL.n389 VSUBS 0.034139f
C1079 VTAIL.n390 VSUBS 0.080711f
C1080 VTAIL.n391 VSUBS 0.014868f
C1081 VTAIL.n392 VSUBS 0.014443f
C1082 VTAIL.n393 VSUBS 0.069472f
C1083 VTAIL.n394 VSUBS 0.040718f
C1084 VTAIL.n395 VSUBS 0.122307f
C1085 VTAIL.n396 VSUBS 0.028966f
C1086 VTAIL.n397 VSUBS 0.026879f
C1087 VTAIL.n398 VSUBS 0.014868f
C1088 VTAIL.n399 VSUBS 0.034139f
C1089 VTAIL.n400 VSUBS 0.014443f
C1090 VTAIL.n401 VSUBS 0.015293f
C1091 VTAIL.n402 VSUBS 0.026879f
C1092 VTAIL.n403 VSUBS 0.014443f
C1093 VTAIL.n404 VSUBS 0.034139f
C1094 VTAIL.n405 VSUBS 0.015293f
C1095 VTAIL.n406 VSUBS 0.026879f
C1096 VTAIL.n407 VSUBS 0.014443f
C1097 VTAIL.n408 VSUBS 0.034139f
C1098 VTAIL.n409 VSUBS 0.015293f
C1099 VTAIL.n410 VSUBS 0.026879f
C1100 VTAIL.n411 VSUBS 0.014443f
C1101 VTAIL.n412 VSUBS 0.034139f
C1102 VTAIL.n413 VSUBS 0.015293f
C1103 VTAIL.n414 VSUBS 0.026879f
C1104 VTAIL.n415 VSUBS 0.014443f
C1105 VTAIL.n416 VSUBS 0.034139f
C1106 VTAIL.n417 VSUBS 0.015293f
C1107 VTAIL.n418 VSUBS 0.026879f
C1108 VTAIL.n419 VSUBS 0.014443f
C1109 VTAIL.n420 VSUBS 0.025604f
C1110 VTAIL.n421 VSUBS 0.021718f
C1111 VTAIL.t6 VSUBS 0.073026f
C1112 VTAIL.n422 VSUBS 0.182495f
C1113 VTAIL.n423 VSUBS 1.60887f
C1114 VTAIL.n424 VSUBS 0.014443f
C1115 VTAIL.n425 VSUBS 0.015293f
C1116 VTAIL.n426 VSUBS 0.034139f
C1117 VTAIL.n427 VSUBS 0.034139f
C1118 VTAIL.n428 VSUBS 0.015293f
C1119 VTAIL.n429 VSUBS 0.014443f
C1120 VTAIL.n430 VSUBS 0.026879f
C1121 VTAIL.n431 VSUBS 0.026879f
C1122 VTAIL.n432 VSUBS 0.014443f
C1123 VTAIL.n433 VSUBS 0.015293f
C1124 VTAIL.n434 VSUBS 0.034139f
C1125 VTAIL.n435 VSUBS 0.034139f
C1126 VTAIL.n436 VSUBS 0.015293f
C1127 VTAIL.n437 VSUBS 0.014443f
C1128 VTAIL.n438 VSUBS 0.026879f
C1129 VTAIL.n439 VSUBS 0.026879f
C1130 VTAIL.n440 VSUBS 0.014443f
C1131 VTAIL.n441 VSUBS 0.015293f
C1132 VTAIL.n442 VSUBS 0.034139f
C1133 VTAIL.n443 VSUBS 0.034139f
C1134 VTAIL.n444 VSUBS 0.015293f
C1135 VTAIL.n445 VSUBS 0.014443f
C1136 VTAIL.n446 VSUBS 0.026879f
C1137 VTAIL.n447 VSUBS 0.026879f
C1138 VTAIL.n448 VSUBS 0.014443f
C1139 VTAIL.n449 VSUBS 0.015293f
C1140 VTAIL.n450 VSUBS 0.034139f
C1141 VTAIL.n451 VSUBS 0.034139f
C1142 VTAIL.n452 VSUBS 0.015293f
C1143 VTAIL.n453 VSUBS 0.014443f
C1144 VTAIL.n454 VSUBS 0.026879f
C1145 VTAIL.n455 VSUBS 0.026879f
C1146 VTAIL.n456 VSUBS 0.014443f
C1147 VTAIL.n457 VSUBS 0.015293f
C1148 VTAIL.n458 VSUBS 0.034139f
C1149 VTAIL.n459 VSUBS 0.034139f
C1150 VTAIL.n460 VSUBS 0.015293f
C1151 VTAIL.n461 VSUBS 0.014443f
C1152 VTAIL.n462 VSUBS 0.026879f
C1153 VTAIL.n463 VSUBS 0.026879f
C1154 VTAIL.n464 VSUBS 0.014443f
C1155 VTAIL.n465 VSUBS 0.015293f
C1156 VTAIL.n466 VSUBS 0.034139f
C1157 VTAIL.n467 VSUBS 0.034139f
C1158 VTAIL.n468 VSUBS 0.080711f
C1159 VTAIL.n469 VSUBS 0.014868f
C1160 VTAIL.n470 VSUBS 0.014443f
C1161 VTAIL.n471 VSUBS 0.069472f
C1162 VTAIL.n472 VSUBS 0.040718f
C1163 VTAIL.n473 VSUBS 0.122307f
C1164 VTAIL.t7 VSUBS 0.299913f
C1165 VTAIL.t2 VSUBS 0.299913f
C1166 VTAIL.n474 VSUBS 2.28811f
C1167 VTAIL.n475 VSUBS 0.706475f
C1168 VTAIL.n476 VSUBS 0.028966f
C1169 VTAIL.n477 VSUBS 0.026879f
C1170 VTAIL.n478 VSUBS 0.014868f
C1171 VTAIL.n479 VSUBS 0.034139f
C1172 VTAIL.n480 VSUBS 0.014443f
C1173 VTAIL.n481 VSUBS 0.015293f
C1174 VTAIL.n482 VSUBS 0.026879f
C1175 VTAIL.n483 VSUBS 0.014443f
C1176 VTAIL.n484 VSUBS 0.034139f
C1177 VTAIL.n485 VSUBS 0.015293f
C1178 VTAIL.n486 VSUBS 0.026879f
C1179 VTAIL.n487 VSUBS 0.014443f
C1180 VTAIL.n488 VSUBS 0.034139f
C1181 VTAIL.n489 VSUBS 0.015293f
C1182 VTAIL.n490 VSUBS 0.026879f
C1183 VTAIL.n491 VSUBS 0.014443f
C1184 VTAIL.n492 VSUBS 0.034139f
C1185 VTAIL.n493 VSUBS 0.015293f
C1186 VTAIL.n494 VSUBS 0.026879f
C1187 VTAIL.n495 VSUBS 0.014443f
C1188 VTAIL.n496 VSUBS 0.034139f
C1189 VTAIL.n497 VSUBS 0.015293f
C1190 VTAIL.n498 VSUBS 0.026879f
C1191 VTAIL.n499 VSUBS 0.014443f
C1192 VTAIL.n500 VSUBS 0.025604f
C1193 VTAIL.n501 VSUBS 0.021718f
C1194 VTAIL.t5 VSUBS 0.073026f
C1195 VTAIL.n502 VSUBS 0.182495f
C1196 VTAIL.n503 VSUBS 1.60887f
C1197 VTAIL.n504 VSUBS 0.014443f
C1198 VTAIL.n505 VSUBS 0.015293f
C1199 VTAIL.n506 VSUBS 0.034139f
C1200 VTAIL.n507 VSUBS 0.034139f
C1201 VTAIL.n508 VSUBS 0.015293f
C1202 VTAIL.n509 VSUBS 0.014443f
C1203 VTAIL.n510 VSUBS 0.026879f
C1204 VTAIL.n511 VSUBS 0.026879f
C1205 VTAIL.n512 VSUBS 0.014443f
C1206 VTAIL.n513 VSUBS 0.015293f
C1207 VTAIL.n514 VSUBS 0.034139f
C1208 VTAIL.n515 VSUBS 0.034139f
C1209 VTAIL.n516 VSUBS 0.015293f
C1210 VTAIL.n517 VSUBS 0.014443f
C1211 VTAIL.n518 VSUBS 0.026879f
C1212 VTAIL.n519 VSUBS 0.026879f
C1213 VTAIL.n520 VSUBS 0.014443f
C1214 VTAIL.n521 VSUBS 0.015293f
C1215 VTAIL.n522 VSUBS 0.034139f
C1216 VTAIL.n523 VSUBS 0.034139f
C1217 VTAIL.n524 VSUBS 0.015293f
C1218 VTAIL.n525 VSUBS 0.014443f
C1219 VTAIL.n526 VSUBS 0.026879f
C1220 VTAIL.n527 VSUBS 0.026879f
C1221 VTAIL.n528 VSUBS 0.014443f
C1222 VTAIL.n529 VSUBS 0.015293f
C1223 VTAIL.n530 VSUBS 0.034139f
C1224 VTAIL.n531 VSUBS 0.034139f
C1225 VTAIL.n532 VSUBS 0.015293f
C1226 VTAIL.n533 VSUBS 0.014443f
C1227 VTAIL.n534 VSUBS 0.026879f
C1228 VTAIL.n535 VSUBS 0.026879f
C1229 VTAIL.n536 VSUBS 0.014443f
C1230 VTAIL.n537 VSUBS 0.015293f
C1231 VTAIL.n538 VSUBS 0.034139f
C1232 VTAIL.n539 VSUBS 0.034139f
C1233 VTAIL.n540 VSUBS 0.015293f
C1234 VTAIL.n541 VSUBS 0.014443f
C1235 VTAIL.n542 VSUBS 0.026879f
C1236 VTAIL.n543 VSUBS 0.026879f
C1237 VTAIL.n544 VSUBS 0.014443f
C1238 VTAIL.n545 VSUBS 0.015293f
C1239 VTAIL.n546 VSUBS 0.034139f
C1240 VTAIL.n547 VSUBS 0.034139f
C1241 VTAIL.n548 VSUBS 0.080711f
C1242 VTAIL.n549 VSUBS 0.014868f
C1243 VTAIL.n550 VSUBS 0.014443f
C1244 VTAIL.n551 VSUBS 0.069472f
C1245 VTAIL.n552 VSUBS 0.040718f
C1246 VTAIL.n553 VSUBS 1.55547f
C1247 VTAIL.n554 VSUBS 0.028966f
C1248 VTAIL.n555 VSUBS 0.026879f
C1249 VTAIL.n556 VSUBS 0.014868f
C1250 VTAIL.n557 VSUBS 0.034139f
C1251 VTAIL.n558 VSUBS 0.015293f
C1252 VTAIL.n559 VSUBS 0.026879f
C1253 VTAIL.n560 VSUBS 0.014443f
C1254 VTAIL.n561 VSUBS 0.034139f
C1255 VTAIL.n562 VSUBS 0.015293f
C1256 VTAIL.n563 VSUBS 0.026879f
C1257 VTAIL.n564 VSUBS 0.014443f
C1258 VTAIL.n565 VSUBS 0.034139f
C1259 VTAIL.n566 VSUBS 0.015293f
C1260 VTAIL.n567 VSUBS 0.026879f
C1261 VTAIL.n568 VSUBS 0.014443f
C1262 VTAIL.n569 VSUBS 0.034139f
C1263 VTAIL.n570 VSUBS 0.015293f
C1264 VTAIL.n571 VSUBS 0.026879f
C1265 VTAIL.n572 VSUBS 0.014443f
C1266 VTAIL.n573 VSUBS 0.034139f
C1267 VTAIL.n574 VSUBS 0.015293f
C1268 VTAIL.n575 VSUBS 0.026879f
C1269 VTAIL.n576 VSUBS 0.014443f
C1270 VTAIL.n577 VSUBS 0.025604f
C1271 VTAIL.n578 VSUBS 0.021718f
C1272 VTAIL.t9 VSUBS 0.073026f
C1273 VTAIL.n579 VSUBS 0.182495f
C1274 VTAIL.n580 VSUBS 1.60887f
C1275 VTAIL.n581 VSUBS 0.014443f
C1276 VTAIL.n582 VSUBS 0.015293f
C1277 VTAIL.n583 VSUBS 0.034139f
C1278 VTAIL.n584 VSUBS 0.034139f
C1279 VTAIL.n585 VSUBS 0.015293f
C1280 VTAIL.n586 VSUBS 0.014443f
C1281 VTAIL.n587 VSUBS 0.026879f
C1282 VTAIL.n588 VSUBS 0.026879f
C1283 VTAIL.n589 VSUBS 0.014443f
C1284 VTAIL.n590 VSUBS 0.015293f
C1285 VTAIL.n591 VSUBS 0.034139f
C1286 VTAIL.n592 VSUBS 0.034139f
C1287 VTAIL.n593 VSUBS 0.015293f
C1288 VTAIL.n594 VSUBS 0.014443f
C1289 VTAIL.n595 VSUBS 0.026879f
C1290 VTAIL.n596 VSUBS 0.026879f
C1291 VTAIL.n597 VSUBS 0.014443f
C1292 VTAIL.n598 VSUBS 0.015293f
C1293 VTAIL.n599 VSUBS 0.034139f
C1294 VTAIL.n600 VSUBS 0.034139f
C1295 VTAIL.n601 VSUBS 0.015293f
C1296 VTAIL.n602 VSUBS 0.014443f
C1297 VTAIL.n603 VSUBS 0.026879f
C1298 VTAIL.n604 VSUBS 0.026879f
C1299 VTAIL.n605 VSUBS 0.014443f
C1300 VTAIL.n606 VSUBS 0.015293f
C1301 VTAIL.n607 VSUBS 0.034139f
C1302 VTAIL.n608 VSUBS 0.034139f
C1303 VTAIL.n609 VSUBS 0.015293f
C1304 VTAIL.n610 VSUBS 0.014443f
C1305 VTAIL.n611 VSUBS 0.026879f
C1306 VTAIL.n612 VSUBS 0.026879f
C1307 VTAIL.n613 VSUBS 0.014443f
C1308 VTAIL.n614 VSUBS 0.015293f
C1309 VTAIL.n615 VSUBS 0.034139f
C1310 VTAIL.n616 VSUBS 0.034139f
C1311 VTAIL.n617 VSUBS 0.015293f
C1312 VTAIL.n618 VSUBS 0.014443f
C1313 VTAIL.n619 VSUBS 0.026879f
C1314 VTAIL.n620 VSUBS 0.026879f
C1315 VTAIL.n621 VSUBS 0.014443f
C1316 VTAIL.n622 VSUBS 0.014443f
C1317 VTAIL.n623 VSUBS 0.015293f
C1318 VTAIL.n624 VSUBS 0.034139f
C1319 VTAIL.n625 VSUBS 0.034139f
C1320 VTAIL.n626 VSUBS 0.080711f
C1321 VTAIL.n627 VSUBS 0.014868f
C1322 VTAIL.n628 VSUBS 0.014443f
C1323 VTAIL.n629 VSUBS 0.069472f
C1324 VTAIL.n630 VSUBS 0.040718f
C1325 VTAIL.n631 VSUBS 1.55043f
C1326 VN.n0 VSUBS 0.21155f
C1327 VN.t7 VSUBS 1.02616f
C1328 VN.n1 VSUBS 0.39331f
C1329 VN.t0 VSUBS 1.01255f
C1330 VN.n2 VSUBS 0.407999f
C1331 VN.t3 VSUBS 1.01255f
C1332 VN.n3 VSUBS 0.407999f
C1333 VN.t5 VSUBS 1.02111f
C1334 VN.n4 VSUBS 0.397884f
C1335 VN.n5 VSUBS 0.048848f
C1336 VN.n6 VSUBS 0.21155f
C1337 VN.t6 VSUBS 1.02111f
C1338 VN.t2 VSUBS 1.01255f
C1339 VN.t4 VSUBS 1.02616f
C1340 VN.n7 VSUBS 0.39331f
C1341 VN.n8 VSUBS 0.407999f
C1342 VN.t1 VSUBS 1.01255f
C1343 VN.n9 VSUBS 0.407999f
C1344 VN.n10 VSUBS 0.397884f
C1345 VN.n11 VSUBS 2.67912f
.ends

