* NGSPICE file created from diff_pair_sample_0576.ext - technology: sky130A

.subckt diff_pair_sample_0576 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t4 VP.t0 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=1.63515 ps=10.24 w=9.91 l=3.43
X1 VDD2.t3 VN.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.63515 pd=10.24 as=3.8649 ps=20.6 w=9.91 l=3.43
X2 VDD1.t3 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.63515 pd=10.24 as=3.8649 ps=20.6 w=9.91 l=3.43
X3 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=0 ps=0 w=9.91 l=3.43
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=0 ps=0 w=9.91 l=3.43
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=0 ps=0 w=9.91 l=3.43
X6 VTAIL.t6 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=1.63515 ps=10.24 w=9.91 l=3.43
X7 VDD2.t1 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.63515 pd=10.24 as=3.8649 ps=20.6 w=9.91 l=3.43
X8 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=1.63515 ps=10.24 w=9.91 l=3.43
X9 VDD1.t2 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.63515 pd=10.24 as=3.8649 ps=20.6 w=9.91 l=3.43
X10 VTAIL.t1 VP.t3 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=1.63515 ps=10.24 w=9.91 l=3.43
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8649 pd=20.6 as=0 ps=0 w=9.91 l=3.43
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n5 VP.t0 103.715
R9 VP.n5 VP.t2 102.513
R10 VP.n7 VP.n6 83.706
R11 VP.n20 VP.n0 83.706
R12 VP.n6 VP.t3 69.6305
R13 VP.n0 VP.t1 69.6305
R14 VP.n12 VP.n2 56.5193
R15 VP.n7 VP.n5 49.5214
R16 VP.n10 VP.n4 24.4675
R17 VP.n11 VP.n10 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n16 VP.n2 24.4675
R20 VP.n17 VP.n16 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n6 VP.n4 6.36192
R23 VP.n18 VP.n0 6.36192
R24 VP.n8 VP.n7 0.354971
R25 VP.n20 VP.n19 0.354971
R26 VP VP.n20 0.26696
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VDD1 VDD1.n1 104.177
R35 VDD1 VDD1.n0 61.7286
R36 VDD1.n0 VDD1.t0 1.99848
R37 VDD1.n0 VDD1.t2 1.99848
R38 VDD1.n1 VDD1.t1 1.99848
R39 VDD1.n1 VDD1.t3 1.99848
R40 VTAIL.n426 VTAIL.n378 289.615
R41 VTAIL.n48 VTAIL.n0 289.615
R42 VTAIL.n102 VTAIL.n54 289.615
R43 VTAIL.n156 VTAIL.n108 289.615
R44 VTAIL.n372 VTAIL.n324 289.615
R45 VTAIL.n318 VTAIL.n270 289.615
R46 VTAIL.n264 VTAIL.n216 289.615
R47 VTAIL.n210 VTAIL.n162 289.615
R48 VTAIL.n394 VTAIL.n393 185
R49 VTAIL.n399 VTAIL.n398 185
R50 VTAIL.n401 VTAIL.n400 185
R51 VTAIL.n390 VTAIL.n389 185
R52 VTAIL.n407 VTAIL.n406 185
R53 VTAIL.n409 VTAIL.n408 185
R54 VTAIL.n386 VTAIL.n385 185
R55 VTAIL.n416 VTAIL.n415 185
R56 VTAIL.n417 VTAIL.n384 185
R57 VTAIL.n419 VTAIL.n418 185
R58 VTAIL.n382 VTAIL.n381 185
R59 VTAIL.n425 VTAIL.n424 185
R60 VTAIL.n427 VTAIL.n426 185
R61 VTAIL.n16 VTAIL.n15 185
R62 VTAIL.n21 VTAIL.n20 185
R63 VTAIL.n23 VTAIL.n22 185
R64 VTAIL.n12 VTAIL.n11 185
R65 VTAIL.n29 VTAIL.n28 185
R66 VTAIL.n31 VTAIL.n30 185
R67 VTAIL.n8 VTAIL.n7 185
R68 VTAIL.n38 VTAIL.n37 185
R69 VTAIL.n39 VTAIL.n6 185
R70 VTAIL.n41 VTAIL.n40 185
R71 VTAIL.n4 VTAIL.n3 185
R72 VTAIL.n47 VTAIL.n46 185
R73 VTAIL.n49 VTAIL.n48 185
R74 VTAIL.n70 VTAIL.n69 185
R75 VTAIL.n75 VTAIL.n74 185
R76 VTAIL.n77 VTAIL.n76 185
R77 VTAIL.n66 VTAIL.n65 185
R78 VTAIL.n83 VTAIL.n82 185
R79 VTAIL.n85 VTAIL.n84 185
R80 VTAIL.n62 VTAIL.n61 185
R81 VTAIL.n92 VTAIL.n91 185
R82 VTAIL.n93 VTAIL.n60 185
R83 VTAIL.n95 VTAIL.n94 185
R84 VTAIL.n58 VTAIL.n57 185
R85 VTAIL.n101 VTAIL.n100 185
R86 VTAIL.n103 VTAIL.n102 185
R87 VTAIL.n124 VTAIL.n123 185
R88 VTAIL.n129 VTAIL.n128 185
R89 VTAIL.n131 VTAIL.n130 185
R90 VTAIL.n120 VTAIL.n119 185
R91 VTAIL.n137 VTAIL.n136 185
R92 VTAIL.n139 VTAIL.n138 185
R93 VTAIL.n116 VTAIL.n115 185
R94 VTAIL.n146 VTAIL.n145 185
R95 VTAIL.n147 VTAIL.n114 185
R96 VTAIL.n149 VTAIL.n148 185
R97 VTAIL.n112 VTAIL.n111 185
R98 VTAIL.n155 VTAIL.n154 185
R99 VTAIL.n157 VTAIL.n156 185
R100 VTAIL.n373 VTAIL.n372 185
R101 VTAIL.n371 VTAIL.n370 185
R102 VTAIL.n328 VTAIL.n327 185
R103 VTAIL.n365 VTAIL.n364 185
R104 VTAIL.n363 VTAIL.n330 185
R105 VTAIL.n362 VTAIL.n361 185
R106 VTAIL.n333 VTAIL.n331 185
R107 VTAIL.n356 VTAIL.n355 185
R108 VTAIL.n354 VTAIL.n353 185
R109 VTAIL.n337 VTAIL.n336 185
R110 VTAIL.n348 VTAIL.n347 185
R111 VTAIL.n346 VTAIL.n345 185
R112 VTAIL.n341 VTAIL.n340 185
R113 VTAIL.n319 VTAIL.n318 185
R114 VTAIL.n317 VTAIL.n316 185
R115 VTAIL.n274 VTAIL.n273 185
R116 VTAIL.n311 VTAIL.n310 185
R117 VTAIL.n309 VTAIL.n276 185
R118 VTAIL.n308 VTAIL.n307 185
R119 VTAIL.n279 VTAIL.n277 185
R120 VTAIL.n302 VTAIL.n301 185
R121 VTAIL.n300 VTAIL.n299 185
R122 VTAIL.n283 VTAIL.n282 185
R123 VTAIL.n294 VTAIL.n293 185
R124 VTAIL.n292 VTAIL.n291 185
R125 VTAIL.n287 VTAIL.n286 185
R126 VTAIL.n265 VTAIL.n264 185
R127 VTAIL.n263 VTAIL.n262 185
R128 VTAIL.n220 VTAIL.n219 185
R129 VTAIL.n257 VTAIL.n256 185
R130 VTAIL.n255 VTAIL.n222 185
R131 VTAIL.n254 VTAIL.n253 185
R132 VTAIL.n225 VTAIL.n223 185
R133 VTAIL.n248 VTAIL.n247 185
R134 VTAIL.n246 VTAIL.n245 185
R135 VTAIL.n229 VTAIL.n228 185
R136 VTAIL.n240 VTAIL.n239 185
R137 VTAIL.n238 VTAIL.n237 185
R138 VTAIL.n233 VTAIL.n232 185
R139 VTAIL.n211 VTAIL.n210 185
R140 VTAIL.n209 VTAIL.n208 185
R141 VTAIL.n166 VTAIL.n165 185
R142 VTAIL.n203 VTAIL.n202 185
R143 VTAIL.n201 VTAIL.n168 185
R144 VTAIL.n200 VTAIL.n199 185
R145 VTAIL.n171 VTAIL.n169 185
R146 VTAIL.n194 VTAIL.n193 185
R147 VTAIL.n192 VTAIL.n191 185
R148 VTAIL.n175 VTAIL.n174 185
R149 VTAIL.n186 VTAIL.n185 185
R150 VTAIL.n184 VTAIL.n183 185
R151 VTAIL.n179 VTAIL.n178 185
R152 VTAIL.n395 VTAIL.t7 149.524
R153 VTAIL.n17 VTAIL.t0 149.524
R154 VTAIL.n71 VTAIL.t3 149.524
R155 VTAIL.n125 VTAIL.t1 149.524
R156 VTAIL.n342 VTAIL.t2 149.524
R157 VTAIL.n288 VTAIL.t4 149.524
R158 VTAIL.n234 VTAIL.t5 149.524
R159 VTAIL.n180 VTAIL.t6 149.524
R160 VTAIL.n399 VTAIL.n393 104.615
R161 VTAIL.n400 VTAIL.n399 104.615
R162 VTAIL.n400 VTAIL.n389 104.615
R163 VTAIL.n407 VTAIL.n389 104.615
R164 VTAIL.n408 VTAIL.n407 104.615
R165 VTAIL.n408 VTAIL.n385 104.615
R166 VTAIL.n416 VTAIL.n385 104.615
R167 VTAIL.n417 VTAIL.n416 104.615
R168 VTAIL.n418 VTAIL.n417 104.615
R169 VTAIL.n418 VTAIL.n381 104.615
R170 VTAIL.n425 VTAIL.n381 104.615
R171 VTAIL.n426 VTAIL.n425 104.615
R172 VTAIL.n21 VTAIL.n15 104.615
R173 VTAIL.n22 VTAIL.n21 104.615
R174 VTAIL.n22 VTAIL.n11 104.615
R175 VTAIL.n29 VTAIL.n11 104.615
R176 VTAIL.n30 VTAIL.n29 104.615
R177 VTAIL.n30 VTAIL.n7 104.615
R178 VTAIL.n38 VTAIL.n7 104.615
R179 VTAIL.n39 VTAIL.n38 104.615
R180 VTAIL.n40 VTAIL.n39 104.615
R181 VTAIL.n40 VTAIL.n3 104.615
R182 VTAIL.n47 VTAIL.n3 104.615
R183 VTAIL.n48 VTAIL.n47 104.615
R184 VTAIL.n75 VTAIL.n69 104.615
R185 VTAIL.n76 VTAIL.n75 104.615
R186 VTAIL.n76 VTAIL.n65 104.615
R187 VTAIL.n83 VTAIL.n65 104.615
R188 VTAIL.n84 VTAIL.n83 104.615
R189 VTAIL.n84 VTAIL.n61 104.615
R190 VTAIL.n92 VTAIL.n61 104.615
R191 VTAIL.n93 VTAIL.n92 104.615
R192 VTAIL.n94 VTAIL.n93 104.615
R193 VTAIL.n94 VTAIL.n57 104.615
R194 VTAIL.n101 VTAIL.n57 104.615
R195 VTAIL.n102 VTAIL.n101 104.615
R196 VTAIL.n129 VTAIL.n123 104.615
R197 VTAIL.n130 VTAIL.n129 104.615
R198 VTAIL.n130 VTAIL.n119 104.615
R199 VTAIL.n137 VTAIL.n119 104.615
R200 VTAIL.n138 VTAIL.n137 104.615
R201 VTAIL.n138 VTAIL.n115 104.615
R202 VTAIL.n146 VTAIL.n115 104.615
R203 VTAIL.n147 VTAIL.n146 104.615
R204 VTAIL.n148 VTAIL.n147 104.615
R205 VTAIL.n148 VTAIL.n111 104.615
R206 VTAIL.n155 VTAIL.n111 104.615
R207 VTAIL.n156 VTAIL.n155 104.615
R208 VTAIL.n372 VTAIL.n371 104.615
R209 VTAIL.n371 VTAIL.n327 104.615
R210 VTAIL.n364 VTAIL.n327 104.615
R211 VTAIL.n364 VTAIL.n363 104.615
R212 VTAIL.n363 VTAIL.n362 104.615
R213 VTAIL.n362 VTAIL.n331 104.615
R214 VTAIL.n355 VTAIL.n331 104.615
R215 VTAIL.n355 VTAIL.n354 104.615
R216 VTAIL.n354 VTAIL.n336 104.615
R217 VTAIL.n347 VTAIL.n336 104.615
R218 VTAIL.n347 VTAIL.n346 104.615
R219 VTAIL.n346 VTAIL.n340 104.615
R220 VTAIL.n318 VTAIL.n317 104.615
R221 VTAIL.n317 VTAIL.n273 104.615
R222 VTAIL.n310 VTAIL.n273 104.615
R223 VTAIL.n310 VTAIL.n309 104.615
R224 VTAIL.n309 VTAIL.n308 104.615
R225 VTAIL.n308 VTAIL.n277 104.615
R226 VTAIL.n301 VTAIL.n277 104.615
R227 VTAIL.n301 VTAIL.n300 104.615
R228 VTAIL.n300 VTAIL.n282 104.615
R229 VTAIL.n293 VTAIL.n282 104.615
R230 VTAIL.n293 VTAIL.n292 104.615
R231 VTAIL.n292 VTAIL.n286 104.615
R232 VTAIL.n264 VTAIL.n263 104.615
R233 VTAIL.n263 VTAIL.n219 104.615
R234 VTAIL.n256 VTAIL.n219 104.615
R235 VTAIL.n256 VTAIL.n255 104.615
R236 VTAIL.n255 VTAIL.n254 104.615
R237 VTAIL.n254 VTAIL.n223 104.615
R238 VTAIL.n247 VTAIL.n223 104.615
R239 VTAIL.n247 VTAIL.n246 104.615
R240 VTAIL.n246 VTAIL.n228 104.615
R241 VTAIL.n239 VTAIL.n228 104.615
R242 VTAIL.n239 VTAIL.n238 104.615
R243 VTAIL.n238 VTAIL.n232 104.615
R244 VTAIL.n210 VTAIL.n209 104.615
R245 VTAIL.n209 VTAIL.n165 104.615
R246 VTAIL.n202 VTAIL.n165 104.615
R247 VTAIL.n202 VTAIL.n201 104.615
R248 VTAIL.n201 VTAIL.n200 104.615
R249 VTAIL.n200 VTAIL.n169 104.615
R250 VTAIL.n193 VTAIL.n169 104.615
R251 VTAIL.n193 VTAIL.n192 104.615
R252 VTAIL.n192 VTAIL.n174 104.615
R253 VTAIL.n185 VTAIL.n174 104.615
R254 VTAIL.n185 VTAIL.n184 104.615
R255 VTAIL.n184 VTAIL.n178 104.615
R256 VTAIL.t7 VTAIL.n393 52.3082
R257 VTAIL.t0 VTAIL.n15 52.3082
R258 VTAIL.t3 VTAIL.n69 52.3082
R259 VTAIL.t1 VTAIL.n123 52.3082
R260 VTAIL.t2 VTAIL.n340 52.3082
R261 VTAIL.t4 VTAIL.n286 52.3082
R262 VTAIL.t5 VTAIL.n232 52.3082
R263 VTAIL.t6 VTAIL.n178 52.3082
R264 VTAIL.n431 VTAIL.n430 31.2157
R265 VTAIL.n53 VTAIL.n52 31.2157
R266 VTAIL.n107 VTAIL.n106 31.2157
R267 VTAIL.n161 VTAIL.n160 31.2157
R268 VTAIL.n377 VTAIL.n376 31.2157
R269 VTAIL.n323 VTAIL.n322 31.2157
R270 VTAIL.n269 VTAIL.n268 31.2157
R271 VTAIL.n215 VTAIL.n214 31.2157
R272 VTAIL.n431 VTAIL.n377 24.1514
R273 VTAIL.n215 VTAIL.n161 24.1514
R274 VTAIL.n419 VTAIL.n384 13.1884
R275 VTAIL.n41 VTAIL.n6 13.1884
R276 VTAIL.n95 VTAIL.n60 13.1884
R277 VTAIL.n149 VTAIL.n114 13.1884
R278 VTAIL.n365 VTAIL.n330 13.1884
R279 VTAIL.n311 VTAIL.n276 13.1884
R280 VTAIL.n257 VTAIL.n222 13.1884
R281 VTAIL.n203 VTAIL.n168 13.1884
R282 VTAIL.n415 VTAIL.n414 12.8005
R283 VTAIL.n420 VTAIL.n382 12.8005
R284 VTAIL.n37 VTAIL.n36 12.8005
R285 VTAIL.n42 VTAIL.n4 12.8005
R286 VTAIL.n91 VTAIL.n90 12.8005
R287 VTAIL.n96 VTAIL.n58 12.8005
R288 VTAIL.n145 VTAIL.n144 12.8005
R289 VTAIL.n150 VTAIL.n112 12.8005
R290 VTAIL.n366 VTAIL.n328 12.8005
R291 VTAIL.n361 VTAIL.n332 12.8005
R292 VTAIL.n312 VTAIL.n274 12.8005
R293 VTAIL.n307 VTAIL.n278 12.8005
R294 VTAIL.n258 VTAIL.n220 12.8005
R295 VTAIL.n253 VTAIL.n224 12.8005
R296 VTAIL.n204 VTAIL.n166 12.8005
R297 VTAIL.n199 VTAIL.n170 12.8005
R298 VTAIL.n413 VTAIL.n386 12.0247
R299 VTAIL.n424 VTAIL.n423 12.0247
R300 VTAIL.n35 VTAIL.n8 12.0247
R301 VTAIL.n46 VTAIL.n45 12.0247
R302 VTAIL.n89 VTAIL.n62 12.0247
R303 VTAIL.n100 VTAIL.n99 12.0247
R304 VTAIL.n143 VTAIL.n116 12.0247
R305 VTAIL.n154 VTAIL.n153 12.0247
R306 VTAIL.n370 VTAIL.n369 12.0247
R307 VTAIL.n360 VTAIL.n333 12.0247
R308 VTAIL.n316 VTAIL.n315 12.0247
R309 VTAIL.n306 VTAIL.n279 12.0247
R310 VTAIL.n262 VTAIL.n261 12.0247
R311 VTAIL.n252 VTAIL.n225 12.0247
R312 VTAIL.n208 VTAIL.n207 12.0247
R313 VTAIL.n198 VTAIL.n171 12.0247
R314 VTAIL.n410 VTAIL.n409 11.249
R315 VTAIL.n427 VTAIL.n380 11.249
R316 VTAIL.n32 VTAIL.n31 11.249
R317 VTAIL.n49 VTAIL.n2 11.249
R318 VTAIL.n86 VTAIL.n85 11.249
R319 VTAIL.n103 VTAIL.n56 11.249
R320 VTAIL.n140 VTAIL.n139 11.249
R321 VTAIL.n157 VTAIL.n110 11.249
R322 VTAIL.n373 VTAIL.n326 11.249
R323 VTAIL.n357 VTAIL.n356 11.249
R324 VTAIL.n319 VTAIL.n272 11.249
R325 VTAIL.n303 VTAIL.n302 11.249
R326 VTAIL.n265 VTAIL.n218 11.249
R327 VTAIL.n249 VTAIL.n248 11.249
R328 VTAIL.n211 VTAIL.n164 11.249
R329 VTAIL.n195 VTAIL.n194 11.249
R330 VTAIL.n406 VTAIL.n388 10.4732
R331 VTAIL.n428 VTAIL.n378 10.4732
R332 VTAIL.n28 VTAIL.n10 10.4732
R333 VTAIL.n50 VTAIL.n0 10.4732
R334 VTAIL.n82 VTAIL.n64 10.4732
R335 VTAIL.n104 VTAIL.n54 10.4732
R336 VTAIL.n136 VTAIL.n118 10.4732
R337 VTAIL.n158 VTAIL.n108 10.4732
R338 VTAIL.n374 VTAIL.n324 10.4732
R339 VTAIL.n353 VTAIL.n335 10.4732
R340 VTAIL.n320 VTAIL.n270 10.4732
R341 VTAIL.n299 VTAIL.n281 10.4732
R342 VTAIL.n266 VTAIL.n216 10.4732
R343 VTAIL.n245 VTAIL.n227 10.4732
R344 VTAIL.n212 VTAIL.n162 10.4732
R345 VTAIL.n191 VTAIL.n173 10.4732
R346 VTAIL.n395 VTAIL.n394 10.2747
R347 VTAIL.n17 VTAIL.n16 10.2747
R348 VTAIL.n71 VTAIL.n70 10.2747
R349 VTAIL.n125 VTAIL.n124 10.2747
R350 VTAIL.n342 VTAIL.n341 10.2747
R351 VTAIL.n288 VTAIL.n287 10.2747
R352 VTAIL.n234 VTAIL.n233 10.2747
R353 VTAIL.n180 VTAIL.n179 10.2747
R354 VTAIL.n405 VTAIL.n390 9.69747
R355 VTAIL.n27 VTAIL.n12 9.69747
R356 VTAIL.n81 VTAIL.n66 9.69747
R357 VTAIL.n135 VTAIL.n120 9.69747
R358 VTAIL.n352 VTAIL.n337 9.69747
R359 VTAIL.n298 VTAIL.n283 9.69747
R360 VTAIL.n244 VTAIL.n229 9.69747
R361 VTAIL.n190 VTAIL.n175 9.69747
R362 VTAIL.n430 VTAIL.n429 9.45567
R363 VTAIL.n52 VTAIL.n51 9.45567
R364 VTAIL.n106 VTAIL.n105 9.45567
R365 VTAIL.n160 VTAIL.n159 9.45567
R366 VTAIL.n376 VTAIL.n375 9.45567
R367 VTAIL.n322 VTAIL.n321 9.45567
R368 VTAIL.n268 VTAIL.n267 9.45567
R369 VTAIL.n214 VTAIL.n213 9.45567
R370 VTAIL.n429 VTAIL.n428 9.3005
R371 VTAIL.n380 VTAIL.n379 9.3005
R372 VTAIL.n423 VTAIL.n422 9.3005
R373 VTAIL.n421 VTAIL.n420 9.3005
R374 VTAIL.n397 VTAIL.n396 9.3005
R375 VTAIL.n392 VTAIL.n391 9.3005
R376 VTAIL.n403 VTAIL.n402 9.3005
R377 VTAIL.n405 VTAIL.n404 9.3005
R378 VTAIL.n388 VTAIL.n387 9.3005
R379 VTAIL.n411 VTAIL.n410 9.3005
R380 VTAIL.n413 VTAIL.n412 9.3005
R381 VTAIL.n414 VTAIL.n383 9.3005
R382 VTAIL.n51 VTAIL.n50 9.3005
R383 VTAIL.n2 VTAIL.n1 9.3005
R384 VTAIL.n45 VTAIL.n44 9.3005
R385 VTAIL.n43 VTAIL.n42 9.3005
R386 VTAIL.n19 VTAIL.n18 9.3005
R387 VTAIL.n14 VTAIL.n13 9.3005
R388 VTAIL.n25 VTAIL.n24 9.3005
R389 VTAIL.n27 VTAIL.n26 9.3005
R390 VTAIL.n10 VTAIL.n9 9.3005
R391 VTAIL.n33 VTAIL.n32 9.3005
R392 VTAIL.n35 VTAIL.n34 9.3005
R393 VTAIL.n36 VTAIL.n5 9.3005
R394 VTAIL.n105 VTAIL.n104 9.3005
R395 VTAIL.n56 VTAIL.n55 9.3005
R396 VTAIL.n99 VTAIL.n98 9.3005
R397 VTAIL.n97 VTAIL.n96 9.3005
R398 VTAIL.n73 VTAIL.n72 9.3005
R399 VTAIL.n68 VTAIL.n67 9.3005
R400 VTAIL.n79 VTAIL.n78 9.3005
R401 VTAIL.n81 VTAIL.n80 9.3005
R402 VTAIL.n64 VTAIL.n63 9.3005
R403 VTAIL.n87 VTAIL.n86 9.3005
R404 VTAIL.n89 VTAIL.n88 9.3005
R405 VTAIL.n90 VTAIL.n59 9.3005
R406 VTAIL.n159 VTAIL.n158 9.3005
R407 VTAIL.n110 VTAIL.n109 9.3005
R408 VTAIL.n153 VTAIL.n152 9.3005
R409 VTAIL.n151 VTAIL.n150 9.3005
R410 VTAIL.n127 VTAIL.n126 9.3005
R411 VTAIL.n122 VTAIL.n121 9.3005
R412 VTAIL.n133 VTAIL.n132 9.3005
R413 VTAIL.n135 VTAIL.n134 9.3005
R414 VTAIL.n118 VTAIL.n117 9.3005
R415 VTAIL.n141 VTAIL.n140 9.3005
R416 VTAIL.n143 VTAIL.n142 9.3005
R417 VTAIL.n144 VTAIL.n113 9.3005
R418 VTAIL.n344 VTAIL.n343 9.3005
R419 VTAIL.n339 VTAIL.n338 9.3005
R420 VTAIL.n350 VTAIL.n349 9.3005
R421 VTAIL.n352 VTAIL.n351 9.3005
R422 VTAIL.n335 VTAIL.n334 9.3005
R423 VTAIL.n358 VTAIL.n357 9.3005
R424 VTAIL.n360 VTAIL.n359 9.3005
R425 VTAIL.n332 VTAIL.n329 9.3005
R426 VTAIL.n375 VTAIL.n374 9.3005
R427 VTAIL.n326 VTAIL.n325 9.3005
R428 VTAIL.n369 VTAIL.n368 9.3005
R429 VTAIL.n367 VTAIL.n366 9.3005
R430 VTAIL.n290 VTAIL.n289 9.3005
R431 VTAIL.n285 VTAIL.n284 9.3005
R432 VTAIL.n296 VTAIL.n295 9.3005
R433 VTAIL.n298 VTAIL.n297 9.3005
R434 VTAIL.n281 VTAIL.n280 9.3005
R435 VTAIL.n304 VTAIL.n303 9.3005
R436 VTAIL.n306 VTAIL.n305 9.3005
R437 VTAIL.n278 VTAIL.n275 9.3005
R438 VTAIL.n321 VTAIL.n320 9.3005
R439 VTAIL.n272 VTAIL.n271 9.3005
R440 VTAIL.n315 VTAIL.n314 9.3005
R441 VTAIL.n313 VTAIL.n312 9.3005
R442 VTAIL.n236 VTAIL.n235 9.3005
R443 VTAIL.n231 VTAIL.n230 9.3005
R444 VTAIL.n242 VTAIL.n241 9.3005
R445 VTAIL.n244 VTAIL.n243 9.3005
R446 VTAIL.n227 VTAIL.n226 9.3005
R447 VTAIL.n250 VTAIL.n249 9.3005
R448 VTAIL.n252 VTAIL.n251 9.3005
R449 VTAIL.n224 VTAIL.n221 9.3005
R450 VTAIL.n267 VTAIL.n266 9.3005
R451 VTAIL.n218 VTAIL.n217 9.3005
R452 VTAIL.n261 VTAIL.n260 9.3005
R453 VTAIL.n259 VTAIL.n258 9.3005
R454 VTAIL.n182 VTAIL.n181 9.3005
R455 VTAIL.n177 VTAIL.n176 9.3005
R456 VTAIL.n188 VTAIL.n187 9.3005
R457 VTAIL.n190 VTAIL.n189 9.3005
R458 VTAIL.n173 VTAIL.n172 9.3005
R459 VTAIL.n196 VTAIL.n195 9.3005
R460 VTAIL.n198 VTAIL.n197 9.3005
R461 VTAIL.n170 VTAIL.n167 9.3005
R462 VTAIL.n213 VTAIL.n212 9.3005
R463 VTAIL.n164 VTAIL.n163 9.3005
R464 VTAIL.n207 VTAIL.n206 9.3005
R465 VTAIL.n205 VTAIL.n204 9.3005
R466 VTAIL.n402 VTAIL.n401 8.92171
R467 VTAIL.n24 VTAIL.n23 8.92171
R468 VTAIL.n78 VTAIL.n77 8.92171
R469 VTAIL.n132 VTAIL.n131 8.92171
R470 VTAIL.n349 VTAIL.n348 8.92171
R471 VTAIL.n295 VTAIL.n294 8.92171
R472 VTAIL.n241 VTAIL.n240 8.92171
R473 VTAIL.n187 VTAIL.n186 8.92171
R474 VTAIL.n398 VTAIL.n392 8.14595
R475 VTAIL.n20 VTAIL.n14 8.14595
R476 VTAIL.n74 VTAIL.n68 8.14595
R477 VTAIL.n128 VTAIL.n122 8.14595
R478 VTAIL.n345 VTAIL.n339 8.14595
R479 VTAIL.n291 VTAIL.n285 8.14595
R480 VTAIL.n237 VTAIL.n231 8.14595
R481 VTAIL.n183 VTAIL.n177 8.14595
R482 VTAIL.n397 VTAIL.n394 7.3702
R483 VTAIL.n19 VTAIL.n16 7.3702
R484 VTAIL.n73 VTAIL.n70 7.3702
R485 VTAIL.n127 VTAIL.n124 7.3702
R486 VTAIL.n344 VTAIL.n341 7.3702
R487 VTAIL.n290 VTAIL.n287 7.3702
R488 VTAIL.n236 VTAIL.n233 7.3702
R489 VTAIL.n182 VTAIL.n179 7.3702
R490 VTAIL.n398 VTAIL.n397 5.81868
R491 VTAIL.n20 VTAIL.n19 5.81868
R492 VTAIL.n74 VTAIL.n73 5.81868
R493 VTAIL.n128 VTAIL.n127 5.81868
R494 VTAIL.n345 VTAIL.n344 5.81868
R495 VTAIL.n291 VTAIL.n290 5.81868
R496 VTAIL.n237 VTAIL.n236 5.81868
R497 VTAIL.n183 VTAIL.n182 5.81868
R498 VTAIL.n401 VTAIL.n392 5.04292
R499 VTAIL.n23 VTAIL.n14 5.04292
R500 VTAIL.n77 VTAIL.n68 5.04292
R501 VTAIL.n131 VTAIL.n122 5.04292
R502 VTAIL.n348 VTAIL.n339 5.04292
R503 VTAIL.n294 VTAIL.n285 5.04292
R504 VTAIL.n240 VTAIL.n231 5.04292
R505 VTAIL.n186 VTAIL.n177 5.04292
R506 VTAIL.n402 VTAIL.n390 4.26717
R507 VTAIL.n24 VTAIL.n12 4.26717
R508 VTAIL.n78 VTAIL.n66 4.26717
R509 VTAIL.n132 VTAIL.n120 4.26717
R510 VTAIL.n349 VTAIL.n337 4.26717
R511 VTAIL.n295 VTAIL.n283 4.26717
R512 VTAIL.n241 VTAIL.n229 4.26717
R513 VTAIL.n187 VTAIL.n175 4.26717
R514 VTAIL.n406 VTAIL.n405 3.49141
R515 VTAIL.n430 VTAIL.n378 3.49141
R516 VTAIL.n28 VTAIL.n27 3.49141
R517 VTAIL.n52 VTAIL.n0 3.49141
R518 VTAIL.n82 VTAIL.n81 3.49141
R519 VTAIL.n106 VTAIL.n54 3.49141
R520 VTAIL.n136 VTAIL.n135 3.49141
R521 VTAIL.n160 VTAIL.n108 3.49141
R522 VTAIL.n376 VTAIL.n324 3.49141
R523 VTAIL.n353 VTAIL.n352 3.49141
R524 VTAIL.n322 VTAIL.n270 3.49141
R525 VTAIL.n299 VTAIL.n298 3.49141
R526 VTAIL.n268 VTAIL.n216 3.49141
R527 VTAIL.n245 VTAIL.n244 3.49141
R528 VTAIL.n214 VTAIL.n162 3.49141
R529 VTAIL.n191 VTAIL.n190 3.49141
R530 VTAIL.n269 VTAIL.n215 3.24188
R531 VTAIL.n377 VTAIL.n323 3.24188
R532 VTAIL.n161 VTAIL.n107 3.24188
R533 VTAIL.n396 VTAIL.n395 2.84303
R534 VTAIL.n18 VTAIL.n17 2.84303
R535 VTAIL.n72 VTAIL.n71 2.84303
R536 VTAIL.n126 VTAIL.n125 2.84303
R537 VTAIL.n343 VTAIL.n342 2.84303
R538 VTAIL.n289 VTAIL.n288 2.84303
R539 VTAIL.n235 VTAIL.n234 2.84303
R540 VTAIL.n181 VTAIL.n180 2.84303
R541 VTAIL.n409 VTAIL.n388 2.71565
R542 VTAIL.n428 VTAIL.n427 2.71565
R543 VTAIL.n31 VTAIL.n10 2.71565
R544 VTAIL.n50 VTAIL.n49 2.71565
R545 VTAIL.n85 VTAIL.n64 2.71565
R546 VTAIL.n104 VTAIL.n103 2.71565
R547 VTAIL.n139 VTAIL.n118 2.71565
R548 VTAIL.n158 VTAIL.n157 2.71565
R549 VTAIL.n374 VTAIL.n373 2.71565
R550 VTAIL.n356 VTAIL.n335 2.71565
R551 VTAIL.n320 VTAIL.n319 2.71565
R552 VTAIL.n302 VTAIL.n281 2.71565
R553 VTAIL.n266 VTAIL.n265 2.71565
R554 VTAIL.n248 VTAIL.n227 2.71565
R555 VTAIL.n212 VTAIL.n211 2.71565
R556 VTAIL.n194 VTAIL.n173 2.71565
R557 VTAIL.n410 VTAIL.n386 1.93989
R558 VTAIL.n424 VTAIL.n380 1.93989
R559 VTAIL.n32 VTAIL.n8 1.93989
R560 VTAIL.n46 VTAIL.n2 1.93989
R561 VTAIL.n86 VTAIL.n62 1.93989
R562 VTAIL.n100 VTAIL.n56 1.93989
R563 VTAIL.n140 VTAIL.n116 1.93989
R564 VTAIL.n154 VTAIL.n110 1.93989
R565 VTAIL.n370 VTAIL.n326 1.93989
R566 VTAIL.n357 VTAIL.n333 1.93989
R567 VTAIL.n316 VTAIL.n272 1.93989
R568 VTAIL.n303 VTAIL.n279 1.93989
R569 VTAIL.n262 VTAIL.n218 1.93989
R570 VTAIL.n249 VTAIL.n225 1.93989
R571 VTAIL.n208 VTAIL.n164 1.93989
R572 VTAIL.n195 VTAIL.n171 1.93989
R573 VTAIL VTAIL.n53 1.67938
R574 VTAIL VTAIL.n431 1.563
R575 VTAIL.n415 VTAIL.n413 1.16414
R576 VTAIL.n423 VTAIL.n382 1.16414
R577 VTAIL.n37 VTAIL.n35 1.16414
R578 VTAIL.n45 VTAIL.n4 1.16414
R579 VTAIL.n91 VTAIL.n89 1.16414
R580 VTAIL.n99 VTAIL.n58 1.16414
R581 VTAIL.n145 VTAIL.n143 1.16414
R582 VTAIL.n153 VTAIL.n112 1.16414
R583 VTAIL.n369 VTAIL.n328 1.16414
R584 VTAIL.n361 VTAIL.n360 1.16414
R585 VTAIL.n315 VTAIL.n274 1.16414
R586 VTAIL.n307 VTAIL.n306 1.16414
R587 VTAIL.n261 VTAIL.n220 1.16414
R588 VTAIL.n253 VTAIL.n252 1.16414
R589 VTAIL.n207 VTAIL.n166 1.16414
R590 VTAIL.n199 VTAIL.n198 1.16414
R591 VTAIL.n323 VTAIL.n269 0.470328
R592 VTAIL.n107 VTAIL.n53 0.470328
R593 VTAIL.n414 VTAIL.n384 0.388379
R594 VTAIL.n420 VTAIL.n419 0.388379
R595 VTAIL.n36 VTAIL.n6 0.388379
R596 VTAIL.n42 VTAIL.n41 0.388379
R597 VTAIL.n90 VTAIL.n60 0.388379
R598 VTAIL.n96 VTAIL.n95 0.388379
R599 VTAIL.n144 VTAIL.n114 0.388379
R600 VTAIL.n150 VTAIL.n149 0.388379
R601 VTAIL.n366 VTAIL.n365 0.388379
R602 VTAIL.n332 VTAIL.n330 0.388379
R603 VTAIL.n312 VTAIL.n311 0.388379
R604 VTAIL.n278 VTAIL.n276 0.388379
R605 VTAIL.n258 VTAIL.n257 0.388379
R606 VTAIL.n224 VTAIL.n222 0.388379
R607 VTAIL.n204 VTAIL.n203 0.388379
R608 VTAIL.n170 VTAIL.n168 0.388379
R609 VTAIL.n396 VTAIL.n391 0.155672
R610 VTAIL.n403 VTAIL.n391 0.155672
R611 VTAIL.n404 VTAIL.n403 0.155672
R612 VTAIL.n404 VTAIL.n387 0.155672
R613 VTAIL.n411 VTAIL.n387 0.155672
R614 VTAIL.n412 VTAIL.n411 0.155672
R615 VTAIL.n412 VTAIL.n383 0.155672
R616 VTAIL.n421 VTAIL.n383 0.155672
R617 VTAIL.n422 VTAIL.n421 0.155672
R618 VTAIL.n422 VTAIL.n379 0.155672
R619 VTAIL.n429 VTAIL.n379 0.155672
R620 VTAIL.n18 VTAIL.n13 0.155672
R621 VTAIL.n25 VTAIL.n13 0.155672
R622 VTAIL.n26 VTAIL.n25 0.155672
R623 VTAIL.n26 VTAIL.n9 0.155672
R624 VTAIL.n33 VTAIL.n9 0.155672
R625 VTAIL.n34 VTAIL.n33 0.155672
R626 VTAIL.n34 VTAIL.n5 0.155672
R627 VTAIL.n43 VTAIL.n5 0.155672
R628 VTAIL.n44 VTAIL.n43 0.155672
R629 VTAIL.n44 VTAIL.n1 0.155672
R630 VTAIL.n51 VTAIL.n1 0.155672
R631 VTAIL.n72 VTAIL.n67 0.155672
R632 VTAIL.n79 VTAIL.n67 0.155672
R633 VTAIL.n80 VTAIL.n79 0.155672
R634 VTAIL.n80 VTAIL.n63 0.155672
R635 VTAIL.n87 VTAIL.n63 0.155672
R636 VTAIL.n88 VTAIL.n87 0.155672
R637 VTAIL.n88 VTAIL.n59 0.155672
R638 VTAIL.n97 VTAIL.n59 0.155672
R639 VTAIL.n98 VTAIL.n97 0.155672
R640 VTAIL.n98 VTAIL.n55 0.155672
R641 VTAIL.n105 VTAIL.n55 0.155672
R642 VTAIL.n126 VTAIL.n121 0.155672
R643 VTAIL.n133 VTAIL.n121 0.155672
R644 VTAIL.n134 VTAIL.n133 0.155672
R645 VTAIL.n134 VTAIL.n117 0.155672
R646 VTAIL.n141 VTAIL.n117 0.155672
R647 VTAIL.n142 VTAIL.n141 0.155672
R648 VTAIL.n142 VTAIL.n113 0.155672
R649 VTAIL.n151 VTAIL.n113 0.155672
R650 VTAIL.n152 VTAIL.n151 0.155672
R651 VTAIL.n152 VTAIL.n109 0.155672
R652 VTAIL.n159 VTAIL.n109 0.155672
R653 VTAIL.n375 VTAIL.n325 0.155672
R654 VTAIL.n368 VTAIL.n325 0.155672
R655 VTAIL.n368 VTAIL.n367 0.155672
R656 VTAIL.n367 VTAIL.n329 0.155672
R657 VTAIL.n359 VTAIL.n329 0.155672
R658 VTAIL.n359 VTAIL.n358 0.155672
R659 VTAIL.n358 VTAIL.n334 0.155672
R660 VTAIL.n351 VTAIL.n334 0.155672
R661 VTAIL.n351 VTAIL.n350 0.155672
R662 VTAIL.n350 VTAIL.n338 0.155672
R663 VTAIL.n343 VTAIL.n338 0.155672
R664 VTAIL.n321 VTAIL.n271 0.155672
R665 VTAIL.n314 VTAIL.n271 0.155672
R666 VTAIL.n314 VTAIL.n313 0.155672
R667 VTAIL.n313 VTAIL.n275 0.155672
R668 VTAIL.n305 VTAIL.n275 0.155672
R669 VTAIL.n305 VTAIL.n304 0.155672
R670 VTAIL.n304 VTAIL.n280 0.155672
R671 VTAIL.n297 VTAIL.n280 0.155672
R672 VTAIL.n297 VTAIL.n296 0.155672
R673 VTAIL.n296 VTAIL.n284 0.155672
R674 VTAIL.n289 VTAIL.n284 0.155672
R675 VTAIL.n267 VTAIL.n217 0.155672
R676 VTAIL.n260 VTAIL.n217 0.155672
R677 VTAIL.n260 VTAIL.n259 0.155672
R678 VTAIL.n259 VTAIL.n221 0.155672
R679 VTAIL.n251 VTAIL.n221 0.155672
R680 VTAIL.n251 VTAIL.n250 0.155672
R681 VTAIL.n250 VTAIL.n226 0.155672
R682 VTAIL.n243 VTAIL.n226 0.155672
R683 VTAIL.n243 VTAIL.n242 0.155672
R684 VTAIL.n242 VTAIL.n230 0.155672
R685 VTAIL.n235 VTAIL.n230 0.155672
R686 VTAIL.n213 VTAIL.n163 0.155672
R687 VTAIL.n206 VTAIL.n163 0.155672
R688 VTAIL.n206 VTAIL.n205 0.155672
R689 VTAIL.n205 VTAIL.n167 0.155672
R690 VTAIL.n197 VTAIL.n167 0.155672
R691 VTAIL.n197 VTAIL.n196 0.155672
R692 VTAIL.n196 VTAIL.n172 0.155672
R693 VTAIL.n189 VTAIL.n172 0.155672
R694 VTAIL.n189 VTAIL.n188 0.155672
R695 VTAIL.n188 VTAIL.n176 0.155672
R696 VTAIL.n181 VTAIL.n176 0.155672
R697 B.n560 B.n356 588.598
R698 B.n121 B.n74 588.598
R699 B.n563 B.n358 588.598
R700 B.n741 B.n76 588.598
R701 B.n741 B.n740 585
R702 B.n279 B.n116 585
R703 B.n278 B.n277 585
R704 B.n276 B.n275 585
R705 B.n274 B.n273 585
R706 B.n272 B.n271 585
R707 B.n270 B.n269 585
R708 B.n268 B.n267 585
R709 B.n266 B.n265 585
R710 B.n264 B.n263 585
R711 B.n262 B.n261 585
R712 B.n260 B.n259 585
R713 B.n258 B.n257 585
R714 B.n256 B.n255 585
R715 B.n254 B.n253 585
R716 B.n252 B.n251 585
R717 B.n250 B.n249 585
R718 B.n248 B.n247 585
R719 B.n246 B.n245 585
R720 B.n244 B.n243 585
R721 B.n242 B.n241 585
R722 B.n240 B.n239 585
R723 B.n238 B.n237 585
R724 B.n236 B.n235 585
R725 B.n234 B.n233 585
R726 B.n232 B.n231 585
R727 B.n230 B.n229 585
R728 B.n228 B.n227 585
R729 B.n226 B.n225 585
R730 B.n224 B.n223 585
R731 B.n222 B.n221 585
R732 B.n220 B.n219 585
R733 B.n218 B.n217 585
R734 B.n216 B.n215 585
R735 B.n214 B.n213 585
R736 B.n211 B.n210 585
R737 B.n209 B.n208 585
R738 B.n207 B.n206 585
R739 B.n205 B.n204 585
R740 B.n203 B.n202 585
R741 B.n201 B.n200 585
R742 B.n199 B.n198 585
R743 B.n197 B.n196 585
R744 B.n195 B.n194 585
R745 B.n193 B.n192 585
R746 B.n190 B.n189 585
R747 B.n188 B.n187 585
R748 B.n186 B.n185 585
R749 B.n184 B.n183 585
R750 B.n182 B.n181 585
R751 B.n180 B.n179 585
R752 B.n178 B.n177 585
R753 B.n176 B.n175 585
R754 B.n174 B.n173 585
R755 B.n172 B.n171 585
R756 B.n170 B.n169 585
R757 B.n168 B.n167 585
R758 B.n166 B.n165 585
R759 B.n164 B.n163 585
R760 B.n162 B.n161 585
R761 B.n160 B.n159 585
R762 B.n158 B.n157 585
R763 B.n156 B.n155 585
R764 B.n154 B.n153 585
R765 B.n152 B.n151 585
R766 B.n150 B.n149 585
R767 B.n148 B.n147 585
R768 B.n146 B.n145 585
R769 B.n144 B.n143 585
R770 B.n142 B.n141 585
R771 B.n140 B.n139 585
R772 B.n138 B.n137 585
R773 B.n136 B.n135 585
R774 B.n134 B.n133 585
R775 B.n132 B.n131 585
R776 B.n130 B.n129 585
R777 B.n128 B.n127 585
R778 B.n126 B.n125 585
R779 B.n124 B.n123 585
R780 B.n122 B.n121 585
R781 B.n739 B.n76 585
R782 B.n744 B.n76 585
R783 B.n738 B.n75 585
R784 B.n745 B.n75 585
R785 B.n737 B.n736 585
R786 B.n736 B.n71 585
R787 B.n735 B.n70 585
R788 B.n751 B.n70 585
R789 B.n734 B.n69 585
R790 B.n752 B.n69 585
R791 B.n733 B.n68 585
R792 B.n753 B.n68 585
R793 B.n732 B.n731 585
R794 B.n731 B.n64 585
R795 B.n730 B.n63 585
R796 B.n759 B.n63 585
R797 B.n729 B.n62 585
R798 B.n760 B.n62 585
R799 B.n728 B.n61 585
R800 B.n761 B.n61 585
R801 B.n727 B.n726 585
R802 B.n726 B.n57 585
R803 B.n725 B.n56 585
R804 B.n767 B.n56 585
R805 B.n724 B.n55 585
R806 B.n768 B.n55 585
R807 B.n723 B.n54 585
R808 B.n769 B.n54 585
R809 B.n722 B.n721 585
R810 B.n721 B.n50 585
R811 B.n720 B.n49 585
R812 B.n775 B.n49 585
R813 B.n719 B.n48 585
R814 B.n776 B.n48 585
R815 B.n718 B.n47 585
R816 B.n777 B.n47 585
R817 B.n717 B.n716 585
R818 B.n716 B.n43 585
R819 B.n715 B.n42 585
R820 B.n783 B.n42 585
R821 B.n714 B.n41 585
R822 B.n784 B.n41 585
R823 B.n713 B.n40 585
R824 B.n785 B.n40 585
R825 B.n712 B.n711 585
R826 B.n711 B.n39 585
R827 B.n710 B.n35 585
R828 B.n791 B.n35 585
R829 B.n709 B.n34 585
R830 B.n792 B.n34 585
R831 B.n708 B.n33 585
R832 B.n793 B.n33 585
R833 B.n707 B.n706 585
R834 B.n706 B.n29 585
R835 B.n705 B.n28 585
R836 B.n799 B.n28 585
R837 B.n704 B.n27 585
R838 B.n800 B.n27 585
R839 B.n703 B.n26 585
R840 B.n801 B.n26 585
R841 B.n702 B.n701 585
R842 B.n701 B.n22 585
R843 B.n700 B.n21 585
R844 B.n807 B.n21 585
R845 B.n699 B.n20 585
R846 B.n808 B.n20 585
R847 B.n698 B.n19 585
R848 B.n809 B.n19 585
R849 B.n697 B.n696 585
R850 B.n696 B.n15 585
R851 B.n695 B.n14 585
R852 B.n815 B.n14 585
R853 B.n694 B.n13 585
R854 B.n816 B.n13 585
R855 B.n693 B.n12 585
R856 B.n817 B.n12 585
R857 B.n692 B.n691 585
R858 B.n691 B.n8 585
R859 B.n690 B.n7 585
R860 B.n823 B.n7 585
R861 B.n689 B.n6 585
R862 B.n824 B.n6 585
R863 B.n688 B.n5 585
R864 B.n825 B.n5 585
R865 B.n687 B.n686 585
R866 B.n686 B.n4 585
R867 B.n685 B.n280 585
R868 B.n685 B.n684 585
R869 B.n675 B.n281 585
R870 B.n282 B.n281 585
R871 B.n677 B.n676 585
R872 B.n678 B.n677 585
R873 B.n674 B.n287 585
R874 B.n287 B.n286 585
R875 B.n673 B.n672 585
R876 B.n672 B.n671 585
R877 B.n289 B.n288 585
R878 B.n290 B.n289 585
R879 B.n664 B.n663 585
R880 B.n665 B.n664 585
R881 B.n662 B.n295 585
R882 B.n295 B.n294 585
R883 B.n661 B.n660 585
R884 B.n660 B.n659 585
R885 B.n297 B.n296 585
R886 B.n298 B.n297 585
R887 B.n652 B.n651 585
R888 B.n653 B.n652 585
R889 B.n650 B.n303 585
R890 B.n303 B.n302 585
R891 B.n649 B.n648 585
R892 B.n648 B.n647 585
R893 B.n305 B.n304 585
R894 B.n306 B.n305 585
R895 B.n640 B.n639 585
R896 B.n641 B.n640 585
R897 B.n638 B.n311 585
R898 B.n311 B.n310 585
R899 B.n637 B.n636 585
R900 B.n636 B.n635 585
R901 B.n313 B.n312 585
R902 B.n628 B.n313 585
R903 B.n627 B.n626 585
R904 B.n629 B.n627 585
R905 B.n625 B.n318 585
R906 B.n318 B.n317 585
R907 B.n624 B.n623 585
R908 B.n623 B.n622 585
R909 B.n320 B.n319 585
R910 B.n321 B.n320 585
R911 B.n615 B.n614 585
R912 B.n616 B.n615 585
R913 B.n613 B.n326 585
R914 B.n326 B.n325 585
R915 B.n612 B.n611 585
R916 B.n611 B.n610 585
R917 B.n328 B.n327 585
R918 B.n329 B.n328 585
R919 B.n603 B.n602 585
R920 B.n604 B.n603 585
R921 B.n601 B.n334 585
R922 B.n334 B.n333 585
R923 B.n600 B.n599 585
R924 B.n599 B.n598 585
R925 B.n336 B.n335 585
R926 B.n337 B.n336 585
R927 B.n591 B.n590 585
R928 B.n592 B.n591 585
R929 B.n589 B.n341 585
R930 B.n345 B.n341 585
R931 B.n588 B.n587 585
R932 B.n587 B.n586 585
R933 B.n343 B.n342 585
R934 B.n344 B.n343 585
R935 B.n579 B.n578 585
R936 B.n580 B.n579 585
R937 B.n577 B.n350 585
R938 B.n350 B.n349 585
R939 B.n576 B.n575 585
R940 B.n575 B.n574 585
R941 B.n352 B.n351 585
R942 B.n353 B.n352 585
R943 B.n567 B.n566 585
R944 B.n568 B.n567 585
R945 B.n565 B.n358 585
R946 B.n358 B.n357 585
R947 B.n560 B.n559 585
R948 B.n558 B.n400 585
R949 B.n557 B.n399 585
R950 B.n562 B.n399 585
R951 B.n556 B.n555 585
R952 B.n554 B.n553 585
R953 B.n552 B.n551 585
R954 B.n550 B.n549 585
R955 B.n548 B.n547 585
R956 B.n546 B.n545 585
R957 B.n544 B.n543 585
R958 B.n542 B.n541 585
R959 B.n540 B.n539 585
R960 B.n538 B.n537 585
R961 B.n536 B.n535 585
R962 B.n534 B.n533 585
R963 B.n532 B.n531 585
R964 B.n530 B.n529 585
R965 B.n528 B.n527 585
R966 B.n526 B.n525 585
R967 B.n524 B.n523 585
R968 B.n522 B.n521 585
R969 B.n520 B.n519 585
R970 B.n518 B.n517 585
R971 B.n516 B.n515 585
R972 B.n514 B.n513 585
R973 B.n512 B.n511 585
R974 B.n510 B.n509 585
R975 B.n508 B.n507 585
R976 B.n506 B.n505 585
R977 B.n504 B.n503 585
R978 B.n502 B.n501 585
R979 B.n500 B.n499 585
R980 B.n498 B.n497 585
R981 B.n496 B.n495 585
R982 B.n494 B.n493 585
R983 B.n492 B.n491 585
R984 B.n490 B.n489 585
R985 B.n488 B.n487 585
R986 B.n486 B.n485 585
R987 B.n484 B.n483 585
R988 B.n482 B.n481 585
R989 B.n480 B.n479 585
R990 B.n478 B.n477 585
R991 B.n476 B.n475 585
R992 B.n474 B.n473 585
R993 B.n472 B.n471 585
R994 B.n470 B.n469 585
R995 B.n468 B.n467 585
R996 B.n466 B.n465 585
R997 B.n464 B.n463 585
R998 B.n462 B.n461 585
R999 B.n460 B.n459 585
R1000 B.n458 B.n457 585
R1001 B.n456 B.n455 585
R1002 B.n454 B.n453 585
R1003 B.n452 B.n451 585
R1004 B.n450 B.n449 585
R1005 B.n448 B.n447 585
R1006 B.n446 B.n445 585
R1007 B.n444 B.n443 585
R1008 B.n442 B.n441 585
R1009 B.n440 B.n439 585
R1010 B.n438 B.n437 585
R1011 B.n436 B.n435 585
R1012 B.n434 B.n433 585
R1013 B.n432 B.n431 585
R1014 B.n430 B.n429 585
R1015 B.n428 B.n427 585
R1016 B.n426 B.n425 585
R1017 B.n424 B.n423 585
R1018 B.n422 B.n421 585
R1019 B.n420 B.n419 585
R1020 B.n418 B.n417 585
R1021 B.n416 B.n415 585
R1022 B.n414 B.n413 585
R1023 B.n412 B.n411 585
R1024 B.n410 B.n409 585
R1025 B.n408 B.n407 585
R1026 B.n360 B.n359 585
R1027 B.n564 B.n563 585
R1028 B.n563 B.n562 585
R1029 B.n356 B.n355 585
R1030 B.n357 B.n356 585
R1031 B.n570 B.n569 585
R1032 B.n569 B.n568 585
R1033 B.n571 B.n354 585
R1034 B.n354 B.n353 585
R1035 B.n573 B.n572 585
R1036 B.n574 B.n573 585
R1037 B.n348 B.n347 585
R1038 B.n349 B.n348 585
R1039 B.n582 B.n581 585
R1040 B.n581 B.n580 585
R1041 B.n583 B.n346 585
R1042 B.n346 B.n344 585
R1043 B.n585 B.n584 585
R1044 B.n586 B.n585 585
R1045 B.n340 B.n339 585
R1046 B.n345 B.n340 585
R1047 B.n594 B.n593 585
R1048 B.n593 B.n592 585
R1049 B.n595 B.n338 585
R1050 B.n338 B.n337 585
R1051 B.n597 B.n596 585
R1052 B.n598 B.n597 585
R1053 B.n332 B.n331 585
R1054 B.n333 B.n332 585
R1055 B.n606 B.n605 585
R1056 B.n605 B.n604 585
R1057 B.n607 B.n330 585
R1058 B.n330 B.n329 585
R1059 B.n609 B.n608 585
R1060 B.n610 B.n609 585
R1061 B.n324 B.n323 585
R1062 B.n325 B.n324 585
R1063 B.n618 B.n617 585
R1064 B.n617 B.n616 585
R1065 B.n619 B.n322 585
R1066 B.n322 B.n321 585
R1067 B.n621 B.n620 585
R1068 B.n622 B.n621 585
R1069 B.n316 B.n315 585
R1070 B.n317 B.n316 585
R1071 B.n631 B.n630 585
R1072 B.n630 B.n629 585
R1073 B.n632 B.n314 585
R1074 B.n628 B.n314 585
R1075 B.n634 B.n633 585
R1076 B.n635 B.n634 585
R1077 B.n309 B.n308 585
R1078 B.n310 B.n309 585
R1079 B.n643 B.n642 585
R1080 B.n642 B.n641 585
R1081 B.n644 B.n307 585
R1082 B.n307 B.n306 585
R1083 B.n646 B.n645 585
R1084 B.n647 B.n646 585
R1085 B.n301 B.n300 585
R1086 B.n302 B.n301 585
R1087 B.n655 B.n654 585
R1088 B.n654 B.n653 585
R1089 B.n656 B.n299 585
R1090 B.n299 B.n298 585
R1091 B.n658 B.n657 585
R1092 B.n659 B.n658 585
R1093 B.n293 B.n292 585
R1094 B.n294 B.n293 585
R1095 B.n667 B.n666 585
R1096 B.n666 B.n665 585
R1097 B.n668 B.n291 585
R1098 B.n291 B.n290 585
R1099 B.n670 B.n669 585
R1100 B.n671 B.n670 585
R1101 B.n285 B.n284 585
R1102 B.n286 B.n285 585
R1103 B.n680 B.n679 585
R1104 B.n679 B.n678 585
R1105 B.n681 B.n283 585
R1106 B.n283 B.n282 585
R1107 B.n683 B.n682 585
R1108 B.n684 B.n683 585
R1109 B.n2 B.n0 585
R1110 B.n4 B.n2 585
R1111 B.n3 B.n1 585
R1112 B.n824 B.n3 585
R1113 B.n822 B.n821 585
R1114 B.n823 B.n822 585
R1115 B.n820 B.n9 585
R1116 B.n9 B.n8 585
R1117 B.n819 B.n818 585
R1118 B.n818 B.n817 585
R1119 B.n11 B.n10 585
R1120 B.n816 B.n11 585
R1121 B.n814 B.n813 585
R1122 B.n815 B.n814 585
R1123 B.n812 B.n16 585
R1124 B.n16 B.n15 585
R1125 B.n811 B.n810 585
R1126 B.n810 B.n809 585
R1127 B.n18 B.n17 585
R1128 B.n808 B.n18 585
R1129 B.n806 B.n805 585
R1130 B.n807 B.n806 585
R1131 B.n804 B.n23 585
R1132 B.n23 B.n22 585
R1133 B.n803 B.n802 585
R1134 B.n802 B.n801 585
R1135 B.n25 B.n24 585
R1136 B.n800 B.n25 585
R1137 B.n798 B.n797 585
R1138 B.n799 B.n798 585
R1139 B.n796 B.n30 585
R1140 B.n30 B.n29 585
R1141 B.n795 B.n794 585
R1142 B.n794 B.n793 585
R1143 B.n32 B.n31 585
R1144 B.n792 B.n32 585
R1145 B.n790 B.n789 585
R1146 B.n791 B.n790 585
R1147 B.n788 B.n36 585
R1148 B.n39 B.n36 585
R1149 B.n787 B.n786 585
R1150 B.n786 B.n785 585
R1151 B.n38 B.n37 585
R1152 B.n784 B.n38 585
R1153 B.n782 B.n781 585
R1154 B.n783 B.n782 585
R1155 B.n780 B.n44 585
R1156 B.n44 B.n43 585
R1157 B.n779 B.n778 585
R1158 B.n778 B.n777 585
R1159 B.n46 B.n45 585
R1160 B.n776 B.n46 585
R1161 B.n774 B.n773 585
R1162 B.n775 B.n774 585
R1163 B.n772 B.n51 585
R1164 B.n51 B.n50 585
R1165 B.n771 B.n770 585
R1166 B.n770 B.n769 585
R1167 B.n53 B.n52 585
R1168 B.n768 B.n53 585
R1169 B.n766 B.n765 585
R1170 B.n767 B.n766 585
R1171 B.n764 B.n58 585
R1172 B.n58 B.n57 585
R1173 B.n763 B.n762 585
R1174 B.n762 B.n761 585
R1175 B.n60 B.n59 585
R1176 B.n760 B.n60 585
R1177 B.n758 B.n757 585
R1178 B.n759 B.n758 585
R1179 B.n756 B.n65 585
R1180 B.n65 B.n64 585
R1181 B.n755 B.n754 585
R1182 B.n754 B.n753 585
R1183 B.n67 B.n66 585
R1184 B.n752 B.n67 585
R1185 B.n750 B.n749 585
R1186 B.n751 B.n750 585
R1187 B.n748 B.n72 585
R1188 B.n72 B.n71 585
R1189 B.n747 B.n746 585
R1190 B.n746 B.n745 585
R1191 B.n74 B.n73 585
R1192 B.n744 B.n74 585
R1193 B.n827 B.n826 585
R1194 B.n826 B.n825 585
R1195 B.n404 B.t11 318.822
R1196 B.n117 B.t6 318.822
R1197 B.n401 B.t14 318.822
R1198 B.n119 B.t16 318.822
R1199 B.n404 B.t8 278.661
R1200 B.n401 B.t12 278.661
R1201 B.n119 B.t15 278.661
R1202 B.n117 B.t4 278.661
R1203 B.n743 B.n742 256.663
R1204 B.n743 B.n115 256.663
R1205 B.n743 B.n114 256.663
R1206 B.n743 B.n113 256.663
R1207 B.n743 B.n112 256.663
R1208 B.n743 B.n111 256.663
R1209 B.n743 B.n110 256.663
R1210 B.n743 B.n109 256.663
R1211 B.n743 B.n108 256.663
R1212 B.n743 B.n107 256.663
R1213 B.n743 B.n106 256.663
R1214 B.n743 B.n105 256.663
R1215 B.n743 B.n104 256.663
R1216 B.n743 B.n103 256.663
R1217 B.n743 B.n102 256.663
R1218 B.n743 B.n101 256.663
R1219 B.n743 B.n100 256.663
R1220 B.n743 B.n99 256.663
R1221 B.n743 B.n98 256.663
R1222 B.n743 B.n97 256.663
R1223 B.n743 B.n96 256.663
R1224 B.n743 B.n95 256.663
R1225 B.n743 B.n94 256.663
R1226 B.n743 B.n93 256.663
R1227 B.n743 B.n92 256.663
R1228 B.n743 B.n91 256.663
R1229 B.n743 B.n90 256.663
R1230 B.n743 B.n89 256.663
R1231 B.n743 B.n88 256.663
R1232 B.n743 B.n87 256.663
R1233 B.n743 B.n86 256.663
R1234 B.n743 B.n85 256.663
R1235 B.n743 B.n84 256.663
R1236 B.n743 B.n83 256.663
R1237 B.n743 B.n82 256.663
R1238 B.n743 B.n81 256.663
R1239 B.n743 B.n80 256.663
R1240 B.n743 B.n79 256.663
R1241 B.n743 B.n78 256.663
R1242 B.n743 B.n77 256.663
R1243 B.n562 B.n561 256.663
R1244 B.n562 B.n361 256.663
R1245 B.n562 B.n362 256.663
R1246 B.n562 B.n363 256.663
R1247 B.n562 B.n364 256.663
R1248 B.n562 B.n365 256.663
R1249 B.n562 B.n366 256.663
R1250 B.n562 B.n367 256.663
R1251 B.n562 B.n368 256.663
R1252 B.n562 B.n369 256.663
R1253 B.n562 B.n370 256.663
R1254 B.n562 B.n371 256.663
R1255 B.n562 B.n372 256.663
R1256 B.n562 B.n373 256.663
R1257 B.n562 B.n374 256.663
R1258 B.n562 B.n375 256.663
R1259 B.n562 B.n376 256.663
R1260 B.n562 B.n377 256.663
R1261 B.n562 B.n378 256.663
R1262 B.n562 B.n379 256.663
R1263 B.n562 B.n380 256.663
R1264 B.n562 B.n381 256.663
R1265 B.n562 B.n382 256.663
R1266 B.n562 B.n383 256.663
R1267 B.n562 B.n384 256.663
R1268 B.n562 B.n385 256.663
R1269 B.n562 B.n386 256.663
R1270 B.n562 B.n387 256.663
R1271 B.n562 B.n388 256.663
R1272 B.n562 B.n389 256.663
R1273 B.n562 B.n390 256.663
R1274 B.n562 B.n391 256.663
R1275 B.n562 B.n392 256.663
R1276 B.n562 B.n393 256.663
R1277 B.n562 B.n394 256.663
R1278 B.n562 B.n395 256.663
R1279 B.n562 B.n396 256.663
R1280 B.n562 B.n397 256.663
R1281 B.n562 B.n398 256.663
R1282 B.n405 B.t10 245.901
R1283 B.n118 B.t7 245.901
R1284 B.n402 B.t13 245.901
R1285 B.n120 B.t17 245.901
R1286 B.n569 B.n356 163.367
R1287 B.n569 B.n354 163.367
R1288 B.n573 B.n354 163.367
R1289 B.n573 B.n348 163.367
R1290 B.n581 B.n348 163.367
R1291 B.n581 B.n346 163.367
R1292 B.n585 B.n346 163.367
R1293 B.n585 B.n340 163.367
R1294 B.n593 B.n340 163.367
R1295 B.n593 B.n338 163.367
R1296 B.n597 B.n338 163.367
R1297 B.n597 B.n332 163.367
R1298 B.n605 B.n332 163.367
R1299 B.n605 B.n330 163.367
R1300 B.n609 B.n330 163.367
R1301 B.n609 B.n324 163.367
R1302 B.n617 B.n324 163.367
R1303 B.n617 B.n322 163.367
R1304 B.n621 B.n322 163.367
R1305 B.n621 B.n316 163.367
R1306 B.n630 B.n316 163.367
R1307 B.n630 B.n314 163.367
R1308 B.n634 B.n314 163.367
R1309 B.n634 B.n309 163.367
R1310 B.n642 B.n309 163.367
R1311 B.n642 B.n307 163.367
R1312 B.n646 B.n307 163.367
R1313 B.n646 B.n301 163.367
R1314 B.n654 B.n301 163.367
R1315 B.n654 B.n299 163.367
R1316 B.n658 B.n299 163.367
R1317 B.n658 B.n293 163.367
R1318 B.n666 B.n293 163.367
R1319 B.n666 B.n291 163.367
R1320 B.n670 B.n291 163.367
R1321 B.n670 B.n285 163.367
R1322 B.n679 B.n285 163.367
R1323 B.n679 B.n283 163.367
R1324 B.n683 B.n283 163.367
R1325 B.n683 B.n2 163.367
R1326 B.n826 B.n2 163.367
R1327 B.n826 B.n3 163.367
R1328 B.n822 B.n3 163.367
R1329 B.n822 B.n9 163.367
R1330 B.n818 B.n9 163.367
R1331 B.n818 B.n11 163.367
R1332 B.n814 B.n11 163.367
R1333 B.n814 B.n16 163.367
R1334 B.n810 B.n16 163.367
R1335 B.n810 B.n18 163.367
R1336 B.n806 B.n18 163.367
R1337 B.n806 B.n23 163.367
R1338 B.n802 B.n23 163.367
R1339 B.n802 B.n25 163.367
R1340 B.n798 B.n25 163.367
R1341 B.n798 B.n30 163.367
R1342 B.n794 B.n30 163.367
R1343 B.n794 B.n32 163.367
R1344 B.n790 B.n32 163.367
R1345 B.n790 B.n36 163.367
R1346 B.n786 B.n36 163.367
R1347 B.n786 B.n38 163.367
R1348 B.n782 B.n38 163.367
R1349 B.n782 B.n44 163.367
R1350 B.n778 B.n44 163.367
R1351 B.n778 B.n46 163.367
R1352 B.n774 B.n46 163.367
R1353 B.n774 B.n51 163.367
R1354 B.n770 B.n51 163.367
R1355 B.n770 B.n53 163.367
R1356 B.n766 B.n53 163.367
R1357 B.n766 B.n58 163.367
R1358 B.n762 B.n58 163.367
R1359 B.n762 B.n60 163.367
R1360 B.n758 B.n60 163.367
R1361 B.n758 B.n65 163.367
R1362 B.n754 B.n65 163.367
R1363 B.n754 B.n67 163.367
R1364 B.n750 B.n67 163.367
R1365 B.n750 B.n72 163.367
R1366 B.n746 B.n72 163.367
R1367 B.n746 B.n74 163.367
R1368 B.n400 B.n399 163.367
R1369 B.n555 B.n399 163.367
R1370 B.n553 B.n552 163.367
R1371 B.n549 B.n548 163.367
R1372 B.n545 B.n544 163.367
R1373 B.n541 B.n540 163.367
R1374 B.n537 B.n536 163.367
R1375 B.n533 B.n532 163.367
R1376 B.n529 B.n528 163.367
R1377 B.n525 B.n524 163.367
R1378 B.n521 B.n520 163.367
R1379 B.n517 B.n516 163.367
R1380 B.n513 B.n512 163.367
R1381 B.n509 B.n508 163.367
R1382 B.n505 B.n504 163.367
R1383 B.n501 B.n500 163.367
R1384 B.n497 B.n496 163.367
R1385 B.n493 B.n492 163.367
R1386 B.n489 B.n488 163.367
R1387 B.n485 B.n484 163.367
R1388 B.n481 B.n480 163.367
R1389 B.n477 B.n476 163.367
R1390 B.n473 B.n472 163.367
R1391 B.n469 B.n468 163.367
R1392 B.n465 B.n464 163.367
R1393 B.n461 B.n460 163.367
R1394 B.n457 B.n456 163.367
R1395 B.n453 B.n452 163.367
R1396 B.n449 B.n448 163.367
R1397 B.n445 B.n444 163.367
R1398 B.n441 B.n440 163.367
R1399 B.n437 B.n436 163.367
R1400 B.n433 B.n432 163.367
R1401 B.n429 B.n428 163.367
R1402 B.n425 B.n424 163.367
R1403 B.n421 B.n420 163.367
R1404 B.n417 B.n416 163.367
R1405 B.n413 B.n412 163.367
R1406 B.n409 B.n408 163.367
R1407 B.n563 B.n360 163.367
R1408 B.n567 B.n358 163.367
R1409 B.n567 B.n352 163.367
R1410 B.n575 B.n352 163.367
R1411 B.n575 B.n350 163.367
R1412 B.n579 B.n350 163.367
R1413 B.n579 B.n343 163.367
R1414 B.n587 B.n343 163.367
R1415 B.n587 B.n341 163.367
R1416 B.n591 B.n341 163.367
R1417 B.n591 B.n336 163.367
R1418 B.n599 B.n336 163.367
R1419 B.n599 B.n334 163.367
R1420 B.n603 B.n334 163.367
R1421 B.n603 B.n328 163.367
R1422 B.n611 B.n328 163.367
R1423 B.n611 B.n326 163.367
R1424 B.n615 B.n326 163.367
R1425 B.n615 B.n320 163.367
R1426 B.n623 B.n320 163.367
R1427 B.n623 B.n318 163.367
R1428 B.n627 B.n318 163.367
R1429 B.n627 B.n313 163.367
R1430 B.n636 B.n313 163.367
R1431 B.n636 B.n311 163.367
R1432 B.n640 B.n311 163.367
R1433 B.n640 B.n305 163.367
R1434 B.n648 B.n305 163.367
R1435 B.n648 B.n303 163.367
R1436 B.n652 B.n303 163.367
R1437 B.n652 B.n297 163.367
R1438 B.n660 B.n297 163.367
R1439 B.n660 B.n295 163.367
R1440 B.n664 B.n295 163.367
R1441 B.n664 B.n289 163.367
R1442 B.n672 B.n289 163.367
R1443 B.n672 B.n287 163.367
R1444 B.n677 B.n287 163.367
R1445 B.n677 B.n281 163.367
R1446 B.n685 B.n281 163.367
R1447 B.n686 B.n685 163.367
R1448 B.n686 B.n5 163.367
R1449 B.n6 B.n5 163.367
R1450 B.n7 B.n6 163.367
R1451 B.n691 B.n7 163.367
R1452 B.n691 B.n12 163.367
R1453 B.n13 B.n12 163.367
R1454 B.n14 B.n13 163.367
R1455 B.n696 B.n14 163.367
R1456 B.n696 B.n19 163.367
R1457 B.n20 B.n19 163.367
R1458 B.n21 B.n20 163.367
R1459 B.n701 B.n21 163.367
R1460 B.n701 B.n26 163.367
R1461 B.n27 B.n26 163.367
R1462 B.n28 B.n27 163.367
R1463 B.n706 B.n28 163.367
R1464 B.n706 B.n33 163.367
R1465 B.n34 B.n33 163.367
R1466 B.n35 B.n34 163.367
R1467 B.n711 B.n35 163.367
R1468 B.n711 B.n40 163.367
R1469 B.n41 B.n40 163.367
R1470 B.n42 B.n41 163.367
R1471 B.n716 B.n42 163.367
R1472 B.n716 B.n47 163.367
R1473 B.n48 B.n47 163.367
R1474 B.n49 B.n48 163.367
R1475 B.n721 B.n49 163.367
R1476 B.n721 B.n54 163.367
R1477 B.n55 B.n54 163.367
R1478 B.n56 B.n55 163.367
R1479 B.n726 B.n56 163.367
R1480 B.n726 B.n61 163.367
R1481 B.n62 B.n61 163.367
R1482 B.n63 B.n62 163.367
R1483 B.n731 B.n63 163.367
R1484 B.n731 B.n68 163.367
R1485 B.n69 B.n68 163.367
R1486 B.n70 B.n69 163.367
R1487 B.n736 B.n70 163.367
R1488 B.n736 B.n75 163.367
R1489 B.n76 B.n75 163.367
R1490 B.n125 B.n124 163.367
R1491 B.n129 B.n128 163.367
R1492 B.n133 B.n132 163.367
R1493 B.n137 B.n136 163.367
R1494 B.n141 B.n140 163.367
R1495 B.n145 B.n144 163.367
R1496 B.n149 B.n148 163.367
R1497 B.n153 B.n152 163.367
R1498 B.n157 B.n156 163.367
R1499 B.n161 B.n160 163.367
R1500 B.n165 B.n164 163.367
R1501 B.n169 B.n168 163.367
R1502 B.n173 B.n172 163.367
R1503 B.n177 B.n176 163.367
R1504 B.n181 B.n180 163.367
R1505 B.n185 B.n184 163.367
R1506 B.n189 B.n188 163.367
R1507 B.n194 B.n193 163.367
R1508 B.n198 B.n197 163.367
R1509 B.n202 B.n201 163.367
R1510 B.n206 B.n205 163.367
R1511 B.n210 B.n209 163.367
R1512 B.n215 B.n214 163.367
R1513 B.n219 B.n218 163.367
R1514 B.n223 B.n222 163.367
R1515 B.n227 B.n226 163.367
R1516 B.n231 B.n230 163.367
R1517 B.n235 B.n234 163.367
R1518 B.n239 B.n238 163.367
R1519 B.n243 B.n242 163.367
R1520 B.n247 B.n246 163.367
R1521 B.n251 B.n250 163.367
R1522 B.n255 B.n254 163.367
R1523 B.n259 B.n258 163.367
R1524 B.n263 B.n262 163.367
R1525 B.n267 B.n266 163.367
R1526 B.n271 B.n270 163.367
R1527 B.n275 B.n274 163.367
R1528 B.n277 B.n116 163.367
R1529 B.n562 B.n357 103.59
R1530 B.n744 B.n743 103.59
R1531 B.n405 B.n404 72.9217
R1532 B.n402 B.n401 72.9217
R1533 B.n120 B.n119 72.9217
R1534 B.n118 B.n117 72.9217
R1535 B.n561 B.n560 71.676
R1536 B.n555 B.n361 71.676
R1537 B.n552 B.n362 71.676
R1538 B.n548 B.n363 71.676
R1539 B.n544 B.n364 71.676
R1540 B.n540 B.n365 71.676
R1541 B.n536 B.n366 71.676
R1542 B.n532 B.n367 71.676
R1543 B.n528 B.n368 71.676
R1544 B.n524 B.n369 71.676
R1545 B.n520 B.n370 71.676
R1546 B.n516 B.n371 71.676
R1547 B.n512 B.n372 71.676
R1548 B.n508 B.n373 71.676
R1549 B.n504 B.n374 71.676
R1550 B.n500 B.n375 71.676
R1551 B.n496 B.n376 71.676
R1552 B.n492 B.n377 71.676
R1553 B.n488 B.n378 71.676
R1554 B.n484 B.n379 71.676
R1555 B.n480 B.n380 71.676
R1556 B.n476 B.n381 71.676
R1557 B.n472 B.n382 71.676
R1558 B.n468 B.n383 71.676
R1559 B.n464 B.n384 71.676
R1560 B.n460 B.n385 71.676
R1561 B.n456 B.n386 71.676
R1562 B.n452 B.n387 71.676
R1563 B.n448 B.n388 71.676
R1564 B.n444 B.n389 71.676
R1565 B.n440 B.n390 71.676
R1566 B.n436 B.n391 71.676
R1567 B.n432 B.n392 71.676
R1568 B.n428 B.n393 71.676
R1569 B.n424 B.n394 71.676
R1570 B.n420 B.n395 71.676
R1571 B.n416 B.n396 71.676
R1572 B.n412 B.n397 71.676
R1573 B.n408 B.n398 71.676
R1574 B.n121 B.n77 71.676
R1575 B.n125 B.n78 71.676
R1576 B.n129 B.n79 71.676
R1577 B.n133 B.n80 71.676
R1578 B.n137 B.n81 71.676
R1579 B.n141 B.n82 71.676
R1580 B.n145 B.n83 71.676
R1581 B.n149 B.n84 71.676
R1582 B.n153 B.n85 71.676
R1583 B.n157 B.n86 71.676
R1584 B.n161 B.n87 71.676
R1585 B.n165 B.n88 71.676
R1586 B.n169 B.n89 71.676
R1587 B.n173 B.n90 71.676
R1588 B.n177 B.n91 71.676
R1589 B.n181 B.n92 71.676
R1590 B.n185 B.n93 71.676
R1591 B.n189 B.n94 71.676
R1592 B.n194 B.n95 71.676
R1593 B.n198 B.n96 71.676
R1594 B.n202 B.n97 71.676
R1595 B.n206 B.n98 71.676
R1596 B.n210 B.n99 71.676
R1597 B.n215 B.n100 71.676
R1598 B.n219 B.n101 71.676
R1599 B.n223 B.n102 71.676
R1600 B.n227 B.n103 71.676
R1601 B.n231 B.n104 71.676
R1602 B.n235 B.n105 71.676
R1603 B.n239 B.n106 71.676
R1604 B.n243 B.n107 71.676
R1605 B.n247 B.n108 71.676
R1606 B.n251 B.n109 71.676
R1607 B.n255 B.n110 71.676
R1608 B.n259 B.n111 71.676
R1609 B.n263 B.n112 71.676
R1610 B.n267 B.n113 71.676
R1611 B.n271 B.n114 71.676
R1612 B.n275 B.n115 71.676
R1613 B.n742 B.n116 71.676
R1614 B.n742 B.n741 71.676
R1615 B.n277 B.n115 71.676
R1616 B.n274 B.n114 71.676
R1617 B.n270 B.n113 71.676
R1618 B.n266 B.n112 71.676
R1619 B.n262 B.n111 71.676
R1620 B.n258 B.n110 71.676
R1621 B.n254 B.n109 71.676
R1622 B.n250 B.n108 71.676
R1623 B.n246 B.n107 71.676
R1624 B.n242 B.n106 71.676
R1625 B.n238 B.n105 71.676
R1626 B.n234 B.n104 71.676
R1627 B.n230 B.n103 71.676
R1628 B.n226 B.n102 71.676
R1629 B.n222 B.n101 71.676
R1630 B.n218 B.n100 71.676
R1631 B.n214 B.n99 71.676
R1632 B.n209 B.n98 71.676
R1633 B.n205 B.n97 71.676
R1634 B.n201 B.n96 71.676
R1635 B.n197 B.n95 71.676
R1636 B.n193 B.n94 71.676
R1637 B.n188 B.n93 71.676
R1638 B.n184 B.n92 71.676
R1639 B.n180 B.n91 71.676
R1640 B.n176 B.n90 71.676
R1641 B.n172 B.n89 71.676
R1642 B.n168 B.n88 71.676
R1643 B.n164 B.n87 71.676
R1644 B.n160 B.n86 71.676
R1645 B.n156 B.n85 71.676
R1646 B.n152 B.n84 71.676
R1647 B.n148 B.n83 71.676
R1648 B.n144 B.n82 71.676
R1649 B.n140 B.n81 71.676
R1650 B.n136 B.n80 71.676
R1651 B.n132 B.n79 71.676
R1652 B.n128 B.n78 71.676
R1653 B.n124 B.n77 71.676
R1654 B.n561 B.n400 71.676
R1655 B.n553 B.n361 71.676
R1656 B.n549 B.n362 71.676
R1657 B.n545 B.n363 71.676
R1658 B.n541 B.n364 71.676
R1659 B.n537 B.n365 71.676
R1660 B.n533 B.n366 71.676
R1661 B.n529 B.n367 71.676
R1662 B.n525 B.n368 71.676
R1663 B.n521 B.n369 71.676
R1664 B.n517 B.n370 71.676
R1665 B.n513 B.n371 71.676
R1666 B.n509 B.n372 71.676
R1667 B.n505 B.n373 71.676
R1668 B.n501 B.n374 71.676
R1669 B.n497 B.n375 71.676
R1670 B.n493 B.n376 71.676
R1671 B.n489 B.n377 71.676
R1672 B.n485 B.n378 71.676
R1673 B.n481 B.n379 71.676
R1674 B.n477 B.n380 71.676
R1675 B.n473 B.n381 71.676
R1676 B.n469 B.n382 71.676
R1677 B.n465 B.n383 71.676
R1678 B.n461 B.n384 71.676
R1679 B.n457 B.n385 71.676
R1680 B.n453 B.n386 71.676
R1681 B.n449 B.n387 71.676
R1682 B.n445 B.n388 71.676
R1683 B.n441 B.n389 71.676
R1684 B.n437 B.n390 71.676
R1685 B.n433 B.n391 71.676
R1686 B.n429 B.n392 71.676
R1687 B.n425 B.n393 71.676
R1688 B.n421 B.n394 71.676
R1689 B.n417 B.n395 71.676
R1690 B.n413 B.n396 71.676
R1691 B.n409 B.n397 71.676
R1692 B.n398 B.n360 71.676
R1693 B.n406 B.n405 59.5399
R1694 B.n403 B.n402 59.5399
R1695 B.n191 B.n120 59.5399
R1696 B.n212 B.n118 59.5399
R1697 B.n568 B.n357 49.2596
R1698 B.n568 B.n353 49.2596
R1699 B.n574 B.n353 49.2596
R1700 B.n574 B.n349 49.2596
R1701 B.n580 B.n349 49.2596
R1702 B.n580 B.n344 49.2596
R1703 B.n586 B.n344 49.2596
R1704 B.n586 B.n345 49.2596
R1705 B.n592 B.n337 49.2596
R1706 B.n598 B.n337 49.2596
R1707 B.n598 B.n333 49.2596
R1708 B.n604 B.n333 49.2596
R1709 B.n604 B.n329 49.2596
R1710 B.n610 B.n329 49.2596
R1711 B.n610 B.n325 49.2596
R1712 B.n616 B.n325 49.2596
R1713 B.n616 B.n321 49.2596
R1714 B.n622 B.n321 49.2596
R1715 B.n622 B.n317 49.2596
R1716 B.n629 B.n317 49.2596
R1717 B.n629 B.n628 49.2596
R1718 B.n635 B.n310 49.2596
R1719 B.n641 B.n310 49.2596
R1720 B.n641 B.n306 49.2596
R1721 B.n647 B.n306 49.2596
R1722 B.n647 B.n302 49.2596
R1723 B.n653 B.n302 49.2596
R1724 B.n653 B.n298 49.2596
R1725 B.n659 B.n298 49.2596
R1726 B.n659 B.n294 49.2596
R1727 B.n665 B.n294 49.2596
R1728 B.n671 B.n290 49.2596
R1729 B.n671 B.n286 49.2596
R1730 B.n678 B.n286 49.2596
R1731 B.n678 B.n282 49.2596
R1732 B.n684 B.n282 49.2596
R1733 B.n684 B.n4 49.2596
R1734 B.n825 B.n4 49.2596
R1735 B.n825 B.n824 49.2596
R1736 B.n824 B.n823 49.2596
R1737 B.n823 B.n8 49.2596
R1738 B.n817 B.n8 49.2596
R1739 B.n817 B.n816 49.2596
R1740 B.n816 B.n815 49.2596
R1741 B.n815 B.n15 49.2596
R1742 B.n809 B.n808 49.2596
R1743 B.n808 B.n807 49.2596
R1744 B.n807 B.n22 49.2596
R1745 B.n801 B.n22 49.2596
R1746 B.n801 B.n800 49.2596
R1747 B.n800 B.n799 49.2596
R1748 B.n799 B.n29 49.2596
R1749 B.n793 B.n29 49.2596
R1750 B.n793 B.n792 49.2596
R1751 B.n792 B.n791 49.2596
R1752 B.n785 B.n39 49.2596
R1753 B.n785 B.n784 49.2596
R1754 B.n784 B.n783 49.2596
R1755 B.n783 B.n43 49.2596
R1756 B.n777 B.n43 49.2596
R1757 B.n777 B.n776 49.2596
R1758 B.n776 B.n775 49.2596
R1759 B.n775 B.n50 49.2596
R1760 B.n769 B.n50 49.2596
R1761 B.n769 B.n768 49.2596
R1762 B.n768 B.n767 49.2596
R1763 B.n767 B.n57 49.2596
R1764 B.n761 B.n57 49.2596
R1765 B.n760 B.n759 49.2596
R1766 B.n759 B.n64 49.2596
R1767 B.n753 B.n64 49.2596
R1768 B.n753 B.n752 49.2596
R1769 B.n752 B.n751 49.2596
R1770 B.n751 B.n71 49.2596
R1771 B.n745 B.n71 49.2596
R1772 B.n745 B.n744 49.2596
R1773 B.n665 B.t3 42.74
R1774 B.n809 B.t0 42.74
R1775 B.n628 B.t1 39.8424
R1776 B.n39 B.t2 39.8424
R1777 B.n122 B.n73 38.2444
R1778 B.n740 B.n739 38.2444
R1779 B.n565 B.n564 38.2444
R1780 B.n559 B.n355 38.2444
R1781 B.n345 B.t9 26.8033
R1782 B.t5 B.n760 26.8033
R1783 B.n592 B.t9 22.4569
R1784 B.n761 B.t5 22.4569
R1785 B B.n827 18.0485
R1786 B.n123 B.n122 10.6151
R1787 B.n126 B.n123 10.6151
R1788 B.n127 B.n126 10.6151
R1789 B.n130 B.n127 10.6151
R1790 B.n131 B.n130 10.6151
R1791 B.n134 B.n131 10.6151
R1792 B.n135 B.n134 10.6151
R1793 B.n138 B.n135 10.6151
R1794 B.n139 B.n138 10.6151
R1795 B.n142 B.n139 10.6151
R1796 B.n143 B.n142 10.6151
R1797 B.n146 B.n143 10.6151
R1798 B.n147 B.n146 10.6151
R1799 B.n150 B.n147 10.6151
R1800 B.n151 B.n150 10.6151
R1801 B.n154 B.n151 10.6151
R1802 B.n155 B.n154 10.6151
R1803 B.n158 B.n155 10.6151
R1804 B.n159 B.n158 10.6151
R1805 B.n162 B.n159 10.6151
R1806 B.n163 B.n162 10.6151
R1807 B.n166 B.n163 10.6151
R1808 B.n167 B.n166 10.6151
R1809 B.n170 B.n167 10.6151
R1810 B.n171 B.n170 10.6151
R1811 B.n174 B.n171 10.6151
R1812 B.n175 B.n174 10.6151
R1813 B.n178 B.n175 10.6151
R1814 B.n179 B.n178 10.6151
R1815 B.n182 B.n179 10.6151
R1816 B.n183 B.n182 10.6151
R1817 B.n186 B.n183 10.6151
R1818 B.n187 B.n186 10.6151
R1819 B.n190 B.n187 10.6151
R1820 B.n195 B.n192 10.6151
R1821 B.n196 B.n195 10.6151
R1822 B.n199 B.n196 10.6151
R1823 B.n200 B.n199 10.6151
R1824 B.n203 B.n200 10.6151
R1825 B.n204 B.n203 10.6151
R1826 B.n207 B.n204 10.6151
R1827 B.n208 B.n207 10.6151
R1828 B.n211 B.n208 10.6151
R1829 B.n216 B.n213 10.6151
R1830 B.n217 B.n216 10.6151
R1831 B.n220 B.n217 10.6151
R1832 B.n221 B.n220 10.6151
R1833 B.n224 B.n221 10.6151
R1834 B.n225 B.n224 10.6151
R1835 B.n228 B.n225 10.6151
R1836 B.n229 B.n228 10.6151
R1837 B.n232 B.n229 10.6151
R1838 B.n233 B.n232 10.6151
R1839 B.n236 B.n233 10.6151
R1840 B.n237 B.n236 10.6151
R1841 B.n240 B.n237 10.6151
R1842 B.n241 B.n240 10.6151
R1843 B.n244 B.n241 10.6151
R1844 B.n245 B.n244 10.6151
R1845 B.n248 B.n245 10.6151
R1846 B.n249 B.n248 10.6151
R1847 B.n252 B.n249 10.6151
R1848 B.n253 B.n252 10.6151
R1849 B.n256 B.n253 10.6151
R1850 B.n257 B.n256 10.6151
R1851 B.n260 B.n257 10.6151
R1852 B.n261 B.n260 10.6151
R1853 B.n264 B.n261 10.6151
R1854 B.n265 B.n264 10.6151
R1855 B.n268 B.n265 10.6151
R1856 B.n269 B.n268 10.6151
R1857 B.n272 B.n269 10.6151
R1858 B.n273 B.n272 10.6151
R1859 B.n276 B.n273 10.6151
R1860 B.n278 B.n276 10.6151
R1861 B.n279 B.n278 10.6151
R1862 B.n740 B.n279 10.6151
R1863 B.n566 B.n565 10.6151
R1864 B.n566 B.n351 10.6151
R1865 B.n576 B.n351 10.6151
R1866 B.n577 B.n576 10.6151
R1867 B.n578 B.n577 10.6151
R1868 B.n578 B.n342 10.6151
R1869 B.n588 B.n342 10.6151
R1870 B.n589 B.n588 10.6151
R1871 B.n590 B.n589 10.6151
R1872 B.n590 B.n335 10.6151
R1873 B.n600 B.n335 10.6151
R1874 B.n601 B.n600 10.6151
R1875 B.n602 B.n601 10.6151
R1876 B.n602 B.n327 10.6151
R1877 B.n612 B.n327 10.6151
R1878 B.n613 B.n612 10.6151
R1879 B.n614 B.n613 10.6151
R1880 B.n614 B.n319 10.6151
R1881 B.n624 B.n319 10.6151
R1882 B.n625 B.n624 10.6151
R1883 B.n626 B.n625 10.6151
R1884 B.n626 B.n312 10.6151
R1885 B.n637 B.n312 10.6151
R1886 B.n638 B.n637 10.6151
R1887 B.n639 B.n638 10.6151
R1888 B.n639 B.n304 10.6151
R1889 B.n649 B.n304 10.6151
R1890 B.n650 B.n649 10.6151
R1891 B.n651 B.n650 10.6151
R1892 B.n651 B.n296 10.6151
R1893 B.n661 B.n296 10.6151
R1894 B.n662 B.n661 10.6151
R1895 B.n663 B.n662 10.6151
R1896 B.n663 B.n288 10.6151
R1897 B.n673 B.n288 10.6151
R1898 B.n674 B.n673 10.6151
R1899 B.n676 B.n674 10.6151
R1900 B.n676 B.n675 10.6151
R1901 B.n675 B.n280 10.6151
R1902 B.n687 B.n280 10.6151
R1903 B.n688 B.n687 10.6151
R1904 B.n689 B.n688 10.6151
R1905 B.n690 B.n689 10.6151
R1906 B.n692 B.n690 10.6151
R1907 B.n693 B.n692 10.6151
R1908 B.n694 B.n693 10.6151
R1909 B.n695 B.n694 10.6151
R1910 B.n697 B.n695 10.6151
R1911 B.n698 B.n697 10.6151
R1912 B.n699 B.n698 10.6151
R1913 B.n700 B.n699 10.6151
R1914 B.n702 B.n700 10.6151
R1915 B.n703 B.n702 10.6151
R1916 B.n704 B.n703 10.6151
R1917 B.n705 B.n704 10.6151
R1918 B.n707 B.n705 10.6151
R1919 B.n708 B.n707 10.6151
R1920 B.n709 B.n708 10.6151
R1921 B.n710 B.n709 10.6151
R1922 B.n712 B.n710 10.6151
R1923 B.n713 B.n712 10.6151
R1924 B.n714 B.n713 10.6151
R1925 B.n715 B.n714 10.6151
R1926 B.n717 B.n715 10.6151
R1927 B.n718 B.n717 10.6151
R1928 B.n719 B.n718 10.6151
R1929 B.n720 B.n719 10.6151
R1930 B.n722 B.n720 10.6151
R1931 B.n723 B.n722 10.6151
R1932 B.n724 B.n723 10.6151
R1933 B.n725 B.n724 10.6151
R1934 B.n727 B.n725 10.6151
R1935 B.n728 B.n727 10.6151
R1936 B.n729 B.n728 10.6151
R1937 B.n730 B.n729 10.6151
R1938 B.n732 B.n730 10.6151
R1939 B.n733 B.n732 10.6151
R1940 B.n734 B.n733 10.6151
R1941 B.n735 B.n734 10.6151
R1942 B.n737 B.n735 10.6151
R1943 B.n738 B.n737 10.6151
R1944 B.n739 B.n738 10.6151
R1945 B.n559 B.n558 10.6151
R1946 B.n558 B.n557 10.6151
R1947 B.n557 B.n556 10.6151
R1948 B.n556 B.n554 10.6151
R1949 B.n554 B.n551 10.6151
R1950 B.n551 B.n550 10.6151
R1951 B.n550 B.n547 10.6151
R1952 B.n547 B.n546 10.6151
R1953 B.n546 B.n543 10.6151
R1954 B.n543 B.n542 10.6151
R1955 B.n542 B.n539 10.6151
R1956 B.n539 B.n538 10.6151
R1957 B.n538 B.n535 10.6151
R1958 B.n535 B.n534 10.6151
R1959 B.n534 B.n531 10.6151
R1960 B.n531 B.n530 10.6151
R1961 B.n530 B.n527 10.6151
R1962 B.n527 B.n526 10.6151
R1963 B.n526 B.n523 10.6151
R1964 B.n523 B.n522 10.6151
R1965 B.n522 B.n519 10.6151
R1966 B.n519 B.n518 10.6151
R1967 B.n518 B.n515 10.6151
R1968 B.n515 B.n514 10.6151
R1969 B.n514 B.n511 10.6151
R1970 B.n511 B.n510 10.6151
R1971 B.n510 B.n507 10.6151
R1972 B.n507 B.n506 10.6151
R1973 B.n506 B.n503 10.6151
R1974 B.n503 B.n502 10.6151
R1975 B.n502 B.n499 10.6151
R1976 B.n499 B.n498 10.6151
R1977 B.n498 B.n495 10.6151
R1978 B.n495 B.n494 10.6151
R1979 B.n491 B.n490 10.6151
R1980 B.n490 B.n487 10.6151
R1981 B.n487 B.n486 10.6151
R1982 B.n486 B.n483 10.6151
R1983 B.n483 B.n482 10.6151
R1984 B.n482 B.n479 10.6151
R1985 B.n479 B.n478 10.6151
R1986 B.n478 B.n475 10.6151
R1987 B.n475 B.n474 10.6151
R1988 B.n471 B.n470 10.6151
R1989 B.n470 B.n467 10.6151
R1990 B.n467 B.n466 10.6151
R1991 B.n466 B.n463 10.6151
R1992 B.n463 B.n462 10.6151
R1993 B.n462 B.n459 10.6151
R1994 B.n459 B.n458 10.6151
R1995 B.n458 B.n455 10.6151
R1996 B.n455 B.n454 10.6151
R1997 B.n454 B.n451 10.6151
R1998 B.n451 B.n450 10.6151
R1999 B.n450 B.n447 10.6151
R2000 B.n447 B.n446 10.6151
R2001 B.n446 B.n443 10.6151
R2002 B.n443 B.n442 10.6151
R2003 B.n442 B.n439 10.6151
R2004 B.n439 B.n438 10.6151
R2005 B.n438 B.n435 10.6151
R2006 B.n435 B.n434 10.6151
R2007 B.n434 B.n431 10.6151
R2008 B.n431 B.n430 10.6151
R2009 B.n430 B.n427 10.6151
R2010 B.n427 B.n426 10.6151
R2011 B.n426 B.n423 10.6151
R2012 B.n423 B.n422 10.6151
R2013 B.n422 B.n419 10.6151
R2014 B.n419 B.n418 10.6151
R2015 B.n418 B.n415 10.6151
R2016 B.n415 B.n414 10.6151
R2017 B.n414 B.n411 10.6151
R2018 B.n411 B.n410 10.6151
R2019 B.n410 B.n407 10.6151
R2020 B.n407 B.n359 10.6151
R2021 B.n564 B.n359 10.6151
R2022 B.n570 B.n355 10.6151
R2023 B.n571 B.n570 10.6151
R2024 B.n572 B.n571 10.6151
R2025 B.n572 B.n347 10.6151
R2026 B.n582 B.n347 10.6151
R2027 B.n583 B.n582 10.6151
R2028 B.n584 B.n583 10.6151
R2029 B.n584 B.n339 10.6151
R2030 B.n594 B.n339 10.6151
R2031 B.n595 B.n594 10.6151
R2032 B.n596 B.n595 10.6151
R2033 B.n596 B.n331 10.6151
R2034 B.n606 B.n331 10.6151
R2035 B.n607 B.n606 10.6151
R2036 B.n608 B.n607 10.6151
R2037 B.n608 B.n323 10.6151
R2038 B.n618 B.n323 10.6151
R2039 B.n619 B.n618 10.6151
R2040 B.n620 B.n619 10.6151
R2041 B.n620 B.n315 10.6151
R2042 B.n631 B.n315 10.6151
R2043 B.n632 B.n631 10.6151
R2044 B.n633 B.n632 10.6151
R2045 B.n633 B.n308 10.6151
R2046 B.n643 B.n308 10.6151
R2047 B.n644 B.n643 10.6151
R2048 B.n645 B.n644 10.6151
R2049 B.n645 B.n300 10.6151
R2050 B.n655 B.n300 10.6151
R2051 B.n656 B.n655 10.6151
R2052 B.n657 B.n656 10.6151
R2053 B.n657 B.n292 10.6151
R2054 B.n667 B.n292 10.6151
R2055 B.n668 B.n667 10.6151
R2056 B.n669 B.n668 10.6151
R2057 B.n669 B.n284 10.6151
R2058 B.n680 B.n284 10.6151
R2059 B.n681 B.n680 10.6151
R2060 B.n682 B.n681 10.6151
R2061 B.n682 B.n0 10.6151
R2062 B.n821 B.n1 10.6151
R2063 B.n821 B.n820 10.6151
R2064 B.n820 B.n819 10.6151
R2065 B.n819 B.n10 10.6151
R2066 B.n813 B.n10 10.6151
R2067 B.n813 B.n812 10.6151
R2068 B.n812 B.n811 10.6151
R2069 B.n811 B.n17 10.6151
R2070 B.n805 B.n17 10.6151
R2071 B.n805 B.n804 10.6151
R2072 B.n804 B.n803 10.6151
R2073 B.n803 B.n24 10.6151
R2074 B.n797 B.n24 10.6151
R2075 B.n797 B.n796 10.6151
R2076 B.n796 B.n795 10.6151
R2077 B.n795 B.n31 10.6151
R2078 B.n789 B.n31 10.6151
R2079 B.n789 B.n788 10.6151
R2080 B.n788 B.n787 10.6151
R2081 B.n787 B.n37 10.6151
R2082 B.n781 B.n37 10.6151
R2083 B.n781 B.n780 10.6151
R2084 B.n780 B.n779 10.6151
R2085 B.n779 B.n45 10.6151
R2086 B.n773 B.n45 10.6151
R2087 B.n773 B.n772 10.6151
R2088 B.n772 B.n771 10.6151
R2089 B.n771 B.n52 10.6151
R2090 B.n765 B.n52 10.6151
R2091 B.n765 B.n764 10.6151
R2092 B.n764 B.n763 10.6151
R2093 B.n763 B.n59 10.6151
R2094 B.n757 B.n59 10.6151
R2095 B.n757 B.n756 10.6151
R2096 B.n756 B.n755 10.6151
R2097 B.n755 B.n66 10.6151
R2098 B.n749 B.n66 10.6151
R2099 B.n749 B.n748 10.6151
R2100 B.n748 B.n747 10.6151
R2101 B.n747 B.n73 10.6151
R2102 B.n635 B.t1 9.41769
R2103 B.n791 B.t2 9.41769
R2104 B.n191 B.n190 9.36635
R2105 B.n213 B.n212 9.36635
R2106 B.n494 B.n403 9.36635
R2107 B.n471 B.n406 9.36635
R2108 B.t3 B.n290 6.52009
R2109 B.t0 B.n15 6.52009
R2110 B.n827 B.n0 2.81026
R2111 B.n827 B.n1 2.81026
R2112 B.n192 B.n191 1.24928
R2113 B.n212 B.n211 1.24928
R2114 B.n491 B.n403 1.24928
R2115 B.n474 B.n406 1.24928
R2116 VN.n0 VN.t3 103.716
R2117 VN.n1 VN.t2 103.716
R2118 VN.n0 VN.t0 102.513
R2119 VN.n1 VN.t1 102.513
R2120 VN VN.n1 49.6867
R2121 VN VN.n0 2.27384
R2122 VDD2.n2 VDD2.n0 103.653
R2123 VDD2.n2 VDD2.n1 61.6705
R2124 VDD2.n1 VDD2.t2 1.99848
R2125 VDD2.n1 VDD2.t1 1.99848
R2126 VDD2.n0 VDD2.t0 1.99848
R2127 VDD2.n0 VDD2.t3 1.99848
R2128 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.149899f
C1 VDD2 VN 4.1525f
C2 VDD1 VP 4.44892f
C3 VP VDD2 0.447269f
C4 VDD1 VTAIL 5.16758f
C5 VTAIL VDD2 5.22735f
C6 VDD1 VDD2 1.22333f
C7 VP VN 6.40639f
C8 VTAIL VN 4.28709f
C9 VTAIL VP 4.3012f
C10 VDD2 B 4.087603f
C11 VDD1 B 8.331511f
C12 VTAIL B 9.268354f
C13 VN B 12.16697f
C14 VP B 10.570698f
C15 VDD2.t0 B 0.215005f
C16 VDD2.t3 B 0.215005f
C17 VDD2.n0 B 2.54847f
C18 VDD2.t2 B 0.215005f
C19 VDD2.t1 B 0.215005f
C20 VDD2.n1 B 1.8909f
C21 VDD2.n2 B 3.80795f
C22 VN.t0 B 2.31523f
C23 VN.t3 B 2.32522f
C24 VN.n0 B 1.39939f
C25 VN.t2 B 2.32522f
C26 VN.t1 B 2.31523f
C27 VN.n1 B 2.73705f
C28 VTAIL.n0 B 0.022873f
C29 VTAIL.n1 B 0.017719f
C30 VTAIL.n2 B 0.009521f
C31 VTAIL.n3 B 0.022505f
C32 VTAIL.n4 B 0.010082f
C33 VTAIL.n5 B 0.017719f
C34 VTAIL.n6 B 0.009801f
C35 VTAIL.n7 B 0.022505f
C36 VTAIL.n8 B 0.010082f
C37 VTAIL.n9 B 0.017719f
C38 VTAIL.n10 B 0.009521f
C39 VTAIL.n11 B 0.022505f
C40 VTAIL.n12 B 0.010082f
C41 VTAIL.n13 B 0.017719f
C42 VTAIL.n14 B 0.009521f
C43 VTAIL.n15 B 0.016879f
C44 VTAIL.n16 B 0.015909f
C45 VTAIL.t0 B 0.037811f
C46 VTAIL.n17 B 0.113536f
C47 VTAIL.n18 B 0.729171f
C48 VTAIL.n19 B 0.009521f
C49 VTAIL.n20 B 0.010082f
C50 VTAIL.n21 B 0.022505f
C51 VTAIL.n22 B 0.022505f
C52 VTAIL.n23 B 0.010082f
C53 VTAIL.n24 B 0.009521f
C54 VTAIL.n25 B 0.017719f
C55 VTAIL.n26 B 0.017719f
C56 VTAIL.n27 B 0.009521f
C57 VTAIL.n28 B 0.010082f
C58 VTAIL.n29 B 0.022505f
C59 VTAIL.n30 B 0.022505f
C60 VTAIL.n31 B 0.010082f
C61 VTAIL.n32 B 0.009521f
C62 VTAIL.n33 B 0.017719f
C63 VTAIL.n34 B 0.017719f
C64 VTAIL.n35 B 0.009521f
C65 VTAIL.n36 B 0.009521f
C66 VTAIL.n37 B 0.010082f
C67 VTAIL.n38 B 0.022505f
C68 VTAIL.n39 B 0.022505f
C69 VTAIL.n40 B 0.022505f
C70 VTAIL.n41 B 0.009801f
C71 VTAIL.n42 B 0.009521f
C72 VTAIL.n43 B 0.017719f
C73 VTAIL.n44 B 0.017719f
C74 VTAIL.n45 B 0.009521f
C75 VTAIL.n46 B 0.010082f
C76 VTAIL.n47 B 0.022505f
C77 VTAIL.n48 B 0.045126f
C78 VTAIL.n49 B 0.010082f
C79 VTAIL.n50 B 0.009521f
C80 VTAIL.n51 B 0.039746f
C81 VTAIL.n52 B 0.024843f
C82 VTAIL.n53 B 0.13713f
C83 VTAIL.n54 B 0.022873f
C84 VTAIL.n55 B 0.017719f
C85 VTAIL.n56 B 0.009521f
C86 VTAIL.n57 B 0.022505f
C87 VTAIL.n58 B 0.010082f
C88 VTAIL.n59 B 0.017719f
C89 VTAIL.n60 B 0.009801f
C90 VTAIL.n61 B 0.022505f
C91 VTAIL.n62 B 0.010082f
C92 VTAIL.n63 B 0.017719f
C93 VTAIL.n64 B 0.009521f
C94 VTAIL.n65 B 0.022505f
C95 VTAIL.n66 B 0.010082f
C96 VTAIL.n67 B 0.017719f
C97 VTAIL.n68 B 0.009521f
C98 VTAIL.n69 B 0.016879f
C99 VTAIL.n70 B 0.015909f
C100 VTAIL.t3 B 0.037811f
C101 VTAIL.n71 B 0.113536f
C102 VTAIL.n72 B 0.729171f
C103 VTAIL.n73 B 0.009521f
C104 VTAIL.n74 B 0.010082f
C105 VTAIL.n75 B 0.022505f
C106 VTAIL.n76 B 0.022505f
C107 VTAIL.n77 B 0.010082f
C108 VTAIL.n78 B 0.009521f
C109 VTAIL.n79 B 0.017719f
C110 VTAIL.n80 B 0.017719f
C111 VTAIL.n81 B 0.009521f
C112 VTAIL.n82 B 0.010082f
C113 VTAIL.n83 B 0.022505f
C114 VTAIL.n84 B 0.022505f
C115 VTAIL.n85 B 0.010082f
C116 VTAIL.n86 B 0.009521f
C117 VTAIL.n87 B 0.017719f
C118 VTAIL.n88 B 0.017719f
C119 VTAIL.n89 B 0.009521f
C120 VTAIL.n90 B 0.009521f
C121 VTAIL.n91 B 0.010082f
C122 VTAIL.n92 B 0.022505f
C123 VTAIL.n93 B 0.022505f
C124 VTAIL.n94 B 0.022505f
C125 VTAIL.n95 B 0.009801f
C126 VTAIL.n96 B 0.009521f
C127 VTAIL.n97 B 0.017719f
C128 VTAIL.n98 B 0.017719f
C129 VTAIL.n99 B 0.009521f
C130 VTAIL.n100 B 0.010082f
C131 VTAIL.n101 B 0.022505f
C132 VTAIL.n102 B 0.045126f
C133 VTAIL.n103 B 0.010082f
C134 VTAIL.n104 B 0.009521f
C135 VTAIL.n105 B 0.039746f
C136 VTAIL.n106 B 0.024843f
C137 VTAIL.n107 B 0.22634f
C138 VTAIL.n108 B 0.022873f
C139 VTAIL.n109 B 0.017719f
C140 VTAIL.n110 B 0.009521f
C141 VTAIL.n111 B 0.022505f
C142 VTAIL.n112 B 0.010082f
C143 VTAIL.n113 B 0.017719f
C144 VTAIL.n114 B 0.009801f
C145 VTAIL.n115 B 0.022505f
C146 VTAIL.n116 B 0.010082f
C147 VTAIL.n117 B 0.017719f
C148 VTAIL.n118 B 0.009521f
C149 VTAIL.n119 B 0.022505f
C150 VTAIL.n120 B 0.010082f
C151 VTAIL.n121 B 0.017719f
C152 VTAIL.n122 B 0.009521f
C153 VTAIL.n123 B 0.016879f
C154 VTAIL.n124 B 0.015909f
C155 VTAIL.t1 B 0.037811f
C156 VTAIL.n125 B 0.113536f
C157 VTAIL.n126 B 0.729171f
C158 VTAIL.n127 B 0.009521f
C159 VTAIL.n128 B 0.010082f
C160 VTAIL.n129 B 0.022505f
C161 VTAIL.n130 B 0.022505f
C162 VTAIL.n131 B 0.010082f
C163 VTAIL.n132 B 0.009521f
C164 VTAIL.n133 B 0.017719f
C165 VTAIL.n134 B 0.017719f
C166 VTAIL.n135 B 0.009521f
C167 VTAIL.n136 B 0.010082f
C168 VTAIL.n137 B 0.022505f
C169 VTAIL.n138 B 0.022505f
C170 VTAIL.n139 B 0.010082f
C171 VTAIL.n140 B 0.009521f
C172 VTAIL.n141 B 0.017719f
C173 VTAIL.n142 B 0.017719f
C174 VTAIL.n143 B 0.009521f
C175 VTAIL.n144 B 0.009521f
C176 VTAIL.n145 B 0.010082f
C177 VTAIL.n146 B 0.022505f
C178 VTAIL.n147 B 0.022505f
C179 VTAIL.n148 B 0.022505f
C180 VTAIL.n149 B 0.009801f
C181 VTAIL.n150 B 0.009521f
C182 VTAIL.n151 B 0.017719f
C183 VTAIL.n152 B 0.017719f
C184 VTAIL.n153 B 0.009521f
C185 VTAIL.n154 B 0.010082f
C186 VTAIL.n155 B 0.022505f
C187 VTAIL.n156 B 0.045126f
C188 VTAIL.n157 B 0.010082f
C189 VTAIL.n158 B 0.009521f
C190 VTAIL.n159 B 0.039746f
C191 VTAIL.n160 B 0.024843f
C192 VTAIL.n161 B 1.11303f
C193 VTAIL.n162 B 0.022873f
C194 VTAIL.n163 B 0.017719f
C195 VTAIL.n164 B 0.009521f
C196 VTAIL.n165 B 0.022505f
C197 VTAIL.n166 B 0.010082f
C198 VTAIL.n167 B 0.017719f
C199 VTAIL.n168 B 0.009801f
C200 VTAIL.n169 B 0.022505f
C201 VTAIL.n170 B 0.009521f
C202 VTAIL.n171 B 0.010082f
C203 VTAIL.n172 B 0.017719f
C204 VTAIL.n173 B 0.009521f
C205 VTAIL.n174 B 0.022505f
C206 VTAIL.n175 B 0.010082f
C207 VTAIL.n176 B 0.017719f
C208 VTAIL.n177 B 0.009521f
C209 VTAIL.n178 B 0.016879f
C210 VTAIL.n179 B 0.015909f
C211 VTAIL.t6 B 0.037811f
C212 VTAIL.n180 B 0.113536f
C213 VTAIL.n181 B 0.729171f
C214 VTAIL.n182 B 0.009521f
C215 VTAIL.n183 B 0.010082f
C216 VTAIL.n184 B 0.022505f
C217 VTAIL.n185 B 0.022505f
C218 VTAIL.n186 B 0.010082f
C219 VTAIL.n187 B 0.009521f
C220 VTAIL.n188 B 0.017719f
C221 VTAIL.n189 B 0.017719f
C222 VTAIL.n190 B 0.009521f
C223 VTAIL.n191 B 0.010082f
C224 VTAIL.n192 B 0.022505f
C225 VTAIL.n193 B 0.022505f
C226 VTAIL.n194 B 0.010082f
C227 VTAIL.n195 B 0.009521f
C228 VTAIL.n196 B 0.017719f
C229 VTAIL.n197 B 0.017719f
C230 VTAIL.n198 B 0.009521f
C231 VTAIL.n199 B 0.010082f
C232 VTAIL.n200 B 0.022505f
C233 VTAIL.n201 B 0.022505f
C234 VTAIL.n202 B 0.022505f
C235 VTAIL.n203 B 0.009801f
C236 VTAIL.n204 B 0.009521f
C237 VTAIL.n205 B 0.017719f
C238 VTAIL.n206 B 0.017719f
C239 VTAIL.n207 B 0.009521f
C240 VTAIL.n208 B 0.010082f
C241 VTAIL.n209 B 0.022505f
C242 VTAIL.n210 B 0.045126f
C243 VTAIL.n211 B 0.010082f
C244 VTAIL.n212 B 0.009521f
C245 VTAIL.n213 B 0.039746f
C246 VTAIL.n214 B 0.024843f
C247 VTAIL.n215 B 1.11303f
C248 VTAIL.n216 B 0.022873f
C249 VTAIL.n217 B 0.017719f
C250 VTAIL.n218 B 0.009521f
C251 VTAIL.n219 B 0.022505f
C252 VTAIL.n220 B 0.010082f
C253 VTAIL.n221 B 0.017719f
C254 VTAIL.n222 B 0.009801f
C255 VTAIL.n223 B 0.022505f
C256 VTAIL.n224 B 0.009521f
C257 VTAIL.n225 B 0.010082f
C258 VTAIL.n226 B 0.017719f
C259 VTAIL.n227 B 0.009521f
C260 VTAIL.n228 B 0.022505f
C261 VTAIL.n229 B 0.010082f
C262 VTAIL.n230 B 0.017719f
C263 VTAIL.n231 B 0.009521f
C264 VTAIL.n232 B 0.016879f
C265 VTAIL.n233 B 0.015909f
C266 VTAIL.t5 B 0.037811f
C267 VTAIL.n234 B 0.113536f
C268 VTAIL.n235 B 0.729171f
C269 VTAIL.n236 B 0.009521f
C270 VTAIL.n237 B 0.010082f
C271 VTAIL.n238 B 0.022505f
C272 VTAIL.n239 B 0.022505f
C273 VTAIL.n240 B 0.010082f
C274 VTAIL.n241 B 0.009521f
C275 VTAIL.n242 B 0.017719f
C276 VTAIL.n243 B 0.017719f
C277 VTAIL.n244 B 0.009521f
C278 VTAIL.n245 B 0.010082f
C279 VTAIL.n246 B 0.022505f
C280 VTAIL.n247 B 0.022505f
C281 VTAIL.n248 B 0.010082f
C282 VTAIL.n249 B 0.009521f
C283 VTAIL.n250 B 0.017719f
C284 VTAIL.n251 B 0.017719f
C285 VTAIL.n252 B 0.009521f
C286 VTAIL.n253 B 0.010082f
C287 VTAIL.n254 B 0.022505f
C288 VTAIL.n255 B 0.022505f
C289 VTAIL.n256 B 0.022505f
C290 VTAIL.n257 B 0.009801f
C291 VTAIL.n258 B 0.009521f
C292 VTAIL.n259 B 0.017719f
C293 VTAIL.n260 B 0.017719f
C294 VTAIL.n261 B 0.009521f
C295 VTAIL.n262 B 0.010082f
C296 VTAIL.n263 B 0.022505f
C297 VTAIL.n264 B 0.045126f
C298 VTAIL.n265 B 0.010082f
C299 VTAIL.n266 B 0.009521f
C300 VTAIL.n267 B 0.039746f
C301 VTAIL.n268 B 0.024843f
C302 VTAIL.n269 B 0.22634f
C303 VTAIL.n270 B 0.022873f
C304 VTAIL.n271 B 0.017719f
C305 VTAIL.n272 B 0.009521f
C306 VTAIL.n273 B 0.022505f
C307 VTAIL.n274 B 0.010082f
C308 VTAIL.n275 B 0.017719f
C309 VTAIL.n276 B 0.009801f
C310 VTAIL.n277 B 0.022505f
C311 VTAIL.n278 B 0.009521f
C312 VTAIL.n279 B 0.010082f
C313 VTAIL.n280 B 0.017719f
C314 VTAIL.n281 B 0.009521f
C315 VTAIL.n282 B 0.022505f
C316 VTAIL.n283 B 0.010082f
C317 VTAIL.n284 B 0.017719f
C318 VTAIL.n285 B 0.009521f
C319 VTAIL.n286 B 0.016879f
C320 VTAIL.n287 B 0.015909f
C321 VTAIL.t4 B 0.037811f
C322 VTAIL.n288 B 0.113536f
C323 VTAIL.n289 B 0.729171f
C324 VTAIL.n290 B 0.009521f
C325 VTAIL.n291 B 0.010082f
C326 VTAIL.n292 B 0.022505f
C327 VTAIL.n293 B 0.022505f
C328 VTAIL.n294 B 0.010082f
C329 VTAIL.n295 B 0.009521f
C330 VTAIL.n296 B 0.017719f
C331 VTAIL.n297 B 0.017719f
C332 VTAIL.n298 B 0.009521f
C333 VTAIL.n299 B 0.010082f
C334 VTAIL.n300 B 0.022505f
C335 VTAIL.n301 B 0.022505f
C336 VTAIL.n302 B 0.010082f
C337 VTAIL.n303 B 0.009521f
C338 VTAIL.n304 B 0.017719f
C339 VTAIL.n305 B 0.017719f
C340 VTAIL.n306 B 0.009521f
C341 VTAIL.n307 B 0.010082f
C342 VTAIL.n308 B 0.022505f
C343 VTAIL.n309 B 0.022505f
C344 VTAIL.n310 B 0.022505f
C345 VTAIL.n311 B 0.009801f
C346 VTAIL.n312 B 0.009521f
C347 VTAIL.n313 B 0.017719f
C348 VTAIL.n314 B 0.017719f
C349 VTAIL.n315 B 0.009521f
C350 VTAIL.n316 B 0.010082f
C351 VTAIL.n317 B 0.022505f
C352 VTAIL.n318 B 0.045126f
C353 VTAIL.n319 B 0.010082f
C354 VTAIL.n320 B 0.009521f
C355 VTAIL.n321 B 0.039746f
C356 VTAIL.n322 B 0.024843f
C357 VTAIL.n323 B 0.22634f
C358 VTAIL.n324 B 0.022873f
C359 VTAIL.n325 B 0.017719f
C360 VTAIL.n326 B 0.009521f
C361 VTAIL.n327 B 0.022505f
C362 VTAIL.n328 B 0.010082f
C363 VTAIL.n329 B 0.017719f
C364 VTAIL.n330 B 0.009801f
C365 VTAIL.n331 B 0.022505f
C366 VTAIL.n332 B 0.009521f
C367 VTAIL.n333 B 0.010082f
C368 VTAIL.n334 B 0.017719f
C369 VTAIL.n335 B 0.009521f
C370 VTAIL.n336 B 0.022505f
C371 VTAIL.n337 B 0.010082f
C372 VTAIL.n338 B 0.017719f
C373 VTAIL.n339 B 0.009521f
C374 VTAIL.n340 B 0.016879f
C375 VTAIL.n341 B 0.015909f
C376 VTAIL.t2 B 0.037811f
C377 VTAIL.n342 B 0.113536f
C378 VTAIL.n343 B 0.729171f
C379 VTAIL.n344 B 0.009521f
C380 VTAIL.n345 B 0.010082f
C381 VTAIL.n346 B 0.022505f
C382 VTAIL.n347 B 0.022505f
C383 VTAIL.n348 B 0.010082f
C384 VTAIL.n349 B 0.009521f
C385 VTAIL.n350 B 0.017719f
C386 VTAIL.n351 B 0.017719f
C387 VTAIL.n352 B 0.009521f
C388 VTAIL.n353 B 0.010082f
C389 VTAIL.n354 B 0.022505f
C390 VTAIL.n355 B 0.022505f
C391 VTAIL.n356 B 0.010082f
C392 VTAIL.n357 B 0.009521f
C393 VTAIL.n358 B 0.017719f
C394 VTAIL.n359 B 0.017719f
C395 VTAIL.n360 B 0.009521f
C396 VTAIL.n361 B 0.010082f
C397 VTAIL.n362 B 0.022505f
C398 VTAIL.n363 B 0.022505f
C399 VTAIL.n364 B 0.022505f
C400 VTAIL.n365 B 0.009801f
C401 VTAIL.n366 B 0.009521f
C402 VTAIL.n367 B 0.017719f
C403 VTAIL.n368 B 0.017719f
C404 VTAIL.n369 B 0.009521f
C405 VTAIL.n370 B 0.010082f
C406 VTAIL.n371 B 0.022505f
C407 VTAIL.n372 B 0.045126f
C408 VTAIL.n373 B 0.010082f
C409 VTAIL.n374 B 0.009521f
C410 VTAIL.n375 B 0.039746f
C411 VTAIL.n376 B 0.024843f
C412 VTAIL.n377 B 1.11303f
C413 VTAIL.n378 B 0.022873f
C414 VTAIL.n379 B 0.017719f
C415 VTAIL.n380 B 0.009521f
C416 VTAIL.n381 B 0.022505f
C417 VTAIL.n382 B 0.010082f
C418 VTAIL.n383 B 0.017719f
C419 VTAIL.n384 B 0.009801f
C420 VTAIL.n385 B 0.022505f
C421 VTAIL.n386 B 0.010082f
C422 VTAIL.n387 B 0.017719f
C423 VTAIL.n388 B 0.009521f
C424 VTAIL.n389 B 0.022505f
C425 VTAIL.n390 B 0.010082f
C426 VTAIL.n391 B 0.017719f
C427 VTAIL.n392 B 0.009521f
C428 VTAIL.n393 B 0.016879f
C429 VTAIL.n394 B 0.015909f
C430 VTAIL.t7 B 0.037811f
C431 VTAIL.n395 B 0.113536f
C432 VTAIL.n396 B 0.729171f
C433 VTAIL.n397 B 0.009521f
C434 VTAIL.n398 B 0.010082f
C435 VTAIL.n399 B 0.022505f
C436 VTAIL.n400 B 0.022505f
C437 VTAIL.n401 B 0.010082f
C438 VTAIL.n402 B 0.009521f
C439 VTAIL.n403 B 0.017719f
C440 VTAIL.n404 B 0.017719f
C441 VTAIL.n405 B 0.009521f
C442 VTAIL.n406 B 0.010082f
C443 VTAIL.n407 B 0.022505f
C444 VTAIL.n408 B 0.022505f
C445 VTAIL.n409 B 0.010082f
C446 VTAIL.n410 B 0.009521f
C447 VTAIL.n411 B 0.017719f
C448 VTAIL.n412 B 0.017719f
C449 VTAIL.n413 B 0.009521f
C450 VTAIL.n414 B 0.009521f
C451 VTAIL.n415 B 0.010082f
C452 VTAIL.n416 B 0.022505f
C453 VTAIL.n417 B 0.022505f
C454 VTAIL.n418 B 0.022505f
C455 VTAIL.n419 B 0.009801f
C456 VTAIL.n420 B 0.009521f
C457 VTAIL.n421 B 0.017719f
C458 VTAIL.n422 B 0.017719f
C459 VTAIL.n423 B 0.009521f
C460 VTAIL.n424 B 0.010082f
C461 VTAIL.n425 B 0.022505f
C462 VTAIL.n426 B 0.045126f
C463 VTAIL.n427 B 0.010082f
C464 VTAIL.n428 B 0.009521f
C465 VTAIL.n429 B 0.039746f
C466 VTAIL.n430 B 0.024843f
C467 VTAIL.n431 B 1.01718f
C468 VDD1.t0 B 0.217236f
C469 VDD1.t2 B 0.217236f
C470 VDD1.n0 B 1.91102f
C471 VDD1.t1 B 0.217236f
C472 VDD1.t3 B 0.217236f
C473 VDD1.n1 B 2.60227f
C474 VP.t1 B 2.06422f
C475 VP.n0 B 0.813034f
C476 VP.n1 B 0.022424f
C477 VP.n2 B 0.032735f
C478 VP.n3 B 0.022424f
C479 VP.n4 B 0.026524f
C480 VP.t0 B 2.36135f
C481 VP.t2 B 2.3512f
C482 VP.n5 B 2.77041f
C483 VP.t3 B 2.06422f
C484 VP.n6 B 0.813034f
C485 VP.n7 B 1.26632f
C486 VP.n8 B 0.036191f
C487 VP.n9 B 0.022424f
C488 VP.n10 B 0.041792f
C489 VP.n11 B 0.041792f
C490 VP.n12 B 0.032735f
C491 VP.n13 B 0.022424f
C492 VP.n14 B 0.022424f
C493 VP.n15 B 0.022424f
C494 VP.n16 B 0.041792f
C495 VP.n17 B 0.041792f
C496 VP.n18 B 0.026524f
C497 VP.n19 B 0.036191f
C498 VP.n20 B 0.062107f
.ends

