* NGSPICE file created from diff_pair_sample_0420.ext - technology: sky130A

.subckt diff_pair_sample_0420 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t3 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=2.30835 pd=14.32 as=5.4561 ps=28.76 w=13.99 l=1.51
X1 VTAIL.t2 VN.t1 VDD2.t2 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=2.30835 ps=14.32 w=13.99 l=1.51
X2 B.t11 B.t9 B.t10 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=0 ps=0 w=13.99 l=1.51
X3 B.t8 B.t6 B.t7 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=0 ps=0 w=13.99 l=1.51
X4 VDD2.t1 VN.t2 VTAIL.t4 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=2.30835 pd=14.32 as=5.4561 ps=28.76 w=13.99 l=1.51
X5 B.t5 B.t3 B.t4 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=0 ps=0 w=13.99 l=1.51
X6 VTAIL.t5 VN.t3 VDD2.t0 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=2.30835 ps=14.32 w=13.99 l=1.51
X7 VTAIL.t7 VP.t0 VDD1.t3 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=2.30835 ps=14.32 w=13.99 l=1.51
X8 VTAIL.t6 VP.t1 VDD1.t2 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=2.30835 ps=14.32 w=13.99 l=1.51
X9 VDD1.t1 VP.t2 VTAIL.t1 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=2.30835 pd=14.32 as=5.4561 ps=28.76 w=13.99 l=1.51
X10 VDD1.t0 VP.t3 VTAIL.t0 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=2.30835 pd=14.32 as=5.4561 ps=28.76 w=13.99 l=1.51
X11 B.t2 B.t0 B.t1 w_n2074_n3766# sky130_fd_pr__pfet_01v8 ad=5.4561 pd=28.76 as=0 ps=0 w=13.99 l=1.51
R0 VN.n0 VN.t1 259.791
R1 VN.n1 VN.t2 259.791
R2 VN.n0 VN.t0 259.474
R3 VN.n1 VN.t3 259.474
R4 VN VN.n1 57.7753
R5 VN VN.n0 13.029
R6 VTAIL.n618 VTAIL.n546 756.745
R7 VTAIL.n72 VTAIL.n0 756.745
R8 VTAIL.n150 VTAIL.n78 756.745
R9 VTAIL.n228 VTAIL.n156 756.745
R10 VTAIL.n540 VTAIL.n468 756.745
R11 VTAIL.n462 VTAIL.n390 756.745
R12 VTAIL.n384 VTAIL.n312 756.745
R13 VTAIL.n306 VTAIL.n234 756.745
R14 VTAIL.n570 VTAIL.n569 585
R15 VTAIL.n575 VTAIL.n574 585
R16 VTAIL.n577 VTAIL.n576 585
R17 VTAIL.n566 VTAIL.n565 585
R18 VTAIL.n583 VTAIL.n582 585
R19 VTAIL.n585 VTAIL.n584 585
R20 VTAIL.n562 VTAIL.n561 585
R21 VTAIL.n591 VTAIL.n590 585
R22 VTAIL.n593 VTAIL.n592 585
R23 VTAIL.n558 VTAIL.n557 585
R24 VTAIL.n599 VTAIL.n598 585
R25 VTAIL.n601 VTAIL.n600 585
R26 VTAIL.n554 VTAIL.n553 585
R27 VTAIL.n607 VTAIL.n606 585
R28 VTAIL.n609 VTAIL.n608 585
R29 VTAIL.n550 VTAIL.n549 585
R30 VTAIL.n616 VTAIL.n615 585
R31 VTAIL.n617 VTAIL.n548 585
R32 VTAIL.n619 VTAIL.n618 585
R33 VTAIL.n24 VTAIL.n23 585
R34 VTAIL.n29 VTAIL.n28 585
R35 VTAIL.n31 VTAIL.n30 585
R36 VTAIL.n20 VTAIL.n19 585
R37 VTAIL.n37 VTAIL.n36 585
R38 VTAIL.n39 VTAIL.n38 585
R39 VTAIL.n16 VTAIL.n15 585
R40 VTAIL.n45 VTAIL.n44 585
R41 VTAIL.n47 VTAIL.n46 585
R42 VTAIL.n12 VTAIL.n11 585
R43 VTAIL.n53 VTAIL.n52 585
R44 VTAIL.n55 VTAIL.n54 585
R45 VTAIL.n8 VTAIL.n7 585
R46 VTAIL.n61 VTAIL.n60 585
R47 VTAIL.n63 VTAIL.n62 585
R48 VTAIL.n4 VTAIL.n3 585
R49 VTAIL.n70 VTAIL.n69 585
R50 VTAIL.n71 VTAIL.n2 585
R51 VTAIL.n73 VTAIL.n72 585
R52 VTAIL.n102 VTAIL.n101 585
R53 VTAIL.n107 VTAIL.n106 585
R54 VTAIL.n109 VTAIL.n108 585
R55 VTAIL.n98 VTAIL.n97 585
R56 VTAIL.n115 VTAIL.n114 585
R57 VTAIL.n117 VTAIL.n116 585
R58 VTAIL.n94 VTAIL.n93 585
R59 VTAIL.n123 VTAIL.n122 585
R60 VTAIL.n125 VTAIL.n124 585
R61 VTAIL.n90 VTAIL.n89 585
R62 VTAIL.n131 VTAIL.n130 585
R63 VTAIL.n133 VTAIL.n132 585
R64 VTAIL.n86 VTAIL.n85 585
R65 VTAIL.n139 VTAIL.n138 585
R66 VTAIL.n141 VTAIL.n140 585
R67 VTAIL.n82 VTAIL.n81 585
R68 VTAIL.n148 VTAIL.n147 585
R69 VTAIL.n149 VTAIL.n80 585
R70 VTAIL.n151 VTAIL.n150 585
R71 VTAIL.n180 VTAIL.n179 585
R72 VTAIL.n185 VTAIL.n184 585
R73 VTAIL.n187 VTAIL.n186 585
R74 VTAIL.n176 VTAIL.n175 585
R75 VTAIL.n193 VTAIL.n192 585
R76 VTAIL.n195 VTAIL.n194 585
R77 VTAIL.n172 VTAIL.n171 585
R78 VTAIL.n201 VTAIL.n200 585
R79 VTAIL.n203 VTAIL.n202 585
R80 VTAIL.n168 VTAIL.n167 585
R81 VTAIL.n209 VTAIL.n208 585
R82 VTAIL.n211 VTAIL.n210 585
R83 VTAIL.n164 VTAIL.n163 585
R84 VTAIL.n217 VTAIL.n216 585
R85 VTAIL.n219 VTAIL.n218 585
R86 VTAIL.n160 VTAIL.n159 585
R87 VTAIL.n226 VTAIL.n225 585
R88 VTAIL.n227 VTAIL.n158 585
R89 VTAIL.n229 VTAIL.n228 585
R90 VTAIL.n541 VTAIL.n540 585
R91 VTAIL.n539 VTAIL.n470 585
R92 VTAIL.n538 VTAIL.n537 585
R93 VTAIL.n473 VTAIL.n471 585
R94 VTAIL.n532 VTAIL.n531 585
R95 VTAIL.n530 VTAIL.n529 585
R96 VTAIL.n477 VTAIL.n476 585
R97 VTAIL.n524 VTAIL.n523 585
R98 VTAIL.n522 VTAIL.n521 585
R99 VTAIL.n481 VTAIL.n480 585
R100 VTAIL.n516 VTAIL.n515 585
R101 VTAIL.n514 VTAIL.n513 585
R102 VTAIL.n485 VTAIL.n484 585
R103 VTAIL.n508 VTAIL.n507 585
R104 VTAIL.n506 VTAIL.n505 585
R105 VTAIL.n489 VTAIL.n488 585
R106 VTAIL.n500 VTAIL.n499 585
R107 VTAIL.n498 VTAIL.n497 585
R108 VTAIL.n493 VTAIL.n492 585
R109 VTAIL.n463 VTAIL.n462 585
R110 VTAIL.n461 VTAIL.n392 585
R111 VTAIL.n460 VTAIL.n459 585
R112 VTAIL.n395 VTAIL.n393 585
R113 VTAIL.n454 VTAIL.n453 585
R114 VTAIL.n452 VTAIL.n451 585
R115 VTAIL.n399 VTAIL.n398 585
R116 VTAIL.n446 VTAIL.n445 585
R117 VTAIL.n444 VTAIL.n443 585
R118 VTAIL.n403 VTAIL.n402 585
R119 VTAIL.n438 VTAIL.n437 585
R120 VTAIL.n436 VTAIL.n435 585
R121 VTAIL.n407 VTAIL.n406 585
R122 VTAIL.n430 VTAIL.n429 585
R123 VTAIL.n428 VTAIL.n427 585
R124 VTAIL.n411 VTAIL.n410 585
R125 VTAIL.n422 VTAIL.n421 585
R126 VTAIL.n420 VTAIL.n419 585
R127 VTAIL.n415 VTAIL.n414 585
R128 VTAIL.n385 VTAIL.n384 585
R129 VTAIL.n383 VTAIL.n314 585
R130 VTAIL.n382 VTAIL.n381 585
R131 VTAIL.n317 VTAIL.n315 585
R132 VTAIL.n376 VTAIL.n375 585
R133 VTAIL.n374 VTAIL.n373 585
R134 VTAIL.n321 VTAIL.n320 585
R135 VTAIL.n368 VTAIL.n367 585
R136 VTAIL.n366 VTAIL.n365 585
R137 VTAIL.n325 VTAIL.n324 585
R138 VTAIL.n360 VTAIL.n359 585
R139 VTAIL.n358 VTAIL.n357 585
R140 VTAIL.n329 VTAIL.n328 585
R141 VTAIL.n352 VTAIL.n351 585
R142 VTAIL.n350 VTAIL.n349 585
R143 VTAIL.n333 VTAIL.n332 585
R144 VTAIL.n344 VTAIL.n343 585
R145 VTAIL.n342 VTAIL.n341 585
R146 VTAIL.n337 VTAIL.n336 585
R147 VTAIL.n307 VTAIL.n306 585
R148 VTAIL.n305 VTAIL.n236 585
R149 VTAIL.n304 VTAIL.n303 585
R150 VTAIL.n239 VTAIL.n237 585
R151 VTAIL.n298 VTAIL.n297 585
R152 VTAIL.n296 VTAIL.n295 585
R153 VTAIL.n243 VTAIL.n242 585
R154 VTAIL.n290 VTAIL.n289 585
R155 VTAIL.n288 VTAIL.n287 585
R156 VTAIL.n247 VTAIL.n246 585
R157 VTAIL.n282 VTAIL.n281 585
R158 VTAIL.n280 VTAIL.n279 585
R159 VTAIL.n251 VTAIL.n250 585
R160 VTAIL.n274 VTAIL.n273 585
R161 VTAIL.n272 VTAIL.n271 585
R162 VTAIL.n255 VTAIL.n254 585
R163 VTAIL.n266 VTAIL.n265 585
R164 VTAIL.n264 VTAIL.n263 585
R165 VTAIL.n259 VTAIL.n258 585
R166 VTAIL.n571 VTAIL.t3 327.466
R167 VTAIL.n25 VTAIL.t2 327.466
R168 VTAIL.n103 VTAIL.t1 327.466
R169 VTAIL.n181 VTAIL.t7 327.466
R170 VTAIL.n494 VTAIL.t0 327.466
R171 VTAIL.n416 VTAIL.t6 327.466
R172 VTAIL.n338 VTAIL.t4 327.466
R173 VTAIL.n260 VTAIL.t5 327.466
R174 VTAIL.n575 VTAIL.n569 171.744
R175 VTAIL.n576 VTAIL.n575 171.744
R176 VTAIL.n576 VTAIL.n565 171.744
R177 VTAIL.n583 VTAIL.n565 171.744
R178 VTAIL.n584 VTAIL.n583 171.744
R179 VTAIL.n584 VTAIL.n561 171.744
R180 VTAIL.n591 VTAIL.n561 171.744
R181 VTAIL.n592 VTAIL.n591 171.744
R182 VTAIL.n592 VTAIL.n557 171.744
R183 VTAIL.n599 VTAIL.n557 171.744
R184 VTAIL.n600 VTAIL.n599 171.744
R185 VTAIL.n600 VTAIL.n553 171.744
R186 VTAIL.n607 VTAIL.n553 171.744
R187 VTAIL.n608 VTAIL.n607 171.744
R188 VTAIL.n608 VTAIL.n549 171.744
R189 VTAIL.n616 VTAIL.n549 171.744
R190 VTAIL.n617 VTAIL.n616 171.744
R191 VTAIL.n618 VTAIL.n617 171.744
R192 VTAIL.n29 VTAIL.n23 171.744
R193 VTAIL.n30 VTAIL.n29 171.744
R194 VTAIL.n30 VTAIL.n19 171.744
R195 VTAIL.n37 VTAIL.n19 171.744
R196 VTAIL.n38 VTAIL.n37 171.744
R197 VTAIL.n38 VTAIL.n15 171.744
R198 VTAIL.n45 VTAIL.n15 171.744
R199 VTAIL.n46 VTAIL.n45 171.744
R200 VTAIL.n46 VTAIL.n11 171.744
R201 VTAIL.n53 VTAIL.n11 171.744
R202 VTAIL.n54 VTAIL.n53 171.744
R203 VTAIL.n54 VTAIL.n7 171.744
R204 VTAIL.n61 VTAIL.n7 171.744
R205 VTAIL.n62 VTAIL.n61 171.744
R206 VTAIL.n62 VTAIL.n3 171.744
R207 VTAIL.n70 VTAIL.n3 171.744
R208 VTAIL.n71 VTAIL.n70 171.744
R209 VTAIL.n72 VTAIL.n71 171.744
R210 VTAIL.n107 VTAIL.n101 171.744
R211 VTAIL.n108 VTAIL.n107 171.744
R212 VTAIL.n108 VTAIL.n97 171.744
R213 VTAIL.n115 VTAIL.n97 171.744
R214 VTAIL.n116 VTAIL.n115 171.744
R215 VTAIL.n116 VTAIL.n93 171.744
R216 VTAIL.n123 VTAIL.n93 171.744
R217 VTAIL.n124 VTAIL.n123 171.744
R218 VTAIL.n124 VTAIL.n89 171.744
R219 VTAIL.n131 VTAIL.n89 171.744
R220 VTAIL.n132 VTAIL.n131 171.744
R221 VTAIL.n132 VTAIL.n85 171.744
R222 VTAIL.n139 VTAIL.n85 171.744
R223 VTAIL.n140 VTAIL.n139 171.744
R224 VTAIL.n140 VTAIL.n81 171.744
R225 VTAIL.n148 VTAIL.n81 171.744
R226 VTAIL.n149 VTAIL.n148 171.744
R227 VTAIL.n150 VTAIL.n149 171.744
R228 VTAIL.n185 VTAIL.n179 171.744
R229 VTAIL.n186 VTAIL.n185 171.744
R230 VTAIL.n186 VTAIL.n175 171.744
R231 VTAIL.n193 VTAIL.n175 171.744
R232 VTAIL.n194 VTAIL.n193 171.744
R233 VTAIL.n194 VTAIL.n171 171.744
R234 VTAIL.n201 VTAIL.n171 171.744
R235 VTAIL.n202 VTAIL.n201 171.744
R236 VTAIL.n202 VTAIL.n167 171.744
R237 VTAIL.n209 VTAIL.n167 171.744
R238 VTAIL.n210 VTAIL.n209 171.744
R239 VTAIL.n210 VTAIL.n163 171.744
R240 VTAIL.n217 VTAIL.n163 171.744
R241 VTAIL.n218 VTAIL.n217 171.744
R242 VTAIL.n218 VTAIL.n159 171.744
R243 VTAIL.n226 VTAIL.n159 171.744
R244 VTAIL.n227 VTAIL.n226 171.744
R245 VTAIL.n228 VTAIL.n227 171.744
R246 VTAIL.n540 VTAIL.n539 171.744
R247 VTAIL.n539 VTAIL.n538 171.744
R248 VTAIL.n538 VTAIL.n471 171.744
R249 VTAIL.n531 VTAIL.n471 171.744
R250 VTAIL.n531 VTAIL.n530 171.744
R251 VTAIL.n530 VTAIL.n476 171.744
R252 VTAIL.n523 VTAIL.n476 171.744
R253 VTAIL.n523 VTAIL.n522 171.744
R254 VTAIL.n522 VTAIL.n480 171.744
R255 VTAIL.n515 VTAIL.n480 171.744
R256 VTAIL.n515 VTAIL.n514 171.744
R257 VTAIL.n514 VTAIL.n484 171.744
R258 VTAIL.n507 VTAIL.n484 171.744
R259 VTAIL.n507 VTAIL.n506 171.744
R260 VTAIL.n506 VTAIL.n488 171.744
R261 VTAIL.n499 VTAIL.n488 171.744
R262 VTAIL.n499 VTAIL.n498 171.744
R263 VTAIL.n498 VTAIL.n492 171.744
R264 VTAIL.n462 VTAIL.n461 171.744
R265 VTAIL.n461 VTAIL.n460 171.744
R266 VTAIL.n460 VTAIL.n393 171.744
R267 VTAIL.n453 VTAIL.n393 171.744
R268 VTAIL.n453 VTAIL.n452 171.744
R269 VTAIL.n452 VTAIL.n398 171.744
R270 VTAIL.n445 VTAIL.n398 171.744
R271 VTAIL.n445 VTAIL.n444 171.744
R272 VTAIL.n444 VTAIL.n402 171.744
R273 VTAIL.n437 VTAIL.n402 171.744
R274 VTAIL.n437 VTAIL.n436 171.744
R275 VTAIL.n436 VTAIL.n406 171.744
R276 VTAIL.n429 VTAIL.n406 171.744
R277 VTAIL.n429 VTAIL.n428 171.744
R278 VTAIL.n428 VTAIL.n410 171.744
R279 VTAIL.n421 VTAIL.n410 171.744
R280 VTAIL.n421 VTAIL.n420 171.744
R281 VTAIL.n420 VTAIL.n414 171.744
R282 VTAIL.n384 VTAIL.n383 171.744
R283 VTAIL.n383 VTAIL.n382 171.744
R284 VTAIL.n382 VTAIL.n315 171.744
R285 VTAIL.n375 VTAIL.n315 171.744
R286 VTAIL.n375 VTAIL.n374 171.744
R287 VTAIL.n374 VTAIL.n320 171.744
R288 VTAIL.n367 VTAIL.n320 171.744
R289 VTAIL.n367 VTAIL.n366 171.744
R290 VTAIL.n366 VTAIL.n324 171.744
R291 VTAIL.n359 VTAIL.n324 171.744
R292 VTAIL.n359 VTAIL.n358 171.744
R293 VTAIL.n358 VTAIL.n328 171.744
R294 VTAIL.n351 VTAIL.n328 171.744
R295 VTAIL.n351 VTAIL.n350 171.744
R296 VTAIL.n350 VTAIL.n332 171.744
R297 VTAIL.n343 VTAIL.n332 171.744
R298 VTAIL.n343 VTAIL.n342 171.744
R299 VTAIL.n342 VTAIL.n336 171.744
R300 VTAIL.n306 VTAIL.n305 171.744
R301 VTAIL.n305 VTAIL.n304 171.744
R302 VTAIL.n304 VTAIL.n237 171.744
R303 VTAIL.n297 VTAIL.n237 171.744
R304 VTAIL.n297 VTAIL.n296 171.744
R305 VTAIL.n296 VTAIL.n242 171.744
R306 VTAIL.n289 VTAIL.n242 171.744
R307 VTAIL.n289 VTAIL.n288 171.744
R308 VTAIL.n288 VTAIL.n246 171.744
R309 VTAIL.n281 VTAIL.n246 171.744
R310 VTAIL.n281 VTAIL.n280 171.744
R311 VTAIL.n280 VTAIL.n250 171.744
R312 VTAIL.n273 VTAIL.n250 171.744
R313 VTAIL.n273 VTAIL.n272 171.744
R314 VTAIL.n272 VTAIL.n254 171.744
R315 VTAIL.n265 VTAIL.n254 171.744
R316 VTAIL.n265 VTAIL.n264 171.744
R317 VTAIL.n264 VTAIL.n258 171.744
R318 VTAIL.t3 VTAIL.n569 85.8723
R319 VTAIL.t2 VTAIL.n23 85.8723
R320 VTAIL.t1 VTAIL.n101 85.8723
R321 VTAIL.t7 VTAIL.n179 85.8723
R322 VTAIL.t0 VTAIL.n492 85.8723
R323 VTAIL.t6 VTAIL.n414 85.8723
R324 VTAIL.t4 VTAIL.n336 85.8723
R325 VTAIL.t5 VTAIL.n258 85.8723
R326 VTAIL.n623 VTAIL.n622 33.5429
R327 VTAIL.n77 VTAIL.n76 33.5429
R328 VTAIL.n155 VTAIL.n154 33.5429
R329 VTAIL.n233 VTAIL.n232 33.5429
R330 VTAIL.n545 VTAIL.n544 33.5429
R331 VTAIL.n467 VTAIL.n466 33.5429
R332 VTAIL.n389 VTAIL.n388 33.5429
R333 VTAIL.n311 VTAIL.n310 33.5429
R334 VTAIL.n623 VTAIL.n545 26.0134
R335 VTAIL.n311 VTAIL.n233 26.0134
R336 VTAIL.n571 VTAIL.n570 16.3895
R337 VTAIL.n25 VTAIL.n24 16.3895
R338 VTAIL.n103 VTAIL.n102 16.3895
R339 VTAIL.n181 VTAIL.n180 16.3895
R340 VTAIL.n494 VTAIL.n493 16.3895
R341 VTAIL.n416 VTAIL.n415 16.3895
R342 VTAIL.n338 VTAIL.n337 16.3895
R343 VTAIL.n260 VTAIL.n259 16.3895
R344 VTAIL.n619 VTAIL.n548 13.1884
R345 VTAIL.n73 VTAIL.n2 13.1884
R346 VTAIL.n151 VTAIL.n80 13.1884
R347 VTAIL.n229 VTAIL.n158 13.1884
R348 VTAIL.n541 VTAIL.n470 13.1884
R349 VTAIL.n463 VTAIL.n392 13.1884
R350 VTAIL.n385 VTAIL.n314 13.1884
R351 VTAIL.n307 VTAIL.n236 13.1884
R352 VTAIL.n574 VTAIL.n573 12.8005
R353 VTAIL.n615 VTAIL.n614 12.8005
R354 VTAIL.n620 VTAIL.n546 12.8005
R355 VTAIL.n28 VTAIL.n27 12.8005
R356 VTAIL.n69 VTAIL.n68 12.8005
R357 VTAIL.n74 VTAIL.n0 12.8005
R358 VTAIL.n106 VTAIL.n105 12.8005
R359 VTAIL.n147 VTAIL.n146 12.8005
R360 VTAIL.n152 VTAIL.n78 12.8005
R361 VTAIL.n184 VTAIL.n183 12.8005
R362 VTAIL.n225 VTAIL.n224 12.8005
R363 VTAIL.n230 VTAIL.n156 12.8005
R364 VTAIL.n542 VTAIL.n468 12.8005
R365 VTAIL.n537 VTAIL.n472 12.8005
R366 VTAIL.n497 VTAIL.n496 12.8005
R367 VTAIL.n464 VTAIL.n390 12.8005
R368 VTAIL.n459 VTAIL.n394 12.8005
R369 VTAIL.n419 VTAIL.n418 12.8005
R370 VTAIL.n386 VTAIL.n312 12.8005
R371 VTAIL.n381 VTAIL.n316 12.8005
R372 VTAIL.n341 VTAIL.n340 12.8005
R373 VTAIL.n308 VTAIL.n234 12.8005
R374 VTAIL.n303 VTAIL.n238 12.8005
R375 VTAIL.n263 VTAIL.n262 12.8005
R376 VTAIL.n577 VTAIL.n568 12.0247
R377 VTAIL.n613 VTAIL.n550 12.0247
R378 VTAIL.n31 VTAIL.n22 12.0247
R379 VTAIL.n67 VTAIL.n4 12.0247
R380 VTAIL.n109 VTAIL.n100 12.0247
R381 VTAIL.n145 VTAIL.n82 12.0247
R382 VTAIL.n187 VTAIL.n178 12.0247
R383 VTAIL.n223 VTAIL.n160 12.0247
R384 VTAIL.n536 VTAIL.n473 12.0247
R385 VTAIL.n500 VTAIL.n491 12.0247
R386 VTAIL.n458 VTAIL.n395 12.0247
R387 VTAIL.n422 VTAIL.n413 12.0247
R388 VTAIL.n380 VTAIL.n317 12.0247
R389 VTAIL.n344 VTAIL.n335 12.0247
R390 VTAIL.n302 VTAIL.n239 12.0247
R391 VTAIL.n266 VTAIL.n257 12.0247
R392 VTAIL.n578 VTAIL.n566 11.249
R393 VTAIL.n610 VTAIL.n609 11.249
R394 VTAIL.n32 VTAIL.n20 11.249
R395 VTAIL.n64 VTAIL.n63 11.249
R396 VTAIL.n110 VTAIL.n98 11.249
R397 VTAIL.n142 VTAIL.n141 11.249
R398 VTAIL.n188 VTAIL.n176 11.249
R399 VTAIL.n220 VTAIL.n219 11.249
R400 VTAIL.n533 VTAIL.n532 11.249
R401 VTAIL.n501 VTAIL.n489 11.249
R402 VTAIL.n455 VTAIL.n454 11.249
R403 VTAIL.n423 VTAIL.n411 11.249
R404 VTAIL.n377 VTAIL.n376 11.249
R405 VTAIL.n345 VTAIL.n333 11.249
R406 VTAIL.n299 VTAIL.n298 11.249
R407 VTAIL.n267 VTAIL.n255 11.249
R408 VTAIL.n582 VTAIL.n581 10.4732
R409 VTAIL.n606 VTAIL.n552 10.4732
R410 VTAIL.n36 VTAIL.n35 10.4732
R411 VTAIL.n60 VTAIL.n6 10.4732
R412 VTAIL.n114 VTAIL.n113 10.4732
R413 VTAIL.n138 VTAIL.n84 10.4732
R414 VTAIL.n192 VTAIL.n191 10.4732
R415 VTAIL.n216 VTAIL.n162 10.4732
R416 VTAIL.n529 VTAIL.n475 10.4732
R417 VTAIL.n505 VTAIL.n504 10.4732
R418 VTAIL.n451 VTAIL.n397 10.4732
R419 VTAIL.n427 VTAIL.n426 10.4732
R420 VTAIL.n373 VTAIL.n319 10.4732
R421 VTAIL.n349 VTAIL.n348 10.4732
R422 VTAIL.n295 VTAIL.n241 10.4732
R423 VTAIL.n271 VTAIL.n270 10.4732
R424 VTAIL.n585 VTAIL.n564 9.69747
R425 VTAIL.n605 VTAIL.n554 9.69747
R426 VTAIL.n39 VTAIL.n18 9.69747
R427 VTAIL.n59 VTAIL.n8 9.69747
R428 VTAIL.n117 VTAIL.n96 9.69747
R429 VTAIL.n137 VTAIL.n86 9.69747
R430 VTAIL.n195 VTAIL.n174 9.69747
R431 VTAIL.n215 VTAIL.n164 9.69747
R432 VTAIL.n528 VTAIL.n477 9.69747
R433 VTAIL.n508 VTAIL.n487 9.69747
R434 VTAIL.n450 VTAIL.n399 9.69747
R435 VTAIL.n430 VTAIL.n409 9.69747
R436 VTAIL.n372 VTAIL.n321 9.69747
R437 VTAIL.n352 VTAIL.n331 9.69747
R438 VTAIL.n294 VTAIL.n243 9.69747
R439 VTAIL.n274 VTAIL.n253 9.69747
R440 VTAIL.n622 VTAIL.n621 9.45567
R441 VTAIL.n76 VTAIL.n75 9.45567
R442 VTAIL.n154 VTAIL.n153 9.45567
R443 VTAIL.n232 VTAIL.n231 9.45567
R444 VTAIL.n544 VTAIL.n543 9.45567
R445 VTAIL.n466 VTAIL.n465 9.45567
R446 VTAIL.n388 VTAIL.n387 9.45567
R447 VTAIL.n310 VTAIL.n309 9.45567
R448 VTAIL.n621 VTAIL.n620 9.3005
R449 VTAIL.n560 VTAIL.n559 9.3005
R450 VTAIL.n589 VTAIL.n588 9.3005
R451 VTAIL.n587 VTAIL.n586 9.3005
R452 VTAIL.n564 VTAIL.n563 9.3005
R453 VTAIL.n581 VTAIL.n580 9.3005
R454 VTAIL.n579 VTAIL.n578 9.3005
R455 VTAIL.n568 VTAIL.n567 9.3005
R456 VTAIL.n573 VTAIL.n572 9.3005
R457 VTAIL.n595 VTAIL.n594 9.3005
R458 VTAIL.n597 VTAIL.n596 9.3005
R459 VTAIL.n556 VTAIL.n555 9.3005
R460 VTAIL.n603 VTAIL.n602 9.3005
R461 VTAIL.n605 VTAIL.n604 9.3005
R462 VTAIL.n552 VTAIL.n551 9.3005
R463 VTAIL.n611 VTAIL.n610 9.3005
R464 VTAIL.n613 VTAIL.n612 9.3005
R465 VTAIL.n614 VTAIL.n547 9.3005
R466 VTAIL.n75 VTAIL.n74 9.3005
R467 VTAIL.n14 VTAIL.n13 9.3005
R468 VTAIL.n43 VTAIL.n42 9.3005
R469 VTAIL.n41 VTAIL.n40 9.3005
R470 VTAIL.n18 VTAIL.n17 9.3005
R471 VTAIL.n35 VTAIL.n34 9.3005
R472 VTAIL.n33 VTAIL.n32 9.3005
R473 VTAIL.n22 VTAIL.n21 9.3005
R474 VTAIL.n27 VTAIL.n26 9.3005
R475 VTAIL.n49 VTAIL.n48 9.3005
R476 VTAIL.n51 VTAIL.n50 9.3005
R477 VTAIL.n10 VTAIL.n9 9.3005
R478 VTAIL.n57 VTAIL.n56 9.3005
R479 VTAIL.n59 VTAIL.n58 9.3005
R480 VTAIL.n6 VTAIL.n5 9.3005
R481 VTAIL.n65 VTAIL.n64 9.3005
R482 VTAIL.n67 VTAIL.n66 9.3005
R483 VTAIL.n68 VTAIL.n1 9.3005
R484 VTAIL.n153 VTAIL.n152 9.3005
R485 VTAIL.n92 VTAIL.n91 9.3005
R486 VTAIL.n121 VTAIL.n120 9.3005
R487 VTAIL.n119 VTAIL.n118 9.3005
R488 VTAIL.n96 VTAIL.n95 9.3005
R489 VTAIL.n113 VTAIL.n112 9.3005
R490 VTAIL.n111 VTAIL.n110 9.3005
R491 VTAIL.n100 VTAIL.n99 9.3005
R492 VTAIL.n105 VTAIL.n104 9.3005
R493 VTAIL.n127 VTAIL.n126 9.3005
R494 VTAIL.n129 VTAIL.n128 9.3005
R495 VTAIL.n88 VTAIL.n87 9.3005
R496 VTAIL.n135 VTAIL.n134 9.3005
R497 VTAIL.n137 VTAIL.n136 9.3005
R498 VTAIL.n84 VTAIL.n83 9.3005
R499 VTAIL.n143 VTAIL.n142 9.3005
R500 VTAIL.n145 VTAIL.n144 9.3005
R501 VTAIL.n146 VTAIL.n79 9.3005
R502 VTAIL.n231 VTAIL.n230 9.3005
R503 VTAIL.n170 VTAIL.n169 9.3005
R504 VTAIL.n199 VTAIL.n198 9.3005
R505 VTAIL.n197 VTAIL.n196 9.3005
R506 VTAIL.n174 VTAIL.n173 9.3005
R507 VTAIL.n191 VTAIL.n190 9.3005
R508 VTAIL.n189 VTAIL.n188 9.3005
R509 VTAIL.n178 VTAIL.n177 9.3005
R510 VTAIL.n183 VTAIL.n182 9.3005
R511 VTAIL.n205 VTAIL.n204 9.3005
R512 VTAIL.n207 VTAIL.n206 9.3005
R513 VTAIL.n166 VTAIL.n165 9.3005
R514 VTAIL.n213 VTAIL.n212 9.3005
R515 VTAIL.n215 VTAIL.n214 9.3005
R516 VTAIL.n162 VTAIL.n161 9.3005
R517 VTAIL.n221 VTAIL.n220 9.3005
R518 VTAIL.n223 VTAIL.n222 9.3005
R519 VTAIL.n224 VTAIL.n157 9.3005
R520 VTAIL.n520 VTAIL.n519 9.3005
R521 VTAIL.n479 VTAIL.n478 9.3005
R522 VTAIL.n526 VTAIL.n525 9.3005
R523 VTAIL.n528 VTAIL.n527 9.3005
R524 VTAIL.n475 VTAIL.n474 9.3005
R525 VTAIL.n534 VTAIL.n533 9.3005
R526 VTAIL.n536 VTAIL.n535 9.3005
R527 VTAIL.n472 VTAIL.n469 9.3005
R528 VTAIL.n543 VTAIL.n542 9.3005
R529 VTAIL.n518 VTAIL.n517 9.3005
R530 VTAIL.n483 VTAIL.n482 9.3005
R531 VTAIL.n512 VTAIL.n511 9.3005
R532 VTAIL.n510 VTAIL.n509 9.3005
R533 VTAIL.n487 VTAIL.n486 9.3005
R534 VTAIL.n504 VTAIL.n503 9.3005
R535 VTAIL.n502 VTAIL.n501 9.3005
R536 VTAIL.n491 VTAIL.n490 9.3005
R537 VTAIL.n496 VTAIL.n495 9.3005
R538 VTAIL.n442 VTAIL.n441 9.3005
R539 VTAIL.n401 VTAIL.n400 9.3005
R540 VTAIL.n448 VTAIL.n447 9.3005
R541 VTAIL.n450 VTAIL.n449 9.3005
R542 VTAIL.n397 VTAIL.n396 9.3005
R543 VTAIL.n456 VTAIL.n455 9.3005
R544 VTAIL.n458 VTAIL.n457 9.3005
R545 VTAIL.n394 VTAIL.n391 9.3005
R546 VTAIL.n465 VTAIL.n464 9.3005
R547 VTAIL.n440 VTAIL.n439 9.3005
R548 VTAIL.n405 VTAIL.n404 9.3005
R549 VTAIL.n434 VTAIL.n433 9.3005
R550 VTAIL.n432 VTAIL.n431 9.3005
R551 VTAIL.n409 VTAIL.n408 9.3005
R552 VTAIL.n426 VTAIL.n425 9.3005
R553 VTAIL.n424 VTAIL.n423 9.3005
R554 VTAIL.n413 VTAIL.n412 9.3005
R555 VTAIL.n418 VTAIL.n417 9.3005
R556 VTAIL.n364 VTAIL.n363 9.3005
R557 VTAIL.n323 VTAIL.n322 9.3005
R558 VTAIL.n370 VTAIL.n369 9.3005
R559 VTAIL.n372 VTAIL.n371 9.3005
R560 VTAIL.n319 VTAIL.n318 9.3005
R561 VTAIL.n378 VTAIL.n377 9.3005
R562 VTAIL.n380 VTAIL.n379 9.3005
R563 VTAIL.n316 VTAIL.n313 9.3005
R564 VTAIL.n387 VTAIL.n386 9.3005
R565 VTAIL.n362 VTAIL.n361 9.3005
R566 VTAIL.n327 VTAIL.n326 9.3005
R567 VTAIL.n356 VTAIL.n355 9.3005
R568 VTAIL.n354 VTAIL.n353 9.3005
R569 VTAIL.n331 VTAIL.n330 9.3005
R570 VTAIL.n348 VTAIL.n347 9.3005
R571 VTAIL.n346 VTAIL.n345 9.3005
R572 VTAIL.n335 VTAIL.n334 9.3005
R573 VTAIL.n340 VTAIL.n339 9.3005
R574 VTAIL.n286 VTAIL.n285 9.3005
R575 VTAIL.n245 VTAIL.n244 9.3005
R576 VTAIL.n292 VTAIL.n291 9.3005
R577 VTAIL.n294 VTAIL.n293 9.3005
R578 VTAIL.n241 VTAIL.n240 9.3005
R579 VTAIL.n300 VTAIL.n299 9.3005
R580 VTAIL.n302 VTAIL.n301 9.3005
R581 VTAIL.n238 VTAIL.n235 9.3005
R582 VTAIL.n309 VTAIL.n308 9.3005
R583 VTAIL.n284 VTAIL.n283 9.3005
R584 VTAIL.n249 VTAIL.n248 9.3005
R585 VTAIL.n278 VTAIL.n277 9.3005
R586 VTAIL.n276 VTAIL.n275 9.3005
R587 VTAIL.n253 VTAIL.n252 9.3005
R588 VTAIL.n270 VTAIL.n269 9.3005
R589 VTAIL.n268 VTAIL.n267 9.3005
R590 VTAIL.n257 VTAIL.n256 9.3005
R591 VTAIL.n262 VTAIL.n261 9.3005
R592 VTAIL.n586 VTAIL.n562 8.92171
R593 VTAIL.n602 VTAIL.n601 8.92171
R594 VTAIL.n40 VTAIL.n16 8.92171
R595 VTAIL.n56 VTAIL.n55 8.92171
R596 VTAIL.n118 VTAIL.n94 8.92171
R597 VTAIL.n134 VTAIL.n133 8.92171
R598 VTAIL.n196 VTAIL.n172 8.92171
R599 VTAIL.n212 VTAIL.n211 8.92171
R600 VTAIL.n525 VTAIL.n524 8.92171
R601 VTAIL.n509 VTAIL.n485 8.92171
R602 VTAIL.n447 VTAIL.n446 8.92171
R603 VTAIL.n431 VTAIL.n407 8.92171
R604 VTAIL.n369 VTAIL.n368 8.92171
R605 VTAIL.n353 VTAIL.n329 8.92171
R606 VTAIL.n291 VTAIL.n290 8.92171
R607 VTAIL.n275 VTAIL.n251 8.92171
R608 VTAIL.n590 VTAIL.n589 8.14595
R609 VTAIL.n598 VTAIL.n556 8.14595
R610 VTAIL.n44 VTAIL.n43 8.14595
R611 VTAIL.n52 VTAIL.n10 8.14595
R612 VTAIL.n122 VTAIL.n121 8.14595
R613 VTAIL.n130 VTAIL.n88 8.14595
R614 VTAIL.n200 VTAIL.n199 8.14595
R615 VTAIL.n208 VTAIL.n166 8.14595
R616 VTAIL.n521 VTAIL.n479 8.14595
R617 VTAIL.n513 VTAIL.n512 8.14595
R618 VTAIL.n443 VTAIL.n401 8.14595
R619 VTAIL.n435 VTAIL.n434 8.14595
R620 VTAIL.n365 VTAIL.n323 8.14595
R621 VTAIL.n357 VTAIL.n356 8.14595
R622 VTAIL.n287 VTAIL.n245 8.14595
R623 VTAIL.n279 VTAIL.n278 8.14595
R624 VTAIL.n593 VTAIL.n560 7.3702
R625 VTAIL.n597 VTAIL.n558 7.3702
R626 VTAIL.n47 VTAIL.n14 7.3702
R627 VTAIL.n51 VTAIL.n12 7.3702
R628 VTAIL.n125 VTAIL.n92 7.3702
R629 VTAIL.n129 VTAIL.n90 7.3702
R630 VTAIL.n203 VTAIL.n170 7.3702
R631 VTAIL.n207 VTAIL.n168 7.3702
R632 VTAIL.n520 VTAIL.n481 7.3702
R633 VTAIL.n516 VTAIL.n483 7.3702
R634 VTAIL.n442 VTAIL.n403 7.3702
R635 VTAIL.n438 VTAIL.n405 7.3702
R636 VTAIL.n364 VTAIL.n325 7.3702
R637 VTAIL.n360 VTAIL.n327 7.3702
R638 VTAIL.n286 VTAIL.n247 7.3702
R639 VTAIL.n282 VTAIL.n249 7.3702
R640 VTAIL.n594 VTAIL.n593 6.59444
R641 VTAIL.n594 VTAIL.n558 6.59444
R642 VTAIL.n48 VTAIL.n47 6.59444
R643 VTAIL.n48 VTAIL.n12 6.59444
R644 VTAIL.n126 VTAIL.n125 6.59444
R645 VTAIL.n126 VTAIL.n90 6.59444
R646 VTAIL.n204 VTAIL.n203 6.59444
R647 VTAIL.n204 VTAIL.n168 6.59444
R648 VTAIL.n517 VTAIL.n481 6.59444
R649 VTAIL.n517 VTAIL.n516 6.59444
R650 VTAIL.n439 VTAIL.n403 6.59444
R651 VTAIL.n439 VTAIL.n438 6.59444
R652 VTAIL.n361 VTAIL.n325 6.59444
R653 VTAIL.n361 VTAIL.n360 6.59444
R654 VTAIL.n283 VTAIL.n247 6.59444
R655 VTAIL.n283 VTAIL.n282 6.59444
R656 VTAIL.n590 VTAIL.n560 5.81868
R657 VTAIL.n598 VTAIL.n597 5.81868
R658 VTAIL.n44 VTAIL.n14 5.81868
R659 VTAIL.n52 VTAIL.n51 5.81868
R660 VTAIL.n122 VTAIL.n92 5.81868
R661 VTAIL.n130 VTAIL.n129 5.81868
R662 VTAIL.n200 VTAIL.n170 5.81868
R663 VTAIL.n208 VTAIL.n207 5.81868
R664 VTAIL.n521 VTAIL.n520 5.81868
R665 VTAIL.n513 VTAIL.n483 5.81868
R666 VTAIL.n443 VTAIL.n442 5.81868
R667 VTAIL.n435 VTAIL.n405 5.81868
R668 VTAIL.n365 VTAIL.n364 5.81868
R669 VTAIL.n357 VTAIL.n327 5.81868
R670 VTAIL.n287 VTAIL.n286 5.81868
R671 VTAIL.n279 VTAIL.n249 5.81868
R672 VTAIL.n589 VTAIL.n562 5.04292
R673 VTAIL.n601 VTAIL.n556 5.04292
R674 VTAIL.n43 VTAIL.n16 5.04292
R675 VTAIL.n55 VTAIL.n10 5.04292
R676 VTAIL.n121 VTAIL.n94 5.04292
R677 VTAIL.n133 VTAIL.n88 5.04292
R678 VTAIL.n199 VTAIL.n172 5.04292
R679 VTAIL.n211 VTAIL.n166 5.04292
R680 VTAIL.n524 VTAIL.n479 5.04292
R681 VTAIL.n512 VTAIL.n485 5.04292
R682 VTAIL.n446 VTAIL.n401 5.04292
R683 VTAIL.n434 VTAIL.n407 5.04292
R684 VTAIL.n368 VTAIL.n323 5.04292
R685 VTAIL.n356 VTAIL.n329 5.04292
R686 VTAIL.n290 VTAIL.n245 5.04292
R687 VTAIL.n278 VTAIL.n251 5.04292
R688 VTAIL.n586 VTAIL.n585 4.26717
R689 VTAIL.n602 VTAIL.n554 4.26717
R690 VTAIL.n40 VTAIL.n39 4.26717
R691 VTAIL.n56 VTAIL.n8 4.26717
R692 VTAIL.n118 VTAIL.n117 4.26717
R693 VTAIL.n134 VTAIL.n86 4.26717
R694 VTAIL.n196 VTAIL.n195 4.26717
R695 VTAIL.n212 VTAIL.n164 4.26717
R696 VTAIL.n525 VTAIL.n477 4.26717
R697 VTAIL.n509 VTAIL.n508 4.26717
R698 VTAIL.n447 VTAIL.n399 4.26717
R699 VTAIL.n431 VTAIL.n430 4.26717
R700 VTAIL.n369 VTAIL.n321 4.26717
R701 VTAIL.n353 VTAIL.n352 4.26717
R702 VTAIL.n291 VTAIL.n243 4.26717
R703 VTAIL.n275 VTAIL.n274 4.26717
R704 VTAIL.n572 VTAIL.n571 3.70982
R705 VTAIL.n26 VTAIL.n25 3.70982
R706 VTAIL.n104 VTAIL.n103 3.70982
R707 VTAIL.n182 VTAIL.n181 3.70982
R708 VTAIL.n495 VTAIL.n494 3.70982
R709 VTAIL.n417 VTAIL.n416 3.70982
R710 VTAIL.n339 VTAIL.n338 3.70982
R711 VTAIL.n261 VTAIL.n260 3.70982
R712 VTAIL.n582 VTAIL.n564 3.49141
R713 VTAIL.n606 VTAIL.n605 3.49141
R714 VTAIL.n36 VTAIL.n18 3.49141
R715 VTAIL.n60 VTAIL.n59 3.49141
R716 VTAIL.n114 VTAIL.n96 3.49141
R717 VTAIL.n138 VTAIL.n137 3.49141
R718 VTAIL.n192 VTAIL.n174 3.49141
R719 VTAIL.n216 VTAIL.n215 3.49141
R720 VTAIL.n529 VTAIL.n528 3.49141
R721 VTAIL.n505 VTAIL.n487 3.49141
R722 VTAIL.n451 VTAIL.n450 3.49141
R723 VTAIL.n427 VTAIL.n409 3.49141
R724 VTAIL.n373 VTAIL.n372 3.49141
R725 VTAIL.n349 VTAIL.n331 3.49141
R726 VTAIL.n295 VTAIL.n294 3.49141
R727 VTAIL.n271 VTAIL.n253 3.49141
R728 VTAIL.n581 VTAIL.n566 2.71565
R729 VTAIL.n609 VTAIL.n552 2.71565
R730 VTAIL.n35 VTAIL.n20 2.71565
R731 VTAIL.n63 VTAIL.n6 2.71565
R732 VTAIL.n113 VTAIL.n98 2.71565
R733 VTAIL.n141 VTAIL.n84 2.71565
R734 VTAIL.n191 VTAIL.n176 2.71565
R735 VTAIL.n219 VTAIL.n162 2.71565
R736 VTAIL.n532 VTAIL.n475 2.71565
R737 VTAIL.n504 VTAIL.n489 2.71565
R738 VTAIL.n454 VTAIL.n397 2.71565
R739 VTAIL.n426 VTAIL.n411 2.71565
R740 VTAIL.n376 VTAIL.n319 2.71565
R741 VTAIL.n348 VTAIL.n333 2.71565
R742 VTAIL.n298 VTAIL.n241 2.71565
R743 VTAIL.n270 VTAIL.n255 2.71565
R744 VTAIL.n578 VTAIL.n577 1.93989
R745 VTAIL.n610 VTAIL.n550 1.93989
R746 VTAIL.n32 VTAIL.n31 1.93989
R747 VTAIL.n64 VTAIL.n4 1.93989
R748 VTAIL.n110 VTAIL.n109 1.93989
R749 VTAIL.n142 VTAIL.n82 1.93989
R750 VTAIL.n188 VTAIL.n187 1.93989
R751 VTAIL.n220 VTAIL.n160 1.93989
R752 VTAIL.n533 VTAIL.n473 1.93989
R753 VTAIL.n501 VTAIL.n500 1.93989
R754 VTAIL.n455 VTAIL.n395 1.93989
R755 VTAIL.n423 VTAIL.n422 1.93989
R756 VTAIL.n377 VTAIL.n317 1.93989
R757 VTAIL.n345 VTAIL.n344 1.93989
R758 VTAIL.n299 VTAIL.n239 1.93989
R759 VTAIL.n267 VTAIL.n266 1.93989
R760 VTAIL.n389 VTAIL.n311 1.58671
R761 VTAIL.n545 VTAIL.n467 1.58671
R762 VTAIL.n233 VTAIL.n155 1.58671
R763 VTAIL.n574 VTAIL.n568 1.16414
R764 VTAIL.n615 VTAIL.n613 1.16414
R765 VTAIL.n622 VTAIL.n546 1.16414
R766 VTAIL.n28 VTAIL.n22 1.16414
R767 VTAIL.n69 VTAIL.n67 1.16414
R768 VTAIL.n76 VTAIL.n0 1.16414
R769 VTAIL.n106 VTAIL.n100 1.16414
R770 VTAIL.n147 VTAIL.n145 1.16414
R771 VTAIL.n154 VTAIL.n78 1.16414
R772 VTAIL.n184 VTAIL.n178 1.16414
R773 VTAIL.n225 VTAIL.n223 1.16414
R774 VTAIL.n232 VTAIL.n156 1.16414
R775 VTAIL.n544 VTAIL.n468 1.16414
R776 VTAIL.n537 VTAIL.n536 1.16414
R777 VTAIL.n497 VTAIL.n491 1.16414
R778 VTAIL.n466 VTAIL.n390 1.16414
R779 VTAIL.n459 VTAIL.n458 1.16414
R780 VTAIL.n419 VTAIL.n413 1.16414
R781 VTAIL.n388 VTAIL.n312 1.16414
R782 VTAIL.n381 VTAIL.n380 1.16414
R783 VTAIL.n341 VTAIL.n335 1.16414
R784 VTAIL.n310 VTAIL.n234 1.16414
R785 VTAIL.n303 VTAIL.n302 1.16414
R786 VTAIL.n263 VTAIL.n257 1.16414
R787 VTAIL VTAIL.n77 0.851793
R788 VTAIL VTAIL.n623 0.735414
R789 VTAIL.n467 VTAIL.n389 0.470328
R790 VTAIL.n155 VTAIL.n77 0.470328
R791 VTAIL.n573 VTAIL.n570 0.388379
R792 VTAIL.n614 VTAIL.n548 0.388379
R793 VTAIL.n620 VTAIL.n619 0.388379
R794 VTAIL.n27 VTAIL.n24 0.388379
R795 VTAIL.n68 VTAIL.n2 0.388379
R796 VTAIL.n74 VTAIL.n73 0.388379
R797 VTAIL.n105 VTAIL.n102 0.388379
R798 VTAIL.n146 VTAIL.n80 0.388379
R799 VTAIL.n152 VTAIL.n151 0.388379
R800 VTAIL.n183 VTAIL.n180 0.388379
R801 VTAIL.n224 VTAIL.n158 0.388379
R802 VTAIL.n230 VTAIL.n229 0.388379
R803 VTAIL.n542 VTAIL.n541 0.388379
R804 VTAIL.n472 VTAIL.n470 0.388379
R805 VTAIL.n496 VTAIL.n493 0.388379
R806 VTAIL.n464 VTAIL.n463 0.388379
R807 VTAIL.n394 VTAIL.n392 0.388379
R808 VTAIL.n418 VTAIL.n415 0.388379
R809 VTAIL.n386 VTAIL.n385 0.388379
R810 VTAIL.n316 VTAIL.n314 0.388379
R811 VTAIL.n340 VTAIL.n337 0.388379
R812 VTAIL.n308 VTAIL.n307 0.388379
R813 VTAIL.n238 VTAIL.n236 0.388379
R814 VTAIL.n262 VTAIL.n259 0.388379
R815 VTAIL.n572 VTAIL.n567 0.155672
R816 VTAIL.n579 VTAIL.n567 0.155672
R817 VTAIL.n580 VTAIL.n579 0.155672
R818 VTAIL.n580 VTAIL.n563 0.155672
R819 VTAIL.n587 VTAIL.n563 0.155672
R820 VTAIL.n588 VTAIL.n587 0.155672
R821 VTAIL.n588 VTAIL.n559 0.155672
R822 VTAIL.n595 VTAIL.n559 0.155672
R823 VTAIL.n596 VTAIL.n595 0.155672
R824 VTAIL.n596 VTAIL.n555 0.155672
R825 VTAIL.n603 VTAIL.n555 0.155672
R826 VTAIL.n604 VTAIL.n603 0.155672
R827 VTAIL.n604 VTAIL.n551 0.155672
R828 VTAIL.n611 VTAIL.n551 0.155672
R829 VTAIL.n612 VTAIL.n611 0.155672
R830 VTAIL.n612 VTAIL.n547 0.155672
R831 VTAIL.n621 VTAIL.n547 0.155672
R832 VTAIL.n26 VTAIL.n21 0.155672
R833 VTAIL.n33 VTAIL.n21 0.155672
R834 VTAIL.n34 VTAIL.n33 0.155672
R835 VTAIL.n34 VTAIL.n17 0.155672
R836 VTAIL.n41 VTAIL.n17 0.155672
R837 VTAIL.n42 VTAIL.n41 0.155672
R838 VTAIL.n42 VTAIL.n13 0.155672
R839 VTAIL.n49 VTAIL.n13 0.155672
R840 VTAIL.n50 VTAIL.n49 0.155672
R841 VTAIL.n50 VTAIL.n9 0.155672
R842 VTAIL.n57 VTAIL.n9 0.155672
R843 VTAIL.n58 VTAIL.n57 0.155672
R844 VTAIL.n58 VTAIL.n5 0.155672
R845 VTAIL.n65 VTAIL.n5 0.155672
R846 VTAIL.n66 VTAIL.n65 0.155672
R847 VTAIL.n66 VTAIL.n1 0.155672
R848 VTAIL.n75 VTAIL.n1 0.155672
R849 VTAIL.n104 VTAIL.n99 0.155672
R850 VTAIL.n111 VTAIL.n99 0.155672
R851 VTAIL.n112 VTAIL.n111 0.155672
R852 VTAIL.n112 VTAIL.n95 0.155672
R853 VTAIL.n119 VTAIL.n95 0.155672
R854 VTAIL.n120 VTAIL.n119 0.155672
R855 VTAIL.n120 VTAIL.n91 0.155672
R856 VTAIL.n127 VTAIL.n91 0.155672
R857 VTAIL.n128 VTAIL.n127 0.155672
R858 VTAIL.n128 VTAIL.n87 0.155672
R859 VTAIL.n135 VTAIL.n87 0.155672
R860 VTAIL.n136 VTAIL.n135 0.155672
R861 VTAIL.n136 VTAIL.n83 0.155672
R862 VTAIL.n143 VTAIL.n83 0.155672
R863 VTAIL.n144 VTAIL.n143 0.155672
R864 VTAIL.n144 VTAIL.n79 0.155672
R865 VTAIL.n153 VTAIL.n79 0.155672
R866 VTAIL.n182 VTAIL.n177 0.155672
R867 VTAIL.n189 VTAIL.n177 0.155672
R868 VTAIL.n190 VTAIL.n189 0.155672
R869 VTAIL.n190 VTAIL.n173 0.155672
R870 VTAIL.n197 VTAIL.n173 0.155672
R871 VTAIL.n198 VTAIL.n197 0.155672
R872 VTAIL.n198 VTAIL.n169 0.155672
R873 VTAIL.n205 VTAIL.n169 0.155672
R874 VTAIL.n206 VTAIL.n205 0.155672
R875 VTAIL.n206 VTAIL.n165 0.155672
R876 VTAIL.n213 VTAIL.n165 0.155672
R877 VTAIL.n214 VTAIL.n213 0.155672
R878 VTAIL.n214 VTAIL.n161 0.155672
R879 VTAIL.n221 VTAIL.n161 0.155672
R880 VTAIL.n222 VTAIL.n221 0.155672
R881 VTAIL.n222 VTAIL.n157 0.155672
R882 VTAIL.n231 VTAIL.n157 0.155672
R883 VTAIL.n543 VTAIL.n469 0.155672
R884 VTAIL.n535 VTAIL.n469 0.155672
R885 VTAIL.n535 VTAIL.n534 0.155672
R886 VTAIL.n534 VTAIL.n474 0.155672
R887 VTAIL.n527 VTAIL.n474 0.155672
R888 VTAIL.n527 VTAIL.n526 0.155672
R889 VTAIL.n526 VTAIL.n478 0.155672
R890 VTAIL.n519 VTAIL.n478 0.155672
R891 VTAIL.n519 VTAIL.n518 0.155672
R892 VTAIL.n518 VTAIL.n482 0.155672
R893 VTAIL.n511 VTAIL.n482 0.155672
R894 VTAIL.n511 VTAIL.n510 0.155672
R895 VTAIL.n510 VTAIL.n486 0.155672
R896 VTAIL.n503 VTAIL.n486 0.155672
R897 VTAIL.n503 VTAIL.n502 0.155672
R898 VTAIL.n502 VTAIL.n490 0.155672
R899 VTAIL.n495 VTAIL.n490 0.155672
R900 VTAIL.n465 VTAIL.n391 0.155672
R901 VTAIL.n457 VTAIL.n391 0.155672
R902 VTAIL.n457 VTAIL.n456 0.155672
R903 VTAIL.n456 VTAIL.n396 0.155672
R904 VTAIL.n449 VTAIL.n396 0.155672
R905 VTAIL.n449 VTAIL.n448 0.155672
R906 VTAIL.n448 VTAIL.n400 0.155672
R907 VTAIL.n441 VTAIL.n400 0.155672
R908 VTAIL.n441 VTAIL.n440 0.155672
R909 VTAIL.n440 VTAIL.n404 0.155672
R910 VTAIL.n433 VTAIL.n404 0.155672
R911 VTAIL.n433 VTAIL.n432 0.155672
R912 VTAIL.n432 VTAIL.n408 0.155672
R913 VTAIL.n425 VTAIL.n408 0.155672
R914 VTAIL.n425 VTAIL.n424 0.155672
R915 VTAIL.n424 VTAIL.n412 0.155672
R916 VTAIL.n417 VTAIL.n412 0.155672
R917 VTAIL.n387 VTAIL.n313 0.155672
R918 VTAIL.n379 VTAIL.n313 0.155672
R919 VTAIL.n379 VTAIL.n378 0.155672
R920 VTAIL.n378 VTAIL.n318 0.155672
R921 VTAIL.n371 VTAIL.n318 0.155672
R922 VTAIL.n371 VTAIL.n370 0.155672
R923 VTAIL.n370 VTAIL.n322 0.155672
R924 VTAIL.n363 VTAIL.n322 0.155672
R925 VTAIL.n363 VTAIL.n362 0.155672
R926 VTAIL.n362 VTAIL.n326 0.155672
R927 VTAIL.n355 VTAIL.n326 0.155672
R928 VTAIL.n355 VTAIL.n354 0.155672
R929 VTAIL.n354 VTAIL.n330 0.155672
R930 VTAIL.n347 VTAIL.n330 0.155672
R931 VTAIL.n347 VTAIL.n346 0.155672
R932 VTAIL.n346 VTAIL.n334 0.155672
R933 VTAIL.n339 VTAIL.n334 0.155672
R934 VTAIL.n309 VTAIL.n235 0.155672
R935 VTAIL.n301 VTAIL.n235 0.155672
R936 VTAIL.n301 VTAIL.n300 0.155672
R937 VTAIL.n300 VTAIL.n240 0.155672
R938 VTAIL.n293 VTAIL.n240 0.155672
R939 VTAIL.n293 VTAIL.n292 0.155672
R940 VTAIL.n292 VTAIL.n244 0.155672
R941 VTAIL.n285 VTAIL.n244 0.155672
R942 VTAIL.n285 VTAIL.n284 0.155672
R943 VTAIL.n284 VTAIL.n248 0.155672
R944 VTAIL.n277 VTAIL.n248 0.155672
R945 VTAIL.n277 VTAIL.n276 0.155672
R946 VTAIL.n276 VTAIL.n252 0.155672
R947 VTAIL.n269 VTAIL.n252 0.155672
R948 VTAIL.n269 VTAIL.n268 0.155672
R949 VTAIL.n268 VTAIL.n256 0.155672
R950 VTAIL.n261 VTAIL.n256 0.155672
R951 VDD2.n2 VDD2.n0 113.225
R952 VDD2.n2 VDD2.n1 72.6917
R953 VDD2.n1 VDD2.t0 2.32395
R954 VDD2.n1 VDD2.t1 2.32395
R955 VDD2.n0 VDD2.t2 2.32395
R956 VDD2.n0 VDD2.t3 2.32395
R957 VDD2 VDD2.n2 0.0586897
R958 B.n355 B.n96 585
R959 B.n354 B.n353 585
R960 B.n352 B.n97 585
R961 B.n351 B.n350 585
R962 B.n349 B.n98 585
R963 B.n348 B.n347 585
R964 B.n346 B.n99 585
R965 B.n345 B.n344 585
R966 B.n343 B.n100 585
R967 B.n342 B.n341 585
R968 B.n340 B.n101 585
R969 B.n339 B.n338 585
R970 B.n337 B.n102 585
R971 B.n336 B.n335 585
R972 B.n334 B.n103 585
R973 B.n333 B.n332 585
R974 B.n331 B.n104 585
R975 B.n330 B.n329 585
R976 B.n328 B.n105 585
R977 B.n327 B.n326 585
R978 B.n325 B.n106 585
R979 B.n324 B.n323 585
R980 B.n322 B.n107 585
R981 B.n321 B.n320 585
R982 B.n319 B.n108 585
R983 B.n318 B.n317 585
R984 B.n316 B.n109 585
R985 B.n315 B.n314 585
R986 B.n313 B.n110 585
R987 B.n312 B.n311 585
R988 B.n310 B.n111 585
R989 B.n309 B.n308 585
R990 B.n307 B.n112 585
R991 B.n306 B.n305 585
R992 B.n304 B.n113 585
R993 B.n303 B.n302 585
R994 B.n301 B.n114 585
R995 B.n300 B.n299 585
R996 B.n298 B.n115 585
R997 B.n297 B.n296 585
R998 B.n295 B.n116 585
R999 B.n294 B.n293 585
R1000 B.n292 B.n117 585
R1001 B.n291 B.n290 585
R1002 B.n289 B.n118 585
R1003 B.n288 B.n287 585
R1004 B.n286 B.n119 585
R1005 B.n285 B.n284 585
R1006 B.n280 B.n120 585
R1007 B.n279 B.n278 585
R1008 B.n277 B.n121 585
R1009 B.n276 B.n275 585
R1010 B.n274 B.n122 585
R1011 B.n273 B.n272 585
R1012 B.n271 B.n123 585
R1013 B.n270 B.n269 585
R1014 B.n268 B.n124 585
R1015 B.n266 B.n265 585
R1016 B.n264 B.n127 585
R1017 B.n263 B.n262 585
R1018 B.n261 B.n128 585
R1019 B.n260 B.n259 585
R1020 B.n258 B.n129 585
R1021 B.n257 B.n256 585
R1022 B.n255 B.n130 585
R1023 B.n254 B.n253 585
R1024 B.n252 B.n131 585
R1025 B.n251 B.n250 585
R1026 B.n249 B.n132 585
R1027 B.n248 B.n247 585
R1028 B.n246 B.n133 585
R1029 B.n245 B.n244 585
R1030 B.n243 B.n134 585
R1031 B.n242 B.n241 585
R1032 B.n240 B.n135 585
R1033 B.n239 B.n238 585
R1034 B.n237 B.n136 585
R1035 B.n236 B.n235 585
R1036 B.n234 B.n137 585
R1037 B.n233 B.n232 585
R1038 B.n231 B.n138 585
R1039 B.n230 B.n229 585
R1040 B.n228 B.n139 585
R1041 B.n227 B.n226 585
R1042 B.n225 B.n140 585
R1043 B.n224 B.n223 585
R1044 B.n222 B.n141 585
R1045 B.n221 B.n220 585
R1046 B.n219 B.n142 585
R1047 B.n218 B.n217 585
R1048 B.n216 B.n143 585
R1049 B.n215 B.n214 585
R1050 B.n213 B.n144 585
R1051 B.n212 B.n211 585
R1052 B.n210 B.n145 585
R1053 B.n209 B.n208 585
R1054 B.n207 B.n146 585
R1055 B.n206 B.n205 585
R1056 B.n204 B.n147 585
R1057 B.n203 B.n202 585
R1058 B.n201 B.n148 585
R1059 B.n200 B.n199 585
R1060 B.n198 B.n149 585
R1061 B.n197 B.n196 585
R1062 B.n357 B.n356 585
R1063 B.n358 B.n95 585
R1064 B.n360 B.n359 585
R1065 B.n361 B.n94 585
R1066 B.n363 B.n362 585
R1067 B.n364 B.n93 585
R1068 B.n366 B.n365 585
R1069 B.n367 B.n92 585
R1070 B.n369 B.n368 585
R1071 B.n370 B.n91 585
R1072 B.n372 B.n371 585
R1073 B.n373 B.n90 585
R1074 B.n375 B.n374 585
R1075 B.n376 B.n89 585
R1076 B.n378 B.n377 585
R1077 B.n379 B.n88 585
R1078 B.n381 B.n380 585
R1079 B.n382 B.n87 585
R1080 B.n384 B.n383 585
R1081 B.n385 B.n86 585
R1082 B.n387 B.n386 585
R1083 B.n388 B.n85 585
R1084 B.n390 B.n389 585
R1085 B.n391 B.n84 585
R1086 B.n393 B.n392 585
R1087 B.n394 B.n83 585
R1088 B.n396 B.n395 585
R1089 B.n397 B.n82 585
R1090 B.n399 B.n398 585
R1091 B.n400 B.n81 585
R1092 B.n402 B.n401 585
R1093 B.n403 B.n80 585
R1094 B.n405 B.n404 585
R1095 B.n406 B.n79 585
R1096 B.n408 B.n407 585
R1097 B.n409 B.n78 585
R1098 B.n411 B.n410 585
R1099 B.n412 B.n77 585
R1100 B.n414 B.n413 585
R1101 B.n415 B.n76 585
R1102 B.n417 B.n416 585
R1103 B.n418 B.n75 585
R1104 B.n420 B.n419 585
R1105 B.n421 B.n74 585
R1106 B.n423 B.n422 585
R1107 B.n424 B.n73 585
R1108 B.n426 B.n425 585
R1109 B.n427 B.n72 585
R1110 B.n429 B.n428 585
R1111 B.n430 B.n71 585
R1112 B.n587 B.n14 585
R1113 B.n586 B.n585 585
R1114 B.n584 B.n15 585
R1115 B.n583 B.n582 585
R1116 B.n581 B.n16 585
R1117 B.n580 B.n579 585
R1118 B.n578 B.n17 585
R1119 B.n577 B.n576 585
R1120 B.n575 B.n18 585
R1121 B.n574 B.n573 585
R1122 B.n572 B.n19 585
R1123 B.n571 B.n570 585
R1124 B.n569 B.n20 585
R1125 B.n568 B.n567 585
R1126 B.n566 B.n21 585
R1127 B.n565 B.n564 585
R1128 B.n563 B.n22 585
R1129 B.n562 B.n561 585
R1130 B.n560 B.n23 585
R1131 B.n559 B.n558 585
R1132 B.n557 B.n24 585
R1133 B.n556 B.n555 585
R1134 B.n554 B.n25 585
R1135 B.n553 B.n552 585
R1136 B.n551 B.n26 585
R1137 B.n550 B.n549 585
R1138 B.n548 B.n27 585
R1139 B.n547 B.n546 585
R1140 B.n545 B.n28 585
R1141 B.n544 B.n543 585
R1142 B.n542 B.n29 585
R1143 B.n541 B.n540 585
R1144 B.n539 B.n30 585
R1145 B.n538 B.n537 585
R1146 B.n536 B.n31 585
R1147 B.n535 B.n534 585
R1148 B.n533 B.n32 585
R1149 B.n532 B.n531 585
R1150 B.n530 B.n33 585
R1151 B.n529 B.n528 585
R1152 B.n527 B.n34 585
R1153 B.n526 B.n525 585
R1154 B.n524 B.n35 585
R1155 B.n523 B.n522 585
R1156 B.n521 B.n36 585
R1157 B.n520 B.n519 585
R1158 B.n518 B.n37 585
R1159 B.n516 B.n515 585
R1160 B.n514 B.n40 585
R1161 B.n513 B.n512 585
R1162 B.n511 B.n41 585
R1163 B.n510 B.n509 585
R1164 B.n508 B.n42 585
R1165 B.n507 B.n506 585
R1166 B.n505 B.n43 585
R1167 B.n504 B.n503 585
R1168 B.n502 B.n44 585
R1169 B.n501 B.n500 585
R1170 B.n499 B.n45 585
R1171 B.n498 B.n497 585
R1172 B.n496 B.n49 585
R1173 B.n495 B.n494 585
R1174 B.n493 B.n50 585
R1175 B.n492 B.n491 585
R1176 B.n490 B.n51 585
R1177 B.n489 B.n488 585
R1178 B.n487 B.n52 585
R1179 B.n486 B.n485 585
R1180 B.n484 B.n53 585
R1181 B.n483 B.n482 585
R1182 B.n481 B.n54 585
R1183 B.n480 B.n479 585
R1184 B.n478 B.n55 585
R1185 B.n477 B.n476 585
R1186 B.n475 B.n56 585
R1187 B.n474 B.n473 585
R1188 B.n472 B.n57 585
R1189 B.n471 B.n470 585
R1190 B.n469 B.n58 585
R1191 B.n468 B.n467 585
R1192 B.n466 B.n59 585
R1193 B.n465 B.n464 585
R1194 B.n463 B.n60 585
R1195 B.n462 B.n461 585
R1196 B.n460 B.n61 585
R1197 B.n459 B.n458 585
R1198 B.n457 B.n62 585
R1199 B.n456 B.n455 585
R1200 B.n454 B.n63 585
R1201 B.n453 B.n452 585
R1202 B.n451 B.n64 585
R1203 B.n450 B.n449 585
R1204 B.n448 B.n65 585
R1205 B.n447 B.n446 585
R1206 B.n445 B.n66 585
R1207 B.n444 B.n443 585
R1208 B.n442 B.n67 585
R1209 B.n441 B.n440 585
R1210 B.n439 B.n68 585
R1211 B.n438 B.n437 585
R1212 B.n436 B.n69 585
R1213 B.n435 B.n434 585
R1214 B.n433 B.n70 585
R1215 B.n432 B.n431 585
R1216 B.n589 B.n588 585
R1217 B.n590 B.n13 585
R1218 B.n592 B.n591 585
R1219 B.n593 B.n12 585
R1220 B.n595 B.n594 585
R1221 B.n596 B.n11 585
R1222 B.n598 B.n597 585
R1223 B.n599 B.n10 585
R1224 B.n601 B.n600 585
R1225 B.n602 B.n9 585
R1226 B.n604 B.n603 585
R1227 B.n605 B.n8 585
R1228 B.n607 B.n606 585
R1229 B.n608 B.n7 585
R1230 B.n610 B.n609 585
R1231 B.n611 B.n6 585
R1232 B.n613 B.n612 585
R1233 B.n614 B.n5 585
R1234 B.n616 B.n615 585
R1235 B.n617 B.n4 585
R1236 B.n619 B.n618 585
R1237 B.n620 B.n3 585
R1238 B.n622 B.n621 585
R1239 B.n623 B.n0 585
R1240 B.n2 B.n1 585
R1241 B.n162 B.n161 585
R1242 B.n164 B.n163 585
R1243 B.n165 B.n160 585
R1244 B.n167 B.n166 585
R1245 B.n168 B.n159 585
R1246 B.n170 B.n169 585
R1247 B.n171 B.n158 585
R1248 B.n173 B.n172 585
R1249 B.n174 B.n157 585
R1250 B.n176 B.n175 585
R1251 B.n177 B.n156 585
R1252 B.n179 B.n178 585
R1253 B.n180 B.n155 585
R1254 B.n182 B.n181 585
R1255 B.n183 B.n154 585
R1256 B.n185 B.n184 585
R1257 B.n186 B.n153 585
R1258 B.n188 B.n187 585
R1259 B.n189 B.n152 585
R1260 B.n191 B.n190 585
R1261 B.n192 B.n151 585
R1262 B.n194 B.n193 585
R1263 B.n195 B.n150 585
R1264 B.n197 B.n150 516.524
R1265 B.n357 B.n96 516.524
R1266 B.n431 B.n430 516.524
R1267 B.n588 B.n587 516.524
R1268 B.n281 B.t1 446.988
R1269 B.n46 B.t8 446.988
R1270 B.n125 B.t4 446.988
R1271 B.n38 B.t11 446.988
R1272 B.n125 B.t3 428.762
R1273 B.n281 B.t0 428.762
R1274 B.n46 B.t6 428.762
R1275 B.n38 B.t9 428.762
R1276 B.n282 B.t2 411.303
R1277 B.n47 B.t7 411.303
R1278 B.n126 B.t5 411.303
R1279 B.n39 B.t10 411.303
R1280 B.n625 B.n624 256.663
R1281 B.n624 B.n623 235.042
R1282 B.n624 B.n2 235.042
R1283 B.n198 B.n197 163.367
R1284 B.n199 B.n198 163.367
R1285 B.n199 B.n148 163.367
R1286 B.n203 B.n148 163.367
R1287 B.n204 B.n203 163.367
R1288 B.n205 B.n204 163.367
R1289 B.n205 B.n146 163.367
R1290 B.n209 B.n146 163.367
R1291 B.n210 B.n209 163.367
R1292 B.n211 B.n210 163.367
R1293 B.n211 B.n144 163.367
R1294 B.n215 B.n144 163.367
R1295 B.n216 B.n215 163.367
R1296 B.n217 B.n216 163.367
R1297 B.n217 B.n142 163.367
R1298 B.n221 B.n142 163.367
R1299 B.n222 B.n221 163.367
R1300 B.n223 B.n222 163.367
R1301 B.n223 B.n140 163.367
R1302 B.n227 B.n140 163.367
R1303 B.n228 B.n227 163.367
R1304 B.n229 B.n228 163.367
R1305 B.n229 B.n138 163.367
R1306 B.n233 B.n138 163.367
R1307 B.n234 B.n233 163.367
R1308 B.n235 B.n234 163.367
R1309 B.n235 B.n136 163.367
R1310 B.n239 B.n136 163.367
R1311 B.n240 B.n239 163.367
R1312 B.n241 B.n240 163.367
R1313 B.n241 B.n134 163.367
R1314 B.n245 B.n134 163.367
R1315 B.n246 B.n245 163.367
R1316 B.n247 B.n246 163.367
R1317 B.n247 B.n132 163.367
R1318 B.n251 B.n132 163.367
R1319 B.n252 B.n251 163.367
R1320 B.n253 B.n252 163.367
R1321 B.n253 B.n130 163.367
R1322 B.n257 B.n130 163.367
R1323 B.n258 B.n257 163.367
R1324 B.n259 B.n258 163.367
R1325 B.n259 B.n128 163.367
R1326 B.n263 B.n128 163.367
R1327 B.n264 B.n263 163.367
R1328 B.n265 B.n264 163.367
R1329 B.n265 B.n124 163.367
R1330 B.n270 B.n124 163.367
R1331 B.n271 B.n270 163.367
R1332 B.n272 B.n271 163.367
R1333 B.n272 B.n122 163.367
R1334 B.n276 B.n122 163.367
R1335 B.n277 B.n276 163.367
R1336 B.n278 B.n277 163.367
R1337 B.n278 B.n120 163.367
R1338 B.n285 B.n120 163.367
R1339 B.n286 B.n285 163.367
R1340 B.n287 B.n286 163.367
R1341 B.n287 B.n118 163.367
R1342 B.n291 B.n118 163.367
R1343 B.n292 B.n291 163.367
R1344 B.n293 B.n292 163.367
R1345 B.n293 B.n116 163.367
R1346 B.n297 B.n116 163.367
R1347 B.n298 B.n297 163.367
R1348 B.n299 B.n298 163.367
R1349 B.n299 B.n114 163.367
R1350 B.n303 B.n114 163.367
R1351 B.n304 B.n303 163.367
R1352 B.n305 B.n304 163.367
R1353 B.n305 B.n112 163.367
R1354 B.n309 B.n112 163.367
R1355 B.n310 B.n309 163.367
R1356 B.n311 B.n310 163.367
R1357 B.n311 B.n110 163.367
R1358 B.n315 B.n110 163.367
R1359 B.n316 B.n315 163.367
R1360 B.n317 B.n316 163.367
R1361 B.n317 B.n108 163.367
R1362 B.n321 B.n108 163.367
R1363 B.n322 B.n321 163.367
R1364 B.n323 B.n322 163.367
R1365 B.n323 B.n106 163.367
R1366 B.n327 B.n106 163.367
R1367 B.n328 B.n327 163.367
R1368 B.n329 B.n328 163.367
R1369 B.n329 B.n104 163.367
R1370 B.n333 B.n104 163.367
R1371 B.n334 B.n333 163.367
R1372 B.n335 B.n334 163.367
R1373 B.n335 B.n102 163.367
R1374 B.n339 B.n102 163.367
R1375 B.n340 B.n339 163.367
R1376 B.n341 B.n340 163.367
R1377 B.n341 B.n100 163.367
R1378 B.n345 B.n100 163.367
R1379 B.n346 B.n345 163.367
R1380 B.n347 B.n346 163.367
R1381 B.n347 B.n98 163.367
R1382 B.n351 B.n98 163.367
R1383 B.n352 B.n351 163.367
R1384 B.n353 B.n352 163.367
R1385 B.n353 B.n96 163.367
R1386 B.n430 B.n429 163.367
R1387 B.n429 B.n72 163.367
R1388 B.n425 B.n72 163.367
R1389 B.n425 B.n424 163.367
R1390 B.n424 B.n423 163.367
R1391 B.n423 B.n74 163.367
R1392 B.n419 B.n74 163.367
R1393 B.n419 B.n418 163.367
R1394 B.n418 B.n417 163.367
R1395 B.n417 B.n76 163.367
R1396 B.n413 B.n76 163.367
R1397 B.n413 B.n412 163.367
R1398 B.n412 B.n411 163.367
R1399 B.n411 B.n78 163.367
R1400 B.n407 B.n78 163.367
R1401 B.n407 B.n406 163.367
R1402 B.n406 B.n405 163.367
R1403 B.n405 B.n80 163.367
R1404 B.n401 B.n80 163.367
R1405 B.n401 B.n400 163.367
R1406 B.n400 B.n399 163.367
R1407 B.n399 B.n82 163.367
R1408 B.n395 B.n82 163.367
R1409 B.n395 B.n394 163.367
R1410 B.n394 B.n393 163.367
R1411 B.n393 B.n84 163.367
R1412 B.n389 B.n84 163.367
R1413 B.n389 B.n388 163.367
R1414 B.n388 B.n387 163.367
R1415 B.n387 B.n86 163.367
R1416 B.n383 B.n86 163.367
R1417 B.n383 B.n382 163.367
R1418 B.n382 B.n381 163.367
R1419 B.n381 B.n88 163.367
R1420 B.n377 B.n88 163.367
R1421 B.n377 B.n376 163.367
R1422 B.n376 B.n375 163.367
R1423 B.n375 B.n90 163.367
R1424 B.n371 B.n90 163.367
R1425 B.n371 B.n370 163.367
R1426 B.n370 B.n369 163.367
R1427 B.n369 B.n92 163.367
R1428 B.n365 B.n92 163.367
R1429 B.n365 B.n364 163.367
R1430 B.n364 B.n363 163.367
R1431 B.n363 B.n94 163.367
R1432 B.n359 B.n94 163.367
R1433 B.n359 B.n358 163.367
R1434 B.n358 B.n357 163.367
R1435 B.n587 B.n586 163.367
R1436 B.n586 B.n15 163.367
R1437 B.n582 B.n15 163.367
R1438 B.n582 B.n581 163.367
R1439 B.n581 B.n580 163.367
R1440 B.n580 B.n17 163.367
R1441 B.n576 B.n17 163.367
R1442 B.n576 B.n575 163.367
R1443 B.n575 B.n574 163.367
R1444 B.n574 B.n19 163.367
R1445 B.n570 B.n19 163.367
R1446 B.n570 B.n569 163.367
R1447 B.n569 B.n568 163.367
R1448 B.n568 B.n21 163.367
R1449 B.n564 B.n21 163.367
R1450 B.n564 B.n563 163.367
R1451 B.n563 B.n562 163.367
R1452 B.n562 B.n23 163.367
R1453 B.n558 B.n23 163.367
R1454 B.n558 B.n557 163.367
R1455 B.n557 B.n556 163.367
R1456 B.n556 B.n25 163.367
R1457 B.n552 B.n25 163.367
R1458 B.n552 B.n551 163.367
R1459 B.n551 B.n550 163.367
R1460 B.n550 B.n27 163.367
R1461 B.n546 B.n27 163.367
R1462 B.n546 B.n545 163.367
R1463 B.n545 B.n544 163.367
R1464 B.n544 B.n29 163.367
R1465 B.n540 B.n29 163.367
R1466 B.n540 B.n539 163.367
R1467 B.n539 B.n538 163.367
R1468 B.n538 B.n31 163.367
R1469 B.n534 B.n31 163.367
R1470 B.n534 B.n533 163.367
R1471 B.n533 B.n532 163.367
R1472 B.n532 B.n33 163.367
R1473 B.n528 B.n33 163.367
R1474 B.n528 B.n527 163.367
R1475 B.n527 B.n526 163.367
R1476 B.n526 B.n35 163.367
R1477 B.n522 B.n35 163.367
R1478 B.n522 B.n521 163.367
R1479 B.n521 B.n520 163.367
R1480 B.n520 B.n37 163.367
R1481 B.n515 B.n37 163.367
R1482 B.n515 B.n514 163.367
R1483 B.n514 B.n513 163.367
R1484 B.n513 B.n41 163.367
R1485 B.n509 B.n41 163.367
R1486 B.n509 B.n508 163.367
R1487 B.n508 B.n507 163.367
R1488 B.n507 B.n43 163.367
R1489 B.n503 B.n43 163.367
R1490 B.n503 B.n502 163.367
R1491 B.n502 B.n501 163.367
R1492 B.n501 B.n45 163.367
R1493 B.n497 B.n45 163.367
R1494 B.n497 B.n496 163.367
R1495 B.n496 B.n495 163.367
R1496 B.n495 B.n50 163.367
R1497 B.n491 B.n50 163.367
R1498 B.n491 B.n490 163.367
R1499 B.n490 B.n489 163.367
R1500 B.n489 B.n52 163.367
R1501 B.n485 B.n52 163.367
R1502 B.n485 B.n484 163.367
R1503 B.n484 B.n483 163.367
R1504 B.n483 B.n54 163.367
R1505 B.n479 B.n54 163.367
R1506 B.n479 B.n478 163.367
R1507 B.n478 B.n477 163.367
R1508 B.n477 B.n56 163.367
R1509 B.n473 B.n56 163.367
R1510 B.n473 B.n472 163.367
R1511 B.n472 B.n471 163.367
R1512 B.n471 B.n58 163.367
R1513 B.n467 B.n58 163.367
R1514 B.n467 B.n466 163.367
R1515 B.n466 B.n465 163.367
R1516 B.n465 B.n60 163.367
R1517 B.n461 B.n60 163.367
R1518 B.n461 B.n460 163.367
R1519 B.n460 B.n459 163.367
R1520 B.n459 B.n62 163.367
R1521 B.n455 B.n62 163.367
R1522 B.n455 B.n454 163.367
R1523 B.n454 B.n453 163.367
R1524 B.n453 B.n64 163.367
R1525 B.n449 B.n64 163.367
R1526 B.n449 B.n448 163.367
R1527 B.n448 B.n447 163.367
R1528 B.n447 B.n66 163.367
R1529 B.n443 B.n66 163.367
R1530 B.n443 B.n442 163.367
R1531 B.n442 B.n441 163.367
R1532 B.n441 B.n68 163.367
R1533 B.n437 B.n68 163.367
R1534 B.n437 B.n436 163.367
R1535 B.n436 B.n435 163.367
R1536 B.n435 B.n70 163.367
R1537 B.n431 B.n70 163.367
R1538 B.n588 B.n13 163.367
R1539 B.n592 B.n13 163.367
R1540 B.n593 B.n592 163.367
R1541 B.n594 B.n593 163.367
R1542 B.n594 B.n11 163.367
R1543 B.n598 B.n11 163.367
R1544 B.n599 B.n598 163.367
R1545 B.n600 B.n599 163.367
R1546 B.n600 B.n9 163.367
R1547 B.n604 B.n9 163.367
R1548 B.n605 B.n604 163.367
R1549 B.n606 B.n605 163.367
R1550 B.n606 B.n7 163.367
R1551 B.n610 B.n7 163.367
R1552 B.n611 B.n610 163.367
R1553 B.n612 B.n611 163.367
R1554 B.n612 B.n5 163.367
R1555 B.n616 B.n5 163.367
R1556 B.n617 B.n616 163.367
R1557 B.n618 B.n617 163.367
R1558 B.n618 B.n3 163.367
R1559 B.n622 B.n3 163.367
R1560 B.n623 B.n622 163.367
R1561 B.n162 B.n2 163.367
R1562 B.n163 B.n162 163.367
R1563 B.n163 B.n160 163.367
R1564 B.n167 B.n160 163.367
R1565 B.n168 B.n167 163.367
R1566 B.n169 B.n168 163.367
R1567 B.n169 B.n158 163.367
R1568 B.n173 B.n158 163.367
R1569 B.n174 B.n173 163.367
R1570 B.n175 B.n174 163.367
R1571 B.n175 B.n156 163.367
R1572 B.n179 B.n156 163.367
R1573 B.n180 B.n179 163.367
R1574 B.n181 B.n180 163.367
R1575 B.n181 B.n154 163.367
R1576 B.n185 B.n154 163.367
R1577 B.n186 B.n185 163.367
R1578 B.n187 B.n186 163.367
R1579 B.n187 B.n152 163.367
R1580 B.n191 B.n152 163.367
R1581 B.n192 B.n191 163.367
R1582 B.n193 B.n192 163.367
R1583 B.n193 B.n150 163.367
R1584 B.n267 B.n126 59.5399
R1585 B.n283 B.n282 59.5399
R1586 B.n48 B.n47 59.5399
R1587 B.n517 B.n39 59.5399
R1588 B.n126 B.n125 35.6853
R1589 B.n282 B.n281 35.6853
R1590 B.n47 B.n46 35.6853
R1591 B.n39 B.n38 35.6853
R1592 B.n589 B.n14 33.5615
R1593 B.n432 B.n71 33.5615
R1594 B.n356 B.n355 33.5615
R1595 B.n196 B.n195 33.5615
R1596 B B.n625 18.0485
R1597 B.n590 B.n589 10.6151
R1598 B.n591 B.n590 10.6151
R1599 B.n591 B.n12 10.6151
R1600 B.n595 B.n12 10.6151
R1601 B.n596 B.n595 10.6151
R1602 B.n597 B.n596 10.6151
R1603 B.n597 B.n10 10.6151
R1604 B.n601 B.n10 10.6151
R1605 B.n602 B.n601 10.6151
R1606 B.n603 B.n602 10.6151
R1607 B.n603 B.n8 10.6151
R1608 B.n607 B.n8 10.6151
R1609 B.n608 B.n607 10.6151
R1610 B.n609 B.n608 10.6151
R1611 B.n609 B.n6 10.6151
R1612 B.n613 B.n6 10.6151
R1613 B.n614 B.n613 10.6151
R1614 B.n615 B.n614 10.6151
R1615 B.n615 B.n4 10.6151
R1616 B.n619 B.n4 10.6151
R1617 B.n620 B.n619 10.6151
R1618 B.n621 B.n620 10.6151
R1619 B.n621 B.n0 10.6151
R1620 B.n585 B.n14 10.6151
R1621 B.n585 B.n584 10.6151
R1622 B.n584 B.n583 10.6151
R1623 B.n583 B.n16 10.6151
R1624 B.n579 B.n16 10.6151
R1625 B.n579 B.n578 10.6151
R1626 B.n578 B.n577 10.6151
R1627 B.n577 B.n18 10.6151
R1628 B.n573 B.n18 10.6151
R1629 B.n573 B.n572 10.6151
R1630 B.n572 B.n571 10.6151
R1631 B.n571 B.n20 10.6151
R1632 B.n567 B.n20 10.6151
R1633 B.n567 B.n566 10.6151
R1634 B.n566 B.n565 10.6151
R1635 B.n565 B.n22 10.6151
R1636 B.n561 B.n22 10.6151
R1637 B.n561 B.n560 10.6151
R1638 B.n560 B.n559 10.6151
R1639 B.n559 B.n24 10.6151
R1640 B.n555 B.n24 10.6151
R1641 B.n555 B.n554 10.6151
R1642 B.n554 B.n553 10.6151
R1643 B.n553 B.n26 10.6151
R1644 B.n549 B.n26 10.6151
R1645 B.n549 B.n548 10.6151
R1646 B.n548 B.n547 10.6151
R1647 B.n547 B.n28 10.6151
R1648 B.n543 B.n28 10.6151
R1649 B.n543 B.n542 10.6151
R1650 B.n542 B.n541 10.6151
R1651 B.n541 B.n30 10.6151
R1652 B.n537 B.n30 10.6151
R1653 B.n537 B.n536 10.6151
R1654 B.n536 B.n535 10.6151
R1655 B.n535 B.n32 10.6151
R1656 B.n531 B.n32 10.6151
R1657 B.n531 B.n530 10.6151
R1658 B.n530 B.n529 10.6151
R1659 B.n529 B.n34 10.6151
R1660 B.n525 B.n34 10.6151
R1661 B.n525 B.n524 10.6151
R1662 B.n524 B.n523 10.6151
R1663 B.n523 B.n36 10.6151
R1664 B.n519 B.n36 10.6151
R1665 B.n519 B.n518 10.6151
R1666 B.n516 B.n40 10.6151
R1667 B.n512 B.n40 10.6151
R1668 B.n512 B.n511 10.6151
R1669 B.n511 B.n510 10.6151
R1670 B.n510 B.n42 10.6151
R1671 B.n506 B.n42 10.6151
R1672 B.n506 B.n505 10.6151
R1673 B.n505 B.n504 10.6151
R1674 B.n504 B.n44 10.6151
R1675 B.n500 B.n499 10.6151
R1676 B.n499 B.n498 10.6151
R1677 B.n498 B.n49 10.6151
R1678 B.n494 B.n49 10.6151
R1679 B.n494 B.n493 10.6151
R1680 B.n493 B.n492 10.6151
R1681 B.n492 B.n51 10.6151
R1682 B.n488 B.n51 10.6151
R1683 B.n488 B.n487 10.6151
R1684 B.n487 B.n486 10.6151
R1685 B.n486 B.n53 10.6151
R1686 B.n482 B.n53 10.6151
R1687 B.n482 B.n481 10.6151
R1688 B.n481 B.n480 10.6151
R1689 B.n480 B.n55 10.6151
R1690 B.n476 B.n55 10.6151
R1691 B.n476 B.n475 10.6151
R1692 B.n475 B.n474 10.6151
R1693 B.n474 B.n57 10.6151
R1694 B.n470 B.n57 10.6151
R1695 B.n470 B.n469 10.6151
R1696 B.n469 B.n468 10.6151
R1697 B.n468 B.n59 10.6151
R1698 B.n464 B.n59 10.6151
R1699 B.n464 B.n463 10.6151
R1700 B.n463 B.n462 10.6151
R1701 B.n462 B.n61 10.6151
R1702 B.n458 B.n61 10.6151
R1703 B.n458 B.n457 10.6151
R1704 B.n457 B.n456 10.6151
R1705 B.n456 B.n63 10.6151
R1706 B.n452 B.n63 10.6151
R1707 B.n452 B.n451 10.6151
R1708 B.n451 B.n450 10.6151
R1709 B.n450 B.n65 10.6151
R1710 B.n446 B.n65 10.6151
R1711 B.n446 B.n445 10.6151
R1712 B.n445 B.n444 10.6151
R1713 B.n444 B.n67 10.6151
R1714 B.n440 B.n67 10.6151
R1715 B.n440 B.n439 10.6151
R1716 B.n439 B.n438 10.6151
R1717 B.n438 B.n69 10.6151
R1718 B.n434 B.n69 10.6151
R1719 B.n434 B.n433 10.6151
R1720 B.n433 B.n432 10.6151
R1721 B.n428 B.n71 10.6151
R1722 B.n428 B.n427 10.6151
R1723 B.n427 B.n426 10.6151
R1724 B.n426 B.n73 10.6151
R1725 B.n422 B.n73 10.6151
R1726 B.n422 B.n421 10.6151
R1727 B.n421 B.n420 10.6151
R1728 B.n420 B.n75 10.6151
R1729 B.n416 B.n75 10.6151
R1730 B.n416 B.n415 10.6151
R1731 B.n415 B.n414 10.6151
R1732 B.n414 B.n77 10.6151
R1733 B.n410 B.n77 10.6151
R1734 B.n410 B.n409 10.6151
R1735 B.n409 B.n408 10.6151
R1736 B.n408 B.n79 10.6151
R1737 B.n404 B.n79 10.6151
R1738 B.n404 B.n403 10.6151
R1739 B.n403 B.n402 10.6151
R1740 B.n402 B.n81 10.6151
R1741 B.n398 B.n81 10.6151
R1742 B.n398 B.n397 10.6151
R1743 B.n397 B.n396 10.6151
R1744 B.n396 B.n83 10.6151
R1745 B.n392 B.n83 10.6151
R1746 B.n392 B.n391 10.6151
R1747 B.n391 B.n390 10.6151
R1748 B.n390 B.n85 10.6151
R1749 B.n386 B.n85 10.6151
R1750 B.n386 B.n385 10.6151
R1751 B.n385 B.n384 10.6151
R1752 B.n384 B.n87 10.6151
R1753 B.n380 B.n87 10.6151
R1754 B.n380 B.n379 10.6151
R1755 B.n379 B.n378 10.6151
R1756 B.n378 B.n89 10.6151
R1757 B.n374 B.n89 10.6151
R1758 B.n374 B.n373 10.6151
R1759 B.n373 B.n372 10.6151
R1760 B.n372 B.n91 10.6151
R1761 B.n368 B.n91 10.6151
R1762 B.n368 B.n367 10.6151
R1763 B.n367 B.n366 10.6151
R1764 B.n366 B.n93 10.6151
R1765 B.n362 B.n93 10.6151
R1766 B.n362 B.n361 10.6151
R1767 B.n361 B.n360 10.6151
R1768 B.n360 B.n95 10.6151
R1769 B.n356 B.n95 10.6151
R1770 B.n161 B.n1 10.6151
R1771 B.n164 B.n161 10.6151
R1772 B.n165 B.n164 10.6151
R1773 B.n166 B.n165 10.6151
R1774 B.n166 B.n159 10.6151
R1775 B.n170 B.n159 10.6151
R1776 B.n171 B.n170 10.6151
R1777 B.n172 B.n171 10.6151
R1778 B.n172 B.n157 10.6151
R1779 B.n176 B.n157 10.6151
R1780 B.n177 B.n176 10.6151
R1781 B.n178 B.n177 10.6151
R1782 B.n178 B.n155 10.6151
R1783 B.n182 B.n155 10.6151
R1784 B.n183 B.n182 10.6151
R1785 B.n184 B.n183 10.6151
R1786 B.n184 B.n153 10.6151
R1787 B.n188 B.n153 10.6151
R1788 B.n189 B.n188 10.6151
R1789 B.n190 B.n189 10.6151
R1790 B.n190 B.n151 10.6151
R1791 B.n194 B.n151 10.6151
R1792 B.n195 B.n194 10.6151
R1793 B.n196 B.n149 10.6151
R1794 B.n200 B.n149 10.6151
R1795 B.n201 B.n200 10.6151
R1796 B.n202 B.n201 10.6151
R1797 B.n202 B.n147 10.6151
R1798 B.n206 B.n147 10.6151
R1799 B.n207 B.n206 10.6151
R1800 B.n208 B.n207 10.6151
R1801 B.n208 B.n145 10.6151
R1802 B.n212 B.n145 10.6151
R1803 B.n213 B.n212 10.6151
R1804 B.n214 B.n213 10.6151
R1805 B.n214 B.n143 10.6151
R1806 B.n218 B.n143 10.6151
R1807 B.n219 B.n218 10.6151
R1808 B.n220 B.n219 10.6151
R1809 B.n220 B.n141 10.6151
R1810 B.n224 B.n141 10.6151
R1811 B.n225 B.n224 10.6151
R1812 B.n226 B.n225 10.6151
R1813 B.n226 B.n139 10.6151
R1814 B.n230 B.n139 10.6151
R1815 B.n231 B.n230 10.6151
R1816 B.n232 B.n231 10.6151
R1817 B.n232 B.n137 10.6151
R1818 B.n236 B.n137 10.6151
R1819 B.n237 B.n236 10.6151
R1820 B.n238 B.n237 10.6151
R1821 B.n238 B.n135 10.6151
R1822 B.n242 B.n135 10.6151
R1823 B.n243 B.n242 10.6151
R1824 B.n244 B.n243 10.6151
R1825 B.n244 B.n133 10.6151
R1826 B.n248 B.n133 10.6151
R1827 B.n249 B.n248 10.6151
R1828 B.n250 B.n249 10.6151
R1829 B.n250 B.n131 10.6151
R1830 B.n254 B.n131 10.6151
R1831 B.n255 B.n254 10.6151
R1832 B.n256 B.n255 10.6151
R1833 B.n256 B.n129 10.6151
R1834 B.n260 B.n129 10.6151
R1835 B.n261 B.n260 10.6151
R1836 B.n262 B.n261 10.6151
R1837 B.n262 B.n127 10.6151
R1838 B.n266 B.n127 10.6151
R1839 B.n269 B.n268 10.6151
R1840 B.n269 B.n123 10.6151
R1841 B.n273 B.n123 10.6151
R1842 B.n274 B.n273 10.6151
R1843 B.n275 B.n274 10.6151
R1844 B.n275 B.n121 10.6151
R1845 B.n279 B.n121 10.6151
R1846 B.n280 B.n279 10.6151
R1847 B.n284 B.n280 10.6151
R1848 B.n288 B.n119 10.6151
R1849 B.n289 B.n288 10.6151
R1850 B.n290 B.n289 10.6151
R1851 B.n290 B.n117 10.6151
R1852 B.n294 B.n117 10.6151
R1853 B.n295 B.n294 10.6151
R1854 B.n296 B.n295 10.6151
R1855 B.n296 B.n115 10.6151
R1856 B.n300 B.n115 10.6151
R1857 B.n301 B.n300 10.6151
R1858 B.n302 B.n301 10.6151
R1859 B.n302 B.n113 10.6151
R1860 B.n306 B.n113 10.6151
R1861 B.n307 B.n306 10.6151
R1862 B.n308 B.n307 10.6151
R1863 B.n308 B.n111 10.6151
R1864 B.n312 B.n111 10.6151
R1865 B.n313 B.n312 10.6151
R1866 B.n314 B.n313 10.6151
R1867 B.n314 B.n109 10.6151
R1868 B.n318 B.n109 10.6151
R1869 B.n319 B.n318 10.6151
R1870 B.n320 B.n319 10.6151
R1871 B.n320 B.n107 10.6151
R1872 B.n324 B.n107 10.6151
R1873 B.n325 B.n324 10.6151
R1874 B.n326 B.n325 10.6151
R1875 B.n326 B.n105 10.6151
R1876 B.n330 B.n105 10.6151
R1877 B.n331 B.n330 10.6151
R1878 B.n332 B.n331 10.6151
R1879 B.n332 B.n103 10.6151
R1880 B.n336 B.n103 10.6151
R1881 B.n337 B.n336 10.6151
R1882 B.n338 B.n337 10.6151
R1883 B.n338 B.n101 10.6151
R1884 B.n342 B.n101 10.6151
R1885 B.n343 B.n342 10.6151
R1886 B.n344 B.n343 10.6151
R1887 B.n344 B.n99 10.6151
R1888 B.n348 B.n99 10.6151
R1889 B.n349 B.n348 10.6151
R1890 B.n350 B.n349 10.6151
R1891 B.n350 B.n97 10.6151
R1892 B.n354 B.n97 10.6151
R1893 B.n355 B.n354 10.6151
R1894 B.n518 B.n517 9.36635
R1895 B.n500 B.n48 9.36635
R1896 B.n267 B.n266 9.36635
R1897 B.n283 B.n119 9.36635
R1898 B.n625 B.n0 8.11757
R1899 B.n625 B.n1 8.11757
R1900 B.n517 B.n516 1.24928
R1901 B.n48 B.n44 1.24928
R1902 B.n268 B.n267 1.24928
R1903 B.n284 B.n283 1.24928
R1904 VP.n2 VP.t1 259.791
R1905 VP.n2 VP.t3 259.474
R1906 VP.n4 VP.t0 223.285
R1907 VP.n11 VP.t2 223.285
R1908 VP.n4 VP.n3 177.448
R1909 VP.n12 VP.n11 177.448
R1910 VP.n10 VP.n0 161.3
R1911 VP.n9 VP.n8 161.3
R1912 VP.n7 VP.n1 161.3
R1913 VP.n6 VP.n5 161.3
R1914 VP.n3 VP.n2 57.3946
R1915 VP.n9 VP.n1 56.5193
R1916 VP.n5 VP.n1 24.4675
R1917 VP.n10 VP.n9 24.4675
R1918 VP.n5 VP.n4 8.31928
R1919 VP.n11 VP.n10 8.31928
R1920 VP.n6 VP.n3 0.189894
R1921 VP.n7 VP.n6 0.189894
R1922 VP.n8 VP.n7 0.189894
R1923 VP.n8 VP.n0 0.189894
R1924 VP.n12 VP.n0 0.189894
R1925 VP VP.n12 0.0516364
R1926 VDD1 VDD1.n1 113.751
R1927 VDD1 VDD1.n0 72.7499
R1928 VDD1.n0 VDD1.t2 2.32395
R1929 VDD1.n0 VDD1.t0 2.32395
R1930 VDD1.n1 VDD1.t3 2.32395
R1931 VDD1.n1 VDD1.t1 2.32395
C0 VDD1 VDD2 0.76218f
C1 VDD1 VP 5.01267f
C2 w_n2074_n3766# VN 3.34862f
C3 VN B 0.925136f
C4 VP VDD2 0.325065f
C5 VDD1 w_n2074_n3766# 1.29307f
C6 VTAIL VN 4.5045f
C7 VDD1 B 1.12347f
C8 w_n2074_n3766# VDD2 1.32485f
C9 VDD1 VTAIL 6.1252f
C10 w_n2074_n3766# VP 3.61248f
C11 VDD2 B 1.15783f
C12 VP B 1.35793f
C13 VTAIL VDD2 6.1721f
C14 VTAIL VP 4.51861f
C15 VDD1 VN 0.148133f
C16 w_n2074_n3766# B 8.462411f
C17 VTAIL w_n2074_n3766# 4.49092f
C18 VDD2 VN 4.8362f
C19 VP VN 5.77469f
C20 VTAIL B 4.97966f
C21 VDD2 VSUBS 0.829149f
C22 VDD1 VSUBS 5.402387f
C23 VTAIL VSUBS 1.144757f
C24 VN VSUBS 5.26214f
C25 VP VSUBS 1.775647f
C26 B VSUBS 3.50201f
C27 w_n2074_n3766# VSUBS 95.8935f
C28 VDD1.t2 VSUBS 0.294755f
C29 VDD1.t0 VSUBS 0.294755f
C30 VDD1.n0 VSUBS 2.37358f
C31 VDD1.t3 VSUBS 0.294755f
C32 VDD1.t1 VSUBS 0.294755f
C33 VDD1.n1 VSUBS 3.11509f
C34 VP.n0 VSUBS 0.043435f
C35 VP.t2 VSUBS 2.51014f
C36 VP.n1 VSUBS 0.063407f
C37 VP.t1 VSUBS 2.66087f
C38 VP.t3 VSUBS 2.65953f
C39 VP.n2 VSUBS 3.61367f
C40 VP.n3 VSUBS 2.50693f
C41 VP.t0 VSUBS 2.51014f
C42 VP.n4 VSUBS 0.983766f
C43 VP.n5 VSUBS 0.054574f
C44 VP.n6 VSUBS 0.043435f
C45 VP.n7 VSUBS 0.043435f
C46 VP.n8 VSUBS 0.043435f
C47 VP.n9 VSUBS 0.063407f
C48 VP.n10 VSUBS 0.054574f
C49 VP.n11 VSUBS 0.983766f
C50 VP.n12 VSUBS 0.042336f
C51 B.n0 VSUBS 0.006385f
C52 B.n1 VSUBS 0.006385f
C53 B.n2 VSUBS 0.009443f
C54 B.n3 VSUBS 0.007237f
C55 B.n4 VSUBS 0.007237f
C56 B.n5 VSUBS 0.007237f
C57 B.n6 VSUBS 0.007237f
C58 B.n7 VSUBS 0.007237f
C59 B.n8 VSUBS 0.007237f
C60 B.n9 VSUBS 0.007237f
C61 B.n10 VSUBS 0.007237f
C62 B.n11 VSUBS 0.007237f
C63 B.n12 VSUBS 0.007237f
C64 B.n13 VSUBS 0.007237f
C65 B.n14 VSUBS 0.017352f
C66 B.n15 VSUBS 0.007237f
C67 B.n16 VSUBS 0.007237f
C68 B.n17 VSUBS 0.007237f
C69 B.n18 VSUBS 0.007237f
C70 B.n19 VSUBS 0.007237f
C71 B.n20 VSUBS 0.007237f
C72 B.n21 VSUBS 0.007237f
C73 B.n22 VSUBS 0.007237f
C74 B.n23 VSUBS 0.007237f
C75 B.n24 VSUBS 0.007237f
C76 B.n25 VSUBS 0.007237f
C77 B.n26 VSUBS 0.007237f
C78 B.n27 VSUBS 0.007237f
C79 B.n28 VSUBS 0.007237f
C80 B.n29 VSUBS 0.007237f
C81 B.n30 VSUBS 0.007237f
C82 B.n31 VSUBS 0.007237f
C83 B.n32 VSUBS 0.007237f
C84 B.n33 VSUBS 0.007237f
C85 B.n34 VSUBS 0.007237f
C86 B.n35 VSUBS 0.007237f
C87 B.n36 VSUBS 0.007237f
C88 B.n37 VSUBS 0.007237f
C89 B.t10 VSUBS 0.264616f
C90 B.t11 VSUBS 0.286433f
C91 B.t9 VSUBS 0.945518f
C92 B.n38 VSUBS 0.423996f
C93 B.n39 VSUBS 0.283597f
C94 B.n40 VSUBS 0.007237f
C95 B.n41 VSUBS 0.007237f
C96 B.n42 VSUBS 0.007237f
C97 B.n43 VSUBS 0.007237f
C98 B.n44 VSUBS 0.004044f
C99 B.n45 VSUBS 0.007237f
C100 B.t7 VSUBS 0.26462f
C101 B.t8 VSUBS 0.286436f
C102 B.t6 VSUBS 0.945518f
C103 B.n46 VSUBS 0.423993f
C104 B.n47 VSUBS 0.283594f
C105 B.n48 VSUBS 0.016766f
C106 B.n49 VSUBS 0.007237f
C107 B.n50 VSUBS 0.007237f
C108 B.n51 VSUBS 0.007237f
C109 B.n52 VSUBS 0.007237f
C110 B.n53 VSUBS 0.007237f
C111 B.n54 VSUBS 0.007237f
C112 B.n55 VSUBS 0.007237f
C113 B.n56 VSUBS 0.007237f
C114 B.n57 VSUBS 0.007237f
C115 B.n58 VSUBS 0.007237f
C116 B.n59 VSUBS 0.007237f
C117 B.n60 VSUBS 0.007237f
C118 B.n61 VSUBS 0.007237f
C119 B.n62 VSUBS 0.007237f
C120 B.n63 VSUBS 0.007237f
C121 B.n64 VSUBS 0.007237f
C122 B.n65 VSUBS 0.007237f
C123 B.n66 VSUBS 0.007237f
C124 B.n67 VSUBS 0.007237f
C125 B.n68 VSUBS 0.007237f
C126 B.n69 VSUBS 0.007237f
C127 B.n70 VSUBS 0.007237f
C128 B.n71 VSUBS 0.017128f
C129 B.n72 VSUBS 0.007237f
C130 B.n73 VSUBS 0.007237f
C131 B.n74 VSUBS 0.007237f
C132 B.n75 VSUBS 0.007237f
C133 B.n76 VSUBS 0.007237f
C134 B.n77 VSUBS 0.007237f
C135 B.n78 VSUBS 0.007237f
C136 B.n79 VSUBS 0.007237f
C137 B.n80 VSUBS 0.007237f
C138 B.n81 VSUBS 0.007237f
C139 B.n82 VSUBS 0.007237f
C140 B.n83 VSUBS 0.007237f
C141 B.n84 VSUBS 0.007237f
C142 B.n85 VSUBS 0.007237f
C143 B.n86 VSUBS 0.007237f
C144 B.n87 VSUBS 0.007237f
C145 B.n88 VSUBS 0.007237f
C146 B.n89 VSUBS 0.007237f
C147 B.n90 VSUBS 0.007237f
C148 B.n91 VSUBS 0.007237f
C149 B.n92 VSUBS 0.007237f
C150 B.n93 VSUBS 0.007237f
C151 B.n94 VSUBS 0.007237f
C152 B.n95 VSUBS 0.007237f
C153 B.n96 VSUBS 0.017352f
C154 B.n97 VSUBS 0.007237f
C155 B.n98 VSUBS 0.007237f
C156 B.n99 VSUBS 0.007237f
C157 B.n100 VSUBS 0.007237f
C158 B.n101 VSUBS 0.007237f
C159 B.n102 VSUBS 0.007237f
C160 B.n103 VSUBS 0.007237f
C161 B.n104 VSUBS 0.007237f
C162 B.n105 VSUBS 0.007237f
C163 B.n106 VSUBS 0.007237f
C164 B.n107 VSUBS 0.007237f
C165 B.n108 VSUBS 0.007237f
C166 B.n109 VSUBS 0.007237f
C167 B.n110 VSUBS 0.007237f
C168 B.n111 VSUBS 0.007237f
C169 B.n112 VSUBS 0.007237f
C170 B.n113 VSUBS 0.007237f
C171 B.n114 VSUBS 0.007237f
C172 B.n115 VSUBS 0.007237f
C173 B.n116 VSUBS 0.007237f
C174 B.n117 VSUBS 0.007237f
C175 B.n118 VSUBS 0.007237f
C176 B.n119 VSUBS 0.006811f
C177 B.n120 VSUBS 0.007237f
C178 B.n121 VSUBS 0.007237f
C179 B.n122 VSUBS 0.007237f
C180 B.n123 VSUBS 0.007237f
C181 B.n124 VSUBS 0.007237f
C182 B.t5 VSUBS 0.264616f
C183 B.t4 VSUBS 0.286433f
C184 B.t3 VSUBS 0.945518f
C185 B.n125 VSUBS 0.423996f
C186 B.n126 VSUBS 0.283597f
C187 B.n127 VSUBS 0.007237f
C188 B.n128 VSUBS 0.007237f
C189 B.n129 VSUBS 0.007237f
C190 B.n130 VSUBS 0.007237f
C191 B.n131 VSUBS 0.007237f
C192 B.n132 VSUBS 0.007237f
C193 B.n133 VSUBS 0.007237f
C194 B.n134 VSUBS 0.007237f
C195 B.n135 VSUBS 0.007237f
C196 B.n136 VSUBS 0.007237f
C197 B.n137 VSUBS 0.007237f
C198 B.n138 VSUBS 0.007237f
C199 B.n139 VSUBS 0.007237f
C200 B.n140 VSUBS 0.007237f
C201 B.n141 VSUBS 0.007237f
C202 B.n142 VSUBS 0.007237f
C203 B.n143 VSUBS 0.007237f
C204 B.n144 VSUBS 0.007237f
C205 B.n145 VSUBS 0.007237f
C206 B.n146 VSUBS 0.007237f
C207 B.n147 VSUBS 0.007237f
C208 B.n148 VSUBS 0.007237f
C209 B.n149 VSUBS 0.007237f
C210 B.n150 VSUBS 0.017128f
C211 B.n151 VSUBS 0.007237f
C212 B.n152 VSUBS 0.007237f
C213 B.n153 VSUBS 0.007237f
C214 B.n154 VSUBS 0.007237f
C215 B.n155 VSUBS 0.007237f
C216 B.n156 VSUBS 0.007237f
C217 B.n157 VSUBS 0.007237f
C218 B.n158 VSUBS 0.007237f
C219 B.n159 VSUBS 0.007237f
C220 B.n160 VSUBS 0.007237f
C221 B.n161 VSUBS 0.007237f
C222 B.n162 VSUBS 0.007237f
C223 B.n163 VSUBS 0.007237f
C224 B.n164 VSUBS 0.007237f
C225 B.n165 VSUBS 0.007237f
C226 B.n166 VSUBS 0.007237f
C227 B.n167 VSUBS 0.007237f
C228 B.n168 VSUBS 0.007237f
C229 B.n169 VSUBS 0.007237f
C230 B.n170 VSUBS 0.007237f
C231 B.n171 VSUBS 0.007237f
C232 B.n172 VSUBS 0.007237f
C233 B.n173 VSUBS 0.007237f
C234 B.n174 VSUBS 0.007237f
C235 B.n175 VSUBS 0.007237f
C236 B.n176 VSUBS 0.007237f
C237 B.n177 VSUBS 0.007237f
C238 B.n178 VSUBS 0.007237f
C239 B.n179 VSUBS 0.007237f
C240 B.n180 VSUBS 0.007237f
C241 B.n181 VSUBS 0.007237f
C242 B.n182 VSUBS 0.007237f
C243 B.n183 VSUBS 0.007237f
C244 B.n184 VSUBS 0.007237f
C245 B.n185 VSUBS 0.007237f
C246 B.n186 VSUBS 0.007237f
C247 B.n187 VSUBS 0.007237f
C248 B.n188 VSUBS 0.007237f
C249 B.n189 VSUBS 0.007237f
C250 B.n190 VSUBS 0.007237f
C251 B.n191 VSUBS 0.007237f
C252 B.n192 VSUBS 0.007237f
C253 B.n193 VSUBS 0.007237f
C254 B.n194 VSUBS 0.007237f
C255 B.n195 VSUBS 0.017128f
C256 B.n196 VSUBS 0.017352f
C257 B.n197 VSUBS 0.017352f
C258 B.n198 VSUBS 0.007237f
C259 B.n199 VSUBS 0.007237f
C260 B.n200 VSUBS 0.007237f
C261 B.n201 VSUBS 0.007237f
C262 B.n202 VSUBS 0.007237f
C263 B.n203 VSUBS 0.007237f
C264 B.n204 VSUBS 0.007237f
C265 B.n205 VSUBS 0.007237f
C266 B.n206 VSUBS 0.007237f
C267 B.n207 VSUBS 0.007237f
C268 B.n208 VSUBS 0.007237f
C269 B.n209 VSUBS 0.007237f
C270 B.n210 VSUBS 0.007237f
C271 B.n211 VSUBS 0.007237f
C272 B.n212 VSUBS 0.007237f
C273 B.n213 VSUBS 0.007237f
C274 B.n214 VSUBS 0.007237f
C275 B.n215 VSUBS 0.007237f
C276 B.n216 VSUBS 0.007237f
C277 B.n217 VSUBS 0.007237f
C278 B.n218 VSUBS 0.007237f
C279 B.n219 VSUBS 0.007237f
C280 B.n220 VSUBS 0.007237f
C281 B.n221 VSUBS 0.007237f
C282 B.n222 VSUBS 0.007237f
C283 B.n223 VSUBS 0.007237f
C284 B.n224 VSUBS 0.007237f
C285 B.n225 VSUBS 0.007237f
C286 B.n226 VSUBS 0.007237f
C287 B.n227 VSUBS 0.007237f
C288 B.n228 VSUBS 0.007237f
C289 B.n229 VSUBS 0.007237f
C290 B.n230 VSUBS 0.007237f
C291 B.n231 VSUBS 0.007237f
C292 B.n232 VSUBS 0.007237f
C293 B.n233 VSUBS 0.007237f
C294 B.n234 VSUBS 0.007237f
C295 B.n235 VSUBS 0.007237f
C296 B.n236 VSUBS 0.007237f
C297 B.n237 VSUBS 0.007237f
C298 B.n238 VSUBS 0.007237f
C299 B.n239 VSUBS 0.007237f
C300 B.n240 VSUBS 0.007237f
C301 B.n241 VSUBS 0.007237f
C302 B.n242 VSUBS 0.007237f
C303 B.n243 VSUBS 0.007237f
C304 B.n244 VSUBS 0.007237f
C305 B.n245 VSUBS 0.007237f
C306 B.n246 VSUBS 0.007237f
C307 B.n247 VSUBS 0.007237f
C308 B.n248 VSUBS 0.007237f
C309 B.n249 VSUBS 0.007237f
C310 B.n250 VSUBS 0.007237f
C311 B.n251 VSUBS 0.007237f
C312 B.n252 VSUBS 0.007237f
C313 B.n253 VSUBS 0.007237f
C314 B.n254 VSUBS 0.007237f
C315 B.n255 VSUBS 0.007237f
C316 B.n256 VSUBS 0.007237f
C317 B.n257 VSUBS 0.007237f
C318 B.n258 VSUBS 0.007237f
C319 B.n259 VSUBS 0.007237f
C320 B.n260 VSUBS 0.007237f
C321 B.n261 VSUBS 0.007237f
C322 B.n262 VSUBS 0.007237f
C323 B.n263 VSUBS 0.007237f
C324 B.n264 VSUBS 0.007237f
C325 B.n265 VSUBS 0.007237f
C326 B.n266 VSUBS 0.006811f
C327 B.n267 VSUBS 0.016766f
C328 B.n268 VSUBS 0.004044f
C329 B.n269 VSUBS 0.007237f
C330 B.n270 VSUBS 0.007237f
C331 B.n271 VSUBS 0.007237f
C332 B.n272 VSUBS 0.007237f
C333 B.n273 VSUBS 0.007237f
C334 B.n274 VSUBS 0.007237f
C335 B.n275 VSUBS 0.007237f
C336 B.n276 VSUBS 0.007237f
C337 B.n277 VSUBS 0.007237f
C338 B.n278 VSUBS 0.007237f
C339 B.n279 VSUBS 0.007237f
C340 B.n280 VSUBS 0.007237f
C341 B.t2 VSUBS 0.26462f
C342 B.t1 VSUBS 0.286436f
C343 B.t0 VSUBS 0.945518f
C344 B.n281 VSUBS 0.423993f
C345 B.n282 VSUBS 0.283594f
C346 B.n283 VSUBS 0.016766f
C347 B.n284 VSUBS 0.004044f
C348 B.n285 VSUBS 0.007237f
C349 B.n286 VSUBS 0.007237f
C350 B.n287 VSUBS 0.007237f
C351 B.n288 VSUBS 0.007237f
C352 B.n289 VSUBS 0.007237f
C353 B.n290 VSUBS 0.007237f
C354 B.n291 VSUBS 0.007237f
C355 B.n292 VSUBS 0.007237f
C356 B.n293 VSUBS 0.007237f
C357 B.n294 VSUBS 0.007237f
C358 B.n295 VSUBS 0.007237f
C359 B.n296 VSUBS 0.007237f
C360 B.n297 VSUBS 0.007237f
C361 B.n298 VSUBS 0.007237f
C362 B.n299 VSUBS 0.007237f
C363 B.n300 VSUBS 0.007237f
C364 B.n301 VSUBS 0.007237f
C365 B.n302 VSUBS 0.007237f
C366 B.n303 VSUBS 0.007237f
C367 B.n304 VSUBS 0.007237f
C368 B.n305 VSUBS 0.007237f
C369 B.n306 VSUBS 0.007237f
C370 B.n307 VSUBS 0.007237f
C371 B.n308 VSUBS 0.007237f
C372 B.n309 VSUBS 0.007237f
C373 B.n310 VSUBS 0.007237f
C374 B.n311 VSUBS 0.007237f
C375 B.n312 VSUBS 0.007237f
C376 B.n313 VSUBS 0.007237f
C377 B.n314 VSUBS 0.007237f
C378 B.n315 VSUBS 0.007237f
C379 B.n316 VSUBS 0.007237f
C380 B.n317 VSUBS 0.007237f
C381 B.n318 VSUBS 0.007237f
C382 B.n319 VSUBS 0.007237f
C383 B.n320 VSUBS 0.007237f
C384 B.n321 VSUBS 0.007237f
C385 B.n322 VSUBS 0.007237f
C386 B.n323 VSUBS 0.007237f
C387 B.n324 VSUBS 0.007237f
C388 B.n325 VSUBS 0.007237f
C389 B.n326 VSUBS 0.007237f
C390 B.n327 VSUBS 0.007237f
C391 B.n328 VSUBS 0.007237f
C392 B.n329 VSUBS 0.007237f
C393 B.n330 VSUBS 0.007237f
C394 B.n331 VSUBS 0.007237f
C395 B.n332 VSUBS 0.007237f
C396 B.n333 VSUBS 0.007237f
C397 B.n334 VSUBS 0.007237f
C398 B.n335 VSUBS 0.007237f
C399 B.n336 VSUBS 0.007237f
C400 B.n337 VSUBS 0.007237f
C401 B.n338 VSUBS 0.007237f
C402 B.n339 VSUBS 0.007237f
C403 B.n340 VSUBS 0.007237f
C404 B.n341 VSUBS 0.007237f
C405 B.n342 VSUBS 0.007237f
C406 B.n343 VSUBS 0.007237f
C407 B.n344 VSUBS 0.007237f
C408 B.n345 VSUBS 0.007237f
C409 B.n346 VSUBS 0.007237f
C410 B.n347 VSUBS 0.007237f
C411 B.n348 VSUBS 0.007237f
C412 B.n349 VSUBS 0.007237f
C413 B.n350 VSUBS 0.007237f
C414 B.n351 VSUBS 0.007237f
C415 B.n352 VSUBS 0.007237f
C416 B.n353 VSUBS 0.007237f
C417 B.n354 VSUBS 0.007237f
C418 B.n355 VSUBS 0.01652f
C419 B.n356 VSUBS 0.017961f
C420 B.n357 VSUBS 0.017128f
C421 B.n358 VSUBS 0.007237f
C422 B.n359 VSUBS 0.007237f
C423 B.n360 VSUBS 0.007237f
C424 B.n361 VSUBS 0.007237f
C425 B.n362 VSUBS 0.007237f
C426 B.n363 VSUBS 0.007237f
C427 B.n364 VSUBS 0.007237f
C428 B.n365 VSUBS 0.007237f
C429 B.n366 VSUBS 0.007237f
C430 B.n367 VSUBS 0.007237f
C431 B.n368 VSUBS 0.007237f
C432 B.n369 VSUBS 0.007237f
C433 B.n370 VSUBS 0.007237f
C434 B.n371 VSUBS 0.007237f
C435 B.n372 VSUBS 0.007237f
C436 B.n373 VSUBS 0.007237f
C437 B.n374 VSUBS 0.007237f
C438 B.n375 VSUBS 0.007237f
C439 B.n376 VSUBS 0.007237f
C440 B.n377 VSUBS 0.007237f
C441 B.n378 VSUBS 0.007237f
C442 B.n379 VSUBS 0.007237f
C443 B.n380 VSUBS 0.007237f
C444 B.n381 VSUBS 0.007237f
C445 B.n382 VSUBS 0.007237f
C446 B.n383 VSUBS 0.007237f
C447 B.n384 VSUBS 0.007237f
C448 B.n385 VSUBS 0.007237f
C449 B.n386 VSUBS 0.007237f
C450 B.n387 VSUBS 0.007237f
C451 B.n388 VSUBS 0.007237f
C452 B.n389 VSUBS 0.007237f
C453 B.n390 VSUBS 0.007237f
C454 B.n391 VSUBS 0.007237f
C455 B.n392 VSUBS 0.007237f
C456 B.n393 VSUBS 0.007237f
C457 B.n394 VSUBS 0.007237f
C458 B.n395 VSUBS 0.007237f
C459 B.n396 VSUBS 0.007237f
C460 B.n397 VSUBS 0.007237f
C461 B.n398 VSUBS 0.007237f
C462 B.n399 VSUBS 0.007237f
C463 B.n400 VSUBS 0.007237f
C464 B.n401 VSUBS 0.007237f
C465 B.n402 VSUBS 0.007237f
C466 B.n403 VSUBS 0.007237f
C467 B.n404 VSUBS 0.007237f
C468 B.n405 VSUBS 0.007237f
C469 B.n406 VSUBS 0.007237f
C470 B.n407 VSUBS 0.007237f
C471 B.n408 VSUBS 0.007237f
C472 B.n409 VSUBS 0.007237f
C473 B.n410 VSUBS 0.007237f
C474 B.n411 VSUBS 0.007237f
C475 B.n412 VSUBS 0.007237f
C476 B.n413 VSUBS 0.007237f
C477 B.n414 VSUBS 0.007237f
C478 B.n415 VSUBS 0.007237f
C479 B.n416 VSUBS 0.007237f
C480 B.n417 VSUBS 0.007237f
C481 B.n418 VSUBS 0.007237f
C482 B.n419 VSUBS 0.007237f
C483 B.n420 VSUBS 0.007237f
C484 B.n421 VSUBS 0.007237f
C485 B.n422 VSUBS 0.007237f
C486 B.n423 VSUBS 0.007237f
C487 B.n424 VSUBS 0.007237f
C488 B.n425 VSUBS 0.007237f
C489 B.n426 VSUBS 0.007237f
C490 B.n427 VSUBS 0.007237f
C491 B.n428 VSUBS 0.007237f
C492 B.n429 VSUBS 0.007237f
C493 B.n430 VSUBS 0.017128f
C494 B.n431 VSUBS 0.017352f
C495 B.n432 VSUBS 0.017352f
C496 B.n433 VSUBS 0.007237f
C497 B.n434 VSUBS 0.007237f
C498 B.n435 VSUBS 0.007237f
C499 B.n436 VSUBS 0.007237f
C500 B.n437 VSUBS 0.007237f
C501 B.n438 VSUBS 0.007237f
C502 B.n439 VSUBS 0.007237f
C503 B.n440 VSUBS 0.007237f
C504 B.n441 VSUBS 0.007237f
C505 B.n442 VSUBS 0.007237f
C506 B.n443 VSUBS 0.007237f
C507 B.n444 VSUBS 0.007237f
C508 B.n445 VSUBS 0.007237f
C509 B.n446 VSUBS 0.007237f
C510 B.n447 VSUBS 0.007237f
C511 B.n448 VSUBS 0.007237f
C512 B.n449 VSUBS 0.007237f
C513 B.n450 VSUBS 0.007237f
C514 B.n451 VSUBS 0.007237f
C515 B.n452 VSUBS 0.007237f
C516 B.n453 VSUBS 0.007237f
C517 B.n454 VSUBS 0.007237f
C518 B.n455 VSUBS 0.007237f
C519 B.n456 VSUBS 0.007237f
C520 B.n457 VSUBS 0.007237f
C521 B.n458 VSUBS 0.007237f
C522 B.n459 VSUBS 0.007237f
C523 B.n460 VSUBS 0.007237f
C524 B.n461 VSUBS 0.007237f
C525 B.n462 VSUBS 0.007237f
C526 B.n463 VSUBS 0.007237f
C527 B.n464 VSUBS 0.007237f
C528 B.n465 VSUBS 0.007237f
C529 B.n466 VSUBS 0.007237f
C530 B.n467 VSUBS 0.007237f
C531 B.n468 VSUBS 0.007237f
C532 B.n469 VSUBS 0.007237f
C533 B.n470 VSUBS 0.007237f
C534 B.n471 VSUBS 0.007237f
C535 B.n472 VSUBS 0.007237f
C536 B.n473 VSUBS 0.007237f
C537 B.n474 VSUBS 0.007237f
C538 B.n475 VSUBS 0.007237f
C539 B.n476 VSUBS 0.007237f
C540 B.n477 VSUBS 0.007237f
C541 B.n478 VSUBS 0.007237f
C542 B.n479 VSUBS 0.007237f
C543 B.n480 VSUBS 0.007237f
C544 B.n481 VSUBS 0.007237f
C545 B.n482 VSUBS 0.007237f
C546 B.n483 VSUBS 0.007237f
C547 B.n484 VSUBS 0.007237f
C548 B.n485 VSUBS 0.007237f
C549 B.n486 VSUBS 0.007237f
C550 B.n487 VSUBS 0.007237f
C551 B.n488 VSUBS 0.007237f
C552 B.n489 VSUBS 0.007237f
C553 B.n490 VSUBS 0.007237f
C554 B.n491 VSUBS 0.007237f
C555 B.n492 VSUBS 0.007237f
C556 B.n493 VSUBS 0.007237f
C557 B.n494 VSUBS 0.007237f
C558 B.n495 VSUBS 0.007237f
C559 B.n496 VSUBS 0.007237f
C560 B.n497 VSUBS 0.007237f
C561 B.n498 VSUBS 0.007237f
C562 B.n499 VSUBS 0.007237f
C563 B.n500 VSUBS 0.006811f
C564 B.n501 VSUBS 0.007237f
C565 B.n502 VSUBS 0.007237f
C566 B.n503 VSUBS 0.007237f
C567 B.n504 VSUBS 0.007237f
C568 B.n505 VSUBS 0.007237f
C569 B.n506 VSUBS 0.007237f
C570 B.n507 VSUBS 0.007237f
C571 B.n508 VSUBS 0.007237f
C572 B.n509 VSUBS 0.007237f
C573 B.n510 VSUBS 0.007237f
C574 B.n511 VSUBS 0.007237f
C575 B.n512 VSUBS 0.007237f
C576 B.n513 VSUBS 0.007237f
C577 B.n514 VSUBS 0.007237f
C578 B.n515 VSUBS 0.007237f
C579 B.n516 VSUBS 0.004044f
C580 B.n517 VSUBS 0.016766f
C581 B.n518 VSUBS 0.006811f
C582 B.n519 VSUBS 0.007237f
C583 B.n520 VSUBS 0.007237f
C584 B.n521 VSUBS 0.007237f
C585 B.n522 VSUBS 0.007237f
C586 B.n523 VSUBS 0.007237f
C587 B.n524 VSUBS 0.007237f
C588 B.n525 VSUBS 0.007237f
C589 B.n526 VSUBS 0.007237f
C590 B.n527 VSUBS 0.007237f
C591 B.n528 VSUBS 0.007237f
C592 B.n529 VSUBS 0.007237f
C593 B.n530 VSUBS 0.007237f
C594 B.n531 VSUBS 0.007237f
C595 B.n532 VSUBS 0.007237f
C596 B.n533 VSUBS 0.007237f
C597 B.n534 VSUBS 0.007237f
C598 B.n535 VSUBS 0.007237f
C599 B.n536 VSUBS 0.007237f
C600 B.n537 VSUBS 0.007237f
C601 B.n538 VSUBS 0.007237f
C602 B.n539 VSUBS 0.007237f
C603 B.n540 VSUBS 0.007237f
C604 B.n541 VSUBS 0.007237f
C605 B.n542 VSUBS 0.007237f
C606 B.n543 VSUBS 0.007237f
C607 B.n544 VSUBS 0.007237f
C608 B.n545 VSUBS 0.007237f
C609 B.n546 VSUBS 0.007237f
C610 B.n547 VSUBS 0.007237f
C611 B.n548 VSUBS 0.007237f
C612 B.n549 VSUBS 0.007237f
C613 B.n550 VSUBS 0.007237f
C614 B.n551 VSUBS 0.007237f
C615 B.n552 VSUBS 0.007237f
C616 B.n553 VSUBS 0.007237f
C617 B.n554 VSUBS 0.007237f
C618 B.n555 VSUBS 0.007237f
C619 B.n556 VSUBS 0.007237f
C620 B.n557 VSUBS 0.007237f
C621 B.n558 VSUBS 0.007237f
C622 B.n559 VSUBS 0.007237f
C623 B.n560 VSUBS 0.007237f
C624 B.n561 VSUBS 0.007237f
C625 B.n562 VSUBS 0.007237f
C626 B.n563 VSUBS 0.007237f
C627 B.n564 VSUBS 0.007237f
C628 B.n565 VSUBS 0.007237f
C629 B.n566 VSUBS 0.007237f
C630 B.n567 VSUBS 0.007237f
C631 B.n568 VSUBS 0.007237f
C632 B.n569 VSUBS 0.007237f
C633 B.n570 VSUBS 0.007237f
C634 B.n571 VSUBS 0.007237f
C635 B.n572 VSUBS 0.007237f
C636 B.n573 VSUBS 0.007237f
C637 B.n574 VSUBS 0.007237f
C638 B.n575 VSUBS 0.007237f
C639 B.n576 VSUBS 0.007237f
C640 B.n577 VSUBS 0.007237f
C641 B.n578 VSUBS 0.007237f
C642 B.n579 VSUBS 0.007237f
C643 B.n580 VSUBS 0.007237f
C644 B.n581 VSUBS 0.007237f
C645 B.n582 VSUBS 0.007237f
C646 B.n583 VSUBS 0.007237f
C647 B.n584 VSUBS 0.007237f
C648 B.n585 VSUBS 0.007237f
C649 B.n586 VSUBS 0.007237f
C650 B.n587 VSUBS 0.017352f
C651 B.n588 VSUBS 0.017128f
C652 B.n589 VSUBS 0.017128f
C653 B.n590 VSUBS 0.007237f
C654 B.n591 VSUBS 0.007237f
C655 B.n592 VSUBS 0.007237f
C656 B.n593 VSUBS 0.007237f
C657 B.n594 VSUBS 0.007237f
C658 B.n595 VSUBS 0.007237f
C659 B.n596 VSUBS 0.007237f
C660 B.n597 VSUBS 0.007237f
C661 B.n598 VSUBS 0.007237f
C662 B.n599 VSUBS 0.007237f
C663 B.n600 VSUBS 0.007237f
C664 B.n601 VSUBS 0.007237f
C665 B.n602 VSUBS 0.007237f
C666 B.n603 VSUBS 0.007237f
C667 B.n604 VSUBS 0.007237f
C668 B.n605 VSUBS 0.007237f
C669 B.n606 VSUBS 0.007237f
C670 B.n607 VSUBS 0.007237f
C671 B.n608 VSUBS 0.007237f
C672 B.n609 VSUBS 0.007237f
C673 B.n610 VSUBS 0.007237f
C674 B.n611 VSUBS 0.007237f
C675 B.n612 VSUBS 0.007237f
C676 B.n613 VSUBS 0.007237f
C677 B.n614 VSUBS 0.007237f
C678 B.n615 VSUBS 0.007237f
C679 B.n616 VSUBS 0.007237f
C680 B.n617 VSUBS 0.007237f
C681 B.n618 VSUBS 0.007237f
C682 B.n619 VSUBS 0.007237f
C683 B.n620 VSUBS 0.007237f
C684 B.n621 VSUBS 0.007237f
C685 B.n622 VSUBS 0.007237f
C686 B.n623 VSUBS 0.009443f
C687 B.n624 VSUBS 0.01006f
C688 B.n625 VSUBS 0.020004f
C689 VDD2.t2 VSUBS 0.294715f
C690 VDD2.t3 VSUBS 0.294715f
C691 VDD2.n0 VSUBS 3.08946f
C692 VDD2.t0 VSUBS 0.294715f
C693 VDD2.t1 VSUBS 0.294715f
C694 VDD2.n1 VSUBS 2.37273f
C695 VDD2.n2 VSUBS 4.21697f
C696 VTAIL.n0 VSUBS 0.022999f
C697 VTAIL.n1 VSUBS 0.022492f
C698 VTAIL.n2 VSUBS 0.012441f
C699 VTAIL.n3 VSUBS 0.028567f
C700 VTAIL.n4 VSUBS 0.012797f
C701 VTAIL.n5 VSUBS 0.022492f
C702 VTAIL.n6 VSUBS 0.012086f
C703 VTAIL.n7 VSUBS 0.028567f
C704 VTAIL.n8 VSUBS 0.012797f
C705 VTAIL.n9 VSUBS 0.022492f
C706 VTAIL.n10 VSUBS 0.012086f
C707 VTAIL.n11 VSUBS 0.028567f
C708 VTAIL.n12 VSUBS 0.012797f
C709 VTAIL.n13 VSUBS 0.022492f
C710 VTAIL.n14 VSUBS 0.012086f
C711 VTAIL.n15 VSUBS 0.028567f
C712 VTAIL.n16 VSUBS 0.012797f
C713 VTAIL.n17 VSUBS 0.022492f
C714 VTAIL.n18 VSUBS 0.012086f
C715 VTAIL.n19 VSUBS 0.028567f
C716 VTAIL.n20 VSUBS 0.012797f
C717 VTAIL.n21 VSUBS 0.022492f
C718 VTAIL.n22 VSUBS 0.012086f
C719 VTAIL.n23 VSUBS 0.021425f
C720 VTAIL.n24 VSUBS 0.018173f
C721 VTAIL.t2 VSUBS 0.0611f
C722 VTAIL.n25 VSUBS 0.151846f
C723 VTAIL.n26 VSUBS 1.333f
C724 VTAIL.n27 VSUBS 0.012086f
C725 VTAIL.n28 VSUBS 0.012797f
C726 VTAIL.n29 VSUBS 0.028567f
C727 VTAIL.n30 VSUBS 0.028567f
C728 VTAIL.n31 VSUBS 0.012797f
C729 VTAIL.n32 VSUBS 0.012086f
C730 VTAIL.n33 VSUBS 0.022492f
C731 VTAIL.n34 VSUBS 0.022492f
C732 VTAIL.n35 VSUBS 0.012086f
C733 VTAIL.n36 VSUBS 0.012797f
C734 VTAIL.n37 VSUBS 0.028567f
C735 VTAIL.n38 VSUBS 0.028567f
C736 VTAIL.n39 VSUBS 0.012797f
C737 VTAIL.n40 VSUBS 0.012086f
C738 VTAIL.n41 VSUBS 0.022492f
C739 VTAIL.n42 VSUBS 0.022492f
C740 VTAIL.n43 VSUBS 0.012086f
C741 VTAIL.n44 VSUBS 0.012797f
C742 VTAIL.n45 VSUBS 0.028567f
C743 VTAIL.n46 VSUBS 0.028567f
C744 VTAIL.n47 VSUBS 0.012797f
C745 VTAIL.n48 VSUBS 0.012086f
C746 VTAIL.n49 VSUBS 0.022492f
C747 VTAIL.n50 VSUBS 0.022492f
C748 VTAIL.n51 VSUBS 0.012086f
C749 VTAIL.n52 VSUBS 0.012797f
C750 VTAIL.n53 VSUBS 0.028567f
C751 VTAIL.n54 VSUBS 0.028567f
C752 VTAIL.n55 VSUBS 0.012797f
C753 VTAIL.n56 VSUBS 0.012086f
C754 VTAIL.n57 VSUBS 0.022492f
C755 VTAIL.n58 VSUBS 0.022492f
C756 VTAIL.n59 VSUBS 0.012086f
C757 VTAIL.n60 VSUBS 0.012797f
C758 VTAIL.n61 VSUBS 0.028567f
C759 VTAIL.n62 VSUBS 0.028567f
C760 VTAIL.n63 VSUBS 0.012797f
C761 VTAIL.n64 VSUBS 0.012086f
C762 VTAIL.n65 VSUBS 0.022492f
C763 VTAIL.n66 VSUBS 0.022492f
C764 VTAIL.n67 VSUBS 0.012086f
C765 VTAIL.n68 VSUBS 0.012086f
C766 VTAIL.n69 VSUBS 0.012797f
C767 VTAIL.n70 VSUBS 0.028567f
C768 VTAIL.n71 VSUBS 0.028567f
C769 VTAIL.n72 VSUBS 0.063316f
C770 VTAIL.n73 VSUBS 0.012441f
C771 VTAIL.n74 VSUBS 0.012086f
C772 VTAIL.n75 VSUBS 0.054139f
C773 VTAIL.n76 VSUBS 0.031647f
C774 VTAIL.n77 VSUBS 0.11617f
C775 VTAIL.n78 VSUBS 0.022999f
C776 VTAIL.n79 VSUBS 0.022492f
C777 VTAIL.n80 VSUBS 0.012441f
C778 VTAIL.n81 VSUBS 0.028567f
C779 VTAIL.n82 VSUBS 0.012797f
C780 VTAIL.n83 VSUBS 0.022492f
C781 VTAIL.n84 VSUBS 0.012086f
C782 VTAIL.n85 VSUBS 0.028567f
C783 VTAIL.n86 VSUBS 0.012797f
C784 VTAIL.n87 VSUBS 0.022492f
C785 VTAIL.n88 VSUBS 0.012086f
C786 VTAIL.n89 VSUBS 0.028567f
C787 VTAIL.n90 VSUBS 0.012797f
C788 VTAIL.n91 VSUBS 0.022492f
C789 VTAIL.n92 VSUBS 0.012086f
C790 VTAIL.n93 VSUBS 0.028567f
C791 VTAIL.n94 VSUBS 0.012797f
C792 VTAIL.n95 VSUBS 0.022492f
C793 VTAIL.n96 VSUBS 0.012086f
C794 VTAIL.n97 VSUBS 0.028567f
C795 VTAIL.n98 VSUBS 0.012797f
C796 VTAIL.n99 VSUBS 0.022492f
C797 VTAIL.n100 VSUBS 0.012086f
C798 VTAIL.n101 VSUBS 0.021425f
C799 VTAIL.n102 VSUBS 0.018173f
C800 VTAIL.t1 VSUBS 0.0611f
C801 VTAIL.n103 VSUBS 0.151846f
C802 VTAIL.n104 VSUBS 1.333f
C803 VTAIL.n105 VSUBS 0.012086f
C804 VTAIL.n106 VSUBS 0.012797f
C805 VTAIL.n107 VSUBS 0.028567f
C806 VTAIL.n108 VSUBS 0.028567f
C807 VTAIL.n109 VSUBS 0.012797f
C808 VTAIL.n110 VSUBS 0.012086f
C809 VTAIL.n111 VSUBS 0.022492f
C810 VTAIL.n112 VSUBS 0.022492f
C811 VTAIL.n113 VSUBS 0.012086f
C812 VTAIL.n114 VSUBS 0.012797f
C813 VTAIL.n115 VSUBS 0.028567f
C814 VTAIL.n116 VSUBS 0.028567f
C815 VTAIL.n117 VSUBS 0.012797f
C816 VTAIL.n118 VSUBS 0.012086f
C817 VTAIL.n119 VSUBS 0.022492f
C818 VTAIL.n120 VSUBS 0.022492f
C819 VTAIL.n121 VSUBS 0.012086f
C820 VTAIL.n122 VSUBS 0.012797f
C821 VTAIL.n123 VSUBS 0.028567f
C822 VTAIL.n124 VSUBS 0.028567f
C823 VTAIL.n125 VSUBS 0.012797f
C824 VTAIL.n126 VSUBS 0.012086f
C825 VTAIL.n127 VSUBS 0.022492f
C826 VTAIL.n128 VSUBS 0.022492f
C827 VTAIL.n129 VSUBS 0.012086f
C828 VTAIL.n130 VSUBS 0.012797f
C829 VTAIL.n131 VSUBS 0.028567f
C830 VTAIL.n132 VSUBS 0.028567f
C831 VTAIL.n133 VSUBS 0.012797f
C832 VTAIL.n134 VSUBS 0.012086f
C833 VTAIL.n135 VSUBS 0.022492f
C834 VTAIL.n136 VSUBS 0.022492f
C835 VTAIL.n137 VSUBS 0.012086f
C836 VTAIL.n138 VSUBS 0.012797f
C837 VTAIL.n139 VSUBS 0.028567f
C838 VTAIL.n140 VSUBS 0.028567f
C839 VTAIL.n141 VSUBS 0.012797f
C840 VTAIL.n142 VSUBS 0.012086f
C841 VTAIL.n143 VSUBS 0.022492f
C842 VTAIL.n144 VSUBS 0.022492f
C843 VTAIL.n145 VSUBS 0.012086f
C844 VTAIL.n146 VSUBS 0.012086f
C845 VTAIL.n147 VSUBS 0.012797f
C846 VTAIL.n148 VSUBS 0.028567f
C847 VTAIL.n149 VSUBS 0.028567f
C848 VTAIL.n150 VSUBS 0.063316f
C849 VTAIL.n151 VSUBS 0.012441f
C850 VTAIL.n152 VSUBS 0.012086f
C851 VTAIL.n153 VSUBS 0.054139f
C852 VTAIL.n154 VSUBS 0.031647f
C853 VTAIL.n155 VSUBS 0.169431f
C854 VTAIL.n156 VSUBS 0.022999f
C855 VTAIL.n157 VSUBS 0.022492f
C856 VTAIL.n158 VSUBS 0.012441f
C857 VTAIL.n159 VSUBS 0.028567f
C858 VTAIL.n160 VSUBS 0.012797f
C859 VTAIL.n161 VSUBS 0.022492f
C860 VTAIL.n162 VSUBS 0.012086f
C861 VTAIL.n163 VSUBS 0.028567f
C862 VTAIL.n164 VSUBS 0.012797f
C863 VTAIL.n165 VSUBS 0.022492f
C864 VTAIL.n166 VSUBS 0.012086f
C865 VTAIL.n167 VSUBS 0.028567f
C866 VTAIL.n168 VSUBS 0.012797f
C867 VTAIL.n169 VSUBS 0.022492f
C868 VTAIL.n170 VSUBS 0.012086f
C869 VTAIL.n171 VSUBS 0.028567f
C870 VTAIL.n172 VSUBS 0.012797f
C871 VTAIL.n173 VSUBS 0.022492f
C872 VTAIL.n174 VSUBS 0.012086f
C873 VTAIL.n175 VSUBS 0.028567f
C874 VTAIL.n176 VSUBS 0.012797f
C875 VTAIL.n177 VSUBS 0.022492f
C876 VTAIL.n178 VSUBS 0.012086f
C877 VTAIL.n179 VSUBS 0.021425f
C878 VTAIL.n180 VSUBS 0.018173f
C879 VTAIL.t7 VSUBS 0.0611f
C880 VTAIL.n181 VSUBS 0.151846f
C881 VTAIL.n182 VSUBS 1.333f
C882 VTAIL.n183 VSUBS 0.012086f
C883 VTAIL.n184 VSUBS 0.012797f
C884 VTAIL.n185 VSUBS 0.028567f
C885 VTAIL.n186 VSUBS 0.028567f
C886 VTAIL.n187 VSUBS 0.012797f
C887 VTAIL.n188 VSUBS 0.012086f
C888 VTAIL.n189 VSUBS 0.022492f
C889 VTAIL.n190 VSUBS 0.022492f
C890 VTAIL.n191 VSUBS 0.012086f
C891 VTAIL.n192 VSUBS 0.012797f
C892 VTAIL.n193 VSUBS 0.028567f
C893 VTAIL.n194 VSUBS 0.028567f
C894 VTAIL.n195 VSUBS 0.012797f
C895 VTAIL.n196 VSUBS 0.012086f
C896 VTAIL.n197 VSUBS 0.022492f
C897 VTAIL.n198 VSUBS 0.022492f
C898 VTAIL.n199 VSUBS 0.012086f
C899 VTAIL.n200 VSUBS 0.012797f
C900 VTAIL.n201 VSUBS 0.028567f
C901 VTAIL.n202 VSUBS 0.028567f
C902 VTAIL.n203 VSUBS 0.012797f
C903 VTAIL.n204 VSUBS 0.012086f
C904 VTAIL.n205 VSUBS 0.022492f
C905 VTAIL.n206 VSUBS 0.022492f
C906 VTAIL.n207 VSUBS 0.012086f
C907 VTAIL.n208 VSUBS 0.012797f
C908 VTAIL.n209 VSUBS 0.028567f
C909 VTAIL.n210 VSUBS 0.028567f
C910 VTAIL.n211 VSUBS 0.012797f
C911 VTAIL.n212 VSUBS 0.012086f
C912 VTAIL.n213 VSUBS 0.022492f
C913 VTAIL.n214 VSUBS 0.022492f
C914 VTAIL.n215 VSUBS 0.012086f
C915 VTAIL.n216 VSUBS 0.012797f
C916 VTAIL.n217 VSUBS 0.028567f
C917 VTAIL.n218 VSUBS 0.028567f
C918 VTAIL.n219 VSUBS 0.012797f
C919 VTAIL.n220 VSUBS 0.012086f
C920 VTAIL.n221 VSUBS 0.022492f
C921 VTAIL.n222 VSUBS 0.022492f
C922 VTAIL.n223 VSUBS 0.012086f
C923 VTAIL.n224 VSUBS 0.012086f
C924 VTAIL.n225 VSUBS 0.012797f
C925 VTAIL.n226 VSUBS 0.028567f
C926 VTAIL.n227 VSUBS 0.028567f
C927 VTAIL.n228 VSUBS 0.063316f
C928 VTAIL.n229 VSUBS 0.012441f
C929 VTAIL.n230 VSUBS 0.012086f
C930 VTAIL.n231 VSUBS 0.054139f
C931 VTAIL.n232 VSUBS 0.031647f
C932 VTAIL.n233 VSUBS 1.42991f
C933 VTAIL.n234 VSUBS 0.022999f
C934 VTAIL.n235 VSUBS 0.022492f
C935 VTAIL.n236 VSUBS 0.012441f
C936 VTAIL.n237 VSUBS 0.028567f
C937 VTAIL.n238 VSUBS 0.012086f
C938 VTAIL.n239 VSUBS 0.012797f
C939 VTAIL.n240 VSUBS 0.022492f
C940 VTAIL.n241 VSUBS 0.012086f
C941 VTAIL.n242 VSUBS 0.028567f
C942 VTAIL.n243 VSUBS 0.012797f
C943 VTAIL.n244 VSUBS 0.022492f
C944 VTAIL.n245 VSUBS 0.012086f
C945 VTAIL.n246 VSUBS 0.028567f
C946 VTAIL.n247 VSUBS 0.012797f
C947 VTAIL.n248 VSUBS 0.022492f
C948 VTAIL.n249 VSUBS 0.012086f
C949 VTAIL.n250 VSUBS 0.028567f
C950 VTAIL.n251 VSUBS 0.012797f
C951 VTAIL.n252 VSUBS 0.022492f
C952 VTAIL.n253 VSUBS 0.012086f
C953 VTAIL.n254 VSUBS 0.028567f
C954 VTAIL.n255 VSUBS 0.012797f
C955 VTAIL.n256 VSUBS 0.022492f
C956 VTAIL.n257 VSUBS 0.012086f
C957 VTAIL.n258 VSUBS 0.021425f
C958 VTAIL.n259 VSUBS 0.018173f
C959 VTAIL.t5 VSUBS 0.0611f
C960 VTAIL.n260 VSUBS 0.151846f
C961 VTAIL.n261 VSUBS 1.333f
C962 VTAIL.n262 VSUBS 0.012086f
C963 VTAIL.n263 VSUBS 0.012797f
C964 VTAIL.n264 VSUBS 0.028567f
C965 VTAIL.n265 VSUBS 0.028567f
C966 VTAIL.n266 VSUBS 0.012797f
C967 VTAIL.n267 VSUBS 0.012086f
C968 VTAIL.n268 VSUBS 0.022492f
C969 VTAIL.n269 VSUBS 0.022492f
C970 VTAIL.n270 VSUBS 0.012086f
C971 VTAIL.n271 VSUBS 0.012797f
C972 VTAIL.n272 VSUBS 0.028567f
C973 VTAIL.n273 VSUBS 0.028567f
C974 VTAIL.n274 VSUBS 0.012797f
C975 VTAIL.n275 VSUBS 0.012086f
C976 VTAIL.n276 VSUBS 0.022492f
C977 VTAIL.n277 VSUBS 0.022492f
C978 VTAIL.n278 VSUBS 0.012086f
C979 VTAIL.n279 VSUBS 0.012797f
C980 VTAIL.n280 VSUBS 0.028567f
C981 VTAIL.n281 VSUBS 0.028567f
C982 VTAIL.n282 VSUBS 0.012797f
C983 VTAIL.n283 VSUBS 0.012086f
C984 VTAIL.n284 VSUBS 0.022492f
C985 VTAIL.n285 VSUBS 0.022492f
C986 VTAIL.n286 VSUBS 0.012086f
C987 VTAIL.n287 VSUBS 0.012797f
C988 VTAIL.n288 VSUBS 0.028567f
C989 VTAIL.n289 VSUBS 0.028567f
C990 VTAIL.n290 VSUBS 0.012797f
C991 VTAIL.n291 VSUBS 0.012086f
C992 VTAIL.n292 VSUBS 0.022492f
C993 VTAIL.n293 VSUBS 0.022492f
C994 VTAIL.n294 VSUBS 0.012086f
C995 VTAIL.n295 VSUBS 0.012797f
C996 VTAIL.n296 VSUBS 0.028567f
C997 VTAIL.n297 VSUBS 0.028567f
C998 VTAIL.n298 VSUBS 0.012797f
C999 VTAIL.n299 VSUBS 0.012086f
C1000 VTAIL.n300 VSUBS 0.022492f
C1001 VTAIL.n301 VSUBS 0.022492f
C1002 VTAIL.n302 VSUBS 0.012086f
C1003 VTAIL.n303 VSUBS 0.012797f
C1004 VTAIL.n304 VSUBS 0.028567f
C1005 VTAIL.n305 VSUBS 0.028567f
C1006 VTAIL.n306 VSUBS 0.063316f
C1007 VTAIL.n307 VSUBS 0.012441f
C1008 VTAIL.n308 VSUBS 0.012086f
C1009 VTAIL.n309 VSUBS 0.054139f
C1010 VTAIL.n310 VSUBS 0.031647f
C1011 VTAIL.n311 VSUBS 1.42991f
C1012 VTAIL.n312 VSUBS 0.022999f
C1013 VTAIL.n313 VSUBS 0.022492f
C1014 VTAIL.n314 VSUBS 0.012441f
C1015 VTAIL.n315 VSUBS 0.028567f
C1016 VTAIL.n316 VSUBS 0.012086f
C1017 VTAIL.n317 VSUBS 0.012797f
C1018 VTAIL.n318 VSUBS 0.022492f
C1019 VTAIL.n319 VSUBS 0.012086f
C1020 VTAIL.n320 VSUBS 0.028567f
C1021 VTAIL.n321 VSUBS 0.012797f
C1022 VTAIL.n322 VSUBS 0.022492f
C1023 VTAIL.n323 VSUBS 0.012086f
C1024 VTAIL.n324 VSUBS 0.028567f
C1025 VTAIL.n325 VSUBS 0.012797f
C1026 VTAIL.n326 VSUBS 0.022492f
C1027 VTAIL.n327 VSUBS 0.012086f
C1028 VTAIL.n328 VSUBS 0.028567f
C1029 VTAIL.n329 VSUBS 0.012797f
C1030 VTAIL.n330 VSUBS 0.022492f
C1031 VTAIL.n331 VSUBS 0.012086f
C1032 VTAIL.n332 VSUBS 0.028567f
C1033 VTAIL.n333 VSUBS 0.012797f
C1034 VTAIL.n334 VSUBS 0.022492f
C1035 VTAIL.n335 VSUBS 0.012086f
C1036 VTAIL.n336 VSUBS 0.021425f
C1037 VTAIL.n337 VSUBS 0.018173f
C1038 VTAIL.t4 VSUBS 0.0611f
C1039 VTAIL.n338 VSUBS 0.151846f
C1040 VTAIL.n339 VSUBS 1.333f
C1041 VTAIL.n340 VSUBS 0.012086f
C1042 VTAIL.n341 VSUBS 0.012797f
C1043 VTAIL.n342 VSUBS 0.028567f
C1044 VTAIL.n343 VSUBS 0.028567f
C1045 VTAIL.n344 VSUBS 0.012797f
C1046 VTAIL.n345 VSUBS 0.012086f
C1047 VTAIL.n346 VSUBS 0.022492f
C1048 VTAIL.n347 VSUBS 0.022492f
C1049 VTAIL.n348 VSUBS 0.012086f
C1050 VTAIL.n349 VSUBS 0.012797f
C1051 VTAIL.n350 VSUBS 0.028567f
C1052 VTAIL.n351 VSUBS 0.028567f
C1053 VTAIL.n352 VSUBS 0.012797f
C1054 VTAIL.n353 VSUBS 0.012086f
C1055 VTAIL.n354 VSUBS 0.022492f
C1056 VTAIL.n355 VSUBS 0.022492f
C1057 VTAIL.n356 VSUBS 0.012086f
C1058 VTAIL.n357 VSUBS 0.012797f
C1059 VTAIL.n358 VSUBS 0.028567f
C1060 VTAIL.n359 VSUBS 0.028567f
C1061 VTAIL.n360 VSUBS 0.012797f
C1062 VTAIL.n361 VSUBS 0.012086f
C1063 VTAIL.n362 VSUBS 0.022492f
C1064 VTAIL.n363 VSUBS 0.022492f
C1065 VTAIL.n364 VSUBS 0.012086f
C1066 VTAIL.n365 VSUBS 0.012797f
C1067 VTAIL.n366 VSUBS 0.028567f
C1068 VTAIL.n367 VSUBS 0.028567f
C1069 VTAIL.n368 VSUBS 0.012797f
C1070 VTAIL.n369 VSUBS 0.012086f
C1071 VTAIL.n370 VSUBS 0.022492f
C1072 VTAIL.n371 VSUBS 0.022492f
C1073 VTAIL.n372 VSUBS 0.012086f
C1074 VTAIL.n373 VSUBS 0.012797f
C1075 VTAIL.n374 VSUBS 0.028567f
C1076 VTAIL.n375 VSUBS 0.028567f
C1077 VTAIL.n376 VSUBS 0.012797f
C1078 VTAIL.n377 VSUBS 0.012086f
C1079 VTAIL.n378 VSUBS 0.022492f
C1080 VTAIL.n379 VSUBS 0.022492f
C1081 VTAIL.n380 VSUBS 0.012086f
C1082 VTAIL.n381 VSUBS 0.012797f
C1083 VTAIL.n382 VSUBS 0.028567f
C1084 VTAIL.n383 VSUBS 0.028567f
C1085 VTAIL.n384 VSUBS 0.063316f
C1086 VTAIL.n385 VSUBS 0.012441f
C1087 VTAIL.n386 VSUBS 0.012086f
C1088 VTAIL.n387 VSUBS 0.054139f
C1089 VTAIL.n388 VSUBS 0.031647f
C1090 VTAIL.n389 VSUBS 0.169431f
C1091 VTAIL.n390 VSUBS 0.022999f
C1092 VTAIL.n391 VSUBS 0.022492f
C1093 VTAIL.n392 VSUBS 0.012441f
C1094 VTAIL.n393 VSUBS 0.028567f
C1095 VTAIL.n394 VSUBS 0.012086f
C1096 VTAIL.n395 VSUBS 0.012797f
C1097 VTAIL.n396 VSUBS 0.022492f
C1098 VTAIL.n397 VSUBS 0.012086f
C1099 VTAIL.n398 VSUBS 0.028567f
C1100 VTAIL.n399 VSUBS 0.012797f
C1101 VTAIL.n400 VSUBS 0.022492f
C1102 VTAIL.n401 VSUBS 0.012086f
C1103 VTAIL.n402 VSUBS 0.028567f
C1104 VTAIL.n403 VSUBS 0.012797f
C1105 VTAIL.n404 VSUBS 0.022492f
C1106 VTAIL.n405 VSUBS 0.012086f
C1107 VTAIL.n406 VSUBS 0.028567f
C1108 VTAIL.n407 VSUBS 0.012797f
C1109 VTAIL.n408 VSUBS 0.022492f
C1110 VTAIL.n409 VSUBS 0.012086f
C1111 VTAIL.n410 VSUBS 0.028567f
C1112 VTAIL.n411 VSUBS 0.012797f
C1113 VTAIL.n412 VSUBS 0.022492f
C1114 VTAIL.n413 VSUBS 0.012086f
C1115 VTAIL.n414 VSUBS 0.021425f
C1116 VTAIL.n415 VSUBS 0.018173f
C1117 VTAIL.t6 VSUBS 0.0611f
C1118 VTAIL.n416 VSUBS 0.151846f
C1119 VTAIL.n417 VSUBS 1.333f
C1120 VTAIL.n418 VSUBS 0.012086f
C1121 VTAIL.n419 VSUBS 0.012797f
C1122 VTAIL.n420 VSUBS 0.028567f
C1123 VTAIL.n421 VSUBS 0.028567f
C1124 VTAIL.n422 VSUBS 0.012797f
C1125 VTAIL.n423 VSUBS 0.012086f
C1126 VTAIL.n424 VSUBS 0.022492f
C1127 VTAIL.n425 VSUBS 0.022492f
C1128 VTAIL.n426 VSUBS 0.012086f
C1129 VTAIL.n427 VSUBS 0.012797f
C1130 VTAIL.n428 VSUBS 0.028567f
C1131 VTAIL.n429 VSUBS 0.028567f
C1132 VTAIL.n430 VSUBS 0.012797f
C1133 VTAIL.n431 VSUBS 0.012086f
C1134 VTAIL.n432 VSUBS 0.022492f
C1135 VTAIL.n433 VSUBS 0.022492f
C1136 VTAIL.n434 VSUBS 0.012086f
C1137 VTAIL.n435 VSUBS 0.012797f
C1138 VTAIL.n436 VSUBS 0.028567f
C1139 VTAIL.n437 VSUBS 0.028567f
C1140 VTAIL.n438 VSUBS 0.012797f
C1141 VTAIL.n439 VSUBS 0.012086f
C1142 VTAIL.n440 VSUBS 0.022492f
C1143 VTAIL.n441 VSUBS 0.022492f
C1144 VTAIL.n442 VSUBS 0.012086f
C1145 VTAIL.n443 VSUBS 0.012797f
C1146 VTAIL.n444 VSUBS 0.028567f
C1147 VTAIL.n445 VSUBS 0.028567f
C1148 VTAIL.n446 VSUBS 0.012797f
C1149 VTAIL.n447 VSUBS 0.012086f
C1150 VTAIL.n448 VSUBS 0.022492f
C1151 VTAIL.n449 VSUBS 0.022492f
C1152 VTAIL.n450 VSUBS 0.012086f
C1153 VTAIL.n451 VSUBS 0.012797f
C1154 VTAIL.n452 VSUBS 0.028567f
C1155 VTAIL.n453 VSUBS 0.028567f
C1156 VTAIL.n454 VSUBS 0.012797f
C1157 VTAIL.n455 VSUBS 0.012086f
C1158 VTAIL.n456 VSUBS 0.022492f
C1159 VTAIL.n457 VSUBS 0.022492f
C1160 VTAIL.n458 VSUBS 0.012086f
C1161 VTAIL.n459 VSUBS 0.012797f
C1162 VTAIL.n460 VSUBS 0.028567f
C1163 VTAIL.n461 VSUBS 0.028567f
C1164 VTAIL.n462 VSUBS 0.063316f
C1165 VTAIL.n463 VSUBS 0.012441f
C1166 VTAIL.n464 VSUBS 0.012086f
C1167 VTAIL.n465 VSUBS 0.054139f
C1168 VTAIL.n466 VSUBS 0.031647f
C1169 VTAIL.n467 VSUBS 0.169431f
C1170 VTAIL.n468 VSUBS 0.022999f
C1171 VTAIL.n469 VSUBS 0.022492f
C1172 VTAIL.n470 VSUBS 0.012441f
C1173 VTAIL.n471 VSUBS 0.028567f
C1174 VTAIL.n472 VSUBS 0.012086f
C1175 VTAIL.n473 VSUBS 0.012797f
C1176 VTAIL.n474 VSUBS 0.022492f
C1177 VTAIL.n475 VSUBS 0.012086f
C1178 VTAIL.n476 VSUBS 0.028567f
C1179 VTAIL.n477 VSUBS 0.012797f
C1180 VTAIL.n478 VSUBS 0.022492f
C1181 VTAIL.n479 VSUBS 0.012086f
C1182 VTAIL.n480 VSUBS 0.028567f
C1183 VTAIL.n481 VSUBS 0.012797f
C1184 VTAIL.n482 VSUBS 0.022492f
C1185 VTAIL.n483 VSUBS 0.012086f
C1186 VTAIL.n484 VSUBS 0.028567f
C1187 VTAIL.n485 VSUBS 0.012797f
C1188 VTAIL.n486 VSUBS 0.022492f
C1189 VTAIL.n487 VSUBS 0.012086f
C1190 VTAIL.n488 VSUBS 0.028567f
C1191 VTAIL.n489 VSUBS 0.012797f
C1192 VTAIL.n490 VSUBS 0.022492f
C1193 VTAIL.n491 VSUBS 0.012086f
C1194 VTAIL.n492 VSUBS 0.021425f
C1195 VTAIL.n493 VSUBS 0.018173f
C1196 VTAIL.t0 VSUBS 0.0611f
C1197 VTAIL.n494 VSUBS 0.151846f
C1198 VTAIL.n495 VSUBS 1.333f
C1199 VTAIL.n496 VSUBS 0.012086f
C1200 VTAIL.n497 VSUBS 0.012797f
C1201 VTAIL.n498 VSUBS 0.028567f
C1202 VTAIL.n499 VSUBS 0.028567f
C1203 VTAIL.n500 VSUBS 0.012797f
C1204 VTAIL.n501 VSUBS 0.012086f
C1205 VTAIL.n502 VSUBS 0.022492f
C1206 VTAIL.n503 VSUBS 0.022492f
C1207 VTAIL.n504 VSUBS 0.012086f
C1208 VTAIL.n505 VSUBS 0.012797f
C1209 VTAIL.n506 VSUBS 0.028567f
C1210 VTAIL.n507 VSUBS 0.028567f
C1211 VTAIL.n508 VSUBS 0.012797f
C1212 VTAIL.n509 VSUBS 0.012086f
C1213 VTAIL.n510 VSUBS 0.022492f
C1214 VTAIL.n511 VSUBS 0.022492f
C1215 VTAIL.n512 VSUBS 0.012086f
C1216 VTAIL.n513 VSUBS 0.012797f
C1217 VTAIL.n514 VSUBS 0.028567f
C1218 VTAIL.n515 VSUBS 0.028567f
C1219 VTAIL.n516 VSUBS 0.012797f
C1220 VTAIL.n517 VSUBS 0.012086f
C1221 VTAIL.n518 VSUBS 0.022492f
C1222 VTAIL.n519 VSUBS 0.022492f
C1223 VTAIL.n520 VSUBS 0.012086f
C1224 VTAIL.n521 VSUBS 0.012797f
C1225 VTAIL.n522 VSUBS 0.028567f
C1226 VTAIL.n523 VSUBS 0.028567f
C1227 VTAIL.n524 VSUBS 0.012797f
C1228 VTAIL.n525 VSUBS 0.012086f
C1229 VTAIL.n526 VSUBS 0.022492f
C1230 VTAIL.n527 VSUBS 0.022492f
C1231 VTAIL.n528 VSUBS 0.012086f
C1232 VTAIL.n529 VSUBS 0.012797f
C1233 VTAIL.n530 VSUBS 0.028567f
C1234 VTAIL.n531 VSUBS 0.028567f
C1235 VTAIL.n532 VSUBS 0.012797f
C1236 VTAIL.n533 VSUBS 0.012086f
C1237 VTAIL.n534 VSUBS 0.022492f
C1238 VTAIL.n535 VSUBS 0.022492f
C1239 VTAIL.n536 VSUBS 0.012086f
C1240 VTAIL.n537 VSUBS 0.012797f
C1241 VTAIL.n538 VSUBS 0.028567f
C1242 VTAIL.n539 VSUBS 0.028567f
C1243 VTAIL.n540 VSUBS 0.063316f
C1244 VTAIL.n541 VSUBS 0.012441f
C1245 VTAIL.n542 VSUBS 0.012086f
C1246 VTAIL.n543 VSUBS 0.054139f
C1247 VTAIL.n544 VSUBS 0.031647f
C1248 VTAIL.n545 VSUBS 1.42991f
C1249 VTAIL.n546 VSUBS 0.022999f
C1250 VTAIL.n547 VSUBS 0.022492f
C1251 VTAIL.n548 VSUBS 0.012441f
C1252 VTAIL.n549 VSUBS 0.028567f
C1253 VTAIL.n550 VSUBS 0.012797f
C1254 VTAIL.n551 VSUBS 0.022492f
C1255 VTAIL.n552 VSUBS 0.012086f
C1256 VTAIL.n553 VSUBS 0.028567f
C1257 VTAIL.n554 VSUBS 0.012797f
C1258 VTAIL.n555 VSUBS 0.022492f
C1259 VTAIL.n556 VSUBS 0.012086f
C1260 VTAIL.n557 VSUBS 0.028567f
C1261 VTAIL.n558 VSUBS 0.012797f
C1262 VTAIL.n559 VSUBS 0.022492f
C1263 VTAIL.n560 VSUBS 0.012086f
C1264 VTAIL.n561 VSUBS 0.028567f
C1265 VTAIL.n562 VSUBS 0.012797f
C1266 VTAIL.n563 VSUBS 0.022492f
C1267 VTAIL.n564 VSUBS 0.012086f
C1268 VTAIL.n565 VSUBS 0.028567f
C1269 VTAIL.n566 VSUBS 0.012797f
C1270 VTAIL.n567 VSUBS 0.022492f
C1271 VTAIL.n568 VSUBS 0.012086f
C1272 VTAIL.n569 VSUBS 0.021425f
C1273 VTAIL.n570 VSUBS 0.018173f
C1274 VTAIL.t3 VSUBS 0.0611f
C1275 VTAIL.n571 VSUBS 0.151846f
C1276 VTAIL.n572 VSUBS 1.333f
C1277 VTAIL.n573 VSUBS 0.012086f
C1278 VTAIL.n574 VSUBS 0.012797f
C1279 VTAIL.n575 VSUBS 0.028567f
C1280 VTAIL.n576 VSUBS 0.028567f
C1281 VTAIL.n577 VSUBS 0.012797f
C1282 VTAIL.n578 VSUBS 0.012086f
C1283 VTAIL.n579 VSUBS 0.022492f
C1284 VTAIL.n580 VSUBS 0.022492f
C1285 VTAIL.n581 VSUBS 0.012086f
C1286 VTAIL.n582 VSUBS 0.012797f
C1287 VTAIL.n583 VSUBS 0.028567f
C1288 VTAIL.n584 VSUBS 0.028567f
C1289 VTAIL.n585 VSUBS 0.012797f
C1290 VTAIL.n586 VSUBS 0.012086f
C1291 VTAIL.n587 VSUBS 0.022492f
C1292 VTAIL.n588 VSUBS 0.022492f
C1293 VTAIL.n589 VSUBS 0.012086f
C1294 VTAIL.n590 VSUBS 0.012797f
C1295 VTAIL.n591 VSUBS 0.028567f
C1296 VTAIL.n592 VSUBS 0.028567f
C1297 VTAIL.n593 VSUBS 0.012797f
C1298 VTAIL.n594 VSUBS 0.012086f
C1299 VTAIL.n595 VSUBS 0.022492f
C1300 VTAIL.n596 VSUBS 0.022492f
C1301 VTAIL.n597 VSUBS 0.012086f
C1302 VTAIL.n598 VSUBS 0.012797f
C1303 VTAIL.n599 VSUBS 0.028567f
C1304 VTAIL.n600 VSUBS 0.028567f
C1305 VTAIL.n601 VSUBS 0.012797f
C1306 VTAIL.n602 VSUBS 0.012086f
C1307 VTAIL.n603 VSUBS 0.022492f
C1308 VTAIL.n604 VSUBS 0.022492f
C1309 VTAIL.n605 VSUBS 0.012086f
C1310 VTAIL.n606 VSUBS 0.012797f
C1311 VTAIL.n607 VSUBS 0.028567f
C1312 VTAIL.n608 VSUBS 0.028567f
C1313 VTAIL.n609 VSUBS 0.012797f
C1314 VTAIL.n610 VSUBS 0.012086f
C1315 VTAIL.n611 VSUBS 0.022492f
C1316 VTAIL.n612 VSUBS 0.022492f
C1317 VTAIL.n613 VSUBS 0.012086f
C1318 VTAIL.n614 VSUBS 0.012086f
C1319 VTAIL.n615 VSUBS 0.012797f
C1320 VTAIL.n616 VSUBS 0.028567f
C1321 VTAIL.n617 VSUBS 0.028567f
C1322 VTAIL.n618 VSUBS 0.063316f
C1323 VTAIL.n619 VSUBS 0.012441f
C1324 VTAIL.n620 VSUBS 0.012086f
C1325 VTAIL.n621 VSUBS 0.054139f
C1326 VTAIL.n622 VSUBS 0.031647f
C1327 VTAIL.n623 VSUBS 1.36821f
C1328 VN.t1 VSUBS 2.58214f
C1329 VN.t0 VSUBS 2.58083f
C1330 VN.n0 VSUBS 1.85258f
C1331 VN.t2 VSUBS 2.58214f
C1332 VN.t3 VSUBS 2.58083f
C1333 VN.n1 VSUBS 3.53131f
.ends

