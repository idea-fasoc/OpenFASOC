* NGSPICE file created from diff_pair_sample_0523.ext - technology: sky130A

.subckt diff_pair_sample_0523 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=1.1484 ps=7.29 w=6.96 l=2.59
X1 VDD2.t1 VN.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=1.1484 ps=7.29 w=6.96 l=2.59
X2 VDD1.t5 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=1.1484 ps=7.29 w=6.96 l=2.59
X3 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=2.59
X4 VDD2.t3 VN.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=2.7144 ps=14.7 w=6.96 l=2.59
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=2.59
X6 VTAIL.t4 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=1.1484 ps=7.29 w=6.96 l=2.59
X7 VDD2.t5 VN.t3 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=1.1484 ps=7.29 w=6.96 l=2.59
X8 VTAIL.t7 VN.t4 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=1.1484 ps=7.29 w=6.96 l=2.59
X9 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=2.59
X10 VDD2.t0 VN.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=2.7144 ps=14.7 w=6.96 l=2.59
X11 VTAIL.t5 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=1.1484 ps=7.29 w=6.96 l=2.59
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=0 ps=0 w=6.96 l=2.59
X13 VDD1.t2 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=2.7144 ps=14.7 w=6.96 l=2.59
X14 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7144 pd=14.7 as=1.1484 ps=7.29 w=6.96 l=2.59
X15 VDD1.t0 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1484 pd=7.29 as=2.7144 ps=14.7 w=6.96 l=2.59
R0 VN.n29 VN.n16 161.3
R1 VN.n28 VN.n27 161.3
R2 VN.n26 VN.n17 161.3
R3 VN.n25 VN.n24 161.3
R4 VN.n23 VN.n18 161.3
R5 VN.n22 VN.n21 161.3
R6 VN.n13 VN.n0 161.3
R7 VN.n12 VN.n11 161.3
R8 VN.n10 VN.n1 161.3
R9 VN.n9 VN.n8 161.3
R10 VN.n7 VN.n2 161.3
R11 VN.n6 VN.n5 161.3
R12 VN.n15 VN.n14 102.547
R13 VN.n31 VN.n30 102.547
R14 VN.n4 VN.t1 97.9633
R15 VN.n20 VN.t5 97.9633
R16 VN.n3 VN.t4 64.7634
R17 VN.n14 VN.t2 64.7634
R18 VN.n19 VN.t0 64.7634
R19 VN.n30 VN.t3 64.7634
R20 VN.n4 VN.n3 60.2807
R21 VN.n20 VN.n19 60.2807
R22 VN.n8 VN.n1 56.5617
R23 VN.n24 VN.n17 56.5617
R24 VN VN.n31 45.0891
R25 VN.n7 VN.n6 24.5923
R26 VN.n8 VN.n7 24.5923
R27 VN.n12 VN.n1 24.5923
R28 VN.n13 VN.n12 24.5923
R29 VN.n24 VN.n23 24.5923
R30 VN.n23 VN.n22 24.5923
R31 VN.n29 VN.n28 24.5923
R32 VN.n28 VN.n17 24.5923
R33 VN.n6 VN.n3 12.2964
R34 VN.n22 VN.n19 12.2964
R35 VN.n14 VN.n13 8.36172
R36 VN.n30 VN.n29 8.36172
R37 VN.n21 VN.n20 6.93618
R38 VN.n5 VN.n4 6.93618
R39 VN.n31 VN.n16 0.278335
R40 VN.n15 VN.n0 0.278335
R41 VN.n27 VN.n16 0.189894
R42 VN.n27 VN.n26 0.189894
R43 VN.n26 VN.n25 0.189894
R44 VN.n25 VN.n18 0.189894
R45 VN.n21 VN.n18 0.189894
R46 VN.n5 VN.n2 0.189894
R47 VN.n9 VN.n2 0.189894
R48 VN.n10 VN.n9 0.189894
R49 VN.n11 VN.n10 0.189894
R50 VN.n11 VN.n0 0.189894
R51 VN VN.n15 0.153485
R52 VDD2.n1 VDD2.t1 67.9612
R53 VDD2.n2 VDD2.t5 66.1288
R54 VDD2.n1 VDD2.n0 63.8579
R55 VDD2 VDD2.n3 63.8549
R56 VDD2.n2 VDD2.n1 37.8963
R57 VDD2.n3 VDD2.t2 2.84533
R58 VDD2.n3 VDD2.t0 2.84533
R59 VDD2.n0 VDD2.t4 2.84533
R60 VDD2.n0 VDD2.t3 2.84533
R61 VDD2 VDD2.n2 1.94662
R62 VTAIL.n7 VTAIL.t6 49.45
R63 VTAIL.n11 VTAIL.t9 49.4498
R64 VTAIL.n2 VTAIL.t0 49.4498
R65 VTAIL.n10 VTAIL.t2 49.4498
R66 VTAIL.n9 VTAIL.n8 46.6052
R67 VTAIL.n6 VTAIL.n5 46.6052
R68 VTAIL.n1 VTAIL.n0 46.6051
R69 VTAIL.n4 VTAIL.n3 46.6051
R70 VTAIL.n6 VTAIL.n4 23.4014
R71 VTAIL.n11 VTAIL.n10 20.8841
R72 VTAIL.n0 VTAIL.t10 2.84533
R73 VTAIL.n0 VTAIL.t7 2.84533
R74 VTAIL.n3 VTAIL.t1 2.84533
R75 VTAIL.n3 VTAIL.t5 2.84533
R76 VTAIL.n8 VTAIL.t3 2.84533
R77 VTAIL.n8 VTAIL.t4 2.84533
R78 VTAIL.n5 VTAIL.t8 2.84533
R79 VTAIL.n5 VTAIL.t11 2.84533
R80 VTAIL.n7 VTAIL.n6 2.51774
R81 VTAIL.n10 VTAIL.n9 2.51774
R82 VTAIL.n4 VTAIL.n2 2.51774
R83 VTAIL VTAIL.n11 1.83024
R84 VTAIL.n9 VTAIL.n7 1.72895
R85 VTAIL.n2 VTAIL.n1 1.72895
R86 VTAIL VTAIL.n1 0.688
R87 B.n543 B.n542 585
R88 B.n543 B.n79 585
R89 B.n546 B.n545 585
R90 B.n547 B.n115 585
R91 B.n549 B.n548 585
R92 B.n551 B.n114 585
R93 B.n554 B.n553 585
R94 B.n555 B.n113 585
R95 B.n557 B.n556 585
R96 B.n559 B.n112 585
R97 B.n562 B.n561 585
R98 B.n563 B.n111 585
R99 B.n565 B.n564 585
R100 B.n567 B.n110 585
R101 B.n570 B.n569 585
R102 B.n571 B.n109 585
R103 B.n573 B.n572 585
R104 B.n575 B.n108 585
R105 B.n578 B.n577 585
R106 B.n579 B.n107 585
R107 B.n581 B.n580 585
R108 B.n583 B.n106 585
R109 B.n586 B.n585 585
R110 B.n587 B.n105 585
R111 B.n589 B.n588 585
R112 B.n591 B.n104 585
R113 B.n594 B.n593 585
R114 B.n595 B.n101 585
R115 B.n598 B.n597 585
R116 B.n600 B.n100 585
R117 B.n603 B.n602 585
R118 B.n604 B.n99 585
R119 B.n606 B.n605 585
R120 B.n608 B.n98 585
R121 B.n611 B.n610 585
R122 B.n612 B.n94 585
R123 B.n614 B.n613 585
R124 B.n616 B.n93 585
R125 B.n619 B.n618 585
R126 B.n620 B.n92 585
R127 B.n622 B.n621 585
R128 B.n624 B.n91 585
R129 B.n627 B.n626 585
R130 B.n628 B.n90 585
R131 B.n630 B.n629 585
R132 B.n632 B.n89 585
R133 B.n635 B.n634 585
R134 B.n636 B.n88 585
R135 B.n638 B.n637 585
R136 B.n640 B.n87 585
R137 B.n643 B.n642 585
R138 B.n644 B.n86 585
R139 B.n646 B.n645 585
R140 B.n648 B.n85 585
R141 B.n651 B.n650 585
R142 B.n652 B.n84 585
R143 B.n654 B.n653 585
R144 B.n656 B.n83 585
R145 B.n659 B.n658 585
R146 B.n660 B.n82 585
R147 B.n662 B.n661 585
R148 B.n664 B.n81 585
R149 B.n667 B.n666 585
R150 B.n668 B.n80 585
R151 B.n541 B.n78 585
R152 B.n671 B.n78 585
R153 B.n540 B.n77 585
R154 B.n672 B.n77 585
R155 B.n539 B.n76 585
R156 B.n673 B.n76 585
R157 B.n538 B.n537 585
R158 B.n537 B.n72 585
R159 B.n536 B.n71 585
R160 B.n679 B.n71 585
R161 B.n535 B.n70 585
R162 B.n680 B.n70 585
R163 B.n534 B.n69 585
R164 B.n681 B.n69 585
R165 B.n533 B.n532 585
R166 B.n532 B.n68 585
R167 B.n531 B.n64 585
R168 B.n687 B.n64 585
R169 B.n530 B.n63 585
R170 B.n688 B.n63 585
R171 B.n529 B.n62 585
R172 B.n689 B.n62 585
R173 B.n528 B.n527 585
R174 B.n527 B.n58 585
R175 B.n526 B.n57 585
R176 B.n695 B.n57 585
R177 B.n525 B.n56 585
R178 B.n696 B.n56 585
R179 B.n524 B.n55 585
R180 B.n697 B.n55 585
R181 B.n523 B.n522 585
R182 B.n522 B.n51 585
R183 B.n521 B.n50 585
R184 B.n703 B.n50 585
R185 B.n520 B.n49 585
R186 B.n704 B.n49 585
R187 B.n519 B.n48 585
R188 B.n705 B.n48 585
R189 B.n518 B.n517 585
R190 B.n517 B.n47 585
R191 B.n516 B.n43 585
R192 B.n711 B.n43 585
R193 B.n515 B.n42 585
R194 B.n712 B.n42 585
R195 B.n514 B.n41 585
R196 B.n713 B.n41 585
R197 B.n513 B.n512 585
R198 B.n512 B.n37 585
R199 B.n511 B.n36 585
R200 B.n719 B.n36 585
R201 B.n510 B.n35 585
R202 B.n720 B.n35 585
R203 B.n509 B.n34 585
R204 B.n721 B.n34 585
R205 B.n508 B.n507 585
R206 B.n507 B.n30 585
R207 B.n506 B.n29 585
R208 B.n727 B.n29 585
R209 B.n505 B.n28 585
R210 B.n728 B.n28 585
R211 B.n504 B.n27 585
R212 B.n729 B.n27 585
R213 B.n503 B.n502 585
R214 B.n502 B.n23 585
R215 B.n501 B.n22 585
R216 B.n735 B.n22 585
R217 B.n500 B.n21 585
R218 B.n736 B.n21 585
R219 B.n499 B.n20 585
R220 B.n737 B.n20 585
R221 B.n498 B.n497 585
R222 B.n497 B.n16 585
R223 B.n496 B.n15 585
R224 B.n743 B.n15 585
R225 B.n495 B.n14 585
R226 B.n744 B.n14 585
R227 B.n494 B.n13 585
R228 B.n745 B.n13 585
R229 B.n493 B.n492 585
R230 B.n492 B.n12 585
R231 B.n491 B.n490 585
R232 B.n491 B.n8 585
R233 B.n489 B.n7 585
R234 B.n752 B.n7 585
R235 B.n488 B.n6 585
R236 B.n753 B.n6 585
R237 B.n487 B.n5 585
R238 B.n754 B.n5 585
R239 B.n486 B.n485 585
R240 B.n485 B.n4 585
R241 B.n484 B.n116 585
R242 B.n484 B.n483 585
R243 B.n474 B.n117 585
R244 B.n118 B.n117 585
R245 B.n476 B.n475 585
R246 B.n477 B.n476 585
R247 B.n473 B.n123 585
R248 B.n123 B.n122 585
R249 B.n472 B.n471 585
R250 B.n471 B.n470 585
R251 B.n125 B.n124 585
R252 B.n126 B.n125 585
R253 B.n463 B.n462 585
R254 B.n464 B.n463 585
R255 B.n461 B.n131 585
R256 B.n131 B.n130 585
R257 B.n460 B.n459 585
R258 B.n459 B.n458 585
R259 B.n133 B.n132 585
R260 B.n134 B.n133 585
R261 B.n451 B.n450 585
R262 B.n452 B.n451 585
R263 B.n449 B.n139 585
R264 B.n139 B.n138 585
R265 B.n448 B.n447 585
R266 B.n447 B.n446 585
R267 B.n141 B.n140 585
R268 B.n142 B.n141 585
R269 B.n439 B.n438 585
R270 B.n440 B.n439 585
R271 B.n437 B.n147 585
R272 B.n147 B.n146 585
R273 B.n436 B.n435 585
R274 B.n435 B.n434 585
R275 B.n149 B.n148 585
R276 B.n150 B.n149 585
R277 B.n427 B.n426 585
R278 B.n428 B.n427 585
R279 B.n425 B.n155 585
R280 B.n155 B.n154 585
R281 B.n424 B.n423 585
R282 B.n423 B.n422 585
R283 B.n157 B.n156 585
R284 B.n415 B.n157 585
R285 B.n414 B.n413 585
R286 B.n416 B.n414 585
R287 B.n412 B.n162 585
R288 B.n162 B.n161 585
R289 B.n411 B.n410 585
R290 B.n410 B.n409 585
R291 B.n164 B.n163 585
R292 B.n165 B.n164 585
R293 B.n402 B.n401 585
R294 B.n403 B.n402 585
R295 B.n400 B.n170 585
R296 B.n170 B.n169 585
R297 B.n399 B.n398 585
R298 B.n398 B.n397 585
R299 B.n172 B.n171 585
R300 B.n173 B.n172 585
R301 B.n390 B.n389 585
R302 B.n391 B.n390 585
R303 B.n388 B.n178 585
R304 B.n178 B.n177 585
R305 B.n387 B.n386 585
R306 B.n386 B.n385 585
R307 B.n180 B.n179 585
R308 B.n378 B.n180 585
R309 B.n377 B.n376 585
R310 B.n379 B.n377 585
R311 B.n375 B.n185 585
R312 B.n185 B.n184 585
R313 B.n374 B.n373 585
R314 B.n373 B.n372 585
R315 B.n187 B.n186 585
R316 B.n188 B.n187 585
R317 B.n365 B.n364 585
R318 B.n366 B.n365 585
R319 B.n363 B.n193 585
R320 B.n193 B.n192 585
R321 B.n362 B.n361 585
R322 B.n361 B.n360 585
R323 B.n357 B.n197 585
R324 B.n356 B.n355 585
R325 B.n353 B.n198 585
R326 B.n353 B.n196 585
R327 B.n352 B.n351 585
R328 B.n350 B.n349 585
R329 B.n348 B.n200 585
R330 B.n346 B.n345 585
R331 B.n344 B.n201 585
R332 B.n343 B.n342 585
R333 B.n340 B.n202 585
R334 B.n338 B.n337 585
R335 B.n336 B.n203 585
R336 B.n335 B.n334 585
R337 B.n332 B.n204 585
R338 B.n330 B.n329 585
R339 B.n328 B.n205 585
R340 B.n327 B.n326 585
R341 B.n324 B.n206 585
R342 B.n322 B.n321 585
R343 B.n320 B.n207 585
R344 B.n319 B.n318 585
R345 B.n316 B.n208 585
R346 B.n314 B.n313 585
R347 B.n312 B.n209 585
R348 B.n311 B.n310 585
R349 B.n308 B.n210 585
R350 B.n306 B.n305 585
R351 B.n303 B.n211 585
R352 B.n302 B.n301 585
R353 B.n299 B.n214 585
R354 B.n297 B.n296 585
R355 B.n295 B.n215 585
R356 B.n294 B.n293 585
R357 B.n291 B.n216 585
R358 B.n289 B.n288 585
R359 B.n287 B.n217 585
R360 B.n285 B.n284 585
R361 B.n282 B.n220 585
R362 B.n280 B.n279 585
R363 B.n278 B.n221 585
R364 B.n277 B.n276 585
R365 B.n274 B.n222 585
R366 B.n272 B.n271 585
R367 B.n270 B.n223 585
R368 B.n269 B.n268 585
R369 B.n266 B.n224 585
R370 B.n264 B.n263 585
R371 B.n262 B.n225 585
R372 B.n261 B.n260 585
R373 B.n258 B.n226 585
R374 B.n256 B.n255 585
R375 B.n254 B.n227 585
R376 B.n253 B.n252 585
R377 B.n250 B.n228 585
R378 B.n248 B.n247 585
R379 B.n246 B.n229 585
R380 B.n245 B.n244 585
R381 B.n242 B.n230 585
R382 B.n240 B.n239 585
R383 B.n238 B.n231 585
R384 B.n237 B.n236 585
R385 B.n234 B.n232 585
R386 B.n195 B.n194 585
R387 B.n359 B.n358 585
R388 B.n360 B.n359 585
R389 B.n191 B.n190 585
R390 B.n192 B.n191 585
R391 B.n368 B.n367 585
R392 B.n367 B.n366 585
R393 B.n369 B.n189 585
R394 B.n189 B.n188 585
R395 B.n371 B.n370 585
R396 B.n372 B.n371 585
R397 B.n183 B.n182 585
R398 B.n184 B.n183 585
R399 B.n381 B.n380 585
R400 B.n380 B.n379 585
R401 B.n382 B.n181 585
R402 B.n378 B.n181 585
R403 B.n384 B.n383 585
R404 B.n385 B.n384 585
R405 B.n176 B.n175 585
R406 B.n177 B.n176 585
R407 B.n393 B.n392 585
R408 B.n392 B.n391 585
R409 B.n394 B.n174 585
R410 B.n174 B.n173 585
R411 B.n396 B.n395 585
R412 B.n397 B.n396 585
R413 B.n168 B.n167 585
R414 B.n169 B.n168 585
R415 B.n405 B.n404 585
R416 B.n404 B.n403 585
R417 B.n406 B.n166 585
R418 B.n166 B.n165 585
R419 B.n408 B.n407 585
R420 B.n409 B.n408 585
R421 B.n160 B.n159 585
R422 B.n161 B.n160 585
R423 B.n418 B.n417 585
R424 B.n417 B.n416 585
R425 B.n419 B.n158 585
R426 B.n415 B.n158 585
R427 B.n421 B.n420 585
R428 B.n422 B.n421 585
R429 B.n153 B.n152 585
R430 B.n154 B.n153 585
R431 B.n430 B.n429 585
R432 B.n429 B.n428 585
R433 B.n431 B.n151 585
R434 B.n151 B.n150 585
R435 B.n433 B.n432 585
R436 B.n434 B.n433 585
R437 B.n145 B.n144 585
R438 B.n146 B.n145 585
R439 B.n442 B.n441 585
R440 B.n441 B.n440 585
R441 B.n443 B.n143 585
R442 B.n143 B.n142 585
R443 B.n445 B.n444 585
R444 B.n446 B.n445 585
R445 B.n137 B.n136 585
R446 B.n138 B.n137 585
R447 B.n454 B.n453 585
R448 B.n453 B.n452 585
R449 B.n455 B.n135 585
R450 B.n135 B.n134 585
R451 B.n457 B.n456 585
R452 B.n458 B.n457 585
R453 B.n129 B.n128 585
R454 B.n130 B.n129 585
R455 B.n466 B.n465 585
R456 B.n465 B.n464 585
R457 B.n467 B.n127 585
R458 B.n127 B.n126 585
R459 B.n469 B.n468 585
R460 B.n470 B.n469 585
R461 B.n121 B.n120 585
R462 B.n122 B.n121 585
R463 B.n479 B.n478 585
R464 B.n478 B.n477 585
R465 B.n480 B.n119 585
R466 B.n119 B.n118 585
R467 B.n482 B.n481 585
R468 B.n483 B.n482 585
R469 B.n3 B.n0 585
R470 B.n4 B.n3 585
R471 B.n751 B.n1 585
R472 B.n752 B.n751 585
R473 B.n750 B.n749 585
R474 B.n750 B.n8 585
R475 B.n748 B.n9 585
R476 B.n12 B.n9 585
R477 B.n747 B.n746 585
R478 B.n746 B.n745 585
R479 B.n11 B.n10 585
R480 B.n744 B.n11 585
R481 B.n742 B.n741 585
R482 B.n743 B.n742 585
R483 B.n740 B.n17 585
R484 B.n17 B.n16 585
R485 B.n739 B.n738 585
R486 B.n738 B.n737 585
R487 B.n19 B.n18 585
R488 B.n736 B.n19 585
R489 B.n734 B.n733 585
R490 B.n735 B.n734 585
R491 B.n732 B.n24 585
R492 B.n24 B.n23 585
R493 B.n731 B.n730 585
R494 B.n730 B.n729 585
R495 B.n26 B.n25 585
R496 B.n728 B.n26 585
R497 B.n726 B.n725 585
R498 B.n727 B.n726 585
R499 B.n724 B.n31 585
R500 B.n31 B.n30 585
R501 B.n723 B.n722 585
R502 B.n722 B.n721 585
R503 B.n33 B.n32 585
R504 B.n720 B.n33 585
R505 B.n718 B.n717 585
R506 B.n719 B.n718 585
R507 B.n716 B.n38 585
R508 B.n38 B.n37 585
R509 B.n715 B.n714 585
R510 B.n714 B.n713 585
R511 B.n40 B.n39 585
R512 B.n712 B.n40 585
R513 B.n710 B.n709 585
R514 B.n711 B.n710 585
R515 B.n708 B.n44 585
R516 B.n47 B.n44 585
R517 B.n707 B.n706 585
R518 B.n706 B.n705 585
R519 B.n46 B.n45 585
R520 B.n704 B.n46 585
R521 B.n702 B.n701 585
R522 B.n703 B.n702 585
R523 B.n700 B.n52 585
R524 B.n52 B.n51 585
R525 B.n699 B.n698 585
R526 B.n698 B.n697 585
R527 B.n54 B.n53 585
R528 B.n696 B.n54 585
R529 B.n694 B.n693 585
R530 B.n695 B.n694 585
R531 B.n692 B.n59 585
R532 B.n59 B.n58 585
R533 B.n691 B.n690 585
R534 B.n690 B.n689 585
R535 B.n61 B.n60 585
R536 B.n688 B.n61 585
R537 B.n686 B.n685 585
R538 B.n687 B.n686 585
R539 B.n684 B.n65 585
R540 B.n68 B.n65 585
R541 B.n683 B.n682 585
R542 B.n682 B.n681 585
R543 B.n67 B.n66 585
R544 B.n680 B.n67 585
R545 B.n678 B.n677 585
R546 B.n679 B.n678 585
R547 B.n676 B.n73 585
R548 B.n73 B.n72 585
R549 B.n675 B.n674 585
R550 B.n674 B.n673 585
R551 B.n75 B.n74 585
R552 B.n672 B.n75 585
R553 B.n670 B.n669 585
R554 B.n671 B.n670 585
R555 B.n755 B.n754 585
R556 B.n753 B.n2 585
R557 B.n670 B.n80 506.916
R558 B.n543 B.n78 506.916
R559 B.n361 B.n195 506.916
R560 B.n359 B.n197 506.916
R561 B.n95 B.t10 272.795
R562 B.n102 B.t6 272.795
R563 B.n218 B.t13 272.795
R564 B.n212 B.t17 272.795
R565 B.n544 B.n79 256.663
R566 B.n550 B.n79 256.663
R567 B.n552 B.n79 256.663
R568 B.n558 B.n79 256.663
R569 B.n560 B.n79 256.663
R570 B.n566 B.n79 256.663
R571 B.n568 B.n79 256.663
R572 B.n574 B.n79 256.663
R573 B.n576 B.n79 256.663
R574 B.n582 B.n79 256.663
R575 B.n584 B.n79 256.663
R576 B.n590 B.n79 256.663
R577 B.n592 B.n79 256.663
R578 B.n599 B.n79 256.663
R579 B.n601 B.n79 256.663
R580 B.n607 B.n79 256.663
R581 B.n609 B.n79 256.663
R582 B.n615 B.n79 256.663
R583 B.n617 B.n79 256.663
R584 B.n623 B.n79 256.663
R585 B.n625 B.n79 256.663
R586 B.n631 B.n79 256.663
R587 B.n633 B.n79 256.663
R588 B.n639 B.n79 256.663
R589 B.n641 B.n79 256.663
R590 B.n647 B.n79 256.663
R591 B.n649 B.n79 256.663
R592 B.n655 B.n79 256.663
R593 B.n657 B.n79 256.663
R594 B.n663 B.n79 256.663
R595 B.n665 B.n79 256.663
R596 B.n354 B.n196 256.663
R597 B.n199 B.n196 256.663
R598 B.n347 B.n196 256.663
R599 B.n341 B.n196 256.663
R600 B.n339 B.n196 256.663
R601 B.n333 B.n196 256.663
R602 B.n331 B.n196 256.663
R603 B.n325 B.n196 256.663
R604 B.n323 B.n196 256.663
R605 B.n317 B.n196 256.663
R606 B.n315 B.n196 256.663
R607 B.n309 B.n196 256.663
R608 B.n307 B.n196 256.663
R609 B.n300 B.n196 256.663
R610 B.n298 B.n196 256.663
R611 B.n292 B.n196 256.663
R612 B.n290 B.n196 256.663
R613 B.n283 B.n196 256.663
R614 B.n281 B.n196 256.663
R615 B.n275 B.n196 256.663
R616 B.n273 B.n196 256.663
R617 B.n267 B.n196 256.663
R618 B.n265 B.n196 256.663
R619 B.n259 B.n196 256.663
R620 B.n257 B.n196 256.663
R621 B.n251 B.n196 256.663
R622 B.n249 B.n196 256.663
R623 B.n243 B.n196 256.663
R624 B.n241 B.n196 256.663
R625 B.n235 B.n196 256.663
R626 B.n233 B.n196 256.663
R627 B.n757 B.n756 256.663
R628 B.n666 B.n664 163.367
R629 B.n662 B.n82 163.367
R630 B.n658 B.n656 163.367
R631 B.n654 B.n84 163.367
R632 B.n650 B.n648 163.367
R633 B.n646 B.n86 163.367
R634 B.n642 B.n640 163.367
R635 B.n638 B.n88 163.367
R636 B.n634 B.n632 163.367
R637 B.n630 B.n90 163.367
R638 B.n626 B.n624 163.367
R639 B.n622 B.n92 163.367
R640 B.n618 B.n616 163.367
R641 B.n614 B.n94 163.367
R642 B.n610 B.n608 163.367
R643 B.n606 B.n99 163.367
R644 B.n602 B.n600 163.367
R645 B.n598 B.n101 163.367
R646 B.n593 B.n591 163.367
R647 B.n589 B.n105 163.367
R648 B.n585 B.n583 163.367
R649 B.n581 B.n107 163.367
R650 B.n577 B.n575 163.367
R651 B.n573 B.n109 163.367
R652 B.n569 B.n567 163.367
R653 B.n565 B.n111 163.367
R654 B.n561 B.n559 163.367
R655 B.n557 B.n113 163.367
R656 B.n553 B.n551 163.367
R657 B.n549 B.n115 163.367
R658 B.n545 B.n543 163.367
R659 B.n361 B.n193 163.367
R660 B.n365 B.n193 163.367
R661 B.n365 B.n187 163.367
R662 B.n373 B.n187 163.367
R663 B.n373 B.n185 163.367
R664 B.n377 B.n185 163.367
R665 B.n377 B.n180 163.367
R666 B.n386 B.n180 163.367
R667 B.n386 B.n178 163.367
R668 B.n390 B.n178 163.367
R669 B.n390 B.n172 163.367
R670 B.n398 B.n172 163.367
R671 B.n398 B.n170 163.367
R672 B.n402 B.n170 163.367
R673 B.n402 B.n164 163.367
R674 B.n410 B.n164 163.367
R675 B.n410 B.n162 163.367
R676 B.n414 B.n162 163.367
R677 B.n414 B.n157 163.367
R678 B.n423 B.n157 163.367
R679 B.n423 B.n155 163.367
R680 B.n427 B.n155 163.367
R681 B.n427 B.n149 163.367
R682 B.n435 B.n149 163.367
R683 B.n435 B.n147 163.367
R684 B.n439 B.n147 163.367
R685 B.n439 B.n141 163.367
R686 B.n447 B.n141 163.367
R687 B.n447 B.n139 163.367
R688 B.n451 B.n139 163.367
R689 B.n451 B.n133 163.367
R690 B.n459 B.n133 163.367
R691 B.n459 B.n131 163.367
R692 B.n463 B.n131 163.367
R693 B.n463 B.n125 163.367
R694 B.n471 B.n125 163.367
R695 B.n471 B.n123 163.367
R696 B.n476 B.n123 163.367
R697 B.n476 B.n117 163.367
R698 B.n484 B.n117 163.367
R699 B.n485 B.n484 163.367
R700 B.n485 B.n5 163.367
R701 B.n6 B.n5 163.367
R702 B.n7 B.n6 163.367
R703 B.n491 B.n7 163.367
R704 B.n492 B.n491 163.367
R705 B.n492 B.n13 163.367
R706 B.n14 B.n13 163.367
R707 B.n15 B.n14 163.367
R708 B.n497 B.n15 163.367
R709 B.n497 B.n20 163.367
R710 B.n21 B.n20 163.367
R711 B.n22 B.n21 163.367
R712 B.n502 B.n22 163.367
R713 B.n502 B.n27 163.367
R714 B.n28 B.n27 163.367
R715 B.n29 B.n28 163.367
R716 B.n507 B.n29 163.367
R717 B.n507 B.n34 163.367
R718 B.n35 B.n34 163.367
R719 B.n36 B.n35 163.367
R720 B.n512 B.n36 163.367
R721 B.n512 B.n41 163.367
R722 B.n42 B.n41 163.367
R723 B.n43 B.n42 163.367
R724 B.n517 B.n43 163.367
R725 B.n517 B.n48 163.367
R726 B.n49 B.n48 163.367
R727 B.n50 B.n49 163.367
R728 B.n522 B.n50 163.367
R729 B.n522 B.n55 163.367
R730 B.n56 B.n55 163.367
R731 B.n57 B.n56 163.367
R732 B.n527 B.n57 163.367
R733 B.n527 B.n62 163.367
R734 B.n63 B.n62 163.367
R735 B.n64 B.n63 163.367
R736 B.n532 B.n64 163.367
R737 B.n532 B.n69 163.367
R738 B.n70 B.n69 163.367
R739 B.n71 B.n70 163.367
R740 B.n537 B.n71 163.367
R741 B.n537 B.n76 163.367
R742 B.n77 B.n76 163.367
R743 B.n78 B.n77 163.367
R744 B.n355 B.n353 163.367
R745 B.n353 B.n352 163.367
R746 B.n349 B.n348 163.367
R747 B.n346 B.n201 163.367
R748 B.n342 B.n340 163.367
R749 B.n338 B.n203 163.367
R750 B.n334 B.n332 163.367
R751 B.n330 B.n205 163.367
R752 B.n326 B.n324 163.367
R753 B.n322 B.n207 163.367
R754 B.n318 B.n316 163.367
R755 B.n314 B.n209 163.367
R756 B.n310 B.n308 163.367
R757 B.n306 B.n211 163.367
R758 B.n301 B.n299 163.367
R759 B.n297 B.n215 163.367
R760 B.n293 B.n291 163.367
R761 B.n289 B.n217 163.367
R762 B.n284 B.n282 163.367
R763 B.n280 B.n221 163.367
R764 B.n276 B.n274 163.367
R765 B.n272 B.n223 163.367
R766 B.n268 B.n266 163.367
R767 B.n264 B.n225 163.367
R768 B.n260 B.n258 163.367
R769 B.n256 B.n227 163.367
R770 B.n252 B.n250 163.367
R771 B.n248 B.n229 163.367
R772 B.n244 B.n242 163.367
R773 B.n240 B.n231 163.367
R774 B.n236 B.n234 163.367
R775 B.n359 B.n191 163.367
R776 B.n367 B.n191 163.367
R777 B.n367 B.n189 163.367
R778 B.n371 B.n189 163.367
R779 B.n371 B.n183 163.367
R780 B.n380 B.n183 163.367
R781 B.n380 B.n181 163.367
R782 B.n384 B.n181 163.367
R783 B.n384 B.n176 163.367
R784 B.n392 B.n176 163.367
R785 B.n392 B.n174 163.367
R786 B.n396 B.n174 163.367
R787 B.n396 B.n168 163.367
R788 B.n404 B.n168 163.367
R789 B.n404 B.n166 163.367
R790 B.n408 B.n166 163.367
R791 B.n408 B.n160 163.367
R792 B.n417 B.n160 163.367
R793 B.n417 B.n158 163.367
R794 B.n421 B.n158 163.367
R795 B.n421 B.n153 163.367
R796 B.n429 B.n153 163.367
R797 B.n429 B.n151 163.367
R798 B.n433 B.n151 163.367
R799 B.n433 B.n145 163.367
R800 B.n441 B.n145 163.367
R801 B.n441 B.n143 163.367
R802 B.n445 B.n143 163.367
R803 B.n445 B.n137 163.367
R804 B.n453 B.n137 163.367
R805 B.n453 B.n135 163.367
R806 B.n457 B.n135 163.367
R807 B.n457 B.n129 163.367
R808 B.n465 B.n129 163.367
R809 B.n465 B.n127 163.367
R810 B.n469 B.n127 163.367
R811 B.n469 B.n121 163.367
R812 B.n478 B.n121 163.367
R813 B.n478 B.n119 163.367
R814 B.n482 B.n119 163.367
R815 B.n482 B.n3 163.367
R816 B.n755 B.n3 163.367
R817 B.n751 B.n2 163.367
R818 B.n751 B.n750 163.367
R819 B.n750 B.n9 163.367
R820 B.n746 B.n9 163.367
R821 B.n746 B.n11 163.367
R822 B.n742 B.n11 163.367
R823 B.n742 B.n17 163.367
R824 B.n738 B.n17 163.367
R825 B.n738 B.n19 163.367
R826 B.n734 B.n19 163.367
R827 B.n734 B.n24 163.367
R828 B.n730 B.n24 163.367
R829 B.n730 B.n26 163.367
R830 B.n726 B.n26 163.367
R831 B.n726 B.n31 163.367
R832 B.n722 B.n31 163.367
R833 B.n722 B.n33 163.367
R834 B.n718 B.n33 163.367
R835 B.n718 B.n38 163.367
R836 B.n714 B.n38 163.367
R837 B.n714 B.n40 163.367
R838 B.n710 B.n40 163.367
R839 B.n710 B.n44 163.367
R840 B.n706 B.n44 163.367
R841 B.n706 B.n46 163.367
R842 B.n702 B.n46 163.367
R843 B.n702 B.n52 163.367
R844 B.n698 B.n52 163.367
R845 B.n698 B.n54 163.367
R846 B.n694 B.n54 163.367
R847 B.n694 B.n59 163.367
R848 B.n690 B.n59 163.367
R849 B.n690 B.n61 163.367
R850 B.n686 B.n61 163.367
R851 B.n686 B.n65 163.367
R852 B.n682 B.n65 163.367
R853 B.n682 B.n67 163.367
R854 B.n678 B.n67 163.367
R855 B.n678 B.n73 163.367
R856 B.n674 B.n73 163.367
R857 B.n674 B.n75 163.367
R858 B.n670 B.n75 163.367
R859 B.n102 B.t8 128.714
R860 B.n218 B.t16 128.714
R861 B.n95 B.t11 128.707
R862 B.n212 B.t19 128.707
R863 B.n360 B.n196 108.787
R864 B.n671 B.n79 108.787
R865 B.n103 B.t9 72.0843
R866 B.n219 B.t15 72.0843
R867 B.n96 B.t12 72.0765
R868 B.n213 B.t18 72.0765
R869 B.n665 B.n80 71.676
R870 B.n664 B.n663 71.676
R871 B.n657 B.n82 71.676
R872 B.n656 B.n655 71.676
R873 B.n649 B.n84 71.676
R874 B.n648 B.n647 71.676
R875 B.n641 B.n86 71.676
R876 B.n640 B.n639 71.676
R877 B.n633 B.n88 71.676
R878 B.n632 B.n631 71.676
R879 B.n625 B.n90 71.676
R880 B.n624 B.n623 71.676
R881 B.n617 B.n92 71.676
R882 B.n616 B.n615 71.676
R883 B.n609 B.n94 71.676
R884 B.n608 B.n607 71.676
R885 B.n601 B.n99 71.676
R886 B.n600 B.n599 71.676
R887 B.n592 B.n101 71.676
R888 B.n591 B.n590 71.676
R889 B.n584 B.n105 71.676
R890 B.n583 B.n582 71.676
R891 B.n576 B.n107 71.676
R892 B.n575 B.n574 71.676
R893 B.n568 B.n109 71.676
R894 B.n567 B.n566 71.676
R895 B.n560 B.n111 71.676
R896 B.n559 B.n558 71.676
R897 B.n552 B.n113 71.676
R898 B.n551 B.n550 71.676
R899 B.n544 B.n115 71.676
R900 B.n545 B.n544 71.676
R901 B.n550 B.n549 71.676
R902 B.n553 B.n552 71.676
R903 B.n558 B.n557 71.676
R904 B.n561 B.n560 71.676
R905 B.n566 B.n565 71.676
R906 B.n569 B.n568 71.676
R907 B.n574 B.n573 71.676
R908 B.n577 B.n576 71.676
R909 B.n582 B.n581 71.676
R910 B.n585 B.n584 71.676
R911 B.n590 B.n589 71.676
R912 B.n593 B.n592 71.676
R913 B.n599 B.n598 71.676
R914 B.n602 B.n601 71.676
R915 B.n607 B.n606 71.676
R916 B.n610 B.n609 71.676
R917 B.n615 B.n614 71.676
R918 B.n618 B.n617 71.676
R919 B.n623 B.n622 71.676
R920 B.n626 B.n625 71.676
R921 B.n631 B.n630 71.676
R922 B.n634 B.n633 71.676
R923 B.n639 B.n638 71.676
R924 B.n642 B.n641 71.676
R925 B.n647 B.n646 71.676
R926 B.n650 B.n649 71.676
R927 B.n655 B.n654 71.676
R928 B.n658 B.n657 71.676
R929 B.n663 B.n662 71.676
R930 B.n666 B.n665 71.676
R931 B.n354 B.n197 71.676
R932 B.n352 B.n199 71.676
R933 B.n348 B.n347 71.676
R934 B.n341 B.n201 71.676
R935 B.n340 B.n339 71.676
R936 B.n333 B.n203 71.676
R937 B.n332 B.n331 71.676
R938 B.n325 B.n205 71.676
R939 B.n324 B.n323 71.676
R940 B.n317 B.n207 71.676
R941 B.n316 B.n315 71.676
R942 B.n309 B.n209 71.676
R943 B.n308 B.n307 71.676
R944 B.n300 B.n211 71.676
R945 B.n299 B.n298 71.676
R946 B.n292 B.n215 71.676
R947 B.n291 B.n290 71.676
R948 B.n283 B.n217 71.676
R949 B.n282 B.n281 71.676
R950 B.n275 B.n221 71.676
R951 B.n274 B.n273 71.676
R952 B.n267 B.n223 71.676
R953 B.n266 B.n265 71.676
R954 B.n259 B.n225 71.676
R955 B.n258 B.n257 71.676
R956 B.n251 B.n227 71.676
R957 B.n250 B.n249 71.676
R958 B.n243 B.n229 71.676
R959 B.n242 B.n241 71.676
R960 B.n235 B.n231 71.676
R961 B.n234 B.n233 71.676
R962 B.n355 B.n354 71.676
R963 B.n349 B.n199 71.676
R964 B.n347 B.n346 71.676
R965 B.n342 B.n341 71.676
R966 B.n339 B.n338 71.676
R967 B.n334 B.n333 71.676
R968 B.n331 B.n330 71.676
R969 B.n326 B.n325 71.676
R970 B.n323 B.n322 71.676
R971 B.n318 B.n317 71.676
R972 B.n315 B.n314 71.676
R973 B.n310 B.n309 71.676
R974 B.n307 B.n306 71.676
R975 B.n301 B.n300 71.676
R976 B.n298 B.n297 71.676
R977 B.n293 B.n292 71.676
R978 B.n290 B.n289 71.676
R979 B.n284 B.n283 71.676
R980 B.n281 B.n280 71.676
R981 B.n276 B.n275 71.676
R982 B.n273 B.n272 71.676
R983 B.n268 B.n267 71.676
R984 B.n265 B.n264 71.676
R985 B.n260 B.n259 71.676
R986 B.n257 B.n256 71.676
R987 B.n252 B.n251 71.676
R988 B.n249 B.n248 71.676
R989 B.n244 B.n243 71.676
R990 B.n241 B.n240 71.676
R991 B.n236 B.n235 71.676
R992 B.n233 B.n195 71.676
R993 B.n756 B.n755 71.676
R994 B.n756 B.n2 71.676
R995 B.n360 B.n192 61.1366
R996 B.n366 B.n192 61.1366
R997 B.n366 B.n188 61.1366
R998 B.n372 B.n188 61.1366
R999 B.n372 B.n184 61.1366
R1000 B.n379 B.n184 61.1366
R1001 B.n379 B.n378 61.1366
R1002 B.n385 B.n177 61.1366
R1003 B.n391 B.n177 61.1366
R1004 B.n391 B.n173 61.1366
R1005 B.n397 B.n173 61.1366
R1006 B.n397 B.n169 61.1366
R1007 B.n403 B.n169 61.1366
R1008 B.n403 B.n165 61.1366
R1009 B.n409 B.n165 61.1366
R1010 B.n409 B.n161 61.1366
R1011 B.n416 B.n161 61.1366
R1012 B.n416 B.n415 61.1366
R1013 B.n422 B.n154 61.1366
R1014 B.n428 B.n154 61.1366
R1015 B.n428 B.n150 61.1366
R1016 B.n434 B.n150 61.1366
R1017 B.n434 B.n146 61.1366
R1018 B.n440 B.n146 61.1366
R1019 B.n440 B.n142 61.1366
R1020 B.n446 B.n142 61.1366
R1021 B.n452 B.n138 61.1366
R1022 B.n452 B.n134 61.1366
R1023 B.n458 B.n134 61.1366
R1024 B.n458 B.n130 61.1366
R1025 B.n464 B.n130 61.1366
R1026 B.n464 B.n126 61.1366
R1027 B.n470 B.n126 61.1366
R1028 B.n477 B.n122 61.1366
R1029 B.n477 B.n118 61.1366
R1030 B.n483 B.n118 61.1366
R1031 B.n483 B.n4 61.1366
R1032 B.n754 B.n4 61.1366
R1033 B.n754 B.n753 61.1366
R1034 B.n753 B.n752 61.1366
R1035 B.n752 B.n8 61.1366
R1036 B.n12 B.n8 61.1366
R1037 B.n745 B.n12 61.1366
R1038 B.n745 B.n744 61.1366
R1039 B.n743 B.n16 61.1366
R1040 B.n737 B.n16 61.1366
R1041 B.n737 B.n736 61.1366
R1042 B.n736 B.n735 61.1366
R1043 B.n735 B.n23 61.1366
R1044 B.n729 B.n23 61.1366
R1045 B.n729 B.n728 61.1366
R1046 B.n727 B.n30 61.1366
R1047 B.n721 B.n30 61.1366
R1048 B.n721 B.n720 61.1366
R1049 B.n720 B.n719 61.1366
R1050 B.n719 B.n37 61.1366
R1051 B.n713 B.n37 61.1366
R1052 B.n713 B.n712 61.1366
R1053 B.n712 B.n711 61.1366
R1054 B.n705 B.n47 61.1366
R1055 B.n705 B.n704 61.1366
R1056 B.n704 B.n703 61.1366
R1057 B.n703 B.n51 61.1366
R1058 B.n697 B.n51 61.1366
R1059 B.n697 B.n696 61.1366
R1060 B.n696 B.n695 61.1366
R1061 B.n695 B.n58 61.1366
R1062 B.n689 B.n58 61.1366
R1063 B.n689 B.n688 61.1366
R1064 B.n688 B.n687 61.1366
R1065 B.n681 B.n68 61.1366
R1066 B.n681 B.n680 61.1366
R1067 B.n680 B.n679 61.1366
R1068 B.n679 B.n72 61.1366
R1069 B.n673 B.n72 61.1366
R1070 B.n673 B.n672 61.1366
R1071 B.n672 B.n671 61.1366
R1072 B.t5 B.n138 60.2375
R1073 B.n728 B.t4 60.2375
R1074 B.n97 B.n96 59.5399
R1075 B.n596 B.n103 59.5399
R1076 B.n286 B.n219 59.5399
R1077 B.n304 B.n213 59.5399
R1078 B.n96 B.n95 56.6308
R1079 B.n103 B.n102 56.6308
R1080 B.n219 B.n218 56.6308
R1081 B.n213 B.n212 56.6308
R1082 B.n378 B.t14 38.6601
R1083 B.n68 B.t7 38.6601
R1084 B.n470 B.t0 36.862
R1085 B.t3 B.n743 36.862
R1086 B.n422 B.t1 35.0638
R1087 B.n711 B.t2 35.0638
R1088 B.n358 B.n357 32.9371
R1089 B.n362 B.n194 32.9371
R1090 B.n542 B.n541 32.9371
R1091 B.n669 B.n668 32.9371
R1092 B.n415 B.t1 26.0732
R1093 B.n47 B.t2 26.0732
R1094 B.t0 B.n122 24.2751
R1095 B.n744 B.t3 24.2751
R1096 B.n385 B.t14 22.477
R1097 B.n687 B.t7 22.477
R1098 B B.n757 18.0485
R1099 B.n358 B.n190 10.6151
R1100 B.n368 B.n190 10.6151
R1101 B.n369 B.n368 10.6151
R1102 B.n370 B.n369 10.6151
R1103 B.n370 B.n182 10.6151
R1104 B.n381 B.n182 10.6151
R1105 B.n382 B.n381 10.6151
R1106 B.n383 B.n382 10.6151
R1107 B.n383 B.n175 10.6151
R1108 B.n393 B.n175 10.6151
R1109 B.n394 B.n393 10.6151
R1110 B.n395 B.n394 10.6151
R1111 B.n395 B.n167 10.6151
R1112 B.n405 B.n167 10.6151
R1113 B.n406 B.n405 10.6151
R1114 B.n407 B.n406 10.6151
R1115 B.n407 B.n159 10.6151
R1116 B.n418 B.n159 10.6151
R1117 B.n419 B.n418 10.6151
R1118 B.n420 B.n419 10.6151
R1119 B.n420 B.n152 10.6151
R1120 B.n430 B.n152 10.6151
R1121 B.n431 B.n430 10.6151
R1122 B.n432 B.n431 10.6151
R1123 B.n432 B.n144 10.6151
R1124 B.n442 B.n144 10.6151
R1125 B.n443 B.n442 10.6151
R1126 B.n444 B.n443 10.6151
R1127 B.n444 B.n136 10.6151
R1128 B.n454 B.n136 10.6151
R1129 B.n455 B.n454 10.6151
R1130 B.n456 B.n455 10.6151
R1131 B.n456 B.n128 10.6151
R1132 B.n466 B.n128 10.6151
R1133 B.n467 B.n466 10.6151
R1134 B.n468 B.n467 10.6151
R1135 B.n468 B.n120 10.6151
R1136 B.n479 B.n120 10.6151
R1137 B.n480 B.n479 10.6151
R1138 B.n481 B.n480 10.6151
R1139 B.n481 B.n0 10.6151
R1140 B.n357 B.n356 10.6151
R1141 B.n356 B.n198 10.6151
R1142 B.n351 B.n198 10.6151
R1143 B.n351 B.n350 10.6151
R1144 B.n350 B.n200 10.6151
R1145 B.n345 B.n200 10.6151
R1146 B.n345 B.n344 10.6151
R1147 B.n344 B.n343 10.6151
R1148 B.n343 B.n202 10.6151
R1149 B.n337 B.n202 10.6151
R1150 B.n337 B.n336 10.6151
R1151 B.n336 B.n335 10.6151
R1152 B.n335 B.n204 10.6151
R1153 B.n329 B.n204 10.6151
R1154 B.n329 B.n328 10.6151
R1155 B.n328 B.n327 10.6151
R1156 B.n327 B.n206 10.6151
R1157 B.n321 B.n206 10.6151
R1158 B.n321 B.n320 10.6151
R1159 B.n320 B.n319 10.6151
R1160 B.n319 B.n208 10.6151
R1161 B.n313 B.n208 10.6151
R1162 B.n313 B.n312 10.6151
R1163 B.n312 B.n311 10.6151
R1164 B.n311 B.n210 10.6151
R1165 B.n305 B.n210 10.6151
R1166 B.n303 B.n302 10.6151
R1167 B.n302 B.n214 10.6151
R1168 B.n296 B.n214 10.6151
R1169 B.n296 B.n295 10.6151
R1170 B.n295 B.n294 10.6151
R1171 B.n294 B.n216 10.6151
R1172 B.n288 B.n216 10.6151
R1173 B.n288 B.n287 10.6151
R1174 B.n285 B.n220 10.6151
R1175 B.n279 B.n220 10.6151
R1176 B.n279 B.n278 10.6151
R1177 B.n278 B.n277 10.6151
R1178 B.n277 B.n222 10.6151
R1179 B.n271 B.n222 10.6151
R1180 B.n271 B.n270 10.6151
R1181 B.n270 B.n269 10.6151
R1182 B.n269 B.n224 10.6151
R1183 B.n263 B.n224 10.6151
R1184 B.n263 B.n262 10.6151
R1185 B.n262 B.n261 10.6151
R1186 B.n261 B.n226 10.6151
R1187 B.n255 B.n226 10.6151
R1188 B.n255 B.n254 10.6151
R1189 B.n254 B.n253 10.6151
R1190 B.n253 B.n228 10.6151
R1191 B.n247 B.n228 10.6151
R1192 B.n247 B.n246 10.6151
R1193 B.n246 B.n245 10.6151
R1194 B.n245 B.n230 10.6151
R1195 B.n239 B.n230 10.6151
R1196 B.n239 B.n238 10.6151
R1197 B.n238 B.n237 10.6151
R1198 B.n237 B.n232 10.6151
R1199 B.n232 B.n194 10.6151
R1200 B.n363 B.n362 10.6151
R1201 B.n364 B.n363 10.6151
R1202 B.n364 B.n186 10.6151
R1203 B.n374 B.n186 10.6151
R1204 B.n375 B.n374 10.6151
R1205 B.n376 B.n375 10.6151
R1206 B.n376 B.n179 10.6151
R1207 B.n387 B.n179 10.6151
R1208 B.n388 B.n387 10.6151
R1209 B.n389 B.n388 10.6151
R1210 B.n389 B.n171 10.6151
R1211 B.n399 B.n171 10.6151
R1212 B.n400 B.n399 10.6151
R1213 B.n401 B.n400 10.6151
R1214 B.n401 B.n163 10.6151
R1215 B.n411 B.n163 10.6151
R1216 B.n412 B.n411 10.6151
R1217 B.n413 B.n412 10.6151
R1218 B.n413 B.n156 10.6151
R1219 B.n424 B.n156 10.6151
R1220 B.n425 B.n424 10.6151
R1221 B.n426 B.n425 10.6151
R1222 B.n426 B.n148 10.6151
R1223 B.n436 B.n148 10.6151
R1224 B.n437 B.n436 10.6151
R1225 B.n438 B.n437 10.6151
R1226 B.n438 B.n140 10.6151
R1227 B.n448 B.n140 10.6151
R1228 B.n449 B.n448 10.6151
R1229 B.n450 B.n449 10.6151
R1230 B.n450 B.n132 10.6151
R1231 B.n460 B.n132 10.6151
R1232 B.n461 B.n460 10.6151
R1233 B.n462 B.n461 10.6151
R1234 B.n462 B.n124 10.6151
R1235 B.n472 B.n124 10.6151
R1236 B.n473 B.n472 10.6151
R1237 B.n475 B.n473 10.6151
R1238 B.n475 B.n474 10.6151
R1239 B.n474 B.n116 10.6151
R1240 B.n486 B.n116 10.6151
R1241 B.n487 B.n486 10.6151
R1242 B.n488 B.n487 10.6151
R1243 B.n489 B.n488 10.6151
R1244 B.n490 B.n489 10.6151
R1245 B.n493 B.n490 10.6151
R1246 B.n494 B.n493 10.6151
R1247 B.n495 B.n494 10.6151
R1248 B.n496 B.n495 10.6151
R1249 B.n498 B.n496 10.6151
R1250 B.n499 B.n498 10.6151
R1251 B.n500 B.n499 10.6151
R1252 B.n501 B.n500 10.6151
R1253 B.n503 B.n501 10.6151
R1254 B.n504 B.n503 10.6151
R1255 B.n505 B.n504 10.6151
R1256 B.n506 B.n505 10.6151
R1257 B.n508 B.n506 10.6151
R1258 B.n509 B.n508 10.6151
R1259 B.n510 B.n509 10.6151
R1260 B.n511 B.n510 10.6151
R1261 B.n513 B.n511 10.6151
R1262 B.n514 B.n513 10.6151
R1263 B.n515 B.n514 10.6151
R1264 B.n516 B.n515 10.6151
R1265 B.n518 B.n516 10.6151
R1266 B.n519 B.n518 10.6151
R1267 B.n520 B.n519 10.6151
R1268 B.n521 B.n520 10.6151
R1269 B.n523 B.n521 10.6151
R1270 B.n524 B.n523 10.6151
R1271 B.n525 B.n524 10.6151
R1272 B.n526 B.n525 10.6151
R1273 B.n528 B.n526 10.6151
R1274 B.n529 B.n528 10.6151
R1275 B.n530 B.n529 10.6151
R1276 B.n531 B.n530 10.6151
R1277 B.n533 B.n531 10.6151
R1278 B.n534 B.n533 10.6151
R1279 B.n535 B.n534 10.6151
R1280 B.n536 B.n535 10.6151
R1281 B.n538 B.n536 10.6151
R1282 B.n539 B.n538 10.6151
R1283 B.n540 B.n539 10.6151
R1284 B.n541 B.n540 10.6151
R1285 B.n749 B.n1 10.6151
R1286 B.n749 B.n748 10.6151
R1287 B.n748 B.n747 10.6151
R1288 B.n747 B.n10 10.6151
R1289 B.n741 B.n10 10.6151
R1290 B.n741 B.n740 10.6151
R1291 B.n740 B.n739 10.6151
R1292 B.n739 B.n18 10.6151
R1293 B.n733 B.n18 10.6151
R1294 B.n733 B.n732 10.6151
R1295 B.n732 B.n731 10.6151
R1296 B.n731 B.n25 10.6151
R1297 B.n725 B.n25 10.6151
R1298 B.n725 B.n724 10.6151
R1299 B.n724 B.n723 10.6151
R1300 B.n723 B.n32 10.6151
R1301 B.n717 B.n32 10.6151
R1302 B.n717 B.n716 10.6151
R1303 B.n716 B.n715 10.6151
R1304 B.n715 B.n39 10.6151
R1305 B.n709 B.n39 10.6151
R1306 B.n709 B.n708 10.6151
R1307 B.n708 B.n707 10.6151
R1308 B.n707 B.n45 10.6151
R1309 B.n701 B.n45 10.6151
R1310 B.n701 B.n700 10.6151
R1311 B.n700 B.n699 10.6151
R1312 B.n699 B.n53 10.6151
R1313 B.n693 B.n53 10.6151
R1314 B.n693 B.n692 10.6151
R1315 B.n692 B.n691 10.6151
R1316 B.n691 B.n60 10.6151
R1317 B.n685 B.n60 10.6151
R1318 B.n685 B.n684 10.6151
R1319 B.n684 B.n683 10.6151
R1320 B.n683 B.n66 10.6151
R1321 B.n677 B.n66 10.6151
R1322 B.n677 B.n676 10.6151
R1323 B.n676 B.n675 10.6151
R1324 B.n675 B.n74 10.6151
R1325 B.n669 B.n74 10.6151
R1326 B.n668 B.n667 10.6151
R1327 B.n667 B.n81 10.6151
R1328 B.n661 B.n81 10.6151
R1329 B.n661 B.n660 10.6151
R1330 B.n660 B.n659 10.6151
R1331 B.n659 B.n83 10.6151
R1332 B.n653 B.n83 10.6151
R1333 B.n653 B.n652 10.6151
R1334 B.n652 B.n651 10.6151
R1335 B.n651 B.n85 10.6151
R1336 B.n645 B.n85 10.6151
R1337 B.n645 B.n644 10.6151
R1338 B.n644 B.n643 10.6151
R1339 B.n643 B.n87 10.6151
R1340 B.n637 B.n87 10.6151
R1341 B.n637 B.n636 10.6151
R1342 B.n636 B.n635 10.6151
R1343 B.n635 B.n89 10.6151
R1344 B.n629 B.n89 10.6151
R1345 B.n629 B.n628 10.6151
R1346 B.n628 B.n627 10.6151
R1347 B.n627 B.n91 10.6151
R1348 B.n621 B.n91 10.6151
R1349 B.n621 B.n620 10.6151
R1350 B.n620 B.n619 10.6151
R1351 B.n619 B.n93 10.6151
R1352 B.n613 B.n612 10.6151
R1353 B.n612 B.n611 10.6151
R1354 B.n611 B.n98 10.6151
R1355 B.n605 B.n98 10.6151
R1356 B.n605 B.n604 10.6151
R1357 B.n604 B.n603 10.6151
R1358 B.n603 B.n100 10.6151
R1359 B.n597 B.n100 10.6151
R1360 B.n595 B.n594 10.6151
R1361 B.n594 B.n104 10.6151
R1362 B.n588 B.n104 10.6151
R1363 B.n588 B.n587 10.6151
R1364 B.n587 B.n586 10.6151
R1365 B.n586 B.n106 10.6151
R1366 B.n580 B.n106 10.6151
R1367 B.n580 B.n579 10.6151
R1368 B.n579 B.n578 10.6151
R1369 B.n578 B.n108 10.6151
R1370 B.n572 B.n108 10.6151
R1371 B.n572 B.n571 10.6151
R1372 B.n571 B.n570 10.6151
R1373 B.n570 B.n110 10.6151
R1374 B.n564 B.n110 10.6151
R1375 B.n564 B.n563 10.6151
R1376 B.n563 B.n562 10.6151
R1377 B.n562 B.n112 10.6151
R1378 B.n556 B.n112 10.6151
R1379 B.n556 B.n555 10.6151
R1380 B.n555 B.n554 10.6151
R1381 B.n554 B.n114 10.6151
R1382 B.n548 B.n114 10.6151
R1383 B.n548 B.n547 10.6151
R1384 B.n547 B.n546 10.6151
R1385 B.n546 B.n542 10.6151
R1386 B.n757 B.n0 8.11757
R1387 B.n757 B.n1 8.11757
R1388 B.n304 B.n303 6.5566
R1389 B.n287 B.n286 6.5566
R1390 B.n613 B.n97 6.5566
R1391 B.n597 B.n596 6.5566
R1392 B.n305 B.n304 4.05904
R1393 B.n286 B.n285 4.05904
R1394 B.n97 B.n93 4.05904
R1395 B.n596 B.n595 4.05904
R1396 B.n446 B.t5 0.89956
R1397 B.t4 B.n727 0.89956
R1398 VP.n13 VP.n12 161.3
R1399 VP.n14 VP.n9 161.3
R1400 VP.n16 VP.n15 161.3
R1401 VP.n17 VP.n8 161.3
R1402 VP.n19 VP.n18 161.3
R1403 VP.n20 VP.n7 161.3
R1404 VP.n42 VP.n0 161.3
R1405 VP.n41 VP.n40 161.3
R1406 VP.n39 VP.n1 161.3
R1407 VP.n38 VP.n37 161.3
R1408 VP.n36 VP.n2 161.3
R1409 VP.n35 VP.n34 161.3
R1410 VP.n33 VP.n32 161.3
R1411 VP.n31 VP.n4 161.3
R1412 VP.n30 VP.n29 161.3
R1413 VP.n28 VP.n5 161.3
R1414 VP.n27 VP.n26 161.3
R1415 VP.n25 VP.n6 161.3
R1416 VP.n24 VP.n23 102.547
R1417 VP.n44 VP.n43 102.547
R1418 VP.n22 VP.n21 102.547
R1419 VP.n11 VP.t0 97.9633
R1420 VP.n24 VP.t4 64.7634
R1421 VP.n3 VP.t2 64.7634
R1422 VP.n43 VP.t3 64.7634
R1423 VP.n21 VP.t5 64.7634
R1424 VP.n10 VP.t1 64.7634
R1425 VP.n11 VP.n10 60.2807
R1426 VP.n30 VP.n5 56.5617
R1427 VP.n37 VP.n1 56.5617
R1428 VP.n15 VP.n8 56.5617
R1429 VP.n23 VP.n22 44.8103
R1430 VP.n26 VP.n25 24.5923
R1431 VP.n26 VP.n5 24.5923
R1432 VP.n31 VP.n30 24.5923
R1433 VP.n32 VP.n31 24.5923
R1434 VP.n36 VP.n35 24.5923
R1435 VP.n37 VP.n36 24.5923
R1436 VP.n41 VP.n1 24.5923
R1437 VP.n42 VP.n41 24.5923
R1438 VP.n19 VP.n8 24.5923
R1439 VP.n20 VP.n19 24.5923
R1440 VP.n14 VP.n13 24.5923
R1441 VP.n15 VP.n14 24.5923
R1442 VP.n32 VP.n3 12.2964
R1443 VP.n35 VP.n3 12.2964
R1444 VP.n13 VP.n10 12.2964
R1445 VP.n25 VP.n24 8.36172
R1446 VP.n43 VP.n42 8.36172
R1447 VP.n21 VP.n20 8.36172
R1448 VP.n12 VP.n11 6.93618
R1449 VP.n22 VP.n7 0.278335
R1450 VP.n23 VP.n6 0.278335
R1451 VP.n44 VP.n0 0.278335
R1452 VP.n12 VP.n9 0.189894
R1453 VP.n16 VP.n9 0.189894
R1454 VP.n17 VP.n16 0.189894
R1455 VP.n18 VP.n17 0.189894
R1456 VP.n18 VP.n7 0.189894
R1457 VP.n27 VP.n6 0.189894
R1458 VP.n28 VP.n27 0.189894
R1459 VP.n29 VP.n28 0.189894
R1460 VP.n29 VP.n4 0.189894
R1461 VP.n33 VP.n4 0.189894
R1462 VP.n34 VP.n33 0.189894
R1463 VP.n34 VP.n2 0.189894
R1464 VP.n38 VP.n2 0.189894
R1465 VP.n39 VP.n38 0.189894
R1466 VP.n40 VP.n39 0.189894
R1467 VP.n40 VP.n0 0.189894
R1468 VP VP.n44 0.153485
R1469 VDD1 VDD1.t5 68.0749
R1470 VDD1.n1 VDD1.t1 67.9612
R1471 VDD1.n1 VDD1.n0 63.8579
R1472 VDD1.n3 VDD1.n2 63.2838
R1473 VDD1.n3 VDD1.n1 39.738
R1474 VDD1.n2 VDD1.t4 2.84533
R1475 VDD1.n2 VDD1.t0 2.84533
R1476 VDD1.n0 VDD1.t3 2.84533
R1477 VDD1.n0 VDD1.t2 2.84533
R1478 VDD1 VDD1.n3 0.571621
C0 VN VDD2 4.05425f
C1 VN VTAIL 4.57145f
C2 VDD1 VDD2 1.40307f
C3 VN VP 5.97881f
C4 VTAIL VDD1 5.8975f
C5 VTAIL VDD2 5.94943f
C6 VDD1 VP 4.35828f
C7 VP VDD2 0.457484f
C8 VTAIL VP 4.58566f
C9 VN VDD1 0.15114f
C10 VDD2 B 5.0913f
C11 VDD1 B 5.415564f
C12 VTAIL B 5.48963f
C13 VN B 12.31596f
C14 VP B 10.979522f
C15 VDD1.t5 B 1.32431f
C16 VDD1.t1 B 1.32347f
C17 VDD1.t3 B 0.122054f
C18 VDD1.t2 B 0.122054f
C19 VDD1.n0 B 1.0377f
C20 VDD1.n1 B 2.40842f
C21 VDD1.t4 B 0.122054f
C22 VDD1.t0 B 0.122054f
C23 VDD1.n2 B 1.03396f
C24 VDD1.n3 B 2.12943f
C25 VP.n0 B 0.034611f
C26 VP.t3 B 1.26279f
C27 VP.n1 B 0.04107f
C28 VP.n2 B 0.026254f
C29 VP.t2 B 1.26279f
C30 VP.n3 B 0.46614f
C31 VP.n4 B 0.026254f
C32 VP.n5 B 0.04107f
C33 VP.n6 B 0.034611f
C34 VP.t4 B 1.26279f
C35 VP.n7 B 0.034611f
C36 VP.t5 B 1.26279f
C37 VP.n8 B 0.04107f
C38 VP.n9 B 0.026254f
C39 VP.t1 B 1.26279f
C40 VP.n10 B 0.54115f
C41 VP.t0 B 1.47517f
C42 VP.n11 B 0.521638f
C43 VP.n12 B 0.253418f
C44 VP.n13 B 0.036668f
C45 VP.n14 B 0.048686f
C46 VP.n15 B 0.035259f
C47 VP.n16 B 0.026254f
C48 VP.n17 B 0.026254f
C49 VP.n18 B 0.026254f
C50 VP.n19 B 0.048686f
C51 VP.n20 B 0.032823f
C52 VP.n21 B 0.550897f
C53 VP.n22 B 1.23876f
C54 VP.n23 B 1.25988f
C55 VP.n24 B 0.550897f
C56 VP.n25 B 0.032823f
C57 VP.n26 B 0.048686f
C58 VP.n27 B 0.026254f
C59 VP.n28 B 0.026254f
C60 VP.n29 B 0.026254f
C61 VP.n30 B 0.035259f
C62 VP.n31 B 0.048686f
C63 VP.n32 B 0.036668f
C64 VP.n33 B 0.026254f
C65 VP.n34 B 0.026254f
C66 VP.n35 B 0.036668f
C67 VP.n36 B 0.048686f
C68 VP.n37 B 0.035259f
C69 VP.n38 B 0.026254f
C70 VP.n39 B 0.026254f
C71 VP.n40 B 0.026254f
C72 VP.n41 B 0.048686f
C73 VP.n42 B 0.032823f
C74 VP.n43 B 0.550897f
C75 VP.n44 B 0.043702f
C76 VTAIL.t10 B 0.144438f
C77 VTAIL.t7 B 0.144438f
C78 VTAIL.n0 B 1.14752f
C79 VTAIL.n1 B 0.4624f
C80 VTAIL.t0 B 1.46106f
C81 VTAIL.n2 B 0.697606f
C82 VTAIL.t1 B 0.144438f
C83 VTAIL.t5 B 0.144438f
C84 VTAIL.n3 B 1.14752f
C85 VTAIL.n4 B 1.76144f
C86 VTAIL.t8 B 0.144438f
C87 VTAIL.t11 B 0.144438f
C88 VTAIL.n5 B 1.14752f
C89 VTAIL.n6 B 1.76144f
C90 VTAIL.t6 B 1.46107f
C91 VTAIL.n7 B 0.6976f
C92 VTAIL.t3 B 0.144438f
C93 VTAIL.t4 B 0.144438f
C94 VTAIL.n8 B 1.14752f
C95 VTAIL.n9 B 0.617231f
C96 VTAIL.t2 B 1.46106f
C97 VTAIL.n10 B 1.62881f
C98 VTAIL.t9 B 1.46106f
C99 VTAIL.n11 B 1.57063f
C100 VDD2.t1 B 1.29523f
C101 VDD2.t4 B 0.119449f
C102 VDD2.t3 B 0.119449f
C103 VDD2.n0 B 1.01555f
C104 VDD2.n1 B 2.25337f
C105 VDD2.t5 B 1.28527f
C106 VDD2.n2 B 2.07991f
C107 VDD2.t2 B 0.119449f
C108 VDD2.t0 B 0.119449f
C109 VDD2.n3 B 1.01552f
C110 VN.n0 B 0.033836f
C111 VN.t2 B 1.2345f
C112 VN.n1 B 0.04015f
C113 VN.n2 B 0.025666f
C114 VN.t4 B 1.2345f
C115 VN.n3 B 0.529025f
C116 VN.t1 B 1.44212f
C117 VN.n4 B 0.50995f
C118 VN.n5 B 0.24774f
C119 VN.n6 B 0.035847f
C120 VN.n7 B 0.047595f
C121 VN.n8 B 0.034469f
C122 VN.n9 B 0.025666f
C123 VN.n10 B 0.025666f
C124 VN.n11 B 0.025666f
C125 VN.n12 B 0.047595f
C126 VN.n13 B 0.032087f
C127 VN.n14 B 0.538554f
C128 VN.n15 B 0.042723f
C129 VN.n16 B 0.033836f
C130 VN.t3 B 1.2345f
C131 VN.n17 B 0.04015f
C132 VN.n18 B 0.025666f
C133 VN.t0 B 1.2345f
C134 VN.n19 B 0.529025f
C135 VN.t5 B 1.44212f
C136 VN.n20 B 0.50995f
C137 VN.n21 B 0.24774f
C138 VN.n22 B 0.035847f
C139 VN.n23 B 0.047595f
C140 VN.n24 B 0.034469f
C141 VN.n25 B 0.025666f
C142 VN.n26 B 0.025666f
C143 VN.n27 B 0.025666f
C144 VN.n28 B 0.047595f
C145 VN.n29 B 0.032087f
C146 VN.n30 B 0.538554f
C147 VN.n31 B 1.22505f
.ends

