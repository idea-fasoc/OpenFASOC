* NGSPICE file created from diff_pair_sample_0412.ext - technology: sky130A

.subckt diff_pair_sample_0412 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=0 ps=0 w=17.75 l=1.08
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=6.9225 ps=36.28 w=17.75 l=1.08
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=6.9225 ps=36.28 w=17.75 l=1.08
X3 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=6.9225 ps=36.28 w=17.75 l=1.08
X4 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=6.9225 ps=36.28 w=17.75 l=1.08
X5 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=0 ps=0 w=17.75 l=1.08
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=0 ps=0 w=17.75 l=1.08
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9225 pd=36.28 as=0 ps=0 w=17.75 l=1.08
R0 B.n101 B.t6 599.529
R1 B.n98 B.t13 599.529
R2 B.n581 B.t2 599.529
R3 B.n418 B.t10 599.529
R4 B.n779 B.n778 585
R5 B.n780 B.n779 585
R6 B.n352 B.n97 585
R7 B.n351 B.n350 585
R8 B.n349 B.n348 585
R9 B.n347 B.n346 585
R10 B.n345 B.n344 585
R11 B.n343 B.n342 585
R12 B.n341 B.n340 585
R13 B.n339 B.n338 585
R14 B.n337 B.n336 585
R15 B.n335 B.n334 585
R16 B.n333 B.n332 585
R17 B.n331 B.n330 585
R18 B.n329 B.n328 585
R19 B.n327 B.n326 585
R20 B.n325 B.n324 585
R21 B.n323 B.n322 585
R22 B.n321 B.n320 585
R23 B.n319 B.n318 585
R24 B.n317 B.n316 585
R25 B.n315 B.n314 585
R26 B.n313 B.n312 585
R27 B.n311 B.n310 585
R28 B.n309 B.n308 585
R29 B.n307 B.n306 585
R30 B.n305 B.n304 585
R31 B.n303 B.n302 585
R32 B.n301 B.n300 585
R33 B.n299 B.n298 585
R34 B.n297 B.n296 585
R35 B.n295 B.n294 585
R36 B.n293 B.n292 585
R37 B.n291 B.n290 585
R38 B.n289 B.n288 585
R39 B.n287 B.n286 585
R40 B.n285 B.n284 585
R41 B.n283 B.n282 585
R42 B.n281 B.n280 585
R43 B.n279 B.n278 585
R44 B.n277 B.n276 585
R45 B.n275 B.n274 585
R46 B.n273 B.n272 585
R47 B.n271 B.n270 585
R48 B.n269 B.n268 585
R49 B.n267 B.n266 585
R50 B.n265 B.n264 585
R51 B.n263 B.n262 585
R52 B.n261 B.n260 585
R53 B.n259 B.n258 585
R54 B.n257 B.n256 585
R55 B.n255 B.n254 585
R56 B.n253 B.n252 585
R57 B.n251 B.n250 585
R58 B.n249 B.n248 585
R59 B.n247 B.n246 585
R60 B.n245 B.n244 585
R61 B.n243 B.n242 585
R62 B.n241 B.n240 585
R63 B.n239 B.n238 585
R64 B.n237 B.n236 585
R65 B.n235 B.n234 585
R66 B.n233 B.n232 585
R67 B.n231 B.n230 585
R68 B.n229 B.n228 585
R69 B.n227 B.n226 585
R70 B.n225 B.n224 585
R71 B.n223 B.n222 585
R72 B.n221 B.n220 585
R73 B.n218 B.n217 585
R74 B.n216 B.n215 585
R75 B.n214 B.n213 585
R76 B.n212 B.n211 585
R77 B.n210 B.n209 585
R78 B.n208 B.n207 585
R79 B.n206 B.n205 585
R80 B.n204 B.n203 585
R81 B.n202 B.n201 585
R82 B.n200 B.n199 585
R83 B.n198 B.n197 585
R84 B.n196 B.n195 585
R85 B.n194 B.n193 585
R86 B.n192 B.n191 585
R87 B.n190 B.n189 585
R88 B.n188 B.n187 585
R89 B.n186 B.n185 585
R90 B.n184 B.n183 585
R91 B.n182 B.n181 585
R92 B.n180 B.n179 585
R93 B.n178 B.n177 585
R94 B.n176 B.n175 585
R95 B.n174 B.n173 585
R96 B.n172 B.n171 585
R97 B.n170 B.n169 585
R98 B.n168 B.n167 585
R99 B.n166 B.n165 585
R100 B.n164 B.n163 585
R101 B.n162 B.n161 585
R102 B.n160 B.n159 585
R103 B.n158 B.n157 585
R104 B.n156 B.n155 585
R105 B.n154 B.n153 585
R106 B.n152 B.n151 585
R107 B.n150 B.n149 585
R108 B.n148 B.n147 585
R109 B.n146 B.n145 585
R110 B.n144 B.n143 585
R111 B.n142 B.n141 585
R112 B.n140 B.n139 585
R113 B.n138 B.n137 585
R114 B.n136 B.n135 585
R115 B.n134 B.n133 585
R116 B.n132 B.n131 585
R117 B.n130 B.n129 585
R118 B.n128 B.n127 585
R119 B.n126 B.n125 585
R120 B.n124 B.n123 585
R121 B.n122 B.n121 585
R122 B.n120 B.n119 585
R123 B.n118 B.n117 585
R124 B.n116 B.n115 585
R125 B.n114 B.n113 585
R126 B.n112 B.n111 585
R127 B.n110 B.n109 585
R128 B.n108 B.n107 585
R129 B.n106 B.n105 585
R130 B.n104 B.n103 585
R131 B.n32 B.n31 585
R132 B.n777 B.n33 585
R133 B.n781 B.n33 585
R134 B.n776 B.n775 585
R135 B.n775 B.n29 585
R136 B.n774 B.n28 585
R137 B.n787 B.n28 585
R138 B.n773 B.n27 585
R139 B.n788 B.n27 585
R140 B.n772 B.n26 585
R141 B.n789 B.n26 585
R142 B.n771 B.n770 585
R143 B.n770 B.n25 585
R144 B.n769 B.n21 585
R145 B.n795 B.n21 585
R146 B.n768 B.n20 585
R147 B.n796 B.n20 585
R148 B.n767 B.n19 585
R149 B.n797 B.n19 585
R150 B.n766 B.n765 585
R151 B.n765 B.n15 585
R152 B.n764 B.n14 585
R153 B.n803 B.n14 585
R154 B.n763 B.n13 585
R155 B.n804 B.n13 585
R156 B.n762 B.n12 585
R157 B.n805 B.n12 585
R158 B.n761 B.n760 585
R159 B.n760 B.n759 585
R160 B.n758 B.n757 585
R161 B.n758 B.n8 585
R162 B.n756 B.n7 585
R163 B.n812 B.n7 585
R164 B.n755 B.n6 585
R165 B.n813 B.n6 585
R166 B.n754 B.n5 585
R167 B.n814 B.n5 585
R168 B.n753 B.n752 585
R169 B.n752 B.n4 585
R170 B.n751 B.n353 585
R171 B.n751 B.n750 585
R172 B.n741 B.n354 585
R173 B.n355 B.n354 585
R174 B.n743 B.n742 585
R175 B.n744 B.n743 585
R176 B.n740 B.n360 585
R177 B.n360 B.n359 585
R178 B.n739 B.n738 585
R179 B.n738 B.n737 585
R180 B.n362 B.n361 585
R181 B.n363 B.n362 585
R182 B.n730 B.n729 585
R183 B.n731 B.n730 585
R184 B.n728 B.n368 585
R185 B.n368 B.n367 585
R186 B.n727 B.n726 585
R187 B.n726 B.n725 585
R188 B.n370 B.n369 585
R189 B.n718 B.n370 585
R190 B.n717 B.n716 585
R191 B.n719 B.n717 585
R192 B.n715 B.n375 585
R193 B.n375 B.n374 585
R194 B.n714 B.n713 585
R195 B.n713 B.n712 585
R196 B.n377 B.n376 585
R197 B.n378 B.n377 585
R198 B.n705 B.n704 585
R199 B.n706 B.n705 585
R200 B.n381 B.n380 585
R201 B.n450 B.n449 585
R202 B.n451 B.n447 585
R203 B.n447 B.n382 585
R204 B.n453 B.n452 585
R205 B.n455 B.n446 585
R206 B.n458 B.n457 585
R207 B.n459 B.n445 585
R208 B.n461 B.n460 585
R209 B.n463 B.n444 585
R210 B.n466 B.n465 585
R211 B.n467 B.n443 585
R212 B.n469 B.n468 585
R213 B.n471 B.n442 585
R214 B.n474 B.n473 585
R215 B.n475 B.n441 585
R216 B.n477 B.n476 585
R217 B.n479 B.n440 585
R218 B.n482 B.n481 585
R219 B.n483 B.n439 585
R220 B.n485 B.n484 585
R221 B.n487 B.n438 585
R222 B.n490 B.n489 585
R223 B.n491 B.n437 585
R224 B.n493 B.n492 585
R225 B.n495 B.n436 585
R226 B.n498 B.n497 585
R227 B.n499 B.n435 585
R228 B.n501 B.n500 585
R229 B.n503 B.n434 585
R230 B.n506 B.n505 585
R231 B.n507 B.n433 585
R232 B.n509 B.n508 585
R233 B.n511 B.n432 585
R234 B.n514 B.n513 585
R235 B.n515 B.n431 585
R236 B.n517 B.n516 585
R237 B.n519 B.n430 585
R238 B.n522 B.n521 585
R239 B.n523 B.n429 585
R240 B.n525 B.n524 585
R241 B.n527 B.n428 585
R242 B.n530 B.n529 585
R243 B.n531 B.n427 585
R244 B.n533 B.n532 585
R245 B.n535 B.n426 585
R246 B.n538 B.n537 585
R247 B.n539 B.n425 585
R248 B.n541 B.n540 585
R249 B.n543 B.n424 585
R250 B.n546 B.n545 585
R251 B.n547 B.n423 585
R252 B.n549 B.n548 585
R253 B.n551 B.n422 585
R254 B.n554 B.n553 585
R255 B.n555 B.n421 585
R256 B.n557 B.n556 585
R257 B.n559 B.n420 585
R258 B.n562 B.n561 585
R259 B.n563 B.n417 585
R260 B.n566 B.n565 585
R261 B.n568 B.n416 585
R262 B.n571 B.n570 585
R263 B.n572 B.n415 585
R264 B.n574 B.n573 585
R265 B.n576 B.n414 585
R266 B.n579 B.n578 585
R267 B.n580 B.n413 585
R268 B.n585 B.n584 585
R269 B.n587 B.n412 585
R270 B.n590 B.n589 585
R271 B.n591 B.n411 585
R272 B.n593 B.n592 585
R273 B.n595 B.n410 585
R274 B.n598 B.n597 585
R275 B.n599 B.n409 585
R276 B.n601 B.n600 585
R277 B.n603 B.n408 585
R278 B.n606 B.n605 585
R279 B.n607 B.n407 585
R280 B.n609 B.n608 585
R281 B.n611 B.n406 585
R282 B.n614 B.n613 585
R283 B.n615 B.n405 585
R284 B.n617 B.n616 585
R285 B.n619 B.n404 585
R286 B.n622 B.n621 585
R287 B.n623 B.n403 585
R288 B.n625 B.n624 585
R289 B.n627 B.n402 585
R290 B.n630 B.n629 585
R291 B.n631 B.n401 585
R292 B.n633 B.n632 585
R293 B.n635 B.n400 585
R294 B.n638 B.n637 585
R295 B.n639 B.n399 585
R296 B.n641 B.n640 585
R297 B.n643 B.n398 585
R298 B.n646 B.n645 585
R299 B.n647 B.n397 585
R300 B.n649 B.n648 585
R301 B.n651 B.n396 585
R302 B.n654 B.n653 585
R303 B.n655 B.n395 585
R304 B.n657 B.n656 585
R305 B.n659 B.n394 585
R306 B.n662 B.n661 585
R307 B.n663 B.n393 585
R308 B.n665 B.n664 585
R309 B.n667 B.n392 585
R310 B.n670 B.n669 585
R311 B.n671 B.n391 585
R312 B.n673 B.n672 585
R313 B.n675 B.n390 585
R314 B.n678 B.n677 585
R315 B.n679 B.n389 585
R316 B.n681 B.n680 585
R317 B.n683 B.n388 585
R318 B.n686 B.n685 585
R319 B.n687 B.n387 585
R320 B.n689 B.n688 585
R321 B.n691 B.n386 585
R322 B.n694 B.n693 585
R323 B.n695 B.n385 585
R324 B.n697 B.n696 585
R325 B.n699 B.n384 585
R326 B.n702 B.n701 585
R327 B.n703 B.n383 585
R328 B.n708 B.n707 585
R329 B.n707 B.n706 585
R330 B.n709 B.n379 585
R331 B.n379 B.n378 585
R332 B.n711 B.n710 585
R333 B.n712 B.n711 585
R334 B.n373 B.n372 585
R335 B.n374 B.n373 585
R336 B.n721 B.n720 585
R337 B.n720 B.n719 585
R338 B.n722 B.n371 585
R339 B.n718 B.n371 585
R340 B.n724 B.n723 585
R341 B.n725 B.n724 585
R342 B.n366 B.n365 585
R343 B.n367 B.n366 585
R344 B.n733 B.n732 585
R345 B.n732 B.n731 585
R346 B.n734 B.n364 585
R347 B.n364 B.n363 585
R348 B.n736 B.n735 585
R349 B.n737 B.n736 585
R350 B.n358 B.n357 585
R351 B.n359 B.n358 585
R352 B.n746 B.n745 585
R353 B.n745 B.n744 585
R354 B.n747 B.n356 585
R355 B.n356 B.n355 585
R356 B.n749 B.n748 585
R357 B.n750 B.n749 585
R358 B.n3 B.n0 585
R359 B.n4 B.n3 585
R360 B.n811 B.n1 585
R361 B.n812 B.n811 585
R362 B.n810 B.n809 585
R363 B.n810 B.n8 585
R364 B.n808 B.n9 585
R365 B.n759 B.n9 585
R366 B.n807 B.n806 585
R367 B.n806 B.n805 585
R368 B.n11 B.n10 585
R369 B.n804 B.n11 585
R370 B.n802 B.n801 585
R371 B.n803 B.n802 585
R372 B.n800 B.n16 585
R373 B.n16 B.n15 585
R374 B.n799 B.n798 585
R375 B.n798 B.n797 585
R376 B.n18 B.n17 585
R377 B.n796 B.n18 585
R378 B.n794 B.n793 585
R379 B.n795 B.n794 585
R380 B.n792 B.n22 585
R381 B.n25 B.n22 585
R382 B.n791 B.n790 585
R383 B.n790 B.n789 585
R384 B.n24 B.n23 585
R385 B.n788 B.n24 585
R386 B.n786 B.n785 585
R387 B.n787 B.n786 585
R388 B.n784 B.n30 585
R389 B.n30 B.n29 585
R390 B.n783 B.n782 585
R391 B.n782 B.n781 585
R392 B.n815 B.n814 585
R393 B.n813 B.n2 585
R394 B.n782 B.n32 463.671
R395 B.n779 B.n33 463.671
R396 B.n705 B.n383 463.671
R397 B.n707 B.n381 463.671
R398 B.n780 B.n96 256.663
R399 B.n780 B.n95 256.663
R400 B.n780 B.n94 256.663
R401 B.n780 B.n93 256.663
R402 B.n780 B.n92 256.663
R403 B.n780 B.n91 256.663
R404 B.n780 B.n90 256.663
R405 B.n780 B.n89 256.663
R406 B.n780 B.n88 256.663
R407 B.n780 B.n87 256.663
R408 B.n780 B.n86 256.663
R409 B.n780 B.n85 256.663
R410 B.n780 B.n84 256.663
R411 B.n780 B.n83 256.663
R412 B.n780 B.n82 256.663
R413 B.n780 B.n81 256.663
R414 B.n780 B.n80 256.663
R415 B.n780 B.n79 256.663
R416 B.n780 B.n78 256.663
R417 B.n780 B.n77 256.663
R418 B.n780 B.n76 256.663
R419 B.n780 B.n75 256.663
R420 B.n780 B.n74 256.663
R421 B.n780 B.n73 256.663
R422 B.n780 B.n72 256.663
R423 B.n780 B.n71 256.663
R424 B.n780 B.n70 256.663
R425 B.n780 B.n69 256.663
R426 B.n780 B.n68 256.663
R427 B.n780 B.n67 256.663
R428 B.n780 B.n66 256.663
R429 B.n780 B.n65 256.663
R430 B.n780 B.n64 256.663
R431 B.n780 B.n63 256.663
R432 B.n780 B.n62 256.663
R433 B.n780 B.n61 256.663
R434 B.n780 B.n60 256.663
R435 B.n780 B.n59 256.663
R436 B.n780 B.n58 256.663
R437 B.n780 B.n57 256.663
R438 B.n780 B.n56 256.663
R439 B.n780 B.n55 256.663
R440 B.n780 B.n54 256.663
R441 B.n780 B.n53 256.663
R442 B.n780 B.n52 256.663
R443 B.n780 B.n51 256.663
R444 B.n780 B.n50 256.663
R445 B.n780 B.n49 256.663
R446 B.n780 B.n48 256.663
R447 B.n780 B.n47 256.663
R448 B.n780 B.n46 256.663
R449 B.n780 B.n45 256.663
R450 B.n780 B.n44 256.663
R451 B.n780 B.n43 256.663
R452 B.n780 B.n42 256.663
R453 B.n780 B.n41 256.663
R454 B.n780 B.n40 256.663
R455 B.n780 B.n39 256.663
R456 B.n780 B.n38 256.663
R457 B.n780 B.n37 256.663
R458 B.n780 B.n36 256.663
R459 B.n780 B.n35 256.663
R460 B.n780 B.n34 256.663
R461 B.n448 B.n382 256.663
R462 B.n454 B.n382 256.663
R463 B.n456 B.n382 256.663
R464 B.n462 B.n382 256.663
R465 B.n464 B.n382 256.663
R466 B.n470 B.n382 256.663
R467 B.n472 B.n382 256.663
R468 B.n478 B.n382 256.663
R469 B.n480 B.n382 256.663
R470 B.n486 B.n382 256.663
R471 B.n488 B.n382 256.663
R472 B.n494 B.n382 256.663
R473 B.n496 B.n382 256.663
R474 B.n502 B.n382 256.663
R475 B.n504 B.n382 256.663
R476 B.n510 B.n382 256.663
R477 B.n512 B.n382 256.663
R478 B.n518 B.n382 256.663
R479 B.n520 B.n382 256.663
R480 B.n526 B.n382 256.663
R481 B.n528 B.n382 256.663
R482 B.n534 B.n382 256.663
R483 B.n536 B.n382 256.663
R484 B.n542 B.n382 256.663
R485 B.n544 B.n382 256.663
R486 B.n550 B.n382 256.663
R487 B.n552 B.n382 256.663
R488 B.n558 B.n382 256.663
R489 B.n560 B.n382 256.663
R490 B.n567 B.n382 256.663
R491 B.n569 B.n382 256.663
R492 B.n575 B.n382 256.663
R493 B.n577 B.n382 256.663
R494 B.n586 B.n382 256.663
R495 B.n588 B.n382 256.663
R496 B.n594 B.n382 256.663
R497 B.n596 B.n382 256.663
R498 B.n602 B.n382 256.663
R499 B.n604 B.n382 256.663
R500 B.n610 B.n382 256.663
R501 B.n612 B.n382 256.663
R502 B.n618 B.n382 256.663
R503 B.n620 B.n382 256.663
R504 B.n626 B.n382 256.663
R505 B.n628 B.n382 256.663
R506 B.n634 B.n382 256.663
R507 B.n636 B.n382 256.663
R508 B.n642 B.n382 256.663
R509 B.n644 B.n382 256.663
R510 B.n650 B.n382 256.663
R511 B.n652 B.n382 256.663
R512 B.n658 B.n382 256.663
R513 B.n660 B.n382 256.663
R514 B.n666 B.n382 256.663
R515 B.n668 B.n382 256.663
R516 B.n674 B.n382 256.663
R517 B.n676 B.n382 256.663
R518 B.n682 B.n382 256.663
R519 B.n684 B.n382 256.663
R520 B.n690 B.n382 256.663
R521 B.n692 B.n382 256.663
R522 B.n698 B.n382 256.663
R523 B.n700 B.n382 256.663
R524 B.n817 B.n816 256.663
R525 B.n105 B.n104 163.367
R526 B.n109 B.n108 163.367
R527 B.n113 B.n112 163.367
R528 B.n117 B.n116 163.367
R529 B.n121 B.n120 163.367
R530 B.n125 B.n124 163.367
R531 B.n129 B.n128 163.367
R532 B.n133 B.n132 163.367
R533 B.n137 B.n136 163.367
R534 B.n141 B.n140 163.367
R535 B.n145 B.n144 163.367
R536 B.n149 B.n148 163.367
R537 B.n153 B.n152 163.367
R538 B.n157 B.n156 163.367
R539 B.n161 B.n160 163.367
R540 B.n165 B.n164 163.367
R541 B.n169 B.n168 163.367
R542 B.n173 B.n172 163.367
R543 B.n177 B.n176 163.367
R544 B.n181 B.n180 163.367
R545 B.n185 B.n184 163.367
R546 B.n189 B.n188 163.367
R547 B.n193 B.n192 163.367
R548 B.n197 B.n196 163.367
R549 B.n201 B.n200 163.367
R550 B.n205 B.n204 163.367
R551 B.n209 B.n208 163.367
R552 B.n213 B.n212 163.367
R553 B.n217 B.n216 163.367
R554 B.n222 B.n221 163.367
R555 B.n226 B.n225 163.367
R556 B.n230 B.n229 163.367
R557 B.n234 B.n233 163.367
R558 B.n238 B.n237 163.367
R559 B.n242 B.n241 163.367
R560 B.n246 B.n245 163.367
R561 B.n250 B.n249 163.367
R562 B.n254 B.n253 163.367
R563 B.n258 B.n257 163.367
R564 B.n262 B.n261 163.367
R565 B.n266 B.n265 163.367
R566 B.n270 B.n269 163.367
R567 B.n274 B.n273 163.367
R568 B.n278 B.n277 163.367
R569 B.n282 B.n281 163.367
R570 B.n286 B.n285 163.367
R571 B.n290 B.n289 163.367
R572 B.n294 B.n293 163.367
R573 B.n298 B.n297 163.367
R574 B.n302 B.n301 163.367
R575 B.n306 B.n305 163.367
R576 B.n310 B.n309 163.367
R577 B.n314 B.n313 163.367
R578 B.n318 B.n317 163.367
R579 B.n322 B.n321 163.367
R580 B.n326 B.n325 163.367
R581 B.n330 B.n329 163.367
R582 B.n334 B.n333 163.367
R583 B.n338 B.n337 163.367
R584 B.n342 B.n341 163.367
R585 B.n346 B.n345 163.367
R586 B.n350 B.n349 163.367
R587 B.n779 B.n97 163.367
R588 B.n705 B.n377 163.367
R589 B.n713 B.n377 163.367
R590 B.n713 B.n375 163.367
R591 B.n717 B.n375 163.367
R592 B.n717 B.n370 163.367
R593 B.n726 B.n370 163.367
R594 B.n726 B.n368 163.367
R595 B.n730 B.n368 163.367
R596 B.n730 B.n362 163.367
R597 B.n738 B.n362 163.367
R598 B.n738 B.n360 163.367
R599 B.n743 B.n360 163.367
R600 B.n743 B.n354 163.367
R601 B.n751 B.n354 163.367
R602 B.n752 B.n751 163.367
R603 B.n752 B.n5 163.367
R604 B.n6 B.n5 163.367
R605 B.n7 B.n6 163.367
R606 B.n758 B.n7 163.367
R607 B.n760 B.n758 163.367
R608 B.n760 B.n12 163.367
R609 B.n13 B.n12 163.367
R610 B.n14 B.n13 163.367
R611 B.n765 B.n14 163.367
R612 B.n765 B.n19 163.367
R613 B.n20 B.n19 163.367
R614 B.n21 B.n20 163.367
R615 B.n770 B.n21 163.367
R616 B.n770 B.n26 163.367
R617 B.n27 B.n26 163.367
R618 B.n28 B.n27 163.367
R619 B.n775 B.n28 163.367
R620 B.n775 B.n33 163.367
R621 B.n449 B.n447 163.367
R622 B.n453 B.n447 163.367
R623 B.n457 B.n455 163.367
R624 B.n461 B.n445 163.367
R625 B.n465 B.n463 163.367
R626 B.n469 B.n443 163.367
R627 B.n473 B.n471 163.367
R628 B.n477 B.n441 163.367
R629 B.n481 B.n479 163.367
R630 B.n485 B.n439 163.367
R631 B.n489 B.n487 163.367
R632 B.n493 B.n437 163.367
R633 B.n497 B.n495 163.367
R634 B.n501 B.n435 163.367
R635 B.n505 B.n503 163.367
R636 B.n509 B.n433 163.367
R637 B.n513 B.n511 163.367
R638 B.n517 B.n431 163.367
R639 B.n521 B.n519 163.367
R640 B.n525 B.n429 163.367
R641 B.n529 B.n527 163.367
R642 B.n533 B.n427 163.367
R643 B.n537 B.n535 163.367
R644 B.n541 B.n425 163.367
R645 B.n545 B.n543 163.367
R646 B.n549 B.n423 163.367
R647 B.n553 B.n551 163.367
R648 B.n557 B.n421 163.367
R649 B.n561 B.n559 163.367
R650 B.n566 B.n417 163.367
R651 B.n570 B.n568 163.367
R652 B.n574 B.n415 163.367
R653 B.n578 B.n576 163.367
R654 B.n585 B.n413 163.367
R655 B.n589 B.n587 163.367
R656 B.n593 B.n411 163.367
R657 B.n597 B.n595 163.367
R658 B.n601 B.n409 163.367
R659 B.n605 B.n603 163.367
R660 B.n609 B.n407 163.367
R661 B.n613 B.n611 163.367
R662 B.n617 B.n405 163.367
R663 B.n621 B.n619 163.367
R664 B.n625 B.n403 163.367
R665 B.n629 B.n627 163.367
R666 B.n633 B.n401 163.367
R667 B.n637 B.n635 163.367
R668 B.n641 B.n399 163.367
R669 B.n645 B.n643 163.367
R670 B.n649 B.n397 163.367
R671 B.n653 B.n651 163.367
R672 B.n657 B.n395 163.367
R673 B.n661 B.n659 163.367
R674 B.n665 B.n393 163.367
R675 B.n669 B.n667 163.367
R676 B.n673 B.n391 163.367
R677 B.n677 B.n675 163.367
R678 B.n681 B.n389 163.367
R679 B.n685 B.n683 163.367
R680 B.n689 B.n387 163.367
R681 B.n693 B.n691 163.367
R682 B.n697 B.n385 163.367
R683 B.n701 B.n699 163.367
R684 B.n707 B.n379 163.367
R685 B.n711 B.n379 163.367
R686 B.n711 B.n373 163.367
R687 B.n720 B.n373 163.367
R688 B.n720 B.n371 163.367
R689 B.n724 B.n371 163.367
R690 B.n724 B.n366 163.367
R691 B.n732 B.n366 163.367
R692 B.n732 B.n364 163.367
R693 B.n736 B.n364 163.367
R694 B.n736 B.n358 163.367
R695 B.n745 B.n358 163.367
R696 B.n745 B.n356 163.367
R697 B.n749 B.n356 163.367
R698 B.n749 B.n3 163.367
R699 B.n815 B.n3 163.367
R700 B.n811 B.n2 163.367
R701 B.n811 B.n810 163.367
R702 B.n810 B.n9 163.367
R703 B.n806 B.n9 163.367
R704 B.n806 B.n11 163.367
R705 B.n802 B.n11 163.367
R706 B.n802 B.n16 163.367
R707 B.n798 B.n16 163.367
R708 B.n798 B.n18 163.367
R709 B.n794 B.n18 163.367
R710 B.n794 B.n22 163.367
R711 B.n790 B.n22 163.367
R712 B.n790 B.n24 163.367
R713 B.n786 B.n24 163.367
R714 B.n786 B.n30 163.367
R715 B.n782 B.n30 163.367
R716 B.n98 B.t14 95.9669
R717 B.n581 B.t5 95.9669
R718 B.n101 B.t8 95.9432
R719 B.n418 B.t12 95.9432
R720 B.n34 B.n32 71.676
R721 B.n105 B.n35 71.676
R722 B.n109 B.n36 71.676
R723 B.n113 B.n37 71.676
R724 B.n117 B.n38 71.676
R725 B.n121 B.n39 71.676
R726 B.n125 B.n40 71.676
R727 B.n129 B.n41 71.676
R728 B.n133 B.n42 71.676
R729 B.n137 B.n43 71.676
R730 B.n141 B.n44 71.676
R731 B.n145 B.n45 71.676
R732 B.n149 B.n46 71.676
R733 B.n153 B.n47 71.676
R734 B.n157 B.n48 71.676
R735 B.n161 B.n49 71.676
R736 B.n165 B.n50 71.676
R737 B.n169 B.n51 71.676
R738 B.n173 B.n52 71.676
R739 B.n177 B.n53 71.676
R740 B.n181 B.n54 71.676
R741 B.n185 B.n55 71.676
R742 B.n189 B.n56 71.676
R743 B.n193 B.n57 71.676
R744 B.n197 B.n58 71.676
R745 B.n201 B.n59 71.676
R746 B.n205 B.n60 71.676
R747 B.n209 B.n61 71.676
R748 B.n213 B.n62 71.676
R749 B.n217 B.n63 71.676
R750 B.n222 B.n64 71.676
R751 B.n226 B.n65 71.676
R752 B.n230 B.n66 71.676
R753 B.n234 B.n67 71.676
R754 B.n238 B.n68 71.676
R755 B.n242 B.n69 71.676
R756 B.n246 B.n70 71.676
R757 B.n250 B.n71 71.676
R758 B.n254 B.n72 71.676
R759 B.n258 B.n73 71.676
R760 B.n262 B.n74 71.676
R761 B.n266 B.n75 71.676
R762 B.n270 B.n76 71.676
R763 B.n274 B.n77 71.676
R764 B.n278 B.n78 71.676
R765 B.n282 B.n79 71.676
R766 B.n286 B.n80 71.676
R767 B.n290 B.n81 71.676
R768 B.n294 B.n82 71.676
R769 B.n298 B.n83 71.676
R770 B.n302 B.n84 71.676
R771 B.n306 B.n85 71.676
R772 B.n310 B.n86 71.676
R773 B.n314 B.n87 71.676
R774 B.n318 B.n88 71.676
R775 B.n322 B.n89 71.676
R776 B.n326 B.n90 71.676
R777 B.n330 B.n91 71.676
R778 B.n334 B.n92 71.676
R779 B.n338 B.n93 71.676
R780 B.n342 B.n94 71.676
R781 B.n346 B.n95 71.676
R782 B.n350 B.n96 71.676
R783 B.n97 B.n96 71.676
R784 B.n349 B.n95 71.676
R785 B.n345 B.n94 71.676
R786 B.n341 B.n93 71.676
R787 B.n337 B.n92 71.676
R788 B.n333 B.n91 71.676
R789 B.n329 B.n90 71.676
R790 B.n325 B.n89 71.676
R791 B.n321 B.n88 71.676
R792 B.n317 B.n87 71.676
R793 B.n313 B.n86 71.676
R794 B.n309 B.n85 71.676
R795 B.n305 B.n84 71.676
R796 B.n301 B.n83 71.676
R797 B.n297 B.n82 71.676
R798 B.n293 B.n81 71.676
R799 B.n289 B.n80 71.676
R800 B.n285 B.n79 71.676
R801 B.n281 B.n78 71.676
R802 B.n277 B.n77 71.676
R803 B.n273 B.n76 71.676
R804 B.n269 B.n75 71.676
R805 B.n265 B.n74 71.676
R806 B.n261 B.n73 71.676
R807 B.n257 B.n72 71.676
R808 B.n253 B.n71 71.676
R809 B.n249 B.n70 71.676
R810 B.n245 B.n69 71.676
R811 B.n241 B.n68 71.676
R812 B.n237 B.n67 71.676
R813 B.n233 B.n66 71.676
R814 B.n229 B.n65 71.676
R815 B.n225 B.n64 71.676
R816 B.n221 B.n63 71.676
R817 B.n216 B.n62 71.676
R818 B.n212 B.n61 71.676
R819 B.n208 B.n60 71.676
R820 B.n204 B.n59 71.676
R821 B.n200 B.n58 71.676
R822 B.n196 B.n57 71.676
R823 B.n192 B.n56 71.676
R824 B.n188 B.n55 71.676
R825 B.n184 B.n54 71.676
R826 B.n180 B.n53 71.676
R827 B.n176 B.n52 71.676
R828 B.n172 B.n51 71.676
R829 B.n168 B.n50 71.676
R830 B.n164 B.n49 71.676
R831 B.n160 B.n48 71.676
R832 B.n156 B.n47 71.676
R833 B.n152 B.n46 71.676
R834 B.n148 B.n45 71.676
R835 B.n144 B.n44 71.676
R836 B.n140 B.n43 71.676
R837 B.n136 B.n42 71.676
R838 B.n132 B.n41 71.676
R839 B.n128 B.n40 71.676
R840 B.n124 B.n39 71.676
R841 B.n120 B.n38 71.676
R842 B.n116 B.n37 71.676
R843 B.n112 B.n36 71.676
R844 B.n108 B.n35 71.676
R845 B.n104 B.n34 71.676
R846 B.n448 B.n381 71.676
R847 B.n454 B.n453 71.676
R848 B.n457 B.n456 71.676
R849 B.n462 B.n461 71.676
R850 B.n465 B.n464 71.676
R851 B.n470 B.n469 71.676
R852 B.n473 B.n472 71.676
R853 B.n478 B.n477 71.676
R854 B.n481 B.n480 71.676
R855 B.n486 B.n485 71.676
R856 B.n489 B.n488 71.676
R857 B.n494 B.n493 71.676
R858 B.n497 B.n496 71.676
R859 B.n502 B.n501 71.676
R860 B.n505 B.n504 71.676
R861 B.n510 B.n509 71.676
R862 B.n513 B.n512 71.676
R863 B.n518 B.n517 71.676
R864 B.n521 B.n520 71.676
R865 B.n526 B.n525 71.676
R866 B.n529 B.n528 71.676
R867 B.n534 B.n533 71.676
R868 B.n537 B.n536 71.676
R869 B.n542 B.n541 71.676
R870 B.n545 B.n544 71.676
R871 B.n550 B.n549 71.676
R872 B.n553 B.n552 71.676
R873 B.n558 B.n557 71.676
R874 B.n561 B.n560 71.676
R875 B.n567 B.n566 71.676
R876 B.n570 B.n569 71.676
R877 B.n575 B.n574 71.676
R878 B.n578 B.n577 71.676
R879 B.n586 B.n585 71.676
R880 B.n589 B.n588 71.676
R881 B.n594 B.n593 71.676
R882 B.n597 B.n596 71.676
R883 B.n602 B.n601 71.676
R884 B.n605 B.n604 71.676
R885 B.n610 B.n609 71.676
R886 B.n613 B.n612 71.676
R887 B.n618 B.n617 71.676
R888 B.n621 B.n620 71.676
R889 B.n626 B.n625 71.676
R890 B.n629 B.n628 71.676
R891 B.n634 B.n633 71.676
R892 B.n637 B.n636 71.676
R893 B.n642 B.n641 71.676
R894 B.n645 B.n644 71.676
R895 B.n650 B.n649 71.676
R896 B.n653 B.n652 71.676
R897 B.n658 B.n657 71.676
R898 B.n661 B.n660 71.676
R899 B.n666 B.n665 71.676
R900 B.n669 B.n668 71.676
R901 B.n674 B.n673 71.676
R902 B.n677 B.n676 71.676
R903 B.n682 B.n681 71.676
R904 B.n685 B.n684 71.676
R905 B.n690 B.n689 71.676
R906 B.n693 B.n692 71.676
R907 B.n698 B.n697 71.676
R908 B.n701 B.n700 71.676
R909 B.n449 B.n448 71.676
R910 B.n455 B.n454 71.676
R911 B.n456 B.n445 71.676
R912 B.n463 B.n462 71.676
R913 B.n464 B.n443 71.676
R914 B.n471 B.n470 71.676
R915 B.n472 B.n441 71.676
R916 B.n479 B.n478 71.676
R917 B.n480 B.n439 71.676
R918 B.n487 B.n486 71.676
R919 B.n488 B.n437 71.676
R920 B.n495 B.n494 71.676
R921 B.n496 B.n435 71.676
R922 B.n503 B.n502 71.676
R923 B.n504 B.n433 71.676
R924 B.n511 B.n510 71.676
R925 B.n512 B.n431 71.676
R926 B.n519 B.n518 71.676
R927 B.n520 B.n429 71.676
R928 B.n527 B.n526 71.676
R929 B.n528 B.n427 71.676
R930 B.n535 B.n534 71.676
R931 B.n536 B.n425 71.676
R932 B.n543 B.n542 71.676
R933 B.n544 B.n423 71.676
R934 B.n551 B.n550 71.676
R935 B.n552 B.n421 71.676
R936 B.n559 B.n558 71.676
R937 B.n560 B.n417 71.676
R938 B.n568 B.n567 71.676
R939 B.n569 B.n415 71.676
R940 B.n576 B.n575 71.676
R941 B.n577 B.n413 71.676
R942 B.n587 B.n586 71.676
R943 B.n588 B.n411 71.676
R944 B.n595 B.n594 71.676
R945 B.n596 B.n409 71.676
R946 B.n603 B.n602 71.676
R947 B.n604 B.n407 71.676
R948 B.n611 B.n610 71.676
R949 B.n612 B.n405 71.676
R950 B.n619 B.n618 71.676
R951 B.n620 B.n403 71.676
R952 B.n627 B.n626 71.676
R953 B.n628 B.n401 71.676
R954 B.n635 B.n634 71.676
R955 B.n636 B.n399 71.676
R956 B.n643 B.n642 71.676
R957 B.n644 B.n397 71.676
R958 B.n651 B.n650 71.676
R959 B.n652 B.n395 71.676
R960 B.n659 B.n658 71.676
R961 B.n660 B.n393 71.676
R962 B.n667 B.n666 71.676
R963 B.n668 B.n391 71.676
R964 B.n675 B.n674 71.676
R965 B.n676 B.n389 71.676
R966 B.n683 B.n682 71.676
R967 B.n684 B.n387 71.676
R968 B.n691 B.n690 71.676
R969 B.n692 B.n385 71.676
R970 B.n699 B.n698 71.676
R971 B.n700 B.n383 71.676
R972 B.n816 B.n815 71.676
R973 B.n816 B.n2 71.676
R974 B.n99 B.t15 68.6215
R975 B.n582 B.t4 68.6215
R976 B.n102 B.t9 68.5977
R977 B.n419 B.t11 68.5977
R978 B.n219 B.n102 59.5399
R979 B.n100 B.n99 59.5399
R980 B.n583 B.n582 59.5399
R981 B.n564 B.n419 59.5399
R982 B.n706 B.n382 55.8478
R983 B.n781 B.n780 55.8478
R984 B.n706 B.n378 32.4587
R985 B.n712 B.n378 32.4587
R986 B.n712 B.n374 32.4587
R987 B.n719 B.n374 32.4587
R988 B.n719 B.n718 32.4587
R989 B.n725 B.n367 32.4587
R990 B.n731 B.n367 32.4587
R991 B.n731 B.n363 32.4587
R992 B.n737 B.n363 32.4587
R993 B.n737 B.n359 32.4587
R994 B.n744 B.n359 32.4587
R995 B.n750 B.n355 32.4587
R996 B.n750 B.n4 32.4587
R997 B.n814 B.n4 32.4587
R998 B.n814 B.n813 32.4587
R999 B.n813 B.n812 32.4587
R1000 B.n812 B.n8 32.4587
R1001 B.n759 B.n8 32.4587
R1002 B.n805 B.n804 32.4587
R1003 B.n804 B.n803 32.4587
R1004 B.n803 B.n15 32.4587
R1005 B.n797 B.n15 32.4587
R1006 B.n797 B.n796 32.4587
R1007 B.n796 B.n795 32.4587
R1008 B.n789 B.n25 32.4587
R1009 B.n789 B.n788 32.4587
R1010 B.n788 B.n787 32.4587
R1011 B.n787 B.n29 32.4587
R1012 B.n781 B.n29 32.4587
R1013 B.n708 B.n380 30.1273
R1014 B.n704 B.n703 30.1273
R1015 B.n778 B.n777 30.1273
R1016 B.n783 B.n31 30.1273
R1017 B.n102 B.n101 27.346
R1018 B.n99 B.n98 27.346
R1019 B.n582 B.n581 27.346
R1020 B.n419 B.n418 27.346
R1021 B.n744 B.t1 26.7308
R1022 B.n805 B.t0 26.7308
R1023 B B.n817 18.0485
R1024 B.n725 B.t3 17.1843
R1025 B.n795 B.t7 17.1843
R1026 B.n718 B.t3 15.275
R1027 B.n25 B.t7 15.275
R1028 B.n709 B.n708 10.6151
R1029 B.n710 B.n709 10.6151
R1030 B.n710 B.n372 10.6151
R1031 B.n721 B.n372 10.6151
R1032 B.n722 B.n721 10.6151
R1033 B.n723 B.n722 10.6151
R1034 B.n723 B.n365 10.6151
R1035 B.n733 B.n365 10.6151
R1036 B.n734 B.n733 10.6151
R1037 B.n735 B.n734 10.6151
R1038 B.n735 B.n357 10.6151
R1039 B.n746 B.n357 10.6151
R1040 B.n747 B.n746 10.6151
R1041 B.n748 B.n747 10.6151
R1042 B.n748 B.n0 10.6151
R1043 B.n450 B.n380 10.6151
R1044 B.n451 B.n450 10.6151
R1045 B.n452 B.n451 10.6151
R1046 B.n452 B.n446 10.6151
R1047 B.n458 B.n446 10.6151
R1048 B.n459 B.n458 10.6151
R1049 B.n460 B.n459 10.6151
R1050 B.n460 B.n444 10.6151
R1051 B.n466 B.n444 10.6151
R1052 B.n467 B.n466 10.6151
R1053 B.n468 B.n467 10.6151
R1054 B.n468 B.n442 10.6151
R1055 B.n474 B.n442 10.6151
R1056 B.n475 B.n474 10.6151
R1057 B.n476 B.n475 10.6151
R1058 B.n476 B.n440 10.6151
R1059 B.n482 B.n440 10.6151
R1060 B.n483 B.n482 10.6151
R1061 B.n484 B.n483 10.6151
R1062 B.n484 B.n438 10.6151
R1063 B.n490 B.n438 10.6151
R1064 B.n491 B.n490 10.6151
R1065 B.n492 B.n491 10.6151
R1066 B.n492 B.n436 10.6151
R1067 B.n498 B.n436 10.6151
R1068 B.n499 B.n498 10.6151
R1069 B.n500 B.n499 10.6151
R1070 B.n500 B.n434 10.6151
R1071 B.n506 B.n434 10.6151
R1072 B.n507 B.n506 10.6151
R1073 B.n508 B.n507 10.6151
R1074 B.n508 B.n432 10.6151
R1075 B.n514 B.n432 10.6151
R1076 B.n515 B.n514 10.6151
R1077 B.n516 B.n515 10.6151
R1078 B.n516 B.n430 10.6151
R1079 B.n522 B.n430 10.6151
R1080 B.n523 B.n522 10.6151
R1081 B.n524 B.n523 10.6151
R1082 B.n524 B.n428 10.6151
R1083 B.n530 B.n428 10.6151
R1084 B.n531 B.n530 10.6151
R1085 B.n532 B.n531 10.6151
R1086 B.n532 B.n426 10.6151
R1087 B.n538 B.n426 10.6151
R1088 B.n539 B.n538 10.6151
R1089 B.n540 B.n539 10.6151
R1090 B.n540 B.n424 10.6151
R1091 B.n546 B.n424 10.6151
R1092 B.n547 B.n546 10.6151
R1093 B.n548 B.n547 10.6151
R1094 B.n548 B.n422 10.6151
R1095 B.n554 B.n422 10.6151
R1096 B.n555 B.n554 10.6151
R1097 B.n556 B.n555 10.6151
R1098 B.n556 B.n420 10.6151
R1099 B.n562 B.n420 10.6151
R1100 B.n563 B.n562 10.6151
R1101 B.n565 B.n416 10.6151
R1102 B.n571 B.n416 10.6151
R1103 B.n572 B.n571 10.6151
R1104 B.n573 B.n572 10.6151
R1105 B.n573 B.n414 10.6151
R1106 B.n579 B.n414 10.6151
R1107 B.n580 B.n579 10.6151
R1108 B.n584 B.n580 10.6151
R1109 B.n590 B.n412 10.6151
R1110 B.n591 B.n590 10.6151
R1111 B.n592 B.n591 10.6151
R1112 B.n592 B.n410 10.6151
R1113 B.n598 B.n410 10.6151
R1114 B.n599 B.n598 10.6151
R1115 B.n600 B.n599 10.6151
R1116 B.n600 B.n408 10.6151
R1117 B.n606 B.n408 10.6151
R1118 B.n607 B.n606 10.6151
R1119 B.n608 B.n607 10.6151
R1120 B.n608 B.n406 10.6151
R1121 B.n614 B.n406 10.6151
R1122 B.n615 B.n614 10.6151
R1123 B.n616 B.n615 10.6151
R1124 B.n616 B.n404 10.6151
R1125 B.n622 B.n404 10.6151
R1126 B.n623 B.n622 10.6151
R1127 B.n624 B.n623 10.6151
R1128 B.n624 B.n402 10.6151
R1129 B.n630 B.n402 10.6151
R1130 B.n631 B.n630 10.6151
R1131 B.n632 B.n631 10.6151
R1132 B.n632 B.n400 10.6151
R1133 B.n638 B.n400 10.6151
R1134 B.n639 B.n638 10.6151
R1135 B.n640 B.n639 10.6151
R1136 B.n640 B.n398 10.6151
R1137 B.n646 B.n398 10.6151
R1138 B.n647 B.n646 10.6151
R1139 B.n648 B.n647 10.6151
R1140 B.n648 B.n396 10.6151
R1141 B.n654 B.n396 10.6151
R1142 B.n655 B.n654 10.6151
R1143 B.n656 B.n655 10.6151
R1144 B.n656 B.n394 10.6151
R1145 B.n662 B.n394 10.6151
R1146 B.n663 B.n662 10.6151
R1147 B.n664 B.n663 10.6151
R1148 B.n664 B.n392 10.6151
R1149 B.n670 B.n392 10.6151
R1150 B.n671 B.n670 10.6151
R1151 B.n672 B.n671 10.6151
R1152 B.n672 B.n390 10.6151
R1153 B.n678 B.n390 10.6151
R1154 B.n679 B.n678 10.6151
R1155 B.n680 B.n679 10.6151
R1156 B.n680 B.n388 10.6151
R1157 B.n686 B.n388 10.6151
R1158 B.n687 B.n686 10.6151
R1159 B.n688 B.n687 10.6151
R1160 B.n688 B.n386 10.6151
R1161 B.n694 B.n386 10.6151
R1162 B.n695 B.n694 10.6151
R1163 B.n696 B.n695 10.6151
R1164 B.n696 B.n384 10.6151
R1165 B.n702 B.n384 10.6151
R1166 B.n703 B.n702 10.6151
R1167 B.n704 B.n376 10.6151
R1168 B.n714 B.n376 10.6151
R1169 B.n715 B.n714 10.6151
R1170 B.n716 B.n715 10.6151
R1171 B.n716 B.n369 10.6151
R1172 B.n727 B.n369 10.6151
R1173 B.n728 B.n727 10.6151
R1174 B.n729 B.n728 10.6151
R1175 B.n729 B.n361 10.6151
R1176 B.n739 B.n361 10.6151
R1177 B.n740 B.n739 10.6151
R1178 B.n742 B.n740 10.6151
R1179 B.n742 B.n741 10.6151
R1180 B.n741 B.n353 10.6151
R1181 B.n753 B.n353 10.6151
R1182 B.n754 B.n753 10.6151
R1183 B.n755 B.n754 10.6151
R1184 B.n756 B.n755 10.6151
R1185 B.n757 B.n756 10.6151
R1186 B.n761 B.n757 10.6151
R1187 B.n762 B.n761 10.6151
R1188 B.n763 B.n762 10.6151
R1189 B.n764 B.n763 10.6151
R1190 B.n766 B.n764 10.6151
R1191 B.n767 B.n766 10.6151
R1192 B.n768 B.n767 10.6151
R1193 B.n769 B.n768 10.6151
R1194 B.n771 B.n769 10.6151
R1195 B.n772 B.n771 10.6151
R1196 B.n773 B.n772 10.6151
R1197 B.n774 B.n773 10.6151
R1198 B.n776 B.n774 10.6151
R1199 B.n777 B.n776 10.6151
R1200 B.n809 B.n1 10.6151
R1201 B.n809 B.n808 10.6151
R1202 B.n808 B.n807 10.6151
R1203 B.n807 B.n10 10.6151
R1204 B.n801 B.n10 10.6151
R1205 B.n801 B.n800 10.6151
R1206 B.n800 B.n799 10.6151
R1207 B.n799 B.n17 10.6151
R1208 B.n793 B.n17 10.6151
R1209 B.n793 B.n792 10.6151
R1210 B.n792 B.n791 10.6151
R1211 B.n791 B.n23 10.6151
R1212 B.n785 B.n23 10.6151
R1213 B.n785 B.n784 10.6151
R1214 B.n784 B.n783 10.6151
R1215 B.n103 B.n31 10.6151
R1216 B.n106 B.n103 10.6151
R1217 B.n107 B.n106 10.6151
R1218 B.n110 B.n107 10.6151
R1219 B.n111 B.n110 10.6151
R1220 B.n114 B.n111 10.6151
R1221 B.n115 B.n114 10.6151
R1222 B.n118 B.n115 10.6151
R1223 B.n119 B.n118 10.6151
R1224 B.n122 B.n119 10.6151
R1225 B.n123 B.n122 10.6151
R1226 B.n126 B.n123 10.6151
R1227 B.n127 B.n126 10.6151
R1228 B.n130 B.n127 10.6151
R1229 B.n131 B.n130 10.6151
R1230 B.n134 B.n131 10.6151
R1231 B.n135 B.n134 10.6151
R1232 B.n138 B.n135 10.6151
R1233 B.n139 B.n138 10.6151
R1234 B.n142 B.n139 10.6151
R1235 B.n143 B.n142 10.6151
R1236 B.n146 B.n143 10.6151
R1237 B.n147 B.n146 10.6151
R1238 B.n150 B.n147 10.6151
R1239 B.n151 B.n150 10.6151
R1240 B.n154 B.n151 10.6151
R1241 B.n155 B.n154 10.6151
R1242 B.n158 B.n155 10.6151
R1243 B.n159 B.n158 10.6151
R1244 B.n162 B.n159 10.6151
R1245 B.n163 B.n162 10.6151
R1246 B.n166 B.n163 10.6151
R1247 B.n167 B.n166 10.6151
R1248 B.n170 B.n167 10.6151
R1249 B.n171 B.n170 10.6151
R1250 B.n174 B.n171 10.6151
R1251 B.n175 B.n174 10.6151
R1252 B.n178 B.n175 10.6151
R1253 B.n179 B.n178 10.6151
R1254 B.n182 B.n179 10.6151
R1255 B.n183 B.n182 10.6151
R1256 B.n186 B.n183 10.6151
R1257 B.n187 B.n186 10.6151
R1258 B.n190 B.n187 10.6151
R1259 B.n191 B.n190 10.6151
R1260 B.n194 B.n191 10.6151
R1261 B.n195 B.n194 10.6151
R1262 B.n198 B.n195 10.6151
R1263 B.n199 B.n198 10.6151
R1264 B.n202 B.n199 10.6151
R1265 B.n203 B.n202 10.6151
R1266 B.n206 B.n203 10.6151
R1267 B.n207 B.n206 10.6151
R1268 B.n210 B.n207 10.6151
R1269 B.n211 B.n210 10.6151
R1270 B.n214 B.n211 10.6151
R1271 B.n215 B.n214 10.6151
R1272 B.n218 B.n215 10.6151
R1273 B.n223 B.n220 10.6151
R1274 B.n224 B.n223 10.6151
R1275 B.n227 B.n224 10.6151
R1276 B.n228 B.n227 10.6151
R1277 B.n231 B.n228 10.6151
R1278 B.n232 B.n231 10.6151
R1279 B.n235 B.n232 10.6151
R1280 B.n236 B.n235 10.6151
R1281 B.n240 B.n239 10.6151
R1282 B.n243 B.n240 10.6151
R1283 B.n244 B.n243 10.6151
R1284 B.n247 B.n244 10.6151
R1285 B.n248 B.n247 10.6151
R1286 B.n251 B.n248 10.6151
R1287 B.n252 B.n251 10.6151
R1288 B.n255 B.n252 10.6151
R1289 B.n256 B.n255 10.6151
R1290 B.n259 B.n256 10.6151
R1291 B.n260 B.n259 10.6151
R1292 B.n263 B.n260 10.6151
R1293 B.n264 B.n263 10.6151
R1294 B.n267 B.n264 10.6151
R1295 B.n268 B.n267 10.6151
R1296 B.n271 B.n268 10.6151
R1297 B.n272 B.n271 10.6151
R1298 B.n275 B.n272 10.6151
R1299 B.n276 B.n275 10.6151
R1300 B.n279 B.n276 10.6151
R1301 B.n280 B.n279 10.6151
R1302 B.n283 B.n280 10.6151
R1303 B.n284 B.n283 10.6151
R1304 B.n287 B.n284 10.6151
R1305 B.n288 B.n287 10.6151
R1306 B.n291 B.n288 10.6151
R1307 B.n292 B.n291 10.6151
R1308 B.n295 B.n292 10.6151
R1309 B.n296 B.n295 10.6151
R1310 B.n299 B.n296 10.6151
R1311 B.n300 B.n299 10.6151
R1312 B.n303 B.n300 10.6151
R1313 B.n304 B.n303 10.6151
R1314 B.n307 B.n304 10.6151
R1315 B.n308 B.n307 10.6151
R1316 B.n311 B.n308 10.6151
R1317 B.n312 B.n311 10.6151
R1318 B.n315 B.n312 10.6151
R1319 B.n316 B.n315 10.6151
R1320 B.n319 B.n316 10.6151
R1321 B.n320 B.n319 10.6151
R1322 B.n323 B.n320 10.6151
R1323 B.n324 B.n323 10.6151
R1324 B.n327 B.n324 10.6151
R1325 B.n328 B.n327 10.6151
R1326 B.n331 B.n328 10.6151
R1327 B.n332 B.n331 10.6151
R1328 B.n335 B.n332 10.6151
R1329 B.n336 B.n335 10.6151
R1330 B.n339 B.n336 10.6151
R1331 B.n340 B.n339 10.6151
R1332 B.n343 B.n340 10.6151
R1333 B.n344 B.n343 10.6151
R1334 B.n347 B.n344 10.6151
R1335 B.n348 B.n347 10.6151
R1336 B.n351 B.n348 10.6151
R1337 B.n352 B.n351 10.6151
R1338 B.n778 B.n352 10.6151
R1339 B.n817 B.n0 8.11757
R1340 B.n817 B.n1 8.11757
R1341 B.n565 B.n564 7.18099
R1342 B.n584 B.n583 7.18099
R1343 B.n220 B.n219 7.18099
R1344 B.n236 B.n100 7.18099
R1345 B.t1 B.n355 5.72842
R1346 B.n759 B.t0 5.72842
R1347 B.n564 B.n563 3.43465
R1348 B.n583 B.n412 3.43465
R1349 B.n219 B.n218 3.43465
R1350 B.n239 B.n100 3.43465
R1351 VN VN.t0 639.361
R1352 VN VN.t1 594.035
R1353 VTAIL.n1 VTAIL.t3 48.9734
R1354 VTAIL.n3 VTAIL.t2 48.9724
R1355 VTAIL.n0 VTAIL.t0 48.9724
R1356 VTAIL.n2 VTAIL.t1 48.9724
R1357 VTAIL.n1 VTAIL.n0 30.1169
R1358 VTAIL.n3 VTAIL.n2 28.9014
R1359 VTAIL.n2 VTAIL.n1 1.07809
R1360 VTAIL VTAIL.n0 0.832397
R1361 VTAIL VTAIL.n3 0.24619
R1362 VDD2.n0 VDD2.t0 107.061
R1363 VDD2.n0 VDD2.t1 65.6512
R1364 VDD2 VDD2.n0 0.362569
R1365 VP.n0 VP.t0 638.981
R1366 VP.n0 VP.t1 593.985
R1367 VP VP.n0 0.0516364
R1368 VDD1 VDD1.t0 107.889
R1369 VDD1 VDD1.t1 66.0133
C0 VDD1 VP 3.38889f
C1 VDD2 VTAIL 7.13886f
C2 VTAIL VN 2.57135f
C3 VDD2 VP 0.271558f
C4 VN VP 5.79814f
C5 VTAIL VP 2.58605f
C6 VDD1 VDD2 0.501765f
C7 VDD1 VN 0.148762f
C8 VDD1 VTAIL 7.10378f
C9 VDD2 VN 3.27159f
C10 VDD2 B 4.929484f
C11 VDD1 B 8.226939f
C12 VTAIL B 8.79491f
C13 VN B 10.71351f
C14 VP B 4.879618f
C15 VDD1.t1 B 3.32277f
C16 VDD1.t0 B 3.95922f
C17 VP.t0 B 3.11521f
C18 VP.t1 B 2.90574f
C19 VP.n0 B 5.75077f
C20 VDD2.t0 B 3.92097f
C21 VDD2.t1 B 3.31343f
C22 VDD2.n0 B 3.10183f
C23 VTAIL.t0 B 3.17092f
C24 VTAIL.n0 B 1.70216f
C25 VTAIL.t3 B 3.17092f
C26 VTAIL.n1 B 1.71782f
C27 VTAIL.t1 B 3.17091f
C28 VTAIL.n2 B 1.64036f
C29 VTAIL.t2 B 3.17092f
C30 VTAIL.n3 B 1.58733f
C31 VN.t1 B 2.86462f
C32 VN.t0 B 3.0749f
.ends

