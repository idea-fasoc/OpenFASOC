* NGSPICE file created from diff_pair_sample_0384.ext - technology: sky130A

.subckt diff_pair_sample_0384 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=2.11
X1 B.t8 B.t6 B.t7 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=2.11
X2 VTAIL.t7 VN.t0 VDD2.t3 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=2.11
X3 B.t5 B.t3 B.t4 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=2.11
X4 VDD1.t3 VP.t0 VTAIL.t0 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=2.11
X5 VDD1.t2 VP.t1 VTAIL.t1 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=2.11
X6 VDD2.t0 VN.t1 VTAIL.t6 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=2.11
X7 VDD2.t2 VN.t2 VTAIL.t5 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=2.11
X8 VTAIL.t2 VP.t2 VDD1.t1 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=2.11
X9 VTAIL.t4 VN.t3 VDD2.t1 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=2.11
X10 B.t2 B.t0 B.t1 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=2.11
X11 VTAIL.t3 VP.t3 VDD1.t0 w_n2434_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=2.11
R0 B.n279 B.n84 585
R1 B.n278 B.n277 585
R2 B.n276 B.n85 585
R3 B.n275 B.n274 585
R4 B.n273 B.n86 585
R5 B.n272 B.n271 585
R6 B.n270 B.n87 585
R7 B.n269 B.n268 585
R8 B.n267 B.n88 585
R9 B.n266 B.n265 585
R10 B.n264 B.n89 585
R11 B.n263 B.n262 585
R12 B.n261 B.n90 585
R13 B.n260 B.n259 585
R14 B.n258 B.n91 585
R15 B.n257 B.n256 585
R16 B.n255 B.n92 585
R17 B.n254 B.n253 585
R18 B.n252 B.n93 585
R19 B.n251 B.n250 585
R20 B.n249 B.n94 585
R21 B.n248 B.n247 585
R22 B.n246 B.n95 585
R23 B.n245 B.n244 585
R24 B.n243 B.n96 585
R25 B.n242 B.n241 585
R26 B.n240 B.n97 585
R27 B.n239 B.n238 585
R28 B.n237 B.n98 585
R29 B.n236 B.n235 585
R30 B.n231 B.n99 585
R31 B.n230 B.n229 585
R32 B.n228 B.n100 585
R33 B.n227 B.n226 585
R34 B.n225 B.n101 585
R35 B.n224 B.n223 585
R36 B.n222 B.n102 585
R37 B.n221 B.n220 585
R38 B.n218 B.n103 585
R39 B.n217 B.n216 585
R40 B.n215 B.n106 585
R41 B.n214 B.n213 585
R42 B.n212 B.n107 585
R43 B.n211 B.n210 585
R44 B.n209 B.n108 585
R45 B.n208 B.n207 585
R46 B.n206 B.n109 585
R47 B.n205 B.n204 585
R48 B.n203 B.n110 585
R49 B.n202 B.n201 585
R50 B.n200 B.n111 585
R51 B.n199 B.n198 585
R52 B.n197 B.n112 585
R53 B.n196 B.n195 585
R54 B.n194 B.n113 585
R55 B.n193 B.n192 585
R56 B.n191 B.n114 585
R57 B.n190 B.n189 585
R58 B.n188 B.n115 585
R59 B.n187 B.n186 585
R60 B.n185 B.n116 585
R61 B.n184 B.n183 585
R62 B.n182 B.n117 585
R63 B.n181 B.n180 585
R64 B.n179 B.n118 585
R65 B.n178 B.n177 585
R66 B.n176 B.n119 585
R67 B.n281 B.n280 585
R68 B.n282 B.n83 585
R69 B.n284 B.n283 585
R70 B.n285 B.n82 585
R71 B.n287 B.n286 585
R72 B.n288 B.n81 585
R73 B.n290 B.n289 585
R74 B.n291 B.n80 585
R75 B.n293 B.n292 585
R76 B.n294 B.n79 585
R77 B.n296 B.n295 585
R78 B.n297 B.n78 585
R79 B.n299 B.n298 585
R80 B.n300 B.n77 585
R81 B.n302 B.n301 585
R82 B.n303 B.n76 585
R83 B.n305 B.n304 585
R84 B.n306 B.n75 585
R85 B.n308 B.n307 585
R86 B.n309 B.n74 585
R87 B.n311 B.n310 585
R88 B.n312 B.n73 585
R89 B.n314 B.n313 585
R90 B.n315 B.n72 585
R91 B.n317 B.n316 585
R92 B.n318 B.n71 585
R93 B.n320 B.n319 585
R94 B.n321 B.n70 585
R95 B.n323 B.n322 585
R96 B.n324 B.n69 585
R97 B.n326 B.n325 585
R98 B.n327 B.n68 585
R99 B.n329 B.n328 585
R100 B.n330 B.n67 585
R101 B.n332 B.n331 585
R102 B.n333 B.n66 585
R103 B.n335 B.n334 585
R104 B.n336 B.n65 585
R105 B.n338 B.n337 585
R106 B.n339 B.n64 585
R107 B.n341 B.n340 585
R108 B.n342 B.n63 585
R109 B.n344 B.n343 585
R110 B.n345 B.n62 585
R111 B.n347 B.n346 585
R112 B.n348 B.n61 585
R113 B.n350 B.n349 585
R114 B.n351 B.n60 585
R115 B.n353 B.n352 585
R116 B.n354 B.n59 585
R117 B.n356 B.n355 585
R118 B.n357 B.n58 585
R119 B.n359 B.n358 585
R120 B.n360 B.n57 585
R121 B.n362 B.n361 585
R122 B.n363 B.n56 585
R123 B.n365 B.n364 585
R124 B.n366 B.n55 585
R125 B.n368 B.n367 585
R126 B.n369 B.n54 585
R127 B.n472 B.n471 585
R128 B.n470 B.n17 585
R129 B.n469 B.n468 585
R130 B.n467 B.n18 585
R131 B.n466 B.n465 585
R132 B.n464 B.n19 585
R133 B.n463 B.n462 585
R134 B.n461 B.n20 585
R135 B.n460 B.n459 585
R136 B.n458 B.n21 585
R137 B.n457 B.n456 585
R138 B.n455 B.n22 585
R139 B.n454 B.n453 585
R140 B.n452 B.n23 585
R141 B.n451 B.n450 585
R142 B.n449 B.n24 585
R143 B.n448 B.n447 585
R144 B.n446 B.n25 585
R145 B.n445 B.n444 585
R146 B.n443 B.n26 585
R147 B.n442 B.n441 585
R148 B.n440 B.n27 585
R149 B.n439 B.n438 585
R150 B.n437 B.n28 585
R151 B.n436 B.n435 585
R152 B.n434 B.n29 585
R153 B.n433 B.n432 585
R154 B.n431 B.n30 585
R155 B.n430 B.n429 585
R156 B.n427 B.n31 585
R157 B.n426 B.n425 585
R158 B.n424 B.n34 585
R159 B.n423 B.n422 585
R160 B.n421 B.n35 585
R161 B.n420 B.n419 585
R162 B.n418 B.n36 585
R163 B.n417 B.n416 585
R164 B.n415 B.n37 585
R165 B.n413 B.n412 585
R166 B.n411 B.n40 585
R167 B.n410 B.n409 585
R168 B.n408 B.n41 585
R169 B.n407 B.n406 585
R170 B.n405 B.n42 585
R171 B.n404 B.n403 585
R172 B.n402 B.n43 585
R173 B.n401 B.n400 585
R174 B.n399 B.n44 585
R175 B.n398 B.n397 585
R176 B.n396 B.n45 585
R177 B.n395 B.n394 585
R178 B.n393 B.n46 585
R179 B.n392 B.n391 585
R180 B.n390 B.n47 585
R181 B.n389 B.n388 585
R182 B.n387 B.n48 585
R183 B.n386 B.n385 585
R184 B.n384 B.n49 585
R185 B.n383 B.n382 585
R186 B.n381 B.n50 585
R187 B.n380 B.n379 585
R188 B.n378 B.n51 585
R189 B.n377 B.n376 585
R190 B.n375 B.n52 585
R191 B.n374 B.n373 585
R192 B.n372 B.n53 585
R193 B.n371 B.n370 585
R194 B.n473 B.n16 585
R195 B.n475 B.n474 585
R196 B.n476 B.n15 585
R197 B.n478 B.n477 585
R198 B.n479 B.n14 585
R199 B.n481 B.n480 585
R200 B.n482 B.n13 585
R201 B.n484 B.n483 585
R202 B.n485 B.n12 585
R203 B.n487 B.n486 585
R204 B.n488 B.n11 585
R205 B.n490 B.n489 585
R206 B.n491 B.n10 585
R207 B.n493 B.n492 585
R208 B.n494 B.n9 585
R209 B.n496 B.n495 585
R210 B.n497 B.n8 585
R211 B.n499 B.n498 585
R212 B.n500 B.n7 585
R213 B.n502 B.n501 585
R214 B.n503 B.n6 585
R215 B.n505 B.n504 585
R216 B.n506 B.n5 585
R217 B.n508 B.n507 585
R218 B.n509 B.n4 585
R219 B.n511 B.n510 585
R220 B.n512 B.n3 585
R221 B.n514 B.n513 585
R222 B.n515 B.n0 585
R223 B.n2 B.n1 585
R224 B.n134 B.n133 585
R225 B.n136 B.n135 585
R226 B.n137 B.n132 585
R227 B.n139 B.n138 585
R228 B.n140 B.n131 585
R229 B.n142 B.n141 585
R230 B.n143 B.n130 585
R231 B.n145 B.n144 585
R232 B.n146 B.n129 585
R233 B.n148 B.n147 585
R234 B.n149 B.n128 585
R235 B.n151 B.n150 585
R236 B.n152 B.n127 585
R237 B.n154 B.n153 585
R238 B.n155 B.n126 585
R239 B.n157 B.n156 585
R240 B.n158 B.n125 585
R241 B.n160 B.n159 585
R242 B.n161 B.n124 585
R243 B.n163 B.n162 585
R244 B.n164 B.n123 585
R245 B.n166 B.n165 585
R246 B.n167 B.n122 585
R247 B.n169 B.n168 585
R248 B.n170 B.n121 585
R249 B.n172 B.n171 585
R250 B.n173 B.n120 585
R251 B.n175 B.n174 585
R252 B.n174 B.n119 559.769
R253 B.n280 B.n279 559.769
R254 B.n370 B.n369 559.769
R255 B.n473 B.n472 559.769
R256 B.n232 B.t9 295.652
R257 B.n38 B.t6 295.652
R258 B.n104 B.t3 295.274
R259 B.n32 B.t0 295.274
R260 B.n517 B.n516 256.663
R261 B.n516 B.n515 235.042
R262 B.n516 B.n2 235.042
R263 B.n178 B.n119 163.367
R264 B.n179 B.n178 163.367
R265 B.n180 B.n179 163.367
R266 B.n180 B.n117 163.367
R267 B.n184 B.n117 163.367
R268 B.n185 B.n184 163.367
R269 B.n186 B.n185 163.367
R270 B.n186 B.n115 163.367
R271 B.n190 B.n115 163.367
R272 B.n191 B.n190 163.367
R273 B.n192 B.n191 163.367
R274 B.n192 B.n113 163.367
R275 B.n196 B.n113 163.367
R276 B.n197 B.n196 163.367
R277 B.n198 B.n197 163.367
R278 B.n198 B.n111 163.367
R279 B.n202 B.n111 163.367
R280 B.n203 B.n202 163.367
R281 B.n204 B.n203 163.367
R282 B.n204 B.n109 163.367
R283 B.n208 B.n109 163.367
R284 B.n209 B.n208 163.367
R285 B.n210 B.n209 163.367
R286 B.n210 B.n107 163.367
R287 B.n214 B.n107 163.367
R288 B.n215 B.n214 163.367
R289 B.n216 B.n215 163.367
R290 B.n216 B.n103 163.367
R291 B.n221 B.n103 163.367
R292 B.n222 B.n221 163.367
R293 B.n223 B.n222 163.367
R294 B.n223 B.n101 163.367
R295 B.n227 B.n101 163.367
R296 B.n228 B.n227 163.367
R297 B.n229 B.n228 163.367
R298 B.n229 B.n99 163.367
R299 B.n236 B.n99 163.367
R300 B.n237 B.n236 163.367
R301 B.n238 B.n237 163.367
R302 B.n238 B.n97 163.367
R303 B.n242 B.n97 163.367
R304 B.n243 B.n242 163.367
R305 B.n244 B.n243 163.367
R306 B.n244 B.n95 163.367
R307 B.n248 B.n95 163.367
R308 B.n249 B.n248 163.367
R309 B.n250 B.n249 163.367
R310 B.n250 B.n93 163.367
R311 B.n254 B.n93 163.367
R312 B.n255 B.n254 163.367
R313 B.n256 B.n255 163.367
R314 B.n256 B.n91 163.367
R315 B.n260 B.n91 163.367
R316 B.n261 B.n260 163.367
R317 B.n262 B.n261 163.367
R318 B.n262 B.n89 163.367
R319 B.n266 B.n89 163.367
R320 B.n267 B.n266 163.367
R321 B.n268 B.n267 163.367
R322 B.n268 B.n87 163.367
R323 B.n272 B.n87 163.367
R324 B.n273 B.n272 163.367
R325 B.n274 B.n273 163.367
R326 B.n274 B.n85 163.367
R327 B.n278 B.n85 163.367
R328 B.n279 B.n278 163.367
R329 B.n369 B.n368 163.367
R330 B.n368 B.n55 163.367
R331 B.n364 B.n55 163.367
R332 B.n364 B.n363 163.367
R333 B.n363 B.n362 163.367
R334 B.n362 B.n57 163.367
R335 B.n358 B.n57 163.367
R336 B.n358 B.n357 163.367
R337 B.n357 B.n356 163.367
R338 B.n356 B.n59 163.367
R339 B.n352 B.n59 163.367
R340 B.n352 B.n351 163.367
R341 B.n351 B.n350 163.367
R342 B.n350 B.n61 163.367
R343 B.n346 B.n61 163.367
R344 B.n346 B.n345 163.367
R345 B.n345 B.n344 163.367
R346 B.n344 B.n63 163.367
R347 B.n340 B.n63 163.367
R348 B.n340 B.n339 163.367
R349 B.n339 B.n338 163.367
R350 B.n338 B.n65 163.367
R351 B.n334 B.n65 163.367
R352 B.n334 B.n333 163.367
R353 B.n333 B.n332 163.367
R354 B.n332 B.n67 163.367
R355 B.n328 B.n67 163.367
R356 B.n328 B.n327 163.367
R357 B.n327 B.n326 163.367
R358 B.n326 B.n69 163.367
R359 B.n322 B.n69 163.367
R360 B.n322 B.n321 163.367
R361 B.n321 B.n320 163.367
R362 B.n320 B.n71 163.367
R363 B.n316 B.n71 163.367
R364 B.n316 B.n315 163.367
R365 B.n315 B.n314 163.367
R366 B.n314 B.n73 163.367
R367 B.n310 B.n73 163.367
R368 B.n310 B.n309 163.367
R369 B.n309 B.n308 163.367
R370 B.n308 B.n75 163.367
R371 B.n304 B.n75 163.367
R372 B.n304 B.n303 163.367
R373 B.n303 B.n302 163.367
R374 B.n302 B.n77 163.367
R375 B.n298 B.n77 163.367
R376 B.n298 B.n297 163.367
R377 B.n297 B.n296 163.367
R378 B.n296 B.n79 163.367
R379 B.n292 B.n79 163.367
R380 B.n292 B.n291 163.367
R381 B.n291 B.n290 163.367
R382 B.n290 B.n81 163.367
R383 B.n286 B.n81 163.367
R384 B.n286 B.n285 163.367
R385 B.n285 B.n284 163.367
R386 B.n284 B.n83 163.367
R387 B.n280 B.n83 163.367
R388 B.n472 B.n17 163.367
R389 B.n468 B.n17 163.367
R390 B.n468 B.n467 163.367
R391 B.n467 B.n466 163.367
R392 B.n466 B.n19 163.367
R393 B.n462 B.n19 163.367
R394 B.n462 B.n461 163.367
R395 B.n461 B.n460 163.367
R396 B.n460 B.n21 163.367
R397 B.n456 B.n21 163.367
R398 B.n456 B.n455 163.367
R399 B.n455 B.n454 163.367
R400 B.n454 B.n23 163.367
R401 B.n450 B.n23 163.367
R402 B.n450 B.n449 163.367
R403 B.n449 B.n448 163.367
R404 B.n448 B.n25 163.367
R405 B.n444 B.n25 163.367
R406 B.n444 B.n443 163.367
R407 B.n443 B.n442 163.367
R408 B.n442 B.n27 163.367
R409 B.n438 B.n27 163.367
R410 B.n438 B.n437 163.367
R411 B.n437 B.n436 163.367
R412 B.n436 B.n29 163.367
R413 B.n432 B.n29 163.367
R414 B.n432 B.n431 163.367
R415 B.n431 B.n430 163.367
R416 B.n430 B.n31 163.367
R417 B.n425 B.n31 163.367
R418 B.n425 B.n424 163.367
R419 B.n424 B.n423 163.367
R420 B.n423 B.n35 163.367
R421 B.n419 B.n35 163.367
R422 B.n419 B.n418 163.367
R423 B.n418 B.n417 163.367
R424 B.n417 B.n37 163.367
R425 B.n412 B.n37 163.367
R426 B.n412 B.n411 163.367
R427 B.n411 B.n410 163.367
R428 B.n410 B.n41 163.367
R429 B.n406 B.n41 163.367
R430 B.n406 B.n405 163.367
R431 B.n405 B.n404 163.367
R432 B.n404 B.n43 163.367
R433 B.n400 B.n43 163.367
R434 B.n400 B.n399 163.367
R435 B.n399 B.n398 163.367
R436 B.n398 B.n45 163.367
R437 B.n394 B.n45 163.367
R438 B.n394 B.n393 163.367
R439 B.n393 B.n392 163.367
R440 B.n392 B.n47 163.367
R441 B.n388 B.n47 163.367
R442 B.n388 B.n387 163.367
R443 B.n387 B.n386 163.367
R444 B.n386 B.n49 163.367
R445 B.n382 B.n49 163.367
R446 B.n382 B.n381 163.367
R447 B.n381 B.n380 163.367
R448 B.n380 B.n51 163.367
R449 B.n376 B.n51 163.367
R450 B.n376 B.n375 163.367
R451 B.n375 B.n374 163.367
R452 B.n374 B.n53 163.367
R453 B.n370 B.n53 163.367
R454 B.n474 B.n473 163.367
R455 B.n474 B.n15 163.367
R456 B.n478 B.n15 163.367
R457 B.n479 B.n478 163.367
R458 B.n480 B.n479 163.367
R459 B.n480 B.n13 163.367
R460 B.n484 B.n13 163.367
R461 B.n485 B.n484 163.367
R462 B.n486 B.n485 163.367
R463 B.n486 B.n11 163.367
R464 B.n490 B.n11 163.367
R465 B.n491 B.n490 163.367
R466 B.n492 B.n491 163.367
R467 B.n492 B.n9 163.367
R468 B.n496 B.n9 163.367
R469 B.n497 B.n496 163.367
R470 B.n498 B.n497 163.367
R471 B.n498 B.n7 163.367
R472 B.n502 B.n7 163.367
R473 B.n503 B.n502 163.367
R474 B.n504 B.n503 163.367
R475 B.n504 B.n5 163.367
R476 B.n508 B.n5 163.367
R477 B.n509 B.n508 163.367
R478 B.n510 B.n509 163.367
R479 B.n510 B.n3 163.367
R480 B.n514 B.n3 163.367
R481 B.n515 B.n514 163.367
R482 B.n133 B.n2 163.367
R483 B.n136 B.n133 163.367
R484 B.n137 B.n136 163.367
R485 B.n138 B.n137 163.367
R486 B.n138 B.n131 163.367
R487 B.n142 B.n131 163.367
R488 B.n143 B.n142 163.367
R489 B.n144 B.n143 163.367
R490 B.n144 B.n129 163.367
R491 B.n148 B.n129 163.367
R492 B.n149 B.n148 163.367
R493 B.n150 B.n149 163.367
R494 B.n150 B.n127 163.367
R495 B.n154 B.n127 163.367
R496 B.n155 B.n154 163.367
R497 B.n156 B.n155 163.367
R498 B.n156 B.n125 163.367
R499 B.n160 B.n125 163.367
R500 B.n161 B.n160 163.367
R501 B.n162 B.n161 163.367
R502 B.n162 B.n123 163.367
R503 B.n166 B.n123 163.367
R504 B.n167 B.n166 163.367
R505 B.n168 B.n167 163.367
R506 B.n168 B.n121 163.367
R507 B.n172 B.n121 163.367
R508 B.n173 B.n172 163.367
R509 B.n174 B.n173 163.367
R510 B.n232 B.t10 160.522
R511 B.n38 B.t8 160.522
R512 B.n104 B.t4 160.513
R513 B.n32 B.t2 160.513
R514 B.n233 B.t11 113.201
R515 B.n39 B.t7 113.201
R516 B.n105 B.t5 113.192
R517 B.n33 B.t1 113.192
R518 B.n219 B.n105 59.5399
R519 B.n234 B.n233 59.5399
R520 B.n414 B.n39 59.5399
R521 B.n428 B.n33 59.5399
R522 B.n105 B.n104 47.3217
R523 B.n233 B.n232 47.3217
R524 B.n39 B.n38 47.3217
R525 B.n33 B.n32 47.3217
R526 B.n471 B.n16 36.3712
R527 B.n371 B.n54 36.3712
R528 B.n176 B.n175 36.3712
R529 B.n281 B.n84 36.3712
R530 B B.n517 18.0485
R531 B.n475 B.n16 10.6151
R532 B.n476 B.n475 10.6151
R533 B.n477 B.n476 10.6151
R534 B.n477 B.n14 10.6151
R535 B.n481 B.n14 10.6151
R536 B.n482 B.n481 10.6151
R537 B.n483 B.n482 10.6151
R538 B.n483 B.n12 10.6151
R539 B.n487 B.n12 10.6151
R540 B.n488 B.n487 10.6151
R541 B.n489 B.n488 10.6151
R542 B.n489 B.n10 10.6151
R543 B.n493 B.n10 10.6151
R544 B.n494 B.n493 10.6151
R545 B.n495 B.n494 10.6151
R546 B.n495 B.n8 10.6151
R547 B.n499 B.n8 10.6151
R548 B.n500 B.n499 10.6151
R549 B.n501 B.n500 10.6151
R550 B.n501 B.n6 10.6151
R551 B.n505 B.n6 10.6151
R552 B.n506 B.n505 10.6151
R553 B.n507 B.n506 10.6151
R554 B.n507 B.n4 10.6151
R555 B.n511 B.n4 10.6151
R556 B.n512 B.n511 10.6151
R557 B.n513 B.n512 10.6151
R558 B.n513 B.n0 10.6151
R559 B.n471 B.n470 10.6151
R560 B.n470 B.n469 10.6151
R561 B.n469 B.n18 10.6151
R562 B.n465 B.n18 10.6151
R563 B.n465 B.n464 10.6151
R564 B.n464 B.n463 10.6151
R565 B.n463 B.n20 10.6151
R566 B.n459 B.n20 10.6151
R567 B.n459 B.n458 10.6151
R568 B.n458 B.n457 10.6151
R569 B.n457 B.n22 10.6151
R570 B.n453 B.n22 10.6151
R571 B.n453 B.n452 10.6151
R572 B.n452 B.n451 10.6151
R573 B.n451 B.n24 10.6151
R574 B.n447 B.n24 10.6151
R575 B.n447 B.n446 10.6151
R576 B.n446 B.n445 10.6151
R577 B.n445 B.n26 10.6151
R578 B.n441 B.n26 10.6151
R579 B.n441 B.n440 10.6151
R580 B.n440 B.n439 10.6151
R581 B.n439 B.n28 10.6151
R582 B.n435 B.n28 10.6151
R583 B.n435 B.n434 10.6151
R584 B.n434 B.n433 10.6151
R585 B.n433 B.n30 10.6151
R586 B.n429 B.n30 10.6151
R587 B.n427 B.n426 10.6151
R588 B.n426 B.n34 10.6151
R589 B.n422 B.n34 10.6151
R590 B.n422 B.n421 10.6151
R591 B.n421 B.n420 10.6151
R592 B.n420 B.n36 10.6151
R593 B.n416 B.n36 10.6151
R594 B.n416 B.n415 10.6151
R595 B.n413 B.n40 10.6151
R596 B.n409 B.n40 10.6151
R597 B.n409 B.n408 10.6151
R598 B.n408 B.n407 10.6151
R599 B.n407 B.n42 10.6151
R600 B.n403 B.n42 10.6151
R601 B.n403 B.n402 10.6151
R602 B.n402 B.n401 10.6151
R603 B.n401 B.n44 10.6151
R604 B.n397 B.n44 10.6151
R605 B.n397 B.n396 10.6151
R606 B.n396 B.n395 10.6151
R607 B.n395 B.n46 10.6151
R608 B.n391 B.n46 10.6151
R609 B.n391 B.n390 10.6151
R610 B.n390 B.n389 10.6151
R611 B.n389 B.n48 10.6151
R612 B.n385 B.n48 10.6151
R613 B.n385 B.n384 10.6151
R614 B.n384 B.n383 10.6151
R615 B.n383 B.n50 10.6151
R616 B.n379 B.n50 10.6151
R617 B.n379 B.n378 10.6151
R618 B.n378 B.n377 10.6151
R619 B.n377 B.n52 10.6151
R620 B.n373 B.n52 10.6151
R621 B.n373 B.n372 10.6151
R622 B.n372 B.n371 10.6151
R623 B.n367 B.n54 10.6151
R624 B.n367 B.n366 10.6151
R625 B.n366 B.n365 10.6151
R626 B.n365 B.n56 10.6151
R627 B.n361 B.n56 10.6151
R628 B.n361 B.n360 10.6151
R629 B.n360 B.n359 10.6151
R630 B.n359 B.n58 10.6151
R631 B.n355 B.n58 10.6151
R632 B.n355 B.n354 10.6151
R633 B.n354 B.n353 10.6151
R634 B.n353 B.n60 10.6151
R635 B.n349 B.n60 10.6151
R636 B.n349 B.n348 10.6151
R637 B.n348 B.n347 10.6151
R638 B.n347 B.n62 10.6151
R639 B.n343 B.n62 10.6151
R640 B.n343 B.n342 10.6151
R641 B.n342 B.n341 10.6151
R642 B.n341 B.n64 10.6151
R643 B.n337 B.n64 10.6151
R644 B.n337 B.n336 10.6151
R645 B.n336 B.n335 10.6151
R646 B.n335 B.n66 10.6151
R647 B.n331 B.n66 10.6151
R648 B.n331 B.n330 10.6151
R649 B.n330 B.n329 10.6151
R650 B.n329 B.n68 10.6151
R651 B.n325 B.n68 10.6151
R652 B.n325 B.n324 10.6151
R653 B.n324 B.n323 10.6151
R654 B.n323 B.n70 10.6151
R655 B.n319 B.n70 10.6151
R656 B.n319 B.n318 10.6151
R657 B.n318 B.n317 10.6151
R658 B.n317 B.n72 10.6151
R659 B.n313 B.n72 10.6151
R660 B.n313 B.n312 10.6151
R661 B.n312 B.n311 10.6151
R662 B.n311 B.n74 10.6151
R663 B.n307 B.n74 10.6151
R664 B.n307 B.n306 10.6151
R665 B.n306 B.n305 10.6151
R666 B.n305 B.n76 10.6151
R667 B.n301 B.n76 10.6151
R668 B.n301 B.n300 10.6151
R669 B.n300 B.n299 10.6151
R670 B.n299 B.n78 10.6151
R671 B.n295 B.n78 10.6151
R672 B.n295 B.n294 10.6151
R673 B.n294 B.n293 10.6151
R674 B.n293 B.n80 10.6151
R675 B.n289 B.n80 10.6151
R676 B.n289 B.n288 10.6151
R677 B.n288 B.n287 10.6151
R678 B.n287 B.n82 10.6151
R679 B.n283 B.n82 10.6151
R680 B.n283 B.n282 10.6151
R681 B.n282 B.n281 10.6151
R682 B.n134 B.n1 10.6151
R683 B.n135 B.n134 10.6151
R684 B.n135 B.n132 10.6151
R685 B.n139 B.n132 10.6151
R686 B.n140 B.n139 10.6151
R687 B.n141 B.n140 10.6151
R688 B.n141 B.n130 10.6151
R689 B.n145 B.n130 10.6151
R690 B.n146 B.n145 10.6151
R691 B.n147 B.n146 10.6151
R692 B.n147 B.n128 10.6151
R693 B.n151 B.n128 10.6151
R694 B.n152 B.n151 10.6151
R695 B.n153 B.n152 10.6151
R696 B.n153 B.n126 10.6151
R697 B.n157 B.n126 10.6151
R698 B.n158 B.n157 10.6151
R699 B.n159 B.n158 10.6151
R700 B.n159 B.n124 10.6151
R701 B.n163 B.n124 10.6151
R702 B.n164 B.n163 10.6151
R703 B.n165 B.n164 10.6151
R704 B.n165 B.n122 10.6151
R705 B.n169 B.n122 10.6151
R706 B.n170 B.n169 10.6151
R707 B.n171 B.n170 10.6151
R708 B.n171 B.n120 10.6151
R709 B.n175 B.n120 10.6151
R710 B.n177 B.n176 10.6151
R711 B.n177 B.n118 10.6151
R712 B.n181 B.n118 10.6151
R713 B.n182 B.n181 10.6151
R714 B.n183 B.n182 10.6151
R715 B.n183 B.n116 10.6151
R716 B.n187 B.n116 10.6151
R717 B.n188 B.n187 10.6151
R718 B.n189 B.n188 10.6151
R719 B.n189 B.n114 10.6151
R720 B.n193 B.n114 10.6151
R721 B.n194 B.n193 10.6151
R722 B.n195 B.n194 10.6151
R723 B.n195 B.n112 10.6151
R724 B.n199 B.n112 10.6151
R725 B.n200 B.n199 10.6151
R726 B.n201 B.n200 10.6151
R727 B.n201 B.n110 10.6151
R728 B.n205 B.n110 10.6151
R729 B.n206 B.n205 10.6151
R730 B.n207 B.n206 10.6151
R731 B.n207 B.n108 10.6151
R732 B.n211 B.n108 10.6151
R733 B.n212 B.n211 10.6151
R734 B.n213 B.n212 10.6151
R735 B.n213 B.n106 10.6151
R736 B.n217 B.n106 10.6151
R737 B.n218 B.n217 10.6151
R738 B.n220 B.n102 10.6151
R739 B.n224 B.n102 10.6151
R740 B.n225 B.n224 10.6151
R741 B.n226 B.n225 10.6151
R742 B.n226 B.n100 10.6151
R743 B.n230 B.n100 10.6151
R744 B.n231 B.n230 10.6151
R745 B.n235 B.n231 10.6151
R746 B.n239 B.n98 10.6151
R747 B.n240 B.n239 10.6151
R748 B.n241 B.n240 10.6151
R749 B.n241 B.n96 10.6151
R750 B.n245 B.n96 10.6151
R751 B.n246 B.n245 10.6151
R752 B.n247 B.n246 10.6151
R753 B.n247 B.n94 10.6151
R754 B.n251 B.n94 10.6151
R755 B.n252 B.n251 10.6151
R756 B.n253 B.n252 10.6151
R757 B.n253 B.n92 10.6151
R758 B.n257 B.n92 10.6151
R759 B.n258 B.n257 10.6151
R760 B.n259 B.n258 10.6151
R761 B.n259 B.n90 10.6151
R762 B.n263 B.n90 10.6151
R763 B.n264 B.n263 10.6151
R764 B.n265 B.n264 10.6151
R765 B.n265 B.n88 10.6151
R766 B.n269 B.n88 10.6151
R767 B.n270 B.n269 10.6151
R768 B.n271 B.n270 10.6151
R769 B.n271 B.n86 10.6151
R770 B.n275 B.n86 10.6151
R771 B.n276 B.n275 10.6151
R772 B.n277 B.n276 10.6151
R773 B.n277 B.n84 10.6151
R774 B.n517 B.n0 8.11757
R775 B.n517 B.n1 8.11757
R776 B.n428 B.n427 6.4005
R777 B.n415 B.n414 6.4005
R778 B.n220 B.n219 6.4005
R779 B.n235 B.n234 6.4005
R780 B.n429 B.n428 4.21513
R781 B.n414 B.n413 4.21513
R782 B.n219 B.n218 4.21513
R783 B.n234 B.n98 4.21513
R784 VN.n0 VN.t0 123.987
R785 VN.n1 VN.t1 123.987
R786 VN.n0 VN.t2 123.439
R787 VN.n1 VN.t3 123.439
R788 VN VN.n1 48.7361
R789 VN VN.n0 6.86868
R790 VDD2.n2 VDD2.n0 118.504
R791 VDD2.n2 VDD2.n1 81.8488
R792 VDD2.n1 VDD2.t1 4.22742
R793 VDD2.n1 VDD2.t0 4.22742
R794 VDD2.n0 VDD2.t3 4.22742
R795 VDD2.n0 VDD2.t2 4.22742
R796 VDD2 VDD2.n2 0.0586897
R797 VTAIL.n6 VTAIL.t1 69.3969
R798 VTAIL.n5 VTAIL.t3 69.3968
R799 VTAIL.n4 VTAIL.t6 69.3968
R800 VTAIL.n3 VTAIL.t4 69.3968
R801 VTAIL.n7 VTAIL.t5 69.3967
R802 VTAIL.n0 VTAIL.t7 69.3967
R803 VTAIL.n1 VTAIL.t0 69.3967
R804 VTAIL.n2 VTAIL.t2 69.3967
R805 VTAIL.n7 VTAIL.n6 21.0996
R806 VTAIL.n3 VTAIL.n2 21.0996
R807 VTAIL.n4 VTAIL.n3 2.10395
R808 VTAIL.n6 VTAIL.n5 2.10395
R809 VTAIL.n2 VTAIL.n1 2.10395
R810 VTAIL VTAIL.n0 1.11041
R811 VTAIL VTAIL.n7 0.994035
R812 VTAIL.n5 VTAIL.n4 0.470328
R813 VTAIL.n1 VTAIL.n0 0.470328
R814 VP.n10 VP.n0 161.3
R815 VP.n9 VP.n8 161.3
R816 VP.n7 VP.n1 161.3
R817 VP.n6 VP.n5 161.3
R818 VP.n2 VP.t3 123.987
R819 VP.n2 VP.t1 123.439
R820 VP.n4 VP.t2 87.8341
R821 VP.n11 VP.t0 87.8341
R822 VP.n4 VP.n3 87.7575
R823 VP.n12 VP.n11 87.7575
R824 VP.n9 VP.n1 56.5193
R825 VP.n3 VP.n2 48.4572
R826 VP.n5 VP.n1 24.4675
R827 VP.n10 VP.n9 24.4675
R828 VP.n5 VP.n4 22.9995
R829 VP.n11 VP.n10 22.9995
R830 VP.n6 VP.n3 0.278367
R831 VP.n12 VP.n0 0.278367
R832 VP.n7 VP.n6 0.189894
R833 VP.n8 VP.n7 0.189894
R834 VP.n8 VP.n0 0.189894
R835 VP VP.n12 0.153454
R836 VDD1 VDD1.n1 119.028
R837 VDD1 VDD1.n0 81.9069
R838 VDD1.n0 VDD1.t0 4.22742
R839 VDD1.n0 VDD1.t2 4.22742
R840 VDD1.n1 VDD1.t1 4.22742
R841 VDD1.n1 VDD1.t3 4.22742
C0 VDD1 w_n2434_n2506# 1.24413f
C1 VDD2 w_n2434_n2506# 1.28929f
C2 VTAIL w_n2434_n2506# 2.98059f
C3 VDD1 VP 3.24323f
C4 VDD2 VP 0.363262f
C5 VTAIL VP 3.07435f
C6 VDD1 B 1.06037f
C7 VDD2 B 1.10448f
C8 VTAIL B 3.34592f
C9 VN VDD1 0.148691f
C10 VDD2 VN 3.02927f
C11 VN VTAIL 3.06024f
C12 VP w_n2434_n2506# 4.26046f
C13 B w_n2434_n2506# 7.44678f
C14 VN w_n2434_n2506# 3.94879f
C15 VP B 1.484f
C16 VN VP 5.03752f
C17 VN B 0.969093f
C18 VDD2 VDD1 0.911354f
C19 VDD1 VTAIL 4.258759f
C20 VDD2 VTAIL 4.30968f
C21 VDD2 VSUBS 0.759314f
C22 VDD1 VSUBS 4.886692f
C23 VTAIL VSUBS 0.949606f
C24 VN VSUBS 5.1193f
C25 VP VSUBS 1.88473f
C26 B VSUBS 3.485525f
C27 w_n2434_n2506# VSUBS 75.7363f
C28 VDD1.t0 VSUBS 0.165731f
C29 VDD1.t2 VSUBS 0.165731f
C30 VDD1.n0 VSUBS 1.16607f
C31 VDD1.t1 VSUBS 0.165731f
C32 VDD1.t3 VSUBS 0.165731f
C33 VDD1.n1 VSUBS 1.6934f
C34 VP.n0 VSUBS 0.056609f
C35 VP.t0 VSUBS 1.86616f
C36 VP.n1 VSUBS 0.062681f
C37 VP.t1 VSUBS 2.13415f
C38 VP.t3 VSUBS 2.1382f
C39 VP.n2 VSUBS 3.22067f
C40 VP.n3 VSUBS 2.11348f
C41 VP.t2 VSUBS 1.86616f
C42 VP.n4 VSUBS 0.837936f
C43 VP.n5 VSUBS 0.077655f
C44 VP.n6 VSUBS 0.056609f
C45 VP.n7 VSUBS 0.042938f
C46 VP.n8 VSUBS 0.042938f
C47 VP.n9 VSUBS 0.062681f
C48 VP.n10 VSUBS 0.077655f
C49 VP.n11 VSUBS 0.837936f
C50 VP.n12 VSUBS 0.04834f
C51 VTAIL.t7 VSUBS 1.31595f
C52 VTAIL.n0 VSUBS 0.730368f
C53 VTAIL.t0 VSUBS 1.31595f
C54 VTAIL.n1 VSUBS 0.811575f
C55 VTAIL.t2 VSUBS 1.31595f
C56 VTAIL.n2 VSUBS 1.83152f
C57 VTAIL.t4 VSUBS 1.31596f
C58 VTAIL.n3 VSUBS 1.83151f
C59 VTAIL.t6 VSUBS 1.31596f
C60 VTAIL.n4 VSUBS 0.811567f
C61 VTAIL.t3 VSUBS 1.31596f
C62 VTAIL.n5 VSUBS 0.811567f
C63 VTAIL.t1 VSUBS 1.31596f
C64 VTAIL.n6 VSUBS 1.83151f
C65 VTAIL.t5 VSUBS 1.31595f
C66 VTAIL.n7 VSUBS 1.7408f
C67 VDD2.t3 VSUBS 0.163508f
C68 VDD2.t2 VSUBS 0.163508f
C69 VDD2.n0 VSUBS 1.64882f
C70 VDD2.t1 VSUBS 0.163508f
C71 VDD2.t0 VSUBS 0.163508f
C72 VDD2.n1 VSUBS 1.14995f
C73 VDD2.n2 VSUBS 3.65904f
C74 VN.t0 VSUBS 2.04803f
C75 VN.t2 VSUBS 2.04415f
C76 VN.n0 VSUBS 1.37448f
C77 VN.t1 VSUBS 2.04803f
C78 VN.t3 VSUBS 2.04415f
C79 VN.n1 VSUBS 3.10609f
C80 B.n0 VSUBS 0.006919f
C81 B.n1 VSUBS 0.006919f
C82 B.n2 VSUBS 0.010233f
C83 B.n3 VSUBS 0.007842f
C84 B.n4 VSUBS 0.007842f
C85 B.n5 VSUBS 0.007842f
C86 B.n6 VSUBS 0.007842f
C87 B.n7 VSUBS 0.007842f
C88 B.n8 VSUBS 0.007842f
C89 B.n9 VSUBS 0.007842f
C90 B.n10 VSUBS 0.007842f
C91 B.n11 VSUBS 0.007842f
C92 B.n12 VSUBS 0.007842f
C93 B.n13 VSUBS 0.007842f
C94 B.n14 VSUBS 0.007842f
C95 B.n15 VSUBS 0.007842f
C96 B.n16 VSUBS 0.019384f
C97 B.n17 VSUBS 0.007842f
C98 B.n18 VSUBS 0.007842f
C99 B.n19 VSUBS 0.007842f
C100 B.n20 VSUBS 0.007842f
C101 B.n21 VSUBS 0.007842f
C102 B.n22 VSUBS 0.007842f
C103 B.n23 VSUBS 0.007842f
C104 B.n24 VSUBS 0.007842f
C105 B.n25 VSUBS 0.007842f
C106 B.n26 VSUBS 0.007842f
C107 B.n27 VSUBS 0.007842f
C108 B.n28 VSUBS 0.007842f
C109 B.n29 VSUBS 0.007842f
C110 B.n30 VSUBS 0.007842f
C111 B.n31 VSUBS 0.007842f
C112 B.t1 VSUBS 0.264086f
C113 B.t2 VSUBS 0.283688f
C114 B.t0 VSUBS 0.838627f
C115 B.n32 VSUBS 0.149774f
C116 B.n33 VSUBS 0.077675f
C117 B.n34 VSUBS 0.007842f
C118 B.n35 VSUBS 0.007842f
C119 B.n36 VSUBS 0.007842f
C120 B.n37 VSUBS 0.007842f
C121 B.t7 VSUBS 0.264084f
C122 B.t8 VSUBS 0.283686f
C123 B.t6 VSUBS 0.838726f
C124 B.n38 VSUBS 0.149677f
C125 B.n39 VSUBS 0.077677f
C126 B.n40 VSUBS 0.007842f
C127 B.n41 VSUBS 0.007842f
C128 B.n42 VSUBS 0.007842f
C129 B.n43 VSUBS 0.007842f
C130 B.n44 VSUBS 0.007842f
C131 B.n45 VSUBS 0.007842f
C132 B.n46 VSUBS 0.007842f
C133 B.n47 VSUBS 0.007842f
C134 B.n48 VSUBS 0.007842f
C135 B.n49 VSUBS 0.007842f
C136 B.n50 VSUBS 0.007842f
C137 B.n51 VSUBS 0.007842f
C138 B.n52 VSUBS 0.007842f
C139 B.n53 VSUBS 0.007842f
C140 B.n54 VSUBS 0.019384f
C141 B.n55 VSUBS 0.007842f
C142 B.n56 VSUBS 0.007842f
C143 B.n57 VSUBS 0.007842f
C144 B.n58 VSUBS 0.007842f
C145 B.n59 VSUBS 0.007842f
C146 B.n60 VSUBS 0.007842f
C147 B.n61 VSUBS 0.007842f
C148 B.n62 VSUBS 0.007842f
C149 B.n63 VSUBS 0.007842f
C150 B.n64 VSUBS 0.007842f
C151 B.n65 VSUBS 0.007842f
C152 B.n66 VSUBS 0.007842f
C153 B.n67 VSUBS 0.007842f
C154 B.n68 VSUBS 0.007842f
C155 B.n69 VSUBS 0.007842f
C156 B.n70 VSUBS 0.007842f
C157 B.n71 VSUBS 0.007842f
C158 B.n72 VSUBS 0.007842f
C159 B.n73 VSUBS 0.007842f
C160 B.n74 VSUBS 0.007842f
C161 B.n75 VSUBS 0.007842f
C162 B.n76 VSUBS 0.007842f
C163 B.n77 VSUBS 0.007842f
C164 B.n78 VSUBS 0.007842f
C165 B.n79 VSUBS 0.007842f
C166 B.n80 VSUBS 0.007842f
C167 B.n81 VSUBS 0.007842f
C168 B.n82 VSUBS 0.007842f
C169 B.n83 VSUBS 0.007842f
C170 B.n84 VSUBS 0.019222f
C171 B.n85 VSUBS 0.007842f
C172 B.n86 VSUBS 0.007842f
C173 B.n87 VSUBS 0.007842f
C174 B.n88 VSUBS 0.007842f
C175 B.n89 VSUBS 0.007842f
C176 B.n90 VSUBS 0.007842f
C177 B.n91 VSUBS 0.007842f
C178 B.n92 VSUBS 0.007842f
C179 B.n93 VSUBS 0.007842f
C180 B.n94 VSUBS 0.007842f
C181 B.n95 VSUBS 0.007842f
C182 B.n96 VSUBS 0.007842f
C183 B.n97 VSUBS 0.007842f
C184 B.n98 VSUBS 0.005478f
C185 B.n99 VSUBS 0.007842f
C186 B.n100 VSUBS 0.007842f
C187 B.n101 VSUBS 0.007842f
C188 B.n102 VSUBS 0.007842f
C189 B.n103 VSUBS 0.007842f
C190 B.t5 VSUBS 0.264086f
C191 B.t4 VSUBS 0.283688f
C192 B.t3 VSUBS 0.838627f
C193 B.n104 VSUBS 0.149774f
C194 B.n105 VSUBS 0.077675f
C195 B.n106 VSUBS 0.007842f
C196 B.n107 VSUBS 0.007842f
C197 B.n108 VSUBS 0.007842f
C198 B.n109 VSUBS 0.007842f
C199 B.n110 VSUBS 0.007842f
C200 B.n111 VSUBS 0.007842f
C201 B.n112 VSUBS 0.007842f
C202 B.n113 VSUBS 0.007842f
C203 B.n114 VSUBS 0.007842f
C204 B.n115 VSUBS 0.007842f
C205 B.n116 VSUBS 0.007842f
C206 B.n117 VSUBS 0.007842f
C207 B.n118 VSUBS 0.007842f
C208 B.n119 VSUBS 0.020054f
C209 B.n120 VSUBS 0.007842f
C210 B.n121 VSUBS 0.007842f
C211 B.n122 VSUBS 0.007842f
C212 B.n123 VSUBS 0.007842f
C213 B.n124 VSUBS 0.007842f
C214 B.n125 VSUBS 0.007842f
C215 B.n126 VSUBS 0.007842f
C216 B.n127 VSUBS 0.007842f
C217 B.n128 VSUBS 0.007842f
C218 B.n129 VSUBS 0.007842f
C219 B.n130 VSUBS 0.007842f
C220 B.n131 VSUBS 0.007842f
C221 B.n132 VSUBS 0.007842f
C222 B.n133 VSUBS 0.007842f
C223 B.n134 VSUBS 0.007842f
C224 B.n135 VSUBS 0.007842f
C225 B.n136 VSUBS 0.007842f
C226 B.n137 VSUBS 0.007842f
C227 B.n138 VSUBS 0.007842f
C228 B.n139 VSUBS 0.007842f
C229 B.n140 VSUBS 0.007842f
C230 B.n141 VSUBS 0.007842f
C231 B.n142 VSUBS 0.007842f
C232 B.n143 VSUBS 0.007842f
C233 B.n144 VSUBS 0.007842f
C234 B.n145 VSUBS 0.007842f
C235 B.n146 VSUBS 0.007842f
C236 B.n147 VSUBS 0.007842f
C237 B.n148 VSUBS 0.007842f
C238 B.n149 VSUBS 0.007842f
C239 B.n150 VSUBS 0.007842f
C240 B.n151 VSUBS 0.007842f
C241 B.n152 VSUBS 0.007842f
C242 B.n153 VSUBS 0.007842f
C243 B.n154 VSUBS 0.007842f
C244 B.n155 VSUBS 0.007842f
C245 B.n156 VSUBS 0.007842f
C246 B.n157 VSUBS 0.007842f
C247 B.n158 VSUBS 0.007842f
C248 B.n159 VSUBS 0.007842f
C249 B.n160 VSUBS 0.007842f
C250 B.n161 VSUBS 0.007842f
C251 B.n162 VSUBS 0.007842f
C252 B.n163 VSUBS 0.007842f
C253 B.n164 VSUBS 0.007842f
C254 B.n165 VSUBS 0.007842f
C255 B.n166 VSUBS 0.007842f
C256 B.n167 VSUBS 0.007842f
C257 B.n168 VSUBS 0.007842f
C258 B.n169 VSUBS 0.007842f
C259 B.n170 VSUBS 0.007842f
C260 B.n171 VSUBS 0.007842f
C261 B.n172 VSUBS 0.007842f
C262 B.n173 VSUBS 0.007842f
C263 B.n174 VSUBS 0.019384f
C264 B.n175 VSUBS 0.019384f
C265 B.n176 VSUBS 0.020054f
C266 B.n177 VSUBS 0.007842f
C267 B.n178 VSUBS 0.007842f
C268 B.n179 VSUBS 0.007842f
C269 B.n180 VSUBS 0.007842f
C270 B.n181 VSUBS 0.007842f
C271 B.n182 VSUBS 0.007842f
C272 B.n183 VSUBS 0.007842f
C273 B.n184 VSUBS 0.007842f
C274 B.n185 VSUBS 0.007842f
C275 B.n186 VSUBS 0.007842f
C276 B.n187 VSUBS 0.007842f
C277 B.n188 VSUBS 0.007842f
C278 B.n189 VSUBS 0.007842f
C279 B.n190 VSUBS 0.007842f
C280 B.n191 VSUBS 0.007842f
C281 B.n192 VSUBS 0.007842f
C282 B.n193 VSUBS 0.007842f
C283 B.n194 VSUBS 0.007842f
C284 B.n195 VSUBS 0.007842f
C285 B.n196 VSUBS 0.007842f
C286 B.n197 VSUBS 0.007842f
C287 B.n198 VSUBS 0.007842f
C288 B.n199 VSUBS 0.007842f
C289 B.n200 VSUBS 0.007842f
C290 B.n201 VSUBS 0.007842f
C291 B.n202 VSUBS 0.007842f
C292 B.n203 VSUBS 0.007842f
C293 B.n204 VSUBS 0.007842f
C294 B.n205 VSUBS 0.007842f
C295 B.n206 VSUBS 0.007842f
C296 B.n207 VSUBS 0.007842f
C297 B.n208 VSUBS 0.007842f
C298 B.n209 VSUBS 0.007842f
C299 B.n210 VSUBS 0.007842f
C300 B.n211 VSUBS 0.007842f
C301 B.n212 VSUBS 0.007842f
C302 B.n213 VSUBS 0.007842f
C303 B.n214 VSUBS 0.007842f
C304 B.n215 VSUBS 0.007842f
C305 B.n216 VSUBS 0.007842f
C306 B.n217 VSUBS 0.007842f
C307 B.n218 VSUBS 0.005478f
C308 B.n219 VSUBS 0.018168f
C309 B.n220 VSUBS 0.006285f
C310 B.n221 VSUBS 0.007842f
C311 B.n222 VSUBS 0.007842f
C312 B.n223 VSUBS 0.007842f
C313 B.n224 VSUBS 0.007842f
C314 B.n225 VSUBS 0.007842f
C315 B.n226 VSUBS 0.007842f
C316 B.n227 VSUBS 0.007842f
C317 B.n228 VSUBS 0.007842f
C318 B.n229 VSUBS 0.007842f
C319 B.n230 VSUBS 0.007842f
C320 B.n231 VSUBS 0.007842f
C321 B.t11 VSUBS 0.264084f
C322 B.t10 VSUBS 0.283686f
C323 B.t9 VSUBS 0.838726f
C324 B.n232 VSUBS 0.149677f
C325 B.n233 VSUBS 0.077677f
C326 B.n234 VSUBS 0.018168f
C327 B.n235 VSUBS 0.006285f
C328 B.n236 VSUBS 0.007842f
C329 B.n237 VSUBS 0.007842f
C330 B.n238 VSUBS 0.007842f
C331 B.n239 VSUBS 0.007842f
C332 B.n240 VSUBS 0.007842f
C333 B.n241 VSUBS 0.007842f
C334 B.n242 VSUBS 0.007842f
C335 B.n243 VSUBS 0.007842f
C336 B.n244 VSUBS 0.007842f
C337 B.n245 VSUBS 0.007842f
C338 B.n246 VSUBS 0.007842f
C339 B.n247 VSUBS 0.007842f
C340 B.n248 VSUBS 0.007842f
C341 B.n249 VSUBS 0.007842f
C342 B.n250 VSUBS 0.007842f
C343 B.n251 VSUBS 0.007842f
C344 B.n252 VSUBS 0.007842f
C345 B.n253 VSUBS 0.007842f
C346 B.n254 VSUBS 0.007842f
C347 B.n255 VSUBS 0.007842f
C348 B.n256 VSUBS 0.007842f
C349 B.n257 VSUBS 0.007842f
C350 B.n258 VSUBS 0.007842f
C351 B.n259 VSUBS 0.007842f
C352 B.n260 VSUBS 0.007842f
C353 B.n261 VSUBS 0.007842f
C354 B.n262 VSUBS 0.007842f
C355 B.n263 VSUBS 0.007842f
C356 B.n264 VSUBS 0.007842f
C357 B.n265 VSUBS 0.007842f
C358 B.n266 VSUBS 0.007842f
C359 B.n267 VSUBS 0.007842f
C360 B.n268 VSUBS 0.007842f
C361 B.n269 VSUBS 0.007842f
C362 B.n270 VSUBS 0.007842f
C363 B.n271 VSUBS 0.007842f
C364 B.n272 VSUBS 0.007842f
C365 B.n273 VSUBS 0.007842f
C366 B.n274 VSUBS 0.007842f
C367 B.n275 VSUBS 0.007842f
C368 B.n276 VSUBS 0.007842f
C369 B.n277 VSUBS 0.007842f
C370 B.n278 VSUBS 0.007842f
C371 B.n279 VSUBS 0.020054f
C372 B.n280 VSUBS 0.019384f
C373 B.n281 VSUBS 0.020216f
C374 B.n282 VSUBS 0.007842f
C375 B.n283 VSUBS 0.007842f
C376 B.n284 VSUBS 0.007842f
C377 B.n285 VSUBS 0.007842f
C378 B.n286 VSUBS 0.007842f
C379 B.n287 VSUBS 0.007842f
C380 B.n288 VSUBS 0.007842f
C381 B.n289 VSUBS 0.007842f
C382 B.n290 VSUBS 0.007842f
C383 B.n291 VSUBS 0.007842f
C384 B.n292 VSUBS 0.007842f
C385 B.n293 VSUBS 0.007842f
C386 B.n294 VSUBS 0.007842f
C387 B.n295 VSUBS 0.007842f
C388 B.n296 VSUBS 0.007842f
C389 B.n297 VSUBS 0.007842f
C390 B.n298 VSUBS 0.007842f
C391 B.n299 VSUBS 0.007842f
C392 B.n300 VSUBS 0.007842f
C393 B.n301 VSUBS 0.007842f
C394 B.n302 VSUBS 0.007842f
C395 B.n303 VSUBS 0.007842f
C396 B.n304 VSUBS 0.007842f
C397 B.n305 VSUBS 0.007842f
C398 B.n306 VSUBS 0.007842f
C399 B.n307 VSUBS 0.007842f
C400 B.n308 VSUBS 0.007842f
C401 B.n309 VSUBS 0.007842f
C402 B.n310 VSUBS 0.007842f
C403 B.n311 VSUBS 0.007842f
C404 B.n312 VSUBS 0.007842f
C405 B.n313 VSUBS 0.007842f
C406 B.n314 VSUBS 0.007842f
C407 B.n315 VSUBS 0.007842f
C408 B.n316 VSUBS 0.007842f
C409 B.n317 VSUBS 0.007842f
C410 B.n318 VSUBS 0.007842f
C411 B.n319 VSUBS 0.007842f
C412 B.n320 VSUBS 0.007842f
C413 B.n321 VSUBS 0.007842f
C414 B.n322 VSUBS 0.007842f
C415 B.n323 VSUBS 0.007842f
C416 B.n324 VSUBS 0.007842f
C417 B.n325 VSUBS 0.007842f
C418 B.n326 VSUBS 0.007842f
C419 B.n327 VSUBS 0.007842f
C420 B.n328 VSUBS 0.007842f
C421 B.n329 VSUBS 0.007842f
C422 B.n330 VSUBS 0.007842f
C423 B.n331 VSUBS 0.007842f
C424 B.n332 VSUBS 0.007842f
C425 B.n333 VSUBS 0.007842f
C426 B.n334 VSUBS 0.007842f
C427 B.n335 VSUBS 0.007842f
C428 B.n336 VSUBS 0.007842f
C429 B.n337 VSUBS 0.007842f
C430 B.n338 VSUBS 0.007842f
C431 B.n339 VSUBS 0.007842f
C432 B.n340 VSUBS 0.007842f
C433 B.n341 VSUBS 0.007842f
C434 B.n342 VSUBS 0.007842f
C435 B.n343 VSUBS 0.007842f
C436 B.n344 VSUBS 0.007842f
C437 B.n345 VSUBS 0.007842f
C438 B.n346 VSUBS 0.007842f
C439 B.n347 VSUBS 0.007842f
C440 B.n348 VSUBS 0.007842f
C441 B.n349 VSUBS 0.007842f
C442 B.n350 VSUBS 0.007842f
C443 B.n351 VSUBS 0.007842f
C444 B.n352 VSUBS 0.007842f
C445 B.n353 VSUBS 0.007842f
C446 B.n354 VSUBS 0.007842f
C447 B.n355 VSUBS 0.007842f
C448 B.n356 VSUBS 0.007842f
C449 B.n357 VSUBS 0.007842f
C450 B.n358 VSUBS 0.007842f
C451 B.n359 VSUBS 0.007842f
C452 B.n360 VSUBS 0.007842f
C453 B.n361 VSUBS 0.007842f
C454 B.n362 VSUBS 0.007842f
C455 B.n363 VSUBS 0.007842f
C456 B.n364 VSUBS 0.007842f
C457 B.n365 VSUBS 0.007842f
C458 B.n366 VSUBS 0.007842f
C459 B.n367 VSUBS 0.007842f
C460 B.n368 VSUBS 0.007842f
C461 B.n369 VSUBS 0.019384f
C462 B.n370 VSUBS 0.020054f
C463 B.n371 VSUBS 0.020054f
C464 B.n372 VSUBS 0.007842f
C465 B.n373 VSUBS 0.007842f
C466 B.n374 VSUBS 0.007842f
C467 B.n375 VSUBS 0.007842f
C468 B.n376 VSUBS 0.007842f
C469 B.n377 VSUBS 0.007842f
C470 B.n378 VSUBS 0.007842f
C471 B.n379 VSUBS 0.007842f
C472 B.n380 VSUBS 0.007842f
C473 B.n381 VSUBS 0.007842f
C474 B.n382 VSUBS 0.007842f
C475 B.n383 VSUBS 0.007842f
C476 B.n384 VSUBS 0.007842f
C477 B.n385 VSUBS 0.007842f
C478 B.n386 VSUBS 0.007842f
C479 B.n387 VSUBS 0.007842f
C480 B.n388 VSUBS 0.007842f
C481 B.n389 VSUBS 0.007842f
C482 B.n390 VSUBS 0.007842f
C483 B.n391 VSUBS 0.007842f
C484 B.n392 VSUBS 0.007842f
C485 B.n393 VSUBS 0.007842f
C486 B.n394 VSUBS 0.007842f
C487 B.n395 VSUBS 0.007842f
C488 B.n396 VSUBS 0.007842f
C489 B.n397 VSUBS 0.007842f
C490 B.n398 VSUBS 0.007842f
C491 B.n399 VSUBS 0.007842f
C492 B.n400 VSUBS 0.007842f
C493 B.n401 VSUBS 0.007842f
C494 B.n402 VSUBS 0.007842f
C495 B.n403 VSUBS 0.007842f
C496 B.n404 VSUBS 0.007842f
C497 B.n405 VSUBS 0.007842f
C498 B.n406 VSUBS 0.007842f
C499 B.n407 VSUBS 0.007842f
C500 B.n408 VSUBS 0.007842f
C501 B.n409 VSUBS 0.007842f
C502 B.n410 VSUBS 0.007842f
C503 B.n411 VSUBS 0.007842f
C504 B.n412 VSUBS 0.007842f
C505 B.n413 VSUBS 0.005478f
C506 B.n414 VSUBS 0.018168f
C507 B.n415 VSUBS 0.006285f
C508 B.n416 VSUBS 0.007842f
C509 B.n417 VSUBS 0.007842f
C510 B.n418 VSUBS 0.007842f
C511 B.n419 VSUBS 0.007842f
C512 B.n420 VSUBS 0.007842f
C513 B.n421 VSUBS 0.007842f
C514 B.n422 VSUBS 0.007842f
C515 B.n423 VSUBS 0.007842f
C516 B.n424 VSUBS 0.007842f
C517 B.n425 VSUBS 0.007842f
C518 B.n426 VSUBS 0.007842f
C519 B.n427 VSUBS 0.006285f
C520 B.n428 VSUBS 0.018168f
C521 B.n429 VSUBS 0.005478f
C522 B.n430 VSUBS 0.007842f
C523 B.n431 VSUBS 0.007842f
C524 B.n432 VSUBS 0.007842f
C525 B.n433 VSUBS 0.007842f
C526 B.n434 VSUBS 0.007842f
C527 B.n435 VSUBS 0.007842f
C528 B.n436 VSUBS 0.007842f
C529 B.n437 VSUBS 0.007842f
C530 B.n438 VSUBS 0.007842f
C531 B.n439 VSUBS 0.007842f
C532 B.n440 VSUBS 0.007842f
C533 B.n441 VSUBS 0.007842f
C534 B.n442 VSUBS 0.007842f
C535 B.n443 VSUBS 0.007842f
C536 B.n444 VSUBS 0.007842f
C537 B.n445 VSUBS 0.007842f
C538 B.n446 VSUBS 0.007842f
C539 B.n447 VSUBS 0.007842f
C540 B.n448 VSUBS 0.007842f
C541 B.n449 VSUBS 0.007842f
C542 B.n450 VSUBS 0.007842f
C543 B.n451 VSUBS 0.007842f
C544 B.n452 VSUBS 0.007842f
C545 B.n453 VSUBS 0.007842f
C546 B.n454 VSUBS 0.007842f
C547 B.n455 VSUBS 0.007842f
C548 B.n456 VSUBS 0.007842f
C549 B.n457 VSUBS 0.007842f
C550 B.n458 VSUBS 0.007842f
C551 B.n459 VSUBS 0.007842f
C552 B.n460 VSUBS 0.007842f
C553 B.n461 VSUBS 0.007842f
C554 B.n462 VSUBS 0.007842f
C555 B.n463 VSUBS 0.007842f
C556 B.n464 VSUBS 0.007842f
C557 B.n465 VSUBS 0.007842f
C558 B.n466 VSUBS 0.007842f
C559 B.n467 VSUBS 0.007842f
C560 B.n468 VSUBS 0.007842f
C561 B.n469 VSUBS 0.007842f
C562 B.n470 VSUBS 0.007842f
C563 B.n471 VSUBS 0.020054f
C564 B.n472 VSUBS 0.020054f
C565 B.n473 VSUBS 0.019384f
C566 B.n474 VSUBS 0.007842f
C567 B.n475 VSUBS 0.007842f
C568 B.n476 VSUBS 0.007842f
C569 B.n477 VSUBS 0.007842f
C570 B.n478 VSUBS 0.007842f
C571 B.n479 VSUBS 0.007842f
C572 B.n480 VSUBS 0.007842f
C573 B.n481 VSUBS 0.007842f
C574 B.n482 VSUBS 0.007842f
C575 B.n483 VSUBS 0.007842f
C576 B.n484 VSUBS 0.007842f
C577 B.n485 VSUBS 0.007842f
C578 B.n486 VSUBS 0.007842f
C579 B.n487 VSUBS 0.007842f
C580 B.n488 VSUBS 0.007842f
C581 B.n489 VSUBS 0.007842f
C582 B.n490 VSUBS 0.007842f
C583 B.n491 VSUBS 0.007842f
C584 B.n492 VSUBS 0.007842f
C585 B.n493 VSUBS 0.007842f
C586 B.n494 VSUBS 0.007842f
C587 B.n495 VSUBS 0.007842f
C588 B.n496 VSUBS 0.007842f
C589 B.n497 VSUBS 0.007842f
C590 B.n498 VSUBS 0.007842f
C591 B.n499 VSUBS 0.007842f
C592 B.n500 VSUBS 0.007842f
C593 B.n501 VSUBS 0.007842f
C594 B.n502 VSUBS 0.007842f
C595 B.n503 VSUBS 0.007842f
C596 B.n504 VSUBS 0.007842f
C597 B.n505 VSUBS 0.007842f
C598 B.n506 VSUBS 0.007842f
C599 B.n507 VSUBS 0.007842f
C600 B.n508 VSUBS 0.007842f
C601 B.n509 VSUBS 0.007842f
C602 B.n510 VSUBS 0.007842f
C603 B.n511 VSUBS 0.007842f
C604 B.n512 VSUBS 0.007842f
C605 B.n513 VSUBS 0.007842f
C606 B.n514 VSUBS 0.007842f
C607 B.n515 VSUBS 0.010233f
C608 B.n516 VSUBS 0.010901f
C609 B.n517 VSUBS 0.021677f
.ends

