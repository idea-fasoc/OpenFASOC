* NGSPICE file created from diff_pair_sample_0710.ext - technology: sky130A

.subckt diff_pair_sample_0710 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t13 VN.t0 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
X1 VTAIL.t1 VP.t0 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
X2 VTAIL.t12 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=2.4024 ps=14.89 w=14.56 l=3.32
X3 VTAIL.t2 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
X4 VTAIL.t0 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=2.4024 ps=14.89 w=14.56 l=3.32
X5 VDD1.t4 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=5.6784 ps=29.9 w=14.56 l=3.32
X6 VDD1.t3 VP.t4 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
X7 VDD2.t1 VN.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
X8 VTAIL.t5 VP.t5 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=2.4024 ps=14.89 w=14.56 l=3.32
X9 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=0 ps=0 w=14.56 l=3.32
X10 VDD1.t1 VP.t6 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=5.6784 ps=29.9 w=14.56 l=3.32
X11 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=0 ps=0 w=14.56 l=3.32
X12 VDD2.t0 VN.t3 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
X13 VDD2.t3 VN.t4 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=5.6784 ps=29.9 w=14.56 l=3.32
X14 VDD2.t2 VN.t5 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=5.6784 ps=29.9 w=14.56 l=3.32
X15 VTAIL.t7 VN.t6 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=0 ps=0 w=14.56 l=3.32
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=0 ps=0 w=14.56 l=3.32
X18 VTAIL.t6 VN.t7 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6784 pd=29.9 as=2.4024 ps=14.89 w=14.56 l=3.32
X19 VDD1.t0 VP.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=14.89 as=2.4024 ps=14.89 w=14.56 l=3.32
R0 VN.n68 VN.n67 161.3
R1 VN.n66 VN.n36 161.3
R2 VN.n65 VN.n64 161.3
R3 VN.n63 VN.n37 161.3
R4 VN.n62 VN.n61 161.3
R5 VN.n60 VN.n38 161.3
R6 VN.n59 VN.n58 161.3
R7 VN.n57 VN.n56 161.3
R8 VN.n55 VN.n40 161.3
R9 VN.n54 VN.n53 161.3
R10 VN.n52 VN.n41 161.3
R11 VN.n51 VN.n50 161.3
R12 VN.n49 VN.n42 161.3
R13 VN.n48 VN.n47 161.3
R14 VN.n46 VN.n43 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n1 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n2 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n25 VN.n3 161.3
R21 VN.n24 VN.n23 161.3
R22 VN.n22 VN.n21 161.3
R23 VN.n20 VN.n5 161.3
R24 VN.n19 VN.n18 161.3
R25 VN.n17 VN.n6 161.3
R26 VN.n16 VN.n15 161.3
R27 VN.n14 VN.n7 161.3
R28 VN.n13 VN.n12 161.3
R29 VN.n11 VN.n8 161.3
R30 VN.n45 VN.t4 137.915
R31 VN.n10 VN.t7 137.915
R32 VN.n9 VN.t3 105.692
R33 VN.n4 VN.t0 105.692
R34 VN.n0 VN.t5 105.692
R35 VN.n44 VN.t6 105.692
R36 VN.n39 VN.t2 105.692
R37 VN.n35 VN.t1 105.692
R38 VN.n34 VN.n0 78.9365
R39 VN.n69 VN.n35 78.9365
R40 VN.n10 VN.n9 70.7064
R41 VN.n45 VN.n44 70.7064
R42 VN.n15 VN.n6 56.4773
R43 VN.n50 VN.n41 56.4773
R44 VN VN.n69 56.4297
R45 VN.n26 VN.n2 50.148
R46 VN.n61 VN.n37 50.148
R47 VN.n30 VN.n2 30.6732
R48 VN.n65 VN.n37 30.6732
R49 VN.n13 VN.n8 24.3439
R50 VN.n14 VN.n13 24.3439
R51 VN.n15 VN.n14 24.3439
R52 VN.n19 VN.n6 24.3439
R53 VN.n20 VN.n19 24.3439
R54 VN.n21 VN.n20 24.3439
R55 VN.n25 VN.n24 24.3439
R56 VN.n26 VN.n25 24.3439
R57 VN.n31 VN.n30 24.3439
R58 VN.n32 VN.n31 24.3439
R59 VN.n50 VN.n49 24.3439
R60 VN.n49 VN.n48 24.3439
R61 VN.n48 VN.n43 24.3439
R62 VN.n61 VN.n60 24.3439
R63 VN.n60 VN.n59 24.3439
R64 VN.n56 VN.n55 24.3439
R65 VN.n55 VN.n54 24.3439
R66 VN.n54 VN.n41 24.3439
R67 VN.n67 VN.n66 24.3439
R68 VN.n66 VN.n65 24.3439
R69 VN.n24 VN.n4 20.6924
R70 VN.n59 VN.n39 20.6924
R71 VN.n32 VN.n0 10.955
R72 VN.n67 VN.n35 10.955
R73 VN.n46 VN.n45 4.36823
R74 VN.n11 VN.n10 4.36823
R75 VN.n9 VN.n8 3.65202
R76 VN.n21 VN.n4 3.65202
R77 VN.n44 VN.n43 3.65202
R78 VN.n56 VN.n39 3.65202
R79 VN.n69 VN.n68 0.355081
R80 VN.n34 VN.n33 0.355081
R81 VN VN.n34 0.26685
R82 VN.n68 VN.n36 0.189894
R83 VN.n64 VN.n36 0.189894
R84 VN.n64 VN.n63 0.189894
R85 VN.n63 VN.n62 0.189894
R86 VN.n62 VN.n38 0.189894
R87 VN.n58 VN.n38 0.189894
R88 VN.n58 VN.n57 0.189894
R89 VN.n57 VN.n40 0.189894
R90 VN.n53 VN.n40 0.189894
R91 VN.n53 VN.n52 0.189894
R92 VN.n52 VN.n51 0.189894
R93 VN.n51 VN.n42 0.189894
R94 VN.n47 VN.n42 0.189894
R95 VN.n47 VN.n46 0.189894
R96 VN.n12 VN.n11 0.189894
R97 VN.n12 VN.n7 0.189894
R98 VN.n16 VN.n7 0.189894
R99 VN.n17 VN.n16 0.189894
R100 VN.n18 VN.n17 0.189894
R101 VN.n18 VN.n5 0.189894
R102 VN.n22 VN.n5 0.189894
R103 VN.n23 VN.n22 0.189894
R104 VN.n23 VN.n3 0.189894
R105 VN.n27 VN.n3 0.189894
R106 VN.n28 VN.n27 0.189894
R107 VN.n29 VN.n28 0.189894
R108 VN.n29 VN.n1 0.189894
R109 VN.n33 VN.n1 0.189894
R110 VDD2.n2 VDD2.n1 61.3389
R111 VDD2.n2 VDD2.n0 61.3389
R112 VDD2 VDD2.n5 61.3361
R113 VDD2.n4 VDD2.n3 59.821
R114 VDD2.n4 VDD2.n2 50.4265
R115 VDD2 VDD2.n4 1.63197
R116 VDD2.n5 VDD2.t5 1.36039
R117 VDD2.n5 VDD2.t3 1.36039
R118 VDD2.n3 VDD2.t6 1.36039
R119 VDD2.n3 VDD2.t1 1.36039
R120 VDD2.n1 VDD2.t7 1.36039
R121 VDD2.n1 VDD2.t2 1.36039
R122 VDD2.n0 VDD2.t4 1.36039
R123 VDD2.n0 VDD2.t0 1.36039
R124 VTAIL.n11 VTAIL.t0 44.5021
R125 VTAIL.n10 VTAIL.t9 44.5021
R126 VTAIL.n7 VTAIL.t12 44.5021
R127 VTAIL.n14 VTAIL.t4 44.502
R128 VTAIL.n15 VTAIL.t8 44.5018
R129 VTAIL.n2 VTAIL.t6 44.5018
R130 VTAIL.n3 VTAIL.t14 44.5018
R131 VTAIL.n6 VTAIL.t5 44.5018
R132 VTAIL.n13 VTAIL.n12 43.1422
R133 VTAIL.n9 VTAIL.n8 43.1422
R134 VTAIL.n1 VTAIL.n0 43.1421
R135 VTAIL.n5 VTAIL.n4 43.1421
R136 VTAIL.n15 VTAIL.n14 28.0652
R137 VTAIL.n7 VTAIL.n6 28.0652
R138 VTAIL.n9 VTAIL.n7 3.14705
R139 VTAIL.n10 VTAIL.n9 3.14705
R140 VTAIL.n13 VTAIL.n11 3.14705
R141 VTAIL.n14 VTAIL.n13 3.14705
R142 VTAIL.n6 VTAIL.n5 3.14705
R143 VTAIL.n5 VTAIL.n3 3.14705
R144 VTAIL.n2 VTAIL.n1 3.14705
R145 VTAIL VTAIL.n15 3.08886
R146 VTAIL.n0 VTAIL.t10 1.36039
R147 VTAIL.n0 VTAIL.t13 1.36039
R148 VTAIL.n4 VTAIL.t3 1.36039
R149 VTAIL.n4 VTAIL.t2 1.36039
R150 VTAIL.n12 VTAIL.t15 1.36039
R151 VTAIL.n12 VTAIL.t1 1.36039
R152 VTAIL.n8 VTAIL.t11 1.36039
R153 VTAIL.n8 VTAIL.t7 1.36039
R154 VTAIL.n11 VTAIL.n10 0.470328
R155 VTAIL.n3 VTAIL.n2 0.470328
R156 VTAIL VTAIL.n1 0.0586897
R157 B.n835 B.n834 585
R158 B.n837 B.n172 585
R159 B.n840 B.n839 585
R160 B.n841 B.n171 585
R161 B.n843 B.n842 585
R162 B.n845 B.n170 585
R163 B.n848 B.n847 585
R164 B.n849 B.n169 585
R165 B.n851 B.n850 585
R166 B.n853 B.n168 585
R167 B.n856 B.n855 585
R168 B.n857 B.n167 585
R169 B.n859 B.n858 585
R170 B.n861 B.n166 585
R171 B.n864 B.n863 585
R172 B.n865 B.n165 585
R173 B.n867 B.n866 585
R174 B.n869 B.n164 585
R175 B.n872 B.n871 585
R176 B.n873 B.n163 585
R177 B.n875 B.n874 585
R178 B.n877 B.n162 585
R179 B.n880 B.n879 585
R180 B.n881 B.n161 585
R181 B.n883 B.n882 585
R182 B.n885 B.n160 585
R183 B.n888 B.n887 585
R184 B.n889 B.n159 585
R185 B.n891 B.n890 585
R186 B.n893 B.n158 585
R187 B.n896 B.n895 585
R188 B.n897 B.n157 585
R189 B.n899 B.n898 585
R190 B.n901 B.n156 585
R191 B.n904 B.n903 585
R192 B.n905 B.n155 585
R193 B.n907 B.n906 585
R194 B.n909 B.n154 585
R195 B.n912 B.n911 585
R196 B.n913 B.n153 585
R197 B.n915 B.n914 585
R198 B.n917 B.n152 585
R199 B.n920 B.n919 585
R200 B.n921 B.n151 585
R201 B.n923 B.n922 585
R202 B.n925 B.n150 585
R203 B.n928 B.n927 585
R204 B.n929 B.n146 585
R205 B.n931 B.n930 585
R206 B.n933 B.n145 585
R207 B.n936 B.n935 585
R208 B.n937 B.n144 585
R209 B.n939 B.n938 585
R210 B.n941 B.n143 585
R211 B.n944 B.n943 585
R212 B.n945 B.n142 585
R213 B.n947 B.n946 585
R214 B.n949 B.n141 585
R215 B.n952 B.n951 585
R216 B.n954 B.n138 585
R217 B.n956 B.n955 585
R218 B.n958 B.n137 585
R219 B.n961 B.n960 585
R220 B.n962 B.n136 585
R221 B.n964 B.n963 585
R222 B.n966 B.n135 585
R223 B.n969 B.n968 585
R224 B.n970 B.n134 585
R225 B.n972 B.n971 585
R226 B.n974 B.n133 585
R227 B.n977 B.n976 585
R228 B.n978 B.n132 585
R229 B.n980 B.n979 585
R230 B.n982 B.n131 585
R231 B.n985 B.n984 585
R232 B.n986 B.n130 585
R233 B.n988 B.n987 585
R234 B.n990 B.n129 585
R235 B.n993 B.n992 585
R236 B.n994 B.n128 585
R237 B.n996 B.n995 585
R238 B.n998 B.n127 585
R239 B.n1001 B.n1000 585
R240 B.n1002 B.n126 585
R241 B.n1004 B.n1003 585
R242 B.n1006 B.n125 585
R243 B.n1009 B.n1008 585
R244 B.n1010 B.n124 585
R245 B.n1012 B.n1011 585
R246 B.n1014 B.n123 585
R247 B.n1017 B.n1016 585
R248 B.n1018 B.n122 585
R249 B.n1020 B.n1019 585
R250 B.n1022 B.n121 585
R251 B.n1025 B.n1024 585
R252 B.n1026 B.n120 585
R253 B.n1028 B.n1027 585
R254 B.n1030 B.n119 585
R255 B.n1033 B.n1032 585
R256 B.n1034 B.n118 585
R257 B.n1036 B.n1035 585
R258 B.n1038 B.n117 585
R259 B.n1041 B.n1040 585
R260 B.n1042 B.n116 585
R261 B.n1044 B.n1043 585
R262 B.n1046 B.n115 585
R263 B.n1049 B.n1048 585
R264 B.n1050 B.n114 585
R265 B.n833 B.n112 585
R266 B.n1053 B.n112 585
R267 B.n832 B.n111 585
R268 B.n1054 B.n111 585
R269 B.n831 B.n110 585
R270 B.n1055 B.n110 585
R271 B.n830 B.n829 585
R272 B.n829 B.n106 585
R273 B.n828 B.n105 585
R274 B.n1061 B.n105 585
R275 B.n827 B.n104 585
R276 B.n1062 B.n104 585
R277 B.n826 B.n103 585
R278 B.n1063 B.n103 585
R279 B.n825 B.n824 585
R280 B.n824 B.n99 585
R281 B.n823 B.n98 585
R282 B.n1069 B.n98 585
R283 B.n822 B.n97 585
R284 B.n1070 B.n97 585
R285 B.n821 B.n96 585
R286 B.n1071 B.n96 585
R287 B.n820 B.n819 585
R288 B.n819 B.n92 585
R289 B.n818 B.n91 585
R290 B.n1077 B.n91 585
R291 B.n817 B.n90 585
R292 B.n1078 B.n90 585
R293 B.n816 B.n89 585
R294 B.n1079 B.n89 585
R295 B.n815 B.n814 585
R296 B.n814 B.n85 585
R297 B.n813 B.n84 585
R298 B.n1085 B.n84 585
R299 B.n812 B.n83 585
R300 B.n1086 B.n83 585
R301 B.n811 B.n82 585
R302 B.n1087 B.n82 585
R303 B.n810 B.n809 585
R304 B.n809 B.n78 585
R305 B.n808 B.n77 585
R306 B.n1093 B.n77 585
R307 B.n807 B.n76 585
R308 B.n1094 B.n76 585
R309 B.n806 B.n75 585
R310 B.n1095 B.n75 585
R311 B.n805 B.n804 585
R312 B.n804 B.n71 585
R313 B.n803 B.n70 585
R314 B.n1101 B.n70 585
R315 B.n802 B.n69 585
R316 B.n1102 B.n69 585
R317 B.n801 B.n68 585
R318 B.n1103 B.n68 585
R319 B.n800 B.n799 585
R320 B.n799 B.n64 585
R321 B.n798 B.n63 585
R322 B.n1109 B.n63 585
R323 B.n797 B.n62 585
R324 B.n1110 B.n62 585
R325 B.n796 B.n61 585
R326 B.n1111 B.n61 585
R327 B.n795 B.n794 585
R328 B.n794 B.n57 585
R329 B.n793 B.n56 585
R330 B.n1117 B.n56 585
R331 B.n792 B.n55 585
R332 B.n1118 B.n55 585
R333 B.n791 B.n54 585
R334 B.n1119 B.n54 585
R335 B.n790 B.n789 585
R336 B.n789 B.n50 585
R337 B.n788 B.n49 585
R338 B.n1125 B.n49 585
R339 B.n787 B.n48 585
R340 B.n1126 B.n48 585
R341 B.n786 B.n47 585
R342 B.n1127 B.n47 585
R343 B.n785 B.n784 585
R344 B.n784 B.n43 585
R345 B.n783 B.n42 585
R346 B.n1133 B.n42 585
R347 B.n782 B.n41 585
R348 B.n1134 B.n41 585
R349 B.n781 B.n40 585
R350 B.n1135 B.n40 585
R351 B.n780 B.n779 585
R352 B.n779 B.n36 585
R353 B.n778 B.n35 585
R354 B.n1141 B.n35 585
R355 B.n777 B.n34 585
R356 B.n1142 B.n34 585
R357 B.n776 B.n33 585
R358 B.n1143 B.n33 585
R359 B.n775 B.n774 585
R360 B.n774 B.n29 585
R361 B.n773 B.n28 585
R362 B.n1149 B.n28 585
R363 B.n772 B.n27 585
R364 B.n1150 B.n27 585
R365 B.n771 B.n26 585
R366 B.n1151 B.n26 585
R367 B.n770 B.n769 585
R368 B.n769 B.n22 585
R369 B.n768 B.n21 585
R370 B.n1157 B.n21 585
R371 B.n767 B.n20 585
R372 B.n1158 B.n20 585
R373 B.n766 B.n19 585
R374 B.n1159 B.n19 585
R375 B.n765 B.n764 585
R376 B.n764 B.n18 585
R377 B.n763 B.n14 585
R378 B.n1165 B.n14 585
R379 B.n762 B.n13 585
R380 B.n1166 B.n13 585
R381 B.n761 B.n12 585
R382 B.n1167 B.n12 585
R383 B.n760 B.n759 585
R384 B.n759 B.n8 585
R385 B.n758 B.n7 585
R386 B.n1173 B.n7 585
R387 B.n757 B.n6 585
R388 B.n1174 B.n6 585
R389 B.n756 B.n5 585
R390 B.n1175 B.n5 585
R391 B.n755 B.n754 585
R392 B.n754 B.n4 585
R393 B.n753 B.n173 585
R394 B.n753 B.n752 585
R395 B.n743 B.n174 585
R396 B.n175 B.n174 585
R397 B.n745 B.n744 585
R398 B.n746 B.n745 585
R399 B.n742 B.n180 585
R400 B.n180 B.n179 585
R401 B.n741 B.n740 585
R402 B.n740 B.n739 585
R403 B.n182 B.n181 585
R404 B.n732 B.n182 585
R405 B.n731 B.n730 585
R406 B.n733 B.n731 585
R407 B.n729 B.n187 585
R408 B.n187 B.n186 585
R409 B.n728 B.n727 585
R410 B.n727 B.n726 585
R411 B.n189 B.n188 585
R412 B.n190 B.n189 585
R413 B.n719 B.n718 585
R414 B.n720 B.n719 585
R415 B.n717 B.n195 585
R416 B.n195 B.n194 585
R417 B.n716 B.n715 585
R418 B.n715 B.n714 585
R419 B.n197 B.n196 585
R420 B.n198 B.n197 585
R421 B.n707 B.n706 585
R422 B.n708 B.n707 585
R423 B.n705 B.n203 585
R424 B.n203 B.n202 585
R425 B.n704 B.n703 585
R426 B.n703 B.n702 585
R427 B.n205 B.n204 585
R428 B.n206 B.n205 585
R429 B.n695 B.n694 585
R430 B.n696 B.n695 585
R431 B.n693 B.n211 585
R432 B.n211 B.n210 585
R433 B.n692 B.n691 585
R434 B.n691 B.n690 585
R435 B.n213 B.n212 585
R436 B.n214 B.n213 585
R437 B.n683 B.n682 585
R438 B.n684 B.n683 585
R439 B.n681 B.n219 585
R440 B.n219 B.n218 585
R441 B.n680 B.n679 585
R442 B.n679 B.n678 585
R443 B.n221 B.n220 585
R444 B.n222 B.n221 585
R445 B.n671 B.n670 585
R446 B.n672 B.n671 585
R447 B.n669 B.n226 585
R448 B.n230 B.n226 585
R449 B.n668 B.n667 585
R450 B.n667 B.n666 585
R451 B.n228 B.n227 585
R452 B.n229 B.n228 585
R453 B.n659 B.n658 585
R454 B.n660 B.n659 585
R455 B.n657 B.n235 585
R456 B.n235 B.n234 585
R457 B.n656 B.n655 585
R458 B.n655 B.n654 585
R459 B.n237 B.n236 585
R460 B.n238 B.n237 585
R461 B.n647 B.n646 585
R462 B.n648 B.n647 585
R463 B.n645 B.n243 585
R464 B.n243 B.n242 585
R465 B.n644 B.n643 585
R466 B.n643 B.n642 585
R467 B.n245 B.n244 585
R468 B.n246 B.n245 585
R469 B.n635 B.n634 585
R470 B.n636 B.n635 585
R471 B.n633 B.n251 585
R472 B.n251 B.n250 585
R473 B.n632 B.n631 585
R474 B.n631 B.n630 585
R475 B.n253 B.n252 585
R476 B.n254 B.n253 585
R477 B.n623 B.n622 585
R478 B.n624 B.n623 585
R479 B.n621 B.n259 585
R480 B.n259 B.n258 585
R481 B.n620 B.n619 585
R482 B.n619 B.n618 585
R483 B.n261 B.n260 585
R484 B.n262 B.n261 585
R485 B.n611 B.n610 585
R486 B.n612 B.n611 585
R487 B.n609 B.n267 585
R488 B.n267 B.n266 585
R489 B.n608 B.n607 585
R490 B.n607 B.n606 585
R491 B.n269 B.n268 585
R492 B.n270 B.n269 585
R493 B.n599 B.n598 585
R494 B.n600 B.n599 585
R495 B.n597 B.n275 585
R496 B.n275 B.n274 585
R497 B.n596 B.n595 585
R498 B.n595 B.n594 585
R499 B.n277 B.n276 585
R500 B.n278 B.n277 585
R501 B.n587 B.n586 585
R502 B.n588 B.n587 585
R503 B.n585 B.n283 585
R504 B.n283 B.n282 585
R505 B.n584 B.n583 585
R506 B.n583 B.n582 585
R507 B.n285 B.n284 585
R508 B.n286 B.n285 585
R509 B.n575 B.n574 585
R510 B.n576 B.n575 585
R511 B.n573 B.n291 585
R512 B.n291 B.n290 585
R513 B.n572 B.n571 585
R514 B.n571 B.n570 585
R515 B.n567 B.n295 585
R516 B.n566 B.n565 585
R517 B.n563 B.n296 585
R518 B.n563 B.n294 585
R519 B.n562 B.n561 585
R520 B.n560 B.n559 585
R521 B.n558 B.n298 585
R522 B.n556 B.n555 585
R523 B.n554 B.n299 585
R524 B.n553 B.n552 585
R525 B.n550 B.n300 585
R526 B.n548 B.n547 585
R527 B.n546 B.n301 585
R528 B.n545 B.n544 585
R529 B.n542 B.n302 585
R530 B.n540 B.n539 585
R531 B.n538 B.n303 585
R532 B.n537 B.n536 585
R533 B.n534 B.n304 585
R534 B.n532 B.n531 585
R535 B.n530 B.n305 585
R536 B.n529 B.n528 585
R537 B.n526 B.n306 585
R538 B.n524 B.n523 585
R539 B.n522 B.n307 585
R540 B.n521 B.n520 585
R541 B.n518 B.n308 585
R542 B.n516 B.n515 585
R543 B.n514 B.n309 585
R544 B.n513 B.n512 585
R545 B.n510 B.n310 585
R546 B.n508 B.n507 585
R547 B.n506 B.n311 585
R548 B.n505 B.n504 585
R549 B.n502 B.n312 585
R550 B.n500 B.n499 585
R551 B.n498 B.n313 585
R552 B.n497 B.n496 585
R553 B.n494 B.n314 585
R554 B.n492 B.n491 585
R555 B.n490 B.n315 585
R556 B.n489 B.n488 585
R557 B.n486 B.n316 585
R558 B.n484 B.n483 585
R559 B.n482 B.n317 585
R560 B.n481 B.n480 585
R561 B.n478 B.n318 585
R562 B.n476 B.n475 585
R563 B.n474 B.n319 585
R564 B.n473 B.n472 585
R565 B.n470 B.n469 585
R566 B.n468 B.n467 585
R567 B.n466 B.n324 585
R568 B.n464 B.n463 585
R569 B.n462 B.n325 585
R570 B.n461 B.n460 585
R571 B.n458 B.n326 585
R572 B.n456 B.n455 585
R573 B.n454 B.n327 585
R574 B.n453 B.n452 585
R575 B.n450 B.n449 585
R576 B.n448 B.n447 585
R577 B.n446 B.n332 585
R578 B.n444 B.n443 585
R579 B.n442 B.n333 585
R580 B.n441 B.n440 585
R581 B.n438 B.n334 585
R582 B.n436 B.n435 585
R583 B.n434 B.n335 585
R584 B.n433 B.n432 585
R585 B.n430 B.n336 585
R586 B.n428 B.n427 585
R587 B.n426 B.n337 585
R588 B.n425 B.n424 585
R589 B.n422 B.n338 585
R590 B.n420 B.n419 585
R591 B.n418 B.n339 585
R592 B.n417 B.n416 585
R593 B.n414 B.n340 585
R594 B.n412 B.n411 585
R595 B.n410 B.n341 585
R596 B.n409 B.n408 585
R597 B.n406 B.n342 585
R598 B.n404 B.n403 585
R599 B.n402 B.n343 585
R600 B.n401 B.n400 585
R601 B.n398 B.n344 585
R602 B.n396 B.n395 585
R603 B.n394 B.n345 585
R604 B.n393 B.n392 585
R605 B.n390 B.n346 585
R606 B.n388 B.n387 585
R607 B.n386 B.n347 585
R608 B.n385 B.n384 585
R609 B.n382 B.n348 585
R610 B.n380 B.n379 585
R611 B.n378 B.n349 585
R612 B.n377 B.n376 585
R613 B.n374 B.n350 585
R614 B.n372 B.n371 585
R615 B.n370 B.n351 585
R616 B.n369 B.n368 585
R617 B.n366 B.n352 585
R618 B.n364 B.n363 585
R619 B.n362 B.n353 585
R620 B.n361 B.n360 585
R621 B.n358 B.n354 585
R622 B.n356 B.n355 585
R623 B.n293 B.n292 585
R624 B.n294 B.n293 585
R625 B.n569 B.n568 585
R626 B.n570 B.n569 585
R627 B.n289 B.n288 585
R628 B.n290 B.n289 585
R629 B.n578 B.n577 585
R630 B.n577 B.n576 585
R631 B.n579 B.n287 585
R632 B.n287 B.n286 585
R633 B.n581 B.n580 585
R634 B.n582 B.n581 585
R635 B.n281 B.n280 585
R636 B.n282 B.n281 585
R637 B.n590 B.n589 585
R638 B.n589 B.n588 585
R639 B.n591 B.n279 585
R640 B.n279 B.n278 585
R641 B.n593 B.n592 585
R642 B.n594 B.n593 585
R643 B.n273 B.n272 585
R644 B.n274 B.n273 585
R645 B.n602 B.n601 585
R646 B.n601 B.n600 585
R647 B.n603 B.n271 585
R648 B.n271 B.n270 585
R649 B.n605 B.n604 585
R650 B.n606 B.n605 585
R651 B.n265 B.n264 585
R652 B.n266 B.n265 585
R653 B.n614 B.n613 585
R654 B.n613 B.n612 585
R655 B.n615 B.n263 585
R656 B.n263 B.n262 585
R657 B.n617 B.n616 585
R658 B.n618 B.n617 585
R659 B.n257 B.n256 585
R660 B.n258 B.n257 585
R661 B.n626 B.n625 585
R662 B.n625 B.n624 585
R663 B.n627 B.n255 585
R664 B.n255 B.n254 585
R665 B.n629 B.n628 585
R666 B.n630 B.n629 585
R667 B.n249 B.n248 585
R668 B.n250 B.n249 585
R669 B.n638 B.n637 585
R670 B.n637 B.n636 585
R671 B.n639 B.n247 585
R672 B.n247 B.n246 585
R673 B.n641 B.n640 585
R674 B.n642 B.n641 585
R675 B.n241 B.n240 585
R676 B.n242 B.n241 585
R677 B.n650 B.n649 585
R678 B.n649 B.n648 585
R679 B.n651 B.n239 585
R680 B.n239 B.n238 585
R681 B.n653 B.n652 585
R682 B.n654 B.n653 585
R683 B.n233 B.n232 585
R684 B.n234 B.n233 585
R685 B.n662 B.n661 585
R686 B.n661 B.n660 585
R687 B.n663 B.n231 585
R688 B.n231 B.n229 585
R689 B.n665 B.n664 585
R690 B.n666 B.n665 585
R691 B.n225 B.n224 585
R692 B.n230 B.n225 585
R693 B.n674 B.n673 585
R694 B.n673 B.n672 585
R695 B.n675 B.n223 585
R696 B.n223 B.n222 585
R697 B.n677 B.n676 585
R698 B.n678 B.n677 585
R699 B.n217 B.n216 585
R700 B.n218 B.n217 585
R701 B.n686 B.n685 585
R702 B.n685 B.n684 585
R703 B.n687 B.n215 585
R704 B.n215 B.n214 585
R705 B.n689 B.n688 585
R706 B.n690 B.n689 585
R707 B.n209 B.n208 585
R708 B.n210 B.n209 585
R709 B.n698 B.n697 585
R710 B.n697 B.n696 585
R711 B.n699 B.n207 585
R712 B.n207 B.n206 585
R713 B.n701 B.n700 585
R714 B.n702 B.n701 585
R715 B.n201 B.n200 585
R716 B.n202 B.n201 585
R717 B.n710 B.n709 585
R718 B.n709 B.n708 585
R719 B.n711 B.n199 585
R720 B.n199 B.n198 585
R721 B.n713 B.n712 585
R722 B.n714 B.n713 585
R723 B.n193 B.n192 585
R724 B.n194 B.n193 585
R725 B.n722 B.n721 585
R726 B.n721 B.n720 585
R727 B.n723 B.n191 585
R728 B.n191 B.n190 585
R729 B.n725 B.n724 585
R730 B.n726 B.n725 585
R731 B.n185 B.n184 585
R732 B.n186 B.n185 585
R733 B.n735 B.n734 585
R734 B.n734 B.n733 585
R735 B.n736 B.n183 585
R736 B.n732 B.n183 585
R737 B.n738 B.n737 585
R738 B.n739 B.n738 585
R739 B.n178 B.n177 585
R740 B.n179 B.n178 585
R741 B.n748 B.n747 585
R742 B.n747 B.n746 585
R743 B.n749 B.n176 585
R744 B.n176 B.n175 585
R745 B.n751 B.n750 585
R746 B.n752 B.n751 585
R747 B.n2 B.n0 585
R748 B.n4 B.n2 585
R749 B.n3 B.n1 585
R750 B.n1174 B.n3 585
R751 B.n1172 B.n1171 585
R752 B.n1173 B.n1172 585
R753 B.n1170 B.n9 585
R754 B.n9 B.n8 585
R755 B.n1169 B.n1168 585
R756 B.n1168 B.n1167 585
R757 B.n11 B.n10 585
R758 B.n1166 B.n11 585
R759 B.n1164 B.n1163 585
R760 B.n1165 B.n1164 585
R761 B.n1162 B.n15 585
R762 B.n18 B.n15 585
R763 B.n1161 B.n1160 585
R764 B.n1160 B.n1159 585
R765 B.n17 B.n16 585
R766 B.n1158 B.n17 585
R767 B.n1156 B.n1155 585
R768 B.n1157 B.n1156 585
R769 B.n1154 B.n23 585
R770 B.n23 B.n22 585
R771 B.n1153 B.n1152 585
R772 B.n1152 B.n1151 585
R773 B.n25 B.n24 585
R774 B.n1150 B.n25 585
R775 B.n1148 B.n1147 585
R776 B.n1149 B.n1148 585
R777 B.n1146 B.n30 585
R778 B.n30 B.n29 585
R779 B.n1145 B.n1144 585
R780 B.n1144 B.n1143 585
R781 B.n32 B.n31 585
R782 B.n1142 B.n32 585
R783 B.n1140 B.n1139 585
R784 B.n1141 B.n1140 585
R785 B.n1138 B.n37 585
R786 B.n37 B.n36 585
R787 B.n1137 B.n1136 585
R788 B.n1136 B.n1135 585
R789 B.n39 B.n38 585
R790 B.n1134 B.n39 585
R791 B.n1132 B.n1131 585
R792 B.n1133 B.n1132 585
R793 B.n1130 B.n44 585
R794 B.n44 B.n43 585
R795 B.n1129 B.n1128 585
R796 B.n1128 B.n1127 585
R797 B.n46 B.n45 585
R798 B.n1126 B.n46 585
R799 B.n1124 B.n1123 585
R800 B.n1125 B.n1124 585
R801 B.n1122 B.n51 585
R802 B.n51 B.n50 585
R803 B.n1121 B.n1120 585
R804 B.n1120 B.n1119 585
R805 B.n53 B.n52 585
R806 B.n1118 B.n53 585
R807 B.n1116 B.n1115 585
R808 B.n1117 B.n1116 585
R809 B.n1114 B.n58 585
R810 B.n58 B.n57 585
R811 B.n1113 B.n1112 585
R812 B.n1112 B.n1111 585
R813 B.n60 B.n59 585
R814 B.n1110 B.n60 585
R815 B.n1108 B.n1107 585
R816 B.n1109 B.n1108 585
R817 B.n1106 B.n65 585
R818 B.n65 B.n64 585
R819 B.n1105 B.n1104 585
R820 B.n1104 B.n1103 585
R821 B.n67 B.n66 585
R822 B.n1102 B.n67 585
R823 B.n1100 B.n1099 585
R824 B.n1101 B.n1100 585
R825 B.n1098 B.n72 585
R826 B.n72 B.n71 585
R827 B.n1097 B.n1096 585
R828 B.n1096 B.n1095 585
R829 B.n74 B.n73 585
R830 B.n1094 B.n74 585
R831 B.n1092 B.n1091 585
R832 B.n1093 B.n1092 585
R833 B.n1090 B.n79 585
R834 B.n79 B.n78 585
R835 B.n1089 B.n1088 585
R836 B.n1088 B.n1087 585
R837 B.n81 B.n80 585
R838 B.n1086 B.n81 585
R839 B.n1084 B.n1083 585
R840 B.n1085 B.n1084 585
R841 B.n1082 B.n86 585
R842 B.n86 B.n85 585
R843 B.n1081 B.n1080 585
R844 B.n1080 B.n1079 585
R845 B.n88 B.n87 585
R846 B.n1078 B.n88 585
R847 B.n1076 B.n1075 585
R848 B.n1077 B.n1076 585
R849 B.n1074 B.n93 585
R850 B.n93 B.n92 585
R851 B.n1073 B.n1072 585
R852 B.n1072 B.n1071 585
R853 B.n95 B.n94 585
R854 B.n1070 B.n95 585
R855 B.n1068 B.n1067 585
R856 B.n1069 B.n1068 585
R857 B.n1066 B.n100 585
R858 B.n100 B.n99 585
R859 B.n1065 B.n1064 585
R860 B.n1064 B.n1063 585
R861 B.n102 B.n101 585
R862 B.n1062 B.n102 585
R863 B.n1060 B.n1059 585
R864 B.n1061 B.n1060 585
R865 B.n1058 B.n107 585
R866 B.n107 B.n106 585
R867 B.n1057 B.n1056 585
R868 B.n1056 B.n1055 585
R869 B.n109 B.n108 585
R870 B.n1054 B.n109 585
R871 B.n1052 B.n1051 585
R872 B.n1053 B.n1052 585
R873 B.n1177 B.n1176 585
R874 B.n1176 B.n1175 585
R875 B.n569 B.n295 454.062
R876 B.n1052 B.n114 454.062
R877 B.n571 B.n293 454.062
R878 B.n835 B.n112 454.062
R879 B.n328 B.t12 314.616
R880 B.n320 B.t16 314.616
R881 B.n139 B.t8 314.616
R882 B.n147 B.t19 314.616
R883 B.n836 B.n113 256.663
R884 B.n838 B.n113 256.663
R885 B.n844 B.n113 256.663
R886 B.n846 B.n113 256.663
R887 B.n852 B.n113 256.663
R888 B.n854 B.n113 256.663
R889 B.n860 B.n113 256.663
R890 B.n862 B.n113 256.663
R891 B.n868 B.n113 256.663
R892 B.n870 B.n113 256.663
R893 B.n876 B.n113 256.663
R894 B.n878 B.n113 256.663
R895 B.n884 B.n113 256.663
R896 B.n886 B.n113 256.663
R897 B.n892 B.n113 256.663
R898 B.n894 B.n113 256.663
R899 B.n900 B.n113 256.663
R900 B.n902 B.n113 256.663
R901 B.n908 B.n113 256.663
R902 B.n910 B.n113 256.663
R903 B.n916 B.n113 256.663
R904 B.n918 B.n113 256.663
R905 B.n924 B.n113 256.663
R906 B.n926 B.n113 256.663
R907 B.n932 B.n113 256.663
R908 B.n934 B.n113 256.663
R909 B.n940 B.n113 256.663
R910 B.n942 B.n113 256.663
R911 B.n948 B.n113 256.663
R912 B.n950 B.n113 256.663
R913 B.n957 B.n113 256.663
R914 B.n959 B.n113 256.663
R915 B.n965 B.n113 256.663
R916 B.n967 B.n113 256.663
R917 B.n973 B.n113 256.663
R918 B.n975 B.n113 256.663
R919 B.n981 B.n113 256.663
R920 B.n983 B.n113 256.663
R921 B.n989 B.n113 256.663
R922 B.n991 B.n113 256.663
R923 B.n997 B.n113 256.663
R924 B.n999 B.n113 256.663
R925 B.n1005 B.n113 256.663
R926 B.n1007 B.n113 256.663
R927 B.n1013 B.n113 256.663
R928 B.n1015 B.n113 256.663
R929 B.n1021 B.n113 256.663
R930 B.n1023 B.n113 256.663
R931 B.n1029 B.n113 256.663
R932 B.n1031 B.n113 256.663
R933 B.n1037 B.n113 256.663
R934 B.n1039 B.n113 256.663
R935 B.n1045 B.n113 256.663
R936 B.n1047 B.n113 256.663
R937 B.n564 B.n294 256.663
R938 B.n297 B.n294 256.663
R939 B.n557 B.n294 256.663
R940 B.n551 B.n294 256.663
R941 B.n549 B.n294 256.663
R942 B.n543 B.n294 256.663
R943 B.n541 B.n294 256.663
R944 B.n535 B.n294 256.663
R945 B.n533 B.n294 256.663
R946 B.n527 B.n294 256.663
R947 B.n525 B.n294 256.663
R948 B.n519 B.n294 256.663
R949 B.n517 B.n294 256.663
R950 B.n511 B.n294 256.663
R951 B.n509 B.n294 256.663
R952 B.n503 B.n294 256.663
R953 B.n501 B.n294 256.663
R954 B.n495 B.n294 256.663
R955 B.n493 B.n294 256.663
R956 B.n487 B.n294 256.663
R957 B.n485 B.n294 256.663
R958 B.n479 B.n294 256.663
R959 B.n477 B.n294 256.663
R960 B.n471 B.n294 256.663
R961 B.n323 B.n294 256.663
R962 B.n465 B.n294 256.663
R963 B.n459 B.n294 256.663
R964 B.n457 B.n294 256.663
R965 B.n451 B.n294 256.663
R966 B.n331 B.n294 256.663
R967 B.n445 B.n294 256.663
R968 B.n439 B.n294 256.663
R969 B.n437 B.n294 256.663
R970 B.n431 B.n294 256.663
R971 B.n429 B.n294 256.663
R972 B.n423 B.n294 256.663
R973 B.n421 B.n294 256.663
R974 B.n415 B.n294 256.663
R975 B.n413 B.n294 256.663
R976 B.n407 B.n294 256.663
R977 B.n405 B.n294 256.663
R978 B.n399 B.n294 256.663
R979 B.n397 B.n294 256.663
R980 B.n391 B.n294 256.663
R981 B.n389 B.n294 256.663
R982 B.n383 B.n294 256.663
R983 B.n381 B.n294 256.663
R984 B.n375 B.n294 256.663
R985 B.n373 B.n294 256.663
R986 B.n367 B.n294 256.663
R987 B.n365 B.n294 256.663
R988 B.n359 B.n294 256.663
R989 B.n357 B.n294 256.663
R990 B.n569 B.n289 163.367
R991 B.n577 B.n289 163.367
R992 B.n577 B.n287 163.367
R993 B.n581 B.n287 163.367
R994 B.n581 B.n281 163.367
R995 B.n589 B.n281 163.367
R996 B.n589 B.n279 163.367
R997 B.n593 B.n279 163.367
R998 B.n593 B.n273 163.367
R999 B.n601 B.n273 163.367
R1000 B.n601 B.n271 163.367
R1001 B.n605 B.n271 163.367
R1002 B.n605 B.n265 163.367
R1003 B.n613 B.n265 163.367
R1004 B.n613 B.n263 163.367
R1005 B.n617 B.n263 163.367
R1006 B.n617 B.n257 163.367
R1007 B.n625 B.n257 163.367
R1008 B.n625 B.n255 163.367
R1009 B.n629 B.n255 163.367
R1010 B.n629 B.n249 163.367
R1011 B.n637 B.n249 163.367
R1012 B.n637 B.n247 163.367
R1013 B.n641 B.n247 163.367
R1014 B.n641 B.n241 163.367
R1015 B.n649 B.n241 163.367
R1016 B.n649 B.n239 163.367
R1017 B.n653 B.n239 163.367
R1018 B.n653 B.n233 163.367
R1019 B.n661 B.n233 163.367
R1020 B.n661 B.n231 163.367
R1021 B.n665 B.n231 163.367
R1022 B.n665 B.n225 163.367
R1023 B.n673 B.n225 163.367
R1024 B.n673 B.n223 163.367
R1025 B.n677 B.n223 163.367
R1026 B.n677 B.n217 163.367
R1027 B.n685 B.n217 163.367
R1028 B.n685 B.n215 163.367
R1029 B.n689 B.n215 163.367
R1030 B.n689 B.n209 163.367
R1031 B.n697 B.n209 163.367
R1032 B.n697 B.n207 163.367
R1033 B.n701 B.n207 163.367
R1034 B.n701 B.n201 163.367
R1035 B.n709 B.n201 163.367
R1036 B.n709 B.n199 163.367
R1037 B.n713 B.n199 163.367
R1038 B.n713 B.n193 163.367
R1039 B.n721 B.n193 163.367
R1040 B.n721 B.n191 163.367
R1041 B.n725 B.n191 163.367
R1042 B.n725 B.n185 163.367
R1043 B.n734 B.n185 163.367
R1044 B.n734 B.n183 163.367
R1045 B.n738 B.n183 163.367
R1046 B.n738 B.n178 163.367
R1047 B.n747 B.n178 163.367
R1048 B.n747 B.n176 163.367
R1049 B.n751 B.n176 163.367
R1050 B.n751 B.n2 163.367
R1051 B.n1176 B.n2 163.367
R1052 B.n1176 B.n3 163.367
R1053 B.n1172 B.n3 163.367
R1054 B.n1172 B.n9 163.367
R1055 B.n1168 B.n9 163.367
R1056 B.n1168 B.n11 163.367
R1057 B.n1164 B.n11 163.367
R1058 B.n1164 B.n15 163.367
R1059 B.n1160 B.n15 163.367
R1060 B.n1160 B.n17 163.367
R1061 B.n1156 B.n17 163.367
R1062 B.n1156 B.n23 163.367
R1063 B.n1152 B.n23 163.367
R1064 B.n1152 B.n25 163.367
R1065 B.n1148 B.n25 163.367
R1066 B.n1148 B.n30 163.367
R1067 B.n1144 B.n30 163.367
R1068 B.n1144 B.n32 163.367
R1069 B.n1140 B.n32 163.367
R1070 B.n1140 B.n37 163.367
R1071 B.n1136 B.n37 163.367
R1072 B.n1136 B.n39 163.367
R1073 B.n1132 B.n39 163.367
R1074 B.n1132 B.n44 163.367
R1075 B.n1128 B.n44 163.367
R1076 B.n1128 B.n46 163.367
R1077 B.n1124 B.n46 163.367
R1078 B.n1124 B.n51 163.367
R1079 B.n1120 B.n51 163.367
R1080 B.n1120 B.n53 163.367
R1081 B.n1116 B.n53 163.367
R1082 B.n1116 B.n58 163.367
R1083 B.n1112 B.n58 163.367
R1084 B.n1112 B.n60 163.367
R1085 B.n1108 B.n60 163.367
R1086 B.n1108 B.n65 163.367
R1087 B.n1104 B.n65 163.367
R1088 B.n1104 B.n67 163.367
R1089 B.n1100 B.n67 163.367
R1090 B.n1100 B.n72 163.367
R1091 B.n1096 B.n72 163.367
R1092 B.n1096 B.n74 163.367
R1093 B.n1092 B.n74 163.367
R1094 B.n1092 B.n79 163.367
R1095 B.n1088 B.n79 163.367
R1096 B.n1088 B.n81 163.367
R1097 B.n1084 B.n81 163.367
R1098 B.n1084 B.n86 163.367
R1099 B.n1080 B.n86 163.367
R1100 B.n1080 B.n88 163.367
R1101 B.n1076 B.n88 163.367
R1102 B.n1076 B.n93 163.367
R1103 B.n1072 B.n93 163.367
R1104 B.n1072 B.n95 163.367
R1105 B.n1068 B.n95 163.367
R1106 B.n1068 B.n100 163.367
R1107 B.n1064 B.n100 163.367
R1108 B.n1064 B.n102 163.367
R1109 B.n1060 B.n102 163.367
R1110 B.n1060 B.n107 163.367
R1111 B.n1056 B.n107 163.367
R1112 B.n1056 B.n109 163.367
R1113 B.n1052 B.n109 163.367
R1114 B.n565 B.n563 163.367
R1115 B.n563 B.n562 163.367
R1116 B.n559 B.n558 163.367
R1117 B.n556 B.n299 163.367
R1118 B.n552 B.n550 163.367
R1119 B.n548 B.n301 163.367
R1120 B.n544 B.n542 163.367
R1121 B.n540 B.n303 163.367
R1122 B.n536 B.n534 163.367
R1123 B.n532 B.n305 163.367
R1124 B.n528 B.n526 163.367
R1125 B.n524 B.n307 163.367
R1126 B.n520 B.n518 163.367
R1127 B.n516 B.n309 163.367
R1128 B.n512 B.n510 163.367
R1129 B.n508 B.n311 163.367
R1130 B.n504 B.n502 163.367
R1131 B.n500 B.n313 163.367
R1132 B.n496 B.n494 163.367
R1133 B.n492 B.n315 163.367
R1134 B.n488 B.n486 163.367
R1135 B.n484 B.n317 163.367
R1136 B.n480 B.n478 163.367
R1137 B.n476 B.n319 163.367
R1138 B.n472 B.n470 163.367
R1139 B.n467 B.n466 163.367
R1140 B.n464 B.n325 163.367
R1141 B.n460 B.n458 163.367
R1142 B.n456 B.n327 163.367
R1143 B.n452 B.n450 163.367
R1144 B.n447 B.n446 163.367
R1145 B.n444 B.n333 163.367
R1146 B.n440 B.n438 163.367
R1147 B.n436 B.n335 163.367
R1148 B.n432 B.n430 163.367
R1149 B.n428 B.n337 163.367
R1150 B.n424 B.n422 163.367
R1151 B.n420 B.n339 163.367
R1152 B.n416 B.n414 163.367
R1153 B.n412 B.n341 163.367
R1154 B.n408 B.n406 163.367
R1155 B.n404 B.n343 163.367
R1156 B.n400 B.n398 163.367
R1157 B.n396 B.n345 163.367
R1158 B.n392 B.n390 163.367
R1159 B.n388 B.n347 163.367
R1160 B.n384 B.n382 163.367
R1161 B.n380 B.n349 163.367
R1162 B.n376 B.n374 163.367
R1163 B.n372 B.n351 163.367
R1164 B.n368 B.n366 163.367
R1165 B.n364 B.n353 163.367
R1166 B.n360 B.n358 163.367
R1167 B.n356 B.n293 163.367
R1168 B.n571 B.n291 163.367
R1169 B.n575 B.n291 163.367
R1170 B.n575 B.n285 163.367
R1171 B.n583 B.n285 163.367
R1172 B.n583 B.n283 163.367
R1173 B.n587 B.n283 163.367
R1174 B.n587 B.n277 163.367
R1175 B.n595 B.n277 163.367
R1176 B.n595 B.n275 163.367
R1177 B.n599 B.n275 163.367
R1178 B.n599 B.n269 163.367
R1179 B.n607 B.n269 163.367
R1180 B.n607 B.n267 163.367
R1181 B.n611 B.n267 163.367
R1182 B.n611 B.n261 163.367
R1183 B.n619 B.n261 163.367
R1184 B.n619 B.n259 163.367
R1185 B.n623 B.n259 163.367
R1186 B.n623 B.n253 163.367
R1187 B.n631 B.n253 163.367
R1188 B.n631 B.n251 163.367
R1189 B.n635 B.n251 163.367
R1190 B.n635 B.n245 163.367
R1191 B.n643 B.n245 163.367
R1192 B.n643 B.n243 163.367
R1193 B.n647 B.n243 163.367
R1194 B.n647 B.n237 163.367
R1195 B.n655 B.n237 163.367
R1196 B.n655 B.n235 163.367
R1197 B.n659 B.n235 163.367
R1198 B.n659 B.n228 163.367
R1199 B.n667 B.n228 163.367
R1200 B.n667 B.n226 163.367
R1201 B.n671 B.n226 163.367
R1202 B.n671 B.n221 163.367
R1203 B.n679 B.n221 163.367
R1204 B.n679 B.n219 163.367
R1205 B.n683 B.n219 163.367
R1206 B.n683 B.n213 163.367
R1207 B.n691 B.n213 163.367
R1208 B.n691 B.n211 163.367
R1209 B.n695 B.n211 163.367
R1210 B.n695 B.n205 163.367
R1211 B.n703 B.n205 163.367
R1212 B.n703 B.n203 163.367
R1213 B.n707 B.n203 163.367
R1214 B.n707 B.n197 163.367
R1215 B.n715 B.n197 163.367
R1216 B.n715 B.n195 163.367
R1217 B.n719 B.n195 163.367
R1218 B.n719 B.n189 163.367
R1219 B.n727 B.n189 163.367
R1220 B.n727 B.n187 163.367
R1221 B.n731 B.n187 163.367
R1222 B.n731 B.n182 163.367
R1223 B.n740 B.n182 163.367
R1224 B.n740 B.n180 163.367
R1225 B.n745 B.n180 163.367
R1226 B.n745 B.n174 163.367
R1227 B.n753 B.n174 163.367
R1228 B.n754 B.n753 163.367
R1229 B.n754 B.n5 163.367
R1230 B.n6 B.n5 163.367
R1231 B.n7 B.n6 163.367
R1232 B.n759 B.n7 163.367
R1233 B.n759 B.n12 163.367
R1234 B.n13 B.n12 163.367
R1235 B.n14 B.n13 163.367
R1236 B.n764 B.n14 163.367
R1237 B.n764 B.n19 163.367
R1238 B.n20 B.n19 163.367
R1239 B.n21 B.n20 163.367
R1240 B.n769 B.n21 163.367
R1241 B.n769 B.n26 163.367
R1242 B.n27 B.n26 163.367
R1243 B.n28 B.n27 163.367
R1244 B.n774 B.n28 163.367
R1245 B.n774 B.n33 163.367
R1246 B.n34 B.n33 163.367
R1247 B.n35 B.n34 163.367
R1248 B.n779 B.n35 163.367
R1249 B.n779 B.n40 163.367
R1250 B.n41 B.n40 163.367
R1251 B.n42 B.n41 163.367
R1252 B.n784 B.n42 163.367
R1253 B.n784 B.n47 163.367
R1254 B.n48 B.n47 163.367
R1255 B.n49 B.n48 163.367
R1256 B.n789 B.n49 163.367
R1257 B.n789 B.n54 163.367
R1258 B.n55 B.n54 163.367
R1259 B.n56 B.n55 163.367
R1260 B.n794 B.n56 163.367
R1261 B.n794 B.n61 163.367
R1262 B.n62 B.n61 163.367
R1263 B.n63 B.n62 163.367
R1264 B.n799 B.n63 163.367
R1265 B.n799 B.n68 163.367
R1266 B.n69 B.n68 163.367
R1267 B.n70 B.n69 163.367
R1268 B.n804 B.n70 163.367
R1269 B.n804 B.n75 163.367
R1270 B.n76 B.n75 163.367
R1271 B.n77 B.n76 163.367
R1272 B.n809 B.n77 163.367
R1273 B.n809 B.n82 163.367
R1274 B.n83 B.n82 163.367
R1275 B.n84 B.n83 163.367
R1276 B.n814 B.n84 163.367
R1277 B.n814 B.n89 163.367
R1278 B.n90 B.n89 163.367
R1279 B.n91 B.n90 163.367
R1280 B.n819 B.n91 163.367
R1281 B.n819 B.n96 163.367
R1282 B.n97 B.n96 163.367
R1283 B.n98 B.n97 163.367
R1284 B.n824 B.n98 163.367
R1285 B.n824 B.n103 163.367
R1286 B.n104 B.n103 163.367
R1287 B.n105 B.n104 163.367
R1288 B.n829 B.n105 163.367
R1289 B.n829 B.n110 163.367
R1290 B.n111 B.n110 163.367
R1291 B.n112 B.n111 163.367
R1292 B.n1048 B.n1046 163.367
R1293 B.n1044 B.n116 163.367
R1294 B.n1040 B.n1038 163.367
R1295 B.n1036 B.n118 163.367
R1296 B.n1032 B.n1030 163.367
R1297 B.n1028 B.n120 163.367
R1298 B.n1024 B.n1022 163.367
R1299 B.n1020 B.n122 163.367
R1300 B.n1016 B.n1014 163.367
R1301 B.n1012 B.n124 163.367
R1302 B.n1008 B.n1006 163.367
R1303 B.n1004 B.n126 163.367
R1304 B.n1000 B.n998 163.367
R1305 B.n996 B.n128 163.367
R1306 B.n992 B.n990 163.367
R1307 B.n988 B.n130 163.367
R1308 B.n984 B.n982 163.367
R1309 B.n980 B.n132 163.367
R1310 B.n976 B.n974 163.367
R1311 B.n972 B.n134 163.367
R1312 B.n968 B.n966 163.367
R1313 B.n964 B.n136 163.367
R1314 B.n960 B.n958 163.367
R1315 B.n956 B.n138 163.367
R1316 B.n951 B.n949 163.367
R1317 B.n947 B.n142 163.367
R1318 B.n943 B.n941 163.367
R1319 B.n939 B.n144 163.367
R1320 B.n935 B.n933 163.367
R1321 B.n931 B.n146 163.367
R1322 B.n927 B.n925 163.367
R1323 B.n923 B.n151 163.367
R1324 B.n919 B.n917 163.367
R1325 B.n915 B.n153 163.367
R1326 B.n911 B.n909 163.367
R1327 B.n907 B.n155 163.367
R1328 B.n903 B.n901 163.367
R1329 B.n899 B.n157 163.367
R1330 B.n895 B.n893 163.367
R1331 B.n891 B.n159 163.367
R1332 B.n887 B.n885 163.367
R1333 B.n883 B.n161 163.367
R1334 B.n879 B.n877 163.367
R1335 B.n875 B.n163 163.367
R1336 B.n871 B.n869 163.367
R1337 B.n867 B.n165 163.367
R1338 B.n863 B.n861 163.367
R1339 B.n859 B.n167 163.367
R1340 B.n855 B.n853 163.367
R1341 B.n851 B.n169 163.367
R1342 B.n847 B.n845 163.367
R1343 B.n843 B.n171 163.367
R1344 B.n839 B.n837 163.367
R1345 B.n328 B.t15 143.721
R1346 B.n147 B.t20 143.721
R1347 B.n320 B.t18 143.702
R1348 B.n139 B.t10 143.702
R1349 B.n329 B.t14 72.9336
R1350 B.n148 B.t21 72.9336
R1351 B.n321 B.t17 72.9149
R1352 B.n140 B.t11 72.9149
R1353 B.n564 B.n295 71.676
R1354 B.n562 B.n297 71.676
R1355 B.n558 B.n557 71.676
R1356 B.n551 B.n299 71.676
R1357 B.n550 B.n549 71.676
R1358 B.n543 B.n301 71.676
R1359 B.n542 B.n541 71.676
R1360 B.n535 B.n303 71.676
R1361 B.n534 B.n533 71.676
R1362 B.n527 B.n305 71.676
R1363 B.n526 B.n525 71.676
R1364 B.n519 B.n307 71.676
R1365 B.n518 B.n517 71.676
R1366 B.n511 B.n309 71.676
R1367 B.n510 B.n509 71.676
R1368 B.n503 B.n311 71.676
R1369 B.n502 B.n501 71.676
R1370 B.n495 B.n313 71.676
R1371 B.n494 B.n493 71.676
R1372 B.n487 B.n315 71.676
R1373 B.n486 B.n485 71.676
R1374 B.n479 B.n317 71.676
R1375 B.n478 B.n477 71.676
R1376 B.n471 B.n319 71.676
R1377 B.n470 B.n323 71.676
R1378 B.n466 B.n465 71.676
R1379 B.n459 B.n325 71.676
R1380 B.n458 B.n457 71.676
R1381 B.n451 B.n327 71.676
R1382 B.n450 B.n331 71.676
R1383 B.n446 B.n445 71.676
R1384 B.n439 B.n333 71.676
R1385 B.n438 B.n437 71.676
R1386 B.n431 B.n335 71.676
R1387 B.n430 B.n429 71.676
R1388 B.n423 B.n337 71.676
R1389 B.n422 B.n421 71.676
R1390 B.n415 B.n339 71.676
R1391 B.n414 B.n413 71.676
R1392 B.n407 B.n341 71.676
R1393 B.n406 B.n405 71.676
R1394 B.n399 B.n343 71.676
R1395 B.n398 B.n397 71.676
R1396 B.n391 B.n345 71.676
R1397 B.n390 B.n389 71.676
R1398 B.n383 B.n347 71.676
R1399 B.n382 B.n381 71.676
R1400 B.n375 B.n349 71.676
R1401 B.n374 B.n373 71.676
R1402 B.n367 B.n351 71.676
R1403 B.n366 B.n365 71.676
R1404 B.n359 B.n353 71.676
R1405 B.n358 B.n357 71.676
R1406 B.n1047 B.n114 71.676
R1407 B.n1046 B.n1045 71.676
R1408 B.n1039 B.n116 71.676
R1409 B.n1038 B.n1037 71.676
R1410 B.n1031 B.n118 71.676
R1411 B.n1030 B.n1029 71.676
R1412 B.n1023 B.n120 71.676
R1413 B.n1022 B.n1021 71.676
R1414 B.n1015 B.n122 71.676
R1415 B.n1014 B.n1013 71.676
R1416 B.n1007 B.n124 71.676
R1417 B.n1006 B.n1005 71.676
R1418 B.n999 B.n126 71.676
R1419 B.n998 B.n997 71.676
R1420 B.n991 B.n128 71.676
R1421 B.n990 B.n989 71.676
R1422 B.n983 B.n130 71.676
R1423 B.n982 B.n981 71.676
R1424 B.n975 B.n132 71.676
R1425 B.n974 B.n973 71.676
R1426 B.n967 B.n134 71.676
R1427 B.n966 B.n965 71.676
R1428 B.n959 B.n136 71.676
R1429 B.n958 B.n957 71.676
R1430 B.n950 B.n138 71.676
R1431 B.n949 B.n948 71.676
R1432 B.n942 B.n142 71.676
R1433 B.n941 B.n940 71.676
R1434 B.n934 B.n144 71.676
R1435 B.n933 B.n932 71.676
R1436 B.n926 B.n146 71.676
R1437 B.n925 B.n924 71.676
R1438 B.n918 B.n151 71.676
R1439 B.n917 B.n916 71.676
R1440 B.n910 B.n153 71.676
R1441 B.n909 B.n908 71.676
R1442 B.n902 B.n155 71.676
R1443 B.n901 B.n900 71.676
R1444 B.n894 B.n157 71.676
R1445 B.n893 B.n892 71.676
R1446 B.n886 B.n159 71.676
R1447 B.n885 B.n884 71.676
R1448 B.n878 B.n161 71.676
R1449 B.n877 B.n876 71.676
R1450 B.n870 B.n163 71.676
R1451 B.n869 B.n868 71.676
R1452 B.n862 B.n165 71.676
R1453 B.n861 B.n860 71.676
R1454 B.n854 B.n167 71.676
R1455 B.n853 B.n852 71.676
R1456 B.n846 B.n169 71.676
R1457 B.n845 B.n844 71.676
R1458 B.n838 B.n171 71.676
R1459 B.n837 B.n836 71.676
R1460 B.n836 B.n835 71.676
R1461 B.n839 B.n838 71.676
R1462 B.n844 B.n843 71.676
R1463 B.n847 B.n846 71.676
R1464 B.n852 B.n851 71.676
R1465 B.n855 B.n854 71.676
R1466 B.n860 B.n859 71.676
R1467 B.n863 B.n862 71.676
R1468 B.n868 B.n867 71.676
R1469 B.n871 B.n870 71.676
R1470 B.n876 B.n875 71.676
R1471 B.n879 B.n878 71.676
R1472 B.n884 B.n883 71.676
R1473 B.n887 B.n886 71.676
R1474 B.n892 B.n891 71.676
R1475 B.n895 B.n894 71.676
R1476 B.n900 B.n899 71.676
R1477 B.n903 B.n902 71.676
R1478 B.n908 B.n907 71.676
R1479 B.n911 B.n910 71.676
R1480 B.n916 B.n915 71.676
R1481 B.n919 B.n918 71.676
R1482 B.n924 B.n923 71.676
R1483 B.n927 B.n926 71.676
R1484 B.n932 B.n931 71.676
R1485 B.n935 B.n934 71.676
R1486 B.n940 B.n939 71.676
R1487 B.n943 B.n942 71.676
R1488 B.n948 B.n947 71.676
R1489 B.n951 B.n950 71.676
R1490 B.n957 B.n956 71.676
R1491 B.n960 B.n959 71.676
R1492 B.n965 B.n964 71.676
R1493 B.n968 B.n967 71.676
R1494 B.n973 B.n972 71.676
R1495 B.n976 B.n975 71.676
R1496 B.n981 B.n980 71.676
R1497 B.n984 B.n983 71.676
R1498 B.n989 B.n988 71.676
R1499 B.n992 B.n991 71.676
R1500 B.n997 B.n996 71.676
R1501 B.n1000 B.n999 71.676
R1502 B.n1005 B.n1004 71.676
R1503 B.n1008 B.n1007 71.676
R1504 B.n1013 B.n1012 71.676
R1505 B.n1016 B.n1015 71.676
R1506 B.n1021 B.n1020 71.676
R1507 B.n1024 B.n1023 71.676
R1508 B.n1029 B.n1028 71.676
R1509 B.n1032 B.n1031 71.676
R1510 B.n1037 B.n1036 71.676
R1511 B.n1040 B.n1039 71.676
R1512 B.n1045 B.n1044 71.676
R1513 B.n1048 B.n1047 71.676
R1514 B.n565 B.n564 71.676
R1515 B.n559 B.n297 71.676
R1516 B.n557 B.n556 71.676
R1517 B.n552 B.n551 71.676
R1518 B.n549 B.n548 71.676
R1519 B.n544 B.n543 71.676
R1520 B.n541 B.n540 71.676
R1521 B.n536 B.n535 71.676
R1522 B.n533 B.n532 71.676
R1523 B.n528 B.n527 71.676
R1524 B.n525 B.n524 71.676
R1525 B.n520 B.n519 71.676
R1526 B.n517 B.n516 71.676
R1527 B.n512 B.n511 71.676
R1528 B.n509 B.n508 71.676
R1529 B.n504 B.n503 71.676
R1530 B.n501 B.n500 71.676
R1531 B.n496 B.n495 71.676
R1532 B.n493 B.n492 71.676
R1533 B.n488 B.n487 71.676
R1534 B.n485 B.n484 71.676
R1535 B.n480 B.n479 71.676
R1536 B.n477 B.n476 71.676
R1537 B.n472 B.n471 71.676
R1538 B.n467 B.n323 71.676
R1539 B.n465 B.n464 71.676
R1540 B.n460 B.n459 71.676
R1541 B.n457 B.n456 71.676
R1542 B.n452 B.n451 71.676
R1543 B.n447 B.n331 71.676
R1544 B.n445 B.n444 71.676
R1545 B.n440 B.n439 71.676
R1546 B.n437 B.n436 71.676
R1547 B.n432 B.n431 71.676
R1548 B.n429 B.n428 71.676
R1549 B.n424 B.n423 71.676
R1550 B.n421 B.n420 71.676
R1551 B.n416 B.n415 71.676
R1552 B.n413 B.n412 71.676
R1553 B.n408 B.n407 71.676
R1554 B.n405 B.n404 71.676
R1555 B.n400 B.n399 71.676
R1556 B.n397 B.n396 71.676
R1557 B.n392 B.n391 71.676
R1558 B.n389 B.n388 71.676
R1559 B.n384 B.n383 71.676
R1560 B.n381 B.n380 71.676
R1561 B.n376 B.n375 71.676
R1562 B.n373 B.n372 71.676
R1563 B.n368 B.n367 71.676
R1564 B.n365 B.n364 71.676
R1565 B.n360 B.n359 71.676
R1566 B.n357 B.n356 71.676
R1567 B.n329 B.n328 70.7884
R1568 B.n321 B.n320 70.7884
R1569 B.n140 B.n139 70.7884
R1570 B.n148 B.n147 70.7884
R1571 B.n570 B.n294 60.4492
R1572 B.n1053 B.n113 60.4492
R1573 B.n330 B.n329 59.5399
R1574 B.n322 B.n321 59.5399
R1575 B.n953 B.n140 59.5399
R1576 B.n149 B.n148 59.5399
R1577 B.n570 B.n290 37.7116
R1578 B.n576 B.n290 37.7116
R1579 B.n576 B.n286 37.7116
R1580 B.n582 B.n286 37.7116
R1581 B.n582 B.n282 37.7116
R1582 B.n588 B.n282 37.7116
R1583 B.n588 B.n278 37.7116
R1584 B.n594 B.n278 37.7116
R1585 B.n600 B.n274 37.7116
R1586 B.n600 B.n270 37.7116
R1587 B.n606 B.n270 37.7116
R1588 B.n606 B.n266 37.7116
R1589 B.n612 B.n266 37.7116
R1590 B.n612 B.n262 37.7116
R1591 B.n618 B.n262 37.7116
R1592 B.n618 B.n258 37.7116
R1593 B.n624 B.n258 37.7116
R1594 B.n624 B.n254 37.7116
R1595 B.n630 B.n254 37.7116
R1596 B.n630 B.n250 37.7116
R1597 B.n636 B.n250 37.7116
R1598 B.n642 B.n246 37.7116
R1599 B.n642 B.n242 37.7116
R1600 B.n648 B.n242 37.7116
R1601 B.n648 B.n238 37.7116
R1602 B.n654 B.n238 37.7116
R1603 B.n654 B.n234 37.7116
R1604 B.n660 B.n234 37.7116
R1605 B.n660 B.n229 37.7116
R1606 B.n666 B.n229 37.7116
R1607 B.n666 B.n230 37.7116
R1608 B.n672 B.n222 37.7116
R1609 B.n678 B.n222 37.7116
R1610 B.n678 B.n218 37.7116
R1611 B.n684 B.n218 37.7116
R1612 B.n684 B.n214 37.7116
R1613 B.n690 B.n214 37.7116
R1614 B.n690 B.n210 37.7116
R1615 B.n696 B.n210 37.7116
R1616 B.n696 B.n206 37.7116
R1617 B.n702 B.n206 37.7116
R1618 B.n708 B.n202 37.7116
R1619 B.n708 B.n198 37.7116
R1620 B.n714 B.n198 37.7116
R1621 B.n714 B.n194 37.7116
R1622 B.n720 B.n194 37.7116
R1623 B.n720 B.n190 37.7116
R1624 B.n726 B.n190 37.7116
R1625 B.n726 B.n186 37.7116
R1626 B.n733 B.n186 37.7116
R1627 B.n733 B.n732 37.7116
R1628 B.n739 B.n179 37.7116
R1629 B.n746 B.n179 37.7116
R1630 B.n746 B.n175 37.7116
R1631 B.n752 B.n175 37.7116
R1632 B.n752 B.n4 37.7116
R1633 B.n1175 B.n4 37.7116
R1634 B.n1175 B.n1174 37.7116
R1635 B.n1174 B.n1173 37.7116
R1636 B.n1173 B.n8 37.7116
R1637 B.n1167 B.n8 37.7116
R1638 B.n1167 B.n1166 37.7116
R1639 B.n1166 B.n1165 37.7116
R1640 B.n1159 B.n18 37.7116
R1641 B.n1159 B.n1158 37.7116
R1642 B.n1158 B.n1157 37.7116
R1643 B.n1157 B.n22 37.7116
R1644 B.n1151 B.n22 37.7116
R1645 B.n1151 B.n1150 37.7116
R1646 B.n1150 B.n1149 37.7116
R1647 B.n1149 B.n29 37.7116
R1648 B.n1143 B.n29 37.7116
R1649 B.n1143 B.n1142 37.7116
R1650 B.n1141 B.n36 37.7116
R1651 B.n1135 B.n36 37.7116
R1652 B.n1135 B.n1134 37.7116
R1653 B.n1134 B.n1133 37.7116
R1654 B.n1133 B.n43 37.7116
R1655 B.n1127 B.n43 37.7116
R1656 B.n1127 B.n1126 37.7116
R1657 B.n1126 B.n1125 37.7116
R1658 B.n1125 B.n50 37.7116
R1659 B.n1119 B.n50 37.7116
R1660 B.n1118 B.n1117 37.7116
R1661 B.n1117 B.n57 37.7116
R1662 B.n1111 B.n57 37.7116
R1663 B.n1111 B.n1110 37.7116
R1664 B.n1110 B.n1109 37.7116
R1665 B.n1109 B.n64 37.7116
R1666 B.n1103 B.n64 37.7116
R1667 B.n1103 B.n1102 37.7116
R1668 B.n1102 B.n1101 37.7116
R1669 B.n1101 B.n71 37.7116
R1670 B.n1095 B.n1094 37.7116
R1671 B.n1094 B.n1093 37.7116
R1672 B.n1093 B.n78 37.7116
R1673 B.n1087 B.n78 37.7116
R1674 B.n1087 B.n1086 37.7116
R1675 B.n1086 B.n1085 37.7116
R1676 B.n1085 B.n85 37.7116
R1677 B.n1079 B.n85 37.7116
R1678 B.n1079 B.n1078 37.7116
R1679 B.n1078 B.n1077 37.7116
R1680 B.n1077 B.n92 37.7116
R1681 B.n1071 B.n92 37.7116
R1682 B.n1071 B.n1070 37.7116
R1683 B.n1069 B.n99 37.7116
R1684 B.n1063 B.n99 37.7116
R1685 B.n1063 B.n1062 37.7116
R1686 B.n1062 B.n1061 37.7116
R1687 B.n1061 B.n106 37.7116
R1688 B.n1055 B.n106 37.7116
R1689 B.n1055 B.n1054 37.7116
R1690 B.n1054 B.n1053 37.7116
R1691 B.n739 B.t6 36.6025
R1692 B.n1165 B.t0 36.6025
R1693 B.n594 B.t13 33.275
R1694 B.t9 B.n1069 33.275
R1695 B.n636 B.t5 31.0567
R1696 B.n1095 B.t4 31.0567
R1697 B.n1051 B.n1050 29.5029
R1698 B.n572 B.n292 29.5029
R1699 B.n568 B.n567 29.5029
R1700 B.n834 B.n833 29.5029
R1701 B.t2 B.n202 26.6201
R1702 B.n1142 B.t7 26.6201
R1703 B.n230 B.t3 21.0744
R1704 B.t1 B.n1118 21.0744
R1705 B B.n1177 18.0485
R1706 B.n672 B.t3 16.6378
R1707 B.n1119 B.t1 16.6378
R1708 B.n702 B.t2 11.092
R1709 B.t7 B.n1141 11.092
R1710 B.n1050 B.n1049 10.6151
R1711 B.n1049 B.n115 10.6151
R1712 B.n1043 B.n115 10.6151
R1713 B.n1043 B.n1042 10.6151
R1714 B.n1042 B.n1041 10.6151
R1715 B.n1041 B.n117 10.6151
R1716 B.n1035 B.n117 10.6151
R1717 B.n1035 B.n1034 10.6151
R1718 B.n1034 B.n1033 10.6151
R1719 B.n1033 B.n119 10.6151
R1720 B.n1027 B.n119 10.6151
R1721 B.n1027 B.n1026 10.6151
R1722 B.n1026 B.n1025 10.6151
R1723 B.n1025 B.n121 10.6151
R1724 B.n1019 B.n121 10.6151
R1725 B.n1019 B.n1018 10.6151
R1726 B.n1018 B.n1017 10.6151
R1727 B.n1017 B.n123 10.6151
R1728 B.n1011 B.n123 10.6151
R1729 B.n1011 B.n1010 10.6151
R1730 B.n1010 B.n1009 10.6151
R1731 B.n1009 B.n125 10.6151
R1732 B.n1003 B.n125 10.6151
R1733 B.n1003 B.n1002 10.6151
R1734 B.n1002 B.n1001 10.6151
R1735 B.n1001 B.n127 10.6151
R1736 B.n995 B.n127 10.6151
R1737 B.n995 B.n994 10.6151
R1738 B.n994 B.n993 10.6151
R1739 B.n993 B.n129 10.6151
R1740 B.n987 B.n129 10.6151
R1741 B.n987 B.n986 10.6151
R1742 B.n986 B.n985 10.6151
R1743 B.n985 B.n131 10.6151
R1744 B.n979 B.n131 10.6151
R1745 B.n979 B.n978 10.6151
R1746 B.n978 B.n977 10.6151
R1747 B.n977 B.n133 10.6151
R1748 B.n971 B.n133 10.6151
R1749 B.n971 B.n970 10.6151
R1750 B.n970 B.n969 10.6151
R1751 B.n969 B.n135 10.6151
R1752 B.n963 B.n135 10.6151
R1753 B.n963 B.n962 10.6151
R1754 B.n962 B.n961 10.6151
R1755 B.n961 B.n137 10.6151
R1756 B.n955 B.n137 10.6151
R1757 B.n955 B.n954 10.6151
R1758 B.n952 B.n141 10.6151
R1759 B.n946 B.n141 10.6151
R1760 B.n946 B.n945 10.6151
R1761 B.n945 B.n944 10.6151
R1762 B.n944 B.n143 10.6151
R1763 B.n938 B.n143 10.6151
R1764 B.n938 B.n937 10.6151
R1765 B.n937 B.n936 10.6151
R1766 B.n936 B.n145 10.6151
R1767 B.n930 B.n929 10.6151
R1768 B.n929 B.n928 10.6151
R1769 B.n928 B.n150 10.6151
R1770 B.n922 B.n150 10.6151
R1771 B.n922 B.n921 10.6151
R1772 B.n921 B.n920 10.6151
R1773 B.n920 B.n152 10.6151
R1774 B.n914 B.n152 10.6151
R1775 B.n914 B.n913 10.6151
R1776 B.n913 B.n912 10.6151
R1777 B.n912 B.n154 10.6151
R1778 B.n906 B.n154 10.6151
R1779 B.n906 B.n905 10.6151
R1780 B.n905 B.n904 10.6151
R1781 B.n904 B.n156 10.6151
R1782 B.n898 B.n156 10.6151
R1783 B.n898 B.n897 10.6151
R1784 B.n897 B.n896 10.6151
R1785 B.n896 B.n158 10.6151
R1786 B.n890 B.n158 10.6151
R1787 B.n890 B.n889 10.6151
R1788 B.n889 B.n888 10.6151
R1789 B.n888 B.n160 10.6151
R1790 B.n882 B.n160 10.6151
R1791 B.n882 B.n881 10.6151
R1792 B.n881 B.n880 10.6151
R1793 B.n880 B.n162 10.6151
R1794 B.n874 B.n162 10.6151
R1795 B.n874 B.n873 10.6151
R1796 B.n873 B.n872 10.6151
R1797 B.n872 B.n164 10.6151
R1798 B.n866 B.n164 10.6151
R1799 B.n866 B.n865 10.6151
R1800 B.n865 B.n864 10.6151
R1801 B.n864 B.n166 10.6151
R1802 B.n858 B.n166 10.6151
R1803 B.n858 B.n857 10.6151
R1804 B.n857 B.n856 10.6151
R1805 B.n856 B.n168 10.6151
R1806 B.n850 B.n168 10.6151
R1807 B.n850 B.n849 10.6151
R1808 B.n849 B.n848 10.6151
R1809 B.n848 B.n170 10.6151
R1810 B.n842 B.n170 10.6151
R1811 B.n842 B.n841 10.6151
R1812 B.n841 B.n840 10.6151
R1813 B.n840 B.n172 10.6151
R1814 B.n834 B.n172 10.6151
R1815 B.n573 B.n572 10.6151
R1816 B.n574 B.n573 10.6151
R1817 B.n574 B.n284 10.6151
R1818 B.n584 B.n284 10.6151
R1819 B.n585 B.n584 10.6151
R1820 B.n586 B.n585 10.6151
R1821 B.n586 B.n276 10.6151
R1822 B.n596 B.n276 10.6151
R1823 B.n597 B.n596 10.6151
R1824 B.n598 B.n597 10.6151
R1825 B.n598 B.n268 10.6151
R1826 B.n608 B.n268 10.6151
R1827 B.n609 B.n608 10.6151
R1828 B.n610 B.n609 10.6151
R1829 B.n610 B.n260 10.6151
R1830 B.n620 B.n260 10.6151
R1831 B.n621 B.n620 10.6151
R1832 B.n622 B.n621 10.6151
R1833 B.n622 B.n252 10.6151
R1834 B.n632 B.n252 10.6151
R1835 B.n633 B.n632 10.6151
R1836 B.n634 B.n633 10.6151
R1837 B.n634 B.n244 10.6151
R1838 B.n644 B.n244 10.6151
R1839 B.n645 B.n644 10.6151
R1840 B.n646 B.n645 10.6151
R1841 B.n646 B.n236 10.6151
R1842 B.n656 B.n236 10.6151
R1843 B.n657 B.n656 10.6151
R1844 B.n658 B.n657 10.6151
R1845 B.n658 B.n227 10.6151
R1846 B.n668 B.n227 10.6151
R1847 B.n669 B.n668 10.6151
R1848 B.n670 B.n669 10.6151
R1849 B.n670 B.n220 10.6151
R1850 B.n680 B.n220 10.6151
R1851 B.n681 B.n680 10.6151
R1852 B.n682 B.n681 10.6151
R1853 B.n682 B.n212 10.6151
R1854 B.n692 B.n212 10.6151
R1855 B.n693 B.n692 10.6151
R1856 B.n694 B.n693 10.6151
R1857 B.n694 B.n204 10.6151
R1858 B.n704 B.n204 10.6151
R1859 B.n705 B.n704 10.6151
R1860 B.n706 B.n705 10.6151
R1861 B.n706 B.n196 10.6151
R1862 B.n716 B.n196 10.6151
R1863 B.n717 B.n716 10.6151
R1864 B.n718 B.n717 10.6151
R1865 B.n718 B.n188 10.6151
R1866 B.n728 B.n188 10.6151
R1867 B.n729 B.n728 10.6151
R1868 B.n730 B.n729 10.6151
R1869 B.n730 B.n181 10.6151
R1870 B.n741 B.n181 10.6151
R1871 B.n742 B.n741 10.6151
R1872 B.n744 B.n742 10.6151
R1873 B.n744 B.n743 10.6151
R1874 B.n743 B.n173 10.6151
R1875 B.n755 B.n173 10.6151
R1876 B.n756 B.n755 10.6151
R1877 B.n757 B.n756 10.6151
R1878 B.n758 B.n757 10.6151
R1879 B.n760 B.n758 10.6151
R1880 B.n761 B.n760 10.6151
R1881 B.n762 B.n761 10.6151
R1882 B.n763 B.n762 10.6151
R1883 B.n765 B.n763 10.6151
R1884 B.n766 B.n765 10.6151
R1885 B.n767 B.n766 10.6151
R1886 B.n768 B.n767 10.6151
R1887 B.n770 B.n768 10.6151
R1888 B.n771 B.n770 10.6151
R1889 B.n772 B.n771 10.6151
R1890 B.n773 B.n772 10.6151
R1891 B.n775 B.n773 10.6151
R1892 B.n776 B.n775 10.6151
R1893 B.n777 B.n776 10.6151
R1894 B.n778 B.n777 10.6151
R1895 B.n780 B.n778 10.6151
R1896 B.n781 B.n780 10.6151
R1897 B.n782 B.n781 10.6151
R1898 B.n783 B.n782 10.6151
R1899 B.n785 B.n783 10.6151
R1900 B.n786 B.n785 10.6151
R1901 B.n787 B.n786 10.6151
R1902 B.n788 B.n787 10.6151
R1903 B.n790 B.n788 10.6151
R1904 B.n791 B.n790 10.6151
R1905 B.n792 B.n791 10.6151
R1906 B.n793 B.n792 10.6151
R1907 B.n795 B.n793 10.6151
R1908 B.n796 B.n795 10.6151
R1909 B.n797 B.n796 10.6151
R1910 B.n798 B.n797 10.6151
R1911 B.n800 B.n798 10.6151
R1912 B.n801 B.n800 10.6151
R1913 B.n802 B.n801 10.6151
R1914 B.n803 B.n802 10.6151
R1915 B.n805 B.n803 10.6151
R1916 B.n806 B.n805 10.6151
R1917 B.n807 B.n806 10.6151
R1918 B.n808 B.n807 10.6151
R1919 B.n810 B.n808 10.6151
R1920 B.n811 B.n810 10.6151
R1921 B.n812 B.n811 10.6151
R1922 B.n813 B.n812 10.6151
R1923 B.n815 B.n813 10.6151
R1924 B.n816 B.n815 10.6151
R1925 B.n817 B.n816 10.6151
R1926 B.n818 B.n817 10.6151
R1927 B.n820 B.n818 10.6151
R1928 B.n821 B.n820 10.6151
R1929 B.n822 B.n821 10.6151
R1930 B.n823 B.n822 10.6151
R1931 B.n825 B.n823 10.6151
R1932 B.n826 B.n825 10.6151
R1933 B.n827 B.n826 10.6151
R1934 B.n828 B.n827 10.6151
R1935 B.n830 B.n828 10.6151
R1936 B.n831 B.n830 10.6151
R1937 B.n832 B.n831 10.6151
R1938 B.n833 B.n832 10.6151
R1939 B.n567 B.n566 10.6151
R1940 B.n566 B.n296 10.6151
R1941 B.n561 B.n296 10.6151
R1942 B.n561 B.n560 10.6151
R1943 B.n560 B.n298 10.6151
R1944 B.n555 B.n298 10.6151
R1945 B.n555 B.n554 10.6151
R1946 B.n554 B.n553 10.6151
R1947 B.n553 B.n300 10.6151
R1948 B.n547 B.n300 10.6151
R1949 B.n547 B.n546 10.6151
R1950 B.n546 B.n545 10.6151
R1951 B.n545 B.n302 10.6151
R1952 B.n539 B.n302 10.6151
R1953 B.n539 B.n538 10.6151
R1954 B.n538 B.n537 10.6151
R1955 B.n537 B.n304 10.6151
R1956 B.n531 B.n304 10.6151
R1957 B.n531 B.n530 10.6151
R1958 B.n530 B.n529 10.6151
R1959 B.n529 B.n306 10.6151
R1960 B.n523 B.n306 10.6151
R1961 B.n523 B.n522 10.6151
R1962 B.n522 B.n521 10.6151
R1963 B.n521 B.n308 10.6151
R1964 B.n515 B.n308 10.6151
R1965 B.n515 B.n514 10.6151
R1966 B.n514 B.n513 10.6151
R1967 B.n513 B.n310 10.6151
R1968 B.n507 B.n310 10.6151
R1969 B.n507 B.n506 10.6151
R1970 B.n506 B.n505 10.6151
R1971 B.n505 B.n312 10.6151
R1972 B.n499 B.n312 10.6151
R1973 B.n499 B.n498 10.6151
R1974 B.n498 B.n497 10.6151
R1975 B.n497 B.n314 10.6151
R1976 B.n491 B.n314 10.6151
R1977 B.n491 B.n490 10.6151
R1978 B.n490 B.n489 10.6151
R1979 B.n489 B.n316 10.6151
R1980 B.n483 B.n316 10.6151
R1981 B.n483 B.n482 10.6151
R1982 B.n482 B.n481 10.6151
R1983 B.n481 B.n318 10.6151
R1984 B.n475 B.n318 10.6151
R1985 B.n475 B.n474 10.6151
R1986 B.n474 B.n473 10.6151
R1987 B.n469 B.n468 10.6151
R1988 B.n468 B.n324 10.6151
R1989 B.n463 B.n324 10.6151
R1990 B.n463 B.n462 10.6151
R1991 B.n462 B.n461 10.6151
R1992 B.n461 B.n326 10.6151
R1993 B.n455 B.n326 10.6151
R1994 B.n455 B.n454 10.6151
R1995 B.n454 B.n453 10.6151
R1996 B.n449 B.n448 10.6151
R1997 B.n448 B.n332 10.6151
R1998 B.n443 B.n332 10.6151
R1999 B.n443 B.n442 10.6151
R2000 B.n442 B.n441 10.6151
R2001 B.n441 B.n334 10.6151
R2002 B.n435 B.n334 10.6151
R2003 B.n435 B.n434 10.6151
R2004 B.n434 B.n433 10.6151
R2005 B.n433 B.n336 10.6151
R2006 B.n427 B.n336 10.6151
R2007 B.n427 B.n426 10.6151
R2008 B.n426 B.n425 10.6151
R2009 B.n425 B.n338 10.6151
R2010 B.n419 B.n338 10.6151
R2011 B.n419 B.n418 10.6151
R2012 B.n418 B.n417 10.6151
R2013 B.n417 B.n340 10.6151
R2014 B.n411 B.n340 10.6151
R2015 B.n411 B.n410 10.6151
R2016 B.n410 B.n409 10.6151
R2017 B.n409 B.n342 10.6151
R2018 B.n403 B.n342 10.6151
R2019 B.n403 B.n402 10.6151
R2020 B.n402 B.n401 10.6151
R2021 B.n401 B.n344 10.6151
R2022 B.n395 B.n344 10.6151
R2023 B.n395 B.n394 10.6151
R2024 B.n394 B.n393 10.6151
R2025 B.n393 B.n346 10.6151
R2026 B.n387 B.n346 10.6151
R2027 B.n387 B.n386 10.6151
R2028 B.n386 B.n385 10.6151
R2029 B.n385 B.n348 10.6151
R2030 B.n379 B.n348 10.6151
R2031 B.n379 B.n378 10.6151
R2032 B.n378 B.n377 10.6151
R2033 B.n377 B.n350 10.6151
R2034 B.n371 B.n350 10.6151
R2035 B.n371 B.n370 10.6151
R2036 B.n370 B.n369 10.6151
R2037 B.n369 B.n352 10.6151
R2038 B.n363 B.n352 10.6151
R2039 B.n363 B.n362 10.6151
R2040 B.n362 B.n361 10.6151
R2041 B.n361 B.n354 10.6151
R2042 B.n355 B.n354 10.6151
R2043 B.n355 B.n292 10.6151
R2044 B.n568 B.n288 10.6151
R2045 B.n578 B.n288 10.6151
R2046 B.n579 B.n578 10.6151
R2047 B.n580 B.n579 10.6151
R2048 B.n580 B.n280 10.6151
R2049 B.n590 B.n280 10.6151
R2050 B.n591 B.n590 10.6151
R2051 B.n592 B.n591 10.6151
R2052 B.n592 B.n272 10.6151
R2053 B.n602 B.n272 10.6151
R2054 B.n603 B.n602 10.6151
R2055 B.n604 B.n603 10.6151
R2056 B.n604 B.n264 10.6151
R2057 B.n614 B.n264 10.6151
R2058 B.n615 B.n614 10.6151
R2059 B.n616 B.n615 10.6151
R2060 B.n616 B.n256 10.6151
R2061 B.n626 B.n256 10.6151
R2062 B.n627 B.n626 10.6151
R2063 B.n628 B.n627 10.6151
R2064 B.n628 B.n248 10.6151
R2065 B.n638 B.n248 10.6151
R2066 B.n639 B.n638 10.6151
R2067 B.n640 B.n639 10.6151
R2068 B.n640 B.n240 10.6151
R2069 B.n650 B.n240 10.6151
R2070 B.n651 B.n650 10.6151
R2071 B.n652 B.n651 10.6151
R2072 B.n652 B.n232 10.6151
R2073 B.n662 B.n232 10.6151
R2074 B.n663 B.n662 10.6151
R2075 B.n664 B.n663 10.6151
R2076 B.n664 B.n224 10.6151
R2077 B.n674 B.n224 10.6151
R2078 B.n675 B.n674 10.6151
R2079 B.n676 B.n675 10.6151
R2080 B.n676 B.n216 10.6151
R2081 B.n686 B.n216 10.6151
R2082 B.n687 B.n686 10.6151
R2083 B.n688 B.n687 10.6151
R2084 B.n688 B.n208 10.6151
R2085 B.n698 B.n208 10.6151
R2086 B.n699 B.n698 10.6151
R2087 B.n700 B.n699 10.6151
R2088 B.n700 B.n200 10.6151
R2089 B.n710 B.n200 10.6151
R2090 B.n711 B.n710 10.6151
R2091 B.n712 B.n711 10.6151
R2092 B.n712 B.n192 10.6151
R2093 B.n722 B.n192 10.6151
R2094 B.n723 B.n722 10.6151
R2095 B.n724 B.n723 10.6151
R2096 B.n724 B.n184 10.6151
R2097 B.n735 B.n184 10.6151
R2098 B.n736 B.n735 10.6151
R2099 B.n737 B.n736 10.6151
R2100 B.n737 B.n177 10.6151
R2101 B.n748 B.n177 10.6151
R2102 B.n749 B.n748 10.6151
R2103 B.n750 B.n749 10.6151
R2104 B.n750 B.n0 10.6151
R2105 B.n1171 B.n1 10.6151
R2106 B.n1171 B.n1170 10.6151
R2107 B.n1170 B.n1169 10.6151
R2108 B.n1169 B.n10 10.6151
R2109 B.n1163 B.n10 10.6151
R2110 B.n1163 B.n1162 10.6151
R2111 B.n1162 B.n1161 10.6151
R2112 B.n1161 B.n16 10.6151
R2113 B.n1155 B.n16 10.6151
R2114 B.n1155 B.n1154 10.6151
R2115 B.n1154 B.n1153 10.6151
R2116 B.n1153 B.n24 10.6151
R2117 B.n1147 B.n24 10.6151
R2118 B.n1147 B.n1146 10.6151
R2119 B.n1146 B.n1145 10.6151
R2120 B.n1145 B.n31 10.6151
R2121 B.n1139 B.n31 10.6151
R2122 B.n1139 B.n1138 10.6151
R2123 B.n1138 B.n1137 10.6151
R2124 B.n1137 B.n38 10.6151
R2125 B.n1131 B.n38 10.6151
R2126 B.n1131 B.n1130 10.6151
R2127 B.n1130 B.n1129 10.6151
R2128 B.n1129 B.n45 10.6151
R2129 B.n1123 B.n45 10.6151
R2130 B.n1123 B.n1122 10.6151
R2131 B.n1122 B.n1121 10.6151
R2132 B.n1121 B.n52 10.6151
R2133 B.n1115 B.n52 10.6151
R2134 B.n1115 B.n1114 10.6151
R2135 B.n1114 B.n1113 10.6151
R2136 B.n1113 B.n59 10.6151
R2137 B.n1107 B.n59 10.6151
R2138 B.n1107 B.n1106 10.6151
R2139 B.n1106 B.n1105 10.6151
R2140 B.n1105 B.n66 10.6151
R2141 B.n1099 B.n66 10.6151
R2142 B.n1099 B.n1098 10.6151
R2143 B.n1098 B.n1097 10.6151
R2144 B.n1097 B.n73 10.6151
R2145 B.n1091 B.n73 10.6151
R2146 B.n1091 B.n1090 10.6151
R2147 B.n1090 B.n1089 10.6151
R2148 B.n1089 B.n80 10.6151
R2149 B.n1083 B.n80 10.6151
R2150 B.n1083 B.n1082 10.6151
R2151 B.n1082 B.n1081 10.6151
R2152 B.n1081 B.n87 10.6151
R2153 B.n1075 B.n87 10.6151
R2154 B.n1075 B.n1074 10.6151
R2155 B.n1074 B.n1073 10.6151
R2156 B.n1073 B.n94 10.6151
R2157 B.n1067 B.n94 10.6151
R2158 B.n1067 B.n1066 10.6151
R2159 B.n1066 B.n1065 10.6151
R2160 B.n1065 B.n101 10.6151
R2161 B.n1059 B.n101 10.6151
R2162 B.n1059 B.n1058 10.6151
R2163 B.n1058 B.n1057 10.6151
R2164 B.n1057 B.n108 10.6151
R2165 B.n1051 B.n108 10.6151
R2166 B.n954 B.n953 9.36635
R2167 B.n930 B.n149 9.36635
R2168 B.n473 B.n322 9.36635
R2169 B.n449 B.n330 9.36635
R2170 B.t5 B.n246 6.6554
R2171 B.t4 B.n71 6.6554
R2172 B.t13 B.n274 4.4371
R2173 B.n1070 B.t9 4.4371
R2174 B.n1177 B.n0 2.81026
R2175 B.n1177 B.n1 2.81026
R2176 B.n953 B.n952 1.24928
R2177 B.n149 B.n145 1.24928
R2178 B.n469 B.n322 1.24928
R2179 B.n453 B.n330 1.24928
R2180 B.n732 B.t6 1.10965
R2181 B.n18 B.t0 1.10965
R2182 VP.n24 VP.n21 161.3
R2183 VP.n26 VP.n25 161.3
R2184 VP.n27 VP.n20 161.3
R2185 VP.n29 VP.n28 161.3
R2186 VP.n30 VP.n19 161.3
R2187 VP.n32 VP.n31 161.3
R2188 VP.n33 VP.n18 161.3
R2189 VP.n35 VP.n34 161.3
R2190 VP.n37 VP.n36 161.3
R2191 VP.n38 VP.n16 161.3
R2192 VP.n40 VP.n39 161.3
R2193 VP.n41 VP.n15 161.3
R2194 VP.n43 VP.n42 161.3
R2195 VP.n44 VP.n14 161.3
R2196 VP.n46 VP.n45 161.3
R2197 VP.n83 VP.n82 161.3
R2198 VP.n81 VP.n1 161.3
R2199 VP.n80 VP.n79 161.3
R2200 VP.n78 VP.n2 161.3
R2201 VP.n77 VP.n76 161.3
R2202 VP.n75 VP.n3 161.3
R2203 VP.n74 VP.n73 161.3
R2204 VP.n72 VP.n71 161.3
R2205 VP.n70 VP.n5 161.3
R2206 VP.n69 VP.n68 161.3
R2207 VP.n67 VP.n6 161.3
R2208 VP.n66 VP.n65 161.3
R2209 VP.n64 VP.n7 161.3
R2210 VP.n63 VP.n62 161.3
R2211 VP.n61 VP.n8 161.3
R2212 VP.n60 VP.n59 161.3
R2213 VP.n57 VP.n9 161.3
R2214 VP.n56 VP.n55 161.3
R2215 VP.n54 VP.n10 161.3
R2216 VP.n53 VP.n52 161.3
R2217 VP.n51 VP.n11 161.3
R2218 VP.n50 VP.n49 161.3
R2219 VP.n23 VP.t2 137.915
R2220 VP.n12 VP.t5 105.692
R2221 VP.n58 VP.t7 105.692
R2222 VP.n4 VP.t1 105.692
R2223 VP.n0 VP.t6 105.692
R2224 VP.n13 VP.t3 105.692
R2225 VP.n17 VP.t0 105.692
R2226 VP.n22 VP.t4 105.692
R2227 VP.n48 VP.n12 78.9365
R2228 VP.n84 VP.n0 78.9365
R2229 VP.n47 VP.n13 78.9365
R2230 VP.n23 VP.n22 70.7064
R2231 VP.n65 VP.n6 56.4773
R2232 VP.n28 VP.n19 56.4773
R2233 VP.n48 VP.n47 56.2643
R2234 VP.n56 VP.n10 50.148
R2235 VP.n76 VP.n2 50.148
R2236 VP.n39 VP.n15 50.148
R2237 VP.n52 VP.n10 30.6732
R2238 VP.n80 VP.n2 30.6732
R2239 VP.n43 VP.n15 30.6732
R2240 VP.n51 VP.n50 24.3439
R2241 VP.n52 VP.n51 24.3439
R2242 VP.n57 VP.n56 24.3439
R2243 VP.n59 VP.n57 24.3439
R2244 VP.n63 VP.n8 24.3439
R2245 VP.n64 VP.n63 24.3439
R2246 VP.n65 VP.n64 24.3439
R2247 VP.n69 VP.n6 24.3439
R2248 VP.n70 VP.n69 24.3439
R2249 VP.n71 VP.n70 24.3439
R2250 VP.n75 VP.n74 24.3439
R2251 VP.n76 VP.n75 24.3439
R2252 VP.n81 VP.n80 24.3439
R2253 VP.n82 VP.n81 24.3439
R2254 VP.n44 VP.n43 24.3439
R2255 VP.n45 VP.n44 24.3439
R2256 VP.n32 VP.n19 24.3439
R2257 VP.n33 VP.n32 24.3439
R2258 VP.n34 VP.n33 24.3439
R2259 VP.n38 VP.n37 24.3439
R2260 VP.n39 VP.n38 24.3439
R2261 VP.n26 VP.n21 24.3439
R2262 VP.n27 VP.n26 24.3439
R2263 VP.n28 VP.n27 24.3439
R2264 VP.n59 VP.n58 20.6924
R2265 VP.n74 VP.n4 20.6924
R2266 VP.n37 VP.n17 20.6924
R2267 VP.n50 VP.n12 10.955
R2268 VP.n82 VP.n0 10.955
R2269 VP.n45 VP.n13 10.955
R2270 VP.n24 VP.n23 4.36821
R2271 VP.n58 VP.n8 3.65202
R2272 VP.n71 VP.n4 3.65202
R2273 VP.n34 VP.n17 3.65202
R2274 VP.n22 VP.n21 3.65202
R2275 VP.n47 VP.n46 0.355081
R2276 VP.n49 VP.n48 0.355081
R2277 VP.n84 VP.n83 0.355081
R2278 VP VP.n84 0.26685
R2279 VP.n25 VP.n24 0.189894
R2280 VP.n25 VP.n20 0.189894
R2281 VP.n29 VP.n20 0.189894
R2282 VP.n30 VP.n29 0.189894
R2283 VP.n31 VP.n30 0.189894
R2284 VP.n31 VP.n18 0.189894
R2285 VP.n35 VP.n18 0.189894
R2286 VP.n36 VP.n35 0.189894
R2287 VP.n36 VP.n16 0.189894
R2288 VP.n40 VP.n16 0.189894
R2289 VP.n41 VP.n40 0.189894
R2290 VP.n42 VP.n41 0.189894
R2291 VP.n42 VP.n14 0.189894
R2292 VP.n46 VP.n14 0.189894
R2293 VP.n49 VP.n11 0.189894
R2294 VP.n53 VP.n11 0.189894
R2295 VP.n54 VP.n53 0.189894
R2296 VP.n55 VP.n54 0.189894
R2297 VP.n55 VP.n9 0.189894
R2298 VP.n60 VP.n9 0.189894
R2299 VP.n61 VP.n60 0.189894
R2300 VP.n62 VP.n61 0.189894
R2301 VP.n62 VP.n7 0.189894
R2302 VP.n66 VP.n7 0.189894
R2303 VP.n67 VP.n66 0.189894
R2304 VP.n68 VP.n67 0.189894
R2305 VP.n68 VP.n5 0.189894
R2306 VP.n72 VP.n5 0.189894
R2307 VP.n73 VP.n72 0.189894
R2308 VP.n73 VP.n3 0.189894
R2309 VP.n77 VP.n3 0.189894
R2310 VP.n78 VP.n77 0.189894
R2311 VP.n79 VP.n78 0.189894
R2312 VP.n79 VP.n1 0.189894
R2313 VP.n83 VP.n1 0.189894
R2314 VDD1 VDD1.n0 61.4524
R2315 VDD1.n3 VDD1.n2 61.3389
R2316 VDD1.n3 VDD1.n1 61.3389
R2317 VDD1.n5 VDD1.n4 59.821
R2318 VDD1.n5 VDD1.n3 51.0095
R2319 VDD1 VDD1.n5 1.51559
R2320 VDD1.n4 VDD1.t7 1.36039
R2321 VDD1.n4 VDD1.t4 1.36039
R2322 VDD1.n0 VDD1.t5 1.36039
R2323 VDD1.n0 VDD1.t3 1.36039
R2324 VDD1.n2 VDD1.t6 1.36039
R2325 VDD1.n2 VDD1.t1 1.36039
R2326 VDD1.n1 VDD1.t2 1.36039
R2327 VDD1.n1 VDD1.t0 1.36039
C0 VDD1 VN 0.15258f
C1 VDD1 VP 11.355f
C2 VDD1 VDD2 2.14903f
C3 VTAIL VN 11.4279f
C4 VTAIL VP 11.441999f
C5 VTAIL VDD2 9.15204f
C6 VP VN 9.02751f
C7 VDD2 VN 10.9135f
C8 VTAIL VDD1 9.092791f
C9 VP VDD2 0.595836f
C10 VDD2 B 6.321f
C11 VDD1 B 6.836056f
C12 VTAIL B 12.523211f
C13 VN B 18.488192f
C14 VP B 17.107962f
C15 VDD1.t5 B 0.311106f
C16 VDD1.t3 B 0.311106f
C17 VDD1.n0 B 2.81687f
C18 VDD1.t2 B 0.311106f
C19 VDD1.t0 B 0.311106f
C20 VDD1.n1 B 2.81545f
C21 VDD1.t6 B 0.311106f
C22 VDD1.t1 B 0.311106f
C23 VDD1.n2 B 2.81545f
C24 VDD1.n3 B 4.23891f
C25 VDD1.t7 B 0.311106f
C26 VDD1.t4 B 0.311106f
C27 VDD1.n4 B 2.79943f
C28 VDD1.n5 B 3.71156f
C29 VP.t6 B 2.46883f
C30 VP.n0 B 0.929562f
C31 VP.n1 B 0.018651f
C32 VP.n2 B 0.017655f
C33 VP.n3 B 0.018651f
C34 VP.t1 B 2.46883f
C35 VP.n4 B 0.859473f
C36 VP.n5 B 0.018651f
C37 VP.n6 B 0.027346f
C38 VP.n7 B 0.018651f
C39 VP.n8 B 0.020274f
C40 VP.n9 B 0.018651f
C41 VP.n10 B 0.017655f
C42 VP.n11 B 0.018651f
C43 VP.t5 B 2.46883f
C44 VP.n12 B 0.929562f
C45 VP.t3 B 2.46883f
C46 VP.n13 B 0.929562f
C47 VP.n14 B 0.018651f
C48 VP.n15 B 0.017655f
C49 VP.n16 B 0.018651f
C50 VP.t0 B 2.46883f
C51 VP.n17 B 0.859473f
C52 VP.n18 B 0.018651f
C53 VP.n19 B 0.027346f
C54 VP.n20 B 0.018651f
C55 VP.n21 B 0.020274f
C56 VP.t2 B 2.70051f
C57 VP.t4 B 2.46883f
C58 VP.n22 B 0.917173f
C59 VP.n23 B 0.881143f
C60 VP.n24 B 0.220872f
C61 VP.n25 B 0.018651f
C62 VP.n26 B 0.034936f
C63 VP.n27 B 0.034936f
C64 VP.n28 B 0.027346f
C65 VP.n29 B 0.018651f
C66 VP.n30 B 0.018651f
C67 VP.n31 B 0.018651f
C68 VP.n32 B 0.034936f
C69 VP.n33 B 0.034936f
C70 VP.n34 B 0.020274f
C71 VP.n35 B 0.018651f
C72 VP.n36 B 0.018651f
C73 VP.n37 B 0.032348f
C74 VP.n38 B 0.034936f
C75 VP.n39 B 0.034403f
C76 VP.n40 B 0.018651f
C77 VP.n41 B 0.018651f
C78 VP.n42 B 0.018651f
C79 VP.n43 B 0.037569f
C80 VP.n44 B 0.034936f
C81 VP.n45 B 0.025449f
C82 VP.n46 B 0.030108f
C83 VP.n47 B 1.25399f
C84 VP.n48 B 1.26588f
C85 VP.n49 B 0.030108f
C86 VP.n50 B 0.025449f
C87 VP.n51 B 0.034936f
C88 VP.n52 B 0.037569f
C89 VP.n53 B 0.018651f
C90 VP.n54 B 0.018651f
C91 VP.n55 B 0.018651f
C92 VP.n56 B 0.034403f
C93 VP.n57 B 0.034936f
C94 VP.t7 B 2.46883f
C95 VP.n58 B 0.859473f
C96 VP.n59 B 0.032348f
C97 VP.n60 B 0.018651f
C98 VP.n61 B 0.018651f
C99 VP.n62 B 0.018651f
C100 VP.n63 B 0.034936f
C101 VP.n64 B 0.034936f
C102 VP.n65 B 0.027346f
C103 VP.n66 B 0.018651f
C104 VP.n67 B 0.018651f
C105 VP.n68 B 0.018651f
C106 VP.n69 B 0.034936f
C107 VP.n70 B 0.034936f
C108 VP.n71 B 0.020274f
C109 VP.n72 B 0.018651f
C110 VP.n73 B 0.018651f
C111 VP.n74 B 0.032348f
C112 VP.n75 B 0.034936f
C113 VP.n76 B 0.034403f
C114 VP.n77 B 0.018651f
C115 VP.n78 B 0.018651f
C116 VP.n79 B 0.018651f
C117 VP.n80 B 0.037569f
C118 VP.n81 B 0.034936f
C119 VP.n82 B 0.025449f
C120 VP.n83 B 0.030108f
C121 VP.n84 B 0.047912f
C122 VTAIL.t10 B 0.225614f
C123 VTAIL.t13 B 0.225614f
C124 VTAIL.n0 B 1.96722f
C125 VTAIL.n1 B 0.405262f
C126 VTAIL.t6 B 2.5105f
C127 VTAIL.n2 B 0.503301f
C128 VTAIL.t14 B 2.5105f
C129 VTAIL.n3 B 0.503301f
C130 VTAIL.t3 B 0.225614f
C131 VTAIL.t2 B 0.225614f
C132 VTAIL.n4 B 1.96722f
C133 VTAIL.n5 B 0.600397f
C134 VTAIL.t5 B 2.5105f
C135 VTAIL.n6 B 1.73186f
C136 VTAIL.t12 B 2.51051f
C137 VTAIL.n7 B 1.73185f
C138 VTAIL.t11 B 0.225614f
C139 VTAIL.t7 B 0.225614f
C140 VTAIL.n8 B 1.96722f
C141 VTAIL.n9 B 0.600398f
C142 VTAIL.t9 B 2.51051f
C143 VTAIL.n10 B 0.503295f
C144 VTAIL.t0 B 2.51051f
C145 VTAIL.n11 B 0.503295f
C146 VTAIL.t15 B 0.225614f
C147 VTAIL.t1 B 0.225614f
C148 VTAIL.n12 B 1.96722f
C149 VTAIL.n13 B 0.600398f
C150 VTAIL.t4 B 2.51051f
C151 VTAIL.n14 B 1.73185f
C152 VTAIL.t8 B 2.5105f
C153 VTAIL.n15 B 1.72818f
C154 VDD2.t4 B 0.306956f
C155 VDD2.t0 B 0.306956f
C156 VDD2.n0 B 2.7779f
C157 VDD2.t7 B 0.306956f
C158 VDD2.t2 B 0.306956f
C159 VDD2.n1 B 2.7779f
C160 VDD2.n2 B 4.1273f
C161 VDD2.t6 B 0.306956f
C162 VDD2.t1 B 0.306956f
C163 VDD2.n3 B 2.76209f
C164 VDD2.n4 B 3.62858f
C165 VDD2.t5 B 0.306956f
C166 VDD2.t3 B 0.306956f
C167 VDD2.n5 B 2.77785f
C168 VN.t5 B 2.42801f
C169 VN.n0 B 0.914192f
C170 VN.n1 B 0.018343f
C171 VN.n2 B 0.017363f
C172 VN.n3 B 0.018343f
C173 VN.t0 B 2.42801f
C174 VN.n4 B 0.845262f
C175 VN.n5 B 0.018343f
C176 VN.n6 B 0.026894f
C177 VN.n7 B 0.018343f
C178 VN.n8 B 0.019939f
C179 VN.t3 B 2.42801f
C180 VN.n9 B 0.902008f
C181 VN.t7 B 2.65586f
C182 VN.n10 B 0.866573f
C183 VN.n11 B 0.21722f
C184 VN.n12 B 0.018343f
C185 VN.n13 B 0.034358f
C186 VN.n14 B 0.034358f
C187 VN.n15 B 0.026894f
C188 VN.n16 B 0.018343f
C189 VN.n17 B 0.018343f
C190 VN.n18 B 0.018343f
C191 VN.n19 B 0.034358f
C192 VN.n20 B 0.034358f
C193 VN.n21 B 0.019939f
C194 VN.n22 B 0.018343f
C195 VN.n23 B 0.018343f
C196 VN.n24 B 0.031813f
C197 VN.n25 B 0.034358f
C198 VN.n26 B 0.033834f
C199 VN.n27 B 0.018343f
C200 VN.n28 B 0.018343f
C201 VN.n29 B 0.018343f
C202 VN.n30 B 0.036948f
C203 VN.n31 B 0.034358f
C204 VN.n32 B 0.025028f
C205 VN.n33 B 0.02961f
C206 VN.n34 B 0.047119f
C207 VN.t1 B 2.42801f
C208 VN.n35 B 0.914192f
C209 VN.n36 B 0.018343f
C210 VN.n37 B 0.017363f
C211 VN.n38 B 0.018343f
C212 VN.t2 B 2.42801f
C213 VN.n39 B 0.845262f
C214 VN.n40 B 0.018343f
C215 VN.n41 B 0.026894f
C216 VN.n42 B 0.018343f
C217 VN.n43 B 0.019939f
C218 VN.t4 B 2.65586f
C219 VN.t6 B 2.42801f
C220 VN.n44 B 0.902008f
C221 VN.n45 B 0.866573f
C222 VN.n46 B 0.21722f
C223 VN.n47 B 0.018343f
C224 VN.n48 B 0.034358f
C225 VN.n49 B 0.034358f
C226 VN.n50 B 0.026894f
C227 VN.n51 B 0.018343f
C228 VN.n52 B 0.018343f
C229 VN.n53 B 0.018343f
C230 VN.n54 B 0.034358f
C231 VN.n55 B 0.034358f
C232 VN.n56 B 0.019939f
C233 VN.n57 B 0.018343f
C234 VN.n58 B 0.018343f
C235 VN.n59 B 0.031813f
C236 VN.n60 B 0.034358f
C237 VN.n61 B 0.033834f
C238 VN.n62 B 0.018343f
C239 VN.n63 B 0.018343f
C240 VN.n64 B 0.018343f
C241 VN.n65 B 0.036948f
C242 VN.n66 B 0.034358f
C243 VN.n67 B 0.025028f
C244 VN.n68 B 0.02961f
C245 VN.n69 B 1.24048f
.ends

