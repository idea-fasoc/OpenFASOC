* NGSPICE file created from diff_pair_sample_0425.ext - technology: sky130A

.subckt diff_pair_sample_0425 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=1.41075 ps=8.88 w=8.55 l=1.66
X1 VDD2.t3 VN.t0 VTAIL.t3 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=1.41075 pd=8.88 as=3.3345 ps=17.88 w=8.55 l=1.66
X2 VDD1.t3 VP.t1 VTAIL.t6 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=1.41075 pd=8.88 as=3.3345 ps=17.88 w=8.55 l=1.66
X3 B.t11 B.t9 B.t10 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=0 ps=0 w=8.55 l=1.66
X4 VDD2.t2 VN.t1 VTAIL.t2 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=1.41075 pd=8.88 as=3.3345 ps=17.88 w=8.55 l=1.66
X5 VDD1.t1 VP.t2 VTAIL.t5 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=1.41075 pd=8.88 as=3.3345 ps=17.88 w=8.55 l=1.66
X6 VTAIL.t4 VP.t3 VDD1.t2 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=1.41075 ps=8.88 w=8.55 l=1.66
X7 B.t8 B.t6 B.t7 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=0 ps=0 w=8.55 l=1.66
X8 B.t5 B.t3 B.t4 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=0 ps=0 w=8.55 l=1.66
X9 VTAIL.t1 VN.t2 VDD2.t1 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=1.41075 ps=8.88 w=8.55 l=1.66
X10 B.t2 B.t0 B.t1 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=0 ps=0 w=8.55 l=1.66
X11 VTAIL.t0 VN.t3 VDD2.t0 w_n2164_n2678# sky130_fd_pr__pfet_01v8 ad=3.3345 pd=17.88 as=1.41075 ps=8.88 w=8.55 l=1.66
R0 VP.n8 VP.n0 161.3
R1 VP.n7 VP.n6 161.3
R2 VP.n5 VP.n1 161.3
R3 VP.n2 VP.t0 158.649
R4 VP.n2 VP.t2 158.232
R5 VP.n3 VP.t3 124.13
R6 VP.n9 VP.t1 124.13
R7 VP.n4 VP.n3 86.5341
R8 VP.n10 VP.n9 86.5341
R9 VP.n4 VP.n2 50.4155
R10 VP.n7 VP.n1 40.4934
R11 VP.n8 VP.n7 40.4934
R12 VP.n3 VP.n1 24.2228
R13 VP.n9 VP.n8 24.2228
R14 VP.n5 VP.n4 0.278367
R15 VP.n10 VP.n0 0.278367
R16 VP.n6 VP.n5 0.189894
R17 VP.n6 VP.n0 0.189894
R18 VP VP.n10 0.153454
R19 VDD1 VDD1.n1 117.642
R20 VDD1 VDD1.n0 80.9441
R21 VDD1.n0 VDD1.t0 3.80225
R22 VDD1.n0 VDD1.t1 3.80225
R23 VDD1.n1 VDD1.t2 3.80225
R24 VDD1.n1 VDD1.t3 3.80225
R25 VTAIL.n362 VTAIL.n322 756.745
R26 VTAIL.n40 VTAIL.n0 756.745
R27 VTAIL.n86 VTAIL.n46 756.745
R28 VTAIL.n132 VTAIL.n92 756.745
R29 VTAIL.n316 VTAIL.n276 756.745
R30 VTAIL.n270 VTAIL.n230 756.745
R31 VTAIL.n224 VTAIL.n184 756.745
R32 VTAIL.n178 VTAIL.n138 756.745
R33 VTAIL.n337 VTAIL.n336 585
R34 VTAIL.n334 VTAIL.n333 585
R35 VTAIL.n343 VTAIL.n342 585
R36 VTAIL.n345 VTAIL.n344 585
R37 VTAIL.n330 VTAIL.n329 585
R38 VTAIL.n351 VTAIL.n350 585
R39 VTAIL.n354 VTAIL.n353 585
R40 VTAIL.n352 VTAIL.n326 585
R41 VTAIL.n359 VTAIL.n325 585
R42 VTAIL.n361 VTAIL.n360 585
R43 VTAIL.n363 VTAIL.n362 585
R44 VTAIL.n15 VTAIL.n14 585
R45 VTAIL.n12 VTAIL.n11 585
R46 VTAIL.n21 VTAIL.n20 585
R47 VTAIL.n23 VTAIL.n22 585
R48 VTAIL.n8 VTAIL.n7 585
R49 VTAIL.n29 VTAIL.n28 585
R50 VTAIL.n32 VTAIL.n31 585
R51 VTAIL.n30 VTAIL.n4 585
R52 VTAIL.n37 VTAIL.n3 585
R53 VTAIL.n39 VTAIL.n38 585
R54 VTAIL.n41 VTAIL.n40 585
R55 VTAIL.n61 VTAIL.n60 585
R56 VTAIL.n58 VTAIL.n57 585
R57 VTAIL.n67 VTAIL.n66 585
R58 VTAIL.n69 VTAIL.n68 585
R59 VTAIL.n54 VTAIL.n53 585
R60 VTAIL.n75 VTAIL.n74 585
R61 VTAIL.n78 VTAIL.n77 585
R62 VTAIL.n76 VTAIL.n50 585
R63 VTAIL.n83 VTAIL.n49 585
R64 VTAIL.n85 VTAIL.n84 585
R65 VTAIL.n87 VTAIL.n86 585
R66 VTAIL.n107 VTAIL.n106 585
R67 VTAIL.n104 VTAIL.n103 585
R68 VTAIL.n113 VTAIL.n112 585
R69 VTAIL.n115 VTAIL.n114 585
R70 VTAIL.n100 VTAIL.n99 585
R71 VTAIL.n121 VTAIL.n120 585
R72 VTAIL.n124 VTAIL.n123 585
R73 VTAIL.n122 VTAIL.n96 585
R74 VTAIL.n129 VTAIL.n95 585
R75 VTAIL.n131 VTAIL.n130 585
R76 VTAIL.n133 VTAIL.n132 585
R77 VTAIL.n317 VTAIL.n316 585
R78 VTAIL.n315 VTAIL.n314 585
R79 VTAIL.n313 VTAIL.n279 585
R80 VTAIL.n283 VTAIL.n280 585
R81 VTAIL.n308 VTAIL.n307 585
R82 VTAIL.n306 VTAIL.n305 585
R83 VTAIL.n285 VTAIL.n284 585
R84 VTAIL.n300 VTAIL.n299 585
R85 VTAIL.n298 VTAIL.n297 585
R86 VTAIL.n289 VTAIL.n288 585
R87 VTAIL.n292 VTAIL.n291 585
R88 VTAIL.n271 VTAIL.n270 585
R89 VTAIL.n269 VTAIL.n268 585
R90 VTAIL.n267 VTAIL.n233 585
R91 VTAIL.n237 VTAIL.n234 585
R92 VTAIL.n262 VTAIL.n261 585
R93 VTAIL.n260 VTAIL.n259 585
R94 VTAIL.n239 VTAIL.n238 585
R95 VTAIL.n254 VTAIL.n253 585
R96 VTAIL.n252 VTAIL.n251 585
R97 VTAIL.n243 VTAIL.n242 585
R98 VTAIL.n246 VTAIL.n245 585
R99 VTAIL.n225 VTAIL.n224 585
R100 VTAIL.n223 VTAIL.n222 585
R101 VTAIL.n221 VTAIL.n187 585
R102 VTAIL.n191 VTAIL.n188 585
R103 VTAIL.n216 VTAIL.n215 585
R104 VTAIL.n214 VTAIL.n213 585
R105 VTAIL.n193 VTAIL.n192 585
R106 VTAIL.n208 VTAIL.n207 585
R107 VTAIL.n206 VTAIL.n205 585
R108 VTAIL.n197 VTAIL.n196 585
R109 VTAIL.n200 VTAIL.n199 585
R110 VTAIL.n179 VTAIL.n178 585
R111 VTAIL.n177 VTAIL.n176 585
R112 VTAIL.n175 VTAIL.n141 585
R113 VTAIL.n145 VTAIL.n142 585
R114 VTAIL.n170 VTAIL.n169 585
R115 VTAIL.n168 VTAIL.n167 585
R116 VTAIL.n147 VTAIL.n146 585
R117 VTAIL.n162 VTAIL.n161 585
R118 VTAIL.n160 VTAIL.n159 585
R119 VTAIL.n151 VTAIL.n150 585
R120 VTAIL.n154 VTAIL.n153 585
R121 VTAIL.t5 VTAIL.n290 329.039
R122 VTAIL.t7 VTAIL.n244 329.039
R123 VTAIL.t2 VTAIL.n198 329.039
R124 VTAIL.t1 VTAIL.n152 329.039
R125 VTAIL.t3 VTAIL.n335 329.038
R126 VTAIL.t0 VTAIL.n13 329.038
R127 VTAIL.t6 VTAIL.n59 329.038
R128 VTAIL.t4 VTAIL.n105 329.038
R129 VTAIL.n336 VTAIL.n333 171.744
R130 VTAIL.n343 VTAIL.n333 171.744
R131 VTAIL.n344 VTAIL.n343 171.744
R132 VTAIL.n344 VTAIL.n329 171.744
R133 VTAIL.n351 VTAIL.n329 171.744
R134 VTAIL.n353 VTAIL.n351 171.744
R135 VTAIL.n353 VTAIL.n352 171.744
R136 VTAIL.n352 VTAIL.n325 171.744
R137 VTAIL.n361 VTAIL.n325 171.744
R138 VTAIL.n362 VTAIL.n361 171.744
R139 VTAIL.n14 VTAIL.n11 171.744
R140 VTAIL.n21 VTAIL.n11 171.744
R141 VTAIL.n22 VTAIL.n21 171.744
R142 VTAIL.n22 VTAIL.n7 171.744
R143 VTAIL.n29 VTAIL.n7 171.744
R144 VTAIL.n31 VTAIL.n29 171.744
R145 VTAIL.n31 VTAIL.n30 171.744
R146 VTAIL.n30 VTAIL.n3 171.744
R147 VTAIL.n39 VTAIL.n3 171.744
R148 VTAIL.n40 VTAIL.n39 171.744
R149 VTAIL.n60 VTAIL.n57 171.744
R150 VTAIL.n67 VTAIL.n57 171.744
R151 VTAIL.n68 VTAIL.n67 171.744
R152 VTAIL.n68 VTAIL.n53 171.744
R153 VTAIL.n75 VTAIL.n53 171.744
R154 VTAIL.n77 VTAIL.n75 171.744
R155 VTAIL.n77 VTAIL.n76 171.744
R156 VTAIL.n76 VTAIL.n49 171.744
R157 VTAIL.n85 VTAIL.n49 171.744
R158 VTAIL.n86 VTAIL.n85 171.744
R159 VTAIL.n106 VTAIL.n103 171.744
R160 VTAIL.n113 VTAIL.n103 171.744
R161 VTAIL.n114 VTAIL.n113 171.744
R162 VTAIL.n114 VTAIL.n99 171.744
R163 VTAIL.n121 VTAIL.n99 171.744
R164 VTAIL.n123 VTAIL.n121 171.744
R165 VTAIL.n123 VTAIL.n122 171.744
R166 VTAIL.n122 VTAIL.n95 171.744
R167 VTAIL.n131 VTAIL.n95 171.744
R168 VTAIL.n132 VTAIL.n131 171.744
R169 VTAIL.n316 VTAIL.n315 171.744
R170 VTAIL.n315 VTAIL.n279 171.744
R171 VTAIL.n283 VTAIL.n279 171.744
R172 VTAIL.n307 VTAIL.n283 171.744
R173 VTAIL.n307 VTAIL.n306 171.744
R174 VTAIL.n306 VTAIL.n284 171.744
R175 VTAIL.n299 VTAIL.n284 171.744
R176 VTAIL.n299 VTAIL.n298 171.744
R177 VTAIL.n298 VTAIL.n288 171.744
R178 VTAIL.n291 VTAIL.n288 171.744
R179 VTAIL.n270 VTAIL.n269 171.744
R180 VTAIL.n269 VTAIL.n233 171.744
R181 VTAIL.n237 VTAIL.n233 171.744
R182 VTAIL.n261 VTAIL.n237 171.744
R183 VTAIL.n261 VTAIL.n260 171.744
R184 VTAIL.n260 VTAIL.n238 171.744
R185 VTAIL.n253 VTAIL.n238 171.744
R186 VTAIL.n253 VTAIL.n252 171.744
R187 VTAIL.n252 VTAIL.n242 171.744
R188 VTAIL.n245 VTAIL.n242 171.744
R189 VTAIL.n224 VTAIL.n223 171.744
R190 VTAIL.n223 VTAIL.n187 171.744
R191 VTAIL.n191 VTAIL.n187 171.744
R192 VTAIL.n215 VTAIL.n191 171.744
R193 VTAIL.n215 VTAIL.n214 171.744
R194 VTAIL.n214 VTAIL.n192 171.744
R195 VTAIL.n207 VTAIL.n192 171.744
R196 VTAIL.n207 VTAIL.n206 171.744
R197 VTAIL.n206 VTAIL.n196 171.744
R198 VTAIL.n199 VTAIL.n196 171.744
R199 VTAIL.n178 VTAIL.n177 171.744
R200 VTAIL.n177 VTAIL.n141 171.744
R201 VTAIL.n145 VTAIL.n141 171.744
R202 VTAIL.n169 VTAIL.n145 171.744
R203 VTAIL.n169 VTAIL.n168 171.744
R204 VTAIL.n168 VTAIL.n146 171.744
R205 VTAIL.n161 VTAIL.n146 171.744
R206 VTAIL.n161 VTAIL.n160 171.744
R207 VTAIL.n160 VTAIL.n150 171.744
R208 VTAIL.n153 VTAIL.n150 171.744
R209 VTAIL.n336 VTAIL.t3 85.8723
R210 VTAIL.n14 VTAIL.t0 85.8723
R211 VTAIL.n60 VTAIL.t6 85.8723
R212 VTAIL.n106 VTAIL.t4 85.8723
R213 VTAIL.n291 VTAIL.t5 85.8723
R214 VTAIL.n245 VTAIL.t7 85.8723
R215 VTAIL.n199 VTAIL.t2 85.8723
R216 VTAIL.n153 VTAIL.t1 85.8723
R217 VTAIL.n367 VTAIL.n366 32.7672
R218 VTAIL.n45 VTAIL.n44 32.7672
R219 VTAIL.n91 VTAIL.n90 32.7672
R220 VTAIL.n137 VTAIL.n136 32.7672
R221 VTAIL.n321 VTAIL.n320 32.7672
R222 VTAIL.n275 VTAIL.n274 32.7672
R223 VTAIL.n229 VTAIL.n228 32.7672
R224 VTAIL.n183 VTAIL.n182 32.7672
R225 VTAIL.n367 VTAIL.n321 21.4531
R226 VTAIL.n183 VTAIL.n137 21.4531
R227 VTAIL.n360 VTAIL.n359 13.1884
R228 VTAIL.n38 VTAIL.n37 13.1884
R229 VTAIL.n84 VTAIL.n83 13.1884
R230 VTAIL.n130 VTAIL.n129 13.1884
R231 VTAIL.n314 VTAIL.n313 13.1884
R232 VTAIL.n268 VTAIL.n267 13.1884
R233 VTAIL.n222 VTAIL.n221 13.1884
R234 VTAIL.n176 VTAIL.n175 13.1884
R235 VTAIL.n358 VTAIL.n326 12.8005
R236 VTAIL.n363 VTAIL.n324 12.8005
R237 VTAIL.n36 VTAIL.n4 12.8005
R238 VTAIL.n41 VTAIL.n2 12.8005
R239 VTAIL.n82 VTAIL.n50 12.8005
R240 VTAIL.n87 VTAIL.n48 12.8005
R241 VTAIL.n128 VTAIL.n96 12.8005
R242 VTAIL.n133 VTAIL.n94 12.8005
R243 VTAIL.n317 VTAIL.n278 12.8005
R244 VTAIL.n312 VTAIL.n280 12.8005
R245 VTAIL.n271 VTAIL.n232 12.8005
R246 VTAIL.n266 VTAIL.n234 12.8005
R247 VTAIL.n225 VTAIL.n186 12.8005
R248 VTAIL.n220 VTAIL.n188 12.8005
R249 VTAIL.n179 VTAIL.n140 12.8005
R250 VTAIL.n174 VTAIL.n142 12.8005
R251 VTAIL.n355 VTAIL.n354 12.0247
R252 VTAIL.n364 VTAIL.n322 12.0247
R253 VTAIL.n33 VTAIL.n32 12.0247
R254 VTAIL.n42 VTAIL.n0 12.0247
R255 VTAIL.n79 VTAIL.n78 12.0247
R256 VTAIL.n88 VTAIL.n46 12.0247
R257 VTAIL.n125 VTAIL.n124 12.0247
R258 VTAIL.n134 VTAIL.n92 12.0247
R259 VTAIL.n318 VTAIL.n276 12.0247
R260 VTAIL.n309 VTAIL.n308 12.0247
R261 VTAIL.n272 VTAIL.n230 12.0247
R262 VTAIL.n263 VTAIL.n262 12.0247
R263 VTAIL.n226 VTAIL.n184 12.0247
R264 VTAIL.n217 VTAIL.n216 12.0247
R265 VTAIL.n180 VTAIL.n138 12.0247
R266 VTAIL.n171 VTAIL.n170 12.0247
R267 VTAIL.n350 VTAIL.n328 11.249
R268 VTAIL.n28 VTAIL.n6 11.249
R269 VTAIL.n74 VTAIL.n52 11.249
R270 VTAIL.n120 VTAIL.n98 11.249
R271 VTAIL.n305 VTAIL.n282 11.249
R272 VTAIL.n259 VTAIL.n236 11.249
R273 VTAIL.n213 VTAIL.n190 11.249
R274 VTAIL.n167 VTAIL.n144 11.249
R275 VTAIL.n337 VTAIL.n335 10.7239
R276 VTAIL.n15 VTAIL.n13 10.7239
R277 VTAIL.n61 VTAIL.n59 10.7239
R278 VTAIL.n107 VTAIL.n105 10.7239
R279 VTAIL.n292 VTAIL.n290 10.7239
R280 VTAIL.n246 VTAIL.n244 10.7239
R281 VTAIL.n200 VTAIL.n198 10.7239
R282 VTAIL.n154 VTAIL.n152 10.7239
R283 VTAIL.n349 VTAIL.n330 10.4732
R284 VTAIL.n27 VTAIL.n8 10.4732
R285 VTAIL.n73 VTAIL.n54 10.4732
R286 VTAIL.n119 VTAIL.n100 10.4732
R287 VTAIL.n304 VTAIL.n285 10.4732
R288 VTAIL.n258 VTAIL.n239 10.4732
R289 VTAIL.n212 VTAIL.n193 10.4732
R290 VTAIL.n166 VTAIL.n147 10.4732
R291 VTAIL.n346 VTAIL.n345 9.69747
R292 VTAIL.n24 VTAIL.n23 9.69747
R293 VTAIL.n70 VTAIL.n69 9.69747
R294 VTAIL.n116 VTAIL.n115 9.69747
R295 VTAIL.n301 VTAIL.n300 9.69747
R296 VTAIL.n255 VTAIL.n254 9.69747
R297 VTAIL.n209 VTAIL.n208 9.69747
R298 VTAIL.n163 VTAIL.n162 9.69747
R299 VTAIL.n366 VTAIL.n365 9.45567
R300 VTAIL.n44 VTAIL.n43 9.45567
R301 VTAIL.n90 VTAIL.n89 9.45567
R302 VTAIL.n136 VTAIL.n135 9.45567
R303 VTAIL.n320 VTAIL.n319 9.45567
R304 VTAIL.n274 VTAIL.n273 9.45567
R305 VTAIL.n228 VTAIL.n227 9.45567
R306 VTAIL.n182 VTAIL.n181 9.45567
R307 VTAIL.n365 VTAIL.n364 9.3005
R308 VTAIL.n324 VTAIL.n323 9.3005
R309 VTAIL.n339 VTAIL.n338 9.3005
R310 VTAIL.n341 VTAIL.n340 9.3005
R311 VTAIL.n332 VTAIL.n331 9.3005
R312 VTAIL.n347 VTAIL.n346 9.3005
R313 VTAIL.n349 VTAIL.n348 9.3005
R314 VTAIL.n328 VTAIL.n327 9.3005
R315 VTAIL.n356 VTAIL.n355 9.3005
R316 VTAIL.n358 VTAIL.n357 9.3005
R317 VTAIL.n43 VTAIL.n42 9.3005
R318 VTAIL.n2 VTAIL.n1 9.3005
R319 VTAIL.n17 VTAIL.n16 9.3005
R320 VTAIL.n19 VTAIL.n18 9.3005
R321 VTAIL.n10 VTAIL.n9 9.3005
R322 VTAIL.n25 VTAIL.n24 9.3005
R323 VTAIL.n27 VTAIL.n26 9.3005
R324 VTAIL.n6 VTAIL.n5 9.3005
R325 VTAIL.n34 VTAIL.n33 9.3005
R326 VTAIL.n36 VTAIL.n35 9.3005
R327 VTAIL.n89 VTAIL.n88 9.3005
R328 VTAIL.n48 VTAIL.n47 9.3005
R329 VTAIL.n63 VTAIL.n62 9.3005
R330 VTAIL.n65 VTAIL.n64 9.3005
R331 VTAIL.n56 VTAIL.n55 9.3005
R332 VTAIL.n71 VTAIL.n70 9.3005
R333 VTAIL.n73 VTAIL.n72 9.3005
R334 VTAIL.n52 VTAIL.n51 9.3005
R335 VTAIL.n80 VTAIL.n79 9.3005
R336 VTAIL.n82 VTAIL.n81 9.3005
R337 VTAIL.n135 VTAIL.n134 9.3005
R338 VTAIL.n94 VTAIL.n93 9.3005
R339 VTAIL.n109 VTAIL.n108 9.3005
R340 VTAIL.n111 VTAIL.n110 9.3005
R341 VTAIL.n102 VTAIL.n101 9.3005
R342 VTAIL.n117 VTAIL.n116 9.3005
R343 VTAIL.n119 VTAIL.n118 9.3005
R344 VTAIL.n98 VTAIL.n97 9.3005
R345 VTAIL.n126 VTAIL.n125 9.3005
R346 VTAIL.n128 VTAIL.n127 9.3005
R347 VTAIL.n294 VTAIL.n293 9.3005
R348 VTAIL.n296 VTAIL.n295 9.3005
R349 VTAIL.n287 VTAIL.n286 9.3005
R350 VTAIL.n302 VTAIL.n301 9.3005
R351 VTAIL.n304 VTAIL.n303 9.3005
R352 VTAIL.n282 VTAIL.n281 9.3005
R353 VTAIL.n310 VTAIL.n309 9.3005
R354 VTAIL.n312 VTAIL.n311 9.3005
R355 VTAIL.n319 VTAIL.n318 9.3005
R356 VTAIL.n278 VTAIL.n277 9.3005
R357 VTAIL.n248 VTAIL.n247 9.3005
R358 VTAIL.n250 VTAIL.n249 9.3005
R359 VTAIL.n241 VTAIL.n240 9.3005
R360 VTAIL.n256 VTAIL.n255 9.3005
R361 VTAIL.n258 VTAIL.n257 9.3005
R362 VTAIL.n236 VTAIL.n235 9.3005
R363 VTAIL.n264 VTAIL.n263 9.3005
R364 VTAIL.n266 VTAIL.n265 9.3005
R365 VTAIL.n273 VTAIL.n272 9.3005
R366 VTAIL.n232 VTAIL.n231 9.3005
R367 VTAIL.n202 VTAIL.n201 9.3005
R368 VTAIL.n204 VTAIL.n203 9.3005
R369 VTAIL.n195 VTAIL.n194 9.3005
R370 VTAIL.n210 VTAIL.n209 9.3005
R371 VTAIL.n212 VTAIL.n211 9.3005
R372 VTAIL.n190 VTAIL.n189 9.3005
R373 VTAIL.n218 VTAIL.n217 9.3005
R374 VTAIL.n220 VTAIL.n219 9.3005
R375 VTAIL.n227 VTAIL.n226 9.3005
R376 VTAIL.n186 VTAIL.n185 9.3005
R377 VTAIL.n156 VTAIL.n155 9.3005
R378 VTAIL.n158 VTAIL.n157 9.3005
R379 VTAIL.n149 VTAIL.n148 9.3005
R380 VTAIL.n164 VTAIL.n163 9.3005
R381 VTAIL.n166 VTAIL.n165 9.3005
R382 VTAIL.n144 VTAIL.n143 9.3005
R383 VTAIL.n172 VTAIL.n171 9.3005
R384 VTAIL.n174 VTAIL.n173 9.3005
R385 VTAIL.n181 VTAIL.n180 9.3005
R386 VTAIL.n140 VTAIL.n139 9.3005
R387 VTAIL.n342 VTAIL.n332 8.92171
R388 VTAIL.n20 VTAIL.n10 8.92171
R389 VTAIL.n66 VTAIL.n56 8.92171
R390 VTAIL.n112 VTAIL.n102 8.92171
R391 VTAIL.n297 VTAIL.n287 8.92171
R392 VTAIL.n251 VTAIL.n241 8.92171
R393 VTAIL.n205 VTAIL.n195 8.92171
R394 VTAIL.n159 VTAIL.n149 8.92171
R395 VTAIL.n341 VTAIL.n334 8.14595
R396 VTAIL.n19 VTAIL.n12 8.14595
R397 VTAIL.n65 VTAIL.n58 8.14595
R398 VTAIL.n111 VTAIL.n104 8.14595
R399 VTAIL.n296 VTAIL.n289 8.14595
R400 VTAIL.n250 VTAIL.n243 8.14595
R401 VTAIL.n204 VTAIL.n197 8.14595
R402 VTAIL.n158 VTAIL.n151 8.14595
R403 VTAIL.n338 VTAIL.n337 7.3702
R404 VTAIL.n16 VTAIL.n15 7.3702
R405 VTAIL.n62 VTAIL.n61 7.3702
R406 VTAIL.n108 VTAIL.n107 7.3702
R407 VTAIL.n293 VTAIL.n292 7.3702
R408 VTAIL.n247 VTAIL.n246 7.3702
R409 VTAIL.n201 VTAIL.n200 7.3702
R410 VTAIL.n155 VTAIL.n154 7.3702
R411 VTAIL.n338 VTAIL.n334 5.81868
R412 VTAIL.n16 VTAIL.n12 5.81868
R413 VTAIL.n62 VTAIL.n58 5.81868
R414 VTAIL.n108 VTAIL.n104 5.81868
R415 VTAIL.n293 VTAIL.n289 5.81868
R416 VTAIL.n247 VTAIL.n243 5.81868
R417 VTAIL.n201 VTAIL.n197 5.81868
R418 VTAIL.n155 VTAIL.n151 5.81868
R419 VTAIL.n342 VTAIL.n341 5.04292
R420 VTAIL.n20 VTAIL.n19 5.04292
R421 VTAIL.n66 VTAIL.n65 5.04292
R422 VTAIL.n112 VTAIL.n111 5.04292
R423 VTAIL.n297 VTAIL.n296 5.04292
R424 VTAIL.n251 VTAIL.n250 5.04292
R425 VTAIL.n205 VTAIL.n204 5.04292
R426 VTAIL.n159 VTAIL.n158 5.04292
R427 VTAIL.n345 VTAIL.n332 4.26717
R428 VTAIL.n23 VTAIL.n10 4.26717
R429 VTAIL.n69 VTAIL.n56 4.26717
R430 VTAIL.n115 VTAIL.n102 4.26717
R431 VTAIL.n300 VTAIL.n287 4.26717
R432 VTAIL.n254 VTAIL.n241 4.26717
R433 VTAIL.n208 VTAIL.n195 4.26717
R434 VTAIL.n162 VTAIL.n149 4.26717
R435 VTAIL.n346 VTAIL.n330 3.49141
R436 VTAIL.n24 VTAIL.n8 3.49141
R437 VTAIL.n70 VTAIL.n54 3.49141
R438 VTAIL.n116 VTAIL.n100 3.49141
R439 VTAIL.n301 VTAIL.n285 3.49141
R440 VTAIL.n255 VTAIL.n239 3.49141
R441 VTAIL.n209 VTAIL.n193 3.49141
R442 VTAIL.n163 VTAIL.n147 3.49141
R443 VTAIL.n350 VTAIL.n349 2.71565
R444 VTAIL.n28 VTAIL.n27 2.71565
R445 VTAIL.n74 VTAIL.n73 2.71565
R446 VTAIL.n120 VTAIL.n119 2.71565
R447 VTAIL.n305 VTAIL.n304 2.71565
R448 VTAIL.n259 VTAIL.n258 2.71565
R449 VTAIL.n213 VTAIL.n212 2.71565
R450 VTAIL.n167 VTAIL.n166 2.71565
R451 VTAIL.n339 VTAIL.n335 2.41285
R452 VTAIL.n17 VTAIL.n13 2.41285
R453 VTAIL.n63 VTAIL.n59 2.41285
R454 VTAIL.n109 VTAIL.n105 2.41285
R455 VTAIL.n294 VTAIL.n290 2.41285
R456 VTAIL.n248 VTAIL.n244 2.41285
R457 VTAIL.n202 VTAIL.n198 2.41285
R458 VTAIL.n156 VTAIL.n152 2.41285
R459 VTAIL.n354 VTAIL.n328 1.93989
R460 VTAIL.n366 VTAIL.n322 1.93989
R461 VTAIL.n32 VTAIL.n6 1.93989
R462 VTAIL.n44 VTAIL.n0 1.93989
R463 VTAIL.n78 VTAIL.n52 1.93989
R464 VTAIL.n90 VTAIL.n46 1.93989
R465 VTAIL.n124 VTAIL.n98 1.93989
R466 VTAIL.n136 VTAIL.n92 1.93989
R467 VTAIL.n320 VTAIL.n276 1.93989
R468 VTAIL.n308 VTAIL.n282 1.93989
R469 VTAIL.n274 VTAIL.n230 1.93989
R470 VTAIL.n262 VTAIL.n236 1.93989
R471 VTAIL.n228 VTAIL.n184 1.93989
R472 VTAIL.n216 VTAIL.n190 1.93989
R473 VTAIL.n182 VTAIL.n138 1.93989
R474 VTAIL.n170 VTAIL.n144 1.93989
R475 VTAIL.n229 VTAIL.n183 1.71602
R476 VTAIL.n321 VTAIL.n275 1.71602
R477 VTAIL.n137 VTAIL.n91 1.71602
R478 VTAIL.n355 VTAIL.n326 1.16414
R479 VTAIL.n364 VTAIL.n363 1.16414
R480 VTAIL.n33 VTAIL.n4 1.16414
R481 VTAIL.n42 VTAIL.n41 1.16414
R482 VTAIL.n79 VTAIL.n50 1.16414
R483 VTAIL.n88 VTAIL.n87 1.16414
R484 VTAIL.n125 VTAIL.n96 1.16414
R485 VTAIL.n134 VTAIL.n133 1.16414
R486 VTAIL.n318 VTAIL.n317 1.16414
R487 VTAIL.n309 VTAIL.n280 1.16414
R488 VTAIL.n272 VTAIL.n271 1.16414
R489 VTAIL.n263 VTAIL.n234 1.16414
R490 VTAIL.n226 VTAIL.n225 1.16414
R491 VTAIL.n217 VTAIL.n188 1.16414
R492 VTAIL.n180 VTAIL.n179 1.16414
R493 VTAIL.n171 VTAIL.n142 1.16414
R494 VTAIL VTAIL.n45 0.916448
R495 VTAIL VTAIL.n367 0.800069
R496 VTAIL.n275 VTAIL.n229 0.470328
R497 VTAIL.n91 VTAIL.n45 0.470328
R498 VTAIL.n359 VTAIL.n358 0.388379
R499 VTAIL.n360 VTAIL.n324 0.388379
R500 VTAIL.n37 VTAIL.n36 0.388379
R501 VTAIL.n38 VTAIL.n2 0.388379
R502 VTAIL.n83 VTAIL.n82 0.388379
R503 VTAIL.n84 VTAIL.n48 0.388379
R504 VTAIL.n129 VTAIL.n128 0.388379
R505 VTAIL.n130 VTAIL.n94 0.388379
R506 VTAIL.n314 VTAIL.n278 0.388379
R507 VTAIL.n313 VTAIL.n312 0.388379
R508 VTAIL.n268 VTAIL.n232 0.388379
R509 VTAIL.n267 VTAIL.n266 0.388379
R510 VTAIL.n222 VTAIL.n186 0.388379
R511 VTAIL.n221 VTAIL.n220 0.388379
R512 VTAIL.n176 VTAIL.n140 0.388379
R513 VTAIL.n175 VTAIL.n174 0.388379
R514 VTAIL.n340 VTAIL.n339 0.155672
R515 VTAIL.n340 VTAIL.n331 0.155672
R516 VTAIL.n347 VTAIL.n331 0.155672
R517 VTAIL.n348 VTAIL.n347 0.155672
R518 VTAIL.n348 VTAIL.n327 0.155672
R519 VTAIL.n356 VTAIL.n327 0.155672
R520 VTAIL.n357 VTAIL.n356 0.155672
R521 VTAIL.n357 VTAIL.n323 0.155672
R522 VTAIL.n365 VTAIL.n323 0.155672
R523 VTAIL.n18 VTAIL.n17 0.155672
R524 VTAIL.n18 VTAIL.n9 0.155672
R525 VTAIL.n25 VTAIL.n9 0.155672
R526 VTAIL.n26 VTAIL.n25 0.155672
R527 VTAIL.n26 VTAIL.n5 0.155672
R528 VTAIL.n34 VTAIL.n5 0.155672
R529 VTAIL.n35 VTAIL.n34 0.155672
R530 VTAIL.n35 VTAIL.n1 0.155672
R531 VTAIL.n43 VTAIL.n1 0.155672
R532 VTAIL.n64 VTAIL.n63 0.155672
R533 VTAIL.n64 VTAIL.n55 0.155672
R534 VTAIL.n71 VTAIL.n55 0.155672
R535 VTAIL.n72 VTAIL.n71 0.155672
R536 VTAIL.n72 VTAIL.n51 0.155672
R537 VTAIL.n80 VTAIL.n51 0.155672
R538 VTAIL.n81 VTAIL.n80 0.155672
R539 VTAIL.n81 VTAIL.n47 0.155672
R540 VTAIL.n89 VTAIL.n47 0.155672
R541 VTAIL.n110 VTAIL.n109 0.155672
R542 VTAIL.n110 VTAIL.n101 0.155672
R543 VTAIL.n117 VTAIL.n101 0.155672
R544 VTAIL.n118 VTAIL.n117 0.155672
R545 VTAIL.n118 VTAIL.n97 0.155672
R546 VTAIL.n126 VTAIL.n97 0.155672
R547 VTAIL.n127 VTAIL.n126 0.155672
R548 VTAIL.n127 VTAIL.n93 0.155672
R549 VTAIL.n135 VTAIL.n93 0.155672
R550 VTAIL.n319 VTAIL.n277 0.155672
R551 VTAIL.n311 VTAIL.n277 0.155672
R552 VTAIL.n311 VTAIL.n310 0.155672
R553 VTAIL.n310 VTAIL.n281 0.155672
R554 VTAIL.n303 VTAIL.n281 0.155672
R555 VTAIL.n303 VTAIL.n302 0.155672
R556 VTAIL.n302 VTAIL.n286 0.155672
R557 VTAIL.n295 VTAIL.n286 0.155672
R558 VTAIL.n295 VTAIL.n294 0.155672
R559 VTAIL.n273 VTAIL.n231 0.155672
R560 VTAIL.n265 VTAIL.n231 0.155672
R561 VTAIL.n265 VTAIL.n264 0.155672
R562 VTAIL.n264 VTAIL.n235 0.155672
R563 VTAIL.n257 VTAIL.n235 0.155672
R564 VTAIL.n257 VTAIL.n256 0.155672
R565 VTAIL.n256 VTAIL.n240 0.155672
R566 VTAIL.n249 VTAIL.n240 0.155672
R567 VTAIL.n249 VTAIL.n248 0.155672
R568 VTAIL.n227 VTAIL.n185 0.155672
R569 VTAIL.n219 VTAIL.n185 0.155672
R570 VTAIL.n219 VTAIL.n218 0.155672
R571 VTAIL.n218 VTAIL.n189 0.155672
R572 VTAIL.n211 VTAIL.n189 0.155672
R573 VTAIL.n211 VTAIL.n210 0.155672
R574 VTAIL.n210 VTAIL.n194 0.155672
R575 VTAIL.n203 VTAIL.n194 0.155672
R576 VTAIL.n203 VTAIL.n202 0.155672
R577 VTAIL.n181 VTAIL.n139 0.155672
R578 VTAIL.n173 VTAIL.n139 0.155672
R579 VTAIL.n173 VTAIL.n172 0.155672
R580 VTAIL.n172 VTAIL.n143 0.155672
R581 VTAIL.n165 VTAIL.n143 0.155672
R582 VTAIL.n165 VTAIL.n164 0.155672
R583 VTAIL.n164 VTAIL.n148 0.155672
R584 VTAIL.n157 VTAIL.n148 0.155672
R585 VTAIL.n157 VTAIL.n156 0.155672
R586 VN.n0 VN.t3 158.649
R587 VN.n1 VN.t1 158.649
R588 VN.n0 VN.t0 158.232
R589 VN.n1 VN.t2 158.232
R590 VN VN.n1 50.6944
R591 VN VN.n0 9.69059
R592 VDD2.n2 VDD2.n0 117.118
R593 VDD2.n2 VDD2.n1 80.8859
R594 VDD2.n1 VDD2.t1 3.80225
R595 VDD2.n1 VDD2.t2 3.80225
R596 VDD2.n0 VDD2.t0 3.80225
R597 VDD2.n0 VDD2.t3 3.80225
R598 VDD2 VDD2.n2 0.0586897
R599 B.n281 B.n82 585
R600 B.n280 B.n279 585
R601 B.n278 B.n83 585
R602 B.n277 B.n276 585
R603 B.n275 B.n84 585
R604 B.n274 B.n273 585
R605 B.n272 B.n85 585
R606 B.n271 B.n270 585
R607 B.n269 B.n86 585
R608 B.n268 B.n267 585
R609 B.n266 B.n87 585
R610 B.n265 B.n264 585
R611 B.n263 B.n88 585
R612 B.n262 B.n261 585
R613 B.n260 B.n89 585
R614 B.n259 B.n258 585
R615 B.n257 B.n90 585
R616 B.n256 B.n255 585
R617 B.n254 B.n91 585
R618 B.n253 B.n252 585
R619 B.n251 B.n92 585
R620 B.n250 B.n249 585
R621 B.n248 B.n93 585
R622 B.n247 B.n246 585
R623 B.n245 B.n94 585
R624 B.n244 B.n243 585
R625 B.n242 B.n95 585
R626 B.n241 B.n240 585
R627 B.n239 B.n96 585
R628 B.n238 B.n237 585
R629 B.n236 B.n97 585
R630 B.n235 B.n234 585
R631 B.n232 B.n98 585
R632 B.n231 B.n230 585
R633 B.n229 B.n101 585
R634 B.n228 B.n227 585
R635 B.n226 B.n102 585
R636 B.n225 B.n224 585
R637 B.n223 B.n103 585
R638 B.n222 B.n221 585
R639 B.n220 B.n104 585
R640 B.n218 B.n217 585
R641 B.n216 B.n107 585
R642 B.n215 B.n214 585
R643 B.n213 B.n108 585
R644 B.n212 B.n211 585
R645 B.n210 B.n109 585
R646 B.n209 B.n208 585
R647 B.n207 B.n110 585
R648 B.n206 B.n205 585
R649 B.n204 B.n111 585
R650 B.n203 B.n202 585
R651 B.n201 B.n112 585
R652 B.n200 B.n199 585
R653 B.n198 B.n113 585
R654 B.n197 B.n196 585
R655 B.n195 B.n114 585
R656 B.n194 B.n193 585
R657 B.n192 B.n115 585
R658 B.n191 B.n190 585
R659 B.n189 B.n116 585
R660 B.n188 B.n187 585
R661 B.n186 B.n117 585
R662 B.n185 B.n184 585
R663 B.n183 B.n118 585
R664 B.n182 B.n181 585
R665 B.n180 B.n119 585
R666 B.n179 B.n178 585
R667 B.n177 B.n120 585
R668 B.n176 B.n175 585
R669 B.n174 B.n121 585
R670 B.n173 B.n172 585
R671 B.n171 B.n122 585
R672 B.n283 B.n282 585
R673 B.n284 B.n81 585
R674 B.n286 B.n285 585
R675 B.n287 B.n80 585
R676 B.n289 B.n288 585
R677 B.n290 B.n79 585
R678 B.n292 B.n291 585
R679 B.n293 B.n78 585
R680 B.n295 B.n294 585
R681 B.n296 B.n77 585
R682 B.n298 B.n297 585
R683 B.n299 B.n76 585
R684 B.n301 B.n300 585
R685 B.n302 B.n75 585
R686 B.n304 B.n303 585
R687 B.n305 B.n74 585
R688 B.n307 B.n306 585
R689 B.n308 B.n73 585
R690 B.n310 B.n309 585
R691 B.n311 B.n72 585
R692 B.n313 B.n312 585
R693 B.n314 B.n71 585
R694 B.n316 B.n315 585
R695 B.n317 B.n70 585
R696 B.n319 B.n318 585
R697 B.n320 B.n69 585
R698 B.n322 B.n321 585
R699 B.n323 B.n68 585
R700 B.n325 B.n324 585
R701 B.n326 B.n67 585
R702 B.n328 B.n327 585
R703 B.n329 B.n66 585
R704 B.n331 B.n330 585
R705 B.n332 B.n65 585
R706 B.n334 B.n333 585
R707 B.n335 B.n64 585
R708 B.n337 B.n336 585
R709 B.n338 B.n63 585
R710 B.n340 B.n339 585
R711 B.n341 B.n62 585
R712 B.n343 B.n342 585
R713 B.n344 B.n61 585
R714 B.n346 B.n345 585
R715 B.n347 B.n60 585
R716 B.n349 B.n348 585
R717 B.n350 B.n59 585
R718 B.n352 B.n351 585
R719 B.n353 B.n58 585
R720 B.n355 B.n354 585
R721 B.n356 B.n57 585
R722 B.n358 B.n357 585
R723 B.n359 B.n56 585
R724 B.n470 B.n469 585
R725 B.n468 B.n15 585
R726 B.n467 B.n466 585
R727 B.n465 B.n16 585
R728 B.n464 B.n463 585
R729 B.n462 B.n17 585
R730 B.n461 B.n460 585
R731 B.n459 B.n18 585
R732 B.n458 B.n457 585
R733 B.n456 B.n19 585
R734 B.n455 B.n454 585
R735 B.n453 B.n20 585
R736 B.n452 B.n451 585
R737 B.n450 B.n21 585
R738 B.n449 B.n448 585
R739 B.n447 B.n22 585
R740 B.n446 B.n445 585
R741 B.n444 B.n23 585
R742 B.n443 B.n442 585
R743 B.n441 B.n24 585
R744 B.n440 B.n439 585
R745 B.n438 B.n25 585
R746 B.n437 B.n436 585
R747 B.n435 B.n26 585
R748 B.n434 B.n433 585
R749 B.n432 B.n27 585
R750 B.n431 B.n430 585
R751 B.n429 B.n28 585
R752 B.n428 B.n427 585
R753 B.n426 B.n29 585
R754 B.n425 B.n424 585
R755 B.n423 B.n30 585
R756 B.n422 B.n421 585
R757 B.n420 B.n31 585
R758 B.n419 B.n418 585
R759 B.n417 B.n35 585
R760 B.n416 B.n415 585
R761 B.n414 B.n36 585
R762 B.n413 B.n412 585
R763 B.n411 B.n37 585
R764 B.n410 B.n409 585
R765 B.n407 B.n38 585
R766 B.n406 B.n405 585
R767 B.n404 B.n41 585
R768 B.n403 B.n402 585
R769 B.n401 B.n42 585
R770 B.n400 B.n399 585
R771 B.n398 B.n43 585
R772 B.n397 B.n396 585
R773 B.n395 B.n44 585
R774 B.n394 B.n393 585
R775 B.n392 B.n45 585
R776 B.n391 B.n390 585
R777 B.n389 B.n46 585
R778 B.n388 B.n387 585
R779 B.n386 B.n47 585
R780 B.n385 B.n384 585
R781 B.n383 B.n48 585
R782 B.n382 B.n381 585
R783 B.n380 B.n49 585
R784 B.n379 B.n378 585
R785 B.n377 B.n50 585
R786 B.n376 B.n375 585
R787 B.n374 B.n51 585
R788 B.n373 B.n372 585
R789 B.n371 B.n52 585
R790 B.n370 B.n369 585
R791 B.n368 B.n53 585
R792 B.n367 B.n366 585
R793 B.n365 B.n54 585
R794 B.n364 B.n363 585
R795 B.n362 B.n55 585
R796 B.n361 B.n360 585
R797 B.n471 B.n14 585
R798 B.n473 B.n472 585
R799 B.n474 B.n13 585
R800 B.n476 B.n475 585
R801 B.n477 B.n12 585
R802 B.n479 B.n478 585
R803 B.n480 B.n11 585
R804 B.n482 B.n481 585
R805 B.n483 B.n10 585
R806 B.n485 B.n484 585
R807 B.n486 B.n9 585
R808 B.n488 B.n487 585
R809 B.n489 B.n8 585
R810 B.n491 B.n490 585
R811 B.n492 B.n7 585
R812 B.n494 B.n493 585
R813 B.n495 B.n6 585
R814 B.n497 B.n496 585
R815 B.n498 B.n5 585
R816 B.n500 B.n499 585
R817 B.n501 B.n4 585
R818 B.n503 B.n502 585
R819 B.n504 B.n3 585
R820 B.n506 B.n505 585
R821 B.n507 B.n0 585
R822 B.n2 B.n1 585
R823 B.n135 B.n134 585
R824 B.n137 B.n136 585
R825 B.n138 B.n133 585
R826 B.n140 B.n139 585
R827 B.n141 B.n132 585
R828 B.n143 B.n142 585
R829 B.n144 B.n131 585
R830 B.n146 B.n145 585
R831 B.n147 B.n130 585
R832 B.n149 B.n148 585
R833 B.n150 B.n129 585
R834 B.n152 B.n151 585
R835 B.n153 B.n128 585
R836 B.n155 B.n154 585
R837 B.n156 B.n127 585
R838 B.n158 B.n157 585
R839 B.n159 B.n126 585
R840 B.n161 B.n160 585
R841 B.n162 B.n125 585
R842 B.n164 B.n163 585
R843 B.n165 B.n124 585
R844 B.n167 B.n166 585
R845 B.n168 B.n123 585
R846 B.n170 B.n169 585
R847 B.n169 B.n122 487.695
R848 B.n283 B.n82 487.695
R849 B.n361 B.n56 487.695
R850 B.n471 B.n470 487.695
R851 B.n99 B.t7 351.967
R852 B.n39 B.t5 351.967
R853 B.n105 B.t10 351.967
R854 B.n32 B.t2 351.967
R855 B.n105 B.t9 330.12
R856 B.n99 B.t6 330.12
R857 B.n39 B.t3 330.12
R858 B.n32 B.t0 330.12
R859 B.n100 B.t8 313.373
R860 B.n40 B.t4 313.373
R861 B.n106 B.t11 313.373
R862 B.n33 B.t1 313.373
R863 B.n509 B.n508 256.663
R864 B.n508 B.n507 235.042
R865 B.n508 B.n2 235.042
R866 B.n173 B.n122 163.367
R867 B.n174 B.n173 163.367
R868 B.n175 B.n174 163.367
R869 B.n175 B.n120 163.367
R870 B.n179 B.n120 163.367
R871 B.n180 B.n179 163.367
R872 B.n181 B.n180 163.367
R873 B.n181 B.n118 163.367
R874 B.n185 B.n118 163.367
R875 B.n186 B.n185 163.367
R876 B.n187 B.n186 163.367
R877 B.n187 B.n116 163.367
R878 B.n191 B.n116 163.367
R879 B.n192 B.n191 163.367
R880 B.n193 B.n192 163.367
R881 B.n193 B.n114 163.367
R882 B.n197 B.n114 163.367
R883 B.n198 B.n197 163.367
R884 B.n199 B.n198 163.367
R885 B.n199 B.n112 163.367
R886 B.n203 B.n112 163.367
R887 B.n204 B.n203 163.367
R888 B.n205 B.n204 163.367
R889 B.n205 B.n110 163.367
R890 B.n209 B.n110 163.367
R891 B.n210 B.n209 163.367
R892 B.n211 B.n210 163.367
R893 B.n211 B.n108 163.367
R894 B.n215 B.n108 163.367
R895 B.n216 B.n215 163.367
R896 B.n217 B.n216 163.367
R897 B.n217 B.n104 163.367
R898 B.n222 B.n104 163.367
R899 B.n223 B.n222 163.367
R900 B.n224 B.n223 163.367
R901 B.n224 B.n102 163.367
R902 B.n228 B.n102 163.367
R903 B.n229 B.n228 163.367
R904 B.n230 B.n229 163.367
R905 B.n230 B.n98 163.367
R906 B.n235 B.n98 163.367
R907 B.n236 B.n235 163.367
R908 B.n237 B.n236 163.367
R909 B.n237 B.n96 163.367
R910 B.n241 B.n96 163.367
R911 B.n242 B.n241 163.367
R912 B.n243 B.n242 163.367
R913 B.n243 B.n94 163.367
R914 B.n247 B.n94 163.367
R915 B.n248 B.n247 163.367
R916 B.n249 B.n248 163.367
R917 B.n249 B.n92 163.367
R918 B.n253 B.n92 163.367
R919 B.n254 B.n253 163.367
R920 B.n255 B.n254 163.367
R921 B.n255 B.n90 163.367
R922 B.n259 B.n90 163.367
R923 B.n260 B.n259 163.367
R924 B.n261 B.n260 163.367
R925 B.n261 B.n88 163.367
R926 B.n265 B.n88 163.367
R927 B.n266 B.n265 163.367
R928 B.n267 B.n266 163.367
R929 B.n267 B.n86 163.367
R930 B.n271 B.n86 163.367
R931 B.n272 B.n271 163.367
R932 B.n273 B.n272 163.367
R933 B.n273 B.n84 163.367
R934 B.n277 B.n84 163.367
R935 B.n278 B.n277 163.367
R936 B.n279 B.n278 163.367
R937 B.n279 B.n82 163.367
R938 B.n357 B.n56 163.367
R939 B.n357 B.n356 163.367
R940 B.n356 B.n355 163.367
R941 B.n355 B.n58 163.367
R942 B.n351 B.n58 163.367
R943 B.n351 B.n350 163.367
R944 B.n350 B.n349 163.367
R945 B.n349 B.n60 163.367
R946 B.n345 B.n60 163.367
R947 B.n345 B.n344 163.367
R948 B.n344 B.n343 163.367
R949 B.n343 B.n62 163.367
R950 B.n339 B.n62 163.367
R951 B.n339 B.n338 163.367
R952 B.n338 B.n337 163.367
R953 B.n337 B.n64 163.367
R954 B.n333 B.n64 163.367
R955 B.n333 B.n332 163.367
R956 B.n332 B.n331 163.367
R957 B.n331 B.n66 163.367
R958 B.n327 B.n66 163.367
R959 B.n327 B.n326 163.367
R960 B.n326 B.n325 163.367
R961 B.n325 B.n68 163.367
R962 B.n321 B.n68 163.367
R963 B.n321 B.n320 163.367
R964 B.n320 B.n319 163.367
R965 B.n319 B.n70 163.367
R966 B.n315 B.n70 163.367
R967 B.n315 B.n314 163.367
R968 B.n314 B.n313 163.367
R969 B.n313 B.n72 163.367
R970 B.n309 B.n72 163.367
R971 B.n309 B.n308 163.367
R972 B.n308 B.n307 163.367
R973 B.n307 B.n74 163.367
R974 B.n303 B.n74 163.367
R975 B.n303 B.n302 163.367
R976 B.n302 B.n301 163.367
R977 B.n301 B.n76 163.367
R978 B.n297 B.n76 163.367
R979 B.n297 B.n296 163.367
R980 B.n296 B.n295 163.367
R981 B.n295 B.n78 163.367
R982 B.n291 B.n78 163.367
R983 B.n291 B.n290 163.367
R984 B.n290 B.n289 163.367
R985 B.n289 B.n80 163.367
R986 B.n285 B.n80 163.367
R987 B.n285 B.n284 163.367
R988 B.n284 B.n283 163.367
R989 B.n470 B.n15 163.367
R990 B.n466 B.n15 163.367
R991 B.n466 B.n465 163.367
R992 B.n465 B.n464 163.367
R993 B.n464 B.n17 163.367
R994 B.n460 B.n17 163.367
R995 B.n460 B.n459 163.367
R996 B.n459 B.n458 163.367
R997 B.n458 B.n19 163.367
R998 B.n454 B.n19 163.367
R999 B.n454 B.n453 163.367
R1000 B.n453 B.n452 163.367
R1001 B.n452 B.n21 163.367
R1002 B.n448 B.n21 163.367
R1003 B.n448 B.n447 163.367
R1004 B.n447 B.n446 163.367
R1005 B.n446 B.n23 163.367
R1006 B.n442 B.n23 163.367
R1007 B.n442 B.n441 163.367
R1008 B.n441 B.n440 163.367
R1009 B.n440 B.n25 163.367
R1010 B.n436 B.n25 163.367
R1011 B.n436 B.n435 163.367
R1012 B.n435 B.n434 163.367
R1013 B.n434 B.n27 163.367
R1014 B.n430 B.n27 163.367
R1015 B.n430 B.n429 163.367
R1016 B.n429 B.n428 163.367
R1017 B.n428 B.n29 163.367
R1018 B.n424 B.n29 163.367
R1019 B.n424 B.n423 163.367
R1020 B.n423 B.n422 163.367
R1021 B.n422 B.n31 163.367
R1022 B.n418 B.n31 163.367
R1023 B.n418 B.n417 163.367
R1024 B.n417 B.n416 163.367
R1025 B.n416 B.n36 163.367
R1026 B.n412 B.n36 163.367
R1027 B.n412 B.n411 163.367
R1028 B.n411 B.n410 163.367
R1029 B.n410 B.n38 163.367
R1030 B.n405 B.n38 163.367
R1031 B.n405 B.n404 163.367
R1032 B.n404 B.n403 163.367
R1033 B.n403 B.n42 163.367
R1034 B.n399 B.n42 163.367
R1035 B.n399 B.n398 163.367
R1036 B.n398 B.n397 163.367
R1037 B.n397 B.n44 163.367
R1038 B.n393 B.n44 163.367
R1039 B.n393 B.n392 163.367
R1040 B.n392 B.n391 163.367
R1041 B.n391 B.n46 163.367
R1042 B.n387 B.n46 163.367
R1043 B.n387 B.n386 163.367
R1044 B.n386 B.n385 163.367
R1045 B.n385 B.n48 163.367
R1046 B.n381 B.n48 163.367
R1047 B.n381 B.n380 163.367
R1048 B.n380 B.n379 163.367
R1049 B.n379 B.n50 163.367
R1050 B.n375 B.n50 163.367
R1051 B.n375 B.n374 163.367
R1052 B.n374 B.n373 163.367
R1053 B.n373 B.n52 163.367
R1054 B.n369 B.n52 163.367
R1055 B.n369 B.n368 163.367
R1056 B.n368 B.n367 163.367
R1057 B.n367 B.n54 163.367
R1058 B.n363 B.n54 163.367
R1059 B.n363 B.n362 163.367
R1060 B.n362 B.n361 163.367
R1061 B.n472 B.n471 163.367
R1062 B.n472 B.n13 163.367
R1063 B.n476 B.n13 163.367
R1064 B.n477 B.n476 163.367
R1065 B.n478 B.n477 163.367
R1066 B.n478 B.n11 163.367
R1067 B.n482 B.n11 163.367
R1068 B.n483 B.n482 163.367
R1069 B.n484 B.n483 163.367
R1070 B.n484 B.n9 163.367
R1071 B.n488 B.n9 163.367
R1072 B.n489 B.n488 163.367
R1073 B.n490 B.n489 163.367
R1074 B.n490 B.n7 163.367
R1075 B.n494 B.n7 163.367
R1076 B.n495 B.n494 163.367
R1077 B.n496 B.n495 163.367
R1078 B.n496 B.n5 163.367
R1079 B.n500 B.n5 163.367
R1080 B.n501 B.n500 163.367
R1081 B.n502 B.n501 163.367
R1082 B.n502 B.n3 163.367
R1083 B.n506 B.n3 163.367
R1084 B.n507 B.n506 163.367
R1085 B.n134 B.n2 163.367
R1086 B.n137 B.n134 163.367
R1087 B.n138 B.n137 163.367
R1088 B.n139 B.n138 163.367
R1089 B.n139 B.n132 163.367
R1090 B.n143 B.n132 163.367
R1091 B.n144 B.n143 163.367
R1092 B.n145 B.n144 163.367
R1093 B.n145 B.n130 163.367
R1094 B.n149 B.n130 163.367
R1095 B.n150 B.n149 163.367
R1096 B.n151 B.n150 163.367
R1097 B.n151 B.n128 163.367
R1098 B.n155 B.n128 163.367
R1099 B.n156 B.n155 163.367
R1100 B.n157 B.n156 163.367
R1101 B.n157 B.n126 163.367
R1102 B.n161 B.n126 163.367
R1103 B.n162 B.n161 163.367
R1104 B.n163 B.n162 163.367
R1105 B.n163 B.n124 163.367
R1106 B.n167 B.n124 163.367
R1107 B.n168 B.n167 163.367
R1108 B.n169 B.n168 163.367
R1109 B.n219 B.n106 59.5399
R1110 B.n233 B.n100 59.5399
R1111 B.n408 B.n40 59.5399
R1112 B.n34 B.n33 59.5399
R1113 B.n106 B.n105 38.5944
R1114 B.n100 B.n99 38.5944
R1115 B.n40 B.n39 38.5944
R1116 B.n33 B.n32 38.5944
R1117 B.n469 B.n14 31.6883
R1118 B.n360 B.n359 31.6883
R1119 B.n282 B.n281 31.6883
R1120 B.n171 B.n170 31.6883
R1121 B B.n509 18.0485
R1122 B.n473 B.n14 10.6151
R1123 B.n474 B.n473 10.6151
R1124 B.n475 B.n474 10.6151
R1125 B.n475 B.n12 10.6151
R1126 B.n479 B.n12 10.6151
R1127 B.n480 B.n479 10.6151
R1128 B.n481 B.n480 10.6151
R1129 B.n481 B.n10 10.6151
R1130 B.n485 B.n10 10.6151
R1131 B.n486 B.n485 10.6151
R1132 B.n487 B.n486 10.6151
R1133 B.n487 B.n8 10.6151
R1134 B.n491 B.n8 10.6151
R1135 B.n492 B.n491 10.6151
R1136 B.n493 B.n492 10.6151
R1137 B.n493 B.n6 10.6151
R1138 B.n497 B.n6 10.6151
R1139 B.n498 B.n497 10.6151
R1140 B.n499 B.n498 10.6151
R1141 B.n499 B.n4 10.6151
R1142 B.n503 B.n4 10.6151
R1143 B.n504 B.n503 10.6151
R1144 B.n505 B.n504 10.6151
R1145 B.n505 B.n0 10.6151
R1146 B.n469 B.n468 10.6151
R1147 B.n468 B.n467 10.6151
R1148 B.n467 B.n16 10.6151
R1149 B.n463 B.n16 10.6151
R1150 B.n463 B.n462 10.6151
R1151 B.n462 B.n461 10.6151
R1152 B.n461 B.n18 10.6151
R1153 B.n457 B.n18 10.6151
R1154 B.n457 B.n456 10.6151
R1155 B.n456 B.n455 10.6151
R1156 B.n455 B.n20 10.6151
R1157 B.n451 B.n20 10.6151
R1158 B.n451 B.n450 10.6151
R1159 B.n450 B.n449 10.6151
R1160 B.n449 B.n22 10.6151
R1161 B.n445 B.n22 10.6151
R1162 B.n445 B.n444 10.6151
R1163 B.n444 B.n443 10.6151
R1164 B.n443 B.n24 10.6151
R1165 B.n439 B.n24 10.6151
R1166 B.n439 B.n438 10.6151
R1167 B.n438 B.n437 10.6151
R1168 B.n437 B.n26 10.6151
R1169 B.n433 B.n26 10.6151
R1170 B.n433 B.n432 10.6151
R1171 B.n432 B.n431 10.6151
R1172 B.n431 B.n28 10.6151
R1173 B.n427 B.n28 10.6151
R1174 B.n427 B.n426 10.6151
R1175 B.n426 B.n425 10.6151
R1176 B.n425 B.n30 10.6151
R1177 B.n421 B.n420 10.6151
R1178 B.n420 B.n419 10.6151
R1179 B.n419 B.n35 10.6151
R1180 B.n415 B.n35 10.6151
R1181 B.n415 B.n414 10.6151
R1182 B.n414 B.n413 10.6151
R1183 B.n413 B.n37 10.6151
R1184 B.n409 B.n37 10.6151
R1185 B.n407 B.n406 10.6151
R1186 B.n406 B.n41 10.6151
R1187 B.n402 B.n41 10.6151
R1188 B.n402 B.n401 10.6151
R1189 B.n401 B.n400 10.6151
R1190 B.n400 B.n43 10.6151
R1191 B.n396 B.n43 10.6151
R1192 B.n396 B.n395 10.6151
R1193 B.n395 B.n394 10.6151
R1194 B.n394 B.n45 10.6151
R1195 B.n390 B.n45 10.6151
R1196 B.n390 B.n389 10.6151
R1197 B.n389 B.n388 10.6151
R1198 B.n388 B.n47 10.6151
R1199 B.n384 B.n47 10.6151
R1200 B.n384 B.n383 10.6151
R1201 B.n383 B.n382 10.6151
R1202 B.n382 B.n49 10.6151
R1203 B.n378 B.n49 10.6151
R1204 B.n378 B.n377 10.6151
R1205 B.n377 B.n376 10.6151
R1206 B.n376 B.n51 10.6151
R1207 B.n372 B.n51 10.6151
R1208 B.n372 B.n371 10.6151
R1209 B.n371 B.n370 10.6151
R1210 B.n370 B.n53 10.6151
R1211 B.n366 B.n53 10.6151
R1212 B.n366 B.n365 10.6151
R1213 B.n365 B.n364 10.6151
R1214 B.n364 B.n55 10.6151
R1215 B.n360 B.n55 10.6151
R1216 B.n359 B.n358 10.6151
R1217 B.n358 B.n57 10.6151
R1218 B.n354 B.n57 10.6151
R1219 B.n354 B.n353 10.6151
R1220 B.n353 B.n352 10.6151
R1221 B.n352 B.n59 10.6151
R1222 B.n348 B.n59 10.6151
R1223 B.n348 B.n347 10.6151
R1224 B.n347 B.n346 10.6151
R1225 B.n346 B.n61 10.6151
R1226 B.n342 B.n61 10.6151
R1227 B.n342 B.n341 10.6151
R1228 B.n341 B.n340 10.6151
R1229 B.n340 B.n63 10.6151
R1230 B.n336 B.n63 10.6151
R1231 B.n336 B.n335 10.6151
R1232 B.n335 B.n334 10.6151
R1233 B.n334 B.n65 10.6151
R1234 B.n330 B.n65 10.6151
R1235 B.n330 B.n329 10.6151
R1236 B.n329 B.n328 10.6151
R1237 B.n328 B.n67 10.6151
R1238 B.n324 B.n67 10.6151
R1239 B.n324 B.n323 10.6151
R1240 B.n323 B.n322 10.6151
R1241 B.n322 B.n69 10.6151
R1242 B.n318 B.n69 10.6151
R1243 B.n318 B.n317 10.6151
R1244 B.n317 B.n316 10.6151
R1245 B.n316 B.n71 10.6151
R1246 B.n312 B.n71 10.6151
R1247 B.n312 B.n311 10.6151
R1248 B.n311 B.n310 10.6151
R1249 B.n310 B.n73 10.6151
R1250 B.n306 B.n73 10.6151
R1251 B.n306 B.n305 10.6151
R1252 B.n305 B.n304 10.6151
R1253 B.n304 B.n75 10.6151
R1254 B.n300 B.n75 10.6151
R1255 B.n300 B.n299 10.6151
R1256 B.n299 B.n298 10.6151
R1257 B.n298 B.n77 10.6151
R1258 B.n294 B.n77 10.6151
R1259 B.n294 B.n293 10.6151
R1260 B.n293 B.n292 10.6151
R1261 B.n292 B.n79 10.6151
R1262 B.n288 B.n79 10.6151
R1263 B.n288 B.n287 10.6151
R1264 B.n287 B.n286 10.6151
R1265 B.n286 B.n81 10.6151
R1266 B.n282 B.n81 10.6151
R1267 B.n135 B.n1 10.6151
R1268 B.n136 B.n135 10.6151
R1269 B.n136 B.n133 10.6151
R1270 B.n140 B.n133 10.6151
R1271 B.n141 B.n140 10.6151
R1272 B.n142 B.n141 10.6151
R1273 B.n142 B.n131 10.6151
R1274 B.n146 B.n131 10.6151
R1275 B.n147 B.n146 10.6151
R1276 B.n148 B.n147 10.6151
R1277 B.n148 B.n129 10.6151
R1278 B.n152 B.n129 10.6151
R1279 B.n153 B.n152 10.6151
R1280 B.n154 B.n153 10.6151
R1281 B.n154 B.n127 10.6151
R1282 B.n158 B.n127 10.6151
R1283 B.n159 B.n158 10.6151
R1284 B.n160 B.n159 10.6151
R1285 B.n160 B.n125 10.6151
R1286 B.n164 B.n125 10.6151
R1287 B.n165 B.n164 10.6151
R1288 B.n166 B.n165 10.6151
R1289 B.n166 B.n123 10.6151
R1290 B.n170 B.n123 10.6151
R1291 B.n172 B.n171 10.6151
R1292 B.n172 B.n121 10.6151
R1293 B.n176 B.n121 10.6151
R1294 B.n177 B.n176 10.6151
R1295 B.n178 B.n177 10.6151
R1296 B.n178 B.n119 10.6151
R1297 B.n182 B.n119 10.6151
R1298 B.n183 B.n182 10.6151
R1299 B.n184 B.n183 10.6151
R1300 B.n184 B.n117 10.6151
R1301 B.n188 B.n117 10.6151
R1302 B.n189 B.n188 10.6151
R1303 B.n190 B.n189 10.6151
R1304 B.n190 B.n115 10.6151
R1305 B.n194 B.n115 10.6151
R1306 B.n195 B.n194 10.6151
R1307 B.n196 B.n195 10.6151
R1308 B.n196 B.n113 10.6151
R1309 B.n200 B.n113 10.6151
R1310 B.n201 B.n200 10.6151
R1311 B.n202 B.n201 10.6151
R1312 B.n202 B.n111 10.6151
R1313 B.n206 B.n111 10.6151
R1314 B.n207 B.n206 10.6151
R1315 B.n208 B.n207 10.6151
R1316 B.n208 B.n109 10.6151
R1317 B.n212 B.n109 10.6151
R1318 B.n213 B.n212 10.6151
R1319 B.n214 B.n213 10.6151
R1320 B.n214 B.n107 10.6151
R1321 B.n218 B.n107 10.6151
R1322 B.n221 B.n220 10.6151
R1323 B.n221 B.n103 10.6151
R1324 B.n225 B.n103 10.6151
R1325 B.n226 B.n225 10.6151
R1326 B.n227 B.n226 10.6151
R1327 B.n227 B.n101 10.6151
R1328 B.n231 B.n101 10.6151
R1329 B.n232 B.n231 10.6151
R1330 B.n234 B.n97 10.6151
R1331 B.n238 B.n97 10.6151
R1332 B.n239 B.n238 10.6151
R1333 B.n240 B.n239 10.6151
R1334 B.n240 B.n95 10.6151
R1335 B.n244 B.n95 10.6151
R1336 B.n245 B.n244 10.6151
R1337 B.n246 B.n245 10.6151
R1338 B.n246 B.n93 10.6151
R1339 B.n250 B.n93 10.6151
R1340 B.n251 B.n250 10.6151
R1341 B.n252 B.n251 10.6151
R1342 B.n252 B.n91 10.6151
R1343 B.n256 B.n91 10.6151
R1344 B.n257 B.n256 10.6151
R1345 B.n258 B.n257 10.6151
R1346 B.n258 B.n89 10.6151
R1347 B.n262 B.n89 10.6151
R1348 B.n263 B.n262 10.6151
R1349 B.n264 B.n263 10.6151
R1350 B.n264 B.n87 10.6151
R1351 B.n268 B.n87 10.6151
R1352 B.n269 B.n268 10.6151
R1353 B.n270 B.n269 10.6151
R1354 B.n270 B.n85 10.6151
R1355 B.n274 B.n85 10.6151
R1356 B.n275 B.n274 10.6151
R1357 B.n276 B.n275 10.6151
R1358 B.n276 B.n83 10.6151
R1359 B.n280 B.n83 10.6151
R1360 B.n281 B.n280 10.6151
R1361 B.n509 B.n0 8.11757
R1362 B.n509 B.n1 8.11757
R1363 B.n421 B.n34 6.5566
R1364 B.n409 B.n408 6.5566
R1365 B.n220 B.n219 6.5566
R1366 B.n233 B.n232 6.5566
R1367 B.n34 B.n30 4.05904
R1368 B.n408 B.n407 4.05904
R1369 B.n219 B.n218 4.05904
R1370 B.n234 B.n233 4.05904
C0 w_n2164_n2678# VDD1 1.17284f
C1 VP VN 4.87872f
C2 VP w_n2164_n2678# 3.71567f
C3 VTAIL VDD2 4.51522f
C4 VDD1 B 1.00354f
C5 VP B 1.34312f
C6 VTAIL VDD1 4.46732f
C7 VP VTAIL 3.08489f
C8 VDD2 VDD1 0.797061f
C9 VP VDD2 0.334311f
C10 VN w_n2164_n2678# 3.43986f
C11 VP VDD1 3.34295f
C12 VN B 0.889794f
C13 w_n2164_n2678# B 7.12179f
C14 VN VTAIL 3.07078f
C15 VTAIL w_n2164_n2678# 3.17954f
C16 VN VDD2 3.15711f
C17 w_n2164_n2678# VDD2 1.20793f
C18 VTAIL B 3.41416f
C19 VDD2 B 1.04034f
C20 VN VDD1 0.14797f
C21 VDD2 VSUBS 0.718772f
C22 VDD1 VSUBS 4.73294f
C23 VTAIL VSUBS 0.90875f
C24 VN VSUBS 5.00124f
C25 VP VSUBS 1.677325f
C26 B VSUBS 3.171383f
C27 w_n2164_n2678# VSUBS 71.8015f
C28 B.n0 VSUBS 0.006988f
C29 B.n1 VSUBS 0.006988f
C30 B.n2 VSUBS 0.010335f
C31 B.n3 VSUBS 0.007919f
C32 B.n4 VSUBS 0.007919f
C33 B.n5 VSUBS 0.007919f
C34 B.n6 VSUBS 0.007919f
C35 B.n7 VSUBS 0.007919f
C36 B.n8 VSUBS 0.007919f
C37 B.n9 VSUBS 0.007919f
C38 B.n10 VSUBS 0.007919f
C39 B.n11 VSUBS 0.007919f
C40 B.n12 VSUBS 0.007919f
C41 B.n13 VSUBS 0.007919f
C42 B.n14 VSUBS 0.01738f
C43 B.n15 VSUBS 0.007919f
C44 B.n16 VSUBS 0.007919f
C45 B.n17 VSUBS 0.007919f
C46 B.n18 VSUBS 0.007919f
C47 B.n19 VSUBS 0.007919f
C48 B.n20 VSUBS 0.007919f
C49 B.n21 VSUBS 0.007919f
C50 B.n22 VSUBS 0.007919f
C51 B.n23 VSUBS 0.007919f
C52 B.n24 VSUBS 0.007919f
C53 B.n25 VSUBS 0.007919f
C54 B.n26 VSUBS 0.007919f
C55 B.n27 VSUBS 0.007919f
C56 B.n28 VSUBS 0.007919f
C57 B.n29 VSUBS 0.007919f
C58 B.n30 VSUBS 0.005474f
C59 B.n31 VSUBS 0.007919f
C60 B.t1 VSUBS 0.155409f
C61 B.t2 VSUBS 0.178593f
C62 B.t0 VSUBS 0.724265f
C63 B.n32 VSUBS 0.295141f
C64 B.n33 VSUBS 0.222723f
C65 B.n34 VSUBS 0.018349f
C66 B.n35 VSUBS 0.007919f
C67 B.n36 VSUBS 0.007919f
C68 B.n37 VSUBS 0.007919f
C69 B.n38 VSUBS 0.007919f
C70 B.t4 VSUBS 0.155412f
C71 B.t5 VSUBS 0.178595f
C72 B.t3 VSUBS 0.724265f
C73 B.n39 VSUBS 0.295138f
C74 B.n40 VSUBS 0.22272f
C75 B.n41 VSUBS 0.007919f
C76 B.n42 VSUBS 0.007919f
C77 B.n43 VSUBS 0.007919f
C78 B.n44 VSUBS 0.007919f
C79 B.n45 VSUBS 0.007919f
C80 B.n46 VSUBS 0.007919f
C81 B.n47 VSUBS 0.007919f
C82 B.n48 VSUBS 0.007919f
C83 B.n49 VSUBS 0.007919f
C84 B.n50 VSUBS 0.007919f
C85 B.n51 VSUBS 0.007919f
C86 B.n52 VSUBS 0.007919f
C87 B.n53 VSUBS 0.007919f
C88 B.n54 VSUBS 0.007919f
C89 B.n55 VSUBS 0.007919f
C90 B.n56 VSUBS 0.01738f
C91 B.n57 VSUBS 0.007919f
C92 B.n58 VSUBS 0.007919f
C93 B.n59 VSUBS 0.007919f
C94 B.n60 VSUBS 0.007919f
C95 B.n61 VSUBS 0.007919f
C96 B.n62 VSUBS 0.007919f
C97 B.n63 VSUBS 0.007919f
C98 B.n64 VSUBS 0.007919f
C99 B.n65 VSUBS 0.007919f
C100 B.n66 VSUBS 0.007919f
C101 B.n67 VSUBS 0.007919f
C102 B.n68 VSUBS 0.007919f
C103 B.n69 VSUBS 0.007919f
C104 B.n70 VSUBS 0.007919f
C105 B.n71 VSUBS 0.007919f
C106 B.n72 VSUBS 0.007919f
C107 B.n73 VSUBS 0.007919f
C108 B.n74 VSUBS 0.007919f
C109 B.n75 VSUBS 0.007919f
C110 B.n76 VSUBS 0.007919f
C111 B.n77 VSUBS 0.007919f
C112 B.n78 VSUBS 0.007919f
C113 B.n79 VSUBS 0.007919f
C114 B.n80 VSUBS 0.007919f
C115 B.n81 VSUBS 0.007919f
C116 B.n82 VSUBS 0.018956f
C117 B.n83 VSUBS 0.007919f
C118 B.n84 VSUBS 0.007919f
C119 B.n85 VSUBS 0.007919f
C120 B.n86 VSUBS 0.007919f
C121 B.n87 VSUBS 0.007919f
C122 B.n88 VSUBS 0.007919f
C123 B.n89 VSUBS 0.007919f
C124 B.n90 VSUBS 0.007919f
C125 B.n91 VSUBS 0.007919f
C126 B.n92 VSUBS 0.007919f
C127 B.n93 VSUBS 0.007919f
C128 B.n94 VSUBS 0.007919f
C129 B.n95 VSUBS 0.007919f
C130 B.n96 VSUBS 0.007919f
C131 B.n97 VSUBS 0.007919f
C132 B.n98 VSUBS 0.007919f
C133 B.t8 VSUBS 0.155412f
C134 B.t7 VSUBS 0.178595f
C135 B.t6 VSUBS 0.724265f
C136 B.n99 VSUBS 0.295138f
C137 B.n100 VSUBS 0.22272f
C138 B.n101 VSUBS 0.007919f
C139 B.n102 VSUBS 0.007919f
C140 B.n103 VSUBS 0.007919f
C141 B.n104 VSUBS 0.007919f
C142 B.t11 VSUBS 0.155409f
C143 B.t10 VSUBS 0.178593f
C144 B.t9 VSUBS 0.724265f
C145 B.n105 VSUBS 0.295141f
C146 B.n106 VSUBS 0.222723f
C147 B.n107 VSUBS 0.007919f
C148 B.n108 VSUBS 0.007919f
C149 B.n109 VSUBS 0.007919f
C150 B.n110 VSUBS 0.007919f
C151 B.n111 VSUBS 0.007919f
C152 B.n112 VSUBS 0.007919f
C153 B.n113 VSUBS 0.007919f
C154 B.n114 VSUBS 0.007919f
C155 B.n115 VSUBS 0.007919f
C156 B.n116 VSUBS 0.007919f
C157 B.n117 VSUBS 0.007919f
C158 B.n118 VSUBS 0.007919f
C159 B.n119 VSUBS 0.007919f
C160 B.n120 VSUBS 0.007919f
C161 B.n121 VSUBS 0.007919f
C162 B.n122 VSUBS 0.018956f
C163 B.n123 VSUBS 0.007919f
C164 B.n124 VSUBS 0.007919f
C165 B.n125 VSUBS 0.007919f
C166 B.n126 VSUBS 0.007919f
C167 B.n127 VSUBS 0.007919f
C168 B.n128 VSUBS 0.007919f
C169 B.n129 VSUBS 0.007919f
C170 B.n130 VSUBS 0.007919f
C171 B.n131 VSUBS 0.007919f
C172 B.n132 VSUBS 0.007919f
C173 B.n133 VSUBS 0.007919f
C174 B.n134 VSUBS 0.007919f
C175 B.n135 VSUBS 0.007919f
C176 B.n136 VSUBS 0.007919f
C177 B.n137 VSUBS 0.007919f
C178 B.n138 VSUBS 0.007919f
C179 B.n139 VSUBS 0.007919f
C180 B.n140 VSUBS 0.007919f
C181 B.n141 VSUBS 0.007919f
C182 B.n142 VSUBS 0.007919f
C183 B.n143 VSUBS 0.007919f
C184 B.n144 VSUBS 0.007919f
C185 B.n145 VSUBS 0.007919f
C186 B.n146 VSUBS 0.007919f
C187 B.n147 VSUBS 0.007919f
C188 B.n148 VSUBS 0.007919f
C189 B.n149 VSUBS 0.007919f
C190 B.n150 VSUBS 0.007919f
C191 B.n151 VSUBS 0.007919f
C192 B.n152 VSUBS 0.007919f
C193 B.n153 VSUBS 0.007919f
C194 B.n154 VSUBS 0.007919f
C195 B.n155 VSUBS 0.007919f
C196 B.n156 VSUBS 0.007919f
C197 B.n157 VSUBS 0.007919f
C198 B.n158 VSUBS 0.007919f
C199 B.n159 VSUBS 0.007919f
C200 B.n160 VSUBS 0.007919f
C201 B.n161 VSUBS 0.007919f
C202 B.n162 VSUBS 0.007919f
C203 B.n163 VSUBS 0.007919f
C204 B.n164 VSUBS 0.007919f
C205 B.n165 VSUBS 0.007919f
C206 B.n166 VSUBS 0.007919f
C207 B.n167 VSUBS 0.007919f
C208 B.n168 VSUBS 0.007919f
C209 B.n169 VSUBS 0.01738f
C210 B.n170 VSUBS 0.01738f
C211 B.n171 VSUBS 0.018956f
C212 B.n172 VSUBS 0.007919f
C213 B.n173 VSUBS 0.007919f
C214 B.n174 VSUBS 0.007919f
C215 B.n175 VSUBS 0.007919f
C216 B.n176 VSUBS 0.007919f
C217 B.n177 VSUBS 0.007919f
C218 B.n178 VSUBS 0.007919f
C219 B.n179 VSUBS 0.007919f
C220 B.n180 VSUBS 0.007919f
C221 B.n181 VSUBS 0.007919f
C222 B.n182 VSUBS 0.007919f
C223 B.n183 VSUBS 0.007919f
C224 B.n184 VSUBS 0.007919f
C225 B.n185 VSUBS 0.007919f
C226 B.n186 VSUBS 0.007919f
C227 B.n187 VSUBS 0.007919f
C228 B.n188 VSUBS 0.007919f
C229 B.n189 VSUBS 0.007919f
C230 B.n190 VSUBS 0.007919f
C231 B.n191 VSUBS 0.007919f
C232 B.n192 VSUBS 0.007919f
C233 B.n193 VSUBS 0.007919f
C234 B.n194 VSUBS 0.007919f
C235 B.n195 VSUBS 0.007919f
C236 B.n196 VSUBS 0.007919f
C237 B.n197 VSUBS 0.007919f
C238 B.n198 VSUBS 0.007919f
C239 B.n199 VSUBS 0.007919f
C240 B.n200 VSUBS 0.007919f
C241 B.n201 VSUBS 0.007919f
C242 B.n202 VSUBS 0.007919f
C243 B.n203 VSUBS 0.007919f
C244 B.n204 VSUBS 0.007919f
C245 B.n205 VSUBS 0.007919f
C246 B.n206 VSUBS 0.007919f
C247 B.n207 VSUBS 0.007919f
C248 B.n208 VSUBS 0.007919f
C249 B.n209 VSUBS 0.007919f
C250 B.n210 VSUBS 0.007919f
C251 B.n211 VSUBS 0.007919f
C252 B.n212 VSUBS 0.007919f
C253 B.n213 VSUBS 0.007919f
C254 B.n214 VSUBS 0.007919f
C255 B.n215 VSUBS 0.007919f
C256 B.n216 VSUBS 0.007919f
C257 B.n217 VSUBS 0.007919f
C258 B.n218 VSUBS 0.005474f
C259 B.n219 VSUBS 0.018349f
C260 B.n220 VSUBS 0.006405f
C261 B.n221 VSUBS 0.007919f
C262 B.n222 VSUBS 0.007919f
C263 B.n223 VSUBS 0.007919f
C264 B.n224 VSUBS 0.007919f
C265 B.n225 VSUBS 0.007919f
C266 B.n226 VSUBS 0.007919f
C267 B.n227 VSUBS 0.007919f
C268 B.n228 VSUBS 0.007919f
C269 B.n229 VSUBS 0.007919f
C270 B.n230 VSUBS 0.007919f
C271 B.n231 VSUBS 0.007919f
C272 B.n232 VSUBS 0.006405f
C273 B.n233 VSUBS 0.018349f
C274 B.n234 VSUBS 0.005474f
C275 B.n235 VSUBS 0.007919f
C276 B.n236 VSUBS 0.007919f
C277 B.n237 VSUBS 0.007919f
C278 B.n238 VSUBS 0.007919f
C279 B.n239 VSUBS 0.007919f
C280 B.n240 VSUBS 0.007919f
C281 B.n241 VSUBS 0.007919f
C282 B.n242 VSUBS 0.007919f
C283 B.n243 VSUBS 0.007919f
C284 B.n244 VSUBS 0.007919f
C285 B.n245 VSUBS 0.007919f
C286 B.n246 VSUBS 0.007919f
C287 B.n247 VSUBS 0.007919f
C288 B.n248 VSUBS 0.007919f
C289 B.n249 VSUBS 0.007919f
C290 B.n250 VSUBS 0.007919f
C291 B.n251 VSUBS 0.007919f
C292 B.n252 VSUBS 0.007919f
C293 B.n253 VSUBS 0.007919f
C294 B.n254 VSUBS 0.007919f
C295 B.n255 VSUBS 0.007919f
C296 B.n256 VSUBS 0.007919f
C297 B.n257 VSUBS 0.007919f
C298 B.n258 VSUBS 0.007919f
C299 B.n259 VSUBS 0.007919f
C300 B.n260 VSUBS 0.007919f
C301 B.n261 VSUBS 0.007919f
C302 B.n262 VSUBS 0.007919f
C303 B.n263 VSUBS 0.007919f
C304 B.n264 VSUBS 0.007919f
C305 B.n265 VSUBS 0.007919f
C306 B.n266 VSUBS 0.007919f
C307 B.n267 VSUBS 0.007919f
C308 B.n268 VSUBS 0.007919f
C309 B.n269 VSUBS 0.007919f
C310 B.n270 VSUBS 0.007919f
C311 B.n271 VSUBS 0.007919f
C312 B.n272 VSUBS 0.007919f
C313 B.n273 VSUBS 0.007919f
C314 B.n274 VSUBS 0.007919f
C315 B.n275 VSUBS 0.007919f
C316 B.n276 VSUBS 0.007919f
C317 B.n277 VSUBS 0.007919f
C318 B.n278 VSUBS 0.007919f
C319 B.n279 VSUBS 0.007919f
C320 B.n280 VSUBS 0.007919f
C321 B.n281 VSUBS 0.017992f
C322 B.n282 VSUBS 0.018345f
C323 B.n283 VSUBS 0.01738f
C324 B.n284 VSUBS 0.007919f
C325 B.n285 VSUBS 0.007919f
C326 B.n286 VSUBS 0.007919f
C327 B.n287 VSUBS 0.007919f
C328 B.n288 VSUBS 0.007919f
C329 B.n289 VSUBS 0.007919f
C330 B.n290 VSUBS 0.007919f
C331 B.n291 VSUBS 0.007919f
C332 B.n292 VSUBS 0.007919f
C333 B.n293 VSUBS 0.007919f
C334 B.n294 VSUBS 0.007919f
C335 B.n295 VSUBS 0.007919f
C336 B.n296 VSUBS 0.007919f
C337 B.n297 VSUBS 0.007919f
C338 B.n298 VSUBS 0.007919f
C339 B.n299 VSUBS 0.007919f
C340 B.n300 VSUBS 0.007919f
C341 B.n301 VSUBS 0.007919f
C342 B.n302 VSUBS 0.007919f
C343 B.n303 VSUBS 0.007919f
C344 B.n304 VSUBS 0.007919f
C345 B.n305 VSUBS 0.007919f
C346 B.n306 VSUBS 0.007919f
C347 B.n307 VSUBS 0.007919f
C348 B.n308 VSUBS 0.007919f
C349 B.n309 VSUBS 0.007919f
C350 B.n310 VSUBS 0.007919f
C351 B.n311 VSUBS 0.007919f
C352 B.n312 VSUBS 0.007919f
C353 B.n313 VSUBS 0.007919f
C354 B.n314 VSUBS 0.007919f
C355 B.n315 VSUBS 0.007919f
C356 B.n316 VSUBS 0.007919f
C357 B.n317 VSUBS 0.007919f
C358 B.n318 VSUBS 0.007919f
C359 B.n319 VSUBS 0.007919f
C360 B.n320 VSUBS 0.007919f
C361 B.n321 VSUBS 0.007919f
C362 B.n322 VSUBS 0.007919f
C363 B.n323 VSUBS 0.007919f
C364 B.n324 VSUBS 0.007919f
C365 B.n325 VSUBS 0.007919f
C366 B.n326 VSUBS 0.007919f
C367 B.n327 VSUBS 0.007919f
C368 B.n328 VSUBS 0.007919f
C369 B.n329 VSUBS 0.007919f
C370 B.n330 VSUBS 0.007919f
C371 B.n331 VSUBS 0.007919f
C372 B.n332 VSUBS 0.007919f
C373 B.n333 VSUBS 0.007919f
C374 B.n334 VSUBS 0.007919f
C375 B.n335 VSUBS 0.007919f
C376 B.n336 VSUBS 0.007919f
C377 B.n337 VSUBS 0.007919f
C378 B.n338 VSUBS 0.007919f
C379 B.n339 VSUBS 0.007919f
C380 B.n340 VSUBS 0.007919f
C381 B.n341 VSUBS 0.007919f
C382 B.n342 VSUBS 0.007919f
C383 B.n343 VSUBS 0.007919f
C384 B.n344 VSUBS 0.007919f
C385 B.n345 VSUBS 0.007919f
C386 B.n346 VSUBS 0.007919f
C387 B.n347 VSUBS 0.007919f
C388 B.n348 VSUBS 0.007919f
C389 B.n349 VSUBS 0.007919f
C390 B.n350 VSUBS 0.007919f
C391 B.n351 VSUBS 0.007919f
C392 B.n352 VSUBS 0.007919f
C393 B.n353 VSUBS 0.007919f
C394 B.n354 VSUBS 0.007919f
C395 B.n355 VSUBS 0.007919f
C396 B.n356 VSUBS 0.007919f
C397 B.n357 VSUBS 0.007919f
C398 B.n358 VSUBS 0.007919f
C399 B.n359 VSUBS 0.01738f
C400 B.n360 VSUBS 0.018956f
C401 B.n361 VSUBS 0.018956f
C402 B.n362 VSUBS 0.007919f
C403 B.n363 VSUBS 0.007919f
C404 B.n364 VSUBS 0.007919f
C405 B.n365 VSUBS 0.007919f
C406 B.n366 VSUBS 0.007919f
C407 B.n367 VSUBS 0.007919f
C408 B.n368 VSUBS 0.007919f
C409 B.n369 VSUBS 0.007919f
C410 B.n370 VSUBS 0.007919f
C411 B.n371 VSUBS 0.007919f
C412 B.n372 VSUBS 0.007919f
C413 B.n373 VSUBS 0.007919f
C414 B.n374 VSUBS 0.007919f
C415 B.n375 VSUBS 0.007919f
C416 B.n376 VSUBS 0.007919f
C417 B.n377 VSUBS 0.007919f
C418 B.n378 VSUBS 0.007919f
C419 B.n379 VSUBS 0.007919f
C420 B.n380 VSUBS 0.007919f
C421 B.n381 VSUBS 0.007919f
C422 B.n382 VSUBS 0.007919f
C423 B.n383 VSUBS 0.007919f
C424 B.n384 VSUBS 0.007919f
C425 B.n385 VSUBS 0.007919f
C426 B.n386 VSUBS 0.007919f
C427 B.n387 VSUBS 0.007919f
C428 B.n388 VSUBS 0.007919f
C429 B.n389 VSUBS 0.007919f
C430 B.n390 VSUBS 0.007919f
C431 B.n391 VSUBS 0.007919f
C432 B.n392 VSUBS 0.007919f
C433 B.n393 VSUBS 0.007919f
C434 B.n394 VSUBS 0.007919f
C435 B.n395 VSUBS 0.007919f
C436 B.n396 VSUBS 0.007919f
C437 B.n397 VSUBS 0.007919f
C438 B.n398 VSUBS 0.007919f
C439 B.n399 VSUBS 0.007919f
C440 B.n400 VSUBS 0.007919f
C441 B.n401 VSUBS 0.007919f
C442 B.n402 VSUBS 0.007919f
C443 B.n403 VSUBS 0.007919f
C444 B.n404 VSUBS 0.007919f
C445 B.n405 VSUBS 0.007919f
C446 B.n406 VSUBS 0.007919f
C447 B.n407 VSUBS 0.005474f
C448 B.n408 VSUBS 0.018349f
C449 B.n409 VSUBS 0.006405f
C450 B.n410 VSUBS 0.007919f
C451 B.n411 VSUBS 0.007919f
C452 B.n412 VSUBS 0.007919f
C453 B.n413 VSUBS 0.007919f
C454 B.n414 VSUBS 0.007919f
C455 B.n415 VSUBS 0.007919f
C456 B.n416 VSUBS 0.007919f
C457 B.n417 VSUBS 0.007919f
C458 B.n418 VSUBS 0.007919f
C459 B.n419 VSUBS 0.007919f
C460 B.n420 VSUBS 0.007919f
C461 B.n421 VSUBS 0.006405f
C462 B.n422 VSUBS 0.007919f
C463 B.n423 VSUBS 0.007919f
C464 B.n424 VSUBS 0.007919f
C465 B.n425 VSUBS 0.007919f
C466 B.n426 VSUBS 0.007919f
C467 B.n427 VSUBS 0.007919f
C468 B.n428 VSUBS 0.007919f
C469 B.n429 VSUBS 0.007919f
C470 B.n430 VSUBS 0.007919f
C471 B.n431 VSUBS 0.007919f
C472 B.n432 VSUBS 0.007919f
C473 B.n433 VSUBS 0.007919f
C474 B.n434 VSUBS 0.007919f
C475 B.n435 VSUBS 0.007919f
C476 B.n436 VSUBS 0.007919f
C477 B.n437 VSUBS 0.007919f
C478 B.n438 VSUBS 0.007919f
C479 B.n439 VSUBS 0.007919f
C480 B.n440 VSUBS 0.007919f
C481 B.n441 VSUBS 0.007919f
C482 B.n442 VSUBS 0.007919f
C483 B.n443 VSUBS 0.007919f
C484 B.n444 VSUBS 0.007919f
C485 B.n445 VSUBS 0.007919f
C486 B.n446 VSUBS 0.007919f
C487 B.n447 VSUBS 0.007919f
C488 B.n448 VSUBS 0.007919f
C489 B.n449 VSUBS 0.007919f
C490 B.n450 VSUBS 0.007919f
C491 B.n451 VSUBS 0.007919f
C492 B.n452 VSUBS 0.007919f
C493 B.n453 VSUBS 0.007919f
C494 B.n454 VSUBS 0.007919f
C495 B.n455 VSUBS 0.007919f
C496 B.n456 VSUBS 0.007919f
C497 B.n457 VSUBS 0.007919f
C498 B.n458 VSUBS 0.007919f
C499 B.n459 VSUBS 0.007919f
C500 B.n460 VSUBS 0.007919f
C501 B.n461 VSUBS 0.007919f
C502 B.n462 VSUBS 0.007919f
C503 B.n463 VSUBS 0.007919f
C504 B.n464 VSUBS 0.007919f
C505 B.n465 VSUBS 0.007919f
C506 B.n466 VSUBS 0.007919f
C507 B.n467 VSUBS 0.007919f
C508 B.n468 VSUBS 0.007919f
C509 B.n469 VSUBS 0.018956f
C510 B.n470 VSUBS 0.018956f
C511 B.n471 VSUBS 0.01738f
C512 B.n472 VSUBS 0.007919f
C513 B.n473 VSUBS 0.007919f
C514 B.n474 VSUBS 0.007919f
C515 B.n475 VSUBS 0.007919f
C516 B.n476 VSUBS 0.007919f
C517 B.n477 VSUBS 0.007919f
C518 B.n478 VSUBS 0.007919f
C519 B.n479 VSUBS 0.007919f
C520 B.n480 VSUBS 0.007919f
C521 B.n481 VSUBS 0.007919f
C522 B.n482 VSUBS 0.007919f
C523 B.n483 VSUBS 0.007919f
C524 B.n484 VSUBS 0.007919f
C525 B.n485 VSUBS 0.007919f
C526 B.n486 VSUBS 0.007919f
C527 B.n487 VSUBS 0.007919f
C528 B.n488 VSUBS 0.007919f
C529 B.n489 VSUBS 0.007919f
C530 B.n490 VSUBS 0.007919f
C531 B.n491 VSUBS 0.007919f
C532 B.n492 VSUBS 0.007919f
C533 B.n493 VSUBS 0.007919f
C534 B.n494 VSUBS 0.007919f
C535 B.n495 VSUBS 0.007919f
C536 B.n496 VSUBS 0.007919f
C537 B.n497 VSUBS 0.007919f
C538 B.n498 VSUBS 0.007919f
C539 B.n499 VSUBS 0.007919f
C540 B.n500 VSUBS 0.007919f
C541 B.n501 VSUBS 0.007919f
C542 B.n502 VSUBS 0.007919f
C543 B.n503 VSUBS 0.007919f
C544 B.n504 VSUBS 0.007919f
C545 B.n505 VSUBS 0.007919f
C546 B.n506 VSUBS 0.007919f
C547 B.n507 VSUBS 0.010335f
C548 B.n508 VSUBS 0.011009f
C549 B.n509 VSUBS 0.021892f
C550 VDD2.t0 VSUBS 0.182231f
C551 VDD2.t3 VSUBS 0.182231f
C552 VDD2.n0 VSUBS 1.84116f
C553 VDD2.t1 VSUBS 0.182231f
C554 VDD2.t2 VSUBS 0.182231f
C555 VDD2.n1 VSUBS 1.33474f
C556 VDD2.n2 VSUBS 3.64028f
C557 VN.t3 VSUBS 1.90468f
C558 VN.t0 VSUBS 1.90241f
C559 VN.n0 VSUBS 1.39021f
C560 VN.t1 VSUBS 1.90468f
C561 VN.t2 VSUBS 1.90241f
C562 VN.n1 VSUBS 3.07501f
C563 VTAIL.n0 VSUBS 0.024964f
C564 VTAIL.n1 VSUBS 0.024414f
C565 VTAIL.n2 VSUBS 0.013119f
C566 VTAIL.n3 VSUBS 0.031009f
C567 VTAIL.n4 VSUBS 0.013891f
C568 VTAIL.n5 VSUBS 0.024414f
C569 VTAIL.n6 VSUBS 0.013119f
C570 VTAIL.n7 VSUBS 0.031009f
C571 VTAIL.n8 VSUBS 0.013891f
C572 VTAIL.n9 VSUBS 0.024414f
C573 VTAIL.n10 VSUBS 0.013119f
C574 VTAIL.n11 VSUBS 0.031009f
C575 VTAIL.n12 VSUBS 0.013891f
C576 VTAIL.n13 VSUBS 0.154234f
C577 VTAIL.t0 VSUBS 0.066587f
C578 VTAIL.n14 VSUBS 0.023256f
C579 VTAIL.n15 VSUBS 0.023326f
C580 VTAIL.n16 VSUBS 0.013119f
C581 VTAIL.n17 VSUBS 0.830384f
C582 VTAIL.n18 VSUBS 0.024414f
C583 VTAIL.n19 VSUBS 0.013119f
C584 VTAIL.n20 VSUBS 0.013891f
C585 VTAIL.n21 VSUBS 0.031009f
C586 VTAIL.n22 VSUBS 0.031009f
C587 VTAIL.n23 VSUBS 0.013891f
C588 VTAIL.n24 VSUBS 0.013119f
C589 VTAIL.n25 VSUBS 0.024414f
C590 VTAIL.n26 VSUBS 0.024414f
C591 VTAIL.n27 VSUBS 0.013119f
C592 VTAIL.n28 VSUBS 0.013891f
C593 VTAIL.n29 VSUBS 0.031009f
C594 VTAIL.n30 VSUBS 0.031009f
C595 VTAIL.n31 VSUBS 0.031009f
C596 VTAIL.n32 VSUBS 0.013891f
C597 VTAIL.n33 VSUBS 0.013119f
C598 VTAIL.n34 VSUBS 0.024414f
C599 VTAIL.n35 VSUBS 0.024414f
C600 VTAIL.n36 VSUBS 0.013119f
C601 VTAIL.n37 VSUBS 0.013505f
C602 VTAIL.n38 VSUBS 0.013505f
C603 VTAIL.n39 VSUBS 0.031009f
C604 VTAIL.n40 VSUBS 0.068728f
C605 VTAIL.n41 VSUBS 0.013891f
C606 VTAIL.n42 VSUBS 0.013119f
C607 VTAIL.n43 VSUBS 0.057432f
C608 VTAIL.n44 VSUBS 0.034312f
C609 VTAIL.n45 VSUBS 0.130431f
C610 VTAIL.n46 VSUBS 0.024964f
C611 VTAIL.n47 VSUBS 0.024414f
C612 VTAIL.n48 VSUBS 0.013119f
C613 VTAIL.n49 VSUBS 0.031009f
C614 VTAIL.n50 VSUBS 0.013891f
C615 VTAIL.n51 VSUBS 0.024414f
C616 VTAIL.n52 VSUBS 0.013119f
C617 VTAIL.n53 VSUBS 0.031009f
C618 VTAIL.n54 VSUBS 0.013891f
C619 VTAIL.n55 VSUBS 0.024414f
C620 VTAIL.n56 VSUBS 0.013119f
C621 VTAIL.n57 VSUBS 0.031009f
C622 VTAIL.n58 VSUBS 0.013891f
C623 VTAIL.n59 VSUBS 0.154234f
C624 VTAIL.t6 VSUBS 0.066587f
C625 VTAIL.n60 VSUBS 0.023256f
C626 VTAIL.n61 VSUBS 0.023326f
C627 VTAIL.n62 VSUBS 0.013119f
C628 VTAIL.n63 VSUBS 0.830384f
C629 VTAIL.n64 VSUBS 0.024414f
C630 VTAIL.n65 VSUBS 0.013119f
C631 VTAIL.n66 VSUBS 0.013891f
C632 VTAIL.n67 VSUBS 0.031009f
C633 VTAIL.n68 VSUBS 0.031009f
C634 VTAIL.n69 VSUBS 0.013891f
C635 VTAIL.n70 VSUBS 0.013119f
C636 VTAIL.n71 VSUBS 0.024414f
C637 VTAIL.n72 VSUBS 0.024414f
C638 VTAIL.n73 VSUBS 0.013119f
C639 VTAIL.n74 VSUBS 0.013891f
C640 VTAIL.n75 VSUBS 0.031009f
C641 VTAIL.n76 VSUBS 0.031009f
C642 VTAIL.n77 VSUBS 0.031009f
C643 VTAIL.n78 VSUBS 0.013891f
C644 VTAIL.n79 VSUBS 0.013119f
C645 VTAIL.n80 VSUBS 0.024414f
C646 VTAIL.n81 VSUBS 0.024414f
C647 VTAIL.n82 VSUBS 0.013119f
C648 VTAIL.n83 VSUBS 0.013505f
C649 VTAIL.n84 VSUBS 0.013505f
C650 VTAIL.n85 VSUBS 0.031009f
C651 VTAIL.n86 VSUBS 0.068728f
C652 VTAIL.n87 VSUBS 0.013891f
C653 VTAIL.n88 VSUBS 0.013119f
C654 VTAIL.n89 VSUBS 0.057432f
C655 VTAIL.n90 VSUBS 0.034312f
C656 VTAIL.n91 VSUBS 0.193331f
C657 VTAIL.n92 VSUBS 0.024964f
C658 VTAIL.n93 VSUBS 0.024414f
C659 VTAIL.n94 VSUBS 0.013119f
C660 VTAIL.n95 VSUBS 0.031009f
C661 VTAIL.n96 VSUBS 0.013891f
C662 VTAIL.n97 VSUBS 0.024414f
C663 VTAIL.n98 VSUBS 0.013119f
C664 VTAIL.n99 VSUBS 0.031009f
C665 VTAIL.n100 VSUBS 0.013891f
C666 VTAIL.n101 VSUBS 0.024414f
C667 VTAIL.n102 VSUBS 0.013119f
C668 VTAIL.n103 VSUBS 0.031009f
C669 VTAIL.n104 VSUBS 0.013891f
C670 VTAIL.n105 VSUBS 0.154234f
C671 VTAIL.t4 VSUBS 0.066587f
C672 VTAIL.n106 VSUBS 0.023256f
C673 VTAIL.n107 VSUBS 0.023326f
C674 VTAIL.n108 VSUBS 0.013119f
C675 VTAIL.n109 VSUBS 0.830384f
C676 VTAIL.n110 VSUBS 0.024414f
C677 VTAIL.n111 VSUBS 0.013119f
C678 VTAIL.n112 VSUBS 0.013891f
C679 VTAIL.n113 VSUBS 0.031009f
C680 VTAIL.n114 VSUBS 0.031009f
C681 VTAIL.n115 VSUBS 0.013891f
C682 VTAIL.n116 VSUBS 0.013119f
C683 VTAIL.n117 VSUBS 0.024414f
C684 VTAIL.n118 VSUBS 0.024414f
C685 VTAIL.n119 VSUBS 0.013119f
C686 VTAIL.n120 VSUBS 0.013891f
C687 VTAIL.n121 VSUBS 0.031009f
C688 VTAIL.n122 VSUBS 0.031009f
C689 VTAIL.n123 VSUBS 0.031009f
C690 VTAIL.n124 VSUBS 0.013891f
C691 VTAIL.n125 VSUBS 0.013119f
C692 VTAIL.n126 VSUBS 0.024414f
C693 VTAIL.n127 VSUBS 0.024414f
C694 VTAIL.n128 VSUBS 0.013119f
C695 VTAIL.n129 VSUBS 0.013505f
C696 VTAIL.n130 VSUBS 0.013505f
C697 VTAIL.n131 VSUBS 0.031009f
C698 VTAIL.n132 VSUBS 0.068728f
C699 VTAIL.n133 VSUBS 0.013891f
C700 VTAIL.n134 VSUBS 0.013119f
C701 VTAIL.n135 VSUBS 0.057432f
C702 VTAIL.n136 VSUBS 0.034312f
C703 VTAIL.n137 VSUBS 1.20279f
C704 VTAIL.n138 VSUBS 0.024964f
C705 VTAIL.n139 VSUBS 0.024414f
C706 VTAIL.n140 VSUBS 0.013119f
C707 VTAIL.n141 VSUBS 0.031009f
C708 VTAIL.n142 VSUBS 0.013891f
C709 VTAIL.n143 VSUBS 0.024414f
C710 VTAIL.n144 VSUBS 0.013119f
C711 VTAIL.n145 VSUBS 0.031009f
C712 VTAIL.n146 VSUBS 0.031009f
C713 VTAIL.n147 VSUBS 0.013891f
C714 VTAIL.n148 VSUBS 0.024414f
C715 VTAIL.n149 VSUBS 0.013119f
C716 VTAIL.n150 VSUBS 0.031009f
C717 VTAIL.n151 VSUBS 0.013891f
C718 VTAIL.n152 VSUBS 0.154234f
C719 VTAIL.t1 VSUBS 0.066587f
C720 VTAIL.n153 VSUBS 0.023256f
C721 VTAIL.n154 VSUBS 0.023326f
C722 VTAIL.n155 VSUBS 0.013119f
C723 VTAIL.n156 VSUBS 0.830384f
C724 VTAIL.n157 VSUBS 0.024414f
C725 VTAIL.n158 VSUBS 0.013119f
C726 VTAIL.n159 VSUBS 0.013891f
C727 VTAIL.n160 VSUBS 0.031009f
C728 VTAIL.n161 VSUBS 0.031009f
C729 VTAIL.n162 VSUBS 0.013891f
C730 VTAIL.n163 VSUBS 0.013119f
C731 VTAIL.n164 VSUBS 0.024414f
C732 VTAIL.n165 VSUBS 0.024414f
C733 VTAIL.n166 VSUBS 0.013119f
C734 VTAIL.n167 VSUBS 0.013891f
C735 VTAIL.n168 VSUBS 0.031009f
C736 VTAIL.n169 VSUBS 0.031009f
C737 VTAIL.n170 VSUBS 0.013891f
C738 VTAIL.n171 VSUBS 0.013119f
C739 VTAIL.n172 VSUBS 0.024414f
C740 VTAIL.n173 VSUBS 0.024414f
C741 VTAIL.n174 VSUBS 0.013119f
C742 VTAIL.n175 VSUBS 0.013505f
C743 VTAIL.n176 VSUBS 0.013505f
C744 VTAIL.n177 VSUBS 0.031009f
C745 VTAIL.n178 VSUBS 0.068728f
C746 VTAIL.n179 VSUBS 0.013891f
C747 VTAIL.n180 VSUBS 0.013119f
C748 VTAIL.n181 VSUBS 0.057432f
C749 VTAIL.n182 VSUBS 0.034312f
C750 VTAIL.n183 VSUBS 1.20279f
C751 VTAIL.n184 VSUBS 0.024964f
C752 VTAIL.n185 VSUBS 0.024414f
C753 VTAIL.n186 VSUBS 0.013119f
C754 VTAIL.n187 VSUBS 0.031009f
C755 VTAIL.n188 VSUBS 0.013891f
C756 VTAIL.n189 VSUBS 0.024414f
C757 VTAIL.n190 VSUBS 0.013119f
C758 VTAIL.n191 VSUBS 0.031009f
C759 VTAIL.n192 VSUBS 0.031009f
C760 VTAIL.n193 VSUBS 0.013891f
C761 VTAIL.n194 VSUBS 0.024414f
C762 VTAIL.n195 VSUBS 0.013119f
C763 VTAIL.n196 VSUBS 0.031009f
C764 VTAIL.n197 VSUBS 0.013891f
C765 VTAIL.n198 VSUBS 0.154234f
C766 VTAIL.t2 VSUBS 0.066587f
C767 VTAIL.n199 VSUBS 0.023256f
C768 VTAIL.n200 VSUBS 0.023326f
C769 VTAIL.n201 VSUBS 0.013119f
C770 VTAIL.n202 VSUBS 0.830384f
C771 VTAIL.n203 VSUBS 0.024414f
C772 VTAIL.n204 VSUBS 0.013119f
C773 VTAIL.n205 VSUBS 0.013891f
C774 VTAIL.n206 VSUBS 0.031009f
C775 VTAIL.n207 VSUBS 0.031009f
C776 VTAIL.n208 VSUBS 0.013891f
C777 VTAIL.n209 VSUBS 0.013119f
C778 VTAIL.n210 VSUBS 0.024414f
C779 VTAIL.n211 VSUBS 0.024414f
C780 VTAIL.n212 VSUBS 0.013119f
C781 VTAIL.n213 VSUBS 0.013891f
C782 VTAIL.n214 VSUBS 0.031009f
C783 VTAIL.n215 VSUBS 0.031009f
C784 VTAIL.n216 VSUBS 0.013891f
C785 VTAIL.n217 VSUBS 0.013119f
C786 VTAIL.n218 VSUBS 0.024414f
C787 VTAIL.n219 VSUBS 0.024414f
C788 VTAIL.n220 VSUBS 0.013119f
C789 VTAIL.n221 VSUBS 0.013505f
C790 VTAIL.n222 VSUBS 0.013505f
C791 VTAIL.n223 VSUBS 0.031009f
C792 VTAIL.n224 VSUBS 0.068728f
C793 VTAIL.n225 VSUBS 0.013891f
C794 VTAIL.n226 VSUBS 0.013119f
C795 VTAIL.n227 VSUBS 0.057432f
C796 VTAIL.n228 VSUBS 0.034312f
C797 VTAIL.n229 VSUBS 0.193331f
C798 VTAIL.n230 VSUBS 0.024964f
C799 VTAIL.n231 VSUBS 0.024414f
C800 VTAIL.n232 VSUBS 0.013119f
C801 VTAIL.n233 VSUBS 0.031009f
C802 VTAIL.n234 VSUBS 0.013891f
C803 VTAIL.n235 VSUBS 0.024414f
C804 VTAIL.n236 VSUBS 0.013119f
C805 VTAIL.n237 VSUBS 0.031009f
C806 VTAIL.n238 VSUBS 0.031009f
C807 VTAIL.n239 VSUBS 0.013891f
C808 VTAIL.n240 VSUBS 0.024414f
C809 VTAIL.n241 VSUBS 0.013119f
C810 VTAIL.n242 VSUBS 0.031009f
C811 VTAIL.n243 VSUBS 0.013891f
C812 VTAIL.n244 VSUBS 0.154234f
C813 VTAIL.t7 VSUBS 0.066587f
C814 VTAIL.n245 VSUBS 0.023256f
C815 VTAIL.n246 VSUBS 0.023326f
C816 VTAIL.n247 VSUBS 0.013119f
C817 VTAIL.n248 VSUBS 0.830384f
C818 VTAIL.n249 VSUBS 0.024414f
C819 VTAIL.n250 VSUBS 0.013119f
C820 VTAIL.n251 VSUBS 0.013891f
C821 VTAIL.n252 VSUBS 0.031009f
C822 VTAIL.n253 VSUBS 0.031009f
C823 VTAIL.n254 VSUBS 0.013891f
C824 VTAIL.n255 VSUBS 0.013119f
C825 VTAIL.n256 VSUBS 0.024414f
C826 VTAIL.n257 VSUBS 0.024414f
C827 VTAIL.n258 VSUBS 0.013119f
C828 VTAIL.n259 VSUBS 0.013891f
C829 VTAIL.n260 VSUBS 0.031009f
C830 VTAIL.n261 VSUBS 0.031009f
C831 VTAIL.n262 VSUBS 0.013891f
C832 VTAIL.n263 VSUBS 0.013119f
C833 VTAIL.n264 VSUBS 0.024414f
C834 VTAIL.n265 VSUBS 0.024414f
C835 VTAIL.n266 VSUBS 0.013119f
C836 VTAIL.n267 VSUBS 0.013505f
C837 VTAIL.n268 VSUBS 0.013505f
C838 VTAIL.n269 VSUBS 0.031009f
C839 VTAIL.n270 VSUBS 0.068728f
C840 VTAIL.n271 VSUBS 0.013891f
C841 VTAIL.n272 VSUBS 0.013119f
C842 VTAIL.n273 VSUBS 0.057432f
C843 VTAIL.n274 VSUBS 0.034312f
C844 VTAIL.n275 VSUBS 0.193331f
C845 VTAIL.n276 VSUBS 0.024964f
C846 VTAIL.n277 VSUBS 0.024414f
C847 VTAIL.n278 VSUBS 0.013119f
C848 VTAIL.n279 VSUBS 0.031009f
C849 VTAIL.n280 VSUBS 0.013891f
C850 VTAIL.n281 VSUBS 0.024414f
C851 VTAIL.n282 VSUBS 0.013119f
C852 VTAIL.n283 VSUBS 0.031009f
C853 VTAIL.n284 VSUBS 0.031009f
C854 VTAIL.n285 VSUBS 0.013891f
C855 VTAIL.n286 VSUBS 0.024414f
C856 VTAIL.n287 VSUBS 0.013119f
C857 VTAIL.n288 VSUBS 0.031009f
C858 VTAIL.n289 VSUBS 0.013891f
C859 VTAIL.n290 VSUBS 0.154234f
C860 VTAIL.t5 VSUBS 0.066587f
C861 VTAIL.n291 VSUBS 0.023256f
C862 VTAIL.n292 VSUBS 0.023326f
C863 VTAIL.n293 VSUBS 0.013119f
C864 VTAIL.n294 VSUBS 0.830384f
C865 VTAIL.n295 VSUBS 0.024414f
C866 VTAIL.n296 VSUBS 0.013119f
C867 VTAIL.n297 VSUBS 0.013891f
C868 VTAIL.n298 VSUBS 0.031009f
C869 VTAIL.n299 VSUBS 0.031009f
C870 VTAIL.n300 VSUBS 0.013891f
C871 VTAIL.n301 VSUBS 0.013119f
C872 VTAIL.n302 VSUBS 0.024414f
C873 VTAIL.n303 VSUBS 0.024414f
C874 VTAIL.n304 VSUBS 0.013119f
C875 VTAIL.n305 VSUBS 0.013891f
C876 VTAIL.n306 VSUBS 0.031009f
C877 VTAIL.n307 VSUBS 0.031009f
C878 VTAIL.n308 VSUBS 0.013891f
C879 VTAIL.n309 VSUBS 0.013119f
C880 VTAIL.n310 VSUBS 0.024414f
C881 VTAIL.n311 VSUBS 0.024414f
C882 VTAIL.n312 VSUBS 0.013119f
C883 VTAIL.n313 VSUBS 0.013505f
C884 VTAIL.n314 VSUBS 0.013505f
C885 VTAIL.n315 VSUBS 0.031009f
C886 VTAIL.n316 VSUBS 0.068728f
C887 VTAIL.n317 VSUBS 0.013891f
C888 VTAIL.n318 VSUBS 0.013119f
C889 VTAIL.n319 VSUBS 0.057432f
C890 VTAIL.n320 VSUBS 0.034312f
C891 VTAIL.n321 VSUBS 1.20279f
C892 VTAIL.n322 VSUBS 0.024964f
C893 VTAIL.n323 VSUBS 0.024414f
C894 VTAIL.n324 VSUBS 0.013119f
C895 VTAIL.n325 VSUBS 0.031009f
C896 VTAIL.n326 VSUBS 0.013891f
C897 VTAIL.n327 VSUBS 0.024414f
C898 VTAIL.n328 VSUBS 0.013119f
C899 VTAIL.n329 VSUBS 0.031009f
C900 VTAIL.n330 VSUBS 0.013891f
C901 VTAIL.n331 VSUBS 0.024414f
C902 VTAIL.n332 VSUBS 0.013119f
C903 VTAIL.n333 VSUBS 0.031009f
C904 VTAIL.n334 VSUBS 0.013891f
C905 VTAIL.n335 VSUBS 0.154234f
C906 VTAIL.t3 VSUBS 0.066587f
C907 VTAIL.n336 VSUBS 0.023256f
C908 VTAIL.n337 VSUBS 0.023326f
C909 VTAIL.n338 VSUBS 0.013119f
C910 VTAIL.n339 VSUBS 0.830384f
C911 VTAIL.n340 VSUBS 0.024414f
C912 VTAIL.n341 VSUBS 0.013119f
C913 VTAIL.n342 VSUBS 0.013891f
C914 VTAIL.n343 VSUBS 0.031009f
C915 VTAIL.n344 VSUBS 0.031009f
C916 VTAIL.n345 VSUBS 0.013891f
C917 VTAIL.n346 VSUBS 0.013119f
C918 VTAIL.n347 VSUBS 0.024414f
C919 VTAIL.n348 VSUBS 0.024414f
C920 VTAIL.n349 VSUBS 0.013119f
C921 VTAIL.n350 VSUBS 0.013891f
C922 VTAIL.n351 VSUBS 0.031009f
C923 VTAIL.n352 VSUBS 0.031009f
C924 VTAIL.n353 VSUBS 0.031009f
C925 VTAIL.n354 VSUBS 0.013891f
C926 VTAIL.n355 VSUBS 0.013119f
C927 VTAIL.n356 VSUBS 0.024414f
C928 VTAIL.n357 VSUBS 0.024414f
C929 VTAIL.n358 VSUBS 0.013119f
C930 VTAIL.n359 VSUBS 0.013505f
C931 VTAIL.n360 VSUBS 0.013505f
C932 VTAIL.n361 VSUBS 0.031009f
C933 VTAIL.n362 VSUBS 0.068728f
C934 VTAIL.n363 VSUBS 0.013891f
C935 VTAIL.n364 VSUBS 0.013119f
C936 VTAIL.n365 VSUBS 0.057432f
C937 VTAIL.n366 VSUBS 0.034312f
C938 VTAIL.n367 VSUBS 1.13074f
C939 VDD1.t0 VSUBS 0.18224f
C940 VDD1.t1 VSUBS 0.18224f
C941 VDD1.n0 VSUBS 1.33526f
C942 VDD1.t2 VSUBS 0.18224f
C943 VDD1.t3 VSUBS 0.18224f
C944 VDD1.n1 VSUBS 1.86334f
C945 VP.n0 VSUBS 0.061265f
C946 VP.t1 VSUBS 1.77628f
C947 VP.n1 VSUBS 0.091928f
C948 VP.t2 VSUBS 1.96305f
C949 VP.t0 VSUBS 1.96539f
C950 VP.n2 VSUBS 3.14981f
C951 VP.t3 VSUBS 1.77628f
C952 VP.n3 VSUBS 0.78911f
C953 VP.n4 VSUBS 2.30465f
C954 VP.n5 VSUBS 0.061265f
C955 VP.n6 VSUBS 0.046469f
C956 VP.n7 VSUBS 0.037566f
C957 VP.n8 VSUBS 0.091928f
C958 VP.n9 VSUBS 0.78911f
C959 VP.n10 VSUBS 0.048461f
.ends

