* NGSPICE file created from diff_pair_sample_1102.ext - technology: sky130A

.subckt diff_pair_sample_1102 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t3 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=1.72
X1 VTAIL.t3 VN.t0 VDD2.t3 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=1.72
X2 B.t11 B.t9 B.t10 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=1.72
X3 B.t8 B.t6 B.t7 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=1.72
X4 VDD1.t1 VP.t1 VTAIL.t6 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=1.72
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=1.72
X6 VDD2.t1 VN.t2 VTAIL.t1 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=1.72
X7 VTAIL.t5 VP.t2 VDD1.t0 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=1.72
X8 VDD1.t2 VP.t3 VTAIL.t4 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=1.72
X9 B.t5 B.t3 B.t4 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=1.72
X10 B.t2 B.t0 B.t1 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=1.72
X11 VTAIL.t2 VN.t3 VDD2.t0 w_n2200_n1868# sky130_fd_pr__pfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=1.72
R0 VP.n5 VP.n4 184.662
R1 VP.n14 VP.n13 184.662
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n3 VP.t0 98.4663
R8 VP.n3 VP.t3 98.0424
R9 VP.n5 VP.t2 63.0528
R10 VP.n13 VP.t1 63.0528
R11 VP.n4 VP.n3 47.2758
R12 VP.n7 VP.n1 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n7 VP.n6 24.5923
R15 VP.n12 VP.n11 24.5923
R16 VP.n6 VP.n5 1.23009
R17 VP.n13 VP.n12 1.23009
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VDD1 VDD1.n1 136.337
R26 VDD1 VDD1.n0 102.975
R27 VDD1.n0 VDD1.t3 7.22383
R28 VDD1.n0 VDD1.t2 7.22383
R29 VDD1.n1 VDD1.t0 7.22383
R30 VDD1.n1 VDD1.t1 7.22383
R31 VTAIL.n186 VTAIL.n168 756.745
R32 VTAIL.n18 VTAIL.n0 756.745
R33 VTAIL.n42 VTAIL.n24 756.745
R34 VTAIL.n66 VTAIL.n48 756.745
R35 VTAIL.n162 VTAIL.n144 756.745
R36 VTAIL.n138 VTAIL.n120 756.745
R37 VTAIL.n114 VTAIL.n96 756.745
R38 VTAIL.n90 VTAIL.n72 756.745
R39 VTAIL.n177 VTAIL.n176 585
R40 VTAIL.n179 VTAIL.n178 585
R41 VTAIL.n172 VTAIL.n171 585
R42 VTAIL.n185 VTAIL.n184 585
R43 VTAIL.n187 VTAIL.n186 585
R44 VTAIL.n9 VTAIL.n8 585
R45 VTAIL.n11 VTAIL.n10 585
R46 VTAIL.n4 VTAIL.n3 585
R47 VTAIL.n17 VTAIL.n16 585
R48 VTAIL.n19 VTAIL.n18 585
R49 VTAIL.n33 VTAIL.n32 585
R50 VTAIL.n35 VTAIL.n34 585
R51 VTAIL.n28 VTAIL.n27 585
R52 VTAIL.n41 VTAIL.n40 585
R53 VTAIL.n43 VTAIL.n42 585
R54 VTAIL.n57 VTAIL.n56 585
R55 VTAIL.n59 VTAIL.n58 585
R56 VTAIL.n52 VTAIL.n51 585
R57 VTAIL.n65 VTAIL.n64 585
R58 VTAIL.n67 VTAIL.n66 585
R59 VTAIL.n163 VTAIL.n162 585
R60 VTAIL.n161 VTAIL.n160 585
R61 VTAIL.n148 VTAIL.n147 585
R62 VTAIL.n155 VTAIL.n154 585
R63 VTAIL.n153 VTAIL.n152 585
R64 VTAIL.n139 VTAIL.n138 585
R65 VTAIL.n137 VTAIL.n136 585
R66 VTAIL.n124 VTAIL.n123 585
R67 VTAIL.n131 VTAIL.n130 585
R68 VTAIL.n129 VTAIL.n128 585
R69 VTAIL.n115 VTAIL.n114 585
R70 VTAIL.n113 VTAIL.n112 585
R71 VTAIL.n100 VTAIL.n99 585
R72 VTAIL.n107 VTAIL.n106 585
R73 VTAIL.n105 VTAIL.n104 585
R74 VTAIL.n91 VTAIL.n90 585
R75 VTAIL.n89 VTAIL.n88 585
R76 VTAIL.n76 VTAIL.n75 585
R77 VTAIL.n83 VTAIL.n82 585
R78 VTAIL.n81 VTAIL.n80 585
R79 VTAIL.n175 VTAIL.t1 328.587
R80 VTAIL.n7 VTAIL.t3 328.587
R81 VTAIL.n31 VTAIL.t6 328.587
R82 VTAIL.n55 VTAIL.t5 328.587
R83 VTAIL.n151 VTAIL.t4 328.587
R84 VTAIL.n127 VTAIL.t7 328.587
R85 VTAIL.n103 VTAIL.t0 328.587
R86 VTAIL.n79 VTAIL.t2 328.587
R87 VTAIL.n178 VTAIL.n177 171.744
R88 VTAIL.n178 VTAIL.n171 171.744
R89 VTAIL.n185 VTAIL.n171 171.744
R90 VTAIL.n186 VTAIL.n185 171.744
R91 VTAIL.n10 VTAIL.n9 171.744
R92 VTAIL.n10 VTAIL.n3 171.744
R93 VTAIL.n17 VTAIL.n3 171.744
R94 VTAIL.n18 VTAIL.n17 171.744
R95 VTAIL.n34 VTAIL.n33 171.744
R96 VTAIL.n34 VTAIL.n27 171.744
R97 VTAIL.n41 VTAIL.n27 171.744
R98 VTAIL.n42 VTAIL.n41 171.744
R99 VTAIL.n58 VTAIL.n57 171.744
R100 VTAIL.n58 VTAIL.n51 171.744
R101 VTAIL.n65 VTAIL.n51 171.744
R102 VTAIL.n66 VTAIL.n65 171.744
R103 VTAIL.n162 VTAIL.n161 171.744
R104 VTAIL.n161 VTAIL.n147 171.744
R105 VTAIL.n154 VTAIL.n147 171.744
R106 VTAIL.n154 VTAIL.n153 171.744
R107 VTAIL.n138 VTAIL.n137 171.744
R108 VTAIL.n137 VTAIL.n123 171.744
R109 VTAIL.n130 VTAIL.n123 171.744
R110 VTAIL.n130 VTAIL.n129 171.744
R111 VTAIL.n114 VTAIL.n113 171.744
R112 VTAIL.n113 VTAIL.n99 171.744
R113 VTAIL.n106 VTAIL.n99 171.744
R114 VTAIL.n106 VTAIL.n105 171.744
R115 VTAIL.n90 VTAIL.n89 171.744
R116 VTAIL.n89 VTAIL.n75 171.744
R117 VTAIL.n82 VTAIL.n75 171.744
R118 VTAIL.n82 VTAIL.n81 171.744
R119 VTAIL.n177 VTAIL.t1 85.8723
R120 VTAIL.n9 VTAIL.t3 85.8723
R121 VTAIL.n33 VTAIL.t6 85.8723
R122 VTAIL.n57 VTAIL.t5 85.8723
R123 VTAIL.n153 VTAIL.t4 85.8723
R124 VTAIL.n129 VTAIL.t7 85.8723
R125 VTAIL.n105 VTAIL.t0 85.8723
R126 VTAIL.n81 VTAIL.t2 85.8723
R127 VTAIL.n191 VTAIL.n190 31.0217
R128 VTAIL.n23 VTAIL.n22 31.0217
R129 VTAIL.n47 VTAIL.n46 31.0217
R130 VTAIL.n71 VTAIL.n70 31.0217
R131 VTAIL.n167 VTAIL.n166 31.0217
R132 VTAIL.n143 VTAIL.n142 31.0217
R133 VTAIL.n119 VTAIL.n118 31.0217
R134 VTAIL.n95 VTAIL.n94 31.0217
R135 VTAIL.n95 VTAIL.n71 18.0134
R136 VTAIL.n191 VTAIL.n167 18.0134
R137 VTAIL.n176 VTAIL.n175 16.3651
R138 VTAIL.n8 VTAIL.n7 16.3651
R139 VTAIL.n32 VTAIL.n31 16.3651
R140 VTAIL.n56 VTAIL.n55 16.3651
R141 VTAIL.n152 VTAIL.n151 16.3651
R142 VTAIL.n128 VTAIL.n127 16.3651
R143 VTAIL.n104 VTAIL.n103 16.3651
R144 VTAIL.n80 VTAIL.n79 16.3651
R145 VTAIL.n179 VTAIL.n174 12.8005
R146 VTAIL.n11 VTAIL.n6 12.8005
R147 VTAIL.n35 VTAIL.n30 12.8005
R148 VTAIL.n59 VTAIL.n54 12.8005
R149 VTAIL.n155 VTAIL.n150 12.8005
R150 VTAIL.n131 VTAIL.n126 12.8005
R151 VTAIL.n107 VTAIL.n102 12.8005
R152 VTAIL.n83 VTAIL.n78 12.8005
R153 VTAIL.n180 VTAIL.n172 12.0247
R154 VTAIL.n12 VTAIL.n4 12.0247
R155 VTAIL.n36 VTAIL.n28 12.0247
R156 VTAIL.n60 VTAIL.n52 12.0247
R157 VTAIL.n156 VTAIL.n148 12.0247
R158 VTAIL.n132 VTAIL.n124 12.0247
R159 VTAIL.n108 VTAIL.n100 12.0247
R160 VTAIL.n84 VTAIL.n76 12.0247
R161 VTAIL.n184 VTAIL.n183 11.249
R162 VTAIL.n16 VTAIL.n15 11.249
R163 VTAIL.n40 VTAIL.n39 11.249
R164 VTAIL.n64 VTAIL.n63 11.249
R165 VTAIL.n160 VTAIL.n159 11.249
R166 VTAIL.n136 VTAIL.n135 11.249
R167 VTAIL.n112 VTAIL.n111 11.249
R168 VTAIL.n88 VTAIL.n87 11.249
R169 VTAIL.n187 VTAIL.n170 10.4732
R170 VTAIL.n19 VTAIL.n2 10.4732
R171 VTAIL.n43 VTAIL.n26 10.4732
R172 VTAIL.n67 VTAIL.n50 10.4732
R173 VTAIL.n163 VTAIL.n146 10.4732
R174 VTAIL.n139 VTAIL.n122 10.4732
R175 VTAIL.n115 VTAIL.n98 10.4732
R176 VTAIL.n91 VTAIL.n74 10.4732
R177 VTAIL.n188 VTAIL.n168 9.69747
R178 VTAIL.n20 VTAIL.n0 9.69747
R179 VTAIL.n44 VTAIL.n24 9.69747
R180 VTAIL.n68 VTAIL.n48 9.69747
R181 VTAIL.n164 VTAIL.n144 9.69747
R182 VTAIL.n140 VTAIL.n120 9.69747
R183 VTAIL.n116 VTAIL.n96 9.69747
R184 VTAIL.n92 VTAIL.n72 9.69747
R185 VTAIL.n190 VTAIL.n189 9.45567
R186 VTAIL.n22 VTAIL.n21 9.45567
R187 VTAIL.n46 VTAIL.n45 9.45567
R188 VTAIL.n70 VTAIL.n69 9.45567
R189 VTAIL.n166 VTAIL.n165 9.45567
R190 VTAIL.n142 VTAIL.n141 9.45567
R191 VTAIL.n118 VTAIL.n117 9.45567
R192 VTAIL.n94 VTAIL.n93 9.45567
R193 VTAIL.n189 VTAIL.n188 9.3005
R194 VTAIL.n170 VTAIL.n169 9.3005
R195 VTAIL.n183 VTAIL.n182 9.3005
R196 VTAIL.n181 VTAIL.n180 9.3005
R197 VTAIL.n174 VTAIL.n173 9.3005
R198 VTAIL.n21 VTAIL.n20 9.3005
R199 VTAIL.n2 VTAIL.n1 9.3005
R200 VTAIL.n15 VTAIL.n14 9.3005
R201 VTAIL.n13 VTAIL.n12 9.3005
R202 VTAIL.n6 VTAIL.n5 9.3005
R203 VTAIL.n45 VTAIL.n44 9.3005
R204 VTAIL.n26 VTAIL.n25 9.3005
R205 VTAIL.n39 VTAIL.n38 9.3005
R206 VTAIL.n37 VTAIL.n36 9.3005
R207 VTAIL.n30 VTAIL.n29 9.3005
R208 VTAIL.n69 VTAIL.n68 9.3005
R209 VTAIL.n50 VTAIL.n49 9.3005
R210 VTAIL.n63 VTAIL.n62 9.3005
R211 VTAIL.n61 VTAIL.n60 9.3005
R212 VTAIL.n54 VTAIL.n53 9.3005
R213 VTAIL.n165 VTAIL.n164 9.3005
R214 VTAIL.n146 VTAIL.n145 9.3005
R215 VTAIL.n159 VTAIL.n158 9.3005
R216 VTAIL.n157 VTAIL.n156 9.3005
R217 VTAIL.n150 VTAIL.n149 9.3005
R218 VTAIL.n141 VTAIL.n140 9.3005
R219 VTAIL.n122 VTAIL.n121 9.3005
R220 VTAIL.n135 VTAIL.n134 9.3005
R221 VTAIL.n133 VTAIL.n132 9.3005
R222 VTAIL.n126 VTAIL.n125 9.3005
R223 VTAIL.n117 VTAIL.n116 9.3005
R224 VTAIL.n98 VTAIL.n97 9.3005
R225 VTAIL.n111 VTAIL.n110 9.3005
R226 VTAIL.n109 VTAIL.n108 9.3005
R227 VTAIL.n102 VTAIL.n101 9.3005
R228 VTAIL.n93 VTAIL.n92 9.3005
R229 VTAIL.n74 VTAIL.n73 9.3005
R230 VTAIL.n87 VTAIL.n86 9.3005
R231 VTAIL.n85 VTAIL.n84 9.3005
R232 VTAIL.n78 VTAIL.n77 9.3005
R233 VTAIL.n190 VTAIL.n168 4.26717
R234 VTAIL.n22 VTAIL.n0 4.26717
R235 VTAIL.n46 VTAIL.n24 4.26717
R236 VTAIL.n70 VTAIL.n48 4.26717
R237 VTAIL.n166 VTAIL.n144 4.26717
R238 VTAIL.n142 VTAIL.n120 4.26717
R239 VTAIL.n118 VTAIL.n96 4.26717
R240 VTAIL.n94 VTAIL.n72 4.26717
R241 VTAIL.n175 VTAIL.n173 3.73474
R242 VTAIL.n7 VTAIL.n5 3.73474
R243 VTAIL.n31 VTAIL.n29 3.73474
R244 VTAIL.n55 VTAIL.n53 3.73474
R245 VTAIL.n151 VTAIL.n149 3.73474
R246 VTAIL.n127 VTAIL.n125 3.73474
R247 VTAIL.n103 VTAIL.n101 3.73474
R248 VTAIL.n79 VTAIL.n77 3.73474
R249 VTAIL.n188 VTAIL.n187 3.49141
R250 VTAIL.n20 VTAIL.n19 3.49141
R251 VTAIL.n44 VTAIL.n43 3.49141
R252 VTAIL.n68 VTAIL.n67 3.49141
R253 VTAIL.n164 VTAIL.n163 3.49141
R254 VTAIL.n140 VTAIL.n139 3.49141
R255 VTAIL.n116 VTAIL.n115 3.49141
R256 VTAIL.n92 VTAIL.n91 3.49141
R257 VTAIL.n184 VTAIL.n170 2.71565
R258 VTAIL.n16 VTAIL.n2 2.71565
R259 VTAIL.n40 VTAIL.n26 2.71565
R260 VTAIL.n64 VTAIL.n50 2.71565
R261 VTAIL.n160 VTAIL.n146 2.71565
R262 VTAIL.n136 VTAIL.n122 2.71565
R263 VTAIL.n112 VTAIL.n98 2.71565
R264 VTAIL.n88 VTAIL.n74 2.71565
R265 VTAIL.n183 VTAIL.n172 1.93989
R266 VTAIL.n15 VTAIL.n4 1.93989
R267 VTAIL.n39 VTAIL.n28 1.93989
R268 VTAIL.n63 VTAIL.n52 1.93989
R269 VTAIL.n159 VTAIL.n148 1.93989
R270 VTAIL.n135 VTAIL.n124 1.93989
R271 VTAIL.n111 VTAIL.n100 1.93989
R272 VTAIL.n87 VTAIL.n76 1.93989
R273 VTAIL.n119 VTAIL.n95 1.76774
R274 VTAIL.n167 VTAIL.n143 1.76774
R275 VTAIL.n71 VTAIL.n47 1.76774
R276 VTAIL.n180 VTAIL.n179 1.16414
R277 VTAIL.n12 VTAIL.n11 1.16414
R278 VTAIL.n36 VTAIL.n35 1.16414
R279 VTAIL.n60 VTAIL.n59 1.16414
R280 VTAIL.n156 VTAIL.n155 1.16414
R281 VTAIL.n132 VTAIL.n131 1.16414
R282 VTAIL.n108 VTAIL.n107 1.16414
R283 VTAIL.n84 VTAIL.n83 1.16414
R284 VTAIL VTAIL.n23 0.94231
R285 VTAIL VTAIL.n191 0.825931
R286 VTAIL.n143 VTAIL.n119 0.470328
R287 VTAIL.n47 VTAIL.n23 0.470328
R288 VTAIL.n176 VTAIL.n174 0.388379
R289 VTAIL.n8 VTAIL.n6 0.388379
R290 VTAIL.n32 VTAIL.n30 0.388379
R291 VTAIL.n56 VTAIL.n54 0.388379
R292 VTAIL.n152 VTAIL.n150 0.388379
R293 VTAIL.n128 VTAIL.n126 0.388379
R294 VTAIL.n104 VTAIL.n102 0.388379
R295 VTAIL.n80 VTAIL.n78 0.388379
R296 VTAIL.n181 VTAIL.n173 0.155672
R297 VTAIL.n182 VTAIL.n181 0.155672
R298 VTAIL.n182 VTAIL.n169 0.155672
R299 VTAIL.n189 VTAIL.n169 0.155672
R300 VTAIL.n13 VTAIL.n5 0.155672
R301 VTAIL.n14 VTAIL.n13 0.155672
R302 VTAIL.n14 VTAIL.n1 0.155672
R303 VTAIL.n21 VTAIL.n1 0.155672
R304 VTAIL.n37 VTAIL.n29 0.155672
R305 VTAIL.n38 VTAIL.n37 0.155672
R306 VTAIL.n38 VTAIL.n25 0.155672
R307 VTAIL.n45 VTAIL.n25 0.155672
R308 VTAIL.n61 VTAIL.n53 0.155672
R309 VTAIL.n62 VTAIL.n61 0.155672
R310 VTAIL.n62 VTAIL.n49 0.155672
R311 VTAIL.n69 VTAIL.n49 0.155672
R312 VTAIL.n165 VTAIL.n145 0.155672
R313 VTAIL.n158 VTAIL.n145 0.155672
R314 VTAIL.n158 VTAIL.n157 0.155672
R315 VTAIL.n157 VTAIL.n149 0.155672
R316 VTAIL.n141 VTAIL.n121 0.155672
R317 VTAIL.n134 VTAIL.n121 0.155672
R318 VTAIL.n134 VTAIL.n133 0.155672
R319 VTAIL.n133 VTAIL.n125 0.155672
R320 VTAIL.n117 VTAIL.n97 0.155672
R321 VTAIL.n110 VTAIL.n97 0.155672
R322 VTAIL.n110 VTAIL.n109 0.155672
R323 VTAIL.n109 VTAIL.n101 0.155672
R324 VTAIL.n93 VTAIL.n73 0.155672
R325 VTAIL.n86 VTAIL.n73 0.155672
R326 VTAIL.n86 VTAIL.n85 0.155672
R327 VTAIL.n85 VTAIL.n77 0.155672
R328 VN.n0 VN.t0 98.4663
R329 VN.n1 VN.t1 98.4663
R330 VN.n0 VN.t2 98.0424
R331 VN.n1 VN.t3 98.0424
R332 VN VN.n1 47.6565
R333 VN VN.n0 9.49365
R334 VDD2.n2 VDD2.n0 135.811
R335 VDD2.n2 VDD2.n1 102.916
R336 VDD2.n1 VDD2.t0 7.22383
R337 VDD2.n1 VDD2.t2 7.22383
R338 VDD2.n0 VDD2.t3 7.22383
R339 VDD2.n0 VDD2.t1 7.22383
R340 VDD2 VDD2.n2 0.0586897
R341 B.n304 B.n43 585
R342 B.n306 B.n305 585
R343 B.n307 B.n42 585
R344 B.n309 B.n308 585
R345 B.n310 B.n41 585
R346 B.n312 B.n311 585
R347 B.n313 B.n40 585
R348 B.n315 B.n314 585
R349 B.n316 B.n39 585
R350 B.n318 B.n317 585
R351 B.n319 B.n38 585
R352 B.n321 B.n320 585
R353 B.n322 B.n37 585
R354 B.n324 B.n323 585
R355 B.n325 B.n36 585
R356 B.n327 B.n326 585
R357 B.n328 B.n35 585
R358 B.n330 B.n329 585
R359 B.n331 B.n34 585
R360 B.n333 B.n332 585
R361 B.n335 B.n31 585
R362 B.n337 B.n336 585
R363 B.n338 B.n30 585
R364 B.n340 B.n339 585
R365 B.n341 B.n29 585
R366 B.n343 B.n342 585
R367 B.n344 B.n28 585
R368 B.n346 B.n345 585
R369 B.n347 B.n25 585
R370 B.n350 B.n349 585
R371 B.n351 B.n24 585
R372 B.n353 B.n352 585
R373 B.n354 B.n23 585
R374 B.n356 B.n355 585
R375 B.n357 B.n22 585
R376 B.n359 B.n358 585
R377 B.n360 B.n21 585
R378 B.n362 B.n361 585
R379 B.n363 B.n20 585
R380 B.n365 B.n364 585
R381 B.n366 B.n19 585
R382 B.n368 B.n367 585
R383 B.n369 B.n18 585
R384 B.n371 B.n370 585
R385 B.n372 B.n17 585
R386 B.n374 B.n373 585
R387 B.n375 B.n16 585
R388 B.n377 B.n376 585
R389 B.n378 B.n15 585
R390 B.n303 B.n302 585
R391 B.n301 B.n44 585
R392 B.n300 B.n299 585
R393 B.n298 B.n45 585
R394 B.n297 B.n296 585
R395 B.n295 B.n46 585
R396 B.n294 B.n293 585
R397 B.n292 B.n47 585
R398 B.n291 B.n290 585
R399 B.n289 B.n48 585
R400 B.n288 B.n287 585
R401 B.n286 B.n49 585
R402 B.n285 B.n284 585
R403 B.n283 B.n50 585
R404 B.n282 B.n281 585
R405 B.n280 B.n51 585
R406 B.n279 B.n278 585
R407 B.n277 B.n52 585
R408 B.n276 B.n275 585
R409 B.n274 B.n53 585
R410 B.n273 B.n272 585
R411 B.n271 B.n54 585
R412 B.n270 B.n269 585
R413 B.n268 B.n55 585
R414 B.n267 B.n266 585
R415 B.n265 B.n56 585
R416 B.n264 B.n263 585
R417 B.n262 B.n57 585
R418 B.n261 B.n260 585
R419 B.n259 B.n58 585
R420 B.n258 B.n257 585
R421 B.n256 B.n59 585
R422 B.n255 B.n254 585
R423 B.n253 B.n60 585
R424 B.n252 B.n251 585
R425 B.n250 B.n61 585
R426 B.n249 B.n248 585
R427 B.n247 B.n62 585
R428 B.n246 B.n245 585
R429 B.n244 B.n63 585
R430 B.n243 B.n242 585
R431 B.n241 B.n64 585
R432 B.n240 B.n239 585
R433 B.n238 B.n65 585
R434 B.n237 B.n236 585
R435 B.n235 B.n66 585
R436 B.n234 B.n233 585
R437 B.n232 B.n67 585
R438 B.n231 B.n230 585
R439 B.n229 B.n68 585
R440 B.n228 B.n227 585
R441 B.n226 B.n69 585
R442 B.n225 B.n224 585
R443 B.n150 B.n149 585
R444 B.n151 B.n98 585
R445 B.n153 B.n152 585
R446 B.n154 B.n97 585
R447 B.n156 B.n155 585
R448 B.n157 B.n96 585
R449 B.n159 B.n158 585
R450 B.n160 B.n95 585
R451 B.n162 B.n161 585
R452 B.n163 B.n94 585
R453 B.n165 B.n164 585
R454 B.n166 B.n93 585
R455 B.n168 B.n167 585
R456 B.n169 B.n92 585
R457 B.n171 B.n170 585
R458 B.n172 B.n91 585
R459 B.n174 B.n173 585
R460 B.n175 B.n90 585
R461 B.n177 B.n176 585
R462 B.n178 B.n87 585
R463 B.n181 B.n180 585
R464 B.n182 B.n86 585
R465 B.n184 B.n183 585
R466 B.n185 B.n85 585
R467 B.n187 B.n186 585
R468 B.n188 B.n84 585
R469 B.n190 B.n189 585
R470 B.n191 B.n83 585
R471 B.n193 B.n192 585
R472 B.n195 B.n194 585
R473 B.n196 B.n79 585
R474 B.n198 B.n197 585
R475 B.n199 B.n78 585
R476 B.n201 B.n200 585
R477 B.n202 B.n77 585
R478 B.n204 B.n203 585
R479 B.n205 B.n76 585
R480 B.n207 B.n206 585
R481 B.n208 B.n75 585
R482 B.n210 B.n209 585
R483 B.n211 B.n74 585
R484 B.n213 B.n212 585
R485 B.n214 B.n73 585
R486 B.n216 B.n215 585
R487 B.n217 B.n72 585
R488 B.n219 B.n218 585
R489 B.n220 B.n71 585
R490 B.n222 B.n221 585
R491 B.n223 B.n70 585
R492 B.n148 B.n99 585
R493 B.n147 B.n146 585
R494 B.n145 B.n100 585
R495 B.n144 B.n143 585
R496 B.n142 B.n101 585
R497 B.n141 B.n140 585
R498 B.n139 B.n102 585
R499 B.n138 B.n137 585
R500 B.n136 B.n103 585
R501 B.n135 B.n134 585
R502 B.n133 B.n104 585
R503 B.n132 B.n131 585
R504 B.n130 B.n105 585
R505 B.n129 B.n128 585
R506 B.n127 B.n106 585
R507 B.n126 B.n125 585
R508 B.n124 B.n107 585
R509 B.n123 B.n122 585
R510 B.n121 B.n108 585
R511 B.n120 B.n119 585
R512 B.n118 B.n109 585
R513 B.n117 B.n116 585
R514 B.n115 B.n110 585
R515 B.n114 B.n113 585
R516 B.n112 B.n111 585
R517 B.n2 B.n0 585
R518 B.n417 B.n1 585
R519 B.n416 B.n415 585
R520 B.n414 B.n3 585
R521 B.n413 B.n412 585
R522 B.n411 B.n4 585
R523 B.n410 B.n409 585
R524 B.n408 B.n5 585
R525 B.n407 B.n406 585
R526 B.n405 B.n6 585
R527 B.n404 B.n403 585
R528 B.n402 B.n7 585
R529 B.n401 B.n400 585
R530 B.n399 B.n8 585
R531 B.n398 B.n397 585
R532 B.n396 B.n9 585
R533 B.n395 B.n394 585
R534 B.n393 B.n10 585
R535 B.n392 B.n391 585
R536 B.n390 B.n11 585
R537 B.n389 B.n388 585
R538 B.n387 B.n12 585
R539 B.n386 B.n385 585
R540 B.n384 B.n13 585
R541 B.n383 B.n382 585
R542 B.n381 B.n14 585
R543 B.n380 B.n379 585
R544 B.n419 B.n418 585
R545 B.n150 B.n99 506.916
R546 B.n380 B.n15 506.916
R547 B.n224 B.n223 506.916
R548 B.n302 B.n43 506.916
R549 B.n80 B.t5 282.163
R550 B.n32 B.t7 282.163
R551 B.n88 B.t11 282.163
R552 B.n26 B.t1 282.163
R553 B.n80 B.t3 269.228
R554 B.n88 B.t9 269.228
R555 B.n26 B.t0 269.228
R556 B.n32 B.t6 269.228
R557 B.n81 B.t4 242.405
R558 B.n33 B.t8 242.405
R559 B.n89 B.t10 242.405
R560 B.n27 B.t2 242.405
R561 B.n146 B.n99 163.367
R562 B.n146 B.n145 163.367
R563 B.n145 B.n144 163.367
R564 B.n144 B.n101 163.367
R565 B.n140 B.n101 163.367
R566 B.n140 B.n139 163.367
R567 B.n139 B.n138 163.367
R568 B.n138 B.n103 163.367
R569 B.n134 B.n103 163.367
R570 B.n134 B.n133 163.367
R571 B.n133 B.n132 163.367
R572 B.n132 B.n105 163.367
R573 B.n128 B.n105 163.367
R574 B.n128 B.n127 163.367
R575 B.n127 B.n126 163.367
R576 B.n126 B.n107 163.367
R577 B.n122 B.n107 163.367
R578 B.n122 B.n121 163.367
R579 B.n121 B.n120 163.367
R580 B.n120 B.n109 163.367
R581 B.n116 B.n109 163.367
R582 B.n116 B.n115 163.367
R583 B.n115 B.n114 163.367
R584 B.n114 B.n111 163.367
R585 B.n111 B.n2 163.367
R586 B.n418 B.n2 163.367
R587 B.n418 B.n417 163.367
R588 B.n417 B.n416 163.367
R589 B.n416 B.n3 163.367
R590 B.n412 B.n3 163.367
R591 B.n412 B.n411 163.367
R592 B.n411 B.n410 163.367
R593 B.n410 B.n5 163.367
R594 B.n406 B.n5 163.367
R595 B.n406 B.n405 163.367
R596 B.n405 B.n404 163.367
R597 B.n404 B.n7 163.367
R598 B.n400 B.n7 163.367
R599 B.n400 B.n399 163.367
R600 B.n399 B.n398 163.367
R601 B.n398 B.n9 163.367
R602 B.n394 B.n9 163.367
R603 B.n394 B.n393 163.367
R604 B.n393 B.n392 163.367
R605 B.n392 B.n11 163.367
R606 B.n388 B.n11 163.367
R607 B.n388 B.n387 163.367
R608 B.n387 B.n386 163.367
R609 B.n386 B.n13 163.367
R610 B.n382 B.n13 163.367
R611 B.n382 B.n381 163.367
R612 B.n381 B.n380 163.367
R613 B.n151 B.n150 163.367
R614 B.n152 B.n151 163.367
R615 B.n152 B.n97 163.367
R616 B.n156 B.n97 163.367
R617 B.n157 B.n156 163.367
R618 B.n158 B.n157 163.367
R619 B.n158 B.n95 163.367
R620 B.n162 B.n95 163.367
R621 B.n163 B.n162 163.367
R622 B.n164 B.n163 163.367
R623 B.n164 B.n93 163.367
R624 B.n168 B.n93 163.367
R625 B.n169 B.n168 163.367
R626 B.n170 B.n169 163.367
R627 B.n170 B.n91 163.367
R628 B.n174 B.n91 163.367
R629 B.n175 B.n174 163.367
R630 B.n176 B.n175 163.367
R631 B.n176 B.n87 163.367
R632 B.n181 B.n87 163.367
R633 B.n182 B.n181 163.367
R634 B.n183 B.n182 163.367
R635 B.n183 B.n85 163.367
R636 B.n187 B.n85 163.367
R637 B.n188 B.n187 163.367
R638 B.n189 B.n188 163.367
R639 B.n189 B.n83 163.367
R640 B.n193 B.n83 163.367
R641 B.n194 B.n193 163.367
R642 B.n194 B.n79 163.367
R643 B.n198 B.n79 163.367
R644 B.n199 B.n198 163.367
R645 B.n200 B.n199 163.367
R646 B.n200 B.n77 163.367
R647 B.n204 B.n77 163.367
R648 B.n205 B.n204 163.367
R649 B.n206 B.n205 163.367
R650 B.n206 B.n75 163.367
R651 B.n210 B.n75 163.367
R652 B.n211 B.n210 163.367
R653 B.n212 B.n211 163.367
R654 B.n212 B.n73 163.367
R655 B.n216 B.n73 163.367
R656 B.n217 B.n216 163.367
R657 B.n218 B.n217 163.367
R658 B.n218 B.n71 163.367
R659 B.n222 B.n71 163.367
R660 B.n223 B.n222 163.367
R661 B.n224 B.n69 163.367
R662 B.n228 B.n69 163.367
R663 B.n229 B.n228 163.367
R664 B.n230 B.n229 163.367
R665 B.n230 B.n67 163.367
R666 B.n234 B.n67 163.367
R667 B.n235 B.n234 163.367
R668 B.n236 B.n235 163.367
R669 B.n236 B.n65 163.367
R670 B.n240 B.n65 163.367
R671 B.n241 B.n240 163.367
R672 B.n242 B.n241 163.367
R673 B.n242 B.n63 163.367
R674 B.n246 B.n63 163.367
R675 B.n247 B.n246 163.367
R676 B.n248 B.n247 163.367
R677 B.n248 B.n61 163.367
R678 B.n252 B.n61 163.367
R679 B.n253 B.n252 163.367
R680 B.n254 B.n253 163.367
R681 B.n254 B.n59 163.367
R682 B.n258 B.n59 163.367
R683 B.n259 B.n258 163.367
R684 B.n260 B.n259 163.367
R685 B.n260 B.n57 163.367
R686 B.n264 B.n57 163.367
R687 B.n265 B.n264 163.367
R688 B.n266 B.n265 163.367
R689 B.n266 B.n55 163.367
R690 B.n270 B.n55 163.367
R691 B.n271 B.n270 163.367
R692 B.n272 B.n271 163.367
R693 B.n272 B.n53 163.367
R694 B.n276 B.n53 163.367
R695 B.n277 B.n276 163.367
R696 B.n278 B.n277 163.367
R697 B.n278 B.n51 163.367
R698 B.n282 B.n51 163.367
R699 B.n283 B.n282 163.367
R700 B.n284 B.n283 163.367
R701 B.n284 B.n49 163.367
R702 B.n288 B.n49 163.367
R703 B.n289 B.n288 163.367
R704 B.n290 B.n289 163.367
R705 B.n290 B.n47 163.367
R706 B.n294 B.n47 163.367
R707 B.n295 B.n294 163.367
R708 B.n296 B.n295 163.367
R709 B.n296 B.n45 163.367
R710 B.n300 B.n45 163.367
R711 B.n301 B.n300 163.367
R712 B.n302 B.n301 163.367
R713 B.n376 B.n15 163.367
R714 B.n376 B.n375 163.367
R715 B.n375 B.n374 163.367
R716 B.n374 B.n17 163.367
R717 B.n370 B.n17 163.367
R718 B.n370 B.n369 163.367
R719 B.n369 B.n368 163.367
R720 B.n368 B.n19 163.367
R721 B.n364 B.n19 163.367
R722 B.n364 B.n363 163.367
R723 B.n363 B.n362 163.367
R724 B.n362 B.n21 163.367
R725 B.n358 B.n21 163.367
R726 B.n358 B.n357 163.367
R727 B.n357 B.n356 163.367
R728 B.n356 B.n23 163.367
R729 B.n352 B.n23 163.367
R730 B.n352 B.n351 163.367
R731 B.n351 B.n350 163.367
R732 B.n350 B.n25 163.367
R733 B.n345 B.n25 163.367
R734 B.n345 B.n344 163.367
R735 B.n344 B.n343 163.367
R736 B.n343 B.n29 163.367
R737 B.n339 B.n29 163.367
R738 B.n339 B.n338 163.367
R739 B.n338 B.n337 163.367
R740 B.n337 B.n31 163.367
R741 B.n332 B.n31 163.367
R742 B.n332 B.n331 163.367
R743 B.n331 B.n330 163.367
R744 B.n330 B.n35 163.367
R745 B.n326 B.n35 163.367
R746 B.n326 B.n325 163.367
R747 B.n325 B.n324 163.367
R748 B.n324 B.n37 163.367
R749 B.n320 B.n37 163.367
R750 B.n320 B.n319 163.367
R751 B.n319 B.n318 163.367
R752 B.n318 B.n39 163.367
R753 B.n314 B.n39 163.367
R754 B.n314 B.n313 163.367
R755 B.n313 B.n312 163.367
R756 B.n312 B.n41 163.367
R757 B.n308 B.n41 163.367
R758 B.n308 B.n307 163.367
R759 B.n307 B.n306 163.367
R760 B.n306 B.n43 163.367
R761 B.n82 B.n81 59.5399
R762 B.n179 B.n89 59.5399
R763 B.n348 B.n27 59.5399
R764 B.n334 B.n33 59.5399
R765 B.n81 B.n80 39.7581
R766 B.n89 B.n88 39.7581
R767 B.n27 B.n26 39.7581
R768 B.n33 B.n32 39.7581
R769 B.n379 B.n378 32.9371
R770 B.n304 B.n303 32.9371
R771 B.n225 B.n70 32.9371
R772 B.n149 B.n148 32.9371
R773 B B.n419 18.0485
R774 B.n378 B.n377 10.6151
R775 B.n377 B.n16 10.6151
R776 B.n373 B.n16 10.6151
R777 B.n373 B.n372 10.6151
R778 B.n372 B.n371 10.6151
R779 B.n371 B.n18 10.6151
R780 B.n367 B.n18 10.6151
R781 B.n367 B.n366 10.6151
R782 B.n366 B.n365 10.6151
R783 B.n365 B.n20 10.6151
R784 B.n361 B.n20 10.6151
R785 B.n361 B.n360 10.6151
R786 B.n360 B.n359 10.6151
R787 B.n359 B.n22 10.6151
R788 B.n355 B.n22 10.6151
R789 B.n355 B.n354 10.6151
R790 B.n354 B.n353 10.6151
R791 B.n353 B.n24 10.6151
R792 B.n349 B.n24 10.6151
R793 B.n347 B.n346 10.6151
R794 B.n346 B.n28 10.6151
R795 B.n342 B.n28 10.6151
R796 B.n342 B.n341 10.6151
R797 B.n341 B.n340 10.6151
R798 B.n340 B.n30 10.6151
R799 B.n336 B.n30 10.6151
R800 B.n336 B.n335 10.6151
R801 B.n333 B.n34 10.6151
R802 B.n329 B.n34 10.6151
R803 B.n329 B.n328 10.6151
R804 B.n328 B.n327 10.6151
R805 B.n327 B.n36 10.6151
R806 B.n323 B.n36 10.6151
R807 B.n323 B.n322 10.6151
R808 B.n322 B.n321 10.6151
R809 B.n321 B.n38 10.6151
R810 B.n317 B.n38 10.6151
R811 B.n317 B.n316 10.6151
R812 B.n316 B.n315 10.6151
R813 B.n315 B.n40 10.6151
R814 B.n311 B.n40 10.6151
R815 B.n311 B.n310 10.6151
R816 B.n310 B.n309 10.6151
R817 B.n309 B.n42 10.6151
R818 B.n305 B.n42 10.6151
R819 B.n305 B.n304 10.6151
R820 B.n226 B.n225 10.6151
R821 B.n227 B.n226 10.6151
R822 B.n227 B.n68 10.6151
R823 B.n231 B.n68 10.6151
R824 B.n232 B.n231 10.6151
R825 B.n233 B.n232 10.6151
R826 B.n233 B.n66 10.6151
R827 B.n237 B.n66 10.6151
R828 B.n238 B.n237 10.6151
R829 B.n239 B.n238 10.6151
R830 B.n239 B.n64 10.6151
R831 B.n243 B.n64 10.6151
R832 B.n244 B.n243 10.6151
R833 B.n245 B.n244 10.6151
R834 B.n245 B.n62 10.6151
R835 B.n249 B.n62 10.6151
R836 B.n250 B.n249 10.6151
R837 B.n251 B.n250 10.6151
R838 B.n251 B.n60 10.6151
R839 B.n255 B.n60 10.6151
R840 B.n256 B.n255 10.6151
R841 B.n257 B.n256 10.6151
R842 B.n257 B.n58 10.6151
R843 B.n261 B.n58 10.6151
R844 B.n262 B.n261 10.6151
R845 B.n263 B.n262 10.6151
R846 B.n263 B.n56 10.6151
R847 B.n267 B.n56 10.6151
R848 B.n268 B.n267 10.6151
R849 B.n269 B.n268 10.6151
R850 B.n269 B.n54 10.6151
R851 B.n273 B.n54 10.6151
R852 B.n274 B.n273 10.6151
R853 B.n275 B.n274 10.6151
R854 B.n275 B.n52 10.6151
R855 B.n279 B.n52 10.6151
R856 B.n280 B.n279 10.6151
R857 B.n281 B.n280 10.6151
R858 B.n281 B.n50 10.6151
R859 B.n285 B.n50 10.6151
R860 B.n286 B.n285 10.6151
R861 B.n287 B.n286 10.6151
R862 B.n287 B.n48 10.6151
R863 B.n291 B.n48 10.6151
R864 B.n292 B.n291 10.6151
R865 B.n293 B.n292 10.6151
R866 B.n293 B.n46 10.6151
R867 B.n297 B.n46 10.6151
R868 B.n298 B.n297 10.6151
R869 B.n299 B.n298 10.6151
R870 B.n299 B.n44 10.6151
R871 B.n303 B.n44 10.6151
R872 B.n149 B.n98 10.6151
R873 B.n153 B.n98 10.6151
R874 B.n154 B.n153 10.6151
R875 B.n155 B.n154 10.6151
R876 B.n155 B.n96 10.6151
R877 B.n159 B.n96 10.6151
R878 B.n160 B.n159 10.6151
R879 B.n161 B.n160 10.6151
R880 B.n161 B.n94 10.6151
R881 B.n165 B.n94 10.6151
R882 B.n166 B.n165 10.6151
R883 B.n167 B.n166 10.6151
R884 B.n167 B.n92 10.6151
R885 B.n171 B.n92 10.6151
R886 B.n172 B.n171 10.6151
R887 B.n173 B.n172 10.6151
R888 B.n173 B.n90 10.6151
R889 B.n177 B.n90 10.6151
R890 B.n178 B.n177 10.6151
R891 B.n180 B.n86 10.6151
R892 B.n184 B.n86 10.6151
R893 B.n185 B.n184 10.6151
R894 B.n186 B.n185 10.6151
R895 B.n186 B.n84 10.6151
R896 B.n190 B.n84 10.6151
R897 B.n191 B.n190 10.6151
R898 B.n192 B.n191 10.6151
R899 B.n196 B.n195 10.6151
R900 B.n197 B.n196 10.6151
R901 B.n197 B.n78 10.6151
R902 B.n201 B.n78 10.6151
R903 B.n202 B.n201 10.6151
R904 B.n203 B.n202 10.6151
R905 B.n203 B.n76 10.6151
R906 B.n207 B.n76 10.6151
R907 B.n208 B.n207 10.6151
R908 B.n209 B.n208 10.6151
R909 B.n209 B.n74 10.6151
R910 B.n213 B.n74 10.6151
R911 B.n214 B.n213 10.6151
R912 B.n215 B.n214 10.6151
R913 B.n215 B.n72 10.6151
R914 B.n219 B.n72 10.6151
R915 B.n220 B.n219 10.6151
R916 B.n221 B.n220 10.6151
R917 B.n221 B.n70 10.6151
R918 B.n148 B.n147 10.6151
R919 B.n147 B.n100 10.6151
R920 B.n143 B.n100 10.6151
R921 B.n143 B.n142 10.6151
R922 B.n142 B.n141 10.6151
R923 B.n141 B.n102 10.6151
R924 B.n137 B.n102 10.6151
R925 B.n137 B.n136 10.6151
R926 B.n136 B.n135 10.6151
R927 B.n135 B.n104 10.6151
R928 B.n131 B.n104 10.6151
R929 B.n131 B.n130 10.6151
R930 B.n130 B.n129 10.6151
R931 B.n129 B.n106 10.6151
R932 B.n125 B.n106 10.6151
R933 B.n125 B.n124 10.6151
R934 B.n124 B.n123 10.6151
R935 B.n123 B.n108 10.6151
R936 B.n119 B.n108 10.6151
R937 B.n119 B.n118 10.6151
R938 B.n118 B.n117 10.6151
R939 B.n117 B.n110 10.6151
R940 B.n113 B.n110 10.6151
R941 B.n113 B.n112 10.6151
R942 B.n112 B.n0 10.6151
R943 B.n415 B.n1 10.6151
R944 B.n415 B.n414 10.6151
R945 B.n414 B.n413 10.6151
R946 B.n413 B.n4 10.6151
R947 B.n409 B.n4 10.6151
R948 B.n409 B.n408 10.6151
R949 B.n408 B.n407 10.6151
R950 B.n407 B.n6 10.6151
R951 B.n403 B.n6 10.6151
R952 B.n403 B.n402 10.6151
R953 B.n402 B.n401 10.6151
R954 B.n401 B.n8 10.6151
R955 B.n397 B.n8 10.6151
R956 B.n397 B.n396 10.6151
R957 B.n396 B.n395 10.6151
R958 B.n395 B.n10 10.6151
R959 B.n391 B.n10 10.6151
R960 B.n391 B.n390 10.6151
R961 B.n390 B.n389 10.6151
R962 B.n389 B.n12 10.6151
R963 B.n385 B.n12 10.6151
R964 B.n385 B.n384 10.6151
R965 B.n384 B.n383 10.6151
R966 B.n383 B.n14 10.6151
R967 B.n379 B.n14 10.6151
R968 B.n348 B.n347 6.5566
R969 B.n335 B.n334 6.5566
R970 B.n180 B.n179 6.5566
R971 B.n192 B.n82 6.5566
R972 B.n349 B.n348 4.05904
R973 B.n334 B.n333 4.05904
R974 B.n179 B.n178 4.05904
R975 B.n195 B.n82 4.05904
R976 B.n419 B.n0 2.81026
R977 B.n419 B.n1 2.81026
C0 VDD1 VTAIL 3.31702f
C1 VN VP 4.172f
C2 B VDD1 0.904917f
C3 w_n2200_n1868# VDD2 1.11128f
C4 VDD2 VTAIL 3.36533f
C5 B VDD2 0.94278f
C6 VP VDD1 2.01656f
C7 VN VDD1 0.152357f
C8 VP VDD2 0.342812f
C9 VN VDD2 1.82699f
C10 w_n2200_n1868# VTAIL 2.21656f
C11 B w_n2200_n1868# 6.06705f
C12 B VTAIL 2.17628f
C13 VDD2 VDD1 0.811921f
C14 VP w_n2200_n1868# 3.70431f
C15 VN w_n2200_n1868# 3.42396f
C16 VP VTAIL 2.03161f
C17 VN VTAIL 2.0175f
C18 B VP 1.32151f
C19 VN B 0.860082f
C20 w_n2200_n1868# VDD1 1.07517f
C21 VDD2 VSUBS 0.567941f
C22 VDD1 VSUBS 4.154968f
C23 VTAIL VSUBS 0.558122f
C24 VN VSUBS 4.48017f
C25 VP VSUBS 1.393223f
C26 B VSUBS 2.740467f
C27 w_n2200_n1868# VSUBS 51.612f
C28 B.n0 VSUBS 0.005945f
C29 B.n1 VSUBS 0.005945f
C30 B.n2 VSUBS 0.009401f
C31 B.n3 VSUBS 0.009401f
C32 B.n4 VSUBS 0.009401f
C33 B.n5 VSUBS 0.009401f
C34 B.n6 VSUBS 0.009401f
C35 B.n7 VSUBS 0.009401f
C36 B.n8 VSUBS 0.009401f
C37 B.n9 VSUBS 0.009401f
C38 B.n10 VSUBS 0.009401f
C39 B.n11 VSUBS 0.009401f
C40 B.n12 VSUBS 0.009401f
C41 B.n13 VSUBS 0.009401f
C42 B.n14 VSUBS 0.009401f
C43 B.n15 VSUBS 0.022967f
C44 B.n16 VSUBS 0.009401f
C45 B.n17 VSUBS 0.009401f
C46 B.n18 VSUBS 0.009401f
C47 B.n19 VSUBS 0.009401f
C48 B.n20 VSUBS 0.009401f
C49 B.n21 VSUBS 0.009401f
C50 B.n22 VSUBS 0.009401f
C51 B.n23 VSUBS 0.009401f
C52 B.n24 VSUBS 0.009401f
C53 B.n25 VSUBS 0.009401f
C54 B.t2 VSUBS 0.086965f
C55 B.t1 VSUBS 0.108409f
C56 B.t0 VSUBS 0.488424f
C57 B.n26 VSUBS 0.194481f
C58 B.n27 VSUBS 0.165599f
C59 B.n28 VSUBS 0.009401f
C60 B.n29 VSUBS 0.009401f
C61 B.n30 VSUBS 0.009401f
C62 B.n31 VSUBS 0.009401f
C63 B.t8 VSUBS 0.086967f
C64 B.t7 VSUBS 0.108411f
C65 B.t6 VSUBS 0.488424f
C66 B.n32 VSUBS 0.19448f
C67 B.n33 VSUBS 0.165597f
C68 B.n34 VSUBS 0.009401f
C69 B.n35 VSUBS 0.009401f
C70 B.n36 VSUBS 0.009401f
C71 B.n37 VSUBS 0.009401f
C72 B.n38 VSUBS 0.009401f
C73 B.n39 VSUBS 0.009401f
C74 B.n40 VSUBS 0.009401f
C75 B.n41 VSUBS 0.009401f
C76 B.n42 VSUBS 0.009401f
C77 B.n43 VSUBS 0.022967f
C78 B.n44 VSUBS 0.009401f
C79 B.n45 VSUBS 0.009401f
C80 B.n46 VSUBS 0.009401f
C81 B.n47 VSUBS 0.009401f
C82 B.n48 VSUBS 0.009401f
C83 B.n49 VSUBS 0.009401f
C84 B.n50 VSUBS 0.009401f
C85 B.n51 VSUBS 0.009401f
C86 B.n52 VSUBS 0.009401f
C87 B.n53 VSUBS 0.009401f
C88 B.n54 VSUBS 0.009401f
C89 B.n55 VSUBS 0.009401f
C90 B.n56 VSUBS 0.009401f
C91 B.n57 VSUBS 0.009401f
C92 B.n58 VSUBS 0.009401f
C93 B.n59 VSUBS 0.009401f
C94 B.n60 VSUBS 0.009401f
C95 B.n61 VSUBS 0.009401f
C96 B.n62 VSUBS 0.009401f
C97 B.n63 VSUBS 0.009401f
C98 B.n64 VSUBS 0.009401f
C99 B.n65 VSUBS 0.009401f
C100 B.n66 VSUBS 0.009401f
C101 B.n67 VSUBS 0.009401f
C102 B.n68 VSUBS 0.009401f
C103 B.n69 VSUBS 0.009401f
C104 B.n70 VSUBS 0.022967f
C105 B.n71 VSUBS 0.009401f
C106 B.n72 VSUBS 0.009401f
C107 B.n73 VSUBS 0.009401f
C108 B.n74 VSUBS 0.009401f
C109 B.n75 VSUBS 0.009401f
C110 B.n76 VSUBS 0.009401f
C111 B.n77 VSUBS 0.009401f
C112 B.n78 VSUBS 0.009401f
C113 B.n79 VSUBS 0.009401f
C114 B.t4 VSUBS 0.086967f
C115 B.t5 VSUBS 0.108411f
C116 B.t3 VSUBS 0.488424f
C117 B.n80 VSUBS 0.19448f
C118 B.n81 VSUBS 0.165597f
C119 B.n82 VSUBS 0.021782f
C120 B.n83 VSUBS 0.009401f
C121 B.n84 VSUBS 0.009401f
C122 B.n85 VSUBS 0.009401f
C123 B.n86 VSUBS 0.009401f
C124 B.n87 VSUBS 0.009401f
C125 B.t10 VSUBS 0.086965f
C126 B.t11 VSUBS 0.108409f
C127 B.t9 VSUBS 0.488424f
C128 B.n88 VSUBS 0.194481f
C129 B.n89 VSUBS 0.165599f
C130 B.n90 VSUBS 0.009401f
C131 B.n91 VSUBS 0.009401f
C132 B.n92 VSUBS 0.009401f
C133 B.n93 VSUBS 0.009401f
C134 B.n94 VSUBS 0.009401f
C135 B.n95 VSUBS 0.009401f
C136 B.n96 VSUBS 0.009401f
C137 B.n97 VSUBS 0.009401f
C138 B.n98 VSUBS 0.009401f
C139 B.n99 VSUBS 0.021275f
C140 B.n100 VSUBS 0.009401f
C141 B.n101 VSUBS 0.009401f
C142 B.n102 VSUBS 0.009401f
C143 B.n103 VSUBS 0.009401f
C144 B.n104 VSUBS 0.009401f
C145 B.n105 VSUBS 0.009401f
C146 B.n106 VSUBS 0.009401f
C147 B.n107 VSUBS 0.009401f
C148 B.n108 VSUBS 0.009401f
C149 B.n109 VSUBS 0.009401f
C150 B.n110 VSUBS 0.009401f
C151 B.n111 VSUBS 0.009401f
C152 B.n112 VSUBS 0.009401f
C153 B.n113 VSUBS 0.009401f
C154 B.n114 VSUBS 0.009401f
C155 B.n115 VSUBS 0.009401f
C156 B.n116 VSUBS 0.009401f
C157 B.n117 VSUBS 0.009401f
C158 B.n118 VSUBS 0.009401f
C159 B.n119 VSUBS 0.009401f
C160 B.n120 VSUBS 0.009401f
C161 B.n121 VSUBS 0.009401f
C162 B.n122 VSUBS 0.009401f
C163 B.n123 VSUBS 0.009401f
C164 B.n124 VSUBS 0.009401f
C165 B.n125 VSUBS 0.009401f
C166 B.n126 VSUBS 0.009401f
C167 B.n127 VSUBS 0.009401f
C168 B.n128 VSUBS 0.009401f
C169 B.n129 VSUBS 0.009401f
C170 B.n130 VSUBS 0.009401f
C171 B.n131 VSUBS 0.009401f
C172 B.n132 VSUBS 0.009401f
C173 B.n133 VSUBS 0.009401f
C174 B.n134 VSUBS 0.009401f
C175 B.n135 VSUBS 0.009401f
C176 B.n136 VSUBS 0.009401f
C177 B.n137 VSUBS 0.009401f
C178 B.n138 VSUBS 0.009401f
C179 B.n139 VSUBS 0.009401f
C180 B.n140 VSUBS 0.009401f
C181 B.n141 VSUBS 0.009401f
C182 B.n142 VSUBS 0.009401f
C183 B.n143 VSUBS 0.009401f
C184 B.n144 VSUBS 0.009401f
C185 B.n145 VSUBS 0.009401f
C186 B.n146 VSUBS 0.009401f
C187 B.n147 VSUBS 0.009401f
C188 B.n148 VSUBS 0.021275f
C189 B.n149 VSUBS 0.022967f
C190 B.n150 VSUBS 0.022967f
C191 B.n151 VSUBS 0.009401f
C192 B.n152 VSUBS 0.009401f
C193 B.n153 VSUBS 0.009401f
C194 B.n154 VSUBS 0.009401f
C195 B.n155 VSUBS 0.009401f
C196 B.n156 VSUBS 0.009401f
C197 B.n157 VSUBS 0.009401f
C198 B.n158 VSUBS 0.009401f
C199 B.n159 VSUBS 0.009401f
C200 B.n160 VSUBS 0.009401f
C201 B.n161 VSUBS 0.009401f
C202 B.n162 VSUBS 0.009401f
C203 B.n163 VSUBS 0.009401f
C204 B.n164 VSUBS 0.009401f
C205 B.n165 VSUBS 0.009401f
C206 B.n166 VSUBS 0.009401f
C207 B.n167 VSUBS 0.009401f
C208 B.n168 VSUBS 0.009401f
C209 B.n169 VSUBS 0.009401f
C210 B.n170 VSUBS 0.009401f
C211 B.n171 VSUBS 0.009401f
C212 B.n172 VSUBS 0.009401f
C213 B.n173 VSUBS 0.009401f
C214 B.n174 VSUBS 0.009401f
C215 B.n175 VSUBS 0.009401f
C216 B.n176 VSUBS 0.009401f
C217 B.n177 VSUBS 0.009401f
C218 B.n178 VSUBS 0.006498f
C219 B.n179 VSUBS 0.021782f
C220 B.n180 VSUBS 0.007604f
C221 B.n181 VSUBS 0.009401f
C222 B.n182 VSUBS 0.009401f
C223 B.n183 VSUBS 0.009401f
C224 B.n184 VSUBS 0.009401f
C225 B.n185 VSUBS 0.009401f
C226 B.n186 VSUBS 0.009401f
C227 B.n187 VSUBS 0.009401f
C228 B.n188 VSUBS 0.009401f
C229 B.n189 VSUBS 0.009401f
C230 B.n190 VSUBS 0.009401f
C231 B.n191 VSUBS 0.009401f
C232 B.n192 VSUBS 0.007604f
C233 B.n193 VSUBS 0.009401f
C234 B.n194 VSUBS 0.009401f
C235 B.n195 VSUBS 0.006498f
C236 B.n196 VSUBS 0.009401f
C237 B.n197 VSUBS 0.009401f
C238 B.n198 VSUBS 0.009401f
C239 B.n199 VSUBS 0.009401f
C240 B.n200 VSUBS 0.009401f
C241 B.n201 VSUBS 0.009401f
C242 B.n202 VSUBS 0.009401f
C243 B.n203 VSUBS 0.009401f
C244 B.n204 VSUBS 0.009401f
C245 B.n205 VSUBS 0.009401f
C246 B.n206 VSUBS 0.009401f
C247 B.n207 VSUBS 0.009401f
C248 B.n208 VSUBS 0.009401f
C249 B.n209 VSUBS 0.009401f
C250 B.n210 VSUBS 0.009401f
C251 B.n211 VSUBS 0.009401f
C252 B.n212 VSUBS 0.009401f
C253 B.n213 VSUBS 0.009401f
C254 B.n214 VSUBS 0.009401f
C255 B.n215 VSUBS 0.009401f
C256 B.n216 VSUBS 0.009401f
C257 B.n217 VSUBS 0.009401f
C258 B.n218 VSUBS 0.009401f
C259 B.n219 VSUBS 0.009401f
C260 B.n220 VSUBS 0.009401f
C261 B.n221 VSUBS 0.009401f
C262 B.n222 VSUBS 0.009401f
C263 B.n223 VSUBS 0.022967f
C264 B.n224 VSUBS 0.021275f
C265 B.n225 VSUBS 0.021275f
C266 B.n226 VSUBS 0.009401f
C267 B.n227 VSUBS 0.009401f
C268 B.n228 VSUBS 0.009401f
C269 B.n229 VSUBS 0.009401f
C270 B.n230 VSUBS 0.009401f
C271 B.n231 VSUBS 0.009401f
C272 B.n232 VSUBS 0.009401f
C273 B.n233 VSUBS 0.009401f
C274 B.n234 VSUBS 0.009401f
C275 B.n235 VSUBS 0.009401f
C276 B.n236 VSUBS 0.009401f
C277 B.n237 VSUBS 0.009401f
C278 B.n238 VSUBS 0.009401f
C279 B.n239 VSUBS 0.009401f
C280 B.n240 VSUBS 0.009401f
C281 B.n241 VSUBS 0.009401f
C282 B.n242 VSUBS 0.009401f
C283 B.n243 VSUBS 0.009401f
C284 B.n244 VSUBS 0.009401f
C285 B.n245 VSUBS 0.009401f
C286 B.n246 VSUBS 0.009401f
C287 B.n247 VSUBS 0.009401f
C288 B.n248 VSUBS 0.009401f
C289 B.n249 VSUBS 0.009401f
C290 B.n250 VSUBS 0.009401f
C291 B.n251 VSUBS 0.009401f
C292 B.n252 VSUBS 0.009401f
C293 B.n253 VSUBS 0.009401f
C294 B.n254 VSUBS 0.009401f
C295 B.n255 VSUBS 0.009401f
C296 B.n256 VSUBS 0.009401f
C297 B.n257 VSUBS 0.009401f
C298 B.n258 VSUBS 0.009401f
C299 B.n259 VSUBS 0.009401f
C300 B.n260 VSUBS 0.009401f
C301 B.n261 VSUBS 0.009401f
C302 B.n262 VSUBS 0.009401f
C303 B.n263 VSUBS 0.009401f
C304 B.n264 VSUBS 0.009401f
C305 B.n265 VSUBS 0.009401f
C306 B.n266 VSUBS 0.009401f
C307 B.n267 VSUBS 0.009401f
C308 B.n268 VSUBS 0.009401f
C309 B.n269 VSUBS 0.009401f
C310 B.n270 VSUBS 0.009401f
C311 B.n271 VSUBS 0.009401f
C312 B.n272 VSUBS 0.009401f
C313 B.n273 VSUBS 0.009401f
C314 B.n274 VSUBS 0.009401f
C315 B.n275 VSUBS 0.009401f
C316 B.n276 VSUBS 0.009401f
C317 B.n277 VSUBS 0.009401f
C318 B.n278 VSUBS 0.009401f
C319 B.n279 VSUBS 0.009401f
C320 B.n280 VSUBS 0.009401f
C321 B.n281 VSUBS 0.009401f
C322 B.n282 VSUBS 0.009401f
C323 B.n283 VSUBS 0.009401f
C324 B.n284 VSUBS 0.009401f
C325 B.n285 VSUBS 0.009401f
C326 B.n286 VSUBS 0.009401f
C327 B.n287 VSUBS 0.009401f
C328 B.n288 VSUBS 0.009401f
C329 B.n289 VSUBS 0.009401f
C330 B.n290 VSUBS 0.009401f
C331 B.n291 VSUBS 0.009401f
C332 B.n292 VSUBS 0.009401f
C333 B.n293 VSUBS 0.009401f
C334 B.n294 VSUBS 0.009401f
C335 B.n295 VSUBS 0.009401f
C336 B.n296 VSUBS 0.009401f
C337 B.n297 VSUBS 0.009401f
C338 B.n298 VSUBS 0.009401f
C339 B.n299 VSUBS 0.009401f
C340 B.n300 VSUBS 0.009401f
C341 B.n301 VSUBS 0.009401f
C342 B.n302 VSUBS 0.021275f
C343 B.n303 VSUBS 0.022376f
C344 B.n304 VSUBS 0.021866f
C345 B.n305 VSUBS 0.009401f
C346 B.n306 VSUBS 0.009401f
C347 B.n307 VSUBS 0.009401f
C348 B.n308 VSUBS 0.009401f
C349 B.n309 VSUBS 0.009401f
C350 B.n310 VSUBS 0.009401f
C351 B.n311 VSUBS 0.009401f
C352 B.n312 VSUBS 0.009401f
C353 B.n313 VSUBS 0.009401f
C354 B.n314 VSUBS 0.009401f
C355 B.n315 VSUBS 0.009401f
C356 B.n316 VSUBS 0.009401f
C357 B.n317 VSUBS 0.009401f
C358 B.n318 VSUBS 0.009401f
C359 B.n319 VSUBS 0.009401f
C360 B.n320 VSUBS 0.009401f
C361 B.n321 VSUBS 0.009401f
C362 B.n322 VSUBS 0.009401f
C363 B.n323 VSUBS 0.009401f
C364 B.n324 VSUBS 0.009401f
C365 B.n325 VSUBS 0.009401f
C366 B.n326 VSUBS 0.009401f
C367 B.n327 VSUBS 0.009401f
C368 B.n328 VSUBS 0.009401f
C369 B.n329 VSUBS 0.009401f
C370 B.n330 VSUBS 0.009401f
C371 B.n331 VSUBS 0.009401f
C372 B.n332 VSUBS 0.009401f
C373 B.n333 VSUBS 0.006498f
C374 B.n334 VSUBS 0.021782f
C375 B.n335 VSUBS 0.007604f
C376 B.n336 VSUBS 0.009401f
C377 B.n337 VSUBS 0.009401f
C378 B.n338 VSUBS 0.009401f
C379 B.n339 VSUBS 0.009401f
C380 B.n340 VSUBS 0.009401f
C381 B.n341 VSUBS 0.009401f
C382 B.n342 VSUBS 0.009401f
C383 B.n343 VSUBS 0.009401f
C384 B.n344 VSUBS 0.009401f
C385 B.n345 VSUBS 0.009401f
C386 B.n346 VSUBS 0.009401f
C387 B.n347 VSUBS 0.007604f
C388 B.n348 VSUBS 0.021782f
C389 B.n349 VSUBS 0.006498f
C390 B.n350 VSUBS 0.009401f
C391 B.n351 VSUBS 0.009401f
C392 B.n352 VSUBS 0.009401f
C393 B.n353 VSUBS 0.009401f
C394 B.n354 VSUBS 0.009401f
C395 B.n355 VSUBS 0.009401f
C396 B.n356 VSUBS 0.009401f
C397 B.n357 VSUBS 0.009401f
C398 B.n358 VSUBS 0.009401f
C399 B.n359 VSUBS 0.009401f
C400 B.n360 VSUBS 0.009401f
C401 B.n361 VSUBS 0.009401f
C402 B.n362 VSUBS 0.009401f
C403 B.n363 VSUBS 0.009401f
C404 B.n364 VSUBS 0.009401f
C405 B.n365 VSUBS 0.009401f
C406 B.n366 VSUBS 0.009401f
C407 B.n367 VSUBS 0.009401f
C408 B.n368 VSUBS 0.009401f
C409 B.n369 VSUBS 0.009401f
C410 B.n370 VSUBS 0.009401f
C411 B.n371 VSUBS 0.009401f
C412 B.n372 VSUBS 0.009401f
C413 B.n373 VSUBS 0.009401f
C414 B.n374 VSUBS 0.009401f
C415 B.n375 VSUBS 0.009401f
C416 B.n376 VSUBS 0.009401f
C417 B.n377 VSUBS 0.009401f
C418 B.n378 VSUBS 0.022967f
C419 B.n379 VSUBS 0.021275f
C420 B.n380 VSUBS 0.021275f
C421 B.n381 VSUBS 0.009401f
C422 B.n382 VSUBS 0.009401f
C423 B.n383 VSUBS 0.009401f
C424 B.n384 VSUBS 0.009401f
C425 B.n385 VSUBS 0.009401f
C426 B.n386 VSUBS 0.009401f
C427 B.n387 VSUBS 0.009401f
C428 B.n388 VSUBS 0.009401f
C429 B.n389 VSUBS 0.009401f
C430 B.n390 VSUBS 0.009401f
C431 B.n391 VSUBS 0.009401f
C432 B.n392 VSUBS 0.009401f
C433 B.n393 VSUBS 0.009401f
C434 B.n394 VSUBS 0.009401f
C435 B.n395 VSUBS 0.009401f
C436 B.n396 VSUBS 0.009401f
C437 B.n397 VSUBS 0.009401f
C438 B.n398 VSUBS 0.009401f
C439 B.n399 VSUBS 0.009401f
C440 B.n400 VSUBS 0.009401f
C441 B.n401 VSUBS 0.009401f
C442 B.n402 VSUBS 0.009401f
C443 B.n403 VSUBS 0.009401f
C444 B.n404 VSUBS 0.009401f
C445 B.n405 VSUBS 0.009401f
C446 B.n406 VSUBS 0.009401f
C447 B.n407 VSUBS 0.009401f
C448 B.n408 VSUBS 0.009401f
C449 B.n409 VSUBS 0.009401f
C450 B.n410 VSUBS 0.009401f
C451 B.n411 VSUBS 0.009401f
C452 B.n412 VSUBS 0.009401f
C453 B.n413 VSUBS 0.009401f
C454 B.n414 VSUBS 0.009401f
C455 B.n415 VSUBS 0.009401f
C456 B.n416 VSUBS 0.009401f
C457 B.n417 VSUBS 0.009401f
C458 B.n418 VSUBS 0.009401f
C459 B.n419 VSUBS 0.021288f
C460 VDD2.t3 VSUBS 0.063596f
C461 VDD2.t1 VSUBS 0.063596f
C462 VDD2.n0 VSUBS 0.596624f
C463 VDD2.t0 VSUBS 0.063596f
C464 VDD2.t2 VSUBS 0.063596f
C465 VDD2.n1 VSUBS 0.386013f
C466 VDD2.n2 VSUBS 2.05729f
C467 VN.t0 VSUBS 1.08126f
C468 VN.t2 VSUBS 1.07883f
C469 VN.n0 VSUBS 0.794276f
C470 VN.t1 VSUBS 1.08126f
C471 VN.t3 VSUBS 1.07883f
C472 VN.n1 VSUBS 2.2557f
C473 VTAIL.n0 VSUBS 0.029139f
C474 VTAIL.n1 VSUBS 0.028146f
C475 VTAIL.n2 VSUBS 0.015125f
C476 VTAIL.n3 VSUBS 0.035749f
C477 VTAIL.n4 VSUBS 0.016014f
C478 VTAIL.n5 VSUBS 0.452841f
C479 VTAIL.n6 VSUBS 0.015125f
C480 VTAIL.t3 VSUBS 0.077362f
C481 VTAIL.n7 VSUBS 0.11247f
C482 VTAIL.n8 VSUBS 0.022647f
C483 VTAIL.n9 VSUBS 0.026812f
C484 VTAIL.n10 VSUBS 0.035749f
C485 VTAIL.n11 VSUBS 0.016014f
C486 VTAIL.n12 VSUBS 0.015125f
C487 VTAIL.n13 VSUBS 0.028146f
C488 VTAIL.n14 VSUBS 0.028146f
C489 VTAIL.n15 VSUBS 0.015125f
C490 VTAIL.n16 VSUBS 0.016014f
C491 VTAIL.n17 VSUBS 0.035749f
C492 VTAIL.n18 VSUBS 0.080454f
C493 VTAIL.n19 VSUBS 0.016014f
C494 VTAIL.n20 VSUBS 0.015125f
C495 VTAIL.n21 VSUBS 0.062752f
C496 VTAIL.n22 VSUBS 0.040117f
C497 VTAIL.n23 VSUBS 0.150765f
C498 VTAIL.n24 VSUBS 0.029139f
C499 VTAIL.n25 VSUBS 0.028146f
C500 VTAIL.n26 VSUBS 0.015125f
C501 VTAIL.n27 VSUBS 0.035749f
C502 VTAIL.n28 VSUBS 0.016014f
C503 VTAIL.n29 VSUBS 0.452841f
C504 VTAIL.n30 VSUBS 0.015125f
C505 VTAIL.t6 VSUBS 0.077362f
C506 VTAIL.n31 VSUBS 0.11247f
C507 VTAIL.n32 VSUBS 0.022647f
C508 VTAIL.n33 VSUBS 0.026812f
C509 VTAIL.n34 VSUBS 0.035749f
C510 VTAIL.n35 VSUBS 0.016014f
C511 VTAIL.n36 VSUBS 0.015125f
C512 VTAIL.n37 VSUBS 0.028146f
C513 VTAIL.n38 VSUBS 0.028146f
C514 VTAIL.n39 VSUBS 0.015125f
C515 VTAIL.n40 VSUBS 0.016014f
C516 VTAIL.n41 VSUBS 0.035749f
C517 VTAIL.n42 VSUBS 0.080454f
C518 VTAIL.n43 VSUBS 0.016014f
C519 VTAIL.n44 VSUBS 0.015125f
C520 VTAIL.n45 VSUBS 0.062752f
C521 VTAIL.n46 VSUBS 0.040117f
C522 VTAIL.n47 VSUBS 0.225626f
C523 VTAIL.n48 VSUBS 0.029139f
C524 VTAIL.n49 VSUBS 0.028146f
C525 VTAIL.n50 VSUBS 0.015125f
C526 VTAIL.n51 VSUBS 0.035749f
C527 VTAIL.n52 VSUBS 0.016014f
C528 VTAIL.n53 VSUBS 0.452841f
C529 VTAIL.n54 VSUBS 0.015125f
C530 VTAIL.t5 VSUBS 0.077362f
C531 VTAIL.n55 VSUBS 0.11247f
C532 VTAIL.n56 VSUBS 0.022647f
C533 VTAIL.n57 VSUBS 0.026812f
C534 VTAIL.n58 VSUBS 0.035749f
C535 VTAIL.n59 VSUBS 0.016014f
C536 VTAIL.n60 VSUBS 0.015125f
C537 VTAIL.n61 VSUBS 0.028146f
C538 VTAIL.n62 VSUBS 0.028146f
C539 VTAIL.n63 VSUBS 0.015125f
C540 VTAIL.n64 VSUBS 0.016014f
C541 VTAIL.n65 VSUBS 0.035749f
C542 VTAIL.n66 VSUBS 0.080454f
C543 VTAIL.n67 VSUBS 0.016014f
C544 VTAIL.n68 VSUBS 0.015125f
C545 VTAIL.n69 VSUBS 0.062752f
C546 VTAIL.n70 VSUBS 0.040117f
C547 VTAIL.n71 VSUBS 1.07746f
C548 VTAIL.n72 VSUBS 0.029139f
C549 VTAIL.n73 VSUBS 0.028146f
C550 VTAIL.n74 VSUBS 0.015125f
C551 VTAIL.n75 VSUBS 0.035749f
C552 VTAIL.n76 VSUBS 0.016014f
C553 VTAIL.n77 VSUBS 0.452841f
C554 VTAIL.n78 VSUBS 0.015125f
C555 VTAIL.t2 VSUBS 0.077362f
C556 VTAIL.n79 VSUBS 0.11247f
C557 VTAIL.n80 VSUBS 0.022647f
C558 VTAIL.n81 VSUBS 0.026812f
C559 VTAIL.n82 VSUBS 0.035749f
C560 VTAIL.n83 VSUBS 0.016014f
C561 VTAIL.n84 VSUBS 0.015125f
C562 VTAIL.n85 VSUBS 0.028146f
C563 VTAIL.n86 VSUBS 0.028146f
C564 VTAIL.n87 VSUBS 0.015125f
C565 VTAIL.n88 VSUBS 0.016014f
C566 VTAIL.n89 VSUBS 0.035749f
C567 VTAIL.n90 VSUBS 0.080454f
C568 VTAIL.n91 VSUBS 0.016014f
C569 VTAIL.n92 VSUBS 0.015125f
C570 VTAIL.n93 VSUBS 0.062752f
C571 VTAIL.n94 VSUBS 0.040117f
C572 VTAIL.n95 VSUBS 1.07746f
C573 VTAIL.n96 VSUBS 0.029139f
C574 VTAIL.n97 VSUBS 0.028146f
C575 VTAIL.n98 VSUBS 0.015125f
C576 VTAIL.n99 VSUBS 0.035749f
C577 VTAIL.n100 VSUBS 0.016014f
C578 VTAIL.n101 VSUBS 0.452841f
C579 VTAIL.n102 VSUBS 0.015125f
C580 VTAIL.t0 VSUBS 0.077362f
C581 VTAIL.n103 VSUBS 0.11247f
C582 VTAIL.n104 VSUBS 0.022647f
C583 VTAIL.n105 VSUBS 0.026812f
C584 VTAIL.n106 VSUBS 0.035749f
C585 VTAIL.n107 VSUBS 0.016014f
C586 VTAIL.n108 VSUBS 0.015125f
C587 VTAIL.n109 VSUBS 0.028146f
C588 VTAIL.n110 VSUBS 0.028146f
C589 VTAIL.n111 VSUBS 0.015125f
C590 VTAIL.n112 VSUBS 0.016014f
C591 VTAIL.n113 VSUBS 0.035749f
C592 VTAIL.n114 VSUBS 0.080454f
C593 VTAIL.n115 VSUBS 0.016014f
C594 VTAIL.n116 VSUBS 0.015125f
C595 VTAIL.n117 VSUBS 0.062752f
C596 VTAIL.n118 VSUBS 0.040117f
C597 VTAIL.n119 VSUBS 0.225626f
C598 VTAIL.n120 VSUBS 0.029139f
C599 VTAIL.n121 VSUBS 0.028146f
C600 VTAIL.n122 VSUBS 0.015125f
C601 VTAIL.n123 VSUBS 0.035749f
C602 VTAIL.n124 VSUBS 0.016014f
C603 VTAIL.n125 VSUBS 0.452841f
C604 VTAIL.n126 VSUBS 0.015125f
C605 VTAIL.t7 VSUBS 0.077362f
C606 VTAIL.n127 VSUBS 0.11247f
C607 VTAIL.n128 VSUBS 0.022647f
C608 VTAIL.n129 VSUBS 0.026812f
C609 VTAIL.n130 VSUBS 0.035749f
C610 VTAIL.n131 VSUBS 0.016014f
C611 VTAIL.n132 VSUBS 0.015125f
C612 VTAIL.n133 VSUBS 0.028146f
C613 VTAIL.n134 VSUBS 0.028146f
C614 VTAIL.n135 VSUBS 0.015125f
C615 VTAIL.n136 VSUBS 0.016014f
C616 VTAIL.n137 VSUBS 0.035749f
C617 VTAIL.n138 VSUBS 0.080454f
C618 VTAIL.n139 VSUBS 0.016014f
C619 VTAIL.n140 VSUBS 0.015125f
C620 VTAIL.n141 VSUBS 0.062752f
C621 VTAIL.n142 VSUBS 0.040117f
C622 VTAIL.n143 VSUBS 0.225626f
C623 VTAIL.n144 VSUBS 0.029139f
C624 VTAIL.n145 VSUBS 0.028146f
C625 VTAIL.n146 VSUBS 0.015125f
C626 VTAIL.n147 VSUBS 0.035749f
C627 VTAIL.n148 VSUBS 0.016014f
C628 VTAIL.n149 VSUBS 0.452841f
C629 VTAIL.n150 VSUBS 0.015125f
C630 VTAIL.t4 VSUBS 0.077362f
C631 VTAIL.n151 VSUBS 0.11247f
C632 VTAIL.n152 VSUBS 0.022647f
C633 VTAIL.n153 VSUBS 0.026812f
C634 VTAIL.n154 VSUBS 0.035749f
C635 VTAIL.n155 VSUBS 0.016014f
C636 VTAIL.n156 VSUBS 0.015125f
C637 VTAIL.n157 VSUBS 0.028146f
C638 VTAIL.n158 VSUBS 0.028146f
C639 VTAIL.n159 VSUBS 0.015125f
C640 VTAIL.n160 VSUBS 0.016014f
C641 VTAIL.n161 VSUBS 0.035749f
C642 VTAIL.n162 VSUBS 0.080454f
C643 VTAIL.n163 VSUBS 0.016014f
C644 VTAIL.n164 VSUBS 0.015125f
C645 VTAIL.n165 VSUBS 0.062752f
C646 VTAIL.n166 VSUBS 0.040117f
C647 VTAIL.n167 VSUBS 1.07746f
C648 VTAIL.n168 VSUBS 0.029139f
C649 VTAIL.n169 VSUBS 0.028146f
C650 VTAIL.n170 VSUBS 0.015125f
C651 VTAIL.n171 VSUBS 0.035749f
C652 VTAIL.n172 VSUBS 0.016014f
C653 VTAIL.n173 VSUBS 0.452841f
C654 VTAIL.n174 VSUBS 0.015125f
C655 VTAIL.t1 VSUBS 0.077362f
C656 VTAIL.n175 VSUBS 0.11247f
C657 VTAIL.n176 VSUBS 0.022647f
C658 VTAIL.n177 VSUBS 0.026812f
C659 VTAIL.n178 VSUBS 0.035749f
C660 VTAIL.n179 VSUBS 0.016014f
C661 VTAIL.n180 VSUBS 0.015125f
C662 VTAIL.n181 VSUBS 0.028146f
C663 VTAIL.n182 VSUBS 0.028146f
C664 VTAIL.n183 VSUBS 0.015125f
C665 VTAIL.n184 VSUBS 0.016014f
C666 VTAIL.n185 VSUBS 0.035749f
C667 VTAIL.n186 VSUBS 0.080454f
C668 VTAIL.n187 VSUBS 0.016014f
C669 VTAIL.n188 VSUBS 0.015125f
C670 VTAIL.n189 VSUBS 0.062752f
C671 VTAIL.n190 VSUBS 0.040117f
C672 VTAIL.n191 VSUBS 0.99204f
C673 VDD1.t3 VSUBS 0.097245f
C674 VDD1.t2 VSUBS 0.097245f
C675 VDD1.n0 VSUBS 0.590585f
C676 VDD1.t0 VSUBS 0.097245f
C677 VDD1.t1 VSUBS 0.097245f
C678 VDD1.n1 VSUBS 0.929842f
C679 VP.n0 VSUBS 0.054644f
C680 VP.t1 VSUBS 1.09748f
C681 VP.n1 VSUBS 0.044134f
C682 VP.n2 VSUBS 0.054644f
C683 VP.t2 VSUBS 1.09748f
C684 VP.t0 VSUBS 1.34896f
C685 VP.t3 VSUBS 1.34593f
C686 VP.n3 VSUBS 2.78164f
C687 VP.n4 VSUBS 2.39775f
C688 VP.n5 VSUBS 0.555039f
C689 VP.n6 VSUBS 0.053808f
C690 VP.n7 VSUBS 0.108032f
C691 VP.n8 VSUBS 0.054644f
C692 VP.n9 VSUBS 0.054644f
C693 VP.n10 VSUBS 0.054644f
C694 VP.n11 VSUBS 0.108032f
C695 VP.n12 VSUBS 0.053808f
C696 VP.n13 VSUBS 0.555039f
C697 VP.n14 VSUBS 0.058268f
.ends

