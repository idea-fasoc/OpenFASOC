* NGSPICE file created from diff_pair_sample_0262.ext - technology: sky130A

.subckt diff_pair_sample_0262 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=3.939 ps=20.98 w=10.1 l=3.55
X1 VDD2.t5 VN.t0 VTAIL.t2 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=1.6665 ps=10.43 w=10.1 l=3.55
X2 B.t11 B.t9 B.t10 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=0 ps=0 w=10.1 l=3.55
X3 VTAIL.t11 VP.t1 VDD1.t4 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=1.6665 ps=10.43 w=10.1 l=3.55
X4 VTAIL.t10 VP.t2 VDD1.t3 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=1.6665 ps=10.43 w=10.1 l=3.55
X5 VDD2.t4 VN.t1 VTAIL.t3 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=3.939 ps=20.98 w=10.1 l=3.55
X6 VDD2.t3 VN.t2 VTAIL.t4 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=1.6665 ps=10.43 w=10.1 l=3.55
X7 VDD1.t2 VP.t3 VTAIL.t7 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=3.939 ps=20.98 w=10.1 l=3.55
X8 VDD2.t2 VN.t3 VTAIL.t1 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=3.939 ps=20.98 w=10.1 l=3.55
X9 VTAIL.t0 VN.t4 VDD2.t1 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=1.6665 ps=10.43 w=10.1 l=3.55
X10 VDD1.t1 VP.t4 VTAIL.t6 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=1.6665 ps=10.43 w=10.1 l=3.55
X11 B.t8 B.t6 B.t7 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=0 ps=0 w=10.1 l=3.55
X12 B.t5 B.t3 B.t4 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=0 ps=0 w=10.1 l=3.55
X13 VTAIL.t5 VN.t5 VDD2.t0 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=1.6665 pd=10.43 as=1.6665 ps=10.43 w=10.1 l=3.55
X14 B.t2 B.t0 B.t1 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=0 ps=0 w=10.1 l=3.55
X15 VDD1.t0 VP.t5 VTAIL.t9 w_n4074_n2988# sky130_fd_pr__pfet_01v8 ad=3.939 pd=20.98 as=1.6665 ps=10.43 w=10.1 l=3.55
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n55 VP.n54 161.3
R9 VP.n53 VP.n1 161.3
R10 VP.n52 VP.n51 161.3
R11 VP.n50 VP.n2 161.3
R12 VP.n49 VP.n48 161.3
R13 VP.n47 VP.n3 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n4 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n40 VP.n5 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n6 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n7 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n31 VP.n8 161.3
R24 VP.n15 VP.t5 101.382
R25 VP.n30 VP.n29 83.8517
R26 VP.n56 VP.n0 83.8517
R27 VP.n28 VP.n9 83.8517
R28 VP.n29 VP.t4 68.5667
R29 VP.n41 VP.t1 68.5667
R30 VP.n0 VP.t0 68.5667
R31 VP.n9 VP.t3 68.5667
R32 VP.n14 VP.t2 68.5667
R33 VP.n15 VP.n14 62.4228
R34 VP.n35 VP.n6 56.5617
R35 VP.n48 VP.n2 56.5617
R36 VP.n20 VP.n11 56.5617
R37 VP.n30 VP.n28 51.0071
R38 VP.n33 VP.n8 24.5923
R39 VP.n34 VP.n33 24.5923
R40 VP.n35 VP.n34 24.5923
R41 VP.n39 VP.n6 24.5923
R42 VP.n40 VP.n39 24.5923
R43 VP.n42 VP.n40 24.5923
R44 VP.n46 VP.n4 24.5923
R45 VP.n47 VP.n46 24.5923
R46 VP.n48 VP.n47 24.5923
R47 VP.n52 VP.n2 24.5923
R48 VP.n53 VP.n52 24.5923
R49 VP.n54 VP.n53 24.5923
R50 VP.n24 VP.n11 24.5923
R51 VP.n25 VP.n24 24.5923
R52 VP.n26 VP.n25 24.5923
R53 VP.n18 VP.n13 24.5923
R54 VP.n19 VP.n18 24.5923
R55 VP.n20 VP.n19 24.5923
R56 VP.n42 VP.n41 12.2964
R57 VP.n41 VP.n4 12.2964
R58 VP.n14 VP.n13 12.2964
R59 VP.n29 VP.n8 6.39438
R60 VP.n54 VP.n0 6.39438
R61 VP.n26 VP.n9 6.39438
R62 VP.n16 VP.n15 3.26267
R63 VP.n28 VP.n27 0.354861
R64 VP.n31 VP.n30 0.354861
R65 VP.n56 VP.n55 0.354861
R66 VP VP.n56 0.267071
R67 VP.n17 VP.n16 0.189894
R68 VP.n17 VP.n12 0.189894
R69 VP.n21 VP.n12 0.189894
R70 VP.n22 VP.n21 0.189894
R71 VP.n23 VP.n22 0.189894
R72 VP.n23 VP.n10 0.189894
R73 VP.n27 VP.n10 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n32 VP.n7 0.189894
R76 VP.n36 VP.n7 0.189894
R77 VP.n37 VP.n36 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n38 VP.n5 0.189894
R80 VP.n43 VP.n5 0.189894
R81 VP.n44 VP.n43 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n45 VP.n3 0.189894
R84 VP.n49 VP.n3 0.189894
R85 VP.n50 VP.n49 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n51 VP.n1 0.189894
R88 VP.n55 VP.n1 0.189894
R89 VTAIL.n218 VTAIL.n170 756.745
R90 VTAIL.n50 VTAIL.n2 756.745
R91 VTAIL.n164 VTAIL.n116 756.745
R92 VTAIL.n108 VTAIL.n60 756.745
R93 VTAIL.n186 VTAIL.n185 585
R94 VTAIL.n191 VTAIL.n190 585
R95 VTAIL.n193 VTAIL.n192 585
R96 VTAIL.n182 VTAIL.n181 585
R97 VTAIL.n199 VTAIL.n198 585
R98 VTAIL.n201 VTAIL.n200 585
R99 VTAIL.n178 VTAIL.n177 585
R100 VTAIL.n208 VTAIL.n207 585
R101 VTAIL.n209 VTAIL.n176 585
R102 VTAIL.n211 VTAIL.n210 585
R103 VTAIL.n174 VTAIL.n173 585
R104 VTAIL.n217 VTAIL.n216 585
R105 VTAIL.n219 VTAIL.n218 585
R106 VTAIL.n18 VTAIL.n17 585
R107 VTAIL.n23 VTAIL.n22 585
R108 VTAIL.n25 VTAIL.n24 585
R109 VTAIL.n14 VTAIL.n13 585
R110 VTAIL.n31 VTAIL.n30 585
R111 VTAIL.n33 VTAIL.n32 585
R112 VTAIL.n10 VTAIL.n9 585
R113 VTAIL.n40 VTAIL.n39 585
R114 VTAIL.n41 VTAIL.n8 585
R115 VTAIL.n43 VTAIL.n42 585
R116 VTAIL.n6 VTAIL.n5 585
R117 VTAIL.n49 VTAIL.n48 585
R118 VTAIL.n51 VTAIL.n50 585
R119 VTAIL.n165 VTAIL.n164 585
R120 VTAIL.n163 VTAIL.n162 585
R121 VTAIL.n120 VTAIL.n119 585
R122 VTAIL.n157 VTAIL.n156 585
R123 VTAIL.n155 VTAIL.n122 585
R124 VTAIL.n154 VTAIL.n153 585
R125 VTAIL.n125 VTAIL.n123 585
R126 VTAIL.n148 VTAIL.n147 585
R127 VTAIL.n146 VTAIL.n145 585
R128 VTAIL.n129 VTAIL.n128 585
R129 VTAIL.n140 VTAIL.n139 585
R130 VTAIL.n138 VTAIL.n137 585
R131 VTAIL.n133 VTAIL.n132 585
R132 VTAIL.n109 VTAIL.n108 585
R133 VTAIL.n107 VTAIL.n106 585
R134 VTAIL.n64 VTAIL.n63 585
R135 VTAIL.n101 VTAIL.n100 585
R136 VTAIL.n99 VTAIL.n66 585
R137 VTAIL.n98 VTAIL.n97 585
R138 VTAIL.n69 VTAIL.n67 585
R139 VTAIL.n92 VTAIL.n91 585
R140 VTAIL.n90 VTAIL.n89 585
R141 VTAIL.n73 VTAIL.n72 585
R142 VTAIL.n84 VTAIL.n83 585
R143 VTAIL.n82 VTAIL.n81 585
R144 VTAIL.n77 VTAIL.n76 585
R145 VTAIL.n187 VTAIL.t1 329.038
R146 VTAIL.n19 VTAIL.t8 329.038
R147 VTAIL.n134 VTAIL.t7 329.038
R148 VTAIL.n78 VTAIL.t3 329.038
R149 VTAIL.n191 VTAIL.n185 171.744
R150 VTAIL.n192 VTAIL.n191 171.744
R151 VTAIL.n192 VTAIL.n181 171.744
R152 VTAIL.n199 VTAIL.n181 171.744
R153 VTAIL.n200 VTAIL.n199 171.744
R154 VTAIL.n200 VTAIL.n177 171.744
R155 VTAIL.n208 VTAIL.n177 171.744
R156 VTAIL.n209 VTAIL.n208 171.744
R157 VTAIL.n210 VTAIL.n209 171.744
R158 VTAIL.n210 VTAIL.n173 171.744
R159 VTAIL.n217 VTAIL.n173 171.744
R160 VTAIL.n218 VTAIL.n217 171.744
R161 VTAIL.n23 VTAIL.n17 171.744
R162 VTAIL.n24 VTAIL.n23 171.744
R163 VTAIL.n24 VTAIL.n13 171.744
R164 VTAIL.n31 VTAIL.n13 171.744
R165 VTAIL.n32 VTAIL.n31 171.744
R166 VTAIL.n32 VTAIL.n9 171.744
R167 VTAIL.n40 VTAIL.n9 171.744
R168 VTAIL.n41 VTAIL.n40 171.744
R169 VTAIL.n42 VTAIL.n41 171.744
R170 VTAIL.n42 VTAIL.n5 171.744
R171 VTAIL.n49 VTAIL.n5 171.744
R172 VTAIL.n50 VTAIL.n49 171.744
R173 VTAIL.n164 VTAIL.n163 171.744
R174 VTAIL.n163 VTAIL.n119 171.744
R175 VTAIL.n156 VTAIL.n119 171.744
R176 VTAIL.n156 VTAIL.n155 171.744
R177 VTAIL.n155 VTAIL.n154 171.744
R178 VTAIL.n154 VTAIL.n123 171.744
R179 VTAIL.n147 VTAIL.n123 171.744
R180 VTAIL.n147 VTAIL.n146 171.744
R181 VTAIL.n146 VTAIL.n128 171.744
R182 VTAIL.n139 VTAIL.n128 171.744
R183 VTAIL.n139 VTAIL.n138 171.744
R184 VTAIL.n138 VTAIL.n132 171.744
R185 VTAIL.n108 VTAIL.n107 171.744
R186 VTAIL.n107 VTAIL.n63 171.744
R187 VTAIL.n100 VTAIL.n63 171.744
R188 VTAIL.n100 VTAIL.n99 171.744
R189 VTAIL.n99 VTAIL.n98 171.744
R190 VTAIL.n98 VTAIL.n67 171.744
R191 VTAIL.n91 VTAIL.n67 171.744
R192 VTAIL.n91 VTAIL.n90 171.744
R193 VTAIL.n90 VTAIL.n72 171.744
R194 VTAIL.n83 VTAIL.n72 171.744
R195 VTAIL.n83 VTAIL.n82 171.744
R196 VTAIL.n82 VTAIL.n76 171.744
R197 VTAIL.t1 VTAIL.n185 85.8723
R198 VTAIL.t8 VTAIL.n17 85.8723
R199 VTAIL.t7 VTAIL.n132 85.8723
R200 VTAIL.t3 VTAIL.n76 85.8723
R201 VTAIL.n115 VTAIL.n114 63.1553
R202 VTAIL.n59 VTAIL.n58 63.1553
R203 VTAIL.n1 VTAIL.n0 63.1551
R204 VTAIL.n57 VTAIL.n56 63.1551
R205 VTAIL.n223 VTAIL.n222 34.9005
R206 VTAIL.n55 VTAIL.n54 34.9005
R207 VTAIL.n169 VTAIL.n168 34.9005
R208 VTAIL.n113 VTAIL.n112 34.9005
R209 VTAIL.n59 VTAIL.n57 27.7634
R210 VTAIL.n223 VTAIL.n169 24.4186
R211 VTAIL.n211 VTAIL.n176 13.1884
R212 VTAIL.n43 VTAIL.n8 13.1884
R213 VTAIL.n157 VTAIL.n122 13.1884
R214 VTAIL.n101 VTAIL.n66 13.1884
R215 VTAIL.n207 VTAIL.n206 12.8005
R216 VTAIL.n212 VTAIL.n174 12.8005
R217 VTAIL.n39 VTAIL.n38 12.8005
R218 VTAIL.n44 VTAIL.n6 12.8005
R219 VTAIL.n158 VTAIL.n120 12.8005
R220 VTAIL.n153 VTAIL.n124 12.8005
R221 VTAIL.n102 VTAIL.n64 12.8005
R222 VTAIL.n97 VTAIL.n68 12.8005
R223 VTAIL.n205 VTAIL.n178 12.0247
R224 VTAIL.n216 VTAIL.n215 12.0247
R225 VTAIL.n37 VTAIL.n10 12.0247
R226 VTAIL.n48 VTAIL.n47 12.0247
R227 VTAIL.n162 VTAIL.n161 12.0247
R228 VTAIL.n152 VTAIL.n125 12.0247
R229 VTAIL.n106 VTAIL.n105 12.0247
R230 VTAIL.n96 VTAIL.n69 12.0247
R231 VTAIL.n202 VTAIL.n201 11.249
R232 VTAIL.n219 VTAIL.n172 11.249
R233 VTAIL.n34 VTAIL.n33 11.249
R234 VTAIL.n51 VTAIL.n4 11.249
R235 VTAIL.n165 VTAIL.n118 11.249
R236 VTAIL.n149 VTAIL.n148 11.249
R237 VTAIL.n109 VTAIL.n62 11.249
R238 VTAIL.n93 VTAIL.n92 11.249
R239 VTAIL.n187 VTAIL.n186 10.7239
R240 VTAIL.n19 VTAIL.n18 10.7239
R241 VTAIL.n134 VTAIL.n133 10.7239
R242 VTAIL.n78 VTAIL.n77 10.7239
R243 VTAIL.n198 VTAIL.n180 10.4732
R244 VTAIL.n220 VTAIL.n170 10.4732
R245 VTAIL.n30 VTAIL.n12 10.4732
R246 VTAIL.n52 VTAIL.n2 10.4732
R247 VTAIL.n166 VTAIL.n116 10.4732
R248 VTAIL.n145 VTAIL.n127 10.4732
R249 VTAIL.n110 VTAIL.n60 10.4732
R250 VTAIL.n89 VTAIL.n71 10.4732
R251 VTAIL.n197 VTAIL.n182 9.69747
R252 VTAIL.n29 VTAIL.n14 9.69747
R253 VTAIL.n144 VTAIL.n129 9.69747
R254 VTAIL.n88 VTAIL.n73 9.69747
R255 VTAIL.n222 VTAIL.n221 9.45567
R256 VTAIL.n54 VTAIL.n53 9.45567
R257 VTAIL.n168 VTAIL.n167 9.45567
R258 VTAIL.n112 VTAIL.n111 9.45567
R259 VTAIL.n221 VTAIL.n220 9.3005
R260 VTAIL.n172 VTAIL.n171 9.3005
R261 VTAIL.n215 VTAIL.n214 9.3005
R262 VTAIL.n213 VTAIL.n212 9.3005
R263 VTAIL.n189 VTAIL.n188 9.3005
R264 VTAIL.n184 VTAIL.n183 9.3005
R265 VTAIL.n195 VTAIL.n194 9.3005
R266 VTAIL.n197 VTAIL.n196 9.3005
R267 VTAIL.n180 VTAIL.n179 9.3005
R268 VTAIL.n203 VTAIL.n202 9.3005
R269 VTAIL.n205 VTAIL.n204 9.3005
R270 VTAIL.n206 VTAIL.n175 9.3005
R271 VTAIL.n53 VTAIL.n52 9.3005
R272 VTAIL.n4 VTAIL.n3 9.3005
R273 VTAIL.n47 VTAIL.n46 9.3005
R274 VTAIL.n45 VTAIL.n44 9.3005
R275 VTAIL.n21 VTAIL.n20 9.3005
R276 VTAIL.n16 VTAIL.n15 9.3005
R277 VTAIL.n27 VTAIL.n26 9.3005
R278 VTAIL.n29 VTAIL.n28 9.3005
R279 VTAIL.n12 VTAIL.n11 9.3005
R280 VTAIL.n35 VTAIL.n34 9.3005
R281 VTAIL.n37 VTAIL.n36 9.3005
R282 VTAIL.n38 VTAIL.n7 9.3005
R283 VTAIL.n136 VTAIL.n135 9.3005
R284 VTAIL.n131 VTAIL.n130 9.3005
R285 VTAIL.n142 VTAIL.n141 9.3005
R286 VTAIL.n144 VTAIL.n143 9.3005
R287 VTAIL.n127 VTAIL.n126 9.3005
R288 VTAIL.n150 VTAIL.n149 9.3005
R289 VTAIL.n152 VTAIL.n151 9.3005
R290 VTAIL.n124 VTAIL.n121 9.3005
R291 VTAIL.n167 VTAIL.n166 9.3005
R292 VTAIL.n118 VTAIL.n117 9.3005
R293 VTAIL.n161 VTAIL.n160 9.3005
R294 VTAIL.n159 VTAIL.n158 9.3005
R295 VTAIL.n80 VTAIL.n79 9.3005
R296 VTAIL.n75 VTAIL.n74 9.3005
R297 VTAIL.n86 VTAIL.n85 9.3005
R298 VTAIL.n88 VTAIL.n87 9.3005
R299 VTAIL.n71 VTAIL.n70 9.3005
R300 VTAIL.n94 VTAIL.n93 9.3005
R301 VTAIL.n96 VTAIL.n95 9.3005
R302 VTAIL.n68 VTAIL.n65 9.3005
R303 VTAIL.n111 VTAIL.n110 9.3005
R304 VTAIL.n62 VTAIL.n61 9.3005
R305 VTAIL.n105 VTAIL.n104 9.3005
R306 VTAIL.n103 VTAIL.n102 9.3005
R307 VTAIL.n194 VTAIL.n193 8.92171
R308 VTAIL.n26 VTAIL.n25 8.92171
R309 VTAIL.n141 VTAIL.n140 8.92171
R310 VTAIL.n85 VTAIL.n84 8.92171
R311 VTAIL.n190 VTAIL.n184 8.14595
R312 VTAIL.n22 VTAIL.n16 8.14595
R313 VTAIL.n137 VTAIL.n131 8.14595
R314 VTAIL.n81 VTAIL.n75 8.14595
R315 VTAIL.n189 VTAIL.n186 7.3702
R316 VTAIL.n21 VTAIL.n18 7.3702
R317 VTAIL.n136 VTAIL.n133 7.3702
R318 VTAIL.n80 VTAIL.n77 7.3702
R319 VTAIL.n190 VTAIL.n189 5.81868
R320 VTAIL.n22 VTAIL.n21 5.81868
R321 VTAIL.n137 VTAIL.n136 5.81868
R322 VTAIL.n81 VTAIL.n80 5.81868
R323 VTAIL.n193 VTAIL.n184 5.04292
R324 VTAIL.n25 VTAIL.n16 5.04292
R325 VTAIL.n140 VTAIL.n131 5.04292
R326 VTAIL.n84 VTAIL.n75 5.04292
R327 VTAIL.n194 VTAIL.n182 4.26717
R328 VTAIL.n26 VTAIL.n14 4.26717
R329 VTAIL.n141 VTAIL.n129 4.26717
R330 VTAIL.n85 VTAIL.n73 4.26717
R331 VTAIL.n198 VTAIL.n197 3.49141
R332 VTAIL.n222 VTAIL.n170 3.49141
R333 VTAIL.n30 VTAIL.n29 3.49141
R334 VTAIL.n54 VTAIL.n2 3.49141
R335 VTAIL.n168 VTAIL.n116 3.49141
R336 VTAIL.n145 VTAIL.n144 3.49141
R337 VTAIL.n112 VTAIL.n60 3.49141
R338 VTAIL.n89 VTAIL.n88 3.49141
R339 VTAIL.n113 VTAIL.n59 3.34533
R340 VTAIL.n169 VTAIL.n115 3.34533
R341 VTAIL.n57 VTAIL.n55 3.34533
R342 VTAIL.n0 VTAIL.t4 3.21882
R343 VTAIL.n0 VTAIL.t0 3.21882
R344 VTAIL.n56 VTAIL.t6 3.21882
R345 VTAIL.n56 VTAIL.t11 3.21882
R346 VTAIL.n114 VTAIL.t9 3.21882
R347 VTAIL.n114 VTAIL.t10 3.21882
R348 VTAIL.n58 VTAIL.t2 3.21882
R349 VTAIL.n58 VTAIL.t5 3.21882
R350 VTAIL.n201 VTAIL.n180 2.71565
R351 VTAIL.n220 VTAIL.n219 2.71565
R352 VTAIL.n33 VTAIL.n12 2.71565
R353 VTAIL.n52 VTAIL.n51 2.71565
R354 VTAIL.n166 VTAIL.n165 2.71565
R355 VTAIL.n148 VTAIL.n127 2.71565
R356 VTAIL.n110 VTAIL.n109 2.71565
R357 VTAIL.n92 VTAIL.n71 2.71565
R358 VTAIL VTAIL.n223 2.45093
R359 VTAIL.n188 VTAIL.n187 2.41283
R360 VTAIL.n20 VTAIL.n19 2.41283
R361 VTAIL.n135 VTAIL.n134 2.41283
R362 VTAIL.n79 VTAIL.n78 2.41283
R363 VTAIL.n115 VTAIL.n113 2.14274
R364 VTAIL.n55 VTAIL.n1 2.14274
R365 VTAIL.n202 VTAIL.n178 1.93989
R366 VTAIL.n216 VTAIL.n172 1.93989
R367 VTAIL.n34 VTAIL.n10 1.93989
R368 VTAIL.n48 VTAIL.n4 1.93989
R369 VTAIL.n162 VTAIL.n118 1.93989
R370 VTAIL.n149 VTAIL.n125 1.93989
R371 VTAIL.n106 VTAIL.n62 1.93989
R372 VTAIL.n93 VTAIL.n69 1.93989
R373 VTAIL.n207 VTAIL.n205 1.16414
R374 VTAIL.n215 VTAIL.n174 1.16414
R375 VTAIL.n39 VTAIL.n37 1.16414
R376 VTAIL.n47 VTAIL.n6 1.16414
R377 VTAIL.n161 VTAIL.n120 1.16414
R378 VTAIL.n153 VTAIL.n152 1.16414
R379 VTAIL.n105 VTAIL.n64 1.16414
R380 VTAIL.n97 VTAIL.n96 1.16414
R381 VTAIL VTAIL.n1 0.894897
R382 VTAIL.n206 VTAIL.n176 0.388379
R383 VTAIL.n212 VTAIL.n211 0.388379
R384 VTAIL.n38 VTAIL.n8 0.388379
R385 VTAIL.n44 VTAIL.n43 0.388379
R386 VTAIL.n158 VTAIL.n157 0.388379
R387 VTAIL.n124 VTAIL.n122 0.388379
R388 VTAIL.n102 VTAIL.n101 0.388379
R389 VTAIL.n68 VTAIL.n66 0.388379
R390 VTAIL.n188 VTAIL.n183 0.155672
R391 VTAIL.n195 VTAIL.n183 0.155672
R392 VTAIL.n196 VTAIL.n195 0.155672
R393 VTAIL.n196 VTAIL.n179 0.155672
R394 VTAIL.n203 VTAIL.n179 0.155672
R395 VTAIL.n204 VTAIL.n203 0.155672
R396 VTAIL.n204 VTAIL.n175 0.155672
R397 VTAIL.n213 VTAIL.n175 0.155672
R398 VTAIL.n214 VTAIL.n213 0.155672
R399 VTAIL.n214 VTAIL.n171 0.155672
R400 VTAIL.n221 VTAIL.n171 0.155672
R401 VTAIL.n20 VTAIL.n15 0.155672
R402 VTAIL.n27 VTAIL.n15 0.155672
R403 VTAIL.n28 VTAIL.n27 0.155672
R404 VTAIL.n28 VTAIL.n11 0.155672
R405 VTAIL.n35 VTAIL.n11 0.155672
R406 VTAIL.n36 VTAIL.n35 0.155672
R407 VTAIL.n36 VTAIL.n7 0.155672
R408 VTAIL.n45 VTAIL.n7 0.155672
R409 VTAIL.n46 VTAIL.n45 0.155672
R410 VTAIL.n46 VTAIL.n3 0.155672
R411 VTAIL.n53 VTAIL.n3 0.155672
R412 VTAIL.n167 VTAIL.n117 0.155672
R413 VTAIL.n160 VTAIL.n117 0.155672
R414 VTAIL.n160 VTAIL.n159 0.155672
R415 VTAIL.n159 VTAIL.n121 0.155672
R416 VTAIL.n151 VTAIL.n121 0.155672
R417 VTAIL.n151 VTAIL.n150 0.155672
R418 VTAIL.n150 VTAIL.n126 0.155672
R419 VTAIL.n143 VTAIL.n126 0.155672
R420 VTAIL.n143 VTAIL.n142 0.155672
R421 VTAIL.n142 VTAIL.n130 0.155672
R422 VTAIL.n135 VTAIL.n130 0.155672
R423 VTAIL.n111 VTAIL.n61 0.155672
R424 VTAIL.n104 VTAIL.n61 0.155672
R425 VTAIL.n104 VTAIL.n103 0.155672
R426 VTAIL.n103 VTAIL.n65 0.155672
R427 VTAIL.n95 VTAIL.n65 0.155672
R428 VTAIL.n95 VTAIL.n94 0.155672
R429 VTAIL.n94 VTAIL.n70 0.155672
R430 VTAIL.n87 VTAIL.n70 0.155672
R431 VTAIL.n87 VTAIL.n86 0.155672
R432 VTAIL.n86 VTAIL.n74 0.155672
R433 VTAIL.n79 VTAIL.n74 0.155672
R434 VDD1.n48 VDD1.n0 756.745
R435 VDD1.n101 VDD1.n53 756.745
R436 VDD1.n49 VDD1.n48 585
R437 VDD1.n47 VDD1.n46 585
R438 VDD1.n4 VDD1.n3 585
R439 VDD1.n41 VDD1.n40 585
R440 VDD1.n39 VDD1.n6 585
R441 VDD1.n38 VDD1.n37 585
R442 VDD1.n9 VDD1.n7 585
R443 VDD1.n32 VDD1.n31 585
R444 VDD1.n30 VDD1.n29 585
R445 VDD1.n13 VDD1.n12 585
R446 VDD1.n24 VDD1.n23 585
R447 VDD1.n22 VDD1.n21 585
R448 VDD1.n17 VDD1.n16 585
R449 VDD1.n69 VDD1.n68 585
R450 VDD1.n74 VDD1.n73 585
R451 VDD1.n76 VDD1.n75 585
R452 VDD1.n65 VDD1.n64 585
R453 VDD1.n82 VDD1.n81 585
R454 VDD1.n84 VDD1.n83 585
R455 VDD1.n61 VDD1.n60 585
R456 VDD1.n91 VDD1.n90 585
R457 VDD1.n92 VDD1.n59 585
R458 VDD1.n94 VDD1.n93 585
R459 VDD1.n57 VDD1.n56 585
R460 VDD1.n100 VDD1.n99 585
R461 VDD1.n102 VDD1.n101 585
R462 VDD1.n70 VDD1.t1 329.038
R463 VDD1.n18 VDD1.t0 329.038
R464 VDD1.n48 VDD1.n47 171.744
R465 VDD1.n47 VDD1.n3 171.744
R466 VDD1.n40 VDD1.n3 171.744
R467 VDD1.n40 VDD1.n39 171.744
R468 VDD1.n39 VDD1.n38 171.744
R469 VDD1.n38 VDD1.n7 171.744
R470 VDD1.n31 VDD1.n7 171.744
R471 VDD1.n31 VDD1.n30 171.744
R472 VDD1.n30 VDD1.n12 171.744
R473 VDD1.n23 VDD1.n12 171.744
R474 VDD1.n23 VDD1.n22 171.744
R475 VDD1.n22 VDD1.n16 171.744
R476 VDD1.n74 VDD1.n68 171.744
R477 VDD1.n75 VDD1.n74 171.744
R478 VDD1.n75 VDD1.n64 171.744
R479 VDD1.n82 VDD1.n64 171.744
R480 VDD1.n83 VDD1.n82 171.744
R481 VDD1.n83 VDD1.n60 171.744
R482 VDD1.n91 VDD1.n60 171.744
R483 VDD1.n92 VDD1.n91 171.744
R484 VDD1.n93 VDD1.n92 171.744
R485 VDD1.n93 VDD1.n56 171.744
R486 VDD1.n100 VDD1.n56 171.744
R487 VDD1.n101 VDD1.n100 171.744
R488 VDD1.t0 VDD1.n16 85.8723
R489 VDD1.t1 VDD1.n68 85.8723
R490 VDD1.n107 VDD1.n106 80.6148
R491 VDD1.n109 VDD1.n108 79.8339
R492 VDD1 VDD1.n52 54.1461
R493 VDD1.n107 VDD1.n105 54.0326
R494 VDD1.n109 VDD1.n107 45.5483
R495 VDD1.n41 VDD1.n6 13.1884
R496 VDD1.n94 VDD1.n59 13.1884
R497 VDD1.n42 VDD1.n4 12.8005
R498 VDD1.n37 VDD1.n8 12.8005
R499 VDD1.n90 VDD1.n89 12.8005
R500 VDD1.n95 VDD1.n57 12.8005
R501 VDD1.n46 VDD1.n45 12.0247
R502 VDD1.n36 VDD1.n9 12.0247
R503 VDD1.n88 VDD1.n61 12.0247
R504 VDD1.n99 VDD1.n98 12.0247
R505 VDD1.n49 VDD1.n2 11.249
R506 VDD1.n33 VDD1.n32 11.249
R507 VDD1.n85 VDD1.n84 11.249
R508 VDD1.n102 VDD1.n55 11.249
R509 VDD1.n18 VDD1.n17 10.7239
R510 VDD1.n70 VDD1.n69 10.7239
R511 VDD1.n50 VDD1.n0 10.4732
R512 VDD1.n29 VDD1.n11 10.4732
R513 VDD1.n81 VDD1.n63 10.4732
R514 VDD1.n103 VDD1.n53 10.4732
R515 VDD1.n28 VDD1.n13 9.69747
R516 VDD1.n80 VDD1.n65 9.69747
R517 VDD1.n52 VDD1.n51 9.45567
R518 VDD1.n105 VDD1.n104 9.45567
R519 VDD1.n20 VDD1.n19 9.3005
R520 VDD1.n15 VDD1.n14 9.3005
R521 VDD1.n26 VDD1.n25 9.3005
R522 VDD1.n28 VDD1.n27 9.3005
R523 VDD1.n11 VDD1.n10 9.3005
R524 VDD1.n34 VDD1.n33 9.3005
R525 VDD1.n36 VDD1.n35 9.3005
R526 VDD1.n8 VDD1.n5 9.3005
R527 VDD1.n51 VDD1.n50 9.3005
R528 VDD1.n2 VDD1.n1 9.3005
R529 VDD1.n45 VDD1.n44 9.3005
R530 VDD1.n43 VDD1.n42 9.3005
R531 VDD1.n104 VDD1.n103 9.3005
R532 VDD1.n55 VDD1.n54 9.3005
R533 VDD1.n98 VDD1.n97 9.3005
R534 VDD1.n96 VDD1.n95 9.3005
R535 VDD1.n72 VDD1.n71 9.3005
R536 VDD1.n67 VDD1.n66 9.3005
R537 VDD1.n78 VDD1.n77 9.3005
R538 VDD1.n80 VDD1.n79 9.3005
R539 VDD1.n63 VDD1.n62 9.3005
R540 VDD1.n86 VDD1.n85 9.3005
R541 VDD1.n88 VDD1.n87 9.3005
R542 VDD1.n89 VDD1.n58 9.3005
R543 VDD1.n25 VDD1.n24 8.92171
R544 VDD1.n77 VDD1.n76 8.92171
R545 VDD1.n21 VDD1.n15 8.14595
R546 VDD1.n73 VDD1.n67 8.14595
R547 VDD1.n20 VDD1.n17 7.3702
R548 VDD1.n72 VDD1.n69 7.3702
R549 VDD1.n21 VDD1.n20 5.81868
R550 VDD1.n73 VDD1.n72 5.81868
R551 VDD1.n24 VDD1.n15 5.04292
R552 VDD1.n76 VDD1.n67 5.04292
R553 VDD1.n25 VDD1.n13 4.26717
R554 VDD1.n77 VDD1.n65 4.26717
R555 VDD1.n52 VDD1.n0 3.49141
R556 VDD1.n29 VDD1.n28 3.49141
R557 VDD1.n81 VDD1.n80 3.49141
R558 VDD1.n105 VDD1.n53 3.49141
R559 VDD1.n108 VDD1.t3 3.21882
R560 VDD1.n108 VDD1.t2 3.21882
R561 VDD1.n106 VDD1.t4 3.21882
R562 VDD1.n106 VDD1.t5 3.21882
R563 VDD1.n50 VDD1.n49 2.71565
R564 VDD1.n32 VDD1.n11 2.71565
R565 VDD1.n84 VDD1.n63 2.71565
R566 VDD1.n103 VDD1.n102 2.71565
R567 VDD1.n19 VDD1.n18 2.41283
R568 VDD1.n71 VDD1.n70 2.41283
R569 VDD1.n46 VDD1.n2 1.93989
R570 VDD1.n33 VDD1.n9 1.93989
R571 VDD1.n85 VDD1.n61 1.93989
R572 VDD1.n99 VDD1.n55 1.93989
R573 VDD1.n45 VDD1.n4 1.16414
R574 VDD1.n37 VDD1.n36 1.16414
R575 VDD1.n90 VDD1.n88 1.16414
R576 VDD1.n98 VDD1.n57 1.16414
R577 VDD1 VDD1.n109 0.778517
R578 VDD1.n42 VDD1.n41 0.388379
R579 VDD1.n8 VDD1.n6 0.388379
R580 VDD1.n89 VDD1.n59 0.388379
R581 VDD1.n95 VDD1.n94 0.388379
R582 VDD1.n51 VDD1.n1 0.155672
R583 VDD1.n44 VDD1.n1 0.155672
R584 VDD1.n44 VDD1.n43 0.155672
R585 VDD1.n43 VDD1.n5 0.155672
R586 VDD1.n35 VDD1.n5 0.155672
R587 VDD1.n35 VDD1.n34 0.155672
R588 VDD1.n34 VDD1.n10 0.155672
R589 VDD1.n27 VDD1.n10 0.155672
R590 VDD1.n27 VDD1.n26 0.155672
R591 VDD1.n26 VDD1.n14 0.155672
R592 VDD1.n19 VDD1.n14 0.155672
R593 VDD1.n71 VDD1.n66 0.155672
R594 VDD1.n78 VDD1.n66 0.155672
R595 VDD1.n79 VDD1.n78 0.155672
R596 VDD1.n79 VDD1.n62 0.155672
R597 VDD1.n86 VDD1.n62 0.155672
R598 VDD1.n87 VDD1.n86 0.155672
R599 VDD1.n87 VDD1.n58 0.155672
R600 VDD1.n96 VDD1.n58 0.155672
R601 VDD1.n97 VDD1.n96 0.155672
R602 VDD1.n97 VDD1.n54 0.155672
R603 VDD1.n104 VDD1.n54 0.155672
R604 VN.n38 VN.n37 161.3
R605 VN.n36 VN.n21 161.3
R606 VN.n35 VN.n34 161.3
R607 VN.n33 VN.n22 161.3
R608 VN.n32 VN.n31 161.3
R609 VN.n30 VN.n23 161.3
R610 VN.n29 VN.n28 161.3
R611 VN.n27 VN.n24 161.3
R612 VN.n18 VN.n17 161.3
R613 VN.n16 VN.n1 161.3
R614 VN.n15 VN.n14 161.3
R615 VN.n13 VN.n2 161.3
R616 VN.n12 VN.n11 161.3
R617 VN.n10 VN.n3 161.3
R618 VN.n9 VN.n8 161.3
R619 VN.n7 VN.n4 161.3
R620 VN.n26 VN.t1 101.382
R621 VN.n6 VN.t2 101.382
R622 VN.n19 VN.n0 83.8517
R623 VN.n39 VN.n20 83.8517
R624 VN.n5 VN.t4 68.5667
R625 VN.n0 VN.t3 68.5667
R626 VN.n25 VN.t5 68.5667
R627 VN.n20 VN.t0 68.5667
R628 VN.n6 VN.n5 62.4228
R629 VN.n26 VN.n25 62.4228
R630 VN.n11 VN.n2 56.5617
R631 VN.n31 VN.n22 56.5617
R632 VN VN.n39 51.1724
R633 VN.n9 VN.n4 24.5923
R634 VN.n10 VN.n9 24.5923
R635 VN.n11 VN.n10 24.5923
R636 VN.n15 VN.n2 24.5923
R637 VN.n16 VN.n15 24.5923
R638 VN.n17 VN.n16 24.5923
R639 VN.n31 VN.n30 24.5923
R640 VN.n30 VN.n29 24.5923
R641 VN.n29 VN.n24 24.5923
R642 VN.n37 VN.n36 24.5923
R643 VN.n36 VN.n35 24.5923
R644 VN.n35 VN.n22 24.5923
R645 VN.n5 VN.n4 12.2964
R646 VN.n25 VN.n24 12.2964
R647 VN.n17 VN.n0 6.39438
R648 VN.n37 VN.n20 6.39438
R649 VN.n27 VN.n26 3.26269
R650 VN.n7 VN.n6 3.26269
R651 VN.n39 VN.n38 0.354861
R652 VN.n19 VN.n18 0.354861
R653 VN VN.n19 0.267071
R654 VN.n38 VN.n21 0.189894
R655 VN.n34 VN.n21 0.189894
R656 VN.n34 VN.n33 0.189894
R657 VN.n33 VN.n32 0.189894
R658 VN.n32 VN.n23 0.189894
R659 VN.n28 VN.n23 0.189894
R660 VN.n28 VN.n27 0.189894
R661 VN.n8 VN.n7 0.189894
R662 VN.n8 VN.n3 0.189894
R663 VN.n12 VN.n3 0.189894
R664 VN.n13 VN.n12 0.189894
R665 VN.n14 VN.n13 0.189894
R666 VN.n14 VN.n1 0.189894
R667 VN.n18 VN.n1 0.189894
R668 VDD2.n103 VDD2.n55 756.745
R669 VDD2.n48 VDD2.n0 756.745
R670 VDD2.n104 VDD2.n103 585
R671 VDD2.n102 VDD2.n101 585
R672 VDD2.n59 VDD2.n58 585
R673 VDD2.n96 VDD2.n95 585
R674 VDD2.n94 VDD2.n61 585
R675 VDD2.n93 VDD2.n92 585
R676 VDD2.n64 VDD2.n62 585
R677 VDD2.n87 VDD2.n86 585
R678 VDD2.n85 VDD2.n84 585
R679 VDD2.n68 VDD2.n67 585
R680 VDD2.n79 VDD2.n78 585
R681 VDD2.n77 VDD2.n76 585
R682 VDD2.n72 VDD2.n71 585
R683 VDD2.n16 VDD2.n15 585
R684 VDD2.n21 VDD2.n20 585
R685 VDD2.n23 VDD2.n22 585
R686 VDD2.n12 VDD2.n11 585
R687 VDD2.n29 VDD2.n28 585
R688 VDD2.n31 VDD2.n30 585
R689 VDD2.n8 VDD2.n7 585
R690 VDD2.n38 VDD2.n37 585
R691 VDD2.n39 VDD2.n6 585
R692 VDD2.n41 VDD2.n40 585
R693 VDD2.n4 VDD2.n3 585
R694 VDD2.n47 VDD2.n46 585
R695 VDD2.n49 VDD2.n48 585
R696 VDD2.n17 VDD2.t3 329.038
R697 VDD2.n73 VDD2.t5 329.038
R698 VDD2.n103 VDD2.n102 171.744
R699 VDD2.n102 VDD2.n58 171.744
R700 VDD2.n95 VDD2.n58 171.744
R701 VDD2.n95 VDD2.n94 171.744
R702 VDD2.n94 VDD2.n93 171.744
R703 VDD2.n93 VDD2.n62 171.744
R704 VDD2.n86 VDD2.n62 171.744
R705 VDD2.n86 VDD2.n85 171.744
R706 VDD2.n85 VDD2.n67 171.744
R707 VDD2.n78 VDD2.n67 171.744
R708 VDD2.n78 VDD2.n77 171.744
R709 VDD2.n77 VDD2.n71 171.744
R710 VDD2.n21 VDD2.n15 171.744
R711 VDD2.n22 VDD2.n21 171.744
R712 VDD2.n22 VDD2.n11 171.744
R713 VDD2.n29 VDD2.n11 171.744
R714 VDD2.n30 VDD2.n29 171.744
R715 VDD2.n30 VDD2.n7 171.744
R716 VDD2.n38 VDD2.n7 171.744
R717 VDD2.n39 VDD2.n38 171.744
R718 VDD2.n40 VDD2.n39 171.744
R719 VDD2.n40 VDD2.n3 171.744
R720 VDD2.n47 VDD2.n3 171.744
R721 VDD2.n48 VDD2.n47 171.744
R722 VDD2.t5 VDD2.n71 85.8723
R723 VDD2.t3 VDD2.n15 85.8723
R724 VDD2.n54 VDD2.n53 80.6148
R725 VDD2 VDD2.n109 80.612
R726 VDD2.n54 VDD2.n52 54.0326
R727 VDD2.n108 VDD2.n107 51.5793
R728 VDD2.n108 VDD2.n54 43.2929
R729 VDD2.n96 VDD2.n61 13.1884
R730 VDD2.n41 VDD2.n6 13.1884
R731 VDD2.n97 VDD2.n59 12.8005
R732 VDD2.n92 VDD2.n63 12.8005
R733 VDD2.n37 VDD2.n36 12.8005
R734 VDD2.n42 VDD2.n4 12.8005
R735 VDD2.n101 VDD2.n100 12.0247
R736 VDD2.n91 VDD2.n64 12.0247
R737 VDD2.n35 VDD2.n8 12.0247
R738 VDD2.n46 VDD2.n45 12.0247
R739 VDD2.n104 VDD2.n57 11.249
R740 VDD2.n88 VDD2.n87 11.249
R741 VDD2.n32 VDD2.n31 11.249
R742 VDD2.n49 VDD2.n2 11.249
R743 VDD2.n73 VDD2.n72 10.7239
R744 VDD2.n17 VDD2.n16 10.7239
R745 VDD2.n105 VDD2.n55 10.4732
R746 VDD2.n84 VDD2.n66 10.4732
R747 VDD2.n28 VDD2.n10 10.4732
R748 VDD2.n50 VDD2.n0 10.4732
R749 VDD2.n83 VDD2.n68 9.69747
R750 VDD2.n27 VDD2.n12 9.69747
R751 VDD2.n107 VDD2.n106 9.45567
R752 VDD2.n52 VDD2.n51 9.45567
R753 VDD2.n75 VDD2.n74 9.3005
R754 VDD2.n70 VDD2.n69 9.3005
R755 VDD2.n81 VDD2.n80 9.3005
R756 VDD2.n83 VDD2.n82 9.3005
R757 VDD2.n66 VDD2.n65 9.3005
R758 VDD2.n89 VDD2.n88 9.3005
R759 VDD2.n91 VDD2.n90 9.3005
R760 VDD2.n63 VDD2.n60 9.3005
R761 VDD2.n106 VDD2.n105 9.3005
R762 VDD2.n57 VDD2.n56 9.3005
R763 VDD2.n100 VDD2.n99 9.3005
R764 VDD2.n98 VDD2.n97 9.3005
R765 VDD2.n51 VDD2.n50 9.3005
R766 VDD2.n2 VDD2.n1 9.3005
R767 VDD2.n45 VDD2.n44 9.3005
R768 VDD2.n43 VDD2.n42 9.3005
R769 VDD2.n19 VDD2.n18 9.3005
R770 VDD2.n14 VDD2.n13 9.3005
R771 VDD2.n25 VDD2.n24 9.3005
R772 VDD2.n27 VDD2.n26 9.3005
R773 VDD2.n10 VDD2.n9 9.3005
R774 VDD2.n33 VDD2.n32 9.3005
R775 VDD2.n35 VDD2.n34 9.3005
R776 VDD2.n36 VDD2.n5 9.3005
R777 VDD2.n80 VDD2.n79 8.92171
R778 VDD2.n24 VDD2.n23 8.92171
R779 VDD2.n76 VDD2.n70 8.14595
R780 VDD2.n20 VDD2.n14 8.14595
R781 VDD2.n75 VDD2.n72 7.3702
R782 VDD2.n19 VDD2.n16 7.3702
R783 VDD2.n76 VDD2.n75 5.81868
R784 VDD2.n20 VDD2.n19 5.81868
R785 VDD2.n79 VDD2.n70 5.04292
R786 VDD2.n23 VDD2.n14 5.04292
R787 VDD2.n80 VDD2.n68 4.26717
R788 VDD2.n24 VDD2.n12 4.26717
R789 VDD2.n107 VDD2.n55 3.49141
R790 VDD2.n84 VDD2.n83 3.49141
R791 VDD2.n28 VDD2.n27 3.49141
R792 VDD2.n52 VDD2.n0 3.49141
R793 VDD2.n109 VDD2.t0 3.21882
R794 VDD2.n109 VDD2.t4 3.21882
R795 VDD2.n53 VDD2.t1 3.21882
R796 VDD2.n53 VDD2.t2 3.21882
R797 VDD2.n105 VDD2.n104 2.71565
R798 VDD2.n87 VDD2.n66 2.71565
R799 VDD2.n31 VDD2.n10 2.71565
R800 VDD2.n50 VDD2.n49 2.71565
R801 VDD2 VDD2.n108 2.56731
R802 VDD2.n74 VDD2.n73 2.41283
R803 VDD2.n18 VDD2.n17 2.41283
R804 VDD2.n101 VDD2.n57 1.93989
R805 VDD2.n88 VDD2.n64 1.93989
R806 VDD2.n32 VDD2.n8 1.93989
R807 VDD2.n46 VDD2.n2 1.93989
R808 VDD2.n100 VDD2.n59 1.16414
R809 VDD2.n92 VDD2.n91 1.16414
R810 VDD2.n37 VDD2.n35 1.16414
R811 VDD2.n45 VDD2.n4 1.16414
R812 VDD2.n97 VDD2.n96 0.388379
R813 VDD2.n63 VDD2.n61 0.388379
R814 VDD2.n36 VDD2.n6 0.388379
R815 VDD2.n42 VDD2.n41 0.388379
R816 VDD2.n106 VDD2.n56 0.155672
R817 VDD2.n99 VDD2.n56 0.155672
R818 VDD2.n99 VDD2.n98 0.155672
R819 VDD2.n98 VDD2.n60 0.155672
R820 VDD2.n90 VDD2.n60 0.155672
R821 VDD2.n90 VDD2.n89 0.155672
R822 VDD2.n89 VDD2.n65 0.155672
R823 VDD2.n82 VDD2.n65 0.155672
R824 VDD2.n82 VDD2.n81 0.155672
R825 VDD2.n81 VDD2.n69 0.155672
R826 VDD2.n74 VDD2.n69 0.155672
R827 VDD2.n18 VDD2.n13 0.155672
R828 VDD2.n25 VDD2.n13 0.155672
R829 VDD2.n26 VDD2.n25 0.155672
R830 VDD2.n26 VDD2.n9 0.155672
R831 VDD2.n33 VDD2.n9 0.155672
R832 VDD2.n34 VDD2.n33 0.155672
R833 VDD2.n34 VDD2.n5 0.155672
R834 VDD2.n43 VDD2.n5 0.155672
R835 VDD2.n44 VDD2.n43 0.155672
R836 VDD2.n44 VDD2.n1 0.155672
R837 VDD2.n51 VDD2.n1 0.155672
R838 B.n402 B.n401 585
R839 B.n400 B.n129 585
R840 B.n399 B.n398 585
R841 B.n397 B.n130 585
R842 B.n396 B.n395 585
R843 B.n394 B.n131 585
R844 B.n393 B.n392 585
R845 B.n391 B.n132 585
R846 B.n390 B.n389 585
R847 B.n388 B.n133 585
R848 B.n387 B.n386 585
R849 B.n385 B.n134 585
R850 B.n384 B.n383 585
R851 B.n382 B.n135 585
R852 B.n381 B.n380 585
R853 B.n379 B.n136 585
R854 B.n378 B.n377 585
R855 B.n376 B.n137 585
R856 B.n375 B.n374 585
R857 B.n373 B.n138 585
R858 B.n372 B.n371 585
R859 B.n370 B.n139 585
R860 B.n369 B.n368 585
R861 B.n367 B.n140 585
R862 B.n366 B.n365 585
R863 B.n364 B.n141 585
R864 B.n363 B.n362 585
R865 B.n361 B.n142 585
R866 B.n360 B.n359 585
R867 B.n358 B.n143 585
R868 B.n357 B.n356 585
R869 B.n355 B.n144 585
R870 B.n354 B.n353 585
R871 B.n352 B.n145 585
R872 B.n351 B.n350 585
R873 B.n349 B.n146 585
R874 B.n347 B.n346 585
R875 B.n345 B.n149 585
R876 B.n344 B.n343 585
R877 B.n342 B.n150 585
R878 B.n341 B.n340 585
R879 B.n339 B.n151 585
R880 B.n338 B.n337 585
R881 B.n336 B.n152 585
R882 B.n335 B.n334 585
R883 B.n333 B.n153 585
R884 B.n332 B.n331 585
R885 B.n327 B.n154 585
R886 B.n326 B.n325 585
R887 B.n324 B.n155 585
R888 B.n323 B.n322 585
R889 B.n321 B.n156 585
R890 B.n320 B.n319 585
R891 B.n318 B.n157 585
R892 B.n317 B.n316 585
R893 B.n315 B.n158 585
R894 B.n314 B.n313 585
R895 B.n312 B.n159 585
R896 B.n311 B.n310 585
R897 B.n309 B.n160 585
R898 B.n308 B.n307 585
R899 B.n306 B.n161 585
R900 B.n305 B.n304 585
R901 B.n303 B.n162 585
R902 B.n302 B.n301 585
R903 B.n300 B.n163 585
R904 B.n299 B.n298 585
R905 B.n297 B.n164 585
R906 B.n296 B.n295 585
R907 B.n294 B.n165 585
R908 B.n293 B.n292 585
R909 B.n291 B.n166 585
R910 B.n290 B.n289 585
R911 B.n288 B.n167 585
R912 B.n287 B.n286 585
R913 B.n285 B.n168 585
R914 B.n284 B.n283 585
R915 B.n282 B.n169 585
R916 B.n281 B.n280 585
R917 B.n279 B.n170 585
R918 B.n278 B.n277 585
R919 B.n276 B.n171 585
R920 B.n403 B.n128 585
R921 B.n405 B.n404 585
R922 B.n406 B.n127 585
R923 B.n408 B.n407 585
R924 B.n409 B.n126 585
R925 B.n411 B.n410 585
R926 B.n412 B.n125 585
R927 B.n414 B.n413 585
R928 B.n415 B.n124 585
R929 B.n417 B.n416 585
R930 B.n418 B.n123 585
R931 B.n420 B.n419 585
R932 B.n421 B.n122 585
R933 B.n423 B.n422 585
R934 B.n424 B.n121 585
R935 B.n426 B.n425 585
R936 B.n427 B.n120 585
R937 B.n429 B.n428 585
R938 B.n430 B.n119 585
R939 B.n432 B.n431 585
R940 B.n433 B.n118 585
R941 B.n435 B.n434 585
R942 B.n436 B.n117 585
R943 B.n438 B.n437 585
R944 B.n439 B.n116 585
R945 B.n441 B.n440 585
R946 B.n442 B.n115 585
R947 B.n444 B.n443 585
R948 B.n445 B.n114 585
R949 B.n447 B.n446 585
R950 B.n448 B.n113 585
R951 B.n450 B.n449 585
R952 B.n451 B.n112 585
R953 B.n453 B.n452 585
R954 B.n454 B.n111 585
R955 B.n456 B.n455 585
R956 B.n457 B.n110 585
R957 B.n459 B.n458 585
R958 B.n460 B.n109 585
R959 B.n462 B.n461 585
R960 B.n463 B.n108 585
R961 B.n465 B.n464 585
R962 B.n466 B.n107 585
R963 B.n468 B.n467 585
R964 B.n469 B.n106 585
R965 B.n471 B.n470 585
R966 B.n472 B.n105 585
R967 B.n474 B.n473 585
R968 B.n475 B.n104 585
R969 B.n477 B.n476 585
R970 B.n478 B.n103 585
R971 B.n480 B.n479 585
R972 B.n481 B.n102 585
R973 B.n483 B.n482 585
R974 B.n484 B.n101 585
R975 B.n486 B.n485 585
R976 B.n487 B.n100 585
R977 B.n489 B.n488 585
R978 B.n490 B.n99 585
R979 B.n492 B.n491 585
R980 B.n493 B.n98 585
R981 B.n495 B.n494 585
R982 B.n496 B.n97 585
R983 B.n498 B.n497 585
R984 B.n499 B.n96 585
R985 B.n501 B.n500 585
R986 B.n502 B.n95 585
R987 B.n504 B.n503 585
R988 B.n505 B.n94 585
R989 B.n507 B.n506 585
R990 B.n508 B.n93 585
R991 B.n510 B.n509 585
R992 B.n511 B.n92 585
R993 B.n513 B.n512 585
R994 B.n514 B.n91 585
R995 B.n516 B.n515 585
R996 B.n517 B.n90 585
R997 B.n519 B.n518 585
R998 B.n520 B.n89 585
R999 B.n522 B.n521 585
R1000 B.n523 B.n88 585
R1001 B.n525 B.n524 585
R1002 B.n526 B.n87 585
R1003 B.n528 B.n527 585
R1004 B.n529 B.n86 585
R1005 B.n531 B.n530 585
R1006 B.n532 B.n85 585
R1007 B.n534 B.n533 585
R1008 B.n535 B.n84 585
R1009 B.n537 B.n536 585
R1010 B.n538 B.n83 585
R1011 B.n540 B.n539 585
R1012 B.n541 B.n82 585
R1013 B.n543 B.n542 585
R1014 B.n544 B.n81 585
R1015 B.n546 B.n545 585
R1016 B.n547 B.n80 585
R1017 B.n549 B.n548 585
R1018 B.n550 B.n79 585
R1019 B.n552 B.n551 585
R1020 B.n553 B.n78 585
R1021 B.n555 B.n554 585
R1022 B.n556 B.n77 585
R1023 B.n558 B.n557 585
R1024 B.n559 B.n76 585
R1025 B.n561 B.n560 585
R1026 B.n562 B.n75 585
R1027 B.n564 B.n563 585
R1028 B.n688 B.n687 585
R1029 B.n686 B.n29 585
R1030 B.n685 B.n684 585
R1031 B.n683 B.n30 585
R1032 B.n682 B.n681 585
R1033 B.n680 B.n31 585
R1034 B.n679 B.n678 585
R1035 B.n677 B.n32 585
R1036 B.n676 B.n675 585
R1037 B.n674 B.n33 585
R1038 B.n673 B.n672 585
R1039 B.n671 B.n34 585
R1040 B.n670 B.n669 585
R1041 B.n668 B.n35 585
R1042 B.n667 B.n666 585
R1043 B.n665 B.n36 585
R1044 B.n664 B.n663 585
R1045 B.n662 B.n37 585
R1046 B.n661 B.n660 585
R1047 B.n659 B.n38 585
R1048 B.n658 B.n657 585
R1049 B.n656 B.n39 585
R1050 B.n655 B.n654 585
R1051 B.n653 B.n40 585
R1052 B.n652 B.n651 585
R1053 B.n650 B.n41 585
R1054 B.n649 B.n648 585
R1055 B.n647 B.n42 585
R1056 B.n646 B.n645 585
R1057 B.n644 B.n43 585
R1058 B.n643 B.n642 585
R1059 B.n641 B.n44 585
R1060 B.n640 B.n639 585
R1061 B.n638 B.n45 585
R1062 B.n637 B.n636 585
R1063 B.n635 B.n46 585
R1064 B.n634 B.n633 585
R1065 B.n632 B.n47 585
R1066 B.n631 B.n630 585
R1067 B.n629 B.n51 585
R1068 B.n628 B.n627 585
R1069 B.n626 B.n52 585
R1070 B.n625 B.n624 585
R1071 B.n623 B.n53 585
R1072 B.n622 B.n621 585
R1073 B.n620 B.n54 585
R1074 B.n618 B.n617 585
R1075 B.n616 B.n57 585
R1076 B.n615 B.n614 585
R1077 B.n613 B.n58 585
R1078 B.n612 B.n611 585
R1079 B.n610 B.n59 585
R1080 B.n609 B.n608 585
R1081 B.n607 B.n60 585
R1082 B.n606 B.n605 585
R1083 B.n604 B.n61 585
R1084 B.n603 B.n602 585
R1085 B.n601 B.n62 585
R1086 B.n600 B.n599 585
R1087 B.n598 B.n63 585
R1088 B.n597 B.n596 585
R1089 B.n595 B.n64 585
R1090 B.n594 B.n593 585
R1091 B.n592 B.n65 585
R1092 B.n591 B.n590 585
R1093 B.n589 B.n66 585
R1094 B.n588 B.n587 585
R1095 B.n586 B.n67 585
R1096 B.n585 B.n584 585
R1097 B.n583 B.n68 585
R1098 B.n582 B.n581 585
R1099 B.n580 B.n69 585
R1100 B.n579 B.n578 585
R1101 B.n577 B.n70 585
R1102 B.n576 B.n575 585
R1103 B.n574 B.n71 585
R1104 B.n573 B.n572 585
R1105 B.n571 B.n72 585
R1106 B.n570 B.n569 585
R1107 B.n568 B.n73 585
R1108 B.n567 B.n566 585
R1109 B.n565 B.n74 585
R1110 B.n689 B.n28 585
R1111 B.n691 B.n690 585
R1112 B.n692 B.n27 585
R1113 B.n694 B.n693 585
R1114 B.n695 B.n26 585
R1115 B.n697 B.n696 585
R1116 B.n698 B.n25 585
R1117 B.n700 B.n699 585
R1118 B.n701 B.n24 585
R1119 B.n703 B.n702 585
R1120 B.n704 B.n23 585
R1121 B.n706 B.n705 585
R1122 B.n707 B.n22 585
R1123 B.n709 B.n708 585
R1124 B.n710 B.n21 585
R1125 B.n712 B.n711 585
R1126 B.n713 B.n20 585
R1127 B.n715 B.n714 585
R1128 B.n716 B.n19 585
R1129 B.n718 B.n717 585
R1130 B.n719 B.n18 585
R1131 B.n721 B.n720 585
R1132 B.n722 B.n17 585
R1133 B.n724 B.n723 585
R1134 B.n725 B.n16 585
R1135 B.n727 B.n726 585
R1136 B.n728 B.n15 585
R1137 B.n730 B.n729 585
R1138 B.n731 B.n14 585
R1139 B.n733 B.n732 585
R1140 B.n734 B.n13 585
R1141 B.n736 B.n735 585
R1142 B.n737 B.n12 585
R1143 B.n739 B.n738 585
R1144 B.n740 B.n11 585
R1145 B.n742 B.n741 585
R1146 B.n743 B.n10 585
R1147 B.n745 B.n744 585
R1148 B.n746 B.n9 585
R1149 B.n748 B.n747 585
R1150 B.n749 B.n8 585
R1151 B.n751 B.n750 585
R1152 B.n752 B.n7 585
R1153 B.n754 B.n753 585
R1154 B.n755 B.n6 585
R1155 B.n757 B.n756 585
R1156 B.n758 B.n5 585
R1157 B.n760 B.n759 585
R1158 B.n761 B.n4 585
R1159 B.n763 B.n762 585
R1160 B.n764 B.n3 585
R1161 B.n766 B.n765 585
R1162 B.n767 B.n0 585
R1163 B.n2 B.n1 585
R1164 B.n198 B.n197 585
R1165 B.n200 B.n199 585
R1166 B.n201 B.n196 585
R1167 B.n203 B.n202 585
R1168 B.n204 B.n195 585
R1169 B.n206 B.n205 585
R1170 B.n207 B.n194 585
R1171 B.n209 B.n208 585
R1172 B.n210 B.n193 585
R1173 B.n212 B.n211 585
R1174 B.n213 B.n192 585
R1175 B.n215 B.n214 585
R1176 B.n216 B.n191 585
R1177 B.n218 B.n217 585
R1178 B.n219 B.n190 585
R1179 B.n221 B.n220 585
R1180 B.n222 B.n189 585
R1181 B.n224 B.n223 585
R1182 B.n225 B.n188 585
R1183 B.n227 B.n226 585
R1184 B.n228 B.n187 585
R1185 B.n230 B.n229 585
R1186 B.n231 B.n186 585
R1187 B.n233 B.n232 585
R1188 B.n234 B.n185 585
R1189 B.n236 B.n235 585
R1190 B.n237 B.n184 585
R1191 B.n239 B.n238 585
R1192 B.n240 B.n183 585
R1193 B.n242 B.n241 585
R1194 B.n243 B.n182 585
R1195 B.n245 B.n244 585
R1196 B.n246 B.n181 585
R1197 B.n248 B.n247 585
R1198 B.n249 B.n180 585
R1199 B.n251 B.n250 585
R1200 B.n252 B.n179 585
R1201 B.n254 B.n253 585
R1202 B.n255 B.n178 585
R1203 B.n257 B.n256 585
R1204 B.n258 B.n177 585
R1205 B.n260 B.n259 585
R1206 B.n261 B.n176 585
R1207 B.n263 B.n262 585
R1208 B.n264 B.n175 585
R1209 B.n266 B.n265 585
R1210 B.n267 B.n174 585
R1211 B.n269 B.n268 585
R1212 B.n270 B.n173 585
R1213 B.n272 B.n271 585
R1214 B.n273 B.n172 585
R1215 B.n275 B.n274 585
R1216 B.n276 B.n275 511.721
R1217 B.n401 B.n128 511.721
R1218 B.n563 B.n74 511.721
R1219 B.n689 B.n688 511.721
R1220 B.n147 B.t10 416.764
R1221 B.n55 B.t8 416.764
R1222 B.n328 B.t1 416.764
R1223 B.n48 B.t5 416.764
R1224 B.n148 B.t11 341.515
R1225 B.n56 B.t7 341.515
R1226 B.n329 B.t2 341.515
R1227 B.n49 B.t4 341.515
R1228 B.n328 B.t0 277.704
R1229 B.n147 B.t9 277.704
R1230 B.n55 B.t6 277.704
R1231 B.n48 B.t3 277.704
R1232 B.n769 B.n768 256.663
R1233 B.n768 B.n767 235.042
R1234 B.n768 B.n2 235.042
R1235 B.n277 B.n276 163.367
R1236 B.n277 B.n170 163.367
R1237 B.n281 B.n170 163.367
R1238 B.n282 B.n281 163.367
R1239 B.n283 B.n282 163.367
R1240 B.n283 B.n168 163.367
R1241 B.n287 B.n168 163.367
R1242 B.n288 B.n287 163.367
R1243 B.n289 B.n288 163.367
R1244 B.n289 B.n166 163.367
R1245 B.n293 B.n166 163.367
R1246 B.n294 B.n293 163.367
R1247 B.n295 B.n294 163.367
R1248 B.n295 B.n164 163.367
R1249 B.n299 B.n164 163.367
R1250 B.n300 B.n299 163.367
R1251 B.n301 B.n300 163.367
R1252 B.n301 B.n162 163.367
R1253 B.n305 B.n162 163.367
R1254 B.n306 B.n305 163.367
R1255 B.n307 B.n306 163.367
R1256 B.n307 B.n160 163.367
R1257 B.n311 B.n160 163.367
R1258 B.n312 B.n311 163.367
R1259 B.n313 B.n312 163.367
R1260 B.n313 B.n158 163.367
R1261 B.n317 B.n158 163.367
R1262 B.n318 B.n317 163.367
R1263 B.n319 B.n318 163.367
R1264 B.n319 B.n156 163.367
R1265 B.n323 B.n156 163.367
R1266 B.n324 B.n323 163.367
R1267 B.n325 B.n324 163.367
R1268 B.n325 B.n154 163.367
R1269 B.n332 B.n154 163.367
R1270 B.n333 B.n332 163.367
R1271 B.n334 B.n333 163.367
R1272 B.n334 B.n152 163.367
R1273 B.n338 B.n152 163.367
R1274 B.n339 B.n338 163.367
R1275 B.n340 B.n339 163.367
R1276 B.n340 B.n150 163.367
R1277 B.n344 B.n150 163.367
R1278 B.n345 B.n344 163.367
R1279 B.n346 B.n345 163.367
R1280 B.n346 B.n146 163.367
R1281 B.n351 B.n146 163.367
R1282 B.n352 B.n351 163.367
R1283 B.n353 B.n352 163.367
R1284 B.n353 B.n144 163.367
R1285 B.n357 B.n144 163.367
R1286 B.n358 B.n357 163.367
R1287 B.n359 B.n358 163.367
R1288 B.n359 B.n142 163.367
R1289 B.n363 B.n142 163.367
R1290 B.n364 B.n363 163.367
R1291 B.n365 B.n364 163.367
R1292 B.n365 B.n140 163.367
R1293 B.n369 B.n140 163.367
R1294 B.n370 B.n369 163.367
R1295 B.n371 B.n370 163.367
R1296 B.n371 B.n138 163.367
R1297 B.n375 B.n138 163.367
R1298 B.n376 B.n375 163.367
R1299 B.n377 B.n376 163.367
R1300 B.n377 B.n136 163.367
R1301 B.n381 B.n136 163.367
R1302 B.n382 B.n381 163.367
R1303 B.n383 B.n382 163.367
R1304 B.n383 B.n134 163.367
R1305 B.n387 B.n134 163.367
R1306 B.n388 B.n387 163.367
R1307 B.n389 B.n388 163.367
R1308 B.n389 B.n132 163.367
R1309 B.n393 B.n132 163.367
R1310 B.n394 B.n393 163.367
R1311 B.n395 B.n394 163.367
R1312 B.n395 B.n130 163.367
R1313 B.n399 B.n130 163.367
R1314 B.n400 B.n399 163.367
R1315 B.n401 B.n400 163.367
R1316 B.n563 B.n562 163.367
R1317 B.n562 B.n561 163.367
R1318 B.n561 B.n76 163.367
R1319 B.n557 B.n76 163.367
R1320 B.n557 B.n556 163.367
R1321 B.n556 B.n555 163.367
R1322 B.n555 B.n78 163.367
R1323 B.n551 B.n78 163.367
R1324 B.n551 B.n550 163.367
R1325 B.n550 B.n549 163.367
R1326 B.n549 B.n80 163.367
R1327 B.n545 B.n80 163.367
R1328 B.n545 B.n544 163.367
R1329 B.n544 B.n543 163.367
R1330 B.n543 B.n82 163.367
R1331 B.n539 B.n82 163.367
R1332 B.n539 B.n538 163.367
R1333 B.n538 B.n537 163.367
R1334 B.n537 B.n84 163.367
R1335 B.n533 B.n84 163.367
R1336 B.n533 B.n532 163.367
R1337 B.n532 B.n531 163.367
R1338 B.n531 B.n86 163.367
R1339 B.n527 B.n86 163.367
R1340 B.n527 B.n526 163.367
R1341 B.n526 B.n525 163.367
R1342 B.n525 B.n88 163.367
R1343 B.n521 B.n88 163.367
R1344 B.n521 B.n520 163.367
R1345 B.n520 B.n519 163.367
R1346 B.n519 B.n90 163.367
R1347 B.n515 B.n90 163.367
R1348 B.n515 B.n514 163.367
R1349 B.n514 B.n513 163.367
R1350 B.n513 B.n92 163.367
R1351 B.n509 B.n92 163.367
R1352 B.n509 B.n508 163.367
R1353 B.n508 B.n507 163.367
R1354 B.n507 B.n94 163.367
R1355 B.n503 B.n94 163.367
R1356 B.n503 B.n502 163.367
R1357 B.n502 B.n501 163.367
R1358 B.n501 B.n96 163.367
R1359 B.n497 B.n96 163.367
R1360 B.n497 B.n496 163.367
R1361 B.n496 B.n495 163.367
R1362 B.n495 B.n98 163.367
R1363 B.n491 B.n98 163.367
R1364 B.n491 B.n490 163.367
R1365 B.n490 B.n489 163.367
R1366 B.n489 B.n100 163.367
R1367 B.n485 B.n100 163.367
R1368 B.n485 B.n484 163.367
R1369 B.n484 B.n483 163.367
R1370 B.n483 B.n102 163.367
R1371 B.n479 B.n102 163.367
R1372 B.n479 B.n478 163.367
R1373 B.n478 B.n477 163.367
R1374 B.n477 B.n104 163.367
R1375 B.n473 B.n104 163.367
R1376 B.n473 B.n472 163.367
R1377 B.n472 B.n471 163.367
R1378 B.n471 B.n106 163.367
R1379 B.n467 B.n106 163.367
R1380 B.n467 B.n466 163.367
R1381 B.n466 B.n465 163.367
R1382 B.n465 B.n108 163.367
R1383 B.n461 B.n108 163.367
R1384 B.n461 B.n460 163.367
R1385 B.n460 B.n459 163.367
R1386 B.n459 B.n110 163.367
R1387 B.n455 B.n110 163.367
R1388 B.n455 B.n454 163.367
R1389 B.n454 B.n453 163.367
R1390 B.n453 B.n112 163.367
R1391 B.n449 B.n112 163.367
R1392 B.n449 B.n448 163.367
R1393 B.n448 B.n447 163.367
R1394 B.n447 B.n114 163.367
R1395 B.n443 B.n114 163.367
R1396 B.n443 B.n442 163.367
R1397 B.n442 B.n441 163.367
R1398 B.n441 B.n116 163.367
R1399 B.n437 B.n116 163.367
R1400 B.n437 B.n436 163.367
R1401 B.n436 B.n435 163.367
R1402 B.n435 B.n118 163.367
R1403 B.n431 B.n118 163.367
R1404 B.n431 B.n430 163.367
R1405 B.n430 B.n429 163.367
R1406 B.n429 B.n120 163.367
R1407 B.n425 B.n120 163.367
R1408 B.n425 B.n424 163.367
R1409 B.n424 B.n423 163.367
R1410 B.n423 B.n122 163.367
R1411 B.n419 B.n122 163.367
R1412 B.n419 B.n418 163.367
R1413 B.n418 B.n417 163.367
R1414 B.n417 B.n124 163.367
R1415 B.n413 B.n124 163.367
R1416 B.n413 B.n412 163.367
R1417 B.n412 B.n411 163.367
R1418 B.n411 B.n126 163.367
R1419 B.n407 B.n126 163.367
R1420 B.n407 B.n406 163.367
R1421 B.n406 B.n405 163.367
R1422 B.n405 B.n128 163.367
R1423 B.n688 B.n29 163.367
R1424 B.n684 B.n29 163.367
R1425 B.n684 B.n683 163.367
R1426 B.n683 B.n682 163.367
R1427 B.n682 B.n31 163.367
R1428 B.n678 B.n31 163.367
R1429 B.n678 B.n677 163.367
R1430 B.n677 B.n676 163.367
R1431 B.n676 B.n33 163.367
R1432 B.n672 B.n33 163.367
R1433 B.n672 B.n671 163.367
R1434 B.n671 B.n670 163.367
R1435 B.n670 B.n35 163.367
R1436 B.n666 B.n35 163.367
R1437 B.n666 B.n665 163.367
R1438 B.n665 B.n664 163.367
R1439 B.n664 B.n37 163.367
R1440 B.n660 B.n37 163.367
R1441 B.n660 B.n659 163.367
R1442 B.n659 B.n658 163.367
R1443 B.n658 B.n39 163.367
R1444 B.n654 B.n39 163.367
R1445 B.n654 B.n653 163.367
R1446 B.n653 B.n652 163.367
R1447 B.n652 B.n41 163.367
R1448 B.n648 B.n41 163.367
R1449 B.n648 B.n647 163.367
R1450 B.n647 B.n646 163.367
R1451 B.n646 B.n43 163.367
R1452 B.n642 B.n43 163.367
R1453 B.n642 B.n641 163.367
R1454 B.n641 B.n640 163.367
R1455 B.n640 B.n45 163.367
R1456 B.n636 B.n45 163.367
R1457 B.n636 B.n635 163.367
R1458 B.n635 B.n634 163.367
R1459 B.n634 B.n47 163.367
R1460 B.n630 B.n47 163.367
R1461 B.n630 B.n629 163.367
R1462 B.n629 B.n628 163.367
R1463 B.n628 B.n52 163.367
R1464 B.n624 B.n52 163.367
R1465 B.n624 B.n623 163.367
R1466 B.n623 B.n622 163.367
R1467 B.n622 B.n54 163.367
R1468 B.n617 B.n54 163.367
R1469 B.n617 B.n616 163.367
R1470 B.n616 B.n615 163.367
R1471 B.n615 B.n58 163.367
R1472 B.n611 B.n58 163.367
R1473 B.n611 B.n610 163.367
R1474 B.n610 B.n609 163.367
R1475 B.n609 B.n60 163.367
R1476 B.n605 B.n60 163.367
R1477 B.n605 B.n604 163.367
R1478 B.n604 B.n603 163.367
R1479 B.n603 B.n62 163.367
R1480 B.n599 B.n62 163.367
R1481 B.n599 B.n598 163.367
R1482 B.n598 B.n597 163.367
R1483 B.n597 B.n64 163.367
R1484 B.n593 B.n64 163.367
R1485 B.n593 B.n592 163.367
R1486 B.n592 B.n591 163.367
R1487 B.n591 B.n66 163.367
R1488 B.n587 B.n66 163.367
R1489 B.n587 B.n586 163.367
R1490 B.n586 B.n585 163.367
R1491 B.n585 B.n68 163.367
R1492 B.n581 B.n68 163.367
R1493 B.n581 B.n580 163.367
R1494 B.n580 B.n579 163.367
R1495 B.n579 B.n70 163.367
R1496 B.n575 B.n70 163.367
R1497 B.n575 B.n574 163.367
R1498 B.n574 B.n573 163.367
R1499 B.n573 B.n72 163.367
R1500 B.n569 B.n72 163.367
R1501 B.n569 B.n568 163.367
R1502 B.n568 B.n567 163.367
R1503 B.n567 B.n74 163.367
R1504 B.n690 B.n689 163.367
R1505 B.n690 B.n27 163.367
R1506 B.n694 B.n27 163.367
R1507 B.n695 B.n694 163.367
R1508 B.n696 B.n695 163.367
R1509 B.n696 B.n25 163.367
R1510 B.n700 B.n25 163.367
R1511 B.n701 B.n700 163.367
R1512 B.n702 B.n701 163.367
R1513 B.n702 B.n23 163.367
R1514 B.n706 B.n23 163.367
R1515 B.n707 B.n706 163.367
R1516 B.n708 B.n707 163.367
R1517 B.n708 B.n21 163.367
R1518 B.n712 B.n21 163.367
R1519 B.n713 B.n712 163.367
R1520 B.n714 B.n713 163.367
R1521 B.n714 B.n19 163.367
R1522 B.n718 B.n19 163.367
R1523 B.n719 B.n718 163.367
R1524 B.n720 B.n719 163.367
R1525 B.n720 B.n17 163.367
R1526 B.n724 B.n17 163.367
R1527 B.n725 B.n724 163.367
R1528 B.n726 B.n725 163.367
R1529 B.n726 B.n15 163.367
R1530 B.n730 B.n15 163.367
R1531 B.n731 B.n730 163.367
R1532 B.n732 B.n731 163.367
R1533 B.n732 B.n13 163.367
R1534 B.n736 B.n13 163.367
R1535 B.n737 B.n736 163.367
R1536 B.n738 B.n737 163.367
R1537 B.n738 B.n11 163.367
R1538 B.n742 B.n11 163.367
R1539 B.n743 B.n742 163.367
R1540 B.n744 B.n743 163.367
R1541 B.n744 B.n9 163.367
R1542 B.n748 B.n9 163.367
R1543 B.n749 B.n748 163.367
R1544 B.n750 B.n749 163.367
R1545 B.n750 B.n7 163.367
R1546 B.n754 B.n7 163.367
R1547 B.n755 B.n754 163.367
R1548 B.n756 B.n755 163.367
R1549 B.n756 B.n5 163.367
R1550 B.n760 B.n5 163.367
R1551 B.n761 B.n760 163.367
R1552 B.n762 B.n761 163.367
R1553 B.n762 B.n3 163.367
R1554 B.n766 B.n3 163.367
R1555 B.n767 B.n766 163.367
R1556 B.n198 B.n2 163.367
R1557 B.n199 B.n198 163.367
R1558 B.n199 B.n196 163.367
R1559 B.n203 B.n196 163.367
R1560 B.n204 B.n203 163.367
R1561 B.n205 B.n204 163.367
R1562 B.n205 B.n194 163.367
R1563 B.n209 B.n194 163.367
R1564 B.n210 B.n209 163.367
R1565 B.n211 B.n210 163.367
R1566 B.n211 B.n192 163.367
R1567 B.n215 B.n192 163.367
R1568 B.n216 B.n215 163.367
R1569 B.n217 B.n216 163.367
R1570 B.n217 B.n190 163.367
R1571 B.n221 B.n190 163.367
R1572 B.n222 B.n221 163.367
R1573 B.n223 B.n222 163.367
R1574 B.n223 B.n188 163.367
R1575 B.n227 B.n188 163.367
R1576 B.n228 B.n227 163.367
R1577 B.n229 B.n228 163.367
R1578 B.n229 B.n186 163.367
R1579 B.n233 B.n186 163.367
R1580 B.n234 B.n233 163.367
R1581 B.n235 B.n234 163.367
R1582 B.n235 B.n184 163.367
R1583 B.n239 B.n184 163.367
R1584 B.n240 B.n239 163.367
R1585 B.n241 B.n240 163.367
R1586 B.n241 B.n182 163.367
R1587 B.n245 B.n182 163.367
R1588 B.n246 B.n245 163.367
R1589 B.n247 B.n246 163.367
R1590 B.n247 B.n180 163.367
R1591 B.n251 B.n180 163.367
R1592 B.n252 B.n251 163.367
R1593 B.n253 B.n252 163.367
R1594 B.n253 B.n178 163.367
R1595 B.n257 B.n178 163.367
R1596 B.n258 B.n257 163.367
R1597 B.n259 B.n258 163.367
R1598 B.n259 B.n176 163.367
R1599 B.n263 B.n176 163.367
R1600 B.n264 B.n263 163.367
R1601 B.n265 B.n264 163.367
R1602 B.n265 B.n174 163.367
R1603 B.n269 B.n174 163.367
R1604 B.n270 B.n269 163.367
R1605 B.n271 B.n270 163.367
R1606 B.n271 B.n172 163.367
R1607 B.n275 B.n172 163.367
R1608 B.n329 B.n328 75.249
R1609 B.n148 B.n147 75.249
R1610 B.n56 B.n55 75.249
R1611 B.n49 B.n48 75.249
R1612 B.n330 B.n329 59.5399
R1613 B.n348 B.n148 59.5399
R1614 B.n619 B.n56 59.5399
R1615 B.n50 B.n49 59.5399
R1616 B.n687 B.n28 33.2493
R1617 B.n565 B.n564 33.2493
R1618 B.n403 B.n402 33.2493
R1619 B.n274 B.n171 33.2493
R1620 B B.n769 18.0485
R1621 B.n691 B.n28 10.6151
R1622 B.n692 B.n691 10.6151
R1623 B.n693 B.n692 10.6151
R1624 B.n693 B.n26 10.6151
R1625 B.n697 B.n26 10.6151
R1626 B.n698 B.n697 10.6151
R1627 B.n699 B.n698 10.6151
R1628 B.n699 B.n24 10.6151
R1629 B.n703 B.n24 10.6151
R1630 B.n704 B.n703 10.6151
R1631 B.n705 B.n704 10.6151
R1632 B.n705 B.n22 10.6151
R1633 B.n709 B.n22 10.6151
R1634 B.n710 B.n709 10.6151
R1635 B.n711 B.n710 10.6151
R1636 B.n711 B.n20 10.6151
R1637 B.n715 B.n20 10.6151
R1638 B.n716 B.n715 10.6151
R1639 B.n717 B.n716 10.6151
R1640 B.n717 B.n18 10.6151
R1641 B.n721 B.n18 10.6151
R1642 B.n722 B.n721 10.6151
R1643 B.n723 B.n722 10.6151
R1644 B.n723 B.n16 10.6151
R1645 B.n727 B.n16 10.6151
R1646 B.n728 B.n727 10.6151
R1647 B.n729 B.n728 10.6151
R1648 B.n729 B.n14 10.6151
R1649 B.n733 B.n14 10.6151
R1650 B.n734 B.n733 10.6151
R1651 B.n735 B.n734 10.6151
R1652 B.n735 B.n12 10.6151
R1653 B.n739 B.n12 10.6151
R1654 B.n740 B.n739 10.6151
R1655 B.n741 B.n740 10.6151
R1656 B.n741 B.n10 10.6151
R1657 B.n745 B.n10 10.6151
R1658 B.n746 B.n745 10.6151
R1659 B.n747 B.n746 10.6151
R1660 B.n747 B.n8 10.6151
R1661 B.n751 B.n8 10.6151
R1662 B.n752 B.n751 10.6151
R1663 B.n753 B.n752 10.6151
R1664 B.n753 B.n6 10.6151
R1665 B.n757 B.n6 10.6151
R1666 B.n758 B.n757 10.6151
R1667 B.n759 B.n758 10.6151
R1668 B.n759 B.n4 10.6151
R1669 B.n763 B.n4 10.6151
R1670 B.n764 B.n763 10.6151
R1671 B.n765 B.n764 10.6151
R1672 B.n765 B.n0 10.6151
R1673 B.n687 B.n686 10.6151
R1674 B.n686 B.n685 10.6151
R1675 B.n685 B.n30 10.6151
R1676 B.n681 B.n30 10.6151
R1677 B.n681 B.n680 10.6151
R1678 B.n680 B.n679 10.6151
R1679 B.n679 B.n32 10.6151
R1680 B.n675 B.n32 10.6151
R1681 B.n675 B.n674 10.6151
R1682 B.n674 B.n673 10.6151
R1683 B.n673 B.n34 10.6151
R1684 B.n669 B.n34 10.6151
R1685 B.n669 B.n668 10.6151
R1686 B.n668 B.n667 10.6151
R1687 B.n667 B.n36 10.6151
R1688 B.n663 B.n36 10.6151
R1689 B.n663 B.n662 10.6151
R1690 B.n662 B.n661 10.6151
R1691 B.n661 B.n38 10.6151
R1692 B.n657 B.n38 10.6151
R1693 B.n657 B.n656 10.6151
R1694 B.n656 B.n655 10.6151
R1695 B.n655 B.n40 10.6151
R1696 B.n651 B.n40 10.6151
R1697 B.n651 B.n650 10.6151
R1698 B.n650 B.n649 10.6151
R1699 B.n649 B.n42 10.6151
R1700 B.n645 B.n42 10.6151
R1701 B.n645 B.n644 10.6151
R1702 B.n644 B.n643 10.6151
R1703 B.n643 B.n44 10.6151
R1704 B.n639 B.n44 10.6151
R1705 B.n639 B.n638 10.6151
R1706 B.n638 B.n637 10.6151
R1707 B.n637 B.n46 10.6151
R1708 B.n633 B.n632 10.6151
R1709 B.n632 B.n631 10.6151
R1710 B.n631 B.n51 10.6151
R1711 B.n627 B.n51 10.6151
R1712 B.n627 B.n626 10.6151
R1713 B.n626 B.n625 10.6151
R1714 B.n625 B.n53 10.6151
R1715 B.n621 B.n53 10.6151
R1716 B.n621 B.n620 10.6151
R1717 B.n618 B.n57 10.6151
R1718 B.n614 B.n57 10.6151
R1719 B.n614 B.n613 10.6151
R1720 B.n613 B.n612 10.6151
R1721 B.n612 B.n59 10.6151
R1722 B.n608 B.n59 10.6151
R1723 B.n608 B.n607 10.6151
R1724 B.n607 B.n606 10.6151
R1725 B.n606 B.n61 10.6151
R1726 B.n602 B.n61 10.6151
R1727 B.n602 B.n601 10.6151
R1728 B.n601 B.n600 10.6151
R1729 B.n600 B.n63 10.6151
R1730 B.n596 B.n63 10.6151
R1731 B.n596 B.n595 10.6151
R1732 B.n595 B.n594 10.6151
R1733 B.n594 B.n65 10.6151
R1734 B.n590 B.n65 10.6151
R1735 B.n590 B.n589 10.6151
R1736 B.n589 B.n588 10.6151
R1737 B.n588 B.n67 10.6151
R1738 B.n584 B.n67 10.6151
R1739 B.n584 B.n583 10.6151
R1740 B.n583 B.n582 10.6151
R1741 B.n582 B.n69 10.6151
R1742 B.n578 B.n69 10.6151
R1743 B.n578 B.n577 10.6151
R1744 B.n577 B.n576 10.6151
R1745 B.n576 B.n71 10.6151
R1746 B.n572 B.n71 10.6151
R1747 B.n572 B.n571 10.6151
R1748 B.n571 B.n570 10.6151
R1749 B.n570 B.n73 10.6151
R1750 B.n566 B.n73 10.6151
R1751 B.n566 B.n565 10.6151
R1752 B.n564 B.n75 10.6151
R1753 B.n560 B.n75 10.6151
R1754 B.n560 B.n559 10.6151
R1755 B.n559 B.n558 10.6151
R1756 B.n558 B.n77 10.6151
R1757 B.n554 B.n77 10.6151
R1758 B.n554 B.n553 10.6151
R1759 B.n553 B.n552 10.6151
R1760 B.n552 B.n79 10.6151
R1761 B.n548 B.n79 10.6151
R1762 B.n548 B.n547 10.6151
R1763 B.n547 B.n546 10.6151
R1764 B.n546 B.n81 10.6151
R1765 B.n542 B.n81 10.6151
R1766 B.n542 B.n541 10.6151
R1767 B.n541 B.n540 10.6151
R1768 B.n540 B.n83 10.6151
R1769 B.n536 B.n83 10.6151
R1770 B.n536 B.n535 10.6151
R1771 B.n535 B.n534 10.6151
R1772 B.n534 B.n85 10.6151
R1773 B.n530 B.n85 10.6151
R1774 B.n530 B.n529 10.6151
R1775 B.n529 B.n528 10.6151
R1776 B.n528 B.n87 10.6151
R1777 B.n524 B.n87 10.6151
R1778 B.n524 B.n523 10.6151
R1779 B.n523 B.n522 10.6151
R1780 B.n522 B.n89 10.6151
R1781 B.n518 B.n89 10.6151
R1782 B.n518 B.n517 10.6151
R1783 B.n517 B.n516 10.6151
R1784 B.n516 B.n91 10.6151
R1785 B.n512 B.n91 10.6151
R1786 B.n512 B.n511 10.6151
R1787 B.n511 B.n510 10.6151
R1788 B.n510 B.n93 10.6151
R1789 B.n506 B.n93 10.6151
R1790 B.n506 B.n505 10.6151
R1791 B.n505 B.n504 10.6151
R1792 B.n504 B.n95 10.6151
R1793 B.n500 B.n95 10.6151
R1794 B.n500 B.n499 10.6151
R1795 B.n499 B.n498 10.6151
R1796 B.n498 B.n97 10.6151
R1797 B.n494 B.n97 10.6151
R1798 B.n494 B.n493 10.6151
R1799 B.n493 B.n492 10.6151
R1800 B.n492 B.n99 10.6151
R1801 B.n488 B.n99 10.6151
R1802 B.n488 B.n487 10.6151
R1803 B.n487 B.n486 10.6151
R1804 B.n486 B.n101 10.6151
R1805 B.n482 B.n101 10.6151
R1806 B.n482 B.n481 10.6151
R1807 B.n481 B.n480 10.6151
R1808 B.n480 B.n103 10.6151
R1809 B.n476 B.n103 10.6151
R1810 B.n476 B.n475 10.6151
R1811 B.n475 B.n474 10.6151
R1812 B.n474 B.n105 10.6151
R1813 B.n470 B.n105 10.6151
R1814 B.n470 B.n469 10.6151
R1815 B.n469 B.n468 10.6151
R1816 B.n468 B.n107 10.6151
R1817 B.n464 B.n107 10.6151
R1818 B.n464 B.n463 10.6151
R1819 B.n463 B.n462 10.6151
R1820 B.n462 B.n109 10.6151
R1821 B.n458 B.n109 10.6151
R1822 B.n458 B.n457 10.6151
R1823 B.n457 B.n456 10.6151
R1824 B.n456 B.n111 10.6151
R1825 B.n452 B.n111 10.6151
R1826 B.n452 B.n451 10.6151
R1827 B.n451 B.n450 10.6151
R1828 B.n450 B.n113 10.6151
R1829 B.n446 B.n113 10.6151
R1830 B.n446 B.n445 10.6151
R1831 B.n445 B.n444 10.6151
R1832 B.n444 B.n115 10.6151
R1833 B.n440 B.n115 10.6151
R1834 B.n440 B.n439 10.6151
R1835 B.n439 B.n438 10.6151
R1836 B.n438 B.n117 10.6151
R1837 B.n434 B.n117 10.6151
R1838 B.n434 B.n433 10.6151
R1839 B.n433 B.n432 10.6151
R1840 B.n432 B.n119 10.6151
R1841 B.n428 B.n119 10.6151
R1842 B.n428 B.n427 10.6151
R1843 B.n427 B.n426 10.6151
R1844 B.n426 B.n121 10.6151
R1845 B.n422 B.n121 10.6151
R1846 B.n422 B.n421 10.6151
R1847 B.n421 B.n420 10.6151
R1848 B.n420 B.n123 10.6151
R1849 B.n416 B.n123 10.6151
R1850 B.n416 B.n415 10.6151
R1851 B.n415 B.n414 10.6151
R1852 B.n414 B.n125 10.6151
R1853 B.n410 B.n125 10.6151
R1854 B.n410 B.n409 10.6151
R1855 B.n409 B.n408 10.6151
R1856 B.n408 B.n127 10.6151
R1857 B.n404 B.n127 10.6151
R1858 B.n404 B.n403 10.6151
R1859 B.n197 B.n1 10.6151
R1860 B.n200 B.n197 10.6151
R1861 B.n201 B.n200 10.6151
R1862 B.n202 B.n201 10.6151
R1863 B.n202 B.n195 10.6151
R1864 B.n206 B.n195 10.6151
R1865 B.n207 B.n206 10.6151
R1866 B.n208 B.n207 10.6151
R1867 B.n208 B.n193 10.6151
R1868 B.n212 B.n193 10.6151
R1869 B.n213 B.n212 10.6151
R1870 B.n214 B.n213 10.6151
R1871 B.n214 B.n191 10.6151
R1872 B.n218 B.n191 10.6151
R1873 B.n219 B.n218 10.6151
R1874 B.n220 B.n219 10.6151
R1875 B.n220 B.n189 10.6151
R1876 B.n224 B.n189 10.6151
R1877 B.n225 B.n224 10.6151
R1878 B.n226 B.n225 10.6151
R1879 B.n226 B.n187 10.6151
R1880 B.n230 B.n187 10.6151
R1881 B.n231 B.n230 10.6151
R1882 B.n232 B.n231 10.6151
R1883 B.n232 B.n185 10.6151
R1884 B.n236 B.n185 10.6151
R1885 B.n237 B.n236 10.6151
R1886 B.n238 B.n237 10.6151
R1887 B.n238 B.n183 10.6151
R1888 B.n242 B.n183 10.6151
R1889 B.n243 B.n242 10.6151
R1890 B.n244 B.n243 10.6151
R1891 B.n244 B.n181 10.6151
R1892 B.n248 B.n181 10.6151
R1893 B.n249 B.n248 10.6151
R1894 B.n250 B.n249 10.6151
R1895 B.n250 B.n179 10.6151
R1896 B.n254 B.n179 10.6151
R1897 B.n255 B.n254 10.6151
R1898 B.n256 B.n255 10.6151
R1899 B.n256 B.n177 10.6151
R1900 B.n260 B.n177 10.6151
R1901 B.n261 B.n260 10.6151
R1902 B.n262 B.n261 10.6151
R1903 B.n262 B.n175 10.6151
R1904 B.n266 B.n175 10.6151
R1905 B.n267 B.n266 10.6151
R1906 B.n268 B.n267 10.6151
R1907 B.n268 B.n173 10.6151
R1908 B.n272 B.n173 10.6151
R1909 B.n273 B.n272 10.6151
R1910 B.n274 B.n273 10.6151
R1911 B.n278 B.n171 10.6151
R1912 B.n279 B.n278 10.6151
R1913 B.n280 B.n279 10.6151
R1914 B.n280 B.n169 10.6151
R1915 B.n284 B.n169 10.6151
R1916 B.n285 B.n284 10.6151
R1917 B.n286 B.n285 10.6151
R1918 B.n286 B.n167 10.6151
R1919 B.n290 B.n167 10.6151
R1920 B.n291 B.n290 10.6151
R1921 B.n292 B.n291 10.6151
R1922 B.n292 B.n165 10.6151
R1923 B.n296 B.n165 10.6151
R1924 B.n297 B.n296 10.6151
R1925 B.n298 B.n297 10.6151
R1926 B.n298 B.n163 10.6151
R1927 B.n302 B.n163 10.6151
R1928 B.n303 B.n302 10.6151
R1929 B.n304 B.n303 10.6151
R1930 B.n304 B.n161 10.6151
R1931 B.n308 B.n161 10.6151
R1932 B.n309 B.n308 10.6151
R1933 B.n310 B.n309 10.6151
R1934 B.n310 B.n159 10.6151
R1935 B.n314 B.n159 10.6151
R1936 B.n315 B.n314 10.6151
R1937 B.n316 B.n315 10.6151
R1938 B.n316 B.n157 10.6151
R1939 B.n320 B.n157 10.6151
R1940 B.n321 B.n320 10.6151
R1941 B.n322 B.n321 10.6151
R1942 B.n322 B.n155 10.6151
R1943 B.n326 B.n155 10.6151
R1944 B.n327 B.n326 10.6151
R1945 B.n331 B.n327 10.6151
R1946 B.n335 B.n153 10.6151
R1947 B.n336 B.n335 10.6151
R1948 B.n337 B.n336 10.6151
R1949 B.n337 B.n151 10.6151
R1950 B.n341 B.n151 10.6151
R1951 B.n342 B.n341 10.6151
R1952 B.n343 B.n342 10.6151
R1953 B.n343 B.n149 10.6151
R1954 B.n347 B.n149 10.6151
R1955 B.n350 B.n349 10.6151
R1956 B.n350 B.n145 10.6151
R1957 B.n354 B.n145 10.6151
R1958 B.n355 B.n354 10.6151
R1959 B.n356 B.n355 10.6151
R1960 B.n356 B.n143 10.6151
R1961 B.n360 B.n143 10.6151
R1962 B.n361 B.n360 10.6151
R1963 B.n362 B.n361 10.6151
R1964 B.n362 B.n141 10.6151
R1965 B.n366 B.n141 10.6151
R1966 B.n367 B.n366 10.6151
R1967 B.n368 B.n367 10.6151
R1968 B.n368 B.n139 10.6151
R1969 B.n372 B.n139 10.6151
R1970 B.n373 B.n372 10.6151
R1971 B.n374 B.n373 10.6151
R1972 B.n374 B.n137 10.6151
R1973 B.n378 B.n137 10.6151
R1974 B.n379 B.n378 10.6151
R1975 B.n380 B.n379 10.6151
R1976 B.n380 B.n135 10.6151
R1977 B.n384 B.n135 10.6151
R1978 B.n385 B.n384 10.6151
R1979 B.n386 B.n385 10.6151
R1980 B.n386 B.n133 10.6151
R1981 B.n390 B.n133 10.6151
R1982 B.n391 B.n390 10.6151
R1983 B.n392 B.n391 10.6151
R1984 B.n392 B.n131 10.6151
R1985 B.n396 B.n131 10.6151
R1986 B.n397 B.n396 10.6151
R1987 B.n398 B.n397 10.6151
R1988 B.n398 B.n129 10.6151
R1989 B.n402 B.n129 10.6151
R1990 B.n50 B.n46 9.36635
R1991 B.n619 B.n618 9.36635
R1992 B.n331 B.n330 9.36635
R1993 B.n349 B.n348 9.36635
R1994 B.n769 B.n0 8.11757
R1995 B.n769 B.n1 8.11757
R1996 B.n633 B.n50 1.24928
R1997 B.n620 B.n619 1.24928
R1998 B.n330 B.n153 1.24928
R1999 B.n348 B.n347 1.24928
C0 B VDD1 2.18741f
C1 VTAIL VDD1 7.42616f
C2 VDD1 VN 0.152466f
C3 VTAIL B 3.60208f
C4 VDD2 VDD1 1.77815f
C5 B VN 1.34993f
C6 VTAIL VN 6.49729f
C7 B VDD2 2.28429f
C8 VTAIL VDD2 7.48449f
C9 VDD2 VN 6.01928f
C10 w_n4074_n2988# VP 8.43442f
C11 VDD1 VP 6.40321f
C12 B VP 2.23854f
C13 VTAIL VP 6.5115f
C14 w_n4074_n2988# VDD1 2.39332f
C15 VN VP 7.49465f
C16 B w_n4074_n2988# 10.455501f
C17 VTAIL w_n4074_n2988# 2.8042f
C18 VDD2 VP 0.539195f
C19 w_n4074_n2988# VN 7.90506f
C20 w_n4074_n2988# VDD2 2.50876f
C21 VDD2 VSUBS 2.106369f
C22 VDD1 VSUBS 2.118851f
C23 VTAIL VSUBS 1.307973f
C24 VN VSUBS 6.72858f
C25 VP VSUBS 3.606997f
C26 B VSUBS 5.416051f
C27 w_n4074_n2988# VSUBS 0.150331p
C28 B.n0 VSUBS 0.008012f
C29 B.n1 VSUBS 0.008012f
C30 B.n2 VSUBS 0.01185f
C31 B.n3 VSUBS 0.009081f
C32 B.n4 VSUBS 0.009081f
C33 B.n5 VSUBS 0.009081f
C34 B.n6 VSUBS 0.009081f
C35 B.n7 VSUBS 0.009081f
C36 B.n8 VSUBS 0.009081f
C37 B.n9 VSUBS 0.009081f
C38 B.n10 VSUBS 0.009081f
C39 B.n11 VSUBS 0.009081f
C40 B.n12 VSUBS 0.009081f
C41 B.n13 VSUBS 0.009081f
C42 B.n14 VSUBS 0.009081f
C43 B.n15 VSUBS 0.009081f
C44 B.n16 VSUBS 0.009081f
C45 B.n17 VSUBS 0.009081f
C46 B.n18 VSUBS 0.009081f
C47 B.n19 VSUBS 0.009081f
C48 B.n20 VSUBS 0.009081f
C49 B.n21 VSUBS 0.009081f
C50 B.n22 VSUBS 0.009081f
C51 B.n23 VSUBS 0.009081f
C52 B.n24 VSUBS 0.009081f
C53 B.n25 VSUBS 0.009081f
C54 B.n26 VSUBS 0.009081f
C55 B.n27 VSUBS 0.009081f
C56 B.n28 VSUBS 0.020613f
C57 B.n29 VSUBS 0.009081f
C58 B.n30 VSUBS 0.009081f
C59 B.n31 VSUBS 0.009081f
C60 B.n32 VSUBS 0.009081f
C61 B.n33 VSUBS 0.009081f
C62 B.n34 VSUBS 0.009081f
C63 B.n35 VSUBS 0.009081f
C64 B.n36 VSUBS 0.009081f
C65 B.n37 VSUBS 0.009081f
C66 B.n38 VSUBS 0.009081f
C67 B.n39 VSUBS 0.009081f
C68 B.n40 VSUBS 0.009081f
C69 B.n41 VSUBS 0.009081f
C70 B.n42 VSUBS 0.009081f
C71 B.n43 VSUBS 0.009081f
C72 B.n44 VSUBS 0.009081f
C73 B.n45 VSUBS 0.009081f
C74 B.n46 VSUBS 0.008547f
C75 B.n47 VSUBS 0.009081f
C76 B.t4 VSUBS 0.22024f
C77 B.t5 VSUBS 0.271382f
C78 B.t3 VSUBS 2.18026f
C79 B.n48 VSUBS 0.436313f
C80 B.n49 VSUBS 0.296199f
C81 B.n50 VSUBS 0.021039f
C82 B.n51 VSUBS 0.009081f
C83 B.n52 VSUBS 0.009081f
C84 B.n53 VSUBS 0.009081f
C85 B.n54 VSUBS 0.009081f
C86 B.t7 VSUBS 0.220244f
C87 B.t8 VSUBS 0.271385f
C88 B.t6 VSUBS 2.18026f
C89 B.n55 VSUBS 0.43631f
C90 B.n56 VSUBS 0.296195f
C91 B.n57 VSUBS 0.009081f
C92 B.n58 VSUBS 0.009081f
C93 B.n59 VSUBS 0.009081f
C94 B.n60 VSUBS 0.009081f
C95 B.n61 VSUBS 0.009081f
C96 B.n62 VSUBS 0.009081f
C97 B.n63 VSUBS 0.009081f
C98 B.n64 VSUBS 0.009081f
C99 B.n65 VSUBS 0.009081f
C100 B.n66 VSUBS 0.009081f
C101 B.n67 VSUBS 0.009081f
C102 B.n68 VSUBS 0.009081f
C103 B.n69 VSUBS 0.009081f
C104 B.n70 VSUBS 0.009081f
C105 B.n71 VSUBS 0.009081f
C106 B.n72 VSUBS 0.009081f
C107 B.n73 VSUBS 0.009081f
C108 B.n74 VSUBS 0.022387f
C109 B.n75 VSUBS 0.009081f
C110 B.n76 VSUBS 0.009081f
C111 B.n77 VSUBS 0.009081f
C112 B.n78 VSUBS 0.009081f
C113 B.n79 VSUBS 0.009081f
C114 B.n80 VSUBS 0.009081f
C115 B.n81 VSUBS 0.009081f
C116 B.n82 VSUBS 0.009081f
C117 B.n83 VSUBS 0.009081f
C118 B.n84 VSUBS 0.009081f
C119 B.n85 VSUBS 0.009081f
C120 B.n86 VSUBS 0.009081f
C121 B.n87 VSUBS 0.009081f
C122 B.n88 VSUBS 0.009081f
C123 B.n89 VSUBS 0.009081f
C124 B.n90 VSUBS 0.009081f
C125 B.n91 VSUBS 0.009081f
C126 B.n92 VSUBS 0.009081f
C127 B.n93 VSUBS 0.009081f
C128 B.n94 VSUBS 0.009081f
C129 B.n95 VSUBS 0.009081f
C130 B.n96 VSUBS 0.009081f
C131 B.n97 VSUBS 0.009081f
C132 B.n98 VSUBS 0.009081f
C133 B.n99 VSUBS 0.009081f
C134 B.n100 VSUBS 0.009081f
C135 B.n101 VSUBS 0.009081f
C136 B.n102 VSUBS 0.009081f
C137 B.n103 VSUBS 0.009081f
C138 B.n104 VSUBS 0.009081f
C139 B.n105 VSUBS 0.009081f
C140 B.n106 VSUBS 0.009081f
C141 B.n107 VSUBS 0.009081f
C142 B.n108 VSUBS 0.009081f
C143 B.n109 VSUBS 0.009081f
C144 B.n110 VSUBS 0.009081f
C145 B.n111 VSUBS 0.009081f
C146 B.n112 VSUBS 0.009081f
C147 B.n113 VSUBS 0.009081f
C148 B.n114 VSUBS 0.009081f
C149 B.n115 VSUBS 0.009081f
C150 B.n116 VSUBS 0.009081f
C151 B.n117 VSUBS 0.009081f
C152 B.n118 VSUBS 0.009081f
C153 B.n119 VSUBS 0.009081f
C154 B.n120 VSUBS 0.009081f
C155 B.n121 VSUBS 0.009081f
C156 B.n122 VSUBS 0.009081f
C157 B.n123 VSUBS 0.009081f
C158 B.n124 VSUBS 0.009081f
C159 B.n125 VSUBS 0.009081f
C160 B.n126 VSUBS 0.009081f
C161 B.n127 VSUBS 0.009081f
C162 B.n128 VSUBS 0.020613f
C163 B.n129 VSUBS 0.009081f
C164 B.n130 VSUBS 0.009081f
C165 B.n131 VSUBS 0.009081f
C166 B.n132 VSUBS 0.009081f
C167 B.n133 VSUBS 0.009081f
C168 B.n134 VSUBS 0.009081f
C169 B.n135 VSUBS 0.009081f
C170 B.n136 VSUBS 0.009081f
C171 B.n137 VSUBS 0.009081f
C172 B.n138 VSUBS 0.009081f
C173 B.n139 VSUBS 0.009081f
C174 B.n140 VSUBS 0.009081f
C175 B.n141 VSUBS 0.009081f
C176 B.n142 VSUBS 0.009081f
C177 B.n143 VSUBS 0.009081f
C178 B.n144 VSUBS 0.009081f
C179 B.n145 VSUBS 0.009081f
C180 B.n146 VSUBS 0.009081f
C181 B.t11 VSUBS 0.220244f
C182 B.t10 VSUBS 0.271385f
C183 B.t9 VSUBS 2.18026f
C184 B.n147 VSUBS 0.43631f
C185 B.n148 VSUBS 0.296195f
C186 B.n149 VSUBS 0.009081f
C187 B.n150 VSUBS 0.009081f
C188 B.n151 VSUBS 0.009081f
C189 B.n152 VSUBS 0.009081f
C190 B.n153 VSUBS 0.005075f
C191 B.n154 VSUBS 0.009081f
C192 B.n155 VSUBS 0.009081f
C193 B.n156 VSUBS 0.009081f
C194 B.n157 VSUBS 0.009081f
C195 B.n158 VSUBS 0.009081f
C196 B.n159 VSUBS 0.009081f
C197 B.n160 VSUBS 0.009081f
C198 B.n161 VSUBS 0.009081f
C199 B.n162 VSUBS 0.009081f
C200 B.n163 VSUBS 0.009081f
C201 B.n164 VSUBS 0.009081f
C202 B.n165 VSUBS 0.009081f
C203 B.n166 VSUBS 0.009081f
C204 B.n167 VSUBS 0.009081f
C205 B.n168 VSUBS 0.009081f
C206 B.n169 VSUBS 0.009081f
C207 B.n170 VSUBS 0.009081f
C208 B.n171 VSUBS 0.022387f
C209 B.n172 VSUBS 0.009081f
C210 B.n173 VSUBS 0.009081f
C211 B.n174 VSUBS 0.009081f
C212 B.n175 VSUBS 0.009081f
C213 B.n176 VSUBS 0.009081f
C214 B.n177 VSUBS 0.009081f
C215 B.n178 VSUBS 0.009081f
C216 B.n179 VSUBS 0.009081f
C217 B.n180 VSUBS 0.009081f
C218 B.n181 VSUBS 0.009081f
C219 B.n182 VSUBS 0.009081f
C220 B.n183 VSUBS 0.009081f
C221 B.n184 VSUBS 0.009081f
C222 B.n185 VSUBS 0.009081f
C223 B.n186 VSUBS 0.009081f
C224 B.n187 VSUBS 0.009081f
C225 B.n188 VSUBS 0.009081f
C226 B.n189 VSUBS 0.009081f
C227 B.n190 VSUBS 0.009081f
C228 B.n191 VSUBS 0.009081f
C229 B.n192 VSUBS 0.009081f
C230 B.n193 VSUBS 0.009081f
C231 B.n194 VSUBS 0.009081f
C232 B.n195 VSUBS 0.009081f
C233 B.n196 VSUBS 0.009081f
C234 B.n197 VSUBS 0.009081f
C235 B.n198 VSUBS 0.009081f
C236 B.n199 VSUBS 0.009081f
C237 B.n200 VSUBS 0.009081f
C238 B.n201 VSUBS 0.009081f
C239 B.n202 VSUBS 0.009081f
C240 B.n203 VSUBS 0.009081f
C241 B.n204 VSUBS 0.009081f
C242 B.n205 VSUBS 0.009081f
C243 B.n206 VSUBS 0.009081f
C244 B.n207 VSUBS 0.009081f
C245 B.n208 VSUBS 0.009081f
C246 B.n209 VSUBS 0.009081f
C247 B.n210 VSUBS 0.009081f
C248 B.n211 VSUBS 0.009081f
C249 B.n212 VSUBS 0.009081f
C250 B.n213 VSUBS 0.009081f
C251 B.n214 VSUBS 0.009081f
C252 B.n215 VSUBS 0.009081f
C253 B.n216 VSUBS 0.009081f
C254 B.n217 VSUBS 0.009081f
C255 B.n218 VSUBS 0.009081f
C256 B.n219 VSUBS 0.009081f
C257 B.n220 VSUBS 0.009081f
C258 B.n221 VSUBS 0.009081f
C259 B.n222 VSUBS 0.009081f
C260 B.n223 VSUBS 0.009081f
C261 B.n224 VSUBS 0.009081f
C262 B.n225 VSUBS 0.009081f
C263 B.n226 VSUBS 0.009081f
C264 B.n227 VSUBS 0.009081f
C265 B.n228 VSUBS 0.009081f
C266 B.n229 VSUBS 0.009081f
C267 B.n230 VSUBS 0.009081f
C268 B.n231 VSUBS 0.009081f
C269 B.n232 VSUBS 0.009081f
C270 B.n233 VSUBS 0.009081f
C271 B.n234 VSUBS 0.009081f
C272 B.n235 VSUBS 0.009081f
C273 B.n236 VSUBS 0.009081f
C274 B.n237 VSUBS 0.009081f
C275 B.n238 VSUBS 0.009081f
C276 B.n239 VSUBS 0.009081f
C277 B.n240 VSUBS 0.009081f
C278 B.n241 VSUBS 0.009081f
C279 B.n242 VSUBS 0.009081f
C280 B.n243 VSUBS 0.009081f
C281 B.n244 VSUBS 0.009081f
C282 B.n245 VSUBS 0.009081f
C283 B.n246 VSUBS 0.009081f
C284 B.n247 VSUBS 0.009081f
C285 B.n248 VSUBS 0.009081f
C286 B.n249 VSUBS 0.009081f
C287 B.n250 VSUBS 0.009081f
C288 B.n251 VSUBS 0.009081f
C289 B.n252 VSUBS 0.009081f
C290 B.n253 VSUBS 0.009081f
C291 B.n254 VSUBS 0.009081f
C292 B.n255 VSUBS 0.009081f
C293 B.n256 VSUBS 0.009081f
C294 B.n257 VSUBS 0.009081f
C295 B.n258 VSUBS 0.009081f
C296 B.n259 VSUBS 0.009081f
C297 B.n260 VSUBS 0.009081f
C298 B.n261 VSUBS 0.009081f
C299 B.n262 VSUBS 0.009081f
C300 B.n263 VSUBS 0.009081f
C301 B.n264 VSUBS 0.009081f
C302 B.n265 VSUBS 0.009081f
C303 B.n266 VSUBS 0.009081f
C304 B.n267 VSUBS 0.009081f
C305 B.n268 VSUBS 0.009081f
C306 B.n269 VSUBS 0.009081f
C307 B.n270 VSUBS 0.009081f
C308 B.n271 VSUBS 0.009081f
C309 B.n272 VSUBS 0.009081f
C310 B.n273 VSUBS 0.009081f
C311 B.n274 VSUBS 0.020613f
C312 B.n275 VSUBS 0.020613f
C313 B.n276 VSUBS 0.022387f
C314 B.n277 VSUBS 0.009081f
C315 B.n278 VSUBS 0.009081f
C316 B.n279 VSUBS 0.009081f
C317 B.n280 VSUBS 0.009081f
C318 B.n281 VSUBS 0.009081f
C319 B.n282 VSUBS 0.009081f
C320 B.n283 VSUBS 0.009081f
C321 B.n284 VSUBS 0.009081f
C322 B.n285 VSUBS 0.009081f
C323 B.n286 VSUBS 0.009081f
C324 B.n287 VSUBS 0.009081f
C325 B.n288 VSUBS 0.009081f
C326 B.n289 VSUBS 0.009081f
C327 B.n290 VSUBS 0.009081f
C328 B.n291 VSUBS 0.009081f
C329 B.n292 VSUBS 0.009081f
C330 B.n293 VSUBS 0.009081f
C331 B.n294 VSUBS 0.009081f
C332 B.n295 VSUBS 0.009081f
C333 B.n296 VSUBS 0.009081f
C334 B.n297 VSUBS 0.009081f
C335 B.n298 VSUBS 0.009081f
C336 B.n299 VSUBS 0.009081f
C337 B.n300 VSUBS 0.009081f
C338 B.n301 VSUBS 0.009081f
C339 B.n302 VSUBS 0.009081f
C340 B.n303 VSUBS 0.009081f
C341 B.n304 VSUBS 0.009081f
C342 B.n305 VSUBS 0.009081f
C343 B.n306 VSUBS 0.009081f
C344 B.n307 VSUBS 0.009081f
C345 B.n308 VSUBS 0.009081f
C346 B.n309 VSUBS 0.009081f
C347 B.n310 VSUBS 0.009081f
C348 B.n311 VSUBS 0.009081f
C349 B.n312 VSUBS 0.009081f
C350 B.n313 VSUBS 0.009081f
C351 B.n314 VSUBS 0.009081f
C352 B.n315 VSUBS 0.009081f
C353 B.n316 VSUBS 0.009081f
C354 B.n317 VSUBS 0.009081f
C355 B.n318 VSUBS 0.009081f
C356 B.n319 VSUBS 0.009081f
C357 B.n320 VSUBS 0.009081f
C358 B.n321 VSUBS 0.009081f
C359 B.n322 VSUBS 0.009081f
C360 B.n323 VSUBS 0.009081f
C361 B.n324 VSUBS 0.009081f
C362 B.n325 VSUBS 0.009081f
C363 B.n326 VSUBS 0.009081f
C364 B.n327 VSUBS 0.009081f
C365 B.t2 VSUBS 0.22024f
C366 B.t1 VSUBS 0.271382f
C367 B.t0 VSUBS 2.18026f
C368 B.n328 VSUBS 0.436313f
C369 B.n329 VSUBS 0.296199f
C370 B.n330 VSUBS 0.021039f
C371 B.n331 VSUBS 0.008547f
C372 B.n332 VSUBS 0.009081f
C373 B.n333 VSUBS 0.009081f
C374 B.n334 VSUBS 0.009081f
C375 B.n335 VSUBS 0.009081f
C376 B.n336 VSUBS 0.009081f
C377 B.n337 VSUBS 0.009081f
C378 B.n338 VSUBS 0.009081f
C379 B.n339 VSUBS 0.009081f
C380 B.n340 VSUBS 0.009081f
C381 B.n341 VSUBS 0.009081f
C382 B.n342 VSUBS 0.009081f
C383 B.n343 VSUBS 0.009081f
C384 B.n344 VSUBS 0.009081f
C385 B.n345 VSUBS 0.009081f
C386 B.n346 VSUBS 0.009081f
C387 B.n347 VSUBS 0.005075f
C388 B.n348 VSUBS 0.021039f
C389 B.n349 VSUBS 0.008547f
C390 B.n350 VSUBS 0.009081f
C391 B.n351 VSUBS 0.009081f
C392 B.n352 VSUBS 0.009081f
C393 B.n353 VSUBS 0.009081f
C394 B.n354 VSUBS 0.009081f
C395 B.n355 VSUBS 0.009081f
C396 B.n356 VSUBS 0.009081f
C397 B.n357 VSUBS 0.009081f
C398 B.n358 VSUBS 0.009081f
C399 B.n359 VSUBS 0.009081f
C400 B.n360 VSUBS 0.009081f
C401 B.n361 VSUBS 0.009081f
C402 B.n362 VSUBS 0.009081f
C403 B.n363 VSUBS 0.009081f
C404 B.n364 VSUBS 0.009081f
C405 B.n365 VSUBS 0.009081f
C406 B.n366 VSUBS 0.009081f
C407 B.n367 VSUBS 0.009081f
C408 B.n368 VSUBS 0.009081f
C409 B.n369 VSUBS 0.009081f
C410 B.n370 VSUBS 0.009081f
C411 B.n371 VSUBS 0.009081f
C412 B.n372 VSUBS 0.009081f
C413 B.n373 VSUBS 0.009081f
C414 B.n374 VSUBS 0.009081f
C415 B.n375 VSUBS 0.009081f
C416 B.n376 VSUBS 0.009081f
C417 B.n377 VSUBS 0.009081f
C418 B.n378 VSUBS 0.009081f
C419 B.n379 VSUBS 0.009081f
C420 B.n380 VSUBS 0.009081f
C421 B.n381 VSUBS 0.009081f
C422 B.n382 VSUBS 0.009081f
C423 B.n383 VSUBS 0.009081f
C424 B.n384 VSUBS 0.009081f
C425 B.n385 VSUBS 0.009081f
C426 B.n386 VSUBS 0.009081f
C427 B.n387 VSUBS 0.009081f
C428 B.n388 VSUBS 0.009081f
C429 B.n389 VSUBS 0.009081f
C430 B.n390 VSUBS 0.009081f
C431 B.n391 VSUBS 0.009081f
C432 B.n392 VSUBS 0.009081f
C433 B.n393 VSUBS 0.009081f
C434 B.n394 VSUBS 0.009081f
C435 B.n395 VSUBS 0.009081f
C436 B.n396 VSUBS 0.009081f
C437 B.n397 VSUBS 0.009081f
C438 B.n398 VSUBS 0.009081f
C439 B.n399 VSUBS 0.009081f
C440 B.n400 VSUBS 0.009081f
C441 B.n401 VSUBS 0.022387f
C442 B.n402 VSUBS 0.021333f
C443 B.n403 VSUBS 0.021667f
C444 B.n404 VSUBS 0.009081f
C445 B.n405 VSUBS 0.009081f
C446 B.n406 VSUBS 0.009081f
C447 B.n407 VSUBS 0.009081f
C448 B.n408 VSUBS 0.009081f
C449 B.n409 VSUBS 0.009081f
C450 B.n410 VSUBS 0.009081f
C451 B.n411 VSUBS 0.009081f
C452 B.n412 VSUBS 0.009081f
C453 B.n413 VSUBS 0.009081f
C454 B.n414 VSUBS 0.009081f
C455 B.n415 VSUBS 0.009081f
C456 B.n416 VSUBS 0.009081f
C457 B.n417 VSUBS 0.009081f
C458 B.n418 VSUBS 0.009081f
C459 B.n419 VSUBS 0.009081f
C460 B.n420 VSUBS 0.009081f
C461 B.n421 VSUBS 0.009081f
C462 B.n422 VSUBS 0.009081f
C463 B.n423 VSUBS 0.009081f
C464 B.n424 VSUBS 0.009081f
C465 B.n425 VSUBS 0.009081f
C466 B.n426 VSUBS 0.009081f
C467 B.n427 VSUBS 0.009081f
C468 B.n428 VSUBS 0.009081f
C469 B.n429 VSUBS 0.009081f
C470 B.n430 VSUBS 0.009081f
C471 B.n431 VSUBS 0.009081f
C472 B.n432 VSUBS 0.009081f
C473 B.n433 VSUBS 0.009081f
C474 B.n434 VSUBS 0.009081f
C475 B.n435 VSUBS 0.009081f
C476 B.n436 VSUBS 0.009081f
C477 B.n437 VSUBS 0.009081f
C478 B.n438 VSUBS 0.009081f
C479 B.n439 VSUBS 0.009081f
C480 B.n440 VSUBS 0.009081f
C481 B.n441 VSUBS 0.009081f
C482 B.n442 VSUBS 0.009081f
C483 B.n443 VSUBS 0.009081f
C484 B.n444 VSUBS 0.009081f
C485 B.n445 VSUBS 0.009081f
C486 B.n446 VSUBS 0.009081f
C487 B.n447 VSUBS 0.009081f
C488 B.n448 VSUBS 0.009081f
C489 B.n449 VSUBS 0.009081f
C490 B.n450 VSUBS 0.009081f
C491 B.n451 VSUBS 0.009081f
C492 B.n452 VSUBS 0.009081f
C493 B.n453 VSUBS 0.009081f
C494 B.n454 VSUBS 0.009081f
C495 B.n455 VSUBS 0.009081f
C496 B.n456 VSUBS 0.009081f
C497 B.n457 VSUBS 0.009081f
C498 B.n458 VSUBS 0.009081f
C499 B.n459 VSUBS 0.009081f
C500 B.n460 VSUBS 0.009081f
C501 B.n461 VSUBS 0.009081f
C502 B.n462 VSUBS 0.009081f
C503 B.n463 VSUBS 0.009081f
C504 B.n464 VSUBS 0.009081f
C505 B.n465 VSUBS 0.009081f
C506 B.n466 VSUBS 0.009081f
C507 B.n467 VSUBS 0.009081f
C508 B.n468 VSUBS 0.009081f
C509 B.n469 VSUBS 0.009081f
C510 B.n470 VSUBS 0.009081f
C511 B.n471 VSUBS 0.009081f
C512 B.n472 VSUBS 0.009081f
C513 B.n473 VSUBS 0.009081f
C514 B.n474 VSUBS 0.009081f
C515 B.n475 VSUBS 0.009081f
C516 B.n476 VSUBS 0.009081f
C517 B.n477 VSUBS 0.009081f
C518 B.n478 VSUBS 0.009081f
C519 B.n479 VSUBS 0.009081f
C520 B.n480 VSUBS 0.009081f
C521 B.n481 VSUBS 0.009081f
C522 B.n482 VSUBS 0.009081f
C523 B.n483 VSUBS 0.009081f
C524 B.n484 VSUBS 0.009081f
C525 B.n485 VSUBS 0.009081f
C526 B.n486 VSUBS 0.009081f
C527 B.n487 VSUBS 0.009081f
C528 B.n488 VSUBS 0.009081f
C529 B.n489 VSUBS 0.009081f
C530 B.n490 VSUBS 0.009081f
C531 B.n491 VSUBS 0.009081f
C532 B.n492 VSUBS 0.009081f
C533 B.n493 VSUBS 0.009081f
C534 B.n494 VSUBS 0.009081f
C535 B.n495 VSUBS 0.009081f
C536 B.n496 VSUBS 0.009081f
C537 B.n497 VSUBS 0.009081f
C538 B.n498 VSUBS 0.009081f
C539 B.n499 VSUBS 0.009081f
C540 B.n500 VSUBS 0.009081f
C541 B.n501 VSUBS 0.009081f
C542 B.n502 VSUBS 0.009081f
C543 B.n503 VSUBS 0.009081f
C544 B.n504 VSUBS 0.009081f
C545 B.n505 VSUBS 0.009081f
C546 B.n506 VSUBS 0.009081f
C547 B.n507 VSUBS 0.009081f
C548 B.n508 VSUBS 0.009081f
C549 B.n509 VSUBS 0.009081f
C550 B.n510 VSUBS 0.009081f
C551 B.n511 VSUBS 0.009081f
C552 B.n512 VSUBS 0.009081f
C553 B.n513 VSUBS 0.009081f
C554 B.n514 VSUBS 0.009081f
C555 B.n515 VSUBS 0.009081f
C556 B.n516 VSUBS 0.009081f
C557 B.n517 VSUBS 0.009081f
C558 B.n518 VSUBS 0.009081f
C559 B.n519 VSUBS 0.009081f
C560 B.n520 VSUBS 0.009081f
C561 B.n521 VSUBS 0.009081f
C562 B.n522 VSUBS 0.009081f
C563 B.n523 VSUBS 0.009081f
C564 B.n524 VSUBS 0.009081f
C565 B.n525 VSUBS 0.009081f
C566 B.n526 VSUBS 0.009081f
C567 B.n527 VSUBS 0.009081f
C568 B.n528 VSUBS 0.009081f
C569 B.n529 VSUBS 0.009081f
C570 B.n530 VSUBS 0.009081f
C571 B.n531 VSUBS 0.009081f
C572 B.n532 VSUBS 0.009081f
C573 B.n533 VSUBS 0.009081f
C574 B.n534 VSUBS 0.009081f
C575 B.n535 VSUBS 0.009081f
C576 B.n536 VSUBS 0.009081f
C577 B.n537 VSUBS 0.009081f
C578 B.n538 VSUBS 0.009081f
C579 B.n539 VSUBS 0.009081f
C580 B.n540 VSUBS 0.009081f
C581 B.n541 VSUBS 0.009081f
C582 B.n542 VSUBS 0.009081f
C583 B.n543 VSUBS 0.009081f
C584 B.n544 VSUBS 0.009081f
C585 B.n545 VSUBS 0.009081f
C586 B.n546 VSUBS 0.009081f
C587 B.n547 VSUBS 0.009081f
C588 B.n548 VSUBS 0.009081f
C589 B.n549 VSUBS 0.009081f
C590 B.n550 VSUBS 0.009081f
C591 B.n551 VSUBS 0.009081f
C592 B.n552 VSUBS 0.009081f
C593 B.n553 VSUBS 0.009081f
C594 B.n554 VSUBS 0.009081f
C595 B.n555 VSUBS 0.009081f
C596 B.n556 VSUBS 0.009081f
C597 B.n557 VSUBS 0.009081f
C598 B.n558 VSUBS 0.009081f
C599 B.n559 VSUBS 0.009081f
C600 B.n560 VSUBS 0.009081f
C601 B.n561 VSUBS 0.009081f
C602 B.n562 VSUBS 0.009081f
C603 B.n563 VSUBS 0.020613f
C604 B.n564 VSUBS 0.020613f
C605 B.n565 VSUBS 0.022387f
C606 B.n566 VSUBS 0.009081f
C607 B.n567 VSUBS 0.009081f
C608 B.n568 VSUBS 0.009081f
C609 B.n569 VSUBS 0.009081f
C610 B.n570 VSUBS 0.009081f
C611 B.n571 VSUBS 0.009081f
C612 B.n572 VSUBS 0.009081f
C613 B.n573 VSUBS 0.009081f
C614 B.n574 VSUBS 0.009081f
C615 B.n575 VSUBS 0.009081f
C616 B.n576 VSUBS 0.009081f
C617 B.n577 VSUBS 0.009081f
C618 B.n578 VSUBS 0.009081f
C619 B.n579 VSUBS 0.009081f
C620 B.n580 VSUBS 0.009081f
C621 B.n581 VSUBS 0.009081f
C622 B.n582 VSUBS 0.009081f
C623 B.n583 VSUBS 0.009081f
C624 B.n584 VSUBS 0.009081f
C625 B.n585 VSUBS 0.009081f
C626 B.n586 VSUBS 0.009081f
C627 B.n587 VSUBS 0.009081f
C628 B.n588 VSUBS 0.009081f
C629 B.n589 VSUBS 0.009081f
C630 B.n590 VSUBS 0.009081f
C631 B.n591 VSUBS 0.009081f
C632 B.n592 VSUBS 0.009081f
C633 B.n593 VSUBS 0.009081f
C634 B.n594 VSUBS 0.009081f
C635 B.n595 VSUBS 0.009081f
C636 B.n596 VSUBS 0.009081f
C637 B.n597 VSUBS 0.009081f
C638 B.n598 VSUBS 0.009081f
C639 B.n599 VSUBS 0.009081f
C640 B.n600 VSUBS 0.009081f
C641 B.n601 VSUBS 0.009081f
C642 B.n602 VSUBS 0.009081f
C643 B.n603 VSUBS 0.009081f
C644 B.n604 VSUBS 0.009081f
C645 B.n605 VSUBS 0.009081f
C646 B.n606 VSUBS 0.009081f
C647 B.n607 VSUBS 0.009081f
C648 B.n608 VSUBS 0.009081f
C649 B.n609 VSUBS 0.009081f
C650 B.n610 VSUBS 0.009081f
C651 B.n611 VSUBS 0.009081f
C652 B.n612 VSUBS 0.009081f
C653 B.n613 VSUBS 0.009081f
C654 B.n614 VSUBS 0.009081f
C655 B.n615 VSUBS 0.009081f
C656 B.n616 VSUBS 0.009081f
C657 B.n617 VSUBS 0.009081f
C658 B.n618 VSUBS 0.008547f
C659 B.n619 VSUBS 0.021039f
C660 B.n620 VSUBS 0.005075f
C661 B.n621 VSUBS 0.009081f
C662 B.n622 VSUBS 0.009081f
C663 B.n623 VSUBS 0.009081f
C664 B.n624 VSUBS 0.009081f
C665 B.n625 VSUBS 0.009081f
C666 B.n626 VSUBS 0.009081f
C667 B.n627 VSUBS 0.009081f
C668 B.n628 VSUBS 0.009081f
C669 B.n629 VSUBS 0.009081f
C670 B.n630 VSUBS 0.009081f
C671 B.n631 VSUBS 0.009081f
C672 B.n632 VSUBS 0.009081f
C673 B.n633 VSUBS 0.005075f
C674 B.n634 VSUBS 0.009081f
C675 B.n635 VSUBS 0.009081f
C676 B.n636 VSUBS 0.009081f
C677 B.n637 VSUBS 0.009081f
C678 B.n638 VSUBS 0.009081f
C679 B.n639 VSUBS 0.009081f
C680 B.n640 VSUBS 0.009081f
C681 B.n641 VSUBS 0.009081f
C682 B.n642 VSUBS 0.009081f
C683 B.n643 VSUBS 0.009081f
C684 B.n644 VSUBS 0.009081f
C685 B.n645 VSUBS 0.009081f
C686 B.n646 VSUBS 0.009081f
C687 B.n647 VSUBS 0.009081f
C688 B.n648 VSUBS 0.009081f
C689 B.n649 VSUBS 0.009081f
C690 B.n650 VSUBS 0.009081f
C691 B.n651 VSUBS 0.009081f
C692 B.n652 VSUBS 0.009081f
C693 B.n653 VSUBS 0.009081f
C694 B.n654 VSUBS 0.009081f
C695 B.n655 VSUBS 0.009081f
C696 B.n656 VSUBS 0.009081f
C697 B.n657 VSUBS 0.009081f
C698 B.n658 VSUBS 0.009081f
C699 B.n659 VSUBS 0.009081f
C700 B.n660 VSUBS 0.009081f
C701 B.n661 VSUBS 0.009081f
C702 B.n662 VSUBS 0.009081f
C703 B.n663 VSUBS 0.009081f
C704 B.n664 VSUBS 0.009081f
C705 B.n665 VSUBS 0.009081f
C706 B.n666 VSUBS 0.009081f
C707 B.n667 VSUBS 0.009081f
C708 B.n668 VSUBS 0.009081f
C709 B.n669 VSUBS 0.009081f
C710 B.n670 VSUBS 0.009081f
C711 B.n671 VSUBS 0.009081f
C712 B.n672 VSUBS 0.009081f
C713 B.n673 VSUBS 0.009081f
C714 B.n674 VSUBS 0.009081f
C715 B.n675 VSUBS 0.009081f
C716 B.n676 VSUBS 0.009081f
C717 B.n677 VSUBS 0.009081f
C718 B.n678 VSUBS 0.009081f
C719 B.n679 VSUBS 0.009081f
C720 B.n680 VSUBS 0.009081f
C721 B.n681 VSUBS 0.009081f
C722 B.n682 VSUBS 0.009081f
C723 B.n683 VSUBS 0.009081f
C724 B.n684 VSUBS 0.009081f
C725 B.n685 VSUBS 0.009081f
C726 B.n686 VSUBS 0.009081f
C727 B.n687 VSUBS 0.022387f
C728 B.n688 VSUBS 0.022387f
C729 B.n689 VSUBS 0.020613f
C730 B.n690 VSUBS 0.009081f
C731 B.n691 VSUBS 0.009081f
C732 B.n692 VSUBS 0.009081f
C733 B.n693 VSUBS 0.009081f
C734 B.n694 VSUBS 0.009081f
C735 B.n695 VSUBS 0.009081f
C736 B.n696 VSUBS 0.009081f
C737 B.n697 VSUBS 0.009081f
C738 B.n698 VSUBS 0.009081f
C739 B.n699 VSUBS 0.009081f
C740 B.n700 VSUBS 0.009081f
C741 B.n701 VSUBS 0.009081f
C742 B.n702 VSUBS 0.009081f
C743 B.n703 VSUBS 0.009081f
C744 B.n704 VSUBS 0.009081f
C745 B.n705 VSUBS 0.009081f
C746 B.n706 VSUBS 0.009081f
C747 B.n707 VSUBS 0.009081f
C748 B.n708 VSUBS 0.009081f
C749 B.n709 VSUBS 0.009081f
C750 B.n710 VSUBS 0.009081f
C751 B.n711 VSUBS 0.009081f
C752 B.n712 VSUBS 0.009081f
C753 B.n713 VSUBS 0.009081f
C754 B.n714 VSUBS 0.009081f
C755 B.n715 VSUBS 0.009081f
C756 B.n716 VSUBS 0.009081f
C757 B.n717 VSUBS 0.009081f
C758 B.n718 VSUBS 0.009081f
C759 B.n719 VSUBS 0.009081f
C760 B.n720 VSUBS 0.009081f
C761 B.n721 VSUBS 0.009081f
C762 B.n722 VSUBS 0.009081f
C763 B.n723 VSUBS 0.009081f
C764 B.n724 VSUBS 0.009081f
C765 B.n725 VSUBS 0.009081f
C766 B.n726 VSUBS 0.009081f
C767 B.n727 VSUBS 0.009081f
C768 B.n728 VSUBS 0.009081f
C769 B.n729 VSUBS 0.009081f
C770 B.n730 VSUBS 0.009081f
C771 B.n731 VSUBS 0.009081f
C772 B.n732 VSUBS 0.009081f
C773 B.n733 VSUBS 0.009081f
C774 B.n734 VSUBS 0.009081f
C775 B.n735 VSUBS 0.009081f
C776 B.n736 VSUBS 0.009081f
C777 B.n737 VSUBS 0.009081f
C778 B.n738 VSUBS 0.009081f
C779 B.n739 VSUBS 0.009081f
C780 B.n740 VSUBS 0.009081f
C781 B.n741 VSUBS 0.009081f
C782 B.n742 VSUBS 0.009081f
C783 B.n743 VSUBS 0.009081f
C784 B.n744 VSUBS 0.009081f
C785 B.n745 VSUBS 0.009081f
C786 B.n746 VSUBS 0.009081f
C787 B.n747 VSUBS 0.009081f
C788 B.n748 VSUBS 0.009081f
C789 B.n749 VSUBS 0.009081f
C790 B.n750 VSUBS 0.009081f
C791 B.n751 VSUBS 0.009081f
C792 B.n752 VSUBS 0.009081f
C793 B.n753 VSUBS 0.009081f
C794 B.n754 VSUBS 0.009081f
C795 B.n755 VSUBS 0.009081f
C796 B.n756 VSUBS 0.009081f
C797 B.n757 VSUBS 0.009081f
C798 B.n758 VSUBS 0.009081f
C799 B.n759 VSUBS 0.009081f
C800 B.n760 VSUBS 0.009081f
C801 B.n761 VSUBS 0.009081f
C802 B.n762 VSUBS 0.009081f
C803 B.n763 VSUBS 0.009081f
C804 B.n764 VSUBS 0.009081f
C805 B.n765 VSUBS 0.009081f
C806 B.n766 VSUBS 0.009081f
C807 B.n767 VSUBS 0.01185f
C808 B.n768 VSUBS 0.012623f
C809 B.n769 VSUBS 0.025103f
C810 VDD2.n0 VSUBS 0.032086f
C811 VDD2.n1 VSUBS 0.029088f
C812 VDD2.n2 VSUBS 0.015631f
C813 VDD2.n3 VSUBS 0.036945f
C814 VDD2.n4 VSUBS 0.01655f
C815 VDD2.n5 VSUBS 0.029088f
C816 VDD2.n6 VSUBS 0.01609f
C817 VDD2.n7 VSUBS 0.036945f
C818 VDD2.n8 VSUBS 0.01655f
C819 VDD2.n9 VSUBS 0.029088f
C820 VDD2.n10 VSUBS 0.015631f
C821 VDD2.n11 VSUBS 0.036945f
C822 VDD2.n12 VSUBS 0.01655f
C823 VDD2.n13 VSUBS 0.029088f
C824 VDD2.n14 VSUBS 0.015631f
C825 VDD2.n15 VSUBS 0.027709f
C826 VDD2.n16 VSUBS 0.027792f
C827 VDD2.t3 VSUBS 0.079454f
C828 VDD2.n17 VSUBS 0.20412f
C829 VDD2.n18 VSUBS 1.18697f
C830 VDD2.n19 VSUBS 0.015631f
C831 VDD2.n20 VSUBS 0.01655f
C832 VDD2.n21 VSUBS 0.036945f
C833 VDD2.n22 VSUBS 0.036945f
C834 VDD2.n23 VSUBS 0.01655f
C835 VDD2.n24 VSUBS 0.015631f
C836 VDD2.n25 VSUBS 0.029088f
C837 VDD2.n26 VSUBS 0.029088f
C838 VDD2.n27 VSUBS 0.015631f
C839 VDD2.n28 VSUBS 0.01655f
C840 VDD2.n29 VSUBS 0.036945f
C841 VDD2.n30 VSUBS 0.036945f
C842 VDD2.n31 VSUBS 0.01655f
C843 VDD2.n32 VSUBS 0.015631f
C844 VDD2.n33 VSUBS 0.029088f
C845 VDD2.n34 VSUBS 0.029088f
C846 VDD2.n35 VSUBS 0.015631f
C847 VDD2.n36 VSUBS 0.015631f
C848 VDD2.n37 VSUBS 0.01655f
C849 VDD2.n38 VSUBS 0.036945f
C850 VDD2.n39 VSUBS 0.036945f
C851 VDD2.n40 VSUBS 0.036945f
C852 VDD2.n41 VSUBS 0.01609f
C853 VDD2.n42 VSUBS 0.015631f
C854 VDD2.n43 VSUBS 0.029088f
C855 VDD2.n44 VSUBS 0.029088f
C856 VDD2.n45 VSUBS 0.015631f
C857 VDD2.n46 VSUBS 0.01655f
C858 VDD2.n47 VSUBS 0.036945f
C859 VDD2.n48 VSUBS 0.089866f
C860 VDD2.n49 VSUBS 0.01655f
C861 VDD2.n50 VSUBS 0.015631f
C862 VDD2.n51 VSUBS 0.072799f
C863 VDD2.n52 VSUBS 0.078562f
C864 VDD2.t1 VSUBS 0.232161f
C865 VDD2.t2 VSUBS 0.232161f
C866 VDD2.n53 VSUBS 1.77397f
C867 VDD2.n54 VSUBS 3.73709f
C868 VDD2.n55 VSUBS 0.032086f
C869 VDD2.n56 VSUBS 0.029088f
C870 VDD2.n57 VSUBS 0.015631f
C871 VDD2.n58 VSUBS 0.036945f
C872 VDD2.n59 VSUBS 0.01655f
C873 VDD2.n60 VSUBS 0.029088f
C874 VDD2.n61 VSUBS 0.01609f
C875 VDD2.n62 VSUBS 0.036945f
C876 VDD2.n63 VSUBS 0.015631f
C877 VDD2.n64 VSUBS 0.01655f
C878 VDD2.n65 VSUBS 0.029088f
C879 VDD2.n66 VSUBS 0.015631f
C880 VDD2.n67 VSUBS 0.036945f
C881 VDD2.n68 VSUBS 0.01655f
C882 VDD2.n69 VSUBS 0.029088f
C883 VDD2.n70 VSUBS 0.015631f
C884 VDD2.n71 VSUBS 0.027709f
C885 VDD2.n72 VSUBS 0.027792f
C886 VDD2.t5 VSUBS 0.079454f
C887 VDD2.n73 VSUBS 0.20412f
C888 VDD2.n74 VSUBS 1.18697f
C889 VDD2.n75 VSUBS 0.015631f
C890 VDD2.n76 VSUBS 0.01655f
C891 VDD2.n77 VSUBS 0.036945f
C892 VDD2.n78 VSUBS 0.036945f
C893 VDD2.n79 VSUBS 0.01655f
C894 VDD2.n80 VSUBS 0.015631f
C895 VDD2.n81 VSUBS 0.029088f
C896 VDD2.n82 VSUBS 0.029088f
C897 VDD2.n83 VSUBS 0.015631f
C898 VDD2.n84 VSUBS 0.01655f
C899 VDD2.n85 VSUBS 0.036945f
C900 VDD2.n86 VSUBS 0.036945f
C901 VDD2.n87 VSUBS 0.01655f
C902 VDD2.n88 VSUBS 0.015631f
C903 VDD2.n89 VSUBS 0.029088f
C904 VDD2.n90 VSUBS 0.029088f
C905 VDD2.n91 VSUBS 0.015631f
C906 VDD2.n92 VSUBS 0.01655f
C907 VDD2.n93 VSUBS 0.036945f
C908 VDD2.n94 VSUBS 0.036945f
C909 VDD2.n95 VSUBS 0.036945f
C910 VDD2.n96 VSUBS 0.01609f
C911 VDD2.n97 VSUBS 0.015631f
C912 VDD2.n98 VSUBS 0.029088f
C913 VDD2.n99 VSUBS 0.029088f
C914 VDD2.n100 VSUBS 0.015631f
C915 VDD2.n101 VSUBS 0.01655f
C916 VDD2.n102 VSUBS 0.036945f
C917 VDD2.n103 VSUBS 0.089866f
C918 VDD2.n104 VSUBS 0.01655f
C919 VDD2.n105 VSUBS 0.015631f
C920 VDD2.n106 VSUBS 0.072799f
C921 VDD2.n107 VSUBS 0.065421f
C922 VDD2.n108 VSUBS 3.11495f
C923 VDD2.t0 VSUBS 0.232161f
C924 VDD2.t4 VSUBS 0.232161f
C925 VDD2.n109 VSUBS 1.77393f
C926 VN.t3 VSUBS 2.65847f
C927 VN.n0 VSUBS 1.04203f
C928 VN.n1 VSUBS 0.02736f
C929 VN.n2 VSUBS 0.044314f
C930 VN.n3 VSUBS 0.02736f
C931 VN.n4 VSUBS 0.038213f
C932 VN.t4 VSUBS 2.65847f
C933 VN.n5 VSUBS 1.03521f
C934 VN.t2 VSUBS 3.02906f
C935 VN.n6 VSUBS 0.983776f
C936 VN.n7 VSUBS 0.341001f
C937 VN.n8 VSUBS 0.02736f
C938 VN.n9 VSUBS 0.050737f
C939 VN.n10 VSUBS 0.050737f
C940 VN.n11 VSUBS 0.03523f
C941 VN.n12 VSUBS 0.02736f
C942 VN.n13 VSUBS 0.02736f
C943 VN.n14 VSUBS 0.02736f
C944 VN.n15 VSUBS 0.050737f
C945 VN.n16 VSUBS 0.050737f
C946 VN.n17 VSUBS 0.032201f
C947 VN.n18 VSUBS 0.044151f
C948 VN.n19 VSUBS 0.077383f
C949 VN.t0 VSUBS 2.65847f
C950 VN.n20 VSUBS 1.04203f
C951 VN.n21 VSUBS 0.02736f
C952 VN.n22 VSUBS 0.044314f
C953 VN.n23 VSUBS 0.02736f
C954 VN.n24 VSUBS 0.038213f
C955 VN.t1 VSUBS 3.02906f
C956 VN.t5 VSUBS 2.65847f
C957 VN.n25 VSUBS 1.03521f
C958 VN.n26 VSUBS 0.983776f
C959 VN.n27 VSUBS 0.341001f
C960 VN.n28 VSUBS 0.02736f
C961 VN.n29 VSUBS 0.050737f
C962 VN.n30 VSUBS 0.050737f
C963 VN.n31 VSUBS 0.03523f
C964 VN.n32 VSUBS 0.02736f
C965 VN.n33 VSUBS 0.02736f
C966 VN.n34 VSUBS 0.02736f
C967 VN.n35 VSUBS 0.050737f
C968 VN.n36 VSUBS 0.050737f
C969 VN.n37 VSUBS 0.032201f
C970 VN.n38 VSUBS 0.044151f
C971 VN.n39 VSUBS 1.62299f
C972 VDD1.n0 VSUBS 0.032074f
C973 VDD1.n1 VSUBS 0.029076f
C974 VDD1.n2 VSUBS 0.015624f
C975 VDD1.n3 VSUBS 0.03693f
C976 VDD1.n4 VSUBS 0.016543f
C977 VDD1.n5 VSUBS 0.029076f
C978 VDD1.n6 VSUBS 0.016084f
C979 VDD1.n7 VSUBS 0.03693f
C980 VDD1.n8 VSUBS 0.015624f
C981 VDD1.n9 VSUBS 0.016543f
C982 VDD1.n10 VSUBS 0.029076f
C983 VDD1.n11 VSUBS 0.015624f
C984 VDD1.n12 VSUBS 0.03693f
C985 VDD1.n13 VSUBS 0.016543f
C986 VDD1.n14 VSUBS 0.029076f
C987 VDD1.n15 VSUBS 0.015624f
C988 VDD1.n16 VSUBS 0.027698f
C989 VDD1.n17 VSUBS 0.027781f
C990 VDD1.t0 VSUBS 0.079422f
C991 VDD1.n18 VSUBS 0.204038f
C992 VDD1.n19 VSUBS 1.18649f
C993 VDD1.n20 VSUBS 0.015624f
C994 VDD1.n21 VSUBS 0.016543f
C995 VDD1.n22 VSUBS 0.03693f
C996 VDD1.n23 VSUBS 0.03693f
C997 VDD1.n24 VSUBS 0.016543f
C998 VDD1.n25 VSUBS 0.015624f
C999 VDD1.n26 VSUBS 0.029076f
C1000 VDD1.n27 VSUBS 0.029076f
C1001 VDD1.n28 VSUBS 0.015624f
C1002 VDD1.n29 VSUBS 0.016543f
C1003 VDD1.n30 VSUBS 0.03693f
C1004 VDD1.n31 VSUBS 0.03693f
C1005 VDD1.n32 VSUBS 0.016543f
C1006 VDD1.n33 VSUBS 0.015624f
C1007 VDD1.n34 VSUBS 0.029076f
C1008 VDD1.n35 VSUBS 0.029076f
C1009 VDD1.n36 VSUBS 0.015624f
C1010 VDD1.n37 VSUBS 0.016543f
C1011 VDD1.n38 VSUBS 0.03693f
C1012 VDD1.n39 VSUBS 0.03693f
C1013 VDD1.n40 VSUBS 0.03693f
C1014 VDD1.n41 VSUBS 0.016084f
C1015 VDD1.n42 VSUBS 0.015624f
C1016 VDD1.n43 VSUBS 0.029076f
C1017 VDD1.n44 VSUBS 0.029076f
C1018 VDD1.n45 VSUBS 0.015624f
C1019 VDD1.n46 VSUBS 0.016543f
C1020 VDD1.n47 VSUBS 0.03693f
C1021 VDD1.n48 VSUBS 0.08983f
C1022 VDD1.n49 VSUBS 0.016543f
C1023 VDD1.n50 VSUBS 0.015624f
C1024 VDD1.n51 VSUBS 0.072769f
C1025 VDD1.n52 VSUBS 0.0796f
C1026 VDD1.n53 VSUBS 0.032074f
C1027 VDD1.n54 VSUBS 0.029076f
C1028 VDD1.n55 VSUBS 0.015624f
C1029 VDD1.n56 VSUBS 0.03693f
C1030 VDD1.n57 VSUBS 0.016543f
C1031 VDD1.n58 VSUBS 0.029076f
C1032 VDD1.n59 VSUBS 0.016084f
C1033 VDD1.n60 VSUBS 0.03693f
C1034 VDD1.n61 VSUBS 0.016543f
C1035 VDD1.n62 VSUBS 0.029076f
C1036 VDD1.n63 VSUBS 0.015624f
C1037 VDD1.n64 VSUBS 0.03693f
C1038 VDD1.n65 VSUBS 0.016543f
C1039 VDD1.n66 VSUBS 0.029076f
C1040 VDD1.n67 VSUBS 0.015624f
C1041 VDD1.n68 VSUBS 0.027698f
C1042 VDD1.n69 VSUBS 0.027781f
C1043 VDD1.t1 VSUBS 0.079422f
C1044 VDD1.n70 VSUBS 0.204038f
C1045 VDD1.n71 VSUBS 1.18649f
C1046 VDD1.n72 VSUBS 0.015624f
C1047 VDD1.n73 VSUBS 0.016543f
C1048 VDD1.n74 VSUBS 0.03693f
C1049 VDD1.n75 VSUBS 0.03693f
C1050 VDD1.n76 VSUBS 0.016543f
C1051 VDD1.n77 VSUBS 0.015624f
C1052 VDD1.n78 VSUBS 0.029076f
C1053 VDD1.n79 VSUBS 0.029076f
C1054 VDD1.n80 VSUBS 0.015624f
C1055 VDD1.n81 VSUBS 0.016543f
C1056 VDD1.n82 VSUBS 0.03693f
C1057 VDD1.n83 VSUBS 0.03693f
C1058 VDD1.n84 VSUBS 0.016543f
C1059 VDD1.n85 VSUBS 0.015624f
C1060 VDD1.n86 VSUBS 0.029076f
C1061 VDD1.n87 VSUBS 0.029076f
C1062 VDD1.n88 VSUBS 0.015624f
C1063 VDD1.n89 VSUBS 0.015624f
C1064 VDD1.n90 VSUBS 0.016543f
C1065 VDD1.n91 VSUBS 0.03693f
C1066 VDD1.n92 VSUBS 0.03693f
C1067 VDD1.n93 VSUBS 0.03693f
C1068 VDD1.n94 VSUBS 0.016084f
C1069 VDD1.n95 VSUBS 0.015624f
C1070 VDD1.n96 VSUBS 0.029076f
C1071 VDD1.n97 VSUBS 0.029076f
C1072 VDD1.n98 VSUBS 0.015624f
C1073 VDD1.n99 VSUBS 0.016543f
C1074 VDD1.n100 VSUBS 0.03693f
C1075 VDD1.n101 VSUBS 0.08983f
C1076 VDD1.n102 VSUBS 0.016543f
C1077 VDD1.n103 VSUBS 0.015624f
C1078 VDD1.n104 VSUBS 0.072769f
C1079 VDD1.n105 VSUBS 0.07853f
C1080 VDD1.t4 VSUBS 0.232067f
C1081 VDD1.t5 VSUBS 0.232067f
C1082 VDD1.n106 VSUBS 1.77326f
C1083 VDD1.n107 VSUBS 3.90719f
C1084 VDD1.t3 VSUBS 0.232067f
C1085 VDD1.t2 VSUBS 0.232067f
C1086 VDD1.n108 VSUBS 1.76438f
C1087 VDD1.n109 VSUBS 3.66556f
C1088 VTAIL.t4 VSUBS 0.245964f
C1089 VTAIL.t0 VSUBS 0.245964f
C1090 VTAIL.n0 VSUBS 1.72665f
C1091 VTAIL.n1 VSUBS 0.951798f
C1092 VTAIL.n2 VSUBS 0.033994f
C1093 VTAIL.n3 VSUBS 0.030817f
C1094 VTAIL.n4 VSUBS 0.01656f
C1095 VTAIL.n5 VSUBS 0.039142f
C1096 VTAIL.n6 VSUBS 0.017534f
C1097 VTAIL.n7 VSUBS 0.030817f
C1098 VTAIL.n8 VSUBS 0.017047f
C1099 VTAIL.n9 VSUBS 0.039142f
C1100 VTAIL.n10 VSUBS 0.017534f
C1101 VTAIL.n11 VSUBS 0.030817f
C1102 VTAIL.n12 VSUBS 0.01656f
C1103 VTAIL.n13 VSUBS 0.039142f
C1104 VTAIL.n14 VSUBS 0.017534f
C1105 VTAIL.n15 VSUBS 0.030817f
C1106 VTAIL.n16 VSUBS 0.01656f
C1107 VTAIL.n17 VSUBS 0.029356f
C1108 VTAIL.n18 VSUBS 0.029444f
C1109 VTAIL.t8 VSUBS 0.084178f
C1110 VTAIL.n19 VSUBS 0.216256f
C1111 VTAIL.n20 VSUBS 1.25754f
C1112 VTAIL.n21 VSUBS 0.01656f
C1113 VTAIL.n22 VSUBS 0.017534f
C1114 VTAIL.n23 VSUBS 0.039142f
C1115 VTAIL.n24 VSUBS 0.039142f
C1116 VTAIL.n25 VSUBS 0.017534f
C1117 VTAIL.n26 VSUBS 0.01656f
C1118 VTAIL.n27 VSUBS 0.030817f
C1119 VTAIL.n28 VSUBS 0.030817f
C1120 VTAIL.n29 VSUBS 0.01656f
C1121 VTAIL.n30 VSUBS 0.017534f
C1122 VTAIL.n31 VSUBS 0.039142f
C1123 VTAIL.n32 VSUBS 0.039142f
C1124 VTAIL.n33 VSUBS 0.017534f
C1125 VTAIL.n34 VSUBS 0.01656f
C1126 VTAIL.n35 VSUBS 0.030817f
C1127 VTAIL.n36 VSUBS 0.030817f
C1128 VTAIL.n37 VSUBS 0.01656f
C1129 VTAIL.n38 VSUBS 0.01656f
C1130 VTAIL.n39 VSUBS 0.017534f
C1131 VTAIL.n40 VSUBS 0.039142f
C1132 VTAIL.n41 VSUBS 0.039142f
C1133 VTAIL.n42 VSUBS 0.039142f
C1134 VTAIL.n43 VSUBS 0.017047f
C1135 VTAIL.n44 VSUBS 0.01656f
C1136 VTAIL.n45 VSUBS 0.030817f
C1137 VTAIL.n46 VSUBS 0.030817f
C1138 VTAIL.n47 VSUBS 0.01656f
C1139 VTAIL.n48 VSUBS 0.017534f
C1140 VTAIL.n49 VSUBS 0.039142f
C1141 VTAIL.n50 VSUBS 0.095209f
C1142 VTAIL.n51 VSUBS 0.017534f
C1143 VTAIL.n52 VSUBS 0.01656f
C1144 VTAIL.n53 VSUBS 0.077127f
C1145 VTAIL.n54 VSUBS 0.048074f
C1146 VTAIL.n55 VSUBS 0.574522f
C1147 VTAIL.t6 VSUBS 0.245964f
C1148 VTAIL.t11 VSUBS 0.245964f
C1149 VTAIL.n56 VSUBS 1.72665f
C1150 VTAIL.n57 VSUBS 2.9299f
C1151 VTAIL.t2 VSUBS 0.245964f
C1152 VTAIL.t5 VSUBS 0.245964f
C1153 VTAIL.n58 VSUBS 1.72666f
C1154 VTAIL.n59 VSUBS 2.92989f
C1155 VTAIL.n60 VSUBS 0.033994f
C1156 VTAIL.n61 VSUBS 0.030817f
C1157 VTAIL.n62 VSUBS 0.01656f
C1158 VTAIL.n63 VSUBS 0.039142f
C1159 VTAIL.n64 VSUBS 0.017534f
C1160 VTAIL.n65 VSUBS 0.030817f
C1161 VTAIL.n66 VSUBS 0.017047f
C1162 VTAIL.n67 VSUBS 0.039142f
C1163 VTAIL.n68 VSUBS 0.01656f
C1164 VTAIL.n69 VSUBS 0.017534f
C1165 VTAIL.n70 VSUBS 0.030817f
C1166 VTAIL.n71 VSUBS 0.01656f
C1167 VTAIL.n72 VSUBS 0.039142f
C1168 VTAIL.n73 VSUBS 0.017534f
C1169 VTAIL.n74 VSUBS 0.030817f
C1170 VTAIL.n75 VSUBS 0.01656f
C1171 VTAIL.n76 VSUBS 0.029356f
C1172 VTAIL.n77 VSUBS 0.029444f
C1173 VTAIL.t3 VSUBS 0.084178f
C1174 VTAIL.n78 VSUBS 0.216256f
C1175 VTAIL.n79 VSUBS 1.25754f
C1176 VTAIL.n80 VSUBS 0.01656f
C1177 VTAIL.n81 VSUBS 0.017534f
C1178 VTAIL.n82 VSUBS 0.039142f
C1179 VTAIL.n83 VSUBS 0.039142f
C1180 VTAIL.n84 VSUBS 0.017534f
C1181 VTAIL.n85 VSUBS 0.01656f
C1182 VTAIL.n86 VSUBS 0.030817f
C1183 VTAIL.n87 VSUBS 0.030817f
C1184 VTAIL.n88 VSUBS 0.01656f
C1185 VTAIL.n89 VSUBS 0.017534f
C1186 VTAIL.n90 VSUBS 0.039142f
C1187 VTAIL.n91 VSUBS 0.039142f
C1188 VTAIL.n92 VSUBS 0.017534f
C1189 VTAIL.n93 VSUBS 0.01656f
C1190 VTAIL.n94 VSUBS 0.030817f
C1191 VTAIL.n95 VSUBS 0.030817f
C1192 VTAIL.n96 VSUBS 0.01656f
C1193 VTAIL.n97 VSUBS 0.017534f
C1194 VTAIL.n98 VSUBS 0.039142f
C1195 VTAIL.n99 VSUBS 0.039142f
C1196 VTAIL.n100 VSUBS 0.039142f
C1197 VTAIL.n101 VSUBS 0.017047f
C1198 VTAIL.n102 VSUBS 0.01656f
C1199 VTAIL.n103 VSUBS 0.030817f
C1200 VTAIL.n104 VSUBS 0.030817f
C1201 VTAIL.n105 VSUBS 0.01656f
C1202 VTAIL.n106 VSUBS 0.017534f
C1203 VTAIL.n107 VSUBS 0.039142f
C1204 VTAIL.n108 VSUBS 0.095209f
C1205 VTAIL.n109 VSUBS 0.017534f
C1206 VTAIL.n110 VSUBS 0.01656f
C1207 VTAIL.n111 VSUBS 0.077127f
C1208 VTAIL.n112 VSUBS 0.048074f
C1209 VTAIL.n113 VSUBS 0.574522f
C1210 VTAIL.t9 VSUBS 0.245964f
C1211 VTAIL.t10 VSUBS 0.245964f
C1212 VTAIL.n114 VSUBS 1.72666f
C1213 VTAIL.n115 VSUBS 1.19512f
C1214 VTAIL.n116 VSUBS 0.033994f
C1215 VTAIL.n117 VSUBS 0.030817f
C1216 VTAIL.n118 VSUBS 0.01656f
C1217 VTAIL.n119 VSUBS 0.039142f
C1218 VTAIL.n120 VSUBS 0.017534f
C1219 VTAIL.n121 VSUBS 0.030817f
C1220 VTAIL.n122 VSUBS 0.017047f
C1221 VTAIL.n123 VSUBS 0.039142f
C1222 VTAIL.n124 VSUBS 0.01656f
C1223 VTAIL.n125 VSUBS 0.017534f
C1224 VTAIL.n126 VSUBS 0.030817f
C1225 VTAIL.n127 VSUBS 0.01656f
C1226 VTAIL.n128 VSUBS 0.039142f
C1227 VTAIL.n129 VSUBS 0.017534f
C1228 VTAIL.n130 VSUBS 0.030817f
C1229 VTAIL.n131 VSUBS 0.01656f
C1230 VTAIL.n132 VSUBS 0.029356f
C1231 VTAIL.n133 VSUBS 0.029444f
C1232 VTAIL.t7 VSUBS 0.084178f
C1233 VTAIL.n134 VSUBS 0.216256f
C1234 VTAIL.n135 VSUBS 1.25754f
C1235 VTAIL.n136 VSUBS 0.01656f
C1236 VTAIL.n137 VSUBS 0.017534f
C1237 VTAIL.n138 VSUBS 0.039142f
C1238 VTAIL.n139 VSUBS 0.039142f
C1239 VTAIL.n140 VSUBS 0.017534f
C1240 VTAIL.n141 VSUBS 0.01656f
C1241 VTAIL.n142 VSUBS 0.030817f
C1242 VTAIL.n143 VSUBS 0.030817f
C1243 VTAIL.n144 VSUBS 0.01656f
C1244 VTAIL.n145 VSUBS 0.017534f
C1245 VTAIL.n146 VSUBS 0.039142f
C1246 VTAIL.n147 VSUBS 0.039142f
C1247 VTAIL.n148 VSUBS 0.017534f
C1248 VTAIL.n149 VSUBS 0.01656f
C1249 VTAIL.n150 VSUBS 0.030817f
C1250 VTAIL.n151 VSUBS 0.030817f
C1251 VTAIL.n152 VSUBS 0.01656f
C1252 VTAIL.n153 VSUBS 0.017534f
C1253 VTAIL.n154 VSUBS 0.039142f
C1254 VTAIL.n155 VSUBS 0.039142f
C1255 VTAIL.n156 VSUBS 0.039142f
C1256 VTAIL.n157 VSUBS 0.017047f
C1257 VTAIL.n158 VSUBS 0.01656f
C1258 VTAIL.n159 VSUBS 0.030817f
C1259 VTAIL.n160 VSUBS 0.030817f
C1260 VTAIL.n161 VSUBS 0.01656f
C1261 VTAIL.n162 VSUBS 0.017534f
C1262 VTAIL.n163 VSUBS 0.039142f
C1263 VTAIL.n164 VSUBS 0.095209f
C1264 VTAIL.n165 VSUBS 0.017534f
C1265 VTAIL.n166 VSUBS 0.01656f
C1266 VTAIL.n167 VSUBS 0.077127f
C1267 VTAIL.n168 VSUBS 0.048074f
C1268 VTAIL.n169 VSUBS 1.97716f
C1269 VTAIL.n170 VSUBS 0.033994f
C1270 VTAIL.n171 VSUBS 0.030817f
C1271 VTAIL.n172 VSUBS 0.01656f
C1272 VTAIL.n173 VSUBS 0.039142f
C1273 VTAIL.n174 VSUBS 0.017534f
C1274 VTAIL.n175 VSUBS 0.030817f
C1275 VTAIL.n176 VSUBS 0.017047f
C1276 VTAIL.n177 VSUBS 0.039142f
C1277 VTAIL.n178 VSUBS 0.017534f
C1278 VTAIL.n179 VSUBS 0.030817f
C1279 VTAIL.n180 VSUBS 0.01656f
C1280 VTAIL.n181 VSUBS 0.039142f
C1281 VTAIL.n182 VSUBS 0.017534f
C1282 VTAIL.n183 VSUBS 0.030817f
C1283 VTAIL.n184 VSUBS 0.01656f
C1284 VTAIL.n185 VSUBS 0.029356f
C1285 VTAIL.n186 VSUBS 0.029444f
C1286 VTAIL.t1 VSUBS 0.084178f
C1287 VTAIL.n187 VSUBS 0.216256f
C1288 VTAIL.n188 VSUBS 1.25754f
C1289 VTAIL.n189 VSUBS 0.01656f
C1290 VTAIL.n190 VSUBS 0.017534f
C1291 VTAIL.n191 VSUBS 0.039142f
C1292 VTAIL.n192 VSUBS 0.039142f
C1293 VTAIL.n193 VSUBS 0.017534f
C1294 VTAIL.n194 VSUBS 0.01656f
C1295 VTAIL.n195 VSUBS 0.030817f
C1296 VTAIL.n196 VSUBS 0.030817f
C1297 VTAIL.n197 VSUBS 0.01656f
C1298 VTAIL.n198 VSUBS 0.017534f
C1299 VTAIL.n199 VSUBS 0.039142f
C1300 VTAIL.n200 VSUBS 0.039142f
C1301 VTAIL.n201 VSUBS 0.017534f
C1302 VTAIL.n202 VSUBS 0.01656f
C1303 VTAIL.n203 VSUBS 0.030817f
C1304 VTAIL.n204 VSUBS 0.030817f
C1305 VTAIL.n205 VSUBS 0.01656f
C1306 VTAIL.n206 VSUBS 0.01656f
C1307 VTAIL.n207 VSUBS 0.017534f
C1308 VTAIL.n208 VSUBS 0.039142f
C1309 VTAIL.n209 VSUBS 0.039142f
C1310 VTAIL.n210 VSUBS 0.039142f
C1311 VTAIL.n211 VSUBS 0.017047f
C1312 VTAIL.n212 VSUBS 0.01656f
C1313 VTAIL.n213 VSUBS 0.030817f
C1314 VTAIL.n214 VSUBS 0.030817f
C1315 VTAIL.n215 VSUBS 0.01656f
C1316 VTAIL.n216 VSUBS 0.017534f
C1317 VTAIL.n217 VSUBS 0.039142f
C1318 VTAIL.n218 VSUBS 0.095209f
C1319 VTAIL.n219 VSUBS 0.017534f
C1320 VTAIL.n220 VSUBS 0.01656f
C1321 VTAIL.n221 VSUBS 0.077127f
C1322 VTAIL.n222 VSUBS 0.048074f
C1323 VTAIL.n223 VSUBS 1.88834f
C1324 VP.t0 VSUBS 2.95793f
C1325 VP.n0 VSUBS 1.15941f
C1326 VP.n1 VSUBS 0.030442f
C1327 VP.n2 VSUBS 0.049306f
C1328 VP.n3 VSUBS 0.030442f
C1329 VP.n4 VSUBS 0.042517f
C1330 VP.n5 VSUBS 0.030442f
C1331 VP.n6 VSUBS 0.039199f
C1332 VP.n7 VSUBS 0.030442f
C1333 VP.n8 VSUBS 0.035829f
C1334 VP.t3 VSUBS 2.95793f
C1335 VP.n9 VSUBS 1.15941f
C1336 VP.n10 VSUBS 0.030442f
C1337 VP.n11 VSUBS 0.049306f
C1338 VP.n12 VSUBS 0.030442f
C1339 VP.n13 VSUBS 0.042517f
C1340 VP.t5 VSUBS 3.37026f
C1341 VP.t2 VSUBS 2.95793f
C1342 VP.n14 VSUBS 1.15182f
C1343 VP.n15 VSUBS 1.09459f
C1344 VP.n16 VSUBS 0.379413f
C1345 VP.n17 VSUBS 0.030442f
C1346 VP.n18 VSUBS 0.056452f
C1347 VP.n19 VSUBS 0.056452f
C1348 VP.n20 VSUBS 0.039199f
C1349 VP.n21 VSUBS 0.030442f
C1350 VP.n22 VSUBS 0.030442f
C1351 VP.n23 VSUBS 0.030442f
C1352 VP.n24 VSUBS 0.056452f
C1353 VP.n25 VSUBS 0.056452f
C1354 VP.n26 VSUBS 0.035829f
C1355 VP.n27 VSUBS 0.049125f
C1356 VP.n28 VSUBS 1.79345f
C1357 VP.t4 VSUBS 2.95793f
C1358 VP.n29 VSUBS 1.15941f
C1359 VP.n30 VSUBS 1.81496f
C1360 VP.n31 VSUBS 0.049125f
C1361 VP.n32 VSUBS 0.030442f
C1362 VP.n33 VSUBS 0.056452f
C1363 VP.n34 VSUBS 0.056452f
C1364 VP.n35 VSUBS 0.049306f
C1365 VP.n36 VSUBS 0.030442f
C1366 VP.n37 VSUBS 0.030442f
C1367 VP.n38 VSUBS 0.030442f
C1368 VP.n39 VSUBS 0.056452f
C1369 VP.n40 VSUBS 0.056452f
C1370 VP.t1 VSUBS 2.95793f
C1371 VP.n41 VSUBS 1.0475f
C1372 VP.n42 VSUBS 0.042517f
C1373 VP.n43 VSUBS 0.030442f
C1374 VP.n44 VSUBS 0.030442f
C1375 VP.n45 VSUBS 0.030442f
C1376 VP.n46 VSUBS 0.056452f
C1377 VP.n47 VSUBS 0.056452f
C1378 VP.n48 VSUBS 0.039199f
C1379 VP.n49 VSUBS 0.030442f
C1380 VP.n50 VSUBS 0.030442f
C1381 VP.n51 VSUBS 0.030442f
C1382 VP.n52 VSUBS 0.056452f
C1383 VP.n53 VSUBS 0.056452f
C1384 VP.n54 VSUBS 0.035829f
C1385 VP.n55 VSUBS 0.049125f
C1386 VP.n56 VSUBS 0.0861f
.ends

