* NGSPICE file created from diff_pair_sample_1669.ext - technology: sky130A

.subckt diff_pair_sample_1669 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=1.74
X1 VDD1.t5 VP.t0 VTAIL.t8 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=1.74
X2 VDD2.t5 VN.t0 VTAIL.t0 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=1.74
X3 B.t8 B.t6 B.t7 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=1.74
X4 VTAIL.t9 VP.t1 VDD1.t4 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=0.47685 ps=3.22 w=2.89 l=1.74
X5 VDD2.t4 VN.t1 VTAIL.t1 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=1.74
X6 VDD1.t3 VP.t2 VTAIL.t10 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=1.74
X7 B.t5 B.t3 B.t4 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=1.74
X8 VTAIL.t5 VN.t2 VDD2.t3 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=0.47685 ps=3.22 w=2.89 l=1.74
X9 VDD2.t2 VN.t3 VTAIL.t4 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=1.1271 ps=6.56 w=2.89 l=1.74
X10 VDD1.t2 VP.t3 VTAIL.t11 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=1.74
X11 VTAIL.t6 VP.t4 VDD1.t1 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=0.47685 ps=3.22 w=2.89 l=1.74
X12 VDD1.t0 VP.t5 VTAIL.t7 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=1.74
X13 B.t2 B.t0 B.t1 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0 ps=0 w=2.89 l=1.74
X14 VDD2.t1 VN.t4 VTAIL.t3 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=1.1271 pd=6.56 as=0.47685 ps=3.22 w=2.89 l=1.74
X15 VTAIL.t2 VN.t5 VDD2.t0 w_n2626_n1546# sky130_fd_pr__pfet_01v8 ad=0.47685 pd=3.22 as=0.47685 ps=3.22 w=2.89 l=1.74
R0 B.n220 B.n75 585
R1 B.n219 B.n218 585
R2 B.n217 B.n76 585
R3 B.n216 B.n215 585
R4 B.n214 B.n77 585
R5 B.n213 B.n212 585
R6 B.n211 B.n78 585
R7 B.n210 B.n209 585
R8 B.n208 B.n79 585
R9 B.n207 B.n206 585
R10 B.n205 B.n80 585
R11 B.n204 B.n203 585
R12 B.n202 B.n81 585
R13 B.n201 B.n200 585
R14 B.n199 B.n82 585
R15 B.n198 B.n197 585
R16 B.n193 B.n83 585
R17 B.n192 B.n191 585
R18 B.n190 B.n84 585
R19 B.n189 B.n188 585
R20 B.n187 B.n85 585
R21 B.n186 B.n185 585
R22 B.n184 B.n86 585
R23 B.n183 B.n182 585
R24 B.n180 B.n87 585
R25 B.n179 B.n178 585
R26 B.n177 B.n90 585
R27 B.n176 B.n175 585
R28 B.n174 B.n91 585
R29 B.n173 B.n172 585
R30 B.n171 B.n92 585
R31 B.n170 B.n169 585
R32 B.n168 B.n93 585
R33 B.n167 B.n166 585
R34 B.n165 B.n94 585
R35 B.n164 B.n163 585
R36 B.n162 B.n95 585
R37 B.n161 B.n160 585
R38 B.n159 B.n96 585
R39 B.n222 B.n221 585
R40 B.n223 B.n74 585
R41 B.n225 B.n224 585
R42 B.n226 B.n73 585
R43 B.n228 B.n227 585
R44 B.n229 B.n72 585
R45 B.n231 B.n230 585
R46 B.n232 B.n71 585
R47 B.n234 B.n233 585
R48 B.n235 B.n70 585
R49 B.n237 B.n236 585
R50 B.n238 B.n69 585
R51 B.n240 B.n239 585
R52 B.n241 B.n68 585
R53 B.n243 B.n242 585
R54 B.n244 B.n67 585
R55 B.n246 B.n245 585
R56 B.n247 B.n66 585
R57 B.n249 B.n248 585
R58 B.n250 B.n65 585
R59 B.n252 B.n251 585
R60 B.n253 B.n64 585
R61 B.n255 B.n254 585
R62 B.n256 B.n63 585
R63 B.n258 B.n257 585
R64 B.n259 B.n62 585
R65 B.n261 B.n260 585
R66 B.n262 B.n61 585
R67 B.n264 B.n263 585
R68 B.n265 B.n60 585
R69 B.n267 B.n266 585
R70 B.n268 B.n59 585
R71 B.n270 B.n269 585
R72 B.n271 B.n58 585
R73 B.n273 B.n272 585
R74 B.n274 B.n57 585
R75 B.n276 B.n275 585
R76 B.n277 B.n56 585
R77 B.n279 B.n278 585
R78 B.n280 B.n55 585
R79 B.n282 B.n281 585
R80 B.n283 B.n54 585
R81 B.n285 B.n284 585
R82 B.n286 B.n53 585
R83 B.n288 B.n287 585
R84 B.n289 B.n52 585
R85 B.n291 B.n290 585
R86 B.n292 B.n51 585
R87 B.n294 B.n293 585
R88 B.n295 B.n50 585
R89 B.n297 B.n296 585
R90 B.n298 B.n49 585
R91 B.n300 B.n299 585
R92 B.n301 B.n48 585
R93 B.n303 B.n302 585
R94 B.n304 B.n47 585
R95 B.n306 B.n305 585
R96 B.n307 B.n46 585
R97 B.n309 B.n308 585
R98 B.n310 B.n45 585
R99 B.n312 B.n311 585
R100 B.n313 B.n44 585
R101 B.n315 B.n314 585
R102 B.n316 B.n43 585
R103 B.n318 B.n317 585
R104 B.n319 B.n42 585
R105 B.n379 B.n18 585
R106 B.n378 B.n377 585
R107 B.n376 B.n19 585
R108 B.n375 B.n374 585
R109 B.n373 B.n20 585
R110 B.n372 B.n371 585
R111 B.n370 B.n21 585
R112 B.n369 B.n368 585
R113 B.n367 B.n22 585
R114 B.n366 B.n365 585
R115 B.n364 B.n23 585
R116 B.n363 B.n362 585
R117 B.n361 B.n24 585
R118 B.n360 B.n359 585
R119 B.n358 B.n25 585
R120 B.n356 B.n355 585
R121 B.n354 B.n28 585
R122 B.n353 B.n352 585
R123 B.n351 B.n29 585
R124 B.n350 B.n349 585
R125 B.n348 B.n30 585
R126 B.n347 B.n346 585
R127 B.n345 B.n31 585
R128 B.n344 B.n343 585
R129 B.n342 B.n341 585
R130 B.n340 B.n35 585
R131 B.n339 B.n338 585
R132 B.n337 B.n36 585
R133 B.n336 B.n335 585
R134 B.n334 B.n37 585
R135 B.n333 B.n332 585
R136 B.n331 B.n38 585
R137 B.n330 B.n329 585
R138 B.n328 B.n39 585
R139 B.n327 B.n326 585
R140 B.n325 B.n40 585
R141 B.n324 B.n323 585
R142 B.n322 B.n41 585
R143 B.n321 B.n320 585
R144 B.n381 B.n380 585
R145 B.n382 B.n17 585
R146 B.n384 B.n383 585
R147 B.n385 B.n16 585
R148 B.n387 B.n386 585
R149 B.n388 B.n15 585
R150 B.n390 B.n389 585
R151 B.n391 B.n14 585
R152 B.n393 B.n392 585
R153 B.n394 B.n13 585
R154 B.n396 B.n395 585
R155 B.n397 B.n12 585
R156 B.n399 B.n398 585
R157 B.n400 B.n11 585
R158 B.n402 B.n401 585
R159 B.n403 B.n10 585
R160 B.n405 B.n404 585
R161 B.n406 B.n9 585
R162 B.n408 B.n407 585
R163 B.n409 B.n8 585
R164 B.n411 B.n410 585
R165 B.n412 B.n7 585
R166 B.n414 B.n413 585
R167 B.n415 B.n6 585
R168 B.n417 B.n416 585
R169 B.n418 B.n5 585
R170 B.n420 B.n419 585
R171 B.n421 B.n4 585
R172 B.n423 B.n422 585
R173 B.n424 B.n3 585
R174 B.n426 B.n425 585
R175 B.n427 B.n0 585
R176 B.n2 B.n1 585
R177 B.n113 B.n112 585
R178 B.n114 B.n111 585
R179 B.n116 B.n115 585
R180 B.n117 B.n110 585
R181 B.n119 B.n118 585
R182 B.n120 B.n109 585
R183 B.n122 B.n121 585
R184 B.n123 B.n108 585
R185 B.n125 B.n124 585
R186 B.n126 B.n107 585
R187 B.n128 B.n127 585
R188 B.n129 B.n106 585
R189 B.n131 B.n130 585
R190 B.n132 B.n105 585
R191 B.n134 B.n133 585
R192 B.n135 B.n104 585
R193 B.n137 B.n136 585
R194 B.n138 B.n103 585
R195 B.n140 B.n139 585
R196 B.n141 B.n102 585
R197 B.n143 B.n142 585
R198 B.n144 B.n101 585
R199 B.n146 B.n145 585
R200 B.n147 B.n100 585
R201 B.n149 B.n148 585
R202 B.n150 B.n99 585
R203 B.n152 B.n151 585
R204 B.n153 B.n98 585
R205 B.n155 B.n154 585
R206 B.n156 B.n97 585
R207 B.n158 B.n157 585
R208 B.n159 B.n158 511.721
R209 B.n222 B.n75 511.721
R210 B.n320 B.n319 511.721
R211 B.n380 B.n379 511.721
R212 B.n429 B.n428 256.663
R213 B.n88 B.t6 246.262
R214 B.n194 B.t0 246.262
R215 B.n32 B.t3 246.262
R216 B.n26 B.t9 246.262
R217 B.n428 B.n427 235.042
R218 B.n428 B.n2 235.042
R219 B.n194 B.t1 183.648
R220 B.n32 B.t5 183.648
R221 B.n88 B.t7 183.645
R222 B.n26 B.t11 183.645
R223 B.n160 B.n159 163.367
R224 B.n160 B.n95 163.367
R225 B.n164 B.n95 163.367
R226 B.n165 B.n164 163.367
R227 B.n166 B.n165 163.367
R228 B.n166 B.n93 163.367
R229 B.n170 B.n93 163.367
R230 B.n171 B.n170 163.367
R231 B.n172 B.n171 163.367
R232 B.n172 B.n91 163.367
R233 B.n176 B.n91 163.367
R234 B.n177 B.n176 163.367
R235 B.n178 B.n177 163.367
R236 B.n178 B.n87 163.367
R237 B.n183 B.n87 163.367
R238 B.n184 B.n183 163.367
R239 B.n185 B.n184 163.367
R240 B.n185 B.n85 163.367
R241 B.n189 B.n85 163.367
R242 B.n190 B.n189 163.367
R243 B.n191 B.n190 163.367
R244 B.n191 B.n83 163.367
R245 B.n198 B.n83 163.367
R246 B.n199 B.n198 163.367
R247 B.n200 B.n199 163.367
R248 B.n200 B.n81 163.367
R249 B.n204 B.n81 163.367
R250 B.n205 B.n204 163.367
R251 B.n206 B.n205 163.367
R252 B.n206 B.n79 163.367
R253 B.n210 B.n79 163.367
R254 B.n211 B.n210 163.367
R255 B.n212 B.n211 163.367
R256 B.n212 B.n77 163.367
R257 B.n216 B.n77 163.367
R258 B.n217 B.n216 163.367
R259 B.n218 B.n217 163.367
R260 B.n218 B.n75 163.367
R261 B.n319 B.n318 163.367
R262 B.n318 B.n43 163.367
R263 B.n314 B.n43 163.367
R264 B.n314 B.n313 163.367
R265 B.n313 B.n312 163.367
R266 B.n312 B.n45 163.367
R267 B.n308 B.n45 163.367
R268 B.n308 B.n307 163.367
R269 B.n307 B.n306 163.367
R270 B.n306 B.n47 163.367
R271 B.n302 B.n47 163.367
R272 B.n302 B.n301 163.367
R273 B.n301 B.n300 163.367
R274 B.n300 B.n49 163.367
R275 B.n296 B.n49 163.367
R276 B.n296 B.n295 163.367
R277 B.n295 B.n294 163.367
R278 B.n294 B.n51 163.367
R279 B.n290 B.n51 163.367
R280 B.n290 B.n289 163.367
R281 B.n289 B.n288 163.367
R282 B.n288 B.n53 163.367
R283 B.n284 B.n53 163.367
R284 B.n284 B.n283 163.367
R285 B.n283 B.n282 163.367
R286 B.n282 B.n55 163.367
R287 B.n278 B.n55 163.367
R288 B.n278 B.n277 163.367
R289 B.n277 B.n276 163.367
R290 B.n276 B.n57 163.367
R291 B.n272 B.n57 163.367
R292 B.n272 B.n271 163.367
R293 B.n271 B.n270 163.367
R294 B.n270 B.n59 163.367
R295 B.n266 B.n59 163.367
R296 B.n266 B.n265 163.367
R297 B.n265 B.n264 163.367
R298 B.n264 B.n61 163.367
R299 B.n260 B.n61 163.367
R300 B.n260 B.n259 163.367
R301 B.n259 B.n258 163.367
R302 B.n258 B.n63 163.367
R303 B.n254 B.n63 163.367
R304 B.n254 B.n253 163.367
R305 B.n253 B.n252 163.367
R306 B.n252 B.n65 163.367
R307 B.n248 B.n65 163.367
R308 B.n248 B.n247 163.367
R309 B.n247 B.n246 163.367
R310 B.n246 B.n67 163.367
R311 B.n242 B.n67 163.367
R312 B.n242 B.n241 163.367
R313 B.n241 B.n240 163.367
R314 B.n240 B.n69 163.367
R315 B.n236 B.n69 163.367
R316 B.n236 B.n235 163.367
R317 B.n235 B.n234 163.367
R318 B.n234 B.n71 163.367
R319 B.n230 B.n71 163.367
R320 B.n230 B.n229 163.367
R321 B.n229 B.n228 163.367
R322 B.n228 B.n73 163.367
R323 B.n224 B.n73 163.367
R324 B.n224 B.n223 163.367
R325 B.n223 B.n222 163.367
R326 B.n379 B.n378 163.367
R327 B.n378 B.n19 163.367
R328 B.n374 B.n19 163.367
R329 B.n374 B.n373 163.367
R330 B.n373 B.n372 163.367
R331 B.n372 B.n21 163.367
R332 B.n368 B.n21 163.367
R333 B.n368 B.n367 163.367
R334 B.n367 B.n366 163.367
R335 B.n366 B.n23 163.367
R336 B.n362 B.n23 163.367
R337 B.n362 B.n361 163.367
R338 B.n361 B.n360 163.367
R339 B.n360 B.n25 163.367
R340 B.n355 B.n25 163.367
R341 B.n355 B.n354 163.367
R342 B.n354 B.n353 163.367
R343 B.n353 B.n29 163.367
R344 B.n349 B.n29 163.367
R345 B.n349 B.n348 163.367
R346 B.n348 B.n347 163.367
R347 B.n347 B.n31 163.367
R348 B.n343 B.n31 163.367
R349 B.n343 B.n342 163.367
R350 B.n342 B.n35 163.367
R351 B.n338 B.n35 163.367
R352 B.n338 B.n337 163.367
R353 B.n337 B.n336 163.367
R354 B.n336 B.n37 163.367
R355 B.n332 B.n37 163.367
R356 B.n332 B.n331 163.367
R357 B.n331 B.n330 163.367
R358 B.n330 B.n39 163.367
R359 B.n326 B.n39 163.367
R360 B.n326 B.n325 163.367
R361 B.n325 B.n324 163.367
R362 B.n324 B.n41 163.367
R363 B.n320 B.n41 163.367
R364 B.n380 B.n17 163.367
R365 B.n384 B.n17 163.367
R366 B.n385 B.n384 163.367
R367 B.n386 B.n385 163.367
R368 B.n386 B.n15 163.367
R369 B.n390 B.n15 163.367
R370 B.n391 B.n390 163.367
R371 B.n392 B.n391 163.367
R372 B.n392 B.n13 163.367
R373 B.n396 B.n13 163.367
R374 B.n397 B.n396 163.367
R375 B.n398 B.n397 163.367
R376 B.n398 B.n11 163.367
R377 B.n402 B.n11 163.367
R378 B.n403 B.n402 163.367
R379 B.n404 B.n403 163.367
R380 B.n404 B.n9 163.367
R381 B.n408 B.n9 163.367
R382 B.n409 B.n408 163.367
R383 B.n410 B.n409 163.367
R384 B.n410 B.n7 163.367
R385 B.n414 B.n7 163.367
R386 B.n415 B.n414 163.367
R387 B.n416 B.n415 163.367
R388 B.n416 B.n5 163.367
R389 B.n420 B.n5 163.367
R390 B.n421 B.n420 163.367
R391 B.n422 B.n421 163.367
R392 B.n422 B.n3 163.367
R393 B.n426 B.n3 163.367
R394 B.n427 B.n426 163.367
R395 B.n112 B.n2 163.367
R396 B.n112 B.n111 163.367
R397 B.n116 B.n111 163.367
R398 B.n117 B.n116 163.367
R399 B.n118 B.n117 163.367
R400 B.n118 B.n109 163.367
R401 B.n122 B.n109 163.367
R402 B.n123 B.n122 163.367
R403 B.n124 B.n123 163.367
R404 B.n124 B.n107 163.367
R405 B.n128 B.n107 163.367
R406 B.n129 B.n128 163.367
R407 B.n130 B.n129 163.367
R408 B.n130 B.n105 163.367
R409 B.n134 B.n105 163.367
R410 B.n135 B.n134 163.367
R411 B.n136 B.n135 163.367
R412 B.n136 B.n103 163.367
R413 B.n140 B.n103 163.367
R414 B.n141 B.n140 163.367
R415 B.n142 B.n141 163.367
R416 B.n142 B.n101 163.367
R417 B.n146 B.n101 163.367
R418 B.n147 B.n146 163.367
R419 B.n148 B.n147 163.367
R420 B.n148 B.n99 163.367
R421 B.n152 B.n99 163.367
R422 B.n153 B.n152 163.367
R423 B.n154 B.n153 163.367
R424 B.n154 B.n97 163.367
R425 B.n158 B.n97 163.367
R426 B.n195 B.t2 143.501
R427 B.n33 B.t4 143.501
R428 B.n89 B.t8 143.5
R429 B.n27 B.t10 143.5
R430 B.n181 B.n89 59.5399
R431 B.n196 B.n195 59.5399
R432 B.n34 B.n33 59.5399
R433 B.n357 B.n27 59.5399
R434 B.n89 B.n88 40.146
R435 B.n195 B.n194 40.146
R436 B.n33 B.n32 40.146
R437 B.n27 B.n26 40.146
R438 B.n381 B.n18 33.2493
R439 B.n321 B.n42 33.2493
R440 B.n221 B.n220 33.2493
R441 B.n157 B.n96 33.2493
R442 B B.n429 18.0485
R443 B.n382 B.n381 10.6151
R444 B.n383 B.n382 10.6151
R445 B.n383 B.n16 10.6151
R446 B.n387 B.n16 10.6151
R447 B.n388 B.n387 10.6151
R448 B.n389 B.n388 10.6151
R449 B.n389 B.n14 10.6151
R450 B.n393 B.n14 10.6151
R451 B.n394 B.n393 10.6151
R452 B.n395 B.n394 10.6151
R453 B.n395 B.n12 10.6151
R454 B.n399 B.n12 10.6151
R455 B.n400 B.n399 10.6151
R456 B.n401 B.n400 10.6151
R457 B.n401 B.n10 10.6151
R458 B.n405 B.n10 10.6151
R459 B.n406 B.n405 10.6151
R460 B.n407 B.n406 10.6151
R461 B.n407 B.n8 10.6151
R462 B.n411 B.n8 10.6151
R463 B.n412 B.n411 10.6151
R464 B.n413 B.n412 10.6151
R465 B.n413 B.n6 10.6151
R466 B.n417 B.n6 10.6151
R467 B.n418 B.n417 10.6151
R468 B.n419 B.n418 10.6151
R469 B.n419 B.n4 10.6151
R470 B.n423 B.n4 10.6151
R471 B.n424 B.n423 10.6151
R472 B.n425 B.n424 10.6151
R473 B.n425 B.n0 10.6151
R474 B.n377 B.n18 10.6151
R475 B.n377 B.n376 10.6151
R476 B.n376 B.n375 10.6151
R477 B.n375 B.n20 10.6151
R478 B.n371 B.n20 10.6151
R479 B.n371 B.n370 10.6151
R480 B.n370 B.n369 10.6151
R481 B.n369 B.n22 10.6151
R482 B.n365 B.n22 10.6151
R483 B.n365 B.n364 10.6151
R484 B.n364 B.n363 10.6151
R485 B.n363 B.n24 10.6151
R486 B.n359 B.n24 10.6151
R487 B.n359 B.n358 10.6151
R488 B.n356 B.n28 10.6151
R489 B.n352 B.n28 10.6151
R490 B.n352 B.n351 10.6151
R491 B.n351 B.n350 10.6151
R492 B.n350 B.n30 10.6151
R493 B.n346 B.n30 10.6151
R494 B.n346 B.n345 10.6151
R495 B.n345 B.n344 10.6151
R496 B.n341 B.n340 10.6151
R497 B.n340 B.n339 10.6151
R498 B.n339 B.n36 10.6151
R499 B.n335 B.n36 10.6151
R500 B.n335 B.n334 10.6151
R501 B.n334 B.n333 10.6151
R502 B.n333 B.n38 10.6151
R503 B.n329 B.n38 10.6151
R504 B.n329 B.n328 10.6151
R505 B.n328 B.n327 10.6151
R506 B.n327 B.n40 10.6151
R507 B.n323 B.n40 10.6151
R508 B.n323 B.n322 10.6151
R509 B.n322 B.n321 10.6151
R510 B.n317 B.n42 10.6151
R511 B.n317 B.n316 10.6151
R512 B.n316 B.n315 10.6151
R513 B.n315 B.n44 10.6151
R514 B.n311 B.n44 10.6151
R515 B.n311 B.n310 10.6151
R516 B.n310 B.n309 10.6151
R517 B.n309 B.n46 10.6151
R518 B.n305 B.n46 10.6151
R519 B.n305 B.n304 10.6151
R520 B.n304 B.n303 10.6151
R521 B.n303 B.n48 10.6151
R522 B.n299 B.n48 10.6151
R523 B.n299 B.n298 10.6151
R524 B.n298 B.n297 10.6151
R525 B.n297 B.n50 10.6151
R526 B.n293 B.n50 10.6151
R527 B.n293 B.n292 10.6151
R528 B.n292 B.n291 10.6151
R529 B.n291 B.n52 10.6151
R530 B.n287 B.n52 10.6151
R531 B.n287 B.n286 10.6151
R532 B.n286 B.n285 10.6151
R533 B.n285 B.n54 10.6151
R534 B.n281 B.n54 10.6151
R535 B.n281 B.n280 10.6151
R536 B.n280 B.n279 10.6151
R537 B.n279 B.n56 10.6151
R538 B.n275 B.n56 10.6151
R539 B.n275 B.n274 10.6151
R540 B.n274 B.n273 10.6151
R541 B.n273 B.n58 10.6151
R542 B.n269 B.n58 10.6151
R543 B.n269 B.n268 10.6151
R544 B.n268 B.n267 10.6151
R545 B.n267 B.n60 10.6151
R546 B.n263 B.n60 10.6151
R547 B.n263 B.n262 10.6151
R548 B.n262 B.n261 10.6151
R549 B.n261 B.n62 10.6151
R550 B.n257 B.n62 10.6151
R551 B.n257 B.n256 10.6151
R552 B.n256 B.n255 10.6151
R553 B.n255 B.n64 10.6151
R554 B.n251 B.n64 10.6151
R555 B.n251 B.n250 10.6151
R556 B.n250 B.n249 10.6151
R557 B.n249 B.n66 10.6151
R558 B.n245 B.n66 10.6151
R559 B.n245 B.n244 10.6151
R560 B.n244 B.n243 10.6151
R561 B.n243 B.n68 10.6151
R562 B.n239 B.n68 10.6151
R563 B.n239 B.n238 10.6151
R564 B.n238 B.n237 10.6151
R565 B.n237 B.n70 10.6151
R566 B.n233 B.n70 10.6151
R567 B.n233 B.n232 10.6151
R568 B.n232 B.n231 10.6151
R569 B.n231 B.n72 10.6151
R570 B.n227 B.n72 10.6151
R571 B.n227 B.n226 10.6151
R572 B.n226 B.n225 10.6151
R573 B.n225 B.n74 10.6151
R574 B.n221 B.n74 10.6151
R575 B.n113 B.n1 10.6151
R576 B.n114 B.n113 10.6151
R577 B.n115 B.n114 10.6151
R578 B.n115 B.n110 10.6151
R579 B.n119 B.n110 10.6151
R580 B.n120 B.n119 10.6151
R581 B.n121 B.n120 10.6151
R582 B.n121 B.n108 10.6151
R583 B.n125 B.n108 10.6151
R584 B.n126 B.n125 10.6151
R585 B.n127 B.n126 10.6151
R586 B.n127 B.n106 10.6151
R587 B.n131 B.n106 10.6151
R588 B.n132 B.n131 10.6151
R589 B.n133 B.n132 10.6151
R590 B.n133 B.n104 10.6151
R591 B.n137 B.n104 10.6151
R592 B.n138 B.n137 10.6151
R593 B.n139 B.n138 10.6151
R594 B.n139 B.n102 10.6151
R595 B.n143 B.n102 10.6151
R596 B.n144 B.n143 10.6151
R597 B.n145 B.n144 10.6151
R598 B.n145 B.n100 10.6151
R599 B.n149 B.n100 10.6151
R600 B.n150 B.n149 10.6151
R601 B.n151 B.n150 10.6151
R602 B.n151 B.n98 10.6151
R603 B.n155 B.n98 10.6151
R604 B.n156 B.n155 10.6151
R605 B.n157 B.n156 10.6151
R606 B.n161 B.n96 10.6151
R607 B.n162 B.n161 10.6151
R608 B.n163 B.n162 10.6151
R609 B.n163 B.n94 10.6151
R610 B.n167 B.n94 10.6151
R611 B.n168 B.n167 10.6151
R612 B.n169 B.n168 10.6151
R613 B.n169 B.n92 10.6151
R614 B.n173 B.n92 10.6151
R615 B.n174 B.n173 10.6151
R616 B.n175 B.n174 10.6151
R617 B.n175 B.n90 10.6151
R618 B.n179 B.n90 10.6151
R619 B.n180 B.n179 10.6151
R620 B.n182 B.n86 10.6151
R621 B.n186 B.n86 10.6151
R622 B.n187 B.n186 10.6151
R623 B.n188 B.n187 10.6151
R624 B.n188 B.n84 10.6151
R625 B.n192 B.n84 10.6151
R626 B.n193 B.n192 10.6151
R627 B.n197 B.n193 10.6151
R628 B.n201 B.n82 10.6151
R629 B.n202 B.n201 10.6151
R630 B.n203 B.n202 10.6151
R631 B.n203 B.n80 10.6151
R632 B.n207 B.n80 10.6151
R633 B.n208 B.n207 10.6151
R634 B.n209 B.n208 10.6151
R635 B.n209 B.n78 10.6151
R636 B.n213 B.n78 10.6151
R637 B.n214 B.n213 10.6151
R638 B.n215 B.n214 10.6151
R639 B.n215 B.n76 10.6151
R640 B.n219 B.n76 10.6151
R641 B.n220 B.n219 10.6151
R642 B.n429 B.n0 8.11757
R643 B.n429 B.n1 8.11757
R644 B.n357 B.n356 6.5566
R645 B.n344 B.n34 6.5566
R646 B.n182 B.n181 6.5566
R647 B.n197 B.n196 6.5566
R648 B.n358 B.n357 4.05904
R649 B.n341 B.n34 4.05904
R650 B.n181 B.n180 4.05904
R651 B.n196 B.n82 4.05904
R652 VP.n18 VP.n17 182.343
R653 VP.n33 VP.n32 182.343
R654 VP.n16 VP.n15 182.343
R655 VP.n10 VP.n9 161.3
R656 VP.n11 VP.n6 161.3
R657 VP.n13 VP.n12 161.3
R658 VP.n14 VP.n5 161.3
R659 VP.n31 VP.n0 161.3
R660 VP.n30 VP.n29 161.3
R661 VP.n28 VP.n1 161.3
R662 VP.n27 VP.n26 161.3
R663 VP.n25 VP.n2 161.3
R664 VP.n24 VP.n23 161.3
R665 VP.n22 VP.n3 161.3
R666 VP.n21 VP.n20 161.3
R667 VP.n19 VP.n4 161.3
R668 VP.n7 VP.t5 74.47
R669 VP.n8 VP.n7 44.5658
R670 VP.n20 VP.n3 43.8928
R671 VP.n30 VP.n1 43.8928
R672 VP.n13 VP.n6 43.8928
R673 VP.n25 VP.t4 40.0287
R674 VP.n18 VP.t3 40.0287
R675 VP.n32 VP.t0 40.0287
R676 VP.n8 VP.t1 40.0287
R677 VP.n15 VP.t2 40.0287
R678 VP.n17 VP.n16 38.2846
R679 VP.n24 VP.n3 37.094
R680 VP.n26 VP.n1 37.094
R681 VP.n9 VP.n6 37.094
R682 VP.n20 VP.n19 24.4675
R683 VP.n25 VP.n24 24.4675
R684 VP.n26 VP.n25 24.4675
R685 VP.n31 VP.n30 24.4675
R686 VP.n14 VP.n13 24.4675
R687 VP.n9 VP.n8 24.4675
R688 VP.n10 VP.n7 12.3021
R689 VP.n19 VP.n18 3.42588
R690 VP.n32 VP.n31 3.42588
R691 VP.n15 VP.n14 3.42588
R692 VP.n11 VP.n10 0.189894
R693 VP.n12 VP.n11 0.189894
R694 VP.n12 VP.n5 0.189894
R695 VP.n16 VP.n5 0.189894
R696 VP.n17 VP.n4 0.189894
R697 VP.n21 VP.n4 0.189894
R698 VP.n22 VP.n21 0.189894
R699 VP.n23 VP.n22 0.189894
R700 VP.n23 VP.n2 0.189894
R701 VP.n27 VP.n2 0.189894
R702 VP.n28 VP.n27 0.189894
R703 VP.n29 VP.n28 0.189894
R704 VP.n29 VP.n0 0.189894
R705 VP.n33 VP.n0 0.189894
R706 VP VP.n33 0.0516364
R707 VTAIL.n7 VTAIL.t1 135.161
R708 VTAIL.n10 VTAIL.t10 135.16
R709 VTAIL.n11 VTAIL.t4 135.16
R710 VTAIL.n2 VTAIL.t8 135.16
R711 VTAIL.n9 VTAIL.n8 123.912
R712 VTAIL.n6 VTAIL.n5 123.912
R713 VTAIL.n1 VTAIL.n0 123.912
R714 VTAIL.n4 VTAIL.n3 123.912
R715 VTAIL.n6 VTAIL.n4 18.4272
R716 VTAIL.n11 VTAIL.n10 16.6427
R717 VTAIL.n0 VTAIL.t0 11.2479
R718 VTAIL.n0 VTAIL.t2 11.2479
R719 VTAIL.n3 VTAIL.t11 11.2479
R720 VTAIL.n3 VTAIL.t6 11.2479
R721 VTAIL.n8 VTAIL.t7 11.2479
R722 VTAIL.n8 VTAIL.t9 11.2479
R723 VTAIL.n5 VTAIL.t3 11.2479
R724 VTAIL.n5 VTAIL.t5 11.2479
R725 VTAIL.n7 VTAIL.n6 1.78498
R726 VTAIL.n10 VTAIL.n9 1.78498
R727 VTAIL.n4 VTAIL.n2 1.78498
R728 VTAIL.n9 VTAIL.n7 1.36257
R729 VTAIL.n2 VTAIL.n1 1.36257
R730 VTAIL VTAIL.n11 1.28067
R731 VTAIL VTAIL.n1 0.50481
R732 VDD1 VDD1.t0 153.236
R733 VDD1.n1 VDD1.t2 153.121
R734 VDD1.n1 VDD1.n0 140.982
R735 VDD1.n3 VDD1.n2 140.591
R736 VDD1.n3 VDD1.n1 33.4815
R737 VDD1.n2 VDD1.t4 11.2479
R738 VDD1.n2 VDD1.t3 11.2479
R739 VDD1.n0 VDD1.t1 11.2479
R740 VDD1.n0 VDD1.t5 11.2479
R741 VDD1 VDD1.n3 0.388431
R742 VN.n11 VN.n10 182.343
R743 VN.n23 VN.n22 182.343
R744 VN.n21 VN.n12 161.3
R745 VN.n20 VN.n19 161.3
R746 VN.n18 VN.n13 161.3
R747 VN.n17 VN.n16 161.3
R748 VN.n9 VN.n0 161.3
R749 VN.n8 VN.n7 161.3
R750 VN.n6 VN.n1 161.3
R751 VN.n5 VN.n4 161.3
R752 VN.n2 VN.t0 74.47
R753 VN.n14 VN.t1 74.47
R754 VN.n15 VN.n14 44.5658
R755 VN.n3 VN.n2 44.5658
R756 VN.n8 VN.n1 43.8928
R757 VN.n20 VN.n13 43.8928
R758 VN.n3 VN.t5 40.0287
R759 VN.n10 VN.t3 40.0287
R760 VN.n15 VN.t2 40.0287
R761 VN.n22 VN.t4 40.0287
R762 VN VN.n23 38.6653
R763 VN.n4 VN.n1 37.094
R764 VN.n16 VN.n13 37.094
R765 VN.n4 VN.n3 24.4675
R766 VN.n9 VN.n8 24.4675
R767 VN.n16 VN.n15 24.4675
R768 VN.n21 VN.n20 24.4675
R769 VN.n17 VN.n14 12.3021
R770 VN.n5 VN.n2 12.3021
R771 VN.n10 VN.n9 3.42588
R772 VN.n22 VN.n21 3.42588
R773 VN.n23 VN.n12 0.189894
R774 VN.n19 VN.n12 0.189894
R775 VN.n19 VN.n18 0.189894
R776 VN.n18 VN.n17 0.189894
R777 VN.n6 VN.n5 0.189894
R778 VN.n7 VN.n6 0.189894
R779 VN.n7 VN.n0 0.189894
R780 VN.n11 VN.n0 0.189894
R781 VN VN.n11 0.0516364
R782 VDD2.n1 VDD2.t5 153.121
R783 VDD2.n2 VDD2.t1 151.839
R784 VDD2.n1 VDD2.n0 140.982
R785 VDD2 VDD2.n3 140.98
R786 VDD2.n2 VDD2.n1 32.0062
R787 VDD2.n3 VDD2.t3 11.2479
R788 VDD2.n3 VDD2.t4 11.2479
R789 VDD2.n0 VDD2.t0 11.2479
R790 VDD2.n0 VDD2.t2 11.2479
R791 VDD2 VDD2.n2 1.39705
C0 VN B 0.875733f
C1 VDD2 VN 1.7616f
C2 VDD1 VTAIL 3.92447f
C3 VDD2 B 1.21322f
C4 VDD1 VP 1.99506f
C5 VDD1 w_n2626_n1546# 1.42849f
C6 VN VTAIL 2.24979f
C7 VP VN 4.41086f
C8 B VTAIL 1.3667f
C9 VDD2 VTAIL 3.97134f
C10 w_n2626_n1546# VN 4.59168f
C11 VP B 1.43379f
C12 VP VDD2 0.390259f
C13 w_n2626_n1546# B 5.94829f
C14 w_n2626_n1546# VDD2 1.48546f
C15 VDD1 VN 0.154655f
C16 VDD1 B 1.15954f
C17 VP VTAIL 2.26396f
C18 VDD1 VDD2 1.09523f
C19 w_n2626_n1546# VTAIL 1.56181f
C20 VP w_n2626_n1546# 4.92628f
C21 VDD2 VSUBS 0.894515f
C22 VDD1 VSUBS 1.248811f
C23 VTAIL VSUBS 0.460945f
C24 VN VSUBS 4.48132f
C25 VP VSUBS 1.75229f
C26 B VSUBS 2.855784f
C27 w_n2626_n1546# VSUBS 51.459103f
C28 VDD2.t5 VSUBS 0.266585f
C29 VDD2.t0 VSUBS 0.035753f
C30 VDD2.t2 VSUBS 0.035753f
C31 VDD2.n0 VSUBS 0.185831f
C32 VDD2.n1 VSUBS 1.36204f
C33 VDD2.t1 VSUBS 0.2642f
C34 VDD2.n2 VSUBS 1.19238f
C35 VDD2.t3 VSUBS 0.035753f
C36 VDD2.t4 VSUBS 0.035753f
C37 VDD2.n3 VSUBS 0.185822f
C38 VN.n0 VSUBS 0.047308f
C39 VN.t3 VSUBS 0.589794f
C40 VN.n1 VSUBS 0.038996f
C41 VN.t0 VSUBS 0.813657f
C42 VN.n2 VSUBS 0.349028f
C43 VN.t5 VSUBS 0.589794f
C44 VN.n3 VSUBS 0.391764f
C45 VN.n4 VSUBS 0.095283f
C46 VN.n5 VSUBS 0.345944f
C47 VN.n6 VSUBS 0.047308f
C48 VN.n7 VSUBS 0.047308f
C49 VN.n8 VSUBS 0.092024f
C50 VN.n9 VSUBS 0.050735f
C51 VN.n10 VSUBS 0.367631f
C52 VN.n11 VSUBS 0.049951f
C53 VN.n12 VSUBS 0.047308f
C54 VN.t4 VSUBS 0.589794f
C55 VN.n13 VSUBS 0.038996f
C56 VN.t1 VSUBS 0.813657f
C57 VN.n14 VSUBS 0.349028f
C58 VN.t2 VSUBS 0.589794f
C59 VN.n15 VSUBS 0.391764f
C60 VN.n16 VSUBS 0.095283f
C61 VN.n17 VSUBS 0.345944f
C62 VN.n18 VSUBS 0.047308f
C63 VN.n19 VSUBS 0.047308f
C64 VN.n20 VSUBS 0.092024f
C65 VN.n21 VSUBS 0.050735f
C66 VN.n22 VSUBS 0.367631f
C67 VN.n23 VSUBS 1.70921f
C68 VDD1.t0 VSUBS 0.256466f
C69 VDD1.t2 VSUBS 0.256217f
C70 VDD1.t1 VSUBS 0.034363f
C71 VDD1.t5 VSUBS 0.034363f
C72 VDD1.n0 VSUBS 0.178604f
C73 VDD1.n1 VSUBS 1.36598f
C74 VDD1.t4 VSUBS 0.034363f
C75 VDD1.t3 VSUBS 0.034363f
C76 VDD1.n2 VSUBS 0.177772f
C77 VDD1.n3 VSUBS 1.16472f
C78 VTAIL.t0 VSUBS 0.0689f
C79 VTAIL.t2 VSUBS 0.0689f
C80 VTAIL.n0 VSUBS 0.306621f
C81 VTAIL.n1 VSUBS 0.56617f
C82 VTAIL.t8 VSUBS 0.45911f
C83 VTAIL.n2 VSUBS 0.726039f
C84 VTAIL.t11 VSUBS 0.0689f
C85 VTAIL.t6 VSUBS 0.0689f
C86 VTAIL.n3 VSUBS 0.306621f
C87 VTAIL.n4 VSUBS 1.55717f
C88 VTAIL.t3 VSUBS 0.0689f
C89 VTAIL.t5 VSUBS 0.0689f
C90 VTAIL.n5 VSUBS 0.306622f
C91 VTAIL.n6 VSUBS 1.55717f
C92 VTAIL.t1 VSUBS 0.459112f
C93 VTAIL.n7 VSUBS 0.726037f
C94 VTAIL.t7 VSUBS 0.0689f
C95 VTAIL.t9 VSUBS 0.0689f
C96 VTAIL.n8 VSUBS 0.306622f
C97 VTAIL.n9 VSUBS 0.690618f
C98 VTAIL.t10 VSUBS 0.45911f
C99 VTAIL.n10 VSUBS 1.41911f
C100 VTAIL.t4 VSUBS 0.45911f
C101 VTAIL.n11 VSUBS 1.37009f
C102 VP.n0 VSUBS 0.04929f
C103 VP.t0 VSUBS 0.614507f
C104 VP.n1 VSUBS 0.04063f
C105 VP.n2 VSUBS 0.04929f
C106 VP.t4 VSUBS 0.614507f
C107 VP.n3 VSUBS 0.04063f
C108 VP.n4 VSUBS 0.04929f
C109 VP.t3 VSUBS 0.614507f
C110 VP.n5 VSUBS 0.04929f
C111 VP.t2 VSUBS 0.614507f
C112 VP.n6 VSUBS 0.04063f
C113 VP.t5 VSUBS 0.84775f
C114 VP.n7 VSUBS 0.363653f
C115 VP.t1 VSUBS 0.614507f
C116 VP.n8 VSUBS 0.408179f
C117 VP.n9 VSUBS 0.099275f
C118 VP.n10 VSUBS 0.360439f
C119 VP.n11 VSUBS 0.04929f
C120 VP.n12 VSUBS 0.04929f
C121 VP.n13 VSUBS 0.09588f
C122 VP.n14 VSUBS 0.05286f
C123 VP.n15 VSUBS 0.383035f
C124 VP.n16 VSUBS 1.74827f
C125 VP.n17 VSUBS 1.79455f
C126 VP.n18 VSUBS 0.383035f
C127 VP.n19 VSUBS 0.05286f
C128 VP.n20 VSUBS 0.09588f
C129 VP.n21 VSUBS 0.04929f
C130 VP.n22 VSUBS 0.04929f
C131 VP.n23 VSUBS 0.04929f
C132 VP.n24 VSUBS 0.099275f
C133 VP.n25 VSUBS 0.323407f
C134 VP.n26 VSUBS 0.099275f
C135 VP.n27 VSUBS 0.04929f
C136 VP.n28 VSUBS 0.04929f
C137 VP.n29 VSUBS 0.04929f
C138 VP.n30 VSUBS 0.09588f
C139 VP.n31 VSUBS 0.05286f
C140 VP.n32 VSUBS 0.383035f
C141 VP.n33 VSUBS 0.052044f
C142 B.n0 VSUBS 0.006932f
C143 B.n1 VSUBS 0.006932f
C144 B.n2 VSUBS 0.010253f
C145 B.n3 VSUBS 0.007857f
C146 B.n4 VSUBS 0.007857f
C147 B.n5 VSUBS 0.007857f
C148 B.n6 VSUBS 0.007857f
C149 B.n7 VSUBS 0.007857f
C150 B.n8 VSUBS 0.007857f
C151 B.n9 VSUBS 0.007857f
C152 B.n10 VSUBS 0.007857f
C153 B.n11 VSUBS 0.007857f
C154 B.n12 VSUBS 0.007857f
C155 B.n13 VSUBS 0.007857f
C156 B.n14 VSUBS 0.007857f
C157 B.n15 VSUBS 0.007857f
C158 B.n16 VSUBS 0.007857f
C159 B.n17 VSUBS 0.007857f
C160 B.n18 VSUBS 0.018925f
C161 B.n19 VSUBS 0.007857f
C162 B.n20 VSUBS 0.007857f
C163 B.n21 VSUBS 0.007857f
C164 B.n22 VSUBS 0.007857f
C165 B.n23 VSUBS 0.007857f
C166 B.n24 VSUBS 0.007857f
C167 B.n25 VSUBS 0.007857f
C168 B.t10 VSUBS 0.077234f
C169 B.t11 VSUBS 0.089779f
C170 B.t9 VSUBS 0.271363f
C171 B.n26 VSUBS 0.082288f
C172 B.n27 VSUBS 0.068593f
C173 B.n28 VSUBS 0.007857f
C174 B.n29 VSUBS 0.007857f
C175 B.n30 VSUBS 0.007857f
C176 B.n31 VSUBS 0.007857f
C177 B.t4 VSUBS 0.077234f
C178 B.t5 VSUBS 0.089779f
C179 B.t3 VSUBS 0.271363f
C180 B.n32 VSUBS 0.082288f
C181 B.n33 VSUBS 0.068593f
C182 B.n34 VSUBS 0.018203f
C183 B.n35 VSUBS 0.007857f
C184 B.n36 VSUBS 0.007857f
C185 B.n37 VSUBS 0.007857f
C186 B.n38 VSUBS 0.007857f
C187 B.n39 VSUBS 0.007857f
C188 B.n40 VSUBS 0.007857f
C189 B.n41 VSUBS 0.007857f
C190 B.n42 VSUBS 0.01828f
C191 B.n43 VSUBS 0.007857f
C192 B.n44 VSUBS 0.007857f
C193 B.n45 VSUBS 0.007857f
C194 B.n46 VSUBS 0.007857f
C195 B.n47 VSUBS 0.007857f
C196 B.n48 VSUBS 0.007857f
C197 B.n49 VSUBS 0.007857f
C198 B.n50 VSUBS 0.007857f
C199 B.n51 VSUBS 0.007857f
C200 B.n52 VSUBS 0.007857f
C201 B.n53 VSUBS 0.007857f
C202 B.n54 VSUBS 0.007857f
C203 B.n55 VSUBS 0.007857f
C204 B.n56 VSUBS 0.007857f
C205 B.n57 VSUBS 0.007857f
C206 B.n58 VSUBS 0.007857f
C207 B.n59 VSUBS 0.007857f
C208 B.n60 VSUBS 0.007857f
C209 B.n61 VSUBS 0.007857f
C210 B.n62 VSUBS 0.007857f
C211 B.n63 VSUBS 0.007857f
C212 B.n64 VSUBS 0.007857f
C213 B.n65 VSUBS 0.007857f
C214 B.n66 VSUBS 0.007857f
C215 B.n67 VSUBS 0.007857f
C216 B.n68 VSUBS 0.007857f
C217 B.n69 VSUBS 0.007857f
C218 B.n70 VSUBS 0.007857f
C219 B.n71 VSUBS 0.007857f
C220 B.n72 VSUBS 0.007857f
C221 B.n73 VSUBS 0.007857f
C222 B.n74 VSUBS 0.007857f
C223 B.n75 VSUBS 0.018925f
C224 B.n76 VSUBS 0.007857f
C225 B.n77 VSUBS 0.007857f
C226 B.n78 VSUBS 0.007857f
C227 B.n79 VSUBS 0.007857f
C228 B.n80 VSUBS 0.007857f
C229 B.n81 VSUBS 0.007857f
C230 B.n82 VSUBS 0.00543f
C231 B.n83 VSUBS 0.007857f
C232 B.n84 VSUBS 0.007857f
C233 B.n85 VSUBS 0.007857f
C234 B.n86 VSUBS 0.007857f
C235 B.n87 VSUBS 0.007857f
C236 B.t8 VSUBS 0.077234f
C237 B.t7 VSUBS 0.089779f
C238 B.t6 VSUBS 0.271363f
C239 B.n88 VSUBS 0.082288f
C240 B.n89 VSUBS 0.068593f
C241 B.n90 VSUBS 0.007857f
C242 B.n91 VSUBS 0.007857f
C243 B.n92 VSUBS 0.007857f
C244 B.n93 VSUBS 0.007857f
C245 B.n94 VSUBS 0.007857f
C246 B.n95 VSUBS 0.007857f
C247 B.n96 VSUBS 0.018925f
C248 B.n97 VSUBS 0.007857f
C249 B.n98 VSUBS 0.007857f
C250 B.n99 VSUBS 0.007857f
C251 B.n100 VSUBS 0.007857f
C252 B.n101 VSUBS 0.007857f
C253 B.n102 VSUBS 0.007857f
C254 B.n103 VSUBS 0.007857f
C255 B.n104 VSUBS 0.007857f
C256 B.n105 VSUBS 0.007857f
C257 B.n106 VSUBS 0.007857f
C258 B.n107 VSUBS 0.007857f
C259 B.n108 VSUBS 0.007857f
C260 B.n109 VSUBS 0.007857f
C261 B.n110 VSUBS 0.007857f
C262 B.n111 VSUBS 0.007857f
C263 B.n112 VSUBS 0.007857f
C264 B.n113 VSUBS 0.007857f
C265 B.n114 VSUBS 0.007857f
C266 B.n115 VSUBS 0.007857f
C267 B.n116 VSUBS 0.007857f
C268 B.n117 VSUBS 0.007857f
C269 B.n118 VSUBS 0.007857f
C270 B.n119 VSUBS 0.007857f
C271 B.n120 VSUBS 0.007857f
C272 B.n121 VSUBS 0.007857f
C273 B.n122 VSUBS 0.007857f
C274 B.n123 VSUBS 0.007857f
C275 B.n124 VSUBS 0.007857f
C276 B.n125 VSUBS 0.007857f
C277 B.n126 VSUBS 0.007857f
C278 B.n127 VSUBS 0.007857f
C279 B.n128 VSUBS 0.007857f
C280 B.n129 VSUBS 0.007857f
C281 B.n130 VSUBS 0.007857f
C282 B.n131 VSUBS 0.007857f
C283 B.n132 VSUBS 0.007857f
C284 B.n133 VSUBS 0.007857f
C285 B.n134 VSUBS 0.007857f
C286 B.n135 VSUBS 0.007857f
C287 B.n136 VSUBS 0.007857f
C288 B.n137 VSUBS 0.007857f
C289 B.n138 VSUBS 0.007857f
C290 B.n139 VSUBS 0.007857f
C291 B.n140 VSUBS 0.007857f
C292 B.n141 VSUBS 0.007857f
C293 B.n142 VSUBS 0.007857f
C294 B.n143 VSUBS 0.007857f
C295 B.n144 VSUBS 0.007857f
C296 B.n145 VSUBS 0.007857f
C297 B.n146 VSUBS 0.007857f
C298 B.n147 VSUBS 0.007857f
C299 B.n148 VSUBS 0.007857f
C300 B.n149 VSUBS 0.007857f
C301 B.n150 VSUBS 0.007857f
C302 B.n151 VSUBS 0.007857f
C303 B.n152 VSUBS 0.007857f
C304 B.n153 VSUBS 0.007857f
C305 B.n154 VSUBS 0.007857f
C306 B.n155 VSUBS 0.007857f
C307 B.n156 VSUBS 0.007857f
C308 B.n157 VSUBS 0.01828f
C309 B.n158 VSUBS 0.01828f
C310 B.n159 VSUBS 0.018925f
C311 B.n160 VSUBS 0.007857f
C312 B.n161 VSUBS 0.007857f
C313 B.n162 VSUBS 0.007857f
C314 B.n163 VSUBS 0.007857f
C315 B.n164 VSUBS 0.007857f
C316 B.n165 VSUBS 0.007857f
C317 B.n166 VSUBS 0.007857f
C318 B.n167 VSUBS 0.007857f
C319 B.n168 VSUBS 0.007857f
C320 B.n169 VSUBS 0.007857f
C321 B.n170 VSUBS 0.007857f
C322 B.n171 VSUBS 0.007857f
C323 B.n172 VSUBS 0.007857f
C324 B.n173 VSUBS 0.007857f
C325 B.n174 VSUBS 0.007857f
C326 B.n175 VSUBS 0.007857f
C327 B.n176 VSUBS 0.007857f
C328 B.n177 VSUBS 0.007857f
C329 B.n178 VSUBS 0.007857f
C330 B.n179 VSUBS 0.007857f
C331 B.n180 VSUBS 0.00543f
C332 B.n181 VSUBS 0.018203f
C333 B.n182 VSUBS 0.006355f
C334 B.n183 VSUBS 0.007857f
C335 B.n184 VSUBS 0.007857f
C336 B.n185 VSUBS 0.007857f
C337 B.n186 VSUBS 0.007857f
C338 B.n187 VSUBS 0.007857f
C339 B.n188 VSUBS 0.007857f
C340 B.n189 VSUBS 0.007857f
C341 B.n190 VSUBS 0.007857f
C342 B.n191 VSUBS 0.007857f
C343 B.n192 VSUBS 0.007857f
C344 B.n193 VSUBS 0.007857f
C345 B.t2 VSUBS 0.077234f
C346 B.t1 VSUBS 0.089779f
C347 B.t0 VSUBS 0.271363f
C348 B.n194 VSUBS 0.082288f
C349 B.n195 VSUBS 0.068593f
C350 B.n196 VSUBS 0.018203f
C351 B.n197 VSUBS 0.006355f
C352 B.n198 VSUBS 0.007857f
C353 B.n199 VSUBS 0.007857f
C354 B.n200 VSUBS 0.007857f
C355 B.n201 VSUBS 0.007857f
C356 B.n202 VSUBS 0.007857f
C357 B.n203 VSUBS 0.007857f
C358 B.n204 VSUBS 0.007857f
C359 B.n205 VSUBS 0.007857f
C360 B.n206 VSUBS 0.007857f
C361 B.n207 VSUBS 0.007857f
C362 B.n208 VSUBS 0.007857f
C363 B.n209 VSUBS 0.007857f
C364 B.n210 VSUBS 0.007857f
C365 B.n211 VSUBS 0.007857f
C366 B.n212 VSUBS 0.007857f
C367 B.n213 VSUBS 0.007857f
C368 B.n214 VSUBS 0.007857f
C369 B.n215 VSUBS 0.007857f
C370 B.n216 VSUBS 0.007857f
C371 B.n217 VSUBS 0.007857f
C372 B.n218 VSUBS 0.007857f
C373 B.n219 VSUBS 0.007857f
C374 B.n220 VSUBS 0.018013f
C375 B.n221 VSUBS 0.019191f
C376 B.n222 VSUBS 0.01828f
C377 B.n223 VSUBS 0.007857f
C378 B.n224 VSUBS 0.007857f
C379 B.n225 VSUBS 0.007857f
C380 B.n226 VSUBS 0.007857f
C381 B.n227 VSUBS 0.007857f
C382 B.n228 VSUBS 0.007857f
C383 B.n229 VSUBS 0.007857f
C384 B.n230 VSUBS 0.007857f
C385 B.n231 VSUBS 0.007857f
C386 B.n232 VSUBS 0.007857f
C387 B.n233 VSUBS 0.007857f
C388 B.n234 VSUBS 0.007857f
C389 B.n235 VSUBS 0.007857f
C390 B.n236 VSUBS 0.007857f
C391 B.n237 VSUBS 0.007857f
C392 B.n238 VSUBS 0.007857f
C393 B.n239 VSUBS 0.007857f
C394 B.n240 VSUBS 0.007857f
C395 B.n241 VSUBS 0.007857f
C396 B.n242 VSUBS 0.007857f
C397 B.n243 VSUBS 0.007857f
C398 B.n244 VSUBS 0.007857f
C399 B.n245 VSUBS 0.007857f
C400 B.n246 VSUBS 0.007857f
C401 B.n247 VSUBS 0.007857f
C402 B.n248 VSUBS 0.007857f
C403 B.n249 VSUBS 0.007857f
C404 B.n250 VSUBS 0.007857f
C405 B.n251 VSUBS 0.007857f
C406 B.n252 VSUBS 0.007857f
C407 B.n253 VSUBS 0.007857f
C408 B.n254 VSUBS 0.007857f
C409 B.n255 VSUBS 0.007857f
C410 B.n256 VSUBS 0.007857f
C411 B.n257 VSUBS 0.007857f
C412 B.n258 VSUBS 0.007857f
C413 B.n259 VSUBS 0.007857f
C414 B.n260 VSUBS 0.007857f
C415 B.n261 VSUBS 0.007857f
C416 B.n262 VSUBS 0.007857f
C417 B.n263 VSUBS 0.007857f
C418 B.n264 VSUBS 0.007857f
C419 B.n265 VSUBS 0.007857f
C420 B.n266 VSUBS 0.007857f
C421 B.n267 VSUBS 0.007857f
C422 B.n268 VSUBS 0.007857f
C423 B.n269 VSUBS 0.007857f
C424 B.n270 VSUBS 0.007857f
C425 B.n271 VSUBS 0.007857f
C426 B.n272 VSUBS 0.007857f
C427 B.n273 VSUBS 0.007857f
C428 B.n274 VSUBS 0.007857f
C429 B.n275 VSUBS 0.007857f
C430 B.n276 VSUBS 0.007857f
C431 B.n277 VSUBS 0.007857f
C432 B.n278 VSUBS 0.007857f
C433 B.n279 VSUBS 0.007857f
C434 B.n280 VSUBS 0.007857f
C435 B.n281 VSUBS 0.007857f
C436 B.n282 VSUBS 0.007857f
C437 B.n283 VSUBS 0.007857f
C438 B.n284 VSUBS 0.007857f
C439 B.n285 VSUBS 0.007857f
C440 B.n286 VSUBS 0.007857f
C441 B.n287 VSUBS 0.007857f
C442 B.n288 VSUBS 0.007857f
C443 B.n289 VSUBS 0.007857f
C444 B.n290 VSUBS 0.007857f
C445 B.n291 VSUBS 0.007857f
C446 B.n292 VSUBS 0.007857f
C447 B.n293 VSUBS 0.007857f
C448 B.n294 VSUBS 0.007857f
C449 B.n295 VSUBS 0.007857f
C450 B.n296 VSUBS 0.007857f
C451 B.n297 VSUBS 0.007857f
C452 B.n298 VSUBS 0.007857f
C453 B.n299 VSUBS 0.007857f
C454 B.n300 VSUBS 0.007857f
C455 B.n301 VSUBS 0.007857f
C456 B.n302 VSUBS 0.007857f
C457 B.n303 VSUBS 0.007857f
C458 B.n304 VSUBS 0.007857f
C459 B.n305 VSUBS 0.007857f
C460 B.n306 VSUBS 0.007857f
C461 B.n307 VSUBS 0.007857f
C462 B.n308 VSUBS 0.007857f
C463 B.n309 VSUBS 0.007857f
C464 B.n310 VSUBS 0.007857f
C465 B.n311 VSUBS 0.007857f
C466 B.n312 VSUBS 0.007857f
C467 B.n313 VSUBS 0.007857f
C468 B.n314 VSUBS 0.007857f
C469 B.n315 VSUBS 0.007857f
C470 B.n316 VSUBS 0.007857f
C471 B.n317 VSUBS 0.007857f
C472 B.n318 VSUBS 0.007857f
C473 B.n319 VSUBS 0.01828f
C474 B.n320 VSUBS 0.018925f
C475 B.n321 VSUBS 0.018925f
C476 B.n322 VSUBS 0.007857f
C477 B.n323 VSUBS 0.007857f
C478 B.n324 VSUBS 0.007857f
C479 B.n325 VSUBS 0.007857f
C480 B.n326 VSUBS 0.007857f
C481 B.n327 VSUBS 0.007857f
C482 B.n328 VSUBS 0.007857f
C483 B.n329 VSUBS 0.007857f
C484 B.n330 VSUBS 0.007857f
C485 B.n331 VSUBS 0.007857f
C486 B.n332 VSUBS 0.007857f
C487 B.n333 VSUBS 0.007857f
C488 B.n334 VSUBS 0.007857f
C489 B.n335 VSUBS 0.007857f
C490 B.n336 VSUBS 0.007857f
C491 B.n337 VSUBS 0.007857f
C492 B.n338 VSUBS 0.007857f
C493 B.n339 VSUBS 0.007857f
C494 B.n340 VSUBS 0.007857f
C495 B.n341 VSUBS 0.00543f
C496 B.n342 VSUBS 0.007857f
C497 B.n343 VSUBS 0.007857f
C498 B.n344 VSUBS 0.006355f
C499 B.n345 VSUBS 0.007857f
C500 B.n346 VSUBS 0.007857f
C501 B.n347 VSUBS 0.007857f
C502 B.n348 VSUBS 0.007857f
C503 B.n349 VSUBS 0.007857f
C504 B.n350 VSUBS 0.007857f
C505 B.n351 VSUBS 0.007857f
C506 B.n352 VSUBS 0.007857f
C507 B.n353 VSUBS 0.007857f
C508 B.n354 VSUBS 0.007857f
C509 B.n355 VSUBS 0.007857f
C510 B.n356 VSUBS 0.006355f
C511 B.n357 VSUBS 0.018203f
C512 B.n358 VSUBS 0.00543f
C513 B.n359 VSUBS 0.007857f
C514 B.n360 VSUBS 0.007857f
C515 B.n361 VSUBS 0.007857f
C516 B.n362 VSUBS 0.007857f
C517 B.n363 VSUBS 0.007857f
C518 B.n364 VSUBS 0.007857f
C519 B.n365 VSUBS 0.007857f
C520 B.n366 VSUBS 0.007857f
C521 B.n367 VSUBS 0.007857f
C522 B.n368 VSUBS 0.007857f
C523 B.n369 VSUBS 0.007857f
C524 B.n370 VSUBS 0.007857f
C525 B.n371 VSUBS 0.007857f
C526 B.n372 VSUBS 0.007857f
C527 B.n373 VSUBS 0.007857f
C528 B.n374 VSUBS 0.007857f
C529 B.n375 VSUBS 0.007857f
C530 B.n376 VSUBS 0.007857f
C531 B.n377 VSUBS 0.007857f
C532 B.n378 VSUBS 0.007857f
C533 B.n379 VSUBS 0.018925f
C534 B.n380 VSUBS 0.01828f
C535 B.n381 VSUBS 0.01828f
C536 B.n382 VSUBS 0.007857f
C537 B.n383 VSUBS 0.007857f
C538 B.n384 VSUBS 0.007857f
C539 B.n385 VSUBS 0.007857f
C540 B.n386 VSUBS 0.007857f
C541 B.n387 VSUBS 0.007857f
C542 B.n388 VSUBS 0.007857f
C543 B.n389 VSUBS 0.007857f
C544 B.n390 VSUBS 0.007857f
C545 B.n391 VSUBS 0.007857f
C546 B.n392 VSUBS 0.007857f
C547 B.n393 VSUBS 0.007857f
C548 B.n394 VSUBS 0.007857f
C549 B.n395 VSUBS 0.007857f
C550 B.n396 VSUBS 0.007857f
C551 B.n397 VSUBS 0.007857f
C552 B.n398 VSUBS 0.007857f
C553 B.n399 VSUBS 0.007857f
C554 B.n400 VSUBS 0.007857f
C555 B.n401 VSUBS 0.007857f
C556 B.n402 VSUBS 0.007857f
C557 B.n403 VSUBS 0.007857f
C558 B.n404 VSUBS 0.007857f
C559 B.n405 VSUBS 0.007857f
C560 B.n406 VSUBS 0.007857f
C561 B.n407 VSUBS 0.007857f
C562 B.n408 VSUBS 0.007857f
C563 B.n409 VSUBS 0.007857f
C564 B.n410 VSUBS 0.007857f
C565 B.n411 VSUBS 0.007857f
C566 B.n412 VSUBS 0.007857f
C567 B.n413 VSUBS 0.007857f
C568 B.n414 VSUBS 0.007857f
C569 B.n415 VSUBS 0.007857f
C570 B.n416 VSUBS 0.007857f
C571 B.n417 VSUBS 0.007857f
C572 B.n418 VSUBS 0.007857f
C573 B.n419 VSUBS 0.007857f
C574 B.n420 VSUBS 0.007857f
C575 B.n421 VSUBS 0.007857f
C576 B.n422 VSUBS 0.007857f
C577 B.n423 VSUBS 0.007857f
C578 B.n424 VSUBS 0.007857f
C579 B.n425 VSUBS 0.007857f
C580 B.n426 VSUBS 0.007857f
C581 B.n427 VSUBS 0.010253f
C582 B.n428 VSUBS 0.010922f
C583 B.n429 VSUBS 0.021719f
.ends

