* NGSPICE file created from diff_pair_sample_0505.ext - technology: sky130A

.subckt diff_pair_sample_0505 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=0.66825 pd=4.38 as=1.5795 ps=8.88 w=4.05 l=3.93
X1 VDD1.t2 VP.t1 VTAIL.t5 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=0.66825 pd=4.38 as=1.5795 ps=8.88 w=4.05 l=3.93
X2 VTAIL.t2 VN.t0 VDD2.t3 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0.66825 ps=4.38 w=4.05 l=3.93
X3 VTAIL.t3 VN.t1 VDD2.t2 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0.66825 ps=4.38 w=4.05 l=3.93
X4 B.t11 B.t9 B.t10 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0 ps=0 w=4.05 l=3.93
X5 B.t8 B.t6 B.t7 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0 ps=0 w=4.05 l=3.93
X6 VDD2.t1 VN.t2 VTAIL.t1 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=0.66825 pd=4.38 as=1.5795 ps=8.88 w=4.05 l=3.93
X7 B.t5 B.t3 B.t4 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0 ps=0 w=4.05 l=3.93
X8 VTAIL.t6 VP.t2 VDD1.t1 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0.66825 ps=4.38 w=4.05 l=3.93
X9 VTAIL.t7 VP.t3 VDD1.t0 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0.66825 ps=4.38 w=4.05 l=3.93
X10 VDD2.t0 VN.t3 VTAIL.t0 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=0.66825 pd=4.38 as=1.5795 ps=8.88 w=4.05 l=3.93
X11 B.t2 B.t0 B.t1 w_n3526_n1778# sky130_fd_pr__pfet_01v8 ad=1.5795 pd=8.88 as=0 ps=0 w=4.05 l=3.93
R0 VP.n18 VP.n0 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n15 VP.n1 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n12 VP.n2 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n3 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n6 VP.n5 63.5869
R9 VP.n20 VP.n19 63.5869
R10 VP.n4 VP.t3 58.6619
R11 VP.n4 VP.t1 57.235
R12 VP.n13 VP.n12 56.5193
R13 VP.n5 VP.n4 46.237
R14 VP.n6 VP.t2 24.8364
R15 VP.n19 VP.t0 24.8364
R16 VP.n7 VP.n3 24.4675
R17 VP.n11 VP.n3 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n13 VP.n1 24.4675
R20 VP.n17 VP.n1 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n7 VP.n6 18.5954
R23 VP.n19 VP.n18 18.5954
R24 VP.n8 VP.n5 0.417535
R25 VP.n20 VP.n0 0.417535
R26 VP VP.n20 0.394291
R27 VP.n9 VP.n8 0.189894
R28 VP.n10 VP.n9 0.189894
R29 VP.n10 VP.n2 0.189894
R30 VP.n14 VP.n2 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VTAIL.n154 VTAIL.n140 756.745
R35 VTAIL.n14 VTAIL.n0 756.745
R36 VTAIL.n34 VTAIL.n20 756.745
R37 VTAIL.n54 VTAIL.n40 756.745
R38 VTAIL.n134 VTAIL.n120 756.745
R39 VTAIL.n114 VTAIL.n100 756.745
R40 VTAIL.n94 VTAIL.n80 756.745
R41 VTAIL.n74 VTAIL.n60 756.745
R42 VTAIL.n147 VTAIL.n146 585
R43 VTAIL.n144 VTAIL.n143 585
R44 VTAIL.n153 VTAIL.n152 585
R45 VTAIL.n155 VTAIL.n154 585
R46 VTAIL.n7 VTAIL.n6 585
R47 VTAIL.n4 VTAIL.n3 585
R48 VTAIL.n13 VTAIL.n12 585
R49 VTAIL.n15 VTAIL.n14 585
R50 VTAIL.n27 VTAIL.n26 585
R51 VTAIL.n24 VTAIL.n23 585
R52 VTAIL.n33 VTAIL.n32 585
R53 VTAIL.n35 VTAIL.n34 585
R54 VTAIL.n47 VTAIL.n46 585
R55 VTAIL.n44 VTAIL.n43 585
R56 VTAIL.n53 VTAIL.n52 585
R57 VTAIL.n55 VTAIL.n54 585
R58 VTAIL.n135 VTAIL.n134 585
R59 VTAIL.n133 VTAIL.n132 585
R60 VTAIL.n124 VTAIL.n123 585
R61 VTAIL.n127 VTAIL.n126 585
R62 VTAIL.n115 VTAIL.n114 585
R63 VTAIL.n113 VTAIL.n112 585
R64 VTAIL.n104 VTAIL.n103 585
R65 VTAIL.n107 VTAIL.n106 585
R66 VTAIL.n95 VTAIL.n94 585
R67 VTAIL.n93 VTAIL.n92 585
R68 VTAIL.n84 VTAIL.n83 585
R69 VTAIL.n87 VTAIL.n86 585
R70 VTAIL.n75 VTAIL.n74 585
R71 VTAIL.n73 VTAIL.n72 585
R72 VTAIL.n64 VTAIL.n63 585
R73 VTAIL.n67 VTAIL.n66 585
R74 VTAIL.t0 VTAIL.n145 330.707
R75 VTAIL.t3 VTAIL.n5 330.707
R76 VTAIL.t4 VTAIL.n25 330.707
R77 VTAIL.t6 VTAIL.n45 330.707
R78 VTAIL.t5 VTAIL.n125 330.707
R79 VTAIL.t7 VTAIL.n105 330.707
R80 VTAIL.t1 VTAIL.n85 330.707
R81 VTAIL.t2 VTAIL.n65 330.707
R82 VTAIL.n146 VTAIL.n143 171.744
R83 VTAIL.n153 VTAIL.n143 171.744
R84 VTAIL.n154 VTAIL.n153 171.744
R85 VTAIL.n6 VTAIL.n3 171.744
R86 VTAIL.n13 VTAIL.n3 171.744
R87 VTAIL.n14 VTAIL.n13 171.744
R88 VTAIL.n26 VTAIL.n23 171.744
R89 VTAIL.n33 VTAIL.n23 171.744
R90 VTAIL.n34 VTAIL.n33 171.744
R91 VTAIL.n46 VTAIL.n43 171.744
R92 VTAIL.n53 VTAIL.n43 171.744
R93 VTAIL.n54 VTAIL.n53 171.744
R94 VTAIL.n134 VTAIL.n133 171.744
R95 VTAIL.n133 VTAIL.n123 171.744
R96 VTAIL.n126 VTAIL.n123 171.744
R97 VTAIL.n114 VTAIL.n113 171.744
R98 VTAIL.n113 VTAIL.n103 171.744
R99 VTAIL.n106 VTAIL.n103 171.744
R100 VTAIL.n94 VTAIL.n93 171.744
R101 VTAIL.n93 VTAIL.n83 171.744
R102 VTAIL.n86 VTAIL.n83 171.744
R103 VTAIL.n74 VTAIL.n73 171.744
R104 VTAIL.n73 VTAIL.n63 171.744
R105 VTAIL.n66 VTAIL.n63 171.744
R106 VTAIL.n146 VTAIL.t0 85.8723
R107 VTAIL.n6 VTAIL.t3 85.8723
R108 VTAIL.n26 VTAIL.t4 85.8723
R109 VTAIL.n46 VTAIL.t6 85.8723
R110 VTAIL.n126 VTAIL.t5 85.8723
R111 VTAIL.n106 VTAIL.t7 85.8723
R112 VTAIL.n86 VTAIL.t1 85.8723
R113 VTAIL.n66 VTAIL.t2 85.8723
R114 VTAIL.n159 VTAIL.n158 36.2581
R115 VTAIL.n19 VTAIL.n18 36.2581
R116 VTAIL.n39 VTAIL.n38 36.2581
R117 VTAIL.n59 VTAIL.n58 36.2581
R118 VTAIL.n139 VTAIL.n138 36.2581
R119 VTAIL.n119 VTAIL.n118 36.2581
R120 VTAIL.n99 VTAIL.n98 36.2581
R121 VTAIL.n79 VTAIL.n78 36.2581
R122 VTAIL.n159 VTAIL.n139 19.5307
R123 VTAIL.n79 VTAIL.n59 19.5307
R124 VTAIL.n147 VTAIL.n145 16.3201
R125 VTAIL.n7 VTAIL.n5 16.3201
R126 VTAIL.n27 VTAIL.n25 16.3201
R127 VTAIL.n47 VTAIL.n45 16.3201
R128 VTAIL.n127 VTAIL.n125 16.3201
R129 VTAIL.n107 VTAIL.n105 16.3201
R130 VTAIL.n87 VTAIL.n85 16.3201
R131 VTAIL.n67 VTAIL.n65 16.3201
R132 VTAIL.n148 VTAIL.n144 12.8005
R133 VTAIL.n8 VTAIL.n4 12.8005
R134 VTAIL.n28 VTAIL.n24 12.8005
R135 VTAIL.n48 VTAIL.n44 12.8005
R136 VTAIL.n128 VTAIL.n124 12.8005
R137 VTAIL.n108 VTAIL.n104 12.8005
R138 VTAIL.n88 VTAIL.n84 12.8005
R139 VTAIL.n68 VTAIL.n64 12.8005
R140 VTAIL.n152 VTAIL.n151 12.0247
R141 VTAIL.n12 VTAIL.n11 12.0247
R142 VTAIL.n32 VTAIL.n31 12.0247
R143 VTAIL.n52 VTAIL.n51 12.0247
R144 VTAIL.n132 VTAIL.n131 12.0247
R145 VTAIL.n112 VTAIL.n111 12.0247
R146 VTAIL.n92 VTAIL.n91 12.0247
R147 VTAIL.n72 VTAIL.n71 12.0247
R148 VTAIL.n155 VTAIL.n142 11.249
R149 VTAIL.n15 VTAIL.n2 11.249
R150 VTAIL.n35 VTAIL.n22 11.249
R151 VTAIL.n55 VTAIL.n42 11.249
R152 VTAIL.n135 VTAIL.n122 11.249
R153 VTAIL.n115 VTAIL.n102 11.249
R154 VTAIL.n95 VTAIL.n82 11.249
R155 VTAIL.n75 VTAIL.n62 11.249
R156 VTAIL.n156 VTAIL.n140 10.4732
R157 VTAIL.n16 VTAIL.n0 10.4732
R158 VTAIL.n36 VTAIL.n20 10.4732
R159 VTAIL.n56 VTAIL.n40 10.4732
R160 VTAIL.n136 VTAIL.n120 10.4732
R161 VTAIL.n116 VTAIL.n100 10.4732
R162 VTAIL.n96 VTAIL.n80 10.4732
R163 VTAIL.n76 VTAIL.n60 10.4732
R164 VTAIL.n158 VTAIL.n157 9.45567
R165 VTAIL.n18 VTAIL.n17 9.45567
R166 VTAIL.n38 VTAIL.n37 9.45567
R167 VTAIL.n58 VTAIL.n57 9.45567
R168 VTAIL.n138 VTAIL.n137 9.45567
R169 VTAIL.n118 VTAIL.n117 9.45567
R170 VTAIL.n98 VTAIL.n97 9.45567
R171 VTAIL.n78 VTAIL.n77 9.45567
R172 VTAIL.n157 VTAIL.n156 9.3005
R173 VTAIL.n142 VTAIL.n141 9.3005
R174 VTAIL.n151 VTAIL.n150 9.3005
R175 VTAIL.n149 VTAIL.n148 9.3005
R176 VTAIL.n17 VTAIL.n16 9.3005
R177 VTAIL.n2 VTAIL.n1 9.3005
R178 VTAIL.n11 VTAIL.n10 9.3005
R179 VTAIL.n9 VTAIL.n8 9.3005
R180 VTAIL.n37 VTAIL.n36 9.3005
R181 VTAIL.n22 VTAIL.n21 9.3005
R182 VTAIL.n31 VTAIL.n30 9.3005
R183 VTAIL.n29 VTAIL.n28 9.3005
R184 VTAIL.n57 VTAIL.n56 9.3005
R185 VTAIL.n42 VTAIL.n41 9.3005
R186 VTAIL.n51 VTAIL.n50 9.3005
R187 VTAIL.n49 VTAIL.n48 9.3005
R188 VTAIL.n137 VTAIL.n136 9.3005
R189 VTAIL.n122 VTAIL.n121 9.3005
R190 VTAIL.n131 VTAIL.n130 9.3005
R191 VTAIL.n129 VTAIL.n128 9.3005
R192 VTAIL.n117 VTAIL.n116 9.3005
R193 VTAIL.n102 VTAIL.n101 9.3005
R194 VTAIL.n111 VTAIL.n110 9.3005
R195 VTAIL.n109 VTAIL.n108 9.3005
R196 VTAIL.n97 VTAIL.n96 9.3005
R197 VTAIL.n82 VTAIL.n81 9.3005
R198 VTAIL.n91 VTAIL.n90 9.3005
R199 VTAIL.n89 VTAIL.n88 9.3005
R200 VTAIL.n77 VTAIL.n76 9.3005
R201 VTAIL.n62 VTAIL.n61 9.3005
R202 VTAIL.n71 VTAIL.n70 9.3005
R203 VTAIL.n69 VTAIL.n68 9.3005
R204 VTAIL.n149 VTAIL.n145 3.78097
R205 VTAIL.n9 VTAIL.n5 3.78097
R206 VTAIL.n29 VTAIL.n25 3.78097
R207 VTAIL.n49 VTAIL.n45 3.78097
R208 VTAIL.n129 VTAIL.n125 3.78097
R209 VTAIL.n109 VTAIL.n105 3.78097
R210 VTAIL.n89 VTAIL.n85 3.78097
R211 VTAIL.n69 VTAIL.n65 3.78097
R212 VTAIL.n99 VTAIL.n79 3.67291
R213 VTAIL.n139 VTAIL.n119 3.67291
R214 VTAIL.n59 VTAIL.n39 3.67291
R215 VTAIL.n158 VTAIL.n140 3.49141
R216 VTAIL.n18 VTAIL.n0 3.49141
R217 VTAIL.n38 VTAIL.n20 3.49141
R218 VTAIL.n58 VTAIL.n40 3.49141
R219 VTAIL.n138 VTAIL.n120 3.49141
R220 VTAIL.n118 VTAIL.n100 3.49141
R221 VTAIL.n98 VTAIL.n80 3.49141
R222 VTAIL.n78 VTAIL.n60 3.49141
R223 VTAIL.n156 VTAIL.n155 2.71565
R224 VTAIL.n16 VTAIL.n15 2.71565
R225 VTAIL.n36 VTAIL.n35 2.71565
R226 VTAIL.n56 VTAIL.n55 2.71565
R227 VTAIL.n136 VTAIL.n135 2.71565
R228 VTAIL.n116 VTAIL.n115 2.71565
R229 VTAIL.n96 VTAIL.n95 2.71565
R230 VTAIL.n76 VTAIL.n75 2.71565
R231 VTAIL.n152 VTAIL.n142 1.93989
R232 VTAIL.n12 VTAIL.n2 1.93989
R233 VTAIL.n32 VTAIL.n22 1.93989
R234 VTAIL.n52 VTAIL.n42 1.93989
R235 VTAIL.n132 VTAIL.n122 1.93989
R236 VTAIL.n112 VTAIL.n102 1.93989
R237 VTAIL.n92 VTAIL.n82 1.93989
R238 VTAIL.n72 VTAIL.n62 1.93989
R239 VTAIL VTAIL.n19 1.8949
R240 VTAIL VTAIL.n159 1.77852
R241 VTAIL.n151 VTAIL.n144 1.16414
R242 VTAIL.n11 VTAIL.n4 1.16414
R243 VTAIL.n31 VTAIL.n24 1.16414
R244 VTAIL.n51 VTAIL.n44 1.16414
R245 VTAIL.n131 VTAIL.n124 1.16414
R246 VTAIL.n111 VTAIL.n104 1.16414
R247 VTAIL.n91 VTAIL.n84 1.16414
R248 VTAIL.n71 VTAIL.n64 1.16414
R249 VTAIL.n119 VTAIL.n99 0.470328
R250 VTAIL.n39 VTAIL.n19 0.470328
R251 VTAIL.n148 VTAIL.n147 0.388379
R252 VTAIL.n8 VTAIL.n7 0.388379
R253 VTAIL.n28 VTAIL.n27 0.388379
R254 VTAIL.n48 VTAIL.n47 0.388379
R255 VTAIL.n128 VTAIL.n127 0.388379
R256 VTAIL.n108 VTAIL.n107 0.388379
R257 VTAIL.n88 VTAIL.n87 0.388379
R258 VTAIL.n68 VTAIL.n67 0.388379
R259 VTAIL.n150 VTAIL.n149 0.155672
R260 VTAIL.n150 VTAIL.n141 0.155672
R261 VTAIL.n157 VTAIL.n141 0.155672
R262 VTAIL.n10 VTAIL.n9 0.155672
R263 VTAIL.n10 VTAIL.n1 0.155672
R264 VTAIL.n17 VTAIL.n1 0.155672
R265 VTAIL.n30 VTAIL.n29 0.155672
R266 VTAIL.n30 VTAIL.n21 0.155672
R267 VTAIL.n37 VTAIL.n21 0.155672
R268 VTAIL.n50 VTAIL.n49 0.155672
R269 VTAIL.n50 VTAIL.n41 0.155672
R270 VTAIL.n57 VTAIL.n41 0.155672
R271 VTAIL.n137 VTAIL.n121 0.155672
R272 VTAIL.n130 VTAIL.n121 0.155672
R273 VTAIL.n130 VTAIL.n129 0.155672
R274 VTAIL.n117 VTAIL.n101 0.155672
R275 VTAIL.n110 VTAIL.n101 0.155672
R276 VTAIL.n110 VTAIL.n109 0.155672
R277 VTAIL.n97 VTAIL.n81 0.155672
R278 VTAIL.n90 VTAIL.n81 0.155672
R279 VTAIL.n90 VTAIL.n89 0.155672
R280 VTAIL.n77 VTAIL.n61 0.155672
R281 VTAIL.n70 VTAIL.n61 0.155672
R282 VTAIL.n70 VTAIL.n69 0.155672
R283 VDD1 VDD1.n1 156.389
R284 VDD1 VDD1.n0 117.7
R285 VDD1.n0 VDD1.t0 8.02643
R286 VDD1.n0 VDD1.t2 8.02643
R287 VDD1.n1 VDD1.t1 8.02643
R288 VDD1.n1 VDD1.t3 8.02643
R289 VN.n0 VN.t1 58.6622
R290 VN.n1 VN.t2 58.6622
R291 VN.n0 VN.t3 57.235
R292 VN.n1 VN.t0 57.235
R293 VN VN.n1 46.275
R294 VN VN.n0 1.78636
R295 VDD2.n2 VDD2.n0 155.864
R296 VDD2.n2 VDD2.n1 117.641
R297 VDD2.n1 VDD2.t3 8.02643
R298 VDD2.n1 VDD2.t1 8.02643
R299 VDD2.n0 VDD2.t2 8.02643
R300 VDD2.n0 VDD2.t0 8.02643
R301 VDD2 VDD2.n2 0.0586897
R302 B.n284 B.n283 585
R303 B.n282 B.n99 585
R304 B.n281 B.n280 585
R305 B.n279 B.n100 585
R306 B.n278 B.n277 585
R307 B.n276 B.n101 585
R308 B.n275 B.n274 585
R309 B.n273 B.n102 585
R310 B.n272 B.n271 585
R311 B.n270 B.n103 585
R312 B.n269 B.n268 585
R313 B.n267 B.n104 585
R314 B.n266 B.n265 585
R315 B.n264 B.n105 585
R316 B.n263 B.n262 585
R317 B.n261 B.n106 585
R318 B.n260 B.n259 585
R319 B.n258 B.n107 585
R320 B.n257 B.n256 585
R321 B.n252 B.n108 585
R322 B.n251 B.n250 585
R323 B.n249 B.n109 585
R324 B.n248 B.n247 585
R325 B.n246 B.n110 585
R326 B.n245 B.n244 585
R327 B.n243 B.n111 585
R328 B.n242 B.n241 585
R329 B.n240 B.n112 585
R330 B.n238 B.n237 585
R331 B.n236 B.n115 585
R332 B.n235 B.n234 585
R333 B.n233 B.n116 585
R334 B.n232 B.n231 585
R335 B.n230 B.n117 585
R336 B.n229 B.n228 585
R337 B.n227 B.n118 585
R338 B.n226 B.n225 585
R339 B.n224 B.n119 585
R340 B.n223 B.n222 585
R341 B.n221 B.n120 585
R342 B.n220 B.n219 585
R343 B.n218 B.n121 585
R344 B.n217 B.n216 585
R345 B.n215 B.n122 585
R346 B.n214 B.n213 585
R347 B.n212 B.n123 585
R348 B.n285 B.n98 585
R349 B.n287 B.n286 585
R350 B.n288 B.n97 585
R351 B.n290 B.n289 585
R352 B.n291 B.n96 585
R353 B.n293 B.n292 585
R354 B.n294 B.n95 585
R355 B.n296 B.n295 585
R356 B.n297 B.n94 585
R357 B.n299 B.n298 585
R358 B.n300 B.n93 585
R359 B.n302 B.n301 585
R360 B.n303 B.n92 585
R361 B.n305 B.n304 585
R362 B.n306 B.n91 585
R363 B.n308 B.n307 585
R364 B.n309 B.n90 585
R365 B.n311 B.n310 585
R366 B.n312 B.n89 585
R367 B.n314 B.n313 585
R368 B.n315 B.n88 585
R369 B.n317 B.n316 585
R370 B.n318 B.n87 585
R371 B.n320 B.n319 585
R372 B.n321 B.n86 585
R373 B.n323 B.n322 585
R374 B.n324 B.n85 585
R375 B.n326 B.n325 585
R376 B.n327 B.n84 585
R377 B.n329 B.n328 585
R378 B.n330 B.n83 585
R379 B.n332 B.n331 585
R380 B.n333 B.n82 585
R381 B.n335 B.n334 585
R382 B.n336 B.n81 585
R383 B.n338 B.n337 585
R384 B.n339 B.n80 585
R385 B.n341 B.n340 585
R386 B.n342 B.n79 585
R387 B.n344 B.n343 585
R388 B.n345 B.n78 585
R389 B.n347 B.n346 585
R390 B.n348 B.n77 585
R391 B.n350 B.n349 585
R392 B.n351 B.n76 585
R393 B.n353 B.n352 585
R394 B.n354 B.n75 585
R395 B.n356 B.n355 585
R396 B.n357 B.n74 585
R397 B.n359 B.n358 585
R398 B.n360 B.n73 585
R399 B.n362 B.n361 585
R400 B.n363 B.n72 585
R401 B.n365 B.n364 585
R402 B.n366 B.n71 585
R403 B.n368 B.n367 585
R404 B.n369 B.n70 585
R405 B.n371 B.n370 585
R406 B.n372 B.n69 585
R407 B.n374 B.n373 585
R408 B.n375 B.n68 585
R409 B.n377 B.n376 585
R410 B.n378 B.n67 585
R411 B.n380 B.n379 585
R412 B.n381 B.n66 585
R413 B.n383 B.n382 585
R414 B.n384 B.n65 585
R415 B.n386 B.n385 585
R416 B.n387 B.n64 585
R417 B.n389 B.n388 585
R418 B.n390 B.n63 585
R419 B.n392 B.n391 585
R420 B.n393 B.n62 585
R421 B.n395 B.n394 585
R422 B.n396 B.n61 585
R423 B.n398 B.n397 585
R424 B.n399 B.n60 585
R425 B.n401 B.n400 585
R426 B.n402 B.n59 585
R427 B.n404 B.n403 585
R428 B.n405 B.n58 585
R429 B.n407 B.n406 585
R430 B.n408 B.n57 585
R431 B.n410 B.n409 585
R432 B.n411 B.n56 585
R433 B.n413 B.n412 585
R434 B.n414 B.n55 585
R435 B.n416 B.n415 585
R436 B.n417 B.n54 585
R437 B.n419 B.n418 585
R438 B.n420 B.n53 585
R439 B.n422 B.n421 585
R440 B.n492 B.n491 585
R441 B.n490 B.n25 585
R442 B.n489 B.n488 585
R443 B.n487 B.n26 585
R444 B.n486 B.n485 585
R445 B.n484 B.n27 585
R446 B.n483 B.n482 585
R447 B.n481 B.n28 585
R448 B.n480 B.n479 585
R449 B.n478 B.n29 585
R450 B.n477 B.n476 585
R451 B.n475 B.n30 585
R452 B.n474 B.n473 585
R453 B.n472 B.n31 585
R454 B.n471 B.n470 585
R455 B.n469 B.n32 585
R456 B.n468 B.n467 585
R457 B.n466 B.n33 585
R458 B.n464 B.n463 585
R459 B.n462 B.n36 585
R460 B.n461 B.n460 585
R461 B.n459 B.n37 585
R462 B.n458 B.n457 585
R463 B.n456 B.n38 585
R464 B.n455 B.n454 585
R465 B.n453 B.n39 585
R466 B.n452 B.n451 585
R467 B.n450 B.n40 585
R468 B.n449 B.n448 585
R469 B.n447 B.n41 585
R470 B.n446 B.n445 585
R471 B.n444 B.n45 585
R472 B.n443 B.n442 585
R473 B.n441 B.n46 585
R474 B.n440 B.n439 585
R475 B.n438 B.n47 585
R476 B.n437 B.n436 585
R477 B.n435 B.n48 585
R478 B.n434 B.n433 585
R479 B.n432 B.n49 585
R480 B.n431 B.n430 585
R481 B.n429 B.n50 585
R482 B.n428 B.n427 585
R483 B.n426 B.n51 585
R484 B.n425 B.n424 585
R485 B.n423 B.n52 585
R486 B.n493 B.n24 585
R487 B.n495 B.n494 585
R488 B.n496 B.n23 585
R489 B.n498 B.n497 585
R490 B.n499 B.n22 585
R491 B.n501 B.n500 585
R492 B.n502 B.n21 585
R493 B.n504 B.n503 585
R494 B.n505 B.n20 585
R495 B.n507 B.n506 585
R496 B.n508 B.n19 585
R497 B.n510 B.n509 585
R498 B.n511 B.n18 585
R499 B.n513 B.n512 585
R500 B.n514 B.n17 585
R501 B.n516 B.n515 585
R502 B.n517 B.n16 585
R503 B.n519 B.n518 585
R504 B.n520 B.n15 585
R505 B.n522 B.n521 585
R506 B.n523 B.n14 585
R507 B.n525 B.n524 585
R508 B.n526 B.n13 585
R509 B.n528 B.n527 585
R510 B.n529 B.n12 585
R511 B.n531 B.n530 585
R512 B.n532 B.n11 585
R513 B.n534 B.n533 585
R514 B.n535 B.n10 585
R515 B.n537 B.n536 585
R516 B.n538 B.n9 585
R517 B.n540 B.n539 585
R518 B.n541 B.n8 585
R519 B.n543 B.n542 585
R520 B.n544 B.n7 585
R521 B.n546 B.n545 585
R522 B.n547 B.n6 585
R523 B.n549 B.n548 585
R524 B.n550 B.n5 585
R525 B.n552 B.n551 585
R526 B.n553 B.n4 585
R527 B.n555 B.n554 585
R528 B.n556 B.n3 585
R529 B.n558 B.n557 585
R530 B.n559 B.n0 585
R531 B.n2 B.n1 585
R532 B.n146 B.n145 585
R533 B.n148 B.n147 585
R534 B.n149 B.n144 585
R535 B.n151 B.n150 585
R536 B.n152 B.n143 585
R537 B.n154 B.n153 585
R538 B.n155 B.n142 585
R539 B.n157 B.n156 585
R540 B.n158 B.n141 585
R541 B.n160 B.n159 585
R542 B.n161 B.n140 585
R543 B.n163 B.n162 585
R544 B.n164 B.n139 585
R545 B.n166 B.n165 585
R546 B.n167 B.n138 585
R547 B.n169 B.n168 585
R548 B.n170 B.n137 585
R549 B.n172 B.n171 585
R550 B.n173 B.n136 585
R551 B.n175 B.n174 585
R552 B.n176 B.n135 585
R553 B.n178 B.n177 585
R554 B.n179 B.n134 585
R555 B.n181 B.n180 585
R556 B.n182 B.n133 585
R557 B.n184 B.n183 585
R558 B.n185 B.n132 585
R559 B.n187 B.n186 585
R560 B.n188 B.n131 585
R561 B.n190 B.n189 585
R562 B.n191 B.n130 585
R563 B.n193 B.n192 585
R564 B.n194 B.n129 585
R565 B.n196 B.n195 585
R566 B.n197 B.n128 585
R567 B.n199 B.n198 585
R568 B.n200 B.n127 585
R569 B.n202 B.n201 585
R570 B.n203 B.n126 585
R571 B.n205 B.n204 585
R572 B.n206 B.n125 585
R573 B.n208 B.n207 585
R574 B.n209 B.n124 585
R575 B.n211 B.n210 585
R576 B.n212 B.n211 535.745
R577 B.n283 B.n98 535.745
R578 B.n421 B.n52 535.745
R579 B.n493 B.n492 535.745
R580 B.n253 B.t10 319.217
R581 B.n42 B.t2 319.217
R582 B.n113 B.t7 319.217
R583 B.n34 B.t5 319.217
R584 B.n561 B.n560 256.663
R585 B.n254 B.t11 236.6
R586 B.n43 B.t1 236.6
R587 B.n114 B.t8 236.6
R588 B.n35 B.t4 236.6
R589 B.n560 B.n559 235.042
R590 B.n560 B.n2 235.042
R591 B.n113 B.t6 234.278
R592 B.n253 B.t9 234.278
R593 B.n42 B.t0 234.278
R594 B.n34 B.t3 234.278
R595 B.n213 B.n212 163.367
R596 B.n213 B.n122 163.367
R597 B.n217 B.n122 163.367
R598 B.n218 B.n217 163.367
R599 B.n219 B.n218 163.367
R600 B.n219 B.n120 163.367
R601 B.n223 B.n120 163.367
R602 B.n224 B.n223 163.367
R603 B.n225 B.n224 163.367
R604 B.n225 B.n118 163.367
R605 B.n229 B.n118 163.367
R606 B.n230 B.n229 163.367
R607 B.n231 B.n230 163.367
R608 B.n231 B.n116 163.367
R609 B.n235 B.n116 163.367
R610 B.n236 B.n235 163.367
R611 B.n237 B.n236 163.367
R612 B.n237 B.n112 163.367
R613 B.n242 B.n112 163.367
R614 B.n243 B.n242 163.367
R615 B.n244 B.n243 163.367
R616 B.n244 B.n110 163.367
R617 B.n248 B.n110 163.367
R618 B.n249 B.n248 163.367
R619 B.n250 B.n249 163.367
R620 B.n250 B.n108 163.367
R621 B.n257 B.n108 163.367
R622 B.n258 B.n257 163.367
R623 B.n259 B.n258 163.367
R624 B.n259 B.n106 163.367
R625 B.n263 B.n106 163.367
R626 B.n264 B.n263 163.367
R627 B.n265 B.n264 163.367
R628 B.n265 B.n104 163.367
R629 B.n269 B.n104 163.367
R630 B.n270 B.n269 163.367
R631 B.n271 B.n270 163.367
R632 B.n271 B.n102 163.367
R633 B.n275 B.n102 163.367
R634 B.n276 B.n275 163.367
R635 B.n277 B.n276 163.367
R636 B.n277 B.n100 163.367
R637 B.n281 B.n100 163.367
R638 B.n282 B.n281 163.367
R639 B.n283 B.n282 163.367
R640 B.n421 B.n420 163.367
R641 B.n420 B.n419 163.367
R642 B.n419 B.n54 163.367
R643 B.n415 B.n54 163.367
R644 B.n415 B.n414 163.367
R645 B.n414 B.n413 163.367
R646 B.n413 B.n56 163.367
R647 B.n409 B.n56 163.367
R648 B.n409 B.n408 163.367
R649 B.n408 B.n407 163.367
R650 B.n407 B.n58 163.367
R651 B.n403 B.n58 163.367
R652 B.n403 B.n402 163.367
R653 B.n402 B.n401 163.367
R654 B.n401 B.n60 163.367
R655 B.n397 B.n60 163.367
R656 B.n397 B.n396 163.367
R657 B.n396 B.n395 163.367
R658 B.n395 B.n62 163.367
R659 B.n391 B.n62 163.367
R660 B.n391 B.n390 163.367
R661 B.n390 B.n389 163.367
R662 B.n389 B.n64 163.367
R663 B.n385 B.n64 163.367
R664 B.n385 B.n384 163.367
R665 B.n384 B.n383 163.367
R666 B.n383 B.n66 163.367
R667 B.n379 B.n66 163.367
R668 B.n379 B.n378 163.367
R669 B.n378 B.n377 163.367
R670 B.n377 B.n68 163.367
R671 B.n373 B.n68 163.367
R672 B.n373 B.n372 163.367
R673 B.n372 B.n371 163.367
R674 B.n371 B.n70 163.367
R675 B.n367 B.n70 163.367
R676 B.n367 B.n366 163.367
R677 B.n366 B.n365 163.367
R678 B.n365 B.n72 163.367
R679 B.n361 B.n72 163.367
R680 B.n361 B.n360 163.367
R681 B.n360 B.n359 163.367
R682 B.n359 B.n74 163.367
R683 B.n355 B.n74 163.367
R684 B.n355 B.n354 163.367
R685 B.n354 B.n353 163.367
R686 B.n353 B.n76 163.367
R687 B.n349 B.n76 163.367
R688 B.n349 B.n348 163.367
R689 B.n348 B.n347 163.367
R690 B.n347 B.n78 163.367
R691 B.n343 B.n78 163.367
R692 B.n343 B.n342 163.367
R693 B.n342 B.n341 163.367
R694 B.n341 B.n80 163.367
R695 B.n337 B.n80 163.367
R696 B.n337 B.n336 163.367
R697 B.n336 B.n335 163.367
R698 B.n335 B.n82 163.367
R699 B.n331 B.n82 163.367
R700 B.n331 B.n330 163.367
R701 B.n330 B.n329 163.367
R702 B.n329 B.n84 163.367
R703 B.n325 B.n84 163.367
R704 B.n325 B.n324 163.367
R705 B.n324 B.n323 163.367
R706 B.n323 B.n86 163.367
R707 B.n319 B.n86 163.367
R708 B.n319 B.n318 163.367
R709 B.n318 B.n317 163.367
R710 B.n317 B.n88 163.367
R711 B.n313 B.n88 163.367
R712 B.n313 B.n312 163.367
R713 B.n312 B.n311 163.367
R714 B.n311 B.n90 163.367
R715 B.n307 B.n90 163.367
R716 B.n307 B.n306 163.367
R717 B.n306 B.n305 163.367
R718 B.n305 B.n92 163.367
R719 B.n301 B.n92 163.367
R720 B.n301 B.n300 163.367
R721 B.n300 B.n299 163.367
R722 B.n299 B.n94 163.367
R723 B.n295 B.n94 163.367
R724 B.n295 B.n294 163.367
R725 B.n294 B.n293 163.367
R726 B.n293 B.n96 163.367
R727 B.n289 B.n96 163.367
R728 B.n289 B.n288 163.367
R729 B.n288 B.n287 163.367
R730 B.n287 B.n98 163.367
R731 B.n492 B.n25 163.367
R732 B.n488 B.n25 163.367
R733 B.n488 B.n487 163.367
R734 B.n487 B.n486 163.367
R735 B.n486 B.n27 163.367
R736 B.n482 B.n27 163.367
R737 B.n482 B.n481 163.367
R738 B.n481 B.n480 163.367
R739 B.n480 B.n29 163.367
R740 B.n476 B.n29 163.367
R741 B.n476 B.n475 163.367
R742 B.n475 B.n474 163.367
R743 B.n474 B.n31 163.367
R744 B.n470 B.n31 163.367
R745 B.n470 B.n469 163.367
R746 B.n469 B.n468 163.367
R747 B.n468 B.n33 163.367
R748 B.n463 B.n33 163.367
R749 B.n463 B.n462 163.367
R750 B.n462 B.n461 163.367
R751 B.n461 B.n37 163.367
R752 B.n457 B.n37 163.367
R753 B.n457 B.n456 163.367
R754 B.n456 B.n455 163.367
R755 B.n455 B.n39 163.367
R756 B.n451 B.n39 163.367
R757 B.n451 B.n450 163.367
R758 B.n450 B.n449 163.367
R759 B.n449 B.n41 163.367
R760 B.n445 B.n41 163.367
R761 B.n445 B.n444 163.367
R762 B.n444 B.n443 163.367
R763 B.n443 B.n46 163.367
R764 B.n439 B.n46 163.367
R765 B.n439 B.n438 163.367
R766 B.n438 B.n437 163.367
R767 B.n437 B.n48 163.367
R768 B.n433 B.n48 163.367
R769 B.n433 B.n432 163.367
R770 B.n432 B.n431 163.367
R771 B.n431 B.n50 163.367
R772 B.n427 B.n50 163.367
R773 B.n427 B.n426 163.367
R774 B.n426 B.n425 163.367
R775 B.n425 B.n52 163.367
R776 B.n494 B.n493 163.367
R777 B.n494 B.n23 163.367
R778 B.n498 B.n23 163.367
R779 B.n499 B.n498 163.367
R780 B.n500 B.n499 163.367
R781 B.n500 B.n21 163.367
R782 B.n504 B.n21 163.367
R783 B.n505 B.n504 163.367
R784 B.n506 B.n505 163.367
R785 B.n506 B.n19 163.367
R786 B.n510 B.n19 163.367
R787 B.n511 B.n510 163.367
R788 B.n512 B.n511 163.367
R789 B.n512 B.n17 163.367
R790 B.n516 B.n17 163.367
R791 B.n517 B.n516 163.367
R792 B.n518 B.n517 163.367
R793 B.n518 B.n15 163.367
R794 B.n522 B.n15 163.367
R795 B.n523 B.n522 163.367
R796 B.n524 B.n523 163.367
R797 B.n524 B.n13 163.367
R798 B.n528 B.n13 163.367
R799 B.n529 B.n528 163.367
R800 B.n530 B.n529 163.367
R801 B.n530 B.n11 163.367
R802 B.n534 B.n11 163.367
R803 B.n535 B.n534 163.367
R804 B.n536 B.n535 163.367
R805 B.n536 B.n9 163.367
R806 B.n540 B.n9 163.367
R807 B.n541 B.n540 163.367
R808 B.n542 B.n541 163.367
R809 B.n542 B.n7 163.367
R810 B.n546 B.n7 163.367
R811 B.n547 B.n546 163.367
R812 B.n548 B.n547 163.367
R813 B.n548 B.n5 163.367
R814 B.n552 B.n5 163.367
R815 B.n553 B.n552 163.367
R816 B.n554 B.n553 163.367
R817 B.n554 B.n3 163.367
R818 B.n558 B.n3 163.367
R819 B.n559 B.n558 163.367
R820 B.n146 B.n2 163.367
R821 B.n147 B.n146 163.367
R822 B.n147 B.n144 163.367
R823 B.n151 B.n144 163.367
R824 B.n152 B.n151 163.367
R825 B.n153 B.n152 163.367
R826 B.n153 B.n142 163.367
R827 B.n157 B.n142 163.367
R828 B.n158 B.n157 163.367
R829 B.n159 B.n158 163.367
R830 B.n159 B.n140 163.367
R831 B.n163 B.n140 163.367
R832 B.n164 B.n163 163.367
R833 B.n165 B.n164 163.367
R834 B.n165 B.n138 163.367
R835 B.n169 B.n138 163.367
R836 B.n170 B.n169 163.367
R837 B.n171 B.n170 163.367
R838 B.n171 B.n136 163.367
R839 B.n175 B.n136 163.367
R840 B.n176 B.n175 163.367
R841 B.n177 B.n176 163.367
R842 B.n177 B.n134 163.367
R843 B.n181 B.n134 163.367
R844 B.n182 B.n181 163.367
R845 B.n183 B.n182 163.367
R846 B.n183 B.n132 163.367
R847 B.n187 B.n132 163.367
R848 B.n188 B.n187 163.367
R849 B.n189 B.n188 163.367
R850 B.n189 B.n130 163.367
R851 B.n193 B.n130 163.367
R852 B.n194 B.n193 163.367
R853 B.n195 B.n194 163.367
R854 B.n195 B.n128 163.367
R855 B.n199 B.n128 163.367
R856 B.n200 B.n199 163.367
R857 B.n201 B.n200 163.367
R858 B.n201 B.n126 163.367
R859 B.n205 B.n126 163.367
R860 B.n206 B.n205 163.367
R861 B.n207 B.n206 163.367
R862 B.n207 B.n124 163.367
R863 B.n211 B.n124 163.367
R864 B.n114 B.n113 82.6187
R865 B.n254 B.n253 82.6187
R866 B.n43 B.n42 82.6187
R867 B.n35 B.n34 82.6187
R868 B.n239 B.n114 59.5399
R869 B.n255 B.n254 59.5399
R870 B.n44 B.n43 59.5399
R871 B.n465 B.n35 59.5399
R872 B.n491 B.n24 34.8103
R873 B.n423 B.n422 34.8103
R874 B.n285 B.n284 34.8103
R875 B.n210 B.n123 34.8103
R876 B B.n561 18.0485
R877 B.n495 B.n24 10.6151
R878 B.n496 B.n495 10.6151
R879 B.n497 B.n496 10.6151
R880 B.n497 B.n22 10.6151
R881 B.n501 B.n22 10.6151
R882 B.n502 B.n501 10.6151
R883 B.n503 B.n502 10.6151
R884 B.n503 B.n20 10.6151
R885 B.n507 B.n20 10.6151
R886 B.n508 B.n507 10.6151
R887 B.n509 B.n508 10.6151
R888 B.n509 B.n18 10.6151
R889 B.n513 B.n18 10.6151
R890 B.n514 B.n513 10.6151
R891 B.n515 B.n514 10.6151
R892 B.n515 B.n16 10.6151
R893 B.n519 B.n16 10.6151
R894 B.n520 B.n519 10.6151
R895 B.n521 B.n520 10.6151
R896 B.n521 B.n14 10.6151
R897 B.n525 B.n14 10.6151
R898 B.n526 B.n525 10.6151
R899 B.n527 B.n526 10.6151
R900 B.n527 B.n12 10.6151
R901 B.n531 B.n12 10.6151
R902 B.n532 B.n531 10.6151
R903 B.n533 B.n532 10.6151
R904 B.n533 B.n10 10.6151
R905 B.n537 B.n10 10.6151
R906 B.n538 B.n537 10.6151
R907 B.n539 B.n538 10.6151
R908 B.n539 B.n8 10.6151
R909 B.n543 B.n8 10.6151
R910 B.n544 B.n543 10.6151
R911 B.n545 B.n544 10.6151
R912 B.n545 B.n6 10.6151
R913 B.n549 B.n6 10.6151
R914 B.n550 B.n549 10.6151
R915 B.n551 B.n550 10.6151
R916 B.n551 B.n4 10.6151
R917 B.n555 B.n4 10.6151
R918 B.n556 B.n555 10.6151
R919 B.n557 B.n556 10.6151
R920 B.n557 B.n0 10.6151
R921 B.n491 B.n490 10.6151
R922 B.n490 B.n489 10.6151
R923 B.n489 B.n26 10.6151
R924 B.n485 B.n26 10.6151
R925 B.n485 B.n484 10.6151
R926 B.n484 B.n483 10.6151
R927 B.n483 B.n28 10.6151
R928 B.n479 B.n28 10.6151
R929 B.n479 B.n478 10.6151
R930 B.n478 B.n477 10.6151
R931 B.n477 B.n30 10.6151
R932 B.n473 B.n30 10.6151
R933 B.n473 B.n472 10.6151
R934 B.n472 B.n471 10.6151
R935 B.n471 B.n32 10.6151
R936 B.n467 B.n32 10.6151
R937 B.n467 B.n466 10.6151
R938 B.n464 B.n36 10.6151
R939 B.n460 B.n36 10.6151
R940 B.n460 B.n459 10.6151
R941 B.n459 B.n458 10.6151
R942 B.n458 B.n38 10.6151
R943 B.n454 B.n38 10.6151
R944 B.n454 B.n453 10.6151
R945 B.n453 B.n452 10.6151
R946 B.n452 B.n40 10.6151
R947 B.n448 B.n447 10.6151
R948 B.n447 B.n446 10.6151
R949 B.n446 B.n45 10.6151
R950 B.n442 B.n45 10.6151
R951 B.n442 B.n441 10.6151
R952 B.n441 B.n440 10.6151
R953 B.n440 B.n47 10.6151
R954 B.n436 B.n47 10.6151
R955 B.n436 B.n435 10.6151
R956 B.n435 B.n434 10.6151
R957 B.n434 B.n49 10.6151
R958 B.n430 B.n49 10.6151
R959 B.n430 B.n429 10.6151
R960 B.n429 B.n428 10.6151
R961 B.n428 B.n51 10.6151
R962 B.n424 B.n51 10.6151
R963 B.n424 B.n423 10.6151
R964 B.n422 B.n53 10.6151
R965 B.n418 B.n53 10.6151
R966 B.n418 B.n417 10.6151
R967 B.n417 B.n416 10.6151
R968 B.n416 B.n55 10.6151
R969 B.n412 B.n55 10.6151
R970 B.n412 B.n411 10.6151
R971 B.n411 B.n410 10.6151
R972 B.n410 B.n57 10.6151
R973 B.n406 B.n57 10.6151
R974 B.n406 B.n405 10.6151
R975 B.n405 B.n404 10.6151
R976 B.n404 B.n59 10.6151
R977 B.n400 B.n59 10.6151
R978 B.n400 B.n399 10.6151
R979 B.n399 B.n398 10.6151
R980 B.n398 B.n61 10.6151
R981 B.n394 B.n61 10.6151
R982 B.n394 B.n393 10.6151
R983 B.n393 B.n392 10.6151
R984 B.n392 B.n63 10.6151
R985 B.n388 B.n63 10.6151
R986 B.n388 B.n387 10.6151
R987 B.n387 B.n386 10.6151
R988 B.n386 B.n65 10.6151
R989 B.n382 B.n65 10.6151
R990 B.n382 B.n381 10.6151
R991 B.n381 B.n380 10.6151
R992 B.n380 B.n67 10.6151
R993 B.n376 B.n67 10.6151
R994 B.n376 B.n375 10.6151
R995 B.n375 B.n374 10.6151
R996 B.n374 B.n69 10.6151
R997 B.n370 B.n69 10.6151
R998 B.n370 B.n369 10.6151
R999 B.n369 B.n368 10.6151
R1000 B.n368 B.n71 10.6151
R1001 B.n364 B.n71 10.6151
R1002 B.n364 B.n363 10.6151
R1003 B.n363 B.n362 10.6151
R1004 B.n362 B.n73 10.6151
R1005 B.n358 B.n73 10.6151
R1006 B.n358 B.n357 10.6151
R1007 B.n357 B.n356 10.6151
R1008 B.n356 B.n75 10.6151
R1009 B.n352 B.n75 10.6151
R1010 B.n352 B.n351 10.6151
R1011 B.n351 B.n350 10.6151
R1012 B.n350 B.n77 10.6151
R1013 B.n346 B.n77 10.6151
R1014 B.n346 B.n345 10.6151
R1015 B.n345 B.n344 10.6151
R1016 B.n344 B.n79 10.6151
R1017 B.n340 B.n79 10.6151
R1018 B.n340 B.n339 10.6151
R1019 B.n339 B.n338 10.6151
R1020 B.n338 B.n81 10.6151
R1021 B.n334 B.n81 10.6151
R1022 B.n334 B.n333 10.6151
R1023 B.n333 B.n332 10.6151
R1024 B.n332 B.n83 10.6151
R1025 B.n328 B.n83 10.6151
R1026 B.n328 B.n327 10.6151
R1027 B.n327 B.n326 10.6151
R1028 B.n326 B.n85 10.6151
R1029 B.n322 B.n85 10.6151
R1030 B.n322 B.n321 10.6151
R1031 B.n321 B.n320 10.6151
R1032 B.n320 B.n87 10.6151
R1033 B.n316 B.n87 10.6151
R1034 B.n316 B.n315 10.6151
R1035 B.n315 B.n314 10.6151
R1036 B.n314 B.n89 10.6151
R1037 B.n310 B.n89 10.6151
R1038 B.n310 B.n309 10.6151
R1039 B.n309 B.n308 10.6151
R1040 B.n308 B.n91 10.6151
R1041 B.n304 B.n91 10.6151
R1042 B.n304 B.n303 10.6151
R1043 B.n303 B.n302 10.6151
R1044 B.n302 B.n93 10.6151
R1045 B.n298 B.n93 10.6151
R1046 B.n298 B.n297 10.6151
R1047 B.n297 B.n296 10.6151
R1048 B.n296 B.n95 10.6151
R1049 B.n292 B.n95 10.6151
R1050 B.n292 B.n291 10.6151
R1051 B.n291 B.n290 10.6151
R1052 B.n290 B.n97 10.6151
R1053 B.n286 B.n97 10.6151
R1054 B.n286 B.n285 10.6151
R1055 B.n145 B.n1 10.6151
R1056 B.n148 B.n145 10.6151
R1057 B.n149 B.n148 10.6151
R1058 B.n150 B.n149 10.6151
R1059 B.n150 B.n143 10.6151
R1060 B.n154 B.n143 10.6151
R1061 B.n155 B.n154 10.6151
R1062 B.n156 B.n155 10.6151
R1063 B.n156 B.n141 10.6151
R1064 B.n160 B.n141 10.6151
R1065 B.n161 B.n160 10.6151
R1066 B.n162 B.n161 10.6151
R1067 B.n162 B.n139 10.6151
R1068 B.n166 B.n139 10.6151
R1069 B.n167 B.n166 10.6151
R1070 B.n168 B.n167 10.6151
R1071 B.n168 B.n137 10.6151
R1072 B.n172 B.n137 10.6151
R1073 B.n173 B.n172 10.6151
R1074 B.n174 B.n173 10.6151
R1075 B.n174 B.n135 10.6151
R1076 B.n178 B.n135 10.6151
R1077 B.n179 B.n178 10.6151
R1078 B.n180 B.n179 10.6151
R1079 B.n180 B.n133 10.6151
R1080 B.n184 B.n133 10.6151
R1081 B.n185 B.n184 10.6151
R1082 B.n186 B.n185 10.6151
R1083 B.n186 B.n131 10.6151
R1084 B.n190 B.n131 10.6151
R1085 B.n191 B.n190 10.6151
R1086 B.n192 B.n191 10.6151
R1087 B.n192 B.n129 10.6151
R1088 B.n196 B.n129 10.6151
R1089 B.n197 B.n196 10.6151
R1090 B.n198 B.n197 10.6151
R1091 B.n198 B.n127 10.6151
R1092 B.n202 B.n127 10.6151
R1093 B.n203 B.n202 10.6151
R1094 B.n204 B.n203 10.6151
R1095 B.n204 B.n125 10.6151
R1096 B.n208 B.n125 10.6151
R1097 B.n209 B.n208 10.6151
R1098 B.n210 B.n209 10.6151
R1099 B.n214 B.n123 10.6151
R1100 B.n215 B.n214 10.6151
R1101 B.n216 B.n215 10.6151
R1102 B.n216 B.n121 10.6151
R1103 B.n220 B.n121 10.6151
R1104 B.n221 B.n220 10.6151
R1105 B.n222 B.n221 10.6151
R1106 B.n222 B.n119 10.6151
R1107 B.n226 B.n119 10.6151
R1108 B.n227 B.n226 10.6151
R1109 B.n228 B.n227 10.6151
R1110 B.n228 B.n117 10.6151
R1111 B.n232 B.n117 10.6151
R1112 B.n233 B.n232 10.6151
R1113 B.n234 B.n233 10.6151
R1114 B.n234 B.n115 10.6151
R1115 B.n238 B.n115 10.6151
R1116 B.n241 B.n240 10.6151
R1117 B.n241 B.n111 10.6151
R1118 B.n245 B.n111 10.6151
R1119 B.n246 B.n245 10.6151
R1120 B.n247 B.n246 10.6151
R1121 B.n247 B.n109 10.6151
R1122 B.n251 B.n109 10.6151
R1123 B.n252 B.n251 10.6151
R1124 B.n256 B.n252 10.6151
R1125 B.n260 B.n107 10.6151
R1126 B.n261 B.n260 10.6151
R1127 B.n262 B.n261 10.6151
R1128 B.n262 B.n105 10.6151
R1129 B.n266 B.n105 10.6151
R1130 B.n267 B.n266 10.6151
R1131 B.n268 B.n267 10.6151
R1132 B.n268 B.n103 10.6151
R1133 B.n272 B.n103 10.6151
R1134 B.n273 B.n272 10.6151
R1135 B.n274 B.n273 10.6151
R1136 B.n274 B.n101 10.6151
R1137 B.n278 B.n101 10.6151
R1138 B.n279 B.n278 10.6151
R1139 B.n280 B.n279 10.6151
R1140 B.n280 B.n99 10.6151
R1141 B.n284 B.n99 10.6151
R1142 B.n466 B.n465 9.36635
R1143 B.n448 B.n44 9.36635
R1144 B.n239 B.n238 9.36635
R1145 B.n255 B.n107 9.36635
R1146 B.n561 B.n0 8.11757
R1147 B.n561 B.n1 8.11757
R1148 B.n465 B.n464 1.24928
R1149 B.n44 B.n40 1.24928
R1150 B.n240 B.n239 1.24928
R1151 B.n256 B.n255 1.24928
C0 B VDD1 1.28335f
C1 VN VTAIL 2.61746f
C2 VP VTAIL 2.63157f
C3 VDD2 VN 1.92658f
C4 VN B 1.27688f
C5 VDD2 VP 0.48385f
C6 w_n3526_n1778# VDD1 1.48869f
C7 B VP 2.04067f
C8 VN w_n3526_n1778# 6.08236f
C9 VDD2 VTAIL 4.22333f
C10 VN VDD1 0.154591f
C11 B VTAIL 2.65456f
C12 VP w_n3526_n1778# 6.53818f
C13 VP VDD1 2.25414f
C14 VDD2 B 1.35771f
C15 VN VP 5.68733f
C16 w_n3526_n1778# VTAIL 2.28145f
C17 VDD1 VTAIL 4.16021f
C18 VDD2 w_n3526_n1778# 1.57375f
C19 VDD2 VDD1 1.35367f
C20 B w_n3526_n1778# 8.680719f
C21 VDD2 VSUBS 0.870233f
C22 VDD1 VSUBS 5.69629f
C23 VTAIL VSUBS 0.760694f
C24 VN VSUBS 5.99882f
C25 VP VSUBS 2.516156f
C26 B VSUBS 4.479791f
C27 w_n3526_n1778# VSUBS 78.9119f
C28 B.n0 VSUBS 0.009345f
C29 B.n1 VSUBS 0.009345f
C30 B.n2 VSUBS 0.013821f
C31 B.n3 VSUBS 0.010591f
C32 B.n4 VSUBS 0.010591f
C33 B.n5 VSUBS 0.010591f
C34 B.n6 VSUBS 0.010591f
C35 B.n7 VSUBS 0.010591f
C36 B.n8 VSUBS 0.010591f
C37 B.n9 VSUBS 0.010591f
C38 B.n10 VSUBS 0.010591f
C39 B.n11 VSUBS 0.010591f
C40 B.n12 VSUBS 0.010591f
C41 B.n13 VSUBS 0.010591f
C42 B.n14 VSUBS 0.010591f
C43 B.n15 VSUBS 0.010591f
C44 B.n16 VSUBS 0.010591f
C45 B.n17 VSUBS 0.010591f
C46 B.n18 VSUBS 0.010591f
C47 B.n19 VSUBS 0.010591f
C48 B.n20 VSUBS 0.010591f
C49 B.n21 VSUBS 0.010591f
C50 B.n22 VSUBS 0.010591f
C51 B.n23 VSUBS 0.010591f
C52 B.n24 VSUBS 0.025125f
C53 B.n25 VSUBS 0.010591f
C54 B.n26 VSUBS 0.010591f
C55 B.n27 VSUBS 0.010591f
C56 B.n28 VSUBS 0.010591f
C57 B.n29 VSUBS 0.010591f
C58 B.n30 VSUBS 0.010591f
C59 B.n31 VSUBS 0.010591f
C60 B.n32 VSUBS 0.010591f
C61 B.n33 VSUBS 0.010591f
C62 B.t4 VSUBS 0.089211f
C63 B.t5 VSUBS 0.133066f
C64 B.t3 VSUBS 1.17338f
C65 B.n34 VSUBS 0.223174f
C66 B.n35 VSUBS 0.18455f
C67 B.n36 VSUBS 0.010591f
C68 B.n37 VSUBS 0.010591f
C69 B.n38 VSUBS 0.010591f
C70 B.n39 VSUBS 0.010591f
C71 B.n40 VSUBS 0.005919f
C72 B.n41 VSUBS 0.010591f
C73 B.t1 VSUBS 0.089213f
C74 B.t2 VSUBS 0.133067f
C75 B.t0 VSUBS 1.17338f
C76 B.n42 VSUBS 0.223173f
C77 B.n43 VSUBS 0.184548f
C78 B.n44 VSUBS 0.024539f
C79 B.n45 VSUBS 0.010591f
C80 B.n46 VSUBS 0.010591f
C81 B.n47 VSUBS 0.010591f
C82 B.n48 VSUBS 0.010591f
C83 B.n49 VSUBS 0.010591f
C84 B.n50 VSUBS 0.010591f
C85 B.n51 VSUBS 0.010591f
C86 B.n52 VSUBS 0.026585f
C87 B.n53 VSUBS 0.010591f
C88 B.n54 VSUBS 0.010591f
C89 B.n55 VSUBS 0.010591f
C90 B.n56 VSUBS 0.010591f
C91 B.n57 VSUBS 0.010591f
C92 B.n58 VSUBS 0.010591f
C93 B.n59 VSUBS 0.010591f
C94 B.n60 VSUBS 0.010591f
C95 B.n61 VSUBS 0.010591f
C96 B.n62 VSUBS 0.010591f
C97 B.n63 VSUBS 0.010591f
C98 B.n64 VSUBS 0.010591f
C99 B.n65 VSUBS 0.010591f
C100 B.n66 VSUBS 0.010591f
C101 B.n67 VSUBS 0.010591f
C102 B.n68 VSUBS 0.010591f
C103 B.n69 VSUBS 0.010591f
C104 B.n70 VSUBS 0.010591f
C105 B.n71 VSUBS 0.010591f
C106 B.n72 VSUBS 0.010591f
C107 B.n73 VSUBS 0.010591f
C108 B.n74 VSUBS 0.010591f
C109 B.n75 VSUBS 0.010591f
C110 B.n76 VSUBS 0.010591f
C111 B.n77 VSUBS 0.010591f
C112 B.n78 VSUBS 0.010591f
C113 B.n79 VSUBS 0.010591f
C114 B.n80 VSUBS 0.010591f
C115 B.n81 VSUBS 0.010591f
C116 B.n82 VSUBS 0.010591f
C117 B.n83 VSUBS 0.010591f
C118 B.n84 VSUBS 0.010591f
C119 B.n85 VSUBS 0.010591f
C120 B.n86 VSUBS 0.010591f
C121 B.n87 VSUBS 0.010591f
C122 B.n88 VSUBS 0.010591f
C123 B.n89 VSUBS 0.010591f
C124 B.n90 VSUBS 0.010591f
C125 B.n91 VSUBS 0.010591f
C126 B.n92 VSUBS 0.010591f
C127 B.n93 VSUBS 0.010591f
C128 B.n94 VSUBS 0.010591f
C129 B.n95 VSUBS 0.010591f
C130 B.n96 VSUBS 0.010591f
C131 B.n97 VSUBS 0.010591f
C132 B.n98 VSUBS 0.025125f
C133 B.n99 VSUBS 0.010591f
C134 B.n100 VSUBS 0.010591f
C135 B.n101 VSUBS 0.010591f
C136 B.n102 VSUBS 0.010591f
C137 B.n103 VSUBS 0.010591f
C138 B.n104 VSUBS 0.010591f
C139 B.n105 VSUBS 0.010591f
C140 B.n106 VSUBS 0.010591f
C141 B.n107 VSUBS 0.009968f
C142 B.n108 VSUBS 0.010591f
C143 B.n109 VSUBS 0.010591f
C144 B.n110 VSUBS 0.010591f
C145 B.n111 VSUBS 0.010591f
C146 B.n112 VSUBS 0.010591f
C147 B.t8 VSUBS 0.089211f
C148 B.t7 VSUBS 0.133066f
C149 B.t6 VSUBS 1.17338f
C150 B.n113 VSUBS 0.223174f
C151 B.n114 VSUBS 0.18455f
C152 B.n115 VSUBS 0.010591f
C153 B.n116 VSUBS 0.010591f
C154 B.n117 VSUBS 0.010591f
C155 B.n118 VSUBS 0.010591f
C156 B.n119 VSUBS 0.010591f
C157 B.n120 VSUBS 0.010591f
C158 B.n121 VSUBS 0.010591f
C159 B.n122 VSUBS 0.010591f
C160 B.n123 VSUBS 0.026585f
C161 B.n124 VSUBS 0.010591f
C162 B.n125 VSUBS 0.010591f
C163 B.n126 VSUBS 0.010591f
C164 B.n127 VSUBS 0.010591f
C165 B.n128 VSUBS 0.010591f
C166 B.n129 VSUBS 0.010591f
C167 B.n130 VSUBS 0.010591f
C168 B.n131 VSUBS 0.010591f
C169 B.n132 VSUBS 0.010591f
C170 B.n133 VSUBS 0.010591f
C171 B.n134 VSUBS 0.010591f
C172 B.n135 VSUBS 0.010591f
C173 B.n136 VSUBS 0.010591f
C174 B.n137 VSUBS 0.010591f
C175 B.n138 VSUBS 0.010591f
C176 B.n139 VSUBS 0.010591f
C177 B.n140 VSUBS 0.010591f
C178 B.n141 VSUBS 0.010591f
C179 B.n142 VSUBS 0.010591f
C180 B.n143 VSUBS 0.010591f
C181 B.n144 VSUBS 0.010591f
C182 B.n145 VSUBS 0.010591f
C183 B.n146 VSUBS 0.010591f
C184 B.n147 VSUBS 0.010591f
C185 B.n148 VSUBS 0.010591f
C186 B.n149 VSUBS 0.010591f
C187 B.n150 VSUBS 0.010591f
C188 B.n151 VSUBS 0.010591f
C189 B.n152 VSUBS 0.010591f
C190 B.n153 VSUBS 0.010591f
C191 B.n154 VSUBS 0.010591f
C192 B.n155 VSUBS 0.010591f
C193 B.n156 VSUBS 0.010591f
C194 B.n157 VSUBS 0.010591f
C195 B.n158 VSUBS 0.010591f
C196 B.n159 VSUBS 0.010591f
C197 B.n160 VSUBS 0.010591f
C198 B.n161 VSUBS 0.010591f
C199 B.n162 VSUBS 0.010591f
C200 B.n163 VSUBS 0.010591f
C201 B.n164 VSUBS 0.010591f
C202 B.n165 VSUBS 0.010591f
C203 B.n166 VSUBS 0.010591f
C204 B.n167 VSUBS 0.010591f
C205 B.n168 VSUBS 0.010591f
C206 B.n169 VSUBS 0.010591f
C207 B.n170 VSUBS 0.010591f
C208 B.n171 VSUBS 0.010591f
C209 B.n172 VSUBS 0.010591f
C210 B.n173 VSUBS 0.010591f
C211 B.n174 VSUBS 0.010591f
C212 B.n175 VSUBS 0.010591f
C213 B.n176 VSUBS 0.010591f
C214 B.n177 VSUBS 0.010591f
C215 B.n178 VSUBS 0.010591f
C216 B.n179 VSUBS 0.010591f
C217 B.n180 VSUBS 0.010591f
C218 B.n181 VSUBS 0.010591f
C219 B.n182 VSUBS 0.010591f
C220 B.n183 VSUBS 0.010591f
C221 B.n184 VSUBS 0.010591f
C222 B.n185 VSUBS 0.010591f
C223 B.n186 VSUBS 0.010591f
C224 B.n187 VSUBS 0.010591f
C225 B.n188 VSUBS 0.010591f
C226 B.n189 VSUBS 0.010591f
C227 B.n190 VSUBS 0.010591f
C228 B.n191 VSUBS 0.010591f
C229 B.n192 VSUBS 0.010591f
C230 B.n193 VSUBS 0.010591f
C231 B.n194 VSUBS 0.010591f
C232 B.n195 VSUBS 0.010591f
C233 B.n196 VSUBS 0.010591f
C234 B.n197 VSUBS 0.010591f
C235 B.n198 VSUBS 0.010591f
C236 B.n199 VSUBS 0.010591f
C237 B.n200 VSUBS 0.010591f
C238 B.n201 VSUBS 0.010591f
C239 B.n202 VSUBS 0.010591f
C240 B.n203 VSUBS 0.010591f
C241 B.n204 VSUBS 0.010591f
C242 B.n205 VSUBS 0.010591f
C243 B.n206 VSUBS 0.010591f
C244 B.n207 VSUBS 0.010591f
C245 B.n208 VSUBS 0.010591f
C246 B.n209 VSUBS 0.010591f
C247 B.n210 VSUBS 0.025125f
C248 B.n211 VSUBS 0.025125f
C249 B.n212 VSUBS 0.026585f
C250 B.n213 VSUBS 0.010591f
C251 B.n214 VSUBS 0.010591f
C252 B.n215 VSUBS 0.010591f
C253 B.n216 VSUBS 0.010591f
C254 B.n217 VSUBS 0.010591f
C255 B.n218 VSUBS 0.010591f
C256 B.n219 VSUBS 0.010591f
C257 B.n220 VSUBS 0.010591f
C258 B.n221 VSUBS 0.010591f
C259 B.n222 VSUBS 0.010591f
C260 B.n223 VSUBS 0.010591f
C261 B.n224 VSUBS 0.010591f
C262 B.n225 VSUBS 0.010591f
C263 B.n226 VSUBS 0.010591f
C264 B.n227 VSUBS 0.010591f
C265 B.n228 VSUBS 0.010591f
C266 B.n229 VSUBS 0.010591f
C267 B.n230 VSUBS 0.010591f
C268 B.n231 VSUBS 0.010591f
C269 B.n232 VSUBS 0.010591f
C270 B.n233 VSUBS 0.010591f
C271 B.n234 VSUBS 0.010591f
C272 B.n235 VSUBS 0.010591f
C273 B.n236 VSUBS 0.010591f
C274 B.n237 VSUBS 0.010591f
C275 B.n238 VSUBS 0.009968f
C276 B.n239 VSUBS 0.024539f
C277 B.n240 VSUBS 0.005919f
C278 B.n241 VSUBS 0.010591f
C279 B.n242 VSUBS 0.010591f
C280 B.n243 VSUBS 0.010591f
C281 B.n244 VSUBS 0.010591f
C282 B.n245 VSUBS 0.010591f
C283 B.n246 VSUBS 0.010591f
C284 B.n247 VSUBS 0.010591f
C285 B.n248 VSUBS 0.010591f
C286 B.n249 VSUBS 0.010591f
C287 B.n250 VSUBS 0.010591f
C288 B.n251 VSUBS 0.010591f
C289 B.n252 VSUBS 0.010591f
C290 B.t11 VSUBS 0.089213f
C291 B.t10 VSUBS 0.133067f
C292 B.t9 VSUBS 1.17338f
C293 B.n253 VSUBS 0.223173f
C294 B.n254 VSUBS 0.184548f
C295 B.n255 VSUBS 0.024539f
C296 B.n256 VSUBS 0.005919f
C297 B.n257 VSUBS 0.010591f
C298 B.n258 VSUBS 0.010591f
C299 B.n259 VSUBS 0.010591f
C300 B.n260 VSUBS 0.010591f
C301 B.n261 VSUBS 0.010591f
C302 B.n262 VSUBS 0.010591f
C303 B.n263 VSUBS 0.010591f
C304 B.n264 VSUBS 0.010591f
C305 B.n265 VSUBS 0.010591f
C306 B.n266 VSUBS 0.010591f
C307 B.n267 VSUBS 0.010591f
C308 B.n268 VSUBS 0.010591f
C309 B.n269 VSUBS 0.010591f
C310 B.n270 VSUBS 0.010591f
C311 B.n271 VSUBS 0.010591f
C312 B.n272 VSUBS 0.010591f
C313 B.n273 VSUBS 0.010591f
C314 B.n274 VSUBS 0.010591f
C315 B.n275 VSUBS 0.010591f
C316 B.n276 VSUBS 0.010591f
C317 B.n277 VSUBS 0.010591f
C318 B.n278 VSUBS 0.010591f
C319 B.n279 VSUBS 0.010591f
C320 B.n280 VSUBS 0.010591f
C321 B.n281 VSUBS 0.010591f
C322 B.n282 VSUBS 0.010591f
C323 B.n283 VSUBS 0.026585f
C324 B.n284 VSUBS 0.025411f
C325 B.n285 VSUBS 0.026299f
C326 B.n286 VSUBS 0.010591f
C327 B.n287 VSUBS 0.010591f
C328 B.n288 VSUBS 0.010591f
C329 B.n289 VSUBS 0.010591f
C330 B.n290 VSUBS 0.010591f
C331 B.n291 VSUBS 0.010591f
C332 B.n292 VSUBS 0.010591f
C333 B.n293 VSUBS 0.010591f
C334 B.n294 VSUBS 0.010591f
C335 B.n295 VSUBS 0.010591f
C336 B.n296 VSUBS 0.010591f
C337 B.n297 VSUBS 0.010591f
C338 B.n298 VSUBS 0.010591f
C339 B.n299 VSUBS 0.010591f
C340 B.n300 VSUBS 0.010591f
C341 B.n301 VSUBS 0.010591f
C342 B.n302 VSUBS 0.010591f
C343 B.n303 VSUBS 0.010591f
C344 B.n304 VSUBS 0.010591f
C345 B.n305 VSUBS 0.010591f
C346 B.n306 VSUBS 0.010591f
C347 B.n307 VSUBS 0.010591f
C348 B.n308 VSUBS 0.010591f
C349 B.n309 VSUBS 0.010591f
C350 B.n310 VSUBS 0.010591f
C351 B.n311 VSUBS 0.010591f
C352 B.n312 VSUBS 0.010591f
C353 B.n313 VSUBS 0.010591f
C354 B.n314 VSUBS 0.010591f
C355 B.n315 VSUBS 0.010591f
C356 B.n316 VSUBS 0.010591f
C357 B.n317 VSUBS 0.010591f
C358 B.n318 VSUBS 0.010591f
C359 B.n319 VSUBS 0.010591f
C360 B.n320 VSUBS 0.010591f
C361 B.n321 VSUBS 0.010591f
C362 B.n322 VSUBS 0.010591f
C363 B.n323 VSUBS 0.010591f
C364 B.n324 VSUBS 0.010591f
C365 B.n325 VSUBS 0.010591f
C366 B.n326 VSUBS 0.010591f
C367 B.n327 VSUBS 0.010591f
C368 B.n328 VSUBS 0.010591f
C369 B.n329 VSUBS 0.010591f
C370 B.n330 VSUBS 0.010591f
C371 B.n331 VSUBS 0.010591f
C372 B.n332 VSUBS 0.010591f
C373 B.n333 VSUBS 0.010591f
C374 B.n334 VSUBS 0.010591f
C375 B.n335 VSUBS 0.010591f
C376 B.n336 VSUBS 0.010591f
C377 B.n337 VSUBS 0.010591f
C378 B.n338 VSUBS 0.010591f
C379 B.n339 VSUBS 0.010591f
C380 B.n340 VSUBS 0.010591f
C381 B.n341 VSUBS 0.010591f
C382 B.n342 VSUBS 0.010591f
C383 B.n343 VSUBS 0.010591f
C384 B.n344 VSUBS 0.010591f
C385 B.n345 VSUBS 0.010591f
C386 B.n346 VSUBS 0.010591f
C387 B.n347 VSUBS 0.010591f
C388 B.n348 VSUBS 0.010591f
C389 B.n349 VSUBS 0.010591f
C390 B.n350 VSUBS 0.010591f
C391 B.n351 VSUBS 0.010591f
C392 B.n352 VSUBS 0.010591f
C393 B.n353 VSUBS 0.010591f
C394 B.n354 VSUBS 0.010591f
C395 B.n355 VSUBS 0.010591f
C396 B.n356 VSUBS 0.010591f
C397 B.n357 VSUBS 0.010591f
C398 B.n358 VSUBS 0.010591f
C399 B.n359 VSUBS 0.010591f
C400 B.n360 VSUBS 0.010591f
C401 B.n361 VSUBS 0.010591f
C402 B.n362 VSUBS 0.010591f
C403 B.n363 VSUBS 0.010591f
C404 B.n364 VSUBS 0.010591f
C405 B.n365 VSUBS 0.010591f
C406 B.n366 VSUBS 0.010591f
C407 B.n367 VSUBS 0.010591f
C408 B.n368 VSUBS 0.010591f
C409 B.n369 VSUBS 0.010591f
C410 B.n370 VSUBS 0.010591f
C411 B.n371 VSUBS 0.010591f
C412 B.n372 VSUBS 0.010591f
C413 B.n373 VSUBS 0.010591f
C414 B.n374 VSUBS 0.010591f
C415 B.n375 VSUBS 0.010591f
C416 B.n376 VSUBS 0.010591f
C417 B.n377 VSUBS 0.010591f
C418 B.n378 VSUBS 0.010591f
C419 B.n379 VSUBS 0.010591f
C420 B.n380 VSUBS 0.010591f
C421 B.n381 VSUBS 0.010591f
C422 B.n382 VSUBS 0.010591f
C423 B.n383 VSUBS 0.010591f
C424 B.n384 VSUBS 0.010591f
C425 B.n385 VSUBS 0.010591f
C426 B.n386 VSUBS 0.010591f
C427 B.n387 VSUBS 0.010591f
C428 B.n388 VSUBS 0.010591f
C429 B.n389 VSUBS 0.010591f
C430 B.n390 VSUBS 0.010591f
C431 B.n391 VSUBS 0.010591f
C432 B.n392 VSUBS 0.010591f
C433 B.n393 VSUBS 0.010591f
C434 B.n394 VSUBS 0.010591f
C435 B.n395 VSUBS 0.010591f
C436 B.n396 VSUBS 0.010591f
C437 B.n397 VSUBS 0.010591f
C438 B.n398 VSUBS 0.010591f
C439 B.n399 VSUBS 0.010591f
C440 B.n400 VSUBS 0.010591f
C441 B.n401 VSUBS 0.010591f
C442 B.n402 VSUBS 0.010591f
C443 B.n403 VSUBS 0.010591f
C444 B.n404 VSUBS 0.010591f
C445 B.n405 VSUBS 0.010591f
C446 B.n406 VSUBS 0.010591f
C447 B.n407 VSUBS 0.010591f
C448 B.n408 VSUBS 0.010591f
C449 B.n409 VSUBS 0.010591f
C450 B.n410 VSUBS 0.010591f
C451 B.n411 VSUBS 0.010591f
C452 B.n412 VSUBS 0.010591f
C453 B.n413 VSUBS 0.010591f
C454 B.n414 VSUBS 0.010591f
C455 B.n415 VSUBS 0.010591f
C456 B.n416 VSUBS 0.010591f
C457 B.n417 VSUBS 0.010591f
C458 B.n418 VSUBS 0.010591f
C459 B.n419 VSUBS 0.010591f
C460 B.n420 VSUBS 0.010591f
C461 B.n421 VSUBS 0.025125f
C462 B.n422 VSUBS 0.025125f
C463 B.n423 VSUBS 0.026585f
C464 B.n424 VSUBS 0.010591f
C465 B.n425 VSUBS 0.010591f
C466 B.n426 VSUBS 0.010591f
C467 B.n427 VSUBS 0.010591f
C468 B.n428 VSUBS 0.010591f
C469 B.n429 VSUBS 0.010591f
C470 B.n430 VSUBS 0.010591f
C471 B.n431 VSUBS 0.010591f
C472 B.n432 VSUBS 0.010591f
C473 B.n433 VSUBS 0.010591f
C474 B.n434 VSUBS 0.010591f
C475 B.n435 VSUBS 0.010591f
C476 B.n436 VSUBS 0.010591f
C477 B.n437 VSUBS 0.010591f
C478 B.n438 VSUBS 0.010591f
C479 B.n439 VSUBS 0.010591f
C480 B.n440 VSUBS 0.010591f
C481 B.n441 VSUBS 0.010591f
C482 B.n442 VSUBS 0.010591f
C483 B.n443 VSUBS 0.010591f
C484 B.n444 VSUBS 0.010591f
C485 B.n445 VSUBS 0.010591f
C486 B.n446 VSUBS 0.010591f
C487 B.n447 VSUBS 0.010591f
C488 B.n448 VSUBS 0.009968f
C489 B.n449 VSUBS 0.010591f
C490 B.n450 VSUBS 0.010591f
C491 B.n451 VSUBS 0.010591f
C492 B.n452 VSUBS 0.010591f
C493 B.n453 VSUBS 0.010591f
C494 B.n454 VSUBS 0.010591f
C495 B.n455 VSUBS 0.010591f
C496 B.n456 VSUBS 0.010591f
C497 B.n457 VSUBS 0.010591f
C498 B.n458 VSUBS 0.010591f
C499 B.n459 VSUBS 0.010591f
C500 B.n460 VSUBS 0.010591f
C501 B.n461 VSUBS 0.010591f
C502 B.n462 VSUBS 0.010591f
C503 B.n463 VSUBS 0.010591f
C504 B.n464 VSUBS 0.005919f
C505 B.n465 VSUBS 0.024539f
C506 B.n466 VSUBS 0.009968f
C507 B.n467 VSUBS 0.010591f
C508 B.n468 VSUBS 0.010591f
C509 B.n469 VSUBS 0.010591f
C510 B.n470 VSUBS 0.010591f
C511 B.n471 VSUBS 0.010591f
C512 B.n472 VSUBS 0.010591f
C513 B.n473 VSUBS 0.010591f
C514 B.n474 VSUBS 0.010591f
C515 B.n475 VSUBS 0.010591f
C516 B.n476 VSUBS 0.010591f
C517 B.n477 VSUBS 0.010591f
C518 B.n478 VSUBS 0.010591f
C519 B.n479 VSUBS 0.010591f
C520 B.n480 VSUBS 0.010591f
C521 B.n481 VSUBS 0.010591f
C522 B.n482 VSUBS 0.010591f
C523 B.n483 VSUBS 0.010591f
C524 B.n484 VSUBS 0.010591f
C525 B.n485 VSUBS 0.010591f
C526 B.n486 VSUBS 0.010591f
C527 B.n487 VSUBS 0.010591f
C528 B.n488 VSUBS 0.010591f
C529 B.n489 VSUBS 0.010591f
C530 B.n490 VSUBS 0.010591f
C531 B.n491 VSUBS 0.026585f
C532 B.n492 VSUBS 0.026585f
C533 B.n493 VSUBS 0.025125f
C534 B.n494 VSUBS 0.010591f
C535 B.n495 VSUBS 0.010591f
C536 B.n496 VSUBS 0.010591f
C537 B.n497 VSUBS 0.010591f
C538 B.n498 VSUBS 0.010591f
C539 B.n499 VSUBS 0.010591f
C540 B.n500 VSUBS 0.010591f
C541 B.n501 VSUBS 0.010591f
C542 B.n502 VSUBS 0.010591f
C543 B.n503 VSUBS 0.010591f
C544 B.n504 VSUBS 0.010591f
C545 B.n505 VSUBS 0.010591f
C546 B.n506 VSUBS 0.010591f
C547 B.n507 VSUBS 0.010591f
C548 B.n508 VSUBS 0.010591f
C549 B.n509 VSUBS 0.010591f
C550 B.n510 VSUBS 0.010591f
C551 B.n511 VSUBS 0.010591f
C552 B.n512 VSUBS 0.010591f
C553 B.n513 VSUBS 0.010591f
C554 B.n514 VSUBS 0.010591f
C555 B.n515 VSUBS 0.010591f
C556 B.n516 VSUBS 0.010591f
C557 B.n517 VSUBS 0.010591f
C558 B.n518 VSUBS 0.010591f
C559 B.n519 VSUBS 0.010591f
C560 B.n520 VSUBS 0.010591f
C561 B.n521 VSUBS 0.010591f
C562 B.n522 VSUBS 0.010591f
C563 B.n523 VSUBS 0.010591f
C564 B.n524 VSUBS 0.010591f
C565 B.n525 VSUBS 0.010591f
C566 B.n526 VSUBS 0.010591f
C567 B.n527 VSUBS 0.010591f
C568 B.n528 VSUBS 0.010591f
C569 B.n529 VSUBS 0.010591f
C570 B.n530 VSUBS 0.010591f
C571 B.n531 VSUBS 0.010591f
C572 B.n532 VSUBS 0.010591f
C573 B.n533 VSUBS 0.010591f
C574 B.n534 VSUBS 0.010591f
C575 B.n535 VSUBS 0.010591f
C576 B.n536 VSUBS 0.010591f
C577 B.n537 VSUBS 0.010591f
C578 B.n538 VSUBS 0.010591f
C579 B.n539 VSUBS 0.010591f
C580 B.n540 VSUBS 0.010591f
C581 B.n541 VSUBS 0.010591f
C582 B.n542 VSUBS 0.010591f
C583 B.n543 VSUBS 0.010591f
C584 B.n544 VSUBS 0.010591f
C585 B.n545 VSUBS 0.010591f
C586 B.n546 VSUBS 0.010591f
C587 B.n547 VSUBS 0.010591f
C588 B.n548 VSUBS 0.010591f
C589 B.n549 VSUBS 0.010591f
C590 B.n550 VSUBS 0.010591f
C591 B.n551 VSUBS 0.010591f
C592 B.n552 VSUBS 0.010591f
C593 B.n553 VSUBS 0.010591f
C594 B.n554 VSUBS 0.010591f
C595 B.n555 VSUBS 0.010591f
C596 B.n556 VSUBS 0.010591f
C597 B.n557 VSUBS 0.010591f
C598 B.n558 VSUBS 0.010591f
C599 B.n559 VSUBS 0.013821f
C600 B.n560 VSUBS 0.014723f
C601 B.n561 VSUBS 0.029278f
C602 VDD2.t2 VSUBS 0.063972f
C603 VDD2.t0 VSUBS 0.063972f
C604 VDD2.n0 VSUBS 0.63012f
C605 VDD2.t3 VSUBS 0.063972f
C606 VDD2.t1 VSUBS 0.063972f
C607 VDD2.n1 VSUBS 0.375587f
C608 VDD2.n2 VSUBS 2.69757f
C609 VN.t1 VSUBS 1.94959f
C610 VN.t3 VSUBS 1.92836f
C611 VN.n0 VSUBS 1.19901f
C612 VN.t2 VSUBS 1.94959f
C613 VN.t0 VSUBS 1.92836f
C614 VN.n1 VSUBS 3.22629f
C615 VDD1.t0 VSUBS 0.097294f
C616 VDD1.t2 VSUBS 0.097294f
C617 VDD1.n0 VSUBS 0.571625f
C618 VDD1.t1 VSUBS 0.097294f
C619 VDD1.t3 VSUBS 0.097294f
C620 VDD1.n1 VSUBS 0.97736f
C621 VTAIL.n0 VSUBS 0.036943f
C622 VTAIL.n1 VSUBS 0.032613f
C623 VTAIL.n2 VSUBS 0.017525f
C624 VTAIL.n3 VSUBS 0.041423f
C625 VTAIL.n4 VSUBS 0.018556f
C626 VTAIL.n5 VSUBS 0.128311f
C627 VTAIL.t3 VSUBS 0.092517f
C628 VTAIL.n6 VSUBS 0.031067f
C629 VTAIL.n7 VSUBS 0.026054f
C630 VTAIL.n8 VSUBS 0.017525f
C631 VTAIL.n9 VSUBS 0.453035f
C632 VTAIL.n10 VSUBS 0.032613f
C633 VTAIL.n11 VSUBS 0.017525f
C634 VTAIL.n12 VSUBS 0.018556f
C635 VTAIL.n13 VSUBS 0.041423f
C636 VTAIL.n14 VSUBS 0.104053f
C637 VTAIL.n15 VSUBS 0.018556f
C638 VTAIL.n16 VSUBS 0.017525f
C639 VTAIL.n17 VSUBS 0.08474f
C640 VTAIL.n18 VSUBS 0.052768f
C641 VTAIL.n19 VSUBS 0.281598f
C642 VTAIL.n20 VSUBS 0.036943f
C643 VTAIL.n21 VSUBS 0.032613f
C644 VTAIL.n22 VSUBS 0.017525f
C645 VTAIL.n23 VSUBS 0.041423f
C646 VTAIL.n24 VSUBS 0.018556f
C647 VTAIL.n25 VSUBS 0.128311f
C648 VTAIL.t4 VSUBS 0.092517f
C649 VTAIL.n26 VSUBS 0.031067f
C650 VTAIL.n27 VSUBS 0.026054f
C651 VTAIL.n28 VSUBS 0.017525f
C652 VTAIL.n29 VSUBS 0.453035f
C653 VTAIL.n30 VSUBS 0.032613f
C654 VTAIL.n31 VSUBS 0.017525f
C655 VTAIL.n32 VSUBS 0.018556f
C656 VTAIL.n33 VSUBS 0.041423f
C657 VTAIL.n34 VSUBS 0.104053f
C658 VTAIL.n35 VSUBS 0.018556f
C659 VTAIL.n36 VSUBS 0.017525f
C660 VTAIL.n37 VSUBS 0.08474f
C661 VTAIL.n38 VSUBS 0.052768f
C662 VTAIL.n39 VSUBS 0.468445f
C663 VTAIL.n40 VSUBS 0.036943f
C664 VTAIL.n41 VSUBS 0.032613f
C665 VTAIL.n42 VSUBS 0.017525f
C666 VTAIL.n43 VSUBS 0.041423f
C667 VTAIL.n44 VSUBS 0.018556f
C668 VTAIL.n45 VSUBS 0.128311f
C669 VTAIL.t6 VSUBS 0.092517f
C670 VTAIL.n46 VSUBS 0.031067f
C671 VTAIL.n47 VSUBS 0.026054f
C672 VTAIL.n48 VSUBS 0.017525f
C673 VTAIL.n49 VSUBS 0.453035f
C674 VTAIL.n50 VSUBS 0.032613f
C675 VTAIL.n51 VSUBS 0.017525f
C676 VTAIL.n52 VSUBS 0.018556f
C677 VTAIL.n53 VSUBS 0.041423f
C678 VTAIL.n54 VSUBS 0.104053f
C679 VTAIL.n55 VSUBS 0.018556f
C680 VTAIL.n56 VSUBS 0.017525f
C681 VTAIL.n57 VSUBS 0.08474f
C682 VTAIL.n58 VSUBS 0.052768f
C683 VTAIL.n59 VSUBS 1.6149f
C684 VTAIL.n60 VSUBS 0.036943f
C685 VTAIL.n61 VSUBS 0.032613f
C686 VTAIL.n62 VSUBS 0.017525f
C687 VTAIL.n63 VSUBS 0.041423f
C688 VTAIL.n64 VSUBS 0.018556f
C689 VTAIL.n65 VSUBS 0.128311f
C690 VTAIL.t2 VSUBS 0.092517f
C691 VTAIL.n66 VSUBS 0.031067f
C692 VTAIL.n67 VSUBS 0.026054f
C693 VTAIL.n68 VSUBS 0.017525f
C694 VTAIL.n69 VSUBS 0.453035f
C695 VTAIL.n70 VSUBS 0.032613f
C696 VTAIL.n71 VSUBS 0.017525f
C697 VTAIL.n72 VSUBS 0.018556f
C698 VTAIL.n73 VSUBS 0.041423f
C699 VTAIL.n74 VSUBS 0.104053f
C700 VTAIL.n75 VSUBS 0.018556f
C701 VTAIL.n76 VSUBS 0.017525f
C702 VTAIL.n77 VSUBS 0.08474f
C703 VTAIL.n78 VSUBS 0.052768f
C704 VTAIL.n79 VSUBS 1.6149f
C705 VTAIL.n80 VSUBS 0.036943f
C706 VTAIL.n81 VSUBS 0.032613f
C707 VTAIL.n82 VSUBS 0.017525f
C708 VTAIL.n83 VSUBS 0.041423f
C709 VTAIL.n84 VSUBS 0.018556f
C710 VTAIL.n85 VSUBS 0.128311f
C711 VTAIL.t1 VSUBS 0.092517f
C712 VTAIL.n86 VSUBS 0.031067f
C713 VTAIL.n87 VSUBS 0.026054f
C714 VTAIL.n88 VSUBS 0.017525f
C715 VTAIL.n89 VSUBS 0.453035f
C716 VTAIL.n90 VSUBS 0.032613f
C717 VTAIL.n91 VSUBS 0.017525f
C718 VTAIL.n92 VSUBS 0.018556f
C719 VTAIL.n93 VSUBS 0.041423f
C720 VTAIL.n94 VSUBS 0.104053f
C721 VTAIL.n95 VSUBS 0.018556f
C722 VTAIL.n96 VSUBS 0.017525f
C723 VTAIL.n97 VSUBS 0.08474f
C724 VTAIL.n98 VSUBS 0.052768f
C725 VTAIL.n99 VSUBS 0.468445f
C726 VTAIL.n100 VSUBS 0.036943f
C727 VTAIL.n101 VSUBS 0.032613f
C728 VTAIL.n102 VSUBS 0.017525f
C729 VTAIL.n103 VSUBS 0.041423f
C730 VTAIL.n104 VSUBS 0.018556f
C731 VTAIL.n105 VSUBS 0.128311f
C732 VTAIL.t7 VSUBS 0.092517f
C733 VTAIL.n106 VSUBS 0.031067f
C734 VTAIL.n107 VSUBS 0.026054f
C735 VTAIL.n108 VSUBS 0.017525f
C736 VTAIL.n109 VSUBS 0.453035f
C737 VTAIL.n110 VSUBS 0.032613f
C738 VTAIL.n111 VSUBS 0.017525f
C739 VTAIL.n112 VSUBS 0.018556f
C740 VTAIL.n113 VSUBS 0.041423f
C741 VTAIL.n114 VSUBS 0.104053f
C742 VTAIL.n115 VSUBS 0.018556f
C743 VTAIL.n116 VSUBS 0.017525f
C744 VTAIL.n117 VSUBS 0.08474f
C745 VTAIL.n118 VSUBS 0.052768f
C746 VTAIL.n119 VSUBS 0.468445f
C747 VTAIL.n120 VSUBS 0.036943f
C748 VTAIL.n121 VSUBS 0.032613f
C749 VTAIL.n122 VSUBS 0.017525f
C750 VTAIL.n123 VSUBS 0.041423f
C751 VTAIL.n124 VSUBS 0.018556f
C752 VTAIL.n125 VSUBS 0.128311f
C753 VTAIL.t5 VSUBS 0.092517f
C754 VTAIL.n126 VSUBS 0.031067f
C755 VTAIL.n127 VSUBS 0.026054f
C756 VTAIL.n128 VSUBS 0.017525f
C757 VTAIL.n129 VSUBS 0.453035f
C758 VTAIL.n130 VSUBS 0.032613f
C759 VTAIL.n131 VSUBS 0.017525f
C760 VTAIL.n132 VSUBS 0.018556f
C761 VTAIL.n133 VSUBS 0.041423f
C762 VTAIL.n134 VSUBS 0.104053f
C763 VTAIL.n135 VSUBS 0.018556f
C764 VTAIL.n136 VSUBS 0.017525f
C765 VTAIL.n137 VSUBS 0.08474f
C766 VTAIL.n138 VSUBS 0.052768f
C767 VTAIL.n139 VSUBS 1.6149f
C768 VTAIL.n140 VSUBS 0.036943f
C769 VTAIL.n141 VSUBS 0.032613f
C770 VTAIL.n142 VSUBS 0.017525f
C771 VTAIL.n143 VSUBS 0.041423f
C772 VTAIL.n144 VSUBS 0.018556f
C773 VTAIL.n145 VSUBS 0.128311f
C774 VTAIL.t0 VSUBS 0.092517f
C775 VTAIL.n146 VSUBS 0.031067f
C776 VTAIL.n147 VSUBS 0.026054f
C777 VTAIL.n148 VSUBS 0.017525f
C778 VTAIL.n149 VSUBS 0.453035f
C779 VTAIL.n150 VSUBS 0.032613f
C780 VTAIL.n151 VSUBS 0.017525f
C781 VTAIL.n152 VSUBS 0.018556f
C782 VTAIL.n153 VSUBS 0.041423f
C783 VTAIL.n154 VSUBS 0.104053f
C784 VTAIL.n155 VSUBS 0.018556f
C785 VTAIL.n156 VSUBS 0.017525f
C786 VTAIL.n157 VSUBS 0.08474f
C787 VTAIL.n158 VSUBS 0.052768f
C788 VTAIL.n159 VSUBS 1.41583f
C789 VP.n0 VSUBS 0.089081f
C790 VP.t0 VSUBS 1.93858f
C791 VP.n1 VSUBS 0.088264f
C792 VP.n2 VSUBS 0.047358f
C793 VP.n3 VSUBS 0.088264f
C794 VP.t1 VSUBS 2.56667f
C795 VP.t3 VSUBS 2.59492f
C796 VP.n4 VSUBS 4.28108f
C797 VP.n5 VSUBS 2.48498f
C798 VP.t2 VSUBS 1.93858f
C799 VP.n6 VSUBS 0.948465f
C800 VP.n7 VSUBS 0.077806f
C801 VP.n8 VSUBS 0.089081f
C802 VP.n9 VSUBS 0.047358f
C803 VP.n10 VSUBS 0.047358f
C804 VP.n11 VSUBS 0.088264f
C805 VP.n12 VSUBS 0.069135f
C806 VP.n13 VSUBS 0.069135f
C807 VP.n14 VSUBS 0.047358f
C808 VP.n15 VSUBS 0.047358f
C809 VP.n16 VSUBS 0.047358f
C810 VP.n17 VSUBS 0.088264f
C811 VP.n18 VSUBS 0.077806f
C812 VP.n19 VSUBS 0.948465f
C813 VP.n20 VSUBS 0.154089f
.ends

