* NGSPICE file created from diff_pair_sample_0765.ext - technology: sky130A

.subckt diff_pair_sample_0765 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t10 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=1.08
X1 B.t15 B.t13 B.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=1.08
X2 VDD1.t5 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=6.0528 ps=31.82 w=15.52 l=1.08
X3 VDD2.t5 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=6.0528 ps=31.82 w=15.52 l=1.08
X4 VDD2.t4 VN.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=2.5608 ps=15.85 w=15.52 l=1.08
X5 VDD1.t4 VP.t1 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=2.5608 ps=15.85 w=15.52 l=1.08
X6 VDD2.t3 VN.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=2.5608 ps=15.85 w=15.52 l=1.08
X7 VTAIL.t11 VN.t3 VDD2.t2 B.t19 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=2.5608 ps=15.85 w=15.52 l=1.08
X8 VDD1.t3 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=6.0528 ps=31.82 w=15.52 l=1.08
X9 VDD2.t1 VN.t4 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=6.0528 ps=31.82 w=15.52 l=1.08
X10 VTAIL.t4 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=2.5608 ps=15.85 w=15.52 l=1.08
X11 VDD1.t1 VP.t4 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=2.5608 ps=15.85 w=15.52 l=1.08
X12 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=1.08
X13 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=1.08
X14 VTAIL.t6 VP.t5 VDD1.t0 B.t19 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=2.5608 ps=15.85 w=15.52 l=1.08
X15 VTAIL.t2 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5608 pd=15.85 as=2.5608 ps=15.85 w=15.52 l=1.08
R0 B.n777 B.n776 585
R1 B.n333 B.n104 585
R2 B.n332 B.n331 585
R3 B.n330 B.n329 585
R4 B.n328 B.n327 585
R5 B.n326 B.n325 585
R6 B.n324 B.n323 585
R7 B.n322 B.n321 585
R8 B.n320 B.n319 585
R9 B.n318 B.n317 585
R10 B.n316 B.n315 585
R11 B.n314 B.n313 585
R12 B.n312 B.n311 585
R13 B.n310 B.n309 585
R14 B.n308 B.n307 585
R15 B.n306 B.n305 585
R16 B.n304 B.n303 585
R17 B.n302 B.n301 585
R18 B.n300 B.n299 585
R19 B.n298 B.n297 585
R20 B.n296 B.n295 585
R21 B.n294 B.n293 585
R22 B.n292 B.n291 585
R23 B.n290 B.n289 585
R24 B.n288 B.n287 585
R25 B.n286 B.n285 585
R26 B.n284 B.n283 585
R27 B.n282 B.n281 585
R28 B.n280 B.n279 585
R29 B.n278 B.n277 585
R30 B.n276 B.n275 585
R31 B.n274 B.n273 585
R32 B.n272 B.n271 585
R33 B.n270 B.n269 585
R34 B.n268 B.n267 585
R35 B.n266 B.n265 585
R36 B.n264 B.n263 585
R37 B.n262 B.n261 585
R38 B.n260 B.n259 585
R39 B.n258 B.n257 585
R40 B.n256 B.n255 585
R41 B.n254 B.n253 585
R42 B.n252 B.n251 585
R43 B.n250 B.n249 585
R44 B.n248 B.n247 585
R45 B.n246 B.n245 585
R46 B.n244 B.n243 585
R47 B.n242 B.n241 585
R48 B.n240 B.n239 585
R49 B.n238 B.n237 585
R50 B.n236 B.n235 585
R51 B.n234 B.n233 585
R52 B.n232 B.n231 585
R53 B.n230 B.n229 585
R54 B.n228 B.n227 585
R55 B.n226 B.n225 585
R56 B.n224 B.n223 585
R57 B.n222 B.n221 585
R58 B.n220 B.n219 585
R59 B.n218 B.n217 585
R60 B.n216 B.n215 585
R61 B.n214 B.n213 585
R62 B.n212 B.n211 585
R63 B.n210 B.n209 585
R64 B.n208 B.n207 585
R65 B.n206 B.n205 585
R66 B.n204 B.n203 585
R67 B.n202 B.n201 585
R68 B.n200 B.n199 585
R69 B.n198 B.n197 585
R70 B.n196 B.n195 585
R71 B.n194 B.n193 585
R72 B.n192 B.n191 585
R73 B.n190 B.n189 585
R74 B.n188 B.n187 585
R75 B.n186 B.n185 585
R76 B.n184 B.n183 585
R77 B.n182 B.n181 585
R78 B.n180 B.n179 585
R79 B.n178 B.n177 585
R80 B.n176 B.n175 585
R81 B.n174 B.n173 585
R82 B.n172 B.n171 585
R83 B.n170 B.n169 585
R84 B.n168 B.n167 585
R85 B.n166 B.n165 585
R86 B.n164 B.n163 585
R87 B.n162 B.n161 585
R88 B.n160 B.n159 585
R89 B.n158 B.n157 585
R90 B.n156 B.n155 585
R91 B.n154 B.n153 585
R92 B.n152 B.n151 585
R93 B.n150 B.n149 585
R94 B.n148 B.n147 585
R95 B.n146 B.n145 585
R96 B.n144 B.n143 585
R97 B.n142 B.n141 585
R98 B.n140 B.n139 585
R99 B.n138 B.n137 585
R100 B.n136 B.n135 585
R101 B.n134 B.n133 585
R102 B.n132 B.n131 585
R103 B.n130 B.n129 585
R104 B.n128 B.n127 585
R105 B.n126 B.n125 585
R106 B.n124 B.n123 585
R107 B.n122 B.n121 585
R108 B.n120 B.n119 585
R109 B.n118 B.n117 585
R110 B.n116 B.n115 585
R111 B.n114 B.n113 585
R112 B.n112 B.n111 585
R113 B.n46 B.n45 585
R114 B.n775 B.n47 585
R115 B.n780 B.n47 585
R116 B.n774 B.n773 585
R117 B.n773 B.n43 585
R118 B.n772 B.n42 585
R119 B.n786 B.n42 585
R120 B.n771 B.n41 585
R121 B.n787 B.n41 585
R122 B.n770 B.n40 585
R123 B.n788 B.n40 585
R124 B.n769 B.n768 585
R125 B.n768 B.n39 585
R126 B.n767 B.n35 585
R127 B.n794 B.n35 585
R128 B.n766 B.n34 585
R129 B.n795 B.n34 585
R130 B.n765 B.n33 585
R131 B.n796 B.n33 585
R132 B.n764 B.n763 585
R133 B.n763 B.n29 585
R134 B.n762 B.n28 585
R135 B.n802 B.n28 585
R136 B.n761 B.n27 585
R137 B.n803 B.n27 585
R138 B.n760 B.n26 585
R139 B.n804 B.n26 585
R140 B.n759 B.n758 585
R141 B.n758 B.n22 585
R142 B.n757 B.n21 585
R143 B.n810 B.n21 585
R144 B.n756 B.n20 585
R145 B.n811 B.n20 585
R146 B.n755 B.n19 585
R147 B.n812 B.n19 585
R148 B.n754 B.n753 585
R149 B.n753 B.n15 585
R150 B.n752 B.n14 585
R151 B.n818 B.n14 585
R152 B.n751 B.n13 585
R153 B.n819 B.n13 585
R154 B.n750 B.n12 585
R155 B.n820 B.n12 585
R156 B.n749 B.n748 585
R157 B.n748 B.n747 585
R158 B.n746 B.n745 585
R159 B.n746 B.n8 585
R160 B.n744 B.n7 585
R161 B.n827 B.n7 585
R162 B.n743 B.n6 585
R163 B.n828 B.n6 585
R164 B.n742 B.n5 585
R165 B.n829 B.n5 585
R166 B.n741 B.n740 585
R167 B.n740 B.n4 585
R168 B.n739 B.n334 585
R169 B.n739 B.n738 585
R170 B.n729 B.n335 585
R171 B.n336 B.n335 585
R172 B.n731 B.n730 585
R173 B.n732 B.n731 585
R174 B.n728 B.n341 585
R175 B.n341 B.n340 585
R176 B.n727 B.n726 585
R177 B.n726 B.n725 585
R178 B.n343 B.n342 585
R179 B.n344 B.n343 585
R180 B.n718 B.n717 585
R181 B.n719 B.n718 585
R182 B.n716 B.n349 585
R183 B.n349 B.n348 585
R184 B.n715 B.n714 585
R185 B.n714 B.n713 585
R186 B.n351 B.n350 585
R187 B.n352 B.n351 585
R188 B.n706 B.n705 585
R189 B.n707 B.n706 585
R190 B.n704 B.n357 585
R191 B.n357 B.n356 585
R192 B.n703 B.n702 585
R193 B.n702 B.n701 585
R194 B.n359 B.n358 585
R195 B.n360 B.n359 585
R196 B.n694 B.n693 585
R197 B.n695 B.n694 585
R198 B.n692 B.n365 585
R199 B.n365 B.n364 585
R200 B.n691 B.n690 585
R201 B.n690 B.n689 585
R202 B.n367 B.n366 585
R203 B.n682 B.n367 585
R204 B.n681 B.n680 585
R205 B.n683 B.n681 585
R206 B.n679 B.n372 585
R207 B.n372 B.n371 585
R208 B.n678 B.n677 585
R209 B.n677 B.n676 585
R210 B.n374 B.n373 585
R211 B.n375 B.n374 585
R212 B.n669 B.n668 585
R213 B.n670 B.n669 585
R214 B.n378 B.n377 585
R215 B.n441 B.n439 585
R216 B.n442 B.n438 585
R217 B.n442 B.n379 585
R218 B.n445 B.n444 585
R219 B.n446 B.n437 585
R220 B.n448 B.n447 585
R221 B.n450 B.n436 585
R222 B.n453 B.n452 585
R223 B.n454 B.n435 585
R224 B.n456 B.n455 585
R225 B.n458 B.n434 585
R226 B.n461 B.n460 585
R227 B.n462 B.n433 585
R228 B.n464 B.n463 585
R229 B.n466 B.n432 585
R230 B.n469 B.n468 585
R231 B.n470 B.n431 585
R232 B.n472 B.n471 585
R233 B.n474 B.n430 585
R234 B.n477 B.n476 585
R235 B.n478 B.n429 585
R236 B.n480 B.n479 585
R237 B.n482 B.n428 585
R238 B.n485 B.n484 585
R239 B.n486 B.n427 585
R240 B.n488 B.n487 585
R241 B.n490 B.n426 585
R242 B.n493 B.n492 585
R243 B.n494 B.n425 585
R244 B.n496 B.n495 585
R245 B.n498 B.n424 585
R246 B.n501 B.n500 585
R247 B.n502 B.n423 585
R248 B.n504 B.n503 585
R249 B.n506 B.n422 585
R250 B.n509 B.n508 585
R251 B.n510 B.n421 585
R252 B.n512 B.n511 585
R253 B.n514 B.n420 585
R254 B.n517 B.n516 585
R255 B.n518 B.n419 585
R256 B.n520 B.n519 585
R257 B.n522 B.n418 585
R258 B.n525 B.n524 585
R259 B.n526 B.n417 585
R260 B.n528 B.n527 585
R261 B.n530 B.n416 585
R262 B.n533 B.n532 585
R263 B.n534 B.n415 585
R264 B.n536 B.n535 585
R265 B.n538 B.n414 585
R266 B.n541 B.n540 585
R267 B.n543 B.n411 585
R268 B.n545 B.n544 585
R269 B.n547 B.n410 585
R270 B.n550 B.n549 585
R271 B.n551 B.n409 585
R272 B.n553 B.n552 585
R273 B.n555 B.n408 585
R274 B.n558 B.n557 585
R275 B.n559 B.n407 585
R276 B.n564 B.n563 585
R277 B.n566 B.n406 585
R278 B.n569 B.n568 585
R279 B.n570 B.n405 585
R280 B.n572 B.n571 585
R281 B.n574 B.n404 585
R282 B.n577 B.n576 585
R283 B.n578 B.n403 585
R284 B.n580 B.n579 585
R285 B.n582 B.n402 585
R286 B.n585 B.n584 585
R287 B.n586 B.n401 585
R288 B.n588 B.n587 585
R289 B.n590 B.n400 585
R290 B.n593 B.n592 585
R291 B.n594 B.n399 585
R292 B.n596 B.n595 585
R293 B.n598 B.n398 585
R294 B.n601 B.n600 585
R295 B.n602 B.n397 585
R296 B.n604 B.n603 585
R297 B.n606 B.n396 585
R298 B.n609 B.n608 585
R299 B.n610 B.n395 585
R300 B.n612 B.n611 585
R301 B.n614 B.n394 585
R302 B.n617 B.n616 585
R303 B.n618 B.n393 585
R304 B.n620 B.n619 585
R305 B.n622 B.n392 585
R306 B.n625 B.n624 585
R307 B.n626 B.n391 585
R308 B.n628 B.n627 585
R309 B.n630 B.n390 585
R310 B.n633 B.n632 585
R311 B.n634 B.n389 585
R312 B.n636 B.n635 585
R313 B.n638 B.n388 585
R314 B.n641 B.n640 585
R315 B.n642 B.n387 585
R316 B.n644 B.n643 585
R317 B.n646 B.n386 585
R318 B.n649 B.n648 585
R319 B.n650 B.n385 585
R320 B.n652 B.n651 585
R321 B.n654 B.n384 585
R322 B.n657 B.n656 585
R323 B.n658 B.n383 585
R324 B.n660 B.n659 585
R325 B.n662 B.n382 585
R326 B.n663 B.n381 585
R327 B.n666 B.n665 585
R328 B.n667 B.n380 585
R329 B.n380 B.n379 585
R330 B.n672 B.n671 585
R331 B.n671 B.n670 585
R332 B.n673 B.n376 585
R333 B.n376 B.n375 585
R334 B.n675 B.n674 585
R335 B.n676 B.n675 585
R336 B.n370 B.n369 585
R337 B.n371 B.n370 585
R338 B.n685 B.n684 585
R339 B.n684 B.n683 585
R340 B.n686 B.n368 585
R341 B.n682 B.n368 585
R342 B.n688 B.n687 585
R343 B.n689 B.n688 585
R344 B.n363 B.n362 585
R345 B.n364 B.n363 585
R346 B.n697 B.n696 585
R347 B.n696 B.n695 585
R348 B.n698 B.n361 585
R349 B.n361 B.n360 585
R350 B.n700 B.n699 585
R351 B.n701 B.n700 585
R352 B.n355 B.n354 585
R353 B.n356 B.n355 585
R354 B.n709 B.n708 585
R355 B.n708 B.n707 585
R356 B.n710 B.n353 585
R357 B.n353 B.n352 585
R358 B.n712 B.n711 585
R359 B.n713 B.n712 585
R360 B.n347 B.n346 585
R361 B.n348 B.n347 585
R362 B.n721 B.n720 585
R363 B.n720 B.n719 585
R364 B.n722 B.n345 585
R365 B.n345 B.n344 585
R366 B.n724 B.n723 585
R367 B.n725 B.n724 585
R368 B.n339 B.n338 585
R369 B.n340 B.n339 585
R370 B.n734 B.n733 585
R371 B.n733 B.n732 585
R372 B.n735 B.n337 585
R373 B.n337 B.n336 585
R374 B.n737 B.n736 585
R375 B.n738 B.n737 585
R376 B.n3 B.n0 585
R377 B.n4 B.n3 585
R378 B.n826 B.n1 585
R379 B.n827 B.n826 585
R380 B.n825 B.n824 585
R381 B.n825 B.n8 585
R382 B.n823 B.n9 585
R383 B.n747 B.n9 585
R384 B.n822 B.n821 585
R385 B.n821 B.n820 585
R386 B.n11 B.n10 585
R387 B.n819 B.n11 585
R388 B.n817 B.n816 585
R389 B.n818 B.n817 585
R390 B.n815 B.n16 585
R391 B.n16 B.n15 585
R392 B.n814 B.n813 585
R393 B.n813 B.n812 585
R394 B.n18 B.n17 585
R395 B.n811 B.n18 585
R396 B.n809 B.n808 585
R397 B.n810 B.n809 585
R398 B.n807 B.n23 585
R399 B.n23 B.n22 585
R400 B.n806 B.n805 585
R401 B.n805 B.n804 585
R402 B.n25 B.n24 585
R403 B.n803 B.n25 585
R404 B.n801 B.n800 585
R405 B.n802 B.n801 585
R406 B.n799 B.n30 585
R407 B.n30 B.n29 585
R408 B.n798 B.n797 585
R409 B.n797 B.n796 585
R410 B.n32 B.n31 585
R411 B.n795 B.n32 585
R412 B.n793 B.n792 585
R413 B.n794 B.n793 585
R414 B.n791 B.n36 585
R415 B.n39 B.n36 585
R416 B.n790 B.n789 585
R417 B.n789 B.n788 585
R418 B.n38 B.n37 585
R419 B.n787 B.n38 585
R420 B.n785 B.n784 585
R421 B.n786 B.n785 585
R422 B.n783 B.n44 585
R423 B.n44 B.n43 585
R424 B.n782 B.n781 585
R425 B.n781 B.n780 585
R426 B.n830 B.n829 585
R427 B.n828 B.n2 585
R428 B.n108 B.t16 549.766
R429 B.n105 B.t9 549.766
R430 B.n560 B.t5 549.766
R431 B.n412 B.t13 549.766
R432 B.n781 B.n46 492.5
R433 B.n777 B.n47 492.5
R434 B.n669 B.n380 492.5
R435 B.n671 B.n378 492.5
R436 B.n105 B.t11 370.243
R437 B.n560 B.t8 370.243
R438 B.n108 B.t17 370.243
R439 B.n412 B.t15 370.243
R440 B.n106 B.t12 342.897
R441 B.n561 B.t7 342.897
R442 B.n109 B.t18 342.897
R443 B.n413 B.t14 342.897
R444 B.n779 B.n778 256.663
R445 B.n779 B.n103 256.663
R446 B.n779 B.n102 256.663
R447 B.n779 B.n101 256.663
R448 B.n779 B.n100 256.663
R449 B.n779 B.n99 256.663
R450 B.n779 B.n98 256.663
R451 B.n779 B.n97 256.663
R452 B.n779 B.n96 256.663
R453 B.n779 B.n95 256.663
R454 B.n779 B.n94 256.663
R455 B.n779 B.n93 256.663
R456 B.n779 B.n92 256.663
R457 B.n779 B.n91 256.663
R458 B.n779 B.n90 256.663
R459 B.n779 B.n89 256.663
R460 B.n779 B.n88 256.663
R461 B.n779 B.n87 256.663
R462 B.n779 B.n86 256.663
R463 B.n779 B.n85 256.663
R464 B.n779 B.n84 256.663
R465 B.n779 B.n83 256.663
R466 B.n779 B.n82 256.663
R467 B.n779 B.n81 256.663
R468 B.n779 B.n80 256.663
R469 B.n779 B.n79 256.663
R470 B.n779 B.n78 256.663
R471 B.n779 B.n77 256.663
R472 B.n779 B.n76 256.663
R473 B.n779 B.n75 256.663
R474 B.n779 B.n74 256.663
R475 B.n779 B.n73 256.663
R476 B.n779 B.n72 256.663
R477 B.n779 B.n71 256.663
R478 B.n779 B.n70 256.663
R479 B.n779 B.n69 256.663
R480 B.n779 B.n68 256.663
R481 B.n779 B.n67 256.663
R482 B.n779 B.n66 256.663
R483 B.n779 B.n65 256.663
R484 B.n779 B.n64 256.663
R485 B.n779 B.n63 256.663
R486 B.n779 B.n62 256.663
R487 B.n779 B.n61 256.663
R488 B.n779 B.n60 256.663
R489 B.n779 B.n59 256.663
R490 B.n779 B.n58 256.663
R491 B.n779 B.n57 256.663
R492 B.n779 B.n56 256.663
R493 B.n779 B.n55 256.663
R494 B.n779 B.n54 256.663
R495 B.n779 B.n53 256.663
R496 B.n779 B.n52 256.663
R497 B.n779 B.n51 256.663
R498 B.n779 B.n50 256.663
R499 B.n779 B.n49 256.663
R500 B.n779 B.n48 256.663
R501 B.n440 B.n379 256.663
R502 B.n443 B.n379 256.663
R503 B.n449 B.n379 256.663
R504 B.n451 B.n379 256.663
R505 B.n457 B.n379 256.663
R506 B.n459 B.n379 256.663
R507 B.n465 B.n379 256.663
R508 B.n467 B.n379 256.663
R509 B.n473 B.n379 256.663
R510 B.n475 B.n379 256.663
R511 B.n481 B.n379 256.663
R512 B.n483 B.n379 256.663
R513 B.n489 B.n379 256.663
R514 B.n491 B.n379 256.663
R515 B.n497 B.n379 256.663
R516 B.n499 B.n379 256.663
R517 B.n505 B.n379 256.663
R518 B.n507 B.n379 256.663
R519 B.n513 B.n379 256.663
R520 B.n515 B.n379 256.663
R521 B.n521 B.n379 256.663
R522 B.n523 B.n379 256.663
R523 B.n529 B.n379 256.663
R524 B.n531 B.n379 256.663
R525 B.n537 B.n379 256.663
R526 B.n539 B.n379 256.663
R527 B.n546 B.n379 256.663
R528 B.n548 B.n379 256.663
R529 B.n554 B.n379 256.663
R530 B.n556 B.n379 256.663
R531 B.n565 B.n379 256.663
R532 B.n567 B.n379 256.663
R533 B.n573 B.n379 256.663
R534 B.n575 B.n379 256.663
R535 B.n581 B.n379 256.663
R536 B.n583 B.n379 256.663
R537 B.n589 B.n379 256.663
R538 B.n591 B.n379 256.663
R539 B.n597 B.n379 256.663
R540 B.n599 B.n379 256.663
R541 B.n605 B.n379 256.663
R542 B.n607 B.n379 256.663
R543 B.n613 B.n379 256.663
R544 B.n615 B.n379 256.663
R545 B.n621 B.n379 256.663
R546 B.n623 B.n379 256.663
R547 B.n629 B.n379 256.663
R548 B.n631 B.n379 256.663
R549 B.n637 B.n379 256.663
R550 B.n639 B.n379 256.663
R551 B.n645 B.n379 256.663
R552 B.n647 B.n379 256.663
R553 B.n653 B.n379 256.663
R554 B.n655 B.n379 256.663
R555 B.n661 B.n379 256.663
R556 B.n664 B.n379 256.663
R557 B.n832 B.n831 256.663
R558 B.n113 B.n112 163.367
R559 B.n117 B.n116 163.367
R560 B.n121 B.n120 163.367
R561 B.n125 B.n124 163.367
R562 B.n129 B.n128 163.367
R563 B.n133 B.n132 163.367
R564 B.n137 B.n136 163.367
R565 B.n141 B.n140 163.367
R566 B.n145 B.n144 163.367
R567 B.n149 B.n148 163.367
R568 B.n153 B.n152 163.367
R569 B.n157 B.n156 163.367
R570 B.n161 B.n160 163.367
R571 B.n165 B.n164 163.367
R572 B.n169 B.n168 163.367
R573 B.n173 B.n172 163.367
R574 B.n177 B.n176 163.367
R575 B.n181 B.n180 163.367
R576 B.n185 B.n184 163.367
R577 B.n189 B.n188 163.367
R578 B.n193 B.n192 163.367
R579 B.n197 B.n196 163.367
R580 B.n201 B.n200 163.367
R581 B.n205 B.n204 163.367
R582 B.n209 B.n208 163.367
R583 B.n213 B.n212 163.367
R584 B.n217 B.n216 163.367
R585 B.n221 B.n220 163.367
R586 B.n225 B.n224 163.367
R587 B.n229 B.n228 163.367
R588 B.n233 B.n232 163.367
R589 B.n237 B.n236 163.367
R590 B.n241 B.n240 163.367
R591 B.n245 B.n244 163.367
R592 B.n249 B.n248 163.367
R593 B.n253 B.n252 163.367
R594 B.n257 B.n256 163.367
R595 B.n261 B.n260 163.367
R596 B.n265 B.n264 163.367
R597 B.n269 B.n268 163.367
R598 B.n273 B.n272 163.367
R599 B.n277 B.n276 163.367
R600 B.n281 B.n280 163.367
R601 B.n285 B.n284 163.367
R602 B.n289 B.n288 163.367
R603 B.n293 B.n292 163.367
R604 B.n297 B.n296 163.367
R605 B.n301 B.n300 163.367
R606 B.n305 B.n304 163.367
R607 B.n309 B.n308 163.367
R608 B.n313 B.n312 163.367
R609 B.n317 B.n316 163.367
R610 B.n321 B.n320 163.367
R611 B.n325 B.n324 163.367
R612 B.n329 B.n328 163.367
R613 B.n331 B.n104 163.367
R614 B.n669 B.n374 163.367
R615 B.n677 B.n374 163.367
R616 B.n677 B.n372 163.367
R617 B.n681 B.n372 163.367
R618 B.n681 B.n367 163.367
R619 B.n690 B.n367 163.367
R620 B.n690 B.n365 163.367
R621 B.n694 B.n365 163.367
R622 B.n694 B.n359 163.367
R623 B.n702 B.n359 163.367
R624 B.n702 B.n357 163.367
R625 B.n706 B.n357 163.367
R626 B.n706 B.n351 163.367
R627 B.n714 B.n351 163.367
R628 B.n714 B.n349 163.367
R629 B.n718 B.n349 163.367
R630 B.n718 B.n343 163.367
R631 B.n726 B.n343 163.367
R632 B.n726 B.n341 163.367
R633 B.n731 B.n341 163.367
R634 B.n731 B.n335 163.367
R635 B.n739 B.n335 163.367
R636 B.n740 B.n739 163.367
R637 B.n740 B.n5 163.367
R638 B.n6 B.n5 163.367
R639 B.n7 B.n6 163.367
R640 B.n746 B.n7 163.367
R641 B.n748 B.n746 163.367
R642 B.n748 B.n12 163.367
R643 B.n13 B.n12 163.367
R644 B.n14 B.n13 163.367
R645 B.n753 B.n14 163.367
R646 B.n753 B.n19 163.367
R647 B.n20 B.n19 163.367
R648 B.n21 B.n20 163.367
R649 B.n758 B.n21 163.367
R650 B.n758 B.n26 163.367
R651 B.n27 B.n26 163.367
R652 B.n28 B.n27 163.367
R653 B.n763 B.n28 163.367
R654 B.n763 B.n33 163.367
R655 B.n34 B.n33 163.367
R656 B.n35 B.n34 163.367
R657 B.n768 B.n35 163.367
R658 B.n768 B.n40 163.367
R659 B.n41 B.n40 163.367
R660 B.n42 B.n41 163.367
R661 B.n773 B.n42 163.367
R662 B.n773 B.n47 163.367
R663 B.n442 B.n441 163.367
R664 B.n444 B.n442 163.367
R665 B.n448 B.n437 163.367
R666 B.n452 B.n450 163.367
R667 B.n456 B.n435 163.367
R668 B.n460 B.n458 163.367
R669 B.n464 B.n433 163.367
R670 B.n468 B.n466 163.367
R671 B.n472 B.n431 163.367
R672 B.n476 B.n474 163.367
R673 B.n480 B.n429 163.367
R674 B.n484 B.n482 163.367
R675 B.n488 B.n427 163.367
R676 B.n492 B.n490 163.367
R677 B.n496 B.n425 163.367
R678 B.n500 B.n498 163.367
R679 B.n504 B.n423 163.367
R680 B.n508 B.n506 163.367
R681 B.n512 B.n421 163.367
R682 B.n516 B.n514 163.367
R683 B.n520 B.n419 163.367
R684 B.n524 B.n522 163.367
R685 B.n528 B.n417 163.367
R686 B.n532 B.n530 163.367
R687 B.n536 B.n415 163.367
R688 B.n540 B.n538 163.367
R689 B.n545 B.n411 163.367
R690 B.n549 B.n547 163.367
R691 B.n553 B.n409 163.367
R692 B.n557 B.n555 163.367
R693 B.n564 B.n407 163.367
R694 B.n568 B.n566 163.367
R695 B.n572 B.n405 163.367
R696 B.n576 B.n574 163.367
R697 B.n580 B.n403 163.367
R698 B.n584 B.n582 163.367
R699 B.n588 B.n401 163.367
R700 B.n592 B.n590 163.367
R701 B.n596 B.n399 163.367
R702 B.n600 B.n598 163.367
R703 B.n604 B.n397 163.367
R704 B.n608 B.n606 163.367
R705 B.n612 B.n395 163.367
R706 B.n616 B.n614 163.367
R707 B.n620 B.n393 163.367
R708 B.n624 B.n622 163.367
R709 B.n628 B.n391 163.367
R710 B.n632 B.n630 163.367
R711 B.n636 B.n389 163.367
R712 B.n640 B.n638 163.367
R713 B.n644 B.n387 163.367
R714 B.n648 B.n646 163.367
R715 B.n652 B.n385 163.367
R716 B.n656 B.n654 163.367
R717 B.n660 B.n383 163.367
R718 B.n663 B.n662 163.367
R719 B.n665 B.n380 163.367
R720 B.n671 B.n376 163.367
R721 B.n675 B.n376 163.367
R722 B.n675 B.n370 163.367
R723 B.n684 B.n370 163.367
R724 B.n684 B.n368 163.367
R725 B.n688 B.n368 163.367
R726 B.n688 B.n363 163.367
R727 B.n696 B.n363 163.367
R728 B.n696 B.n361 163.367
R729 B.n700 B.n361 163.367
R730 B.n700 B.n355 163.367
R731 B.n708 B.n355 163.367
R732 B.n708 B.n353 163.367
R733 B.n712 B.n353 163.367
R734 B.n712 B.n347 163.367
R735 B.n720 B.n347 163.367
R736 B.n720 B.n345 163.367
R737 B.n724 B.n345 163.367
R738 B.n724 B.n339 163.367
R739 B.n733 B.n339 163.367
R740 B.n733 B.n337 163.367
R741 B.n737 B.n337 163.367
R742 B.n737 B.n3 163.367
R743 B.n830 B.n3 163.367
R744 B.n826 B.n2 163.367
R745 B.n826 B.n825 163.367
R746 B.n825 B.n9 163.367
R747 B.n821 B.n9 163.367
R748 B.n821 B.n11 163.367
R749 B.n817 B.n11 163.367
R750 B.n817 B.n16 163.367
R751 B.n813 B.n16 163.367
R752 B.n813 B.n18 163.367
R753 B.n809 B.n18 163.367
R754 B.n809 B.n23 163.367
R755 B.n805 B.n23 163.367
R756 B.n805 B.n25 163.367
R757 B.n801 B.n25 163.367
R758 B.n801 B.n30 163.367
R759 B.n797 B.n30 163.367
R760 B.n797 B.n32 163.367
R761 B.n793 B.n32 163.367
R762 B.n793 B.n36 163.367
R763 B.n789 B.n36 163.367
R764 B.n789 B.n38 163.367
R765 B.n785 B.n38 163.367
R766 B.n785 B.n44 163.367
R767 B.n781 B.n44 163.367
R768 B.n670 B.n379 72.4698
R769 B.n780 B.n779 72.4698
R770 B.n48 B.n46 71.676
R771 B.n113 B.n49 71.676
R772 B.n117 B.n50 71.676
R773 B.n121 B.n51 71.676
R774 B.n125 B.n52 71.676
R775 B.n129 B.n53 71.676
R776 B.n133 B.n54 71.676
R777 B.n137 B.n55 71.676
R778 B.n141 B.n56 71.676
R779 B.n145 B.n57 71.676
R780 B.n149 B.n58 71.676
R781 B.n153 B.n59 71.676
R782 B.n157 B.n60 71.676
R783 B.n161 B.n61 71.676
R784 B.n165 B.n62 71.676
R785 B.n169 B.n63 71.676
R786 B.n173 B.n64 71.676
R787 B.n177 B.n65 71.676
R788 B.n181 B.n66 71.676
R789 B.n185 B.n67 71.676
R790 B.n189 B.n68 71.676
R791 B.n193 B.n69 71.676
R792 B.n197 B.n70 71.676
R793 B.n201 B.n71 71.676
R794 B.n205 B.n72 71.676
R795 B.n209 B.n73 71.676
R796 B.n213 B.n74 71.676
R797 B.n217 B.n75 71.676
R798 B.n221 B.n76 71.676
R799 B.n225 B.n77 71.676
R800 B.n229 B.n78 71.676
R801 B.n233 B.n79 71.676
R802 B.n237 B.n80 71.676
R803 B.n241 B.n81 71.676
R804 B.n245 B.n82 71.676
R805 B.n249 B.n83 71.676
R806 B.n253 B.n84 71.676
R807 B.n257 B.n85 71.676
R808 B.n261 B.n86 71.676
R809 B.n265 B.n87 71.676
R810 B.n269 B.n88 71.676
R811 B.n273 B.n89 71.676
R812 B.n277 B.n90 71.676
R813 B.n281 B.n91 71.676
R814 B.n285 B.n92 71.676
R815 B.n289 B.n93 71.676
R816 B.n293 B.n94 71.676
R817 B.n297 B.n95 71.676
R818 B.n301 B.n96 71.676
R819 B.n305 B.n97 71.676
R820 B.n309 B.n98 71.676
R821 B.n313 B.n99 71.676
R822 B.n317 B.n100 71.676
R823 B.n321 B.n101 71.676
R824 B.n325 B.n102 71.676
R825 B.n329 B.n103 71.676
R826 B.n778 B.n104 71.676
R827 B.n778 B.n777 71.676
R828 B.n331 B.n103 71.676
R829 B.n328 B.n102 71.676
R830 B.n324 B.n101 71.676
R831 B.n320 B.n100 71.676
R832 B.n316 B.n99 71.676
R833 B.n312 B.n98 71.676
R834 B.n308 B.n97 71.676
R835 B.n304 B.n96 71.676
R836 B.n300 B.n95 71.676
R837 B.n296 B.n94 71.676
R838 B.n292 B.n93 71.676
R839 B.n288 B.n92 71.676
R840 B.n284 B.n91 71.676
R841 B.n280 B.n90 71.676
R842 B.n276 B.n89 71.676
R843 B.n272 B.n88 71.676
R844 B.n268 B.n87 71.676
R845 B.n264 B.n86 71.676
R846 B.n260 B.n85 71.676
R847 B.n256 B.n84 71.676
R848 B.n252 B.n83 71.676
R849 B.n248 B.n82 71.676
R850 B.n244 B.n81 71.676
R851 B.n240 B.n80 71.676
R852 B.n236 B.n79 71.676
R853 B.n232 B.n78 71.676
R854 B.n228 B.n77 71.676
R855 B.n224 B.n76 71.676
R856 B.n220 B.n75 71.676
R857 B.n216 B.n74 71.676
R858 B.n212 B.n73 71.676
R859 B.n208 B.n72 71.676
R860 B.n204 B.n71 71.676
R861 B.n200 B.n70 71.676
R862 B.n196 B.n69 71.676
R863 B.n192 B.n68 71.676
R864 B.n188 B.n67 71.676
R865 B.n184 B.n66 71.676
R866 B.n180 B.n65 71.676
R867 B.n176 B.n64 71.676
R868 B.n172 B.n63 71.676
R869 B.n168 B.n62 71.676
R870 B.n164 B.n61 71.676
R871 B.n160 B.n60 71.676
R872 B.n156 B.n59 71.676
R873 B.n152 B.n58 71.676
R874 B.n148 B.n57 71.676
R875 B.n144 B.n56 71.676
R876 B.n140 B.n55 71.676
R877 B.n136 B.n54 71.676
R878 B.n132 B.n53 71.676
R879 B.n128 B.n52 71.676
R880 B.n124 B.n51 71.676
R881 B.n120 B.n50 71.676
R882 B.n116 B.n49 71.676
R883 B.n112 B.n48 71.676
R884 B.n440 B.n378 71.676
R885 B.n444 B.n443 71.676
R886 B.n449 B.n448 71.676
R887 B.n452 B.n451 71.676
R888 B.n457 B.n456 71.676
R889 B.n460 B.n459 71.676
R890 B.n465 B.n464 71.676
R891 B.n468 B.n467 71.676
R892 B.n473 B.n472 71.676
R893 B.n476 B.n475 71.676
R894 B.n481 B.n480 71.676
R895 B.n484 B.n483 71.676
R896 B.n489 B.n488 71.676
R897 B.n492 B.n491 71.676
R898 B.n497 B.n496 71.676
R899 B.n500 B.n499 71.676
R900 B.n505 B.n504 71.676
R901 B.n508 B.n507 71.676
R902 B.n513 B.n512 71.676
R903 B.n516 B.n515 71.676
R904 B.n521 B.n520 71.676
R905 B.n524 B.n523 71.676
R906 B.n529 B.n528 71.676
R907 B.n532 B.n531 71.676
R908 B.n537 B.n536 71.676
R909 B.n540 B.n539 71.676
R910 B.n546 B.n545 71.676
R911 B.n549 B.n548 71.676
R912 B.n554 B.n553 71.676
R913 B.n557 B.n556 71.676
R914 B.n565 B.n564 71.676
R915 B.n568 B.n567 71.676
R916 B.n573 B.n572 71.676
R917 B.n576 B.n575 71.676
R918 B.n581 B.n580 71.676
R919 B.n584 B.n583 71.676
R920 B.n589 B.n588 71.676
R921 B.n592 B.n591 71.676
R922 B.n597 B.n596 71.676
R923 B.n600 B.n599 71.676
R924 B.n605 B.n604 71.676
R925 B.n608 B.n607 71.676
R926 B.n613 B.n612 71.676
R927 B.n616 B.n615 71.676
R928 B.n621 B.n620 71.676
R929 B.n624 B.n623 71.676
R930 B.n629 B.n628 71.676
R931 B.n632 B.n631 71.676
R932 B.n637 B.n636 71.676
R933 B.n640 B.n639 71.676
R934 B.n645 B.n644 71.676
R935 B.n648 B.n647 71.676
R936 B.n653 B.n652 71.676
R937 B.n656 B.n655 71.676
R938 B.n661 B.n660 71.676
R939 B.n664 B.n663 71.676
R940 B.n441 B.n440 71.676
R941 B.n443 B.n437 71.676
R942 B.n450 B.n449 71.676
R943 B.n451 B.n435 71.676
R944 B.n458 B.n457 71.676
R945 B.n459 B.n433 71.676
R946 B.n466 B.n465 71.676
R947 B.n467 B.n431 71.676
R948 B.n474 B.n473 71.676
R949 B.n475 B.n429 71.676
R950 B.n482 B.n481 71.676
R951 B.n483 B.n427 71.676
R952 B.n490 B.n489 71.676
R953 B.n491 B.n425 71.676
R954 B.n498 B.n497 71.676
R955 B.n499 B.n423 71.676
R956 B.n506 B.n505 71.676
R957 B.n507 B.n421 71.676
R958 B.n514 B.n513 71.676
R959 B.n515 B.n419 71.676
R960 B.n522 B.n521 71.676
R961 B.n523 B.n417 71.676
R962 B.n530 B.n529 71.676
R963 B.n531 B.n415 71.676
R964 B.n538 B.n537 71.676
R965 B.n539 B.n411 71.676
R966 B.n547 B.n546 71.676
R967 B.n548 B.n409 71.676
R968 B.n555 B.n554 71.676
R969 B.n556 B.n407 71.676
R970 B.n566 B.n565 71.676
R971 B.n567 B.n405 71.676
R972 B.n574 B.n573 71.676
R973 B.n575 B.n403 71.676
R974 B.n582 B.n581 71.676
R975 B.n583 B.n401 71.676
R976 B.n590 B.n589 71.676
R977 B.n591 B.n399 71.676
R978 B.n598 B.n597 71.676
R979 B.n599 B.n397 71.676
R980 B.n606 B.n605 71.676
R981 B.n607 B.n395 71.676
R982 B.n614 B.n613 71.676
R983 B.n615 B.n393 71.676
R984 B.n622 B.n621 71.676
R985 B.n623 B.n391 71.676
R986 B.n630 B.n629 71.676
R987 B.n631 B.n389 71.676
R988 B.n638 B.n637 71.676
R989 B.n639 B.n387 71.676
R990 B.n646 B.n645 71.676
R991 B.n647 B.n385 71.676
R992 B.n654 B.n653 71.676
R993 B.n655 B.n383 71.676
R994 B.n662 B.n661 71.676
R995 B.n665 B.n664 71.676
R996 B.n831 B.n830 71.676
R997 B.n831 B.n2 71.676
R998 B.n110 B.n109 59.5399
R999 B.n107 B.n106 59.5399
R1000 B.n562 B.n561 59.5399
R1001 B.n542 B.n413 59.5399
R1002 B.n670 B.n375 35.9707
R1003 B.n676 B.n375 35.9707
R1004 B.n676 B.n371 35.9707
R1005 B.n683 B.n371 35.9707
R1006 B.n683 B.n682 35.9707
R1007 B.n689 B.n364 35.9707
R1008 B.n695 B.n364 35.9707
R1009 B.n695 B.n360 35.9707
R1010 B.n701 B.n360 35.9707
R1011 B.n701 B.n356 35.9707
R1012 B.n707 B.n356 35.9707
R1013 B.n713 B.n352 35.9707
R1014 B.n713 B.n348 35.9707
R1015 B.n719 B.n348 35.9707
R1016 B.n725 B.n344 35.9707
R1017 B.n725 B.n340 35.9707
R1018 B.n732 B.n340 35.9707
R1019 B.n738 B.n336 35.9707
R1020 B.n738 B.n4 35.9707
R1021 B.n829 B.n4 35.9707
R1022 B.n829 B.n828 35.9707
R1023 B.n828 B.n827 35.9707
R1024 B.n827 B.n8 35.9707
R1025 B.n747 B.n8 35.9707
R1026 B.n820 B.n819 35.9707
R1027 B.n819 B.n818 35.9707
R1028 B.n818 B.n15 35.9707
R1029 B.n812 B.n811 35.9707
R1030 B.n811 B.n810 35.9707
R1031 B.n810 B.n22 35.9707
R1032 B.n804 B.n803 35.9707
R1033 B.n803 B.n802 35.9707
R1034 B.n802 B.n29 35.9707
R1035 B.n796 B.n29 35.9707
R1036 B.n796 B.n795 35.9707
R1037 B.n795 B.n794 35.9707
R1038 B.n788 B.n39 35.9707
R1039 B.n788 B.n787 35.9707
R1040 B.n787 B.n786 35.9707
R1041 B.n786 B.n43 35.9707
R1042 B.n780 B.n43 35.9707
R1043 B.n672 B.n377 32.0005
R1044 B.n668 B.n667 32.0005
R1045 B.n776 B.n775 32.0005
R1046 B.n782 B.n45 32.0005
R1047 B.n689 B.t6 29.623
R1048 B.n732 B.t0 29.623
R1049 B.n820 B.t3 29.623
R1050 B.n794 B.t10 29.623
R1051 B.n109 B.n108 27.346
R1052 B.n106 B.n105 27.346
R1053 B.n561 B.n560 27.346
R1054 B.n413 B.n412 27.346
R1055 B.n719 B.t19 24.3333
R1056 B.n812 B.t2 24.3333
R1057 B.n707 B.t4 19.0435
R1058 B.n804 B.t1 19.0435
R1059 B B.n832 18.0485
R1060 B.t4 B.n352 16.9276
R1061 B.t1 B.n22 16.9276
R1062 B.t19 B.n344 11.6379
R1063 B.t2 B.n15 11.6379
R1064 B.n673 B.n672 10.6151
R1065 B.n674 B.n673 10.6151
R1066 B.n674 B.n369 10.6151
R1067 B.n685 B.n369 10.6151
R1068 B.n686 B.n685 10.6151
R1069 B.n687 B.n686 10.6151
R1070 B.n687 B.n362 10.6151
R1071 B.n697 B.n362 10.6151
R1072 B.n698 B.n697 10.6151
R1073 B.n699 B.n698 10.6151
R1074 B.n699 B.n354 10.6151
R1075 B.n709 B.n354 10.6151
R1076 B.n710 B.n709 10.6151
R1077 B.n711 B.n710 10.6151
R1078 B.n711 B.n346 10.6151
R1079 B.n721 B.n346 10.6151
R1080 B.n722 B.n721 10.6151
R1081 B.n723 B.n722 10.6151
R1082 B.n723 B.n338 10.6151
R1083 B.n734 B.n338 10.6151
R1084 B.n735 B.n734 10.6151
R1085 B.n736 B.n735 10.6151
R1086 B.n736 B.n0 10.6151
R1087 B.n439 B.n377 10.6151
R1088 B.n439 B.n438 10.6151
R1089 B.n445 B.n438 10.6151
R1090 B.n446 B.n445 10.6151
R1091 B.n447 B.n446 10.6151
R1092 B.n447 B.n436 10.6151
R1093 B.n453 B.n436 10.6151
R1094 B.n454 B.n453 10.6151
R1095 B.n455 B.n454 10.6151
R1096 B.n455 B.n434 10.6151
R1097 B.n461 B.n434 10.6151
R1098 B.n462 B.n461 10.6151
R1099 B.n463 B.n462 10.6151
R1100 B.n463 B.n432 10.6151
R1101 B.n469 B.n432 10.6151
R1102 B.n470 B.n469 10.6151
R1103 B.n471 B.n470 10.6151
R1104 B.n471 B.n430 10.6151
R1105 B.n477 B.n430 10.6151
R1106 B.n478 B.n477 10.6151
R1107 B.n479 B.n478 10.6151
R1108 B.n479 B.n428 10.6151
R1109 B.n485 B.n428 10.6151
R1110 B.n486 B.n485 10.6151
R1111 B.n487 B.n486 10.6151
R1112 B.n487 B.n426 10.6151
R1113 B.n493 B.n426 10.6151
R1114 B.n494 B.n493 10.6151
R1115 B.n495 B.n494 10.6151
R1116 B.n495 B.n424 10.6151
R1117 B.n501 B.n424 10.6151
R1118 B.n502 B.n501 10.6151
R1119 B.n503 B.n502 10.6151
R1120 B.n503 B.n422 10.6151
R1121 B.n509 B.n422 10.6151
R1122 B.n510 B.n509 10.6151
R1123 B.n511 B.n510 10.6151
R1124 B.n511 B.n420 10.6151
R1125 B.n517 B.n420 10.6151
R1126 B.n518 B.n517 10.6151
R1127 B.n519 B.n518 10.6151
R1128 B.n519 B.n418 10.6151
R1129 B.n525 B.n418 10.6151
R1130 B.n526 B.n525 10.6151
R1131 B.n527 B.n526 10.6151
R1132 B.n527 B.n416 10.6151
R1133 B.n533 B.n416 10.6151
R1134 B.n534 B.n533 10.6151
R1135 B.n535 B.n534 10.6151
R1136 B.n535 B.n414 10.6151
R1137 B.n541 B.n414 10.6151
R1138 B.n544 B.n543 10.6151
R1139 B.n544 B.n410 10.6151
R1140 B.n550 B.n410 10.6151
R1141 B.n551 B.n550 10.6151
R1142 B.n552 B.n551 10.6151
R1143 B.n552 B.n408 10.6151
R1144 B.n558 B.n408 10.6151
R1145 B.n559 B.n558 10.6151
R1146 B.n563 B.n559 10.6151
R1147 B.n569 B.n406 10.6151
R1148 B.n570 B.n569 10.6151
R1149 B.n571 B.n570 10.6151
R1150 B.n571 B.n404 10.6151
R1151 B.n577 B.n404 10.6151
R1152 B.n578 B.n577 10.6151
R1153 B.n579 B.n578 10.6151
R1154 B.n579 B.n402 10.6151
R1155 B.n585 B.n402 10.6151
R1156 B.n586 B.n585 10.6151
R1157 B.n587 B.n586 10.6151
R1158 B.n587 B.n400 10.6151
R1159 B.n593 B.n400 10.6151
R1160 B.n594 B.n593 10.6151
R1161 B.n595 B.n594 10.6151
R1162 B.n595 B.n398 10.6151
R1163 B.n601 B.n398 10.6151
R1164 B.n602 B.n601 10.6151
R1165 B.n603 B.n602 10.6151
R1166 B.n603 B.n396 10.6151
R1167 B.n609 B.n396 10.6151
R1168 B.n610 B.n609 10.6151
R1169 B.n611 B.n610 10.6151
R1170 B.n611 B.n394 10.6151
R1171 B.n617 B.n394 10.6151
R1172 B.n618 B.n617 10.6151
R1173 B.n619 B.n618 10.6151
R1174 B.n619 B.n392 10.6151
R1175 B.n625 B.n392 10.6151
R1176 B.n626 B.n625 10.6151
R1177 B.n627 B.n626 10.6151
R1178 B.n627 B.n390 10.6151
R1179 B.n633 B.n390 10.6151
R1180 B.n634 B.n633 10.6151
R1181 B.n635 B.n634 10.6151
R1182 B.n635 B.n388 10.6151
R1183 B.n641 B.n388 10.6151
R1184 B.n642 B.n641 10.6151
R1185 B.n643 B.n642 10.6151
R1186 B.n643 B.n386 10.6151
R1187 B.n649 B.n386 10.6151
R1188 B.n650 B.n649 10.6151
R1189 B.n651 B.n650 10.6151
R1190 B.n651 B.n384 10.6151
R1191 B.n657 B.n384 10.6151
R1192 B.n658 B.n657 10.6151
R1193 B.n659 B.n658 10.6151
R1194 B.n659 B.n382 10.6151
R1195 B.n382 B.n381 10.6151
R1196 B.n666 B.n381 10.6151
R1197 B.n667 B.n666 10.6151
R1198 B.n668 B.n373 10.6151
R1199 B.n678 B.n373 10.6151
R1200 B.n679 B.n678 10.6151
R1201 B.n680 B.n679 10.6151
R1202 B.n680 B.n366 10.6151
R1203 B.n691 B.n366 10.6151
R1204 B.n692 B.n691 10.6151
R1205 B.n693 B.n692 10.6151
R1206 B.n693 B.n358 10.6151
R1207 B.n703 B.n358 10.6151
R1208 B.n704 B.n703 10.6151
R1209 B.n705 B.n704 10.6151
R1210 B.n705 B.n350 10.6151
R1211 B.n715 B.n350 10.6151
R1212 B.n716 B.n715 10.6151
R1213 B.n717 B.n716 10.6151
R1214 B.n717 B.n342 10.6151
R1215 B.n727 B.n342 10.6151
R1216 B.n728 B.n727 10.6151
R1217 B.n730 B.n728 10.6151
R1218 B.n730 B.n729 10.6151
R1219 B.n729 B.n334 10.6151
R1220 B.n741 B.n334 10.6151
R1221 B.n742 B.n741 10.6151
R1222 B.n743 B.n742 10.6151
R1223 B.n744 B.n743 10.6151
R1224 B.n745 B.n744 10.6151
R1225 B.n749 B.n745 10.6151
R1226 B.n750 B.n749 10.6151
R1227 B.n751 B.n750 10.6151
R1228 B.n752 B.n751 10.6151
R1229 B.n754 B.n752 10.6151
R1230 B.n755 B.n754 10.6151
R1231 B.n756 B.n755 10.6151
R1232 B.n757 B.n756 10.6151
R1233 B.n759 B.n757 10.6151
R1234 B.n760 B.n759 10.6151
R1235 B.n761 B.n760 10.6151
R1236 B.n762 B.n761 10.6151
R1237 B.n764 B.n762 10.6151
R1238 B.n765 B.n764 10.6151
R1239 B.n766 B.n765 10.6151
R1240 B.n767 B.n766 10.6151
R1241 B.n769 B.n767 10.6151
R1242 B.n770 B.n769 10.6151
R1243 B.n771 B.n770 10.6151
R1244 B.n772 B.n771 10.6151
R1245 B.n774 B.n772 10.6151
R1246 B.n775 B.n774 10.6151
R1247 B.n824 B.n1 10.6151
R1248 B.n824 B.n823 10.6151
R1249 B.n823 B.n822 10.6151
R1250 B.n822 B.n10 10.6151
R1251 B.n816 B.n10 10.6151
R1252 B.n816 B.n815 10.6151
R1253 B.n815 B.n814 10.6151
R1254 B.n814 B.n17 10.6151
R1255 B.n808 B.n17 10.6151
R1256 B.n808 B.n807 10.6151
R1257 B.n807 B.n806 10.6151
R1258 B.n806 B.n24 10.6151
R1259 B.n800 B.n24 10.6151
R1260 B.n800 B.n799 10.6151
R1261 B.n799 B.n798 10.6151
R1262 B.n798 B.n31 10.6151
R1263 B.n792 B.n31 10.6151
R1264 B.n792 B.n791 10.6151
R1265 B.n791 B.n790 10.6151
R1266 B.n790 B.n37 10.6151
R1267 B.n784 B.n37 10.6151
R1268 B.n784 B.n783 10.6151
R1269 B.n783 B.n782 10.6151
R1270 B.n111 B.n45 10.6151
R1271 B.n114 B.n111 10.6151
R1272 B.n115 B.n114 10.6151
R1273 B.n118 B.n115 10.6151
R1274 B.n119 B.n118 10.6151
R1275 B.n122 B.n119 10.6151
R1276 B.n123 B.n122 10.6151
R1277 B.n126 B.n123 10.6151
R1278 B.n127 B.n126 10.6151
R1279 B.n130 B.n127 10.6151
R1280 B.n131 B.n130 10.6151
R1281 B.n134 B.n131 10.6151
R1282 B.n135 B.n134 10.6151
R1283 B.n138 B.n135 10.6151
R1284 B.n139 B.n138 10.6151
R1285 B.n142 B.n139 10.6151
R1286 B.n143 B.n142 10.6151
R1287 B.n146 B.n143 10.6151
R1288 B.n147 B.n146 10.6151
R1289 B.n150 B.n147 10.6151
R1290 B.n151 B.n150 10.6151
R1291 B.n154 B.n151 10.6151
R1292 B.n155 B.n154 10.6151
R1293 B.n158 B.n155 10.6151
R1294 B.n159 B.n158 10.6151
R1295 B.n162 B.n159 10.6151
R1296 B.n163 B.n162 10.6151
R1297 B.n166 B.n163 10.6151
R1298 B.n167 B.n166 10.6151
R1299 B.n170 B.n167 10.6151
R1300 B.n171 B.n170 10.6151
R1301 B.n174 B.n171 10.6151
R1302 B.n175 B.n174 10.6151
R1303 B.n178 B.n175 10.6151
R1304 B.n179 B.n178 10.6151
R1305 B.n182 B.n179 10.6151
R1306 B.n183 B.n182 10.6151
R1307 B.n186 B.n183 10.6151
R1308 B.n187 B.n186 10.6151
R1309 B.n190 B.n187 10.6151
R1310 B.n191 B.n190 10.6151
R1311 B.n194 B.n191 10.6151
R1312 B.n195 B.n194 10.6151
R1313 B.n198 B.n195 10.6151
R1314 B.n199 B.n198 10.6151
R1315 B.n202 B.n199 10.6151
R1316 B.n203 B.n202 10.6151
R1317 B.n206 B.n203 10.6151
R1318 B.n207 B.n206 10.6151
R1319 B.n210 B.n207 10.6151
R1320 B.n211 B.n210 10.6151
R1321 B.n215 B.n214 10.6151
R1322 B.n218 B.n215 10.6151
R1323 B.n219 B.n218 10.6151
R1324 B.n222 B.n219 10.6151
R1325 B.n223 B.n222 10.6151
R1326 B.n226 B.n223 10.6151
R1327 B.n227 B.n226 10.6151
R1328 B.n230 B.n227 10.6151
R1329 B.n231 B.n230 10.6151
R1330 B.n235 B.n234 10.6151
R1331 B.n238 B.n235 10.6151
R1332 B.n239 B.n238 10.6151
R1333 B.n242 B.n239 10.6151
R1334 B.n243 B.n242 10.6151
R1335 B.n246 B.n243 10.6151
R1336 B.n247 B.n246 10.6151
R1337 B.n250 B.n247 10.6151
R1338 B.n251 B.n250 10.6151
R1339 B.n254 B.n251 10.6151
R1340 B.n255 B.n254 10.6151
R1341 B.n258 B.n255 10.6151
R1342 B.n259 B.n258 10.6151
R1343 B.n262 B.n259 10.6151
R1344 B.n263 B.n262 10.6151
R1345 B.n266 B.n263 10.6151
R1346 B.n267 B.n266 10.6151
R1347 B.n270 B.n267 10.6151
R1348 B.n271 B.n270 10.6151
R1349 B.n274 B.n271 10.6151
R1350 B.n275 B.n274 10.6151
R1351 B.n278 B.n275 10.6151
R1352 B.n279 B.n278 10.6151
R1353 B.n282 B.n279 10.6151
R1354 B.n283 B.n282 10.6151
R1355 B.n286 B.n283 10.6151
R1356 B.n287 B.n286 10.6151
R1357 B.n290 B.n287 10.6151
R1358 B.n291 B.n290 10.6151
R1359 B.n294 B.n291 10.6151
R1360 B.n295 B.n294 10.6151
R1361 B.n298 B.n295 10.6151
R1362 B.n299 B.n298 10.6151
R1363 B.n302 B.n299 10.6151
R1364 B.n303 B.n302 10.6151
R1365 B.n306 B.n303 10.6151
R1366 B.n307 B.n306 10.6151
R1367 B.n310 B.n307 10.6151
R1368 B.n311 B.n310 10.6151
R1369 B.n314 B.n311 10.6151
R1370 B.n315 B.n314 10.6151
R1371 B.n318 B.n315 10.6151
R1372 B.n319 B.n318 10.6151
R1373 B.n322 B.n319 10.6151
R1374 B.n323 B.n322 10.6151
R1375 B.n326 B.n323 10.6151
R1376 B.n327 B.n326 10.6151
R1377 B.n330 B.n327 10.6151
R1378 B.n332 B.n330 10.6151
R1379 B.n333 B.n332 10.6151
R1380 B.n776 B.n333 10.6151
R1381 B.n542 B.n541 9.36635
R1382 B.n562 B.n406 9.36635
R1383 B.n211 B.n110 9.36635
R1384 B.n234 B.n107 9.36635
R1385 B.n832 B.n0 8.11757
R1386 B.n832 B.n1 8.11757
R1387 B.n682 B.t6 6.34818
R1388 B.t0 B.n336 6.34818
R1389 B.n747 B.t3 6.34818
R1390 B.n39 B.t10 6.34818
R1391 B.n543 B.n542 1.24928
R1392 B.n563 B.n562 1.24928
R1393 B.n214 B.n110 1.24928
R1394 B.n231 B.n107 1.24928
R1395 VP.n3 VP.t4 405.647
R1396 VP.n8 VP.t1 382.7
R1397 VP.n14 VP.t0 382.7
R1398 VP.n6 VP.t2 382.7
R1399 VP.n12 VP.t5 346.327
R1400 VP.n4 VP.t3 346.327
R1401 VP.n5 VP.n2 161.3
R1402 VP.n13 VP.n0 161.3
R1403 VP.n12 VP.n11 161.3
R1404 VP.n10 VP.n1 161.3
R1405 VP.n7 VP.n6 80.6037
R1406 VP.n15 VP.n14 80.6037
R1407 VP.n9 VP.n8 80.6037
R1408 VP.n8 VP.n1 50.1678
R1409 VP.n14 VP.n13 50.1678
R1410 VP.n6 VP.n5 50.1678
R1411 VP.n9 VP.n7 45.5506
R1412 VP.n4 VP.n3 32.6313
R1413 VP.n3 VP.n2 28.168
R1414 VP.n12 VP.n1 24.5923
R1415 VP.n13 VP.n12 24.5923
R1416 VP.n5 VP.n4 24.5923
R1417 VP.n7 VP.n2 0.285035
R1418 VP.n10 VP.n9 0.285035
R1419 VP.n15 VP.n0 0.285035
R1420 VP.n11 VP.n10 0.189894
R1421 VP.n11 VP.n0 0.189894
R1422 VP VP.n15 0.146778
R1423 VTAIL.n346 VTAIL.n266 289.615
R1424 VTAIL.n82 VTAIL.n2 289.615
R1425 VTAIL.n260 VTAIL.n180 289.615
R1426 VTAIL.n172 VTAIL.n92 289.615
R1427 VTAIL.n295 VTAIL.n294 185
R1428 VTAIL.n297 VTAIL.n296 185
R1429 VTAIL.n290 VTAIL.n289 185
R1430 VTAIL.n303 VTAIL.n302 185
R1431 VTAIL.n305 VTAIL.n304 185
R1432 VTAIL.n286 VTAIL.n285 185
R1433 VTAIL.n311 VTAIL.n310 185
R1434 VTAIL.n313 VTAIL.n312 185
R1435 VTAIL.n282 VTAIL.n281 185
R1436 VTAIL.n319 VTAIL.n318 185
R1437 VTAIL.n321 VTAIL.n320 185
R1438 VTAIL.n278 VTAIL.n277 185
R1439 VTAIL.n327 VTAIL.n326 185
R1440 VTAIL.n329 VTAIL.n328 185
R1441 VTAIL.n274 VTAIL.n273 185
R1442 VTAIL.n336 VTAIL.n335 185
R1443 VTAIL.n337 VTAIL.n272 185
R1444 VTAIL.n339 VTAIL.n338 185
R1445 VTAIL.n270 VTAIL.n269 185
R1446 VTAIL.n345 VTAIL.n344 185
R1447 VTAIL.n347 VTAIL.n346 185
R1448 VTAIL.n31 VTAIL.n30 185
R1449 VTAIL.n33 VTAIL.n32 185
R1450 VTAIL.n26 VTAIL.n25 185
R1451 VTAIL.n39 VTAIL.n38 185
R1452 VTAIL.n41 VTAIL.n40 185
R1453 VTAIL.n22 VTAIL.n21 185
R1454 VTAIL.n47 VTAIL.n46 185
R1455 VTAIL.n49 VTAIL.n48 185
R1456 VTAIL.n18 VTAIL.n17 185
R1457 VTAIL.n55 VTAIL.n54 185
R1458 VTAIL.n57 VTAIL.n56 185
R1459 VTAIL.n14 VTAIL.n13 185
R1460 VTAIL.n63 VTAIL.n62 185
R1461 VTAIL.n65 VTAIL.n64 185
R1462 VTAIL.n10 VTAIL.n9 185
R1463 VTAIL.n72 VTAIL.n71 185
R1464 VTAIL.n73 VTAIL.n8 185
R1465 VTAIL.n75 VTAIL.n74 185
R1466 VTAIL.n6 VTAIL.n5 185
R1467 VTAIL.n81 VTAIL.n80 185
R1468 VTAIL.n83 VTAIL.n82 185
R1469 VTAIL.n261 VTAIL.n260 185
R1470 VTAIL.n259 VTAIL.n258 185
R1471 VTAIL.n184 VTAIL.n183 185
R1472 VTAIL.n188 VTAIL.n186 185
R1473 VTAIL.n253 VTAIL.n252 185
R1474 VTAIL.n251 VTAIL.n250 185
R1475 VTAIL.n190 VTAIL.n189 185
R1476 VTAIL.n245 VTAIL.n244 185
R1477 VTAIL.n243 VTAIL.n242 185
R1478 VTAIL.n194 VTAIL.n193 185
R1479 VTAIL.n237 VTAIL.n236 185
R1480 VTAIL.n235 VTAIL.n234 185
R1481 VTAIL.n198 VTAIL.n197 185
R1482 VTAIL.n229 VTAIL.n228 185
R1483 VTAIL.n227 VTAIL.n226 185
R1484 VTAIL.n202 VTAIL.n201 185
R1485 VTAIL.n221 VTAIL.n220 185
R1486 VTAIL.n219 VTAIL.n218 185
R1487 VTAIL.n206 VTAIL.n205 185
R1488 VTAIL.n213 VTAIL.n212 185
R1489 VTAIL.n211 VTAIL.n210 185
R1490 VTAIL.n173 VTAIL.n172 185
R1491 VTAIL.n171 VTAIL.n170 185
R1492 VTAIL.n96 VTAIL.n95 185
R1493 VTAIL.n100 VTAIL.n98 185
R1494 VTAIL.n165 VTAIL.n164 185
R1495 VTAIL.n163 VTAIL.n162 185
R1496 VTAIL.n102 VTAIL.n101 185
R1497 VTAIL.n157 VTAIL.n156 185
R1498 VTAIL.n155 VTAIL.n154 185
R1499 VTAIL.n106 VTAIL.n105 185
R1500 VTAIL.n149 VTAIL.n148 185
R1501 VTAIL.n147 VTAIL.n146 185
R1502 VTAIL.n110 VTAIL.n109 185
R1503 VTAIL.n141 VTAIL.n140 185
R1504 VTAIL.n139 VTAIL.n138 185
R1505 VTAIL.n114 VTAIL.n113 185
R1506 VTAIL.n133 VTAIL.n132 185
R1507 VTAIL.n131 VTAIL.n130 185
R1508 VTAIL.n118 VTAIL.n117 185
R1509 VTAIL.n125 VTAIL.n124 185
R1510 VTAIL.n123 VTAIL.n122 185
R1511 VTAIL.n293 VTAIL.t0 147.659
R1512 VTAIL.n29 VTAIL.t3 147.659
R1513 VTAIL.n209 VTAIL.t5 147.659
R1514 VTAIL.n121 VTAIL.t1 147.659
R1515 VTAIL.n296 VTAIL.n295 104.615
R1516 VTAIL.n296 VTAIL.n289 104.615
R1517 VTAIL.n303 VTAIL.n289 104.615
R1518 VTAIL.n304 VTAIL.n303 104.615
R1519 VTAIL.n304 VTAIL.n285 104.615
R1520 VTAIL.n311 VTAIL.n285 104.615
R1521 VTAIL.n312 VTAIL.n311 104.615
R1522 VTAIL.n312 VTAIL.n281 104.615
R1523 VTAIL.n319 VTAIL.n281 104.615
R1524 VTAIL.n320 VTAIL.n319 104.615
R1525 VTAIL.n320 VTAIL.n277 104.615
R1526 VTAIL.n327 VTAIL.n277 104.615
R1527 VTAIL.n328 VTAIL.n327 104.615
R1528 VTAIL.n328 VTAIL.n273 104.615
R1529 VTAIL.n336 VTAIL.n273 104.615
R1530 VTAIL.n337 VTAIL.n336 104.615
R1531 VTAIL.n338 VTAIL.n337 104.615
R1532 VTAIL.n338 VTAIL.n269 104.615
R1533 VTAIL.n345 VTAIL.n269 104.615
R1534 VTAIL.n346 VTAIL.n345 104.615
R1535 VTAIL.n32 VTAIL.n31 104.615
R1536 VTAIL.n32 VTAIL.n25 104.615
R1537 VTAIL.n39 VTAIL.n25 104.615
R1538 VTAIL.n40 VTAIL.n39 104.615
R1539 VTAIL.n40 VTAIL.n21 104.615
R1540 VTAIL.n47 VTAIL.n21 104.615
R1541 VTAIL.n48 VTAIL.n47 104.615
R1542 VTAIL.n48 VTAIL.n17 104.615
R1543 VTAIL.n55 VTAIL.n17 104.615
R1544 VTAIL.n56 VTAIL.n55 104.615
R1545 VTAIL.n56 VTAIL.n13 104.615
R1546 VTAIL.n63 VTAIL.n13 104.615
R1547 VTAIL.n64 VTAIL.n63 104.615
R1548 VTAIL.n64 VTAIL.n9 104.615
R1549 VTAIL.n72 VTAIL.n9 104.615
R1550 VTAIL.n73 VTAIL.n72 104.615
R1551 VTAIL.n74 VTAIL.n73 104.615
R1552 VTAIL.n74 VTAIL.n5 104.615
R1553 VTAIL.n81 VTAIL.n5 104.615
R1554 VTAIL.n82 VTAIL.n81 104.615
R1555 VTAIL.n260 VTAIL.n259 104.615
R1556 VTAIL.n259 VTAIL.n183 104.615
R1557 VTAIL.n188 VTAIL.n183 104.615
R1558 VTAIL.n252 VTAIL.n188 104.615
R1559 VTAIL.n252 VTAIL.n251 104.615
R1560 VTAIL.n251 VTAIL.n189 104.615
R1561 VTAIL.n244 VTAIL.n189 104.615
R1562 VTAIL.n244 VTAIL.n243 104.615
R1563 VTAIL.n243 VTAIL.n193 104.615
R1564 VTAIL.n236 VTAIL.n193 104.615
R1565 VTAIL.n236 VTAIL.n235 104.615
R1566 VTAIL.n235 VTAIL.n197 104.615
R1567 VTAIL.n228 VTAIL.n197 104.615
R1568 VTAIL.n228 VTAIL.n227 104.615
R1569 VTAIL.n227 VTAIL.n201 104.615
R1570 VTAIL.n220 VTAIL.n201 104.615
R1571 VTAIL.n220 VTAIL.n219 104.615
R1572 VTAIL.n219 VTAIL.n205 104.615
R1573 VTAIL.n212 VTAIL.n205 104.615
R1574 VTAIL.n212 VTAIL.n211 104.615
R1575 VTAIL.n172 VTAIL.n171 104.615
R1576 VTAIL.n171 VTAIL.n95 104.615
R1577 VTAIL.n100 VTAIL.n95 104.615
R1578 VTAIL.n164 VTAIL.n100 104.615
R1579 VTAIL.n164 VTAIL.n163 104.615
R1580 VTAIL.n163 VTAIL.n101 104.615
R1581 VTAIL.n156 VTAIL.n101 104.615
R1582 VTAIL.n156 VTAIL.n155 104.615
R1583 VTAIL.n155 VTAIL.n105 104.615
R1584 VTAIL.n148 VTAIL.n105 104.615
R1585 VTAIL.n148 VTAIL.n147 104.615
R1586 VTAIL.n147 VTAIL.n109 104.615
R1587 VTAIL.n140 VTAIL.n109 104.615
R1588 VTAIL.n140 VTAIL.n139 104.615
R1589 VTAIL.n139 VTAIL.n113 104.615
R1590 VTAIL.n132 VTAIL.n113 104.615
R1591 VTAIL.n132 VTAIL.n131 104.615
R1592 VTAIL.n131 VTAIL.n117 104.615
R1593 VTAIL.n124 VTAIL.n117 104.615
R1594 VTAIL.n124 VTAIL.n123 104.615
R1595 VTAIL.n295 VTAIL.t0 52.3082
R1596 VTAIL.n31 VTAIL.t3 52.3082
R1597 VTAIL.n211 VTAIL.t5 52.3082
R1598 VTAIL.n123 VTAIL.t1 52.3082
R1599 VTAIL.n179 VTAIL.n178 47.2668
R1600 VTAIL.n91 VTAIL.n90 47.2668
R1601 VTAIL.n1 VTAIL.n0 47.2666
R1602 VTAIL.n89 VTAIL.n88 47.2666
R1603 VTAIL.n351 VTAIL.n350 35.2884
R1604 VTAIL.n87 VTAIL.n86 35.2884
R1605 VTAIL.n265 VTAIL.n264 35.2884
R1606 VTAIL.n177 VTAIL.n176 35.2884
R1607 VTAIL.n91 VTAIL.n89 28.1772
R1608 VTAIL.n351 VTAIL.n265 26.9617
R1609 VTAIL.n294 VTAIL.n293 15.6677
R1610 VTAIL.n30 VTAIL.n29 15.6677
R1611 VTAIL.n210 VTAIL.n209 15.6677
R1612 VTAIL.n122 VTAIL.n121 15.6677
R1613 VTAIL.n339 VTAIL.n270 13.1884
R1614 VTAIL.n75 VTAIL.n6 13.1884
R1615 VTAIL.n186 VTAIL.n184 13.1884
R1616 VTAIL.n98 VTAIL.n96 13.1884
R1617 VTAIL.n297 VTAIL.n292 12.8005
R1618 VTAIL.n340 VTAIL.n272 12.8005
R1619 VTAIL.n344 VTAIL.n343 12.8005
R1620 VTAIL.n33 VTAIL.n28 12.8005
R1621 VTAIL.n76 VTAIL.n8 12.8005
R1622 VTAIL.n80 VTAIL.n79 12.8005
R1623 VTAIL.n258 VTAIL.n257 12.8005
R1624 VTAIL.n254 VTAIL.n253 12.8005
R1625 VTAIL.n213 VTAIL.n208 12.8005
R1626 VTAIL.n170 VTAIL.n169 12.8005
R1627 VTAIL.n166 VTAIL.n165 12.8005
R1628 VTAIL.n125 VTAIL.n120 12.8005
R1629 VTAIL.n298 VTAIL.n290 12.0247
R1630 VTAIL.n335 VTAIL.n334 12.0247
R1631 VTAIL.n347 VTAIL.n268 12.0247
R1632 VTAIL.n34 VTAIL.n26 12.0247
R1633 VTAIL.n71 VTAIL.n70 12.0247
R1634 VTAIL.n83 VTAIL.n4 12.0247
R1635 VTAIL.n261 VTAIL.n182 12.0247
R1636 VTAIL.n250 VTAIL.n187 12.0247
R1637 VTAIL.n214 VTAIL.n206 12.0247
R1638 VTAIL.n173 VTAIL.n94 12.0247
R1639 VTAIL.n162 VTAIL.n99 12.0247
R1640 VTAIL.n126 VTAIL.n118 12.0247
R1641 VTAIL.n302 VTAIL.n301 11.249
R1642 VTAIL.n333 VTAIL.n274 11.249
R1643 VTAIL.n348 VTAIL.n266 11.249
R1644 VTAIL.n38 VTAIL.n37 11.249
R1645 VTAIL.n69 VTAIL.n10 11.249
R1646 VTAIL.n84 VTAIL.n2 11.249
R1647 VTAIL.n262 VTAIL.n180 11.249
R1648 VTAIL.n249 VTAIL.n190 11.249
R1649 VTAIL.n218 VTAIL.n217 11.249
R1650 VTAIL.n174 VTAIL.n92 11.249
R1651 VTAIL.n161 VTAIL.n102 11.249
R1652 VTAIL.n130 VTAIL.n129 11.249
R1653 VTAIL.n305 VTAIL.n288 10.4732
R1654 VTAIL.n330 VTAIL.n329 10.4732
R1655 VTAIL.n41 VTAIL.n24 10.4732
R1656 VTAIL.n66 VTAIL.n65 10.4732
R1657 VTAIL.n246 VTAIL.n245 10.4732
R1658 VTAIL.n221 VTAIL.n204 10.4732
R1659 VTAIL.n158 VTAIL.n157 10.4732
R1660 VTAIL.n133 VTAIL.n116 10.4732
R1661 VTAIL.n306 VTAIL.n286 9.69747
R1662 VTAIL.n326 VTAIL.n276 9.69747
R1663 VTAIL.n42 VTAIL.n22 9.69747
R1664 VTAIL.n62 VTAIL.n12 9.69747
R1665 VTAIL.n242 VTAIL.n192 9.69747
R1666 VTAIL.n222 VTAIL.n202 9.69747
R1667 VTAIL.n154 VTAIL.n104 9.69747
R1668 VTAIL.n134 VTAIL.n114 9.69747
R1669 VTAIL.n350 VTAIL.n349 9.45567
R1670 VTAIL.n86 VTAIL.n85 9.45567
R1671 VTAIL.n264 VTAIL.n263 9.45567
R1672 VTAIL.n176 VTAIL.n175 9.45567
R1673 VTAIL.n349 VTAIL.n348 9.3005
R1674 VTAIL.n268 VTAIL.n267 9.3005
R1675 VTAIL.n343 VTAIL.n342 9.3005
R1676 VTAIL.n315 VTAIL.n314 9.3005
R1677 VTAIL.n284 VTAIL.n283 9.3005
R1678 VTAIL.n309 VTAIL.n308 9.3005
R1679 VTAIL.n307 VTAIL.n306 9.3005
R1680 VTAIL.n288 VTAIL.n287 9.3005
R1681 VTAIL.n301 VTAIL.n300 9.3005
R1682 VTAIL.n299 VTAIL.n298 9.3005
R1683 VTAIL.n292 VTAIL.n291 9.3005
R1684 VTAIL.n317 VTAIL.n316 9.3005
R1685 VTAIL.n280 VTAIL.n279 9.3005
R1686 VTAIL.n323 VTAIL.n322 9.3005
R1687 VTAIL.n325 VTAIL.n324 9.3005
R1688 VTAIL.n276 VTAIL.n275 9.3005
R1689 VTAIL.n331 VTAIL.n330 9.3005
R1690 VTAIL.n333 VTAIL.n332 9.3005
R1691 VTAIL.n334 VTAIL.n271 9.3005
R1692 VTAIL.n341 VTAIL.n340 9.3005
R1693 VTAIL.n85 VTAIL.n84 9.3005
R1694 VTAIL.n4 VTAIL.n3 9.3005
R1695 VTAIL.n79 VTAIL.n78 9.3005
R1696 VTAIL.n51 VTAIL.n50 9.3005
R1697 VTAIL.n20 VTAIL.n19 9.3005
R1698 VTAIL.n45 VTAIL.n44 9.3005
R1699 VTAIL.n43 VTAIL.n42 9.3005
R1700 VTAIL.n24 VTAIL.n23 9.3005
R1701 VTAIL.n37 VTAIL.n36 9.3005
R1702 VTAIL.n35 VTAIL.n34 9.3005
R1703 VTAIL.n28 VTAIL.n27 9.3005
R1704 VTAIL.n53 VTAIL.n52 9.3005
R1705 VTAIL.n16 VTAIL.n15 9.3005
R1706 VTAIL.n59 VTAIL.n58 9.3005
R1707 VTAIL.n61 VTAIL.n60 9.3005
R1708 VTAIL.n12 VTAIL.n11 9.3005
R1709 VTAIL.n67 VTAIL.n66 9.3005
R1710 VTAIL.n69 VTAIL.n68 9.3005
R1711 VTAIL.n70 VTAIL.n7 9.3005
R1712 VTAIL.n77 VTAIL.n76 9.3005
R1713 VTAIL.n196 VTAIL.n195 9.3005
R1714 VTAIL.n239 VTAIL.n238 9.3005
R1715 VTAIL.n241 VTAIL.n240 9.3005
R1716 VTAIL.n192 VTAIL.n191 9.3005
R1717 VTAIL.n247 VTAIL.n246 9.3005
R1718 VTAIL.n249 VTAIL.n248 9.3005
R1719 VTAIL.n187 VTAIL.n185 9.3005
R1720 VTAIL.n255 VTAIL.n254 9.3005
R1721 VTAIL.n263 VTAIL.n262 9.3005
R1722 VTAIL.n182 VTAIL.n181 9.3005
R1723 VTAIL.n257 VTAIL.n256 9.3005
R1724 VTAIL.n233 VTAIL.n232 9.3005
R1725 VTAIL.n231 VTAIL.n230 9.3005
R1726 VTAIL.n200 VTAIL.n199 9.3005
R1727 VTAIL.n225 VTAIL.n224 9.3005
R1728 VTAIL.n223 VTAIL.n222 9.3005
R1729 VTAIL.n204 VTAIL.n203 9.3005
R1730 VTAIL.n217 VTAIL.n216 9.3005
R1731 VTAIL.n215 VTAIL.n214 9.3005
R1732 VTAIL.n208 VTAIL.n207 9.3005
R1733 VTAIL.n108 VTAIL.n107 9.3005
R1734 VTAIL.n151 VTAIL.n150 9.3005
R1735 VTAIL.n153 VTAIL.n152 9.3005
R1736 VTAIL.n104 VTAIL.n103 9.3005
R1737 VTAIL.n159 VTAIL.n158 9.3005
R1738 VTAIL.n161 VTAIL.n160 9.3005
R1739 VTAIL.n99 VTAIL.n97 9.3005
R1740 VTAIL.n167 VTAIL.n166 9.3005
R1741 VTAIL.n175 VTAIL.n174 9.3005
R1742 VTAIL.n94 VTAIL.n93 9.3005
R1743 VTAIL.n169 VTAIL.n168 9.3005
R1744 VTAIL.n145 VTAIL.n144 9.3005
R1745 VTAIL.n143 VTAIL.n142 9.3005
R1746 VTAIL.n112 VTAIL.n111 9.3005
R1747 VTAIL.n137 VTAIL.n136 9.3005
R1748 VTAIL.n135 VTAIL.n134 9.3005
R1749 VTAIL.n116 VTAIL.n115 9.3005
R1750 VTAIL.n129 VTAIL.n128 9.3005
R1751 VTAIL.n127 VTAIL.n126 9.3005
R1752 VTAIL.n120 VTAIL.n119 9.3005
R1753 VTAIL.n310 VTAIL.n309 8.92171
R1754 VTAIL.n325 VTAIL.n278 8.92171
R1755 VTAIL.n46 VTAIL.n45 8.92171
R1756 VTAIL.n61 VTAIL.n14 8.92171
R1757 VTAIL.n241 VTAIL.n194 8.92171
R1758 VTAIL.n226 VTAIL.n225 8.92171
R1759 VTAIL.n153 VTAIL.n106 8.92171
R1760 VTAIL.n138 VTAIL.n137 8.92171
R1761 VTAIL.n313 VTAIL.n284 8.14595
R1762 VTAIL.n322 VTAIL.n321 8.14595
R1763 VTAIL.n49 VTAIL.n20 8.14595
R1764 VTAIL.n58 VTAIL.n57 8.14595
R1765 VTAIL.n238 VTAIL.n237 8.14595
R1766 VTAIL.n229 VTAIL.n200 8.14595
R1767 VTAIL.n150 VTAIL.n149 8.14595
R1768 VTAIL.n141 VTAIL.n112 8.14595
R1769 VTAIL.n314 VTAIL.n282 7.3702
R1770 VTAIL.n318 VTAIL.n280 7.3702
R1771 VTAIL.n50 VTAIL.n18 7.3702
R1772 VTAIL.n54 VTAIL.n16 7.3702
R1773 VTAIL.n234 VTAIL.n196 7.3702
R1774 VTAIL.n230 VTAIL.n198 7.3702
R1775 VTAIL.n146 VTAIL.n108 7.3702
R1776 VTAIL.n142 VTAIL.n110 7.3702
R1777 VTAIL.n317 VTAIL.n282 6.59444
R1778 VTAIL.n318 VTAIL.n317 6.59444
R1779 VTAIL.n53 VTAIL.n18 6.59444
R1780 VTAIL.n54 VTAIL.n53 6.59444
R1781 VTAIL.n234 VTAIL.n233 6.59444
R1782 VTAIL.n233 VTAIL.n198 6.59444
R1783 VTAIL.n146 VTAIL.n145 6.59444
R1784 VTAIL.n145 VTAIL.n110 6.59444
R1785 VTAIL.n314 VTAIL.n313 5.81868
R1786 VTAIL.n321 VTAIL.n280 5.81868
R1787 VTAIL.n50 VTAIL.n49 5.81868
R1788 VTAIL.n57 VTAIL.n16 5.81868
R1789 VTAIL.n237 VTAIL.n196 5.81868
R1790 VTAIL.n230 VTAIL.n229 5.81868
R1791 VTAIL.n149 VTAIL.n108 5.81868
R1792 VTAIL.n142 VTAIL.n141 5.81868
R1793 VTAIL.n310 VTAIL.n284 5.04292
R1794 VTAIL.n322 VTAIL.n278 5.04292
R1795 VTAIL.n46 VTAIL.n20 5.04292
R1796 VTAIL.n58 VTAIL.n14 5.04292
R1797 VTAIL.n238 VTAIL.n194 5.04292
R1798 VTAIL.n226 VTAIL.n200 5.04292
R1799 VTAIL.n150 VTAIL.n106 5.04292
R1800 VTAIL.n138 VTAIL.n112 5.04292
R1801 VTAIL.n293 VTAIL.n291 4.38563
R1802 VTAIL.n29 VTAIL.n27 4.38563
R1803 VTAIL.n209 VTAIL.n207 4.38563
R1804 VTAIL.n121 VTAIL.n119 4.38563
R1805 VTAIL.n309 VTAIL.n286 4.26717
R1806 VTAIL.n326 VTAIL.n325 4.26717
R1807 VTAIL.n45 VTAIL.n22 4.26717
R1808 VTAIL.n62 VTAIL.n61 4.26717
R1809 VTAIL.n242 VTAIL.n241 4.26717
R1810 VTAIL.n225 VTAIL.n202 4.26717
R1811 VTAIL.n154 VTAIL.n153 4.26717
R1812 VTAIL.n137 VTAIL.n114 4.26717
R1813 VTAIL.n306 VTAIL.n305 3.49141
R1814 VTAIL.n329 VTAIL.n276 3.49141
R1815 VTAIL.n42 VTAIL.n41 3.49141
R1816 VTAIL.n65 VTAIL.n12 3.49141
R1817 VTAIL.n245 VTAIL.n192 3.49141
R1818 VTAIL.n222 VTAIL.n221 3.49141
R1819 VTAIL.n157 VTAIL.n104 3.49141
R1820 VTAIL.n134 VTAIL.n133 3.49141
R1821 VTAIL.n302 VTAIL.n288 2.71565
R1822 VTAIL.n330 VTAIL.n274 2.71565
R1823 VTAIL.n350 VTAIL.n266 2.71565
R1824 VTAIL.n38 VTAIL.n24 2.71565
R1825 VTAIL.n66 VTAIL.n10 2.71565
R1826 VTAIL.n86 VTAIL.n2 2.71565
R1827 VTAIL.n264 VTAIL.n180 2.71565
R1828 VTAIL.n246 VTAIL.n190 2.71565
R1829 VTAIL.n218 VTAIL.n204 2.71565
R1830 VTAIL.n176 VTAIL.n92 2.71565
R1831 VTAIL.n158 VTAIL.n102 2.71565
R1832 VTAIL.n130 VTAIL.n116 2.71565
R1833 VTAIL.n301 VTAIL.n290 1.93989
R1834 VTAIL.n335 VTAIL.n333 1.93989
R1835 VTAIL.n348 VTAIL.n347 1.93989
R1836 VTAIL.n37 VTAIL.n26 1.93989
R1837 VTAIL.n71 VTAIL.n69 1.93989
R1838 VTAIL.n84 VTAIL.n83 1.93989
R1839 VTAIL.n262 VTAIL.n261 1.93989
R1840 VTAIL.n250 VTAIL.n249 1.93989
R1841 VTAIL.n217 VTAIL.n206 1.93989
R1842 VTAIL.n174 VTAIL.n173 1.93989
R1843 VTAIL.n162 VTAIL.n161 1.93989
R1844 VTAIL.n129 VTAIL.n118 1.93989
R1845 VTAIL.n0 VTAIL.t10 1.27627
R1846 VTAIL.n0 VTAIL.t2 1.27627
R1847 VTAIL.n88 VTAIL.t7 1.27627
R1848 VTAIL.n88 VTAIL.t6 1.27627
R1849 VTAIL.n178 VTAIL.t8 1.27627
R1850 VTAIL.n178 VTAIL.t4 1.27627
R1851 VTAIL.n90 VTAIL.t9 1.27627
R1852 VTAIL.n90 VTAIL.t11 1.27627
R1853 VTAIL.n177 VTAIL.n91 1.21602
R1854 VTAIL.n265 VTAIL.n179 1.21602
R1855 VTAIL.n89 VTAIL.n87 1.21602
R1856 VTAIL.n298 VTAIL.n297 1.16414
R1857 VTAIL.n334 VTAIL.n272 1.16414
R1858 VTAIL.n344 VTAIL.n268 1.16414
R1859 VTAIL.n34 VTAIL.n33 1.16414
R1860 VTAIL.n70 VTAIL.n8 1.16414
R1861 VTAIL.n80 VTAIL.n4 1.16414
R1862 VTAIL.n258 VTAIL.n182 1.16414
R1863 VTAIL.n253 VTAIL.n187 1.16414
R1864 VTAIL.n214 VTAIL.n213 1.16414
R1865 VTAIL.n170 VTAIL.n94 1.16414
R1866 VTAIL.n165 VTAIL.n99 1.16414
R1867 VTAIL.n126 VTAIL.n125 1.16414
R1868 VTAIL.n179 VTAIL.n177 1.07809
R1869 VTAIL.n87 VTAIL.n1 1.07809
R1870 VTAIL VTAIL.n351 0.853948
R1871 VTAIL.n294 VTAIL.n292 0.388379
R1872 VTAIL.n340 VTAIL.n339 0.388379
R1873 VTAIL.n343 VTAIL.n270 0.388379
R1874 VTAIL.n30 VTAIL.n28 0.388379
R1875 VTAIL.n76 VTAIL.n75 0.388379
R1876 VTAIL.n79 VTAIL.n6 0.388379
R1877 VTAIL.n257 VTAIL.n184 0.388379
R1878 VTAIL.n254 VTAIL.n186 0.388379
R1879 VTAIL.n210 VTAIL.n208 0.388379
R1880 VTAIL.n169 VTAIL.n96 0.388379
R1881 VTAIL.n166 VTAIL.n98 0.388379
R1882 VTAIL.n122 VTAIL.n120 0.388379
R1883 VTAIL VTAIL.n1 0.362569
R1884 VTAIL.n299 VTAIL.n291 0.155672
R1885 VTAIL.n300 VTAIL.n299 0.155672
R1886 VTAIL.n300 VTAIL.n287 0.155672
R1887 VTAIL.n307 VTAIL.n287 0.155672
R1888 VTAIL.n308 VTAIL.n307 0.155672
R1889 VTAIL.n308 VTAIL.n283 0.155672
R1890 VTAIL.n315 VTAIL.n283 0.155672
R1891 VTAIL.n316 VTAIL.n315 0.155672
R1892 VTAIL.n316 VTAIL.n279 0.155672
R1893 VTAIL.n323 VTAIL.n279 0.155672
R1894 VTAIL.n324 VTAIL.n323 0.155672
R1895 VTAIL.n324 VTAIL.n275 0.155672
R1896 VTAIL.n331 VTAIL.n275 0.155672
R1897 VTAIL.n332 VTAIL.n331 0.155672
R1898 VTAIL.n332 VTAIL.n271 0.155672
R1899 VTAIL.n341 VTAIL.n271 0.155672
R1900 VTAIL.n342 VTAIL.n341 0.155672
R1901 VTAIL.n342 VTAIL.n267 0.155672
R1902 VTAIL.n349 VTAIL.n267 0.155672
R1903 VTAIL.n35 VTAIL.n27 0.155672
R1904 VTAIL.n36 VTAIL.n35 0.155672
R1905 VTAIL.n36 VTAIL.n23 0.155672
R1906 VTAIL.n43 VTAIL.n23 0.155672
R1907 VTAIL.n44 VTAIL.n43 0.155672
R1908 VTAIL.n44 VTAIL.n19 0.155672
R1909 VTAIL.n51 VTAIL.n19 0.155672
R1910 VTAIL.n52 VTAIL.n51 0.155672
R1911 VTAIL.n52 VTAIL.n15 0.155672
R1912 VTAIL.n59 VTAIL.n15 0.155672
R1913 VTAIL.n60 VTAIL.n59 0.155672
R1914 VTAIL.n60 VTAIL.n11 0.155672
R1915 VTAIL.n67 VTAIL.n11 0.155672
R1916 VTAIL.n68 VTAIL.n67 0.155672
R1917 VTAIL.n68 VTAIL.n7 0.155672
R1918 VTAIL.n77 VTAIL.n7 0.155672
R1919 VTAIL.n78 VTAIL.n77 0.155672
R1920 VTAIL.n78 VTAIL.n3 0.155672
R1921 VTAIL.n85 VTAIL.n3 0.155672
R1922 VTAIL.n263 VTAIL.n181 0.155672
R1923 VTAIL.n256 VTAIL.n181 0.155672
R1924 VTAIL.n256 VTAIL.n255 0.155672
R1925 VTAIL.n255 VTAIL.n185 0.155672
R1926 VTAIL.n248 VTAIL.n185 0.155672
R1927 VTAIL.n248 VTAIL.n247 0.155672
R1928 VTAIL.n247 VTAIL.n191 0.155672
R1929 VTAIL.n240 VTAIL.n191 0.155672
R1930 VTAIL.n240 VTAIL.n239 0.155672
R1931 VTAIL.n239 VTAIL.n195 0.155672
R1932 VTAIL.n232 VTAIL.n195 0.155672
R1933 VTAIL.n232 VTAIL.n231 0.155672
R1934 VTAIL.n231 VTAIL.n199 0.155672
R1935 VTAIL.n224 VTAIL.n199 0.155672
R1936 VTAIL.n224 VTAIL.n223 0.155672
R1937 VTAIL.n223 VTAIL.n203 0.155672
R1938 VTAIL.n216 VTAIL.n203 0.155672
R1939 VTAIL.n216 VTAIL.n215 0.155672
R1940 VTAIL.n215 VTAIL.n207 0.155672
R1941 VTAIL.n175 VTAIL.n93 0.155672
R1942 VTAIL.n168 VTAIL.n93 0.155672
R1943 VTAIL.n168 VTAIL.n167 0.155672
R1944 VTAIL.n167 VTAIL.n97 0.155672
R1945 VTAIL.n160 VTAIL.n97 0.155672
R1946 VTAIL.n160 VTAIL.n159 0.155672
R1947 VTAIL.n159 VTAIL.n103 0.155672
R1948 VTAIL.n152 VTAIL.n103 0.155672
R1949 VTAIL.n152 VTAIL.n151 0.155672
R1950 VTAIL.n151 VTAIL.n107 0.155672
R1951 VTAIL.n144 VTAIL.n107 0.155672
R1952 VTAIL.n144 VTAIL.n143 0.155672
R1953 VTAIL.n143 VTAIL.n111 0.155672
R1954 VTAIL.n136 VTAIL.n111 0.155672
R1955 VTAIL.n136 VTAIL.n135 0.155672
R1956 VTAIL.n135 VTAIL.n115 0.155672
R1957 VTAIL.n128 VTAIL.n115 0.155672
R1958 VTAIL.n128 VTAIL.n127 0.155672
R1959 VTAIL.n127 VTAIL.n119 0.155672
R1960 VDD1.n80 VDD1.n0 289.615
R1961 VDD1.n165 VDD1.n85 289.615
R1962 VDD1.n81 VDD1.n80 185
R1963 VDD1.n79 VDD1.n78 185
R1964 VDD1.n4 VDD1.n3 185
R1965 VDD1.n8 VDD1.n6 185
R1966 VDD1.n73 VDD1.n72 185
R1967 VDD1.n71 VDD1.n70 185
R1968 VDD1.n10 VDD1.n9 185
R1969 VDD1.n65 VDD1.n64 185
R1970 VDD1.n63 VDD1.n62 185
R1971 VDD1.n14 VDD1.n13 185
R1972 VDD1.n57 VDD1.n56 185
R1973 VDD1.n55 VDD1.n54 185
R1974 VDD1.n18 VDD1.n17 185
R1975 VDD1.n49 VDD1.n48 185
R1976 VDD1.n47 VDD1.n46 185
R1977 VDD1.n22 VDD1.n21 185
R1978 VDD1.n41 VDD1.n40 185
R1979 VDD1.n39 VDD1.n38 185
R1980 VDD1.n26 VDD1.n25 185
R1981 VDD1.n33 VDD1.n32 185
R1982 VDD1.n31 VDD1.n30 185
R1983 VDD1.n114 VDD1.n113 185
R1984 VDD1.n116 VDD1.n115 185
R1985 VDD1.n109 VDD1.n108 185
R1986 VDD1.n122 VDD1.n121 185
R1987 VDD1.n124 VDD1.n123 185
R1988 VDD1.n105 VDD1.n104 185
R1989 VDD1.n130 VDD1.n129 185
R1990 VDD1.n132 VDD1.n131 185
R1991 VDD1.n101 VDD1.n100 185
R1992 VDD1.n138 VDD1.n137 185
R1993 VDD1.n140 VDD1.n139 185
R1994 VDD1.n97 VDD1.n96 185
R1995 VDD1.n146 VDD1.n145 185
R1996 VDD1.n148 VDD1.n147 185
R1997 VDD1.n93 VDD1.n92 185
R1998 VDD1.n155 VDD1.n154 185
R1999 VDD1.n156 VDD1.n91 185
R2000 VDD1.n158 VDD1.n157 185
R2001 VDD1.n89 VDD1.n88 185
R2002 VDD1.n164 VDD1.n163 185
R2003 VDD1.n166 VDD1.n165 185
R2004 VDD1.n29 VDD1.t1 147.659
R2005 VDD1.n112 VDD1.t4 147.659
R2006 VDD1.n80 VDD1.n79 104.615
R2007 VDD1.n79 VDD1.n3 104.615
R2008 VDD1.n8 VDD1.n3 104.615
R2009 VDD1.n72 VDD1.n8 104.615
R2010 VDD1.n72 VDD1.n71 104.615
R2011 VDD1.n71 VDD1.n9 104.615
R2012 VDD1.n64 VDD1.n9 104.615
R2013 VDD1.n64 VDD1.n63 104.615
R2014 VDD1.n63 VDD1.n13 104.615
R2015 VDD1.n56 VDD1.n13 104.615
R2016 VDD1.n56 VDD1.n55 104.615
R2017 VDD1.n55 VDD1.n17 104.615
R2018 VDD1.n48 VDD1.n17 104.615
R2019 VDD1.n48 VDD1.n47 104.615
R2020 VDD1.n47 VDD1.n21 104.615
R2021 VDD1.n40 VDD1.n21 104.615
R2022 VDD1.n40 VDD1.n39 104.615
R2023 VDD1.n39 VDD1.n25 104.615
R2024 VDD1.n32 VDD1.n25 104.615
R2025 VDD1.n32 VDD1.n31 104.615
R2026 VDD1.n115 VDD1.n114 104.615
R2027 VDD1.n115 VDD1.n108 104.615
R2028 VDD1.n122 VDD1.n108 104.615
R2029 VDD1.n123 VDD1.n122 104.615
R2030 VDD1.n123 VDD1.n104 104.615
R2031 VDD1.n130 VDD1.n104 104.615
R2032 VDD1.n131 VDD1.n130 104.615
R2033 VDD1.n131 VDD1.n100 104.615
R2034 VDD1.n138 VDD1.n100 104.615
R2035 VDD1.n139 VDD1.n138 104.615
R2036 VDD1.n139 VDD1.n96 104.615
R2037 VDD1.n146 VDD1.n96 104.615
R2038 VDD1.n147 VDD1.n146 104.615
R2039 VDD1.n147 VDD1.n92 104.615
R2040 VDD1.n155 VDD1.n92 104.615
R2041 VDD1.n156 VDD1.n155 104.615
R2042 VDD1.n157 VDD1.n156 104.615
R2043 VDD1.n157 VDD1.n88 104.615
R2044 VDD1.n164 VDD1.n88 104.615
R2045 VDD1.n165 VDD1.n164 104.615
R2046 VDD1.n171 VDD1.n170 64.194
R2047 VDD1.n173 VDD1.n172 63.9454
R2048 VDD1 VDD1.n84 52.937
R2049 VDD1.n171 VDD1.n169 52.8235
R2050 VDD1.n31 VDD1.t1 52.3082
R2051 VDD1.n114 VDD1.t4 52.3082
R2052 VDD1.n173 VDD1.n171 42.2358
R2053 VDD1.n30 VDD1.n29 15.6677
R2054 VDD1.n113 VDD1.n112 15.6677
R2055 VDD1.n6 VDD1.n4 13.1884
R2056 VDD1.n158 VDD1.n89 13.1884
R2057 VDD1.n78 VDD1.n77 12.8005
R2058 VDD1.n74 VDD1.n73 12.8005
R2059 VDD1.n33 VDD1.n28 12.8005
R2060 VDD1.n116 VDD1.n111 12.8005
R2061 VDD1.n159 VDD1.n91 12.8005
R2062 VDD1.n163 VDD1.n162 12.8005
R2063 VDD1.n81 VDD1.n2 12.0247
R2064 VDD1.n70 VDD1.n7 12.0247
R2065 VDD1.n34 VDD1.n26 12.0247
R2066 VDD1.n117 VDD1.n109 12.0247
R2067 VDD1.n154 VDD1.n153 12.0247
R2068 VDD1.n166 VDD1.n87 12.0247
R2069 VDD1.n82 VDD1.n0 11.249
R2070 VDD1.n69 VDD1.n10 11.249
R2071 VDD1.n38 VDD1.n37 11.249
R2072 VDD1.n121 VDD1.n120 11.249
R2073 VDD1.n152 VDD1.n93 11.249
R2074 VDD1.n167 VDD1.n85 11.249
R2075 VDD1.n66 VDD1.n65 10.4732
R2076 VDD1.n41 VDD1.n24 10.4732
R2077 VDD1.n124 VDD1.n107 10.4732
R2078 VDD1.n149 VDD1.n148 10.4732
R2079 VDD1.n62 VDD1.n12 9.69747
R2080 VDD1.n42 VDD1.n22 9.69747
R2081 VDD1.n125 VDD1.n105 9.69747
R2082 VDD1.n145 VDD1.n95 9.69747
R2083 VDD1.n84 VDD1.n83 9.45567
R2084 VDD1.n169 VDD1.n168 9.45567
R2085 VDD1.n16 VDD1.n15 9.3005
R2086 VDD1.n59 VDD1.n58 9.3005
R2087 VDD1.n61 VDD1.n60 9.3005
R2088 VDD1.n12 VDD1.n11 9.3005
R2089 VDD1.n67 VDD1.n66 9.3005
R2090 VDD1.n69 VDD1.n68 9.3005
R2091 VDD1.n7 VDD1.n5 9.3005
R2092 VDD1.n75 VDD1.n74 9.3005
R2093 VDD1.n83 VDD1.n82 9.3005
R2094 VDD1.n2 VDD1.n1 9.3005
R2095 VDD1.n77 VDD1.n76 9.3005
R2096 VDD1.n53 VDD1.n52 9.3005
R2097 VDD1.n51 VDD1.n50 9.3005
R2098 VDD1.n20 VDD1.n19 9.3005
R2099 VDD1.n45 VDD1.n44 9.3005
R2100 VDD1.n43 VDD1.n42 9.3005
R2101 VDD1.n24 VDD1.n23 9.3005
R2102 VDD1.n37 VDD1.n36 9.3005
R2103 VDD1.n35 VDD1.n34 9.3005
R2104 VDD1.n28 VDD1.n27 9.3005
R2105 VDD1.n168 VDD1.n167 9.3005
R2106 VDD1.n87 VDD1.n86 9.3005
R2107 VDD1.n162 VDD1.n161 9.3005
R2108 VDD1.n134 VDD1.n133 9.3005
R2109 VDD1.n103 VDD1.n102 9.3005
R2110 VDD1.n128 VDD1.n127 9.3005
R2111 VDD1.n126 VDD1.n125 9.3005
R2112 VDD1.n107 VDD1.n106 9.3005
R2113 VDD1.n120 VDD1.n119 9.3005
R2114 VDD1.n118 VDD1.n117 9.3005
R2115 VDD1.n111 VDD1.n110 9.3005
R2116 VDD1.n136 VDD1.n135 9.3005
R2117 VDD1.n99 VDD1.n98 9.3005
R2118 VDD1.n142 VDD1.n141 9.3005
R2119 VDD1.n144 VDD1.n143 9.3005
R2120 VDD1.n95 VDD1.n94 9.3005
R2121 VDD1.n150 VDD1.n149 9.3005
R2122 VDD1.n152 VDD1.n151 9.3005
R2123 VDD1.n153 VDD1.n90 9.3005
R2124 VDD1.n160 VDD1.n159 9.3005
R2125 VDD1.n61 VDD1.n14 8.92171
R2126 VDD1.n46 VDD1.n45 8.92171
R2127 VDD1.n129 VDD1.n128 8.92171
R2128 VDD1.n144 VDD1.n97 8.92171
R2129 VDD1.n58 VDD1.n57 8.14595
R2130 VDD1.n49 VDD1.n20 8.14595
R2131 VDD1.n132 VDD1.n103 8.14595
R2132 VDD1.n141 VDD1.n140 8.14595
R2133 VDD1.n54 VDD1.n16 7.3702
R2134 VDD1.n50 VDD1.n18 7.3702
R2135 VDD1.n133 VDD1.n101 7.3702
R2136 VDD1.n137 VDD1.n99 7.3702
R2137 VDD1.n54 VDD1.n53 6.59444
R2138 VDD1.n53 VDD1.n18 6.59444
R2139 VDD1.n136 VDD1.n101 6.59444
R2140 VDD1.n137 VDD1.n136 6.59444
R2141 VDD1.n57 VDD1.n16 5.81868
R2142 VDD1.n50 VDD1.n49 5.81868
R2143 VDD1.n133 VDD1.n132 5.81868
R2144 VDD1.n140 VDD1.n99 5.81868
R2145 VDD1.n58 VDD1.n14 5.04292
R2146 VDD1.n46 VDD1.n20 5.04292
R2147 VDD1.n129 VDD1.n103 5.04292
R2148 VDD1.n141 VDD1.n97 5.04292
R2149 VDD1.n29 VDD1.n27 4.38563
R2150 VDD1.n112 VDD1.n110 4.38563
R2151 VDD1.n62 VDD1.n61 4.26717
R2152 VDD1.n45 VDD1.n22 4.26717
R2153 VDD1.n128 VDD1.n105 4.26717
R2154 VDD1.n145 VDD1.n144 4.26717
R2155 VDD1.n65 VDD1.n12 3.49141
R2156 VDD1.n42 VDD1.n41 3.49141
R2157 VDD1.n125 VDD1.n124 3.49141
R2158 VDD1.n148 VDD1.n95 3.49141
R2159 VDD1.n84 VDD1.n0 2.71565
R2160 VDD1.n66 VDD1.n10 2.71565
R2161 VDD1.n38 VDD1.n24 2.71565
R2162 VDD1.n121 VDD1.n107 2.71565
R2163 VDD1.n149 VDD1.n93 2.71565
R2164 VDD1.n169 VDD1.n85 2.71565
R2165 VDD1.n82 VDD1.n81 1.93989
R2166 VDD1.n70 VDD1.n69 1.93989
R2167 VDD1.n37 VDD1.n26 1.93989
R2168 VDD1.n120 VDD1.n109 1.93989
R2169 VDD1.n154 VDD1.n152 1.93989
R2170 VDD1.n167 VDD1.n166 1.93989
R2171 VDD1.n172 VDD1.t2 1.27627
R2172 VDD1.n172 VDD1.t3 1.27627
R2173 VDD1.n170 VDD1.t0 1.27627
R2174 VDD1.n170 VDD1.t5 1.27627
R2175 VDD1.n78 VDD1.n2 1.16414
R2176 VDD1.n73 VDD1.n7 1.16414
R2177 VDD1.n34 VDD1.n33 1.16414
R2178 VDD1.n117 VDD1.n116 1.16414
R2179 VDD1.n153 VDD1.n91 1.16414
R2180 VDD1.n163 VDD1.n87 1.16414
R2181 VDD1.n77 VDD1.n4 0.388379
R2182 VDD1.n74 VDD1.n6 0.388379
R2183 VDD1.n30 VDD1.n28 0.388379
R2184 VDD1.n113 VDD1.n111 0.388379
R2185 VDD1.n159 VDD1.n158 0.388379
R2186 VDD1.n162 VDD1.n89 0.388379
R2187 VDD1 VDD1.n173 0.24619
R2188 VDD1.n83 VDD1.n1 0.155672
R2189 VDD1.n76 VDD1.n1 0.155672
R2190 VDD1.n76 VDD1.n75 0.155672
R2191 VDD1.n75 VDD1.n5 0.155672
R2192 VDD1.n68 VDD1.n5 0.155672
R2193 VDD1.n68 VDD1.n67 0.155672
R2194 VDD1.n67 VDD1.n11 0.155672
R2195 VDD1.n60 VDD1.n11 0.155672
R2196 VDD1.n60 VDD1.n59 0.155672
R2197 VDD1.n59 VDD1.n15 0.155672
R2198 VDD1.n52 VDD1.n15 0.155672
R2199 VDD1.n52 VDD1.n51 0.155672
R2200 VDD1.n51 VDD1.n19 0.155672
R2201 VDD1.n44 VDD1.n19 0.155672
R2202 VDD1.n44 VDD1.n43 0.155672
R2203 VDD1.n43 VDD1.n23 0.155672
R2204 VDD1.n36 VDD1.n23 0.155672
R2205 VDD1.n36 VDD1.n35 0.155672
R2206 VDD1.n35 VDD1.n27 0.155672
R2207 VDD1.n118 VDD1.n110 0.155672
R2208 VDD1.n119 VDD1.n118 0.155672
R2209 VDD1.n119 VDD1.n106 0.155672
R2210 VDD1.n126 VDD1.n106 0.155672
R2211 VDD1.n127 VDD1.n126 0.155672
R2212 VDD1.n127 VDD1.n102 0.155672
R2213 VDD1.n134 VDD1.n102 0.155672
R2214 VDD1.n135 VDD1.n134 0.155672
R2215 VDD1.n135 VDD1.n98 0.155672
R2216 VDD1.n142 VDD1.n98 0.155672
R2217 VDD1.n143 VDD1.n142 0.155672
R2218 VDD1.n143 VDD1.n94 0.155672
R2219 VDD1.n150 VDD1.n94 0.155672
R2220 VDD1.n151 VDD1.n150 0.155672
R2221 VDD1.n151 VDD1.n90 0.155672
R2222 VDD1.n160 VDD1.n90 0.155672
R2223 VDD1.n161 VDD1.n160 0.155672
R2224 VDD1.n161 VDD1.n86 0.155672
R2225 VDD1.n168 VDD1.n86 0.155672
R2226 VN.n1 VN.t1 405.647
R2227 VN.n7 VN.t4 405.647
R2228 VN.n4 VN.t0 382.7
R2229 VN.n10 VN.t2 382.7
R2230 VN.n2 VN.t5 346.327
R2231 VN.n8 VN.t3 346.327
R2232 VN.n9 VN.n6 161.3
R2233 VN.n3 VN.n0 161.3
R2234 VN.n11 VN.n10 80.6037
R2235 VN.n5 VN.n4 80.6037
R2236 VN.n4 VN.n3 50.1678
R2237 VN.n10 VN.n9 50.1678
R2238 VN VN.n11 45.8362
R2239 VN.n2 VN.n1 32.6313
R2240 VN.n8 VN.n7 32.6313
R2241 VN.n7 VN.n6 28.168
R2242 VN.n1 VN.n0 28.168
R2243 VN.n3 VN.n2 24.5923
R2244 VN.n9 VN.n8 24.5923
R2245 VN.n11 VN.n6 0.285035
R2246 VN.n5 VN.n0 0.285035
R2247 VN VN.n5 0.146778
R2248 VDD2.n167 VDD2.n87 289.615
R2249 VDD2.n80 VDD2.n0 289.615
R2250 VDD2.n168 VDD2.n167 185
R2251 VDD2.n166 VDD2.n165 185
R2252 VDD2.n91 VDD2.n90 185
R2253 VDD2.n95 VDD2.n93 185
R2254 VDD2.n160 VDD2.n159 185
R2255 VDD2.n158 VDD2.n157 185
R2256 VDD2.n97 VDD2.n96 185
R2257 VDD2.n152 VDD2.n151 185
R2258 VDD2.n150 VDD2.n149 185
R2259 VDD2.n101 VDD2.n100 185
R2260 VDD2.n144 VDD2.n143 185
R2261 VDD2.n142 VDD2.n141 185
R2262 VDD2.n105 VDD2.n104 185
R2263 VDD2.n136 VDD2.n135 185
R2264 VDD2.n134 VDD2.n133 185
R2265 VDD2.n109 VDD2.n108 185
R2266 VDD2.n128 VDD2.n127 185
R2267 VDD2.n126 VDD2.n125 185
R2268 VDD2.n113 VDD2.n112 185
R2269 VDD2.n120 VDD2.n119 185
R2270 VDD2.n118 VDD2.n117 185
R2271 VDD2.n29 VDD2.n28 185
R2272 VDD2.n31 VDD2.n30 185
R2273 VDD2.n24 VDD2.n23 185
R2274 VDD2.n37 VDD2.n36 185
R2275 VDD2.n39 VDD2.n38 185
R2276 VDD2.n20 VDD2.n19 185
R2277 VDD2.n45 VDD2.n44 185
R2278 VDD2.n47 VDD2.n46 185
R2279 VDD2.n16 VDD2.n15 185
R2280 VDD2.n53 VDD2.n52 185
R2281 VDD2.n55 VDD2.n54 185
R2282 VDD2.n12 VDD2.n11 185
R2283 VDD2.n61 VDD2.n60 185
R2284 VDD2.n63 VDD2.n62 185
R2285 VDD2.n8 VDD2.n7 185
R2286 VDD2.n70 VDD2.n69 185
R2287 VDD2.n71 VDD2.n6 185
R2288 VDD2.n73 VDD2.n72 185
R2289 VDD2.n4 VDD2.n3 185
R2290 VDD2.n79 VDD2.n78 185
R2291 VDD2.n81 VDD2.n80 185
R2292 VDD2.n116 VDD2.t3 147.659
R2293 VDD2.n27 VDD2.t4 147.659
R2294 VDD2.n167 VDD2.n166 104.615
R2295 VDD2.n166 VDD2.n90 104.615
R2296 VDD2.n95 VDD2.n90 104.615
R2297 VDD2.n159 VDD2.n95 104.615
R2298 VDD2.n159 VDD2.n158 104.615
R2299 VDD2.n158 VDD2.n96 104.615
R2300 VDD2.n151 VDD2.n96 104.615
R2301 VDD2.n151 VDD2.n150 104.615
R2302 VDD2.n150 VDD2.n100 104.615
R2303 VDD2.n143 VDD2.n100 104.615
R2304 VDD2.n143 VDD2.n142 104.615
R2305 VDD2.n142 VDD2.n104 104.615
R2306 VDD2.n135 VDD2.n104 104.615
R2307 VDD2.n135 VDD2.n134 104.615
R2308 VDD2.n134 VDD2.n108 104.615
R2309 VDD2.n127 VDD2.n108 104.615
R2310 VDD2.n127 VDD2.n126 104.615
R2311 VDD2.n126 VDD2.n112 104.615
R2312 VDD2.n119 VDD2.n112 104.615
R2313 VDD2.n119 VDD2.n118 104.615
R2314 VDD2.n30 VDD2.n29 104.615
R2315 VDD2.n30 VDD2.n23 104.615
R2316 VDD2.n37 VDD2.n23 104.615
R2317 VDD2.n38 VDD2.n37 104.615
R2318 VDD2.n38 VDD2.n19 104.615
R2319 VDD2.n45 VDD2.n19 104.615
R2320 VDD2.n46 VDD2.n45 104.615
R2321 VDD2.n46 VDD2.n15 104.615
R2322 VDD2.n53 VDD2.n15 104.615
R2323 VDD2.n54 VDD2.n53 104.615
R2324 VDD2.n54 VDD2.n11 104.615
R2325 VDD2.n61 VDD2.n11 104.615
R2326 VDD2.n62 VDD2.n61 104.615
R2327 VDD2.n62 VDD2.n7 104.615
R2328 VDD2.n70 VDD2.n7 104.615
R2329 VDD2.n71 VDD2.n70 104.615
R2330 VDD2.n72 VDD2.n71 104.615
R2331 VDD2.n72 VDD2.n3 104.615
R2332 VDD2.n79 VDD2.n3 104.615
R2333 VDD2.n80 VDD2.n79 104.615
R2334 VDD2.n86 VDD2.n85 64.194
R2335 VDD2 VDD2.n173 64.1911
R2336 VDD2.n86 VDD2.n84 52.8235
R2337 VDD2.n118 VDD2.t3 52.3082
R2338 VDD2.n29 VDD2.t4 52.3082
R2339 VDD2.n172 VDD2.n171 51.9672
R2340 VDD2.n172 VDD2.n86 41.045
R2341 VDD2.n117 VDD2.n116 15.6677
R2342 VDD2.n28 VDD2.n27 15.6677
R2343 VDD2.n93 VDD2.n91 13.1884
R2344 VDD2.n73 VDD2.n4 13.1884
R2345 VDD2.n165 VDD2.n164 12.8005
R2346 VDD2.n161 VDD2.n160 12.8005
R2347 VDD2.n120 VDD2.n115 12.8005
R2348 VDD2.n31 VDD2.n26 12.8005
R2349 VDD2.n74 VDD2.n6 12.8005
R2350 VDD2.n78 VDD2.n77 12.8005
R2351 VDD2.n168 VDD2.n89 12.0247
R2352 VDD2.n157 VDD2.n94 12.0247
R2353 VDD2.n121 VDD2.n113 12.0247
R2354 VDD2.n32 VDD2.n24 12.0247
R2355 VDD2.n69 VDD2.n68 12.0247
R2356 VDD2.n81 VDD2.n2 12.0247
R2357 VDD2.n169 VDD2.n87 11.249
R2358 VDD2.n156 VDD2.n97 11.249
R2359 VDD2.n125 VDD2.n124 11.249
R2360 VDD2.n36 VDD2.n35 11.249
R2361 VDD2.n67 VDD2.n8 11.249
R2362 VDD2.n82 VDD2.n0 11.249
R2363 VDD2.n153 VDD2.n152 10.4732
R2364 VDD2.n128 VDD2.n111 10.4732
R2365 VDD2.n39 VDD2.n22 10.4732
R2366 VDD2.n64 VDD2.n63 10.4732
R2367 VDD2.n149 VDD2.n99 9.69747
R2368 VDD2.n129 VDD2.n109 9.69747
R2369 VDD2.n40 VDD2.n20 9.69747
R2370 VDD2.n60 VDD2.n10 9.69747
R2371 VDD2.n171 VDD2.n170 9.45567
R2372 VDD2.n84 VDD2.n83 9.45567
R2373 VDD2.n103 VDD2.n102 9.3005
R2374 VDD2.n146 VDD2.n145 9.3005
R2375 VDD2.n148 VDD2.n147 9.3005
R2376 VDD2.n99 VDD2.n98 9.3005
R2377 VDD2.n154 VDD2.n153 9.3005
R2378 VDD2.n156 VDD2.n155 9.3005
R2379 VDD2.n94 VDD2.n92 9.3005
R2380 VDD2.n162 VDD2.n161 9.3005
R2381 VDD2.n170 VDD2.n169 9.3005
R2382 VDD2.n89 VDD2.n88 9.3005
R2383 VDD2.n164 VDD2.n163 9.3005
R2384 VDD2.n140 VDD2.n139 9.3005
R2385 VDD2.n138 VDD2.n137 9.3005
R2386 VDD2.n107 VDD2.n106 9.3005
R2387 VDD2.n132 VDD2.n131 9.3005
R2388 VDD2.n130 VDD2.n129 9.3005
R2389 VDD2.n111 VDD2.n110 9.3005
R2390 VDD2.n124 VDD2.n123 9.3005
R2391 VDD2.n122 VDD2.n121 9.3005
R2392 VDD2.n115 VDD2.n114 9.3005
R2393 VDD2.n83 VDD2.n82 9.3005
R2394 VDD2.n2 VDD2.n1 9.3005
R2395 VDD2.n77 VDD2.n76 9.3005
R2396 VDD2.n49 VDD2.n48 9.3005
R2397 VDD2.n18 VDD2.n17 9.3005
R2398 VDD2.n43 VDD2.n42 9.3005
R2399 VDD2.n41 VDD2.n40 9.3005
R2400 VDD2.n22 VDD2.n21 9.3005
R2401 VDD2.n35 VDD2.n34 9.3005
R2402 VDD2.n33 VDD2.n32 9.3005
R2403 VDD2.n26 VDD2.n25 9.3005
R2404 VDD2.n51 VDD2.n50 9.3005
R2405 VDD2.n14 VDD2.n13 9.3005
R2406 VDD2.n57 VDD2.n56 9.3005
R2407 VDD2.n59 VDD2.n58 9.3005
R2408 VDD2.n10 VDD2.n9 9.3005
R2409 VDD2.n65 VDD2.n64 9.3005
R2410 VDD2.n67 VDD2.n66 9.3005
R2411 VDD2.n68 VDD2.n5 9.3005
R2412 VDD2.n75 VDD2.n74 9.3005
R2413 VDD2.n148 VDD2.n101 8.92171
R2414 VDD2.n133 VDD2.n132 8.92171
R2415 VDD2.n44 VDD2.n43 8.92171
R2416 VDD2.n59 VDD2.n12 8.92171
R2417 VDD2.n145 VDD2.n144 8.14595
R2418 VDD2.n136 VDD2.n107 8.14595
R2419 VDD2.n47 VDD2.n18 8.14595
R2420 VDD2.n56 VDD2.n55 8.14595
R2421 VDD2.n141 VDD2.n103 7.3702
R2422 VDD2.n137 VDD2.n105 7.3702
R2423 VDD2.n48 VDD2.n16 7.3702
R2424 VDD2.n52 VDD2.n14 7.3702
R2425 VDD2.n141 VDD2.n140 6.59444
R2426 VDD2.n140 VDD2.n105 6.59444
R2427 VDD2.n51 VDD2.n16 6.59444
R2428 VDD2.n52 VDD2.n51 6.59444
R2429 VDD2.n144 VDD2.n103 5.81868
R2430 VDD2.n137 VDD2.n136 5.81868
R2431 VDD2.n48 VDD2.n47 5.81868
R2432 VDD2.n55 VDD2.n14 5.81868
R2433 VDD2.n145 VDD2.n101 5.04292
R2434 VDD2.n133 VDD2.n107 5.04292
R2435 VDD2.n44 VDD2.n18 5.04292
R2436 VDD2.n56 VDD2.n12 5.04292
R2437 VDD2.n116 VDD2.n114 4.38563
R2438 VDD2.n27 VDD2.n25 4.38563
R2439 VDD2.n149 VDD2.n148 4.26717
R2440 VDD2.n132 VDD2.n109 4.26717
R2441 VDD2.n43 VDD2.n20 4.26717
R2442 VDD2.n60 VDD2.n59 4.26717
R2443 VDD2.n152 VDD2.n99 3.49141
R2444 VDD2.n129 VDD2.n128 3.49141
R2445 VDD2.n40 VDD2.n39 3.49141
R2446 VDD2.n63 VDD2.n10 3.49141
R2447 VDD2.n171 VDD2.n87 2.71565
R2448 VDD2.n153 VDD2.n97 2.71565
R2449 VDD2.n125 VDD2.n111 2.71565
R2450 VDD2.n36 VDD2.n22 2.71565
R2451 VDD2.n64 VDD2.n8 2.71565
R2452 VDD2.n84 VDD2.n0 2.71565
R2453 VDD2.n169 VDD2.n168 1.93989
R2454 VDD2.n157 VDD2.n156 1.93989
R2455 VDD2.n124 VDD2.n113 1.93989
R2456 VDD2.n35 VDD2.n24 1.93989
R2457 VDD2.n69 VDD2.n67 1.93989
R2458 VDD2.n82 VDD2.n81 1.93989
R2459 VDD2.n173 VDD2.t2 1.27627
R2460 VDD2.n173 VDD2.t1 1.27627
R2461 VDD2.n85 VDD2.t0 1.27627
R2462 VDD2.n85 VDD2.t5 1.27627
R2463 VDD2.n165 VDD2.n89 1.16414
R2464 VDD2.n160 VDD2.n94 1.16414
R2465 VDD2.n121 VDD2.n120 1.16414
R2466 VDD2.n32 VDD2.n31 1.16414
R2467 VDD2.n68 VDD2.n6 1.16414
R2468 VDD2.n78 VDD2.n2 1.16414
R2469 VDD2 VDD2.n172 0.970328
R2470 VDD2.n164 VDD2.n91 0.388379
R2471 VDD2.n161 VDD2.n93 0.388379
R2472 VDD2.n117 VDD2.n115 0.388379
R2473 VDD2.n28 VDD2.n26 0.388379
R2474 VDD2.n74 VDD2.n73 0.388379
R2475 VDD2.n77 VDD2.n4 0.388379
R2476 VDD2.n170 VDD2.n88 0.155672
R2477 VDD2.n163 VDD2.n88 0.155672
R2478 VDD2.n163 VDD2.n162 0.155672
R2479 VDD2.n162 VDD2.n92 0.155672
R2480 VDD2.n155 VDD2.n92 0.155672
R2481 VDD2.n155 VDD2.n154 0.155672
R2482 VDD2.n154 VDD2.n98 0.155672
R2483 VDD2.n147 VDD2.n98 0.155672
R2484 VDD2.n147 VDD2.n146 0.155672
R2485 VDD2.n146 VDD2.n102 0.155672
R2486 VDD2.n139 VDD2.n102 0.155672
R2487 VDD2.n139 VDD2.n138 0.155672
R2488 VDD2.n138 VDD2.n106 0.155672
R2489 VDD2.n131 VDD2.n106 0.155672
R2490 VDD2.n131 VDD2.n130 0.155672
R2491 VDD2.n130 VDD2.n110 0.155672
R2492 VDD2.n123 VDD2.n110 0.155672
R2493 VDD2.n123 VDD2.n122 0.155672
R2494 VDD2.n122 VDD2.n114 0.155672
R2495 VDD2.n33 VDD2.n25 0.155672
R2496 VDD2.n34 VDD2.n33 0.155672
R2497 VDD2.n34 VDD2.n21 0.155672
R2498 VDD2.n41 VDD2.n21 0.155672
R2499 VDD2.n42 VDD2.n41 0.155672
R2500 VDD2.n42 VDD2.n17 0.155672
R2501 VDD2.n49 VDD2.n17 0.155672
R2502 VDD2.n50 VDD2.n49 0.155672
R2503 VDD2.n50 VDD2.n13 0.155672
R2504 VDD2.n57 VDD2.n13 0.155672
R2505 VDD2.n58 VDD2.n57 0.155672
R2506 VDD2.n58 VDD2.n9 0.155672
R2507 VDD2.n65 VDD2.n9 0.155672
R2508 VDD2.n66 VDD2.n65 0.155672
R2509 VDD2.n66 VDD2.n5 0.155672
R2510 VDD2.n75 VDD2.n5 0.155672
R2511 VDD2.n76 VDD2.n75 0.155672
R2512 VDD2.n76 VDD2.n1 0.155672
R2513 VDD2.n83 VDD2.n1 0.155672
C0 VTAIL VP 6.352951f
C1 VTAIL VDD1 10.5036f
C2 VTAIL VN 6.33833f
C3 VTAIL VDD2 10.539901f
C4 VDD1 VP 6.85931f
C5 VP VN 6.09786f
C6 VDD1 VN 0.149055f
C7 VDD2 VP 0.330547f
C8 VDD1 VDD2 0.85125f
C9 VDD2 VN 6.68292f
C10 VDD2 B 5.414504f
C11 VDD1 B 5.466732f
C12 VTAIL B 8.047722f
C13 VN B 9.07068f
C14 VP B 7.162646f
C15 VDD2.n0 B 0.031115f
C16 VDD2.n1 B 0.022137f
C17 VDD2.n2 B 0.011895f
C18 VDD2.n3 B 0.028117f
C19 VDD2.n4 B 0.012245f
C20 VDD2.n5 B 0.022137f
C21 VDD2.n6 B 0.012595f
C22 VDD2.n7 B 0.028117f
C23 VDD2.n8 B 0.012595f
C24 VDD2.n9 B 0.022137f
C25 VDD2.n10 B 0.011895f
C26 VDD2.n11 B 0.028117f
C27 VDD2.n12 B 0.012595f
C28 VDD2.n13 B 0.022137f
C29 VDD2.n14 B 0.011895f
C30 VDD2.n15 B 0.028117f
C31 VDD2.n16 B 0.012595f
C32 VDD2.n17 B 0.022137f
C33 VDD2.n18 B 0.011895f
C34 VDD2.n19 B 0.028117f
C35 VDD2.n20 B 0.012595f
C36 VDD2.n21 B 0.022137f
C37 VDD2.n22 B 0.011895f
C38 VDD2.n23 B 0.028117f
C39 VDD2.n24 B 0.012595f
C40 VDD2.n25 B 1.49302f
C41 VDD2.n26 B 0.011895f
C42 VDD2.t4 B 0.0464f
C43 VDD2.n27 B 0.147268f
C44 VDD2.n28 B 0.016609f
C45 VDD2.n29 B 0.021087f
C46 VDD2.n30 B 0.028117f
C47 VDD2.n31 B 0.012595f
C48 VDD2.n32 B 0.011895f
C49 VDD2.n33 B 0.022137f
C50 VDD2.n34 B 0.022137f
C51 VDD2.n35 B 0.011895f
C52 VDD2.n36 B 0.012595f
C53 VDD2.n37 B 0.028117f
C54 VDD2.n38 B 0.028117f
C55 VDD2.n39 B 0.012595f
C56 VDD2.n40 B 0.011895f
C57 VDD2.n41 B 0.022137f
C58 VDD2.n42 B 0.022137f
C59 VDD2.n43 B 0.011895f
C60 VDD2.n44 B 0.012595f
C61 VDD2.n45 B 0.028117f
C62 VDD2.n46 B 0.028117f
C63 VDD2.n47 B 0.012595f
C64 VDD2.n48 B 0.011895f
C65 VDD2.n49 B 0.022137f
C66 VDD2.n50 B 0.022137f
C67 VDD2.n51 B 0.011895f
C68 VDD2.n52 B 0.012595f
C69 VDD2.n53 B 0.028117f
C70 VDD2.n54 B 0.028117f
C71 VDD2.n55 B 0.012595f
C72 VDD2.n56 B 0.011895f
C73 VDD2.n57 B 0.022137f
C74 VDD2.n58 B 0.022137f
C75 VDD2.n59 B 0.011895f
C76 VDD2.n60 B 0.012595f
C77 VDD2.n61 B 0.028117f
C78 VDD2.n62 B 0.028117f
C79 VDD2.n63 B 0.012595f
C80 VDD2.n64 B 0.011895f
C81 VDD2.n65 B 0.022137f
C82 VDD2.n66 B 0.022137f
C83 VDD2.n67 B 0.011895f
C84 VDD2.n68 B 0.011895f
C85 VDD2.n69 B 0.012595f
C86 VDD2.n70 B 0.028117f
C87 VDD2.n71 B 0.028117f
C88 VDD2.n72 B 0.028117f
C89 VDD2.n73 B 0.012245f
C90 VDD2.n74 B 0.011895f
C91 VDD2.n75 B 0.022137f
C92 VDD2.n76 B 0.022137f
C93 VDD2.n77 B 0.011895f
C94 VDD2.n78 B 0.012595f
C95 VDD2.n79 B 0.028117f
C96 VDD2.n80 B 0.060867f
C97 VDD2.n81 B 0.012595f
C98 VDD2.n82 B 0.011895f
C99 VDD2.n83 B 0.056007f
C100 VDD2.n84 B 0.051187f
C101 VDD2.t0 B 0.271496f
C102 VDD2.t5 B 0.271496f
C103 VDD2.n85 B 2.46196f
C104 VDD2.n86 B 1.97852f
C105 VDD2.n87 B 0.031115f
C106 VDD2.n88 B 0.022137f
C107 VDD2.n89 B 0.011895f
C108 VDD2.n90 B 0.028117f
C109 VDD2.n91 B 0.012245f
C110 VDD2.n92 B 0.022137f
C111 VDD2.n93 B 0.012245f
C112 VDD2.n94 B 0.011895f
C113 VDD2.n95 B 0.028117f
C114 VDD2.n96 B 0.028117f
C115 VDD2.n97 B 0.012595f
C116 VDD2.n98 B 0.022137f
C117 VDD2.n99 B 0.011895f
C118 VDD2.n100 B 0.028117f
C119 VDD2.n101 B 0.012595f
C120 VDD2.n102 B 0.022137f
C121 VDD2.n103 B 0.011895f
C122 VDD2.n104 B 0.028117f
C123 VDD2.n105 B 0.012595f
C124 VDD2.n106 B 0.022137f
C125 VDD2.n107 B 0.011895f
C126 VDD2.n108 B 0.028117f
C127 VDD2.n109 B 0.012595f
C128 VDD2.n110 B 0.022137f
C129 VDD2.n111 B 0.011895f
C130 VDD2.n112 B 0.028117f
C131 VDD2.n113 B 0.012595f
C132 VDD2.n114 B 1.49302f
C133 VDD2.n115 B 0.011895f
C134 VDD2.t3 B 0.0464f
C135 VDD2.n116 B 0.147268f
C136 VDD2.n117 B 0.016609f
C137 VDD2.n118 B 0.021087f
C138 VDD2.n119 B 0.028117f
C139 VDD2.n120 B 0.012595f
C140 VDD2.n121 B 0.011895f
C141 VDD2.n122 B 0.022137f
C142 VDD2.n123 B 0.022137f
C143 VDD2.n124 B 0.011895f
C144 VDD2.n125 B 0.012595f
C145 VDD2.n126 B 0.028117f
C146 VDD2.n127 B 0.028117f
C147 VDD2.n128 B 0.012595f
C148 VDD2.n129 B 0.011895f
C149 VDD2.n130 B 0.022137f
C150 VDD2.n131 B 0.022137f
C151 VDD2.n132 B 0.011895f
C152 VDD2.n133 B 0.012595f
C153 VDD2.n134 B 0.028117f
C154 VDD2.n135 B 0.028117f
C155 VDD2.n136 B 0.012595f
C156 VDD2.n137 B 0.011895f
C157 VDD2.n138 B 0.022137f
C158 VDD2.n139 B 0.022137f
C159 VDD2.n140 B 0.011895f
C160 VDD2.n141 B 0.012595f
C161 VDD2.n142 B 0.028117f
C162 VDD2.n143 B 0.028117f
C163 VDD2.n144 B 0.012595f
C164 VDD2.n145 B 0.011895f
C165 VDD2.n146 B 0.022137f
C166 VDD2.n147 B 0.022137f
C167 VDD2.n148 B 0.011895f
C168 VDD2.n149 B 0.012595f
C169 VDD2.n150 B 0.028117f
C170 VDD2.n151 B 0.028117f
C171 VDD2.n152 B 0.012595f
C172 VDD2.n153 B 0.011895f
C173 VDD2.n154 B 0.022137f
C174 VDD2.n155 B 0.022137f
C175 VDD2.n156 B 0.011895f
C176 VDD2.n157 B 0.012595f
C177 VDD2.n158 B 0.028117f
C178 VDD2.n159 B 0.028117f
C179 VDD2.n160 B 0.012595f
C180 VDD2.n161 B 0.011895f
C181 VDD2.n162 B 0.022137f
C182 VDD2.n163 B 0.022137f
C183 VDD2.n164 B 0.011895f
C184 VDD2.n165 B 0.012595f
C185 VDD2.n166 B 0.028117f
C186 VDD2.n167 B 0.060867f
C187 VDD2.n168 B 0.012595f
C188 VDD2.n169 B 0.011895f
C189 VDD2.n170 B 0.056007f
C190 VDD2.n171 B 0.049451f
C191 VDD2.n172 B 2.14508f
C192 VDD2.t2 B 0.271496f
C193 VDD2.t1 B 0.271496f
C194 VDD2.n173 B 2.46194f
C195 VN.n0 B 0.209788f
C196 VN.t5 B 1.74307f
C197 VN.t1 B 1.84507f
C198 VN.n1 B 0.676304f
C199 VN.n2 B 0.68976f
C200 VN.n3 B 0.048464f
C201 VN.t0 B 1.80543f
C202 VN.n4 B 0.691294f
C203 VN.n5 B 0.035515f
C204 VN.n6 B 0.209788f
C205 VN.t3 B 1.74307f
C206 VN.t4 B 1.84507f
C207 VN.n7 B 0.676304f
C208 VN.n8 B 0.68976f
C209 VN.n9 B 0.048464f
C210 VN.t2 B 1.80543f
C211 VN.n10 B 0.691294f
C212 VN.n11 B 1.82015f
C213 VDD1.n0 B 0.031328f
C214 VDD1.n1 B 0.022288f
C215 VDD1.n2 B 0.011977f
C216 VDD1.n3 B 0.028309f
C217 VDD1.n4 B 0.012329f
C218 VDD1.n5 B 0.022288f
C219 VDD1.n6 B 0.012329f
C220 VDD1.n7 B 0.011977f
C221 VDD1.n8 B 0.028309f
C222 VDD1.n9 B 0.028309f
C223 VDD1.n10 B 0.012681f
C224 VDD1.n11 B 0.022288f
C225 VDD1.n12 B 0.011977f
C226 VDD1.n13 B 0.028309f
C227 VDD1.n14 B 0.012681f
C228 VDD1.n15 B 0.022288f
C229 VDD1.n16 B 0.011977f
C230 VDD1.n17 B 0.028309f
C231 VDD1.n18 B 0.012681f
C232 VDD1.n19 B 0.022288f
C233 VDD1.n20 B 0.011977f
C234 VDD1.n21 B 0.028309f
C235 VDD1.n22 B 0.012681f
C236 VDD1.n23 B 0.022288f
C237 VDD1.n24 B 0.011977f
C238 VDD1.n25 B 0.028309f
C239 VDD1.n26 B 0.012681f
C240 VDD1.n27 B 1.50323f
C241 VDD1.n28 B 0.011977f
C242 VDD1.t1 B 0.046718f
C243 VDD1.n29 B 0.148276f
C244 VDD1.n30 B 0.016723f
C245 VDD1.n31 B 0.021232f
C246 VDD1.n32 B 0.028309f
C247 VDD1.n33 B 0.012681f
C248 VDD1.n34 B 0.011977f
C249 VDD1.n35 B 0.022288f
C250 VDD1.n36 B 0.022288f
C251 VDD1.n37 B 0.011977f
C252 VDD1.n38 B 0.012681f
C253 VDD1.n39 B 0.028309f
C254 VDD1.n40 B 0.028309f
C255 VDD1.n41 B 0.012681f
C256 VDD1.n42 B 0.011977f
C257 VDD1.n43 B 0.022288f
C258 VDD1.n44 B 0.022288f
C259 VDD1.n45 B 0.011977f
C260 VDD1.n46 B 0.012681f
C261 VDD1.n47 B 0.028309f
C262 VDD1.n48 B 0.028309f
C263 VDD1.n49 B 0.012681f
C264 VDD1.n50 B 0.011977f
C265 VDD1.n51 B 0.022288f
C266 VDD1.n52 B 0.022288f
C267 VDD1.n53 B 0.011977f
C268 VDD1.n54 B 0.012681f
C269 VDD1.n55 B 0.028309f
C270 VDD1.n56 B 0.028309f
C271 VDD1.n57 B 0.012681f
C272 VDD1.n58 B 0.011977f
C273 VDD1.n59 B 0.022288f
C274 VDD1.n60 B 0.022288f
C275 VDD1.n61 B 0.011977f
C276 VDD1.n62 B 0.012681f
C277 VDD1.n63 B 0.028309f
C278 VDD1.n64 B 0.028309f
C279 VDD1.n65 B 0.012681f
C280 VDD1.n66 B 0.011977f
C281 VDD1.n67 B 0.022288f
C282 VDD1.n68 B 0.022288f
C283 VDD1.n69 B 0.011977f
C284 VDD1.n70 B 0.012681f
C285 VDD1.n71 B 0.028309f
C286 VDD1.n72 B 0.028309f
C287 VDD1.n73 B 0.012681f
C288 VDD1.n74 B 0.011977f
C289 VDD1.n75 B 0.022288f
C290 VDD1.n76 B 0.022288f
C291 VDD1.n77 B 0.011977f
C292 VDD1.n78 B 0.012681f
C293 VDD1.n79 B 0.028309f
C294 VDD1.n80 B 0.061284f
C295 VDD1.n81 B 0.012681f
C296 VDD1.n82 B 0.011977f
C297 VDD1.n83 B 0.05639f
C298 VDD1.n84 B 0.051903f
C299 VDD1.n85 B 0.031328f
C300 VDD1.n86 B 0.022288f
C301 VDD1.n87 B 0.011977f
C302 VDD1.n88 B 0.028309f
C303 VDD1.n89 B 0.012329f
C304 VDD1.n90 B 0.022288f
C305 VDD1.n91 B 0.012681f
C306 VDD1.n92 B 0.028309f
C307 VDD1.n93 B 0.012681f
C308 VDD1.n94 B 0.022288f
C309 VDD1.n95 B 0.011977f
C310 VDD1.n96 B 0.028309f
C311 VDD1.n97 B 0.012681f
C312 VDD1.n98 B 0.022288f
C313 VDD1.n99 B 0.011977f
C314 VDD1.n100 B 0.028309f
C315 VDD1.n101 B 0.012681f
C316 VDD1.n102 B 0.022288f
C317 VDD1.n103 B 0.011977f
C318 VDD1.n104 B 0.028309f
C319 VDD1.n105 B 0.012681f
C320 VDD1.n106 B 0.022288f
C321 VDD1.n107 B 0.011977f
C322 VDD1.n108 B 0.028309f
C323 VDD1.n109 B 0.012681f
C324 VDD1.n110 B 1.50323f
C325 VDD1.n111 B 0.011977f
C326 VDD1.t4 B 0.046718f
C327 VDD1.n112 B 0.148276f
C328 VDD1.n113 B 0.016723f
C329 VDD1.n114 B 0.021232f
C330 VDD1.n115 B 0.028309f
C331 VDD1.n116 B 0.012681f
C332 VDD1.n117 B 0.011977f
C333 VDD1.n118 B 0.022288f
C334 VDD1.n119 B 0.022288f
C335 VDD1.n120 B 0.011977f
C336 VDD1.n121 B 0.012681f
C337 VDD1.n122 B 0.028309f
C338 VDD1.n123 B 0.028309f
C339 VDD1.n124 B 0.012681f
C340 VDD1.n125 B 0.011977f
C341 VDD1.n126 B 0.022288f
C342 VDD1.n127 B 0.022288f
C343 VDD1.n128 B 0.011977f
C344 VDD1.n129 B 0.012681f
C345 VDD1.n130 B 0.028309f
C346 VDD1.n131 B 0.028309f
C347 VDD1.n132 B 0.012681f
C348 VDD1.n133 B 0.011977f
C349 VDD1.n134 B 0.022288f
C350 VDD1.n135 B 0.022288f
C351 VDD1.n136 B 0.011977f
C352 VDD1.n137 B 0.012681f
C353 VDD1.n138 B 0.028309f
C354 VDD1.n139 B 0.028309f
C355 VDD1.n140 B 0.012681f
C356 VDD1.n141 B 0.011977f
C357 VDD1.n142 B 0.022288f
C358 VDD1.n143 B 0.022288f
C359 VDD1.n144 B 0.011977f
C360 VDD1.n145 B 0.012681f
C361 VDD1.n146 B 0.028309f
C362 VDD1.n147 B 0.028309f
C363 VDD1.n148 B 0.012681f
C364 VDD1.n149 B 0.011977f
C365 VDD1.n150 B 0.022288f
C366 VDD1.n151 B 0.022288f
C367 VDD1.n152 B 0.011977f
C368 VDD1.n153 B 0.011977f
C369 VDD1.n154 B 0.012681f
C370 VDD1.n155 B 0.028309f
C371 VDD1.n156 B 0.028309f
C372 VDD1.n157 B 0.028309f
C373 VDD1.n158 B 0.012329f
C374 VDD1.n159 B 0.011977f
C375 VDD1.n160 B 0.022288f
C376 VDD1.n161 B 0.022288f
C377 VDD1.n162 B 0.011977f
C378 VDD1.n163 B 0.012681f
C379 VDD1.n164 B 0.028309f
C380 VDD1.n165 B 0.061284f
C381 VDD1.n166 B 0.012681f
C382 VDD1.n167 B 0.011977f
C383 VDD1.n168 B 0.05639f
C384 VDD1.n169 B 0.051537f
C385 VDD1.t0 B 0.273353f
C386 VDD1.t5 B 0.273353f
C387 VDD1.n170 B 2.4788f
C388 VDD1.n171 B 2.07002f
C389 VDD1.t2 B 0.273353f
C390 VDD1.t3 B 0.273353f
C391 VDD1.n172 B 2.47765f
C392 VDD1.n173 B 2.34273f
C393 VTAIL.t10 B 0.281073f
C394 VTAIL.t2 B 0.281073f
C395 VTAIL.n0 B 2.48383f
C396 VTAIL.n1 B 0.324097f
C397 VTAIL.n2 B 0.032213f
C398 VTAIL.n3 B 0.022918f
C399 VTAIL.n4 B 0.012315f
C400 VTAIL.n5 B 0.029108f
C401 VTAIL.n6 B 0.012677f
C402 VTAIL.n7 B 0.022918f
C403 VTAIL.n8 B 0.01304f
C404 VTAIL.n9 B 0.029108f
C405 VTAIL.n10 B 0.01304f
C406 VTAIL.n11 B 0.022918f
C407 VTAIL.n12 B 0.012315f
C408 VTAIL.n13 B 0.029108f
C409 VTAIL.n14 B 0.01304f
C410 VTAIL.n15 B 0.022918f
C411 VTAIL.n16 B 0.012315f
C412 VTAIL.n17 B 0.029108f
C413 VTAIL.n18 B 0.01304f
C414 VTAIL.n19 B 0.022918f
C415 VTAIL.n20 B 0.012315f
C416 VTAIL.n21 B 0.029108f
C417 VTAIL.n22 B 0.01304f
C418 VTAIL.n23 B 0.022918f
C419 VTAIL.n24 B 0.012315f
C420 VTAIL.n25 B 0.029108f
C421 VTAIL.n26 B 0.01304f
C422 VTAIL.n27 B 1.54568f
C423 VTAIL.n28 B 0.012315f
C424 VTAIL.t3 B 0.048037f
C425 VTAIL.n29 B 0.152463f
C426 VTAIL.n30 B 0.017195f
C427 VTAIL.n31 B 0.021831f
C428 VTAIL.n32 B 0.029108f
C429 VTAIL.n33 B 0.01304f
C430 VTAIL.n34 B 0.012315f
C431 VTAIL.n35 B 0.022918f
C432 VTAIL.n36 B 0.022918f
C433 VTAIL.n37 B 0.012315f
C434 VTAIL.n38 B 0.01304f
C435 VTAIL.n39 B 0.029108f
C436 VTAIL.n40 B 0.029108f
C437 VTAIL.n41 B 0.01304f
C438 VTAIL.n42 B 0.012315f
C439 VTAIL.n43 B 0.022918f
C440 VTAIL.n44 B 0.022918f
C441 VTAIL.n45 B 0.012315f
C442 VTAIL.n46 B 0.01304f
C443 VTAIL.n47 B 0.029108f
C444 VTAIL.n48 B 0.029108f
C445 VTAIL.n49 B 0.01304f
C446 VTAIL.n50 B 0.012315f
C447 VTAIL.n51 B 0.022918f
C448 VTAIL.n52 B 0.022918f
C449 VTAIL.n53 B 0.012315f
C450 VTAIL.n54 B 0.01304f
C451 VTAIL.n55 B 0.029108f
C452 VTAIL.n56 B 0.029108f
C453 VTAIL.n57 B 0.01304f
C454 VTAIL.n58 B 0.012315f
C455 VTAIL.n59 B 0.022918f
C456 VTAIL.n60 B 0.022918f
C457 VTAIL.n61 B 0.012315f
C458 VTAIL.n62 B 0.01304f
C459 VTAIL.n63 B 0.029108f
C460 VTAIL.n64 B 0.029108f
C461 VTAIL.n65 B 0.01304f
C462 VTAIL.n66 B 0.012315f
C463 VTAIL.n67 B 0.022918f
C464 VTAIL.n68 B 0.022918f
C465 VTAIL.n69 B 0.012315f
C466 VTAIL.n70 B 0.012315f
C467 VTAIL.n71 B 0.01304f
C468 VTAIL.n72 B 0.029108f
C469 VTAIL.n73 B 0.029108f
C470 VTAIL.n74 B 0.029108f
C471 VTAIL.n75 B 0.012677f
C472 VTAIL.n76 B 0.012315f
C473 VTAIL.n77 B 0.022918f
C474 VTAIL.n78 B 0.022918f
C475 VTAIL.n79 B 0.012315f
C476 VTAIL.n80 B 0.01304f
C477 VTAIL.n81 B 0.029108f
C478 VTAIL.n82 B 0.063014f
C479 VTAIL.n83 B 0.01304f
C480 VTAIL.n84 B 0.012315f
C481 VTAIL.n85 B 0.057983f
C482 VTAIL.n86 B 0.035407f
C483 VTAIL.n87 B 0.191744f
C484 VTAIL.t7 B 0.281073f
C485 VTAIL.t6 B 0.281073f
C486 VTAIL.n88 B 2.48383f
C487 VTAIL.n89 B 1.78639f
C488 VTAIL.t9 B 0.281073f
C489 VTAIL.t11 B 0.281073f
C490 VTAIL.n90 B 2.48384f
C491 VTAIL.n91 B 1.78638f
C492 VTAIL.n92 B 0.032213f
C493 VTAIL.n93 B 0.022918f
C494 VTAIL.n94 B 0.012315f
C495 VTAIL.n95 B 0.029108f
C496 VTAIL.n96 B 0.012677f
C497 VTAIL.n97 B 0.022918f
C498 VTAIL.n98 B 0.012677f
C499 VTAIL.n99 B 0.012315f
C500 VTAIL.n100 B 0.029108f
C501 VTAIL.n101 B 0.029108f
C502 VTAIL.n102 B 0.01304f
C503 VTAIL.n103 B 0.022918f
C504 VTAIL.n104 B 0.012315f
C505 VTAIL.n105 B 0.029108f
C506 VTAIL.n106 B 0.01304f
C507 VTAIL.n107 B 0.022918f
C508 VTAIL.n108 B 0.012315f
C509 VTAIL.n109 B 0.029108f
C510 VTAIL.n110 B 0.01304f
C511 VTAIL.n111 B 0.022918f
C512 VTAIL.n112 B 0.012315f
C513 VTAIL.n113 B 0.029108f
C514 VTAIL.n114 B 0.01304f
C515 VTAIL.n115 B 0.022918f
C516 VTAIL.n116 B 0.012315f
C517 VTAIL.n117 B 0.029108f
C518 VTAIL.n118 B 0.01304f
C519 VTAIL.n119 B 1.54568f
C520 VTAIL.n120 B 0.012315f
C521 VTAIL.t1 B 0.048037f
C522 VTAIL.n121 B 0.152463f
C523 VTAIL.n122 B 0.017195f
C524 VTAIL.n123 B 0.021831f
C525 VTAIL.n124 B 0.029108f
C526 VTAIL.n125 B 0.01304f
C527 VTAIL.n126 B 0.012315f
C528 VTAIL.n127 B 0.022918f
C529 VTAIL.n128 B 0.022918f
C530 VTAIL.n129 B 0.012315f
C531 VTAIL.n130 B 0.01304f
C532 VTAIL.n131 B 0.029108f
C533 VTAIL.n132 B 0.029108f
C534 VTAIL.n133 B 0.01304f
C535 VTAIL.n134 B 0.012315f
C536 VTAIL.n135 B 0.022918f
C537 VTAIL.n136 B 0.022918f
C538 VTAIL.n137 B 0.012315f
C539 VTAIL.n138 B 0.01304f
C540 VTAIL.n139 B 0.029108f
C541 VTAIL.n140 B 0.029108f
C542 VTAIL.n141 B 0.01304f
C543 VTAIL.n142 B 0.012315f
C544 VTAIL.n143 B 0.022918f
C545 VTAIL.n144 B 0.022918f
C546 VTAIL.n145 B 0.012315f
C547 VTAIL.n146 B 0.01304f
C548 VTAIL.n147 B 0.029108f
C549 VTAIL.n148 B 0.029108f
C550 VTAIL.n149 B 0.01304f
C551 VTAIL.n150 B 0.012315f
C552 VTAIL.n151 B 0.022918f
C553 VTAIL.n152 B 0.022918f
C554 VTAIL.n153 B 0.012315f
C555 VTAIL.n154 B 0.01304f
C556 VTAIL.n155 B 0.029108f
C557 VTAIL.n156 B 0.029108f
C558 VTAIL.n157 B 0.01304f
C559 VTAIL.n158 B 0.012315f
C560 VTAIL.n159 B 0.022918f
C561 VTAIL.n160 B 0.022918f
C562 VTAIL.n161 B 0.012315f
C563 VTAIL.n162 B 0.01304f
C564 VTAIL.n163 B 0.029108f
C565 VTAIL.n164 B 0.029108f
C566 VTAIL.n165 B 0.01304f
C567 VTAIL.n166 B 0.012315f
C568 VTAIL.n167 B 0.022918f
C569 VTAIL.n168 B 0.022918f
C570 VTAIL.n169 B 0.012315f
C571 VTAIL.n170 B 0.01304f
C572 VTAIL.n171 B 0.029108f
C573 VTAIL.n172 B 0.063014f
C574 VTAIL.n173 B 0.01304f
C575 VTAIL.n174 B 0.012315f
C576 VTAIL.n175 B 0.057983f
C577 VTAIL.n176 B 0.035407f
C578 VTAIL.n177 B 0.191744f
C579 VTAIL.t8 B 0.281073f
C580 VTAIL.t4 B 0.281073f
C581 VTAIL.n178 B 2.48384f
C582 VTAIL.n179 B 0.38711f
C583 VTAIL.n180 B 0.032213f
C584 VTAIL.n181 B 0.022918f
C585 VTAIL.n182 B 0.012315f
C586 VTAIL.n183 B 0.029108f
C587 VTAIL.n184 B 0.012677f
C588 VTAIL.n185 B 0.022918f
C589 VTAIL.n186 B 0.012677f
C590 VTAIL.n187 B 0.012315f
C591 VTAIL.n188 B 0.029108f
C592 VTAIL.n189 B 0.029108f
C593 VTAIL.n190 B 0.01304f
C594 VTAIL.n191 B 0.022918f
C595 VTAIL.n192 B 0.012315f
C596 VTAIL.n193 B 0.029108f
C597 VTAIL.n194 B 0.01304f
C598 VTAIL.n195 B 0.022918f
C599 VTAIL.n196 B 0.012315f
C600 VTAIL.n197 B 0.029108f
C601 VTAIL.n198 B 0.01304f
C602 VTAIL.n199 B 0.022918f
C603 VTAIL.n200 B 0.012315f
C604 VTAIL.n201 B 0.029108f
C605 VTAIL.n202 B 0.01304f
C606 VTAIL.n203 B 0.022918f
C607 VTAIL.n204 B 0.012315f
C608 VTAIL.n205 B 0.029108f
C609 VTAIL.n206 B 0.01304f
C610 VTAIL.n207 B 1.54568f
C611 VTAIL.n208 B 0.012315f
C612 VTAIL.t5 B 0.048037f
C613 VTAIL.n209 B 0.152463f
C614 VTAIL.n210 B 0.017195f
C615 VTAIL.n211 B 0.021831f
C616 VTAIL.n212 B 0.029108f
C617 VTAIL.n213 B 0.01304f
C618 VTAIL.n214 B 0.012315f
C619 VTAIL.n215 B 0.022918f
C620 VTAIL.n216 B 0.022918f
C621 VTAIL.n217 B 0.012315f
C622 VTAIL.n218 B 0.01304f
C623 VTAIL.n219 B 0.029108f
C624 VTAIL.n220 B 0.029108f
C625 VTAIL.n221 B 0.01304f
C626 VTAIL.n222 B 0.012315f
C627 VTAIL.n223 B 0.022918f
C628 VTAIL.n224 B 0.022918f
C629 VTAIL.n225 B 0.012315f
C630 VTAIL.n226 B 0.01304f
C631 VTAIL.n227 B 0.029108f
C632 VTAIL.n228 B 0.029108f
C633 VTAIL.n229 B 0.01304f
C634 VTAIL.n230 B 0.012315f
C635 VTAIL.n231 B 0.022918f
C636 VTAIL.n232 B 0.022918f
C637 VTAIL.n233 B 0.012315f
C638 VTAIL.n234 B 0.01304f
C639 VTAIL.n235 B 0.029108f
C640 VTAIL.n236 B 0.029108f
C641 VTAIL.n237 B 0.01304f
C642 VTAIL.n238 B 0.012315f
C643 VTAIL.n239 B 0.022918f
C644 VTAIL.n240 B 0.022918f
C645 VTAIL.n241 B 0.012315f
C646 VTAIL.n242 B 0.01304f
C647 VTAIL.n243 B 0.029108f
C648 VTAIL.n244 B 0.029108f
C649 VTAIL.n245 B 0.01304f
C650 VTAIL.n246 B 0.012315f
C651 VTAIL.n247 B 0.022918f
C652 VTAIL.n248 B 0.022918f
C653 VTAIL.n249 B 0.012315f
C654 VTAIL.n250 B 0.01304f
C655 VTAIL.n251 B 0.029108f
C656 VTAIL.n252 B 0.029108f
C657 VTAIL.n253 B 0.01304f
C658 VTAIL.n254 B 0.012315f
C659 VTAIL.n255 B 0.022918f
C660 VTAIL.n256 B 0.022918f
C661 VTAIL.n257 B 0.012315f
C662 VTAIL.n258 B 0.01304f
C663 VTAIL.n259 B 0.029108f
C664 VTAIL.n260 B 0.063014f
C665 VTAIL.n261 B 0.01304f
C666 VTAIL.n262 B 0.012315f
C667 VTAIL.n263 B 0.057983f
C668 VTAIL.n264 B 0.035407f
C669 VTAIL.n265 B 1.50125f
C670 VTAIL.n266 B 0.032213f
C671 VTAIL.n267 B 0.022918f
C672 VTAIL.n268 B 0.012315f
C673 VTAIL.n269 B 0.029108f
C674 VTAIL.n270 B 0.012677f
C675 VTAIL.n271 B 0.022918f
C676 VTAIL.n272 B 0.01304f
C677 VTAIL.n273 B 0.029108f
C678 VTAIL.n274 B 0.01304f
C679 VTAIL.n275 B 0.022918f
C680 VTAIL.n276 B 0.012315f
C681 VTAIL.n277 B 0.029108f
C682 VTAIL.n278 B 0.01304f
C683 VTAIL.n279 B 0.022918f
C684 VTAIL.n280 B 0.012315f
C685 VTAIL.n281 B 0.029108f
C686 VTAIL.n282 B 0.01304f
C687 VTAIL.n283 B 0.022918f
C688 VTAIL.n284 B 0.012315f
C689 VTAIL.n285 B 0.029108f
C690 VTAIL.n286 B 0.01304f
C691 VTAIL.n287 B 0.022918f
C692 VTAIL.n288 B 0.012315f
C693 VTAIL.n289 B 0.029108f
C694 VTAIL.n290 B 0.01304f
C695 VTAIL.n291 B 1.54568f
C696 VTAIL.n292 B 0.012315f
C697 VTAIL.t0 B 0.048037f
C698 VTAIL.n293 B 0.152463f
C699 VTAIL.n294 B 0.017195f
C700 VTAIL.n295 B 0.021831f
C701 VTAIL.n296 B 0.029108f
C702 VTAIL.n297 B 0.01304f
C703 VTAIL.n298 B 0.012315f
C704 VTAIL.n299 B 0.022918f
C705 VTAIL.n300 B 0.022918f
C706 VTAIL.n301 B 0.012315f
C707 VTAIL.n302 B 0.01304f
C708 VTAIL.n303 B 0.029108f
C709 VTAIL.n304 B 0.029108f
C710 VTAIL.n305 B 0.01304f
C711 VTAIL.n306 B 0.012315f
C712 VTAIL.n307 B 0.022918f
C713 VTAIL.n308 B 0.022918f
C714 VTAIL.n309 B 0.012315f
C715 VTAIL.n310 B 0.01304f
C716 VTAIL.n311 B 0.029108f
C717 VTAIL.n312 B 0.029108f
C718 VTAIL.n313 B 0.01304f
C719 VTAIL.n314 B 0.012315f
C720 VTAIL.n315 B 0.022918f
C721 VTAIL.n316 B 0.022918f
C722 VTAIL.n317 B 0.012315f
C723 VTAIL.n318 B 0.01304f
C724 VTAIL.n319 B 0.029108f
C725 VTAIL.n320 B 0.029108f
C726 VTAIL.n321 B 0.01304f
C727 VTAIL.n322 B 0.012315f
C728 VTAIL.n323 B 0.022918f
C729 VTAIL.n324 B 0.022918f
C730 VTAIL.n325 B 0.012315f
C731 VTAIL.n326 B 0.01304f
C732 VTAIL.n327 B 0.029108f
C733 VTAIL.n328 B 0.029108f
C734 VTAIL.n329 B 0.01304f
C735 VTAIL.n330 B 0.012315f
C736 VTAIL.n331 B 0.022918f
C737 VTAIL.n332 B 0.022918f
C738 VTAIL.n333 B 0.012315f
C739 VTAIL.n334 B 0.012315f
C740 VTAIL.n335 B 0.01304f
C741 VTAIL.n336 B 0.029108f
C742 VTAIL.n337 B 0.029108f
C743 VTAIL.n338 B 0.029108f
C744 VTAIL.n339 B 0.012677f
C745 VTAIL.n340 B 0.012315f
C746 VTAIL.n341 B 0.022918f
C747 VTAIL.n342 B 0.022918f
C748 VTAIL.n343 B 0.012315f
C749 VTAIL.n344 B 0.01304f
C750 VTAIL.n345 B 0.029108f
C751 VTAIL.n346 B 0.063014f
C752 VTAIL.n347 B 0.01304f
C753 VTAIL.n348 B 0.012315f
C754 VTAIL.n349 B 0.057983f
C755 VTAIL.n350 B 0.035407f
C756 VTAIL.n351 B 1.47452f
C757 VP.n0 B 0.05154f
C758 VP.t5 B 1.7754f
C759 VP.n1 B 0.049363f
C760 VP.n2 B 0.21368f
C761 VP.t2 B 1.83892f
C762 VP.t3 B 1.7754f
C763 VP.t4 B 1.8793f
C764 VP.n3 B 0.688849f
C765 VP.n4 B 0.702555f
C766 VP.n5 B 0.049363f
C767 VP.n6 B 0.704117f
C768 VP.n7 B 1.83254f
C769 VP.t1 B 1.83892f
C770 VP.n8 B 0.704117f
C771 VP.n9 B 1.86311f
C772 VP.n10 B 0.05154f
C773 VP.n11 B 0.038625f
C774 VP.n12 B 0.676416f
C775 VP.n13 B 0.049363f
C776 VP.t0 B 1.83892f
C777 VP.n14 B 0.704117f
C778 VP.n15 B 0.036174f
.ends

