* NGSPICE file created from diff_pair_sample_0097.ext - technology: sky130A

.subckt diff_pair_sample_0097 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t4 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X1 VTAIL.t19 VP.t0 VDD1.t9 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X2 VDD1.t8 VP.t1 VTAIL.t1 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=2.04105 ps=12.7 w=12.37 l=2
X3 B.t11 B.t9 B.t10 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=0 ps=0 w=12.37 l=2
X4 VDD2.t2 VN.t1 VTAIL.t17 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=2.04105 ps=12.7 w=12.37 l=2
X5 VDD2.t8 VN.t2 VTAIL.t16 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=4.8243 ps=25.52 w=12.37 l=2
X6 VDD2.t5 VN.t3 VTAIL.t15 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X7 VTAIL.t14 VN.t4 VDD2.t6 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X8 B.t8 B.t6 B.t7 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=0 ps=0 w=12.37 l=2
X9 VTAIL.t8 VP.t2 VDD1.t7 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X10 VTAIL.t13 VN.t5 VDD2.t0 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X11 VDD1.t6 VP.t3 VTAIL.t2 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X12 VTAIL.t5 VP.t4 VDD1.t5 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X13 VTAIL.t3 VP.t5 VDD1.t4 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X14 VDD1.t3 VP.t6 VTAIL.t0 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=2.04105 ps=12.7 w=12.37 l=2
X15 VDD2.t1 VN.t6 VTAIL.t12 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X16 B.t5 B.t3 B.t4 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=0 ps=0 w=12.37 l=2
X17 VDD2.t9 VN.t7 VTAIL.t11 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=4.8243 ps=25.52 w=12.37 l=2
X18 VDD1.t2 VP.t7 VTAIL.t4 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=4.8243 ps=25.52 w=12.37 l=2
X19 VDD2.t3 VN.t8 VTAIL.t10 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=2.04105 ps=12.7 w=12.37 l=2
X20 VDD1.t1 VP.t8 VTAIL.t6 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X21 VDD1.t0 VP.t9 VTAIL.t7 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=4.8243 ps=25.52 w=12.37 l=2
X22 VTAIL.t9 VN.t9 VDD2.t7 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=2.04105 pd=12.7 as=2.04105 ps=12.7 w=12.37 l=2
X23 B.t2 B.t0 B.t1 w_n3766_n3442# sky130_fd_pr__pfet_01v8 ad=4.8243 pd=25.52 as=0 ps=0 w=12.37 l=2
R0 VN.n8 VN.t8 179.425
R1 VN.n42 VN.t2 179.425
R2 VN.n65 VN.n34 161.3
R3 VN.n64 VN.n63 161.3
R4 VN.n62 VN.n35 161.3
R5 VN.n61 VN.n60 161.3
R6 VN.n58 VN.n36 161.3
R7 VN.n57 VN.n56 161.3
R8 VN.n55 VN.n37 161.3
R9 VN.n54 VN.n53 161.3
R10 VN.n52 VN.n38 161.3
R11 VN.n50 VN.n49 161.3
R12 VN.n48 VN.n39 161.3
R13 VN.n47 VN.n46 161.3
R14 VN.n45 VN.n40 161.3
R15 VN.n44 VN.n43 161.3
R16 VN.n31 VN.n0 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n1 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n24 VN.n2 161.3
R21 VN.n23 VN.n22 161.3
R22 VN.n21 VN.n3 161.3
R23 VN.n20 VN.n19 161.3
R24 VN.n18 VN.n4 161.3
R25 VN.n16 VN.n15 161.3
R26 VN.n14 VN.n5 161.3
R27 VN.n13 VN.n12 161.3
R28 VN.n11 VN.n6 161.3
R29 VN.n10 VN.n9 161.3
R30 VN.n7 VN.t5 149.06
R31 VN.n17 VN.t6 149.06
R32 VN.n25 VN.t4 149.06
R33 VN.n32 VN.t7 149.06
R34 VN.n41 VN.t0 149.06
R35 VN.n51 VN.t3 149.06
R36 VN.n59 VN.t9 149.06
R37 VN.n66 VN.t1 149.06
R38 VN.n33 VN.n32 90.6935
R39 VN.n67 VN.n66 90.6935
R40 VN.n8 VN.n7 65.9005
R41 VN.n42 VN.n41 65.9005
R42 VN.n30 VN.n1 56.5193
R43 VN.n64 VN.n35 56.5193
R44 VN VN.n67 50.4413
R45 VN.n12 VN.n5 48.7492
R46 VN.n19 VN.n3 48.7492
R47 VN.n46 VN.n39 48.7492
R48 VN.n53 VN.n37 48.7492
R49 VN.n12 VN.n11 32.2376
R50 VN.n23 VN.n3 32.2376
R51 VN.n46 VN.n45 32.2376
R52 VN.n57 VN.n37 32.2376
R53 VN.n11 VN.n10 24.4675
R54 VN.n16 VN.n5 24.4675
R55 VN.n19 VN.n18 24.4675
R56 VN.n24 VN.n23 24.4675
R57 VN.n26 VN.n1 24.4675
R58 VN.n31 VN.n30 24.4675
R59 VN.n45 VN.n44 24.4675
R60 VN.n53 VN.n52 24.4675
R61 VN.n50 VN.n39 24.4675
R62 VN.n60 VN.n35 24.4675
R63 VN.n58 VN.n57 24.4675
R64 VN.n65 VN.n64 24.4675
R65 VN.n26 VN.n25 20.5528
R66 VN.n60 VN.n59 20.5528
R67 VN.n32 VN.n31 20.0634
R68 VN.n66 VN.n65 20.0634
R69 VN.n43 VN.n42 13.2957
R70 VN.n9 VN.n8 13.2957
R71 VN.n17 VN.n16 12.234
R72 VN.n18 VN.n17 12.234
R73 VN.n52 VN.n51 12.234
R74 VN.n51 VN.n50 12.234
R75 VN.n10 VN.n7 3.91522
R76 VN.n25 VN.n24 3.91522
R77 VN.n44 VN.n41 3.91522
R78 VN.n59 VN.n58 3.91522
R79 VN.n67 VN.n34 0.278367
R80 VN.n33 VN.n0 0.278367
R81 VN.n63 VN.n34 0.189894
R82 VN.n63 VN.n62 0.189894
R83 VN.n62 VN.n61 0.189894
R84 VN.n61 VN.n36 0.189894
R85 VN.n56 VN.n36 0.189894
R86 VN.n56 VN.n55 0.189894
R87 VN.n55 VN.n54 0.189894
R88 VN.n54 VN.n38 0.189894
R89 VN.n49 VN.n38 0.189894
R90 VN.n49 VN.n48 0.189894
R91 VN.n48 VN.n47 0.189894
R92 VN.n47 VN.n40 0.189894
R93 VN.n43 VN.n40 0.189894
R94 VN.n9 VN.n6 0.189894
R95 VN.n13 VN.n6 0.189894
R96 VN.n14 VN.n13 0.189894
R97 VN.n15 VN.n14 0.189894
R98 VN.n15 VN.n4 0.189894
R99 VN.n20 VN.n4 0.189894
R100 VN.n21 VN.n20 0.189894
R101 VN.n22 VN.n21 0.189894
R102 VN.n22 VN.n2 0.189894
R103 VN.n27 VN.n2 0.189894
R104 VN.n28 VN.n27 0.189894
R105 VN.n29 VN.n28 0.189894
R106 VN.n29 VN.n0 0.189894
R107 VN VN.n33 0.153454
R108 VDD2.n1 VDD2.t3 75.9146
R109 VDD2.n4 VDD2.t2 73.9061
R110 VDD2.n3 VDD2.n2 72.7293
R111 VDD2 VDD2.n7 72.7265
R112 VDD2.n6 VDD2.n5 71.2784
R113 VDD2.n1 VDD2.n0 71.2782
R114 VDD2.n4 VDD2.n3 43.92
R115 VDD2.n7 VDD2.t4 2.62823
R116 VDD2.n7 VDD2.t8 2.62823
R117 VDD2.n5 VDD2.t7 2.62823
R118 VDD2.n5 VDD2.t5 2.62823
R119 VDD2.n2 VDD2.t6 2.62823
R120 VDD2.n2 VDD2.t9 2.62823
R121 VDD2.n0 VDD2.t0 2.62823
R122 VDD2.n0 VDD2.t1 2.62823
R123 VDD2.n6 VDD2.n4 2.00912
R124 VDD2 VDD2.n6 0.560845
R125 VDD2.n3 VDD2.n1 0.447309
R126 VTAIL.n11 VTAIL.t16 57.2273
R127 VTAIL.n17 VTAIL.t11 57.2272
R128 VTAIL.n2 VTAIL.t7 57.2272
R129 VTAIL.n16 VTAIL.t4 57.2272
R130 VTAIL.n15 VTAIL.n14 54.5996
R131 VTAIL.n13 VTAIL.n12 54.5996
R132 VTAIL.n10 VTAIL.n9 54.5996
R133 VTAIL.n8 VTAIL.n7 54.5996
R134 VTAIL.n19 VTAIL.n18 54.5994
R135 VTAIL.n1 VTAIL.n0 54.5994
R136 VTAIL.n4 VTAIL.n3 54.5994
R137 VTAIL.n6 VTAIL.n5 54.5994
R138 VTAIL.n8 VTAIL.n6 27.0479
R139 VTAIL.n17 VTAIL.n16 25.0393
R140 VTAIL.n18 VTAIL.t12 2.62823
R141 VTAIL.n18 VTAIL.t14 2.62823
R142 VTAIL.n0 VTAIL.t10 2.62823
R143 VTAIL.n0 VTAIL.t13 2.62823
R144 VTAIL.n3 VTAIL.t2 2.62823
R145 VTAIL.n3 VTAIL.t3 2.62823
R146 VTAIL.n5 VTAIL.t0 2.62823
R147 VTAIL.n5 VTAIL.t19 2.62823
R148 VTAIL.n14 VTAIL.t6 2.62823
R149 VTAIL.n14 VTAIL.t8 2.62823
R150 VTAIL.n12 VTAIL.t1 2.62823
R151 VTAIL.n12 VTAIL.t5 2.62823
R152 VTAIL.n9 VTAIL.t15 2.62823
R153 VTAIL.n9 VTAIL.t18 2.62823
R154 VTAIL.n7 VTAIL.t17 2.62823
R155 VTAIL.n7 VTAIL.t9 2.62823
R156 VTAIL.n10 VTAIL.n8 2.00912
R157 VTAIL.n11 VTAIL.n10 2.00912
R158 VTAIL.n15 VTAIL.n13 2.00912
R159 VTAIL.n16 VTAIL.n15 2.00912
R160 VTAIL.n6 VTAIL.n4 2.00912
R161 VTAIL.n4 VTAIL.n2 2.00912
R162 VTAIL.n19 VTAIL.n17 2.00912
R163 VTAIL VTAIL.n1 1.56516
R164 VTAIL.n13 VTAIL.n11 1.47464
R165 VTAIL.n2 VTAIL.n1 1.47464
R166 VTAIL VTAIL.n19 0.444466
R167 VP.n18 VP.t1 179.425
R168 VP.n20 VP.n19 161.3
R169 VP.n21 VP.n16 161.3
R170 VP.n23 VP.n22 161.3
R171 VP.n24 VP.n15 161.3
R172 VP.n26 VP.n25 161.3
R173 VP.n28 VP.n14 161.3
R174 VP.n30 VP.n29 161.3
R175 VP.n31 VP.n13 161.3
R176 VP.n33 VP.n32 161.3
R177 VP.n34 VP.n12 161.3
R178 VP.n37 VP.n36 161.3
R179 VP.n38 VP.n11 161.3
R180 VP.n40 VP.n39 161.3
R181 VP.n41 VP.n10 161.3
R182 VP.n74 VP.n0 161.3
R183 VP.n73 VP.n72 161.3
R184 VP.n71 VP.n1 161.3
R185 VP.n70 VP.n69 161.3
R186 VP.n67 VP.n2 161.3
R187 VP.n66 VP.n65 161.3
R188 VP.n64 VP.n3 161.3
R189 VP.n63 VP.n62 161.3
R190 VP.n61 VP.n4 161.3
R191 VP.n59 VP.n58 161.3
R192 VP.n57 VP.n5 161.3
R193 VP.n56 VP.n55 161.3
R194 VP.n54 VP.n6 161.3
R195 VP.n53 VP.n52 161.3
R196 VP.n51 VP.n50 161.3
R197 VP.n49 VP.n8 161.3
R198 VP.n48 VP.n47 161.3
R199 VP.n46 VP.n9 161.3
R200 VP.n44 VP.t6 149.06
R201 VP.n7 VP.t0 149.06
R202 VP.n60 VP.t3 149.06
R203 VP.n68 VP.t5 149.06
R204 VP.n75 VP.t9 149.06
R205 VP.n42 VP.t7 149.06
R206 VP.n35 VP.t2 149.06
R207 VP.n27 VP.t8 149.06
R208 VP.n17 VP.t4 149.06
R209 VP.n45 VP.n44 90.6935
R210 VP.n76 VP.n75 90.6935
R211 VP.n43 VP.n42 90.6935
R212 VP.n18 VP.n17 65.9005
R213 VP.n49 VP.n48 56.5193
R214 VP.n73 VP.n1 56.5193
R215 VP.n40 VP.n11 56.5193
R216 VP.n45 VP.n43 50.1625
R217 VP.n55 VP.n5 48.7492
R218 VP.n62 VP.n3 48.7492
R219 VP.n29 VP.n13 48.7492
R220 VP.n22 VP.n15 48.7492
R221 VP.n55 VP.n54 32.2376
R222 VP.n66 VP.n3 32.2376
R223 VP.n33 VP.n13 32.2376
R224 VP.n22 VP.n21 32.2376
R225 VP.n48 VP.n9 24.4675
R226 VP.n50 VP.n49 24.4675
R227 VP.n54 VP.n53 24.4675
R228 VP.n59 VP.n5 24.4675
R229 VP.n62 VP.n61 24.4675
R230 VP.n67 VP.n66 24.4675
R231 VP.n69 VP.n1 24.4675
R232 VP.n74 VP.n73 24.4675
R233 VP.n41 VP.n40 24.4675
R234 VP.n34 VP.n33 24.4675
R235 VP.n36 VP.n11 24.4675
R236 VP.n26 VP.n15 24.4675
R237 VP.n29 VP.n28 24.4675
R238 VP.n21 VP.n20 24.4675
R239 VP.n50 VP.n7 20.5528
R240 VP.n69 VP.n68 20.5528
R241 VP.n36 VP.n35 20.5528
R242 VP.n44 VP.n9 20.0634
R243 VP.n75 VP.n74 20.0634
R244 VP.n42 VP.n41 20.0634
R245 VP.n19 VP.n18 13.2957
R246 VP.n60 VP.n59 12.234
R247 VP.n61 VP.n60 12.234
R248 VP.n27 VP.n26 12.234
R249 VP.n28 VP.n27 12.234
R250 VP.n53 VP.n7 3.91522
R251 VP.n68 VP.n67 3.91522
R252 VP.n35 VP.n34 3.91522
R253 VP.n20 VP.n17 3.91522
R254 VP.n43 VP.n10 0.278367
R255 VP.n46 VP.n45 0.278367
R256 VP.n76 VP.n0 0.278367
R257 VP.n19 VP.n16 0.189894
R258 VP.n23 VP.n16 0.189894
R259 VP.n24 VP.n23 0.189894
R260 VP.n25 VP.n24 0.189894
R261 VP.n25 VP.n14 0.189894
R262 VP.n30 VP.n14 0.189894
R263 VP.n31 VP.n30 0.189894
R264 VP.n32 VP.n31 0.189894
R265 VP.n32 VP.n12 0.189894
R266 VP.n37 VP.n12 0.189894
R267 VP.n38 VP.n37 0.189894
R268 VP.n39 VP.n38 0.189894
R269 VP.n39 VP.n10 0.189894
R270 VP.n47 VP.n46 0.189894
R271 VP.n47 VP.n8 0.189894
R272 VP.n51 VP.n8 0.189894
R273 VP.n52 VP.n51 0.189894
R274 VP.n52 VP.n6 0.189894
R275 VP.n56 VP.n6 0.189894
R276 VP.n57 VP.n56 0.189894
R277 VP.n58 VP.n57 0.189894
R278 VP.n58 VP.n4 0.189894
R279 VP.n63 VP.n4 0.189894
R280 VP.n64 VP.n63 0.189894
R281 VP.n65 VP.n64 0.189894
R282 VP.n65 VP.n2 0.189894
R283 VP.n70 VP.n2 0.189894
R284 VP.n71 VP.n70 0.189894
R285 VP.n72 VP.n71 0.189894
R286 VP.n72 VP.n0 0.189894
R287 VP VP.n76 0.153454
R288 VDD1.n1 VDD1.t8 75.9147
R289 VDD1.n3 VDD1.t3 75.9146
R290 VDD1.n5 VDD1.n4 72.7293
R291 VDD1.n1 VDD1.n0 71.2784
R292 VDD1.n7 VDD1.n6 71.2782
R293 VDD1.n3 VDD1.n2 71.2782
R294 VDD1.n7 VDD1.n5 45.5074
R295 VDD1.n6 VDD1.t7 2.62823
R296 VDD1.n6 VDD1.t2 2.62823
R297 VDD1.n0 VDD1.t5 2.62823
R298 VDD1.n0 VDD1.t1 2.62823
R299 VDD1.n4 VDD1.t4 2.62823
R300 VDD1.n4 VDD1.t0 2.62823
R301 VDD1.n2 VDD1.t9 2.62823
R302 VDD1.n2 VDD1.t6 2.62823
R303 VDD1 VDD1.n7 1.44878
R304 VDD1 VDD1.n1 0.560845
R305 VDD1.n5 VDD1.n3 0.447309
R306 B.n569 B.n78 585
R307 B.n571 B.n570 585
R308 B.n572 B.n77 585
R309 B.n574 B.n573 585
R310 B.n575 B.n76 585
R311 B.n577 B.n576 585
R312 B.n578 B.n75 585
R313 B.n580 B.n579 585
R314 B.n581 B.n74 585
R315 B.n583 B.n582 585
R316 B.n584 B.n73 585
R317 B.n586 B.n585 585
R318 B.n587 B.n72 585
R319 B.n589 B.n588 585
R320 B.n590 B.n71 585
R321 B.n592 B.n591 585
R322 B.n593 B.n70 585
R323 B.n595 B.n594 585
R324 B.n596 B.n69 585
R325 B.n598 B.n597 585
R326 B.n599 B.n68 585
R327 B.n601 B.n600 585
R328 B.n602 B.n67 585
R329 B.n604 B.n603 585
R330 B.n605 B.n66 585
R331 B.n607 B.n606 585
R332 B.n608 B.n65 585
R333 B.n610 B.n609 585
R334 B.n611 B.n64 585
R335 B.n613 B.n612 585
R336 B.n614 B.n63 585
R337 B.n616 B.n615 585
R338 B.n617 B.n62 585
R339 B.n619 B.n618 585
R340 B.n620 B.n61 585
R341 B.n622 B.n621 585
R342 B.n623 B.n60 585
R343 B.n625 B.n624 585
R344 B.n626 B.n59 585
R345 B.n628 B.n627 585
R346 B.n629 B.n58 585
R347 B.n631 B.n630 585
R348 B.n632 B.n55 585
R349 B.n635 B.n634 585
R350 B.n636 B.n54 585
R351 B.n638 B.n637 585
R352 B.n639 B.n53 585
R353 B.n641 B.n640 585
R354 B.n642 B.n52 585
R355 B.n644 B.n643 585
R356 B.n645 B.n51 585
R357 B.n647 B.n646 585
R358 B.n649 B.n648 585
R359 B.n650 B.n47 585
R360 B.n652 B.n651 585
R361 B.n653 B.n46 585
R362 B.n655 B.n654 585
R363 B.n656 B.n45 585
R364 B.n658 B.n657 585
R365 B.n659 B.n44 585
R366 B.n661 B.n660 585
R367 B.n662 B.n43 585
R368 B.n664 B.n663 585
R369 B.n665 B.n42 585
R370 B.n667 B.n666 585
R371 B.n668 B.n41 585
R372 B.n670 B.n669 585
R373 B.n671 B.n40 585
R374 B.n673 B.n672 585
R375 B.n674 B.n39 585
R376 B.n676 B.n675 585
R377 B.n677 B.n38 585
R378 B.n679 B.n678 585
R379 B.n680 B.n37 585
R380 B.n682 B.n681 585
R381 B.n683 B.n36 585
R382 B.n685 B.n684 585
R383 B.n686 B.n35 585
R384 B.n688 B.n687 585
R385 B.n689 B.n34 585
R386 B.n691 B.n690 585
R387 B.n692 B.n33 585
R388 B.n694 B.n693 585
R389 B.n695 B.n32 585
R390 B.n697 B.n696 585
R391 B.n698 B.n31 585
R392 B.n700 B.n699 585
R393 B.n701 B.n30 585
R394 B.n703 B.n702 585
R395 B.n704 B.n29 585
R396 B.n706 B.n705 585
R397 B.n707 B.n28 585
R398 B.n709 B.n708 585
R399 B.n710 B.n27 585
R400 B.n712 B.n711 585
R401 B.n568 B.n567 585
R402 B.n566 B.n79 585
R403 B.n565 B.n564 585
R404 B.n563 B.n80 585
R405 B.n562 B.n561 585
R406 B.n560 B.n81 585
R407 B.n559 B.n558 585
R408 B.n557 B.n82 585
R409 B.n556 B.n555 585
R410 B.n554 B.n83 585
R411 B.n553 B.n552 585
R412 B.n551 B.n84 585
R413 B.n550 B.n549 585
R414 B.n548 B.n85 585
R415 B.n547 B.n546 585
R416 B.n545 B.n86 585
R417 B.n544 B.n543 585
R418 B.n542 B.n87 585
R419 B.n541 B.n540 585
R420 B.n539 B.n88 585
R421 B.n538 B.n537 585
R422 B.n536 B.n89 585
R423 B.n535 B.n534 585
R424 B.n533 B.n90 585
R425 B.n532 B.n531 585
R426 B.n530 B.n91 585
R427 B.n529 B.n528 585
R428 B.n527 B.n92 585
R429 B.n526 B.n525 585
R430 B.n524 B.n93 585
R431 B.n523 B.n522 585
R432 B.n521 B.n94 585
R433 B.n520 B.n519 585
R434 B.n518 B.n95 585
R435 B.n517 B.n516 585
R436 B.n515 B.n96 585
R437 B.n514 B.n513 585
R438 B.n512 B.n97 585
R439 B.n511 B.n510 585
R440 B.n509 B.n98 585
R441 B.n508 B.n507 585
R442 B.n506 B.n99 585
R443 B.n505 B.n504 585
R444 B.n503 B.n100 585
R445 B.n502 B.n501 585
R446 B.n500 B.n101 585
R447 B.n499 B.n498 585
R448 B.n497 B.n102 585
R449 B.n496 B.n495 585
R450 B.n494 B.n103 585
R451 B.n493 B.n492 585
R452 B.n491 B.n104 585
R453 B.n490 B.n489 585
R454 B.n488 B.n105 585
R455 B.n487 B.n486 585
R456 B.n485 B.n106 585
R457 B.n484 B.n483 585
R458 B.n482 B.n107 585
R459 B.n481 B.n480 585
R460 B.n479 B.n108 585
R461 B.n478 B.n477 585
R462 B.n476 B.n109 585
R463 B.n475 B.n474 585
R464 B.n473 B.n110 585
R465 B.n472 B.n471 585
R466 B.n470 B.n111 585
R467 B.n469 B.n468 585
R468 B.n467 B.n112 585
R469 B.n466 B.n465 585
R470 B.n464 B.n113 585
R471 B.n463 B.n462 585
R472 B.n461 B.n114 585
R473 B.n460 B.n459 585
R474 B.n458 B.n115 585
R475 B.n457 B.n456 585
R476 B.n455 B.n116 585
R477 B.n454 B.n453 585
R478 B.n452 B.n117 585
R479 B.n451 B.n450 585
R480 B.n449 B.n118 585
R481 B.n448 B.n447 585
R482 B.n446 B.n119 585
R483 B.n445 B.n444 585
R484 B.n443 B.n120 585
R485 B.n442 B.n441 585
R486 B.n440 B.n121 585
R487 B.n439 B.n438 585
R488 B.n437 B.n122 585
R489 B.n436 B.n435 585
R490 B.n434 B.n123 585
R491 B.n433 B.n432 585
R492 B.n431 B.n124 585
R493 B.n430 B.n429 585
R494 B.n428 B.n125 585
R495 B.n427 B.n426 585
R496 B.n425 B.n126 585
R497 B.n424 B.n423 585
R498 B.n422 B.n127 585
R499 B.n421 B.n420 585
R500 B.n277 B.n276 585
R501 B.n278 B.n179 585
R502 B.n280 B.n279 585
R503 B.n281 B.n178 585
R504 B.n283 B.n282 585
R505 B.n284 B.n177 585
R506 B.n286 B.n285 585
R507 B.n287 B.n176 585
R508 B.n289 B.n288 585
R509 B.n290 B.n175 585
R510 B.n292 B.n291 585
R511 B.n293 B.n174 585
R512 B.n295 B.n294 585
R513 B.n296 B.n173 585
R514 B.n298 B.n297 585
R515 B.n299 B.n172 585
R516 B.n301 B.n300 585
R517 B.n302 B.n171 585
R518 B.n304 B.n303 585
R519 B.n305 B.n170 585
R520 B.n307 B.n306 585
R521 B.n308 B.n169 585
R522 B.n310 B.n309 585
R523 B.n311 B.n168 585
R524 B.n313 B.n312 585
R525 B.n314 B.n167 585
R526 B.n316 B.n315 585
R527 B.n317 B.n166 585
R528 B.n319 B.n318 585
R529 B.n320 B.n165 585
R530 B.n322 B.n321 585
R531 B.n323 B.n164 585
R532 B.n325 B.n324 585
R533 B.n326 B.n163 585
R534 B.n328 B.n327 585
R535 B.n329 B.n162 585
R536 B.n331 B.n330 585
R537 B.n332 B.n161 585
R538 B.n334 B.n333 585
R539 B.n335 B.n160 585
R540 B.n337 B.n336 585
R541 B.n338 B.n159 585
R542 B.n340 B.n339 585
R543 B.n342 B.n341 585
R544 B.n343 B.n155 585
R545 B.n345 B.n344 585
R546 B.n346 B.n154 585
R547 B.n348 B.n347 585
R548 B.n349 B.n153 585
R549 B.n351 B.n350 585
R550 B.n352 B.n152 585
R551 B.n354 B.n353 585
R552 B.n356 B.n149 585
R553 B.n358 B.n357 585
R554 B.n359 B.n148 585
R555 B.n361 B.n360 585
R556 B.n362 B.n147 585
R557 B.n364 B.n363 585
R558 B.n365 B.n146 585
R559 B.n367 B.n366 585
R560 B.n368 B.n145 585
R561 B.n370 B.n369 585
R562 B.n371 B.n144 585
R563 B.n373 B.n372 585
R564 B.n374 B.n143 585
R565 B.n376 B.n375 585
R566 B.n377 B.n142 585
R567 B.n379 B.n378 585
R568 B.n380 B.n141 585
R569 B.n382 B.n381 585
R570 B.n383 B.n140 585
R571 B.n385 B.n384 585
R572 B.n386 B.n139 585
R573 B.n388 B.n387 585
R574 B.n389 B.n138 585
R575 B.n391 B.n390 585
R576 B.n392 B.n137 585
R577 B.n394 B.n393 585
R578 B.n395 B.n136 585
R579 B.n397 B.n396 585
R580 B.n398 B.n135 585
R581 B.n400 B.n399 585
R582 B.n401 B.n134 585
R583 B.n403 B.n402 585
R584 B.n404 B.n133 585
R585 B.n406 B.n405 585
R586 B.n407 B.n132 585
R587 B.n409 B.n408 585
R588 B.n410 B.n131 585
R589 B.n412 B.n411 585
R590 B.n413 B.n130 585
R591 B.n415 B.n414 585
R592 B.n416 B.n129 585
R593 B.n418 B.n417 585
R594 B.n419 B.n128 585
R595 B.n275 B.n180 585
R596 B.n274 B.n273 585
R597 B.n272 B.n181 585
R598 B.n271 B.n270 585
R599 B.n269 B.n182 585
R600 B.n268 B.n267 585
R601 B.n266 B.n183 585
R602 B.n265 B.n264 585
R603 B.n263 B.n184 585
R604 B.n262 B.n261 585
R605 B.n260 B.n185 585
R606 B.n259 B.n258 585
R607 B.n257 B.n186 585
R608 B.n256 B.n255 585
R609 B.n254 B.n187 585
R610 B.n253 B.n252 585
R611 B.n251 B.n188 585
R612 B.n250 B.n249 585
R613 B.n248 B.n189 585
R614 B.n247 B.n246 585
R615 B.n245 B.n190 585
R616 B.n244 B.n243 585
R617 B.n242 B.n191 585
R618 B.n241 B.n240 585
R619 B.n239 B.n192 585
R620 B.n238 B.n237 585
R621 B.n236 B.n193 585
R622 B.n235 B.n234 585
R623 B.n233 B.n194 585
R624 B.n232 B.n231 585
R625 B.n230 B.n195 585
R626 B.n229 B.n228 585
R627 B.n227 B.n196 585
R628 B.n226 B.n225 585
R629 B.n224 B.n197 585
R630 B.n223 B.n222 585
R631 B.n221 B.n198 585
R632 B.n220 B.n219 585
R633 B.n218 B.n199 585
R634 B.n217 B.n216 585
R635 B.n215 B.n200 585
R636 B.n214 B.n213 585
R637 B.n212 B.n201 585
R638 B.n211 B.n210 585
R639 B.n209 B.n202 585
R640 B.n208 B.n207 585
R641 B.n206 B.n203 585
R642 B.n205 B.n204 585
R643 B.n2 B.n0 585
R644 B.n785 B.n1 585
R645 B.n784 B.n783 585
R646 B.n782 B.n3 585
R647 B.n781 B.n780 585
R648 B.n779 B.n4 585
R649 B.n778 B.n777 585
R650 B.n776 B.n5 585
R651 B.n775 B.n774 585
R652 B.n773 B.n6 585
R653 B.n772 B.n771 585
R654 B.n770 B.n7 585
R655 B.n769 B.n768 585
R656 B.n767 B.n8 585
R657 B.n766 B.n765 585
R658 B.n764 B.n9 585
R659 B.n763 B.n762 585
R660 B.n761 B.n10 585
R661 B.n760 B.n759 585
R662 B.n758 B.n11 585
R663 B.n757 B.n756 585
R664 B.n755 B.n12 585
R665 B.n754 B.n753 585
R666 B.n752 B.n13 585
R667 B.n751 B.n750 585
R668 B.n749 B.n14 585
R669 B.n748 B.n747 585
R670 B.n746 B.n15 585
R671 B.n745 B.n744 585
R672 B.n743 B.n16 585
R673 B.n742 B.n741 585
R674 B.n740 B.n17 585
R675 B.n739 B.n738 585
R676 B.n737 B.n18 585
R677 B.n736 B.n735 585
R678 B.n734 B.n19 585
R679 B.n733 B.n732 585
R680 B.n731 B.n20 585
R681 B.n730 B.n729 585
R682 B.n728 B.n21 585
R683 B.n727 B.n726 585
R684 B.n725 B.n22 585
R685 B.n724 B.n723 585
R686 B.n722 B.n23 585
R687 B.n721 B.n720 585
R688 B.n719 B.n24 585
R689 B.n718 B.n717 585
R690 B.n716 B.n25 585
R691 B.n715 B.n714 585
R692 B.n713 B.n26 585
R693 B.n787 B.n786 585
R694 B.n276 B.n275 535.745
R695 B.n713 B.n712 535.745
R696 B.n420 B.n419 535.745
R697 B.n569 B.n568 535.745
R698 B.n150 B.t3 355.976
R699 B.n156 B.t9 355.976
R700 B.n48 B.t6 355.976
R701 B.n56 B.t0 355.976
R702 B.n275 B.n274 163.367
R703 B.n274 B.n181 163.367
R704 B.n270 B.n181 163.367
R705 B.n270 B.n269 163.367
R706 B.n269 B.n268 163.367
R707 B.n268 B.n183 163.367
R708 B.n264 B.n183 163.367
R709 B.n264 B.n263 163.367
R710 B.n263 B.n262 163.367
R711 B.n262 B.n185 163.367
R712 B.n258 B.n185 163.367
R713 B.n258 B.n257 163.367
R714 B.n257 B.n256 163.367
R715 B.n256 B.n187 163.367
R716 B.n252 B.n187 163.367
R717 B.n252 B.n251 163.367
R718 B.n251 B.n250 163.367
R719 B.n250 B.n189 163.367
R720 B.n246 B.n189 163.367
R721 B.n246 B.n245 163.367
R722 B.n245 B.n244 163.367
R723 B.n244 B.n191 163.367
R724 B.n240 B.n191 163.367
R725 B.n240 B.n239 163.367
R726 B.n239 B.n238 163.367
R727 B.n238 B.n193 163.367
R728 B.n234 B.n193 163.367
R729 B.n234 B.n233 163.367
R730 B.n233 B.n232 163.367
R731 B.n232 B.n195 163.367
R732 B.n228 B.n195 163.367
R733 B.n228 B.n227 163.367
R734 B.n227 B.n226 163.367
R735 B.n226 B.n197 163.367
R736 B.n222 B.n197 163.367
R737 B.n222 B.n221 163.367
R738 B.n221 B.n220 163.367
R739 B.n220 B.n199 163.367
R740 B.n216 B.n199 163.367
R741 B.n216 B.n215 163.367
R742 B.n215 B.n214 163.367
R743 B.n214 B.n201 163.367
R744 B.n210 B.n201 163.367
R745 B.n210 B.n209 163.367
R746 B.n209 B.n208 163.367
R747 B.n208 B.n203 163.367
R748 B.n204 B.n203 163.367
R749 B.n204 B.n2 163.367
R750 B.n786 B.n2 163.367
R751 B.n786 B.n785 163.367
R752 B.n785 B.n784 163.367
R753 B.n784 B.n3 163.367
R754 B.n780 B.n3 163.367
R755 B.n780 B.n779 163.367
R756 B.n779 B.n778 163.367
R757 B.n778 B.n5 163.367
R758 B.n774 B.n5 163.367
R759 B.n774 B.n773 163.367
R760 B.n773 B.n772 163.367
R761 B.n772 B.n7 163.367
R762 B.n768 B.n7 163.367
R763 B.n768 B.n767 163.367
R764 B.n767 B.n766 163.367
R765 B.n766 B.n9 163.367
R766 B.n762 B.n9 163.367
R767 B.n762 B.n761 163.367
R768 B.n761 B.n760 163.367
R769 B.n760 B.n11 163.367
R770 B.n756 B.n11 163.367
R771 B.n756 B.n755 163.367
R772 B.n755 B.n754 163.367
R773 B.n754 B.n13 163.367
R774 B.n750 B.n13 163.367
R775 B.n750 B.n749 163.367
R776 B.n749 B.n748 163.367
R777 B.n748 B.n15 163.367
R778 B.n744 B.n15 163.367
R779 B.n744 B.n743 163.367
R780 B.n743 B.n742 163.367
R781 B.n742 B.n17 163.367
R782 B.n738 B.n17 163.367
R783 B.n738 B.n737 163.367
R784 B.n737 B.n736 163.367
R785 B.n736 B.n19 163.367
R786 B.n732 B.n19 163.367
R787 B.n732 B.n731 163.367
R788 B.n731 B.n730 163.367
R789 B.n730 B.n21 163.367
R790 B.n726 B.n21 163.367
R791 B.n726 B.n725 163.367
R792 B.n725 B.n724 163.367
R793 B.n724 B.n23 163.367
R794 B.n720 B.n23 163.367
R795 B.n720 B.n719 163.367
R796 B.n719 B.n718 163.367
R797 B.n718 B.n25 163.367
R798 B.n714 B.n25 163.367
R799 B.n714 B.n713 163.367
R800 B.n276 B.n179 163.367
R801 B.n280 B.n179 163.367
R802 B.n281 B.n280 163.367
R803 B.n282 B.n281 163.367
R804 B.n282 B.n177 163.367
R805 B.n286 B.n177 163.367
R806 B.n287 B.n286 163.367
R807 B.n288 B.n287 163.367
R808 B.n288 B.n175 163.367
R809 B.n292 B.n175 163.367
R810 B.n293 B.n292 163.367
R811 B.n294 B.n293 163.367
R812 B.n294 B.n173 163.367
R813 B.n298 B.n173 163.367
R814 B.n299 B.n298 163.367
R815 B.n300 B.n299 163.367
R816 B.n300 B.n171 163.367
R817 B.n304 B.n171 163.367
R818 B.n305 B.n304 163.367
R819 B.n306 B.n305 163.367
R820 B.n306 B.n169 163.367
R821 B.n310 B.n169 163.367
R822 B.n311 B.n310 163.367
R823 B.n312 B.n311 163.367
R824 B.n312 B.n167 163.367
R825 B.n316 B.n167 163.367
R826 B.n317 B.n316 163.367
R827 B.n318 B.n317 163.367
R828 B.n318 B.n165 163.367
R829 B.n322 B.n165 163.367
R830 B.n323 B.n322 163.367
R831 B.n324 B.n323 163.367
R832 B.n324 B.n163 163.367
R833 B.n328 B.n163 163.367
R834 B.n329 B.n328 163.367
R835 B.n330 B.n329 163.367
R836 B.n330 B.n161 163.367
R837 B.n334 B.n161 163.367
R838 B.n335 B.n334 163.367
R839 B.n336 B.n335 163.367
R840 B.n336 B.n159 163.367
R841 B.n340 B.n159 163.367
R842 B.n341 B.n340 163.367
R843 B.n341 B.n155 163.367
R844 B.n345 B.n155 163.367
R845 B.n346 B.n345 163.367
R846 B.n347 B.n346 163.367
R847 B.n347 B.n153 163.367
R848 B.n351 B.n153 163.367
R849 B.n352 B.n351 163.367
R850 B.n353 B.n352 163.367
R851 B.n353 B.n149 163.367
R852 B.n358 B.n149 163.367
R853 B.n359 B.n358 163.367
R854 B.n360 B.n359 163.367
R855 B.n360 B.n147 163.367
R856 B.n364 B.n147 163.367
R857 B.n365 B.n364 163.367
R858 B.n366 B.n365 163.367
R859 B.n366 B.n145 163.367
R860 B.n370 B.n145 163.367
R861 B.n371 B.n370 163.367
R862 B.n372 B.n371 163.367
R863 B.n372 B.n143 163.367
R864 B.n376 B.n143 163.367
R865 B.n377 B.n376 163.367
R866 B.n378 B.n377 163.367
R867 B.n378 B.n141 163.367
R868 B.n382 B.n141 163.367
R869 B.n383 B.n382 163.367
R870 B.n384 B.n383 163.367
R871 B.n384 B.n139 163.367
R872 B.n388 B.n139 163.367
R873 B.n389 B.n388 163.367
R874 B.n390 B.n389 163.367
R875 B.n390 B.n137 163.367
R876 B.n394 B.n137 163.367
R877 B.n395 B.n394 163.367
R878 B.n396 B.n395 163.367
R879 B.n396 B.n135 163.367
R880 B.n400 B.n135 163.367
R881 B.n401 B.n400 163.367
R882 B.n402 B.n401 163.367
R883 B.n402 B.n133 163.367
R884 B.n406 B.n133 163.367
R885 B.n407 B.n406 163.367
R886 B.n408 B.n407 163.367
R887 B.n408 B.n131 163.367
R888 B.n412 B.n131 163.367
R889 B.n413 B.n412 163.367
R890 B.n414 B.n413 163.367
R891 B.n414 B.n129 163.367
R892 B.n418 B.n129 163.367
R893 B.n419 B.n418 163.367
R894 B.n420 B.n127 163.367
R895 B.n424 B.n127 163.367
R896 B.n425 B.n424 163.367
R897 B.n426 B.n425 163.367
R898 B.n426 B.n125 163.367
R899 B.n430 B.n125 163.367
R900 B.n431 B.n430 163.367
R901 B.n432 B.n431 163.367
R902 B.n432 B.n123 163.367
R903 B.n436 B.n123 163.367
R904 B.n437 B.n436 163.367
R905 B.n438 B.n437 163.367
R906 B.n438 B.n121 163.367
R907 B.n442 B.n121 163.367
R908 B.n443 B.n442 163.367
R909 B.n444 B.n443 163.367
R910 B.n444 B.n119 163.367
R911 B.n448 B.n119 163.367
R912 B.n449 B.n448 163.367
R913 B.n450 B.n449 163.367
R914 B.n450 B.n117 163.367
R915 B.n454 B.n117 163.367
R916 B.n455 B.n454 163.367
R917 B.n456 B.n455 163.367
R918 B.n456 B.n115 163.367
R919 B.n460 B.n115 163.367
R920 B.n461 B.n460 163.367
R921 B.n462 B.n461 163.367
R922 B.n462 B.n113 163.367
R923 B.n466 B.n113 163.367
R924 B.n467 B.n466 163.367
R925 B.n468 B.n467 163.367
R926 B.n468 B.n111 163.367
R927 B.n472 B.n111 163.367
R928 B.n473 B.n472 163.367
R929 B.n474 B.n473 163.367
R930 B.n474 B.n109 163.367
R931 B.n478 B.n109 163.367
R932 B.n479 B.n478 163.367
R933 B.n480 B.n479 163.367
R934 B.n480 B.n107 163.367
R935 B.n484 B.n107 163.367
R936 B.n485 B.n484 163.367
R937 B.n486 B.n485 163.367
R938 B.n486 B.n105 163.367
R939 B.n490 B.n105 163.367
R940 B.n491 B.n490 163.367
R941 B.n492 B.n491 163.367
R942 B.n492 B.n103 163.367
R943 B.n496 B.n103 163.367
R944 B.n497 B.n496 163.367
R945 B.n498 B.n497 163.367
R946 B.n498 B.n101 163.367
R947 B.n502 B.n101 163.367
R948 B.n503 B.n502 163.367
R949 B.n504 B.n503 163.367
R950 B.n504 B.n99 163.367
R951 B.n508 B.n99 163.367
R952 B.n509 B.n508 163.367
R953 B.n510 B.n509 163.367
R954 B.n510 B.n97 163.367
R955 B.n514 B.n97 163.367
R956 B.n515 B.n514 163.367
R957 B.n516 B.n515 163.367
R958 B.n516 B.n95 163.367
R959 B.n520 B.n95 163.367
R960 B.n521 B.n520 163.367
R961 B.n522 B.n521 163.367
R962 B.n522 B.n93 163.367
R963 B.n526 B.n93 163.367
R964 B.n527 B.n526 163.367
R965 B.n528 B.n527 163.367
R966 B.n528 B.n91 163.367
R967 B.n532 B.n91 163.367
R968 B.n533 B.n532 163.367
R969 B.n534 B.n533 163.367
R970 B.n534 B.n89 163.367
R971 B.n538 B.n89 163.367
R972 B.n539 B.n538 163.367
R973 B.n540 B.n539 163.367
R974 B.n540 B.n87 163.367
R975 B.n544 B.n87 163.367
R976 B.n545 B.n544 163.367
R977 B.n546 B.n545 163.367
R978 B.n546 B.n85 163.367
R979 B.n550 B.n85 163.367
R980 B.n551 B.n550 163.367
R981 B.n552 B.n551 163.367
R982 B.n552 B.n83 163.367
R983 B.n556 B.n83 163.367
R984 B.n557 B.n556 163.367
R985 B.n558 B.n557 163.367
R986 B.n558 B.n81 163.367
R987 B.n562 B.n81 163.367
R988 B.n563 B.n562 163.367
R989 B.n564 B.n563 163.367
R990 B.n564 B.n79 163.367
R991 B.n568 B.n79 163.367
R992 B.n712 B.n27 163.367
R993 B.n708 B.n27 163.367
R994 B.n708 B.n707 163.367
R995 B.n707 B.n706 163.367
R996 B.n706 B.n29 163.367
R997 B.n702 B.n29 163.367
R998 B.n702 B.n701 163.367
R999 B.n701 B.n700 163.367
R1000 B.n700 B.n31 163.367
R1001 B.n696 B.n31 163.367
R1002 B.n696 B.n695 163.367
R1003 B.n695 B.n694 163.367
R1004 B.n694 B.n33 163.367
R1005 B.n690 B.n33 163.367
R1006 B.n690 B.n689 163.367
R1007 B.n689 B.n688 163.367
R1008 B.n688 B.n35 163.367
R1009 B.n684 B.n35 163.367
R1010 B.n684 B.n683 163.367
R1011 B.n683 B.n682 163.367
R1012 B.n682 B.n37 163.367
R1013 B.n678 B.n37 163.367
R1014 B.n678 B.n677 163.367
R1015 B.n677 B.n676 163.367
R1016 B.n676 B.n39 163.367
R1017 B.n672 B.n39 163.367
R1018 B.n672 B.n671 163.367
R1019 B.n671 B.n670 163.367
R1020 B.n670 B.n41 163.367
R1021 B.n666 B.n41 163.367
R1022 B.n666 B.n665 163.367
R1023 B.n665 B.n664 163.367
R1024 B.n664 B.n43 163.367
R1025 B.n660 B.n43 163.367
R1026 B.n660 B.n659 163.367
R1027 B.n659 B.n658 163.367
R1028 B.n658 B.n45 163.367
R1029 B.n654 B.n45 163.367
R1030 B.n654 B.n653 163.367
R1031 B.n653 B.n652 163.367
R1032 B.n652 B.n47 163.367
R1033 B.n648 B.n47 163.367
R1034 B.n648 B.n647 163.367
R1035 B.n647 B.n51 163.367
R1036 B.n643 B.n51 163.367
R1037 B.n643 B.n642 163.367
R1038 B.n642 B.n641 163.367
R1039 B.n641 B.n53 163.367
R1040 B.n637 B.n53 163.367
R1041 B.n637 B.n636 163.367
R1042 B.n636 B.n635 163.367
R1043 B.n635 B.n55 163.367
R1044 B.n630 B.n55 163.367
R1045 B.n630 B.n629 163.367
R1046 B.n629 B.n628 163.367
R1047 B.n628 B.n59 163.367
R1048 B.n624 B.n59 163.367
R1049 B.n624 B.n623 163.367
R1050 B.n623 B.n622 163.367
R1051 B.n622 B.n61 163.367
R1052 B.n618 B.n61 163.367
R1053 B.n618 B.n617 163.367
R1054 B.n617 B.n616 163.367
R1055 B.n616 B.n63 163.367
R1056 B.n612 B.n63 163.367
R1057 B.n612 B.n611 163.367
R1058 B.n611 B.n610 163.367
R1059 B.n610 B.n65 163.367
R1060 B.n606 B.n65 163.367
R1061 B.n606 B.n605 163.367
R1062 B.n605 B.n604 163.367
R1063 B.n604 B.n67 163.367
R1064 B.n600 B.n67 163.367
R1065 B.n600 B.n599 163.367
R1066 B.n599 B.n598 163.367
R1067 B.n598 B.n69 163.367
R1068 B.n594 B.n69 163.367
R1069 B.n594 B.n593 163.367
R1070 B.n593 B.n592 163.367
R1071 B.n592 B.n71 163.367
R1072 B.n588 B.n71 163.367
R1073 B.n588 B.n587 163.367
R1074 B.n587 B.n586 163.367
R1075 B.n586 B.n73 163.367
R1076 B.n582 B.n73 163.367
R1077 B.n582 B.n581 163.367
R1078 B.n581 B.n580 163.367
R1079 B.n580 B.n75 163.367
R1080 B.n576 B.n75 163.367
R1081 B.n576 B.n575 163.367
R1082 B.n575 B.n574 163.367
R1083 B.n574 B.n77 163.367
R1084 B.n570 B.n77 163.367
R1085 B.n570 B.n569 163.367
R1086 B.n150 B.t5 154.732
R1087 B.n56 B.t1 154.732
R1088 B.n156 B.t11 154.716
R1089 B.n48 B.t7 154.716
R1090 B.n151 B.t4 109.543
R1091 B.n57 B.t2 109.543
R1092 B.n157 B.t10 109.528
R1093 B.n49 B.t8 109.528
R1094 B.n355 B.n151 59.5399
R1095 B.n158 B.n157 59.5399
R1096 B.n50 B.n49 59.5399
R1097 B.n633 B.n57 59.5399
R1098 B.n151 B.n150 45.1884
R1099 B.n157 B.n156 45.1884
R1100 B.n49 B.n48 45.1884
R1101 B.n57 B.n56 45.1884
R1102 B.n711 B.n26 34.8103
R1103 B.n567 B.n78 34.8103
R1104 B.n421 B.n128 34.8103
R1105 B.n277 B.n180 34.8103
R1106 B B.n787 18.0485
R1107 B.n711 B.n710 10.6151
R1108 B.n710 B.n709 10.6151
R1109 B.n709 B.n28 10.6151
R1110 B.n705 B.n28 10.6151
R1111 B.n705 B.n704 10.6151
R1112 B.n704 B.n703 10.6151
R1113 B.n703 B.n30 10.6151
R1114 B.n699 B.n30 10.6151
R1115 B.n699 B.n698 10.6151
R1116 B.n698 B.n697 10.6151
R1117 B.n697 B.n32 10.6151
R1118 B.n693 B.n32 10.6151
R1119 B.n693 B.n692 10.6151
R1120 B.n692 B.n691 10.6151
R1121 B.n691 B.n34 10.6151
R1122 B.n687 B.n34 10.6151
R1123 B.n687 B.n686 10.6151
R1124 B.n686 B.n685 10.6151
R1125 B.n685 B.n36 10.6151
R1126 B.n681 B.n36 10.6151
R1127 B.n681 B.n680 10.6151
R1128 B.n680 B.n679 10.6151
R1129 B.n679 B.n38 10.6151
R1130 B.n675 B.n38 10.6151
R1131 B.n675 B.n674 10.6151
R1132 B.n674 B.n673 10.6151
R1133 B.n673 B.n40 10.6151
R1134 B.n669 B.n40 10.6151
R1135 B.n669 B.n668 10.6151
R1136 B.n668 B.n667 10.6151
R1137 B.n667 B.n42 10.6151
R1138 B.n663 B.n42 10.6151
R1139 B.n663 B.n662 10.6151
R1140 B.n662 B.n661 10.6151
R1141 B.n661 B.n44 10.6151
R1142 B.n657 B.n44 10.6151
R1143 B.n657 B.n656 10.6151
R1144 B.n656 B.n655 10.6151
R1145 B.n655 B.n46 10.6151
R1146 B.n651 B.n46 10.6151
R1147 B.n651 B.n650 10.6151
R1148 B.n650 B.n649 10.6151
R1149 B.n646 B.n645 10.6151
R1150 B.n645 B.n644 10.6151
R1151 B.n644 B.n52 10.6151
R1152 B.n640 B.n52 10.6151
R1153 B.n640 B.n639 10.6151
R1154 B.n639 B.n638 10.6151
R1155 B.n638 B.n54 10.6151
R1156 B.n634 B.n54 10.6151
R1157 B.n632 B.n631 10.6151
R1158 B.n631 B.n58 10.6151
R1159 B.n627 B.n58 10.6151
R1160 B.n627 B.n626 10.6151
R1161 B.n626 B.n625 10.6151
R1162 B.n625 B.n60 10.6151
R1163 B.n621 B.n60 10.6151
R1164 B.n621 B.n620 10.6151
R1165 B.n620 B.n619 10.6151
R1166 B.n619 B.n62 10.6151
R1167 B.n615 B.n62 10.6151
R1168 B.n615 B.n614 10.6151
R1169 B.n614 B.n613 10.6151
R1170 B.n613 B.n64 10.6151
R1171 B.n609 B.n64 10.6151
R1172 B.n609 B.n608 10.6151
R1173 B.n608 B.n607 10.6151
R1174 B.n607 B.n66 10.6151
R1175 B.n603 B.n66 10.6151
R1176 B.n603 B.n602 10.6151
R1177 B.n602 B.n601 10.6151
R1178 B.n601 B.n68 10.6151
R1179 B.n597 B.n68 10.6151
R1180 B.n597 B.n596 10.6151
R1181 B.n596 B.n595 10.6151
R1182 B.n595 B.n70 10.6151
R1183 B.n591 B.n70 10.6151
R1184 B.n591 B.n590 10.6151
R1185 B.n590 B.n589 10.6151
R1186 B.n589 B.n72 10.6151
R1187 B.n585 B.n72 10.6151
R1188 B.n585 B.n584 10.6151
R1189 B.n584 B.n583 10.6151
R1190 B.n583 B.n74 10.6151
R1191 B.n579 B.n74 10.6151
R1192 B.n579 B.n578 10.6151
R1193 B.n578 B.n577 10.6151
R1194 B.n577 B.n76 10.6151
R1195 B.n573 B.n76 10.6151
R1196 B.n573 B.n572 10.6151
R1197 B.n572 B.n571 10.6151
R1198 B.n571 B.n78 10.6151
R1199 B.n422 B.n421 10.6151
R1200 B.n423 B.n422 10.6151
R1201 B.n423 B.n126 10.6151
R1202 B.n427 B.n126 10.6151
R1203 B.n428 B.n427 10.6151
R1204 B.n429 B.n428 10.6151
R1205 B.n429 B.n124 10.6151
R1206 B.n433 B.n124 10.6151
R1207 B.n434 B.n433 10.6151
R1208 B.n435 B.n434 10.6151
R1209 B.n435 B.n122 10.6151
R1210 B.n439 B.n122 10.6151
R1211 B.n440 B.n439 10.6151
R1212 B.n441 B.n440 10.6151
R1213 B.n441 B.n120 10.6151
R1214 B.n445 B.n120 10.6151
R1215 B.n446 B.n445 10.6151
R1216 B.n447 B.n446 10.6151
R1217 B.n447 B.n118 10.6151
R1218 B.n451 B.n118 10.6151
R1219 B.n452 B.n451 10.6151
R1220 B.n453 B.n452 10.6151
R1221 B.n453 B.n116 10.6151
R1222 B.n457 B.n116 10.6151
R1223 B.n458 B.n457 10.6151
R1224 B.n459 B.n458 10.6151
R1225 B.n459 B.n114 10.6151
R1226 B.n463 B.n114 10.6151
R1227 B.n464 B.n463 10.6151
R1228 B.n465 B.n464 10.6151
R1229 B.n465 B.n112 10.6151
R1230 B.n469 B.n112 10.6151
R1231 B.n470 B.n469 10.6151
R1232 B.n471 B.n470 10.6151
R1233 B.n471 B.n110 10.6151
R1234 B.n475 B.n110 10.6151
R1235 B.n476 B.n475 10.6151
R1236 B.n477 B.n476 10.6151
R1237 B.n477 B.n108 10.6151
R1238 B.n481 B.n108 10.6151
R1239 B.n482 B.n481 10.6151
R1240 B.n483 B.n482 10.6151
R1241 B.n483 B.n106 10.6151
R1242 B.n487 B.n106 10.6151
R1243 B.n488 B.n487 10.6151
R1244 B.n489 B.n488 10.6151
R1245 B.n489 B.n104 10.6151
R1246 B.n493 B.n104 10.6151
R1247 B.n494 B.n493 10.6151
R1248 B.n495 B.n494 10.6151
R1249 B.n495 B.n102 10.6151
R1250 B.n499 B.n102 10.6151
R1251 B.n500 B.n499 10.6151
R1252 B.n501 B.n500 10.6151
R1253 B.n501 B.n100 10.6151
R1254 B.n505 B.n100 10.6151
R1255 B.n506 B.n505 10.6151
R1256 B.n507 B.n506 10.6151
R1257 B.n507 B.n98 10.6151
R1258 B.n511 B.n98 10.6151
R1259 B.n512 B.n511 10.6151
R1260 B.n513 B.n512 10.6151
R1261 B.n513 B.n96 10.6151
R1262 B.n517 B.n96 10.6151
R1263 B.n518 B.n517 10.6151
R1264 B.n519 B.n518 10.6151
R1265 B.n519 B.n94 10.6151
R1266 B.n523 B.n94 10.6151
R1267 B.n524 B.n523 10.6151
R1268 B.n525 B.n524 10.6151
R1269 B.n525 B.n92 10.6151
R1270 B.n529 B.n92 10.6151
R1271 B.n530 B.n529 10.6151
R1272 B.n531 B.n530 10.6151
R1273 B.n531 B.n90 10.6151
R1274 B.n535 B.n90 10.6151
R1275 B.n536 B.n535 10.6151
R1276 B.n537 B.n536 10.6151
R1277 B.n537 B.n88 10.6151
R1278 B.n541 B.n88 10.6151
R1279 B.n542 B.n541 10.6151
R1280 B.n543 B.n542 10.6151
R1281 B.n543 B.n86 10.6151
R1282 B.n547 B.n86 10.6151
R1283 B.n548 B.n547 10.6151
R1284 B.n549 B.n548 10.6151
R1285 B.n549 B.n84 10.6151
R1286 B.n553 B.n84 10.6151
R1287 B.n554 B.n553 10.6151
R1288 B.n555 B.n554 10.6151
R1289 B.n555 B.n82 10.6151
R1290 B.n559 B.n82 10.6151
R1291 B.n560 B.n559 10.6151
R1292 B.n561 B.n560 10.6151
R1293 B.n561 B.n80 10.6151
R1294 B.n565 B.n80 10.6151
R1295 B.n566 B.n565 10.6151
R1296 B.n567 B.n566 10.6151
R1297 B.n278 B.n277 10.6151
R1298 B.n279 B.n278 10.6151
R1299 B.n279 B.n178 10.6151
R1300 B.n283 B.n178 10.6151
R1301 B.n284 B.n283 10.6151
R1302 B.n285 B.n284 10.6151
R1303 B.n285 B.n176 10.6151
R1304 B.n289 B.n176 10.6151
R1305 B.n290 B.n289 10.6151
R1306 B.n291 B.n290 10.6151
R1307 B.n291 B.n174 10.6151
R1308 B.n295 B.n174 10.6151
R1309 B.n296 B.n295 10.6151
R1310 B.n297 B.n296 10.6151
R1311 B.n297 B.n172 10.6151
R1312 B.n301 B.n172 10.6151
R1313 B.n302 B.n301 10.6151
R1314 B.n303 B.n302 10.6151
R1315 B.n303 B.n170 10.6151
R1316 B.n307 B.n170 10.6151
R1317 B.n308 B.n307 10.6151
R1318 B.n309 B.n308 10.6151
R1319 B.n309 B.n168 10.6151
R1320 B.n313 B.n168 10.6151
R1321 B.n314 B.n313 10.6151
R1322 B.n315 B.n314 10.6151
R1323 B.n315 B.n166 10.6151
R1324 B.n319 B.n166 10.6151
R1325 B.n320 B.n319 10.6151
R1326 B.n321 B.n320 10.6151
R1327 B.n321 B.n164 10.6151
R1328 B.n325 B.n164 10.6151
R1329 B.n326 B.n325 10.6151
R1330 B.n327 B.n326 10.6151
R1331 B.n327 B.n162 10.6151
R1332 B.n331 B.n162 10.6151
R1333 B.n332 B.n331 10.6151
R1334 B.n333 B.n332 10.6151
R1335 B.n333 B.n160 10.6151
R1336 B.n337 B.n160 10.6151
R1337 B.n338 B.n337 10.6151
R1338 B.n339 B.n338 10.6151
R1339 B.n343 B.n342 10.6151
R1340 B.n344 B.n343 10.6151
R1341 B.n344 B.n154 10.6151
R1342 B.n348 B.n154 10.6151
R1343 B.n349 B.n348 10.6151
R1344 B.n350 B.n349 10.6151
R1345 B.n350 B.n152 10.6151
R1346 B.n354 B.n152 10.6151
R1347 B.n357 B.n356 10.6151
R1348 B.n357 B.n148 10.6151
R1349 B.n361 B.n148 10.6151
R1350 B.n362 B.n361 10.6151
R1351 B.n363 B.n362 10.6151
R1352 B.n363 B.n146 10.6151
R1353 B.n367 B.n146 10.6151
R1354 B.n368 B.n367 10.6151
R1355 B.n369 B.n368 10.6151
R1356 B.n369 B.n144 10.6151
R1357 B.n373 B.n144 10.6151
R1358 B.n374 B.n373 10.6151
R1359 B.n375 B.n374 10.6151
R1360 B.n375 B.n142 10.6151
R1361 B.n379 B.n142 10.6151
R1362 B.n380 B.n379 10.6151
R1363 B.n381 B.n380 10.6151
R1364 B.n381 B.n140 10.6151
R1365 B.n385 B.n140 10.6151
R1366 B.n386 B.n385 10.6151
R1367 B.n387 B.n386 10.6151
R1368 B.n387 B.n138 10.6151
R1369 B.n391 B.n138 10.6151
R1370 B.n392 B.n391 10.6151
R1371 B.n393 B.n392 10.6151
R1372 B.n393 B.n136 10.6151
R1373 B.n397 B.n136 10.6151
R1374 B.n398 B.n397 10.6151
R1375 B.n399 B.n398 10.6151
R1376 B.n399 B.n134 10.6151
R1377 B.n403 B.n134 10.6151
R1378 B.n404 B.n403 10.6151
R1379 B.n405 B.n404 10.6151
R1380 B.n405 B.n132 10.6151
R1381 B.n409 B.n132 10.6151
R1382 B.n410 B.n409 10.6151
R1383 B.n411 B.n410 10.6151
R1384 B.n411 B.n130 10.6151
R1385 B.n415 B.n130 10.6151
R1386 B.n416 B.n415 10.6151
R1387 B.n417 B.n416 10.6151
R1388 B.n417 B.n128 10.6151
R1389 B.n273 B.n180 10.6151
R1390 B.n273 B.n272 10.6151
R1391 B.n272 B.n271 10.6151
R1392 B.n271 B.n182 10.6151
R1393 B.n267 B.n182 10.6151
R1394 B.n267 B.n266 10.6151
R1395 B.n266 B.n265 10.6151
R1396 B.n265 B.n184 10.6151
R1397 B.n261 B.n184 10.6151
R1398 B.n261 B.n260 10.6151
R1399 B.n260 B.n259 10.6151
R1400 B.n259 B.n186 10.6151
R1401 B.n255 B.n186 10.6151
R1402 B.n255 B.n254 10.6151
R1403 B.n254 B.n253 10.6151
R1404 B.n253 B.n188 10.6151
R1405 B.n249 B.n188 10.6151
R1406 B.n249 B.n248 10.6151
R1407 B.n248 B.n247 10.6151
R1408 B.n247 B.n190 10.6151
R1409 B.n243 B.n190 10.6151
R1410 B.n243 B.n242 10.6151
R1411 B.n242 B.n241 10.6151
R1412 B.n241 B.n192 10.6151
R1413 B.n237 B.n192 10.6151
R1414 B.n237 B.n236 10.6151
R1415 B.n236 B.n235 10.6151
R1416 B.n235 B.n194 10.6151
R1417 B.n231 B.n194 10.6151
R1418 B.n231 B.n230 10.6151
R1419 B.n230 B.n229 10.6151
R1420 B.n229 B.n196 10.6151
R1421 B.n225 B.n196 10.6151
R1422 B.n225 B.n224 10.6151
R1423 B.n224 B.n223 10.6151
R1424 B.n223 B.n198 10.6151
R1425 B.n219 B.n198 10.6151
R1426 B.n219 B.n218 10.6151
R1427 B.n218 B.n217 10.6151
R1428 B.n217 B.n200 10.6151
R1429 B.n213 B.n200 10.6151
R1430 B.n213 B.n212 10.6151
R1431 B.n212 B.n211 10.6151
R1432 B.n211 B.n202 10.6151
R1433 B.n207 B.n202 10.6151
R1434 B.n207 B.n206 10.6151
R1435 B.n206 B.n205 10.6151
R1436 B.n205 B.n0 10.6151
R1437 B.n783 B.n1 10.6151
R1438 B.n783 B.n782 10.6151
R1439 B.n782 B.n781 10.6151
R1440 B.n781 B.n4 10.6151
R1441 B.n777 B.n4 10.6151
R1442 B.n777 B.n776 10.6151
R1443 B.n776 B.n775 10.6151
R1444 B.n775 B.n6 10.6151
R1445 B.n771 B.n6 10.6151
R1446 B.n771 B.n770 10.6151
R1447 B.n770 B.n769 10.6151
R1448 B.n769 B.n8 10.6151
R1449 B.n765 B.n8 10.6151
R1450 B.n765 B.n764 10.6151
R1451 B.n764 B.n763 10.6151
R1452 B.n763 B.n10 10.6151
R1453 B.n759 B.n10 10.6151
R1454 B.n759 B.n758 10.6151
R1455 B.n758 B.n757 10.6151
R1456 B.n757 B.n12 10.6151
R1457 B.n753 B.n12 10.6151
R1458 B.n753 B.n752 10.6151
R1459 B.n752 B.n751 10.6151
R1460 B.n751 B.n14 10.6151
R1461 B.n747 B.n14 10.6151
R1462 B.n747 B.n746 10.6151
R1463 B.n746 B.n745 10.6151
R1464 B.n745 B.n16 10.6151
R1465 B.n741 B.n16 10.6151
R1466 B.n741 B.n740 10.6151
R1467 B.n740 B.n739 10.6151
R1468 B.n739 B.n18 10.6151
R1469 B.n735 B.n18 10.6151
R1470 B.n735 B.n734 10.6151
R1471 B.n734 B.n733 10.6151
R1472 B.n733 B.n20 10.6151
R1473 B.n729 B.n20 10.6151
R1474 B.n729 B.n728 10.6151
R1475 B.n728 B.n727 10.6151
R1476 B.n727 B.n22 10.6151
R1477 B.n723 B.n22 10.6151
R1478 B.n723 B.n722 10.6151
R1479 B.n722 B.n721 10.6151
R1480 B.n721 B.n24 10.6151
R1481 B.n717 B.n24 10.6151
R1482 B.n717 B.n716 10.6151
R1483 B.n716 B.n715 10.6151
R1484 B.n715 B.n26 10.6151
R1485 B.n646 B.n50 6.5566
R1486 B.n634 B.n633 6.5566
R1487 B.n342 B.n158 6.5566
R1488 B.n355 B.n354 6.5566
R1489 B.n649 B.n50 4.05904
R1490 B.n633 B.n632 4.05904
R1491 B.n339 B.n158 4.05904
R1492 B.n356 B.n355 4.05904
R1493 B.n787 B.n0 2.81026
R1494 B.n787 B.n1 2.81026
C0 B VP 1.95309f
C1 VDD2 B 2.36701f
C2 VP VTAIL 10.7394f
C3 VDD2 VTAIL 10.6875f
C4 B VN 1.13503f
C5 VN VTAIL 10.724999f
C6 VDD1 VP 10.699f
C7 VDD2 VDD1 1.78411f
C8 VDD1 VN 0.151987f
C9 VP w_n3766_n3442# 8.37039f
C10 VDD2 w_n3766_n3442# 2.69915f
C11 w_n3766_n3442# VN 7.88192f
C12 B VTAIL 3.54476f
C13 VDD1 B 2.27246f
C14 VDD1 VTAIL 10.6414f
C15 B w_n3766_n3442# 9.6417f
C16 w_n3766_n3442# VTAIL 3.18728f
C17 VDD2 VP 0.507109f
C18 VP VN 7.58398f
C19 VDD2 VN 10.3478f
C20 VDD1 w_n3766_n3442# 2.58669f
C21 VDD2 VSUBS 1.918848f
C22 VDD1 VSUBS 1.712694f
C23 VTAIL VSUBS 1.171056f
C24 VN VSUBS 6.72599f
C25 VP VSUBS 3.491589f
C26 B VSUBS 4.652433f
C27 w_n3766_n3442# VSUBS 0.159483p
C28 B.n0 VSUBS 0.005443f
C29 B.n1 VSUBS 0.005443f
C30 B.n2 VSUBS 0.008608f
C31 B.n3 VSUBS 0.008608f
C32 B.n4 VSUBS 0.008608f
C33 B.n5 VSUBS 0.008608f
C34 B.n6 VSUBS 0.008608f
C35 B.n7 VSUBS 0.008608f
C36 B.n8 VSUBS 0.008608f
C37 B.n9 VSUBS 0.008608f
C38 B.n10 VSUBS 0.008608f
C39 B.n11 VSUBS 0.008608f
C40 B.n12 VSUBS 0.008608f
C41 B.n13 VSUBS 0.008608f
C42 B.n14 VSUBS 0.008608f
C43 B.n15 VSUBS 0.008608f
C44 B.n16 VSUBS 0.008608f
C45 B.n17 VSUBS 0.008608f
C46 B.n18 VSUBS 0.008608f
C47 B.n19 VSUBS 0.008608f
C48 B.n20 VSUBS 0.008608f
C49 B.n21 VSUBS 0.008608f
C50 B.n22 VSUBS 0.008608f
C51 B.n23 VSUBS 0.008608f
C52 B.n24 VSUBS 0.008608f
C53 B.n25 VSUBS 0.008608f
C54 B.n26 VSUBS 0.020373f
C55 B.n27 VSUBS 0.008608f
C56 B.n28 VSUBS 0.008608f
C57 B.n29 VSUBS 0.008608f
C58 B.n30 VSUBS 0.008608f
C59 B.n31 VSUBS 0.008608f
C60 B.n32 VSUBS 0.008608f
C61 B.n33 VSUBS 0.008608f
C62 B.n34 VSUBS 0.008608f
C63 B.n35 VSUBS 0.008608f
C64 B.n36 VSUBS 0.008608f
C65 B.n37 VSUBS 0.008608f
C66 B.n38 VSUBS 0.008608f
C67 B.n39 VSUBS 0.008608f
C68 B.n40 VSUBS 0.008608f
C69 B.n41 VSUBS 0.008608f
C70 B.n42 VSUBS 0.008608f
C71 B.n43 VSUBS 0.008608f
C72 B.n44 VSUBS 0.008608f
C73 B.n45 VSUBS 0.008608f
C74 B.n46 VSUBS 0.008608f
C75 B.n47 VSUBS 0.008608f
C76 B.t8 VSUBS 0.497302f
C77 B.t7 VSUBS 0.518618f
C78 B.t6 VSUBS 1.35737f
C79 B.n48 VSUBS 0.252421f
C80 B.n49 VSUBS 0.08526f
C81 B.n50 VSUBS 0.019943f
C82 B.n51 VSUBS 0.008608f
C83 B.n52 VSUBS 0.008608f
C84 B.n53 VSUBS 0.008608f
C85 B.n54 VSUBS 0.008608f
C86 B.n55 VSUBS 0.008608f
C87 B.t2 VSUBS 0.497292f
C88 B.t1 VSUBS 0.518609f
C89 B.t0 VSUBS 1.35737f
C90 B.n56 VSUBS 0.25243f
C91 B.n57 VSUBS 0.08527f
C92 B.n58 VSUBS 0.008608f
C93 B.n59 VSUBS 0.008608f
C94 B.n60 VSUBS 0.008608f
C95 B.n61 VSUBS 0.008608f
C96 B.n62 VSUBS 0.008608f
C97 B.n63 VSUBS 0.008608f
C98 B.n64 VSUBS 0.008608f
C99 B.n65 VSUBS 0.008608f
C100 B.n66 VSUBS 0.008608f
C101 B.n67 VSUBS 0.008608f
C102 B.n68 VSUBS 0.008608f
C103 B.n69 VSUBS 0.008608f
C104 B.n70 VSUBS 0.008608f
C105 B.n71 VSUBS 0.008608f
C106 B.n72 VSUBS 0.008608f
C107 B.n73 VSUBS 0.008608f
C108 B.n74 VSUBS 0.008608f
C109 B.n75 VSUBS 0.008608f
C110 B.n76 VSUBS 0.008608f
C111 B.n77 VSUBS 0.008608f
C112 B.n78 VSUBS 0.020699f
C113 B.n79 VSUBS 0.008608f
C114 B.n80 VSUBS 0.008608f
C115 B.n81 VSUBS 0.008608f
C116 B.n82 VSUBS 0.008608f
C117 B.n83 VSUBS 0.008608f
C118 B.n84 VSUBS 0.008608f
C119 B.n85 VSUBS 0.008608f
C120 B.n86 VSUBS 0.008608f
C121 B.n87 VSUBS 0.008608f
C122 B.n88 VSUBS 0.008608f
C123 B.n89 VSUBS 0.008608f
C124 B.n90 VSUBS 0.008608f
C125 B.n91 VSUBS 0.008608f
C126 B.n92 VSUBS 0.008608f
C127 B.n93 VSUBS 0.008608f
C128 B.n94 VSUBS 0.008608f
C129 B.n95 VSUBS 0.008608f
C130 B.n96 VSUBS 0.008608f
C131 B.n97 VSUBS 0.008608f
C132 B.n98 VSUBS 0.008608f
C133 B.n99 VSUBS 0.008608f
C134 B.n100 VSUBS 0.008608f
C135 B.n101 VSUBS 0.008608f
C136 B.n102 VSUBS 0.008608f
C137 B.n103 VSUBS 0.008608f
C138 B.n104 VSUBS 0.008608f
C139 B.n105 VSUBS 0.008608f
C140 B.n106 VSUBS 0.008608f
C141 B.n107 VSUBS 0.008608f
C142 B.n108 VSUBS 0.008608f
C143 B.n109 VSUBS 0.008608f
C144 B.n110 VSUBS 0.008608f
C145 B.n111 VSUBS 0.008608f
C146 B.n112 VSUBS 0.008608f
C147 B.n113 VSUBS 0.008608f
C148 B.n114 VSUBS 0.008608f
C149 B.n115 VSUBS 0.008608f
C150 B.n116 VSUBS 0.008608f
C151 B.n117 VSUBS 0.008608f
C152 B.n118 VSUBS 0.008608f
C153 B.n119 VSUBS 0.008608f
C154 B.n120 VSUBS 0.008608f
C155 B.n121 VSUBS 0.008608f
C156 B.n122 VSUBS 0.008608f
C157 B.n123 VSUBS 0.008608f
C158 B.n124 VSUBS 0.008608f
C159 B.n125 VSUBS 0.008608f
C160 B.n126 VSUBS 0.008608f
C161 B.n127 VSUBS 0.008608f
C162 B.n128 VSUBS 0.021653f
C163 B.n129 VSUBS 0.008608f
C164 B.n130 VSUBS 0.008608f
C165 B.n131 VSUBS 0.008608f
C166 B.n132 VSUBS 0.008608f
C167 B.n133 VSUBS 0.008608f
C168 B.n134 VSUBS 0.008608f
C169 B.n135 VSUBS 0.008608f
C170 B.n136 VSUBS 0.008608f
C171 B.n137 VSUBS 0.008608f
C172 B.n138 VSUBS 0.008608f
C173 B.n139 VSUBS 0.008608f
C174 B.n140 VSUBS 0.008608f
C175 B.n141 VSUBS 0.008608f
C176 B.n142 VSUBS 0.008608f
C177 B.n143 VSUBS 0.008608f
C178 B.n144 VSUBS 0.008608f
C179 B.n145 VSUBS 0.008608f
C180 B.n146 VSUBS 0.008608f
C181 B.n147 VSUBS 0.008608f
C182 B.n148 VSUBS 0.008608f
C183 B.n149 VSUBS 0.008608f
C184 B.t4 VSUBS 0.497292f
C185 B.t5 VSUBS 0.518609f
C186 B.t3 VSUBS 1.35737f
C187 B.n150 VSUBS 0.25243f
C188 B.n151 VSUBS 0.08527f
C189 B.n152 VSUBS 0.008608f
C190 B.n153 VSUBS 0.008608f
C191 B.n154 VSUBS 0.008608f
C192 B.n155 VSUBS 0.008608f
C193 B.t10 VSUBS 0.497302f
C194 B.t11 VSUBS 0.518618f
C195 B.t9 VSUBS 1.35737f
C196 B.n156 VSUBS 0.252421f
C197 B.n157 VSUBS 0.08526f
C198 B.n158 VSUBS 0.019943f
C199 B.n159 VSUBS 0.008608f
C200 B.n160 VSUBS 0.008608f
C201 B.n161 VSUBS 0.008608f
C202 B.n162 VSUBS 0.008608f
C203 B.n163 VSUBS 0.008608f
C204 B.n164 VSUBS 0.008608f
C205 B.n165 VSUBS 0.008608f
C206 B.n166 VSUBS 0.008608f
C207 B.n167 VSUBS 0.008608f
C208 B.n168 VSUBS 0.008608f
C209 B.n169 VSUBS 0.008608f
C210 B.n170 VSUBS 0.008608f
C211 B.n171 VSUBS 0.008608f
C212 B.n172 VSUBS 0.008608f
C213 B.n173 VSUBS 0.008608f
C214 B.n174 VSUBS 0.008608f
C215 B.n175 VSUBS 0.008608f
C216 B.n176 VSUBS 0.008608f
C217 B.n177 VSUBS 0.008608f
C218 B.n178 VSUBS 0.008608f
C219 B.n179 VSUBS 0.008608f
C220 B.n180 VSUBS 0.020373f
C221 B.n181 VSUBS 0.008608f
C222 B.n182 VSUBS 0.008608f
C223 B.n183 VSUBS 0.008608f
C224 B.n184 VSUBS 0.008608f
C225 B.n185 VSUBS 0.008608f
C226 B.n186 VSUBS 0.008608f
C227 B.n187 VSUBS 0.008608f
C228 B.n188 VSUBS 0.008608f
C229 B.n189 VSUBS 0.008608f
C230 B.n190 VSUBS 0.008608f
C231 B.n191 VSUBS 0.008608f
C232 B.n192 VSUBS 0.008608f
C233 B.n193 VSUBS 0.008608f
C234 B.n194 VSUBS 0.008608f
C235 B.n195 VSUBS 0.008608f
C236 B.n196 VSUBS 0.008608f
C237 B.n197 VSUBS 0.008608f
C238 B.n198 VSUBS 0.008608f
C239 B.n199 VSUBS 0.008608f
C240 B.n200 VSUBS 0.008608f
C241 B.n201 VSUBS 0.008608f
C242 B.n202 VSUBS 0.008608f
C243 B.n203 VSUBS 0.008608f
C244 B.n204 VSUBS 0.008608f
C245 B.n205 VSUBS 0.008608f
C246 B.n206 VSUBS 0.008608f
C247 B.n207 VSUBS 0.008608f
C248 B.n208 VSUBS 0.008608f
C249 B.n209 VSUBS 0.008608f
C250 B.n210 VSUBS 0.008608f
C251 B.n211 VSUBS 0.008608f
C252 B.n212 VSUBS 0.008608f
C253 B.n213 VSUBS 0.008608f
C254 B.n214 VSUBS 0.008608f
C255 B.n215 VSUBS 0.008608f
C256 B.n216 VSUBS 0.008608f
C257 B.n217 VSUBS 0.008608f
C258 B.n218 VSUBS 0.008608f
C259 B.n219 VSUBS 0.008608f
C260 B.n220 VSUBS 0.008608f
C261 B.n221 VSUBS 0.008608f
C262 B.n222 VSUBS 0.008608f
C263 B.n223 VSUBS 0.008608f
C264 B.n224 VSUBS 0.008608f
C265 B.n225 VSUBS 0.008608f
C266 B.n226 VSUBS 0.008608f
C267 B.n227 VSUBS 0.008608f
C268 B.n228 VSUBS 0.008608f
C269 B.n229 VSUBS 0.008608f
C270 B.n230 VSUBS 0.008608f
C271 B.n231 VSUBS 0.008608f
C272 B.n232 VSUBS 0.008608f
C273 B.n233 VSUBS 0.008608f
C274 B.n234 VSUBS 0.008608f
C275 B.n235 VSUBS 0.008608f
C276 B.n236 VSUBS 0.008608f
C277 B.n237 VSUBS 0.008608f
C278 B.n238 VSUBS 0.008608f
C279 B.n239 VSUBS 0.008608f
C280 B.n240 VSUBS 0.008608f
C281 B.n241 VSUBS 0.008608f
C282 B.n242 VSUBS 0.008608f
C283 B.n243 VSUBS 0.008608f
C284 B.n244 VSUBS 0.008608f
C285 B.n245 VSUBS 0.008608f
C286 B.n246 VSUBS 0.008608f
C287 B.n247 VSUBS 0.008608f
C288 B.n248 VSUBS 0.008608f
C289 B.n249 VSUBS 0.008608f
C290 B.n250 VSUBS 0.008608f
C291 B.n251 VSUBS 0.008608f
C292 B.n252 VSUBS 0.008608f
C293 B.n253 VSUBS 0.008608f
C294 B.n254 VSUBS 0.008608f
C295 B.n255 VSUBS 0.008608f
C296 B.n256 VSUBS 0.008608f
C297 B.n257 VSUBS 0.008608f
C298 B.n258 VSUBS 0.008608f
C299 B.n259 VSUBS 0.008608f
C300 B.n260 VSUBS 0.008608f
C301 B.n261 VSUBS 0.008608f
C302 B.n262 VSUBS 0.008608f
C303 B.n263 VSUBS 0.008608f
C304 B.n264 VSUBS 0.008608f
C305 B.n265 VSUBS 0.008608f
C306 B.n266 VSUBS 0.008608f
C307 B.n267 VSUBS 0.008608f
C308 B.n268 VSUBS 0.008608f
C309 B.n269 VSUBS 0.008608f
C310 B.n270 VSUBS 0.008608f
C311 B.n271 VSUBS 0.008608f
C312 B.n272 VSUBS 0.008608f
C313 B.n273 VSUBS 0.008608f
C314 B.n274 VSUBS 0.008608f
C315 B.n275 VSUBS 0.020373f
C316 B.n276 VSUBS 0.021653f
C317 B.n277 VSUBS 0.021653f
C318 B.n278 VSUBS 0.008608f
C319 B.n279 VSUBS 0.008608f
C320 B.n280 VSUBS 0.008608f
C321 B.n281 VSUBS 0.008608f
C322 B.n282 VSUBS 0.008608f
C323 B.n283 VSUBS 0.008608f
C324 B.n284 VSUBS 0.008608f
C325 B.n285 VSUBS 0.008608f
C326 B.n286 VSUBS 0.008608f
C327 B.n287 VSUBS 0.008608f
C328 B.n288 VSUBS 0.008608f
C329 B.n289 VSUBS 0.008608f
C330 B.n290 VSUBS 0.008608f
C331 B.n291 VSUBS 0.008608f
C332 B.n292 VSUBS 0.008608f
C333 B.n293 VSUBS 0.008608f
C334 B.n294 VSUBS 0.008608f
C335 B.n295 VSUBS 0.008608f
C336 B.n296 VSUBS 0.008608f
C337 B.n297 VSUBS 0.008608f
C338 B.n298 VSUBS 0.008608f
C339 B.n299 VSUBS 0.008608f
C340 B.n300 VSUBS 0.008608f
C341 B.n301 VSUBS 0.008608f
C342 B.n302 VSUBS 0.008608f
C343 B.n303 VSUBS 0.008608f
C344 B.n304 VSUBS 0.008608f
C345 B.n305 VSUBS 0.008608f
C346 B.n306 VSUBS 0.008608f
C347 B.n307 VSUBS 0.008608f
C348 B.n308 VSUBS 0.008608f
C349 B.n309 VSUBS 0.008608f
C350 B.n310 VSUBS 0.008608f
C351 B.n311 VSUBS 0.008608f
C352 B.n312 VSUBS 0.008608f
C353 B.n313 VSUBS 0.008608f
C354 B.n314 VSUBS 0.008608f
C355 B.n315 VSUBS 0.008608f
C356 B.n316 VSUBS 0.008608f
C357 B.n317 VSUBS 0.008608f
C358 B.n318 VSUBS 0.008608f
C359 B.n319 VSUBS 0.008608f
C360 B.n320 VSUBS 0.008608f
C361 B.n321 VSUBS 0.008608f
C362 B.n322 VSUBS 0.008608f
C363 B.n323 VSUBS 0.008608f
C364 B.n324 VSUBS 0.008608f
C365 B.n325 VSUBS 0.008608f
C366 B.n326 VSUBS 0.008608f
C367 B.n327 VSUBS 0.008608f
C368 B.n328 VSUBS 0.008608f
C369 B.n329 VSUBS 0.008608f
C370 B.n330 VSUBS 0.008608f
C371 B.n331 VSUBS 0.008608f
C372 B.n332 VSUBS 0.008608f
C373 B.n333 VSUBS 0.008608f
C374 B.n334 VSUBS 0.008608f
C375 B.n335 VSUBS 0.008608f
C376 B.n336 VSUBS 0.008608f
C377 B.n337 VSUBS 0.008608f
C378 B.n338 VSUBS 0.008608f
C379 B.n339 VSUBS 0.005949f
C380 B.n340 VSUBS 0.008608f
C381 B.n341 VSUBS 0.008608f
C382 B.n342 VSUBS 0.006962f
C383 B.n343 VSUBS 0.008608f
C384 B.n344 VSUBS 0.008608f
C385 B.n345 VSUBS 0.008608f
C386 B.n346 VSUBS 0.008608f
C387 B.n347 VSUBS 0.008608f
C388 B.n348 VSUBS 0.008608f
C389 B.n349 VSUBS 0.008608f
C390 B.n350 VSUBS 0.008608f
C391 B.n351 VSUBS 0.008608f
C392 B.n352 VSUBS 0.008608f
C393 B.n353 VSUBS 0.008608f
C394 B.n354 VSUBS 0.006962f
C395 B.n355 VSUBS 0.019943f
C396 B.n356 VSUBS 0.005949f
C397 B.n357 VSUBS 0.008608f
C398 B.n358 VSUBS 0.008608f
C399 B.n359 VSUBS 0.008608f
C400 B.n360 VSUBS 0.008608f
C401 B.n361 VSUBS 0.008608f
C402 B.n362 VSUBS 0.008608f
C403 B.n363 VSUBS 0.008608f
C404 B.n364 VSUBS 0.008608f
C405 B.n365 VSUBS 0.008608f
C406 B.n366 VSUBS 0.008608f
C407 B.n367 VSUBS 0.008608f
C408 B.n368 VSUBS 0.008608f
C409 B.n369 VSUBS 0.008608f
C410 B.n370 VSUBS 0.008608f
C411 B.n371 VSUBS 0.008608f
C412 B.n372 VSUBS 0.008608f
C413 B.n373 VSUBS 0.008608f
C414 B.n374 VSUBS 0.008608f
C415 B.n375 VSUBS 0.008608f
C416 B.n376 VSUBS 0.008608f
C417 B.n377 VSUBS 0.008608f
C418 B.n378 VSUBS 0.008608f
C419 B.n379 VSUBS 0.008608f
C420 B.n380 VSUBS 0.008608f
C421 B.n381 VSUBS 0.008608f
C422 B.n382 VSUBS 0.008608f
C423 B.n383 VSUBS 0.008608f
C424 B.n384 VSUBS 0.008608f
C425 B.n385 VSUBS 0.008608f
C426 B.n386 VSUBS 0.008608f
C427 B.n387 VSUBS 0.008608f
C428 B.n388 VSUBS 0.008608f
C429 B.n389 VSUBS 0.008608f
C430 B.n390 VSUBS 0.008608f
C431 B.n391 VSUBS 0.008608f
C432 B.n392 VSUBS 0.008608f
C433 B.n393 VSUBS 0.008608f
C434 B.n394 VSUBS 0.008608f
C435 B.n395 VSUBS 0.008608f
C436 B.n396 VSUBS 0.008608f
C437 B.n397 VSUBS 0.008608f
C438 B.n398 VSUBS 0.008608f
C439 B.n399 VSUBS 0.008608f
C440 B.n400 VSUBS 0.008608f
C441 B.n401 VSUBS 0.008608f
C442 B.n402 VSUBS 0.008608f
C443 B.n403 VSUBS 0.008608f
C444 B.n404 VSUBS 0.008608f
C445 B.n405 VSUBS 0.008608f
C446 B.n406 VSUBS 0.008608f
C447 B.n407 VSUBS 0.008608f
C448 B.n408 VSUBS 0.008608f
C449 B.n409 VSUBS 0.008608f
C450 B.n410 VSUBS 0.008608f
C451 B.n411 VSUBS 0.008608f
C452 B.n412 VSUBS 0.008608f
C453 B.n413 VSUBS 0.008608f
C454 B.n414 VSUBS 0.008608f
C455 B.n415 VSUBS 0.008608f
C456 B.n416 VSUBS 0.008608f
C457 B.n417 VSUBS 0.008608f
C458 B.n418 VSUBS 0.008608f
C459 B.n419 VSUBS 0.021653f
C460 B.n420 VSUBS 0.020373f
C461 B.n421 VSUBS 0.020373f
C462 B.n422 VSUBS 0.008608f
C463 B.n423 VSUBS 0.008608f
C464 B.n424 VSUBS 0.008608f
C465 B.n425 VSUBS 0.008608f
C466 B.n426 VSUBS 0.008608f
C467 B.n427 VSUBS 0.008608f
C468 B.n428 VSUBS 0.008608f
C469 B.n429 VSUBS 0.008608f
C470 B.n430 VSUBS 0.008608f
C471 B.n431 VSUBS 0.008608f
C472 B.n432 VSUBS 0.008608f
C473 B.n433 VSUBS 0.008608f
C474 B.n434 VSUBS 0.008608f
C475 B.n435 VSUBS 0.008608f
C476 B.n436 VSUBS 0.008608f
C477 B.n437 VSUBS 0.008608f
C478 B.n438 VSUBS 0.008608f
C479 B.n439 VSUBS 0.008608f
C480 B.n440 VSUBS 0.008608f
C481 B.n441 VSUBS 0.008608f
C482 B.n442 VSUBS 0.008608f
C483 B.n443 VSUBS 0.008608f
C484 B.n444 VSUBS 0.008608f
C485 B.n445 VSUBS 0.008608f
C486 B.n446 VSUBS 0.008608f
C487 B.n447 VSUBS 0.008608f
C488 B.n448 VSUBS 0.008608f
C489 B.n449 VSUBS 0.008608f
C490 B.n450 VSUBS 0.008608f
C491 B.n451 VSUBS 0.008608f
C492 B.n452 VSUBS 0.008608f
C493 B.n453 VSUBS 0.008608f
C494 B.n454 VSUBS 0.008608f
C495 B.n455 VSUBS 0.008608f
C496 B.n456 VSUBS 0.008608f
C497 B.n457 VSUBS 0.008608f
C498 B.n458 VSUBS 0.008608f
C499 B.n459 VSUBS 0.008608f
C500 B.n460 VSUBS 0.008608f
C501 B.n461 VSUBS 0.008608f
C502 B.n462 VSUBS 0.008608f
C503 B.n463 VSUBS 0.008608f
C504 B.n464 VSUBS 0.008608f
C505 B.n465 VSUBS 0.008608f
C506 B.n466 VSUBS 0.008608f
C507 B.n467 VSUBS 0.008608f
C508 B.n468 VSUBS 0.008608f
C509 B.n469 VSUBS 0.008608f
C510 B.n470 VSUBS 0.008608f
C511 B.n471 VSUBS 0.008608f
C512 B.n472 VSUBS 0.008608f
C513 B.n473 VSUBS 0.008608f
C514 B.n474 VSUBS 0.008608f
C515 B.n475 VSUBS 0.008608f
C516 B.n476 VSUBS 0.008608f
C517 B.n477 VSUBS 0.008608f
C518 B.n478 VSUBS 0.008608f
C519 B.n479 VSUBS 0.008608f
C520 B.n480 VSUBS 0.008608f
C521 B.n481 VSUBS 0.008608f
C522 B.n482 VSUBS 0.008608f
C523 B.n483 VSUBS 0.008608f
C524 B.n484 VSUBS 0.008608f
C525 B.n485 VSUBS 0.008608f
C526 B.n486 VSUBS 0.008608f
C527 B.n487 VSUBS 0.008608f
C528 B.n488 VSUBS 0.008608f
C529 B.n489 VSUBS 0.008608f
C530 B.n490 VSUBS 0.008608f
C531 B.n491 VSUBS 0.008608f
C532 B.n492 VSUBS 0.008608f
C533 B.n493 VSUBS 0.008608f
C534 B.n494 VSUBS 0.008608f
C535 B.n495 VSUBS 0.008608f
C536 B.n496 VSUBS 0.008608f
C537 B.n497 VSUBS 0.008608f
C538 B.n498 VSUBS 0.008608f
C539 B.n499 VSUBS 0.008608f
C540 B.n500 VSUBS 0.008608f
C541 B.n501 VSUBS 0.008608f
C542 B.n502 VSUBS 0.008608f
C543 B.n503 VSUBS 0.008608f
C544 B.n504 VSUBS 0.008608f
C545 B.n505 VSUBS 0.008608f
C546 B.n506 VSUBS 0.008608f
C547 B.n507 VSUBS 0.008608f
C548 B.n508 VSUBS 0.008608f
C549 B.n509 VSUBS 0.008608f
C550 B.n510 VSUBS 0.008608f
C551 B.n511 VSUBS 0.008608f
C552 B.n512 VSUBS 0.008608f
C553 B.n513 VSUBS 0.008608f
C554 B.n514 VSUBS 0.008608f
C555 B.n515 VSUBS 0.008608f
C556 B.n516 VSUBS 0.008608f
C557 B.n517 VSUBS 0.008608f
C558 B.n518 VSUBS 0.008608f
C559 B.n519 VSUBS 0.008608f
C560 B.n520 VSUBS 0.008608f
C561 B.n521 VSUBS 0.008608f
C562 B.n522 VSUBS 0.008608f
C563 B.n523 VSUBS 0.008608f
C564 B.n524 VSUBS 0.008608f
C565 B.n525 VSUBS 0.008608f
C566 B.n526 VSUBS 0.008608f
C567 B.n527 VSUBS 0.008608f
C568 B.n528 VSUBS 0.008608f
C569 B.n529 VSUBS 0.008608f
C570 B.n530 VSUBS 0.008608f
C571 B.n531 VSUBS 0.008608f
C572 B.n532 VSUBS 0.008608f
C573 B.n533 VSUBS 0.008608f
C574 B.n534 VSUBS 0.008608f
C575 B.n535 VSUBS 0.008608f
C576 B.n536 VSUBS 0.008608f
C577 B.n537 VSUBS 0.008608f
C578 B.n538 VSUBS 0.008608f
C579 B.n539 VSUBS 0.008608f
C580 B.n540 VSUBS 0.008608f
C581 B.n541 VSUBS 0.008608f
C582 B.n542 VSUBS 0.008608f
C583 B.n543 VSUBS 0.008608f
C584 B.n544 VSUBS 0.008608f
C585 B.n545 VSUBS 0.008608f
C586 B.n546 VSUBS 0.008608f
C587 B.n547 VSUBS 0.008608f
C588 B.n548 VSUBS 0.008608f
C589 B.n549 VSUBS 0.008608f
C590 B.n550 VSUBS 0.008608f
C591 B.n551 VSUBS 0.008608f
C592 B.n552 VSUBS 0.008608f
C593 B.n553 VSUBS 0.008608f
C594 B.n554 VSUBS 0.008608f
C595 B.n555 VSUBS 0.008608f
C596 B.n556 VSUBS 0.008608f
C597 B.n557 VSUBS 0.008608f
C598 B.n558 VSUBS 0.008608f
C599 B.n559 VSUBS 0.008608f
C600 B.n560 VSUBS 0.008608f
C601 B.n561 VSUBS 0.008608f
C602 B.n562 VSUBS 0.008608f
C603 B.n563 VSUBS 0.008608f
C604 B.n564 VSUBS 0.008608f
C605 B.n565 VSUBS 0.008608f
C606 B.n566 VSUBS 0.008608f
C607 B.n567 VSUBS 0.021327f
C608 B.n568 VSUBS 0.020373f
C609 B.n569 VSUBS 0.021653f
C610 B.n570 VSUBS 0.008608f
C611 B.n571 VSUBS 0.008608f
C612 B.n572 VSUBS 0.008608f
C613 B.n573 VSUBS 0.008608f
C614 B.n574 VSUBS 0.008608f
C615 B.n575 VSUBS 0.008608f
C616 B.n576 VSUBS 0.008608f
C617 B.n577 VSUBS 0.008608f
C618 B.n578 VSUBS 0.008608f
C619 B.n579 VSUBS 0.008608f
C620 B.n580 VSUBS 0.008608f
C621 B.n581 VSUBS 0.008608f
C622 B.n582 VSUBS 0.008608f
C623 B.n583 VSUBS 0.008608f
C624 B.n584 VSUBS 0.008608f
C625 B.n585 VSUBS 0.008608f
C626 B.n586 VSUBS 0.008608f
C627 B.n587 VSUBS 0.008608f
C628 B.n588 VSUBS 0.008608f
C629 B.n589 VSUBS 0.008608f
C630 B.n590 VSUBS 0.008608f
C631 B.n591 VSUBS 0.008608f
C632 B.n592 VSUBS 0.008608f
C633 B.n593 VSUBS 0.008608f
C634 B.n594 VSUBS 0.008608f
C635 B.n595 VSUBS 0.008608f
C636 B.n596 VSUBS 0.008608f
C637 B.n597 VSUBS 0.008608f
C638 B.n598 VSUBS 0.008608f
C639 B.n599 VSUBS 0.008608f
C640 B.n600 VSUBS 0.008608f
C641 B.n601 VSUBS 0.008608f
C642 B.n602 VSUBS 0.008608f
C643 B.n603 VSUBS 0.008608f
C644 B.n604 VSUBS 0.008608f
C645 B.n605 VSUBS 0.008608f
C646 B.n606 VSUBS 0.008608f
C647 B.n607 VSUBS 0.008608f
C648 B.n608 VSUBS 0.008608f
C649 B.n609 VSUBS 0.008608f
C650 B.n610 VSUBS 0.008608f
C651 B.n611 VSUBS 0.008608f
C652 B.n612 VSUBS 0.008608f
C653 B.n613 VSUBS 0.008608f
C654 B.n614 VSUBS 0.008608f
C655 B.n615 VSUBS 0.008608f
C656 B.n616 VSUBS 0.008608f
C657 B.n617 VSUBS 0.008608f
C658 B.n618 VSUBS 0.008608f
C659 B.n619 VSUBS 0.008608f
C660 B.n620 VSUBS 0.008608f
C661 B.n621 VSUBS 0.008608f
C662 B.n622 VSUBS 0.008608f
C663 B.n623 VSUBS 0.008608f
C664 B.n624 VSUBS 0.008608f
C665 B.n625 VSUBS 0.008608f
C666 B.n626 VSUBS 0.008608f
C667 B.n627 VSUBS 0.008608f
C668 B.n628 VSUBS 0.008608f
C669 B.n629 VSUBS 0.008608f
C670 B.n630 VSUBS 0.008608f
C671 B.n631 VSUBS 0.008608f
C672 B.n632 VSUBS 0.005949f
C673 B.n633 VSUBS 0.019943f
C674 B.n634 VSUBS 0.006962f
C675 B.n635 VSUBS 0.008608f
C676 B.n636 VSUBS 0.008608f
C677 B.n637 VSUBS 0.008608f
C678 B.n638 VSUBS 0.008608f
C679 B.n639 VSUBS 0.008608f
C680 B.n640 VSUBS 0.008608f
C681 B.n641 VSUBS 0.008608f
C682 B.n642 VSUBS 0.008608f
C683 B.n643 VSUBS 0.008608f
C684 B.n644 VSUBS 0.008608f
C685 B.n645 VSUBS 0.008608f
C686 B.n646 VSUBS 0.006962f
C687 B.n647 VSUBS 0.008608f
C688 B.n648 VSUBS 0.008608f
C689 B.n649 VSUBS 0.005949f
C690 B.n650 VSUBS 0.008608f
C691 B.n651 VSUBS 0.008608f
C692 B.n652 VSUBS 0.008608f
C693 B.n653 VSUBS 0.008608f
C694 B.n654 VSUBS 0.008608f
C695 B.n655 VSUBS 0.008608f
C696 B.n656 VSUBS 0.008608f
C697 B.n657 VSUBS 0.008608f
C698 B.n658 VSUBS 0.008608f
C699 B.n659 VSUBS 0.008608f
C700 B.n660 VSUBS 0.008608f
C701 B.n661 VSUBS 0.008608f
C702 B.n662 VSUBS 0.008608f
C703 B.n663 VSUBS 0.008608f
C704 B.n664 VSUBS 0.008608f
C705 B.n665 VSUBS 0.008608f
C706 B.n666 VSUBS 0.008608f
C707 B.n667 VSUBS 0.008608f
C708 B.n668 VSUBS 0.008608f
C709 B.n669 VSUBS 0.008608f
C710 B.n670 VSUBS 0.008608f
C711 B.n671 VSUBS 0.008608f
C712 B.n672 VSUBS 0.008608f
C713 B.n673 VSUBS 0.008608f
C714 B.n674 VSUBS 0.008608f
C715 B.n675 VSUBS 0.008608f
C716 B.n676 VSUBS 0.008608f
C717 B.n677 VSUBS 0.008608f
C718 B.n678 VSUBS 0.008608f
C719 B.n679 VSUBS 0.008608f
C720 B.n680 VSUBS 0.008608f
C721 B.n681 VSUBS 0.008608f
C722 B.n682 VSUBS 0.008608f
C723 B.n683 VSUBS 0.008608f
C724 B.n684 VSUBS 0.008608f
C725 B.n685 VSUBS 0.008608f
C726 B.n686 VSUBS 0.008608f
C727 B.n687 VSUBS 0.008608f
C728 B.n688 VSUBS 0.008608f
C729 B.n689 VSUBS 0.008608f
C730 B.n690 VSUBS 0.008608f
C731 B.n691 VSUBS 0.008608f
C732 B.n692 VSUBS 0.008608f
C733 B.n693 VSUBS 0.008608f
C734 B.n694 VSUBS 0.008608f
C735 B.n695 VSUBS 0.008608f
C736 B.n696 VSUBS 0.008608f
C737 B.n697 VSUBS 0.008608f
C738 B.n698 VSUBS 0.008608f
C739 B.n699 VSUBS 0.008608f
C740 B.n700 VSUBS 0.008608f
C741 B.n701 VSUBS 0.008608f
C742 B.n702 VSUBS 0.008608f
C743 B.n703 VSUBS 0.008608f
C744 B.n704 VSUBS 0.008608f
C745 B.n705 VSUBS 0.008608f
C746 B.n706 VSUBS 0.008608f
C747 B.n707 VSUBS 0.008608f
C748 B.n708 VSUBS 0.008608f
C749 B.n709 VSUBS 0.008608f
C750 B.n710 VSUBS 0.008608f
C751 B.n711 VSUBS 0.021653f
C752 B.n712 VSUBS 0.021653f
C753 B.n713 VSUBS 0.020373f
C754 B.n714 VSUBS 0.008608f
C755 B.n715 VSUBS 0.008608f
C756 B.n716 VSUBS 0.008608f
C757 B.n717 VSUBS 0.008608f
C758 B.n718 VSUBS 0.008608f
C759 B.n719 VSUBS 0.008608f
C760 B.n720 VSUBS 0.008608f
C761 B.n721 VSUBS 0.008608f
C762 B.n722 VSUBS 0.008608f
C763 B.n723 VSUBS 0.008608f
C764 B.n724 VSUBS 0.008608f
C765 B.n725 VSUBS 0.008608f
C766 B.n726 VSUBS 0.008608f
C767 B.n727 VSUBS 0.008608f
C768 B.n728 VSUBS 0.008608f
C769 B.n729 VSUBS 0.008608f
C770 B.n730 VSUBS 0.008608f
C771 B.n731 VSUBS 0.008608f
C772 B.n732 VSUBS 0.008608f
C773 B.n733 VSUBS 0.008608f
C774 B.n734 VSUBS 0.008608f
C775 B.n735 VSUBS 0.008608f
C776 B.n736 VSUBS 0.008608f
C777 B.n737 VSUBS 0.008608f
C778 B.n738 VSUBS 0.008608f
C779 B.n739 VSUBS 0.008608f
C780 B.n740 VSUBS 0.008608f
C781 B.n741 VSUBS 0.008608f
C782 B.n742 VSUBS 0.008608f
C783 B.n743 VSUBS 0.008608f
C784 B.n744 VSUBS 0.008608f
C785 B.n745 VSUBS 0.008608f
C786 B.n746 VSUBS 0.008608f
C787 B.n747 VSUBS 0.008608f
C788 B.n748 VSUBS 0.008608f
C789 B.n749 VSUBS 0.008608f
C790 B.n750 VSUBS 0.008608f
C791 B.n751 VSUBS 0.008608f
C792 B.n752 VSUBS 0.008608f
C793 B.n753 VSUBS 0.008608f
C794 B.n754 VSUBS 0.008608f
C795 B.n755 VSUBS 0.008608f
C796 B.n756 VSUBS 0.008608f
C797 B.n757 VSUBS 0.008608f
C798 B.n758 VSUBS 0.008608f
C799 B.n759 VSUBS 0.008608f
C800 B.n760 VSUBS 0.008608f
C801 B.n761 VSUBS 0.008608f
C802 B.n762 VSUBS 0.008608f
C803 B.n763 VSUBS 0.008608f
C804 B.n764 VSUBS 0.008608f
C805 B.n765 VSUBS 0.008608f
C806 B.n766 VSUBS 0.008608f
C807 B.n767 VSUBS 0.008608f
C808 B.n768 VSUBS 0.008608f
C809 B.n769 VSUBS 0.008608f
C810 B.n770 VSUBS 0.008608f
C811 B.n771 VSUBS 0.008608f
C812 B.n772 VSUBS 0.008608f
C813 B.n773 VSUBS 0.008608f
C814 B.n774 VSUBS 0.008608f
C815 B.n775 VSUBS 0.008608f
C816 B.n776 VSUBS 0.008608f
C817 B.n777 VSUBS 0.008608f
C818 B.n778 VSUBS 0.008608f
C819 B.n779 VSUBS 0.008608f
C820 B.n780 VSUBS 0.008608f
C821 B.n781 VSUBS 0.008608f
C822 B.n782 VSUBS 0.008608f
C823 B.n783 VSUBS 0.008608f
C824 B.n784 VSUBS 0.008608f
C825 B.n785 VSUBS 0.008608f
C826 B.n786 VSUBS 0.008608f
C827 B.n787 VSUBS 0.019491f
C828 VDD1.t8 VSUBS 2.76339f
C829 VDD1.t5 VSUBS 0.268919f
C830 VDD1.t1 VSUBS 0.268919f
C831 VDD1.n0 VSUBS 2.09973f
C832 VDD1.n1 VSUBS 1.54478f
C833 VDD1.t3 VSUBS 2.76338f
C834 VDD1.t9 VSUBS 0.268919f
C835 VDD1.t6 VSUBS 0.268919f
C836 VDD1.n2 VSUBS 2.09972f
C837 VDD1.n3 VSUBS 1.53616f
C838 VDD1.t4 VSUBS 0.268919f
C839 VDD1.t0 VSUBS 0.268919f
C840 VDD1.n4 VSUBS 2.11663f
C841 VDD1.n5 VSUBS 3.295f
C842 VDD1.t7 VSUBS 0.268919f
C843 VDD1.t2 VSUBS 0.268919f
C844 VDD1.n6 VSUBS 2.09972f
C845 VDD1.n7 VSUBS 3.55209f
C846 VP.n0 VSUBS 0.043429f
C847 VP.t9 VSUBS 2.22234f
C848 VP.n1 VSUBS 0.047632f
C849 VP.n2 VSUBS 0.032941f
C850 VP.t5 VSUBS 2.22234f
C851 VP.n3 VSUBS 0.02982f
C852 VP.n4 VSUBS 0.032941f
C853 VP.t3 VSUBS 2.22234f
C854 VP.n5 VSUBS 0.061393f
C855 VP.n6 VSUBS 0.032941f
C856 VP.t0 VSUBS 2.22234f
C857 VP.n7 VSUBS 0.791606f
C858 VP.n8 VSUBS 0.032941f
C859 VP.n9 VSUBS 0.055937f
C860 VP.n10 VSUBS 0.043429f
C861 VP.t7 VSUBS 2.22234f
C862 VP.n11 VSUBS 0.047632f
C863 VP.n12 VSUBS 0.032941f
C864 VP.t2 VSUBS 2.22234f
C865 VP.n13 VSUBS 0.02982f
C866 VP.n14 VSUBS 0.032941f
C867 VP.t8 VSUBS 2.22234f
C868 VP.n15 VSUBS 0.061393f
C869 VP.n16 VSUBS 0.032941f
C870 VP.t4 VSUBS 2.22234f
C871 VP.n17 VSUBS 0.860821f
C872 VP.t1 VSUBS 2.38361f
C873 VP.n18 VSUBS 0.877584f
C874 VP.n19 VSUBS 0.246614f
C875 VP.n20 VSUBS 0.035933f
C876 VP.n21 VSUBS 0.066361f
C877 VP.n22 VSUBS 0.02982f
C878 VP.n23 VSUBS 0.032941f
C879 VP.n24 VSUBS 0.032941f
C880 VP.n25 VSUBS 0.032941f
C881 VP.n26 VSUBS 0.046238f
C882 VP.n27 VSUBS 0.791606f
C883 VP.n28 VSUBS 0.046238f
C884 VP.n29 VSUBS 0.061393f
C885 VP.n30 VSUBS 0.032941f
C886 VP.n31 VSUBS 0.032941f
C887 VP.n32 VSUBS 0.032941f
C888 VP.n33 VSUBS 0.066361f
C889 VP.n34 VSUBS 0.035933f
C890 VP.n35 VSUBS 0.791606f
C891 VP.n36 VSUBS 0.056544f
C892 VP.n37 VSUBS 0.032941f
C893 VP.n38 VSUBS 0.032941f
C894 VP.n39 VSUBS 0.032941f
C895 VP.n40 VSUBS 0.04855f
C896 VP.n41 VSUBS 0.055937f
C897 VP.n42 VSUBS 0.893115f
C898 VP.n43 VSUBS 1.82699f
C899 VP.t6 VSUBS 2.22234f
C900 VP.n44 VSUBS 0.893115f
C901 VP.n45 VSUBS 1.8506f
C902 VP.n46 VSUBS 0.043429f
C903 VP.n47 VSUBS 0.032941f
C904 VP.n48 VSUBS 0.04855f
C905 VP.n49 VSUBS 0.047632f
C906 VP.n50 VSUBS 0.056544f
C907 VP.n51 VSUBS 0.032941f
C908 VP.n52 VSUBS 0.032941f
C909 VP.n53 VSUBS 0.035933f
C910 VP.n54 VSUBS 0.066361f
C911 VP.n55 VSUBS 0.02982f
C912 VP.n56 VSUBS 0.032941f
C913 VP.n57 VSUBS 0.032941f
C914 VP.n58 VSUBS 0.032941f
C915 VP.n59 VSUBS 0.046238f
C916 VP.n60 VSUBS 0.791606f
C917 VP.n61 VSUBS 0.046238f
C918 VP.n62 VSUBS 0.061393f
C919 VP.n63 VSUBS 0.032941f
C920 VP.n64 VSUBS 0.032941f
C921 VP.n65 VSUBS 0.032941f
C922 VP.n66 VSUBS 0.066361f
C923 VP.n67 VSUBS 0.035933f
C924 VP.n68 VSUBS 0.791606f
C925 VP.n69 VSUBS 0.056544f
C926 VP.n70 VSUBS 0.032941f
C927 VP.n71 VSUBS 0.032941f
C928 VP.n72 VSUBS 0.032941f
C929 VP.n73 VSUBS 0.04855f
C930 VP.n74 VSUBS 0.055937f
C931 VP.n75 VSUBS 0.893115f
C932 VP.n76 VSUBS 0.039725f
C933 VTAIL.t10 VSUBS 0.276479f
C934 VTAIL.t13 VSUBS 0.276479f
C935 VTAIL.n0 VSUBS 1.99423f
C936 VTAIL.n1 VSUBS 0.946988f
C937 VTAIL.t7 VSUBS 2.63476f
C938 VTAIL.n2 VSUBS 1.10095f
C939 VTAIL.t2 VSUBS 0.276479f
C940 VTAIL.t3 VSUBS 0.276479f
C941 VTAIL.n3 VSUBS 1.99423f
C942 VTAIL.n4 VSUBS 1.03616f
C943 VTAIL.t0 VSUBS 0.276479f
C944 VTAIL.t19 VSUBS 0.276479f
C945 VTAIL.n5 VSUBS 1.99423f
C946 VTAIL.n6 VSUBS 2.57529f
C947 VTAIL.t17 VSUBS 0.276479f
C948 VTAIL.t9 VSUBS 0.276479f
C949 VTAIL.n7 VSUBS 1.99423f
C950 VTAIL.n8 VSUBS 2.57528f
C951 VTAIL.t15 VSUBS 0.276479f
C952 VTAIL.t18 VSUBS 0.276479f
C953 VTAIL.n9 VSUBS 1.99423f
C954 VTAIL.n10 VSUBS 1.03615f
C955 VTAIL.t16 VSUBS 2.63477f
C956 VTAIL.n11 VSUBS 1.10093f
C957 VTAIL.t1 VSUBS 0.276479f
C958 VTAIL.t5 VSUBS 0.276479f
C959 VTAIL.n12 VSUBS 1.99423f
C960 VTAIL.n13 VSUBS 0.98744f
C961 VTAIL.t6 VSUBS 0.276479f
C962 VTAIL.t8 VSUBS 0.276479f
C963 VTAIL.n14 VSUBS 1.99423f
C964 VTAIL.n15 VSUBS 1.03615f
C965 VTAIL.t4 VSUBS 2.63476f
C966 VTAIL.n16 VSUBS 2.50573f
C967 VTAIL.t11 VSUBS 2.63476f
C968 VTAIL.n17 VSUBS 2.50573f
C969 VTAIL.t12 VSUBS 0.276479f
C970 VTAIL.t14 VSUBS 0.276479f
C971 VTAIL.n18 VSUBS 1.99423f
C972 VTAIL.n19 VSUBS 0.893563f
C973 VDD2.t3 VSUBS 2.76355f
C974 VDD2.t0 VSUBS 0.268936f
C975 VDD2.t1 VSUBS 0.268936f
C976 VDD2.n0 VSUBS 2.09985f
C977 VDD2.n1 VSUBS 1.53625f
C978 VDD2.t6 VSUBS 0.268936f
C979 VDD2.t9 VSUBS 0.268936f
C980 VDD2.n2 VSUBS 2.11676f
C981 VDD2.n3 VSUBS 3.17477f
C982 VDD2.t2 VSUBS 2.74215f
C983 VDD2.n4 VSUBS 3.53389f
C984 VDD2.t7 VSUBS 0.268936f
C985 VDD2.t5 VSUBS 0.268936f
C986 VDD2.n5 VSUBS 2.09986f
C987 VDD2.n6 VSUBS 0.756854f
C988 VDD2.t4 VSUBS 0.268936f
C989 VDD2.t8 VSUBS 0.268936f
C990 VDD2.n7 VSUBS 2.11671f
C991 VN.n0 VSUBS 0.042332f
C992 VN.t7 VSUBS 2.16618f
C993 VN.n1 VSUBS 0.046428f
C994 VN.n2 VSUBS 0.032108f
C995 VN.t4 VSUBS 2.16618f
C996 VN.n3 VSUBS 0.029067f
C997 VN.n4 VSUBS 0.032108f
C998 VN.t6 VSUBS 2.16618f
C999 VN.n5 VSUBS 0.059842f
C1000 VN.n6 VSUBS 0.032108f
C1001 VN.t5 VSUBS 2.16618f
C1002 VN.n7 VSUBS 0.839067f
C1003 VN.t8 VSUBS 2.32338f
C1004 VN.n8 VSUBS 0.855407f
C1005 VN.n9 VSUBS 0.240382f
C1006 VN.n10 VSUBS 0.035025f
C1007 VN.n11 VSUBS 0.064684f
C1008 VN.n12 VSUBS 0.029067f
C1009 VN.n13 VSUBS 0.032108f
C1010 VN.n14 VSUBS 0.032108f
C1011 VN.n15 VSUBS 0.032108f
C1012 VN.n16 VSUBS 0.04507f
C1013 VN.n17 VSUBS 0.771601f
C1014 VN.n18 VSUBS 0.04507f
C1015 VN.n19 VSUBS 0.059842f
C1016 VN.n20 VSUBS 0.032108f
C1017 VN.n21 VSUBS 0.032108f
C1018 VN.n22 VSUBS 0.032108f
C1019 VN.n23 VSUBS 0.064684f
C1020 VN.n24 VSUBS 0.035025f
C1021 VN.n25 VSUBS 0.771601f
C1022 VN.n26 VSUBS 0.055115f
C1023 VN.n27 VSUBS 0.032108f
C1024 VN.n28 VSUBS 0.032108f
C1025 VN.n29 VSUBS 0.032108f
C1026 VN.n30 VSUBS 0.047323f
C1027 VN.n31 VSUBS 0.054524f
C1028 VN.n32 VSUBS 0.870545f
C1029 VN.n33 VSUBS 0.038721f
C1030 VN.n34 VSUBS 0.042332f
C1031 VN.t1 VSUBS 2.16618f
C1032 VN.n35 VSUBS 0.046428f
C1033 VN.n36 VSUBS 0.032108f
C1034 VN.t9 VSUBS 2.16618f
C1035 VN.n37 VSUBS 0.029067f
C1036 VN.n38 VSUBS 0.032108f
C1037 VN.t3 VSUBS 2.16618f
C1038 VN.n39 VSUBS 0.059842f
C1039 VN.n40 VSUBS 0.032108f
C1040 VN.t0 VSUBS 2.16618f
C1041 VN.n41 VSUBS 0.839067f
C1042 VN.t2 VSUBS 2.32338f
C1043 VN.n42 VSUBS 0.855407f
C1044 VN.n43 VSUBS 0.240382f
C1045 VN.n44 VSUBS 0.035025f
C1046 VN.n45 VSUBS 0.064684f
C1047 VN.n46 VSUBS 0.029067f
C1048 VN.n47 VSUBS 0.032108f
C1049 VN.n48 VSUBS 0.032108f
C1050 VN.n49 VSUBS 0.032108f
C1051 VN.n50 VSUBS 0.04507f
C1052 VN.n51 VSUBS 0.771601f
C1053 VN.n52 VSUBS 0.04507f
C1054 VN.n53 VSUBS 0.059842f
C1055 VN.n54 VSUBS 0.032108f
C1056 VN.n55 VSUBS 0.032108f
C1057 VN.n56 VSUBS 0.032108f
C1058 VN.n57 VSUBS 0.064684f
C1059 VN.n58 VSUBS 0.035025f
C1060 VN.n59 VSUBS 0.771601f
C1061 VN.n60 VSUBS 0.055115f
C1062 VN.n61 VSUBS 0.032108f
C1063 VN.n62 VSUBS 0.032108f
C1064 VN.n63 VSUBS 0.032108f
C1065 VN.n64 VSUBS 0.047323f
C1066 VN.n65 VSUBS 0.054524f
C1067 VN.n66 VSUBS 0.870545f
C1068 VN.n67 VSUBS 1.79807f
.ends

