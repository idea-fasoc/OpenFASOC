* NGSPICE file created from diff_pair_sample_0170.ext - technology: sky130A

.subckt diff_pair_sample_0170 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0 ps=0 w=4.07 l=3.49
X1 VDD1.t5 VP.t0 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0.67155 ps=4.4 w=4.07 l=3.49
X2 VDD2.t5 VN.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0.67155 ps=4.4 w=4.07 l=3.49
X3 VTAIL.t3 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=0.67155 ps=4.4 w=4.07 l=3.49
X4 VDD1.t4 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=1.5873 ps=8.92 w=4.07 l=3.49
X5 VDD1.t3 VP.t2 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0.67155 ps=4.4 w=4.07 l=3.49
X6 VTAIL.t7 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=0.67155 ps=4.4 w=4.07 l=3.49
X7 VDD2.t3 VN.t2 VTAIL.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0.67155 ps=4.4 w=4.07 l=3.49
X8 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0 ps=0 w=4.07 l=3.49
X9 VDD2.t2 VN.t3 VTAIL.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=1.5873 ps=8.92 w=4.07 l=3.49
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0 ps=0 w=4.07 l=3.49
X11 VDD2.t1 VN.t4 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=1.5873 ps=8.92 w=4.07 l=3.49
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5873 pd=8.92 as=0 ps=0 w=4.07 l=3.49
X13 VDD1.t1 VP.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=1.5873 ps=8.92 w=4.07 l=3.49
X14 VTAIL.t9 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=0.67155 ps=4.4 w=4.07 l=3.49
X15 VTAIL.t5 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.67155 pd=4.4 as=0.67155 ps=4.4 w=4.07 l=3.49
R0 B.n667 B.n666 585
R1 B.n215 B.n120 585
R2 B.n214 B.n213 585
R3 B.n212 B.n211 585
R4 B.n210 B.n209 585
R5 B.n208 B.n207 585
R6 B.n206 B.n205 585
R7 B.n204 B.n203 585
R8 B.n202 B.n201 585
R9 B.n200 B.n199 585
R10 B.n198 B.n197 585
R11 B.n196 B.n195 585
R12 B.n194 B.n193 585
R13 B.n192 B.n191 585
R14 B.n190 B.n189 585
R15 B.n188 B.n187 585
R16 B.n186 B.n185 585
R17 B.n184 B.n183 585
R18 B.n182 B.n181 585
R19 B.n180 B.n179 585
R20 B.n178 B.n177 585
R21 B.n176 B.n175 585
R22 B.n174 B.n173 585
R23 B.n172 B.n171 585
R24 B.n170 B.n169 585
R25 B.n168 B.n167 585
R26 B.n166 B.n165 585
R27 B.n164 B.n163 585
R28 B.n162 B.n161 585
R29 B.n160 B.n159 585
R30 B.n158 B.n157 585
R31 B.n156 B.n155 585
R32 B.n154 B.n153 585
R33 B.n152 B.n151 585
R34 B.n150 B.n149 585
R35 B.n148 B.n147 585
R36 B.n146 B.n145 585
R37 B.n144 B.n143 585
R38 B.n142 B.n141 585
R39 B.n140 B.n139 585
R40 B.n138 B.n137 585
R41 B.n136 B.n135 585
R42 B.n134 B.n133 585
R43 B.n132 B.n131 585
R44 B.n130 B.n129 585
R45 B.n128 B.n127 585
R46 B.n665 B.n97 585
R47 B.n670 B.n97 585
R48 B.n664 B.n96 585
R49 B.n671 B.n96 585
R50 B.n663 B.n662 585
R51 B.n662 B.n92 585
R52 B.n661 B.n91 585
R53 B.n677 B.n91 585
R54 B.n660 B.n90 585
R55 B.n678 B.n90 585
R56 B.n659 B.n89 585
R57 B.n679 B.n89 585
R58 B.n658 B.n657 585
R59 B.n657 B.n85 585
R60 B.n656 B.n84 585
R61 B.n685 B.n84 585
R62 B.n655 B.n83 585
R63 B.n686 B.n83 585
R64 B.n654 B.n82 585
R65 B.n687 B.n82 585
R66 B.n653 B.n652 585
R67 B.n652 B.n78 585
R68 B.n651 B.n77 585
R69 B.n693 B.n77 585
R70 B.n650 B.n76 585
R71 B.n694 B.n76 585
R72 B.n649 B.n75 585
R73 B.n695 B.n75 585
R74 B.n648 B.n647 585
R75 B.n647 B.n71 585
R76 B.n646 B.n70 585
R77 B.n701 B.n70 585
R78 B.n645 B.n69 585
R79 B.n702 B.n69 585
R80 B.n644 B.n68 585
R81 B.n703 B.n68 585
R82 B.n643 B.n642 585
R83 B.n642 B.n64 585
R84 B.n641 B.n63 585
R85 B.n709 B.n63 585
R86 B.n640 B.n62 585
R87 B.n710 B.n62 585
R88 B.n639 B.n61 585
R89 B.n711 B.n61 585
R90 B.n638 B.n637 585
R91 B.n637 B.n57 585
R92 B.n636 B.n56 585
R93 B.n717 B.n56 585
R94 B.n635 B.n55 585
R95 B.n718 B.n55 585
R96 B.n634 B.n54 585
R97 B.n719 B.n54 585
R98 B.n633 B.n632 585
R99 B.n632 B.n50 585
R100 B.n631 B.n49 585
R101 B.n725 B.n49 585
R102 B.n630 B.n48 585
R103 B.n726 B.n48 585
R104 B.n629 B.n47 585
R105 B.n727 B.n47 585
R106 B.n628 B.n627 585
R107 B.n627 B.n43 585
R108 B.n626 B.n42 585
R109 B.n733 B.n42 585
R110 B.n625 B.n41 585
R111 B.n734 B.n41 585
R112 B.n624 B.n40 585
R113 B.n735 B.n40 585
R114 B.n623 B.n622 585
R115 B.n622 B.n39 585
R116 B.n621 B.n35 585
R117 B.n741 B.n35 585
R118 B.n620 B.n34 585
R119 B.n742 B.n34 585
R120 B.n619 B.n33 585
R121 B.n743 B.n33 585
R122 B.n618 B.n617 585
R123 B.n617 B.n29 585
R124 B.n616 B.n28 585
R125 B.n749 B.n28 585
R126 B.n615 B.n27 585
R127 B.n750 B.n27 585
R128 B.n614 B.n26 585
R129 B.n751 B.n26 585
R130 B.n613 B.n612 585
R131 B.n612 B.n22 585
R132 B.n611 B.n21 585
R133 B.n757 B.n21 585
R134 B.n610 B.n20 585
R135 B.n758 B.n20 585
R136 B.n609 B.n19 585
R137 B.n759 B.n19 585
R138 B.n608 B.n607 585
R139 B.n607 B.n15 585
R140 B.n606 B.n14 585
R141 B.n765 B.n14 585
R142 B.n605 B.n13 585
R143 B.n766 B.n13 585
R144 B.n604 B.n12 585
R145 B.n767 B.n12 585
R146 B.n603 B.n602 585
R147 B.n602 B.n8 585
R148 B.n601 B.n7 585
R149 B.n773 B.n7 585
R150 B.n600 B.n6 585
R151 B.n774 B.n6 585
R152 B.n599 B.n5 585
R153 B.n775 B.n5 585
R154 B.n598 B.n597 585
R155 B.n597 B.n4 585
R156 B.n596 B.n216 585
R157 B.n596 B.n595 585
R158 B.n586 B.n217 585
R159 B.n218 B.n217 585
R160 B.n588 B.n587 585
R161 B.n589 B.n588 585
R162 B.n585 B.n223 585
R163 B.n223 B.n222 585
R164 B.n584 B.n583 585
R165 B.n583 B.n582 585
R166 B.n225 B.n224 585
R167 B.n226 B.n225 585
R168 B.n575 B.n574 585
R169 B.n576 B.n575 585
R170 B.n573 B.n231 585
R171 B.n231 B.n230 585
R172 B.n572 B.n571 585
R173 B.n571 B.n570 585
R174 B.n233 B.n232 585
R175 B.n234 B.n233 585
R176 B.n563 B.n562 585
R177 B.n564 B.n563 585
R178 B.n561 B.n239 585
R179 B.n239 B.n238 585
R180 B.n560 B.n559 585
R181 B.n559 B.n558 585
R182 B.n241 B.n240 585
R183 B.n242 B.n241 585
R184 B.n551 B.n550 585
R185 B.n552 B.n551 585
R186 B.n549 B.n247 585
R187 B.n247 B.n246 585
R188 B.n548 B.n547 585
R189 B.n547 B.n546 585
R190 B.n249 B.n248 585
R191 B.n539 B.n249 585
R192 B.n538 B.n537 585
R193 B.n540 B.n538 585
R194 B.n536 B.n254 585
R195 B.n254 B.n253 585
R196 B.n535 B.n534 585
R197 B.n534 B.n533 585
R198 B.n256 B.n255 585
R199 B.n257 B.n256 585
R200 B.n526 B.n525 585
R201 B.n527 B.n526 585
R202 B.n524 B.n262 585
R203 B.n262 B.n261 585
R204 B.n523 B.n522 585
R205 B.n522 B.n521 585
R206 B.n264 B.n263 585
R207 B.n265 B.n264 585
R208 B.n514 B.n513 585
R209 B.n515 B.n514 585
R210 B.n512 B.n270 585
R211 B.n270 B.n269 585
R212 B.n511 B.n510 585
R213 B.n510 B.n509 585
R214 B.n272 B.n271 585
R215 B.n273 B.n272 585
R216 B.n502 B.n501 585
R217 B.n503 B.n502 585
R218 B.n500 B.n278 585
R219 B.n278 B.n277 585
R220 B.n499 B.n498 585
R221 B.n498 B.n497 585
R222 B.n280 B.n279 585
R223 B.n281 B.n280 585
R224 B.n490 B.n489 585
R225 B.n491 B.n490 585
R226 B.n488 B.n286 585
R227 B.n286 B.n285 585
R228 B.n487 B.n486 585
R229 B.n486 B.n485 585
R230 B.n288 B.n287 585
R231 B.n289 B.n288 585
R232 B.n478 B.n477 585
R233 B.n479 B.n478 585
R234 B.n476 B.n294 585
R235 B.n294 B.n293 585
R236 B.n475 B.n474 585
R237 B.n474 B.n473 585
R238 B.n296 B.n295 585
R239 B.n297 B.n296 585
R240 B.n466 B.n465 585
R241 B.n467 B.n466 585
R242 B.n464 B.n301 585
R243 B.n305 B.n301 585
R244 B.n463 B.n462 585
R245 B.n462 B.n461 585
R246 B.n303 B.n302 585
R247 B.n304 B.n303 585
R248 B.n454 B.n453 585
R249 B.n455 B.n454 585
R250 B.n452 B.n310 585
R251 B.n310 B.n309 585
R252 B.n451 B.n450 585
R253 B.n450 B.n449 585
R254 B.n312 B.n311 585
R255 B.n313 B.n312 585
R256 B.n442 B.n441 585
R257 B.n443 B.n442 585
R258 B.n440 B.n318 585
R259 B.n318 B.n317 585
R260 B.n435 B.n434 585
R261 B.n433 B.n343 585
R262 B.n432 B.n342 585
R263 B.n437 B.n342 585
R264 B.n431 B.n430 585
R265 B.n429 B.n428 585
R266 B.n427 B.n426 585
R267 B.n425 B.n424 585
R268 B.n423 B.n422 585
R269 B.n421 B.n420 585
R270 B.n419 B.n418 585
R271 B.n417 B.n416 585
R272 B.n415 B.n414 585
R273 B.n413 B.n412 585
R274 B.n411 B.n410 585
R275 B.n409 B.n408 585
R276 B.n407 B.n406 585
R277 B.n405 B.n404 585
R278 B.n403 B.n402 585
R279 B.n400 B.n399 585
R280 B.n398 B.n397 585
R281 B.n396 B.n395 585
R282 B.n394 B.n393 585
R283 B.n392 B.n391 585
R284 B.n390 B.n389 585
R285 B.n388 B.n387 585
R286 B.n386 B.n385 585
R287 B.n384 B.n383 585
R288 B.n382 B.n381 585
R289 B.n379 B.n378 585
R290 B.n377 B.n376 585
R291 B.n375 B.n374 585
R292 B.n373 B.n372 585
R293 B.n371 B.n370 585
R294 B.n369 B.n368 585
R295 B.n367 B.n366 585
R296 B.n365 B.n364 585
R297 B.n363 B.n362 585
R298 B.n361 B.n360 585
R299 B.n359 B.n358 585
R300 B.n357 B.n356 585
R301 B.n355 B.n354 585
R302 B.n353 B.n352 585
R303 B.n351 B.n350 585
R304 B.n349 B.n348 585
R305 B.n320 B.n319 585
R306 B.n439 B.n438 585
R307 B.n438 B.n437 585
R308 B.n316 B.n315 585
R309 B.n317 B.n316 585
R310 B.n445 B.n444 585
R311 B.n444 B.n443 585
R312 B.n446 B.n314 585
R313 B.n314 B.n313 585
R314 B.n448 B.n447 585
R315 B.n449 B.n448 585
R316 B.n308 B.n307 585
R317 B.n309 B.n308 585
R318 B.n457 B.n456 585
R319 B.n456 B.n455 585
R320 B.n458 B.n306 585
R321 B.n306 B.n304 585
R322 B.n460 B.n459 585
R323 B.n461 B.n460 585
R324 B.n300 B.n299 585
R325 B.n305 B.n300 585
R326 B.n469 B.n468 585
R327 B.n468 B.n467 585
R328 B.n470 B.n298 585
R329 B.n298 B.n297 585
R330 B.n472 B.n471 585
R331 B.n473 B.n472 585
R332 B.n292 B.n291 585
R333 B.n293 B.n292 585
R334 B.n481 B.n480 585
R335 B.n480 B.n479 585
R336 B.n482 B.n290 585
R337 B.n290 B.n289 585
R338 B.n484 B.n483 585
R339 B.n485 B.n484 585
R340 B.n284 B.n283 585
R341 B.n285 B.n284 585
R342 B.n493 B.n492 585
R343 B.n492 B.n491 585
R344 B.n494 B.n282 585
R345 B.n282 B.n281 585
R346 B.n496 B.n495 585
R347 B.n497 B.n496 585
R348 B.n276 B.n275 585
R349 B.n277 B.n276 585
R350 B.n505 B.n504 585
R351 B.n504 B.n503 585
R352 B.n506 B.n274 585
R353 B.n274 B.n273 585
R354 B.n508 B.n507 585
R355 B.n509 B.n508 585
R356 B.n268 B.n267 585
R357 B.n269 B.n268 585
R358 B.n517 B.n516 585
R359 B.n516 B.n515 585
R360 B.n518 B.n266 585
R361 B.n266 B.n265 585
R362 B.n520 B.n519 585
R363 B.n521 B.n520 585
R364 B.n260 B.n259 585
R365 B.n261 B.n260 585
R366 B.n529 B.n528 585
R367 B.n528 B.n527 585
R368 B.n530 B.n258 585
R369 B.n258 B.n257 585
R370 B.n532 B.n531 585
R371 B.n533 B.n532 585
R372 B.n252 B.n251 585
R373 B.n253 B.n252 585
R374 B.n542 B.n541 585
R375 B.n541 B.n540 585
R376 B.n543 B.n250 585
R377 B.n539 B.n250 585
R378 B.n545 B.n544 585
R379 B.n546 B.n545 585
R380 B.n245 B.n244 585
R381 B.n246 B.n245 585
R382 B.n554 B.n553 585
R383 B.n553 B.n552 585
R384 B.n555 B.n243 585
R385 B.n243 B.n242 585
R386 B.n557 B.n556 585
R387 B.n558 B.n557 585
R388 B.n237 B.n236 585
R389 B.n238 B.n237 585
R390 B.n566 B.n565 585
R391 B.n565 B.n564 585
R392 B.n567 B.n235 585
R393 B.n235 B.n234 585
R394 B.n569 B.n568 585
R395 B.n570 B.n569 585
R396 B.n229 B.n228 585
R397 B.n230 B.n229 585
R398 B.n578 B.n577 585
R399 B.n577 B.n576 585
R400 B.n579 B.n227 585
R401 B.n227 B.n226 585
R402 B.n581 B.n580 585
R403 B.n582 B.n581 585
R404 B.n221 B.n220 585
R405 B.n222 B.n221 585
R406 B.n591 B.n590 585
R407 B.n590 B.n589 585
R408 B.n592 B.n219 585
R409 B.n219 B.n218 585
R410 B.n594 B.n593 585
R411 B.n595 B.n594 585
R412 B.n2 B.n0 585
R413 B.n4 B.n2 585
R414 B.n3 B.n1 585
R415 B.n774 B.n3 585
R416 B.n772 B.n771 585
R417 B.n773 B.n772 585
R418 B.n770 B.n9 585
R419 B.n9 B.n8 585
R420 B.n769 B.n768 585
R421 B.n768 B.n767 585
R422 B.n11 B.n10 585
R423 B.n766 B.n11 585
R424 B.n764 B.n763 585
R425 B.n765 B.n764 585
R426 B.n762 B.n16 585
R427 B.n16 B.n15 585
R428 B.n761 B.n760 585
R429 B.n760 B.n759 585
R430 B.n18 B.n17 585
R431 B.n758 B.n18 585
R432 B.n756 B.n755 585
R433 B.n757 B.n756 585
R434 B.n754 B.n23 585
R435 B.n23 B.n22 585
R436 B.n753 B.n752 585
R437 B.n752 B.n751 585
R438 B.n25 B.n24 585
R439 B.n750 B.n25 585
R440 B.n748 B.n747 585
R441 B.n749 B.n748 585
R442 B.n746 B.n30 585
R443 B.n30 B.n29 585
R444 B.n745 B.n744 585
R445 B.n744 B.n743 585
R446 B.n32 B.n31 585
R447 B.n742 B.n32 585
R448 B.n740 B.n739 585
R449 B.n741 B.n740 585
R450 B.n738 B.n36 585
R451 B.n39 B.n36 585
R452 B.n737 B.n736 585
R453 B.n736 B.n735 585
R454 B.n38 B.n37 585
R455 B.n734 B.n38 585
R456 B.n732 B.n731 585
R457 B.n733 B.n732 585
R458 B.n730 B.n44 585
R459 B.n44 B.n43 585
R460 B.n729 B.n728 585
R461 B.n728 B.n727 585
R462 B.n46 B.n45 585
R463 B.n726 B.n46 585
R464 B.n724 B.n723 585
R465 B.n725 B.n724 585
R466 B.n722 B.n51 585
R467 B.n51 B.n50 585
R468 B.n721 B.n720 585
R469 B.n720 B.n719 585
R470 B.n53 B.n52 585
R471 B.n718 B.n53 585
R472 B.n716 B.n715 585
R473 B.n717 B.n716 585
R474 B.n714 B.n58 585
R475 B.n58 B.n57 585
R476 B.n713 B.n712 585
R477 B.n712 B.n711 585
R478 B.n60 B.n59 585
R479 B.n710 B.n60 585
R480 B.n708 B.n707 585
R481 B.n709 B.n708 585
R482 B.n706 B.n65 585
R483 B.n65 B.n64 585
R484 B.n705 B.n704 585
R485 B.n704 B.n703 585
R486 B.n67 B.n66 585
R487 B.n702 B.n67 585
R488 B.n700 B.n699 585
R489 B.n701 B.n700 585
R490 B.n698 B.n72 585
R491 B.n72 B.n71 585
R492 B.n697 B.n696 585
R493 B.n696 B.n695 585
R494 B.n74 B.n73 585
R495 B.n694 B.n74 585
R496 B.n692 B.n691 585
R497 B.n693 B.n692 585
R498 B.n690 B.n79 585
R499 B.n79 B.n78 585
R500 B.n689 B.n688 585
R501 B.n688 B.n687 585
R502 B.n81 B.n80 585
R503 B.n686 B.n81 585
R504 B.n684 B.n683 585
R505 B.n685 B.n684 585
R506 B.n682 B.n86 585
R507 B.n86 B.n85 585
R508 B.n681 B.n680 585
R509 B.n680 B.n679 585
R510 B.n88 B.n87 585
R511 B.n678 B.n88 585
R512 B.n676 B.n675 585
R513 B.n677 B.n676 585
R514 B.n674 B.n93 585
R515 B.n93 B.n92 585
R516 B.n673 B.n672 585
R517 B.n672 B.n671 585
R518 B.n95 B.n94 585
R519 B.n670 B.n95 585
R520 B.n777 B.n776 585
R521 B.n776 B.n775 585
R522 B.n435 B.n316 521.33
R523 B.n127 B.n95 521.33
R524 B.n438 B.n318 521.33
R525 B.n667 B.n97 521.33
R526 B.n669 B.n668 256.663
R527 B.n669 B.n119 256.663
R528 B.n669 B.n118 256.663
R529 B.n669 B.n117 256.663
R530 B.n669 B.n116 256.663
R531 B.n669 B.n115 256.663
R532 B.n669 B.n114 256.663
R533 B.n669 B.n113 256.663
R534 B.n669 B.n112 256.663
R535 B.n669 B.n111 256.663
R536 B.n669 B.n110 256.663
R537 B.n669 B.n109 256.663
R538 B.n669 B.n108 256.663
R539 B.n669 B.n107 256.663
R540 B.n669 B.n106 256.663
R541 B.n669 B.n105 256.663
R542 B.n669 B.n104 256.663
R543 B.n669 B.n103 256.663
R544 B.n669 B.n102 256.663
R545 B.n669 B.n101 256.663
R546 B.n669 B.n100 256.663
R547 B.n669 B.n99 256.663
R548 B.n669 B.n98 256.663
R549 B.n437 B.n436 256.663
R550 B.n437 B.n321 256.663
R551 B.n437 B.n322 256.663
R552 B.n437 B.n323 256.663
R553 B.n437 B.n324 256.663
R554 B.n437 B.n325 256.663
R555 B.n437 B.n326 256.663
R556 B.n437 B.n327 256.663
R557 B.n437 B.n328 256.663
R558 B.n437 B.n329 256.663
R559 B.n437 B.n330 256.663
R560 B.n437 B.n331 256.663
R561 B.n437 B.n332 256.663
R562 B.n437 B.n333 256.663
R563 B.n437 B.n334 256.663
R564 B.n437 B.n335 256.663
R565 B.n437 B.n336 256.663
R566 B.n437 B.n337 256.663
R567 B.n437 B.n338 256.663
R568 B.n437 B.n339 256.663
R569 B.n437 B.n340 256.663
R570 B.n437 B.n341 256.663
R571 B.n346 B.t17 237.19
R572 B.n344 B.t10 237.19
R573 B.n124 B.t6 237.19
R574 B.n121 B.t14 237.19
R575 B.n346 B.t19 220.702
R576 B.n121 B.t15 220.702
R577 B.n344 B.t13 220.702
R578 B.n124 B.t8 220.702
R579 B.n444 B.n316 163.367
R580 B.n444 B.n314 163.367
R581 B.n448 B.n314 163.367
R582 B.n448 B.n308 163.367
R583 B.n456 B.n308 163.367
R584 B.n456 B.n306 163.367
R585 B.n460 B.n306 163.367
R586 B.n460 B.n300 163.367
R587 B.n468 B.n300 163.367
R588 B.n468 B.n298 163.367
R589 B.n472 B.n298 163.367
R590 B.n472 B.n292 163.367
R591 B.n480 B.n292 163.367
R592 B.n480 B.n290 163.367
R593 B.n484 B.n290 163.367
R594 B.n484 B.n284 163.367
R595 B.n492 B.n284 163.367
R596 B.n492 B.n282 163.367
R597 B.n496 B.n282 163.367
R598 B.n496 B.n276 163.367
R599 B.n504 B.n276 163.367
R600 B.n504 B.n274 163.367
R601 B.n508 B.n274 163.367
R602 B.n508 B.n268 163.367
R603 B.n516 B.n268 163.367
R604 B.n516 B.n266 163.367
R605 B.n520 B.n266 163.367
R606 B.n520 B.n260 163.367
R607 B.n528 B.n260 163.367
R608 B.n528 B.n258 163.367
R609 B.n532 B.n258 163.367
R610 B.n532 B.n252 163.367
R611 B.n541 B.n252 163.367
R612 B.n541 B.n250 163.367
R613 B.n545 B.n250 163.367
R614 B.n545 B.n245 163.367
R615 B.n553 B.n245 163.367
R616 B.n553 B.n243 163.367
R617 B.n557 B.n243 163.367
R618 B.n557 B.n237 163.367
R619 B.n565 B.n237 163.367
R620 B.n565 B.n235 163.367
R621 B.n569 B.n235 163.367
R622 B.n569 B.n229 163.367
R623 B.n577 B.n229 163.367
R624 B.n577 B.n227 163.367
R625 B.n581 B.n227 163.367
R626 B.n581 B.n221 163.367
R627 B.n590 B.n221 163.367
R628 B.n590 B.n219 163.367
R629 B.n594 B.n219 163.367
R630 B.n594 B.n2 163.367
R631 B.n776 B.n2 163.367
R632 B.n776 B.n3 163.367
R633 B.n772 B.n3 163.367
R634 B.n772 B.n9 163.367
R635 B.n768 B.n9 163.367
R636 B.n768 B.n11 163.367
R637 B.n764 B.n11 163.367
R638 B.n764 B.n16 163.367
R639 B.n760 B.n16 163.367
R640 B.n760 B.n18 163.367
R641 B.n756 B.n18 163.367
R642 B.n756 B.n23 163.367
R643 B.n752 B.n23 163.367
R644 B.n752 B.n25 163.367
R645 B.n748 B.n25 163.367
R646 B.n748 B.n30 163.367
R647 B.n744 B.n30 163.367
R648 B.n744 B.n32 163.367
R649 B.n740 B.n32 163.367
R650 B.n740 B.n36 163.367
R651 B.n736 B.n36 163.367
R652 B.n736 B.n38 163.367
R653 B.n732 B.n38 163.367
R654 B.n732 B.n44 163.367
R655 B.n728 B.n44 163.367
R656 B.n728 B.n46 163.367
R657 B.n724 B.n46 163.367
R658 B.n724 B.n51 163.367
R659 B.n720 B.n51 163.367
R660 B.n720 B.n53 163.367
R661 B.n716 B.n53 163.367
R662 B.n716 B.n58 163.367
R663 B.n712 B.n58 163.367
R664 B.n712 B.n60 163.367
R665 B.n708 B.n60 163.367
R666 B.n708 B.n65 163.367
R667 B.n704 B.n65 163.367
R668 B.n704 B.n67 163.367
R669 B.n700 B.n67 163.367
R670 B.n700 B.n72 163.367
R671 B.n696 B.n72 163.367
R672 B.n696 B.n74 163.367
R673 B.n692 B.n74 163.367
R674 B.n692 B.n79 163.367
R675 B.n688 B.n79 163.367
R676 B.n688 B.n81 163.367
R677 B.n684 B.n81 163.367
R678 B.n684 B.n86 163.367
R679 B.n680 B.n86 163.367
R680 B.n680 B.n88 163.367
R681 B.n676 B.n88 163.367
R682 B.n676 B.n93 163.367
R683 B.n672 B.n93 163.367
R684 B.n672 B.n95 163.367
R685 B.n343 B.n342 163.367
R686 B.n430 B.n342 163.367
R687 B.n428 B.n427 163.367
R688 B.n424 B.n423 163.367
R689 B.n420 B.n419 163.367
R690 B.n416 B.n415 163.367
R691 B.n412 B.n411 163.367
R692 B.n408 B.n407 163.367
R693 B.n404 B.n403 163.367
R694 B.n399 B.n398 163.367
R695 B.n395 B.n394 163.367
R696 B.n391 B.n390 163.367
R697 B.n387 B.n386 163.367
R698 B.n383 B.n382 163.367
R699 B.n378 B.n377 163.367
R700 B.n374 B.n373 163.367
R701 B.n370 B.n369 163.367
R702 B.n366 B.n365 163.367
R703 B.n362 B.n361 163.367
R704 B.n358 B.n357 163.367
R705 B.n354 B.n353 163.367
R706 B.n350 B.n349 163.367
R707 B.n438 B.n320 163.367
R708 B.n442 B.n318 163.367
R709 B.n442 B.n312 163.367
R710 B.n450 B.n312 163.367
R711 B.n450 B.n310 163.367
R712 B.n454 B.n310 163.367
R713 B.n454 B.n303 163.367
R714 B.n462 B.n303 163.367
R715 B.n462 B.n301 163.367
R716 B.n466 B.n301 163.367
R717 B.n466 B.n296 163.367
R718 B.n474 B.n296 163.367
R719 B.n474 B.n294 163.367
R720 B.n478 B.n294 163.367
R721 B.n478 B.n288 163.367
R722 B.n486 B.n288 163.367
R723 B.n486 B.n286 163.367
R724 B.n490 B.n286 163.367
R725 B.n490 B.n280 163.367
R726 B.n498 B.n280 163.367
R727 B.n498 B.n278 163.367
R728 B.n502 B.n278 163.367
R729 B.n502 B.n272 163.367
R730 B.n510 B.n272 163.367
R731 B.n510 B.n270 163.367
R732 B.n514 B.n270 163.367
R733 B.n514 B.n264 163.367
R734 B.n522 B.n264 163.367
R735 B.n522 B.n262 163.367
R736 B.n526 B.n262 163.367
R737 B.n526 B.n256 163.367
R738 B.n534 B.n256 163.367
R739 B.n534 B.n254 163.367
R740 B.n538 B.n254 163.367
R741 B.n538 B.n249 163.367
R742 B.n547 B.n249 163.367
R743 B.n547 B.n247 163.367
R744 B.n551 B.n247 163.367
R745 B.n551 B.n241 163.367
R746 B.n559 B.n241 163.367
R747 B.n559 B.n239 163.367
R748 B.n563 B.n239 163.367
R749 B.n563 B.n233 163.367
R750 B.n571 B.n233 163.367
R751 B.n571 B.n231 163.367
R752 B.n575 B.n231 163.367
R753 B.n575 B.n225 163.367
R754 B.n583 B.n225 163.367
R755 B.n583 B.n223 163.367
R756 B.n588 B.n223 163.367
R757 B.n588 B.n217 163.367
R758 B.n596 B.n217 163.367
R759 B.n597 B.n596 163.367
R760 B.n597 B.n5 163.367
R761 B.n6 B.n5 163.367
R762 B.n7 B.n6 163.367
R763 B.n602 B.n7 163.367
R764 B.n602 B.n12 163.367
R765 B.n13 B.n12 163.367
R766 B.n14 B.n13 163.367
R767 B.n607 B.n14 163.367
R768 B.n607 B.n19 163.367
R769 B.n20 B.n19 163.367
R770 B.n21 B.n20 163.367
R771 B.n612 B.n21 163.367
R772 B.n612 B.n26 163.367
R773 B.n27 B.n26 163.367
R774 B.n28 B.n27 163.367
R775 B.n617 B.n28 163.367
R776 B.n617 B.n33 163.367
R777 B.n34 B.n33 163.367
R778 B.n35 B.n34 163.367
R779 B.n622 B.n35 163.367
R780 B.n622 B.n40 163.367
R781 B.n41 B.n40 163.367
R782 B.n42 B.n41 163.367
R783 B.n627 B.n42 163.367
R784 B.n627 B.n47 163.367
R785 B.n48 B.n47 163.367
R786 B.n49 B.n48 163.367
R787 B.n632 B.n49 163.367
R788 B.n632 B.n54 163.367
R789 B.n55 B.n54 163.367
R790 B.n56 B.n55 163.367
R791 B.n637 B.n56 163.367
R792 B.n637 B.n61 163.367
R793 B.n62 B.n61 163.367
R794 B.n63 B.n62 163.367
R795 B.n642 B.n63 163.367
R796 B.n642 B.n68 163.367
R797 B.n69 B.n68 163.367
R798 B.n70 B.n69 163.367
R799 B.n647 B.n70 163.367
R800 B.n647 B.n75 163.367
R801 B.n76 B.n75 163.367
R802 B.n77 B.n76 163.367
R803 B.n652 B.n77 163.367
R804 B.n652 B.n82 163.367
R805 B.n83 B.n82 163.367
R806 B.n84 B.n83 163.367
R807 B.n657 B.n84 163.367
R808 B.n657 B.n89 163.367
R809 B.n90 B.n89 163.367
R810 B.n91 B.n90 163.367
R811 B.n662 B.n91 163.367
R812 B.n662 B.n96 163.367
R813 B.n97 B.n96 163.367
R814 B.n131 B.n130 163.367
R815 B.n135 B.n134 163.367
R816 B.n139 B.n138 163.367
R817 B.n143 B.n142 163.367
R818 B.n147 B.n146 163.367
R819 B.n151 B.n150 163.367
R820 B.n155 B.n154 163.367
R821 B.n159 B.n158 163.367
R822 B.n163 B.n162 163.367
R823 B.n167 B.n166 163.367
R824 B.n171 B.n170 163.367
R825 B.n175 B.n174 163.367
R826 B.n179 B.n178 163.367
R827 B.n183 B.n182 163.367
R828 B.n187 B.n186 163.367
R829 B.n191 B.n190 163.367
R830 B.n195 B.n194 163.367
R831 B.n199 B.n198 163.367
R832 B.n203 B.n202 163.367
R833 B.n207 B.n206 163.367
R834 B.n211 B.n210 163.367
R835 B.n213 B.n120 163.367
R836 B.n437 B.n317 149.493
R837 B.n670 B.n669 149.493
R838 B.n347 B.t18 146.618
R839 B.n122 B.t16 146.618
R840 B.n345 B.t12 146.618
R841 B.n125 B.t9 146.618
R842 B.n443 B.n317 80.0433
R843 B.n443 B.n313 80.0433
R844 B.n449 B.n313 80.0433
R845 B.n449 B.n309 80.0433
R846 B.n455 B.n309 80.0433
R847 B.n455 B.n304 80.0433
R848 B.n461 B.n304 80.0433
R849 B.n461 B.n305 80.0433
R850 B.n467 B.n297 80.0433
R851 B.n473 B.n297 80.0433
R852 B.n473 B.n293 80.0433
R853 B.n479 B.n293 80.0433
R854 B.n479 B.n289 80.0433
R855 B.n485 B.n289 80.0433
R856 B.n485 B.n285 80.0433
R857 B.n491 B.n285 80.0433
R858 B.n491 B.n281 80.0433
R859 B.n497 B.n281 80.0433
R860 B.n497 B.n277 80.0433
R861 B.n503 B.n277 80.0433
R862 B.n503 B.n273 80.0433
R863 B.n509 B.n273 80.0433
R864 B.n515 B.n269 80.0433
R865 B.n515 B.n265 80.0433
R866 B.n521 B.n265 80.0433
R867 B.n521 B.n261 80.0433
R868 B.n527 B.n261 80.0433
R869 B.n527 B.n257 80.0433
R870 B.n533 B.n257 80.0433
R871 B.n533 B.n253 80.0433
R872 B.n540 B.n253 80.0433
R873 B.n540 B.n539 80.0433
R874 B.n546 B.n246 80.0433
R875 B.n552 B.n246 80.0433
R876 B.n552 B.n242 80.0433
R877 B.n558 B.n242 80.0433
R878 B.n558 B.n238 80.0433
R879 B.n564 B.n238 80.0433
R880 B.n564 B.n234 80.0433
R881 B.n570 B.n234 80.0433
R882 B.n570 B.n230 80.0433
R883 B.n576 B.n230 80.0433
R884 B.n582 B.n226 80.0433
R885 B.n582 B.n222 80.0433
R886 B.n589 B.n222 80.0433
R887 B.n589 B.n218 80.0433
R888 B.n595 B.n218 80.0433
R889 B.n595 B.n4 80.0433
R890 B.n775 B.n4 80.0433
R891 B.n775 B.n774 80.0433
R892 B.n774 B.n773 80.0433
R893 B.n773 B.n8 80.0433
R894 B.n767 B.n8 80.0433
R895 B.n767 B.n766 80.0433
R896 B.n766 B.n765 80.0433
R897 B.n765 B.n15 80.0433
R898 B.n759 B.n758 80.0433
R899 B.n758 B.n757 80.0433
R900 B.n757 B.n22 80.0433
R901 B.n751 B.n22 80.0433
R902 B.n751 B.n750 80.0433
R903 B.n750 B.n749 80.0433
R904 B.n749 B.n29 80.0433
R905 B.n743 B.n29 80.0433
R906 B.n743 B.n742 80.0433
R907 B.n742 B.n741 80.0433
R908 B.n735 B.n39 80.0433
R909 B.n735 B.n734 80.0433
R910 B.n734 B.n733 80.0433
R911 B.n733 B.n43 80.0433
R912 B.n727 B.n43 80.0433
R913 B.n727 B.n726 80.0433
R914 B.n726 B.n725 80.0433
R915 B.n725 B.n50 80.0433
R916 B.n719 B.n50 80.0433
R917 B.n719 B.n718 80.0433
R918 B.n717 B.n57 80.0433
R919 B.n711 B.n57 80.0433
R920 B.n711 B.n710 80.0433
R921 B.n710 B.n709 80.0433
R922 B.n709 B.n64 80.0433
R923 B.n703 B.n64 80.0433
R924 B.n703 B.n702 80.0433
R925 B.n702 B.n701 80.0433
R926 B.n701 B.n71 80.0433
R927 B.n695 B.n71 80.0433
R928 B.n695 B.n694 80.0433
R929 B.n694 B.n693 80.0433
R930 B.n693 B.n78 80.0433
R931 B.n687 B.n78 80.0433
R932 B.n686 B.n685 80.0433
R933 B.n685 B.n85 80.0433
R934 B.n679 B.n85 80.0433
R935 B.n679 B.n678 80.0433
R936 B.n678 B.n677 80.0433
R937 B.n677 B.n92 80.0433
R938 B.n671 B.n92 80.0433
R939 B.n671 B.n670 80.0433
R940 B.n347 B.n346 74.0854
R941 B.n345 B.n344 74.0854
R942 B.n125 B.n124 74.0854
R943 B.n122 B.n121 74.0854
R944 B.n436 B.n435 71.676
R945 B.n430 B.n321 71.676
R946 B.n427 B.n322 71.676
R947 B.n423 B.n323 71.676
R948 B.n419 B.n324 71.676
R949 B.n415 B.n325 71.676
R950 B.n411 B.n326 71.676
R951 B.n407 B.n327 71.676
R952 B.n403 B.n328 71.676
R953 B.n398 B.n329 71.676
R954 B.n394 B.n330 71.676
R955 B.n390 B.n331 71.676
R956 B.n386 B.n332 71.676
R957 B.n382 B.n333 71.676
R958 B.n377 B.n334 71.676
R959 B.n373 B.n335 71.676
R960 B.n369 B.n336 71.676
R961 B.n365 B.n337 71.676
R962 B.n361 B.n338 71.676
R963 B.n357 B.n339 71.676
R964 B.n353 B.n340 71.676
R965 B.n349 B.n341 71.676
R966 B.n127 B.n98 71.676
R967 B.n131 B.n99 71.676
R968 B.n135 B.n100 71.676
R969 B.n139 B.n101 71.676
R970 B.n143 B.n102 71.676
R971 B.n147 B.n103 71.676
R972 B.n151 B.n104 71.676
R973 B.n155 B.n105 71.676
R974 B.n159 B.n106 71.676
R975 B.n163 B.n107 71.676
R976 B.n167 B.n108 71.676
R977 B.n171 B.n109 71.676
R978 B.n175 B.n110 71.676
R979 B.n179 B.n111 71.676
R980 B.n183 B.n112 71.676
R981 B.n187 B.n113 71.676
R982 B.n191 B.n114 71.676
R983 B.n195 B.n115 71.676
R984 B.n199 B.n116 71.676
R985 B.n203 B.n117 71.676
R986 B.n207 B.n118 71.676
R987 B.n211 B.n119 71.676
R988 B.n668 B.n120 71.676
R989 B.n668 B.n667 71.676
R990 B.n213 B.n119 71.676
R991 B.n210 B.n118 71.676
R992 B.n206 B.n117 71.676
R993 B.n202 B.n116 71.676
R994 B.n198 B.n115 71.676
R995 B.n194 B.n114 71.676
R996 B.n190 B.n113 71.676
R997 B.n186 B.n112 71.676
R998 B.n182 B.n111 71.676
R999 B.n178 B.n110 71.676
R1000 B.n174 B.n109 71.676
R1001 B.n170 B.n108 71.676
R1002 B.n166 B.n107 71.676
R1003 B.n162 B.n106 71.676
R1004 B.n158 B.n105 71.676
R1005 B.n154 B.n104 71.676
R1006 B.n150 B.n103 71.676
R1007 B.n146 B.n102 71.676
R1008 B.n142 B.n101 71.676
R1009 B.n138 B.n100 71.676
R1010 B.n134 B.n99 71.676
R1011 B.n130 B.n98 71.676
R1012 B.n436 B.n343 71.676
R1013 B.n428 B.n321 71.676
R1014 B.n424 B.n322 71.676
R1015 B.n420 B.n323 71.676
R1016 B.n416 B.n324 71.676
R1017 B.n412 B.n325 71.676
R1018 B.n408 B.n326 71.676
R1019 B.n404 B.n327 71.676
R1020 B.n399 B.n328 71.676
R1021 B.n395 B.n329 71.676
R1022 B.n391 B.n330 71.676
R1023 B.n387 B.n331 71.676
R1024 B.n383 B.n332 71.676
R1025 B.n378 B.n333 71.676
R1026 B.n374 B.n334 71.676
R1027 B.n370 B.n335 71.676
R1028 B.n366 B.n336 71.676
R1029 B.n362 B.n337 71.676
R1030 B.n358 B.n338 71.676
R1031 B.n354 B.n339 71.676
R1032 B.n350 B.n340 71.676
R1033 B.n341 B.n320 71.676
R1034 B.n305 B.t11 69.4494
R1035 B.t7 B.n686 69.4494
R1036 B.n576 B.t5 62.3868
R1037 B.n759 B.t4 62.3868
R1038 B.n380 B.n347 59.5399
R1039 B.n401 B.n345 59.5399
R1040 B.n126 B.n125 59.5399
R1041 B.n123 B.n122 59.5399
R1042 B.t0 B.n269 55.3242
R1043 B.n718 B.t3 55.3242
R1044 B.n539 B.t2 43.5532
R1045 B.n39 B.t1 43.5532
R1046 B.n546 B.t2 36.4906
R1047 B.n741 B.t1 36.4906
R1048 B.n128 B.n94 33.8737
R1049 B.n666 B.n665 33.8737
R1050 B.n440 B.n439 33.8737
R1051 B.n434 B.n315 33.8737
R1052 B.n509 B.t0 24.7196
R1053 B.t3 B.n717 24.7196
R1054 B B.n777 18.0485
R1055 B.t5 B.n226 17.657
R1056 B.t4 B.n15 17.657
R1057 B.n129 B.n128 10.6151
R1058 B.n132 B.n129 10.6151
R1059 B.n133 B.n132 10.6151
R1060 B.n136 B.n133 10.6151
R1061 B.n137 B.n136 10.6151
R1062 B.n140 B.n137 10.6151
R1063 B.n141 B.n140 10.6151
R1064 B.n144 B.n141 10.6151
R1065 B.n145 B.n144 10.6151
R1066 B.n148 B.n145 10.6151
R1067 B.n149 B.n148 10.6151
R1068 B.n152 B.n149 10.6151
R1069 B.n153 B.n152 10.6151
R1070 B.n156 B.n153 10.6151
R1071 B.n157 B.n156 10.6151
R1072 B.n160 B.n157 10.6151
R1073 B.n161 B.n160 10.6151
R1074 B.n165 B.n164 10.6151
R1075 B.n168 B.n165 10.6151
R1076 B.n169 B.n168 10.6151
R1077 B.n172 B.n169 10.6151
R1078 B.n173 B.n172 10.6151
R1079 B.n176 B.n173 10.6151
R1080 B.n177 B.n176 10.6151
R1081 B.n180 B.n177 10.6151
R1082 B.n181 B.n180 10.6151
R1083 B.n185 B.n184 10.6151
R1084 B.n188 B.n185 10.6151
R1085 B.n189 B.n188 10.6151
R1086 B.n192 B.n189 10.6151
R1087 B.n193 B.n192 10.6151
R1088 B.n196 B.n193 10.6151
R1089 B.n197 B.n196 10.6151
R1090 B.n200 B.n197 10.6151
R1091 B.n201 B.n200 10.6151
R1092 B.n204 B.n201 10.6151
R1093 B.n205 B.n204 10.6151
R1094 B.n208 B.n205 10.6151
R1095 B.n209 B.n208 10.6151
R1096 B.n212 B.n209 10.6151
R1097 B.n214 B.n212 10.6151
R1098 B.n215 B.n214 10.6151
R1099 B.n666 B.n215 10.6151
R1100 B.n441 B.n440 10.6151
R1101 B.n441 B.n311 10.6151
R1102 B.n451 B.n311 10.6151
R1103 B.n452 B.n451 10.6151
R1104 B.n453 B.n452 10.6151
R1105 B.n453 B.n302 10.6151
R1106 B.n463 B.n302 10.6151
R1107 B.n464 B.n463 10.6151
R1108 B.n465 B.n464 10.6151
R1109 B.n465 B.n295 10.6151
R1110 B.n475 B.n295 10.6151
R1111 B.n476 B.n475 10.6151
R1112 B.n477 B.n476 10.6151
R1113 B.n477 B.n287 10.6151
R1114 B.n487 B.n287 10.6151
R1115 B.n488 B.n487 10.6151
R1116 B.n489 B.n488 10.6151
R1117 B.n489 B.n279 10.6151
R1118 B.n499 B.n279 10.6151
R1119 B.n500 B.n499 10.6151
R1120 B.n501 B.n500 10.6151
R1121 B.n501 B.n271 10.6151
R1122 B.n511 B.n271 10.6151
R1123 B.n512 B.n511 10.6151
R1124 B.n513 B.n512 10.6151
R1125 B.n513 B.n263 10.6151
R1126 B.n523 B.n263 10.6151
R1127 B.n524 B.n523 10.6151
R1128 B.n525 B.n524 10.6151
R1129 B.n525 B.n255 10.6151
R1130 B.n535 B.n255 10.6151
R1131 B.n536 B.n535 10.6151
R1132 B.n537 B.n536 10.6151
R1133 B.n537 B.n248 10.6151
R1134 B.n548 B.n248 10.6151
R1135 B.n549 B.n548 10.6151
R1136 B.n550 B.n549 10.6151
R1137 B.n550 B.n240 10.6151
R1138 B.n560 B.n240 10.6151
R1139 B.n561 B.n560 10.6151
R1140 B.n562 B.n561 10.6151
R1141 B.n562 B.n232 10.6151
R1142 B.n572 B.n232 10.6151
R1143 B.n573 B.n572 10.6151
R1144 B.n574 B.n573 10.6151
R1145 B.n574 B.n224 10.6151
R1146 B.n584 B.n224 10.6151
R1147 B.n585 B.n584 10.6151
R1148 B.n587 B.n585 10.6151
R1149 B.n587 B.n586 10.6151
R1150 B.n586 B.n216 10.6151
R1151 B.n598 B.n216 10.6151
R1152 B.n599 B.n598 10.6151
R1153 B.n600 B.n599 10.6151
R1154 B.n601 B.n600 10.6151
R1155 B.n603 B.n601 10.6151
R1156 B.n604 B.n603 10.6151
R1157 B.n605 B.n604 10.6151
R1158 B.n606 B.n605 10.6151
R1159 B.n608 B.n606 10.6151
R1160 B.n609 B.n608 10.6151
R1161 B.n610 B.n609 10.6151
R1162 B.n611 B.n610 10.6151
R1163 B.n613 B.n611 10.6151
R1164 B.n614 B.n613 10.6151
R1165 B.n615 B.n614 10.6151
R1166 B.n616 B.n615 10.6151
R1167 B.n618 B.n616 10.6151
R1168 B.n619 B.n618 10.6151
R1169 B.n620 B.n619 10.6151
R1170 B.n621 B.n620 10.6151
R1171 B.n623 B.n621 10.6151
R1172 B.n624 B.n623 10.6151
R1173 B.n625 B.n624 10.6151
R1174 B.n626 B.n625 10.6151
R1175 B.n628 B.n626 10.6151
R1176 B.n629 B.n628 10.6151
R1177 B.n630 B.n629 10.6151
R1178 B.n631 B.n630 10.6151
R1179 B.n633 B.n631 10.6151
R1180 B.n634 B.n633 10.6151
R1181 B.n635 B.n634 10.6151
R1182 B.n636 B.n635 10.6151
R1183 B.n638 B.n636 10.6151
R1184 B.n639 B.n638 10.6151
R1185 B.n640 B.n639 10.6151
R1186 B.n641 B.n640 10.6151
R1187 B.n643 B.n641 10.6151
R1188 B.n644 B.n643 10.6151
R1189 B.n645 B.n644 10.6151
R1190 B.n646 B.n645 10.6151
R1191 B.n648 B.n646 10.6151
R1192 B.n649 B.n648 10.6151
R1193 B.n650 B.n649 10.6151
R1194 B.n651 B.n650 10.6151
R1195 B.n653 B.n651 10.6151
R1196 B.n654 B.n653 10.6151
R1197 B.n655 B.n654 10.6151
R1198 B.n656 B.n655 10.6151
R1199 B.n658 B.n656 10.6151
R1200 B.n659 B.n658 10.6151
R1201 B.n660 B.n659 10.6151
R1202 B.n661 B.n660 10.6151
R1203 B.n663 B.n661 10.6151
R1204 B.n664 B.n663 10.6151
R1205 B.n665 B.n664 10.6151
R1206 B.n434 B.n433 10.6151
R1207 B.n433 B.n432 10.6151
R1208 B.n432 B.n431 10.6151
R1209 B.n431 B.n429 10.6151
R1210 B.n429 B.n426 10.6151
R1211 B.n426 B.n425 10.6151
R1212 B.n425 B.n422 10.6151
R1213 B.n422 B.n421 10.6151
R1214 B.n421 B.n418 10.6151
R1215 B.n418 B.n417 10.6151
R1216 B.n417 B.n414 10.6151
R1217 B.n414 B.n413 10.6151
R1218 B.n413 B.n410 10.6151
R1219 B.n410 B.n409 10.6151
R1220 B.n409 B.n406 10.6151
R1221 B.n406 B.n405 10.6151
R1222 B.n405 B.n402 10.6151
R1223 B.n400 B.n397 10.6151
R1224 B.n397 B.n396 10.6151
R1225 B.n396 B.n393 10.6151
R1226 B.n393 B.n392 10.6151
R1227 B.n392 B.n389 10.6151
R1228 B.n389 B.n388 10.6151
R1229 B.n388 B.n385 10.6151
R1230 B.n385 B.n384 10.6151
R1231 B.n384 B.n381 10.6151
R1232 B.n379 B.n376 10.6151
R1233 B.n376 B.n375 10.6151
R1234 B.n375 B.n372 10.6151
R1235 B.n372 B.n371 10.6151
R1236 B.n371 B.n368 10.6151
R1237 B.n368 B.n367 10.6151
R1238 B.n367 B.n364 10.6151
R1239 B.n364 B.n363 10.6151
R1240 B.n363 B.n360 10.6151
R1241 B.n360 B.n359 10.6151
R1242 B.n359 B.n356 10.6151
R1243 B.n356 B.n355 10.6151
R1244 B.n355 B.n352 10.6151
R1245 B.n352 B.n351 10.6151
R1246 B.n351 B.n348 10.6151
R1247 B.n348 B.n319 10.6151
R1248 B.n439 B.n319 10.6151
R1249 B.n445 B.n315 10.6151
R1250 B.n446 B.n445 10.6151
R1251 B.n447 B.n446 10.6151
R1252 B.n447 B.n307 10.6151
R1253 B.n457 B.n307 10.6151
R1254 B.n458 B.n457 10.6151
R1255 B.n459 B.n458 10.6151
R1256 B.n459 B.n299 10.6151
R1257 B.n469 B.n299 10.6151
R1258 B.n470 B.n469 10.6151
R1259 B.n471 B.n470 10.6151
R1260 B.n471 B.n291 10.6151
R1261 B.n481 B.n291 10.6151
R1262 B.n482 B.n481 10.6151
R1263 B.n483 B.n482 10.6151
R1264 B.n483 B.n283 10.6151
R1265 B.n493 B.n283 10.6151
R1266 B.n494 B.n493 10.6151
R1267 B.n495 B.n494 10.6151
R1268 B.n495 B.n275 10.6151
R1269 B.n505 B.n275 10.6151
R1270 B.n506 B.n505 10.6151
R1271 B.n507 B.n506 10.6151
R1272 B.n507 B.n267 10.6151
R1273 B.n517 B.n267 10.6151
R1274 B.n518 B.n517 10.6151
R1275 B.n519 B.n518 10.6151
R1276 B.n519 B.n259 10.6151
R1277 B.n529 B.n259 10.6151
R1278 B.n530 B.n529 10.6151
R1279 B.n531 B.n530 10.6151
R1280 B.n531 B.n251 10.6151
R1281 B.n542 B.n251 10.6151
R1282 B.n543 B.n542 10.6151
R1283 B.n544 B.n543 10.6151
R1284 B.n544 B.n244 10.6151
R1285 B.n554 B.n244 10.6151
R1286 B.n555 B.n554 10.6151
R1287 B.n556 B.n555 10.6151
R1288 B.n556 B.n236 10.6151
R1289 B.n566 B.n236 10.6151
R1290 B.n567 B.n566 10.6151
R1291 B.n568 B.n567 10.6151
R1292 B.n568 B.n228 10.6151
R1293 B.n578 B.n228 10.6151
R1294 B.n579 B.n578 10.6151
R1295 B.n580 B.n579 10.6151
R1296 B.n580 B.n220 10.6151
R1297 B.n591 B.n220 10.6151
R1298 B.n592 B.n591 10.6151
R1299 B.n593 B.n592 10.6151
R1300 B.n593 B.n0 10.6151
R1301 B.n771 B.n1 10.6151
R1302 B.n771 B.n770 10.6151
R1303 B.n770 B.n769 10.6151
R1304 B.n769 B.n10 10.6151
R1305 B.n763 B.n10 10.6151
R1306 B.n763 B.n762 10.6151
R1307 B.n762 B.n761 10.6151
R1308 B.n761 B.n17 10.6151
R1309 B.n755 B.n17 10.6151
R1310 B.n755 B.n754 10.6151
R1311 B.n754 B.n753 10.6151
R1312 B.n753 B.n24 10.6151
R1313 B.n747 B.n24 10.6151
R1314 B.n747 B.n746 10.6151
R1315 B.n746 B.n745 10.6151
R1316 B.n745 B.n31 10.6151
R1317 B.n739 B.n31 10.6151
R1318 B.n739 B.n738 10.6151
R1319 B.n738 B.n737 10.6151
R1320 B.n737 B.n37 10.6151
R1321 B.n731 B.n37 10.6151
R1322 B.n731 B.n730 10.6151
R1323 B.n730 B.n729 10.6151
R1324 B.n729 B.n45 10.6151
R1325 B.n723 B.n45 10.6151
R1326 B.n723 B.n722 10.6151
R1327 B.n722 B.n721 10.6151
R1328 B.n721 B.n52 10.6151
R1329 B.n715 B.n52 10.6151
R1330 B.n715 B.n714 10.6151
R1331 B.n714 B.n713 10.6151
R1332 B.n713 B.n59 10.6151
R1333 B.n707 B.n59 10.6151
R1334 B.n707 B.n706 10.6151
R1335 B.n706 B.n705 10.6151
R1336 B.n705 B.n66 10.6151
R1337 B.n699 B.n66 10.6151
R1338 B.n699 B.n698 10.6151
R1339 B.n698 B.n697 10.6151
R1340 B.n697 B.n73 10.6151
R1341 B.n691 B.n73 10.6151
R1342 B.n691 B.n690 10.6151
R1343 B.n690 B.n689 10.6151
R1344 B.n689 B.n80 10.6151
R1345 B.n683 B.n80 10.6151
R1346 B.n683 B.n682 10.6151
R1347 B.n682 B.n681 10.6151
R1348 B.n681 B.n87 10.6151
R1349 B.n675 B.n87 10.6151
R1350 B.n675 B.n674 10.6151
R1351 B.n674 B.n673 10.6151
R1352 B.n673 B.n94 10.6151
R1353 B.n467 B.t11 10.5944
R1354 B.n687 B.t7 10.5944
R1355 B.n161 B.n126 9.36635
R1356 B.n184 B.n123 9.36635
R1357 B.n402 B.n401 9.36635
R1358 B.n380 B.n379 9.36635
R1359 B.n777 B.n0 2.81026
R1360 B.n777 B.n1 2.81026
R1361 B.n164 B.n126 1.24928
R1362 B.n181 B.n123 1.24928
R1363 B.n401 B.n400 1.24928
R1364 B.n381 B.n380 1.24928
R1365 VP.n16 VP.n13 161.3
R1366 VP.n18 VP.n17 161.3
R1367 VP.n19 VP.n12 161.3
R1368 VP.n21 VP.n20 161.3
R1369 VP.n22 VP.n11 161.3
R1370 VP.n24 VP.n23 161.3
R1371 VP.n25 VP.n10 161.3
R1372 VP.n27 VP.n26 161.3
R1373 VP.n55 VP.n54 161.3
R1374 VP.n53 VP.n1 161.3
R1375 VP.n52 VP.n51 161.3
R1376 VP.n50 VP.n2 161.3
R1377 VP.n49 VP.n48 161.3
R1378 VP.n47 VP.n3 161.3
R1379 VP.n46 VP.n45 161.3
R1380 VP.n44 VP.n4 161.3
R1381 VP.n43 VP.n42 161.3
R1382 VP.n40 VP.n5 161.3
R1383 VP.n39 VP.n38 161.3
R1384 VP.n37 VP.n6 161.3
R1385 VP.n36 VP.n35 161.3
R1386 VP.n34 VP.n7 161.3
R1387 VP.n33 VP.n32 161.3
R1388 VP.n31 VP.n8 161.3
R1389 VP.n30 VP.n29 86.642
R1390 VP.n56 VP.n0 86.642
R1391 VP.n28 VP.n9 86.642
R1392 VP.n15 VP.n14 62.1829
R1393 VP.n15 VP.t0 60.1672
R1394 VP.n35 VP.n6 56.0336
R1395 VP.n48 VP.n2 56.0336
R1396 VP.n20 VP.n11 56.0336
R1397 VP.n30 VP.n28 46.1433
R1398 VP.n29 VP.t2 28.1057
R1399 VP.n41 VP.t5 28.1057
R1400 VP.n0 VP.t4 28.1057
R1401 VP.n9 VP.t1 28.1057
R1402 VP.n14 VP.t3 28.1057
R1403 VP.n39 VP.n6 24.9531
R1404 VP.n48 VP.n47 24.9531
R1405 VP.n20 VP.n19 24.9531
R1406 VP.n33 VP.n8 24.4675
R1407 VP.n34 VP.n33 24.4675
R1408 VP.n35 VP.n34 24.4675
R1409 VP.n40 VP.n39 24.4675
R1410 VP.n42 VP.n40 24.4675
R1411 VP.n46 VP.n4 24.4675
R1412 VP.n47 VP.n46 24.4675
R1413 VP.n52 VP.n2 24.4675
R1414 VP.n53 VP.n52 24.4675
R1415 VP.n54 VP.n53 24.4675
R1416 VP.n24 VP.n11 24.4675
R1417 VP.n25 VP.n24 24.4675
R1418 VP.n26 VP.n25 24.4675
R1419 VP.n18 VP.n13 24.4675
R1420 VP.n19 VP.n18 24.4675
R1421 VP.n42 VP.n41 12.234
R1422 VP.n41 VP.n4 12.234
R1423 VP.n14 VP.n13 12.234
R1424 VP.n29 VP.n8 3.42588
R1425 VP.n54 VP.n0 3.42588
R1426 VP.n26 VP.n9 3.42588
R1427 VP.n16 VP.n15 3.37057
R1428 VP.n28 VP.n27 0.354971
R1429 VP.n31 VP.n30 0.354971
R1430 VP.n56 VP.n55 0.354971
R1431 VP VP.n56 0.26696
R1432 VP.n17 VP.n16 0.189894
R1433 VP.n17 VP.n12 0.189894
R1434 VP.n21 VP.n12 0.189894
R1435 VP.n22 VP.n21 0.189894
R1436 VP.n23 VP.n22 0.189894
R1437 VP.n23 VP.n10 0.189894
R1438 VP.n27 VP.n10 0.189894
R1439 VP.n32 VP.n31 0.189894
R1440 VP.n32 VP.n7 0.189894
R1441 VP.n36 VP.n7 0.189894
R1442 VP.n37 VP.n36 0.189894
R1443 VP.n38 VP.n37 0.189894
R1444 VP.n38 VP.n5 0.189894
R1445 VP.n43 VP.n5 0.189894
R1446 VP.n44 VP.n43 0.189894
R1447 VP.n45 VP.n44 0.189894
R1448 VP.n45 VP.n3 0.189894
R1449 VP.n49 VP.n3 0.189894
R1450 VP.n50 VP.n49 0.189894
R1451 VP.n51 VP.n50 0.189894
R1452 VP.n51 VP.n1 0.189894
R1453 VP.n55 VP.n1 0.189894
R1454 VTAIL.n82 VTAIL.n68 289.615
R1455 VTAIL.n16 VTAIL.n2 289.615
R1456 VTAIL.n62 VTAIL.n48 289.615
R1457 VTAIL.n40 VTAIL.n26 289.615
R1458 VTAIL.n75 VTAIL.n74 185
R1459 VTAIL.n72 VTAIL.n71 185
R1460 VTAIL.n81 VTAIL.n80 185
R1461 VTAIL.n83 VTAIL.n82 185
R1462 VTAIL.n9 VTAIL.n8 185
R1463 VTAIL.n6 VTAIL.n5 185
R1464 VTAIL.n15 VTAIL.n14 185
R1465 VTAIL.n17 VTAIL.n16 185
R1466 VTAIL.n63 VTAIL.n62 185
R1467 VTAIL.n61 VTAIL.n60 185
R1468 VTAIL.n52 VTAIL.n51 185
R1469 VTAIL.n55 VTAIL.n54 185
R1470 VTAIL.n41 VTAIL.n40 185
R1471 VTAIL.n39 VTAIL.n38 185
R1472 VTAIL.n30 VTAIL.n29 185
R1473 VTAIL.n33 VTAIL.n32 185
R1474 VTAIL.t2 VTAIL.n73 147.888
R1475 VTAIL.t11 VTAIL.n7 147.888
R1476 VTAIL.t6 VTAIL.n53 147.888
R1477 VTAIL.t0 VTAIL.n31 147.888
R1478 VTAIL.n74 VTAIL.n71 104.615
R1479 VTAIL.n81 VTAIL.n71 104.615
R1480 VTAIL.n82 VTAIL.n81 104.615
R1481 VTAIL.n8 VTAIL.n5 104.615
R1482 VTAIL.n15 VTAIL.n5 104.615
R1483 VTAIL.n16 VTAIL.n15 104.615
R1484 VTAIL.n62 VTAIL.n61 104.615
R1485 VTAIL.n61 VTAIL.n51 104.615
R1486 VTAIL.n54 VTAIL.n51 104.615
R1487 VTAIL.n40 VTAIL.n39 104.615
R1488 VTAIL.n39 VTAIL.n29 104.615
R1489 VTAIL.n32 VTAIL.n29 104.615
R1490 VTAIL.n47 VTAIL.n46 61.2459
R1491 VTAIL.n25 VTAIL.n24 61.2459
R1492 VTAIL.n1 VTAIL.n0 61.2458
R1493 VTAIL.n23 VTAIL.n22 61.2458
R1494 VTAIL.n74 VTAIL.t2 52.3082
R1495 VTAIL.n8 VTAIL.t11 52.3082
R1496 VTAIL.n54 VTAIL.t6 52.3082
R1497 VTAIL.n32 VTAIL.t0 52.3082
R1498 VTAIL.n87 VTAIL.n86 36.646
R1499 VTAIL.n21 VTAIL.n20 36.646
R1500 VTAIL.n67 VTAIL.n66 36.646
R1501 VTAIL.n45 VTAIL.n44 36.646
R1502 VTAIL.n25 VTAIL.n23 22.4617
R1503 VTAIL.n87 VTAIL.n67 19.1686
R1504 VTAIL.n75 VTAIL.n73 15.6496
R1505 VTAIL.n9 VTAIL.n7 15.6496
R1506 VTAIL.n55 VTAIL.n53 15.6496
R1507 VTAIL.n33 VTAIL.n31 15.6496
R1508 VTAIL.n76 VTAIL.n72 12.8005
R1509 VTAIL.n10 VTAIL.n6 12.8005
R1510 VTAIL.n56 VTAIL.n52 12.8005
R1511 VTAIL.n34 VTAIL.n30 12.8005
R1512 VTAIL.n80 VTAIL.n79 12.0247
R1513 VTAIL.n14 VTAIL.n13 12.0247
R1514 VTAIL.n60 VTAIL.n59 12.0247
R1515 VTAIL.n38 VTAIL.n37 12.0247
R1516 VTAIL.n83 VTAIL.n70 11.249
R1517 VTAIL.n17 VTAIL.n4 11.249
R1518 VTAIL.n63 VTAIL.n50 11.249
R1519 VTAIL.n41 VTAIL.n28 11.249
R1520 VTAIL.n84 VTAIL.n68 10.4732
R1521 VTAIL.n18 VTAIL.n2 10.4732
R1522 VTAIL.n64 VTAIL.n48 10.4732
R1523 VTAIL.n42 VTAIL.n26 10.4732
R1524 VTAIL.n86 VTAIL.n85 9.45567
R1525 VTAIL.n20 VTAIL.n19 9.45567
R1526 VTAIL.n66 VTAIL.n65 9.45567
R1527 VTAIL.n44 VTAIL.n43 9.45567
R1528 VTAIL.n85 VTAIL.n84 9.3005
R1529 VTAIL.n70 VTAIL.n69 9.3005
R1530 VTAIL.n79 VTAIL.n78 9.3005
R1531 VTAIL.n77 VTAIL.n76 9.3005
R1532 VTAIL.n19 VTAIL.n18 9.3005
R1533 VTAIL.n4 VTAIL.n3 9.3005
R1534 VTAIL.n13 VTAIL.n12 9.3005
R1535 VTAIL.n11 VTAIL.n10 9.3005
R1536 VTAIL.n65 VTAIL.n64 9.3005
R1537 VTAIL.n50 VTAIL.n49 9.3005
R1538 VTAIL.n59 VTAIL.n58 9.3005
R1539 VTAIL.n57 VTAIL.n56 9.3005
R1540 VTAIL.n43 VTAIL.n42 9.3005
R1541 VTAIL.n28 VTAIL.n27 9.3005
R1542 VTAIL.n37 VTAIL.n36 9.3005
R1543 VTAIL.n35 VTAIL.n34 9.3005
R1544 VTAIL.n0 VTAIL.t1 4.86536
R1545 VTAIL.n0 VTAIL.t3 4.86536
R1546 VTAIL.n22 VTAIL.t10 4.86536
R1547 VTAIL.n22 VTAIL.t9 4.86536
R1548 VTAIL.n46 VTAIL.t8 4.86536
R1549 VTAIL.n46 VTAIL.t7 4.86536
R1550 VTAIL.n24 VTAIL.t4 4.86536
R1551 VTAIL.n24 VTAIL.t5 4.86536
R1552 VTAIL.n77 VTAIL.n73 4.40546
R1553 VTAIL.n11 VTAIL.n7 4.40546
R1554 VTAIL.n57 VTAIL.n53 4.40546
R1555 VTAIL.n35 VTAIL.n31 4.40546
R1556 VTAIL.n86 VTAIL.n68 3.49141
R1557 VTAIL.n20 VTAIL.n2 3.49141
R1558 VTAIL.n66 VTAIL.n48 3.49141
R1559 VTAIL.n44 VTAIL.n26 3.49141
R1560 VTAIL.n45 VTAIL.n25 3.2936
R1561 VTAIL.n67 VTAIL.n47 3.2936
R1562 VTAIL.n23 VTAIL.n21 3.2936
R1563 VTAIL.n84 VTAIL.n83 2.71565
R1564 VTAIL.n18 VTAIL.n17 2.71565
R1565 VTAIL.n64 VTAIL.n63 2.71565
R1566 VTAIL.n42 VTAIL.n41 2.71565
R1567 VTAIL VTAIL.n87 2.41214
R1568 VTAIL.n47 VTAIL.n45 2.11688
R1569 VTAIL.n21 VTAIL.n1 2.11688
R1570 VTAIL.n80 VTAIL.n70 1.93989
R1571 VTAIL.n14 VTAIL.n4 1.93989
R1572 VTAIL.n60 VTAIL.n50 1.93989
R1573 VTAIL.n38 VTAIL.n28 1.93989
R1574 VTAIL.n79 VTAIL.n72 1.16414
R1575 VTAIL.n13 VTAIL.n6 1.16414
R1576 VTAIL.n59 VTAIL.n52 1.16414
R1577 VTAIL.n37 VTAIL.n30 1.16414
R1578 VTAIL VTAIL.n1 0.881965
R1579 VTAIL.n76 VTAIL.n75 0.388379
R1580 VTAIL.n10 VTAIL.n9 0.388379
R1581 VTAIL.n56 VTAIL.n55 0.388379
R1582 VTAIL.n34 VTAIL.n33 0.388379
R1583 VTAIL.n78 VTAIL.n77 0.155672
R1584 VTAIL.n78 VTAIL.n69 0.155672
R1585 VTAIL.n85 VTAIL.n69 0.155672
R1586 VTAIL.n12 VTAIL.n11 0.155672
R1587 VTAIL.n12 VTAIL.n3 0.155672
R1588 VTAIL.n19 VTAIL.n3 0.155672
R1589 VTAIL.n65 VTAIL.n49 0.155672
R1590 VTAIL.n58 VTAIL.n49 0.155672
R1591 VTAIL.n58 VTAIL.n57 0.155672
R1592 VTAIL.n43 VTAIL.n27 0.155672
R1593 VTAIL.n36 VTAIL.n27 0.155672
R1594 VTAIL.n36 VTAIL.n35 0.155672
R1595 VDD1.n14 VDD1.n0 289.615
R1596 VDD1.n33 VDD1.n19 289.615
R1597 VDD1.n15 VDD1.n14 185
R1598 VDD1.n13 VDD1.n12 185
R1599 VDD1.n4 VDD1.n3 185
R1600 VDD1.n7 VDD1.n6 185
R1601 VDD1.n26 VDD1.n25 185
R1602 VDD1.n23 VDD1.n22 185
R1603 VDD1.n32 VDD1.n31 185
R1604 VDD1.n34 VDD1.n33 185
R1605 VDD1.t5 VDD1.n5 147.888
R1606 VDD1.t3 VDD1.n24 147.888
R1607 VDD1.n14 VDD1.n13 104.615
R1608 VDD1.n13 VDD1.n3 104.615
R1609 VDD1.n6 VDD1.n3 104.615
R1610 VDD1.n25 VDD1.n22 104.615
R1611 VDD1.n32 VDD1.n22 104.615
R1612 VDD1.n33 VDD1.n32 104.615
R1613 VDD1.n39 VDD1.n38 78.6925
R1614 VDD1.n41 VDD1.n40 77.9246
R1615 VDD1 VDD1.n18 55.8528
R1616 VDD1.n39 VDD1.n37 55.7392
R1617 VDD1.n6 VDD1.t5 52.3082
R1618 VDD1.n25 VDD1.t3 52.3082
R1619 VDD1.n41 VDD1.n39 40.1561
R1620 VDD1.n7 VDD1.n5 15.6496
R1621 VDD1.n26 VDD1.n24 15.6496
R1622 VDD1.n8 VDD1.n4 12.8005
R1623 VDD1.n27 VDD1.n23 12.8005
R1624 VDD1.n12 VDD1.n11 12.0247
R1625 VDD1.n31 VDD1.n30 12.0247
R1626 VDD1.n15 VDD1.n2 11.249
R1627 VDD1.n34 VDD1.n21 11.249
R1628 VDD1.n16 VDD1.n0 10.4732
R1629 VDD1.n35 VDD1.n19 10.4732
R1630 VDD1.n18 VDD1.n17 9.45567
R1631 VDD1.n37 VDD1.n36 9.45567
R1632 VDD1.n17 VDD1.n16 9.3005
R1633 VDD1.n2 VDD1.n1 9.3005
R1634 VDD1.n11 VDD1.n10 9.3005
R1635 VDD1.n9 VDD1.n8 9.3005
R1636 VDD1.n36 VDD1.n35 9.3005
R1637 VDD1.n21 VDD1.n20 9.3005
R1638 VDD1.n30 VDD1.n29 9.3005
R1639 VDD1.n28 VDD1.n27 9.3005
R1640 VDD1.n40 VDD1.t2 4.86536
R1641 VDD1.n40 VDD1.t4 4.86536
R1642 VDD1.n38 VDD1.t0 4.86536
R1643 VDD1.n38 VDD1.t1 4.86536
R1644 VDD1.n9 VDD1.n5 4.40546
R1645 VDD1.n28 VDD1.n24 4.40546
R1646 VDD1.n18 VDD1.n0 3.49141
R1647 VDD1.n37 VDD1.n19 3.49141
R1648 VDD1.n16 VDD1.n15 2.71565
R1649 VDD1.n35 VDD1.n34 2.71565
R1650 VDD1.n12 VDD1.n2 1.93989
R1651 VDD1.n31 VDD1.n21 1.93989
R1652 VDD1.n11 VDD1.n4 1.16414
R1653 VDD1.n30 VDD1.n23 1.16414
R1654 VDD1 VDD1.n41 0.765586
R1655 VDD1.n8 VDD1.n7 0.388379
R1656 VDD1.n27 VDD1.n26 0.388379
R1657 VDD1.n17 VDD1.n1 0.155672
R1658 VDD1.n10 VDD1.n1 0.155672
R1659 VDD1.n10 VDD1.n9 0.155672
R1660 VDD1.n29 VDD1.n28 0.155672
R1661 VDD1.n29 VDD1.n20 0.155672
R1662 VDD1.n36 VDD1.n20 0.155672
R1663 VN.n38 VN.n37 161.3
R1664 VN.n36 VN.n21 161.3
R1665 VN.n35 VN.n34 161.3
R1666 VN.n33 VN.n22 161.3
R1667 VN.n32 VN.n31 161.3
R1668 VN.n30 VN.n23 161.3
R1669 VN.n29 VN.n28 161.3
R1670 VN.n27 VN.n24 161.3
R1671 VN.n18 VN.n17 161.3
R1672 VN.n16 VN.n1 161.3
R1673 VN.n15 VN.n14 161.3
R1674 VN.n13 VN.n2 161.3
R1675 VN.n12 VN.n11 161.3
R1676 VN.n10 VN.n3 161.3
R1677 VN.n9 VN.n8 161.3
R1678 VN.n7 VN.n4 161.3
R1679 VN.n19 VN.n0 86.642
R1680 VN.n39 VN.n20 86.642
R1681 VN.n6 VN.n5 62.1829
R1682 VN.n26 VN.n25 62.1829
R1683 VN.n6 VN.t2 60.1673
R1684 VN.n26 VN.t3 60.1673
R1685 VN.n11 VN.n2 56.0336
R1686 VN.n31 VN.n22 56.0336
R1687 VN VN.n39 46.3086
R1688 VN.n5 VN.t1 28.1057
R1689 VN.n0 VN.t4 28.1057
R1690 VN.n25 VN.t5 28.1057
R1691 VN.n20 VN.t0 28.1057
R1692 VN.n11 VN.n10 24.9531
R1693 VN.n31 VN.n30 24.9531
R1694 VN.n9 VN.n4 24.4675
R1695 VN.n10 VN.n9 24.4675
R1696 VN.n15 VN.n2 24.4675
R1697 VN.n16 VN.n15 24.4675
R1698 VN.n17 VN.n16 24.4675
R1699 VN.n30 VN.n29 24.4675
R1700 VN.n29 VN.n24 24.4675
R1701 VN.n37 VN.n36 24.4675
R1702 VN.n36 VN.n35 24.4675
R1703 VN.n35 VN.n22 24.4675
R1704 VN.n5 VN.n4 12.234
R1705 VN.n25 VN.n24 12.234
R1706 VN.n17 VN.n0 3.42588
R1707 VN.n37 VN.n20 3.42588
R1708 VN.n27 VN.n26 3.37058
R1709 VN.n7 VN.n6 3.37058
R1710 VN.n39 VN.n38 0.354971
R1711 VN.n19 VN.n18 0.354971
R1712 VN VN.n19 0.26696
R1713 VN.n38 VN.n21 0.189894
R1714 VN.n34 VN.n21 0.189894
R1715 VN.n34 VN.n33 0.189894
R1716 VN.n33 VN.n32 0.189894
R1717 VN.n32 VN.n23 0.189894
R1718 VN.n28 VN.n23 0.189894
R1719 VN.n28 VN.n27 0.189894
R1720 VN.n8 VN.n7 0.189894
R1721 VN.n8 VN.n3 0.189894
R1722 VN.n12 VN.n3 0.189894
R1723 VN.n13 VN.n12 0.189894
R1724 VN.n14 VN.n13 0.189894
R1725 VN.n14 VN.n1 0.189894
R1726 VN.n18 VN.n1 0.189894
R1727 VDD2.n35 VDD2.n21 289.615
R1728 VDD2.n14 VDD2.n0 289.615
R1729 VDD2.n36 VDD2.n35 185
R1730 VDD2.n34 VDD2.n33 185
R1731 VDD2.n25 VDD2.n24 185
R1732 VDD2.n28 VDD2.n27 185
R1733 VDD2.n7 VDD2.n6 185
R1734 VDD2.n4 VDD2.n3 185
R1735 VDD2.n13 VDD2.n12 185
R1736 VDD2.n15 VDD2.n14 185
R1737 VDD2.t5 VDD2.n26 147.888
R1738 VDD2.t3 VDD2.n5 147.888
R1739 VDD2.n35 VDD2.n34 104.615
R1740 VDD2.n34 VDD2.n24 104.615
R1741 VDD2.n27 VDD2.n24 104.615
R1742 VDD2.n6 VDD2.n3 104.615
R1743 VDD2.n13 VDD2.n3 104.615
R1744 VDD2.n14 VDD2.n13 104.615
R1745 VDD2.n20 VDD2.n19 78.6925
R1746 VDD2 VDD2.n41 78.6897
R1747 VDD2.n20 VDD2.n18 55.7392
R1748 VDD2.n40 VDD2.n39 53.3247
R1749 VDD2.n27 VDD2.t5 52.3082
R1750 VDD2.n6 VDD2.t3 52.3082
R1751 VDD2.n40 VDD2.n20 37.9265
R1752 VDD2.n28 VDD2.n26 15.6496
R1753 VDD2.n7 VDD2.n5 15.6496
R1754 VDD2.n29 VDD2.n25 12.8005
R1755 VDD2.n8 VDD2.n4 12.8005
R1756 VDD2.n33 VDD2.n32 12.0247
R1757 VDD2.n12 VDD2.n11 12.0247
R1758 VDD2.n36 VDD2.n23 11.249
R1759 VDD2.n15 VDD2.n2 11.249
R1760 VDD2.n37 VDD2.n21 10.4732
R1761 VDD2.n16 VDD2.n0 10.4732
R1762 VDD2.n39 VDD2.n38 9.45567
R1763 VDD2.n18 VDD2.n17 9.45567
R1764 VDD2.n38 VDD2.n37 9.3005
R1765 VDD2.n23 VDD2.n22 9.3005
R1766 VDD2.n32 VDD2.n31 9.3005
R1767 VDD2.n30 VDD2.n29 9.3005
R1768 VDD2.n17 VDD2.n16 9.3005
R1769 VDD2.n2 VDD2.n1 9.3005
R1770 VDD2.n11 VDD2.n10 9.3005
R1771 VDD2.n9 VDD2.n8 9.3005
R1772 VDD2.n41 VDD2.t0 4.86536
R1773 VDD2.n41 VDD2.t2 4.86536
R1774 VDD2.n19 VDD2.t4 4.86536
R1775 VDD2.n19 VDD2.t1 4.86536
R1776 VDD2.n30 VDD2.n26 4.40546
R1777 VDD2.n9 VDD2.n5 4.40546
R1778 VDD2.n39 VDD2.n21 3.49141
R1779 VDD2.n18 VDD2.n0 3.49141
R1780 VDD2.n37 VDD2.n36 2.71565
R1781 VDD2.n16 VDD2.n15 2.71565
R1782 VDD2 VDD2.n40 2.52852
R1783 VDD2.n33 VDD2.n23 1.93989
R1784 VDD2.n12 VDD2.n2 1.93989
R1785 VDD2.n32 VDD2.n25 1.16414
R1786 VDD2.n11 VDD2.n4 1.16414
R1787 VDD2.n29 VDD2.n28 0.388379
R1788 VDD2.n8 VDD2.n7 0.388379
R1789 VDD2.n38 VDD2.n22 0.155672
R1790 VDD2.n31 VDD2.n22 0.155672
R1791 VDD2.n31 VDD2.n30 0.155672
R1792 VDD2.n10 VDD2.n9 0.155672
R1793 VDD2.n10 VDD2.n1 0.155672
R1794 VDD2.n17 VDD2.n1 0.155672
C0 VDD2 VDD1 1.75407f
C1 VTAIL VDD2 5.48309f
C2 VN VDD1 0.15627f
C3 VDD1 VP 3.03976f
C4 VTAIL VN 3.62856f
C5 VN VDD2 2.66055f
C6 VTAIL VP 3.64271f
C7 VDD2 VP 0.538205f
C8 VN VP 6.33419f
C9 VTAIL VDD1 5.42417f
C10 VDD2 B 5.262958f
C11 VDD1 B 5.434056f
C12 VTAIL B 4.738874f
C13 VN B 14.798719f
C14 VP B 13.435296f
C15 VDD2.n0 B 0.033052f
C16 VDD2.n1 B 0.022336f
C17 VDD2.n2 B 0.012002f
C18 VDD2.n3 B 0.028369f
C19 VDD2.n4 B 0.012708f
C20 VDD2.n5 B 0.087148f
C21 VDD2.t3 B 0.0474f
C22 VDD2.n6 B 0.021277f
C23 VDD2.n7 B 0.016697f
C24 VDD2.n8 B 0.012002f
C25 VDD2.n9 B 0.330265f
C26 VDD2.n10 B 0.022336f
C27 VDD2.n11 B 0.012002f
C28 VDD2.n12 B 0.012708f
C29 VDD2.n13 B 0.028369f
C30 VDD2.n14 B 0.064345f
C31 VDD2.n15 B 0.012708f
C32 VDD2.n16 B 0.012002f
C33 VDD2.n17 B 0.058645f
C34 VDD2.n18 B 0.061457f
C35 VDD2.t4 B 0.071836f
C36 VDD2.t1 B 0.071836f
C37 VDD2.n19 B 0.569886f
C38 VDD2.n20 B 2.30276f
C39 VDD2.n21 B 0.033052f
C40 VDD2.n22 B 0.022336f
C41 VDD2.n23 B 0.012002f
C42 VDD2.n24 B 0.028369f
C43 VDD2.n25 B 0.012708f
C44 VDD2.n26 B 0.087148f
C45 VDD2.t5 B 0.0474f
C46 VDD2.n27 B 0.021277f
C47 VDD2.n28 B 0.016697f
C48 VDD2.n29 B 0.012002f
C49 VDD2.n30 B 0.330265f
C50 VDD2.n31 B 0.022336f
C51 VDD2.n32 B 0.012002f
C52 VDD2.n33 B 0.012708f
C53 VDD2.n34 B 0.028369f
C54 VDD2.n35 B 0.064345f
C55 VDD2.n36 B 0.012708f
C56 VDD2.n37 B 0.012002f
C57 VDD2.n38 B 0.058645f
C58 VDD2.n39 B 0.051883f
C59 VDD2.n40 B 1.95548f
C60 VDD2.t0 B 0.071836f
C61 VDD2.t2 B 0.071836f
C62 VDD2.n41 B 0.569861f
C63 VN.t4 B 0.889515f
C64 VN.n0 B 0.430296f
C65 VN.n1 B 0.024339f
C66 VN.n2 B 0.041575f
C67 VN.n3 B 0.024339f
C68 VN.n4 B 0.034164f
C69 VN.t1 B 0.889515f
C70 VN.n5 B 0.428686f
C71 VN.t2 B 1.16925f
C72 VN.n6 B 0.425379f
C73 VN.n7 B 0.302462f
C74 VN.n8 B 0.024339f
C75 VN.n9 B 0.045362f
C76 VN.n10 B 0.045788f
C77 VN.n11 B 0.02906f
C78 VN.n12 B 0.024339f
C79 VN.n13 B 0.024339f
C80 VN.n14 B 0.024339f
C81 VN.n15 B 0.045362f
C82 VN.n16 B 0.045362f
C83 VN.n17 B 0.026102f
C84 VN.n18 B 0.039283f
C85 VN.n19 B 0.070216f
C86 VN.t0 B 0.889515f
C87 VN.n20 B 0.430296f
C88 VN.n21 B 0.024339f
C89 VN.n22 B 0.041575f
C90 VN.n23 B 0.024339f
C91 VN.n24 B 0.034164f
C92 VN.t3 B 1.16926f
C93 VN.t5 B 0.889515f
C94 VN.n25 B 0.428686f
C95 VN.n26 B 0.425379f
C96 VN.n27 B 0.302462f
C97 VN.n28 B 0.024339f
C98 VN.n29 B 0.045362f
C99 VN.n30 B 0.045788f
C100 VN.n31 B 0.02906f
C101 VN.n32 B 0.024339f
C102 VN.n33 B 0.024339f
C103 VN.n34 B 0.024339f
C104 VN.n35 B 0.045362f
C105 VN.n36 B 0.045362f
C106 VN.n37 B 0.026102f
C107 VN.n38 B 0.039283f
C108 VN.n39 B 1.25047f
C109 VDD1.n0 B 0.033521f
C110 VDD1.n1 B 0.022652f
C111 VDD1.n2 B 0.012172f
C112 VDD1.n3 B 0.028771f
C113 VDD1.n4 B 0.012889f
C114 VDD1.n5 B 0.088384f
C115 VDD1.t5 B 0.048072f
C116 VDD1.n6 B 0.021578f
C117 VDD1.n7 B 0.016934f
C118 VDD1.n8 B 0.012172f
C119 VDD1.n9 B 0.33495f
C120 VDD1.n10 B 0.022652f
C121 VDD1.n11 B 0.012172f
C122 VDD1.n12 B 0.012889f
C123 VDD1.n13 B 0.028771f
C124 VDD1.n14 B 0.065258f
C125 VDD1.n15 B 0.012889f
C126 VDD1.n16 B 0.012172f
C127 VDD1.n17 B 0.059478f
C128 VDD1.n18 B 0.06313f
C129 VDD1.n19 B 0.033521f
C130 VDD1.n20 B 0.022652f
C131 VDD1.n21 B 0.012172f
C132 VDD1.n22 B 0.028771f
C133 VDD1.n23 B 0.012889f
C134 VDD1.n24 B 0.088384f
C135 VDD1.t3 B 0.048072f
C136 VDD1.n25 B 0.021578f
C137 VDD1.n26 B 0.016934f
C138 VDD1.n27 B 0.012172f
C139 VDD1.n28 B 0.33495f
C140 VDD1.n29 B 0.022652f
C141 VDD1.n30 B 0.012172f
C142 VDD1.n31 B 0.012889f
C143 VDD1.n32 B 0.028771f
C144 VDD1.n33 B 0.065258f
C145 VDD1.n34 B 0.012889f
C146 VDD1.n35 B 0.012172f
C147 VDD1.n36 B 0.059478f
C148 VDD1.n37 B 0.062329f
C149 VDD1.t0 B 0.072856f
C150 VDD1.t1 B 0.072856f
C151 VDD1.n38 B 0.577971f
C152 VDD1.n39 B 2.46115f
C153 VDD1.t2 B 0.072856f
C154 VDD1.t4 B 0.072856f
C155 VDD1.n40 B 0.573249f
C156 VDD1.n41 B 2.19192f
C157 VTAIL.t1 B 0.098582f
C158 VTAIL.t3 B 0.098582f
C159 VTAIL.n0 B 0.711808f
C160 VTAIL.n1 B 0.558628f
C161 VTAIL.n2 B 0.045358f
C162 VTAIL.n3 B 0.030651f
C163 VTAIL.n4 B 0.016471f
C164 VTAIL.n5 B 0.038931f
C165 VTAIL.n6 B 0.017439f
C166 VTAIL.n7 B 0.119593f
C167 VTAIL.t11 B 0.065047f
C168 VTAIL.n8 B 0.029198f
C169 VTAIL.n9 B 0.022913f
C170 VTAIL.n10 B 0.016471f
C171 VTAIL.n11 B 0.453225f
C172 VTAIL.n12 B 0.030651f
C173 VTAIL.n13 B 0.016471f
C174 VTAIL.n14 B 0.017439f
C175 VTAIL.n15 B 0.038931f
C176 VTAIL.n16 B 0.088301f
C177 VTAIL.n17 B 0.017439f
C178 VTAIL.n18 B 0.016471f
C179 VTAIL.n19 B 0.08048f
C180 VTAIL.n20 B 0.050101f
C181 VTAIL.n21 B 0.5659f
C182 VTAIL.t10 B 0.098582f
C183 VTAIL.t9 B 0.098582f
C184 VTAIL.n22 B 0.711808f
C185 VTAIL.n23 B 2.00117f
C186 VTAIL.t4 B 0.098582f
C187 VTAIL.t5 B 0.098582f
C188 VTAIL.n24 B 0.711813f
C189 VTAIL.n25 B 2.00116f
C190 VTAIL.n26 B 0.045358f
C191 VTAIL.n27 B 0.030651f
C192 VTAIL.n28 B 0.016471f
C193 VTAIL.n29 B 0.038931f
C194 VTAIL.n30 B 0.017439f
C195 VTAIL.n31 B 0.119593f
C196 VTAIL.t0 B 0.065047f
C197 VTAIL.n32 B 0.029198f
C198 VTAIL.n33 B 0.022913f
C199 VTAIL.n34 B 0.016471f
C200 VTAIL.n35 B 0.453225f
C201 VTAIL.n36 B 0.030651f
C202 VTAIL.n37 B 0.016471f
C203 VTAIL.n38 B 0.017439f
C204 VTAIL.n39 B 0.038931f
C205 VTAIL.n40 B 0.088301f
C206 VTAIL.n41 B 0.017439f
C207 VTAIL.n42 B 0.016471f
C208 VTAIL.n43 B 0.08048f
C209 VTAIL.n44 B 0.050101f
C210 VTAIL.n45 B 0.5659f
C211 VTAIL.t8 B 0.098582f
C212 VTAIL.t7 B 0.098582f
C213 VTAIL.n46 B 0.711813f
C214 VTAIL.n47 B 0.79681f
C215 VTAIL.n48 B 0.045358f
C216 VTAIL.n49 B 0.030651f
C217 VTAIL.n50 B 0.016471f
C218 VTAIL.n51 B 0.038931f
C219 VTAIL.n52 B 0.017439f
C220 VTAIL.n53 B 0.119593f
C221 VTAIL.t6 B 0.065047f
C222 VTAIL.n54 B 0.029198f
C223 VTAIL.n55 B 0.022913f
C224 VTAIL.n56 B 0.016471f
C225 VTAIL.n57 B 0.453225f
C226 VTAIL.n58 B 0.030651f
C227 VTAIL.n59 B 0.016471f
C228 VTAIL.n60 B 0.017439f
C229 VTAIL.n61 B 0.038931f
C230 VTAIL.n62 B 0.088301f
C231 VTAIL.n63 B 0.017439f
C232 VTAIL.n64 B 0.016471f
C233 VTAIL.n65 B 0.08048f
C234 VTAIL.n66 B 0.050101f
C235 VTAIL.n67 B 1.44501f
C236 VTAIL.n68 B 0.045358f
C237 VTAIL.n69 B 0.030651f
C238 VTAIL.n70 B 0.016471f
C239 VTAIL.n71 B 0.038931f
C240 VTAIL.n72 B 0.017439f
C241 VTAIL.n73 B 0.119593f
C242 VTAIL.t2 B 0.065047f
C243 VTAIL.n74 B 0.029198f
C244 VTAIL.n75 B 0.022913f
C245 VTAIL.n76 B 0.016471f
C246 VTAIL.n77 B 0.453225f
C247 VTAIL.n78 B 0.030651f
C248 VTAIL.n79 B 0.016471f
C249 VTAIL.n80 B 0.017439f
C250 VTAIL.n81 B 0.038931f
C251 VTAIL.n82 B 0.088301f
C252 VTAIL.n83 B 0.017439f
C253 VTAIL.n84 B 0.016471f
C254 VTAIL.n85 B 0.08048f
C255 VTAIL.n86 B 0.050101f
C256 VTAIL.n87 B 1.35795f
C257 VP.t4 B 0.913174f
C258 VP.n0 B 0.441741f
C259 VP.n1 B 0.024986f
C260 VP.n2 B 0.042681f
C261 VP.n3 B 0.024986f
C262 VP.n4 B 0.035073f
C263 VP.n5 B 0.024986f
C264 VP.n6 B 0.029833f
C265 VP.n7 B 0.024986f
C266 VP.n8 B 0.026796f
C267 VP.t1 B 0.913174f
C268 VP.n9 B 0.441741f
C269 VP.n10 B 0.024986f
C270 VP.n11 B 0.042681f
C271 VP.n12 B 0.024986f
C272 VP.n13 B 0.035073f
C273 VP.t0 B 1.20035f
C274 VP.t3 B 0.913174f
C275 VP.n14 B 0.440087f
C276 VP.n15 B 0.436693f
C277 VP.n16 B 0.310507f
C278 VP.n17 B 0.024986f
C279 VP.n18 B 0.046568f
C280 VP.n19 B 0.047006f
C281 VP.n20 B 0.029833f
C282 VP.n21 B 0.024986f
C283 VP.n22 B 0.024986f
C284 VP.n23 B 0.024986f
C285 VP.n24 B 0.046568f
C286 VP.n25 B 0.046568f
C287 VP.n26 B 0.026796f
C288 VP.n27 B 0.040327f
C289 VP.n28 B 1.2732f
C290 VP.t2 B 0.913174f
C291 VP.n29 B 0.441741f
C292 VP.n30 B 1.29267f
C293 VP.n31 B 0.040327f
C294 VP.n32 B 0.024986f
C295 VP.n33 B 0.046568f
C296 VP.n34 B 0.046568f
C297 VP.n35 B 0.042681f
C298 VP.n36 B 0.024986f
C299 VP.n37 B 0.024986f
C300 VP.n38 B 0.024986f
C301 VP.n39 B 0.047006f
C302 VP.n40 B 0.046568f
C303 VP.t5 B 0.913174f
C304 VP.n41 B 0.354536f
C305 VP.n42 B 0.035073f
C306 VP.n43 B 0.024986f
C307 VP.n44 B 0.024986f
C308 VP.n45 B 0.024986f
C309 VP.n46 B 0.046568f
C310 VP.n47 B 0.047006f
C311 VP.n48 B 0.029833f
C312 VP.n49 B 0.024986f
C313 VP.n50 B 0.024986f
C314 VP.n51 B 0.024986f
C315 VP.n52 B 0.046568f
C316 VP.n53 B 0.046568f
C317 VP.n54 B 0.026796f
C318 VP.n55 B 0.040327f
C319 VP.n56 B 0.072084f
.ends

