* NGSPICE file created from diff_pair_sample_0888.ext - technology: sky130A

.subckt diff_pair_sample_0888 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X1 VDD2.t8 VN.t1 VTAIL.t18 B.t23 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X2 VTAIL.t3 VP.t0 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X3 VDD1.t8 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=6.6729 ps=35 w=17.11 l=0.31
X4 VTAIL.t17 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X5 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=0 ps=0 w=17.11 l=0.31
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=0 ps=0 w=17.11 l=0.31
X7 VDD2.t6 VN.t3 VTAIL.t16 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=2.82315 ps=17.44 w=17.11 l=0.31
X8 VDD2.t5 VN.t4 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=2.82315 ps=17.44 w=17.11 l=0.31
X9 VTAIL.t6 VP.t2 VDD1.t7 B.t20 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X10 VDD1.t6 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=2.82315 ps=17.44 w=17.11 l=0.31
X11 VTAIL.t4 VP.t4 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X12 VDD1.t4 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X13 VTAIL.t8 VP.t6 VDD1.t3 B.t22 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X14 VDD1.t2 VP.t7 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=2.82315 ps=17.44 w=17.11 l=0.31
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=0 ps=0 w=17.11 l=0.31
X16 VDD2.t4 VN.t5 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=6.6729 ps=35 w=17.11 l=0.31
X17 VDD1.t1 VP.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=6.6729 ps=35 w=17.11 l=0.31
X18 VTAIL.t13 VN.t6 VDD2.t1 B.t22 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X19 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6729 pd=35 as=0 ps=0 w=17.11 l=0.31
X20 VDD1.t0 VP.t9 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X21 VDD2.t0 VN.t7 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X22 VTAIL.t11 VN.t8 VDD2.t3 B.t20 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=2.82315 ps=17.44 w=17.11 l=0.31
X23 VDD2.t2 VN.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.82315 pd=17.44 as=6.6729 ps=35 w=17.11 l=0.31
R0 VN.n9 VN.t9 1472.9
R1 VN.n3 VN.t4 1472.9
R2 VN.n20 VN.t3 1472.9
R3 VN.n14 VN.t5 1472.9
R4 VN.n6 VN.t1 1432.01
R5 VN.n8 VN.t8 1432.01
R6 VN.n2 VN.t0 1432.01
R7 VN.n17 VN.t7 1432.01
R8 VN.n19 VN.t6 1432.01
R9 VN.n13 VN.t2 1432.01
R10 VN.n15 VN.n14 161.489
R11 VN.n4 VN.n3 161.489
R12 VN.n10 VN.n9 161.3
R13 VN.n21 VN.n20 161.3
R14 VN.n18 VN.n11 161.3
R15 VN.n17 VN.n16 161.3
R16 VN.n15 VN.n12 161.3
R17 VN.n7 VN.n0 161.3
R18 VN.n6 VN.n5 161.3
R19 VN.n4 VN.n1 161.3
R20 VN.n6 VN.n1 73.0308
R21 VN.n7 VN.n6 73.0308
R22 VN.n18 VN.n17 73.0308
R23 VN.n17 VN.n12 73.0308
R24 VN.n3 VN.n2 52.5823
R25 VN.n9 VN.n8 52.5823
R26 VN.n20 VN.n19 52.5823
R27 VN.n14 VN.n13 52.5823
R28 VN VN.n21 44.9872
R29 VN.n2 VN.n1 20.449
R30 VN.n8 VN.n7 20.449
R31 VN.n19 VN.n18 20.449
R32 VN.n13 VN.n12 20.449
R33 VN.n21 VN.n11 0.189894
R34 VN.n16 VN.n11 0.189894
R35 VN.n16 VN.n15 0.189894
R36 VN.n5 VN.n4 0.189894
R37 VN.n5 VN.n0 0.189894
R38 VN.n10 VN.n0 0.189894
R39 VN VN.n10 0.0516364
R40 VDD2.n1 VDD2.t5 61.4411
R41 VDD2.n4 VDD2.t6 60.8895
R42 VDD2.n3 VDD2.n2 60.0906
R43 VDD2 VDD2.n7 60.0878
R44 VDD2.n6 VDD2.n5 59.7324
R45 VDD2.n1 VDD2.n0 59.7321
R46 VDD2.n4 VDD2.n3 41.086
R47 VDD2.n7 VDD2.t7 1.15772
R48 VDD2.n7 VDD2.t4 1.15772
R49 VDD2.n5 VDD2.t1 1.15772
R50 VDD2.n5 VDD2.t0 1.15772
R51 VDD2.n2 VDD2.t3 1.15772
R52 VDD2.n2 VDD2.t2 1.15772
R53 VDD2.n0 VDD2.t9 1.15772
R54 VDD2.n0 VDD2.t8 1.15772
R55 VDD2.n6 VDD2.n4 0.552224
R56 VDD2 VDD2.n6 0.196621
R57 VDD2.n3 VDD2.n1 0.083085
R58 VTAIL.n11 VTAIL.t14 44.2107
R59 VTAIL.n17 VTAIL.t10 44.2106
R60 VTAIL.n2 VTAIL.t0 44.2106
R61 VTAIL.n16 VTAIL.t2 44.2106
R62 VTAIL.n15 VTAIL.n14 43.0536
R63 VTAIL.n13 VTAIL.n12 43.0536
R64 VTAIL.n10 VTAIL.n9 43.0536
R65 VTAIL.n8 VTAIL.n7 43.0536
R66 VTAIL.n19 VTAIL.n18 43.0533
R67 VTAIL.n1 VTAIL.n0 43.0533
R68 VTAIL.n4 VTAIL.n3 43.0533
R69 VTAIL.n6 VTAIL.n5 43.0533
R70 VTAIL.n8 VTAIL.n6 28.2203
R71 VTAIL.n17 VTAIL.n16 27.6686
R72 VTAIL.n18 VTAIL.t18 1.15772
R73 VTAIL.n18 VTAIL.t11 1.15772
R74 VTAIL.n0 VTAIL.t15 1.15772
R75 VTAIL.n0 VTAIL.t19 1.15772
R76 VTAIL.n3 VTAIL.t5 1.15772
R77 VTAIL.n3 VTAIL.t4 1.15772
R78 VTAIL.n5 VTAIL.t1 1.15772
R79 VTAIL.n5 VTAIL.t8 1.15772
R80 VTAIL.n14 VTAIL.t9 1.15772
R81 VTAIL.n14 VTAIL.t6 1.15772
R82 VTAIL.n12 VTAIL.t7 1.15772
R83 VTAIL.n12 VTAIL.t3 1.15772
R84 VTAIL.n9 VTAIL.t12 1.15772
R85 VTAIL.n9 VTAIL.t17 1.15772
R86 VTAIL.n7 VTAIL.t16 1.15772
R87 VTAIL.n7 VTAIL.t13 1.15772
R88 VTAIL.n13 VTAIL.n11 0.74619
R89 VTAIL.n2 VTAIL.n1 0.74619
R90 VTAIL.n10 VTAIL.n8 0.552224
R91 VTAIL.n11 VTAIL.n10 0.552224
R92 VTAIL.n15 VTAIL.n13 0.552224
R93 VTAIL.n16 VTAIL.n15 0.552224
R94 VTAIL.n6 VTAIL.n4 0.552224
R95 VTAIL.n4 VTAIL.n2 0.552224
R96 VTAIL.n19 VTAIL.n17 0.552224
R97 VTAIL VTAIL.n1 0.472483
R98 VTAIL VTAIL.n19 0.0802414
R99 B.n105 B.t14 1545.14
R100 B.n102 B.t10 1545.14
R101 B.n447 B.t17 1545.14
R102 B.n444 B.t6 1545.14
R103 B.n781 B.n780 585
R104 B.n782 B.n781 585
R105 B.n346 B.n100 585
R106 B.n345 B.n344 585
R107 B.n343 B.n342 585
R108 B.n341 B.n340 585
R109 B.n339 B.n338 585
R110 B.n337 B.n336 585
R111 B.n335 B.n334 585
R112 B.n333 B.n332 585
R113 B.n331 B.n330 585
R114 B.n329 B.n328 585
R115 B.n327 B.n326 585
R116 B.n325 B.n324 585
R117 B.n323 B.n322 585
R118 B.n321 B.n320 585
R119 B.n319 B.n318 585
R120 B.n317 B.n316 585
R121 B.n315 B.n314 585
R122 B.n313 B.n312 585
R123 B.n311 B.n310 585
R124 B.n309 B.n308 585
R125 B.n307 B.n306 585
R126 B.n305 B.n304 585
R127 B.n303 B.n302 585
R128 B.n301 B.n300 585
R129 B.n299 B.n298 585
R130 B.n297 B.n296 585
R131 B.n295 B.n294 585
R132 B.n293 B.n292 585
R133 B.n291 B.n290 585
R134 B.n289 B.n288 585
R135 B.n287 B.n286 585
R136 B.n285 B.n284 585
R137 B.n283 B.n282 585
R138 B.n281 B.n280 585
R139 B.n279 B.n278 585
R140 B.n277 B.n276 585
R141 B.n275 B.n274 585
R142 B.n273 B.n272 585
R143 B.n271 B.n270 585
R144 B.n269 B.n268 585
R145 B.n267 B.n266 585
R146 B.n265 B.n264 585
R147 B.n263 B.n262 585
R148 B.n261 B.n260 585
R149 B.n259 B.n258 585
R150 B.n257 B.n256 585
R151 B.n255 B.n254 585
R152 B.n253 B.n252 585
R153 B.n251 B.n250 585
R154 B.n249 B.n248 585
R155 B.n247 B.n246 585
R156 B.n245 B.n244 585
R157 B.n243 B.n242 585
R158 B.n241 B.n240 585
R159 B.n239 B.n238 585
R160 B.n237 B.n236 585
R161 B.n235 B.n234 585
R162 B.n233 B.n232 585
R163 B.n231 B.n230 585
R164 B.n229 B.n228 585
R165 B.n227 B.n226 585
R166 B.n225 B.n224 585
R167 B.n223 B.n222 585
R168 B.n221 B.n220 585
R169 B.n219 B.n218 585
R170 B.n216 B.n215 585
R171 B.n214 B.n213 585
R172 B.n212 B.n211 585
R173 B.n210 B.n209 585
R174 B.n208 B.n207 585
R175 B.n206 B.n205 585
R176 B.n204 B.n203 585
R177 B.n202 B.n201 585
R178 B.n200 B.n199 585
R179 B.n198 B.n197 585
R180 B.n196 B.n195 585
R181 B.n194 B.n193 585
R182 B.n192 B.n191 585
R183 B.n190 B.n189 585
R184 B.n188 B.n187 585
R185 B.n186 B.n185 585
R186 B.n184 B.n183 585
R187 B.n182 B.n181 585
R188 B.n180 B.n179 585
R189 B.n178 B.n177 585
R190 B.n176 B.n175 585
R191 B.n174 B.n173 585
R192 B.n172 B.n171 585
R193 B.n170 B.n169 585
R194 B.n168 B.n167 585
R195 B.n166 B.n165 585
R196 B.n164 B.n163 585
R197 B.n162 B.n161 585
R198 B.n160 B.n159 585
R199 B.n158 B.n157 585
R200 B.n156 B.n155 585
R201 B.n154 B.n153 585
R202 B.n152 B.n151 585
R203 B.n150 B.n149 585
R204 B.n148 B.n147 585
R205 B.n146 B.n145 585
R206 B.n144 B.n143 585
R207 B.n142 B.n141 585
R208 B.n140 B.n139 585
R209 B.n138 B.n137 585
R210 B.n136 B.n135 585
R211 B.n134 B.n133 585
R212 B.n132 B.n131 585
R213 B.n130 B.n129 585
R214 B.n128 B.n127 585
R215 B.n126 B.n125 585
R216 B.n124 B.n123 585
R217 B.n122 B.n121 585
R218 B.n120 B.n119 585
R219 B.n118 B.n117 585
R220 B.n116 B.n115 585
R221 B.n114 B.n113 585
R222 B.n112 B.n111 585
R223 B.n110 B.n109 585
R224 B.n108 B.n107 585
R225 B.n39 B.n38 585
R226 B.n785 B.n784 585
R227 B.n779 B.n101 585
R228 B.n101 B.n36 585
R229 B.n778 B.n35 585
R230 B.n789 B.n35 585
R231 B.n777 B.n34 585
R232 B.n790 B.n34 585
R233 B.n776 B.n33 585
R234 B.n791 B.n33 585
R235 B.n775 B.n774 585
R236 B.n774 B.n32 585
R237 B.n773 B.n28 585
R238 B.n797 B.n28 585
R239 B.n772 B.n27 585
R240 B.n798 B.n27 585
R241 B.n771 B.n26 585
R242 B.n799 B.n26 585
R243 B.n770 B.n769 585
R244 B.n769 B.n22 585
R245 B.n768 B.n21 585
R246 B.n805 B.n21 585
R247 B.n767 B.n20 585
R248 B.n806 B.n20 585
R249 B.n766 B.n19 585
R250 B.n807 B.n19 585
R251 B.n765 B.n764 585
R252 B.n764 B.n15 585
R253 B.n763 B.n14 585
R254 B.n813 B.n14 585
R255 B.n762 B.n13 585
R256 B.n814 B.n13 585
R257 B.n761 B.n12 585
R258 B.n815 B.n12 585
R259 B.n760 B.n759 585
R260 B.n759 B.n758 585
R261 B.n757 B.n756 585
R262 B.n757 B.n8 585
R263 B.n755 B.n7 585
R264 B.n822 B.n7 585
R265 B.n754 B.n6 585
R266 B.n823 B.n6 585
R267 B.n753 B.n5 585
R268 B.n824 B.n5 585
R269 B.n752 B.n751 585
R270 B.n751 B.n4 585
R271 B.n750 B.n347 585
R272 B.n750 B.n749 585
R273 B.n739 B.n348 585
R274 B.n742 B.n348 585
R275 B.n741 B.n740 585
R276 B.n743 B.n741 585
R277 B.n738 B.n353 585
R278 B.n353 B.n352 585
R279 B.n737 B.n736 585
R280 B.n736 B.n735 585
R281 B.n355 B.n354 585
R282 B.n356 B.n355 585
R283 B.n728 B.n727 585
R284 B.n729 B.n728 585
R285 B.n726 B.n361 585
R286 B.n361 B.n360 585
R287 B.n725 B.n724 585
R288 B.n724 B.n723 585
R289 B.n363 B.n362 585
R290 B.n364 B.n363 585
R291 B.n716 B.n715 585
R292 B.n717 B.n716 585
R293 B.n714 B.n369 585
R294 B.n369 B.n368 585
R295 B.n713 B.n712 585
R296 B.n712 B.n711 585
R297 B.n371 B.n370 585
R298 B.n704 B.n371 585
R299 B.n703 B.n702 585
R300 B.n705 B.n703 585
R301 B.n701 B.n376 585
R302 B.n376 B.n375 585
R303 B.n700 B.n699 585
R304 B.n699 B.n698 585
R305 B.n378 B.n377 585
R306 B.n379 B.n378 585
R307 B.n694 B.n693 585
R308 B.n382 B.n381 585
R309 B.n690 B.n689 585
R310 B.n691 B.n690 585
R311 B.n688 B.n443 585
R312 B.n687 B.n686 585
R313 B.n685 B.n684 585
R314 B.n683 B.n682 585
R315 B.n681 B.n680 585
R316 B.n679 B.n678 585
R317 B.n677 B.n676 585
R318 B.n675 B.n674 585
R319 B.n673 B.n672 585
R320 B.n671 B.n670 585
R321 B.n669 B.n668 585
R322 B.n667 B.n666 585
R323 B.n665 B.n664 585
R324 B.n663 B.n662 585
R325 B.n661 B.n660 585
R326 B.n659 B.n658 585
R327 B.n657 B.n656 585
R328 B.n655 B.n654 585
R329 B.n653 B.n652 585
R330 B.n651 B.n650 585
R331 B.n649 B.n648 585
R332 B.n647 B.n646 585
R333 B.n645 B.n644 585
R334 B.n643 B.n642 585
R335 B.n641 B.n640 585
R336 B.n639 B.n638 585
R337 B.n637 B.n636 585
R338 B.n635 B.n634 585
R339 B.n633 B.n632 585
R340 B.n631 B.n630 585
R341 B.n629 B.n628 585
R342 B.n627 B.n626 585
R343 B.n625 B.n624 585
R344 B.n623 B.n622 585
R345 B.n621 B.n620 585
R346 B.n619 B.n618 585
R347 B.n617 B.n616 585
R348 B.n615 B.n614 585
R349 B.n613 B.n612 585
R350 B.n611 B.n610 585
R351 B.n609 B.n608 585
R352 B.n607 B.n606 585
R353 B.n605 B.n604 585
R354 B.n603 B.n602 585
R355 B.n601 B.n600 585
R356 B.n599 B.n598 585
R357 B.n597 B.n596 585
R358 B.n595 B.n594 585
R359 B.n593 B.n592 585
R360 B.n591 B.n590 585
R361 B.n589 B.n588 585
R362 B.n587 B.n586 585
R363 B.n585 B.n584 585
R364 B.n583 B.n582 585
R365 B.n581 B.n580 585
R366 B.n579 B.n578 585
R367 B.n577 B.n576 585
R368 B.n575 B.n574 585
R369 B.n573 B.n572 585
R370 B.n571 B.n570 585
R371 B.n569 B.n568 585
R372 B.n567 B.n566 585
R373 B.n565 B.n564 585
R374 B.n562 B.n561 585
R375 B.n560 B.n559 585
R376 B.n558 B.n557 585
R377 B.n556 B.n555 585
R378 B.n554 B.n553 585
R379 B.n552 B.n551 585
R380 B.n550 B.n549 585
R381 B.n548 B.n547 585
R382 B.n546 B.n545 585
R383 B.n544 B.n543 585
R384 B.n542 B.n541 585
R385 B.n540 B.n539 585
R386 B.n538 B.n537 585
R387 B.n536 B.n535 585
R388 B.n534 B.n533 585
R389 B.n532 B.n531 585
R390 B.n530 B.n529 585
R391 B.n528 B.n527 585
R392 B.n526 B.n525 585
R393 B.n524 B.n523 585
R394 B.n522 B.n521 585
R395 B.n520 B.n519 585
R396 B.n518 B.n517 585
R397 B.n516 B.n515 585
R398 B.n514 B.n513 585
R399 B.n512 B.n511 585
R400 B.n510 B.n509 585
R401 B.n508 B.n507 585
R402 B.n506 B.n505 585
R403 B.n504 B.n503 585
R404 B.n502 B.n501 585
R405 B.n500 B.n499 585
R406 B.n498 B.n497 585
R407 B.n496 B.n495 585
R408 B.n494 B.n493 585
R409 B.n492 B.n491 585
R410 B.n490 B.n489 585
R411 B.n488 B.n487 585
R412 B.n486 B.n485 585
R413 B.n484 B.n483 585
R414 B.n482 B.n481 585
R415 B.n480 B.n479 585
R416 B.n478 B.n477 585
R417 B.n476 B.n475 585
R418 B.n474 B.n473 585
R419 B.n472 B.n471 585
R420 B.n470 B.n469 585
R421 B.n468 B.n467 585
R422 B.n466 B.n465 585
R423 B.n464 B.n463 585
R424 B.n462 B.n461 585
R425 B.n460 B.n459 585
R426 B.n458 B.n457 585
R427 B.n456 B.n455 585
R428 B.n454 B.n453 585
R429 B.n452 B.n451 585
R430 B.n450 B.n449 585
R431 B.n695 B.n380 585
R432 B.n380 B.n379 585
R433 B.n697 B.n696 585
R434 B.n698 B.n697 585
R435 B.n374 B.n373 585
R436 B.n375 B.n374 585
R437 B.n707 B.n706 585
R438 B.n706 B.n705 585
R439 B.n708 B.n372 585
R440 B.n704 B.n372 585
R441 B.n710 B.n709 585
R442 B.n711 B.n710 585
R443 B.n367 B.n366 585
R444 B.n368 B.n367 585
R445 B.n719 B.n718 585
R446 B.n718 B.n717 585
R447 B.n720 B.n365 585
R448 B.n365 B.n364 585
R449 B.n722 B.n721 585
R450 B.n723 B.n722 585
R451 B.n359 B.n358 585
R452 B.n360 B.n359 585
R453 B.n731 B.n730 585
R454 B.n730 B.n729 585
R455 B.n732 B.n357 585
R456 B.n357 B.n356 585
R457 B.n734 B.n733 585
R458 B.n735 B.n734 585
R459 B.n351 B.n350 585
R460 B.n352 B.n351 585
R461 B.n745 B.n744 585
R462 B.n744 B.n743 585
R463 B.n746 B.n349 585
R464 B.n742 B.n349 585
R465 B.n748 B.n747 585
R466 B.n749 B.n748 585
R467 B.n3 B.n0 585
R468 B.n4 B.n3 585
R469 B.n821 B.n1 585
R470 B.n822 B.n821 585
R471 B.n820 B.n819 585
R472 B.n820 B.n8 585
R473 B.n818 B.n9 585
R474 B.n758 B.n9 585
R475 B.n817 B.n816 585
R476 B.n816 B.n815 585
R477 B.n11 B.n10 585
R478 B.n814 B.n11 585
R479 B.n812 B.n811 585
R480 B.n813 B.n812 585
R481 B.n810 B.n16 585
R482 B.n16 B.n15 585
R483 B.n809 B.n808 585
R484 B.n808 B.n807 585
R485 B.n18 B.n17 585
R486 B.n806 B.n18 585
R487 B.n804 B.n803 585
R488 B.n805 B.n804 585
R489 B.n802 B.n23 585
R490 B.n23 B.n22 585
R491 B.n801 B.n800 585
R492 B.n800 B.n799 585
R493 B.n25 B.n24 585
R494 B.n798 B.n25 585
R495 B.n796 B.n795 585
R496 B.n797 B.n796 585
R497 B.n794 B.n29 585
R498 B.n32 B.n29 585
R499 B.n793 B.n792 585
R500 B.n792 B.n791 585
R501 B.n31 B.n30 585
R502 B.n790 B.n31 585
R503 B.n788 B.n787 585
R504 B.n789 B.n788 585
R505 B.n786 B.n37 585
R506 B.n37 B.n36 585
R507 B.n825 B.n824 585
R508 B.n823 B.n2 585
R509 B.n784 B.n37 473.281
R510 B.n781 B.n101 473.281
R511 B.n449 B.n378 473.281
R512 B.n693 B.n380 473.281
R513 B.n782 B.n99 256.663
R514 B.n782 B.n98 256.663
R515 B.n782 B.n97 256.663
R516 B.n782 B.n96 256.663
R517 B.n782 B.n95 256.663
R518 B.n782 B.n94 256.663
R519 B.n782 B.n93 256.663
R520 B.n782 B.n92 256.663
R521 B.n782 B.n91 256.663
R522 B.n782 B.n90 256.663
R523 B.n782 B.n89 256.663
R524 B.n782 B.n88 256.663
R525 B.n782 B.n87 256.663
R526 B.n782 B.n86 256.663
R527 B.n782 B.n85 256.663
R528 B.n782 B.n84 256.663
R529 B.n782 B.n83 256.663
R530 B.n782 B.n82 256.663
R531 B.n782 B.n81 256.663
R532 B.n782 B.n80 256.663
R533 B.n782 B.n79 256.663
R534 B.n782 B.n78 256.663
R535 B.n782 B.n77 256.663
R536 B.n782 B.n76 256.663
R537 B.n782 B.n75 256.663
R538 B.n782 B.n74 256.663
R539 B.n782 B.n73 256.663
R540 B.n782 B.n72 256.663
R541 B.n782 B.n71 256.663
R542 B.n782 B.n70 256.663
R543 B.n782 B.n69 256.663
R544 B.n782 B.n68 256.663
R545 B.n782 B.n67 256.663
R546 B.n782 B.n66 256.663
R547 B.n782 B.n65 256.663
R548 B.n782 B.n64 256.663
R549 B.n782 B.n63 256.663
R550 B.n782 B.n62 256.663
R551 B.n782 B.n61 256.663
R552 B.n782 B.n60 256.663
R553 B.n782 B.n59 256.663
R554 B.n782 B.n58 256.663
R555 B.n782 B.n57 256.663
R556 B.n782 B.n56 256.663
R557 B.n782 B.n55 256.663
R558 B.n782 B.n54 256.663
R559 B.n782 B.n53 256.663
R560 B.n782 B.n52 256.663
R561 B.n782 B.n51 256.663
R562 B.n782 B.n50 256.663
R563 B.n782 B.n49 256.663
R564 B.n782 B.n48 256.663
R565 B.n782 B.n47 256.663
R566 B.n782 B.n46 256.663
R567 B.n782 B.n45 256.663
R568 B.n782 B.n44 256.663
R569 B.n782 B.n43 256.663
R570 B.n782 B.n42 256.663
R571 B.n782 B.n41 256.663
R572 B.n782 B.n40 256.663
R573 B.n783 B.n782 256.663
R574 B.n692 B.n691 256.663
R575 B.n691 B.n383 256.663
R576 B.n691 B.n384 256.663
R577 B.n691 B.n385 256.663
R578 B.n691 B.n386 256.663
R579 B.n691 B.n387 256.663
R580 B.n691 B.n388 256.663
R581 B.n691 B.n389 256.663
R582 B.n691 B.n390 256.663
R583 B.n691 B.n391 256.663
R584 B.n691 B.n392 256.663
R585 B.n691 B.n393 256.663
R586 B.n691 B.n394 256.663
R587 B.n691 B.n395 256.663
R588 B.n691 B.n396 256.663
R589 B.n691 B.n397 256.663
R590 B.n691 B.n398 256.663
R591 B.n691 B.n399 256.663
R592 B.n691 B.n400 256.663
R593 B.n691 B.n401 256.663
R594 B.n691 B.n402 256.663
R595 B.n691 B.n403 256.663
R596 B.n691 B.n404 256.663
R597 B.n691 B.n405 256.663
R598 B.n691 B.n406 256.663
R599 B.n691 B.n407 256.663
R600 B.n691 B.n408 256.663
R601 B.n691 B.n409 256.663
R602 B.n691 B.n410 256.663
R603 B.n691 B.n411 256.663
R604 B.n691 B.n412 256.663
R605 B.n691 B.n413 256.663
R606 B.n691 B.n414 256.663
R607 B.n691 B.n415 256.663
R608 B.n691 B.n416 256.663
R609 B.n691 B.n417 256.663
R610 B.n691 B.n418 256.663
R611 B.n691 B.n419 256.663
R612 B.n691 B.n420 256.663
R613 B.n691 B.n421 256.663
R614 B.n691 B.n422 256.663
R615 B.n691 B.n423 256.663
R616 B.n691 B.n424 256.663
R617 B.n691 B.n425 256.663
R618 B.n691 B.n426 256.663
R619 B.n691 B.n427 256.663
R620 B.n691 B.n428 256.663
R621 B.n691 B.n429 256.663
R622 B.n691 B.n430 256.663
R623 B.n691 B.n431 256.663
R624 B.n691 B.n432 256.663
R625 B.n691 B.n433 256.663
R626 B.n691 B.n434 256.663
R627 B.n691 B.n435 256.663
R628 B.n691 B.n436 256.663
R629 B.n691 B.n437 256.663
R630 B.n691 B.n438 256.663
R631 B.n691 B.n439 256.663
R632 B.n691 B.n440 256.663
R633 B.n691 B.n441 256.663
R634 B.n691 B.n442 256.663
R635 B.n827 B.n826 256.663
R636 B.n107 B.n39 163.367
R637 B.n111 B.n110 163.367
R638 B.n115 B.n114 163.367
R639 B.n119 B.n118 163.367
R640 B.n123 B.n122 163.367
R641 B.n127 B.n126 163.367
R642 B.n131 B.n130 163.367
R643 B.n135 B.n134 163.367
R644 B.n139 B.n138 163.367
R645 B.n143 B.n142 163.367
R646 B.n147 B.n146 163.367
R647 B.n151 B.n150 163.367
R648 B.n155 B.n154 163.367
R649 B.n159 B.n158 163.367
R650 B.n163 B.n162 163.367
R651 B.n167 B.n166 163.367
R652 B.n171 B.n170 163.367
R653 B.n175 B.n174 163.367
R654 B.n179 B.n178 163.367
R655 B.n183 B.n182 163.367
R656 B.n187 B.n186 163.367
R657 B.n191 B.n190 163.367
R658 B.n195 B.n194 163.367
R659 B.n199 B.n198 163.367
R660 B.n203 B.n202 163.367
R661 B.n207 B.n206 163.367
R662 B.n211 B.n210 163.367
R663 B.n215 B.n214 163.367
R664 B.n220 B.n219 163.367
R665 B.n224 B.n223 163.367
R666 B.n228 B.n227 163.367
R667 B.n232 B.n231 163.367
R668 B.n236 B.n235 163.367
R669 B.n240 B.n239 163.367
R670 B.n244 B.n243 163.367
R671 B.n248 B.n247 163.367
R672 B.n252 B.n251 163.367
R673 B.n256 B.n255 163.367
R674 B.n260 B.n259 163.367
R675 B.n264 B.n263 163.367
R676 B.n268 B.n267 163.367
R677 B.n272 B.n271 163.367
R678 B.n276 B.n275 163.367
R679 B.n280 B.n279 163.367
R680 B.n284 B.n283 163.367
R681 B.n288 B.n287 163.367
R682 B.n292 B.n291 163.367
R683 B.n296 B.n295 163.367
R684 B.n300 B.n299 163.367
R685 B.n304 B.n303 163.367
R686 B.n308 B.n307 163.367
R687 B.n312 B.n311 163.367
R688 B.n316 B.n315 163.367
R689 B.n320 B.n319 163.367
R690 B.n324 B.n323 163.367
R691 B.n328 B.n327 163.367
R692 B.n332 B.n331 163.367
R693 B.n336 B.n335 163.367
R694 B.n340 B.n339 163.367
R695 B.n344 B.n343 163.367
R696 B.n781 B.n100 163.367
R697 B.n699 B.n378 163.367
R698 B.n699 B.n376 163.367
R699 B.n703 B.n376 163.367
R700 B.n703 B.n371 163.367
R701 B.n712 B.n371 163.367
R702 B.n712 B.n369 163.367
R703 B.n716 B.n369 163.367
R704 B.n716 B.n363 163.367
R705 B.n724 B.n363 163.367
R706 B.n724 B.n361 163.367
R707 B.n728 B.n361 163.367
R708 B.n728 B.n355 163.367
R709 B.n736 B.n355 163.367
R710 B.n736 B.n353 163.367
R711 B.n741 B.n353 163.367
R712 B.n741 B.n348 163.367
R713 B.n750 B.n348 163.367
R714 B.n751 B.n750 163.367
R715 B.n751 B.n5 163.367
R716 B.n6 B.n5 163.367
R717 B.n7 B.n6 163.367
R718 B.n757 B.n7 163.367
R719 B.n759 B.n757 163.367
R720 B.n759 B.n12 163.367
R721 B.n13 B.n12 163.367
R722 B.n14 B.n13 163.367
R723 B.n764 B.n14 163.367
R724 B.n764 B.n19 163.367
R725 B.n20 B.n19 163.367
R726 B.n21 B.n20 163.367
R727 B.n769 B.n21 163.367
R728 B.n769 B.n26 163.367
R729 B.n27 B.n26 163.367
R730 B.n28 B.n27 163.367
R731 B.n774 B.n28 163.367
R732 B.n774 B.n33 163.367
R733 B.n34 B.n33 163.367
R734 B.n35 B.n34 163.367
R735 B.n101 B.n35 163.367
R736 B.n690 B.n382 163.367
R737 B.n690 B.n443 163.367
R738 B.n686 B.n685 163.367
R739 B.n682 B.n681 163.367
R740 B.n678 B.n677 163.367
R741 B.n674 B.n673 163.367
R742 B.n670 B.n669 163.367
R743 B.n666 B.n665 163.367
R744 B.n662 B.n661 163.367
R745 B.n658 B.n657 163.367
R746 B.n654 B.n653 163.367
R747 B.n650 B.n649 163.367
R748 B.n646 B.n645 163.367
R749 B.n642 B.n641 163.367
R750 B.n638 B.n637 163.367
R751 B.n634 B.n633 163.367
R752 B.n630 B.n629 163.367
R753 B.n626 B.n625 163.367
R754 B.n622 B.n621 163.367
R755 B.n618 B.n617 163.367
R756 B.n614 B.n613 163.367
R757 B.n610 B.n609 163.367
R758 B.n606 B.n605 163.367
R759 B.n602 B.n601 163.367
R760 B.n598 B.n597 163.367
R761 B.n594 B.n593 163.367
R762 B.n590 B.n589 163.367
R763 B.n586 B.n585 163.367
R764 B.n582 B.n581 163.367
R765 B.n578 B.n577 163.367
R766 B.n574 B.n573 163.367
R767 B.n570 B.n569 163.367
R768 B.n566 B.n565 163.367
R769 B.n561 B.n560 163.367
R770 B.n557 B.n556 163.367
R771 B.n553 B.n552 163.367
R772 B.n549 B.n548 163.367
R773 B.n545 B.n544 163.367
R774 B.n541 B.n540 163.367
R775 B.n537 B.n536 163.367
R776 B.n533 B.n532 163.367
R777 B.n529 B.n528 163.367
R778 B.n525 B.n524 163.367
R779 B.n521 B.n520 163.367
R780 B.n517 B.n516 163.367
R781 B.n513 B.n512 163.367
R782 B.n509 B.n508 163.367
R783 B.n505 B.n504 163.367
R784 B.n501 B.n500 163.367
R785 B.n497 B.n496 163.367
R786 B.n493 B.n492 163.367
R787 B.n489 B.n488 163.367
R788 B.n485 B.n484 163.367
R789 B.n481 B.n480 163.367
R790 B.n477 B.n476 163.367
R791 B.n473 B.n472 163.367
R792 B.n469 B.n468 163.367
R793 B.n465 B.n464 163.367
R794 B.n461 B.n460 163.367
R795 B.n457 B.n456 163.367
R796 B.n453 B.n452 163.367
R797 B.n697 B.n380 163.367
R798 B.n697 B.n374 163.367
R799 B.n706 B.n374 163.367
R800 B.n706 B.n372 163.367
R801 B.n710 B.n372 163.367
R802 B.n710 B.n367 163.367
R803 B.n718 B.n367 163.367
R804 B.n718 B.n365 163.367
R805 B.n722 B.n365 163.367
R806 B.n722 B.n359 163.367
R807 B.n730 B.n359 163.367
R808 B.n730 B.n357 163.367
R809 B.n734 B.n357 163.367
R810 B.n734 B.n351 163.367
R811 B.n744 B.n351 163.367
R812 B.n744 B.n349 163.367
R813 B.n748 B.n349 163.367
R814 B.n748 B.n3 163.367
R815 B.n825 B.n3 163.367
R816 B.n821 B.n2 163.367
R817 B.n821 B.n820 163.367
R818 B.n820 B.n9 163.367
R819 B.n816 B.n9 163.367
R820 B.n816 B.n11 163.367
R821 B.n812 B.n11 163.367
R822 B.n812 B.n16 163.367
R823 B.n808 B.n16 163.367
R824 B.n808 B.n18 163.367
R825 B.n804 B.n18 163.367
R826 B.n804 B.n23 163.367
R827 B.n800 B.n23 163.367
R828 B.n800 B.n25 163.367
R829 B.n796 B.n25 163.367
R830 B.n796 B.n29 163.367
R831 B.n792 B.n29 163.367
R832 B.n792 B.n31 163.367
R833 B.n788 B.n31 163.367
R834 B.n788 B.n37 163.367
R835 B.n102 B.t12 81.8501
R836 B.n447 B.t19 81.8501
R837 B.n105 B.t15 81.8273
R838 B.n444 B.t9 81.8273
R839 B.n784 B.n783 71.676
R840 B.n107 B.n40 71.676
R841 B.n111 B.n41 71.676
R842 B.n115 B.n42 71.676
R843 B.n119 B.n43 71.676
R844 B.n123 B.n44 71.676
R845 B.n127 B.n45 71.676
R846 B.n131 B.n46 71.676
R847 B.n135 B.n47 71.676
R848 B.n139 B.n48 71.676
R849 B.n143 B.n49 71.676
R850 B.n147 B.n50 71.676
R851 B.n151 B.n51 71.676
R852 B.n155 B.n52 71.676
R853 B.n159 B.n53 71.676
R854 B.n163 B.n54 71.676
R855 B.n167 B.n55 71.676
R856 B.n171 B.n56 71.676
R857 B.n175 B.n57 71.676
R858 B.n179 B.n58 71.676
R859 B.n183 B.n59 71.676
R860 B.n187 B.n60 71.676
R861 B.n191 B.n61 71.676
R862 B.n195 B.n62 71.676
R863 B.n199 B.n63 71.676
R864 B.n203 B.n64 71.676
R865 B.n207 B.n65 71.676
R866 B.n211 B.n66 71.676
R867 B.n215 B.n67 71.676
R868 B.n220 B.n68 71.676
R869 B.n224 B.n69 71.676
R870 B.n228 B.n70 71.676
R871 B.n232 B.n71 71.676
R872 B.n236 B.n72 71.676
R873 B.n240 B.n73 71.676
R874 B.n244 B.n74 71.676
R875 B.n248 B.n75 71.676
R876 B.n252 B.n76 71.676
R877 B.n256 B.n77 71.676
R878 B.n260 B.n78 71.676
R879 B.n264 B.n79 71.676
R880 B.n268 B.n80 71.676
R881 B.n272 B.n81 71.676
R882 B.n276 B.n82 71.676
R883 B.n280 B.n83 71.676
R884 B.n284 B.n84 71.676
R885 B.n288 B.n85 71.676
R886 B.n292 B.n86 71.676
R887 B.n296 B.n87 71.676
R888 B.n300 B.n88 71.676
R889 B.n304 B.n89 71.676
R890 B.n308 B.n90 71.676
R891 B.n312 B.n91 71.676
R892 B.n316 B.n92 71.676
R893 B.n320 B.n93 71.676
R894 B.n324 B.n94 71.676
R895 B.n328 B.n95 71.676
R896 B.n332 B.n96 71.676
R897 B.n336 B.n97 71.676
R898 B.n340 B.n98 71.676
R899 B.n344 B.n99 71.676
R900 B.n100 B.n99 71.676
R901 B.n343 B.n98 71.676
R902 B.n339 B.n97 71.676
R903 B.n335 B.n96 71.676
R904 B.n331 B.n95 71.676
R905 B.n327 B.n94 71.676
R906 B.n323 B.n93 71.676
R907 B.n319 B.n92 71.676
R908 B.n315 B.n91 71.676
R909 B.n311 B.n90 71.676
R910 B.n307 B.n89 71.676
R911 B.n303 B.n88 71.676
R912 B.n299 B.n87 71.676
R913 B.n295 B.n86 71.676
R914 B.n291 B.n85 71.676
R915 B.n287 B.n84 71.676
R916 B.n283 B.n83 71.676
R917 B.n279 B.n82 71.676
R918 B.n275 B.n81 71.676
R919 B.n271 B.n80 71.676
R920 B.n267 B.n79 71.676
R921 B.n263 B.n78 71.676
R922 B.n259 B.n77 71.676
R923 B.n255 B.n76 71.676
R924 B.n251 B.n75 71.676
R925 B.n247 B.n74 71.676
R926 B.n243 B.n73 71.676
R927 B.n239 B.n72 71.676
R928 B.n235 B.n71 71.676
R929 B.n231 B.n70 71.676
R930 B.n227 B.n69 71.676
R931 B.n223 B.n68 71.676
R932 B.n219 B.n67 71.676
R933 B.n214 B.n66 71.676
R934 B.n210 B.n65 71.676
R935 B.n206 B.n64 71.676
R936 B.n202 B.n63 71.676
R937 B.n198 B.n62 71.676
R938 B.n194 B.n61 71.676
R939 B.n190 B.n60 71.676
R940 B.n186 B.n59 71.676
R941 B.n182 B.n58 71.676
R942 B.n178 B.n57 71.676
R943 B.n174 B.n56 71.676
R944 B.n170 B.n55 71.676
R945 B.n166 B.n54 71.676
R946 B.n162 B.n53 71.676
R947 B.n158 B.n52 71.676
R948 B.n154 B.n51 71.676
R949 B.n150 B.n50 71.676
R950 B.n146 B.n49 71.676
R951 B.n142 B.n48 71.676
R952 B.n138 B.n47 71.676
R953 B.n134 B.n46 71.676
R954 B.n130 B.n45 71.676
R955 B.n126 B.n44 71.676
R956 B.n122 B.n43 71.676
R957 B.n118 B.n42 71.676
R958 B.n114 B.n41 71.676
R959 B.n110 B.n40 71.676
R960 B.n783 B.n39 71.676
R961 B.n693 B.n692 71.676
R962 B.n443 B.n383 71.676
R963 B.n685 B.n384 71.676
R964 B.n681 B.n385 71.676
R965 B.n677 B.n386 71.676
R966 B.n673 B.n387 71.676
R967 B.n669 B.n388 71.676
R968 B.n665 B.n389 71.676
R969 B.n661 B.n390 71.676
R970 B.n657 B.n391 71.676
R971 B.n653 B.n392 71.676
R972 B.n649 B.n393 71.676
R973 B.n645 B.n394 71.676
R974 B.n641 B.n395 71.676
R975 B.n637 B.n396 71.676
R976 B.n633 B.n397 71.676
R977 B.n629 B.n398 71.676
R978 B.n625 B.n399 71.676
R979 B.n621 B.n400 71.676
R980 B.n617 B.n401 71.676
R981 B.n613 B.n402 71.676
R982 B.n609 B.n403 71.676
R983 B.n605 B.n404 71.676
R984 B.n601 B.n405 71.676
R985 B.n597 B.n406 71.676
R986 B.n593 B.n407 71.676
R987 B.n589 B.n408 71.676
R988 B.n585 B.n409 71.676
R989 B.n581 B.n410 71.676
R990 B.n577 B.n411 71.676
R991 B.n573 B.n412 71.676
R992 B.n569 B.n413 71.676
R993 B.n565 B.n414 71.676
R994 B.n560 B.n415 71.676
R995 B.n556 B.n416 71.676
R996 B.n552 B.n417 71.676
R997 B.n548 B.n418 71.676
R998 B.n544 B.n419 71.676
R999 B.n540 B.n420 71.676
R1000 B.n536 B.n421 71.676
R1001 B.n532 B.n422 71.676
R1002 B.n528 B.n423 71.676
R1003 B.n524 B.n424 71.676
R1004 B.n520 B.n425 71.676
R1005 B.n516 B.n426 71.676
R1006 B.n512 B.n427 71.676
R1007 B.n508 B.n428 71.676
R1008 B.n504 B.n429 71.676
R1009 B.n500 B.n430 71.676
R1010 B.n496 B.n431 71.676
R1011 B.n492 B.n432 71.676
R1012 B.n488 B.n433 71.676
R1013 B.n484 B.n434 71.676
R1014 B.n480 B.n435 71.676
R1015 B.n476 B.n436 71.676
R1016 B.n472 B.n437 71.676
R1017 B.n468 B.n438 71.676
R1018 B.n464 B.n439 71.676
R1019 B.n460 B.n440 71.676
R1020 B.n456 B.n441 71.676
R1021 B.n452 B.n442 71.676
R1022 B.n692 B.n382 71.676
R1023 B.n686 B.n383 71.676
R1024 B.n682 B.n384 71.676
R1025 B.n678 B.n385 71.676
R1026 B.n674 B.n386 71.676
R1027 B.n670 B.n387 71.676
R1028 B.n666 B.n388 71.676
R1029 B.n662 B.n389 71.676
R1030 B.n658 B.n390 71.676
R1031 B.n654 B.n391 71.676
R1032 B.n650 B.n392 71.676
R1033 B.n646 B.n393 71.676
R1034 B.n642 B.n394 71.676
R1035 B.n638 B.n395 71.676
R1036 B.n634 B.n396 71.676
R1037 B.n630 B.n397 71.676
R1038 B.n626 B.n398 71.676
R1039 B.n622 B.n399 71.676
R1040 B.n618 B.n400 71.676
R1041 B.n614 B.n401 71.676
R1042 B.n610 B.n402 71.676
R1043 B.n606 B.n403 71.676
R1044 B.n602 B.n404 71.676
R1045 B.n598 B.n405 71.676
R1046 B.n594 B.n406 71.676
R1047 B.n590 B.n407 71.676
R1048 B.n586 B.n408 71.676
R1049 B.n582 B.n409 71.676
R1050 B.n578 B.n410 71.676
R1051 B.n574 B.n411 71.676
R1052 B.n570 B.n412 71.676
R1053 B.n566 B.n413 71.676
R1054 B.n561 B.n414 71.676
R1055 B.n557 B.n415 71.676
R1056 B.n553 B.n416 71.676
R1057 B.n549 B.n417 71.676
R1058 B.n545 B.n418 71.676
R1059 B.n541 B.n419 71.676
R1060 B.n537 B.n420 71.676
R1061 B.n533 B.n421 71.676
R1062 B.n529 B.n422 71.676
R1063 B.n525 B.n423 71.676
R1064 B.n521 B.n424 71.676
R1065 B.n517 B.n425 71.676
R1066 B.n513 B.n426 71.676
R1067 B.n509 B.n427 71.676
R1068 B.n505 B.n428 71.676
R1069 B.n501 B.n429 71.676
R1070 B.n497 B.n430 71.676
R1071 B.n493 B.n431 71.676
R1072 B.n489 B.n432 71.676
R1073 B.n485 B.n433 71.676
R1074 B.n481 B.n434 71.676
R1075 B.n477 B.n435 71.676
R1076 B.n473 B.n436 71.676
R1077 B.n469 B.n437 71.676
R1078 B.n465 B.n438 71.676
R1079 B.n461 B.n439 71.676
R1080 B.n457 B.n440 71.676
R1081 B.n453 B.n441 71.676
R1082 B.n449 B.n442 71.676
R1083 B.n826 B.n825 71.676
R1084 B.n826 B.n2 71.676
R1085 B.n103 B.t13 69.4379
R1086 B.n448 B.t18 69.4379
R1087 B.n106 B.t16 69.4152
R1088 B.n445 B.t8 69.4152
R1089 B.n217 B.n106 59.5399
R1090 B.n104 B.n103 59.5399
R1091 B.n563 B.n448 59.5399
R1092 B.n446 B.n445 59.5399
R1093 B.n691 B.n379 57.4944
R1094 B.n782 B.n36 57.4944
R1095 B.n698 B.n379 33.4157
R1096 B.n698 B.n375 33.4157
R1097 B.n705 B.n375 33.4157
R1098 B.n705 B.n704 33.4157
R1099 B.n711 B.n368 33.4157
R1100 B.n717 B.n368 33.4157
R1101 B.n717 B.n364 33.4157
R1102 B.n723 B.n364 33.4157
R1103 B.n729 B.n360 33.4157
R1104 B.n735 B.n356 33.4157
R1105 B.n743 B.n352 33.4157
R1106 B.n749 B.n4 33.4157
R1107 B.n824 B.n4 33.4157
R1108 B.n824 B.n823 33.4157
R1109 B.n823 B.n822 33.4157
R1110 B.n822 B.n8 33.4157
R1111 B.n815 B.n814 33.4157
R1112 B.n813 B.n15 33.4157
R1113 B.n807 B.n806 33.4157
R1114 B.n805 B.n22 33.4157
R1115 B.n799 B.n22 33.4157
R1116 B.n799 B.n798 33.4157
R1117 B.n798 B.n797 33.4157
R1118 B.n791 B.n32 33.4157
R1119 B.n791 B.n790 33.4157
R1120 B.n790 B.n789 33.4157
R1121 B.n789 B.n36 33.4157
R1122 B.n742 B.t0 31.9415
R1123 B.n758 B.t21 31.9415
R1124 B.t4 B.n742 30.9587
R1125 B.n758 B.t3 30.9587
R1126 B.n695 B.n694 30.7517
R1127 B.n450 B.n377 30.7517
R1128 B.n780 B.n779 30.7517
R1129 B.n786 B.n785 30.7517
R1130 B.t5 B.n352 27.0275
R1131 B.n814 B.t23 27.0275
R1132 B.t22 B.n356 23.0963
R1133 B.t20 B.n15 23.0963
R1134 B.n711 B.t7 22.1135
R1135 B.n797 B.t11 22.1135
R1136 B.t1 B.n360 19.1651
R1137 B.n806 B.t2 19.1651
R1138 B B.n827 18.0485
R1139 B.n723 B.t1 14.2511
R1140 B.t2 B.n805 14.2511
R1141 B.n106 B.n105 12.4126
R1142 B.n103 B.n102 12.4126
R1143 B.n448 B.n447 12.4126
R1144 B.n445 B.n444 12.4126
R1145 B.n704 B.t7 11.3027
R1146 B.n32 B.t11 11.3027
R1147 B.n696 B.n695 10.6151
R1148 B.n696 B.n373 10.6151
R1149 B.n707 B.n373 10.6151
R1150 B.n708 B.n707 10.6151
R1151 B.n709 B.n708 10.6151
R1152 B.n709 B.n366 10.6151
R1153 B.n719 B.n366 10.6151
R1154 B.n720 B.n719 10.6151
R1155 B.n721 B.n720 10.6151
R1156 B.n721 B.n358 10.6151
R1157 B.n731 B.n358 10.6151
R1158 B.n732 B.n731 10.6151
R1159 B.n733 B.n732 10.6151
R1160 B.n733 B.n350 10.6151
R1161 B.n745 B.n350 10.6151
R1162 B.n746 B.n745 10.6151
R1163 B.n747 B.n746 10.6151
R1164 B.n747 B.n0 10.6151
R1165 B.n694 B.n381 10.6151
R1166 B.n689 B.n381 10.6151
R1167 B.n689 B.n688 10.6151
R1168 B.n688 B.n687 10.6151
R1169 B.n687 B.n684 10.6151
R1170 B.n684 B.n683 10.6151
R1171 B.n683 B.n680 10.6151
R1172 B.n680 B.n679 10.6151
R1173 B.n679 B.n676 10.6151
R1174 B.n676 B.n675 10.6151
R1175 B.n675 B.n672 10.6151
R1176 B.n672 B.n671 10.6151
R1177 B.n671 B.n668 10.6151
R1178 B.n668 B.n667 10.6151
R1179 B.n667 B.n664 10.6151
R1180 B.n664 B.n663 10.6151
R1181 B.n663 B.n660 10.6151
R1182 B.n660 B.n659 10.6151
R1183 B.n659 B.n656 10.6151
R1184 B.n656 B.n655 10.6151
R1185 B.n655 B.n652 10.6151
R1186 B.n652 B.n651 10.6151
R1187 B.n651 B.n648 10.6151
R1188 B.n648 B.n647 10.6151
R1189 B.n647 B.n644 10.6151
R1190 B.n644 B.n643 10.6151
R1191 B.n643 B.n640 10.6151
R1192 B.n640 B.n639 10.6151
R1193 B.n639 B.n636 10.6151
R1194 B.n636 B.n635 10.6151
R1195 B.n635 B.n632 10.6151
R1196 B.n632 B.n631 10.6151
R1197 B.n631 B.n628 10.6151
R1198 B.n628 B.n627 10.6151
R1199 B.n627 B.n624 10.6151
R1200 B.n624 B.n623 10.6151
R1201 B.n623 B.n620 10.6151
R1202 B.n620 B.n619 10.6151
R1203 B.n619 B.n616 10.6151
R1204 B.n616 B.n615 10.6151
R1205 B.n615 B.n612 10.6151
R1206 B.n612 B.n611 10.6151
R1207 B.n611 B.n608 10.6151
R1208 B.n608 B.n607 10.6151
R1209 B.n607 B.n604 10.6151
R1210 B.n604 B.n603 10.6151
R1211 B.n603 B.n600 10.6151
R1212 B.n600 B.n599 10.6151
R1213 B.n599 B.n596 10.6151
R1214 B.n596 B.n595 10.6151
R1215 B.n595 B.n592 10.6151
R1216 B.n592 B.n591 10.6151
R1217 B.n591 B.n588 10.6151
R1218 B.n588 B.n587 10.6151
R1219 B.n587 B.n584 10.6151
R1220 B.n584 B.n583 10.6151
R1221 B.n580 B.n579 10.6151
R1222 B.n579 B.n576 10.6151
R1223 B.n576 B.n575 10.6151
R1224 B.n575 B.n572 10.6151
R1225 B.n572 B.n571 10.6151
R1226 B.n571 B.n568 10.6151
R1227 B.n568 B.n567 10.6151
R1228 B.n567 B.n564 10.6151
R1229 B.n562 B.n559 10.6151
R1230 B.n559 B.n558 10.6151
R1231 B.n558 B.n555 10.6151
R1232 B.n555 B.n554 10.6151
R1233 B.n554 B.n551 10.6151
R1234 B.n551 B.n550 10.6151
R1235 B.n550 B.n547 10.6151
R1236 B.n547 B.n546 10.6151
R1237 B.n546 B.n543 10.6151
R1238 B.n543 B.n542 10.6151
R1239 B.n542 B.n539 10.6151
R1240 B.n539 B.n538 10.6151
R1241 B.n538 B.n535 10.6151
R1242 B.n535 B.n534 10.6151
R1243 B.n534 B.n531 10.6151
R1244 B.n531 B.n530 10.6151
R1245 B.n530 B.n527 10.6151
R1246 B.n527 B.n526 10.6151
R1247 B.n526 B.n523 10.6151
R1248 B.n523 B.n522 10.6151
R1249 B.n522 B.n519 10.6151
R1250 B.n519 B.n518 10.6151
R1251 B.n518 B.n515 10.6151
R1252 B.n515 B.n514 10.6151
R1253 B.n514 B.n511 10.6151
R1254 B.n511 B.n510 10.6151
R1255 B.n510 B.n507 10.6151
R1256 B.n507 B.n506 10.6151
R1257 B.n506 B.n503 10.6151
R1258 B.n503 B.n502 10.6151
R1259 B.n502 B.n499 10.6151
R1260 B.n499 B.n498 10.6151
R1261 B.n498 B.n495 10.6151
R1262 B.n495 B.n494 10.6151
R1263 B.n494 B.n491 10.6151
R1264 B.n491 B.n490 10.6151
R1265 B.n490 B.n487 10.6151
R1266 B.n487 B.n486 10.6151
R1267 B.n486 B.n483 10.6151
R1268 B.n483 B.n482 10.6151
R1269 B.n482 B.n479 10.6151
R1270 B.n479 B.n478 10.6151
R1271 B.n478 B.n475 10.6151
R1272 B.n475 B.n474 10.6151
R1273 B.n474 B.n471 10.6151
R1274 B.n471 B.n470 10.6151
R1275 B.n470 B.n467 10.6151
R1276 B.n467 B.n466 10.6151
R1277 B.n466 B.n463 10.6151
R1278 B.n463 B.n462 10.6151
R1279 B.n462 B.n459 10.6151
R1280 B.n459 B.n458 10.6151
R1281 B.n458 B.n455 10.6151
R1282 B.n455 B.n454 10.6151
R1283 B.n454 B.n451 10.6151
R1284 B.n451 B.n450 10.6151
R1285 B.n700 B.n377 10.6151
R1286 B.n701 B.n700 10.6151
R1287 B.n702 B.n701 10.6151
R1288 B.n702 B.n370 10.6151
R1289 B.n713 B.n370 10.6151
R1290 B.n714 B.n713 10.6151
R1291 B.n715 B.n714 10.6151
R1292 B.n715 B.n362 10.6151
R1293 B.n725 B.n362 10.6151
R1294 B.n726 B.n725 10.6151
R1295 B.n727 B.n726 10.6151
R1296 B.n727 B.n354 10.6151
R1297 B.n737 B.n354 10.6151
R1298 B.n738 B.n737 10.6151
R1299 B.n740 B.n738 10.6151
R1300 B.n740 B.n739 10.6151
R1301 B.n739 B.n347 10.6151
R1302 B.n752 B.n347 10.6151
R1303 B.n753 B.n752 10.6151
R1304 B.n754 B.n753 10.6151
R1305 B.n755 B.n754 10.6151
R1306 B.n756 B.n755 10.6151
R1307 B.n760 B.n756 10.6151
R1308 B.n761 B.n760 10.6151
R1309 B.n762 B.n761 10.6151
R1310 B.n763 B.n762 10.6151
R1311 B.n765 B.n763 10.6151
R1312 B.n766 B.n765 10.6151
R1313 B.n767 B.n766 10.6151
R1314 B.n768 B.n767 10.6151
R1315 B.n770 B.n768 10.6151
R1316 B.n771 B.n770 10.6151
R1317 B.n772 B.n771 10.6151
R1318 B.n773 B.n772 10.6151
R1319 B.n775 B.n773 10.6151
R1320 B.n776 B.n775 10.6151
R1321 B.n777 B.n776 10.6151
R1322 B.n778 B.n777 10.6151
R1323 B.n779 B.n778 10.6151
R1324 B.n819 B.n1 10.6151
R1325 B.n819 B.n818 10.6151
R1326 B.n818 B.n817 10.6151
R1327 B.n817 B.n10 10.6151
R1328 B.n811 B.n10 10.6151
R1329 B.n811 B.n810 10.6151
R1330 B.n810 B.n809 10.6151
R1331 B.n809 B.n17 10.6151
R1332 B.n803 B.n17 10.6151
R1333 B.n803 B.n802 10.6151
R1334 B.n802 B.n801 10.6151
R1335 B.n801 B.n24 10.6151
R1336 B.n795 B.n24 10.6151
R1337 B.n795 B.n794 10.6151
R1338 B.n794 B.n793 10.6151
R1339 B.n793 B.n30 10.6151
R1340 B.n787 B.n30 10.6151
R1341 B.n787 B.n786 10.6151
R1342 B.n785 B.n38 10.6151
R1343 B.n108 B.n38 10.6151
R1344 B.n109 B.n108 10.6151
R1345 B.n112 B.n109 10.6151
R1346 B.n113 B.n112 10.6151
R1347 B.n116 B.n113 10.6151
R1348 B.n117 B.n116 10.6151
R1349 B.n120 B.n117 10.6151
R1350 B.n121 B.n120 10.6151
R1351 B.n124 B.n121 10.6151
R1352 B.n125 B.n124 10.6151
R1353 B.n128 B.n125 10.6151
R1354 B.n129 B.n128 10.6151
R1355 B.n132 B.n129 10.6151
R1356 B.n133 B.n132 10.6151
R1357 B.n136 B.n133 10.6151
R1358 B.n137 B.n136 10.6151
R1359 B.n140 B.n137 10.6151
R1360 B.n141 B.n140 10.6151
R1361 B.n144 B.n141 10.6151
R1362 B.n145 B.n144 10.6151
R1363 B.n148 B.n145 10.6151
R1364 B.n149 B.n148 10.6151
R1365 B.n152 B.n149 10.6151
R1366 B.n153 B.n152 10.6151
R1367 B.n156 B.n153 10.6151
R1368 B.n157 B.n156 10.6151
R1369 B.n160 B.n157 10.6151
R1370 B.n161 B.n160 10.6151
R1371 B.n164 B.n161 10.6151
R1372 B.n165 B.n164 10.6151
R1373 B.n168 B.n165 10.6151
R1374 B.n169 B.n168 10.6151
R1375 B.n172 B.n169 10.6151
R1376 B.n173 B.n172 10.6151
R1377 B.n176 B.n173 10.6151
R1378 B.n177 B.n176 10.6151
R1379 B.n180 B.n177 10.6151
R1380 B.n181 B.n180 10.6151
R1381 B.n184 B.n181 10.6151
R1382 B.n185 B.n184 10.6151
R1383 B.n188 B.n185 10.6151
R1384 B.n189 B.n188 10.6151
R1385 B.n192 B.n189 10.6151
R1386 B.n193 B.n192 10.6151
R1387 B.n196 B.n193 10.6151
R1388 B.n197 B.n196 10.6151
R1389 B.n200 B.n197 10.6151
R1390 B.n201 B.n200 10.6151
R1391 B.n204 B.n201 10.6151
R1392 B.n205 B.n204 10.6151
R1393 B.n208 B.n205 10.6151
R1394 B.n209 B.n208 10.6151
R1395 B.n212 B.n209 10.6151
R1396 B.n213 B.n212 10.6151
R1397 B.n216 B.n213 10.6151
R1398 B.n221 B.n218 10.6151
R1399 B.n222 B.n221 10.6151
R1400 B.n225 B.n222 10.6151
R1401 B.n226 B.n225 10.6151
R1402 B.n229 B.n226 10.6151
R1403 B.n230 B.n229 10.6151
R1404 B.n233 B.n230 10.6151
R1405 B.n234 B.n233 10.6151
R1406 B.n238 B.n237 10.6151
R1407 B.n241 B.n238 10.6151
R1408 B.n242 B.n241 10.6151
R1409 B.n245 B.n242 10.6151
R1410 B.n246 B.n245 10.6151
R1411 B.n249 B.n246 10.6151
R1412 B.n250 B.n249 10.6151
R1413 B.n253 B.n250 10.6151
R1414 B.n254 B.n253 10.6151
R1415 B.n257 B.n254 10.6151
R1416 B.n258 B.n257 10.6151
R1417 B.n261 B.n258 10.6151
R1418 B.n262 B.n261 10.6151
R1419 B.n265 B.n262 10.6151
R1420 B.n266 B.n265 10.6151
R1421 B.n269 B.n266 10.6151
R1422 B.n270 B.n269 10.6151
R1423 B.n273 B.n270 10.6151
R1424 B.n274 B.n273 10.6151
R1425 B.n277 B.n274 10.6151
R1426 B.n278 B.n277 10.6151
R1427 B.n281 B.n278 10.6151
R1428 B.n282 B.n281 10.6151
R1429 B.n285 B.n282 10.6151
R1430 B.n286 B.n285 10.6151
R1431 B.n289 B.n286 10.6151
R1432 B.n290 B.n289 10.6151
R1433 B.n293 B.n290 10.6151
R1434 B.n294 B.n293 10.6151
R1435 B.n297 B.n294 10.6151
R1436 B.n298 B.n297 10.6151
R1437 B.n301 B.n298 10.6151
R1438 B.n302 B.n301 10.6151
R1439 B.n305 B.n302 10.6151
R1440 B.n306 B.n305 10.6151
R1441 B.n309 B.n306 10.6151
R1442 B.n310 B.n309 10.6151
R1443 B.n313 B.n310 10.6151
R1444 B.n314 B.n313 10.6151
R1445 B.n317 B.n314 10.6151
R1446 B.n318 B.n317 10.6151
R1447 B.n321 B.n318 10.6151
R1448 B.n322 B.n321 10.6151
R1449 B.n325 B.n322 10.6151
R1450 B.n326 B.n325 10.6151
R1451 B.n329 B.n326 10.6151
R1452 B.n330 B.n329 10.6151
R1453 B.n333 B.n330 10.6151
R1454 B.n334 B.n333 10.6151
R1455 B.n337 B.n334 10.6151
R1456 B.n338 B.n337 10.6151
R1457 B.n341 B.n338 10.6151
R1458 B.n342 B.n341 10.6151
R1459 B.n345 B.n342 10.6151
R1460 B.n346 B.n345 10.6151
R1461 B.n780 B.n346 10.6151
R1462 B.n729 B.t22 10.3199
R1463 B.n807 B.t20 10.3199
R1464 B.n827 B.n0 8.11757
R1465 B.n827 B.n1 8.11757
R1466 B.n580 B.n446 6.5566
R1467 B.n564 B.n563 6.5566
R1468 B.n218 B.n217 6.5566
R1469 B.n234 B.n104 6.5566
R1470 B.n735 B.t5 6.38871
R1471 B.t23 B.n813 6.38871
R1472 B.n583 B.n446 4.05904
R1473 B.n563 B.n562 4.05904
R1474 B.n217 B.n216 4.05904
R1475 B.n237 B.n104 4.05904
R1476 B.n743 B.t4 2.4575
R1477 B.n815 B.t3 2.4575
R1478 B.n749 B.t0 1.4747
R1479 B.t21 B.n8 1.4747
R1480 VP.n21 VP.t8 1472.9
R1481 VP.n14 VP.t3 1472.9
R1482 VP.n5 VP.t7 1472.9
R1483 VP.n11 VP.t1 1472.9
R1484 VP.n18 VP.t5 1432.01
R1485 VP.n20 VP.t4 1432.01
R1486 VP.n13 VP.t6 1432.01
R1487 VP.n8 VP.t9 1432.01
R1488 VP.n4 VP.t0 1432.01
R1489 VP.n10 VP.t2 1432.01
R1490 VP.n6 VP.n5 161.489
R1491 VP.n22 VP.n21 161.3
R1492 VP.n6 VP.n3 161.3
R1493 VP.n8 VP.n7 161.3
R1494 VP.n9 VP.n2 161.3
R1495 VP.n12 VP.n11 161.3
R1496 VP.n19 VP.n0 161.3
R1497 VP.n18 VP.n17 161.3
R1498 VP.n16 VP.n1 161.3
R1499 VP.n15 VP.n14 161.3
R1500 VP.n18 VP.n1 73.0308
R1501 VP.n19 VP.n18 73.0308
R1502 VP.n8 VP.n3 73.0308
R1503 VP.n9 VP.n8 73.0308
R1504 VP.n14 VP.n13 52.5823
R1505 VP.n21 VP.n20 52.5823
R1506 VP.n5 VP.n4 52.5823
R1507 VP.n11 VP.n10 52.5823
R1508 VP.n15 VP.n12 44.6066
R1509 VP.n13 VP.n1 20.449
R1510 VP.n20 VP.n19 20.449
R1511 VP.n4 VP.n3 20.449
R1512 VP.n10 VP.n9 20.449
R1513 VP.n7 VP.n6 0.189894
R1514 VP.n7 VP.n2 0.189894
R1515 VP.n12 VP.n2 0.189894
R1516 VP.n16 VP.n15 0.189894
R1517 VP.n17 VP.n16 0.189894
R1518 VP.n17 VP.n0 0.189894
R1519 VP.n22 VP.n0 0.189894
R1520 VP VP.n22 0.0516364
R1521 VDD1.n1 VDD1.t2 61.4413
R1522 VDD1.n3 VDD1.t6 61.4411
R1523 VDD1.n5 VDD1.n4 60.0906
R1524 VDD1.n1 VDD1.n0 59.7324
R1525 VDD1.n7 VDD1.n6 59.7322
R1526 VDD1.n3 VDD1.n2 59.7321
R1527 VDD1.n7 VDD1.n5 41.9449
R1528 VDD1.n6 VDD1.t7 1.15772
R1529 VDD1.n6 VDD1.t8 1.15772
R1530 VDD1.n0 VDD1.t9 1.15772
R1531 VDD1.n0 VDD1.t0 1.15772
R1532 VDD1.n4 VDD1.t5 1.15772
R1533 VDD1.n4 VDD1.t1 1.15772
R1534 VDD1.n2 VDD1.t3 1.15772
R1535 VDD1.n2 VDD1.t4 1.15772
R1536 VDD1 VDD1.n7 0.356103
R1537 VDD1 VDD1.n1 0.196621
R1538 VDD1.n5 VDD1.n3 0.083085
C0 VDD2 VDD1 0.733253f
C1 VP VTAIL 5.05257f
C2 VP VN 5.96833f
C3 VP VDD2 0.292854f
C4 VP VDD1 5.77534f
C5 VN VTAIL 5.03754f
C6 VDD2 VTAIL 28.4943f
C7 VDD1 VTAIL 28.4681f
C8 VN VDD2 5.63777f
C9 VN VDD1 0.148018f
C10 VDD2 B 5.462409f
C11 VDD1 B 5.31894f
C12 VTAIL B 7.829703f
C13 VN B 8.51637f
C14 VP B 5.967411f
C15 VDD1.t2 B 4.67936f
C16 VDD1.t9 B 0.402785f
C17 VDD1.t0 B 0.402785f
C18 VDD1.n0 B 3.66007f
C19 VDD1.n1 B 0.712536f
C20 VDD1.t6 B 4.67934f
C21 VDD1.t3 B 0.402785f
C22 VDD1.t4 B 0.402785f
C23 VDD1.n2 B 3.66007f
C24 VDD1.n3 B 0.710024f
C25 VDD1.t5 B 0.402785f
C26 VDD1.t1 B 0.402785f
C27 VDD1.n4 B 3.66216f
C28 VDD1.n5 B 2.47625f
C29 VDD1.t7 B 0.402785f
C30 VDD1.t8 B 0.402785f
C31 VDD1.n6 B 3.66006f
C32 VDD1.n7 B 3.1249f
C33 VP.n0 B 0.05442f
C34 VP.t4 B 0.813811f
C35 VP.t5 B 0.813811f
C36 VP.n1 B 0.02275f
C37 VP.n2 B 0.05442f
C38 VP.t2 B 0.813811f
C39 VP.t9 B 0.813811f
C40 VP.n3 B 0.02275f
C41 VP.t7 B 0.822421f
C42 VP.t0 B 0.813811f
C43 VP.n4 B 0.307063f
C44 VP.n5 B 0.324301f
C45 VP.n6 B 0.121175f
C46 VP.n7 B 0.05442f
C47 VP.n8 B 0.325115f
C48 VP.n9 B 0.02275f
C49 VP.n10 B 0.307063f
C50 VP.t1 B 0.822421f
C51 VP.n11 B 0.324223f
C52 VP.n12 B 2.47852f
C53 VP.t3 B 0.822421f
C54 VP.t6 B 0.813811f
C55 VP.n13 B 0.307063f
C56 VP.n14 B 0.324223f
C57 VP.n15 B 2.52238f
C58 VP.n16 B 0.05442f
C59 VP.n17 B 0.05442f
C60 VP.n18 B 0.325115f
C61 VP.n19 B 0.02275f
C62 VP.n20 B 0.307063f
C63 VP.t8 B 0.822421f
C64 VP.n21 B 0.324223f
C65 VP.n22 B 0.042173f
C66 VTAIL.t15 B 0.409582f
C67 VTAIL.t19 B 0.409582f
C68 VTAIL.n0 B 3.62626f
C69 VTAIL.n1 B 0.42574f
C70 VTAIL.t0 B 4.62985f
C71 VTAIL.n2 B 0.546972f
C72 VTAIL.t5 B 0.409582f
C73 VTAIL.t4 B 0.409582f
C74 VTAIL.n3 B 3.62626f
C75 VTAIL.n4 B 0.41459f
C76 VTAIL.t1 B 0.409582f
C77 VTAIL.t8 B 0.409582f
C78 VTAIL.n5 B 3.62626f
C79 VTAIL.n6 B 2.31968f
C80 VTAIL.t16 B 0.409582f
C81 VTAIL.t13 B 0.409582f
C82 VTAIL.n7 B 3.62626f
C83 VTAIL.n8 B 2.31967f
C84 VTAIL.t12 B 0.409582f
C85 VTAIL.t17 B 0.409582f
C86 VTAIL.n9 B 3.62626f
C87 VTAIL.n10 B 0.414585f
C88 VTAIL.t14 B 4.62988f
C89 VTAIL.n11 B 0.546943f
C90 VTAIL.t7 B 0.409582f
C91 VTAIL.t3 B 0.409582f
C92 VTAIL.n12 B 3.62626f
C93 VTAIL.n13 B 0.433518f
C94 VTAIL.t9 B 0.409582f
C95 VTAIL.t6 B 0.409582f
C96 VTAIL.n14 B 3.62626f
C97 VTAIL.n15 B 0.414585f
C98 VTAIL.t2 B 4.62985f
C99 VTAIL.n16 B 2.37927f
C100 VTAIL.t10 B 4.62985f
C101 VTAIL.n17 B 2.37927f
C102 VTAIL.t18 B 0.409582f
C103 VTAIL.t11 B 0.409582f
C104 VTAIL.n18 B 3.62626f
C105 VTAIL.n19 B 0.36852f
C106 VDD2.t5 B 4.66702f
C107 VDD2.t9 B 0.401725f
C108 VDD2.t8 B 0.401725f
C109 VDD2.n0 B 3.65044f
C110 VDD2.n1 B 0.708156f
C111 VDD2.t3 B 0.401725f
C112 VDD2.t2 B 0.401725f
C113 VDD2.n2 B 3.65252f
C114 VDD2.n3 B 2.38794f
C115 VDD2.t6 B 4.6635f
C116 VDD2.n4 B 3.13723f
C117 VDD2.t1 B 0.401725f
C118 VDD2.t0 B 0.401725f
C119 VDD2.n5 B 3.65044f
C120 VDD2.n6 B 0.31923f
C121 VDD2.t7 B 0.401725f
C122 VDD2.t4 B 0.401725f
C123 VDD2.n7 B 3.65248f
C124 VN.n0 B 0.053213f
C125 VN.t8 B 0.795763f
C126 VN.t1 B 0.795763f
C127 VN.n1 B 0.022246f
C128 VN.t4 B 0.804181f
C129 VN.t0 B 0.795763f
C130 VN.n2 B 0.300253f
C131 VN.n3 B 0.317109f
C132 VN.n4 B 0.118488f
C133 VN.n5 B 0.053213f
C134 VN.n6 B 0.317905f
C135 VN.n7 B 0.022246f
C136 VN.n8 B 0.300253f
C137 VN.t9 B 0.804181f
C138 VN.n9 B 0.317032f
C139 VN.n10 B 0.041238f
C140 VN.n11 B 0.053213f
C141 VN.t3 B 0.804181f
C142 VN.t6 B 0.795763f
C143 VN.t7 B 0.795763f
C144 VN.n12 B 0.022246f
C145 VN.t2 B 0.795763f
C146 VN.n13 B 0.300253f
C147 VN.t5 B 0.804181f
C148 VN.n14 B 0.317109f
C149 VN.n15 B 0.118488f
C150 VN.n16 B 0.053213f
C151 VN.n17 B 0.317905f
C152 VN.n18 B 0.022246f
C153 VN.n19 B 0.300253f
C154 VN.n20 B 0.317032f
C155 VN.n21 B 2.45836f
.ends

