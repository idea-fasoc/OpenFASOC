* NGSPICE file created from diff_pair_sample_1158.ext - technology: sky130A

.subckt diff_pair_sample_1158 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
X1 VTAIL.t0 VP.t0 VDD1.t7 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=1.65165 ps=10.34 w=10.01 l=2.42
X2 VDD1.t6 VP.t1 VTAIL.t1 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
X3 B.t11 B.t9 B.t10 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=0 ps=0 w=10.01 l=2.42
X4 VDD2.t6 VN.t1 VTAIL.t10 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
X5 B.t8 B.t6 B.t7 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=0 ps=0 w=10.01 l=2.42
X6 B.t5 B.t3 B.t4 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=0 ps=0 w=10.01 l=2.42
X7 VDD1.t5 VP.t2 VTAIL.t2 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
X8 B.t2 B.t0 B.t1 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=0 ps=0 w=10.01 l=2.42
X9 VDD2.t5 VN.t2 VTAIL.t13 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=3.9039 ps=20.8 w=10.01 l=2.42
X10 VTAIL.t12 VN.t3 VDD2.t4 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=1.65165 ps=10.34 w=10.01 l=2.42
X11 VDD1.t4 VP.t3 VTAIL.t3 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=3.9039 ps=20.8 w=10.01 l=2.42
X12 VDD1.t3 VP.t4 VTAIL.t5 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=3.9039 ps=20.8 w=10.01 l=2.42
X13 VTAIL.t15 VN.t4 VDD2.t3 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
X14 VTAIL.t11 VN.t5 VDD2.t2 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
X15 VTAIL.t6 VP.t5 VDD1.t2 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
X16 VTAIL.t9 VN.t6 VDD2.t1 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=1.65165 ps=10.34 w=10.01 l=2.42
X17 VTAIL.t4 VP.t6 VDD1.t1 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=3.9039 pd=20.8 as=1.65165 ps=10.34 w=10.01 l=2.42
X18 VDD2.t0 VN.t7 VTAIL.t14 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=3.9039 ps=20.8 w=10.01 l=2.42
X19 VTAIL.t7 VP.t7 VDD1.t0 w_n3720_n2970# sky130_fd_pr__pfet_01v8 ad=1.65165 pd=10.34 as=1.65165 ps=10.34 w=10.01 l=2.42
R0 VN.n51 VN.n27 161.3
R1 VN.n50 VN.n49 161.3
R2 VN.n48 VN.n28 161.3
R3 VN.n47 VN.n46 161.3
R4 VN.n45 VN.n29 161.3
R5 VN.n44 VN.n43 161.3
R6 VN.n42 VN.n41 161.3
R7 VN.n40 VN.n31 161.3
R8 VN.n39 VN.n38 161.3
R9 VN.n37 VN.n32 161.3
R10 VN.n36 VN.n35 161.3
R11 VN.n24 VN.n0 161.3
R12 VN.n23 VN.n22 161.3
R13 VN.n21 VN.n1 161.3
R14 VN.n20 VN.n19 161.3
R15 VN.n18 VN.n2 161.3
R16 VN.n17 VN.n16 161.3
R17 VN.n15 VN.n14 161.3
R18 VN.n13 VN.n4 161.3
R19 VN.n12 VN.n11 161.3
R20 VN.n10 VN.n5 161.3
R21 VN.n9 VN.n8 161.3
R22 VN.n6 VN.t6 132.111
R23 VN.n33 VN.t2 132.111
R24 VN.n26 VN.n25 104.639
R25 VN.n53 VN.n52 104.639
R26 VN.n7 VN.t0 99.6869
R27 VN.n3 VN.t5 99.6869
R28 VN.n25 VN.t7 99.6869
R29 VN.n34 VN.t4 99.6869
R30 VN.n30 VN.t1 99.6869
R31 VN.n52 VN.t3 99.6869
R32 VN.n19 VN.n1 56.5193
R33 VN.n46 VN.n28 56.5193
R34 VN.n7 VN.n6 53.8585
R35 VN.n34 VN.n33 53.8585
R36 VN VN.n53 48.7406
R37 VN.n12 VN.n5 40.4934
R38 VN.n13 VN.n12 40.4934
R39 VN.n39 VN.n32 40.4934
R40 VN.n40 VN.n39 40.4934
R41 VN.n8 VN.n5 24.4675
R42 VN.n14 VN.n13 24.4675
R43 VN.n18 VN.n17 24.4675
R44 VN.n19 VN.n18 24.4675
R45 VN.n23 VN.n1 24.4675
R46 VN.n24 VN.n23 24.4675
R47 VN.n35 VN.n32 24.4675
R48 VN.n46 VN.n45 24.4675
R49 VN.n45 VN.n44 24.4675
R50 VN.n41 VN.n40 24.4675
R51 VN.n51 VN.n50 24.4675
R52 VN.n50 VN.n28 24.4675
R53 VN.n8 VN.n7 18.3508
R54 VN.n14 VN.n3 18.3508
R55 VN.n35 VN.n34 18.3508
R56 VN.n41 VN.n30 18.3508
R57 VN.n36 VN.n33 7.09421
R58 VN.n9 VN.n6 7.09421
R59 VN.n17 VN.n3 6.11725
R60 VN.n25 VN.n24 6.11725
R61 VN.n44 VN.n30 6.11725
R62 VN.n52 VN.n51 6.11725
R63 VN.n53 VN.n27 0.278367
R64 VN.n26 VN.n0 0.278367
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n43 VN.n29 0.189894
R70 VN.n43 VN.n42 0.189894
R71 VN.n42 VN.n31 0.189894
R72 VN.n38 VN.n31 0.189894
R73 VN.n38 VN.n37 0.189894
R74 VN.n37 VN.n36 0.189894
R75 VN.n10 VN.n9 0.189894
R76 VN.n11 VN.n10 0.189894
R77 VN.n11 VN.n4 0.189894
R78 VN.n15 VN.n4 0.189894
R79 VN.n16 VN.n15 0.189894
R80 VN.n16 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153454
R86 VTAIL.n434 VTAIL.n386 756.745
R87 VTAIL.n50 VTAIL.n2 756.745
R88 VTAIL.n104 VTAIL.n56 756.745
R89 VTAIL.n160 VTAIL.n112 756.745
R90 VTAIL.n380 VTAIL.n332 756.745
R91 VTAIL.n324 VTAIL.n276 756.745
R92 VTAIL.n270 VTAIL.n222 756.745
R93 VTAIL.n214 VTAIL.n166 756.745
R94 VTAIL.n402 VTAIL.n401 585
R95 VTAIL.n407 VTAIL.n406 585
R96 VTAIL.n409 VTAIL.n408 585
R97 VTAIL.n398 VTAIL.n397 585
R98 VTAIL.n415 VTAIL.n414 585
R99 VTAIL.n417 VTAIL.n416 585
R100 VTAIL.n394 VTAIL.n393 585
R101 VTAIL.n424 VTAIL.n423 585
R102 VTAIL.n425 VTAIL.n392 585
R103 VTAIL.n427 VTAIL.n426 585
R104 VTAIL.n390 VTAIL.n389 585
R105 VTAIL.n433 VTAIL.n432 585
R106 VTAIL.n435 VTAIL.n434 585
R107 VTAIL.n18 VTAIL.n17 585
R108 VTAIL.n23 VTAIL.n22 585
R109 VTAIL.n25 VTAIL.n24 585
R110 VTAIL.n14 VTAIL.n13 585
R111 VTAIL.n31 VTAIL.n30 585
R112 VTAIL.n33 VTAIL.n32 585
R113 VTAIL.n10 VTAIL.n9 585
R114 VTAIL.n40 VTAIL.n39 585
R115 VTAIL.n41 VTAIL.n8 585
R116 VTAIL.n43 VTAIL.n42 585
R117 VTAIL.n6 VTAIL.n5 585
R118 VTAIL.n49 VTAIL.n48 585
R119 VTAIL.n51 VTAIL.n50 585
R120 VTAIL.n72 VTAIL.n71 585
R121 VTAIL.n77 VTAIL.n76 585
R122 VTAIL.n79 VTAIL.n78 585
R123 VTAIL.n68 VTAIL.n67 585
R124 VTAIL.n85 VTAIL.n84 585
R125 VTAIL.n87 VTAIL.n86 585
R126 VTAIL.n64 VTAIL.n63 585
R127 VTAIL.n94 VTAIL.n93 585
R128 VTAIL.n95 VTAIL.n62 585
R129 VTAIL.n97 VTAIL.n96 585
R130 VTAIL.n60 VTAIL.n59 585
R131 VTAIL.n103 VTAIL.n102 585
R132 VTAIL.n105 VTAIL.n104 585
R133 VTAIL.n128 VTAIL.n127 585
R134 VTAIL.n133 VTAIL.n132 585
R135 VTAIL.n135 VTAIL.n134 585
R136 VTAIL.n124 VTAIL.n123 585
R137 VTAIL.n141 VTAIL.n140 585
R138 VTAIL.n143 VTAIL.n142 585
R139 VTAIL.n120 VTAIL.n119 585
R140 VTAIL.n150 VTAIL.n149 585
R141 VTAIL.n151 VTAIL.n118 585
R142 VTAIL.n153 VTAIL.n152 585
R143 VTAIL.n116 VTAIL.n115 585
R144 VTAIL.n159 VTAIL.n158 585
R145 VTAIL.n161 VTAIL.n160 585
R146 VTAIL.n381 VTAIL.n380 585
R147 VTAIL.n379 VTAIL.n378 585
R148 VTAIL.n336 VTAIL.n335 585
R149 VTAIL.n373 VTAIL.n372 585
R150 VTAIL.n371 VTAIL.n338 585
R151 VTAIL.n370 VTAIL.n369 585
R152 VTAIL.n341 VTAIL.n339 585
R153 VTAIL.n364 VTAIL.n363 585
R154 VTAIL.n362 VTAIL.n361 585
R155 VTAIL.n345 VTAIL.n344 585
R156 VTAIL.n356 VTAIL.n355 585
R157 VTAIL.n354 VTAIL.n353 585
R158 VTAIL.n349 VTAIL.n348 585
R159 VTAIL.n325 VTAIL.n324 585
R160 VTAIL.n323 VTAIL.n322 585
R161 VTAIL.n280 VTAIL.n279 585
R162 VTAIL.n317 VTAIL.n316 585
R163 VTAIL.n315 VTAIL.n282 585
R164 VTAIL.n314 VTAIL.n313 585
R165 VTAIL.n285 VTAIL.n283 585
R166 VTAIL.n308 VTAIL.n307 585
R167 VTAIL.n306 VTAIL.n305 585
R168 VTAIL.n289 VTAIL.n288 585
R169 VTAIL.n300 VTAIL.n299 585
R170 VTAIL.n298 VTAIL.n297 585
R171 VTAIL.n293 VTAIL.n292 585
R172 VTAIL.n271 VTAIL.n270 585
R173 VTAIL.n269 VTAIL.n268 585
R174 VTAIL.n226 VTAIL.n225 585
R175 VTAIL.n263 VTAIL.n262 585
R176 VTAIL.n261 VTAIL.n228 585
R177 VTAIL.n260 VTAIL.n259 585
R178 VTAIL.n231 VTAIL.n229 585
R179 VTAIL.n254 VTAIL.n253 585
R180 VTAIL.n252 VTAIL.n251 585
R181 VTAIL.n235 VTAIL.n234 585
R182 VTAIL.n246 VTAIL.n245 585
R183 VTAIL.n244 VTAIL.n243 585
R184 VTAIL.n239 VTAIL.n238 585
R185 VTAIL.n215 VTAIL.n214 585
R186 VTAIL.n213 VTAIL.n212 585
R187 VTAIL.n170 VTAIL.n169 585
R188 VTAIL.n207 VTAIL.n206 585
R189 VTAIL.n205 VTAIL.n172 585
R190 VTAIL.n204 VTAIL.n203 585
R191 VTAIL.n175 VTAIL.n173 585
R192 VTAIL.n198 VTAIL.n197 585
R193 VTAIL.n196 VTAIL.n195 585
R194 VTAIL.n179 VTAIL.n178 585
R195 VTAIL.n190 VTAIL.n189 585
R196 VTAIL.n188 VTAIL.n187 585
R197 VTAIL.n183 VTAIL.n182 585
R198 VTAIL.n403 VTAIL.t14 329.038
R199 VTAIL.n19 VTAIL.t9 329.038
R200 VTAIL.n73 VTAIL.t3 329.038
R201 VTAIL.n129 VTAIL.t4 329.038
R202 VTAIL.n350 VTAIL.t5 329.038
R203 VTAIL.n294 VTAIL.t0 329.038
R204 VTAIL.n240 VTAIL.t13 329.038
R205 VTAIL.n184 VTAIL.t12 329.038
R206 VTAIL.n407 VTAIL.n401 171.744
R207 VTAIL.n408 VTAIL.n407 171.744
R208 VTAIL.n408 VTAIL.n397 171.744
R209 VTAIL.n415 VTAIL.n397 171.744
R210 VTAIL.n416 VTAIL.n415 171.744
R211 VTAIL.n416 VTAIL.n393 171.744
R212 VTAIL.n424 VTAIL.n393 171.744
R213 VTAIL.n425 VTAIL.n424 171.744
R214 VTAIL.n426 VTAIL.n425 171.744
R215 VTAIL.n426 VTAIL.n389 171.744
R216 VTAIL.n433 VTAIL.n389 171.744
R217 VTAIL.n434 VTAIL.n433 171.744
R218 VTAIL.n23 VTAIL.n17 171.744
R219 VTAIL.n24 VTAIL.n23 171.744
R220 VTAIL.n24 VTAIL.n13 171.744
R221 VTAIL.n31 VTAIL.n13 171.744
R222 VTAIL.n32 VTAIL.n31 171.744
R223 VTAIL.n32 VTAIL.n9 171.744
R224 VTAIL.n40 VTAIL.n9 171.744
R225 VTAIL.n41 VTAIL.n40 171.744
R226 VTAIL.n42 VTAIL.n41 171.744
R227 VTAIL.n42 VTAIL.n5 171.744
R228 VTAIL.n49 VTAIL.n5 171.744
R229 VTAIL.n50 VTAIL.n49 171.744
R230 VTAIL.n77 VTAIL.n71 171.744
R231 VTAIL.n78 VTAIL.n77 171.744
R232 VTAIL.n78 VTAIL.n67 171.744
R233 VTAIL.n85 VTAIL.n67 171.744
R234 VTAIL.n86 VTAIL.n85 171.744
R235 VTAIL.n86 VTAIL.n63 171.744
R236 VTAIL.n94 VTAIL.n63 171.744
R237 VTAIL.n95 VTAIL.n94 171.744
R238 VTAIL.n96 VTAIL.n95 171.744
R239 VTAIL.n96 VTAIL.n59 171.744
R240 VTAIL.n103 VTAIL.n59 171.744
R241 VTAIL.n104 VTAIL.n103 171.744
R242 VTAIL.n133 VTAIL.n127 171.744
R243 VTAIL.n134 VTAIL.n133 171.744
R244 VTAIL.n134 VTAIL.n123 171.744
R245 VTAIL.n141 VTAIL.n123 171.744
R246 VTAIL.n142 VTAIL.n141 171.744
R247 VTAIL.n142 VTAIL.n119 171.744
R248 VTAIL.n150 VTAIL.n119 171.744
R249 VTAIL.n151 VTAIL.n150 171.744
R250 VTAIL.n152 VTAIL.n151 171.744
R251 VTAIL.n152 VTAIL.n115 171.744
R252 VTAIL.n159 VTAIL.n115 171.744
R253 VTAIL.n160 VTAIL.n159 171.744
R254 VTAIL.n380 VTAIL.n379 171.744
R255 VTAIL.n379 VTAIL.n335 171.744
R256 VTAIL.n372 VTAIL.n335 171.744
R257 VTAIL.n372 VTAIL.n371 171.744
R258 VTAIL.n371 VTAIL.n370 171.744
R259 VTAIL.n370 VTAIL.n339 171.744
R260 VTAIL.n363 VTAIL.n339 171.744
R261 VTAIL.n363 VTAIL.n362 171.744
R262 VTAIL.n362 VTAIL.n344 171.744
R263 VTAIL.n355 VTAIL.n344 171.744
R264 VTAIL.n355 VTAIL.n354 171.744
R265 VTAIL.n354 VTAIL.n348 171.744
R266 VTAIL.n324 VTAIL.n323 171.744
R267 VTAIL.n323 VTAIL.n279 171.744
R268 VTAIL.n316 VTAIL.n279 171.744
R269 VTAIL.n316 VTAIL.n315 171.744
R270 VTAIL.n315 VTAIL.n314 171.744
R271 VTAIL.n314 VTAIL.n283 171.744
R272 VTAIL.n307 VTAIL.n283 171.744
R273 VTAIL.n307 VTAIL.n306 171.744
R274 VTAIL.n306 VTAIL.n288 171.744
R275 VTAIL.n299 VTAIL.n288 171.744
R276 VTAIL.n299 VTAIL.n298 171.744
R277 VTAIL.n298 VTAIL.n292 171.744
R278 VTAIL.n270 VTAIL.n269 171.744
R279 VTAIL.n269 VTAIL.n225 171.744
R280 VTAIL.n262 VTAIL.n225 171.744
R281 VTAIL.n262 VTAIL.n261 171.744
R282 VTAIL.n261 VTAIL.n260 171.744
R283 VTAIL.n260 VTAIL.n229 171.744
R284 VTAIL.n253 VTAIL.n229 171.744
R285 VTAIL.n253 VTAIL.n252 171.744
R286 VTAIL.n252 VTAIL.n234 171.744
R287 VTAIL.n245 VTAIL.n234 171.744
R288 VTAIL.n245 VTAIL.n244 171.744
R289 VTAIL.n244 VTAIL.n238 171.744
R290 VTAIL.n214 VTAIL.n213 171.744
R291 VTAIL.n213 VTAIL.n169 171.744
R292 VTAIL.n206 VTAIL.n169 171.744
R293 VTAIL.n206 VTAIL.n205 171.744
R294 VTAIL.n205 VTAIL.n204 171.744
R295 VTAIL.n204 VTAIL.n173 171.744
R296 VTAIL.n197 VTAIL.n173 171.744
R297 VTAIL.n197 VTAIL.n196 171.744
R298 VTAIL.n196 VTAIL.n178 171.744
R299 VTAIL.n189 VTAIL.n178 171.744
R300 VTAIL.n189 VTAIL.n188 171.744
R301 VTAIL.n188 VTAIL.n182 171.744
R302 VTAIL.t14 VTAIL.n401 85.8723
R303 VTAIL.t9 VTAIL.n17 85.8723
R304 VTAIL.t3 VTAIL.n71 85.8723
R305 VTAIL.t4 VTAIL.n127 85.8723
R306 VTAIL.t5 VTAIL.n348 85.8723
R307 VTAIL.t0 VTAIL.n292 85.8723
R308 VTAIL.t13 VTAIL.n238 85.8723
R309 VTAIL.t12 VTAIL.n182 85.8723
R310 VTAIL.n331 VTAIL.n330 61.4099
R311 VTAIL.n221 VTAIL.n220 61.4099
R312 VTAIL.n1 VTAIL.n0 61.4097
R313 VTAIL.n111 VTAIL.n110 61.4097
R314 VTAIL.n439 VTAIL.n438 33.155
R315 VTAIL.n55 VTAIL.n54 33.155
R316 VTAIL.n109 VTAIL.n108 33.155
R317 VTAIL.n165 VTAIL.n164 33.155
R318 VTAIL.n385 VTAIL.n384 33.155
R319 VTAIL.n329 VTAIL.n328 33.155
R320 VTAIL.n275 VTAIL.n274 33.155
R321 VTAIL.n219 VTAIL.n218 33.155
R322 VTAIL.n439 VTAIL.n385 23.3669
R323 VTAIL.n219 VTAIL.n165 23.3669
R324 VTAIL.n427 VTAIL.n392 13.1884
R325 VTAIL.n43 VTAIL.n8 13.1884
R326 VTAIL.n97 VTAIL.n62 13.1884
R327 VTAIL.n153 VTAIL.n118 13.1884
R328 VTAIL.n373 VTAIL.n338 13.1884
R329 VTAIL.n317 VTAIL.n282 13.1884
R330 VTAIL.n263 VTAIL.n228 13.1884
R331 VTAIL.n207 VTAIL.n172 13.1884
R332 VTAIL.n423 VTAIL.n422 12.8005
R333 VTAIL.n428 VTAIL.n390 12.8005
R334 VTAIL.n39 VTAIL.n38 12.8005
R335 VTAIL.n44 VTAIL.n6 12.8005
R336 VTAIL.n93 VTAIL.n92 12.8005
R337 VTAIL.n98 VTAIL.n60 12.8005
R338 VTAIL.n149 VTAIL.n148 12.8005
R339 VTAIL.n154 VTAIL.n116 12.8005
R340 VTAIL.n374 VTAIL.n336 12.8005
R341 VTAIL.n369 VTAIL.n340 12.8005
R342 VTAIL.n318 VTAIL.n280 12.8005
R343 VTAIL.n313 VTAIL.n284 12.8005
R344 VTAIL.n264 VTAIL.n226 12.8005
R345 VTAIL.n259 VTAIL.n230 12.8005
R346 VTAIL.n208 VTAIL.n170 12.8005
R347 VTAIL.n203 VTAIL.n174 12.8005
R348 VTAIL.n421 VTAIL.n394 12.0247
R349 VTAIL.n432 VTAIL.n431 12.0247
R350 VTAIL.n37 VTAIL.n10 12.0247
R351 VTAIL.n48 VTAIL.n47 12.0247
R352 VTAIL.n91 VTAIL.n64 12.0247
R353 VTAIL.n102 VTAIL.n101 12.0247
R354 VTAIL.n147 VTAIL.n120 12.0247
R355 VTAIL.n158 VTAIL.n157 12.0247
R356 VTAIL.n378 VTAIL.n377 12.0247
R357 VTAIL.n368 VTAIL.n341 12.0247
R358 VTAIL.n322 VTAIL.n321 12.0247
R359 VTAIL.n312 VTAIL.n285 12.0247
R360 VTAIL.n268 VTAIL.n267 12.0247
R361 VTAIL.n258 VTAIL.n231 12.0247
R362 VTAIL.n212 VTAIL.n211 12.0247
R363 VTAIL.n202 VTAIL.n175 12.0247
R364 VTAIL.n418 VTAIL.n417 11.249
R365 VTAIL.n435 VTAIL.n388 11.249
R366 VTAIL.n34 VTAIL.n33 11.249
R367 VTAIL.n51 VTAIL.n4 11.249
R368 VTAIL.n88 VTAIL.n87 11.249
R369 VTAIL.n105 VTAIL.n58 11.249
R370 VTAIL.n144 VTAIL.n143 11.249
R371 VTAIL.n161 VTAIL.n114 11.249
R372 VTAIL.n381 VTAIL.n334 11.249
R373 VTAIL.n365 VTAIL.n364 11.249
R374 VTAIL.n325 VTAIL.n278 11.249
R375 VTAIL.n309 VTAIL.n308 11.249
R376 VTAIL.n271 VTAIL.n224 11.249
R377 VTAIL.n255 VTAIL.n254 11.249
R378 VTAIL.n215 VTAIL.n168 11.249
R379 VTAIL.n199 VTAIL.n198 11.249
R380 VTAIL.n403 VTAIL.n402 10.7239
R381 VTAIL.n19 VTAIL.n18 10.7239
R382 VTAIL.n73 VTAIL.n72 10.7239
R383 VTAIL.n129 VTAIL.n128 10.7239
R384 VTAIL.n350 VTAIL.n349 10.7239
R385 VTAIL.n294 VTAIL.n293 10.7239
R386 VTAIL.n240 VTAIL.n239 10.7239
R387 VTAIL.n184 VTAIL.n183 10.7239
R388 VTAIL.n414 VTAIL.n396 10.4732
R389 VTAIL.n436 VTAIL.n386 10.4732
R390 VTAIL.n30 VTAIL.n12 10.4732
R391 VTAIL.n52 VTAIL.n2 10.4732
R392 VTAIL.n84 VTAIL.n66 10.4732
R393 VTAIL.n106 VTAIL.n56 10.4732
R394 VTAIL.n140 VTAIL.n122 10.4732
R395 VTAIL.n162 VTAIL.n112 10.4732
R396 VTAIL.n382 VTAIL.n332 10.4732
R397 VTAIL.n361 VTAIL.n343 10.4732
R398 VTAIL.n326 VTAIL.n276 10.4732
R399 VTAIL.n305 VTAIL.n287 10.4732
R400 VTAIL.n272 VTAIL.n222 10.4732
R401 VTAIL.n251 VTAIL.n233 10.4732
R402 VTAIL.n216 VTAIL.n166 10.4732
R403 VTAIL.n195 VTAIL.n177 10.4732
R404 VTAIL.n413 VTAIL.n398 9.69747
R405 VTAIL.n29 VTAIL.n14 9.69747
R406 VTAIL.n83 VTAIL.n68 9.69747
R407 VTAIL.n139 VTAIL.n124 9.69747
R408 VTAIL.n360 VTAIL.n345 9.69747
R409 VTAIL.n304 VTAIL.n289 9.69747
R410 VTAIL.n250 VTAIL.n235 9.69747
R411 VTAIL.n194 VTAIL.n179 9.69747
R412 VTAIL.n438 VTAIL.n437 9.45567
R413 VTAIL.n54 VTAIL.n53 9.45567
R414 VTAIL.n108 VTAIL.n107 9.45567
R415 VTAIL.n164 VTAIL.n163 9.45567
R416 VTAIL.n384 VTAIL.n383 9.45567
R417 VTAIL.n328 VTAIL.n327 9.45567
R418 VTAIL.n274 VTAIL.n273 9.45567
R419 VTAIL.n218 VTAIL.n217 9.45567
R420 VTAIL.n437 VTAIL.n436 9.3005
R421 VTAIL.n388 VTAIL.n387 9.3005
R422 VTAIL.n431 VTAIL.n430 9.3005
R423 VTAIL.n429 VTAIL.n428 9.3005
R424 VTAIL.n405 VTAIL.n404 9.3005
R425 VTAIL.n400 VTAIL.n399 9.3005
R426 VTAIL.n411 VTAIL.n410 9.3005
R427 VTAIL.n413 VTAIL.n412 9.3005
R428 VTAIL.n396 VTAIL.n395 9.3005
R429 VTAIL.n419 VTAIL.n418 9.3005
R430 VTAIL.n421 VTAIL.n420 9.3005
R431 VTAIL.n422 VTAIL.n391 9.3005
R432 VTAIL.n53 VTAIL.n52 9.3005
R433 VTAIL.n4 VTAIL.n3 9.3005
R434 VTAIL.n47 VTAIL.n46 9.3005
R435 VTAIL.n45 VTAIL.n44 9.3005
R436 VTAIL.n21 VTAIL.n20 9.3005
R437 VTAIL.n16 VTAIL.n15 9.3005
R438 VTAIL.n27 VTAIL.n26 9.3005
R439 VTAIL.n29 VTAIL.n28 9.3005
R440 VTAIL.n12 VTAIL.n11 9.3005
R441 VTAIL.n35 VTAIL.n34 9.3005
R442 VTAIL.n37 VTAIL.n36 9.3005
R443 VTAIL.n38 VTAIL.n7 9.3005
R444 VTAIL.n107 VTAIL.n106 9.3005
R445 VTAIL.n58 VTAIL.n57 9.3005
R446 VTAIL.n101 VTAIL.n100 9.3005
R447 VTAIL.n99 VTAIL.n98 9.3005
R448 VTAIL.n75 VTAIL.n74 9.3005
R449 VTAIL.n70 VTAIL.n69 9.3005
R450 VTAIL.n81 VTAIL.n80 9.3005
R451 VTAIL.n83 VTAIL.n82 9.3005
R452 VTAIL.n66 VTAIL.n65 9.3005
R453 VTAIL.n89 VTAIL.n88 9.3005
R454 VTAIL.n91 VTAIL.n90 9.3005
R455 VTAIL.n92 VTAIL.n61 9.3005
R456 VTAIL.n163 VTAIL.n162 9.3005
R457 VTAIL.n114 VTAIL.n113 9.3005
R458 VTAIL.n157 VTAIL.n156 9.3005
R459 VTAIL.n155 VTAIL.n154 9.3005
R460 VTAIL.n131 VTAIL.n130 9.3005
R461 VTAIL.n126 VTAIL.n125 9.3005
R462 VTAIL.n137 VTAIL.n136 9.3005
R463 VTAIL.n139 VTAIL.n138 9.3005
R464 VTAIL.n122 VTAIL.n121 9.3005
R465 VTAIL.n145 VTAIL.n144 9.3005
R466 VTAIL.n147 VTAIL.n146 9.3005
R467 VTAIL.n148 VTAIL.n117 9.3005
R468 VTAIL.n352 VTAIL.n351 9.3005
R469 VTAIL.n347 VTAIL.n346 9.3005
R470 VTAIL.n358 VTAIL.n357 9.3005
R471 VTAIL.n360 VTAIL.n359 9.3005
R472 VTAIL.n343 VTAIL.n342 9.3005
R473 VTAIL.n366 VTAIL.n365 9.3005
R474 VTAIL.n368 VTAIL.n367 9.3005
R475 VTAIL.n340 VTAIL.n337 9.3005
R476 VTAIL.n383 VTAIL.n382 9.3005
R477 VTAIL.n334 VTAIL.n333 9.3005
R478 VTAIL.n377 VTAIL.n376 9.3005
R479 VTAIL.n375 VTAIL.n374 9.3005
R480 VTAIL.n296 VTAIL.n295 9.3005
R481 VTAIL.n291 VTAIL.n290 9.3005
R482 VTAIL.n302 VTAIL.n301 9.3005
R483 VTAIL.n304 VTAIL.n303 9.3005
R484 VTAIL.n287 VTAIL.n286 9.3005
R485 VTAIL.n310 VTAIL.n309 9.3005
R486 VTAIL.n312 VTAIL.n311 9.3005
R487 VTAIL.n284 VTAIL.n281 9.3005
R488 VTAIL.n327 VTAIL.n326 9.3005
R489 VTAIL.n278 VTAIL.n277 9.3005
R490 VTAIL.n321 VTAIL.n320 9.3005
R491 VTAIL.n319 VTAIL.n318 9.3005
R492 VTAIL.n242 VTAIL.n241 9.3005
R493 VTAIL.n237 VTAIL.n236 9.3005
R494 VTAIL.n248 VTAIL.n247 9.3005
R495 VTAIL.n250 VTAIL.n249 9.3005
R496 VTAIL.n233 VTAIL.n232 9.3005
R497 VTAIL.n256 VTAIL.n255 9.3005
R498 VTAIL.n258 VTAIL.n257 9.3005
R499 VTAIL.n230 VTAIL.n227 9.3005
R500 VTAIL.n273 VTAIL.n272 9.3005
R501 VTAIL.n224 VTAIL.n223 9.3005
R502 VTAIL.n267 VTAIL.n266 9.3005
R503 VTAIL.n265 VTAIL.n264 9.3005
R504 VTAIL.n186 VTAIL.n185 9.3005
R505 VTAIL.n181 VTAIL.n180 9.3005
R506 VTAIL.n192 VTAIL.n191 9.3005
R507 VTAIL.n194 VTAIL.n193 9.3005
R508 VTAIL.n177 VTAIL.n176 9.3005
R509 VTAIL.n200 VTAIL.n199 9.3005
R510 VTAIL.n202 VTAIL.n201 9.3005
R511 VTAIL.n174 VTAIL.n171 9.3005
R512 VTAIL.n217 VTAIL.n216 9.3005
R513 VTAIL.n168 VTAIL.n167 9.3005
R514 VTAIL.n211 VTAIL.n210 9.3005
R515 VTAIL.n209 VTAIL.n208 9.3005
R516 VTAIL.n410 VTAIL.n409 8.92171
R517 VTAIL.n26 VTAIL.n25 8.92171
R518 VTAIL.n80 VTAIL.n79 8.92171
R519 VTAIL.n136 VTAIL.n135 8.92171
R520 VTAIL.n357 VTAIL.n356 8.92171
R521 VTAIL.n301 VTAIL.n300 8.92171
R522 VTAIL.n247 VTAIL.n246 8.92171
R523 VTAIL.n191 VTAIL.n190 8.92171
R524 VTAIL.n406 VTAIL.n400 8.14595
R525 VTAIL.n22 VTAIL.n16 8.14595
R526 VTAIL.n76 VTAIL.n70 8.14595
R527 VTAIL.n132 VTAIL.n126 8.14595
R528 VTAIL.n353 VTAIL.n347 8.14595
R529 VTAIL.n297 VTAIL.n291 8.14595
R530 VTAIL.n243 VTAIL.n237 8.14595
R531 VTAIL.n187 VTAIL.n181 8.14595
R532 VTAIL.n405 VTAIL.n402 7.3702
R533 VTAIL.n21 VTAIL.n18 7.3702
R534 VTAIL.n75 VTAIL.n72 7.3702
R535 VTAIL.n131 VTAIL.n128 7.3702
R536 VTAIL.n352 VTAIL.n349 7.3702
R537 VTAIL.n296 VTAIL.n293 7.3702
R538 VTAIL.n242 VTAIL.n239 7.3702
R539 VTAIL.n186 VTAIL.n183 7.3702
R540 VTAIL.n406 VTAIL.n405 5.81868
R541 VTAIL.n22 VTAIL.n21 5.81868
R542 VTAIL.n76 VTAIL.n75 5.81868
R543 VTAIL.n132 VTAIL.n131 5.81868
R544 VTAIL.n353 VTAIL.n352 5.81868
R545 VTAIL.n297 VTAIL.n296 5.81868
R546 VTAIL.n243 VTAIL.n242 5.81868
R547 VTAIL.n187 VTAIL.n186 5.81868
R548 VTAIL.n409 VTAIL.n400 5.04292
R549 VTAIL.n25 VTAIL.n16 5.04292
R550 VTAIL.n79 VTAIL.n70 5.04292
R551 VTAIL.n135 VTAIL.n126 5.04292
R552 VTAIL.n356 VTAIL.n347 5.04292
R553 VTAIL.n300 VTAIL.n291 5.04292
R554 VTAIL.n246 VTAIL.n237 5.04292
R555 VTAIL.n190 VTAIL.n181 5.04292
R556 VTAIL.n410 VTAIL.n398 4.26717
R557 VTAIL.n26 VTAIL.n14 4.26717
R558 VTAIL.n80 VTAIL.n68 4.26717
R559 VTAIL.n136 VTAIL.n124 4.26717
R560 VTAIL.n357 VTAIL.n345 4.26717
R561 VTAIL.n301 VTAIL.n289 4.26717
R562 VTAIL.n247 VTAIL.n235 4.26717
R563 VTAIL.n191 VTAIL.n179 4.26717
R564 VTAIL.n414 VTAIL.n413 3.49141
R565 VTAIL.n438 VTAIL.n386 3.49141
R566 VTAIL.n30 VTAIL.n29 3.49141
R567 VTAIL.n54 VTAIL.n2 3.49141
R568 VTAIL.n84 VTAIL.n83 3.49141
R569 VTAIL.n108 VTAIL.n56 3.49141
R570 VTAIL.n140 VTAIL.n139 3.49141
R571 VTAIL.n164 VTAIL.n112 3.49141
R572 VTAIL.n384 VTAIL.n332 3.49141
R573 VTAIL.n361 VTAIL.n360 3.49141
R574 VTAIL.n328 VTAIL.n276 3.49141
R575 VTAIL.n305 VTAIL.n304 3.49141
R576 VTAIL.n274 VTAIL.n222 3.49141
R577 VTAIL.n251 VTAIL.n250 3.49141
R578 VTAIL.n218 VTAIL.n166 3.49141
R579 VTAIL.n195 VTAIL.n194 3.49141
R580 VTAIL.n0 VTAIL.t8 3.24775
R581 VTAIL.n0 VTAIL.t11 3.24775
R582 VTAIL.n110 VTAIL.t2 3.24775
R583 VTAIL.n110 VTAIL.t7 3.24775
R584 VTAIL.n330 VTAIL.t1 3.24775
R585 VTAIL.n330 VTAIL.t6 3.24775
R586 VTAIL.n220 VTAIL.t10 3.24775
R587 VTAIL.n220 VTAIL.t15 3.24775
R588 VTAIL.n417 VTAIL.n396 2.71565
R589 VTAIL.n436 VTAIL.n435 2.71565
R590 VTAIL.n33 VTAIL.n12 2.71565
R591 VTAIL.n52 VTAIL.n51 2.71565
R592 VTAIL.n87 VTAIL.n66 2.71565
R593 VTAIL.n106 VTAIL.n105 2.71565
R594 VTAIL.n143 VTAIL.n122 2.71565
R595 VTAIL.n162 VTAIL.n161 2.71565
R596 VTAIL.n382 VTAIL.n381 2.71565
R597 VTAIL.n364 VTAIL.n343 2.71565
R598 VTAIL.n326 VTAIL.n325 2.71565
R599 VTAIL.n308 VTAIL.n287 2.71565
R600 VTAIL.n272 VTAIL.n271 2.71565
R601 VTAIL.n254 VTAIL.n233 2.71565
R602 VTAIL.n216 VTAIL.n215 2.71565
R603 VTAIL.n198 VTAIL.n177 2.71565
R604 VTAIL.n404 VTAIL.n403 2.41283
R605 VTAIL.n20 VTAIL.n19 2.41283
R606 VTAIL.n74 VTAIL.n73 2.41283
R607 VTAIL.n130 VTAIL.n129 2.41283
R608 VTAIL.n351 VTAIL.n350 2.41283
R609 VTAIL.n295 VTAIL.n294 2.41283
R610 VTAIL.n241 VTAIL.n240 2.41283
R611 VTAIL.n185 VTAIL.n184 2.41283
R612 VTAIL.n221 VTAIL.n219 2.37119
R613 VTAIL.n275 VTAIL.n221 2.37119
R614 VTAIL.n331 VTAIL.n329 2.37119
R615 VTAIL.n385 VTAIL.n331 2.37119
R616 VTAIL.n165 VTAIL.n111 2.37119
R617 VTAIL.n111 VTAIL.n109 2.37119
R618 VTAIL.n55 VTAIL.n1 2.37119
R619 VTAIL VTAIL.n439 2.313
R620 VTAIL.n418 VTAIL.n394 1.93989
R621 VTAIL.n432 VTAIL.n388 1.93989
R622 VTAIL.n34 VTAIL.n10 1.93989
R623 VTAIL.n48 VTAIL.n4 1.93989
R624 VTAIL.n88 VTAIL.n64 1.93989
R625 VTAIL.n102 VTAIL.n58 1.93989
R626 VTAIL.n144 VTAIL.n120 1.93989
R627 VTAIL.n158 VTAIL.n114 1.93989
R628 VTAIL.n378 VTAIL.n334 1.93989
R629 VTAIL.n365 VTAIL.n341 1.93989
R630 VTAIL.n322 VTAIL.n278 1.93989
R631 VTAIL.n309 VTAIL.n285 1.93989
R632 VTAIL.n268 VTAIL.n224 1.93989
R633 VTAIL.n255 VTAIL.n231 1.93989
R634 VTAIL.n212 VTAIL.n168 1.93989
R635 VTAIL.n199 VTAIL.n175 1.93989
R636 VTAIL.n423 VTAIL.n421 1.16414
R637 VTAIL.n431 VTAIL.n390 1.16414
R638 VTAIL.n39 VTAIL.n37 1.16414
R639 VTAIL.n47 VTAIL.n6 1.16414
R640 VTAIL.n93 VTAIL.n91 1.16414
R641 VTAIL.n101 VTAIL.n60 1.16414
R642 VTAIL.n149 VTAIL.n147 1.16414
R643 VTAIL.n157 VTAIL.n116 1.16414
R644 VTAIL.n377 VTAIL.n336 1.16414
R645 VTAIL.n369 VTAIL.n368 1.16414
R646 VTAIL.n321 VTAIL.n280 1.16414
R647 VTAIL.n313 VTAIL.n312 1.16414
R648 VTAIL.n267 VTAIL.n226 1.16414
R649 VTAIL.n259 VTAIL.n258 1.16414
R650 VTAIL.n211 VTAIL.n170 1.16414
R651 VTAIL.n203 VTAIL.n202 1.16414
R652 VTAIL.n329 VTAIL.n275 0.470328
R653 VTAIL.n109 VTAIL.n55 0.470328
R654 VTAIL.n422 VTAIL.n392 0.388379
R655 VTAIL.n428 VTAIL.n427 0.388379
R656 VTAIL.n38 VTAIL.n8 0.388379
R657 VTAIL.n44 VTAIL.n43 0.388379
R658 VTAIL.n92 VTAIL.n62 0.388379
R659 VTAIL.n98 VTAIL.n97 0.388379
R660 VTAIL.n148 VTAIL.n118 0.388379
R661 VTAIL.n154 VTAIL.n153 0.388379
R662 VTAIL.n374 VTAIL.n373 0.388379
R663 VTAIL.n340 VTAIL.n338 0.388379
R664 VTAIL.n318 VTAIL.n317 0.388379
R665 VTAIL.n284 VTAIL.n282 0.388379
R666 VTAIL.n264 VTAIL.n263 0.388379
R667 VTAIL.n230 VTAIL.n228 0.388379
R668 VTAIL.n208 VTAIL.n207 0.388379
R669 VTAIL.n174 VTAIL.n172 0.388379
R670 VTAIL.n404 VTAIL.n399 0.155672
R671 VTAIL.n411 VTAIL.n399 0.155672
R672 VTAIL.n412 VTAIL.n411 0.155672
R673 VTAIL.n412 VTAIL.n395 0.155672
R674 VTAIL.n419 VTAIL.n395 0.155672
R675 VTAIL.n420 VTAIL.n419 0.155672
R676 VTAIL.n420 VTAIL.n391 0.155672
R677 VTAIL.n429 VTAIL.n391 0.155672
R678 VTAIL.n430 VTAIL.n429 0.155672
R679 VTAIL.n430 VTAIL.n387 0.155672
R680 VTAIL.n437 VTAIL.n387 0.155672
R681 VTAIL.n20 VTAIL.n15 0.155672
R682 VTAIL.n27 VTAIL.n15 0.155672
R683 VTAIL.n28 VTAIL.n27 0.155672
R684 VTAIL.n28 VTAIL.n11 0.155672
R685 VTAIL.n35 VTAIL.n11 0.155672
R686 VTAIL.n36 VTAIL.n35 0.155672
R687 VTAIL.n36 VTAIL.n7 0.155672
R688 VTAIL.n45 VTAIL.n7 0.155672
R689 VTAIL.n46 VTAIL.n45 0.155672
R690 VTAIL.n46 VTAIL.n3 0.155672
R691 VTAIL.n53 VTAIL.n3 0.155672
R692 VTAIL.n74 VTAIL.n69 0.155672
R693 VTAIL.n81 VTAIL.n69 0.155672
R694 VTAIL.n82 VTAIL.n81 0.155672
R695 VTAIL.n82 VTAIL.n65 0.155672
R696 VTAIL.n89 VTAIL.n65 0.155672
R697 VTAIL.n90 VTAIL.n89 0.155672
R698 VTAIL.n90 VTAIL.n61 0.155672
R699 VTAIL.n99 VTAIL.n61 0.155672
R700 VTAIL.n100 VTAIL.n99 0.155672
R701 VTAIL.n100 VTAIL.n57 0.155672
R702 VTAIL.n107 VTAIL.n57 0.155672
R703 VTAIL.n130 VTAIL.n125 0.155672
R704 VTAIL.n137 VTAIL.n125 0.155672
R705 VTAIL.n138 VTAIL.n137 0.155672
R706 VTAIL.n138 VTAIL.n121 0.155672
R707 VTAIL.n145 VTAIL.n121 0.155672
R708 VTAIL.n146 VTAIL.n145 0.155672
R709 VTAIL.n146 VTAIL.n117 0.155672
R710 VTAIL.n155 VTAIL.n117 0.155672
R711 VTAIL.n156 VTAIL.n155 0.155672
R712 VTAIL.n156 VTAIL.n113 0.155672
R713 VTAIL.n163 VTAIL.n113 0.155672
R714 VTAIL.n383 VTAIL.n333 0.155672
R715 VTAIL.n376 VTAIL.n333 0.155672
R716 VTAIL.n376 VTAIL.n375 0.155672
R717 VTAIL.n375 VTAIL.n337 0.155672
R718 VTAIL.n367 VTAIL.n337 0.155672
R719 VTAIL.n367 VTAIL.n366 0.155672
R720 VTAIL.n366 VTAIL.n342 0.155672
R721 VTAIL.n359 VTAIL.n342 0.155672
R722 VTAIL.n359 VTAIL.n358 0.155672
R723 VTAIL.n358 VTAIL.n346 0.155672
R724 VTAIL.n351 VTAIL.n346 0.155672
R725 VTAIL.n327 VTAIL.n277 0.155672
R726 VTAIL.n320 VTAIL.n277 0.155672
R727 VTAIL.n320 VTAIL.n319 0.155672
R728 VTAIL.n319 VTAIL.n281 0.155672
R729 VTAIL.n311 VTAIL.n281 0.155672
R730 VTAIL.n311 VTAIL.n310 0.155672
R731 VTAIL.n310 VTAIL.n286 0.155672
R732 VTAIL.n303 VTAIL.n286 0.155672
R733 VTAIL.n303 VTAIL.n302 0.155672
R734 VTAIL.n302 VTAIL.n290 0.155672
R735 VTAIL.n295 VTAIL.n290 0.155672
R736 VTAIL.n273 VTAIL.n223 0.155672
R737 VTAIL.n266 VTAIL.n223 0.155672
R738 VTAIL.n266 VTAIL.n265 0.155672
R739 VTAIL.n265 VTAIL.n227 0.155672
R740 VTAIL.n257 VTAIL.n227 0.155672
R741 VTAIL.n257 VTAIL.n256 0.155672
R742 VTAIL.n256 VTAIL.n232 0.155672
R743 VTAIL.n249 VTAIL.n232 0.155672
R744 VTAIL.n249 VTAIL.n248 0.155672
R745 VTAIL.n248 VTAIL.n236 0.155672
R746 VTAIL.n241 VTAIL.n236 0.155672
R747 VTAIL.n217 VTAIL.n167 0.155672
R748 VTAIL.n210 VTAIL.n167 0.155672
R749 VTAIL.n210 VTAIL.n209 0.155672
R750 VTAIL.n209 VTAIL.n171 0.155672
R751 VTAIL.n201 VTAIL.n171 0.155672
R752 VTAIL.n201 VTAIL.n200 0.155672
R753 VTAIL.n200 VTAIL.n176 0.155672
R754 VTAIL.n193 VTAIL.n176 0.155672
R755 VTAIL.n193 VTAIL.n192 0.155672
R756 VTAIL.n192 VTAIL.n180 0.155672
R757 VTAIL.n185 VTAIL.n180 0.155672
R758 VTAIL VTAIL.n1 0.0586897
R759 VDD2.n2 VDD2.n1 79.2185
R760 VDD2.n2 VDD2.n0 79.2185
R761 VDD2 VDD2.n5 79.2156
R762 VDD2.n4 VDD2.n3 78.0887
R763 VDD2.n4 VDD2.n2 43.0127
R764 VDD2.n5 VDD2.t3 3.24775
R765 VDD2.n5 VDD2.t5 3.24775
R766 VDD2.n3 VDD2.t4 3.24775
R767 VDD2.n3 VDD2.t6 3.24775
R768 VDD2.n1 VDD2.t2 3.24775
R769 VDD2.n1 VDD2.t0 3.24775
R770 VDD2.n0 VDD2.t1 3.24775
R771 VDD2.n0 VDD2.t7 3.24775
R772 VDD2 VDD2.n4 1.24403
R773 VP.n19 VP.n18 161.3
R774 VP.n20 VP.n15 161.3
R775 VP.n22 VP.n21 161.3
R776 VP.n23 VP.n14 161.3
R777 VP.n25 VP.n24 161.3
R778 VP.n27 VP.n26 161.3
R779 VP.n28 VP.n12 161.3
R780 VP.n30 VP.n29 161.3
R781 VP.n31 VP.n11 161.3
R782 VP.n33 VP.n32 161.3
R783 VP.n34 VP.n10 161.3
R784 VP.n64 VP.n0 161.3
R785 VP.n63 VP.n62 161.3
R786 VP.n61 VP.n1 161.3
R787 VP.n60 VP.n59 161.3
R788 VP.n58 VP.n2 161.3
R789 VP.n57 VP.n56 161.3
R790 VP.n55 VP.n54 161.3
R791 VP.n53 VP.n4 161.3
R792 VP.n52 VP.n51 161.3
R793 VP.n50 VP.n5 161.3
R794 VP.n49 VP.n48 161.3
R795 VP.n46 VP.n6 161.3
R796 VP.n45 VP.n44 161.3
R797 VP.n43 VP.n7 161.3
R798 VP.n42 VP.n41 161.3
R799 VP.n40 VP.n8 161.3
R800 VP.n39 VP.n38 161.3
R801 VP.n16 VP.t0 132.111
R802 VP.n37 VP.n9 104.639
R803 VP.n66 VP.n65 104.639
R804 VP.n36 VP.n35 104.639
R805 VP.n9 VP.t6 99.6869
R806 VP.n47 VP.t2 99.6869
R807 VP.n3 VP.t7 99.6869
R808 VP.n65 VP.t3 99.6869
R809 VP.n35 VP.t4 99.6869
R810 VP.n13 VP.t5 99.6869
R811 VP.n17 VP.t1 99.6869
R812 VP.n41 VP.n7 56.5193
R813 VP.n59 VP.n1 56.5193
R814 VP.n29 VP.n11 56.5193
R815 VP.n17 VP.n16 53.8585
R816 VP.n37 VP.n36 48.4617
R817 VP.n52 VP.n5 40.4934
R818 VP.n53 VP.n52 40.4934
R819 VP.n23 VP.n22 40.4934
R820 VP.n22 VP.n15 40.4934
R821 VP.n40 VP.n39 24.4675
R822 VP.n41 VP.n40 24.4675
R823 VP.n45 VP.n7 24.4675
R824 VP.n46 VP.n45 24.4675
R825 VP.n48 VP.n5 24.4675
R826 VP.n54 VP.n53 24.4675
R827 VP.n58 VP.n57 24.4675
R828 VP.n59 VP.n58 24.4675
R829 VP.n63 VP.n1 24.4675
R830 VP.n64 VP.n63 24.4675
R831 VP.n33 VP.n11 24.4675
R832 VP.n34 VP.n33 24.4675
R833 VP.n24 VP.n23 24.4675
R834 VP.n28 VP.n27 24.4675
R835 VP.n29 VP.n28 24.4675
R836 VP.n18 VP.n15 24.4675
R837 VP.n48 VP.n47 18.3508
R838 VP.n54 VP.n3 18.3508
R839 VP.n24 VP.n13 18.3508
R840 VP.n18 VP.n17 18.3508
R841 VP.n19 VP.n16 7.09421
R842 VP.n39 VP.n9 6.11725
R843 VP.n47 VP.n46 6.11725
R844 VP.n57 VP.n3 6.11725
R845 VP.n65 VP.n64 6.11725
R846 VP.n35 VP.n34 6.11725
R847 VP.n27 VP.n13 6.11725
R848 VP.n36 VP.n10 0.278367
R849 VP.n38 VP.n37 0.278367
R850 VP.n66 VP.n0 0.278367
R851 VP.n20 VP.n19 0.189894
R852 VP.n21 VP.n20 0.189894
R853 VP.n21 VP.n14 0.189894
R854 VP.n25 VP.n14 0.189894
R855 VP.n26 VP.n25 0.189894
R856 VP.n26 VP.n12 0.189894
R857 VP.n30 VP.n12 0.189894
R858 VP.n31 VP.n30 0.189894
R859 VP.n32 VP.n31 0.189894
R860 VP.n32 VP.n10 0.189894
R861 VP.n38 VP.n8 0.189894
R862 VP.n42 VP.n8 0.189894
R863 VP.n43 VP.n42 0.189894
R864 VP.n44 VP.n43 0.189894
R865 VP.n44 VP.n6 0.189894
R866 VP.n49 VP.n6 0.189894
R867 VP.n50 VP.n49 0.189894
R868 VP.n51 VP.n50 0.189894
R869 VP.n51 VP.n4 0.189894
R870 VP.n55 VP.n4 0.189894
R871 VP.n56 VP.n55 0.189894
R872 VP.n56 VP.n2 0.189894
R873 VP.n60 VP.n2 0.189894
R874 VP.n61 VP.n60 0.189894
R875 VP.n62 VP.n61 0.189894
R876 VP.n62 VP.n0 0.189894
R877 VP VP.n66 0.153454
R878 VDD1 VDD1.n0 79.3322
R879 VDD1.n3 VDD1.n2 79.2185
R880 VDD1.n3 VDD1.n1 79.2185
R881 VDD1.n5 VDD1.n4 78.0885
R882 VDD1.n5 VDD1.n3 43.5957
R883 VDD1.n4 VDD1.t2 3.24775
R884 VDD1.n4 VDD1.t3 3.24775
R885 VDD1.n0 VDD1.t7 3.24775
R886 VDD1.n0 VDD1.t6 3.24775
R887 VDD1.n2 VDD1.t0 3.24775
R888 VDD1.n2 VDD1.t4 3.24775
R889 VDD1.n1 VDD1.t1 3.24775
R890 VDD1.n1 VDD1.t5 3.24775
R891 VDD1 VDD1.n5 1.12766
R892 B.n381 B.n120 585
R893 B.n380 B.n379 585
R894 B.n378 B.n121 585
R895 B.n377 B.n376 585
R896 B.n375 B.n122 585
R897 B.n374 B.n373 585
R898 B.n372 B.n123 585
R899 B.n371 B.n370 585
R900 B.n369 B.n124 585
R901 B.n368 B.n367 585
R902 B.n366 B.n125 585
R903 B.n365 B.n364 585
R904 B.n363 B.n126 585
R905 B.n362 B.n361 585
R906 B.n360 B.n127 585
R907 B.n359 B.n358 585
R908 B.n357 B.n128 585
R909 B.n356 B.n355 585
R910 B.n354 B.n129 585
R911 B.n353 B.n352 585
R912 B.n351 B.n130 585
R913 B.n350 B.n349 585
R914 B.n348 B.n131 585
R915 B.n347 B.n346 585
R916 B.n345 B.n132 585
R917 B.n344 B.n343 585
R918 B.n342 B.n133 585
R919 B.n341 B.n340 585
R920 B.n339 B.n134 585
R921 B.n338 B.n337 585
R922 B.n336 B.n135 585
R923 B.n335 B.n334 585
R924 B.n333 B.n136 585
R925 B.n332 B.n331 585
R926 B.n330 B.n137 585
R927 B.n329 B.n328 585
R928 B.n327 B.n326 585
R929 B.n325 B.n141 585
R930 B.n324 B.n323 585
R931 B.n322 B.n142 585
R932 B.n321 B.n320 585
R933 B.n319 B.n143 585
R934 B.n318 B.n317 585
R935 B.n316 B.n144 585
R936 B.n315 B.n314 585
R937 B.n312 B.n145 585
R938 B.n311 B.n310 585
R939 B.n309 B.n148 585
R940 B.n308 B.n307 585
R941 B.n306 B.n149 585
R942 B.n305 B.n304 585
R943 B.n303 B.n150 585
R944 B.n302 B.n301 585
R945 B.n300 B.n151 585
R946 B.n299 B.n298 585
R947 B.n297 B.n152 585
R948 B.n296 B.n295 585
R949 B.n294 B.n153 585
R950 B.n293 B.n292 585
R951 B.n291 B.n154 585
R952 B.n290 B.n289 585
R953 B.n288 B.n155 585
R954 B.n287 B.n286 585
R955 B.n285 B.n156 585
R956 B.n284 B.n283 585
R957 B.n282 B.n157 585
R958 B.n281 B.n280 585
R959 B.n279 B.n158 585
R960 B.n278 B.n277 585
R961 B.n276 B.n159 585
R962 B.n275 B.n274 585
R963 B.n273 B.n160 585
R964 B.n272 B.n271 585
R965 B.n270 B.n161 585
R966 B.n269 B.n268 585
R967 B.n267 B.n162 585
R968 B.n266 B.n265 585
R969 B.n264 B.n163 585
R970 B.n263 B.n262 585
R971 B.n261 B.n164 585
R972 B.n260 B.n259 585
R973 B.n383 B.n382 585
R974 B.n384 B.n119 585
R975 B.n386 B.n385 585
R976 B.n387 B.n118 585
R977 B.n389 B.n388 585
R978 B.n390 B.n117 585
R979 B.n392 B.n391 585
R980 B.n393 B.n116 585
R981 B.n395 B.n394 585
R982 B.n396 B.n115 585
R983 B.n398 B.n397 585
R984 B.n399 B.n114 585
R985 B.n401 B.n400 585
R986 B.n402 B.n113 585
R987 B.n404 B.n403 585
R988 B.n405 B.n112 585
R989 B.n407 B.n406 585
R990 B.n408 B.n111 585
R991 B.n410 B.n409 585
R992 B.n411 B.n110 585
R993 B.n413 B.n412 585
R994 B.n414 B.n109 585
R995 B.n416 B.n415 585
R996 B.n417 B.n108 585
R997 B.n419 B.n418 585
R998 B.n420 B.n107 585
R999 B.n422 B.n421 585
R1000 B.n423 B.n106 585
R1001 B.n425 B.n424 585
R1002 B.n426 B.n105 585
R1003 B.n428 B.n427 585
R1004 B.n429 B.n104 585
R1005 B.n431 B.n430 585
R1006 B.n432 B.n103 585
R1007 B.n434 B.n433 585
R1008 B.n435 B.n102 585
R1009 B.n437 B.n436 585
R1010 B.n438 B.n101 585
R1011 B.n440 B.n439 585
R1012 B.n441 B.n100 585
R1013 B.n443 B.n442 585
R1014 B.n444 B.n99 585
R1015 B.n446 B.n445 585
R1016 B.n447 B.n98 585
R1017 B.n449 B.n448 585
R1018 B.n450 B.n97 585
R1019 B.n452 B.n451 585
R1020 B.n453 B.n96 585
R1021 B.n455 B.n454 585
R1022 B.n456 B.n95 585
R1023 B.n458 B.n457 585
R1024 B.n459 B.n94 585
R1025 B.n461 B.n460 585
R1026 B.n462 B.n93 585
R1027 B.n464 B.n463 585
R1028 B.n465 B.n92 585
R1029 B.n467 B.n466 585
R1030 B.n468 B.n91 585
R1031 B.n470 B.n469 585
R1032 B.n471 B.n90 585
R1033 B.n473 B.n472 585
R1034 B.n474 B.n89 585
R1035 B.n476 B.n475 585
R1036 B.n477 B.n88 585
R1037 B.n479 B.n478 585
R1038 B.n480 B.n87 585
R1039 B.n482 B.n481 585
R1040 B.n483 B.n86 585
R1041 B.n485 B.n484 585
R1042 B.n486 B.n85 585
R1043 B.n488 B.n487 585
R1044 B.n489 B.n84 585
R1045 B.n491 B.n490 585
R1046 B.n492 B.n83 585
R1047 B.n494 B.n493 585
R1048 B.n495 B.n82 585
R1049 B.n497 B.n496 585
R1050 B.n498 B.n81 585
R1051 B.n500 B.n499 585
R1052 B.n501 B.n80 585
R1053 B.n503 B.n502 585
R1054 B.n504 B.n79 585
R1055 B.n506 B.n505 585
R1056 B.n507 B.n78 585
R1057 B.n509 B.n508 585
R1058 B.n510 B.n77 585
R1059 B.n512 B.n511 585
R1060 B.n513 B.n76 585
R1061 B.n515 B.n514 585
R1062 B.n516 B.n75 585
R1063 B.n518 B.n517 585
R1064 B.n519 B.n74 585
R1065 B.n521 B.n520 585
R1066 B.n522 B.n73 585
R1067 B.n524 B.n523 585
R1068 B.n525 B.n72 585
R1069 B.n527 B.n526 585
R1070 B.n528 B.n71 585
R1071 B.n651 B.n26 585
R1072 B.n650 B.n649 585
R1073 B.n648 B.n27 585
R1074 B.n647 B.n646 585
R1075 B.n645 B.n28 585
R1076 B.n644 B.n643 585
R1077 B.n642 B.n29 585
R1078 B.n641 B.n640 585
R1079 B.n639 B.n30 585
R1080 B.n638 B.n637 585
R1081 B.n636 B.n31 585
R1082 B.n635 B.n634 585
R1083 B.n633 B.n32 585
R1084 B.n632 B.n631 585
R1085 B.n630 B.n33 585
R1086 B.n629 B.n628 585
R1087 B.n627 B.n34 585
R1088 B.n626 B.n625 585
R1089 B.n624 B.n35 585
R1090 B.n623 B.n622 585
R1091 B.n621 B.n36 585
R1092 B.n620 B.n619 585
R1093 B.n618 B.n37 585
R1094 B.n617 B.n616 585
R1095 B.n615 B.n38 585
R1096 B.n614 B.n613 585
R1097 B.n612 B.n39 585
R1098 B.n611 B.n610 585
R1099 B.n609 B.n40 585
R1100 B.n608 B.n607 585
R1101 B.n606 B.n41 585
R1102 B.n605 B.n604 585
R1103 B.n603 B.n42 585
R1104 B.n602 B.n601 585
R1105 B.n600 B.n43 585
R1106 B.n599 B.n598 585
R1107 B.n597 B.n596 585
R1108 B.n595 B.n47 585
R1109 B.n594 B.n593 585
R1110 B.n592 B.n48 585
R1111 B.n591 B.n590 585
R1112 B.n589 B.n49 585
R1113 B.n588 B.n587 585
R1114 B.n586 B.n50 585
R1115 B.n585 B.n584 585
R1116 B.n582 B.n51 585
R1117 B.n581 B.n580 585
R1118 B.n579 B.n54 585
R1119 B.n578 B.n577 585
R1120 B.n576 B.n55 585
R1121 B.n575 B.n574 585
R1122 B.n573 B.n56 585
R1123 B.n572 B.n571 585
R1124 B.n570 B.n57 585
R1125 B.n569 B.n568 585
R1126 B.n567 B.n58 585
R1127 B.n566 B.n565 585
R1128 B.n564 B.n59 585
R1129 B.n563 B.n562 585
R1130 B.n561 B.n60 585
R1131 B.n560 B.n559 585
R1132 B.n558 B.n61 585
R1133 B.n557 B.n556 585
R1134 B.n555 B.n62 585
R1135 B.n554 B.n553 585
R1136 B.n552 B.n63 585
R1137 B.n551 B.n550 585
R1138 B.n549 B.n64 585
R1139 B.n548 B.n547 585
R1140 B.n546 B.n65 585
R1141 B.n545 B.n544 585
R1142 B.n543 B.n66 585
R1143 B.n542 B.n541 585
R1144 B.n540 B.n67 585
R1145 B.n539 B.n538 585
R1146 B.n537 B.n68 585
R1147 B.n536 B.n535 585
R1148 B.n534 B.n69 585
R1149 B.n533 B.n532 585
R1150 B.n531 B.n70 585
R1151 B.n530 B.n529 585
R1152 B.n653 B.n652 585
R1153 B.n654 B.n25 585
R1154 B.n656 B.n655 585
R1155 B.n657 B.n24 585
R1156 B.n659 B.n658 585
R1157 B.n660 B.n23 585
R1158 B.n662 B.n661 585
R1159 B.n663 B.n22 585
R1160 B.n665 B.n664 585
R1161 B.n666 B.n21 585
R1162 B.n668 B.n667 585
R1163 B.n669 B.n20 585
R1164 B.n671 B.n670 585
R1165 B.n672 B.n19 585
R1166 B.n674 B.n673 585
R1167 B.n675 B.n18 585
R1168 B.n677 B.n676 585
R1169 B.n678 B.n17 585
R1170 B.n680 B.n679 585
R1171 B.n681 B.n16 585
R1172 B.n683 B.n682 585
R1173 B.n684 B.n15 585
R1174 B.n686 B.n685 585
R1175 B.n687 B.n14 585
R1176 B.n689 B.n688 585
R1177 B.n690 B.n13 585
R1178 B.n692 B.n691 585
R1179 B.n693 B.n12 585
R1180 B.n695 B.n694 585
R1181 B.n696 B.n11 585
R1182 B.n698 B.n697 585
R1183 B.n699 B.n10 585
R1184 B.n701 B.n700 585
R1185 B.n702 B.n9 585
R1186 B.n704 B.n703 585
R1187 B.n705 B.n8 585
R1188 B.n707 B.n706 585
R1189 B.n708 B.n7 585
R1190 B.n710 B.n709 585
R1191 B.n711 B.n6 585
R1192 B.n713 B.n712 585
R1193 B.n714 B.n5 585
R1194 B.n716 B.n715 585
R1195 B.n717 B.n4 585
R1196 B.n719 B.n718 585
R1197 B.n720 B.n3 585
R1198 B.n722 B.n721 585
R1199 B.n723 B.n0 585
R1200 B.n2 B.n1 585
R1201 B.n189 B.n188 585
R1202 B.n191 B.n190 585
R1203 B.n192 B.n187 585
R1204 B.n194 B.n193 585
R1205 B.n195 B.n186 585
R1206 B.n197 B.n196 585
R1207 B.n198 B.n185 585
R1208 B.n200 B.n199 585
R1209 B.n201 B.n184 585
R1210 B.n203 B.n202 585
R1211 B.n204 B.n183 585
R1212 B.n206 B.n205 585
R1213 B.n207 B.n182 585
R1214 B.n209 B.n208 585
R1215 B.n210 B.n181 585
R1216 B.n212 B.n211 585
R1217 B.n213 B.n180 585
R1218 B.n215 B.n214 585
R1219 B.n216 B.n179 585
R1220 B.n218 B.n217 585
R1221 B.n219 B.n178 585
R1222 B.n221 B.n220 585
R1223 B.n222 B.n177 585
R1224 B.n224 B.n223 585
R1225 B.n225 B.n176 585
R1226 B.n227 B.n226 585
R1227 B.n228 B.n175 585
R1228 B.n230 B.n229 585
R1229 B.n231 B.n174 585
R1230 B.n233 B.n232 585
R1231 B.n234 B.n173 585
R1232 B.n236 B.n235 585
R1233 B.n237 B.n172 585
R1234 B.n239 B.n238 585
R1235 B.n240 B.n171 585
R1236 B.n242 B.n241 585
R1237 B.n243 B.n170 585
R1238 B.n245 B.n244 585
R1239 B.n246 B.n169 585
R1240 B.n248 B.n247 585
R1241 B.n249 B.n168 585
R1242 B.n251 B.n250 585
R1243 B.n252 B.n167 585
R1244 B.n254 B.n253 585
R1245 B.n255 B.n166 585
R1246 B.n257 B.n256 585
R1247 B.n258 B.n165 585
R1248 B.n260 B.n165 516.524
R1249 B.n382 B.n381 516.524
R1250 B.n530 B.n71 516.524
R1251 B.n652 B.n651 516.524
R1252 B.n138 B.t4 393.103
R1253 B.n52 B.t11 393.103
R1254 B.n146 B.t1 393.103
R1255 B.n44 B.t8 393.103
R1256 B.n139 B.t5 339.771
R1257 B.n53 B.t10 339.771
R1258 B.n147 B.t2 339.771
R1259 B.n45 B.t7 339.771
R1260 B.n146 B.t0 307.445
R1261 B.n138 B.t3 307.445
R1262 B.n52 B.t9 307.445
R1263 B.n44 B.t6 307.445
R1264 B.n725 B.n724 256.663
R1265 B.n724 B.n723 235.042
R1266 B.n724 B.n2 235.042
R1267 B.n261 B.n260 163.367
R1268 B.n262 B.n261 163.367
R1269 B.n262 B.n163 163.367
R1270 B.n266 B.n163 163.367
R1271 B.n267 B.n266 163.367
R1272 B.n268 B.n267 163.367
R1273 B.n268 B.n161 163.367
R1274 B.n272 B.n161 163.367
R1275 B.n273 B.n272 163.367
R1276 B.n274 B.n273 163.367
R1277 B.n274 B.n159 163.367
R1278 B.n278 B.n159 163.367
R1279 B.n279 B.n278 163.367
R1280 B.n280 B.n279 163.367
R1281 B.n280 B.n157 163.367
R1282 B.n284 B.n157 163.367
R1283 B.n285 B.n284 163.367
R1284 B.n286 B.n285 163.367
R1285 B.n286 B.n155 163.367
R1286 B.n290 B.n155 163.367
R1287 B.n291 B.n290 163.367
R1288 B.n292 B.n291 163.367
R1289 B.n292 B.n153 163.367
R1290 B.n296 B.n153 163.367
R1291 B.n297 B.n296 163.367
R1292 B.n298 B.n297 163.367
R1293 B.n298 B.n151 163.367
R1294 B.n302 B.n151 163.367
R1295 B.n303 B.n302 163.367
R1296 B.n304 B.n303 163.367
R1297 B.n304 B.n149 163.367
R1298 B.n308 B.n149 163.367
R1299 B.n309 B.n308 163.367
R1300 B.n310 B.n309 163.367
R1301 B.n310 B.n145 163.367
R1302 B.n315 B.n145 163.367
R1303 B.n316 B.n315 163.367
R1304 B.n317 B.n316 163.367
R1305 B.n317 B.n143 163.367
R1306 B.n321 B.n143 163.367
R1307 B.n322 B.n321 163.367
R1308 B.n323 B.n322 163.367
R1309 B.n323 B.n141 163.367
R1310 B.n327 B.n141 163.367
R1311 B.n328 B.n327 163.367
R1312 B.n328 B.n137 163.367
R1313 B.n332 B.n137 163.367
R1314 B.n333 B.n332 163.367
R1315 B.n334 B.n333 163.367
R1316 B.n334 B.n135 163.367
R1317 B.n338 B.n135 163.367
R1318 B.n339 B.n338 163.367
R1319 B.n340 B.n339 163.367
R1320 B.n340 B.n133 163.367
R1321 B.n344 B.n133 163.367
R1322 B.n345 B.n344 163.367
R1323 B.n346 B.n345 163.367
R1324 B.n346 B.n131 163.367
R1325 B.n350 B.n131 163.367
R1326 B.n351 B.n350 163.367
R1327 B.n352 B.n351 163.367
R1328 B.n352 B.n129 163.367
R1329 B.n356 B.n129 163.367
R1330 B.n357 B.n356 163.367
R1331 B.n358 B.n357 163.367
R1332 B.n358 B.n127 163.367
R1333 B.n362 B.n127 163.367
R1334 B.n363 B.n362 163.367
R1335 B.n364 B.n363 163.367
R1336 B.n364 B.n125 163.367
R1337 B.n368 B.n125 163.367
R1338 B.n369 B.n368 163.367
R1339 B.n370 B.n369 163.367
R1340 B.n370 B.n123 163.367
R1341 B.n374 B.n123 163.367
R1342 B.n375 B.n374 163.367
R1343 B.n376 B.n375 163.367
R1344 B.n376 B.n121 163.367
R1345 B.n380 B.n121 163.367
R1346 B.n381 B.n380 163.367
R1347 B.n526 B.n71 163.367
R1348 B.n526 B.n525 163.367
R1349 B.n525 B.n524 163.367
R1350 B.n524 B.n73 163.367
R1351 B.n520 B.n73 163.367
R1352 B.n520 B.n519 163.367
R1353 B.n519 B.n518 163.367
R1354 B.n518 B.n75 163.367
R1355 B.n514 B.n75 163.367
R1356 B.n514 B.n513 163.367
R1357 B.n513 B.n512 163.367
R1358 B.n512 B.n77 163.367
R1359 B.n508 B.n77 163.367
R1360 B.n508 B.n507 163.367
R1361 B.n507 B.n506 163.367
R1362 B.n506 B.n79 163.367
R1363 B.n502 B.n79 163.367
R1364 B.n502 B.n501 163.367
R1365 B.n501 B.n500 163.367
R1366 B.n500 B.n81 163.367
R1367 B.n496 B.n81 163.367
R1368 B.n496 B.n495 163.367
R1369 B.n495 B.n494 163.367
R1370 B.n494 B.n83 163.367
R1371 B.n490 B.n83 163.367
R1372 B.n490 B.n489 163.367
R1373 B.n489 B.n488 163.367
R1374 B.n488 B.n85 163.367
R1375 B.n484 B.n85 163.367
R1376 B.n484 B.n483 163.367
R1377 B.n483 B.n482 163.367
R1378 B.n482 B.n87 163.367
R1379 B.n478 B.n87 163.367
R1380 B.n478 B.n477 163.367
R1381 B.n477 B.n476 163.367
R1382 B.n476 B.n89 163.367
R1383 B.n472 B.n89 163.367
R1384 B.n472 B.n471 163.367
R1385 B.n471 B.n470 163.367
R1386 B.n470 B.n91 163.367
R1387 B.n466 B.n91 163.367
R1388 B.n466 B.n465 163.367
R1389 B.n465 B.n464 163.367
R1390 B.n464 B.n93 163.367
R1391 B.n460 B.n93 163.367
R1392 B.n460 B.n459 163.367
R1393 B.n459 B.n458 163.367
R1394 B.n458 B.n95 163.367
R1395 B.n454 B.n95 163.367
R1396 B.n454 B.n453 163.367
R1397 B.n453 B.n452 163.367
R1398 B.n452 B.n97 163.367
R1399 B.n448 B.n97 163.367
R1400 B.n448 B.n447 163.367
R1401 B.n447 B.n446 163.367
R1402 B.n446 B.n99 163.367
R1403 B.n442 B.n99 163.367
R1404 B.n442 B.n441 163.367
R1405 B.n441 B.n440 163.367
R1406 B.n440 B.n101 163.367
R1407 B.n436 B.n101 163.367
R1408 B.n436 B.n435 163.367
R1409 B.n435 B.n434 163.367
R1410 B.n434 B.n103 163.367
R1411 B.n430 B.n103 163.367
R1412 B.n430 B.n429 163.367
R1413 B.n429 B.n428 163.367
R1414 B.n428 B.n105 163.367
R1415 B.n424 B.n105 163.367
R1416 B.n424 B.n423 163.367
R1417 B.n423 B.n422 163.367
R1418 B.n422 B.n107 163.367
R1419 B.n418 B.n107 163.367
R1420 B.n418 B.n417 163.367
R1421 B.n417 B.n416 163.367
R1422 B.n416 B.n109 163.367
R1423 B.n412 B.n109 163.367
R1424 B.n412 B.n411 163.367
R1425 B.n411 B.n410 163.367
R1426 B.n410 B.n111 163.367
R1427 B.n406 B.n111 163.367
R1428 B.n406 B.n405 163.367
R1429 B.n405 B.n404 163.367
R1430 B.n404 B.n113 163.367
R1431 B.n400 B.n113 163.367
R1432 B.n400 B.n399 163.367
R1433 B.n399 B.n398 163.367
R1434 B.n398 B.n115 163.367
R1435 B.n394 B.n115 163.367
R1436 B.n394 B.n393 163.367
R1437 B.n393 B.n392 163.367
R1438 B.n392 B.n117 163.367
R1439 B.n388 B.n117 163.367
R1440 B.n388 B.n387 163.367
R1441 B.n387 B.n386 163.367
R1442 B.n386 B.n119 163.367
R1443 B.n382 B.n119 163.367
R1444 B.n651 B.n650 163.367
R1445 B.n650 B.n27 163.367
R1446 B.n646 B.n27 163.367
R1447 B.n646 B.n645 163.367
R1448 B.n645 B.n644 163.367
R1449 B.n644 B.n29 163.367
R1450 B.n640 B.n29 163.367
R1451 B.n640 B.n639 163.367
R1452 B.n639 B.n638 163.367
R1453 B.n638 B.n31 163.367
R1454 B.n634 B.n31 163.367
R1455 B.n634 B.n633 163.367
R1456 B.n633 B.n632 163.367
R1457 B.n632 B.n33 163.367
R1458 B.n628 B.n33 163.367
R1459 B.n628 B.n627 163.367
R1460 B.n627 B.n626 163.367
R1461 B.n626 B.n35 163.367
R1462 B.n622 B.n35 163.367
R1463 B.n622 B.n621 163.367
R1464 B.n621 B.n620 163.367
R1465 B.n620 B.n37 163.367
R1466 B.n616 B.n37 163.367
R1467 B.n616 B.n615 163.367
R1468 B.n615 B.n614 163.367
R1469 B.n614 B.n39 163.367
R1470 B.n610 B.n39 163.367
R1471 B.n610 B.n609 163.367
R1472 B.n609 B.n608 163.367
R1473 B.n608 B.n41 163.367
R1474 B.n604 B.n41 163.367
R1475 B.n604 B.n603 163.367
R1476 B.n603 B.n602 163.367
R1477 B.n602 B.n43 163.367
R1478 B.n598 B.n43 163.367
R1479 B.n598 B.n597 163.367
R1480 B.n597 B.n47 163.367
R1481 B.n593 B.n47 163.367
R1482 B.n593 B.n592 163.367
R1483 B.n592 B.n591 163.367
R1484 B.n591 B.n49 163.367
R1485 B.n587 B.n49 163.367
R1486 B.n587 B.n586 163.367
R1487 B.n586 B.n585 163.367
R1488 B.n585 B.n51 163.367
R1489 B.n580 B.n51 163.367
R1490 B.n580 B.n579 163.367
R1491 B.n579 B.n578 163.367
R1492 B.n578 B.n55 163.367
R1493 B.n574 B.n55 163.367
R1494 B.n574 B.n573 163.367
R1495 B.n573 B.n572 163.367
R1496 B.n572 B.n57 163.367
R1497 B.n568 B.n57 163.367
R1498 B.n568 B.n567 163.367
R1499 B.n567 B.n566 163.367
R1500 B.n566 B.n59 163.367
R1501 B.n562 B.n59 163.367
R1502 B.n562 B.n561 163.367
R1503 B.n561 B.n560 163.367
R1504 B.n560 B.n61 163.367
R1505 B.n556 B.n61 163.367
R1506 B.n556 B.n555 163.367
R1507 B.n555 B.n554 163.367
R1508 B.n554 B.n63 163.367
R1509 B.n550 B.n63 163.367
R1510 B.n550 B.n549 163.367
R1511 B.n549 B.n548 163.367
R1512 B.n548 B.n65 163.367
R1513 B.n544 B.n65 163.367
R1514 B.n544 B.n543 163.367
R1515 B.n543 B.n542 163.367
R1516 B.n542 B.n67 163.367
R1517 B.n538 B.n67 163.367
R1518 B.n538 B.n537 163.367
R1519 B.n537 B.n536 163.367
R1520 B.n536 B.n69 163.367
R1521 B.n532 B.n69 163.367
R1522 B.n532 B.n531 163.367
R1523 B.n531 B.n530 163.367
R1524 B.n652 B.n25 163.367
R1525 B.n656 B.n25 163.367
R1526 B.n657 B.n656 163.367
R1527 B.n658 B.n657 163.367
R1528 B.n658 B.n23 163.367
R1529 B.n662 B.n23 163.367
R1530 B.n663 B.n662 163.367
R1531 B.n664 B.n663 163.367
R1532 B.n664 B.n21 163.367
R1533 B.n668 B.n21 163.367
R1534 B.n669 B.n668 163.367
R1535 B.n670 B.n669 163.367
R1536 B.n670 B.n19 163.367
R1537 B.n674 B.n19 163.367
R1538 B.n675 B.n674 163.367
R1539 B.n676 B.n675 163.367
R1540 B.n676 B.n17 163.367
R1541 B.n680 B.n17 163.367
R1542 B.n681 B.n680 163.367
R1543 B.n682 B.n681 163.367
R1544 B.n682 B.n15 163.367
R1545 B.n686 B.n15 163.367
R1546 B.n687 B.n686 163.367
R1547 B.n688 B.n687 163.367
R1548 B.n688 B.n13 163.367
R1549 B.n692 B.n13 163.367
R1550 B.n693 B.n692 163.367
R1551 B.n694 B.n693 163.367
R1552 B.n694 B.n11 163.367
R1553 B.n698 B.n11 163.367
R1554 B.n699 B.n698 163.367
R1555 B.n700 B.n699 163.367
R1556 B.n700 B.n9 163.367
R1557 B.n704 B.n9 163.367
R1558 B.n705 B.n704 163.367
R1559 B.n706 B.n705 163.367
R1560 B.n706 B.n7 163.367
R1561 B.n710 B.n7 163.367
R1562 B.n711 B.n710 163.367
R1563 B.n712 B.n711 163.367
R1564 B.n712 B.n5 163.367
R1565 B.n716 B.n5 163.367
R1566 B.n717 B.n716 163.367
R1567 B.n718 B.n717 163.367
R1568 B.n718 B.n3 163.367
R1569 B.n722 B.n3 163.367
R1570 B.n723 B.n722 163.367
R1571 B.n189 B.n2 163.367
R1572 B.n190 B.n189 163.367
R1573 B.n190 B.n187 163.367
R1574 B.n194 B.n187 163.367
R1575 B.n195 B.n194 163.367
R1576 B.n196 B.n195 163.367
R1577 B.n196 B.n185 163.367
R1578 B.n200 B.n185 163.367
R1579 B.n201 B.n200 163.367
R1580 B.n202 B.n201 163.367
R1581 B.n202 B.n183 163.367
R1582 B.n206 B.n183 163.367
R1583 B.n207 B.n206 163.367
R1584 B.n208 B.n207 163.367
R1585 B.n208 B.n181 163.367
R1586 B.n212 B.n181 163.367
R1587 B.n213 B.n212 163.367
R1588 B.n214 B.n213 163.367
R1589 B.n214 B.n179 163.367
R1590 B.n218 B.n179 163.367
R1591 B.n219 B.n218 163.367
R1592 B.n220 B.n219 163.367
R1593 B.n220 B.n177 163.367
R1594 B.n224 B.n177 163.367
R1595 B.n225 B.n224 163.367
R1596 B.n226 B.n225 163.367
R1597 B.n226 B.n175 163.367
R1598 B.n230 B.n175 163.367
R1599 B.n231 B.n230 163.367
R1600 B.n232 B.n231 163.367
R1601 B.n232 B.n173 163.367
R1602 B.n236 B.n173 163.367
R1603 B.n237 B.n236 163.367
R1604 B.n238 B.n237 163.367
R1605 B.n238 B.n171 163.367
R1606 B.n242 B.n171 163.367
R1607 B.n243 B.n242 163.367
R1608 B.n244 B.n243 163.367
R1609 B.n244 B.n169 163.367
R1610 B.n248 B.n169 163.367
R1611 B.n249 B.n248 163.367
R1612 B.n250 B.n249 163.367
R1613 B.n250 B.n167 163.367
R1614 B.n254 B.n167 163.367
R1615 B.n255 B.n254 163.367
R1616 B.n256 B.n255 163.367
R1617 B.n256 B.n165 163.367
R1618 B.n313 B.n147 59.5399
R1619 B.n140 B.n139 59.5399
R1620 B.n583 B.n53 59.5399
R1621 B.n46 B.n45 59.5399
R1622 B.n147 B.n146 53.3338
R1623 B.n139 B.n138 53.3338
R1624 B.n53 B.n52 53.3338
R1625 B.n45 B.n44 53.3338
R1626 B.n653 B.n26 33.5615
R1627 B.n529 B.n528 33.5615
R1628 B.n383 B.n120 33.5615
R1629 B.n259 B.n258 33.5615
R1630 B B.n725 18.0485
R1631 B.n654 B.n653 10.6151
R1632 B.n655 B.n654 10.6151
R1633 B.n655 B.n24 10.6151
R1634 B.n659 B.n24 10.6151
R1635 B.n660 B.n659 10.6151
R1636 B.n661 B.n660 10.6151
R1637 B.n661 B.n22 10.6151
R1638 B.n665 B.n22 10.6151
R1639 B.n666 B.n665 10.6151
R1640 B.n667 B.n666 10.6151
R1641 B.n667 B.n20 10.6151
R1642 B.n671 B.n20 10.6151
R1643 B.n672 B.n671 10.6151
R1644 B.n673 B.n672 10.6151
R1645 B.n673 B.n18 10.6151
R1646 B.n677 B.n18 10.6151
R1647 B.n678 B.n677 10.6151
R1648 B.n679 B.n678 10.6151
R1649 B.n679 B.n16 10.6151
R1650 B.n683 B.n16 10.6151
R1651 B.n684 B.n683 10.6151
R1652 B.n685 B.n684 10.6151
R1653 B.n685 B.n14 10.6151
R1654 B.n689 B.n14 10.6151
R1655 B.n690 B.n689 10.6151
R1656 B.n691 B.n690 10.6151
R1657 B.n691 B.n12 10.6151
R1658 B.n695 B.n12 10.6151
R1659 B.n696 B.n695 10.6151
R1660 B.n697 B.n696 10.6151
R1661 B.n697 B.n10 10.6151
R1662 B.n701 B.n10 10.6151
R1663 B.n702 B.n701 10.6151
R1664 B.n703 B.n702 10.6151
R1665 B.n703 B.n8 10.6151
R1666 B.n707 B.n8 10.6151
R1667 B.n708 B.n707 10.6151
R1668 B.n709 B.n708 10.6151
R1669 B.n709 B.n6 10.6151
R1670 B.n713 B.n6 10.6151
R1671 B.n714 B.n713 10.6151
R1672 B.n715 B.n714 10.6151
R1673 B.n715 B.n4 10.6151
R1674 B.n719 B.n4 10.6151
R1675 B.n720 B.n719 10.6151
R1676 B.n721 B.n720 10.6151
R1677 B.n721 B.n0 10.6151
R1678 B.n649 B.n26 10.6151
R1679 B.n649 B.n648 10.6151
R1680 B.n648 B.n647 10.6151
R1681 B.n647 B.n28 10.6151
R1682 B.n643 B.n28 10.6151
R1683 B.n643 B.n642 10.6151
R1684 B.n642 B.n641 10.6151
R1685 B.n641 B.n30 10.6151
R1686 B.n637 B.n30 10.6151
R1687 B.n637 B.n636 10.6151
R1688 B.n636 B.n635 10.6151
R1689 B.n635 B.n32 10.6151
R1690 B.n631 B.n32 10.6151
R1691 B.n631 B.n630 10.6151
R1692 B.n630 B.n629 10.6151
R1693 B.n629 B.n34 10.6151
R1694 B.n625 B.n34 10.6151
R1695 B.n625 B.n624 10.6151
R1696 B.n624 B.n623 10.6151
R1697 B.n623 B.n36 10.6151
R1698 B.n619 B.n36 10.6151
R1699 B.n619 B.n618 10.6151
R1700 B.n618 B.n617 10.6151
R1701 B.n617 B.n38 10.6151
R1702 B.n613 B.n38 10.6151
R1703 B.n613 B.n612 10.6151
R1704 B.n612 B.n611 10.6151
R1705 B.n611 B.n40 10.6151
R1706 B.n607 B.n40 10.6151
R1707 B.n607 B.n606 10.6151
R1708 B.n606 B.n605 10.6151
R1709 B.n605 B.n42 10.6151
R1710 B.n601 B.n42 10.6151
R1711 B.n601 B.n600 10.6151
R1712 B.n600 B.n599 10.6151
R1713 B.n596 B.n595 10.6151
R1714 B.n595 B.n594 10.6151
R1715 B.n594 B.n48 10.6151
R1716 B.n590 B.n48 10.6151
R1717 B.n590 B.n589 10.6151
R1718 B.n589 B.n588 10.6151
R1719 B.n588 B.n50 10.6151
R1720 B.n584 B.n50 10.6151
R1721 B.n582 B.n581 10.6151
R1722 B.n581 B.n54 10.6151
R1723 B.n577 B.n54 10.6151
R1724 B.n577 B.n576 10.6151
R1725 B.n576 B.n575 10.6151
R1726 B.n575 B.n56 10.6151
R1727 B.n571 B.n56 10.6151
R1728 B.n571 B.n570 10.6151
R1729 B.n570 B.n569 10.6151
R1730 B.n569 B.n58 10.6151
R1731 B.n565 B.n58 10.6151
R1732 B.n565 B.n564 10.6151
R1733 B.n564 B.n563 10.6151
R1734 B.n563 B.n60 10.6151
R1735 B.n559 B.n60 10.6151
R1736 B.n559 B.n558 10.6151
R1737 B.n558 B.n557 10.6151
R1738 B.n557 B.n62 10.6151
R1739 B.n553 B.n62 10.6151
R1740 B.n553 B.n552 10.6151
R1741 B.n552 B.n551 10.6151
R1742 B.n551 B.n64 10.6151
R1743 B.n547 B.n64 10.6151
R1744 B.n547 B.n546 10.6151
R1745 B.n546 B.n545 10.6151
R1746 B.n545 B.n66 10.6151
R1747 B.n541 B.n66 10.6151
R1748 B.n541 B.n540 10.6151
R1749 B.n540 B.n539 10.6151
R1750 B.n539 B.n68 10.6151
R1751 B.n535 B.n68 10.6151
R1752 B.n535 B.n534 10.6151
R1753 B.n534 B.n533 10.6151
R1754 B.n533 B.n70 10.6151
R1755 B.n529 B.n70 10.6151
R1756 B.n528 B.n527 10.6151
R1757 B.n527 B.n72 10.6151
R1758 B.n523 B.n72 10.6151
R1759 B.n523 B.n522 10.6151
R1760 B.n522 B.n521 10.6151
R1761 B.n521 B.n74 10.6151
R1762 B.n517 B.n74 10.6151
R1763 B.n517 B.n516 10.6151
R1764 B.n516 B.n515 10.6151
R1765 B.n515 B.n76 10.6151
R1766 B.n511 B.n76 10.6151
R1767 B.n511 B.n510 10.6151
R1768 B.n510 B.n509 10.6151
R1769 B.n509 B.n78 10.6151
R1770 B.n505 B.n78 10.6151
R1771 B.n505 B.n504 10.6151
R1772 B.n504 B.n503 10.6151
R1773 B.n503 B.n80 10.6151
R1774 B.n499 B.n80 10.6151
R1775 B.n499 B.n498 10.6151
R1776 B.n498 B.n497 10.6151
R1777 B.n497 B.n82 10.6151
R1778 B.n493 B.n82 10.6151
R1779 B.n493 B.n492 10.6151
R1780 B.n492 B.n491 10.6151
R1781 B.n491 B.n84 10.6151
R1782 B.n487 B.n84 10.6151
R1783 B.n487 B.n486 10.6151
R1784 B.n486 B.n485 10.6151
R1785 B.n485 B.n86 10.6151
R1786 B.n481 B.n86 10.6151
R1787 B.n481 B.n480 10.6151
R1788 B.n480 B.n479 10.6151
R1789 B.n479 B.n88 10.6151
R1790 B.n475 B.n88 10.6151
R1791 B.n475 B.n474 10.6151
R1792 B.n474 B.n473 10.6151
R1793 B.n473 B.n90 10.6151
R1794 B.n469 B.n90 10.6151
R1795 B.n469 B.n468 10.6151
R1796 B.n468 B.n467 10.6151
R1797 B.n467 B.n92 10.6151
R1798 B.n463 B.n92 10.6151
R1799 B.n463 B.n462 10.6151
R1800 B.n462 B.n461 10.6151
R1801 B.n461 B.n94 10.6151
R1802 B.n457 B.n94 10.6151
R1803 B.n457 B.n456 10.6151
R1804 B.n456 B.n455 10.6151
R1805 B.n455 B.n96 10.6151
R1806 B.n451 B.n96 10.6151
R1807 B.n451 B.n450 10.6151
R1808 B.n450 B.n449 10.6151
R1809 B.n449 B.n98 10.6151
R1810 B.n445 B.n98 10.6151
R1811 B.n445 B.n444 10.6151
R1812 B.n444 B.n443 10.6151
R1813 B.n443 B.n100 10.6151
R1814 B.n439 B.n100 10.6151
R1815 B.n439 B.n438 10.6151
R1816 B.n438 B.n437 10.6151
R1817 B.n437 B.n102 10.6151
R1818 B.n433 B.n102 10.6151
R1819 B.n433 B.n432 10.6151
R1820 B.n432 B.n431 10.6151
R1821 B.n431 B.n104 10.6151
R1822 B.n427 B.n104 10.6151
R1823 B.n427 B.n426 10.6151
R1824 B.n426 B.n425 10.6151
R1825 B.n425 B.n106 10.6151
R1826 B.n421 B.n106 10.6151
R1827 B.n421 B.n420 10.6151
R1828 B.n420 B.n419 10.6151
R1829 B.n419 B.n108 10.6151
R1830 B.n415 B.n108 10.6151
R1831 B.n415 B.n414 10.6151
R1832 B.n414 B.n413 10.6151
R1833 B.n413 B.n110 10.6151
R1834 B.n409 B.n110 10.6151
R1835 B.n409 B.n408 10.6151
R1836 B.n408 B.n407 10.6151
R1837 B.n407 B.n112 10.6151
R1838 B.n403 B.n112 10.6151
R1839 B.n403 B.n402 10.6151
R1840 B.n402 B.n401 10.6151
R1841 B.n401 B.n114 10.6151
R1842 B.n397 B.n114 10.6151
R1843 B.n397 B.n396 10.6151
R1844 B.n396 B.n395 10.6151
R1845 B.n395 B.n116 10.6151
R1846 B.n391 B.n116 10.6151
R1847 B.n391 B.n390 10.6151
R1848 B.n390 B.n389 10.6151
R1849 B.n389 B.n118 10.6151
R1850 B.n385 B.n118 10.6151
R1851 B.n385 B.n384 10.6151
R1852 B.n384 B.n383 10.6151
R1853 B.n188 B.n1 10.6151
R1854 B.n191 B.n188 10.6151
R1855 B.n192 B.n191 10.6151
R1856 B.n193 B.n192 10.6151
R1857 B.n193 B.n186 10.6151
R1858 B.n197 B.n186 10.6151
R1859 B.n198 B.n197 10.6151
R1860 B.n199 B.n198 10.6151
R1861 B.n199 B.n184 10.6151
R1862 B.n203 B.n184 10.6151
R1863 B.n204 B.n203 10.6151
R1864 B.n205 B.n204 10.6151
R1865 B.n205 B.n182 10.6151
R1866 B.n209 B.n182 10.6151
R1867 B.n210 B.n209 10.6151
R1868 B.n211 B.n210 10.6151
R1869 B.n211 B.n180 10.6151
R1870 B.n215 B.n180 10.6151
R1871 B.n216 B.n215 10.6151
R1872 B.n217 B.n216 10.6151
R1873 B.n217 B.n178 10.6151
R1874 B.n221 B.n178 10.6151
R1875 B.n222 B.n221 10.6151
R1876 B.n223 B.n222 10.6151
R1877 B.n223 B.n176 10.6151
R1878 B.n227 B.n176 10.6151
R1879 B.n228 B.n227 10.6151
R1880 B.n229 B.n228 10.6151
R1881 B.n229 B.n174 10.6151
R1882 B.n233 B.n174 10.6151
R1883 B.n234 B.n233 10.6151
R1884 B.n235 B.n234 10.6151
R1885 B.n235 B.n172 10.6151
R1886 B.n239 B.n172 10.6151
R1887 B.n240 B.n239 10.6151
R1888 B.n241 B.n240 10.6151
R1889 B.n241 B.n170 10.6151
R1890 B.n245 B.n170 10.6151
R1891 B.n246 B.n245 10.6151
R1892 B.n247 B.n246 10.6151
R1893 B.n247 B.n168 10.6151
R1894 B.n251 B.n168 10.6151
R1895 B.n252 B.n251 10.6151
R1896 B.n253 B.n252 10.6151
R1897 B.n253 B.n166 10.6151
R1898 B.n257 B.n166 10.6151
R1899 B.n258 B.n257 10.6151
R1900 B.n259 B.n164 10.6151
R1901 B.n263 B.n164 10.6151
R1902 B.n264 B.n263 10.6151
R1903 B.n265 B.n264 10.6151
R1904 B.n265 B.n162 10.6151
R1905 B.n269 B.n162 10.6151
R1906 B.n270 B.n269 10.6151
R1907 B.n271 B.n270 10.6151
R1908 B.n271 B.n160 10.6151
R1909 B.n275 B.n160 10.6151
R1910 B.n276 B.n275 10.6151
R1911 B.n277 B.n276 10.6151
R1912 B.n277 B.n158 10.6151
R1913 B.n281 B.n158 10.6151
R1914 B.n282 B.n281 10.6151
R1915 B.n283 B.n282 10.6151
R1916 B.n283 B.n156 10.6151
R1917 B.n287 B.n156 10.6151
R1918 B.n288 B.n287 10.6151
R1919 B.n289 B.n288 10.6151
R1920 B.n289 B.n154 10.6151
R1921 B.n293 B.n154 10.6151
R1922 B.n294 B.n293 10.6151
R1923 B.n295 B.n294 10.6151
R1924 B.n295 B.n152 10.6151
R1925 B.n299 B.n152 10.6151
R1926 B.n300 B.n299 10.6151
R1927 B.n301 B.n300 10.6151
R1928 B.n301 B.n150 10.6151
R1929 B.n305 B.n150 10.6151
R1930 B.n306 B.n305 10.6151
R1931 B.n307 B.n306 10.6151
R1932 B.n307 B.n148 10.6151
R1933 B.n311 B.n148 10.6151
R1934 B.n312 B.n311 10.6151
R1935 B.n314 B.n144 10.6151
R1936 B.n318 B.n144 10.6151
R1937 B.n319 B.n318 10.6151
R1938 B.n320 B.n319 10.6151
R1939 B.n320 B.n142 10.6151
R1940 B.n324 B.n142 10.6151
R1941 B.n325 B.n324 10.6151
R1942 B.n326 B.n325 10.6151
R1943 B.n330 B.n329 10.6151
R1944 B.n331 B.n330 10.6151
R1945 B.n331 B.n136 10.6151
R1946 B.n335 B.n136 10.6151
R1947 B.n336 B.n335 10.6151
R1948 B.n337 B.n336 10.6151
R1949 B.n337 B.n134 10.6151
R1950 B.n341 B.n134 10.6151
R1951 B.n342 B.n341 10.6151
R1952 B.n343 B.n342 10.6151
R1953 B.n343 B.n132 10.6151
R1954 B.n347 B.n132 10.6151
R1955 B.n348 B.n347 10.6151
R1956 B.n349 B.n348 10.6151
R1957 B.n349 B.n130 10.6151
R1958 B.n353 B.n130 10.6151
R1959 B.n354 B.n353 10.6151
R1960 B.n355 B.n354 10.6151
R1961 B.n355 B.n128 10.6151
R1962 B.n359 B.n128 10.6151
R1963 B.n360 B.n359 10.6151
R1964 B.n361 B.n360 10.6151
R1965 B.n361 B.n126 10.6151
R1966 B.n365 B.n126 10.6151
R1967 B.n366 B.n365 10.6151
R1968 B.n367 B.n366 10.6151
R1969 B.n367 B.n124 10.6151
R1970 B.n371 B.n124 10.6151
R1971 B.n372 B.n371 10.6151
R1972 B.n373 B.n372 10.6151
R1973 B.n373 B.n122 10.6151
R1974 B.n377 B.n122 10.6151
R1975 B.n378 B.n377 10.6151
R1976 B.n379 B.n378 10.6151
R1977 B.n379 B.n120 10.6151
R1978 B.n725 B.n0 8.11757
R1979 B.n725 B.n1 8.11757
R1980 B.n596 B.n46 6.5566
R1981 B.n584 B.n583 6.5566
R1982 B.n314 B.n313 6.5566
R1983 B.n326 B.n140 6.5566
R1984 B.n599 B.n46 4.05904
R1985 B.n583 B.n582 4.05904
R1986 B.n313 B.n312 4.05904
R1987 B.n329 B.n140 4.05904
C0 VDD2 VDD1 1.68443f
C1 B VN 1.15999f
C2 VTAIL VN 7.64781f
C3 B VDD2 1.63253f
C4 VTAIL VDD2 7.41208f
C5 VDD2 VN 7.21494f
C6 w_n3720_n2970# VP 7.97594f
C7 VDD1 VP 7.56275f
C8 B VP 1.9677f
C9 VTAIL VP 7.66192f
C10 w_n3720_n2970# VDD1 1.84555f
C11 VN VP 7.07819f
C12 B w_n3720_n2970# 9.28242f
C13 VTAIL w_n3720_n2970# 3.74149f
C14 VDD2 VP 0.500617f
C15 w_n3720_n2970# VN 7.493529f
C16 w_n3720_n2970# VDD2 1.95271f
C17 B VDD1 1.54217f
C18 VTAIL VDD1 7.35887f
C19 VDD1 VN 0.151502f
C20 VTAIL B 4.25354f
C21 VDD2 VSUBS 1.669347f
C22 VDD1 VSUBS 2.295449f
C23 VTAIL VSUBS 1.215728f
C24 VN VSUBS 6.4347f
C25 VP VSUBS 3.323056f
C26 B VSUBS 4.629606f
C27 w_n3720_n2970# VSUBS 0.136464p
C28 B.n0 VSUBS 0.00632f
C29 B.n1 VSUBS 0.00632f
C30 B.n2 VSUBS 0.009347f
C31 B.n3 VSUBS 0.007163f
C32 B.n4 VSUBS 0.007163f
C33 B.n5 VSUBS 0.007163f
C34 B.n6 VSUBS 0.007163f
C35 B.n7 VSUBS 0.007163f
C36 B.n8 VSUBS 0.007163f
C37 B.n9 VSUBS 0.007163f
C38 B.n10 VSUBS 0.007163f
C39 B.n11 VSUBS 0.007163f
C40 B.n12 VSUBS 0.007163f
C41 B.n13 VSUBS 0.007163f
C42 B.n14 VSUBS 0.007163f
C43 B.n15 VSUBS 0.007163f
C44 B.n16 VSUBS 0.007163f
C45 B.n17 VSUBS 0.007163f
C46 B.n18 VSUBS 0.007163f
C47 B.n19 VSUBS 0.007163f
C48 B.n20 VSUBS 0.007163f
C49 B.n21 VSUBS 0.007163f
C50 B.n22 VSUBS 0.007163f
C51 B.n23 VSUBS 0.007163f
C52 B.n24 VSUBS 0.007163f
C53 B.n25 VSUBS 0.007163f
C54 B.n26 VSUBS 0.017457f
C55 B.n27 VSUBS 0.007163f
C56 B.n28 VSUBS 0.007163f
C57 B.n29 VSUBS 0.007163f
C58 B.n30 VSUBS 0.007163f
C59 B.n31 VSUBS 0.007163f
C60 B.n32 VSUBS 0.007163f
C61 B.n33 VSUBS 0.007163f
C62 B.n34 VSUBS 0.007163f
C63 B.n35 VSUBS 0.007163f
C64 B.n36 VSUBS 0.007163f
C65 B.n37 VSUBS 0.007163f
C66 B.n38 VSUBS 0.007163f
C67 B.n39 VSUBS 0.007163f
C68 B.n40 VSUBS 0.007163f
C69 B.n41 VSUBS 0.007163f
C70 B.n42 VSUBS 0.007163f
C71 B.n43 VSUBS 0.007163f
C72 B.t7 VSUBS 0.171623f
C73 B.t8 VSUBS 0.20112f
C74 B.t6 VSUBS 1.13617f
C75 B.n44 VSUBS 0.325429f
C76 B.n45 VSUBS 0.227632f
C77 B.n46 VSUBS 0.016596f
C78 B.n47 VSUBS 0.007163f
C79 B.n48 VSUBS 0.007163f
C80 B.n49 VSUBS 0.007163f
C81 B.n50 VSUBS 0.007163f
C82 B.n51 VSUBS 0.007163f
C83 B.t10 VSUBS 0.171626f
C84 B.t11 VSUBS 0.201123f
C85 B.t9 VSUBS 1.13617f
C86 B.n52 VSUBS 0.325427f
C87 B.n53 VSUBS 0.22763f
C88 B.n54 VSUBS 0.007163f
C89 B.n55 VSUBS 0.007163f
C90 B.n56 VSUBS 0.007163f
C91 B.n57 VSUBS 0.007163f
C92 B.n58 VSUBS 0.007163f
C93 B.n59 VSUBS 0.007163f
C94 B.n60 VSUBS 0.007163f
C95 B.n61 VSUBS 0.007163f
C96 B.n62 VSUBS 0.007163f
C97 B.n63 VSUBS 0.007163f
C98 B.n64 VSUBS 0.007163f
C99 B.n65 VSUBS 0.007163f
C100 B.n66 VSUBS 0.007163f
C101 B.n67 VSUBS 0.007163f
C102 B.n68 VSUBS 0.007163f
C103 B.n69 VSUBS 0.007163f
C104 B.n70 VSUBS 0.007163f
C105 B.n71 VSUBS 0.016673f
C106 B.n72 VSUBS 0.007163f
C107 B.n73 VSUBS 0.007163f
C108 B.n74 VSUBS 0.007163f
C109 B.n75 VSUBS 0.007163f
C110 B.n76 VSUBS 0.007163f
C111 B.n77 VSUBS 0.007163f
C112 B.n78 VSUBS 0.007163f
C113 B.n79 VSUBS 0.007163f
C114 B.n80 VSUBS 0.007163f
C115 B.n81 VSUBS 0.007163f
C116 B.n82 VSUBS 0.007163f
C117 B.n83 VSUBS 0.007163f
C118 B.n84 VSUBS 0.007163f
C119 B.n85 VSUBS 0.007163f
C120 B.n86 VSUBS 0.007163f
C121 B.n87 VSUBS 0.007163f
C122 B.n88 VSUBS 0.007163f
C123 B.n89 VSUBS 0.007163f
C124 B.n90 VSUBS 0.007163f
C125 B.n91 VSUBS 0.007163f
C126 B.n92 VSUBS 0.007163f
C127 B.n93 VSUBS 0.007163f
C128 B.n94 VSUBS 0.007163f
C129 B.n95 VSUBS 0.007163f
C130 B.n96 VSUBS 0.007163f
C131 B.n97 VSUBS 0.007163f
C132 B.n98 VSUBS 0.007163f
C133 B.n99 VSUBS 0.007163f
C134 B.n100 VSUBS 0.007163f
C135 B.n101 VSUBS 0.007163f
C136 B.n102 VSUBS 0.007163f
C137 B.n103 VSUBS 0.007163f
C138 B.n104 VSUBS 0.007163f
C139 B.n105 VSUBS 0.007163f
C140 B.n106 VSUBS 0.007163f
C141 B.n107 VSUBS 0.007163f
C142 B.n108 VSUBS 0.007163f
C143 B.n109 VSUBS 0.007163f
C144 B.n110 VSUBS 0.007163f
C145 B.n111 VSUBS 0.007163f
C146 B.n112 VSUBS 0.007163f
C147 B.n113 VSUBS 0.007163f
C148 B.n114 VSUBS 0.007163f
C149 B.n115 VSUBS 0.007163f
C150 B.n116 VSUBS 0.007163f
C151 B.n117 VSUBS 0.007163f
C152 B.n118 VSUBS 0.007163f
C153 B.n119 VSUBS 0.007163f
C154 B.n120 VSUBS 0.016633f
C155 B.n121 VSUBS 0.007163f
C156 B.n122 VSUBS 0.007163f
C157 B.n123 VSUBS 0.007163f
C158 B.n124 VSUBS 0.007163f
C159 B.n125 VSUBS 0.007163f
C160 B.n126 VSUBS 0.007163f
C161 B.n127 VSUBS 0.007163f
C162 B.n128 VSUBS 0.007163f
C163 B.n129 VSUBS 0.007163f
C164 B.n130 VSUBS 0.007163f
C165 B.n131 VSUBS 0.007163f
C166 B.n132 VSUBS 0.007163f
C167 B.n133 VSUBS 0.007163f
C168 B.n134 VSUBS 0.007163f
C169 B.n135 VSUBS 0.007163f
C170 B.n136 VSUBS 0.007163f
C171 B.n137 VSUBS 0.007163f
C172 B.t5 VSUBS 0.171626f
C173 B.t4 VSUBS 0.201123f
C174 B.t3 VSUBS 1.13617f
C175 B.n138 VSUBS 0.325427f
C176 B.n139 VSUBS 0.22763f
C177 B.n140 VSUBS 0.016596f
C178 B.n141 VSUBS 0.007163f
C179 B.n142 VSUBS 0.007163f
C180 B.n143 VSUBS 0.007163f
C181 B.n144 VSUBS 0.007163f
C182 B.n145 VSUBS 0.007163f
C183 B.t2 VSUBS 0.171623f
C184 B.t1 VSUBS 0.20112f
C185 B.t0 VSUBS 1.13617f
C186 B.n146 VSUBS 0.325429f
C187 B.n147 VSUBS 0.227632f
C188 B.n148 VSUBS 0.007163f
C189 B.n149 VSUBS 0.007163f
C190 B.n150 VSUBS 0.007163f
C191 B.n151 VSUBS 0.007163f
C192 B.n152 VSUBS 0.007163f
C193 B.n153 VSUBS 0.007163f
C194 B.n154 VSUBS 0.007163f
C195 B.n155 VSUBS 0.007163f
C196 B.n156 VSUBS 0.007163f
C197 B.n157 VSUBS 0.007163f
C198 B.n158 VSUBS 0.007163f
C199 B.n159 VSUBS 0.007163f
C200 B.n160 VSUBS 0.007163f
C201 B.n161 VSUBS 0.007163f
C202 B.n162 VSUBS 0.007163f
C203 B.n163 VSUBS 0.007163f
C204 B.n164 VSUBS 0.007163f
C205 B.n165 VSUBS 0.016673f
C206 B.n166 VSUBS 0.007163f
C207 B.n167 VSUBS 0.007163f
C208 B.n168 VSUBS 0.007163f
C209 B.n169 VSUBS 0.007163f
C210 B.n170 VSUBS 0.007163f
C211 B.n171 VSUBS 0.007163f
C212 B.n172 VSUBS 0.007163f
C213 B.n173 VSUBS 0.007163f
C214 B.n174 VSUBS 0.007163f
C215 B.n175 VSUBS 0.007163f
C216 B.n176 VSUBS 0.007163f
C217 B.n177 VSUBS 0.007163f
C218 B.n178 VSUBS 0.007163f
C219 B.n179 VSUBS 0.007163f
C220 B.n180 VSUBS 0.007163f
C221 B.n181 VSUBS 0.007163f
C222 B.n182 VSUBS 0.007163f
C223 B.n183 VSUBS 0.007163f
C224 B.n184 VSUBS 0.007163f
C225 B.n185 VSUBS 0.007163f
C226 B.n186 VSUBS 0.007163f
C227 B.n187 VSUBS 0.007163f
C228 B.n188 VSUBS 0.007163f
C229 B.n189 VSUBS 0.007163f
C230 B.n190 VSUBS 0.007163f
C231 B.n191 VSUBS 0.007163f
C232 B.n192 VSUBS 0.007163f
C233 B.n193 VSUBS 0.007163f
C234 B.n194 VSUBS 0.007163f
C235 B.n195 VSUBS 0.007163f
C236 B.n196 VSUBS 0.007163f
C237 B.n197 VSUBS 0.007163f
C238 B.n198 VSUBS 0.007163f
C239 B.n199 VSUBS 0.007163f
C240 B.n200 VSUBS 0.007163f
C241 B.n201 VSUBS 0.007163f
C242 B.n202 VSUBS 0.007163f
C243 B.n203 VSUBS 0.007163f
C244 B.n204 VSUBS 0.007163f
C245 B.n205 VSUBS 0.007163f
C246 B.n206 VSUBS 0.007163f
C247 B.n207 VSUBS 0.007163f
C248 B.n208 VSUBS 0.007163f
C249 B.n209 VSUBS 0.007163f
C250 B.n210 VSUBS 0.007163f
C251 B.n211 VSUBS 0.007163f
C252 B.n212 VSUBS 0.007163f
C253 B.n213 VSUBS 0.007163f
C254 B.n214 VSUBS 0.007163f
C255 B.n215 VSUBS 0.007163f
C256 B.n216 VSUBS 0.007163f
C257 B.n217 VSUBS 0.007163f
C258 B.n218 VSUBS 0.007163f
C259 B.n219 VSUBS 0.007163f
C260 B.n220 VSUBS 0.007163f
C261 B.n221 VSUBS 0.007163f
C262 B.n222 VSUBS 0.007163f
C263 B.n223 VSUBS 0.007163f
C264 B.n224 VSUBS 0.007163f
C265 B.n225 VSUBS 0.007163f
C266 B.n226 VSUBS 0.007163f
C267 B.n227 VSUBS 0.007163f
C268 B.n228 VSUBS 0.007163f
C269 B.n229 VSUBS 0.007163f
C270 B.n230 VSUBS 0.007163f
C271 B.n231 VSUBS 0.007163f
C272 B.n232 VSUBS 0.007163f
C273 B.n233 VSUBS 0.007163f
C274 B.n234 VSUBS 0.007163f
C275 B.n235 VSUBS 0.007163f
C276 B.n236 VSUBS 0.007163f
C277 B.n237 VSUBS 0.007163f
C278 B.n238 VSUBS 0.007163f
C279 B.n239 VSUBS 0.007163f
C280 B.n240 VSUBS 0.007163f
C281 B.n241 VSUBS 0.007163f
C282 B.n242 VSUBS 0.007163f
C283 B.n243 VSUBS 0.007163f
C284 B.n244 VSUBS 0.007163f
C285 B.n245 VSUBS 0.007163f
C286 B.n246 VSUBS 0.007163f
C287 B.n247 VSUBS 0.007163f
C288 B.n248 VSUBS 0.007163f
C289 B.n249 VSUBS 0.007163f
C290 B.n250 VSUBS 0.007163f
C291 B.n251 VSUBS 0.007163f
C292 B.n252 VSUBS 0.007163f
C293 B.n253 VSUBS 0.007163f
C294 B.n254 VSUBS 0.007163f
C295 B.n255 VSUBS 0.007163f
C296 B.n256 VSUBS 0.007163f
C297 B.n257 VSUBS 0.007163f
C298 B.n258 VSUBS 0.016673f
C299 B.n259 VSUBS 0.017457f
C300 B.n260 VSUBS 0.017457f
C301 B.n261 VSUBS 0.007163f
C302 B.n262 VSUBS 0.007163f
C303 B.n263 VSUBS 0.007163f
C304 B.n264 VSUBS 0.007163f
C305 B.n265 VSUBS 0.007163f
C306 B.n266 VSUBS 0.007163f
C307 B.n267 VSUBS 0.007163f
C308 B.n268 VSUBS 0.007163f
C309 B.n269 VSUBS 0.007163f
C310 B.n270 VSUBS 0.007163f
C311 B.n271 VSUBS 0.007163f
C312 B.n272 VSUBS 0.007163f
C313 B.n273 VSUBS 0.007163f
C314 B.n274 VSUBS 0.007163f
C315 B.n275 VSUBS 0.007163f
C316 B.n276 VSUBS 0.007163f
C317 B.n277 VSUBS 0.007163f
C318 B.n278 VSUBS 0.007163f
C319 B.n279 VSUBS 0.007163f
C320 B.n280 VSUBS 0.007163f
C321 B.n281 VSUBS 0.007163f
C322 B.n282 VSUBS 0.007163f
C323 B.n283 VSUBS 0.007163f
C324 B.n284 VSUBS 0.007163f
C325 B.n285 VSUBS 0.007163f
C326 B.n286 VSUBS 0.007163f
C327 B.n287 VSUBS 0.007163f
C328 B.n288 VSUBS 0.007163f
C329 B.n289 VSUBS 0.007163f
C330 B.n290 VSUBS 0.007163f
C331 B.n291 VSUBS 0.007163f
C332 B.n292 VSUBS 0.007163f
C333 B.n293 VSUBS 0.007163f
C334 B.n294 VSUBS 0.007163f
C335 B.n295 VSUBS 0.007163f
C336 B.n296 VSUBS 0.007163f
C337 B.n297 VSUBS 0.007163f
C338 B.n298 VSUBS 0.007163f
C339 B.n299 VSUBS 0.007163f
C340 B.n300 VSUBS 0.007163f
C341 B.n301 VSUBS 0.007163f
C342 B.n302 VSUBS 0.007163f
C343 B.n303 VSUBS 0.007163f
C344 B.n304 VSUBS 0.007163f
C345 B.n305 VSUBS 0.007163f
C346 B.n306 VSUBS 0.007163f
C347 B.n307 VSUBS 0.007163f
C348 B.n308 VSUBS 0.007163f
C349 B.n309 VSUBS 0.007163f
C350 B.n310 VSUBS 0.007163f
C351 B.n311 VSUBS 0.007163f
C352 B.n312 VSUBS 0.004951f
C353 B.n313 VSUBS 0.016596f
C354 B.n314 VSUBS 0.005794f
C355 B.n315 VSUBS 0.007163f
C356 B.n316 VSUBS 0.007163f
C357 B.n317 VSUBS 0.007163f
C358 B.n318 VSUBS 0.007163f
C359 B.n319 VSUBS 0.007163f
C360 B.n320 VSUBS 0.007163f
C361 B.n321 VSUBS 0.007163f
C362 B.n322 VSUBS 0.007163f
C363 B.n323 VSUBS 0.007163f
C364 B.n324 VSUBS 0.007163f
C365 B.n325 VSUBS 0.007163f
C366 B.n326 VSUBS 0.005794f
C367 B.n327 VSUBS 0.007163f
C368 B.n328 VSUBS 0.007163f
C369 B.n329 VSUBS 0.004951f
C370 B.n330 VSUBS 0.007163f
C371 B.n331 VSUBS 0.007163f
C372 B.n332 VSUBS 0.007163f
C373 B.n333 VSUBS 0.007163f
C374 B.n334 VSUBS 0.007163f
C375 B.n335 VSUBS 0.007163f
C376 B.n336 VSUBS 0.007163f
C377 B.n337 VSUBS 0.007163f
C378 B.n338 VSUBS 0.007163f
C379 B.n339 VSUBS 0.007163f
C380 B.n340 VSUBS 0.007163f
C381 B.n341 VSUBS 0.007163f
C382 B.n342 VSUBS 0.007163f
C383 B.n343 VSUBS 0.007163f
C384 B.n344 VSUBS 0.007163f
C385 B.n345 VSUBS 0.007163f
C386 B.n346 VSUBS 0.007163f
C387 B.n347 VSUBS 0.007163f
C388 B.n348 VSUBS 0.007163f
C389 B.n349 VSUBS 0.007163f
C390 B.n350 VSUBS 0.007163f
C391 B.n351 VSUBS 0.007163f
C392 B.n352 VSUBS 0.007163f
C393 B.n353 VSUBS 0.007163f
C394 B.n354 VSUBS 0.007163f
C395 B.n355 VSUBS 0.007163f
C396 B.n356 VSUBS 0.007163f
C397 B.n357 VSUBS 0.007163f
C398 B.n358 VSUBS 0.007163f
C399 B.n359 VSUBS 0.007163f
C400 B.n360 VSUBS 0.007163f
C401 B.n361 VSUBS 0.007163f
C402 B.n362 VSUBS 0.007163f
C403 B.n363 VSUBS 0.007163f
C404 B.n364 VSUBS 0.007163f
C405 B.n365 VSUBS 0.007163f
C406 B.n366 VSUBS 0.007163f
C407 B.n367 VSUBS 0.007163f
C408 B.n368 VSUBS 0.007163f
C409 B.n369 VSUBS 0.007163f
C410 B.n370 VSUBS 0.007163f
C411 B.n371 VSUBS 0.007163f
C412 B.n372 VSUBS 0.007163f
C413 B.n373 VSUBS 0.007163f
C414 B.n374 VSUBS 0.007163f
C415 B.n375 VSUBS 0.007163f
C416 B.n376 VSUBS 0.007163f
C417 B.n377 VSUBS 0.007163f
C418 B.n378 VSUBS 0.007163f
C419 B.n379 VSUBS 0.007163f
C420 B.n380 VSUBS 0.007163f
C421 B.n381 VSUBS 0.017457f
C422 B.n382 VSUBS 0.016673f
C423 B.n383 VSUBS 0.017497f
C424 B.n384 VSUBS 0.007163f
C425 B.n385 VSUBS 0.007163f
C426 B.n386 VSUBS 0.007163f
C427 B.n387 VSUBS 0.007163f
C428 B.n388 VSUBS 0.007163f
C429 B.n389 VSUBS 0.007163f
C430 B.n390 VSUBS 0.007163f
C431 B.n391 VSUBS 0.007163f
C432 B.n392 VSUBS 0.007163f
C433 B.n393 VSUBS 0.007163f
C434 B.n394 VSUBS 0.007163f
C435 B.n395 VSUBS 0.007163f
C436 B.n396 VSUBS 0.007163f
C437 B.n397 VSUBS 0.007163f
C438 B.n398 VSUBS 0.007163f
C439 B.n399 VSUBS 0.007163f
C440 B.n400 VSUBS 0.007163f
C441 B.n401 VSUBS 0.007163f
C442 B.n402 VSUBS 0.007163f
C443 B.n403 VSUBS 0.007163f
C444 B.n404 VSUBS 0.007163f
C445 B.n405 VSUBS 0.007163f
C446 B.n406 VSUBS 0.007163f
C447 B.n407 VSUBS 0.007163f
C448 B.n408 VSUBS 0.007163f
C449 B.n409 VSUBS 0.007163f
C450 B.n410 VSUBS 0.007163f
C451 B.n411 VSUBS 0.007163f
C452 B.n412 VSUBS 0.007163f
C453 B.n413 VSUBS 0.007163f
C454 B.n414 VSUBS 0.007163f
C455 B.n415 VSUBS 0.007163f
C456 B.n416 VSUBS 0.007163f
C457 B.n417 VSUBS 0.007163f
C458 B.n418 VSUBS 0.007163f
C459 B.n419 VSUBS 0.007163f
C460 B.n420 VSUBS 0.007163f
C461 B.n421 VSUBS 0.007163f
C462 B.n422 VSUBS 0.007163f
C463 B.n423 VSUBS 0.007163f
C464 B.n424 VSUBS 0.007163f
C465 B.n425 VSUBS 0.007163f
C466 B.n426 VSUBS 0.007163f
C467 B.n427 VSUBS 0.007163f
C468 B.n428 VSUBS 0.007163f
C469 B.n429 VSUBS 0.007163f
C470 B.n430 VSUBS 0.007163f
C471 B.n431 VSUBS 0.007163f
C472 B.n432 VSUBS 0.007163f
C473 B.n433 VSUBS 0.007163f
C474 B.n434 VSUBS 0.007163f
C475 B.n435 VSUBS 0.007163f
C476 B.n436 VSUBS 0.007163f
C477 B.n437 VSUBS 0.007163f
C478 B.n438 VSUBS 0.007163f
C479 B.n439 VSUBS 0.007163f
C480 B.n440 VSUBS 0.007163f
C481 B.n441 VSUBS 0.007163f
C482 B.n442 VSUBS 0.007163f
C483 B.n443 VSUBS 0.007163f
C484 B.n444 VSUBS 0.007163f
C485 B.n445 VSUBS 0.007163f
C486 B.n446 VSUBS 0.007163f
C487 B.n447 VSUBS 0.007163f
C488 B.n448 VSUBS 0.007163f
C489 B.n449 VSUBS 0.007163f
C490 B.n450 VSUBS 0.007163f
C491 B.n451 VSUBS 0.007163f
C492 B.n452 VSUBS 0.007163f
C493 B.n453 VSUBS 0.007163f
C494 B.n454 VSUBS 0.007163f
C495 B.n455 VSUBS 0.007163f
C496 B.n456 VSUBS 0.007163f
C497 B.n457 VSUBS 0.007163f
C498 B.n458 VSUBS 0.007163f
C499 B.n459 VSUBS 0.007163f
C500 B.n460 VSUBS 0.007163f
C501 B.n461 VSUBS 0.007163f
C502 B.n462 VSUBS 0.007163f
C503 B.n463 VSUBS 0.007163f
C504 B.n464 VSUBS 0.007163f
C505 B.n465 VSUBS 0.007163f
C506 B.n466 VSUBS 0.007163f
C507 B.n467 VSUBS 0.007163f
C508 B.n468 VSUBS 0.007163f
C509 B.n469 VSUBS 0.007163f
C510 B.n470 VSUBS 0.007163f
C511 B.n471 VSUBS 0.007163f
C512 B.n472 VSUBS 0.007163f
C513 B.n473 VSUBS 0.007163f
C514 B.n474 VSUBS 0.007163f
C515 B.n475 VSUBS 0.007163f
C516 B.n476 VSUBS 0.007163f
C517 B.n477 VSUBS 0.007163f
C518 B.n478 VSUBS 0.007163f
C519 B.n479 VSUBS 0.007163f
C520 B.n480 VSUBS 0.007163f
C521 B.n481 VSUBS 0.007163f
C522 B.n482 VSUBS 0.007163f
C523 B.n483 VSUBS 0.007163f
C524 B.n484 VSUBS 0.007163f
C525 B.n485 VSUBS 0.007163f
C526 B.n486 VSUBS 0.007163f
C527 B.n487 VSUBS 0.007163f
C528 B.n488 VSUBS 0.007163f
C529 B.n489 VSUBS 0.007163f
C530 B.n490 VSUBS 0.007163f
C531 B.n491 VSUBS 0.007163f
C532 B.n492 VSUBS 0.007163f
C533 B.n493 VSUBS 0.007163f
C534 B.n494 VSUBS 0.007163f
C535 B.n495 VSUBS 0.007163f
C536 B.n496 VSUBS 0.007163f
C537 B.n497 VSUBS 0.007163f
C538 B.n498 VSUBS 0.007163f
C539 B.n499 VSUBS 0.007163f
C540 B.n500 VSUBS 0.007163f
C541 B.n501 VSUBS 0.007163f
C542 B.n502 VSUBS 0.007163f
C543 B.n503 VSUBS 0.007163f
C544 B.n504 VSUBS 0.007163f
C545 B.n505 VSUBS 0.007163f
C546 B.n506 VSUBS 0.007163f
C547 B.n507 VSUBS 0.007163f
C548 B.n508 VSUBS 0.007163f
C549 B.n509 VSUBS 0.007163f
C550 B.n510 VSUBS 0.007163f
C551 B.n511 VSUBS 0.007163f
C552 B.n512 VSUBS 0.007163f
C553 B.n513 VSUBS 0.007163f
C554 B.n514 VSUBS 0.007163f
C555 B.n515 VSUBS 0.007163f
C556 B.n516 VSUBS 0.007163f
C557 B.n517 VSUBS 0.007163f
C558 B.n518 VSUBS 0.007163f
C559 B.n519 VSUBS 0.007163f
C560 B.n520 VSUBS 0.007163f
C561 B.n521 VSUBS 0.007163f
C562 B.n522 VSUBS 0.007163f
C563 B.n523 VSUBS 0.007163f
C564 B.n524 VSUBS 0.007163f
C565 B.n525 VSUBS 0.007163f
C566 B.n526 VSUBS 0.007163f
C567 B.n527 VSUBS 0.007163f
C568 B.n528 VSUBS 0.016673f
C569 B.n529 VSUBS 0.017457f
C570 B.n530 VSUBS 0.017457f
C571 B.n531 VSUBS 0.007163f
C572 B.n532 VSUBS 0.007163f
C573 B.n533 VSUBS 0.007163f
C574 B.n534 VSUBS 0.007163f
C575 B.n535 VSUBS 0.007163f
C576 B.n536 VSUBS 0.007163f
C577 B.n537 VSUBS 0.007163f
C578 B.n538 VSUBS 0.007163f
C579 B.n539 VSUBS 0.007163f
C580 B.n540 VSUBS 0.007163f
C581 B.n541 VSUBS 0.007163f
C582 B.n542 VSUBS 0.007163f
C583 B.n543 VSUBS 0.007163f
C584 B.n544 VSUBS 0.007163f
C585 B.n545 VSUBS 0.007163f
C586 B.n546 VSUBS 0.007163f
C587 B.n547 VSUBS 0.007163f
C588 B.n548 VSUBS 0.007163f
C589 B.n549 VSUBS 0.007163f
C590 B.n550 VSUBS 0.007163f
C591 B.n551 VSUBS 0.007163f
C592 B.n552 VSUBS 0.007163f
C593 B.n553 VSUBS 0.007163f
C594 B.n554 VSUBS 0.007163f
C595 B.n555 VSUBS 0.007163f
C596 B.n556 VSUBS 0.007163f
C597 B.n557 VSUBS 0.007163f
C598 B.n558 VSUBS 0.007163f
C599 B.n559 VSUBS 0.007163f
C600 B.n560 VSUBS 0.007163f
C601 B.n561 VSUBS 0.007163f
C602 B.n562 VSUBS 0.007163f
C603 B.n563 VSUBS 0.007163f
C604 B.n564 VSUBS 0.007163f
C605 B.n565 VSUBS 0.007163f
C606 B.n566 VSUBS 0.007163f
C607 B.n567 VSUBS 0.007163f
C608 B.n568 VSUBS 0.007163f
C609 B.n569 VSUBS 0.007163f
C610 B.n570 VSUBS 0.007163f
C611 B.n571 VSUBS 0.007163f
C612 B.n572 VSUBS 0.007163f
C613 B.n573 VSUBS 0.007163f
C614 B.n574 VSUBS 0.007163f
C615 B.n575 VSUBS 0.007163f
C616 B.n576 VSUBS 0.007163f
C617 B.n577 VSUBS 0.007163f
C618 B.n578 VSUBS 0.007163f
C619 B.n579 VSUBS 0.007163f
C620 B.n580 VSUBS 0.007163f
C621 B.n581 VSUBS 0.007163f
C622 B.n582 VSUBS 0.004951f
C623 B.n583 VSUBS 0.016596f
C624 B.n584 VSUBS 0.005794f
C625 B.n585 VSUBS 0.007163f
C626 B.n586 VSUBS 0.007163f
C627 B.n587 VSUBS 0.007163f
C628 B.n588 VSUBS 0.007163f
C629 B.n589 VSUBS 0.007163f
C630 B.n590 VSUBS 0.007163f
C631 B.n591 VSUBS 0.007163f
C632 B.n592 VSUBS 0.007163f
C633 B.n593 VSUBS 0.007163f
C634 B.n594 VSUBS 0.007163f
C635 B.n595 VSUBS 0.007163f
C636 B.n596 VSUBS 0.005794f
C637 B.n597 VSUBS 0.007163f
C638 B.n598 VSUBS 0.007163f
C639 B.n599 VSUBS 0.004951f
C640 B.n600 VSUBS 0.007163f
C641 B.n601 VSUBS 0.007163f
C642 B.n602 VSUBS 0.007163f
C643 B.n603 VSUBS 0.007163f
C644 B.n604 VSUBS 0.007163f
C645 B.n605 VSUBS 0.007163f
C646 B.n606 VSUBS 0.007163f
C647 B.n607 VSUBS 0.007163f
C648 B.n608 VSUBS 0.007163f
C649 B.n609 VSUBS 0.007163f
C650 B.n610 VSUBS 0.007163f
C651 B.n611 VSUBS 0.007163f
C652 B.n612 VSUBS 0.007163f
C653 B.n613 VSUBS 0.007163f
C654 B.n614 VSUBS 0.007163f
C655 B.n615 VSUBS 0.007163f
C656 B.n616 VSUBS 0.007163f
C657 B.n617 VSUBS 0.007163f
C658 B.n618 VSUBS 0.007163f
C659 B.n619 VSUBS 0.007163f
C660 B.n620 VSUBS 0.007163f
C661 B.n621 VSUBS 0.007163f
C662 B.n622 VSUBS 0.007163f
C663 B.n623 VSUBS 0.007163f
C664 B.n624 VSUBS 0.007163f
C665 B.n625 VSUBS 0.007163f
C666 B.n626 VSUBS 0.007163f
C667 B.n627 VSUBS 0.007163f
C668 B.n628 VSUBS 0.007163f
C669 B.n629 VSUBS 0.007163f
C670 B.n630 VSUBS 0.007163f
C671 B.n631 VSUBS 0.007163f
C672 B.n632 VSUBS 0.007163f
C673 B.n633 VSUBS 0.007163f
C674 B.n634 VSUBS 0.007163f
C675 B.n635 VSUBS 0.007163f
C676 B.n636 VSUBS 0.007163f
C677 B.n637 VSUBS 0.007163f
C678 B.n638 VSUBS 0.007163f
C679 B.n639 VSUBS 0.007163f
C680 B.n640 VSUBS 0.007163f
C681 B.n641 VSUBS 0.007163f
C682 B.n642 VSUBS 0.007163f
C683 B.n643 VSUBS 0.007163f
C684 B.n644 VSUBS 0.007163f
C685 B.n645 VSUBS 0.007163f
C686 B.n646 VSUBS 0.007163f
C687 B.n647 VSUBS 0.007163f
C688 B.n648 VSUBS 0.007163f
C689 B.n649 VSUBS 0.007163f
C690 B.n650 VSUBS 0.007163f
C691 B.n651 VSUBS 0.017457f
C692 B.n652 VSUBS 0.016673f
C693 B.n653 VSUBS 0.016673f
C694 B.n654 VSUBS 0.007163f
C695 B.n655 VSUBS 0.007163f
C696 B.n656 VSUBS 0.007163f
C697 B.n657 VSUBS 0.007163f
C698 B.n658 VSUBS 0.007163f
C699 B.n659 VSUBS 0.007163f
C700 B.n660 VSUBS 0.007163f
C701 B.n661 VSUBS 0.007163f
C702 B.n662 VSUBS 0.007163f
C703 B.n663 VSUBS 0.007163f
C704 B.n664 VSUBS 0.007163f
C705 B.n665 VSUBS 0.007163f
C706 B.n666 VSUBS 0.007163f
C707 B.n667 VSUBS 0.007163f
C708 B.n668 VSUBS 0.007163f
C709 B.n669 VSUBS 0.007163f
C710 B.n670 VSUBS 0.007163f
C711 B.n671 VSUBS 0.007163f
C712 B.n672 VSUBS 0.007163f
C713 B.n673 VSUBS 0.007163f
C714 B.n674 VSUBS 0.007163f
C715 B.n675 VSUBS 0.007163f
C716 B.n676 VSUBS 0.007163f
C717 B.n677 VSUBS 0.007163f
C718 B.n678 VSUBS 0.007163f
C719 B.n679 VSUBS 0.007163f
C720 B.n680 VSUBS 0.007163f
C721 B.n681 VSUBS 0.007163f
C722 B.n682 VSUBS 0.007163f
C723 B.n683 VSUBS 0.007163f
C724 B.n684 VSUBS 0.007163f
C725 B.n685 VSUBS 0.007163f
C726 B.n686 VSUBS 0.007163f
C727 B.n687 VSUBS 0.007163f
C728 B.n688 VSUBS 0.007163f
C729 B.n689 VSUBS 0.007163f
C730 B.n690 VSUBS 0.007163f
C731 B.n691 VSUBS 0.007163f
C732 B.n692 VSUBS 0.007163f
C733 B.n693 VSUBS 0.007163f
C734 B.n694 VSUBS 0.007163f
C735 B.n695 VSUBS 0.007163f
C736 B.n696 VSUBS 0.007163f
C737 B.n697 VSUBS 0.007163f
C738 B.n698 VSUBS 0.007163f
C739 B.n699 VSUBS 0.007163f
C740 B.n700 VSUBS 0.007163f
C741 B.n701 VSUBS 0.007163f
C742 B.n702 VSUBS 0.007163f
C743 B.n703 VSUBS 0.007163f
C744 B.n704 VSUBS 0.007163f
C745 B.n705 VSUBS 0.007163f
C746 B.n706 VSUBS 0.007163f
C747 B.n707 VSUBS 0.007163f
C748 B.n708 VSUBS 0.007163f
C749 B.n709 VSUBS 0.007163f
C750 B.n710 VSUBS 0.007163f
C751 B.n711 VSUBS 0.007163f
C752 B.n712 VSUBS 0.007163f
C753 B.n713 VSUBS 0.007163f
C754 B.n714 VSUBS 0.007163f
C755 B.n715 VSUBS 0.007163f
C756 B.n716 VSUBS 0.007163f
C757 B.n717 VSUBS 0.007163f
C758 B.n718 VSUBS 0.007163f
C759 B.n719 VSUBS 0.007163f
C760 B.n720 VSUBS 0.007163f
C761 B.n721 VSUBS 0.007163f
C762 B.n722 VSUBS 0.007163f
C763 B.n723 VSUBS 0.009347f
C764 B.n724 VSUBS 0.009957f
C765 B.n725 VSUBS 0.019801f
C766 VDD1.t7 VSUBS 0.196142f
C767 VDD1.t6 VSUBS 0.196142f
C768 VDD1.n0 VSUBS 1.49557f
C769 VDD1.t1 VSUBS 0.196142f
C770 VDD1.t5 VSUBS 0.196142f
C771 VDD1.n1 VSUBS 1.4944f
C772 VDD1.t0 VSUBS 0.196142f
C773 VDD1.t4 VSUBS 0.196142f
C774 VDD1.n2 VSUBS 1.4944f
C775 VDD1.n3 VSUBS 3.55622f
C776 VDD1.t2 VSUBS 0.196142f
C777 VDD1.t3 VSUBS 0.196142f
C778 VDD1.n4 VSUBS 1.4839f
C779 VDD1.n5 VSUBS 2.98436f
C780 VP.n0 VSUBS 0.043342f
C781 VP.t3 VSUBS 2.15747f
C782 VP.n1 VSUBS 0.047991f
C783 VP.n2 VSUBS 0.032875f
C784 VP.t7 VSUBS 2.15747f
C785 VP.n3 VSUBS 0.774176f
C786 VP.n4 VSUBS 0.032875f
C787 VP.n5 VSUBS 0.065338f
C788 VP.n6 VSUBS 0.032875f
C789 VP.t2 VSUBS 2.15747f
C790 VP.n7 VSUBS 0.047991f
C791 VP.n8 VSUBS 0.032875f
C792 VP.t6 VSUBS 2.15747f
C793 VP.n9 VSUBS 0.8697f
C794 VP.n10 VSUBS 0.043342f
C795 VP.t4 VSUBS 2.15747f
C796 VP.n11 VSUBS 0.047991f
C797 VP.n12 VSUBS 0.032875f
C798 VP.t5 VSUBS 2.15747f
C799 VP.n13 VSUBS 0.774176f
C800 VP.n14 VSUBS 0.032875f
C801 VP.n15 VSUBS 0.065338f
C802 VP.t0 VSUBS 2.39447f
C803 VP.n16 VSUBS 0.847251f
C804 VP.t1 VSUBS 2.15747f
C805 VP.n17 VSUBS 0.873115f
C806 VP.n18 VSUBS 0.053707f
C807 VP.n19 VSUBS 0.311253f
C808 VP.n20 VSUBS 0.032875f
C809 VP.n21 VSUBS 0.032875f
C810 VP.n22 VSUBS 0.026576f
C811 VP.n23 VSUBS 0.065338f
C812 VP.n24 VSUBS 0.053707f
C813 VP.n25 VSUBS 0.032875f
C814 VP.n26 VSUBS 0.032875f
C815 VP.n27 VSUBS 0.038582f
C816 VP.n28 VSUBS 0.06127f
C817 VP.n29 VSUBS 0.047991f
C818 VP.n30 VSUBS 0.032875f
C819 VP.n31 VSUBS 0.032875f
C820 VP.n32 VSUBS 0.032875f
C821 VP.n33 VSUBS 0.06127f
C822 VP.n34 VSUBS 0.038582f
C823 VP.n35 VSUBS 0.8697f
C824 VP.n36 VSUBS 1.74586f
C825 VP.n37 VSUBS 1.77024f
C826 VP.n38 VSUBS 0.043342f
C827 VP.n39 VSUBS 0.038582f
C828 VP.n40 VSUBS 0.06127f
C829 VP.n41 VSUBS 0.047991f
C830 VP.n42 VSUBS 0.032875f
C831 VP.n43 VSUBS 0.032875f
C832 VP.n44 VSUBS 0.032875f
C833 VP.n45 VSUBS 0.06127f
C834 VP.n46 VSUBS 0.038582f
C835 VP.n47 VSUBS 0.774176f
C836 VP.n48 VSUBS 0.053707f
C837 VP.n49 VSUBS 0.032875f
C838 VP.n50 VSUBS 0.032875f
C839 VP.n51 VSUBS 0.032875f
C840 VP.n52 VSUBS 0.026576f
C841 VP.n53 VSUBS 0.065338f
C842 VP.n54 VSUBS 0.053707f
C843 VP.n55 VSUBS 0.032875f
C844 VP.n56 VSUBS 0.032875f
C845 VP.n57 VSUBS 0.038582f
C846 VP.n58 VSUBS 0.06127f
C847 VP.n59 VSUBS 0.047991f
C848 VP.n60 VSUBS 0.032875f
C849 VP.n61 VSUBS 0.032875f
C850 VP.n62 VSUBS 0.032875f
C851 VP.n63 VSUBS 0.06127f
C852 VP.n64 VSUBS 0.038582f
C853 VP.n65 VSUBS 0.8697f
C854 VP.n66 VSUBS 0.05439f
C855 VDD2.t1 VSUBS 0.192085f
C856 VDD2.t7 VSUBS 0.192085f
C857 VDD2.n0 VSUBS 1.46348f
C858 VDD2.t2 VSUBS 0.192085f
C859 VDD2.t0 VSUBS 0.192085f
C860 VDD2.n1 VSUBS 1.46348f
C861 VDD2.n2 VSUBS 3.4319f
C862 VDD2.t4 VSUBS 0.192085f
C863 VDD2.t6 VSUBS 0.192085f
C864 VDD2.n3 VSUBS 1.45321f
C865 VDD2.n4 VSUBS 2.89278f
C866 VDD2.t3 VSUBS 0.192085f
C867 VDD2.t5 VSUBS 0.192085f
C868 VDD2.n5 VSUBS 1.46344f
C869 VTAIL.t8 VSUBS 0.203953f
C870 VTAIL.t11 VSUBS 0.203953f
C871 VTAIL.n0 VSUBS 1.41851f
C872 VTAIL.n1 VSUBS 0.754497f
C873 VTAIL.n2 VSUBS 0.027458f
C874 VTAIL.n3 VSUBS 0.025784f
C875 VTAIL.n4 VSUBS 0.013855f
C876 VTAIL.n5 VSUBS 0.032748f
C877 VTAIL.n6 VSUBS 0.01467f
C878 VTAIL.n7 VSUBS 0.025784f
C879 VTAIL.n8 VSUBS 0.014262f
C880 VTAIL.n9 VSUBS 0.032748f
C881 VTAIL.n10 VSUBS 0.01467f
C882 VTAIL.n11 VSUBS 0.025784f
C883 VTAIL.n12 VSUBS 0.013855f
C884 VTAIL.n13 VSUBS 0.032748f
C885 VTAIL.n14 VSUBS 0.01467f
C886 VTAIL.n15 VSUBS 0.025784f
C887 VTAIL.n16 VSUBS 0.013855f
C888 VTAIL.n17 VSUBS 0.024561f
C889 VTAIL.n18 VSUBS 0.024635f
C890 VTAIL.t9 VSUBS 0.070415f
C891 VTAIL.n19 VSUBS 0.179878f
C892 VTAIL.n20 VSUBS 1.04197f
C893 VTAIL.n21 VSUBS 0.013855f
C894 VTAIL.n22 VSUBS 0.01467f
C895 VTAIL.n23 VSUBS 0.032748f
C896 VTAIL.n24 VSUBS 0.032748f
C897 VTAIL.n25 VSUBS 0.01467f
C898 VTAIL.n26 VSUBS 0.013855f
C899 VTAIL.n27 VSUBS 0.025784f
C900 VTAIL.n28 VSUBS 0.025784f
C901 VTAIL.n29 VSUBS 0.013855f
C902 VTAIL.n30 VSUBS 0.01467f
C903 VTAIL.n31 VSUBS 0.032748f
C904 VTAIL.n32 VSUBS 0.032748f
C905 VTAIL.n33 VSUBS 0.01467f
C906 VTAIL.n34 VSUBS 0.013855f
C907 VTAIL.n35 VSUBS 0.025784f
C908 VTAIL.n36 VSUBS 0.025784f
C909 VTAIL.n37 VSUBS 0.013855f
C910 VTAIL.n38 VSUBS 0.013855f
C911 VTAIL.n39 VSUBS 0.01467f
C912 VTAIL.n40 VSUBS 0.032748f
C913 VTAIL.n41 VSUBS 0.032748f
C914 VTAIL.n42 VSUBS 0.032748f
C915 VTAIL.n43 VSUBS 0.014262f
C916 VTAIL.n44 VSUBS 0.013855f
C917 VTAIL.n45 VSUBS 0.025784f
C918 VTAIL.n46 VSUBS 0.025784f
C919 VTAIL.n47 VSUBS 0.013855f
C920 VTAIL.n48 VSUBS 0.01467f
C921 VTAIL.n49 VSUBS 0.032748f
C922 VTAIL.n50 VSUBS 0.076306f
C923 VTAIL.n51 VSUBS 0.01467f
C924 VTAIL.n52 VSUBS 0.013855f
C925 VTAIL.n53 VSUBS 0.061359f
C926 VTAIL.n54 VSUBS 0.038295f
C927 VTAIL.n55 VSUBS 0.259007f
C928 VTAIL.n56 VSUBS 0.027458f
C929 VTAIL.n57 VSUBS 0.025784f
C930 VTAIL.n58 VSUBS 0.013855f
C931 VTAIL.n59 VSUBS 0.032748f
C932 VTAIL.n60 VSUBS 0.01467f
C933 VTAIL.n61 VSUBS 0.025784f
C934 VTAIL.n62 VSUBS 0.014262f
C935 VTAIL.n63 VSUBS 0.032748f
C936 VTAIL.n64 VSUBS 0.01467f
C937 VTAIL.n65 VSUBS 0.025784f
C938 VTAIL.n66 VSUBS 0.013855f
C939 VTAIL.n67 VSUBS 0.032748f
C940 VTAIL.n68 VSUBS 0.01467f
C941 VTAIL.n69 VSUBS 0.025784f
C942 VTAIL.n70 VSUBS 0.013855f
C943 VTAIL.n71 VSUBS 0.024561f
C944 VTAIL.n72 VSUBS 0.024635f
C945 VTAIL.t3 VSUBS 0.070415f
C946 VTAIL.n73 VSUBS 0.179878f
C947 VTAIL.n74 VSUBS 1.04197f
C948 VTAIL.n75 VSUBS 0.013855f
C949 VTAIL.n76 VSUBS 0.01467f
C950 VTAIL.n77 VSUBS 0.032748f
C951 VTAIL.n78 VSUBS 0.032748f
C952 VTAIL.n79 VSUBS 0.01467f
C953 VTAIL.n80 VSUBS 0.013855f
C954 VTAIL.n81 VSUBS 0.025784f
C955 VTAIL.n82 VSUBS 0.025784f
C956 VTAIL.n83 VSUBS 0.013855f
C957 VTAIL.n84 VSUBS 0.01467f
C958 VTAIL.n85 VSUBS 0.032748f
C959 VTAIL.n86 VSUBS 0.032748f
C960 VTAIL.n87 VSUBS 0.01467f
C961 VTAIL.n88 VSUBS 0.013855f
C962 VTAIL.n89 VSUBS 0.025784f
C963 VTAIL.n90 VSUBS 0.025784f
C964 VTAIL.n91 VSUBS 0.013855f
C965 VTAIL.n92 VSUBS 0.013855f
C966 VTAIL.n93 VSUBS 0.01467f
C967 VTAIL.n94 VSUBS 0.032748f
C968 VTAIL.n95 VSUBS 0.032748f
C969 VTAIL.n96 VSUBS 0.032748f
C970 VTAIL.n97 VSUBS 0.014262f
C971 VTAIL.n98 VSUBS 0.013855f
C972 VTAIL.n99 VSUBS 0.025784f
C973 VTAIL.n100 VSUBS 0.025784f
C974 VTAIL.n101 VSUBS 0.013855f
C975 VTAIL.n102 VSUBS 0.01467f
C976 VTAIL.n103 VSUBS 0.032748f
C977 VTAIL.n104 VSUBS 0.076306f
C978 VTAIL.n105 VSUBS 0.01467f
C979 VTAIL.n106 VSUBS 0.013855f
C980 VTAIL.n107 VSUBS 0.061359f
C981 VTAIL.n108 VSUBS 0.038295f
C982 VTAIL.n109 VSUBS 0.259007f
C983 VTAIL.t2 VSUBS 0.203953f
C984 VTAIL.t7 VSUBS 0.203953f
C985 VTAIL.n110 VSUBS 1.41851f
C986 VTAIL.n111 VSUBS 0.946621f
C987 VTAIL.n112 VSUBS 0.027458f
C988 VTAIL.n113 VSUBS 0.025784f
C989 VTAIL.n114 VSUBS 0.013855f
C990 VTAIL.n115 VSUBS 0.032748f
C991 VTAIL.n116 VSUBS 0.01467f
C992 VTAIL.n117 VSUBS 0.025784f
C993 VTAIL.n118 VSUBS 0.014262f
C994 VTAIL.n119 VSUBS 0.032748f
C995 VTAIL.n120 VSUBS 0.01467f
C996 VTAIL.n121 VSUBS 0.025784f
C997 VTAIL.n122 VSUBS 0.013855f
C998 VTAIL.n123 VSUBS 0.032748f
C999 VTAIL.n124 VSUBS 0.01467f
C1000 VTAIL.n125 VSUBS 0.025784f
C1001 VTAIL.n126 VSUBS 0.013855f
C1002 VTAIL.n127 VSUBS 0.024561f
C1003 VTAIL.n128 VSUBS 0.024635f
C1004 VTAIL.t4 VSUBS 0.070415f
C1005 VTAIL.n129 VSUBS 0.179878f
C1006 VTAIL.n130 VSUBS 1.04197f
C1007 VTAIL.n131 VSUBS 0.013855f
C1008 VTAIL.n132 VSUBS 0.01467f
C1009 VTAIL.n133 VSUBS 0.032748f
C1010 VTAIL.n134 VSUBS 0.032748f
C1011 VTAIL.n135 VSUBS 0.01467f
C1012 VTAIL.n136 VSUBS 0.013855f
C1013 VTAIL.n137 VSUBS 0.025784f
C1014 VTAIL.n138 VSUBS 0.025784f
C1015 VTAIL.n139 VSUBS 0.013855f
C1016 VTAIL.n140 VSUBS 0.01467f
C1017 VTAIL.n141 VSUBS 0.032748f
C1018 VTAIL.n142 VSUBS 0.032748f
C1019 VTAIL.n143 VSUBS 0.01467f
C1020 VTAIL.n144 VSUBS 0.013855f
C1021 VTAIL.n145 VSUBS 0.025784f
C1022 VTAIL.n146 VSUBS 0.025784f
C1023 VTAIL.n147 VSUBS 0.013855f
C1024 VTAIL.n148 VSUBS 0.013855f
C1025 VTAIL.n149 VSUBS 0.01467f
C1026 VTAIL.n150 VSUBS 0.032748f
C1027 VTAIL.n151 VSUBS 0.032748f
C1028 VTAIL.n152 VSUBS 0.032748f
C1029 VTAIL.n153 VSUBS 0.014262f
C1030 VTAIL.n154 VSUBS 0.013855f
C1031 VTAIL.n155 VSUBS 0.025784f
C1032 VTAIL.n156 VSUBS 0.025784f
C1033 VTAIL.n157 VSUBS 0.013855f
C1034 VTAIL.n158 VSUBS 0.01467f
C1035 VTAIL.n159 VSUBS 0.032748f
C1036 VTAIL.n160 VSUBS 0.076306f
C1037 VTAIL.n161 VSUBS 0.01467f
C1038 VTAIL.n162 VSUBS 0.013855f
C1039 VTAIL.n163 VSUBS 0.061359f
C1040 VTAIL.n164 VSUBS 0.038295f
C1041 VTAIL.n165 VSUBS 1.4841f
C1042 VTAIL.n166 VSUBS 0.027458f
C1043 VTAIL.n167 VSUBS 0.025784f
C1044 VTAIL.n168 VSUBS 0.013855f
C1045 VTAIL.n169 VSUBS 0.032748f
C1046 VTAIL.n170 VSUBS 0.01467f
C1047 VTAIL.n171 VSUBS 0.025784f
C1048 VTAIL.n172 VSUBS 0.014262f
C1049 VTAIL.n173 VSUBS 0.032748f
C1050 VTAIL.n174 VSUBS 0.013855f
C1051 VTAIL.n175 VSUBS 0.01467f
C1052 VTAIL.n176 VSUBS 0.025784f
C1053 VTAIL.n177 VSUBS 0.013855f
C1054 VTAIL.n178 VSUBS 0.032748f
C1055 VTAIL.n179 VSUBS 0.01467f
C1056 VTAIL.n180 VSUBS 0.025784f
C1057 VTAIL.n181 VSUBS 0.013855f
C1058 VTAIL.n182 VSUBS 0.024561f
C1059 VTAIL.n183 VSUBS 0.024635f
C1060 VTAIL.t12 VSUBS 0.070415f
C1061 VTAIL.n184 VSUBS 0.179878f
C1062 VTAIL.n185 VSUBS 1.04197f
C1063 VTAIL.n186 VSUBS 0.013855f
C1064 VTAIL.n187 VSUBS 0.01467f
C1065 VTAIL.n188 VSUBS 0.032748f
C1066 VTAIL.n189 VSUBS 0.032748f
C1067 VTAIL.n190 VSUBS 0.01467f
C1068 VTAIL.n191 VSUBS 0.013855f
C1069 VTAIL.n192 VSUBS 0.025784f
C1070 VTAIL.n193 VSUBS 0.025784f
C1071 VTAIL.n194 VSUBS 0.013855f
C1072 VTAIL.n195 VSUBS 0.01467f
C1073 VTAIL.n196 VSUBS 0.032748f
C1074 VTAIL.n197 VSUBS 0.032748f
C1075 VTAIL.n198 VSUBS 0.01467f
C1076 VTAIL.n199 VSUBS 0.013855f
C1077 VTAIL.n200 VSUBS 0.025784f
C1078 VTAIL.n201 VSUBS 0.025784f
C1079 VTAIL.n202 VSUBS 0.013855f
C1080 VTAIL.n203 VSUBS 0.01467f
C1081 VTAIL.n204 VSUBS 0.032748f
C1082 VTAIL.n205 VSUBS 0.032748f
C1083 VTAIL.n206 VSUBS 0.032748f
C1084 VTAIL.n207 VSUBS 0.014262f
C1085 VTAIL.n208 VSUBS 0.013855f
C1086 VTAIL.n209 VSUBS 0.025784f
C1087 VTAIL.n210 VSUBS 0.025784f
C1088 VTAIL.n211 VSUBS 0.013855f
C1089 VTAIL.n212 VSUBS 0.01467f
C1090 VTAIL.n213 VSUBS 0.032748f
C1091 VTAIL.n214 VSUBS 0.076306f
C1092 VTAIL.n215 VSUBS 0.01467f
C1093 VTAIL.n216 VSUBS 0.013855f
C1094 VTAIL.n217 VSUBS 0.061359f
C1095 VTAIL.n218 VSUBS 0.038295f
C1096 VTAIL.n219 VSUBS 1.4841f
C1097 VTAIL.t10 VSUBS 0.203953f
C1098 VTAIL.t15 VSUBS 0.203953f
C1099 VTAIL.n220 VSUBS 1.41852f
C1100 VTAIL.n221 VSUBS 0.946611f
C1101 VTAIL.n222 VSUBS 0.027458f
C1102 VTAIL.n223 VSUBS 0.025784f
C1103 VTAIL.n224 VSUBS 0.013855f
C1104 VTAIL.n225 VSUBS 0.032748f
C1105 VTAIL.n226 VSUBS 0.01467f
C1106 VTAIL.n227 VSUBS 0.025784f
C1107 VTAIL.n228 VSUBS 0.014262f
C1108 VTAIL.n229 VSUBS 0.032748f
C1109 VTAIL.n230 VSUBS 0.013855f
C1110 VTAIL.n231 VSUBS 0.01467f
C1111 VTAIL.n232 VSUBS 0.025784f
C1112 VTAIL.n233 VSUBS 0.013855f
C1113 VTAIL.n234 VSUBS 0.032748f
C1114 VTAIL.n235 VSUBS 0.01467f
C1115 VTAIL.n236 VSUBS 0.025784f
C1116 VTAIL.n237 VSUBS 0.013855f
C1117 VTAIL.n238 VSUBS 0.024561f
C1118 VTAIL.n239 VSUBS 0.024635f
C1119 VTAIL.t13 VSUBS 0.070415f
C1120 VTAIL.n240 VSUBS 0.179878f
C1121 VTAIL.n241 VSUBS 1.04197f
C1122 VTAIL.n242 VSUBS 0.013855f
C1123 VTAIL.n243 VSUBS 0.01467f
C1124 VTAIL.n244 VSUBS 0.032748f
C1125 VTAIL.n245 VSUBS 0.032748f
C1126 VTAIL.n246 VSUBS 0.01467f
C1127 VTAIL.n247 VSUBS 0.013855f
C1128 VTAIL.n248 VSUBS 0.025784f
C1129 VTAIL.n249 VSUBS 0.025784f
C1130 VTAIL.n250 VSUBS 0.013855f
C1131 VTAIL.n251 VSUBS 0.01467f
C1132 VTAIL.n252 VSUBS 0.032748f
C1133 VTAIL.n253 VSUBS 0.032748f
C1134 VTAIL.n254 VSUBS 0.01467f
C1135 VTAIL.n255 VSUBS 0.013855f
C1136 VTAIL.n256 VSUBS 0.025784f
C1137 VTAIL.n257 VSUBS 0.025784f
C1138 VTAIL.n258 VSUBS 0.013855f
C1139 VTAIL.n259 VSUBS 0.01467f
C1140 VTAIL.n260 VSUBS 0.032748f
C1141 VTAIL.n261 VSUBS 0.032748f
C1142 VTAIL.n262 VSUBS 0.032748f
C1143 VTAIL.n263 VSUBS 0.014262f
C1144 VTAIL.n264 VSUBS 0.013855f
C1145 VTAIL.n265 VSUBS 0.025784f
C1146 VTAIL.n266 VSUBS 0.025784f
C1147 VTAIL.n267 VSUBS 0.013855f
C1148 VTAIL.n268 VSUBS 0.01467f
C1149 VTAIL.n269 VSUBS 0.032748f
C1150 VTAIL.n270 VSUBS 0.076306f
C1151 VTAIL.n271 VSUBS 0.01467f
C1152 VTAIL.n272 VSUBS 0.013855f
C1153 VTAIL.n273 VSUBS 0.061359f
C1154 VTAIL.n274 VSUBS 0.038295f
C1155 VTAIL.n275 VSUBS 0.259007f
C1156 VTAIL.n276 VSUBS 0.027458f
C1157 VTAIL.n277 VSUBS 0.025784f
C1158 VTAIL.n278 VSUBS 0.013855f
C1159 VTAIL.n279 VSUBS 0.032748f
C1160 VTAIL.n280 VSUBS 0.01467f
C1161 VTAIL.n281 VSUBS 0.025784f
C1162 VTAIL.n282 VSUBS 0.014262f
C1163 VTAIL.n283 VSUBS 0.032748f
C1164 VTAIL.n284 VSUBS 0.013855f
C1165 VTAIL.n285 VSUBS 0.01467f
C1166 VTAIL.n286 VSUBS 0.025784f
C1167 VTAIL.n287 VSUBS 0.013855f
C1168 VTAIL.n288 VSUBS 0.032748f
C1169 VTAIL.n289 VSUBS 0.01467f
C1170 VTAIL.n290 VSUBS 0.025784f
C1171 VTAIL.n291 VSUBS 0.013855f
C1172 VTAIL.n292 VSUBS 0.024561f
C1173 VTAIL.n293 VSUBS 0.024635f
C1174 VTAIL.t0 VSUBS 0.070415f
C1175 VTAIL.n294 VSUBS 0.179878f
C1176 VTAIL.n295 VSUBS 1.04197f
C1177 VTAIL.n296 VSUBS 0.013855f
C1178 VTAIL.n297 VSUBS 0.01467f
C1179 VTAIL.n298 VSUBS 0.032748f
C1180 VTAIL.n299 VSUBS 0.032748f
C1181 VTAIL.n300 VSUBS 0.01467f
C1182 VTAIL.n301 VSUBS 0.013855f
C1183 VTAIL.n302 VSUBS 0.025784f
C1184 VTAIL.n303 VSUBS 0.025784f
C1185 VTAIL.n304 VSUBS 0.013855f
C1186 VTAIL.n305 VSUBS 0.01467f
C1187 VTAIL.n306 VSUBS 0.032748f
C1188 VTAIL.n307 VSUBS 0.032748f
C1189 VTAIL.n308 VSUBS 0.01467f
C1190 VTAIL.n309 VSUBS 0.013855f
C1191 VTAIL.n310 VSUBS 0.025784f
C1192 VTAIL.n311 VSUBS 0.025784f
C1193 VTAIL.n312 VSUBS 0.013855f
C1194 VTAIL.n313 VSUBS 0.01467f
C1195 VTAIL.n314 VSUBS 0.032748f
C1196 VTAIL.n315 VSUBS 0.032748f
C1197 VTAIL.n316 VSUBS 0.032748f
C1198 VTAIL.n317 VSUBS 0.014262f
C1199 VTAIL.n318 VSUBS 0.013855f
C1200 VTAIL.n319 VSUBS 0.025784f
C1201 VTAIL.n320 VSUBS 0.025784f
C1202 VTAIL.n321 VSUBS 0.013855f
C1203 VTAIL.n322 VSUBS 0.01467f
C1204 VTAIL.n323 VSUBS 0.032748f
C1205 VTAIL.n324 VSUBS 0.076306f
C1206 VTAIL.n325 VSUBS 0.01467f
C1207 VTAIL.n326 VSUBS 0.013855f
C1208 VTAIL.n327 VSUBS 0.061359f
C1209 VTAIL.n328 VSUBS 0.038295f
C1210 VTAIL.n329 VSUBS 0.259007f
C1211 VTAIL.t1 VSUBS 0.203953f
C1212 VTAIL.t6 VSUBS 0.203953f
C1213 VTAIL.n330 VSUBS 1.41852f
C1214 VTAIL.n331 VSUBS 0.946611f
C1215 VTAIL.n332 VSUBS 0.027458f
C1216 VTAIL.n333 VSUBS 0.025784f
C1217 VTAIL.n334 VSUBS 0.013855f
C1218 VTAIL.n335 VSUBS 0.032748f
C1219 VTAIL.n336 VSUBS 0.01467f
C1220 VTAIL.n337 VSUBS 0.025784f
C1221 VTAIL.n338 VSUBS 0.014262f
C1222 VTAIL.n339 VSUBS 0.032748f
C1223 VTAIL.n340 VSUBS 0.013855f
C1224 VTAIL.n341 VSUBS 0.01467f
C1225 VTAIL.n342 VSUBS 0.025784f
C1226 VTAIL.n343 VSUBS 0.013855f
C1227 VTAIL.n344 VSUBS 0.032748f
C1228 VTAIL.n345 VSUBS 0.01467f
C1229 VTAIL.n346 VSUBS 0.025784f
C1230 VTAIL.n347 VSUBS 0.013855f
C1231 VTAIL.n348 VSUBS 0.024561f
C1232 VTAIL.n349 VSUBS 0.024635f
C1233 VTAIL.t5 VSUBS 0.070415f
C1234 VTAIL.n350 VSUBS 0.179878f
C1235 VTAIL.n351 VSUBS 1.04197f
C1236 VTAIL.n352 VSUBS 0.013855f
C1237 VTAIL.n353 VSUBS 0.01467f
C1238 VTAIL.n354 VSUBS 0.032748f
C1239 VTAIL.n355 VSUBS 0.032748f
C1240 VTAIL.n356 VSUBS 0.01467f
C1241 VTAIL.n357 VSUBS 0.013855f
C1242 VTAIL.n358 VSUBS 0.025784f
C1243 VTAIL.n359 VSUBS 0.025784f
C1244 VTAIL.n360 VSUBS 0.013855f
C1245 VTAIL.n361 VSUBS 0.01467f
C1246 VTAIL.n362 VSUBS 0.032748f
C1247 VTAIL.n363 VSUBS 0.032748f
C1248 VTAIL.n364 VSUBS 0.01467f
C1249 VTAIL.n365 VSUBS 0.013855f
C1250 VTAIL.n366 VSUBS 0.025784f
C1251 VTAIL.n367 VSUBS 0.025784f
C1252 VTAIL.n368 VSUBS 0.013855f
C1253 VTAIL.n369 VSUBS 0.01467f
C1254 VTAIL.n370 VSUBS 0.032748f
C1255 VTAIL.n371 VSUBS 0.032748f
C1256 VTAIL.n372 VSUBS 0.032748f
C1257 VTAIL.n373 VSUBS 0.014262f
C1258 VTAIL.n374 VSUBS 0.013855f
C1259 VTAIL.n375 VSUBS 0.025784f
C1260 VTAIL.n376 VSUBS 0.025784f
C1261 VTAIL.n377 VSUBS 0.013855f
C1262 VTAIL.n378 VSUBS 0.01467f
C1263 VTAIL.n379 VSUBS 0.032748f
C1264 VTAIL.n380 VSUBS 0.076306f
C1265 VTAIL.n381 VSUBS 0.01467f
C1266 VTAIL.n382 VSUBS 0.013855f
C1267 VTAIL.n383 VSUBS 0.061359f
C1268 VTAIL.n384 VSUBS 0.038295f
C1269 VTAIL.n385 VSUBS 1.4841f
C1270 VTAIL.n386 VSUBS 0.027458f
C1271 VTAIL.n387 VSUBS 0.025784f
C1272 VTAIL.n388 VSUBS 0.013855f
C1273 VTAIL.n389 VSUBS 0.032748f
C1274 VTAIL.n390 VSUBS 0.01467f
C1275 VTAIL.n391 VSUBS 0.025784f
C1276 VTAIL.n392 VSUBS 0.014262f
C1277 VTAIL.n393 VSUBS 0.032748f
C1278 VTAIL.n394 VSUBS 0.01467f
C1279 VTAIL.n395 VSUBS 0.025784f
C1280 VTAIL.n396 VSUBS 0.013855f
C1281 VTAIL.n397 VSUBS 0.032748f
C1282 VTAIL.n398 VSUBS 0.01467f
C1283 VTAIL.n399 VSUBS 0.025784f
C1284 VTAIL.n400 VSUBS 0.013855f
C1285 VTAIL.n401 VSUBS 0.024561f
C1286 VTAIL.n402 VSUBS 0.024635f
C1287 VTAIL.t14 VSUBS 0.070415f
C1288 VTAIL.n403 VSUBS 0.179878f
C1289 VTAIL.n404 VSUBS 1.04197f
C1290 VTAIL.n405 VSUBS 0.013855f
C1291 VTAIL.n406 VSUBS 0.01467f
C1292 VTAIL.n407 VSUBS 0.032748f
C1293 VTAIL.n408 VSUBS 0.032748f
C1294 VTAIL.n409 VSUBS 0.01467f
C1295 VTAIL.n410 VSUBS 0.013855f
C1296 VTAIL.n411 VSUBS 0.025784f
C1297 VTAIL.n412 VSUBS 0.025784f
C1298 VTAIL.n413 VSUBS 0.013855f
C1299 VTAIL.n414 VSUBS 0.01467f
C1300 VTAIL.n415 VSUBS 0.032748f
C1301 VTAIL.n416 VSUBS 0.032748f
C1302 VTAIL.n417 VSUBS 0.01467f
C1303 VTAIL.n418 VSUBS 0.013855f
C1304 VTAIL.n419 VSUBS 0.025784f
C1305 VTAIL.n420 VSUBS 0.025784f
C1306 VTAIL.n421 VSUBS 0.013855f
C1307 VTAIL.n422 VSUBS 0.013855f
C1308 VTAIL.n423 VSUBS 0.01467f
C1309 VTAIL.n424 VSUBS 0.032748f
C1310 VTAIL.n425 VSUBS 0.032748f
C1311 VTAIL.n426 VSUBS 0.032748f
C1312 VTAIL.n427 VSUBS 0.014262f
C1313 VTAIL.n428 VSUBS 0.013855f
C1314 VTAIL.n429 VSUBS 0.025784f
C1315 VTAIL.n430 VSUBS 0.025784f
C1316 VTAIL.n431 VSUBS 0.013855f
C1317 VTAIL.n432 VSUBS 0.01467f
C1318 VTAIL.n433 VSUBS 0.032748f
C1319 VTAIL.n434 VSUBS 0.076306f
C1320 VTAIL.n435 VSUBS 0.01467f
C1321 VTAIL.n436 VSUBS 0.013855f
C1322 VTAIL.n437 VSUBS 0.061359f
C1323 VTAIL.n438 VSUBS 0.038295f
C1324 VTAIL.n439 VSUBS 1.47926f
C1325 VN.n0 VSUBS 0.041853f
C1326 VN.t7 VSUBS 2.08333f
C1327 VN.n1 VSUBS 0.046342f
C1328 VN.n2 VSUBS 0.031745f
C1329 VN.t5 VSUBS 2.08333f
C1330 VN.n3 VSUBS 0.747574f
C1331 VN.n4 VSUBS 0.031745f
C1332 VN.n5 VSUBS 0.063093f
C1333 VN.t6 VSUBS 2.31219f
C1334 VN.n6 VSUBS 0.818137f
C1335 VN.t0 VSUBS 2.08333f
C1336 VN.n7 VSUBS 0.843112f
C1337 VN.n8 VSUBS 0.051861f
C1338 VN.n9 VSUBS 0.300557f
C1339 VN.n10 VSUBS 0.031745f
C1340 VN.n11 VSUBS 0.031745f
C1341 VN.n12 VSUBS 0.025663f
C1342 VN.n13 VSUBS 0.063093f
C1343 VN.n14 VSUBS 0.051861f
C1344 VN.n15 VSUBS 0.031745f
C1345 VN.n16 VSUBS 0.031745f
C1346 VN.n17 VSUBS 0.037256f
C1347 VN.n18 VSUBS 0.059165f
C1348 VN.n19 VSUBS 0.046342f
C1349 VN.n20 VSUBS 0.031745f
C1350 VN.n21 VSUBS 0.031745f
C1351 VN.n22 VSUBS 0.031745f
C1352 VN.n23 VSUBS 0.059165f
C1353 VN.n24 VSUBS 0.037256f
C1354 VN.n25 VSUBS 0.839814f
C1355 VN.n26 VSUBS 0.052521f
C1356 VN.n27 VSUBS 0.041853f
C1357 VN.t3 VSUBS 2.08333f
C1358 VN.n28 VSUBS 0.046342f
C1359 VN.n29 VSUBS 0.031745f
C1360 VN.t1 VSUBS 2.08333f
C1361 VN.n30 VSUBS 0.747574f
C1362 VN.n31 VSUBS 0.031745f
C1363 VN.n32 VSUBS 0.063093f
C1364 VN.t2 VSUBS 2.31219f
C1365 VN.n33 VSUBS 0.818137f
C1366 VN.t4 VSUBS 2.08333f
C1367 VN.n34 VSUBS 0.843112f
C1368 VN.n35 VSUBS 0.051861f
C1369 VN.n36 VSUBS 0.300557f
C1370 VN.n37 VSUBS 0.031745f
C1371 VN.n38 VSUBS 0.031745f
C1372 VN.n39 VSUBS 0.025663f
C1373 VN.n40 VSUBS 0.063093f
C1374 VN.n41 VSUBS 0.051861f
C1375 VN.n42 VSUBS 0.031745f
C1376 VN.n43 VSUBS 0.031745f
C1377 VN.n44 VSUBS 0.037256f
C1378 VN.n45 VSUBS 0.059165f
C1379 VN.n46 VSUBS 0.046342f
C1380 VN.n47 VSUBS 0.031745f
C1381 VN.n48 VSUBS 0.031745f
C1382 VN.n49 VSUBS 0.031745f
C1383 VN.n50 VSUBS 0.059165f
C1384 VN.n51 VSUBS 0.037256f
C1385 VN.n52 VSUBS 0.839814f
C1386 VN.n53 VSUBS 1.70301f
.ends

