* NGSPICE file created from diff_pair_sample_0937.ext - technology: sky130A

.subckt diff_pair_sample_0937 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t7 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X1 B.t11 B.t9 B.t10 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=2.8
X2 VTAIL.t10 VN.t1 VDD2.t6 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X3 VDD2.t5 VN.t2 VTAIL.t9 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=2.8
X4 VDD2.t4 VN.t3 VTAIL.t12 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X5 VDD1.t7 VP.t0 VTAIL.t3 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X6 VTAIL.t13 VN.t4 VDD2.t3 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X7 B.t8 B.t6 B.t7 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=2.8
X8 VDD1.t6 VP.t1 VTAIL.t15 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X9 VDD1.t5 VP.t2 VTAIL.t5 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=2.8
X10 VTAIL.t2 VP.t3 VDD1.t4 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=2.8
X11 VDD2.t2 VN.t5 VTAIL.t11 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=2.8
X12 B.t5 B.t3 B.t4 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=2.8
X13 VTAIL.t1 VP.t4 VDD1.t3 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X14 VDD1.t2 VP.t5 VTAIL.t0 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=2.8
X15 VTAIL.t6 VP.t6 VDD1.t1 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=2.8
X16 B.t2 B.t0 B.t1 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=2.8
X17 VTAIL.t8 VN.t6 VDD2.t1 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=2.8
X18 VTAIL.t4 VP.t7 VDD1.t0 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=2.8
X19 VTAIL.t14 VN.t7 VDD2.t0 w_n4100_n1574# sky130_fd_pr__pfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=2.8
R0 VN.n56 VN.n55 161.3
R1 VN.n54 VN.n30 161.3
R2 VN.n53 VN.n52 161.3
R3 VN.n51 VN.n31 161.3
R4 VN.n50 VN.n49 161.3
R5 VN.n48 VN.n32 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n27 VN.n26 161.3
R13 VN.n25 VN.n1 161.3
R14 VN.n24 VN.n23 161.3
R15 VN.n22 VN.n2 161.3
R16 VN.n21 VN.n20 161.3
R17 VN.n19 VN.n3 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n28 VN.n0 68.2918
R25 VN.n57 VN.n29 68.2918
R26 VN.n8 VN.n7 58.2301
R27 VN.n37 VN.n36 58.2301
R28 VN.n37 VN.t5 57.9638
R29 VN.n8 VN.t7 57.9638
R30 VN.n13 VN.n12 56.5193
R31 VN.n42 VN.n41 56.5193
R32 VN.n24 VN.n2 52.1486
R33 VN.n53 VN.n31 52.1486
R34 VN VN.n57 45.3011
R35 VN.n25 VN.n24 28.8382
R36 VN.n54 VN.n53 28.8382
R37 VN.n7 VN.t3 26.0801
R38 VN.n18 VN.t1 26.0801
R39 VN.n0 VN.t2 26.0801
R40 VN.n36 VN.t4 26.0801
R41 VN.n47 VN.t0 26.0801
R42 VN.n29 VN.t6 26.0801
R43 VN.n11 VN.n6 24.4675
R44 VN.n12 VN.n11 24.4675
R45 VN.n13 VN.n4 24.4675
R46 VN.n17 VN.n4 24.4675
R47 VN.n20 VN.n19 24.4675
R48 VN.n20 VN.n2 24.4675
R49 VN.n26 VN.n25 24.4675
R50 VN.n41 VN.n40 24.4675
R51 VN.n40 VN.n35 24.4675
R52 VN.n49 VN.n31 24.4675
R53 VN.n49 VN.n48 24.4675
R54 VN.n46 VN.n33 24.4675
R55 VN.n42 VN.n33 24.4675
R56 VN.n55 VN.n54 24.4675
R57 VN.n26 VN.n0 21.7761
R58 VN.n55 VN.n29 21.7761
R59 VN.n7 VN.n6 15.4147
R60 VN.n18 VN.n17 15.4147
R61 VN.n36 VN.n35 15.4147
R62 VN.n47 VN.n46 15.4147
R63 VN.n19 VN.n18 9.05329
R64 VN.n48 VN.n47 9.05329
R65 VN.n38 VN.n37 5.40755
R66 VN.n9 VN.n8 5.40755
R67 VN.n57 VN.n56 0.354971
R68 VN.n28 VN.n27 0.354971
R69 VN VN.n28 0.26696
R70 VN.n56 VN.n30 0.189894
R71 VN.n52 VN.n30 0.189894
R72 VN.n52 VN.n51 0.189894
R73 VN.n51 VN.n50 0.189894
R74 VN.n50 VN.n32 0.189894
R75 VN.n45 VN.n32 0.189894
R76 VN.n45 VN.n44 0.189894
R77 VN.n44 VN.n43 0.189894
R78 VN.n43 VN.n34 0.189894
R79 VN.n39 VN.n34 0.189894
R80 VN.n39 VN.n38 0.189894
R81 VN.n10 VN.n9 0.189894
R82 VN.n10 VN.n5 0.189894
R83 VN.n14 VN.n5 0.189894
R84 VN.n15 VN.n14 0.189894
R85 VN.n16 VN.n15 0.189894
R86 VN.n16 VN.n3 0.189894
R87 VN.n21 VN.n3 0.189894
R88 VN.n22 VN.n21 0.189894
R89 VN.n23 VN.n22 0.189894
R90 VN.n23 VN.n1 0.189894
R91 VN.n27 VN.n1 0.189894
R92 VTAIL.n14 VTAIL.t0 131.593
R93 VTAIL.n11 VTAIL.t6 131.593
R94 VTAIL.n10 VTAIL.t11 131.593
R95 VTAIL.n7 VTAIL.t8 131.593
R96 VTAIL.n15 VTAIL.t9 131.593
R97 VTAIL.n2 VTAIL.t14 131.593
R98 VTAIL.n3 VTAIL.t5 131.593
R99 VTAIL.n6 VTAIL.t2 131.593
R100 VTAIL.n13 VTAIL.n12 120.865
R101 VTAIL.n9 VTAIL.n8 120.865
R102 VTAIL.n1 VTAIL.n0 120.865
R103 VTAIL.n5 VTAIL.n4 120.865
R104 VTAIL.n15 VTAIL.n14 17.6772
R105 VTAIL.n7 VTAIL.n6 17.6772
R106 VTAIL.n0 VTAIL.t12 10.7282
R107 VTAIL.n0 VTAIL.t10 10.7282
R108 VTAIL.n4 VTAIL.t3 10.7282
R109 VTAIL.n4 VTAIL.t1 10.7282
R110 VTAIL.n12 VTAIL.t15 10.7282
R111 VTAIL.n12 VTAIL.t4 10.7282
R112 VTAIL.n8 VTAIL.t7 10.7282
R113 VTAIL.n8 VTAIL.t13 10.7282
R114 VTAIL.n9 VTAIL.n7 2.69878
R115 VTAIL.n10 VTAIL.n9 2.69878
R116 VTAIL.n13 VTAIL.n11 2.69878
R117 VTAIL.n14 VTAIL.n13 2.69878
R118 VTAIL.n6 VTAIL.n5 2.69878
R119 VTAIL.n5 VTAIL.n3 2.69878
R120 VTAIL.n2 VTAIL.n1 2.69878
R121 VTAIL VTAIL.n15 2.64059
R122 VTAIL.n11 VTAIL.n10 0.470328
R123 VTAIL.n3 VTAIL.n2 0.470328
R124 VTAIL VTAIL.n1 0.0586897
R125 VDD2.n2 VDD2.n1 138.838
R126 VDD2.n2 VDD2.n0 138.838
R127 VDD2 VDD2.n5 138.834
R128 VDD2.n4 VDD2.n3 137.543
R129 VDD2.n4 VDD2.n2 38.4696
R130 VDD2.n5 VDD2.t3 10.7282
R131 VDD2.n5 VDD2.t2 10.7282
R132 VDD2.n3 VDD2.t1 10.7282
R133 VDD2.n3 VDD2.t7 10.7282
R134 VDD2.n1 VDD2.t6 10.7282
R135 VDD2.n1 VDD2.t5 10.7282
R136 VDD2.n0 VDD2.t0 10.7282
R137 VDD2.n0 VDD2.t4 10.7282
R138 VDD2 VDD2.n4 1.40783
R139 B.n465 B.n464 585
R140 B.n466 B.n53 585
R141 B.n468 B.n467 585
R142 B.n469 B.n52 585
R143 B.n471 B.n470 585
R144 B.n472 B.n51 585
R145 B.n474 B.n473 585
R146 B.n475 B.n50 585
R147 B.n477 B.n476 585
R148 B.n478 B.n49 585
R149 B.n480 B.n479 585
R150 B.n481 B.n48 585
R151 B.n483 B.n482 585
R152 B.n484 B.n47 585
R153 B.n486 B.n485 585
R154 B.n488 B.n44 585
R155 B.n490 B.n489 585
R156 B.n491 B.n43 585
R157 B.n493 B.n492 585
R158 B.n494 B.n42 585
R159 B.n496 B.n495 585
R160 B.n497 B.n41 585
R161 B.n499 B.n498 585
R162 B.n500 B.n37 585
R163 B.n502 B.n501 585
R164 B.n503 B.n36 585
R165 B.n505 B.n504 585
R166 B.n506 B.n35 585
R167 B.n508 B.n507 585
R168 B.n509 B.n34 585
R169 B.n511 B.n510 585
R170 B.n512 B.n33 585
R171 B.n514 B.n513 585
R172 B.n515 B.n32 585
R173 B.n517 B.n516 585
R174 B.n518 B.n31 585
R175 B.n520 B.n519 585
R176 B.n521 B.n30 585
R177 B.n523 B.n522 585
R178 B.n524 B.n29 585
R179 B.n463 B.n54 585
R180 B.n462 B.n461 585
R181 B.n460 B.n55 585
R182 B.n459 B.n458 585
R183 B.n457 B.n56 585
R184 B.n456 B.n455 585
R185 B.n454 B.n57 585
R186 B.n453 B.n452 585
R187 B.n451 B.n58 585
R188 B.n450 B.n449 585
R189 B.n448 B.n59 585
R190 B.n447 B.n446 585
R191 B.n445 B.n60 585
R192 B.n444 B.n443 585
R193 B.n442 B.n61 585
R194 B.n441 B.n440 585
R195 B.n439 B.n62 585
R196 B.n438 B.n437 585
R197 B.n436 B.n63 585
R198 B.n435 B.n434 585
R199 B.n433 B.n64 585
R200 B.n432 B.n431 585
R201 B.n430 B.n65 585
R202 B.n429 B.n428 585
R203 B.n427 B.n66 585
R204 B.n426 B.n425 585
R205 B.n424 B.n67 585
R206 B.n423 B.n422 585
R207 B.n421 B.n68 585
R208 B.n420 B.n419 585
R209 B.n418 B.n69 585
R210 B.n417 B.n416 585
R211 B.n415 B.n70 585
R212 B.n414 B.n413 585
R213 B.n412 B.n71 585
R214 B.n411 B.n410 585
R215 B.n409 B.n72 585
R216 B.n408 B.n407 585
R217 B.n406 B.n73 585
R218 B.n405 B.n404 585
R219 B.n403 B.n74 585
R220 B.n402 B.n401 585
R221 B.n400 B.n75 585
R222 B.n399 B.n398 585
R223 B.n397 B.n76 585
R224 B.n396 B.n395 585
R225 B.n394 B.n77 585
R226 B.n393 B.n392 585
R227 B.n391 B.n78 585
R228 B.n390 B.n389 585
R229 B.n388 B.n79 585
R230 B.n387 B.n386 585
R231 B.n385 B.n80 585
R232 B.n384 B.n383 585
R233 B.n382 B.n81 585
R234 B.n381 B.n380 585
R235 B.n379 B.n82 585
R236 B.n378 B.n377 585
R237 B.n376 B.n83 585
R238 B.n375 B.n374 585
R239 B.n373 B.n84 585
R240 B.n372 B.n371 585
R241 B.n370 B.n85 585
R242 B.n369 B.n368 585
R243 B.n367 B.n86 585
R244 B.n366 B.n365 585
R245 B.n364 B.n87 585
R246 B.n363 B.n362 585
R247 B.n361 B.n88 585
R248 B.n360 B.n359 585
R249 B.n358 B.n89 585
R250 B.n357 B.n356 585
R251 B.n355 B.n90 585
R252 B.n354 B.n353 585
R253 B.n352 B.n91 585
R254 B.n351 B.n350 585
R255 B.n349 B.n92 585
R256 B.n348 B.n347 585
R257 B.n346 B.n93 585
R258 B.n345 B.n344 585
R259 B.n343 B.n94 585
R260 B.n342 B.n341 585
R261 B.n340 B.n95 585
R262 B.n339 B.n338 585
R263 B.n337 B.n96 585
R264 B.n336 B.n335 585
R265 B.n334 B.n97 585
R266 B.n333 B.n332 585
R267 B.n331 B.n98 585
R268 B.n330 B.n329 585
R269 B.n328 B.n99 585
R270 B.n327 B.n326 585
R271 B.n325 B.n100 585
R272 B.n324 B.n323 585
R273 B.n322 B.n101 585
R274 B.n321 B.n320 585
R275 B.n319 B.n102 585
R276 B.n318 B.n317 585
R277 B.n316 B.n103 585
R278 B.n315 B.n314 585
R279 B.n313 B.n104 585
R280 B.n312 B.n311 585
R281 B.n310 B.n105 585
R282 B.n309 B.n308 585
R283 B.n307 B.n106 585
R284 B.n306 B.n305 585
R285 B.n304 B.n107 585
R286 B.n303 B.n302 585
R287 B.n301 B.n108 585
R288 B.n240 B.n239 585
R289 B.n241 B.n132 585
R290 B.n243 B.n242 585
R291 B.n244 B.n131 585
R292 B.n246 B.n245 585
R293 B.n247 B.n130 585
R294 B.n249 B.n248 585
R295 B.n250 B.n129 585
R296 B.n252 B.n251 585
R297 B.n253 B.n128 585
R298 B.n255 B.n254 585
R299 B.n256 B.n127 585
R300 B.n258 B.n257 585
R301 B.n259 B.n126 585
R302 B.n261 B.n260 585
R303 B.n263 B.n262 585
R304 B.n264 B.n122 585
R305 B.n266 B.n265 585
R306 B.n267 B.n121 585
R307 B.n269 B.n268 585
R308 B.n270 B.n120 585
R309 B.n272 B.n271 585
R310 B.n273 B.n119 585
R311 B.n275 B.n274 585
R312 B.n276 B.n116 585
R313 B.n279 B.n278 585
R314 B.n280 B.n115 585
R315 B.n282 B.n281 585
R316 B.n283 B.n114 585
R317 B.n285 B.n284 585
R318 B.n286 B.n113 585
R319 B.n288 B.n287 585
R320 B.n289 B.n112 585
R321 B.n291 B.n290 585
R322 B.n292 B.n111 585
R323 B.n294 B.n293 585
R324 B.n295 B.n110 585
R325 B.n297 B.n296 585
R326 B.n298 B.n109 585
R327 B.n300 B.n299 585
R328 B.n238 B.n133 585
R329 B.n237 B.n236 585
R330 B.n235 B.n134 585
R331 B.n234 B.n233 585
R332 B.n232 B.n135 585
R333 B.n231 B.n230 585
R334 B.n229 B.n136 585
R335 B.n228 B.n227 585
R336 B.n226 B.n137 585
R337 B.n225 B.n224 585
R338 B.n223 B.n138 585
R339 B.n222 B.n221 585
R340 B.n220 B.n139 585
R341 B.n219 B.n218 585
R342 B.n217 B.n140 585
R343 B.n216 B.n215 585
R344 B.n214 B.n141 585
R345 B.n213 B.n212 585
R346 B.n211 B.n142 585
R347 B.n210 B.n209 585
R348 B.n208 B.n143 585
R349 B.n207 B.n206 585
R350 B.n205 B.n144 585
R351 B.n204 B.n203 585
R352 B.n202 B.n145 585
R353 B.n201 B.n200 585
R354 B.n199 B.n146 585
R355 B.n198 B.n197 585
R356 B.n196 B.n147 585
R357 B.n195 B.n194 585
R358 B.n193 B.n148 585
R359 B.n192 B.n191 585
R360 B.n190 B.n149 585
R361 B.n189 B.n188 585
R362 B.n187 B.n150 585
R363 B.n186 B.n185 585
R364 B.n184 B.n151 585
R365 B.n183 B.n182 585
R366 B.n181 B.n152 585
R367 B.n180 B.n179 585
R368 B.n178 B.n153 585
R369 B.n177 B.n176 585
R370 B.n175 B.n154 585
R371 B.n174 B.n173 585
R372 B.n172 B.n155 585
R373 B.n171 B.n170 585
R374 B.n169 B.n156 585
R375 B.n168 B.n167 585
R376 B.n166 B.n157 585
R377 B.n165 B.n164 585
R378 B.n163 B.n158 585
R379 B.n162 B.n161 585
R380 B.n160 B.n159 585
R381 B.n2 B.n0 585
R382 B.n605 B.n1 585
R383 B.n604 B.n603 585
R384 B.n602 B.n3 585
R385 B.n601 B.n600 585
R386 B.n599 B.n4 585
R387 B.n598 B.n597 585
R388 B.n596 B.n5 585
R389 B.n595 B.n594 585
R390 B.n593 B.n6 585
R391 B.n592 B.n591 585
R392 B.n590 B.n7 585
R393 B.n589 B.n588 585
R394 B.n587 B.n8 585
R395 B.n586 B.n585 585
R396 B.n584 B.n9 585
R397 B.n583 B.n582 585
R398 B.n581 B.n10 585
R399 B.n580 B.n579 585
R400 B.n578 B.n11 585
R401 B.n577 B.n576 585
R402 B.n575 B.n12 585
R403 B.n574 B.n573 585
R404 B.n572 B.n13 585
R405 B.n571 B.n570 585
R406 B.n569 B.n14 585
R407 B.n568 B.n567 585
R408 B.n566 B.n15 585
R409 B.n565 B.n564 585
R410 B.n563 B.n16 585
R411 B.n562 B.n561 585
R412 B.n560 B.n17 585
R413 B.n559 B.n558 585
R414 B.n557 B.n18 585
R415 B.n556 B.n555 585
R416 B.n554 B.n19 585
R417 B.n553 B.n552 585
R418 B.n551 B.n20 585
R419 B.n550 B.n549 585
R420 B.n548 B.n21 585
R421 B.n547 B.n546 585
R422 B.n545 B.n22 585
R423 B.n544 B.n543 585
R424 B.n542 B.n23 585
R425 B.n541 B.n540 585
R426 B.n539 B.n24 585
R427 B.n538 B.n537 585
R428 B.n536 B.n25 585
R429 B.n535 B.n534 585
R430 B.n533 B.n26 585
R431 B.n532 B.n531 585
R432 B.n530 B.n27 585
R433 B.n529 B.n528 585
R434 B.n527 B.n28 585
R435 B.n526 B.n525 585
R436 B.n607 B.n606 585
R437 B.n239 B.n238 526.135
R438 B.n526 B.n29 526.135
R439 B.n299 B.n108 526.135
R440 B.n465 B.n54 526.135
R441 B.n117 B.t3 234.41
R442 B.n123 B.t9 234.41
R443 B.n38 B.t0 234.41
R444 B.n45 B.t6 234.41
R445 B.n117 B.t5 206.4
R446 B.n45 B.t7 206.4
R447 B.n123 B.t11 206.399
R448 B.n38 B.t1 206.399
R449 B.n238 B.n237 163.367
R450 B.n237 B.n134 163.367
R451 B.n233 B.n134 163.367
R452 B.n233 B.n232 163.367
R453 B.n232 B.n231 163.367
R454 B.n231 B.n136 163.367
R455 B.n227 B.n136 163.367
R456 B.n227 B.n226 163.367
R457 B.n226 B.n225 163.367
R458 B.n225 B.n138 163.367
R459 B.n221 B.n138 163.367
R460 B.n221 B.n220 163.367
R461 B.n220 B.n219 163.367
R462 B.n219 B.n140 163.367
R463 B.n215 B.n140 163.367
R464 B.n215 B.n214 163.367
R465 B.n214 B.n213 163.367
R466 B.n213 B.n142 163.367
R467 B.n209 B.n142 163.367
R468 B.n209 B.n208 163.367
R469 B.n208 B.n207 163.367
R470 B.n207 B.n144 163.367
R471 B.n203 B.n144 163.367
R472 B.n203 B.n202 163.367
R473 B.n202 B.n201 163.367
R474 B.n201 B.n146 163.367
R475 B.n197 B.n146 163.367
R476 B.n197 B.n196 163.367
R477 B.n196 B.n195 163.367
R478 B.n195 B.n148 163.367
R479 B.n191 B.n148 163.367
R480 B.n191 B.n190 163.367
R481 B.n190 B.n189 163.367
R482 B.n189 B.n150 163.367
R483 B.n185 B.n150 163.367
R484 B.n185 B.n184 163.367
R485 B.n184 B.n183 163.367
R486 B.n183 B.n152 163.367
R487 B.n179 B.n152 163.367
R488 B.n179 B.n178 163.367
R489 B.n178 B.n177 163.367
R490 B.n177 B.n154 163.367
R491 B.n173 B.n154 163.367
R492 B.n173 B.n172 163.367
R493 B.n172 B.n171 163.367
R494 B.n171 B.n156 163.367
R495 B.n167 B.n156 163.367
R496 B.n167 B.n166 163.367
R497 B.n166 B.n165 163.367
R498 B.n165 B.n158 163.367
R499 B.n161 B.n158 163.367
R500 B.n161 B.n160 163.367
R501 B.n160 B.n2 163.367
R502 B.n606 B.n2 163.367
R503 B.n606 B.n605 163.367
R504 B.n605 B.n604 163.367
R505 B.n604 B.n3 163.367
R506 B.n600 B.n3 163.367
R507 B.n600 B.n599 163.367
R508 B.n599 B.n598 163.367
R509 B.n598 B.n5 163.367
R510 B.n594 B.n5 163.367
R511 B.n594 B.n593 163.367
R512 B.n593 B.n592 163.367
R513 B.n592 B.n7 163.367
R514 B.n588 B.n7 163.367
R515 B.n588 B.n587 163.367
R516 B.n587 B.n586 163.367
R517 B.n586 B.n9 163.367
R518 B.n582 B.n9 163.367
R519 B.n582 B.n581 163.367
R520 B.n581 B.n580 163.367
R521 B.n580 B.n11 163.367
R522 B.n576 B.n11 163.367
R523 B.n576 B.n575 163.367
R524 B.n575 B.n574 163.367
R525 B.n574 B.n13 163.367
R526 B.n570 B.n13 163.367
R527 B.n570 B.n569 163.367
R528 B.n569 B.n568 163.367
R529 B.n568 B.n15 163.367
R530 B.n564 B.n15 163.367
R531 B.n564 B.n563 163.367
R532 B.n563 B.n562 163.367
R533 B.n562 B.n17 163.367
R534 B.n558 B.n17 163.367
R535 B.n558 B.n557 163.367
R536 B.n557 B.n556 163.367
R537 B.n556 B.n19 163.367
R538 B.n552 B.n19 163.367
R539 B.n552 B.n551 163.367
R540 B.n551 B.n550 163.367
R541 B.n550 B.n21 163.367
R542 B.n546 B.n21 163.367
R543 B.n546 B.n545 163.367
R544 B.n545 B.n544 163.367
R545 B.n544 B.n23 163.367
R546 B.n540 B.n23 163.367
R547 B.n540 B.n539 163.367
R548 B.n539 B.n538 163.367
R549 B.n538 B.n25 163.367
R550 B.n534 B.n25 163.367
R551 B.n534 B.n533 163.367
R552 B.n533 B.n532 163.367
R553 B.n532 B.n27 163.367
R554 B.n528 B.n27 163.367
R555 B.n528 B.n527 163.367
R556 B.n527 B.n526 163.367
R557 B.n239 B.n132 163.367
R558 B.n243 B.n132 163.367
R559 B.n244 B.n243 163.367
R560 B.n245 B.n244 163.367
R561 B.n245 B.n130 163.367
R562 B.n249 B.n130 163.367
R563 B.n250 B.n249 163.367
R564 B.n251 B.n250 163.367
R565 B.n251 B.n128 163.367
R566 B.n255 B.n128 163.367
R567 B.n256 B.n255 163.367
R568 B.n257 B.n256 163.367
R569 B.n257 B.n126 163.367
R570 B.n261 B.n126 163.367
R571 B.n262 B.n261 163.367
R572 B.n262 B.n122 163.367
R573 B.n266 B.n122 163.367
R574 B.n267 B.n266 163.367
R575 B.n268 B.n267 163.367
R576 B.n268 B.n120 163.367
R577 B.n272 B.n120 163.367
R578 B.n273 B.n272 163.367
R579 B.n274 B.n273 163.367
R580 B.n274 B.n116 163.367
R581 B.n279 B.n116 163.367
R582 B.n280 B.n279 163.367
R583 B.n281 B.n280 163.367
R584 B.n281 B.n114 163.367
R585 B.n285 B.n114 163.367
R586 B.n286 B.n285 163.367
R587 B.n287 B.n286 163.367
R588 B.n287 B.n112 163.367
R589 B.n291 B.n112 163.367
R590 B.n292 B.n291 163.367
R591 B.n293 B.n292 163.367
R592 B.n293 B.n110 163.367
R593 B.n297 B.n110 163.367
R594 B.n298 B.n297 163.367
R595 B.n299 B.n298 163.367
R596 B.n303 B.n108 163.367
R597 B.n304 B.n303 163.367
R598 B.n305 B.n304 163.367
R599 B.n305 B.n106 163.367
R600 B.n309 B.n106 163.367
R601 B.n310 B.n309 163.367
R602 B.n311 B.n310 163.367
R603 B.n311 B.n104 163.367
R604 B.n315 B.n104 163.367
R605 B.n316 B.n315 163.367
R606 B.n317 B.n316 163.367
R607 B.n317 B.n102 163.367
R608 B.n321 B.n102 163.367
R609 B.n322 B.n321 163.367
R610 B.n323 B.n322 163.367
R611 B.n323 B.n100 163.367
R612 B.n327 B.n100 163.367
R613 B.n328 B.n327 163.367
R614 B.n329 B.n328 163.367
R615 B.n329 B.n98 163.367
R616 B.n333 B.n98 163.367
R617 B.n334 B.n333 163.367
R618 B.n335 B.n334 163.367
R619 B.n335 B.n96 163.367
R620 B.n339 B.n96 163.367
R621 B.n340 B.n339 163.367
R622 B.n341 B.n340 163.367
R623 B.n341 B.n94 163.367
R624 B.n345 B.n94 163.367
R625 B.n346 B.n345 163.367
R626 B.n347 B.n346 163.367
R627 B.n347 B.n92 163.367
R628 B.n351 B.n92 163.367
R629 B.n352 B.n351 163.367
R630 B.n353 B.n352 163.367
R631 B.n353 B.n90 163.367
R632 B.n357 B.n90 163.367
R633 B.n358 B.n357 163.367
R634 B.n359 B.n358 163.367
R635 B.n359 B.n88 163.367
R636 B.n363 B.n88 163.367
R637 B.n364 B.n363 163.367
R638 B.n365 B.n364 163.367
R639 B.n365 B.n86 163.367
R640 B.n369 B.n86 163.367
R641 B.n370 B.n369 163.367
R642 B.n371 B.n370 163.367
R643 B.n371 B.n84 163.367
R644 B.n375 B.n84 163.367
R645 B.n376 B.n375 163.367
R646 B.n377 B.n376 163.367
R647 B.n377 B.n82 163.367
R648 B.n381 B.n82 163.367
R649 B.n382 B.n381 163.367
R650 B.n383 B.n382 163.367
R651 B.n383 B.n80 163.367
R652 B.n387 B.n80 163.367
R653 B.n388 B.n387 163.367
R654 B.n389 B.n388 163.367
R655 B.n389 B.n78 163.367
R656 B.n393 B.n78 163.367
R657 B.n394 B.n393 163.367
R658 B.n395 B.n394 163.367
R659 B.n395 B.n76 163.367
R660 B.n399 B.n76 163.367
R661 B.n400 B.n399 163.367
R662 B.n401 B.n400 163.367
R663 B.n401 B.n74 163.367
R664 B.n405 B.n74 163.367
R665 B.n406 B.n405 163.367
R666 B.n407 B.n406 163.367
R667 B.n407 B.n72 163.367
R668 B.n411 B.n72 163.367
R669 B.n412 B.n411 163.367
R670 B.n413 B.n412 163.367
R671 B.n413 B.n70 163.367
R672 B.n417 B.n70 163.367
R673 B.n418 B.n417 163.367
R674 B.n419 B.n418 163.367
R675 B.n419 B.n68 163.367
R676 B.n423 B.n68 163.367
R677 B.n424 B.n423 163.367
R678 B.n425 B.n424 163.367
R679 B.n425 B.n66 163.367
R680 B.n429 B.n66 163.367
R681 B.n430 B.n429 163.367
R682 B.n431 B.n430 163.367
R683 B.n431 B.n64 163.367
R684 B.n435 B.n64 163.367
R685 B.n436 B.n435 163.367
R686 B.n437 B.n436 163.367
R687 B.n437 B.n62 163.367
R688 B.n441 B.n62 163.367
R689 B.n442 B.n441 163.367
R690 B.n443 B.n442 163.367
R691 B.n443 B.n60 163.367
R692 B.n447 B.n60 163.367
R693 B.n448 B.n447 163.367
R694 B.n449 B.n448 163.367
R695 B.n449 B.n58 163.367
R696 B.n453 B.n58 163.367
R697 B.n454 B.n453 163.367
R698 B.n455 B.n454 163.367
R699 B.n455 B.n56 163.367
R700 B.n459 B.n56 163.367
R701 B.n460 B.n459 163.367
R702 B.n461 B.n460 163.367
R703 B.n461 B.n54 163.367
R704 B.n522 B.n29 163.367
R705 B.n522 B.n521 163.367
R706 B.n521 B.n520 163.367
R707 B.n520 B.n31 163.367
R708 B.n516 B.n31 163.367
R709 B.n516 B.n515 163.367
R710 B.n515 B.n514 163.367
R711 B.n514 B.n33 163.367
R712 B.n510 B.n33 163.367
R713 B.n510 B.n509 163.367
R714 B.n509 B.n508 163.367
R715 B.n508 B.n35 163.367
R716 B.n504 B.n35 163.367
R717 B.n504 B.n503 163.367
R718 B.n503 B.n502 163.367
R719 B.n502 B.n37 163.367
R720 B.n498 B.n37 163.367
R721 B.n498 B.n497 163.367
R722 B.n497 B.n496 163.367
R723 B.n496 B.n42 163.367
R724 B.n492 B.n42 163.367
R725 B.n492 B.n491 163.367
R726 B.n491 B.n490 163.367
R727 B.n490 B.n44 163.367
R728 B.n485 B.n44 163.367
R729 B.n485 B.n484 163.367
R730 B.n484 B.n483 163.367
R731 B.n483 B.n48 163.367
R732 B.n479 B.n48 163.367
R733 B.n479 B.n478 163.367
R734 B.n478 B.n477 163.367
R735 B.n477 B.n50 163.367
R736 B.n473 B.n50 163.367
R737 B.n473 B.n472 163.367
R738 B.n472 B.n471 163.367
R739 B.n471 B.n52 163.367
R740 B.n467 B.n52 163.367
R741 B.n467 B.n466 163.367
R742 B.n466 B.n465 163.367
R743 B.n118 B.t4 145.697
R744 B.n46 B.t8 145.697
R745 B.n124 B.t10 145.696
R746 B.n39 B.t2 145.696
R747 B.n118 B.n117 60.7035
R748 B.n124 B.n123 60.7035
R749 B.n39 B.n38 60.7035
R750 B.n46 B.n45 60.7035
R751 B.n277 B.n118 59.5399
R752 B.n125 B.n124 59.5399
R753 B.n40 B.n39 59.5399
R754 B.n487 B.n46 59.5399
R755 B.n525 B.n524 34.1859
R756 B.n464 B.n463 34.1859
R757 B.n301 B.n300 34.1859
R758 B.n240 B.n133 34.1859
R759 B B.n607 18.0485
R760 B.n524 B.n523 10.6151
R761 B.n523 B.n30 10.6151
R762 B.n519 B.n30 10.6151
R763 B.n519 B.n518 10.6151
R764 B.n518 B.n517 10.6151
R765 B.n517 B.n32 10.6151
R766 B.n513 B.n32 10.6151
R767 B.n513 B.n512 10.6151
R768 B.n512 B.n511 10.6151
R769 B.n511 B.n34 10.6151
R770 B.n507 B.n34 10.6151
R771 B.n507 B.n506 10.6151
R772 B.n506 B.n505 10.6151
R773 B.n505 B.n36 10.6151
R774 B.n501 B.n500 10.6151
R775 B.n500 B.n499 10.6151
R776 B.n499 B.n41 10.6151
R777 B.n495 B.n41 10.6151
R778 B.n495 B.n494 10.6151
R779 B.n494 B.n493 10.6151
R780 B.n493 B.n43 10.6151
R781 B.n489 B.n43 10.6151
R782 B.n489 B.n488 10.6151
R783 B.n486 B.n47 10.6151
R784 B.n482 B.n47 10.6151
R785 B.n482 B.n481 10.6151
R786 B.n481 B.n480 10.6151
R787 B.n480 B.n49 10.6151
R788 B.n476 B.n49 10.6151
R789 B.n476 B.n475 10.6151
R790 B.n475 B.n474 10.6151
R791 B.n474 B.n51 10.6151
R792 B.n470 B.n51 10.6151
R793 B.n470 B.n469 10.6151
R794 B.n469 B.n468 10.6151
R795 B.n468 B.n53 10.6151
R796 B.n464 B.n53 10.6151
R797 B.n302 B.n301 10.6151
R798 B.n302 B.n107 10.6151
R799 B.n306 B.n107 10.6151
R800 B.n307 B.n306 10.6151
R801 B.n308 B.n307 10.6151
R802 B.n308 B.n105 10.6151
R803 B.n312 B.n105 10.6151
R804 B.n313 B.n312 10.6151
R805 B.n314 B.n313 10.6151
R806 B.n314 B.n103 10.6151
R807 B.n318 B.n103 10.6151
R808 B.n319 B.n318 10.6151
R809 B.n320 B.n319 10.6151
R810 B.n320 B.n101 10.6151
R811 B.n324 B.n101 10.6151
R812 B.n325 B.n324 10.6151
R813 B.n326 B.n325 10.6151
R814 B.n326 B.n99 10.6151
R815 B.n330 B.n99 10.6151
R816 B.n331 B.n330 10.6151
R817 B.n332 B.n331 10.6151
R818 B.n332 B.n97 10.6151
R819 B.n336 B.n97 10.6151
R820 B.n337 B.n336 10.6151
R821 B.n338 B.n337 10.6151
R822 B.n338 B.n95 10.6151
R823 B.n342 B.n95 10.6151
R824 B.n343 B.n342 10.6151
R825 B.n344 B.n343 10.6151
R826 B.n344 B.n93 10.6151
R827 B.n348 B.n93 10.6151
R828 B.n349 B.n348 10.6151
R829 B.n350 B.n349 10.6151
R830 B.n350 B.n91 10.6151
R831 B.n354 B.n91 10.6151
R832 B.n355 B.n354 10.6151
R833 B.n356 B.n355 10.6151
R834 B.n356 B.n89 10.6151
R835 B.n360 B.n89 10.6151
R836 B.n361 B.n360 10.6151
R837 B.n362 B.n361 10.6151
R838 B.n362 B.n87 10.6151
R839 B.n366 B.n87 10.6151
R840 B.n367 B.n366 10.6151
R841 B.n368 B.n367 10.6151
R842 B.n368 B.n85 10.6151
R843 B.n372 B.n85 10.6151
R844 B.n373 B.n372 10.6151
R845 B.n374 B.n373 10.6151
R846 B.n374 B.n83 10.6151
R847 B.n378 B.n83 10.6151
R848 B.n379 B.n378 10.6151
R849 B.n380 B.n379 10.6151
R850 B.n380 B.n81 10.6151
R851 B.n384 B.n81 10.6151
R852 B.n385 B.n384 10.6151
R853 B.n386 B.n385 10.6151
R854 B.n386 B.n79 10.6151
R855 B.n390 B.n79 10.6151
R856 B.n391 B.n390 10.6151
R857 B.n392 B.n391 10.6151
R858 B.n392 B.n77 10.6151
R859 B.n396 B.n77 10.6151
R860 B.n397 B.n396 10.6151
R861 B.n398 B.n397 10.6151
R862 B.n398 B.n75 10.6151
R863 B.n402 B.n75 10.6151
R864 B.n403 B.n402 10.6151
R865 B.n404 B.n403 10.6151
R866 B.n404 B.n73 10.6151
R867 B.n408 B.n73 10.6151
R868 B.n409 B.n408 10.6151
R869 B.n410 B.n409 10.6151
R870 B.n410 B.n71 10.6151
R871 B.n414 B.n71 10.6151
R872 B.n415 B.n414 10.6151
R873 B.n416 B.n415 10.6151
R874 B.n416 B.n69 10.6151
R875 B.n420 B.n69 10.6151
R876 B.n421 B.n420 10.6151
R877 B.n422 B.n421 10.6151
R878 B.n422 B.n67 10.6151
R879 B.n426 B.n67 10.6151
R880 B.n427 B.n426 10.6151
R881 B.n428 B.n427 10.6151
R882 B.n428 B.n65 10.6151
R883 B.n432 B.n65 10.6151
R884 B.n433 B.n432 10.6151
R885 B.n434 B.n433 10.6151
R886 B.n434 B.n63 10.6151
R887 B.n438 B.n63 10.6151
R888 B.n439 B.n438 10.6151
R889 B.n440 B.n439 10.6151
R890 B.n440 B.n61 10.6151
R891 B.n444 B.n61 10.6151
R892 B.n445 B.n444 10.6151
R893 B.n446 B.n445 10.6151
R894 B.n446 B.n59 10.6151
R895 B.n450 B.n59 10.6151
R896 B.n451 B.n450 10.6151
R897 B.n452 B.n451 10.6151
R898 B.n452 B.n57 10.6151
R899 B.n456 B.n57 10.6151
R900 B.n457 B.n456 10.6151
R901 B.n458 B.n457 10.6151
R902 B.n458 B.n55 10.6151
R903 B.n462 B.n55 10.6151
R904 B.n463 B.n462 10.6151
R905 B.n241 B.n240 10.6151
R906 B.n242 B.n241 10.6151
R907 B.n242 B.n131 10.6151
R908 B.n246 B.n131 10.6151
R909 B.n247 B.n246 10.6151
R910 B.n248 B.n247 10.6151
R911 B.n248 B.n129 10.6151
R912 B.n252 B.n129 10.6151
R913 B.n253 B.n252 10.6151
R914 B.n254 B.n253 10.6151
R915 B.n254 B.n127 10.6151
R916 B.n258 B.n127 10.6151
R917 B.n259 B.n258 10.6151
R918 B.n260 B.n259 10.6151
R919 B.n264 B.n263 10.6151
R920 B.n265 B.n264 10.6151
R921 B.n265 B.n121 10.6151
R922 B.n269 B.n121 10.6151
R923 B.n270 B.n269 10.6151
R924 B.n271 B.n270 10.6151
R925 B.n271 B.n119 10.6151
R926 B.n275 B.n119 10.6151
R927 B.n276 B.n275 10.6151
R928 B.n278 B.n115 10.6151
R929 B.n282 B.n115 10.6151
R930 B.n283 B.n282 10.6151
R931 B.n284 B.n283 10.6151
R932 B.n284 B.n113 10.6151
R933 B.n288 B.n113 10.6151
R934 B.n289 B.n288 10.6151
R935 B.n290 B.n289 10.6151
R936 B.n290 B.n111 10.6151
R937 B.n294 B.n111 10.6151
R938 B.n295 B.n294 10.6151
R939 B.n296 B.n295 10.6151
R940 B.n296 B.n109 10.6151
R941 B.n300 B.n109 10.6151
R942 B.n236 B.n133 10.6151
R943 B.n236 B.n235 10.6151
R944 B.n235 B.n234 10.6151
R945 B.n234 B.n135 10.6151
R946 B.n230 B.n135 10.6151
R947 B.n230 B.n229 10.6151
R948 B.n229 B.n228 10.6151
R949 B.n228 B.n137 10.6151
R950 B.n224 B.n137 10.6151
R951 B.n224 B.n223 10.6151
R952 B.n223 B.n222 10.6151
R953 B.n222 B.n139 10.6151
R954 B.n218 B.n139 10.6151
R955 B.n218 B.n217 10.6151
R956 B.n217 B.n216 10.6151
R957 B.n216 B.n141 10.6151
R958 B.n212 B.n141 10.6151
R959 B.n212 B.n211 10.6151
R960 B.n211 B.n210 10.6151
R961 B.n210 B.n143 10.6151
R962 B.n206 B.n143 10.6151
R963 B.n206 B.n205 10.6151
R964 B.n205 B.n204 10.6151
R965 B.n204 B.n145 10.6151
R966 B.n200 B.n145 10.6151
R967 B.n200 B.n199 10.6151
R968 B.n199 B.n198 10.6151
R969 B.n198 B.n147 10.6151
R970 B.n194 B.n147 10.6151
R971 B.n194 B.n193 10.6151
R972 B.n193 B.n192 10.6151
R973 B.n192 B.n149 10.6151
R974 B.n188 B.n149 10.6151
R975 B.n188 B.n187 10.6151
R976 B.n187 B.n186 10.6151
R977 B.n186 B.n151 10.6151
R978 B.n182 B.n151 10.6151
R979 B.n182 B.n181 10.6151
R980 B.n181 B.n180 10.6151
R981 B.n180 B.n153 10.6151
R982 B.n176 B.n153 10.6151
R983 B.n176 B.n175 10.6151
R984 B.n175 B.n174 10.6151
R985 B.n174 B.n155 10.6151
R986 B.n170 B.n155 10.6151
R987 B.n170 B.n169 10.6151
R988 B.n169 B.n168 10.6151
R989 B.n168 B.n157 10.6151
R990 B.n164 B.n157 10.6151
R991 B.n164 B.n163 10.6151
R992 B.n163 B.n162 10.6151
R993 B.n162 B.n159 10.6151
R994 B.n159 B.n0 10.6151
R995 B.n603 B.n1 10.6151
R996 B.n603 B.n602 10.6151
R997 B.n602 B.n601 10.6151
R998 B.n601 B.n4 10.6151
R999 B.n597 B.n4 10.6151
R1000 B.n597 B.n596 10.6151
R1001 B.n596 B.n595 10.6151
R1002 B.n595 B.n6 10.6151
R1003 B.n591 B.n6 10.6151
R1004 B.n591 B.n590 10.6151
R1005 B.n590 B.n589 10.6151
R1006 B.n589 B.n8 10.6151
R1007 B.n585 B.n8 10.6151
R1008 B.n585 B.n584 10.6151
R1009 B.n584 B.n583 10.6151
R1010 B.n583 B.n10 10.6151
R1011 B.n579 B.n10 10.6151
R1012 B.n579 B.n578 10.6151
R1013 B.n578 B.n577 10.6151
R1014 B.n577 B.n12 10.6151
R1015 B.n573 B.n12 10.6151
R1016 B.n573 B.n572 10.6151
R1017 B.n572 B.n571 10.6151
R1018 B.n571 B.n14 10.6151
R1019 B.n567 B.n14 10.6151
R1020 B.n567 B.n566 10.6151
R1021 B.n566 B.n565 10.6151
R1022 B.n565 B.n16 10.6151
R1023 B.n561 B.n16 10.6151
R1024 B.n561 B.n560 10.6151
R1025 B.n560 B.n559 10.6151
R1026 B.n559 B.n18 10.6151
R1027 B.n555 B.n18 10.6151
R1028 B.n555 B.n554 10.6151
R1029 B.n554 B.n553 10.6151
R1030 B.n553 B.n20 10.6151
R1031 B.n549 B.n20 10.6151
R1032 B.n549 B.n548 10.6151
R1033 B.n548 B.n547 10.6151
R1034 B.n547 B.n22 10.6151
R1035 B.n543 B.n22 10.6151
R1036 B.n543 B.n542 10.6151
R1037 B.n542 B.n541 10.6151
R1038 B.n541 B.n24 10.6151
R1039 B.n537 B.n24 10.6151
R1040 B.n537 B.n536 10.6151
R1041 B.n536 B.n535 10.6151
R1042 B.n535 B.n26 10.6151
R1043 B.n531 B.n26 10.6151
R1044 B.n531 B.n530 10.6151
R1045 B.n530 B.n529 10.6151
R1046 B.n529 B.n28 10.6151
R1047 B.n525 B.n28 10.6151
R1048 B.n40 B.n36 9.36635
R1049 B.n487 B.n486 9.36635
R1050 B.n260 B.n125 9.36635
R1051 B.n278 B.n277 9.36635
R1052 B.n607 B.n0 2.81026
R1053 B.n607 B.n1 2.81026
R1054 B.n501 B.n40 1.24928
R1055 B.n488 B.n487 1.24928
R1056 B.n263 B.n125 1.24928
R1057 B.n277 B.n276 1.24928
R1058 VP.n19 VP.n16 161.3
R1059 VP.n21 VP.n20 161.3
R1060 VP.n22 VP.n15 161.3
R1061 VP.n24 VP.n23 161.3
R1062 VP.n25 VP.n14 161.3
R1063 VP.n27 VP.n26 161.3
R1064 VP.n29 VP.n13 161.3
R1065 VP.n31 VP.n30 161.3
R1066 VP.n32 VP.n12 161.3
R1067 VP.n34 VP.n33 161.3
R1068 VP.n35 VP.n11 161.3
R1069 VP.n37 VP.n36 161.3
R1070 VP.n69 VP.n68 161.3
R1071 VP.n67 VP.n1 161.3
R1072 VP.n66 VP.n65 161.3
R1073 VP.n64 VP.n2 161.3
R1074 VP.n63 VP.n62 161.3
R1075 VP.n61 VP.n3 161.3
R1076 VP.n59 VP.n58 161.3
R1077 VP.n57 VP.n4 161.3
R1078 VP.n56 VP.n55 161.3
R1079 VP.n54 VP.n5 161.3
R1080 VP.n53 VP.n52 161.3
R1081 VP.n51 VP.n6 161.3
R1082 VP.n50 VP.n49 161.3
R1083 VP.n47 VP.n7 161.3
R1084 VP.n46 VP.n45 161.3
R1085 VP.n44 VP.n8 161.3
R1086 VP.n43 VP.n42 161.3
R1087 VP.n41 VP.n9 161.3
R1088 VP.n40 VP.n39 68.2918
R1089 VP.n70 VP.n0 68.2918
R1090 VP.n38 VP.n10 68.2918
R1091 VP.n18 VP.n17 58.2302
R1092 VP.n18 VP.t6 57.9635
R1093 VP.n55 VP.n54 56.5193
R1094 VP.n23 VP.n22 56.5193
R1095 VP.n46 VP.n8 52.1486
R1096 VP.n66 VP.n2 52.1486
R1097 VP.n34 VP.n12 52.1486
R1098 VP.n39 VP.n38 45.1357
R1099 VP.n42 VP.n8 28.8382
R1100 VP.n67 VP.n66 28.8382
R1101 VP.n35 VP.n34 28.8382
R1102 VP.n40 VP.t3 26.0801
R1103 VP.n48 VP.t0 26.0801
R1104 VP.n60 VP.t4 26.0801
R1105 VP.n0 VP.t2 26.0801
R1106 VP.n10 VP.t5 26.0801
R1107 VP.n28 VP.t7 26.0801
R1108 VP.n17 VP.t1 26.0801
R1109 VP.n42 VP.n41 24.4675
R1110 VP.n47 VP.n46 24.4675
R1111 VP.n49 VP.n47 24.4675
R1112 VP.n53 VP.n6 24.4675
R1113 VP.n54 VP.n53 24.4675
R1114 VP.n55 VP.n4 24.4675
R1115 VP.n59 VP.n4 24.4675
R1116 VP.n62 VP.n61 24.4675
R1117 VP.n62 VP.n2 24.4675
R1118 VP.n68 VP.n67 24.4675
R1119 VP.n36 VP.n35 24.4675
R1120 VP.n23 VP.n14 24.4675
R1121 VP.n27 VP.n14 24.4675
R1122 VP.n30 VP.n29 24.4675
R1123 VP.n30 VP.n12 24.4675
R1124 VP.n21 VP.n16 24.4675
R1125 VP.n22 VP.n21 24.4675
R1126 VP.n41 VP.n40 21.7761
R1127 VP.n68 VP.n0 21.7761
R1128 VP.n36 VP.n10 21.7761
R1129 VP.n48 VP.n6 15.4147
R1130 VP.n60 VP.n59 15.4147
R1131 VP.n28 VP.n27 15.4147
R1132 VP.n17 VP.n16 15.4147
R1133 VP.n49 VP.n48 9.05329
R1134 VP.n61 VP.n60 9.05329
R1135 VP.n29 VP.n28 9.05329
R1136 VP.n19 VP.n18 5.40752
R1137 VP.n38 VP.n37 0.354971
R1138 VP.n39 VP.n9 0.354971
R1139 VP.n70 VP.n69 0.354971
R1140 VP VP.n70 0.26696
R1141 VP.n20 VP.n19 0.189894
R1142 VP.n20 VP.n15 0.189894
R1143 VP.n24 VP.n15 0.189894
R1144 VP.n25 VP.n24 0.189894
R1145 VP.n26 VP.n25 0.189894
R1146 VP.n26 VP.n13 0.189894
R1147 VP.n31 VP.n13 0.189894
R1148 VP.n32 VP.n31 0.189894
R1149 VP.n33 VP.n32 0.189894
R1150 VP.n33 VP.n11 0.189894
R1151 VP.n37 VP.n11 0.189894
R1152 VP.n43 VP.n9 0.189894
R1153 VP.n44 VP.n43 0.189894
R1154 VP.n45 VP.n44 0.189894
R1155 VP.n45 VP.n7 0.189894
R1156 VP.n50 VP.n7 0.189894
R1157 VP.n51 VP.n50 0.189894
R1158 VP.n52 VP.n51 0.189894
R1159 VP.n52 VP.n5 0.189894
R1160 VP.n56 VP.n5 0.189894
R1161 VP.n57 VP.n56 0.189894
R1162 VP.n58 VP.n57 0.189894
R1163 VP.n58 VP.n3 0.189894
R1164 VP.n63 VP.n3 0.189894
R1165 VP.n64 VP.n63 0.189894
R1166 VP.n65 VP.n64 0.189894
R1167 VP.n65 VP.n1 0.189894
R1168 VP.n69 VP.n1 0.189894
R1169 VDD1 VDD1.n0 138.952
R1170 VDD1.n3 VDD1.n2 138.838
R1171 VDD1.n3 VDD1.n1 138.838
R1172 VDD1.n5 VDD1.n4 137.543
R1173 VDD1.n5 VDD1.n3 39.0526
R1174 VDD1.n4 VDD1.t0 10.7282
R1175 VDD1.n4 VDD1.t2 10.7282
R1176 VDD1.n0 VDD1.t1 10.7282
R1177 VDD1.n0 VDD1.t6 10.7282
R1178 VDD1.n2 VDD1.t3 10.7282
R1179 VDD1.n2 VDD1.t5 10.7282
R1180 VDD1.n1 VDD1.t4 10.7282
R1181 VDD1.n1 VDD1.t7 10.7282
R1182 VDD1 VDD1.n5 1.29145
C0 VDD2 B 1.56986f
C1 VN VDD1 0.156954f
C2 VDD1 VP 2.95703f
C3 VN w_n4100_n1574# 8.253691f
C4 VP w_n4100_n1574# 8.784269f
C5 B VTAIL 2.03196f
C6 VN VDD2 2.56987f
C7 VDD2 VP 0.546664f
C8 VDD1 w_n4100_n1574# 1.77567f
C9 VN VTAIL 3.68258f
C10 VP VTAIL 3.69668f
C11 VDD1 VDD2 1.88109f
C12 VDD2 w_n4100_n1574# 1.89827f
C13 VN B 1.18399f
C14 B VP 2.07788f
C15 VDD1 VTAIL 5.2257f
C16 w_n4100_n1574# VTAIL 2.19808f
C17 VDD1 B 1.46731f
C18 B w_n4100_n1574# 7.94263f
C19 VN VP 6.25674f
C20 VDD2 VTAIL 5.28146f
C21 VDD2 VSUBS 1.491013f
C22 VDD1 VSUBS 2.188208f
C23 VTAIL VSUBS 0.636999f
C24 VN VSUBS 6.94403f
C25 VP VSUBS 3.2206f
C26 B VSUBS 4.202252f
C27 w_n4100_n1574# VSUBS 81.72121f
C28 VDD1.t1 VSUBS 0.059681f
C29 VDD1.t6 VSUBS 0.059681f
C30 VDD1.n0 VSUBS 0.308363f
C31 VDD1.t4 VSUBS 0.059681f
C32 VDD1.t7 VSUBS 0.059681f
C33 VDD1.n1 VSUBS 0.307739f
C34 VDD1.t3 VSUBS 0.059681f
C35 VDD1.t5 VSUBS 0.059681f
C36 VDD1.n2 VSUBS 0.307739f
C37 VDD1.n3 VSUBS 3.14618f
C38 VDD1.t0 VSUBS 0.059681f
C39 VDD1.t2 VSUBS 0.059681f
C40 VDD1.n4 VSUBS 0.301582f
C41 VDD1.n5 VSUBS 2.47152f
C42 VP.t2 VSUBS 1.10629f
C43 VP.n0 VSUBS 0.663033f
C44 VP.n1 VSUBS 0.052281f
C45 VP.n2 VSUBS 0.093859f
C46 VP.n3 VSUBS 0.052281f
C47 VP.t4 VSUBS 1.10629f
C48 VP.n4 VSUBS 0.097438f
C49 VP.n5 VSUBS 0.052281f
C50 VP.n6 VSUBS 0.079637f
C51 VP.n7 VSUBS 0.052281f
C52 VP.n8 VSUBS 0.052807f
C53 VP.n9 VSUBS 0.08438f
C54 VP.t3 VSUBS 1.10629f
C55 VP.t5 VSUBS 1.10629f
C56 VP.n10 VSUBS 0.663033f
C57 VP.n11 VSUBS 0.052281f
C58 VP.n12 VSUBS 0.093859f
C59 VP.n13 VSUBS 0.052281f
C60 VP.t7 VSUBS 1.10629f
C61 VP.n14 VSUBS 0.097438f
C62 VP.n15 VSUBS 0.052281f
C63 VP.n16 VSUBS 0.079637f
C64 VP.t6 VSUBS 1.54717f
C65 VP.t1 VSUBS 1.10629f
C66 VP.n17 VSUBS 0.628965f
C67 VP.n18 VSUBS 0.60694f
C68 VP.n19 VSUBS 0.551608f
C69 VP.n20 VSUBS 0.052281f
C70 VP.n21 VSUBS 0.097438f
C71 VP.n22 VSUBS 0.07632f
C72 VP.n23 VSUBS 0.07632f
C73 VP.n24 VSUBS 0.052281f
C74 VP.n25 VSUBS 0.052281f
C75 VP.n26 VSUBS 0.052281f
C76 VP.n27 VSUBS 0.079637f
C77 VP.n28 VSUBS 0.462446f
C78 VP.n29 VSUBS 0.067129f
C79 VP.n30 VSUBS 0.097438f
C80 VP.n31 VSUBS 0.052281f
C81 VP.n32 VSUBS 0.052281f
C82 VP.n33 VSUBS 0.052281f
C83 VP.n34 VSUBS 0.052807f
C84 VP.n35 VSUBS 0.103414f
C85 VP.n36 VSUBS 0.092144f
C86 VP.n37 VSUBS 0.08438f
C87 VP.n38 VSUBS 2.52939f
C88 VP.n39 VSUBS 2.57102f
C89 VP.n40 VSUBS 0.663033f
C90 VP.n41 VSUBS 0.092144f
C91 VP.n42 VSUBS 0.103414f
C92 VP.n43 VSUBS 0.052281f
C93 VP.n44 VSUBS 0.052281f
C94 VP.n45 VSUBS 0.052281f
C95 VP.n46 VSUBS 0.093859f
C96 VP.n47 VSUBS 0.097438f
C97 VP.t0 VSUBS 1.10629f
C98 VP.n48 VSUBS 0.462446f
C99 VP.n49 VSUBS 0.067129f
C100 VP.n50 VSUBS 0.052281f
C101 VP.n51 VSUBS 0.052281f
C102 VP.n52 VSUBS 0.052281f
C103 VP.n53 VSUBS 0.097438f
C104 VP.n54 VSUBS 0.07632f
C105 VP.n55 VSUBS 0.07632f
C106 VP.n56 VSUBS 0.052281f
C107 VP.n57 VSUBS 0.052281f
C108 VP.n58 VSUBS 0.052281f
C109 VP.n59 VSUBS 0.079637f
C110 VP.n60 VSUBS 0.462446f
C111 VP.n61 VSUBS 0.067129f
C112 VP.n62 VSUBS 0.097438f
C113 VP.n63 VSUBS 0.052281f
C114 VP.n64 VSUBS 0.052281f
C115 VP.n65 VSUBS 0.052281f
C116 VP.n66 VSUBS 0.052807f
C117 VP.n67 VSUBS 0.103414f
C118 VP.n68 VSUBS 0.092144f
C119 VP.n69 VSUBS 0.08438f
C120 VP.n70 VSUBS 0.101309f
C121 B.n0 VSUBS 0.007278f
C122 B.n1 VSUBS 0.007278f
C123 B.n2 VSUBS 0.011509f
C124 B.n3 VSUBS 0.011509f
C125 B.n4 VSUBS 0.011509f
C126 B.n5 VSUBS 0.011509f
C127 B.n6 VSUBS 0.011509f
C128 B.n7 VSUBS 0.011509f
C129 B.n8 VSUBS 0.011509f
C130 B.n9 VSUBS 0.011509f
C131 B.n10 VSUBS 0.011509f
C132 B.n11 VSUBS 0.011509f
C133 B.n12 VSUBS 0.011509f
C134 B.n13 VSUBS 0.011509f
C135 B.n14 VSUBS 0.011509f
C136 B.n15 VSUBS 0.011509f
C137 B.n16 VSUBS 0.011509f
C138 B.n17 VSUBS 0.011509f
C139 B.n18 VSUBS 0.011509f
C140 B.n19 VSUBS 0.011509f
C141 B.n20 VSUBS 0.011509f
C142 B.n21 VSUBS 0.011509f
C143 B.n22 VSUBS 0.011509f
C144 B.n23 VSUBS 0.011509f
C145 B.n24 VSUBS 0.011509f
C146 B.n25 VSUBS 0.011509f
C147 B.n26 VSUBS 0.011509f
C148 B.n27 VSUBS 0.011509f
C149 B.n28 VSUBS 0.011509f
C150 B.n29 VSUBS 0.028503f
C151 B.n30 VSUBS 0.011509f
C152 B.n31 VSUBS 0.011509f
C153 B.n32 VSUBS 0.011509f
C154 B.n33 VSUBS 0.011509f
C155 B.n34 VSUBS 0.011509f
C156 B.n35 VSUBS 0.011509f
C157 B.n36 VSUBS 0.010832f
C158 B.n37 VSUBS 0.011509f
C159 B.t2 VSUBS 0.119805f
C160 B.t1 VSUBS 0.147141f
C161 B.t0 VSUBS 0.679427f
C162 B.n38 VSUBS 0.138289f
C163 B.n39 VSUBS 0.10936f
C164 B.n40 VSUBS 0.026666f
C165 B.n41 VSUBS 0.011509f
C166 B.n42 VSUBS 0.011509f
C167 B.n43 VSUBS 0.011509f
C168 B.n44 VSUBS 0.011509f
C169 B.t8 VSUBS 0.119805f
C170 B.t7 VSUBS 0.147141f
C171 B.t6 VSUBS 0.679427f
C172 B.n45 VSUBS 0.13829f
C173 B.n46 VSUBS 0.10936f
C174 B.n47 VSUBS 0.011509f
C175 B.n48 VSUBS 0.011509f
C176 B.n49 VSUBS 0.011509f
C177 B.n50 VSUBS 0.011509f
C178 B.n51 VSUBS 0.011509f
C179 B.n52 VSUBS 0.011509f
C180 B.n53 VSUBS 0.011509f
C181 B.n54 VSUBS 0.027014f
C182 B.n55 VSUBS 0.011509f
C183 B.n56 VSUBS 0.011509f
C184 B.n57 VSUBS 0.011509f
C185 B.n58 VSUBS 0.011509f
C186 B.n59 VSUBS 0.011509f
C187 B.n60 VSUBS 0.011509f
C188 B.n61 VSUBS 0.011509f
C189 B.n62 VSUBS 0.011509f
C190 B.n63 VSUBS 0.011509f
C191 B.n64 VSUBS 0.011509f
C192 B.n65 VSUBS 0.011509f
C193 B.n66 VSUBS 0.011509f
C194 B.n67 VSUBS 0.011509f
C195 B.n68 VSUBS 0.011509f
C196 B.n69 VSUBS 0.011509f
C197 B.n70 VSUBS 0.011509f
C198 B.n71 VSUBS 0.011509f
C199 B.n72 VSUBS 0.011509f
C200 B.n73 VSUBS 0.011509f
C201 B.n74 VSUBS 0.011509f
C202 B.n75 VSUBS 0.011509f
C203 B.n76 VSUBS 0.011509f
C204 B.n77 VSUBS 0.011509f
C205 B.n78 VSUBS 0.011509f
C206 B.n79 VSUBS 0.011509f
C207 B.n80 VSUBS 0.011509f
C208 B.n81 VSUBS 0.011509f
C209 B.n82 VSUBS 0.011509f
C210 B.n83 VSUBS 0.011509f
C211 B.n84 VSUBS 0.011509f
C212 B.n85 VSUBS 0.011509f
C213 B.n86 VSUBS 0.011509f
C214 B.n87 VSUBS 0.011509f
C215 B.n88 VSUBS 0.011509f
C216 B.n89 VSUBS 0.011509f
C217 B.n90 VSUBS 0.011509f
C218 B.n91 VSUBS 0.011509f
C219 B.n92 VSUBS 0.011509f
C220 B.n93 VSUBS 0.011509f
C221 B.n94 VSUBS 0.011509f
C222 B.n95 VSUBS 0.011509f
C223 B.n96 VSUBS 0.011509f
C224 B.n97 VSUBS 0.011509f
C225 B.n98 VSUBS 0.011509f
C226 B.n99 VSUBS 0.011509f
C227 B.n100 VSUBS 0.011509f
C228 B.n101 VSUBS 0.011509f
C229 B.n102 VSUBS 0.011509f
C230 B.n103 VSUBS 0.011509f
C231 B.n104 VSUBS 0.011509f
C232 B.n105 VSUBS 0.011509f
C233 B.n106 VSUBS 0.011509f
C234 B.n107 VSUBS 0.011509f
C235 B.n108 VSUBS 0.027014f
C236 B.n109 VSUBS 0.011509f
C237 B.n110 VSUBS 0.011509f
C238 B.n111 VSUBS 0.011509f
C239 B.n112 VSUBS 0.011509f
C240 B.n113 VSUBS 0.011509f
C241 B.n114 VSUBS 0.011509f
C242 B.n115 VSUBS 0.011509f
C243 B.n116 VSUBS 0.011509f
C244 B.t4 VSUBS 0.119805f
C245 B.t5 VSUBS 0.147141f
C246 B.t3 VSUBS 0.679427f
C247 B.n117 VSUBS 0.13829f
C248 B.n118 VSUBS 0.10936f
C249 B.n119 VSUBS 0.011509f
C250 B.n120 VSUBS 0.011509f
C251 B.n121 VSUBS 0.011509f
C252 B.n122 VSUBS 0.011509f
C253 B.t10 VSUBS 0.119805f
C254 B.t11 VSUBS 0.147141f
C255 B.t9 VSUBS 0.679427f
C256 B.n123 VSUBS 0.138289f
C257 B.n124 VSUBS 0.10936f
C258 B.n125 VSUBS 0.026666f
C259 B.n126 VSUBS 0.011509f
C260 B.n127 VSUBS 0.011509f
C261 B.n128 VSUBS 0.011509f
C262 B.n129 VSUBS 0.011509f
C263 B.n130 VSUBS 0.011509f
C264 B.n131 VSUBS 0.011509f
C265 B.n132 VSUBS 0.011509f
C266 B.n133 VSUBS 0.027014f
C267 B.n134 VSUBS 0.011509f
C268 B.n135 VSUBS 0.011509f
C269 B.n136 VSUBS 0.011509f
C270 B.n137 VSUBS 0.011509f
C271 B.n138 VSUBS 0.011509f
C272 B.n139 VSUBS 0.011509f
C273 B.n140 VSUBS 0.011509f
C274 B.n141 VSUBS 0.011509f
C275 B.n142 VSUBS 0.011509f
C276 B.n143 VSUBS 0.011509f
C277 B.n144 VSUBS 0.011509f
C278 B.n145 VSUBS 0.011509f
C279 B.n146 VSUBS 0.011509f
C280 B.n147 VSUBS 0.011509f
C281 B.n148 VSUBS 0.011509f
C282 B.n149 VSUBS 0.011509f
C283 B.n150 VSUBS 0.011509f
C284 B.n151 VSUBS 0.011509f
C285 B.n152 VSUBS 0.011509f
C286 B.n153 VSUBS 0.011509f
C287 B.n154 VSUBS 0.011509f
C288 B.n155 VSUBS 0.011509f
C289 B.n156 VSUBS 0.011509f
C290 B.n157 VSUBS 0.011509f
C291 B.n158 VSUBS 0.011509f
C292 B.n159 VSUBS 0.011509f
C293 B.n160 VSUBS 0.011509f
C294 B.n161 VSUBS 0.011509f
C295 B.n162 VSUBS 0.011509f
C296 B.n163 VSUBS 0.011509f
C297 B.n164 VSUBS 0.011509f
C298 B.n165 VSUBS 0.011509f
C299 B.n166 VSUBS 0.011509f
C300 B.n167 VSUBS 0.011509f
C301 B.n168 VSUBS 0.011509f
C302 B.n169 VSUBS 0.011509f
C303 B.n170 VSUBS 0.011509f
C304 B.n171 VSUBS 0.011509f
C305 B.n172 VSUBS 0.011509f
C306 B.n173 VSUBS 0.011509f
C307 B.n174 VSUBS 0.011509f
C308 B.n175 VSUBS 0.011509f
C309 B.n176 VSUBS 0.011509f
C310 B.n177 VSUBS 0.011509f
C311 B.n178 VSUBS 0.011509f
C312 B.n179 VSUBS 0.011509f
C313 B.n180 VSUBS 0.011509f
C314 B.n181 VSUBS 0.011509f
C315 B.n182 VSUBS 0.011509f
C316 B.n183 VSUBS 0.011509f
C317 B.n184 VSUBS 0.011509f
C318 B.n185 VSUBS 0.011509f
C319 B.n186 VSUBS 0.011509f
C320 B.n187 VSUBS 0.011509f
C321 B.n188 VSUBS 0.011509f
C322 B.n189 VSUBS 0.011509f
C323 B.n190 VSUBS 0.011509f
C324 B.n191 VSUBS 0.011509f
C325 B.n192 VSUBS 0.011509f
C326 B.n193 VSUBS 0.011509f
C327 B.n194 VSUBS 0.011509f
C328 B.n195 VSUBS 0.011509f
C329 B.n196 VSUBS 0.011509f
C330 B.n197 VSUBS 0.011509f
C331 B.n198 VSUBS 0.011509f
C332 B.n199 VSUBS 0.011509f
C333 B.n200 VSUBS 0.011509f
C334 B.n201 VSUBS 0.011509f
C335 B.n202 VSUBS 0.011509f
C336 B.n203 VSUBS 0.011509f
C337 B.n204 VSUBS 0.011509f
C338 B.n205 VSUBS 0.011509f
C339 B.n206 VSUBS 0.011509f
C340 B.n207 VSUBS 0.011509f
C341 B.n208 VSUBS 0.011509f
C342 B.n209 VSUBS 0.011509f
C343 B.n210 VSUBS 0.011509f
C344 B.n211 VSUBS 0.011509f
C345 B.n212 VSUBS 0.011509f
C346 B.n213 VSUBS 0.011509f
C347 B.n214 VSUBS 0.011509f
C348 B.n215 VSUBS 0.011509f
C349 B.n216 VSUBS 0.011509f
C350 B.n217 VSUBS 0.011509f
C351 B.n218 VSUBS 0.011509f
C352 B.n219 VSUBS 0.011509f
C353 B.n220 VSUBS 0.011509f
C354 B.n221 VSUBS 0.011509f
C355 B.n222 VSUBS 0.011509f
C356 B.n223 VSUBS 0.011509f
C357 B.n224 VSUBS 0.011509f
C358 B.n225 VSUBS 0.011509f
C359 B.n226 VSUBS 0.011509f
C360 B.n227 VSUBS 0.011509f
C361 B.n228 VSUBS 0.011509f
C362 B.n229 VSUBS 0.011509f
C363 B.n230 VSUBS 0.011509f
C364 B.n231 VSUBS 0.011509f
C365 B.n232 VSUBS 0.011509f
C366 B.n233 VSUBS 0.011509f
C367 B.n234 VSUBS 0.011509f
C368 B.n235 VSUBS 0.011509f
C369 B.n236 VSUBS 0.011509f
C370 B.n237 VSUBS 0.011509f
C371 B.n238 VSUBS 0.027014f
C372 B.n239 VSUBS 0.028503f
C373 B.n240 VSUBS 0.028503f
C374 B.n241 VSUBS 0.011509f
C375 B.n242 VSUBS 0.011509f
C376 B.n243 VSUBS 0.011509f
C377 B.n244 VSUBS 0.011509f
C378 B.n245 VSUBS 0.011509f
C379 B.n246 VSUBS 0.011509f
C380 B.n247 VSUBS 0.011509f
C381 B.n248 VSUBS 0.011509f
C382 B.n249 VSUBS 0.011509f
C383 B.n250 VSUBS 0.011509f
C384 B.n251 VSUBS 0.011509f
C385 B.n252 VSUBS 0.011509f
C386 B.n253 VSUBS 0.011509f
C387 B.n254 VSUBS 0.011509f
C388 B.n255 VSUBS 0.011509f
C389 B.n256 VSUBS 0.011509f
C390 B.n257 VSUBS 0.011509f
C391 B.n258 VSUBS 0.011509f
C392 B.n259 VSUBS 0.011509f
C393 B.n260 VSUBS 0.010832f
C394 B.n261 VSUBS 0.011509f
C395 B.n262 VSUBS 0.011509f
C396 B.n263 VSUBS 0.006432f
C397 B.n264 VSUBS 0.011509f
C398 B.n265 VSUBS 0.011509f
C399 B.n266 VSUBS 0.011509f
C400 B.n267 VSUBS 0.011509f
C401 B.n268 VSUBS 0.011509f
C402 B.n269 VSUBS 0.011509f
C403 B.n270 VSUBS 0.011509f
C404 B.n271 VSUBS 0.011509f
C405 B.n272 VSUBS 0.011509f
C406 B.n273 VSUBS 0.011509f
C407 B.n274 VSUBS 0.011509f
C408 B.n275 VSUBS 0.011509f
C409 B.n276 VSUBS 0.006432f
C410 B.n277 VSUBS 0.026666f
C411 B.n278 VSUBS 0.010832f
C412 B.n279 VSUBS 0.011509f
C413 B.n280 VSUBS 0.011509f
C414 B.n281 VSUBS 0.011509f
C415 B.n282 VSUBS 0.011509f
C416 B.n283 VSUBS 0.011509f
C417 B.n284 VSUBS 0.011509f
C418 B.n285 VSUBS 0.011509f
C419 B.n286 VSUBS 0.011509f
C420 B.n287 VSUBS 0.011509f
C421 B.n288 VSUBS 0.011509f
C422 B.n289 VSUBS 0.011509f
C423 B.n290 VSUBS 0.011509f
C424 B.n291 VSUBS 0.011509f
C425 B.n292 VSUBS 0.011509f
C426 B.n293 VSUBS 0.011509f
C427 B.n294 VSUBS 0.011509f
C428 B.n295 VSUBS 0.011509f
C429 B.n296 VSUBS 0.011509f
C430 B.n297 VSUBS 0.011509f
C431 B.n298 VSUBS 0.011509f
C432 B.n299 VSUBS 0.028503f
C433 B.n300 VSUBS 0.028503f
C434 B.n301 VSUBS 0.027014f
C435 B.n302 VSUBS 0.011509f
C436 B.n303 VSUBS 0.011509f
C437 B.n304 VSUBS 0.011509f
C438 B.n305 VSUBS 0.011509f
C439 B.n306 VSUBS 0.011509f
C440 B.n307 VSUBS 0.011509f
C441 B.n308 VSUBS 0.011509f
C442 B.n309 VSUBS 0.011509f
C443 B.n310 VSUBS 0.011509f
C444 B.n311 VSUBS 0.011509f
C445 B.n312 VSUBS 0.011509f
C446 B.n313 VSUBS 0.011509f
C447 B.n314 VSUBS 0.011509f
C448 B.n315 VSUBS 0.011509f
C449 B.n316 VSUBS 0.011509f
C450 B.n317 VSUBS 0.011509f
C451 B.n318 VSUBS 0.011509f
C452 B.n319 VSUBS 0.011509f
C453 B.n320 VSUBS 0.011509f
C454 B.n321 VSUBS 0.011509f
C455 B.n322 VSUBS 0.011509f
C456 B.n323 VSUBS 0.011509f
C457 B.n324 VSUBS 0.011509f
C458 B.n325 VSUBS 0.011509f
C459 B.n326 VSUBS 0.011509f
C460 B.n327 VSUBS 0.011509f
C461 B.n328 VSUBS 0.011509f
C462 B.n329 VSUBS 0.011509f
C463 B.n330 VSUBS 0.011509f
C464 B.n331 VSUBS 0.011509f
C465 B.n332 VSUBS 0.011509f
C466 B.n333 VSUBS 0.011509f
C467 B.n334 VSUBS 0.011509f
C468 B.n335 VSUBS 0.011509f
C469 B.n336 VSUBS 0.011509f
C470 B.n337 VSUBS 0.011509f
C471 B.n338 VSUBS 0.011509f
C472 B.n339 VSUBS 0.011509f
C473 B.n340 VSUBS 0.011509f
C474 B.n341 VSUBS 0.011509f
C475 B.n342 VSUBS 0.011509f
C476 B.n343 VSUBS 0.011509f
C477 B.n344 VSUBS 0.011509f
C478 B.n345 VSUBS 0.011509f
C479 B.n346 VSUBS 0.011509f
C480 B.n347 VSUBS 0.011509f
C481 B.n348 VSUBS 0.011509f
C482 B.n349 VSUBS 0.011509f
C483 B.n350 VSUBS 0.011509f
C484 B.n351 VSUBS 0.011509f
C485 B.n352 VSUBS 0.011509f
C486 B.n353 VSUBS 0.011509f
C487 B.n354 VSUBS 0.011509f
C488 B.n355 VSUBS 0.011509f
C489 B.n356 VSUBS 0.011509f
C490 B.n357 VSUBS 0.011509f
C491 B.n358 VSUBS 0.011509f
C492 B.n359 VSUBS 0.011509f
C493 B.n360 VSUBS 0.011509f
C494 B.n361 VSUBS 0.011509f
C495 B.n362 VSUBS 0.011509f
C496 B.n363 VSUBS 0.011509f
C497 B.n364 VSUBS 0.011509f
C498 B.n365 VSUBS 0.011509f
C499 B.n366 VSUBS 0.011509f
C500 B.n367 VSUBS 0.011509f
C501 B.n368 VSUBS 0.011509f
C502 B.n369 VSUBS 0.011509f
C503 B.n370 VSUBS 0.011509f
C504 B.n371 VSUBS 0.011509f
C505 B.n372 VSUBS 0.011509f
C506 B.n373 VSUBS 0.011509f
C507 B.n374 VSUBS 0.011509f
C508 B.n375 VSUBS 0.011509f
C509 B.n376 VSUBS 0.011509f
C510 B.n377 VSUBS 0.011509f
C511 B.n378 VSUBS 0.011509f
C512 B.n379 VSUBS 0.011509f
C513 B.n380 VSUBS 0.011509f
C514 B.n381 VSUBS 0.011509f
C515 B.n382 VSUBS 0.011509f
C516 B.n383 VSUBS 0.011509f
C517 B.n384 VSUBS 0.011509f
C518 B.n385 VSUBS 0.011509f
C519 B.n386 VSUBS 0.011509f
C520 B.n387 VSUBS 0.011509f
C521 B.n388 VSUBS 0.011509f
C522 B.n389 VSUBS 0.011509f
C523 B.n390 VSUBS 0.011509f
C524 B.n391 VSUBS 0.011509f
C525 B.n392 VSUBS 0.011509f
C526 B.n393 VSUBS 0.011509f
C527 B.n394 VSUBS 0.011509f
C528 B.n395 VSUBS 0.011509f
C529 B.n396 VSUBS 0.011509f
C530 B.n397 VSUBS 0.011509f
C531 B.n398 VSUBS 0.011509f
C532 B.n399 VSUBS 0.011509f
C533 B.n400 VSUBS 0.011509f
C534 B.n401 VSUBS 0.011509f
C535 B.n402 VSUBS 0.011509f
C536 B.n403 VSUBS 0.011509f
C537 B.n404 VSUBS 0.011509f
C538 B.n405 VSUBS 0.011509f
C539 B.n406 VSUBS 0.011509f
C540 B.n407 VSUBS 0.011509f
C541 B.n408 VSUBS 0.011509f
C542 B.n409 VSUBS 0.011509f
C543 B.n410 VSUBS 0.011509f
C544 B.n411 VSUBS 0.011509f
C545 B.n412 VSUBS 0.011509f
C546 B.n413 VSUBS 0.011509f
C547 B.n414 VSUBS 0.011509f
C548 B.n415 VSUBS 0.011509f
C549 B.n416 VSUBS 0.011509f
C550 B.n417 VSUBS 0.011509f
C551 B.n418 VSUBS 0.011509f
C552 B.n419 VSUBS 0.011509f
C553 B.n420 VSUBS 0.011509f
C554 B.n421 VSUBS 0.011509f
C555 B.n422 VSUBS 0.011509f
C556 B.n423 VSUBS 0.011509f
C557 B.n424 VSUBS 0.011509f
C558 B.n425 VSUBS 0.011509f
C559 B.n426 VSUBS 0.011509f
C560 B.n427 VSUBS 0.011509f
C561 B.n428 VSUBS 0.011509f
C562 B.n429 VSUBS 0.011509f
C563 B.n430 VSUBS 0.011509f
C564 B.n431 VSUBS 0.011509f
C565 B.n432 VSUBS 0.011509f
C566 B.n433 VSUBS 0.011509f
C567 B.n434 VSUBS 0.011509f
C568 B.n435 VSUBS 0.011509f
C569 B.n436 VSUBS 0.011509f
C570 B.n437 VSUBS 0.011509f
C571 B.n438 VSUBS 0.011509f
C572 B.n439 VSUBS 0.011509f
C573 B.n440 VSUBS 0.011509f
C574 B.n441 VSUBS 0.011509f
C575 B.n442 VSUBS 0.011509f
C576 B.n443 VSUBS 0.011509f
C577 B.n444 VSUBS 0.011509f
C578 B.n445 VSUBS 0.011509f
C579 B.n446 VSUBS 0.011509f
C580 B.n447 VSUBS 0.011509f
C581 B.n448 VSUBS 0.011509f
C582 B.n449 VSUBS 0.011509f
C583 B.n450 VSUBS 0.011509f
C584 B.n451 VSUBS 0.011509f
C585 B.n452 VSUBS 0.011509f
C586 B.n453 VSUBS 0.011509f
C587 B.n454 VSUBS 0.011509f
C588 B.n455 VSUBS 0.011509f
C589 B.n456 VSUBS 0.011509f
C590 B.n457 VSUBS 0.011509f
C591 B.n458 VSUBS 0.011509f
C592 B.n459 VSUBS 0.011509f
C593 B.n460 VSUBS 0.011509f
C594 B.n461 VSUBS 0.011509f
C595 B.n462 VSUBS 0.011509f
C596 B.n463 VSUBS 0.028313f
C597 B.n464 VSUBS 0.027204f
C598 B.n465 VSUBS 0.028503f
C599 B.n466 VSUBS 0.011509f
C600 B.n467 VSUBS 0.011509f
C601 B.n468 VSUBS 0.011509f
C602 B.n469 VSUBS 0.011509f
C603 B.n470 VSUBS 0.011509f
C604 B.n471 VSUBS 0.011509f
C605 B.n472 VSUBS 0.011509f
C606 B.n473 VSUBS 0.011509f
C607 B.n474 VSUBS 0.011509f
C608 B.n475 VSUBS 0.011509f
C609 B.n476 VSUBS 0.011509f
C610 B.n477 VSUBS 0.011509f
C611 B.n478 VSUBS 0.011509f
C612 B.n479 VSUBS 0.011509f
C613 B.n480 VSUBS 0.011509f
C614 B.n481 VSUBS 0.011509f
C615 B.n482 VSUBS 0.011509f
C616 B.n483 VSUBS 0.011509f
C617 B.n484 VSUBS 0.011509f
C618 B.n485 VSUBS 0.011509f
C619 B.n486 VSUBS 0.010832f
C620 B.n487 VSUBS 0.026666f
C621 B.n488 VSUBS 0.006432f
C622 B.n489 VSUBS 0.011509f
C623 B.n490 VSUBS 0.011509f
C624 B.n491 VSUBS 0.011509f
C625 B.n492 VSUBS 0.011509f
C626 B.n493 VSUBS 0.011509f
C627 B.n494 VSUBS 0.011509f
C628 B.n495 VSUBS 0.011509f
C629 B.n496 VSUBS 0.011509f
C630 B.n497 VSUBS 0.011509f
C631 B.n498 VSUBS 0.011509f
C632 B.n499 VSUBS 0.011509f
C633 B.n500 VSUBS 0.011509f
C634 B.n501 VSUBS 0.006432f
C635 B.n502 VSUBS 0.011509f
C636 B.n503 VSUBS 0.011509f
C637 B.n504 VSUBS 0.011509f
C638 B.n505 VSUBS 0.011509f
C639 B.n506 VSUBS 0.011509f
C640 B.n507 VSUBS 0.011509f
C641 B.n508 VSUBS 0.011509f
C642 B.n509 VSUBS 0.011509f
C643 B.n510 VSUBS 0.011509f
C644 B.n511 VSUBS 0.011509f
C645 B.n512 VSUBS 0.011509f
C646 B.n513 VSUBS 0.011509f
C647 B.n514 VSUBS 0.011509f
C648 B.n515 VSUBS 0.011509f
C649 B.n516 VSUBS 0.011509f
C650 B.n517 VSUBS 0.011509f
C651 B.n518 VSUBS 0.011509f
C652 B.n519 VSUBS 0.011509f
C653 B.n520 VSUBS 0.011509f
C654 B.n521 VSUBS 0.011509f
C655 B.n522 VSUBS 0.011509f
C656 B.n523 VSUBS 0.011509f
C657 B.n524 VSUBS 0.028503f
C658 B.n525 VSUBS 0.027014f
C659 B.n526 VSUBS 0.027014f
C660 B.n527 VSUBS 0.011509f
C661 B.n528 VSUBS 0.011509f
C662 B.n529 VSUBS 0.011509f
C663 B.n530 VSUBS 0.011509f
C664 B.n531 VSUBS 0.011509f
C665 B.n532 VSUBS 0.011509f
C666 B.n533 VSUBS 0.011509f
C667 B.n534 VSUBS 0.011509f
C668 B.n535 VSUBS 0.011509f
C669 B.n536 VSUBS 0.011509f
C670 B.n537 VSUBS 0.011509f
C671 B.n538 VSUBS 0.011509f
C672 B.n539 VSUBS 0.011509f
C673 B.n540 VSUBS 0.011509f
C674 B.n541 VSUBS 0.011509f
C675 B.n542 VSUBS 0.011509f
C676 B.n543 VSUBS 0.011509f
C677 B.n544 VSUBS 0.011509f
C678 B.n545 VSUBS 0.011509f
C679 B.n546 VSUBS 0.011509f
C680 B.n547 VSUBS 0.011509f
C681 B.n548 VSUBS 0.011509f
C682 B.n549 VSUBS 0.011509f
C683 B.n550 VSUBS 0.011509f
C684 B.n551 VSUBS 0.011509f
C685 B.n552 VSUBS 0.011509f
C686 B.n553 VSUBS 0.011509f
C687 B.n554 VSUBS 0.011509f
C688 B.n555 VSUBS 0.011509f
C689 B.n556 VSUBS 0.011509f
C690 B.n557 VSUBS 0.011509f
C691 B.n558 VSUBS 0.011509f
C692 B.n559 VSUBS 0.011509f
C693 B.n560 VSUBS 0.011509f
C694 B.n561 VSUBS 0.011509f
C695 B.n562 VSUBS 0.011509f
C696 B.n563 VSUBS 0.011509f
C697 B.n564 VSUBS 0.011509f
C698 B.n565 VSUBS 0.011509f
C699 B.n566 VSUBS 0.011509f
C700 B.n567 VSUBS 0.011509f
C701 B.n568 VSUBS 0.011509f
C702 B.n569 VSUBS 0.011509f
C703 B.n570 VSUBS 0.011509f
C704 B.n571 VSUBS 0.011509f
C705 B.n572 VSUBS 0.011509f
C706 B.n573 VSUBS 0.011509f
C707 B.n574 VSUBS 0.011509f
C708 B.n575 VSUBS 0.011509f
C709 B.n576 VSUBS 0.011509f
C710 B.n577 VSUBS 0.011509f
C711 B.n578 VSUBS 0.011509f
C712 B.n579 VSUBS 0.011509f
C713 B.n580 VSUBS 0.011509f
C714 B.n581 VSUBS 0.011509f
C715 B.n582 VSUBS 0.011509f
C716 B.n583 VSUBS 0.011509f
C717 B.n584 VSUBS 0.011509f
C718 B.n585 VSUBS 0.011509f
C719 B.n586 VSUBS 0.011509f
C720 B.n587 VSUBS 0.011509f
C721 B.n588 VSUBS 0.011509f
C722 B.n589 VSUBS 0.011509f
C723 B.n590 VSUBS 0.011509f
C724 B.n591 VSUBS 0.011509f
C725 B.n592 VSUBS 0.011509f
C726 B.n593 VSUBS 0.011509f
C727 B.n594 VSUBS 0.011509f
C728 B.n595 VSUBS 0.011509f
C729 B.n596 VSUBS 0.011509f
C730 B.n597 VSUBS 0.011509f
C731 B.n598 VSUBS 0.011509f
C732 B.n599 VSUBS 0.011509f
C733 B.n600 VSUBS 0.011509f
C734 B.n601 VSUBS 0.011509f
C735 B.n602 VSUBS 0.011509f
C736 B.n603 VSUBS 0.011509f
C737 B.n604 VSUBS 0.011509f
C738 B.n605 VSUBS 0.011509f
C739 B.n606 VSUBS 0.011509f
C740 B.n607 VSUBS 0.026061f
C741 VDD2.t0 VSUBS 0.058151f
C742 VDD2.t4 VSUBS 0.058151f
C743 VDD2.n0 VSUBS 0.299846f
C744 VDD2.t6 VSUBS 0.058151f
C745 VDD2.t5 VSUBS 0.058151f
C746 VDD2.n1 VSUBS 0.299846f
C747 VDD2.n2 VSUBS 3.01482f
C748 VDD2.t1 VSUBS 0.058151f
C749 VDD2.t7 VSUBS 0.058151f
C750 VDD2.n3 VSUBS 0.293847f
C751 VDD2.n4 VSUBS 2.37822f
C752 VDD2.t3 VSUBS 0.058151f
C753 VDD2.t2 VSUBS 0.058151f
C754 VDD2.n5 VSUBS 0.299828f
C755 VTAIL.t12 VSUBS 0.084401f
C756 VTAIL.t10 VSUBS 0.084401f
C757 VTAIL.n0 VSUBS 0.363074f
C758 VTAIL.n1 VSUBS 0.794876f
C759 VTAIL.t14 VSUBS 0.551774f
C760 VTAIL.n2 VSUBS 0.883113f
C761 VTAIL.t5 VSUBS 0.551774f
C762 VTAIL.n3 VSUBS 0.883113f
C763 VTAIL.t3 VSUBS 0.084401f
C764 VTAIL.t1 VSUBS 0.084401f
C765 VTAIL.n4 VSUBS 0.363074f
C766 VTAIL.n5 VSUBS 1.09474f
C767 VTAIL.t2 VSUBS 0.551774f
C768 VTAIL.n6 VSUBS 1.91172f
C769 VTAIL.t8 VSUBS 0.551776f
C770 VTAIL.n7 VSUBS 1.91172f
C771 VTAIL.t7 VSUBS 0.084401f
C772 VTAIL.t13 VSUBS 0.084401f
C773 VTAIL.n8 VSUBS 0.363076f
C774 VTAIL.n9 VSUBS 1.09474f
C775 VTAIL.t11 VSUBS 0.551776f
C776 VTAIL.n10 VSUBS 0.883111f
C777 VTAIL.t6 VSUBS 0.551776f
C778 VTAIL.n11 VSUBS 0.883111f
C779 VTAIL.t15 VSUBS 0.084401f
C780 VTAIL.t4 VSUBS 0.084401f
C781 VTAIL.n12 VSUBS 0.363076f
C782 VTAIL.n13 VSUBS 1.09474f
C783 VTAIL.t0 VSUBS 0.551776f
C784 VTAIL.n14 VSUBS 1.91172f
C785 VTAIL.t9 VSUBS 0.551774f
C786 VTAIL.n15 VSUBS 1.90511f
C787 VN.t2 VSUBS 0.964458f
C788 VN.n0 VSUBS 0.578029f
C789 VN.n1 VSUBS 0.045578f
C790 VN.n2 VSUBS 0.081826f
C791 VN.n3 VSUBS 0.045578f
C792 VN.t1 VSUBS 0.964458f
C793 VN.n4 VSUBS 0.084946f
C794 VN.n5 VSUBS 0.045578f
C795 VN.n6 VSUBS 0.069427f
C796 VN.t3 VSUBS 0.964458f
C797 VN.n7 VSUBS 0.54833f
C798 VN.t7 VSUBS 1.34882f
C799 VN.n8 VSUBS 0.529127f
C800 VN.n9 VSUBS 0.480889f
C801 VN.n10 VSUBS 0.045578f
C802 VN.n11 VSUBS 0.084946f
C803 VN.n12 VSUBS 0.066536f
C804 VN.n13 VSUBS 0.066536f
C805 VN.n14 VSUBS 0.045578f
C806 VN.n15 VSUBS 0.045578f
C807 VN.n16 VSUBS 0.045578f
C808 VN.n17 VSUBS 0.069427f
C809 VN.n18 VSUBS 0.403159f
C810 VN.n19 VSUBS 0.058523f
C811 VN.n20 VSUBS 0.084946f
C812 VN.n21 VSUBS 0.045578f
C813 VN.n22 VSUBS 0.045578f
C814 VN.n23 VSUBS 0.045578f
C815 VN.n24 VSUBS 0.046037f
C816 VN.n25 VSUBS 0.090156f
C817 VN.n26 VSUBS 0.080331f
C818 VN.n27 VSUBS 0.073562f
C819 VN.n28 VSUBS 0.088321f
C820 VN.t6 VSUBS 0.964458f
C821 VN.n29 VSUBS 0.578029f
C822 VN.n30 VSUBS 0.045578f
C823 VN.n31 VSUBS 0.081826f
C824 VN.n32 VSUBS 0.045578f
C825 VN.t0 VSUBS 0.964458f
C826 VN.n33 VSUBS 0.084946f
C827 VN.n34 VSUBS 0.045578f
C828 VN.n35 VSUBS 0.069427f
C829 VN.t5 VSUBS 1.34882f
C830 VN.t4 VSUBS 0.964458f
C831 VN.n36 VSUBS 0.54833f
C832 VN.n37 VSUBS 0.529127f
C833 VN.n38 VSUBS 0.480889f
C834 VN.n39 VSUBS 0.045578f
C835 VN.n40 VSUBS 0.084946f
C836 VN.n41 VSUBS 0.066536f
C837 VN.n42 VSUBS 0.066536f
C838 VN.n43 VSUBS 0.045578f
C839 VN.n44 VSUBS 0.045578f
C840 VN.n45 VSUBS 0.045578f
C841 VN.n46 VSUBS 0.069427f
C842 VN.n47 VSUBS 0.403159f
C843 VN.n48 VSUBS 0.058523f
C844 VN.n49 VSUBS 0.084946f
C845 VN.n50 VSUBS 0.045578f
C846 VN.n51 VSUBS 0.045578f
C847 VN.n52 VSUBS 0.045578f
C848 VN.n53 VSUBS 0.046037f
C849 VN.n54 VSUBS 0.090156f
C850 VN.n55 VSUBS 0.080331f
C851 VN.n56 VSUBS 0.073562f
C852 VN.n57 VSUBS 2.22447f
.ends

