* NGSPICE file created from diff_pair_sample_0257.ext - technology: sky130A

.subckt diff_pair_sample_0257 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.25
X1 VDD1.t5 VP.t0 VTAIL.t1 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.25
X2 B.t11 B.t9 B.t10 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.25
X3 B.t8 B.t6 B.t7 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.25
X4 B.t5 B.t3 B.t4 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.25
X5 VTAIL.t2 VP.t1 VDD1.t4 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.25
X6 VDD2.t4 VN.t1 VTAIL.t6 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.25
X7 B.t2 B.t0 B.t1 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=0 ps=0 w=15.81 l=2.25
X8 VDD1.t3 VP.t2 VTAIL.t0 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.25
X9 VTAIL.t3 VP.t3 VDD1.t2 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.25
X10 VTAIL.t7 VN.t2 VDD2.t3 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.25
X11 VDD1.t1 VP.t4 VTAIL.t10 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.25
X12 VTAIL.t4 VN.t3 VDD2.t2 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=2.60865 ps=16.14 w=15.81 l=2.25
X13 VDD1.t0 VP.t5 VTAIL.t11 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.25
X14 VDD2.t1 VN.t4 VTAIL.t9 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=6.1659 pd=32.4 as=2.60865 ps=16.14 w=15.81 l=2.25
X15 VDD2.t0 VN.t5 VTAIL.t5 w_n3034_n4130# sky130_fd_pr__pfet_01v8 ad=2.60865 pd=16.14 as=6.1659 ps=32.4 w=15.81 l=2.25
R0 VN.n3 VN.t4 202.423
R1 VN.n17 VN.t1 202.423
R2 VN.n4 VN.t2 169.344
R3 VN.n12 VN.t5 169.344
R4 VN.n18 VN.t3 169.344
R5 VN.n26 VN.t0 169.344
R6 VN.n25 VN.n14 161.3
R7 VN.n24 VN.n23 161.3
R8 VN.n22 VN.n15 161.3
R9 VN.n21 VN.n20 161.3
R10 VN.n19 VN.n16 161.3
R11 VN.n11 VN.n0 161.3
R12 VN.n10 VN.n9 161.3
R13 VN.n8 VN.n1 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n13 VN.n12 94.6082
R17 VN.n27 VN.n26 94.6082
R18 VN.n4 VN.n3 59.2533
R19 VN.n18 VN.n17 59.2533
R20 VN VN.n27 50.4982
R21 VN.n10 VN.n1 44.3785
R22 VN.n24 VN.n15 44.3785
R23 VN.n6 VN.n1 36.6083
R24 VN.n20 VN.n15 36.6083
R25 VN.n6 VN.n5 24.4675
R26 VN.n11 VN.n10 24.4675
R27 VN.n20 VN.n19 24.4675
R28 VN.n25 VN.n24 24.4675
R29 VN.n12 VN.n11 16.1487
R30 VN.n26 VN.n25 16.1487
R31 VN.n5 VN.n4 12.234
R32 VN.n19 VN.n18 12.234
R33 VN.n17 VN.n16 9.34402
R34 VN.n3 VN.n2 9.34402
R35 VN.n27 VN.n14 0.278367
R36 VN.n13 VN.n0 0.278367
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153454
R46 VTAIL.n7 VTAIL.t6 57.1463
R47 VTAIL.n11 VTAIL.t5 57.1462
R48 VTAIL.n2 VTAIL.t1 57.1462
R49 VTAIL.n10 VTAIL.t0 57.1462
R50 VTAIL.n9 VTAIL.n8 55.0904
R51 VTAIL.n6 VTAIL.n5 55.0904
R52 VTAIL.n1 VTAIL.n0 55.0902
R53 VTAIL.n4 VTAIL.n3 55.0902
R54 VTAIL.n6 VTAIL.n4 30.4445
R55 VTAIL.n11 VTAIL.n10 28.2203
R56 VTAIL.n7 VTAIL.n6 2.22464
R57 VTAIL.n10 VTAIL.n9 2.22464
R58 VTAIL.n4 VTAIL.n2 2.22464
R59 VTAIL.n0 VTAIL.t9 2.05648
R60 VTAIL.n0 VTAIL.t7 2.05648
R61 VTAIL.n3 VTAIL.t10 2.05648
R62 VTAIL.n3 VTAIL.t3 2.05648
R63 VTAIL.n8 VTAIL.t11 2.05648
R64 VTAIL.n8 VTAIL.t2 2.05648
R65 VTAIL.n5 VTAIL.t8 2.05648
R66 VTAIL.n5 VTAIL.t4 2.05648
R67 VTAIL VTAIL.n11 1.61041
R68 VTAIL.n9 VTAIL.n7 1.5824
R69 VTAIL.n2 VTAIL.n1 1.5824
R70 VTAIL VTAIL.n1 0.614724
R71 VDD2.n1 VDD2.t1 75.4378
R72 VDD2.n2 VDD2.t5 73.8251
R73 VDD2.n1 VDD2.n0 72.2697
R74 VDD2 VDD2.n3 72.2669
R75 VDD2.n2 VDD2.n1 44.5731
R76 VDD2.n3 VDD2.t2 2.05648
R77 VDD2.n3 VDD2.t4 2.05648
R78 VDD2.n0 VDD2.t3 2.05648
R79 VDD2.n0 VDD2.t0 2.05648
R80 VDD2 VDD2.n2 1.72679
R81 VP.n9 VP.t5 202.423
R82 VP.n5 VP.t4 169.344
R83 VP.n29 VP.t3 169.344
R84 VP.n37 VP.t0 169.344
R85 VP.n18 VP.t2 169.344
R86 VP.n10 VP.t1 169.344
R87 VP.n11 VP.n8 161.3
R88 VP.n13 VP.n12 161.3
R89 VP.n14 VP.n7 161.3
R90 VP.n16 VP.n15 161.3
R91 VP.n17 VP.n6 161.3
R92 VP.n36 VP.n0 161.3
R93 VP.n35 VP.n34 161.3
R94 VP.n33 VP.n1 161.3
R95 VP.n32 VP.n31 161.3
R96 VP.n30 VP.n2 161.3
R97 VP.n28 VP.n27 161.3
R98 VP.n26 VP.n3 161.3
R99 VP.n25 VP.n24 161.3
R100 VP.n23 VP.n4 161.3
R101 VP.n22 VP.n21 161.3
R102 VP.n20 VP.n5 94.6082
R103 VP.n38 VP.n37 94.6082
R104 VP.n19 VP.n18 94.6082
R105 VP.n10 VP.n9 59.2533
R106 VP.n20 VP.n19 50.2193
R107 VP.n24 VP.n23 44.3785
R108 VP.n35 VP.n1 44.3785
R109 VP.n16 VP.n7 44.3785
R110 VP.n24 VP.n3 36.6083
R111 VP.n31 VP.n1 36.6083
R112 VP.n12 VP.n7 36.6083
R113 VP.n23 VP.n22 24.4675
R114 VP.n28 VP.n3 24.4675
R115 VP.n31 VP.n30 24.4675
R116 VP.n36 VP.n35 24.4675
R117 VP.n17 VP.n16 24.4675
R118 VP.n12 VP.n11 24.4675
R119 VP.n22 VP.n5 16.1487
R120 VP.n37 VP.n36 16.1487
R121 VP.n18 VP.n17 16.1487
R122 VP.n29 VP.n28 12.234
R123 VP.n30 VP.n29 12.234
R124 VP.n11 VP.n10 12.234
R125 VP.n9 VP.n8 9.34402
R126 VP.n19 VP.n6 0.278367
R127 VP.n21 VP.n20 0.278367
R128 VP.n38 VP.n0 0.278367
R129 VP.n13 VP.n8 0.189894
R130 VP.n14 VP.n13 0.189894
R131 VP.n15 VP.n14 0.189894
R132 VP.n15 VP.n6 0.189894
R133 VP.n21 VP.n4 0.189894
R134 VP.n25 VP.n4 0.189894
R135 VP.n26 VP.n25 0.189894
R136 VP.n27 VP.n26 0.189894
R137 VP.n27 VP.n2 0.189894
R138 VP.n32 VP.n2 0.189894
R139 VP.n33 VP.n32 0.189894
R140 VP.n34 VP.n33 0.189894
R141 VP.n34 VP.n0 0.189894
R142 VP VP.n38 0.153454
R143 VDD1 VDD1.t0 75.5514
R144 VDD1.n1 VDD1.t1 75.4378
R145 VDD1.n1 VDD1.n0 72.2697
R146 VDD1.n3 VDD1.n2 71.769
R147 VDD1.n3 VDD1.n1 46.2681
R148 VDD1.n2 VDD1.t4 2.05648
R149 VDD1.n2 VDD1.t3 2.05648
R150 VDD1.n0 VDD1.t2 2.05648
R151 VDD1.n0 VDD1.t5 2.05648
R152 VDD1 VDD1.n3 0.498345
R153 B.n431 B.n122 585
R154 B.n430 B.n429 585
R155 B.n428 B.n123 585
R156 B.n427 B.n426 585
R157 B.n425 B.n124 585
R158 B.n424 B.n423 585
R159 B.n422 B.n125 585
R160 B.n421 B.n420 585
R161 B.n419 B.n126 585
R162 B.n418 B.n417 585
R163 B.n416 B.n127 585
R164 B.n415 B.n414 585
R165 B.n413 B.n128 585
R166 B.n412 B.n411 585
R167 B.n410 B.n129 585
R168 B.n409 B.n408 585
R169 B.n407 B.n130 585
R170 B.n406 B.n405 585
R171 B.n404 B.n131 585
R172 B.n403 B.n402 585
R173 B.n401 B.n132 585
R174 B.n400 B.n399 585
R175 B.n398 B.n133 585
R176 B.n397 B.n396 585
R177 B.n395 B.n134 585
R178 B.n394 B.n393 585
R179 B.n392 B.n135 585
R180 B.n391 B.n390 585
R181 B.n389 B.n136 585
R182 B.n388 B.n387 585
R183 B.n386 B.n137 585
R184 B.n385 B.n384 585
R185 B.n383 B.n138 585
R186 B.n382 B.n381 585
R187 B.n380 B.n139 585
R188 B.n379 B.n378 585
R189 B.n377 B.n140 585
R190 B.n376 B.n375 585
R191 B.n374 B.n141 585
R192 B.n373 B.n372 585
R193 B.n371 B.n142 585
R194 B.n370 B.n369 585
R195 B.n368 B.n143 585
R196 B.n367 B.n366 585
R197 B.n365 B.n144 585
R198 B.n364 B.n363 585
R199 B.n362 B.n145 585
R200 B.n361 B.n360 585
R201 B.n359 B.n146 585
R202 B.n358 B.n357 585
R203 B.n356 B.n147 585
R204 B.n355 B.n354 585
R205 B.n353 B.n148 585
R206 B.n352 B.n351 585
R207 B.n347 B.n149 585
R208 B.n346 B.n345 585
R209 B.n344 B.n150 585
R210 B.n343 B.n342 585
R211 B.n341 B.n151 585
R212 B.n340 B.n339 585
R213 B.n338 B.n152 585
R214 B.n337 B.n336 585
R215 B.n334 B.n153 585
R216 B.n333 B.n332 585
R217 B.n331 B.n156 585
R218 B.n330 B.n329 585
R219 B.n328 B.n157 585
R220 B.n327 B.n326 585
R221 B.n325 B.n158 585
R222 B.n324 B.n323 585
R223 B.n322 B.n159 585
R224 B.n321 B.n320 585
R225 B.n319 B.n160 585
R226 B.n318 B.n317 585
R227 B.n316 B.n161 585
R228 B.n315 B.n314 585
R229 B.n313 B.n162 585
R230 B.n312 B.n311 585
R231 B.n310 B.n163 585
R232 B.n309 B.n308 585
R233 B.n307 B.n164 585
R234 B.n306 B.n305 585
R235 B.n304 B.n165 585
R236 B.n303 B.n302 585
R237 B.n301 B.n166 585
R238 B.n300 B.n299 585
R239 B.n298 B.n167 585
R240 B.n297 B.n296 585
R241 B.n295 B.n168 585
R242 B.n294 B.n293 585
R243 B.n292 B.n169 585
R244 B.n291 B.n290 585
R245 B.n289 B.n170 585
R246 B.n288 B.n287 585
R247 B.n286 B.n171 585
R248 B.n285 B.n284 585
R249 B.n283 B.n172 585
R250 B.n282 B.n281 585
R251 B.n280 B.n173 585
R252 B.n279 B.n278 585
R253 B.n277 B.n174 585
R254 B.n276 B.n275 585
R255 B.n274 B.n175 585
R256 B.n273 B.n272 585
R257 B.n271 B.n176 585
R258 B.n270 B.n269 585
R259 B.n268 B.n177 585
R260 B.n267 B.n266 585
R261 B.n265 B.n178 585
R262 B.n264 B.n263 585
R263 B.n262 B.n179 585
R264 B.n261 B.n260 585
R265 B.n259 B.n180 585
R266 B.n258 B.n257 585
R267 B.n256 B.n181 585
R268 B.n433 B.n432 585
R269 B.n434 B.n121 585
R270 B.n436 B.n435 585
R271 B.n437 B.n120 585
R272 B.n439 B.n438 585
R273 B.n440 B.n119 585
R274 B.n442 B.n441 585
R275 B.n443 B.n118 585
R276 B.n445 B.n444 585
R277 B.n446 B.n117 585
R278 B.n448 B.n447 585
R279 B.n449 B.n116 585
R280 B.n451 B.n450 585
R281 B.n452 B.n115 585
R282 B.n454 B.n453 585
R283 B.n455 B.n114 585
R284 B.n457 B.n456 585
R285 B.n458 B.n113 585
R286 B.n460 B.n459 585
R287 B.n461 B.n112 585
R288 B.n463 B.n462 585
R289 B.n464 B.n111 585
R290 B.n466 B.n465 585
R291 B.n467 B.n110 585
R292 B.n469 B.n468 585
R293 B.n470 B.n109 585
R294 B.n472 B.n471 585
R295 B.n473 B.n108 585
R296 B.n475 B.n474 585
R297 B.n476 B.n107 585
R298 B.n478 B.n477 585
R299 B.n479 B.n106 585
R300 B.n481 B.n480 585
R301 B.n482 B.n105 585
R302 B.n484 B.n483 585
R303 B.n485 B.n104 585
R304 B.n487 B.n486 585
R305 B.n488 B.n103 585
R306 B.n490 B.n489 585
R307 B.n491 B.n102 585
R308 B.n493 B.n492 585
R309 B.n494 B.n101 585
R310 B.n496 B.n495 585
R311 B.n497 B.n100 585
R312 B.n499 B.n498 585
R313 B.n500 B.n99 585
R314 B.n502 B.n501 585
R315 B.n503 B.n98 585
R316 B.n505 B.n504 585
R317 B.n506 B.n97 585
R318 B.n508 B.n507 585
R319 B.n509 B.n96 585
R320 B.n511 B.n510 585
R321 B.n512 B.n95 585
R322 B.n514 B.n513 585
R323 B.n515 B.n94 585
R324 B.n517 B.n516 585
R325 B.n518 B.n93 585
R326 B.n520 B.n519 585
R327 B.n521 B.n92 585
R328 B.n523 B.n522 585
R329 B.n524 B.n91 585
R330 B.n526 B.n525 585
R331 B.n527 B.n90 585
R332 B.n529 B.n528 585
R333 B.n530 B.n89 585
R334 B.n532 B.n531 585
R335 B.n533 B.n88 585
R336 B.n535 B.n534 585
R337 B.n536 B.n87 585
R338 B.n538 B.n537 585
R339 B.n539 B.n86 585
R340 B.n541 B.n540 585
R341 B.n542 B.n85 585
R342 B.n544 B.n543 585
R343 B.n545 B.n84 585
R344 B.n547 B.n546 585
R345 B.n548 B.n83 585
R346 B.n722 B.n21 585
R347 B.n721 B.n720 585
R348 B.n719 B.n22 585
R349 B.n718 B.n717 585
R350 B.n716 B.n23 585
R351 B.n715 B.n714 585
R352 B.n713 B.n24 585
R353 B.n712 B.n711 585
R354 B.n710 B.n25 585
R355 B.n709 B.n708 585
R356 B.n707 B.n26 585
R357 B.n706 B.n705 585
R358 B.n704 B.n27 585
R359 B.n703 B.n702 585
R360 B.n701 B.n28 585
R361 B.n700 B.n699 585
R362 B.n698 B.n29 585
R363 B.n697 B.n696 585
R364 B.n695 B.n30 585
R365 B.n694 B.n693 585
R366 B.n692 B.n31 585
R367 B.n691 B.n690 585
R368 B.n689 B.n32 585
R369 B.n688 B.n687 585
R370 B.n686 B.n33 585
R371 B.n685 B.n684 585
R372 B.n683 B.n34 585
R373 B.n682 B.n681 585
R374 B.n680 B.n35 585
R375 B.n679 B.n678 585
R376 B.n677 B.n36 585
R377 B.n676 B.n675 585
R378 B.n674 B.n37 585
R379 B.n673 B.n672 585
R380 B.n671 B.n38 585
R381 B.n670 B.n669 585
R382 B.n668 B.n39 585
R383 B.n667 B.n666 585
R384 B.n665 B.n40 585
R385 B.n664 B.n663 585
R386 B.n662 B.n41 585
R387 B.n661 B.n660 585
R388 B.n659 B.n42 585
R389 B.n658 B.n657 585
R390 B.n656 B.n43 585
R391 B.n655 B.n654 585
R392 B.n653 B.n44 585
R393 B.n652 B.n651 585
R394 B.n650 B.n45 585
R395 B.n649 B.n648 585
R396 B.n647 B.n46 585
R397 B.n646 B.n645 585
R398 B.n644 B.n47 585
R399 B.n642 B.n641 585
R400 B.n640 B.n50 585
R401 B.n639 B.n638 585
R402 B.n637 B.n51 585
R403 B.n636 B.n635 585
R404 B.n634 B.n52 585
R405 B.n633 B.n632 585
R406 B.n631 B.n53 585
R407 B.n630 B.n629 585
R408 B.n628 B.n627 585
R409 B.n626 B.n57 585
R410 B.n625 B.n624 585
R411 B.n623 B.n58 585
R412 B.n622 B.n621 585
R413 B.n620 B.n59 585
R414 B.n619 B.n618 585
R415 B.n617 B.n60 585
R416 B.n616 B.n615 585
R417 B.n614 B.n61 585
R418 B.n613 B.n612 585
R419 B.n611 B.n62 585
R420 B.n610 B.n609 585
R421 B.n608 B.n63 585
R422 B.n607 B.n606 585
R423 B.n605 B.n64 585
R424 B.n604 B.n603 585
R425 B.n602 B.n65 585
R426 B.n601 B.n600 585
R427 B.n599 B.n66 585
R428 B.n598 B.n597 585
R429 B.n596 B.n67 585
R430 B.n595 B.n594 585
R431 B.n593 B.n68 585
R432 B.n592 B.n591 585
R433 B.n590 B.n69 585
R434 B.n589 B.n588 585
R435 B.n587 B.n70 585
R436 B.n586 B.n585 585
R437 B.n584 B.n71 585
R438 B.n583 B.n582 585
R439 B.n581 B.n72 585
R440 B.n580 B.n579 585
R441 B.n578 B.n73 585
R442 B.n577 B.n576 585
R443 B.n575 B.n74 585
R444 B.n574 B.n573 585
R445 B.n572 B.n75 585
R446 B.n571 B.n570 585
R447 B.n569 B.n76 585
R448 B.n568 B.n567 585
R449 B.n566 B.n77 585
R450 B.n565 B.n564 585
R451 B.n563 B.n78 585
R452 B.n562 B.n561 585
R453 B.n560 B.n79 585
R454 B.n559 B.n558 585
R455 B.n557 B.n80 585
R456 B.n556 B.n555 585
R457 B.n554 B.n81 585
R458 B.n553 B.n552 585
R459 B.n551 B.n82 585
R460 B.n550 B.n549 585
R461 B.n724 B.n723 585
R462 B.n725 B.n20 585
R463 B.n727 B.n726 585
R464 B.n728 B.n19 585
R465 B.n730 B.n729 585
R466 B.n731 B.n18 585
R467 B.n733 B.n732 585
R468 B.n734 B.n17 585
R469 B.n736 B.n735 585
R470 B.n737 B.n16 585
R471 B.n739 B.n738 585
R472 B.n740 B.n15 585
R473 B.n742 B.n741 585
R474 B.n743 B.n14 585
R475 B.n745 B.n744 585
R476 B.n746 B.n13 585
R477 B.n748 B.n747 585
R478 B.n749 B.n12 585
R479 B.n751 B.n750 585
R480 B.n752 B.n11 585
R481 B.n754 B.n753 585
R482 B.n755 B.n10 585
R483 B.n757 B.n756 585
R484 B.n758 B.n9 585
R485 B.n760 B.n759 585
R486 B.n761 B.n8 585
R487 B.n763 B.n762 585
R488 B.n764 B.n7 585
R489 B.n766 B.n765 585
R490 B.n767 B.n6 585
R491 B.n769 B.n768 585
R492 B.n770 B.n5 585
R493 B.n772 B.n771 585
R494 B.n773 B.n4 585
R495 B.n775 B.n774 585
R496 B.n776 B.n3 585
R497 B.n778 B.n777 585
R498 B.n779 B.n0 585
R499 B.n2 B.n1 585
R500 B.n201 B.n200 585
R501 B.n202 B.n199 585
R502 B.n204 B.n203 585
R503 B.n205 B.n198 585
R504 B.n207 B.n206 585
R505 B.n208 B.n197 585
R506 B.n210 B.n209 585
R507 B.n211 B.n196 585
R508 B.n213 B.n212 585
R509 B.n214 B.n195 585
R510 B.n216 B.n215 585
R511 B.n217 B.n194 585
R512 B.n219 B.n218 585
R513 B.n220 B.n193 585
R514 B.n222 B.n221 585
R515 B.n223 B.n192 585
R516 B.n225 B.n224 585
R517 B.n226 B.n191 585
R518 B.n228 B.n227 585
R519 B.n229 B.n190 585
R520 B.n231 B.n230 585
R521 B.n232 B.n189 585
R522 B.n234 B.n233 585
R523 B.n235 B.n188 585
R524 B.n237 B.n236 585
R525 B.n238 B.n187 585
R526 B.n240 B.n239 585
R527 B.n241 B.n186 585
R528 B.n243 B.n242 585
R529 B.n244 B.n185 585
R530 B.n246 B.n245 585
R531 B.n247 B.n184 585
R532 B.n249 B.n248 585
R533 B.n250 B.n183 585
R534 B.n252 B.n251 585
R535 B.n253 B.n182 585
R536 B.n255 B.n254 585
R537 B.n254 B.n181 511.721
R538 B.n432 B.n431 511.721
R539 B.n550 B.n83 511.721
R540 B.n724 B.n21 511.721
R541 B.n348 B.t3 377.45
R542 B.n54 B.t0 377.45
R543 B.n154 B.t9 377.087
R544 B.n48 B.t6 377.087
R545 B.n781 B.n780 256.663
R546 B.n780 B.n779 235.042
R547 B.n780 B.n2 235.042
R548 B.n258 B.n181 163.367
R549 B.n259 B.n258 163.367
R550 B.n260 B.n259 163.367
R551 B.n260 B.n179 163.367
R552 B.n264 B.n179 163.367
R553 B.n265 B.n264 163.367
R554 B.n266 B.n265 163.367
R555 B.n266 B.n177 163.367
R556 B.n270 B.n177 163.367
R557 B.n271 B.n270 163.367
R558 B.n272 B.n271 163.367
R559 B.n272 B.n175 163.367
R560 B.n276 B.n175 163.367
R561 B.n277 B.n276 163.367
R562 B.n278 B.n277 163.367
R563 B.n278 B.n173 163.367
R564 B.n282 B.n173 163.367
R565 B.n283 B.n282 163.367
R566 B.n284 B.n283 163.367
R567 B.n284 B.n171 163.367
R568 B.n288 B.n171 163.367
R569 B.n289 B.n288 163.367
R570 B.n290 B.n289 163.367
R571 B.n290 B.n169 163.367
R572 B.n294 B.n169 163.367
R573 B.n295 B.n294 163.367
R574 B.n296 B.n295 163.367
R575 B.n296 B.n167 163.367
R576 B.n300 B.n167 163.367
R577 B.n301 B.n300 163.367
R578 B.n302 B.n301 163.367
R579 B.n302 B.n165 163.367
R580 B.n306 B.n165 163.367
R581 B.n307 B.n306 163.367
R582 B.n308 B.n307 163.367
R583 B.n308 B.n163 163.367
R584 B.n312 B.n163 163.367
R585 B.n313 B.n312 163.367
R586 B.n314 B.n313 163.367
R587 B.n314 B.n161 163.367
R588 B.n318 B.n161 163.367
R589 B.n319 B.n318 163.367
R590 B.n320 B.n319 163.367
R591 B.n320 B.n159 163.367
R592 B.n324 B.n159 163.367
R593 B.n325 B.n324 163.367
R594 B.n326 B.n325 163.367
R595 B.n326 B.n157 163.367
R596 B.n330 B.n157 163.367
R597 B.n331 B.n330 163.367
R598 B.n332 B.n331 163.367
R599 B.n332 B.n153 163.367
R600 B.n337 B.n153 163.367
R601 B.n338 B.n337 163.367
R602 B.n339 B.n338 163.367
R603 B.n339 B.n151 163.367
R604 B.n343 B.n151 163.367
R605 B.n344 B.n343 163.367
R606 B.n345 B.n344 163.367
R607 B.n345 B.n149 163.367
R608 B.n352 B.n149 163.367
R609 B.n353 B.n352 163.367
R610 B.n354 B.n353 163.367
R611 B.n354 B.n147 163.367
R612 B.n358 B.n147 163.367
R613 B.n359 B.n358 163.367
R614 B.n360 B.n359 163.367
R615 B.n360 B.n145 163.367
R616 B.n364 B.n145 163.367
R617 B.n365 B.n364 163.367
R618 B.n366 B.n365 163.367
R619 B.n366 B.n143 163.367
R620 B.n370 B.n143 163.367
R621 B.n371 B.n370 163.367
R622 B.n372 B.n371 163.367
R623 B.n372 B.n141 163.367
R624 B.n376 B.n141 163.367
R625 B.n377 B.n376 163.367
R626 B.n378 B.n377 163.367
R627 B.n378 B.n139 163.367
R628 B.n382 B.n139 163.367
R629 B.n383 B.n382 163.367
R630 B.n384 B.n383 163.367
R631 B.n384 B.n137 163.367
R632 B.n388 B.n137 163.367
R633 B.n389 B.n388 163.367
R634 B.n390 B.n389 163.367
R635 B.n390 B.n135 163.367
R636 B.n394 B.n135 163.367
R637 B.n395 B.n394 163.367
R638 B.n396 B.n395 163.367
R639 B.n396 B.n133 163.367
R640 B.n400 B.n133 163.367
R641 B.n401 B.n400 163.367
R642 B.n402 B.n401 163.367
R643 B.n402 B.n131 163.367
R644 B.n406 B.n131 163.367
R645 B.n407 B.n406 163.367
R646 B.n408 B.n407 163.367
R647 B.n408 B.n129 163.367
R648 B.n412 B.n129 163.367
R649 B.n413 B.n412 163.367
R650 B.n414 B.n413 163.367
R651 B.n414 B.n127 163.367
R652 B.n418 B.n127 163.367
R653 B.n419 B.n418 163.367
R654 B.n420 B.n419 163.367
R655 B.n420 B.n125 163.367
R656 B.n424 B.n125 163.367
R657 B.n425 B.n424 163.367
R658 B.n426 B.n425 163.367
R659 B.n426 B.n123 163.367
R660 B.n430 B.n123 163.367
R661 B.n431 B.n430 163.367
R662 B.n546 B.n83 163.367
R663 B.n546 B.n545 163.367
R664 B.n545 B.n544 163.367
R665 B.n544 B.n85 163.367
R666 B.n540 B.n85 163.367
R667 B.n540 B.n539 163.367
R668 B.n539 B.n538 163.367
R669 B.n538 B.n87 163.367
R670 B.n534 B.n87 163.367
R671 B.n534 B.n533 163.367
R672 B.n533 B.n532 163.367
R673 B.n532 B.n89 163.367
R674 B.n528 B.n89 163.367
R675 B.n528 B.n527 163.367
R676 B.n527 B.n526 163.367
R677 B.n526 B.n91 163.367
R678 B.n522 B.n91 163.367
R679 B.n522 B.n521 163.367
R680 B.n521 B.n520 163.367
R681 B.n520 B.n93 163.367
R682 B.n516 B.n93 163.367
R683 B.n516 B.n515 163.367
R684 B.n515 B.n514 163.367
R685 B.n514 B.n95 163.367
R686 B.n510 B.n95 163.367
R687 B.n510 B.n509 163.367
R688 B.n509 B.n508 163.367
R689 B.n508 B.n97 163.367
R690 B.n504 B.n97 163.367
R691 B.n504 B.n503 163.367
R692 B.n503 B.n502 163.367
R693 B.n502 B.n99 163.367
R694 B.n498 B.n99 163.367
R695 B.n498 B.n497 163.367
R696 B.n497 B.n496 163.367
R697 B.n496 B.n101 163.367
R698 B.n492 B.n101 163.367
R699 B.n492 B.n491 163.367
R700 B.n491 B.n490 163.367
R701 B.n490 B.n103 163.367
R702 B.n486 B.n103 163.367
R703 B.n486 B.n485 163.367
R704 B.n485 B.n484 163.367
R705 B.n484 B.n105 163.367
R706 B.n480 B.n105 163.367
R707 B.n480 B.n479 163.367
R708 B.n479 B.n478 163.367
R709 B.n478 B.n107 163.367
R710 B.n474 B.n107 163.367
R711 B.n474 B.n473 163.367
R712 B.n473 B.n472 163.367
R713 B.n472 B.n109 163.367
R714 B.n468 B.n109 163.367
R715 B.n468 B.n467 163.367
R716 B.n467 B.n466 163.367
R717 B.n466 B.n111 163.367
R718 B.n462 B.n111 163.367
R719 B.n462 B.n461 163.367
R720 B.n461 B.n460 163.367
R721 B.n460 B.n113 163.367
R722 B.n456 B.n113 163.367
R723 B.n456 B.n455 163.367
R724 B.n455 B.n454 163.367
R725 B.n454 B.n115 163.367
R726 B.n450 B.n115 163.367
R727 B.n450 B.n449 163.367
R728 B.n449 B.n448 163.367
R729 B.n448 B.n117 163.367
R730 B.n444 B.n117 163.367
R731 B.n444 B.n443 163.367
R732 B.n443 B.n442 163.367
R733 B.n442 B.n119 163.367
R734 B.n438 B.n119 163.367
R735 B.n438 B.n437 163.367
R736 B.n437 B.n436 163.367
R737 B.n436 B.n121 163.367
R738 B.n432 B.n121 163.367
R739 B.n720 B.n21 163.367
R740 B.n720 B.n719 163.367
R741 B.n719 B.n718 163.367
R742 B.n718 B.n23 163.367
R743 B.n714 B.n23 163.367
R744 B.n714 B.n713 163.367
R745 B.n713 B.n712 163.367
R746 B.n712 B.n25 163.367
R747 B.n708 B.n25 163.367
R748 B.n708 B.n707 163.367
R749 B.n707 B.n706 163.367
R750 B.n706 B.n27 163.367
R751 B.n702 B.n27 163.367
R752 B.n702 B.n701 163.367
R753 B.n701 B.n700 163.367
R754 B.n700 B.n29 163.367
R755 B.n696 B.n29 163.367
R756 B.n696 B.n695 163.367
R757 B.n695 B.n694 163.367
R758 B.n694 B.n31 163.367
R759 B.n690 B.n31 163.367
R760 B.n690 B.n689 163.367
R761 B.n689 B.n688 163.367
R762 B.n688 B.n33 163.367
R763 B.n684 B.n33 163.367
R764 B.n684 B.n683 163.367
R765 B.n683 B.n682 163.367
R766 B.n682 B.n35 163.367
R767 B.n678 B.n35 163.367
R768 B.n678 B.n677 163.367
R769 B.n677 B.n676 163.367
R770 B.n676 B.n37 163.367
R771 B.n672 B.n37 163.367
R772 B.n672 B.n671 163.367
R773 B.n671 B.n670 163.367
R774 B.n670 B.n39 163.367
R775 B.n666 B.n39 163.367
R776 B.n666 B.n665 163.367
R777 B.n665 B.n664 163.367
R778 B.n664 B.n41 163.367
R779 B.n660 B.n41 163.367
R780 B.n660 B.n659 163.367
R781 B.n659 B.n658 163.367
R782 B.n658 B.n43 163.367
R783 B.n654 B.n43 163.367
R784 B.n654 B.n653 163.367
R785 B.n653 B.n652 163.367
R786 B.n652 B.n45 163.367
R787 B.n648 B.n45 163.367
R788 B.n648 B.n647 163.367
R789 B.n647 B.n646 163.367
R790 B.n646 B.n47 163.367
R791 B.n641 B.n47 163.367
R792 B.n641 B.n640 163.367
R793 B.n640 B.n639 163.367
R794 B.n639 B.n51 163.367
R795 B.n635 B.n51 163.367
R796 B.n635 B.n634 163.367
R797 B.n634 B.n633 163.367
R798 B.n633 B.n53 163.367
R799 B.n629 B.n53 163.367
R800 B.n629 B.n628 163.367
R801 B.n628 B.n57 163.367
R802 B.n624 B.n57 163.367
R803 B.n624 B.n623 163.367
R804 B.n623 B.n622 163.367
R805 B.n622 B.n59 163.367
R806 B.n618 B.n59 163.367
R807 B.n618 B.n617 163.367
R808 B.n617 B.n616 163.367
R809 B.n616 B.n61 163.367
R810 B.n612 B.n61 163.367
R811 B.n612 B.n611 163.367
R812 B.n611 B.n610 163.367
R813 B.n610 B.n63 163.367
R814 B.n606 B.n63 163.367
R815 B.n606 B.n605 163.367
R816 B.n605 B.n604 163.367
R817 B.n604 B.n65 163.367
R818 B.n600 B.n65 163.367
R819 B.n600 B.n599 163.367
R820 B.n599 B.n598 163.367
R821 B.n598 B.n67 163.367
R822 B.n594 B.n67 163.367
R823 B.n594 B.n593 163.367
R824 B.n593 B.n592 163.367
R825 B.n592 B.n69 163.367
R826 B.n588 B.n69 163.367
R827 B.n588 B.n587 163.367
R828 B.n587 B.n586 163.367
R829 B.n586 B.n71 163.367
R830 B.n582 B.n71 163.367
R831 B.n582 B.n581 163.367
R832 B.n581 B.n580 163.367
R833 B.n580 B.n73 163.367
R834 B.n576 B.n73 163.367
R835 B.n576 B.n575 163.367
R836 B.n575 B.n574 163.367
R837 B.n574 B.n75 163.367
R838 B.n570 B.n75 163.367
R839 B.n570 B.n569 163.367
R840 B.n569 B.n568 163.367
R841 B.n568 B.n77 163.367
R842 B.n564 B.n77 163.367
R843 B.n564 B.n563 163.367
R844 B.n563 B.n562 163.367
R845 B.n562 B.n79 163.367
R846 B.n558 B.n79 163.367
R847 B.n558 B.n557 163.367
R848 B.n557 B.n556 163.367
R849 B.n556 B.n81 163.367
R850 B.n552 B.n81 163.367
R851 B.n552 B.n551 163.367
R852 B.n551 B.n550 163.367
R853 B.n725 B.n724 163.367
R854 B.n726 B.n725 163.367
R855 B.n726 B.n19 163.367
R856 B.n730 B.n19 163.367
R857 B.n731 B.n730 163.367
R858 B.n732 B.n731 163.367
R859 B.n732 B.n17 163.367
R860 B.n736 B.n17 163.367
R861 B.n737 B.n736 163.367
R862 B.n738 B.n737 163.367
R863 B.n738 B.n15 163.367
R864 B.n742 B.n15 163.367
R865 B.n743 B.n742 163.367
R866 B.n744 B.n743 163.367
R867 B.n744 B.n13 163.367
R868 B.n748 B.n13 163.367
R869 B.n749 B.n748 163.367
R870 B.n750 B.n749 163.367
R871 B.n750 B.n11 163.367
R872 B.n754 B.n11 163.367
R873 B.n755 B.n754 163.367
R874 B.n756 B.n755 163.367
R875 B.n756 B.n9 163.367
R876 B.n760 B.n9 163.367
R877 B.n761 B.n760 163.367
R878 B.n762 B.n761 163.367
R879 B.n762 B.n7 163.367
R880 B.n766 B.n7 163.367
R881 B.n767 B.n766 163.367
R882 B.n768 B.n767 163.367
R883 B.n768 B.n5 163.367
R884 B.n772 B.n5 163.367
R885 B.n773 B.n772 163.367
R886 B.n774 B.n773 163.367
R887 B.n774 B.n3 163.367
R888 B.n778 B.n3 163.367
R889 B.n779 B.n778 163.367
R890 B.n200 B.n2 163.367
R891 B.n200 B.n199 163.367
R892 B.n204 B.n199 163.367
R893 B.n205 B.n204 163.367
R894 B.n206 B.n205 163.367
R895 B.n206 B.n197 163.367
R896 B.n210 B.n197 163.367
R897 B.n211 B.n210 163.367
R898 B.n212 B.n211 163.367
R899 B.n212 B.n195 163.367
R900 B.n216 B.n195 163.367
R901 B.n217 B.n216 163.367
R902 B.n218 B.n217 163.367
R903 B.n218 B.n193 163.367
R904 B.n222 B.n193 163.367
R905 B.n223 B.n222 163.367
R906 B.n224 B.n223 163.367
R907 B.n224 B.n191 163.367
R908 B.n228 B.n191 163.367
R909 B.n229 B.n228 163.367
R910 B.n230 B.n229 163.367
R911 B.n230 B.n189 163.367
R912 B.n234 B.n189 163.367
R913 B.n235 B.n234 163.367
R914 B.n236 B.n235 163.367
R915 B.n236 B.n187 163.367
R916 B.n240 B.n187 163.367
R917 B.n241 B.n240 163.367
R918 B.n242 B.n241 163.367
R919 B.n242 B.n185 163.367
R920 B.n246 B.n185 163.367
R921 B.n247 B.n246 163.367
R922 B.n248 B.n247 163.367
R923 B.n248 B.n183 163.367
R924 B.n252 B.n183 163.367
R925 B.n253 B.n252 163.367
R926 B.n254 B.n253 163.367
R927 B.n348 B.t4 159.978
R928 B.n54 B.t2 159.978
R929 B.n154 B.t10 159.958
R930 B.n48 B.t8 159.958
R931 B.n349 B.t5 109.942
R932 B.n55 B.t1 109.942
R933 B.n155 B.t11 109.922
R934 B.n49 B.t7 109.922
R935 B.n335 B.n155 59.5399
R936 B.n350 B.n349 59.5399
R937 B.n56 B.n55 59.5399
R938 B.n643 B.n49 59.5399
R939 B.n155 B.n154 50.0369
R940 B.n349 B.n348 50.0369
R941 B.n55 B.n54 50.0369
R942 B.n49 B.n48 50.0369
R943 B.n723 B.n722 33.2493
R944 B.n549 B.n548 33.2493
R945 B.n433 B.n122 33.2493
R946 B.n256 B.n255 33.2493
R947 B B.n781 18.0485
R948 B.n723 B.n20 10.6151
R949 B.n727 B.n20 10.6151
R950 B.n728 B.n727 10.6151
R951 B.n729 B.n728 10.6151
R952 B.n729 B.n18 10.6151
R953 B.n733 B.n18 10.6151
R954 B.n734 B.n733 10.6151
R955 B.n735 B.n734 10.6151
R956 B.n735 B.n16 10.6151
R957 B.n739 B.n16 10.6151
R958 B.n740 B.n739 10.6151
R959 B.n741 B.n740 10.6151
R960 B.n741 B.n14 10.6151
R961 B.n745 B.n14 10.6151
R962 B.n746 B.n745 10.6151
R963 B.n747 B.n746 10.6151
R964 B.n747 B.n12 10.6151
R965 B.n751 B.n12 10.6151
R966 B.n752 B.n751 10.6151
R967 B.n753 B.n752 10.6151
R968 B.n753 B.n10 10.6151
R969 B.n757 B.n10 10.6151
R970 B.n758 B.n757 10.6151
R971 B.n759 B.n758 10.6151
R972 B.n759 B.n8 10.6151
R973 B.n763 B.n8 10.6151
R974 B.n764 B.n763 10.6151
R975 B.n765 B.n764 10.6151
R976 B.n765 B.n6 10.6151
R977 B.n769 B.n6 10.6151
R978 B.n770 B.n769 10.6151
R979 B.n771 B.n770 10.6151
R980 B.n771 B.n4 10.6151
R981 B.n775 B.n4 10.6151
R982 B.n776 B.n775 10.6151
R983 B.n777 B.n776 10.6151
R984 B.n777 B.n0 10.6151
R985 B.n722 B.n721 10.6151
R986 B.n721 B.n22 10.6151
R987 B.n717 B.n22 10.6151
R988 B.n717 B.n716 10.6151
R989 B.n716 B.n715 10.6151
R990 B.n715 B.n24 10.6151
R991 B.n711 B.n24 10.6151
R992 B.n711 B.n710 10.6151
R993 B.n710 B.n709 10.6151
R994 B.n709 B.n26 10.6151
R995 B.n705 B.n26 10.6151
R996 B.n705 B.n704 10.6151
R997 B.n704 B.n703 10.6151
R998 B.n703 B.n28 10.6151
R999 B.n699 B.n28 10.6151
R1000 B.n699 B.n698 10.6151
R1001 B.n698 B.n697 10.6151
R1002 B.n697 B.n30 10.6151
R1003 B.n693 B.n30 10.6151
R1004 B.n693 B.n692 10.6151
R1005 B.n692 B.n691 10.6151
R1006 B.n691 B.n32 10.6151
R1007 B.n687 B.n32 10.6151
R1008 B.n687 B.n686 10.6151
R1009 B.n686 B.n685 10.6151
R1010 B.n685 B.n34 10.6151
R1011 B.n681 B.n34 10.6151
R1012 B.n681 B.n680 10.6151
R1013 B.n680 B.n679 10.6151
R1014 B.n679 B.n36 10.6151
R1015 B.n675 B.n36 10.6151
R1016 B.n675 B.n674 10.6151
R1017 B.n674 B.n673 10.6151
R1018 B.n673 B.n38 10.6151
R1019 B.n669 B.n38 10.6151
R1020 B.n669 B.n668 10.6151
R1021 B.n668 B.n667 10.6151
R1022 B.n667 B.n40 10.6151
R1023 B.n663 B.n40 10.6151
R1024 B.n663 B.n662 10.6151
R1025 B.n662 B.n661 10.6151
R1026 B.n661 B.n42 10.6151
R1027 B.n657 B.n42 10.6151
R1028 B.n657 B.n656 10.6151
R1029 B.n656 B.n655 10.6151
R1030 B.n655 B.n44 10.6151
R1031 B.n651 B.n44 10.6151
R1032 B.n651 B.n650 10.6151
R1033 B.n650 B.n649 10.6151
R1034 B.n649 B.n46 10.6151
R1035 B.n645 B.n46 10.6151
R1036 B.n645 B.n644 10.6151
R1037 B.n642 B.n50 10.6151
R1038 B.n638 B.n50 10.6151
R1039 B.n638 B.n637 10.6151
R1040 B.n637 B.n636 10.6151
R1041 B.n636 B.n52 10.6151
R1042 B.n632 B.n52 10.6151
R1043 B.n632 B.n631 10.6151
R1044 B.n631 B.n630 10.6151
R1045 B.n627 B.n626 10.6151
R1046 B.n626 B.n625 10.6151
R1047 B.n625 B.n58 10.6151
R1048 B.n621 B.n58 10.6151
R1049 B.n621 B.n620 10.6151
R1050 B.n620 B.n619 10.6151
R1051 B.n619 B.n60 10.6151
R1052 B.n615 B.n60 10.6151
R1053 B.n615 B.n614 10.6151
R1054 B.n614 B.n613 10.6151
R1055 B.n613 B.n62 10.6151
R1056 B.n609 B.n62 10.6151
R1057 B.n609 B.n608 10.6151
R1058 B.n608 B.n607 10.6151
R1059 B.n607 B.n64 10.6151
R1060 B.n603 B.n64 10.6151
R1061 B.n603 B.n602 10.6151
R1062 B.n602 B.n601 10.6151
R1063 B.n601 B.n66 10.6151
R1064 B.n597 B.n66 10.6151
R1065 B.n597 B.n596 10.6151
R1066 B.n596 B.n595 10.6151
R1067 B.n595 B.n68 10.6151
R1068 B.n591 B.n68 10.6151
R1069 B.n591 B.n590 10.6151
R1070 B.n590 B.n589 10.6151
R1071 B.n589 B.n70 10.6151
R1072 B.n585 B.n70 10.6151
R1073 B.n585 B.n584 10.6151
R1074 B.n584 B.n583 10.6151
R1075 B.n583 B.n72 10.6151
R1076 B.n579 B.n72 10.6151
R1077 B.n579 B.n578 10.6151
R1078 B.n578 B.n577 10.6151
R1079 B.n577 B.n74 10.6151
R1080 B.n573 B.n74 10.6151
R1081 B.n573 B.n572 10.6151
R1082 B.n572 B.n571 10.6151
R1083 B.n571 B.n76 10.6151
R1084 B.n567 B.n76 10.6151
R1085 B.n567 B.n566 10.6151
R1086 B.n566 B.n565 10.6151
R1087 B.n565 B.n78 10.6151
R1088 B.n561 B.n78 10.6151
R1089 B.n561 B.n560 10.6151
R1090 B.n560 B.n559 10.6151
R1091 B.n559 B.n80 10.6151
R1092 B.n555 B.n80 10.6151
R1093 B.n555 B.n554 10.6151
R1094 B.n554 B.n553 10.6151
R1095 B.n553 B.n82 10.6151
R1096 B.n549 B.n82 10.6151
R1097 B.n548 B.n547 10.6151
R1098 B.n547 B.n84 10.6151
R1099 B.n543 B.n84 10.6151
R1100 B.n543 B.n542 10.6151
R1101 B.n542 B.n541 10.6151
R1102 B.n541 B.n86 10.6151
R1103 B.n537 B.n86 10.6151
R1104 B.n537 B.n536 10.6151
R1105 B.n536 B.n535 10.6151
R1106 B.n535 B.n88 10.6151
R1107 B.n531 B.n88 10.6151
R1108 B.n531 B.n530 10.6151
R1109 B.n530 B.n529 10.6151
R1110 B.n529 B.n90 10.6151
R1111 B.n525 B.n90 10.6151
R1112 B.n525 B.n524 10.6151
R1113 B.n524 B.n523 10.6151
R1114 B.n523 B.n92 10.6151
R1115 B.n519 B.n92 10.6151
R1116 B.n519 B.n518 10.6151
R1117 B.n518 B.n517 10.6151
R1118 B.n517 B.n94 10.6151
R1119 B.n513 B.n94 10.6151
R1120 B.n513 B.n512 10.6151
R1121 B.n512 B.n511 10.6151
R1122 B.n511 B.n96 10.6151
R1123 B.n507 B.n96 10.6151
R1124 B.n507 B.n506 10.6151
R1125 B.n506 B.n505 10.6151
R1126 B.n505 B.n98 10.6151
R1127 B.n501 B.n98 10.6151
R1128 B.n501 B.n500 10.6151
R1129 B.n500 B.n499 10.6151
R1130 B.n499 B.n100 10.6151
R1131 B.n495 B.n100 10.6151
R1132 B.n495 B.n494 10.6151
R1133 B.n494 B.n493 10.6151
R1134 B.n493 B.n102 10.6151
R1135 B.n489 B.n102 10.6151
R1136 B.n489 B.n488 10.6151
R1137 B.n488 B.n487 10.6151
R1138 B.n487 B.n104 10.6151
R1139 B.n483 B.n104 10.6151
R1140 B.n483 B.n482 10.6151
R1141 B.n482 B.n481 10.6151
R1142 B.n481 B.n106 10.6151
R1143 B.n477 B.n106 10.6151
R1144 B.n477 B.n476 10.6151
R1145 B.n476 B.n475 10.6151
R1146 B.n475 B.n108 10.6151
R1147 B.n471 B.n108 10.6151
R1148 B.n471 B.n470 10.6151
R1149 B.n470 B.n469 10.6151
R1150 B.n469 B.n110 10.6151
R1151 B.n465 B.n110 10.6151
R1152 B.n465 B.n464 10.6151
R1153 B.n464 B.n463 10.6151
R1154 B.n463 B.n112 10.6151
R1155 B.n459 B.n112 10.6151
R1156 B.n459 B.n458 10.6151
R1157 B.n458 B.n457 10.6151
R1158 B.n457 B.n114 10.6151
R1159 B.n453 B.n114 10.6151
R1160 B.n453 B.n452 10.6151
R1161 B.n452 B.n451 10.6151
R1162 B.n451 B.n116 10.6151
R1163 B.n447 B.n116 10.6151
R1164 B.n447 B.n446 10.6151
R1165 B.n446 B.n445 10.6151
R1166 B.n445 B.n118 10.6151
R1167 B.n441 B.n118 10.6151
R1168 B.n441 B.n440 10.6151
R1169 B.n440 B.n439 10.6151
R1170 B.n439 B.n120 10.6151
R1171 B.n435 B.n120 10.6151
R1172 B.n435 B.n434 10.6151
R1173 B.n434 B.n433 10.6151
R1174 B.n201 B.n1 10.6151
R1175 B.n202 B.n201 10.6151
R1176 B.n203 B.n202 10.6151
R1177 B.n203 B.n198 10.6151
R1178 B.n207 B.n198 10.6151
R1179 B.n208 B.n207 10.6151
R1180 B.n209 B.n208 10.6151
R1181 B.n209 B.n196 10.6151
R1182 B.n213 B.n196 10.6151
R1183 B.n214 B.n213 10.6151
R1184 B.n215 B.n214 10.6151
R1185 B.n215 B.n194 10.6151
R1186 B.n219 B.n194 10.6151
R1187 B.n220 B.n219 10.6151
R1188 B.n221 B.n220 10.6151
R1189 B.n221 B.n192 10.6151
R1190 B.n225 B.n192 10.6151
R1191 B.n226 B.n225 10.6151
R1192 B.n227 B.n226 10.6151
R1193 B.n227 B.n190 10.6151
R1194 B.n231 B.n190 10.6151
R1195 B.n232 B.n231 10.6151
R1196 B.n233 B.n232 10.6151
R1197 B.n233 B.n188 10.6151
R1198 B.n237 B.n188 10.6151
R1199 B.n238 B.n237 10.6151
R1200 B.n239 B.n238 10.6151
R1201 B.n239 B.n186 10.6151
R1202 B.n243 B.n186 10.6151
R1203 B.n244 B.n243 10.6151
R1204 B.n245 B.n244 10.6151
R1205 B.n245 B.n184 10.6151
R1206 B.n249 B.n184 10.6151
R1207 B.n250 B.n249 10.6151
R1208 B.n251 B.n250 10.6151
R1209 B.n251 B.n182 10.6151
R1210 B.n255 B.n182 10.6151
R1211 B.n257 B.n256 10.6151
R1212 B.n257 B.n180 10.6151
R1213 B.n261 B.n180 10.6151
R1214 B.n262 B.n261 10.6151
R1215 B.n263 B.n262 10.6151
R1216 B.n263 B.n178 10.6151
R1217 B.n267 B.n178 10.6151
R1218 B.n268 B.n267 10.6151
R1219 B.n269 B.n268 10.6151
R1220 B.n269 B.n176 10.6151
R1221 B.n273 B.n176 10.6151
R1222 B.n274 B.n273 10.6151
R1223 B.n275 B.n274 10.6151
R1224 B.n275 B.n174 10.6151
R1225 B.n279 B.n174 10.6151
R1226 B.n280 B.n279 10.6151
R1227 B.n281 B.n280 10.6151
R1228 B.n281 B.n172 10.6151
R1229 B.n285 B.n172 10.6151
R1230 B.n286 B.n285 10.6151
R1231 B.n287 B.n286 10.6151
R1232 B.n287 B.n170 10.6151
R1233 B.n291 B.n170 10.6151
R1234 B.n292 B.n291 10.6151
R1235 B.n293 B.n292 10.6151
R1236 B.n293 B.n168 10.6151
R1237 B.n297 B.n168 10.6151
R1238 B.n298 B.n297 10.6151
R1239 B.n299 B.n298 10.6151
R1240 B.n299 B.n166 10.6151
R1241 B.n303 B.n166 10.6151
R1242 B.n304 B.n303 10.6151
R1243 B.n305 B.n304 10.6151
R1244 B.n305 B.n164 10.6151
R1245 B.n309 B.n164 10.6151
R1246 B.n310 B.n309 10.6151
R1247 B.n311 B.n310 10.6151
R1248 B.n311 B.n162 10.6151
R1249 B.n315 B.n162 10.6151
R1250 B.n316 B.n315 10.6151
R1251 B.n317 B.n316 10.6151
R1252 B.n317 B.n160 10.6151
R1253 B.n321 B.n160 10.6151
R1254 B.n322 B.n321 10.6151
R1255 B.n323 B.n322 10.6151
R1256 B.n323 B.n158 10.6151
R1257 B.n327 B.n158 10.6151
R1258 B.n328 B.n327 10.6151
R1259 B.n329 B.n328 10.6151
R1260 B.n329 B.n156 10.6151
R1261 B.n333 B.n156 10.6151
R1262 B.n334 B.n333 10.6151
R1263 B.n336 B.n152 10.6151
R1264 B.n340 B.n152 10.6151
R1265 B.n341 B.n340 10.6151
R1266 B.n342 B.n341 10.6151
R1267 B.n342 B.n150 10.6151
R1268 B.n346 B.n150 10.6151
R1269 B.n347 B.n346 10.6151
R1270 B.n351 B.n347 10.6151
R1271 B.n355 B.n148 10.6151
R1272 B.n356 B.n355 10.6151
R1273 B.n357 B.n356 10.6151
R1274 B.n357 B.n146 10.6151
R1275 B.n361 B.n146 10.6151
R1276 B.n362 B.n361 10.6151
R1277 B.n363 B.n362 10.6151
R1278 B.n363 B.n144 10.6151
R1279 B.n367 B.n144 10.6151
R1280 B.n368 B.n367 10.6151
R1281 B.n369 B.n368 10.6151
R1282 B.n369 B.n142 10.6151
R1283 B.n373 B.n142 10.6151
R1284 B.n374 B.n373 10.6151
R1285 B.n375 B.n374 10.6151
R1286 B.n375 B.n140 10.6151
R1287 B.n379 B.n140 10.6151
R1288 B.n380 B.n379 10.6151
R1289 B.n381 B.n380 10.6151
R1290 B.n381 B.n138 10.6151
R1291 B.n385 B.n138 10.6151
R1292 B.n386 B.n385 10.6151
R1293 B.n387 B.n386 10.6151
R1294 B.n387 B.n136 10.6151
R1295 B.n391 B.n136 10.6151
R1296 B.n392 B.n391 10.6151
R1297 B.n393 B.n392 10.6151
R1298 B.n393 B.n134 10.6151
R1299 B.n397 B.n134 10.6151
R1300 B.n398 B.n397 10.6151
R1301 B.n399 B.n398 10.6151
R1302 B.n399 B.n132 10.6151
R1303 B.n403 B.n132 10.6151
R1304 B.n404 B.n403 10.6151
R1305 B.n405 B.n404 10.6151
R1306 B.n405 B.n130 10.6151
R1307 B.n409 B.n130 10.6151
R1308 B.n410 B.n409 10.6151
R1309 B.n411 B.n410 10.6151
R1310 B.n411 B.n128 10.6151
R1311 B.n415 B.n128 10.6151
R1312 B.n416 B.n415 10.6151
R1313 B.n417 B.n416 10.6151
R1314 B.n417 B.n126 10.6151
R1315 B.n421 B.n126 10.6151
R1316 B.n422 B.n421 10.6151
R1317 B.n423 B.n422 10.6151
R1318 B.n423 B.n124 10.6151
R1319 B.n427 B.n124 10.6151
R1320 B.n428 B.n427 10.6151
R1321 B.n429 B.n428 10.6151
R1322 B.n429 B.n122 10.6151
R1323 B.n781 B.n0 8.11757
R1324 B.n781 B.n1 8.11757
R1325 B.n643 B.n642 6.4005
R1326 B.n630 B.n56 6.4005
R1327 B.n336 B.n335 6.4005
R1328 B.n351 B.n350 6.4005
R1329 B.n644 B.n643 4.21513
R1330 B.n627 B.n56 4.21513
R1331 B.n335 B.n334 4.21513
R1332 B.n350 B.n148 4.21513
C0 VN VTAIL 8.40186f
C1 VP VDD2 0.428871f
C2 B VN 1.14226f
C3 VDD1 VTAIL 9.163691f
C4 B VDD1 2.29918f
C5 VDD2 w_n3034_n4130# 2.54384f
C6 B VTAIL 4.38006f
C7 VN VDD2 8.4885f
C8 VP w_n3034_n4130# 6.13737f
C9 VDD2 VDD1 1.27013f
C10 VP VN 7.29248f
C11 VDD2 VTAIL 9.21075f
C12 VP VDD1 8.76319f
C13 B VDD2 2.36488f
C14 VN w_n3034_n4130# 5.74609f
C15 VP VTAIL 8.41625f
C16 VDD1 w_n3034_n4130# 2.46991f
C17 B VP 1.79378f
C18 VN VDD1 0.150125f
C19 VTAIL w_n3034_n4130# 3.47557f
C20 B w_n3034_n4130# 10.272599f
C21 VDD2 VSUBS 1.925736f
C22 VDD1 VSUBS 2.384128f
C23 VTAIL VSUBS 1.262635f
C24 VN VSUBS 5.6758f
C25 VP VSUBS 2.804684f
C26 B VSUBS 4.61266f
C27 w_n3034_n4130# VSUBS 0.153533p
C28 B.n0 VSUBS 0.006798f
C29 B.n1 VSUBS 0.006798f
C30 B.n2 VSUBS 0.010053f
C31 B.n3 VSUBS 0.007704f
C32 B.n4 VSUBS 0.007704f
C33 B.n5 VSUBS 0.007704f
C34 B.n6 VSUBS 0.007704f
C35 B.n7 VSUBS 0.007704f
C36 B.n8 VSUBS 0.007704f
C37 B.n9 VSUBS 0.007704f
C38 B.n10 VSUBS 0.007704f
C39 B.n11 VSUBS 0.007704f
C40 B.n12 VSUBS 0.007704f
C41 B.n13 VSUBS 0.007704f
C42 B.n14 VSUBS 0.007704f
C43 B.n15 VSUBS 0.007704f
C44 B.n16 VSUBS 0.007704f
C45 B.n17 VSUBS 0.007704f
C46 B.n18 VSUBS 0.007704f
C47 B.n19 VSUBS 0.007704f
C48 B.n20 VSUBS 0.007704f
C49 B.n21 VSUBS 0.018557f
C50 B.n22 VSUBS 0.007704f
C51 B.n23 VSUBS 0.007704f
C52 B.n24 VSUBS 0.007704f
C53 B.n25 VSUBS 0.007704f
C54 B.n26 VSUBS 0.007704f
C55 B.n27 VSUBS 0.007704f
C56 B.n28 VSUBS 0.007704f
C57 B.n29 VSUBS 0.007704f
C58 B.n30 VSUBS 0.007704f
C59 B.n31 VSUBS 0.007704f
C60 B.n32 VSUBS 0.007704f
C61 B.n33 VSUBS 0.007704f
C62 B.n34 VSUBS 0.007704f
C63 B.n35 VSUBS 0.007704f
C64 B.n36 VSUBS 0.007704f
C65 B.n37 VSUBS 0.007704f
C66 B.n38 VSUBS 0.007704f
C67 B.n39 VSUBS 0.007704f
C68 B.n40 VSUBS 0.007704f
C69 B.n41 VSUBS 0.007704f
C70 B.n42 VSUBS 0.007704f
C71 B.n43 VSUBS 0.007704f
C72 B.n44 VSUBS 0.007704f
C73 B.n45 VSUBS 0.007704f
C74 B.n46 VSUBS 0.007704f
C75 B.n47 VSUBS 0.007704f
C76 B.t7 VSUBS 0.581854f
C77 B.t8 VSUBS 0.602709f
C78 B.t6 VSUBS 1.73309f
C79 B.n48 VSUBS 0.308214f
C80 B.n49 VSUBS 0.077659f
C81 B.n50 VSUBS 0.007704f
C82 B.n51 VSUBS 0.007704f
C83 B.n52 VSUBS 0.007704f
C84 B.n53 VSUBS 0.007704f
C85 B.t1 VSUBS 0.581836f
C86 B.t2 VSUBS 0.602694f
C87 B.t0 VSUBS 1.73332f
C88 B.n54 VSUBS 0.308001f
C89 B.n55 VSUBS 0.077677f
C90 B.n56 VSUBS 0.01785f
C91 B.n57 VSUBS 0.007704f
C92 B.n58 VSUBS 0.007704f
C93 B.n59 VSUBS 0.007704f
C94 B.n60 VSUBS 0.007704f
C95 B.n61 VSUBS 0.007704f
C96 B.n62 VSUBS 0.007704f
C97 B.n63 VSUBS 0.007704f
C98 B.n64 VSUBS 0.007704f
C99 B.n65 VSUBS 0.007704f
C100 B.n66 VSUBS 0.007704f
C101 B.n67 VSUBS 0.007704f
C102 B.n68 VSUBS 0.007704f
C103 B.n69 VSUBS 0.007704f
C104 B.n70 VSUBS 0.007704f
C105 B.n71 VSUBS 0.007704f
C106 B.n72 VSUBS 0.007704f
C107 B.n73 VSUBS 0.007704f
C108 B.n74 VSUBS 0.007704f
C109 B.n75 VSUBS 0.007704f
C110 B.n76 VSUBS 0.007704f
C111 B.n77 VSUBS 0.007704f
C112 B.n78 VSUBS 0.007704f
C113 B.n79 VSUBS 0.007704f
C114 B.n80 VSUBS 0.007704f
C115 B.n81 VSUBS 0.007704f
C116 B.n82 VSUBS 0.007704f
C117 B.n83 VSUBS 0.017924f
C118 B.n84 VSUBS 0.007704f
C119 B.n85 VSUBS 0.007704f
C120 B.n86 VSUBS 0.007704f
C121 B.n87 VSUBS 0.007704f
C122 B.n88 VSUBS 0.007704f
C123 B.n89 VSUBS 0.007704f
C124 B.n90 VSUBS 0.007704f
C125 B.n91 VSUBS 0.007704f
C126 B.n92 VSUBS 0.007704f
C127 B.n93 VSUBS 0.007704f
C128 B.n94 VSUBS 0.007704f
C129 B.n95 VSUBS 0.007704f
C130 B.n96 VSUBS 0.007704f
C131 B.n97 VSUBS 0.007704f
C132 B.n98 VSUBS 0.007704f
C133 B.n99 VSUBS 0.007704f
C134 B.n100 VSUBS 0.007704f
C135 B.n101 VSUBS 0.007704f
C136 B.n102 VSUBS 0.007704f
C137 B.n103 VSUBS 0.007704f
C138 B.n104 VSUBS 0.007704f
C139 B.n105 VSUBS 0.007704f
C140 B.n106 VSUBS 0.007704f
C141 B.n107 VSUBS 0.007704f
C142 B.n108 VSUBS 0.007704f
C143 B.n109 VSUBS 0.007704f
C144 B.n110 VSUBS 0.007704f
C145 B.n111 VSUBS 0.007704f
C146 B.n112 VSUBS 0.007704f
C147 B.n113 VSUBS 0.007704f
C148 B.n114 VSUBS 0.007704f
C149 B.n115 VSUBS 0.007704f
C150 B.n116 VSUBS 0.007704f
C151 B.n117 VSUBS 0.007704f
C152 B.n118 VSUBS 0.007704f
C153 B.n119 VSUBS 0.007704f
C154 B.n120 VSUBS 0.007704f
C155 B.n121 VSUBS 0.007704f
C156 B.n122 VSUBS 0.017663f
C157 B.n123 VSUBS 0.007704f
C158 B.n124 VSUBS 0.007704f
C159 B.n125 VSUBS 0.007704f
C160 B.n126 VSUBS 0.007704f
C161 B.n127 VSUBS 0.007704f
C162 B.n128 VSUBS 0.007704f
C163 B.n129 VSUBS 0.007704f
C164 B.n130 VSUBS 0.007704f
C165 B.n131 VSUBS 0.007704f
C166 B.n132 VSUBS 0.007704f
C167 B.n133 VSUBS 0.007704f
C168 B.n134 VSUBS 0.007704f
C169 B.n135 VSUBS 0.007704f
C170 B.n136 VSUBS 0.007704f
C171 B.n137 VSUBS 0.007704f
C172 B.n138 VSUBS 0.007704f
C173 B.n139 VSUBS 0.007704f
C174 B.n140 VSUBS 0.007704f
C175 B.n141 VSUBS 0.007704f
C176 B.n142 VSUBS 0.007704f
C177 B.n143 VSUBS 0.007704f
C178 B.n144 VSUBS 0.007704f
C179 B.n145 VSUBS 0.007704f
C180 B.n146 VSUBS 0.007704f
C181 B.n147 VSUBS 0.007704f
C182 B.n148 VSUBS 0.005381f
C183 B.n149 VSUBS 0.007704f
C184 B.n150 VSUBS 0.007704f
C185 B.n151 VSUBS 0.007704f
C186 B.n152 VSUBS 0.007704f
C187 B.n153 VSUBS 0.007704f
C188 B.t11 VSUBS 0.581854f
C189 B.t10 VSUBS 0.602709f
C190 B.t9 VSUBS 1.73309f
C191 B.n154 VSUBS 0.308214f
C192 B.n155 VSUBS 0.077659f
C193 B.n156 VSUBS 0.007704f
C194 B.n157 VSUBS 0.007704f
C195 B.n158 VSUBS 0.007704f
C196 B.n159 VSUBS 0.007704f
C197 B.n160 VSUBS 0.007704f
C198 B.n161 VSUBS 0.007704f
C199 B.n162 VSUBS 0.007704f
C200 B.n163 VSUBS 0.007704f
C201 B.n164 VSUBS 0.007704f
C202 B.n165 VSUBS 0.007704f
C203 B.n166 VSUBS 0.007704f
C204 B.n167 VSUBS 0.007704f
C205 B.n168 VSUBS 0.007704f
C206 B.n169 VSUBS 0.007704f
C207 B.n170 VSUBS 0.007704f
C208 B.n171 VSUBS 0.007704f
C209 B.n172 VSUBS 0.007704f
C210 B.n173 VSUBS 0.007704f
C211 B.n174 VSUBS 0.007704f
C212 B.n175 VSUBS 0.007704f
C213 B.n176 VSUBS 0.007704f
C214 B.n177 VSUBS 0.007704f
C215 B.n178 VSUBS 0.007704f
C216 B.n179 VSUBS 0.007704f
C217 B.n180 VSUBS 0.007704f
C218 B.n181 VSUBS 0.018557f
C219 B.n182 VSUBS 0.007704f
C220 B.n183 VSUBS 0.007704f
C221 B.n184 VSUBS 0.007704f
C222 B.n185 VSUBS 0.007704f
C223 B.n186 VSUBS 0.007704f
C224 B.n187 VSUBS 0.007704f
C225 B.n188 VSUBS 0.007704f
C226 B.n189 VSUBS 0.007704f
C227 B.n190 VSUBS 0.007704f
C228 B.n191 VSUBS 0.007704f
C229 B.n192 VSUBS 0.007704f
C230 B.n193 VSUBS 0.007704f
C231 B.n194 VSUBS 0.007704f
C232 B.n195 VSUBS 0.007704f
C233 B.n196 VSUBS 0.007704f
C234 B.n197 VSUBS 0.007704f
C235 B.n198 VSUBS 0.007704f
C236 B.n199 VSUBS 0.007704f
C237 B.n200 VSUBS 0.007704f
C238 B.n201 VSUBS 0.007704f
C239 B.n202 VSUBS 0.007704f
C240 B.n203 VSUBS 0.007704f
C241 B.n204 VSUBS 0.007704f
C242 B.n205 VSUBS 0.007704f
C243 B.n206 VSUBS 0.007704f
C244 B.n207 VSUBS 0.007704f
C245 B.n208 VSUBS 0.007704f
C246 B.n209 VSUBS 0.007704f
C247 B.n210 VSUBS 0.007704f
C248 B.n211 VSUBS 0.007704f
C249 B.n212 VSUBS 0.007704f
C250 B.n213 VSUBS 0.007704f
C251 B.n214 VSUBS 0.007704f
C252 B.n215 VSUBS 0.007704f
C253 B.n216 VSUBS 0.007704f
C254 B.n217 VSUBS 0.007704f
C255 B.n218 VSUBS 0.007704f
C256 B.n219 VSUBS 0.007704f
C257 B.n220 VSUBS 0.007704f
C258 B.n221 VSUBS 0.007704f
C259 B.n222 VSUBS 0.007704f
C260 B.n223 VSUBS 0.007704f
C261 B.n224 VSUBS 0.007704f
C262 B.n225 VSUBS 0.007704f
C263 B.n226 VSUBS 0.007704f
C264 B.n227 VSUBS 0.007704f
C265 B.n228 VSUBS 0.007704f
C266 B.n229 VSUBS 0.007704f
C267 B.n230 VSUBS 0.007704f
C268 B.n231 VSUBS 0.007704f
C269 B.n232 VSUBS 0.007704f
C270 B.n233 VSUBS 0.007704f
C271 B.n234 VSUBS 0.007704f
C272 B.n235 VSUBS 0.007704f
C273 B.n236 VSUBS 0.007704f
C274 B.n237 VSUBS 0.007704f
C275 B.n238 VSUBS 0.007704f
C276 B.n239 VSUBS 0.007704f
C277 B.n240 VSUBS 0.007704f
C278 B.n241 VSUBS 0.007704f
C279 B.n242 VSUBS 0.007704f
C280 B.n243 VSUBS 0.007704f
C281 B.n244 VSUBS 0.007704f
C282 B.n245 VSUBS 0.007704f
C283 B.n246 VSUBS 0.007704f
C284 B.n247 VSUBS 0.007704f
C285 B.n248 VSUBS 0.007704f
C286 B.n249 VSUBS 0.007704f
C287 B.n250 VSUBS 0.007704f
C288 B.n251 VSUBS 0.007704f
C289 B.n252 VSUBS 0.007704f
C290 B.n253 VSUBS 0.007704f
C291 B.n254 VSUBS 0.017924f
C292 B.n255 VSUBS 0.017924f
C293 B.n256 VSUBS 0.018557f
C294 B.n257 VSUBS 0.007704f
C295 B.n258 VSUBS 0.007704f
C296 B.n259 VSUBS 0.007704f
C297 B.n260 VSUBS 0.007704f
C298 B.n261 VSUBS 0.007704f
C299 B.n262 VSUBS 0.007704f
C300 B.n263 VSUBS 0.007704f
C301 B.n264 VSUBS 0.007704f
C302 B.n265 VSUBS 0.007704f
C303 B.n266 VSUBS 0.007704f
C304 B.n267 VSUBS 0.007704f
C305 B.n268 VSUBS 0.007704f
C306 B.n269 VSUBS 0.007704f
C307 B.n270 VSUBS 0.007704f
C308 B.n271 VSUBS 0.007704f
C309 B.n272 VSUBS 0.007704f
C310 B.n273 VSUBS 0.007704f
C311 B.n274 VSUBS 0.007704f
C312 B.n275 VSUBS 0.007704f
C313 B.n276 VSUBS 0.007704f
C314 B.n277 VSUBS 0.007704f
C315 B.n278 VSUBS 0.007704f
C316 B.n279 VSUBS 0.007704f
C317 B.n280 VSUBS 0.007704f
C318 B.n281 VSUBS 0.007704f
C319 B.n282 VSUBS 0.007704f
C320 B.n283 VSUBS 0.007704f
C321 B.n284 VSUBS 0.007704f
C322 B.n285 VSUBS 0.007704f
C323 B.n286 VSUBS 0.007704f
C324 B.n287 VSUBS 0.007704f
C325 B.n288 VSUBS 0.007704f
C326 B.n289 VSUBS 0.007704f
C327 B.n290 VSUBS 0.007704f
C328 B.n291 VSUBS 0.007704f
C329 B.n292 VSUBS 0.007704f
C330 B.n293 VSUBS 0.007704f
C331 B.n294 VSUBS 0.007704f
C332 B.n295 VSUBS 0.007704f
C333 B.n296 VSUBS 0.007704f
C334 B.n297 VSUBS 0.007704f
C335 B.n298 VSUBS 0.007704f
C336 B.n299 VSUBS 0.007704f
C337 B.n300 VSUBS 0.007704f
C338 B.n301 VSUBS 0.007704f
C339 B.n302 VSUBS 0.007704f
C340 B.n303 VSUBS 0.007704f
C341 B.n304 VSUBS 0.007704f
C342 B.n305 VSUBS 0.007704f
C343 B.n306 VSUBS 0.007704f
C344 B.n307 VSUBS 0.007704f
C345 B.n308 VSUBS 0.007704f
C346 B.n309 VSUBS 0.007704f
C347 B.n310 VSUBS 0.007704f
C348 B.n311 VSUBS 0.007704f
C349 B.n312 VSUBS 0.007704f
C350 B.n313 VSUBS 0.007704f
C351 B.n314 VSUBS 0.007704f
C352 B.n315 VSUBS 0.007704f
C353 B.n316 VSUBS 0.007704f
C354 B.n317 VSUBS 0.007704f
C355 B.n318 VSUBS 0.007704f
C356 B.n319 VSUBS 0.007704f
C357 B.n320 VSUBS 0.007704f
C358 B.n321 VSUBS 0.007704f
C359 B.n322 VSUBS 0.007704f
C360 B.n323 VSUBS 0.007704f
C361 B.n324 VSUBS 0.007704f
C362 B.n325 VSUBS 0.007704f
C363 B.n326 VSUBS 0.007704f
C364 B.n327 VSUBS 0.007704f
C365 B.n328 VSUBS 0.007704f
C366 B.n329 VSUBS 0.007704f
C367 B.n330 VSUBS 0.007704f
C368 B.n331 VSUBS 0.007704f
C369 B.n332 VSUBS 0.007704f
C370 B.n333 VSUBS 0.007704f
C371 B.n334 VSUBS 0.005381f
C372 B.n335 VSUBS 0.01785f
C373 B.n336 VSUBS 0.006175f
C374 B.n337 VSUBS 0.007704f
C375 B.n338 VSUBS 0.007704f
C376 B.n339 VSUBS 0.007704f
C377 B.n340 VSUBS 0.007704f
C378 B.n341 VSUBS 0.007704f
C379 B.n342 VSUBS 0.007704f
C380 B.n343 VSUBS 0.007704f
C381 B.n344 VSUBS 0.007704f
C382 B.n345 VSUBS 0.007704f
C383 B.n346 VSUBS 0.007704f
C384 B.n347 VSUBS 0.007704f
C385 B.t5 VSUBS 0.581836f
C386 B.t4 VSUBS 0.602694f
C387 B.t3 VSUBS 1.73332f
C388 B.n348 VSUBS 0.308001f
C389 B.n349 VSUBS 0.077677f
C390 B.n350 VSUBS 0.01785f
C391 B.n351 VSUBS 0.006175f
C392 B.n352 VSUBS 0.007704f
C393 B.n353 VSUBS 0.007704f
C394 B.n354 VSUBS 0.007704f
C395 B.n355 VSUBS 0.007704f
C396 B.n356 VSUBS 0.007704f
C397 B.n357 VSUBS 0.007704f
C398 B.n358 VSUBS 0.007704f
C399 B.n359 VSUBS 0.007704f
C400 B.n360 VSUBS 0.007704f
C401 B.n361 VSUBS 0.007704f
C402 B.n362 VSUBS 0.007704f
C403 B.n363 VSUBS 0.007704f
C404 B.n364 VSUBS 0.007704f
C405 B.n365 VSUBS 0.007704f
C406 B.n366 VSUBS 0.007704f
C407 B.n367 VSUBS 0.007704f
C408 B.n368 VSUBS 0.007704f
C409 B.n369 VSUBS 0.007704f
C410 B.n370 VSUBS 0.007704f
C411 B.n371 VSUBS 0.007704f
C412 B.n372 VSUBS 0.007704f
C413 B.n373 VSUBS 0.007704f
C414 B.n374 VSUBS 0.007704f
C415 B.n375 VSUBS 0.007704f
C416 B.n376 VSUBS 0.007704f
C417 B.n377 VSUBS 0.007704f
C418 B.n378 VSUBS 0.007704f
C419 B.n379 VSUBS 0.007704f
C420 B.n380 VSUBS 0.007704f
C421 B.n381 VSUBS 0.007704f
C422 B.n382 VSUBS 0.007704f
C423 B.n383 VSUBS 0.007704f
C424 B.n384 VSUBS 0.007704f
C425 B.n385 VSUBS 0.007704f
C426 B.n386 VSUBS 0.007704f
C427 B.n387 VSUBS 0.007704f
C428 B.n388 VSUBS 0.007704f
C429 B.n389 VSUBS 0.007704f
C430 B.n390 VSUBS 0.007704f
C431 B.n391 VSUBS 0.007704f
C432 B.n392 VSUBS 0.007704f
C433 B.n393 VSUBS 0.007704f
C434 B.n394 VSUBS 0.007704f
C435 B.n395 VSUBS 0.007704f
C436 B.n396 VSUBS 0.007704f
C437 B.n397 VSUBS 0.007704f
C438 B.n398 VSUBS 0.007704f
C439 B.n399 VSUBS 0.007704f
C440 B.n400 VSUBS 0.007704f
C441 B.n401 VSUBS 0.007704f
C442 B.n402 VSUBS 0.007704f
C443 B.n403 VSUBS 0.007704f
C444 B.n404 VSUBS 0.007704f
C445 B.n405 VSUBS 0.007704f
C446 B.n406 VSUBS 0.007704f
C447 B.n407 VSUBS 0.007704f
C448 B.n408 VSUBS 0.007704f
C449 B.n409 VSUBS 0.007704f
C450 B.n410 VSUBS 0.007704f
C451 B.n411 VSUBS 0.007704f
C452 B.n412 VSUBS 0.007704f
C453 B.n413 VSUBS 0.007704f
C454 B.n414 VSUBS 0.007704f
C455 B.n415 VSUBS 0.007704f
C456 B.n416 VSUBS 0.007704f
C457 B.n417 VSUBS 0.007704f
C458 B.n418 VSUBS 0.007704f
C459 B.n419 VSUBS 0.007704f
C460 B.n420 VSUBS 0.007704f
C461 B.n421 VSUBS 0.007704f
C462 B.n422 VSUBS 0.007704f
C463 B.n423 VSUBS 0.007704f
C464 B.n424 VSUBS 0.007704f
C465 B.n425 VSUBS 0.007704f
C466 B.n426 VSUBS 0.007704f
C467 B.n427 VSUBS 0.007704f
C468 B.n428 VSUBS 0.007704f
C469 B.n429 VSUBS 0.007704f
C470 B.n430 VSUBS 0.007704f
C471 B.n431 VSUBS 0.018557f
C472 B.n432 VSUBS 0.017924f
C473 B.n433 VSUBS 0.018818f
C474 B.n434 VSUBS 0.007704f
C475 B.n435 VSUBS 0.007704f
C476 B.n436 VSUBS 0.007704f
C477 B.n437 VSUBS 0.007704f
C478 B.n438 VSUBS 0.007704f
C479 B.n439 VSUBS 0.007704f
C480 B.n440 VSUBS 0.007704f
C481 B.n441 VSUBS 0.007704f
C482 B.n442 VSUBS 0.007704f
C483 B.n443 VSUBS 0.007704f
C484 B.n444 VSUBS 0.007704f
C485 B.n445 VSUBS 0.007704f
C486 B.n446 VSUBS 0.007704f
C487 B.n447 VSUBS 0.007704f
C488 B.n448 VSUBS 0.007704f
C489 B.n449 VSUBS 0.007704f
C490 B.n450 VSUBS 0.007704f
C491 B.n451 VSUBS 0.007704f
C492 B.n452 VSUBS 0.007704f
C493 B.n453 VSUBS 0.007704f
C494 B.n454 VSUBS 0.007704f
C495 B.n455 VSUBS 0.007704f
C496 B.n456 VSUBS 0.007704f
C497 B.n457 VSUBS 0.007704f
C498 B.n458 VSUBS 0.007704f
C499 B.n459 VSUBS 0.007704f
C500 B.n460 VSUBS 0.007704f
C501 B.n461 VSUBS 0.007704f
C502 B.n462 VSUBS 0.007704f
C503 B.n463 VSUBS 0.007704f
C504 B.n464 VSUBS 0.007704f
C505 B.n465 VSUBS 0.007704f
C506 B.n466 VSUBS 0.007704f
C507 B.n467 VSUBS 0.007704f
C508 B.n468 VSUBS 0.007704f
C509 B.n469 VSUBS 0.007704f
C510 B.n470 VSUBS 0.007704f
C511 B.n471 VSUBS 0.007704f
C512 B.n472 VSUBS 0.007704f
C513 B.n473 VSUBS 0.007704f
C514 B.n474 VSUBS 0.007704f
C515 B.n475 VSUBS 0.007704f
C516 B.n476 VSUBS 0.007704f
C517 B.n477 VSUBS 0.007704f
C518 B.n478 VSUBS 0.007704f
C519 B.n479 VSUBS 0.007704f
C520 B.n480 VSUBS 0.007704f
C521 B.n481 VSUBS 0.007704f
C522 B.n482 VSUBS 0.007704f
C523 B.n483 VSUBS 0.007704f
C524 B.n484 VSUBS 0.007704f
C525 B.n485 VSUBS 0.007704f
C526 B.n486 VSUBS 0.007704f
C527 B.n487 VSUBS 0.007704f
C528 B.n488 VSUBS 0.007704f
C529 B.n489 VSUBS 0.007704f
C530 B.n490 VSUBS 0.007704f
C531 B.n491 VSUBS 0.007704f
C532 B.n492 VSUBS 0.007704f
C533 B.n493 VSUBS 0.007704f
C534 B.n494 VSUBS 0.007704f
C535 B.n495 VSUBS 0.007704f
C536 B.n496 VSUBS 0.007704f
C537 B.n497 VSUBS 0.007704f
C538 B.n498 VSUBS 0.007704f
C539 B.n499 VSUBS 0.007704f
C540 B.n500 VSUBS 0.007704f
C541 B.n501 VSUBS 0.007704f
C542 B.n502 VSUBS 0.007704f
C543 B.n503 VSUBS 0.007704f
C544 B.n504 VSUBS 0.007704f
C545 B.n505 VSUBS 0.007704f
C546 B.n506 VSUBS 0.007704f
C547 B.n507 VSUBS 0.007704f
C548 B.n508 VSUBS 0.007704f
C549 B.n509 VSUBS 0.007704f
C550 B.n510 VSUBS 0.007704f
C551 B.n511 VSUBS 0.007704f
C552 B.n512 VSUBS 0.007704f
C553 B.n513 VSUBS 0.007704f
C554 B.n514 VSUBS 0.007704f
C555 B.n515 VSUBS 0.007704f
C556 B.n516 VSUBS 0.007704f
C557 B.n517 VSUBS 0.007704f
C558 B.n518 VSUBS 0.007704f
C559 B.n519 VSUBS 0.007704f
C560 B.n520 VSUBS 0.007704f
C561 B.n521 VSUBS 0.007704f
C562 B.n522 VSUBS 0.007704f
C563 B.n523 VSUBS 0.007704f
C564 B.n524 VSUBS 0.007704f
C565 B.n525 VSUBS 0.007704f
C566 B.n526 VSUBS 0.007704f
C567 B.n527 VSUBS 0.007704f
C568 B.n528 VSUBS 0.007704f
C569 B.n529 VSUBS 0.007704f
C570 B.n530 VSUBS 0.007704f
C571 B.n531 VSUBS 0.007704f
C572 B.n532 VSUBS 0.007704f
C573 B.n533 VSUBS 0.007704f
C574 B.n534 VSUBS 0.007704f
C575 B.n535 VSUBS 0.007704f
C576 B.n536 VSUBS 0.007704f
C577 B.n537 VSUBS 0.007704f
C578 B.n538 VSUBS 0.007704f
C579 B.n539 VSUBS 0.007704f
C580 B.n540 VSUBS 0.007704f
C581 B.n541 VSUBS 0.007704f
C582 B.n542 VSUBS 0.007704f
C583 B.n543 VSUBS 0.007704f
C584 B.n544 VSUBS 0.007704f
C585 B.n545 VSUBS 0.007704f
C586 B.n546 VSUBS 0.007704f
C587 B.n547 VSUBS 0.007704f
C588 B.n548 VSUBS 0.017924f
C589 B.n549 VSUBS 0.018557f
C590 B.n550 VSUBS 0.018557f
C591 B.n551 VSUBS 0.007704f
C592 B.n552 VSUBS 0.007704f
C593 B.n553 VSUBS 0.007704f
C594 B.n554 VSUBS 0.007704f
C595 B.n555 VSUBS 0.007704f
C596 B.n556 VSUBS 0.007704f
C597 B.n557 VSUBS 0.007704f
C598 B.n558 VSUBS 0.007704f
C599 B.n559 VSUBS 0.007704f
C600 B.n560 VSUBS 0.007704f
C601 B.n561 VSUBS 0.007704f
C602 B.n562 VSUBS 0.007704f
C603 B.n563 VSUBS 0.007704f
C604 B.n564 VSUBS 0.007704f
C605 B.n565 VSUBS 0.007704f
C606 B.n566 VSUBS 0.007704f
C607 B.n567 VSUBS 0.007704f
C608 B.n568 VSUBS 0.007704f
C609 B.n569 VSUBS 0.007704f
C610 B.n570 VSUBS 0.007704f
C611 B.n571 VSUBS 0.007704f
C612 B.n572 VSUBS 0.007704f
C613 B.n573 VSUBS 0.007704f
C614 B.n574 VSUBS 0.007704f
C615 B.n575 VSUBS 0.007704f
C616 B.n576 VSUBS 0.007704f
C617 B.n577 VSUBS 0.007704f
C618 B.n578 VSUBS 0.007704f
C619 B.n579 VSUBS 0.007704f
C620 B.n580 VSUBS 0.007704f
C621 B.n581 VSUBS 0.007704f
C622 B.n582 VSUBS 0.007704f
C623 B.n583 VSUBS 0.007704f
C624 B.n584 VSUBS 0.007704f
C625 B.n585 VSUBS 0.007704f
C626 B.n586 VSUBS 0.007704f
C627 B.n587 VSUBS 0.007704f
C628 B.n588 VSUBS 0.007704f
C629 B.n589 VSUBS 0.007704f
C630 B.n590 VSUBS 0.007704f
C631 B.n591 VSUBS 0.007704f
C632 B.n592 VSUBS 0.007704f
C633 B.n593 VSUBS 0.007704f
C634 B.n594 VSUBS 0.007704f
C635 B.n595 VSUBS 0.007704f
C636 B.n596 VSUBS 0.007704f
C637 B.n597 VSUBS 0.007704f
C638 B.n598 VSUBS 0.007704f
C639 B.n599 VSUBS 0.007704f
C640 B.n600 VSUBS 0.007704f
C641 B.n601 VSUBS 0.007704f
C642 B.n602 VSUBS 0.007704f
C643 B.n603 VSUBS 0.007704f
C644 B.n604 VSUBS 0.007704f
C645 B.n605 VSUBS 0.007704f
C646 B.n606 VSUBS 0.007704f
C647 B.n607 VSUBS 0.007704f
C648 B.n608 VSUBS 0.007704f
C649 B.n609 VSUBS 0.007704f
C650 B.n610 VSUBS 0.007704f
C651 B.n611 VSUBS 0.007704f
C652 B.n612 VSUBS 0.007704f
C653 B.n613 VSUBS 0.007704f
C654 B.n614 VSUBS 0.007704f
C655 B.n615 VSUBS 0.007704f
C656 B.n616 VSUBS 0.007704f
C657 B.n617 VSUBS 0.007704f
C658 B.n618 VSUBS 0.007704f
C659 B.n619 VSUBS 0.007704f
C660 B.n620 VSUBS 0.007704f
C661 B.n621 VSUBS 0.007704f
C662 B.n622 VSUBS 0.007704f
C663 B.n623 VSUBS 0.007704f
C664 B.n624 VSUBS 0.007704f
C665 B.n625 VSUBS 0.007704f
C666 B.n626 VSUBS 0.007704f
C667 B.n627 VSUBS 0.005381f
C668 B.n628 VSUBS 0.007704f
C669 B.n629 VSUBS 0.007704f
C670 B.n630 VSUBS 0.006175f
C671 B.n631 VSUBS 0.007704f
C672 B.n632 VSUBS 0.007704f
C673 B.n633 VSUBS 0.007704f
C674 B.n634 VSUBS 0.007704f
C675 B.n635 VSUBS 0.007704f
C676 B.n636 VSUBS 0.007704f
C677 B.n637 VSUBS 0.007704f
C678 B.n638 VSUBS 0.007704f
C679 B.n639 VSUBS 0.007704f
C680 B.n640 VSUBS 0.007704f
C681 B.n641 VSUBS 0.007704f
C682 B.n642 VSUBS 0.006175f
C683 B.n643 VSUBS 0.01785f
C684 B.n644 VSUBS 0.005381f
C685 B.n645 VSUBS 0.007704f
C686 B.n646 VSUBS 0.007704f
C687 B.n647 VSUBS 0.007704f
C688 B.n648 VSUBS 0.007704f
C689 B.n649 VSUBS 0.007704f
C690 B.n650 VSUBS 0.007704f
C691 B.n651 VSUBS 0.007704f
C692 B.n652 VSUBS 0.007704f
C693 B.n653 VSUBS 0.007704f
C694 B.n654 VSUBS 0.007704f
C695 B.n655 VSUBS 0.007704f
C696 B.n656 VSUBS 0.007704f
C697 B.n657 VSUBS 0.007704f
C698 B.n658 VSUBS 0.007704f
C699 B.n659 VSUBS 0.007704f
C700 B.n660 VSUBS 0.007704f
C701 B.n661 VSUBS 0.007704f
C702 B.n662 VSUBS 0.007704f
C703 B.n663 VSUBS 0.007704f
C704 B.n664 VSUBS 0.007704f
C705 B.n665 VSUBS 0.007704f
C706 B.n666 VSUBS 0.007704f
C707 B.n667 VSUBS 0.007704f
C708 B.n668 VSUBS 0.007704f
C709 B.n669 VSUBS 0.007704f
C710 B.n670 VSUBS 0.007704f
C711 B.n671 VSUBS 0.007704f
C712 B.n672 VSUBS 0.007704f
C713 B.n673 VSUBS 0.007704f
C714 B.n674 VSUBS 0.007704f
C715 B.n675 VSUBS 0.007704f
C716 B.n676 VSUBS 0.007704f
C717 B.n677 VSUBS 0.007704f
C718 B.n678 VSUBS 0.007704f
C719 B.n679 VSUBS 0.007704f
C720 B.n680 VSUBS 0.007704f
C721 B.n681 VSUBS 0.007704f
C722 B.n682 VSUBS 0.007704f
C723 B.n683 VSUBS 0.007704f
C724 B.n684 VSUBS 0.007704f
C725 B.n685 VSUBS 0.007704f
C726 B.n686 VSUBS 0.007704f
C727 B.n687 VSUBS 0.007704f
C728 B.n688 VSUBS 0.007704f
C729 B.n689 VSUBS 0.007704f
C730 B.n690 VSUBS 0.007704f
C731 B.n691 VSUBS 0.007704f
C732 B.n692 VSUBS 0.007704f
C733 B.n693 VSUBS 0.007704f
C734 B.n694 VSUBS 0.007704f
C735 B.n695 VSUBS 0.007704f
C736 B.n696 VSUBS 0.007704f
C737 B.n697 VSUBS 0.007704f
C738 B.n698 VSUBS 0.007704f
C739 B.n699 VSUBS 0.007704f
C740 B.n700 VSUBS 0.007704f
C741 B.n701 VSUBS 0.007704f
C742 B.n702 VSUBS 0.007704f
C743 B.n703 VSUBS 0.007704f
C744 B.n704 VSUBS 0.007704f
C745 B.n705 VSUBS 0.007704f
C746 B.n706 VSUBS 0.007704f
C747 B.n707 VSUBS 0.007704f
C748 B.n708 VSUBS 0.007704f
C749 B.n709 VSUBS 0.007704f
C750 B.n710 VSUBS 0.007704f
C751 B.n711 VSUBS 0.007704f
C752 B.n712 VSUBS 0.007704f
C753 B.n713 VSUBS 0.007704f
C754 B.n714 VSUBS 0.007704f
C755 B.n715 VSUBS 0.007704f
C756 B.n716 VSUBS 0.007704f
C757 B.n717 VSUBS 0.007704f
C758 B.n718 VSUBS 0.007704f
C759 B.n719 VSUBS 0.007704f
C760 B.n720 VSUBS 0.007704f
C761 B.n721 VSUBS 0.007704f
C762 B.n722 VSUBS 0.018557f
C763 B.n723 VSUBS 0.017924f
C764 B.n724 VSUBS 0.017924f
C765 B.n725 VSUBS 0.007704f
C766 B.n726 VSUBS 0.007704f
C767 B.n727 VSUBS 0.007704f
C768 B.n728 VSUBS 0.007704f
C769 B.n729 VSUBS 0.007704f
C770 B.n730 VSUBS 0.007704f
C771 B.n731 VSUBS 0.007704f
C772 B.n732 VSUBS 0.007704f
C773 B.n733 VSUBS 0.007704f
C774 B.n734 VSUBS 0.007704f
C775 B.n735 VSUBS 0.007704f
C776 B.n736 VSUBS 0.007704f
C777 B.n737 VSUBS 0.007704f
C778 B.n738 VSUBS 0.007704f
C779 B.n739 VSUBS 0.007704f
C780 B.n740 VSUBS 0.007704f
C781 B.n741 VSUBS 0.007704f
C782 B.n742 VSUBS 0.007704f
C783 B.n743 VSUBS 0.007704f
C784 B.n744 VSUBS 0.007704f
C785 B.n745 VSUBS 0.007704f
C786 B.n746 VSUBS 0.007704f
C787 B.n747 VSUBS 0.007704f
C788 B.n748 VSUBS 0.007704f
C789 B.n749 VSUBS 0.007704f
C790 B.n750 VSUBS 0.007704f
C791 B.n751 VSUBS 0.007704f
C792 B.n752 VSUBS 0.007704f
C793 B.n753 VSUBS 0.007704f
C794 B.n754 VSUBS 0.007704f
C795 B.n755 VSUBS 0.007704f
C796 B.n756 VSUBS 0.007704f
C797 B.n757 VSUBS 0.007704f
C798 B.n758 VSUBS 0.007704f
C799 B.n759 VSUBS 0.007704f
C800 B.n760 VSUBS 0.007704f
C801 B.n761 VSUBS 0.007704f
C802 B.n762 VSUBS 0.007704f
C803 B.n763 VSUBS 0.007704f
C804 B.n764 VSUBS 0.007704f
C805 B.n765 VSUBS 0.007704f
C806 B.n766 VSUBS 0.007704f
C807 B.n767 VSUBS 0.007704f
C808 B.n768 VSUBS 0.007704f
C809 B.n769 VSUBS 0.007704f
C810 B.n770 VSUBS 0.007704f
C811 B.n771 VSUBS 0.007704f
C812 B.n772 VSUBS 0.007704f
C813 B.n773 VSUBS 0.007704f
C814 B.n774 VSUBS 0.007704f
C815 B.n775 VSUBS 0.007704f
C816 B.n776 VSUBS 0.007704f
C817 B.n777 VSUBS 0.007704f
C818 B.n778 VSUBS 0.007704f
C819 B.n779 VSUBS 0.010053f
C820 B.n780 VSUBS 0.010709f
C821 B.n781 VSUBS 0.021297f
C822 VDD1.t0 VSUBS 3.65408f
C823 VDD1.t1 VSUBS 3.65271f
C824 VDD1.t2 VSUBS 0.341632f
C825 VDD1.t5 VSUBS 0.341632f
C826 VDD1.n0 VSUBS 2.8043f
C827 VDD1.n1 VSUBS 4.00935f
C828 VDD1.t4 VSUBS 0.341632f
C829 VDD1.t3 VSUBS 0.341632f
C830 VDD1.n2 VSUBS 2.79893f
C831 VDD1.n3 VSUBS 3.55712f
C832 VP.n0 VSUBS 0.041478f
C833 VP.t0 VSUBS 3.06889f
C834 VP.n1 VSUBS 0.026086f
C835 VP.n2 VSUBS 0.031461f
C836 VP.t3 VSUBS 3.06889f
C837 VP.n3 VSUBS 0.063433f
C838 VP.n4 VSUBS 0.031461f
C839 VP.t4 VSUBS 3.06889f
C840 VP.n5 VSUBS 1.17568f
C841 VP.n6 VSUBS 0.041478f
C842 VP.t2 VSUBS 3.06889f
C843 VP.n7 VSUBS 0.026086f
C844 VP.n8 VSUBS 0.269427f
C845 VP.t1 VSUBS 3.06889f
C846 VP.t5 VSUBS 3.27289f
C847 VP.n9 VSUBS 1.14368f
C848 VP.n10 VSUBS 1.15666f
C849 VP.n11 VSUBS 0.044161f
C850 VP.n12 VSUBS 0.063433f
C851 VP.n13 VSUBS 0.031461f
C852 VP.n14 VSUBS 0.031461f
C853 VP.n15 VSUBS 0.031461f
C854 VP.n16 VSUBS 0.06097f
C855 VP.n17 VSUBS 0.048792f
C856 VP.n18 VSUBS 1.17568f
C857 VP.n19 VSUBS 1.75332f
C858 VP.n20 VSUBS 1.77584f
C859 VP.n21 VSUBS 0.041478f
C860 VP.n22 VSUBS 0.048792f
C861 VP.n23 VSUBS 0.06097f
C862 VP.n24 VSUBS 0.026086f
C863 VP.n25 VSUBS 0.031461f
C864 VP.n26 VSUBS 0.031461f
C865 VP.n27 VSUBS 0.031461f
C866 VP.n28 VSUBS 0.044161f
C867 VP.n29 VSUBS 1.07439f
C868 VP.n30 VSUBS 0.044161f
C869 VP.n31 VSUBS 0.063433f
C870 VP.n32 VSUBS 0.031461f
C871 VP.n33 VSUBS 0.031461f
C872 VP.n34 VSUBS 0.031461f
C873 VP.n35 VSUBS 0.06097f
C874 VP.n36 VSUBS 0.048792f
C875 VP.n37 VSUBS 1.17568f
C876 VP.n38 VSUBS 0.042986f
C877 VDD2.t1 VSUBS 3.63678f
C878 VDD2.t3 VSUBS 0.340142f
C879 VDD2.t0 VSUBS 0.340142f
C880 VDD2.n0 VSUBS 2.79206f
C881 VDD2.n1 VSUBS 3.86388f
C882 VDD2.t5 VSUBS 3.62043f
C883 VDD2.n2 VSUBS 3.57563f
C884 VDD2.t2 VSUBS 0.340142f
C885 VDD2.t4 VSUBS 0.340142f
C886 VDD2.n3 VSUBS 2.79202f
C887 VTAIL.t9 VSUBS 0.347969f
C888 VTAIL.t7 VSUBS 0.347969f
C889 VTAIL.n0 VSUBS 2.69169f
C890 VTAIL.n1 VSUBS 0.849384f
C891 VTAIL.t1 VSUBS 3.52222f
C892 VTAIL.n2 VSUBS 1.11234f
C893 VTAIL.t10 VSUBS 0.347969f
C894 VTAIL.t3 VSUBS 0.347969f
C895 VTAIL.n3 VSUBS 2.69169f
C896 VTAIL.n4 VSUBS 2.85261f
C897 VTAIL.t8 VSUBS 0.347969f
C898 VTAIL.t4 VSUBS 0.347969f
C899 VTAIL.n5 VSUBS 2.6917f
C900 VTAIL.n6 VSUBS 2.8526f
C901 VTAIL.t6 VSUBS 3.52225f
C902 VTAIL.n7 VSUBS 1.11231f
C903 VTAIL.t11 VSUBS 0.347969f
C904 VTAIL.t2 VSUBS 0.347969f
C905 VTAIL.n8 VSUBS 2.6917f
C906 VTAIL.n9 VSUBS 0.99386f
C907 VTAIL.t0 VSUBS 3.52222f
C908 VTAIL.n10 VSUBS 2.77148f
C909 VTAIL.t5 VSUBS 3.52222f
C910 VTAIL.n11 VSUBS 2.71635f
C911 VN.n0 VSUBS 0.04047f
C912 VN.t5 VSUBS 2.99436f
C913 VN.n1 VSUBS 0.025452f
C914 VN.n2 VSUBS 0.262883f
C915 VN.t2 VSUBS 2.99436f
C916 VN.t4 VSUBS 3.1934f
C917 VN.n3 VSUBS 1.11591f
C918 VN.n4 VSUBS 1.12857f
C919 VN.n5 VSUBS 0.043088f
C920 VN.n6 VSUBS 0.061892f
C921 VN.n7 VSUBS 0.030697f
C922 VN.n8 VSUBS 0.030697f
C923 VN.n9 VSUBS 0.030697f
C924 VN.n10 VSUBS 0.059489f
C925 VN.n11 VSUBS 0.047607f
C926 VN.n12 VSUBS 1.14713f
C927 VN.n13 VSUBS 0.041942f
C928 VN.n14 VSUBS 0.04047f
C929 VN.t0 VSUBS 2.99436f
C930 VN.n15 VSUBS 0.025452f
C931 VN.n16 VSUBS 0.262883f
C932 VN.t3 VSUBS 2.99436f
C933 VN.t1 VSUBS 3.1934f
C934 VN.n17 VSUBS 1.11591f
C935 VN.n18 VSUBS 1.12857f
C936 VN.n19 VSUBS 0.043088f
C937 VN.n20 VSUBS 0.061892f
C938 VN.n21 VSUBS 0.030697f
C939 VN.n22 VSUBS 0.030697f
C940 VN.n23 VSUBS 0.030697f
C941 VN.n24 VSUBS 0.059489f
C942 VN.n25 VSUBS 0.047607f
C943 VN.n26 VSUBS 1.14713f
C944 VN.n27 VSUBS 1.72722f
.ends

