* NGSPICE file created from opamp_sample_0009.ext - technology: sky130A

.subckt opamp_sample_0009 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 GND.t80 CS_BIAS.t18 CS_BIAS.t19 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X1 a_n7516_558.t24 DIFFPAIR_BIAS.t4 GND.t87 GND.t86 sky130_fd_pr__nfet_01v8 ad=2.5128 pd=8.42 as=2.5128 ps=8.42 w=3.49 l=2.02
X2 GND.t185 GND.t183 GND.t184 GND.t110 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X3 GND.t79 CS_BIAS.t16 CS_BIAS.t17 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X4 a_n11545_9494.t25 a_n11545_9494.t24 a_n11689_9690.t11 VDD.t92 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X5 VDD.t67 VDD.t65 VDD.t66 VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X6 GND.t182 GND.t180 GND.t181 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X7 a_n11545_9494.t7 VP.t0 a_n7516_558.t13 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X8 VOUT.t54 CS_BIAS.t20 GND.t78 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X9 VOUT.t53 CS_BIAS.t21 GND.t77 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X10 CS_BIAS.t15 CS_BIAS.t14 GND.t75 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X11 VOUT.t52 CS_BIAS.t22 GND.t76 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X12 a_n11545_9494.t26 VP.t1 a_n7516_558.t22 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X13 VDD.t108 a_n11545_9494.t28 a_n11689_9690.t12 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X14 a_n17362_8608.t18 a_n11545_9494.t29 a_n7386_8166.t0 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X15 a_n17362_8608.t17 a_n11545_9494.t30 a_n7386_8166.t2 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X16 a_n11689_9690.t14 a_n11545_9494.t31 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X17 GND.t74 CS_BIAS.t23 VOUT.t51 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X18 VDD.t64 VDD.t62 VDD.t63 VDD.t50 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X19 a_n11689_9690.t10 a_n11545_9494.t18 a_n11545_9494.t19 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X20 GND.t179 GND.t177 GND.t178 GND.t147 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.42
X21 VDD.t61 VDD.t59 VDD.t60 VDD.t17 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X22 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t187 GND.t186 sky130_fd_pr__nfet_01v8 ad=2.5128 pd=8.42 as=2.5128 ps=8.42 w=3.49 l=2.02
X23 GND.t176 GND.t174 GND.t175 GND.t134 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X24 VDD.t58 VDD.t56 VDD.t57 VDD.t13 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X25 a_n17362_8608.t19 VN.t0 a_n7516_558.t21 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X26 VOUT.t50 CS_BIAS.t24 GND.t73 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X27 VOUT.t49 CS_BIAS.t25 GND.t72 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X28 a_n11689_9690.t13 a_n11545_9494.t32 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X29 VOUT.t48 CS_BIAS.t26 GND.t71 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X30 GND.t70 CS_BIAS.t27 VOUT.t47 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X31 GND.t69 CS_BIAS.t28 VOUT.t46 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X32 a_n17362_8608.t10 VN.t1 a_n7516_558.t20 GND.t85 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.42
X33 VOUT.t45 CS_BIAS.t29 GND.t64 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X34 VOUT.t44 CS_BIAS.t30 GND.t65 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X35 GND.t68 CS_BIAS.t31 VOUT.t43 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X36 VOUT.t42 CS_BIAS.t32 GND.t67 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X37 GND.t66 CS_BIAS.t33 VOUT.t41 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X38 a_n7516_558.t19 VN.t2 a_n17362_8608.t9 GND.t10 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.42
X39 VDD.t55 VDD.t53 VDD.t54 VDD.t37 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X40 a_n7516_558.t4 VP.t2 a_n11545_9494.t1 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X41 VOUT.t58 a_n7386_8166.t16 sky130_fd_pr__cap_mim_m3_1 l=14.21 w=18.87
X42 a_n17362_8608.t8 VN.t3 a_n7516_558.t18 GND.t81 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X43 CS_BIAS.t7 CS_BIAS.t6 GND.t63 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X44 a_n7386_8166.t13 a_n11545_9494.t33 a_n17362_8608.t16 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X45 VOUT.t40 CS_BIAS.t34 GND.t62 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X46 GND.t173 GND.t171 GND.t172 GND.t126 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X47 VOUT.t56 a_n17362_8608.t20 VDD.t11 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.2507 pd=4.45 as=2.7288 ps=9.02 w=3.79 l=4.11
X48 VDD.t52 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X49 VOUT.t39 CS_BIAS.t35 GND.t61 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X50 VDD.t48 VDD.t46 VDD.t47 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X51 a_n7516_558.t17 VN.t4 a_n17362_8608.t7 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X52 VDD.t101 a_n11545_9494.t34 a_n11689_9690.t3 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X53 VOUT.t55 a_n17362_8608.t21 VDD.t10 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.2507 pd=4.45 as=2.7288 ps=9.02 w=3.79 l=4.11
X54 GND.t170 GND.t168 GND.t169 GND.t134 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X55 GND.t167 GND.t165 GND.t166 GND.t134 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X56 GND.t164 GND.t162 GND.t163 GND.t134 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X57 CS_BIAS.t5 CS_BIAS.t4 GND.t58 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X58 a_n11545_9494.t23 a_n11545_9494.t22 a_n11689_9690.t9 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X59 GND.t161 GND.t159 GND.t160 GND.t110 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X60 a_n17362_8608.t6 VN.t5 a_n7516_558.t16 GND.t84 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.42
X61 a_n7516_558.t6 VN.t6 a_n17362_8608.t4 GND.t5 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.42
X62 VDD.t45 VDD.t43 VDD.t44 VDD.t29 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X63 a_n13259_9690# a_n13259_9690# a_n13259_9690# VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=2.9952 ps=11.2 w=2.08 l=5.77
X64 a_n7386_8166.t12 a_n11545_9494.t35 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X65 GND.t60 CS_BIAS.t36 VOUT.t38 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X66 VOUT.t37 CS_BIAS.t37 GND.t59 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X67 GND.t57 CS_BIAS.t38 VOUT.t36 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X68 GND.t56 CS_BIAS.t39 VOUT.t35 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X69 VOUT.t34 CS_BIAS.t40 GND.t55 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X70 VOUT.t33 CS_BIAS.t41 GND.t54 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X71 VOUT.t32 CS_BIAS.t42 GND.t53 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X72 CS_BIAS.t3 CS_BIAS.t2 GND.t52 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X73 GND.t158 GND.t156 GND.t157 GND.t134 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X74 CS_BIAS.t1 CS_BIAS.t0 GND.t51 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X75 a_n11689_9690.t8 a_n11545_9494.t20 a_n11545_9494.t21 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X76 a_n7516_558.t10 VP.t3 a_n11545_9494.t4 GND.t10 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.42
X77 GND.t155 GND.t153 GND.t154 GND.t126 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X78 VDD.t97 a_n11545_9494.t36 a_n7386_8166.t11 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X79 VDD.t42 VDD.t40 VDD.t41 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X80 VDD.t39 VDD.t36 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X81 GND.t152 GND.t150 GND.t151 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X82 GND.t149 GND.t146 GND.t148 GND.t147 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.42
X83 GND.t145 GND.t143 GND.t144 GND.t126 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X84 GND.t50 CS_BIAS.t43 VOUT.t31 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X85 GND.t142 GND.t140 GND.t141 GND.t126 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X86 GND.t139 GND.t137 GND.t138 GND.t126 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X87 a_n7386_8166.t15 a_n11545_9494.t37 a_n17362_8608.t15 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X88 a_n11689_9690.t15 a_n11545_9494.t38 VDD.t94 VDD.t93 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X89 GND.t49 CS_BIAS.t44 VOUT.t30 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X90 a_n7386_8166.t3 a_n11545_9494.t39 a_n17362_8608.t14 VDD.t92 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X91 VOUT.t29 CS_BIAS.t45 GND.t48 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X92 VOUT.t28 CS_BIAS.t46 GND.t47 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X93 VOUT.t27 CS_BIAS.t47 GND.t46 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X94 GND.t45 CS_BIAS.t48 VOUT.t26 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X95 VOUT.t25 CS_BIAS.t49 GND.t43 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X96 VDD.t109 a_n17362_8608.t22 VOUT.t57 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=1.2507 ps=4.45 w=3.79 l=4.11
X97 VOUT.t24 CS_BIAS.t50 GND.t42 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X98 a_n7516_558.t7 VN.t7 a_n17362_8608.t5 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X99 a_n7516_558.t0 VN.t8 a_n17362_8608.t0 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X100 a_n17362_8608.t1 VN.t9 a_n7516_558.t1 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X101 a_n11545_9494.t27 VP.t4 a_n7516_558.t25 GND.t85 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.42
X102 a_n11545_9494.t17 a_n11545_9494.t16 a_n11689_9690.t7 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X103 VDD.t35 VDD.t32 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X104 a_n7386_8166.t4 a_n11545_9494.t40 a_n17362_8608.t13 VDD.t83 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X105 VDD.t31 VDD.t28 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X106 a_n11689_9690.t6 a_n11545_9494.t10 a_n11545_9494.t11 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X107 VDD.t89 a_n11545_9494.t41 a_n11689_9690.t0 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X108 GND.t41 CS_BIAS.t12 CS_BIAS.t13 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X109 a_n7516_558.t5 VN.t10 a_n17362_8608.t3 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X110 a_n7516_558.t3 VP.t5 a_n11545_9494.t0 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X111 a_n17362_8608.t12 a_n11545_9494.t42 a_n7386_8166.t14 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X112 a_n7516_558.t9 VP.t6 a_n11545_9494.t3 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X113 GND.t136 GND.t133 GND.t135 GND.t134 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X114 VOUT.t4 a_n17362_8608.t23 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.2507 pd=4.45 as=2.7288 ps=9.02 w=3.79 l=4.11
X115 VOUT.t59 a_n7386_8166.t16 sky130_fd_pr__cap_mim_m3_1 l=14.21 w=18.87
X116 VDD.t87 a_n11545_9494.t43 a_n11689_9690.t1 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X117 a_n7386_8166.t10 a_n11545_9494.t44 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X118 CS_BIAS.t11 CS_BIAS.t10 GND.t40 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X119 a_n11545_9494.t13 a_n11545_9494.t12 a_n11689_9690.t5 VDD.t83 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.77
X120 a_n17362_8608.t2 VN.t11 a_n7516_558.t2 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X121 GND.t39 CS_BIAS.t51 VOUT.t23 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X122 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t83 GND.t82 sky130_fd_pr__nfet_01v8 ad=2.5128 pd=8.42 as=2.5128 ps=8.42 w=3.49 l=2.02
X123 VDD.t82 a_n11545_9494.t45 a_n7386_8166.t9 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X124 VDD.t80 a_n11545_9494.t46 a_n7386_8166.t8 VDD.t79 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.77
X125 a_11817_9690# a_11817_9690# a_11817_9690# VDD.t68 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=2.9952 ps=11.2 w=2.08 l=5.77
X126 GND.t38 CS_BIAS.t52 VOUT.t22 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X127 GND.t37 CS_BIAS.t8 CS_BIAS.t9 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X128 GND.t132 GND.t129 GND.t131 GND.t130 sky130_fd_pr__nfet_01v8 ad=2.5128 pd=8.42 as=0 ps=0 w=3.49 l=2.02
X129 GND.t36 CS_BIAS.t53 VOUT.t21 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X130 VOUT.t20 CS_BIAS.t54 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X131 a_n11545_9494.t8 VP.t7 a_n7516_558.t14 GND.t84 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.42
X132 VDD.t27 VDD.t24 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X133 GND.t128 GND.t125 GND.t127 GND.t126 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X134 a_n17362_8608.t11 a_n11545_9494.t47 a_n7386_8166.t1 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X135 GND.t124 GND.t122 GND.t123 GND.t110 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X136 GND.t121 GND.t119 GND.t120 GND.t110 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X137 VDD.t23 VDD.t20 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X138 GND.t118 GND.t116 GND.t117 GND.t110 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X139 VDD.t2 a_n17362_8608.t24 VOUT.t0 VDD.t1 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=1.2507 ps=4.45 w=3.79 l=4.11
X140 VOUT.t1 a_n17362_8608.t25 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.2507 pd=4.45 as=2.7288 ps=9.02 w=3.79 l=4.11
X141 VDD.t19 VDD.t16 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.77
X142 VDD.t77 a_n11545_9494.t48 a_n7386_8166.t7 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X143 VOUT.t19 CS_BIAS.t55 GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X144 GND.t31 CS_BIAS.t56 VOUT.t18 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X145 a_n7516_558.t11 VP.t8 a_n11545_9494.t5 GND.t5 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.42
X146 a_n11689_9690.t2 a_n11545_9494.t49 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X147 GND.t115 GND.t113 GND.t114 GND.t106 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.42
X148 GND.t112 GND.t109 GND.t111 GND.t110 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X149 a_n11545_9494.t6 VP.t9 a_n7516_558.t12 GND.t81 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X150 GND.t29 CS_BIAS.t57 VOUT.t17 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X151 a_n11689_9690.t4 a_n11545_9494.t14 a_n11545_9494.t15 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X152 VOUT.t16 CS_BIAS.t58 GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X153 GND.t28 CS_BIAS.t59 VOUT.t15 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X154 GND.t27 CS_BIAS.t60 VOUT.t14 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X155 GND.t108 GND.t105 GND.t107 GND.t106 sky130_fd_pr__nfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.42
X156 VDD.t7 a_n17362_8608.t26 VOUT.t3 VDD.t1 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=1.2507 ps=4.45 w=3.79 l=4.11
X157 GND.t24 CS_BIAS.t61 VOUT.t13 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X158 VOUT.t12 CS_BIAS.t62 GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=1.4976 ps=5.6 w=2.08 l=5.72
X159 GND.t104 GND.t102 GND.t103 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X160 GND.t101 GND.t99 GND.t100 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X161 GND.t98 GND.t96 GND.t97 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X162 VOUT.t11 CS_BIAS.t63 GND.t18 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X163 GND.t20 CS_BIAS.t64 VOUT.t10 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.72
X164 VOUT.t9 CS_BIAS.t65 GND.t17 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X165 VOUT.t8 CS_BIAS.t66 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X166 a_n7386_8166.t6 a_n11545_9494.t50 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X167 GND.t95 GND.t92 GND.t94 GND.t93 sky130_fd_pr__nfet_01v8 ad=2.5128 pd=8.42 as=0 ps=0 w=3.49 l=2.02
X168 a_n7516_558.t23 DIFFPAIR_BIAS.t5 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=2.5128 pd=8.42 as=2.5128 ps=8.42 w=3.49 l=2.02
X169 VDD.t15 VDD.t12 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=0 ps=0 w=3.79 l=4.11
X170 a_n11545_9494.t2 VP.t10 a_n7516_558.t8 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X171 a_n7386_8166.t5 a_n11545_9494.t51 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8 ad=0.6864 pd=2.74 as=0.6864 ps=2.74 w=2.08 l=5.77
X172 VDD.t6 a_n17362_8608.t27 VOUT.t2 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.7288 pd=9.02 as=1.2507 ps=4.45 w=3.79 l=4.11
X173 VOUT.t7 CS_BIAS.t67 GND.t14 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X174 GND.t91 GND.t88 GND.t90 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0 ps=0 w=2.08 l=5.72
X175 a_n7516_558.t15 VP.t11 a_n11545_9494.t9 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.42
X176 VOUT.t6 CS_BIAS.t68 GND.t13 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
X177 VOUT.t5 CS_BIAS.t69 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=5.6 as=0.6864 ps=2.74 w=2.08 l=5.72
R0 CS_BIAS.n511 CS_BIAS.n510 161.3
R1 CS_BIAS.n509 CS_BIAS.n430 161.3
R2 CS_BIAS.n508 CS_BIAS.n507 161.3
R3 CS_BIAS.n506 CS_BIAS.n431 161.3
R4 CS_BIAS.n505 CS_BIAS.n504 161.3
R5 CS_BIAS.n503 CS_BIAS.n432 161.3
R6 CS_BIAS.n502 CS_BIAS.n501 161.3
R7 CS_BIAS.n500 CS_BIAS.n433 161.3
R8 CS_BIAS.n499 CS_BIAS.n498 161.3
R9 CS_BIAS.n497 CS_BIAS.n434 161.3
R10 CS_BIAS.n496 CS_BIAS.n495 161.3
R11 CS_BIAS.n494 CS_BIAS.n435 161.3
R12 CS_BIAS.n493 CS_BIAS.n492 161.3
R13 CS_BIAS.n490 CS_BIAS.n436 161.3
R14 CS_BIAS.n489 CS_BIAS.n488 161.3
R15 CS_BIAS.n487 CS_BIAS.n437 161.3
R16 CS_BIAS.n486 CS_BIAS.n485 161.3
R17 CS_BIAS.n484 CS_BIAS.n438 161.3
R18 CS_BIAS.n483 CS_BIAS.n482 161.3
R19 CS_BIAS.n481 CS_BIAS.n439 161.3
R20 CS_BIAS.n480 CS_BIAS.n479 161.3
R21 CS_BIAS.n478 CS_BIAS.n440 161.3
R22 CS_BIAS.n477 CS_BIAS.n476 161.3
R23 CS_BIAS.n475 CS_BIAS.n441 161.3
R24 CS_BIAS.n474 CS_BIAS.n473 161.3
R25 CS_BIAS.n472 CS_BIAS.n442 161.3
R26 CS_BIAS.n470 CS_BIAS.n469 161.3
R27 CS_BIAS.n468 CS_BIAS.n443 161.3
R28 CS_BIAS.n467 CS_BIAS.n466 161.3
R29 CS_BIAS.n465 CS_BIAS.n444 161.3
R30 CS_BIAS.n464 CS_BIAS.n463 161.3
R31 CS_BIAS.n462 CS_BIAS.n445 161.3
R32 CS_BIAS.n461 CS_BIAS.n460 161.3
R33 CS_BIAS.n459 CS_BIAS.n446 161.3
R34 CS_BIAS.n458 CS_BIAS.n457 161.3
R35 CS_BIAS.n456 CS_BIAS.n447 161.3
R36 CS_BIAS.n455 CS_BIAS.n454 161.3
R37 CS_BIAS.n453 CS_BIAS.n448 161.3
R38 CS_BIAS.n452 CS_BIAS.n451 161.3
R39 CS_BIAS.n367 CS_BIAS.n366 161.3
R40 CS_BIAS.n368 CS_BIAS.n363 161.3
R41 CS_BIAS.n370 CS_BIAS.n369 161.3
R42 CS_BIAS.n371 CS_BIAS.n362 161.3
R43 CS_BIAS.n373 CS_BIAS.n372 161.3
R44 CS_BIAS.n374 CS_BIAS.n361 161.3
R45 CS_BIAS.n376 CS_BIAS.n375 161.3
R46 CS_BIAS.n377 CS_BIAS.n360 161.3
R47 CS_BIAS.n379 CS_BIAS.n378 161.3
R48 CS_BIAS.n380 CS_BIAS.n359 161.3
R49 CS_BIAS.n382 CS_BIAS.n381 161.3
R50 CS_BIAS.n383 CS_BIAS.n358 161.3
R51 CS_BIAS.n385 CS_BIAS.n384 161.3
R52 CS_BIAS.n387 CS_BIAS.n357 161.3
R53 CS_BIAS.n389 CS_BIAS.n388 161.3
R54 CS_BIAS.n390 CS_BIAS.n356 161.3
R55 CS_BIAS.n392 CS_BIAS.n391 161.3
R56 CS_BIAS.n393 CS_BIAS.n355 161.3
R57 CS_BIAS.n395 CS_BIAS.n394 161.3
R58 CS_BIAS.n396 CS_BIAS.n354 161.3
R59 CS_BIAS.n398 CS_BIAS.n397 161.3
R60 CS_BIAS.n399 CS_BIAS.n353 161.3
R61 CS_BIAS.n401 CS_BIAS.n400 161.3
R62 CS_BIAS.n402 CS_BIAS.n352 161.3
R63 CS_BIAS.n404 CS_BIAS.n403 161.3
R64 CS_BIAS.n405 CS_BIAS.n351 161.3
R65 CS_BIAS.n408 CS_BIAS.n407 161.3
R66 CS_BIAS.n409 CS_BIAS.n350 161.3
R67 CS_BIAS.n411 CS_BIAS.n410 161.3
R68 CS_BIAS.n412 CS_BIAS.n349 161.3
R69 CS_BIAS.n414 CS_BIAS.n413 161.3
R70 CS_BIAS.n415 CS_BIAS.n348 161.3
R71 CS_BIAS.n417 CS_BIAS.n416 161.3
R72 CS_BIAS.n418 CS_BIAS.n347 161.3
R73 CS_BIAS.n420 CS_BIAS.n419 161.3
R74 CS_BIAS.n421 CS_BIAS.n346 161.3
R75 CS_BIAS.n423 CS_BIAS.n422 161.3
R76 CS_BIAS.n424 CS_BIAS.n345 161.3
R77 CS_BIAS.n426 CS_BIAS.n425 161.3
R78 CS_BIAS.n282 CS_BIAS.n281 161.3
R79 CS_BIAS.n283 CS_BIAS.n278 161.3
R80 CS_BIAS.n285 CS_BIAS.n284 161.3
R81 CS_BIAS.n286 CS_BIAS.n277 161.3
R82 CS_BIAS.n288 CS_BIAS.n287 161.3
R83 CS_BIAS.n289 CS_BIAS.n276 161.3
R84 CS_BIAS.n291 CS_BIAS.n290 161.3
R85 CS_BIAS.n292 CS_BIAS.n275 161.3
R86 CS_BIAS.n294 CS_BIAS.n293 161.3
R87 CS_BIAS.n295 CS_BIAS.n274 161.3
R88 CS_BIAS.n297 CS_BIAS.n296 161.3
R89 CS_BIAS.n298 CS_BIAS.n273 161.3
R90 CS_BIAS.n300 CS_BIAS.n299 161.3
R91 CS_BIAS.n302 CS_BIAS.n272 161.3
R92 CS_BIAS.n304 CS_BIAS.n303 161.3
R93 CS_BIAS.n305 CS_BIAS.n271 161.3
R94 CS_BIAS.n307 CS_BIAS.n306 161.3
R95 CS_BIAS.n308 CS_BIAS.n270 161.3
R96 CS_BIAS.n310 CS_BIAS.n309 161.3
R97 CS_BIAS.n311 CS_BIAS.n269 161.3
R98 CS_BIAS.n313 CS_BIAS.n312 161.3
R99 CS_BIAS.n314 CS_BIAS.n268 161.3
R100 CS_BIAS.n316 CS_BIAS.n315 161.3
R101 CS_BIAS.n317 CS_BIAS.n267 161.3
R102 CS_BIAS.n319 CS_BIAS.n318 161.3
R103 CS_BIAS.n320 CS_BIAS.n266 161.3
R104 CS_BIAS.n323 CS_BIAS.n322 161.3
R105 CS_BIAS.n324 CS_BIAS.n265 161.3
R106 CS_BIAS.n326 CS_BIAS.n325 161.3
R107 CS_BIAS.n327 CS_BIAS.n264 161.3
R108 CS_BIAS.n329 CS_BIAS.n328 161.3
R109 CS_BIAS.n330 CS_BIAS.n263 161.3
R110 CS_BIAS.n332 CS_BIAS.n331 161.3
R111 CS_BIAS.n333 CS_BIAS.n262 161.3
R112 CS_BIAS.n335 CS_BIAS.n334 161.3
R113 CS_BIAS.n336 CS_BIAS.n261 161.3
R114 CS_BIAS.n338 CS_BIAS.n337 161.3
R115 CS_BIAS.n339 CS_BIAS.n260 161.3
R116 CS_BIAS.n341 CS_BIAS.n340 161.3
R117 CS_BIAS.n197 CS_BIAS.n196 161.3
R118 CS_BIAS.n198 CS_BIAS.n193 161.3
R119 CS_BIAS.n200 CS_BIAS.n199 161.3
R120 CS_BIAS.n201 CS_BIAS.n192 161.3
R121 CS_BIAS.n203 CS_BIAS.n202 161.3
R122 CS_BIAS.n204 CS_BIAS.n191 161.3
R123 CS_BIAS.n206 CS_BIAS.n205 161.3
R124 CS_BIAS.n207 CS_BIAS.n190 161.3
R125 CS_BIAS.n209 CS_BIAS.n208 161.3
R126 CS_BIAS.n210 CS_BIAS.n189 161.3
R127 CS_BIAS.n212 CS_BIAS.n211 161.3
R128 CS_BIAS.n213 CS_BIAS.n188 161.3
R129 CS_BIAS.n215 CS_BIAS.n214 161.3
R130 CS_BIAS.n217 CS_BIAS.n187 161.3
R131 CS_BIAS.n219 CS_BIAS.n218 161.3
R132 CS_BIAS.n220 CS_BIAS.n186 161.3
R133 CS_BIAS.n222 CS_BIAS.n221 161.3
R134 CS_BIAS.n223 CS_BIAS.n185 161.3
R135 CS_BIAS.n225 CS_BIAS.n224 161.3
R136 CS_BIAS.n226 CS_BIAS.n184 161.3
R137 CS_BIAS.n228 CS_BIAS.n227 161.3
R138 CS_BIAS.n229 CS_BIAS.n183 161.3
R139 CS_BIAS.n231 CS_BIAS.n230 161.3
R140 CS_BIAS.n232 CS_BIAS.n182 161.3
R141 CS_BIAS.n234 CS_BIAS.n233 161.3
R142 CS_BIAS.n235 CS_BIAS.n181 161.3
R143 CS_BIAS.n238 CS_BIAS.n237 161.3
R144 CS_BIAS.n239 CS_BIAS.n180 161.3
R145 CS_BIAS.n241 CS_BIAS.n240 161.3
R146 CS_BIAS.n242 CS_BIAS.n179 161.3
R147 CS_BIAS.n244 CS_BIAS.n243 161.3
R148 CS_BIAS.n245 CS_BIAS.n178 161.3
R149 CS_BIAS.n247 CS_BIAS.n246 161.3
R150 CS_BIAS.n248 CS_BIAS.n177 161.3
R151 CS_BIAS.n250 CS_BIAS.n249 161.3
R152 CS_BIAS.n251 CS_BIAS.n176 161.3
R153 CS_BIAS.n253 CS_BIAS.n252 161.3
R154 CS_BIAS.n254 CS_BIAS.n175 161.3
R155 CS_BIAS.n256 CS_BIAS.n255 161.3
R156 CS_BIAS.n38 CS_BIAS.n37 161.3
R157 CS_BIAS.n39 CS_BIAS.n34 161.3
R158 CS_BIAS.n41 CS_BIAS.n40 161.3
R159 CS_BIAS.n42 CS_BIAS.n33 161.3
R160 CS_BIAS.n44 CS_BIAS.n43 161.3
R161 CS_BIAS.n45 CS_BIAS.n32 161.3
R162 CS_BIAS.n47 CS_BIAS.n46 161.3
R163 CS_BIAS.n48 CS_BIAS.n31 161.3
R164 CS_BIAS.n50 CS_BIAS.n49 161.3
R165 CS_BIAS.n51 CS_BIAS.n30 161.3
R166 CS_BIAS.n53 CS_BIAS.n52 161.3
R167 CS_BIAS.n54 CS_BIAS.n29 161.3
R168 CS_BIAS.n56 CS_BIAS.n55 161.3
R169 CS_BIAS.n58 CS_BIAS.n28 161.3
R170 CS_BIAS.n60 CS_BIAS.n59 161.3
R171 CS_BIAS.n61 CS_BIAS.n27 161.3
R172 CS_BIAS.n63 CS_BIAS.n62 161.3
R173 CS_BIAS.n64 CS_BIAS.n26 161.3
R174 CS_BIAS.n66 CS_BIAS.n65 161.3
R175 CS_BIAS.n67 CS_BIAS.n25 161.3
R176 CS_BIAS.n69 CS_BIAS.n68 161.3
R177 CS_BIAS.n70 CS_BIAS.n24 161.3
R178 CS_BIAS.n72 CS_BIAS.n71 161.3
R179 CS_BIAS.n73 CS_BIAS.n23 161.3
R180 CS_BIAS.n75 CS_BIAS.n74 161.3
R181 CS_BIAS.n76 CS_BIAS.n22 161.3
R182 CS_BIAS.n79 CS_BIAS.n78 161.3
R183 CS_BIAS.n80 CS_BIAS.n21 161.3
R184 CS_BIAS.n82 CS_BIAS.n81 161.3
R185 CS_BIAS.n83 CS_BIAS.n20 161.3
R186 CS_BIAS.n85 CS_BIAS.n84 161.3
R187 CS_BIAS.n86 CS_BIAS.n19 161.3
R188 CS_BIAS.n88 CS_BIAS.n87 161.3
R189 CS_BIAS.n89 CS_BIAS.n18 161.3
R190 CS_BIAS.n91 CS_BIAS.n90 161.3
R191 CS_BIAS.n92 CS_BIAS.n17 161.3
R192 CS_BIAS.n94 CS_BIAS.n93 161.3
R193 CS_BIAS.n95 CS_BIAS.n16 161.3
R194 CS_BIAS.n97 CS_BIAS.n96 161.3
R195 CS_BIAS.n113 CS_BIAS.n112 161.3
R196 CS_BIAS.n114 CS_BIAS.n109 161.3
R197 CS_BIAS.n116 CS_BIAS.n115 161.3
R198 CS_BIAS.n117 CS_BIAS.n108 161.3
R199 CS_BIAS.n119 CS_BIAS.n118 161.3
R200 CS_BIAS.n120 CS_BIAS.n107 161.3
R201 CS_BIAS.n122 CS_BIAS.n121 161.3
R202 CS_BIAS.n123 CS_BIAS.n106 161.3
R203 CS_BIAS.n125 CS_BIAS.n124 161.3
R204 CS_BIAS.n126 CS_BIAS.n105 161.3
R205 CS_BIAS.n128 CS_BIAS.n127 161.3
R206 CS_BIAS.n129 CS_BIAS.n14 161.3
R207 CS_BIAS.n131 CS_BIAS.n130 161.3
R208 CS_BIAS.n133 CS_BIAS.n13 161.3
R209 CS_BIAS.n135 CS_BIAS.n134 161.3
R210 CS_BIAS.n136 CS_BIAS.n12 161.3
R211 CS_BIAS.n138 CS_BIAS.n137 161.3
R212 CS_BIAS.n139 CS_BIAS.n11 161.3
R213 CS_BIAS.n141 CS_BIAS.n140 161.3
R214 CS_BIAS.n142 CS_BIAS.n10 161.3
R215 CS_BIAS.n144 CS_BIAS.n143 161.3
R216 CS_BIAS.n145 CS_BIAS.n9 161.3
R217 CS_BIAS.n147 CS_BIAS.n146 161.3
R218 CS_BIAS.n148 CS_BIAS.n8 161.3
R219 CS_BIAS.n150 CS_BIAS.n149 161.3
R220 CS_BIAS.n151 CS_BIAS.n7 161.3
R221 CS_BIAS.n154 CS_BIAS.n153 161.3
R222 CS_BIAS.n155 CS_BIAS.n6 161.3
R223 CS_BIAS.n157 CS_BIAS.n156 161.3
R224 CS_BIAS.n158 CS_BIAS.n5 161.3
R225 CS_BIAS.n160 CS_BIAS.n159 161.3
R226 CS_BIAS.n161 CS_BIAS.n4 161.3
R227 CS_BIAS.n163 CS_BIAS.n162 161.3
R228 CS_BIAS.n164 CS_BIAS.n3 161.3
R229 CS_BIAS.n166 CS_BIAS.n165 161.3
R230 CS_BIAS.n167 CS_BIAS.n2 161.3
R231 CS_BIAS.n169 CS_BIAS.n168 161.3
R232 CS_BIAS.n170 CS_BIAS.n1 161.3
R233 CS_BIAS.n172 CS_BIAS.n171 161.3
R234 CS_BIAS.n1025 CS_BIAS.n1024 161.3
R235 CS_BIAS.n1023 CS_BIAS.n944 161.3
R236 CS_BIAS.n1022 CS_BIAS.n1021 161.3
R237 CS_BIAS.n1020 CS_BIAS.n945 161.3
R238 CS_BIAS.n1019 CS_BIAS.n1018 161.3
R239 CS_BIAS.n1017 CS_BIAS.n946 161.3
R240 CS_BIAS.n1016 CS_BIAS.n1015 161.3
R241 CS_BIAS.n1014 CS_BIAS.n947 161.3
R242 CS_BIAS.n1013 CS_BIAS.n1012 161.3
R243 CS_BIAS.n1011 CS_BIAS.n948 161.3
R244 CS_BIAS.n1010 CS_BIAS.n1009 161.3
R245 CS_BIAS.n1008 CS_BIAS.n949 161.3
R246 CS_BIAS.n1007 CS_BIAS.n1006 161.3
R247 CS_BIAS.n1004 CS_BIAS.n950 161.3
R248 CS_BIAS.n1003 CS_BIAS.n1002 161.3
R249 CS_BIAS.n1001 CS_BIAS.n951 161.3
R250 CS_BIAS.n1000 CS_BIAS.n999 161.3
R251 CS_BIAS.n998 CS_BIAS.n952 161.3
R252 CS_BIAS.n997 CS_BIAS.n996 161.3
R253 CS_BIAS.n995 CS_BIAS.n953 161.3
R254 CS_BIAS.n994 CS_BIAS.n993 161.3
R255 CS_BIAS.n992 CS_BIAS.n954 161.3
R256 CS_BIAS.n991 CS_BIAS.n990 161.3
R257 CS_BIAS.n989 CS_BIAS.n955 161.3
R258 CS_BIAS.n988 CS_BIAS.n987 161.3
R259 CS_BIAS.n986 CS_BIAS.n956 161.3
R260 CS_BIAS.n984 CS_BIAS.n983 161.3
R261 CS_BIAS.n982 CS_BIAS.n957 161.3
R262 CS_BIAS.n981 CS_BIAS.n980 161.3
R263 CS_BIAS.n979 CS_BIAS.n958 161.3
R264 CS_BIAS.n978 CS_BIAS.n977 161.3
R265 CS_BIAS.n976 CS_BIAS.n959 161.3
R266 CS_BIAS.n975 CS_BIAS.n974 161.3
R267 CS_BIAS.n973 CS_BIAS.n960 161.3
R268 CS_BIAS.n972 CS_BIAS.n971 161.3
R269 CS_BIAS.n970 CS_BIAS.n961 161.3
R270 CS_BIAS.n969 CS_BIAS.n968 161.3
R271 CS_BIAS.n967 CS_BIAS.n962 161.3
R272 CS_BIAS.n966 CS_BIAS.n965 161.3
R273 CS_BIAS.n940 CS_BIAS.n939 161.3
R274 CS_BIAS.n938 CS_BIAS.n859 161.3
R275 CS_BIAS.n937 CS_BIAS.n936 161.3
R276 CS_BIAS.n935 CS_BIAS.n860 161.3
R277 CS_BIAS.n934 CS_BIAS.n933 161.3
R278 CS_BIAS.n932 CS_BIAS.n861 161.3
R279 CS_BIAS.n931 CS_BIAS.n930 161.3
R280 CS_BIAS.n929 CS_BIAS.n862 161.3
R281 CS_BIAS.n928 CS_BIAS.n927 161.3
R282 CS_BIAS.n926 CS_BIAS.n863 161.3
R283 CS_BIAS.n925 CS_BIAS.n924 161.3
R284 CS_BIAS.n923 CS_BIAS.n864 161.3
R285 CS_BIAS.n922 CS_BIAS.n921 161.3
R286 CS_BIAS.n919 CS_BIAS.n865 161.3
R287 CS_BIAS.n918 CS_BIAS.n917 161.3
R288 CS_BIAS.n916 CS_BIAS.n866 161.3
R289 CS_BIAS.n915 CS_BIAS.n914 161.3
R290 CS_BIAS.n913 CS_BIAS.n867 161.3
R291 CS_BIAS.n912 CS_BIAS.n911 161.3
R292 CS_BIAS.n910 CS_BIAS.n868 161.3
R293 CS_BIAS.n909 CS_BIAS.n908 161.3
R294 CS_BIAS.n907 CS_BIAS.n869 161.3
R295 CS_BIAS.n906 CS_BIAS.n905 161.3
R296 CS_BIAS.n904 CS_BIAS.n870 161.3
R297 CS_BIAS.n903 CS_BIAS.n902 161.3
R298 CS_BIAS.n901 CS_BIAS.n871 161.3
R299 CS_BIAS.n899 CS_BIAS.n898 161.3
R300 CS_BIAS.n897 CS_BIAS.n872 161.3
R301 CS_BIAS.n896 CS_BIAS.n895 161.3
R302 CS_BIAS.n894 CS_BIAS.n873 161.3
R303 CS_BIAS.n893 CS_BIAS.n892 161.3
R304 CS_BIAS.n891 CS_BIAS.n874 161.3
R305 CS_BIAS.n890 CS_BIAS.n889 161.3
R306 CS_BIAS.n888 CS_BIAS.n875 161.3
R307 CS_BIAS.n887 CS_BIAS.n886 161.3
R308 CS_BIAS.n885 CS_BIAS.n876 161.3
R309 CS_BIAS.n884 CS_BIAS.n883 161.3
R310 CS_BIAS.n882 CS_BIAS.n877 161.3
R311 CS_BIAS.n881 CS_BIAS.n880 161.3
R312 CS_BIAS.n855 CS_BIAS.n854 161.3
R313 CS_BIAS.n853 CS_BIAS.n774 161.3
R314 CS_BIAS.n852 CS_BIAS.n851 161.3
R315 CS_BIAS.n850 CS_BIAS.n775 161.3
R316 CS_BIAS.n849 CS_BIAS.n848 161.3
R317 CS_BIAS.n847 CS_BIAS.n776 161.3
R318 CS_BIAS.n846 CS_BIAS.n845 161.3
R319 CS_BIAS.n844 CS_BIAS.n777 161.3
R320 CS_BIAS.n843 CS_BIAS.n842 161.3
R321 CS_BIAS.n841 CS_BIAS.n778 161.3
R322 CS_BIAS.n840 CS_BIAS.n839 161.3
R323 CS_BIAS.n838 CS_BIAS.n779 161.3
R324 CS_BIAS.n837 CS_BIAS.n836 161.3
R325 CS_BIAS.n834 CS_BIAS.n780 161.3
R326 CS_BIAS.n833 CS_BIAS.n832 161.3
R327 CS_BIAS.n831 CS_BIAS.n781 161.3
R328 CS_BIAS.n830 CS_BIAS.n829 161.3
R329 CS_BIAS.n828 CS_BIAS.n782 161.3
R330 CS_BIAS.n827 CS_BIAS.n826 161.3
R331 CS_BIAS.n825 CS_BIAS.n783 161.3
R332 CS_BIAS.n824 CS_BIAS.n823 161.3
R333 CS_BIAS.n822 CS_BIAS.n784 161.3
R334 CS_BIAS.n821 CS_BIAS.n820 161.3
R335 CS_BIAS.n819 CS_BIAS.n785 161.3
R336 CS_BIAS.n818 CS_BIAS.n817 161.3
R337 CS_BIAS.n816 CS_BIAS.n786 161.3
R338 CS_BIAS.n814 CS_BIAS.n813 161.3
R339 CS_BIAS.n812 CS_BIAS.n787 161.3
R340 CS_BIAS.n811 CS_BIAS.n810 161.3
R341 CS_BIAS.n809 CS_BIAS.n788 161.3
R342 CS_BIAS.n808 CS_BIAS.n807 161.3
R343 CS_BIAS.n806 CS_BIAS.n789 161.3
R344 CS_BIAS.n805 CS_BIAS.n804 161.3
R345 CS_BIAS.n803 CS_BIAS.n790 161.3
R346 CS_BIAS.n802 CS_BIAS.n801 161.3
R347 CS_BIAS.n800 CS_BIAS.n791 161.3
R348 CS_BIAS.n799 CS_BIAS.n798 161.3
R349 CS_BIAS.n797 CS_BIAS.n792 161.3
R350 CS_BIAS.n796 CS_BIAS.n795 161.3
R351 CS_BIAS.n770 CS_BIAS.n769 161.3
R352 CS_BIAS.n768 CS_BIAS.n689 161.3
R353 CS_BIAS.n767 CS_BIAS.n766 161.3
R354 CS_BIAS.n765 CS_BIAS.n690 161.3
R355 CS_BIAS.n764 CS_BIAS.n763 161.3
R356 CS_BIAS.n762 CS_BIAS.n691 161.3
R357 CS_BIAS.n761 CS_BIAS.n760 161.3
R358 CS_BIAS.n759 CS_BIAS.n692 161.3
R359 CS_BIAS.n758 CS_BIAS.n757 161.3
R360 CS_BIAS.n756 CS_BIAS.n693 161.3
R361 CS_BIAS.n755 CS_BIAS.n754 161.3
R362 CS_BIAS.n753 CS_BIAS.n694 161.3
R363 CS_BIAS.n752 CS_BIAS.n751 161.3
R364 CS_BIAS.n749 CS_BIAS.n695 161.3
R365 CS_BIAS.n748 CS_BIAS.n747 161.3
R366 CS_BIAS.n746 CS_BIAS.n696 161.3
R367 CS_BIAS.n745 CS_BIAS.n744 161.3
R368 CS_BIAS.n743 CS_BIAS.n697 161.3
R369 CS_BIAS.n742 CS_BIAS.n741 161.3
R370 CS_BIAS.n740 CS_BIAS.n698 161.3
R371 CS_BIAS.n739 CS_BIAS.n738 161.3
R372 CS_BIAS.n737 CS_BIAS.n699 161.3
R373 CS_BIAS.n736 CS_BIAS.n735 161.3
R374 CS_BIAS.n734 CS_BIAS.n700 161.3
R375 CS_BIAS.n733 CS_BIAS.n732 161.3
R376 CS_BIAS.n731 CS_BIAS.n701 161.3
R377 CS_BIAS.n729 CS_BIAS.n728 161.3
R378 CS_BIAS.n727 CS_BIAS.n702 161.3
R379 CS_BIAS.n726 CS_BIAS.n725 161.3
R380 CS_BIAS.n724 CS_BIAS.n703 161.3
R381 CS_BIAS.n723 CS_BIAS.n722 161.3
R382 CS_BIAS.n721 CS_BIAS.n704 161.3
R383 CS_BIAS.n720 CS_BIAS.n719 161.3
R384 CS_BIAS.n718 CS_BIAS.n705 161.3
R385 CS_BIAS.n717 CS_BIAS.n716 161.3
R386 CS_BIAS.n715 CS_BIAS.n706 161.3
R387 CS_BIAS.n714 CS_BIAS.n713 161.3
R388 CS_BIAS.n712 CS_BIAS.n707 161.3
R389 CS_BIAS.n711 CS_BIAS.n710 161.3
R390 CS_BIAS.n638 CS_BIAS.n637 161.3
R391 CS_BIAS.n636 CS_BIAS.n557 161.3
R392 CS_BIAS.n635 CS_BIAS.n634 161.3
R393 CS_BIAS.n633 CS_BIAS.n558 161.3
R394 CS_BIAS.n632 CS_BIAS.n631 161.3
R395 CS_BIAS.n630 CS_BIAS.n559 161.3
R396 CS_BIAS.n629 CS_BIAS.n628 161.3
R397 CS_BIAS.n627 CS_BIAS.n560 161.3
R398 CS_BIAS.n626 CS_BIAS.n625 161.3
R399 CS_BIAS.n624 CS_BIAS.n561 161.3
R400 CS_BIAS.n623 CS_BIAS.n622 161.3
R401 CS_BIAS.n621 CS_BIAS.n562 161.3
R402 CS_BIAS.n620 CS_BIAS.n619 161.3
R403 CS_BIAS.n617 CS_BIAS.n563 161.3
R404 CS_BIAS.n616 CS_BIAS.n615 161.3
R405 CS_BIAS.n614 CS_BIAS.n564 161.3
R406 CS_BIAS.n613 CS_BIAS.n612 161.3
R407 CS_BIAS.n611 CS_BIAS.n565 161.3
R408 CS_BIAS.n610 CS_BIAS.n609 161.3
R409 CS_BIAS.n608 CS_BIAS.n566 161.3
R410 CS_BIAS.n607 CS_BIAS.n606 161.3
R411 CS_BIAS.n605 CS_BIAS.n567 161.3
R412 CS_BIAS.n604 CS_BIAS.n603 161.3
R413 CS_BIAS.n602 CS_BIAS.n568 161.3
R414 CS_BIAS.n601 CS_BIAS.n600 161.3
R415 CS_BIAS.n599 CS_BIAS.n569 161.3
R416 CS_BIAS.n597 CS_BIAS.n596 161.3
R417 CS_BIAS.n595 CS_BIAS.n570 161.3
R418 CS_BIAS.n594 CS_BIAS.n593 161.3
R419 CS_BIAS.n592 CS_BIAS.n571 161.3
R420 CS_BIAS.n591 CS_BIAS.n590 161.3
R421 CS_BIAS.n589 CS_BIAS.n572 161.3
R422 CS_BIAS.n588 CS_BIAS.n587 161.3
R423 CS_BIAS.n586 CS_BIAS.n573 161.3
R424 CS_BIAS.n585 CS_BIAS.n584 161.3
R425 CS_BIAS.n583 CS_BIAS.n574 161.3
R426 CS_BIAS.n582 CS_BIAS.n581 161.3
R427 CS_BIAS.n580 CS_BIAS.n575 161.3
R428 CS_BIAS.n579 CS_BIAS.n578 161.3
R429 CS_BIAS.n645 CS_BIAS.n644 161.3
R430 CS_BIAS.n553 CS_BIAS.n528 161.3
R431 CS_BIAS.n552 CS_BIAS.n551 161.3
R432 CS_BIAS.n550 CS_BIAS.n529 161.3
R433 CS_BIAS.n549 CS_BIAS.n548 161.3
R434 CS_BIAS.n547 CS_BIAS.n530 161.3
R435 CS_BIAS.n546 CS_BIAS.n545 161.3
R436 CS_BIAS.n544 CS_BIAS.n531 161.3
R437 CS_BIAS.n543 CS_BIAS.n542 161.3
R438 CS_BIAS.n541 CS_BIAS.n532 161.3
R439 CS_BIAS.n540 CS_BIAS.n539 161.3
R440 CS_BIAS.n538 CS_BIAS.n533 161.3
R441 CS_BIAS.n537 CS_BIAS.n536 161.3
R442 CS_BIAS.n686 CS_BIAS.n685 161.3
R443 CS_BIAS.n684 CS_BIAS.n515 161.3
R444 CS_BIAS.n683 CS_BIAS.n682 161.3
R445 CS_BIAS.n681 CS_BIAS.n516 161.3
R446 CS_BIAS.n680 CS_BIAS.n679 161.3
R447 CS_BIAS.n678 CS_BIAS.n517 161.3
R448 CS_BIAS.n677 CS_BIAS.n676 161.3
R449 CS_BIAS.n675 CS_BIAS.n518 161.3
R450 CS_BIAS.n674 CS_BIAS.n673 161.3
R451 CS_BIAS.n672 CS_BIAS.n519 161.3
R452 CS_BIAS.n671 CS_BIAS.n670 161.3
R453 CS_BIAS.n669 CS_BIAS.n520 161.3
R454 CS_BIAS.n668 CS_BIAS.n667 161.3
R455 CS_BIAS.n665 CS_BIAS.n521 161.3
R456 CS_BIAS.n664 CS_BIAS.n663 161.3
R457 CS_BIAS.n662 CS_BIAS.n522 161.3
R458 CS_BIAS.n661 CS_BIAS.n660 161.3
R459 CS_BIAS.n659 CS_BIAS.n523 161.3
R460 CS_BIAS.n658 CS_BIAS.n657 161.3
R461 CS_BIAS.n656 CS_BIAS.n524 161.3
R462 CS_BIAS.n655 CS_BIAS.n654 161.3
R463 CS_BIAS.n653 CS_BIAS.n525 161.3
R464 CS_BIAS.n652 CS_BIAS.n651 161.3
R465 CS_BIAS.n650 CS_BIAS.n526 161.3
R466 CS_BIAS.n649 CS_BIAS.n648 161.3
R467 CS_BIAS.n647 CS_BIAS.n527 161.3
R468 CS_BIAS.n555 CS_BIAS.t11 107.871
R469 CS_BIAS.n99 CS_BIAS.t15 106.037
R470 CS_BIAS.n103 CS_BIAS.n102 88.3741
R471 CS_BIAS.n101 CS_BIAS.n100 86.9991
R472 CS_BIAS.n641 CS_BIAS.n640 86.9991
R473 CS_BIAS.n555 CS_BIAS.n554 86.9991
R474 CS_BIAS.n512 CS_BIAS.n429 78.5377
R475 CS_BIAS.n427 CS_BIAS.n344 78.5377
R476 CS_BIAS.n342 CS_BIAS.n259 78.5377
R477 CS_BIAS.n257 CS_BIAS.n174 78.5377
R478 CS_BIAS.n98 CS_BIAS.n15 78.5377
R479 CS_BIAS.n173 CS_BIAS.n0 78.5377
R480 CS_BIAS.n1026 CS_BIAS.n943 78.5377
R481 CS_BIAS.n941 CS_BIAS.n858 78.5377
R482 CS_BIAS.n856 CS_BIAS.n773 78.5377
R483 CS_BIAS.n771 CS_BIAS.n688 78.5377
R484 CS_BIAS.n639 CS_BIAS.n556 78.5377
R485 CS_BIAS.n687 CS_BIAS.n514 78.5377
R486 CS_BIAS.n502 CS_BIAS.n433 73.0308
R487 CS_BIAS.n417 CS_BIAS.n348 73.0308
R488 CS_BIAS.n332 CS_BIAS.n263 73.0308
R489 CS_BIAS.n247 CS_BIAS.n178 73.0308
R490 CS_BIAS.n88 CS_BIAS.n19 73.0308
R491 CS_BIAS.n163 CS_BIAS.n4 73.0308
R492 CS_BIAS.n1016 CS_BIAS.n947 73.0308
R493 CS_BIAS.n931 CS_BIAS.n862 73.0308
R494 CS_BIAS.n846 CS_BIAS.n777 73.0308
R495 CS_BIAS.n761 CS_BIAS.n692 73.0308
R496 CS_BIAS.n629 CS_BIAS.n560 73.0308
R497 CS_BIAS.n677 CS_BIAS.n518 73.0308
R498 CS_BIAS.n450 CS_BIAS.n449 69.9188
R499 CS_BIAS.n365 CS_BIAS.n364 69.9188
R500 CS_BIAS.n280 CS_BIAS.n279 69.9188
R501 CS_BIAS.n195 CS_BIAS.n194 69.9188
R502 CS_BIAS.n36 CS_BIAS.n35 69.9188
R503 CS_BIAS.n111 CS_BIAS.n110 69.9188
R504 CS_BIAS.n964 CS_BIAS.n963 69.9188
R505 CS_BIAS.n879 CS_BIAS.n878 69.9188
R506 CS_BIAS.n794 CS_BIAS.n793 69.9188
R507 CS_BIAS.n709 CS_BIAS.n708 69.9188
R508 CS_BIAS.n577 CS_BIAS.n576 69.9188
R509 CS_BIAS.n535 CS_BIAS.n534 69.9188
R510 CS_BIAS.n460 CS_BIAS.n445 62.3743
R511 CS_BIAS.n479 CS_BIAS.n439 62.3743
R512 CS_BIAS.n394 CS_BIAS.n354 62.3743
R513 CS_BIAS.n375 CS_BIAS.n360 62.3743
R514 CS_BIAS.n309 CS_BIAS.n269 62.3743
R515 CS_BIAS.n290 CS_BIAS.n275 62.3743
R516 CS_BIAS.n224 CS_BIAS.n184 62.3743
R517 CS_BIAS.n205 CS_BIAS.n190 62.3743
R518 CS_BIAS.n65 CS_BIAS.n25 62.3743
R519 CS_BIAS.n46 CS_BIAS.n31 62.3743
R520 CS_BIAS.n140 CS_BIAS.n10 62.3743
R521 CS_BIAS.n121 CS_BIAS.n106 62.3743
R522 CS_BIAS.n974 CS_BIAS.n959 62.3743
R523 CS_BIAS.n993 CS_BIAS.n953 62.3743
R524 CS_BIAS.n889 CS_BIAS.n874 62.3743
R525 CS_BIAS.n908 CS_BIAS.n868 62.3743
R526 CS_BIAS.n804 CS_BIAS.n789 62.3743
R527 CS_BIAS.n823 CS_BIAS.n783 62.3743
R528 CS_BIAS.n719 CS_BIAS.n704 62.3743
R529 CS_BIAS.n738 CS_BIAS.n698 62.3743
R530 CS_BIAS.n587 CS_BIAS.n572 62.3743
R531 CS_BIAS.n606 CS_BIAS.n566 62.3743
R532 CS_BIAS.n654 CS_BIAS.n524 62.3743
R533 CS_BIAS.n545 CS_BIAS.n530 62.3743
R534 CS_BIAS.n460 CS_BIAS.n459 50.7491
R535 CS_BIAS.n483 CS_BIAS.n439 50.7491
R536 CS_BIAS.n398 CS_BIAS.n354 50.7491
R537 CS_BIAS.n375 CS_BIAS.n374 50.7491
R538 CS_BIAS.n313 CS_BIAS.n269 50.7491
R539 CS_BIAS.n290 CS_BIAS.n289 50.7491
R540 CS_BIAS.n228 CS_BIAS.n184 50.7491
R541 CS_BIAS.n205 CS_BIAS.n204 50.7491
R542 CS_BIAS.n69 CS_BIAS.n25 50.7491
R543 CS_BIAS.n46 CS_BIAS.n45 50.7491
R544 CS_BIAS.n144 CS_BIAS.n10 50.7491
R545 CS_BIAS.n121 CS_BIAS.n120 50.7491
R546 CS_BIAS.n974 CS_BIAS.n973 50.7491
R547 CS_BIAS.n997 CS_BIAS.n953 50.7491
R548 CS_BIAS.n889 CS_BIAS.n888 50.7491
R549 CS_BIAS.n912 CS_BIAS.n868 50.7491
R550 CS_BIAS.n804 CS_BIAS.n803 50.7491
R551 CS_BIAS.n827 CS_BIAS.n783 50.7491
R552 CS_BIAS.n719 CS_BIAS.n718 50.7491
R553 CS_BIAS.n742 CS_BIAS.n698 50.7491
R554 CS_BIAS.n587 CS_BIAS.n586 50.7491
R555 CS_BIAS.n610 CS_BIAS.n566 50.7491
R556 CS_BIAS.n658 CS_BIAS.n524 50.7491
R557 CS_BIAS.n545 CS_BIAS.n544 50.7491
R558 CS_BIAS.n964 CS_BIAS.t63 41.5421
R559 CS_BIAS.n879 CS_BIAS.t66 41.5421
R560 CS_BIAS.n794 CS_BIAS.t65 41.5421
R561 CS_BIAS.n709 CS_BIAS.t35 41.5421
R562 CS_BIAS.n577 CS_BIAS.t10 41.5421
R563 CS_BIAS.n535 CS_BIAS.t24 41.5421
R564 CS_BIAS.n450 CS_BIAS.t45 41.5421
R565 CS_BIAS.n365 CS_BIAS.t46 41.5421
R566 CS_BIAS.n280 CS_BIAS.t47 41.5421
R567 CS_BIAS.n195 CS_BIAS.t49 41.5421
R568 CS_BIAS.n36 CS_BIAS.t0 41.5421
R569 CS_BIAS.n111 CS_BIAS.t62 41.5421
R570 CS_BIAS.n503 CS_BIAS.n502 39.1239
R571 CS_BIAS.n418 CS_BIAS.n417 39.1239
R572 CS_BIAS.n333 CS_BIAS.n332 39.1239
R573 CS_BIAS.n248 CS_BIAS.n247 39.1239
R574 CS_BIAS.n89 CS_BIAS.n88 39.1239
R575 CS_BIAS.n164 CS_BIAS.n163 39.1239
R576 CS_BIAS.n1017 CS_BIAS.n1016 39.1239
R577 CS_BIAS.n932 CS_BIAS.n931 39.1239
R578 CS_BIAS.n847 CS_BIAS.n846 39.1239
R579 CS_BIAS.n762 CS_BIAS.n761 39.1239
R580 CS_BIAS.n630 CS_BIAS.n629 39.1239
R581 CS_BIAS.n678 CS_BIAS.n677 39.1239
R582 CS_BIAS.n498 CS_BIAS.n433 25.5611
R583 CS_BIAS.n413 CS_BIAS.n348 25.5611
R584 CS_BIAS.n328 CS_BIAS.n263 25.5611
R585 CS_BIAS.n243 CS_BIAS.n178 25.5611
R586 CS_BIAS.n84 CS_BIAS.n19 25.5611
R587 CS_BIAS.n159 CS_BIAS.n4 25.5611
R588 CS_BIAS.n1012 CS_BIAS.n947 25.5611
R589 CS_BIAS.n927 CS_BIAS.n862 25.5611
R590 CS_BIAS.n842 CS_BIAS.n777 25.5611
R591 CS_BIAS.n757 CS_BIAS.n692 25.5611
R592 CS_BIAS.n625 CS_BIAS.n560 25.5611
R593 CS_BIAS.n673 CS_BIAS.n518 25.5611
R594 CS_BIAS.n459 CS_BIAS.n458 24.5923
R595 CS_BIAS.n458 CS_BIAS.n447 24.5923
R596 CS_BIAS.n454 CS_BIAS.n447 24.5923
R597 CS_BIAS.n454 CS_BIAS.n453 24.5923
R598 CS_BIAS.n453 CS_BIAS.n452 24.5923
R599 CS_BIAS.n479 CS_BIAS.n478 24.5923
R600 CS_BIAS.n478 CS_BIAS.n477 24.5923
R601 CS_BIAS.n477 CS_BIAS.n441 24.5923
R602 CS_BIAS.n473 CS_BIAS.n441 24.5923
R603 CS_BIAS.n473 CS_BIAS.n472 24.5923
R604 CS_BIAS.n470 CS_BIAS.n443 24.5923
R605 CS_BIAS.n466 CS_BIAS.n443 24.5923
R606 CS_BIAS.n466 CS_BIAS.n465 24.5923
R607 CS_BIAS.n465 CS_BIAS.n464 24.5923
R608 CS_BIAS.n464 CS_BIAS.n445 24.5923
R609 CS_BIAS.n498 CS_BIAS.n497 24.5923
R610 CS_BIAS.n497 CS_BIAS.n496 24.5923
R611 CS_BIAS.n496 CS_BIAS.n435 24.5923
R612 CS_BIAS.n492 CS_BIAS.n435 24.5923
R613 CS_BIAS.n490 CS_BIAS.n489 24.5923
R614 CS_BIAS.n489 CS_BIAS.n437 24.5923
R615 CS_BIAS.n485 CS_BIAS.n437 24.5923
R616 CS_BIAS.n485 CS_BIAS.n484 24.5923
R617 CS_BIAS.n484 CS_BIAS.n483 24.5923
R618 CS_BIAS.n510 CS_BIAS.n509 24.5923
R619 CS_BIAS.n509 CS_BIAS.n508 24.5923
R620 CS_BIAS.n508 CS_BIAS.n431 24.5923
R621 CS_BIAS.n504 CS_BIAS.n431 24.5923
R622 CS_BIAS.n504 CS_BIAS.n503 24.5923
R623 CS_BIAS.n425 CS_BIAS.n424 24.5923
R624 CS_BIAS.n424 CS_BIAS.n423 24.5923
R625 CS_BIAS.n423 CS_BIAS.n346 24.5923
R626 CS_BIAS.n419 CS_BIAS.n346 24.5923
R627 CS_BIAS.n419 CS_BIAS.n418 24.5923
R628 CS_BIAS.n413 CS_BIAS.n412 24.5923
R629 CS_BIAS.n412 CS_BIAS.n411 24.5923
R630 CS_BIAS.n411 CS_BIAS.n350 24.5923
R631 CS_BIAS.n407 CS_BIAS.n350 24.5923
R632 CS_BIAS.n405 CS_BIAS.n404 24.5923
R633 CS_BIAS.n404 CS_BIAS.n352 24.5923
R634 CS_BIAS.n400 CS_BIAS.n352 24.5923
R635 CS_BIAS.n400 CS_BIAS.n399 24.5923
R636 CS_BIAS.n399 CS_BIAS.n398 24.5923
R637 CS_BIAS.n394 CS_BIAS.n393 24.5923
R638 CS_BIAS.n393 CS_BIAS.n392 24.5923
R639 CS_BIAS.n392 CS_BIAS.n356 24.5923
R640 CS_BIAS.n388 CS_BIAS.n356 24.5923
R641 CS_BIAS.n388 CS_BIAS.n387 24.5923
R642 CS_BIAS.n385 CS_BIAS.n358 24.5923
R643 CS_BIAS.n381 CS_BIAS.n358 24.5923
R644 CS_BIAS.n381 CS_BIAS.n380 24.5923
R645 CS_BIAS.n380 CS_BIAS.n379 24.5923
R646 CS_BIAS.n379 CS_BIAS.n360 24.5923
R647 CS_BIAS.n374 CS_BIAS.n373 24.5923
R648 CS_BIAS.n373 CS_BIAS.n362 24.5923
R649 CS_BIAS.n369 CS_BIAS.n362 24.5923
R650 CS_BIAS.n369 CS_BIAS.n368 24.5923
R651 CS_BIAS.n368 CS_BIAS.n367 24.5923
R652 CS_BIAS.n340 CS_BIAS.n339 24.5923
R653 CS_BIAS.n339 CS_BIAS.n338 24.5923
R654 CS_BIAS.n338 CS_BIAS.n261 24.5923
R655 CS_BIAS.n334 CS_BIAS.n261 24.5923
R656 CS_BIAS.n334 CS_BIAS.n333 24.5923
R657 CS_BIAS.n328 CS_BIAS.n327 24.5923
R658 CS_BIAS.n327 CS_BIAS.n326 24.5923
R659 CS_BIAS.n326 CS_BIAS.n265 24.5923
R660 CS_BIAS.n322 CS_BIAS.n265 24.5923
R661 CS_BIAS.n320 CS_BIAS.n319 24.5923
R662 CS_BIAS.n319 CS_BIAS.n267 24.5923
R663 CS_BIAS.n315 CS_BIAS.n267 24.5923
R664 CS_BIAS.n315 CS_BIAS.n314 24.5923
R665 CS_BIAS.n314 CS_BIAS.n313 24.5923
R666 CS_BIAS.n309 CS_BIAS.n308 24.5923
R667 CS_BIAS.n308 CS_BIAS.n307 24.5923
R668 CS_BIAS.n307 CS_BIAS.n271 24.5923
R669 CS_BIAS.n303 CS_BIAS.n271 24.5923
R670 CS_BIAS.n303 CS_BIAS.n302 24.5923
R671 CS_BIAS.n300 CS_BIAS.n273 24.5923
R672 CS_BIAS.n296 CS_BIAS.n273 24.5923
R673 CS_BIAS.n296 CS_BIAS.n295 24.5923
R674 CS_BIAS.n295 CS_BIAS.n294 24.5923
R675 CS_BIAS.n294 CS_BIAS.n275 24.5923
R676 CS_BIAS.n289 CS_BIAS.n288 24.5923
R677 CS_BIAS.n288 CS_BIAS.n277 24.5923
R678 CS_BIAS.n284 CS_BIAS.n277 24.5923
R679 CS_BIAS.n284 CS_BIAS.n283 24.5923
R680 CS_BIAS.n283 CS_BIAS.n282 24.5923
R681 CS_BIAS.n255 CS_BIAS.n254 24.5923
R682 CS_BIAS.n254 CS_BIAS.n253 24.5923
R683 CS_BIAS.n253 CS_BIAS.n176 24.5923
R684 CS_BIAS.n249 CS_BIAS.n176 24.5923
R685 CS_BIAS.n249 CS_BIAS.n248 24.5923
R686 CS_BIAS.n243 CS_BIAS.n242 24.5923
R687 CS_BIAS.n242 CS_BIAS.n241 24.5923
R688 CS_BIAS.n241 CS_BIAS.n180 24.5923
R689 CS_BIAS.n237 CS_BIAS.n180 24.5923
R690 CS_BIAS.n235 CS_BIAS.n234 24.5923
R691 CS_BIAS.n234 CS_BIAS.n182 24.5923
R692 CS_BIAS.n230 CS_BIAS.n182 24.5923
R693 CS_BIAS.n230 CS_BIAS.n229 24.5923
R694 CS_BIAS.n229 CS_BIAS.n228 24.5923
R695 CS_BIAS.n224 CS_BIAS.n223 24.5923
R696 CS_BIAS.n223 CS_BIAS.n222 24.5923
R697 CS_BIAS.n222 CS_BIAS.n186 24.5923
R698 CS_BIAS.n218 CS_BIAS.n186 24.5923
R699 CS_BIAS.n218 CS_BIAS.n217 24.5923
R700 CS_BIAS.n215 CS_BIAS.n188 24.5923
R701 CS_BIAS.n211 CS_BIAS.n188 24.5923
R702 CS_BIAS.n211 CS_BIAS.n210 24.5923
R703 CS_BIAS.n210 CS_BIAS.n209 24.5923
R704 CS_BIAS.n209 CS_BIAS.n190 24.5923
R705 CS_BIAS.n204 CS_BIAS.n203 24.5923
R706 CS_BIAS.n203 CS_BIAS.n192 24.5923
R707 CS_BIAS.n199 CS_BIAS.n192 24.5923
R708 CS_BIAS.n199 CS_BIAS.n198 24.5923
R709 CS_BIAS.n198 CS_BIAS.n197 24.5923
R710 CS_BIAS.n96 CS_BIAS.n95 24.5923
R711 CS_BIAS.n95 CS_BIAS.n94 24.5923
R712 CS_BIAS.n94 CS_BIAS.n17 24.5923
R713 CS_BIAS.n90 CS_BIAS.n17 24.5923
R714 CS_BIAS.n90 CS_BIAS.n89 24.5923
R715 CS_BIAS.n84 CS_BIAS.n83 24.5923
R716 CS_BIAS.n83 CS_BIAS.n82 24.5923
R717 CS_BIAS.n82 CS_BIAS.n21 24.5923
R718 CS_BIAS.n78 CS_BIAS.n21 24.5923
R719 CS_BIAS.n76 CS_BIAS.n75 24.5923
R720 CS_BIAS.n75 CS_BIAS.n23 24.5923
R721 CS_BIAS.n71 CS_BIAS.n23 24.5923
R722 CS_BIAS.n71 CS_BIAS.n70 24.5923
R723 CS_BIAS.n70 CS_BIAS.n69 24.5923
R724 CS_BIAS.n65 CS_BIAS.n64 24.5923
R725 CS_BIAS.n64 CS_BIAS.n63 24.5923
R726 CS_BIAS.n63 CS_BIAS.n27 24.5923
R727 CS_BIAS.n59 CS_BIAS.n27 24.5923
R728 CS_BIAS.n59 CS_BIAS.n58 24.5923
R729 CS_BIAS.n56 CS_BIAS.n29 24.5923
R730 CS_BIAS.n52 CS_BIAS.n29 24.5923
R731 CS_BIAS.n52 CS_BIAS.n51 24.5923
R732 CS_BIAS.n51 CS_BIAS.n50 24.5923
R733 CS_BIAS.n50 CS_BIAS.n31 24.5923
R734 CS_BIAS.n45 CS_BIAS.n44 24.5923
R735 CS_BIAS.n44 CS_BIAS.n33 24.5923
R736 CS_BIAS.n40 CS_BIAS.n33 24.5923
R737 CS_BIAS.n40 CS_BIAS.n39 24.5923
R738 CS_BIAS.n39 CS_BIAS.n38 24.5923
R739 CS_BIAS.n171 CS_BIAS.n170 24.5923
R740 CS_BIAS.n170 CS_BIAS.n169 24.5923
R741 CS_BIAS.n169 CS_BIAS.n2 24.5923
R742 CS_BIAS.n165 CS_BIAS.n2 24.5923
R743 CS_BIAS.n165 CS_BIAS.n164 24.5923
R744 CS_BIAS.n159 CS_BIAS.n158 24.5923
R745 CS_BIAS.n158 CS_BIAS.n157 24.5923
R746 CS_BIAS.n157 CS_BIAS.n6 24.5923
R747 CS_BIAS.n153 CS_BIAS.n6 24.5923
R748 CS_BIAS.n151 CS_BIAS.n150 24.5923
R749 CS_BIAS.n150 CS_BIAS.n8 24.5923
R750 CS_BIAS.n146 CS_BIAS.n8 24.5923
R751 CS_BIAS.n146 CS_BIAS.n145 24.5923
R752 CS_BIAS.n145 CS_BIAS.n144 24.5923
R753 CS_BIAS.n140 CS_BIAS.n139 24.5923
R754 CS_BIAS.n139 CS_BIAS.n138 24.5923
R755 CS_BIAS.n138 CS_BIAS.n12 24.5923
R756 CS_BIAS.n134 CS_BIAS.n12 24.5923
R757 CS_BIAS.n134 CS_BIAS.n133 24.5923
R758 CS_BIAS.n131 CS_BIAS.n14 24.5923
R759 CS_BIAS.n127 CS_BIAS.n14 24.5923
R760 CS_BIAS.n127 CS_BIAS.n126 24.5923
R761 CS_BIAS.n126 CS_BIAS.n125 24.5923
R762 CS_BIAS.n125 CS_BIAS.n106 24.5923
R763 CS_BIAS.n120 CS_BIAS.n119 24.5923
R764 CS_BIAS.n119 CS_BIAS.n108 24.5923
R765 CS_BIAS.n115 CS_BIAS.n108 24.5923
R766 CS_BIAS.n115 CS_BIAS.n114 24.5923
R767 CS_BIAS.n114 CS_BIAS.n113 24.5923
R768 CS_BIAS.n967 CS_BIAS.n966 24.5923
R769 CS_BIAS.n968 CS_BIAS.n967 24.5923
R770 CS_BIAS.n968 CS_BIAS.n961 24.5923
R771 CS_BIAS.n972 CS_BIAS.n961 24.5923
R772 CS_BIAS.n973 CS_BIAS.n972 24.5923
R773 CS_BIAS.n978 CS_BIAS.n959 24.5923
R774 CS_BIAS.n979 CS_BIAS.n978 24.5923
R775 CS_BIAS.n980 CS_BIAS.n979 24.5923
R776 CS_BIAS.n980 CS_BIAS.n957 24.5923
R777 CS_BIAS.n984 CS_BIAS.n957 24.5923
R778 CS_BIAS.n987 CS_BIAS.n986 24.5923
R779 CS_BIAS.n987 CS_BIAS.n955 24.5923
R780 CS_BIAS.n991 CS_BIAS.n955 24.5923
R781 CS_BIAS.n992 CS_BIAS.n991 24.5923
R782 CS_BIAS.n993 CS_BIAS.n992 24.5923
R783 CS_BIAS.n998 CS_BIAS.n997 24.5923
R784 CS_BIAS.n999 CS_BIAS.n998 24.5923
R785 CS_BIAS.n999 CS_BIAS.n951 24.5923
R786 CS_BIAS.n1003 CS_BIAS.n951 24.5923
R787 CS_BIAS.n1004 CS_BIAS.n1003 24.5923
R788 CS_BIAS.n1006 CS_BIAS.n949 24.5923
R789 CS_BIAS.n1010 CS_BIAS.n949 24.5923
R790 CS_BIAS.n1011 CS_BIAS.n1010 24.5923
R791 CS_BIAS.n1012 CS_BIAS.n1011 24.5923
R792 CS_BIAS.n1018 CS_BIAS.n1017 24.5923
R793 CS_BIAS.n1018 CS_BIAS.n945 24.5923
R794 CS_BIAS.n1022 CS_BIAS.n945 24.5923
R795 CS_BIAS.n1023 CS_BIAS.n1022 24.5923
R796 CS_BIAS.n1024 CS_BIAS.n1023 24.5923
R797 CS_BIAS.n882 CS_BIAS.n881 24.5923
R798 CS_BIAS.n883 CS_BIAS.n882 24.5923
R799 CS_BIAS.n883 CS_BIAS.n876 24.5923
R800 CS_BIAS.n887 CS_BIAS.n876 24.5923
R801 CS_BIAS.n888 CS_BIAS.n887 24.5923
R802 CS_BIAS.n893 CS_BIAS.n874 24.5923
R803 CS_BIAS.n894 CS_BIAS.n893 24.5923
R804 CS_BIAS.n895 CS_BIAS.n894 24.5923
R805 CS_BIAS.n895 CS_BIAS.n872 24.5923
R806 CS_BIAS.n899 CS_BIAS.n872 24.5923
R807 CS_BIAS.n902 CS_BIAS.n901 24.5923
R808 CS_BIAS.n902 CS_BIAS.n870 24.5923
R809 CS_BIAS.n906 CS_BIAS.n870 24.5923
R810 CS_BIAS.n907 CS_BIAS.n906 24.5923
R811 CS_BIAS.n908 CS_BIAS.n907 24.5923
R812 CS_BIAS.n913 CS_BIAS.n912 24.5923
R813 CS_BIAS.n914 CS_BIAS.n913 24.5923
R814 CS_BIAS.n914 CS_BIAS.n866 24.5923
R815 CS_BIAS.n918 CS_BIAS.n866 24.5923
R816 CS_BIAS.n919 CS_BIAS.n918 24.5923
R817 CS_BIAS.n921 CS_BIAS.n864 24.5923
R818 CS_BIAS.n925 CS_BIAS.n864 24.5923
R819 CS_BIAS.n926 CS_BIAS.n925 24.5923
R820 CS_BIAS.n927 CS_BIAS.n926 24.5923
R821 CS_BIAS.n933 CS_BIAS.n932 24.5923
R822 CS_BIAS.n933 CS_BIAS.n860 24.5923
R823 CS_BIAS.n937 CS_BIAS.n860 24.5923
R824 CS_BIAS.n938 CS_BIAS.n937 24.5923
R825 CS_BIAS.n939 CS_BIAS.n938 24.5923
R826 CS_BIAS.n797 CS_BIAS.n796 24.5923
R827 CS_BIAS.n798 CS_BIAS.n797 24.5923
R828 CS_BIAS.n798 CS_BIAS.n791 24.5923
R829 CS_BIAS.n802 CS_BIAS.n791 24.5923
R830 CS_BIAS.n803 CS_BIAS.n802 24.5923
R831 CS_BIAS.n808 CS_BIAS.n789 24.5923
R832 CS_BIAS.n809 CS_BIAS.n808 24.5923
R833 CS_BIAS.n810 CS_BIAS.n809 24.5923
R834 CS_BIAS.n810 CS_BIAS.n787 24.5923
R835 CS_BIAS.n814 CS_BIAS.n787 24.5923
R836 CS_BIAS.n817 CS_BIAS.n816 24.5923
R837 CS_BIAS.n817 CS_BIAS.n785 24.5923
R838 CS_BIAS.n821 CS_BIAS.n785 24.5923
R839 CS_BIAS.n822 CS_BIAS.n821 24.5923
R840 CS_BIAS.n823 CS_BIAS.n822 24.5923
R841 CS_BIAS.n828 CS_BIAS.n827 24.5923
R842 CS_BIAS.n829 CS_BIAS.n828 24.5923
R843 CS_BIAS.n829 CS_BIAS.n781 24.5923
R844 CS_BIAS.n833 CS_BIAS.n781 24.5923
R845 CS_BIAS.n834 CS_BIAS.n833 24.5923
R846 CS_BIAS.n836 CS_BIAS.n779 24.5923
R847 CS_BIAS.n840 CS_BIAS.n779 24.5923
R848 CS_BIAS.n841 CS_BIAS.n840 24.5923
R849 CS_BIAS.n842 CS_BIAS.n841 24.5923
R850 CS_BIAS.n848 CS_BIAS.n847 24.5923
R851 CS_BIAS.n848 CS_BIAS.n775 24.5923
R852 CS_BIAS.n852 CS_BIAS.n775 24.5923
R853 CS_BIAS.n853 CS_BIAS.n852 24.5923
R854 CS_BIAS.n854 CS_BIAS.n853 24.5923
R855 CS_BIAS.n712 CS_BIAS.n711 24.5923
R856 CS_BIAS.n713 CS_BIAS.n712 24.5923
R857 CS_BIAS.n713 CS_BIAS.n706 24.5923
R858 CS_BIAS.n717 CS_BIAS.n706 24.5923
R859 CS_BIAS.n718 CS_BIAS.n717 24.5923
R860 CS_BIAS.n723 CS_BIAS.n704 24.5923
R861 CS_BIAS.n724 CS_BIAS.n723 24.5923
R862 CS_BIAS.n725 CS_BIAS.n724 24.5923
R863 CS_BIAS.n725 CS_BIAS.n702 24.5923
R864 CS_BIAS.n729 CS_BIAS.n702 24.5923
R865 CS_BIAS.n732 CS_BIAS.n731 24.5923
R866 CS_BIAS.n732 CS_BIAS.n700 24.5923
R867 CS_BIAS.n736 CS_BIAS.n700 24.5923
R868 CS_BIAS.n737 CS_BIAS.n736 24.5923
R869 CS_BIAS.n738 CS_BIAS.n737 24.5923
R870 CS_BIAS.n743 CS_BIAS.n742 24.5923
R871 CS_BIAS.n744 CS_BIAS.n743 24.5923
R872 CS_BIAS.n744 CS_BIAS.n696 24.5923
R873 CS_BIAS.n748 CS_BIAS.n696 24.5923
R874 CS_BIAS.n749 CS_BIAS.n748 24.5923
R875 CS_BIAS.n751 CS_BIAS.n694 24.5923
R876 CS_BIAS.n755 CS_BIAS.n694 24.5923
R877 CS_BIAS.n756 CS_BIAS.n755 24.5923
R878 CS_BIAS.n757 CS_BIAS.n756 24.5923
R879 CS_BIAS.n763 CS_BIAS.n762 24.5923
R880 CS_BIAS.n763 CS_BIAS.n690 24.5923
R881 CS_BIAS.n767 CS_BIAS.n690 24.5923
R882 CS_BIAS.n768 CS_BIAS.n767 24.5923
R883 CS_BIAS.n769 CS_BIAS.n768 24.5923
R884 CS_BIAS.n580 CS_BIAS.n579 24.5923
R885 CS_BIAS.n581 CS_BIAS.n580 24.5923
R886 CS_BIAS.n581 CS_BIAS.n574 24.5923
R887 CS_BIAS.n585 CS_BIAS.n574 24.5923
R888 CS_BIAS.n586 CS_BIAS.n585 24.5923
R889 CS_BIAS.n591 CS_BIAS.n572 24.5923
R890 CS_BIAS.n592 CS_BIAS.n591 24.5923
R891 CS_BIAS.n593 CS_BIAS.n592 24.5923
R892 CS_BIAS.n593 CS_BIAS.n570 24.5923
R893 CS_BIAS.n597 CS_BIAS.n570 24.5923
R894 CS_BIAS.n600 CS_BIAS.n599 24.5923
R895 CS_BIAS.n600 CS_BIAS.n568 24.5923
R896 CS_BIAS.n604 CS_BIAS.n568 24.5923
R897 CS_BIAS.n605 CS_BIAS.n604 24.5923
R898 CS_BIAS.n606 CS_BIAS.n605 24.5923
R899 CS_BIAS.n611 CS_BIAS.n610 24.5923
R900 CS_BIAS.n612 CS_BIAS.n611 24.5923
R901 CS_BIAS.n612 CS_BIAS.n564 24.5923
R902 CS_BIAS.n616 CS_BIAS.n564 24.5923
R903 CS_BIAS.n617 CS_BIAS.n616 24.5923
R904 CS_BIAS.n619 CS_BIAS.n562 24.5923
R905 CS_BIAS.n623 CS_BIAS.n562 24.5923
R906 CS_BIAS.n624 CS_BIAS.n623 24.5923
R907 CS_BIAS.n625 CS_BIAS.n624 24.5923
R908 CS_BIAS.n631 CS_BIAS.n630 24.5923
R909 CS_BIAS.n631 CS_BIAS.n558 24.5923
R910 CS_BIAS.n635 CS_BIAS.n558 24.5923
R911 CS_BIAS.n636 CS_BIAS.n635 24.5923
R912 CS_BIAS.n637 CS_BIAS.n636 24.5923
R913 CS_BIAS.n679 CS_BIAS.n678 24.5923
R914 CS_BIAS.n679 CS_BIAS.n516 24.5923
R915 CS_BIAS.n683 CS_BIAS.n516 24.5923
R916 CS_BIAS.n684 CS_BIAS.n683 24.5923
R917 CS_BIAS.n685 CS_BIAS.n684 24.5923
R918 CS_BIAS.n659 CS_BIAS.n658 24.5923
R919 CS_BIAS.n660 CS_BIAS.n659 24.5923
R920 CS_BIAS.n660 CS_BIAS.n522 24.5923
R921 CS_BIAS.n664 CS_BIAS.n522 24.5923
R922 CS_BIAS.n665 CS_BIAS.n664 24.5923
R923 CS_BIAS.n667 CS_BIAS.n520 24.5923
R924 CS_BIAS.n671 CS_BIAS.n520 24.5923
R925 CS_BIAS.n672 CS_BIAS.n671 24.5923
R926 CS_BIAS.n673 CS_BIAS.n672 24.5923
R927 CS_BIAS.n538 CS_BIAS.n537 24.5923
R928 CS_BIAS.n539 CS_BIAS.n538 24.5923
R929 CS_BIAS.n539 CS_BIAS.n532 24.5923
R930 CS_BIAS.n543 CS_BIAS.n532 24.5923
R931 CS_BIAS.n544 CS_BIAS.n543 24.5923
R932 CS_BIAS.n549 CS_BIAS.n530 24.5923
R933 CS_BIAS.n550 CS_BIAS.n549 24.5923
R934 CS_BIAS.n551 CS_BIAS.n550 24.5923
R935 CS_BIAS.n551 CS_BIAS.n528 24.5923
R936 CS_BIAS.n645 CS_BIAS.n528 24.5923
R937 CS_BIAS.n648 CS_BIAS.n647 24.5923
R938 CS_BIAS.n648 CS_BIAS.n526 24.5923
R939 CS_BIAS.n652 CS_BIAS.n526 24.5923
R940 CS_BIAS.n653 CS_BIAS.n652 24.5923
R941 CS_BIAS.n654 CS_BIAS.n653 24.5923
R942 CS_BIAS.n102 CS_BIAS.t17 19.039
R943 CS_BIAS.n102 CS_BIAS.t1 19.039
R944 CS_BIAS.n100 CS_BIAS.t19 19.039
R945 CS_BIAS.n100 CS_BIAS.t3 19.039
R946 CS_BIAS.n640 CS_BIAS.t9 19.039
R947 CS_BIAS.n640 CS_BIAS.t5 19.039
R948 CS_BIAS.n554 CS_BIAS.t13 19.039
R949 CS_BIAS.n554 CS_BIAS.t7 19.039
R950 CS_BIAS.n492 CS_BIAS.n491 18.1985
R951 CS_BIAS.n407 CS_BIAS.n406 18.1985
R952 CS_BIAS.n322 CS_BIAS.n321 18.1985
R953 CS_BIAS.n237 CS_BIAS.n236 18.1985
R954 CS_BIAS.n78 CS_BIAS.n77 18.1985
R955 CS_BIAS.n153 CS_BIAS.n152 18.1985
R956 CS_BIAS.n1006 CS_BIAS.n1005 18.1985
R957 CS_BIAS.n921 CS_BIAS.n920 18.1985
R958 CS_BIAS.n836 CS_BIAS.n835 18.1985
R959 CS_BIAS.n751 CS_BIAS.n750 18.1985
R960 CS_BIAS.n619 CS_BIAS.n618 18.1985
R961 CS_BIAS.n667 CS_BIAS.n666 18.1985
R962 CS_BIAS.n641 CS_BIAS.n639 12.3394
R963 CS_BIAS.n472 CS_BIAS.n471 12.2964
R964 CS_BIAS.n471 CS_BIAS.n470 12.2964
R965 CS_BIAS.n387 CS_BIAS.n386 12.2964
R966 CS_BIAS.n386 CS_BIAS.n385 12.2964
R967 CS_BIAS.n302 CS_BIAS.n301 12.2964
R968 CS_BIAS.n301 CS_BIAS.n300 12.2964
R969 CS_BIAS.n217 CS_BIAS.n216 12.2964
R970 CS_BIAS.n216 CS_BIAS.n215 12.2964
R971 CS_BIAS.n58 CS_BIAS.n57 12.2964
R972 CS_BIAS.n57 CS_BIAS.n56 12.2964
R973 CS_BIAS.n133 CS_BIAS.n132 12.2964
R974 CS_BIAS.n132 CS_BIAS.n131 12.2964
R975 CS_BIAS.n985 CS_BIAS.n984 12.2964
R976 CS_BIAS.n986 CS_BIAS.n985 12.2964
R977 CS_BIAS.n900 CS_BIAS.n899 12.2964
R978 CS_BIAS.n901 CS_BIAS.n900 12.2964
R979 CS_BIAS.n815 CS_BIAS.n814 12.2964
R980 CS_BIAS.n816 CS_BIAS.n815 12.2964
R981 CS_BIAS.n730 CS_BIAS.n729 12.2964
R982 CS_BIAS.n731 CS_BIAS.n730 12.2964
R983 CS_BIAS.n598 CS_BIAS.n597 12.2964
R984 CS_BIAS.n599 CS_BIAS.n598 12.2964
R985 CS_BIAS.n646 CS_BIAS.n645 12.2964
R986 CS_BIAS.n647 CS_BIAS.n646 12.2964
R987 CS_BIAS.n99 CS_BIAS.n98 11.4227
R988 CS_BIAS.n1028 CS_BIAS.n513 9.83298
R989 CS_BIAS.n104 CS_BIAS.n103 9.50363
R990 CS_BIAS.n643 CS_BIAS.n642 9.50363
R991 CS_BIAS.n449 CS_BIAS.t51 8.76414
R992 CS_BIAS.n471 CS_BIAS.t26 8.76414
R993 CS_BIAS.n491 CS_BIAS.t36 8.76414
R994 CS_BIAS.n429 CS_BIAS.t67 8.76414
R995 CS_BIAS.n344 CS_BIAS.t68 8.76414
R996 CS_BIAS.n406 CS_BIAS.t38 8.76414
R997 CS_BIAS.n386 CS_BIAS.t29 8.76414
R998 CS_BIAS.n364 CS_BIAS.t52 8.76414
R999 CS_BIAS.n259 CS_BIAS.t69 8.76414
R1000 CS_BIAS.n321 CS_BIAS.t39 8.76414
R1001 CS_BIAS.n301 CS_BIAS.t30 8.76414
R1002 CS_BIAS.n279 CS_BIAS.t53 8.76414
R1003 CS_BIAS.n174 CS_BIAS.t42 8.76414
R1004 CS_BIAS.n236 CS_BIAS.t48 8.76414
R1005 CS_BIAS.n216 CS_BIAS.t32 8.76414
R1006 CS_BIAS.n194 CS_BIAS.t61 8.76414
R1007 CS_BIAS.n15 CS_BIAS.t14 8.76414
R1008 CS_BIAS.n77 CS_BIAS.t18 8.76414
R1009 CS_BIAS.n57 CS_BIAS.t2 8.76414
R1010 CS_BIAS.n35 CS_BIAS.t16 8.76414
R1011 CS_BIAS.n0 CS_BIAS.t50 8.76414
R1012 CS_BIAS.n152 CS_BIAS.t43 8.76414
R1013 CS_BIAS.n132 CS_BIAS.t58 8.76414
R1014 CS_BIAS.n110 CS_BIAS.t44 8.76414
R1015 CS_BIAS.n963 CS_BIAS.t57 8.76414
R1016 CS_BIAS.n985 CS_BIAS.t21 8.76414
R1017 CS_BIAS.n1005 CS_BIAS.t28 8.76414
R1018 CS_BIAS.n943 CS_BIAS.t37 8.76414
R1019 CS_BIAS.n878 CS_BIAS.t59 8.76414
R1020 CS_BIAS.n900 CS_BIAS.t20 8.76414
R1021 CS_BIAS.n920 CS_BIAS.t27 8.76414
R1022 CS_BIAS.n858 CS_BIAS.t41 8.76414
R1023 CS_BIAS.n793 CS_BIAS.t60 8.76414
R1024 CS_BIAS.n815 CS_BIAS.t22 8.76414
R1025 CS_BIAS.n835 CS_BIAS.t31 8.76414
R1026 CS_BIAS.n773 CS_BIAS.t40 8.76414
R1027 CS_BIAS.n708 CS_BIAS.t64 8.76414
R1028 CS_BIAS.n730 CS_BIAS.t34 8.76414
R1029 CS_BIAS.n750 CS_BIAS.t56 8.76414
R1030 CS_BIAS.n688 CS_BIAS.t25 8.76414
R1031 CS_BIAS.n576 CS_BIAS.t12 8.76414
R1032 CS_BIAS.n598 CS_BIAS.t6 8.76414
R1033 CS_BIAS.n618 CS_BIAS.t8 8.76414
R1034 CS_BIAS.n556 CS_BIAS.t4 8.76414
R1035 CS_BIAS.n514 CS_BIAS.t55 8.76414
R1036 CS_BIAS.n666 CS_BIAS.t33 8.76414
R1037 CS_BIAS.n534 CS_BIAS.t23 8.76414
R1038 CS_BIAS.n646 CS_BIAS.t54 8.76414
R1039 CS_BIAS.n258 CS_BIAS.n173 7.46183
R1040 CS_BIAS.n772 CS_BIAS.n687 7.46183
R1041 CS_BIAS.n452 CS_BIAS.n449 6.39438
R1042 CS_BIAS.n491 CS_BIAS.n490 6.39438
R1043 CS_BIAS.n406 CS_BIAS.n405 6.39438
R1044 CS_BIAS.n367 CS_BIAS.n364 6.39438
R1045 CS_BIAS.n321 CS_BIAS.n320 6.39438
R1046 CS_BIAS.n282 CS_BIAS.n279 6.39438
R1047 CS_BIAS.n236 CS_BIAS.n235 6.39438
R1048 CS_BIAS.n197 CS_BIAS.n194 6.39438
R1049 CS_BIAS.n77 CS_BIAS.n76 6.39438
R1050 CS_BIAS.n38 CS_BIAS.n35 6.39438
R1051 CS_BIAS.n152 CS_BIAS.n151 6.39438
R1052 CS_BIAS.n113 CS_BIAS.n110 6.39438
R1053 CS_BIAS.n966 CS_BIAS.n963 6.39438
R1054 CS_BIAS.n1005 CS_BIAS.n1004 6.39438
R1055 CS_BIAS.n881 CS_BIAS.n878 6.39438
R1056 CS_BIAS.n920 CS_BIAS.n919 6.39438
R1057 CS_BIAS.n796 CS_BIAS.n793 6.39438
R1058 CS_BIAS.n835 CS_BIAS.n834 6.39438
R1059 CS_BIAS.n711 CS_BIAS.n708 6.39438
R1060 CS_BIAS.n750 CS_BIAS.n749 6.39438
R1061 CS_BIAS.n579 CS_BIAS.n576 6.39438
R1062 CS_BIAS.n618 CS_BIAS.n617 6.39438
R1063 CS_BIAS.n666 CS_BIAS.n665 6.39438
R1064 CS_BIAS.n537 CS_BIAS.n534 6.39438
R1065 CS_BIAS.n1028 CS_BIAS.n1027 6.18891
R1066 CS_BIAS.n513 CS_BIAS.n512 5.41448
R1067 CS_BIAS.n428 CS_BIAS.n427 5.41448
R1068 CS_BIAS.n343 CS_BIAS.n342 5.41448
R1069 CS_BIAS.n258 CS_BIAS.n257 5.41448
R1070 CS_BIAS.n1027 CS_BIAS.n1026 5.41448
R1071 CS_BIAS.n942 CS_BIAS.n941 5.41448
R1072 CS_BIAS.n857 CS_BIAS.n856 5.41448
R1073 CS_BIAS.n772 CS_BIAS.n771 5.41448
R1074 CS_BIAS CS_BIAS.n1028 4.37075
R1075 CS_BIAS.n343 CS_BIAS.n258 2.04785
R1076 CS_BIAS.n428 CS_BIAS.n343 2.04785
R1077 CS_BIAS.n513 CS_BIAS.n428 2.04785
R1078 CS_BIAS.n857 CS_BIAS.n772 2.04785
R1079 CS_BIAS.n942 CS_BIAS.n857 2.04785
R1080 CS_BIAS.n1027 CS_BIAS.n942 2.04785
R1081 CS_BIAS.n101 CS_BIAS.n99 1.83383
R1082 CS_BIAS.n642 CS_BIAS.n641 1.3755
R1083 CS_BIAS.n965 CS_BIAS.n964 0.881314
R1084 CS_BIAS.n880 CS_BIAS.n879 0.881314
R1085 CS_BIAS.n795 CS_BIAS.n794 0.881314
R1086 CS_BIAS.n710 CS_BIAS.n709 0.881314
R1087 CS_BIAS.n578 CS_BIAS.n577 0.881314
R1088 CS_BIAS.n536 CS_BIAS.n535 0.881314
R1089 CS_BIAS.n451 CS_BIAS.n450 0.881314
R1090 CS_BIAS.n366 CS_BIAS.n365 0.881313
R1091 CS_BIAS.n281 CS_BIAS.n280 0.881313
R1092 CS_BIAS.n196 CS_BIAS.n195 0.881313
R1093 CS_BIAS.n37 CS_BIAS.n36 0.881313
R1094 CS_BIAS.n112 CS_BIAS.n111 0.881313
R1095 CS_BIAS.n510 CS_BIAS.n429 0.492337
R1096 CS_BIAS.n425 CS_BIAS.n344 0.492337
R1097 CS_BIAS.n340 CS_BIAS.n259 0.492337
R1098 CS_BIAS.n255 CS_BIAS.n174 0.492337
R1099 CS_BIAS.n96 CS_BIAS.n15 0.492337
R1100 CS_BIAS.n171 CS_BIAS.n0 0.492337
R1101 CS_BIAS.n1024 CS_BIAS.n943 0.492337
R1102 CS_BIAS.n939 CS_BIAS.n858 0.492337
R1103 CS_BIAS.n854 CS_BIAS.n773 0.492337
R1104 CS_BIAS.n769 CS_BIAS.n688 0.492337
R1105 CS_BIAS.n637 CS_BIAS.n556 0.492337
R1106 CS_BIAS.n685 CS_BIAS.n514 0.492337
R1107 CS_BIAS.n512 CS_BIAS.n511 0.46582
R1108 CS_BIAS.n427 CS_BIAS.n426 0.46582
R1109 CS_BIAS.n342 CS_BIAS.n341 0.46582
R1110 CS_BIAS.n257 CS_BIAS.n256 0.46582
R1111 CS_BIAS.n98 CS_BIAS.n97 0.46582
R1112 CS_BIAS.n173 CS_BIAS.n172 0.46582
R1113 CS_BIAS.n1026 CS_BIAS.n1025 0.46582
R1114 CS_BIAS.n941 CS_BIAS.n940 0.46582
R1115 CS_BIAS.n856 CS_BIAS.n855 0.46582
R1116 CS_BIAS.n771 CS_BIAS.n770 0.46582
R1117 CS_BIAS.n639 CS_BIAS.n638 0.46582
R1118 CS_BIAS.n687 CS_BIAS.n686 0.46582
R1119 CS_BIAS.n103 CS_BIAS.n101 0.458833
R1120 CS_BIAS.n642 CS_BIAS.n555 0.458833
R1121 CS_BIAS.n511 CS_BIAS.n430 0.189894
R1122 CS_BIAS.n507 CS_BIAS.n430 0.189894
R1123 CS_BIAS.n507 CS_BIAS.n506 0.189894
R1124 CS_BIAS.n506 CS_BIAS.n505 0.189894
R1125 CS_BIAS.n505 CS_BIAS.n432 0.189894
R1126 CS_BIAS.n501 CS_BIAS.n432 0.189894
R1127 CS_BIAS.n501 CS_BIAS.n500 0.189894
R1128 CS_BIAS.n500 CS_BIAS.n499 0.189894
R1129 CS_BIAS.n499 CS_BIAS.n434 0.189894
R1130 CS_BIAS.n495 CS_BIAS.n434 0.189894
R1131 CS_BIAS.n495 CS_BIAS.n494 0.189894
R1132 CS_BIAS.n494 CS_BIAS.n493 0.189894
R1133 CS_BIAS.n493 CS_BIAS.n436 0.189894
R1134 CS_BIAS.n488 CS_BIAS.n436 0.189894
R1135 CS_BIAS.n488 CS_BIAS.n487 0.189894
R1136 CS_BIAS.n487 CS_BIAS.n486 0.189894
R1137 CS_BIAS.n486 CS_BIAS.n438 0.189894
R1138 CS_BIAS.n482 CS_BIAS.n438 0.189894
R1139 CS_BIAS.n482 CS_BIAS.n481 0.189894
R1140 CS_BIAS.n481 CS_BIAS.n480 0.189894
R1141 CS_BIAS.n480 CS_BIAS.n440 0.189894
R1142 CS_BIAS.n476 CS_BIAS.n440 0.189894
R1143 CS_BIAS.n476 CS_BIAS.n475 0.189894
R1144 CS_BIAS.n475 CS_BIAS.n474 0.189894
R1145 CS_BIAS.n474 CS_BIAS.n442 0.189894
R1146 CS_BIAS.n469 CS_BIAS.n442 0.189894
R1147 CS_BIAS.n469 CS_BIAS.n468 0.189894
R1148 CS_BIAS.n468 CS_BIAS.n467 0.189894
R1149 CS_BIAS.n467 CS_BIAS.n444 0.189894
R1150 CS_BIAS.n463 CS_BIAS.n444 0.189894
R1151 CS_BIAS.n463 CS_BIAS.n462 0.189894
R1152 CS_BIAS.n462 CS_BIAS.n461 0.189894
R1153 CS_BIAS.n461 CS_BIAS.n446 0.189894
R1154 CS_BIAS.n457 CS_BIAS.n446 0.189894
R1155 CS_BIAS.n457 CS_BIAS.n456 0.189894
R1156 CS_BIAS.n456 CS_BIAS.n455 0.189894
R1157 CS_BIAS.n455 CS_BIAS.n448 0.189894
R1158 CS_BIAS.n451 CS_BIAS.n448 0.189894
R1159 CS_BIAS.n426 CS_BIAS.n345 0.189894
R1160 CS_BIAS.n422 CS_BIAS.n345 0.189894
R1161 CS_BIAS.n422 CS_BIAS.n421 0.189894
R1162 CS_BIAS.n421 CS_BIAS.n420 0.189894
R1163 CS_BIAS.n420 CS_BIAS.n347 0.189894
R1164 CS_BIAS.n416 CS_BIAS.n347 0.189894
R1165 CS_BIAS.n416 CS_BIAS.n415 0.189894
R1166 CS_BIAS.n415 CS_BIAS.n414 0.189894
R1167 CS_BIAS.n414 CS_BIAS.n349 0.189894
R1168 CS_BIAS.n410 CS_BIAS.n349 0.189894
R1169 CS_BIAS.n410 CS_BIAS.n409 0.189894
R1170 CS_BIAS.n409 CS_BIAS.n408 0.189894
R1171 CS_BIAS.n408 CS_BIAS.n351 0.189894
R1172 CS_BIAS.n403 CS_BIAS.n351 0.189894
R1173 CS_BIAS.n403 CS_BIAS.n402 0.189894
R1174 CS_BIAS.n402 CS_BIAS.n401 0.189894
R1175 CS_BIAS.n401 CS_BIAS.n353 0.189894
R1176 CS_BIAS.n397 CS_BIAS.n353 0.189894
R1177 CS_BIAS.n397 CS_BIAS.n396 0.189894
R1178 CS_BIAS.n396 CS_BIAS.n395 0.189894
R1179 CS_BIAS.n395 CS_BIAS.n355 0.189894
R1180 CS_BIAS.n391 CS_BIAS.n355 0.189894
R1181 CS_BIAS.n391 CS_BIAS.n390 0.189894
R1182 CS_BIAS.n390 CS_BIAS.n389 0.189894
R1183 CS_BIAS.n389 CS_BIAS.n357 0.189894
R1184 CS_BIAS.n384 CS_BIAS.n357 0.189894
R1185 CS_BIAS.n384 CS_BIAS.n383 0.189894
R1186 CS_BIAS.n383 CS_BIAS.n382 0.189894
R1187 CS_BIAS.n382 CS_BIAS.n359 0.189894
R1188 CS_BIAS.n378 CS_BIAS.n359 0.189894
R1189 CS_BIAS.n378 CS_BIAS.n377 0.189894
R1190 CS_BIAS.n377 CS_BIAS.n376 0.189894
R1191 CS_BIAS.n376 CS_BIAS.n361 0.189894
R1192 CS_BIAS.n372 CS_BIAS.n361 0.189894
R1193 CS_BIAS.n372 CS_BIAS.n371 0.189894
R1194 CS_BIAS.n371 CS_BIAS.n370 0.189894
R1195 CS_BIAS.n370 CS_BIAS.n363 0.189894
R1196 CS_BIAS.n366 CS_BIAS.n363 0.189894
R1197 CS_BIAS.n341 CS_BIAS.n260 0.189894
R1198 CS_BIAS.n337 CS_BIAS.n260 0.189894
R1199 CS_BIAS.n337 CS_BIAS.n336 0.189894
R1200 CS_BIAS.n336 CS_BIAS.n335 0.189894
R1201 CS_BIAS.n335 CS_BIAS.n262 0.189894
R1202 CS_BIAS.n331 CS_BIAS.n262 0.189894
R1203 CS_BIAS.n331 CS_BIAS.n330 0.189894
R1204 CS_BIAS.n330 CS_BIAS.n329 0.189894
R1205 CS_BIAS.n329 CS_BIAS.n264 0.189894
R1206 CS_BIAS.n325 CS_BIAS.n264 0.189894
R1207 CS_BIAS.n325 CS_BIAS.n324 0.189894
R1208 CS_BIAS.n324 CS_BIAS.n323 0.189894
R1209 CS_BIAS.n323 CS_BIAS.n266 0.189894
R1210 CS_BIAS.n318 CS_BIAS.n266 0.189894
R1211 CS_BIAS.n318 CS_BIAS.n317 0.189894
R1212 CS_BIAS.n317 CS_BIAS.n316 0.189894
R1213 CS_BIAS.n316 CS_BIAS.n268 0.189894
R1214 CS_BIAS.n312 CS_BIAS.n268 0.189894
R1215 CS_BIAS.n312 CS_BIAS.n311 0.189894
R1216 CS_BIAS.n311 CS_BIAS.n310 0.189894
R1217 CS_BIAS.n310 CS_BIAS.n270 0.189894
R1218 CS_BIAS.n306 CS_BIAS.n270 0.189894
R1219 CS_BIAS.n306 CS_BIAS.n305 0.189894
R1220 CS_BIAS.n305 CS_BIAS.n304 0.189894
R1221 CS_BIAS.n304 CS_BIAS.n272 0.189894
R1222 CS_BIAS.n299 CS_BIAS.n272 0.189894
R1223 CS_BIAS.n299 CS_BIAS.n298 0.189894
R1224 CS_BIAS.n298 CS_BIAS.n297 0.189894
R1225 CS_BIAS.n297 CS_BIAS.n274 0.189894
R1226 CS_BIAS.n293 CS_BIAS.n274 0.189894
R1227 CS_BIAS.n293 CS_BIAS.n292 0.189894
R1228 CS_BIAS.n292 CS_BIAS.n291 0.189894
R1229 CS_BIAS.n291 CS_BIAS.n276 0.189894
R1230 CS_BIAS.n287 CS_BIAS.n276 0.189894
R1231 CS_BIAS.n287 CS_BIAS.n286 0.189894
R1232 CS_BIAS.n286 CS_BIAS.n285 0.189894
R1233 CS_BIAS.n285 CS_BIAS.n278 0.189894
R1234 CS_BIAS.n281 CS_BIAS.n278 0.189894
R1235 CS_BIAS.n256 CS_BIAS.n175 0.189894
R1236 CS_BIAS.n252 CS_BIAS.n175 0.189894
R1237 CS_BIAS.n252 CS_BIAS.n251 0.189894
R1238 CS_BIAS.n251 CS_BIAS.n250 0.189894
R1239 CS_BIAS.n250 CS_BIAS.n177 0.189894
R1240 CS_BIAS.n246 CS_BIAS.n177 0.189894
R1241 CS_BIAS.n246 CS_BIAS.n245 0.189894
R1242 CS_BIAS.n245 CS_BIAS.n244 0.189894
R1243 CS_BIAS.n244 CS_BIAS.n179 0.189894
R1244 CS_BIAS.n240 CS_BIAS.n179 0.189894
R1245 CS_BIAS.n240 CS_BIAS.n239 0.189894
R1246 CS_BIAS.n239 CS_BIAS.n238 0.189894
R1247 CS_BIAS.n238 CS_BIAS.n181 0.189894
R1248 CS_BIAS.n233 CS_BIAS.n181 0.189894
R1249 CS_BIAS.n233 CS_BIAS.n232 0.189894
R1250 CS_BIAS.n232 CS_BIAS.n231 0.189894
R1251 CS_BIAS.n231 CS_BIAS.n183 0.189894
R1252 CS_BIAS.n227 CS_BIAS.n183 0.189894
R1253 CS_BIAS.n227 CS_BIAS.n226 0.189894
R1254 CS_BIAS.n226 CS_BIAS.n225 0.189894
R1255 CS_BIAS.n225 CS_BIAS.n185 0.189894
R1256 CS_BIAS.n221 CS_BIAS.n185 0.189894
R1257 CS_BIAS.n221 CS_BIAS.n220 0.189894
R1258 CS_BIAS.n220 CS_BIAS.n219 0.189894
R1259 CS_BIAS.n219 CS_BIAS.n187 0.189894
R1260 CS_BIAS.n214 CS_BIAS.n187 0.189894
R1261 CS_BIAS.n214 CS_BIAS.n213 0.189894
R1262 CS_BIAS.n213 CS_BIAS.n212 0.189894
R1263 CS_BIAS.n212 CS_BIAS.n189 0.189894
R1264 CS_BIAS.n208 CS_BIAS.n189 0.189894
R1265 CS_BIAS.n208 CS_BIAS.n207 0.189894
R1266 CS_BIAS.n207 CS_BIAS.n206 0.189894
R1267 CS_BIAS.n206 CS_BIAS.n191 0.189894
R1268 CS_BIAS.n202 CS_BIAS.n191 0.189894
R1269 CS_BIAS.n202 CS_BIAS.n201 0.189894
R1270 CS_BIAS.n201 CS_BIAS.n200 0.189894
R1271 CS_BIAS.n200 CS_BIAS.n193 0.189894
R1272 CS_BIAS.n196 CS_BIAS.n193 0.189894
R1273 CS_BIAS.n97 CS_BIAS.n16 0.189894
R1274 CS_BIAS.n93 CS_BIAS.n16 0.189894
R1275 CS_BIAS.n93 CS_BIAS.n92 0.189894
R1276 CS_BIAS.n92 CS_BIAS.n91 0.189894
R1277 CS_BIAS.n91 CS_BIAS.n18 0.189894
R1278 CS_BIAS.n87 CS_BIAS.n18 0.189894
R1279 CS_BIAS.n87 CS_BIAS.n86 0.189894
R1280 CS_BIAS.n86 CS_BIAS.n85 0.189894
R1281 CS_BIAS.n85 CS_BIAS.n20 0.189894
R1282 CS_BIAS.n81 CS_BIAS.n20 0.189894
R1283 CS_BIAS.n81 CS_BIAS.n80 0.189894
R1284 CS_BIAS.n80 CS_BIAS.n79 0.189894
R1285 CS_BIAS.n79 CS_BIAS.n22 0.189894
R1286 CS_BIAS.n74 CS_BIAS.n22 0.189894
R1287 CS_BIAS.n74 CS_BIAS.n73 0.189894
R1288 CS_BIAS.n73 CS_BIAS.n72 0.189894
R1289 CS_BIAS.n72 CS_BIAS.n24 0.189894
R1290 CS_BIAS.n68 CS_BIAS.n24 0.189894
R1291 CS_BIAS.n68 CS_BIAS.n67 0.189894
R1292 CS_BIAS.n67 CS_BIAS.n66 0.189894
R1293 CS_BIAS.n66 CS_BIAS.n26 0.189894
R1294 CS_BIAS.n62 CS_BIAS.n26 0.189894
R1295 CS_BIAS.n62 CS_BIAS.n61 0.189894
R1296 CS_BIAS.n61 CS_BIAS.n60 0.189894
R1297 CS_BIAS.n60 CS_BIAS.n28 0.189894
R1298 CS_BIAS.n55 CS_BIAS.n28 0.189894
R1299 CS_BIAS.n55 CS_BIAS.n54 0.189894
R1300 CS_BIAS.n54 CS_BIAS.n53 0.189894
R1301 CS_BIAS.n53 CS_BIAS.n30 0.189894
R1302 CS_BIAS.n49 CS_BIAS.n30 0.189894
R1303 CS_BIAS.n49 CS_BIAS.n48 0.189894
R1304 CS_BIAS.n48 CS_BIAS.n47 0.189894
R1305 CS_BIAS.n47 CS_BIAS.n32 0.189894
R1306 CS_BIAS.n43 CS_BIAS.n32 0.189894
R1307 CS_BIAS.n43 CS_BIAS.n42 0.189894
R1308 CS_BIAS.n42 CS_BIAS.n41 0.189894
R1309 CS_BIAS.n41 CS_BIAS.n34 0.189894
R1310 CS_BIAS.n37 CS_BIAS.n34 0.189894
R1311 CS_BIAS.n130 CS_BIAS.n129 0.189894
R1312 CS_BIAS.n129 CS_BIAS.n128 0.189894
R1313 CS_BIAS.n128 CS_BIAS.n105 0.189894
R1314 CS_BIAS.n124 CS_BIAS.n105 0.189894
R1315 CS_BIAS.n124 CS_BIAS.n123 0.189894
R1316 CS_BIAS.n123 CS_BIAS.n122 0.189894
R1317 CS_BIAS.n122 CS_BIAS.n107 0.189894
R1318 CS_BIAS.n118 CS_BIAS.n107 0.189894
R1319 CS_BIAS.n118 CS_BIAS.n117 0.189894
R1320 CS_BIAS.n117 CS_BIAS.n116 0.189894
R1321 CS_BIAS.n116 CS_BIAS.n109 0.189894
R1322 CS_BIAS.n112 CS_BIAS.n109 0.189894
R1323 CS_BIAS.n172 CS_BIAS.n1 0.189894
R1324 CS_BIAS.n168 CS_BIAS.n1 0.189894
R1325 CS_BIAS.n168 CS_BIAS.n167 0.189894
R1326 CS_BIAS.n167 CS_BIAS.n166 0.189894
R1327 CS_BIAS.n166 CS_BIAS.n3 0.189894
R1328 CS_BIAS.n162 CS_BIAS.n3 0.189894
R1329 CS_BIAS.n162 CS_BIAS.n161 0.189894
R1330 CS_BIAS.n161 CS_BIAS.n160 0.189894
R1331 CS_BIAS.n160 CS_BIAS.n5 0.189894
R1332 CS_BIAS.n156 CS_BIAS.n5 0.189894
R1333 CS_BIAS.n156 CS_BIAS.n155 0.189894
R1334 CS_BIAS.n155 CS_BIAS.n154 0.189894
R1335 CS_BIAS.n154 CS_BIAS.n7 0.189894
R1336 CS_BIAS.n149 CS_BIAS.n7 0.189894
R1337 CS_BIAS.n149 CS_BIAS.n148 0.189894
R1338 CS_BIAS.n148 CS_BIAS.n147 0.189894
R1339 CS_BIAS.n147 CS_BIAS.n9 0.189894
R1340 CS_BIAS.n143 CS_BIAS.n9 0.189894
R1341 CS_BIAS.n143 CS_BIAS.n142 0.189894
R1342 CS_BIAS.n142 CS_BIAS.n141 0.189894
R1343 CS_BIAS.n141 CS_BIAS.n11 0.189894
R1344 CS_BIAS.n137 CS_BIAS.n11 0.189894
R1345 CS_BIAS.n137 CS_BIAS.n136 0.189894
R1346 CS_BIAS.n136 CS_BIAS.n135 0.189894
R1347 CS_BIAS.n135 CS_BIAS.n13 0.189894
R1348 CS_BIAS.n965 CS_BIAS.n962 0.189894
R1349 CS_BIAS.n969 CS_BIAS.n962 0.189894
R1350 CS_BIAS.n970 CS_BIAS.n969 0.189894
R1351 CS_BIAS.n971 CS_BIAS.n970 0.189894
R1352 CS_BIAS.n971 CS_BIAS.n960 0.189894
R1353 CS_BIAS.n975 CS_BIAS.n960 0.189894
R1354 CS_BIAS.n976 CS_BIAS.n975 0.189894
R1355 CS_BIAS.n977 CS_BIAS.n976 0.189894
R1356 CS_BIAS.n977 CS_BIAS.n958 0.189894
R1357 CS_BIAS.n981 CS_BIAS.n958 0.189894
R1358 CS_BIAS.n982 CS_BIAS.n981 0.189894
R1359 CS_BIAS.n983 CS_BIAS.n982 0.189894
R1360 CS_BIAS.n983 CS_BIAS.n956 0.189894
R1361 CS_BIAS.n988 CS_BIAS.n956 0.189894
R1362 CS_BIAS.n989 CS_BIAS.n988 0.189894
R1363 CS_BIAS.n990 CS_BIAS.n989 0.189894
R1364 CS_BIAS.n990 CS_BIAS.n954 0.189894
R1365 CS_BIAS.n994 CS_BIAS.n954 0.189894
R1366 CS_BIAS.n995 CS_BIAS.n994 0.189894
R1367 CS_BIAS.n996 CS_BIAS.n995 0.189894
R1368 CS_BIAS.n996 CS_BIAS.n952 0.189894
R1369 CS_BIAS.n1000 CS_BIAS.n952 0.189894
R1370 CS_BIAS.n1001 CS_BIAS.n1000 0.189894
R1371 CS_BIAS.n1002 CS_BIAS.n1001 0.189894
R1372 CS_BIAS.n1002 CS_BIAS.n950 0.189894
R1373 CS_BIAS.n1007 CS_BIAS.n950 0.189894
R1374 CS_BIAS.n1008 CS_BIAS.n1007 0.189894
R1375 CS_BIAS.n1009 CS_BIAS.n1008 0.189894
R1376 CS_BIAS.n1009 CS_BIAS.n948 0.189894
R1377 CS_BIAS.n1013 CS_BIAS.n948 0.189894
R1378 CS_BIAS.n1014 CS_BIAS.n1013 0.189894
R1379 CS_BIAS.n1015 CS_BIAS.n1014 0.189894
R1380 CS_BIAS.n1015 CS_BIAS.n946 0.189894
R1381 CS_BIAS.n1019 CS_BIAS.n946 0.189894
R1382 CS_BIAS.n1020 CS_BIAS.n1019 0.189894
R1383 CS_BIAS.n1021 CS_BIAS.n1020 0.189894
R1384 CS_BIAS.n1021 CS_BIAS.n944 0.189894
R1385 CS_BIAS.n1025 CS_BIAS.n944 0.189894
R1386 CS_BIAS.n880 CS_BIAS.n877 0.189894
R1387 CS_BIAS.n884 CS_BIAS.n877 0.189894
R1388 CS_BIAS.n885 CS_BIAS.n884 0.189894
R1389 CS_BIAS.n886 CS_BIAS.n885 0.189894
R1390 CS_BIAS.n886 CS_BIAS.n875 0.189894
R1391 CS_BIAS.n890 CS_BIAS.n875 0.189894
R1392 CS_BIAS.n891 CS_BIAS.n890 0.189894
R1393 CS_BIAS.n892 CS_BIAS.n891 0.189894
R1394 CS_BIAS.n892 CS_BIAS.n873 0.189894
R1395 CS_BIAS.n896 CS_BIAS.n873 0.189894
R1396 CS_BIAS.n897 CS_BIAS.n896 0.189894
R1397 CS_BIAS.n898 CS_BIAS.n897 0.189894
R1398 CS_BIAS.n898 CS_BIAS.n871 0.189894
R1399 CS_BIAS.n903 CS_BIAS.n871 0.189894
R1400 CS_BIAS.n904 CS_BIAS.n903 0.189894
R1401 CS_BIAS.n905 CS_BIAS.n904 0.189894
R1402 CS_BIAS.n905 CS_BIAS.n869 0.189894
R1403 CS_BIAS.n909 CS_BIAS.n869 0.189894
R1404 CS_BIAS.n910 CS_BIAS.n909 0.189894
R1405 CS_BIAS.n911 CS_BIAS.n910 0.189894
R1406 CS_BIAS.n911 CS_BIAS.n867 0.189894
R1407 CS_BIAS.n915 CS_BIAS.n867 0.189894
R1408 CS_BIAS.n916 CS_BIAS.n915 0.189894
R1409 CS_BIAS.n917 CS_BIAS.n916 0.189894
R1410 CS_BIAS.n917 CS_BIAS.n865 0.189894
R1411 CS_BIAS.n922 CS_BIAS.n865 0.189894
R1412 CS_BIAS.n923 CS_BIAS.n922 0.189894
R1413 CS_BIAS.n924 CS_BIAS.n923 0.189894
R1414 CS_BIAS.n924 CS_BIAS.n863 0.189894
R1415 CS_BIAS.n928 CS_BIAS.n863 0.189894
R1416 CS_BIAS.n929 CS_BIAS.n928 0.189894
R1417 CS_BIAS.n930 CS_BIAS.n929 0.189894
R1418 CS_BIAS.n930 CS_BIAS.n861 0.189894
R1419 CS_BIAS.n934 CS_BIAS.n861 0.189894
R1420 CS_BIAS.n935 CS_BIAS.n934 0.189894
R1421 CS_BIAS.n936 CS_BIAS.n935 0.189894
R1422 CS_BIAS.n936 CS_BIAS.n859 0.189894
R1423 CS_BIAS.n940 CS_BIAS.n859 0.189894
R1424 CS_BIAS.n795 CS_BIAS.n792 0.189894
R1425 CS_BIAS.n799 CS_BIAS.n792 0.189894
R1426 CS_BIAS.n800 CS_BIAS.n799 0.189894
R1427 CS_BIAS.n801 CS_BIAS.n800 0.189894
R1428 CS_BIAS.n801 CS_BIAS.n790 0.189894
R1429 CS_BIAS.n805 CS_BIAS.n790 0.189894
R1430 CS_BIAS.n806 CS_BIAS.n805 0.189894
R1431 CS_BIAS.n807 CS_BIAS.n806 0.189894
R1432 CS_BIAS.n807 CS_BIAS.n788 0.189894
R1433 CS_BIAS.n811 CS_BIAS.n788 0.189894
R1434 CS_BIAS.n812 CS_BIAS.n811 0.189894
R1435 CS_BIAS.n813 CS_BIAS.n812 0.189894
R1436 CS_BIAS.n813 CS_BIAS.n786 0.189894
R1437 CS_BIAS.n818 CS_BIAS.n786 0.189894
R1438 CS_BIAS.n819 CS_BIAS.n818 0.189894
R1439 CS_BIAS.n820 CS_BIAS.n819 0.189894
R1440 CS_BIAS.n820 CS_BIAS.n784 0.189894
R1441 CS_BIAS.n824 CS_BIAS.n784 0.189894
R1442 CS_BIAS.n825 CS_BIAS.n824 0.189894
R1443 CS_BIAS.n826 CS_BIAS.n825 0.189894
R1444 CS_BIAS.n826 CS_BIAS.n782 0.189894
R1445 CS_BIAS.n830 CS_BIAS.n782 0.189894
R1446 CS_BIAS.n831 CS_BIAS.n830 0.189894
R1447 CS_BIAS.n832 CS_BIAS.n831 0.189894
R1448 CS_BIAS.n832 CS_BIAS.n780 0.189894
R1449 CS_BIAS.n837 CS_BIAS.n780 0.189894
R1450 CS_BIAS.n838 CS_BIAS.n837 0.189894
R1451 CS_BIAS.n839 CS_BIAS.n838 0.189894
R1452 CS_BIAS.n839 CS_BIAS.n778 0.189894
R1453 CS_BIAS.n843 CS_BIAS.n778 0.189894
R1454 CS_BIAS.n844 CS_BIAS.n843 0.189894
R1455 CS_BIAS.n845 CS_BIAS.n844 0.189894
R1456 CS_BIAS.n845 CS_BIAS.n776 0.189894
R1457 CS_BIAS.n849 CS_BIAS.n776 0.189894
R1458 CS_BIAS.n850 CS_BIAS.n849 0.189894
R1459 CS_BIAS.n851 CS_BIAS.n850 0.189894
R1460 CS_BIAS.n851 CS_BIAS.n774 0.189894
R1461 CS_BIAS.n855 CS_BIAS.n774 0.189894
R1462 CS_BIAS.n710 CS_BIAS.n707 0.189894
R1463 CS_BIAS.n714 CS_BIAS.n707 0.189894
R1464 CS_BIAS.n715 CS_BIAS.n714 0.189894
R1465 CS_BIAS.n716 CS_BIAS.n715 0.189894
R1466 CS_BIAS.n716 CS_BIAS.n705 0.189894
R1467 CS_BIAS.n720 CS_BIAS.n705 0.189894
R1468 CS_BIAS.n721 CS_BIAS.n720 0.189894
R1469 CS_BIAS.n722 CS_BIAS.n721 0.189894
R1470 CS_BIAS.n722 CS_BIAS.n703 0.189894
R1471 CS_BIAS.n726 CS_BIAS.n703 0.189894
R1472 CS_BIAS.n727 CS_BIAS.n726 0.189894
R1473 CS_BIAS.n728 CS_BIAS.n727 0.189894
R1474 CS_BIAS.n728 CS_BIAS.n701 0.189894
R1475 CS_BIAS.n733 CS_BIAS.n701 0.189894
R1476 CS_BIAS.n734 CS_BIAS.n733 0.189894
R1477 CS_BIAS.n735 CS_BIAS.n734 0.189894
R1478 CS_BIAS.n735 CS_BIAS.n699 0.189894
R1479 CS_BIAS.n739 CS_BIAS.n699 0.189894
R1480 CS_BIAS.n740 CS_BIAS.n739 0.189894
R1481 CS_BIAS.n741 CS_BIAS.n740 0.189894
R1482 CS_BIAS.n741 CS_BIAS.n697 0.189894
R1483 CS_BIAS.n745 CS_BIAS.n697 0.189894
R1484 CS_BIAS.n746 CS_BIAS.n745 0.189894
R1485 CS_BIAS.n747 CS_BIAS.n746 0.189894
R1486 CS_BIAS.n747 CS_BIAS.n695 0.189894
R1487 CS_BIAS.n752 CS_BIAS.n695 0.189894
R1488 CS_BIAS.n753 CS_BIAS.n752 0.189894
R1489 CS_BIAS.n754 CS_BIAS.n753 0.189894
R1490 CS_BIAS.n754 CS_BIAS.n693 0.189894
R1491 CS_BIAS.n758 CS_BIAS.n693 0.189894
R1492 CS_BIAS.n759 CS_BIAS.n758 0.189894
R1493 CS_BIAS.n760 CS_BIAS.n759 0.189894
R1494 CS_BIAS.n760 CS_BIAS.n691 0.189894
R1495 CS_BIAS.n764 CS_BIAS.n691 0.189894
R1496 CS_BIAS.n765 CS_BIAS.n764 0.189894
R1497 CS_BIAS.n766 CS_BIAS.n765 0.189894
R1498 CS_BIAS.n766 CS_BIAS.n689 0.189894
R1499 CS_BIAS.n770 CS_BIAS.n689 0.189894
R1500 CS_BIAS.n578 CS_BIAS.n575 0.189894
R1501 CS_BIAS.n582 CS_BIAS.n575 0.189894
R1502 CS_BIAS.n583 CS_BIAS.n582 0.189894
R1503 CS_BIAS.n584 CS_BIAS.n583 0.189894
R1504 CS_BIAS.n584 CS_BIAS.n573 0.189894
R1505 CS_BIAS.n588 CS_BIAS.n573 0.189894
R1506 CS_BIAS.n589 CS_BIAS.n588 0.189894
R1507 CS_BIAS.n590 CS_BIAS.n589 0.189894
R1508 CS_BIAS.n590 CS_BIAS.n571 0.189894
R1509 CS_BIAS.n594 CS_BIAS.n571 0.189894
R1510 CS_BIAS.n595 CS_BIAS.n594 0.189894
R1511 CS_BIAS.n596 CS_BIAS.n595 0.189894
R1512 CS_BIAS.n596 CS_BIAS.n569 0.189894
R1513 CS_BIAS.n601 CS_BIAS.n569 0.189894
R1514 CS_BIAS.n602 CS_BIAS.n601 0.189894
R1515 CS_BIAS.n603 CS_BIAS.n602 0.189894
R1516 CS_BIAS.n603 CS_BIAS.n567 0.189894
R1517 CS_BIAS.n607 CS_BIAS.n567 0.189894
R1518 CS_BIAS.n608 CS_BIAS.n607 0.189894
R1519 CS_BIAS.n609 CS_BIAS.n608 0.189894
R1520 CS_BIAS.n609 CS_BIAS.n565 0.189894
R1521 CS_BIAS.n613 CS_BIAS.n565 0.189894
R1522 CS_BIAS.n614 CS_BIAS.n613 0.189894
R1523 CS_BIAS.n615 CS_BIAS.n614 0.189894
R1524 CS_BIAS.n615 CS_BIAS.n563 0.189894
R1525 CS_BIAS.n620 CS_BIAS.n563 0.189894
R1526 CS_BIAS.n621 CS_BIAS.n620 0.189894
R1527 CS_BIAS.n622 CS_BIAS.n621 0.189894
R1528 CS_BIAS.n622 CS_BIAS.n561 0.189894
R1529 CS_BIAS.n626 CS_BIAS.n561 0.189894
R1530 CS_BIAS.n627 CS_BIAS.n626 0.189894
R1531 CS_BIAS.n628 CS_BIAS.n627 0.189894
R1532 CS_BIAS.n628 CS_BIAS.n559 0.189894
R1533 CS_BIAS.n632 CS_BIAS.n559 0.189894
R1534 CS_BIAS.n633 CS_BIAS.n632 0.189894
R1535 CS_BIAS.n634 CS_BIAS.n633 0.189894
R1536 CS_BIAS.n634 CS_BIAS.n557 0.189894
R1537 CS_BIAS.n638 CS_BIAS.n557 0.189894
R1538 CS_BIAS.n536 CS_BIAS.n533 0.189894
R1539 CS_BIAS.n540 CS_BIAS.n533 0.189894
R1540 CS_BIAS.n541 CS_BIAS.n540 0.189894
R1541 CS_BIAS.n542 CS_BIAS.n541 0.189894
R1542 CS_BIAS.n542 CS_BIAS.n531 0.189894
R1543 CS_BIAS.n546 CS_BIAS.n531 0.189894
R1544 CS_BIAS.n547 CS_BIAS.n546 0.189894
R1545 CS_BIAS.n548 CS_BIAS.n547 0.189894
R1546 CS_BIAS.n548 CS_BIAS.n529 0.189894
R1547 CS_BIAS.n552 CS_BIAS.n529 0.189894
R1548 CS_BIAS.n553 CS_BIAS.n552 0.189894
R1549 CS_BIAS.n644 CS_BIAS.n553 0.189894
R1550 CS_BIAS.n649 CS_BIAS.n527 0.189894
R1551 CS_BIAS.n650 CS_BIAS.n649 0.189894
R1552 CS_BIAS.n651 CS_BIAS.n650 0.189894
R1553 CS_BIAS.n651 CS_BIAS.n525 0.189894
R1554 CS_BIAS.n655 CS_BIAS.n525 0.189894
R1555 CS_BIAS.n656 CS_BIAS.n655 0.189894
R1556 CS_BIAS.n657 CS_BIAS.n656 0.189894
R1557 CS_BIAS.n657 CS_BIAS.n523 0.189894
R1558 CS_BIAS.n661 CS_BIAS.n523 0.189894
R1559 CS_BIAS.n662 CS_BIAS.n661 0.189894
R1560 CS_BIAS.n663 CS_BIAS.n662 0.189894
R1561 CS_BIAS.n663 CS_BIAS.n521 0.189894
R1562 CS_BIAS.n668 CS_BIAS.n521 0.189894
R1563 CS_BIAS.n669 CS_BIAS.n668 0.189894
R1564 CS_BIAS.n670 CS_BIAS.n669 0.189894
R1565 CS_BIAS.n670 CS_BIAS.n519 0.189894
R1566 CS_BIAS.n674 CS_BIAS.n519 0.189894
R1567 CS_BIAS.n675 CS_BIAS.n674 0.189894
R1568 CS_BIAS.n676 CS_BIAS.n675 0.189894
R1569 CS_BIAS.n676 CS_BIAS.n517 0.189894
R1570 CS_BIAS.n680 CS_BIAS.n517 0.189894
R1571 CS_BIAS.n681 CS_BIAS.n680 0.189894
R1572 CS_BIAS.n682 CS_BIAS.n681 0.189894
R1573 CS_BIAS.n682 CS_BIAS.n515 0.189894
R1574 CS_BIAS.n686 CS_BIAS.n515 0.189894
R1575 CS_BIAS.n130 CS_BIAS.n104 0.0762576
R1576 CS_BIAS.n104 CS_BIAS.n13 0.0762576
R1577 CS_BIAS.n644 CS_BIAS.n643 0.0762576
R1578 CS_BIAS.n643 CS_BIAS.n527 0.0762576
R1579 GND.n2976 GND.n2975 5638.7
R1580 GND.n3960 GND.n3779 1822.22
R1581 GND.n8447 GND.n384 788
R1582 GND.n8329 GND.n8328 788
R1583 GND.n7711 GND.n669 788
R1584 GND.n7699 GND.n671 788
R1585 GND.n6281 GND.n1632 788
R1586 GND.n6287 GND.n1629 788
R1587 GND.n2541 GND.n2540 788
R1588 GND.n2973 GND.n2466 788
R1589 GND.n4729 GND.n3022 783.196
R1590 GND.n3961 GND.n3780 783.196
R1591 GND.n8457 GND.n344 783.196
R1592 GND.n4845 GND.n2427 783.196
R1593 GND.n6983 GND.n1177 778.39
R1594 GND.n6932 GND.n1174 778.39
R1595 GND.n6376 GND.n6375 778.39
R1596 GND.n6315 GND.n6314 778.39
R1597 GND.n451 GND.n351 763.976
R1598 GND.n8217 GND.n8216 763.976
R1599 GND.n711 GND.n673 763.976
R1600 GND.n1225 GND.n672 763.976
R1601 GND.n2864 GND.n2863 763.976
R1602 GND.n6285 GND.n6284 763.976
R1603 GND.n2604 GND.n2462 763.976
R1604 GND.n1660 GND.n1633 763.976
R1605 GND.n6284 GND.n1618 589.749
R1606 GND.n1660 GND.n1623 589.052
R1607 GND.n1204 GND.n711 589.052
R1608 GND.n4729 GND.n4728 585
R1609 GND.n4731 GND.n3021 585
R1610 GND.n4734 GND.n4733 585
R1611 GND.n3019 GND.n3018 585
R1612 GND.n4739 GND.n4738 585
R1613 GND.n4741 GND.n3017 585
R1614 GND.n4744 GND.n4743 585
R1615 GND.n3015 GND.n3014 585
R1616 GND.n4749 GND.n4748 585
R1617 GND.n4751 GND.n3013 585
R1618 GND.n4754 GND.n4753 585
R1619 GND.n3011 GND.n3010 585
R1620 GND.n4759 GND.n4758 585
R1621 GND.n4761 GND.n3009 585
R1622 GND.n4764 GND.n4763 585
R1623 GND.n3007 GND.n3006 585
R1624 GND.n4769 GND.n4768 585
R1625 GND.n4771 GND.n3005 585
R1626 GND.n4774 GND.n4773 585
R1627 GND.n3003 GND.n3002 585
R1628 GND.n4779 GND.n4778 585
R1629 GND.n4781 GND.n3001 585
R1630 GND.n4784 GND.n4783 585
R1631 GND.n2999 GND.n2998 585
R1632 GND.n4789 GND.n4788 585
R1633 GND.n4791 GND.n2997 585
R1634 GND.n4794 GND.n4793 585
R1635 GND.n2995 GND.n2994 585
R1636 GND.n4799 GND.n4798 585
R1637 GND.n4801 GND.n2993 585
R1638 GND.n4804 GND.n4803 585
R1639 GND.n2991 GND.n2990 585
R1640 GND.n4809 GND.n4808 585
R1641 GND.n4811 GND.n2989 585
R1642 GND.n4814 GND.n4813 585
R1643 GND.n2987 GND.n2986 585
R1644 GND.n4819 GND.n4818 585
R1645 GND.n4821 GND.n2985 585
R1646 GND.n4824 GND.n4823 585
R1647 GND.n2983 GND.n2982 585
R1648 GND.n4829 GND.n4828 585
R1649 GND.n4831 GND.n2981 585
R1650 GND.n4834 GND.n4833 585
R1651 GND.n2979 GND.n2978 585
R1652 GND.n4840 GND.n4839 585
R1653 GND.n4842 GND.n2977 585
R1654 GND.n4843 GND.n2430 585
R1655 GND.n4846 GND.n4845 585
R1656 GND.n4725 GND.n3022 585
R1657 GND.n3026 GND.n3022 585
R1658 GND.n4724 GND.n4723 585
R1659 GND.n4723 GND.n4722 585
R1660 GND.n3025 GND.n3024 585
R1661 GND.n4721 GND.n3025 585
R1662 GND.n4719 GND.n4718 585
R1663 GND.n4720 GND.n4719 585
R1664 GND.n4717 GND.n3028 585
R1665 GND.n3028 GND.n3027 585
R1666 GND.n4716 GND.n4715 585
R1667 GND.n4715 GND.n4714 585
R1668 GND.n3034 GND.n3033 585
R1669 GND.n4713 GND.n3034 585
R1670 GND.n4711 GND.n4710 585
R1671 GND.n4712 GND.n4711 585
R1672 GND.n4709 GND.n3036 585
R1673 GND.n3036 GND.n3035 585
R1674 GND.n4708 GND.n4707 585
R1675 GND.n4707 GND.n4706 585
R1676 GND.n3042 GND.n3041 585
R1677 GND.n4705 GND.n3042 585
R1678 GND.n4703 GND.n4702 585
R1679 GND.n4704 GND.n4703 585
R1680 GND.n4701 GND.n3044 585
R1681 GND.n3044 GND.n3043 585
R1682 GND.n4700 GND.n4699 585
R1683 GND.n4699 GND.n4698 585
R1684 GND.n3050 GND.n3049 585
R1685 GND.n4697 GND.n3050 585
R1686 GND.n4695 GND.n4694 585
R1687 GND.n4696 GND.n4695 585
R1688 GND.n4693 GND.n3052 585
R1689 GND.n3052 GND.n3051 585
R1690 GND.n4692 GND.n4691 585
R1691 GND.n4691 GND.n4690 585
R1692 GND.n3058 GND.n3057 585
R1693 GND.n4689 GND.n3058 585
R1694 GND.n4687 GND.n4686 585
R1695 GND.n4688 GND.n4687 585
R1696 GND.n4685 GND.n3060 585
R1697 GND.n3060 GND.n3059 585
R1698 GND.n4684 GND.n4683 585
R1699 GND.n4683 GND.n4682 585
R1700 GND.n3066 GND.n3065 585
R1701 GND.n4681 GND.n3066 585
R1702 GND.n4679 GND.n4678 585
R1703 GND.n4680 GND.n4679 585
R1704 GND.n4677 GND.n3068 585
R1705 GND.n3068 GND.n3067 585
R1706 GND.n4676 GND.n4675 585
R1707 GND.n4675 GND.n4674 585
R1708 GND.n3074 GND.n3073 585
R1709 GND.n4673 GND.n3074 585
R1710 GND.n4671 GND.n4670 585
R1711 GND.n4672 GND.n4671 585
R1712 GND.n4669 GND.n3076 585
R1713 GND.n3076 GND.n3075 585
R1714 GND.n4668 GND.n4667 585
R1715 GND.n4667 GND.n4666 585
R1716 GND.n3082 GND.n3081 585
R1717 GND.n4665 GND.n3082 585
R1718 GND.n4663 GND.n4662 585
R1719 GND.n4664 GND.n4663 585
R1720 GND.n4661 GND.n3084 585
R1721 GND.n3084 GND.n3083 585
R1722 GND.n4660 GND.n4659 585
R1723 GND.n4659 GND.n4658 585
R1724 GND.n3090 GND.n3089 585
R1725 GND.n4657 GND.n3090 585
R1726 GND.n4655 GND.n4654 585
R1727 GND.n4656 GND.n4655 585
R1728 GND.n4653 GND.n3092 585
R1729 GND.n3092 GND.n3091 585
R1730 GND.n4652 GND.n4651 585
R1731 GND.n4651 GND.n4650 585
R1732 GND.n3098 GND.n3097 585
R1733 GND.n4649 GND.n3098 585
R1734 GND.n4647 GND.n4646 585
R1735 GND.n4648 GND.n4647 585
R1736 GND.n4645 GND.n3100 585
R1737 GND.n3100 GND.n3099 585
R1738 GND.n4644 GND.n4643 585
R1739 GND.n4643 GND.n4642 585
R1740 GND.n3106 GND.n3105 585
R1741 GND.n4641 GND.n3106 585
R1742 GND.n4639 GND.n4638 585
R1743 GND.n4640 GND.n4639 585
R1744 GND.n4637 GND.n3108 585
R1745 GND.n3108 GND.n3107 585
R1746 GND.n4636 GND.n4635 585
R1747 GND.n4635 GND.n4634 585
R1748 GND.n3114 GND.n3113 585
R1749 GND.n4633 GND.n3114 585
R1750 GND.n4631 GND.n4630 585
R1751 GND.n4632 GND.n4631 585
R1752 GND.n4629 GND.n3116 585
R1753 GND.n3116 GND.n3115 585
R1754 GND.n4628 GND.n4627 585
R1755 GND.n4627 GND.n4626 585
R1756 GND.n3122 GND.n3121 585
R1757 GND.n4625 GND.n3122 585
R1758 GND.n4623 GND.n4622 585
R1759 GND.n4624 GND.n4623 585
R1760 GND.n4621 GND.n3124 585
R1761 GND.n3124 GND.n3123 585
R1762 GND.n4620 GND.n4619 585
R1763 GND.n4619 GND.n4618 585
R1764 GND.n3130 GND.n3129 585
R1765 GND.n4617 GND.n3130 585
R1766 GND.n4615 GND.n4614 585
R1767 GND.n4616 GND.n4615 585
R1768 GND.n4613 GND.n3132 585
R1769 GND.n3132 GND.n3131 585
R1770 GND.n4612 GND.n4611 585
R1771 GND.n4611 GND.n4610 585
R1772 GND.n3138 GND.n3137 585
R1773 GND.n4609 GND.n3138 585
R1774 GND.n4607 GND.n4606 585
R1775 GND.n4608 GND.n4607 585
R1776 GND.n4605 GND.n3140 585
R1777 GND.n3140 GND.n3139 585
R1778 GND.n4604 GND.n4603 585
R1779 GND.n4603 GND.n4602 585
R1780 GND.n3146 GND.n3145 585
R1781 GND.n4601 GND.n3146 585
R1782 GND.n4599 GND.n4598 585
R1783 GND.n4600 GND.n4599 585
R1784 GND.n4597 GND.n3148 585
R1785 GND.n3148 GND.n3147 585
R1786 GND.n4596 GND.n4595 585
R1787 GND.n4595 GND.n4594 585
R1788 GND.n3154 GND.n3153 585
R1789 GND.n4593 GND.n3154 585
R1790 GND.n4591 GND.n4590 585
R1791 GND.n4592 GND.n4591 585
R1792 GND.n4589 GND.n3156 585
R1793 GND.n3156 GND.n3155 585
R1794 GND.n4588 GND.n4587 585
R1795 GND.n4587 GND.n4586 585
R1796 GND.n3162 GND.n3161 585
R1797 GND.n4585 GND.n3162 585
R1798 GND.n4583 GND.n4582 585
R1799 GND.n4584 GND.n4583 585
R1800 GND.n4581 GND.n3164 585
R1801 GND.n3164 GND.n3163 585
R1802 GND.n4580 GND.n4579 585
R1803 GND.n4579 GND.n4578 585
R1804 GND.n3170 GND.n3169 585
R1805 GND.n4577 GND.n3170 585
R1806 GND.n4575 GND.n4574 585
R1807 GND.n4576 GND.n4575 585
R1808 GND.n4573 GND.n3172 585
R1809 GND.n3172 GND.n3171 585
R1810 GND.n4572 GND.n4571 585
R1811 GND.n4571 GND.n4570 585
R1812 GND.n3178 GND.n3177 585
R1813 GND.n4569 GND.n3178 585
R1814 GND.n4567 GND.n4566 585
R1815 GND.n4568 GND.n4567 585
R1816 GND.n4565 GND.n3180 585
R1817 GND.n3180 GND.n3179 585
R1818 GND.n4564 GND.n4563 585
R1819 GND.n4563 GND.n4562 585
R1820 GND.n3186 GND.n3185 585
R1821 GND.n4561 GND.n3186 585
R1822 GND.n4559 GND.n4558 585
R1823 GND.n4560 GND.n4559 585
R1824 GND.n4557 GND.n3188 585
R1825 GND.n3188 GND.n3187 585
R1826 GND.n4556 GND.n4555 585
R1827 GND.n4555 GND.n4554 585
R1828 GND.n3194 GND.n3193 585
R1829 GND.n4553 GND.n3194 585
R1830 GND.n4551 GND.n4550 585
R1831 GND.n4552 GND.n4551 585
R1832 GND.n4549 GND.n3196 585
R1833 GND.n3196 GND.n3195 585
R1834 GND.n4548 GND.n4547 585
R1835 GND.n4547 GND.n4546 585
R1836 GND.n3202 GND.n3201 585
R1837 GND.n4545 GND.n3202 585
R1838 GND.n4543 GND.n4542 585
R1839 GND.n4544 GND.n4543 585
R1840 GND.n4541 GND.n3204 585
R1841 GND.n3204 GND.n3203 585
R1842 GND.n4540 GND.n4539 585
R1843 GND.n4539 GND.n4538 585
R1844 GND.n3210 GND.n3209 585
R1845 GND.n4537 GND.n3210 585
R1846 GND.n4535 GND.n4534 585
R1847 GND.n4536 GND.n4535 585
R1848 GND.n4533 GND.n3212 585
R1849 GND.n3212 GND.n3211 585
R1850 GND.n4532 GND.n4531 585
R1851 GND.n4531 GND.n4530 585
R1852 GND.n3218 GND.n3217 585
R1853 GND.n4529 GND.n3218 585
R1854 GND.n4527 GND.n4526 585
R1855 GND.n4528 GND.n4527 585
R1856 GND.n4525 GND.n3220 585
R1857 GND.n3220 GND.n3219 585
R1858 GND.n4524 GND.n4523 585
R1859 GND.n4523 GND.n4522 585
R1860 GND.n3226 GND.n3225 585
R1861 GND.n4521 GND.n3226 585
R1862 GND.n4519 GND.n4518 585
R1863 GND.n4520 GND.n4519 585
R1864 GND.n4517 GND.n3228 585
R1865 GND.n3228 GND.n3227 585
R1866 GND.n4516 GND.n4515 585
R1867 GND.n4515 GND.n4514 585
R1868 GND.n3234 GND.n3233 585
R1869 GND.n4513 GND.n3234 585
R1870 GND.n4511 GND.n4510 585
R1871 GND.n4512 GND.n4511 585
R1872 GND.n4509 GND.n3236 585
R1873 GND.n3236 GND.n3235 585
R1874 GND.n4508 GND.n4507 585
R1875 GND.n4507 GND.n4506 585
R1876 GND.n3242 GND.n3241 585
R1877 GND.n4505 GND.n3242 585
R1878 GND.n4503 GND.n4502 585
R1879 GND.n4504 GND.n4503 585
R1880 GND.n4501 GND.n3244 585
R1881 GND.n3244 GND.n3243 585
R1882 GND.n4500 GND.n4499 585
R1883 GND.n4499 GND.n4498 585
R1884 GND.n3250 GND.n3249 585
R1885 GND.n4497 GND.n3250 585
R1886 GND.n4495 GND.n4494 585
R1887 GND.n4496 GND.n4495 585
R1888 GND.n4493 GND.n3252 585
R1889 GND.n3252 GND.n3251 585
R1890 GND.n4492 GND.n4491 585
R1891 GND.n4491 GND.n4490 585
R1892 GND.n3258 GND.n3257 585
R1893 GND.n4489 GND.n3258 585
R1894 GND.n4487 GND.n4486 585
R1895 GND.n4488 GND.n4487 585
R1896 GND.n4485 GND.n3260 585
R1897 GND.n3260 GND.n3259 585
R1898 GND.n4484 GND.n4483 585
R1899 GND.n4483 GND.n4482 585
R1900 GND.n3266 GND.n3265 585
R1901 GND.n4481 GND.n3266 585
R1902 GND.n4479 GND.n4478 585
R1903 GND.n4480 GND.n4479 585
R1904 GND.n4477 GND.n3268 585
R1905 GND.n3268 GND.n3267 585
R1906 GND.n4476 GND.n4475 585
R1907 GND.n4475 GND.n4474 585
R1908 GND.n3274 GND.n3273 585
R1909 GND.n4473 GND.n3274 585
R1910 GND.n4471 GND.n4470 585
R1911 GND.n4472 GND.n4471 585
R1912 GND.n4469 GND.n3276 585
R1913 GND.n3276 GND.n3275 585
R1914 GND.n4468 GND.n4467 585
R1915 GND.n4467 GND.n4466 585
R1916 GND.n3282 GND.n3281 585
R1917 GND.n4465 GND.n3282 585
R1918 GND.n4463 GND.n4462 585
R1919 GND.n4464 GND.n4463 585
R1920 GND.n4461 GND.n3284 585
R1921 GND.n3284 GND.n3283 585
R1922 GND.n4460 GND.n4459 585
R1923 GND.n4459 GND.n4458 585
R1924 GND.n3290 GND.n3289 585
R1925 GND.n4457 GND.n3290 585
R1926 GND.n4455 GND.n4454 585
R1927 GND.n4456 GND.n4455 585
R1928 GND.n4453 GND.n3292 585
R1929 GND.n3292 GND.n3291 585
R1930 GND.n4452 GND.n4451 585
R1931 GND.n4451 GND.n4450 585
R1932 GND.n3298 GND.n3297 585
R1933 GND.n4449 GND.n3298 585
R1934 GND.n4447 GND.n4446 585
R1935 GND.n4448 GND.n4447 585
R1936 GND.n4445 GND.n3300 585
R1937 GND.n3300 GND.n3299 585
R1938 GND.n4444 GND.n4443 585
R1939 GND.n4443 GND.n4442 585
R1940 GND.n3306 GND.n3305 585
R1941 GND.n4441 GND.n3306 585
R1942 GND.n4439 GND.n4438 585
R1943 GND.n4440 GND.n4439 585
R1944 GND.n4437 GND.n3308 585
R1945 GND.n3308 GND.n3307 585
R1946 GND.n4436 GND.n4435 585
R1947 GND.n4435 GND.n4434 585
R1948 GND.n3314 GND.n3313 585
R1949 GND.n4433 GND.n3314 585
R1950 GND.n4431 GND.n4430 585
R1951 GND.n4432 GND.n4431 585
R1952 GND.n4429 GND.n3316 585
R1953 GND.n3316 GND.n3315 585
R1954 GND.n4428 GND.n4427 585
R1955 GND.n4427 GND.n4426 585
R1956 GND.n3322 GND.n3321 585
R1957 GND.n4425 GND.n3322 585
R1958 GND.n4423 GND.n4422 585
R1959 GND.n4424 GND.n4423 585
R1960 GND.n4421 GND.n3324 585
R1961 GND.n3324 GND.n3323 585
R1962 GND.n4420 GND.n4419 585
R1963 GND.n4419 GND.n4418 585
R1964 GND.n3330 GND.n3329 585
R1965 GND.n4417 GND.n3330 585
R1966 GND.n4415 GND.n4414 585
R1967 GND.n4416 GND.n4415 585
R1968 GND.n4413 GND.n3332 585
R1969 GND.n3332 GND.n3331 585
R1970 GND.n4412 GND.n4411 585
R1971 GND.n4411 GND.n4410 585
R1972 GND.n3338 GND.n3337 585
R1973 GND.n4409 GND.n3338 585
R1974 GND.n4407 GND.n4406 585
R1975 GND.n4408 GND.n4407 585
R1976 GND.n4405 GND.n3340 585
R1977 GND.n3340 GND.n3339 585
R1978 GND.n4404 GND.n4403 585
R1979 GND.n4403 GND.n4402 585
R1980 GND.n3346 GND.n3345 585
R1981 GND.n4401 GND.n3346 585
R1982 GND.n4399 GND.n4398 585
R1983 GND.n4400 GND.n4399 585
R1984 GND.n4397 GND.n3348 585
R1985 GND.n3348 GND.n3347 585
R1986 GND.n4396 GND.n4395 585
R1987 GND.n4395 GND.n4394 585
R1988 GND.n3354 GND.n3353 585
R1989 GND.n4393 GND.n3354 585
R1990 GND.n4391 GND.n4390 585
R1991 GND.n4392 GND.n4391 585
R1992 GND.n4389 GND.n3356 585
R1993 GND.n3356 GND.n3355 585
R1994 GND.n4388 GND.n4387 585
R1995 GND.n4387 GND.n4386 585
R1996 GND.n3362 GND.n3361 585
R1997 GND.n4385 GND.n3362 585
R1998 GND.n4383 GND.n4382 585
R1999 GND.n4384 GND.n4383 585
R2000 GND.n4381 GND.n3364 585
R2001 GND.n3364 GND.n3363 585
R2002 GND.n4380 GND.n4379 585
R2003 GND.n4379 GND.n4378 585
R2004 GND.n3370 GND.n3369 585
R2005 GND.n4377 GND.n3370 585
R2006 GND.n4375 GND.n4374 585
R2007 GND.n4376 GND.n4375 585
R2008 GND.n4373 GND.n3372 585
R2009 GND.n3372 GND.n3371 585
R2010 GND.n4372 GND.n4371 585
R2011 GND.n4371 GND.n4370 585
R2012 GND.n3378 GND.n3377 585
R2013 GND.n4369 GND.n3378 585
R2014 GND.n4367 GND.n4366 585
R2015 GND.n4368 GND.n4367 585
R2016 GND.n4365 GND.n3380 585
R2017 GND.n3380 GND.n3379 585
R2018 GND.n4364 GND.n4363 585
R2019 GND.n4363 GND.n4362 585
R2020 GND.n3386 GND.n3385 585
R2021 GND.n4361 GND.n3386 585
R2022 GND.n4359 GND.n4358 585
R2023 GND.n4360 GND.n4359 585
R2024 GND.n4357 GND.n3388 585
R2025 GND.n3388 GND.n3387 585
R2026 GND.n4356 GND.n4355 585
R2027 GND.n4355 GND.n4354 585
R2028 GND.n3394 GND.n3393 585
R2029 GND.n4353 GND.n3394 585
R2030 GND.n4351 GND.n4350 585
R2031 GND.n4352 GND.n4351 585
R2032 GND.n4349 GND.n3396 585
R2033 GND.n3396 GND.n3395 585
R2034 GND.n4348 GND.n4347 585
R2035 GND.n4347 GND.n4346 585
R2036 GND.n3402 GND.n3401 585
R2037 GND.n4345 GND.n3402 585
R2038 GND.n4343 GND.n4342 585
R2039 GND.n4344 GND.n4343 585
R2040 GND.n4341 GND.n3404 585
R2041 GND.n3404 GND.n3403 585
R2042 GND.n4340 GND.n4339 585
R2043 GND.n4339 GND.n4338 585
R2044 GND.n3410 GND.n3409 585
R2045 GND.n4337 GND.n3410 585
R2046 GND.n4335 GND.n4334 585
R2047 GND.n4336 GND.n4335 585
R2048 GND.n4333 GND.n3412 585
R2049 GND.n3412 GND.n3411 585
R2050 GND.n4332 GND.n4331 585
R2051 GND.n4331 GND.n4330 585
R2052 GND.n3418 GND.n3417 585
R2053 GND.n4329 GND.n3418 585
R2054 GND.n4327 GND.n4326 585
R2055 GND.n4328 GND.n4327 585
R2056 GND.n4325 GND.n3420 585
R2057 GND.n3420 GND.n3419 585
R2058 GND.n4324 GND.n4323 585
R2059 GND.n4323 GND.n4322 585
R2060 GND.n3426 GND.n3425 585
R2061 GND.n4321 GND.n3426 585
R2062 GND.n4319 GND.n4318 585
R2063 GND.n4320 GND.n4319 585
R2064 GND.n4317 GND.n3428 585
R2065 GND.n3428 GND.n3427 585
R2066 GND.n4316 GND.n4315 585
R2067 GND.n4315 GND.n4314 585
R2068 GND.n3434 GND.n3433 585
R2069 GND.n4313 GND.n3434 585
R2070 GND.n4311 GND.n4310 585
R2071 GND.n4312 GND.n4311 585
R2072 GND.n4309 GND.n3436 585
R2073 GND.n3436 GND.n3435 585
R2074 GND.n4308 GND.n4307 585
R2075 GND.n4307 GND.n4306 585
R2076 GND.n3442 GND.n3441 585
R2077 GND.n4305 GND.n3442 585
R2078 GND.n4303 GND.n4302 585
R2079 GND.n4304 GND.n4303 585
R2080 GND.n4301 GND.n3444 585
R2081 GND.n3444 GND.n3443 585
R2082 GND.n4300 GND.n4299 585
R2083 GND.n4299 GND.n4298 585
R2084 GND.n3450 GND.n3449 585
R2085 GND.n4297 GND.n3450 585
R2086 GND.n4295 GND.n4294 585
R2087 GND.n4296 GND.n4295 585
R2088 GND.n4293 GND.n3452 585
R2089 GND.n3452 GND.n3451 585
R2090 GND.n4292 GND.n4291 585
R2091 GND.n4291 GND.n4290 585
R2092 GND.n3458 GND.n3457 585
R2093 GND.n4289 GND.n3458 585
R2094 GND.n4287 GND.n4286 585
R2095 GND.n4288 GND.n4287 585
R2096 GND.n4285 GND.n3460 585
R2097 GND.n3460 GND.n3459 585
R2098 GND.n4284 GND.n4283 585
R2099 GND.n4283 GND.n4282 585
R2100 GND.n3466 GND.n3465 585
R2101 GND.n4281 GND.n3466 585
R2102 GND.n4279 GND.n4278 585
R2103 GND.n4280 GND.n4279 585
R2104 GND.n4277 GND.n3468 585
R2105 GND.n3468 GND.n3467 585
R2106 GND.n4276 GND.n4275 585
R2107 GND.n4275 GND.n4274 585
R2108 GND.n3474 GND.n3473 585
R2109 GND.n4273 GND.n3474 585
R2110 GND.n4271 GND.n4270 585
R2111 GND.n4272 GND.n4271 585
R2112 GND.n4269 GND.n3476 585
R2113 GND.n3476 GND.n3475 585
R2114 GND.n4268 GND.n4267 585
R2115 GND.n4267 GND.n4266 585
R2116 GND.n3482 GND.n3481 585
R2117 GND.n4265 GND.n3482 585
R2118 GND.n4263 GND.n4262 585
R2119 GND.n4264 GND.n4263 585
R2120 GND.n4261 GND.n3484 585
R2121 GND.n3484 GND.n3483 585
R2122 GND.n4260 GND.n4259 585
R2123 GND.n4259 GND.n4258 585
R2124 GND.n3490 GND.n3489 585
R2125 GND.n4257 GND.n3490 585
R2126 GND.n4255 GND.n4254 585
R2127 GND.n4256 GND.n4255 585
R2128 GND.n4253 GND.n3492 585
R2129 GND.n3492 GND.n3491 585
R2130 GND.n4252 GND.n4251 585
R2131 GND.n4251 GND.n4250 585
R2132 GND.n3498 GND.n3497 585
R2133 GND.n4249 GND.n3498 585
R2134 GND.n4247 GND.n4246 585
R2135 GND.n4248 GND.n4247 585
R2136 GND.n4245 GND.n3500 585
R2137 GND.n3500 GND.n3499 585
R2138 GND.n4244 GND.n4243 585
R2139 GND.n4243 GND.n4242 585
R2140 GND.n3506 GND.n3505 585
R2141 GND.n4241 GND.n3506 585
R2142 GND.n4239 GND.n4238 585
R2143 GND.n4240 GND.n4239 585
R2144 GND.n4237 GND.n3508 585
R2145 GND.n3508 GND.n3507 585
R2146 GND.n4236 GND.n4235 585
R2147 GND.n4235 GND.n4234 585
R2148 GND.n3514 GND.n3513 585
R2149 GND.n4233 GND.n3514 585
R2150 GND.n4231 GND.n4230 585
R2151 GND.n4232 GND.n4231 585
R2152 GND.n4229 GND.n3516 585
R2153 GND.n3516 GND.n3515 585
R2154 GND.n4228 GND.n4227 585
R2155 GND.n4227 GND.n4226 585
R2156 GND.n3522 GND.n3521 585
R2157 GND.n4225 GND.n3522 585
R2158 GND.n4223 GND.n4222 585
R2159 GND.n4224 GND.n4223 585
R2160 GND.n4221 GND.n3524 585
R2161 GND.n3524 GND.n3523 585
R2162 GND.n4220 GND.n4219 585
R2163 GND.n4219 GND.n4218 585
R2164 GND.n3530 GND.n3529 585
R2165 GND.n4217 GND.n3530 585
R2166 GND.n4215 GND.n4214 585
R2167 GND.n4216 GND.n4215 585
R2168 GND.n4213 GND.n3532 585
R2169 GND.n3532 GND.n3531 585
R2170 GND.n4212 GND.n4211 585
R2171 GND.n4211 GND.n4210 585
R2172 GND.n3538 GND.n3537 585
R2173 GND.n4209 GND.n3538 585
R2174 GND.n4207 GND.n4206 585
R2175 GND.n4208 GND.n4207 585
R2176 GND.n4205 GND.n3540 585
R2177 GND.n3540 GND.n3539 585
R2178 GND.n4204 GND.n4203 585
R2179 GND.n4203 GND.n4202 585
R2180 GND.n3546 GND.n3545 585
R2181 GND.n4201 GND.n3546 585
R2182 GND.n4199 GND.n4198 585
R2183 GND.n4200 GND.n4199 585
R2184 GND.n4197 GND.n3548 585
R2185 GND.n3548 GND.n3547 585
R2186 GND.n4196 GND.n4195 585
R2187 GND.n4195 GND.n4194 585
R2188 GND.n3554 GND.n3553 585
R2189 GND.n4193 GND.n3554 585
R2190 GND.n4191 GND.n4190 585
R2191 GND.n4192 GND.n4191 585
R2192 GND.n4189 GND.n3556 585
R2193 GND.n3556 GND.n3555 585
R2194 GND.n4188 GND.n4187 585
R2195 GND.n4187 GND.n4186 585
R2196 GND.n3562 GND.n3561 585
R2197 GND.n4185 GND.n3562 585
R2198 GND.n4183 GND.n4182 585
R2199 GND.n4184 GND.n4183 585
R2200 GND.n4181 GND.n3564 585
R2201 GND.n3564 GND.n3563 585
R2202 GND.n4180 GND.n4179 585
R2203 GND.n4179 GND.n4178 585
R2204 GND.n3570 GND.n3569 585
R2205 GND.n4177 GND.n3570 585
R2206 GND.n4175 GND.n4174 585
R2207 GND.n4176 GND.n4175 585
R2208 GND.n4173 GND.n3572 585
R2209 GND.n3572 GND.n3571 585
R2210 GND.n4172 GND.n4171 585
R2211 GND.n4171 GND.n4170 585
R2212 GND.n3578 GND.n3577 585
R2213 GND.n4169 GND.n3578 585
R2214 GND.n4167 GND.n4166 585
R2215 GND.n4168 GND.n4167 585
R2216 GND.n4165 GND.n3580 585
R2217 GND.n3580 GND.n3579 585
R2218 GND.n4164 GND.n4163 585
R2219 GND.n4163 GND.n4162 585
R2220 GND.n3586 GND.n3585 585
R2221 GND.n4161 GND.n3586 585
R2222 GND.n4159 GND.n4158 585
R2223 GND.n4160 GND.n4159 585
R2224 GND.n4157 GND.n3588 585
R2225 GND.n3588 GND.n3587 585
R2226 GND.n4156 GND.n4155 585
R2227 GND.n4155 GND.n4154 585
R2228 GND.n3594 GND.n3593 585
R2229 GND.n4153 GND.n3594 585
R2230 GND.n4151 GND.n4150 585
R2231 GND.n4152 GND.n4151 585
R2232 GND.n4149 GND.n3596 585
R2233 GND.n3596 GND.n3595 585
R2234 GND.n4148 GND.n4147 585
R2235 GND.n4147 GND.n4146 585
R2236 GND.n3602 GND.n3601 585
R2237 GND.n4145 GND.n3602 585
R2238 GND.n4143 GND.n4142 585
R2239 GND.n4144 GND.n4143 585
R2240 GND.n4141 GND.n3604 585
R2241 GND.n3604 GND.n3603 585
R2242 GND.n4140 GND.n4139 585
R2243 GND.n4139 GND.n4138 585
R2244 GND.n3610 GND.n3609 585
R2245 GND.n4137 GND.n3610 585
R2246 GND.n4135 GND.n4134 585
R2247 GND.n4136 GND.n4135 585
R2248 GND.n4133 GND.n3612 585
R2249 GND.n3612 GND.n3611 585
R2250 GND.n4132 GND.n4131 585
R2251 GND.n4131 GND.n4130 585
R2252 GND.n3618 GND.n3617 585
R2253 GND.n4129 GND.n3618 585
R2254 GND.n4127 GND.n4126 585
R2255 GND.n4128 GND.n4127 585
R2256 GND.n4125 GND.n3620 585
R2257 GND.n3620 GND.n3619 585
R2258 GND.n4124 GND.n4123 585
R2259 GND.n4123 GND.n4122 585
R2260 GND.n3626 GND.n3625 585
R2261 GND.n4121 GND.n3626 585
R2262 GND.n4119 GND.n4118 585
R2263 GND.n4120 GND.n4119 585
R2264 GND.n4117 GND.n3628 585
R2265 GND.n3628 GND.n3627 585
R2266 GND.n4116 GND.n4115 585
R2267 GND.n4115 GND.n4114 585
R2268 GND.n3634 GND.n3633 585
R2269 GND.n4113 GND.n3634 585
R2270 GND.n4111 GND.n4110 585
R2271 GND.n4112 GND.n4111 585
R2272 GND.n4109 GND.n3636 585
R2273 GND.n3636 GND.n3635 585
R2274 GND.n4108 GND.n4107 585
R2275 GND.n4107 GND.n4106 585
R2276 GND.n3642 GND.n3641 585
R2277 GND.n4105 GND.n3642 585
R2278 GND.n4103 GND.n4102 585
R2279 GND.n4104 GND.n4103 585
R2280 GND.n4101 GND.n3644 585
R2281 GND.n3644 GND.n3643 585
R2282 GND.n4100 GND.n4099 585
R2283 GND.n4099 GND.n4098 585
R2284 GND.n3650 GND.n3649 585
R2285 GND.n4097 GND.n3650 585
R2286 GND.n4095 GND.n4094 585
R2287 GND.n4096 GND.n4095 585
R2288 GND.n4093 GND.n3652 585
R2289 GND.n3652 GND.n3651 585
R2290 GND.n4092 GND.n4091 585
R2291 GND.n4091 GND.n4090 585
R2292 GND.n3658 GND.n3657 585
R2293 GND.n4089 GND.n3658 585
R2294 GND.n4087 GND.n4086 585
R2295 GND.n4088 GND.n4087 585
R2296 GND.n4085 GND.n3660 585
R2297 GND.n3660 GND.n3659 585
R2298 GND.n4084 GND.n4083 585
R2299 GND.n4083 GND.n4082 585
R2300 GND.n3666 GND.n3665 585
R2301 GND.n4081 GND.n3666 585
R2302 GND.n4079 GND.n4078 585
R2303 GND.n4080 GND.n4079 585
R2304 GND.n4077 GND.n3668 585
R2305 GND.n3668 GND.n3667 585
R2306 GND.n4076 GND.n4075 585
R2307 GND.n4075 GND.n4074 585
R2308 GND.n3674 GND.n3673 585
R2309 GND.n4073 GND.n3674 585
R2310 GND.n4071 GND.n4070 585
R2311 GND.n4072 GND.n4071 585
R2312 GND.n4069 GND.n3676 585
R2313 GND.n3676 GND.n3675 585
R2314 GND.n4068 GND.n4067 585
R2315 GND.n4067 GND.n4066 585
R2316 GND.n3682 GND.n3681 585
R2317 GND.n4065 GND.n3682 585
R2318 GND.n4063 GND.n4062 585
R2319 GND.n4064 GND.n4063 585
R2320 GND.n4061 GND.n3684 585
R2321 GND.n3684 GND.n3683 585
R2322 GND.n4060 GND.n4059 585
R2323 GND.n4059 GND.n4058 585
R2324 GND.n3690 GND.n3689 585
R2325 GND.n4057 GND.n3690 585
R2326 GND.n4055 GND.n4054 585
R2327 GND.n4056 GND.n4055 585
R2328 GND.n4053 GND.n3692 585
R2329 GND.n3692 GND.n3691 585
R2330 GND.n4052 GND.n4051 585
R2331 GND.n4051 GND.n4050 585
R2332 GND.n3698 GND.n3697 585
R2333 GND.n4049 GND.n3698 585
R2334 GND.n4047 GND.n4046 585
R2335 GND.n4048 GND.n4047 585
R2336 GND.n4045 GND.n3700 585
R2337 GND.n3700 GND.n3699 585
R2338 GND.n4044 GND.n4043 585
R2339 GND.n4043 GND.n4042 585
R2340 GND.n3706 GND.n3705 585
R2341 GND.n4041 GND.n3706 585
R2342 GND.n4039 GND.n4038 585
R2343 GND.n4040 GND.n4039 585
R2344 GND.n4037 GND.n3708 585
R2345 GND.n3708 GND.n3707 585
R2346 GND.n4036 GND.n4035 585
R2347 GND.n4035 GND.n4034 585
R2348 GND.n3714 GND.n3713 585
R2349 GND.n4033 GND.n3714 585
R2350 GND.n4031 GND.n4030 585
R2351 GND.n4032 GND.n4031 585
R2352 GND.n4029 GND.n3716 585
R2353 GND.n3716 GND.n3715 585
R2354 GND.n4028 GND.n4027 585
R2355 GND.n4027 GND.n4026 585
R2356 GND.n3722 GND.n3721 585
R2357 GND.n4025 GND.n3722 585
R2358 GND.n4023 GND.n4022 585
R2359 GND.n4024 GND.n4023 585
R2360 GND.n4021 GND.n3724 585
R2361 GND.n3724 GND.n3723 585
R2362 GND.n4020 GND.n4019 585
R2363 GND.n4019 GND.n4018 585
R2364 GND.n3730 GND.n3729 585
R2365 GND.n4017 GND.n3730 585
R2366 GND.n4015 GND.n4014 585
R2367 GND.n4016 GND.n4015 585
R2368 GND.n4013 GND.n3732 585
R2369 GND.n3732 GND.n3731 585
R2370 GND.n4012 GND.n4011 585
R2371 GND.n4011 GND.n4010 585
R2372 GND.n3738 GND.n3737 585
R2373 GND.n4009 GND.n3738 585
R2374 GND.n4007 GND.n4006 585
R2375 GND.n4008 GND.n4007 585
R2376 GND.n4005 GND.n3740 585
R2377 GND.n3740 GND.n3739 585
R2378 GND.n4004 GND.n4003 585
R2379 GND.n4003 GND.n4002 585
R2380 GND.n3746 GND.n3745 585
R2381 GND.n4001 GND.n3746 585
R2382 GND.n3999 GND.n3998 585
R2383 GND.n4000 GND.n3999 585
R2384 GND.n3997 GND.n3748 585
R2385 GND.n3748 GND.n3747 585
R2386 GND.n3996 GND.n3995 585
R2387 GND.n3995 GND.n3994 585
R2388 GND.n3754 GND.n3753 585
R2389 GND.n3993 GND.n3754 585
R2390 GND.n3991 GND.n3990 585
R2391 GND.n3992 GND.n3991 585
R2392 GND.n3989 GND.n3756 585
R2393 GND.n3756 GND.n3755 585
R2394 GND.n3988 GND.n3987 585
R2395 GND.n3987 GND.n3986 585
R2396 GND.n3762 GND.n3761 585
R2397 GND.n3985 GND.n3762 585
R2398 GND.n3983 GND.n3982 585
R2399 GND.n3984 GND.n3983 585
R2400 GND.n3981 GND.n3764 585
R2401 GND.n3764 GND.n3763 585
R2402 GND.n3980 GND.n3979 585
R2403 GND.n3979 GND.n3978 585
R2404 GND.n3770 GND.n3769 585
R2405 GND.n3977 GND.n3770 585
R2406 GND.n3975 GND.n3974 585
R2407 GND.n3976 GND.n3975 585
R2408 GND.n3973 GND.n3772 585
R2409 GND.n3772 GND.n3771 585
R2410 GND.n3972 GND.n3971 585
R2411 GND.n3971 GND.n3970 585
R2412 GND.n3778 GND.n3777 585
R2413 GND.n3969 GND.n3778 585
R2414 GND.n3967 GND.n3966 585
R2415 GND.n3968 GND.n3967 585
R2416 GND.n3965 GND.n3780 585
R2417 GND.n3780 GND.n3779 585
R2418 GND.n8453 GND.n344 585
R2419 GND.n8449 GND.n344 585
R2420 GND.n8452 GND.n8451 585
R2421 GND.n8451 GND.n8450 585
R2422 GND.n348 GND.n347 585
R2423 GND.n349 GND.n348 585
R2424 GND.n3874 GND.n3873 585
R2425 GND.n3873 GND.n3872 585
R2426 GND.n3875 GND.n3866 585
R2427 GND.n3866 GND.n3865 585
R2428 GND.n3877 GND.n3876 585
R2429 GND.n3878 GND.n3877 585
R2430 GND.n3864 GND.n3863 585
R2431 GND.n3879 GND.n3864 585
R2432 GND.n3882 GND.n3881 585
R2433 GND.n3881 GND.n3880 585
R2434 GND.n3883 GND.n3858 585
R2435 GND.n3858 GND.n3857 585
R2436 GND.n3885 GND.n3884 585
R2437 GND.n3886 GND.n3885 585
R2438 GND.n3856 GND.n3855 585
R2439 GND.n3887 GND.n3856 585
R2440 GND.n3890 GND.n3889 585
R2441 GND.n3889 GND.n3888 585
R2442 GND.n3891 GND.n3850 585
R2443 GND.n3850 GND.n3849 585
R2444 GND.n3893 GND.n3892 585
R2445 GND.n3894 GND.n3893 585
R2446 GND.n3848 GND.n3847 585
R2447 GND.n3895 GND.n3848 585
R2448 GND.n3898 GND.n3897 585
R2449 GND.n3897 GND.n3896 585
R2450 GND.n3899 GND.n3842 585
R2451 GND.n3842 GND.n3841 585
R2452 GND.n3901 GND.n3900 585
R2453 GND.n3902 GND.n3901 585
R2454 GND.n3840 GND.n3839 585
R2455 GND.n3903 GND.n3840 585
R2456 GND.n3906 GND.n3905 585
R2457 GND.n3905 GND.n3904 585
R2458 GND.n3907 GND.n3834 585
R2459 GND.n3834 GND.n3833 585
R2460 GND.n3909 GND.n3908 585
R2461 GND.n3910 GND.n3909 585
R2462 GND.n3832 GND.n3831 585
R2463 GND.n3911 GND.n3832 585
R2464 GND.n3914 GND.n3913 585
R2465 GND.n3913 GND.n3912 585
R2466 GND.n3915 GND.n3826 585
R2467 GND.n3826 GND.n3825 585
R2468 GND.n3917 GND.n3916 585
R2469 GND.n3918 GND.n3917 585
R2470 GND.n3824 GND.n3823 585
R2471 GND.n3919 GND.n3824 585
R2472 GND.n3922 GND.n3921 585
R2473 GND.n3921 GND.n3920 585
R2474 GND.n3923 GND.n3818 585
R2475 GND.n3818 GND.n3817 585
R2476 GND.n3925 GND.n3924 585
R2477 GND.n3926 GND.n3925 585
R2478 GND.n3816 GND.n3815 585
R2479 GND.n3927 GND.n3816 585
R2480 GND.n3930 GND.n3929 585
R2481 GND.n3929 GND.n3928 585
R2482 GND.n3931 GND.n3810 585
R2483 GND.n3810 GND.n3809 585
R2484 GND.n3933 GND.n3932 585
R2485 GND.n3934 GND.n3933 585
R2486 GND.n3808 GND.n3807 585
R2487 GND.n3935 GND.n3808 585
R2488 GND.n3938 GND.n3937 585
R2489 GND.n3937 GND.n3936 585
R2490 GND.n3939 GND.n3802 585
R2491 GND.n3802 GND.n3801 585
R2492 GND.n3941 GND.n3940 585
R2493 GND.n3942 GND.n3941 585
R2494 GND.n3800 GND.n3799 585
R2495 GND.n3943 GND.n3800 585
R2496 GND.n3946 GND.n3945 585
R2497 GND.n3945 GND.n3944 585
R2498 GND.n3947 GND.n3794 585
R2499 GND.n3794 GND.n3793 585
R2500 GND.n3949 GND.n3948 585
R2501 GND.n3950 GND.n3949 585
R2502 GND.n3792 GND.n3791 585
R2503 GND.n3951 GND.n3792 585
R2504 GND.n3954 GND.n3953 585
R2505 GND.n3953 GND.n3952 585
R2506 GND.n3955 GND.n3787 585
R2507 GND.n3787 GND.n3786 585
R2508 GND.n3957 GND.n3956 585
R2509 GND.n3958 GND.n3957 585
R2510 GND.n3785 GND.n3784 585
R2511 GND.n3959 GND.n3785 585
R2512 GND.n3962 GND.n3961 585
R2513 GND.n3961 GND.n3960 585
R2514 GND.n451 GND.n446 585
R2515 GND.n451 GND.n350 585
R2516 GND.n8312 GND.n452 585
R2517 GND.n8326 GND.n452 585
R2518 GND.n8313 GND.n8224 585
R2519 GND.n8224 GND.n449 585
R2520 GND.n8315 GND.n8314 585
R2521 GND.n8316 GND.n8315 585
R2522 GND.n8225 GND.n8223 585
R2523 GND.n8223 GND.n8069 585
R2524 GND.n8304 GND.n8303 585
R2525 GND.n8303 GND.n342 585
R2526 GND.n8302 GND.n341 585
R2527 GND.n8458 GND.n341 585
R2528 GND.n8301 GND.n8300 585
R2529 GND.n8300 GND.n332 585
R2530 GND.n8299 GND.n331 585
R2531 GND.n8464 GND.n331 585
R2532 GND.n8298 GND.n8297 585
R2533 GND.n8297 GND.n321 585
R2534 GND.n8295 GND.n320 585
R2535 GND.n8470 GND.n320 585
R2536 GND.n8294 GND.n8293 585
R2537 GND.n8293 GND.n311 585
R2538 GND.n8292 GND.n310 585
R2539 GND.n8476 GND.n310 585
R2540 GND.n8291 GND.n8290 585
R2541 GND.n8290 GND.n300 585
R2542 GND.n8288 GND.n299 585
R2543 GND.n8482 GND.n299 585
R2544 GND.n8287 GND.n8286 585
R2545 GND.n8286 GND.n290 585
R2546 GND.n8285 GND.n289 585
R2547 GND.n8488 GND.n289 585
R2548 GND.n8284 GND.n8283 585
R2549 GND.n8283 GND.n279 585
R2550 GND.n8281 GND.n278 585
R2551 GND.n8494 GND.n278 585
R2552 GND.n8280 GND.n8279 585
R2553 GND.n8279 GND.n269 585
R2554 GND.n8278 GND.n268 585
R2555 GND.n8500 GND.n268 585
R2556 GND.n8277 GND.n8276 585
R2557 GND.n8276 GND.n258 585
R2558 GND.n8274 GND.n257 585
R2559 GND.n8506 GND.n257 585
R2560 GND.n8273 GND.n8272 585
R2561 GND.n8272 GND.n248 585
R2562 GND.n8271 GND.n247 585
R2563 GND.n8512 GND.n247 585
R2564 GND.n8270 GND.n8269 585
R2565 GND.n8269 GND.n237 585
R2566 GND.n8267 GND.n236 585
R2567 GND.n8518 GND.n236 585
R2568 GND.n8266 GND.n8265 585
R2569 GND.n8265 GND.n227 585
R2570 GND.n8264 GND.n226 585
R2571 GND.n8524 GND.n226 585
R2572 GND.n8263 GND.n8262 585
R2573 GND.n8262 GND.n216 585
R2574 GND.n8260 GND.n215 585
R2575 GND.n8530 GND.n215 585
R2576 GND.n8259 GND.n8258 585
R2577 GND.n8258 GND.n206 585
R2578 GND.n8257 GND.n205 585
R2579 GND.n8536 GND.n205 585
R2580 GND.n8256 GND.n8255 585
R2581 GND.n8255 GND.n195 585
R2582 GND.n8253 GND.n194 585
R2583 GND.n8542 GND.n194 585
R2584 GND.n8252 GND.n8251 585
R2585 GND.n8251 GND.n192 585
R2586 GND.n8250 GND.n184 585
R2587 GND.n8548 GND.n184 585
R2588 GND.n8249 GND.n8248 585
R2589 GND.n8248 GND.n174 585
R2590 GND.n8246 GND.n173 585
R2591 GND.n8554 GND.n173 585
R2592 GND.n8245 GND.n8244 585
R2593 GND.n8244 GND.n164 585
R2594 GND.n8243 GND.n163 585
R2595 GND.n8560 GND.n163 585
R2596 GND.n8242 GND.n8241 585
R2597 GND.n8241 GND.n154 585
R2598 GND.n8239 GND.n153 585
R2599 GND.n8566 GND.n153 585
R2600 GND.n8238 GND.n8237 585
R2601 GND.n8237 GND.n142 585
R2602 GND.n8236 GND.n141 585
R2603 GND.n8572 GND.n141 585
R2604 GND.n8235 GND.n134 585
R2605 GND.n136 GND.n134 585
R2606 GND.n8580 GND.n133 585
R2607 GND.n8580 GND.n8579 585
R2608 GND.n8582 GND.n8581 585
R2609 GND.n8581 GND.n71 585
R2610 GND.n8583 GND.n72 585
R2611 GND.t25 GND.n72 585
R2612 GND.n8585 GND.n8584 585
R2613 GND.n8585 GND.n68 585
R2614 GND.n8587 GND.n8586 585
R2615 GND.n8586 GND.n103 585
R2616 GND.n8588 GND.n102 585
R2617 GND.n8624 GND.n102 585
R2618 GND.n8590 GND.n8589 585
R2619 GND.n8589 GND.n91 585
R2620 GND.n8591 GND.n90 585
R2621 GND.n8630 GND.n90 585
R2622 GND.n8593 GND.n8592 585
R2623 GND.n8592 GND.n88 585
R2624 GND.n128 GND.n112 585
R2625 GND.n8608 GND.n112 585
R2626 GND.n7939 GND.n7938 585
R2627 GND.n7938 GND.n110 585
R2628 GND.n7940 GND.n121 585
R2629 GND.n8600 GND.n121 585
R2630 GND.n7942 GND.n7941 585
R2631 GND.n7941 GND.n119 585
R2632 GND.n7937 GND.n481 585
R2633 GND.n7957 GND.n481 585
R2634 GND.n7936 GND.n7935 585
R2635 GND.n7935 GND.n480 585
R2636 GND.n7934 GND.n491 585
R2637 GND.n7949 GND.n491 585
R2638 GND.n7933 GND.n7932 585
R2639 GND.n7932 GND.n489 585
R2640 GND.n7931 GND.n498 585
R2641 GND.n7931 GND.n7930 585
R2642 GND.n7915 GND.n500 585
R2643 GND.n501 GND.n500 585
R2644 GND.n7914 GND.n512 585
R2645 GND.n7922 GND.n512 585
R2646 GND.n7913 GND.n7912 585
R2647 GND.n7912 GND.n510 585
R2648 GND.n7911 GND.n518 585
R2649 GND.n7911 GND.n7910 585
R2650 GND.n7895 GND.n520 585
R2651 GND.n521 GND.n520 585
R2652 GND.n7894 GND.n532 585
R2653 GND.n7902 GND.n532 585
R2654 GND.n7893 GND.n7892 585
R2655 GND.n7892 GND.n530 585
R2656 GND.n7891 GND.n538 585
R2657 GND.n7891 GND.n7890 585
R2658 GND.n7875 GND.n540 585
R2659 GND.n541 GND.n540 585
R2660 GND.n7874 GND.n551 585
R2661 GND.n7882 GND.n551 585
R2662 GND.n7873 GND.n7872 585
R2663 GND.n7872 GND.n7871 585
R2664 GND.n559 GND.n557 585
R2665 GND.n560 GND.n559 585
R2666 GND.n7799 GND.n569 585
R2667 GND.n7818 GND.n569 585
R2668 GND.n7798 GND.n7797 585
R2669 GND.n7797 GND.n567 585
R2670 GND.n7796 GND.n579 585
R2671 GND.n7808 GND.n579 585
R2672 GND.n7795 GND.n7794 585
R2673 GND.n7794 GND.n577 585
R2674 GND.n7793 GND.n586 585
R2675 GND.n7793 GND.n7792 585
R2676 GND.n7777 GND.n588 585
R2677 GND.n589 GND.n588 585
R2678 GND.n7776 GND.n600 585
R2679 GND.n7784 GND.n600 585
R2680 GND.n7775 GND.n7774 585
R2681 GND.n7774 GND.n598 585
R2682 GND.n7773 GND.n606 585
R2683 GND.n7773 GND.n7772 585
R2684 GND.n7757 GND.n608 585
R2685 GND.n609 GND.n608 585
R2686 GND.n7756 GND.n620 585
R2687 GND.n7764 GND.n620 585
R2688 GND.n7755 GND.n7754 585
R2689 GND.n7754 GND.n618 585
R2690 GND.n7753 GND.n626 585
R2691 GND.n7753 GND.n7752 585
R2692 GND.n7737 GND.n628 585
R2693 GND.n629 GND.n628 585
R2694 GND.n7736 GND.n640 585
R2695 GND.n7744 GND.n640 585
R2696 GND.n7735 GND.n7734 585
R2697 GND.n7734 GND.n638 585
R2698 GND.n7733 GND.n646 585
R2699 GND.n7733 GND.n7732 585
R2700 GND.n7717 GND.n648 585
R2701 GND.n649 GND.n648 585
R2702 GND.n7716 GND.n660 585
R2703 GND.n7724 GND.n660 585
R2704 GND.n7715 GND.n667 585
R2705 GND.n667 GND.n658 585
R2706 GND.n672 GND.n666 585
R2707 GND.n7710 GND.n672 585
R2708 GND.n1226 GND.n1225 585
R2709 GND.n1224 GND.n1223 585
R2710 GND.n1222 GND.n1221 585
R2711 GND.n1220 GND.n1219 585
R2712 GND.n1218 GND.n1217 585
R2713 GND.n1216 GND.n1215 585
R2714 GND.n1214 GND.n1213 585
R2715 GND.n1212 GND.n1211 585
R2716 GND.n1210 GND.n1209 585
R2717 GND.n1208 GND.n1205 585
R2718 GND.n7701 GND.n711 585
R2719 GND.n8216 GND.n8215 585
R2720 GND.n8209 GND.n8186 585
R2721 GND.n8211 GND.n8210 585
R2722 GND.n8208 GND.n8207 585
R2723 GND.n8206 GND.n8205 585
R2724 GND.n8199 GND.n8188 585
R2725 GND.n8201 GND.n8200 585
R2726 GND.n8198 GND.n8197 585
R2727 GND.n8196 GND.n8195 585
R2728 GND.n8192 GND.n8191 585
R2729 GND.n8190 GND.n351 585
R2730 GND.n8448 GND.n351 585
R2731 GND.n8218 GND.n8217 585
R2732 GND.n8217 GND.n350 585
R2733 GND.n8219 GND.n450 585
R2734 GND.n8326 GND.n450 585
R2735 GND.n8220 GND.n8072 585
R2736 GND.n8072 GND.n449 585
R2737 GND.n8222 GND.n8221 585
R2738 GND.n8316 GND.n8222 585
R2739 GND.n8073 GND.n8071 585
R2740 GND.n8071 GND.n8069 585
R2741 GND.n8177 GND.n8176 585
R2742 GND.n8176 GND.n342 585
R2743 GND.n8175 GND.n343 585
R2744 GND.n8458 GND.n343 585
R2745 GND.n8174 GND.n8173 585
R2746 GND.n8173 GND.n332 585
R2747 GND.n8075 GND.n333 585
R2748 GND.n8464 GND.n333 585
R2749 GND.n8169 GND.n8168 585
R2750 GND.n8168 GND.n321 585
R2751 GND.n8167 GND.n322 585
R2752 GND.n8470 GND.n322 585
R2753 GND.n8166 GND.n8165 585
R2754 GND.n8165 GND.n311 585
R2755 GND.n8077 GND.n312 585
R2756 GND.n8476 GND.n312 585
R2757 GND.n8161 GND.n8160 585
R2758 GND.n8160 GND.n300 585
R2759 GND.n8159 GND.n301 585
R2760 GND.n8482 GND.n301 585
R2761 GND.n8158 GND.n8157 585
R2762 GND.n8157 GND.n290 585
R2763 GND.n8079 GND.n291 585
R2764 GND.n8488 GND.n291 585
R2765 GND.n8153 GND.n8152 585
R2766 GND.n8152 GND.n279 585
R2767 GND.n8151 GND.n280 585
R2768 GND.n8494 GND.n280 585
R2769 GND.n8150 GND.n8149 585
R2770 GND.n8149 GND.n269 585
R2771 GND.n8081 GND.n270 585
R2772 GND.n8500 GND.n270 585
R2773 GND.n8145 GND.n8144 585
R2774 GND.n8144 GND.n258 585
R2775 GND.n8143 GND.n259 585
R2776 GND.n8506 GND.n259 585
R2777 GND.n8142 GND.n8141 585
R2778 GND.n8141 GND.n248 585
R2779 GND.n8083 GND.n249 585
R2780 GND.n8512 GND.n249 585
R2781 GND.n8137 GND.n8136 585
R2782 GND.n8136 GND.n237 585
R2783 GND.n8135 GND.n238 585
R2784 GND.n8518 GND.n238 585
R2785 GND.n8134 GND.n8133 585
R2786 GND.n8133 GND.n227 585
R2787 GND.n8085 GND.n228 585
R2788 GND.n8524 GND.n228 585
R2789 GND.n8129 GND.n8128 585
R2790 GND.n8128 GND.n216 585
R2791 GND.n8127 GND.n217 585
R2792 GND.n8530 GND.n217 585
R2793 GND.n8126 GND.n8125 585
R2794 GND.n8125 GND.n206 585
R2795 GND.n8087 GND.n207 585
R2796 GND.n8536 GND.n207 585
R2797 GND.n8121 GND.n8120 585
R2798 GND.n8120 GND.n195 585
R2799 GND.n8119 GND.n196 585
R2800 GND.n8542 GND.n196 585
R2801 GND.n8118 GND.n8117 585
R2802 GND.n8117 GND.n192 585
R2803 GND.n8089 GND.n185 585
R2804 GND.n8548 GND.n185 585
R2805 GND.n8113 GND.n8112 585
R2806 GND.n8112 GND.n174 585
R2807 GND.n8111 GND.n175 585
R2808 GND.n8554 GND.n175 585
R2809 GND.n8110 GND.n8109 585
R2810 GND.n8109 GND.n164 585
R2811 GND.n8091 GND.n165 585
R2812 GND.n8560 GND.n165 585
R2813 GND.n8105 GND.n8104 585
R2814 GND.n8104 GND.n154 585
R2815 GND.n8103 GND.n155 585
R2816 GND.n8566 GND.n155 585
R2817 GND.n8102 GND.n8101 585
R2818 GND.n8101 GND.n142 585
R2819 GND.n8093 GND.n143 585
R2820 GND.n8572 GND.n143 585
R2821 GND.n8097 GND.n8096 585
R2822 GND.n8096 GND.n136 585
R2823 GND.n8095 GND.n137 585
R2824 GND.n8579 GND.n137 585
R2825 GND.n67 GND.n65 585
R2826 GND.n71 GND.n67 585
R2827 GND.n8638 GND.n8637 585
R2828 GND.n8637 GND.t25 585
R2829 GND.n66 GND.n64 585
R2830 GND.n68 GND.n66 585
R2831 GND.n8617 GND.n105 585
R2832 GND.n105 GND.n103 585
R2833 GND.n8619 GND.n8618 585
R2834 GND.n8624 GND.n8619 585
R2835 GND.n106 GND.n104 585
R2836 GND.n104 GND.n91 585
R2837 GND.n8612 GND.n92 585
R2838 GND.n8630 GND.n92 585
R2839 GND.n8611 GND.n8610 585
R2840 GND.n8610 GND.n88 585
R2841 GND.n8609 GND.n108 585
R2842 GND.n8609 GND.n8608 585
R2843 GND.n7843 GND.n109 585
R2844 GND.n110 GND.n109 585
R2845 GND.n7844 GND.n122 585
R2846 GND.n8600 GND.n122 585
R2847 GND.n7846 GND.n7845 585
R2848 GND.n7845 GND.n119 585
R2849 GND.n7847 GND.n482 585
R2850 GND.n7957 GND.n482 585
R2851 GND.n7849 GND.n7848 585
R2852 GND.n7848 GND.n480 585
R2853 GND.n7850 GND.n492 585
R2854 GND.n7949 GND.n492 585
R2855 GND.n7852 GND.n7851 585
R2856 GND.n7851 GND.n489 585
R2857 GND.n7853 GND.n503 585
R2858 GND.n7930 GND.n503 585
R2859 GND.n7855 GND.n7854 585
R2860 GND.n7854 GND.n501 585
R2861 GND.n7856 GND.n513 585
R2862 GND.n7922 GND.n513 585
R2863 GND.n7858 GND.n7857 585
R2864 GND.n7857 GND.n510 585
R2865 GND.n7859 GND.n523 585
R2866 GND.n7910 GND.n523 585
R2867 GND.n7861 GND.n7860 585
R2868 GND.n7860 GND.n521 585
R2869 GND.n7862 GND.n533 585
R2870 GND.n7902 GND.n533 585
R2871 GND.n7864 GND.n7863 585
R2872 GND.n7863 GND.n530 585
R2873 GND.n7865 GND.n543 585
R2874 GND.n7890 GND.n543 585
R2875 GND.n7867 GND.n7866 585
R2876 GND.n7866 GND.n541 585
R2877 GND.n7868 GND.n552 585
R2878 GND.n7882 GND.n552 585
R2879 GND.n7870 GND.n7869 585
R2880 GND.n7871 GND.n7870 585
R2881 GND.n563 GND.n562 585
R2882 GND.n562 GND.n560 585
R2883 GND.n7820 GND.n7819 585
R2884 GND.n7819 GND.n7818 585
R2885 GND.n566 GND.n565 585
R2886 GND.n567 GND.n566 585
R2887 GND.n1246 GND.n580 585
R2888 GND.n7808 GND.n580 585
R2889 GND.n1248 GND.n1247 585
R2890 GND.n1247 GND.n577 585
R2891 GND.n1249 GND.n591 585
R2892 GND.n7792 GND.n591 585
R2893 GND.n1251 GND.n1250 585
R2894 GND.n1250 GND.n589 585
R2895 GND.n1252 GND.n601 585
R2896 GND.n7784 GND.n601 585
R2897 GND.n1254 GND.n1253 585
R2898 GND.n1253 GND.n598 585
R2899 GND.n1255 GND.n611 585
R2900 GND.n7772 GND.n611 585
R2901 GND.n1257 GND.n1256 585
R2902 GND.n1256 GND.n609 585
R2903 GND.n1258 GND.n621 585
R2904 GND.n7764 GND.n621 585
R2905 GND.n1260 GND.n1259 585
R2906 GND.n1259 GND.n618 585
R2907 GND.n1261 GND.n631 585
R2908 GND.n7752 GND.n631 585
R2909 GND.n1263 GND.n1262 585
R2910 GND.n1262 GND.n629 585
R2911 GND.n1264 GND.n641 585
R2912 GND.n7744 GND.n641 585
R2913 GND.n1266 GND.n1265 585
R2914 GND.n1265 GND.n638 585
R2915 GND.n1267 GND.n651 585
R2916 GND.n7732 GND.n651 585
R2917 GND.n1269 GND.n1268 585
R2918 GND.n1268 GND.n649 585
R2919 GND.n1270 GND.n661 585
R2920 GND.n7724 GND.n661 585
R2921 GND.n1271 GND.n1228 585
R2922 GND.n1228 GND.n658 585
R2923 GND.n1272 GND.n673 585
R2924 GND.n7710 GND.n673 585
R2925 GND.n6983 GND.n6982 585
R2926 GND.n6984 GND.n6983 585
R2927 GND.n1178 GND.n1176 585
R2928 GND.n6925 GND.n1176 585
R2929 GND.n6868 GND.n6867 585
R2930 GND.n6867 GND.n1295 585
R2931 GND.n6869 GND.n1323 585
R2932 GND.n6807 GND.n1323 585
R2933 GND.n6871 GND.n6870 585
R2934 GND.n6872 GND.n6871 585
R2935 GND.n1324 GND.n1322 585
R2936 GND.n1322 GND.n1310 585
R2937 GND.n6861 GND.n6860 585
R2938 GND.n6860 GND.n1315 585
R2939 GND.n6859 GND.n1326 585
R2940 GND.n6859 GND.n1314 585
R2941 GND.n6858 GND.n1328 585
R2942 GND.n6858 GND.n6857 585
R2943 GND.n6837 GND.n1327 585
R2944 GND.n6849 GND.n1327 585
R2945 GND.n6839 GND.n6838 585
R2946 GND.n6840 GND.n6839 585
R2947 GND.n1345 GND.n1344 585
R2948 GND.n6821 GND.n1344 585
R2949 GND.n6831 GND.n6830 585
R2950 GND.n6830 GND.n6829 585
R2951 GND.n1348 GND.n1347 585
R2952 GND.n6790 GND.n1348 585
R2953 GND.n6769 GND.n1375 585
R2954 GND.n1375 GND.n1364 585
R2955 GND.n6771 GND.n6770 585
R2956 GND.n6772 GND.n6771 585
R2957 GND.n1376 GND.n1374 585
R2958 GND.t5 GND.n1374 585
R2959 GND.n6764 GND.n6763 585
R2960 GND.n6763 GND.n6762 585
R2961 GND.n1379 GND.n1378 585
R2962 GND.n6754 GND.n1379 585
R2963 GND.n6701 GND.n1406 585
R2964 GND.n1406 GND.n1397 585
R2965 GND.n6703 GND.n6702 585
R2966 GND.n6704 GND.n6703 585
R2967 GND.n1407 GND.n1405 585
R2968 GND.n1405 GND.n1401 585
R2969 GND.n6696 GND.n6695 585
R2970 GND.n6695 GND.n6694 585
R2971 GND.n1410 GND.n1409 585
R2972 GND.n1421 GND.n1410 585
R2973 GND.n6642 GND.n1437 585
R2974 GND.n1437 GND.n1419 585
R2975 GND.n6644 GND.n6643 585
R2976 GND.n6645 GND.n6644 585
R2977 GND.n1438 GND.n1436 585
R2978 GND.n1461 GND.n1436 585
R2979 GND.n6637 GND.n6636 585
R2980 GND.n6636 GND.n6635 585
R2981 GND.n1441 GND.n1440 585
R2982 GND.n1467 GND.n1441 585
R2983 GND.n6604 GND.n6603 585
R2984 GND.n6605 GND.n6604 585
R2985 GND.n1478 GND.n1477 585
R2986 GND.n6573 GND.n1477 585
R2987 GND.n6599 GND.n6598 585
R2988 GND.n6598 GND.t84 585
R2989 GND.n1481 GND.n1480 585
R2990 GND.n6581 GND.n1481 585
R2991 GND.n6552 GND.n6551 585
R2992 GND.n6553 GND.n6552 585
R2993 GND.n1504 GND.n1503 585
R2994 GND.n1525 GND.n1503 585
R2995 GND.n6547 GND.n6546 585
R2996 GND.n6546 GND.n6545 585
R2997 GND.n1507 GND.n1506 585
R2998 GND.n1519 GND.n1507 585
R2999 GND.n6491 GND.n6490 585
R3000 GND.n6490 GND.n1517 585
R3001 GND.n6492 GND.n1539 585
R3002 GND.n1539 GND.n1530 585
R3003 GND.n6494 GND.n6493 585
R3004 GND.n6495 GND.n6494 585
R3005 GND.n1540 GND.n1538 585
R3006 GND.n1547 GND.n1538 585
R3007 GND.n6484 GND.n6483 585
R3008 GND.n6483 GND.n6482 585
R3009 GND.n1543 GND.n1542 585
R3010 GND.n6467 GND.n1543 585
R3011 GND.n6456 GND.n6455 585
R3012 GND.n6457 GND.n6456 585
R3013 GND.n1567 GND.n1566 585
R3014 GND.n6407 GND.n1566 585
R3015 GND.n6451 GND.n6450 585
R3016 GND.n6450 GND.n6449 585
R3017 GND.n1570 GND.n1569 585
R3018 GND.n1578 GND.n1570 585
R3019 GND.n6314 GND.n6313 585
R3020 GND.n6314 GND.n1588 585
R3021 GND.n6315 GND.n6311 585
R3022 GND.n6318 GND.n6317 585
R3023 GND.n6309 GND.n6308 585
R3024 GND.n6308 GND.n1592 585
R3025 GND.n6323 GND.n6322 585
R3026 GND.n6325 GND.n6307 585
R3027 GND.n6328 GND.n6327 585
R3028 GND.n6305 GND.n6304 585
R3029 GND.n6334 GND.n6333 585
R3030 GND.n6336 GND.n6302 585
R3031 GND.n6339 GND.n6338 585
R3032 GND.n6340 GND.n6301 585
R3033 GND.n6342 GND.n6341 585
R3034 GND.n6345 GND.n6344 585
R3035 GND.n6347 GND.n6346 585
R3036 GND.n6350 GND.n6349 585
R3037 GND.n6352 GND.n6351 585
R3038 GND.n6355 GND.n6354 585
R3039 GND.n6357 GND.n6356 585
R3040 GND.n6360 GND.n6359 585
R3041 GND.n6362 GND.n6361 585
R3042 GND.n6364 GND.n6300 585
R3043 GND.n6367 GND.n6366 585
R3044 GND.n1615 GND.n1614 585
R3045 GND.n6373 GND.n6372 585
R3046 GND.n6375 GND.n1613 585
R3047 GND.n6932 GND.n6931 585
R3048 GND.n6934 GND.n1284 585
R3049 GND.n6936 GND.n6935 585
R3050 GND.n6938 GND.n1283 585
R3051 GND.n6943 GND.n6942 585
R3052 GND.n6945 GND.n1282 585
R3053 GND.n6947 GND.n6946 585
R3054 GND.n6948 GND.n1279 585
R3055 GND.n6951 GND.n6950 585
R3056 GND.n6953 GND.n1278 585
R3057 GND.n6955 GND.n6954 585
R3058 GND.n6956 GND.n1198 585
R3059 GND.n6958 GND.n6957 585
R3060 GND.n6960 GND.n1196 585
R3061 GND.n6962 GND.n6961 585
R3062 GND.n6963 GND.n1191 585
R3063 GND.n6965 GND.n6964 585
R3064 GND.n6967 GND.n1189 585
R3065 GND.n6969 GND.n6968 585
R3066 GND.n6970 GND.n1183 585
R3067 GND.n6972 GND.n6971 585
R3068 GND.n6974 GND.n1182 585
R3069 GND.n6975 GND.n1181 585
R3070 GND.n6978 GND.n6977 585
R3071 GND.n6979 GND.n1177 585
R3072 GND.n1177 GND.n1161 585
R3073 GND.n6928 GND.n1174 585
R3074 GND.n6984 GND.n1174 585
R3075 GND.n6927 GND.n6926 585
R3076 GND.n6926 GND.n6925 585
R3077 GND.n1289 GND.n1288 585
R3078 GND.n1295 GND.n1289 585
R3079 GND.n6809 GND.n6808 585
R3080 GND.n6808 GND.n6807 585
R3081 GND.n6810 GND.n1321 585
R3082 GND.n6872 GND.n1321 585
R3083 GND.n6812 GND.n6811 585
R3084 GND.n6812 GND.n1310 585
R3085 GND.n6813 GND.n6800 585
R3086 GND.n6813 GND.n1315 585
R3087 GND.n6815 GND.n6814 585
R3088 GND.n6814 GND.n1314 585
R3089 GND.n6816 GND.n1330 585
R3090 GND.n6857 GND.n1330 585
R3091 GND.n6817 GND.n1339 585
R3092 GND.n6849 GND.n1339 585
R3093 GND.n6818 GND.n1343 585
R3094 GND.n6840 GND.n1343 585
R3095 GND.n6820 GND.n6819 585
R3096 GND.n6821 GND.n6820 585
R3097 GND.n1356 GND.n1350 585
R3098 GND.n6829 GND.n1350 585
R3099 GND.n6792 GND.n6791 585
R3100 GND.n6791 GND.n6790 585
R3101 GND.n1359 GND.n1358 585
R3102 GND.n1364 GND.n1359 585
R3103 GND.n6662 GND.n1372 585
R3104 GND.n6772 GND.n1372 585
R3105 GND.n6664 GND.n6663 585
R3106 GND.t5 GND.n6664 585
R3107 GND.n1426 GND.n1381 585
R3108 GND.n6762 GND.n1381 585
R3109 GND.n6657 GND.n1389 585
R3110 GND.n6754 GND.n1389 585
R3111 GND.n6656 GND.n6655 585
R3112 GND.n6655 GND.n1397 585
R3113 GND.n6654 GND.n1404 585
R3114 GND.n6704 GND.n1404 585
R3115 GND.n1429 GND.n1428 585
R3116 GND.n1428 GND.n1401 585
R3117 GND.n6650 GND.n1412 585
R3118 GND.n6694 GND.n1412 585
R3119 GND.n6649 GND.n6648 585
R3120 GND.n6648 GND.n1421 585
R3121 GND.n6647 GND.n1431 585
R3122 GND.n6647 GND.n1419 585
R3123 GND.n6646 GND.n1433 585
R3124 GND.n6646 GND.n6645 585
R3125 GND.n6566 GND.n1432 585
R3126 GND.n1461 GND.n1432 585
R3127 GND.n6567 GND.n1442 585
R3128 GND.n6635 GND.n1442 585
R3129 GND.n6569 GND.n6568 585
R3130 GND.n6568 GND.n1467 585
R3131 GND.n6570 GND.n1475 585
R3132 GND.n6605 GND.n1475 585
R3133 GND.n6572 GND.n6571 585
R3134 GND.n6573 GND.n6572 585
R3135 GND.n1498 GND.n1483 585
R3136 GND.t84 GND.n1483 585
R3137 GND.n6556 GND.n1492 585
R3138 GND.n6581 GND.n1492 585
R3139 GND.n6555 GND.n6554 585
R3140 GND.n6554 GND.n6553 585
R3141 GND.n1501 GND.n1500 585
R3142 GND.n1525 GND.n1501 585
R3143 GND.n6393 GND.n1509 585
R3144 GND.n6545 GND.n1509 585
R3145 GND.n6395 GND.n6394 585
R3146 GND.n6395 GND.n1519 585
R3147 GND.n6396 GND.n6388 585
R3148 GND.n6396 GND.n1517 585
R3149 GND.n6398 GND.n6397 585
R3150 GND.n6397 GND.n1530 585
R3151 GND.n6399 GND.n1536 585
R3152 GND.n6495 GND.n1536 585
R3153 GND.n6401 GND.n6400 585
R3154 GND.n6400 GND.n1547 585
R3155 GND.n6402 GND.n1545 585
R3156 GND.n6482 GND.n1545 585
R3157 GND.n6403 GND.n1556 585
R3158 GND.n6467 GND.n1556 585
R3159 GND.n6404 GND.n1565 585
R3160 GND.n6457 GND.n1565 585
R3161 GND.n6406 GND.n6405 585
R3162 GND.n6407 GND.n6406 585
R3163 GND.n1610 GND.n1572 585
R3164 GND.n6449 GND.n1572 585
R3165 GND.n6378 GND.n6377 585
R3166 GND.n6377 GND.n1578 585
R3167 GND.n6376 GND.n1612 585
R3168 GND.n6376 GND.n1588 585
R3169 GND.n7510 GND.n862 585
R3170 GND.n7506 GND.n862 585
R3171 GND.n7509 GND.n7508 585
R3172 GND.n7508 GND.n7507 585
R3173 GND.n865 GND.n864 585
R3174 GND.n7483 GND.n865 585
R3175 GND.n7427 GND.n881 585
R3176 GND.n881 GND.n875 585
R3177 GND.n7429 GND.n7428 585
R3178 GND.n7430 GND.n7429 585
R3179 GND.n7426 GND.n880 585
R3180 GND.n886 GND.n880 585
R3181 GND.n7425 GND.n7424 585
R3182 GND.n7424 GND.n7423 585
R3183 GND.n883 GND.n882 585
R3184 GND.n884 GND.n883 585
R3185 GND.n7412 GND.n7411 585
R3186 GND.n7413 GND.n7412 585
R3187 GND.n7410 GND.n895 585
R3188 GND.n895 GND.n892 585
R3189 GND.n7409 GND.n7408 585
R3190 GND.n7408 GND.n7407 585
R3191 GND.n897 GND.n896 585
R3192 GND.n898 GND.n897 585
R3193 GND.n7395 GND.n7394 585
R3194 GND.n7396 GND.n7395 585
R3195 GND.n7393 GND.n904 585
R3196 GND.n7389 GND.n904 585
R3197 GND.n7392 GND.n7391 585
R3198 GND.n7391 GND.n7390 585
R3199 GND.n906 GND.n905 585
R3200 GND.n7377 GND.n906 585
R3201 GND.n7367 GND.n921 585
R3202 GND.n921 GND.n915 585
R3203 GND.n7369 GND.n7368 585
R3204 GND.n7370 GND.n7369 585
R3205 GND.n7366 GND.n920 585
R3206 GND.n926 GND.n920 585
R3207 GND.n7365 GND.n7364 585
R3208 GND.n7364 GND.n7363 585
R3209 GND.n923 GND.n922 585
R3210 GND.n924 GND.n923 585
R3211 GND.n7352 GND.n7351 585
R3212 GND.n7353 GND.n7352 585
R3213 GND.n7350 GND.n935 585
R3214 GND.n935 GND.n932 585
R3215 GND.n7349 GND.n7348 585
R3216 GND.n7348 GND.n7347 585
R3217 GND.n937 GND.n936 585
R3218 GND.n944 GND.n937 585
R3219 GND.n7335 GND.n7334 585
R3220 GND.n7336 GND.n7335 585
R3221 GND.n7333 GND.n946 585
R3222 GND.n946 GND.n943 585
R3223 GND.n7332 GND.n7331 585
R3224 GND.n7331 GND.n7330 585
R3225 GND.n948 GND.n947 585
R3226 GND.n959 GND.n948 585
R3227 GND.n7317 GND.n7316 585
R3228 GND.n7318 GND.n7317 585
R3229 GND.n7315 GND.n960 585
R3230 GND.n960 GND.n957 585
R3231 GND.n7314 GND.n7313 585
R3232 GND.n7313 GND.n7312 585
R3233 GND.n962 GND.n961 585
R3234 GND.n963 GND.n962 585
R3235 GND.n7299 GND.n7298 585
R3236 GND.n7300 GND.n7299 585
R3237 GND.n7297 GND.n970 585
R3238 GND.n974 GND.n970 585
R3239 GND.n7296 GND.n7295 585
R3240 GND.n7295 GND.n7294 585
R3241 GND.n972 GND.n971 585
R3242 GND.n973 GND.n972 585
R3243 GND.n7279 GND.n7278 585
R3244 GND.n7280 GND.n7279 585
R3245 GND.n7277 GND.n985 585
R3246 GND.n985 GND.n982 585
R3247 GND.n7276 GND.n7275 585
R3248 GND.n7275 GND.n7274 585
R3249 GND.n987 GND.n986 585
R3250 GND.n994 GND.n987 585
R3251 GND.n7262 GND.n7261 585
R3252 GND.n7263 GND.n7262 585
R3253 GND.n7260 GND.n996 585
R3254 GND.n996 GND.n993 585
R3255 GND.n7259 GND.n7258 585
R3256 GND.n7258 GND.n7257 585
R3257 GND.n998 GND.n997 585
R3258 GND.n1009 GND.n998 585
R3259 GND.n7244 GND.n7243 585
R3260 GND.n7245 GND.n7244 585
R3261 GND.n7242 GND.n1010 585
R3262 GND.n1010 GND.n1007 585
R3263 GND.n7241 GND.n7240 585
R3264 GND.n7240 GND.n7239 585
R3265 GND.n1012 GND.n1011 585
R3266 GND.n1013 GND.n1012 585
R3267 GND.n7226 GND.n7225 585
R3268 GND.n7227 GND.n7226 585
R3269 GND.n7224 GND.n1020 585
R3270 GND.n7220 GND.n1020 585
R3271 GND.n7223 GND.n7222 585
R3272 GND.n7222 GND.n7221 585
R3273 GND.n1022 GND.n1021 585
R3274 GND.n1028 GND.n1022 585
R3275 GND.n7213 GND.n7212 585
R3276 GND.n7214 GND.n7213 585
R3277 GND.n7211 GND.n1030 585
R3278 GND.n1030 GND.n1027 585
R3279 GND.n7210 GND.n7209 585
R3280 GND.n7209 GND.n7208 585
R3281 GND.n1032 GND.n1031 585
R3282 GND.n1043 GND.n1032 585
R3283 GND.n7186 GND.n7185 585
R3284 GND.n7187 GND.n7186 585
R3285 GND.n7184 GND.n1044 585
R3286 GND.n1044 GND.n1041 585
R3287 GND.n7183 GND.n7182 585
R3288 GND.n7182 GND.n7181 585
R3289 GND.n1046 GND.n1045 585
R3290 GND.n1047 GND.n1046 585
R3291 GND.n7168 GND.n7167 585
R3292 GND.n7169 GND.n7168 585
R3293 GND.n7166 GND.n1053 585
R3294 GND.n1058 GND.n1053 585
R3295 GND.n7165 GND.n7164 585
R3296 GND.n7164 GND.n7163 585
R3297 GND.n1055 GND.n1054 585
R3298 GND.n1056 GND.n1055 585
R3299 GND.n7147 GND.n7146 585
R3300 GND.n7148 GND.n7147 585
R3301 GND.n7145 GND.n1068 585
R3302 GND.n1068 GND.n1065 585
R3303 GND.n7144 GND.n7143 585
R3304 GND.n7143 GND.n7142 585
R3305 GND.n1070 GND.n1069 585
R3306 GND.n1077 GND.n1070 585
R3307 GND.n7130 GND.n7129 585
R3308 GND.n7131 GND.n7130 585
R3309 GND.n7128 GND.n1079 585
R3310 GND.n1079 GND.n1076 585
R3311 GND.n7127 GND.n7126 585
R3312 GND.n7126 GND.n7125 585
R3313 GND.n1081 GND.n1080 585
R3314 GND.n1092 GND.n1081 585
R3315 GND.n7112 GND.n7111 585
R3316 GND.n7113 GND.n7112 585
R3317 GND.n7110 GND.n1093 585
R3318 GND.n1093 GND.n1090 585
R3319 GND.n7109 GND.n7108 585
R3320 GND.n7108 GND.n7107 585
R3321 GND.n1095 GND.n1094 585
R3322 GND.n1096 GND.n1095 585
R3323 GND.n7094 GND.n7093 585
R3324 GND.n7095 GND.n7094 585
R3325 GND.n7092 GND.n1103 585
R3326 GND.n7088 GND.n1103 585
R3327 GND.n7091 GND.n7090 585
R3328 GND.n7090 GND.n7089 585
R3329 GND.n1105 GND.n1104 585
R3330 GND.n1111 GND.n1105 585
R3331 GND.n7081 GND.n7080 585
R3332 GND.n7082 GND.n7081 585
R3333 GND.n7079 GND.n1113 585
R3334 GND.n1113 GND.n1110 585
R3335 GND.n7078 GND.n7077 585
R3336 GND.n7077 GND.n7076 585
R3337 GND.n1115 GND.n1114 585
R3338 GND.n1126 GND.n1115 585
R3339 GND.n7044 GND.n1125 585
R3340 GND.n7056 GND.n1125 585
R3341 GND.n7045 GND.n1134 585
R3342 GND.n1134 GND.n1124 585
R3343 GND.n7047 GND.n7046 585
R3344 GND.n7048 GND.n7047 585
R3345 GND.n7043 GND.n1133 585
R3346 GND.n7039 GND.n1133 585
R3347 GND.n7042 GND.n7041 585
R3348 GND.n7041 GND.n7040 585
R3349 GND.n1136 GND.n1135 585
R3350 GND.n1142 GND.n1136 585
R3351 GND.n7032 GND.n7031 585
R3352 GND.n7033 GND.n7032 585
R3353 GND.n7030 GND.n1144 585
R3354 GND.n1144 GND.n1141 585
R3355 GND.n7029 GND.n7028 585
R3356 GND.n7028 GND.n7027 585
R3357 GND.n1146 GND.n1145 585
R3358 GND.n1157 GND.n1146 585
R3359 GND.n7008 GND.n7007 585
R3360 GND.n7009 GND.n7008 585
R3361 GND.n7006 GND.n1158 585
R3362 GND.n1158 GND.n1155 585
R3363 GND.n7005 GND.n7004 585
R3364 GND.n7004 GND.n7003 585
R3365 GND.n1160 GND.n1159 585
R3366 GND.n1167 GND.n1160 585
R3367 GND.n6990 GND.n6989 585
R3368 GND.n6991 GND.n6990 585
R3369 GND.n6988 GND.n1169 585
R3370 GND.n1175 GND.n1169 585
R3371 GND.n6987 GND.n6986 585
R3372 GND.n6986 GND.n6985 585
R3373 GND.n1171 GND.n1170 585
R3374 GND.n6924 GND.n1171 585
R3375 GND.n6914 GND.n1298 585
R3376 GND.n1298 GND.n1297 585
R3377 GND.n6916 GND.n6915 585
R3378 GND.n6917 GND.n6916 585
R3379 GND.n6913 GND.n1296 585
R3380 GND.n6806 GND.n1296 585
R3381 GND.n6912 GND.n6911 585
R3382 GND.n6911 GND.n6910 585
R3383 GND.n1300 GND.n1299 585
R3384 GND.n6873 GND.n1300 585
R3385 GND.n6885 GND.n6884 585
R3386 GND.n6886 GND.n6885 585
R3387 GND.n6883 GND.n1311 585
R3388 GND.n1311 GND.n1308 585
R3389 GND.n6882 GND.n6881 585
R3390 GND.n6881 GND.n6880 585
R3391 GND.n1313 GND.n1312 585
R3392 GND.n1332 GND.n1313 585
R3393 GND.n6855 GND.n6854 585
R3394 GND.n6856 GND.n6855 585
R3395 GND.n6853 GND.n1334 585
R3396 GND.n6848 GND.n1334 585
R3397 GND.n6852 GND.n6851 585
R3398 GND.n6851 GND.n6850 585
R3399 GND.n1336 GND.n1335 585
R3400 GND.n6841 GND.n1336 585
R3401 GND.n6824 GND.n6823 585
R3402 GND.n6823 GND.n6822 585
R3403 GND.n6825 GND.n1353 585
R3404 GND.n1355 GND.n1353 585
R3405 GND.n6827 GND.n6826 585
R3406 GND.n6828 GND.n6827 585
R3407 GND.n1354 GND.n1352 585
R3408 GND.n6789 GND.n1352 585
R3409 GND.n6777 GND.n1367 585
R3410 GND.n1367 GND.n1360 585
R3411 GND.n6779 GND.n6778 585
R3412 GND.n6780 GND.n6779 585
R3413 GND.n6776 GND.n1366 585
R3414 GND.n1373 GND.n1366 585
R3415 GND.n6775 GND.n6774 585
R3416 GND.n6774 GND.n6773 585
R3417 GND.n1369 GND.n1368 585
R3418 GND.n6665 GND.n1369 585
R3419 GND.n6760 GND.n6759 585
R3420 GND.n6761 GND.n6760 585
R3421 GND.n6758 GND.n1384 585
R3422 GND.n1384 GND.n1380 585
R3423 GND.n6757 GND.n6756 585
R3424 GND.n6756 GND.n6755 585
R3425 GND.n1386 GND.n1385 585
R3426 GND.n6672 GND.n1386 585
R3427 GND.n6712 GND.n6711 585
R3428 GND.n6713 GND.n6712 585
R3429 GND.n6710 GND.n1398 585
R3430 GND.n6705 GND.n1398 585
R3431 GND.n6709 GND.n6708 585
R3432 GND.n6708 GND.n6707 585
R3433 GND.n1400 GND.n1399 585
R3434 GND.n1413 GND.n1400 585
R3435 GND.n1450 GND.n1449 585
R3436 GND.n1450 GND.n1411 585
R3437 GND.n1454 GND.n1453 585
R3438 GND.n1453 GND.n1452 585
R3439 GND.n1455 GND.n1420 585
R3440 GND.n6685 GND.n1420 585
R3441 GND.n1459 GND.n1456 585
R3442 GND.n1459 GND.n1458 585
R3443 GND.n1460 GND.n1448 585
R3444 GND.n1460 GND.n1435 585
R3445 GND.n6630 GND.n6629 585
R3446 GND.n6629 GND.n6628 585
R3447 GND.n6631 GND.n1446 585
R3448 GND.n1462 GND.n1446 585
R3449 GND.n6633 GND.n6632 585
R3450 GND.n6634 GND.n6633 585
R3451 GND.n1447 GND.n1445 585
R3452 GND.n6620 GND.n1445 585
R3453 GND.n6590 GND.n6587 585
R3454 GND.n6590 GND.n6589 585
R3455 GND.n6591 GND.n6586 585
R3456 GND.n6591 GND.n1476 585
R3457 GND.n6593 GND.n6592 585
R3458 GND.n6592 GND.n1474 585
R3459 GND.n6594 GND.n1487 585
R3460 GND.n6574 GND.n1487 585
R3461 GND.n6596 GND.n6595 585
R3462 GND.n6597 GND.n6596 585
R3463 GND.n6585 GND.n1486 585
R3464 GND.n6580 GND.n1486 585
R3465 GND.n6584 GND.n6583 585
R3466 GND.n6583 GND.n6582 585
R3467 GND.n1489 GND.n1488 585
R3468 GND.n1502 GND.n1489 585
R3469 GND.n6520 GND.n1524 585
R3470 GND.n6520 GND.n6519 585
R3471 GND.n6521 GND.n1523 585
R3472 GND.n6521 GND.n1510 585
R3473 GND.n6523 GND.n6522 585
R3474 GND.n6522 GND.n1508 585
R3475 GND.n6524 GND.n1521 585
R3476 GND.n6510 GND.n1521 585
R3477 GND.n6526 GND.n6525 585
R3478 GND.n6527 GND.n6526 585
R3479 GND.n1522 GND.n1520 585
R3480 GND.n6504 GND.n1520 585
R3481 GND.n6501 GND.n6500 585
R3482 GND.n6502 GND.n6501 585
R3483 GND.n6499 GND.n1531 585
R3484 GND.n1596 GND.n1531 585
R3485 GND.n6498 GND.n6497 585
R3486 GND.n6497 GND.n6496 585
R3487 GND.n1533 GND.n1532 585
R3488 GND.n1600 GND.n1533 585
R3489 GND.n6462 GND.n1546 585
R3490 GND.n6481 GND.n1546 585
R3491 GND.n6463 GND.n1560 585
R3492 GND.n1560 GND.n1544 585
R3493 GND.n6465 GND.n6464 585
R3494 GND.n6466 GND.n6465 585
R3495 GND.n6461 GND.n1559 585
R3496 GND.n1559 GND.n1555 585
R3497 GND.n6460 GND.n6459 585
R3498 GND.n6459 GND.n6458 585
R3499 GND.n1562 GND.n1561 585
R3500 GND.n6408 GND.n1562 585
R3501 GND.n6447 GND.n6446 585
R3502 GND.n6448 GND.n6447 585
R3503 GND.n6445 GND.n1575 585
R3504 GND.n1575 GND.n1571 585
R3505 GND.n6444 GND.n6443 585
R3506 GND.n6443 GND.n6442 585
R3507 GND.n1577 GND.n1576 585
R3508 GND.n6416 GND.n1577 585
R3509 GND.n6429 GND.n6428 585
R3510 GND.n6430 GND.n6429 585
R3511 GND.n6427 GND.n1589 585
R3512 GND.n1589 GND.n1586 585
R3513 GND.n6426 GND.n6425 585
R3514 GND.n6425 GND.n6424 585
R3515 GND.n1591 GND.n1590 585
R3516 GND.n5951 GND.n1591 585
R3517 GND.n5930 GND.n5929 585
R3518 GND.n5950 GND.n5930 585
R3519 GND.n5963 GND.n5962 585
R3520 GND.n5962 GND.n5961 585
R3521 GND.n5964 GND.n5927 585
R3522 GND.n5931 GND.n5927 585
R3523 GND.n5966 GND.n5965 585
R3524 GND.n5967 GND.n5966 585
R3525 GND.n5928 GND.n5926 585
R3526 GND.n5926 GND.n5923 585
R3527 GND.n5939 GND.n5938 585
R3528 GND.n5940 GND.n5939 585
R3529 GND.n5909 GND.n5908 585
R3530 GND.n5912 GND.n5909 585
R3531 GND.n5977 GND.n5976 585
R3532 GND.n5976 GND.n5975 585
R3533 GND.n5978 GND.n5903 585
R3534 GND.n5910 GND.n5903 585
R3535 GND.n5980 GND.n5979 585
R3536 GND.n5981 GND.n5980 585
R3537 GND.n5907 GND.n5902 585
R3538 GND.n5902 GND.n5848 585
R3539 GND.n5906 GND.n5847 585
R3540 GND.n5987 GND.n5847 585
R3541 GND.n5905 GND.n5904 585
R3542 GND.n5904 GND.n5846 585
R3543 GND.n5834 GND.n5833 585
R3544 GND.n5837 GND.n5834 585
R3545 GND.n5996 GND.n5995 585
R3546 GND.n5995 GND.n5994 585
R3547 GND.n5997 GND.n5831 585
R3548 GND.n5835 GND.n5831 585
R3549 GND.n5999 GND.n5998 585
R3550 GND.n6000 GND.n5999 585
R3551 GND.n5832 GND.n5830 585
R3552 GND.n5830 GND.n5827 585
R3553 GND.n5886 GND.n5885 585
R3554 GND.n5887 GND.n5886 585
R3555 GND.n5816 GND.n5815 585
R3556 GND.n5819 GND.n5816 585
R3557 GND.n6010 GND.n6009 585
R3558 GND.n6009 GND.n6008 585
R3559 GND.n6011 GND.n5813 585
R3560 GND.n5817 GND.n5813 585
R3561 GND.n6013 GND.n6012 585
R3562 GND.n6014 GND.n6013 585
R3563 GND.n5814 GND.n5812 585
R3564 GND.n5812 GND.n5809 585
R3565 GND.n5873 GND.n5872 585
R3566 GND.n5874 GND.n5873 585
R3567 GND.n5799 GND.n5798 585
R3568 GND.n5870 GND.n5799 585
R3569 GND.n6024 GND.n6023 585
R3570 GND.n6023 GND.n6022 585
R3571 GND.n6025 GND.n5796 585
R3572 GND.n5800 GND.n5796 585
R3573 GND.n6027 GND.n6026 585
R3574 GND.n6028 GND.n6027 585
R3575 GND.n5797 GND.n5795 585
R3576 GND.n5795 GND.n5792 585
R3577 GND.n5859 GND.n5858 585
R3578 GND.n5860 GND.n5859 585
R3579 GND.n5778 GND.n5777 585
R3580 GND.n5781 GND.n5778 585
R3581 GND.n6038 GND.n6037 585
R3582 GND.n6037 GND.n6036 585
R3583 GND.n6039 GND.n5772 585
R3584 GND.n5779 GND.n5772 585
R3585 GND.n6041 GND.n6040 585
R3586 GND.n6042 GND.n6041 585
R3587 GND.n5776 GND.n5771 585
R3588 GND.n5771 GND.n5718 585
R3589 GND.n5775 GND.n5717 585
R3590 GND.n6048 GND.n5717 585
R3591 GND.n5774 GND.n5773 585
R3592 GND.n5773 GND.n5716 585
R3593 GND.n5704 GND.n5703 585
R3594 GND.n5707 GND.n5704 585
R3595 GND.n6057 GND.n6056 585
R3596 GND.n6056 GND.n6055 585
R3597 GND.n6058 GND.n5701 585
R3598 GND.n5705 GND.n5701 585
R3599 GND.n6060 GND.n6059 585
R3600 GND.n6061 GND.n6060 585
R3601 GND.n5702 GND.n5700 585
R3602 GND.n5700 GND.n5697 585
R3603 GND.n5755 GND.n5754 585
R3604 GND.n5756 GND.n5755 585
R3605 GND.n5686 GND.n5685 585
R3606 GND.n5689 GND.n5686 585
R3607 GND.n6071 GND.n6070 585
R3608 GND.n6070 GND.n6069 585
R3609 GND.n6072 GND.n5683 585
R3610 GND.n5687 GND.n5683 585
R3611 GND.n6074 GND.n6073 585
R3612 GND.n6075 GND.n6074 585
R3613 GND.n5684 GND.n5682 585
R3614 GND.n5682 GND.n5679 585
R3615 GND.n5742 GND.n5741 585
R3616 GND.n5743 GND.n5742 585
R3617 GND.n5668 GND.n5667 585
R3618 GND.n5671 GND.n5668 585
R3619 GND.n6085 GND.n6084 585
R3620 GND.n6084 GND.n6083 585
R3621 GND.n6086 GND.n5665 585
R3622 GND.n5669 GND.n5665 585
R3623 GND.n6088 GND.n6087 585
R3624 GND.n6089 GND.n6088 585
R3625 GND.n5666 GND.n5664 585
R3626 GND.n5664 GND.n5661 585
R3627 GND.n5729 GND.n5728 585
R3628 GND.n5730 GND.n5729 585
R3629 GND.n5647 GND.n5646 585
R3630 GND.n5650 GND.n5647 585
R3631 GND.n6099 GND.n6098 585
R3632 GND.n6098 GND.n6097 585
R3633 GND.n6100 GND.n5639 585
R3634 GND.n5648 GND.n5639 585
R3635 GND.n6102 GND.n6101 585
R3636 GND.n6103 GND.n6102 585
R3637 GND.n5645 GND.n5638 585
R3638 GND.n5638 GND.n5585 585
R3639 GND.n5644 GND.n5584 585
R3640 GND.n6109 GND.n5584 585
R3641 GND.n5643 GND.n5642 585
R3642 GND.n5642 GND.n5641 585
R3643 GND.n5573 GND.n5572 585
R3644 GND.n5576 GND.n5573 585
R3645 GND.n6118 GND.n6117 585
R3646 GND.n6117 GND.n6116 585
R3647 GND.n6119 GND.n5570 585
R3648 GND.n5574 GND.n5570 585
R3649 GND.n6121 GND.n6120 585
R3650 GND.n6122 GND.n6121 585
R3651 GND.n5571 GND.n5569 585
R3652 GND.n5569 GND.n5566 585
R3653 GND.n5622 GND.n5621 585
R3654 GND.n5623 GND.n5622 585
R3655 GND.n5555 GND.n5554 585
R3656 GND.n5558 GND.n5555 585
R3657 GND.n6132 GND.n6131 585
R3658 GND.n6131 GND.n6130 585
R3659 GND.n6133 GND.n5552 585
R3660 GND.n5556 GND.n5552 585
R3661 GND.n6135 GND.n6134 585
R3662 GND.n6136 GND.n6135 585
R3663 GND.n5553 GND.n5551 585
R3664 GND.n5551 GND.n5548 585
R3665 GND.n5609 GND.n5608 585
R3666 GND.n5610 GND.n5609 585
R3667 GND.n5537 GND.n5536 585
R3668 GND.n5540 GND.n5537 585
R3669 GND.n6146 GND.n6145 585
R3670 GND.n6145 GND.n6144 585
R3671 GND.n6147 GND.n5534 585
R3672 GND.n5538 GND.n5534 585
R3673 GND.n6149 GND.n6148 585
R3674 GND.n6150 GND.n6149 585
R3675 GND.n5535 GND.n5533 585
R3676 GND.n5533 GND.n5530 585
R3677 GND.n5596 GND.n5595 585
R3678 GND.n5597 GND.n5596 585
R3679 GND.n5515 GND.n5514 585
R3680 GND.n5518 GND.n5515 585
R3681 GND.n6160 GND.n6159 585
R3682 GND.n6159 GND.n6158 585
R3683 GND.n6161 GND.n5509 585
R3684 GND.n5516 GND.n5509 585
R3685 GND.n6163 GND.n6162 585
R3686 GND.n6164 GND.n6163 585
R3687 GND.n5513 GND.n5508 585
R3688 GND.n5508 GND.n5437 585
R3689 GND.n5512 GND.n5436 585
R3690 GND.n6170 GND.n5436 585
R3691 GND.n5511 GND.n5510 585
R3692 GND.n5510 GND.n5435 585
R3693 GND.n5423 GND.n5422 585
R3694 GND.n5426 GND.n5423 585
R3695 GND.n6179 GND.n6178 585
R3696 GND.n6178 GND.n6177 585
R3697 GND.n6180 GND.n5420 585
R3698 GND.n5424 GND.n5420 585
R3699 GND.n6182 GND.n6181 585
R3700 GND.n6183 GND.n6182 585
R3701 GND.n5421 GND.n5419 585
R3702 GND.n5419 GND.n5416 585
R3703 GND.n5493 GND.n5492 585
R3704 GND.n5494 GND.n5493 585
R3705 GND.n1851 GND.n1850 585
R3706 GND.n1854 GND.n1851 585
R3707 GND.n6193 GND.n6192 585
R3708 GND.n6192 GND.n6191 585
R3709 GND.n6194 GND.n1849 585
R3710 GND.n1852 GND.n1849 585
R3711 GND.n6235 GND.n6234 585
R3712 GND.n6233 GND.n1848 585
R3713 GND.n6232 GND.n1847 585
R3714 GND.n6237 GND.n1847 585
R3715 GND.n6231 GND.n6230 585
R3716 GND.n6229 GND.n6228 585
R3717 GND.n6227 GND.n6226 585
R3718 GND.n6225 GND.n6224 585
R3719 GND.n6223 GND.n6222 585
R3720 GND.n6221 GND.n6220 585
R3721 GND.n6219 GND.n6218 585
R3722 GND.n6217 GND.n6216 585
R3723 GND.n6215 GND.n6214 585
R3724 GND.n6213 GND.n6212 585
R3725 GND.n6211 GND.n6210 585
R3726 GND.n6209 GND.n6208 585
R3727 GND.n6207 GND.n6206 585
R3728 GND.n6205 GND.n6204 585
R3729 GND.n6203 GND.n6202 585
R3730 GND.n6200 GND.n6199 585
R3731 GND.n6198 GND.n6197 585
R3732 GND.n1823 GND.n1822 585
R3733 GND.n6240 GND.n6239 585
R3734 GND.n5443 GND.n1820 585
R3735 GND.n5445 GND.n5444 585
R3736 GND.n5447 GND.n5446 585
R3737 GND.n5449 GND.n5448 585
R3738 GND.n5452 GND.n5451 585
R3739 GND.n5454 GND.n5453 585
R3740 GND.n5456 GND.n5455 585
R3741 GND.n5458 GND.n5457 585
R3742 GND.n5460 GND.n5459 585
R3743 GND.n5462 GND.n5461 585
R3744 GND.n5464 GND.n5463 585
R3745 GND.n5466 GND.n5465 585
R3746 GND.n5468 GND.n5467 585
R3747 GND.n5470 GND.n5469 585
R3748 GND.n5472 GND.n5471 585
R3749 GND.n5474 GND.n5473 585
R3750 GND.n5476 GND.n5475 585
R3751 GND.n5478 GND.n5477 585
R3752 GND.n5480 GND.n5479 585
R3753 GND.n5482 GND.n5481 585
R3754 GND.n5484 GND.n5483 585
R3755 GND.n5485 GND.n1845 585
R3756 GND.n6237 GND.n1845 585
R3757 GND.n7478 GND.n7477 585
R3758 GND.n7476 GND.n7475 585
R3759 GND.n7474 GND.n7473 585
R3760 GND.n7472 GND.n7471 585
R3761 GND.n7470 GND.n7469 585
R3762 GND.n7468 GND.n7467 585
R3763 GND.n7466 GND.n7465 585
R3764 GND.n7464 GND.n7463 585
R3765 GND.n7462 GND.n7461 585
R3766 GND.n7460 GND.n7459 585
R3767 GND.n7458 GND.n7457 585
R3768 GND.n7456 GND.n7455 585
R3769 GND.n7454 GND.n7453 585
R3770 GND.n7452 GND.n7451 585
R3771 GND.n7450 GND.n7449 585
R3772 GND.n7448 GND.n7447 585
R3773 GND.n7446 GND.n7445 585
R3774 GND.n7444 GND.n7443 585
R3775 GND.n7442 GND.n7441 585
R3776 GND.n7440 GND.n7439 585
R3777 GND.n7438 GND.n7437 585
R3778 GND.n838 GND.n836 585
R3779 GND.n7557 GND.n7556 585
R3780 GND.n7513 GND.n835 585
R3781 GND.n7515 GND.n7514 585
R3782 GND.n7517 GND.n7516 585
R3783 GND.n7519 GND.n7518 585
R3784 GND.n7522 GND.n7521 585
R3785 GND.n7524 GND.n7523 585
R3786 GND.n7526 GND.n7525 585
R3787 GND.n7528 GND.n7527 585
R3788 GND.n7530 GND.n7529 585
R3789 GND.n7532 GND.n7531 585
R3790 GND.n7534 GND.n7533 585
R3791 GND.n7536 GND.n7535 585
R3792 GND.n7538 GND.n7537 585
R3793 GND.n7540 GND.n7539 585
R3794 GND.n7542 GND.n7541 585
R3795 GND.n7544 GND.n7543 585
R3796 GND.n7546 GND.n7545 585
R3797 GND.n7548 GND.n7547 585
R3798 GND.n7550 GND.n7549 585
R3799 GND.n7552 GND.n7551 585
R3800 GND.n7553 GND.n863 585
R3801 GND.n7555 GND.n7554 585
R3802 GND.n7556 GND.n7555 585
R3803 GND.n7479 GND.n868 585
R3804 GND.n7506 GND.n868 585
R3805 GND.n7480 GND.n867 585
R3806 GND.n7507 GND.n867 585
R3807 GND.n7482 GND.n7481 585
R3808 GND.n7483 GND.n7482 585
R3809 GND.n7433 GND.n876 585
R3810 GND.n876 GND.n875 585
R3811 GND.n7432 GND.n7431 585
R3812 GND.n7431 GND.n7430 585
R3813 GND.n878 GND.n877 585
R3814 GND.n886 GND.n878 585
R3815 GND.n7400 GND.n885 585
R3816 GND.n7423 GND.n885 585
R3817 GND.n7402 GND.n7401 585
R3818 GND.n7401 GND.n884 585
R3819 GND.n7403 GND.n893 585
R3820 GND.n7413 GND.n893 585
R3821 GND.n7404 GND.n900 585
R3822 GND.n900 GND.n892 585
R3823 GND.n7406 GND.n7405 585
R3824 GND.n7407 GND.n7406 585
R3825 GND.n7399 GND.n899 585
R3826 GND.n899 GND.n898 585
R3827 GND.n7398 GND.n7397 585
R3828 GND.n7397 GND.n7396 585
R3829 GND.n902 GND.n901 585
R3830 GND.n7389 GND.n902 585
R3831 GND.n7374 GND.n908 585
R3832 GND.n7390 GND.n908 585
R3833 GND.n7376 GND.n7375 585
R3834 GND.n7377 GND.n7376 585
R3835 GND.n7373 GND.n916 585
R3836 GND.n916 GND.n915 585
R3837 GND.n7372 GND.n7371 585
R3838 GND.n7371 GND.n7370 585
R3839 GND.n918 GND.n917 585
R3840 GND.n926 GND.n918 585
R3841 GND.n7340 GND.n925 585
R3842 GND.n7363 GND.n925 585
R3843 GND.n7342 GND.n7341 585
R3844 GND.n7341 GND.n924 585
R3845 GND.n7343 GND.n933 585
R3846 GND.n7353 GND.n933 585
R3847 GND.n7344 GND.n940 585
R3848 GND.n940 GND.n932 585
R3849 GND.n7346 GND.n7345 585
R3850 GND.n7347 GND.n7346 585
R3851 GND.n7339 GND.n939 585
R3852 GND.n944 GND.n939 585
R3853 GND.n7338 GND.n7337 585
R3854 GND.n7337 GND.n7336 585
R3855 GND.n942 GND.n941 585
R3856 GND.n943 GND.n942 585
R3857 GND.n7304 GND.n950 585
R3858 GND.n7330 GND.n950 585
R3859 GND.n7306 GND.n7305 585
R3860 GND.n7305 GND.n959 585
R3861 GND.n7307 GND.n958 585
R3862 GND.n7318 GND.n958 585
R3863 GND.n7308 GND.n965 585
R3864 GND.n965 GND.n957 585
R3865 GND.n7310 GND.n7309 585
R3866 GND.n7312 GND.n7310 585
R3867 GND.n7303 GND.n964 585
R3868 GND.n964 GND.n963 585
R3869 GND.n7302 GND.n7301 585
R3870 GND.n7301 GND.n7300 585
R3871 GND.n967 GND.n966 585
R3872 GND.n974 GND.n967 585
R3873 GND.n7267 GND.n975 585
R3874 GND.n7294 GND.n975 585
R3875 GND.n7269 GND.n7268 585
R3876 GND.n7268 GND.n973 585
R3877 GND.n7270 GND.n983 585
R3878 GND.n7280 GND.n983 585
R3879 GND.n7271 GND.n990 585
R3880 GND.n990 GND.n982 585
R3881 GND.n7273 GND.n7272 585
R3882 GND.n7274 GND.n7273 585
R3883 GND.n7266 GND.n989 585
R3884 GND.n994 GND.n989 585
R3885 GND.n7265 GND.n7264 585
R3886 GND.n7264 GND.n7263 585
R3887 GND.n992 GND.n991 585
R3888 GND.n993 GND.n992 585
R3889 GND.n7231 GND.n1000 585
R3890 GND.n7257 GND.n1000 585
R3891 GND.n7233 GND.n7232 585
R3892 GND.n7232 GND.n1009 585
R3893 GND.n7234 GND.n1008 585
R3894 GND.n7245 GND.n1008 585
R3895 GND.n7235 GND.n1015 585
R3896 GND.n1015 GND.n1007 585
R3897 GND.n7237 GND.n7236 585
R3898 GND.n7239 GND.n7237 585
R3899 GND.n7230 GND.n1014 585
R3900 GND.n1014 GND.n1013 585
R3901 GND.n7229 GND.n7228 585
R3902 GND.n7228 GND.n7227 585
R3903 GND.n1017 GND.n1016 585
R3904 GND.n7220 GND.n1017 585
R3905 GND.n7219 GND.n7218 585
R3906 GND.n7221 GND.n7219 585
R3907 GND.n7217 GND.n1024 585
R3908 GND.n1028 GND.n1024 585
R3909 GND.n7216 GND.n7215 585
R3910 GND.n7215 GND.n7214 585
R3911 GND.n1026 GND.n1025 585
R3912 GND.n1027 GND.n1026 585
R3913 GND.n7173 GND.n1034 585
R3914 GND.n7208 GND.n1034 585
R3915 GND.n7175 GND.n7174 585
R3916 GND.n7174 GND.n1043 585
R3917 GND.n7176 GND.n1042 585
R3918 GND.n7187 GND.n1042 585
R3919 GND.n7177 GND.n1049 585
R3920 GND.n1049 GND.n1041 585
R3921 GND.n7179 GND.n7178 585
R3922 GND.n7181 GND.n7179 585
R3923 GND.n7172 GND.n1048 585
R3924 GND.n1048 GND.n1047 585
R3925 GND.n7171 GND.n7170 585
R3926 GND.n7170 GND.n7169 585
R3927 GND.n1051 GND.n1050 585
R3928 GND.n1058 GND.n1051 585
R3929 GND.n7135 GND.n1057 585
R3930 GND.n7163 GND.n1057 585
R3931 GND.n7137 GND.n7136 585
R3932 GND.n7136 GND.n1056 585
R3933 GND.n7138 GND.n1066 585
R3934 GND.n7148 GND.n1066 585
R3935 GND.n7139 GND.n1073 585
R3936 GND.n1073 GND.n1065 585
R3937 GND.n7141 GND.n7140 585
R3938 GND.n7142 GND.n7141 585
R3939 GND.n7134 GND.n1072 585
R3940 GND.n1077 GND.n1072 585
R3941 GND.n7133 GND.n7132 585
R3942 GND.n7132 GND.n7131 585
R3943 GND.n1075 GND.n1074 585
R3944 GND.n1076 GND.n1075 585
R3945 GND.n7099 GND.n1083 585
R3946 GND.n7125 GND.n1083 585
R3947 GND.n7101 GND.n7100 585
R3948 GND.n7100 GND.n1092 585
R3949 GND.n7102 GND.n1091 585
R3950 GND.n7113 GND.n1091 585
R3951 GND.n7103 GND.n1098 585
R3952 GND.n1098 GND.n1090 585
R3953 GND.n7105 GND.n7104 585
R3954 GND.n7107 GND.n7105 585
R3955 GND.n7098 GND.n1097 585
R3956 GND.n1097 GND.n1096 585
R3957 GND.n7097 GND.n7096 585
R3958 GND.n7096 GND.n7095 585
R3959 GND.n1100 GND.n1099 585
R3960 GND.n7088 GND.n1100 585
R3961 GND.n7087 GND.n7086 585
R3962 GND.n7089 GND.n7087 585
R3963 GND.n7085 GND.n1107 585
R3964 GND.n1111 GND.n1107 585
R3965 GND.n7084 GND.n7083 585
R3966 GND.n7083 GND.n7082 585
R3967 GND.n1109 GND.n1108 585
R3968 GND.n1110 GND.n1109 585
R3969 GND.n7052 GND.n1117 585
R3970 GND.n7076 GND.n1117 585
R3971 GND.n7053 GND.n1128 585
R3972 GND.n1128 GND.n1126 585
R3973 GND.n7055 GND.n7054 585
R3974 GND.n7056 GND.n7055 585
R3975 GND.n7051 GND.n1127 585
R3976 GND.n1127 GND.n1124 585
R3977 GND.n7050 GND.n7049 585
R3978 GND.n7049 GND.n7048 585
R3979 GND.n1130 GND.n1129 585
R3980 GND.n7039 GND.n1130 585
R3981 GND.n7038 GND.n7037 585
R3982 GND.n7040 GND.n7038 585
R3983 GND.n7036 GND.n1138 585
R3984 GND.n1142 GND.n1138 585
R3985 GND.n7035 GND.n7034 585
R3986 GND.n7034 GND.n7033 585
R3987 GND.n1140 GND.n1139 585
R3988 GND.n1141 GND.n1140 585
R3989 GND.n6995 GND.n1148 585
R3990 GND.n7027 GND.n1148 585
R3991 GND.n6997 GND.n6996 585
R3992 GND.n6996 GND.n1157 585
R3993 GND.n6998 GND.n1156 585
R3994 GND.n7009 GND.n1156 585
R3995 GND.n6999 GND.n1163 585
R3996 GND.n1163 GND.n1155 585
R3997 GND.n7001 GND.n7000 585
R3998 GND.n7003 GND.n7001 585
R3999 GND.n6994 GND.n1162 585
R4000 GND.n1167 GND.n1162 585
R4001 GND.n6993 GND.n6992 585
R4002 GND.n6992 GND.n6991 585
R4003 GND.n1165 GND.n1164 585
R4004 GND.n1175 GND.n1165 585
R4005 GND.n6921 GND.n1173 585
R4006 GND.n6985 GND.n1173 585
R4007 GND.n6923 GND.n6922 585
R4008 GND.n6924 GND.n6923 585
R4009 GND.n6920 GND.n1291 585
R4010 GND.n1297 GND.n1291 585
R4011 GND.n6919 GND.n6918 585
R4012 GND.n6918 GND.n6917 585
R4013 GND.n1293 GND.n1292 585
R4014 GND.n6806 GND.n1293 585
R4015 GND.n1319 GND.n1301 585
R4016 GND.n6910 GND.n1301 585
R4017 GND.n6875 GND.n6874 585
R4018 GND.n6874 GND.n6873 585
R4019 GND.n6876 GND.n1309 585
R4020 GND.n6886 GND.n1309 585
R4021 GND.n6877 GND.n1317 585
R4022 GND.n1317 GND.n1308 585
R4023 GND.n6879 GND.n6878 585
R4024 GND.n6880 GND.n6879 585
R4025 GND.n1318 GND.n1316 585
R4026 GND.n1332 GND.n1316 585
R4027 GND.n6845 GND.n1331 585
R4028 GND.n6856 GND.n1331 585
R4029 GND.n6847 GND.n6846 585
R4030 GND.n6848 GND.n6847 585
R4031 GND.n6844 GND.n1338 585
R4032 GND.n6850 GND.n1338 585
R4033 GND.n6843 GND.n6842 585
R4034 GND.n6842 GND.n6841 585
R4035 GND.n1341 GND.n1340 585
R4036 GND.n6822 GND.n1341 585
R4037 GND.n6785 GND.n6784 585
R4038 GND.n6784 GND.n1355 585
R4039 GND.n6786 GND.n1351 585
R4040 GND.n6828 GND.n1351 585
R4041 GND.n6788 GND.n6787 585
R4042 GND.n6789 GND.n6788 585
R4043 GND.n6783 GND.n1361 585
R4044 GND.n1361 GND.n1360 585
R4045 GND.n6782 GND.n6781 585
R4046 GND.n6781 GND.n6780 585
R4047 GND.n1363 GND.n1362 585
R4048 GND.n1373 GND.n1363 585
R4049 GND.n1425 GND.n1371 585
R4050 GND.n6773 GND.n1371 585
R4051 GND.n6667 GND.n6666 585
R4052 GND.n6666 GND.n6665 585
R4053 GND.n6668 GND.n1382 585
R4054 GND.n6761 GND.n1382 585
R4055 GND.n6670 GND.n6669 585
R4056 GND.n6669 GND.n1380 585
R4057 GND.n6671 GND.n1388 585
R4058 GND.n6755 GND.n1388 585
R4059 GND.n6674 GND.n6673 585
R4060 GND.n6673 GND.n6672 585
R4061 GND.n6675 GND.n1396 585
R4062 GND.n6713 GND.n1396 585
R4063 GND.n6676 GND.n1403 585
R4064 GND.n6705 GND.n1403 585
R4065 GND.n6677 GND.n1402 585
R4066 GND.n6707 GND.n1402 585
R4067 GND.n6679 GND.n6678 585
R4068 GND.n6679 GND.n1413 585
R4069 GND.n6681 GND.n6680 585
R4070 GND.n6680 GND.n1411 585
R4071 GND.n6682 GND.n1423 585
R4072 GND.n1452 GND.n1423 585
R4073 GND.n6684 GND.n6683 585
R4074 GND.n6685 GND.n6684 585
R4075 GND.n1424 GND.n1422 585
R4076 GND.n1458 GND.n1422 585
R4077 GND.n6625 GND.n1464 585
R4078 GND.n1464 GND.n1435 585
R4079 GND.n6627 GND.n6626 585
R4080 GND.n6628 GND.n6627 585
R4081 GND.n6624 GND.n1463 585
R4082 GND.n1463 GND.n1462 585
R4083 GND.n6623 GND.n1443 585
R4084 GND.n6634 GND.n1443 585
R4085 GND.n6622 GND.n6621 585
R4086 GND.n6621 GND.n6620 585
R4087 GND.n1466 GND.n1465 585
R4088 GND.n6589 GND.n1466 585
R4089 GND.n1496 GND.n1495 585
R4090 GND.n1496 GND.n1476 585
R4091 GND.n1497 GND.n1494 585
R4092 GND.n1497 GND.n1474 585
R4093 GND.n6576 GND.n6575 585
R4094 GND.n6575 GND.n6574 585
R4095 GND.n6577 GND.n1484 585
R4096 GND.n6597 GND.n1484 585
R4097 GND.n6579 GND.n6578 585
R4098 GND.n6580 GND.n6579 585
R4099 GND.n1493 GND.n1491 585
R4100 GND.n6582 GND.n1491 585
R4101 GND.n6515 GND.n1527 585
R4102 GND.n1527 GND.n1502 585
R4103 GND.n6517 GND.n6516 585
R4104 GND.n6519 GND.n6517 585
R4105 GND.n6514 GND.n1526 585
R4106 GND.n1526 GND.n1510 585
R4107 GND.n6513 GND.n6512 585
R4108 GND.n6512 GND.n1508 585
R4109 GND.n6511 GND.n6508 585
R4110 GND.n6511 GND.n6510 585
R4111 GND.n6507 GND.n1518 585
R4112 GND.n6527 GND.n1518 585
R4113 GND.n6506 GND.n6505 585
R4114 GND.n6505 GND.n6504 585
R4115 GND.n1529 GND.n1528 585
R4116 GND.n6502 GND.n1529 585
R4117 GND.n1598 GND.n1597 585
R4118 GND.n1597 GND.n1596 585
R4119 GND.n1599 GND.n1535 585
R4120 GND.n6496 GND.n1535 585
R4121 GND.n1602 GND.n1601 585
R4122 GND.n1601 GND.n1600 585
R4123 GND.n1603 GND.n1548 585
R4124 GND.n6481 GND.n1548 585
R4125 GND.n1605 GND.n1604 585
R4126 GND.n1604 GND.n1544 585
R4127 GND.n1606 GND.n1557 585
R4128 GND.n6466 GND.n1557 585
R4129 GND.n1608 GND.n1607 585
R4130 GND.n1607 GND.n1555 585
R4131 GND.n1609 GND.n1564 585
R4132 GND.n6458 GND.n1564 585
R4133 GND.n6410 GND.n6409 585
R4134 GND.n6409 GND.n6408 585
R4135 GND.n6411 GND.n1573 585
R4136 GND.n6448 GND.n1573 585
R4137 GND.n6413 GND.n6412 585
R4138 GND.n6412 GND.n1571 585
R4139 GND.n6414 GND.n1579 585
R4140 GND.n6442 GND.n1579 585
R4141 GND.n6418 GND.n6417 585
R4142 GND.n6417 GND.n6416 585
R4143 GND.n6419 GND.n1587 585
R4144 GND.n6430 GND.n1587 585
R4145 GND.n6420 GND.n1594 585
R4146 GND.n1594 GND.n1586 585
R4147 GND.n6422 GND.n6421 585
R4148 GND.n6424 GND.n6422 585
R4149 GND.n1595 GND.n1593 585
R4150 GND.n5951 GND.n1593 585
R4151 GND.n5949 GND.n5948 585
R4152 GND.n5950 GND.n5949 585
R4153 GND.n5947 GND.n5932 585
R4154 GND.n5961 GND.n5932 585
R4155 GND.n5946 GND.n5945 585
R4156 GND.n5945 GND.n5931 585
R4157 GND.n5944 GND.n5924 585
R4158 GND.n5967 GND.n5924 585
R4159 GND.n5943 GND.n5942 585
R4160 GND.n5942 GND.n5923 585
R4161 GND.n5941 GND.n5933 585
R4162 GND.n5941 GND.n5940 585
R4163 GND.n5936 GND.n5935 585
R4164 GND.n5936 GND.n5912 585
R4165 GND.n5934 GND.n5911 585
R4166 GND.n5975 GND.n5911 585
R4167 GND.n5899 GND.n5898 585
R4168 GND.n5910 GND.n5899 585
R4169 GND.n5983 GND.n5982 585
R4170 GND.n5982 GND.n5981 585
R4171 GND.n5984 GND.n5850 585
R4172 GND.n5850 GND.n5848 585
R4173 GND.n5986 GND.n5985 585
R4174 GND.n5987 GND.n5986 585
R4175 GND.n5897 GND.n5849 585
R4176 GND.n5849 GND.n5846 585
R4177 GND.n5896 GND.n5895 585
R4178 GND.n5895 GND.n5837 585
R4179 GND.n5894 GND.n5836 585
R4180 GND.n5994 GND.n5836 585
R4181 GND.n5893 GND.n5892 585
R4182 GND.n5892 GND.n5835 585
R4183 GND.n5891 GND.n5828 585
R4184 GND.n6000 GND.n5828 585
R4185 GND.n5890 GND.n5889 585
R4186 GND.n5889 GND.n5827 585
R4187 GND.n5888 GND.n5851 585
R4188 GND.n5888 GND.n5887 585
R4189 GND.n5883 GND.n5882 585
R4190 GND.n5883 GND.n5819 585
R4191 GND.n5881 GND.n5818 585
R4192 GND.n6008 GND.n5818 585
R4193 GND.n5880 GND.n5879 585
R4194 GND.n5879 GND.n5817 585
R4195 GND.n5878 GND.n5810 585
R4196 GND.n6014 GND.n5810 585
R4197 GND.n5877 GND.n5876 585
R4198 GND.n5876 GND.n5809 585
R4199 GND.n5875 GND.n5852 585
R4200 GND.n5875 GND.n5874 585
R4201 GND.n5869 GND.n5868 585
R4202 GND.n5870 GND.n5869 585
R4203 GND.n5867 GND.n5801 585
R4204 GND.n6022 GND.n5801 585
R4205 GND.n5866 GND.n5865 585
R4206 GND.n5865 GND.n5800 585
R4207 GND.n5864 GND.n5793 585
R4208 GND.n6028 GND.n5793 585
R4209 GND.n5863 GND.n5862 585
R4210 GND.n5862 GND.n5792 585
R4211 GND.n5861 GND.n5853 585
R4212 GND.n5861 GND.n5860 585
R4213 GND.n5856 GND.n5855 585
R4214 GND.n5856 GND.n5781 585
R4215 GND.n5854 GND.n5780 585
R4216 GND.n6036 GND.n5780 585
R4217 GND.n5768 GND.n5767 585
R4218 GND.n5779 GND.n5768 585
R4219 GND.n6044 GND.n6043 585
R4220 GND.n6043 GND.n6042 585
R4221 GND.n6045 GND.n5720 585
R4222 GND.n5720 GND.n5718 585
R4223 GND.n6047 GND.n6046 585
R4224 GND.n6048 GND.n6047 585
R4225 GND.n5766 GND.n5719 585
R4226 GND.n5719 GND.n5716 585
R4227 GND.n5765 GND.n5764 585
R4228 GND.n5764 GND.n5707 585
R4229 GND.n5763 GND.n5706 585
R4230 GND.n6055 GND.n5706 585
R4231 GND.n5762 GND.n5761 585
R4232 GND.n5761 GND.n5705 585
R4233 GND.n5760 GND.n5698 585
R4234 GND.n6061 GND.n5698 585
R4235 GND.n5759 GND.n5758 585
R4236 GND.n5758 GND.n5697 585
R4237 GND.n5757 GND.n5721 585
R4238 GND.n5757 GND.n5756 585
R4239 GND.n5752 GND.n5751 585
R4240 GND.n5752 GND.n5689 585
R4241 GND.n5750 GND.n5688 585
R4242 GND.n6069 GND.n5688 585
R4243 GND.n5749 GND.n5748 585
R4244 GND.n5748 GND.n5687 585
R4245 GND.n5747 GND.n5680 585
R4246 GND.n6075 GND.n5680 585
R4247 GND.n5746 GND.n5745 585
R4248 GND.n5745 GND.n5679 585
R4249 GND.n5744 GND.n5722 585
R4250 GND.n5744 GND.n5743 585
R4251 GND.n5739 GND.n5738 585
R4252 GND.n5739 GND.n5671 585
R4253 GND.n5737 GND.n5670 585
R4254 GND.n6083 GND.n5670 585
R4255 GND.n5736 GND.n5735 585
R4256 GND.n5735 GND.n5669 585
R4257 GND.n5734 GND.n5662 585
R4258 GND.n6089 GND.n5662 585
R4259 GND.n5733 GND.n5732 585
R4260 GND.n5732 GND.n5661 585
R4261 GND.n5731 GND.n5723 585
R4262 GND.n5731 GND.n5730 585
R4263 GND.n5726 GND.n5725 585
R4264 GND.n5726 GND.n5650 585
R4265 GND.n5724 GND.n5649 585
R4266 GND.n6097 GND.n5649 585
R4267 GND.n5635 GND.n5634 585
R4268 GND.n5648 GND.n5635 585
R4269 GND.n6105 GND.n6104 585
R4270 GND.n6104 GND.n6103 585
R4271 GND.n6106 GND.n5587 585
R4272 GND.n5587 GND.n5585 585
R4273 GND.n6108 GND.n6107 585
R4274 GND.n6109 GND.n6108 585
R4275 GND.n5633 GND.n5586 585
R4276 GND.n5641 GND.n5586 585
R4277 GND.n5632 GND.n5631 585
R4278 GND.n5631 GND.n5576 585
R4279 GND.n5630 GND.n5575 585
R4280 GND.n6116 GND.n5575 585
R4281 GND.n5629 GND.n5628 585
R4282 GND.n5628 GND.n5574 585
R4283 GND.n5627 GND.n5567 585
R4284 GND.n6122 GND.n5567 585
R4285 GND.n5626 GND.n5625 585
R4286 GND.n5625 GND.n5566 585
R4287 GND.n5624 GND.n5588 585
R4288 GND.n5624 GND.n5623 585
R4289 GND.n5619 GND.n5618 585
R4290 GND.n5619 GND.n5558 585
R4291 GND.n5617 GND.n5557 585
R4292 GND.n6130 GND.n5557 585
R4293 GND.n5616 GND.n5615 585
R4294 GND.n5615 GND.n5556 585
R4295 GND.n5614 GND.n5549 585
R4296 GND.n6136 GND.n5549 585
R4297 GND.n5613 GND.n5612 585
R4298 GND.n5612 GND.n5548 585
R4299 GND.n5611 GND.n5589 585
R4300 GND.n5611 GND.n5610 585
R4301 GND.n5606 GND.n5605 585
R4302 GND.n5606 GND.n5540 585
R4303 GND.n5604 GND.n5539 585
R4304 GND.n6144 GND.n5539 585
R4305 GND.n5603 GND.n5602 585
R4306 GND.n5602 GND.n5538 585
R4307 GND.n5601 GND.n5531 585
R4308 GND.n6150 GND.n5531 585
R4309 GND.n5600 GND.n5599 585
R4310 GND.n5599 GND.n5530 585
R4311 GND.n5598 GND.n5590 585
R4312 GND.n5598 GND.n5597 585
R4313 GND.n5593 GND.n5592 585
R4314 GND.n5593 GND.n5518 585
R4315 GND.n5591 GND.n5517 585
R4316 GND.n6158 GND.n5517 585
R4317 GND.n5506 GND.n5505 585
R4318 GND.n5516 GND.n5506 585
R4319 GND.n6166 GND.n6165 585
R4320 GND.n6165 GND.n6164 585
R4321 GND.n6167 GND.n5439 585
R4322 GND.n5439 GND.n5437 585
R4323 GND.n6169 GND.n6168 585
R4324 GND.n6170 GND.n6169 585
R4325 GND.n5504 GND.n5438 585
R4326 GND.n5438 GND.n5435 585
R4327 GND.n5503 GND.n5502 585
R4328 GND.n5502 GND.n5426 585
R4329 GND.n5501 GND.n5425 585
R4330 GND.n6177 GND.n5425 585
R4331 GND.n5500 GND.n5499 585
R4332 GND.n5499 GND.n5424 585
R4333 GND.n5498 GND.n5417 585
R4334 GND.n6183 GND.n5417 585
R4335 GND.n5497 GND.n5496 585
R4336 GND.n5496 GND.n5416 585
R4337 GND.n5495 GND.n5440 585
R4338 GND.n5495 GND.n5494 585
R4339 GND.n5490 GND.n5489 585
R4340 GND.n5490 GND.n1854 585
R4341 GND.n5488 GND.n1853 585
R4342 GND.n6191 GND.n1853 585
R4343 GND.n5487 GND.n5486 585
R4344 GND.n5486 GND.n1852 585
R4345 GND.n2134 GND.n1632 585
R4346 GND.n6286 GND.n1632 585
R4347 GND.n2136 GND.n2135 585
R4348 GND.n2135 GND.n1630 585
R4349 GND.n2137 GND.n1870 585
R4350 GND.n5387 GND.n1870 585
R4351 GND.n2139 GND.n2138 585
R4352 GND.n2138 GND.n1869 585
R4353 GND.n2140 GND.n1879 585
R4354 GND.n5378 GND.n1879 585
R4355 GND.n2142 GND.n2141 585
R4356 GND.n2141 GND.n1878 585
R4357 GND.n2143 GND.n1887 585
R4358 GND.n5368 GND.n1887 585
R4359 GND.n2144 GND.n1898 585
R4360 GND.n5357 GND.n1898 585
R4361 GND.n2146 GND.n2145 585
R4362 GND.n2145 GND.n1897 585
R4363 GND.n2147 GND.n1905 585
R4364 GND.n5333 GND.n1905 585
R4365 GND.n2149 GND.n2148 585
R4366 GND.n2148 GND.n1904 585
R4367 GND.n2150 GND.n1915 585
R4368 GND.n5323 GND.n1915 585
R4369 GND.n2152 GND.n2151 585
R4370 GND.n2151 GND.n1914 585
R4371 GND.n2153 GND.n1926 585
R4372 GND.n5306 GND.n1926 585
R4373 GND.n2155 GND.n2154 585
R4374 GND.n2154 GND.n1925 585
R4375 GND.n2156 GND.n1935 585
R4376 GND.n5298 GND.n1935 585
R4377 GND.n2158 GND.n2157 585
R4378 GND.n2157 GND.n1934 585
R4379 GND.n2159 GND.n1946 585
R4380 GND.n5286 GND.n1946 585
R4381 GND.n2161 GND.n2160 585
R4382 GND.n2160 GND.n1945 585
R4383 GND.n2162 GND.n1955 585
R4384 GND.n5278 GND.n1955 585
R4385 GND.n2164 GND.n2163 585
R4386 GND.n2163 GND.n1954 585
R4387 GND.n2165 GND.n1966 585
R4388 GND.n5266 GND.n1966 585
R4389 GND.n2167 GND.n2166 585
R4390 GND.n2166 GND.n1965 585
R4391 GND.n2168 GND.n1975 585
R4392 GND.n5258 GND.n1975 585
R4393 GND.n2170 GND.n2169 585
R4394 GND.n2169 GND.n1974 585
R4395 GND.n2171 GND.n1986 585
R4396 GND.n5246 GND.n1986 585
R4397 GND.n2173 GND.n2172 585
R4398 GND.n2172 GND.n1985 585
R4399 GND.n2174 GND.n1995 585
R4400 GND.n5238 GND.n1995 585
R4401 GND.n2176 GND.n2175 585
R4402 GND.n2175 GND.n1994 585
R4403 GND.n2177 GND.n2006 585
R4404 GND.n5226 GND.n2006 585
R4405 GND.n2179 GND.n2178 585
R4406 GND.n2178 GND.n2005 585
R4407 GND.n2180 GND.n2015 585
R4408 GND.n5218 GND.n2015 585
R4409 GND.n2182 GND.n2181 585
R4410 GND.n2181 GND.n2014 585
R4411 GND.n2183 GND.n2026 585
R4412 GND.n5206 GND.n2026 585
R4413 GND.n2185 GND.n2184 585
R4414 GND.n2184 GND.n2025 585
R4415 GND.n2186 GND.n2034 585
R4416 GND.n5198 GND.n2034 585
R4417 GND.n2187 GND.n2045 585
R4418 GND.n5187 GND.n2045 585
R4419 GND.n2189 GND.n2188 585
R4420 GND.n2188 GND.n2044 585
R4421 GND.n2190 GND.n2052 585
R4422 GND.n5117 GND.n2052 585
R4423 GND.n2192 GND.n2191 585
R4424 GND.n2191 GND.n2051 585
R4425 GND.n2193 GND.n2062 585
R4426 GND.n5107 GND.n2062 585
R4427 GND.n2195 GND.n2194 585
R4428 GND.n2194 GND.n2061 585
R4429 GND.n2196 GND.n2073 585
R4430 GND.n5090 GND.n2073 585
R4431 GND.n5084 GND.n5083 585
R4432 GND.n5083 GND.n2072 585
R4433 GND.n5082 GND.n2092 585
R4434 GND.n5082 GND.n5081 585
R4435 GND.n2206 GND.n2197 585
R4436 GND.n2198 GND.n2197 585
R4437 GND.n2208 GND.n2207 585
R4438 GND.n5075 GND.n2208 585
R4439 GND.n2220 GND.n2219 585
R4440 GND.n2219 GND.n2205 585
R4441 GND.n2222 GND.n2221 585
R4442 GND.t34 GND.n2222 585
R4443 GND.n2229 GND.n2228 585
R4444 GND.n2228 GND.n2218 585
R4445 GND.n2231 GND.n2230 585
R4446 GND.n5050 GND.n2231 585
R4447 GND.n2243 GND.n2242 585
R4448 GND.n2242 GND.n2227 585
R4449 GND.n2245 GND.n2244 585
R4450 GND.n5038 GND.n2245 585
R4451 GND.n2657 GND.n2656 585
R4452 GND.n2657 GND.n2241 585
R4453 GND.n2659 GND.n2658 585
R4454 GND.n2658 GND.n2255 585
R4455 GND.n2660 GND.n2253 585
R4456 GND.n5030 GND.n2253 585
R4457 GND.n2662 GND.n2661 585
R4458 GND.n2661 GND.n2252 585
R4459 GND.n2663 GND.n2265 585
R4460 GND.n5013 GND.n2265 585
R4461 GND.n2665 GND.n2664 585
R4462 GND.n2664 GND.n2264 585
R4463 GND.n2666 GND.n2274 585
R4464 GND.n5004 GND.n2274 585
R4465 GND.n2668 GND.n2667 585
R4466 GND.n2667 GND.n2273 585
R4467 GND.n2669 GND.n2285 585
R4468 GND.n4992 GND.n2285 585
R4469 GND.n2671 GND.n2670 585
R4470 GND.n2670 GND.n2284 585
R4471 GND.n2672 GND.n2294 585
R4472 GND.n4984 GND.n2294 585
R4473 GND.n2674 GND.n2673 585
R4474 GND.n2673 GND.n2293 585
R4475 GND.n2675 GND.n2305 585
R4476 GND.n4972 GND.n2305 585
R4477 GND.n2677 GND.n2676 585
R4478 GND.n2676 GND.n2304 585
R4479 GND.n2678 GND.n2314 585
R4480 GND.n4964 GND.n2314 585
R4481 GND.n2680 GND.n2679 585
R4482 GND.n2679 GND.n2313 585
R4483 GND.n2681 GND.n2325 585
R4484 GND.n4952 GND.n2325 585
R4485 GND.n2683 GND.n2682 585
R4486 GND.n2682 GND.n2324 585
R4487 GND.n2684 GND.n2334 585
R4488 GND.n4944 GND.n2334 585
R4489 GND.n2686 GND.n2685 585
R4490 GND.n2685 GND.n2333 585
R4491 GND.n2687 GND.n2344 585
R4492 GND.n4932 GND.n2344 585
R4493 GND.n2689 GND.n2688 585
R4494 GND.n2688 GND.n2355 585
R4495 GND.n2690 GND.n2353 585
R4496 GND.n4924 GND.n2353 585
R4497 GND.n2692 GND.n2691 585
R4498 GND.n2691 GND.n2352 585
R4499 GND.n2693 GND.n2365 585
R4500 GND.n4912 GND.n2365 585
R4501 GND.n2695 GND.n2694 585
R4502 GND.n2694 GND.n2364 585
R4503 GND.n2696 GND.n2374 585
R4504 GND.n4904 GND.n2374 585
R4505 GND.n2698 GND.n2697 585
R4506 GND.n2697 GND.n2373 585
R4507 GND.n2699 GND.n2385 585
R4508 GND.n4892 GND.n2385 585
R4509 GND.n2701 GND.n2700 585
R4510 GND.n2700 GND.n2384 585
R4511 GND.n2702 GND.n2394 585
R4512 GND.n4884 GND.n2394 585
R4513 GND.n2704 GND.n2703 585
R4514 GND.n2703 GND.n2393 585
R4515 GND.n2705 GND.n2405 585
R4516 GND.n4872 GND.n2405 585
R4517 GND.n2707 GND.n2706 585
R4518 GND.n2706 GND.n2404 585
R4519 GND.n2708 GND.n2414 585
R4520 GND.n4864 GND.n2414 585
R4521 GND.n2710 GND.n2709 585
R4522 GND.n2709 GND.n2413 585
R4523 GND.n2711 GND.n2424 585
R4524 GND.n4852 GND.n2424 585
R4525 GND.n2712 GND.n2553 585
R4526 GND.n2848 GND.n2553 585
R4527 GND.n2713 GND.n2565 585
R4528 GND.n2565 GND.n2552 585
R4529 GND.n2715 GND.n2714 585
R4530 GND.n2716 GND.n2715 585
R4531 GND.n2566 GND.n2564 585
R4532 GND.n2564 GND.n2560 585
R4533 GND.n2615 GND.n2614 585
R4534 GND.n2614 GND.n2613 585
R4535 GND.n2571 GND.n2570 585
R4536 GND.n2572 GND.n2571 585
R4537 GND.n2569 GND.n2466 585
R4538 GND.n2466 GND.n2463 585
R4539 GND.n2973 GND.n2972 585
R4540 GND.n2971 GND.n2465 585
R4541 GND.n2970 GND.n2464 585
R4542 GND.n2975 GND.n2464 585
R4543 GND.n2969 GND.n2968 585
R4544 GND.n2967 GND.n2966 585
R4545 GND.n2965 GND.n2964 585
R4546 GND.n2963 GND.n2962 585
R4547 GND.n2961 GND.n2960 585
R4548 GND.n2959 GND.n2958 585
R4549 GND.n2957 GND.n2956 585
R4550 GND.n2955 GND.n2954 585
R4551 GND.n2953 GND.n2952 585
R4552 GND.n2951 GND.n2950 585
R4553 GND.n2949 GND.n2948 585
R4554 GND.n2947 GND.n2946 585
R4555 GND.n2945 GND.n2944 585
R4556 GND.n2943 GND.n2942 585
R4557 GND.n2941 GND.n2940 585
R4558 GND.n2939 GND.n2938 585
R4559 GND.n2937 GND.n2936 585
R4560 GND.n2935 GND.n2489 585
R4561 GND.n2934 GND.n2933 585
R4562 GND.n2932 GND.n2931 585
R4563 GND.n2930 GND.n2929 585
R4564 GND.n2928 GND.n2927 585
R4565 GND.n2926 GND.n2925 585
R4566 GND.n2924 GND.n2923 585
R4567 GND.n2922 GND.n2921 585
R4568 GND.n2920 GND.n2919 585
R4569 GND.n2918 GND.n2917 585
R4570 GND.n2916 GND.n2915 585
R4571 GND.n2914 GND.n2913 585
R4572 GND.n2912 GND.n2911 585
R4573 GND.n2910 GND.n2909 585
R4574 GND.n2908 GND.n2907 585
R4575 GND.n2906 GND.n2905 585
R4576 GND.n2904 GND.n2903 585
R4577 GND.n2902 GND.n2901 585
R4578 GND.n2900 GND.n2899 585
R4579 GND.n2898 GND.n2897 585
R4580 GND.n2896 GND.n2895 585
R4581 GND.n2894 GND.n2893 585
R4582 GND.n2892 GND.n2516 585
R4583 GND.n2891 GND.n2890 585
R4584 GND.n2889 GND.n2888 585
R4585 GND.n2887 GND.n2886 585
R4586 GND.n2885 GND.n2884 585
R4587 GND.n2883 GND.n2882 585
R4588 GND.n2881 GND.n2880 585
R4589 GND.n2879 GND.n2878 585
R4590 GND.n2877 GND.n2876 585
R4591 GND.n2875 GND.n2874 585
R4592 GND.n2873 GND.n2872 585
R4593 GND.n2871 GND.n2870 585
R4594 GND.n2540 GND.n2530 585
R4595 GND.n1776 GND.n1629 585
R4596 GND.n1777 GND.n1775 585
R4597 GND.n1774 GND.n1771 585
R4598 GND.n1781 GND.n1770 585
R4599 GND.n1782 GND.n1769 585
R4600 GND.n1783 GND.n1768 585
R4601 GND.n1767 GND.n1765 585
R4602 GND.n1787 GND.n1764 585
R4603 GND.n1788 GND.n1763 585
R4604 GND.n1789 GND.n1762 585
R4605 GND.n1761 GND.n1759 585
R4606 GND.n1793 GND.n1758 585
R4607 GND.n1794 GND.n1757 585
R4608 GND.n1795 GND.n1753 585
R4609 GND.n1796 GND.n1752 585
R4610 GND.n1750 GND.n1749 585
R4611 GND.n1800 GND.n1748 585
R4612 GND.n1801 GND.n1747 585
R4613 GND.n1802 GND.n1746 585
R4614 GND.n1744 GND.n1743 585
R4615 GND.n1806 GND.n1742 585
R4616 GND.n1807 GND.n1741 585
R4617 GND.n1808 GND.n1740 585
R4618 GND.n1738 GND.n1737 585
R4619 GND.n1812 GND.n1734 585
R4620 GND.n1813 GND.n1733 585
R4621 GND.n1814 GND.n1732 585
R4622 GND.n1730 GND.n1729 585
R4623 GND.n1818 GND.n1728 585
R4624 GND.n6245 GND.n6244 585
R4625 GND.n6243 GND.n1726 585
R4626 GND.n6249 GND.n1725 585
R4627 GND.n6250 GND.n1724 585
R4628 GND.n6251 GND.n1720 585
R4629 GND.n6252 GND.n1719 585
R4630 GND.n1717 GND.n1716 585
R4631 GND.n6256 GND.n1715 585
R4632 GND.n6257 GND.n1714 585
R4633 GND.n6258 GND.n1713 585
R4634 GND.n1711 GND.n1710 585
R4635 GND.n6262 GND.n1709 585
R4636 GND.n6263 GND.n1708 585
R4637 GND.n6264 GND.n1707 585
R4638 GND.n1705 GND.n1704 585
R4639 GND.n6268 GND.n1701 585
R4640 GND.n6269 GND.n1700 585
R4641 GND.n6270 GND.n1699 585
R4642 GND.n1697 GND.n1696 585
R4643 GND.n6274 GND.n1695 585
R4644 GND.n6275 GND.n1694 585
R4645 GND.n6276 GND.n1693 585
R4646 GND.n1690 GND.n1689 585
R4647 GND.n6281 GND.n6280 585
R4648 GND.n6282 GND.n6281 585
R4649 GND.n6288 GND.n6287 585
R4650 GND.n6287 GND.n6286 585
R4651 GND.n1628 GND.n1627 585
R4652 GND.n1630 GND.n1628 585
R4653 GND.n5386 GND.n5385 585
R4654 GND.n5387 GND.n5386 585
R4655 GND.n1874 GND.n1873 585
R4656 GND.n1873 GND.n1869 585
R4657 GND.n5362 GND.n1881 585
R4658 GND.n5378 GND.n1881 585
R4659 GND.n1893 GND.n1891 585
R4660 GND.n1891 GND.n1878 585
R4661 GND.n5367 GND.n5366 585
R4662 GND.n5368 GND.n5367 585
R4663 GND.n1892 GND.n1890 585
R4664 GND.n5357 GND.n1890 585
R4665 GND.n5316 GND.n5315 585
R4666 GND.n5315 GND.n1897 585
R4667 GND.n5317 GND.n1907 585
R4668 GND.n5333 GND.n1907 585
R4669 GND.n1921 GND.n1919 585
R4670 GND.n1919 GND.n1904 585
R4671 GND.n5322 GND.n5321 585
R4672 GND.n5323 GND.n5322 585
R4673 GND.n1920 GND.n1918 585
R4674 GND.n1918 GND.n1914 585
R4675 GND.n5292 GND.n1928 585
R4676 GND.n5306 GND.n1928 585
R4677 GND.n1941 GND.n1939 585
R4678 GND.n1939 GND.n1925 585
R4679 GND.n5297 GND.n5296 585
R4680 GND.n5298 GND.n5297 585
R4681 GND.n1940 GND.n1938 585
R4682 GND.n1938 GND.n1934 585
R4683 GND.n5272 GND.n1948 585
R4684 GND.n5286 GND.n1948 585
R4685 GND.n1961 GND.n1959 585
R4686 GND.n1959 GND.n1945 585
R4687 GND.n5277 GND.n5276 585
R4688 GND.n5278 GND.n5277 585
R4689 GND.n1960 GND.n1958 585
R4690 GND.n1958 GND.n1954 585
R4691 GND.n5252 GND.n1968 585
R4692 GND.n5266 GND.n1968 585
R4693 GND.n1981 GND.n1979 585
R4694 GND.n1979 GND.n1965 585
R4695 GND.n5257 GND.n5256 585
R4696 GND.n5258 GND.n5257 585
R4697 GND.n1980 GND.n1978 585
R4698 GND.n1978 GND.n1974 585
R4699 GND.n5232 GND.n1988 585
R4700 GND.n5246 GND.n1988 585
R4701 GND.n2001 GND.n1999 585
R4702 GND.n1999 GND.n1985 585
R4703 GND.n5237 GND.n5236 585
R4704 GND.n5238 GND.n5237 585
R4705 GND.n2000 GND.n1998 585
R4706 GND.n1998 GND.n1994 585
R4707 GND.n5212 GND.n2008 585
R4708 GND.n5226 GND.n2008 585
R4709 GND.n2021 GND.n2019 585
R4710 GND.n2019 GND.n2005 585
R4711 GND.n5217 GND.n5216 585
R4712 GND.n5218 GND.n5217 585
R4713 GND.n2020 GND.n2018 585
R4714 GND.n2018 GND.n2014 585
R4715 GND.n5192 GND.n2028 585
R4716 GND.n5206 GND.n2028 585
R4717 GND.n2040 GND.n2038 585
R4718 GND.n2038 GND.n2025 585
R4719 GND.n5197 GND.n5196 585
R4720 GND.n5198 GND.n5197 585
R4721 GND.n2039 GND.n2037 585
R4722 GND.n5187 GND.n2037 585
R4723 GND.n5100 GND.n5099 585
R4724 GND.n5099 GND.n2044 585
R4725 GND.n5101 GND.n2054 585
R4726 GND.n5117 GND.n2054 585
R4727 GND.n2068 GND.n2066 585
R4728 GND.n2066 GND.n2051 585
R4729 GND.n5106 GND.n5105 585
R4730 GND.n5107 GND.n5106 585
R4731 GND.n2067 GND.n2065 585
R4732 GND.n2065 GND.n2061 585
R4733 GND.n5067 GND.n2075 585
R4734 GND.n5090 GND.n2075 585
R4735 GND.n5068 GND.n5065 585
R4736 GND.n5065 GND.n2072 585
R4737 GND.n5069 GND.n2201 585
R4738 GND.n5081 GND.n2201 585
R4739 GND.n2214 GND.n2212 585
R4740 GND.n2212 GND.n2198 585
R4741 GND.n5074 GND.n5073 585
R4742 GND.n5075 GND.n5074 585
R4743 GND.n2213 GND.n2211 585
R4744 GND.n2211 GND.n2205 585
R4745 GND.n5044 GND.n2223 585
R4746 GND.t34 GND.n2223 585
R4747 GND.n2237 GND.n2235 585
R4748 GND.n2235 GND.n2218 585
R4749 GND.n5049 GND.n5048 585
R4750 GND.n5050 GND.n5049 585
R4751 GND.n2236 GND.n2234 585
R4752 GND.n2234 GND.n2227 585
R4753 GND.n5023 GND.n2247 585
R4754 GND.n5038 GND.n2247 585
R4755 GND.n5024 GND.n5022 585
R4756 GND.n5022 GND.n2241 585
R4757 GND.n2260 GND.n2258 585
R4758 GND.n2258 GND.n2255 585
R4759 GND.n5029 GND.n5028 585
R4760 GND.n5030 GND.n5029 585
R4761 GND.n2259 GND.n2257 585
R4762 GND.n2257 GND.n2252 585
R4763 GND.n4998 GND.n2267 585
R4764 GND.n5013 GND.n2267 585
R4765 GND.n2280 GND.n2278 585
R4766 GND.n2278 GND.n2264 585
R4767 GND.n5003 GND.n5002 585
R4768 GND.n5004 GND.n5003 585
R4769 GND.n2279 GND.n2277 585
R4770 GND.n2277 GND.n2273 585
R4771 GND.n4978 GND.n2287 585
R4772 GND.n4992 GND.n2287 585
R4773 GND.n2300 GND.n2298 585
R4774 GND.n2298 GND.n2284 585
R4775 GND.n4983 GND.n4982 585
R4776 GND.n4984 GND.n4983 585
R4777 GND.n2299 GND.n2297 585
R4778 GND.n2297 GND.n2293 585
R4779 GND.n4958 GND.n2307 585
R4780 GND.n4972 GND.n2307 585
R4781 GND.n2320 GND.n2318 585
R4782 GND.n2318 GND.n2304 585
R4783 GND.n4963 GND.n4962 585
R4784 GND.n4964 GND.n4963 585
R4785 GND.n2319 GND.n2317 585
R4786 GND.n2317 GND.n2313 585
R4787 GND.n4938 GND.n2327 585
R4788 GND.n4952 GND.n2327 585
R4789 GND.n2340 GND.n2338 585
R4790 GND.n2338 GND.n2324 585
R4791 GND.n4943 GND.n4942 585
R4792 GND.n4944 GND.n4943 585
R4793 GND.n2339 GND.n2337 585
R4794 GND.n2337 GND.n2333 585
R4795 GND.n4918 GND.n2346 585
R4796 GND.n4932 GND.n2346 585
R4797 GND.n2360 GND.n2358 585
R4798 GND.n2358 GND.n2355 585
R4799 GND.n4923 GND.n4922 585
R4800 GND.n4924 GND.n4923 585
R4801 GND.n2359 GND.n2357 585
R4802 GND.n2357 GND.n2352 585
R4803 GND.n4898 GND.n2367 585
R4804 GND.n4912 GND.n2367 585
R4805 GND.n2380 GND.n2378 585
R4806 GND.n2378 GND.n2364 585
R4807 GND.n4903 GND.n4902 585
R4808 GND.n4904 GND.n4903 585
R4809 GND.n2379 GND.n2377 585
R4810 GND.n2377 GND.n2373 585
R4811 GND.n4878 GND.n2387 585
R4812 GND.n4892 GND.n2387 585
R4813 GND.n2400 GND.n2398 585
R4814 GND.n2398 GND.n2384 585
R4815 GND.n4883 GND.n4882 585
R4816 GND.n4884 GND.n4883 585
R4817 GND.n2399 GND.n2397 585
R4818 GND.n2397 GND.n2393 585
R4819 GND.n4858 GND.n2407 585
R4820 GND.n4872 GND.n2407 585
R4821 GND.n2420 GND.n2418 585
R4822 GND.n2418 GND.n2404 585
R4823 GND.n4863 GND.n4862 585
R4824 GND.n4864 GND.n4863 585
R4825 GND.n2419 GND.n2417 585
R4826 GND.n2417 GND.n2413 585
R4827 GND.n2851 GND.n2426 585
R4828 GND.n4852 GND.n2426 585
R4829 GND.n2852 GND.n2849 585
R4830 GND.n2849 GND.n2848 585
R4831 GND.n2853 GND.n2551 585
R4832 GND.n2552 GND.n2551 585
R4833 GND.n2561 GND.n2545 585
R4834 GND.n2716 GND.n2561 585
R4835 GND.n2857 GND.n2544 585
R4836 GND.n2560 GND.n2544 585
R4837 GND.n2858 GND.n2543 585
R4838 GND.n2613 GND.n2543 585
R4839 GND.n2859 GND.n2542 585
R4840 GND.n2572 GND.n2542 585
R4841 GND.n2541 GND.n2539 585
R4842 GND.n2541 GND.n2463 585
R4843 GND.n8323 GND.n384 585
R4844 GND.n384 GND.n350 585
R4845 GND.n8325 GND.n8324 585
R4846 GND.n8326 GND.n8325 585
R4847 GND.n454 GND.n453 585
R4848 GND.n453 GND.n449 585
R4849 GND.n8318 GND.n8317 585
R4850 GND.n8317 GND.n8316 585
R4851 GND.n8068 GND.n456 585
R4852 GND.n8069 GND.n8068 585
R4853 GND.n8067 GND.n8066 585
R4854 GND.n8067 GND.n342 585
R4855 GND.n457 GND.n340 585
R4856 GND.n8458 GND.n340 585
R4857 GND.n8062 GND.n8061 585
R4858 GND.n8061 GND.n332 585
R4859 GND.n8060 GND.n330 585
R4860 GND.n8464 GND.n330 585
R4861 GND.n8059 GND.n8058 585
R4862 GND.n8058 GND.n321 585
R4863 GND.n459 GND.n319 585
R4864 GND.n8470 GND.n319 585
R4865 GND.n8054 GND.n8053 585
R4866 GND.n8053 GND.n311 585
R4867 GND.n8052 GND.n309 585
R4868 GND.n8476 GND.n309 585
R4869 GND.n8051 GND.n8050 585
R4870 GND.n8050 GND.n300 585
R4871 GND.n461 GND.n298 585
R4872 GND.n8482 GND.n298 585
R4873 GND.n8046 GND.n8045 585
R4874 GND.n8045 GND.n290 585
R4875 GND.n8044 GND.n288 585
R4876 GND.n8488 GND.n288 585
R4877 GND.n8043 GND.n8042 585
R4878 GND.n8042 GND.n279 585
R4879 GND.n463 GND.n277 585
R4880 GND.n8494 GND.n277 585
R4881 GND.n8038 GND.n8037 585
R4882 GND.n8037 GND.n269 585
R4883 GND.n8036 GND.n267 585
R4884 GND.n8500 GND.n267 585
R4885 GND.n8035 GND.n8034 585
R4886 GND.n8034 GND.n258 585
R4887 GND.n465 GND.n256 585
R4888 GND.n8506 GND.n256 585
R4889 GND.n8030 GND.n8029 585
R4890 GND.n8029 GND.n248 585
R4891 GND.n8028 GND.n246 585
R4892 GND.n8512 GND.n246 585
R4893 GND.n8027 GND.n8026 585
R4894 GND.n8026 GND.n237 585
R4895 GND.n467 GND.n235 585
R4896 GND.n8518 GND.n235 585
R4897 GND.n8022 GND.n8021 585
R4898 GND.n8021 GND.n227 585
R4899 GND.n8020 GND.n225 585
R4900 GND.n8524 GND.n225 585
R4901 GND.n8019 GND.n8018 585
R4902 GND.n8018 GND.n216 585
R4903 GND.n469 GND.n214 585
R4904 GND.n8530 GND.n214 585
R4905 GND.n8014 GND.n8013 585
R4906 GND.n8013 GND.n206 585
R4907 GND.n8012 GND.n204 585
R4908 GND.n8536 GND.n204 585
R4909 GND.n8011 GND.n8010 585
R4910 GND.n8010 GND.n195 585
R4911 GND.n471 GND.n193 585
R4912 GND.n8542 GND.n193 585
R4913 GND.n8006 GND.n8005 585
R4914 GND.n8005 GND.n192 585
R4915 GND.n8004 GND.n183 585
R4916 GND.n8548 GND.n183 585
R4917 GND.n8003 GND.n8002 585
R4918 GND.n8002 GND.n174 585
R4919 GND.n473 GND.n172 585
R4920 GND.n8554 GND.n172 585
R4921 GND.n7998 GND.n7997 585
R4922 GND.n7997 GND.n164 585
R4923 GND.n7996 GND.n162 585
R4924 GND.n8560 GND.n162 585
R4925 GND.n7995 GND.n7994 585
R4926 GND.n7994 GND.n154 585
R4927 GND.n7991 GND.n152 585
R4928 GND.n8566 GND.n152 585
R4929 GND.n7990 GND.n7989 585
R4930 GND.n7989 GND.n142 585
R4931 GND.n7988 GND.n140 585
R4932 GND.n8572 GND.n140 585
R4933 GND.n7986 GND.n7985 585
R4934 GND.n7985 GND.n136 585
R4935 GND.n7984 GND.n135 585
R4936 GND.n8579 GND.n135 585
R4937 GND.n7982 GND.n7981 585
R4938 GND.n7981 GND.n71 585
R4939 GND.n7980 GND.n69 585
R4940 GND.t25 GND.n69 585
R4941 GND.n7978 GND.n7977 585
R4942 GND.n7977 GND.n68 585
R4943 GND.n7976 GND.n7975 585
R4944 GND.n7976 GND.n103 585
R4945 GND.n7973 GND.n101 585
R4946 GND.n8624 GND.n101 585
R4947 GND.n7972 GND.n7971 585
R4948 GND.n7971 GND.n91 585
R4949 GND.n7969 GND.n89 585
R4950 GND.n8630 GND.n89 585
R4951 GND.n7968 GND.n7967 585
R4952 GND.n7967 GND.n88 585
R4953 GND.n475 GND.n111 585
R4954 GND.n8608 GND.n111 585
R4955 GND.n7963 GND.n7962 585
R4956 GND.n7962 GND.n110 585
R4957 GND.n7961 GND.n120 585
R4958 GND.n8600 GND.n120 585
R4959 GND.n7960 GND.n7959 585
R4960 GND.n7959 GND.n119 585
R4961 GND.n7958 GND.n477 585
R4962 GND.n7958 GND.n7957 585
R4963 GND.n751 GND.n479 585
R4964 GND.n480 GND.n479 585
R4965 GND.n752 GND.n490 585
R4966 GND.n7949 GND.n490 585
R4967 GND.n754 GND.n753 585
R4968 GND.n753 GND.n489 585
R4969 GND.n755 GND.n502 585
R4970 GND.n7930 GND.n502 585
R4971 GND.n757 GND.n756 585
R4972 GND.n756 GND.n501 585
R4973 GND.n758 GND.n511 585
R4974 GND.n7922 GND.n511 585
R4975 GND.n760 GND.n759 585
R4976 GND.n759 GND.n510 585
R4977 GND.n761 GND.n522 585
R4978 GND.n7910 GND.n522 585
R4979 GND.n763 GND.n762 585
R4980 GND.n762 GND.n521 585
R4981 GND.n764 GND.n531 585
R4982 GND.n7902 GND.n531 585
R4983 GND.n766 GND.n765 585
R4984 GND.n765 GND.n530 585
R4985 GND.n767 GND.n542 585
R4986 GND.n7890 GND.n542 585
R4987 GND.n769 GND.n768 585
R4988 GND.n768 GND.n541 585
R4989 GND.n770 GND.n550 585
R4990 GND.n7882 GND.n550 585
R4991 GND.n771 GND.n561 585
R4992 GND.n7871 GND.n561 585
R4993 GND.n773 GND.n772 585
R4994 GND.n772 GND.n560 585
R4995 GND.n774 GND.n568 585
R4996 GND.n7818 GND.n568 585
R4997 GND.n776 GND.n775 585
R4998 GND.n775 GND.n567 585
R4999 GND.n777 GND.n578 585
R5000 GND.n7808 GND.n578 585
R5001 GND.n779 GND.n778 585
R5002 GND.n778 GND.n577 585
R5003 GND.n780 GND.n590 585
R5004 GND.n7792 GND.n590 585
R5005 GND.n782 GND.n781 585
R5006 GND.n781 GND.n589 585
R5007 GND.n783 GND.n599 585
R5008 GND.n7784 GND.n599 585
R5009 GND.n785 GND.n784 585
R5010 GND.n784 GND.n598 585
R5011 GND.n786 GND.n610 585
R5012 GND.n7772 GND.n610 585
R5013 GND.n788 GND.n787 585
R5014 GND.n787 GND.n609 585
R5015 GND.n789 GND.n619 585
R5016 GND.n7764 GND.n619 585
R5017 GND.n791 GND.n790 585
R5018 GND.n790 GND.n618 585
R5019 GND.n792 GND.n630 585
R5020 GND.n7752 GND.n630 585
R5021 GND.n794 GND.n793 585
R5022 GND.n793 GND.n629 585
R5023 GND.n795 GND.n639 585
R5024 GND.n7744 GND.n639 585
R5025 GND.n797 GND.n796 585
R5026 GND.n796 GND.n638 585
R5027 GND.n798 GND.n650 585
R5028 GND.n7732 GND.n650 585
R5029 GND.n800 GND.n799 585
R5030 GND.n799 GND.n649 585
R5031 GND.n801 GND.n659 585
R5032 GND.n7724 GND.n659 585
R5033 GND.n803 GND.n802 585
R5034 GND.n802 GND.n658 585
R5035 GND.n804 GND.n671 585
R5036 GND.n7710 GND.n671 585
R5037 GND.n7699 GND.n7698 585
R5038 GND.n7697 GND.n713 585
R5039 GND.n7696 GND.n712 585
R5040 GND.n7701 GND.n712 585
R5041 GND.n7695 GND.n7694 585
R5042 GND.n7693 GND.n7692 585
R5043 GND.n7691 GND.n7690 585
R5044 GND.n7689 GND.n7688 585
R5045 GND.n7687 GND.n7686 585
R5046 GND.n7685 GND.n7684 585
R5047 GND.n7683 GND.n7682 585
R5048 GND.n7681 GND.n7680 585
R5049 GND.n7679 GND.n7678 585
R5050 GND.n7677 GND.n7676 585
R5051 GND.n7675 GND.n7674 585
R5052 GND.n7673 GND.n7672 585
R5053 GND.n7671 GND.n7670 585
R5054 GND.n7669 GND.n7668 585
R5055 GND.n7667 GND.n7666 585
R5056 GND.n7665 GND.n7664 585
R5057 GND.n7663 GND.n7662 585
R5058 GND.n7661 GND.n828 585
R5059 GND.n7660 GND.n7659 585
R5060 GND.n7658 GND.n7657 585
R5061 GND.n7656 GND.n7655 585
R5062 GND.n7653 GND.n7652 585
R5063 GND.n7651 GND.n7650 585
R5064 GND.n7649 GND.n7648 585
R5065 GND.n7647 GND.n7646 585
R5066 GND.n7645 GND.n7644 585
R5067 GND.n7643 GND.n7642 585
R5068 GND.n7641 GND.n7640 585
R5069 GND.n7639 GND.n7638 585
R5070 GND.n7637 GND.n7636 585
R5071 GND.n7635 GND.n7634 585
R5072 GND.n7633 GND.n7632 585
R5073 GND.n7631 GND.n7630 585
R5074 GND.n7629 GND.n7628 585
R5075 GND.n7627 GND.n7626 585
R5076 GND.n7625 GND.n7624 585
R5077 GND.n7623 GND.n7622 585
R5078 GND.n7621 GND.n7580 585
R5079 GND.n7620 GND.n7619 585
R5080 GND.n7618 GND.n7617 585
R5081 GND.n7616 GND.n7615 585
R5082 GND.n7614 GND.n7613 585
R5083 GND.n7612 GND.n7611 585
R5084 GND.n7610 GND.n7609 585
R5085 GND.n7608 GND.n7607 585
R5086 GND.n7606 GND.n7605 585
R5087 GND.n7604 GND.n7603 585
R5088 GND.n7602 GND.n7601 585
R5089 GND.n7600 GND.n7599 585
R5090 GND.n7594 GND.n669 585
R5091 GND.n8328 GND.n441 585
R5092 GND.n8336 GND.n8335 585
R5093 GND.n8338 GND.n8337 585
R5094 GND.n8340 GND.n8339 585
R5095 GND.n8342 GND.n8341 585
R5096 GND.n8344 GND.n8343 585
R5097 GND.n8346 GND.n8345 585
R5098 GND.n8348 GND.n8347 585
R5099 GND.n8350 GND.n8349 585
R5100 GND.n8352 GND.n8351 585
R5101 GND.n8354 GND.n8353 585
R5102 GND.n431 GND.n428 585
R5103 GND.n8358 GND.n432 585
R5104 GND.n8360 GND.n8359 585
R5105 GND.n8362 GND.n8361 585
R5106 GND.n8364 GND.n8363 585
R5107 GND.n8366 GND.n8365 585
R5108 GND.n8368 GND.n8367 585
R5109 GND.n8370 GND.n8369 585
R5110 GND.n8372 GND.n8371 585
R5111 GND.n8374 GND.n8373 585
R5112 GND.n8377 GND.n8376 585
R5113 GND.n8375 GND.n417 585
R5114 GND.n8382 GND.n8381 585
R5115 GND.n8384 GND.n8383 585
R5116 GND.n8386 GND.n8385 585
R5117 GND.n8388 GND.n8387 585
R5118 GND.n8390 GND.n8389 585
R5119 GND.n8392 GND.n8391 585
R5120 GND.n8394 GND.n8393 585
R5121 GND.n8396 GND.n8395 585
R5122 GND.n8398 GND.n8397 585
R5123 GND.n8400 GND.n8399 585
R5124 GND.n407 GND.n404 585
R5125 GND.n8404 GND.n408 585
R5126 GND.n8406 GND.n8405 585
R5127 GND.n8408 GND.n8407 585
R5128 GND.n8410 GND.n8409 585
R5129 GND.n8412 GND.n8411 585
R5130 GND.n8414 GND.n8413 585
R5131 GND.n8416 GND.n8415 585
R5132 GND.n8418 GND.n8417 585
R5133 GND.n8420 GND.n8419 585
R5134 GND.n8423 GND.n8422 585
R5135 GND.n8421 GND.n393 585
R5136 GND.n8428 GND.n8427 585
R5137 GND.n8430 GND.n8429 585
R5138 GND.n8432 GND.n8431 585
R5139 GND.n8434 GND.n8433 585
R5140 GND.n8436 GND.n8435 585
R5141 GND.n8438 GND.n8437 585
R5142 GND.n8441 GND.n8440 585
R5143 GND.n8439 GND.n387 585
R5144 GND.n8445 GND.n385 585
R5145 GND.n8447 GND.n8446 585
R5146 GND.n8448 GND.n8447 585
R5147 GND.n8330 GND.n8329 585
R5148 GND.n8329 GND.n350 585
R5149 GND.n8327 GND.n447 585
R5150 GND.n8327 GND.n8326 585
R5151 GND.n8310 GND.n448 585
R5152 GND.n449 GND.n448 585
R5153 GND.n8309 GND.n8070 585
R5154 GND.n8316 GND.n8070 585
R5155 GND.n8308 GND.n8307 585
R5156 GND.n8307 GND.n8069 585
R5157 GND.n339 GND.n338 585
R5158 GND.n342 GND.n339 585
R5159 GND.n8460 GND.n8459 585
R5160 GND.n8459 GND.n8458 585
R5161 GND.n8461 GND.n334 585
R5162 GND.n334 GND.n332 585
R5163 GND.n8463 GND.n8462 585
R5164 GND.n8464 GND.n8463 585
R5165 GND.n318 GND.n317 585
R5166 GND.n321 GND.n318 585
R5167 GND.n8472 GND.n8471 585
R5168 GND.n8471 GND.n8470 585
R5169 GND.n8473 GND.n313 585
R5170 GND.n313 GND.n311 585
R5171 GND.n8475 GND.n8474 585
R5172 GND.n8476 GND.n8475 585
R5173 GND.n297 GND.n296 585
R5174 GND.n300 GND.n297 585
R5175 GND.n8484 GND.n8483 585
R5176 GND.n8483 GND.n8482 585
R5177 GND.n8485 GND.n292 585
R5178 GND.n292 GND.n290 585
R5179 GND.n8487 GND.n8486 585
R5180 GND.n8488 GND.n8487 585
R5181 GND.n276 GND.n275 585
R5182 GND.n279 GND.n276 585
R5183 GND.n8496 GND.n8495 585
R5184 GND.n8495 GND.n8494 585
R5185 GND.n8497 GND.n271 585
R5186 GND.n271 GND.n269 585
R5187 GND.n8499 GND.n8498 585
R5188 GND.n8500 GND.n8499 585
R5189 GND.n255 GND.n254 585
R5190 GND.n258 GND.n255 585
R5191 GND.n8508 GND.n8507 585
R5192 GND.n8507 GND.n8506 585
R5193 GND.n8509 GND.n250 585
R5194 GND.n250 GND.n248 585
R5195 GND.n8511 GND.n8510 585
R5196 GND.n8512 GND.n8511 585
R5197 GND.n234 GND.n233 585
R5198 GND.n237 GND.n234 585
R5199 GND.n8520 GND.n8519 585
R5200 GND.n8519 GND.n8518 585
R5201 GND.n8521 GND.n229 585
R5202 GND.n229 GND.n227 585
R5203 GND.n8523 GND.n8522 585
R5204 GND.n8524 GND.n8523 585
R5205 GND.n213 GND.n212 585
R5206 GND.n216 GND.n213 585
R5207 GND.n8532 GND.n8531 585
R5208 GND.n8531 GND.n8530 585
R5209 GND.n8533 GND.n208 585
R5210 GND.n208 GND.n206 585
R5211 GND.n8535 GND.n8534 585
R5212 GND.n8536 GND.n8535 585
R5213 GND.n191 GND.n190 585
R5214 GND.n195 GND.n191 585
R5215 GND.n8544 GND.n8543 585
R5216 GND.n8543 GND.n8542 585
R5217 GND.n8545 GND.n186 585
R5218 GND.n192 GND.n186 585
R5219 GND.n8547 GND.n8546 585
R5220 GND.n8548 GND.n8547 585
R5221 GND.n171 GND.n170 585
R5222 GND.n174 GND.n171 585
R5223 GND.n8556 GND.n8555 585
R5224 GND.n8555 GND.n8554 585
R5225 GND.n8557 GND.n166 585
R5226 GND.n166 GND.n164 585
R5227 GND.n8559 GND.n8558 585
R5228 GND.n8560 GND.n8559 585
R5229 GND.n151 GND.n150 585
R5230 GND.n154 GND.n151 585
R5231 GND.n8568 GND.n8567 585
R5232 GND.n8567 GND.n8566 585
R5233 GND.n8569 GND.n145 585
R5234 GND.n145 GND.n142 585
R5235 GND.n8571 GND.n8570 585
R5236 GND.n8572 GND.n8571 585
R5237 GND.n146 GND.n144 585
R5238 GND.n144 GND.n136 585
R5239 GND.n8232 GND.n138 585
R5240 GND.n8579 GND.n138 585
R5241 GND.n8231 GND.n8230 585
R5242 GND.n8230 GND.n71 585
R5243 GND.n8229 GND.n70 585
R5244 GND.t25 GND.n70 585
R5245 GND.n8228 GND.n8227 585
R5246 GND.n8227 GND.n68 585
R5247 GND.n100 GND.n99 585
R5248 GND.n103 GND.n100 585
R5249 GND.n8626 GND.n8625 585
R5250 GND.n8625 GND.n8624 585
R5251 GND.n8627 GND.n94 585
R5252 GND.n94 GND.n91 585
R5253 GND.n8629 GND.n8628 585
R5254 GND.n8630 GND.n8629 585
R5255 GND.n95 GND.n93 585
R5256 GND.n93 GND.n88 585
R5257 GND.n8596 GND.n113 585
R5258 GND.n8608 GND.n113 585
R5259 GND.n8597 GND.n124 585
R5260 GND.n124 GND.n110 585
R5261 GND.n8599 GND.n8598 585
R5262 GND.n8600 GND.n8599 585
R5263 GND.n125 GND.n123 585
R5264 GND.n123 GND.n119 585
R5265 GND.n7945 GND.n483 585
R5266 GND.n7957 GND.n483 585
R5267 GND.n7946 GND.n494 585
R5268 GND.n494 GND.n480 585
R5269 GND.n7948 GND.n7947 585
R5270 GND.n7949 GND.n7948 585
R5271 GND.n495 GND.n493 585
R5272 GND.n493 GND.n489 585
R5273 GND.n7918 GND.n504 585
R5274 GND.n7930 GND.n504 585
R5275 GND.n7919 GND.n515 585
R5276 GND.n515 GND.n501 585
R5277 GND.n7921 GND.n7920 585
R5278 GND.n7922 GND.n7921 585
R5279 GND.n516 GND.n514 585
R5280 GND.n514 GND.n510 585
R5281 GND.n7898 GND.n524 585
R5282 GND.n7910 GND.n524 585
R5283 GND.n7899 GND.n535 585
R5284 GND.n535 GND.n521 585
R5285 GND.n7901 GND.n7900 585
R5286 GND.n7902 GND.n7901 585
R5287 GND.n536 GND.n534 585
R5288 GND.n534 GND.n530 585
R5289 GND.n7878 GND.n544 585
R5290 GND.n7890 GND.n544 585
R5291 GND.n7879 GND.n554 585
R5292 GND.n554 GND.n541 585
R5293 GND.n7881 GND.n7880 585
R5294 GND.n7882 GND.n7881 585
R5295 GND.n555 GND.n553 585
R5296 GND.n7871 GND.n553 585
R5297 GND.n7803 GND.n7802 585
R5298 GND.n7802 GND.n560 585
R5299 GND.n7804 GND.n570 585
R5300 GND.n7818 GND.n570 585
R5301 GND.n7805 GND.n582 585
R5302 GND.n582 GND.n567 585
R5303 GND.n7807 GND.n7806 585
R5304 GND.n7808 GND.n7807 585
R5305 GND.n583 GND.n581 585
R5306 GND.n581 GND.n577 585
R5307 GND.n7780 GND.n592 585
R5308 GND.n7792 GND.n592 585
R5309 GND.n7781 GND.n603 585
R5310 GND.n603 GND.n589 585
R5311 GND.n7783 GND.n7782 585
R5312 GND.n7784 GND.n7783 585
R5313 GND.n604 GND.n602 585
R5314 GND.n602 GND.n598 585
R5315 GND.n7760 GND.n612 585
R5316 GND.n7772 GND.n612 585
R5317 GND.n7761 GND.n623 585
R5318 GND.n623 GND.n609 585
R5319 GND.n7763 GND.n7762 585
R5320 GND.n7764 GND.n7763 585
R5321 GND.n624 GND.n622 585
R5322 GND.n622 GND.n618 585
R5323 GND.n7740 GND.n632 585
R5324 GND.n7752 GND.n632 585
R5325 GND.n7741 GND.n643 585
R5326 GND.n643 GND.n629 585
R5327 GND.n7743 GND.n7742 585
R5328 GND.n7744 GND.n7743 585
R5329 GND.n644 GND.n642 585
R5330 GND.n642 GND.n638 585
R5331 GND.n7720 GND.n652 585
R5332 GND.n7732 GND.n652 585
R5333 GND.n7721 GND.n663 585
R5334 GND.n663 GND.n649 585
R5335 GND.n7723 GND.n7722 585
R5336 GND.n7724 GND.n7723 585
R5337 GND.n664 GND.n662 585
R5338 GND.n662 GND.n658 585
R5339 GND.n7712 GND.n7711 585
R5340 GND.n7711 GND.n7710 585
R5341 GND.n8457 GND.n8456 585
R5342 GND.n8458 GND.n8457 585
R5343 GND.n329 GND.n328 585
R5344 GND.n332 GND.n329 585
R5345 GND.n8466 GND.n8465 585
R5346 GND.n8465 GND.n8464 585
R5347 GND.n8467 GND.n323 585
R5348 GND.n323 GND.n321 585
R5349 GND.n8469 GND.n8468 585
R5350 GND.n8470 GND.n8469 585
R5351 GND.n308 GND.n307 585
R5352 GND.n311 GND.n308 585
R5353 GND.n8478 GND.n8477 585
R5354 GND.n8477 GND.n8476 585
R5355 GND.n8479 GND.n302 585
R5356 GND.n302 GND.n300 585
R5357 GND.n8481 GND.n8480 585
R5358 GND.n8482 GND.n8481 585
R5359 GND.n287 GND.n286 585
R5360 GND.n290 GND.n287 585
R5361 GND.n8490 GND.n8489 585
R5362 GND.n8489 GND.n8488 585
R5363 GND.n8491 GND.n281 585
R5364 GND.n281 GND.n279 585
R5365 GND.n8493 GND.n8492 585
R5366 GND.n8494 GND.n8493 585
R5367 GND.n266 GND.n265 585
R5368 GND.n269 GND.n266 585
R5369 GND.n8502 GND.n8501 585
R5370 GND.n8501 GND.n8500 585
R5371 GND.n8503 GND.n260 585
R5372 GND.n260 GND.n258 585
R5373 GND.n8505 GND.n8504 585
R5374 GND.n8506 GND.n8505 585
R5375 GND.n245 GND.n244 585
R5376 GND.n248 GND.n245 585
R5377 GND.n8514 GND.n8513 585
R5378 GND.n8513 GND.n8512 585
R5379 GND.n8515 GND.n239 585
R5380 GND.n239 GND.n237 585
R5381 GND.n8517 GND.n8516 585
R5382 GND.n8518 GND.n8517 585
R5383 GND.n224 GND.n223 585
R5384 GND.n227 GND.n224 585
R5385 GND.n8526 GND.n8525 585
R5386 GND.n8525 GND.n8524 585
R5387 GND.n8527 GND.n218 585
R5388 GND.n218 GND.n216 585
R5389 GND.n8529 GND.n8528 585
R5390 GND.n8530 GND.n8529 585
R5391 GND.n203 GND.n202 585
R5392 GND.n206 GND.n203 585
R5393 GND.n8538 GND.n8537 585
R5394 GND.n8537 GND.n8536 585
R5395 GND.n8539 GND.n197 585
R5396 GND.n197 GND.n195 585
R5397 GND.n8541 GND.n8540 585
R5398 GND.n8542 GND.n8541 585
R5399 GND.n182 GND.n181 585
R5400 GND.n192 GND.n182 585
R5401 GND.n8550 GND.n8549 585
R5402 GND.n8549 GND.n8548 585
R5403 GND.n8551 GND.n176 585
R5404 GND.n176 GND.n174 585
R5405 GND.n8553 GND.n8552 585
R5406 GND.n8554 GND.n8553 585
R5407 GND.n161 GND.n160 585
R5408 GND.n164 GND.n161 585
R5409 GND.n8562 GND.n8561 585
R5410 GND.n8561 GND.n8560 585
R5411 GND.n8563 GND.n156 585
R5412 GND.n156 GND.n154 585
R5413 GND.n8565 GND.n8564 585
R5414 GND.n8566 GND.n8565 585
R5415 GND.n157 GND.n139 585
R5416 GND.n142 GND.n139 585
R5417 GND.n8574 GND.n8573 585
R5418 GND.n8573 GND.n8572 585
R5419 GND.n8576 GND.n8575 585
R5420 GND.n8576 GND.n136 585
R5421 GND.n8578 GND.n8577 585
R5422 GND.n8579 GND.n8578 585
R5423 GND.n76 GND.n74 585
R5424 GND.n74 GND.n71 585
R5425 GND.n8636 GND.n8635 585
R5426 GND.t25 GND.n8636 585
R5427 GND.n75 GND.n73 585
R5428 GND.n73 GND.n68 585
R5429 GND.n8621 GND.n8620 585
R5430 GND.n8620 GND.n103 585
R5431 GND.n8623 GND.n8622 585
R5432 GND.n8624 GND.n8623 585
R5433 GND.n87 GND.n85 585
R5434 GND.n91 GND.n87 585
R5435 GND.n8632 GND.n8631 585
R5436 GND.n8631 GND.n8630 585
R5437 GND.n86 GND.n84 585
R5438 GND.n88 GND.n86 585
R5439 GND.n8607 GND.n8606 585
R5440 GND.n8608 GND.n8607 585
R5441 GND.n115 GND.n114 585
R5442 GND.n114 GND.n110 585
R5443 GND.n8602 GND.n8601 585
R5444 GND.n8601 GND.n8600 585
R5445 GND.n118 GND.n117 585
R5446 GND.n119 GND.n118 585
R5447 GND.n7956 GND.n7955 585
R5448 GND.n7957 GND.n7956 585
R5449 GND.n485 GND.n484 585
R5450 GND.n484 GND.n480 585
R5451 GND.n7951 GND.n7950 585
R5452 GND.n7950 GND.n7949 585
R5453 GND.n488 GND.n487 585
R5454 GND.n489 GND.n488 585
R5455 GND.n7929 GND.n7928 585
R5456 GND.n7930 GND.n7929 585
R5457 GND.n506 GND.n505 585
R5458 GND.n505 GND.n501 585
R5459 GND.n7924 GND.n7923 585
R5460 GND.n7923 GND.n7922 585
R5461 GND.n509 GND.n508 585
R5462 GND.n510 GND.n509 585
R5463 GND.n7909 GND.n7908 585
R5464 GND.n7910 GND.n7909 585
R5465 GND.n526 GND.n525 585
R5466 GND.n525 GND.n521 585
R5467 GND.n7904 GND.n7903 585
R5468 GND.n7903 GND.n7902 585
R5469 GND.n529 GND.n528 585
R5470 GND.n530 GND.n529 585
R5471 GND.n7889 GND.n7888 585
R5472 GND.n7890 GND.n7889 585
R5473 GND.n546 GND.n545 585
R5474 GND.n545 GND.n541 585
R5475 GND.n7884 GND.n7883 585
R5476 GND.n7883 GND.n7882 585
R5477 GND.n549 GND.n548 585
R5478 GND.n7871 GND.n549 585
R5479 GND.n7815 GND.n572 585
R5480 GND.n572 GND.n560 585
R5481 GND.n7817 GND.n7816 585
R5482 GND.n7818 GND.n7817 585
R5483 GND.n573 GND.n571 585
R5484 GND.n571 GND.n567 585
R5485 GND.n7810 GND.n7809 585
R5486 GND.n7809 GND.n7808 585
R5487 GND.n576 GND.n575 585
R5488 GND.n577 GND.n576 585
R5489 GND.n7791 GND.n7790 585
R5490 GND.n7792 GND.n7791 585
R5491 GND.n594 GND.n593 585
R5492 GND.n593 GND.n589 585
R5493 GND.n7786 GND.n7785 585
R5494 GND.n7785 GND.n7784 585
R5495 GND.n597 GND.n596 585
R5496 GND.n598 GND.n597 585
R5497 GND.n7771 GND.n7770 585
R5498 GND.n7772 GND.n7771 585
R5499 GND.n614 GND.n613 585
R5500 GND.n613 GND.n609 585
R5501 GND.n7766 GND.n7765 585
R5502 GND.n7765 GND.n7764 585
R5503 GND.n617 GND.n616 585
R5504 GND.n618 GND.n617 585
R5505 GND.n7751 GND.n7750 585
R5506 GND.n7752 GND.n7751 585
R5507 GND.n634 GND.n633 585
R5508 GND.n633 GND.n629 585
R5509 GND.n7746 GND.n7745 585
R5510 GND.n7745 GND.n7744 585
R5511 GND.n637 GND.n636 585
R5512 GND.n638 GND.n637 585
R5513 GND.n7731 GND.n7730 585
R5514 GND.n7732 GND.n7731 585
R5515 GND.n654 GND.n653 585
R5516 GND.n653 GND.n649 585
R5517 GND.n7726 GND.n7725 585
R5518 GND.n7725 GND.n7724 585
R5519 GND.n657 GND.n656 585
R5520 GND.n658 GND.n657 585
R5521 GND.n7709 GND.n7708 585
R5522 GND.n7710 GND.n7709 585
R5523 GND.n675 GND.n674 585
R5524 GND.n674 GND.n670 585
R5525 GND.n7704 GND.n7703 585
R5526 GND.n7703 GND.n7702 585
R5527 GND.n678 GND.n677 585
R5528 GND.n679 GND.n678 585
R5529 GND.n7496 GND.n7495 585
R5530 GND.n7497 GND.n7496 585
R5531 GND.n7499 GND.n7492 585
R5532 GND.n7499 GND.n7498 585
R5533 GND.n7501 GND.n7500 585
R5534 GND.n7500 GND.n851 585
R5535 GND.n7502 GND.n870 585
R5536 GND.n870 GND.n839 585
R5537 GND.n7504 GND.n7503 585
R5538 GND.n7505 GND.n7504 585
R5539 GND.n871 GND.n869 585
R5540 GND.n869 GND.n866 585
R5541 GND.n7486 GND.n7485 585
R5542 GND.n7485 GND.n7484 585
R5543 GND.n874 GND.n873 585
R5544 GND.n879 GND.n874 585
R5545 GND.n7421 GND.n7420 585
R5546 GND.n7422 GND.n7421 585
R5547 GND.n888 GND.n887 585
R5548 GND.n894 GND.n887 585
R5549 GND.n7416 GND.n7415 585
R5550 GND.n7415 GND.n7414 585
R5551 GND.n891 GND.n890 585
R5552 GND.n7407 GND.n891 585
R5553 GND.n7385 GND.n910 585
R5554 GND.n910 GND.n903 585
R5555 GND.n7387 GND.n7386 585
R5556 GND.n7388 GND.n7387 585
R5557 GND.n911 GND.n909 585
R5558 GND.n909 GND.n907 585
R5559 GND.n7380 GND.n7379 585
R5560 GND.n7379 GND.n7378 585
R5561 GND.n914 GND.n913 585
R5562 GND.n919 GND.n914 585
R5563 GND.n7361 GND.n7360 585
R5564 GND.n7362 GND.n7361 585
R5565 GND.n928 GND.n927 585
R5566 GND.n934 GND.n927 585
R5567 GND.n7356 GND.n7355 585
R5568 GND.n7355 GND.n7354 585
R5569 GND.n931 GND.n930 585
R5570 GND.n938 GND.n931 585
R5571 GND.n7326 GND.n952 585
R5572 GND.n952 GND.n945 585
R5573 GND.n7328 GND.n7327 585
R5574 GND.n7329 GND.n7328 585
R5575 GND.n953 GND.n951 585
R5576 GND.n951 GND.n949 585
R5577 GND.n7321 GND.n7320 585
R5578 GND.n7320 GND.n7319 585
R5579 GND.n956 GND.n955 585
R5580 GND.n7311 GND.n956 585
R5581 GND.n7290 GND.n7289 585
R5582 GND.n7289 GND.n969 585
R5583 GND.n7291 GND.n977 585
R5584 GND.n977 GND.n968 585
R5585 GND.n7293 GND.n7292 585
R5586 GND.n7294 GND.n7293 585
R5587 GND.n978 GND.n976 585
R5588 GND.n984 GND.n976 585
R5589 GND.n7283 GND.n7282 585
R5590 GND.n7282 GND.n7281 585
R5591 GND.n981 GND.n980 585
R5592 GND.n988 GND.n981 585
R5593 GND.n7253 GND.n1002 585
R5594 GND.n1002 GND.n995 585
R5595 GND.n7255 GND.n7254 585
R5596 GND.n7256 GND.n7255 585
R5597 GND.n1003 GND.n1001 585
R5598 GND.n1001 GND.n999 585
R5599 GND.n7248 GND.n7247 585
R5600 GND.n7247 GND.n7246 585
R5601 GND.n1006 GND.n1005 585
R5602 GND.n7238 GND.n1006 585
R5603 GND.n7200 GND.n7199 585
R5604 GND.n7200 GND.n1019 585
R5605 GND.n7201 GND.n7196 585
R5606 GND.n7201 GND.n1018 585
R5607 GND.n7203 GND.n7202 585
R5608 GND.n7202 GND.n1023 585
R5609 GND.n7204 GND.n1036 585
R5610 GND.n1036 GND.n1029 585
R5611 GND.n7206 GND.n7205 585
R5612 GND.n7207 GND.n7206 585
R5613 GND.n1037 GND.n1035 585
R5614 GND.n1035 GND.n1033 585
R5615 GND.n7190 GND.n7189 585
R5616 GND.n7189 GND.n7188 585
R5617 GND.n1040 GND.n1039 585
R5618 GND.n7180 GND.n1040 585
R5619 GND.n7158 GND.n7157 585
R5620 GND.n7157 GND.n1047 585
R5621 GND.n7159 GND.n1060 585
R5622 GND.n1060 GND.n1052 585
R5623 GND.n7161 GND.n7160 585
R5624 GND.n7162 GND.n7161 585
R5625 GND.n1061 GND.n1059 585
R5626 GND.n1067 GND.n1059 585
R5627 GND.n7151 GND.n7150 585
R5628 GND.n7150 GND.n7149 585
R5629 GND.n1064 GND.n1063 585
R5630 GND.n1071 GND.n1064 585
R5631 GND.n7121 GND.n1085 585
R5632 GND.n1085 GND.n1078 585
R5633 GND.n7123 GND.n7122 585
R5634 GND.n7124 GND.n7123 585
R5635 GND.n1086 GND.n1084 585
R5636 GND.n1084 GND.n1082 585
R5637 GND.n7116 GND.n7115 585
R5638 GND.n7115 GND.n7114 585
R5639 GND.n1089 GND.n1088 585
R5640 GND.n7106 GND.n1089 585
R5641 GND.n7068 GND.n7067 585
R5642 GND.n7068 GND.n1102 585
R5643 GND.n7069 GND.n7064 585
R5644 GND.n7069 GND.n1101 585
R5645 GND.n7071 GND.n7070 585
R5646 GND.n7070 GND.n1106 585
R5647 GND.n7072 GND.n1119 585
R5648 GND.n1119 GND.n1112 585
R5649 GND.n7074 GND.n7073 585
R5650 GND.n7075 GND.n7074 585
R5651 GND.n1120 GND.n1118 585
R5652 GND.n1118 GND.n1116 585
R5653 GND.n7058 GND.n7057 585
R5654 GND.n7057 GND.n7056 585
R5655 GND.n1123 GND.n1122 585
R5656 GND.n1132 GND.n1123 585
R5657 GND.n7020 GND.n7019 585
R5658 GND.n7020 GND.n1131 585
R5659 GND.n7022 GND.n7021 585
R5660 GND.n7021 GND.n1137 585
R5661 GND.n7023 GND.n1150 585
R5662 GND.n1150 GND.n1143 585
R5663 GND.n7025 GND.n7024 585
R5664 GND.n7026 GND.n7025 585
R5665 GND.n1151 GND.n1149 585
R5666 GND.n1149 GND.n1147 585
R5667 GND.n7012 GND.n7011 585
R5668 GND.n7011 GND.n7010 585
R5669 GND.n1154 GND.n1153 585
R5670 GND.n7002 GND.n1154 585
R5671 GND.n6900 GND.n6896 585
R5672 GND.n6896 GND.n1168 585
R5673 GND.n6902 GND.n6901 585
R5674 GND.n6902 GND.n1166 585
R5675 GND.n6903 GND.n6895 585
R5676 GND.n6903 GND.n1172 585
R5677 GND.n6905 GND.n6904 585
R5678 GND.n6904 GND.n1290 585
R5679 GND.n6906 GND.n1303 585
R5680 GND.n1303 GND.n1294 585
R5681 GND.n6908 GND.n6907 585
R5682 GND.n6909 GND.n6908 585
R5683 GND.n1304 GND.n1302 585
R5684 GND.n1320 GND.n1302 585
R5685 GND.n6889 GND.n6888 585
R5686 GND.n6888 GND.n6887 585
R5687 GND.n1307 GND.n1306 585
R5688 GND.n6880 GND.n1307 585
R5689 GND.n6735 GND.n6734 585
R5690 GND.n6734 GND.n1333 585
R5691 GND.n6736 GND.n6729 585
R5692 GND.n6729 GND.n1329 585
R5693 GND.n6738 GND.n6737 585
R5694 GND.n6738 GND.n1337 585
R5695 GND.n6739 GND.n6728 585
R5696 GND.n6739 GND.n1342 585
R5697 GND.n6742 GND.n6741 585
R5698 GND.n6741 GND.n6740 585
R5699 GND.n6743 GND.n6723 585
R5700 GND.n6723 GND.n1349 585
R5701 GND.n6745 GND.n6744 585
R5702 GND.n6745 GND.n1365 585
R5703 GND.n6747 GND.n6722 585
R5704 GND.n6747 GND.n6746 585
R5705 GND.n6749 GND.n6748 585
R5706 GND.n6748 GND.n1370 585
R5707 GND.n6750 GND.n1391 585
R5708 GND.n1391 GND.n1383 585
R5709 GND.n6752 GND.n6751 585
R5710 GND.n6753 GND.n6752 585
R5711 GND.n1392 GND.n1390 585
R5712 GND.n1390 GND.n1387 585
R5713 GND.n6716 GND.n6715 585
R5714 GND.n6715 GND.n6714 585
R5715 GND.n1395 GND.n1394 585
R5716 GND.n6706 GND.n1395 585
R5717 GND.n6692 GND.n6691 585
R5718 GND.n6693 GND.n6692 585
R5719 GND.n1415 GND.n1414 585
R5720 GND.n1451 GND.n1414 585
R5721 GND.n6687 GND.n6686 585
R5722 GND.n6686 GND.n6685 585
R5723 GND.n1418 GND.n1417 585
R5724 GND.n1457 GND.n1418 585
R5725 GND.n6615 GND.n6614 585
R5726 GND.n6614 GND.n1434 585
R5727 GND.n6616 GND.n1469 585
R5728 GND.n1469 GND.n1444 585
R5729 GND.n6618 GND.n6617 585
R5730 GND.n6619 GND.n6618 585
R5731 GND.n1470 GND.n1468 585
R5732 GND.n6588 GND.n1468 585
R5733 GND.n6608 GND.n6607 585
R5734 GND.n6607 GND.n6606 585
R5735 GND.n1473 GND.n1472 585
R5736 GND.n1485 GND.n1473 585
R5737 GND.n6538 GND.n6537 585
R5738 GND.n6538 GND.n1482 585
R5739 GND.n6540 GND.n6539 585
R5740 GND.n6539 GND.n1490 585
R5741 GND.n6541 GND.n1512 585
R5742 GND.n6518 GND.n1512 585
R5743 GND.n6543 GND.n6542 585
R5744 GND.n6544 GND.n6543 585
R5745 GND.n1513 GND.n1511 585
R5746 GND.n6509 GND.n1511 585
R5747 GND.n6530 GND.n6529 585
R5748 GND.n6529 GND.n6528 585
R5749 GND.n1516 GND.n1515 585
R5750 GND.n6503 GND.n1516 585
R5751 GND.n6477 GND.n6476 585
R5752 GND.n6476 GND.n1537 585
R5753 GND.n6478 GND.n1550 585
R5754 GND.n1550 GND.n1534 585
R5755 GND.n6480 GND.n6479 585
R5756 GND.n6481 GND.n6480 585
R5757 GND.n1551 GND.n1549 585
R5758 GND.n1558 GND.n1549 585
R5759 GND.n6470 GND.n6469 585
R5760 GND.n6469 GND.n6468 585
R5761 GND.n1554 GND.n1553 585
R5762 GND.n1563 GND.n1554 585
R5763 GND.n6438 GND.n1581 585
R5764 GND.n1581 GND.n1574 585
R5765 GND.n6440 GND.n6439 585
R5766 GND.n6441 GND.n6440 585
R5767 GND.n1582 GND.n1580 585
R5768 GND.n6415 GND.n1580 585
R5769 GND.n6433 GND.n6432 585
R5770 GND.n6432 GND.n6431 585
R5771 GND.n1585 GND.n1584 585
R5772 GND.n6423 GND.n1585 585
R5773 GND.n5957 GND.n5953 585
R5774 GND.n5953 GND.n5952 585
R5775 GND.n5959 GND.n5958 585
R5776 GND.n5960 GND.n5959 585
R5777 GND.n5922 GND.n5921 585
R5778 GND.n5925 GND.n5922 585
R5779 GND.n5970 GND.n5969 585
R5780 GND.n5969 GND.n5968 585
R5781 GND.n5971 GND.n5914 585
R5782 GND.n5937 GND.n5914 585
R5783 GND.n5973 GND.n5972 585
R5784 GND.n5974 GND.n5973 585
R5785 GND.n5915 GND.n5913 585
R5786 GND.n5913 GND.n5901 585
R5787 GND.n5844 GND.n5843 585
R5788 GND.n5900 GND.n5844 585
R5789 GND.n5989 GND.n5988 585
R5790 GND.n5988 GND.n5987 585
R5791 GND.n5990 GND.n5838 585
R5792 GND.n5845 GND.n5838 585
R5793 GND.n5992 GND.n5991 585
R5794 GND.n5993 GND.n5992 585
R5795 GND.n5826 GND.n5825 585
R5796 GND.n5829 GND.n5826 585
R5797 GND.n6003 GND.n6002 585
R5798 GND.n6002 GND.n6001 585
R5799 GND.n6004 GND.n5820 585
R5800 GND.n5884 GND.n5820 585
R5801 GND.n6006 GND.n6005 585
R5802 GND.n6007 GND.n6006 585
R5803 GND.n5808 GND.n5807 585
R5804 GND.n5811 GND.n5808 585
R5805 GND.n6017 GND.n6016 585
R5806 GND.n6016 GND.n6015 585
R5807 GND.n6018 GND.n5802 585
R5808 GND.n5871 GND.n5802 585
R5809 GND.n6020 GND.n6019 585
R5810 GND.n6021 GND.n6020 585
R5811 GND.n5791 GND.n5790 585
R5812 GND.n5794 GND.n5791 585
R5813 GND.n6031 GND.n6030 585
R5814 GND.n6030 GND.n6029 585
R5815 GND.n6032 GND.n5783 585
R5816 GND.n5857 GND.n5783 585
R5817 GND.n6034 GND.n6033 585
R5818 GND.n6035 GND.n6034 585
R5819 GND.n5784 GND.n5782 585
R5820 GND.n5782 GND.n5770 585
R5821 GND.n5714 GND.n5713 585
R5822 GND.n5769 GND.n5714 585
R5823 GND.n6050 GND.n6049 585
R5824 GND.n6049 GND.n6048 585
R5825 GND.n6051 GND.n5708 585
R5826 GND.n5715 GND.n5708 585
R5827 GND.n6053 GND.n6052 585
R5828 GND.n6054 GND.n6053 585
R5829 GND.n5696 GND.n5695 585
R5830 GND.n5699 GND.n5696 585
R5831 GND.n6064 GND.n6063 585
R5832 GND.n6063 GND.n6062 585
R5833 GND.n6065 GND.n5690 585
R5834 GND.n5753 GND.n5690 585
R5835 GND.n6067 GND.n6066 585
R5836 GND.n6068 GND.n6067 585
R5837 GND.n5678 GND.n5677 585
R5838 GND.n5681 GND.n5678 585
R5839 GND.n6078 GND.n6077 585
R5840 GND.n6077 GND.n6076 585
R5841 GND.n6079 GND.n5672 585
R5842 GND.n5740 GND.n5672 585
R5843 GND.n6081 GND.n6080 585
R5844 GND.n6082 GND.n6081 585
R5845 GND.n5660 GND.n5659 585
R5846 GND.n5663 GND.n5660 585
R5847 GND.n6092 GND.n6091 585
R5848 GND.n6091 GND.n6090 585
R5849 GND.n6093 GND.n5652 585
R5850 GND.n5727 GND.n5652 585
R5851 GND.n6095 GND.n6094 585
R5852 GND.n6096 GND.n6095 585
R5853 GND.n5653 GND.n5651 585
R5854 GND.n5651 GND.n5637 585
R5855 GND.n5583 GND.n5582 585
R5856 GND.n5636 GND.n5583 585
R5857 GND.n6111 GND.n6110 585
R5858 GND.n6110 GND.n6109 585
R5859 GND.n6112 GND.n5577 585
R5860 GND.n5640 GND.n5577 585
R5861 GND.n6114 GND.n6113 585
R5862 GND.n6115 GND.n6114 585
R5863 GND.n5565 GND.n5564 585
R5864 GND.n5568 GND.n5565 585
R5865 GND.n6125 GND.n6124 585
R5866 GND.n6124 GND.n6123 585
R5867 GND.n6126 GND.n5559 585
R5868 GND.n5620 GND.n5559 585
R5869 GND.n6128 GND.n6127 585
R5870 GND.n6129 GND.n6128 585
R5871 GND.n5547 GND.n5546 585
R5872 GND.n5550 GND.n5547 585
R5873 GND.n6139 GND.n6138 585
R5874 GND.n6138 GND.n6137 585
R5875 GND.n6140 GND.n5541 585
R5876 GND.n5607 GND.n5541 585
R5877 GND.n6142 GND.n6141 585
R5878 GND.n6143 GND.n6142 585
R5879 GND.n5529 GND.n5528 585
R5880 GND.n5532 GND.n5529 585
R5881 GND.n6153 GND.n6152 585
R5882 GND.n6152 GND.n6151 585
R5883 GND.n6154 GND.n5521 585
R5884 GND.n5594 GND.n5521 585
R5885 GND.n6156 GND.n6155 585
R5886 GND.n6157 GND.n6156 585
R5887 GND.n5522 GND.n5520 585
R5888 GND.n5520 GND.n5519 585
R5889 GND.n5433 GND.n5432 585
R5890 GND.n5507 GND.n5433 585
R5891 GND.n6172 GND.n6171 585
R5892 GND.n6171 GND.n6170 585
R5893 GND.n6173 GND.n5427 585
R5894 GND.n5434 GND.n5427 585
R5895 GND.n6175 GND.n6174 585
R5896 GND.n6176 GND.n6175 585
R5897 GND.n5415 GND.n5414 585
R5898 GND.n5418 GND.n5415 585
R5899 GND.n6186 GND.n6185 585
R5900 GND.n6185 GND.n6184 585
R5901 GND.n6187 GND.n1857 585
R5902 GND.n5491 GND.n1857 585
R5903 GND.n6189 GND.n6188 585
R5904 GND.n6190 GND.n6189 585
R5905 GND.n1858 GND.n1856 585
R5906 GND.n1856 GND.n1855 585
R5907 GND.n5408 GND.n5407 585
R5908 GND.n5407 GND.n1846 585
R5909 GND.n5406 GND.n1860 585
R5910 GND.n5406 GND.n1824 585
R5911 GND.n5405 GND.n5402 585
R5912 GND.n5405 GND.n5404 585
R5913 GND.n1862 GND.n1861 585
R5914 GND.n5403 GND.n1861 585
R5915 GND.n5398 GND.n5397 585
R5916 GND.n5397 GND.n1661 585
R5917 GND.n5396 GND.n1864 585
R5918 GND.n5396 GND.n1637 585
R5919 GND.n5395 GND.n5394 585
R5920 GND.n5395 GND.n1634 585
R5921 GND.n1865 GND.n1631 585
R5922 GND.n6286 GND.n1631 585
R5923 GND.n5390 GND.n5389 585
R5924 GND.n5389 GND.n1630 585
R5925 GND.n5388 GND.n1867 585
R5926 GND.n5388 GND.n5387 585
R5927 GND.n5375 GND.n1868 585
R5928 GND.n1869 GND.n1868 585
R5929 GND.n5377 GND.n5376 585
R5930 GND.n5378 GND.n5377 585
R5931 GND.n1883 GND.n1882 585
R5932 GND.n1882 GND.n1878 585
R5933 GND.n5370 GND.n5369 585
R5934 GND.n5369 GND.n5368 585
R5935 GND.n1886 GND.n1885 585
R5936 GND.n5357 GND.n1886 585
R5937 GND.n5330 GND.n1909 585
R5938 GND.n1909 GND.n1897 585
R5939 GND.n5332 GND.n5331 585
R5940 GND.n5333 GND.n5332 585
R5941 GND.n1910 GND.n1908 585
R5942 GND.n1908 GND.n1904 585
R5943 GND.n5325 GND.n5324 585
R5944 GND.n5324 GND.n5323 585
R5945 GND.n1913 GND.n1912 585
R5946 GND.n1914 GND.n1913 585
R5947 GND.n5305 GND.n5304 585
R5948 GND.n5306 GND.n5305 585
R5949 GND.n1930 GND.n1929 585
R5950 GND.n1929 GND.n1925 585
R5951 GND.n5300 GND.n5299 585
R5952 GND.n5299 GND.n5298 585
R5953 GND.n1933 GND.n1932 585
R5954 GND.n1934 GND.n1933 585
R5955 GND.n5285 GND.n5284 585
R5956 GND.n5286 GND.n5285 585
R5957 GND.n1950 GND.n1949 585
R5958 GND.n1949 GND.n1945 585
R5959 GND.n5280 GND.n5279 585
R5960 GND.n5279 GND.n5278 585
R5961 GND.n1953 GND.n1952 585
R5962 GND.n1954 GND.n1953 585
R5963 GND.n5265 GND.n5264 585
R5964 GND.n5266 GND.n5265 585
R5965 GND.n1970 GND.n1969 585
R5966 GND.n1969 GND.n1965 585
R5967 GND.n5260 GND.n5259 585
R5968 GND.n5259 GND.n5258 585
R5969 GND.n1973 GND.n1972 585
R5970 GND.n1974 GND.n1973 585
R5971 GND.n5245 GND.n5244 585
R5972 GND.n5246 GND.n5245 585
R5973 GND.n1990 GND.n1989 585
R5974 GND.n1989 GND.n1985 585
R5975 GND.n5240 GND.n5239 585
R5976 GND.n5239 GND.n5238 585
R5977 GND.n1993 GND.n1992 585
R5978 GND.n1994 GND.n1993 585
R5979 GND.n5225 GND.n5224 585
R5980 GND.n5226 GND.n5225 585
R5981 GND.n2010 GND.n2009 585
R5982 GND.n2009 GND.n2005 585
R5983 GND.n5220 GND.n5219 585
R5984 GND.n5219 GND.n5218 585
R5985 GND.n2013 GND.n2012 585
R5986 GND.n2014 GND.n2013 585
R5987 GND.n5205 GND.n5204 585
R5988 GND.n5206 GND.n5205 585
R5989 GND.n2030 GND.n2029 585
R5990 GND.n2029 GND.n2025 585
R5991 GND.n5200 GND.n5199 585
R5992 GND.n5199 GND.n5198 585
R5993 GND.n2033 GND.n2032 585
R5994 GND.n5187 GND.n2033 585
R5995 GND.n5114 GND.n2056 585
R5996 GND.n2056 GND.n2044 585
R5997 GND.n5116 GND.n5115 585
R5998 GND.n5117 GND.n5116 585
R5999 GND.n2057 GND.n2055 585
R6000 GND.n2055 GND.n2051 585
R6001 GND.n5109 GND.n5108 585
R6002 GND.n5108 GND.n5107 585
R6003 GND.n2060 GND.n2059 585
R6004 GND.n2061 GND.n2060 585
R6005 GND.n5089 GND.n5088 585
R6006 GND.n5090 GND.n5089 585
R6007 GND.n2077 GND.n2076 585
R6008 GND.n2076 GND.n2072 585
R6009 GND.n5080 GND.n5079 585
R6010 GND.n5081 GND.n5080 585
R6011 GND.n5078 GND.n5077 585
R6012 GND.n5077 GND.n2198 585
R6013 GND.n5076 GND.n2204 585
R6014 GND.n5076 GND.n5075 585
R6015 GND.n2203 GND.n2202 585
R6016 GND.n2205 GND.n2202 585
R6017 GND.n5055 GND.n5054 585
R6018 GND.t34 GND.n5055 585
R6019 GND.n5053 GND.n5052 585
R6020 GND.n5052 GND.n2218 585
R6021 GND.n5051 GND.n2226 585
R6022 GND.n5051 GND.n5050 585
R6023 GND.n2225 GND.n2084 585
R6024 GND.n2227 GND.n2225 585
R6025 GND.n5037 GND.n5036 585
R6026 GND.n5038 GND.n5037 585
R6027 GND.n5035 GND.n5034 585
R6028 GND.n5035 GND.n2241 585
R6029 GND.n5033 GND.n2248 585
R6030 GND.n2255 GND.n2248 585
R6031 GND.n5032 GND.n5031 585
R6032 GND.n5031 GND.n5030 585
R6033 GND.n2251 GND.n2249 585
R6034 GND.n2252 GND.n2251 585
R6035 GND.n5012 GND.n5011 585
R6036 GND.n5013 GND.n5012 585
R6037 GND.n2269 GND.n2268 585
R6038 GND.n2268 GND.n2264 585
R6039 GND.n5006 GND.n5005 585
R6040 GND.n5005 GND.n5004 585
R6041 GND.n2272 GND.n2271 585
R6042 GND.n2273 GND.n2272 585
R6043 GND.n4991 GND.n4990 585
R6044 GND.n4992 GND.n4991 585
R6045 GND.n2289 GND.n2288 585
R6046 GND.n2288 GND.n2284 585
R6047 GND.n4986 GND.n4985 585
R6048 GND.n4985 GND.n4984 585
R6049 GND.n2292 GND.n2291 585
R6050 GND.n2293 GND.n2292 585
R6051 GND.n4971 GND.n4970 585
R6052 GND.n4972 GND.n4971 585
R6053 GND.n2309 GND.n2308 585
R6054 GND.n2308 GND.n2304 585
R6055 GND.n4966 GND.n4965 585
R6056 GND.n4965 GND.n4964 585
R6057 GND.n2312 GND.n2311 585
R6058 GND.n2313 GND.n2312 585
R6059 GND.n4951 GND.n4950 585
R6060 GND.n4952 GND.n4951 585
R6061 GND.n2329 GND.n2328 585
R6062 GND.n2328 GND.n2324 585
R6063 GND.n4946 GND.n4945 585
R6064 GND.n4945 GND.n4944 585
R6065 GND.n2332 GND.n2331 585
R6066 GND.n2333 GND.n2332 585
R6067 GND.n4931 GND.n4930 585
R6068 GND.n4932 GND.n4931 585
R6069 GND.n2348 GND.n2347 585
R6070 GND.n2355 GND.n2347 585
R6071 GND.n4926 GND.n4925 585
R6072 GND.n4925 GND.n4924 585
R6073 GND.n2351 GND.n2350 585
R6074 GND.n2352 GND.n2351 585
R6075 GND.n4911 GND.n4910 585
R6076 GND.n4912 GND.n4911 585
R6077 GND.n2369 GND.n2368 585
R6078 GND.n2368 GND.n2364 585
R6079 GND.n4906 GND.n4905 585
R6080 GND.n4905 GND.n4904 585
R6081 GND.n2372 GND.n2371 585
R6082 GND.n2373 GND.n2372 585
R6083 GND.n4891 GND.n4890 585
R6084 GND.n4892 GND.n4891 585
R6085 GND.n2389 GND.n2388 585
R6086 GND.n2388 GND.n2384 585
R6087 GND.n4886 GND.n4885 585
R6088 GND.n4885 GND.n4884 585
R6089 GND.n2392 GND.n2391 585
R6090 GND.n2393 GND.n2392 585
R6091 GND.n4871 GND.n4870 585
R6092 GND.n4872 GND.n4871 585
R6093 GND.n2409 GND.n2408 585
R6094 GND.n2408 GND.n2404 585
R6095 GND.n4866 GND.n4865 585
R6096 GND.n4865 GND.n4864 585
R6097 GND.n2412 GND.n2411 585
R6098 GND.n2413 GND.n2412 585
R6099 GND.n4851 GND.n4850 585
R6100 GND.n4852 GND.n4851 585
R6101 GND.n2428 GND.n2427 585
R6102 GND.n2848 GND.n2427 585
R6103 GND.n6285 GND.n1626 585
R6104 GND.n6286 GND.n6285 585
R6105 GND.n5382 GND.n1635 585
R6106 GND.n1635 GND.n1630 585
R6107 GND.n5383 GND.n1871 585
R6108 GND.n5387 GND.n1871 585
R6109 GND.n5381 GND.n5380 585
R6110 GND.n5380 GND.n1869 585
R6111 GND.n5379 GND.n1876 585
R6112 GND.n5379 GND.n5378 585
R6113 GND.n5361 GND.n1877 585
R6114 GND.n1878 GND.n1877 585
R6115 GND.n5360 GND.n1888 585
R6116 GND.n5368 GND.n1888 585
R6117 GND.n5359 GND.n5358 585
R6118 GND.n5358 GND.n5357 585
R6119 GND.n1896 GND.n1895 585
R6120 GND.n1897 GND.n1896 585
R6121 GND.n5313 GND.n1906 585
R6122 GND.n5333 GND.n1906 585
R6123 GND.n5312 GND.n5311 585
R6124 GND.n5311 GND.n1904 585
R6125 GND.n5310 GND.n1916 585
R6126 GND.n5323 GND.n1916 585
R6127 GND.n5309 GND.n5308 585
R6128 GND.n5308 GND.n1914 585
R6129 GND.n5307 GND.n1923 585
R6130 GND.n5307 GND.n5306 585
R6131 GND.n5291 GND.n1924 585
R6132 GND.n1925 GND.n1924 585
R6133 GND.n5290 GND.n1936 585
R6134 GND.n5298 GND.n1936 585
R6135 GND.n5289 GND.n5288 585
R6136 GND.n5288 GND.n1934 585
R6137 GND.n5287 GND.n1943 585
R6138 GND.n5287 GND.n5286 585
R6139 GND.n5271 GND.n1944 585
R6140 GND.n1945 GND.n1944 585
R6141 GND.n5270 GND.n1956 585
R6142 GND.n5278 GND.n1956 585
R6143 GND.n5269 GND.n5268 585
R6144 GND.n5268 GND.n1954 585
R6145 GND.n5267 GND.n1963 585
R6146 GND.n5267 GND.n5266 585
R6147 GND.n5251 GND.n1964 585
R6148 GND.n1965 GND.n1964 585
R6149 GND.n5250 GND.n1976 585
R6150 GND.n5258 GND.n1976 585
R6151 GND.n5249 GND.n5248 585
R6152 GND.n5248 GND.n1974 585
R6153 GND.n5247 GND.n1983 585
R6154 GND.n5247 GND.n5246 585
R6155 GND.n5231 GND.n1984 585
R6156 GND.n1985 GND.n1984 585
R6157 GND.n5230 GND.n1996 585
R6158 GND.n5238 GND.n1996 585
R6159 GND.n5229 GND.n5228 585
R6160 GND.n5228 GND.n1994 585
R6161 GND.n5227 GND.n2003 585
R6162 GND.n5227 GND.n5226 585
R6163 GND.n5211 GND.n2004 585
R6164 GND.n2005 GND.n2004 585
R6165 GND.n5210 GND.n2016 585
R6166 GND.n5218 GND.n2016 585
R6167 GND.n5209 GND.n5208 585
R6168 GND.n5208 GND.n2014 585
R6169 GND.n5207 GND.n2023 585
R6170 GND.n5207 GND.n5206 585
R6171 GND.n5191 GND.n2024 585
R6172 GND.n2025 GND.n2024 585
R6173 GND.n5190 GND.n2035 585
R6174 GND.n5198 GND.n2035 585
R6175 GND.n5189 GND.n5188 585
R6176 GND.n5188 GND.n5187 585
R6177 GND.n2043 GND.n2042 585
R6178 GND.n2044 GND.n2043 585
R6179 GND.n5097 GND.n2053 585
R6180 GND.n5117 GND.n2053 585
R6181 GND.n5096 GND.n5095 585
R6182 GND.n5095 GND.n2051 585
R6183 GND.n5094 GND.n2063 585
R6184 GND.n5107 GND.n2063 585
R6185 GND.n5093 GND.n5092 585
R6186 GND.n5092 GND.n2061 585
R6187 GND.n5091 GND.n2070 585
R6188 GND.n5091 GND.n5090 585
R6189 GND.n5063 GND.n2071 585
R6190 GND.n2072 GND.n2071 585
R6191 GND.n5062 GND.n2199 585
R6192 GND.n5081 GND.n2199 585
R6193 GND.n5061 GND.n5060 585
R6194 GND.n5060 GND.n2198 585
R6195 GND.n5059 GND.n2209 585
R6196 GND.n5075 GND.n2209 585
R6197 GND.n5058 GND.n5057 585
R6198 GND.n5057 GND.n2205 585
R6199 GND.n5056 GND.n2216 585
R6200 GND.n5056 GND.t34 585
R6201 GND.n5043 GND.n2217 585
R6202 GND.n2218 GND.n2217 585
R6203 GND.n5042 GND.n2232 585
R6204 GND.n5050 GND.n2232 585
R6205 GND.n5041 GND.n5040 585
R6206 GND.n5040 GND.n2227 585
R6207 GND.n5039 GND.n2239 585
R6208 GND.n5039 GND.n5038 585
R6209 GND.n5020 GND.n2240 585
R6210 GND.n2241 GND.n2240 585
R6211 GND.n5019 GND.n5018 585
R6212 GND.n5018 GND.n2255 585
R6213 GND.n5017 GND.n2254 585
R6214 GND.n5030 GND.n2254 585
R6215 GND.n5016 GND.n5015 585
R6216 GND.n5015 GND.n2252 585
R6217 GND.n5014 GND.n2262 585
R6218 GND.n5014 GND.n5013 585
R6219 GND.n4997 GND.n2263 585
R6220 GND.n2264 GND.n2263 585
R6221 GND.n4996 GND.n2275 585
R6222 GND.n5004 GND.n2275 585
R6223 GND.n4995 GND.n4994 585
R6224 GND.n4994 GND.n2273 585
R6225 GND.n4993 GND.n2282 585
R6226 GND.n4993 GND.n4992 585
R6227 GND.n4977 GND.n2283 585
R6228 GND.n2284 GND.n2283 585
R6229 GND.n4976 GND.n2295 585
R6230 GND.n4984 GND.n2295 585
R6231 GND.n4975 GND.n4974 585
R6232 GND.n4974 GND.n2293 585
R6233 GND.n4973 GND.n2302 585
R6234 GND.n4973 GND.n4972 585
R6235 GND.n4957 GND.n2303 585
R6236 GND.n2304 GND.n2303 585
R6237 GND.n4956 GND.n2315 585
R6238 GND.n4964 GND.n2315 585
R6239 GND.n4955 GND.n4954 585
R6240 GND.n4954 GND.n2313 585
R6241 GND.n4953 GND.n2322 585
R6242 GND.n4953 GND.n4952 585
R6243 GND.n4937 GND.n2323 585
R6244 GND.n2324 GND.n2323 585
R6245 GND.n4936 GND.n2335 585
R6246 GND.n4944 GND.n2335 585
R6247 GND.n4935 GND.n4934 585
R6248 GND.n4934 GND.n2333 585
R6249 GND.n4933 GND.n2342 585
R6250 GND.n4933 GND.n4932 585
R6251 GND.n4917 GND.n2343 585
R6252 GND.n2355 GND.n2343 585
R6253 GND.n4916 GND.n2354 585
R6254 GND.n4924 GND.n2354 585
R6255 GND.n4915 GND.n4914 585
R6256 GND.n4914 GND.n2352 585
R6257 GND.n4913 GND.n2362 585
R6258 GND.n4913 GND.n4912 585
R6259 GND.n4897 GND.n2363 585
R6260 GND.n2364 GND.n2363 585
R6261 GND.n4896 GND.n2375 585
R6262 GND.n4904 GND.n2375 585
R6263 GND.n4895 GND.n4894 585
R6264 GND.n4894 GND.n2373 585
R6265 GND.n4893 GND.n2382 585
R6266 GND.n4893 GND.n4892 585
R6267 GND.n4877 GND.n2383 585
R6268 GND.n2384 GND.n2383 585
R6269 GND.n4876 GND.n2395 585
R6270 GND.n4884 GND.n2395 585
R6271 GND.n4875 GND.n4874 585
R6272 GND.n4874 GND.n2393 585
R6273 GND.n4873 GND.n2402 585
R6274 GND.n4873 GND.n4872 585
R6275 GND.n4857 GND.n2403 585
R6276 GND.n2404 GND.n2403 585
R6277 GND.n4856 GND.n2415 585
R6278 GND.n4864 GND.n2415 585
R6279 GND.n4855 GND.n4854 585
R6280 GND.n4854 GND.n2413 585
R6281 GND.n4853 GND.n2422 585
R6282 GND.n4853 GND.n4852 585
R6283 GND.n2549 GND.n2423 585
R6284 GND.n2848 GND.n2423 585
R6285 GND.n2562 GND.n2548 585
R6286 GND.n2562 GND.n2552 585
R6287 GND.n2563 GND.n2547 585
R6288 GND.n2716 GND.n2563 585
R6289 GND.n2611 GND.n2546 585
R6290 GND.n2611 GND.n2560 585
R6291 GND.n2612 GND.n2537 585
R6292 GND.n2613 GND.n2612 585
R6293 GND.n2861 GND.n2536 585
R6294 GND.n2572 GND.n2536 585
R6295 GND.n2863 GND.n2862 585
R6296 GND.n2863 GND.n2463 585
R6297 GND.n2865 GND.n2864 585
R6298 GND.n2586 GND.n2535 585
R6299 GND.n2588 GND.n2587 585
R6300 GND.n2584 GND.n2583 585
R6301 GND.n2592 GND.n2585 585
R6302 GND.n2594 GND.n2593 585
R6303 GND.n2596 GND.n2595 585
R6304 GND.n2580 GND.n2579 585
R6305 GND.n2600 GND.n2581 585
R6306 GND.n2601 GND.n2576 585
R6307 GND.n2602 GND.n2462 585
R6308 GND.n2975 GND.n2462 585
R6309 GND.n5345 GND.n1633 585
R6310 GND.n6286 GND.n1633 585
R6311 GND.n5347 GND.n5346 585
R6312 GND.n5346 GND.n1630 585
R6313 GND.n5348 GND.n1872 585
R6314 GND.n5387 GND.n1872 585
R6315 GND.n5350 GND.n5349 585
R6316 GND.n5349 GND.n1869 585
R6317 GND.n5351 GND.n1880 585
R6318 GND.n5378 GND.n1880 585
R6319 GND.n5353 GND.n5352 585
R6320 GND.n5352 GND.n1878 585
R6321 GND.n5354 GND.n1889 585
R6322 GND.n5368 GND.n1889 585
R6323 GND.n5356 GND.n5355 585
R6324 GND.n5357 GND.n5356 585
R6325 GND.n1900 GND.n1899 585
R6326 GND.n1899 GND.n1897 585
R6327 GND.n5335 GND.n5334 585
R6328 GND.n5334 GND.n5333 585
R6329 GND.n1903 GND.n1902 585
R6330 GND.n1904 GND.n1903 585
R6331 GND.n5148 GND.n1917 585
R6332 GND.n5323 GND.n1917 585
R6333 GND.n5150 GND.n5149 585
R6334 GND.n5149 GND.n1914 585
R6335 GND.n5151 GND.n1927 585
R6336 GND.n5306 GND.n1927 585
R6337 GND.n5153 GND.n5152 585
R6338 GND.n5152 GND.n1925 585
R6339 GND.n5154 GND.n1937 585
R6340 GND.n5298 GND.n1937 585
R6341 GND.n5156 GND.n5155 585
R6342 GND.n5155 GND.n1934 585
R6343 GND.n5157 GND.n1947 585
R6344 GND.n5286 GND.n1947 585
R6345 GND.n5159 GND.n5158 585
R6346 GND.n5158 GND.n1945 585
R6347 GND.n5160 GND.n1957 585
R6348 GND.n5278 GND.n1957 585
R6349 GND.n5162 GND.n5161 585
R6350 GND.n5161 GND.n1954 585
R6351 GND.n5163 GND.n1967 585
R6352 GND.n5266 GND.n1967 585
R6353 GND.n5165 GND.n5164 585
R6354 GND.n5164 GND.n1965 585
R6355 GND.n5166 GND.n1977 585
R6356 GND.n5258 GND.n1977 585
R6357 GND.n5168 GND.n5167 585
R6358 GND.n5167 GND.n1974 585
R6359 GND.n5169 GND.n1987 585
R6360 GND.n5246 GND.n1987 585
R6361 GND.n5171 GND.n5170 585
R6362 GND.n5170 GND.n1985 585
R6363 GND.n5172 GND.n1997 585
R6364 GND.n5238 GND.n1997 585
R6365 GND.n5174 GND.n5173 585
R6366 GND.n5173 GND.n1994 585
R6367 GND.n5175 GND.n2007 585
R6368 GND.n5226 GND.n2007 585
R6369 GND.n5177 GND.n5176 585
R6370 GND.n5176 GND.n2005 585
R6371 GND.n5178 GND.n2017 585
R6372 GND.n5218 GND.n2017 585
R6373 GND.n5180 GND.n5179 585
R6374 GND.n5179 GND.n2014 585
R6375 GND.n5181 GND.n2027 585
R6376 GND.n5206 GND.n2027 585
R6377 GND.n5183 GND.n5182 585
R6378 GND.n5182 GND.n2025 585
R6379 GND.n5184 GND.n2036 585
R6380 GND.n5198 GND.n2036 585
R6381 GND.n5186 GND.n5185 585
R6382 GND.n5187 GND.n5186 585
R6383 GND.n2047 GND.n2046 585
R6384 GND.n2046 GND.n2044 585
R6385 GND.n5119 GND.n5118 585
R6386 GND.n5118 GND.n5117 585
R6387 GND.n2050 GND.n2049 585
R6388 GND.n2051 GND.n2050 585
R6389 GND.n2770 GND.n2064 585
R6390 GND.n5107 GND.n2064 585
R6391 GND.n2772 GND.n2771 585
R6392 GND.n2771 GND.n2061 585
R6393 GND.n2773 GND.n2074 585
R6394 GND.n5090 GND.n2074 585
R6395 GND.n2775 GND.n2774 585
R6396 GND.n2774 GND.n2072 585
R6397 GND.n2776 GND.n2200 585
R6398 GND.n5081 GND.n2200 585
R6399 GND.n2778 GND.n2777 585
R6400 GND.n2777 GND.n2198 585
R6401 GND.n2779 GND.n2210 585
R6402 GND.n5075 GND.n2210 585
R6403 GND.n2781 GND.n2780 585
R6404 GND.n2780 GND.n2205 585
R6405 GND.n2762 GND.n2224 585
R6406 GND.t34 GND.n2224 585
R6407 GND.n2761 GND.n2760 585
R6408 GND.n2760 GND.n2218 585
R6409 GND.n2786 GND.n2233 585
R6410 GND.n5050 GND.n2233 585
R6411 GND.n2787 GND.n2759 585
R6412 GND.n2759 GND.n2227 585
R6413 GND.n2788 GND.n2246 585
R6414 GND.n5038 GND.n2246 585
R6415 GND.n2757 GND.n2756 585
R6416 GND.n2756 GND.n2241 585
R6417 GND.n2792 GND.n2755 585
R6418 GND.n2755 GND.n2255 585
R6419 GND.n2793 GND.n2256 585
R6420 GND.n5030 GND.n2256 585
R6421 GND.n2794 GND.n2754 585
R6422 GND.n2754 GND.n2252 585
R6423 GND.n2752 GND.n2266 585
R6424 GND.n5013 GND.n2266 585
R6425 GND.n2798 GND.n2751 585
R6426 GND.n2751 GND.n2264 585
R6427 GND.n2799 GND.n2276 585
R6428 GND.n5004 GND.n2276 585
R6429 GND.n2800 GND.n2750 585
R6430 GND.n2750 GND.n2273 585
R6431 GND.n2748 GND.n2286 585
R6432 GND.n4992 GND.n2286 585
R6433 GND.n2804 GND.n2747 585
R6434 GND.n2747 GND.n2284 585
R6435 GND.n2805 GND.n2296 585
R6436 GND.n4984 GND.n2296 585
R6437 GND.n2806 GND.n2746 585
R6438 GND.n2746 GND.n2293 585
R6439 GND.n2744 GND.n2306 585
R6440 GND.n4972 GND.n2306 585
R6441 GND.n2810 GND.n2743 585
R6442 GND.n2743 GND.n2304 585
R6443 GND.n2811 GND.n2316 585
R6444 GND.n4964 GND.n2316 585
R6445 GND.n2812 GND.n2742 585
R6446 GND.n2742 GND.n2313 585
R6447 GND.n2740 GND.n2326 585
R6448 GND.n4952 GND.n2326 585
R6449 GND.n2816 GND.n2739 585
R6450 GND.n2739 GND.n2324 585
R6451 GND.n2817 GND.n2336 585
R6452 GND.n4944 GND.n2336 585
R6453 GND.n2818 GND.n2738 585
R6454 GND.n2738 GND.n2333 585
R6455 GND.n2736 GND.n2345 585
R6456 GND.n4932 GND.n2345 585
R6457 GND.n2822 GND.n2735 585
R6458 GND.n2735 GND.n2355 585
R6459 GND.n2823 GND.n2356 585
R6460 GND.n4924 GND.n2356 585
R6461 GND.n2824 GND.n2734 585
R6462 GND.n2734 GND.n2352 585
R6463 GND.n2732 GND.n2366 585
R6464 GND.n4912 GND.n2366 585
R6465 GND.n2828 GND.n2731 585
R6466 GND.n2731 GND.n2364 585
R6467 GND.n2829 GND.n2376 585
R6468 GND.n4904 GND.n2376 585
R6469 GND.n2830 GND.n2730 585
R6470 GND.n2730 GND.n2373 585
R6471 GND.n2728 GND.n2386 585
R6472 GND.n4892 GND.n2386 585
R6473 GND.n2834 GND.n2727 585
R6474 GND.n2727 GND.n2384 585
R6475 GND.n2835 GND.n2396 585
R6476 GND.n4884 GND.n2396 585
R6477 GND.n2836 GND.n2726 585
R6478 GND.n2726 GND.n2393 585
R6479 GND.n2724 GND.n2406 585
R6480 GND.n4872 GND.n2406 585
R6481 GND.n2840 GND.n2723 585
R6482 GND.n2723 GND.n2404 585
R6483 GND.n2841 GND.n2416 585
R6484 GND.n4864 GND.n2416 585
R6485 GND.n2842 GND.n2722 585
R6486 GND.n2722 GND.n2413 585
R6487 GND.n2556 GND.n2425 585
R6488 GND.n4852 GND.n2425 585
R6489 GND.n2847 GND.n2846 585
R6490 GND.n2848 GND.n2847 585
R6491 GND.n2555 GND.n2554 585
R6492 GND.n2554 GND.n2552 585
R6493 GND.n2718 GND.n2717 585
R6494 GND.n2717 GND.n2716 585
R6495 GND.n2559 GND.n2558 585
R6496 GND.n2560 GND.n2559 585
R6497 GND.n2610 GND.n2609 585
R6498 GND.n2613 GND.n2610 585
R6499 GND.n2574 GND.n2573 585
R6500 GND.n2573 GND.n2572 585
R6501 GND.n2605 GND.n2604 585
R6502 GND.n2604 GND.n2463 585
R6503 GND.n6282 GND.n1660 585
R6504 GND.n1659 GND.n1658 585
R6505 GND.n1654 GND.n1622 585
R6506 GND.n1653 GND.n1652 585
R6507 GND.n1650 GND.n1649 585
R6508 GND.n1648 GND.n1647 585
R6509 GND.n1645 GND.n1644 585
R6510 GND.n1643 GND.n1642 585
R6511 GND.n1640 GND.n1639 585
R6512 GND.n1638 GND.n1636 585
R6513 GND.n7555 GND.n862 550.159
R6514 GND.n7477 GND.n868 550.159
R6515 GND.n5486 GND.n1845 550.159
R6516 GND.n6235 GND.n1849 550.159
R6517 GND.n4722 GND.n3026 280.613
R6518 GND.n4722 GND.n4721 280.613
R6519 GND.n4721 GND.n4720 280.613
R6520 GND.n4720 GND.n3027 280.613
R6521 GND.n4714 GND.n3027 280.613
R6522 GND.n4714 GND.n4713 280.613
R6523 GND.n4713 GND.n4712 280.613
R6524 GND.n4712 GND.n3035 280.613
R6525 GND.n4706 GND.n3035 280.613
R6526 GND.n4706 GND.n4705 280.613
R6527 GND.n4705 GND.n4704 280.613
R6528 GND.n4704 GND.n3043 280.613
R6529 GND.n4698 GND.n3043 280.613
R6530 GND.n4698 GND.n4697 280.613
R6531 GND.n4697 GND.n4696 280.613
R6532 GND.n4696 GND.n3051 280.613
R6533 GND.n4690 GND.n3051 280.613
R6534 GND.n4690 GND.n4689 280.613
R6535 GND.n4689 GND.n4688 280.613
R6536 GND.n4688 GND.n3059 280.613
R6537 GND.n4682 GND.n3059 280.613
R6538 GND.n4682 GND.n4681 280.613
R6539 GND.n4681 GND.n4680 280.613
R6540 GND.n4680 GND.n3067 280.613
R6541 GND.n4674 GND.n3067 280.613
R6542 GND.n4674 GND.n4673 280.613
R6543 GND.n4673 GND.n4672 280.613
R6544 GND.n4672 GND.n3075 280.613
R6545 GND.n4666 GND.n3075 280.613
R6546 GND.n4666 GND.n4665 280.613
R6547 GND.n4665 GND.n4664 280.613
R6548 GND.n4664 GND.n3083 280.613
R6549 GND.n4658 GND.n3083 280.613
R6550 GND.n4658 GND.n4657 280.613
R6551 GND.n4657 GND.n4656 280.613
R6552 GND.n4656 GND.n3091 280.613
R6553 GND.n4650 GND.n3091 280.613
R6554 GND.n4650 GND.n4649 280.613
R6555 GND.n4649 GND.n4648 280.613
R6556 GND.n4648 GND.n3099 280.613
R6557 GND.n4642 GND.n3099 280.613
R6558 GND.n4642 GND.n4641 280.613
R6559 GND.n4641 GND.n4640 280.613
R6560 GND.n4640 GND.n3107 280.613
R6561 GND.n4634 GND.n3107 280.613
R6562 GND.n4634 GND.n4633 280.613
R6563 GND.n4633 GND.n4632 280.613
R6564 GND.n4632 GND.n3115 280.613
R6565 GND.n4626 GND.n3115 280.613
R6566 GND.n4626 GND.n4625 280.613
R6567 GND.n4625 GND.n4624 280.613
R6568 GND.n4624 GND.n3123 280.613
R6569 GND.n4618 GND.n3123 280.613
R6570 GND.n4618 GND.n4617 280.613
R6571 GND.n4617 GND.n4616 280.613
R6572 GND.n4616 GND.n3131 280.613
R6573 GND.n4610 GND.n3131 280.613
R6574 GND.n4610 GND.n4609 280.613
R6575 GND.n4609 GND.n4608 280.613
R6576 GND.n4608 GND.n3139 280.613
R6577 GND.n4602 GND.n3139 280.613
R6578 GND.n4602 GND.n4601 280.613
R6579 GND.n4601 GND.n4600 280.613
R6580 GND.n4600 GND.n3147 280.613
R6581 GND.n4594 GND.n3147 280.613
R6582 GND.n4594 GND.n4593 280.613
R6583 GND.n4593 GND.n4592 280.613
R6584 GND.n4592 GND.n3155 280.613
R6585 GND.n4586 GND.n3155 280.613
R6586 GND.n4586 GND.n4585 280.613
R6587 GND.n4585 GND.n4584 280.613
R6588 GND.n4584 GND.n3163 280.613
R6589 GND.n4578 GND.n3163 280.613
R6590 GND.n4578 GND.n4577 280.613
R6591 GND.n4577 GND.n4576 280.613
R6592 GND.n4576 GND.n3171 280.613
R6593 GND.n4570 GND.n3171 280.613
R6594 GND.n4570 GND.n4569 280.613
R6595 GND.n4569 GND.n4568 280.613
R6596 GND.n4568 GND.n3179 280.613
R6597 GND.n4562 GND.n3179 280.613
R6598 GND.n4562 GND.n4561 280.613
R6599 GND.n4561 GND.n4560 280.613
R6600 GND.n4560 GND.n3187 280.613
R6601 GND.n4554 GND.n3187 280.613
R6602 GND.n4554 GND.n4553 280.613
R6603 GND.n4553 GND.n4552 280.613
R6604 GND.n4552 GND.n3195 280.613
R6605 GND.n4546 GND.n3195 280.613
R6606 GND.n4546 GND.n4545 280.613
R6607 GND.n4545 GND.n4544 280.613
R6608 GND.n4544 GND.n3203 280.613
R6609 GND.n4538 GND.n3203 280.613
R6610 GND.n4538 GND.n4537 280.613
R6611 GND.n4537 GND.n4536 280.613
R6612 GND.n4536 GND.n3211 280.613
R6613 GND.n4530 GND.n3211 280.613
R6614 GND.n4530 GND.n4529 280.613
R6615 GND.n4529 GND.n4528 280.613
R6616 GND.n4528 GND.n3219 280.613
R6617 GND.n4522 GND.n3219 280.613
R6618 GND.n4522 GND.n4521 280.613
R6619 GND.n4521 GND.n4520 280.613
R6620 GND.n4520 GND.n3227 280.613
R6621 GND.n4514 GND.n3227 280.613
R6622 GND.n4514 GND.n4513 280.613
R6623 GND.n4513 GND.n4512 280.613
R6624 GND.n4512 GND.n3235 280.613
R6625 GND.n4506 GND.n3235 280.613
R6626 GND.n4506 GND.n4505 280.613
R6627 GND.n4505 GND.n4504 280.613
R6628 GND.n4504 GND.n3243 280.613
R6629 GND.n4498 GND.n3243 280.613
R6630 GND.n4498 GND.n4497 280.613
R6631 GND.n4497 GND.n4496 280.613
R6632 GND.n4496 GND.n3251 280.613
R6633 GND.n4490 GND.n3251 280.613
R6634 GND.n4490 GND.n4489 280.613
R6635 GND.n4489 GND.n4488 280.613
R6636 GND.n4488 GND.n3259 280.613
R6637 GND.n4482 GND.n3259 280.613
R6638 GND.n4482 GND.n4481 280.613
R6639 GND.n4481 GND.n4480 280.613
R6640 GND.n4480 GND.n3267 280.613
R6641 GND.n4474 GND.n3267 280.613
R6642 GND.n4474 GND.n4473 280.613
R6643 GND.n4473 GND.n4472 280.613
R6644 GND.n4472 GND.n3275 280.613
R6645 GND.n4466 GND.n3275 280.613
R6646 GND.n4466 GND.n4465 280.613
R6647 GND.n4465 GND.n4464 280.613
R6648 GND.n4464 GND.n3283 280.613
R6649 GND.n4458 GND.n3283 280.613
R6650 GND.n4458 GND.n4457 280.613
R6651 GND.n4457 GND.n4456 280.613
R6652 GND.n4456 GND.n3291 280.613
R6653 GND.n4450 GND.n3291 280.613
R6654 GND.n4450 GND.n4449 280.613
R6655 GND.n4449 GND.n4448 280.613
R6656 GND.n4448 GND.n3299 280.613
R6657 GND.n4442 GND.n3299 280.613
R6658 GND.n4442 GND.n4441 280.613
R6659 GND.n4441 GND.n4440 280.613
R6660 GND.n4440 GND.n3307 280.613
R6661 GND.n4434 GND.n3307 280.613
R6662 GND.n4434 GND.n4433 280.613
R6663 GND.n4433 GND.n4432 280.613
R6664 GND.n4432 GND.n3315 280.613
R6665 GND.n4426 GND.n3315 280.613
R6666 GND.n4426 GND.n4425 280.613
R6667 GND.n4425 GND.n4424 280.613
R6668 GND.n4424 GND.n3323 280.613
R6669 GND.n4418 GND.n3323 280.613
R6670 GND.n4418 GND.n4417 280.613
R6671 GND.n4417 GND.n4416 280.613
R6672 GND.n4416 GND.n3331 280.613
R6673 GND.n4410 GND.n3331 280.613
R6674 GND.n4410 GND.n4409 280.613
R6675 GND.n4409 GND.n4408 280.613
R6676 GND.n4408 GND.n3339 280.613
R6677 GND.n4402 GND.n3339 280.613
R6678 GND.n4402 GND.n4401 280.613
R6679 GND.n4401 GND.n4400 280.613
R6680 GND.n4400 GND.n3347 280.613
R6681 GND.n4394 GND.n3347 280.613
R6682 GND.n4394 GND.n4393 280.613
R6683 GND.n4393 GND.n4392 280.613
R6684 GND.n4392 GND.n3355 280.613
R6685 GND.n4386 GND.n3355 280.613
R6686 GND.n4386 GND.n4385 280.613
R6687 GND.n4385 GND.n4384 280.613
R6688 GND.n4384 GND.n3363 280.613
R6689 GND.n4378 GND.n3363 280.613
R6690 GND.n4378 GND.n4377 280.613
R6691 GND.n4377 GND.n4376 280.613
R6692 GND.n4376 GND.n3371 280.613
R6693 GND.n4370 GND.n3371 280.613
R6694 GND.n4370 GND.n4369 280.613
R6695 GND.n4369 GND.n4368 280.613
R6696 GND.n4368 GND.n3379 280.613
R6697 GND.n4362 GND.n3379 280.613
R6698 GND.n4362 GND.n4361 280.613
R6699 GND.n4361 GND.n4360 280.613
R6700 GND.n4360 GND.n3387 280.613
R6701 GND.n4354 GND.n3387 280.613
R6702 GND.n4354 GND.n4353 280.613
R6703 GND.n4353 GND.n4352 280.613
R6704 GND.n4352 GND.n3395 280.613
R6705 GND.n4346 GND.n3395 280.613
R6706 GND.n4346 GND.n4345 280.613
R6707 GND.n4345 GND.n4344 280.613
R6708 GND.n4344 GND.n3403 280.613
R6709 GND.n4338 GND.n3403 280.613
R6710 GND.n4338 GND.n4337 280.613
R6711 GND.n4337 GND.n4336 280.613
R6712 GND.n4336 GND.n3411 280.613
R6713 GND.n4330 GND.n3411 280.613
R6714 GND.n4330 GND.n4329 280.613
R6715 GND.n4329 GND.n4328 280.613
R6716 GND.n4328 GND.n3419 280.613
R6717 GND.n4322 GND.n3419 280.613
R6718 GND.n4322 GND.n4321 280.613
R6719 GND.n4321 GND.n4320 280.613
R6720 GND.n4320 GND.n3427 280.613
R6721 GND.n4314 GND.n3427 280.613
R6722 GND.n4314 GND.n4313 280.613
R6723 GND.n4313 GND.n4312 280.613
R6724 GND.n4312 GND.n3435 280.613
R6725 GND.n4306 GND.n3435 280.613
R6726 GND.n4306 GND.n4305 280.613
R6727 GND.n4305 GND.n4304 280.613
R6728 GND.n4304 GND.n3443 280.613
R6729 GND.n4298 GND.n3443 280.613
R6730 GND.n4298 GND.n4297 280.613
R6731 GND.n4297 GND.n4296 280.613
R6732 GND.n4296 GND.n3451 280.613
R6733 GND.n4290 GND.n3451 280.613
R6734 GND.n4290 GND.n4289 280.613
R6735 GND.n4289 GND.n4288 280.613
R6736 GND.n4288 GND.n3459 280.613
R6737 GND.n4282 GND.n3459 280.613
R6738 GND.n4282 GND.n4281 280.613
R6739 GND.n4281 GND.n4280 280.613
R6740 GND.n4280 GND.n3467 280.613
R6741 GND.n4274 GND.n3467 280.613
R6742 GND.n4274 GND.n4273 280.613
R6743 GND.n4273 GND.n4272 280.613
R6744 GND.n4272 GND.n3475 280.613
R6745 GND.n4266 GND.n3475 280.613
R6746 GND.n4266 GND.n4265 280.613
R6747 GND.n4265 GND.n4264 280.613
R6748 GND.n4264 GND.n3483 280.613
R6749 GND.n4258 GND.n3483 280.613
R6750 GND.n4258 GND.n4257 280.613
R6751 GND.n4257 GND.n4256 280.613
R6752 GND.n4256 GND.n3491 280.613
R6753 GND.n4250 GND.n3491 280.613
R6754 GND.n4250 GND.n4249 280.613
R6755 GND.n4249 GND.n4248 280.613
R6756 GND.n4248 GND.n3499 280.613
R6757 GND.n4242 GND.n3499 280.613
R6758 GND.n4242 GND.n4241 280.613
R6759 GND.n4241 GND.n4240 280.613
R6760 GND.n4240 GND.n3507 280.613
R6761 GND.n4234 GND.n3507 280.613
R6762 GND.n4234 GND.n4233 280.613
R6763 GND.n4233 GND.n4232 280.613
R6764 GND.n4232 GND.n3515 280.613
R6765 GND.n4226 GND.n3515 280.613
R6766 GND.n4226 GND.n4225 280.613
R6767 GND.n4225 GND.n4224 280.613
R6768 GND.n4224 GND.n3523 280.613
R6769 GND.n4218 GND.n3523 280.613
R6770 GND.n4218 GND.n4217 280.613
R6771 GND.n4217 GND.n4216 280.613
R6772 GND.n4216 GND.n3531 280.613
R6773 GND.n4210 GND.n3531 280.613
R6774 GND.n4210 GND.n4209 280.613
R6775 GND.n4209 GND.n4208 280.613
R6776 GND.n4208 GND.n3539 280.613
R6777 GND.n4202 GND.n3539 280.613
R6778 GND.n4202 GND.n4201 280.613
R6779 GND.n4201 GND.n4200 280.613
R6780 GND.n4200 GND.n3547 280.613
R6781 GND.n4194 GND.n3547 280.613
R6782 GND.n4194 GND.n4193 280.613
R6783 GND.n4193 GND.n4192 280.613
R6784 GND.n4192 GND.n3555 280.613
R6785 GND.n4186 GND.n3555 280.613
R6786 GND.n4186 GND.n4185 280.613
R6787 GND.n4185 GND.n4184 280.613
R6788 GND.n4184 GND.n3563 280.613
R6789 GND.n4178 GND.n3563 280.613
R6790 GND.n4178 GND.n4177 280.613
R6791 GND.n4177 GND.n4176 280.613
R6792 GND.n4176 GND.n3571 280.613
R6793 GND.n4170 GND.n3571 280.613
R6794 GND.n4170 GND.n4169 280.613
R6795 GND.n4169 GND.n4168 280.613
R6796 GND.n4168 GND.n3579 280.613
R6797 GND.n4162 GND.n3579 280.613
R6798 GND.n4162 GND.n4161 280.613
R6799 GND.n4161 GND.n4160 280.613
R6800 GND.n4160 GND.n3587 280.613
R6801 GND.n4154 GND.n3587 280.613
R6802 GND.n4154 GND.n4153 280.613
R6803 GND.n4153 GND.n4152 280.613
R6804 GND.n4152 GND.n3595 280.613
R6805 GND.n4146 GND.n3595 280.613
R6806 GND.n4146 GND.n4145 280.613
R6807 GND.n4145 GND.n4144 280.613
R6808 GND.n4144 GND.n3603 280.613
R6809 GND.n4138 GND.n3603 280.613
R6810 GND.n4138 GND.n4137 280.613
R6811 GND.n4137 GND.n4136 280.613
R6812 GND.n4136 GND.n3611 280.613
R6813 GND.n4130 GND.n3611 280.613
R6814 GND.n4130 GND.n4129 280.613
R6815 GND.n4129 GND.n4128 280.613
R6816 GND.n4128 GND.n3619 280.613
R6817 GND.n4122 GND.n3619 280.613
R6818 GND.n4122 GND.n4121 280.613
R6819 GND.n4121 GND.n4120 280.613
R6820 GND.n4120 GND.n3627 280.613
R6821 GND.n4114 GND.n3627 280.613
R6822 GND.n4114 GND.n4113 280.613
R6823 GND.n4113 GND.n4112 280.613
R6824 GND.n4112 GND.n3635 280.613
R6825 GND.n4106 GND.n3635 280.613
R6826 GND.n4106 GND.n4105 280.613
R6827 GND.n4105 GND.n4104 280.613
R6828 GND.n4104 GND.n3643 280.613
R6829 GND.n4098 GND.n3643 280.613
R6830 GND.n4098 GND.n4097 280.613
R6831 GND.n4097 GND.n4096 280.613
R6832 GND.n4096 GND.n3651 280.613
R6833 GND.n4090 GND.n3651 280.613
R6834 GND.n4090 GND.n4089 280.613
R6835 GND.n4089 GND.n4088 280.613
R6836 GND.n4088 GND.n3659 280.613
R6837 GND.n4082 GND.n3659 280.613
R6838 GND.n4082 GND.n4081 280.613
R6839 GND.n4081 GND.n4080 280.613
R6840 GND.n4080 GND.n3667 280.613
R6841 GND.n4074 GND.n3667 280.613
R6842 GND.n4074 GND.n4073 280.613
R6843 GND.n4073 GND.n4072 280.613
R6844 GND.n4072 GND.n3675 280.613
R6845 GND.n4066 GND.n3675 280.613
R6846 GND.n4066 GND.n4065 280.613
R6847 GND.n4065 GND.n4064 280.613
R6848 GND.n4064 GND.n3683 280.613
R6849 GND.n4058 GND.n3683 280.613
R6850 GND.n4058 GND.n4057 280.613
R6851 GND.n4057 GND.n4056 280.613
R6852 GND.n4056 GND.n3691 280.613
R6853 GND.n4050 GND.n3691 280.613
R6854 GND.n4050 GND.n4049 280.613
R6855 GND.n4049 GND.n4048 280.613
R6856 GND.n4048 GND.n3699 280.613
R6857 GND.n4042 GND.n3699 280.613
R6858 GND.n4042 GND.n4041 280.613
R6859 GND.n4041 GND.n4040 280.613
R6860 GND.n4040 GND.n3707 280.613
R6861 GND.n4034 GND.n3707 280.613
R6862 GND.n4034 GND.n4033 280.613
R6863 GND.n4033 GND.n4032 280.613
R6864 GND.n4032 GND.n3715 280.613
R6865 GND.n4026 GND.n3715 280.613
R6866 GND.n4026 GND.n4025 280.613
R6867 GND.n4025 GND.n4024 280.613
R6868 GND.n4024 GND.n3723 280.613
R6869 GND.n4018 GND.n3723 280.613
R6870 GND.n4018 GND.n4017 280.613
R6871 GND.n4017 GND.n4016 280.613
R6872 GND.n4016 GND.n3731 280.613
R6873 GND.n4010 GND.n3731 280.613
R6874 GND.n4010 GND.n4009 280.613
R6875 GND.n4009 GND.n4008 280.613
R6876 GND.n4008 GND.n3739 280.613
R6877 GND.n4002 GND.n3739 280.613
R6878 GND.n4002 GND.n4001 280.613
R6879 GND.n4001 GND.n4000 280.613
R6880 GND.n4000 GND.n3747 280.613
R6881 GND.n3994 GND.n3747 280.613
R6882 GND.n3994 GND.n3993 280.613
R6883 GND.n3993 GND.n3992 280.613
R6884 GND.n3992 GND.n3755 280.613
R6885 GND.n3986 GND.n3755 280.613
R6886 GND.n3986 GND.n3985 280.613
R6887 GND.n3985 GND.n3984 280.613
R6888 GND.n3984 GND.n3763 280.613
R6889 GND.n3978 GND.n3763 280.613
R6890 GND.n3978 GND.n3977 280.613
R6891 GND.n3977 GND.n3976 280.613
R6892 GND.n3976 GND.n3771 280.613
R6893 GND.n3970 GND.n3771 280.613
R6894 GND.n3970 GND.n3969 280.613
R6895 GND.n3969 GND.n3968 280.613
R6896 GND.n3968 GND.n3779 280.613
R6897 GND.n6237 GND.n6236 256.663
R6898 GND.n6237 GND.n1825 256.663
R6899 GND.n6237 GND.n1826 256.663
R6900 GND.n6237 GND.n1827 256.663
R6901 GND.n6237 GND.n1828 256.663
R6902 GND.n6237 GND.n1829 256.663
R6903 GND.n6237 GND.n1830 256.663
R6904 GND.n6237 GND.n1831 256.663
R6905 GND.n6237 GND.n1832 256.663
R6906 GND.n6237 GND.n1833 256.663
R6907 GND.n6238 GND.n6237 256.663
R6908 GND.n6241 GND.n1821 256.663
R6909 GND.n6237 GND.n1834 256.663
R6910 GND.n6237 GND.n1835 256.663
R6911 GND.n6237 GND.n1836 256.663
R6912 GND.n6237 GND.n1837 256.663
R6913 GND.n6237 GND.n1838 256.663
R6914 GND.n6237 GND.n1839 256.663
R6915 GND.n6237 GND.n1840 256.663
R6916 GND.n6237 GND.n1841 256.663
R6917 GND.n6237 GND.n1842 256.663
R6918 GND.n6237 GND.n1843 256.663
R6919 GND.n6237 GND.n1844 256.663
R6920 GND.n7556 GND.n850 256.663
R6921 GND.n7556 GND.n849 256.663
R6922 GND.n7556 GND.n848 256.663
R6923 GND.n7556 GND.n847 256.663
R6924 GND.n7556 GND.n846 256.663
R6925 GND.n7556 GND.n845 256.663
R6926 GND.n7556 GND.n844 256.663
R6927 GND.n7556 GND.n843 256.663
R6928 GND.n7556 GND.n842 256.663
R6929 GND.n7556 GND.n841 256.663
R6930 GND.n7556 GND.n840 256.663
R6931 GND.n7559 GND.n7558 256.663
R6932 GND.n7556 GND.n837 256.663
R6933 GND.n7556 GND.n852 256.663
R6934 GND.n7556 GND.n853 256.663
R6935 GND.n7556 GND.n854 256.663
R6936 GND.n7556 GND.n855 256.663
R6937 GND.n7556 GND.n856 256.663
R6938 GND.n7556 GND.n857 256.663
R6939 GND.n7556 GND.n858 256.663
R6940 GND.n7556 GND.n859 256.663
R6941 GND.n7556 GND.n860 256.663
R6942 GND.n7556 GND.n861 256.663
R6943 GND.n6297 GND.t92 248.602
R6944 GND.n6939 GND.t129 248.602
R6945 GND.n4730 GND.n2976 242.672
R6946 GND.n4732 GND.n2976 242.672
R6947 GND.n4740 GND.n2976 242.672
R6948 GND.n4742 GND.n2976 242.672
R6949 GND.n4750 GND.n2976 242.672
R6950 GND.n4752 GND.n2976 242.672
R6951 GND.n4760 GND.n2976 242.672
R6952 GND.n4762 GND.n2976 242.672
R6953 GND.n4770 GND.n2976 242.672
R6954 GND.n4772 GND.n2976 242.672
R6955 GND.n4780 GND.n2976 242.672
R6956 GND.n4782 GND.n2976 242.672
R6957 GND.n4790 GND.n2976 242.672
R6958 GND.n4792 GND.n2976 242.672
R6959 GND.n4800 GND.n2976 242.672
R6960 GND.n4802 GND.n2976 242.672
R6961 GND.n4810 GND.n2976 242.672
R6962 GND.n4812 GND.n2976 242.672
R6963 GND.n4820 GND.n2976 242.672
R6964 GND.n4822 GND.n2976 242.672
R6965 GND.n4830 GND.n2976 242.672
R6966 GND.n4832 GND.n2976 242.672
R6967 GND.n4841 GND.n2976 242.672
R6968 GND.n4844 GND.n2976 242.672
R6969 GND.n7701 GND.n706 242.672
R6970 GND.n7701 GND.n707 242.672
R6971 GND.n7701 GND.n708 242.672
R6972 GND.n7701 GND.n709 242.672
R6973 GND.n7701 GND.n710 242.672
R6974 GND.n8448 GND.n356 242.672
R6975 GND.n8448 GND.n355 242.672
R6976 GND.n8448 GND.n354 242.672
R6977 GND.n8448 GND.n353 242.672
R6978 GND.n8448 GND.n352 242.672
R6979 GND.n6316 GND.n1592 242.672
R6980 GND.n6324 GND.n1592 242.672
R6981 GND.n6326 GND.n1592 242.672
R6982 GND.n6335 GND.n1592 242.672
R6983 GND.n6337 GND.n1592 242.672
R6984 GND.n6343 GND.n1592 242.672
R6985 GND.n6348 GND.n1592 242.672
R6986 GND.n6353 GND.n1592 242.672
R6987 GND.n6358 GND.n1592 242.672
R6988 GND.n6363 GND.n1592 242.672
R6989 GND.n6365 GND.n1592 242.672
R6990 GND.n6374 GND.n1592 242.672
R6991 GND.n6933 GND.n1161 242.672
R6992 GND.n1285 GND.n1161 242.672
R6993 GND.n6944 GND.n1161 242.672
R6994 GND.n1281 GND.n1161 242.672
R6995 GND.n6952 GND.n1161 242.672
R6996 GND.n1277 GND.n1161 242.672
R6997 GND.n6959 GND.n1161 242.672
R6998 GND.n1197 GND.n1161 242.672
R6999 GND.n6966 GND.n1161 242.672
R7000 GND.n1190 GND.n1161 242.672
R7001 GND.n6973 GND.n1161 242.672
R7002 GND.n6976 GND.n1161 242.672
R7003 GND.n2975 GND.n2974 242.672
R7004 GND.n2975 GND.n2431 242.672
R7005 GND.n2975 GND.n2432 242.672
R7006 GND.n2975 GND.n2433 242.672
R7007 GND.n2975 GND.n2434 242.672
R7008 GND.n2975 GND.n2435 242.672
R7009 GND.n2975 GND.n2436 242.672
R7010 GND.n2975 GND.n2437 242.672
R7011 GND.n2975 GND.n2438 242.672
R7012 GND.n2975 GND.n2439 242.672
R7013 GND.n2975 GND.n2440 242.672
R7014 GND.n2975 GND.n2441 242.672
R7015 GND.n2975 GND.n2442 242.672
R7016 GND.n2975 GND.n2443 242.672
R7017 GND.n2975 GND.n2444 242.672
R7018 GND.n2975 GND.n2445 242.672
R7019 GND.n2975 GND.n2446 242.672
R7020 GND.n2975 GND.n2447 242.672
R7021 GND.n2975 GND.n2448 242.672
R7022 GND.n2975 GND.n2449 242.672
R7023 GND.n2975 GND.n2450 242.672
R7024 GND.n2975 GND.n2451 242.672
R7025 GND.n2975 GND.n2452 242.672
R7026 GND.n2975 GND.n2453 242.672
R7027 GND.n2975 GND.n2454 242.672
R7028 GND.n2975 GND.n2455 242.672
R7029 GND.n2975 GND.n2456 242.672
R7030 GND.n6282 GND.n1662 242.672
R7031 GND.n6282 GND.n1663 242.672
R7032 GND.n6282 GND.n1664 242.672
R7033 GND.n6282 GND.n1665 242.672
R7034 GND.n6282 GND.n1666 242.672
R7035 GND.n6282 GND.n1667 242.672
R7036 GND.n6282 GND.n1668 242.672
R7037 GND.n6282 GND.n1669 242.672
R7038 GND.n6282 GND.n1670 242.672
R7039 GND.n6282 GND.n1671 242.672
R7040 GND.n6282 GND.n1672 242.672
R7041 GND.n6282 GND.n1673 242.672
R7042 GND.n6282 GND.n1674 242.672
R7043 GND.n6282 GND.n1675 242.672
R7044 GND.n6282 GND.n1676 242.672
R7045 GND.n6242 GND.n1819 242.672
R7046 GND.n6282 GND.n1677 242.672
R7047 GND.n6282 GND.n1678 242.672
R7048 GND.n6282 GND.n1679 242.672
R7049 GND.n6282 GND.n1680 242.672
R7050 GND.n6282 GND.n1681 242.672
R7051 GND.n6282 GND.n1682 242.672
R7052 GND.n6282 GND.n1683 242.672
R7053 GND.n6282 GND.n1684 242.672
R7054 GND.n6282 GND.n1685 242.672
R7055 GND.n6282 GND.n1686 242.672
R7056 GND.n6282 GND.n1687 242.672
R7057 GND.n6282 GND.n1688 242.672
R7058 GND.n7701 GND.n7700 242.672
R7059 GND.n7701 GND.n680 242.672
R7060 GND.n7701 GND.n681 242.672
R7061 GND.n7701 GND.n682 242.672
R7062 GND.n7701 GND.n683 242.672
R7063 GND.n7701 GND.n684 242.672
R7064 GND.n7701 GND.n685 242.672
R7065 GND.n7701 GND.n686 242.672
R7066 GND.n7701 GND.n687 242.672
R7067 GND.n7701 GND.n688 242.672
R7068 GND.n7701 GND.n689 242.672
R7069 GND.n7701 GND.n690 242.672
R7070 GND.n7654 GND.n7560 242.672
R7071 GND.n7701 GND.n691 242.672
R7072 GND.n7701 GND.n692 242.672
R7073 GND.n7701 GND.n693 242.672
R7074 GND.n7701 GND.n694 242.672
R7075 GND.n7701 GND.n695 242.672
R7076 GND.n7701 GND.n696 242.672
R7077 GND.n7701 GND.n697 242.672
R7078 GND.n7701 GND.n698 242.672
R7079 GND.n7701 GND.n699 242.672
R7080 GND.n7701 GND.n700 242.672
R7081 GND.n7701 GND.n701 242.672
R7082 GND.n7701 GND.n702 242.672
R7083 GND.n7701 GND.n703 242.672
R7084 GND.n7701 GND.n704 242.672
R7085 GND.n7701 GND.n705 242.672
R7086 GND.n8448 GND.n357 242.672
R7087 GND.n8448 GND.n358 242.672
R7088 GND.n8448 GND.n359 242.672
R7089 GND.n8448 GND.n360 242.672
R7090 GND.n8448 GND.n361 242.672
R7091 GND.n8448 GND.n362 242.672
R7092 GND.n8448 GND.n363 242.672
R7093 GND.n8448 GND.n364 242.672
R7094 GND.n8448 GND.n365 242.672
R7095 GND.n8448 GND.n366 242.672
R7096 GND.n8448 GND.n367 242.672
R7097 GND.n8448 GND.n368 242.672
R7098 GND.n8448 GND.n369 242.672
R7099 GND.n8448 GND.n370 242.672
R7100 GND.n8448 GND.n371 242.672
R7101 GND.n8448 GND.n372 242.672
R7102 GND.n8448 GND.n373 242.672
R7103 GND.n8448 GND.n374 242.672
R7104 GND.n8448 GND.n375 242.672
R7105 GND.n8448 GND.n376 242.672
R7106 GND.n8448 GND.n377 242.672
R7107 GND.n8448 GND.n378 242.672
R7108 GND.n8448 GND.n379 242.672
R7109 GND.n8448 GND.n380 242.672
R7110 GND.n8448 GND.n381 242.672
R7111 GND.n8448 GND.n382 242.672
R7112 GND.n8448 GND.n383 242.672
R7113 GND.n2975 GND.n2457 242.672
R7114 GND.n2975 GND.n2458 242.672
R7115 GND.n2975 GND.n2459 242.672
R7116 GND.n2975 GND.n2460 242.672
R7117 GND.n2975 GND.n2461 242.672
R7118 GND.n6282 GND.n1655 242.672
R7119 GND.n6282 GND.n1651 242.672
R7120 GND.n6282 GND.n1646 242.672
R7121 GND.n6282 GND.n1641 242.672
R7122 GND.n6283 GND.n6282 242.672
R7123 GND.n8447 GND.n385 240.244
R7124 GND.n8440 GND.n8439 240.244
R7125 GND.n8437 GND.n8436 240.244
R7126 GND.n8433 GND.n8432 240.244
R7127 GND.n8429 GND.n8428 240.244
R7128 GND.n8422 GND.n8421 240.244
R7129 GND.n8419 GND.n8418 240.244
R7130 GND.n8415 GND.n8414 240.244
R7131 GND.n8411 GND.n8410 240.244
R7132 GND.n8407 GND.n8406 240.244
R7133 GND.n408 GND.n407 240.244
R7134 GND.n8399 GND.n8398 240.244
R7135 GND.n8395 GND.n8394 240.244
R7136 GND.n8391 GND.n8390 240.244
R7137 GND.n8387 GND.n8386 240.244
R7138 GND.n8383 GND.n8382 240.244
R7139 GND.n8376 GND.n8375 240.244
R7140 GND.n8373 GND.n8372 240.244
R7141 GND.n8369 GND.n8368 240.244
R7142 GND.n8365 GND.n8364 240.244
R7143 GND.n8361 GND.n8360 240.244
R7144 GND.n432 GND.n431 240.244
R7145 GND.n8353 GND.n8352 240.244
R7146 GND.n8349 GND.n8348 240.244
R7147 GND.n8345 GND.n8344 240.244
R7148 GND.n8341 GND.n8340 240.244
R7149 GND.n8337 GND.n8336 240.244
R7150 GND.n7711 GND.n662 240.244
R7151 GND.n7723 GND.n662 240.244
R7152 GND.n7723 GND.n663 240.244
R7153 GND.n663 GND.n652 240.244
R7154 GND.n652 GND.n642 240.244
R7155 GND.n7743 GND.n642 240.244
R7156 GND.n7743 GND.n643 240.244
R7157 GND.n643 GND.n632 240.244
R7158 GND.n632 GND.n622 240.244
R7159 GND.n7763 GND.n622 240.244
R7160 GND.n7763 GND.n623 240.244
R7161 GND.n623 GND.n612 240.244
R7162 GND.n612 GND.n602 240.244
R7163 GND.n7783 GND.n602 240.244
R7164 GND.n7783 GND.n603 240.244
R7165 GND.n603 GND.n592 240.244
R7166 GND.n592 GND.n581 240.244
R7167 GND.n7807 GND.n581 240.244
R7168 GND.n7807 GND.n582 240.244
R7169 GND.n582 GND.n570 240.244
R7170 GND.n7802 GND.n570 240.244
R7171 GND.n7802 GND.n553 240.244
R7172 GND.n7881 GND.n553 240.244
R7173 GND.n7881 GND.n554 240.244
R7174 GND.n554 GND.n544 240.244
R7175 GND.n544 GND.n534 240.244
R7176 GND.n7901 GND.n534 240.244
R7177 GND.n7901 GND.n535 240.244
R7178 GND.n535 GND.n524 240.244
R7179 GND.n524 GND.n514 240.244
R7180 GND.n7921 GND.n514 240.244
R7181 GND.n7921 GND.n515 240.244
R7182 GND.n515 GND.n504 240.244
R7183 GND.n504 GND.n493 240.244
R7184 GND.n7948 GND.n493 240.244
R7185 GND.n7948 GND.n494 240.244
R7186 GND.n494 GND.n483 240.244
R7187 GND.n483 GND.n123 240.244
R7188 GND.n8599 GND.n123 240.244
R7189 GND.n8599 GND.n124 240.244
R7190 GND.n124 GND.n113 240.244
R7191 GND.n113 GND.n93 240.244
R7192 GND.n8629 GND.n93 240.244
R7193 GND.n8629 GND.n94 240.244
R7194 GND.n8625 GND.n94 240.244
R7195 GND.n8625 GND.n100 240.244
R7196 GND.n8227 GND.n100 240.244
R7197 GND.n8227 GND.n70 240.244
R7198 GND.n8230 GND.n70 240.244
R7199 GND.n8230 GND.n138 240.244
R7200 GND.n144 GND.n138 240.244
R7201 GND.n8571 GND.n144 240.244
R7202 GND.n8571 GND.n145 240.244
R7203 GND.n8567 GND.n145 240.244
R7204 GND.n8567 GND.n151 240.244
R7205 GND.n8559 GND.n151 240.244
R7206 GND.n8559 GND.n166 240.244
R7207 GND.n8555 GND.n166 240.244
R7208 GND.n8555 GND.n171 240.244
R7209 GND.n8547 GND.n171 240.244
R7210 GND.n8547 GND.n186 240.244
R7211 GND.n8543 GND.n186 240.244
R7212 GND.n8543 GND.n191 240.244
R7213 GND.n8535 GND.n191 240.244
R7214 GND.n8535 GND.n208 240.244
R7215 GND.n8531 GND.n208 240.244
R7216 GND.n8531 GND.n213 240.244
R7217 GND.n8523 GND.n213 240.244
R7218 GND.n8523 GND.n229 240.244
R7219 GND.n8519 GND.n229 240.244
R7220 GND.n8519 GND.n234 240.244
R7221 GND.n8511 GND.n234 240.244
R7222 GND.n8511 GND.n250 240.244
R7223 GND.n8507 GND.n250 240.244
R7224 GND.n8507 GND.n255 240.244
R7225 GND.n8499 GND.n255 240.244
R7226 GND.n8499 GND.n271 240.244
R7227 GND.n8495 GND.n271 240.244
R7228 GND.n8495 GND.n276 240.244
R7229 GND.n8487 GND.n276 240.244
R7230 GND.n8487 GND.n292 240.244
R7231 GND.n8483 GND.n292 240.244
R7232 GND.n8483 GND.n297 240.244
R7233 GND.n8475 GND.n297 240.244
R7234 GND.n8475 GND.n313 240.244
R7235 GND.n8471 GND.n313 240.244
R7236 GND.n8471 GND.n318 240.244
R7237 GND.n8463 GND.n318 240.244
R7238 GND.n8463 GND.n334 240.244
R7239 GND.n8459 GND.n334 240.244
R7240 GND.n8459 GND.n339 240.244
R7241 GND.n8307 GND.n339 240.244
R7242 GND.n8307 GND.n8070 240.244
R7243 GND.n8070 GND.n448 240.244
R7244 GND.n8327 GND.n448 240.244
R7245 GND.n8329 GND.n8327 240.244
R7246 GND.n713 GND.n712 240.244
R7247 GND.n7694 GND.n712 240.244
R7248 GND.n7692 GND.n7691 240.244
R7249 GND.n7688 GND.n7687 240.244
R7250 GND.n7684 GND.n7683 240.244
R7251 GND.n7680 GND.n7679 240.244
R7252 GND.n7676 GND.n7675 240.244
R7253 GND.n7672 GND.n7671 240.244
R7254 GND.n7668 GND.n7667 240.244
R7255 GND.n7664 GND.n7663 240.244
R7256 GND.n7659 GND.n828 240.244
R7257 GND.n7657 GND.n7656 240.244
R7258 GND.n7652 GND.n7651 240.244
R7259 GND.n7648 GND.n7647 240.244
R7260 GND.n7644 GND.n7643 240.244
R7261 GND.n7640 GND.n7639 240.244
R7262 GND.n7636 GND.n7635 240.244
R7263 GND.n7632 GND.n7631 240.244
R7264 GND.n7628 GND.n7627 240.244
R7265 GND.n7624 GND.n7623 240.244
R7266 GND.n7619 GND.n7580 240.244
R7267 GND.n7617 GND.n7616 240.244
R7268 GND.n7613 GND.n7612 240.244
R7269 GND.n7609 GND.n7608 240.244
R7270 GND.n7605 GND.n7604 240.244
R7271 GND.n7601 GND.n7600 240.244
R7272 GND.n802 GND.n671 240.244
R7273 GND.n802 GND.n659 240.244
R7274 GND.n799 GND.n659 240.244
R7275 GND.n799 GND.n650 240.244
R7276 GND.n796 GND.n650 240.244
R7277 GND.n796 GND.n639 240.244
R7278 GND.n793 GND.n639 240.244
R7279 GND.n793 GND.n630 240.244
R7280 GND.n790 GND.n630 240.244
R7281 GND.n790 GND.n619 240.244
R7282 GND.n787 GND.n619 240.244
R7283 GND.n787 GND.n610 240.244
R7284 GND.n784 GND.n610 240.244
R7285 GND.n784 GND.n599 240.244
R7286 GND.n781 GND.n599 240.244
R7287 GND.n781 GND.n590 240.244
R7288 GND.n778 GND.n590 240.244
R7289 GND.n778 GND.n578 240.244
R7290 GND.n775 GND.n578 240.244
R7291 GND.n775 GND.n568 240.244
R7292 GND.n772 GND.n568 240.244
R7293 GND.n772 GND.n561 240.244
R7294 GND.n561 GND.n550 240.244
R7295 GND.n768 GND.n550 240.244
R7296 GND.n768 GND.n542 240.244
R7297 GND.n765 GND.n542 240.244
R7298 GND.n765 GND.n531 240.244
R7299 GND.n762 GND.n531 240.244
R7300 GND.n762 GND.n522 240.244
R7301 GND.n759 GND.n522 240.244
R7302 GND.n759 GND.n511 240.244
R7303 GND.n756 GND.n511 240.244
R7304 GND.n756 GND.n502 240.244
R7305 GND.n753 GND.n502 240.244
R7306 GND.n753 GND.n490 240.244
R7307 GND.n490 GND.n479 240.244
R7308 GND.n7958 GND.n479 240.244
R7309 GND.n7959 GND.n7958 240.244
R7310 GND.n7959 GND.n120 240.244
R7311 GND.n7962 GND.n120 240.244
R7312 GND.n7962 GND.n111 240.244
R7313 GND.n7967 GND.n111 240.244
R7314 GND.n7967 GND.n89 240.244
R7315 GND.n7971 GND.n89 240.244
R7316 GND.n7971 GND.n101 240.244
R7317 GND.n7976 GND.n101 240.244
R7318 GND.n7977 GND.n7976 240.244
R7319 GND.n7977 GND.n69 240.244
R7320 GND.n7981 GND.n69 240.244
R7321 GND.n7981 GND.n135 240.244
R7322 GND.n7985 GND.n135 240.244
R7323 GND.n7985 GND.n140 240.244
R7324 GND.n7989 GND.n140 240.244
R7325 GND.n7989 GND.n152 240.244
R7326 GND.n7994 GND.n152 240.244
R7327 GND.n7994 GND.n162 240.244
R7328 GND.n7997 GND.n162 240.244
R7329 GND.n7997 GND.n172 240.244
R7330 GND.n8002 GND.n172 240.244
R7331 GND.n8002 GND.n183 240.244
R7332 GND.n8005 GND.n183 240.244
R7333 GND.n8005 GND.n193 240.244
R7334 GND.n8010 GND.n193 240.244
R7335 GND.n8010 GND.n204 240.244
R7336 GND.n8013 GND.n204 240.244
R7337 GND.n8013 GND.n214 240.244
R7338 GND.n8018 GND.n214 240.244
R7339 GND.n8018 GND.n225 240.244
R7340 GND.n8021 GND.n225 240.244
R7341 GND.n8021 GND.n235 240.244
R7342 GND.n8026 GND.n235 240.244
R7343 GND.n8026 GND.n246 240.244
R7344 GND.n8029 GND.n246 240.244
R7345 GND.n8029 GND.n256 240.244
R7346 GND.n8034 GND.n256 240.244
R7347 GND.n8034 GND.n267 240.244
R7348 GND.n8037 GND.n267 240.244
R7349 GND.n8037 GND.n277 240.244
R7350 GND.n8042 GND.n277 240.244
R7351 GND.n8042 GND.n288 240.244
R7352 GND.n8045 GND.n288 240.244
R7353 GND.n8045 GND.n298 240.244
R7354 GND.n8050 GND.n298 240.244
R7355 GND.n8050 GND.n309 240.244
R7356 GND.n8053 GND.n309 240.244
R7357 GND.n8053 GND.n319 240.244
R7358 GND.n8058 GND.n319 240.244
R7359 GND.n8058 GND.n330 240.244
R7360 GND.n8061 GND.n330 240.244
R7361 GND.n8061 GND.n340 240.244
R7362 GND.n8067 GND.n340 240.244
R7363 GND.n8068 GND.n8067 240.244
R7364 GND.n8317 GND.n8068 240.244
R7365 GND.n8317 GND.n453 240.244
R7366 GND.n8325 GND.n453 240.244
R7367 GND.n8325 GND.n384 240.244
R7368 GND.n6281 GND.n1689 240.244
R7369 GND.n1694 GND.n1693 240.244
R7370 GND.n1696 GND.n1695 240.244
R7371 GND.n1700 GND.n1699 240.244
R7372 GND.n1704 GND.n1701 240.244
R7373 GND.n1708 GND.n1707 240.244
R7374 GND.n1710 GND.n1709 240.244
R7375 GND.n1714 GND.n1713 240.244
R7376 GND.n1716 GND.n1715 240.244
R7377 GND.n1720 GND.n1719 240.244
R7378 GND.n1725 GND.n1724 240.244
R7379 GND.n6244 GND.n6243 240.244
R7380 GND.n1729 GND.n1728 240.244
R7381 GND.n1733 GND.n1732 240.244
R7382 GND.n1737 GND.n1734 240.244
R7383 GND.n1741 GND.n1740 240.244
R7384 GND.n1743 GND.n1742 240.244
R7385 GND.n1747 GND.n1746 240.244
R7386 GND.n1749 GND.n1748 240.244
R7387 GND.n1753 GND.n1752 240.244
R7388 GND.n1758 GND.n1757 240.244
R7389 GND.n1762 GND.n1761 240.244
R7390 GND.n1764 GND.n1763 240.244
R7391 GND.n1768 GND.n1767 240.244
R7392 GND.n1770 GND.n1769 240.244
R7393 GND.n1775 GND.n1774 240.244
R7394 GND.n2542 GND.n2541 240.244
R7395 GND.n2543 GND.n2542 240.244
R7396 GND.n2544 GND.n2543 240.244
R7397 GND.n2561 GND.n2544 240.244
R7398 GND.n2561 GND.n2551 240.244
R7399 GND.n2849 GND.n2551 240.244
R7400 GND.n2849 GND.n2426 240.244
R7401 GND.n2426 GND.n2417 240.244
R7402 GND.n4863 GND.n2417 240.244
R7403 GND.n4863 GND.n2418 240.244
R7404 GND.n2418 GND.n2407 240.244
R7405 GND.n2407 GND.n2397 240.244
R7406 GND.n4883 GND.n2397 240.244
R7407 GND.n4883 GND.n2398 240.244
R7408 GND.n2398 GND.n2387 240.244
R7409 GND.n2387 GND.n2377 240.244
R7410 GND.n4903 GND.n2377 240.244
R7411 GND.n4903 GND.n2378 240.244
R7412 GND.n2378 GND.n2367 240.244
R7413 GND.n2367 GND.n2357 240.244
R7414 GND.n4923 GND.n2357 240.244
R7415 GND.n4923 GND.n2358 240.244
R7416 GND.n2358 GND.n2346 240.244
R7417 GND.n2346 GND.n2337 240.244
R7418 GND.n4943 GND.n2337 240.244
R7419 GND.n4943 GND.n2338 240.244
R7420 GND.n2338 GND.n2327 240.244
R7421 GND.n2327 GND.n2317 240.244
R7422 GND.n4963 GND.n2317 240.244
R7423 GND.n4963 GND.n2318 240.244
R7424 GND.n2318 GND.n2307 240.244
R7425 GND.n2307 GND.n2297 240.244
R7426 GND.n4983 GND.n2297 240.244
R7427 GND.n4983 GND.n2298 240.244
R7428 GND.n2298 GND.n2287 240.244
R7429 GND.n2287 GND.n2277 240.244
R7430 GND.n5003 GND.n2277 240.244
R7431 GND.n5003 GND.n2278 240.244
R7432 GND.n2278 GND.n2267 240.244
R7433 GND.n2267 GND.n2257 240.244
R7434 GND.n5029 GND.n2257 240.244
R7435 GND.n5029 GND.n2258 240.244
R7436 GND.n5022 GND.n2258 240.244
R7437 GND.n5022 GND.n2247 240.244
R7438 GND.n2247 GND.n2234 240.244
R7439 GND.n5049 GND.n2234 240.244
R7440 GND.n5049 GND.n2235 240.244
R7441 GND.n2235 GND.n2223 240.244
R7442 GND.n2223 GND.n2211 240.244
R7443 GND.n5074 GND.n2211 240.244
R7444 GND.n5074 GND.n2212 240.244
R7445 GND.n2212 GND.n2201 240.244
R7446 GND.n5065 GND.n2201 240.244
R7447 GND.n5065 GND.n2075 240.244
R7448 GND.n2075 GND.n2065 240.244
R7449 GND.n5106 GND.n2065 240.244
R7450 GND.n5106 GND.n2066 240.244
R7451 GND.n2066 GND.n2054 240.244
R7452 GND.n5099 GND.n2054 240.244
R7453 GND.n5099 GND.n2037 240.244
R7454 GND.n5197 GND.n2037 240.244
R7455 GND.n5197 GND.n2038 240.244
R7456 GND.n2038 GND.n2028 240.244
R7457 GND.n2028 GND.n2018 240.244
R7458 GND.n5217 GND.n2018 240.244
R7459 GND.n5217 GND.n2019 240.244
R7460 GND.n2019 GND.n2008 240.244
R7461 GND.n2008 GND.n1998 240.244
R7462 GND.n5237 GND.n1998 240.244
R7463 GND.n5237 GND.n1999 240.244
R7464 GND.n1999 GND.n1988 240.244
R7465 GND.n1988 GND.n1978 240.244
R7466 GND.n5257 GND.n1978 240.244
R7467 GND.n5257 GND.n1979 240.244
R7468 GND.n1979 GND.n1968 240.244
R7469 GND.n1968 GND.n1958 240.244
R7470 GND.n5277 GND.n1958 240.244
R7471 GND.n5277 GND.n1959 240.244
R7472 GND.n1959 GND.n1948 240.244
R7473 GND.n1948 GND.n1938 240.244
R7474 GND.n5297 GND.n1938 240.244
R7475 GND.n5297 GND.n1939 240.244
R7476 GND.n1939 GND.n1928 240.244
R7477 GND.n1928 GND.n1918 240.244
R7478 GND.n5322 GND.n1918 240.244
R7479 GND.n5322 GND.n1919 240.244
R7480 GND.n1919 GND.n1907 240.244
R7481 GND.n5315 GND.n1907 240.244
R7482 GND.n5315 GND.n1890 240.244
R7483 GND.n5367 GND.n1890 240.244
R7484 GND.n5367 GND.n1891 240.244
R7485 GND.n1891 GND.n1881 240.244
R7486 GND.n1881 GND.n1873 240.244
R7487 GND.n5386 GND.n1873 240.244
R7488 GND.n5386 GND.n1628 240.244
R7489 GND.n6287 GND.n1628 240.244
R7490 GND.n2465 GND.n2464 240.244
R7491 GND.n2968 GND.n2464 240.244
R7492 GND.n2966 GND.n2965 240.244
R7493 GND.n2962 GND.n2961 240.244
R7494 GND.n2958 GND.n2957 240.244
R7495 GND.n2954 GND.n2953 240.244
R7496 GND.n2950 GND.n2949 240.244
R7497 GND.n2946 GND.n2945 240.244
R7498 GND.n2942 GND.n2941 240.244
R7499 GND.n2938 GND.n2937 240.244
R7500 GND.n2933 GND.n2489 240.244
R7501 GND.n2931 GND.n2930 240.244
R7502 GND.n2927 GND.n2926 240.244
R7503 GND.n2923 GND.n2922 240.244
R7504 GND.n2919 GND.n2918 240.244
R7505 GND.n2915 GND.n2914 240.244
R7506 GND.n2911 GND.n2910 240.244
R7507 GND.n2907 GND.n2906 240.244
R7508 GND.n2903 GND.n2902 240.244
R7509 GND.n2899 GND.n2898 240.244
R7510 GND.n2895 GND.n2894 240.244
R7511 GND.n2890 GND.n2516 240.244
R7512 GND.n2888 GND.n2887 240.244
R7513 GND.n2884 GND.n2883 240.244
R7514 GND.n2880 GND.n2879 240.244
R7515 GND.n2876 GND.n2875 240.244
R7516 GND.n2872 GND.n2871 240.244
R7517 GND.n2571 GND.n2466 240.244
R7518 GND.n2614 GND.n2571 240.244
R7519 GND.n2614 GND.n2564 240.244
R7520 GND.n2715 GND.n2564 240.244
R7521 GND.n2715 GND.n2565 240.244
R7522 GND.n2565 GND.n2553 240.244
R7523 GND.n2553 GND.n2424 240.244
R7524 GND.n2709 GND.n2424 240.244
R7525 GND.n2709 GND.n2414 240.244
R7526 GND.n2706 GND.n2414 240.244
R7527 GND.n2706 GND.n2405 240.244
R7528 GND.n2703 GND.n2405 240.244
R7529 GND.n2703 GND.n2394 240.244
R7530 GND.n2700 GND.n2394 240.244
R7531 GND.n2700 GND.n2385 240.244
R7532 GND.n2697 GND.n2385 240.244
R7533 GND.n2697 GND.n2374 240.244
R7534 GND.n2694 GND.n2374 240.244
R7535 GND.n2694 GND.n2365 240.244
R7536 GND.n2691 GND.n2365 240.244
R7537 GND.n2691 GND.n2353 240.244
R7538 GND.n2688 GND.n2353 240.244
R7539 GND.n2688 GND.n2344 240.244
R7540 GND.n2685 GND.n2344 240.244
R7541 GND.n2685 GND.n2334 240.244
R7542 GND.n2682 GND.n2334 240.244
R7543 GND.n2682 GND.n2325 240.244
R7544 GND.n2679 GND.n2325 240.244
R7545 GND.n2679 GND.n2314 240.244
R7546 GND.n2676 GND.n2314 240.244
R7547 GND.n2676 GND.n2305 240.244
R7548 GND.n2673 GND.n2305 240.244
R7549 GND.n2673 GND.n2294 240.244
R7550 GND.n2670 GND.n2294 240.244
R7551 GND.n2670 GND.n2285 240.244
R7552 GND.n2667 GND.n2285 240.244
R7553 GND.n2667 GND.n2274 240.244
R7554 GND.n2664 GND.n2274 240.244
R7555 GND.n2664 GND.n2265 240.244
R7556 GND.n2661 GND.n2265 240.244
R7557 GND.n2661 GND.n2253 240.244
R7558 GND.n2658 GND.n2253 240.244
R7559 GND.n2658 GND.n2657 240.244
R7560 GND.n2657 GND.n2245 240.244
R7561 GND.n2245 GND.n2242 240.244
R7562 GND.n2242 GND.n2231 240.244
R7563 GND.n2231 GND.n2228 240.244
R7564 GND.n2228 GND.n2222 240.244
R7565 GND.n2222 GND.n2219 240.244
R7566 GND.n2219 GND.n2208 240.244
R7567 GND.n2208 GND.n2197 240.244
R7568 GND.n5082 GND.n2197 240.244
R7569 GND.n5083 GND.n5082 240.244
R7570 GND.n5083 GND.n2073 240.244
R7571 GND.n2194 GND.n2073 240.244
R7572 GND.n2194 GND.n2062 240.244
R7573 GND.n2191 GND.n2062 240.244
R7574 GND.n2191 GND.n2052 240.244
R7575 GND.n2188 GND.n2052 240.244
R7576 GND.n2188 GND.n2045 240.244
R7577 GND.n2045 GND.n2034 240.244
R7578 GND.n2184 GND.n2034 240.244
R7579 GND.n2184 GND.n2026 240.244
R7580 GND.n2181 GND.n2026 240.244
R7581 GND.n2181 GND.n2015 240.244
R7582 GND.n2178 GND.n2015 240.244
R7583 GND.n2178 GND.n2006 240.244
R7584 GND.n2175 GND.n2006 240.244
R7585 GND.n2175 GND.n1995 240.244
R7586 GND.n2172 GND.n1995 240.244
R7587 GND.n2172 GND.n1986 240.244
R7588 GND.n2169 GND.n1986 240.244
R7589 GND.n2169 GND.n1975 240.244
R7590 GND.n2166 GND.n1975 240.244
R7591 GND.n2166 GND.n1966 240.244
R7592 GND.n2163 GND.n1966 240.244
R7593 GND.n2163 GND.n1955 240.244
R7594 GND.n2160 GND.n1955 240.244
R7595 GND.n2160 GND.n1946 240.244
R7596 GND.n2157 GND.n1946 240.244
R7597 GND.n2157 GND.n1935 240.244
R7598 GND.n2154 GND.n1935 240.244
R7599 GND.n2154 GND.n1926 240.244
R7600 GND.n2151 GND.n1926 240.244
R7601 GND.n2151 GND.n1915 240.244
R7602 GND.n2148 GND.n1915 240.244
R7603 GND.n2148 GND.n1905 240.244
R7604 GND.n2145 GND.n1905 240.244
R7605 GND.n2145 GND.n1898 240.244
R7606 GND.n1898 GND.n1887 240.244
R7607 GND.n2141 GND.n1887 240.244
R7608 GND.n2141 GND.n1879 240.244
R7609 GND.n2138 GND.n1879 240.244
R7610 GND.n2138 GND.n1870 240.244
R7611 GND.n2135 GND.n1870 240.244
R7612 GND.n2135 GND.n1632 240.244
R7613 GND.n6977 GND.n1177 240.244
R7614 GND.n6975 GND.n6974 240.244
R7615 GND.n6972 GND.n1183 240.244
R7616 GND.n6968 GND.n6967 240.244
R7617 GND.n6965 GND.n1191 240.244
R7618 GND.n6961 GND.n6960 240.244
R7619 GND.n6958 GND.n1198 240.244
R7620 GND.n6954 GND.n6953 240.244
R7621 GND.n6951 GND.n1279 240.244
R7622 GND.n6946 GND.n6945 240.244
R7623 GND.n6943 GND.n1283 240.244
R7624 GND.n6935 GND.n6934 240.244
R7625 GND.n6377 GND.n6376 240.244
R7626 GND.n6377 GND.n1572 240.244
R7627 GND.n6406 GND.n1572 240.244
R7628 GND.n6406 GND.n1565 240.244
R7629 GND.n1565 GND.n1556 240.244
R7630 GND.n1556 GND.n1545 240.244
R7631 GND.n6400 GND.n1545 240.244
R7632 GND.n6400 GND.n1536 240.244
R7633 GND.n6397 GND.n1536 240.244
R7634 GND.n6397 GND.n6396 240.244
R7635 GND.n6396 GND.n6395 240.244
R7636 GND.n6395 GND.n1509 240.244
R7637 GND.n1509 GND.n1501 240.244
R7638 GND.n6554 GND.n1501 240.244
R7639 GND.n6554 GND.n1492 240.244
R7640 GND.n1492 GND.n1483 240.244
R7641 GND.n6572 GND.n1483 240.244
R7642 GND.n6572 GND.n1475 240.244
R7643 GND.n6568 GND.n1475 240.244
R7644 GND.n6568 GND.n1442 240.244
R7645 GND.n1442 GND.n1432 240.244
R7646 GND.n6646 GND.n1432 240.244
R7647 GND.n6647 GND.n6646 240.244
R7648 GND.n6648 GND.n6647 240.244
R7649 GND.n6648 GND.n1412 240.244
R7650 GND.n1428 GND.n1412 240.244
R7651 GND.n1428 GND.n1404 240.244
R7652 GND.n6655 GND.n1404 240.244
R7653 GND.n6655 GND.n1389 240.244
R7654 GND.n1389 GND.n1381 240.244
R7655 GND.n6664 GND.n1381 240.244
R7656 GND.n6664 GND.n1372 240.244
R7657 GND.n1372 GND.n1359 240.244
R7658 GND.n6791 GND.n1359 240.244
R7659 GND.n6791 GND.n1350 240.244
R7660 GND.n6820 GND.n1350 240.244
R7661 GND.n6820 GND.n1343 240.244
R7662 GND.n1343 GND.n1339 240.244
R7663 GND.n1339 GND.n1330 240.244
R7664 GND.n6814 GND.n1330 240.244
R7665 GND.n6814 GND.n6813 240.244
R7666 GND.n6813 GND.n6812 240.244
R7667 GND.n6812 GND.n1321 240.244
R7668 GND.n6808 GND.n1321 240.244
R7669 GND.n6808 GND.n1289 240.244
R7670 GND.n6926 GND.n1289 240.244
R7671 GND.n6926 GND.n1174 240.244
R7672 GND.n6317 GND.n6308 240.244
R7673 GND.n6323 GND.n6308 240.244
R7674 GND.n6327 GND.n6325 240.244
R7675 GND.n6334 GND.n6304 240.244
R7676 GND.n6338 GND.n6336 240.244
R7677 GND.n6342 GND.n6301 240.244
R7678 GND.n6347 GND.n6344 240.244
R7679 GND.n6352 GND.n6349 240.244
R7680 GND.n6357 GND.n6354 240.244
R7681 GND.n6362 GND.n6359 240.244
R7682 GND.n6366 GND.n6364 240.244
R7683 GND.n6373 GND.n1614 240.244
R7684 GND.n6314 GND.n1570 240.244
R7685 GND.n6450 GND.n1570 240.244
R7686 GND.n6450 GND.n1566 240.244
R7687 GND.n6456 GND.n1566 240.244
R7688 GND.n6456 GND.n1543 240.244
R7689 GND.n6483 GND.n1543 240.244
R7690 GND.n6483 GND.n1538 240.244
R7691 GND.n6494 GND.n1538 240.244
R7692 GND.n6494 GND.n1539 240.244
R7693 GND.n6490 GND.n1539 240.244
R7694 GND.n6490 GND.n1507 240.244
R7695 GND.n6546 GND.n1507 240.244
R7696 GND.n6546 GND.n1503 240.244
R7697 GND.n6552 GND.n1503 240.244
R7698 GND.n6552 GND.n1481 240.244
R7699 GND.n6598 GND.n1481 240.244
R7700 GND.n6598 GND.n1477 240.244
R7701 GND.n6604 GND.n1477 240.244
R7702 GND.n6604 GND.n1441 240.244
R7703 GND.n6636 GND.n1441 240.244
R7704 GND.n6636 GND.n1436 240.244
R7705 GND.n6644 GND.n1436 240.244
R7706 GND.n6644 GND.n1437 240.244
R7707 GND.n1437 GND.n1410 240.244
R7708 GND.n6695 GND.n1410 240.244
R7709 GND.n6695 GND.n1405 240.244
R7710 GND.n6703 GND.n1405 240.244
R7711 GND.n6703 GND.n1406 240.244
R7712 GND.n1406 GND.n1379 240.244
R7713 GND.n6763 GND.n1379 240.244
R7714 GND.n6763 GND.n1374 240.244
R7715 GND.n6771 GND.n1374 240.244
R7716 GND.n6771 GND.n1375 240.244
R7717 GND.n1375 GND.n1348 240.244
R7718 GND.n6830 GND.n1348 240.244
R7719 GND.n6830 GND.n1344 240.244
R7720 GND.n6839 GND.n1344 240.244
R7721 GND.n6839 GND.n1327 240.244
R7722 GND.n6858 GND.n1327 240.244
R7723 GND.n6859 GND.n6858 240.244
R7724 GND.n6860 GND.n6859 240.244
R7725 GND.n6860 GND.n1322 240.244
R7726 GND.n6871 GND.n1322 240.244
R7727 GND.n6871 GND.n1323 240.244
R7728 GND.n6867 GND.n1323 240.244
R7729 GND.n6867 GND.n1176 240.244
R7730 GND.n6983 GND.n1176 240.244
R7731 GND.n8191 GND.n351 240.244
R7732 GND.n8197 GND.n8196 240.244
R7733 GND.n8200 GND.n8199 240.244
R7734 GND.n8207 GND.n8206 240.244
R7735 GND.n8210 GND.n8209 240.244
R7736 GND.n1228 GND.n673 240.244
R7737 GND.n1228 GND.n661 240.244
R7738 GND.n1268 GND.n661 240.244
R7739 GND.n1268 GND.n651 240.244
R7740 GND.n1265 GND.n651 240.244
R7741 GND.n1265 GND.n641 240.244
R7742 GND.n1262 GND.n641 240.244
R7743 GND.n1262 GND.n631 240.244
R7744 GND.n1259 GND.n631 240.244
R7745 GND.n1259 GND.n621 240.244
R7746 GND.n1256 GND.n621 240.244
R7747 GND.n1256 GND.n611 240.244
R7748 GND.n1253 GND.n611 240.244
R7749 GND.n1253 GND.n601 240.244
R7750 GND.n1250 GND.n601 240.244
R7751 GND.n1250 GND.n591 240.244
R7752 GND.n1247 GND.n591 240.244
R7753 GND.n1247 GND.n580 240.244
R7754 GND.n580 GND.n566 240.244
R7755 GND.n7819 GND.n566 240.244
R7756 GND.n7819 GND.n562 240.244
R7757 GND.n7870 GND.n562 240.244
R7758 GND.n7870 GND.n552 240.244
R7759 GND.n7866 GND.n552 240.244
R7760 GND.n7866 GND.n543 240.244
R7761 GND.n7863 GND.n543 240.244
R7762 GND.n7863 GND.n533 240.244
R7763 GND.n7860 GND.n533 240.244
R7764 GND.n7860 GND.n523 240.244
R7765 GND.n7857 GND.n523 240.244
R7766 GND.n7857 GND.n513 240.244
R7767 GND.n7854 GND.n513 240.244
R7768 GND.n7854 GND.n503 240.244
R7769 GND.n7851 GND.n503 240.244
R7770 GND.n7851 GND.n492 240.244
R7771 GND.n7848 GND.n492 240.244
R7772 GND.n7848 GND.n482 240.244
R7773 GND.n7845 GND.n482 240.244
R7774 GND.n7845 GND.n122 240.244
R7775 GND.n122 GND.n109 240.244
R7776 GND.n8609 GND.n109 240.244
R7777 GND.n8610 GND.n8609 240.244
R7778 GND.n8610 GND.n92 240.244
R7779 GND.n104 GND.n92 240.244
R7780 GND.n8619 GND.n104 240.244
R7781 GND.n8619 GND.n105 240.244
R7782 GND.n105 GND.n66 240.244
R7783 GND.n8637 GND.n66 240.244
R7784 GND.n8637 GND.n67 240.244
R7785 GND.n137 GND.n67 240.244
R7786 GND.n8096 GND.n137 240.244
R7787 GND.n8096 GND.n143 240.244
R7788 GND.n8101 GND.n143 240.244
R7789 GND.n8101 GND.n155 240.244
R7790 GND.n8104 GND.n155 240.244
R7791 GND.n8104 GND.n165 240.244
R7792 GND.n8109 GND.n165 240.244
R7793 GND.n8109 GND.n175 240.244
R7794 GND.n8112 GND.n175 240.244
R7795 GND.n8112 GND.n185 240.244
R7796 GND.n8117 GND.n185 240.244
R7797 GND.n8117 GND.n196 240.244
R7798 GND.n8120 GND.n196 240.244
R7799 GND.n8120 GND.n207 240.244
R7800 GND.n8125 GND.n207 240.244
R7801 GND.n8125 GND.n217 240.244
R7802 GND.n8128 GND.n217 240.244
R7803 GND.n8128 GND.n228 240.244
R7804 GND.n8133 GND.n228 240.244
R7805 GND.n8133 GND.n238 240.244
R7806 GND.n8136 GND.n238 240.244
R7807 GND.n8136 GND.n249 240.244
R7808 GND.n8141 GND.n249 240.244
R7809 GND.n8141 GND.n259 240.244
R7810 GND.n8144 GND.n259 240.244
R7811 GND.n8144 GND.n270 240.244
R7812 GND.n8149 GND.n270 240.244
R7813 GND.n8149 GND.n280 240.244
R7814 GND.n8152 GND.n280 240.244
R7815 GND.n8152 GND.n291 240.244
R7816 GND.n8157 GND.n291 240.244
R7817 GND.n8157 GND.n301 240.244
R7818 GND.n8160 GND.n301 240.244
R7819 GND.n8160 GND.n312 240.244
R7820 GND.n8165 GND.n312 240.244
R7821 GND.n8165 GND.n322 240.244
R7822 GND.n8168 GND.n322 240.244
R7823 GND.n8168 GND.n333 240.244
R7824 GND.n8173 GND.n333 240.244
R7825 GND.n8173 GND.n343 240.244
R7826 GND.n8176 GND.n343 240.244
R7827 GND.n8176 GND.n8071 240.244
R7828 GND.n8222 GND.n8071 240.244
R7829 GND.n8222 GND.n8072 240.244
R7830 GND.n8072 GND.n450 240.244
R7831 GND.n8217 GND.n450 240.244
R7832 GND.n1223 GND.n1222 240.244
R7833 GND.n1219 GND.n1218 240.244
R7834 GND.n1215 GND.n1214 240.244
R7835 GND.n1211 GND.n1210 240.244
R7836 GND.n1205 GND.n711 240.244
R7837 GND.n672 GND.n667 240.244
R7838 GND.n667 GND.n660 240.244
R7839 GND.n660 GND.n648 240.244
R7840 GND.n7733 GND.n648 240.244
R7841 GND.n7734 GND.n7733 240.244
R7842 GND.n7734 GND.n640 240.244
R7843 GND.n640 GND.n628 240.244
R7844 GND.n7753 GND.n628 240.244
R7845 GND.n7754 GND.n7753 240.244
R7846 GND.n7754 GND.n620 240.244
R7847 GND.n620 GND.n608 240.244
R7848 GND.n7773 GND.n608 240.244
R7849 GND.n7774 GND.n7773 240.244
R7850 GND.n7774 GND.n600 240.244
R7851 GND.n600 GND.n588 240.244
R7852 GND.n7793 GND.n588 240.244
R7853 GND.n7794 GND.n7793 240.244
R7854 GND.n7794 GND.n579 240.244
R7855 GND.n7797 GND.n579 240.244
R7856 GND.n7797 GND.n569 240.244
R7857 GND.n569 GND.n559 240.244
R7858 GND.n7872 GND.n559 240.244
R7859 GND.n7872 GND.n551 240.244
R7860 GND.n551 GND.n540 240.244
R7861 GND.n7891 GND.n540 240.244
R7862 GND.n7892 GND.n7891 240.244
R7863 GND.n7892 GND.n532 240.244
R7864 GND.n532 GND.n520 240.244
R7865 GND.n7911 GND.n520 240.244
R7866 GND.n7912 GND.n7911 240.244
R7867 GND.n7912 GND.n512 240.244
R7868 GND.n512 GND.n500 240.244
R7869 GND.n7931 GND.n500 240.244
R7870 GND.n7932 GND.n7931 240.244
R7871 GND.n7932 GND.n491 240.244
R7872 GND.n7935 GND.n491 240.244
R7873 GND.n7935 GND.n481 240.244
R7874 GND.n7941 GND.n481 240.244
R7875 GND.n7941 GND.n121 240.244
R7876 GND.n7938 GND.n121 240.244
R7877 GND.n7938 GND.n112 240.244
R7878 GND.n8592 GND.n112 240.244
R7879 GND.n8592 GND.n90 240.244
R7880 GND.n8589 GND.n90 240.244
R7881 GND.n8589 GND.n102 240.244
R7882 GND.n8586 GND.n102 240.244
R7883 GND.n8586 GND.n8585 240.244
R7884 GND.n8585 GND.n72 240.244
R7885 GND.n8581 GND.n72 240.244
R7886 GND.n8581 GND.n8580 240.244
R7887 GND.n8580 GND.n134 240.244
R7888 GND.n141 GND.n134 240.244
R7889 GND.n8237 GND.n141 240.244
R7890 GND.n8237 GND.n153 240.244
R7891 GND.n8241 GND.n153 240.244
R7892 GND.n8241 GND.n163 240.244
R7893 GND.n8244 GND.n163 240.244
R7894 GND.n8244 GND.n173 240.244
R7895 GND.n8248 GND.n173 240.244
R7896 GND.n8248 GND.n184 240.244
R7897 GND.n8251 GND.n184 240.244
R7898 GND.n8251 GND.n194 240.244
R7899 GND.n8255 GND.n194 240.244
R7900 GND.n8255 GND.n205 240.244
R7901 GND.n8258 GND.n205 240.244
R7902 GND.n8258 GND.n215 240.244
R7903 GND.n8262 GND.n215 240.244
R7904 GND.n8262 GND.n226 240.244
R7905 GND.n8265 GND.n226 240.244
R7906 GND.n8265 GND.n236 240.244
R7907 GND.n8269 GND.n236 240.244
R7908 GND.n8269 GND.n247 240.244
R7909 GND.n8272 GND.n247 240.244
R7910 GND.n8272 GND.n257 240.244
R7911 GND.n8276 GND.n257 240.244
R7912 GND.n8276 GND.n268 240.244
R7913 GND.n8279 GND.n268 240.244
R7914 GND.n8279 GND.n278 240.244
R7915 GND.n8283 GND.n278 240.244
R7916 GND.n8283 GND.n289 240.244
R7917 GND.n8286 GND.n289 240.244
R7918 GND.n8286 GND.n299 240.244
R7919 GND.n8290 GND.n299 240.244
R7920 GND.n8290 GND.n310 240.244
R7921 GND.n8293 GND.n310 240.244
R7922 GND.n8293 GND.n320 240.244
R7923 GND.n8297 GND.n320 240.244
R7924 GND.n8297 GND.n331 240.244
R7925 GND.n8300 GND.n331 240.244
R7926 GND.n8300 GND.n341 240.244
R7927 GND.n8303 GND.n341 240.244
R7928 GND.n8303 GND.n8223 240.244
R7929 GND.n8315 GND.n8223 240.244
R7930 GND.n8315 GND.n8224 240.244
R7931 GND.n8224 GND.n452 240.244
R7932 GND.n452 GND.n451 240.244
R7933 GND.n4723 GND.n3022 240.244
R7934 GND.n4723 GND.n3025 240.244
R7935 GND.n4719 GND.n3025 240.244
R7936 GND.n4719 GND.n3028 240.244
R7937 GND.n4715 GND.n3028 240.244
R7938 GND.n4715 GND.n3034 240.244
R7939 GND.n4711 GND.n3034 240.244
R7940 GND.n4711 GND.n3036 240.244
R7941 GND.n4707 GND.n3036 240.244
R7942 GND.n4707 GND.n3042 240.244
R7943 GND.n4703 GND.n3042 240.244
R7944 GND.n4703 GND.n3044 240.244
R7945 GND.n4699 GND.n3044 240.244
R7946 GND.n4699 GND.n3050 240.244
R7947 GND.n4695 GND.n3050 240.244
R7948 GND.n4695 GND.n3052 240.244
R7949 GND.n4691 GND.n3052 240.244
R7950 GND.n4691 GND.n3058 240.244
R7951 GND.n4687 GND.n3058 240.244
R7952 GND.n4687 GND.n3060 240.244
R7953 GND.n4683 GND.n3060 240.244
R7954 GND.n4683 GND.n3066 240.244
R7955 GND.n4679 GND.n3066 240.244
R7956 GND.n4679 GND.n3068 240.244
R7957 GND.n4675 GND.n3068 240.244
R7958 GND.n4675 GND.n3074 240.244
R7959 GND.n4671 GND.n3074 240.244
R7960 GND.n4671 GND.n3076 240.244
R7961 GND.n4667 GND.n3076 240.244
R7962 GND.n4667 GND.n3082 240.244
R7963 GND.n4663 GND.n3082 240.244
R7964 GND.n4663 GND.n3084 240.244
R7965 GND.n4659 GND.n3084 240.244
R7966 GND.n4659 GND.n3090 240.244
R7967 GND.n4655 GND.n3090 240.244
R7968 GND.n4655 GND.n3092 240.244
R7969 GND.n4651 GND.n3092 240.244
R7970 GND.n4651 GND.n3098 240.244
R7971 GND.n4647 GND.n3098 240.244
R7972 GND.n4647 GND.n3100 240.244
R7973 GND.n4643 GND.n3100 240.244
R7974 GND.n4643 GND.n3106 240.244
R7975 GND.n4639 GND.n3106 240.244
R7976 GND.n4639 GND.n3108 240.244
R7977 GND.n4635 GND.n3108 240.244
R7978 GND.n4635 GND.n3114 240.244
R7979 GND.n4631 GND.n3114 240.244
R7980 GND.n4631 GND.n3116 240.244
R7981 GND.n4627 GND.n3116 240.244
R7982 GND.n4627 GND.n3122 240.244
R7983 GND.n4623 GND.n3122 240.244
R7984 GND.n4623 GND.n3124 240.244
R7985 GND.n4619 GND.n3124 240.244
R7986 GND.n4619 GND.n3130 240.244
R7987 GND.n4615 GND.n3130 240.244
R7988 GND.n4615 GND.n3132 240.244
R7989 GND.n4611 GND.n3132 240.244
R7990 GND.n4611 GND.n3138 240.244
R7991 GND.n4607 GND.n3138 240.244
R7992 GND.n4607 GND.n3140 240.244
R7993 GND.n4603 GND.n3140 240.244
R7994 GND.n4603 GND.n3146 240.244
R7995 GND.n4599 GND.n3146 240.244
R7996 GND.n4599 GND.n3148 240.244
R7997 GND.n4595 GND.n3148 240.244
R7998 GND.n4595 GND.n3154 240.244
R7999 GND.n4591 GND.n3154 240.244
R8000 GND.n4591 GND.n3156 240.244
R8001 GND.n4587 GND.n3156 240.244
R8002 GND.n4587 GND.n3162 240.244
R8003 GND.n4583 GND.n3162 240.244
R8004 GND.n4583 GND.n3164 240.244
R8005 GND.n4579 GND.n3164 240.244
R8006 GND.n4579 GND.n3170 240.244
R8007 GND.n4575 GND.n3170 240.244
R8008 GND.n4575 GND.n3172 240.244
R8009 GND.n4571 GND.n3172 240.244
R8010 GND.n4571 GND.n3178 240.244
R8011 GND.n4567 GND.n3178 240.244
R8012 GND.n4567 GND.n3180 240.244
R8013 GND.n4563 GND.n3180 240.244
R8014 GND.n4563 GND.n3186 240.244
R8015 GND.n4559 GND.n3186 240.244
R8016 GND.n4559 GND.n3188 240.244
R8017 GND.n4555 GND.n3188 240.244
R8018 GND.n4555 GND.n3194 240.244
R8019 GND.n4551 GND.n3194 240.244
R8020 GND.n4551 GND.n3196 240.244
R8021 GND.n4547 GND.n3196 240.244
R8022 GND.n4547 GND.n3202 240.244
R8023 GND.n4543 GND.n3202 240.244
R8024 GND.n4543 GND.n3204 240.244
R8025 GND.n4539 GND.n3204 240.244
R8026 GND.n4539 GND.n3210 240.244
R8027 GND.n4535 GND.n3210 240.244
R8028 GND.n4535 GND.n3212 240.244
R8029 GND.n4531 GND.n3212 240.244
R8030 GND.n4531 GND.n3218 240.244
R8031 GND.n4527 GND.n3218 240.244
R8032 GND.n4527 GND.n3220 240.244
R8033 GND.n4523 GND.n3220 240.244
R8034 GND.n4523 GND.n3226 240.244
R8035 GND.n4519 GND.n3226 240.244
R8036 GND.n4519 GND.n3228 240.244
R8037 GND.n4515 GND.n3228 240.244
R8038 GND.n4515 GND.n3234 240.244
R8039 GND.n4511 GND.n3234 240.244
R8040 GND.n4511 GND.n3236 240.244
R8041 GND.n4507 GND.n3236 240.244
R8042 GND.n4507 GND.n3242 240.244
R8043 GND.n4503 GND.n3242 240.244
R8044 GND.n4503 GND.n3244 240.244
R8045 GND.n4499 GND.n3244 240.244
R8046 GND.n4499 GND.n3250 240.244
R8047 GND.n4495 GND.n3250 240.244
R8048 GND.n4495 GND.n3252 240.244
R8049 GND.n4491 GND.n3252 240.244
R8050 GND.n4491 GND.n3258 240.244
R8051 GND.n4487 GND.n3258 240.244
R8052 GND.n4487 GND.n3260 240.244
R8053 GND.n4483 GND.n3260 240.244
R8054 GND.n4483 GND.n3266 240.244
R8055 GND.n4479 GND.n3266 240.244
R8056 GND.n4479 GND.n3268 240.244
R8057 GND.n4475 GND.n3268 240.244
R8058 GND.n4475 GND.n3274 240.244
R8059 GND.n4471 GND.n3274 240.244
R8060 GND.n4471 GND.n3276 240.244
R8061 GND.n4467 GND.n3276 240.244
R8062 GND.n4467 GND.n3282 240.244
R8063 GND.n4463 GND.n3282 240.244
R8064 GND.n4463 GND.n3284 240.244
R8065 GND.n4459 GND.n3284 240.244
R8066 GND.n4459 GND.n3290 240.244
R8067 GND.n4455 GND.n3290 240.244
R8068 GND.n4455 GND.n3292 240.244
R8069 GND.n4451 GND.n3292 240.244
R8070 GND.n4451 GND.n3298 240.244
R8071 GND.n4447 GND.n3298 240.244
R8072 GND.n4447 GND.n3300 240.244
R8073 GND.n4443 GND.n3300 240.244
R8074 GND.n4443 GND.n3306 240.244
R8075 GND.n4439 GND.n3306 240.244
R8076 GND.n4439 GND.n3308 240.244
R8077 GND.n4435 GND.n3308 240.244
R8078 GND.n4435 GND.n3314 240.244
R8079 GND.n4431 GND.n3314 240.244
R8080 GND.n4431 GND.n3316 240.244
R8081 GND.n4427 GND.n3316 240.244
R8082 GND.n4427 GND.n3322 240.244
R8083 GND.n4423 GND.n3322 240.244
R8084 GND.n4423 GND.n3324 240.244
R8085 GND.n4419 GND.n3324 240.244
R8086 GND.n4419 GND.n3330 240.244
R8087 GND.n4415 GND.n3330 240.244
R8088 GND.n4415 GND.n3332 240.244
R8089 GND.n4411 GND.n3332 240.244
R8090 GND.n4411 GND.n3338 240.244
R8091 GND.n4407 GND.n3338 240.244
R8092 GND.n4407 GND.n3340 240.244
R8093 GND.n4403 GND.n3340 240.244
R8094 GND.n4403 GND.n3346 240.244
R8095 GND.n4399 GND.n3346 240.244
R8096 GND.n4399 GND.n3348 240.244
R8097 GND.n4395 GND.n3348 240.244
R8098 GND.n4395 GND.n3354 240.244
R8099 GND.n4391 GND.n3354 240.244
R8100 GND.n4391 GND.n3356 240.244
R8101 GND.n4387 GND.n3356 240.244
R8102 GND.n4387 GND.n3362 240.244
R8103 GND.n4383 GND.n3362 240.244
R8104 GND.n4383 GND.n3364 240.244
R8105 GND.n4379 GND.n3364 240.244
R8106 GND.n4379 GND.n3370 240.244
R8107 GND.n4375 GND.n3370 240.244
R8108 GND.n4375 GND.n3372 240.244
R8109 GND.n4371 GND.n3372 240.244
R8110 GND.n4371 GND.n3378 240.244
R8111 GND.n4367 GND.n3378 240.244
R8112 GND.n4367 GND.n3380 240.244
R8113 GND.n4363 GND.n3380 240.244
R8114 GND.n4363 GND.n3386 240.244
R8115 GND.n4359 GND.n3386 240.244
R8116 GND.n4359 GND.n3388 240.244
R8117 GND.n4355 GND.n3388 240.244
R8118 GND.n4355 GND.n3394 240.244
R8119 GND.n4351 GND.n3394 240.244
R8120 GND.n4351 GND.n3396 240.244
R8121 GND.n4347 GND.n3396 240.244
R8122 GND.n4347 GND.n3402 240.244
R8123 GND.n4343 GND.n3402 240.244
R8124 GND.n4343 GND.n3404 240.244
R8125 GND.n4339 GND.n3404 240.244
R8126 GND.n4339 GND.n3410 240.244
R8127 GND.n4335 GND.n3410 240.244
R8128 GND.n4335 GND.n3412 240.244
R8129 GND.n4331 GND.n3412 240.244
R8130 GND.n4331 GND.n3418 240.244
R8131 GND.n4327 GND.n3418 240.244
R8132 GND.n4327 GND.n3420 240.244
R8133 GND.n4323 GND.n3420 240.244
R8134 GND.n4323 GND.n3426 240.244
R8135 GND.n4319 GND.n3426 240.244
R8136 GND.n4319 GND.n3428 240.244
R8137 GND.n4315 GND.n3428 240.244
R8138 GND.n4315 GND.n3434 240.244
R8139 GND.n4311 GND.n3434 240.244
R8140 GND.n4311 GND.n3436 240.244
R8141 GND.n4307 GND.n3436 240.244
R8142 GND.n4307 GND.n3442 240.244
R8143 GND.n4303 GND.n3442 240.244
R8144 GND.n4303 GND.n3444 240.244
R8145 GND.n4299 GND.n3444 240.244
R8146 GND.n4299 GND.n3450 240.244
R8147 GND.n4295 GND.n3450 240.244
R8148 GND.n4295 GND.n3452 240.244
R8149 GND.n4291 GND.n3452 240.244
R8150 GND.n4291 GND.n3458 240.244
R8151 GND.n4287 GND.n3458 240.244
R8152 GND.n4287 GND.n3460 240.244
R8153 GND.n4283 GND.n3460 240.244
R8154 GND.n4283 GND.n3466 240.244
R8155 GND.n4279 GND.n3466 240.244
R8156 GND.n4279 GND.n3468 240.244
R8157 GND.n4275 GND.n3468 240.244
R8158 GND.n4275 GND.n3474 240.244
R8159 GND.n4271 GND.n3474 240.244
R8160 GND.n4271 GND.n3476 240.244
R8161 GND.n4267 GND.n3476 240.244
R8162 GND.n4267 GND.n3482 240.244
R8163 GND.n4263 GND.n3482 240.244
R8164 GND.n4263 GND.n3484 240.244
R8165 GND.n4259 GND.n3484 240.244
R8166 GND.n4259 GND.n3490 240.244
R8167 GND.n4255 GND.n3490 240.244
R8168 GND.n4255 GND.n3492 240.244
R8169 GND.n4251 GND.n3492 240.244
R8170 GND.n4251 GND.n3498 240.244
R8171 GND.n4247 GND.n3498 240.244
R8172 GND.n4247 GND.n3500 240.244
R8173 GND.n4243 GND.n3500 240.244
R8174 GND.n4243 GND.n3506 240.244
R8175 GND.n4239 GND.n3506 240.244
R8176 GND.n4239 GND.n3508 240.244
R8177 GND.n4235 GND.n3508 240.244
R8178 GND.n4235 GND.n3514 240.244
R8179 GND.n4231 GND.n3514 240.244
R8180 GND.n4231 GND.n3516 240.244
R8181 GND.n4227 GND.n3516 240.244
R8182 GND.n4227 GND.n3522 240.244
R8183 GND.n4223 GND.n3522 240.244
R8184 GND.n4223 GND.n3524 240.244
R8185 GND.n4219 GND.n3524 240.244
R8186 GND.n4219 GND.n3530 240.244
R8187 GND.n4215 GND.n3530 240.244
R8188 GND.n4215 GND.n3532 240.244
R8189 GND.n4211 GND.n3532 240.244
R8190 GND.n4211 GND.n3538 240.244
R8191 GND.n4207 GND.n3538 240.244
R8192 GND.n4207 GND.n3540 240.244
R8193 GND.n4203 GND.n3540 240.244
R8194 GND.n4203 GND.n3546 240.244
R8195 GND.n4199 GND.n3546 240.244
R8196 GND.n4199 GND.n3548 240.244
R8197 GND.n4195 GND.n3548 240.244
R8198 GND.n4195 GND.n3554 240.244
R8199 GND.n4191 GND.n3554 240.244
R8200 GND.n4191 GND.n3556 240.244
R8201 GND.n4187 GND.n3556 240.244
R8202 GND.n4187 GND.n3562 240.244
R8203 GND.n4183 GND.n3562 240.244
R8204 GND.n4183 GND.n3564 240.244
R8205 GND.n4179 GND.n3564 240.244
R8206 GND.n4179 GND.n3570 240.244
R8207 GND.n4175 GND.n3570 240.244
R8208 GND.n4175 GND.n3572 240.244
R8209 GND.n4171 GND.n3572 240.244
R8210 GND.n4171 GND.n3578 240.244
R8211 GND.n4167 GND.n3578 240.244
R8212 GND.n4167 GND.n3580 240.244
R8213 GND.n4163 GND.n3580 240.244
R8214 GND.n4163 GND.n3586 240.244
R8215 GND.n4159 GND.n3586 240.244
R8216 GND.n4159 GND.n3588 240.244
R8217 GND.n4155 GND.n3588 240.244
R8218 GND.n4155 GND.n3594 240.244
R8219 GND.n4151 GND.n3594 240.244
R8220 GND.n4151 GND.n3596 240.244
R8221 GND.n4147 GND.n3596 240.244
R8222 GND.n4147 GND.n3602 240.244
R8223 GND.n4143 GND.n3602 240.244
R8224 GND.n4143 GND.n3604 240.244
R8225 GND.n4139 GND.n3604 240.244
R8226 GND.n4139 GND.n3610 240.244
R8227 GND.n4135 GND.n3610 240.244
R8228 GND.n4135 GND.n3612 240.244
R8229 GND.n4131 GND.n3612 240.244
R8230 GND.n4131 GND.n3618 240.244
R8231 GND.n4127 GND.n3618 240.244
R8232 GND.n4127 GND.n3620 240.244
R8233 GND.n4123 GND.n3620 240.244
R8234 GND.n4123 GND.n3626 240.244
R8235 GND.n4119 GND.n3626 240.244
R8236 GND.n4119 GND.n3628 240.244
R8237 GND.n4115 GND.n3628 240.244
R8238 GND.n4115 GND.n3634 240.244
R8239 GND.n4111 GND.n3634 240.244
R8240 GND.n4111 GND.n3636 240.244
R8241 GND.n4107 GND.n3636 240.244
R8242 GND.n4107 GND.n3642 240.244
R8243 GND.n4103 GND.n3642 240.244
R8244 GND.n4103 GND.n3644 240.244
R8245 GND.n4099 GND.n3644 240.244
R8246 GND.n4099 GND.n3650 240.244
R8247 GND.n4095 GND.n3650 240.244
R8248 GND.n4095 GND.n3652 240.244
R8249 GND.n4091 GND.n3652 240.244
R8250 GND.n4091 GND.n3658 240.244
R8251 GND.n4087 GND.n3658 240.244
R8252 GND.n4087 GND.n3660 240.244
R8253 GND.n4083 GND.n3660 240.244
R8254 GND.n4083 GND.n3666 240.244
R8255 GND.n4079 GND.n3666 240.244
R8256 GND.n4079 GND.n3668 240.244
R8257 GND.n4075 GND.n3668 240.244
R8258 GND.n4075 GND.n3674 240.244
R8259 GND.n4071 GND.n3674 240.244
R8260 GND.n4071 GND.n3676 240.244
R8261 GND.n4067 GND.n3676 240.244
R8262 GND.n4067 GND.n3682 240.244
R8263 GND.n4063 GND.n3682 240.244
R8264 GND.n4063 GND.n3684 240.244
R8265 GND.n4059 GND.n3684 240.244
R8266 GND.n4059 GND.n3690 240.244
R8267 GND.n4055 GND.n3690 240.244
R8268 GND.n4055 GND.n3692 240.244
R8269 GND.n4051 GND.n3692 240.244
R8270 GND.n4051 GND.n3698 240.244
R8271 GND.n4047 GND.n3698 240.244
R8272 GND.n4047 GND.n3700 240.244
R8273 GND.n4043 GND.n3700 240.244
R8274 GND.n4043 GND.n3706 240.244
R8275 GND.n4039 GND.n3706 240.244
R8276 GND.n4039 GND.n3708 240.244
R8277 GND.n4035 GND.n3708 240.244
R8278 GND.n4035 GND.n3714 240.244
R8279 GND.n4031 GND.n3714 240.244
R8280 GND.n4031 GND.n3716 240.244
R8281 GND.n4027 GND.n3716 240.244
R8282 GND.n4027 GND.n3722 240.244
R8283 GND.n4023 GND.n3722 240.244
R8284 GND.n4023 GND.n3724 240.244
R8285 GND.n4019 GND.n3724 240.244
R8286 GND.n4019 GND.n3730 240.244
R8287 GND.n4015 GND.n3730 240.244
R8288 GND.n4015 GND.n3732 240.244
R8289 GND.n4011 GND.n3732 240.244
R8290 GND.n4011 GND.n3738 240.244
R8291 GND.n4007 GND.n3738 240.244
R8292 GND.n4007 GND.n3740 240.244
R8293 GND.n4003 GND.n3740 240.244
R8294 GND.n4003 GND.n3746 240.244
R8295 GND.n3999 GND.n3746 240.244
R8296 GND.n3999 GND.n3748 240.244
R8297 GND.n3995 GND.n3748 240.244
R8298 GND.n3995 GND.n3754 240.244
R8299 GND.n3991 GND.n3754 240.244
R8300 GND.n3991 GND.n3756 240.244
R8301 GND.n3987 GND.n3756 240.244
R8302 GND.n3987 GND.n3762 240.244
R8303 GND.n3983 GND.n3762 240.244
R8304 GND.n3983 GND.n3764 240.244
R8305 GND.n3979 GND.n3764 240.244
R8306 GND.n3979 GND.n3770 240.244
R8307 GND.n3975 GND.n3770 240.244
R8308 GND.n3975 GND.n3772 240.244
R8309 GND.n3971 GND.n3772 240.244
R8310 GND.n3971 GND.n3778 240.244
R8311 GND.n3967 GND.n3778 240.244
R8312 GND.n3967 GND.n3780 240.244
R8313 GND.n3961 GND.n3785 240.244
R8314 GND.n3957 GND.n3785 240.244
R8315 GND.n3957 GND.n3787 240.244
R8316 GND.n3953 GND.n3787 240.244
R8317 GND.n3953 GND.n3792 240.244
R8318 GND.n3949 GND.n3792 240.244
R8319 GND.n3949 GND.n3794 240.244
R8320 GND.n3945 GND.n3794 240.244
R8321 GND.n3945 GND.n3800 240.244
R8322 GND.n3941 GND.n3800 240.244
R8323 GND.n3941 GND.n3802 240.244
R8324 GND.n3937 GND.n3802 240.244
R8325 GND.n3937 GND.n3808 240.244
R8326 GND.n3933 GND.n3808 240.244
R8327 GND.n3933 GND.n3810 240.244
R8328 GND.n3929 GND.n3810 240.244
R8329 GND.n3929 GND.n3816 240.244
R8330 GND.n3925 GND.n3816 240.244
R8331 GND.n3925 GND.n3818 240.244
R8332 GND.n3921 GND.n3818 240.244
R8333 GND.n3921 GND.n3824 240.244
R8334 GND.n3917 GND.n3824 240.244
R8335 GND.n3917 GND.n3826 240.244
R8336 GND.n3913 GND.n3826 240.244
R8337 GND.n3913 GND.n3832 240.244
R8338 GND.n3909 GND.n3832 240.244
R8339 GND.n3909 GND.n3834 240.244
R8340 GND.n3905 GND.n3834 240.244
R8341 GND.n3905 GND.n3840 240.244
R8342 GND.n3901 GND.n3840 240.244
R8343 GND.n3901 GND.n3842 240.244
R8344 GND.n3897 GND.n3842 240.244
R8345 GND.n3897 GND.n3848 240.244
R8346 GND.n3893 GND.n3848 240.244
R8347 GND.n3893 GND.n3850 240.244
R8348 GND.n3889 GND.n3850 240.244
R8349 GND.n3889 GND.n3856 240.244
R8350 GND.n3885 GND.n3856 240.244
R8351 GND.n3885 GND.n3858 240.244
R8352 GND.n3881 GND.n3858 240.244
R8353 GND.n3881 GND.n3864 240.244
R8354 GND.n3877 GND.n3864 240.244
R8355 GND.n3877 GND.n3866 240.244
R8356 GND.n3873 GND.n3866 240.244
R8357 GND.n3873 GND.n348 240.244
R8358 GND.n8451 GND.n348 240.244
R8359 GND.n8451 GND.n344 240.244
R8360 GND.n4851 GND.n2427 240.244
R8361 GND.n4851 GND.n2412 240.244
R8362 GND.n4865 GND.n2412 240.244
R8363 GND.n4865 GND.n2408 240.244
R8364 GND.n4871 GND.n2408 240.244
R8365 GND.n4871 GND.n2392 240.244
R8366 GND.n4885 GND.n2392 240.244
R8367 GND.n4885 GND.n2388 240.244
R8368 GND.n4891 GND.n2388 240.244
R8369 GND.n4891 GND.n2372 240.244
R8370 GND.n4905 GND.n2372 240.244
R8371 GND.n4905 GND.n2368 240.244
R8372 GND.n4911 GND.n2368 240.244
R8373 GND.n4911 GND.n2351 240.244
R8374 GND.n4925 GND.n2351 240.244
R8375 GND.n4925 GND.n2347 240.244
R8376 GND.n4931 GND.n2347 240.244
R8377 GND.n4931 GND.n2332 240.244
R8378 GND.n4945 GND.n2332 240.244
R8379 GND.n4945 GND.n2328 240.244
R8380 GND.n4951 GND.n2328 240.244
R8381 GND.n4951 GND.n2312 240.244
R8382 GND.n4965 GND.n2312 240.244
R8383 GND.n4965 GND.n2308 240.244
R8384 GND.n4971 GND.n2308 240.244
R8385 GND.n4971 GND.n2292 240.244
R8386 GND.n4985 GND.n2292 240.244
R8387 GND.n4985 GND.n2288 240.244
R8388 GND.n4991 GND.n2288 240.244
R8389 GND.n4991 GND.n2272 240.244
R8390 GND.n5005 GND.n2272 240.244
R8391 GND.n5005 GND.n2268 240.244
R8392 GND.n5012 GND.n2268 240.244
R8393 GND.n5012 GND.n2251 240.244
R8394 GND.n5031 GND.n2251 240.244
R8395 GND.n5031 GND.n2248 240.244
R8396 GND.n5035 GND.n2248 240.244
R8397 GND.n5037 GND.n5035 240.244
R8398 GND.n5037 GND.n2225 240.244
R8399 GND.n5051 GND.n2225 240.244
R8400 GND.n5052 GND.n5051 240.244
R8401 GND.n5055 GND.n5052 240.244
R8402 GND.n5055 GND.n2202 240.244
R8403 GND.n5076 GND.n2202 240.244
R8404 GND.n5077 GND.n5076 240.244
R8405 GND.n5080 GND.n5077 240.244
R8406 GND.n5080 GND.n2076 240.244
R8407 GND.n5089 GND.n2076 240.244
R8408 GND.n5089 GND.n2060 240.244
R8409 GND.n5108 GND.n2060 240.244
R8410 GND.n5108 GND.n2055 240.244
R8411 GND.n5116 GND.n2055 240.244
R8412 GND.n5116 GND.n2056 240.244
R8413 GND.n2056 GND.n2033 240.244
R8414 GND.n5199 GND.n2033 240.244
R8415 GND.n5199 GND.n2029 240.244
R8416 GND.n5205 GND.n2029 240.244
R8417 GND.n5205 GND.n2013 240.244
R8418 GND.n5219 GND.n2013 240.244
R8419 GND.n5219 GND.n2009 240.244
R8420 GND.n5225 GND.n2009 240.244
R8421 GND.n5225 GND.n1993 240.244
R8422 GND.n5239 GND.n1993 240.244
R8423 GND.n5239 GND.n1989 240.244
R8424 GND.n5245 GND.n1989 240.244
R8425 GND.n5245 GND.n1973 240.244
R8426 GND.n5259 GND.n1973 240.244
R8427 GND.n5259 GND.n1969 240.244
R8428 GND.n5265 GND.n1969 240.244
R8429 GND.n5265 GND.n1953 240.244
R8430 GND.n5279 GND.n1953 240.244
R8431 GND.n5279 GND.n1949 240.244
R8432 GND.n5285 GND.n1949 240.244
R8433 GND.n5285 GND.n1933 240.244
R8434 GND.n5299 GND.n1933 240.244
R8435 GND.n5299 GND.n1929 240.244
R8436 GND.n5305 GND.n1929 240.244
R8437 GND.n5305 GND.n1913 240.244
R8438 GND.n5324 GND.n1913 240.244
R8439 GND.n5324 GND.n1908 240.244
R8440 GND.n5332 GND.n1908 240.244
R8441 GND.n5332 GND.n1909 240.244
R8442 GND.n1909 GND.n1886 240.244
R8443 GND.n5369 GND.n1886 240.244
R8444 GND.n5369 GND.n1882 240.244
R8445 GND.n5377 GND.n1882 240.244
R8446 GND.n5377 GND.n1868 240.244
R8447 GND.n5388 GND.n1868 240.244
R8448 GND.n5389 GND.n5388 240.244
R8449 GND.n5389 GND.n1631 240.244
R8450 GND.n5395 GND.n1631 240.244
R8451 GND.n5396 GND.n5395 240.244
R8452 GND.n5397 GND.n5396 240.244
R8453 GND.n5397 GND.n1861 240.244
R8454 GND.n5405 GND.n1861 240.244
R8455 GND.n5406 GND.n5405 240.244
R8456 GND.n5407 GND.n5406 240.244
R8457 GND.n5407 GND.n1856 240.244
R8458 GND.n6189 GND.n1856 240.244
R8459 GND.n6189 GND.n1857 240.244
R8460 GND.n6185 GND.n1857 240.244
R8461 GND.n6185 GND.n5415 240.244
R8462 GND.n6175 GND.n5415 240.244
R8463 GND.n6175 GND.n5427 240.244
R8464 GND.n6171 GND.n5427 240.244
R8465 GND.n6171 GND.n5433 240.244
R8466 GND.n5520 GND.n5433 240.244
R8467 GND.n6156 GND.n5520 240.244
R8468 GND.n6156 GND.n5521 240.244
R8469 GND.n6152 GND.n5521 240.244
R8470 GND.n6152 GND.n5529 240.244
R8471 GND.n6142 GND.n5529 240.244
R8472 GND.n6142 GND.n5541 240.244
R8473 GND.n6138 GND.n5541 240.244
R8474 GND.n6138 GND.n5547 240.244
R8475 GND.n6128 GND.n5547 240.244
R8476 GND.n6128 GND.n5559 240.244
R8477 GND.n6124 GND.n5559 240.244
R8478 GND.n6124 GND.n5565 240.244
R8479 GND.n6114 GND.n5565 240.244
R8480 GND.n6114 GND.n5577 240.244
R8481 GND.n6110 GND.n5577 240.244
R8482 GND.n6110 GND.n5583 240.244
R8483 GND.n5651 GND.n5583 240.244
R8484 GND.n6095 GND.n5651 240.244
R8485 GND.n6095 GND.n5652 240.244
R8486 GND.n6091 GND.n5652 240.244
R8487 GND.n6091 GND.n5660 240.244
R8488 GND.n6081 GND.n5660 240.244
R8489 GND.n6081 GND.n5672 240.244
R8490 GND.n6077 GND.n5672 240.244
R8491 GND.n6077 GND.n5678 240.244
R8492 GND.n6067 GND.n5678 240.244
R8493 GND.n6067 GND.n5690 240.244
R8494 GND.n6063 GND.n5690 240.244
R8495 GND.n6063 GND.n5696 240.244
R8496 GND.n6053 GND.n5696 240.244
R8497 GND.n6053 GND.n5708 240.244
R8498 GND.n6049 GND.n5708 240.244
R8499 GND.n6049 GND.n5714 240.244
R8500 GND.n5782 GND.n5714 240.244
R8501 GND.n6034 GND.n5782 240.244
R8502 GND.n6034 GND.n5783 240.244
R8503 GND.n6030 GND.n5783 240.244
R8504 GND.n6030 GND.n5791 240.244
R8505 GND.n6020 GND.n5791 240.244
R8506 GND.n6020 GND.n5802 240.244
R8507 GND.n6016 GND.n5802 240.244
R8508 GND.n6016 GND.n5808 240.244
R8509 GND.n6006 GND.n5808 240.244
R8510 GND.n6006 GND.n5820 240.244
R8511 GND.n6002 GND.n5820 240.244
R8512 GND.n6002 GND.n5826 240.244
R8513 GND.n5992 GND.n5826 240.244
R8514 GND.n5992 GND.n5838 240.244
R8515 GND.n5988 GND.n5838 240.244
R8516 GND.n5988 GND.n5844 240.244
R8517 GND.n5913 GND.n5844 240.244
R8518 GND.n5973 GND.n5913 240.244
R8519 GND.n5973 GND.n5914 240.244
R8520 GND.n5969 GND.n5914 240.244
R8521 GND.n5969 GND.n5922 240.244
R8522 GND.n5959 GND.n5922 240.244
R8523 GND.n5959 GND.n5953 240.244
R8524 GND.n5953 GND.n1585 240.244
R8525 GND.n6432 GND.n1585 240.244
R8526 GND.n6432 GND.n1580 240.244
R8527 GND.n6440 GND.n1580 240.244
R8528 GND.n6440 GND.n1581 240.244
R8529 GND.n1581 GND.n1554 240.244
R8530 GND.n6469 GND.n1554 240.244
R8531 GND.n6469 GND.n1549 240.244
R8532 GND.n6480 GND.n1549 240.244
R8533 GND.n6480 GND.n1550 240.244
R8534 GND.n6476 GND.n1550 240.244
R8535 GND.n6476 GND.n1516 240.244
R8536 GND.n6529 GND.n1516 240.244
R8537 GND.n6529 GND.n1511 240.244
R8538 GND.n6543 GND.n1511 240.244
R8539 GND.n6543 GND.n1512 240.244
R8540 GND.n6539 GND.n1512 240.244
R8541 GND.n6539 GND.n6538 240.244
R8542 GND.n6538 GND.n1473 240.244
R8543 GND.n6607 GND.n1473 240.244
R8544 GND.n6607 GND.n1468 240.244
R8545 GND.n6618 GND.n1468 240.244
R8546 GND.n6618 GND.n1469 240.244
R8547 GND.n6614 GND.n1469 240.244
R8548 GND.n6614 GND.n1418 240.244
R8549 GND.n6686 GND.n1418 240.244
R8550 GND.n6686 GND.n1414 240.244
R8551 GND.n6692 GND.n1414 240.244
R8552 GND.n6692 GND.n1395 240.244
R8553 GND.n6715 GND.n1395 240.244
R8554 GND.n6715 GND.n1390 240.244
R8555 GND.n6752 GND.n1390 240.244
R8556 GND.n6752 GND.n1391 240.244
R8557 GND.n6748 GND.n1391 240.244
R8558 GND.n6748 GND.n6747 240.244
R8559 GND.n6747 GND.n6745 240.244
R8560 GND.n6745 GND.n6723 240.244
R8561 GND.n6741 GND.n6723 240.244
R8562 GND.n6741 GND.n6739 240.244
R8563 GND.n6739 GND.n6738 240.244
R8564 GND.n6738 GND.n6729 240.244
R8565 GND.n6734 GND.n6729 240.244
R8566 GND.n6734 GND.n1307 240.244
R8567 GND.n6888 GND.n1307 240.244
R8568 GND.n6888 GND.n1302 240.244
R8569 GND.n6908 GND.n1302 240.244
R8570 GND.n6908 GND.n1303 240.244
R8571 GND.n6904 GND.n1303 240.244
R8572 GND.n6904 GND.n6903 240.244
R8573 GND.n6903 GND.n6902 240.244
R8574 GND.n6902 GND.n6896 240.244
R8575 GND.n6896 GND.n1154 240.244
R8576 GND.n7011 GND.n1154 240.244
R8577 GND.n7011 GND.n1149 240.244
R8578 GND.n7025 GND.n1149 240.244
R8579 GND.n7025 GND.n1150 240.244
R8580 GND.n7021 GND.n1150 240.244
R8581 GND.n7021 GND.n7020 240.244
R8582 GND.n7020 GND.n1123 240.244
R8583 GND.n7057 GND.n1123 240.244
R8584 GND.n7057 GND.n1118 240.244
R8585 GND.n7074 GND.n1118 240.244
R8586 GND.n7074 GND.n1119 240.244
R8587 GND.n7070 GND.n1119 240.244
R8588 GND.n7070 GND.n7069 240.244
R8589 GND.n7069 GND.n7068 240.244
R8590 GND.n7068 GND.n1089 240.244
R8591 GND.n7115 GND.n1089 240.244
R8592 GND.n7115 GND.n1084 240.244
R8593 GND.n7123 GND.n1084 240.244
R8594 GND.n7123 GND.n1085 240.244
R8595 GND.n1085 GND.n1064 240.244
R8596 GND.n7150 GND.n1064 240.244
R8597 GND.n7150 GND.n1059 240.244
R8598 GND.n7161 GND.n1059 240.244
R8599 GND.n7161 GND.n1060 240.244
R8600 GND.n7157 GND.n1060 240.244
R8601 GND.n7157 GND.n1040 240.244
R8602 GND.n7189 GND.n1040 240.244
R8603 GND.n7189 GND.n1035 240.244
R8604 GND.n7206 GND.n1035 240.244
R8605 GND.n7206 GND.n1036 240.244
R8606 GND.n7202 GND.n1036 240.244
R8607 GND.n7202 GND.n7201 240.244
R8608 GND.n7201 GND.n7200 240.244
R8609 GND.n7200 GND.n1006 240.244
R8610 GND.n7247 GND.n1006 240.244
R8611 GND.n7247 GND.n1001 240.244
R8612 GND.n7255 GND.n1001 240.244
R8613 GND.n7255 GND.n1002 240.244
R8614 GND.n1002 GND.n981 240.244
R8615 GND.n7282 GND.n981 240.244
R8616 GND.n7282 GND.n976 240.244
R8617 GND.n7293 GND.n976 240.244
R8618 GND.n7293 GND.n977 240.244
R8619 GND.n7289 GND.n977 240.244
R8620 GND.n7289 GND.n956 240.244
R8621 GND.n7320 GND.n956 240.244
R8622 GND.n7320 GND.n951 240.244
R8623 GND.n7328 GND.n951 240.244
R8624 GND.n7328 GND.n952 240.244
R8625 GND.n952 GND.n931 240.244
R8626 GND.n7355 GND.n931 240.244
R8627 GND.n7355 GND.n927 240.244
R8628 GND.n7361 GND.n927 240.244
R8629 GND.n7361 GND.n914 240.244
R8630 GND.n7379 GND.n914 240.244
R8631 GND.n7379 GND.n909 240.244
R8632 GND.n7387 GND.n909 240.244
R8633 GND.n7387 GND.n910 240.244
R8634 GND.n910 GND.n891 240.244
R8635 GND.n7415 GND.n891 240.244
R8636 GND.n7415 GND.n887 240.244
R8637 GND.n7421 GND.n887 240.244
R8638 GND.n7421 GND.n874 240.244
R8639 GND.n7485 GND.n874 240.244
R8640 GND.n7485 GND.n869 240.244
R8641 GND.n7504 GND.n869 240.244
R8642 GND.n7504 GND.n870 240.244
R8643 GND.n7500 GND.n870 240.244
R8644 GND.n7500 GND.n7499 240.244
R8645 GND.n7499 GND.n7496 240.244
R8646 GND.n7496 GND.n678 240.244
R8647 GND.n7703 GND.n678 240.244
R8648 GND.n7703 GND.n674 240.244
R8649 GND.n7709 GND.n674 240.244
R8650 GND.n7709 GND.n657 240.244
R8651 GND.n7725 GND.n657 240.244
R8652 GND.n7725 GND.n653 240.244
R8653 GND.n7731 GND.n653 240.244
R8654 GND.n7731 GND.n637 240.244
R8655 GND.n7745 GND.n637 240.244
R8656 GND.n7745 GND.n633 240.244
R8657 GND.n7751 GND.n633 240.244
R8658 GND.n7751 GND.n617 240.244
R8659 GND.n7765 GND.n617 240.244
R8660 GND.n7765 GND.n613 240.244
R8661 GND.n7771 GND.n613 240.244
R8662 GND.n7771 GND.n597 240.244
R8663 GND.n7785 GND.n597 240.244
R8664 GND.n7785 GND.n593 240.244
R8665 GND.n7791 GND.n593 240.244
R8666 GND.n7791 GND.n576 240.244
R8667 GND.n7809 GND.n576 240.244
R8668 GND.n7809 GND.n571 240.244
R8669 GND.n7817 GND.n571 240.244
R8670 GND.n7817 GND.n572 240.244
R8671 GND.n572 GND.n549 240.244
R8672 GND.n7883 GND.n549 240.244
R8673 GND.n7883 GND.n545 240.244
R8674 GND.n7889 GND.n545 240.244
R8675 GND.n7889 GND.n529 240.244
R8676 GND.n7903 GND.n529 240.244
R8677 GND.n7903 GND.n525 240.244
R8678 GND.n7909 GND.n525 240.244
R8679 GND.n7909 GND.n509 240.244
R8680 GND.n7923 GND.n509 240.244
R8681 GND.n7923 GND.n505 240.244
R8682 GND.n7929 GND.n505 240.244
R8683 GND.n7929 GND.n488 240.244
R8684 GND.n7950 GND.n488 240.244
R8685 GND.n7950 GND.n484 240.244
R8686 GND.n7956 GND.n484 240.244
R8687 GND.n7956 GND.n118 240.244
R8688 GND.n8601 GND.n118 240.244
R8689 GND.n8601 GND.n114 240.244
R8690 GND.n8607 GND.n114 240.244
R8691 GND.n8607 GND.n86 240.244
R8692 GND.n8631 GND.n86 240.244
R8693 GND.n8631 GND.n87 240.244
R8694 GND.n8623 GND.n87 240.244
R8695 GND.n8623 GND.n8620 240.244
R8696 GND.n8620 GND.n73 240.244
R8697 GND.n8636 GND.n73 240.244
R8698 GND.n8636 GND.n74 240.244
R8699 GND.n8578 GND.n74 240.244
R8700 GND.n8578 GND.n8576 240.244
R8701 GND.n8576 GND.n8573 240.244
R8702 GND.n8573 GND.n139 240.244
R8703 GND.n8565 GND.n139 240.244
R8704 GND.n8565 GND.n156 240.244
R8705 GND.n8561 GND.n156 240.244
R8706 GND.n8561 GND.n161 240.244
R8707 GND.n8553 GND.n161 240.244
R8708 GND.n8553 GND.n176 240.244
R8709 GND.n8549 GND.n176 240.244
R8710 GND.n8549 GND.n182 240.244
R8711 GND.n8541 GND.n182 240.244
R8712 GND.n8541 GND.n197 240.244
R8713 GND.n8537 GND.n197 240.244
R8714 GND.n8537 GND.n203 240.244
R8715 GND.n8529 GND.n203 240.244
R8716 GND.n8529 GND.n218 240.244
R8717 GND.n8525 GND.n218 240.244
R8718 GND.n8525 GND.n224 240.244
R8719 GND.n8517 GND.n224 240.244
R8720 GND.n8517 GND.n239 240.244
R8721 GND.n8513 GND.n239 240.244
R8722 GND.n8513 GND.n245 240.244
R8723 GND.n8505 GND.n245 240.244
R8724 GND.n8505 GND.n260 240.244
R8725 GND.n8501 GND.n260 240.244
R8726 GND.n8501 GND.n266 240.244
R8727 GND.n8493 GND.n266 240.244
R8728 GND.n8493 GND.n281 240.244
R8729 GND.n8489 GND.n281 240.244
R8730 GND.n8489 GND.n287 240.244
R8731 GND.n8481 GND.n287 240.244
R8732 GND.n8481 GND.n302 240.244
R8733 GND.n8477 GND.n302 240.244
R8734 GND.n8477 GND.n308 240.244
R8735 GND.n8469 GND.n308 240.244
R8736 GND.n8469 GND.n323 240.244
R8737 GND.n8465 GND.n323 240.244
R8738 GND.n8465 GND.n329 240.244
R8739 GND.n8457 GND.n329 240.244
R8740 GND.n4733 GND.n4731 240.244
R8741 GND.n4739 GND.n3018 240.244
R8742 GND.n4743 GND.n4741 240.244
R8743 GND.n4749 GND.n3014 240.244
R8744 GND.n4753 GND.n4751 240.244
R8745 GND.n4759 GND.n3010 240.244
R8746 GND.n4763 GND.n4761 240.244
R8747 GND.n4769 GND.n3006 240.244
R8748 GND.n4773 GND.n4771 240.244
R8749 GND.n4779 GND.n3002 240.244
R8750 GND.n4783 GND.n4781 240.244
R8751 GND.n4789 GND.n2998 240.244
R8752 GND.n4793 GND.n4791 240.244
R8753 GND.n4799 GND.n2994 240.244
R8754 GND.n4803 GND.n4801 240.244
R8755 GND.n4809 GND.n2990 240.244
R8756 GND.n4813 GND.n4811 240.244
R8757 GND.n4819 GND.n2986 240.244
R8758 GND.n4823 GND.n4821 240.244
R8759 GND.n4829 GND.n2982 240.244
R8760 GND.n4833 GND.n4831 240.244
R8761 GND.n4840 GND.n2978 240.244
R8762 GND.n4843 GND.n4842 240.244
R8763 GND.n2863 GND.n2536 240.244
R8764 GND.n2612 GND.n2536 240.244
R8765 GND.n2612 GND.n2611 240.244
R8766 GND.n2611 GND.n2563 240.244
R8767 GND.n2563 GND.n2562 240.244
R8768 GND.n2562 GND.n2423 240.244
R8769 GND.n4853 GND.n2423 240.244
R8770 GND.n4854 GND.n4853 240.244
R8771 GND.n4854 GND.n2415 240.244
R8772 GND.n2415 GND.n2403 240.244
R8773 GND.n4873 GND.n2403 240.244
R8774 GND.n4874 GND.n4873 240.244
R8775 GND.n4874 GND.n2395 240.244
R8776 GND.n2395 GND.n2383 240.244
R8777 GND.n4893 GND.n2383 240.244
R8778 GND.n4894 GND.n4893 240.244
R8779 GND.n4894 GND.n2375 240.244
R8780 GND.n2375 GND.n2363 240.244
R8781 GND.n4913 GND.n2363 240.244
R8782 GND.n4914 GND.n4913 240.244
R8783 GND.n4914 GND.n2354 240.244
R8784 GND.n2354 GND.n2343 240.244
R8785 GND.n4933 GND.n2343 240.244
R8786 GND.n4934 GND.n4933 240.244
R8787 GND.n4934 GND.n2335 240.244
R8788 GND.n2335 GND.n2323 240.244
R8789 GND.n4953 GND.n2323 240.244
R8790 GND.n4954 GND.n4953 240.244
R8791 GND.n4954 GND.n2315 240.244
R8792 GND.n2315 GND.n2303 240.244
R8793 GND.n4973 GND.n2303 240.244
R8794 GND.n4974 GND.n4973 240.244
R8795 GND.n4974 GND.n2295 240.244
R8796 GND.n2295 GND.n2283 240.244
R8797 GND.n4993 GND.n2283 240.244
R8798 GND.n4994 GND.n4993 240.244
R8799 GND.n4994 GND.n2275 240.244
R8800 GND.n2275 GND.n2263 240.244
R8801 GND.n5014 GND.n2263 240.244
R8802 GND.n5015 GND.n5014 240.244
R8803 GND.n5015 GND.n2254 240.244
R8804 GND.n5018 GND.n2254 240.244
R8805 GND.n5018 GND.n2240 240.244
R8806 GND.n5039 GND.n2240 240.244
R8807 GND.n5040 GND.n5039 240.244
R8808 GND.n5040 GND.n2232 240.244
R8809 GND.n2232 GND.n2217 240.244
R8810 GND.n5056 GND.n2217 240.244
R8811 GND.n5057 GND.n5056 240.244
R8812 GND.n5057 GND.n2209 240.244
R8813 GND.n5060 GND.n2209 240.244
R8814 GND.n5060 GND.n2199 240.244
R8815 GND.n2199 GND.n2071 240.244
R8816 GND.n5091 GND.n2071 240.244
R8817 GND.n5092 GND.n5091 240.244
R8818 GND.n5092 GND.n2063 240.244
R8819 GND.n5095 GND.n2063 240.244
R8820 GND.n5095 GND.n2053 240.244
R8821 GND.n2053 GND.n2043 240.244
R8822 GND.n5188 GND.n2043 240.244
R8823 GND.n5188 GND.n2035 240.244
R8824 GND.n2035 GND.n2024 240.244
R8825 GND.n5207 GND.n2024 240.244
R8826 GND.n5208 GND.n5207 240.244
R8827 GND.n5208 GND.n2016 240.244
R8828 GND.n2016 GND.n2004 240.244
R8829 GND.n5227 GND.n2004 240.244
R8830 GND.n5228 GND.n5227 240.244
R8831 GND.n5228 GND.n1996 240.244
R8832 GND.n1996 GND.n1984 240.244
R8833 GND.n5247 GND.n1984 240.244
R8834 GND.n5248 GND.n5247 240.244
R8835 GND.n5248 GND.n1976 240.244
R8836 GND.n1976 GND.n1964 240.244
R8837 GND.n5267 GND.n1964 240.244
R8838 GND.n5268 GND.n5267 240.244
R8839 GND.n5268 GND.n1956 240.244
R8840 GND.n1956 GND.n1944 240.244
R8841 GND.n5287 GND.n1944 240.244
R8842 GND.n5288 GND.n5287 240.244
R8843 GND.n5288 GND.n1936 240.244
R8844 GND.n1936 GND.n1924 240.244
R8845 GND.n5307 GND.n1924 240.244
R8846 GND.n5308 GND.n5307 240.244
R8847 GND.n5308 GND.n1916 240.244
R8848 GND.n5311 GND.n1916 240.244
R8849 GND.n5311 GND.n1906 240.244
R8850 GND.n1906 GND.n1896 240.244
R8851 GND.n5358 GND.n1896 240.244
R8852 GND.n5358 GND.n1888 240.244
R8853 GND.n1888 GND.n1877 240.244
R8854 GND.n5379 GND.n1877 240.244
R8855 GND.n5380 GND.n5379 240.244
R8856 GND.n5380 GND.n1871 240.244
R8857 GND.n1871 GND.n1635 240.244
R8858 GND.n6285 GND.n1635 240.244
R8859 GND.n2587 GND.n2586 240.244
R8860 GND.n2585 GND.n2584 240.244
R8861 GND.n2595 GND.n2594 240.244
R8862 GND.n2581 GND.n2580 240.244
R8863 GND.n2576 GND.n2462 240.244
R8864 GND.n2604 GND.n2573 240.244
R8865 GND.n2610 GND.n2573 240.244
R8866 GND.n2610 GND.n2559 240.244
R8867 GND.n2717 GND.n2559 240.244
R8868 GND.n2717 GND.n2554 240.244
R8869 GND.n2847 GND.n2554 240.244
R8870 GND.n2847 GND.n2425 240.244
R8871 GND.n2722 GND.n2425 240.244
R8872 GND.n2722 GND.n2416 240.244
R8873 GND.n2723 GND.n2416 240.244
R8874 GND.n2723 GND.n2406 240.244
R8875 GND.n2726 GND.n2406 240.244
R8876 GND.n2726 GND.n2396 240.244
R8877 GND.n2727 GND.n2396 240.244
R8878 GND.n2727 GND.n2386 240.244
R8879 GND.n2730 GND.n2386 240.244
R8880 GND.n2730 GND.n2376 240.244
R8881 GND.n2731 GND.n2376 240.244
R8882 GND.n2731 GND.n2366 240.244
R8883 GND.n2734 GND.n2366 240.244
R8884 GND.n2734 GND.n2356 240.244
R8885 GND.n2735 GND.n2356 240.244
R8886 GND.n2735 GND.n2345 240.244
R8887 GND.n2738 GND.n2345 240.244
R8888 GND.n2738 GND.n2336 240.244
R8889 GND.n2739 GND.n2336 240.244
R8890 GND.n2739 GND.n2326 240.244
R8891 GND.n2742 GND.n2326 240.244
R8892 GND.n2742 GND.n2316 240.244
R8893 GND.n2743 GND.n2316 240.244
R8894 GND.n2743 GND.n2306 240.244
R8895 GND.n2746 GND.n2306 240.244
R8896 GND.n2746 GND.n2296 240.244
R8897 GND.n2747 GND.n2296 240.244
R8898 GND.n2747 GND.n2286 240.244
R8899 GND.n2750 GND.n2286 240.244
R8900 GND.n2750 GND.n2276 240.244
R8901 GND.n2751 GND.n2276 240.244
R8902 GND.n2751 GND.n2266 240.244
R8903 GND.n2754 GND.n2266 240.244
R8904 GND.n2754 GND.n2256 240.244
R8905 GND.n2755 GND.n2256 240.244
R8906 GND.n2756 GND.n2755 240.244
R8907 GND.n2756 GND.n2246 240.244
R8908 GND.n2759 GND.n2246 240.244
R8909 GND.n2759 GND.n2233 240.244
R8910 GND.n2760 GND.n2233 240.244
R8911 GND.n2760 GND.n2224 240.244
R8912 GND.n2780 GND.n2224 240.244
R8913 GND.n2780 GND.n2210 240.244
R8914 GND.n2777 GND.n2210 240.244
R8915 GND.n2777 GND.n2200 240.244
R8916 GND.n2774 GND.n2200 240.244
R8917 GND.n2774 GND.n2074 240.244
R8918 GND.n2771 GND.n2074 240.244
R8919 GND.n2771 GND.n2064 240.244
R8920 GND.n2064 GND.n2050 240.244
R8921 GND.n5118 GND.n2050 240.244
R8922 GND.n5118 GND.n2046 240.244
R8923 GND.n5186 GND.n2046 240.244
R8924 GND.n5186 GND.n2036 240.244
R8925 GND.n5182 GND.n2036 240.244
R8926 GND.n5182 GND.n2027 240.244
R8927 GND.n5179 GND.n2027 240.244
R8928 GND.n5179 GND.n2017 240.244
R8929 GND.n5176 GND.n2017 240.244
R8930 GND.n5176 GND.n2007 240.244
R8931 GND.n5173 GND.n2007 240.244
R8932 GND.n5173 GND.n1997 240.244
R8933 GND.n5170 GND.n1997 240.244
R8934 GND.n5170 GND.n1987 240.244
R8935 GND.n5167 GND.n1987 240.244
R8936 GND.n5167 GND.n1977 240.244
R8937 GND.n5164 GND.n1977 240.244
R8938 GND.n5164 GND.n1967 240.244
R8939 GND.n5161 GND.n1967 240.244
R8940 GND.n5161 GND.n1957 240.244
R8941 GND.n5158 GND.n1957 240.244
R8942 GND.n5158 GND.n1947 240.244
R8943 GND.n5155 GND.n1947 240.244
R8944 GND.n5155 GND.n1937 240.244
R8945 GND.n5152 GND.n1937 240.244
R8946 GND.n5152 GND.n1927 240.244
R8947 GND.n5149 GND.n1927 240.244
R8948 GND.n5149 GND.n1917 240.244
R8949 GND.n1917 GND.n1903 240.244
R8950 GND.n5334 GND.n1903 240.244
R8951 GND.n5334 GND.n1899 240.244
R8952 GND.n5356 GND.n1899 240.244
R8953 GND.n5356 GND.n1889 240.244
R8954 GND.n5352 GND.n1889 240.244
R8955 GND.n5352 GND.n1880 240.244
R8956 GND.n5349 GND.n1880 240.244
R8957 GND.n5349 GND.n1872 240.244
R8958 GND.n5346 GND.n1872 240.244
R8959 GND.n5346 GND.n1633 240.244
R8960 GND.n1640 GND.n1636 240.244
R8961 GND.n1645 GND.n1642 240.244
R8962 GND.n1650 GND.n1647 240.244
R8963 GND.n1654 GND.n1653 240.244
R8964 GND.n1660 GND.n1659 240.244
R8965 GND.n7511 GND.t105 223.19
R8966 GND.n6195 GND.t177 223.19
R8967 GND.n5441 GND.t146 223.19
R8968 GND.n7434 GND.t113 223.19
R8969 GND.n8449 GND.n8448 212.637
R8970 GND.n2577 GND.t88 210.603
R8971 GND.n1702 GND.t143 210.603
R8972 GND.n1721 GND.t137 210.603
R8973 GND.n1735 GND.t140 210.603
R8974 GND.n1754 GND.t153 210.603
R8975 GND.n1772 GND.t125 210.603
R8976 GND.n816 GND.t168 210.603
R8977 GND.n830 GND.t165 210.603
R8978 GND.n7568 GND.t162 210.603
R8979 GND.n7582 GND.t156 210.603
R8980 GND.n7595 GND.t174 210.603
R8981 GND.n442 GND.t109 210.603
R8982 GND.n429 GND.t183 210.603
R8983 GND.n418 GND.t116 210.603
R8984 GND.n405 GND.t119 210.603
R8985 GND.n394 GND.t122 210.603
R8986 GND.n8184 GND.t159 210.603
R8987 GND.n1206 GND.t133 210.603
R8988 GND.n2477 GND.t102 210.603
R8989 GND.n2491 GND.t99 210.603
R8990 GND.n2504 GND.t96 210.603
R8991 GND.n2518 GND.t180 210.603
R8992 GND.n2531 GND.t150 210.603
R8993 GND.n1656 GND.t171 210.603
R8994 GND.n3960 GND.n3959 207.156
R8995 GND.n3959 GND.n3958 207.156
R8996 GND.n3958 GND.n3786 207.156
R8997 GND.n3952 GND.n3786 207.156
R8998 GND.n3952 GND.n3951 207.156
R8999 GND.n3951 GND.n3950 207.156
R9000 GND.n3950 GND.n3793 207.156
R9001 GND.n3944 GND.n3793 207.156
R9002 GND.n3944 GND.n3943 207.156
R9003 GND.n3943 GND.n3942 207.156
R9004 GND.n3942 GND.n3801 207.156
R9005 GND.n3936 GND.n3801 207.156
R9006 GND.n3936 GND.n3935 207.156
R9007 GND.n3935 GND.n3934 207.156
R9008 GND.n3934 GND.n3809 207.156
R9009 GND.n3928 GND.n3809 207.156
R9010 GND.n3928 GND.n3927 207.156
R9011 GND.n3927 GND.n3926 207.156
R9012 GND.n3926 GND.n3817 207.156
R9013 GND.n3920 GND.n3817 207.156
R9014 GND.n3920 GND.n3919 207.156
R9015 GND.n3919 GND.n3918 207.156
R9016 GND.n3918 GND.n3825 207.156
R9017 GND.n3912 GND.n3825 207.156
R9018 GND.n3912 GND.n3911 207.156
R9019 GND.n3911 GND.n3910 207.156
R9020 GND.n3910 GND.n3833 207.156
R9021 GND.n3904 GND.n3833 207.156
R9022 GND.n3904 GND.n3903 207.156
R9023 GND.n3903 GND.n3902 207.156
R9024 GND.n3902 GND.n3841 207.156
R9025 GND.n3896 GND.n3841 207.156
R9026 GND.n3896 GND.n3895 207.156
R9027 GND.n3895 GND.n3894 207.156
R9028 GND.n3894 GND.n3849 207.156
R9029 GND.n3888 GND.n3849 207.156
R9030 GND.n3888 GND.n3887 207.156
R9031 GND.n3887 GND.n3886 207.156
R9032 GND.n3886 GND.n3857 207.156
R9033 GND.n3880 GND.n3857 207.156
R9034 GND.n3880 GND.n3879 207.156
R9035 GND.n3879 GND.n3878 207.156
R9036 GND.n3878 GND.n3865 207.156
R9037 GND.n3872 GND.n3865 207.156
R9038 GND.n3872 GND.n349 207.156
R9039 GND.n8450 GND.n349 207.156
R9040 GND.n8450 GND.n8449 207.156
R9041 GND.n7560 GND.n690 199.319
R9042 GND.n7560 GND.n691 199.319
R9043 GND.n1819 GND.n1677 199.319
R9044 GND.n1819 GND.n1676 199.319
R9045 GND.n7568 GND.t164 198.947
R9046 GND.n7582 GND.t158 198.947
R9047 GND.n429 GND.t184 198.947
R9048 GND.n2577 GND.t91 189.347
R9049 GND.n1702 GND.t144 189.347
R9050 GND.n1721 GND.t138 189.347
R9051 GND.n1735 GND.t141 189.347
R9052 GND.n1754 GND.t154 189.347
R9053 GND.n1772 GND.t127 189.347
R9054 GND.n816 GND.t170 189.347
R9055 GND.n830 GND.t167 189.347
R9056 GND.n7595 GND.t176 189.347
R9057 GND.n442 GND.t111 189.347
R9058 GND.n418 GND.t117 189.347
R9059 GND.n405 GND.t120 189.347
R9060 GND.n394 GND.t123 189.347
R9061 GND.n8184 GND.t160 189.347
R9062 GND.n1206 GND.t136 189.347
R9063 GND.n2477 GND.t104 189.347
R9064 GND.n2491 GND.t101 189.347
R9065 GND.n2504 GND.t98 189.347
R9066 GND.n2518 GND.t182 189.347
R9067 GND.n2531 GND.t152 189.347
R9068 GND.n1656 GND.t172 189.347
R9069 GND.n3026 GND.n2976 181.487
R9070 GND.n5441 GND.t149 172.393
R9071 GND.n7434 GND.t114 172.393
R9072 GND.n7511 GND.t107 172.392
R9073 GND.n6195 GND.t179 172.392
R9074 GND.n7555 GND.n863 163.367
R9075 GND.n7551 GND.n7550 163.367
R9076 GND.n7547 GND.n7546 163.367
R9077 GND.n7543 GND.n7542 163.367
R9078 GND.n7539 GND.n7538 163.367
R9079 GND.n7535 GND.n7534 163.367
R9080 GND.n7531 GND.n7530 163.367
R9081 GND.n7527 GND.n7526 163.367
R9082 GND.n7523 GND.n7522 163.367
R9083 GND.n7518 GND.n7517 163.367
R9084 GND.n7514 GND.n7513 163.367
R9085 GND.n7557 GND.n838 163.367
R9086 GND.n7439 GND.n7438 163.367
R9087 GND.n7443 GND.n7442 163.367
R9088 GND.n7447 GND.n7446 163.367
R9089 GND.n7451 GND.n7450 163.367
R9090 GND.n7455 GND.n7454 163.367
R9091 GND.n7459 GND.n7458 163.367
R9092 GND.n7463 GND.n7462 163.367
R9093 GND.n7467 GND.n7466 163.367
R9094 GND.n7471 GND.n7470 163.367
R9095 GND.n7475 GND.n7474 163.367
R9096 GND.n5486 GND.n1853 163.367
R9097 GND.n5490 GND.n1853 163.367
R9098 GND.n5495 GND.n5490 163.367
R9099 GND.n5496 GND.n5495 163.367
R9100 GND.n5496 GND.n5417 163.367
R9101 GND.n5499 GND.n5417 163.367
R9102 GND.n5499 GND.n5425 163.367
R9103 GND.n5502 GND.n5425 163.367
R9104 GND.n5502 GND.n5438 163.367
R9105 GND.n6169 GND.n5438 163.367
R9106 GND.n6169 GND.n5439 163.367
R9107 GND.n6165 GND.n5439 163.367
R9108 GND.n6165 GND.n5506 163.367
R9109 GND.n5517 GND.n5506 163.367
R9110 GND.n5593 GND.n5517 163.367
R9111 GND.n5598 GND.n5593 163.367
R9112 GND.n5599 GND.n5598 163.367
R9113 GND.n5599 GND.n5531 163.367
R9114 GND.n5602 GND.n5531 163.367
R9115 GND.n5602 GND.n5539 163.367
R9116 GND.n5606 GND.n5539 163.367
R9117 GND.n5611 GND.n5606 163.367
R9118 GND.n5612 GND.n5611 163.367
R9119 GND.n5612 GND.n5549 163.367
R9120 GND.n5615 GND.n5549 163.367
R9121 GND.n5615 GND.n5557 163.367
R9122 GND.n5619 GND.n5557 163.367
R9123 GND.n5624 GND.n5619 163.367
R9124 GND.n5625 GND.n5624 163.367
R9125 GND.n5625 GND.n5567 163.367
R9126 GND.n5628 GND.n5567 163.367
R9127 GND.n5628 GND.n5575 163.367
R9128 GND.n5631 GND.n5575 163.367
R9129 GND.n5631 GND.n5586 163.367
R9130 GND.n6108 GND.n5586 163.367
R9131 GND.n6108 GND.n5587 163.367
R9132 GND.n6104 GND.n5587 163.367
R9133 GND.n6104 GND.n5635 163.367
R9134 GND.n5649 GND.n5635 163.367
R9135 GND.n5726 GND.n5649 163.367
R9136 GND.n5731 GND.n5726 163.367
R9137 GND.n5732 GND.n5731 163.367
R9138 GND.n5732 GND.n5662 163.367
R9139 GND.n5735 GND.n5662 163.367
R9140 GND.n5735 GND.n5670 163.367
R9141 GND.n5739 GND.n5670 163.367
R9142 GND.n5744 GND.n5739 163.367
R9143 GND.n5745 GND.n5744 163.367
R9144 GND.n5745 GND.n5680 163.367
R9145 GND.n5748 GND.n5680 163.367
R9146 GND.n5748 GND.n5688 163.367
R9147 GND.n5752 GND.n5688 163.367
R9148 GND.n5757 GND.n5752 163.367
R9149 GND.n5758 GND.n5757 163.367
R9150 GND.n5758 GND.n5698 163.367
R9151 GND.n5761 GND.n5698 163.367
R9152 GND.n5761 GND.n5706 163.367
R9153 GND.n5764 GND.n5706 163.367
R9154 GND.n5764 GND.n5719 163.367
R9155 GND.n6047 GND.n5719 163.367
R9156 GND.n6047 GND.n5720 163.367
R9157 GND.n6043 GND.n5720 163.367
R9158 GND.n6043 GND.n5768 163.367
R9159 GND.n5780 GND.n5768 163.367
R9160 GND.n5856 GND.n5780 163.367
R9161 GND.n5861 GND.n5856 163.367
R9162 GND.n5862 GND.n5861 163.367
R9163 GND.n5862 GND.n5793 163.367
R9164 GND.n5865 GND.n5793 163.367
R9165 GND.n5865 GND.n5801 163.367
R9166 GND.n5869 GND.n5801 163.367
R9167 GND.n5875 GND.n5869 163.367
R9168 GND.n5876 GND.n5875 163.367
R9169 GND.n5876 GND.n5810 163.367
R9170 GND.n5879 GND.n5810 163.367
R9171 GND.n5879 GND.n5818 163.367
R9172 GND.n5883 GND.n5818 163.367
R9173 GND.n5888 GND.n5883 163.367
R9174 GND.n5889 GND.n5888 163.367
R9175 GND.n5889 GND.n5828 163.367
R9176 GND.n5892 GND.n5828 163.367
R9177 GND.n5892 GND.n5836 163.367
R9178 GND.n5895 GND.n5836 163.367
R9179 GND.n5895 GND.n5849 163.367
R9180 GND.n5986 GND.n5849 163.367
R9181 GND.n5986 GND.n5850 163.367
R9182 GND.n5982 GND.n5850 163.367
R9183 GND.n5982 GND.n5899 163.367
R9184 GND.n5911 GND.n5899 163.367
R9185 GND.n5936 GND.n5911 163.367
R9186 GND.n5941 GND.n5936 163.367
R9187 GND.n5942 GND.n5941 163.367
R9188 GND.n5942 GND.n5924 163.367
R9189 GND.n5945 GND.n5924 163.367
R9190 GND.n5945 GND.n5932 163.367
R9191 GND.n5949 GND.n5932 163.367
R9192 GND.n5949 GND.n1593 163.367
R9193 GND.n6422 GND.n1593 163.367
R9194 GND.n6422 GND.n1594 163.367
R9195 GND.n1594 GND.n1587 163.367
R9196 GND.n6417 GND.n1587 163.367
R9197 GND.n6417 GND.n1579 163.367
R9198 GND.n6412 GND.n1579 163.367
R9199 GND.n6412 GND.n1573 163.367
R9200 GND.n6409 GND.n1573 163.367
R9201 GND.n6409 GND.n1564 163.367
R9202 GND.n1607 GND.n1564 163.367
R9203 GND.n1607 GND.n1557 163.367
R9204 GND.n1604 GND.n1557 163.367
R9205 GND.n1604 GND.n1548 163.367
R9206 GND.n1601 GND.n1548 163.367
R9207 GND.n1601 GND.n1535 163.367
R9208 GND.n1597 GND.n1535 163.367
R9209 GND.n1597 GND.n1529 163.367
R9210 GND.n6505 GND.n1529 163.367
R9211 GND.n6505 GND.n1518 163.367
R9212 GND.n6511 GND.n1518 163.367
R9213 GND.n6512 GND.n6511 163.367
R9214 GND.n6512 GND.n1526 163.367
R9215 GND.n6517 GND.n1526 163.367
R9216 GND.n6517 GND.n1527 163.367
R9217 GND.n1527 GND.n1491 163.367
R9218 GND.n6579 GND.n1491 163.367
R9219 GND.n6579 GND.n1484 163.367
R9220 GND.n6575 GND.n1484 163.367
R9221 GND.n6575 GND.n1497 163.367
R9222 GND.n1497 GND.n1496 163.367
R9223 GND.n1496 GND.n1466 163.367
R9224 GND.n6621 GND.n1466 163.367
R9225 GND.n6621 GND.n1443 163.367
R9226 GND.n1463 GND.n1443 163.367
R9227 GND.n6627 GND.n1463 163.367
R9228 GND.n6627 GND.n1464 163.367
R9229 GND.n1464 GND.n1422 163.367
R9230 GND.n6684 GND.n1422 163.367
R9231 GND.n6684 GND.n1423 163.367
R9232 GND.n6680 GND.n1423 163.367
R9233 GND.n6680 GND.n6679 163.367
R9234 GND.n6679 GND.n1402 163.367
R9235 GND.n1403 GND.n1402 163.367
R9236 GND.n1403 GND.n1396 163.367
R9237 GND.n6673 GND.n1396 163.367
R9238 GND.n6673 GND.n1388 163.367
R9239 GND.n6669 GND.n1388 163.367
R9240 GND.n6669 GND.n1382 163.367
R9241 GND.n6666 GND.n1382 163.367
R9242 GND.n6666 GND.n1371 163.367
R9243 GND.n1371 GND.n1363 163.367
R9244 GND.n6781 GND.n1363 163.367
R9245 GND.n6781 GND.n1361 163.367
R9246 GND.n6788 GND.n1361 163.367
R9247 GND.n6788 GND.n1351 163.367
R9248 GND.n6784 GND.n1351 163.367
R9249 GND.n6784 GND.n1341 163.367
R9250 GND.n6842 GND.n1341 163.367
R9251 GND.n6842 GND.n1338 163.367
R9252 GND.n6847 GND.n1338 163.367
R9253 GND.n6847 GND.n1331 163.367
R9254 GND.n1331 GND.n1316 163.367
R9255 GND.n6879 GND.n1316 163.367
R9256 GND.n6879 GND.n1317 163.367
R9257 GND.n1317 GND.n1309 163.367
R9258 GND.n6874 GND.n1309 163.367
R9259 GND.n6874 GND.n1301 163.367
R9260 GND.n1301 GND.n1293 163.367
R9261 GND.n6918 GND.n1293 163.367
R9262 GND.n6918 GND.n1291 163.367
R9263 GND.n6923 GND.n1291 163.367
R9264 GND.n6923 GND.n1173 163.367
R9265 GND.n1173 GND.n1165 163.367
R9266 GND.n6992 GND.n1165 163.367
R9267 GND.n6992 GND.n1162 163.367
R9268 GND.n7001 GND.n1162 163.367
R9269 GND.n7001 GND.n1163 163.367
R9270 GND.n1163 GND.n1156 163.367
R9271 GND.n6996 GND.n1156 163.367
R9272 GND.n6996 GND.n1148 163.367
R9273 GND.n1148 GND.n1140 163.367
R9274 GND.n7034 GND.n1140 163.367
R9275 GND.n7034 GND.n1138 163.367
R9276 GND.n7038 GND.n1138 163.367
R9277 GND.n7038 GND.n1130 163.367
R9278 GND.n7049 GND.n1130 163.367
R9279 GND.n7049 GND.n1127 163.367
R9280 GND.n7055 GND.n1127 163.367
R9281 GND.n7055 GND.n1128 163.367
R9282 GND.n1128 GND.n1117 163.367
R9283 GND.n1117 GND.n1109 163.367
R9284 GND.n7083 GND.n1109 163.367
R9285 GND.n7083 GND.n1107 163.367
R9286 GND.n7087 GND.n1107 163.367
R9287 GND.n7087 GND.n1100 163.367
R9288 GND.n7096 GND.n1100 163.367
R9289 GND.n7096 GND.n1097 163.367
R9290 GND.n7105 GND.n1097 163.367
R9291 GND.n7105 GND.n1098 163.367
R9292 GND.n1098 GND.n1091 163.367
R9293 GND.n7100 GND.n1091 163.367
R9294 GND.n7100 GND.n1083 163.367
R9295 GND.n1083 GND.n1075 163.367
R9296 GND.n7132 GND.n1075 163.367
R9297 GND.n7132 GND.n1072 163.367
R9298 GND.n7141 GND.n1072 163.367
R9299 GND.n7141 GND.n1073 163.367
R9300 GND.n1073 GND.n1066 163.367
R9301 GND.n7136 GND.n1066 163.367
R9302 GND.n7136 GND.n1057 163.367
R9303 GND.n1057 GND.n1051 163.367
R9304 GND.n7170 GND.n1051 163.367
R9305 GND.n7170 GND.n1048 163.367
R9306 GND.n7179 GND.n1048 163.367
R9307 GND.n7179 GND.n1049 163.367
R9308 GND.n1049 GND.n1042 163.367
R9309 GND.n7174 GND.n1042 163.367
R9310 GND.n7174 GND.n1034 163.367
R9311 GND.n1034 GND.n1026 163.367
R9312 GND.n7215 GND.n1026 163.367
R9313 GND.n7215 GND.n1024 163.367
R9314 GND.n7219 GND.n1024 163.367
R9315 GND.n7219 GND.n1017 163.367
R9316 GND.n7228 GND.n1017 163.367
R9317 GND.n7228 GND.n1014 163.367
R9318 GND.n7237 GND.n1014 163.367
R9319 GND.n7237 GND.n1015 163.367
R9320 GND.n1015 GND.n1008 163.367
R9321 GND.n7232 GND.n1008 163.367
R9322 GND.n7232 GND.n1000 163.367
R9323 GND.n1000 GND.n992 163.367
R9324 GND.n7264 GND.n992 163.367
R9325 GND.n7264 GND.n989 163.367
R9326 GND.n7273 GND.n989 163.367
R9327 GND.n7273 GND.n990 163.367
R9328 GND.n990 GND.n983 163.367
R9329 GND.n7268 GND.n983 163.367
R9330 GND.n7268 GND.n975 163.367
R9331 GND.n975 GND.n967 163.367
R9332 GND.n7301 GND.n967 163.367
R9333 GND.n7301 GND.n964 163.367
R9334 GND.n7310 GND.n964 163.367
R9335 GND.n7310 GND.n965 163.367
R9336 GND.n965 GND.n958 163.367
R9337 GND.n7305 GND.n958 163.367
R9338 GND.n7305 GND.n950 163.367
R9339 GND.n950 GND.n942 163.367
R9340 GND.n7337 GND.n942 163.367
R9341 GND.n7337 GND.n939 163.367
R9342 GND.n7346 GND.n939 163.367
R9343 GND.n7346 GND.n940 163.367
R9344 GND.n940 GND.n933 163.367
R9345 GND.n7341 GND.n933 163.367
R9346 GND.n7341 GND.n925 163.367
R9347 GND.n925 GND.n918 163.367
R9348 GND.n7371 GND.n918 163.367
R9349 GND.n7371 GND.n916 163.367
R9350 GND.n7376 GND.n916 163.367
R9351 GND.n7376 GND.n908 163.367
R9352 GND.n908 GND.n902 163.367
R9353 GND.n7397 GND.n902 163.367
R9354 GND.n7397 GND.n899 163.367
R9355 GND.n7406 GND.n899 163.367
R9356 GND.n7406 GND.n900 163.367
R9357 GND.n900 GND.n893 163.367
R9358 GND.n7401 GND.n893 163.367
R9359 GND.n7401 GND.n885 163.367
R9360 GND.n885 GND.n878 163.367
R9361 GND.n7431 GND.n878 163.367
R9362 GND.n7431 GND.n876 163.367
R9363 GND.n7482 GND.n876 163.367
R9364 GND.n7482 GND.n867 163.367
R9365 GND.n868 GND.n867 163.367
R9366 GND.n1848 GND.n1847 163.367
R9367 GND.n6230 GND.n1847 163.367
R9368 GND.n6228 GND.n6227 163.367
R9369 GND.n6224 GND.n6223 163.367
R9370 GND.n6220 GND.n6219 163.367
R9371 GND.n6216 GND.n6215 163.367
R9372 GND.n6212 GND.n6211 163.367
R9373 GND.n6208 GND.n6207 163.367
R9374 GND.n6204 GND.n6203 163.367
R9375 GND.n6199 GND.n6198 163.367
R9376 GND.n6239 GND.n1823 163.367
R9377 GND.n5444 GND.n5443 163.367
R9378 GND.n5448 GND.n5447 163.367
R9379 GND.n5453 GND.n5452 163.367
R9380 GND.n5457 GND.n5456 163.367
R9381 GND.n5461 GND.n5460 163.367
R9382 GND.n5465 GND.n5464 163.367
R9383 GND.n5469 GND.n5468 163.367
R9384 GND.n5473 GND.n5472 163.367
R9385 GND.n5477 GND.n5476 163.367
R9386 GND.n5481 GND.n5480 163.367
R9387 GND.n5483 GND.n1845 163.367
R9388 GND.n6192 GND.n1849 163.367
R9389 GND.n6192 GND.n1851 163.367
R9390 GND.n5493 GND.n1851 163.367
R9391 GND.n5493 GND.n5419 163.367
R9392 GND.n6182 GND.n5419 163.367
R9393 GND.n6182 GND.n5420 163.367
R9394 GND.n6178 GND.n5420 163.367
R9395 GND.n6178 GND.n5423 163.367
R9396 GND.n5510 GND.n5423 163.367
R9397 GND.n5510 GND.n5436 163.367
R9398 GND.n5508 GND.n5436 163.367
R9399 GND.n6163 GND.n5508 163.367
R9400 GND.n6163 GND.n5509 163.367
R9401 GND.n6159 GND.n5509 163.367
R9402 GND.n6159 GND.n5515 163.367
R9403 GND.n5596 GND.n5515 163.367
R9404 GND.n5596 GND.n5533 163.367
R9405 GND.n6149 GND.n5533 163.367
R9406 GND.n6149 GND.n5534 163.367
R9407 GND.n6145 GND.n5534 163.367
R9408 GND.n6145 GND.n5537 163.367
R9409 GND.n5609 GND.n5537 163.367
R9410 GND.n5609 GND.n5551 163.367
R9411 GND.n6135 GND.n5551 163.367
R9412 GND.n6135 GND.n5552 163.367
R9413 GND.n6131 GND.n5552 163.367
R9414 GND.n6131 GND.n5555 163.367
R9415 GND.n5622 GND.n5555 163.367
R9416 GND.n5622 GND.n5569 163.367
R9417 GND.n6121 GND.n5569 163.367
R9418 GND.n6121 GND.n5570 163.367
R9419 GND.n6117 GND.n5570 163.367
R9420 GND.n6117 GND.n5573 163.367
R9421 GND.n5642 GND.n5573 163.367
R9422 GND.n5642 GND.n5584 163.367
R9423 GND.n5638 GND.n5584 163.367
R9424 GND.n6102 GND.n5638 163.367
R9425 GND.n6102 GND.n5639 163.367
R9426 GND.n6098 GND.n5639 163.367
R9427 GND.n6098 GND.n5647 163.367
R9428 GND.n5729 GND.n5647 163.367
R9429 GND.n5729 GND.n5664 163.367
R9430 GND.n6088 GND.n5664 163.367
R9431 GND.n6088 GND.n5665 163.367
R9432 GND.n6084 GND.n5665 163.367
R9433 GND.n6084 GND.n5668 163.367
R9434 GND.n5742 GND.n5668 163.367
R9435 GND.n5742 GND.n5682 163.367
R9436 GND.n6074 GND.n5682 163.367
R9437 GND.n6074 GND.n5683 163.367
R9438 GND.n6070 GND.n5683 163.367
R9439 GND.n6070 GND.n5686 163.367
R9440 GND.n5755 GND.n5686 163.367
R9441 GND.n5755 GND.n5700 163.367
R9442 GND.n6060 GND.n5700 163.367
R9443 GND.n6060 GND.n5701 163.367
R9444 GND.n6056 GND.n5701 163.367
R9445 GND.n6056 GND.n5704 163.367
R9446 GND.n5773 GND.n5704 163.367
R9447 GND.n5773 GND.n5717 163.367
R9448 GND.n5771 GND.n5717 163.367
R9449 GND.n6041 GND.n5771 163.367
R9450 GND.n6041 GND.n5772 163.367
R9451 GND.n6037 GND.n5772 163.367
R9452 GND.n6037 GND.n5778 163.367
R9453 GND.n5859 GND.n5778 163.367
R9454 GND.n5859 GND.n5795 163.367
R9455 GND.n6027 GND.n5795 163.367
R9456 GND.n6027 GND.n5796 163.367
R9457 GND.n6023 GND.n5796 163.367
R9458 GND.n6023 GND.n5799 163.367
R9459 GND.n5873 GND.n5799 163.367
R9460 GND.n5873 GND.n5812 163.367
R9461 GND.n6013 GND.n5812 163.367
R9462 GND.n6013 GND.n5813 163.367
R9463 GND.n6009 GND.n5813 163.367
R9464 GND.n6009 GND.n5816 163.367
R9465 GND.n5886 GND.n5816 163.367
R9466 GND.n5886 GND.n5830 163.367
R9467 GND.n5999 GND.n5830 163.367
R9468 GND.n5999 GND.n5831 163.367
R9469 GND.n5995 GND.n5831 163.367
R9470 GND.n5995 GND.n5834 163.367
R9471 GND.n5904 GND.n5834 163.367
R9472 GND.n5904 GND.n5847 163.367
R9473 GND.n5902 GND.n5847 163.367
R9474 GND.n5980 GND.n5902 163.367
R9475 GND.n5980 GND.n5903 163.367
R9476 GND.n5976 GND.n5903 163.367
R9477 GND.n5976 GND.n5909 163.367
R9478 GND.n5939 GND.n5909 163.367
R9479 GND.n5939 GND.n5926 163.367
R9480 GND.n5966 GND.n5926 163.367
R9481 GND.n5966 GND.n5927 163.367
R9482 GND.n5962 GND.n5927 163.367
R9483 GND.n5962 GND.n5930 163.367
R9484 GND.n5930 GND.n1591 163.367
R9485 GND.n6425 GND.n1591 163.367
R9486 GND.n6425 GND.n1589 163.367
R9487 GND.n6429 GND.n1589 163.367
R9488 GND.n6429 GND.n1577 163.367
R9489 GND.n6443 GND.n1577 163.367
R9490 GND.n6443 GND.n1575 163.367
R9491 GND.n6447 GND.n1575 163.367
R9492 GND.n6447 GND.n1562 163.367
R9493 GND.n6459 GND.n1562 163.367
R9494 GND.n6459 GND.n1559 163.367
R9495 GND.n6465 GND.n1559 163.367
R9496 GND.n6465 GND.n1560 163.367
R9497 GND.n1560 GND.n1546 163.367
R9498 GND.n1546 GND.n1533 163.367
R9499 GND.n6497 GND.n1533 163.367
R9500 GND.n6497 GND.n1531 163.367
R9501 GND.n6501 GND.n1531 163.367
R9502 GND.n6501 GND.n1520 163.367
R9503 GND.n6526 GND.n1520 163.367
R9504 GND.n6526 GND.n1521 163.367
R9505 GND.n6522 GND.n1521 163.367
R9506 GND.n6522 GND.n6521 163.367
R9507 GND.n6521 GND.n6520 163.367
R9508 GND.n6520 GND.n1489 163.367
R9509 GND.n6583 GND.n1489 163.367
R9510 GND.n6583 GND.n1486 163.367
R9511 GND.n6596 GND.n1486 163.367
R9512 GND.n6596 GND.n1487 163.367
R9513 GND.n6592 GND.n1487 163.367
R9514 GND.n6592 GND.n6591 163.367
R9515 GND.n6591 GND.n6590 163.367
R9516 GND.n6590 GND.n1445 163.367
R9517 GND.n6633 GND.n1445 163.367
R9518 GND.n6633 GND.n1446 163.367
R9519 GND.n6629 GND.n1446 163.367
R9520 GND.n6629 GND.n1460 163.367
R9521 GND.n1460 GND.n1459 163.367
R9522 GND.n1459 GND.n1420 163.367
R9523 GND.n1453 GND.n1420 163.367
R9524 GND.n1453 GND.n1450 163.367
R9525 GND.n1450 GND.n1400 163.367
R9526 GND.n6708 GND.n1400 163.367
R9527 GND.n6708 GND.n1398 163.367
R9528 GND.n6712 GND.n1398 163.367
R9529 GND.n6712 GND.n1386 163.367
R9530 GND.n6756 GND.n1386 163.367
R9531 GND.n6756 GND.n1384 163.367
R9532 GND.n6760 GND.n1384 163.367
R9533 GND.n6760 GND.n1369 163.367
R9534 GND.n6774 GND.n1369 163.367
R9535 GND.n6774 GND.n1366 163.367
R9536 GND.n6779 GND.n1366 163.367
R9537 GND.n6779 GND.n1367 163.367
R9538 GND.n1367 GND.n1352 163.367
R9539 GND.n6827 GND.n1352 163.367
R9540 GND.n6827 GND.n1353 163.367
R9541 GND.n6823 GND.n1353 163.367
R9542 GND.n6823 GND.n1336 163.367
R9543 GND.n6851 GND.n1336 163.367
R9544 GND.n6851 GND.n1334 163.367
R9545 GND.n6855 GND.n1334 163.367
R9546 GND.n6855 GND.n1313 163.367
R9547 GND.n6881 GND.n1313 163.367
R9548 GND.n6881 GND.n1311 163.367
R9549 GND.n6885 GND.n1311 163.367
R9550 GND.n6885 GND.n1300 163.367
R9551 GND.n6911 GND.n1300 163.367
R9552 GND.n6911 GND.n1296 163.367
R9553 GND.n6916 GND.n1296 163.367
R9554 GND.n6916 GND.n1298 163.367
R9555 GND.n1298 GND.n1171 163.367
R9556 GND.n6986 GND.n1171 163.367
R9557 GND.n6986 GND.n1169 163.367
R9558 GND.n6990 GND.n1169 163.367
R9559 GND.n6990 GND.n1160 163.367
R9560 GND.n7004 GND.n1160 163.367
R9561 GND.n7004 GND.n1158 163.367
R9562 GND.n7008 GND.n1158 163.367
R9563 GND.n7008 GND.n1146 163.367
R9564 GND.n7028 GND.n1146 163.367
R9565 GND.n7028 GND.n1144 163.367
R9566 GND.n7032 GND.n1144 163.367
R9567 GND.n7032 GND.n1136 163.367
R9568 GND.n7041 GND.n1136 163.367
R9569 GND.n7041 GND.n1133 163.367
R9570 GND.n7047 GND.n1133 163.367
R9571 GND.n7047 GND.n1134 163.367
R9572 GND.n1134 GND.n1125 163.367
R9573 GND.n1125 GND.n1115 163.367
R9574 GND.n7077 GND.n1115 163.367
R9575 GND.n7077 GND.n1113 163.367
R9576 GND.n7081 GND.n1113 163.367
R9577 GND.n7081 GND.n1105 163.367
R9578 GND.n7090 GND.n1105 163.367
R9579 GND.n7090 GND.n1103 163.367
R9580 GND.n7094 GND.n1103 163.367
R9581 GND.n7094 GND.n1095 163.367
R9582 GND.n7108 GND.n1095 163.367
R9583 GND.n7108 GND.n1093 163.367
R9584 GND.n7112 GND.n1093 163.367
R9585 GND.n7112 GND.n1081 163.367
R9586 GND.n7126 GND.n1081 163.367
R9587 GND.n7126 GND.n1079 163.367
R9588 GND.n7130 GND.n1079 163.367
R9589 GND.n7130 GND.n1070 163.367
R9590 GND.n7143 GND.n1070 163.367
R9591 GND.n7143 GND.n1068 163.367
R9592 GND.n7147 GND.n1068 163.367
R9593 GND.n7147 GND.n1055 163.367
R9594 GND.n7164 GND.n1055 163.367
R9595 GND.n7164 GND.n1053 163.367
R9596 GND.n7168 GND.n1053 163.367
R9597 GND.n7168 GND.n1046 163.367
R9598 GND.n7182 GND.n1046 163.367
R9599 GND.n7182 GND.n1044 163.367
R9600 GND.n7186 GND.n1044 163.367
R9601 GND.n7186 GND.n1032 163.367
R9602 GND.n7209 GND.n1032 163.367
R9603 GND.n7209 GND.n1030 163.367
R9604 GND.n7213 GND.n1030 163.367
R9605 GND.n7213 GND.n1022 163.367
R9606 GND.n7222 GND.n1022 163.367
R9607 GND.n7222 GND.n1020 163.367
R9608 GND.n7226 GND.n1020 163.367
R9609 GND.n7226 GND.n1012 163.367
R9610 GND.n7240 GND.n1012 163.367
R9611 GND.n7240 GND.n1010 163.367
R9612 GND.n7244 GND.n1010 163.367
R9613 GND.n7244 GND.n998 163.367
R9614 GND.n7258 GND.n998 163.367
R9615 GND.n7258 GND.n996 163.367
R9616 GND.n7262 GND.n996 163.367
R9617 GND.n7262 GND.n987 163.367
R9618 GND.n7275 GND.n987 163.367
R9619 GND.n7275 GND.n985 163.367
R9620 GND.n7279 GND.n985 163.367
R9621 GND.n7279 GND.n972 163.367
R9622 GND.n7295 GND.n972 163.367
R9623 GND.n7295 GND.n970 163.367
R9624 GND.n7299 GND.n970 163.367
R9625 GND.n7299 GND.n962 163.367
R9626 GND.n7313 GND.n962 163.367
R9627 GND.n7313 GND.n960 163.367
R9628 GND.n7317 GND.n960 163.367
R9629 GND.n7317 GND.n948 163.367
R9630 GND.n7331 GND.n948 163.367
R9631 GND.n7331 GND.n946 163.367
R9632 GND.n7335 GND.n946 163.367
R9633 GND.n7335 GND.n937 163.367
R9634 GND.n7348 GND.n937 163.367
R9635 GND.n7348 GND.n935 163.367
R9636 GND.n7352 GND.n935 163.367
R9637 GND.n7352 GND.n923 163.367
R9638 GND.n7364 GND.n923 163.367
R9639 GND.n7364 GND.n920 163.367
R9640 GND.n7369 GND.n920 163.367
R9641 GND.n7369 GND.n921 163.367
R9642 GND.n921 GND.n906 163.367
R9643 GND.n7391 GND.n906 163.367
R9644 GND.n7391 GND.n904 163.367
R9645 GND.n7395 GND.n904 163.367
R9646 GND.n7395 GND.n897 163.367
R9647 GND.n7408 GND.n897 163.367
R9648 GND.n7408 GND.n895 163.367
R9649 GND.n7412 GND.n895 163.367
R9650 GND.n7412 GND.n883 163.367
R9651 GND.n7424 GND.n883 163.367
R9652 GND.n7424 GND.n880 163.367
R9653 GND.n7429 GND.n880 163.367
R9654 GND.n7429 GND.n881 163.367
R9655 GND.n881 GND.n865 163.367
R9656 GND.n7508 GND.n865 163.367
R9657 GND.n7508 GND.n862 163.367
R9658 GND.n7558 GND.n837 143.351
R9659 GND.n6238 GND.n1821 143.351
R9660 GND.n1834 GND.n1821 143.351
R9661 GND.n30 GND.t87 141.24
R9662 GND.n30 GND.t9 140.468
R9663 GND.n7569 GND.n7568 123.734
R9664 GND.n7583 GND.n7582 123.734
R9665 GND.n430 GND.n429 123.734
R9666 GND.n2578 GND.n2577 110.933
R9667 GND.n1703 GND.n1702 110.933
R9668 GND.n1722 GND.n1721 110.933
R9669 GND.n1736 GND.n1735 110.933
R9670 GND.n1755 GND.n1754 110.933
R9671 GND.n1773 GND.n1772 110.933
R9672 GND.n817 GND.n816 110.933
R9673 GND.n831 GND.n830 110.933
R9674 GND.n7596 GND.n7595 110.933
R9675 GND.n443 GND.n442 110.933
R9676 GND.n419 GND.n418 110.933
R9677 GND.n406 GND.n405 110.933
R9678 GND.n395 GND.n394 110.933
R9679 GND.n8185 GND.n8184 110.933
R9680 GND.n1207 GND.n1206 110.933
R9681 GND.n2478 GND.n2477 110.933
R9682 GND.n2492 GND.n2491 110.933
R9683 GND.n2505 GND.n2504 110.933
R9684 GND.n2519 GND.n2518 110.933
R9685 GND.n2532 GND.n2531 110.933
R9686 GND.n1657 GND.n1656 110.933
R9687 GND.n7512 GND.n7511 105.115
R9688 GND.n6196 GND.n6195 105.115
R9689 GND.n5442 GND.n5441 105.115
R9690 GND.n7435 GND.n7434 105.115
R9691 GND.n6297 GND.t95 100.264
R9692 GND.n6939 GND.t131 100.264
R9693 GND.n8439 GND.n383 99.6594
R9694 GND.n8437 GND.n382 99.6594
R9695 GND.n8433 GND.n381 99.6594
R9696 GND.n8429 GND.n380 99.6594
R9697 GND.n8421 GND.n379 99.6594
R9698 GND.n8419 GND.n378 99.6594
R9699 GND.n8415 GND.n377 99.6594
R9700 GND.n8411 GND.n376 99.6594
R9701 GND.n8407 GND.n375 99.6594
R9702 GND.n408 GND.n374 99.6594
R9703 GND.n8399 GND.n373 99.6594
R9704 GND.n8395 GND.n372 99.6594
R9705 GND.n8391 GND.n371 99.6594
R9706 GND.n8387 GND.n370 99.6594
R9707 GND.n8383 GND.n369 99.6594
R9708 GND.n8375 GND.n368 99.6594
R9709 GND.n8373 GND.n367 99.6594
R9710 GND.n8369 GND.n366 99.6594
R9711 GND.n8365 GND.n365 99.6594
R9712 GND.n8361 GND.n364 99.6594
R9713 GND.n432 GND.n363 99.6594
R9714 GND.n8353 GND.n362 99.6594
R9715 GND.n8349 GND.n361 99.6594
R9716 GND.n8345 GND.n360 99.6594
R9717 GND.n8341 GND.n359 99.6594
R9718 GND.n8337 GND.n358 99.6594
R9719 GND.n8328 GND.n357 99.6594
R9720 GND.n7700 GND.n7699 99.6594
R9721 GND.n7694 GND.n680 99.6594
R9722 GND.n7691 GND.n681 99.6594
R9723 GND.n7687 GND.n682 99.6594
R9724 GND.n7683 GND.n683 99.6594
R9725 GND.n7679 GND.n684 99.6594
R9726 GND.n7675 GND.n685 99.6594
R9727 GND.n7671 GND.n686 99.6594
R9728 GND.n7667 GND.n687 99.6594
R9729 GND.n7663 GND.n688 99.6594
R9730 GND.n7659 GND.n689 99.6594
R9731 GND.n7656 GND.n690 99.6594
R9732 GND.n7651 GND.n692 99.6594
R9733 GND.n7647 GND.n693 99.6594
R9734 GND.n7643 GND.n694 99.6594
R9735 GND.n7639 GND.n695 99.6594
R9736 GND.n7635 GND.n696 99.6594
R9737 GND.n7631 GND.n697 99.6594
R9738 GND.n7627 GND.n698 99.6594
R9739 GND.n7623 GND.n699 99.6594
R9740 GND.n7619 GND.n700 99.6594
R9741 GND.n7616 GND.n701 99.6594
R9742 GND.n7612 GND.n702 99.6594
R9743 GND.n7608 GND.n703 99.6594
R9744 GND.n7604 GND.n704 99.6594
R9745 GND.n7600 GND.n705 99.6594
R9746 GND.n1693 GND.n1688 99.6594
R9747 GND.n1695 GND.n1687 99.6594
R9748 GND.n1699 GND.n1686 99.6594
R9749 GND.n1701 GND.n1685 99.6594
R9750 GND.n1707 GND.n1684 99.6594
R9751 GND.n1709 GND.n1683 99.6594
R9752 GND.n1713 GND.n1682 99.6594
R9753 GND.n1715 GND.n1681 99.6594
R9754 GND.n1719 GND.n1680 99.6594
R9755 GND.n1724 GND.n1679 99.6594
R9756 GND.n6243 GND.n1678 99.6594
R9757 GND.n1728 GND.n1676 99.6594
R9758 GND.n1732 GND.n1675 99.6594
R9759 GND.n1734 GND.n1674 99.6594
R9760 GND.n1740 GND.n1673 99.6594
R9761 GND.n1742 GND.n1672 99.6594
R9762 GND.n1746 GND.n1671 99.6594
R9763 GND.n1748 GND.n1670 99.6594
R9764 GND.n1752 GND.n1669 99.6594
R9765 GND.n1757 GND.n1668 99.6594
R9766 GND.n1761 GND.n1667 99.6594
R9767 GND.n1763 GND.n1666 99.6594
R9768 GND.n1767 GND.n1665 99.6594
R9769 GND.n1769 GND.n1664 99.6594
R9770 GND.n1774 GND.n1663 99.6594
R9771 GND.n1662 GND.n1629 99.6594
R9772 GND.n2974 GND.n2973 99.6594
R9773 GND.n2968 GND.n2431 99.6594
R9774 GND.n2965 GND.n2432 99.6594
R9775 GND.n2961 GND.n2433 99.6594
R9776 GND.n2957 GND.n2434 99.6594
R9777 GND.n2953 GND.n2435 99.6594
R9778 GND.n2949 GND.n2436 99.6594
R9779 GND.n2945 GND.n2437 99.6594
R9780 GND.n2941 GND.n2438 99.6594
R9781 GND.n2937 GND.n2439 99.6594
R9782 GND.n2933 GND.n2440 99.6594
R9783 GND.n2930 GND.n2441 99.6594
R9784 GND.n2926 GND.n2442 99.6594
R9785 GND.n2922 GND.n2443 99.6594
R9786 GND.n2918 GND.n2444 99.6594
R9787 GND.n2914 GND.n2445 99.6594
R9788 GND.n2910 GND.n2446 99.6594
R9789 GND.n2906 GND.n2447 99.6594
R9790 GND.n2902 GND.n2448 99.6594
R9791 GND.n2898 GND.n2449 99.6594
R9792 GND.n2894 GND.n2450 99.6594
R9793 GND.n2890 GND.n2451 99.6594
R9794 GND.n2887 GND.n2452 99.6594
R9795 GND.n2883 GND.n2453 99.6594
R9796 GND.n2879 GND.n2454 99.6594
R9797 GND.n2875 GND.n2455 99.6594
R9798 GND.n2871 GND.n2456 99.6594
R9799 GND.n6976 GND.n6975 99.6594
R9800 GND.n6973 GND.n6972 99.6594
R9801 GND.n6968 GND.n1190 99.6594
R9802 GND.n6966 GND.n6965 99.6594
R9803 GND.n6961 GND.n1197 99.6594
R9804 GND.n6959 GND.n6958 99.6594
R9805 GND.n6954 GND.n1277 99.6594
R9806 GND.n6952 GND.n6951 99.6594
R9807 GND.n6946 GND.n1281 99.6594
R9808 GND.n6944 GND.n6943 99.6594
R9809 GND.n6935 GND.n1285 99.6594
R9810 GND.n6933 GND.n6932 99.6594
R9811 GND.n6316 GND.n6315 99.6594
R9812 GND.n6324 GND.n6323 99.6594
R9813 GND.n6327 GND.n6326 99.6594
R9814 GND.n6335 GND.n6334 99.6594
R9815 GND.n6338 GND.n6337 99.6594
R9816 GND.n6343 GND.n6342 99.6594
R9817 GND.n6348 GND.n6347 99.6594
R9818 GND.n6353 GND.n6352 99.6594
R9819 GND.n6358 GND.n6357 99.6594
R9820 GND.n6363 GND.n6362 99.6594
R9821 GND.n6366 GND.n6365 99.6594
R9822 GND.n6374 GND.n6373 99.6594
R9823 GND.n8196 GND.n352 99.6594
R9824 GND.n8200 GND.n353 99.6594
R9825 GND.n8206 GND.n354 99.6594
R9826 GND.n8210 GND.n355 99.6594
R9827 GND.n8216 GND.n356 99.6594
R9828 GND.n1225 GND.n706 99.6594
R9829 GND.n1222 GND.n707 99.6594
R9830 GND.n1218 GND.n708 99.6594
R9831 GND.n1214 GND.n709 99.6594
R9832 GND.n1210 GND.n710 99.6594
R9833 GND.n4730 GND.n4729 99.6594
R9834 GND.n4733 GND.n4732 99.6594
R9835 GND.n4740 GND.n4739 99.6594
R9836 GND.n4743 GND.n4742 99.6594
R9837 GND.n4750 GND.n4749 99.6594
R9838 GND.n4753 GND.n4752 99.6594
R9839 GND.n4760 GND.n4759 99.6594
R9840 GND.n4763 GND.n4762 99.6594
R9841 GND.n4770 GND.n4769 99.6594
R9842 GND.n4773 GND.n4772 99.6594
R9843 GND.n4780 GND.n4779 99.6594
R9844 GND.n4783 GND.n4782 99.6594
R9845 GND.n4790 GND.n4789 99.6594
R9846 GND.n4793 GND.n4792 99.6594
R9847 GND.n4800 GND.n4799 99.6594
R9848 GND.n4803 GND.n4802 99.6594
R9849 GND.n4810 GND.n4809 99.6594
R9850 GND.n4813 GND.n4812 99.6594
R9851 GND.n4820 GND.n4819 99.6594
R9852 GND.n4823 GND.n4822 99.6594
R9853 GND.n4830 GND.n4829 99.6594
R9854 GND.n4833 GND.n4832 99.6594
R9855 GND.n4841 GND.n4840 99.6594
R9856 GND.n4844 GND.n4843 99.6594
R9857 GND.n4731 GND.n4730 99.6594
R9858 GND.n4732 GND.n3018 99.6594
R9859 GND.n4741 GND.n4740 99.6594
R9860 GND.n4742 GND.n3014 99.6594
R9861 GND.n4751 GND.n4750 99.6594
R9862 GND.n4752 GND.n3010 99.6594
R9863 GND.n4761 GND.n4760 99.6594
R9864 GND.n4762 GND.n3006 99.6594
R9865 GND.n4771 GND.n4770 99.6594
R9866 GND.n4772 GND.n3002 99.6594
R9867 GND.n4781 GND.n4780 99.6594
R9868 GND.n4782 GND.n2998 99.6594
R9869 GND.n4791 GND.n4790 99.6594
R9870 GND.n4792 GND.n2994 99.6594
R9871 GND.n4801 GND.n4800 99.6594
R9872 GND.n4802 GND.n2990 99.6594
R9873 GND.n4811 GND.n4810 99.6594
R9874 GND.n4812 GND.n2986 99.6594
R9875 GND.n4821 GND.n4820 99.6594
R9876 GND.n4822 GND.n2982 99.6594
R9877 GND.n4831 GND.n4830 99.6594
R9878 GND.n4832 GND.n2978 99.6594
R9879 GND.n4842 GND.n4841 99.6594
R9880 GND.n4845 GND.n4844 99.6594
R9881 GND.n1223 GND.n706 99.6594
R9882 GND.n1219 GND.n707 99.6594
R9883 GND.n1215 GND.n708 99.6594
R9884 GND.n1211 GND.n709 99.6594
R9885 GND.n1205 GND.n710 99.6594
R9886 GND.n8209 GND.n356 99.6594
R9887 GND.n8207 GND.n355 99.6594
R9888 GND.n8199 GND.n354 99.6594
R9889 GND.n8197 GND.n353 99.6594
R9890 GND.n8191 GND.n352 99.6594
R9891 GND.n6317 GND.n6316 99.6594
R9892 GND.n6325 GND.n6324 99.6594
R9893 GND.n6326 GND.n6304 99.6594
R9894 GND.n6336 GND.n6335 99.6594
R9895 GND.n6337 GND.n6301 99.6594
R9896 GND.n6344 GND.n6343 99.6594
R9897 GND.n6349 GND.n6348 99.6594
R9898 GND.n6354 GND.n6353 99.6594
R9899 GND.n6359 GND.n6358 99.6594
R9900 GND.n6364 GND.n6363 99.6594
R9901 GND.n6365 GND.n1614 99.6594
R9902 GND.n6375 GND.n6374 99.6594
R9903 GND.n6934 GND.n6933 99.6594
R9904 GND.n1285 GND.n1283 99.6594
R9905 GND.n6945 GND.n6944 99.6594
R9906 GND.n1281 GND.n1279 99.6594
R9907 GND.n6953 GND.n6952 99.6594
R9908 GND.n1277 GND.n1198 99.6594
R9909 GND.n6960 GND.n6959 99.6594
R9910 GND.n1197 GND.n1191 99.6594
R9911 GND.n6967 GND.n6966 99.6594
R9912 GND.n1190 GND.n1183 99.6594
R9913 GND.n6974 GND.n6973 99.6594
R9914 GND.n6977 GND.n6976 99.6594
R9915 GND.n2974 GND.n2465 99.6594
R9916 GND.n2966 GND.n2431 99.6594
R9917 GND.n2962 GND.n2432 99.6594
R9918 GND.n2958 GND.n2433 99.6594
R9919 GND.n2954 GND.n2434 99.6594
R9920 GND.n2950 GND.n2435 99.6594
R9921 GND.n2946 GND.n2436 99.6594
R9922 GND.n2942 GND.n2437 99.6594
R9923 GND.n2938 GND.n2438 99.6594
R9924 GND.n2489 GND.n2439 99.6594
R9925 GND.n2931 GND.n2440 99.6594
R9926 GND.n2927 GND.n2441 99.6594
R9927 GND.n2923 GND.n2442 99.6594
R9928 GND.n2919 GND.n2443 99.6594
R9929 GND.n2915 GND.n2444 99.6594
R9930 GND.n2911 GND.n2445 99.6594
R9931 GND.n2907 GND.n2446 99.6594
R9932 GND.n2903 GND.n2447 99.6594
R9933 GND.n2899 GND.n2448 99.6594
R9934 GND.n2895 GND.n2449 99.6594
R9935 GND.n2516 GND.n2450 99.6594
R9936 GND.n2888 GND.n2451 99.6594
R9937 GND.n2884 GND.n2452 99.6594
R9938 GND.n2880 GND.n2453 99.6594
R9939 GND.n2876 GND.n2454 99.6594
R9940 GND.n2872 GND.n2455 99.6594
R9941 GND.n2540 GND.n2456 99.6594
R9942 GND.n1775 GND.n1662 99.6594
R9943 GND.n1770 GND.n1663 99.6594
R9944 GND.n1768 GND.n1664 99.6594
R9945 GND.n1764 GND.n1665 99.6594
R9946 GND.n1762 GND.n1666 99.6594
R9947 GND.n1758 GND.n1667 99.6594
R9948 GND.n1753 GND.n1668 99.6594
R9949 GND.n1749 GND.n1669 99.6594
R9950 GND.n1747 GND.n1670 99.6594
R9951 GND.n1743 GND.n1671 99.6594
R9952 GND.n1741 GND.n1672 99.6594
R9953 GND.n1737 GND.n1673 99.6594
R9954 GND.n1733 GND.n1674 99.6594
R9955 GND.n1729 GND.n1675 99.6594
R9956 GND.n6244 GND.n1677 99.6594
R9957 GND.n1725 GND.n1678 99.6594
R9958 GND.n1720 GND.n1679 99.6594
R9959 GND.n1716 GND.n1680 99.6594
R9960 GND.n1714 GND.n1681 99.6594
R9961 GND.n1710 GND.n1682 99.6594
R9962 GND.n1708 GND.n1683 99.6594
R9963 GND.n1704 GND.n1684 99.6594
R9964 GND.n1700 GND.n1685 99.6594
R9965 GND.n1696 GND.n1686 99.6594
R9966 GND.n1694 GND.n1687 99.6594
R9967 GND.n1689 GND.n1688 99.6594
R9968 GND.n7700 GND.n713 99.6594
R9969 GND.n7692 GND.n680 99.6594
R9970 GND.n7688 GND.n681 99.6594
R9971 GND.n7684 GND.n682 99.6594
R9972 GND.n7680 GND.n683 99.6594
R9973 GND.n7676 GND.n684 99.6594
R9974 GND.n7672 GND.n685 99.6594
R9975 GND.n7668 GND.n686 99.6594
R9976 GND.n7664 GND.n687 99.6594
R9977 GND.n828 GND.n688 99.6594
R9978 GND.n7657 GND.n689 99.6594
R9979 GND.n7652 GND.n691 99.6594
R9980 GND.n7648 GND.n692 99.6594
R9981 GND.n7644 GND.n693 99.6594
R9982 GND.n7640 GND.n694 99.6594
R9983 GND.n7636 GND.n695 99.6594
R9984 GND.n7632 GND.n696 99.6594
R9985 GND.n7628 GND.n697 99.6594
R9986 GND.n7624 GND.n698 99.6594
R9987 GND.n7580 GND.n699 99.6594
R9988 GND.n7617 GND.n700 99.6594
R9989 GND.n7613 GND.n701 99.6594
R9990 GND.n7609 GND.n702 99.6594
R9991 GND.n7605 GND.n703 99.6594
R9992 GND.n7601 GND.n704 99.6594
R9993 GND.n705 GND.n669 99.6594
R9994 GND.n8336 GND.n357 99.6594
R9995 GND.n8340 GND.n358 99.6594
R9996 GND.n8344 GND.n359 99.6594
R9997 GND.n8348 GND.n360 99.6594
R9998 GND.n8352 GND.n361 99.6594
R9999 GND.n431 GND.n362 99.6594
R10000 GND.n8360 GND.n363 99.6594
R10001 GND.n8364 GND.n364 99.6594
R10002 GND.n8368 GND.n365 99.6594
R10003 GND.n8372 GND.n366 99.6594
R10004 GND.n8376 GND.n367 99.6594
R10005 GND.n8382 GND.n368 99.6594
R10006 GND.n8386 GND.n369 99.6594
R10007 GND.n8390 GND.n370 99.6594
R10008 GND.n8394 GND.n371 99.6594
R10009 GND.n8398 GND.n372 99.6594
R10010 GND.n407 GND.n373 99.6594
R10011 GND.n8406 GND.n374 99.6594
R10012 GND.n8410 GND.n375 99.6594
R10013 GND.n8414 GND.n376 99.6594
R10014 GND.n8418 GND.n377 99.6594
R10015 GND.n8422 GND.n378 99.6594
R10016 GND.n8428 GND.n379 99.6594
R10017 GND.n8432 GND.n380 99.6594
R10018 GND.n8436 GND.n381 99.6594
R10019 GND.n8440 GND.n382 99.6594
R10020 GND.n385 GND.n383 99.6594
R10021 GND.n2864 GND.n2457 99.6594
R10022 GND.n2587 GND.n2458 99.6594
R10023 GND.n2585 GND.n2459 99.6594
R10024 GND.n2595 GND.n2460 99.6594
R10025 GND.n2581 GND.n2461 99.6594
R10026 GND.n2586 GND.n2457 99.6594
R10027 GND.n2584 GND.n2458 99.6594
R10028 GND.n2594 GND.n2459 99.6594
R10029 GND.n2580 GND.n2460 99.6594
R10030 GND.n2576 GND.n2461 99.6594
R10031 GND.n6284 GND.n6283 99.6594
R10032 GND.n1641 GND.n1640 99.6594
R10033 GND.n1646 GND.n1645 99.6594
R10034 GND.n1651 GND.n1650 99.6594
R10035 GND.n1655 GND.n1654 99.6594
R10036 GND.n1659 GND.n1655 99.6594
R10037 GND.n1653 GND.n1651 99.6594
R10038 GND.n1647 GND.n1646 99.6594
R10039 GND.n1642 GND.n1641 99.6594
R10040 GND.n6283 GND.n1636 99.6594
R10041 GND.n5 GND.t59 88.2828
R10042 GND.n9 GND.t54 88.2828
R10043 GND.n14 GND.t55 88.2828
R10044 GND.n19 GND.t72 88.2828
R10045 GND.n24 GND.t33 88.2828
R10046 GND.n1 GND.t58 88.2828
R10047 GND.n36 GND.t48 86.4495
R10048 GND.n40 GND.t47 86.4495
R10049 GND.n45 GND.t46 86.4495
R10050 GND.n50 GND.t43 86.4495
R10051 GND.n55 GND.t22 86.4495
R10052 GND.n60 GND.t51 86.4495
R10053 GND.n2578 GND.t90 78.4142
R10054 GND.n1703 GND.t145 78.4142
R10055 GND.n1722 GND.t139 78.4142
R10056 GND.n1736 GND.t142 78.4142
R10057 GND.n1755 GND.t155 78.4142
R10058 GND.n1773 GND.t128 78.4142
R10059 GND.n817 GND.t169 78.4142
R10060 GND.n831 GND.t166 78.4142
R10061 GND.n7596 GND.t175 78.4142
R10062 GND.n443 GND.t112 78.4142
R10063 GND.n419 GND.t118 78.4142
R10064 GND.n406 GND.t121 78.4142
R10065 GND.n395 GND.t124 78.4142
R10066 GND.n8185 GND.t161 78.4142
R10067 GND.n1207 GND.t135 78.4142
R10068 GND.n2478 GND.t103 78.4142
R10069 GND.n2492 GND.t100 78.4142
R10070 GND.n2505 GND.t97 78.4142
R10071 GND.n2519 GND.t181 78.4142
R10072 GND.n2532 GND.t151 78.4142
R10073 GND.n1657 GND.t173 78.4142
R10074 GND.n7569 GND.t163 75.2142
R10075 GND.n7583 GND.t157 75.2142
R10076 GND.n430 GND.t185 75.2142
R10077 GND.n31 GND.t187 73.7497
R10078 GND.n31 GND.t83 72.9764
R10079 GND.n7551 GND.n861 71.676
R10080 GND.n7547 GND.n860 71.676
R10081 GND.n7543 GND.n859 71.676
R10082 GND.n7539 GND.n858 71.676
R10083 GND.n7535 GND.n857 71.676
R10084 GND.n7531 GND.n856 71.676
R10085 GND.n7527 GND.n855 71.676
R10086 GND.n7523 GND.n854 71.676
R10087 GND.n7518 GND.n853 71.676
R10088 GND.n7514 GND.n852 71.676
R10089 GND.n7558 GND.n7557 71.676
R10090 GND.n7438 GND.n840 71.676
R10091 GND.n7442 GND.n841 71.676
R10092 GND.n7446 GND.n842 71.676
R10093 GND.n7450 GND.n843 71.676
R10094 GND.n7454 GND.n844 71.676
R10095 GND.n7458 GND.n845 71.676
R10096 GND.n7462 GND.n846 71.676
R10097 GND.n7466 GND.n847 71.676
R10098 GND.n7470 GND.n848 71.676
R10099 GND.n7474 GND.n849 71.676
R10100 GND.n7477 GND.n850 71.676
R10101 GND.n6236 GND.n6235 71.676
R10102 GND.n6230 GND.n1825 71.676
R10103 GND.n6227 GND.n1826 71.676
R10104 GND.n6223 GND.n1827 71.676
R10105 GND.n6219 GND.n1828 71.676
R10106 GND.n6215 GND.n1829 71.676
R10107 GND.n6211 GND.n1830 71.676
R10108 GND.n6207 GND.n1831 71.676
R10109 GND.n6203 GND.n1832 71.676
R10110 GND.n6198 GND.n1833 71.676
R10111 GND.n6239 GND.n6238 71.676
R10112 GND.n5444 GND.n1835 71.676
R10113 GND.n5448 GND.n1836 71.676
R10114 GND.n5453 GND.n1837 71.676
R10115 GND.n5457 GND.n1838 71.676
R10116 GND.n5461 GND.n1839 71.676
R10117 GND.n5465 GND.n1840 71.676
R10118 GND.n5469 GND.n1841 71.676
R10119 GND.n5473 GND.n1842 71.676
R10120 GND.n5477 GND.n1843 71.676
R10121 GND.n5481 GND.n1844 71.676
R10122 GND.n6236 GND.n1848 71.676
R10123 GND.n6228 GND.n1825 71.676
R10124 GND.n6224 GND.n1826 71.676
R10125 GND.n6220 GND.n1827 71.676
R10126 GND.n6216 GND.n1828 71.676
R10127 GND.n6212 GND.n1829 71.676
R10128 GND.n6208 GND.n1830 71.676
R10129 GND.n6204 GND.n1831 71.676
R10130 GND.n6199 GND.n1832 71.676
R10131 GND.n1833 GND.n1823 71.676
R10132 GND.n5443 GND.n1834 71.676
R10133 GND.n5447 GND.n1835 71.676
R10134 GND.n5452 GND.n1836 71.676
R10135 GND.n5456 GND.n1837 71.676
R10136 GND.n5460 GND.n1838 71.676
R10137 GND.n5464 GND.n1839 71.676
R10138 GND.n5468 GND.n1840 71.676
R10139 GND.n5472 GND.n1841 71.676
R10140 GND.n5476 GND.n1842 71.676
R10141 GND.n5480 GND.n1843 71.676
R10142 GND.n5483 GND.n1844 71.676
R10143 GND.n7475 GND.n850 71.676
R10144 GND.n7471 GND.n849 71.676
R10145 GND.n7467 GND.n848 71.676
R10146 GND.n7463 GND.n847 71.676
R10147 GND.n7459 GND.n846 71.676
R10148 GND.n7455 GND.n845 71.676
R10149 GND.n7451 GND.n844 71.676
R10150 GND.n7447 GND.n843 71.676
R10151 GND.n7443 GND.n842 71.676
R10152 GND.n7439 GND.n841 71.676
R10153 GND.n840 GND.n838 71.676
R10154 GND.n7513 GND.n837 71.676
R10155 GND.n7517 GND.n852 71.676
R10156 GND.n7522 GND.n853 71.676
R10157 GND.n7526 GND.n854 71.676
R10158 GND.n7530 GND.n855 71.676
R10159 GND.n7534 GND.n856 71.676
R10160 GND.n7538 GND.n857 71.676
R10161 GND.n7542 GND.n858 71.676
R10162 GND.n7546 GND.n859 71.676
R10163 GND.n7550 GND.n860 71.676
R10164 GND.n863 GND.n861 71.676
R10165 GND.n2975 GND.n2463 71.0366
R10166 GND.n8448 GND.n350 71.0366
R10167 GND.n35 GND.n33 69.2446
R10168 GND.n39 GND.n37 69.2446
R10169 GND.n44 GND.n42 69.2446
R10170 GND.n49 GND.n47 69.2446
R10171 GND.n54 GND.n52 69.2446
R10172 GND.n59 GND.n57 69.2446
R10173 GND.n5 GND.n4 67.4112
R10174 GND.n7 GND.n6 67.4112
R10175 GND.n9 GND.n8 67.4112
R10176 GND.n11 GND.n10 67.4112
R10177 GND.n14 GND.n13 67.4112
R10178 GND.n16 GND.n15 67.4112
R10179 GND.n19 GND.n18 67.4112
R10180 GND.n21 GND.n20 67.4112
R10181 GND.n24 GND.n23 67.4112
R10182 GND.n26 GND.n25 67.4112
R10183 GND.n1 GND.n0 67.4112
R10184 GND.n3 GND.n2 67.4112
R10185 GND.n35 GND.n34 67.4112
R10186 GND.n39 GND.n38 67.4112
R10187 GND.n44 GND.n43 67.4112
R10188 GND.n49 GND.n48 67.4112
R10189 GND.n54 GND.n53 67.4112
R10190 GND.n59 GND.n58 67.4112
R10191 GND.n5442 GND.t148 67.2784
R10192 GND.n7435 GND.t115 67.2784
R10193 GND.n7512 GND.t108 67.2767
R10194 GND.n6196 GND.t178 67.2767
R10195 GND.n6298 GND.t94 61.0883
R10196 GND.n6940 GND.t132 61.0883
R10197 GND.n7520 GND.n7512 53.1399
R10198 GND.n6201 GND.n6196 53.1399
R10199 GND.n5450 GND.n5442 53.1399
R10200 GND.n7436 GND.n7435 53.1399
R10201 GND.n7642 GND.n7569 48.6793
R10202 GND.n7621 GND.n7583 48.6793
R10203 GND.n8358 GND.n430 48.6793
R10204 GND.n6298 GND.n6297 39.1763
R10205 GND.n6940 GND.n6939 39.1763
R10206 GND.n2601 GND.n2578 35.8793
R10207 GND.n1705 GND.n1703 35.8793
R10208 GND.n6250 GND.n1722 35.8793
R10209 GND.n1738 GND.n1736 35.8793
R10210 GND.n1794 GND.n1755 35.8793
R10211 GND.n1777 GND.n1773 35.8793
R10212 GND.n7682 GND.n817 35.8793
R10213 GND.n7661 GND.n831 35.8793
R10214 GND.n7599 GND.n7596 35.8793
R10215 GND.n8335 GND.n443 35.8793
R10216 GND.n8381 GND.n419 35.8793
R10217 GND.n8404 GND.n406 35.8793
R10218 GND.n8427 GND.n395 35.8793
R10219 GND.n8186 GND.n8185 35.8793
R10220 GND.n6299 GND.n6298 35.8793
R10221 GND.n6941 GND.n6940 35.8793
R10222 GND.n1208 GND.n1207 35.8793
R10223 GND.n2956 GND.n2478 35.8793
R10224 GND.n2935 GND.n2492 35.8793
R10225 GND.n2913 GND.n2505 35.8793
R10226 GND.n2892 GND.n2519 35.8793
R10227 GND.n2870 GND.n2532 35.8793
R10228 GND.n1658 GND.n1657 35.8793
R10229 GND.n7479 GND.n7478 35.7468
R10230 GND.n7554 GND.n7510 35.7468
R10231 GND.n5487 GND.n5485 35.7468
R10232 GND.n6234 GND.n6194 35.7468
R10233 GND.n2572 GND.n2463 35.3419
R10234 GND.n2613 GND.n2572 35.3419
R10235 GND.n2613 GND.n2560 35.3419
R10236 GND.n2716 GND.n2560 35.3419
R10237 GND.n2716 GND.n2552 35.3419
R10238 GND.n2848 GND.n2552 35.3419
R10239 GND.n4852 GND.n2413 35.3419
R10240 GND.n4864 GND.n2413 35.3419
R10241 GND.n4864 GND.n2404 35.3419
R10242 GND.n4872 GND.n2404 35.3419
R10243 GND.n4872 GND.n2393 35.3419
R10244 GND.n4884 GND.n2393 35.3419
R10245 GND.n4884 GND.n2384 35.3419
R10246 GND.n4892 GND.n2384 35.3419
R10247 GND.n4892 GND.n2373 35.3419
R10248 GND.n4904 GND.n2373 35.3419
R10249 GND.n4904 GND.n2364 35.3419
R10250 GND.n4912 GND.n2364 35.3419
R10251 GND.n4912 GND.n2352 35.3419
R10252 GND.n4924 GND.n2352 35.3419
R10253 GND.n4924 GND.n2355 35.3419
R10254 GND.n4932 GND.n2333 35.3419
R10255 GND.n4944 GND.n2333 35.3419
R10256 GND.n4944 GND.n2324 35.3419
R10257 GND.n4952 GND.n2324 35.3419
R10258 GND.n4952 GND.n2313 35.3419
R10259 GND.n4964 GND.n2313 35.3419
R10260 GND.n4964 GND.n2304 35.3419
R10261 GND.n4972 GND.n2304 35.3419
R10262 GND.n4972 GND.n2293 35.3419
R10263 GND.n4984 GND.n2293 35.3419
R10264 GND.n4984 GND.n2284 35.3419
R10265 GND.n4992 GND.n2284 35.3419
R10266 GND.n5004 GND.n2273 35.3419
R10267 GND.n5004 GND.n2264 35.3419
R10268 GND.n5013 GND.n2264 35.3419
R10269 GND.n5013 GND.n2252 35.3419
R10270 GND.n5030 GND.n2252 35.3419
R10271 GND.n5030 GND.n2255 35.3419
R10272 GND.n2255 GND.n2241 35.3419
R10273 GND.n5038 GND.n2241 35.3419
R10274 GND.n5038 GND.n2227 35.3419
R10275 GND.n5050 GND.n2227 35.3419
R10276 GND.n5050 GND.n2218 35.3419
R10277 GND.t34 GND.n2218 35.3419
R10278 GND.t34 GND.n2205 35.3419
R10279 GND.n5075 GND.n2205 35.3419
R10280 GND.n5075 GND.n2198 35.3419
R10281 GND.n5081 GND.n2198 35.3419
R10282 GND.n5081 GND.n2072 35.3419
R10283 GND.n5090 GND.n2072 35.3419
R10284 GND.n5090 GND.n2061 35.3419
R10285 GND.n5107 GND.n2061 35.3419
R10286 GND.n5107 GND.n2051 35.3419
R10287 GND.n5117 GND.n2051 35.3419
R10288 GND.n5117 GND.n2044 35.3419
R10289 GND.n5187 GND.n2044 35.3419
R10290 GND.n5198 GND.n2025 35.3419
R10291 GND.n5206 GND.n2025 35.3419
R10292 GND.n5206 GND.n2014 35.3419
R10293 GND.n5218 GND.n2014 35.3419
R10294 GND.n5218 GND.n2005 35.3419
R10295 GND.n5226 GND.n2005 35.3419
R10296 GND.n5226 GND.n1994 35.3419
R10297 GND.n5238 GND.n1994 35.3419
R10298 GND.n5238 GND.n1985 35.3419
R10299 GND.n5246 GND.n1985 35.3419
R10300 GND.n5246 GND.n1974 35.3419
R10301 GND.n5258 GND.n1974 35.3419
R10302 GND.n5266 GND.n1965 35.3419
R10303 GND.n5266 GND.n1954 35.3419
R10304 GND.n5278 GND.n1954 35.3419
R10305 GND.n5278 GND.n1945 35.3419
R10306 GND.n5286 GND.n1945 35.3419
R10307 GND.n5286 GND.n1934 35.3419
R10308 GND.n5298 GND.n1934 35.3419
R10309 GND.n5298 GND.n1925 35.3419
R10310 GND.n5306 GND.n1925 35.3419
R10311 GND.n5306 GND.n1914 35.3419
R10312 GND.n5323 GND.n1914 35.3419
R10313 GND.n5323 GND.n1904 35.3419
R10314 GND.n5333 GND.n1904 35.3419
R10315 GND.n5333 GND.n1897 35.3419
R10316 GND.n5357 GND.n1897 35.3419
R10317 GND.n5368 GND.n1878 35.3419
R10318 GND.n5378 GND.n1878 35.3419
R10319 GND.n5378 GND.n1869 35.3419
R10320 GND.n5387 GND.n1869 35.3419
R10321 GND.n5387 GND.n1630 35.3419
R10322 GND.n6286 GND.n1630 35.3419
R10323 GND.n6286 GND.n1634 35.3419
R10324 GND.n1637 GND.n1634 35.3419
R10325 GND.n5403 GND.n1661 35.3419
R10326 GND.n5404 GND.n5403 35.3419
R10327 GND.n5404 GND.n1824 35.3419
R10328 GND.n1855 GND.n1846 35.3419
R10329 GND.n7505 GND.n839 35.3419
R10330 GND.n7498 GND.n851 35.3419
R10331 GND.n7498 GND.n7497 35.3419
R10332 GND.n7497 GND.n679 35.3419
R10333 GND.n7702 GND.n670 35.3419
R10334 GND.n7710 GND.n670 35.3419
R10335 GND.n7710 GND.n658 35.3419
R10336 GND.n7724 GND.n658 35.3419
R10337 GND.n7724 GND.n649 35.3419
R10338 GND.n7732 GND.n649 35.3419
R10339 GND.n7732 GND.n638 35.3419
R10340 GND.n7744 GND.n638 35.3419
R10341 GND.n7752 GND.n629 35.3419
R10342 GND.n7752 GND.n618 35.3419
R10343 GND.n7764 GND.n618 35.3419
R10344 GND.n7764 GND.n609 35.3419
R10345 GND.n7772 GND.n609 35.3419
R10346 GND.n7772 GND.n598 35.3419
R10347 GND.n7784 GND.n598 35.3419
R10348 GND.n7784 GND.n589 35.3419
R10349 GND.n7792 GND.n589 35.3419
R10350 GND.n7792 GND.n577 35.3419
R10351 GND.n7808 GND.n577 35.3419
R10352 GND.n7808 GND.n567 35.3419
R10353 GND.n7818 GND.n567 35.3419
R10354 GND.n7818 GND.n560 35.3419
R10355 GND.n7871 GND.n560 35.3419
R10356 GND.n7882 GND.n541 35.3419
R10357 GND.n7890 GND.n541 35.3419
R10358 GND.n7890 GND.n530 35.3419
R10359 GND.n7902 GND.n530 35.3419
R10360 GND.n7902 GND.n521 35.3419
R10361 GND.n7910 GND.n521 35.3419
R10362 GND.n7910 GND.n510 35.3419
R10363 GND.n7922 GND.n510 35.3419
R10364 GND.n7922 GND.n501 35.3419
R10365 GND.n7930 GND.n501 35.3419
R10366 GND.n7930 GND.n489 35.3419
R10367 GND.n7949 GND.n489 35.3419
R10368 GND.n7957 GND.n480 35.3419
R10369 GND.n7957 GND.n119 35.3419
R10370 GND.n8600 GND.n119 35.3419
R10371 GND.n8600 GND.n110 35.3419
R10372 GND.n8608 GND.n110 35.3419
R10373 GND.n8608 GND.n88 35.3419
R10374 GND.n8630 GND.n88 35.3419
R10375 GND.n8630 GND.n91 35.3419
R10376 GND.n8624 GND.n91 35.3419
R10377 GND.n8624 GND.n103 35.3419
R10378 GND.n103 GND.n68 35.3419
R10379 GND.t25 GND.n68 35.3419
R10380 GND.t25 GND.n71 35.3419
R10381 GND.n8579 GND.n71 35.3419
R10382 GND.n8579 GND.n136 35.3419
R10383 GND.n8572 GND.n136 35.3419
R10384 GND.n8572 GND.n142 35.3419
R10385 GND.n8566 GND.n142 35.3419
R10386 GND.n8566 GND.n154 35.3419
R10387 GND.n8560 GND.n154 35.3419
R10388 GND.n8560 GND.n164 35.3419
R10389 GND.n8554 GND.n164 35.3419
R10390 GND.n8554 GND.n174 35.3419
R10391 GND.n8548 GND.n174 35.3419
R10392 GND.n8542 GND.n192 35.3419
R10393 GND.n8542 GND.n195 35.3419
R10394 GND.n8536 GND.n195 35.3419
R10395 GND.n8536 GND.n206 35.3419
R10396 GND.n8530 GND.n206 35.3419
R10397 GND.n8530 GND.n216 35.3419
R10398 GND.n8524 GND.n216 35.3419
R10399 GND.n8524 GND.n227 35.3419
R10400 GND.n8518 GND.n227 35.3419
R10401 GND.n8518 GND.n237 35.3419
R10402 GND.n8512 GND.n237 35.3419
R10403 GND.n8512 GND.n248 35.3419
R10404 GND.n8506 GND.n258 35.3419
R10405 GND.n8500 GND.n258 35.3419
R10406 GND.n8500 GND.n269 35.3419
R10407 GND.n8494 GND.n269 35.3419
R10408 GND.n8494 GND.n279 35.3419
R10409 GND.n8488 GND.n279 35.3419
R10410 GND.n8488 GND.n290 35.3419
R10411 GND.n8482 GND.n290 35.3419
R10412 GND.n8482 GND.n300 35.3419
R10413 GND.n8476 GND.n300 35.3419
R10414 GND.n8476 GND.n311 35.3419
R10415 GND.n8470 GND.n311 35.3419
R10416 GND.n8470 GND.n321 35.3419
R10417 GND.n8464 GND.n321 35.3419
R10418 GND.n8464 GND.n332 35.3419
R10419 GND.n8458 GND.n342 35.3419
R10420 GND.n8069 GND.n342 35.3419
R10421 GND.n8316 GND.n8069 35.3419
R10422 GND.n8316 GND.n449 35.3419
R10423 GND.n8326 GND.n449 35.3419
R10424 GND.n8326 GND.n350 35.3419
R10425 GND.n6282 GND.n1661 34.9885
R10426 GND.n7701 GND.n679 34.9885
R10427 GND.n2848 GND.t89 31.1009
R10428 GND.n5368 GND.t126 31.1009
R10429 GND.n7744 GND.t134 31.1009
R10430 GND.n8458 GND.t110 31.1009
R10431 GND.n6242 GND.n6241 30.7205
R10432 GND.n7654 GND.n7559 30.7205
R10433 GND.n6237 GND.n1824 28.627
R10434 GND.n7556 GND.n851 28.627
R10435 GND.t19 GND.n2273 26.8599
R10436 GND.n5187 GND.t30 26.8599
R10437 GND.t44 GND.n480 26.8599
R10438 GND.n8548 GND.t23 26.8599
R10439 GND.n6191 GND.n1852 24.0326
R10440 GND.n5494 GND.n5416 24.0326
R10441 GND.n6177 GND.n5424 24.0326
R10442 GND.n6170 GND.n5435 24.0326
R10443 GND.n6170 GND.n5437 24.0326
R10444 GND.n6158 GND.n5516 24.0326
R10445 GND.n5597 GND.n5530 24.0326
R10446 GND.n6144 GND.n5538 24.0326
R10447 GND.n5610 GND.n5548 24.0326
R10448 GND.n6130 GND.n5556 24.0326
R10449 GND.n5623 GND.n5566 24.0326
R10450 GND.n6116 GND.n5574 24.0326
R10451 GND.n6109 GND.n5585 24.0326
R10452 GND.n6097 GND.n5648 24.0326
R10453 GND.n5730 GND.n5661 24.0326
R10454 GND.n6083 GND.n5669 24.0326
R10455 GND.n5743 GND.n5679 24.0326
R10456 GND.n6069 GND.n5687 24.0326
R10457 GND.n5756 GND.n5697 24.0326
R10458 GND.n6055 GND.n5705 24.0326
R10459 GND.n6048 GND.n5716 24.0326
R10460 GND.n6048 GND.n5718 24.0326
R10461 GND.n6036 GND.n5779 24.0326
R10462 GND.n5860 GND.n5792 24.0326
R10463 GND.n6022 GND.n5800 24.0326
R10464 GND.n5874 GND.n5809 24.0326
R10465 GND.n6008 GND.n5817 24.0326
R10466 GND.n5887 GND.n5827 24.0326
R10467 GND.n5994 GND.n5835 24.0326
R10468 GND.n5987 GND.n5846 24.0326
R10469 GND.n5987 GND.n5848 24.0326
R10470 GND.n5940 GND.n5923 24.0326
R10471 GND.n5961 GND.n5931 24.0326
R10472 GND.n7009 GND.n1157 24.0326
R10473 GND.n7033 GND.n1141 24.0326
R10474 GND.n7056 GND.n1124 24.0326
R10475 GND.n7056 GND.n1126 24.0326
R10476 GND.n7082 GND.n1110 24.0326
R10477 GND.n7089 GND.n7088 24.0326
R10478 GND.n7107 GND.n1096 24.0326
R10479 GND.n7113 GND.n1092 24.0326
R10480 GND.n7131 GND.n1076 24.0326
R10481 GND.n7142 GND.n1065 24.0326
R10482 GND.n7163 GND.n1056 24.0326
R10483 GND.n7169 GND.n1047 24.0326
R10484 GND.n7181 GND.n1047 24.0326
R10485 GND.n7187 GND.n1043 24.0326
R10486 GND.n7214 GND.n1027 24.0326
R10487 GND.n7221 GND.n7220 24.0326
R10488 GND.n7239 GND.n1013 24.0326
R10489 GND.n7245 GND.n1009 24.0326
R10490 GND.n7263 GND.n993 24.0326
R10491 GND.n7274 GND.n982 24.0326
R10492 GND.n7294 GND.n973 24.0326
R10493 GND.n7312 GND.n963 24.0326
R10494 GND.n7318 GND.n959 24.0326
R10495 GND.n7336 GND.n943 24.0326
R10496 GND.n7347 GND.n932 24.0326
R10497 GND.n7363 GND.n924 24.0326
R10498 GND.n7370 GND.n915 24.0326
R10499 GND.n7390 GND.n7389 24.0326
R10500 GND.n7407 GND.n898 24.0326
R10501 GND.n7407 GND.n892 24.0326
R10502 GND.n7423 GND.n884 24.0326
R10503 GND.n7430 GND.n875 24.0326
R10504 GND.n7507 GND.n7506 24.0326
R10505 GND.n6176 GND.n5426 22.619
R10506 GND.n6115 GND.n5576 22.619
R10507 GND.n6103 GND.n5637 22.619
R10508 GND.n6054 GND.n5707 22.619
R10509 GND.n6042 GND.n5770 22.619
R10510 GND.n5993 GND.n5837 22.619
R10511 GND.n5981 GND.n5901 22.619
R10512 GND.n7048 GND.n1131 22.619
R10513 GND.n7076 GND.n7075 22.619
R10514 GND.n7162 GND.n1058 22.619
R10515 GND.n7188 GND.n1041 22.619
R10516 GND.n7281 GND.n7280 22.619
R10517 GND.n7300 GND.n969 22.619
R10518 GND.n7413 GND.n894 22.619
R10519 GND.n6184 GND.n6183 21.2053
R10520 GND.n5594 GND.n5518 21.2053
R10521 GND.n6123 GND.n6122 21.2053
R10522 GND.n5727 GND.n5650 21.2053
R10523 GND.n6062 GND.n6061 21.2053
R10524 GND.n5857 GND.n5781 21.2053
R10525 GND.n6001 GND.n6000 21.2053
R10526 GND.n5937 GND.n5912 21.2053
R10527 GND.n1143 GND.n1142 21.2053
R10528 GND.n1111 GND.n1106 21.2053
R10529 GND.n7149 GND.n7148 21.2053
R10530 GND.n7208 GND.n7207 21.2053
R10531 GND.n995 GND.n994 21.2053
R10532 GND.n7319 GND.n957 21.2053
R10533 GND.n7378 GND.n7377 21.2053
R10534 GND.n886 GND.n879 21.2053
R10535 GND.n6190 GND.n1854 19.7917
R10536 GND.n6150 GND.n5532 19.7917
R10537 GND.n6129 GND.n5558 19.7917
R10538 GND.n6089 GND.n5663 19.7917
R10539 GND.n6068 GND.n5689 19.7917
R10540 GND.n6028 GND.n5794 19.7917
R10541 GND.n6007 GND.n5819 19.7917
R10542 GND.n5967 GND.n5925 19.7917
R10543 GND.n7027 GND.n1147 19.7917
R10544 GND.n7095 GND.n1102 19.7917
R10545 GND.n1078 GND.n1077 19.7917
R10546 GND.n1028 GND.n1023 19.7917
R10547 GND.n7257 GND.n999 19.7917
R10548 GND.n7330 GND.n7329 19.7917
R10549 GND.n7362 GND.n926 19.7917
R10550 GND.n7483 GND.n866 19.7917
R10551 GND.n2605 GND.n2574 19.3944
R10552 GND.n2609 GND.n2574 19.3944
R10553 GND.n2609 GND.n2558 19.3944
R10554 GND.n2718 GND.n2558 19.3944
R10555 GND.n2718 GND.n2555 19.3944
R10556 GND.n2846 GND.n2555 19.3944
R10557 GND.n2846 GND.n2556 19.3944
R10558 GND.n2842 GND.n2556 19.3944
R10559 GND.n2842 GND.n2841 19.3944
R10560 GND.n2841 GND.n2840 19.3944
R10561 GND.n2840 GND.n2724 19.3944
R10562 GND.n2836 GND.n2724 19.3944
R10563 GND.n2836 GND.n2835 19.3944
R10564 GND.n2835 GND.n2834 19.3944
R10565 GND.n2834 GND.n2728 19.3944
R10566 GND.n2830 GND.n2728 19.3944
R10567 GND.n2830 GND.n2829 19.3944
R10568 GND.n2829 GND.n2828 19.3944
R10569 GND.n2828 GND.n2732 19.3944
R10570 GND.n2824 GND.n2732 19.3944
R10571 GND.n2824 GND.n2823 19.3944
R10572 GND.n2823 GND.n2822 19.3944
R10573 GND.n2822 GND.n2736 19.3944
R10574 GND.n2818 GND.n2736 19.3944
R10575 GND.n2818 GND.n2817 19.3944
R10576 GND.n2817 GND.n2816 19.3944
R10577 GND.n2816 GND.n2740 19.3944
R10578 GND.n2812 GND.n2740 19.3944
R10579 GND.n2812 GND.n2811 19.3944
R10580 GND.n2811 GND.n2810 19.3944
R10581 GND.n2810 GND.n2744 19.3944
R10582 GND.n2806 GND.n2744 19.3944
R10583 GND.n2806 GND.n2805 19.3944
R10584 GND.n2805 GND.n2804 19.3944
R10585 GND.n2804 GND.n2748 19.3944
R10586 GND.n2800 GND.n2748 19.3944
R10587 GND.n2800 GND.n2799 19.3944
R10588 GND.n2799 GND.n2798 19.3944
R10589 GND.n2798 GND.n2752 19.3944
R10590 GND.n2794 GND.n2752 19.3944
R10591 GND.n2794 GND.n2793 19.3944
R10592 GND.n2793 GND.n2792 19.3944
R10593 GND.n2792 GND.n2757 19.3944
R10594 GND.n2788 GND.n2757 19.3944
R10595 GND.n2788 GND.n2787 19.3944
R10596 GND.n2787 GND.n2786 19.3944
R10597 GND.n2786 GND.n2761 19.3944
R10598 GND.n2762 GND.n2761 19.3944
R10599 GND.n2781 GND.n2762 19.3944
R10600 GND.n2781 GND.n2779 19.3944
R10601 GND.n2779 GND.n2778 19.3944
R10602 GND.n2778 GND.n2776 19.3944
R10603 GND.n2776 GND.n2775 19.3944
R10604 GND.n2775 GND.n2773 19.3944
R10605 GND.n2773 GND.n2772 19.3944
R10606 GND.n2772 GND.n2770 19.3944
R10607 GND.n2770 GND.n2049 19.3944
R10608 GND.n5119 GND.n2049 19.3944
R10609 GND.n5119 GND.n2047 19.3944
R10610 GND.n5185 GND.n2047 19.3944
R10611 GND.n5185 GND.n5184 19.3944
R10612 GND.n5184 GND.n5183 19.3944
R10613 GND.n5183 GND.n5181 19.3944
R10614 GND.n5181 GND.n5180 19.3944
R10615 GND.n5180 GND.n5178 19.3944
R10616 GND.n5178 GND.n5177 19.3944
R10617 GND.n5177 GND.n5175 19.3944
R10618 GND.n5175 GND.n5174 19.3944
R10619 GND.n5174 GND.n5172 19.3944
R10620 GND.n5172 GND.n5171 19.3944
R10621 GND.n5171 GND.n5169 19.3944
R10622 GND.n5169 GND.n5168 19.3944
R10623 GND.n5168 GND.n5166 19.3944
R10624 GND.n5166 GND.n5165 19.3944
R10625 GND.n5165 GND.n5163 19.3944
R10626 GND.n5163 GND.n5162 19.3944
R10627 GND.n5162 GND.n5160 19.3944
R10628 GND.n5160 GND.n5159 19.3944
R10629 GND.n5159 GND.n5157 19.3944
R10630 GND.n5157 GND.n5156 19.3944
R10631 GND.n5156 GND.n5154 19.3944
R10632 GND.n5154 GND.n5153 19.3944
R10633 GND.n5153 GND.n5151 19.3944
R10634 GND.n5151 GND.n5150 19.3944
R10635 GND.n5150 GND.n5148 19.3944
R10636 GND.n5148 GND.n1902 19.3944
R10637 GND.n5335 GND.n1902 19.3944
R10638 GND.n5335 GND.n1900 19.3944
R10639 GND.n5355 GND.n1900 19.3944
R10640 GND.n5355 GND.n5354 19.3944
R10641 GND.n5354 GND.n5353 19.3944
R10642 GND.n5353 GND.n5351 19.3944
R10643 GND.n5351 GND.n5350 19.3944
R10644 GND.n5350 GND.n5348 19.3944
R10645 GND.n5348 GND.n5347 19.3944
R10646 GND.n5347 GND.n5345 19.3944
R10647 GND.n2865 GND.n2535 19.3944
R10648 GND.n2588 GND.n2535 19.3944
R10649 GND.n2588 GND.n2583 19.3944
R10650 GND.n2592 GND.n2583 19.3944
R10651 GND.n2593 GND.n2592 19.3944
R10652 GND.n2596 GND.n2593 19.3944
R10653 GND.n2596 GND.n2579 19.3944
R10654 GND.n2600 GND.n2579 19.3944
R10655 GND.n2859 GND.n2539 19.3944
R10656 GND.n2859 GND.n2858 19.3944
R10657 GND.n2858 GND.n2857 19.3944
R10658 GND.n2857 GND.n2545 19.3944
R10659 GND.n2853 GND.n2545 19.3944
R10660 GND.n2853 GND.n2852 19.3944
R10661 GND.n2852 GND.n2851 19.3944
R10662 GND.n2851 GND.n2419 19.3944
R10663 GND.n4862 GND.n2419 19.3944
R10664 GND.n4862 GND.n2420 19.3944
R10665 GND.n4858 GND.n2420 19.3944
R10666 GND.n4858 GND.n2399 19.3944
R10667 GND.n4882 GND.n2399 19.3944
R10668 GND.n4882 GND.n2400 19.3944
R10669 GND.n4878 GND.n2400 19.3944
R10670 GND.n4878 GND.n2379 19.3944
R10671 GND.n4902 GND.n2379 19.3944
R10672 GND.n4902 GND.n2380 19.3944
R10673 GND.n4898 GND.n2380 19.3944
R10674 GND.n4898 GND.n2359 19.3944
R10675 GND.n4922 GND.n2359 19.3944
R10676 GND.n4922 GND.n2360 19.3944
R10677 GND.n4918 GND.n2360 19.3944
R10678 GND.n4918 GND.n2339 19.3944
R10679 GND.n4942 GND.n2339 19.3944
R10680 GND.n4942 GND.n2340 19.3944
R10681 GND.n4938 GND.n2340 19.3944
R10682 GND.n4938 GND.n2319 19.3944
R10683 GND.n4962 GND.n2319 19.3944
R10684 GND.n4962 GND.n2320 19.3944
R10685 GND.n4958 GND.n2320 19.3944
R10686 GND.n4958 GND.n2299 19.3944
R10687 GND.n4982 GND.n2299 19.3944
R10688 GND.n4982 GND.n2300 19.3944
R10689 GND.n4978 GND.n2300 19.3944
R10690 GND.n4978 GND.n2279 19.3944
R10691 GND.n5002 GND.n2279 19.3944
R10692 GND.n5002 GND.n2280 19.3944
R10693 GND.n4998 GND.n2280 19.3944
R10694 GND.n4998 GND.n2259 19.3944
R10695 GND.n5028 GND.n2259 19.3944
R10696 GND.n5028 GND.n2260 19.3944
R10697 GND.n5024 GND.n2260 19.3944
R10698 GND.n5024 GND.n5023 19.3944
R10699 GND.n5023 GND.n2236 19.3944
R10700 GND.n5048 GND.n2236 19.3944
R10701 GND.n5048 GND.n2237 19.3944
R10702 GND.n5044 GND.n2237 19.3944
R10703 GND.n5044 GND.n2213 19.3944
R10704 GND.n5073 GND.n2213 19.3944
R10705 GND.n5073 GND.n2214 19.3944
R10706 GND.n5069 GND.n2214 19.3944
R10707 GND.n5069 GND.n5068 19.3944
R10708 GND.n5068 GND.n5067 19.3944
R10709 GND.n5067 GND.n2067 19.3944
R10710 GND.n5105 GND.n2067 19.3944
R10711 GND.n5105 GND.n2068 19.3944
R10712 GND.n5101 GND.n2068 19.3944
R10713 GND.n5101 GND.n5100 19.3944
R10714 GND.n5100 GND.n2039 19.3944
R10715 GND.n5196 GND.n2039 19.3944
R10716 GND.n5196 GND.n2040 19.3944
R10717 GND.n5192 GND.n2040 19.3944
R10718 GND.n5192 GND.n2020 19.3944
R10719 GND.n5216 GND.n2020 19.3944
R10720 GND.n5216 GND.n2021 19.3944
R10721 GND.n5212 GND.n2021 19.3944
R10722 GND.n5212 GND.n2000 19.3944
R10723 GND.n5236 GND.n2000 19.3944
R10724 GND.n5236 GND.n2001 19.3944
R10725 GND.n5232 GND.n2001 19.3944
R10726 GND.n5232 GND.n1980 19.3944
R10727 GND.n5256 GND.n1980 19.3944
R10728 GND.n5256 GND.n1981 19.3944
R10729 GND.n5252 GND.n1981 19.3944
R10730 GND.n5252 GND.n1960 19.3944
R10731 GND.n5276 GND.n1960 19.3944
R10732 GND.n5276 GND.n1961 19.3944
R10733 GND.n5272 GND.n1961 19.3944
R10734 GND.n5272 GND.n1940 19.3944
R10735 GND.n5296 GND.n1940 19.3944
R10736 GND.n5296 GND.n1941 19.3944
R10737 GND.n5292 GND.n1941 19.3944
R10738 GND.n5292 GND.n1920 19.3944
R10739 GND.n5321 GND.n1920 19.3944
R10740 GND.n5321 GND.n1921 19.3944
R10741 GND.n5317 GND.n1921 19.3944
R10742 GND.n5317 GND.n5316 19.3944
R10743 GND.n5316 GND.n1892 19.3944
R10744 GND.n5366 GND.n1892 19.3944
R10745 GND.n5366 GND.n1893 19.3944
R10746 GND.n5362 GND.n1893 19.3944
R10747 GND.n5362 GND.n1874 19.3944
R10748 GND.n5385 GND.n1874 19.3944
R10749 GND.n5385 GND.n1627 19.3944
R10750 GND.n6288 GND.n1627 19.3944
R10751 GND.n6280 GND.n1690 19.3944
R10752 GND.n6276 GND.n1690 19.3944
R10753 GND.n6276 GND.n6275 19.3944
R10754 GND.n6275 GND.n6274 19.3944
R10755 GND.n6274 GND.n1697 19.3944
R10756 GND.n6270 GND.n1697 19.3944
R10757 GND.n6270 GND.n6269 19.3944
R10758 GND.n6269 GND.n6268 19.3944
R10759 GND.n6264 GND.n6263 19.3944
R10760 GND.n6263 GND.n6262 19.3944
R10761 GND.n6262 GND.n1711 19.3944
R10762 GND.n6258 GND.n1711 19.3944
R10763 GND.n6258 GND.n6257 19.3944
R10764 GND.n6257 GND.n6256 19.3944
R10765 GND.n6256 GND.n1717 19.3944
R10766 GND.n6252 GND.n1717 19.3944
R10767 GND.n6252 GND.n6251 19.3944
R10768 GND.n6249 GND.n1726 19.3944
R10769 GND.n6245 GND.n1726 19.3944
R10770 GND.n1818 GND.n1730 19.3944
R10771 GND.n1814 GND.n1730 19.3944
R10772 GND.n1814 GND.n1813 19.3944
R10773 GND.n1813 GND.n1812 19.3944
R10774 GND.n1808 GND.n1807 19.3944
R10775 GND.n1807 GND.n1806 19.3944
R10776 GND.n1806 GND.n1744 19.3944
R10777 GND.n1802 GND.n1744 19.3944
R10778 GND.n1802 GND.n1801 19.3944
R10779 GND.n1801 GND.n1800 19.3944
R10780 GND.n1800 GND.n1750 19.3944
R10781 GND.n1796 GND.n1750 19.3944
R10782 GND.n1796 GND.n1795 19.3944
R10783 GND.n1793 GND.n1759 19.3944
R10784 GND.n1789 GND.n1759 19.3944
R10785 GND.n1789 GND.n1788 19.3944
R10786 GND.n1788 GND.n1787 19.3944
R10787 GND.n1787 GND.n1765 19.3944
R10788 GND.n1783 GND.n1765 19.3944
R10789 GND.n1783 GND.n1782 19.3944
R10790 GND.n1782 GND.n1781 19.3944
R10791 GND.n1781 GND.n1771 19.3944
R10792 GND.n3962 GND.n3784 19.3944
R10793 GND.n3956 GND.n3784 19.3944
R10794 GND.n3956 GND.n3955 19.3944
R10795 GND.n3955 GND.n3954 19.3944
R10796 GND.n3954 GND.n3791 19.3944
R10797 GND.n3948 GND.n3791 19.3944
R10798 GND.n3948 GND.n3947 19.3944
R10799 GND.n3947 GND.n3946 19.3944
R10800 GND.n3946 GND.n3799 19.3944
R10801 GND.n3940 GND.n3799 19.3944
R10802 GND.n3940 GND.n3939 19.3944
R10803 GND.n3939 GND.n3938 19.3944
R10804 GND.n3938 GND.n3807 19.3944
R10805 GND.n3932 GND.n3807 19.3944
R10806 GND.n3932 GND.n3931 19.3944
R10807 GND.n3931 GND.n3930 19.3944
R10808 GND.n3930 GND.n3815 19.3944
R10809 GND.n3924 GND.n3815 19.3944
R10810 GND.n3924 GND.n3923 19.3944
R10811 GND.n3923 GND.n3922 19.3944
R10812 GND.n3922 GND.n3823 19.3944
R10813 GND.n3916 GND.n3823 19.3944
R10814 GND.n3916 GND.n3915 19.3944
R10815 GND.n3915 GND.n3914 19.3944
R10816 GND.n3914 GND.n3831 19.3944
R10817 GND.n3908 GND.n3831 19.3944
R10818 GND.n3908 GND.n3907 19.3944
R10819 GND.n3907 GND.n3906 19.3944
R10820 GND.n3906 GND.n3839 19.3944
R10821 GND.n3900 GND.n3839 19.3944
R10822 GND.n3900 GND.n3899 19.3944
R10823 GND.n3899 GND.n3898 19.3944
R10824 GND.n3898 GND.n3847 19.3944
R10825 GND.n3892 GND.n3847 19.3944
R10826 GND.n3892 GND.n3891 19.3944
R10827 GND.n3891 GND.n3890 19.3944
R10828 GND.n3890 GND.n3855 19.3944
R10829 GND.n3884 GND.n3855 19.3944
R10830 GND.n3884 GND.n3883 19.3944
R10831 GND.n3883 GND.n3882 19.3944
R10832 GND.n3882 GND.n3863 19.3944
R10833 GND.n3876 GND.n3863 19.3944
R10834 GND.n3876 GND.n3875 19.3944
R10835 GND.n3875 GND.n3874 19.3944
R10836 GND.n3874 GND.n347 19.3944
R10837 GND.n8452 GND.n347 19.3944
R10838 GND.n8453 GND.n8452 19.3944
R10839 GND.n4725 GND.n4724 19.3944
R10840 GND.n4724 GND.n3024 19.3944
R10841 GND.n4718 GND.n3024 19.3944
R10842 GND.n4718 GND.n4717 19.3944
R10843 GND.n4717 GND.n4716 19.3944
R10844 GND.n4716 GND.n3033 19.3944
R10845 GND.n4710 GND.n3033 19.3944
R10846 GND.n4710 GND.n4709 19.3944
R10847 GND.n4709 GND.n4708 19.3944
R10848 GND.n4708 GND.n3041 19.3944
R10849 GND.n4702 GND.n3041 19.3944
R10850 GND.n4702 GND.n4701 19.3944
R10851 GND.n4701 GND.n4700 19.3944
R10852 GND.n4700 GND.n3049 19.3944
R10853 GND.n4694 GND.n3049 19.3944
R10854 GND.n4694 GND.n4693 19.3944
R10855 GND.n4693 GND.n4692 19.3944
R10856 GND.n4692 GND.n3057 19.3944
R10857 GND.n4686 GND.n3057 19.3944
R10858 GND.n4686 GND.n4685 19.3944
R10859 GND.n4685 GND.n4684 19.3944
R10860 GND.n4684 GND.n3065 19.3944
R10861 GND.n4678 GND.n3065 19.3944
R10862 GND.n4678 GND.n4677 19.3944
R10863 GND.n4677 GND.n4676 19.3944
R10864 GND.n4676 GND.n3073 19.3944
R10865 GND.n4670 GND.n3073 19.3944
R10866 GND.n4670 GND.n4669 19.3944
R10867 GND.n4669 GND.n4668 19.3944
R10868 GND.n4668 GND.n3081 19.3944
R10869 GND.n4662 GND.n3081 19.3944
R10870 GND.n4662 GND.n4661 19.3944
R10871 GND.n4661 GND.n4660 19.3944
R10872 GND.n4660 GND.n3089 19.3944
R10873 GND.n4654 GND.n3089 19.3944
R10874 GND.n4654 GND.n4653 19.3944
R10875 GND.n4653 GND.n4652 19.3944
R10876 GND.n4652 GND.n3097 19.3944
R10877 GND.n4646 GND.n3097 19.3944
R10878 GND.n4646 GND.n4645 19.3944
R10879 GND.n4645 GND.n4644 19.3944
R10880 GND.n4644 GND.n3105 19.3944
R10881 GND.n4638 GND.n3105 19.3944
R10882 GND.n4638 GND.n4637 19.3944
R10883 GND.n4637 GND.n4636 19.3944
R10884 GND.n4636 GND.n3113 19.3944
R10885 GND.n4630 GND.n3113 19.3944
R10886 GND.n4630 GND.n4629 19.3944
R10887 GND.n4629 GND.n4628 19.3944
R10888 GND.n4628 GND.n3121 19.3944
R10889 GND.n4622 GND.n3121 19.3944
R10890 GND.n4622 GND.n4621 19.3944
R10891 GND.n4621 GND.n4620 19.3944
R10892 GND.n4620 GND.n3129 19.3944
R10893 GND.n4614 GND.n3129 19.3944
R10894 GND.n4614 GND.n4613 19.3944
R10895 GND.n4613 GND.n4612 19.3944
R10896 GND.n4612 GND.n3137 19.3944
R10897 GND.n4606 GND.n3137 19.3944
R10898 GND.n4606 GND.n4605 19.3944
R10899 GND.n4605 GND.n4604 19.3944
R10900 GND.n4604 GND.n3145 19.3944
R10901 GND.n4598 GND.n3145 19.3944
R10902 GND.n4598 GND.n4597 19.3944
R10903 GND.n4597 GND.n4596 19.3944
R10904 GND.n4596 GND.n3153 19.3944
R10905 GND.n4590 GND.n3153 19.3944
R10906 GND.n4590 GND.n4589 19.3944
R10907 GND.n4589 GND.n4588 19.3944
R10908 GND.n4588 GND.n3161 19.3944
R10909 GND.n4582 GND.n3161 19.3944
R10910 GND.n4582 GND.n4581 19.3944
R10911 GND.n4581 GND.n4580 19.3944
R10912 GND.n4580 GND.n3169 19.3944
R10913 GND.n4574 GND.n3169 19.3944
R10914 GND.n4574 GND.n4573 19.3944
R10915 GND.n4573 GND.n4572 19.3944
R10916 GND.n4572 GND.n3177 19.3944
R10917 GND.n4566 GND.n3177 19.3944
R10918 GND.n4566 GND.n4565 19.3944
R10919 GND.n4565 GND.n4564 19.3944
R10920 GND.n4564 GND.n3185 19.3944
R10921 GND.n4558 GND.n3185 19.3944
R10922 GND.n4558 GND.n4557 19.3944
R10923 GND.n4557 GND.n4556 19.3944
R10924 GND.n4556 GND.n3193 19.3944
R10925 GND.n4550 GND.n3193 19.3944
R10926 GND.n4550 GND.n4549 19.3944
R10927 GND.n4549 GND.n4548 19.3944
R10928 GND.n4548 GND.n3201 19.3944
R10929 GND.n4542 GND.n3201 19.3944
R10930 GND.n4542 GND.n4541 19.3944
R10931 GND.n4541 GND.n4540 19.3944
R10932 GND.n4540 GND.n3209 19.3944
R10933 GND.n4534 GND.n3209 19.3944
R10934 GND.n4534 GND.n4533 19.3944
R10935 GND.n4533 GND.n4532 19.3944
R10936 GND.n4532 GND.n3217 19.3944
R10937 GND.n4526 GND.n3217 19.3944
R10938 GND.n4526 GND.n4525 19.3944
R10939 GND.n4525 GND.n4524 19.3944
R10940 GND.n4524 GND.n3225 19.3944
R10941 GND.n4518 GND.n3225 19.3944
R10942 GND.n4518 GND.n4517 19.3944
R10943 GND.n4517 GND.n4516 19.3944
R10944 GND.n4516 GND.n3233 19.3944
R10945 GND.n4510 GND.n3233 19.3944
R10946 GND.n4510 GND.n4509 19.3944
R10947 GND.n4509 GND.n4508 19.3944
R10948 GND.n4508 GND.n3241 19.3944
R10949 GND.n4502 GND.n3241 19.3944
R10950 GND.n4502 GND.n4501 19.3944
R10951 GND.n4501 GND.n4500 19.3944
R10952 GND.n4500 GND.n3249 19.3944
R10953 GND.n4494 GND.n3249 19.3944
R10954 GND.n4494 GND.n4493 19.3944
R10955 GND.n4493 GND.n4492 19.3944
R10956 GND.n4492 GND.n3257 19.3944
R10957 GND.n4486 GND.n3257 19.3944
R10958 GND.n4486 GND.n4485 19.3944
R10959 GND.n4485 GND.n4484 19.3944
R10960 GND.n4484 GND.n3265 19.3944
R10961 GND.n4478 GND.n3265 19.3944
R10962 GND.n4478 GND.n4477 19.3944
R10963 GND.n4477 GND.n4476 19.3944
R10964 GND.n4476 GND.n3273 19.3944
R10965 GND.n4470 GND.n3273 19.3944
R10966 GND.n4470 GND.n4469 19.3944
R10967 GND.n4469 GND.n4468 19.3944
R10968 GND.n4468 GND.n3281 19.3944
R10969 GND.n4462 GND.n3281 19.3944
R10970 GND.n4462 GND.n4461 19.3944
R10971 GND.n4461 GND.n4460 19.3944
R10972 GND.n4460 GND.n3289 19.3944
R10973 GND.n4454 GND.n3289 19.3944
R10974 GND.n4454 GND.n4453 19.3944
R10975 GND.n4453 GND.n4452 19.3944
R10976 GND.n4452 GND.n3297 19.3944
R10977 GND.n4446 GND.n3297 19.3944
R10978 GND.n4446 GND.n4445 19.3944
R10979 GND.n4445 GND.n4444 19.3944
R10980 GND.n4444 GND.n3305 19.3944
R10981 GND.n4438 GND.n3305 19.3944
R10982 GND.n4438 GND.n4437 19.3944
R10983 GND.n4437 GND.n4436 19.3944
R10984 GND.n4436 GND.n3313 19.3944
R10985 GND.n4430 GND.n3313 19.3944
R10986 GND.n4430 GND.n4429 19.3944
R10987 GND.n4429 GND.n4428 19.3944
R10988 GND.n4428 GND.n3321 19.3944
R10989 GND.n4422 GND.n3321 19.3944
R10990 GND.n4422 GND.n4421 19.3944
R10991 GND.n4421 GND.n4420 19.3944
R10992 GND.n4420 GND.n3329 19.3944
R10993 GND.n4414 GND.n3329 19.3944
R10994 GND.n4414 GND.n4413 19.3944
R10995 GND.n4413 GND.n4412 19.3944
R10996 GND.n4412 GND.n3337 19.3944
R10997 GND.n4406 GND.n3337 19.3944
R10998 GND.n4406 GND.n4405 19.3944
R10999 GND.n4405 GND.n4404 19.3944
R11000 GND.n4404 GND.n3345 19.3944
R11001 GND.n4398 GND.n3345 19.3944
R11002 GND.n4398 GND.n4397 19.3944
R11003 GND.n4397 GND.n4396 19.3944
R11004 GND.n4396 GND.n3353 19.3944
R11005 GND.n4390 GND.n3353 19.3944
R11006 GND.n4390 GND.n4389 19.3944
R11007 GND.n4389 GND.n4388 19.3944
R11008 GND.n4388 GND.n3361 19.3944
R11009 GND.n4382 GND.n3361 19.3944
R11010 GND.n4382 GND.n4381 19.3944
R11011 GND.n4381 GND.n4380 19.3944
R11012 GND.n4380 GND.n3369 19.3944
R11013 GND.n4374 GND.n3369 19.3944
R11014 GND.n4374 GND.n4373 19.3944
R11015 GND.n4373 GND.n4372 19.3944
R11016 GND.n4372 GND.n3377 19.3944
R11017 GND.n4366 GND.n3377 19.3944
R11018 GND.n4366 GND.n4365 19.3944
R11019 GND.n4365 GND.n4364 19.3944
R11020 GND.n4364 GND.n3385 19.3944
R11021 GND.n4358 GND.n3385 19.3944
R11022 GND.n4358 GND.n4357 19.3944
R11023 GND.n4357 GND.n4356 19.3944
R11024 GND.n4356 GND.n3393 19.3944
R11025 GND.n4350 GND.n3393 19.3944
R11026 GND.n4350 GND.n4349 19.3944
R11027 GND.n4349 GND.n4348 19.3944
R11028 GND.n4348 GND.n3401 19.3944
R11029 GND.n4342 GND.n3401 19.3944
R11030 GND.n4342 GND.n4341 19.3944
R11031 GND.n4341 GND.n4340 19.3944
R11032 GND.n4340 GND.n3409 19.3944
R11033 GND.n4334 GND.n3409 19.3944
R11034 GND.n4334 GND.n4333 19.3944
R11035 GND.n4333 GND.n4332 19.3944
R11036 GND.n4332 GND.n3417 19.3944
R11037 GND.n4326 GND.n3417 19.3944
R11038 GND.n4326 GND.n4325 19.3944
R11039 GND.n4325 GND.n4324 19.3944
R11040 GND.n4324 GND.n3425 19.3944
R11041 GND.n4318 GND.n3425 19.3944
R11042 GND.n4318 GND.n4317 19.3944
R11043 GND.n4317 GND.n4316 19.3944
R11044 GND.n4316 GND.n3433 19.3944
R11045 GND.n4310 GND.n3433 19.3944
R11046 GND.n4310 GND.n4309 19.3944
R11047 GND.n4309 GND.n4308 19.3944
R11048 GND.n4308 GND.n3441 19.3944
R11049 GND.n4302 GND.n3441 19.3944
R11050 GND.n4302 GND.n4301 19.3944
R11051 GND.n4301 GND.n4300 19.3944
R11052 GND.n4300 GND.n3449 19.3944
R11053 GND.n4294 GND.n3449 19.3944
R11054 GND.n4294 GND.n4293 19.3944
R11055 GND.n4293 GND.n4292 19.3944
R11056 GND.n4292 GND.n3457 19.3944
R11057 GND.n4286 GND.n3457 19.3944
R11058 GND.n4286 GND.n4285 19.3944
R11059 GND.n4285 GND.n4284 19.3944
R11060 GND.n4284 GND.n3465 19.3944
R11061 GND.n4278 GND.n3465 19.3944
R11062 GND.n4278 GND.n4277 19.3944
R11063 GND.n4277 GND.n4276 19.3944
R11064 GND.n4276 GND.n3473 19.3944
R11065 GND.n4270 GND.n3473 19.3944
R11066 GND.n4270 GND.n4269 19.3944
R11067 GND.n4269 GND.n4268 19.3944
R11068 GND.n4268 GND.n3481 19.3944
R11069 GND.n4262 GND.n3481 19.3944
R11070 GND.n4262 GND.n4261 19.3944
R11071 GND.n4261 GND.n4260 19.3944
R11072 GND.n4260 GND.n3489 19.3944
R11073 GND.n4254 GND.n3489 19.3944
R11074 GND.n4254 GND.n4253 19.3944
R11075 GND.n4253 GND.n4252 19.3944
R11076 GND.n4252 GND.n3497 19.3944
R11077 GND.n4246 GND.n3497 19.3944
R11078 GND.n4246 GND.n4245 19.3944
R11079 GND.n4245 GND.n4244 19.3944
R11080 GND.n4244 GND.n3505 19.3944
R11081 GND.n4238 GND.n3505 19.3944
R11082 GND.n4238 GND.n4237 19.3944
R11083 GND.n4237 GND.n4236 19.3944
R11084 GND.n4236 GND.n3513 19.3944
R11085 GND.n4230 GND.n3513 19.3944
R11086 GND.n4230 GND.n4229 19.3944
R11087 GND.n4229 GND.n4228 19.3944
R11088 GND.n4228 GND.n3521 19.3944
R11089 GND.n4222 GND.n3521 19.3944
R11090 GND.n4222 GND.n4221 19.3944
R11091 GND.n4221 GND.n4220 19.3944
R11092 GND.n4220 GND.n3529 19.3944
R11093 GND.n4214 GND.n3529 19.3944
R11094 GND.n4214 GND.n4213 19.3944
R11095 GND.n4213 GND.n4212 19.3944
R11096 GND.n4212 GND.n3537 19.3944
R11097 GND.n4206 GND.n3537 19.3944
R11098 GND.n4206 GND.n4205 19.3944
R11099 GND.n4205 GND.n4204 19.3944
R11100 GND.n4204 GND.n3545 19.3944
R11101 GND.n4198 GND.n3545 19.3944
R11102 GND.n4198 GND.n4197 19.3944
R11103 GND.n4197 GND.n4196 19.3944
R11104 GND.n4196 GND.n3553 19.3944
R11105 GND.n4190 GND.n3553 19.3944
R11106 GND.n4190 GND.n4189 19.3944
R11107 GND.n4189 GND.n4188 19.3944
R11108 GND.n4188 GND.n3561 19.3944
R11109 GND.n4182 GND.n3561 19.3944
R11110 GND.n4182 GND.n4181 19.3944
R11111 GND.n4181 GND.n4180 19.3944
R11112 GND.n4180 GND.n3569 19.3944
R11113 GND.n4174 GND.n3569 19.3944
R11114 GND.n4174 GND.n4173 19.3944
R11115 GND.n4173 GND.n4172 19.3944
R11116 GND.n4172 GND.n3577 19.3944
R11117 GND.n4166 GND.n3577 19.3944
R11118 GND.n4166 GND.n4165 19.3944
R11119 GND.n4165 GND.n4164 19.3944
R11120 GND.n4164 GND.n3585 19.3944
R11121 GND.n4158 GND.n3585 19.3944
R11122 GND.n4158 GND.n4157 19.3944
R11123 GND.n4157 GND.n4156 19.3944
R11124 GND.n4156 GND.n3593 19.3944
R11125 GND.n4150 GND.n3593 19.3944
R11126 GND.n4150 GND.n4149 19.3944
R11127 GND.n4149 GND.n4148 19.3944
R11128 GND.n4148 GND.n3601 19.3944
R11129 GND.n4142 GND.n3601 19.3944
R11130 GND.n4142 GND.n4141 19.3944
R11131 GND.n4141 GND.n4140 19.3944
R11132 GND.n4140 GND.n3609 19.3944
R11133 GND.n4134 GND.n3609 19.3944
R11134 GND.n4134 GND.n4133 19.3944
R11135 GND.n4133 GND.n4132 19.3944
R11136 GND.n4132 GND.n3617 19.3944
R11137 GND.n4126 GND.n3617 19.3944
R11138 GND.n4126 GND.n4125 19.3944
R11139 GND.n4125 GND.n4124 19.3944
R11140 GND.n4124 GND.n3625 19.3944
R11141 GND.n4118 GND.n3625 19.3944
R11142 GND.n4118 GND.n4117 19.3944
R11143 GND.n4117 GND.n4116 19.3944
R11144 GND.n4116 GND.n3633 19.3944
R11145 GND.n4110 GND.n3633 19.3944
R11146 GND.n4110 GND.n4109 19.3944
R11147 GND.n4109 GND.n4108 19.3944
R11148 GND.n4108 GND.n3641 19.3944
R11149 GND.n4102 GND.n3641 19.3944
R11150 GND.n4102 GND.n4101 19.3944
R11151 GND.n4101 GND.n4100 19.3944
R11152 GND.n4100 GND.n3649 19.3944
R11153 GND.n4094 GND.n3649 19.3944
R11154 GND.n4094 GND.n4093 19.3944
R11155 GND.n4093 GND.n4092 19.3944
R11156 GND.n4092 GND.n3657 19.3944
R11157 GND.n4086 GND.n3657 19.3944
R11158 GND.n4086 GND.n4085 19.3944
R11159 GND.n4085 GND.n4084 19.3944
R11160 GND.n4084 GND.n3665 19.3944
R11161 GND.n4078 GND.n3665 19.3944
R11162 GND.n4078 GND.n4077 19.3944
R11163 GND.n4077 GND.n4076 19.3944
R11164 GND.n4076 GND.n3673 19.3944
R11165 GND.n4070 GND.n3673 19.3944
R11166 GND.n4070 GND.n4069 19.3944
R11167 GND.n4069 GND.n4068 19.3944
R11168 GND.n4068 GND.n3681 19.3944
R11169 GND.n4062 GND.n3681 19.3944
R11170 GND.n4062 GND.n4061 19.3944
R11171 GND.n4061 GND.n4060 19.3944
R11172 GND.n4060 GND.n3689 19.3944
R11173 GND.n4054 GND.n3689 19.3944
R11174 GND.n4054 GND.n4053 19.3944
R11175 GND.n4053 GND.n4052 19.3944
R11176 GND.n4052 GND.n3697 19.3944
R11177 GND.n4046 GND.n3697 19.3944
R11178 GND.n4046 GND.n4045 19.3944
R11179 GND.n4045 GND.n4044 19.3944
R11180 GND.n4044 GND.n3705 19.3944
R11181 GND.n4038 GND.n3705 19.3944
R11182 GND.n4038 GND.n4037 19.3944
R11183 GND.n4037 GND.n4036 19.3944
R11184 GND.n4036 GND.n3713 19.3944
R11185 GND.n4030 GND.n3713 19.3944
R11186 GND.n4030 GND.n4029 19.3944
R11187 GND.n4029 GND.n4028 19.3944
R11188 GND.n4028 GND.n3721 19.3944
R11189 GND.n4022 GND.n3721 19.3944
R11190 GND.n4022 GND.n4021 19.3944
R11191 GND.n4021 GND.n4020 19.3944
R11192 GND.n4020 GND.n3729 19.3944
R11193 GND.n4014 GND.n3729 19.3944
R11194 GND.n4014 GND.n4013 19.3944
R11195 GND.n4013 GND.n4012 19.3944
R11196 GND.n4012 GND.n3737 19.3944
R11197 GND.n4006 GND.n3737 19.3944
R11198 GND.n4006 GND.n4005 19.3944
R11199 GND.n4005 GND.n4004 19.3944
R11200 GND.n4004 GND.n3745 19.3944
R11201 GND.n3998 GND.n3745 19.3944
R11202 GND.n3998 GND.n3997 19.3944
R11203 GND.n3997 GND.n3996 19.3944
R11204 GND.n3996 GND.n3753 19.3944
R11205 GND.n3990 GND.n3753 19.3944
R11206 GND.n3990 GND.n3989 19.3944
R11207 GND.n3989 GND.n3988 19.3944
R11208 GND.n3988 GND.n3761 19.3944
R11209 GND.n3982 GND.n3761 19.3944
R11210 GND.n3982 GND.n3981 19.3944
R11211 GND.n3981 GND.n3980 19.3944
R11212 GND.n3980 GND.n3769 19.3944
R11213 GND.n3974 GND.n3769 19.3944
R11214 GND.n3974 GND.n3973 19.3944
R11215 GND.n3973 GND.n3972 19.3944
R11216 GND.n3972 GND.n3777 19.3944
R11217 GND.n3966 GND.n3777 19.3944
R11218 GND.n3966 GND.n3965 19.3944
R11219 GND.n7698 GND.n7697 19.3944
R11220 GND.n7697 GND.n7696 19.3944
R11221 GND.n7696 GND.n7695 19.3944
R11222 GND.n7695 GND.n7693 19.3944
R11223 GND.n7693 GND.n7690 19.3944
R11224 GND.n7690 GND.n7689 19.3944
R11225 GND.n7689 GND.n7686 19.3944
R11226 GND.n7686 GND.n7685 19.3944
R11227 GND.n7681 GND.n7678 19.3944
R11228 GND.n7678 GND.n7677 19.3944
R11229 GND.n7677 GND.n7674 19.3944
R11230 GND.n7674 GND.n7673 19.3944
R11231 GND.n7673 GND.n7670 19.3944
R11232 GND.n7670 GND.n7669 19.3944
R11233 GND.n7669 GND.n7666 19.3944
R11234 GND.n7666 GND.n7665 19.3944
R11235 GND.n7665 GND.n7662 19.3944
R11236 GND.n7660 GND.n7658 19.3944
R11237 GND.n7658 GND.n7655 19.3944
R11238 GND.n7653 GND.n7650 19.3944
R11239 GND.n7650 GND.n7649 19.3944
R11240 GND.n7649 GND.n7646 19.3944
R11241 GND.n7646 GND.n7645 19.3944
R11242 GND.n7641 GND.n7638 19.3944
R11243 GND.n7638 GND.n7637 19.3944
R11244 GND.n7637 GND.n7634 19.3944
R11245 GND.n7634 GND.n7633 19.3944
R11246 GND.n7633 GND.n7630 19.3944
R11247 GND.n7630 GND.n7629 19.3944
R11248 GND.n7629 GND.n7626 19.3944
R11249 GND.n7626 GND.n7625 19.3944
R11250 GND.n7625 GND.n7622 19.3944
R11251 GND.n7620 GND.n7618 19.3944
R11252 GND.n7618 GND.n7615 19.3944
R11253 GND.n7615 GND.n7614 19.3944
R11254 GND.n7614 GND.n7611 19.3944
R11255 GND.n7611 GND.n7610 19.3944
R11256 GND.n7610 GND.n7607 19.3944
R11257 GND.n7607 GND.n7606 19.3944
R11258 GND.n7606 GND.n7603 19.3944
R11259 GND.n7603 GND.n7602 19.3944
R11260 GND.n7712 GND.n664 19.3944
R11261 GND.n7722 GND.n664 19.3944
R11262 GND.n7722 GND.n7721 19.3944
R11263 GND.n7721 GND.n7720 19.3944
R11264 GND.n7720 GND.n644 19.3944
R11265 GND.n7742 GND.n644 19.3944
R11266 GND.n7742 GND.n7741 19.3944
R11267 GND.n7741 GND.n7740 19.3944
R11268 GND.n7740 GND.n624 19.3944
R11269 GND.n7762 GND.n624 19.3944
R11270 GND.n7762 GND.n7761 19.3944
R11271 GND.n7761 GND.n7760 19.3944
R11272 GND.n7760 GND.n604 19.3944
R11273 GND.n7782 GND.n604 19.3944
R11274 GND.n7782 GND.n7781 19.3944
R11275 GND.n7781 GND.n7780 19.3944
R11276 GND.n7780 GND.n583 19.3944
R11277 GND.n7806 GND.n583 19.3944
R11278 GND.n7806 GND.n7805 19.3944
R11279 GND.n7805 GND.n7804 19.3944
R11280 GND.n7804 GND.n7803 19.3944
R11281 GND.n7803 GND.n555 19.3944
R11282 GND.n7880 GND.n555 19.3944
R11283 GND.n7880 GND.n7879 19.3944
R11284 GND.n7879 GND.n7878 19.3944
R11285 GND.n7878 GND.n536 19.3944
R11286 GND.n7900 GND.n536 19.3944
R11287 GND.n7900 GND.n7899 19.3944
R11288 GND.n7899 GND.n7898 19.3944
R11289 GND.n7898 GND.n516 19.3944
R11290 GND.n7920 GND.n516 19.3944
R11291 GND.n7920 GND.n7919 19.3944
R11292 GND.n7919 GND.n7918 19.3944
R11293 GND.n7918 GND.n495 19.3944
R11294 GND.n7947 GND.n495 19.3944
R11295 GND.n7947 GND.n7946 19.3944
R11296 GND.n7946 GND.n7945 19.3944
R11297 GND.n7945 GND.n125 19.3944
R11298 GND.n8598 GND.n125 19.3944
R11299 GND.n8598 GND.n8597 19.3944
R11300 GND.n8597 GND.n8596 19.3944
R11301 GND.n8596 GND.n95 19.3944
R11302 GND.n8628 GND.n95 19.3944
R11303 GND.n8628 GND.n8627 19.3944
R11304 GND.n8627 GND.n8626 19.3944
R11305 GND.n8626 GND.n99 19.3944
R11306 GND.n8228 GND.n99 19.3944
R11307 GND.n8229 GND.n8228 19.3944
R11308 GND.n8231 GND.n8229 19.3944
R11309 GND.n8232 GND.n8231 19.3944
R11310 GND.n8232 GND.n146 19.3944
R11311 GND.n8570 GND.n146 19.3944
R11312 GND.n8570 GND.n8569 19.3944
R11313 GND.n8569 GND.n8568 19.3944
R11314 GND.n8568 GND.n150 19.3944
R11315 GND.n8558 GND.n150 19.3944
R11316 GND.n8558 GND.n8557 19.3944
R11317 GND.n8557 GND.n8556 19.3944
R11318 GND.n8556 GND.n170 19.3944
R11319 GND.n8546 GND.n170 19.3944
R11320 GND.n8546 GND.n8545 19.3944
R11321 GND.n8545 GND.n8544 19.3944
R11322 GND.n8544 GND.n190 19.3944
R11323 GND.n8534 GND.n190 19.3944
R11324 GND.n8534 GND.n8533 19.3944
R11325 GND.n8533 GND.n8532 19.3944
R11326 GND.n8532 GND.n212 19.3944
R11327 GND.n8522 GND.n212 19.3944
R11328 GND.n8522 GND.n8521 19.3944
R11329 GND.n8521 GND.n8520 19.3944
R11330 GND.n8520 GND.n233 19.3944
R11331 GND.n8510 GND.n233 19.3944
R11332 GND.n8510 GND.n8509 19.3944
R11333 GND.n8509 GND.n8508 19.3944
R11334 GND.n8508 GND.n254 19.3944
R11335 GND.n8498 GND.n254 19.3944
R11336 GND.n8498 GND.n8497 19.3944
R11337 GND.n8497 GND.n8496 19.3944
R11338 GND.n8496 GND.n275 19.3944
R11339 GND.n8486 GND.n275 19.3944
R11340 GND.n8486 GND.n8485 19.3944
R11341 GND.n8485 GND.n8484 19.3944
R11342 GND.n8484 GND.n296 19.3944
R11343 GND.n8474 GND.n296 19.3944
R11344 GND.n8474 GND.n8473 19.3944
R11345 GND.n8473 GND.n8472 19.3944
R11346 GND.n8472 GND.n317 19.3944
R11347 GND.n8462 GND.n317 19.3944
R11348 GND.n8462 GND.n8461 19.3944
R11349 GND.n8461 GND.n8460 19.3944
R11350 GND.n8460 GND.n338 19.3944
R11351 GND.n8308 GND.n338 19.3944
R11352 GND.n8309 GND.n8308 19.3944
R11353 GND.n8310 GND.n8309 19.3944
R11354 GND.n8310 GND.n447 19.3944
R11355 GND.n8330 GND.n447 19.3944
R11356 GND.n7715 GND.n666 19.3944
R11357 GND.n7716 GND.n7715 19.3944
R11358 GND.n7717 GND.n7716 19.3944
R11359 GND.n7717 GND.n646 19.3944
R11360 GND.n7735 GND.n646 19.3944
R11361 GND.n7736 GND.n7735 19.3944
R11362 GND.n7737 GND.n7736 19.3944
R11363 GND.n7737 GND.n626 19.3944
R11364 GND.n7755 GND.n626 19.3944
R11365 GND.n7756 GND.n7755 19.3944
R11366 GND.n7757 GND.n7756 19.3944
R11367 GND.n7757 GND.n606 19.3944
R11368 GND.n7775 GND.n606 19.3944
R11369 GND.n7776 GND.n7775 19.3944
R11370 GND.n7777 GND.n7776 19.3944
R11371 GND.n7777 GND.n586 19.3944
R11372 GND.n7795 GND.n586 19.3944
R11373 GND.n7796 GND.n7795 19.3944
R11374 GND.n7798 GND.n7796 19.3944
R11375 GND.n7799 GND.n7798 19.3944
R11376 GND.n7799 GND.n557 19.3944
R11377 GND.n7873 GND.n557 19.3944
R11378 GND.n7874 GND.n7873 19.3944
R11379 GND.n7875 GND.n7874 19.3944
R11380 GND.n7875 GND.n538 19.3944
R11381 GND.n7893 GND.n538 19.3944
R11382 GND.n7894 GND.n7893 19.3944
R11383 GND.n7895 GND.n7894 19.3944
R11384 GND.n7895 GND.n518 19.3944
R11385 GND.n7913 GND.n518 19.3944
R11386 GND.n7914 GND.n7913 19.3944
R11387 GND.n7915 GND.n7914 19.3944
R11388 GND.n7915 GND.n498 19.3944
R11389 GND.n7933 GND.n498 19.3944
R11390 GND.n7934 GND.n7933 19.3944
R11391 GND.n7936 GND.n7934 19.3944
R11392 GND.n7937 GND.n7936 19.3944
R11393 GND.n7942 GND.n7937 19.3944
R11394 GND.n7942 GND.n7940 19.3944
R11395 GND.n7940 GND.n7939 19.3944
R11396 GND.n7939 GND.n128 19.3944
R11397 GND.n8593 GND.n128 19.3944
R11398 GND.n8593 GND.n8591 19.3944
R11399 GND.n8591 GND.n8590 19.3944
R11400 GND.n8590 GND.n8588 19.3944
R11401 GND.n8588 GND.n8587 19.3944
R11402 GND.n8587 GND.n8584 19.3944
R11403 GND.n8584 GND.n8583 19.3944
R11404 GND.n8583 GND.n8582 19.3944
R11405 GND.n8582 GND.n133 19.3944
R11406 GND.n8235 GND.n133 19.3944
R11407 GND.n8236 GND.n8235 19.3944
R11408 GND.n8238 GND.n8236 19.3944
R11409 GND.n8239 GND.n8238 19.3944
R11410 GND.n8242 GND.n8239 19.3944
R11411 GND.n8243 GND.n8242 19.3944
R11412 GND.n8245 GND.n8243 19.3944
R11413 GND.n8246 GND.n8245 19.3944
R11414 GND.n8249 GND.n8246 19.3944
R11415 GND.n8250 GND.n8249 19.3944
R11416 GND.n8252 GND.n8250 19.3944
R11417 GND.n8253 GND.n8252 19.3944
R11418 GND.n8256 GND.n8253 19.3944
R11419 GND.n8257 GND.n8256 19.3944
R11420 GND.n8259 GND.n8257 19.3944
R11421 GND.n8260 GND.n8259 19.3944
R11422 GND.n8263 GND.n8260 19.3944
R11423 GND.n8264 GND.n8263 19.3944
R11424 GND.n8266 GND.n8264 19.3944
R11425 GND.n8267 GND.n8266 19.3944
R11426 GND.n8270 GND.n8267 19.3944
R11427 GND.n8271 GND.n8270 19.3944
R11428 GND.n8273 GND.n8271 19.3944
R11429 GND.n8274 GND.n8273 19.3944
R11430 GND.n8277 GND.n8274 19.3944
R11431 GND.n8278 GND.n8277 19.3944
R11432 GND.n8280 GND.n8278 19.3944
R11433 GND.n8281 GND.n8280 19.3944
R11434 GND.n8284 GND.n8281 19.3944
R11435 GND.n8285 GND.n8284 19.3944
R11436 GND.n8287 GND.n8285 19.3944
R11437 GND.n8288 GND.n8287 19.3944
R11438 GND.n8291 GND.n8288 19.3944
R11439 GND.n8292 GND.n8291 19.3944
R11440 GND.n8294 GND.n8292 19.3944
R11441 GND.n8295 GND.n8294 19.3944
R11442 GND.n8298 GND.n8295 19.3944
R11443 GND.n8299 GND.n8298 19.3944
R11444 GND.n8301 GND.n8299 19.3944
R11445 GND.n8302 GND.n8301 19.3944
R11446 GND.n8304 GND.n8302 19.3944
R11447 GND.n8304 GND.n8225 19.3944
R11448 GND.n8314 GND.n8225 19.3944
R11449 GND.n8314 GND.n8313 19.3944
R11450 GND.n8313 GND.n8312 19.3944
R11451 GND.n8312 GND.n446 19.3944
R11452 GND.n8354 GND.n428 19.3944
R11453 GND.n8354 GND.n8351 19.3944
R11454 GND.n8351 GND.n8350 19.3944
R11455 GND.n8350 GND.n8347 19.3944
R11456 GND.n8347 GND.n8346 19.3944
R11457 GND.n8346 GND.n8343 19.3944
R11458 GND.n8343 GND.n8342 19.3944
R11459 GND.n8342 GND.n8339 19.3944
R11460 GND.n8339 GND.n8338 19.3944
R11461 GND.n8377 GND.n417 19.3944
R11462 GND.n8377 GND.n8374 19.3944
R11463 GND.n8374 GND.n8371 19.3944
R11464 GND.n8371 GND.n8370 19.3944
R11465 GND.n8370 GND.n8367 19.3944
R11466 GND.n8367 GND.n8366 19.3944
R11467 GND.n8366 GND.n8363 19.3944
R11468 GND.n8363 GND.n8362 19.3944
R11469 GND.n8362 GND.n8359 19.3944
R11470 GND.n8400 GND.n404 19.3944
R11471 GND.n8400 GND.n8397 19.3944
R11472 GND.n8397 GND.n8396 19.3944
R11473 GND.n8396 GND.n8393 19.3944
R11474 GND.n8393 GND.n8392 19.3944
R11475 GND.n8392 GND.n8389 19.3944
R11476 GND.n8389 GND.n8388 19.3944
R11477 GND.n8388 GND.n8385 19.3944
R11478 GND.n8385 GND.n8384 19.3944
R11479 GND.n8423 GND.n393 19.3944
R11480 GND.n8423 GND.n8420 19.3944
R11481 GND.n8420 GND.n8417 19.3944
R11482 GND.n8417 GND.n8416 19.3944
R11483 GND.n8416 GND.n8413 19.3944
R11484 GND.n8413 GND.n8412 19.3944
R11485 GND.n8412 GND.n8409 19.3944
R11486 GND.n8409 GND.n8408 19.3944
R11487 GND.n8408 GND.n8405 19.3944
R11488 GND.n8446 GND.n8445 19.3944
R11489 GND.n8445 GND.n387 19.3944
R11490 GND.n8441 GND.n387 19.3944
R11491 GND.n8441 GND.n8438 19.3944
R11492 GND.n8438 GND.n8435 19.3944
R11493 GND.n8435 GND.n8434 19.3944
R11494 GND.n8434 GND.n8431 19.3944
R11495 GND.n8431 GND.n8430 19.3944
R11496 GND.n8192 GND.n8190 19.3944
R11497 GND.n8195 GND.n8192 19.3944
R11498 GND.n8198 GND.n8195 19.3944
R11499 GND.n8201 GND.n8198 19.3944
R11500 GND.n8201 GND.n8188 19.3944
R11501 GND.n8205 GND.n8188 19.3944
R11502 GND.n8208 GND.n8205 19.3944
R11503 GND.n8211 GND.n8208 19.3944
R11504 GND.n1272 GND.n1271 19.3944
R11505 GND.n1271 GND.n1270 19.3944
R11506 GND.n1270 GND.n1269 19.3944
R11507 GND.n1269 GND.n1267 19.3944
R11508 GND.n1267 GND.n1266 19.3944
R11509 GND.n1266 GND.n1264 19.3944
R11510 GND.n1264 GND.n1263 19.3944
R11511 GND.n1263 GND.n1261 19.3944
R11512 GND.n1261 GND.n1260 19.3944
R11513 GND.n1260 GND.n1258 19.3944
R11514 GND.n1258 GND.n1257 19.3944
R11515 GND.n1257 GND.n1255 19.3944
R11516 GND.n1255 GND.n1254 19.3944
R11517 GND.n1254 GND.n1252 19.3944
R11518 GND.n1252 GND.n1251 19.3944
R11519 GND.n1251 GND.n1249 19.3944
R11520 GND.n1249 GND.n1248 19.3944
R11521 GND.n1248 GND.n1246 19.3944
R11522 GND.n1246 GND.n565 19.3944
R11523 GND.n7820 GND.n565 19.3944
R11524 GND.n7820 GND.n563 19.3944
R11525 GND.n7869 GND.n563 19.3944
R11526 GND.n7869 GND.n7868 19.3944
R11527 GND.n7868 GND.n7867 19.3944
R11528 GND.n7867 GND.n7865 19.3944
R11529 GND.n7865 GND.n7864 19.3944
R11530 GND.n7864 GND.n7862 19.3944
R11531 GND.n7862 GND.n7861 19.3944
R11532 GND.n7861 GND.n7859 19.3944
R11533 GND.n7859 GND.n7858 19.3944
R11534 GND.n7858 GND.n7856 19.3944
R11535 GND.n7856 GND.n7855 19.3944
R11536 GND.n7855 GND.n7853 19.3944
R11537 GND.n7853 GND.n7852 19.3944
R11538 GND.n7852 GND.n7850 19.3944
R11539 GND.n7850 GND.n7849 19.3944
R11540 GND.n7849 GND.n7847 19.3944
R11541 GND.n7847 GND.n7846 19.3944
R11542 GND.n7846 GND.n7844 19.3944
R11543 GND.n7844 GND.n7843 19.3944
R11544 GND.n7843 GND.n108 19.3944
R11545 GND.n8611 GND.n108 19.3944
R11546 GND.n8612 GND.n8611 19.3944
R11547 GND.n8612 GND.n106 19.3944
R11548 GND.n8618 GND.n106 19.3944
R11549 GND.n8618 GND.n8617 19.3944
R11550 GND.n8617 GND.n64 19.3944
R11551 GND.n8638 GND.n64 19.3944
R11552 GND.n8638 GND.n65 19.3944
R11553 GND.n8095 GND.n65 19.3944
R11554 GND.n8097 GND.n8095 19.3944
R11555 GND.n8097 GND.n8093 19.3944
R11556 GND.n8102 GND.n8093 19.3944
R11557 GND.n8103 GND.n8102 19.3944
R11558 GND.n8105 GND.n8103 19.3944
R11559 GND.n8105 GND.n8091 19.3944
R11560 GND.n8110 GND.n8091 19.3944
R11561 GND.n8111 GND.n8110 19.3944
R11562 GND.n8113 GND.n8111 19.3944
R11563 GND.n8113 GND.n8089 19.3944
R11564 GND.n8118 GND.n8089 19.3944
R11565 GND.n8119 GND.n8118 19.3944
R11566 GND.n8121 GND.n8119 19.3944
R11567 GND.n8121 GND.n8087 19.3944
R11568 GND.n8126 GND.n8087 19.3944
R11569 GND.n8127 GND.n8126 19.3944
R11570 GND.n8129 GND.n8127 19.3944
R11571 GND.n8129 GND.n8085 19.3944
R11572 GND.n8134 GND.n8085 19.3944
R11573 GND.n8135 GND.n8134 19.3944
R11574 GND.n8137 GND.n8135 19.3944
R11575 GND.n8137 GND.n8083 19.3944
R11576 GND.n8142 GND.n8083 19.3944
R11577 GND.n8143 GND.n8142 19.3944
R11578 GND.n8145 GND.n8143 19.3944
R11579 GND.n8145 GND.n8081 19.3944
R11580 GND.n8150 GND.n8081 19.3944
R11581 GND.n8151 GND.n8150 19.3944
R11582 GND.n8153 GND.n8151 19.3944
R11583 GND.n8153 GND.n8079 19.3944
R11584 GND.n8158 GND.n8079 19.3944
R11585 GND.n8159 GND.n8158 19.3944
R11586 GND.n8161 GND.n8159 19.3944
R11587 GND.n8161 GND.n8077 19.3944
R11588 GND.n8166 GND.n8077 19.3944
R11589 GND.n8167 GND.n8166 19.3944
R11590 GND.n8169 GND.n8167 19.3944
R11591 GND.n8169 GND.n8075 19.3944
R11592 GND.n8174 GND.n8075 19.3944
R11593 GND.n8175 GND.n8174 19.3944
R11594 GND.n8177 GND.n8175 19.3944
R11595 GND.n8177 GND.n8073 19.3944
R11596 GND.n8221 GND.n8073 19.3944
R11597 GND.n8221 GND.n8220 19.3944
R11598 GND.n8220 GND.n8219 19.3944
R11599 GND.n8219 GND.n8218 19.3944
R11600 GND.n6378 GND.n1612 19.3944
R11601 GND.n6378 GND.n1610 19.3944
R11602 GND.n6405 GND.n1610 19.3944
R11603 GND.n6405 GND.n6404 19.3944
R11604 GND.n6404 GND.n6403 19.3944
R11605 GND.n6403 GND.n6402 19.3944
R11606 GND.n6402 GND.n6401 19.3944
R11607 GND.n6401 GND.n6399 19.3944
R11608 GND.n6399 GND.n6398 19.3944
R11609 GND.n6398 GND.n6388 19.3944
R11610 GND.n6394 GND.n6388 19.3944
R11611 GND.n6394 GND.n6393 19.3944
R11612 GND.n6393 GND.n1500 19.3944
R11613 GND.n6555 GND.n1500 19.3944
R11614 GND.n6556 GND.n6555 19.3944
R11615 GND.n6556 GND.n1498 19.3944
R11616 GND.n6571 GND.n1498 19.3944
R11617 GND.n6571 GND.n6570 19.3944
R11618 GND.n6570 GND.n6569 19.3944
R11619 GND.n6569 GND.n6567 19.3944
R11620 GND.n6567 GND.n6566 19.3944
R11621 GND.n6566 GND.n1433 19.3944
R11622 GND.n1433 GND.n1431 19.3944
R11623 GND.n6649 GND.n1431 19.3944
R11624 GND.n6650 GND.n6649 19.3944
R11625 GND.n6650 GND.n1429 19.3944
R11626 GND.n6654 GND.n1429 19.3944
R11627 GND.n6656 GND.n6654 19.3944
R11628 GND.n6657 GND.n6656 19.3944
R11629 GND.n6657 GND.n1426 19.3944
R11630 GND.n6663 GND.n1426 19.3944
R11631 GND.n6663 GND.n6662 19.3944
R11632 GND.n6662 GND.n1358 19.3944
R11633 GND.n6792 GND.n1358 19.3944
R11634 GND.n6792 GND.n1356 19.3944
R11635 GND.n6819 GND.n1356 19.3944
R11636 GND.n6819 GND.n6818 19.3944
R11637 GND.n6818 GND.n6817 19.3944
R11638 GND.n6817 GND.n6816 19.3944
R11639 GND.n6816 GND.n6815 19.3944
R11640 GND.n6815 GND.n6800 19.3944
R11641 GND.n6811 GND.n6800 19.3944
R11642 GND.n6811 GND.n6810 19.3944
R11643 GND.n6810 GND.n6809 19.3944
R11644 GND.n6809 GND.n1288 19.3944
R11645 GND.n6927 GND.n1288 19.3944
R11646 GND.n6928 GND.n6927 19.3944
R11647 GND.n6313 GND.n1569 19.3944
R11648 GND.n6451 GND.n1569 19.3944
R11649 GND.n6451 GND.n1567 19.3944
R11650 GND.n6455 GND.n1567 19.3944
R11651 GND.n6455 GND.n1542 19.3944
R11652 GND.n6484 GND.n1542 19.3944
R11653 GND.n6484 GND.n1540 19.3944
R11654 GND.n6493 GND.n1540 19.3944
R11655 GND.n6493 GND.n6492 19.3944
R11656 GND.n6492 GND.n6491 19.3944
R11657 GND.n6491 GND.n1506 19.3944
R11658 GND.n6547 GND.n1506 19.3944
R11659 GND.n6547 GND.n1504 19.3944
R11660 GND.n6551 GND.n1504 19.3944
R11661 GND.n6551 GND.n1480 19.3944
R11662 GND.n6599 GND.n1480 19.3944
R11663 GND.n6599 GND.n1478 19.3944
R11664 GND.n6603 GND.n1478 19.3944
R11665 GND.n6603 GND.n1440 19.3944
R11666 GND.n6637 GND.n1440 19.3944
R11667 GND.n6637 GND.n1438 19.3944
R11668 GND.n6643 GND.n1438 19.3944
R11669 GND.n6643 GND.n6642 19.3944
R11670 GND.n6642 GND.n1409 19.3944
R11671 GND.n6696 GND.n1409 19.3944
R11672 GND.n6696 GND.n1407 19.3944
R11673 GND.n6702 GND.n1407 19.3944
R11674 GND.n6702 GND.n6701 19.3944
R11675 GND.n6701 GND.n1378 19.3944
R11676 GND.n6764 GND.n1378 19.3944
R11677 GND.n6764 GND.n1376 19.3944
R11678 GND.n6770 GND.n1376 19.3944
R11679 GND.n6770 GND.n6769 19.3944
R11680 GND.n6769 GND.n1347 19.3944
R11681 GND.n6831 GND.n1347 19.3944
R11682 GND.n6831 GND.n1345 19.3944
R11683 GND.n6838 GND.n1345 19.3944
R11684 GND.n6838 GND.n6837 19.3944
R11685 GND.n6837 GND.n1328 19.3944
R11686 GND.n1328 GND.n1326 19.3944
R11687 GND.n6861 GND.n1326 19.3944
R11688 GND.n6861 GND.n1324 19.3944
R11689 GND.n6870 GND.n1324 19.3944
R11690 GND.n6870 GND.n6869 19.3944
R11691 GND.n6869 GND.n6868 19.3944
R11692 GND.n6868 GND.n1178 19.3944
R11693 GND.n6982 GND.n1178 19.3944
R11694 GND.n6318 GND.n6311 19.3944
R11695 GND.n6318 GND.n6309 19.3944
R11696 GND.n6322 GND.n6309 19.3944
R11697 GND.n6322 GND.n6307 19.3944
R11698 GND.n6328 GND.n6307 19.3944
R11699 GND.n6328 GND.n6305 19.3944
R11700 GND.n6333 GND.n6305 19.3944
R11701 GND.n6333 GND.n6302 19.3944
R11702 GND.n6339 GND.n6302 19.3944
R11703 GND.n6340 GND.n6339 19.3944
R11704 GND.n6341 GND.n6340 19.3944
R11705 GND.n6346 GND.n6345 19.3944
R11706 GND.n6351 GND.n6350 19.3944
R11707 GND.n6356 GND.n6355 19.3944
R11708 GND.n6361 GND.n6360 19.3944
R11709 GND.n6372 GND.n1615 19.3944
R11710 GND.n6372 GND.n1613 19.3944
R11711 GND.n6936 GND.n1284 19.3944
R11712 GND.n6931 GND.n1284 19.3944
R11713 GND.n6979 GND.n6978 19.3944
R11714 GND.n6978 GND.n1181 19.3944
R11715 GND.n1182 GND.n1181 19.3944
R11716 GND.n6971 GND.n1182 19.3944
R11717 GND.n6971 GND.n6970 19.3944
R11718 GND.n6970 GND.n6969 19.3944
R11719 GND.n6969 GND.n1189 19.3944
R11720 GND.n6964 GND.n1189 19.3944
R11721 GND.n6964 GND.n6963 19.3944
R11722 GND.n6963 GND.n6962 19.3944
R11723 GND.n6962 GND.n1196 19.3944
R11724 GND.n6957 GND.n6956 19.3944
R11725 GND.n6956 GND.n6955 19.3944
R11726 GND.n6950 GND.n1278 19.3944
R11727 GND.n6948 GND.n6947 19.3944
R11728 GND.n6942 GND.n1282 19.3944
R11729 GND.n1226 GND.n1224 19.3944
R11730 GND.n1221 GND.n1220 19.3944
R11731 GND.n1217 GND.n1216 19.3944
R11732 GND.n1213 GND.n1212 19.3944
R11733 GND.n804 GND.n803 19.3944
R11734 GND.n803 GND.n801 19.3944
R11735 GND.n801 GND.n800 19.3944
R11736 GND.n800 GND.n798 19.3944
R11737 GND.n798 GND.n797 19.3944
R11738 GND.n797 GND.n795 19.3944
R11739 GND.n795 GND.n794 19.3944
R11740 GND.n794 GND.n792 19.3944
R11741 GND.n792 GND.n791 19.3944
R11742 GND.n791 GND.n789 19.3944
R11743 GND.n789 GND.n788 19.3944
R11744 GND.n788 GND.n786 19.3944
R11745 GND.n786 GND.n785 19.3944
R11746 GND.n785 GND.n783 19.3944
R11747 GND.n783 GND.n782 19.3944
R11748 GND.n782 GND.n780 19.3944
R11749 GND.n780 GND.n779 19.3944
R11750 GND.n779 GND.n777 19.3944
R11751 GND.n777 GND.n776 19.3944
R11752 GND.n776 GND.n774 19.3944
R11753 GND.n774 GND.n773 19.3944
R11754 GND.n773 GND.n771 19.3944
R11755 GND.n771 GND.n770 19.3944
R11756 GND.n770 GND.n769 19.3944
R11757 GND.n769 GND.n767 19.3944
R11758 GND.n767 GND.n766 19.3944
R11759 GND.n766 GND.n764 19.3944
R11760 GND.n764 GND.n763 19.3944
R11761 GND.n763 GND.n761 19.3944
R11762 GND.n761 GND.n760 19.3944
R11763 GND.n760 GND.n758 19.3944
R11764 GND.n758 GND.n757 19.3944
R11765 GND.n757 GND.n755 19.3944
R11766 GND.n755 GND.n754 19.3944
R11767 GND.n754 GND.n752 19.3944
R11768 GND.n752 GND.n751 19.3944
R11769 GND.n751 GND.n477 19.3944
R11770 GND.n7960 GND.n477 19.3944
R11771 GND.n7961 GND.n7960 19.3944
R11772 GND.n7963 GND.n7961 19.3944
R11773 GND.n7963 GND.n475 19.3944
R11774 GND.n7968 GND.n475 19.3944
R11775 GND.n7969 GND.n7968 19.3944
R11776 GND.n7973 GND.n7972 19.3944
R11777 GND.n7978 GND.n7975 19.3944
R11778 GND.n7982 GND.n7980 19.3944
R11779 GND.n7986 GND.n7984 19.3944
R11780 GND.n7990 GND.n7988 19.3944
R11781 GND.n7991 GND.n7990 19.3944
R11782 GND.n7995 GND.n7991 19.3944
R11783 GND.n7996 GND.n7995 19.3944
R11784 GND.n7998 GND.n7996 19.3944
R11785 GND.n7998 GND.n473 19.3944
R11786 GND.n8003 GND.n473 19.3944
R11787 GND.n8004 GND.n8003 19.3944
R11788 GND.n8006 GND.n8004 19.3944
R11789 GND.n8006 GND.n471 19.3944
R11790 GND.n8011 GND.n471 19.3944
R11791 GND.n8012 GND.n8011 19.3944
R11792 GND.n8014 GND.n8012 19.3944
R11793 GND.n8014 GND.n469 19.3944
R11794 GND.n8019 GND.n469 19.3944
R11795 GND.n8020 GND.n8019 19.3944
R11796 GND.n8022 GND.n8020 19.3944
R11797 GND.n8022 GND.n467 19.3944
R11798 GND.n8027 GND.n467 19.3944
R11799 GND.n8028 GND.n8027 19.3944
R11800 GND.n8030 GND.n8028 19.3944
R11801 GND.n8030 GND.n465 19.3944
R11802 GND.n8035 GND.n465 19.3944
R11803 GND.n8036 GND.n8035 19.3944
R11804 GND.n8038 GND.n8036 19.3944
R11805 GND.n8038 GND.n463 19.3944
R11806 GND.n8043 GND.n463 19.3944
R11807 GND.n8044 GND.n8043 19.3944
R11808 GND.n8046 GND.n8044 19.3944
R11809 GND.n8046 GND.n461 19.3944
R11810 GND.n8051 GND.n461 19.3944
R11811 GND.n8052 GND.n8051 19.3944
R11812 GND.n8054 GND.n8052 19.3944
R11813 GND.n8054 GND.n459 19.3944
R11814 GND.n8059 GND.n459 19.3944
R11815 GND.n8060 GND.n8059 19.3944
R11816 GND.n8062 GND.n8060 19.3944
R11817 GND.n8062 GND.n457 19.3944
R11818 GND.n8066 GND.n457 19.3944
R11819 GND.n8066 GND.n456 19.3944
R11820 GND.n8318 GND.n456 19.3944
R11821 GND.n8318 GND.n454 19.3944
R11822 GND.n8324 GND.n454 19.3944
R11823 GND.n8324 GND.n8323 19.3944
R11824 GND.n2972 GND.n2971 19.3944
R11825 GND.n2971 GND.n2970 19.3944
R11826 GND.n2970 GND.n2969 19.3944
R11827 GND.n2969 GND.n2967 19.3944
R11828 GND.n2967 GND.n2964 19.3944
R11829 GND.n2964 GND.n2963 19.3944
R11830 GND.n2963 GND.n2960 19.3944
R11831 GND.n2960 GND.n2959 19.3944
R11832 GND.n2955 GND.n2952 19.3944
R11833 GND.n2952 GND.n2951 19.3944
R11834 GND.n2951 GND.n2948 19.3944
R11835 GND.n2948 GND.n2947 19.3944
R11836 GND.n2947 GND.n2944 19.3944
R11837 GND.n2944 GND.n2943 19.3944
R11838 GND.n2943 GND.n2940 19.3944
R11839 GND.n2940 GND.n2939 19.3944
R11840 GND.n2939 GND.n2936 19.3944
R11841 GND.n2934 GND.n2932 19.3944
R11842 GND.n2932 GND.n2929 19.3944
R11843 GND.n2929 GND.n2928 19.3944
R11844 GND.n2928 GND.n2925 19.3944
R11845 GND.n2925 GND.n2924 19.3944
R11846 GND.n2924 GND.n2921 19.3944
R11847 GND.n2921 GND.n2920 19.3944
R11848 GND.n2920 GND.n2917 19.3944
R11849 GND.n2917 GND.n2916 19.3944
R11850 GND.n2912 GND.n2909 19.3944
R11851 GND.n2909 GND.n2908 19.3944
R11852 GND.n2908 GND.n2905 19.3944
R11853 GND.n2905 GND.n2904 19.3944
R11854 GND.n2904 GND.n2901 19.3944
R11855 GND.n2901 GND.n2900 19.3944
R11856 GND.n2900 GND.n2897 19.3944
R11857 GND.n2897 GND.n2896 19.3944
R11858 GND.n2896 GND.n2893 19.3944
R11859 GND.n2891 GND.n2889 19.3944
R11860 GND.n2889 GND.n2886 19.3944
R11861 GND.n2886 GND.n2885 19.3944
R11862 GND.n2885 GND.n2882 19.3944
R11863 GND.n2882 GND.n2881 19.3944
R11864 GND.n2881 GND.n2878 19.3944
R11865 GND.n2878 GND.n2877 19.3944
R11866 GND.n2877 GND.n2874 19.3944
R11867 GND.n2874 GND.n2873 19.3944
R11868 GND.n2570 GND.n2569 19.3944
R11869 GND.n2615 GND.n2570 19.3944
R11870 GND.n2615 GND.n2566 19.3944
R11871 GND.n2714 GND.n2566 19.3944
R11872 GND.n2714 GND.n2713 19.3944
R11873 GND.n2713 GND.n2712 19.3944
R11874 GND.n2712 GND.n2711 19.3944
R11875 GND.n2711 GND.n2710 19.3944
R11876 GND.n2710 GND.n2708 19.3944
R11877 GND.n2708 GND.n2707 19.3944
R11878 GND.n2707 GND.n2705 19.3944
R11879 GND.n2705 GND.n2704 19.3944
R11880 GND.n2704 GND.n2702 19.3944
R11881 GND.n2702 GND.n2701 19.3944
R11882 GND.n2701 GND.n2699 19.3944
R11883 GND.n2699 GND.n2698 19.3944
R11884 GND.n2698 GND.n2696 19.3944
R11885 GND.n2696 GND.n2695 19.3944
R11886 GND.n2695 GND.n2693 19.3944
R11887 GND.n2693 GND.n2692 19.3944
R11888 GND.n2692 GND.n2690 19.3944
R11889 GND.n2690 GND.n2689 19.3944
R11890 GND.n2689 GND.n2687 19.3944
R11891 GND.n2687 GND.n2686 19.3944
R11892 GND.n2686 GND.n2684 19.3944
R11893 GND.n2684 GND.n2683 19.3944
R11894 GND.n2683 GND.n2681 19.3944
R11895 GND.n2681 GND.n2680 19.3944
R11896 GND.n2680 GND.n2678 19.3944
R11897 GND.n2678 GND.n2677 19.3944
R11898 GND.n2677 GND.n2675 19.3944
R11899 GND.n2675 GND.n2674 19.3944
R11900 GND.n2674 GND.n2672 19.3944
R11901 GND.n2672 GND.n2671 19.3944
R11902 GND.n2671 GND.n2669 19.3944
R11903 GND.n2669 GND.n2668 19.3944
R11904 GND.n2668 GND.n2666 19.3944
R11905 GND.n2666 GND.n2665 19.3944
R11906 GND.n2665 GND.n2663 19.3944
R11907 GND.n2663 GND.n2662 19.3944
R11908 GND.n2662 GND.n2660 19.3944
R11909 GND.n2660 GND.n2659 19.3944
R11910 GND.n2659 GND.n2656 19.3944
R11911 GND.n2244 GND.n2243 19.3944
R11912 GND.n2230 GND.n2229 19.3944
R11913 GND.n2221 GND.n2220 19.3944
R11914 GND.n2207 GND.n2206 19.3944
R11915 GND.n5084 GND.n2092 19.3944
R11916 GND.n5084 GND.n2196 19.3944
R11917 GND.n2196 GND.n2195 19.3944
R11918 GND.n2195 GND.n2193 19.3944
R11919 GND.n2193 GND.n2192 19.3944
R11920 GND.n2192 GND.n2190 19.3944
R11921 GND.n2190 GND.n2189 19.3944
R11922 GND.n2189 GND.n2187 19.3944
R11923 GND.n2187 GND.n2186 19.3944
R11924 GND.n2186 GND.n2185 19.3944
R11925 GND.n2185 GND.n2183 19.3944
R11926 GND.n2183 GND.n2182 19.3944
R11927 GND.n2182 GND.n2180 19.3944
R11928 GND.n2180 GND.n2179 19.3944
R11929 GND.n2179 GND.n2177 19.3944
R11930 GND.n2177 GND.n2176 19.3944
R11931 GND.n2176 GND.n2174 19.3944
R11932 GND.n2174 GND.n2173 19.3944
R11933 GND.n2173 GND.n2171 19.3944
R11934 GND.n2171 GND.n2170 19.3944
R11935 GND.n2170 GND.n2168 19.3944
R11936 GND.n2168 GND.n2167 19.3944
R11937 GND.n2167 GND.n2165 19.3944
R11938 GND.n2165 GND.n2164 19.3944
R11939 GND.n2164 GND.n2162 19.3944
R11940 GND.n2162 GND.n2161 19.3944
R11941 GND.n2161 GND.n2159 19.3944
R11942 GND.n2159 GND.n2158 19.3944
R11943 GND.n2158 GND.n2156 19.3944
R11944 GND.n2156 GND.n2155 19.3944
R11945 GND.n2155 GND.n2153 19.3944
R11946 GND.n2153 GND.n2152 19.3944
R11947 GND.n2152 GND.n2150 19.3944
R11948 GND.n2150 GND.n2149 19.3944
R11949 GND.n2149 GND.n2147 19.3944
R11950 GND.n2147 GND.n2146 19.3944
R11951 GND.n2146 GND.n2144 19.3944
R11952 GND.n2144 GND.n2143 19.3944
R11953 GND.n2143 GND.n2142 19.3944
R11954 GND.n2142 GND.n2140 19.3944
R11955 GND.n2140 GND.n2139 19.3944
R11956 GND.n2139 GND.n2137 19.3944
R11957 GND.n2137 GND.n2136 19.3944
R11958 GND.n2136 GND.n2134 19.3944
R11959 GND.n4850 GND.n2428 19.3944
R11960 GND.n4850 GND.n2411 19.3944
R11961 GND.n4866 GND.n2411 19.3944
R11962 GND.n4866 GND.n2409 19.3944
R11963 GND.n4870 GND.n2409 19.3944
R11964 GND.n4870 GND.n2391 19.3944
R11965 GND.n4886 GND.n2391 19.3944
R11966 GND.n4886 GND.n2389 19.3944
R11967 GND.n4890 GND.n2389 19.3944
R11968 GND.n4890 GND.n2371 19.3944
R11969 GND.n4906 GND.n2371 19.3944
R11970 GND.n4906 GND.n2369 19.3944
R11971 GND.n4910 GND.n2369 19.3944
R11972 GND.n4910 GND.n2350 19.3944
R11973 GND.n4926 GND.n2350 19.3944
R11974 GND.n4926 GND.n2348 19.3944
R11975 GND.n4930 GND.n2348 19.3944
R11976 GND.n4930 GND.n2331 19.3944
R11977 GND.n4946 GND.n2331 19.3944
R11978 GND.n4946 GND.n2329 19.3944
R11979 GND.n4950 GND.n2329 19.3944
R11980 GND.n4950 GND.n2311 19.3944
R11981 GND.n4966 GND.n2311 19.3944
R11982 GND.n4966 GND.n2309 19.3944
R11983 GND.n4970 GND.n2309 19.3944
R11984 GND.n4970 GND.n2291 19.3944
R11985 GND.n4986 GND.n2291 19.3944
R11986 GND.n4986 GND.n2289 19.3944
R11987 GND.n4990 GND.n2289 19.3944
R11988 GND.n4990 GND.n2271 19.3944
R11989 GND.n5006 GND.n2271 19.3944
R11990 GND.n5006 GND.n2269 19.3944
R11991 GND.n5011 GND.n2269 19.3944
R11992 GND.n5011 GND.n2249 19.3944
R11993 GND.n5032 GND.n2249 19.3944
R11994 GND.n5033 GND.n5032 19.3944
R11995 GND.n5034 GND.n5033 19.3944
R11996 GND.n5036 GND.n2084 19.3944
R11997 GND.n2226 GND.n2084 19.3944
R11998 GND.n5054 GND.n5053 19.3944
R11999 GND.n2204 GND.n2203 19.3944
R12000 GND.n5079 GND.n5078 19.3944
R12001 GND.n5088 GND.n2077 19.3944
R12002 GND.n5088 GND.n2059 19.3944
R12003 GND.n5109 GND.n2059 19.3944
R12004 GND.n5109 GND.n2057 19.3944
R12005 GND.n5115 GND.n2057 19.3944
R12006 GND.n5115 GND.n5114 19.3944
R12007 GND.n5114 GND.n2032 19.3944
R12008 GND.n5200 GND.n2032 19.3944
R12009 GND.n5200 GND.n2030 19.3944
R12010 GND.n5204 GND.n2030 19.3944
R12011 GND.n5204 GND.n2012 19.3944
R12012 GND.n5220 GND.n2012 19.3944
R12013 GND.n5220 GND.n2010 19.3944
R12014 GND.n5224 GND.n2010 19.3944
R12015 GND.n5224 GND.n1992 19.3944
R12016 GND.n5240 GND.n1992 19.3944
R12017 GND.n5240 GND.n1990 19.3944
R12018 GND.n5244 GND.n1990 19.3944
R12019 GND.n5244 GND.n1972 19.3944
R12020 GND.n5260 GND.n1972 19.3944
R12021 GND.n5260 GND.n1970 19.3944
R12022 GND.n5264 GND.n1970 19.3944
R12023 GND.n5264 GND.n1952 19.3944
R12024 GND.n5280 GND.n1952 19.3944
R12025 GND.n5280 GND.n1950 19.3944
R12026 GND.n5284 GND.n1950 19.3944
R12027 GND.n5284 GND.n1932 19.3944
R12028 GND.n5300 GND.n1932 19.3944
R12029 GND.n5300 GND.n1930 19.3944
R12030 GND.n5304 GND.n1930 19.3944
R12031 GND.n5304 GND.n1912 19.3944
R12032 GND.n5325 GND.n1912 19.3944
R12033 GND.n5325 GND.n1910 19.3944
R12034 GND.n5331 GND.n1910 19.3944
R12035 GND.n5331 GND.n5330 19.3944
R12036 GND.n5330 GND.n1885 19.3944
R12037 GND.n5370 GND.n1885 19.3944
R12038 GND.n5370 GND.n1883 19.3944
R12039 GND.n5376 GND.n1883 19.3944
R12040 GND.n5376 GND.n5375 19.3944
R12041 GND.n5375 GND.n1867 19.3944
R12042 GND.n5390 GND.n1867 19.3944
R12043 GND.n5390 GND.n1865 19.3944
R12044 GND.n5394 GND.n1865 19.3944
R12045 GND.n5394 GND.n1864 19.3944
R12046 GND.n5398 GND.n1864 19.3944
R12047 GND.n5398 GND.n1862 19.3944
R12048 GND.n5402 GND.n1862 19.3944
R12049 GND.n5402 GND.n1860 19.3944
R12050 GND.n5408 GND.n1860 19.3944
R12051 GND.n5408 GND.n1858 19.3944
R12052 GND.n6188 GND.n1858 19.3944
R12053 GND.n6188 GND.n6187 19.3944
R12054 GND.n6187 GND.n6186 19.3944
R12055 GND.n6186 GND.n5414 19.3944
R12056 GND.n6174 GND.n5414 19.3944
R12057 GND.n6174 GND.n6173 19.3944
R12058 GND.n6173 GND.n6172 19.3944
R12059 GND.n6172 GND.n5432 19.3944
R12060 GND.n5522 GND.n5432 19.3944
R12061 GND.n6155 GND.n5522 19.3944
R12062 GND.n6155 GND.n6154 19.3944
R12063 GND.n6154 GND.n6153 19.3944
R12064 GND.n6153 GND.n5528 19.3944
R12065 GND.n6141 GND.n5528 19.3944
R12066 GND.n6141 GND.n6140 19.3944
R12067 GND.n6140 GND.n6139 19.3944
R12068 GND.n6139 GND.n5546 19.3944
R12069 GND.n6127 GND.n5546 19.3944
R12070 GND.n6127 GND.n6126 19.3944
R12071 GND.n6126 GND.n6125 19.3944
R12072 GND.n6125 GND.n5564 19.3944
R12073 GND.n6113 GND.n5564 19.3944
R12074 GND.n6113 GND.n6112 19.3944
R12075 GND.n6112 GND.n6111 19.3944
R12076 GND.n6111 GND.n5582 19.3944
R12077 GND.n5653 GND.n5582 19.3944
R12078 GND.n6094 GND.n5653 19.3944
R12079 GND.n6094 GND.n6093 19.3944
R12080 GND.n6093 GND.n6092 19.3944
R12081 GND.n6092 GND.n5659 19.3944
R12082 GND.n6080 GND.n5659 19.3944
R12083 GND.n6080 GND.n6079 19.3944
R12084 GND.n6079 GND.n6078 19.3944
R12085 GND.n6078 GND.n5677 19.3944
R12086 GND.n6066 GND.n5677 19.3944
R12087 GND.n6066 GND.n6065 19.3944
R12088 GND.n6065 GND.n6064 19.3944
R12089 GND.n6064 GND.n5695 19.3944
R12090 GND.n6052 GND.n5695 19.3944
R12091 GND.n6052 GND.n6051 19.3944
R12092 GND.n6051 GND.n6050 19.3944
R12093 GND.n6050 GND.n5713 19.3944
R12094 GND.n5784 GND.n5713 19.3944
R12095 GND.n6033 GND.n5784 19.3944
R12096 GND.n6033 GND.n6032 19.3944
R12097 GND.n6032 GND.n6031 19.3944
R12098 GND.n6031 GND.n5790 19.3944
R12099 GND.n6019 GND.n5790 19.3944
R12100 GND.n6019 GND.n6018 19.3944
R12101 GND.n6018 GND.n6017 19.3944
R12102 GND.n6017 GND.n5807 19.3944
R12103 GND.n6005 GND.n5807 19.3944
R12104 GND.n6005 GND.n6004 19.3944
R12105 GND.n6004 GND.n6003 19.3944
R12106 GND.n6003 GND.n5825 19.3944
R12107 GND.n5991 GND.n5825 19.3944
R12108 GND.n5991 GND.n5990 19.3944
R12109 GND.n5990 GND.n5989 19.3944
R12110 GND.n5989 GND.n5843 19.3944
R12111 GND.n5915 GND.n5843 19.3944
R12112 GND.n5972 GND.n5915 19.3944
R12113 GND.n5972 GND.n5971 19.3944
R12114 GND.n5971 GND.n5970 19.3944
R12115 GND.n5970 GND.n5921 19.3944
R12116 GND.n5958 GND.n5921 19.3944
R12117 GND.n5958 GND.n5957 19.3944
R12118 GND.n5957 GND.n1584 19.3944
R12119 GND.n6433 GND.n1584 19.3944
R12120 GND.n6433 GND.n1582 19.3944
R12121 GND.n6439 GND.n1582 19.3944
R12122 GND.n6439 GND.n6438 19.3944
R12123 GND.n6438 GND.n1553 19.3944
R12124 GND.n6470 GND.n1553 19.3944
R12125 GND.n6470 GND.n1551 19.3944
R12126 GND.n6479 GND.n1551 19.3944
R12127 GND.n6479 GND.n6478 19.3944
R12128 GND.n6478 GND.n6477 19.3944
R12129 GND.n6477 GND.n1515 19.3944
R12130 GND.n6530 GND.n1515 19.3944
R12131 GND.n6530 GND.n1513 19.3944
R12132 GND.n6542 GND.n1513 19.3944
R12133 GND.n6542 GND.n6541 19.3944
R12134 GND.n6541 GND.n6540 19.3944
R12135 GND.n6540 GND.n6537 19.3944
R12136 GND.n6537 GND.n1472 19.3944
R12137 GND.n6608 GND.n1472 19.3944
R12138 GND.n6608 GND.n1470 19.3944
R12139 GND.n6617 GND.n1470 19.3944
R12140 GND.n6617 GND.n6616 19.3944
R12141 GND.n6616 GND.n6615 19.3944
R12142 GND.n6615 GND.n1417 19.3944
R12143 GND.n6687 GND.n1417 19.3944
R12144 GND.n6687 GND.n1415 19.3944
R12145 GND.n6691 GND.n1415 19.3944
R12146 GND.n6691 GND.n1394 19.3944
R12147 GND.n6716 GND.n1394 19.3944
R12148 GND.n6716 GND.n1392 19.3944
R12149 GND.n6751 GND.n1392 19.3944
R12150 GND.n6751 GND.n6750 19.3944
R12151 GND.n6750 GND.n6749 19.3944
R12152 GND.n6749 GND.n6722 19.3944
R12153 GND.n6744 GND.n6722 19.3944
R12154 GND.n6744 GND.n6743 19.3944
R12155 GND.n6743 GND.n6742 19.3944
R12156 GND.n6742 GND.n6728 19.3944
R12157 GND.n6737 GND.n6728 19.3944
R12158 GND.n6737 GND.n6736 19.3944
R12159 GND.n6736 GND.n6735 19.3944
R12160 GND.n6735 GND.n1306 19.3944
R12161 GND.n6889 GND.n1306 19.3944
R12162 GND.n6889 GND.n1304 19.3944
R12163 GND.n6907 GND.n1304 19.3944
R12164 GND.n6907 GND.n6906 19.3944
R12165 GND.n6906 GND.n6905 19.3944
R12166 GND.n6905 GND.n6895 19.3944
R12167 GND.n6901 GND.n6895 19.3944
R12168 GND.n6901 GND.n6900 19.3944
R12169 GND.n6900 GND.n1153 19.3944
R12170 GND.n7012 GND.n1153 19.3944
R12171 GND.n7012 GND.n1151 19.3944
R12172 GND.n7024 GND.n1151 19.3944
R12173 GND.n7024 GND.n7023 19.3944
R12174 GND.n7023 GND.n7022 19.3944
R12175 GND.n7022 GND.n7019 19.3944
R12176 GND.n7019 GND.n1122 19.3944
R12177 GND.n7058 GND.n1122 19.3944
R12178 GND.n7058 GND.n1120 19.3944
R12179 GND.n7073 GND.n1120 19.3944
R12180 GND.n7073 GND.n7072 19.3944
R12181 GND.n7072 GND.n7071 19.3944
R12182 GND.n7071 GND.n7064 19.3944
R12183 GND.n7067 GND.n7064 19.3944
R12184 GND.n7067 GND.n1088 19.3944
R12185 GND.n7116 GND.n1088 19.3944
R12186 GND.n7116 GND.n1086 19.3944
R12187 GND.n7122 GND.n1086 19.3944
R12188 GND.n7122 GND.n7121 19.3944
R12189 GND.n7121 GND.n1063 19.3944
R12190 GND.n7151 GND.n1063 19.3944
R12191 GND.n7151 GND.n1061 19.3944
R12192 GND.n7160 GND.n1061 19.3944
R12193 GND.n7160 GND.n7159 19.3944
R12194 GND.n7159 GND.n7158 19.3944
R12195 GND.n7158 GND.n1039 19.3944
R12196 GND.n7190 GND.n1039 19.3944
R12197 GND.n7190 GND.n1037 19.3944
R12198 GND.n7205 GND.n1037 19.3944
R12199 GND.n7205 GND.n7204 19.3944
R12200 GND.n7204 GND.n7203 19.3944
R12201 GND.n7203 GND.n7196 19.3944
R12202 GND.n7199 GND.n7196 19.3944
R12203 GND.n7199 GND.n1005 19.3944
R12204 GND.n7248 GND.n1005 19.3944
R12205 GND.n7248 GND.n1003 19.3944
R12206 GND.n7254 GND.n1003 19.3944
R12207 GND.n7254 GND.n7253 19.3944
R12208 GND.n7253 GND.n980 19.3944
R12209 GND.n7283 GND.n980 19.3944
R12210 GND.n7283 GND.n978 19.3944
R12211 GND.n7292 GND.n978 19.3944
R12212 GND.n7292 GND.n7291 19.3944
R12213 GND.n7291 GND.n7290 19.3944
R12214 GND.n7290 GND.n955 19.3944
R12215 GND.n7321 GND.n955 19.3944
R12216 GND.n7321 GND.n953 19.3944
R12217 GND.n7327 GND.n953 19.3944
R12218 GND.n7327 GND.n7326 19.3944
R12219 GND.n7326 GND.n930 19.3944
R12220 GND.n7356 GND.n930 19.3944
R12221 GND.n7356 GND.n928 19.3944
R12222 GND.n7360 GND.n928 19.3944
R12223 GND.n7360 GND.n913 19.3944
R12224 GND.n7380 GND.n913 19.3944
R12225 GND.n7380 GND.n911 19.3944
R12226 GND.n7386 GND.n911 19.3944
R12227 GND.n7386 GND.n7385 19.3944
R12228 GND.n7385 GND.n890 19.3944
R12229 GND.n7416 GND.n890 19.3944
R12230 GND.n7416 GND.n888 19.3944
R12231 GND.n7420 GND.n888 19.3944
R12232 GND.n7420 GND.n873 19.3944
R12233 GND.n7486 GND.n873 19.3944
R12234 GND.n7486 GND.n871 19.3944
R12235 GND.n7503 GND.n871 19.3944
R12236 GND.n7503 GND.n7502 19.3944
R12237 GND.n7502 GND.n7501 19.3944
R12238 GND.n7501 GND.n7492 19.3944
R12239 GND.n7495 GND.n7492 19.3944
R12240 GND.n7495 GND.n677 19.3944
R12241 GND.n7704 GND.n677 19.3944
R12242 GND.n7704 GND.n675 19.3944
R12243 GND.n7708 GND.n675 19.3944
R12244 GND.n7708 GND.n656 19.3944
R12245 GND.n7726 GND.n656 19.3944
R12246 GND.n7726 GND.n654 19.3944
R12247 GND.n7730 GND.n654 19.3944
R12248 GND.n7730 GND.n636 19.3944
R12249 GND.n7746 GND.n636 19.3944
R12250 GND.n7746 GND.n634 19.3944
R12251 GND.n7750 GND.n634 19.3944
R12252 GND.n7750 GND.n616 19.3944
R12253 GND.n7766 GND.n616 19.3944
R12254 GND.n7766 GND.n614 19.3944
R12255 GND.n7770 GND.n614 19.3944
R12256 GND.n7770 GND.n596 19.3944
R12257 GND.n7786 GND.n596 19.3944
R12258 GND.n7786 GND.n594 19.3944
R12259 GND.n7790 GND.n594 19.3944
R12260 GND.n7790 GND.n575 19.3944
R12261 GND.n7810 GND.n575 19.3944
R12262 GND.n7810 GND.n573 19.3944
R12263 GND.n7816 GND.n573 19.3944
R12264 GND.n7816 GND.n7815 19.3944
R12265 GND.n7815 GND.n548 19.3944
R12266 GND.n7884 GND.n548 19.3944
R12267 GND.n7884 GND.n546 19.3944
R12268 GND.n7888 GND.n546 19.3944
R12269 GND.n7888 GND.n528 19.3944
R12270 GND.n7904 GND.n528 19.3944
R12271 GND.n7904 GND.n526 19.3944
R12272 GND.n7908 GND.n526 19.3944
R12273 GND.n7908 GND.n508 19.3944
R12274 GND.n7924 GND.n508 19.3944
R12275 GND.n7924 GND.n506 19.3944
R12276 GND.n7928 GND.n506 19.3944
R12277 GND.n7928 GND.n487 19.3944
R12278 GND.n7951 GND.n487 19.3944
R12279 GND.n7951 GND.n485 19.3944
R12280 GND.n7955 GND.n485 19.3944
R12281 GND.n7955 GND.n117 19.3944
R12282 GND.n8602 GND.n117 19.3944
R12283 GND.n8602 GND.n115 19.3944
R12284 GND.n8606 GND.n115 19.3944
R12285 GND.n8606 GND.n84 19.3944
R12286 GND.n8632 GND.n84 19.3944
R12287 GND.n8632 GND.n85 19.3944
R12288 GND.n8622 GND.n8621 19.3944
R12289 GND.n8635 GND.n75 19.3944
R12290 GND.n8577 GND.n76 19.3944
R12291 GND.n8575 GND.n8574 19.3944
R12292 GND.n8564 GND.n157 19.3944
R12293 GND.n8564 GND.n8563 19.3944
R12294 GND.n8563 GND.n8562 19.3944
R12295 GND.n8562 GND.n160 19.3944
R12296 GND.n8552 GND.n160 19.3944
R12297 GND.n8552 GND.n8551 19.3944
R12298 GND.n8551 GND.n8550 19.3944
R12299 GND.n8550 GND.n181 19.3944
R12300 GND.n8540 GND.n181 19.3944
R12301 GND.n8540 GND.n8539 19.3944
R12302 GND.n8539 GND.n8538 19.3944
R12303 GND.n8538 GND.n202 19.3944
R12304 GND.n8528 GND.n202 19.3944
R12305 GND.n8528 GND.n8527 19.3944
R12306 GND.n8527 GND.n8526 19.3944
R12307 GND.n8526 GND.n223 19.3944
R12308 GND.n8516 GND.n223 19.3944
R12309 GND.n8516 GND.n8515 19.3944
R12310 GND.n8515 GND.n8514 19.3944
R12311 GND.n8514 GND.n244 19.3944
R12312 GND.n8504 GND.n244 19.3944
R12313 GND.n8504 GND.n8503 19.3944
R12314 GND.n8503 GND.n8502 19.3944
R12315 GND.n8502 GND.n265 19.3944
R12316 GND.n8492 GND.n265 19.3944
R12317 GND.n8492 GND.n8491 19.3944
R12318 GND.n8491 GND.n8490 19.3944
R12319 GND.n8490 GND.n286 19.3944
R12320 GND.n8480 GND.n286 19.3944
R12321 GND.n8480 GND.n8479 19.3944
R12322 GND.n8479 GND.n8478 19.3944
R12323 GND.n8478 GND.n307 19.3944
R12324 GND.n8468 GND.n307 19.3944
R12325 GND.n8468 GND.n8467 19.3944
R12326 GND.n8467 GND.n8466 19.3944
R12327 GND.n8466 GND.n328 19.3944
R12328 GND.n8456 GND.n328 19.3944
R12329 GND.n4728 GND.n3021 19.3944
R12330 GND.n4734 GND.n3021 19.3944
R12331 GND.n4734 GND.n3019 19.3944
R12332 GND.n4738 GND.n3019 19.3944
R12333 GND.n4738 GND.n3017 19.3944
R12334 GND.n4744 GND.n3017 19.3944
R12335 GND.n4744 GND.n3015 19.3944
R12336 GND.n4748 GND.n3015 19.3944
R12337 GND.n4748 GND.n3013 19.3944
R12338 GND.n4754 GND.n3013 19.3944
R12339 GND.n4754 GND.n3011 19.3944
R12340 GND.n4758 GND.n3011 19.3944
R12341 GND.n4758 GND.n3009 19.3944
R12342 GND.n4764 GND.n3009 19.3944
R12343 GND.n4764 GND.n3007 19.3944
R12344 GND.n4768 GND.n3007 19.3944
R12345 GND.n4768 GND.n3005 19.3944
R12346 GND.n4774 GND.n3005 19.3944
R12347 GND.n4774 GND.n3003 19.3944
R12348 GND.n4778 GND.n3003 19.3944
R12349 GND.n4778 GND.n3001 19.3944
R12350 GND.n4784 GND.n3001 19.3944
R12351 GND.n4784 GND.n2999 19.3944
R12352 GND.n4788 GND.n2999 19.3944
R12353 GND.n4788 GND.n2997 19.3944
R12354 GND.n4794 GND.n2997 19.3944
R12355 GND.n4794 GND.n2995 19.3944
R12356 GND.n4798 GND.n2995 19.3944
R12357 GND.n4798 GND.n2993 19.3944
R12358 GND.n4804 GND.n2993 19.3944
R12359 GND.n4804 GND.n2991 19.3944
R12360 GND.n4808 GND.n2991 19.3944
R12361 GND.n4808 GND.n2989 19.3944
R12362 GND.n4814 GND.n2989 19.3944
R12363 GND.n4814 GND.n2987 19.3944
R12364 GND.n4818 GND.n2987 19.3944
R12365 GND.n4818 GND.n2985 19.3944
R12366 GND.n4824 GND.n2985 19.3944
R12367 GND.n4824 GND.n2983 19.3944
R12368 GND.n4828 GND.n2983 19.3944
R12369 GND.n4828 GND.n2981 19.3944
R12370 GND.n4834 GND.n2981 19.3944
R12371 GND.n4834 GND.n2979 19.3944
R12372 GND.n4839 GND.n2979 19.3944
R12373 GND.n4839 GND.n2977 19.3944
R12374 GND.n2977 GND.n2430 19.3944
R12375 GND.n4846 GND.n2430 19.3944
R12376 GND.n2862 GND.n2861 19.3944
R12377 GND.n2861 GND.n2537 19.3944
R12378 GND.n2546 GND.n2537 19.3944
R12379 GND.n2547 GND.n2546 19.3944
R12380 GND.n2548 GND.n2547 19.3944
R12381 GND.n2549 GND.n2548 19.3944
R12382 GND.n2549 GND.n2422 19.3944
R12383 GND.n4855 GND.n2422 19.3944
R12384 GND.n4856 GND.n4855 19.3944
R12385 GND.n4857 GND.n4856 19.3944
R12386 GND.n4857 GND.n2402 19.3944
R12387 GND.n4875 GND.n2402 19.3944
R12388 GND.n4876 GND.n4875 19.3944
R12389 GND.n4877 GND.n4876 19.3944
R12390 GND.n4877 GND.n2382 19.3944
R12391 GND.n4895 GND.n2382 19.3944
R12392 GND.n4896 GND.n4895 19.3944
R12393 GND.n4897 GND.n4896 19.3944
R12394 GND.n4897 GND.n2362 19.3944
R12395 GND.n4915 GND.n2362 19.3944
R12396 GND.n4916 GND.n4915 19.3944
R12397 GND.n4917 GND.n4916 19.3944
R12398 GND.n4917 GND.n2342 19.3944
R12399 GND.n4935 GND.n2342 19.3944
R12400 GND.n4936 GND.n4935 19.3944
R12401 GND.n4937 GND.n4936 19.3944
R12402 GND.n4937 GND.n2322 19.3944
R12403 GND.n4955 GND.n2322 19.3944
R12404 GND.n4956 GND.n4955 19.3944
R12405 GND.n4957 GND.n4956 19.3944
R12406 GND.n4957 GND.n2302 19.3944
R12407 GND.n4975 GND.n2302 19.3944
R12408 GND.n4976 GND.n4975 19.3944
R12409 GND.n4977 GND.n4976 19.3944
R12410 GND.n4977 GND.n2282 19.3944
R12411 GND.n4995 GND.n2282 19.3944
R12412 GND.n4996 GND.n4995 19.3944
R12413 GND.n4997 GND.n4996 19.3944
R12414 GND.n4997 GND.n2262 19.3944
R12415 GND.n5016 GND.n2262 19.3944
R12416 GND.n5017 GND.n5016 19.3944
R12417 GND.n5019 GND.n5017 19.3944
R12418 GND.n5020 GND.n5019 19.3944
R12419 GND.n5020 GND.n2239 19.3944
R12420 GND.n5041 GND.n2239 19.3944
R12421 GND.n5042 GND.n5041 19.3944
R12422 GND.n5043 GND.n5042 19.3944
R12423 GND.n5043 GND.n2216 19.3944
R12424 GND.n5058 GND.n2216 19.3944
R12425 GND.n5059 GND.n5058 19.3944
R12426 GND.n5061 GND.n5059 19.3944
R12427 GND.n5062 GND.n5061 19.3944
R12428 GND.n5063 GND.n5062 19.3944
R12429 GND.n5063 GND.n2070 19.3944
R12430 GND.n5093 GND.n2070 19.3944
R12431 GND.n5094 GND.n5093 19.3944
R12432 GND.n5096 GND.n5094 19.3944
R12433 GND.n5097 GND.n5096 19.3944
R12434 GND.n5097 GND.n2042 19.3944
R12435 GND.n5189 GND.n2042 19.3944
R12436 GND.n5190 GND.n5189 19.3944
R12437 GND.n5191 GND.n5190 19.3944
R12438 GND.n5191 GND.n2023 19.3944
R12439 GND.n5209 GND.n2023 19.3944
R12440 GND.n5210 GND.n5209 19.3944
R12441 GND.n5211 GND.n5210 19.3944
R12442 GND.n5211 GND.n2003 19.3944
R12443 GND.n5229 GND.n2003 19.3944
R12444 GND.n5230 GND.n5229 19.3944
R12445 GND.n5231 GND.n5230 19.3944
R12446 GND.n5231 GND.n1983 19.3944
R12447 GND.n5249 GND.n1983 19.3944
R12448 GND.n5250 GND.n5249 19.3944
R12449 GND.n5251 GND.n5250 19.3944
R12450 GND.n5251 GND.n1963 19.3944
R12451 GND.n5269 GND.n1963 19.3944
R12452 GND.n5270 GND.n5269 19.3944
R12453 GND.n5271 GND.n5270 19.3944
R12454 GND.n5271 GND.n1943 19.3944
R12455 GND.n5289 GND.n1943 19.3944
R12456 GND.n5290 GND.n5289 19.3944
R12457 GND.n5291 GND.n5290 19.3944
R12458 GND.n5291 GND.n1923 19.3944
R12459 GND.n5309 GND.n1923 19.3944
R12460 GND.n5310 GND.n5309 19.3944
R12461 GND.n5312 GND.n5310 19.3944
R12462 GND.n5313 GND.n5312 19.3944
R12463 GND.n5313 GND.n1895 19.3944
R12464 GND.n5359 GND.n1895 19.3944
R12465 GND.n5360 GND.n5359 19.3944
R12466 GND.n5361 GND.n5360 19.3944
R12467 GND.n5361 GND.n1876 19.3944
R12468 GND.n5381 GND.n1876 19.3944
R12469 GND.n5383 GND.n5381 19.3944
R12470 GND.n5383 GND.n5382 19.3944
R12471 GND.n5382 GND.n1626 19.3944
R12472 GND.n1639 GND.n1638 19.3944
R12473 GND.n1644 GND.n1643 19.3944
R12474 GND.n1649 GND.n1648 19.3944
R12475 GND.n1652 GND.n1622 19.3944
R12476 GND.n5975 GND.t1 19.0848
R12477 GND.n7040 GND.t0 19.0848
R12478 GND.n4 GND.t77 19.039
R12479 GND.n4 GND.t69 19.039
R12480 GND.n6 GND.t18 19.039
R12481 GND.n6 GND.t29 19.039
R12482 GND.n8 GND.t78 19.039
R12483 GND.n8 GND.t70 19.039
R12484 GND.n10 GND.t16 19.039
R12485 GND.n10 GND.t28 19.039
R12486 GND.n13 GND.t76 19.039
R12487 GND.n13 GND.t68 19.039
R12488 GND.n15 GND.t17 19.039
R12489 GND.n15 GND.t27 19.039
R12490 GND.n18 GND.t62 19.039
R12491 GND.n18 GND.t31 19.039
R12492 GND.n20 GND.t61 19.039
R12493 GND.n20 GND.t20 19.039
R12494 GND.n23 GND.t35 19.039
R12495 GND.n23 GND.t66 19.039
R12496 GND.n25 GND.t73 19.039
R12497 GND.n25 GND.t74 19.039
R12498 GND.n0 GND.t63 19.039
R12499 GND.n0 GND.t37 19.039
R12500 GND.n2 GND.t40 19.039
R12501 GND.n2 GND.t41 19.039
R12502 GND.n34 GND.t71 19.039
R12503 GND.n34 GND.t39 19.039
R12504 GND.n33 GND.t14 19.039
R12505 GND.n33 GND.t60 19.039
R12506 GND.n38 GND.t64 19.039
R12507 GND.n38 GND.t38 19.039
R12508 GND.n37 GND.t13 19.039
R12509 GND.n37 GND.t57 19.039
R12510 GND.n43 GND.t65 19.039
R12511 GND.n43 GND.t36 19.039
R12512 GND.n42 GND.t12 19.039
R12513 GND.n42 GND.t56 19.039
R12514 GND.n48 GND.t67 19.039
R12515 GND.n48 GND.t24 19.039
R12516 GND.n47 GND.t53 19.039
R12517 GND.n47 GND.t45 19.039
R12518 GND.n53 GND.t26 19.039
R12519 GND.n53 GND.t49 19.039
R12520 GND.n52 GND.t42 19.039
R12521 GND.n52 GND.t50 19.039
R12522 GND.n58 GND.t52 19.039
R12523 GND.n58 GND.t79 19.039
R12524 GND.n57 GND.t75 19.039
R12525 GND.n57 GND.t80 19.039
R12526 GND.n6245 GND.n6242 18.6187
R12527 GND.n7655 GND.n7654 18.6187
R12528 GND.n4932 GND.t15 18.378
R12529 GND.n5258 GND.t32 18.378
R12530 GND.n5607 GND.n5540 18.378
R12531 GND.n6137 GND.n6136 18.378
R12532 GND.n5740 GND.n5671 18.378
R12533 GND.n6076 GND.n6075 18.378
R12534 GND.n5871 GND.n5870 18.378
R12535 GND.n6015 GND.n6014 18.378
R12536 GND.n5952 GND.n5950 18.378
R12537 GND.n6423 GND.n1586 18.378
R12538 GND.n6991 GND.n1168 18.378
R12539 GND.n7002 GND.n1155 18.378
R12540 GND.n7114 GND.n1090 18.378
R12541 GND.n7125 GND.n1082 18.378
R12542 GND.n7227 GND.n1019 18.378
R12543 GND.n7238 GND.n1007 18.378
R12544 GND.n944 GND.n938 18.378
R12545 GND.n7354 GND.n7353 18.378
R12546 GND.n7882 GND.t11 18.378
R12547 GND.t21 GND.n248 18.378
R12548 GND.n6415 GND.n1578 17.6712
R12549 GND.n6407 GND.n1574 17.6712
R12550 GND.n6468 GND.n6467 17.6712
R12551 GND.n6482 GND.n6481 17.6712
R12552 GND.n6481 GND.n1547 17.6712
R12553 GND.n6495 GND.n1537 17.6712
R12554 GND.n6528 GND.n1517 17.6712
R12555 GND.n6545 GND.n6544 17.6712
R12556 GND.n6553 GND.n1490 17.6712
R12557 GND.t84 GND.n1482 17.6712
R12558 GND.n6606 GND.n6605 17.6712
R12559 GND.n6645 GND.n1434 17.6712
R12560 GND.n6685 GND.n1419 17.6712
R12561 GND.n6685 GND.n1421 17.6712
R12562 GND.n6694 GND.n6693 17.6712
R12563 GND.n6754 GND.n6753 17.6712
R12564 GND.t5 GND.n1370 17.6712
R12565 GND.n6746 GND.n1364 17.6712
R12566 GND.n6829 GND.n1349 17.6712
R12567 GND.n6840 GND.n1342 17.6712
R12568 GND.n6857 GND.n1329 17.6712
R12569 GND.n6880 GND.n1314 17.6712
R12570 GND.n6880 GND.n1315 17.6712
R12571 GND.n1320 GND.n1310 17.6712
R12572 GND.n6807 GND.n1294 17.6712
R12573 GND.n6925 GND.n1172 17.6712
R12574 GND.n6635 GND.t186 17.3178
R12575 GND.n6704 GND.t8 17.3178
R12576 GND.n2355 GND.t15 16.9644
R12577 GND.t32 GND.n1965 16.9644
R12578 GND.n6143 GND.n5540 16.9644
R12579 GND.n6136 GND.n5550 16.9644
R12580 GND.n6082 GND.n5671 16.9644
R12581 GND.n6075 GND.n5681 16.9644
R12582 GND.n6014 GND.n5811 16.9644
R12583 GND.n5960 GND.n5950 16.9644
R12584 GND.n5951 GND.n1592 16.9644
R12585 GND.n6431 GND.n1586 16.9644
R12586 GND.n6518 GND.n1502 16.9644
R12587 GND.n6597 GND.n1485 16.9644
R12588 GND.n6665 GND.n1383 16.9644
R12589 GND.n6780 GND.n1365 16.9644
R12590 GND.n6991 GND.n1166 16.9644
R12591 GND.n7003 GND.n1161 16.9644
R12592 GND.n7010 GND.n1155 16.9644
R12593 GND.n7106 GND.n1090 16.9644
R12594 GND.n7227 GND.n1018 16.9644
R12595 GND.n7246 GND.n1007 16.9644
R12596 GND.n945 GND.n944 16.9644
R12597 GND.n7353 GND.n934 16.9644
R12598 GND.n7871 GND.t11 16.9644
R12599 GND.n8506 GND.t21 16.9644
R12600 GND.n6264 GND.n1705 16.2914
R12601 GND.n7682 GND.n7681 16.2914
R12602 GND.n8427 GND.n393 16.2914
R12603 GND.n2956 GND.n2955 16.2914
R12604 GND.n5870 GND.t6 16.2575
R12605 GND.n6457 GND.n1555 16.2575
R12606 GND.n1596 GND.n1530 16.2575
R12607 GND.n6628 GND.n1461 16.2575
R12608 GND.n1413 GND.n1401 16.2575
R12609 GND.n6849 GND.n6848 16.2575
R12610 GND.n6873 GND.n6872 16.2575
R12611 GND.n7125 GND.t7 16.2575
R12612 GND.n6250 GND.n6249 16.0975
R12613 GND.n7661 GND.n7660 16.0975
R12614 GND.n8404 GND.n404 16.0975
R12615 GND.n2935 GND.n2934 16.0975
R12616 GND.n1808 GND.n1738 15.9035
R12617 GND.n7642 GND.n7641 15.9035
R12618 GND.n8381 GND.n417 15.9035
R12619 GND.n2913 GND.n2912 15.9035
R12620 GND.n1794 GND.n1793 15.7096
R12621 GND.n7621 GND.n7620 15.7096
R12622 GND.n8358 GND.n428 15.7096
R12623 GND.n2892 GND.n2891 15.7096
R12624 GND.n5491 GND.n1854 15.5507
R12625 GND.n6151 GND.n6150 15.5507
R12626 GND.n5620 GND.n5558 15.5507
R12627 GND.n6090 GND.n6089 15.5507
R12628 GND.n6029 GND.n6028 15.5507
R12629 GND.n5884 GND.n5819 15.5507
R12630 GND.n5968 GND.n5967 15.5507
R12631 GND.n6442 GND.n6441 15.5507
R12632 GND.n6588 GND.n1476 15.5507
R12633 GND.n6755 GND.n1387 15.5507
R12634 GND.n6924 GND.n1290 15.5507
R12635 GND.n7027 GND.n7026 15.5507
R12636 GND.n7095 GND.n1101 15.5507
R12637 GND.n1077 GND.n1071 15.5507
R12638 GND.n7257 GND.n7256 15.5507
R12639 GND.n7330 GND.n949 15.5507
R12640 GND.n926 GND.n919 15.5507
R12641 GND.n7484 GND.n7483 15.5507
R12642 GND.n1777 GND.n1776 15.5157
R12643 GND.n7599 GND.n7594 15.5157
R12644 GND.n8335 GND.n441 15.5157
R12645 GND.n2870 GND.n2530 15.5157
R12646 GND.n6449 GND.n6448 14.8439
R12647 GND.n6527 GND.n1519 14.8439
R12648 GND.n6620 GND.n1467 14.8439
R12649 GND.n6713 GND.n1397 14.8439
R12650 GND.n6822 GND.n6821 14.8439
R12651 GND.n6917 GND.n1295 14.8439
R12652 GND.t86 GND.n1508 14.4905
R12653 GND.n6828 GND.t82 14.4905
R12654 GND.n2602 GND.n2601 14.352
R12655 GND.n8215 GND.n8186 14.352
R12656 GND.n6183 GND.n5418 14.137
R12657 GND.n6157 GND.n5518 14.137
R12658 GND.n6122 GND.n5568 14.137
R12659 GND.n6096 GND.n5650 14.137
R12660 GND.n6061 GND.n5699 14.137
R12661 GND.n6035 GND.n5781 14.137
R12662 GND.n6000 GND.n5829 14.137
R12663 GND.n5974 GND.n5912 14.137
R12664 GND.n6504 GND.n6503 14.137
R12665 GND.n6634 GND.n1444 14.137
R12666 GND.n6706 GND.n6705 14.137
R12667 GND.n6841 GND.n1337 14.137
R12668 GND.n1142 GND.n1137 14.137
R12669 GND.n1112 GND.n1111 14.137
R12670 GND.n7148 GND.n1067 14.137
R12671 GND.n7208 GND.n1033 14.137
R12672 GND.n994 GND.n988 14.137
R12673 GND.n7311 GND.n957 14.137
R12674 GND.n7377 GND.n907 14.137
R12675 GND.n7422 GND.n886 14.137
R12676 GND.n5641 GND.t10 13.4302
R12677 GND.n6416 GND.n1588 13.4302
R12678 GND.n1525 GND.n1510 13.4302
R12679 GND.n6573 GND.n1474 13.4302
R12680 GND.n6762 GND.n1380 13.4302
R12681 GND.n6790 GND.n6789 13.4302
R12682 GND.n6985 GND.n6984 13.4302
R12683 GND.t85 GND.n974 13.4302
R12684 GND.n5434 GND.n5426 12.7234
R12685 GND.n6164 GND.n5507 12.7234
R12686 GND.n5640 GND.n5576 12.7234
R12687 GND.n6103 GND.n5636 12.7234
R12688 GND.n5715 GND.n5707 12.7234
R12689 GND.n6042 GND.n5769 12.7234
R12690 GND.n5845 GND.n5837 12.7234
R12691 GND.n5981 GND.n5900 12.7234
R12692 GND.n6466 GND.n1558 12.7234
R12693 GND.n6496 GND.n1534 12.7234
R12694 GND.n1457 GND.n1435 12.7234
R12695 GND.n1451 GND.n1411 12.7234
R12696 GND.n6856 GND.n1333 12.7234
R12697 GND.n6887 GND.n6886 12.7234
R12698 GND.n7048 GND.n1132 12.7234
R12699 GND.n7076 GND.n1116 12.7234
R12700 GND.n1058 GND.n1052 12.7234
R12701 GND.n7180 GND.n1041 12.7234
R12702 GND.n7280 GND.n984 12.7234
R12703 GND.n7300 GND.n968 12.7234
R12704 GND.n7396 GND.n903 12.7234
R12705 GND.n7414 GND.n7413 12.7234
R12706 GND.n6164 GND.t147 12.0166
R12707 GND.n6582 GND.n6581 12.0166
R12708 GND.n6581 GND.n6580 12.0166
R12709 GND.n6773 GND.n6772 12.0166
R12710 GND.n6772 GND.n1373 12.0166
R12711 GND.n7396 GND.t106 12.0166
R12712 GND.n2601 GND.n2600 11.6369
R12713 GND.n8211 GND.n8186 11.6369
R12714 GND.n1209 GND.n1208 11.6369
R12715 GND.n1658 GND.n1622 11.6369
R12716 GND.n5435 GND.n5434 11.3097
R12717 GND.n5507 GND.n5437 11.3097
R12718 GND.n5641 GND.n5640 11.3097
R12719 GND.n5636 GND.n5585 11.3097
R12720 GND.n5716 GND.n5715 11.3097
R12721 GND.n5769 GND.n5718 11.3097
R12722 GND.n5846 GND.n5845 11.3097
R12723 GND.n5900 GND.n5848 11.3097
R12724 GND.n1558 GND.n1544 11.3097
R12725 GND.n1600 GND.n1534 11.3097
R12726 GND.n1458 GND.n1457 11.3097
R12727 GND.n1452 GND.n1451 11.3097
R12728 GND.n1333 GND.n1332 11.3097
R12729 GND.n6887 GND.n1308 11.3097
R12730 GND.n1132 GND.n1124 11.3097
R12731 GND.n1126 GND.n1116 11.3097
R12732 GND.n7169 GND.n1052 11.3097
R12733 GND.n7181 GND.n7180 11.3097
R12734 GND.n984 GND.n973 11.3097
R12735 GND.n974 GND.n968 11.3097
R12736 GND.n903 GND.n898 11.3097
R12737 GND.n7414 GND.n892 11.3097
R12738 GND.n7554 GND.n7553 10.6151
R12739 GND.n7553 GND.n7552 10.6151
R12740 GND.n7552 GND.n7549 10.6151
R12741 GND.n7549 GND.n7548 10.6151
R12742 GND.n7548 GND.n7545 10.6151
R12743 GND.n7545 GND.n7544 10.6151
R12744 GND.n7544 GND.n7541 10.6151
R12745 GND.n7541 GND.n7540 10.6151
R12746 GND.n7540 GND.n7537 10.6151
R12747 GND.n7537 GND.n7536 10.6151
R12748 GND.n7536 GND.n7533 10.6151
R12749 GND.n7533 GND.n7532 10.6151
R12750 GND.n7532 GND.n7529 10.6151
R12751 GND.n7529 GND.n7528 10.6151
R12752 GND.n7528 GND.n7525 10.6151
R12753 GND.n7525 GND.n7524 10.6151
R12754 GND.n7524 GND.n7521 10.6151
R12755 GND.n7519 GND.n7516 10.6151
R12756 GND.n7516 GND.n7515 10.6151
R12757 GND.n7515 GND.n835 10.6151
R12758 GND.n7437 GND.n836 10.6151
R12759 GND.n7440 GND.n7437 10.6151
R12760 GND.n7441 GND.n7440 10.6151
R12761 GND.n7445 GND.n7444 10.6151
R12762 GND.n7448 GND.n7445 10.6151
R12763 GND.n7449 GND.n7448 10.6151
R12764 GND.n7452 GND.n7449 10.6151
R12765 GND.n7453 GND.n7452 10.6151
R12766 GND.n7456 GND.n7453 10.6151
R12767 GND.n7457 GND.n7456 10.6151
R12768 GND.n7460 GND.n7457 10.6151
R12769 GND.n7461 GND.n7460 10.6151
R12770 GND.n7464 GND.n7461 10.6151
R12771 GND.n7465 GND.n7464 10.6151
R12772 GND.n7468 GND.n7465 10.6151
R12773 GND.n7469 GND.n7468 10.6151
R12774 GND.n7472 GND.n7469 10.6151
R12775 GND.n7473 GND.n7472 10.6151
R12776 GND.n7476 GND.n7473 10.6151
R12777 GND.n7478 GND.n7476 10.6151
R12778 GND.n5488 GND.n5487 10.6151
R12779 GND.n5489 GND.n5488 10.6151
R12780 GND.n5489 GND.n5440 10.6151
R12781 GND.n5497 GND.n5440 10.6151
R12782 GND.n5498 GND.n5497 10.6151
R12783 GND.n5500 GND.n5498 10.6151
R12784 GND.n5501 GND.n5500 10.6151
R12785 GND.n5503 GND.n5501 10.6151
R12786 GND.n5504 GND.n5503 10.6151
R12787 GND.n6168 GND.n5504 10.6151
R12788 GND.n6168 GND.n6167 10.6151
R12789 GND.n6167 GND.n6166 10.6151
R12790 GND.n6166 GND.n5505 10.6151
R12791 GND.n5591 GND.n5505 10.6151
R12792 GND.n5592 GND.n5591 10.6151
R12793 GND.n5592 GND.n5590 10.6151
R12794 GND.n5600 GND.n5590 10.6151
R12795 GND.n5601 GND.n5600 10.6151
R12796 GND.n5603 GND.n5601 10.6151
R12797 GND.n5604 GND.n5603 10.6151
R12798 GND.n5605 GND.n5604 10.6151
R12799 GND.n5605 GND.n5589 10.6151
R12800 GND.n5613 GND.n5589 10.6151
R12801 GND.n5614 GND.n5613 10.6151
R12802 GND.n5616 GND.n5614 10.6151
R12803 GND.n5617 GND.n5616 10.6151
R12804 GND.n5618 GND.n5617 10.6151
R12805 GND.n5618 GND.n5588 10.6151
R12806 GND.n5626 GND.n5588 10.6151
R12807 GND.n5627 GND.n5626 10.6151
R12808 GND.n5629 GND.n5627 10.6151
R12809 GND.n5630 GND.n5629 10.6151
R12810 GND.n5632 GND.n5630 10.6151
R12811 GND.n5633 GND.n5632 10.6151
R12812 GND.n6107 GND.n5633 10.6151
R12813 GND.n6107 GND.n6106 10.6151
R12814 GND.n6106 GND.n6105 10.6151
R12815 GND.n6105 GND.n5634 10.6151
R12816 GND.n5724 GND.n5634 10.6151
R12817 GND.n5725 GND.n5724 10.6151
R12818 GND.n5725 GND.n5723 10.6151
R12819 GND.n5733 GND.n5723 10.6151
R12820 GND.n5734 GND.n5733 10.6151
R12821 GND.n5736 GND.n5734 10.6151
R12822 GND.n5737 GND.n5736 10.6151
R12823 GND.n5738 GND.n5737 10.6151
R12824 GND.n5738 GND.n5722 10.6151
R12825 GND.n5746 GND.n5722 10.6151
R12826 GND.n5747 GND.n5746 10.6151
R12827 GND.n5749 GND.n5747 10.6151
R12828 GND.n5750 GND.n5749 10.6151
R12829 GND.n5751 GND.n5750 10.6151
R12830 GND.n5751 GND.n5721 10.6151
R12831 GND.n5759 GND.n5721 10.6151
R12832 GND.n5760 GND.n5759 10.6151
R12833 GND.n5762 GND.n5760 10.6151
R12834 GND.n5763 GND.n5762 10.6151
R12835 GND.n5765 GND.n5763 10.6151
R12836 GND.n5766 GND.n5765 10.6151
R12837 GND.n6046 GND.n5766 10.6151
R12838 GND.n6046 GND.n6045 10.6151
R12839 GND.n6045 GND.n6044 10.6151
R12840 GND.n6044 GND.n5767 10.6151
R12841 GND.n5854 GND.n5767 10.6151
R12842 GND.n5855 GND.n5854 10.6151
R12843 GND.n5855 GND.n5853 10.6151
R12844 GND.n5863 GND.n5853 10.6151
R12845 GND.n5864 GND.n5863 10.6151
R12846 GND.n5866 GND.n5864 10.6151
R12847 GND.n5867 GND.n5866 10.6151
R12848 GND.n5868 GND.n5867 10.6151
R12849 GND.n5868 GND.n5852 10.6151
R12850 GND.n5877 GND.n5852 10.6151
R12851 GND.n5878 GND.n5877 10.6151
R12852 GND.n5880 GND.n5878 10.6151
R12853 GND.n5881 GND.n5880 10.6151
R12854 GND.n5882 GND.n5881 10.6151
R12855 GND.n5882 GND.n5851 10.6151
R12856 GND.n5890 GND.n5851 10.6151
R12857 GND.n5891 GND.n5890 10.6151
R12858 GND.n5893 GND.n5891 10.6151
R12859 GND.n5894 GND.n5893 10.6151
R12860 GND.n5896 GND.n5894 10.6151
R12861 GND.n5897 GND.n5896 10.6151
R12862 GND.n5985 GND.n5897 10.6151
R12863 GND.n5985 GND.n5984 10.6151
R12864 GND.n5984 GND.n5983 10.6151
R12865 GND.n5983 GND.n5898 10.6151
R12866 GND.n5934 GND.n5898 10.6151
R12867 GND.n5935 GND.n5934 10.6151
R12868 GND.n5935 GND.n5933 10.6151
R12869 GND.n5943 GND.n5933 10.6151
R12870 GND.n5944 GND.n5943 10.6151
R12871 GND.n5946 GND.n5944 10.6151
R12872 GND.n5947 GND.n5946 10.6151
R12873 GND.n5948 GND.n5947 10.6151
R12874 GND.n5948 GND.n1595 10.6151
R12875 GND.n6421 GND.n1595 10.6151
R12876 GND.n6421 GND.n6420 10.6151
R12877 GND.n6420 GND.n6419 10.6151
R12878 GND.n6419 GND.n6418 10.6151
R12879 GND.n6418 GND.n6414 10.6151
R12880 GND.n6414 GND.n6413 10.6151
R12881 GND.n6413 GND.n6411 10.6151
R12882 GND.n6411 GND.n6410 10.6151
R12883 GND.n6410 GND.n1609 10.6151
R12884 GND.n1609 GND.n1608 10.6151
R12885 GND.n1608 GND.n1606 10.6151
R12886 GND.n1606 GND.n1605 10.6151
R12887 GND.n1605 GND.n1603 10.6151
R12888 GND.n1603 GND.n1602 10.6151
R12889 GND.n1602 GND.n1599 10.6151
R12890 GND.n1599 GND.n1598 10.6151
R12891 GND.n1598 GND.n1528 10.6151
R12892 GND.n6506 GND.n1528 10.6151
R12893 GND.n6507 GND.n6506 10.6151
R12894 GND.n6508 GND.n6507 10.6151
R12895 GND.n6513 GND.n6508 10.6151
R12896 GND.n6514 GND.n6513 10.6151
R12897 GND.n6516 GND.n6514 10.6151
R12898 GND.n6516 GND.n6515 10.6151
R12899 GND.n6515 GND.n1493 10.6151
R12900 GND.n6578 GND.n1493 10.6151
R12901 GND.n6578 GND.n6577 10.6151
R12902 GND.n6577 GND.n6576 10.6151
R12903 GND.n6576 GND.n1494 10.6151
R12904 GND.n1495 GND.n1494 10.6151
R12905 GND.n1495 GND.n1465 10.6151
R12906 GND.n6622 GND.n1465 10.6151
R12907 GND.n6623 GND.n6622 10.6151
R12908 GND.n6624 GND.n6623 10.6151
R12909 GND.n6626 GND.n6624 10.6151
R12910 GND.n6626 GND.n6625 10.6151
R12911 GND.n6625 GND.n1424 10.6151
R12912 GND.n6683 GND.n1424 10.6151
R12913 GND.n6683 GND.n6682 10.6151
R12914 GND.n6682 GND.n6681 10.6151
R12915 GND.n6681 GND.n6678 10.6151
R12916 GND.n6678 GND.n6677 10.6151
R12917 GND.n6677 GND.n6676 10.6151
R12918 GND.n6676 GND.n6675 10.6151
R12919 GND.n6675 GND.n6674 10.6151
R12920 GND.n6674 GND.n6671 10.6151
R12921 GND.n6671 GND.n6670 10.6151
R12922 GND.n6670 GND.n6668 10.6151
R12923 GND.n6668 GND.n6667 10.6151
R12924 GND.n6667 GND.n1425 10.6151
R12925 GND.n1425 GND.n1362 10.6151
R12926 GND.n6782 GND.n1362 10.6151
R12927 GND.n6783 GND.n6782 10.6151
R12928 GND.n6787 GND.n6783 10.6151
R12929 GND.n6787 GND.n6786 10.6151
R12930 GND.n6786 GND.n6785 10.6151
R12931 GND.n6785 GND.n1340 10.6151
R12932 GND.n6843 GND.n1340 10.6151
R12933 GND.n6844 GND.n6843 10.6151
R12934 GND.n6846 GND.n6844 10.6151
R12935 GND.n6846 GND.n6845 10.6151
R12936 GND.n6845 GND.n1318 10.6151
R12937 GND.n6878 GND.n1318 10.6151
R12938 GND.n6878 GND.n6877 10.6151
R12939 GND.n6877 GND.n6876 10.6151
R12940 GND.n6876 GND.n6875 10.6151
R12941 GND.n6875 GND.n1319 10.6151
R12942 GND.n1319 GND.n1292 10.6151
R12943 GND.n6919 GND.n1292 10.6151
R12944 GND.n6920 GND.n6919 10.6151
R12945 GND.n6922 GND.n6920 10.6151
R12946 GND.n6922 GND.n6921 10.6151
R12947 GND.n6921 GND.n1164 10.6151
R12948 GND.n6993 GND.n1164 10.6151
R12949 GND.n6994 GND.n6993 10.6151
R12950 GND.n7000 GND.n6994 10.6151
R12951 GND.n7000 GND.n6999 10.6151
R12952 GND.n6999 GND.n6998 10.6151
R12953 GND.n6998 GND.n6997 10.6151
R12954 GND.n6997 GND.n6995 10.6151
R12955 GND.n6995 GND.n1139 10.6151
R12956 GND.n7035 GND.n1139 10.6151
R12957 GND.n7036 GND.n7035 10.6151
R12958 GND.n7037 GND.n7036 10.6151
R12959 GND.n7037 GND.n1129 10.6151
R12960 GND.n7050 GND.n1129 10.6151
R12961 GND.n7051 GND.n7050 10.6151
R12962 GND.n7054 GND.n7051 10.6151
R12963 GND.n7054 GND.n7053 10.6151
R12964 GND.n7053 GND.n7052 10.6151
R12965 GND.n7052 GND.n1108 10.6151
R12966 GND.n7084 GND.n1108 10.6151
R12967 GND.n7085 GND.n7084 10.6151
R12968 GND.n7086 GND.n7085 10.6151
R12969 GND.n7086 GND.n1099 10.6151
R12970 GND.n7097 GND.n1099 10.6151
R12971 GND.n7098 GND.n7097 10.6151
R12972 GND.n7104 GND.n7098 10.6151
R12973 GND.n7104 GND.n7103 10.6151
R12974 GND.n7103 GND.n7102 10.6151
R12975 GND.n7102 GND.n7101 10.6151
R12976 GND.n7101 GND.n7099 10.6151
R12977 GND.n7099 GND.n1074 10.6151
R12978 GND.n7133 GND.n1074 10.6151
R12979 GND.n7134 GND.n7133 10.6151
R12980 GND.n7140 GND.n7134 10.6151
R12981 GND.n7140 GND.n7139 10.6151
R12982 GND.n7139 GND.n7138 10.6151
R12983 GND.n7138 GND.n7137 10.6151
R12984 GND.n7137 GND.n7135 10.6151
R12985 GND.n7135 GND.n1050 10.6151
R12986 GND.n7171 GND.n1050 10.6151
R12987 GND.n7172 GND.n7171 10.6151
R12988 GND.n7178 GND.n7172 10.6151
R12989 GND.n7178 GND.n7177 10.6151
R12990 GND.n7177 GND.n7176 10.6151
R12991 GND.n7176 GND.n7175 10.6151
R12992 GND.n7175 GND.n7173 10.6151
R12993 GND.n7173 GND.n1025 10.6151
R12994 GND.n7216 GND.n1025 10.6151
R12995 GND.n7217 GND.n7216 10.6151
R12996 GND.n7218 GND.n7217 10.6151
R12997 GND.n7218 GND.n1016 10.6151
R12998 GND.n7229 GND.n1016 10.6151
R12999 GND.n7230 GND.n7229 10.6151
R13000 GND.n7236 GND.n7230 10.6151
R13001 GND.n7236 GND.n7235 10.6151
R13002 GND.n7235 GND.n7234 10.6151
R13003 GND.n7234 GND.n7233 10.6151
R13004 GND.n7233 GND.n7231 10.6151
R13005 GND.n7231 GND.n991 10.6151
R13006 GND.n7265 GND.n991 10.6151
R13007 GND.n7266 GND.n7265 10.6151
R13008 GND.n7272 GND.n7266 10.6151
R13009 GND.n7272 GND.n7271 10.6151
R13010 GND.n7271 GND.n7270 10.6151
R13011 GND.n7270 GND.n7269 10.6151
R13012 GND.n7269 GND.n7267 10.6151
R13013 GND.n7267 GND.n966 10.6151
R13014 GND.n7302 GND.n966 10.6151
R13015 GND.n7303 GND.n7302 10.6151
R13016 GND.n7309 GND.n7303 10.6151
R13017 GND.n7309 GND.n7308 10.6151
R13018 GND.n7308 GND.n7307 10.6151
R13019 GND.n7307 GND.n7306 10.6151
R13020 GND.n7306 GND.n7304 10.6151
R13021 GND.n7304 GND.n941 10.6151
R13022 GND.n7338 GND.n941 10.6151
R13023 GND.n7339 GND.n7338 10.6151
R13024 GND.n7345 GND.n7339 10.6151
R13025 GND.n7345 GND.n7344 10.6151
R13026 GND.n7344 GND.n7343 10.6151
R13027 GND.n7343 GND.n7342 10.6151
R13028 GND.n7342 GND.n7340 10.6151
R13029 GND.n7340 GND.n917 10.6151
R13030 GND.n7372 GND.n917 10.6151
R13031 GND.n7373 GND.n7372 10.6151
R13032 GND.n7375 GND.n7373 10.6151
R13033 GND.n7375 GND.n7374 10.6151
R13034 GND.n7374 GND.n901 10.6151
R13035 GND.n7398 GND.n901 10.6151
R13036 GND.n7399 GND.n7398 10.6151
R13037 GND.n7405 GND.n7399 10.6151
R13038 GND.n7405 GND.n7404 10.6151
R13039 GND.n7404 GND.n7403 10.6151
R13040 GND.n7403 GND.n7402 10.6151
R13041 GND.n7402 GND.n7400 10.6151
R13042 GND.n7400 GND.n877 10.6151
R13043 GND.n7432 GND.n877 10.6151
R13044 GND.n7433 GND.n7432 10.6151
R13045 GND.n7481 GND.n7433 10.6151
R13046 GND.n7481 GND.n7480 10.6151
R13047 GND.n7480 GND.n7479 10.6151
R13048 GND.n5445 GND.n1820 10.6151
R13049 GND.n5446 GND.n5445 10.6151
R13050 GND.n5449 GND.n5446 10.6151
R13051 GND.n5454 GND.n5451 10.6151
R13052 GND.n5455 GND.n5454 10.6151
R13053 GND.n5458 GND.n5455 10.6151
R13054 GND.n5459 GND.n5458 10.6151
R13055 GND.n5462 GND.n5459 10.6151
R13056 GND.n5463 GND.n5462 10.6151
R13057 GND.n5466 GND.n5463 10.6151
R13058 GND.n5467 GND.n5466 10.6151
R13059 GND.n5470 GND.n5467 10.6151
R13060 GND.n5471 GND.n5470 10.6151
R13061 GND.n5474 GND.n5471 10.6151
R13062 GND.n5475 GND.n5474 10.6151
R13063 GND.n5478 GND.n5475 10.6151
R13064 GND.n5479 GND.n5478 10.6151
R13065 GND.n5482 GND.n5479 10.6151
R13066 GND.n5484 GND.n5482 10.6151
R13067 GND.n5485 GND.n5484 10.6151
R13068 GND.n6234 GND.n6233 10.6151
R13069 GND.n6233 GND.n6232 10.6151
R13070 GND.n6232 GND.n6231 10.6151
R13071 GND.n6231 GND.n6229 10.6151
R13072 GND.n6229 GND.n6226 10.6151
R13073 GND.n6226 GND.n6225 10.6151
R13074 GND.n6225 GND.n6222 10.6151
R13075 GND.n6222 GND.n6221 10.6151
R13076 GND.n6221 GND.n6218 10.6151
R13077 GND.n6218 GND.n6217 10.6151
R13078 GND.n6217 GND.n6214 10.6151
R13079 GND.n6214 GND.n6213 10.6151
R13080 GND.n6213 GND.n6210 10.6151
R13081 GND.n6210 GND.n6209 10.6151
R13082 GND.n6209 GND.n6206 10.6151
R13083 GND.n6206 GND.n6205 10.6151
R13084 GND.n6205 GND.n6202 10.6151
R13085 GND.n6200 GND.n6197 10.6151
R13086 GND.n6197 GND.n1822 10.6151
R13087 GND.n6240 GND.n1822 10.6151
R13088 GND.n6194 GND.n6193 10.6151
R13089 GND.n6193 GND.n1850 10.6151
R13090 GND.n5492 GND.n1850 10.6151
R13091 GND.n5492 GND.n5421 10.6151
R13092 GND.n6181 GND.n5421 10.6151
R13093 GND.n6181 GND.n6180 10.6151
R13094 GND.n6180 GND.n6179 10.6151
R13095 GND.n6179 GND.n5422 10.6151
R13096 GND.n5511 GND.n5422 10.6151
R13097 GND.n5512 GND.n5511 10.6151
R13098 GND.n5513 GND.n5512 10.6151
R13099 GND.n6162 GND.n5513 10.6151
R13100 GND.n6162 GND.n6161 10.6151
R13101 GND.n6161 GND.n6160 10.6151
R13102 GND.n6160 GND.n5514 10.6151
R13103 GND.n5595 GND.n5514 10.6151
R13104 GND.n5595 GND.n5535 10.6151
R13105 GND.n6148 GND.n5535 10.6151
R13106 GND.n6148 GND.n6147 10.6151
R13107 GND.n6147 GND.n6146 10.6151
R13108 GND.n6146 GND.n5536 10.6151
R13109 GND.n5608 GND.n5536 10.6151
R13110 GND.n5608 GND.n5553 10.6151
R13111 GND.n6134 GND.n5553 10.6151
R13112 GND.n6134 GND.n6133 10.6151
R13113 GND.n6133 GND.n6132 10.6151
R13114 GND.n6132 GND.n5554 10.6151
R13115 GND.n5621 GND.n5554 10.6151
R13116 GND.n5621 GND.n5571 10.6151
R13117 GND.n6120 GND.n5571 10.6151
R13118 GND.n6120 GND.n6119 10.6151
R13119 GND.n6119 GND.n6118 10.6151
R13120 GND.n6118 GND.n5572 10.6151
R13121 GND.n5643 GND.n5572 10.6151
R13122 GND.n5644 GND.n5643 10.6151
R13123 GND.n5645 GND.n5644 10.6151
R13124 GND.n6101 GND.n5645 10.6151
R13125 GND.n6101 GND.n6100 10.6151
R13126 GND.n6100 GND.n6099 10.6151
R13127 GND.n6099 GND.n5646 10.6151
R13128 GND.n5728 GND.n5646 10.6151
R13129 GND.n5728 GND.n5666 10.6151
R13130 GND.n6087 GND.n5666 10.6151
R13131 GND.n6087 GND.n6086 10.6151
R13132 GND.n6086 GND.n6085 10.6151
R13133 GND.n6085 GND.n5667 10.6151
R13134 GND.n5741 GND.n5667 10.6151
R13135 GND.n5741 GND.n5684 10.6151
R13136 GND.n6073 GND.n5684 10.6151
R13137 GND.n6073 GND.n6072 10.6151
R13138 GND.n6072 GND.n6071 10.6151
R13139 GND.n6071 GND.n5685 10.6151
R13140 GND.n5754 GND.n5685 10.6151
R13141 GND.n5754 GND.n5702 10.6151
R13142 GND.n6059 GND.n5702 10.6151
R13143 GND.n6059 GND.n6058 10.6151
R13144 GND.n6058 GND.n6057 10.6151
R13145 GND.n6057 GND.n5703 10.6151
R13146 GND.n5774 GND.n5703 10.6151
R13147 GND.n5775 GND.n5774 10.6151
R13148 GND.n5776 GND.n5775 10.6151
R13149 GND.n6040 GND.n5776 10.6151
R13150 GND.n6040 GND.n6039 10.6151
R13151 GND.n6039 GND.n6038 10.6151
R13152 GND.n6038 GND.n5777 10.6151
R13153 GND.n5858 GND.n5777 10.6151
R13154 GND.n5858 GND.n5797 10.6151
R13155 GND.n6026 GND.n5797 10.6151
R13156 GND.n6026 GND.n6025 10.6151
R13157 GND.n6025 GND.n6024 10.6151
R13158 GND.n6024 GND.n5798 10.6151
R13159 GND.n5872 GND.n5798 10.6151
R13160 GND.n5872 GND.n5814 10.6151
R13161 GND.n6012 GND.n5814 10.6151
R13162 GND.n6012 GND.n6011 10.6151
R13163 GND.n6011 GND.n6010 10.6151
R13164 GND.n6010 GND.n5815 10.6151
R13165 GND.n5885 GND.n5815 10.6151
R13166 GND.n5885 GND.n5832 10.6151
R13167 GND.n5998 GND.n5832 10.6151
R13168 GND.n5998 GND.n5997 10.6151
R13169 GND.n5997 GND.n5996 10.6151
R13170 GND.n5996 GND.n5833 10.6151
R13171 GND.n5905 GND.n5833 10.6151
R13172 GND.n5906 GND.n5905 10.6151
R13173 GND.n5907 GND.n5906 10.6151
R13174 GND.n5979 GND.n5907 10.6151
R13175 GND.n5979 GND.n5978 10.6151
R13176 GND.n5978 GND.n5977 10.6151
R13177 GND.n5977 GND.n5908 10.6151
R13178 GND.n5938 GND.n5908 10.6151
R13179 GND.n5938 GND.n5928 10.6151
R13180 GND.n5965 GND.n5928 10.6151
R13181 GND.n5965 GND.n5964 10.6151
R13182 GND.n5964 GND.n5963 10.6151
R13183 GND.n5963 GND.n5929 10.6151
R13184 GND.n5929 GND.n1590 10.6151
R13185 GND.n6426 GND.n1590 10.6151
R13186 GND.n6427 GND.n6426 10.6151
R13187 GND.n6428 GND.n6427 10.6151
R13188 GND.n6428 GND.n1576 10.6151
R13189 GND.n6444 GND.n1576 10.6151
R13190 GND.n6445 GND.n6444 10.6151
R13191 GND.n6446 GND.n6445 10.6151
R13192 GND.n6446 GND.n1561 10.6151
R13193 GND.n6460 GND.n1561 10.6151
R13194 GND.n6461 GND.n6460 10.6151
R13195 GND.n6464 GND.n6461 10.6151
R13196 GND.n6464 GND.n6463 10.6151
R13197 GND.n6463 GND.n6462 10.6151
R13198 GND.n6462 GND.n1532 10.6151
R13199 GND.n6498 GND.n1532 10.6151
R13200 GND.n6499 GND.n6498 10.6151
R13201 GND.n6500 GND.n6499 10.6151
R13202 GND.n6500 GND.n1522 10.6151
R13203 GND.n6525 GND.n1522 10.6151
R13204 GND.n6525 GND.n6524 10.6151
R13205 GND.n6524 GND.n6523 10.6151
R13206 GND.n6523 GND.n1523 10.6151
R13207 GND.n1524 GND.n1523 10.6151
R13208 GND.n1524 GND.n1488 10.6151
R13209 GND.n6584 GND.n1488 10.6151
R13210 GND.n6585 GND.n6584 10.6151
R13211 GND.n6595 GND.n6585 10.6151
R13212 GND.n6595 GND.n6594 10.6151
R13213 GND.n6594 GND.n6593 10.6151
R13214 GND.n6593 GND.n6586 10.6151
R13215 GND.n6587 GND.n6586 10.6151
R13216 GND.n6587 GND.n1447 10.6151
R13217 GND.n6632 GND.n1447 10.6151
R13218 GND.n6632 GND.n6631 10.6151
R13219 GND.n6631 GND.n6630 10.6151
R13220 GND.n6630 GND.n1448 10.6151
R13221 GND.n1456 GND.n1448 10.6151
R13222 GND.n1456 GND.n1455 10.6151
R13223 GND.n1455 GND.n1454 10.6151
R13224 GND.n1454 GND.n1449 10.6151
R13225 GND.n1449 GND.n1399 10.6151
R13226 GND.n6709 GND.n1399 10.6151
R13227 GND.n6710 GND.n6709 10.6151
R13228 GND.n6711 GND.n6710 10.6151
R13229 GND.n6711 GND.n1385 10.6151
R13230 GND.n6757 GND.n1385 10.6151
R13231 GND.n6758 GND.n6757 10.6151
R13232 GND.n6759 GND.n6758 10.6151
R13233 GND.n6759 GND.n1368 10.6151
R13234 GND.n6775 GND.n1368 10.6151
R13235 GND.n6776 GND.n6775 10.6151
R13236 GND.n6778 GND.n6776 10.6151
R13237 GND.n6778 GND.n6777 10.6151
R13238 GND.n6777 GND.n1354 10.6151
R13239 GND.n6826 GND.n1354 10.6151
R13240 GND.n6826 GND.n6825 10.6151
R13241 GND.n6825 GND.n6824 10.6151
R13242 GND.n6824 GND.n1335 10.6151
R13243 GND.n6852 GND.n1335 10.6151
R13244 GND.n6853 GND.n6852 10.6151
R13245 GND.n6854 GND.n6853 10.6151
R13246 GND.n6854 GND.n1312 10.6151
R13247 GND.n6882 GND.n1312 10.6151
R13248 GND.n6883 GND.n6882 10.6151
R13249 GND.n6884 GND.n6883 10.6151
R13250 GND.n6884 GND.n1299 10.6151
R13251 GND.n6912 GND.n1299 10.6151
R13252 GND.n6913 GND.n6912 10.6151
R13253 GND.n6915 GND.n6913 10.6151
R13254 GND.n6915 GND.n6914 10.6151
R13255 GND.n6914 GND.n1170 10.6151
R13256 GND.n6987 GND.n1170 10.6151
R13257 GND.n6988 GND.n6987 10.6151
R13258 GND.n6989 GND.n6988 10.6151
R13259 GND.n6989 GND.n1159 10.6151
R13260 GND.n7005 GND.n1159 10.6151
R13261 GND.n7006 GND.n7005 10.6151
R13262 GND.n7007 GND.n7006 10.6151
R13263 GND.n7007 GND.n1145 10.6151
R13264 GND.n7029 GND.n1145 10.6151
R13265 GND.n7030 GND.n7029 10.6151
R13266 GND.n7031 GND.n7030 10.6151
R13267 GND.n7031 GND.n1135 10.6151
R13268 GND.n7042 GND.n1135 10.6151
R13269 GND.n7043 GND.n7042 10.6151
R13270 GND.n7046 GND.n7043 10.6151
R13271 GND.n7046 GND.n7045 10.6151
R13272 GND.n7045 GND.n7044 10.6151
R13273 GND.n7044 GND.n1114 10.6151
R13274 GND.n7078 GND.n1114 10.6151
R13275 GND.n7079 GND.n7078 10.6151
R13276 GND.n7080 GND.n7079 10.6151
R13277 GND.n7080 GND.n1104 10.6151
R13278 GND.n7091 GND.n1104 10.6151
R13279 GND.n7092 GND.n7091 10.6151
R13280 GND.n7093 GND.n7092 10.6151
R13281 GND.n7093 GND.n1094 10.6151
R13282 GND.n7109 GND.n1094 10.6151
R13283 GND.n7110 GND.n7109 10.6151
R13284 GND.n7111 GND.n7110 10.6151
R13285 GND.n7111 GND.n1080 10.6151
R13286 GND.n7127 GND.n1080 10.6151
R13287 GND.n7128 GND.n7127 10.6151
R13288 GND.n7129 GND.n7128 10.6151
R13289 GND.n7129 GND.n1069 10.6151
R13290 GND.n7144 GND.n1069 10.6151
R13291 GND.n7145 GND.n7144 10.6151
R13292 GND.n7146 GND.n7145 10.6151
R13293 GND.n7146 GND.n1054 10.6151
R13294 GND.n7165 GND.n1054 10.6151
R13295 GND.n7166 GND.n7165 10.6151
R13296 GND.n7167 GND.n7166 10.6151
R13297 GND.n7167 GND.n1045 10.6151
R13298 GND.n7183 GND.n1045 10.6151
R13299 GND.n7184 GND.n7183 10.6151
R13300 GND.n7185 GND.n7184 10.6151
R13301 GND.n7185 GND.n1031 10.6151
R13302 GND.n7210 GND.n1031 10.6151
R13303 GND.n7211 GND.n7210 10.6151
R13304 GND.n7212 GND.n7211 10.6151
R13305 GND.n7212 GND.n1021 10.6151
R13306 GND.n7223 GND.n1021 10.6151
R13307 GND.n7224 GND.n7223 10.6151
R13308 GND.n7225 GND.n7224 10.6151
R13309 GND.n7225 GND.n1011 10.6151
R13310 GND.n7241 GND.n1011 10.6151
R13311 GND.n7242 GND.n7241 10.6151
R13312 GND.n7243 GND.n7242 10.6151
R13313 GND.n7243 GND.n997 10.6151
R13314 GND.n7259 GND.n997 10.6151
R13315 GND.n7260 GND.n7259 10.6151
R13316 GND.n7261 GND.n7260 10.6151
R13317 GND.n7261 GND.n986 10.6151
R13318 GND.n7276 GND.n986 10.6151
R13319 GND.n7277 GND.n7276 10.6151
R13320 GND.n7278 GND.n7277 10.6151
R13321 GND.n7278 GND.n971 10.6151
R13322 GND.n7296 GND.n971 10.6151
R13323 GND.n7297 GND.n7296 10.6151
R13324 GND.n7298 GND.n7297 10.6151
R13325 GND.n7298 GND.n961 10.6151
R13326 GND.n7314 GND.n961 10.6151
R13327 GND.n7315 GND.n7314 10.6151
R13328 GND.n7316 GND.n7315 10.6151
R13329 GND.n7316 GND.n947 10.6151
R13330 GND.n7332 GND.n947 10.6151
R13331 GND.n7333 GND.n7332 10.6151
R13332 GND.n7334 GND.n7333 10.6151
R13333 GND.n7334 GND.n936 10.6151
R13334 GND.n7349 GND.n936 10.6151
R13335 GND.n7350 GND.n7349 10.6151
R13336 GND.n7351 GND.n7350 10.6151
R13337 GND.n7351 GND.n922 10.6151
R13338 GND.n7365 GND.n922 10.6151
R13339 GND.n7366 GND.n7365 10.6151
R13340 GND.n7368 GND.n7366 10.6151
R13341 GND.n7368 GND.n7367 10.6151
R13342 GND.n7367 GND.n905 10.6151
R13343 GND.n7392 GND.n905 10.6151
R13344 GND.n7393 GND.n7392 10.6151
R13345 GND.n7394 GND.n7393 10.6151
R13346 GND.n7394 GND.n896 10.6151
R13347 GND.n7409 GND.n896 10.6151
R13348 GND.n7410 GND.n7409 10.6151
R13349 GND.n7411 GND.n7410 10.6151
R13350 GND.n7411 GND.n882 10.6151
R13351 GND.n7425 GND.n882 10.6151
R13352 GND.n7426 GND.n7425 10.6151
R13353 GND.n7428 GND.n7426 10.6151
R13354 GND.n7428 GND.n7427 10.6151
R13355 GND.n7427 GND.n864 10.6151
R13356 GND.n7509 GND.n864 10.6151
R13357 GND.n7510 GND.n7509 10.6151
R13358 GND.n5519 GND.t147 10.6029
R13359 GND.n6109 GND.t10 10.6029
R13360 GND.t81 GND.n5689 10.6029
R13361 GND.n6430 GND.n1588 10.6029
R13362 GND.n6519 GND.n1525 10.6029
R13363 GND.n6574 GND.n6573 10.6029
R13364 GND.n6762 GND.n6761 10.6029
R13365 GND.n6790 GND.n1360 10.6029
R13366 GND.n6984 GND.n1175 10.6029
R13367 GND.t3 GND.n1028 10.6029
R13368 GND.n7294 GND.t85 10.6029
R13369 GND.n7388 GND.t106 10.6029
R13370 GND.n1777 GND.n1771 10.4732
R13371 GND.n7602 GND.n7599 10.4732
R13372 GND.n8338 GND.n8335 10.4732
R13373 GND.n2873 GND.n2870 10.4732
R13374 GND.n1795 GND.n1794 10.2793
R13375 GND.n7622 GND.n7621 10.2793
R13376 GND.n8359 GND.n8358 10.2793
R13377 GND.n2893 GND.n2892 10.2793
R13378 GND.n1812 GND.n1738 10.0853
R13379 GND.n7645 GND.n7642 10.0853
R13380 GND.n8384 GND.n8381 10.0853
R13381 GND.n2916 GND.n2913 10.0853
R13382 GND.n5424 GND.n5418 9.89608
R13383 GND.n6158 GND.n6157 9.89608
R13384 GND.n5574 GND.n5568 9.89608
R13385 GND.n6097 GND.n6096 9.89608
R13386 GND.n5705 GND.n5699 9.89608
R13387 GND.n6036 GND.n6035 9.89608
R13388 GND.n5835 GND.n5829 9.89608
R13389 GND.n5975 GND.n5974 9.89608
R13390 GND.n6458 GND.n1563 9.89608
R13391 GND.n6503 GND.n6502 9.89608
R13392 GND.n1462 GND.n1444 9.89608
R13393 GND.n6707 GND.n6706 9.89608
R13394 GND.n6850 GND.n1337 9.89608
R13395 GND.n6910 GND.n6909 9.89608
R13396 GND.n7040 GND.n1137 9.89608
R13397 GND.n7082 GND.n1112 9.89608
R13398 GND.n1067 GND.n1056 9.89608
R13399 GND.n1043 GND.n1033 9.89608
R13400 GND.n7274 GND.n988 9.89608
R13401 GND.n7312 GND.n7311 9.89608
R13402 GND.n7390 GND.n907 9.89608
R13403 GND.n7423 GND.n7422 9.89608
R13404 GND.n6251 GND.n6250 9.89141
R13405 GND.n7662 GND.n7661 9.89141
R13406 GND.n8405 GND.n8404 9.89141
R13407 GND.n2936 GND.n2935 9.89141
R13408 GND.n6268 GND.n1705 9.69747
R13409 GND.n7685 GND.n7682 9.69747
R13410 GND.n8430 GND.n8427 9.69747
R13411 GND.n2959 GND.n2956 9.69747
R13412 GND.n7521 GND.n7520 9.36635
R13413 GND.n7444 GND.n7436 9.36635
R13414 GND.n5451 GND.n5450 9.36635
R13415 GND.n6202 GND.n6201 9.36635
R13416 GND.n2782 GND.n2781 9.3005
R13417 GND.n2779 GND.n2763 9.3005
R13418 GND.n2778 GND.n2764 9.3005
R13419 GND.n2776 GND.n2765 9.3005
R13420 GND.n2775 GND.n2766 9.3005
R13421 GND.n2773 GND.n2767 9.3005
R13422 GND.n2772 GND.n2768 9.3005
R13423 GND.n2770 GND.n2769 9.3005
R13424 GND.n2049 GND.n2048 9.3005
R13425 GND.n5120 GND.n5119 9.3005
R13426 GND.n5121 GND.n2047 9.3005
R13427 GND.n5185 GND.n5122 9.3005
R13428 GND.n5184 GND.n5123 9.3005
R13429 GND.n5183 GND.n5124 9.3005
R13430 GND.n5181 GND.n5125 9.3005
R13431 GND.n5180 GND.n5126 9.3005
R13432 GND.n5178 GND.n5127 9.3005
R13433 GND.n5177 GND.n5128 9.3005
R13434 GND.n5175 GND.n5129 9.3005
R13435 GND.n5174 GND.n5130 9.3005
R13436 GND.n5172 GND.n5131 9.3005
R13437 GND.n5171 GND.n5132 9.3005
R13438 GND.n5169 GND.n5133 9.3005
R13439 GND.n5168 GND.n5134 9.3005
R13440 GND.n5166 GND.n5135 9.3005
R13441 GND.n5165 GND.n5136 9.3005
R13442 GND.n5163 GND.n5137 9.3005
R13443 GND.n5162 GND.n5138 9.3005
R13444 GND.n5160 GND.n5139 9.3005
R13445 GND.n5159 GND.n5140 9.3005
R13446 GND.n5157 GND.n5141 9.3005
R13447 GND.n5156 GND.n5142 9.3005
R13448 GND.n5154 GND.n5143 9.3005
R13449 GND.n5153 GND.n5144 9.3005
R13450 GND.n5151 GND.n5145 9.3005
R13451 GND.n5150 GND.n5146 9.3005
R13452 GND.n5148 GND.n5147 9.3005
R13453 GND.n1902 GND.n1901 9.3005
R13454 GND.n5336 GND.n5335 9.3005
R13455 GND.n5337 GND.n1900 9.3005
R13456 GND.n5355 GND.n5338 9.3005
R13457 GND.n5354 GND.n5339 9.3005
R13458 GND.n5353 GND.n5340 9.3005
R13459 GND.n5351 GND.n5341 9.3005
R13460 GND.n5350 GND.n5342 9.3005
R13461 GND.n5348 GND.n5343 9.3005
R13462 GND.n5347 GND.n5344 9.3005
R13463 GND.n5345 GND.n1617 9.3005
R13464 GND.n4726 GND.n4725 9.3005
R13465 GND.n4724 GND.n3023 9.3005
R13466 GND.n3029 GND.n3024 9.3005
R13467 GND.n4718 GND.n3030 9.3005
R13468 GND.n4717 GND.n3031 9.3005
R13469 GND.n4716 GND.n3032 9.3005
R13470 GND.n3037 GND.n3033 9.3005
R13471 GND.n4710 GND.n3038 9.3005
R13472 GND.n4709 GND.n3039 9.3005
R13473 GND.n4708 GND.n3040 9.3005
R13474 GND.n3045 GND.n3041 9.3005
R13475 GND.n4702 GND.n3046 9.3005
R13476 GND.n4701 GND.n3047 9.3005
R13477 GND.n4700 GND.n3048 9.3005
R13478 GND.n3053 GND.n3049 9.3005
R13479 GND.n4694 GND.n3054 9.3005
R13480 GND.n4693 GND.n3055 9.3005
R13481 GND.n4692 GND.n3056 9.3005
R13482 GND.n3061 GND.n3057 9.3005
R13483 GND.n4686 GND.n3062 9.3005
R13484 GND.n4685 GND.n3063 9.3005
R13485 GND.n4684 GND.n3064 9.3005
R13486 GND.n3069 GND.n3065 9.3005
R13487 GND.n4678 GND.n3070 9.3005
R13488 GND.n4677 GND.n3071 9.3005
R13489 GND.n4676 GND.n3072 9.3005
R13490 GND.n3077 GND.n3073 9.3005
R13491 GND.n4670 GND.n3078 9.3005
R13492 GND.n4669 GND.n3079 9.3005
R13493 GND.n4668 GND.n3080 9.3005
R13494 GND.n3085 GND.n3081 9.3005
R13495 GND.n4662 GND.n3086 9.3005
R13496 GND.n4661 GND.n3087 9.3005
R13497 GND.n4660 GND.n3088 9.3005
R13498 GND.n3093 GND.n3089 9.3005
R13499 GND.n4654 GND.n3094 9.3005
R13500 GND.n4653 GND.n3095 9.3005
R13501 GND.n4652 GND.n3096 9.3005
R13502 GND.n3101 GND.n3097 9.3005
R13503 GND.n4646 GND.n3102 9.3005
R13504 GND.n4645 GND.n3103 9.3005
R13505 GND.n4644 GND.n3104 9.3005
R13506 GND.n3109 GND.n3105 9.3005
R13507 GND.n4638 GND.n3110 9.3005
R13508 GND.n4637 GND.n3111 9.3005
R13509 GND.n4636 GND.n3112 9.3005
R13510 GND.n3117 GND.n3113 9.3005
R13511 GND.n4630 GND.n3118 9.3005
R13512 GND.n4629 GND.n3119 9.3005
R13513 GND.n4628 GND.n3120 9.3005
R13514 GND.n3125 GND.n3121 9.3005
R13515 GND.n4622 GND.n3126 9.3005
R13516 GND.n4621 GND.n3127 9.3005
R13517 GND.n4620 GND.n3128 9.3005
R13518 GND.n3133 GND.n3129 9.3005
R13519 GND.n4614 GND.n3134 9.3005
R13520 GND.n4613 GND.n3135 9.3005
R13521 GND.n4612 GND.n3136 9.3005
R13522 GND.n3141 GND.n3137 9.3005
R13523 GND.n4606 GND.n3142 9.3005
R13524 GND.n4605 GND.n3143 9.3005
R13525 GND.n4604 GND.n3144 9.3005
R13526 GND.n3149 GND.n3145 9.3005
R13527 GND.n4598 GND.n3150 9.3005
R13528 GND.n4597 GND.n3151 9.3005
R13529 GND.n4596 GND.n3152 9.3005
R13530 GND.n3157 GND.n3153 9.3005
R13531 GND.n4590 GND.n3158 9.3005
R13532 GND.n4589 GND.n3159 9.3005
R13533 GND.n4588 GND.n3160 9.3005
R13534 GND.n3165 GND.n3161 9.3005
R13535 GND.n4582 GND.n3166 9.3005
R13536 GND.n4581 GND.n3167 9.3005
R13537 GND.n4580 GND.n3168 9.3005
R13538 GND.n3173 GND.n3169 9.3005
R13539 GND.n4574 GND.n3174 9.3005
R13540 GND.n4573 GND.n3175 9.3005
R13541 GND.n4572 GND.n3176 9.3005
R13542 GND.n3181 GND.n3177 9.3005
R13543 GND.n4566 GND.n3182 9.3005
R13544 GND.n4565 GND.n3183 9.3005
R13545 GND.n4564 GND.n3184 9.3005
R13546 GND.n3189 GND.n3185 9.3005
R13547 GND.n4558 GND.n3190 9.3005
R13548 GND.n4557 GND.n3191 9.3005
R13549 GND.n4556 GND.n3192 9.3005
R13550 GND.n3197 GND.n3193 9.3005
R13551 GND.n4550 GND.n3198 9.3005
R13552 GND.n4549 GND.n3199 9.3005
R13553 GND.n4548 GND.n3200 9.3005
R13554 GND.n3205 GND.n3201 9.3005
R13555 GND.n4542 GND.n3206 9.3005
R13556 GND.n4541 GND.n3207 9.3005
R13557 GND.n4540 GND.n3208 9.3005
R13558 GND.n3213 GND.n3209 9.3005
R13559 GND.n4534 GND.n3214 9.3005
R13560 GND.n4533 GND.n3215 9.3005
R13561 GND.n4532 GND.n3216 9.3005
R13562 GND.n3221 GND.n3217 9.3005
R13563 GND.n4526 GND.n3222 9.3005
R13564 GND.n4525 GND.n3223 9.3005
R13565 GND.n4524 GND.n3224 9.3005
R13566 GND.n3229 GND.n3225 9.3005
R13567 GND.n4518 GND.n3230 9.3005
R13568 GND.n4517 GND.n3231 9.3005
R13569 GND.n4516 GND.n3232 9.3005
R13570 GND.n3237 GND.n3233 9.3005
R13571 GND.n4510 GND.n3238 9.3005
R13572 GND.n4509 GND.n3239 9.3005
R13573 GND.n4508 GND.n3240 9.3005
R13574 GND.n3245 GND.n3241 9.3005
R13575 GND.n4502 GND.n3246 9.3005
R13576 GND.n4501 GND.n3247 9.3005
R13577 GND.n4500 GND.n3248 9.3005
R13578 GND.n3253 GND.n3249 9.3005
R13579 GND.n4494 GND.n3254 9.3005
R13580 GND.n4493 GND.n3255 9.3005
R13581 GND.n4492 GND.n3256 9.3005
R13582 GND.n3261 GND.n3257 9.3005
R13583 GND.n4486 GND.n3262 9.3005
R13584 GND.n4485 GND.n3263 9.3005
R13585 GND.n4484 GND.n3264 9.3005
R13586 GND.n3269 GND.n3265 9.3005
R13587 GND.n4478 GND.n3270 9.3005
R13588 GND.n4477 GND.n3271 9.3005
R13589 GND.n4476 GND.n3272 9.3005
R13590 GND.n3277 GND.n3273 9.3005
R13591 GND.n4470 GND.n3278 9.3005
R13592 GND.n4469 GND.n3279 9.3005
R13593 GND.n4468 GND.n3280 9.3005
R13594 GND.n3285 GND.n3281 9.3005
R13595 GND.n4462 GND.n3286 9.3005
R13596 GND.n4461 GND.n3287 9.3005
R13597 GND.n4460 GND.n3288 9.3005
R13598 GND.n3293 GND.n3289 9.3005
R13599 GND.n4454 GND.n3294 9.3005
R13600 GND.n4453 GND.n3295 9.3005
R13601 GND.n4452 GND.n3296 9.3005
R13602 GND.n3301 GND.n3297 9.3005
R13603 GND.n4446 GND.n3302 9.3005
R13604 GND.n4445 GND.n3303 9.3005
R13605 GND.n4444 GND.n3304 9.3005
R13606 GND.n3309 GND.n3305 9.3005
R13607 GND.n4438 GND.n3310 9.3005
R13608 GND.n4437 GND.n3311 9.3005
R13609 GND.n4436 GND.n3312 9.3005
R13610 GND.n3317 GND.n3313 9.3005
R13611 GND.n4430 GND.n3318 9.3005
R13612 GND.n4429 GND.n3319 9.3005
R13613 GND.n4428 GND.n3320 9.3005
R13614 GND.n3325 GND.n3321 9.3005
R13615 GND.n4422 GND.n3326 9.3005
R13616 GND.n4421 GND.n3327 9.3005
R13617 GND.n4420 GND.n3328 9.3005
R13618 GND.n3333 GND.n3329 9.3005
R13619 GND.n4414 GND.n3334 9.3005
R13620 GND.n4413 GND.n3335 9.3005
R13621 GND.n4412 GND.n3336 9.3005
R13622 GND.n3341 GND.n3337 9.3005
R13623 GND.n4406 GND.n3342 9.3005
R13624 GND.n4405 GND.n3343 9.3005
R13625 GND.n4404 GND.n3344 9.3005
R13626 GND.n3349 GND.n3345 9.3005
R13627 GND.n4398 GND.n3350 9.3005
R13628 GND.n4397 GND.n3351 9.3005
R13629 GND.n4396 GND.n3352 9.3005
R13630 GND.n3357 GND.n3353 9.3005
R13631 GND.n4390 GND.n3358 9.3005
R13632 GND.n4389 GND.n3359 9.3005
R13633 GND.n4388 GND.n3360 9.3005
R13634 GND.n3365 GND.n3361 9.3005
R13635 GND.n4382 GND.n3366 9.3005
R13636 GND.n4381 GND.n3367 9.3005
R13637 GND.n4380 GND.n3368 9.3005
R13638 GND.n3373 GND.n3369 9.3005
R13639 GND.n4374 GND.n3374 9.3005
R13640 GND.n4373 GND.n3375 9.3005
R13641 GND.n4372 GND.n3376 9.3005
R13642 GND.n3381 GND.n3377 9.3005
R13643 GND.n4366 GND.n3382 9.3005
R13644 GND.n4365 GND.n3383 9.3005
R13645 GND.n4364 GND.n3384 9.3005
R13646 GND.n3389 GND.n3385 9.3005
R13647 GND.n4358 GND.n3390 9.3005
R13648 GND.n4357 GND.n3391 9.3005
R13649 GND.n4356 GND.n3392 9.3005
R13650 GND.n3397 GND.n3393 9.3005
R13651 GND.n4350 GND.n3398 9.3005
R13652 GND.n4349 GND.n3399 9.3005
R13653 GND.n4348 GND.n3400 9.3005
R13654 GND.n3405 GND.n3401 9.3005
R13655 GND.n4342 GND.n3406 9.3005
R13656 GND.n4341 GND.n3407 9.3005
R13657 GND.n4340 GND.n3408 9.3005
R13658 GND.n3413 GND.n3409 9.3005
R13659 GND.n4334 GND.n3414 9.3005
R13660 GND.n4333 GND.n3415 9.3005
R13661 GND.n4332 GND.n3416 9.3005
R13662 GND.n3421 GND.n3417 9.3005
R13663 GND.n4326 GND.n3422 9.3005
R13664 GND.n4325 GND.n3423 9.3005
R13665 GND.n4324 GND.n3424 9.3005
R13666 GND.n3429 GND.n3425 9.3005
R13667 GND.n4318 GND.n3430 9.3005
R13668 GND.n4317 GND.n3431 9.3005
R13669 GND.n4316 GND.n3432 9.3005
R13670 GND.n3437 GND.n3433 9.3005
R13671 GND.n4310 GND.n3438 9.3005
R13672 GND.n4309 GND.n3439 9.3005
R13673 GND.n4308 GND.n3440 9.3005
R13674 GND.n3445 GND.n3441 9.3005
R13675 GND.n4302 GND.n3446 9.3005
R13676 GND.n4301 GND.n3447 9.3005
R13677 GND.n4300 GND.n3448 9.3005
R13678 GND.n3453 GND.n3449 9.3005
R13679 GND.n4294 GND.n3454 9.3005
R13680 GND.n4293 GND.n3455 9.3005
R13681 GND.n4292 GND.n3456 9.3005
R13682 GND.n3461 GND.n3457 9.3005
R13683 GND.n4286 GND.n3462 9.3005
R13684 GND.n4285 GND.n3463 9.3005
R13685 GND.n4284 GND.n3464 9.3005
R13686 GND.n3469 GND.n3465 9.3005
R13687 GND.n4278 GND.n3470 9.3005
R13688 GND.n4277 GND.n3471 9.3005
R13689 GND.n4276 GND.n3472 9.3005
R13690 GND.n3477 GND.n3473 9.3005
R13691 GND.n4270 GND.n3478 9.3005
R13692 GND.n4269 GND.n3479 9.3005
R13693 GND.n4268 GND.n3480 9.3005
R13694 GND.n3485 GND.n3481 9.3005
R13695 GND.n4262 GND.n3486 9.3005
R13696 GND.n4261 GND.n3487 9.3005
R13697 GND.n4260 GND.n3488 9.3005
R13698 GND.n3493 GND.n3489 9.3005
R13699 GND.n4254 GND.n3494 9.3005
R13700 GND.n4253 GND.n3495 9.3005
R13701 GND.n4252 GND.n3496 9.3005
R13702 GND.n3501 GND.n3497 9.3005
R13703 GND.n4246 GND.n3502 9.3005
R13704 GND.n4245 GND.n3503 9.3005
R13705 GND.n4244 GND.n3504 9.3005
R13706 GND.n3509 GND.n3505 9.3005
R13707 GND.n4238 GND.n3510 9.3005
R13708 GND.n4237 GND.n3511 9.3005
R13709 GND.n4236 GND.n3512 9.3005
R13710 GND.n3517 GND.n3513 9.3005
R13711 GND.n4230 GND.n3518 9.3005
R13712 GND.n4229 GND.n3519 9.3005
R13713 GND.n4228 GND.n3520 9.3005
R13714 GND.n3525 GND.n3521 9.3005
R13715 GND.n4222 GND.n3526 9.3005
R13716 GND.n4221 GND.n3527 9.3005
R13717 GND.n4220 GND.n3528 9.3005
R13718 GND.n3533 GND.n3529 9.3005
R13719 GND.n4214 GND.n3534 9.3005
R13720 GND.n4213 GND.n3535 9.3005
R13721 GND.n4212 GND.n3536 9.3005
R13722 GND.n3541 GND.n3537 9.3005
R13723 GND.n4206 GND.n3542 9.3005
R13724 GND.n4205 GND.n3543 9.3005
R13725 GND.n4204 GND.n3544 9.3005
R13726 GND.n3549 GND.n3545 9.3005
R13727 GND.n4198 GND.n3550 9.3005
R13728 GND.n4197 GND.n3551 9.3005
R13729 GND.n4196 GND.n3552 9.3005
R13730 GND.n3557 GND.n3553 9.3005
R13731 GND.n4190 GND.n3558 9.3005
R13732 GND.n4189 GND.n3559 9.3005
R13733 GND.n4188 GND.n3560 9.3005
R13734 GND.n3565 GND.n3561 9.3005
R13735 GND.n4182 GND.n3566 9.3005
R13736 GND.n4181 GND.n3567 9.3005
R13737 GND.n4180 GND.n3568 9.3005
R13738 GND.n3573 GND.n3569 9.3005
R13739 GND.n4174 GND.n3574 9.3005
R13740 GND.n4173 GND.n3575 9.3005
R13741 GND.n4172 GND.n3576 9.3005
R13742 GND.n3581 GND.n3577 9.3005
R13743 GND.n4166 GND.n3582 9.3005
R13744 GND.n4165 GND.n3583 9.3005
R13745 GND.n4164 GND.n3584 9.3005
R13746 GND.n3589 GND.n3585 9.3005
R13747 GND.n4158 GND.n3590 9.3005
R13748 GND.n4157 GND.n3591 9.3005
R13749 GND.n4156 GND.n3592 9.3005
R13750 GND.n3597 GND.n3593 9.3005
R13751 GND.n4150 GND.n3598 9.3005
R13752 GND.n4149 GND.n3599 9.3005
R13753 GND.n4148 GND.n3600 9.3005
R13754 GND.n3605 GND.n3601 9.3005
R13755 GND.n4142 GND.n3606 9.3005
R13756 GND.n4141 GND.n3607 9.3005
R13757 GND.n4140 GND.n3608 9.3005
R13758 GND.n3613 GND.n3609 9.3005
R13759 GND.n4134 GND.n3614 9.3005
R13760 GND.n4133 GND.n3615 9.3005
R13761 GND.n4132 GND.n3616 9.3005
R13762 GND.n3621 GND.n3617 9.3005
R13763 GND.n4126 GND.n3622 9.3005
R13764 GND.n4125 GND.n3623 9.3005
R13765 GND.n4124 GND.n3624 9.3005
R13766 GND.n3629 GND.n3625 9.3005
R13767 GND.n4118 GND.n3630 9.3005
R13768 GND.n4117 GND.n3631 9.3005
R13769 GND.n4116 GND.n3632 9.3005
R13770 GND.n3637 GND.n3633 9.3005
R13771 GND.n4110 GND.n3638 9.3005
R13772 GND.n4109 GND.n3639 9.3005
R13773 GND.n4108 GND.n3640 9.3005
R13774 GND.n3645 GND.n3641 9.3005
R13775 GND.n4102 GND.n3646 9.3005
R13776 GND.n4101 GND.n3647 9.3005
R13777 GND.n4100 GND.n3648 9.3005
R13778 GND.n3653 GND.n3649 9.3005
R13779 GND.n4094 GND.n3654 9.3005
R13780 GND.n4093 GND.n3655 9.3005
R13781 GND.n4092 GND.n3656 9.3005
R13782 GND.n3661 GND.n3657 9.3005
R13783 GND.n4086 GND.n3662 9.3005
R13784 GND.n4085 GND.n3663 9.3005
R13785 GND.n4084 GND.n3664 9.3005
R13786 GND.n3669 GND.n3665 9.3005
R13787 GND.n4078 GND.n3670 9.3005
R13788 GND.n4077 GND.n3671 9.3005
R13789 GND.n4076 GND.n3672 9.3005
R13790 GND.n3677 GND.n3673 9.3005
R13791 GND.n4070 GND.n3678 9.3005
R13792 GND.n4069 GND.n3679 9.3005
R13793 GND.n4068 GND.n3680 9.3005
R13794 GND.n3685 GND.n3681 9.3005
R13795 GND.n4062 GND.n3686 9.3005
R13796 GND.n4061 GND.n3687 9.3005
R13797 GND.n4060 GND.n3688 9.3005
R13798 GND.n3693 GND.n3689 9.3005
R13799 GND.n4054 GND.n3694 9.3005
R13800 GND.n4053 GND.n3695 9.3005
R13801 GND.n4052 GND.n3696 9.3005
R13802 GND.n3701 GND.n3697 9.3005
R13803 GND.n4046 GND.n3702 9.3005
R13804 GND.n4045 GND.n3703 9.3005
R13805 GND.n4044 GND.n3704 9.3005
R13806 GND.n3709 GND.n3705 9.3005
R13807 GND.n4038 GND.n3710 9.3005
R13808 GND.n4037 GND.n3711 9.3005
R13809 GND.n4036 GND.n3712 9.3005
R13810 GND.n3717 GND.n3713 9.3005
R13811 GND.n4030 GND.n3718 9.3005
R13812 GND.n4029 GND.n3719 9.3005
R13813 GND.n4028 GND.n3720 9.3005
R13814 GND.n3725 GND.n3721 9.3005
R13815 GND.n4022 GND.n3726 9.3005
R13816 GND.n4021 GND.n3727 9.3005
R13817 GND.n4020 GND.n3728 9.3005
R13818 GND.n3733 GND.n3729 9.3005
R13819 GND.n4014 GND.n3734 9.3005
R13820 GND.n4013 GND.n3735 9.3005
R13821 GND.n4012 GND.n3736 9.3005
R13822 GND.n3741 GND.n3737 9.3005
R13823 GND.n4006 GND.n3742 9.3005
R13824 GND.n4005 GND.n3743 9.3005
R13825 GND.n4004 GND.n3744 9.3005
R13826 GND.n3749 GND.n3745 9.3005
R13827 GND.n3998 GND.n3750 9.3005
R13828 GND.n3997 GND.n3751 9.3005
R13829 GND.n3996 GND.n3752 9.3005
R13830 GND.n3757 GND.n3753 9.3005
R13831 GND.n3990 GND.n3758 9.3005
R13832 GND.n3989 GND.n3759 9.3005
R13833 GND.n3988 GND.n3760 9.3005
R13834 GND.n3765 GND.n3761 9.3005
R13835 GND.n3982 GND.n3766 9.3005
R13836 GND.n3981 GND.n3767 9.3005
R13837 GND.n3980 GND.n3768 9.3005
R13838 GND.n3773 GND.n3769 9.3005
R13839 GND.n3974 GND.n3774 9.3005
R13840 GND.n3973 GND.n3775 9.3005
R13841 GND.n3972 GND.n3776 9.3005
R13842 GND.n3781 GND.n3777 9.3005
R13843 GND.n3966 GND.n3782 9.3005
R13844 GND.n3965 GND.n3964 9.3005
R13845 GND.n3784 GND.n3783 9.3005
R13846 GND.n3956 GND.n3788 9.3005
R13847 GND.n3955 GND.n3789 9.3005
R13848 GND.n3954 GND.n3790 9.3005
R13849 GND.n3795 GND.n3791 9.3005
R13850 GND.n3948 GND.n3796 9.3005
R13851 GND.n3947 GND.n3797 9.3005
R13852 GND.n3946 GND.n3798 9.3005
R13853 GND.n3803 GND.n3799 9.3005
R13854 GND.n3940 GND.n3804 9.3005
R13855 GND.n3939 GND.n3805 9.3005
R13856 GND.n3938 GND.n3806 9.3005
R13857 GND.n3811 GND.n3807 9.3005
R13858 GND.n3932 GND.n3812 9.3005
R13859 GND.n3931 GND.n3813 9.3005
R13860 GND.n3930 GND.n3814 9.3005
R13861 GND.n3819 GND.n3815 9.3005
R13862 GND.n3924 GND.n3820 9.3005
R13863 GND.n3923 GND.n3821 9.3005
R13864 GND.n3922 GND.n3822 9.3005
R13865 GND.n3827 GND.n3823 9.3005
R13866 GND.n3916 GND.n3828 9.3005
R13867 GND.n3915 GND.n3829 9.3005
R13868 GND.n3914 GND.n3830 9.3005
R13869 GND.n3835 GND.n3831 9.3005
R13870 GND.n3908 GND.n3836 9.3005
R13871 GND.n3907 GND.n3837 9.3005
R13872 GND.n3906 GND.n3838 9.3005
R13873 GND.n3843 GND.n3839 9.3005
R13874 GND.n3900 GND.n3844 9.3005
R13875 GND.n3899 GND.n3845 9.3005
R13876 GND.n3898 GND.n3846 9.3005
R13877 GND.n3851 GND.n3847 9.3005
R13878 GND.n3892 GND.n3852 9.3005
R13879 GND.n3891 GND.n3853 9.3005
R13880 GND.n3890 GND.n3854 9.3005
R13881 GND.n3859 GND.n3855 9.3005
R13882 GND.n3884 GND.n3860 9.3005
R13883 GND.n3883 GND.n3861 9.3005
R13884 GND.n3882 GND.n3862 9.3005
R13885 GND.n3867 GND.n3863 9.3005
R13886 GND.n3876 GND.n3868 9.3005
R13887 GND.n3875 GND.n3869 9.3005
R13888 GND.n3874 GND.n3871 9.3005
R13889 GND.n3870 GND.n347 9.3005
R13890 GND.n8452 GND.n346 9.3005
R13891 GND.n8454 GND.n8453 9.3005
R13892 GND.n3963 GND.n3962 9.3005
R13893 GND.n1569 GND.n1568 9.3005
R13894 GND.n6452 GND.n6451 9.3005
R13895 GND.n6453 GND.n1567 9.3005
R13896 GND.n6455 GND.n6454 9.3005
R13897 GND.n1542 GND.n1541 9.3005
R13898 GND.n6485 GND.n6484 9.3005
R13899 GND.n6486 GND.n1540 9.3005
R13900 GND.n6493 GND.n6487 9.3005
R13901 GND.n6492 GND.n6488 9.3005
R13902 GND.n6491 GND.n6489 9.3005
R13903 GND.n1506 GND.n1505 9.3005
R13904 GND.n6548 GND.n6547 9.3005
R13905 GND.n6549 GND.n1504 9.3005
R13906 GND.n6551 GND.n6550 9.3005
R13907 GND.n1480 GND.n1479 9.3005
R13908 GND.n6600 GND.n6599 9.3005
R13909 GND.n6601 GND.n1478 9.3005
R13910 GND.n6603 GND.n6602 9.3005
R13911 GND.n1440 GND.n1439 9.3005
R13912 GND.n6638 GND.n6637 9.3005
R13913 GND.n6639 GND.n1438 9.3005
R13914 GND.n6643 GND.n6640 9.3005
R13915 GND.n6642 GND.n6641 9.3005
R13916 GND.n1409 GND.n1408 9.3005
R13917 GND.n6697 GND.n6696 9.3005
R13918 GND.n6698 GND.n1407 9.3005
R13919 GND.n6702 GND.n6699 9.3005
R13920 GND.n6701 GND.n6700 9.3005
R13921 GND.n1378 GND.n1377 9.3005
R13922 GND.n6765 GND.n6764 9.3005
R13923 GND.n6766 GND.n1376 9.3005
R13924 GND.n6770 GND.n6767 9.3005
R13925 GND.n6769 GND.n6768 9.3005
R13926 GND.n1347 GND.n1346 9.3005
R13927 GND.n6832 GND.n6831 9.3005
R13928 GND.n6833 GND.n1345 9.3005
R13929 GND.n6838 GND.n6834 9.3005
R13930 GND.n6837 GND.n6836 9.3005
R13931 GND.n6835 GND.n1328 9.3005
R13932 GND.n1326 GND.n1325 9.3005
R13933 GND.n6862 GND.n6861 9.3005
R13934 GND.n6863 GND.n1324 9.3005
R13935 GND.n6870 GND.n6864 9.3005
R13936 GND.n6869 GND.n6865 9.3005
R13937 GND.n6868 GND.n6866 9.3005
R13938 GND.n1179 GND.n1178 9.3005
R13939 GND.n6982 GND.n6981 9.3005
R13940 GND.n6313 GND.n6312 9.3005
R13941 GND.n6340 GND.n1616 9.3005
R13942 GND.n6339 GND.n6303 9.3005
R13943 GND.n6331 GND.n6302 9.3005
R13944 GND.n6333 GND.n6332 9.3005
R13945 GND.n6330 GND.n6305 9.3005
R13946 GND.n6329 GND.n6328 9.3005
R13947 GND.n6307 GND.n6306 9.3005
R13948 GND.n6322 GND.n6321 9.3005
R13949 GND.n6320 GND.n6309 9.3005
R13950 GND.n6319 GND.n6318 9.3005
R13951 GND.n6311 GND.n6310 9.3005
R13952 GND.n6372 GND.n6371 9.3005
R13953 GND.n6370 GND.n1613 9.3005
R13954 GND.n6379 GND.n6378 9.3005
R13955 GND.n6380 GND.n1610 9.3005
R13956 GND.n6405 GND.n6381 9.3005
R13957 GND.n6404 GND.n6382 9.3005
R13958 GND.n6403 GND.n6383 9.3005
R13959 GND.n6402 GND.n6384 9.3005
R13960 GND.n6401 GND.n6385 9.3005
R13961 GND.n6399 GND.n6386 9.3005
R13962 GND.n6398 GND.n6387 9.3005
R13963 GND.n6389 GND.n6388 9.3005
R13964 GND.n6394 GND.n6390 9.3005
R13965 GND.n6393 GND.n6392 9.3005
R13966 GND.n6391 GND.n1500 9.3005
R13967 GND.n6555 GND.n1499 9.3005
R13968 GND.n6557 GND.n6556 9.3005
R13969 GND.n6558 GND.n1498 9.3005
R13970 GND.n6571 GND.n6559 9.3005
R13971 GND.n6570 GND.n6560 9.3005
R13972 GND.n6569 GND.n6561 9.3005
R13973 GND.n6567 GND.n6562 9.3005
R13974 GND.n6566 GND.n6565 9.3005
R13975 GND.n6564 GND.n1433 9.3005
R13976 GND.n6563 GND.n1431 9.3005
R13977 GND.n6649 GND.n1430 9.3005
R13978 GND.n6651 GND.n6650 9.3005
R13979 GND.n6652 GND.n1429 9.3005
R13980 GND.n6654 GND.n6653 9.3005
R13981 GND.n6656 GND.n1427 9.3005
R13982 GND.n6658 GND.n6657 9.3005
R13983 GND.n6659 GND.n1426 9.3005
R13984 GND.n6663 GND.n6660 9.3005
R13985 GND.n6662 GND.n6661 9.3005
R13986 GND.n1358 GND.n1357 9.3005
R13987 GND.n6793 GND.n6792 9.3005
R13988 GND.n6794 GND.n1356 9.3005
R13989 GND.n6819 GND.n6795 9.3005
R13990 GND.n6818 GND.n6796 9.3005
R13991 GND.n6817 GND.n6797 9.3005
R13992 GND.n6816 GND.n6798 9.3005
R13993 GND.n6815 GND.n6799 9.3005
R13994 GND.n6801 GND.n6800 9.3005
R13995 GND.n6811 GND.n6802 9.3005
R13996 GND.n6810 GND.n6803 9.3005
R13997 GND.n6809 GND.n6805 9.3005
R13998 GND.n6804 GND.n1288 9.3005
R13999 GND.n6927 GND.n1287 9.3005
R14000 GND.n6929 GND.n6928 9.3005
R14001 GND.n1612 GND.n1611 9.3005
R14002 GND.n1286 GND.n1284 9.3005
R14003 GND.n6931 GND.n6930 9.3005
R14004 GND.n6978 GND.n1180 9.3005
R14005 GND.n1184 GND.n1181 9.3005
R14006 GND.n1185 GND.n1182 9.3005
R14007 GND.n6971 GND.n1186 9.3005
R14008 GND.n6970 GND.n1187 9.3005
R14009 GND.n6969 GND.n1188 9.3005
R14010 GND.n1192 GND.n1189 9.3005
R14011 GND.n6964 GND.n1193 9.3005
R14012 GND.n6963 GND.n1194 9.3005
R14013 GND.n6962 GND.n1195 9.3005
R14014 GND.n6980 GND.n6979 9.3005
R14015 GND.n1274 GND.n1226 9.3005
R14016 GND.n6956 GND.n1275 9.3005
R14017 GND.n6942 GND.n1275 9.3005
R14018 GND.n1271 GND.n1227 9.3005
R14019 GND.n1270 GND.n1229 9.3005
R14020 GND.n1269 GND.n1230 9.3005
R14021 GND.n1267 GND.n1231 9.3005
R14022 GND.n1266 GND.n1232 9.3005
R14023 GND.n1264 GND.n1233 9.3005
R14024 GND.n1263 GND.n1234 9.3005
R14025 GND.n1261 GND.n1235 9.3005
R14026 GND.n1260 GND.n1236 9.3005
R14027 GND.n1258 GND.n1237 9.3005
R14028 GND.n1257 GND.n1238 9.3005
R14029 GND.n1255 GND.n1239 9.3005
R14030 GND.n1254 GND.n1240 9.3005
R14031 GND.n1252 GND.n1241 9.3005
R14032 GND.n1251 GND.n1242 9.3005
R14033 GND.n1249 GND.n1243 9.3005
R14034 GND.n1248 GND.n1244 9.3005
R14035 GND.n1246 GND.n1245 9.3005
R14036 GND.n565 GND.n564 9.3005
R14037 GND.n7821 GND.n7820 9.3005
R14038 GND.n7822 GND.n563 9.3005
R14039 GND.n7869 GND.n7823 9.3005
R14040 GND.n7868 GND.n7824 9.3005
R14041 GND.n7867 GND.n7825 9.3005
R14042 GND.n7865 GND.n7826 9.3005
R14043 GND.n7864 GND.n7827 9.3005
R14044 GND.n7862 GND.n7828 9.3005
R14045 GND.n7861 GND.n7829 9.3005
R14046 GND.n7859 GND.n7830 9.3005
R14047 GND.n7858 GND.n7831 9.3005
R14048 GND.n7856 GND.n7832 9.3005
R14049 GND.n7855 GND.n7833 9.3005
R14050 GND.n7853 GND.n7834 9.3005
R14051 GND.n7852 GND.n7835 9.3005
R14052 GND.n7850 GND.n7836 9.3005
R14053 GND.n7849 GND.n7837 9.3005
R14054 GND.n7847 GND.n7838 9.3005
R14055 GND.n7846 GND.n7839 9.3005
R14056 GND.n7844 GND.n7840 9.3005
R14057 GND.n7843 GND.n7842 9.3005
R14058 GND.n7841 GND.n108 9.3005
R14059 GND.n8611 GND.n107 9.3005
R14060 GND.n8613 GND.n8612 9.3005
R14061 GND.n8614 GND.n106 9.3005
R14062 GND.n8618 GND.n8615 9.3005
R14063 GND.n8617 GND.n8616 9.3005
R14064 GND.n64 GND.n62 9.3005
R14065 GND.n1273 GND.n1272 9.3005
R14066 GND.n8639 GND.n8638 9.3005
R14067 GND.n65 GND.n63 9.3005
R14068 GND.n8095 GND.n8094 9.3005
R14069 GND.n8098 GND.n8097 9.3005
R14070 GND.n8099 GND.n8093 9.3005
R14071 GND.n8102 GND.n8100 9.3005
R14072 GND.n8103 GND.n8092 9.3005
R14073 GND.n8106 GND.n8105 9.3005
R14074 GND.n8107 GND.n8091 9.3005
R14075 GND.n8110 GND.n8108 9.3005
R14076 GND.n8111 GND.n8090 9.3005
R14077 GND.n8114 GND.n8113 9.3005
R14078 GND.n8115 GND.n8089 9.3005
R14079 GND.n8118 GND.n8116 9.3005
R14080 GND.n8119 GND.n8088 9.3005
R14081 GND.n8122 GND.n8121 9.3005
R14082 GND.n8123 GND.n8087 9.3005
R14083 GND.n8126 GND.n8124 9.3005
R14084 GND.n8127 GND.n8086 9.3005
R14085 GND.n8130 GND.n8129 9.3005
R14086 GND.n8131 GND.n8085 9.3005
R14087 GND.n8134 GND.n8132 9.3005
R14088 GND.n8135 GND.n8084 9.3005
R14089 GND.n8138 GND.n8137 9.3005
R14090 GND.n8139 GND.n8083 9.3005
R14091 GND.n8142 GND.n8140 9.3005
R14092 GND.n8143 GND.n8082 9.3005
R14093 GND.n8146 GND.n8145 9.3005
R14094 GND.n8147 GND.n8081 9.3005
R14095 GND.n8150 GND.n8148 9.3005
R14096 GND.n8151 GND.n8080 9.3005
R14097 GND.n8154 GND.n8153 9.3005
R14098 GND.n8155 GND.n8079 9.3005
R14099 GND.n8158 GND.n8156 9.3005
R14100 GND.n8159 GND.n8078 9.3005
R14101 GND.n8162 GND.n8161 9.3005
R14102 GND.n8163 GND.n8077 9.3005
R14103 GND.n8166 GND.n8164 9.3005
R14104 GND.n8167 GND.n8076 9.3005
R14105 GND.n8170 GND.n8169 9.3005
R14106 GND.n8171 GND.n8075 9.3005
R14107 GND.n8174 GND.n8172 9.3005
R14108 GND.n8175 GND.n8074 9.3005
R14109 GND.n8178 GND.n8177 9.3005
R14110 GND.n8179 GND.n8073 9.3005
R14111 GND.n8221 GND.n8180 9.3005
R14112 GND.n8220 GND.n8181 9.3005
R14113 GND.n8219 GND.n8182 9.3005
R14114 GND.n8218 GND.n8183 9.3005
R14115 GND.n8193 GND.n8192 9.3005
R14116 GND.n8195 GND.n8194 9.3005
R14117 GND.n8198 GND.n8189 9.3005
R14118 GND.n8202 GND.n8201 9.3005
R14119 GND.n8203 GND.n8188 9.3005
R14120 GND.n8205 GND.n8204 9.3005
R14121 GND.n8208 GND.n8187 9.3005
R14122 GND.n8212 GND.n8211 9.3005
R14123 GND.n8213 GND.n8186 9.3005
R14124 GND.n8215 GND.n8214 9.3005
R14125 GND.n8190 GND.n444 9.3005
R14126 GND.n8445 GND.n8444 9.3005
R14127 GND.n8443 GND.n387 9.3005
R14128 GND.n8442 GND.n8441 9.3005
R14129 GND.n8438 GND.n388 9.3005
R14130 GND.n8435 GND.n389 9.3005
R14131 GND.n8434 GND.n390 9.3005
R14132 GND.n8431 GND.n391 9.3005
R14133 GND.n8430 GND.n392 9.3005
R14134 GND.n8427 GND.n8426 9.3005
R14135 GND.n8425 GND.n393 9.3005
R14136 GND.n8424 GND.n8423 9.3005
R14137 GND.n8420 GND.n396 9.3005
R14138 GND.n8417 GND.n397 9.3005
R14139 GND.n8416 GND.n398 9.3005
R14140 GND.n8413 GND.n399 9.3005
R14141 GND.n8412 GND.n400 9.3005
R14142 GND.n8409 GND.n401 9.3005
R14143 GND.n8408 GND.n402 9.3005
R14144 GND.n8405 GND.n403 9.3005
R14145 GND.n8404 GND.n8403 9.3005
R14146 GND.n8402 GND.n404 9.3005
R14147 GND.n8401 GND.n8400 9.3005
R14148 GND.n8397 GND.n409 9.3005
R14149 GND.n8396 GND.n410 9.3005
R14150 GND.n8393 GND.n411 9.3005
R14151 GND.n8392 GND.n412 9.3005
R14152 GND.n8389 GND.n413 9.3005
R14153 GND.n8388 GND.n414 9.3005
R14154 GND.n8385 GND.n415 9.3005
R14155 GND.n8384 GND.n416 9.3005
R14156 GND.n8381 GND.n8380 9.3005
R14157 GND.n8379 GND.n417 9.3005
R14158 GND.n8378 GND.n8377 9.3005
R14159 GND.n8374 GND.n420 9.3005
R14160 GND.n8371 GND.n421 9.3005
R14161 GND.n8370 GND.n422 9.3005
R14162 GND.n8367 GND.n423 9.3005
R14163 GND.n8366 GND.n424 9.3005
R14164 GND.n8363 GND.n425 9.3005
R14165 GND.n8362 GND.n426 9.3005
R14166 GND.n8359 GND.n427 9.3005
R14167 GND.n8358 GND.n8357 9.3005
R14168 GND.n8356 GND.n428 9.3005
R14169 GND.n8355 GND.n8354 9.3005
R14170 GND.n8351 GND.n433 9.3005
R14171 GND.n8350 GND.n434 9.3005
R14172 GND.n8347 GND.n435 9.3005
R14173 GND.n8346 GND.n436 9.3005
R14174 GND.n8343 GND.n437 9.3005
R14175 GND.n8342 GND.n438 9.3005
R14176 GND.n8339 GND.n439 9.3005
R14177 GND.n8338 GND.n440 9.3005
R14178 GND.n8335 GND.n8334 9.3005
R14179 GND.n8333 GND.n441 9.3005
R14180 GND.n8446 GND.n386 9.3005
R14181 GND.n7715 GND.n7714 9.3005
R14182 GND.n7716 GND.n665 9.3005
R14183 GND.n7718 GND.n7717 9.3005
R14184 GND.n7719 GND.n646 9.3005
R14185 GND.n7735 GND.n647 9.3005
R14186 GND.n7736 GND.n645 9.3005
R14187 GND.n7738 GND.n7737 9.3005
R14188 GND.n7739 GND.n626 9.3005
R14189 GND.n7755 GND.n627 9.3005
R14190 GND.n7756 GND.n625 9.3005
R14191 GND.n7758 GND.n7757 9.3005
R14192 GND.n7759 GND.n606 9.3005
R14193 GND.n7775 GND.n607 9.3005
R14194 GND.n7776 GND.n605 9.3005
R14195 GND.n7778 GND.n7777 9.3005
R14196 GND.n7779 GND.n586 9.3005
R14197 GND.n7795 GND.n587 9.3005
R14198 GND.n7796 GND.n584 9.3005
R14199 GND.n7798 GND.n585 9.3005
R14200 GND.n7800 GND.n7799 9.3005
R14201 GND.n7801 GND.n557 9.3005
R14202 GND.n7873 GND.n558 9.3005
R14203 GND.n7874 GND.n556 9.3005
R14204 GND.n7876 GND.n7875 9.3005
R14205 GND.n7877 GND.n538 9.3005
R14206 GND.n7893 GND.n539 9.3005
R14207 GND.n7894 GND.n537 9.3005
R14208 GND.n7896 GND.n7895 9.3005
R14209 GND.n7897 GND.n518 9.3005
R14210 GND.n7913 GND.n519 9.3005
R14211 GND.n7914 GND.n517 9.3005
R14212 GND.n7916 GND.n7915 9.3005
R14213 GND.n7917 GND.n498 9.3005
R14214 GND.n7933 GND.n499 9.3005
R14215 GND.n7934 GND.n496 9.3005
R14216 GND.n7936 GND.n497 9.3005
R14217 GND.n7944 GND.n7937 9.3005
R14218 GND.n7943 GND.n7942 9.3005
R14219 GND.n7940 GND.n126 9.3005
R14220 GND.n7939 GND.n127 9.3005
R14221 GND.n8595 GND.n128 9.3005
R14222 GND.n8594 GND.n8593 9.3005
R14223 GND.n8591 GND.n96 9.3005
R14224 GND.n8590 GND.n97 9.3005
R14225 GND.n8588 GND.n98 9.3005
R14226 GND.n8587 GND.n129 9.3005
R14227 GND.n8584 GND.n130 9.3005
R14228 GND.n8583 GND.n131 9.3005
R14229 GND.n8582 GND.n132 9.3005
R14230 GND.n8233 GND.n133 9.3005
R14231 GND.n8235 GND.n8234 9.3005
R14232 GND.n8236 GND.n147 9.3005
R14233 GND.n8238 GND.n148 9.3005
R14234 GND.n8239 GND.n149 9.3005
R14235 GND.n8242 GND.n8240 9.3005
R14236 GND.n8243 GND.n167 9.3005
R14237 GND.n8245 GND.n168 9.3005
R14238 GND.n8246 GND.n169 9.3005
R14239 GND.n8249 GND.n8247 9.3005
R14240 GND.n8250 GND.n187 9.3005
R14241 GND.n8252 GND.n188 9.3005
R14242 GND.n8253 GND.n189 9.3005
R14243 GND.n8256 GND.n8254 9.3005
R14244 GND.n8257 GND.n209 9.3005
R14245 GND.n8259 GND.n210 9.3005
R14246 GND.n8260 GND.n211 9.3005
R14247 GND.n8263 GND.n8261 9.3005
R14248 GND.n8264 GND.n230 9.3005
R14249 GND.n8266 GND.n231 9.3005
R14250 GND.n8267 GND.n232 9.3005
R14251 GND.n8270 GND.n8268 9.3005
R14252 GND.n8271 GND.n251 9.3005
R14253 GND.n8273 GND.n252 9.3005
R14254 GND.n8274 GND.n253 9.3005
R14255 GND.n8277 GND.n8275 9.3005
R14256 GND.n8278 GND.n272 9.3005
R14257 GND.n8280 GND.n273 9.3005
R14258 GND.n8281 GND.n274 9.3005
R14259 GND.n8284 GND.n8282 9.3005
R14260 GND.n8285 GND.n293 9.3005
R14261 GND.n8287 GND.n294 9.3005
R14262 GND.n8288 GND.n295 9.3005
R14263 GND.n8291 GND.n8289 9.3005
R14264 GND.n8292 GND.n314 9.3005
R14265 GND.n8294 GND.n315 9.3005
R14266 GND.n8295 GND.n316 9.3005
R14267 GND.n8298 GND.n8296 9.3005
R14268 GND.n8299 GND.n335 9.3005
R14269 GND.n8301 GND.n336 9.3005
R14270 GND.n8302 GND.n337 9.3005
R14271 GND.n8305 GND.n8304 9.3005
R14272 GND.n8306 GND.n8225 9.3005
R14273 GND.n8314 GND.n8226 9.3005
R14274 GND.n8313 GND.n8311 9.3005
R14275 GND.n8312 GND.n445 9.3005
R14276 GND.n8331 GND.n446 9.3005
R14277 GND.n7713 GND.n666 9.3005
R14278 GND.n7714 GND.n664 9.3005
R14279 GND.n7722 GND.n665 9.3005
R14280 GND.n7721 GND.n7718 9.3005
R14281 GND.n7720 GND.n7719 9.3005
R14282 GND.n647 GND.n644 9.3005
R14283 GND.n7742 GND.n645 9.3005
R14284 GND.n7741 GND.n7738 9.3005
R14285 GND.n7740 GND.n7739 9.3005
R14286 GND.n627 GND.n624 9.3005
R14287 GND.n7762 GND.n625 9.3005
R14288 GND.n7761 GND.n7758 9.3005
R14289 GND.n7760 GND.n7759 9.3005
R14290 GND.n607 GND.n604 9.3005
R14291 GND.n7782 GND.n605 9.3005
R14292 GND.n7781 GND.n7778 9.3005
R14293 GND.n7780 GND.n7779 9.3005
R14294 GND.n587 GND.n583 9.3005
R14295 GND.n7806 GND.n584 9.3005
R14296 GND.n7805 GND.n585 9.3005
R14297 GND.n7804 GND.n7800 9.3005
R14298 GND.n7803 GND.n7801 9.3005
R14299 GND.n558 GND.n555 9.3005
R14300 GND.n7880 GND.n556 9.3005
R14301 GND.n7879 GND.n7876 9.3005
R14302 GND.n7878 GND.n7877 9.3005
R14303 GND.n539 GND.n536 9.3005
R14304 GND.n7900 GND.n537 9.3005
R14305 GND.n7899 GND.n7896 9.3005
R14306 GND.n7898 GND.n7897 9.3005
R14307 GND.n519 GND.n516 9.3005
R14308 GND.n7920 GND.n517 9.3005
R14309 GND.n7919 GND.n7916 9.3005
R14310 GND.n7918 GND.n7917 9.3005
R14311 GND.n499 GND.n495 9.3005
R14312 GND.n7947 GND.n496 9.3005
R14313 GND.n7946 GND.n497 9.3005
R14314 GND.n7945 GND.n7944 9.3005
R14315 GND.n7943 GND.n125 9.3005
R14316 GND.n8598 GND.n126 9.3005
R14317 GND.n8597 GND.n127 9.3005
R14318 GND.n8596 GND.n8595 9.3005
R14319 GND.n8594 GND.n95 9.3005
R14320 GND.n8628 GND.n96 9.3005
R14321 GND.n8627 GND.n97 9.3005
R14322 GND.n8626 GND.n98 9.3005
R14323 GND.n129 GND.n99 9.3005
R14324 GND.n8228 GND.n130 9.3005
R14325 GND.n8229 GND.n131 9.3005
R14326 GND.n8231 GND.n132 9.3005
R14327 GND.n8233 GND.n8232 9.3005
R14328 GND.n8234 GND.n146 9.3005
R14329 GND.n8570 GND.n147 9.3005
R14330 GND.n8569 GND.n148 9.3005
R14331 GND.n8568 GND.n149 9.3005
R14332 GND.n8240 GND.n150 9.3005
R14333 GND.n8558 GND.n167 9.3005
R14334 GND.n8557 GND.n168 9.3005
R14335 GND.n8556 GND.n169 9.3005
R14336 GND.n8247 GND.n170 9.3005
R14337 GND.n8546 GND.n187 9.3005
R14338 GND.n8545 GND.n188 9.3005
R14339 GND.n8544 GND.n189 9.3005
R14340 GND.n8254 GND.n190 9.3005
R14341 GND.n8534 GND.n209 9.3005
R14342 GND.n8533 GND.n210 9.3005
R14343 GND.n8532 GND.n211 9.3005
R14344 GND.n8261 GND.n212 9.3005
R14345 GND.n8522 GND.n230 9.3005
R14346 GND.n8521 GND.n231 9.3005
R14347 GND.n8520 GND.n232 9.3005
R14348 GND.n8268 GND.n233 9.3005
R14349 GND.n8510 GND.n251 9.3005
R14350 GND.n8509 GND.n252 9.3005
R14351 GND.n8508 GND.n253 9.3005
R14352 GND.n8275 GND.n254 9.3005
R14353 GND.n8498 GND.n272 9.3005
R14354 GND.n8497 GND.n273 9.3005
R14355 GND.n8496 GND.n274 9.3005
R14356 GND.n8282 GND.n275 9.3005
R14357 GND.n8486 GND.n293 9.3005
R14358 GND.n8485 GND.n294 9.3005
R14359 GND.n8484 GND.n295 9.3005
R14360 GND.n8289 GND.n296 9.3005
R14361 GND.n8474 GND.n314 9.3005
R14362 GND.n8473 GND.n315 9.3005
R14363 GND.n8472 GND.n316 9.3005
R14364 GND.n8296 GND.n317 9.3005
R14365 GND.n8462 GND.n335 9.3005
R14366 GND.n8461 GND.n336 9.3005
R14367 GND.n8460 GND.n337 9.3005
R14368 GND.n8305 GND.n338 9.3005
R14369 GND.n8308 GND.n8306 9.3005
R14370 GND.n8309 GND.n8226 9.3005
R14371 GND.n8311 GND.n8310 9.3005
R14372 GND.n447 GND.n445 9.3005
R14373 GND.n8331 GND.n8330 9.3005
R14374 GND.n7713 GND.n7712 9.3005
R14375 GND.n7599 GND.n7598 9.3005
R14376 GND.n7602 GND.n7593 9.3005
R14377 GND.n7603 GND.n7592 9.3005
R14378 GND.n7606 GND.n7591 9.3005
R14379 GND.n7607 GND.n7590 9.3005
R14380 GND.n7610 GND.n7589 9.3005
R14381 GND.n7611 GND.n7588 9.3005
R14382 GND.n7614 GND.n7587 9.3005
R14383 GND.n7615 GND.n7586 9.3005
R14384 GND.n7618 GND.n7585 9.3005
R14385 GND.n7620 GND.n7584 9.3005
R14386 GND.n7621 GND.n7581 9.3005
R14387 GND.n7622 GND.n7579 9.3005
R14388 GND.n7625 GND.n7578 9.3005
R14389 GND.n7626 GND.n7577 9.3005
R14390 GND.n7629 GND.n7576 9.3005
R14391 GND.n7630 GND.n7575 9.3005
R14392 GND.n7633 GND.n7574 9.3005
R14393 GND.n7634 GND.n7573 9.3005
R14394 GND.n7637 GND.n7572 9.3005
R14395 GND.n7638 GND.n7571 9.3005
R14396 GND.n7641 GND.n7570 9.3005
R14397 GND.n7642 GND.n7567 9.3005
R14398 GND.n7645 GND.n7566 9.3005
R14399 GND.n7646 GND.n7565 9.3005
R14400 GND.n7649 GND.n7564 9.3005
R14401 GND.n7650 GND.n7563 9.3005
R14402 GND.n7653 GND.n7562 9.3005
R14403 GND.n7655 GND.n834 9.3005
R14404 GND.n7658 GND.n833 9.3005
R14405 GND.n7660 GND.n832 9.3005
R14406 GND.n7661 GND.n829 9.3005
R14407 GND.n7662 GND.n827 9.3005
R14408 GND.n7665 GND.n826 9.3005
R14409 GND.n7666 GND.n825 9.3005
R14410 GND.n7669 GND.n824 9.3005
R14411 GND.n7670 GND.n823 9.3005
R14412 GND.n7673 GND.n822 9.3005
R14413 GND.n7674 GND.n821 9.3005
R14414 GND.n7677 GND.n820 9.3005
R14415 GND.n7678 GND.n819 9.3005
R14416 GND.n7681 GND.n818 9.3005
R14417 GND.n7682 GND.n815 9.3005
R14418 GND.n7685 GND.n814 9.3005
R14419 GND.n7686 GND.n813 9.3005
R14420 GND.n7689 GND.n812 9.3005
R14421 GND.n7690 GND.n811 9.3005
R14422 GND.n7693 GND.n810 9.3005
R14423 GND.n7695 GND.n809 9.3005
R14424 GND.n7696 GND.n808 9.3005
R14425 GND.n7697 GND.n807 9.3005
R14426 GND.n7698 GND.n806 9.3005
R14427 GND.n7597 GND.n7594 9.3005
R14428 GND.n803 GND.n714 9.3005
R14429 GND.n801 GND.n715 9.3005
R14430 GND.n800 GND.n716 9.3005
R14431 GND.n798 GND.n717 9.3005
R14432 GND.n797 GND.n718 9.3005
R14433 GND.n795 GND.n719 9.3005
R14434 GND.n794 GND.n720 9.3005
R14435 GND.n792 GND.n721 9.3005
R14436 GND.n791 GND.n722 9.3005
R14437 GND.n789 GND.n723 9.3005
R14438 GND.n788 GND.n724 9.3005
R14439 GND.n786 GND.n725 9.3005
R14440 GND.n785 GND.n726 9.3005
R14441 GND.n783 GND.n727 9.3005
R14442 GND.n782 GND.n728 9.3005
R14443 GND.n780 GND.n729 9.3005
R14444 GND.n779 GND.n730 9.3005
R14445 GND.n777 GND.n731 9.3005
R14446 GND.n776 GND.n732 9.3005
R14447 GND.n774 GND.n733 9.3005
R14448 GND.n773 GND.n734 9.3005
R14449 GND.n771 GND.n735 9.3005
R14450 GND.n770 GND.n736 9.3005
R14451 GND.n769 GND.n737 9.3005
R14452 GND.n767 GND.n738 9.3005
R14453 GND.n766 GND.n739 9.3005
R14454 GND.n764 GND.n740 9.3005
R14455 GND.n763 GND.n741 9.3005
R14456 GND.n761 GND.n742 9.3005
R14457 GND.n760 GND.n743 9.3005
R14458 GND.n758 GND.n744 9.3005
R14459 GND.n757 GND.n745 9.3005
R14460 GND.n755 GND.n746 9.3005
R14461 GND.n754 GND.n747 9.3005
R14462 GND.n752 GND.n748 9.3005
R14463 GND.n751 GND.n750 9.3005
R14464 GND.n749 GND.n477 9.3005
R14465 GND.n7960 GND.n478 9.3005
R14466 GND.n7961 GND.n476 9.3005
R14467 GND.n7964 GND.n7963 9.3005
R14468 GND.n7965 GND.n475 9.3005
R14469 GND.n7968 GND.n7966 9.3005
R14470 GND.n7992 GND.n7991 9.3005
R14471 GND.n7995 GND.n7993 9.3005
R14472 GND.n7996 GND.n474 9.3005
R14473 GND.n7999 GND.n7998 9.3005
R14474 GND.n8000 GND.n473 9.3005
R14475 GND.n8003 GND.n8001 9.3005
R14476 GND.n8004 GND.n472 9.3005
R14477 GND.n8007 GND.n8006 9.3005
R14478 GND.n8008 GND.n471 9.3005
R14479 GND.n8011 GND.n8009 9.3005
R14480 GND.n8012 GND.n470 9.3005
R14481 GND.n8015 GND.n8014 9.3005
R14482 GND.n8016 GND.n469 9.3005
R14483 GND.n8019 GND.n8017 9.3005
R14484 GND.n8020 GND.n468 9.3005
R14485 GND.n8023 GND.n8022 9.3005
R14486 GND.n8024 GND.n467 9.3005
R14487 GND.n8027 GND.n8025 9.3005
R14488 GND.n8028 GND.n466 9.3005
R14489 GND.n8031 GND.n8030 9.3005
R14490 GND.n8032 GND.n465 9.3005
R14491 GND.n8035 GND.n8033 9.3005
R14492 GND.n8036 GND.n464 9.3005
R14493 GND.n8039 GND.n8038 9.3005
R14494 GND.n8040 GND.n463 9.3005
R14495 GND.n8043 GND.n8041 9.3005
R14496 GND.n8044 GND.n462 9.3005
R14497 GND.n8047 GND.n8046 9.3005
R14498 GND.n8048 GND.n461 9.3005
R14499 GND.n8051 GND.n8049 9.3005
R14500 GND.n8052 GND.n460 9.3005
R14501 GND.n8055 GND.n8054 9.3005
R14502 GND.n8056 GND.n459 9.3005
R14503 GND.n8059 GND.n8057 9.3005
R14504 GND.n8060 GND.n458 9.3005
R14505 GND.n8063 GND.n8062 9.3005
R14506 GND.n8064 GND.n457 9.3005
R14507 GND.n8066 GND.n8065 9.3005
R14508 GND.n456 GND.n455 9.3005
R14509 GND.n8319 GND.n8318 9.3005
R14510 GND.n8320 GND.n454 9.3005
R14511 GND.n8324 GND.n8321 9.3005
R14512 GND.n8323 GND.n8322 9.3005
R14513 GND.n805 GND.n804 9.3005
R14514 GND.n7990 GND.n82 9.3005
R14515 GND.n2870 GND.n2869 9.3005
R14516 GND.n2873 GND.n2529 9.3005
R14517 GND.n2874 GND.n2528 9.3005
R14518 GND.n2877 GND.n2527 9.3005
R14519 GND.n2878 GND.n2526 9.3005
R14520 GND.n2881 GND.n2525 9.3005
R14521 GND.n2882 GND.n2524 9.3005
R14522 GND.n2885 GND.n2523 9.3005
R14523 GND.n2886 GND.n2522 9.3005
R14524 GND.n2889 GND.n2521 9.3005
R14525 GND.n2891 GND.n2520 9.3005
R14526 GND.n2892 GND.n2517 9.3005
R14527 GND.n2893 GND.n2515 9.3005
R14528 GND.n2896 GND.n2514 9.3005
R14529 GND.n2897 GND.n2513 9.3005
R14530 GND.n2900 GND.n2512 9.3005
R14531 GND.n2901 GND.n2511 9.3005
R14532 GND.n2904 GND.n2510 9.3005
R14533 GND.n2905 GND.n2509 9.3005
R14534 GND.n2908 GND.n2508 9.3005
R14535 GND.n2909 GND.n2507 9.3005
R14536 GND.n2912 GND.n2506 9.3005
R14537 GND.n2913 GND.n2503 9.3005
R14538 GND.n2916 GND.n2502 9.3005
R14539 GND.n2917 GND.n2501 9.3005
R14540 GND.n2920 GND.n2500 9.3005
R14541 GND.n2921 GND.n2499 9.3005
R14542 GND.n2924 GND.n2498 9.3005
R14543 GND.n2925 GND.n2497 9.3005
R14544 GND.n2928 GND.n2496 9.3005
R14545 GND.n2929 GND.n2495 9.3005
R14546 GND.n2932 GND.n2494 9.3005
R14547 GND.n2934 GND.n2493 9.3005
R14548 GND.n2935 GND.n2490 9.3005
R14549 GND.n2936 GND.n2488 9.3005
R14550 GND.n2939 GND.n2487 9.3005
R14551 GND.n2940 GND.n2486 9.3005
R14552 GND.n2943 GND.n2485 9.3005
R14553 GND.n2944 GND.n2484 9.3005
R14554 GND.n2947 GND.n2483 9.3005
R14555 GND.n2948 GND.n2482 9.3005
R14556 GND.n2951 GND.n2481 9.3005
R14557 GND.n2952 GND.n2480 9.3005
R14558 GND.n2955 GND.n2479 9.3005
R14559 GND.n2956 GND.n2476 9.3005
R14560 GND.n2959 GND.n2475 9.3005
R14561 GND.n2960 GND.n2474 9.3005
R14562 GND.n2963 GND.n2473 9.3005
R14563 GND.n2964 GND.n2472 9.3005
R14564 GND.n2967 GND.n2471 9.3005
R14565 GND.n2969 GND.n2470 9.3005
R14566 GND.n2970 GND.n2469 9.3005
R14567 GND.n2971 GND.n2468 9.3005
R14568 GND.n2972 GND.n2467 9.3005
R14569 GND.n2868 GND.n2530 9.3005
R14570 GND.n2570 GND.n2567 9.3005
R14571 GND.n2616 GND.n2615 9.3005
R14572 GND.n2617 GND.n2566 9.3005
R14573 GND.n2714 GND.n2618 9.3005
R14574 GND.n2713 GND.n2619 9.3005
R14575 GND.n2712 GND.n2620 9.3005
R14576 GND.n2711 GND.n2621 9.3005
R14577 GND.n2710 GND.n2622 9.3005
R14578 GND.n2708 GND.n2623 9.3005
R14579 GND.n2707 GND.n2624 9.3005
R14580 GND.n2705 GND.n2625 9.3005
R14581 GND.n2704 GND.n2626 9.3005
R14582 GND.n2702 GND.n2627 9.3005
R14583 GND.n2701 GND.n2628 9.3005
R14584 GND.n2699 GND.n2629 9.3005
R14585 GND.n2698 GND.n2630 9.3005
R14586 GND.n2696 GND.n2631 9.3005
R14587 GND.n2695 GND.n2632 9.3005
R14588 GND.n2693 GND.n2633 9.3005
R14589 GND.n2692 GND.n2634 9.3005
R14590 GND.n2690 GND.n2635 9.3005
R14591 GND.n2689 GND.n2636 9.3005
R14592 GND.n2687 GND.n2637 9.3005
R14593 GND.n2686 GND.n2638 9.3005
R14594 GND.n2684 GND.n2639 9.3005
R14595 GND.n2683 GND.n2640 9.3005
R14596 GND.n2681 GND.n2641 9.3005
R14597 GND.n2680 GND.n2642 9.3005
R14598 GND.n2678 GND.n2643 9.3005
R14599 GND.n2677 GND.n2644 9.3005
R14600 GND.n2675 GND.n2645 9.3005
R14601 GND.n2674 GND.n2646 9.3005
R14602 GND.n2672 GND.n2647 9.3005
R14603 GND.n2671 GND.n2648 9.3005
R14604 GND.n2669 GND.n2649 9.3005
R14605 GND.n2668 GND.n2650 9.3005
R14606 GND.n2666 GND.n2651 9.3005
R14607 GND.n2665 GND.n2652 9.3005
R14608 GND.n2663 GND.n2653 9.3005
R14609 GND.n2662 GND.n2654 9.3005
R14610 GND.n2660 GND.n2655 9.3005
R14611 GND.n2659 GND.n2086 9.3005
R14612 GND.n2196 GND.n2085 9.3005
R14613 GND.n2195 GND.n2093 9.3005
R14614 GND.n2193 GND.n2094 9.3005
R14615 GND.n2192 GND.n2095 9.3005
R14616 GND.n2190 GND.n2096 9.3005
R14617 GND.n2189 GND.n2097 9.3005
R14618 GND.n2187 GND.n2098 9.3005
R14619 GND.n2186 GND.n2099 9.3005
R14620 GND.n2185 GND.n2100 9.3005
R14621 GND.n2183 GND.n2101 9.3005
R14622 GND.n2182 GND.n2102 9.3005
R14623 GND.n2180 GND.n2103 9.3005
R14624 GND.n2179 GND.n2104 9.3005
R14625 GND.n2177 GND.n2105 9.3005
R14626 GND.n2176 GND.n2106 9.3005
R14627 GND.n2174 GND.n2107 9.3005
R14628 GND.n2173 GND.n2108 9.3005
R14629 GND.n2171 GND.n2109 9.3005
R14630 GND.n2170 GND.n2110 9.3005
R14631 GND.n2168 GND.n2111 9.3005
R14632 GND.n2167 GND.n2112 9.3005
R14633 GND.n2165 GND.n2113 9.3005
R14634 GND.n2164 GND.n2114 9.3005
R14635 GND.n2162 GND.n2115 9.3005
R14636 GND.n2161 GND.n2116 9.3005
R14637 GND.n2159 GND.n2117 9.3005
R14638 GND.n2158 GND.n2118 9.3005
R14639 GND.n2156 GND.n2119 9.3005
R14640 GND.n2155 GND.n2120 9.3005
R14641 GND.n2153 GND.n2121 9.3005
R14642 GND.n2152 GND.n2122 9.3005
R14643 GND.n2150 GND.n2123 9.3005
R14644 GND.n2149 GND.n2124 9.3005
R14645 GND.n2147 GND.n2125 9.3005
R14646 GND.n2146 GND.n2126 9.3005
R14647 GND.n2144 GND.n2127 9.3005
R14648 GND.n2143 GND.n2128 9.3005
R14649 GND.n2142 GND.n2129 9.3005
R14650 GND.n2140 GND.n2130 9.3005
R14651 GND.n2139 GND.n2131 9.3005
R14652 GND.n2137 GND.n2132 9.3005
R14653 GND.n2136 GND.n2133 9.3005
R14654 GND.n2134 GND.n1691 9.3005
R14655 GND.n2569 GND.n2568 9.3005
R14656 GND.n5085 GND.n5084 9.3005
R14657 GND.n5086 GND.n2084 9.3005
R14658 GND.n5088 GND.n5087 9.3005
R14659 GND.n2059 GND.n2058 9.3005
R14660 GND.n5110 GND.n5109 9.3005
R14661 GND.n5111 GND.n2057 9.3005
R14662 GND.n5115 GND.n5112 9.3005
R14663 GND.n5114 GND.n5113 9.3005
R14664 GND.n2032 GND.n2031 9.3005
R14665 GND.n5201 GND.n5200 9.3005
R14666 GND.n5202 GND.n2030 9.3005
R14667 GND.n5204 GND.n5203 9.3005
R14668 GND.n2012 GND.n2011 9.3005
R14669 GND.n5221 GND.n5220 9.3005
R14670 GND.n5222 GND.n2010 9.3005
R14671 GND.n5224 GND.n5223 9.3005
R14672 GND.n1992 GND.n1991 9.3005
R14673 GND.n5241 GND.n5240 9.3005
R14674 GND.n5242 GND.n1990 9.3005
R14675 GND.n5244 GND.n5243 9.3005
R14676 GND.n1972 GND.n1971 9.3005
R14677 GND.n5261 GND.n5260 9.3005
R14678 GND.n5262 GND.n1970 9.3005
R14679 GND.n5264 GND.n5263 9.3005
R14680 GND.n1952 GND.n1951 9.3005
R14681 GND.n5281 GND.n5280 9.3005
R14682 GND.n5282 GND.n1950 9.3005
R14683 GND.n5284 GND.n5283 9.3005
R14684 GND.n1932 GND.n1931 9.3005
R14685 GND.n5301 GND.n5300 9.3005
R14686 GND.n5302 GND.n1930 9.3005
R14687 GND.n5304 GND.n5303 9.3005
R14688 GND.n1912 GND.n1911 9.3005
R14689 GND.n5326 GND.n5325 9.3005
R14690 GND.n5327 GND.n1910 9.3005
R14691 GND.n5331 GND.n5328 9.3005
R14692 GND.n5330 GND.n5329 9.3005
R14693 GND.n1885 GND.n1884 9.3005
R14694 GND.n5371 GND.n5370 9.3005
R14695 GND.n5372 GND.n1883 9.3005
R14696 GND.n5376 GND.n5373 9.3005
R14697 GND.n5375 GND.n5374 9.3005
R14698 GND.n1867 GND.n1866 9.3005
R14699 GND.n5391 GND.n5390 9.3005
R14700 GND.n5392 GND.n1865 9.3005
R14701 GND.n5394 GND.n5393 9.3005
R14702 GND.n1864 GND.n1863 9.3005
R14703 GND.n5399 GND.n5398 9.3005
R14704 GND.n5400 GND.n1862 9.3005
R14705 GND.n5402 GND.n5401 9.3005
R14706 GND.n1860 GND.n1859 9.3005
R14707 GND.n5409 GND.n5408 9.3005
R14708 GND.n5410 GND.n1858 9.3005
R14709 GND.n6188 GND.n5411 9.3005
R14710 GND.n6187 GND.n5412 9.3005
R14711 GND.n6186 GND.n5413 9.3005
R14712 GND.n5428 GND.n5414 9.3005
R14713 GND.n6174 GND.n5429 9.3005
R14714 GND.n6173 GND.n5430 9.3005
R14715 GND.n6172 GND.n5431 9.3005
R14716 GND.n5523 GND.n5432 9.3005
R14717 GND.n5524 GND.n5522 9.3005
R14718 GND.n6155 GND.n5525 9.3005
R14719 GND.n6154 GND.n5526 9.3005
R14720 GND.n6153 GND.n5527 9.3005
R14721 GND.n5542 GND.n5528 9.3005
R14722 GND.n6141 GND.n5543 9.3005
R14723 GND.n6140 GND.n5544 9.3005
R14724 GND.n6139 GND.n5545 9.3005
R14725 GND.n5560 GND.n5546 9.3005
R14726 GND.n6127 GND.n5561 9.3005
R14727 GND.n6126 GND.n5562 9.3005
R14728 GND.n6125 GND.n5563 9.3005
R14729 GND.n5578 GND.n5564 9.3005
R14730 GND.n6113 GND.n5579 9.3005
R14731 GND.n6112 GND.n5580 9.3005
R14732 GND.n6111 GND.n5581 9.3005
R14733 GND.n5654 GND.n5582 9.3005
R14734 GND.n5655 GND.n5653 9.3005
R14735 GND.n6094 GND.n5656 9.3005
R14736 GND.n6093 GND.n5657 9.3005
R14737 GND.n6092 GND.n5658 9.3005
R14738 GND.n5673 GND.n5659 9.3005
R14739 GND.n6080 GND.n5674 9.3005
R14740 GND.n6079 GND.n5675 9.3005
R14741 GND.n6078 GND.n5676 9.3005
R14742 GND.n5691 GND.n5677 9.3005
R14743 GND.n6066 GND.n5692 9.3005
R14744 GND.n6065 GND.n5693 9.3005
R14745 GND.n6064 GND.n5694 9.3005
R14746 GND.n5709 GND.n5695 9.3005
R14747 GND.n6052 GND.n5710 9.3005
R14748 GND.n6051 GND.n5711 9.3005
R14749 GND.n6050 GND.n5712 9.3005
R14750 GND.n5785 GND.n5713 9.3005
R14751 GND.n5786 GND.n5784 9.3005
R14752 GND.n6033 GND.n5787 9.3005
R14753 GND.n6032 GND.n5788 9.3005
R14754 GND.n6031 GND.n5789 9.3005
R14755 GND.n5803 GND.n5790 9.3005
R14756 GND.n6019 GND.n5804 9.3005
R14757 GND.n6018 GND.n5805 9.3005
R14758 GND.n6017 GND.n5806 9.3005
R14759 GND.n5821 GND.n5807 9.3005
R14760 GND.n6005 GND.n5822 9.3005
R14761 GND.n6004 GND.n5823 9.3005
R14762 GND.n6003 GND.n5824 9.3005
R14763 GND.n5839 GND.n5825 9.3005
R14764 GND.n5991 GND.n5840 9.3005
R14765 GND.n5990 GND.n5841 9.3005
R14766 GND.n5989 GND.n5842 9.3005
R14767 GND.n5916 GND.n5843 9.3005
R14768 GND.n5917 GND.n5915 9.3005
R14769 GND.n5972 GND.n5918 9.3005
R14770 GND.n5971 GND.n5919 9.3005
R14771 GND.n5970 GND.n5920 9.3005
R14772 GND.n5954 GND.n5921 9.3005
R14773 GND.n5958 GND.n5955 9.3005
R14774 GND.n5957 GND.n5956 9.3005
R14775 GND.n1584 GND.n1583 9.3005
R14776 GND.n6434 GND.n6433 9.3005
R14777 GND.n6435 GND.n1582 9.3005
R14778 GND.n6439 GND.n6436 9.3005
R14779 GND.n6438 GND.n6437 9.3005
R14780 GND.n1553 GND.n1552 9.3005
R14781 GND.n6471 GND.n6470 9.3005
R14782 GND.n6472 GND.n1551 9.3005
R14783 GND.n6479 GND.n6473 9.3005
R14784 GND.n6478 GND.n6474 9.3005
R14785 GND.n6477 GND.n6475 9.3005
R14786 GND.n1515 GND.n1514 9.3005
R14787 GND.n6531 GND.n6530 9.3005
R14788 GND.n6532 GND.n1513 9.3005
R14789 GND.n6542 GND.n6533 9.3005
R14790 GND.n6541 GND.n6534 9.3005
R14791 GND.n6540 GND.n6535 9.3005
R14792 GND.n6537 GND.n6536 9.3005
R14793 GND.n1472 GND.n1471 9.3005
R14794 GND.n6609 GND.n6608 9.3005
R14795 GND.n6610 GND.n1470 9.3005
R14796 GND.n6617 GND.n6611 9.3005
R14797 GND.n6616 GND.n6612 9.3005
R14798 GND.n6615 GND.n6613 9.3005
R14799 GND.n1417 GND.n1416 9.3005
R14800 GND.n6688 GND.n6687 9.3005
R14801 GND.n6689 GND.n1415 9.3005
R14802 GND.n6691 GND.n6690 9.3005
R14803 GND.n1394 GND.n1393 9.3005
R14804 GND.n6717 GND.n6716 9.3005
R14805 GND.n6718 GND.n1392 9.3005
R14806 GND.n6751 GND.n6719 9.3005
R14807 GND.n6750 GND.n6720 9.3005
R14808 GND.n6749 GND.n6721 9.3005
R14809 GND.n6724 GND.n6722 9.3005
R14810 GND.n6744 GND.n6725 9.3005
R14811 GND.n6743 GND.n6726 9.3005
R14812 GND.n6742 GND.n6727 9.3005
R14813 GND.n6730 GND.n6728 9.3005
R14814 GND.n6737 GND.n6731 9.3005
R14815 GND.n6736 GND.n6732 9.3005
R14816 GND.n6735 GND.n6733 9.3005
R14817 GND.n1306 GND.n1305 9.3005
R14818 GND.n6890 GND.n6889 9.3005
R14819 GND.n6891 GND.n1304 9.3005
R14820 GND.n6907 GND.n6892 9.3005
R14821 GND.n6906 GND.n6893 9.3005
R14822 GND.n6905 GND.n6894 9.3005
R14823 GND.n6897 GND.n6895 9.3005
R14824 GND.n6901 GND.n6898 9.3005
R14825 GND.n6900 GND.n6899 9.3005
R14826 GND.n1153 GND.n1152 9.3005
R14827 GND.n7013 GND.n7012 9.3005
R14828 GND.n7014 GND.n1151 9.3005
R14829 GND.n7024 GND.n7015 9.3005
R14830 GND.n7023 GND.n7016 9.3005
R14831 GND.n7022 GND.n7017 9.3005
R14832 GND.n7019 GND.n7018 9.3005
R14833 GND.n1122 GND.n1121 9.3005
R14834 GND.n7059 GND.n7058 9.3005
R14835 GND.n7060 GND.n1120 9.3005
R14836 GND.n7073 GND.n7061 9.3005
R14837 GND.n7072 GND.n7062 9.3005
R14838 GND.n7071 GND.n7063 9.3005
R14839 GND.n7065 GND.n7064 9.3005
R14840 GND.n7067 GND.n7066 9.3005
R14841 GND.n1088 GND.n1087 9.3005
R14842 GND.n7117 GND.n7116 9.3005
R14843 GND.n7118 GND.n1086 9.3005
R14844 GND.n7122 GND.n7119 9.3005
R14845 GND.n7121 GND.n7120 9.3005
R14846 GND.n1063 GND.n1062 9.3005
R14847 GND.n7152 GND.n7151 9.3005
R14848 GND.n7153 GND.n1061 9.3005
R14849 GND.n7160 GND.n7154 9.3005
R14850 GND.n7159 GND.n7155 9.3005
R14851 GND.n7158 GND.n7156 9.3005
R14852 GND.n1039 GND.n1038 9.3005
R14853 GND.n7191 GND.n7190 9.3005
R14854 GND.n7192 GND.n1037 9.3005
R14855 GND.n7205 GND.n7193 9.3005
R14856 GND.n7204 GND.n7194 9.3005
R14857 GND.n7203 GND.n7195 9.3005
R14858 GND.n7197 GND.n7196 9.3005
R14859 GND.n7199 GND.n7198 9.3005
R14860 GND.n1005 GND.n1004 9.3005
R14861 GND.n7249 GND.n7248 9.3005
R14862 GND.n7250 GND.n1003 9.3005
R14863 GND.n7254 GND.n7251 9.3005
R14864 GND.n7253 GND.n7252 9.3005
R14865 GND.n980 GND.n979 9.3005
R14866 GND.n7284 GND.n7283 9.3005
R14867 GND.n7285 GND.n978 9.3005
R14868 GND.n7292 GND.n7286 9.3005
R14869 GND.n7291 GND.n7287 9.3005
R14870 GND.n7290 GND.n7288 9.3005
R14871 GND.n955 GND.n954 9.3005
R14872 GND.n7322 GND.n7321 9.3005
R14873 GND.n7323 GND.n953 9.3005
R14874 GND.n7327 GND.n7324 9.3005
R14875 GND.n7326 GND.n7325 9.3005
R14876 GND.n930 GND.n929 9.3005
R14877 GND.n7357 GND.n7356 9.3005
R14878 GND.n7358 GND.n928 9.3005
R14879 GND.n7360 GND.n7359 9.3005
R14880 GND.n913 GND.n912 9.3005
R14881 GND.n7381 GND.n7380 9.3005
R14882 GND.n7382 GND.n911 9.3005
R14883 GND.n7386 GND.n7383 9.3005
R14884 GND.n7385 GND.n7384 9.3005
R14885 GND.n890 GND.n889 9.3005
R14886 GND.n7417 GND.n7416 9.3005
R14887 GND.n7418 GND.n888 9.3005
R14888 GND.n7420 GND.n7419 9.3005
R14889 GND.n873 GND.n872 9.3005
R14890 GND.n7487 GND.n7486 9.3005
R14891 GND.n7488 GND.n871 9.3005
R14892 GND.n7503 GND.n7489 9.3005
R14893 GND.n7502 GND.n7490 9.3005
R14894 GND.n7501 GND.n7491 9.3005
R14895 GND.n7493 GND.n7492 9.3005
R14896 GND.n7495 GND.n7494 9.3005
R14897 GND.n677 GND.n676 9.3005
R14898 GND.n7705 GND.n7704 9.3005
R14899 GND.n7706 GND.n675 9.3005
R14900 GND.n7708 GND.n7707 9.3005
R14901 GND.n656 GND.n655 9.3005
R14902 GND.n7727 GND.n7726 9.3005
R14903 GND.n7728 GND.n654 9.3005
R14904 GND.n7730 GND.n7729 9.3005
R14905 GND.n636 GND.n635 9.3005
R14906 GND.n7747 GND.n7746 9.3005
R14907 GND.n7748 GND.n634 9.3005
R14908 GND.n7750 GND.n7749 9.3005
R14909 GND.n616 GND.n615 9.3005
R14910 GND.n7767 GND.n7766 9.3005
R14911 GND.n7768 GND.n614 9.3005
R14912 GND.n7770 GND.n7769 9.3005
R14913 GND.n596 GND.n595 9.3005
R14914 GND.n7787 GND.n7786 9.3005
R14915 GND.n7788 GND.n594 9.3005
R14916 GND.n7790 GND.n7789 9.3005
R14917 GND.n575 GND.n574 9.3005
R14918 GND.n7811 GND.n7810 9.3005
R14919 GND.n7812 GND.n573 9.3005
R14920 GND.n7816 GND.n7813 9.3005
R14921 GND.n7815 GND.n7814 9.3005
R14922 GND.n548 GND.n547 9.3005
R14923 GND.n7885 GND.n7884 9.3005
R14924 GND.n7886 GND.n546 9.3005
R14925 GND.n7888 GND.n7887 9.3005
R14926 GND.n528 GND.n527 9.3005
R14927 GND.n7905 GND.n7904 9.3005
R14928 GND.n7906 GND.n526 9.3005
R14929 GND.n7908 GND.n7907 9.3005
R14930 GND.n508 GND.n507 9.3005
R14931 GND.n7925 GND.n7924 9.3005
R14932 GND.n7926 GND.n506 9.3005
R14933 GND.n7928 GND.n7927 9.3005
R14934 GND.n487 GND.n486 9.3005
R14935 GND.n7952 GND.n7951 9.3005
R14936 GND.n7953 GND.n485 9.3005
R14937 GND.n7955 GND.n7954 9.3005
R14938 GND.n117 GND.n116 9.3005
R14939 GND.n8603 GND.n8602 9.3005
R14940 GND.n8604 GND.n115 9.3005
R14941 GND.n8606 GND.n8605 9.3005
R14942 GND.n84 GND.n83 9.3005
R14943 GND.n8633 GND.n8632 9.3005
R14944 GND.n8564 GND.n77 9.3005
R14945 GND.n8563 GND.n158 9.3005
R14946 GND.n8562 GND.n159 9.3005
R14947 GND.n177 GND.n160 9.3005
R14948 GND.n8552 GND.n178 9.3005
R14949 GND.n8551 GND.n179 9.3005
R14950 GND.n8550 GND.n180 9.3005
R14951 GND.n198 GND.n181 9.3005
R14952 GND.n8540 GND.n199 9.3005
R14953 GND.n8539 GND.n200 9.3005
R14954 GND.n8538 GND.n201 9.3005
R14955 GND.n219 GND.n202 9.3005
R14956 GND.n8528 GND.n220 9.3005
R14957 GND.n8527 GND.n221 9.3005
R14958 GND.n8526 GND.n222 9.3005
R14959 GND.n240 GND.n223 9.3005
R14960 GND.n8516 GND.n241 9.3005
R14961 GND.n8515 GND.n242 9.3005
R14962 GND.n8514 GND.n243 9.3005
R14963 GND.n261 GND.n244 9.3005
R14964 GND.n8504 GND.n262 9.3005
R14965 GND.n8503 GND.n263 9.3005
R14966 GND.n8502 GND.n264 9.3005
R14967 GND.n282 GND.n265 9.3005
R14968 GND.n8492 GND.n283 9.3005
R14969 GND.n8491 GND.n284 9.3005
R14970 GND.n8490 GND.n285 9.3005
R14971 GND.n303 GND.n286 9.3005
R14972 GND.n8480 GND.n304 9.3005
R14973 GND.n8479 GND.n305 9.3005
R14974 GND.n8478 GND.n306 9.3005
R14975 GND.n324 GND.n307 9.3005
R14976 GND.n8468 GND.n325 9.3005
R14977 GND.n8467 GND.n326 9.3005
R14978 GND.n8466 GND.n327 9.3005
R14979 GND.n345 GND.n328 9.3005
R14980 GND.n8456 GND.n8455 9.3005
R14981 GND.n4850 GND.n4849 9.3005
R14982 GND.n2411 GND.n2410 9.3005
R14983 GND.n4867 GND.n4866 9.3005
R14984 GND.n4868 GND.n2409 9.3005
R14985 GND.n4870 GND.n4869 9.3005
R14986 GND.n2391 GND.n2390 9.3005
R14987 GND.n4887 GND.n4886 9.3005
R14988 GND.n4888 GND.n2389 9.3005
R14989 GND.n4890 GND.n4889 9.3005
R14990 GND.n2371 GND.n2370 9.3005
R14991 GND.n4907 GND.n4906 9.3005
R14992 GND.n4908 GND.n2369 9.3005
R14993 GND.n4910 GND.n4909 9.3005
R14994 GND.n2350 GND.n2349 9.3005
R14995 GND.n4927 GND.n4926 9.3005
R14996 GND.n4928 GND.n2348 9.3005
R14997 GND.n4930 GND.n4929 9.3005
R14998 GND.n2331 GND.n2330 9.3005
R14999 GND.n4947 GND.n4946 9.3005
R15000 GND.n4948 GND.n2329 9.3005
R15001 GND.n4950 GND.n4949 9.3005
R15002 GND.n2311 GND.n2310 9.3005
R15003 GND.n4967 GND.n4966 9.3005
R15004 GND.n4968 GND.n2309 9.3005
R15005 GND.n4970 GND.n4969 9.3005
R15006 GND.n2291 GND.n2290 9.3005
R15007 GND.n4987 GND.n4986 9.3005
R15008 GND.n4988 GND.n2289 9.3005
R15009 GND.n4990 GND.n4989 9.3005
R15010 GND.n2271 GND.n2270 9.3005
R15011 GND.n5007 GND.n5006 9.3005
R15012 GND.n5008 GND.n2269 9.3005
R15013 GND.n5011 GND.n5010 9.3005
R15014 GND.n5009 GND.n2249 9.3005
R15015 GND.n5032 GND.n2250 9.3005
R15016 GND.n5033 GND.n2079 9.3005
R15017 GND.n4848 GND.n2428 9.3005
R15018 GND.n2430 GND.n2429 9.3005
R15019 GND.n4837 GND.n2977 9.3005
R15020 GND.n4839 GND.n4838 9.3005
R15021 GND.n4836 GND.n2979 9.3005
R15022 GND.n4835 GND.n4834 9.3005
R15023 GND.n2981 GND.n2980 9.3005
R15024 GND.n4828 GND.n4827 9.3005
R15025 GND.n4826 GND.n2983 9.3005
R15026 GND.n4825 GND.n4824 9.3005
R15027 GND.n2985 GND.n2984 9.3005
R15028 GND.n4818 GND.n4817 9.3005
R15029 GND.n4816 GND.n2987 9.3005
R15030 GND.n4815 GND.n4814 9.3005
R15031 GND.n2989 GND.n2988 9.3005
R15032 GND.n4808 GND.n4807 9.3005
R15033 GND.n4806 GND.n2991 9.3005
R15034 GND.n4805 GND.n4804 9.3005
R15035 GND.n2993 GND.n2992 9.3005
R15036 GND.n4798 GND.n4797 9.3005
R15037 GND.n4796 GND.n2995 9.3005
R15038 GND.n4795 GND.n4794 9.3005
R15039 GND.n2997 GND.n2996 9.3005
R15040 GND.n4788 GND.n4787 9.3005
R15041 GND.n4786 GND.n2999 9.3005
R15042 GND.n4785 GND.n4784 9.3005
R15043 GND.n3001 GND.n3000 9.3005
R15044 GND.n4778 GND.n4777 9.3005
R15045 GND.n4776 GND.n3003 9.3005
R15046 GND.n4775 GND.n4774 9.3005
R15047 GND.n3005 GND.n3004 9.3005
R15048 GND.n4768 GND.n4767 9.3005
R15049 GND.n4766 GND.n3007 9.3005
R15050 GND.n4765 GND.n4764 9.3005
R15051 GND.n3009 GND.n3008 9.3005
R15052 GND.n4758 GND.n4757 9.3005
R15053 GND.n4756 GND.n3011 9.3005
R15054 GND.n4755 GND.n4754 9.3005
R15055 GND.n3013 GND.n3012 9.3005
R15056 GND.n4748 GND.n4747 9.3005
R15057 GND.n4746 GND.n3015 9.3005
R15058 GND.n4745 GND.n4744 9.3005
R15059 GND.n3017 GND.n3016 9.3005
R15060 GND.n4738 GND.n4737 9.3005
R15061 GND.n4736 GND.n3019 9.3005
R15062 GND.n4735 GND.n4734 9.3005
R15063 GND.n3021 GND.n3020 9.3005
R15064 GND.n4728 GND.n4727 9.3005
R15065 GND.n4847 GND.n4846 9.3005
R15066 GND.n6291 GND.n1622 9.3005
R15067 GND.n6246 GND.n6245 9.3005
R15068 GND.n6247 GND.n1726 9.3005
R15069 GND.n6249 GND.n6248 9.3005
R15070 GND.n6250 GND.n1723 9.3005
R15071 GND.n6251 GND.n1718 9.3005
R15072 GND.n6253 GND.n6252 9.3005
R15073 GND.n6254 GND.n1717 9.3005
R15074 GND.n6256 GND.n6255 9.3005
R15075 GND.n6257 GND.n1712 9.3005
R15076 GND.n6259 GND.n6258 9.3005
R15077 GND.n6260 GND.n1711 9.3005
R15078 GND.n6262 GND.n6261 9.3005
R15079 GND.n6263 GND.n1706 9.3005
R15080 GND.n6265 GND.n6264 9.3005
R15081 GND.n6266 GND.n1705 9.3005
R15082 GND.n6268 GND.n6267 9.3005
R15083 GND.n6269 GND.n1698 9.3005
R15084 GND.n6271 GND.n6270 9.3005
R15085 GND.n6272 GND.n1697 9.3005
R15086 GND.n6274 GND.n6273 9.3005
R15087 GND.n6275 GND.n1692 9.3005
R15088 GND.n6277 GND.n6276 9.3005
R15089 GND.n6278 GND.n1690 9.3005
R15090 GND.n6280 GND.n6279 9.3005
R15091 GND.n1818 GND.n1817 9.3005
R15092 GND.n1816 GND.n1730 9.3005
R15093 GND.n1815 GND.n1814 9.3005
R15094 GND.n1813 GND.n1731 9.3005
R15095 GND.n1812 GND.n1811 9.3005
R15096 GND.n1810 GND.n1738 9.3005
R15097 GND.n1809 GND.n1808 9.3005
R15098 GND.n1807 GND.n1739 9.3005
R15099 GND.n1806 GND.n1805 9.3005
R15100 GND.n1804 GND.n1744 9.3005
R15101 GND.n1803 GND.n1802 9.3005
R15102 GND.n1801 GND.n1745 9.3005
R15103 GND.n1800 GND.n1799 9.3005
R15104 GND.n1798 GND.n1750 9.3005
R15105 GND.n1797 GND.n1796 9.3005
R15106 GND.n1795 GND.n1751 9.3005
R15107 GND.n1794 GND.n1756 9.3005
R15108 GND.n1793 GND.n1792 9.3005
R15109 GND.n1791 GND.n1759 9.3005
R15110 GND.n1790 GND.n1789 9.3005
R15111 GND.n1788 GND.n1760 9.3005
R15112 GND.n1787 GND.n1786 9.3005
R15113 GND.n1785 GND.n1765 9.3005
R15114 GND.n1784 GND.n1783 9.3005
R15115 GND.n1782 GND.n1766 9.3005
R15116 GND.n1781 GND.n1780 9.3005
R15117 GND.n1779 GND.n1771 9.3005
R15118 GND.n1778 GND.n1777 9.3005
R15119 GND.n1776 GND.n1624 9.3005
R15120 GND.n2861 GND.n2860 9.3005
R15121 GND.n2538 GND.n2537 9.3005
R15122 GND.n2856 GND.n2546 9.3005
R15123 GND.n2855 GND.n2547 9.3005
R15124 GND.n2854 GND.n2548 9.3005
R15125 GND.n2550 GND.n2549 9.3005
R15126 GND.n2850 GND.n2422 9.3005
R15127 GND.n4855 GND.n2421 9.3005
R15128 GND.n4861 GND.n4856 9.3005
R15129 GND.n4860 GND.n4857 9.3005
R15130 GND.n4859 GND.n2402 9.3005
R15131 GND.n4875 GND.n2401 9.3005
R15132 GND.n4881 GND.n4876 9.3005
R15133 GND.n4880 GND.n4877 9.3005
R15134 GND.n4879 GND.n2382 9.3005
R15135 GND.n4895 GND.n2381 9.3005
R15136 GND.n4901 GND.n4896 9.3005
R15137 GND.n4900 GND.n4897 9.3005
R15138 GND.n4899 GND.n2362 9.3005
R15139 GND.n4915 GND.n2361 9.3005
R15140 GND.n4921 GND.n4916 9.3005
R15141 GND.n4920 GND.n4917 9.3005
R15142 GND.n4919 GND.n2342 9.3005
R15143 GND.n4935 GND.n2341 9.3005
R15144 GND.n4941 GND.n4936 9.3005
R15145 GND.n4940 GND.n4937 9.3005
R15146 GND.n4939 GND.n2322 9.3005
R15147 GND.n4955 GND.n2321 9.3005
R15148 GND.n4961 GND.n4956 9.3005
R15149 GND.n4960 GND.n4957 9.3005
R15150 GND.n4959 GND.n2302 9.3005
R15151 GND.n4975 GND.n2301 9.3005
R15152 GND.n4981 GND.n4976 9.3005
R15153 GND.n4980 GND.n4977 9.3005
R15154 GND.n4979 GND.n2282 9.3005
R15155 GND.n4995 GND.n2281 9.3005
R15156 GND.n5001 GND.n4996 9.3005
R15157 GND.n5000 GND.n4997 9.3005
R15158 GND.n4999 GND.n2262 9.3005
R15159 GND.n5016 GND.n2261 9.3005
R15160 GND.n5027 GND.n5017 9.3005
R15161 GND.n5026 GND.n5019 9.3005
R15162 GND.n5025 GND.n5020 9.3005
R15163 GND.n5021 GND.n2239 9.3005
R15164 GND.n5041 GND.n2238 9.3005
R15165 GND.n5047 GND.n5042 9.3005
R15166 GND.n5046 GND.n5043 9.3005
R15167 GND.n5045 GND.n2216 9.3005
R15168 GND.n5058 GND.n2215 9.3005
R15169 GND.n5072 GND.n5059 9.3005
R15170 GND.n5071 GND.n5061 9.3005
R15171 GND.n5070 GND.n5062 9.3005
R15172 GND.n5064 GND.n5063 9.3005
R15173 GND.n5066 GND.n2070 9.3005
R15174 GND.n5093 GND.n2069 9.3005
R15175 GND.n5104 GND.n5094 9.3005
R15176 GND.n5103 GND.n5096 9.3005
R15177 GND.n5102 GND.n5097 9.3005
R15178 GND.n5098 GND.n2042 9.3005
R15179 GND.n5189 GND.n2041 9.3005
R15180 GND.n5195 GND.n5190 9.3005
R15181 GND.n5194 GND.n5191 9.3005
R15182 GND.n5193 GND.n2023 9.3005
R15183 GND.n5209 GND.n2022 9.3005
R15184 GND.n5215 GND.n5210 9.3005
R15185 GND.n5214 GND.n5211 9.3005
R15186 GND.n5213 GND.n2003 9.3005
R15187 GND.n5229 GND.n2002 9.3005
R15188 GND.n5235 GND.n5230 9.3005
R15189 GND.n5234 GND.n5231 9.3005
R15190 GND.n5233 GND.n1983 9.3005
R15191 GND.n5249 GND.n1982 9.3005
R15192 GND.n5255 GND.n5250 9.3005
R15193 GND.n5254 GND.n5251 9.3005
R15194 GND.n5253 GND.n1963 9.3005
R15195 GND.n5269 GND.n1962 9.3005
R15196 GND.n5275 GND.n5270 9.3005
R15197 GND.n5274 GND.n5271 9.3005
R15198 GND.n5273 GND.n1943 9.3005
R15199 GND.n5289 GND.n1942 9.3005
R15200 GND.n5295 GND.n5290 9.3005
R15201 GND.n5294 GND.n5291 9.3005
R15202 GND.n5293 GND.n1923 9.3005
R15203 GND.n5309 GND.n1922 9.3005
R15204 GND.n5320 GND.n5310 9.3005
R15205 GND.n5319 GND.n5312 9.3005
R15206 GND.n5318 GND.n5313 9.3005
R15207 GND.n5314 GND.n1895 9.3005
R15208 GND.n5359 GND.n1894 9.3005
R15209 GND.n5365 GND.n5360 9.3005
R15210 GND.n5364 GND.n5361 9.3005
R15211 GND.n5363 GND.n1876 9.3005
R15212 GND.n5381 GND.n1875 9.3005
R15213 GND.n5384 GND.n5383 9.3005
R15214 GND.n5382 GND.n1625 9.3005
R15215 GND.n6289 GND.n1626 9.3005
R15216 GND.n2862 GND.n2533 9.3005
R15217 GND.n2860 GND.n2859 9.3005
R15218 GND.n2858 GND.n2538 9.3005
R15219 GND.n2857 GND.n2856 9.3005
R15220 GND.n2855 GND.n2545 9.3005
R15221 GND.n2854 GND.n2853 9.3005
R15222 GND.n2852 GND.n2550 9.3005
R15223 GND.n2851 GND.n2850 9.3005
R15224 GND.n2421 GND.n2419 9.3005
R15225 GND.n4862 GND.n4861 9.3005
R15226 GND.n4860 GND.n2420 9.3005
R15227 GND.n4859 GND.n4858 9.3005
R15228 GND.n2401 GND.n2399 9.3005
R15229 GND.n4882 GND.n4881 9.3005
R15230 GND.n4880 GND.n2400 9.3005
R15231 GND.n4879 GND.n4878 9.3005
R15232 GND.n2381 GND.n2379 9.3005
R15233 GND.n4902 GND.n4901 9.3005
R15234 GND.n4900 GND.n2380 9.3005
R15235 GND.n4899 GND.n4898 9.3005
R15236 GND.n2361 GND.n2359 9.3005
R15237 GND.n4922 GND.n4921 9.3005
R15238 GND.n4920 GND.n2360 9.3005
R15239 GND.n4919 GND.n4918 9.3005
R15240 GND.n2341 GND.n2339 9.3005
R15241 GND.n4942 GND.n4941 9.3005
R15242 GND.n4940 GND.n2340 9.3005
R15243 GND.n4939 GND.n4938 9.3005
R15244 GND.n2321 GND.n2319 9.3005
R15245 GND.n4962 GND.n4961 9.3005
R15246 GND.n4960 GND.n2320 9.3005
R15247 GND.n4959 GND.n4958 9.3005
R15248 GND.n2301 GND.n2299 9.3005
R15249 GND.n4982 GND.n4981 9.3005
R15250 GND.n4980 GND.n2300 9.3005
R15251 GND.n4979 GND.n4978 9.3005
R15252 GND.n2281 GND.n2279 9.3005
R15253 GND.n5002 GND.n5001 9.3005
R15254 GND.n5000 GND.n2280 9.3005
R15255 GND.n4999 GND.n4998 9.3005
R15256 GND.n2261 GND.n2259 9.3005
R15257 GND.n5028 GND.n5027 9.3005
R15258 GND.n5026 GND.n2260 9.3005
R15259 GND.n5025 GND.n5024 9.3005
R15260 GND.n5023 GND.n5021 9.3005
R15261 GND.n2238 GND.n2236 9.3005
R15262 GND.n5048 GND.n5047 9.3005
R15263 GND.n5046 GND.n2237 9.3005
R15264 GND.n5045 GND.n5044 9.3005
R15265 GND.n2215 GND.n2213 9.3005
R15266 GND.n5073 GND.n5072 9.3005
R15267 GND.n5071 GND.n2214 9.3005
R15268 GND.n5070 GND.n5069 9.3005
R15269 GND.n5068 GND.n5064 9.3005
R15270 GND.n5067 GND.n5066 9.3005
R15271 GND.n2069 GND.n2067 9.3005
R15272 GND.n5105 GND.n5104 9.3005
R15273 GND.n5103 GND.n2068 9.3005
R15274 GND.n5102 GND.n5101 9.3005
R15275 GND.n5100 GND.n5098 9.3005
R15276 GND.n2041 GND.n2039 9.3005
R15277 GND.n5196 GND.n5195 9.3005
R15278 GND.n5194 GND.n2040 9.3005
R15279 GND.n5193 GND.n5192 9.3005
R15280 GND.n2022 GND.n2020 9.3005
R15281 GND.n5216 GND.n5215 9.3005
R15282 GND.n5214 GND.n2021 9.3005
R15283 GND.n5213 GND.n5212 9.3005
R15284 GND.n2002 GND.n2000 9.3005
R15285 GND.n5236 GND.n5235 9.3005
R15286 GND.n5234 GND.n2001 9.3005
R15287 GND.n5233 GND.n5232 9.3005
R15288 GND.n1982 GND.n1980 9.3005
R15289 GND.n5256 GND.n5255 9.3005
R15290 GND.n5254 GND.n1981 9.3005
R15291 GND.n5253 GND.n5252 9.3005
R15292 GND.n1962 GND.n1960 9.3005
R15293 GND.n5276 GND.n5275 9.3005
R15294 GND.n5274 GND.n1961 9.3005
R15295 GND.n5273 GND.n5272 9.3005
R15296 GND.n1942 GND.n1940 9.3005
R15297 GND.n5296 GND.n5295 9.3005
R15298 GND.n5294 GND.n1941 9.3005
R15299 GND.n5293 GND.n5292 9.3005
R15300 GND.n1922 GND.n1920 9.3005
R15301 GND.n5321 GND.n5320 9.3005
R15302 GND.n5319 GND.n1921 9.3005
R15303 GND.n5318 GND.n5317 9.3005
R15304 GND.n5316 GND.n5314 9.3005
R15305 GND.n1894 GND.n1892 9.3005
R15306 GND.n5366 GND.n5365 9.3005
R15307 GND.n5364 GND.n1893 9.3005
R15308 GND.n5363 GND.n5362 9.3005
R15309 GND.n1875 GND.n1874 9.3005
R15310 GND.n5385 GND.n5384 9.3005
R15311 GND.n1627 GND.n1625 9.3005
R15312 GND.n6289 GND.n6288 9.3005
R15313 GND.n2539 GND.n2533 9.3005
R15314 GND.n2601 GND.n2575 9.3005
R15315 GND.n2600 GND.n2599 9.3005
R15316 GND.n2598 GND.n2579 9.3005
R15317 GND.n2597 GND.n2596 9.3005
R15318 GND.n2593 GND.n2582 9.3005
R15319 GND.n2592 GND.n2591 9.3005
R15320 GND.n2590 GND.n2583 9.3005
R15321 GND.n2589 GND.n2588 9.3005
R15322 GND.n2535 GND.n2534 9.3005
R15323 GND.n2866 GND.n2865 9.3005
R15324 GND.n2603 GND.n2602 9.3005
R15325 GND.n2607 GND.n2574 9.3005
R15326 GND.n2609 GND.n2608 9.3005
R15327 GND.n2558 GND.n2557 9.3005
R15328 GND.n2719 GND.n2718 9.3005
R15329 GND.n2720 GND.n2555 9.3005
R15330 GND.n2846 GND.n2845 9.3005
R15331 GND.n2844 GND.n2556 9.3005
R15332 GND.n2843 GND.n2842 9.3005
R15333 GND.n2841 GND.n2721 9.3005
R15334 GND.n2840 GND.n2839 9.3005
R15335 GND.n2838 GND.n2724 9.3005
R15336 GND.n2837 GND.n2836 9.3005
R15337 GND.n2835 GND.n2725 9.3005
R15338 GND.n2834 GND.n2833 9.3005
R15339 GND.n2832 GND.n2728 9.3005
R15340 GND.n2831 GND.n2830 9.3005
R15341 GND.n2829 GND.n2729 9.3005
R15342 GND.n2828 GND.n2827 9.3005
R15343 GND.n2826 GND.n2732 9.3005
R15344 GND.n2825 GND.n2824 9.3005
R15345 GND.n2823 GND.n2733 9.3005
R15346 GND.n2822 GND.n2821 9.3005
R15347 GND.n2820 GND.n2736 9.3005
R15348 GND.n2819 GND.n2818 9.3005
R15349 GND.n2817 GND.n2737 9.3005
R15350 GND.n2816 GND.n2815 9.3005
R15351 GND.n2814 GND.n2740 9.3005
R15352 GND.n2813 GND.n2812 9.3005
R15353 GND.n2811 GND.n2741 9.3005
R15354 GND.n2810 GND.n2809 9.3005
R15355 GND.n2808 GND.n2744 9.3005
R15356 GND.n2807 GND.n2806 9.3005
R15357 GND.n2805 GND.n2745 9.3005
R15358 GND.n2804 GND.n2803 9.3005
R15359 GND.n2802 GND.n2748 9.3005
R15360 GND.n2801 GND.n2800 9.3005
R15361 GND.n2799 GND.n2749 9.3005
R15362 GND.n2798 GND.n2797 9.3005
R15363 GND.n2796 GND.n2752 9.3005
R15364 GND.n2795 GND.n2794 9.3005
R15365 GND.n2793 GND.n2753 9.3005
R15366 GND.n2792 GND.n2791 9.3005
R15367 GND.n2790 GND.n2757 9.3005
R15368 GND.n2789 GND.n2788 9.3005
R15369 GND.n2787 GND.n2758 9.3005
R15370 GND.n2786 GND.n2785 9.3005
R15371 GND.n2784 GND.n2761 9.3005
R15372 GND.n2606 GND.n2605 9.3005
R15373 GND.n2783 GND.n2762 9.3005
R15374 GND.n6449 GND.n1571 9.18926
R15375 GND.n6510 GND.n1519 9.18926
R15376 GND.n6589 GND.n1467 9.18926
R15377 GND.n6672 GND.n1397 9.18926
R15378 GND.n6821 GND.n1355 9.18926
R15379 GND.n1297 GND.n1295 9.18926
R15380 GND.n4992 GND.t19 8.48243
R15381 GND.n5198 GND.t30 8.48243
R15382 GND.n5494 GND.n5491 8.48243
R15383 GND.n6151 GND.n5530 8.48243
R15384 GND.n5623 GND.n5620 8.48243
R15385 GND.n6090 GND.n5661 8.48243
R15386 GND.n5756 GND.n5753 8.48243
R15387 GND.n6029 GND.n5792 8.48243
R15388 GND.n5887 GND.n5884 8.48243
R15389 GND.n5968 GND.n5923 8.48243
R15390 GND.n6441 GND.n1571 8.48243
R15391 GND.n6510 GND.n6509 8.48243
R15392 GND.n6589 GND.n6588 8.48243
R15393 GND.n6672 GND.n1387 8.48243
R15394 GND.n6740 GND.n1355 8.48243
R15395 GND.n1297 GND.n1290 8.48243
R15396 GND.n7026 GND.n1141 8.48243
R15397 GND.n7088 GND.n1101 8.48243
R15398 GND.n7142 GND.n1071 8.48243
R15399 GND.n7214 GND.n1029 8.48243
R15400 GND.n7256 GND.n993 8.48243
R15401 GND.n959 GND.n949 8.48243
R15402 GND.n7370 GND.n919 8.48243
R15403 GND.n7484 GND.n875 8.48243
R15404 GND.n7949 GND.t44 8.48243
R15405 GND.n192 GND.t23 8.48243
R15406 GND.n8640 GND.n8639 8.14362
R15407 GND.n2783 GND.n29 8.14362
R15408 GND.n6408 GND.t93 8.12901
R15409 GND.n6806 GND.t130 8.12901
R15410 GND.n6502 GND.n1530 7.7756
R15411 GND.n1462 GND.n1461 7.7756
R15412 GND.n6707 GND.n1401 7.7756
R15413 GND.n6850 GND.n6849 7.7756
R15414 GND.n1855 GND.n1852 7.06877
R15415 GND.n6144 GND.n6143 7.06877
R15416 GND.n5556 GND.n5550 7.06877
R15417 GND.n6083 GND.n6082 7.06877
R15418 GND.n5687 GND.n5681 7.06877
R15419 GND.n6022 GND.n6021 7.06877
R15420 GND.n5817 GND.n5811 7.06877
R15421 GND.n5961 GND.n5960 7.06877
R15422 GND.n6424 GND.n1592 7.06877
R15423 GND.n6431 GND.n6430 7.06877
R15424 GND.n6519 GND.n6518 7.06877
R15425 GND.n6574 GND.n1485 7.06877
R15426 GND.n6761 GND.n1383 7.06877
R15427 GND.n1365 GND.n1360 7.06877
R15428 GND.n1175 GND.n1166 7.06877
R15429 GND.n1167 GND.n1161 7.06877
R15430 GND.n7010 GND.n7009 7.06877
R15431 GND.n7107 GND.n7106 7.06877
R15432 GND.n7124 GND.n1076 7.06877
R15433 GND.n7220 GND.n1018 7.06877
R15434 GND.n7246 GND.n7245 7.06877
R15435 GND.n7336 GND.n945 7.06877
R15436 GND.n934 GND.n924 7.06877
R15437 GND.n7506 GND.n7505 7.06877
R15438 GND.n6237 GND.n1846 6.71536
R15439 GND.n7556 GND.n839 6.71536
R15440 GND.n6482 GND.n1544 6.36195
R15441 GND.n1600 GND.n1547 6.36195
R15442 GND.n1458 GND.n1419 6.36195
R15443 GND.n1452 GND.n1421 6.36195
R15444 GND.n1332 GND.n1314 6.36195
R15445 GND.n1315 GND.n1308 6.36195
R15446 GND.n12 GND.n7 6.34605
R15447 GND.t93 GND.n1563 6.00853
R15448 GND.n6909 GND.t130 6.00853
R15449 GND.n5610 GND.n5607 5.65512
R15450 GND.n6137 GND.n5548 5.65512
R15451 GND.n5743 GND.n5740 5.65512
R15452 GND.n6076 GND.n5679 5.65512
R15453 GND.n5874 GND.n5871 5.65512
R15454 GND.n6015 GND.n5809 5.65512
R15455 GND.n5952 GND.n5951 5.65512
R15456 GND.n6424 GND.n6423 5.65512
R15457 GND.t4 GND.n6457 5.65512
R15458 GND.n6582 GND.n1490 5.65512
R15459 GND.n6580 GND.n1482 5.65512
R15460 GND.n6773 GND.n1370 5.65512
R15461 GND.n6746 GND.n1373 5.65512
R15462 GND.n6872 GND.t2 5.65512
R15463 GND.n1168 GND.n1167 5.65512
R15464 GND.n7003 GND.n7002 5.65512
R15465 GND.n7114 GND.n7113 5.65512
R15466 GND.n1092 GND.n1082 5.65512
R15467 GND.n1019 GND.n1013 5.65512
R15468 GND.n7239 GND.n7238 5.65512
R15469 GND.n7347 GND.n938 5.65512
R15470 GND.n7354 GND.n932 5.65512
R15471 GND.n28 GND.n3 5.6176
R15472 GND.n12 GND.n11 5.5551
R15473 GND.n17 GND.n16 5.5551
R15474 GND.n22 GND.n21 5.5551
R15475 GND.n27 GND.n26 5.5551
R15476 GND.n41 GND.n36 5.42938
R15477 GND.n6300 GND.n6299 5.23686
R15478 GND.n6942 GND.n6941 5.23686
R15479 GND.n5753 GND.t81 4.94829
R15480 GND.t1 GND.n5910 4.94829
R15481 GND.n6467 GND.n6466 4.94829
R15482 GND.n6496 GND.n6495 4.94829
R15483 GND.n6645 GND.n1435 4.94829
R15484 GND.n6694 GND.n1411 4.94829
R15485 GND.n6857 GND.n6856 4.94829
R15486 GND.n6886 GND.n1310 4.94829
R15487 GND.t0 GND.n7039 4.94829
R15488 GND.n1029 GND.t3 4.94829
R15489 GND.n29 GND.n28 4.93126
R15490 GND.n8640 GND.n61 4.93126
R15491 GND.n6345 GND.n6292 4.74817
R15492 GND.n6350 GND.n6293 4.74817
R15493 GND.n6355 GND.n6294 4.74817
R15494 GND.n6360 GND.n6295 4.74817
R15495 GND.n6300 GND.n6296 4.74817
R15496 GND.n6368 GND.n1615 4.74817
R15497 GND.n6938 GND.n6937 4.74817
R15498 GND.n1199 GND.n1196 4.74817
R15499 GND.n1278 GND.n1276 4.74817
R15500 GND.n6949 GND.n6948 4.74817
R15501 GND.n1282 GND.n1280 4.74817
R15502 GND.n1224 GND.n1200 4.74817
R15503 GND.n1220 GND.n1201 4.74817
R15504 GND.n1216 GND.n1202 4.74817
R15505 GND.n1212 GND.n1203 4.74817
R15506 GND.n1209 GND.n1203 4.74817
R15507 GND.n1213 GND.n1202 4.74817
R15508 GND.n1217 GND.n1201 4.74817
R15509 GND.n1221 GND.n1200 4.74817
R15510 GND.n6957 GND.n1199 4.74817
R15511 GND.n6955 GND.n1276 4.74817
R15512 GND.n6950 GND.n6949 4.74817
R15513 GND.n6947 GND.n1280 4.74817
R15514 GND.n6937 GND.n6936 4.74817
R15515 GND.n7972 GND.n7970 4.74817
R15516 GND.n7975 GND.n7974 4.74817
R15517 GND.n7980 GND.n7979 4.74817
R15518 GND.n7984 GND.n7983 4.74817
R15519 GND.n7988 GND.n7987 4.74817
R15520 GND.n7970 GND.n7969 4.74817
R15521 GND.n7974 GND.n7973 4.74817
R15522 GND.n7979 GND.n7978 4.74817
R15523 GND.n7983 GND.n7982 4.74817
R15524 GND.n7987 GND.n7986 4.74817
R15525 GND.n2244 GND.n2091 4.74817
R15526 GND.n2230 GND.n2090 4.74817
R15527 GND.n2221 GND.n2089 4.74817
R15528 GND.n2207 GND.n2088 4.74817
R15529 GND.n2092 GND.n2087 4.74817
R15530 GND.n2656 GND.n2091 4.74817
R15531 GND.n2243 GND.n2090 4.74817
R15532 GND.n2229 GND.n2089 4.74817
R15533 GND.n2220 GND.n2088 4.74817
R15534 GND.n2206 GND.n2087 4.74817
R15535 GND.n5034 GND.n2078 4.74817
R15536 GND.n5053 GND.n2083 4.74817
R15537 GND.n2203 GND.n2082 4.74817
R15538 GND.n5078 GND.n2081 4.74817
R15539 GND.n2080 GND.n2077 4.74817
R15540 GND.n8622 GND.n81 4.74817
R15541 GND.n80 GND.n75 4.74817
R15542 GND.n8634 GND.n76 4.74817
R15543 GND.n8575 GND.n79 4.74817
R15544 GND.n157 GND.n78 4.74817
R15545 GND.n5036 GND.n2078 4.74817
R15546 GND.n2226 GND.n2083 4.74817
R15547 GND.n5054 GND.n2082 4.74817
R15548 GND.n2204 GND.n2081 4.74817
R15549 GND.n5079 GND.n2080 4.74817
R15550 GND.n85 GND.n81 4.74817
R15551 GND.n8621 GND.n80 4.74817
R15552 GND.n8635 GND.n8634 4.74817
R15553 GND.n8577 GND.n79 4.74817
R15554 GND.n8574 GND.n78 4.74817
R15555 GND.n1638 GND.n1618 4.74817
R15556 GND.n1639 GND.n1619 4.74817
R15557 GND.n1644 GND.n1620 4.74817
R15558 GND.n1649 GND.n1621 4.74817
R15559 GND.n1643 GND.n1619 4.74817
R15560 GND.n1648 GND.n1620 4.74817
R15561 GND.n1652 GND.n1621 4.74817
R15562 GND.n6368 GND.n6367 4.74817
R15563 GND.n6361 GND.n6296 4.74817
R15564 GND.n6356 GND.n6295 4.74817
R15565 GND.n6351 GND.n6294 4.74817
R15566 GND.n6346 GND.n6293 4.74817
R15567 GND.n6341 GND.n6292 4.74817
R15568 GND.n61 GND.n60 4.70093
R15569 GND.n41 GND.n40 4.63843
R15570 GND.n46 GND.n45 4.63843
R15571 GND.n51 GND.n50 4.63843
R15572 GND.n56 GND.n55 4.63843
R15573 GND.n7654 GND.n7561 4.6132
R15574 GND.n6242 GND.n1727 4.6132
R15575 GND.n4852 GND.t89 4.24146
R15576 GND.n5357 GND.t126 4.24146
R15577 GND.n6191 GND.n6190 4.24146
R15578 GND.n5538 GND.n5532 4.24146
R15579 GND.n6130 GND.n6129 4.24146
R15580 GND.n5669 GND.n5663 4.24146
R15581 GND.n6069 GND.n6068 4.24146
R15582 GND.n5800 GND.n5794 4.24146
R15583 GND.n6008 GND.n6007 4.24146
R15584 GND.n5931 GND.n5925 4.24146
R15585 GND.n6416 GND.n6415 4.24146
R15586 GND.n6544 GND.n1510 4.24146
R15587 GND.n6606 GND.n1474 4.24146
R15588 GND.n6753 GND.n1380 4.24146
R15589 GND.n6789 GND.n1349 4.24146
R15590 GND.n6985 GND.n1172 4.24146
R15591 GND.n1157 GND.n1147 4.24146
R15592 GND.n1102 GND.n1096 4.24146
R15593 GND.n7131 GND.n1078 4.24146
R15594 GND.n7221 GND.n1023 4.24146
R15595 GND.n1009 GND.n999 4.24146
R15596 GND.n7329 GND.n943 4.24146
R15597 GND.n7363 GND.n7362 4.24146
R15598 GND.n7507 GND.n866 4.24146
R15599 GND.t134 GND.n629 4.24146
R15600 GND.t110 GND.n332 4.24146
R15601 GND.n1208 GND.n1204 4.05147
R15602 GND.n1658 GND.n1623 4.05147
R15603 GND.n32 GND.n30 4.02701
R15604 GND.n32 GND.n31 3.53792
R15605 GND.n6408 GND.n6407 3.53464
R15606 GND.n6504 GND.n1517 3.53464
R15607 GND.n6635 GND.n6634 3.53464
R15608 GND.n6705 GND.n6704 3.53464
R15609 GND.n6841 GND.n6840 3.53464
R15610 GND.n6807 GND.n6806 3.53464
R15611 GND.n6184 GND.n5416 2.82781
R15612 GND.n5597 GND.n5594 2.82781
R15613 GND.n6123 GND.n5566 2.82781
R15614 GND.n5730 GND.n5727 2.82781
R15615 GND.n6062 GND.n5697 2.82781
R15616 GND.n5860 GND.n5857 2.82781
R15617 GND.n6001 GND.n5827 2.82781
R15618 GND.n5940 GND.n5937 2.82781
R15619 GND.n6448 GND.n1574 2.82781
R15620 GND.n6528 GND.n6527 2.82781
R15621 GND.n6620 GND.n6619 2.82781
R15622 GND.n6714 GND.n6713 2.82781
R15623 GND.n6822 GND.n1342 2.82781
R15624 GND.n6917 GND.n1294 2.82781
R15625 GND.n7033 GND.n1143 2.82781
R15626 GND.n7089 GND.n1106 2.82781
R15627 GND.n7149 GND.n1065 2.82781
R15628 GND.n7207 GND.n1027 2.82781
R15629 GND.n7263 GND.n995 2.82781
R15630 GND.n7319 GND.n7318 2.82781
R15631 GND.n7378 GND.n915 2.82781
R15632 GND.n7430 GND.n879 2.82781
R15633 GND.n1274 GND.n1204 2.62577
R15634 GND.n6291 GND.n1623 2.62577
R15635 GND GND.n29 2.29567
R15636 GND.n1274 GND.n1203 2.27742
R15637 GND.n1274 GND.n1202 2.27742
R15638 GND.n1274 GND.n1201 2.27742
R15639 GND.n1274 GND.n1200 2.27742
R15640 GND.n1275 GND.n1199 2.27742
R15641 GND.n1276 GND.n1275 2.27742
R15642 GND.n6949 GND.n1275 2.27742
R15643 GND.n1280 GND.n1275 2.27742
R15644 GND.n6937 GND.n1275 2.27742
R15645 GND.n7970 GND.n82 2.27742
R15646 GND.n7974 GND.n82 2.27742
R15647 GND.n7979 GND.n82 2.27742
R15648 GND.n7983 GND.n82 2.27742
R15649 GND.n7987 GND.n82 2.27742
R15650 GND.n5085 GND.n2091 2.27742
R15651 GND.n5085 GND.n2090 2.27742
R15652 GND.n5085 GND.n2089 2.27742
R15653 GND.n5085 GND.n2088 2.27742
R15654 GND.n5085 GND.n2087 2.27742
R15655 GND.n5086 GND.n2083 2.27742
R15656 GND.n5086 GND.n2082 2.27742
R15657 GND.n5086 GND.n2081 2.27742
R15658 GND.n5086 GND.n2080 2.27742
R15659 GND.n8633 GND.n81 2.27742
R15660 GND.n8633 GND.n80 2.27742
R15661 GND.n8634 GND.n8633 2.27742
R15662 GND.n8633 GND.n79 2.27742
R15663 GND.n8633 GND.n78 2.27742
R15664 GND.n5086 GND.n2078 2.27742
R15665 GND.n6291 GND.n1618 2.27742
R15666 GND.n6291 GND.n1619 2.27742
R15667 GND.n6291 GND.n1620 2.27742
R15668 GND.n6291 GND.n1621 2.27742
R15669 GND.n6369 GND.n6368 2.27742
R15670 GND.n6369 GND.n6296 2.27742
R15671 GND.n6369 GND.n6295 2.27742
R15672 GND.n6369 GND.n6294 2.27742
R15673 GND.n6369 GND.n6293 2.27742
R15674 GND.n6369 GND.n6292 2.27742
R15675 GND.n6442 GND.n1578 2.12098
R15676 GND.n6458 GND.t4 2.12098
R15677 GND.n6545 GND.n1508 2.12098
R15678 GND.n6605 GND.n1476 2.12098
R15679 GND.n6755 GND.n6754 2.12098
R15680 GND.n6829 GND.n6828 2.12098
R15681 GND.n6910 GND.t2 2.12098
R15682 GND.n6925 GND.n6924 2.12098
R15683 GND.n8641 GND.n8640 2.04453
R15684 GND.n7 GND.n5 1.83383
R15685 GND.n11 GND.n9 1.83383
R15686 GND.n16 GND.n14 1.83383
R15687 GND.n21 GND.n19 1.83383
R15688 GND.n26 GND.n24 1.83383
R15689 GND.n3 GND.n1 1.83383
R15690 GND.n36 GND.n35 1.83383
R15691 GND.n40 GND.n39 1.83383
R15692 GND.n45 GND.n44 1.83383
R15693 GND.n50 GND.n49 1.83383
R15694 GND.n55 GND.n54 1.83383
R15695 GND.n60 GND.n59 1.83383
R15696 GND.n6177 GND.n6176 1.41415
R15697 GND.n5519 GND.n5516 1.41415
R15698 GND.n6116 GND.n6115 1.41415
R15699 GND.n5648 GND.n5637 1.41415
R15700 GND.n6055 GND.n6054 1.41415
R15701 GND.n5779 GND.n5770 1.41415
R15702 GND.n5994 GND.n5993 1.41415
R15703 GND.n5910 GND.n5901 1.41415
R15704 GND.n6468 GND.n1555 1.41415
R15705 GND.n1596 GND.n1537 1.41415
R15706 GND.n6628 GND.n1434 1.41415
R15707 GND.n6693 GND.n1413 1.41415
R15708 GND.n6848 GND.n1329 1.41415
R15709 GND.n6873 GND.n1320 1.41415
R15710 GND.n7039 GND.n1131 1.41415
R15711 GND.n7075 GND.n1110 1.41415
R15712 GND.n7163 GND.n7162 1.41415
R15713 GND.n7188 GND.n7187 1.41415
R15714 GND.n7281 GND.n982 1.41415
R15715 GND.n969 GND.n963 1.41415
R15716 GND.n7389 GND.n7388 1.41415
R15717 GND.n894 GND.n884 1.41415
R15718 GND.n6367 GND.n6299 1.35808
R15719 GND.n6941 GND.n6938 1.35808
R15720 GND.n7520 GND.n7519 1.24928
R15721 GND.n7441 GND.n7436 1.24928
R15722 GND.n5450 GND.n5449 1.24928
R15723 GND.n6201 GND.n6200 1.24928
R15724 GND.n28 GND.n27 1.13125
R15725 GND.n61 GND.n56 1.13125
R15726 GND.n6509 GND.t86 1.06074
R15727 GND.n6740 GND.t82 1.06074
R15728 GND.n17 GND.n12 0.791448
R15729 GND.n22 GND.n17 0.791448
R15730 GND.n27 GND.n22 0.791448
R15731 GND.n46 GND.n41 0.791448
R15732 GND.n51 GND.n46 0.791448
R15733 GND.n56 GND.n51 0.791448
R15734 GND.n6242 GND.n1818 0.776258
R15735 GND.n7654 GND.n7653 0.776258
R15736 GND.n1275 GND.n1274 0.736217
R15737 GND.n6369 GND.n6291 0.736217
R15738 GND.n6021 GND.t6 0.707327
R15739 GND.n6553 GND.n1502 0.707327
R15740 GND.t84 GND.n6597 0.707327
R15741 GND.n6665 GND.t5 0.707327
R15742 GND.n6780 GND.n1364 0.707327
R15743 GND.t7 GND.n7124 0.707327
R15744 GND.n8322 GND.n386 0.5005
R15745 GND.n806 GND.n805 0.5005
R15746 GND.n6279 GND.n1691 0.5005
R15747 GND.n2568 GND.n2467 0.5005
R15748 GND.n4727 GND.n4726 0.497451
R15749 GND.n3964 GND.n3963 0.497451
R15750 GND.n8455 GND.n8454 0.497451
R15751 GND.n4848 GND.n4847 0.497451
R15752 GND.n6981 GND.n6980 0.494402
R15753 GND.n6312 GND.n6310 0.494402
R15754 GND.n6370 GND.n1611 0.494402
R15755 GND.n6930 GND.n6929 0.494402
R15756 GND.n8214 GND.n8183 0.485256
R15757 GND.n2606 GND.n2603 0.485256
R15758 GND.n8633 GND.n82 0.407
R15759 GND.n5086 GND.n5085 0.407
R15760 GND.n6282 GND.n1637 0.353914
R15761 GND.n6619 GND.t186 0.353914
R15762 GND.n6714 GND.t8 0.353914
R15763 GND.n7702 GND.n7701 0.353914
R15764 GND.n7559 GND.n835 0.312695
R15765 GND.n7559 GND.n836 0.312695
R15766 GND.n6241 GND.n1820 0.312695
R15767 GND.n6241 GND.n6240 0.312695
R15768 GND.n6291 GND.n1617 0.306902
R15769 GND.n1274 GND.n1273 0.306902
R15770 GND.n8641 GND.n32 0.263073
R15771 GND.n8333 GND.n8332 0.256598
R15772 GND.n7597 GND.n668 0.256598
R15773 GND.n2868 GND.n2867 0.256598
R15774 GND.n6290 GND.n1624 0.256598
R15775 GND.n8332 GND.n444 0.241354
R15776 GND.n2867 GND.n2866 0.241354
R15777 GND.n7561 GND.n834 0.229039
R15778 GND.n7562 GND.n7561 0.229039
R15779 GND.n6246 GND.n1727 0.229039
R15780 GND.n1817 GND.n1727 0.229039
R15781 GND.n2782 GND.n2763 0.152939
R15782 GND.n2764 GND.n2763 0.152939
R15783 GND.n2765 GND.n2764 0.152939
R15784 GND.n2766 GND.n2765 0.152939
R15785 GND.n2767 GND.n2766 0.152939
R15786 GND.n2768 GND.n2767 0.152939
R15787 GND.n2769 GND.n2768 0.152939
R15788 GND.n2769 GND.n2048 0.152939
R15789 GND.n5120 GND.n2048 0.152939
R15790 GND.n5121 GND.n5120 0.152939
R15791 GND.n5122 GND.n5121 0.152939
R15792 GND.n5123 GND.n5122 0.152939
R15793 GND.n5124 GND.n5123 0.152939
R15794 GND.n5125 GND.n5124 0.152939
R15795 GND.n5126 GND.n5125 0.152939
R15796 GND.n5127 GND.n5126 0.152939
R15797 GND.n5128 GND.n5127 0.152939
R15798 GND.n5129 GND.n5128 0.152939
R15799 GND.n5130 GND.n5129 0.152939
R15800 GND.n5131 GND.n5130 0.152939
R15801 GND.n5132 GND.n5131 0.152939
R15802 GND.n5133 GND.n5132 0.152939
R15803 GND.n5134 GND.n5133 0.152939
R15804 GND.n5135 GND.n5134 0.152939
R15805 GND.n5136 GND.n5135 0.152939
R15806 GND.n5137 GND.n5136 0.152939
R15807 GND.n5138 GND.n5137 0.152939
R15808 GND.n5139 GND.n5138 0.152939
R15809 GND.n5140 GND.n5139 0.152939
R15810 GND.n5141 GND.n5140 0.152939
R15811 GND.n5142 GND.n5141 0.152939
R15812 GND.n5143 GND.n5142 0.152939
R15813 GND.n5144 GND.n5143 0.152939
R15814 GND.n5145 GND.n5144 0.152939
R15815 GND.n5146 GND.n5145 0.152939
R15816 GND.n5147 GND.n5146 0.152939
R15817 GND.n5147 GND.n1901 0.152939
R15818 GND.n5336 GND.n1901 0.152939
R15819 GND.n5337 GND.n5336 0.152939
R15820 GND.n5338 GND.n5337 0.152939
R15821 GND.n5339 GND.n5338 0.152939
R15822 GND.n5340 GND.n5339 0.152939
R15823 GND.n5341 GND.n5340 0.152939
R15824 GND.n5342 GND.n5341 0.152939
R15825 GND.n5343 GND.n5342 0.152939
R15826 GND.n5344 GND.n5343 0.152939
R15827 GND.n5344 GND.n1617 0.152939
R15828 GND.n4726 GND.n3023 0.152939
R15829 GND.n3029 GND.n3023 0.152939
R15830 GND.n3030 GND.n3029 0.152939
R15831 GND.n3031 GND.n3030 0.152939
R15832 GND.n3032 GND.n3031 0.152939
R15833 GND.n3037 GND.n3032 0.152939
R15834 GND.n3038 GND.n3037 0.152939
R15835 GND.n3039 GND.n3038 0.152939
R15836 GND.n3040 GND.n3039 0.152939
R15837 GND.n3045 GND.n3040 0.152939
R15838 GND.n3046 GND.n3045 0.152939
R15839 GND.n3047 GND.n3046 0.152939
R15840 GND.n3048 GND.n3047 0.152939
R15841 GND.n3053 GND.n3048 0.152939
R15842 GND.n3054 GND.n3053 0.152939
R15843 GND.n3055 GND.n3054 0.152939
R15844 GND.n3056 GND.n3055 0.152939
R15845 GND.n3061 GND.n3056 0.152939
R15846 GND.n3062 GND.n3061 0.152939
R15847 GND.n3063 GND.n3062 0.152939
R15848 GND.n3064 GND.n3063 0.152939
R15849 GND.n3069 GND.n3064 0.152939
R15850 GND.n3070 GND.n3069 0.152939
R15851 GND.n3071 GND.n3070 0.152939
R15852 GND.n3072 GND.n3071 0.152939
R15853 GND.n3077 GND.n3072 0.152939
R15854 GND.n3078 GND.n3077 0.152939
R15855 GND.n3079 GND.n3078 0.152939
R15856 GND.n3080 GND.n3079 0.152939
R15857 GND.n3085 GND.n3080 0.152939
R15858 GND.n3086 GND.n3085 0.152939
R15859 GND.n3087 GND.n3086 0.152939
R15860 GND.n3088 GND.n3087 0.152939
R15861 GND.n3093 GND.n3088 0.152939
R15862 GND.n3094 GND.n3093 0.152939
R15863 GND.n3095 GND.n3094 0.152939
R15864 GND.n3096 GND.n3095 0.152939
R15865 GND.n3101 GND.n3096 0.152939
R15866 GND.n3102 GND.n3101 0.152939
R15867 GND.n3103 GND.n3102 0.152939
R15868 GND.n3104 GND.n3103 0.152939
R15869 GND.n3109 GND.n3104 0.152939
R15870 GND.n3110 GND.n3109 0.152939
R15871 GND.n3111 GND.n3110 0.152939
R15872 GND.n3112 GND.n3111 0.152939
R15873 GND.n3117 GND.n3112 0.152939
R15874 GND.n3118 GND.n3117 0.152939
R15875 GND.n3119 GND.n3118 0.152939
R15876 GND.n3120 GND.n3119 0.152939
R15877 GND.n3125 GND.n3120 0.152939
R15878 GND.n3126 GND.n3125 0.152939
R15879 GND.n3127 GND.n3126 0.152939
R15880 GND.n3128 GND.n3127 0.152939
R15881 GND.n3133 GND.n3128 0.152939
R15882 GND.n3134 GND.n3133 0.152939
R15883 GND.n3135 GND.n3134 0.152939
R15884 GND.n3136 GND.n3135 0.152939
R15885 GND.n3141 GND.n3136 0.152939
R15886 GND.n3142 GND.n3141 0.152939
R15887 GND.n3143 GND.n3142 0.152939
R15888 GND.n3144 GND.n3143 0.152939
R15889 GND.n3149 GND.n3144 0.152939
R15890 GND.n3150 GND.n3149 0.152939
R15891 GND.n3151 GND.n3150 0.152939
R15892 GND.n3152 GND.n3151 0.152939
R15893 GND.n3157 GND.n3152 0.152939
R15894 GND.n3158 GND.n3157 0.152939
R15895 GND.n3159 GND.n3158 0.152939
R15896 GND.n3160 GND.n3159 0.152939
R15897 GND.n3165 GND.n3160 0.152939
R15898 GND.n3166 GND.n3165 0.152939
R15899 GND.n3167 GND.n3166 0.152939
R15900 GND.n3168 GND.n3167 0.152939
R15901 GND.n3173 GND.n3168 0.152939
R15902 GND.n3174 GND.n3173 0.152939
R15903 GND.n3175 GND.n3174 0.152939
R15904 GND.n3176 GND.n3175 0.152939
R15905 GND.n3181 GND.n3176 0.152939
R15906 GND.n3182 GND.n3181 0.152939
R15907 GND.n3183 GND.n3182 0.152939
R15908 GND.n3184 GND.n3183 0.152939
R15909 GND.n3189 GND.n3184 0.152939
R15910 GND.n3190 GND.n3189 0.152939
R15911 GND.n3191 GND.n3190 0.152939
R15912 GND.n3192 GND.n3191 0.152939
R15913 GND.n3197 GND.n3192 0.152939
R15914 GND.n3198 GND.n3197 0.152939
R15915 GND.n3199 GND.n3198 0.152939
R15916 GND.n3200 GND.n3199 0.152939
R15917 GND.n3205 GND.n3200 0.152939
R15918 GND.n3206 GND.n3205 0.152939
R15919 GND.n3207 GND.n3206 0.152939
R15920 GND.n3208 GND.n3207 0.152939
R15921 GND.n3213 GND.n3208 0.152939
R15922 GND.n3214 GND.n3213 0.152939
R15923 GND.n3215 GND.n3214 0.152939
R15924 GND.n3216 GND.n3215 0.152939
R15925 GND.n3221 GND.n3216 0.152939
R15926 GND.n3222 GND.n3221 0.152939
R15927 GND.n3223 GND.n3222 0.152939
R15928 GND.n3224 GND.n3223 0.152939
R15929 GND.n3229 GND.n3224 0.152939
R15930 GND.n3230 GND.n3229 0.152939
R15931 GND.n3231 GND.n3230 0.152939
R15932 GND.n3232 GND.n3231 0.152939
R15933 GND.n3237 GND.n3232 0.152939
R15934 GND.n3238 GND.n3237 0.152939
R15935 GND.n3239 GND.n3238 0.152939
R15936 GND.n3240 GND.n3239 0.152939
R15937 GND.n3245 GND.n3240 0.152939
R15938 GND.n3246 GND.n3245 0.152939
R15939 GND.n3247 GND.n3246 0.152939
R15940 GND.n3248 GND.n3247 0.152939
R15941 GND.n3253 GND.n3248 0.152939
R15942 GND.n3254 GND.n3253 0.152939
R15943 GND.n3255 GND.n3254 0.152939
R15944 GND.n3256 GND.n3255 0.152939
R15945 GND.n3261 GND.n3256 0.152939
R15946 GND.n3262 GND.n3261 0.152939
R15947 GND.n3263 GND.n3262 0.152939
R15948 GND.n3264 GND.n3263 0.152939
R15949 GND.n3269 GND.n3264 0.152939
R15950 GND.n3270 GND.n3269 0.152939
R15951 GND.n3271 GND.n3270 0.152939
R15952 GND.n3272 GND.n3271 0.152939
R15953 GND.n3277 GND.n3272 0.152939
R15954 GND.n3278 GND.n3277 0.152939
R15955 GND.n3279 GND.n3278 0.152939
R15956 GND.n3280 GND.n3279 0.152939
R15957 GND.n3285 GND.n3280 0.152939
R15958 GND.n3286 GND.n3285 0.152939
R15959 GND.n3287 GND.n3286 0.152939
R15960 GND.n3288 GND.n3287 0.152939
R15961 GND.n3293 GND.n3288 0.152939
R15962 GND.n3294 GND.n3293 0.152939
R15963 GND.n3295 GND.n3294 0.152939
R15964 GND.n3296 GND.n3295 0.152939
R15965 GND.n3301 GND.n3296 0.152939
R15966 GND.n3302 GND.n3301 0.152939
R15967 GND.n3303 GND.n3302 0.152939
R15968 GND.n3304 GND.n3303 0.152939
R15969 GND.n3309 GND.n3304 0.152939
R15970 GND.n3310 GND.n3309 0.152939
R15971 GND.n3311 GND.n3310 0.152939
R15972 GND.n3312 GND.n3311 0.152939
R15973 GND.n3317 GND.n3312 0.152939
R15974 GND.n3318 GND.n3317 0.152939
R15975 GND.n3319 GND.n3318 0.152939
R15976 GND.n3320 GND.n3319 0.152939
R15977 GND.n3325 GND.n3320 0.152939
R15978 GND.n3326 GND.n3325 0.152939
R15979 GND.n3327 GND.n3326 0.152939
R15980 GND.n3328 GND.n3327 0.152939
R15981 GND.n3333 GND.n3328 0.152939
R15982 GND.n3334 GND.n3333 0.152939
R15983 GND.n3335 GND.n3334 0.152939
R15984 GND.n3336 GND.n3335 0.152939
R15985 GND.n3341 GND.n3336 0.152939
R15986 GND.n3342 GND.n3341 0.152939
R15987 GND.n3343 GND.n3342 0.152939
R15988 GND.n3344 GND.n3343 0.152939
R15989 GND.n3349 GND.n3344 0.152939
R15990 GND.n3350 GND.n3349 0.152939
R15991 GND.n3351 GND.n3350 0.152939
R15992 GND.n3352 GND.n3351 0.152939
R15993 GND.n3357 GND.n3352 0.152939
R15994 GND.n3358 GND.n3357 0.152939
R15995 GND.n3359 GND.n3358 0.152939
R15996 GND.n3360 GND.n3359 0.152939
R15997 GND.n3365 GND.n3360 0.152939
R15998 GND.n3366 GND.n3365 0.152939
R15999 GND.n3367 GND.n3366 0.152939
R16000 GND.n3368 GND.n3367 0.152939
R16001 GND.n3373 GND.n3368 0.152939
R16002 GND.n3374 GND.n3373 0.152939
R16003 GND.n3375 GND.n3374 0.152939
R16004 GND.n3376 GND.n3375 0.152939
R16005 GND.n3381 GND.n3376 0.152939
R16006 GND.n3382 GND.n3381 0.152939
R16007 GND.n3383 GND.n3382 0.152939
R16008 GND.n3384 GND.n3383 0.152939
R16009 GND.n3389 GND.n3384 0.152939
R16010 GND.n3390 GND.n3389 0.152939
R16011 GND.n3391 GND.n3390 0.152939
R16012 GND.n3392 GND.n3391 0.152939
R16013 GND.n3397 GND.n3392 0.152939
R16014 GND.n3398 GND.n3397 0.152939
R16015 GND.n3399 GND.n3398 0.152939
R16016 GND.n3400 GND.n3399 0.152939
R16017 GND.n3405 GND.n3400 0.152939
R16018 GND.n3406 GND.n3405 0.152939
R16019 GND.n3407 GND.n3406 0.152939
R16020 GND.n3408 GND.n3407 0.152939
R16021 GND.n3413 GND.n3408 0.152939
R16022 GND.n3414 GND.n3413 0.152939
R16023 GND.n3415 GND.n3414 0.152939
R16024 GND.n3416 GND.n3415 0.152939
R16025 GND.n3421 GND.n3416 0.152939
R16026 GND.n3422 GND.n3421 0.152939
R16027 GND.n3423 GND.n3422 0.152939
R16028 GND.n3424 GND.n3423 0.152939
R16029 GND.n3429 GND.n3424 0.152939
R16030 GND.n3430 GND.n3429 0.152939
R16031 GND.n3431 GND.n3430 0.152939
R16032 GND.n3432 GND.n3431 0.152939
R16033 GND.n3437 GND.n3432 0.152939
R16034 GND.n3438 GND.n3437 0.152939
R16035 GND.n3439 GND.n3438 0.152939
R16036 GND.n3440 GND.n3439 0.152939
R16037 GND.n3445 GND.n3440 0.152939
R16038 GND.n3446 GND.n3445 0.152939
R16039 GND.n3447 GND.n3446 0.152939
R16040 GND.n3448 GND.n3447 0.152939
R16041 GND.n3453 GND.n3448 0.152939
R16042 GND.n3454 GND.n3453 0.152939
R16043 GND.n3455 GND.n3454 0.152939
R16044 GND.n3456 GND.n3455 0.152939
R16045 GND.n3461 GND.n3456 0.152939
R16046 GND.n3462 GND.n3461 0.152939
R16047 GND.n3463 GND.n3462 0.152939
R16048 GND.n3464 GND.n3463 0.152939
R16049 GND.n3469 GND.n3464 0.152939
R16050 GND.n3470 GND.n3469 0.152939
R16051 GND.n3471 GND.n3470 0.152939
R16052 GND.n3472 GND.n3471 0.152939
R16053 GND.n3477 GND.n3472 0.152939
R16054 GND.n3478 GND.n3477 0.152939
R16055 GND.n3479 GND.n3478 0.152939
R16056 GND.n3480 GND.n3479 0.152939
R16057 GND.n3485 GND.n3480 0.152939
R16058 GND.n3486 GND.n3485 0.152939
R16059 GND.n3487 GND.n3486 0.152939
R16060 GND.n3488 GND.n3487 0.152939
R16061 GND.n3493 GND.n3488 0.152939
R16062 GND.n3494 GND.n3493 0.152939
R16063 GND.n3495 GND.n3494 0.152939
R16064 GND.n3496 GND.n3495 0.152939
R16065 GND.n3501 GND.n3496 0.152939
R16066 GND.n3502 GND.n3501 0.152939
R16067 GND.n3503 GND.n3502 0.152939
R16068 GND.n3504 GND.n3503 0.152939
R16069 GND.n3509 GND.n3504 0.152939
R16070 GND.n3510 GND.n3509 0.152939
R16071 GND.n3511 GND.n3510 0.152939
R16072 GND.n3512 GND.n3511 0.152939
R16073 GND.n3517 GND.n3512 0.152939
R16074 GND.n3518 GND.n3517 0.152939
R16075 GND.n3519 GND.n3518 0.152939
R16076 GND.n3520 GND.n3519 0.152939
R16077 GND.n3525 GND.n3520 0.152939
R16078 GND.n3526 GND.n3525 0.152939
R16079 GND.n3527 GND.n3526 0.152939
R16080 GND.n3528 GND.n3527 0.152939
R16081 GND.n3533 GND.n3528 0.152939
R16082 GND.n3534 GND.n3533 0.152939
R16083 GND.n3535 GND.n3534 0.152939
R16084 GND.n3536 GND.n3535 0.152939
R16085 GND.n3541 GND.n3536 0.152939
R16086 GND.n3542 GND.n3541 0.152939
R16087 GND.n3543 GND.n3542 0.152939
R16088 GND.n3544 GND.n3543 0.152939
R16089 GND.n3549 GND.n3544 0.152939
R16090 GND.n3550 GND.n3549 0.152939
R16091 GND.n3551 GND.n3550 0.152939
R16092 GND.n3552 GND.n3551 0.152939
R16093 GND.n3557 GND.n3552 0.152939
R16094 GND.n3558 GND.n3557 0.152939
R16095 GND.n3559 GND.n3558 0.152939
R16096 GND.n3560 GND.n3559 0.152939
R16097 GND.n3565 GND.n3560 0.152939
R16098 GND.n3566 GND.n3565 0.152939
R16099 GND.n3567 GND.n3566 0.152939
R16100 GND.n3568 GND.n3567 0.152939
R16101 GND.n3573 GND.n3568 0.152939
R16102 GND.n3574 GND.n3573 0.152939
R16103 GND.n3575 GND.n3574 0.152939
R16104 GND.n3576 GND.n3575 0.152939
R16105 GND.n3581 GND.n3576 0.152939
R16106 GND.n3582 GND.n3581 0.152939
R16107 GND.n3583 GND.n3582 0.152939
R16108 GND.n3584 GND.n3583 0.152939
R16109 GND.n3589 GND.n3584 0.152939
R16110 GND.n3590 GND.n3589 0.152939
R16111 GND.n3591 GND.n3590 0.152939
R16112 GND.n3592 GND.n3591 0.152939
R16113 GND.n3597 GND.n3592 0.152939
R16114 GND.n3598 GND.n3597 0.152939
R16115 GND.n3599 GND.n3598 0.152939
R16116 GND.n3600 GND.n3599 0.152939
R16117 GND.n3605 GND.n3600 0.152939
R16118 GND.n3606 GND.n3605 0.152939
R16119 GND.n3607 GND.n3606 0.152939
R16120 GND.n3608 GND.n3607 0.152939
R16121 GND.n3613 GND.n3608 0.152939
R16122 GND.n3614 GND.n3613 0.152939
R16123 GND.n3615 GND.n3614 0.152939
R16124 GND.n3616 GND.n3615 0.152939
R16125 GND.n3621 GND.n3616 0.152939
R16126 GND.n3622 GND.n3621 0.152939
R16127 GND.n3623 GND.n3622 0.152939
R16128 GND.n3624 GND.n3623 0.152939
R16129 GND.n3629 GND.n3624 0.152939
R16130 GND.n3630 GND.n3629 0.152939
R16131 GND.n3631 GND.n3630 0.152939
R16132 GND.n3632 GND.n3631 0.152939
R16133 GND.n3637 GND.n3632 0.152939
R16134 GND.n3638 GND.n3637 0.152939
R16135 GND.n3639 GND.n3638 0.152939
R16136 GND.n3640 GND.n3639 0.152939
R16137 GND.n3645 GND.n3640 0.152939
R16138 GND.n3646 GND.n3645 0.152939
R16139 GND.n3647 GND.n3646 0.152939
R16140 GND.n3648 GND.n3647 0.152939
R16141 GND.n3653 GND.n3648 0.152939
R16142 GND.n3654 GND.n3653 0.152939
R16143 GND.n3655 GND.n3654 0.152939
R16144 GND.n3656 GND.n3655 0.152939
R16145 GND.n3661 GND.n3656 0.152939
R16146 GND.n3662 GND.n3661 0.152939
R16147 GND.n3663 GND.n3662 0.152939
R16148 GND.n3664 GND.n3663 0.152939
R16149 GND.n3669 GND.n3664 0.152939
R16150 GND.n3670 GND.n3669 0.152939
R16151 GND.n3671 GND.n3670 0.152939
R16152 GND.n3672 GND.n3671 0.152939
R16153 GND.n3677 GND.n3672 0.152939
R16154 GND.n3678 GND.n3677 0.152939
R16155 GND.n3679 GND.n3678 0.152939
R16156 GND.n3680 GND.n3679 0.152939
R16157 GND.n3685 GND.n3680 0.152939
R16158 GND.n3686 GND.n3685 0.152939
R16159 GND.n3687 GND.n3686 0.152939
R16160 GND.n3688 GND.n3687 0.152939
R16161 GND.n3693 GND.n3688 0.152939
R16162 GND.n3694 GND.n3693 0.152939
R16163 GND.n3695 GND.n3694 0.152939
R16164 GND.n3696 GND.n3695 0.152939
R16165 GND.n3701 GND.n3696 0.152939
R16166 GND.n3702 GND.n3701 0.152939
R16167 GND.n3703 GND.n3702 0.152939
R16168 GND.n3704 GND.n3703 0.152939
R16169 GND.n3709 GND.n3704 0.152939
R16170 GND.n3710 GND.n3709 0.152939
R16171 GND.n3711 GND.n3710 0.152939
R16172 GND.n3712 GND.n3711 0.152939
R16173 GND.n3717 GND.n3712 0.152939
R16174 GND.n3718 GND.n3717 0.152939
R16175 GND.n3719 GND.n3718 0.152939
R16176 GND.n3720 GND.n3719 0.152939
R16177 GND.n3725 GND.n3720 0.152939
R16178 GND.n3726 GND.n3725 0.152939
R16179 GND.n3727 GND.n3726 0.152939
R16180 GND.n3728 GND.n3727 0.152939
R16181 GND.n3733 GND.n3728 0.152939
R16182 GND.n3734 GND.n3733 0.152939
R16183 GND.n3735 GND.n3734 0.152939
R16184 GND.n3736 GND.n3735 0.152939
R16185 GND.n3741 GND.n3736 0.152939
R16186 GND.n3742 GND.n3741 0.152939
R16187 GND.n3743 GND.n3742 0.152939
R16188 GND.n3744 GND.n3743 0.152939
R16189 GND.n3749 GND.n3744 0.152939
R16190 GND.n3750 GND.n3749 0.152939
R16191 GND.n3751 GND.n3750 0.152939
R16192 GND.n3752 GND.n3751 0.152939
R16193 GND.n3757 GND.n3752 0.152939
R16194 GND.n3758 GND.n3757 0.152939
R16195 GND.n3759 GND.n3758 0.152939
R16196 GND.n3760 GND.n3759 0.152939
R16197 GND.n3765 GND.n3760 0.152939
R16198 GND.n3766 GND.n3765 0.152939
R16199 GND.n3767 GND.n3766 0.152939
R16200 GND.n3768 GND.n3767 0.152939
R16201 GND.n3773 GND.n3768 0.152939
R16202 GND.n3774 GND.n3773 0.152939
R16203 GND.n3775 GND.n3774 0.152939
R16204 GND.n3776 GND.n3775 0.152939
R16205 GND.n3781 GND.n3776 0.152939
R16206 GND.n3782 GND.n3781 0.152939
R16207 GND.n3964 GND.n3782 0.152939
R16208 GND.n3963 GND.n3783 0.152939
R16209 GND.n3788 GND.n3783 0.152939
R16210 GND.n3789 GND.n3788 0.152939
R16211 GND.n3790 GND.n3789 0.152939
R16212 GND.n3795 GND.n3790 0.152939
R16213 GND.n3796 GND.n3795 0.152939
R16214 GND.n3797 GND.n3796 0.152939
R16215 GND.n3798 GND.n3797 0.152939
R16216 GND.n3803 GND.n3798 0.152939
R16217 GND.n3804 GND.n3803 0.152939
R16218 GND.n3805 GND.n3804 0.152939
R16219 GND.n3806 GND.n3805 0.152939
R16220 GND.n3811 GND.n3806 0.152939
R16221 GND.n3812 GND.n3811 0.152939
R16222 GND.n3813 GND.n3812 0.152939
R16223 GND.n3814 GND.n3813 0.152939
R16224 GND.n3819 GND.n3814 0.152939
R16225 GND.n3820 GND.n3819 0.152939
R16226 GND.n3821 GND.n3820 0.152939
R16227 GND.n3822 GND.n3821 0.152939
R16228 GND.n3827 GND.n3822 0.152939
R16229 GND.n3828 GND.n3827 0.152939
R16230 GND.n3829 GND.n3828 0.152939
R16231 GND.n3830 GND.n3829 0.152939
R16232 GND.n3835 GND.n3830 0.152939
R16233 GND.n3836 GND.n3835 0.152939
R16234 GND.n3837 GND.n3836 0.152939
R16235 GND.n3838 GND.n3837 0.152939
R16236 GND.n3843 GND.n3838 0.152939
R16237 GND.n3844 GND.n3843 0.152939
R16238 GND.n3845 GND.n3844 0.152939
R16239 GND.n3846 GND.n3845 0.152939
R16240 GND.n3851 GND.n3846 0.152939
R16241 GND.n3852 GND.n3851 0.152939
R16242 GND.n3853 GND.n3852 0.152939
R16243 GND.n3854 GND.n3853 0.152939
R16244 GND.n3859 GND.n3854 0.152939
R16245 GND.n3860 GND.n3859 0.152939
R16246 GND.n3861 GND.n3860 0.152939
R16247 GND.n3862 GND.n3861 0.152939
R16248 GND.n3867 GND.n3862 0.152939
R16249 GND.n3868 GND.n3867 0.152939
R16250 GND.n3869 GND.n3868 0.152939
R16251 GND.n3871 GND.n3869 0.152939
R16252 GND.n3871 GND.n3870 0.152939
R16253 GND.n3870 GND.n346 0.152939
R16254 GND.n8454 GND.n346 0.152939
R16255 GND.n8633 GND.n77 0.152939
R16256 GND.n158 GND.n77 0.152939
R16257 GND.n159 GND.n158 0.152939
R16258 GND.n177 GND.n159 0.152939
R16259 GND.n178 GND.n177 0.152939
R16260 GND.n179 GND.n178 0.152939
R16261 GND.n180 GND.n179 0.152939
R16262 GND.n198 GND.n180 0.152939
R16263 GND.n199 GND.n198 0.152939
R16264 GND.n200 GND.n199 0.152939
R16265 GND.n201 GND.n200 0.152939
R16266 GND.n219 GND.n201 0.152939
R16267 GND.n220 GND.n219 0.152939
R16268 GND.n221 GND.n220 0.152939
R16269 GND.n222 GND.n221 0.152939
R16270 GND.n240 GND.n222 0.152939
R16271 GND.n241 GND.n240 0.152939
R16272 GND.n242 GND.n241 0.152939
R16273 GND.n243 GND.n242 0.152939
R16274 GND.n261 GND.n243 0.152939
R16275 GND.n262 GND.n261 0.152939
R16276 GND.n263 GND.n262 0.152939
R16277 GND.n264 GND.n263 0.152939
R16278 GND.n282 GND.n264 0.152939
R16279 GND.n283 GND.n282 0.152939
R16280 GND.n284 GND.n283 0.152939
R16281 GND.n285 GND.n284 0.152939
R16282 GND.n303 GND.n285 0.152939
R16283 GND.n304 GND.n303 0.152939
R16284 GND.n305 GND.n304 0.152939
R16285 GND.n306 GND.n305 0.152939
R16286 GND.n324 GND.n306 0.152939
R16287 GND.n325 GND.n324 0.152939
R16288 GND.n326 GND.n325 0.152939
R16289 GND.n327 GND.n326 0.152939
R16290 GND.n345 GND.n327 0.152939
R16291 GND.n8455 GND.n345 0.152939
R16292 GND.n7992 GND.n82 0.152939
R16293 GND.n7993 GND.n7992 0.152939
R16294 GND.n7993 GND.n474 0.152939
R16295 GND.n7999 GND.n474 0.152939
R16296 GND.n8000 GND.n7999 0.152939
R16297 GND.n8001 GND.n8000 0.152939
R16298 GND.n8001 GND.n472 0.152939
R16299 GND.n8007 GND.n472 0.152939
R16300 GND.n8008 GND.n8007 0.152939
R16301 GND.n8009 GND.n8008 0.152939
R16302 GND.n8009 GND.n470 0.152939
R16303 GND.n8015 GND.n470 0.152939
R16304 GND.n8016 GND.n8015 0.152939
R16305 GND.n8017 GND.n8016 0.152939
R16306 GND.n8017 GND.n468 0.152939
R16307 GND.n8023 GND.n468 0.152939
R16308 GND.n8024 GND.n8023 0.152939
R16309 GND.n8025 GND.n8024 0.152939
R16310 GND.n8025 GND.n466 0.152939
R16311 GND.n8031 GND.n466 0.152939
R16312 GND.n8032 GND.n8031 0.152939
R16313 GND.n8033 GND.n8032 0.152939
R16314 GND.n8033 GND.n464 0.152939
R16315 GND.n8039 GND.n464 0.152939
R16316 GND.n8040 GND.n8039 0.152939
R16317 GND.n8041 GND.n8040 0.152939
R16318 GND.n8041 GND.n462 0.152939
R16319 GND.n8047 GND.n462 0.152939
R16320 GND.n8048 GND.n8047 0.152939
R16321 GND.n8049 GND.n8048 0.152939
R16322 GND.n8049 GND.n460 0.152939
R16323 GND.n8055 GND.n460 0.152939
R16324 GND.n8056 GND.n8055 0.152939
R16325 GND.n8057 GND.n8056 0.152939
R16326 GND.n8057 GND.n458 0.152939
R16327 GND.n8063 GND.n458 0.152939
R16328 GND.n8064 GND.n8063 0.152939
R16329 GND.n8065 GND.n8064 0.152939
R16330 GND.n8065 GND.n455 0.152939
R16331 GND.n8319 GND.n455 0.152939
R16332 GND.n8320 GND.n8319 0.152939
R16333 GND.n8321 GND.n8320 0.152939
R16334 GND.n8322 GND.n8321 0.152939
R16335 GND.n6980 GND.n1180 0.152939
R16336 GND.n1184 GND.n1180 0.152939
R16337 GND.n1185 GND.n1184 0.152939
R16338 GND.n1186 GND.n1185 0.152939
R16339 GND.n1187 GND.n1186 0.152939
R16340 GND.n1188 GND.n1187 0.152939
R16341 GND.n1192 GND.n1188 0.152939
R16342 GND.n1193 GND.n1192 0.152939
R16343 GND.n1194 GND.n1193 0.152939
R16344 GND.n1195 GND.n1194 0.152939
R16345 GND.n6312 GND.n1568 0.152939
R16346 GND.n6452 GND.n1568 0.152939
R16347 GND.n6453 GND.n6452 0.152939
R16348 GND.n6454 GND.n6453 0.152939
R16349 GND.n6454 GND.n1541 0.152939
R16350 GND.n6485 GND.n1541 0.152939
R16351 GND.n6486 GND.n6485 0.152939
R16352 GND.n6487 GND.n6486 0.152939
R16353 GND.n6488 GND.n6487 0.152939
R16354 GND.n6489 GND.n6488 0.152939
R16355 GND.n6489 GND.n1505 0.152939
R16356 GND.n6548 GND.n1505 0.152939
R16357 GND.n6549 GND.n6548 0.152939
R16358 GND.n6550 GND.n6549 0.152939
R16359 GND.n6550 GND.n1479 0.152939
R16360 GND.n6600 GND.n1479 0.152939
R16361 GND.n6601 GND.n6600 0.152939
R16362 GND.n6602 GND.n6601 0.152939
R16363 GND.n6602 GND.n1439 0.152939
R16364 GND.n6638 GND.n1439 0.152939
R16365 GND.n6639 GND.n6638 0.152939
R16366 GND.n6640 GND.n6639 0.152939
R16367 GND.n6641 GND.n6640 0.152939
R16368 GND.n6641 GND.n1408 0.152939
R16369 GND.n6697 GND.n1408 0.152939
R16370 GND.n6698 GND.n6697 0.152939
R16371 GND.n6699 GND.n6698 0.152939
R16372 GND.n6700 GND.n6699 0.152939
R16373 GND.n6700 GND.n1377 0.152939
R16374 GND.n6765 GND.n1377 0.152939
R16375 GND.n6766 GND.n6765 0.152939
R16376 GND.n6767 GND.n6766 0.152939
R16377 GND.n6768 GND.n6767 0.152939
R16378 GND.n6768 GND.n1346 0.152939
R16379 GND.n6832 GND.n1346 0.152939
R16380 GND.n6833 GND.n6832 0.152939
R16381 GND.n6834 GND.n6833 0.152939
R16382 GND.n6836 GND.n6834 0.152939
R16383 GND.n6836 GND.n6835 0.152939
R16384 GND.n6835 GND.n1325 0.152939
R16385 GND.n6862 GND.n1325 0.152939
R16386 GND.n6863 GND.n6862 0.152939
R16387 GND.n6864 GND.n6863 0.152939
R16388 GND.n6865 GND.n6864 0.152939
R16389 GND.n6866 GND.n6865 0.152939
R16390 GND.n6866 GND.n1179 0.152939
R16391 GND.n6981 GND.n1179 0.152939
R16392 GND.n6319 GND.n6310 0.152939
R16393 GND.n6320 GND.n6319 0.152939
R16394 GND.n6321 GND.n6320 0.152939
R16395 GND.n6321 GND.n6306 0.152939
R16396 GND.n6329 GND.n6306 0.152939
R16397 GND.n6330 GND.n6329 0.152939
R16398 GND.n6332 GND.n6330 0.152939
R16399 GND.n6332 GND.n6331 0.152939
R16400 GND.n6331 GND.n6303 0.152939
R16401 GND.n6303 GND.n1616 0.152939
R16402 GND.n6371 GND.n6370 0.152939
R16403 GND.n6379 GND.n1611 0.152939
R16404 GND.n6380 GND.n6379 0.152939
R16405 GND.n6381 GND.n6380 0.152939
R16406 GND.n6382 GND.n6381 0.152939
R16407 GND.n6383 GND.n6382 0.152939
R16408 GND.n6384 GND.n6383 0.152939
R16409 GND.n6385 GND.n6384 0.152939
R16410 GND.n6386 GND.n6385 0.152939
R16411 GND.n6387 GND.n6386 0.152939
R16412 GND.n6389 GND.n6387 0.152939
R16413 GND.n6390 GND.n6389 0.152939
R16414 GND.n6392 GND.n6390 0.152939
R16415 GND.n6392 GND.n6391 0.152939
R16416 GND.n6391 GND.n1499 0.152939
R16417 GND.n6557 GND.n1499 0.152939
R16418 GND.n6558 GND.n6557 0.152939
R16419 GND.n6559 GND.n6558 0.152939
R16420 GND.n6560 GND.n6559 0.152939
R16421 GND.n6561 GND.n6560 0.152939
R16422 GND.n6562 GND.n6561 0.152939
R16423 GND.n6565 GND.n6562 0.152939
R16424 GND.n6565 GND.n6564 0.152939
R16425 GND.n6564 GND.n6563 0.152939
R16426 GND.n6563 GND.n1430 0.152939
R16427 GND.n6651 GND.n1430 0.152939
R16428 GND.n6652 GND.n6651 0.152939
R16429 GND.n6653 GND.n6652 0.152939
R16430 GND.n6653 GND.n1427 0.152939
R16431 GND.n6658 GND.n1427 0.152939
R16432 GND.n6659 GND.n6658 0.152939
R16433 GND.n6660 GND.n6659 0.152939
R16434 GND.n6661 GND.n6660 0.152939
R16435 GND.n6661 GND.n1357 0.152939
R16436 GND.n6793 GND.n1357 0.152939
R16437 GND.n6794 GND.n6793 0.152939
R16438 GND.n6795 GND.n6794 0.152939
R16439 GND.n6796 GND.n6795 0.152939
R16440 GND.n6797 GND.n6796 0.152939
R16441 GND.n6798 GND.n6797 0.152939
R16442 GND.n6799 GND.n6798 0.152939
R16443 GND.n6801 GND.n6799 0.152939
R16444 GND.n6802 GND.n6801 0.152939
R16445 GND.n6803 GND.n6802 0.152939
R16446 GND.n6805 GND.n6803 0.152939
R16447 GND.n6805 GND.n6804 0.152939
R16448 GND.n6804 GND.n1287 0.152939
R16449 GND.n6929 GND.n1287 0.152939
R16450 GND.n6930 GND.n1286 0.152939
R16451 GND.n1273 GND.n1227 0.152939
R16452 GND.n1229 GND.n1227 0.152939
R16453 GND.n1230 GND.n1229 0.152939
R16454 GND.n1231 GND.n1230 0.152939
R16455 GND.n1232 GND.n1231 0.152939
R16456 GND.n1233 GND.n1232 0.152939
R16457 GND.n1234 GND.n1233 0.152939
R16458 GND.n1235 GND.n1234 0.152939
R16459 GND.n1236 GND.n1235 0.152939
R16460 GND.n1237 GND.n1236 0.152939
R16461 GND.n1238 GND.n1237 0.152939
R16462 GND.n1239 GND.n1238 0.152939
R16463 GND.n1240 GND.n1239 0.152939
R16464 GND.n1241 GND.n1240 0.152939
R16465 GND.n1242 GND.n1241 0.152939
R16466 GND.n1243 GND.n1242 0.152939
R16467 GND.n1244 GND.n1243 0.152939
R16468 GND.n1245 GND.n1244 0.152939
R16469 GND.n1245 GND.n564 0.152939
R16470 GND.n7821 GND.n564 0.152939
R16471 GND.n7822 GND.n7821 0.152939
R16472 GND.n7823 GND.n7822 0.152939
R16473 GND.n7824 GND.n7823 0.152939
R16474 GND.n7825 GND.n7824 0.152939
R16475 GND.n7826 GND.n7825 0.152939
R16476 GND.n7827 GND.n7826 0.152939
R16477 GND.n7828 GND.n7827 0.152939
R16478 GND.n7829 GND.n7828 0.152939
R16479 GND.n7830 GND.n7829 0.152939
R16480 GND.n7831 GND.n7830 0.152939
R16481 GND.n7832 GND.n7831 0.152939
R16482 GND.n7833 GND.n7832 0.152939
R16483 GND.n7834 GND.n7833 0.152939
R16484 GND.n7835 GND.n7834 0.152939
R16485 GND.n7836 GND.n7835 0.152939
R16486 GND.n7837 GND.n7836 0.152939
R16487 GND.n7838 GND.n7837 0.152939
R16488 GND.n7839 GND.n7838 0.152939
R16489 GND.n7840 GND.n7839 0.152939
R16490 GND.n7842 GND.n7840 0.152939
R16491 GND.n7842 GND.n7841 0.152939
R16492 GND.n7841 GND.n107 0.152939
R16493 GND.n8613 GND.n107 0.152939
R16494 GND.n8614 GND.n8613 0.152939
R16495 GND.n8615 GND.n8614 0.152939
R16496 GND.n8616 GND.n8615 0.152939
R16497 GND.n8616 GND.n62 0.152939
R16498 GND.n8094 GND.n63 0.152939
R16499 GND.n8098 GND.n8094 0.152939
R16500 GND.n8099 GND.n8098 0.152939
R16501 GND.n8100 GND.n8099 0.152939
R16502 GND.n8100 GND.n8092 0.152939
R16503 GND.n8106 GND.n8092 0.152939
R16504 GND.n8107 GND.n8106 0.152939
R16505 GND.n8108 GND.n8107 0.152939
R16506 GND.n8108 GND.n8090 0.152939
R16507 GND.n8114 GND.n8090 0.152939
R16508 GND.n8115 GND.n8114 0.152939
R16509 GND.n8116 GND.n8115 0.152939
R16510 GND.n8116 GND.n8088 0.152939
R16511 GND.n8122 GND.n8088 0.152939
R16512 GND.n8123 GND.n8122 0.152939
R16513 GND.n8124 GND.n8123 0.152939
R16514 GND.n8124 GND.n8086 0.152939
R16515 GND.n8130 GND.n8086 0.152939
R16516 GND.n8131 GND.n8130 0.152939
R16517 GND.n8132 GND.n8131 0.152939
R16518 GND.n8132 GND.n8084 0.152939
R16519 GND.n8138 GND.n8084 0.152939
R16520 GND.n8139 GND.n8138 0.152939
R16521 GND.n8140 GND.n8139 0.152939
R16522 GND.n8140 GND.n8082 0.152939
R16523 GND.n8146 GND.n8082 0.152939
R16524 GND.n8147 GND.n8146 0.152939
R16525 GND.n8148 GND.n8147 0.152939
R16526 GND.n8148 GND.n8080 0.152939
R16527 GND.n8154 GND.n8080 0.152939
R16528 GND.n8155 GND.n8154 0.152939
R16529 GND.n8156 GND.n8155 0.152939
R16530 GND.n8156 GND.n8078 0.152939
R16531 GND.n8162 GND.n8078 0.152939
R16532 GND.n8163 GND.n8162 0.152939
R16533 GND.n8164 GND.n8163 0.152939
R16534 GND.n8164 GND.n8076 0.152939
R16535 GND.n8170 GND.n8076 0.152939
R16536 GND.n8171 GND.n8170 0.152939
R16537 GND.n8172 GND.n8171 0.152939
R16538 GND.n8172 GND.n8074 0.152939
R16539 GND.n8178 GND.n8074 0.152939
R16540 GND.n8179 GND.n8178 0.152939
R16541 GND.n8180 GND.n8179 0.152939
R16542 GND.n8181 GND.n8180 0.152939
R16543 GND.n8182 GND.n8181 0.152939
R16544 GND.n8183 GND.n8182 0.152939
R16545 GND.n8193 GND.n444 0.152939
R16546 GND.n8194 GND.n8193 0.152939
R16547 GND.n8194 GND.n8189 0.152939
R16548 GND.n8202 GND.n8189 0.152939
R16549 GND.n8203 GND.n8202 0.152939
R16550 GND.n8204 GND.n8203 0.152939
R16551 GND.n8204 GND.n8187 0.152939
R16552 GND.n8212 GND.n8187 0.152939
R16553 GND.n8213 GND.n8212 0.152939
R16554 GND.n8214 GND.n8213 0.152939
R16555 GND.n8444 GND.n386 0.152939
R16556 GND.n8444 GND.n8443 0.152939
R16557 GND.n8443 GND.n8442 0.152939
R16558 GND.n8442 GND.n388 0.152939
R16559 GND.n389 GND.n388 0.152939
R16560 GND.n390 GND.n389 0.152939
R16561 GND.n391 GND.n390 0.152939
R16562 GND.n392 GND.n391 0.152939
R16563 GND.n8426 GND.n392 0.152939
R16564 GND.n8426 GND.n8425 0.152939
R16565 GND.n8425 GND.n8424 0.152939
R16566 GND.n8424 GND.n396 0.152939
R16567 GND.n397 GND.n396 0.152939
R16568 GND.n398 GND.n397 0.152939
R16569 GND.n399 GND.n398 0.152939
R16570 GND.n400 GND.n399 0.152939
R16571 GND.n401 GND.n400 0.152939
R16572 GND.n402 GND.n401 0.152939
R16573 GND.n403 GND.n402 0.152939
R16574 GND.n8403 GND.n403 0.152939
R16575 GND.n8403 GND.n8402 0.152939
R16576 GND.n8402 GND.n8401 0.152939
R16577 GND.n8401 GND.n409 0.152939
R16578 GND.n410 GND.n409 0.152939
R16579 GND.n411 GND.n410 0.152939
R16580 GND.n412 GND.n411 0.152939
R16581 GND.n413 GND.n412 0.152939
R16582 GND.n414 GND.n413 0.152939
R16583 GND.n415 GND.n414 0.152939
R16584 GND.n416 GND.n415 0.152939
R16585 GND.n8380 GND.n416 0.152939
R16586 GND.n8380 GND.n8379 0.152939
R16587 GND.n8379 GND.n8378 0.152939
R16588 GND.n8378 GND.n420 0.152939
R16589 GND.n421 GND.n420 0.152939
R16590 GND.n422 GND.n421 0.152939
R16591 GND.n423 GND.n422 0.152939
R16592 GND.n424 GND.n423 0.152939
R16593 GND.n425 GND.n424 0.152939
R16594 GND.n426 GND.n425 0.152939
R16595 GND.n427 GND.n426 0.152939
R16596 GND.n8357 GND.n427 0.152939
R16597 GND.n8357 GND.n8356 0.152939
R16598 GND.n8356 GND.n8355 0.152939
R16599 GND.n8355 GND.n433 0.152939
R16600 GND.n434 GND.n433 0.152939
R16601 GND.n435 GND.n434 0.152939
R16602 GND.n436 GND.n435 0.152939
R16603 GND.n437 GND.n436 0.152939
R16604 GND.n438 GND.n437 0.152939
R16605 GND.n439 GND.n438 0.152939
R16606 GND.n440 GND.n439 0.152939
R16607 GND.n8334 GND.n440 0.152939
R16608 GND.n8334 GND.n8333 0.152939
R16609 GND.n807 GND.n806 0.152939
R16610 GND.n808 GND.n807 0.152939
R16611 GND.n809 GND.n808 0.152939
R16612 GND.n810 GND.n809 0.152939
R16613 GND.n811 GND.n810 0.152939
R16614 GND.n812 GND.n811 0.152939
R16615 GND.n813 GND.n812 0.152939
R16616 GND.n814 GND.n813 0.152939
R16617 GND.n815 GND.n814 0.152939
R16618 GND.n818 GND.n815 0.152939
R16619 GND.n819 GND.n818 0.152939
R16620 GND.n820 GND.n819 0.152939
R16621 GND.n821 GND.n820 0.152939
R16622 GND.n822 GND.n821 0.152939
R16623 GND.n823 GND.n822 0.152939
R16624 GND.n824 GND.n823 0.152939
R16625 GND.n825 GND.n824 0.152939
R16626 GND.n826 GND.n825 0.152939
R16627 GND.n827 GND.n826 0.152939
R16628 GND.n829 GND.n827 0.152939
R16629 GND.n832 GND.n829 0.152939
R16630 GND.n833 GND.n832 0.152939
R16631 GND.n834 GND.n833 0.152939
R16632 GND.n7563 GND.n7562 0.152939
R16633 GND.n7564 GND.n7563 0.152939
R16634 GND.n7565 GND.n7564 0.152939
R16635 GND.n7566 GND.n7565 0.152939
R16636 GND.n7567 GND.n7566 0.152939
R16637 GND.n7570 GND.n7567 0.152939
R16638 GND.n7571 GND.n7570 0.152939
R16639 GND.n7572 GND.n7571 0.152939
R16640 GND.n7573 GND.n7572 0.152939
R16641 GND.n7574 GND.n7573 0.152939
R16642 GND.n7575 GND.n7574 0.152939
R16643 GND.n7576 GND.n7575 0.152939
R16644 GND.n7577 GND.n7576 0.152939
R16645 GND.n7578 GND.n7577 0.152939
R16646 GND.n7579 GND.n7578 0.152939
R16647 GND.n7581 GND.n7579 0.152939
R16648 GND.n7584 GND.n7581 0.152939
R16649 GND.n7585 GND.n7584 0.152939
R16650 GND.n7586 GND.n7585 0.152939
R16651 GND.n7587 GND.n7586 0.152939
R16652 GND.n7588 GND.n7587 0.152939
R16653 GND.n7589 GND.n7588 0.152939
R16654 GND.n7590 GND.n7589 0.152939
R16655 GND.n7591 GND.n7590 0.152939
R16656 GND.n7592 GND.n7591 0.152939
R16657 GND.n7593 GND.n7592 0.152939
R16658 GND.n7598 GND.n7593 0.152939
R16659 GND.n7598 GND.n7597 0.152939
R16660 GND.n805 GND.n714 0.152939
R16661 GND.n715 GND.n714 0.152939
R16662 GND.n716 GND.n715 0.152939
R16663 GND.n717 GND.n716 0.152939
R16664 GND.n718 GND.n717 0.152939
R16665 GND.n719 GND.n718 0.152939
R16666 GND.n720 GND.n719 0.152939
R16667 GND.n721 GND.n720 0.152939
R16668 GND.n722 GND.n721 0.152939
R16669 GND.n723 GND.n722 0.152939
R16670 GND.n724 GND.n723 0.152939
R16671 GND.n725 GND.n724 0.152939
R16672 GND.n726 GND.n725 0.152939
R16673 GND.n727 GND.n726 0.152939
R16674 GND.n728 GND.n727 0.152939
R16675 GND.n729 GND.n728 0.152939
R16676 GND.n730 GND.n729 0.152939
R16677 GND.n731 GND.n730 0.152939
R16678 GND.n732 GND.n731 0.152939
R16679 GND.n733 GND.n732 0.152939
R16680 GND.n734 GND.n733 0.152939
R16681 GND.n735 GND.n734 0.152939
R16682 GND.n736 GND.n735 0.152939
R16683 GND.n737 GND.n736 0.152939
R16684 GND.n738 GND.n737 0.152939
R16685 GND.n739 GND.n738 0.152939
R16686 GND.n740 GND.n739 0.152939
R16687 GND.n741 GND.n740 0.152939
R16688 GND.n742 GND.n741 0.152939
R16689 GND.n743 GND.n742 0.152939
R16690 GND.n744 GND.n743 0.152939
R16691 GND.n745 GND.n744 0.152939
R16692 GND.n746 GND.n745 0.152939
R16693 GND.n747 GND.n746 0.152939
R16694 GND.n748 GND.n747 0.152939
R16695 GND.n750 GND.n748 0.152939
R16696 GND.n750 GND.n749 0.152939
R16697 GND.n749 GND.n478 0.152939
R16698 GND.n478 GND.n476 0.152939
R16699 GND.n7964 GND.n476 0.152939
R16700 GND.n7965 GND.n7964 0.152939
R16701 GND.n7966 GND.n7965 0.152939
R16702 GND.n7966 GND.n82 0.152939
R16703 GND.n5087 GND.n5086 0.152939
R16704 GND.n5087 GND.n2058 0.152939
R16705 GND.n5110 GND.n2058 0.152939
R16706 GND.n5111 GND.n5110 0.152939
R16707 GND.n5112 GND.n5111 0.152939
R16708 GND.n5113 GND.n5112 0.152939
R16709 GND.n5113 GND.n2031 0.152939
R16710 GND.n5201 GND.n2031 0.152939
R16711 GND.n5202 GND.n5201 0.152939
R16712 GND.n5203 GND.n5202 0.152939
R16713 GND.n5203 GND.n2011 0.152939
R16714 GND.n5221 GND.n2011 0.152939
R16715 GND.n5222 GND.n5221 0.152939
R16716 GND.n5223 GND.n5222 0.152939
R16717 GND.n5223 GND.n1991 0.152939
R16718 GND.n5241 GND.n1991 0.152939
R16719 GND.n5242 GND.n5241 0.152939
R16720 GND.n5243 GND.n5242 0.152939
R16721 GND.n5243 GND.n1971 0.152939
R16722 GND.n5261 GND.n1971 0.152939
R16723 GND.n5262 GND.n5261 0.152939
R16724 GND.n5263 GND.n5262 0.152939
R16725 GND.n5263 GND.n1951 0.152939
R16726 GND.n5281 GND.n1951 0.152939
R16727 GND.n5282 GND.n5281 0.152939
R16728 GND.n5283 GND.n5282 0.152939
R16729 GND.n5283 GND.n1931 0.152939
R16730 GND.n5301 GND.n1931 0.152939
R16731 GND.n5302 GND.n5301 0.152939
R16732 GND.n5303 GND.n5302 0.152939
R16733 GND.n5303 GND.n1911 0.152939
R16734 GND.n5326 GND.n1911 0.152939
R16735 GND.n5327 GND.n5326 0.152939
R16736 GND.n5328 GND.n5327 0.152939
R16737 GND.n5329 GND.n5328 0.152939
R16738 GND.n5329 GND.n1884 0.152939
R16739 GND.n5371 GND.n1884 0.152939
R16740 GND.n5372 GND.n5371 0.152939
R16741 GND.n5373 GND.n5372 0.152939
R16742 GND.n5374 GND.n5373 0.152939
R16743 GND.n5374 GND.n1866 0.152939
R16744 GND.n5391 GND.n1866 0.152939
R16745 GND.n5392 GND.n5391 0.152939
R16746 GND.n5393 GND.n5392 0.152939
R16747 GND.n5393 GND.n1863 0.152939
R16748 GND.n5399 GND.n1863 0.152939
R16749 GND.n5400 GND.n5399 0.152939
R16750 GND.n5401 GND.n5400 0.152939
R16751 GND.n5401 GND.n1859 0.152939
R16752 GND.n5409 GND.n1859 0.152939
R16753 GND.n5410 GND.n5409 0.152939
R16754 GND.n5411 GND.n5410 0.152939
R16755 GND.n5412 GND.n5411 0.152939
R16756 GND.n5413 GND.n5412 0.152939
R16757 GND.n5428 GND.n5413 0.152939
R16758 GND.n5429 GND.n5428 0.152939
R16759 GND.n5430 GND.n5429 0.152939
R16760 GND.n5431 GND.n5430 0.152939
R16761 GND.n5523 GND.n5431 0.152939
R16762 GND.n5524 GND.n5523 0.152939
R16763 GND.n5525 GND.n5524 0.152939
R16764 GND.n5526 GND.n5525 0.152939
R16765 GND.n5527 GND.n5526 0.152939
R16766 GND.n5542 GND.n5527 0.152939
R16767 GND.n5543 GND.n5542 0.152939
R16768 GND.n5544 GND.n5543 0.152939
R16769 GND.n5545 GND.n5544 0.152939
R16770 GND.n5560 GND.n5545 0.152939
R16771 GND.n5561 GND.n5560 0.152939
R16772 GND.n5562 GND.n5561 0.152939
R16773 GND.n5563 GND.n5562 0.152939
R16774 GND.n5578 GND.n5563 0.152939
R16775 GND.n5579 GND.n5578 0.152939
R16776 GND.n5580 GND.n5579 0.152939
R16777 GND.n5581 GND.n5580 0.152939
R16778 GND.n5654 GND.n5581 0.152939
R16779 GND.n5655 GND.n5654 0.152939
R16780 GND.n5656 GND.n5655 0.152939
R16781 GND.n5657 GND.n5656 0.152939
R16782 GND.n5658 GND.n5657 0.152939
R16783 GND.n5673 GND.n5658 0.152939
R16784 GND.n5674 GND.n5673 0.152939
R16785 GND.n5675 GND.n5674 0.152939
R16786 GND.n5676 GND.n5675 0.152939
R16787 GND.n5691 GND.n5676 0.152939
R16788 GND.n5692 GND.n5691 0.152939
R16789 GND.n5693 GND.n5692 0.152939
R16790 GND.n5694 GND.n5693 0.152939
R16791 GND.n5709 GND.n5694 0.152939
R16792 GND.n5710 GND.n5709 0.152939
R16793 GND.n5711 GND.n5710 0.152939
R16794 GND.n5712 GND.n5711 0.152939
R16795 GND.n5785 GND.n5712 0.152939
R16796 GND.n5786 GND.n5785 0.152939
R16797 GND.n5787 GND.n5786 0.152939
R16798 GND.n5788 GND.n5787 0.152939
R16799 GND.n5789 GND.n5788 0.152939
R16800 GND.n5803 GND.n5789 0.152939
R16801 GND.n5804 GND.n5803 0.152939
R16802 GND.n5805 GND.n5804 0.152939
R16803 GND.n5806 GND.n5805 0.152939
R16804 GND.n5821 GND.n5806 0.152939
R16805 GND.n5822 GND.n5821 0.152939
R16806 GND.n5823 GND.n5822 0.152939
R16807 GND.n5824 GND.n5823 0.152939
R16808 GND.n5839 GND.n5824 0.152939
R16809 GND.n5840 GND.n5839 0.152939
R16810 GND.n5841 GND.n5840 0.152939
R16811 GND.n5842 GND.n5841 0.152939
R16812 GND.n5916 GND.n5842 0.152939
R16813 GND.n5917 GND.n5916 0.152939
R16814 GND.n5918 GND.n5917 0.152939
R16815 GND.n5919 GND.n5918 0.152939
R16816 GND.n5920 GND.n5919 0.152939
R16817 GND.n5954 GND.n5920 0.152939
R16818 GND.n5955 GND.n5954 0.152939
R16819 GND.n5956 GND.n5955 0.152939
R16820 GND.n5956 GND.n1583 0.152939
R16821 GND.n6434 GND.n1583 0.152939
R16822 GND.n6435 GND.n6434 0.152939
R16823 GND.n6436 GND.n6435 0.152939
R16824 GND.n6437 GND.n6436 0.152939
R16825 GND.n6437 GND.n1552 0.152939
R16826 GND.n6471 GND.n1552 0.152939
R16827 GND.n6472 GND.n6471 0.152939
R16828 GND.n6473 GND.n6472 0.152939
R16829 GND.n6474 GND.n6473 0.152939
R16830 GND.n6475 GND.n6474 0.152939
R16831 GND.n6475 GND.n1514 0.152939
R16832 GND.n6531 GND.n1514 0.152939
R16833 GND.n6532 GND.n6531 0.152939
R16834 GND.n6533 GND.n6532 0.152939
R16835 GND.n6534 GND.n6533 0.152939
R16836 GND.n6535 GND.n6534 0.152939
R16837 GND.n6536 GND.n6535 0.152939
R16838 GND.n6536 GND.n1471 0.152939
R16839 GND.n6609 GND.n1471 0.152939
R16840 GND.n6610 GND.n6609 0.152939
R16841 GND.n6611 GND.n6610 0.152939
R16842 GND.n6612 GND.n6611 0.152939
R16843 GND.n6613 GND.n6612 0.152939
R16844 GND.n6613 GND.n1416 0.152939
R16845 GND.n6688 GND.n1416 0.152939
R16846 GND.n6689 GND.n6688 0.152939
R16847 GND.n6690 GND.n6689 0.152939
R16848 GND.n6690 GND.n1393 0.152939
R16849 GND.n6717 GND.n1393 0.152939
R16850 GND.n6718 GND.n6717 0.152939
R16851 GND.n6719 GND.n6718 0.152939
R16852 GND.n6720 GND.n6719 0.152939
R16853 GND.n6721 GND.n6720 0.152939
R16854 GND.n6724 GND.n6721 0.152939
R16855 GND.n6725 GND.n6724 0.152939
R16856 GND.n6726 GND.n6725 0.152939
R16857 GND.n6727 GND.n6726 0.152939
R16858 GND.n6730 GND.n6727 0.152939
R16859 GND.n6731 GND.n6730 0.152939
R16860 GND.n6732 GND.n6731 0.152939
R16861 GND.n6733 GND.n6732 0.152939
R16862 GND.n6733 GND.n1305 0.152939
R16863 GND.n6890 GND.n1305 0.152939
R16864 GND.n6891 GND.n6890 0.152939
R16865 GND.n6892 GND.n6891 0.152939
R16866 GND.n6893 GND.n6892 0.152939
R16867 GND.n6894 GND.n6893 0.152939
R16868 GND.n6897 GND.n6894 0.152939
R16869 GND.n6898 GND.n6897 0.152939
R16870 GND.n6899 GND.n6898 0.152939
R16871 GND.n6899 GND.n1152 0.152939
R16872 GND.n7013 GND.n1152 0.152939
R16873 GND.n7014 GND.n7013 0.152939
R16874 GND.n7015 GND.n7014 0.152939
R16875 GND.n7016 GND.n7015 0.152939
R16876 GND.n7017 GND.n7016 0.152939
R16877 GND.n7018 GND.n7017 0.152939
R16878 GND.n7018 GND.n1121 0.152939
R16879 GND.n7059 GND.n1121 0.152939
R16880 GND.n7060 GND.n7059 0.152939
R16881 GND.n7061 GND.n7060 0.152939
R16882 GND.n7062 GND.n7061 0.152939
R16883 GND.n7063 GND.n7062 0.152939
R16884 GND.n7065 GND.n7063 0.152939
R16885 GND.n7066 GND.n7065 0.152939
R16886 GND.n7066 GND.n1087 0.152939
R16887 GND.n7117 GND.n1087 0.152939
R16888 GND.n7118 GND.n7117 0.152939
R16889 GND.n7119 GND.n7118 0.152939
R16890 GND.n7120 GND.n7119 0.152939
R16891 GND.n7120 GND.n1062 0.152939
R16892 GND.n7152 GND.n1062 0.152939
R16893 GND.n7153 GND.n7152 0.152939
R16894 GND.n7154 GND.n7153 0.152939
R16895 GND.n7155 GND.n7154 0.152939
R16896 GND.n7156 GND.n7155 0.152939
R16897 GND.n7156 GND.n1038 0.152939
R16898 GND.n7191 GND.n1038 0.152939
R16899 GND.n7192 GND.n7191 0.152939
R16900 GND.n7193 GND.n7192 0.152939
R16901 GND.n7194 GND.n7193 0.152939
R16902 GND.n7195 GND.n7194 0.152939
R16903 GND.n7197 GND.n7195 0.152939
R16904 GND.n7198 GND.n7197 0.152939
R16905 GND.n7198 GND.n1004 0.152939
R16906 GND.n7249 GND.n1004 0.152939
R16907 GND.n7250 GND.n7249 0.152939
R16908 GND.n7251 GND.n7250 0.152939
R16909 GND.n7252 GND.n7251 0.152939
R16910 GND.n7252 GND.n979 0.152939
R16911 GND.n7284 GND.n979 0.152939
R16912 GND.n7285 GND.n7284 0.152939
R16913 GND.n7286 GND.n7285 0.152939
R16914 GND.n7287 GND.n7286 0.152939
R16915 GND.n7288 GND.n7287 0.152939
R16916 GND.n7288 GND.n954 0.152939
R16917 GND.n7322 GND.n954 0.152939
R16918 GND.n7323 GND.n7322 0.152939
R16919 GND.n7324 GND.n7323 0.152939
R16920 GND.n7325 GND.n7324 0.152939
R16921 GND.n7325 GND.n929 0.152939
R16922 GND.n7357 GND.n929 0.152939
R16923 GND.n7358 GND.n7357 0.152939
R16924 GND.n7359 GND.n7358 0.152939
R16925 GND.n7359 GND.n912 0.152939
R16926 GND.n7381 GND.n912 0.152939
R16927 GND.n7382 GND.n7381 0.152939
R16928 GND.n7383 GND.n7382 0.152939
R16929 GND.n7384 GND.n7383 0.152939
R16930 GND.n7384 GND.n889 0.152939
R16931 GND.n7417 GND.n889 0.152939
R16932 GND.n7418 GND.n7417 0.152939
R16933 GND.n7419 GND.n7418 0.152939
R16934 GND.n7419 GND.n872 0.152939
R16935 GND.n7487 GND.n872 0.152939
R16936 GND.n7488 GND.n7487 0.152939
R16937 GND.n7489 GND.n7488 0.152939
R16938 GND.n7490 GND.n7489 0.152939
R16939 GND.n7491 GND.n7490 0.152939
R16940 GND.n7493 GND.n7491 0.152939
R16941 GND.n7494 GND.n7493 0.152939
R16942 GND.n7494 GND.n676 0.152939
R16943 GND.n7705 GND.n676 0.152939
R16944 GND.n7706 GND.n7705 0.152939
R16945 GND.n7707 GND.n7706 0.152939
R16946 GND.n7707 GND.n655 0.152939
R16947 GND.n7727 GND.n655 0.152939
R16948 GND.n7728 GND.n7727 0.152939
R16949 GND.n7729 GND.n7728 0.152939
R16950 GND.n7729 GND.n635 0.152939
R16951 GND.n7747 GND.n635 0.152939
R16952 GND.n7748 GND.n7747 0.152939
R16953 GND.n7749 GND.n7748 0.152939
R16954 GND.n7749 GND.n615 0.152939
R16955 GND.n7767 GND.n615 0.152939
R16956 GND.n7768 GND.n7767 0.152939
R16957 GND.n7769 GND.n7768 0.152939
R16958 GND.n7769 GND.n595 0.152939
R16959 GND.n7787 GND.n595 0.152939
R16960 GND.n7788 GND.n7787 0.152939
R16961 GND.n7789 GND.n7788 0.152939
R16962 GND.n7789 GND.n574 0.152939
R16963 GND.n7811 GND.n574 0.152939
R16964 GND.n7812 GND.n7811 0.152939
R16965 GND.n7813 GND.n7812 0.152939
R16966 GND.n7814 GND.n7813 0.152939
R16967 GND.n7814 GND.n547 0.152939
R16968 GND.n7885 GND.n547 0.152939
R16969 GND.n7886 GND.n7885 0.152939
R16970 GND.n7887 GND.n7886 0.152939
R16971 GND.n7887 GND.n527 0.152939
R16972 GND.n7905 GND.n527 0.152939
R16973 GND.n7906 GND.n7905 0.152939
R16974 GND.n7907 GND.n7906 0.152939
R16975 GND.n7907 GND.n507 0.152939
R16976 GND.n7925 GND.n507 0.152939
R16977 GND.n7926 GND.n7925 0.152939
R16978 GND.n7927 GND.n7926 0.152939
R16979 GND.n7927 GND.n486 0.152939
R16980 GND.n7952 GND.n486 0.152939
R16981 GND.n7953 GND.n7952 0.152939
R16982 GND.n7954 GND.n7953 0.152939
R16983 GND.n7954 GND.n116 0.152939
R16984 GND.n8603 GND.n116 0.152939
R16985 GND.n8604 GND.n8603 0.152939
R16986 GND.n8605 GND.n8604 0.152939
R16987 GND.n8605 GND.n83 0.152939
R16988 GND.n8633 GND.n83 0.152939
R16989 GND.n5085 GND.n2085 0.152939
R16990 GND.n2093 GND.n2085 0.152939
R16991 GND.n2094 GND.n2093 0.152939
R16992 GND.n2095 GND.n2094 0.152939
R16993 GND.n2096 GND.n2095 0.152939
R16994 GND.n2097 GND.n2096 0.152939
R16995 GND.n2098 GND.n2097 0.152939
R16996 GND.n2099 GND.n2098 0.152939
R16997 GND.n2100 GND.n2099 0.152939
R16998 GND.n2101 GND.n2100 0.152939
R16999 GND.n2102 GND.n2101 0.152939
R17000 GND.n2103 GND.n2102 0.152939
R17001 GND.n2104 GND.n2103 0.152939
R17002 GND.n2105 GND.n2104 0.152939
R17003 GND.n2106 GND.n2105 0.152939
R17004 GND.n2107 GND.n2106 0.152939
R17005 GND.n2108 GND.n2107 0.152939
R17006 GND.n2109 GND.n2108 0.152939
R17007 GND.n2110 GND.n2109 0.152939
R17008 GND.n2111 GND.n2110 0.152939
R17009 GND.n2112 GND.n2111 0.152939
R17010 GND.n2113 GND.n2112 0.152939
R17011 GND.n2114 GND.n2113 0.152939
R17012 GND.n2115 GND.n2114 0.152939
R17013 GND.n2116 GND.n2115 0.152939
R17014 GND.n2117 GND.n2116 0.152939
R17015 GND.n2118 GND.n2117 0.152939
R17016 GND.n2119 GND.n2118 0.152939
R17017 GND.n2120 GND.n2119 0.152939
R17018 GND.n2121 GND.n2120 0.152939
R17019 GND.n2122 GND.n2121 0.152939
R17020 GND.n2123 GND.n2122 0.152939
R17021 GND.n2124 GND.n2123 0.152939
R17022 GND.n2125 GND.n2124 0.152939
R17023 GND.n2126 GND.n2125 0.152939
R17024 GND.n2127 GND.n2126 0.152939
R17025 GND.n2128 GND.n2127 0.152939
R17026 GND.n2129 GND.n2128 0.152939
R17027 GND.n2130 GND.n2129 0.152939
R17028 GND.n2131 GND.n2130 0.152939
R17029 GND.n2132 GND.n2131 0.152939
R17030 GND.n2133 GND.n2132 0.152939
R17031 GND.n2133 GND.n1691 0.152939
R17032 GND.n2468 GND.n2467 0.152939
R17033 GND.n2469 GND.n2468 0.152939
R17034 GND.n2470 GND.n2469 0.152939
R17035 GND.n2471 GND.n2470 0.152939
R17036 GND.n2472 GND.n2471 0.152939
R17037 GND.n2473 GND.n2472 0.152939
R17038 GND.n2474 GND.n2473 0.152939
R17039 GND.n2475 GND.n2474 0.152939
R17040 GND.n2476 GND.n2475 0.152939
R17041 GND.n2479 GND.n2476 0.152939
R17042 GND.n2480 GND.n2479 0.152939
R17043 GND.n2481 GND.n2480 0.152939
R17044 GND.n2482 GND.n2481 0.152939
R17045 GND.n2483 GND.n2482 0.152939
R17046 GND.n2484 GND.n2483 0.152939
R17047 GND.n2485 GND.n2484 0.152939
R17048 GND.n2486 GND.n2485 0.152939
R17049 GND.n2487 GND.n2486 0.152939
R17050 GND.n2488 GND.n2487 0.152939
R17051 GND.n2490 GND.n2488 0.152939
R17052 GND.n2493 GND.n2490 0.152939
R17053 GND.n2494 GND.n2493 0.152939
R17054 GND.n2495 GND.n2494 0.152939
R17055 GND.n2496 GND.n2495 0.152939
R17056 GND.n2497 GND.n2496 0.152939
R17057 GND.n2498 GND.n2497 0.152939
R17058 GND.n2499 GND.n2498 0.152939
R17059 GND.n2500 GND.n2499 0.152939
R17060 GND.n2501 GND.n2500 0.152939
R17061 GND.n2502 GND.n2501 0.152939
R17062 GND.n2503 GND.n2502 0.152939
R17063 GND.n2506 GND.n2503 0.152939
R17064 GND.n2507 GND.n2506 0.152939
R17065 GND.n2508 GND.n2507 0.152939
R17066 GND.n2509 GND.n2508 0.152939
R17067 GND.n2510 GND.n2509 0.152939
R17068 GND.n2511 GND.n2510 0.152939
R17069 GND.n2512 GND.n2511 0.152939
R17070 GND.n2513 GND.n2512 0.152939
R17071 GND.n2514 GND.n2513 0.152939
R17072 GND.n2515 GND.n2514 0.152939
R17073 GND.n2517 GND.n2515 0.152939
R17074 GND.n2520 GND.n2517 0.152939
R17075 GND.n2521 GND.n2520 0.152939
R17076 GND.n2522 GND.n2521 0.152939
R17077 GND.n2523 GND.n2522 0.152939
R17078 GND.n2524 GND.n2523 0.152939
R17079 GND.n2525 GND.n2524 0.152939
R17080 GND.n2526 GND.n2525 0.152939
R17081 GND.n2527 GND.n2526 0.152939
R17082 GND.n2528 GND.n2527 0.152939
R17083 GND.n2529 GND.n2528 0.152939
R17084 GND.n2869 GND.n2529 0.152939
R17085 GND.n2869 GND.n2868 0.152939
R17086 GND.n2568 GND.n2567 0.152939
R17087 GND.n2616 GND.n2567 0.152939
R17088 GND.n2617 GND.n2616 0.152939
R17089 GND.n2618 GND.n2617 0.152939
R17090 GND.n2619 GND.n2618 0.152939
R17091 GND.n2620 GND.n2619 0.152939
R17092 GND.n2621 GND.n2620 0.152939
R17093 GND.n2622 GND.n2621 0.152939
R17094 GND.n2623 GND.n2622 0.152939
R17095 GND.n2624 GND.n2623 0.152939
R17096 GND.n2625 GND.n2624 0.152939
R17097 GND.n2626 GND.n2625 0.152939
R17098 GND.n2627 GND.n2626 0.152939
R17099 GND.n2628 GND.n2627 0.152939
R17100 GND.n2629 GND.n2628 0.152939
R17101 GND.n2630 GND.n2629 0.152939
R17102 GND.n2631 GND.n2630 0.152939
R17103 GND.n2632 GND.n2631 0.152939
R17104 GND.n2633 GND.n2632 0.152939
R17105 GND.n2634 GND.n2633 0.152939
R17106 GND.n2635 GND.n2634 0.152939
R17107 GND.n2636 GND.n2635 0.152939
R17108 GND.n2637 GND.n2636 0.152939
R17109 GND.n2638 GND.n2637 0.152939
R17110 GND.n2639 GND.n2638 0.152939
R17111 GND.n2640 GND.n2639 0.152939
R17112 GND.n2641 GND.n2640 0.152939
R17113 GND.n2642 GND.n2641 0.152939
R17114 GND.n2643 GND.n2642 0.152939
R17115 GND.n2644 GND.n2643 0.152939
R17116 GND.n2645 GND.n2644 0.152939
R17117 GND.n2646 GND.n2645 0.152939
R17118 GND.n2647 GND.n2646 0.152939
R17119 GND.n2648 GND.n2647 0.152939
R17120 GND.n2649 GND.n2648 0.152939
R17121 GND.n2650 GND.n2649 0.152939
R17122 GND.n2651 GND.n2650 0.152939
R17123 GND.n2652 GND.n2651 0.152939
R17124 GND.n2653 GND.n2652 0.152939
R17125 GND.n2654 GND.n2653 0.152939
R17126 GND.n2655 GND.n2654 0.152939
R17127 GND.n2655 GND.n2086 0.152939
R17128 GND.n5085 GND.n2086 0.152939
R17129 GND.n4849 GND.n4848 0.152939
R17130 GND.n4849 GND.n2410 0.152939
R17131 GND.n4867 GND.n2410 0.152939
R17132 GND.n4868 GND.n4867 0.152939
R17133 GND.n4869 GND.n4868 0.152939
R17134 GND.n4869 GND.n2390 0.152939
R17135 GND.n4887 GND.n2390 0.152939
R17136 GND.n4888 GND.n4887 0.152939
R17137 GND.n4889 GND.n4888 0.152939
R17138 GND.n4889 GND.n2370 0.152939
R17139 GND.n4907 GND.n2370 0.152939
R17140 GND.n4908 GND.n4907 0.152939
R17141 GND.n4909 GND.n4908 0.152939
R17142 GND.n4909 GND.n2349 0.152939
R17143 GND.n4927 GND.n2349 0.152939
R17144 GND.n4928 GND.n4927 0.152939
R17145 GND.n4929 GND.n4928 0.152939
R17146 GND.n4929 GND.n2330 0.152939
R17147 GND.n4947 GND.n2330 0.152939
R17148 GND.n4948 GND.n4947 0.152939
R17149 GND.n4949 GND.n4948 0.152939
R17150 GND.n4949 GND.n2310 0.152939
R17151 GND.n4967 GND.n2310 0.152939
R17152 GND.n4968 GND.n4967 0.152939
R17153 GND.n4969 GND.n4968 0.152939
R17154 GND.n4969 GND.n2290 0.152939
R17155 GND.n4987 GND.n2290 0.152939
R17156 GND.n4988 GND.n4987 0.152939
R17157 GND.n4989 GND.n4988 0.152939
R17158 GND.n4989 GND.n2270 0.152939
R17159 GND.n5007 GND.n2270 0.152939
R17160 GND.n5008 GND.n5007 0.152939
R17161 GND.n5010 GND.n5008 0.152939
R17162 GND.n5010 GND.n5009 0.152939
R17163 GND.n5009 GND.n2250 0.152939
R17164 GND.n2250 GND.n2079 0.152939
R17165 GND.n5086 GND.n2079 0.152939
R17166 GND.n4727 GND.n3020 0.152939
R17167 GND.n4735 GND.n3020 0.152939
R17168 GND.n4736 GND.n4735 0.152939
R17169 GND.n4737 GND.n4736 0.152939
R17170 GND.n4737 GND.n3016 0.152939
R17171 GND.n4745 GND.n3016 0.152939
R17172 GND.n4746 GND.n4745 0.152939
R17173 GND.n4747 GND.n4746 0.152939
R17174 GND.n4747 GND.n3012 0.152939
R17175 GND.n4755 GND.n3012 0.152939
R17176 GND.n4756 GND.n4755 0.152939
R17177 GND.n4757 GND.n4756 0.152939
R17178 GND.n4757 GND.n3008 0.152939
R17179 GND.n4765 GND.n3008 0.152939
R17180 GND.n4766 GND.n4765 0.152939
R17181 GND.n4767 GND.n4766 0.152939
R17182 GND.n4767 GND.n3004 0.152939
R17183 GND.n4775 GND.n3004 0.152939
R17184 GND.n4776 GND.n4775 0.152939
R17185 GND.n4777 GND.n4776 0.152939
R17186 GND.n4777 GND.n3000 0.152939
R17187 GND.n4785 GND.n3000 0.152939
R17188 GND.n4786 GND.n4785 0.152939
R17189 GND.n4787 GND.n4786 0.152939
R17190 GND.n4787 GND.n2996 0.152939
R17191 GND.n4795 GND.n2996 0.152939
R17192 GND.n4796 GND.n4795 0.152939
R17193 GND.n4797 GND.n4796 0.152939
R17194 GND.n4797 GND.n2992 0.152939
R17195 GND.n4805 GND.n2992 0.152939
R17196 GND.n4806 GND.n4805 0.152939
R17197 GND.n4807 GND.n4806 0.152939
R17198 GND.n4807 GND.n2988 0.152939
R17199 GND.n4815 GND.n2988 0.152939
R17200 GND.n4816 GND.n4815 0.152939
R17201 GND.n4817 GND.n4816 0.152939
R17202 GND.n4817 GND.n2984 0.152939
R17203 GND.n4825 GND.n2984 0.152939
R17204 GND.n4826 GND.n4825 0.152939
R17205 GND.n4827 GND.n4826 0.152939
R17206 GND.n4827 GND.n2980 0.152939
R17207 GND.n4835 GND.n2980 0.152939
R17208 GND.n4836 GND.n4835 0.152939
R17209 GND.n4838 GND.n4836 0.152939
R17210 GND.n4838 GND.n4837 0.152939
R17211 GND.n4837 GND.n2429 0.152939
R17212 GND.n4847 GND.n2429 0.152939
R17213 GND.n6279 GND.n6278 0.152939
R17214 GND.n6278 GND.n6277 0.152939
R17215 GND.n6277 GND.n1692 0.152939
R17216 GND.n6273 GND.n1692 0.152939
R17217 GND.n6273 GND.n6272 0.152939
R17218 GND.n6272 GND.n6271 0.152939
R17219 GND.n6271 GND.n1698 0.152939
R17220 GND.n6267 GND.n1698 0.152939
R17221 GND.n6267 GND.n6266 0.152939
R17222 GND.n6266 GND.n6265 0.152939
R17223 GND.n6265 GND.n1706 0.152939
R17224 GND.n6261 GND.n1706 0.152939
R17225 GND.n6261 GND.n6260 0.152939
R17226 GND.n6260 GND.n6259 0.152939
R17227 GND.n6259 GND.n1712 0.152939
R17228 GND.n6255 GND.n1712 0.152939
R17229 GND.n6255 GND.n6254 0.152939
R17230 GND.n6254 GND.n6253 0.152939
R17231 GND.n6253 GND.n1718 0.152939
R17232 GND.n1723 GND.n1718 0.152939
R17233 GND.n6248 GND.n1723 0.152939
R17234 GND.n6248 GND.n6247 0.152939
R17235 GND.n6247 GND.n6246 0.152939
R17236 GND.n1817 GND.n1816 0.152939
R17237 GND.n1816 GND.n1815 0.152939
R17238 GND.n1815 GND.n1731 0.152939
R17239 GND.n1811 GND.n1731 0.152939
R17240 GND.n1811 GND.n1810 0.152939
R17241 GND.n1810 GND.n1809 0.152939
R17242 GND.n1809 GND.n1739 0.152939
R17243 GND.n1805 GND.n1739 0.152939
R17244 GND.n1805 GND.n1804 0.152939
R17245 GND.n1804 GND.n1803 0.152939
R17246 GND.n1803 GND.n1745 0.152939
R17247 GND.n1799 GND.n1745 0.152939
R17248 GND.n1799 GND.n1798 0.152939
R17249 GND.n1798 GND.n1797 0.152939
R17250 GND.n1797 GND.n1751 0.152939
R17251 GND.n1756 GND.n1751 0.152939
R17252 GND.n1792 GND.n1756 0.152939
R17253 GND.n1792 GND.n1791 0.152939
R17254 GND.n1791 GND.n1790 0.152939
R17255 GND.n1790 GND.n1760 0.152939
R17256 GND.n1786 GND.n1760 0.152939
R17257 GND.n1786 GND.n1785 0.152939
R17258 GND.n1785 GND.n1784 0.152939
R17259 GND.n1784 GND.n1766 0.152939
R17260 GND.n1780 GND.n1766 0.152939
R17261 GND.n1780 GND.n1779 0.152939
R17262 GND.n1779 GND.n1778 0.152939
R17263 GND.n1778 GND.n1624 0.152939
R17264 GND.n2866 GND.n2534 0.152939
R17265 GND.n2589 GND.n2534 0.152939
R17266 GND.n2590 GND.n2589 0.152939
R17267 GND.n2591 GND.n2590 0.152939
R17268 GND.n2591 GND.n2582 0.152939
R17269 GND.n2597 GND.n2582 0.152939
R17270 GND.n2598 GND.n2597 0.152939
R17271 GND.n2599 GND.n2598 0.152939
R17272 GND.n2599 GND.n2575 0.152939
R17273 GND.n2603 GND.n2575 0.152939
R17274 GND.n2607 GND.n2606 0.152939
R17275 GND.n2608 GND.n2607 0.152939
R17276 GND.n2608 GND.n2557 0.152939
R17277 GND.n2719 GND.n2557 0.152939
R17278 GND.n2720 GND.n2719 0.152939
R17279 GND.n2845 GND.n2720 0.152939
R17280 GND.n2845 GND.n2844 0.152939
R17281 GND.n2844 GND.n2843 0.152939
R17282 GND.n2843 GND.n2721 0.152939
R17283 GND.n2839 GND.n2721 0.152939
R17284 GND.n2839 GND.n2838 0.152939
R17285 GND.n2838 GND.n2837 0.152939
R17286 GND.n2837 GND.n2725 0.152939
R17287 GND.n2833 GND.n2725 0.152939
R17288 GND.n2833 GND.n2832 0.152939
R17289 GND.n2832 GND.n2831 0.152939
R17290 GND.n2831 GND.n2729 0.152939
R17291 GND.n2827 GND.n2729 0.152939
R17292 GND.n2827 GND.n2826 0.152939
R17293 GND.n2826 GND.n2825 0.152939
R17294 GND.n2825 GND.n2733 0.152939
R17295 GND.n2821 GND.n2733 0.152939
R17296 GND.n2821 GND.n2820 0.152939
R17297 GND.n2820 GND.n2819 0.152939
R17298 GND.n2819 GND.n2737 0.152939
R17299 GND.n2815 GND.n2737 0.152939
R17300 GND.n2815 GND.n2814 0.152939
R17301 GND.n2814 GND.n2813 0.152939
R17302 GND.n2813 GND.n2741 0.152939
R17303 GND.n2809 GND.n2741 0.152939
R17304 GND.n2809 GND.n2808 0.152939
R17305 GND.n2808 GND.n2807 0.152939
R17306 GND.n2807 GND.n2745 0.152939
R17307 GND.n2803 GND.n2745 0.152939
R17308 GND.n2803 GND.n2802 0.152939
R17309 GND.n2802 GND.n2801 0.152939
R17310 GND.n2801 GND.n2749 0.152939
R17311 GND.n2797 GND.n2749 0.152939
R17312 GND.n2797 GND.n2796 0.152939
R17313 GND.n2796 GND.n2795 0.152939
R17314 GND.n2795 GND.n2753 0.152939
R17315 GND.n2791 GND.n2753 0.152939
R17316 GND.n2791 GND.n2790 0.152939
R17317 GND.n2790 GND.n2789 0.152939
R17318 GND.n2789 GND.n2758 0.152939
R17319 GND.n2785 GND.n2758 0.152939
R17320 GND.n2785 GND.n2784 0.152939
R17321 GND.n2783 GND.n2782 0.145814
R17322 GND.n8639 GND.n62 0.145814
R17323 GND.n8639 GND.n63 0.145814
R17324 GND.n2784 GND.n2783 0.145814
R17325 GND GND.n8641 0.128027
R17326 GND.n1275 GND.n1195 0.0767195
R17327 GND.n6369 GND.n1616 0.0767195
R17328 GND.n1274 GND.n668 0.063
R17329 GND.n6291 GND.n6290 0.063
R17330 GND.n7713 GND.n668 0.0548478
R17331 GND.n8332 GND.n8331 0.0548478
R17332 GND.n2867 GND.n2533 0.0548478
R17333 GND.n6290 GND.n6289 0.0548478
R17334 GND.n7714 GND.n7713 0.0344674
R17335 GND.n7714 GND.n665 0.0344674
R17336 GND.n7718 GND.n665 0.0344674
R17337 GND.n7719 GND.n7718 0.0344674
R17338 GND.n7719 GND.n647 0.0344674
R17339 GND.n647 GND.n645 0.0344674
R17340 GND.n7738 GND.n645 0.0344674
R17341 GND.n7739 GND.n7738 0.0344674
R17342 GND.n7739 GND.n627 0.0344674
R17343 GND.n627 GND.n625 0.0344674
R17344 GND.n7758 GND.n625 0.0344674
R17345 GND.n7759 GND.n7758 0.0344674
R17346 GND.n7759 GND.n607 0.0344674
R17347 GND.n607 GND.n605 0.0344674
R17348 GND.n7778 GND.n605 0.0344674
R17349 GND.n7779 GND.n7778 0.0344674
R17350 GND.n7779 GND.n587 0.0344674
R17351 GND.n587 GND.n584 0.0344674
R17352 GND.n585 GND.n584 0.0344674
R17353 GND.n7800 GND.n585 0.0344674
R17354 GND.n7801 GND.n7800 0.0344674
R17355 GND.n7801 GND.n558 0.0344674
R17356 GND.n558 GND.n556 0.0344674
R17357 GND.n7876 GND.n556 0.0344674
R17358 GND.n7877 GND.n7876 0.0344674
R17359 GND.n7877 GND.n539 0.0344674
R17360 GND.n539 GND.n537 0.0344674
R17361 GND.n7896 GND.n537 0.0344674
R17362 GND.n7897 GND.n7896 0.0344674
R17363 GND.n7897 GND.n519 0.0344674
R17364 GND.n519 GND.n517 0.0344674
R17365 GND.n7916 GND.n517 0.0344674
R17366 GND.n7917 GND.n7916 0.0344674
R17367 GND.n7917 GND.n499 0.0344674
R17368 GND.n499 GND.n496 0.0344674
R17369 GND.n497 GND.n496 0.0344674
R17370 GND.n7944 GND.n497 0.0344674
R17371 GND.n7944 GND.n7943 0.0344674
R17372 GND.n7943 GND.n126 0.0344674
R17373 GND.n127 GND.n126 0.0344674
R17374 GND.n8595 GND.n127 0.0344674
R17375 GND.n8595 GND.n8594 0.0344674
R17376 GND.n8594 GND.n96 0.0344674
R17377 GND.n97 GND.n96 0.0344674
R17378 GND.n98 GND.n97 0.0344674
R17379 GND.n129 GND.n98 0.0344674
R17380 GND.n130 GND.n129 0.0344674
R17381 GND.n131 GND.n130 0.0344674
R17382 GND.n132 GND.n131 0.0344674
R17383 GND.n8233 GND.n132 0.0344674
R17384 GND.n8234 GND.n8233 0.0344674
R17385 GND.n8234 GND.n147 0.0344674
R17386 GND.n148 GND.n147 0.0344674
R17387 GND.n149 GND.n148 0.0344674
R17388 GND.n8240 GND.n149 0.0344674
R17389 GND.n8240 GND.n167 0.0344674
R17390 GND.n168 GND.n167 0.0344674
R17391 GND.n169 GND.n168 0.0344674
R17392 GND.n8247 GND.n169 0.0344674
R17393 GND.n8247 GND.n187 0.0344674
R17394 GND.n188 GND.n187 0.0344674
R17395 GND.n189 GND.n188 0.0344674
R17396 GND.n8254 GND.n189 0.0344674
R17397 GND.n8254 GND.n209 0.0344674
R17398 GND.n210 GND.n209 0.0344674
R17399 GND.n211 GND.n210 0.0344674
R17400 GND.n8261 GND.n211 0.0344674
R17401 GND.n8261 GND.n230 0.0344674
R17402 GND.n231 GND.n230 0.0344674
R17403 GND.n232 GND.n231 0.0344674
R17404 GND.n8268 GND.n232 0.0344674
R17405 GND.n8268 GND.n251 0.0344674
R17406 GND.n252 GND.n251 0.0344674
R17407 GND.n253 GND.n252 0.0344674
R17408 GND.n8275 GND.n253 0.0344674
R17409 GND.n8275 GND.n272 0.0344674
R17410 GND.n273 GND.n272 0.0344674
R17411 GND.n274 GND.n273 0.0344674
R17412 GND.n8282 GND.n274 0.0344674
R17413 GND.n8282 GND.n293 0.0344674
R17414 GND.n294 GND.n293 0.0344674
R17415 GND.n295 GND.n294 0.0344674
R17416 GND.n8289 GND.n295 0.0344674
R17417 GND.n8289 GND.n314 0.0344674
R17418 GND.n315 GND.n314 0.0344674
R17419 GND.n316 GND.n315 0.0344674
R17420 GND.n8296 GND.n316 0.0344674
R17421 GND.n8296 GND.n335 0.0344674
R17422 GND.n336 GND.n335 0.0344674
R17423 GND.n337 GND.n336 0.0344674
R17424 GND.n8305 GND.n337 0.0344674
R17425 GND.n8306 GND.n8305 0.0344674
R17426 GND.n8306 GND.n8226 0.0344674
R17427 GND.n8311 GND.n8226 0.0344674
R17428 GND.n8311 GND.n445 0.0344674
R17429 GND.n8331 GND.n445 0.0344674
R17430 GND.n2860 GND.n2533 0.0344674
R17431 GND.n2860 GND.n2538 0.0344674
R17432 GND.n2856 GND.n2538 0.0344674
R17433 GND.n2856 GND.n2855 0.0344674
R17434 GND.n2855 GND.n2854 0.0344674
R17435 GND.n2854 GND.n2550 0.0344674
R17436 GND.n2850 GND.n2550 0.0344674
R17437 GND.n2850 GND.n2421 0.0344674
R17438 GND.n4861 GND.n2421 0.0344674
R17439 GND.n4861 GND.n4860 0.0344674
R17440 GND.n4860 GND.n4859 0.0344674
R17441 GND.n4859 GND.n2401 0.0344674
R17442 GND.n4881 GND.n2401 0.0344674
R17443 GND.n4881 GND.n4880 0.0344674
R17444 GND.n4880 GND.n4879 0.0344674
R17445 GND.n4879 GND.n2381 0.0344674
R17446 GND.n4901 GND.n2381 0.0344674
R17447 GND.n4901 GND.n4900 0.0344674
R17448 GND.n4900 GND.n4899 0.0344674
R17449 GND.n4899 GND.n2361 0.0344674
R17450 GND.n4921 GND.n2361 0.0344674
R17451 GND.n4921 GND.n4920 0.0344674
R17452 GND.n4920 GND.n4919 0.0344674
R17453 GND.n4919 GND.n2341 0.0344674
R17454 GND.n4941 GND.n2341 0.0344674
R17455 GND.n4941 GND.n4940 0.0344674
R17456 GND.n4940 GND.n4939 0.0344674
R17457 GND.n4939 GND.n2321 0.0344674
R17458 GND.n4961 GND.n2321 0.0344674
R17459 GND.n4961 GND.n4960 0.0344674
R17460 GND.n4960 GND.n4959 0.0344674
R17461 GND.n4959 GND.n2301 0.0344674
R17462 GND.n4981 GND.n2301 0.0344674
R17463 GND.n4981 GND.n4980 0.0344674
R17464 GND.n4980 GND.n4979 0.0344674
R17465 GND.n4979 GND.n2281 0.0344674
R17466 GND.n5001 GND.n2281 0.0344674
R17467 GND.n5001 GND.n5000 0.0344674
R17468 GND.n5000 GND.n4999 0.0344674
R17469 GND.n4999 GND.n2261 0.0344674
R17470 GND.n5027 GND.n2261 0.0344674
R17471 GND.n5027 GND.n5026 0.0344674
R17472 GND.n5026 GND.n5025 0.0344674
R17473 GND.n5025 GND.n5021 0.0344674
R17474 GND.n5021 GND.n2238 0.0344674
R17475 GND.n5047 GND.n2238 0.0344674
R17476 GND.n5047 GND.n5046 0.0344674
R17477 GND.n5046 GND.n5045 0.0344674
R17478 GND.n5045 GND.n2215 0.0344674
R17479 GND.n5072 GND.n2215 0.0344674
R17480 GND.n5072 GND.n5071 0.0344674
R17481 GND.n5071 GND.n5070 0.0344674
R17482 GND.n5070 GND.n5064 0.0344674
R17483 GND.n5066 GND.n5064 0.0344674
R17484 GND.n5066 GND.n2069 0.0344674
R17485 GND.n5104 GND.n2069 0.0344674
R17486 GND.n5104 GND.n5103 0.0344674
R17487 GND.n5103 GND.n5102 0.0344674
R17488 GND.n5102 GND.n5098 0.0344674
R17489 GND.n5098 GND.n2041 0.0344674
R17490 GND.n5195 GND.n2041 0.0344674
R17491 GND.n5195 GND.n5194 0.0344674
R17492 GND.n5194 GND.n5193 0.0344674
R17493 GND.n5193 GND.n2022 0.0344674
R17494 GND.n5215 GND.n2022 0.0344674
R17495 GND.n5215 GND.n5214 0.0344674
R17496 GND.n5214 GND.n5213 0.0344674
R17497 GND.n5213 GND.n2002 0.0344674
R17498 GND.n5235 GND.n2002 0.0344674
R17499 GND.n5235 GND.n5234 0.0344674
R17500 GND.n5234 GND.n5233 0.0344674
R17501 GND.n5233 GND.n1982 0.0344674
R17502 GND.n5255 GND.n1982 0.0344674
R17503 GND.n5255 GND.n5254 0.0344674
R17504 GND.n5254 GND.n5253 0.0344674
R17505 GND.n5253 GND.n1962 0.0344674
R17506 GND.n5275 GND.n1962 0.0344674
R17507 GND.n5275 GND.n5274 0.0344674
R17508 GND.n5274 GND.n5273 0.0344674
R17509 GND.n5273 GND.n1942 0.0344674
R17510 GND.n5295 GND.n1942 0.0344674
R17511 GND.n5295 GND.n5294 0.0344674
R17512 GND.n5294 GND.n5293 0.0344674
R17513 GND.n5293 GND.n1922 0.0344674
R17514 GND.n5320 GND.n1922 0.0344674
R17515 GND.n5320 GND.n5319 0.0344674
R17516 GND.n5319 GND.n5318 0.0344674
R17517 GND.n5318 GND.n5314 0.0344674
R17518 GND.n5314 GND.n1894 0.0344674
R17519 GND.n5365 GND.n1894 0.0344674
R17520 GND.n5365 GND.n5364 0.0344674
R17521 GND.n5364 GND.n5363 0.0344674
R17522 GND.n5363 GND.n1875 0.0344674
R17523 GND.n5384 GND.n1875 0.0344674
R17524 GND.n5384 GND.n1625 0.0344674
R17525 GND.n6289 GND.n1625 0.0344674
R17526 GND.n6371 GND.n6369 0.0248902
R17527 GND.n1286 GND.n1275 0.0248902
R17528 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t5 146.422
R17529 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t4 145.986
R17530 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t1 104.198
R17531 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t3 103.424
R17532 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t0 102.09
R17533 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t2 99.7677
R17534 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 5.41005
R17535 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 4.28744
R17536 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n0 4.16686
R17537 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 1.59564
R17538 DIFFPAIR_BIAS DIFFPAIR_BIAS.n4 0.683625
R17539 a_n7516_558.t24 a_n7516_558.n7 170.916
R17540 a_n7516_558.n7 a_n7516_558.t23 170.916
R17541 a_n7516_558.n1 a_n7516_558.t6 72.1419
R17542 a_n7516_558.n1 a_n7516_558.t14 72.1419
R17543 a_n7516_558.n3 a_n7516_558.t10 72.1419
R17544 a_n7516_558.n6 a_n7516_558.t25 72.1416
R17545 a_n7516_558.n0 a_n7516_558.t11 72.1416
R17546 a_n7516_558.n0 a_n7516_558.t16 72.1416
R17547 a_n7516_558.n5 a_n7516_558.t19 72.1416
R17548 a_n7516_558.n4 a_n7516_558.t20 72.1416
R17549 a_n7516_558.n4 a_n7516_558.n11 58.5336
R17550 a_n7516_558.n1 a_n7516_558.n10 58.5336
R17551 a_n7516_558.n1 a_n7516_558.n9 58.5336
R17552 a_n7516_558.n3 a_n7516_558.n8 58.5336
R17553 a_n7516_558.n6 a_n7516_558.n15 58.5334
R17554 a_n7516_558.n0 a_n7516_558.n14 58.5334
R17555 a_n7516_558.n0 a_n7516_558.n13 58.5334
R17556 a_n7516_558.n5 a_n7516_558.n12 58.5334
R17557 a_n7516_558.n15 a_n7516_558.t8 13.6087
R17558 a_n7516_558.n15 a_n7516_558.t3 13.6087
R17559 a_n7516_558.n14 a_n7516_558.t13 13.6087
R17560 a_n7516_558.n14 a_n7516_558.t15 13.6087
R17561 a_n7516_558.n13 a_n7516_558.t1 13.6087
R17562 a_n7516_558.n13 a_n7516_558.t5 13.6087
R17563 a_n7516_558.n12 a_n7516_558.t18 13.6087
R17564 a_n7516_558.n12 a_n7516_558.t7 13.6087
R17565 a_n7516_558.n11 a_n7516_558.t21 13.6087
R17566 a_n7516_558.n11 a_n7516_558.t17 13.6087
R17567 a_n7516_558.n10 a_n7516_558.t2 13.6087
R17568 a_n7516_558.n10 a_n7516_558.t0 13.6087
R17569 a_n7516_558.n9 a_n7516_558.t22 13.6087
R17570 a_n7516_558.n9 a_n7516_558.t4 13.6087
R17571 a_n7516_558.n8 a_n7516_558.t12 13.6087
R17572 a_n7516_558.n8 a_n7516_558.t9 13.6087
R17573 a_n7516_558.n3 a_n7516_558.n2 9.69061
R17574 a_n7516_558.n16 a_n7516_558.n4 9.69061
R17575 a_n7516_558.n7 a_n7516_558.n2 6.88079
R17576 a_n7516_558.n7 a_n7516_558.n16 6.75385
R17577 a_n7516_558.n5 a_n7516_558.n2 5.70955
R17578 a_n7516_558.n16 a_n7516_558.n6 5.70955
R17579 a_n7516_558.n4 a_n7516_558.n1 5.4459
R17580 a_n7516_558.n6 a_n7516_558.n0 5.4459
R17581 a_n7516_558.n0 a_n7516_558.n5 5.24188
R17582 a_n7516_558.n1 a_n7516_558.n3 5.24188
R17583 a_n11545_9494.n1 a_n11545_9494.t25 180.57
R17584 a_n11545_9494.n2 a_n11545_9494.t19 180.57
R17585 a_n11545_9494.n1 a_n11545_9494.t11 178.721
R17586 a_n11545_9494.n2 a_n11545_9494.t13 178.721
R17587 a_n11545_9494.n1 a_n11545_9494.n13 147.466
R17588 a_n11545_9494.n2 a_n11545_9494.n15 147.466
R17589 a_n11545_9494.t27 a_n11545_9494.n16 79.8687
R17590 a_n11545_9494.n12 a_n11545_9494.t1 79.8686
R17591 a_n11545_9494.n16 a_n11545_9494.t5 79.8684
R17592 a_n11545_9494.n12 a_n11545_9494.t3 78.1215
R17593 a_n11545_9494.n12 a_n11545_9494.t4 78.1215
R17594 a_n11545_9494.n16 a_n11545_9494.t9 78.1213
R17595 a_n11545_9494.n11 a_n11545_9494.n10 1.0888
R17596 a_n11545_9494.n16 a_n11545_9494.n12 35.6967
R17597 a_n11545_9494.n13 a_n11545_9494.t21 31.2553
R17598 a_n11545_9494.n13 a_n11545_9494.t17 31.2553
R17599 a_n11545_9494.n15 a_n11545_9494.t15 31.2553
R17600 a_n11545_9494.n15 a_n11545_9494.t23 31.2553
R17601 a_n11545_9494.n0 a_n11545_9494.t31 18.0625
R17602 a_n11545_9494.t43 a_n11545_9494.n0 34.165
R17603 a_n11545_9494.n0 a_n11545_9494.t38 18.0625
R17604 a_n11545_9494.t34 a_n11545_9494.n0 34.165
R17605 a_n11545_9494.n0 a_n11545_9494.t44 18.0625
R17606 a_n11545_9494.t45 a_n11545_9494.n0 34.165
R17607 a_n11545_9494.n0 a_n11545_9494.t35 18.0625
R17608 a_n11545_9494.t46 a_n11545_9494.n0 34.165
R17609 a_n11545_9494.n3 a_n11545_9494.n6 2.27663
R17610 a_n11545_9494.t10 a_n11545_9494.n3 34.165
R17611 a_n11545_9494.n4 a_n11545_9494.n5 2.27663
R17612 a_n11545_9494.t30 a_n11545_9494.n4 34.165
R17613 a_n11545_9494.n7 a_n11545_9494.n8 2.27663
R17614 a_n11545_9494.t29 a_n11545_9494.n7 34.165
R17615 a_n11545_9494.n9 a_n11545_9494.n14 64.2347
R17616 a_n11545_9494.n11 a_n11545_9494.n14 68.2777
R17617 a_n11545_9494.n11 a_n11545_9494.t18 31.6112
R17618 a_n11545_9494.n2 a_n11545_9494.n4 19.9107
R17619 a_n11545_9494.n7 a_n11545_9494.n0 19.4864
R17620 a_n11545_9494.n10 a_n11545_9494.n9 2.1671
R17621 a_n11545_9494.t9 a_n11545_9494.t2 13.6087
R17622 a_n11545_9494.t1 a_n11545_9494.t8 13.6087
R17623 a_n11545_9494.t3 a_n11545_9494.t26 13.6087
R17624 a_n11545_9494.t4 a_n11545_9494.t6 13.6087
R17625 a_n11545_9494.t5 a_n11545_9494.t7 13.6087
R17626 a_n11545_9494.t0 a_n11545_9494.t27 13.6087
R17627 a_n11545_9494.n4 a_n11545_9494.n3 9.81709
R17628 a_n11545_9494.n10 a_n11545_9494.n7 9.81709
R17629 a_n11545_9494.n0 a_n11545_9494.t41 42.7341
R17630 a_n11545_9494.n0 a_n11545_9494.t32 39.6989
R17631 a_n11545_9494.n0 a_n11545_9494.t28 42.8653
R17632 a_n11545_9494.n0 a_n11545_9494.t49 39.6315
R17633 a_n11545_9494.n0 a_n11545_9494.t36 42.7341
R17634 a_n11545_9494.n0 a_n11545_9494.t50 39.6989
R17635 a_n11545_9494.n0 a_n11545_9494.t48 42.8653
R17636 a_n11545_9494.n0 a_n11545_9494.t51 39.6315
R17637 a_n11545_9494.n6 a_n11545_9494.t20 43.001
R17638 a_n11545_9494.n6 a_n11545_9494.t16 39.5619
R17639 a_n11545_9494.n5 a_n11545_9494.t42 43.001
R17640 a_n11545_9494.n5 a_n11545_9494.t37 39.5619
R17641 a_n11545_9494.n8 a_n11545_9494.t47 43.001
R17642 a_n11545_9494.n8 a_n11545_9494.t33 39.5619
R17643 a_n11545_9494.n9 a_n11545_9494.t14 39.9643
R17644 a_n11545_9494.n14 a_n11545_9494.t22 8.6882
R17645 a_n11545_9494.n3 a_n11545_9494.t24 32.2029
R17646 a_n11545_9494.n4 a_n11545_9494.t40 32.2029
R17647 a_n11545_9494.n7 a_n11545_9494.t39 32.2029
R17648 a_n11545_9494.n12 a_n11545_9494.n10 25.7305
R17649 a_n11545_9494.n10 a_n11545_9494.t12 31.8746
R17650 a_n11545_9494.n3 a_n11545_9494.n0 28.7282
R17651 a_n11545_9494.n2 a_n11545_9494.n10 28.5036
R17652 a_n11545_9494.n0 a_n11545_9494.n1 23.6384
R17653 a_n11545_9494.n0 a_n11545_9494.n2 17.9267
R17654 a_n11689_9690.n0 a_n11689_9690.t15 180.57
R17655 a_n11689_9690.n1 a_n11689_9690.t1 178.721
R17656 a_n11689_9690.n0 a_n11689_9690.t14 178.721
R17657 a_n11689_9690.n0 a_n11689_9690.t3 178.721
R17658 a_n11689_9690.n10 a_n11689_9690.n9 168.901
R17659 a_n11689_9690.n4 a_n11689_9690.n2 167.858
R17660 a_n11689_9690.n4 a_n11689_9690.n3 167.054
R17661 a_n11689_9690.n9 a_n11689_9690.n8 167.054
R17662 a_n11689_9690.n1 a_n11689_9690.n6 147.466
R17663 a_n11689_9690.n0 a_n11689_9690.n5 147.466
R17664 a_n11689_9690.n8 a_n11689_9690.t7 31.2553
R17665 a_n11689_9690.n8 a_n11689_9690.t6 31.2553
R17666 a_n11689_9690.n6 a_n11689_9690.t0 31.2553
R17667 a_n11689_9690.n6 a_n11689_9690.t13 31.2553
R17668 a_n11689_9690.n5 a_n11689_9690.t12 31.2553
R17669 a_n11689_9690.n5 a_n11689_9690.t2 31.2553
R17670 a_n11689_9690.n3 a_n11689_9690.t9 31.2553
R17671 a_n11689_9690.n3 a_n11689_9690.t10 31.2553
R17672 a_n11689_9690.n2 a_n11689_9690.t5 31.2553
R17673 a_n11689_9690.n2 a_n11689_9690.t4 31.2553
R17674 a_n11689_9690.t11 a_n11689_9690.n10 31.2553
R17675 a_n11689_9690.n10 a_n11689_9690.t8 31.2553
R17676 a_n11689_9690.n7 a_n11689_9690.n4 18.1752
R17677 a_n11689_9690.n9 a_n11689_9690.n7 13.3361
R17678 a_n11689_9690.n1 a_n11689_9690.n0 5.98829
R17679 a_n11689_9690.n7 a_n11689_9690.n1 5.8324
R17680 VDD.n117 VDD.n80 452.195
R17681 VDD.n3661 VDD.n82 452.195
R17682 VDD.n276 VDD.n255 452.195
R17683 VDD.n3520 VDD.n257 452.195
R17684 VDD.n1632 VDD.n1631 452.195
R17685 VDD.n1673 VDD.n1182 452.195
R17686 VDD.n1358 VDD.n1339 452.195
R17687 VDD.n1442 VDD.n1341 452.195
R17688 VDD.t68 VDD.t98 310.212
R17689 VDD.t86 VDD.t0 310.212
R17690 VDD.n3013 VDD.n709 307.317
R17691 VDD.n3438 VDD.n326 307.317
R17692 VDD.n3411 VDD.n3410 307.317
R17693 VDD.n2781 VDD.n2559 307.317
R17694 VDD.n2545 VDD.n735 307.317
R17695 VDD.n2515 VDD.n2514 307.317
R17696 VDD.n1712 VDD.n1109 307.317
R17697 VDD.n2105 VDD.n1107 307.317
R17698 VDD.n3388 VDD.n3387 307.317
R17699 VDD.n3448 VDD.n318 307.317
R17700 VDD.n2978 VDD.n2782 307.317
R17701 VDD.n3011 VDD.n2783 307.317
R17702 VDD.n2493 VDD.n2492 307.317
R17703 VDD.n2555 VDD.n727 307.317
R17704 VDD.n2069 VDD.n1110 307.317
R17705 VDD.n2103 VDD.n1111 307.317
R17706 VDD.n1671 VDD.t68 300.135
R17707 VDD.n3518 VDD.t0 300.135
R17708 VDD.n2790 VDD.t35 282.913
R17709 VDD.n335 VDD.t22 282.913
R17710 VDD.n2588 VDD.t48 282.913
R17711 VDD.n314 VDD.t41 282.913
R17712 VDD.n1119 VDD.t67 282.913
R17713 VDD.n1137 VDD.t27 282.913
R17714 VDD.n737 VDD.t60 282.913
R17715 VDD.n2462 VDD.t18 282.913
R17716 VDD.t98 VDD.t76 254.097
R17717 VDD.t102 VDD.t86 254.097
R17718 VDD.n1396 VDD.t36 231.792
R17719 VDD.n1420 VDD.t53 231.792
R17720 VDD.n290 VDD.t62 231.792
R17721 VDD.n305 VDD.t49 231.792
R17722 VDD.n97 VDD.t56 231.792
R17723 VDD.n107 VDD.t12 231.792
R17724 VDD.n1192 VDD.t43 231.792
R17725 VDD.n1179 VDD.t28 231.792
R17726 VDD.n2790 VDD.t32 210.619
R17727 VDD.n335 VDD.t20 210.619
R17728 VDD.n2588 VDD.t46 210.619
R17729 VDD.n314 VDD.t40 210.619
R17730 VDD.n1119 VDD.t65 210.619
R17731 VDD.n1137 VDD.t24 210.619
R17732 VDD.n737 VDD.t59 210.619
R17733 VDD.n2462 VDD.t16 210.619
R17734 VDD.n1396 VDD.t39 187.812
R17735 VDD.n1420 VDD.t55 187.812
R17736 VDD.n290 VDD.t64 187.812
R17737 VDD.n305 VDD.t52 187.812
R17738 VDD.n97 VDD.t57 187.812
R17739 VDD.n107 VDD.t14 187.812
R17740 VDD.n1192 VDD.t44 187.812
R17741 VDD.n1179 VDD.t30 187.812
R17742 VDD.n2494 VDD.n2493 185
R17743 VDD.n2493 VDD.n710 185
R17744 VDD.n2495 VDD.n733 185
R17745 VDD.n2550 VDD.n733 185
R17746 VDD.n2497 VDD.n2496 185
R17747 VDD.n2496 VDD.n731 185
R17748 VDD.n2498 VDD.n744 185
R17749 VDD.n2508 VDD.n744 185
R17750 VDD.n2499 VDD.n752 185
R17751 VDD.n752 VDD.n742 185
R17752 VDD.n2501 VDD.n2500 185
R17753 VDD.n2502 VDD.n2501 185
R17754 VDD.n2461 VDD.n751 185
R17755 VDD.n751 VDD.n748 185
R17756 VDD.n2460 VDD.n2459 185
R17757 VDD.n2459 VDD.n2458 185
R17758 VDD.n754 VDD.n753 185
R17759 VDD.n755 VDD.n754 185
R17760 VDD.n2451 VDD.n2450 185
R17761 VDD.n2452 VDD.n2451 185
R17762 VDD.n2449 VDD.n764 185
R17763 VDD.n764 VDD.n761 185
R17764 VDD.n2448 VDD.n2447 185
R17765 VDD.n2447 VDD.n2446 185
R17766 VDD.n766 VDD.n765 185
R17767 VDD.n1896 VDD.n766 185
R17768 VDD.n2439 VDD.n2438 185
R17769 VDD.n2440 VDD.n2439 185
R17770 VDD.n2437 VDD.n775 185
R17771 VDD.n775 VDD.n772 185
R17772 VDD.n2436 VDD.n2435 185
R17773 VDD.n2435 VDD.n2434 185
R17774 VDD.n777 VDD.n776 185
R17775 VDD.n778 VDD.n777 185
R17776 VDD.n2427 VDD.n2426 185
R17777 VDD.n2428 VDD.n2427 185
R17778 VDD.n2425 VDD.n787 185
R17779 VDD.n787 VDD.n784 185
R17780 VDD.n2424 VDD.n2423 185
R17781 VDD.n2423 VDD.n2422 185
R17782 VDD.n789 VDD.n788 185
R17783 VDD.n790 VDD.n789 185
R17784 VDD.n2415 VDD.n2414 185
R17785 VDD.n2416 VDD.n2415 185
R17786 VDD.n2413 VDD.n799 185
R17787 VDD.n799 VDD.n796 185
R17788 VDD.n2412 VDD.n2411 185
R17789 VDD.n2411 VDD.n2410 185
R17790 VDD.n801 VDD.n800 185
R17791 VDD.n802 VDD.n801 185
R17792 VDD.n2403 VDD.n2402 185
R17793 VDD.n2404 VDD.n2403 185
R17794 VDD.n2401 VDD.n811 185
R17795 VDD.n811 VDD.n808 185
R17796 VDD.n2400 VDD.n2399 185
R17797 VDD.n2399 VDD.n2398 185
R17798 VDD.n813 VDD.n812 185
R17799 VDD.n814 VDD.n813 185
R17800 VDD.n2391 VDD.n2390 185
R17801 VDD.n2392 VDD.n2391 185
R17802 VDD.n2389 VDD.n823 185
R17803 VDD.n823 VDD.n820 185
R17804 VDD.n2388 VDD.n2387 185
R17805 VDD.n2387 VDD.n2386 185
R17806 VDD.n825 VDD.n824 185
R17807 VDD.n834 VDD.n825 185
R17808 VDD.n2379 VDD.n2378 185
R17809 VDD.n2380 VDD.n2379 185
R17810 VDD.n2377 VDD.n835 185
R17811 VDD.n835 VDD.n831 185
R17812 VDD.n2376 VDD.n2375 185
R17813 VDD.n2375 VDD.n2374 185
R17814 VDD.n837 VDD.n836 185
R17815 VDD.n838 VDD.n837 185
R17816 VDD.n2367 VDD.n2366 185
R17817 VDD.n2368 VDD.n2367 185
R17818 VDD.n2365 VDD.n847 185
R17819 VDD.n847 VDD.n844 185
R17820 VDD.n2364 VDD.n2363 185
R17821 VDD.n2363 VDD.n2362 185
R17822 VDD.n849 VDD.n848 185
R17823 VDD.n850 VDD.n849 185
R17824 VDD.n2355 VDD.n2354 185
R17825 VDD.n2356 VDD.n2355 185
R17826 VDD.n2353 VDD.n859 185
R17827 VDD.n859 VDD.n856 185
R17828 VDD.n2352 VDD.n2351 185
R17829 VDD.n2351 VDD.n2350 185
R17830 VDD.n861 VDD.n860 185
R17831 VDD.n862 VDD.n861 185
R17832 VDD.n2343 VDD.n2342 185
R17833 VDD.n2344 VDD.n2343 185
R17834 VDD.n2341 VDD.n871 185
R17835 VDD.n871 VDD.n868 185
R17836 VDD.n2340 VDD.n2339 185
R17837 VDD.n2339 VDD.n2338 185
R17838 VDD.n873 VDD.n872 185
R17839 VDD.n874 VDD.n873 185
R17840 VDD.n2331 VDD.n2330 185
R17841 VDD.n2332 VDD.n2331 185
R17842 VDD.n2329 VDD.n883 185
R17843 VDD.n883 VDD.n880 185
R17844 VDD.n2328 VDD.n2327 185
R17845 VDD.n2327 VDD.n2326 185
R17846 VDD.n885 VDD.n884 185
R17847 VDD.n886 VDD.n885 185
R17848 VDD.n2319 VDD.n2318 185
R17849 VDD.n2320 VDD.n2319 185
R17850 VDD.n2317 VDD.n894 185
R17851 VDD.n900 VDD.n894 185
R17852 VDD.n2316 VDD.n2315 185
R17853 VDD.n2315 VDD.n2314 185
R17854 VDD.n896 VDD.n895 185
R17855 VDD.n897 VDD.n896 185
R17856 VDD.n2307 VDD.n2306 185
R17857 VDD.n2308 VDD.n2307 185
R17858 VDD.n2305 VDD.n907 185
R17859 VDD.n907 VDD.n904 185
R17860 VDD.n2304 VDD.n2303 185
R17861 VDD.n2303 VDD.n2302 185
R17862 VDD.n909 VDD.n908 185
R17863 VDD.n910 VDD.n909 185
R17864 VDD.n2295 VDD.n2294 185
R17865 VDD.n2296 VDD.n2295 185
R17866 VDD.n2293 VDD.n919 185
R17867 VDD.n919 VDD.n916 185
R17868 VDD.n2292 VDD.n2291 185
R17869 VDD.n2291 VDD.n2290 185
R17870 VDD.n921 VDD.n920 185
R17871 VDD.n922 VDD.n921 185
R17872 VDD.n2283 VDD.n2282 185
R17873 VDD.n2284 VDD.n2283 185
R17874 VDD.n2281 VDD.n931 185
R17875 VDD.n931 VDD.n928 185
R17876 VDD.n2280 VDD.n2279 185
R17877 VDD.n2279 VDD.n2278 185
R17878 VDD.n933 VDD.n932 185
R17879 VDD.n934 VDD.n933 185
R17880 VDD.n2271 VDD.n2270 185
R17881 VDD.n2272 VDD.n2271 185
R17882 VDD.n2269 VDD.n942 185
R17883 VDD.n947 VDD.n942 185
R17884 VDD.n2268 VDD.n2267 185
R17885 VDD.n2267 VDD.n2266 185
R17886 VDD.n944 VDD.n943 185
R17887 VDD.n954 VDD.n944 185
R17888 VDD.n2259 VDD.n2258 185
R17889 VDD.n2260 VDD.n2259 185
R17890 VDD.n2257 VDD.n955 185
R17891 VDD.n955 VDD.n951 185
R17892 VDD.n2256 VDD.n2255 185
R17893 VDD.n2255 VDD.n2254 185
R17894 VDD.n957 VDD.n956 185
R17895 VDD.n958 VDD.n957 185
R17896 VDD.n2247 VDD.n2246 185
R17897 VDD.n2248 VDD.n2247 185
R17898 VDD.n2245 VDD.n967 185
R17899 VDD.n967 VDD.n964 185
R17900 VDD.n2244 VDD.n2243 185
R17901 VDD.n2243 VDD.n2242 185
R17902 VDD.n969 VDD.n968 185
R17903 VDD.n970 VDD.n969 185
R17904 VDD.n2235 VDD.n2234 185
R17905 VDD.n2236 VDD.n2235 185
R17906 VDD.n2233 VDD.n979 185
R17907 VDD.n979 VDD.n976 185
R17908 VDD.n2232 VDD.n2231 185
R17909 VDD.n2231 VDD.n2230 185
R17910 VDD.n981 VDD.n980 185
R17911 VDD.n982 VDD.n981 185
R17912 VDD.n2223 VDD.n2222 185
R17913 VDD.n2224 VDD.n2223 185
R17914 VDD.n2221 VDD.n991 185
R17915 VDD.n991 VDD.n988 185
R17916 VDD.n2220 VDD.n2219 185
R17917 VDD.n2219 VDD.n2218 185
R17918 VDD.n993 VDD.n992 185
R17919 VDD.n994 VDD.n993 185
R17920 VDD.n2211 VDD.n2210 185
R17921 VDD.n2212 VDD.n2211 185
R17922 VDD.n2209 VDD.n1003 185
R17923 VDD.n1003 VDD.n1000 185
R17924 VDD.n2208 VDD.n2207 185
R17925 VDD.n2207 VDD.n2206 185
R17926 VDD.n1005 VDD.n1004 185
R17927 VDD.n1006 VDD.n1005 185
R17928 VDD.n2199 VDD.n2198 185
R17929 VDD.n2200 VDD.n2199 185
R17930 VDD.n2197 VDD.n1015 185
R17931 VDD.n1015 VDD.n1012 185
R17932 VDD.n2196 VDD.n2195 185
R17933 VDD.n2195 VDD.n2194 185
R17934 VDD.n1017 VDD.n1016 185
R17935 VDD.n1018 VDD.n1017 185
R17936 VDD.n2187 VDD.n2186 185
R17937 VDD.n2188 VDD.n2187 185
R17938 VDD.n2185 VDD.n1026 185
R17939 VDD.n1032 VDD.n1026 185
R17940 VDD.n2184 VDD.n2183 185
R17941 VDD.n2183 VDD.n2182 185
R17942 VDD.n1028 VDD.n1027 185
R17943 VDD.n1029 VDD.n1028 185
R17944 VDD.n2175 VDD.n2174 185
R17945 VDD.n2176 VDD.n2175 185
R17946 VDD.n2173 VDD.n1039 185
R17947 VDD.n1039 VDD.n1036 185
R17948 VDD.n2172 VDD.n2171 185
R17949 VDD.n2171 VDD.n2170 185
R17950 VDD.n1041 VDD.n1040 185
R17951 VDD.n1042 VDD.n1041 185
R17952 VDD.n2163 VDD.n2162 185
R17953 VDD.n2164 VDD.n2163 185
R17954 VDD.n2161 VDD.n1051 185
R17955 VDD.n1051 VDD.n1048 185
R17956 VDD.n2160 VDD.n2159 185
R17957 VDD.n2159 VDD.n2158 185
R17958 VDD.n1053 VDD.n1052 185
R17959 VDD.n1054 VDD.n1053 185
R17960 VDD.n2151 VDD.n2150 185
R17961 VDD.n2152 VDD.n2151 185
R17962 VDD.n2149 VDD.n1063 185
R17963 VDD.n1063 VDD.n1060 185
R17964 VDD.n2148 VDD.n2147 185
R17965 VDD.n2147 VDD.n2146 185
R17966 VDD.n1065 VDD.n1064 185
R17967 VDD.n1066 VDD.n1065 185
R17968 VDD.n2139 VDD.n2138 185
R17969 VDD.n2140 VDD.n2139 185
R17970 VDD.n2137 VDD.n1074 185
R17971 VDD.n1080 VDD.n1074 185
R17972 VDD.n2136 VDD.n2135 185
R17973 VDD.n2135 VDD.n2134 185
R17974 VDD.n1076 VDD.n1075 185
R17975 VDD.n1077 VDD.n1076 185
R17976 VDD.n2127 VDD.n2126 185
R17977 VDD.n2128 VDD.n2127 185
R17978 VDD.n2125 VDD.n1087 185
R17979 VDD.n1087 VDD.n1084 185
R17980 VDD.n2124 VDD.n2123 185
R17981 VDD.n2123 VDD.n2122 185
R17982 VDD.n1089 VDD.n1088 185
R17983 VDD.n1090 VDD.n1089 185
R17984 VDD.n2115 VDD.n2114 185
R17985 VDD.n2116 VDD.n2115 185
R17986 VDD.n2113 VDD.n1099 185
R17987 VDD.n1099 VDD.n1096 185
R17988 VDD.n2112 VDD.n2111 185
R17989 VDD.n2111 VDD.n2110 185
R17990 VDD.n1101 VDD.n1100 185
R17991 VDD.n1102 VDD.n1101 185
R17992 VDD.n2103 VDD.n2102 185
R17993 VDD.n2104 VDD.n2103 185
R17994 VDD.n2101 VDD.n1111 185
R17995 VDD.n2100 VDD.n2099 185
R17996 VDD.n2097 VDD.n1112 185
R17997 VDD.n2095 VDD.n2094 185
R17998 VDD.n2093 VDD.n1113 185
R17999 VDD.n2092 VDD.n2091 185
R18000 VDD.n2089 VDD.n1114 185
R18001 VDD.n2087 VDD.n2086 185
R18002 VDD.n2084 VDD.n1115 185
R18003 VDD.n2083 VDD.n2082 185
R18004 VDD.n2080 VDD.n1117 185
R18005 VDD.n2078 VDD.n2077 185
R18006 VDD.n2075 VDD.n1118 185
R18007 VDD.n2074 VDD.n2073 185
R18008 VDD.n2071 VDD.n1121 185
R18009 VDD.n2069 VDD.n2068 185
R18010 VDD.n2555 VDD.n2554 185
R18011 VDD.n728 VDD.n726 185
R18012 VDD.n2466 VDD.n2465 185
R18013 VDD.n2468 VDD.n2467 185
R18014 VDD.n2470 VDD.n2469 185
R18015 VDD.n2472 VDD.n2471 185
R18016 VDD.n2474 VDD.n2473 185
R18017 VDD.n2476 VDD.n2475 185
R18018 VDD.n2478 VDD.n2477 185
R18019 VDD.n2480 VDD.n2479 185
R18020 VDD.n2482 VDD.n2481 185
R18021 VDD.n2484 VDD.n2483 185
R18022 VDD.n2486 VDD.n2485 185
R18023 VDD.n2488 VDD.n2487 185
R18024 VDD.n2490 VDD.n2489 185
R18025 VDD.n2492 VDD.n2491 185
R18026 VDD.n2553 VDD.n727 185
R18027 VDD.n727 VDD.n710 185
R18028 VDD.n2552 VDD.n2551 185
R18029 VDD.n2551 VDD.n2550 185
R18030 VDD.n730 VDD.n729 185
R18031 VDD.n731 VDD.n730 185
R18032 VDD.n1122 VDD.n743 185
R18033 VDD.n2508 VDD.n743 185
R18034 VDD.n1124 VDD.n1123 185
R18035 VDD.n1123 VDD.n742 185
R18036 VDD.n1125 VDD.n750 185
R18037 VDD.n2502 VDD.n750 185
R18038 VDD.n1127 VDD.n1126 185
R18039 VDD.n1126 VDD.n748 185
R18040 VDD.n1128 VDD.n757 185
R18041 VDD.n2458 VDD.n757 185
R18042 VDD.n1130 VDD.n1129 185
R18043 VDD.n1129 VDD.n755 185
R18044 VDD.n1131 VDD.n763 185
R18045 VDD.n2452 VDD.n763 185
R18046 VDD.n1133 VDD.n1132 185
R18047 VDD.n1132 VDD.n761 185
R18048 VDD.n1134 VDD.n768 185
R18049 VDD.n2446 VDD.n768 185
R18050 VDD.n1898 VDD.n1897 185
R18051 VDD.n1897 VDD.n1896 185
R18052 VDD.n1899 VDD.n774 185
R18053 VDD.n2440 VDD.n774 185
R18054 VDD.n1901 VDD.n1900 185
R18055 VDD.n1900 VDD.n772 185
R18056 VDD.n1902 VDD.n780 185
R18057 VDD.n2434 VDD.n780 185
R18058 VDD.n1904 VDD.n1903 185
R18059 VDD.n1903 VDD.n778 185
R18060 VDD.n1905 VDD.n786 185
R18061 VDD.n2428 VDD.n786 185
R18062 VDD.n1907 VDD.n1906 185
R18063 VDD.n1906 VDD.n784 185
R18064 VDD.n1908 VDD.n792 185
R18065 VDD.n2422 VDD.n792 185
R18066 VDD.n1910 VDD.n1909 185
R18067 VDD.n1909 VDD.n790 185
R18068 VDD.n1911 VDD.n798 185
R18069 VDD.n2416 VDD.n798 185
R18070 VDD.n1913 VDD.n1912 185
R18071 VDD.n1912 VDD.n796 185
R18072 VDD.n1914 VDD.n804 185
R18073 VDD.n2410 VDD.n804 185
R18074 VDD.n1916 VDD.n1915 185
R18075 VDD.n1915 VDD.n802 185
R18076 VDD.n1917 VDD.n810 185
R18077 VDD.n2404 VDD.n810 185
R18078 VDD.n1919 VDD.n1918 185
R18079 VDD.n1918 VDD.n808 185
R18080 VDD.n1920 VDD.n816 185
R18081 VDD.n2398 VDD.n816 185
R18082 VDD.n1922 VDD.n1921 185
R18083 VDD.n1921 VDD.n814 185
R18084 VDD.n1923 VDD.n822 185
R18085 VDD.n2392 VDD.n822 185
R18086 VDD.n1925 VDD.n1924 185
R18087 VDD.n1924 VDD.n820 185
R18088 VDD.n1926 VDD.n827 185
R18089 VDD.n2386 VDD.n827 185
R18090 VDD.n1928 VDD.n1927 185
R18091 VDD.n1927 VDD.n834 185
R18092 VDD.n1929 VDD.n833 185
R18093 VDD.n2380 VDD.n833 185
R18094 VDD.n1931 VDD.n1930 185
R18095 VDD.n1930 VDD.n831 185
R18096 VDD.n1932 VDD.n840 185
R18097 VDD.n2374 VDD.n840 185
R18098 VDD.n1934 VDD.n1933 185
R18099 VDD.n1933 VDD.n838 185
R18100 VDD.n1935 VDD.n846 185
R18101 VDD.n2368 VDD.n846 185
R18102 VDD.n1937 VDD.n1936 185
R18103 VDD.n1936 VDD.n844 185
R18104 VDD.n1938 VDD.n852 185
R18105 VDD.n2362 VDD.n852 185
R18106 VDD.n1940 VDD.n1939 185
R18107 VDD.n1939 VDD.n850 185
R18108 VDD.n1941 VDD.n858 185
R18109 VDD.n2356 VDD.n858 185
R18110 VDD.n1943 VDD.n1942 185
R18111 VDD.n1942 VDD.n856 185
R18112 VDD.n1944 VDD.n864 185
R18113 VDD.n2350 VDD.n864 185
R18114 VDD.n1946 VDD.n1945 185
R18115 VDD.n1945 VDD.n862 185
R18116 VDD.n1947 VDD.n870 185
R18117 VDD.n2344 VDD.n870 185
R18118 VDD.n1949 VDD.n1948 185
R18119 VDD.n1948 VDD.n868 185
R18120 VDD.n1950 VDD.n876 185
R18121 VDD.n2338 VDD.n876 185
R18122 VDD.n1952 VDD.n1951 185
R18123 VDD.n1951 VDD.n874 185
R18124 VDD.n1953 VDD.n882 185
R18125 VDD.n2332 VDD.n882 185
R18126 VDD.n1955 VDD.n1954 185
R18127 VDD.n1954 VDD.n880 185
R18128 VDD.n1956 VDD.n888 185
R18129 VDD.n2326 VDD.n888 185
R18130 VDD.n1958 VDD.n1957 185
R18131 VDD.n1957 VDD.n886 185
R18132 VDD.n1959 VDD.n893 185
R18133 VDD.n2320 VDD.n893 185
R18134 VDD.n1961 VDD.n1960 185
R18135 VDD.n1960 VDD.n900 185
R18136 VDD.n1962 VDD.n899 185
R18137 VDD.n2314 VDD.n899 185
R18138 VDD.n1964 VDD.n1963 185
R18139 VDD.n1963 VDD.n897 185
R18140 VDD.n1965 VDD.n906 185
R18141 VDD.n2308 VDD.n906 185
R18142 VDD.n1967 VDD.n1966 185
R18143 VDD.n1966 VDD.n904 185
R18144 VDD.n1968 VDD.n912 185
R18145 VDD.n2302 VDD.n912 185
R18146 VDD.n1970 VDD.n1969 185
R18147 VDD.n1969 VDD.n910 185
R18148 VDD.n1971 VDD.n918 185
R18149 VDD.n2296 VDD.n918 185
R18150 VDD.n1973 VDD.n1972 185
R18151 VDD.n1972 VDD.n916 185
R18152 VDD.n1974 VDD.n924 185
R18153 VDD.n2290 VDD.n924 185
R18154 VDD.n1976 VDD.n1975 185
R18155 VDD.n1975 VDD.n922 185
R18156 VDD.n1977 VDD.n930 185
R18157 VDD.n2284 VDD.n930 185
R18158 VDD.n1979 VDD.n1978 185
R18159 VDD.n1978 VDD.n928 185
R18160 VDD.n1980 VDD.n936 185
R18161 VDD.n2278 VDD.n936 185
R18162 VDD.n1982 VDD.n1981 185
R18163 VDD.n1981 VDD.n934 185
R18164 VDD.n1983 VDD.n941 185
R18165 VDD.n2272 VDD.n941 185
R18166 VDD.n1985 VDD.n1984 185
R18167 VDD.n1984 VDD.n947 185
R18168 VDD.n1986 VDD.n946 185
R18169 VDD.n2266 VDD.n946 185
R18170 VDD.n1988 VDD.n1987 185
R18171 VDD.n1987 VDD.n954 185
R18172 VDD.n1989 VDD.n953 185
R18173 VDD.n2260 VDD.n953 185
R18174 VDD.n1991 VDD.n1990 185
R18175 VDD.n1990 VDD.n951 185
R18176 VDD.n1992 VDD.n960 185
R18177 VDD.n2254 VDD.n960 185
R18178 VDD.n1994 VDD.n1993 185
R18179 VDD.n1993 VDD.n958 185
R18180 VDD.n1995 VDD.n966 185
R18181 VDD.n2248 VDD.n966 185
R18182 VDD.n1997 VDD.n1996 185
R18183 VDD.n1996 VDD.n964 185
R18184 VDD.n1998 VDD.n972 185
R18185 VDD.n2242 VDD.n972 185
R18186 VDD.n2000 VDD.n1999 185
R18187 VDD.n1999 VDD.n970 185
R18188 VDD.n2001 VDD.n978 185
R18189 VDD.n2236 VDD.n978 185
R18190 VDD.n2003 VDD.n2002 185
R18191 VDD.n2002 VDD.n976 185
R18192 VDD.n2004 VDD.n984 185
R18193 VDD.n2230 VDD.n984 185
R18194 VDD.n2006 VDD.n2005 185
R18195 VDD.n2005 VDD.n982 185
R18196 VDD.n2007 VDD.n990 185
R18197 VDD.n2224 VDD.n990 185
R18198 VDD.n2009 VDD.n2008 185
R18199 VDD.n2008 VDD.n988 185
R18200 VDD.n2010 VDD.n996 185
R18201 VDD.n2218 VDD.n996 185
R18202 VDD.n2012 VDD.n2011 185
R18203 VDD.n2011 VDD.n994 185
R18204 VDD.n2013 VDD.n1002 185
R18205 VDD.n2212 VDD.n1002 185
R18206 VDD.n2015 VDD.n2014 185
R18207 VDD.n2014 VDD.n1000 185
R18208 VDD.n2016 VDD.n1008 185
R18209 VDD.n2206 VDD.n1008 185
R18210 VDD.n2018 VDD.n2017 185
R18211 VDD.n2017 VDD.n1006 185
R18212 VDD.n2019 VDD.n1014 185
R18213 VDD.n2200 VDD.n1014 185
R18214 VDD.n2021 VDD.n2020 185
R18215 VDD.n2020 VDD.n1012 185
R18216 VDD.n2022 VDD.n1020 185
R18217 VDD.n2194 VDD.n1020 185
R18218 VDD.n2024 VDD.n2023 185
R18219 VDD.n2023 VDD.n1018 185
R18220 VDD.n2025 VDD.n1025 185
R18221 VDD.n2188 VDD.n1025 185
R18222 VDD.n2027 VDD.n2026 185
R18223 VDD.n2026 VDD.n1032 185
R18224 VDD.n2028 VDD.n1031 185
R18225 VDD.n2182 VDD.n1031 185
R18226 VDD.n2030 VDD.n2029 185
R18227 VDD.n2029 VDD.n1029 185
R18228 VDD.n2031 VDD.n1038 185
R18229 VDD.n2176 VDD.n1038 185
R18230 VDD.n2033 VDD.n2032 185
R18231 VDD.n2032 VDD.n1036 185
R18232 VDD.n2034 VDD.n1044 185
R18233 VDD.n2170 VDD.n1044 185
R18234 VDD.n2036 VDD.n2035 185
R18235 VDD.n2035 VDD.n1042 185
R18236 VDD.n2037 VDD.n1050 185
R18237 VDD.n2164 VDD.n1050 185
R18238 VDD.n2039 VDD.n2038 185
R18239 VDD.n2038 VDD.n1048 185
R18240 VDD.n2040 VDD.n1056 185
R18241 VDD.n2158 VDD.n1056 185
R18242 VDD.n2042 VDD.n2041 185
R18243 VDD.n2041 VDD.n1054 185
R18244 VDD.n2043 VDD.n1062 185
R18245 VDD.n2152 VDD.n1062 185
R18246 VDD.n2045 VDD.n2044 185
R18247 VDD.n2044 VDD.n1060 185
R18248 VDD.n2046 VDD.n1068 185
R18249 VDD.n2146 VDD.n1068 185
R18250 VDD.n2048 VDD.n2047 185
R18251 VDD.n2047 VDD.n1066 185
R18252 VDD.n2049 VDD.n1073 185
R18253 VDD.n2140 VDD.n1073 185
R18254 VDD.n2051 VDD.n2050 185
R18255 VDD.n2050 VDD.n1080 185
R18256 VDD.n2052 VDD.n1079 185
R18257 VDD.n2134 VDD.n1079 185
R18258 VDD.n2054 VDD.n2053 185
R18259 VDD.n2053 VDD.n1077 185
R18260 VDD.n2055 VDD.n1086 185
R18261 VDD.n2128 VDD.n1086 185
R18262 VDD.n2057 VDD.n2056 185
R18263 VDD.n2056 VDD.n1084 185
R18264 VDD.n2058 VDD.n1092 185
R18265 VDD.n2122 VDD.n1092 185
R18266 VDD.n2060 VDD.n2059 185
R18267 VDD.n2059 VDD.n1090 185
R18268 VDD.n2061 VDD.n1098 185
R18269 VDD.n2116 VDD.n1098 185
R18270 VDD.n2063 VDD.n2062 185
R18271 VDD.n2062 VDD.n1096 185
R18272 VDD.n2064 VDD.n1104 185
R18273 VDD.n2110 VDD.n1104 185
R18274 VDD.n2066 VDD.n2065 185
R18275 VDD.n2065 VDD.n1102 185
R18276 VDD.n2067 VDD.n1110 185
R18277 VDD.n2104 VDD.n1110 185
R18278 VDD.n3389 VDD.n3388 185
R18279 VDD.n3388 VDD.n323 185
R18280 VDD.n3390 VDD.n324 185
R18281 VDD.n3443 VDD.n324 185
R18282 VDD.n3392 VDD.n3391 185
R18283 VDD.n3391 VDD.n321 185
R18284 VDD.n3393 VDD.n345 185
R18285 VDD.n3403 VDD.n345 185
R18286 VDD.n3394 VDD.n353 185
R18287 VDD.n353 VDD.n343 185
R18288 VDD.n3396 VDD.n3395 185
R18289 VDD.n3397 VDD.n3396 185
R18290 VDD.n3369 VDD.n352 185
R18291 VDD.n352 VDD.n349 185
R18292 VDD.n3368 VDD.n3367 185
R18293 VDD.n3367 VDD.n3366 185
R18294 VDD.n355 VDD.n354 185
R18295 VDD.n356 VDD.n355 185
R18296 VDD.n3359 VDD.n3358 185
R18297 VDD.n3360 VDD.n3359 185
R18298 VDD.n3357 VDD.n365 185
R18299 VDD.n365 VDD.n362 185
R18300 VDD.n3356 VDD.n3355 185
R18301 VDD.n3355 VDD.n3354 185
R18302 VDD.n367 VDD.n366 185
R18303 VDD.n376 VDD.n367 185
R18304 VDD.n3347 VDD.n3346 185
R18305 VDD.n3348 VDD.n3347 185
R18306 VDD.n3345 VDD.n377 185
R18307 VDD.n377 VDD.n373 185
R18308 VDD.n3344 VDD.n3343 185
R18309 VDD.n3343 VDD.n3342 185
R18310 VDD.n379 VDD.n378 185
R18311 VDD.n380 VDD.n379 185
R18312 VDD.n3335 VDD.n3334 185
R18313 VDD.n3336 VDD.n3335 185
R18314 VDD.n3333 VDD.n389 185
R18315 VDD.n389 VDD.n386 185
R18316 VDD.n3332 VDD.n3331 185
R18317 VDD.n3331 VDD.n3330 185
R18318 VDD.n391 VDD.n390 185
R18319 VDD.n392 VDD.n391 185
R18320 VDD.n3323 VDD.n3322 185
R18321 VDD.n3324 VDD.n3323 185
R18322 VDD.n3321 VDD.n401 185
R18323 VDD.n401 VDD.n398 185
R18324 VDD.n3320 VDD.n3319 185
R18325 VDD.n3319 VDD.n3318 185
R18326 VDD.n403 VDD.n402 185
R18327 VDD.n404 VDD.n403 185
R18328 VDD.n3311 VDD.n3310 185
R18329 VDD.n3312 VDD.n3311 185
R18330 VDD.n3309 VDD.n413 185
R18331 VDD.n413 VDD.n410 185
R18332 VDD.n3308 VDD.n3307 185
R18333 VDD.n3307 VDD.n3306 185
R18334 VDD.n415 VDD.n414 185
R18335 VDD.n424 VDD.n415 185
R18336 VDD.n3299 VDD.n3298 185
R18337 VDD.n3300 VDD.n3299 185
R18338 VDD.n3297 VDD.n425 185
R18339 VDD.n425 VDD.n421 185
R18340 VDD.n3296 VDD.n3295 185
R18341 VDD.n3295 VDD.n3294 185
R18342 VDD.n427 VDD.n426 185
R18343 VDD.n428 VDD.n427 185
R18344 VDD.n3287 VDD.n3286 185
R18345 VDD.n3288 VDD.n3287 185
R18346 VDD.n3285 VDD.n437 185
R18347 VDD.n437 VDD.n434 185
R18348 VDD.n3284 VDD.n3283 185
R18349 VDD.n3283 VDD.n3282 185
R18350 VDD.n439 VDD.n438 185
R18351 VDD.n440 VDD.n439 185
R18352 VDD.n3275 VDD.n3274 185
R18353 VDD.n3276 VDD.n3275 185
R18354 VDD.n3273 VDD.n449 185
R18355 VDD.n449 VDD.n446 185
R18356 VDD.n3272 VDD.n3271 185
R18357 VDD.n3271 VDD.n3270 185
R18358 VDD.n451 VDD.n450 185
R18359 VDD.n452 VDD.n451 185
R18360 VDD.n3263 VDD.n3262 185
R18361 VDD.n3264 VDD.n3263 185
R18362 VDD.n3261 VDD.n461 185
R18363 VDD.n461 VDD.n458 185
R18364 VDD.n3260 VDD.n3259 185
R18365 VDD.n3259 VDD.n3258 185
R18366 VDD.n463 VDD.n462 185
R18367 VDD.n464 VDD.n463 185
R18368 VDD.n3251 VDD.n3250 185
R18369 VDD.n3252 VDD.n3251 185
R18370 VDD.n3249 VDD.n473 185
R18371 VDD.n473 VDD.n470 185
R18372 VDD.n3248 VDD.n3247 185
R18373 VDD.n3247 VDD.n3246 185
R18374 VDD.n475 VDD.n474 185
R18375 VDD.n476 VDD.n475 185
R18376 VDD.n3239 VDD.n3238 185
R18377 VDD.n3240 VDD.n3239 185
R18378 VDD.n3237 VDD.n485 185
R18379 VDD.n485 VDD.n482 185
R18380 VDD.n3236 VDD.n3235 185
R18381 VDD.n3235 VDD.n3234 185
R18382 VDD.n487 VDD.n486 185
R18383 VDD.n488 VDD.n487 185
R18384 VDD.n3227 VDD.n3226 185
R18385 VDD.n3228 VDD.n3227 185
R18386 VDD.n3225 VDD.n496 185
R18387 VDD.n501 VDD.n496 185
R18388 VDD.n3224 VDD.n3223 185
R18389 VDD.n3223 VDD.n3222 185
R18390 VDD.n498 VDD.n497 185
R18391 VDD.n508 VDD.n498 185
R18392 VDD.n3215 VDD.n3214 185
R18393 VDD.n3216 VDD.n3215 185
R18394 VDD.n3213 VDD.n509 185
R18395 VDD.n509 VDD.n505 185
R18396 VDD.n3212 VDD.n3211 185
R18397 VDD.n3211 VDD.n3210 185
R18398 VDD.n511 VDD.n510 185
R18399 VDD.n512 VDD.n511 185
R18400 VDD.n3203 VDD.n3202 185
R18401 VDD.n3204 VDD.n3203 185
R18402 VDD.n3201 VDD.n521 185
R18403 VDD.n521 VDD.n518 185
R18404 VDD.n3200 VDD.n3199 185
R18405 VDD.n3199 VDD.n3198 185
R18406 VDD.n523 VDD.n522 185
R18407 VDD.n524 VDD.n523 185
R18408 VDD.n3191 VDD.n3190 185
R18409 VDD.n3192 VDD.n3191 185
R18410 VDD.n3189 VDD.n533 185
R18411 VDD.n533 VDD.n530 185
R18412 VDD.n3188 VDD.n3187 185
R18413 VDD.n3187 VDD.n3186 185
R18414 VDD.n535 VDD.n534 185
R18415 VDD.n536 VDD.n535 185
R18416 VDD.n3179 VDD.n3178 185
R18417 VDD.n3180 VDD.n3179 185
R18418 VDD.n3177 VDD.n545 185
R18419 VDD.n545 VDD.n542 185
R18420 VDD.n3176 VDD.n3175 185
R18421 VDD.n3175 VDD.n3174 185
R18422 VDD.n547 VDD.n546 185
R18423 VDD.n556 VDD.n547 185
R18424 VDD.n3167 VDD.n3166 185
R18425 VDD.n3168 VDD.n3167 185
R18426 VDD.n3165 VDD.n557 185
R18427 VDD.n557 VDD.n553 185
R18428 VDD.n3164 VDD.n3163 185
R18429 VDD.n3163 VDD.n3162 185
R18430 VDD.n559 VDD.n558 185
R18431 VDD.n560 VDD.n559 185
R18432 VDD.n3155 VDD.n3154 185
R18433 VDD.n3156 VDD.n3155 185
R18434 VDD.n3153 VDD.n569 185
R18435 VDD.n569 VDD.n566 185
R18436 VDD.n3152 VDD.n3151 185
R18437 VDD.n3151 VDD.n3150 185
R18438 VDD.n571 VDD.n570 185
R18439 VDD.n572 VDD.n571 185
R18440 VDD.n3143 VDD.n3142 185
R18441 VDD.n3144 VDD.n3143 185
R18442 VDD.n3141 VDD.n581 185
R18443 VDD.n581 VDD.n578 185
R18444 VDD.n3140 VDD.n3139 185
R18445 VDD.n3139 VDD.n3138 185
R18446 VDD.n583 VDD.n582 185
R18447 VDD.n584 VDD.n583 185
R18448 VDD.n3131 VDD.n3130 185
R18449 VDD.n3132 VDD.n3131 185
R18450 VDD.n3129 VDD.n593 185
R18451 VDD.n593 VDD.n590 185
R18452 VDD.n3128 VDD.n3127 185
R18453 VDD.n3127 VDD.n3126 185
R18454 VDD.n595 VDD.n594 185
R18455 VDD.n596 VDD.n595 185
R18456 VDD.n3119 VDD.n3118 185
R18457 VDD.n3120 VDD.n3119 185
R18458 VDD.n3117 VDD.n605 185
R18459 VDD.n605 VDD.n602 185
R18460 VDD.n3116 VDD.n3115 185
R18461 VDD.n3115 VDD.n3114 185
R18462 VDD.n607 VDD.n606 185
R18463 VDD.n608 VDD.n607 185
R18464 VDD.n3107 VDD.n3106 185
R18465 VDD.n3108 VDD.n3107 185
R18466 VDD.n3105 VDD.n616 185
R18467 VDD.n622 VDD.n616 185
R18468 VDD.n3104 VDD.n3103 185
R18469 VDD.n3103 VDD.n3102 185
R18470 VDD.n618 VDD.n617 185
R18471 VDD.n619 VDD.n618 185
R18472 VDD.n3095 VDD.n3094 185
R18473 VDD.n3096 VDD.n3095 185
R18474 VDD.n3093 VDD.n629 185
R18475 VDD.n629 VDD.n626 185
R18476 VDD.n3092 VDD.n3091 185
R18477 VDD.n3091 VDD.n3090 185
R18478 VDD.n631 VDD.n630 185
R18479 VDD.n632 VDD.n631 185
R18480 VDD.n3083 VDD.n3082 185
R18481 VDD.n3084 VDD.n3083 185
R18482 VDD.n3081 VDD.n641 185
R18483 VDD.n641 VDD.n638 185
R18484 VDD.n3080 VDD.n3079 185
R18485 VDD.n3079 VDD.n3078 185
R18486 VDD.n643 VDD.n642 185
R18487 VDD.n644 VDD.n643 185
R18488 VDD.n3071 VDD.n3070 185
R18489 VDD.n3072 VDD.n3071 185
R18490 VDD.n3069 VDD.n653 185
R18491 VDD.n653 VDD.n650 185
R18492 VDD.n3068 VDD.n3067 185
R18493 VDD.n3067 VDD.n3066 185
R18494 VDD.n655 VDD.n654 185
R18495 VDD.n656 VDD.n655 185
R18496 VDD.n3059 VDD.n3058 185
R18497 VDD.n3060 VDD.n3059 185
R18498 VDD.n3057 VDD.n665 185
R18499 VDD.n665 VDD.n662 185
R18500 VDD.n3056 VDD.n3055 185
R18501 VDD.n3055 VDD.n3054 185
R18502 VDD.n667 VDD.n666 185
R18503 VDD.n668 VDD.n667 185
R18504 VDD.n3047 VDD.n3046 185
R18505 VDD.n3048 VDD.n3047 185
R18506 VDD.n3045 VDD.n676 185
R18507 VDD.n682 VDD.n676 185
R18508 VDD.n3044 VDD.n3043 185
R18509 VDD.n3043 VDD.n3042 185
R18510 VDD.n678 VDD.n677 185
R18511 VDD.n679 VDD.n678 185
R18512 VDD.n3035 VDD.n3034 185
R18513 VDD.n3036 VDD.n3035 185
R18514 VDD.n3033 VDD.n689 185
R18515 VDD.n689 VDD.n686 185
R18516 VDD.n3032 VDD.n3031 185
R18517 VDD.n3031 VDD.n3030 185
R18518 VDD.n691 VDD.n690 185
R18519 VDD.n692 VDD.n691 185
R18520 VDD.n3023 VDD.n3022 185
R18521 VDD.n3024 VDD.n3023 185
R18522 VDD.n3021 VDD.n701 185
R18523 VDD.n701 VDD.n698 185
R18524 VDD.n3020 VDD.n3019 185
R18525 VDD.n3019 VDD.n3018 185
R18526 VDD.n703 VDD.n702 185
R18527 VDD.n704 VDD.n703 185
R18528 VDD.n3011 VDD.n3010 185
R18529 VDD.n3012 VDD.n3011 185
R18530 VDD.n3009 VDD.n2783 185
R18531 VDD.n3008 VDD.n3007 185
R18532 VDD.n3005 VDD.n2784 185
R18533 VDD.n3003 VDD.n3002 185
R18534 VDD.n3001 VDD.n2785 185
R18535 VDD.n3000 VDD.n2999 185
R18536 VDD.n2997 VDD.n2786 185
R18537 VDD.n2995 VDD.n2994 185
R18538 VDD.n2993 VDD.n2787 185
R18539 VDD.n2992 VDD.n2991 185
R18540 VDD.n2989 VDD.n2788 185
R18541 VDD.n2987 VDD.n2986 185
R18542 VDD.n2984 VDD.n2789 185
R18543 VDD.n2983 VDD.n2982 185
R18544 VDD.n2980 VDD.n2792 185
R18545 VDD.n2978 VDD.n2977 185
R18546 VDD.n3448 VDD.n3447 185
R18547 VDD.n3450 VDD.n316 185
R18548 VDD.n3452 VDD.n3451 185
R18549 VDD.n3453 VDD.n313 185
R18550 VDD.n3456 VDD.n3455 185
R18551 VDD.n3458 VDD.n312 185
R18552 VDD.n3459 VDD.n309 185
R18553 VDD.n3462 VDD.n3461 185
R18554 VDD.n310 VDD.n308 185
R18555 VDD.n3376 VDD.n3375 185
R18556 VDD.n3378 VDD.n3377 185
R18557 VDD.n3380 VDD.n3372 185
R18558 VDD.n3382 VDD.n3381 185
R18559 VDD.n3383 VDD.n3371 185
R18560 VDD.n3385 VDD.n3384 185
R18561 VDD.n3387 VDD.n3370 185
R18562 VDD.n3446 VDD.n318 185
R18563 VDD.n323 VDD.n318 185
R18564 VDD.n3445 VDD.n3444 185
R18565 VDD.n3444 VDD.n3443 185
R18566 VDD.n320 VDD.n319 185
R18567 VDD.n321 VDD.n320 185
R18568 VDD.n2793 VDD.n344 185
R18569 VDD.n3403 VDD.n344 185
R18570 VDD.n2795 VDD.n2794 185
R18571 VDD.n2794 VDD.n343 185
R18572 VDD.n2796 VDD.n351 185
R18573 VDD.n3397 VDD.n351 185
R18574 VDD.n2798 VDD.n2797 185
R18575 VDD.n2797 VDD.n349 185
R18576 VDD.n2799 VDD.n358 185
R18577 VDD.n3366 VDD.n358 185
R18578 VDD.n2801 VDD.n2800 185
R18579 VDD.n2800 VDD.n356 185
R18580 VDD.n2802 VDD.n364 185
R18581 VDD.n3360 VDD.n364 185
R18582 VDD.n2804 VDD.n2803 185
R18583 VDD.n2803 VDD.n362 185
R18584 VDD.n2805 VDD.n369 185
R18585 VDD.n3354 VDD.n369 185
R18586 VDD.n2807 VDD.n2806 185
R18587 VDD.n2806 VDD.n376 185
R18588 VDD.n2808 VDD.n375 185
R18589 VDD.n3348 VDD.n375 185
R18590 VDD.n2810 VDD.n2809 185
R18591 VDD.n2809 VDD.n373 185
R18592 VDD.n2811 VDD.n382 185
R18593 VDD.n3342 VDD.n382 185
R18594 VDD.n2813 VDD.n2812 185
R18595 VDD.n2812 VDD.n380 185
R18596 VDD.n2814 VDD.n388 185
R18597 VDD.n3336 VDD.n388 185
R18598 VDD.n2816 VDD.n2815 185
R18599 VDD.n2815 VDD.n386 185
R18600 VDD.n2817 VDD.n394 185
R18601 VDD.n3330 VDD.n394 185
R18602 VDD.n2819 VDD.n2818 185
R18603 VDD.n2818 VDD.n392 185
R18604 VDD.n2820 VDD.n400 185
R18605 VDD.n3324 VDD.n400 185
R18606 VDD.n2822 VDD.n2821 185
R18607 VDD.n2821 VDD.n398 185
R18608 VDD.n2823 VDD.n406 185
R18609 VDD.n3318 VDD.n406 185
R18610 VDD.n2825 VDD.n2824 185
R18611 VDD.n2824 VDD.n404 185
R18612 VDD.n2826 VDD.n412 185
R18613 VDD.n3312 VDD.n412 185
R18614 VDD.n2828 VDD.n2827 185
R18615 VDD.n2827 VDD.n410 185
R18616 VDD.n2829 VDD.n417 185
R18617 VDD.n3306 VDD.n417 185
R18618 VDD.n2831 VDD.n2830 185
R18619 VDD.n2830 VDD.n424 185
R18620 VDD.n2832 VDD.n423 185
R18621 VDD.n3300 VDD.n423 185
R18622 VDD.n2834 VDD.n2833 185
R18623 VDD.n2833 VDD.n421 185
R18624 VDD.n2835 VDD.n430 185
R18625 VDD.n3294 VDD.n430 185
R18626 VDD.n2837 VDD.n2836 185
R18627 VDD.n2836 VDD.n428 185
R18628 VDD.n2838 VDD.n436 185
R18629 VDD.n3288 VDD.n436 185
R18630 VDD.n2840 VDD.n2839 185
R18631 VDD.n2839 VDD.n434 185
R18632 VDD.n2841 VDD.n442 185
R18633 VDD.n3282 VDD.n442 185
R18634 VDD.n2843 VDD.n2842 185
R18635 VDD.n2842 VDD.n440 185
R18636 VDD.n2844 VDD.n448 185
R18637 VDD.n3276 VDD.n448 185
R18638 VDD.n2846 VDD.n2845 185
R18639 VDD.n2845 VDD.n446 185
R18640 VDD.n2847 VDD.n454 185
R18641 VDD.n3270 VDD.n454 185
R18642 VDD.n2849 VDD.n2848 185
R18643 VDD.n2848 VDD.n452 185
R18644 VDD.n2850 VDD.n460 185
R18645 VDD.n3264 VDD.n460 185
R18646 VDD.n2852 VDD.n2851 185
R18647 VDD.n2851 VDD.n458 185
R18648 VDD.n2853 VDD.n466 185
R18649 VDD.n3258 VDD.n466 185
R18650 VDD.n2855 VDD.n2854 185
R18651 VDD.n2854 VDD.n464 185
R18652 VDD.n2856 VDD.n472 185
R18653 VDD.n3252 VDD.n472 185
R18654 VDD.n2858 VDD.n2857 185
R18655 VDD.n2857 VDD.n470 185
R18656 VDD.n2859 VDD.n478 185
R18657 VDD.n3246 VDD.n478 185
R18658 VDD.n2861 VDD.n2860 185
R18659 VDD.n2860 VDD.n476 185
R18660 VDD.n2862 VDD.n484 185
R18661 VDD.n3240 VDD.n484 185
R18662 VDD.n2864 VDD.n2863 185
R18663 VDD.n2863 VDD.n482 185
R18664 VDD.n2865 VDD.n490 185
R18665 VDD.n3234 VDD.n490 185
R18666 VDD.n2867 VDD.n2866 185
R18667 VDD.n2866 VDD.n488 185
R18668 VDD.n2868 VDD.n495 185
R18669 VDD.n3228 VDD.n495 185
R18670 VDD.n2870 VDD.n2869 185
R18671 VDD.n2869 VDD.n501 185
R18672 VDD.n2871 VDD.n500 185
R18673 VDD.n3222 VDD.n500 185
R18674 VDD.n2873 VDD.n2872 185
R18675 VDD.n2872 VDD.n508 185
R18676 VDD.n2874 VDD.n507 185
R18677 VDD.n3216 VDD.n507 185
R18678 VDD.n2876 VDD.n2875 185
R18679 VDD.n2875 VDD.n505 185
R18680 VDD.n2877 VDD.n514 185
R18681 VDD.n3210 VDD.n514 185
R18682 VDD.n2879 VDD.n2878 185
R18683 VDD.n2878 VDD.n512 185
R18684 VDD.n2880 VDD.n520 185
R18685 VDD.n3204 VDD.n520 185
R18686 VDD.n2882 VDD.n2881 185
R18687 VDD.n2881 VDD.n518 185
R18688 VDD.n2883 VDD.n526 185
R18689 VDD.n3198 VDD.n526 185
R18690 VDD.n2885 VDD.n2884 185
R18691 VDD.n2884 VDD.n524 185
R18692 VDD.n2886 VDD.n532 185
R18693 VDD.n3192 VDD.n532 185
R18694 VDD.n2888 VDD.n2887 185
R18695 VDD.n2887 VDD.n530 185
R18696 VDD.n2889 VDD.n538 185
R18697 VDD.n3186 VDD.n538 185
R18698 VDD.n2891 VDD.n2890 185
R18699 VDD.n2890 VDD.n536 185
R18700 VDD.n2892 VDD.n544 185
R18701 VDD.n3180 VDD.n544 185
R18702 VDD.n2894 VDD.n2893 185
R18703 VDD.n2893 VDD.n542 185
R18704 VDD.n2895 VDD.n549 185
R18705 VDD.n3174 VDD.n549 185
R18706 VDD.n2897 VDD.n2896 185
R18707 VDD.n2896 VDD.n556 185
R18708 VDD.n2898 VDD.n555 185
R18709 VDD.n3168 VDD.n555 185
R18710 VDD.n2900 VDD.n2899 185
R18711 VDD.n2899 VDD.n553 185
R18712 VDD.n2901 VDD.n562 185
R18713 VDD.n3162 VDD.n562 185
R18714 VDD.n2903 VDD.n2902 185
R18715 VDD.n2902 VDD.n560 185
R18716 VDD.n2904 VDD.n568 185
R18717 VDD.n3156 VDD.n568 185
R18718 VDD.n2906 VDD.n2905 185
R18719 VDD.n2905 VDD.n566 185
R18720 VDD.n2907 VDD.n574 185
R18721 VDD.n3150 VDD.n574 185
R18722 VDD.n2909 VDD.n2908 185
R18723 VDD.n2908 VDD.n572 185
R18724 VDD.n2910 VDD.n580 185
R18725 VDD.n3144 VDD.n580 185
R18726 VDD.n2912 VDD.n2911 185
R18727 VDD.n2911 VDD.n578 185
R18728 VDD.n2913 VDD.n586 185
R18729 VDD.n3138 VDD.n586 185
R18730 VDD.n2915 VDD.n2914 185
R18731 VDD.n2914 VDD.n584 185
R18732 VDD.n2916 VDD.n592 185
R18733 VDD.n3132 VDD.n592 185
R18734 VDD.n2918 VDD.n2917 185
R18735 VDD.n2917 VDD.n590 185
R18736 VDD.n2919 VDD.n598 185
R18737 VDD.n3126 VDD.n598 185
R18738 VDD.n2921 VDD.n2920 185
R18739 VDD.n2920 VDD.n596 185
R18740 VDD.n2922 VDD.n604 185
R18741 VDD.n3120 VDD.n604 185
R18742 VDD.n2924 VDD.n2923 185
R18743 VDD.n2923 VDD.n602 185
R18744 VDD.n2925 VDD.n610 185
R18745 VDD.n3114 VDD.n610 185
R18746 VDD.n2927 VDD.n2926 185
R18747 VDD.n2926 VDD.n608 185
R18748 VDD.n2928 VDD.n615 185
R18749 VDD.n3108 VDD.n615 185
R18750 VDD.n2930 VDD.n2929 185
R18751 VDD.n2929 VDD.n622 185
R18752 VDD.n2931 VDD.n621 185
R18753 VDD.n3102 VDD.n621 185
R18754 VDD.n2933 VDD.n2932 185
R18755 VDD.n2932 VDD.n619 185
R18756 VDD.n2934 VDD.n628 185
R18757 VDD.n3096 VDD.n628 185
R18758 VDD.n2936 VDD.n2935 185
R18759 VDD.n2935 VDD.n626 185
R18760 VDD.n2937 VDD.n634 185
R18761 VDD.n3090 VDD.n634 185
R18762 VDD.n2939 VDD.n2938 185
R18763 VDD.n2938 VDD.n632 185
R18764 VDD.n2940 VDD.n640 185
R18765 VDD.n3084 VDD.n640 185
R18766 VDD.n2942 VDD.n2941 185
R18767 VDD.n2941 VDD.n638 185
R18768 VDD.n2943 VDD.n646 185
R18769 VDD.n3078 VDD.n646 185
R18770 VDD.n2945 VDD.n2944 185
R18771 VDD.n2944 VDD.n644 185
R18772 VDD.n2946 VDD.n652 185
R18773 VDD.n3072 VDD.n652 185
R18774 VDD.n2948 VDD.n2947 185
R18775 VDD.n2947 VDD.n650 185
R18776 VDD.n2949 VDD.n658 185
R18777 VDD.n3066 VDD.n658 185
R18778 VDD.n2951 VDD.n2950 185
R18779 VDD.n2950 VDD.n656 185
R18780 VDD.n2952 VDD.n664 185
R18781 VDD.n3060 VDD.n664 185
R18782 VDD.n2954 VDD.n2953 185
R18783 VDD.n2953 VDD.n662 185
R18784 VDD.n2955 VDD.n670 185
R18785 VDD.n3054 VDD.n670 185
R18786 VDD.n2957 VDD.n2956 185
R18787 VDD.n2956 VDD.n668 185
R18788 VDD.n2958 VDD.n675 185
R18789 VDD.n3048 VDD.n675 185
R18790 VDD.n2960 VDD.n2959 185
R18791 VDD.n2959 VDD.n682 185
R18792 VDD.n2961 VDD.n681 185
R18793 VDD.n3042 VDD.n681 185
R18794 VDD.n2963 VDD.n2962 185
R18795 VDD.n2962 VDD.n679 185
R18796 VDD.n2964 VDD.n688 185
R18797 VDD.n3036 VDD.n688 185
R18798 VDD.n2966 VDD.n2965 185
R18799 VDD.n2965 VDD.n686 185
R18800 VDD.n2967 VDD.n694 185
R18801 VDD.n3030 VDD.n694 185
R18802 VDD.n2969 VDD.n2968 185
R18803 VDD.n2968 VDD.n692 185
R18804 VDD.n2970 VDD.n700 185
R18805 VDD.n3024 VDD.n700 185
R18806 VDD.n2972 VDD.n2971 185
R18807 VDD.n2971 VDD.n698 185
R18808 VDD.n2973 VDD.n706 185
R18809 VDD.n3018 VDD.n706 185
R18810 VDD.n2975 VDD.n2974 185
R18811 VDD.n2974 VDD.n704 185
R18812 VDD.n2976 VDD.n2782 185
R18813 VDD.n3012 VDD.n2782 185
R18814 VDD.n2547 VDD.n735 185
R18815 VDD.n735 VDD.n710 185
R18816 VDD.n2549 VDD.n2548 185
R18817 VDD.n2550 VDD.n2549 185
R18818 VDD.n736 VDD.n734 185
R18819 VDD.n734 VDD.n731 185
R18820 VDD.n2507 VDD.n2506 185
R18821 VDD.n2508 VDD.n2507 185
R18822 VDD.n2505 VDD.n745 185
R18823 VDD.n745 VDD.n742 185
R18824 VDD.n2504 VDD.n2503 185
R18825 VDD.n2503 VDD.n2502 185
R18826 VDD.n747 VDD.n746 185
R18827 VDD.n748 VDD.n747 185
R18828 VDD.n2457 VDD.n2456 185
R18829 VDD.n2458 VDD.n2457 185
R18830 VDD.n2455 VDD.n758 185
R18831 VDD.n758 VDD.n755 185
R18832 VDD.n2454 VDD.n2453 185
R18833 VDD.n2453 VDD.n2452 185
R18834 VDD.n760 VDD.n759 185
R18835 VDD.n761 VDD.n760 185
R18836 VDD.n2445 VDD.n2444 185
R18837 VDD.n2446 VDD.n2445 185
R18838 VDD.n2443 VDD.n769 185
R18839 VDD.n1896 VDD.n769 185
R18840 VDD.n2442 VDD.n2441 185
R18841 VDD.n2441 VDD.n2440 185
R18842 VDD.n771 VDD.n770 185
R18843 VDD.n772 VDD.n771 185
R18844 VDD.n2433 VDD.n2432 185
R18845 VDD.n2434 VDD.n2433 185
R18846 VDD.n2431 VDD.n781 185
R18847 VDD.n781 VDD.n778 185
R18848 VDD.n2430 VDD.n2429 185
R18849 VDD.n2429 VDD.n2428 185
R18850 VDD.n783 VDD.n782 185
R18851 VDD.n784 VDD.n783 185
R18852 VDD.n2421 VDD.n2420 185
R18853 VDD.n2422 VDD.n2421 185
R18854 VDD.n2419 VDD.n793 185
R18855 VDD.n793 VDD.n790 185
R18856 VDD.n2418 VDD.n2417 185
R18857 VDD.n2417 VDD.n2416 185
R18858 VDD.n795 VDD.n794 185
R18859 VDD.n796 VDD.n795 185
R18860 VDD.n2409 VDD.n2408 185
R18861 VDD.n2410 VDD.n2409 185
R18862 VDD.n2407 VDD.n805 185
R18863 VDD.n805 VDD.n802 185
R18864 VDD.n2406 VDD.n2405 185
R18865 VDD.n2405 VDD.n2404 185
R18866 VDD.n807 VDD.n806 185
R18867 VDD.n808 VDD.n807 185
R18868 VDD.n2397 VDD.n2396 185
R18869 VDD.n2398 VDD.n2397 185
R18870 VDD.n2395 VDD.n817 185
R18871 VDD.n817 VDD.n814 185
R18872 VDD.n2394 VDD.n2393 185
R18873 VDD.n2393 VDD.n2392 185
R18874 VDD.n819 VDD.n818 185
R18875 VDD.n820 VDD.n819 185
R18876 VDD.n2385 VDD.n2384 185
R18877 VDD.n2386 VDD.n2385 185
R18878 VDD.n2383 VDD.n828 185
R18879 VDD.n834 VDD.n828 185
R18880 VDD.n2382 VDD.n2381 185
R18881 VDD.n2381 VDD.n2380 185
R18882 VDD.n830 VDD.n829 185
R18883 VDD.n831 VDD.n830 185
R18884 VDD.n2373 VDD.n2372 185
R18885 VDD.n2374 VDD.n2373 185
R18886 VDD.n2371 VDD.n841 185
R18887 VDD.n841 VDD.n838 185
R18888 VDD.n2370 VDD.n2369 185
R18889 VDD.n2369 VDD.n2368 185
R18890 VDD.n843 VDD.n842 185
R18891 VDD.n844 VDD.n843 185
R18892 VDD.n2361 VDD.n2360 185
R18893 VDD.n2362 VDD.n2361 185
R18894 VDD.n2359 VDD.n853 185
R18895 VDD.n853 VDD.n850 185
R18896 VDD.n2358 VDD.n2357 185
R18897 VDD.n2357 VDD.n2356 185
R18898 VDD.n855 VDD.n854 185
R18899 VDD.n856 VDD.n855 185
R18900 VDD.n2349 VDD.n2348 185
R18901 VDD.n2350 VDD.n2349 185
R18902 VDD.n2347 VDD.n865 185
R18903 VDD.n865 VDD.n862 185
R18904 VDD.n2346 VDD.n2345 185
R18905 VDD.n2345 VDD.n2344 185
R18906 VDD.n867 VDD.n866 185
R18907 VDD.n868 VDD.n867 185
R18908 VDD.n2337 VDD.n2336 185
R18909 VDD.n2338 VDD.n2337 185
R18910 VDD.n2335 VDD.n877 185
R18911 VDD.n877 VDD.n874 185
R18912 VDD.n2334 VDD.n2333 185
R18913 VDD.n2333 VDD.n2332 185
R18914 VDD.n879 VDD.n878 185
R18915 VDD.n880 VDD.n879 185
R18916 VDD.n2325 VDD.n2324 185
R18917 VDD.n2326 VDD.n2325 185
R18918 VDD.n2323 VDD.n889 185
R18919 VDD.n889 VDD.n886 185
R18920 VDD.n2322 VDD.n2321 185
R18921 VDD.n2321 VDD.n2320 185
R18922 VDD.n891 VDD.n890 185
R18923 VDD.n900 VDD.n891 185
R18924 VDD.n2313 VDD.n2312 185
R18925 VDD.n2314 VDD.n2313 185
R18926 VDD.n2311 VDD.n901 185
R18927 VDD.n901 VDD.n897 185
R18928 VDD.n2310 VDD.n2309 185
R18929 VDD.n2309 VDD.n2308 185
R18930 VDD.n903 VDD.n902 185
R18931 VDD.n904 VDD.n903 185
R18932 VDD.n2301 VDD.n2300 185
R18933 VDD.n2302 VDD.n2301 185
R18934 VDD.n2299 VDD.n913 185
R18935 VDD.n913 VDD.n910 185
R18936 VDD.n2298 VDD.n2297 185
R18937 VDD.n2297 VDD.n2296 185
R18938 VDD.n915 VDD.n914 185
R18939 VDD.n916 VDD.n915 185
R18940 VDD.n2289 VDD.n2288 185
R18941 VDD.n2290 VDD.n2289 185
R18942 VDD.n2287 VDD.n925 185
R18943 VDD.n925 VDD.n922 185
R18944 VDD.n2286 VDD.n2285 185
R18945 VDD.n2285 VDD.n2284 185
R18946 VDD.n927 VDD.n926 185
R18947 VDD.n928 VDD.n927 185
R18948 VDD.n2277 VDD.n2276 185
R18949 VDD.n2278 VDD.n2277 185
R18950 VDD.n2275 VDD.n937 185
R18951 VDD.n937 VDD.n934 185
R18952 VDD.n2274 VDD.n2273 185
R18953 VDD.n2273 VDD.n2272 185
R18954 VDD.n939 VDD.n938 185
R18955 VDD.n947 VDD.n939 185
R18956 VDD.n2265 VDD.n2264 185
R18957 VDD.n2266 VDD.n2265 185
R18958 VDD.n2263 VDD.n948 185
R18959 VDD.n954 VDD.n948 185
R18960 VDD.n2262 VDD.n2261 185
R18961 VDD.n2261 VDD.n2260 185
R18962 VDD.n950 VDD.n949 185
R18963 VDD.n951 VDD.n950 185
R18964 VDD.n2253 VDD.n2252 185
R18965 VDD.n2254 VDD.n2253 185
R18966 VDD.n2251 VDD.n961 185
R18967 VDD.n961 VDD.n958 185
R18968 VDD.n2250 VDD.n2249 185
R18969 VDD.n2249 VDD.n2248 185
R18970 VDD.n963 VDD.n962 185
R18971 VDD.n964 VDD.n963 185
R18972 VDD.n2241 VDD.n2240 185
R18973 VDD.n2242 VDD.n2241 185
R18974 VDD.n2239 VDD.n973 185
R18975 VDD.n973 VDD.n970 185
R18976 VDD.n2238 VDD.n2237 185
R18977 VDD.n2237 VDD.n2236 185
R18978 VDD.n975 VDD.n974 185
R18979 VDD.n976 VDD.n975 185
R18980 VDD.n2229 VDD.n2228 185
R18981 VDD.n2230 VDD.n2229 185
R18982 VDD.n2227 VDD.n985 185
R18983 VDD.n985 VDD.n982 185
R18984 VDD.n2226 VDD.n2225 185
R18985 VDD.n2225 VDD.n2224 185
R18986 VDD.n987 VDD.n986 185
R18987 VDD.n988 VDD.n987 185
R18988 VDD.n2217 VDD.n2216 185
R18989 VDD.n2218 VDD.n2217 185
R18990 VDD.n2215 VDD.n997 185
R18991 VDD.n997 VDD.n994 185
R18992 VDD.n2214 VDD.n2213 185
R18993 VDD.n2213 VDD.n2212 185
R18994 VDD.n999 VDD.n998 185
R18995 VDD.n1000 VDD.n999 185
R18996 VDD.n2205 VDD.n2204 185
R18997 VDD.n2206 VDD.n2205 185
R18998 VDD.n2203 VDD.n1009 185
R18999 VDD.n1009 VDD.n1006 185
R19000 VDD.n2202 VDD.n2201 185
R19001 VDD.n2201 VDD.n2200 185
R19002 VDD.n1011 VDD.n1010 185
R19003 VDD.n1012 VDD.n1011 185
R19004 VDD.n2193 VDD.n2192 185
R19005 VDD.n2194 VDD.n2193 185
R19006 VDD.n2191 VDD.n1021 185
R19007 VDD.n1021 VDD.n1018 185
R19008 VDD.n2190 VDD.n2189 185
R19009 VDD.n2189 VDD.n2188 185
R19010 VDD.n1023 VDD.n1022 185
R19011 VDD.n1032 VDD.n1023 185
R19012 VDD.n2181 VDD.n2180 185
R19013 VDD.n2182 VDD.n2181 185
R19014 VDD.n2179 VDD.n1033 185
R19015 VDD.n1033 VDD.n1029 185
R19016 VDD.n2178 VDD.n2177 185
R19017 VDD.n2177 VDD.n2176 185
R19018 VDD.n1035 VDD.n1034 185
R19019 VDD.n1036 VDD.n1035 185
R19020 VDD.n2169 VDD.n2168 185
R19021 VDD.n2170 VDD.n2169 185
R19022 VDD.n2167 VDD.n1045 185
R19023 VDD.n1045 VDD.n1042 185
R19024 VDD.n2166 VDD.n2165 185
R19025 VDD.n2165 VDD.n2164 185
R19026 VDD.n1047 VDD.n1046 185
R19027 VDD.n1048 VDD.n1047 185
R19028 VDD.n2157 VDD.n2156 185
R19029 VDD.n2158 VDD.n2157 185
R19030 VDD.n2155 VDD.n1057 185
R19031 VDD.n1057 VDD.n1054 185
R19032 VDD.n2154 VDD.n2153 185
R19033 VDD.n2153 VDD.n2152 185
R19034 VDD.n1059 VDD.n1058 185
R19035 VDD.n1060 VDD.n1059 185
R19036 VDD.n2145 VDD.n2144 185
R19037 VDD.n2146 VDD.n2145 185
R19038 VDD.n2143 VDD.n1069 185
R19039 VDD.n1069 VDD.n1066 185
R19040 VDD.n2142 VDD.n2141 185
R19041 VDD.n2141 VDD.n2140 185
R19042 VDD.n1071 VDD.n1070 185
R19043 VDD.n1080 VDD.n1071 185
R19044 VDD.n2133 VDD.n2132 185
R19045 VDD.n2134 VDD.n2133 185
R19046 VDD.n2131 VDD.n1081 185
R19047 VDD.n1081 VDD.n1077 185
R19048 VDD.n2130 VDD.n2129 185
R19049 VDD.n2129 VDD.n2128 185
R19050 VDD.n1083 VDD.n1082 185
R19051 VDD.n1084 VDD.n1083 185
R19052 VDD.n2121 VDD.n2120 185
R19053 VDD.n2122 VDD.n2121 185
R19054 VDD.n2119 VDD.n1093 185
R19055 VDD.n1093 VDD.n1090 185
R19056 VDD.n2118 VDD.n2117 185
R19057 VDD.n2117 VDD.n2116 185
R19058 VDD.n1095 VDD.n1094 185
R19059 VDD.n1096 VDD.n1095 185
R19060 VDD.n2109 VDD.n2108 185
R19061 VDD.n2110 VDD.n2109 185
R19062 VDD.n2107 VDD.n1105 185
R19063 VDD.n1105 VDD.n1102 185
R19064 VDD.n2106 VDD.n2105 185
R19065 VDD.n2105 VDD.n2104 185
R19066 VDD.n1107 VDD.n1106 185
R19067 VDD.n1146 VDD.n1144 185
R19068 VDD.n1147 VDD.n1143 185
R19069 VDD.n1147 VDD.n1108 185
R19070 VDD.n1150 VDD.n1149 185
R19071 VDD.n1151 VDD.n1142 185
R19072 VDD.n1153 VDD.n1152 185
R19073 VDD.n1155 VDD.n1141 185
R19074 VDD.n1158 VDD.n1157 185
R19075 VDD.n1698 VDD.n1140 185
R19076 VDD.n1700 VDD.n1699 185
R19077 VDD.n1702 VDD.n1139 185
R19078 VDD.n1705 VDD.n1704 185
R19079 VDD.n1707 VDD.n1136 185
R19080 VDD.n1709 VDD.n1708 185
R19081 VDD.n1711 VDD.n1135 185
R19082 VDD.n1713 VDD.n1712 185
R19083 VDD.n1712 VDD.n1108 185
R19084 VDD.n2516 VDD.n2515 185
R19085 VDD.n2518 VDD.n2517 185
R19086 VDD.n2520 VDD.n2519 185
R19087 VDD.n2522 VDD.n2521 185
R19088 VDD.n2524 VDD.n2523 185
R19089 VDD.n2526 VDD.n2525 185
R19090 VDD.n2528 VDD.n2527 185
R19091 VDD.n2530 VDD.n2529 185
R19092 VDD.n2532 VDD.n2531 185
R19093 VDD.n2534 VDD.n2533 185
R19094 VDD.n2536 VDD.n2535 185
R19095 VDD.n2538 VDD.n2537 185
R19096 VDD.n2540 VDD.n2539 185
R19097 VDD.n2542 VDD.n2541 185
R19098 VDD.n2544 VDD.n2543 185
R19099 VDD.n2546 VDD.n2545 185
R19100 VDD.n2514 VDD.n2513 185
R19101 VDD.n2514 VDD.n710 185
R19102 VDD.n2512 VDD.n732 185
R19103 VDD.n2550 VDD.n732 185
R19104 VDD.n2511 VDD.n2510 185
R19105 VDD.n2510 VDD.n731 185
R19106 VDD.n2509 VDD.n740 185
R19107 VDD.n2509 VDD.n2508 185
R19108 VDD.n1883 VDD.n741 185
R19109 VDD.n742 VDD.n741 185
R19110 VDD.n1884 VDD.n749 185
R19111 VDD.n2502 VDD.n749 185
R19112 VDD.n1886 VDD.n1885 185
R19113 VDD.n1885 VDD.n748 185
R19114 VDD.n1887 VDD.n756 185
R19115 VDD.n2458 VDD.n756 185
R19116 VDD.n1889 VDD.n1888 185
R19117 VDD.n1888 VDD.n755 185
R19118 VDD.n1890 VDD.n762 185
R19119 VDD.n2452 VDD.n762 185
R19120 VDD.n1892 VDD.n1891 185
R19121 VDD.n1891 VDD.n761 185
R19122 VDD.n1893 VDD.n767 185
R19123 VDD.n2446 VDD.n767 185
R19124 VDD.n1895 VDD.n1894 185
R19125 VDD.n1896 VDD.n1895 185
R19126 VDD.n1882 VDD.n773 185
R19127 VDD.n2440 VDD.n773 185
R19128 VDD.n1881 VDD.n1880 185
R19129 VDD.n1880 VDD.n772 185
R19130 VDD.n1879 VDD.n779 185
R19131 VDD.n2434 VDD.n779 185
R19132 VDD.n1878 VDD.n1877 185
R19133 VDD.n1877 VDD.n778 185
R19134 VDD.n1876 VDD.n785 185
R19135 VDD.n2428 VDD.n785 185
R19136 VDD.n1875 VDD.n1874 185
R19137 VDD.n1874 VDD.n784 185
R19138 VDD.n1873 VDD.n791 185
R19139 VDD.n2422 VDD.n791 185
R19140 VDD.n1872 VDD.n1871 185
R19141 VDD.n1871 VDD.n790 185
R19142 VDD.n1870 VDD.n797 185
R19143 VDD.n2416 VDD.n797 185
R19144 VDD.n1869 VDD.n1868 185
R19145 VDD.n1868 VDD.n796 185
R19146 VDD.n1867 VDD.n803 185
R19147 VDD.n2410 VDD.n803 185
R19148 VDD.n1866 VDD.n1865 185
R19149 VDD.n1865 VDD.n802 185
R19150 VDD.n1864 VDD.n809 185
R19151 VDD.n2404 VDD.n809 185
R19152 VDD.n1863 VDD.n1862 185
R19153 VDD.n1862 VDD.n808 185
R19154 VDD.n1861 VDD.n815 185
R19155 VDD.n2398 VDD.n815 185
R19156 VDD.n1860 VDD.n1859 185
R19157 VDD.n1859 VDD.n814 185
R19158 VDD.n1858 VDD.n821 185
R19159 VDD.n2392 VDD.n821 185
R19160 VDD.n1857 VDD.n1856 185
R19161 VDD.n1856 VDD.n820 185
R19162 VDD.n1855 VDD.n826 185
R19163 VDD.n2386 VDD.n826 185
R19164 VDD.n1854 VDD.n1853 185
R19165 VDD.n1853 VDD.n834 185
R19166 VDD.n1852 VDD.n832 185
R19167 VDD.n2380 VDD.n832 185
R19168 VDD.n1851 VDD.n1850 185
R19169 VDD.n1850 VDD.n831 185
R19170 VDD.n1849 VDD.n839 185
R19171 VDD.n2374 VDD.n839 185
R19172 VDD.n1848 VDD.n1847 185
R19173 VDD.n1847 VDD.n838 185
R19174 VDD.n1846 VDD.n845 185
R19175 VDD.n2368 VDD.n845 185
R19176 VDD.n1845 VDD.n1844 185
R19177 VDD.n1844 VDD.n844 185
R19178 VDD.n1843 VDD.n851 185
R19179 VDD.n2362 VDD.n851 185
R19180 VDD.n1842 VDD.n1841 185
R19181 VDD.n1841 VDD.n850 185
R19182 VDD.n1840 VDD.n857 185
R19183 VDD.n2356 VDD.n857 185
R19184 VDD.n1839 VDD.n1838 185
R19185 VDD.n1838 VDD.n856 185
R19186 VDD.n1837 VDD.n863 185
R19187 VDD.n2350 VDD.n863 185
R19188 VDD.n1836 VDD.n1835 185
R19189 VDD.n1835 VDD.n862 185
R19190 VDD.n1834 VDD.n869 185
R19191 VDD.n2344 VDD.n869 185
R19192 VDD.n1833 VDD.n1832 185
R19193 VDD.n1832 VDD.n868 185
R19194 VDD.n1831 VDD.n875 185
R19195 VDD.n2338 VDD.n875 185
R19196 VDD.n1830 VDD.n1829 185
R19197 VDD.n1829 VDD.n874 185
R19198 VDD.n1828 VDD.n881 185
R19199 VDD.n2332 VDD.n881 185
R19200 VDD.n1827 VDD.n1826 185
R19201 VDD.n1826 VDD.n880 185
R19202 VDD.n1825 VDD.n887 185
R19203 VDD.n2326 VDD.n887 185
R19204 VDD.n1824 VDD.n1823 185
R19205 VDD.n1823 VDD.n886 185
R19206 VDD.n1822 VDD.n892 185
R19207 VDD.n2320 VDD.n892 185
R19208 VDD.n1821 VDD.n1820 185
R19209 VDD.n1820 VDD.n900 185
R19210 VDD.n1819 VDD.n898 185
R19211 VDD.n2314 VDD.n898 185
R19212 VDD.n1818 VDD.n1817 185
R19213 VDD.n1817 VDD.n897 185
R19214 VDD.n1816 VDD.n905 185
R19215 VDD.n2308 VDD.n905 185
R19216 VDD.n1815 VDD.n1814 185
R19217 VDD.n1814 VDD.n904 185
R19218 VDD.n1813 VDD.n911 185
R19219 VDD.n2302 VDD.n911 185
R19220 VDD.n1812 VDD.n1811 185
R19221 VDD.n1811 VDD.n910 185
R19222 VDD.n1810 VDD.n917 185
R19223 VDD.n2296 VDD.n917 185
R19224 VDD.n1809 VDD.n1808 185
R19225 VDD.n1808 VDD.n916 185
R19226 VDD.n1807 VDD.n923 185
R19227 VDD.n2290 VDD.n923 185
R19228 VDD.n1806 VDD.n1805 185
R19229 VDD.n1805 VDD.n922 185
R19230 VDD.n1804 VDD.n929 185
R19231 VDD.n2284 VDD.n929 185
R19232 VDD.n1803 VDD.n1802 185
R19233 VDD.n1802 VDD.n928 185
R19234 VDD.n1801 VDD.n935 185
R19235 VDD.n2278 VDD.n935 185
R19236 VDD.n1800 VDD.n1799 185
R19237 VDD.n1799 VDD.n934 185
R19238 VDD.n1798 VDD.n940 185
R19239 VDD.n2272 VDD.n940 185
R19240 VDD.n1797 VDD.n1796 185
R19241 VDD.n1796 VDD.n947 185
R19242 VDD.n1795 VDD.n945 185
R19243 VDD.n2266 VDD.n945 185
R19244 VDD.n1794 VDD.n1793 185
R19245 VDD.n1793 VDD.n954 185
R19246 VDD.n1792 VDD.n952 185
R19247 VDD.n2260 VDD.n952 185
R19248 VDD.n1791 VDD.n1790 185
R19249 VDD.n1790 VDD.n951 185
R19250 VDD.n1789 VDD.n959 185
R19251 VDD.n2254 VDD.n959 185
R19252 VDD.n1788 VDD.n1787 185
R19253 VDD.n1787 VDD.n958 185
R19254 VDD.n1786 VDD.n965 185
R19255 VDD.n2248 VDD.n965 185
R19256 VDD.n1785 VDD.n1784 185
R19257 VDD.n1784 VDD.n964 185
R19258 VDD.n1783 VDD.n971 185
R19259 VDD.n2242 VDD.n971 185
R19260 VDD.n1782 VDD.n1781 185
R19261 VDD.n1781 VDD.n970 185
R19262 VDD.n1780 VDD.n977 185
R19263 VDD.n2236 VDD.n977 185
R19264 VDD.n1779 VDD.n1778 185
R19265 VDD.n1778 VDD.n976 185
R19266 VDD.n1777 VDD.n983 185
R19267 VDD.n2230 VDD.n983 185
R19268 VDD.n1776 VDD.n1775 185
R19269 VDD.n1775 VDD.n982 185
R19270 VDD.n1774 VDD.n989 185
R19271 VDD.n2224 VDD.n989 185
R19272 VDD.n1773 VDD.n1772 185
R19273 VDD.n1772 VDD.n988 185
R19274 VDD.n1771 VDD.n995 185
R19275 VDD.n2218 VDD.n995 185
R19276 VDD.n1770 VDD.n1769 185
R19277 VDD.n1769 VDD.n994 185
R19278 VDD.n1768 VDD.n1001 185
R19279 VDD.n2212 VDD.n1001 185
R19280 VDD.n1767 VDD.n1766 185
R19281 VDD.n1766 VDD.n1000 185
R19282 VDD.n1765 VDD.n1007 185
R19283 VDD.n2206 VDD.n1007 185
R19284 VDD.n1764 VDD.n1763 185
R19285 VDD.n1763 VDD.n1006 185
R19286 VDD.n1762 VDD.n1013 185
R19287 VDD.n2200 VDD.n1013 185
R19288 VDD.n1761 VDD.n1760 185
R19289 VDD.n1760 VDD.n1012 185
R19290 VDD.n1759 VDD.n1019 185
R19291 VDD.n2194 VDD.n1019 185
R19292 VDD.n1758 VDD.n1757 185
R19293 VDD.n1757 VDD.n1018 185
R19294 VDD.n1756 VDD.n1024 185
R19295 VDD.n2188 VDD.n1024 185
R19296 VDD.n1755 VDD.n1754 185
R19297 VDD.n1754 VDD.n1032 185
R19298 VDD.n1753 VDD.n1030 185
R19299 VDD.n2182 VDD.n1030 185
R19300 VDD.n1752 VDD.n1751 185
R19301 VDD.n1751 VDD.n1029 185
R19302 VDD.n1750 VDD.n1037 185
R19303 VDD.n2176 VDD.n1037 185
R19304 VDD.n1749 VDD.n1748 185
R19305 VDD.n1748 VDD.n1036 185
R19306 VDD.n1747 VDD.n1043 185
R19307 VDD.n2170 VDD.n1043 185
R19308 VDD.n1746 VDD.n1745 185
R19309 VDD.n1745 VDD.n1042 185
R19310 VDD.n1744 VDD.n1049 185
R19311 VDD.n2164 VDD.n1049 185
R19312 VDD.n1743 VDD.n1742 185
R19313 VDD.n1742 VDD.n1048 185
R19314 VDD.n1741 VDD.n1055 185
R19315 VDD.n2158 VDD.n1055 185
R19316 VDD.n1740 VDD.n1739 185
R19317 VDD.n1739 VDD.n1054 185
R19318 VDD.n1738 VDD.n1061 185
R19319 VDD.n2152 VDD.n1061 185
R19320 VDD.n1737 VDD.n1736 185
R19321 VDD.n1736 VDD.n1060 185
R19322 VDD.n1735 VDD.n1067 185
R19323 VDD.n2146 VDD.n1067 185
R19324 VDD.n1734 VDD.n1733 185
R19325 VDD.n1733 VDD.n1066 185
R19326 VDD.n1732 VDD.n1072 185
R19327 VDD.n2140 VDD.n1072 185
R19328 VDD.n1731 VDD.n1730 185
R19329 VDD.n1730 VDD.n1080 185
R19330 VDD.n1729 VDD.n1078 185
R19331 VDD.n2134 VDD.n1078 185
R19332 VDD.n1728 VDD.n1727 185
R19333 VDD.n1727 VDD.n1077 185
R19334 VDD.n1726 VDD.n1085 185
R19335 VDD.n2128 VDD.n1085 185
R19336 VDD.n1725 VDD.n1724 185
R19337 VDD.n1724 VDD.n1084 185
R19338 VDD.n1723 VDD.n1091 185
R19339 VDD.n2122 VDD.n1091 185
R19340 VDD.n1722 VDD.n1721 185
R19341 VDD.n1721 VDD.n1090 185
R19342 VDD.n1720 VDD.n1097 185
R19343 VDD.n2116 VDD.n1097 185
R19344 VDD.n1719 VDD.n1718 185
R19345 VDD.n1718 VDD.n1096 185
R19346 VDD.n1717 VDD.n1103 185
R19347 VDD.n2110 VDD.n1103 185
R19348 VDD.n1716 VDD.n1715 185
R19349 VDD.n1715 VDD.n1102 185
R19350 VDD.n1714 VDD.n1109 185
R19351 VDD.n2104 VDD.n1109 185
R19352 VDD.n80 VDD.n79 185
R19353 VDD.n3664 VDD.n80 185
R19354 VDD.n3667 VDD.n3666 185
R19355 VDD.n3666 VDD.n3665 185
R19356 VDD.n3668 VDD.n74 185
R19357 VDD.n74 VDD.n73 185
R19358 VDD.n3670 VDD.n3669 185
R19359 VDD.n3671 VDD.n3670 185
R19360 VDD.n69 VDD.n68 185
R19361 VDD.n3672 VDD.n69 185
R19362 VDD.n3675 VDD.n3674 185
R19363 VDD.n3674 VDD.n3673 185
R19364 VDD.n3676 VDD.n63 185
R19365 VDD.n63 VDD.n62 185
R19366 VDD.n3678 VDD.n3677 185
R19367 VDD.n3679 VDD.n3678 185
R19368 VDD.n58 VDD.n57 185
R19369 VDD.n3680 VDD.n58 185
R19370 VDD.n3683 VDD.n3682 185
R19371 VDD.n3682 VDD.n3681 185
R19372 VDD.n3684 VDD.n52 185
R19373 VDD.n52 VDD.n51 185
R19374 VDD.n3686 VDD.n3685 185
R19375 VDD.n3687 VDD.n3686 185
R19376 VDD.n47 VDD.n46 185
R19377 VDD.n3688 VDD.n47 185
R19378 VDD.n3691 VDD.n3690 185
R19379 VDD.n3690 VDD.n3689 185
R19380 VDD.n3692 VDD.n41 185
R19381 VDD.n41 VDD.n40 185
R19382 VDD.n3694 VDD.n3693 185
R19383 VDD.n3695 VDD.n3694 185
R19384 VDD.n36 VDD.n35 185
R19385 VDD.n3696 VDD.n36 185
R19386 VDD.n3699 VDD.n3698 185
R19387 VDD.n3698 VDD.n3697 185
R19388 VDD.n3700 VDD.n30 185
R19389 VDD.n30 VDD.n29 185
R19390 VDD.n3702 VDD.n3701 185
R19391 VDD.n3703 VDD.n3702 185
R19392 VDD.n24 VDD.n23 185
R19393 VDD.n3704 VDD.n24 185
R19394 VDD.n3707 VDD.n3706 185
R19395 VDD.n3706 VDD.n3705 185
R19396 VDD.n3708 VDD.n22 185
R19397 VDD.n25 VDD.n22 185
R19398 VDD.n3616 VDD.n21 185
R19399 VDD.n3617 VDD.n3616 185
R19400 VDD.n3615 VDD.n3614 185
R19401 VDD.n3615 VDD.n196 185
R19402 VDD.n198 VDD.n197 185
R19403 VDD.n3607 VDD.n197 185
R19404 VDD.n3610 VDD.n3609 185
R19405 VDD.n3609 VDD.n3608 185
R19406 VDD.n201 VDD.n200 185
R19407 VDD.n202 VDD.n201 185
R19408 VDD.n3594 VDD.n3593 185
R19409 VDD.n3595 VDD.n3594 185
R19410 VDD.n210 VDD.n209 185
R19411 VDD.n209 VDD.n208 185
R19412 VDD.n3589 VDD.n3588 185
R19413 VDD.n3588 VDD.n3587 185
R19414 VDD.n213 VDD.n212 185
R19415 VDD.n214 VDD.n213 185
R19416 VDD.n3576 VDD.n3575 185
R19417 VDD.n3577 VDD.n3576 185
R19418 VDD.n222 VDD.n221 185
R19419 VDD.n221 VDD.n220 185
R19420 VDD.n3571 VDD.n3570 185
R19421 VDD.n3570 VDD.n3569 185
R19422 VDD.n225 VDD.n224 185
R19423 VDD.n226 VDD.n225 185
R19424 VDD.n3560 VDD.n3559 185
R19425 VDD.n3561 VDD.n3560 185
R19426 VDD.n234 VDD.n233 185
R19427 VDD.n233 VDD.n232 185
R19428 VDD.n3555 VDD.n3554 185
R19429 VDD.n3554 VDD.n3553 185
R19430 VDD.n237 VDD.n236 185
R19431 VDD.n238 VDD.n237 185
R19432 VDD.n3544 VDD.n3543 185
R19433 VDD.n3545 VDD.n3544 185
R19434 VDD.n246 VDD.n245 185
R19435 VDD.n245 VDD.n244 185
R19436 VDD.n3539 VDD.n3538 185
R19437 VDD.n3538 VDD.n3537 185
R19438 VDD.n249 VDD.n248 185
R19439 VDD.n250 VDD.n249 185
R19440 VDD.n3528 VDD.n3527 185
R19441 VDD.n3529 VDD.n3528 185
R19442 VDD.n258 VDD.n257 185
R19443 VDD.n257 VDD.n256 185
R19444 VDD.n3521 VDD.n3520 185
R19445 VDD.n263 VDD.n262 185
R19446 VDD.n3517 VDD.n3516 185
R19447 VDD.n3518 VDD.n3517 185
R19448 VDD.n3515 VDD.n277 185
R19449 VDD.n3514 VDD.n3513 185
R19450 VDD.n3512 VDD.n3511 185
R19451 VDD.n3510 VDD.n3509 185
R19452 VDD.n3508 VDD.n3507 185
R19453 VDD.n3506 VDD.n3505 185
R19454 VDD.n3504 VDD.n3503 185
R19455 VDD.n3502 VDD.n3501 185
R19456 VDD.n3500 VDD.n3499 185
R19457 VDD.n3498 VDD.n288 185
R19458 VDD.n3497 VDD.n3496 185
R19459 VDD.n3495 VDD.n3494 185
R19460 VDD.n3493 VDD.n3492 185
R19461 VDD.n3491 VDD.n3490 185
R19462 VDD.n3489 VDD.n3488 185
R19463 VDD.n3487 VDD.n3486 185
R19464 VDD.n3485 VDD.n3484 185
R19465 VDD.n3483 VDD.n3482 185
R19466 VDD.n3481 VDD.n3480 185
R19467 VDD.n3479 VDD.n3478 185
R19468 VDD.n3477 VDD.n3476 185
R19469 VDD.n3475 VDD.n3474 185
R19470 VDD.n3473 VDD.n3472 185
R19471 VDD.n307 VDD.n304 185
R19472 VDD.n3468 VDD.n276 185
R19473 VDD.n3518 VDD.n276 185
R19474 VDD.n3661 VDD.n3660 185
R19475 VDD.n99 VDD.n96 185
R19476 VDD.n179 VDD.n178 185
R19477 VDD.n177 VDD.n176 185
R19478 VDD.n175 VDD.n174 185
R19479 VDD.n168 VDD.n101 185
R19480 VDD.n170 VDD.n169 185
R19481 VDD.n167 VDD.n166 185
R19482 VDD.n165 VDD.n164 185
R19483 VDD.n158 VDD.n103 185
R19484 VDD.n160 VDD.n159 185
R19485 VDD.n157 VDD.n156 185
R19486 VDD.n155 VDD.n154 185
R19487 VDD.n148 VDD.n105 185
R19488 VDD.n150 VDD.n149 185
R19489 VDD.n147 VDD.n109 185
R19490 VDD.n146 VDD.n145 185
R19491 VDD.n139 VDD.n110 185
R19492 VDD.n141 VDD.n140 185
R19493 VDD.n138 VDD.n137 185
R19494 VDD.n136 VDD.n135 185
R19495 VDD.n129 VDD.n112 185
R19496 VDD.n131 VDD.n130 185
R19497 VDD.n128 VDD.n127 185
R19498 VDD.n126 VDD.n125 185
R19499 VDD.n119 VDD.n114 185
R19500 VDD.n121 VDD.n120 185
R19501 VDD.n118 VDD.n117 185
R19502 VDD.n3657 VDD.n82 185
R19503 VDD.n3664 VDD.n82 185
R19504 VDD.n3656 VDD.n81 185
R19505 VDD.n3665 VDD.n81 185
R19506 VDD.n3655 VDD.n3654 185
R19507 VDD.n3654 VDD.n73 185
R19508 VDD.n183 VDD.n72 185
R19509 VDD.n3671 VDD.n72 185
R19510 VDD.n3650 VDD.n71 185
R19511 VDD.n3672 VDD.n71 185
R19512 VDD.n3649 VDD.n70 185
R19513 VDD.n3673 VDD.n70 185
R19514 VDD.n3648 VDD.n3647 185
R19515 VDD.n3647 VDD.n62 185
R19516 VDD.n185 VDD.n61 185
R19517 VDD.n3679 VDD.n61 185
R19518 VDD.n3643 VDD.n60 185
R19519 VDD.n3680 VDD.n60 185
R19520 VDD.n3642 VDD.n59 185
R19521 VDD.n3681 VDD.n59 185
R19522 VDD.n3641 VDD.n3640 185
R19523 VDD.n3640 VDD.n51 185
R19524 VDD.n187 VDD.n50 185
R19525 VDD.n3687 VDD.n50 185
R19526 VDD.n3636 VDD.n49 185
R19527 VDD.n3688 VDD.n49 185
R19528 VDD.n3635 VDD.n48 185
R19529 VDD.n3689 VDD.n48 185
R19530 VDD.n3634 VDD.n3633 185
R19531 VDD.n3633 VDD.n40 185
R19532 VDD.n189 VDD.n39 185
R19533 VDD.n3695 VDD.n39 185
R19534 VDD.n3629 VDD.n38 185
R19535 VDD.n3696 VDD.n38 185
R19536 VDD.n3628 VDD.n37 185
R19537 VDD.n3697 VDD.n37 185
R19538 VDD.n3627 VDD.n3626 185
R19539 VDD.n3626 VDD.n29 185
R19540 VDD.n191 VDD.n28 185
R19541 VDD.n3703 VDD.n28 185
R19542 VDD.n3622 VDD.n27 185
R19543 VDD.n3704 VDD.n27 185
R19544 VDD.n3621 VDD.n26 185
R19545 VDD.n3705 VDD.n26 185
R19546 VDD.n3620 VDD.n3619 185
R19547 VDD.n3619 VDD.n25 185
R19548 VDD.n3618 VDD.n193 185
R19549 VDD.n3618 VDD.n3617 185
R19550 VDD.n3604 VDD.n195 185
R19551 VDD.n196 VDD.n195 185
R19552 VDD.n3606 VDD.n3605 185
R19553 VDD.n3607 VDD.n3606 185
R19554 VDD.n204 VDD.n203 185
R19555 VDD.n3608 VDD.n203 185
R19556 VDD.n3598 VDD.n3597 185
R19557 VDD.n3597 VDD.n202 185
R19558 VDD.n3596 VDD.n206 185
R19559 VDD.n3596 VDD.n3595 185
R19560 VDD.n3584 VDD.n207 185
R19561 VDD.n208 VDD.n207 185
R19562 VDD.n3586 VDD.n3585 185
R19563 VDD.n3587 VDD.n3586 185
R19564 VDD.n216 VDD.n215 185
R19565 VDD.n215 VDD.n214 185
R19566 VDD.n3579 VDD.n3578 185
R19567 VDD.n3578 VDD.n3577 185
R19568 VDD.n219 VDD.n218 185
R19569 VDD.n220 VDD.n219 185
R19570 VDD.n3568 VDD.n3567 185
R19571 VDD.n3569 VDD.n3568 185
R19572 VDD.n228 VDD.n227 185
R19573 VDD.n227 VDD.n226 185
R19574 VDD.n3563 VDD.n3562 185
R19575 VDD.n3562 VDD.n3561 185
R19576 VDD.n231 VDD.n230 185
R19577 VDD.n232 VDD.n231 185
R19578 VDD.n3552 VDD.n3551 185
R19579 VDD.n3553 VDD.n3552 185
R19580 VDD.n240 VDD.n239 185
R19581 VDD.n239 VDD.n238 185
R19582 VDD.n3547 VDD.n3546 185
R19583 VDD.n3546 VDD.n3545 185
R19584 VDD.n243 VDD.n242 185
R19585 VDD.n244 VDD.n243 185
R19586 VDD.n3536 VDD.n3535 185
R19587 VDD.n3537 VDD.n3536 185
R19588 VDD.n252 VDD.n251 185
R19589 VDD.n251 VDD.n250 185
R19590 VDD.n3531 VDD.n3530 185
R19591 VDD.n3530 VDD.n3529 185
R19592 VDD.n255 VDD.n254 185
R19593 VDD.n256 VDD.n255 185
R19594 VDD.n709 VDD.n708 185
R19595 VDD.n2570 VDD.n2569 185
R19596 VDD.n2571 VDD.n2567 185
R19597 VDD.n2567 VDD.n2558 185
R19598 VDD.n2573 VDD.n2572 185
R19599 VDD.n2575 VDD.n2566 185
R19600 VDD.n2578 VDD.n2577 185
R19601 VDD.n2579 VDD.n2565 185
R19602 VDD.n2581 VDD.n2580 185
R19603 VDD.n2583 VDD.n2564 185
R19604 VDD.n2586 VDD.n2585 185
R19605 VDD.n2587 VDD.n2563 185
R19606 VDD.n2592 VDD.n2591 185
R19607 VDD.n2594 VDD.n2562 185
R19608 VDD.n2595 VDD.n2561 185
R19609 VDD.n2598 VDD.n2597 185
R19610 VDD.n2599 VDD.n2559 185
R19611 VDD.n2559 VDD.n2558 185
R19612 VDD.n3412 VDD.n3411 185
R19613 VDD.n3413 VDD.n340 185
R19614 VDD.n3415 VDD.n3414 185
R19615 VDD.n3417 VDD.n339 185
R19616 VDD.n3419 VDD.n3418 185
R19617 VDD.n3420 VDD.n334 185
R19618 VDD.n3422 VDD.n3421 185
R19619 VDD.n3424 VDD.n333 185
R19620 VDD.n3426 VDD.n3425 185
R19621 VDD.n3428 VDD.n331 185
R19622 VDD.n3430 VDD.n3429 185
R19623 VDD.n3431 VDD.n330 185
R19624 VDD.n3433 VDD.n3432 185
R19625 VDD.n3435 VDD.n329 185
R19626 VDD.n3436 VDD.n328 185
R19627 VDD.n3439 VDD.n3438 185
R19628 VDD.n3410 VDD.n3408 185
R19629 VDD.n3410 VDD.n323 185
R19630 VDD.n3407 VDD.n322 185
R19631 VDD.n3443 VDD.n322 185
R19632 VDD.n3406 VDD.n3405 185
R19633 VDD.n3405 VDD.n321 185
R19634 VDD.n3404 VDD.n341 185
R19635 VDD.n3404 VDD.n3403 185
R19636 VDD.n2600 VDD.n342 185
R19637 VDD.n343 VDD.n342 185
R19638 VDD.n2601 VDD.n350 185
R19639 VDD.n3397 VDD.n350 185
R19640 VDD.n2603 VDD.n2602 185
R19641 VDD.n2602 VDD.n349 185
R19642 VDD.n2604 VDD.n357 185
R19643 VDD.n3366 VDD.n357 185
R19644 VDD.n2606 VDD.n2605 185
R19645 VDD.n2605 VDD.n356 185
R19646 VDD.n2607 VDD.n363 185
R19647 VDD.n3360 VDD.n363 185
R19648 VDD.n2609 VDD.n2608 185
R19649 VDD.n2608 VDD.n362 185
R19650 VDD.n2610 VDD.n368 185
R19651 VDD.n3354 VDD.n368 185
R19652 VDD.n2612 VDD.n2611 185
R19653 VDD.n2611 VDD.n376 185
R19654 VDD.n2613 VDD.n374 185
R19655 VDD.n3348 VDD.n374 185
R19656 VDD.n2615 VDD.n2614 185
R19657 VDD.n2614 VDD.n373 185
R19658 VDD.n2616 VDD.n381 185
R19659 VDD.n3342 VDD.n381 185
R19660 VDD.n2618 VDD.n2617 185
R19661 VDD.n2617 VDD.n380 185
R19662 VDD.n2619 VDD.n387 185
R19663 VDD.n3336 VDD.n387 185
R19664 VDD.n2621 VDD.n2620 185
R19665 VDD.n2620 VDD.n386 185
R19666 VDD.n2622 VDD.n393 185
R19667 VDD.n3330 VDD.n393 185
R19668 VDD.n2624 VDD.n2623 185
R19669 VDD.n2623 VDD.n392 185
R19670 VDD.n2625 VDD.n399 185
R19671 VDD.n3324 VDD.n399 185
R19672 VDD.n2627 VDD.n2626 185
R19673 VDD.n2626 VDD.n398 185
R19674 VDD.n2628 VDD.n405 185
R19675 VDD.n3318 VDD.n405 185
R19676 VDD.n2630 VDD.n2629 185
R19677 VDD.n2629 VDD.n404 185
R19678 VDD.n2631 VDD.n411 185
R19679 VDD.n3312 VDD.n411 185
R19680 VDD.n2633 VDD.n2632 185
R19681 VDD.n2632 VDD.n410 185
R19682 VDD.n2634 VDD.n416 185
R19683 VDD.n3306 VDD.n416 185
R19684 VDD.n2636 VDD.n2635 185
R19685 VDD.n2635 VDD.n424 185
R19686 VDD.n2637 VDD.n422 185
R19687 VDD.n3300 VDD.n422 185
R19688 VDD.n2639 VDD.n2638 185
R19689 VDD.n2638 VDD.n421 185
R19690 VDD.n2640 VDD.n429 185
R19691 VDD.n3294 VDD.n429 185
R19692 VDD.n2642 VDD.n2641 185
R19693 VDD.n2641 VDD.n428 185
R19694 VDD.n2643 VDD.n435 185
R19695 VDD.n3288 VDD.n435 185
R19696 VDD.n2645 VDD.n2644 185
R19697 VDD.n2644 VDD.n434 185
R19698 VDD.n2646 VDD.n441 185
R19699 VDD.n3282 VDD.n441 185
R19700 VDD.n2648 VDD.n2647 185
R19701 VDD.n2647 VDD.n440 185
R19702 VDD.n2649 VDD.n447 185
R19703 VDD.n3276 VDD.n447 185
R19704 VDD.n2651 VDD.n2650 185
R19705 VDD.n2650 VDD.n446 185
R19706 VDD.n2652 VDD.n453 185
R19707 VDD.n3270 VDD.n453 185
R19708 VDD.n2654 VDD.n2653 185
R19709 VDD.n2653 VDD.n452 185
R19710 VDD.n2655 VDD.n459 185
R19711 VDD.n3264 VDD.n459 185
R19712 VDD.n2657 VDD.n2656 185
R19713 VDD.n2656 VDD.n458 185
R19714 VDD.n2658 VDD.n465 185
R19715 VDD.n3258 VDD.n465 185
R19716 VDD.n2660 VDD.n2659 185
R19717 VDD.n2659 VDD.n464 185
R19718 VDD.n2661 VDD.n471 185
R19719 VDD.n3252 VDD.n471 185
R19720 VDD.n2663 VDD.n2662 185
R19721 VDD.n2662 VDD.n470 185
R19722 VDD.n2664 VDD.n477 185
R19723 VDD.n3246 VDD.n477 185
R19724 VDD.n2666 VDD.n2665 185
R19725 VDD.n2665 VDD.n476 185
R19726 VDD.n2667 VDD.n483 185
R19727 VDD.n3240 VDD.n483 185
R19728 VDD.n2669 VDD.n2668 185
R19729 VDD.n2668 VDD.n482 185
R19730 VDD.n2670 VDD.n489 185
R19731 VDD.n3234 VDD.n489 185
R19732 VDD.n2672 VDD.n2671 185
R19733 VDD.n2671 VDD.n488 185
R19734 VDD.n2673 VDD.n494 185
R19735 VDD.n3228 VDD.n494 185
R19736 VDD.n2675 VDD.n2674 185
R19737 VDD.n2674 VDD.n501 185
R19738 VDD.n2676 VDD.n499 185
R19739 VDD.n3222 VDD.n499 185
R19740 VDD.n2678 VDD.n2677 185
R19741 VDD.n2677 VDD.n508 185
R19742 VDD.n2679 VDD.n506 185
R19743 VDD.n3216 VDD.n506 185
R19744 VDD.n2681 VDD.n2680 185
R19745 VDD.n2680 VDD.n505 185
R19746 VDD.n2682 VDD.n513 185
R19747 VDD.n3210 VDD.n513 185
R19748 VDD.n2684 VDD.n2683 185
R19749 VDD.n2683 VDD.n512 185
R19750 VDD.n2685 VDD.n519 185
R19751 VDD.n3204 VDD.n519 185
R19752 VDD.n2687 VDD.n2686 185
R19753 VDD.n2686 VDD.n518 185
R19754 VDD.n2688 VDD.n525 185
R19755 VDD.n3198 VDD.n525 185
R19756 VDD.n2690 VDD.n2689 185
R19757 VDD.n2689 VDD.n524 185
R19758 VDD.n2691 VDD.n531 185
R19759 VDD.n3192 VDD.n531 185
R19760 VDD.n2693 VDD.n2692 185
R19761 VDD.n2692 VDD.n530 185
R19762 VDD.n2694 VDD.n537 185
R19763 VDD.n3186 VDD.n537 185
R19764 VDD.n2696 VDD.n2695 185
R19765 VDD.n2695 VDD.n536 185
R19766 VDD.n2697 VDD.n543 185
R19767 VDD.n3180 VDD.n543 185
R19768 VDD.n2699 VDD.n2698 185
R19769 VDD.n2698 VDD.n542 185
R19770 VDD.n2700 VDD.n548 185
R19771 VDD.n3174 VDD.n548 185
R19772 VDD.n2702 VDD.n2701 185
R19773 VDD.n2701 VDD.n556 185
R19774 VDD.n2703 VDD.n554 185
R19775 VDD.n3168 VDD.n554 185
R19776 VDD.n2705 VDD.n2704 185
R19777 VDD.n2704 VDD.n553 185
R19778 VDD.n2706 VDD.n561 185
R19779 VDD.n3162 VDD.n561 185
R19780 VDD.n2708 VDD.n2707 185
R19781 VDD.n2707 VDD.n560 185
R19782 VDD.n2709 VDD.n567 185
R19783 VDD.n3156 VDD.n567 185
R19784 VDD.n2711 VDD.n2710 185
R19785 VDD.n2710 VDD.n566 185
R19786 VDD.n2712 VDD.n573 185
R19787 VDD.n3150 VDD.n573 185
R19788 VDD.n2714 VDD.n2713 185
R19789 VDD.n2713 VDD.n572 185
R19790 VDD.n2715 VDD.n579 185
R19791 VDD.n3144 VDD.n579 185
R19792 VDD.n2717 VDD.n2716 185
R19793 VDD.n2716 VDD.n578 185
R19794 VDD.n2718 VDD.n585 185
R19795 VDD.n3138 VDD.n585 185
R19796 VDD.n2720 VDD.n2719 185
R19797 VDD.n2719 VDD.n584 185
R19798 VDD.n2721 VDD.n591 185
R19799 VDD.n3132 VDD.n591 185
R19800 VDD.n2723 VDD.n2722 185
R19801 VDD.n2722 VDD.n590 185
R19802 VDD.n2724 VDD.n597 185
R19803 VDD.n3126 VDD.n597 185
R19804 VDD.n2726 VDD.n2725 185
R19805 VDD.n2725 VDD.n596 185
R19806 VDD.n2727 VDD.n603 185
R19807 VDD.n3120 VDD.n603 185
R19808 VDD.n2729 VDD.n2728 185
R19809 VDD.n2728 VDD.n602 185
R19810 VDD.n2730 VDD.n609 185
R19811 VDD.n3114 VDD.n609 185
R19812 VDD.n2732 VDD.n2731 185
R19813 VDD.n2731 VDD.n608 185
R19814 VDD.n2733 VDD.n614 185
R19815 VDD.n3108 VDD.n614 185
R19816 VDD.n2735 VDD.n2734 185
R19817 VDD.n2734 VDD.n622 185
R19818 VDD.n2736 VDD.n620 185
R19819 VDD.n3102 VDD.n620 185
R19820 VDD.n2738 VDD.n2737 185
R19821 VDD.n2737 VDD.n619 185
R19822 VDD.n2739 VDD.n627 185
R19823 VDD.n3096 VDD.n627 185
R19824 VDD.n2741 VDD.n2740 185
R19825 VDD.n2740 VDD.n626 185
R19826 VDD.n2742 VDD.n633 185
R19827 VDD.n3090 VDD.n633 185
R19828 VDD.n2744 VDD.n2743 185
R19829 VDD.n2743 VDD.n632 185
R19830 VDD.n2745 VDD.n639 185
R19831 VDD.n3084 VDD.n639 185
R19832 VDD.n2747 VDD.n2746 185
R19833 VDD.n2746 VDD.n638 185
R19834 VDD.n2748 VDD.n645 185
R19835 VDD.n3078 VDD.n645 185
R19836 VDD.n2750 VDD.n2749 185
R19837 VDD.n2749 VDD.n644 185
R19838 VDD.n2751 VDD.n651 185
R19839 VDD.n3072 VDD.n651 185
R19840 VDD.n2753 VDD.n2752 185
R19841 VDD.n2752 VDD.n650 185
R19842 VDD.n2754 VDD.n657 185
R19843 VDD.n3066 VDD.n657 185
R19844 VDD.n2756 VDD.n2755 185
R19845 VDD.n2755 VDD.n656 185
R19846 VDD.n2757 VDD.n663 185
R19847 VDD.n3060 VDD.n663 185
R19848 VDD.n2759 VDD.n2758 185
R19849 VDD.n2758 VDD.n662 185
R19850 VDD.n2760 VDD.n669 185
R19851 VDD.n3054 VDD.n669 185
R19852 VDD.n2762 VDD.n2761 185
R19853 VDD.n2761 VDD.n668 185
R19854 VDD.n2763 VDD.n674 185
R19855 VDD.n3048 VDD.n674 185
R19856 VDD.n2765 VDD.n2764 185
R19857 VDD.n2764 VDD.n682 185
R19858 VDD.n2766 VDD.n680 185
R19859 VDD.n3042 VDD.n680 185
R19860 VDD.n2768 VDD.n2767 185
R19861 VDD.n2767 VDD.n679 185
R19862 VDD.n2769 VDD.n687 185
R19863 VDD.n3036 VDD.n687 185
R19864 VDD.n2771 VDD.n2770 185
R19865 VDD.n2770 VDD.n686 185
R19866 VDD.n2772 VDD.n693 185
R19867 VDD.n3030 VDD.n693 185
R19868 VDD.n2774 VDD.n2773 185
R19869 VDD.n2773 VDD.n692 185
R19870 VDD.n2775 VDD.n699 185
R19871 VDD.n3024 VDD.n699 185
R19872 VDD.n2777 VDD.n2776 185
R19873 VDD.n2776 VDD.n698 185
R19874 VDD.n2778 VDD.n705 185
R19875 VDD.n3018 VDD.n705 185
R19876 VDD.n2779 VDD.n2560 185
R19877 VDD.n2560 VDD.n704 185
R19878 VDD.n2781 VDD.n2780 185
R19879 VDD.n3012 VDD.n2781 185
R19880 VDD.n3014 VDD.n3013 185
R19881 VDD.n3013 VDD.n3012 185
R19882 VDD.n3015 VDD.n707 185
R19883 VDD.n707 VDD.n704 185
R19884 VDD.n3017 VDD.n3016 185
R19885 VDD.n3018 VDD.n3017 185
R19886 VDD.n697 VDD.n696 185
R19887 VDD.n698 VDD.n697 185
R19888 VDD.n3026 VDD.n3025 185
R19889 VDD.n3025 VDD.n3024 185
R19890 VDD.n3027 VDD.n695 185
R19891 VDD.n695 VDD.n692 185
R19892 VDD.n3029 VDD.n3028 185
R19893 VDD.n3030 VDD.n3029 185
R19894 VDD.n685 VDD.n684 185
R19895 VDD.n686 VDD.n685 185
R19896 VDD.n3038 VDD.n3037 185
R19897 VDD.n3037 VDD.n3036 185
R19898 VDD.n3039 VDD.n683 185
R19899 VDD.n683 VDD.n679 185
R19900 VDD.n3041 VDD.n3040 185
R19901 VDD.n3042 VDD.n3041 185
R19902 VDD.n673 VDD.n672 185
R19903 VDD.n682 VDD.n673 185
R19904 VDD.n3050 VDD.n3049 185
R19905 VDD.n3049 VDD.n3048 185
R19906 VDD.n3051 VDD.n671 185
R19907 VDD.n671 VDD.n668 185
R19908 VDD.n3053 VDD.n3052 185
R19909 VDD.n3054 VDD.n3053 185
R19910 VDD.n661 VDD.n660 185
R19911 VDD.n662 VDD.n661 185
R19912 VDD.n3062 VDD.n3061 185
R19913 VDD.n3061 VDD.n3060 185
R19914 VDD.n3063 VDD.n659 185
R19915 VDD.n659 VDD.n656 185
R19916 VDD.n3065 VDD.n3064 185
R19917 VDD.n3066 VDD.n3065 185
R19918 VDD.n649 VDD.n648 185
R19919 VDD.n650 VDD.n649 185
R19920 VDD.n3074 VDD.n3073 185
R19921 VDD.n3073 VDD.n3072 185
R19922 VDD.n3075 VDD.n647 185
R19923 VDD.n647 VDD.n644 185
R19924 VDD.n3077 VDD.n3076 185
R19925 VDD.n3078 VDD.n3077 185
R19926 VDD.n637 VDD.n636 185
R19927 VDD.n638 VDD.n637 185
R19928 VDD.n3086 VDD.n3085 185
R19929 VDD.n3085 VDD.n3084 185
R19930 VDD.n3087 VDD.n635 185
R19931 VDD.n635 VDD.n632 185
R19932 VDD.n3089 VDD.n3088 185
R19933 VDD.n3090 VDD.n3089 185
R19934 VDD.n625 VDD.n624 185
R19935 VDD.n626 VDD.n625 185
R19936 VDD.n3098 VDD.n3097 185
R19937 VDD.n3097 VDD.n3096 185
R19938 VDD.n3099 VDD.n623 185
R19939 VDD.n623 VDD.n619 185
R19940 VDD.n3101 VDD.n3100 185
R19941 VDD.n3102 VDD.n3101 185
R19942 VDD.n613 VDD.n612 185
R19943 VDD.n622 VDD.n613 185
R19944 VDD.n3110 VDD.n3109 185
R19945 VDD.n3109 VDD.n3108 185
R19946 VDD.n3111 VDD.n611 185
R19947 VDD.n611 VDD.n608 185
R19948 VDD.n3113 VDD.n3112 185
R19949 VDD.n3114 VDD.n3113 185
R19950 VDD.n601 VDD.n600 185
R19951 VDD.n602 VDD.n601 185
R19952 VDD.n3122 VDD.n3121 185
R19953 VDD.n3121 VDD.n3120 185
R19954 VDD.n3123 VDD.n599 185
R19955 VDD.n599 VDD.n596 185
R19956 VDD.n3125 VDD.n3124 185
R19957 VDD.n3126 VDD.n3125 185
R19958 VDD.n589 VDD.n588 185
R19959 VDD.n590 VDD.n589 185
R19960 VDD.n3134 VDD.n3133 185
R19961 VDD.n3133 VDD.n3132 185
R19962 VDD.n3135 VDD.n587 185
R19963 VDD.n587 VDD.n584 185
R19964 VDD.n3137 VDD.n3136 185
R19965 VDD.n3138 VDD.n3137 185
R19966 VDD.n577 VDD.n576 185
R19967 VDD.n578 VDD.n577 185
R19968 VDD.n3146 VDD.n3145 185
R19969 VDD.n3145 VDD.n3144 185
R19970 VDD.n3147 VDD.n575 185
R19971 VDD.n575 VDD.n572 185
R19972 VDD.n3149 VDD.n3148 185
R19973 VDD.n3150 VDD.n3149 185
R19974 VDD.n565 VDD.n564 185
R19975 VDD.n566 VDD.n565 185
R19976 VDD.n3158 VDD.n3157 185
R19977 VDD.n3157 VDD.n3156 185
R19978 VDD.n3159 VDD.n563 185
R19979 VDD.n563 VDD.n560 185
R19980 VDD.n3161 VDD.n3160 185
R19981 VDD.n3162 VDD.n3161 185
R19982 VDD.n552 VDD.n551 185
R19983 VDD.n553 VDD.n552 185
R19984 VDD.n3170 VDD.n3169 185
R19985 VDD.n3169 VDD.n3168 185
R19986 VDD.n3171 VDD.n550 185
R19987 VDD.n556 VDD.n550 185
R19988 VDD.n3173 VDD.n3172 185
R19989 VDD.n3174 VDD.n3173 185
R19990 VDD.n541 VDD.n540 185
R19991 VDD.n542 VDD.n541 185
R19992 VDD.n3182 VDD.n3181 185
R19993 VDD.n3181 VDD.n3180 185
R19994 VDD.n3183 VDD.n539 185
R19995 VDD.n539 VDD.n536 185
R19996 VDD.n3185 VDD.n3184 185
R19997 VDD.n3186 VDD.n3185 185
R19998 VDD.n529 VDD.n528 185
R19999 VDD.n530 VDD.n529 185
R20000 VDD.n3194 VDD.n3193 185
R20001 VDD.n3193 VDD.n3192 185
R20002 VDD.n3195 VDD.n527 185
R20003 VDD.n527 VDD.n524 185
R20004 VDD.n3197 VDD.n3196 185
R20005 VDD.n3198 VDD.n3197 185
R20006 VDD.n517 VDD.n516 185
R20007 VDD.n518 VDD.n517 185
R20008 VDD.n3206 VDD.n3205 185
R20009 VDD.n3205 VDD.n3204 185
R20010 VDD.n3207 VDD.n515 185
R20011 VDD.n515 VDD.n512 185
R20012 VDD.n3209 VDD.n3208 185
R20013 VDD.n3210 VDD.n3209 185
R20014 VDD.n504 VDD.n503 185
R20015 VDD.n505 VDD.n504 185
R20016 VDD.n3218 VDD.n3217 185
R20017 VDD.n3217 VDD.n3216 185
R20018 VDD.n3219 VDD.n502 185
R20019 VDD.n508 VDD.n502 185
R20020 VDD.n3221 VDD.n3220 185
R20021 VDD.n3222 VDD.n3221 185
R20022 VDD.n493 VDD.n492 185
R20023 VDD.n501 VDD.n493 185
R20024 VDD.n3230 VDD.n3229 185
R20025 VDD.n3229 VDD.n3228 185
R20026 VDD.n3231 VDD.n491 185
R20027 VDD.n491 VDD.n488 185
R20028 VDD.n3233 VDD.n3232 185
R20029 VDD.n3234 VDD.n3233 185
R20030 VDD.n481 VDD.n480 185
R20031 VDD.n482 VDD.n481 185
R20032 VDD.n3242 VDD.n3241 185
R20033 VDD.n3241 VDD.n3240 185
R20034 VDD.n3243 VDD.n479 185
R20035 VDD.n479 VDD.n476 185
R20036 VDD.n3245 VDD.n3244 185
R20037 VDD.n3246 VDD.n3245 185
R20038 VDD.n469 VDD.n468 185
R20039 VDD.n470 VDD.n469 185
R20040 VDD.n3254 VDD.n3253 185
R20041 VDD.n3253 VDD.n3252 185
R20042 VDD.n3255 VDD.n467 185
R20043 VDD.n467 VDD.n464 185
R20044 VDD.n3257 VDD.n3256 185
R20045 VDD.n3258 VDD.n3257 185
R20046 VDD.n457 VDD.n456 185
R20047 VDD.n458 VDD.n457 185
R20048 VDD.n3266 VDD.n3265 185
R20049 VDD.n3265 VDD.n3264 185
R20050 VDD.n3267 VDD.n455 185
R20051 VDD.n455 VDD.n452 185
R20052 VDD.n3269 VDD.n3268 185
R20053 VDD.n3270 VDD.n3269 185
R20054 VDD.n445 VDD.n444 185
R20055 VDD.n446 VDD.n445 185
R20056 VDD.n3278 VDD.n3277 185
R20057 VDD.n3277 VDD.n3276 185
R20058 VDD.n3279 VDD.n443 185
R20059 VDD.n443 VDD.n440 185
R20060 VDD.n3281 VDD.n3280 185
R20061 VDD.n3282 VDD.n3281 185
R20062 VDD.n433 VDD.n432 185
R20063 VDD.n434 VDD.n433 185
R20064 VDD.n3290 VDD.n3289 185
R20065 VDD.n3289 VDD.n3288 185
R20066 VDD.n3291 VDD.n431 185
R20067 VDD.n431 VDD.n428 185
R20068 VDD.n3293 VDD.n3292 185
R20069 VDD.n3294 VDD.n3293 185
R20070 VDD.n420 VDD.n419 185
R20071 VDD.n421 VDD.n420 185
R20072 VDD.n3302 VDD.n3301 185
R20073 VDD.n3301 VDD.n3300 185
R20074 VDD.n3303 VDD.n418 185
R20075 VDD.n424 VDD.n418 185
R20076 VDD.n3305 VDD.n3304 185
R20077 VDD.n3306 VDD.n3305 185
R20078 VDD.n409 VDD.n408 185
R20079 VDD.n410 VDD.n409 185
R20080 VDD.n3314 VDD.n3313 185
R20081 VDD.n3313 VDD.n3312 185
R20082 VDD.n3315 VDD.n407 185
R20083 VDD.n407 VDD.n404 185
R20084 VDD.n3317 VDD.n3316 185
R20085 VDD.n3318 VDD.n3317 185
R20086 VDD.n397 VDD.n396 185
R20087 VDD.n398 VDD.n397 185
R20088 VDD.n3326 VDD.n3325 185
R20089 VDD.n3325 VDD.n3324 185
R20090 VDD.n3327 VDD.n395 185
R20091 VDD.n395 VDD.n392 185
R20092 VDD.n3329 VDD.n3328 185
R20093 VDD.n3330 VDD.n3329 185
R20094 VDD.n385 VDD.n384 185
R20095 VDD.n386 VDD.n385 185
R20096 VDD.n3338 VDD.n3337 185
R20097 VDD.n3337 VDD.n3336 185
R20098 VDD.n3339 VDD.n383 185
R20099 VDD.n383 VDD.n380 185
R20100 VDD.n3341 VDD.n3340 185
R20101 VDD.n3342 VDD.n3341 185
R20102 VDD.n372 VDD.n371 185
R20103 VDD.n373 VDD.n372 185
R20104 VDD.n3350 VDD.n3349 185
R20105 VDD.n3349 VDD.n3348 185
R20106 VDD.n3351 VDD.n370 185
R20107 VDD.n376 VDD.n370 185
R20108 VDD.n3353 VDD.n3352 185
R20109 VDD.n3354 VDD.n3353 185
R20110 VDD.n361 VDD.n360 185
R20111 VDD.n362 VDD.n361 185
R20112 VDD.n3362 VDD.n3361 185
R20113 VDD.n3361 VDD.n3360 185
R20114 VDD.n3363 VDD.n359 185
R20115 VDD.n359 VDD.n356 185
R20116 VDD.n3365 VDD.n3364 185
R20117 VDD.n3366 VDD.n3365 185
R20118 VDD.n348 VDD.n347 185
R20119 VDD.n349 VDD.n348 185
R20120 VDD.n3399 VDD.n3398 185
R20121 VDD.n3398 VDD.n3397 185
R20122 VDD.n3400 VDD.n346 185
R20123 VDD.n346 VDD.n343 185
R20124 VDD.n3402 VDD.n3401 185
R20125 VDD.n3403 VDD.n3402 185
R20126 VDD.n327 VDD.n325 185
R20127 VDD.n325 VDD.n321 185
R20128 VDD.n3442 VDD.n3441 185
R20129 VDD.n3443 VDD.n3442 185
R20130 VDD.n3440 VDD.n326 185
R20131 VDD.n326 VDD.n323 185
R20132 VDD.n1674 VDD.n1673 185
R20133 VDD.n1675 VDD.n1181 185
R20134 VDD.n1669 VDD.n1177 185
R20135 VDD.n1679 VDD.n1176 185
R20136 VDD.n1680 VDD.n1175 185
R20137 VDD.n1681 VDD.n1174 185
R20138 VDD.n1666 VDD.n1172 185
R20139 VDD.n1685 VDD.n1171 185
R20140 VDD.n1686 VDD.n1170 185
R20141 VDD.n1687 VDD.n1169 185
R20142 VDD.n1663 VDD.n1167 185
R20143 VDD.n1691 VDD.n1166 185
R20144 VDD.n1692 VDD.n1165 185
R20145 VDD.n1693 VDD.n1164 185
R20146 VDD.n1660 VDD.n1163 185
R20147 VDD.n1659 VDD.n1658 185
R20148 VDD.n1191 VDD.n1190 185
R20149 VDD.n1654 VDD.n1653 185
R20150 VDD.n1652 VDD.n1651 185
R20151 VDD.n1650 VDD.n1197 185
R20152 VDD.n1196 VDD.n1195 185
R20153 VDD.n1646 VDD.n1645 185
R20154 VDD.n1644 VDD.n1643 185
R20155 VDD.n1642 VDD.n1201 185
R20156 VDD.n1200 VDD.n1199 185
R20157 VDD.n1638 VDD.n1637 185
R20158 VDD.n1636 VDD.n1635 185
R20159 VDD.n1634 VDD.n1632 185
R20160 VDD.n1211 VDD.n1182 185
R20161 VDD.n1183 VDD.n1182 185
R20162 VDD.n1622 VDD.n1621 185
R20163 VDD.n1623 VDD.n1622 185
R20164 VDD.n1210 VDD.n1209 185
R20165 VDD.n1624 VDD.n1209 185
R20166 VDD.n1614 VDD.n1613 185
R20167 VDD.n1613 VDD.n1208 185
R20168 VDD.n1612 VDD.n1213 185
R20169 VDD.n1612 VDD.n1611 185
R20170 VDD.n1224 VDD.n1214 185
R20171 VDD.n1215 VDD.n1214 185
R20172 VDD.n1602 VDD.n1601 185
R20173 VDD.n1603 VDD.n1602 185
R20174 VDD.n1223 VDD.n1222 185
R20175 VDD.n1222 VDD.n1221 185
R20176 VDD.n1596 VDD.n1595 185
R20177 VDD.n1595 VDD.n1594 185
R20178 VDD.n1227 VDD.n1226 185
R20179 VDD.n1228 VDD.n1227 185
R20180 VDD.n1585 VDD.n1584 185
R20181 VDD.n1586 VDD.n1585 185
R20182 VDD.n1236 VDD.n1235 185
R20183 VDD.n1235 VDD.n1234 185
R20184 VDD.n1580 VDD.n1579 185
R20185 VDD.n1579 VDD.n1578 185
R20186 VDD.n1239 VDD.n1238 185
R20187 VDD.n1240 VDD.n1239 185
R20188 VDD.n1569 VDD.n1568 185
R20189 VDD.n1570 VDD.n1569 185
R20190 VDD.n1248 VDD.n1247 185
R20191 VDD.n1247 VDD.n1246 185
R20192 VDD.n1564 VDD.n1563 185
R20193 VDD.n1563 VDD.n1562 185
R20194 VDD.n1251 VDD.n1250 185
R20195 VDD.n1252 VDD.n1251 185
R20196 VDD.n1553 VDD.n1552 185
R20197 VDD.n1554 VDD.n1553 185
R20198 VDD.n1260 VDD.n1259 185
R20199 VDD.n1259 VDD.n1258 185
R20200 VDD.n1548 VDD.n1547 185
R20201 VDD.n1547 VDD.n1546 185
R20202 VDD.n1263 VDD.n1262 185
R20203 VDD.n1264 VDD.n1263 185
R20204 VDD.n1537 VDD.n1536 185
R20205 VDD.n1538 VDD.n1537 185
R20206 VDD.n1276 VDD.n1275 185
R20207 VDD.n1275 VDD.n1274 185
R20208 VDD.n1532 VDD.n1531 185
R20209 VDD.n1531 VDD.n1530 185
R20210 VDD.n1279 VDD.n1278 185
R20211 VDD.n1280 VDD.n1279 185
R20212 VDD.n1520 VDD.n1519 185
R20213 VDD.n1521 VDD.n1520 185
R20214 VDD.n1288 VDD.n1287 185
R20215 VDD.n1287 VDD.n1286 185
R20216 VDD.n1515 VDD.n1514 185
R20217 VDD.n1514 VDD.n1513 185
R20218 VDD.n1291 VDD.n1290 185
R20219 VDD.n1292 VDD.n1291 185
R20220 VDD.n1504 VDD.n1503 185
R20221 VDD.n1505 VDD.n1504 185
R20222 VDD.n1300 VDD.n1299 185
R20223 VDD.n1299 VDD.n1298 185
R20224 VDD.n1499 VDD.n1498 185
R20225 VDD.n1498 VDD.n1497 185
R20226 VDD.n1303 VDD.n1302 185
R20227 VDD.n1304 VDD.n1303 185
R20228 VDD.n1488 VDD.n1487 185
R20229 VDD.n1489 VDD.n1488 185
R20230 VDD.n1312 VDD.n1311 185
R20231 VDD.n1311 VDD.n1310 185
R20232 VDD.n1483 VDD.n1482 185
R20233 VDD.n1482 VDD.n1481 185
R20234 VDD.n1315 VDD.n1314 185
R20235 VDD.n1316 VDD.n1315 185
R20236 VDD.n1472 VDD.n1471 185
R20237 VDD.n1473 VDD.n1472 185
R20238 VDD.n1324 VDD.n1323 185
R20239 VDD.n1323 VDD.n1322 185
R20240 VDD.n1467 VDD.n1466 185
R20241 VDD.n1466 VDD.n1465 185
R20242 VDD.n1327 VDD.n1326 185
R20243 VDD.n1328 VDD.n1327 185
R20244 VDD.n1456 VDD.n1455 185
R20245 VDD.n1457 VDD.n1456 185
R20246 VDD.n1336 VDD.n1335 185
R20247 VDD.n1335 VDD.n1334 185
R20248 VDD.n1451 VDD.n1450 185
R20249 VDD.n1450 VDD.n1449 185
R20250 VDD.n1339 VDD.n1338 185
R20251 VDD.n1340 VDD.n1339 185
R20252 VDD.n1443 VDD.n1442 185
R20253 VDD.n1345 VDD.n1344 185
R20254 VDD.n1439 VDD.n1438 185
R20255 VDD.n1440 VDD.n1439 185
R20256 VDD.n1360 VDD.n1359 185
R20257 VDD.n1434 VDD.n1362 185
R20258 VDD.n1433 VDD.n1363 185
R20259 VDD.n1432 VDD.n1364 185
R20260 VDD.n1366 VDD.n1365 185
R20261 VDD.n1428 VDD.n1368 185
R20262 VDD.n1427 VDD.n1369 185
R20263 VDD.n1426 VDD.n1370 185
R20264 VDD.n1372 VDD.n1371 185
R20265 VDD.n1422 VDD.n1419 185
R20266 VDD.n1418 VDD.n1417 185
R20267 VDD.n1416 VDD.n1374 185
R20268 VDD.n1376 VDD.n1375 185
R20269 VDD.n1412 VDD.n1378 185
R20270 VDD.n1411 VDD.n1379 185
R20271 VDD.n1410 VDD.n1380 185
R20272 VDD.n1382 VDD.n1381 185
R20273 VDD.n1406 VDD.n1384 185
R20274 VDD.n1405 VDD.n1385 185
R20275 VDD.n1404 VDD.n1386 185
R20276 VDD.n1388 VDD.n1387 185
R20277 VDD.n1400 VDD.n1390 185
R20278 VDD.n1399 VDD.n1391 185
R20279 VDD.n1398 VDD.n1395 185
R20280 VDD.n1392 VDD.n1358 185
R20281 VDD.n1440 VDD.n1358 185
R20282 VDD.n1631 VDD.n1630 185
R20283 VDD.n1631 VDD.n1183 185
R20284 VDD.n1204 VDD.n1203 185
R20285 VDD.n1623 VDD.n1203 185
R20286 VDD.n1626 VDD.n1625 185
R20287 VDD.n1625 VDD.n1624 185
R20288 VDD.n1207 VDD.n1206 185
R20289 VDD.n1208 VDD.n1207 185
R20290 VDD.n1610 VDD.n1609 185
R20291 VDD.n1611 VDD.n1610 185
R20292 VDD.n1217 VDD.n1216 185
R20293 VDD.n1216 VDD.n1215 185
R20294 VDD.n1605 VDD.n1604 185
R20295 VDD.n1604 VDD.n1603 185
R20296 VDD.n1220 VDD.n1219 185
R20297 VDD.n1221 VDD.n1220 185
R20298 VDD.n1593 VDD.n1592 185
R20299 VDD.n1594 VDD.n1593 185
R20300 VDD.n1230 VDD.n1229 185
R20301 VDD.n1229 VDD.n1228 185
R20302 VDD.n1588 VDD.n1587 185
R20303 VDD.n1587 VDD.n1586 185
R20304 VDD.n1233 VDD.n1232 185
R20305 VDD.n1234 VDD.n1233 185
R20306 VDD.n1577 VDD.n1576 185
R20307 VDD.n1578 VDD.n1577 185
R20308 VDD.n1242 VDD.n1241 185
R20309 VDD.n1241 VDD.n1240 185
R20310 VDD.n1572 VDD.n1571 185
R20311 VDD.n1571 VDD.n1570 185
R20312 VDD.n1245 VDD.n1244 185
R20313 VDD.n1246 VDD.n1245 185
R20314 VDD.n1561 VDD.n1560 185
R20315 VDD.n1562 VDD.n1561 185
R20316 VDD.n1254 VDD.n1253 185
R20317 VDD.n1253 VDD.n1252 185
R20318 VDD.n1556 VDD.n1555 185
R20319 VDD.n1555 VDD.n1554 185
R20320 VDD.n1257 VDD.n1256 185
R20321 VDD.n1258 VDD.n1257 185
R20322 VDD.n1545 VDD.n1544 185
R20323 VDD.n1546 VDD.n1545 185
R20324 VDD.n1266 VDD.n1265 185
R20325 VDD.n1265 VDD.n1264 185
R20326 VDD.n1540 VDD.n1539 185
R20327 VDD.n1539 VDD.n1538 185
R20328 VDD.n1273 VDD.n1272 185
R20329 VDD.n1274 VDD.n1273 185
R20330 VDD.n1529 VDD.n1528 185
R20331 VDD.n1530 VDD.n1529 185
R20332 VDD.n1282 VDD.n1281 185
R20333 VDD.n1281 VDD.n1280 185
R20334 VDD.n1523 VDD.n1522 185
R20335 VDD.n1522 VDD.n1521 185
R20336 VDD.n1285 VDD.n1284 185
R20337 VDD.n1286 VDD.n1285 185
R20338 VDD.n1512 VDD.n1511 185
R20339 VDD.n1513 VDD.n1512 185
R20340 VDD.n1294 VDD.n1293 185
R20341 VDD.n1293 VDD.n1292 185
R20342 VDD.n1507 VDD.n1506 185
R20343 VDD.n1506 VDD.n1505 185
R20344 VDD.n1297 VDD.n1296 185
R20345 VDD.n1298 VDD.n1297 185
R20346 VDD.n1496 VDD.n1495 185
R20347 VDD.n1497 VDD.n1496 185
R20348 VDD.n1306 VDD.n1305 185
R20349 VDD.n1305 VDD.n1304 185
R20350 VDD.n1491 VDD.n1490 185
R20351 VDD.n1490 VDD.n1489 185
R20352 VDD.n1309 VDD.n1308 185
R20353 VDD.n1310 VDD.n1309 185
R20354 VDD.n1480 VDD.n1479 185
R20355 VDD.n1481 VDD.n1480 185
R20356 VDD.n1318 VDD.n1317 185
R20357 VDD.n1317 VDD.n1316 185
R20358 VDD.n1475 VDD.n1474 185
R20359 VDD.n1474 VDD.n1473 185
R20360 VDD.n1321 VDD.n1320 185
R20361 VDD.n1322 VDD.n1321 185
R20362 VDD.n1464 VDD.n1463 185
R20363 VDD.n1465 VDD.n1464 185
R20364 VDD.n1330 VDD.n1329 185
R20365 VDD.n1329 VDD.n1328 185
R20366 VDD.n1459 VDD.n1458 185
R20367 VDD.n1458 VDD.n1457 185
R20368 VDD.n1333 VDD.n1332 185
R20369 VDD.n1334 VDD.n1333 185
R20370 VDD.n1448 VDD.n1447 185
R20371 VDD.n1449 VDD.n1448 185
R20372 VDD.n1342 VDD.n1341 185
R20373 VDD.n1341 VDD.n1340 185
R20374 VDD.n2791 VDD.t34 171.01
R20375 VDD.n336 VDD.t23 171.01
R20376 VDD.n2589 VDD.t47 171.01
R20377 VDD.n315 VDD.t42 171.01
R20378 VDD.n1120 VDD.t66 171.01
R20379 VDD.n1138 VDD.t26 171.01
R20380 VDD.n738 VDD.t61 171.01
R20381 VDD.n2463 VDD.t19 171.01
R20382 VDD.n9 VDD.n7 168.903
R20383 VDD.n2 VDD.n0 168.903
R20384 VDD.n9 VDD.n8 167.054
R20385 VDD.n11 VDD.n10 167.054
R20386 VDD.n13 VDD.n12 167.054
R20387 VDD.n6 VDD.n5 167.054
R20388 VDD.n4 VDD.n3 167.054
R20389 VDD.n2 VDD.n1 167.054
R20390 VDD.n120 VDD.n119 146.341
R20391 VDD.n127 VDD.n126 146.341
R20392 VDD.n130 VDD.n129 146.341
R20393 VDD.n137 VDD.n136 146.341
R20394 VDD.n140 VDD.n139 146.341
R20395 VDD.n145 VDD.n109 146.341
R20396 VDD.n149 VDD.n148 146.341
R20397 VDD.n156 VDD.n155 146.341
R20398 VDD.n159 VDD.n158 146.341
R20399 VDD.n166 VDD.n165 146.341
R20400 VDD.n169 VDD.n168 146.341
R20401 VDD.n176 VDD.n175 146.341
R20402 VDD.n178 VDD.n96 146.341
R20403 VDD.n3530 VDD.n255 146.341
R20404 VDD.n3530 VDD.n251 146.341
R20405 VDD.n3536 VDD.n251 146.341
R20406 VDD.n3536 VDD.n243 146.341
R20407 VDD.n3546 VDD.n243 146.341
R20408 VDD.n3546 VDD.n239 146.341
R20409 VDD.n3552 VDD.n239 146.341
R20410 VDD.n3552 VDD.n231 146.341
R20411 VDD.n3562 VDD.n231 146.341
R20412 VDD.n3562 VDD.n227 146.341
R20413 VDD.n3568 VDD.n227 146.341
R20414 VDD.n3568 VDD.n219 146.341
R20415 VDD.n3578 VDD.n219 146.341
R20416 VDD.n3578 VDD.n215 146.341
R20417 VDD.n3586 VDD.n215 146.341
R20418 VDD.n3586 VDD.n207 146.341
R20419 VDD.n3596 VDD.n207 146.341
R20420 VDD.n3597 VDD.n3596 146.341
R20421 VDD.n3597 VDD.n203 146.341
R20422 VDD.n3606 VDD.n203 146.341
R20423 VDD.n3606 VDD.n195 146.341
R20424 VDD.n3618 VDD.n195 146.341
R20425 VDD.n3619 VDD.n3618 146.341
R20426 VDD.n3619 VDD.n26 146.341
R20427 VDD.n27 VDD.n26 146.341
R20428 VDD.n28 VDD.n27 146.341
R20429 VDD.n3626 VDD.n28 146.341
R20430 VDD.n3626 VDD.n37 146.341
R20431 VDD.n38 VDD.n37 146.341
R20432 VDD.n39 VDD.n38 146.341
R20433 VDD.n3633 VDD.n39 146.341
R20434 VDD.n3633 VDD.n48 146.341
R20435 VDD.n49 VDD.n48 146.341
R20436 VDD.n50 VDD.n49 146.341
R20437 VDD.n3640 VDD.n50 146.341
R20438 VDD.n3640 VDD.n59 146.341
R20439 VDD.n60 VDD.n59 146.341
R20440 VDD.n61 VDD.n60 146.341
R20441 VDD.n3647 VDD.n61 146.341
R20442 VDD.n3647 VDD.n70 146.341
R20443 VDD.n71 VDD.n70 146.341
R20444 VDD.n72 VDD.n71 146.341
R20445 VDD.n3654 VDD.n72 146.341
R20446 VDD.n3654 VDD.n81 146.341
R20447 VDD.n82 VDD.n81 146.341
R20448 VDD.n3517 VDD.n263 146.341
R20449 VDD.n3517 VDD.n277 146.341
R20450 VDD.n3513 VDD.n3512 146.341
R20451 VDD.n3509 VDD.n3508 146.341
R20452 VDD.n3505 VDD.n3504 146.341
R20453 VDD.n3501 VDD.n3500 146.341
R20454 VDD.n3496 VDD.n288 146.341
R20455 VDD.n3494 VDD.n3493 146.341
R20456 VDD.n3490 VDD.n3489 146.341
R20457 VDD.n3486 VDD.n3485 146.341
R20458 VDD.n3482 VDD.n3481 146.341
R20459 VDD.n3478 VDD.n3477 146.341
R20460 VDD.n3474 VDD.n3473 146.341
R20461 VDD.n304 VDD.n276 146.341
R20462 VDD.n3528 VDD.n257 146.341
R20463 VDD.n3528 VDD.n249 146.341
R20464 VDD.n3538 VDD.n249 146.341
R20465 VDD.n3538 VDD.n245 146.341
R20466 VDD.n3544 VDD.n245 146.341
R20467 VDD.n3544 VDD.n237 146.341
R20468 VDD.n3554 VDD.n237 146.341
R20469 VDD.n3554 VDD.n233 146.341
R20470 VDD.n3560 VDD.n233 146.341
R20471 VDD.n3560 VDD.n225 146.341
R20472 VDD.n3570 VDD.n225 146.341
R20473 VDD.n3570 VDD.n221 146.341
R20474 VDD.n3576 VDD.n221 146.341
R20475 VDD.n3576 VDD.n213 146.341
R20476 VDD.n3588 VDD.n213 146.341
R20477 VDD.n3588 VDD.n209 146.341
R20478 VDD.n3594 VDD.n209 146.341
R20479 VDD.n3594 VDD.n201 146.341
R20480 VDD.n3609 VDD.n201 146.341
R20481 VDD.n3609 VDD.n197 146.341
R20482 VDD.n3615 VDD.n197 146.341
R20483 VDD.n3616 VDD.n3615 146.341
R20484 VDD.n3616 VDD.n22 146.341
R20485 VDD.n3706 VDD.n22 146.341
R20486 VDD.n3706 VDD.n24 146.341
R20487 VDD.n3702 VDD.n24 146.341
R20488 VDD.n3702 VDD.n30 146.341
R20489 VDD.n3698 VDD.n30 146.341
R20490 VDD.n3698 VDD.n36 146.341
R20491 VDD.n3694 VDD.n36 146.341
R20492 VDD.n3694 VDD.n41 146.341
R20493 VDD.n3690 VDD.n41 146.341
R20494 VDD.n3690 VDD.n47 146.341
R20495 VDD.n3686 VDD.n47 146.341
R20496 VDD.n3686 VDD.n52 146.341
R20497 VDD.n3682 VDD.n52 146.341
R20498 VDD.n3682 VDD.n58 146.341
R20499 VDD.n3678 VDD.n58 146.341
R20500 VDD.n3678 VDD.n63 146.341
R20501 VDD.n3674 VDD.n63 146.341
R20502 VDD.n3674 VDD.n69 146.341
R20503 VDD.n3670 VDD.n69 146.341
R20504 VDD.n3670 VDD.n74 146.341
R20505 VDD.n3666 VDD.n74 146.341
R20506 VDD.n3666 VDD.n80 146.341
R20507 VDD.n1637 VDD.n1636 146.341
R20508 VDD.n1201 VDD.n1200 146.341
R20509 VDD.n1645 VDD.n1644 146.341
R20510 VDD.n1197 VDD.n1196 146.341
R20511 VDD.n1653 VDD.n1652 146.341
R20512 VDD.n1659 VDD.n1190 146.341
R20513 VDD.n1660 VDD.n1164 146.341
R20514 VDD.n1166 VDD.n1165 146.341
R20515 VDD.n1663 VDD.n1169 146.341
R20516 VDD.n1171 VDD.n1170 146.341
R20517 VDD.n1666 VDD.n1174 146.341
R20518 VDD.n1176 VDD.n1175 146.341
R20519 VDD.n1669 VDD.n1181 146.341
R20520 VDD.n1450 VDD.n1339 146.341
R20521 VDD.n1450 VDD.n1335 146.341
R20522 VDD.n1456 VDD.n1335 146.341
R20523 VDD.n1456 VDD.n1327 146.341
R20524 VDD.n1466 VDD.n1327 146.341
R20525 VDD.n1466 VDD.n1323 146.341
R20526 VDD.n1472 VDD.n1323 146.341
R20527 VDD.n1472 VDD.n1315 146.341
R20528 VDD.n1482 VDD.n1315 146.341
R20529 VDD.n1482 VDD.n1311 146.341
R20530 VDD.n1488 VDD.n1311 146.341
R20531 VDD.n1488 VDD.n1303 146.341
R20532 VDD.n1498 VDD.n1303 146.341
R20533 VDD.n1498 VDD.n1299 146.341
R20534 VDD.n1504 VDD.n1299 146.341
R20535 VDD.n1504 VDD.n1291 146.341
R20536 VDD.n1514 VDD.n1291 146.341
R20537 VDD.n1514 VDD.n1287 146.341
R20538 VDD.n1520 VDD.n1287 146.341
R20539 VDD.n1520 VDD.n1279 146.341
R20540 VDD.n1531 VDD.n1279 146.341
R20541 VDD.n1531 VDD.n1275 146.341
R20542 VDD.n1537 VDD.n1275 146.341
R20543 VDD.n1537 VDD.n1263 146.341
R20544 VDD.n1547 VDD.n1263 146.341
R20545 VDD.n1547 VDD.n1259 146.341
R20546 VDD.n1553 VDD.n1259 146.341
R20547 VDD.n1553 VDD.n1251 146.341
R20548 VDD.n1563 VDD.n1251 146.341
R20549 VDD.n1563 VDD.n1247 146.341
R20550 VDD.n1569 VDD.n1247 146.341
R20551 VDD.n1569 VDD.n1239 146.341
R20552 VDD.n1579 VDD.n1239 146.341
R20553 VDD.n1579 VDD.n1235 146.341
R20554 VDD.n1585 VDD.n1235 146.341
R20555 VDD.n1585 VDD.n1227 146.341
R20556 VDD.n1595 VDD.n1227 146.341
R20557 VDD.n1595 VDD.n1222 146.341
R20558 VDD.n1602 VDD.n1222 146.341
R20559 VDD.n1602 VDD.n1214 146.341
R20560 VDD.n1612 VDD.n1214 146.341
R20561 VDD.n1613 VDD.n1612 146.341
R20562 VDD.n1613 VDD.n1209 146.341
R20563 VDD.n1622 VDD.n1209 146.341
R20564 VDD.n1622 VDD.n1182 146.341
R20565 VDD.n1439 VDD.n1345 146.341
R20566 VDD.n1439 VDD.n1359 146.341
R20567 VDD.n1363 VDD.n1362 146.341
R20568 VDD.n1365 VDD.n1364 146.341
R20569 VDD.n1369 VDD.n1368 146.341
R20570 VDD.n1371 VDD.n1370 146.341
R20571 VDD.n1419 VDD.n1418 146.341
R20572 VDD.n1375 VDD.n1374 146.341
R20573 VDD.n1379 VDD.n1378 146.341
R20574 VDD.n1381 VDD.n1380 146.341
R20575 VDD.n1385 VDD.n1384 146.341
R20576 VDD.n1387 VDD.n1386 146.341
R20577 VDD.n1391 VDD.n1390 146.341
R20578 VDD.n1395 VDD.n1358 146.341
R20579 VDD.n1448 VDD.n1341 146.341
R20580 VDD.n1448 VDD.n1333 146.341
R20581 VDD.n1458 VDD.n1333 146.341
R20582 VDD.n1458 VDD.n1329 146.341
R20583 VDD.n1464 VDD.n1329 146.341
R20584 VDD.n1464 VDD.n1321 146.341
R20585 VDD.n1474 VDD.n1321 146.341
R20586 VDD.n1474 VDD.n1317 146.341
R20587 VDD.n1480 VDD.n1317 146.341
R20588 VDD.n1480 VDD.n1309 146.341
R20589 VDD.n1490 VDD.n1309 146.341
R20590 VDD.n1490 VDD.n1305 146.341
R20591 VDD.n1496 VDD.n1305 146.341
R20592 VDD.n1496 VDD.n1297 146.341
R20593 VDD.n1506 VDD.n1297 146.341
R20594 VDD.n1506 VDD.n1293 146.341
R20595 VDD.n1512 VDD.n1293 146.341
R20596 VDD.n1512 VDD.n1285 146.341
R20597 VDD.n1522 VDD.n1285 146.341
R20598 VDD.n1522 VDD.n1281 146.341
R20599 VDD.n1529 VDD.n1281 146.341
R20600 VDD.n1529 VDD.n1273 146.341
R20601 VDD.n1539 VDD.n1273 146.341
R20602 VDD.n1539 VDD.n1265 146.341
R20603 VDD.n1545 VDD.n1265 146.341
R20604 VDD.n1545 VDD.n1257 146.341
R20605 VDD.n1555 VDD.n1257 146.341
R20606 VDD.n1555 VDD.n1253 146.341
R20607 VDD.n1561 VDD.n1253 146.341
R20608 VDD.n1561 VDD.n1245 146.341
R20609 VDD.n1571 VDD.n1245 146.341
R20610 VDD.n1571 VDD.n1241 146.341
R20611 VDD.n1577 VDD.n1241 146.341
R20612 VDD.n1577 VDD.n1233 146.341
R20613 VDD.n1587 VDD.n1233 146.341
R20614 VDD.n1587 VDD.n1229 146.341
R20615 VDD.n1593 VDD.n1229 146.341
R20616 VDD.n1593 VDD.n1220 146.341
R20617 VDD.n1604 VDD.n1220 146.341
R20618 VDD.n1604 VDD.n1216 146.341
R20619 VDD.n1610 VDD.n1216 146.341
R20620 VDD.n1610 VDD.n1207 146.341
R20621 VDD.n1625 VDD.n1207 146.341
R20622 VDD.n1625 VDD.n1203 146.341
R20623 VDD.n1631 VDD.n1203 146.341
R20624 VDD.n2558 VDD.n2557 143.448
R20625 VDD.t76 VDD.n1108 113.219
R20626 VDD.n311 VDD.t102 113.219
R20627 VDD.n2791 VDD.n2790 111.903
R20628 VDD.n336 VDD.n335 111.903
R20629 VDD.n2589 VDD.n2588 111.903
R20630 VDD.n315 VDD.n314 111.903
R20631 VDD.n1120 VDD.n1119 111.903
R20632 VDD.n1138 VDD.n1137 111.903
R20633 VDD.n738 VDD.n737 111.903
R20634 VDD.n2463 VDD.n2462 111.903
R20635 VDD.n1397 VDD.t38 108.103
R20636 VDD.n1421 VDD.t54 108.103
R20637 VDD.n291 VDD.t63 108.103
R20638 VDD.n306 VDD.t51 108.103
R20639 VDD.n98 VDD.t58 108.103
R20640 VDD.n108 VDD.t15 108.103
R20641 VDD.n1193 VDD.t45 108.103
R20642 VDD.n1180 VDD.t31 108.103
R20643 VDD.n17 VDD.t7 107.823
R20644 VDD.n16 VDD.t2 107.823
R20645 VDD.n1268 VDD.t4 107.823
R20646 VDD.n1267 VDD.t10 107.823
R20647 VDD.n17 VDD.t11 106.451
R20648 VDD.n16 VDD.t9 106.451
R20649 VDD.n1268 VDD.t109 106.451
R20650 VDD.n1267 VDD.t6 106.451
R20651 VDD.n3013 VDD.n707 99.5127
R20652 VDD.n3017 VDD.n707 99.5127
R20653 VDD.n3017 VDD.n697 99.5127
R20654 VDD.n3025 VDD.n697 99.5127
R20655 VDD.n3025 VDD.n695 99.5127
R20656 VDD.n3029 VDD.n695 99.5127
R20657 VDD.n3029 VDD.n685 99.5127
R20658 VDD.n3037 VDD.n685 99.5127
R20659 VDD.n3037 VDD.n683 99.5127
R20660 VDD.n3041 VDD.n683 99.5127
R20661 VDD.n3041 VDD.n673 99.5127
R20662 VDD.n3049 VDD.n673 99.5127
R20663 VDD.n3049 VDD.n671 99.5127
R20664 VDD.n3053 VDD.n671 99.5127
R20665 VDD.n3053 VDD.n661 99.5127
R20666 VDD.n3061 VDD.n661 99.5127
R20667 VDD.n3061 VDD.n659 99.5127
R20668 VDD.n3065 VDD.n659 99.5127
R20669 VDD.n3065 VDD.n649 99.5127
R20670 VDD.n3073 VDD.n649 99.5127
R20671 VDD.n3073 VDD.n647 99.5127
R20672 VDD.n3077 VDD.n647 99.5127
R20673 VDD.n3077 VDD.n637 99.5127
R20674 VDD.n3085 VDD.n637 99.5127
R20675 VDD.n3085 VDD.n635 99.5127
R20676 VDD.n3089 VDD.n635 99.5127
R20677 VDD.n3089 VDD.n625 99.5127
R20678 VDD.n3097 VDD.n625 99.5127
R20679 VDD.n3097 VDD.n623 99.5127
R20680 VDD.n3101 VDD.n623 99.5127
R20681 VDD.n3101 VDD.n613 99.5127
R20682 VDD.n3109 VDD.n613 99.5127
R20683 VDD.n3109 VDD.n611 99.5127
R20684 VDD.n3113 VDD.n611 99.5127
R20685 VDD.n3113 VDD.n601 99.5127
R20686 VDD.n3121 VDD.n601 99.5127
R20687 VDD.n3121 VDD.n599 99.5127
R20688 VDD.n3125 VDD.n599 99.5127
R20689 VDD.n3125 VDD.n589 99.5127
R20690 VDD.n3133 VDD.n589 99.5127
R20691 VDD.n3133 VDD.n587 99.5127
R20692 VDD.n3137 VDD.n587 99.5127
R20693 VDD.n3137 VDD.n577 99.5127
R20694 VDD.n3145 VDD.n577 99.5127
R20695 VDD.n3145 VDD.n575 99.5127
R20696 VDD.n3149 VDD.n575 99.5127
R20697 VDD.n3149 VDD.n565 99.5127
R20698 VDD.n3157 VDD.n565 99.5127
R20699 VDD.n3157 VDD.n563 99.5127
R20700 VDD.n3161 VDD.n563 99.5127
R20701 VDD.n3161 VDD.n552 99.5127
R20702 VDD.n3169 VDD.n552 99.5127
R20703 VDD.n3169 VDD.n550 99.5127
R20704 VDD.n3173 VDD.n550 99.5127
R20705 VDD.n3173 VDD.n541 99.5127
R20706 VDD.n3181 VDD.n541 99.5127
R20707 VDD.n3181 VDD.n539 99.5127
R20708 VDD.n3185 VDD.n539 99.5127
R20709 VDD.n3185 VDD.n529 99.5127
R20710 VDD.n3193 VDD.n529 99.5127
R20711 VDD.n3193 VDD.n527 99.5127
R20712 VDD.n3197 VDD.n527 99.5127
R20713 VDD.n3197 VDD.n517 99.5127
R20714 VDD.n3205 VDD.n517 99.5127
R20715 VDD.n3205 VDD.n515 99.5127
R20716 VDD.n3209 VDD.n515 99.5127
R20717 VDD.n3209 VDD.n504 99.5127
R20718 VDD.n3217 VDD.n504 99.5127
R20719 VDD.n3217 VDD.n502 99.5127
R20720 VDD.n3221 VDD.n502 99.5127
R20721 VDD.n3221 VDD.n493 99.5127
R20722 VDD.n3229 VDD.n493 99.5127
R20723 VDD.n3229 VDD.n491 99.5127
R20724 VDD.n3233 VDD.n491 99.5127
R20725 VDD.n3233 VDD.n481 99.5127
R20726 VDD.n3241 VDD.n481 99.5127
R20727 VDD.n3241 VDD.n479 99.5127
R20728 VDD.n3245 VDD.n479 99.5127
R20729 VDD.n3245 VDD.n469 99.5127
R20730 VDD.n3253 VDD.n469 99.5127
R20731 VDD.n3253 VDD.n467 99.5127
R20732 VDD.n3257 VDD.n467 99.5127
R20733 VDD.n3257 VDD.n457 99.5127
R20734 VDD.n3265 VDD.n457 99.5127
R20735 VDD.n3265 VDD.n455 99.5127
R20736 VDD.n3269 VDD.n455 99.5127
R20737 VDD.n3269 VDD.n445 99.5127
R20738 VDD.n3277 VDD.n445 99.5127
R20739 VDD.n3277 VDD.n443 99.5127
R20740 VDD.n3281 VDD.n443 99.5127
R20741 VDD.n3281 VDD.n433 99.5127
R20742 VDD.n3289 VDD.n433 99.5127
R20743 VDD.n3289 VDD.n431 99.5127
R20744 VDD.n3293 VDD.n431 99.5127
R20745 VDD.n3293 VDD.n420 99.5127
R20746 VDD.n3301 VDD.n420 99.5127
R20747 VDD.n3301 VDD.n418 99.5127
R20748 VDD.n3305 VDD.n418 99.5127
R20749 VDD.n3305 VDD.n409 99.5127
R20750 VDD.n3313 VDD.n409 99.5127
R20751 VDD.n3313 VDD.n407 99.5127
R20752 VDD.n3317 VDD.n407 99.5127
R20753 VDD.n3317 VDD.n397 99.5127
R20754 VDD.n3325 VDD.n397 99.5127
R20755 VDD.n3325 VDD.n395 99.5127
R20756 VDD.n3329 VDD.n395 99.5127
R20757 VDD.n3329 VDD.n385 99.5127
R20758 VDD.n3337 VDD.n385 99.5127
R20759 VDD.n3337 VDD.n383 99.5127
R20760 VDD.n3341 VDD.n383 99.5127
R20761 VDD.n3341 VDD.n372 99.5127
R20762 VDD.n3349 VDD.n372 99.5127
R20763 VDD.n3349 VDD.n370 99.5127
R20764 VDD.n3353 VDD.n370 99.5127
R20765 VDD.n3353 VDD.n361 99.5127
R20766 VDD.n3361 VDD.n361 99.5127
R20767 VDD.n3361 VDD.n359 99.5127
R20768 VDD.n3365 VDD.n359 99.5127
R20769 VDD.n3365 VDD.n348 99.5127
R20770 VDD.n3398 VDD.n348 99.5127
R20771 VDD.n3398 VDD.n346 99.5127
R20772 VDD.n3402 VDD.n346 99.5127
R20773 VDD.n3402 VDD.n325 99.5127
R20774 VDD.n3442 VDD.n325 99.5127
R20775 VDD.n3442 VDD.n326 99.5127
R20776 VDD.n3436 VDD.n3435 99.5127
R20777 VDD.n3433 VDD.n330 99.5127
R20778 VDD.n3429 VDD.n3428 99.5127
R20779 VDD.n3426 VDD.n3424 99.5127
R20780 VDD.n3422 VDD.n334 99.5127
R20781 VDD.n3418 VDD.n3417 99.5127
R20782 VDD.n3415 VDD.n340 99.5127
R20783 VDD.n2781 VDD.n2560 99.5127
R20784 VDD.n2560 VDD.n705 99.5127
R20785 VDD.n2776 VDD.n705 99.5127
R20786 VDD.n2776 VDD.n699 99.5127
R20787 VDD.n2773 VDD.n699 99.5127
R20788 VDD.n2773 VDD.n693 99.5127
R20789 VDD.n2770 VDD.n693 99.5127
R20790 VDD.n2770 VDD.n687 99.5127
R20791 VDD.n2767 VDD.n687 99.5127
R20792 VDD.n2767 VDD.n680 99.5127
R20793 VDD.n2764 VDD.n680 99.5127
R20794 VDD.n2764 VDD.n674 99.5127
R20795 VDD.n2761 VDD.n674 99.5127
R20796 VDD.n2761 VDD.n669 99.5127
R20797 VDD.n2758 VDD.n669 99.5127
R20798 VDD.n2758 VDD.n663 99.5127
R20799 VDD.n2755 VDD.n663 99.5127
R20800 VDD.n2755 VDD.n657 99.5127
R20801 VDD.n2752 VDD.n657 99.5127
R20802 VDD.n2752 VDD.n651 99.5127
R20803 VDD.n2749 VDD.n651 99.5127
R20804 VDD.n2749 VDD.n645 99.5127
R20805 VDD.n2746 VDD.n645 99.5127
R20806 VDD.n2746 VDD.n639 99.5127
R20807 VDD.n2743 VDD.n639 99.5127
R20808 VDD.n2743 VDD.n633 99.5127
R20809 VDD.n2740 VDD.n633 99.5127
R20810 VDD.n2740 VDD.n627 99.5127
R20811 VDD.n2737 VDD.n627 99.5127
R20812 VDD.n2737 VDD.n620 99.5127
R20813 VDD.n2734 VDD.n620 99.5127
R20814 VDD.n2734 VDD.n614 99.5127
R20815 VDD.n2731 VDD.n614 99.5127
R20816 VDD.n2731 VDD.n609 99.5127
R20817 VDD.n2728 VDD.n609 99.5127
R20818 VDD.n2728 VDD.n603 99.5127
R20819 VDD.n2725 VDD.n603 99.5127
R20820 VDD.n2725 VDD.n597 99.5127
R20821 VDD.n2722 VDD.n597 99.5127
R20822 VDD.n2722 VDD.n591 99.5127
R20823 VDD.n2719 VDD.n591 99.5127
R20824 VDD.n2719 VDD.n585 99.5127
R20825 VDD.n2716 VDD.n585 99.5127
R20826 VDD.n2716 VDD.n579 99.5127
R20827 VDD.n2713 VDD.n579 99.5127
R20828 VDD.n2713 VDD.n573 99.5127
R20829 VDD.n2710 VDD.n573 99.5127
R20830 VDD.n2710 VDD.n567 99.5127
R20831 VDD.n2707 VDD.n567 99.5127
R20832 VDD.n2707 VDD.n561 99.5127
R20833 VDD.n2704 VDD.n561 99.5127
R20834 VDD.n2704 VDD.n554 99.5127
R20835 VDD.n2701 VDD.n554 99.5127
R20836 VDD.n2701 VDD.n548 99.5127
R20837 VDD.n2698 VDD.n548 99.5127
R20838 VDD.n2698 VDD.n543 99.5127
R20839 VDD.n2695 VDD.n543 99.5127
R20840 VDD.n2695 VDD.n537 99.5127
R20841 VDD.n2692 VDD.n537 99.5127
R20842 VDD.n2692 VDD.n531 99.5127
R20843 VDD.n2689 VDD.n531 99.5127
R20844 VDD.n2689 VDD.n525 99.5127
R20845 VDD.n2686 VDD.n525 99.5127
R20846 VDD.n2686 VDD.n519 99.5127
R20847 VDD.n2683 VDD.n519 99.5127
R20848 VDD.n2683 VDD.n513 99.5127
R20849 VDD.n2680 VDD.n513 99.5127
R20850 VDD.n2680 VDD.n506 99.5127
R20851 VDD.n2677 VDD.n506 99.5127
R20852 VDD.n2677 VDD.n499 99.5127
R20853 VDD.n2674 VDD.n499 99.5127
R20854 VDD.n2674 VDD.n494 99.5127
R20855 VDD.n2671 VDD.n494 99.5127
R20856 VDD.n2671 VDD.n489 99.5127
R20857 VDD.n2668 VDD.n489 99.5127
R20858 VDD.n2668 VDD.n483 99.5127
R20859 VDD.n2665 VDD.n483 99.5127
R20860 VDD.n2665 VDD.n477 99.5127
R20861 VDD.n2662 VDD.n477 99.5127
R20862 VDD.n2662 VDD.n471 99.5127
R20863 VDD.n2659 VDD.n471 99.5127
R20864 VDD.n2659 VDD.n465 99.5127
R20865 VDD.n2656 VDD.n465 99.5127
R20866 VDD.n2656 VDD.n459 99.5127
R20867 VDD.n2653 VDD.n459 99.5127
R20868 VDD.n2653 VDD.n453 99.5127
R20869 VDD.n2650 VDD.n453 99.5127
R20870 VDD.n2650 VDD.n447 99.5127
R20871 VDD.n2647 VDD.n447 99.5127
R20872 VDD.n2647 VDD.n441 99.5127
R20873 VDD.n2644 VDD.n441 99.5127
R20874 VDD.n2644 VDD.n435 99.5127
R20875 VDD.n2641 VDD.n435 99.5127
R20876 VDD.n2641 VDD.n429 99.5127
R20877 VDD.n2638 VDD.n429 99.5127
R20878 VDD.n2638 VDD.n422 99.5127
R20879 VDD.n2635 VDD.n422 99.5127
R20880 VDD.n2635 VDD.n416 99.5127
R20881 VDD.n2632 VDD.n416 99.5127
R20882 VDD.n2632 VDD.n411 99.5127
R20883 VDD.n2629 VDD.n411 99.5127
R20884 VDD.n2629 VDD.n405 99.5127
R20885 VDD.n2626 VDD.n405 99.5127
R20886 VDD.n2626 VDD.n399 99.5127
R20887 VDD.n2623 VDD.n399 99.5127
R20888 VDD.n2623 VDD.n393 99.5127
R20889 VDD.n2620 VDD.n393 99.5127
R20890 VDD.n2620 VDD.n387 99.5127
R20891 VDD.n2617 VDD.n387 99.5127
R20892 VDD.n2617 VDD.n381 99.5127
R20893 VDD.n2614 VDD.n381 99.5127
R20894 VDD.n2614 VDD.n374 99.5127
R20895 VDD.n2611 VDD.n374 99.5127
R20896 VDD.n2611 VDD.n368 99.5127
R20897 VDD.n2608 VDD.n368 99.5127
R20898 VDD.n2608 VDD.n363 99.5127
R20899 VDD.n2605 VDD.n363 99.5127
R20900 VDD.n2605 VDD.n357 99.5127
R20901 VDD.n2602 VDD.n357 99.5127
R20902 VDD.n2602 VDD.n350 99.5127
R20903 VDD.n350 VDD.n342 99.5127
R20904 VDD.n3404 VDD.n342 99.5127
R20905 VDD.n3405 VDD.n3404 99.5127
R20906 VDD.n3405 VDD.n322 99.5127
R20907 VDD.n3410 VDD.n322 99.5127
R20908 VDD.n2569 VDD.n2567 99.5127
R20909 VDD.n2573 VDD.n2567 99.5127
R20910 VDD.n2577 VDD.n2575 99.5127
R20911 VDD.n2581 VDD.n2565 99.5127
R20912 VDD.n2585 VDD.n2583 99.5127
R20913 VDD.n2592 VDD.n2563 99.5127
R20914 VDD.n2595 VDD.n2594 99.5127
R20915 VDD.n2597 VDD.n2559 99.5127
R20916 VDD.n2543 VDD.n2542 99.5127
R20917 VDD.n2539 VDD.n2538 99.5127
R20918 VDD.n2535 VDD.n2534 99.5127
R20919 VDD.n2531 VDD.n2530 99.5127
R20920 VDD.n2527 VDD.n2526 99.5127
R20921 VDD.n2523 VDD.n2522 99.5127
R20922 VDD.n2519 VDD.n2518 99.5127
R20923 VDD.n1715 VDD.n1109 99.5127
R20924 VDD.n1715 VDD.n1103 99.5127
R20925 VDD.n1718 VDD.n1103 99.5127
R20926 VDD.n1718 VDD.n1097 99.5127
R20927 VDD.n1721 VDD.n1097 99.5127
R20928 VDD.n1721 VDD.n1091 99.5127
R20929 VDD.n1724 VDD.n1091 99.5127
R20930 VDD.n1724 VDD.n1085 99.5127
R20931 VDD.n1727 VDD.n1085 99.5127
R20932 VDD.n1727 VDD.n1078 99.5127
R20933 VDD.n1730 VDD.n1078 99.5127
R20934 VDD.n1730 VDD.n1072 99.5127
R20935 VDD.n1733 VDD.n1072 99.5127
R20936 VDD.n1733 VDD.n1067 99.5127
R20937 VDD.n1736 VDD.n1067 99.5127
R20938 VDD.n1736 VDD.n1061 99.5127
R20939 VDD.n1739 VDD.n1061 99.5127
R20940 VDD.n1739 VDD.n1055 99.5127
R20941 VDD.n1742 VDD.n1055 99.5127
R20942 VDD.n1742 VDD.n1049 99.5127
R20943 VDD.n1745 VDD.n1049 99.5127
R20944 VDD.n1745 VDD.n1043 99.5127
R20945 VDD.n1748 VDD.n1043 99.5127
R20946 VDD.n1748 VDD.n1037 99.5127
R20947 VDD.n1751 VDD.n1037 99.5127
R20948 VDD.n1751 VDD.n1030 99.5127
R20949 VDD.n1754 VDD.n1030 99.5127
R20950 VDD.n1754 VDD.n1024 99.5127
R20951 VDD.n1757 VDD.n1024 99.5127
R20952 VDD.n1757 VDD.n1019 99.5127
R20953 VDD.n1760 VDD.n1019 99.5127
R20954 VDD.n1760 VDD.n1013 99.5127
R20955 VDD.n1763 VDD.n1013 99.5127
R20956 VDD.n1763 VDD.n1007 99.5127
R20957 VDD.n1766 VDD.n1007 99.5127
R20958 VDD.n1766 VDD.n1001 99.5127
R20959 VDD.n1769 VDD.n1001 99.5127
R20960 VDD.n1769 VDD.n995 99.5127
R20961 VDD.n1772 VDD.n995 99.5127
R20962 VDD.n1772 VDD.n989 99.5127
R20963 VDD.n1775 VDD.n989 99.5127
R20964 VDD.n1775 VDD.n983 99.5127
R20965 VDD.n1778 VDD.n983 99.5127
R20966 VDD.n1778 VDD.n977 99.5127
R20967 VDD.n1781 VDD.n977 99.5127
R20968 VDD.n1781 VDD.n971 99.5127
R20969 VDD.n1784 VDD.n971 99.5127
R20970 VDD.n1784 VDD.n965 99.5127
R20971 VDD.n1787 VDD.n965 99.5127
R20972 VDD.n1787 VDD.n959 99.5127
R20973 VDD.n1790 VDD.n959 99.5127
R20974 VDD.n1790 VDD.n952 99.5127
R20975 VDD.n1793 VDD.n952 99.5127
R20976 VDD.n1793 VDD.n945 99.5127
R20977 VDD.n1796 VDD.n945 99.5127
R20978 VDD.n1796 VDD.n940 99.5127
R20979 VDD.n1799 VDD.n940 99.5127
R20980 VDD.n1799 VDD.n935 99.5127
R20981 VDD.n1802 VDD.n935 99.5127
R20982 VDD.n1802 VDD.n929 99.5127
R20983 VDD.n1805 VDD.n929 99.5127
R20984 VDD.n1805 VDD.n923 99.5127
R20985 VDD.n1808 VDD.n923 99.5127
R20986 VDD.n1808 VDD.n917 99.5127
R20987 VDD.n1811 VDD.n917 99.5127
R20988 VDD.n1811 VDD.n911 99.5127
R20989 VDD.n1814 VDD.n911 99.5127
R20990 VDD.n1814 VDD.n905 99.5127
R20991 VDD.n1817 VDD.n905 99.5127
R20992 VDD.n1817 VDD.n898 99.5127
R20993 VDD.n1820 VDD.n898 99.5127
R20994 VDD.n1820 VDD.n892 99.5127
R20995 VDD.n1823 VDD.n892 99.5127
R20996 VDD.n1823 VDD.n887 99.5127
R20997 VDD.n1826 VDD.n887 99.5127
R20998 VDD.n1826 VDD.n881 99.5127
R20999 VDD.n1829 VDD.n881 99.5127
R21000 VDD.n1829 VDD.n875 99.5127
R21001 VDD.n1832 VDD.n875 99.5127
R21002 VDD.n1832 VDD.n869 99.5127
R21003 VDD.n1835 VDD.n869 99.5127
R21004 VDD.n1835 VDD.n863 99.5127
R21005 VDD.n1838 VDD.n863 99.5127
R21006 VDD.n1838 VDD.n857 99.5127
R21007 VDD.n1841 VDD.n857 99.5127
R21008 VDD.n1841 VDD.n851 99.5127
R21009 VDD.n1844 VDD.n851 99.5127
R21010 VDD.n1844 VDD.n845 99.5127
R21011 VDD.n1847 VDD.n845 99.5127
R21012 VDD.n1847 VDD.n839 99.5127
R21013 VDD.n1850 VDD.n839 99.5127
R21014 VDD.n1850 VDD.n832 99.5127
R21015 VDD.n1853 VDD.n832 99.5127
R21016 VDD.n1853 VDD.n826 99.5127
R21017 VDD.n1856 VDD.n826 99.5127
R21018 VDD.n1856 VDD.n821 99.5127
R21019 VDD.n1859 VDD.n821 99.5127
R21020 VDD.n1859 VDD.n815 99.5127
R21021 VDD.n1862 VDD.n815 99.5127
R21022 VDD.n1862 VDD.n809 99.5127
R21023 VDD.n1865 VDD.n809 99.5127
R21024 VDD.n1865 VDD.n803 99.5127
R21025 VDD.n1868 VDD.n803 99.5127
R21026 VDD.n1868 VDD.n797 99.5127
R21027 VDD.n1871 VDD.n797 99.5127
R21028 VDD.n1871 VDD.n791 99.5127
R21029 VDD.n1874 VDD.n791 99.5127
R21030 VDD.n1874 VDD.n785 99.5127
R21031 VDD.n1877 VDD.n785 99.5127
R21032 VDD.n1877 VDD.n779 99.5127
R21033 VDD.n1880 VDD.n779 99.5127
R21034 VDD.n1880 VDD.n773 99.5127
R21035 VDD.n1895 VDD.n773 99.5127
R21036 VDD.n1895 VDD.n767 99.5127
R21037 VDD.n1891 VDD.n767 99.5127
R21038 VDD.n1891 VDD.n762 99.5127
R21039 VDD.n1888 VDD.n762 99.5127
R21040 VDD.n1888 VDD.n756 99.5127
R21041 VDD.n1885 VDD.n756 99.5127
R21042 VDD.n1885 VDD.n749 99.5127
R21043 VDD.n749 VDD.n741 99.5127
R21044 VDD.n2509 VDD.n741 99.5127
R21045 VDD.n2510 VDD.n2509 99.5127
R21046 VDD.n2510 VDD.n732 99.5127
R21047 VDD.n2514 VDD.n732 99.5127
R21048 VDD.n1147 VDD.n1146 99.5127
R21049 VDD.n1149 VDD.n1147 99.5127
R21050 VDD.n1153 VDD.n1142 99.5127
R21051 VDD.n1157 VDD.n1155 99.5127
R21052 VDD.n1700 VDD.n1140 99.5127
R21053 VDD.n1704 VDD.n1702 99.5127
R21054 VDD.n1709 VDD.n1136 99.5127
R21055 VDD.n1712 VDD.n1711 99.5127
R21056 VDD.n2105 VDD.n1105 99.5127
R21057 VDD.n2109 VDD.n1105 99.5127
R21058 VDD.n2109 VDD.n1095 99.5127
R21059 VDD.n2117 VDD.n1095 99.5127
R21060 VDD.n2117 VDD.n1093 99.5127
R21061 VDD.n2121 VDD.n1093 99.5127
R21062 VDD.n2121 VDD.n1083 99.5127
R21063 VDD.n2129 VDD.n1083 99.5127
R21064 VDD.n2129 VDD.n1081 99.5127
R21065 VDD.n2133 VDD.n1081 99.5127
R21066 VDD.n2133 VDD.n1071 99.5127
R21067 VDD.n2141 VDD.n1071 99.5127
R21068 VDD.n2141 VDD.n1069 99.5127
R21069 VDD.n2145 VDD.n1069 99.5127
R21070 VDD.n2145 VDD.n1059 99.5127
R21071 VDD.n2153 VDD.n1059 99.5127
R21072 VDD.n2153 VDD.n1057 99.5127
R21073 VDD.n2157 VDD.n1057 99.5127
R21074 VDD.n2157 VDD.n1047 99.5127
R21075 VDD.n2165 VDD.n1047 99.5127
R21076 VDD.n2165 VDD.n1045 99.5127
R21077 VDD.n2169 VDD.n1045 99.5127
R21078 VDD.n2169 VDD.n1035 99.5127
R21079 VDD.n2177 VDD.n1035 99.5127
R21080 VDD.n2177 VDD.n1033 99.5127
R21081 VDD.n2181 VDD.n1033 99.5127
R21082 VDD.n2181 VDD.n1023 99.5127
R21083 VDD.n2189 VDD.n1023 99.5127
R21084 VDD.n2189 VDD.n1021 99.5127
R21085 VDD.n2193 VDD.n1021 99.5127
R21086 VDD.n2193 VDD.n1011 99.5127
R21087 VDD.n2201 VDD.n1011 99.5127
R21088 VDD.n2201 VDD.n1009 99.5127
R21089 VDD.n2205 VDD.n1009 99.5127
R21090 VDD.n2205 VDD.n999 99.5127
R21091 VDD.n2213 VDD.n999 99.5127
R21092 VDD.n2213 VDD.n997 99.5127
R21093 VDD.n2217 VDD.n997 99.5127
R21094 VDD.n2217 VDD.n987 99.5127
R21095 VDD.n2225 VDD.n987 99.5127
R21096 VDD.n2225 VDD.n985 99.5127
R21097 VDD.n2229 VDD.n985 99.5127
R21098 VDD.n2229 VDD.n975 99.5127
R21099 VDD.n2237 VDD.n975 99.5127
R21100 VDD.n2237 VDD.n973 99.5127
R21101 VDD.n2241 VDD.n973 99.5127
R21102 VDD.n2241 VDD.n963 99.5127
R21103 VDD.n2249 VDD.n963 99.5127
R21104 VDD.n2249 VDD.n961 99.5127
R21105 VDD.n2253 VDD.n961 99.5127
R21106 VDD.n2253 VDD.n950 99.5127
R21107 VDD.n2261 VDD.n950 99.5127
R21108 VDD.n2261 VDD.n948 99.5127
R21109 VDD.n2265 VDD.n948 99.5127
R21110 VDD.n2265 VDD.n939 99.5127
R21111 VDD.n2273 VDD.n939 99.5127
R21112 VDD.n2273 VDD.n937 99.5127
R21113 VDD.n2277 VDD.n937 99.5127
R21114 VDD.n2277 VDD.n927 99.5127
R21115 VDD.n2285 VDD.n927 99.5127
R21116 VDD.n2285 VDD.n925 99.5127
R21117 VDD.n2289 VDD.n925 99.5127
R21118 VDD.n2289 VDD.n915 99.5127
R21119 VDD.n2297 VDD.n915 99.5127
R21120 VDD.n2297 VDD.n913 99.5127
R21121 VDD.n2301 VDD.n913 99.5127
R21122 VDD.n2301 VDD.n903 99.5127
R21123 VDD.n2309 VDD.n903 99.5127
R21124 VDD.n2309 VDD.n901 99.5127
R21125 VDD.n2313 VDD.n901 99.5127
R21126 VDD.n2313 VDD.n891 99.5127
R21127 VDD.n2321 VDD.n891 99.5127
R21128 VDD.n2321 VDD.n889 99.5127
R21129 VDD.n2325 VDD.n889 99.5127
R21130 VDD.n2325 VDD.n879 99.5127
R21131 VDD.n2333 VDD.n879 99.5127
R21132 VDD.n2333 VDD.n877 99.5127
R21133 VDD.n2337 VDD.n877 99.5127
R21134 VDD.n2337 VDD.n867 99.5127
R21135 VDD.n2345 VDD.n867 99.5127
R21136 VDD.n2345 VDD.n865 99.5127
R21137 VDD.n2349 VDD.n865 99.5127
R21138 VDD.n2349 VDD.n855 99.5127
R21139 VDD.n2357 VDD.n855 99.5127
R21140 VDD.n2357 VDD.n853 99.5127
R21141 VDD.n2361 VDD.n853 99.5127
R21142 VDD.n2361 VDD.n843 99.5127
R21143 VDD.n2369 VDD.n843 99.5127
R21144 VDD.n2369 VDD.n841 99.5127
R21145 VDD.n2373 VDD.n841 99.5127
R21146 VDD.n2373 VDD.n830 99.5127
R21147 VDD.n2381 VDD.n830 99.5127
R21148 VDD.n2381 VDD.n828 99.5127
R21149 VDD.n2385 VDD.n828 99.5127
R21150 VDD.n2385 VDD.n819 99.5127
R21151 VDD.n2393 VDD.n819 99.5127
R21152 VDD.n2393 VDD.n817 99.5127
R21153 VDD.n2397 VDD.n817 99.5127
R21154 VDD.n2397 VDD.n807 99.5127
R21155 VDD.n2405 VDD.n807 99.5127
R21156 VDD.n2405 VDD.n805 99.5127
R21157 VDD.n2409 VDD.n805 99.5127
R21158 VDD.n2409 VDD.n795 99.5127
R21159 VDD.n2417 VDD.n795 99.5127
R21160 VDD.n2417 VDD.n793 99.5127
R21161 VDD.n2421 VDD.n793 99.5127
R21162 VDD.n2421 VDD.n783 99.5127
R21163 VDD.n2429 VDD.n783 99.5127
R21164 VDD.n2429 VDD.n781 99.5127
R21165 VDD.n2433 VDD.n781 99.5127
R21166 VDD.n2433 VDD.n771 99.5127
R21167 VDD.n2441 VDD.n771 99.5127
R21168 VDD.n2441 VDD.n769 99.5127
R21169 VDD.n2445 VDD.n769 99.5127
R21170 VDD.n2445 VDD.n760 99.5127
R21171 VDD.n2453 VDD.n760 99.5127
R21172 VDD.n2453 VDD.n758 99.5127
R21173 VDD.n2457 VDD.n758 99.5127
R21174 VDD.n2457 VDD.n747 99.5127
R21175 VDD.n2503 VDD.n747 99.5127
R21176 VDD.n2503 VDD.n745 99.5127
R21177 VDD.n2507 VDD.n745 99.5127
R21178 VDD.n2507 VDD.n734 99.5127
R21179 VDD.n2549 VDD.n734 99.5127
R21180 VDD.n2549 VDD.n735 99.5127
R21181 VDD.n3385 VDD.n3371 99.5127
R21182 VDD.n3381 VDD.n3380 99.5127
R21183 VDD.n3378 VDD.n3375 99.5127
R21184 VDD.n3461 VDD.n310 99.5127
R21185 VDD.n3459 VDD.n3458 99.5127
R21186 VDD.n3456 VDD.n313 99.5127
R21187 VDD.n3451 VDD.n3450 99.5127
R21188 VDD.n2974 VDD.n2782 99.5127
R21189 VDD.n2974 VDD.n706 99.5127
R21190 VDD.n2971 VDD.n706 99.5127
R21191 VDD.n2971 VDD.n700 99.5127
R21192 VDD.n2968 VDD.n700 99.5127
R21193 VDD.n2968 VDD.n694 99.5127
R21194 VDD.n2965 VDD.n694 99.5127
R21195 VDD.n2965 VDD.n688 99.5127
R21196 VDD.n2962 VDD.n688 99.5127
R21197 VDD.n2962 VDD.n681 99.5127
R21198 VDD.n2959 VDD.n681 99.5127
R21199 VDD.n2959 VDD.n675 99.5127
R21200 VDD.n2956 VDD.n675 99.5127
R21201 VDD.n2956 VDD.n670 99.5127
R21202 VDD.n2953 VDD.n670 99.5127
R21203 VDD.n2953 VDD.n664 99.5127
R21204 VDD.n2950 VDD.n664 99.5127
R21205 VDD.n2950 VDD.n658 99.5127
R21206 VDD.n2947 VDD.n658 99.5127
R21207 VDD.n2947 VDD.n652 99.5127
R21208 VDD.n2944 VDD.n652 99.5127
R21209 VDD.n2944 VDD.n646 99.5127
R21210 VDD.n2941 VDD.n646 99.5127
R21211 VDD.n2941 VDD.n640 99.5127
R21212 VDD.n2938 VDD.n640 99.5127
R21213 VDD.n2938 VDD.n634 99.5127
R21214 VDD.n2935 VDD.n634 99.5127
R21215 VDD.n2935 VDD.n628 99.5127
R21216 VDD.n2932 VDD.n628 99.5127
R21217 VDD.n2932 VDD.n621 99.5127
R21218 VDD.n2929 VDD.n621 99.5127
R21219 VDD.n2929 VDD.n615 99.5127
R21220 VDD.n2926 VDD.n615 99.5127
R21221 VDD.n2926 VDD.n610 99.5127
R21222 VDD.n2923 VDD.n610 99.5127
R21223 VDD.n2923 VDD.n604 99.5127
R21224 VDD.n2920 VDD.n604 99.5127
R21225 VDD.n2920 VDD.n598 99.5127
R21226 VDD.n2917 VDD.n598 99.5127
R21227 VDD.n2917 VDD.n592 99.5127
R21228 VDD.n2914 VDD.n592 99.5127
R21229 VDD.n2914 VDD.n586 99.5127
R21230 VDD.n2911 VDD.n586 99.5127
R21231 VDD.n2911 VDD.n580 99.5127
R21232 VDD.n2908 VDD.n580 99.5127
R21233 VDD.n2908 VDD.n574 99.5127
R21234 VDD.n2905 VDD.n574 99.5127
R21235 VDD.n2905 VDD.n568 99.5127
R21236 VDD.n2902 VDD.n568 99.5127
R21237 VDD.n2902 VDD.n562 99.5127
R21238 VDD.n2899 VDD.n562 99.5127
R21239 VDD.n2899 VDD.n555 99.5127
R21240 VDD.n2896 VDD.n555 99.5127
R21241 VDD.n2896 VDD.n549 99.5127
R21242 VDD.n2893 VDD.n549 99.5127
R21243 VDD.n2893 VDD.n544 99.5127
R21244 VDD.n2890 VDD.n544 99.5127
R21245 VDD.n2890 VDD.n538 99.5127
R21246 VDD.n2887 VDD.n538 99.5127
R21247 VDD.n2887 VDD.n532 99.5127
R21248 VDD.n2884 VDD.n532 99.5127
R21249 VDD.n2884 VDD.n526 99.5127
R21250 VDD.n2881 VDD.n526 99.5127
R21251 VDD.n2881 VDD.n520 99.5127
R21252 VDD.n2878 VDD.n520 99.5127
R21253 VDD.n2878 VDD.n514 99.5127
R21254 VDD.n2875 VDD.n514 99.5127
R21255 VDD.n2875 VDD.n507 99.5127
R21256 VDD.n2872 VDD.n507 99.5127
R21257 VDD.n2872 VDD.n500 99.5127
R21258 VDD.n2869 VDD.n500 99.5127
R21259 VDD.n2869 VDD.n495 99.5127
R21260 VDD.n2866 VDD.n495 99.5127
R21261 VDD.n2866 VDD.n490 99.5127
R21262 VDD.n2863 VDD.n490 99.5127
R21263 VDD.n2863 VDD.n484 99.5127
R21264 VDD.n2860 VDD.n484 99.5127
R21265 VDD.n2860 VDD.n478 99.5127
R21266 VDD.n2857 VDD.n478 99.5127
R21267 VDD.n2857 VDD.n472 99.5127
R21268 VDD.n2854 VDD.n472 99.5127
R21269 VDD.n2854 VDD.n466 99.5127
R21270 VDD.n2851 VDD.n466 99.5127
R21271 VDD.n2851 VDD.n460 99.5127
R21272 VDD.n2848 VDD.n460 99.5127
R21273 VDD.n2848 VDD.n454 99.5127
R21274 VDD.n2845 VDD.n454 99.5127
R21275 VDD.n2845 VDD.n448 99.5127
R21276 VDD.n2842 VDD.n448 99.5127
R21277 VDD.n2842 VDD.n442 99.5127
R21278 VDD.n2839 VDD.n442 99.5127
R21279 VDD.n2839 VDD.n436 99.5127
R21280 VDD.n2836 VDD.n436 99.5127
R21281 VDD.n2836 VDD.n430 99.5127
R21282 VDD.n2833 VDD.n430 99.5127
R21283 VDD.n2833 VDD.n423 99.5127
R21284 VDD.n2830 VDD.n423 99.5127
R21285 VDD.n2830 VDD.n417 99.5127
R21286 VDD.n2827 VDD.n417 99.5127
R21287 VDD.n2827 VDD.n412 99.5127
R21288 VDD.n2824 VDD.n412 99.5127
R21289 VDD.n2824 VDD.n406 99.5127
R21290 VDD.n2821 VDD.n406 99.5127
R21291 VDD.n2821 VDD.n400 99.5127
R21292 VDD.n2818 VDD.n400 99.5127
R21293 VDD.n2818 VDD.n394 99.5127
R21294 VDD.n2815 VDD.n394 99.5127
R21295 VDD.n2815 VDD.n388 99.5127
R21296 VDD.n2812 VDD.n388 99.5127
R21297 VDD.n2812 VDD.n382 99.5127
R21298 VDD.n2809 VDD.n382 99.5127
R21299 VDD.n2809 VDD.n375 99.5127
R21300 VDD.n2806 VDD.n375 99.5127
R21301 VDD.n2806 VDD.n369 99.5127
R21302 VDD.n2803 VDD.n369 99.5127
R21303 VDD.n2803 VDD.n364 99.5127
R21304 VDD.n2800 VDD.n364 99.5127
R21305 VDD.n2800 VDD.n358 99.5127
R21306 VDD.n2797 VDD.n358 99.5127
R21307 VDD.n2797 VDD.n351 99.5127
R21308 VDD.n2794 VDD.n351 99.5127
R21309 VDD.n2794 VDD.n344 99.5127
R21310 VDD.n344 VDD.n320 99.5127
R21311 VDD.n3444 VDD.n320 99.5127
R21312 VDD.n3444 VDD.n318 99.5127
R21313 VDD.n3007 VDD.n3005 99.5127
R21314 VDD.n3003 VDD.n2785 99.5127
R21315 VDD.n2999 VDD.n2997 99.5127
R21316 VDD.n2995 VDD.n2787 99.5127
R21317 VDD.n2991 VDD.n2989 99.5127
R21318 VDD.n2987 VDD.n2789 99.5127
R21319 VDD.n2982 VDD.n2980 99.5127
R21320 VDD.n3011 VDD.n703 99.5127
R21321 VDD.n3019 VDD.n703 99.5127
R21322 VDD.n3019 VDD.n701 99.5127
R21323 VDD.n3023 VDD.n701 99.5127
R21324 VDD.n3023 VDD.n691 99.5127
R21325 VDD.n3031 VDD.n691 99.5127
R21326 VDD.n3031 VDD.n689 99.5127
R21327 VDD.n3035 VDD.n689 99.5127
R21328 VDD.n3035 VDD.n678 99.5127
R21329 VDD.n3043 VDD.n678 99.5127
R21330 VDD.n3043 VDD.n676 99.5127
R21331 VDD.n3047 VDD.n676 99.5127
R21332 VDD.n3047 VDD.n667 99.5127
R21333 VDD.n3055 VDD.n667 99.5127
R21334 VDD.n3055 VDD.n665 99.5127
R21335 VDD.n3059 VDD.n665 99.5127
R21336 VDD.n3059 VDD.n655 99.5127
R21337 VDD.n3067 VDD.n655 99.5127
R21338 VDD.n3067 VDD.n653 99.5127
R21339 VDD.n3071 VDD.n653 99.5127
R21340 VDD.n3071 VDD.n643 99.5127
R21341 VDD.n3079 VDD.n643 99.5127
R21342 VDD.n3079 VDD.n641 99.5127
R21343 VDD.n3083 VDD.n641 99.5127
R21344 VDD.n3083 VDD.n631 99.5127
R21345 VDD.n3091 VDD.n631 99.5127
R21346 VDD.n3091 VDD.n629 99.5127
R21347 VDD.n3095 VDD.n629 99.5127
R21348 VDD.n3095 VDD.n618 99.5127
R21349 VDD.n3103 VDD.n618 99.5127
R21350 VDD.n3103 VDD.n616 99.5127
R21351 VDD.n3107 VDD.n616 99.5127
R21352 VDD.n3107 VDD.n607 99.5127
R21353 VDD.n3115 VDD.n607 99.5127
R21354 VDD.n3115 VDD.n605 99.5127
R21355 VDD.n3119 VDD.n605 99.5127
R21356 VDD.n3119 VDD.n595 99.5127
R21357 VDD.n3127 VDD.n595 99.5127
R21358 VDD.n3127 VDD.n593 99.5127
R21359 VDD.n3131 VDD.n593 99.5127
R21360 VDD.n3131 VDD.n583 99.5127
R21361 VDD.n3139 VDD.n583 99.5127
R21362 VDD.n3139 VDD.n581 99.5127
R21363 VDD.n3143 VDD.n581 99.5127
R21364 VDD.n3143 VDD.n571 99.5127
R21365 VDD.n3151 VDD.n571 99.5127
R21366 VDD.n3151 VDD.n569 99.5127
R21367 VDD.n3155 VDD.n569 99.5127
R21368 VDD.n3155 VDD.n559 99.5127
R21369 VDD.n3163 VDD.n559 99.5127
R21370 VDD.n3163 VDD.n557 99.5127
R21371 VDD.n3167 VDD.n557 99.5127
R21372 VDD.n3167 VDD.n547 99.5127
R21373 VDD.n3175 VDD.n547 99.5127
R21374 VDD.n3175 VDD.n545 99.5127
R21375 VDD.n3179 VDD.n545 99.5127
R21376 VDD.n3179 VDD.n535 99.5127
R21377 VDD.n3187 VDD.n535 99.5127
R21378 VDD.n3187 VDD.n533 99.5127
R21379 VDD.n3191 VDD.n533 99.5127
R21380 VDD.n3191 VDD.n523 99.5127
R21381 VDD.n3199 VDD.n523 99.5127
R21382 VDD.n3199 VDD.n521 99.5127
R21383 VDD.n3203 VDD.n521 99.5127
R21384 VDD.n3203 VDD.n511 99.5127
R21385 VDD.n3211 VDD.n511 99.5127
R21386 VDD.n3211 VDD.n509 99.5127
R21387 VDD.n3215 VDD.n509 99.5127
R21388 VDD.n3215 VDD.n498 99.5127
R21389 VDD.n3223 VDD.n498 99.5127
R21390 VDD.n3223 VDD.n496 99.5127
R21391 VDD.n3227 VDD.n496 99.5127
R21392 VDD.n3227 VDD.n487 99.5127
R21393 VDD.n3235 VDD.n487 99.5127
R21394 VDD.n3235 VDD.n485 99.5127
R21395 VDD.n3239 VDD.n485 99.5127
R21396 VDD.n3239 VDD.n475 99.5127
R21397 VDD.n3247 VDD.n475 99.5127
R21398 VDD.n3247 VDD.n473 99.5127
R21399 VDD.n3251 VDD.n473 99.5127
R21400 VDD.n3251 VDD.n463 99.5127
R21401 VDD.n3259 VDD.n463 99.5127
R21402 VDD.n3259 VDD.n461 99.5127
R21403 VDD.n3263 VDD.n461 99.5127
R21404 VDD.n3263 VDD.n451 99.5127
R21405 VDD.n3271 VDD.n451 99.5127
R21406 VDD.n3271 VDD.n449 99.5127
R21407 VDD.n3275 VDD.n449 99.5127
R21408 VDD.n3275 VDD.n439 99.5127
R21409 VDD.n3283 VDD.n439 99.5127
R21410 VDD.n3283 VDD.n437 99.5127
R21411 VDD.n3287 VDD.n437 99.5127
R21412 VDD.n3287 VDD.n427 99.5127
R21413 VDD.n3295 VDD.n427 99.5127
R21414 VDD.n3295 VDD.n425 99.5127
R21415 VDD.n3299 VDD.n425 99.5127
R21416 VDD.n3299 VDD.n415 99.5127
R21417 VDD.n3307 VDD.n415 99.5127
R21418 VDD.n3307 VDD.n413 99.5127
R21419 VDD.n3311 VDD.n413 99.5127
R21420 VDD.n3311 VDD.n403 99.5127
R21421 VDD.n3319 VDD.n403 99.5127
R21422 VDD.n3319 VDD.n401 99.5127
R21423 VDD.n3323 VDD.n401 99.5127
R21424 VDD.n3323 VDD.n391 99.5127
R21425 VDD.n3331 VDD.n391 99.5127
R21426 VDD.n3331 VDD.n389 99.5127
R21427 VDD.n3335 VDD.n389 99.5127
R21428 VDD.n3335 VDD.n379 99.5127
R21429 VDD.n3343 VDD.n379 99.5127
R21430 VDD.n3343 VDD.n377 99.5127
R21431 VDD.n3347 VDD.n377 99.5127
R21432 VDD.n3347 VDD.n367 99.5127
R21433 VDD.n3355 VDD.n367 99.5127
R21434 VDD.n3355 VDD.n365 99.5127
R21435 VDD.n3359 VDD.n365 99.5127
R21436 VDD.n3359 VDD.n355 99.5127
R21437 VDD.n3367 VDD.n355 99.5127
R21438 VDD.n3367 VDD.n352 99.5127
R21439 VDD.n3396 VDD.n352 99.5127
R21440 VDD.n3396 VDD.n353 99.5127
R21441 VDD.n353 VDD.n345 99.5127
R21442 VDD.n3391 VDD.n345 99.5127
R21443 VDD.n3391 VDD.n324 99.5127
R21444 VDD.n3388 VDD.n324 99.5127
R21445 VDD.n2489 VDD.n2488 99.5127
R21446 VDD.n2485 VDD.n2484 99.5127
R21447 VDD.n2481 VDD.n2480 99.5127
R21448 VDD.n2477 VDD.n2476 99.5127
R21449 VDD.n2473 VDD.n2472 99.5127
R21450 VDD.n2469 VDD.n2468 99.5127
R21451 VDD.n2465 VDD.n726 99.5127
R21452 VDD.n2065 VDD.n1110 99.5127
R21453 VDD.n2065 VDD.n1104 99.5127
R21454 VDD.n2062 VDD.n1104 99.5127
R21455 VDD.n2062 VDD.n1098 99.5127
R21456 VDD.n2059 VDD.n1098 99.5127
R21457 VDD.n2059 VDD.n1092 99.5127
R21458 VDD.n2056 VDD.n1092 99.5127
R21459 VDD.n2056 VDD.n1086 99.5127
R21460 VDD.n2053 VDD.n1086 99.5127
R21461 VDD.n2053 VDD.n1079 99.5127
R21462 VDD.n2050 VDD.n1079 99.5127
R21463 VDD.n2050 VDD.n1073 99.5127
R21464 VDD.n2047 VDD.n1073 99.5127
R21465 VDD.n2047 VDD.n1068 99.5127
R21466 VDD.n2044 VDD.n1068 99.5127
R21467 VDD.n2044 VDD.n1062 99.5127
R21468 VDD.n2041 VDD.n1062 99.5127
R21469 VDD.n2041 VDD.n1056 99.5127
R21470 VDD.n2038 VDD.n1056 99.5127
R21471 VDD.n2038 VDD.n1050 99.5127
R21472 VDD.n2035 VDD.n1050 99.5127
R21473 VDD.n2035 VDD.n1044 99.5127
R21474 VDD.n2032 VDD.n1044 99.5127
R21475 VDD.n2032 VDD.n1038 99.5127
R21476 VDD.n2029 VDD.n1038 99.5127
R21477 VDD.n2029 VDD.n1031 99.5127
R21478 VDD.n2026 VDD.n1031 99.5127
R21479 VDD.n2026 VDD.n1025 99.5127
R21480 VDD.n2023 VDD.n1025 99.5127
R21481 VDD.n2023 VDD.n1020 99.5127
R21482 VDD.n2020 VDD.n1020 99.5127
R21483 VDD.n2020 VDD.n1014 99.5127
R21484 VDD.n2017 VDD.n1014 99.5127
R21485 VDD.n2017 VDD.n1008 99.5127
R21486 VDD.n2014 VDD.n1008 99.5127
R21487 VDD.n2014 VDD.n1002 99.5127
R21488 VDD.n2011 VDD.n1002 99.5127
R21489 VDD.n2011 VDD.n996 99.5127
R21490 VDD.n2008 VDD.n996 99.5127
R21491 VDD.n2008 VDD.n990 99.5127
R21492 VDD.n2005 VDD.n990 99.5127
R21493 VDD.n2005 VDD.n984 99.5127
R21494 VDD.n2002 VDD.n984 99.5127
R21495 VDD.n2002 VDD.n978 99.5127
R21496 VDD.n1999 VDD.n978 99.5127
R21497 VDD.n1999 VDD.n972 99.5127
R21498 VDD.n1996 VDD.n972 99.5127
R21499 VDD.n1996 VDD.n966 99.5127
R21500 VDD.n1993 VDD.n966 99.5127
R21501 VDD.n1993 VDD.n960 99.5127
R21502 VDD.n1990 VDD.n960 99.5127
R21503 VDD.n1990 VDD.n953 99.5127
R21504 VDD.n1987 VDD.n953 99.5127
R21505 VDD.n1987 VDD.n946 99.5127
R21506 VDD.n1984 VDD.n946 99.5127
R21507 VDD.n1984 VDD.n941 99.5127
R21508 VDD.n1981 VDD.n941 99.5127
R21509 VDD.n1981 VDD.n936 99.5127
R21510 VDD.n1978 VDD.n936 99.5127
R21511 VDD.n1978 VDD.n930 99.5127
R21512 VDD.n1975 VDD.n930 99.5127
R21513 VDD.n1975 VDD.n924 99.5127
R21514 VDD.n1972 VDD.n924 99.5127
R21515 VDD.n1972 VDD.n918 99.5127
R21516 VDD.n1969 VDD.n918 99.5127
R21517 VDD.n1969 VDD.n912 99.5127
R21518 VDD.n1966 VDD.n912 99.5127
R21519 VDD.n1966 VDD.n906 99.5127
R21520 VDD.n1963 VDD.n906 99.5127
R21521 VDD.n1963 VDD.n899 99.5127
R21522 VDD.n1960 VDD.n899 99.5127
R21523 VDD.n1960 VDD.n893 99.5127
R21524 VDD.n1957 VDD.n893 99.5127
R21525 VDD.n1957 VDD.n888 99.5127
R21526 VDD.n1954 VDD.n888 99.5127
R21527 VDD.n1954 VDD.n882 99.5127
R21528 VDD.n1951 VDD.n882 99.5127
R21529 VDD.n1951 VDD.n876 99.5127
R21530 VDD.n1948 VDD.n876 99.5127
R21531 VDD.n1948 VDD.n870 99.5127
R21532 VDD.n1945 VDD.n870 99.5127
R21533 VDD.n1945 VDD.n864 99.5127
R21534 VDD.n1942 VDD.n864 99.5127
R21535 VDD.n1942 VDD.n858 99.5127
R21536 VDD.n1939 VDD.n858 99.5127
R21537 VDD.n1939 VDD.n852 99.5127
R21538 VDD.n1936 VDD.n852 99.5127
R21539 VDD.n1936 VDD.n846 99.5127
R21540 VDD.n1933 VDD.n846 99.5127
R21541 VDD.n1933 VDD.n840 99.5127
R21542 VDD.n1930 VDD.n840 99.5127
R21543 VDD.n1930 VDD.n833 99.5127
R21544 VDD.n1927 VDD.n833 99.5127
R21545 VDD.n1927 VDD.n827 99.5127
R21546 VDD.n1924 VDD.n827 99.5127
R21547 VDD.n1924 VDD.n822 99.5127
R21548 VDD.n1921 VDD.n822 99.5127
R21549 VDD.n1921 VDD.n816 99.5127
R21550 VDD.n1918 VDD.n816 99.5127
R21551 VDD.n1918 VDD.n810 99.5127
R21552 VDD.n1915 VDD.n810 99.5127
R21553 VDD.n1915 VDD.n804 99.5127
R21554 VDD.n1912 VDD.n804 99.5127
R21555 VDD.n1912 VDD.n798 99.5127
R21556 VDD.n1909 VDD.n798 99.5127
R21557 VDD.n1909 VDD.n792 99.5127
R21558 VDD.n1906 VDD.n792 99.5127
R21559 VDD.n1906 VDD.n786 99.5127
R21560 VDD.n1903 VDD.n786 99.5127
R21561 VDD.n1903 VDD.n780 99.5127
R21562 VDD.n1900 VDD.n780 99.5127
R21563 VDD.n1900 VDD.n774 99.5127
R21564 VDD.n1897 VDD.n774 99.5127
R21565 VDD.n1897 VDD.n768 99.5127
R21566 VDD.n1132 VDD.n768 99.5127
R21567 VDD.n1132 VDD.n763 99.5127
R21568 VDD.n1129 VDD.n763 99.5127
R21569 VDD.n1129 VDD.n757 99.5127
R21570 VDD.n1126 VDD.n757 99.5127
R21571 VDD.n1126 VDD.n750 99.5127
R21572 VDD.n1123 VDD.n750 99.5127
R21573 VDD.n1123 VDD.n743 99.5127
R21574 VDD.n743 VDD.n730 99.5127
R21575 VDD.n2551 VDD.n730 99.5127
R21576 VDD.n2551 VDD.n727 99.5127
R21577 VDD.n2099 VDD.n2097 99.5127
R21578 VDD.n2095 VDD.n1113 99.5127
R21579 VDD.n2091 VDD.n2089 99.5127
R21580 VDD.n2087 VDD.n1115 99.5127
R21581 VDD.n2082 VDD.n2080 99.5127
R21582 VDD.n2078 VDD.n1118 99.5127
R21583 VDD.n2073 VDD.n2071 99.5127
R21584 VDD.n2103 VDD.n1101 99.5127
R21585 VDD.n2111 VDD.n1101 99.5127
R21586 VDD.n2111 VDD.n1099 99.5127
R21587 VDD.n2115 VDD.n1099 99.5127
R21588 VDD.n2115 VDD.n1089 99.5127
R21589 VDD.n2123 VDD.n1089 99.5127
R21590 VDD.n2123 VDD.n1087 99.5127
R21591 VDD.n2127 VDD.n1087 99.5127
R21592 VDD.n2127 VDD.n1076 99.5127
R21593 VDD.n2135 VDD.n1076 99.5127
R21594 VDD.n2135 VDD.n1074 99.5127
R21595 VDD.n2139 VDD.n1074 99.5127
R21596 VDD.n2139 VDD.n1065 99.5127
R21597 VDD.n2147 VDD.n1065 99.5127
R21598 VDD.n2147 VDD.n1063 99.5127
R21599 VDD.n2151 VDD.n1063 99.5127
R21600 VDD.n2151 VDD.n1053 99.5127
R21601 VDD.n2159 VDD.n1053 99.5127
R21602 VDD.n2159 VDD.n1051 99.5127
R21603 VDD.n2163 VDD.n1051 99.5127
R21604 VDD.n2163 VDD.n1041 99.5127
R21605 VDD.n2171 VDD.n1041 99.5127
R21606 VDD.n2171 VDD.n1039 99.5127
R21607 VDD.n2175 VDD.n1039 99.5127
R21608 VDD.n2175 VDD.n1028 99.5127
R21609 VDD.n2183 VDD.n1028 99.5127
R21610 VDD.n2183 VDD.n1026 99.5127
R21611 VDD.n2187 VDD.n1026 99.5127
R21612 VDD.n2187 VDD.n1017 99.5127
R21613 VDD.n2195 VDD.n1017 99.5127
R21614 VDD.n2195 VDD.n1015 99.5127
R21615 VDD.n2199 VDD.n1015 99.5127
R21616 VDD.n2199 VDD.n1005 99.5127
R21617 VDD.n2207 VDD.n1005 99.5127
R21618 VDD.n2207 VDD.n1003 99.5127
R21619 VDD.n2211 VDD.n1003 99.5127
R21620 VDD.n2211 VDD.n993 99.5127
R21621 VDD.n2219 VDD.n993 99.5127
R21622 VDD.n2219 VDD.n991 99.5127
R21623 VDD.n2223 VDD.n991 99.5127
R21624 VDD.n2223 VDD.n981 99.5127
R21625 VDD.n2231 VDD.n981 99.5127
R21626 VDD.n2231 VDD.n979 99.5127
R21627 VDD.n2235 VDD.n979 99.5127
R21628 VDD.n2235 VDD.n969 99.5127
R21629 VDD.n2243 VDD.n969 99.5127
R21630 VDD.n2243 VDD.n967 99.5127
R21631 VDD.n2247 VDD.n967 99.5127
R21632 VDD.n2247 VDD.n957 99.5127
R21633 VDD.n2255 VDD.n957 99.5127
R21634 VDD.n2255 VDD.n955 99.5127
R21635 VDD.n2259 VDD.n955 99.5127
R21636 VDD.n2259 VDD.n944 99.5127
R21637 VDD.n2267 VDD.n944 99.5127
R21638 VDD.n2267 VDD.n942 99.5127
R21639 VDD.n2271 VDD.n942 99.5127
R21640 VDD.n2271 VDD.n933 99.5127
R21641 VDD.n2279 VDD.n933 99.5127
R21642 VDD.n2279 VDD.n931 99.5127
R21643 VDD.n2283 VDD.n931 99.5127
R21644 VDD.n2283 VDD.n921 99.5127
R21645 VDD.n2291 VDD.n921 99.5127
R21646 VDD.n2291 VDD.n919 99.5127
R21647 VDD.n2295 VDD.n919 99.5127
R21648 VDD.n2295 VDD.n909 99.5127
R21649 VDD.n2303 VDD.n909 99.5127
R21650 VDD.n2303 VDD.n907 99.5127
R21651 VDD.n2307 VDD.n907 99.5127
R21652 VDD.n2307 VDD.n896 99.5127
R21653 VDD.n2315 VDD.n896 99.5127
R21654 VDD.n2315 VDD.n894 99.5127
R21655 VDD.n2319 VDD.n894 99.5127
R21656 VDD.n2319 VDD.n885 99.5127
R21657 VDD.n2327 VDD.n885 99.5127
R21658 VDD.n2327 VDD.n883 99.5127
R21659 VDD.n2331 VDD.n883 99.5127
R21660 VDD.n2331 VDD.n873 99.5127
R21661 VDD.n2339 VDD.n873 99.5127
R21662 VDD.n2339 VDD.n871 99.5127
R21663 VDD.n2343 VDD.n871 99.5127
R21664 VDD.n2343 VDD.n861 99.5127
R21665 VDD.n2351 VDD.n861 99.5127
R21666 VDD.n2351 VDD.n859 99.5127
R21667 VDD.n2355 VDD.n859 99.5127
R21668 VDD.n2355 VDD.n849 99.5127
R21669 VDD.n2363 VDD.n849 99.5127
R21670 VDD.n2363 VDD.n847 99.5127
R21671 VDD.n2367 VDD.n847 99.5127
R21672 VDD.n2367 VDD.n837 99.5127
R21673 VDD.n2375 VDD.n837 99.5127
R21674 VDD.n2375 VDD.n835 99.5127
R21675 VDD.n2379 VDD.n835 99.5127
R21676 VDD.n2379 VDD.n825 99.5127
R21677 VDD.n2387 VDD.n825 99.5127
R21678 VDD.n2387 VDD.n823 99.5127
R21679 VDD.n2391 VDD.n823 99.5127
R21680 VDD.n2391 VDD.n813 99.5127
R21681 VDD.n2399 VDD.n813 99.5127
R21682 VDD.n2399 VDD.n811 99.5127
R21683 VDD.n2403 VDD.n811 99.5127
R21684 VDD.n2403 VDD.n801 99.5127
R21685 VDD.n2411 VDD.n801 99.5127
R21686 VDD.n2411 VDD.n799 99.5127
R21687 VDD.n2415 VDD.n799 99.5127
R21688 VDD.n2415 VDD.n789 99.5127
R21689 VDD.n2423 VDD.n789 99.5127
R21690 VDD.n2423 VDD.n787 99.5127
R21691 VDD.n2427 VDD.n787 99.5127
R21692 VDD.n2427 VDD.n777 99.5127
R21693 VDD.n2435 VDD.n777 99.5127
R21694 VDD.n2435 VDD.n775 99.5127
R21695 VDD.n2439 VDD.n775 99.5127
R21696 VDD.n2439 VDD.n766 99.5127
R21697 VDD.n2447 VDD.n766 99.5127
R21698 VDD.n2447 VDD.n764 99.5127
R21699 VDD.n2451 VDD.n764 99.5127
R21700 VDD.n2451 VDD.n754 99.5127
R21701 VDD.n2459 VDD.n754 99.5127
R21702 VDD.n2459 VDD.n751 99.5127
R21703 VDD.n2501 VDD.n751 99.5127
R21704 VDD.n2501 VDD.n752 99.5127
R21705 VDD.n752 VDD.n744 99.5127
R21706 VDD.n2496 VDD.n744 99.5127
R21707 VDD.n2496 VDD.n733 99.5127
R21708 VDD.n2493 VDD.n733 99.5127
R21709 VDD.n1397 VDD.n1396 79.7096
R21710 VDD.n1421 VDD.n1420 79.7096
R21711 VDD.n291 VDD.n290 79.7096
R21712 VDD.n306 VDD.n305 79.7096
R21713 VDD.n98 VDD.n97 79.7096
R21714 VDD.n108 VDD.n107 79.7096
R21715 VDD.n1193 VDD.n1192 79.7096
R21716 VDD.n1180 VDD.n1179 79.7096
R21717 VDD.n2098 VDD.n1108 72.8958
R21718 VDD.n2096 VDD.n1108 72.8958
R21719 VDD.n2090 VDD.n1108 72.8958
R21720 VDD.n2088 VDD.n1108 72.8958
R21721 VDD.n2081 VDD.n1108 72.8958
R21722 VDD.n2079 VDD.n1108 72.8958
R21723 VDD.n2072 VDD.n1108 72.8958
R21724 VDD.n2070 VDD.n1108 72.8958
R21725 VDD.n2557 VDD.n2556 72.8958
R21726 VDD.n2557 VDD.n725 72.8958
R21727 VDD.n2557 VDD.n724 72.8958
R21728 VDD.n2557 VDD.n723 72.8958
R21729 VDD.n2557 VDD.n722 72.8958
R21730 VDD.n2557 VDD.n721 72.8958
R21731 VDD.n2557 VDD.n720 72.8958
R21732 VDD.n2557 VDD.n719 72.8958
R21733 VDD.n3006 VDD.n2558 72.8958
R21734 VDD.n3004 VDD.n2558 72.8958
R21735 VDD.n2998 VDD.n2558 72.8958
R21736 VDD.n2996 VDD.n2558 72.8958
R21737 VDD.n2990 VDD.n2558 72.8958
R21738 VDD.n2988 VDD.n2558 72.8958
R21739 VDD.n2981 VDD.n2558 72.8958
R21740 VDD.n2979 VDD.n2558 72.8958
R21741 VDD.n3449 VDD.n311 72.8958
R21742 VDD.n317 VDD.n311 72.8958
R21743 VDD.n3457 VDD.n311 72.8958
R21744 VDD.n3460 VDD.n311 72.8958
R21745 VDD.n3374 VDD.n311 72.8958
R21746 VDD.n3379 VDD.n311 72.8958
R21747 VDD.n3373 VDD.n311 72.8958
R21748 VDD.n3386 VDD.n311 72.8958
R21749 VDD.n1145 VDD.n1108 72.8958
R21750 VDD.n1148 VDD.n1108 72.8958
R21751 VDD.n1154 VDD.n1108 72.8958
R21752 VDD.n1156 VDD.n1108 72.8958
R21753 VDD.n1701 VDD.n1108 72.8958
R21754 VDD.n1703 VDD.n1108 72.8958
R21755 VDD.n1710 VDD.n1108 72.8958
R21756 VDD.n2557 VDD.n718 72.8958
R21757 VDD.n2557 VDD.n717 72.8958
R21758 VDD.n2557 VDD.n716 72.8958
R21759 VDD.n2557 VDD.n715 72.8958
R21760 VDD.n2557 VDD.n714 72.8958
R21761 VDD.n2557 VDD.n713 72.8958
R21762 VDD.n2557 VDD.n712 72.8958
R21763 VDD.n2557 VDD.n711 72.8958
R21764 VDD.n2568 VDD.n2558 72.8958
R21765 VDD.n2574 VDD.n2558 72.8958
R21766 VDD.n2576 VDD.n2558 72.8958
R21767 VDD.n2582 VDD.n2558 72.8958
R21768 VDD.n2584 VDD.n2558 72.8958
R21769 VDD.n2593 VDD.n2558 72.8958
R21770 VDD.n2596 VDD.n2558 72.8958
R21771 VDD.n3409 VDD.n311 72.8958
R21772 VDD.n3416 VDD.n311 72.8958
R21773 VDD.n338 VDD.n311 72.8958
R21774 VDD.n3423 VDD.n311 72.8958
R21775 VDD.n3427 VDD.n311 72.8958
R21776 VDD.n332 VDD.n311 72.8958
R21777 VDD.n3434 VDD.n311 72.8958
R21778 VDD.n3437 VDD.n311 72.8958
R21779 VDD.n3519 VDD.n3518 66.2847
R21780 VDD.n3518 VDD.n264 66.2847
R21781 VDD.n3518 VDD.n265 66.2847
R21782 VDD.n3518 VDD.n266 66.2847
R21783 VDD.n3518 VDD.n267 66.2847
R21784 VDD.n3518 VDD.n268 66.2847
R21785 VDD.n3518 VDD.n269 66.2847
R21786 VDD.n3518 VDD.n270 66.2847
R21787 VDD.n3518 VDD.n271 66.2847
R21788 VDD.n3518 VDD.n272 66.2847
R21789 VDD.n3518 VDD.n273 66.2847
R21790 VDD.n3518 VDD.n274 66.2847
R21791 VDD.n3518 VDD.n275 66.2847
R21792 VDD.n3663 VDD.n3662 66.2847
R21793 VDD.n3663 VDD.n95 66.2847
R21794 VDD.n3663 VDD.n94 66.2847
R21795 VDD.n3663 VDD.n93 66.2847
R21796 VDD.n3663 VDD.n92 66.2847
R21797 VDD.n3663 VDD.n91 66.2847
R21798 VDD.n3663 VDD.n90 66.2847
R21799 VDD.n3663 VDD.n89 66.2847
R21800 VDD.n3663 VDD.n88 66.2847
R21801 VDD.n3663 VDD.n87 66.2847
R21802 VDD.n3663 VDD.n86 66.2847
R21803 VDD.n3663 VDD.n85 66.2847
R21804 VDD.n3663 VDD.n84 66.2847
R21805 VDD.n3663 VDD.n83 66.2847
R21806 VDD.n1672 VDD.n1671 66.2847
R21807 VDD.n1671 VDD.n1670 66.2847
R21808 VDD.n1671 VDD.n1668 66.2847
R21809 VDD.n1671 VDD.n1667 66.2847
R21810 VDD.n1671 VDD.n1665 66.2847
R21811 VDD.n1671 VDD.n1664 66.2847
R21812 VDD.n1671 VDD.n1662 66.2847
R21813 VDD.n1671 VDD.n1661 66.2847
R21814 VDD.n1671 VDD.n1189 66.2847
R21815 VDD.n1671 VDD.n1188 66.2847
R21816 VDD.n1671 VDD.n1187 66.2847
R21817 VDD.n1671 VDD.n1186 66.2847
R21818 VDD.n1671 VDD.n1185 66.2847
R21819 VDD.n1671 VDD.n1184 66.2847
R21820 VDD.n1441 VDD.n1440 66.2847
R21821 VDD.n1440 VDD.n1346 66.2847
R21822 VDD.n1440 VDD.n1347 66.2847
R21823 VDD.n1440 VDD.n1348 66.2847
R21824 VDD.n1440 VDD.n1349 66.2847
R21825 VDD.n1440 VDD.n1350 66.2847
R21826 VDD.n1440 VDD.n1351 66.2847
R21827 VDD.n1440 VDD.n1352 66.2847
R21828 VDD.n1440 VDD.n1353 66.2847
R21829 VDD.n1440 VDD.n1354 66.2847
R21830 VDD.n1440 VDD.n1355 66.2847
R21831 VDD.n1440 VDD.n1356 66.2847
R21832 VDD.n1440 VDD.n1357 66.2847
R21833 VDD.n120 VDD.n83 52.4337
R21834 VDD.n126 VDD.n84 52.4337
R21835 VDD.n130 VDD.n85 52.4337
R21836 VDD.n136 VDD.n86 52.4337
R21837 VDD.n140 VDD.n87 52.4337
R21838 VDD.n145 VDD.n88 52.4337
R21839 VDD.n149 VDD.n89 52.4337
R21840 VDD.n155 VDD.n90 52.4337
R21841 VDD.n159 VDD.n91 52.4337
R21842 VDD.n165 VDD.n92 52.4337
R21843 VDD.n169 VDD.n93 52.4337
R21844 VDD.n175 VDD.n94 52.4337
R21845 VDD.n178 VDD.n95 52.4337
R21846 VDD.n3662 VDD.n3661 52.4337
R21847 VDD.n3520 VDD.n3519 52.4337
R21848 VDD.n277 VDD.n264 52.4337
R21849 VDD.n3512 VDD.n265 52.4337
R21850 VDD.n3508 VDD.n266 52.4337
R21851 VDD.n3504 VDD.n267 52.4337
R21852 VDD.n3500 VDD.n268 52.4337
R21853 VDD.n3496 VDD.n269 52.4337
R21854 VDD.n3493 VDD.n270 52.4337
R21855 VDD.n3489 VDD.n271 52.4337
R21856 VDD.n3485 VDD.n272 52.4337
R21857 VDD.n3481 VDD.n273 52.4337
R21858 VDD.n3477 VDD.n274 52.4337
R21859 VDD.n3473 VDD.n275 52.4337
R21860 VDD.n3519 VDD.n263 52.4337
R21861 VDD.n3513 VDD.n264 52.4337
R21862 VDD.n3509 VDD.n265 52.4337
R21863 VDD.n3505 VDD.n266 52.4337
R21864 VDD.n3501 VDD.n267 52.4337
R21865 VDD.n288 VDD.n268 52.4337
R21866 VDD.n3494 VDD.n269 52.4337
R21867 VDD.n3490 VDD.n270 52.4337
R21868 VDD.n3486 VDD.n271 52.4337
R21869 VDD.n3482 VDD.n272 52.4337
R21870 VDD.n3478 VDD.n273 52.4337
R21871 VDD.n3474 VDD.n274 52.4337
R21872 VDD.n304 VDD.n275 52.4337
R21873 VDD.n3662 VDD.n96 52.4337
R21874 VDD.n176 VDD.n95 52.4337
R21875 VDD.n168 VDD.n94 52.4337
R21876 VDD.n166 VDD.n93 52.4337
R21877 VDD.n158 VDD.n92 52.4337
R21878 VDD.n156 VDD.n91 52.4337
R21879 VDD.n148 VDD.n90 52.4337
R21880 VDD.n109 VDD.n89 52.4337
R21881 VDD.n139 VDD.n88 52.4337
R21882 VDD.n137 VDD.n87 52.4337
R21883 VDD.n129 VDD.n86 52.4337
R21884 VDD.n127 VDD.n85 52.4337
R21885 VDD.n119 VDD.n84 52.4337
R21886 VDD.n117 VDD.n83 52.4337
R21887 VDD.n1632 VDD.n1184 52.4337
R21888 VDD.n1637 VDD.n1185 52.4337
R21889 VDD.n1201 VDD.n1186 52.4337
R21890 VDD.n1645 VDD.n1187 52.4337
R21891 VDD.n1197 VDD.n1188 52.4337
R21892 VDD.n1653 VDD.n1189 52.4337
R21893 VDD.n1661 VDD.n1659 52.4337
R21894 VDD.n1662 VDD.n1164 52.4337
R21895 VDD.n1664 VDD.n1166 52.4337
R21896 VDD.n1665 VDD.n1169 52.4337
R21897 VDD.n1667 VDD.n1171 52.4337
R21898 VDD.n1668 VDD.n1174 52.4337
R21899 VDD.n1670 VDD.n1176 52.4337
R21900 VDD.n1672 VDD.n1181 52.4337
R21901 VDD.n1673 VDD.n1672 52.4337
R21902 VDD.n1670 VDD.n1669 52.4337
R21903 VDD.n1668 VDD.n1175 52.4337
R21904 VDD.n1667 VDD.n1666 52.4337
R21905 VDD.n1665 VDD.n1170 52.4337
R21906 VDD.n1664 VDD.n1663 52.4337
R21907 VDD.n1662 VDD.n1165 52.4337
R21908 VDD.n1661 VDD.n1660 52.4337
R21909 VDD.n1190 VDD.n1189 52.4337
R21910 VDD.n1652 VDD.n1188 52.4337
R21911 VDD.n1196 VDD.n1187 52.4337
R21912 VDD.n1644 VDD.n1186 52.4337
R21913 VDD.n1200 VDD.n1185 52.4337
R21914 VDD.n1636 VDD.n1184 52.4337
R21915 VDD.n1442 VDD.n1441 52.4337
R21916 VDD.n1359 VDD.n1346 52.4337
R21917 VDD.n1363 VDD.n1347 52.4337
R21918 VDD.n1365 VDD.n1348 52.4337
R21919 VDD.n1369 VDD.n1349 52.4337
R21920 VDD.n1371 VDD.n1350 52.4337
R21921 VDD.n1418 VDD.n1351 52.4337
R21922 VDD.n1375 VDD.n1352 52.4337
R21923 VDD.n1379 VDD.n1353 52.4337
R21924 VDD.n1381 VDD.n1354 52.4337
R21925 VDD.n1385 VDD.n1355 52.4337
R21926 VDD.n1387 VDD.n1356 52.4337
R21927 VDD.n1391 VDD.n1357 52.4337
R21928 VDD.n1441 VDD.n1345 52.4337
R21929 VDD.n1362 VDD.n1346 52.4337
R21930 VDD.n1364 VDD.n1347 52.4337
R21931 VDD.n1368 VDD.n1348 52.4337
R21932 VDD.n1370 VDD.n1349 52.4337
R21933 VDD.n1419 VDD.n1350 52.4337
R21934 VDD.n1374 VDD.n1351 52.4337
R21935 VDD.n1378 VDD.n1352 52.4337
R21936 VDD.n1380 VDD.n1353 52.4337
R21937 VDD.n1384 VDD.n1354 52.4337
R21938 VDD.n1386 VDD.n1355 52.4337
R21939 VDD.n1390 VDD.n1356 52.4337
R21940 VDD.n1395 VDD.n1357 52.4337
R21941 VDD.n3437 VDD.n3436 39.2114
R21942 VDD.n3434 VDD.n3433 39.2114
R21943 VDD.n3429 VDD.n332 39.2114
R21944 VDD.n3427 VDD.n3426 39.2114
R21945 VDD.n3423 VDD.n3422 39.2114
R21946 VDD.n3418 VDD.n338 39.2114
R21947 VDD.n3416 VDD.n3415 39.2114
R21948 VDD.n3411 VDD.n3409 39.2114
R21949 VDD.n2568 VDD.n709 39.2114
R21950 VDD.n2574 VDD.n2573 39.2114
R21951 VDD.n2577 VDD.n2576 39.2114
R21952 VDD.n2582 VDD.n2581 39.2114
R21953 VDD.n2585 VDD.n2584 39.2114
R21954 VDD.n2593 VDD.n2592 39.2114
R21955 VDD.n2596 VDD.n2595 39.2114
R21956 VDD.n2543 VDD.n711 39.2114
R21957 VDD.n2539 VDD.n712 39.2114
R21958 VDD.n2535 VDD.n713 39.2114
R21959 VDD.n2531 VDD.n714 39.2114
R21960 VDD.n2527 VDD.n715 39.2114
R21961 VDD.n2523 VDD.n716 39.2114
R21962 VDD.n2519 VDD.n717 39.2114
R21963 VDD.n2515 VDD.n718 39.2114
R21964 VDD.n1145 VDD.n1107 39.2114
R21965 VDD.n1149 VDD.n1148 39.2114
R21966 VDD.n1154 VDD.n1153 39.2114
R21967 VDD.n1157 VDD.n1156 39.2114
R21968 VDD.n1701 VDD.n1700 39.2114
R21969 VDD.n1704 VDD.n1703 39.2114
R21970 VDD.n1710 VDD.n1709 39.2114
R21971 VDD.n3386 VDD.n3385 39.2114
R21972 VDD.n3381 VDD.n3373 39.2114
R21973 VDD.n3379 VDD.n3378 39.2114
R21974 VDD.n3374 VDD.n310 39.2114
R21975 VDD.n3460 VDD.n3459 39.2114
R21976 VDD.n3457 VDD.n3456 39.2114
R21977 VDD.n3451 VDD.n317 39.2114
R21978 VDD.n3449 VDD.n3448 39.2114
R21979 VDD.n3006 VDD.n2783 39.2114
R21980 VDD.n3005 VDD.n3004 39.2114
R21981 VDD.n2998 VDD.n2785 39.2114
R21982 VDD.n2997 VDD.n2996 39.2114
R21983 VDD.n2990 VDD.n2787 39.2114
R21984 VDD.n2989 VDD.n2988 39.2114
R21985 VDD.n2981 VDD.n2789 39.2114
R21986 VDD.n2980 VDD.n2979 39.2114
R21987 VDD.n2489 VDD.n719 39.2114
R21988 VDD.n2485 VDD.n720 39.2114
R21989 VDD.n2481 VDD.n721 39.2114
R21990 VDD.n2477 VDD.n722 39.2114
R21991 VDD.n2473 VDD.n723 39.2114
R21992 VDD.n2469 VDD.n724 39.2114
R21993 VDD.n2465 VDD.n725 39.2114
R21994 VDD.n2556 VDD.n2555 39.2114
R21995 VDD.n2098 VDD.n1111 39.2114
R21996 VDD.n2097 VDD.n2096 39.2114
R21997 VDD.n2090 VDD.n1113 39.2114
R21998 VDD.n2089 VDD.n2088 39.2114
R21999 VDD.n2081 VDD.n1115 39.2114
R22000 VDD.n2080 VDD.n2079 39.2114
R22001 VDD.n2072 VDD.n1118 39.2114
R22002 VDD.n2071 VDD.n2070 39.2114
R22003 VDD.n2099 VDD.n2098 39.2114
R22004 VDD.n2096 VDD.n2095 39.2114
R22005 VDD.n2091 VDD.n2090 39.2114
R22006 VDD.n2088 VDD.n2087 39.2114
R22007 VDD.n2082 VDD.n2081 39.2114
R22008 VDD.n2079 VDD.n2078 39.2114
R22009 VDD.n2073 VDD.n2072 39.2114
R22010 VDD.n2070 VDD.n2069 39.2114
R22011 VDD.n2556 VDD.n726 39.2114
R22012 VDD.n2468 VDD.n725 39.2114
R22013 VDD.n2472 VDD.n724 39.2114
R22014 VDD.n2476 VDD.n723 39.2114
R22015 VDD.n2480 VDD.n722 39.2114
R22016 VDD.n2484 VDD.n721 39.2114
R22017 VDD.n2488 VDD.n720 39.2114
R22018 VDD.n2492 VDD.n719 39.2114
R22019 VDD.n3007 VDD.n3006 39.2114
R22020 VDD.n3004 VDD.n3003 39.2114
R22021 VDD.n2999 VDD.n2998 39.2114
R22022 VDD.n2996 VDD.n2995 39.2114
R22023 VDD.n2991 VDD.n2990 39.2114
R22024 VDD.n2988 VDD.n2987 39.2114
R22025 VDD.n2982 VDD.n2981 39.2114
R22026 VDD.n2979 VDD.n2978 39.2114
R22027 VDD.n3450 VDD.n3449 39.2114
R22028 VDD.n317 VDD.n313 39.2114
R22029 VDD.n3458 VDD.n3457 39.2114
R22030 VDD.n3461 VDD.n3460 39.2114
R22031 VDD.n3375 VDD.n3374 39.2114
R22032 VDD.n3380 VDD.n3379 39.2114
R22033 VDD.n3373 VDD.n3371 39.2114
R22034 VDD.n3387 VDD.n3386 39.2114
R22035 VDD.n1146 VDD.n1145 39.2114
R22036 VDD.n1148 VDD.n1142 39.2114
R22037 VDD.n1155 VDD.n1154 39.2114
R22038 VDD.n1156 VDD.n1140 39.2114
R22039 VDD.n1702 VDD.n1701 39.2114
R22040 VDD.n1703 VDD.n1136 39.2114
R22041 VDD.n1711 VDD.n1710 39.2114
R22042 VDD.n2518 VDD.n718 39.2114
R22043 VDD.n2522 VDD.n717 39.2114
R22044 VDD.n2526 VDD.n716 39.2114
R22045 VDD.n2530 VDD.n715 39.2114
R22046 VDD.n2534 VDD.n714 39.2114
R22047 VDD.n2538 VDD.n713 39.2114
R22048 VDD.n2542 VDD.n712 39.2114
R22049 VDD.n2545 VDD.n711 39.2114
R22050 VDD.n2569 VDD.n2568 39.2114
R22051 VDD.n2575 VDD.n2574 39.2114
R22052 VDD.n2576 VDD.n2565 39.2114
R22053 VDD.n2583 VDD.n2582 39.2114
R22054 VDD.n2584 VDD.n2563 39.2114
R22055 VDD.n2594 VDD.n2593 39.2114
R22056 VDD.n2597 VDD.n2596 39.2114
R22057 VDD.n3409 VDD.n340 39.2114
R22058 VDD.n3417 VDD.n3416 39.2114
R22059 VDD.n338 VDD.n334 39.2114
R22060 VDD.n3424 VDD.n3423 39.2114
R22061 VDD.n3428 VDD.n3427 39.2114
R22062 VDD.n332 VDD.n330 39.2114
R22063 VDD.n3435 VDD.n3434 39.2114
R22064 VDD.n3438 VDD.n3437 39.2114
R22065 VDD.n1440 VDD.n1340 32.9976
R22066 VDD.n1671 VDD.n1183 32.9976
R22067 VDD.n3518 VDD.n256 32.9976
R22068 VDD.n3664 VDD.n3663 32.9976
R22069 VDD.n2780 VDD.n2599 32.781
R22070 VDD.n3412 VDD.n3408 32.781
R22071 VDD.n3014 VDD.n708 32.781
R22072 VDD.n3440 VDD.n3439 32.781
R22073 VDD.n3389 VDD.n3370 32.781
R22074 VDD.n3447 VDD.n3446 32.781
R22075 VDD.n2977 VDD.n2976 32.781
R22076 VDD.n3010 VDD.n3009 32.781
R22077 VDD.n2106 VDD.n1106 32.781
R22078 VDD.n2547 VDD.n2546 32.781
R22079 VDD.n2516 VDD.n2513 32.781
R22080 VDD.n1714 VDD.n1713 32.781
R22081 VDD.n2494 VDD.n2491 32.781
R22082 VDD.n2554 VDD.n2553 32.781
R22083 VDD.n2068 VDD.n2067 32.781
R22084 VDD.n2102 VDD.n2101 32.781
R22085 VDD.n7 VDD.t103 31.2553
R22086 VDD.n7 VDD.t87 31.2553
R22087 VDD.n8 VDD.t106 31.2553
R22088 VDD.n8 VDD.t89 31.2553
R22089 VDD.n10 VDD.t75 31.2553
R22090 VDD.n10 VDD.t101 31.2553
R22091 VDD.n12 VDD.t94 31.2553
R22092 VDD.n12 VDD.t108 31.2553
R22093 VDD.n5 VDD.t72 31.2553
R22094 VDD.n5 VDD.t82 31.2553
R22095 VDD.n3 VDD.t85 31.2553
R22096 VDD.n3 VDD.t97 31.2553
R22097 VDD.n1 VDD.t70 31.2553
R22098 VDD.n1 VDD.t80 31.2553
R22099 VDD.n0 VDD.t99 31.2553
R22100 VDD.n0 VDD.t77 31.2553
R22101 VDD.n1398 VDD.n1397 30.8369
R22102 VDD.n1422 VDD.n1421 30.8369
R22103 VDD.n3498 VDD.n291 30.8369
R22104 VDD.n307 VDD.n306 30.8369
R22105 VDD.n99 VDD.n98 30.8369
R22106 VDD.n147 VDD.n108 30.8369
R22107 VDD.n1658 VDD.n1193 30.8369
R22108 VDD.n1675 VDD.n1180 30.8369
R22109 VDD.n2104 VDD.n1108 24.3037
R22110 VDD.n2557 VDD.n710 24.3037
R22111 VDD.n3012 VDD.n2558 24.3037
R22112 VDD.n323 VDD.n311 24.3037
R22113 VDD.n2985 VDD.n2791 24.049
R22114 VDD.n337 VDD.n336 24.049
R22115 VDD.n2590 VDD.n2589 24.049
R22116 VDD.n3454 VDD.n315 24.049
R22117 VDD.n2076 VDD.n1120 24.049
R22118 VDD.n1706 VDD.n1138 24.049
R22119 VDD.n739 VDD.n738 24.049
R22120 VDD.n2464 VDD.n2463 24.049
R22121 VDD.n1449 VDD.n1340 19.7592
R22122 VDD.n1449 VDD.n1334 19.7592
R22123 VDD.n1457 VDD.n1334 19.7592
R22124 VDD.n1457 VDD.n1328 19.7592
R22125 VDD.n1465 VDD.n1328 19.7592
R22126 VDD.n1473 VDD.n1322 19.7592
R22127 VDD.n1473 VDD.n1316 19.7592
R22128 VDD.n1481 VDD.n1316 19.7592
R22129 VDD.n1481 VDD.n1310 19.7592
R22130 VDD.n1489 VDD.n1310 19.7592
R22131 VDD.n1489 VDD.n1304 19.7592
R22132 VDD.n1497 VDD.n1304 19.7592
R22133 VDD.n1497 VDD.n1298 19.7592
R22134 VDD.n1505 VDD.n1298 19.7592
R22135 VDD.n1505 VDD.n1292 19.7592
R22136 VDD.n1513 VDD.n1292 19.7592
R22137 VDD.n1521 VDD.n1286 19.7592
R22138 VDD.n1521 VDD.n1280 19.7592
R22139 VDD.n1530 VDD.n1280 19.7592
R22140 VDD.n1530 VDD.n1274 19.7592
R22141 VDD.n1538 VDD.n1274 19.7592
R22142 VDD.n1538 VDD.n1264 19.7592
R22143 VDD.n1546 VDD.n1264 19.7592
R22144 VDD.n1546 VDD.n1258 19.7592
R22145 VDD.n1554 VDD.n1258 19.7592
R22146 VDD.n1562 VDD.n1252 19.7592
R22147 VDD.n1562 VDD.n1246 19.7592
R22148 VDD.n1570 VDD.n1246 19.7592
R22149 VDD.n1570 VDD.n1240 19.7592
R22150 VDD.n1578 VDD.n1240 19.7592
R22151 VDD.n1578 VDD.n1234 19.7592
R22152 VDD.n1586 VDD.n1234 19.7592
R22153 VDD.n1586 VDD.n1228 19.7592
R22154 VDD.n1594 VDD.n1228 19.7592
R22155 VDD.n1594 VDD.n1221 19.7592
R22156 VDD.n1603 VDD.n1221 19.7592
R22157 VDD.n1611 VDD.n1215 19.7592
R22158 VDD.n1611 VDD.n1208 19.7592
R22159 VDD.n1624 VDD.n1208 19.7592
R22160 VDD.n1624 VDD.n1623 19.7592
R22161 VDD.n1623 VDD.n1183 19.7592
R22162 VDD.n3529 VDD.n256 19.7592
R22163 VDD.n3529 VDD.n250 19.7592
R22164 VDD.n3537 VDD.n250 19.7592
R22165 VDD.n3537 VDD.n244 19.7592
R22166 VDD.n3545 VDD.n244 19.7592
R22167 VDD.n3553 VDD.n238 19.7592
R22168 VDD.n3553 VDD.n232 19.7592
R22169 VDD.n3561 VDD.n232 19.7592
R22170 VDD.n3561 VDD.n226 19.7592
R22171 VDD.n3569 VDD.n226 19.7592
R22172 VDD.n3569 VDD.n220 19.7592
R22173 VDD.n3577 VDD.n220 19.7592
R22174 VDD.n3577 VDD.n214 19.7592
R22175 VDD.n3587 VDD.n214 19.7592
R22176 VDD.n3587 VDD.n208 19.7592
R22177 VDD.n3595 VDD.n208 19.7592
R22178 VDD.n3608 VDD.n202 19.7592
R22179 VDD.n3608 VDD.n3607 19.7592
R22180 VDD.n3607 VDD.n196 19.7592
R22181 VDD.n3617 VDD.n196 19.7592
R22182 VDD.n3617 VDD.n25 19.7592
R22183 VDD.n3705 VDD.n25 19.7592
R22184 VDD.n3705 VDD.n3704 19.7592
R22185 VDD.n3704 VDD.n3703 19.7592
R22186 VDD.n3703 VDD.n29 19.7592
R22187 VDD.n3697 VDD.n3696 19.7592
R22188 VDD.n3696 VDD.n3695 19.7592
R22189 VDD.n3695 VDD.n40 19.7592
R22190 VDD.n3689 VDD.n40 19.7592
R22191 VDD.n3689 VDD.n3688 19.7592
R22192 VDD.n3688 VDD.n3687 19.7592
R22193 VDD.n3687 VDD.n51 19.7592
R22194 VDD.n3681 VDD.n51 19.7592
R22195 VDD.n3681 VDD.n3680 19.7592
R22196 VDD.n3680 VDD.n3679 19.7592
R22197 VDD.n3679 VDD.n62 19.7592
R22198 VDD.n3673 VDD.n3672 19.7592
R22199 VDD.n3672 VDD.n3671 19.7592
R22200 VDD.n3671 VDD.n73 19.7592
R22201 VDD.n3665 VDD.n73 19.7592
R22202 VDD.n3665 VDD.n3664 19.7592
R22203 VDD.n1417 VDD.n1416 19.3944
R22204 VDD.n1416 VDD.n1376 19.3944
R22205 VDD.n1412 VDD.n1376 19.3944
R22206 VDD.n1412 VDD.n1411 19.3944
R22207 VDD.n1411 VDD.n1410 19.3944
R22208 VDD.n1410 VDD.n1382 19.3944
R22209 VDD.n1406 VDD.n1382 19.3944
R22210 VDD.n1406 VDD.n1405 19.3944
R22211 VDD.n1405 VDD.n1404 19.3944
R22212 VDD.n1404 VDD.n1388 19.3944
R22213 VDD.n1400 VDD.n1388 19.3944
R22214 VDD.n1400 VDD.n1399 19.3944
R22215 VDD.n1443 VDD.n1344 19.3944
R22216 VDD.n1438 VDD.n1344 19.3944
R22217 VDD.n1438 VDD.n1360 19.3944
R22218 VDD.n1434 VDD.n1360 19.3944
R22219 VDD.n1434 VDD.n1433 19.3944
R22220 VDD.n1433 VDD.n1432 19.3944
R22221 VDD.n1432 VDD.n1366 19.3944
R22222 VDD.n1428 VDD.n1366 19.3944
R22223 VDD.n1428 VDD.n1427 19.3944
R22224 VDD.n1427 VDD.n1426 19.3944
R22225 VDD.n1426 VDD.n1372 19.3944
R22226 VDD.n1451 VDD.n1338 19.3944
R22227 VDD.n1451 VDD.n1336 19.3944
R22228 VDD.n1455 VDD.n1336 19.3944
R22229 VDD.n1455 VDD.n1326 19.3944
R22230 VDD.n1467 VDD.n1326 19.3944
R22231 VDD.n1467 VDD.n1324 19.3944
R22232 VDD.n1471 VDD.n1324 19.3944
R22233 VDD.n1471 VDD.n1314 19.3944
R22234 VDD.n1483 VDD.n1314 19.3944
R22235 VDD.n1483 VDD.n1312 19.3944
R22236 VDD.n1487 VDD.n1312 19.3944
R22237 VDD.n1487 VDD.n1302 19.3944
R22238 VDD.n1499 VDD.n1302 19.3944
R22239 VDD.n1499 VDD.n1300 19.3944
R22240 VDD.n1503 VDD.n1300 19.3944
R22241 VDD.n1503 VDD.n1290 19.3944
R22242 VDD.n1515 VDD.n1290 19.3944
R22243 VDD.n1515 VDD.n1288 19.3944
R22244 VDD.n1519 VDD.n1288 19.3944
R22245 VDD.n1519 VDD.n1278 19.3944
R22246 VDD.n1532 VDD.n1278 19.3944
R22247 VDD.n1532 VDD.n1276 19.3944
R22248 VDD.n1536 VDD.n1276 19.3944
R22249 VDD.n1536 VDD.n1262 19.3944
R22250 VDD.n1548 VDD.n1262 19.3944
R22251 VDD.n1548 VDD.n1260 19.3944
R22252 VDD.n1552 VDD.n1260 19.3944
R22253 VDD.n1552 VDD.n1250 19.3944
R22254 VDD.n1564 VDD.n1250 19.3944
R22255 VDD.n1564 VDD.n1248 19.3944
R22256 VDD.n1568 VDD.n1248 19.3944
R22257 VDD.n1568 VDD.n1238 19.3944
R22258 VDD.n1580 VDD.n1238 19.3944
R22259 VDD.n1580 VDD.n1236 19.3944
R22260 VDD.n1584 VDD.n1236 19.3944
R22261 VDD.n1584 VDD.n1226 19.3944
R22262 VDD.n1596 VDD.n1226 19.3944
R22263 VDD.n1596 VDD.n1223 19.3944
R22264 VDD.n1601 VDD.n1223 19.3944
R22265 VDD.n1601 VDD.n1224 19.3944
R22266 VDD.n1224 VDD.n1213 19.3944
R22267 VDD.n1614 VDD.n1213 19.3944
R22268 VDD.n1614 VDD.n1210 19.3944
R22269 VDD.n1621 VDD.n1210 19.3944
R22270 VDD.n1621 VDD.n1211 19.3944
R22271 VDD.n3521 VDD.n262 19.3944
R22272 VDD.n3516 VDD.n262 19.3944
R22273 VDD.n3516 VDD.n3515 19.3944
R22274 VDD.n3515 VDD.n3514 19.3944
R22275 VDD.n3514 VDD.n3511 19.3944
R22276 VDD.n3511 VDD.n3510 19.3944
R22277 VDD.n3510 VDD.n3507 19.3944
R22278 VDD.n3507 VDD.n3506 19.3944
R22279 VDD.n3506 VDD.n3503 19.3944
R22280 VDD.n3503 VDD.n3502 19.3944
R22281 VDD.n3502 VDD.n3499 19.3944
R22282 VDD.n3497 VDD.n3495 19.3944
R22283 VDD.n3495 VDD.n3492 19.3944
R22284 VDD.n3492 VDD.n3491 19.3944
R22285 VDD.n3491 VDD.n3488 19.3944
R22286 VDD.n3488 VDD.n3487 19.3944
R22287 VDD.n3487 VDD.n3484 19.3944
R22288 VDD.n3484 VDD.n3483 19.3944
R22289 VDD.n3483 VDD.n3480 19.3944
R22290 VDD.n3480 VDD.n3479 19.3944
R22291 VDD.n3479 VDD.n3476 19.3944
R22292 VDD.n3476 VDD.n3475 19.3944
R22293 VDD.n3475 VDD.n3472 19.3944
R22294 VDD.n3527 VDD.n258 19.3944
R22295 VDD.n3527 VDD.n248 19.3944
R22296 VDD.n3539 VDD.n248 19.3944
R22297 VDD.n3539 VDD.n246 19.3944
R22298 VDD.n3543 VDD.n246 19.3944
R22299 VDD.n3543 VDD.n236 19.3944
R22300 VDD.n3555 VDD.n236 19.3944
R22301 VDD.n3555 VDD.n234 19.3944
R22302 VDD.n3559 VDD.n234 19.3944
R22303 VDD.n3559 VDD.n224 19.3944
R22304 VDD.n3571 VDD.n224 19.3944
R22305 VDD.n3571 VDD.n222 19.3944
R22306 VDD.n3575 VDD.n222 19.3944
R22307 VDD.n3575 VDD.n212 19.3944
R22308 VDD.n3589 VDD.n212 19.3944
R22309 VDD.n3589 VDD.n210 19.3944
R22310 VDD.n3593 VDD.n210 19.3944
R22311 VDD.n3593 VDD.n200 19.3944
R22312 VDD.n3610 VDD.n200 19.3944
R22313 VDD.n3610 VDD.n198 19.3944
R22314 VDD.n3614 VDD.n198 19.3944
R22315 VDD.n3614 VDD.n21 19.3944
R22316 VDD.n3708 VDD.n21 19.3944
R22317 VDD.n3708 VDD.n3707 19.3944
R22318 VDD.n3707 VDD.n23 19.3944
R22319 VDD.n3701 VDD.n23 19.3944
R22320 VDD.n3701 VDD.n3700 19.3944
R22321 VDD.n3700 VDD.n3699 19.3944
R22322 VDD.n3699 VDD.n35 19.3944
R22323 VDD.n3693 VDD.n35 19.3944
R22324 VDD.n3693 VDD.n3692 19.3944
R22325 VDD.n3692 VDD.n3691 19.3944
R22326 VDD.n3691 VDD.n46 19.3944
R22327 VDD.n3685 VDD.n46 19.3944
R22328 VDD.n3685 VDD.n3684 19.3944
R22329 VDD.n3684 VDD.n3683 19.3944
R22330 VDD.n3683 VDD.n57 19.3944
R22331 VDD.n3677 VDD.n57 19.3944
R22332 VDD.n3677 VDD.n3676 19.3944
R22333 VDD.n3676 VDD.n3675 19.3944
R22334 VDD.n3675 VDD.n68 19.3944
R22335 VDD.n3669 VDD.n68 19.3944
R22336 VDD.n3669 VDD.n3668 19.3944
R22337 VDD.n3668 VDD.n3667 19.3944
R22338 VDD.n3667 VDD.n79 19.3944
R22339 VDD.n150 VDD.n105 19.3944
R22340 VDD.n154 VDD.n105 19.3944
R22341 VDD.n157 VDD.n154 19.3944
R22342 VDD.n160 VDD.n157 19.3944
R22343 VDD.n160 VDD.n103 19.3944
R22344 VDD.n164 VDD.n103 19.3944
R22345 VDD.n167 VDD.n164 19.3944
R22346 VDD.n170 VDD.n167 19.3944
R22347 VDD.n170 VDD.n101 19.3944
R22348 VDD.n174 VDD.n101 19.3944
R22349 VDD.n177 VDD.n174 19.3944
R22350 VDD.n179 VDD.n177 19.3944
R22351 VDD.n121 VDD.n118 19.3944
R22352 VDD.n121 VDD.n114 19.3944
R22353 VDD.n125 VDD.n114 19.3944
R22354 VDD.n128 VDD.n125 19.3944
R22355 VDD.n131 VDD.n128 19.3944
R22356 VDD.n131 VDD.n112 19.3944
R22357 VDD.n135 VDD.n112 19.3944
R22358 VDD.n138 VDD.n135 19.3944
R22359 VDD.n141 VDD.n138 19.3944
R22360 VDD.n141 VDD.n110 19.3944
R22361 VDD.n146 VDD.n110 19.3944
R22362 VDD.n3531 VDD.n254 19.3944
R22363 VDD.n3531 VDD.n252 19.3944
R22364 VDD.n3535 VDD.n252 19.3944
R22365 VDD.n3535 VDD.n242 19.3944
R22366 VDD.n3547 VDD.n242 19.3944
R22367 VDD.n3547 VDD.n240 19.3944
R22368 VDD.n3551 VDD.n240 19.3944
R22369 VDD.n3551 VDD.n230 19.3944
R22370 VDD.n3563 VDD.n230 19.3944
R22371 VDD.n3563 VDD.n228 19.3944
R22372 VDD.n3567 VDD.n228 19.3944
R22373 VDD.n3567 VDD.n218 19.3944
R22374 VDD.n3579 VDD.n218 19.3944
R22375 VDD.n3579 VDD.n216 19.3944
R22376 VDD.n3585 VDD.n216 19.3944
R22377 VDD.n3585 VDD.n3584 19.3944
R22378 VDD.n3584 VDD.n206 19.3944
R22379 VDD.n3598 VDD.n206 19.3944
R22380 VDD.n3598 VDD.n204 19.3944
R22381 VDD.n3605 VDD.n204 19.3944
R22382 VDD.n3605 VDD.n3604 19.3944
R22383 VDD.n3604 VDD.n193 19.3944
R22384 VDD.n3620 VDD.n193 19.3944
R22385 VDD.n3621 VDD.n3620 19.3944
R22386 VDD.n3622 VDD.n3621 19.3944
R22387 VDD.n3622 VDD.n191 19.3944
R22388 VDD.n3627 VDD.n191 19.3944
R22389 VDD.n3628 VDD.n3627 19.3944
R22390 VDD.n3629 VDD.n3628 19.3944
R22391 VDD.n3629 VDD.n189 19.3944
R22392 VDD.n3634 VDD.n189 19.3944
R22393 VDD.n3635 VDD.n3634 19.3944
R22394 VDD.n3636 VDD.n3635 19.3944
R22395 VDD.n3636 VDD.n187 19.3944
R22396 VDD.n3641 VDD.n187 19.3944
R22397 VDD.n3642 VDD.n3641 19.3944
R22398 VDD.n3643 VDD.n3642 19.3944
R22399 VDD.n3643 VDD.n185 19.3944
R22400 VDD.n3648 VDD.n185 19.3944
R22401 VDD.n3649 VDD.n3648 19.3944
R22402 VDD.n3650 VDD.n3649 19.3944
R22403 VDD.n3650 VDD.n183 19.3944
R22404 VDD.n3655 VDD.n183 19.3944
R22405 VDD.n3656 VDD.n3655 19.3944
R22406 VDD.n3657 VDD.n3656 19.3944
R22407 VDD.n1635 VDD.n1634 19.3944
R22408 VDD.n1638 VDD.n1635 19.3944
R22409 VDD.n1638 VDD.n1199 19.3944
R22410 VDD.n1642 VDD.n1199 19.3944
R22411 VDD.n1643 VDD.n1642 19.3944
R22412 VDD.n1646 VDD.n1643 19.3944
R22413 VDD.n1646 VDD.n1195 19.3944
R22414 VDD.n1650 VDD.n1195 19.3944
R22415 VDD.n1651 VDD.n1650 19.3944
R22416 VDD.n1654 VDD.n1651 19.3944
R22417 VDD.n1654 VDD.n1191 19.3944
R22418 VDD.n1693 VDD.n1163 19.3944
R22419 VDD.n1693 VDD.n1692 19.3944
R22420 VDD.n1692 VDD.n1691 19.3944
R22421 VDD.n1691 VDD.n1167 19.3944
R22422 VDD.n1687 VDD.n1167 19.3944
R22423 VDD.n1687 VDD.n1686 19.3944
R22424 VDD.n1686 VDD.n1685 19.3944
R22425 VDD.n1685 VDD.n1172 19.3944
R22426 VDD.n1681 VDD.n1172 19.3944
R22427 VDD.n1681 VDD.n1680 19.3944
R22428 VDD.n1680 VDD.n1679 19.3944
R22429 VDD.n1679 VDD.n1177 19.3944
R22430 VDD.n1447 VDD.n1342 19.3944
R22431 VDD.n1447 VDD.n1332 19.3944
R22432 VDD.n1459 VDD.n1332 19.3944
R22433 VDD.n1459 VDD.n1330 19.3944
R22434 VDD.n1463 VDD.n1330 19.3944
R22435 VDD.n1463 VDD.n1320 19.3944
R22436 VDD.n1475 VDD.n1320 19.3944
R22437 VDD.n1475 VDD.n1318 19.3944
R22438 VDD.n1479 VDD.n1318 19.3944
R22439 VDD.n1479 VDD.n1308 19.3944
R22440 VDD.n1491 VDD.n1308 19.3944
R22441 VDD.n1491 VDD.n1306 19.3944
R22442 VDD.n1495 VDD.n1306 19.3944
R22443 VDD.n1495 VDD.n1296 19.3944
R22444 VDD.n1507 VDD.n1296 19.3944
R22445 VDD.n1507 VDD.n1294 19.3944
R22446 VDD.n1511 VDD.n1294 19.3944
R22447 VDD.n1511 VDD.n1284 19.3944
R22448 VDD.n1523 VDD.n1284 19.3944
R22449 VDD.n1523 VDD.n1282 19.3944
R22450 VDD.n1528 VDD.n1282 19.3944
R22451 VDD.n1528 VDD.n1272 19.3944
R22452 VDD.n1540 VDD.n1272 19.3944
R22453 VDD.n1540 VDD.n1266 19.3944
R22454 VDD.n1544 VDD.n1266 19.3944
R22455 VDD.n1544 VDD.n1256 19.3944
R22456 VDD.n1556 VDD.n1256 19.3944
R22457 VDD.n1556 VDD.n1254 19.3944
R22458 VDD.n1560 VDD.n1254 19.3944
R22459 VDD.n1560 VDD.n1244 19.3944
R22460 VDD.n1572 VDD.n1244 19.3944
R22461 VDD.n1572 VDD.n1242 19.3944
R22462 VDD.n1576 VDD.n1242 19.3944
R22463 VDD.n1576 VDD.n1232 19.3944
R22464 VDD.n1588 VDD.n1232 19.3944
R22465 VDD.n1588 VDD.n1230 19.3944
R22466 VDD.n1592 VDD.n1230 19.3944
R22467 VDD.n1592 VDD.n1219 19.3944
R22468 VDD.n1605 VDD.n1219 19.3944
R22469 VDD.n1605 VDD.n1217 19.3944
R22470 VDD.n1609 VDD.n1217 19.3944
R22471 VDD.n1609 VDD.n1206 19.3944
R22472 VDD.n1626 VDD.n1206 19.3944
R22473 VDD.n1626 VDD.n1204 19.3944
R22474 VDD.n1630 VDD.n1204 19.3944
R22475 VDD.n1399 VDD.n1398 18.4247
R22476 VDD.n3472 VDD.n307 18.4247
R22477 VDD.n179 VDD.n99 18.4247
R22478 VDD.n1675 VDD.n1177 18.4247
R22479 VDD.n1422 VDD.n1417 16.0975
R22480 VDD.n3498 VDD.n3497 16.0975
R22481 VDD.n150 VDD.n147 16.0975
R22482 VDD.n1658 VDD.n1163 16.0975
R22483 VDD.n3464 VDD.n3463 14.5893
R22484 VDD.n2085 VDD.n1116 14.5871
R22485 VDD.n1513 VDD.t5 14.4244
R22486 VDD.t3 VDD.n1252 14.4244
R22487 VDD.n3595 VDD.t1 14.4244
R22488 VDD.n3697 VDD.t8 14.4244
R22489 VDD.n2104 VDD.n1102 13.4364
R22490 VDD.n2110 VDD.n1102 13.4364
R22491 VDD.n2110 VDD.n1096 13.4364
R22492 VDD.n2116 VDD.n1096 13.4364
R22493 VDD.n2116 VDD.n1090 13.4364
R22494 VDD.n2122 VDD.n1090 13.4364
R22495 VDD.n2122 VDD.n1084 13.4364
R22496 VDD.n2128 VDD.n1084 13.4364
R22497 VDD.n2134 VDD.n1077 13.4364
R22498 VDD.n2134 VDD.n1080 13.4364
R22499 VDD.n2140 VDD.n1066 13.4364
R22500 VDD.n2146 VDD.n1066 13.4364
R22501 VDD.n2146 VDD.n1060 13.4364
R22502 VDD.n2152 VDD.n1060 13.4364
R22503 VDD.n2152 VDD.n1054 13.4364
R22504 VDD.n2158 VDD.n1054 13.4364
R22505 VDD.n2158 VDD.n1048 13.4364
R22506 VDD.n2164 VDD.n1048 13.4364
R22507 VDD.n2164 VDD.n1042 13.4364
R22508 VDD.n2170 VDD.n1042 13.4364
R22509 VDD.n2170 VDD.n1036 13.4364
R22510 VDD.n2176 VDD.n1036 13.4364
R22511 VDD.n2176 VDD.n1029 13.4364
R22512 VDD.n2182 VDD.n1029 13.4364
R22513 VDD.n2182 VDD.n1032 13.4364
R22514 VDD.n2188 VDD.n1018 13.4364
R22515 VDD.n2194 VDD.n1018 13.4364
R22516 VDD.n2194 VDD.n1012 13.4364
R22517 VDD.n2200 VDD.n1012 13.4364
R22518 VDD.n2200 VDD.n1006 13.4364
R22519 VDD.n2206 VDD.n1006 13.4364
R22520 VDD.n2212 VDD.n1000 13.4364
R22521 VDD.n2212 VDD.n994 13.4364
R22522 VDD.n2218 VDD.n994 13.4364
R22523 VDD.n2218 VDD.n988 13.4364
R22524 VDD.n2224 VDD.n988 13.4364
R22525 VDD.n2224 VDD.n982 13.4364
R22526 VDD.n2230 VDD.n982 13.4364
R22527 VDD.n2230 VDD.n976 13.4364
R22528 VDD.n2236 VDD.n976 13.4364
R22529 VDD.n2236 VDD.n970 13.4364
R22530 VDD.n2242 VDD.n970 13.4364
R22531 VDD.n2242 VDD.n964 13.4364
R22532 VDD.n2248 VDD.n964 13.4364
R22533 VDD.n2248 VDD.n958 13.4364
R22534 VDD.n2254 VDD.n958 13.4364
R22535 VDD.n2254 VDD.n951 13.4364
R22536 VDD.n2260 VDD.n951 13.4364
R22537 VDD.n2260 VDD.n954 13.4364
R22538 VDD.n2266 VDD.n947 13.4364
R22539 VDD.n2272 VDD.n934 13.4364
R22540 VDD.n2278 VDD.n934 13.4364
R22541 VDD.n2278 VDD.n928 13.4364
R22542 VDD.n2284 VDD.n928 13.4364
R22543 VDD.n2284 VDD.n922 13.4364
R22544 VDD.n2290 VDD.n922 13.4364
R22545 VDD.n2290 VDD.n916 13.4364
R22546 VDD.n2296 VDD.n916 13.4364
R22547 VDD.n2296 VDD.n910 13.4364
R22548 VDD.n2302 VDD.n910 13.4364
R22549 VDD.n2302 VDD.n904 13.4364
R22550 VDD.n2308 VDD.n904 13.4364
R22551 VDD.n2308 VDD.n897 13.4364
R22552 VDD.n2314 VDD.n897 13.4364
R22553 VDD.n2314 VDD.n900 13.4364
R22554 VDD.n2320 VDD.n886 13.4364
R22555 VDD.n2326 VDD.n886 13.4364
R22556 VDD.n2332 VDD.n880 13.4364
R22557 VDD.n2332 VDD.n874 13.4364
R22558 VDD.n2338 VDD.n874 13.4364
R22559 VDD.n2338 VDD.n868 13.4364
R22560 VDD.n2344 VDD.n868 13.4364
R22561 VDD.n2344 VDD.n862 13.4364
R22562 VDD.n2350 VDD.n862 13.4364
R22563 VDD.n2350 VDD.n856 13.4364
R22564 VDD.n2356 VDD.n856 13.4364
R22565 VDD.n2356 VDD.n850 13.4364
R22566 VDD.n2362 VDD.n850 13.4364
R22567 VDD.n2362 VDD.n844 13.4364
R22568 VDD.n2368 VDD.n844 13.4364
R22569 VDD.n2368 VDD.n838 13.4364
R22570 VDD.n2374 VDD.n838 13.4364
R22571 VDD.n2380 VDD.n831 13.4364
R22572 VDD.n2380 VDD.n834 13.4364
R22573 VDD.n2386 VDD.n820 13.4364
R22574 VDD.n2392 VDD.n820 13.4364
R22575 VDD.n2392 VDD.n814 13.4364
R22576 VDD.n2398 VDD.n814 13.4364
R22577 VDD.n2398 VDD.n808 13.4364
R22578 VDD.n2404 VDD.n808 13.4364
R22579 VDD.n2404 VDD.n802 13.4364
R22580 VDD.n2410 VDD.n802 13.4364
R22581 VDD.n2410 VDD.n796 13.4364
R22582 VDD.n2416 VDD.n796 13.4364
R22583 VDD.n2416 VDD.n790 13.4364
R22584 VDD.n2422 VDD.n790 13.4364
R22585 VDD.n2422 VDD.n784 13.4364
R22586 VDD.n2428 VDD.n784 13.4364
R22587 VDD.n2428 VDD.n778 13.4364
R22588 VDD.n2434 VDD.n778 13.4364
R22589 VDD.n2434 VDD.n772 13.4364
R22590 VDD.n2440 VDD.n772 13.4364
R22591 VDD.n2446 VDD.n761 13.4364
R22592 VDD.n2452 VDD.n761 13.4364
R22593 VDD.n2452 VDD.n755 13.4364
R22594 VDD.n2458 VDD.n755 13.4364
R22595 VDD.n2458 VDD.n748 13.4364
R22596 VDD.n2502 VDD.n748 13.4364
R22597 VDD.n2502 VDD.n742 13.4364
R22598 VDD.n2508 VDD.n742 13.4364
R22599 VDD.n2508 VDD.n731 13.4364
R22600 VDD.n2550 VDD.n731 13.4364
R22601 VDD.n2550 VDD.n710 13.4364
R22602 VDD.n3012 VDD.n704 13.4364
R22603 VDD.n3018 VDD.n704 13.4364
R22604 VDD.n3018 VDD.n698 13.4364
R22605 VDD.n3024 VDD.n698 13.4364
R22606 VDD.n3024 VDD.n692 13.4364
R22607 VDD.n3030 VDD.n692 13.4364
R22608 VDD.n3030 VDD.n686 13.4364
R22609 VDD.n3036 VDD.n686 13.4364
R22610 VDD.n3036 VDD.n679 13.4364
R22611 VDD.n3042 VDD.n679 13.4364
R22612 VDD.n3042 VDD.n682 13.4364
R22613 VDD.n3054 VDD.n668 13.4364
R22614 VDD.n3054 VDD.n662 13.4364
R22615 VDD.n3060 VDD.n662 13.4364
R22616 VDD.n3060 VDD.n656 13.4364
R22617 VDD.n3066 VDD.n656 13.4364
R22618 VDD.n3066 VDD.n650 13.4364
R22619 VDD.n3072 VDD.n650 13.4364
R22620 VDD.n3072 VDD.n644 13.4364
R22621 VDD.n3078 VDD.n644 13.4364
R22622 VDD.n3078 VDD.n638 13.4364
R22623 VDD.n3084 VDD.n638 13.4364
R22624 VDD.n3084 VDD.n632 13.4364
R22625 VDD.n3090 VDD.n632 13.4364
R22626 VDD.n3090 VDD.n626 13.4364
R22627 VDD.n3096 VDD.n626 13.4364
R22628 VDD.n3096 VDD.n619 13.4364
R22629 VDD.n3102 VDD.n619 13.4364
R22630 VDD.n3102 VDD.n622 13.4364
R22631 VDD.n3108 VDD.n608 13.4364
R22632 VDD.n3114 VDD.n608 13.4364
R22633 VDD.n3120 VDD.n602 13.4364
R22634 VDD.n3120 VDD.n596 13.4364
R22635 VDD.n3126 VDD.n596 13.4364
R22636 VDD.n3126 VDD.n590 13.4364
R22637 VDD.n3132 VDD.n590 13.4364
R22638 VDD.n3132 VDD.n584 13.4364
R22639 VDD.n3138 VDD.n584 13.4364
R22640 VDD.n3138 VDD.n578 13.4364
R22641 VDD.n3144 VDD.n578 13.4364
R22642 VDD.n3144 VDD.n572 13.4364
R22643 VDD.n3150 VDD.n572 13.4364
R22644 VDD.n3150 VDD.n566 13.4364
R22645 VDD.n3156 VDD.n566 13.4364
R22646 VDD.n3156 VDD.n560 13.4364
R22647 VDD.n3162 VDD.n560 13.4364
R22648 VDD.n3168 VDD.n553 13.4364
R22649 VDD.n3168 VDD.n556 13.4364
R22650 VDD.n3174 VDD.n542 13.4364
R22651 VDD.n3180 VDD.n542 13.4364
R22652 VDD.n3180 VDD.n536 13.4364
R22653 VDD.n3186 VDD.n536 13.4364
R22654 VDD.n3186 VDD.n530 13.4364
R22655 VDD.n3192 VDD.n530 13.4364
R22656 VDD.n3192 VDD.n524 13.4364
R22657 VDD.n3198 VDD.n524 13.4364
R22658 VDD.n3198 VDD.n518 13.4364
R22659 VDD.n3204 VDD.n518 13.4364
R22660 VDD.n3204 VDD.n512 13.4364
R22661 VDD.n3210 VDD.n512 13.4364
R22662 VDD.n3210 VDD.n505 13.4364
R22663 VDD.n3216 VDD.n505 13.4364
R22664 VDD.n3216 VDD.n508 13.4364
R22665 VDD.n3222 VDD.n501 13.4364
R22666 VDD.n3228 VDD.n488 13.4364
R22667 VDD.n3234 VDD.n488 13.4364
R22668 VDD.n3234 VDD.n482 13.4364
R22669 VDD.n3240 VDD.n482 13.4364
R22670 VDD.n3240 VDD.n476 13.4364
R22671 VDD.n3246 VDD.n476 13.4364
R22672 VDD.n3246 VDD.n470 13.4364
R22673 VDD.n3252 VDD.n470 13.4364
R22674 VDD.n3252 VDD.n464 13.4364
R22675 VDD.n3258 VDD.n464 13.4364
R22676 VDD.n3258 VDD.n458 13.4364
R22677 VDD.n3264 VDD.n458 13.4364
R22678 VDD.n3264 VDD.n452 13.4364
R22679 VDD.n3270 VDD.n452 13.4364
R22680 VDD.n3270 VDD.n446 13.4364
R22681 VDD.n3276 VDD.n446 13.4364
R22682 VDD.n3276 VDD.n440 13.4364
R22683 VDD.n3282 VDD.n440 13.4364
R22684 VDD.n3288 VDD.n434 13.4364
R22685 VDD.n3288 VDD.n428 13.4364
R22686 VDD.n3294 VDD.n428 13.4364
R22687 VDD.n3294 VDD.n421 13.4364
R22688 VDD.n3300 VDD.n421 13.4364
R22689 VDD.n3300 VDD.n424 13.4364
R22690 VDD.n3306 VDD.n410 13.4364
R22691 VDD.n3312 VDD.n410 13.4364
R22692 VDD.n3312 VDD.n404 13.4364
R22693 VDD.n3318 VDD.n404 13.4364
R22694 VDD.n3318 VDD.n398 13.4364
R22695 VDD.n3324 VDD.n398 13.4364
R22696 VDD.n3324 VDD.n392 13.4364
R22697 VDD.n3330 VDD.n392 13.4364
R22698 VDD.n3330 VDD.n386 13.4364
R22699 VDD.n3336 VDD.n386 13.4364
R22700 VDD.n3336 VDD.n380 13.4364
R22701 VDD.n3342 VDD.n380 13.4364
R22702 VDD.n3342 VDD.n373 13.4364
R22703 VDD.n3348 VDD.n373 13.4364
R22704 VDD.n3348 VDD.n376 13.4364
R22705 VDD.n3354 VDD.n362 13.4364
R22706 VDD.n3360 VDD.n362 13.4364
R22707 VDD.n3366 VDD.n356 13.4364
R22708 VDD.n3366 VDD.n349 13.4364
R22709 VDD.n3397 VDD.n349 13.4364
R22710 VDD.n3397 VDD.n343 13.4364
R22711 VDD.n3403 VDD.n343 13.4364
R22712 VDD.n3403 VDD.n321 13.4364
R22713 VDD.n3443 VDD.n321 13.4364
R22714 VDD.n3443 VDD.n323 13.4364
R22715 VDD.t37 VDD.n1322 12.8437
R22716 VDD.n1603 VDD.t29 12.8437
R22717 VDD.n2140 VDD.t25 12.8437
R22718 VDD.n2266 VDD.t73 12.8437
R22719 VDD.n900 VDD.t95 12.8437
R22720 VDD.n1896 VDD.t17 12.8437
R22721 VDD.n3048 VDD.t33 12.8437
R22722 VDD.n3174 VDD.t78 12.8437
R22723 VDD.n501 VDD.t91 12.8437
R22724 VDD.n376 VDD.t21 12.8437
R22725 VDD.t50 VDD.n238 12.8437
R22726 VDD.t13 VDD.n62 12.8437
R22727 VDD.t83 VDD.n1000 11.6582
R22728 VDD.n2374 VDD.t104 11.6582
R22729 VDD.t92 VDD.n602 11.6582
R22730 VDD.n3282 VDD.t90 11.6582
R22731 VDD.n3523 VDD.n260 10.8277
R22732 VDD.n1697 VDD.n1696 10.8274
R22733 VDD.n2780 VDD.n2779 10.6151
R22734 VDD.n2779 VDD.n2778 10.6151
R22735 VDD.n2778 VDD.n2777 10.6151
R22736 VDD.n2777 VDD.n2775 10.6151
R22737 VDD.n2775 VDD.n2774 10.6151
R22738 VDD.n2774 VDD.n2772 10.6151
R22739 VDD.n2772 VDD.n2771 10.6151
R22740 VDD.n2771 VDD.n2769 10.6151
R22741 VDD.n2769 VDD.n2768 10.6151
R22742 VDD.n2768 VDD.n2766 10.6151
R22743 VDD.n2766 VDD.n2765 10.6151
R22744 VDD.n2765 VDD.n2763 10.6151
R22745 VDD.n2763 VDD.n2762 10.6151
R22746 VDD.n2762 VDD.n2760 10.6151
R22747 VDD.n2760 VDD.n2759 10.6151
R22748 VDD.n2759 VDD.n2757 10.6151
R22749 VDD.n2757 VDD.n2756 10.6151
R22750 VDD.n2756 VDD.n2754 10.6151
R22751 VDD.n2754 VDD.n2753 10.6151
R22752 VDD.n2753 VDD.n2751 10.6151
R22753 VDD.n2751 VDD.n2750 10.6151
R22754 VDD.n2750 VDD.n2748 10.6151
R22755 VDD.n2748 VDD.n2747 10.6151
R22756 VDD.n2747 VDD.n2745 10.6151
R22757 VDD.n2745 VDD.n2744 10.6151
R22758 VDD.n2744 VDD.n2742 10.6151
R22759 VDD.n2742 VDD.n2741 10.6151
R22760 VDD.n2741 VDD.n2739 10.6151
R22761 VDD.n2739 VDD.n2738 10.6151
R22762 VDD.n2738 VDD.n2736 10.6151
R22763 VDD.n2736 VDD.n2735 10.6151
R22764 VDD.n2735 VDD.n2733 10.6151
R22765 VDD.n2733 VDD.n2732 10.6151
R22766 VDD.n2732 VDD.n2730 10.6151
R22767 VDD.n2730 VDD.n2729 10.6151
R22768 VDD.n2729 VDD.n2727 10.6151
R22769 VDD.n2727 VDD.n2726 10.6151
R22770 VDD.n2726 VDD.n2724 10.6151
R22771 VDD.n2724 VDD.n2723 10.6151
R22772 VDD.n2723 VDD.n2721 10.6151
R22773 VDD.n2721 VDD.n2720 10.6151
R22774 VDD.n2720 VDD.n2718 10.6151
R22775 VDD.n2718 VDD.n2717 10.6151
R22776 VDD.n2717 VDD.n2715 10.6151
R22777 VDD.n2715 VDD.n2714 10.6151
R22778 VDD.n2714 VDD.n2712 10.6151
R22779 VDD.n2712 VDD.n2711 10.6151
R22780 VDD.n2711 VDD.n2709 10.6151
R22781 VDD.n2709 VDD.n2708 10.6151
R22782 VDD.n2708 VDD.n2706 10.6151
R22783 VDD.n2706 VDD.n2705 10.6151
R22784 VDD.n2705 VDD.n2703 10.6151
R22785 VDD.n2703 VDD.n2702 10.6151
R22786 VDD.n2702 VDD.n2700 10.6151
R22787 VDD.n2700 VDD.n2699 10.6151
R22788 VDD.n2699 VDD.n2697 10.6151
R22789 VDD.n2697 VDD.n2696 10.6151
R22790 VDD.n2696 VDD.n2694 10.6151
R22791 VDD.n2694 VDD.n2693 10.6151
R22792 VDD.n2693 VDD.n2691 10.6151
R22793 VDD.n2691 VDD.n2690 10.6151
R22794 VDD.n2690 VDD.n2688 10.6151
R22795 VDD.n2688 VDD.n2687 10.6151
R22796 VDD.n2687 VDD.n2685 10.6151
R22797 VDD.n2685 VDD.n2684 10.6151
R22798 VDD.n2684 VDD.n2682 10.6151
R22799 VDD.n2682 VDD.n2681 10.6151
R22800 VDD.n2681 VDD.n2679 10.6151
R22801 VDD.n2679 VDD.n2678 10.6151
R22802 VDD.n2678 VDD.n2676 10.6151
R22803 VDD.n2676 VDD.n2675 10.6151
R22804 VDD.n2675 VDD.n2673 10.6151
R22805 VDD.n2673 VDD.n2672 10.6151
R22806 VDD.n2672 VDD.n2670 10.6151
R22807 VDD.n2670 VDD.n2669 10.6151
R22808 VDD.n2669 VDD.n2667 10.6151
R22809 VDD.n2667 VDD.n2666 10.6151
R22810 VDD.n2666 VDD.n2664 10.6151
R22811 VDD.n2664 VDD.n2663 10.6151
R22812 VDD.n2663 VDD.n2661 10.6151
R22813 VDD.n2661 VDD.n2660 10.6151
R22814 VDD.n2660 VDD.n2658 10.6151
R22815 VDD.n2658 VDD.n2657 10.6151
R22816 VDD.n2657 VDD.n2655 10.6151
R22817 VDD.n2655 VDD.n2654 10.6151
R22818 VDD.n2654 VDD.n2652 10.6151
R22819 VDD.n2652 VDD.n2651 10.6151
R22820 VDD.n2651 VDD.n2649 10.6151
R22821 VDD.n2649 VDD.n2648 10.6151
R22822 VDD.n2648 VDD.n2646 10.6151
R22823 VDD.n2646 VDD.n2645 10.6151
R22824 VDD.n2645 VDD.n2643 10.6151
R22825 VDD.n2643 VDD.n2642 10.6151
R22826 VDD.n2642 VDD.n2640 10.6151
R22827 VDD.n2640 VDD.n2639 10.6151
R22828 VDD.n2639 VDD.n2637 10.6151
R22829 VDD.n2637 VDD.n2636 10.6151
R22830 VDD.n2636 VDD.n2634 10.6151
R22831 VDD.n2634 VDD.n2633 10.6151
R22832 VDD.n2633 VDD.n2631 10.6151
R22833 VDD.n2631 VDD.n2630 10.6151
R22834 VDD.n2630 VDD.n2628 10.6151
R22835 VDD.n2628 VDD.n2627 10.6151
R22836 VDD.n2627 VDD.n2625 10.6151
R22837 VDD.n2625 VDD.n2624 10.6151
R22838 VDD.n2624 VDD.n2622 10.6151
R22839 VDD.n2622 VDD.n2621 10.6151
R22840 VDD.n2621 VDD.n2619 10.6151
R22841 VDD.n2619 VDD.n2618 10.6151
R22842 VDD.n2618 VDD.n2616 10.6151
R22843 VDD.n2616 VDD.n2615 10.6151
R22844 VDD.n2615 VDD.n2613 10.6151
R22845 VDD.n2613 VDD.n2612 10.6151
R22846 VDD.n2612 VDD.n2610 10.6151
R22847 VDD.n2610 VDD.n2609 10.6151
R22848 VDD.n2609 VDD.n2607 10.6151
R22849 VDD.n2607 VDD.n2606 10.6151
R22850 VDD.n2606 VDD.n2604 10.6151
R22851 VDD.n2604 VDD.n2603 10.6151
R22852 VDD.n2603 VDD.n2601 10.6151
R22853 VDD.n2601 VDD.n2600 10.6151
R22854 VDD.n2600 VDD.n341 10.6151
R22855 VDD.n3406 VDD.n341 10.6151
R22856 VDD.n3407 VDD.n3406 10.6151
R22857 VDD.n3408 VDD.n3407 10.6151
R22858 VDD.n2570 VDD.n708 10.6151
R22859 VDD.n2571 VDD.n2570 10.6151
R22860 VDD.n2572 VDD.n2571 10.6151
R22861 VDD.n2572 VDD.n2566 10.6151
R22862 VDD.n2578 VDD.n2566 10.6151
R22863 VDD.n2579 VDD.n2578 10.6151
R22864 VDD.n2580 VDD.n2579 10.6151
R22865 VDD.n2580 VDD.n2564 10.6151
R22866 VDD.n2586 VDD.n2564 10.6151
R22867 VDD.n2587 VDD.n2586 10.6151
R22868 VDD.n2591 VDD.n2587 10.6151
R22869 VDD.n2562 VDD.n2561 10.6151
R22870 VDD.n2598 VDD.n2561 10.6151
R22871 VDD.n2599 VDD.n2598 10.6151
R22872 VDD.n3015 VDD.n3014 10.6151
R22873 VDD.n3016 VDD.n3015 10.6151
R22874 VDD.n3016 VDD.n696 10.6151
R22875 VDD.n3026 VDD.n696 10.6151
R22876 VDD.n3027 VDD.n3026 10.6151
R22877 VDD.n3028 VDD.n3027 10.6151
R22878 VDD.n3028 VDD.n684 10.6151
R22879 VDD.n3038 VDD.n684 10.6151
R22880 VDD.n3039 VDD.n3038 10.6151
R22881 VDD.n3040 VDD.n3039 10.6151
R22882 VDD.n3040 VDD.n672 10.6151
R22883 VDD.n3050 VDD.n672 10.6151
R22884 VDD.n3051 VDD.n3050 10.6151
R22885 VDD.n3052 VDD.n3051 10.6151
R22886 VDD.n3052 VDD.n660 10.6151
R22887 VDD.n3062 VDD.n660 10.6151
R22888 VDD.n3063 VDD.n3062 10.6151
R22889 VDD.n3064 VDD.n3063 10.6151
R22890 VDD.n3064 VDD.n648 10.6151
R22891 VDD.n3074 VDD.n648 10.6151
R22892 VDD.n3075 VDD.n3074 10.6151
R22893 VDD.n3076 VDD.n3075 10.6151
R22894 VDD.n3076 VDD.n636 10.6151
R22895 VDD.n3086 VDD.n636 10.6151
R22896 VDD.n3087 VDD.n3086 10.6151
R22897 VDD.n3088 VDD.n3087 10.6151
R22898 VDD.n3088 VDD.n624 10.6151
R22899 VDD.n3098 VDD.n624 10.6151
R22900 VDD.n3099 VDD.n3098 10.6151
R22901 VDD.n3100 VDD.n3099 10.6151
R22902 VDD.n3100 VDD.n612 10.6151
R22903 VDD.n3110 VDD.n612 10.6151
R22904 VDD.n3111 VDD.n3110 10.6151
R22905 VDD.n3112 VDD.n3111 10.6151
R22906 VDD.n3112 VDD.n600 10.6151
R22907 VDD.n3122 VDD.n600 10.6151
R22908 VDD.n3123 VDD.n3122 10.6151
R22909 VDD.n3124 VDD.n3123 10.6151
R22910 VDD.n3124 VDD.n588 10.6151
R22911 VDD.n3134 VDD.n588 10.6151
R22912 VDD.n3135 VDD.n3134 10.6151
R22913 VDD.n3136 VDD.n3135 10.6151
R22914 VDD.n3136 VDD.n576 10.6151
R22915 VDD.n3146 VDD.n576 10.6151
R22916 VDD.n3147 VDD.n3146 10.6151
R22917 VDD.n3148 VDD.n3147 10.6151
R22918 VDD.n3148 VDD.n564 10.6151
R22919 VDD.n3158 VDD.n564 10.6151
R22920 VDD.n3159 VDD.n3158 10.6151
R22921 VDD.n3160 VDD.n3159 10.6151
R22922 VDD.n3160 VDD.n551 10.6151
R22923 VDD.n3170 VDD.n551 10.6151
R22924 VDD.n3171 VDD.n3170 10.6151
R22925 VDD.n3172 VDD.n3171 10.6151
R22926 VDD.n3172 VDD.n540 10.6151
R22927 VDD.n3182 VDD.n540 10.6151
R22928 VDD.n3183 VDD.n3182 10.6151
R22929 VDD.n3184 VDD.n3183 10.6151
R22930 VDD.n3184 VDD.n528 10.6151
R22931 VDD.n3194 VDD.n528 10.6151
R22932 VDD.n3195 VDD.n3194 10.6151
R22933 VDD.n3196 VDD.n3195 10.6151
R22934 VDD.n3196 VDD.n516 10.6151
R22935 VDD.n3206 VDD.n516 10.6151
R22936 VDD.n3207 VDD.n3206 10.6151
R22937 VDD.n3208 VDD.n3207 10.6151
R22938 VDD.n3208 VDD.n503 10.6151
R22939 VDD.n3218 VDD.n503 10.6151
R22940 VDD.n3219 VDD.n3218 10.6151
R22941 VDD.n3220 VDD.n3219 10.6151
R22942 VDD.n3220 VDD.n492 10.6151
R22943 VDD.n3230 VDD.n492 10.6151
R22944 VDD.n3231 VDD.n3230 10.6151
R22945 VDD.n3232 VDD.n3231 10.6151
R22946 VDD.n3232 VDD.n480 10.6151
R22947 VDD.n3242 VDD.n480 10.6151
R22948 VDD.n3243 VDD.n3242 10.6151
R22949 VDD.n3244 VDD.n3243 10.6151
R22950 VDD.n3244 VDD.n468 10.6151
R22951 VDD.n3254 VDD.n468 10.6151
R22952 VDD.n3255 VDD.n3254 10.6151
R22953 VDD.n3256 VDD.n3255 10.6151
R22954 VDD.n3256 VDD.n456 10.6151
R22955 VDD.n3266 VDD.n456 10.6151
R22956 VDD.n3267 VDD.n3266 10.6151
R22957 VDD.n3268 VDD.n3267 10.6151
R22958 VDD.n3268 VDD.n444 10.6151
R22959 VDD.n3278 VDD.n444 10.6151
R22960 VDD.n3279 VDD.n3278 10.6151
R22961 VDD.n3280 VDD.n3279 10.6151
R22962 VDD.n3280 VDD.n432 10.6151
R22963 VDD.n3290 VDD.n432 10.6151
R22964 VDD.n3291 VDD.n3290 10.6151
R22965 VDD.n3292 VDD.n3291 10.6151
R22966 VDD.n3292 VDD.n419 10.6151
R22967 VDD.n3302 VDD.n419 10.6151
R22968 VDD.n3303 VDD.n3302 10.6151
R22969 VDD.n3304 VDD.n3303 10.6151
R22970 VDD.n3304 VDD.n408 10.6151
R22971 VDD.n3314 VDD.n408 10.6151
R22972 VDD.n3315 VDD.n3314 10.6151
R22973 VDD.n3316 VDD.n3315 10.6151
R22974 VDD.n3316 VDD.n396 10.6151
R22975 VDD.n3326 VDD.n396 10.6151
R22976 VDD.n3327 VDD.n3326 10.6151
R22977 VDD.n3328 VDD.n3327 10.6151
R22978 VDD.n3328 VDD.n384 10.6151
R22979 VDD.n3338 VDD.n384 10.6151
R22980 VDD.n3339 VDD.n3338 10.6151
R22981 VDD.n3340 VDD.n3339 10.6151
R22982 VDD.n3340 VDD.n371 10.6151
R22983 VDD.n3350 VDD.n371 10.6151
R22984 VDD.n3351 VDD.n3350 10.6151
R22985 VDD.n3352 VDD.n3351 10.6151
R22986 VDD.n3352 VDD.n360 10.6151
R22987 VDD.n3362 VDD.n360 10.6151
R22988 VDD.n3363 VDD.n3362 10.6151
R22989 VDD.n3364 VDD.n3363 10.6151
R22990 VDD.n3364 VDD.n347 10.6151
R22991 VDD.n3399 VDD.n347 10.6151
R22992 VDD.n3400 VDD.n3399 10.6151
R22993 VDD.n3401 VDD.n3400 10.6151
R22994 VDD.n3401 VDD.n327 10.6151
R22995 VDD.n3441 VDD.n327 10.6151
R22996 VDD.n3441 VDD.n3440 10.6151
R22997 VDD.n3439 VDD.n328 10.6151
R22998 VDD.n329 VDD.n328 10.6151
R22999 VDD.n3432 VDD.n329 10.6151
R23000 VDD.n3432 VDD.n3431 10.6151
R23001 VDD.n3431 VDD.n3430 10.6151
R23002 VDD.n3430 VDD.n331 10.6151
R23003 VDD.n3425 VDD.n331 10.6151
R23004 VDD.n3421 VDD.n333 10.6151
R23005 VDD.n3421 VDD.n3420 10.6151
R23006 VDD.n3420 VDD.n3419 10.6151
R23007 VDD.n3414 VDD.n339 10.6151
R23008 VDD.n3414 VDD.n3413 10.6151
R23009 VDD.n3413 VDD.n3412 10.6151
R23010 VDD.n3384 VDD.n3370 10.6151
R23011 VDD.n3384 VDD.n3383 10.6151
R23012 VDD.n3383 VDD.n3382 10.6151
R23013 VDD.n3382 VDD.n3372 10.6151
R23014 VDD.n3377 VDD.n3372 10.6151
R23015 VDD.n3377 VDD.n3376 10.6151
R23016 VDD.n3376 VDD.n308 10.6151
R23017 VDD.n3462 VDD.n309 10.6151
R23018 VDD.n312 VDD.n309 10.6151
R23019 VDD.n3455 VDD.n312 10.6151
R23020 VDD.n3453 VDD.n3452 10.6151
R23021 VDD.n3452 VDD.n316 10.6151
R23022 VDD.n3447 VDD.n316 10.6151
R23023 VDD.n2976 VDD.n2975 10.6151
R23024 VDD.n2975 VDD.n2973 10.6151
R23025 VDD.n2973 VDD.n2972 10.6151
R23026 VDD.n2972 VDD.n2970 10.6151
R23027 VDD.n2970 VDD.n2969 10.6151
R23028 VDD.n2969 VDD.n2967 10.6151
R23029 VDD.n2967 VDD.n2966 10.6151
R23030 VDD.n2966 VDD.n2964 10.6151
R23031 VDD.n2964 VDD.n2963 10.6151
R23032 VDD.n2963 VDD.n2961 10.6151
R23033 VDD.n2961 VDD.n2960 10.6151
R23034 VDD.n2960 VDD.n2958 10.6151
R23035 VDD.n2958 VDD.n2957 10.6151
R23036 VDD.n2957 VDD.n2955 10.6151
R23037 VDD.n2955 VDD.n2954 10.6151
R23038 VDD.n2954 VDD.n2952 10.6151
R23039 VDD.n2952 VDD.n2951 10.6151
R23040 VDD.n2951 VDD.n2949 10.6151
R23041 VDD.n2949 VDD.n2948 10.6151
R23042 VDD.n2948 VDD.n2946 10.6151
R23043 VDD.n2946 VDD.n2945 10.6151
R23044 VDD.n2945 VDD.n2943 10.6151
R23045 VDD.n2943 VDD.n2942 10.6151
R23046 VDD.n2942 VDD.n2940 10.6151
R23047 VDD.n2940 VDD.n2939 10.6151
R23048 VDD.n2939 VDD.n2937 10.6151
R23049 VDD.n2937 VDD.n2936 10.6151
R23050 VDD.n2936 VDD.n2934 10.6151
R23051 VDD.n2934 VDD.n2933 10.6151
R23052 VDD.n2933 VDD.n2931 10.6151
R23053 VDD.n2931 VDD.n2930 10.6151
R23054 VDD.n2930 VDD.n2928 10.6151
R23055 VDD.n2928 VDD.n2927 10.6151
R23056 VDD.n2927 VDD.n2925 10.6151
R23057 VDD.n2925 VDD.n2924 10.6151
R23058 VDD.n2924 VDD.n2922 10.6151
R23059 VDD.n2922 VDD.n2921 10.6151
R23060 VDD.n2921 VDD.n2919 10.6151
R23061 VDD.n2919 VDD.n2918 10.6151
R23062 VDD.n2918 VDD.n2916 10.6151
R23063 VDD.n2916 VDD.n2915 10.6151
R23064 VDD.n2915 VDD.n2913 10.6151
R23065 VDD.n2913 VDD.n2912 10.6151
R23066 VDD.n2912 VDD.n2910 10.6151
R23067 VDD.n2910 VDD.n2909 10.6151
R23068 VDD.n2909 VDD.n2907 10.6151
R23069 VDD.n2907 VDD.n2906 10.6151
R23070 VDD.n2906 VDD.n2904 10.6151
R23071 VDD.n2904 VDD.n2903 10.6151
R23072 VDD.n2903 VDD.n2901 10.6151
R23073 VDD.n2901 VDD.n2900 10.6151
R23074 VDD.n2900 VDD.n2898 10.6151
R23075 VDD.n2898 VDD.n2897 10.6151
R23076 VDD.n2897 VDD.n2895 10.6151
R23077 VDD.n2895 VDD.n2894 10.6151
R23078 VDD.n2894 VDD.n2892 10.6151
R23079 VDD.n2892 VDD.n2891 10.6151
R23080 VDD.n2891 VDD.n2889 10.6151
R23081 VDD.n2889 VDD.n2888 10.6151
R23082 VDD.n2888 VDD.n2886 10.6151
R23083 VDD.n2886 VDD.n2885 10.6151
R23084 VDD.n2885 VDD.n2883 10.6151
R23085 VDD.n2883 VDD.n2882 10.6151
R23086 VDD.n2882 VDD.n2880 10.6151
R23087 VDD.n2880 VDD.n2879 10.6151
R23088 VDD.n2879 VDD.n2877 10.6151
R23089 VDD.n2877 VDD.n2876 10.6151
R23090 VDD.n2876 VDD.n2874 10.6151
R23091 VDD.n2874 VDD.n2873 10.6151
R23092 VDD.n2873 VDD.n2871 10.6151
R23093 VDD.n2871 VDD.n2870 10.6151
R23094 VDD.n2870 VDD.n2868 10.6151
R23095 VDD.n2868 VDD.n2867 10.6151
R23096 VDD.n2867 VDD.n2865 10.6151
R23097 VDD.n2865 VDD.n2864 10.6151
R23098 VDD.n2864 VDD.n2862 10.6151
R23099 VDD.n2862 VDD.n2861 10.6151
R23100 VDD.n2861 VDD.n2859 10.6151
R23101 VDD.n2859 VDD.n2858 10.6151
R23102 VDD.n2858 VDD.n2856 10.6151
R23103 VDD.n2856 VDD.n2855 10.6151
R23104 VDD.n2855 VDD.n2853 10.6151
R23105 VDD.n2853 VDD.n2852 10.6151
R23106 VDD.n2852 VDD.n2850 10.6151
R23107 VDD.n2850 VDD.n2849 10.6151
R23108 VDD.n2849 VDD.n2847 10.6151
R23109 VDD.n2847 VDD.n2846 10.6151
R23110 VDD.n2846 VDD.n2844 10.6151
R23111 VDD.n2844 VDD.n2843 10.6151
R23112 VDD.n2843 VDD.n2841 10.6151
R23113 VDD.n2841 VDD.n2840 10.6151
R23114 VDD.n2840 VDD.n2838 10.6151
R23115 VDD.n2838 VDD.n2837 10.6151
R23116 VDD.n2837 VDD.n2835 10.6151
R23117 VDD.n2835 VDD.n2834 10.6151
R23118 VDD.n2834 VDD.n2832 10.6151
R23119 VDD.n2832 VDD.n2831 10.6151
R23120 VDD.n2831 VDD.n2829 10.6151
R23121 VDD.n2829 VDD.n2828 10.6151
R23122 VDD.n2828 VDD.n2826 10.6151
R23123 VDD.n2826 VDD.n2825 10.6151
R23124 VDD.n2825 VDD.n2823 10.6151
R23125 VDD.n2823 VDD.n2822 10.6151
R23126 VDD.n2822 VDD.n2820 10.6151
R23127 VDD.n2820 VDD.n2819 10.6151
R23128 VDD.n2819 VDD.n2817 10.6151
R23129 VDD.n2817 VDD.n2816 10.6151
R23130 VDD.n2816 VDD.n2814 10.6151
R23131 VDD.n2814 VDD.n2813 10.6151
R23132 VDD.n2813 VDD.n2811 10.6151
R23133 VDD.n2811 VDD.n2810 10.6151
R23134 VDD.n2810 VDD.n2808 10.6151
R23135 VDD.n2808 VDD.n2807 10.6151
R23136 VDD.n2807 VDD.n2805 10.6151
R23137 VDD.n2805 VDD.n2804 10.6151
R23138 VDD.n2804 VDD.n2802 10.6151
R23139 VDD.n2802 VDD.n2801 10.6151
R23140 VDD.n2801 VDD.n2799 10.6151
R23141 VDD.n2799 VDD.n2798 10.6151
R23142 VDD.n2798 VDD.n2796 10.6151
R23143 VDD.n2796 VDD.n2795 10.6151
R23144 VDD.n2795 VDD.n2793 10.6151
R23145 VDD.n2793 VDD.n319 10.6151
R23146 VDD.n3445 VDD.n319 10.6151
R23147 VDD.n3446 VDD.n3445 10.6151
R23148 VDD.n3009 VDD.n3008 10.6151
R23149 VDD.n3008 VDD.n2784 10.6151
R23150 VDD.n3002 VDD.n2784 10.6151
R23151 VDD.n3002 VDD.n3001 10.6151
R23152 VDD.n3001 VDD.n3000 10.6151
R23153 VDD.n3000 VDD.n2786 10.6151
R23154 VDD.n2994 VDD.n2786 10.6151
R23155 VDD.n2994 VDD.n2993 10.6151
R23156 VDD.n2993 VDD.n2992 10.6151
R23157 VDD.n2992 VDD.n2788 10.6151
R23158 VDD.n2986 VDD.n2788 10.6151
R23159 VDD.n2984 VDD.n2983 10.6151
R23160 VDD.n2983 VDD.n2792 10.6151
R23161 VDD.n2977 VDD.n2792 10.6151
R23162 VDD.n3010 VDD.n702 10.6151
R23163 VDD.n3020 VDD.n702 10.6151
R23164 VDD.n3021 VDD.n3020 10.6151
R23165 VDD.n3022 VDD.n3021 10.6151
R23166 VDD.n3022 VDD.n690 10.6151
R23167 VDD.n3032 VDD.n690 10.6151
R23168 VDD.n3033 VDD.n3032 10.6151
R23169 VDD.n3034 VDD.n3033 10.6151
R23170 VDD.n3034 VDD.n677 10.6151
R23171 VDD.n3044 VDD.n677 10.6151
R23172 VDD.n3045 VDD.n3044 10.6151
R23173 VDD.n3046 VDD.n3045 10.6151
R23174 VDD.n3046 VDD.n666 10.6151
R23175 VDD.n3056 VDD.n666 10.6151
R23176 VDD.n3057 VDD.n3056 10.6151
R23177 VDD.n3058 VDD.n3057 10.6151
R23178 VDD.n3058 VDD.n654 10.6151
R23179 VDD.n3068 VDD.n654 10.6151
R23180 VDD.n3069 VDD.n3068 10.6151
R23181 VDD.n3070 VDD.n3069 10.6151
R23182 VDD.n3070 VDD.n642 10.6151
R23183 VDD.n3080 VDD.n642 10.6151
R23184 VDD.n3081 VDD.n3080 10.6151
R23185 VDD.n3082 VDD.n3081 10.6151
R23186 VDD.n3082 VDD.n630 10.6151
R23187 VDD.n3092 VDD.n630 10.6151
R23188 VDD.n3093 VDD.n3092 10.6151
R23189 VDD.n3094 VDD.n3093 10.6151
R23190 VDD.n3094 VDD.n617 10.6151
R23191 VDD.n3104 VDD.n617 10.6151
R23192 VDD.n3105 VDD.n3104 10.6151
R23193 VDD.n3106 VDD.n3105 10.6151
R23194 VDD.n3106 VDD.n606 10.6151
R23195 VDD.n3116 VDD.n606 10.6151
R23196 VDD.n3117 VDD.n3116 10.6151
R23197 VDD.n3118 VDD.n3117 10.6151
R23198 VDD.n3118 VDD.n594 10.6151
R23199 VDD.n3128 VDD.n594 10.6151
R23200 VDD.n3129 VDD.n3128 10.6151
R23201 VDD.n3130 VDD.n3129 10.6151
R23202 VDD.n3130 VDD.n582 10.6151
R23203 VDD.n3140 VDD.n582 10.6151
R23204 VDD.n3141 VDD.n3140 10.6151
R23205 VDD.n3142 VDD.n3141 10.6151
R23206 VDD.n3142 VDD.n570 10.6151
R23207 VDD.n3152 VDD.n570 10.6151
R23208 VDD.n3153 VDD.n3152 10.6151
R23209 VDD.n3154 VDD.n3153 10.6151
R23210 VDD.n3154 VDD.n558 10.6151
R23211 VDD.n3164 VDD.n558 10.6151
R23212 VDD.n3165 VDD.n3164 10.6151
R23213 VDD.n3166 VDD.n3165 10.6151
R23214 VDD.n3166 VDD.n546 10.6151
R23215 VDD.n3176 VDD.n546 10.6151
R23216 VDD.n3177 VDD.n3176 10.6151
R23217 VDD.n3178 VDD.n3177 10.6151
R23218 VDD.n3178 VDD.n534 10.6151
R23219 VDD.n3188 VDD.n534 10.6151
R23220 VDD.n3189 VDD.n3188 10.6151
R23221 VDD.n3190 VDD.n3189 10.6151
R23222 VDD.n3190 VDD.n522 10.6151
R23223 VDD.n3200 VDD.n522 10.6151
R23224 VDD.n3201 VDD.n3200 10.6151
R23225 VDD.n3202 VDD.n3201 10.6151
R23226 VDD.n3202 VDD.n510 10.6151
R23227 VDD.n3212 VDD.n510 10.6151
R23228 VDD.n3213 VDD.n3212 10.6151
R23229 VDD.n3214 VDD.n3213 10.6151
R23230 VDD.n3214 VDD.n497 10.6151
R23231 VDD.n3224 VDD.n497 10.6151
R23232 VDD.n3225 VDD.n3224 10.6151
R23233 VDD.n3226 VDD.n3225 10.6151
R23234 VDD.n3226 VDD.n486 10.6151
R23235 VDD.n3236 VDD.n486 10.6151
R23236 VDD.n3237 VDD.n3236 10.6151
R23237 VDD.n3238 VDD.n3237 10.6151
R23238 VDD.n3238 VDD.n474 10.6151
R23239 VDD.n3248 VDD.n474 10.6151
R23240 VDD.n3249 VDD.n3248 10.6151
R23241 VDD.n3250 VDD.n3249 10.6151
R23242 VDD.n3250 VDD.n462 10.6151
R23243 VDD.n3260 VDD.n462 10.6151
R23244 VDD.n3261 VDD.n3260 10.6151
R23245 VDD.n3262 VDD.n3261 10.6151
R23246 VDD.n3262 VDD.n450 10.6151
R23247 VDD.n3272 VDD.n450 10.6151
R23248 VDD.n3273 VDD.n3272 10.6151
R23249 VDD.n3274 VDD.n3273 10.6151
R23250 VDD.n3274 VDD.n438 10.6151
R23251 VDD.n3284 VDD.n438 10.6151
R23252 VDD.n3285 VDD.n3284 10.6151
R23253 VDD.n3286 VDD.n3285 10.6151
R23254 VDD.n3286 VDD.n426 10.6151
R23255 VDD.n3296 VDD.n426 10.6151
R23256 VDD.n3297 VDD.n3296 10.6151
R23257 VDD.n3298 VDD.n3297 10.6151
R23258 VDD.n3298 VDD.n414 10.6151
R23259 VDD.n3308 VDD.n414 10.6151
R23260 VDD.n3309 VDD.n3308 10.6151
R23261 VDD.n3310 VDD.n3309 10.6151
R23262 VDD.n3310 VDD.n402 10.6151
R23263 VDD.n3320 VDD.n402 10.6151
R23264 VDD.n3321 VDD.n3320 10.6151
R23265 VDD.n3322 VDD.n3321 10.6151
R23266 VDD.n3322 VDD.n390 10.6151
R23267 VDD.n3332 VDD.n390 10.6151
R23268 VDD.n3333 VDD.n3332 10.6151
R23269 VDD.n3334 VDD.n3333 10.6151
R23270 VDD.n3334 VDD.n378 10.6151
R23271 VDD.n3344 VDD.n378 10.6151
R23272 VDD.n3345 VDD.n3344 10.6151
R23273 VDD.n3346 VDD.n3345 10.6151
R23274 VDD.n3346 VDD.n366 10.6151
R23275 VDD.n3356 VDD.n366 10.6151
R23276 VDD.n3357 VDD.n3356 10.6151
R23277 VDD.n3358 VDD.n3357 10.6151
R23278 VDD.n3358 VDD.n354 10.6151
R23279 VDD.n3368 VDD.n354 10.6151
R23280 VDD.n3369 VDD.n3368 10.6151
R23281 VDD.n3395 VDD.n3369 10.6151
R23282 VDD.n3395 VDD.n3394 10.6151
R23283 VDD.n3394 VDD.n3393 10.6151
R23284 VDD.n3393 VDD.n3392 10.6151
R23285 VDD.n3392 VDD.n3390 10.6151
R23286 VDD.n3390 VDD.n3389 10.6151
R23287 VDD.n2107 VDD.n2106 10.6151
R23288 VDD.n2108 VDD.n2107 10.6151
R23289 VDD.n2108 VDD.n1094 10.6151
R23290 VDD.n2118 VDD.n1094 10.6151
R23291 VDD.n2119 VDD.n2118 10.6151
R23292 VDD.n2120 VDD.n2119 10.6151
R23293 VDD.n2120 VDD.n1082 10.6151
R23294 VDD.n2130 VDD.n1082 10.6151
R23295 VDD.n2131 VDD.n2130 10.6151
R23296 VDD.n2132 VDD.n2131 10.6151
R23297 VDD.n2132 VDD.n1070 10.6151
R23298 VDD.n2142 VDD.n1070 10.6151
R23299 VDD.n2143 VDD.n2142 10.6151
R23300 VDD.n2144 VDD.n2143 10.6151
R23301 VDD.n2144 VDD.n1058 10.6151
R23302 VDD.n2154 VDD.n1058 10.6151
R23303 VDD.n2155 VDD.n2154 10.6151
R23304 VDD.n2156 VDD.n2155 10.6151
R23305 VDD.n2156 VDD.n1046 10.6151
R23306 VDD.n2166 VDD.n1046 10.6151
R23307 VDD.n2167 VDD.n2166 10.6151
R23308 VDD.n2168 VDD.n2167 10.6151
R23309 VDD.n2168 VDD.n1034 10.6151
R23310 VDD.n2178 VDD.n1034 10.6151
R23311 VDD.n2179 VDD.n2178 10.6151
R23312 VDD.n2180 VDD.n2179 10.6151
R23313 VDD.n2180 VDD.n1022 10.6151
R23314 VDD.n2190 VDD.n1022 10.6151
R23315 VDD.n2191 VDD.n2190 10.6151
R23316 VDD.n2192 VDD.n2191 10.6151
R23317 VDD.n2192 VDD.n1010 10.6151
R23318 VDD.n2202 VDD.n1010 10.6151
R23319 VDD.n2203 VDD.n2202 10.6151
R23320 VDD.n2204 VDD.n2203 10.6151
R23321 VDD.n2204 VDD.n998 10.6151
R23322 VDD.n2214 VDD.n998 10.6151
R23323 VDD.n2215 VDD.n2214 10.6151
R23324 VDD.n2216 VDD.n2215 10.6151
R23325 VDD.n2216 VDD.n986 10.6151
R23326 VDD.n2226 VDD.n986 10.6151
R23327 VDD.n2227 VDD.n2226 10.6151
R23328 VDD.n2228 VDD.n2227 10.6151
R23329 VDD.n2228 VDD.n974 10.6151
R23330 VDD.n2238 VDD.n974 10.6151
R23331 VDD.n2239 VDD.n2238 10.6151
R23332 VDD.n2240 VDD.n2239 10.6151
R23333 VDD.n2240 VDD.n962 10.6151
R23334 VDD.n2250 VDD.n962 10.6151
R23335 VDD.n2251 VDD.n2250 10.6151
R23336 VDD.n2252 VDD.n2251 10.6151
R23337 VDD.n2252 VDD.n949 10.6151
R23338 VDD.n2262 VDD.n949 10.6151
R23339 VDD.n2263 VDD.n2262 10.6151
R23340 VDD.n2264 VDD.n2263 10.6151
R23341 VDD.n2264 VDD.n938 10.6151
R23342 VDD.n2274 VDD.n938 10.6151
R23343 VDD.n2275 VDD.n2274 10.6151
R23344 VDD.n2276 VDD.n2275 10.6151
R23345 VDD.n2276 VDD.n926 10.6151
R23346 VDD.n2286 VDD.n926 10.6151
R23347 VDD.n2287 VDD.n2286 10.6151
R23348 VDD.n2288 VDD.n2287 10.6151
R23349 VDD.n2288 VDD.n914 10.6151
R23350 VDD.n2298 VDD.n914 10.6151
R23351 VDD.n2299 VDD.n2298 10.6151
R23352 VDD.n2300 VDD.n2299 10.6151
R23353 VDD.n2300 VDD.n902 10.6151
R23354 VDD.n2310 VDD.n902 10.6151
R23355 VDD.n2311 VDD.n2310 10.6151
R23356 VDD.n2312 VDD.n2311 10.6151
R23357 VDD.n2312 VDD.n890 10.6151
R23358 VDD.n2322 VDD.n890 10.6151
R23359 VDD.n2323 VDD.n2322 10.6151
R23360 VDD.n2324 VDD.n2323 10.6151
R23361 VDD.n2324 VDD.n878 10.6151
R23362 VDD.n2334 VDD.n878 10.6151
R23363 VDD.n2335 VDD.n2334 10.6151
R23364 VDD.n2336 VDD.n2335 10.6151
R23365 VDD.n2336 VDD.n866 10.6151
R23366 VDD.n2346 VDD.n866 10.6151
R23367 VDD.n2347 VDD.n2346 10.6151
R23368 VDD.n2348 VDD.n2347 10.6151
R23369 VDD.n2348 VDD.n854 10.6151
R23370 VDD.n2358 VDD.n854 10.6151
R23371 VDD.n2359 VDD.n2358 10.6151
R23372 VDD.n2360 VDD.n2359 10.6151
R23373 VDD.n2360 VDD.n842 10.6151
R23374 VDD.n2370 VDD.n842 10.6151
R23375 VDD.n2371 VDD.n2370 10.6151
R23376 VDD.n2372 VDD.n2371 10.6151
R23377 VDD.n2372 VDD.n829 10.6151
R23378 VDD.n2382 VDD.n829 10.6151
R23379 VDD.n2383 VDD.n2382 10.6151
R23380 VDD.n2384 VDD.n2383 10.6151
R23381 VDD.n2384 VDD.n818 10.6151
R23382 VDD.n2394 VDD.n818 10.6151
R23383 VDD.n2395 VDD.n2394 10.6151
R23384 VDD.n2396 VDD.n2395 10.6151
R23385 VDD.n2396 VDD.n806 10.6151
R23386 VDD.n2406 VDD.n806 10.6151
R23387 VDD.n2407 VDD.n2406 10.6151
R23388 VDD.n2408 VDD.n2407 10.6151
R23389 VDD.n2408 VDD.n794 10.6151
R23390 VDD.n2418 VDD.n794 10.6151
R23391 VDD.n2419 VDD.n2418 10.6151
R23392 VDD.n2420 VDD.n2419 10.6151
R23393 VDD.n2420 VDD.n782 10.6151
R23394 VDD.n2430 VDD.n782 10.6151
R23395 VDD.n2431 VDD.n2430 10.6151
R23396 VDD.n2432 VDD.n2431 10.6151
R23397 VDD.n2432 VDD.n770 10.6151
R23398 VDD.n2442 VDD.n770 10.6151
R23399 VDD.n2443 VDD.n2442 10.6151
R23400 VDD.n2444 VDD.n2443 10.6151
R23401 VDD.n2444 VDD.n759 10.6151
R23402 VDD.n2454 VDD.n759 10.6151
R23403 VDD.n2455 VDD.n2454 10.6151
R23404 VDD.n2456 VDD.n2455 10.6151
R23405 VDD.n2456 VDD.n746 10.6151
R23406 VDD.n2504 VDD.n746 10.6151
R23407 VDD.n2505 VDD.n2504 10.6151
R23408 VDD.n2506 VDD.n2505 10.6151
R23409 VDD.n2506 VDD.n736 10.6151
R23410 VDD.n2548 VDD.n736 10.6151
R23411 VDD.n2548 VDD.n2547 10.6151
R23412 VDD.n2546 VDD.n2544 10.6151
R23413 VDD.n2544 VDD.n2541 10.6151
R23414 VDD.n2541 VDD.n2540 10.6151
R23415 VDD.n2540 VDD.n2537 10.6151
R23416 VDD.n2537 VDD.n2536 10.6151
R23417 VDD.n2536 VDD.n2533 10.6151
R23418 VDD.n2533 VDD.n2532 10.6151
R23419 VDD.n2532 VDD.n2529 10.6151
R23420 VDD.n2529 VDD.n2528 10.6151
R23421 VDD.n2528 VDD.n2525 10.6151
R23422 VDD.n2525 VDD.n2524 10.6151
R23423 VDD.n2521 VDD.n2520 10.6151
R23424 VDD.n2520 VDD.n2517 10.6151
R23425 VDD.n2517 VDD.n2516 10.6151
R23426 VDD.n1716 VDD.n1714 10.6151
R23427 VDD.n1717 VDD.n1716 10.6151
R23428 VDD.n1719 VDD.n1717 10.6151
R23429 VDD.n1720 VDD.n1719 10.6151
R23430 VDD.n1722 VDD.n1720 10.6151
R23431 VDD.n1723 VDD.n1722 10.6151
R23432 VDD.n1725 VDD.n1723 10.6151
R23433 VDD.n1726 VDD.n1725 10.6151
R23434 VDD.n1728 VDD.n1726 10.6151
R23435 VDD.n1729 VDD.n1728 10.6151
R23436 VDD.n1731 VDD.n1729 10.6151
R23437 VDD.n1732 VDD.n1731 10.6151
R23438 VDD.n1734 VDD.n1732 10.6151
R23439 VDD.n1735 VDD.n1734 10.6151
R23440 VDD.n1737 VDD.n1735 10.6151
R23441 VDD.n1738 VDD.n1737 10.6151
R23442 VDD.n1740 VDD.n1738 10.6151
R23443 VDD.n1741 VDD.n1740 10.6151
R23444 VDD.n1743 VDD.n1741 10.6151
R23445 VDD.n1744 VDD.n1743 10.6151
R23446 VDD.n1746 VDD.n1744 10.6151
R23447 VDD.n1747 VDD.n1746 10.6151
R23448 VDD.n1749 VDD.n1747 10.6151
R23449 VDD.n1750 VDD.n1749 10.6151
R23450 VDD.n1752 VDD.n1750 10.6151
R23451 VDD.n1753 VDD.n1752 10.6151
R23452 VDD.n1755 VDD.n1753 10.6151
R23453 VDD.n1756 VDD.n1755 10.6151
R23454 VDD.n1758 VDD.n1756 10.6151
R23455 VDD.n1759 VDD.n1758 10.6151
R23456 VDD.n1761 VDD.n1759 10.6151
R23457 VDD.n1762 VDD.n1761 10.6151
R23458 VDD.n1764 VDD.n1762 10.6151
R23459 VDD.n1765 VDD.n1764 10.6151
R23460 VDD.n1767 VDD.n1765 10.6151
R23461 VDD.n1768 VDD.n1767 10.6151
R23462 VDD.n1770 VDD.n1768 10.6151
R23463 VDD.n1771 VDD.n1770 10.6151
R23464 VDD.n1773 VDD.n1771 10.6151
R23465 VDD.n1774 VDD.n1773 10.6151
R23466 VDD.n1776 VDD.n1774 10.6151
R23467 VDD.n1777 VDD.n1776 10.6151
R23468 VDD.n1779 VDD.n1777 10.6151
R23469 VDD.n1780 VDD.n1779 10.6151
R23470 VDD.n1782 VDD.n1780 10.6151
R23471 VDD.n1783 VDD.n1782 10.6151
R23472 VDD.n1785 VDD.n1783 10.6151
R23473 VDD.n1786 VDD.n1785 10.6151
R23474 VDD.n1788 VDD.n1786 10.6151
R23475 VDD.n1789 VDD.n1788 10.6151
R23476 VDD.n1791 VDD.n1789 10.6151
R23477 VDD.n1792 VDD.n1791 10.6151
R23478 VDD.n1794 VDD.n1792 10.6151
R23479 VDD.n1795 VDD.n1794 10.6151
R23480 VDD.n1797 VDD.n1795 10.6151
R23481 VDD.n1798 VDD.n1797 10.6151
R23482 VDD.n1800 VDD.n1798 10.6151
R23483 VDD.n1801 VDD.n1800 10.6151
R23484 VDD.n1803 VDD.n1801 10.6151
R23485 VDD.n1804 VDD.n1803 10.6151
R23486 VDD.n1806 VDD.n1804 10.6151
R23487 VDD.n1807 VDD.n1806 10.6151
R23488 VDD.n1809 VDD.n1807 10.6151
R23489 VDD.n1810 VDD.n1809 10.6151
R23490 VDD.n1812 VDD.n1810 10.6151
R23491 VDD.n1813 VDD.n1812 10.6151
R23492 VDD.n1815 VDD.n1813 10.6151
R23493 VDD.n1816 VDD.n1815 10.6151
R23494 VDD.n1818 VDD.n1816 10.6151
R23495 VDD.n1819 VDD.n1818 10.6151
R23496 VDD.n1821 VDD.n1819 10.6151
R23497 VDD.n1822 VDD.n1821 10.6151
R23498 VDD.n1824 VDD.n1822 10.6151
R23499 VDD.n1825 VDD.n1824 10.6151
R23500 VDD.n1827 VDD.n1825 10.6151
R23501 VDD.n1828 VDD.n1827 10.6151
R23502 VDD.n1830 VDD.n1828 10.6151
R23503 VDD.n1831 VDD.n1830 10.6151
R23504 VDD.n1833 VDD.n1831 10.6151
R23505 VDD.n1834 VDD.n1833 10.6151
R23506 VDD.n1836 VDD.n1834 10.6151
R23507 VDD.n1837 VDD.n1836 10.6151
R23508 VDD.n1839 VDD.n1837 10.6151
R23509 VDD.n1840 VDD.n1839 10.6151
R23510 VDD.n1842 VDD.n1840 10.6151
R23511 VDD.n1843 VDD.n1842 10.6151
R23512 VDD.n1845 VDD.n1843 10.6151
R23513 VDD.n1846 VDD.n1845 10.6151
R23514 VDD.n1848 VDD.n1846 10.6151
R23515 VDD.n1849 VDD.n1848 10.6151
R23516 VDD.n1851 VDD.n1849 10.6151
R23517 VDD.n1852 VDD.n1851 10.6151
R23518 VDD.n1854 VDD.n1852 10.6151
R23519 VDD.n1855 VDD.n1854 10.6151
R23520 VDD.n1857 VDD.n1855 10.6151
R23521 VDD.n1858 VDD.n1857 10.6151
R23522 VDD.n1860 VDD.n1858 10.6151
R23523 VDD.n1861 VDD.n1860 10.6151
R23524 VDD.n1863 VDD.n1861 10.6151
R23525 VDD.n1864 VDD.n1863 10.6151
R23526 VDD.n1866 VDD.n1864 10.6151
R23527 VDD.n1867 VDD.n1866 10.6151
R23528 VDD.n1869 VDD.n1867 10.6151
R23529 VDD.n1870 VDD.n1869 10.6151
R23530 VDD.n1872 VDD.n1870 10.6151
R23531 VDD.n1873 VDD.n1872 10.6151
R23532 VDD.n1875 VDD.n1873 10.6151
R23533 VDD.n1876 VDD.n1875 10.6151
R23534 VDD.n1878 VDD.n1876 10.6151
R23535 VDD.n1879 VDD.n1878 10.6151
R23536 VDD.n1881 VDD.n1879 10.6151
R23537 VDD.n1882 VDD.n1881 10.6151
R23538 VDD.n1894 VDD.n1882 10.6151
R23539 VDD.n1894 VDD.n1893 10.6151
R23540 VDD.n1893 VDD.n1892 10.6151
R23541 VDD.n1892 VDD.n1890 10.6151
R23542 VDD.n1890 VDD.n1889 10.6151
R23543 VDD.n1889 VDD.n1887 10.6151
R23544 VDD.n1887 VDD.n1886 10.6151
R23545 VDD.n1886 VDD.n1884 10.6151
R23546 VDD.n1884 VDD.n1883 10.6151
R23547 VDD.n1883 VDD.n740 10.6151
R23548 VDD.n2511 VDD.n740 10.6151
R23549 VDD.n2512 VDD.n2511 10.6151
R23550 VDD.n2513 VDD.n2512 10.6151
R23551 VDD.n1144 VDD.n1106 10.6151
R23552 VDD.n1144 VDD.n1143 10.6151
R23553 VDD.n1150 VDD.n1143 10.6151
R23554 VDD.n1151 VDD.n1150 10.6151
R23555 VDD.n1152 VDD.n1151 10.6151
R23556 VDD.n1152 VDD.n1141 10.6151
R23557 VDD.n1158 VDD.n1141 10.6151
R23558 VDD.n1699 VDD.n1698 10.6151
R23559 VDD.n1699 VDD.n1139 10.6151
R23560 VDD.n1705 VDD.n1139 10.6151
R23561 VDD.n1708 VDD.n1707 10.6151
R23562 VDD.n1708 VDD.n1135 10.6151
R23563 VDD.n1713 VDD.n1135 10.6151
R23564 VDD.n2491 VDD.n2490 10.6151
R23565 VDD.n2490 VDD.n2487 10.6151
R23566 VDD.n2487 VDD.n2486 10.6151
R23567 VDD.n2486 VDD.n2483 10.6151
R23568 VDD.n2483 VDD.n2482 10.6151
R23569 VDD.n2482 VDD.n2479 10.6151
R23570 VDD.n2479 VDD.n2478 10.6151
R23571 VDD.n2478 VDD.n2475 10.6151
R23572 VDD.n2475 VDD.n2474 10.6151
R23573 VDD.n2474 VDD.n2471 10.6151
R23574 VDD.n2471 VDD.n2470 10.6151
R23575 VDD.n2467 VDD.n2466 10.6151
R23576 VDD.n2466 VDD.n728 10.6151
R23577 VDD.n2554 VDD.n728 10.6151
R23578 VDD.n2067 VDD.n2066 10.6151
R23579 VDD.n2066 VDD.n2064 10.6151
R23580 VDD.n2064 VDD.n2063 10.6151
R23581 VDD.n2063 VDD.n2061 10.6151
R23582 VDD.n2061 VDD.n2060 10.6151
R23583 VDD.n2060 VDD.n2058 10.6151
R23584 VDD.n2058 VDD.n2057 10.6151
R23585 VDD.n2057 VDD.n2055 10.6151
R23586 VDD.n2055 VDD.n2054 10.6151
R23587 VDD.n2054 VDD.n2052 10.6151
R23588 VDD.n2052 VDD.n2051 10.6151
R23589 VDD.n2051 VDD.n2049 10.6151
R23590 VDD.n2049 VDD.n2048 10.6151
R23591 VDD.n2048 VDD.n2046 10.6151
R23592 VDD.n2046 VDD.n2045 10.6151
R23593 VDD.n2045 VDD.n2043 10.6151
R23594 VDD.n2043 VDD.n2042 10.6151
R23595 VDD.n2042 VDD.n2040 10.6151
R23596 VDD.n2040 VDD.n2039 10.6151
R23597 VDD.n2039 VDD.n2037 10.6151
R23598 VDD.n2037 VDD.n2036 10.6151
R23599 VDD.n2036 VDD.n2034 10.6151
R23600 VDD.n2034 VDD.n2033 10.6151
R23601 VDD.n2033 VDD.n2031 10.6151
R23602 VDD.n2031 VDD.n2030 10.6151
R23603 VDD.n2030 VDD.n2028 10.6151
R23604 VDD.n2028 VDD.n2027 10.6151
R23605 VDD.n2027 VDD.n2025 10.6151
R23606 VDD.n2025 VDD.n2024 10.6151
R23607 VDD.n2024 VDD.n2022 10.6151
R23608 VDD.n2022 VDD.n2021 10.6151
R23609 VDD.n2021 VDD.n2019 10.6151
R23610 VDD.n2019 VDD.n2018 10.6151
R23611 VDD.n2018 VDD.n2016 10.6151
R23612 VDD.n2016 VDD.n2015 10.6151
R23613 VDD.n2015 VDD.n2013 10.6151
R23614 VDD.n2013 VDD.n2012 10.6151
R23615 VDD.n2012 VDD.n2010 10.6151
R23616 VDD.n2010 VDD.n2009 10.6151
R23617 VDD.n2009 VDD.n2007 10.6151
R23618 VDD.n2007 VDD.n2006 10.6151
R23619 VDD.n2006 VDD.n2004 10.6151
R23620 VDD.n2004 VDD.n2003 10.6151
R23621 VDD.n2003 VDD.n2001 10.6151
R23622 VDD.n2001 VDD.n2000 10.6151
R23623 VDD.n2000 VDD.n1998 10.6151
R23624 VDD.n1998 VDD.n1997 10.6151
R23625 VDD.n1997 VDD.n1995 10.6151
R23626 VDD.n1995 VDD.n1994 10.6151
R23627 VDD.n1994 VDD.n1992 10.6151
R23628 VDD.n1992 VDD.n1991 10.6151
R23629 VDD.n1991 VDD.n1989 10.6151
R23630 VDD.n1989 VDD.n1988 10.6151
R23631 VDD.n1988 VDD.n1986 10.6151
R23632 VDD.n1986 VDD.n1985 10.6151
R23633 VDD.n1985 VDD.n1983 10.6151
R23634 VDD.n1983 VDD.n1982 10.6151
R23635 VDD.n1982 VDD.n1980 10.6151
R23636 VDD.n1980 VDD.n1979 10.6151
R23637 VDD.n1979 VDD.n1977 10.6151
R23638 VDD.n1977 VDD.n1976 10.6151
R23639 VDD.n1976 VDD.n1974 10.6151
R23640 VDD.n1974 VDD.n1973 10.6151
R23641 VDD.n1973 VDD.n1971 10.6151
R23642 VDD.n1971 VDD.n1970 10.6151
R23643 VDD.n1970 VDD.n1968 10.6151
R23644 VDD.n1968 VDD.n1967 10.6151
R23645 VDD.n1967 VDD.n1965 10.6151
R23646 VDD.n1965 VDD.n1964 10.6151
R23647 VDD.n1964 VDD.n1962 10.6151
R23648 VDD.n1962 VDD.n1961 10.6151
R23649 VDD.n1961 VDD.n1959 10.6151
R23650 VDD.n1959 VDD.n1958 10.6151
R23651 VDD.n1958 VDD.n1956 10.6151
R23652 VDD.n1956 VDD.n1955 10.6151
R23653 VDD.n1955 VDD.n1953 10.6151
R23654 VDD.n1953 VDD.n1952 10.6151
R23655 VDD.n1952 VDD.n1950 10.6151
R23656 VDD.n1950 VDD.n1949 10.6151
R23657 VDD.n1949 VDD.n1947 10.6151
R23658 VDD.n1947 VDD.n1946 10.6151
R23659 VDD.n1946 VDD.n1944 10.6151
R23660 VDD.n1944 VDD.n1943 10.6151
R23661 VDD.n1943 VDD.n1941 10.6151
R23662 VDD.n1941 VDD.n1940 10.6151
R23663 VDD.n1940 VDD.n1938 10.6151
R23664 VDD.n1938 VDD.n1937 10.6151
R23665 VDD.n1937 VDD.n1935 10.6151
R23666 VDD.n1935 VDD.n1934 10.6151
R23667 VDD.n1934 VDD.n1932 10.6151
R23668 VDD.n1932 VDD.n1931 10.6151
R23669 VDD.n1931 VDD.n1929 10.6151
R23670 VDD.n1929 VDD.n1928 10.6151
R23671 VDD.n1928 VDD.n1926 10.6151
R23672 VDD.n1926 VDD.n1925 10.6151
R23673 VDD.n1925 VDD.n1923 10.6151
R23674 VDD.n1923 VDD.n1922 10.6151
R23675 VDD.n1922 VDD.n1920 10.6151
R23676 VDD.n1920 VDD.n1919 10.6151
R23677 VDD.n1919 VDD.n1917 10.6151
R23678 VDD.n1917 VDD.n1916 10.6151
R23679 VDD.n1916 VDD.n1914 10.6151
R23680 VDD.n1914 VDD.n1913 10.6151
R23681 VDD.n1913 VDD.n1911 10.6151
R23682 VDD.n1911 VDD.n1910 10.6151
R23683 VDD.n1910 VDD.n1908 10.6151
R23684 VDD.n1908 VDD.n1907 10.6151
R23685 VDD.n1907 VDD.n1905 10.6151
R23686 VDD.n1905 VDD.n1904 10.6151
R23687 VDD.n1904 VDD.n1902 10.6151
R23688 VDD.n1902 VDD.n1901 10.6151
R23689 VDD.n1901 VDD.n1899 10.6151
R23690 VDD.n1899 VDD.n1898 10.6151
R23691 VDD.n1898 VDD.n1134 10.6151
R23692 VDD.n1134 VDD.n1133 10.6151
R23693 VDD.n1133 VDD.n1131 10.6151
R23694 VDD.n1131 VDD.n1130 10.6151
R23695 VDD.n1130 VDD.n1128 10.6151
R23696 VDD.n1128 VDD.n1127 10.6151
R23697 VDD.n1127 VDD.n1125 10.6151
R23698 VDD.n1125 VDD.n1124 10.6151
R23699 VDD.n1124 VDD.n1122 10.6151
R23700 VDD.n1122 VDD.n729 10.6151
R23701 VDD.n2552 VDD.n729 10.6151
R23702 VDD.n2553 VDD.n2552 10.6151
R23703 VDD.n2101 VDD.n2100 10.6151
R23704 VDD.n2100 VDD.n1112 10.6151
R23705 VDD.n2094 VDD.n1112 10.6151
R23706 VDD.n2094 VDD.n2093 10.6151
R23707 VDD.n2093 VDD.n2092 10.6151
R23708 VDD.n2092 VDD.n1114 10.6151
R23709 VDD.n2086 VDD.n1114 10.6151
R23710 VDD.n2084 VDD.n2083 10.6151
R23711 VDD.n2083 VDD.n1117 10.6151
R23712 VDD.n2077 VDD.n1117 10.6151
R23713 VDD.n2075 VDD.n2074 10.6151
R23714 VDD.n2074 VDD.n1121 10.6151
R23715 VDD.n2068 VDD.n1121 10.6151
R23716 VDD.n2102 VDD.n1100 10.6151
R23717 VDD.n2112 VDD.n1100 10.6151
R23718 VDD.n2113 VDD.n2112 10.6151
R23719 VDD.n2114 VDD.n2113 10.6151
R23720 VDD.n2114 VDD.n1088 10.6151
R23721 VDD.n2124 VDD.n1088 10.6151
R23722 VDD.n2125 VDD.n2124 10.6151
R23723 VDD.n2126 VDD.n2125 10.6151
R23724 VDD.n2126 VDD.n1075 10.6151
R23725 VDD.n2136 VDD.n1075 10.6151
R23726 VDD.n2137 VDD.n2136 10.6151
R23727 VDD.n2138 VDD.n2137 10.6151
R23728 VDD.n2138 VDD.n1064 10.6151
R23729 VDD.n2148 VDD.n1064 10.6151
R23730 VDD.n2149 VDD.n2148 10.6151
R23731 VDD.n2150 VDD.n2149 10.6151
R23732 VDD.n2150 VDD.n1052 10.6151
R23733 VDD.n2160 VDD.n1052 10.6151
R23734 VDD.n2161 VDD.n2160 10.6151
R23735 VDD.n2162 VDD.n2161 10.6151
R23736 VDD.n2162 VDD.n1040 10.6151
R23737 VDD.n2172 VDD.n1040 10.6151
R23738 VDD.n2173 VDD.n2172 10.6151
R23739 VDD.n2174 VDD.n2173 10.6151
R23740 VDD.n2174 VDD.n1027 10.6151
R23741 VDD.n2184 VDD.n1027 10.6151
R23742 VDD.n2185 VDD.n2184 10.6151
R23743 VDD.n2186 VDD.n2185 10.6151
R23744 VDD.n2186 VDD.n1016 10.6151
R23745 VDD.n2196 VDD.n1016 10.6151
R23746 VDD.n2197 VDD.n2196 10.6151
R23747 VDD.n2198 VDD.n2197 10.6151
R23748 VDD.n2198 VDD.n1004 10.6151
R23749 VDD.n2208 VDD.n1004 10.6151
R23750 VDD.n2209 VDD.n2208 10.6151
R23751 VDD.n2210 VDD.n2209 10.6151
R23752 VDD.n2210 VDD.n992 10.6151
R23753 VDD.n2220 VDD.n992 10.6151
R23754 VDD.n2221 VDD.n2220 10.6151
R23755 VDD.n2222 VDD.n2221 10.6151
R23756 VDD.n2222 VDD.n980 10.6151
R23757 VDD.n2232 VDD.n980 10.6151
R23758 VDD.n2233 VDD.n2232 10.6151
R23759 VDD.n2234 VDD.n2233 10.6151
R23760 VDD.n2234 VDD.n968 10.6151
R23761 VDD.n2244 VDD.n968 10.6151
R23762 VDD.n2245 VDD.n2244 10.6151
R23763 VDD.n2246 VDD.n2245 10.6151
R23764 VDD.n2246 VDD.n956 10.6151
R23765 VDD.n2256 VDD.n956 10.6151
R23766 VDD.n2257 VDD.n2256 10.6151
R23767 VDD.n2258 VDD.n2257 10.6151
R23768 VDD.n2258 VDD.n943 10.6151
R23769 VDD.n2268 VDD.n943 10.6151
R23770 VDD.n2269 VDD.n2268 10.6151
R23771 VDD.n2270 VDD.n2269 10.6151
R23772 VDD.n2270 VDD.n932 10.6151
R23773 VDD.n2280 VDD.n932 10.6151
R23774 VDD.n2281 VDD.n2280 10.6151
R23775 VDD.n2282 VDD.n2281 10.6151
R23776 VDD.n2282 VDD.n920 10.6151
R23777 VDD.n2292 VDD.n920 10.6151
R23778 VDD.n2293 VDD.n2292 10.6151
R23779 VDD.n2294 VDD.n2293 10.6151
R23780 VDD.n2294 VDD.n908 10.6151
R23781 VDD.n2304 VDD.n908 10.6151
R23782 VDD.n2305 VDD.n2304 10.6151
R23783 VDD.n2306 VDD.n2305 10.6151
R23784 VDD.n2306 VDD.n895 10.6151
R23785 VDD.n2316 VDD.n895 10.6151
R23786 VDD.n2317 VDD.n2316 10.6151
R23787 VDD.n2318 VDD.n2317 10.6151
R23788 VDD.n2318 VDD.n884 10.6151
R23789 VDD.n2328 VDD.n884 10.6151
R23790 VDD.n2329 VDD.n2328 10.6151
R23791 VDD.n2330 VDD.n2329 10.6151
R23792 VDD.n2330 VDD.n872 10.6151
R23793 VDD.n2340 VDD.n872 10.6151
R23794 VDD.n2341 VDD.n2340 10.6151
R23795 VDD.n2342 VDD.n2341 10.6151
R23796 VDD.n2342 VDD.n860 10.6151
R23797 VDD.n2352 VDD.n860 10.6151
R23798 VDD.n2353 VDD.n2352 10.6151
R23799 VDD.n2354 VDD.n2353 10.6151
R23800 VDD.n2354 VDD.n848 10.6151
R23801 VDD.n2364 VDD.n848 10.6151
R23802 VDD.n2365 VDD.n2364 10.6151
R23803 VDD.n2366 VDD.n2365 10.6151
R23804 VDD.n2366 VDD.n836 10.6151
R23805 VDD.n2376 VDD.n836 10.6151
R23806 VDD.n2377 VDD.n2376 10.6151
R23807 VDD.n2378 VDD.n2377 10.6151
R23808 VDD.n2378 VDD.n824 10.6151
R23809 VDD.n2388 VDD.n824 10.6151
R23810 VDD.n2389 VDD.n2388 10.6151
R23811 VDD.n2390 VDD.n2389 10.6151
R23812 VDD.n2390 VDD.n812 10.6151
R23813 VDD.n2400 VDD.n812 10.6151
R23814 VDD.n2401 VDD.n2400 10.6151
R23815 VDD.n2402 VDD.n2401 10.6151
R23816 VDD.n2402 VDD.n800 10.6151
R23817 VDD.n2412 VDD.n800 10.6151
R23818 VDD.n2413 VDD.n2412 10.6151
R23819 VDD.n2414 VDD.n2413 10.6151
R23820 VDD.n2414 VDD.n788 10.6151
R23821 VDD.n2424 VDD.n788 10.6151
R23822 VDD.n2425 VDD.n2424 10.6151
R23823 VDD.n2426 VDD.n2425 10.6151
R23824 VDD.n2426 VDD.n776 10.6151
R23825 VDD.n2436 VDD.n776 10.6151
R23826 VDD.n2437 VDD.n2436 10.6151
R23827 VDD.n2438 VDD.n2437 10.6151
R23828 VDD.n2438 VDD.n765 10.6151
R23829 VDD.n2448 VDD.n765 10.6151
R23830 VDD.n2449 VDD.n2448 10.6151
R23831 VDD.n2450 VDD.n2449 10.6151
R23832 VDD.n2450 VDD.n753 10.6151
R23833 VDD.n2460 VDD.n753 10.6151
R23834 VDD.n2461 VDD.n2460 10.6151
R23835 VDD.n2500 VDD.n2461 10.6151
R23836 VDD.n2500 VDD.n2499 10.6151
R23837 VDD.n2499 VDD.n2498 10.6151
R23838 VDD.n2498 VDD.n2497 10.6151
R23839 VDD.n2497 VDD.n2495 10.6151
R23840 VDD.n2495 VDD.n2494 10.6151
R23841 VDD.n1422 VDD.n1372 9.89141
R23842 VDD.n3499 VDD.n3498 9.89141
R23843 VDD.n147 VDD.n146 9.89141
R23844 VDD.n1658 VDD.n1191 9.89141
R23845 VDD.n3532 VDD.n3531 9.3005
R23846 VDD.n3533 VDD.n252 9.3005
R23847 VDD.n3535 VDD.n3534 9.3005
R23848 VDD.n242 VDD.n241 9.3005
R23849 VDD.n3548 VDD.n3547 9.3005
R23850 VDD.n3549 VDD.n240 9.3005
R23851 VDD.n3551 VDD.n3550 9.3005
R23852 VDD.n230 VDD.n229 9.3005
R23853 VDD.n3564 VDD.n3563 9.3005
R23854 VDD.n3565 VDD.n228 9.3005
R23855 VDD.n3567 VDD.n3566 9.3005
R23856 VDD.n218 VDD.n217 9.3005
R23857 VDD.n3580 VDD.n3579 9.3005
R23858 VDD.n3581 VDD.n216 9.3005
R23859 VDD.n3585 VDD.n3582 9.3005
R23860 VDD.n3584 VDD.n3583 9.3005
R23861 VDD.n206 VDD.n205 9.3005
R23862 VDD.n3599 VDD.n3598 9.3005
R23863 VDD.n3600 VDD.n204 9.3005
R23864 VDD.n3605 VDD.n3601 9.3005
R23865 VDD.n3604 VDD.n3603 9.3005
R23866 VDD.n3602 VDD.n193 9.3005
R23867 VDD.n3620 VDD.n194 9.3005
R23868 VDD.n3621 VDD.n192 9.3005
R23869 VDD.n3623 VDD.n3622 9.3005
R23870 VDD.n3624 VDD.n191 9.3005
R23871 VDD.n3627 VDD.n3625 9.3005
R23872 VDD.n3628 VDD.n190 9.3005
R23873 VDD.n3630 VDD.n3629 9.3005
R23874 VDD.n3631 VDD.n189 9.3005
R23875 VDD.n3634 VDD.n3632 9.3005
R23876 VDD.n3635 VDD.n188 9.3005
R23877 VDD.n3637 VDD.n3636 9.3005
R23878 VDD.n3638 VDD.n187 9.3005
R23879 VDD.n3641 VDD.n3639 9.3005
R23880 VDD.n3642 VDD.n186 9.3005
R23881 VDD.n3644 VDD.n3643 9.3005
R23882 VDD.n3645 VDD.n185 9.3005
R23883 VDD.n3648 VDD.n3646 9.3005
R23884 VDD.n3649 VDD.n184 9.3005
R23885 VDD.n3651 VDD.n3650 9.3005
R23886 VDD.n3652 VDD.n183 9.3005
R23887 VDD.n3655 VDD.n3653 9.3005
R23888 VDD.n3656 VDD.n182 9.3005
R23889 VDD.n3658 VDD.n3657 9.3005
R23890 VDD.n254 VDD.n253 9.3005
R23891 VDD.n122 VDD.n121 9.3005
R23892 VDD.n123 VDD.n114 9.3005
R23893 VDD.n125 VDD.n124 9.3005
R23894 VDD.n128 VDD.n113 9.3005
R23895 VDD.n132 VDD.n131 9.3005
R23896 VDD.n133 VDD.n112 9.3005
R23897 VDD.n135 VDD.n134 9.3005
R23898 VDD.n138 VDD.n111 9.3005
R23899 VDD.n142 VDD.n141 9.3005
R23900 VDD.n143 VDD.n110 9.3005
R23901 VDD.n146 VDD.n144 9.3005
R23902 VDD.n147 VDD.n106 9.3005
R23903 VDD.n151 VDD.n150 9.3005
R23904 VDD.n152 VDD.n105 9.3005
R23905 VDD.n154 VDD.n153 9.3005
R23906 VDD.n157 VDD.n104 9.3005
R23907 VDD.n161 VDD.n160 9.3005
R23908 VDD.n162 VDD.n103 9.3005
R23909 VDD.n164 VDD.n163 9.3005
R23910 VDD.n167 VDD.n102 9.3005
R23911 VDD.n171 VDD.n170 9.3005
R23912 VDD.n172 VDD.n101 9.3005
R23913 VDD.n174 VDD.n173 9.3005
R23914 VDD.n177 VDD.n100 9.3005
R23915 VDD.n180 VDD.n179 9.3005
R23916 VDD.n181 VDD.n99 9.3005
R23917 VDD.n3660 VDD.n3659 9.3005
R23918 VDD.n118 VDD.n116 9.3005
R23919 VDD.n3709 VDD.n3708 9.3005
R23920 VDD.n3707 VDD.n20 9.3005
R23921 VDD.n31 VDD.n23 9.3005
R23922 VDD.n3701 VDD.n32 9.3005
R23923 VDD.n3700 VDD.n33 9.3005
R23924 VDD.n3699 VDD.n34 9.3005
R23925 VDD.n42 VDD.n35 9.3005
R23926 VDD.n3693 VDD.n43 9.3005
R23927 VDD.n3692 VDD.n44 9.3005
R23928 VDD.n3691 VDD.n45 9.3005
R23929 VDD.n53 VDD.n46 9.3005
R23930 VDD.n3685 VDD.n54 9.3005
R23931 VDD.n3684 VDD.n55 9.3005
R23932 VDD.n3683 VDD.n56 9.3005
R23933 VDD.n64 VDD.n57 9.3005
R23934 VDD.n3677 VDD.n65 9.3005
R23935 VDD.n3676 VDD.n66 9.3005
R23936 VDD.n3675 VDD.n67 9.3005
R23937 VDD.n75 VDD.n68 9.3005
R23938 VDD.n3669 VDD.n76 9.3005
R23939 VDD.n3668 VDD.n77 9.3005
R23940 VDD.n3667 VDD.n78 9.3005
R23941 VDD.n115 VDD.n79 9.3005
R23942 VDD.n3527 VDD.n3526 9.3005
R23943 VDD.n248 VDD.n247 9.3005
R23944 VDD.n3540 VDD.n3539 9.3005
R23945 VDD.n3541 VDD.n246 9.3005
R23946 VDD.n3543 VDD.n3542 9.3005
R23947 VDD.n236 VDD.n235 9.3005
R23948 VDD.n3556 VDD.n3555 9.3005
R23949 VDD.n3557 VDD.n234 9.3005
R23950 VDD.n3559 VDD.n3558 9.3005
R23951 VDD.n224 VDD.n223 9.3005
R23952 VDD.n3572 VDD.n3571 9.3005
R23953 VDD.n3573 VDD.n222 9.3005
R23954 VDD.n3575 VDD.n3574 9.3005
R23955 VDD.n212 VDD.n211 9.3005
R23956 VDD.n3590 VDD.n3589 9.3005
R23957 VDD.n3591 VDD.n210 9.3005
R23958 VDD.n3593 VDD.n3592 9.3005
R23959 VDD.n200 VDD.n199 9.3005
R23960 VDD.n3611 VDD.n3610 9.3005
R23961 VDD.n3612 VDD.n198 9.3005
R23962 VDD.n3614 VDD.n3613 9.3005
R23963 VDD.n21 VDD.n19 9.3005
R23964 VDD.n3525 VDD.n258 9.3005
R23965 VDD.n3472 VDD.n3471 9.3005
R23966 VDD.n3475 VDD.n303 9.3005
R23967 VDD.n3476 VDD.n302 9.3005
R23968 VDD.n3479 VDD.n301 9.3005
R23969 VDD.n3480 VDD.n300 9.3005
R23970 VDD.n3483 VDD.n299 9.3005
R23971 VDD.n3484 VDD.n298 9.3005
R23972 VDD.n3487 VDD.n297 9.3005
R23973 VDD.n3488 VDD.n296 9.3005
R23974 VDD.n3491 VDD.n295 9.3005
R23975 VDD.n3492 VDD.n294 9.3005
R23976 VDD.n3495 VDD.n293 9.3005
R23977 VDD.n3497 VDD.n292 9.3005
R23978 VDD.n3498 VDD.n289 9.3005
R23979 VDD.n3499 VDD.n287 9.3005
R23980 VDD.n3502 VDD.n286 9.3005
R23981 VDD.n3503 VDD.n285 9.3005
R23982 VDD.n3506 VDD.n284 9.3005
R23983 VDD.n3507 VDD.n283 9.3005
R23984 VDD.n3510 VDD.n282 9.3005
R23985 VDD.n3511 VDD.n281 9.3005
R23986 VDD.n3514 VDD.n280 9.3005
R23987 VDD.n3515 VDD.n279 9.3005
R23988 VDD.n3516 VDD.n278 9.3005
R23989 VDD.n262 VDD.n261 9.3005
R23990 VDD.n3522 VDD.n3521 9.3005
R23991 VDD.n3470 VDD.n307 9.3005
R23992 VDD.n3469 VDD.n3468 9.3005
R23993 VDD.n1541 VDD.n1540 9.3005
R23994 VDD.n1542 VDD.n1266 9.3005
R23995 VDD.n1544 VDD.n1543 9.3005
R23996 VDD.n1256 VDD.n1255 9.3005
R23997 VDD.n1557 VDD.n1556 9.3005
R23998 VDD.n1558 VDD.n1254 9.3005
R23999 VDD.n1560 VDD.n1559 9.3005
R24000 VDD.n1244 VDD.n1243 9.3005
R24001 VDD.n1573 VDD.n1572 9.3005
R24002 VDD.n1574 VDD.n1242 9.3005
R24003 VDD.n1576 VDD.n1575 9.3005
R24004 VDD.n1232 VDD.n1231 9.3005
R24005 VDD.n1589 VDD.n1588 9.3005
R24006 VDD.n1590 VDD.n1230 9.3005
R24007 VDD.n1592 VDD.n1591 9.3005
R24008 VDD.n1219 VDD.n1218 9.3005
R24009 VDD.n1606 VDD.n1605 9.3005
R24010 VDD.n1607 VDD.n1217 9.3005
R24011 VDD.n1609 VDD.n1608 9.3005
R24012 VDD.n1206 VDD.n1205 9.3005
R24013 VDD.n1627 VDD.n1626 9.3005
R24014 VDD.n1628 VDD.n1204 9.3005
R24015 VDD.n1630 VDD.n1629 9.3005
R24016 VDD.n1635 VDD.n1202 9.3005
R24017 VDD.n1639 VDD.n1638 9.3005
R24018 VDD.n1640 VDD.n1199 9.3005
R24019 VDD.n1642 VDD.n1641 9.3005
R24020 VDD.n1643 VDD.n1198 9.3005
R24021 VDD.n1647 VDD.n1646 9.3005
R24022 VDD.n1648 VDD.n1195 9.3005
R24023 VDD.n1650 VDD.n1649 9.3005
R24024 VDD.n1651 VDD.n1194 9.3005
R24025 VDD.n1655 VDD.n1654 9.3005
R24026 VDD.n1656 VDD.n1191 9.3005
R24027 VDD.n1658 VDD.n1657 9.3005
R24028 VDD.n1163 VDD.n1161 9.3005
R24029 VDD.n1694 VDD.n1693 9.3005
R24030 VDD.n1692 VDD.n1162 9.3005
R24031 VDD.n1691 VDD.n1690 9.3005
R24032 VDD.n1689 VDD.n1167 9.3005
R24033 VDD.n1688 VDD.n1687 9.3005
R24034 VDD.n1686 VDD.n1168 9.3005
R24035 VDD.n1685 VDD.n1684 9.3005
R24036 VDD.n1683 VDD.n1172 9.3005
R24037 VDD.n1682 VDD.n1681 9.3005
R24038 VDD.n1680 VDD.n1173 9.3005
R24039 VDD.n1679 VDD.n1678 9.3005
R24040 VDD.n1677 VDD.n1177 9.3005
R24041 VDD.n1676 VDD.n1675 9.3005
R24042 VDD.n1674 VDD.n1178 9.3005
R24043 VDD.n1634 VDD.n1633 9.3005
R24044 VDD.n1452 VDD.n1451 9.3005
R24045 VDD.n1453 VDD.n1336 9.3005
R24046 VDD.n1455 VDD.n1454 9.3005
R24047 VDD.n1326 VDD.n1325 9.3005
R24048 VDD.n1468 VDD.n1467 9.3005
R24049 VDD.n1469 VDD.n1324 9.3005
R24050 VDD.n1471 VDD.n1470 9.3005
R24051 VDD.n1314 VDD.n1313 9.3005
R24052 VDD.n1484 VDD.n1483 9.3005
R24053 VDD.n1485 VDD.n1312 9.3005
R24054 VDD.n1487 VDD.n1486 9.3005
R24055 VDD.n1302 VDD.n1301 9.3005
R24056 VDD.n1500 VDD.n1499 9.3005
R24057 VDD.n1501 VDD.n1300 9.3005
R24058 VDD.n1503 VDD.n1502 9.3005
R24059 VDD.n1290 VDD.n1289 9.3005
R24060 VDD.n1516 VDD.n1515 9.3005
R24061 VDD.n1517 VDD.n1288 9.3005
R24062 VDD.n1519 VDD.n1518 9.3005
R24063 VDD.n1278 VDD.n1277 9.3005
R24064 VDD.n1533 VDD.n1532 9.3005
R24065 VDD.n1534 VDD.n1276 9.3005
R24066 VDD.n1536 VDD.n1535 9.3005
R24067 VDD.n1262 VDD.n1261 9.3005
R24068 VDD.n1549 VDD.n1548 9.3005
R24069 VDD.n1550 VDD.n1260 9.3005
R24070 VDD.n1552 VDD.n1551 9.3005
R24071 VDD.n1250 VDD.n1249 9.3005
R24072 VDD.n1565 VDD.n1564 9.3005
R24073 VDD.n1566 VDD.n1248 9.3005
R24074 VDD.n1568 VDD.n1567 9.3005
R24075 VDD.n1238 VDD.n1237 9.3005
R24076 VDD.n1581 VDD.n1580 9.3005
R24077 VDD.n1582 VDD.n1236 9.3005
R24078 VDD.n1584 VDD.n1583 9.3005
R24079 VDD.n1226 VDD.n1225 9.3005
R24080 VDD.n1597 VDD.n1596 9.3005
R24081 VDD.n1598 VDD.n1223 9.3005
R24082 VDD.n1601 VDD.n1600 9.3005
R24083 VDD.n1599 VDD.n1224 9.3005
R24084 VDD.n1213 VDD.n1212 9.3005
R24085 VDD.n1615 VDD.n1614 9.3005
R24086 VDD.n1616 VDD.n1210 9.3005
R24087 VDD.n1621 VDD.n1620 9.3005
R24088 VDD.n1619 VDD.n1211 9.3005
R24089 VDD.n1338 VDD.n1337 9.3005
R24090 VDD.n1399 VDD.n1389 9.3005
R24091 VDD.n1401 VDD.n1400 9.3005
R24092 VDD.n1402 VDD.n1388 9.3005
R24093 VDD.n1404 VDD.n1403 9.3005
R24094 VDD.n1405 VDD.n1383 9.3005
R24095 VDD.n1407 VDD.n1406 9.3005
R24096 VDD.n1408 VDD.n1382 9.3005
R24097 VDD.n1410 VDD.n1409 9.3005
R24098 VDD.n1411 VDD.n1377 9.3005
R24099 VDD.n1413 VDD.n1412 9.3005
R24100 VDD.n1414 VDD.n1376 9.3005
R24101 VDD.n1416 VDD.n1415 9.3005
R24102 VDD.n1417 VDD.n1373 9.3005
R24103 VDD.n1423 VDD.n1422 9.3005
R24104 VDD.n1424 VDD.n1372 9.3005
R24105 VDD.n1426 VDD.n1425 9.3005
R24106 VDD.n1427 VDD.n1367 9.3005
R24107 VDD.n1429 VDD.n1428 9.3005
R24108 VDD.n1430 VDD.n1366 9.3005
R24109 VDD.n1432 VDD.n1431 9.3005
R24110 VDD.n1433 VDD.n1361 9.3005
R24111 VDD.n1435 VDD.n1434 9.3005
R24112 VDD.n1436 VDD.n1360 9.3005
R24113 VDD.n1438 VDD.n1437 9.3005
R24114 VDD.n1344 VDD.n1343 9.3005
R24115 VDD.n1444 VDD.n1443 9.3005
R24116 VDD.n1398 VDD.n1394 9.3005
R24117 VDD.n1393 VDD.n1392 9.3005
R24118 VDD.n1447 VDD.n1446 9.3005
R24119 VDD.n1332 VDD.n1331 9.3005
R24120 VDD.n1460 VDD.n1459 9.3005
R24121 VDD.n1461 VDD.n1330 9.3005
R24122 VDD.n1463 VDD.n1462 9.3005
R24123 VDD.n1320 VDD.n1319 9.3005
R24124 VDD.n1476 VDD.n1475 9.3005
R24125 VDD.n1477 VDD.n1318 9.3005
R24126 VDD.n1479 VDD.n1478 9.3005
R24127 VDD.n1308 VDD.n1307 9.3005
R24128 VDD.n1492 VDD.n1491 9.3005
R24129 VDD.n1493 VDD.n1306 9.3005
R24130 VDD.n1495 VDD.n1494 9.3005
R24131 VDD.n1296 VDD.n1295 9.3005
R24132 VDD.n1508 VDD.n1507 9.3005
R24133 VDD.n1509 VDD.n1294 9.3005
R24134 VDD.n1511 VDD.n1510 9.3005
R24135 VDD.n1284 VDD.n1283 9.3005
R24136 VDD.n1524 VDD.n1523 9.3005
R24137 VDD.n1525 VDD.n1282 9.3005
R24138 VDD.n1528 VDD.n1527 9.3005
R24139 VDD.n1526 VDD.n1272 9.3005
R24140 VDD.n1445 VDD.n1342 9.3005
R24141 VDD.n2128 VDD.t69 9.08952
R24142 VDD.t88 VDD.n356 9.08952
R24143 VDD.n1896 VDD.t81 8.89193
R24144 VDD.n3048 VDD.t93 8.89193
R24145 VDD.n2591 VDD.n2590 8.27367
R24146 VDD.n3419 VDD.n337 8.27367
R24147 VDD.n3455 VDD.n3454 8.27367
R24148 VDD.n2986 VDD.n2985 8.27367
R24149 VDD.n2524 VDD.n739 8.27367
R24150 VDD.n1706 VDD.n1705 8.27367
R24151 VDD.n2470 VDD.n2464 8.27367
R24152 VDD.n2077 VDD.n2076 8.27367
R24153 VDD.n15 VDD.n14 8.24655
R24154 VDD.n3711 VDD.n3710 8.16525
R24155 VDD.n1271 VDD.n1270 8.16525
R24156 VDD.n947 VDD.t84 8.10158
R24157 VDD.n3222 VDD.t100 8.10158
R24158 VDD.n1032 VDD.t79 7.90399
R24159 VDD.n3306 VDD.t105 7.90399
R24160 VDD.n2386 VDD.t71 7.70641
R24161 VDD.n622 VDD.t107 7.70641
R24162 VDD.n1398 VDD.n1392 7.56414
R24163 VDD.n3468 VDD.n307 7.56414
R24164 VDD.n3660 VDD.n99 7.56414
R24165 VDD.n1675 VDD.n1674 7.56414
R24166 VDD.n1465 VDD.t37 6.91606
R24167 VDD.t29 VDD.n1215 6.91606
R24168 VDD.n2326 VDD.t96 6.91606
R24169 VDD.t74 VDD.n553 6.91606
R24170 VDD.n3545 VDD.t50 6.91606
R24171 VDD.n3673 VDD.t13 6.91606
R24172 VDD.t96 VDD.n880 6.52088
R24173 VDD.n3162 VDD.t74 6.52088
R24174 VDD.n834 VDD.t71 5.73053
R24175 VDD.n3108 VDD.t107 5.73053
R24176 VDD.n18 VDD.n16 5.67579
R24177 VDD.n1269 VDD.n1267 5.67579
R24178 VDD.n2188 VDD.t79 5.53295
R24179 VDD.n424 VDD.t105 5.53295
R24180 VDD.t5 VDD.n1286 5.33536
R24181 VDD.n1554 VDD.t3 5.33536
R24182 VDD.n2272 VDD.t84 5.33536
R24183 VDD.n508 VDD.t100 5.33536
R24184 VDD.t1 VDD.n202 5.33536
R24185 VDD.t8 VDD.n29 5.33536
R24186 VDD.n3425 VDD.n260 5.30782
R24187 VDD.n333 VDD.n260 5.30782
R24188 VDD.n3463 VDD.n308 5.30782
R24189 VDD.n3463 VDD.n3462 5.30782
R24190 VDD.n1697 VDD.n1158 5.30782
R24191 VDD.n1698 VDD.n1697 5.30782
R24192 VDD.n2086 VDD.n2085 5.30782
R24193 VDD.n2085 VDD.n2084 5.30782
R24194 VDD.n3711 VDD.n18 4.74396
R24195 VDD.n1270 VDD.n1269 4.74396
R24196 VDD.n18 VDD.n17 4.63843
R24197 VDD.n1269 VDD.n1268 4.63843
R24198 VDD.n3466 VDD.n259 4.61026
R24199 VDD.n3524 VDD.n259 4.57367
R24200 VDD.n2440 VDD.t81 4.54501
R24201 VDD.t93 VDD.n668 4.54501
R24202 VDD.n1696 VDD.n1695 4.34806
R24203 VDD.n1695 VDD.n1160 4.34806
R24204 VDD.t69 VDD.n1077 4.34742
R24205 VDD.n3360 VDD.t88 4.34742
R24206 VDD.n1270 VDD.n15 2.54226
R24207 VDD VDD.n3711 2.53443
R24208 VDD.n2590 VDD.n2562 2.34196
R24209 VDD.n339 VDD.n337 2.34196
R24210 VDD.n3454 VDD.n3453 2.34196
R24211 VDD.n2985 VDD.n2984 2.34196
R24212 VDD.n2521 VDD.n739 2.34196
R24213 VDD.n1707 VDD.n1706 2.34196
R24214 VDD.n2467 VDD.n2464 2.34196
R24215 VDD.n2076 VDD.n2075 2.34196
R24216 VDD.n4 VDD.n2 2.29289
R24217 VDD.n11 VDD.n9 2.29289
R24218 VDD.n6 VDD.n4 1.8482
R24219 VDD.n13 VDD.n11 1.8482
R24220 VDD.n1618 VDD.n1116 1.81083
R24221 VDD.n3465 VDD.n3464 1.80928
R24222 VDD.n3467 VDD.n3464 1.77901
R24223 VDD.n1160 VDD.n1116 1.77901
R24224 VDD.n2206 VDD.t83 1.77879
R24225 VDD.t104 VDD.n831 1.77879
R24226 VDD.n3114 VDD.t92 1.77879
R24227 VDD.t90 VDD.n434 1.77879
R24228 VDD.n14 VDD.n6 1.4301
R24229 VDD.n14 VDD.n13 1.4301
R24230 VDD.n1080 VDD.t25 0.593262
R24231 VDD.n954 VDD.t73 0.593262
R24232 VDD.n2320 VDD.t95 0.593262
R24233 VDD.n2446 VDD.t17 0.593262
R24234 VDD.n682 VDD.t33 0.593262
R24235 VDD.n556 VDD.t78 0.593262
R24236 VDD.n3228 VDD.t91 0.593262
R24237 VDD.n3354 VDD.t21 0.593262
R24238 VDD.n1617 VDD.n1178 0.494402
R24239 VDD.n3659 VDD.n3658 0.471537
R24240 VDD.n116 VDD.n115 0.471537
R24241 VDD.n1393 VDD.n1337 0.471537
R24242 VDD.n1445 VDD.n1444 0.471537
R24243 VDD.n1633 VDD.n1159 0.457817
R24244 VDD.n3522 VDD.n261 0.305378
R24245 VDD.n278 VDD.n261 0.305378
R24246 VDD.n279 VDD.n278 0.305378
R24247 VDD.n280 VDD.n279 0.305378
R24248 VDD.n281 VDD.n280 0.305378
R24249 VDD.n282 VDD.n281 0.305378
R24250 VDD.n283 VDD.n282 0.305378
R24251 VDD.n284 VDD.n283 0.305378
R24252 VDD.n285 VDD.n284 0.305378
R24253 VDD.n286 VDD.n285 0.305378
R24254 VDD.n287 VDD.n286 0.305378
R24255 VDD.n289 VDD.n287 0.305378
R24256 VDD.n292 VDD.n289 0.305378
R24257 VDD.n294 VDD.n293 0.305378
R24258 VDD.n295 VDD.n294 0.305378
R24259 VDD.n296 VDD.n295 0.305378
R24260 VDD.n297 VDD.n296 0.305378
R24261 VDD.n298 VDD.n297 0.305378
R24262 VDD.n299 VDD.n298 0.305378
R24263 VDD.n300 VDD.n299 0.305378
R24264 VDD.n301 VDD.n300 0.305378
R24265 VDD.n302 VDD.n301 0.305378
R24266 VDD.n303 VDD.n302 0.305378
R24267 VDD.n3471 VDD.n303 0.305378
R24268 VDD.n3471 VDD.n3470 0.305378
R24269 VDD.n3470 VDD.n3469 0.305378
R24270 VDD.n1633 VDD.n1202 0.305378
R24271 VDD.n1639 VDD.n1202 0.305378
R24272 VDD.n1640 VDD.n1639 0.305378
R24273 VDD.n1641 VDD.n1640 0.305378
R24274 VDD.n1641 VDD.n1198 0.305378
R24275 VDD.n1647 VDD.n1198 0.305378
R24276 VDD.n1648 VDD.n1647 0.305378
R24277 VDD.n1649 VDD.n1648 0.305378
R24278 VDD.n1649 VDD.n1194 0.305378
R24279 VDD.n1655 VDD.n1194 0.305378
R24280 VDD.n1656 VDD.n1655 0.305378
R24281 VDD.n1657 VDD.n1656 0.305378
R24282 VDD.n1657 VDD.n1161 0.305378
R24283 VDD.n1694 VDD.n1162 0.305378
R24284 VDD.n1690 VDD.n1162 0.305378
R24285 VDD.n1690 VDD.n1689 0.305378
R24286 VDD.n1689 VDD.n1688 0.305378
R24287 VDD.n1688 VDD.n1168 0.305378
R24288 VDD.n1684 VDD.n1168 0.305378
R24289 VDD.n1684 VDD.n1683 0.305378
R24290 VDD.n1683 VDD.n1682 0.305378
R24291 VDD.n1682 VDD.n1173 0.305378
R24292 VDD.n1678 VDD.n1173 0.305378
R24293 VDD.n1678 VDD.n1677 0.305378
R24294 VDD.n1677 VDD.n1676 0.305378
R24295 VDD.n1676 VDD.n1178 0.305378
R24296 VDD.n3525 VDD.n3524 0.293183
R24297 VDD.n1629 VDD.n1159 0.293183
R24298 VDD.n3523 VDD.n3522 0.232207
R24299 VDD.n3469 VDD.n3467 0.232207
R24300 VDD.n3465 VDD.n253 0.192573
R24301 VDD.n1619 VDD.n1618 0.192573
R24302 VDD.n3532 VDD.n253 0.152939
R24303 VDD.n3533 VDD.n3532 0.152939
R24304 VDD.n3534 VDD.n3533 0.152939
R24305 VDD.n3534 VDD.n241 0.152939
R24306 VDD.n3548 VDD.n241 0.152939
R24307 VDD.n3549 VDD.n3548 0.152939
R24308 VDD.n3550 VDD.n3549 0.152939
R24309 VDD.n3550 VDD.n229 0.152939
R24310 VDD.n3564 VDD.n229 0.152939
R24311 VDD.n3565 VDD.n3564 0.152939
R24312 VDD.n3566 VDD.n3565 0.152939
R24313 VDD.n3566 VDD.n217 0.152939
R24314 VDD.n3580 VDD.n217 0.152939
R24315 VDD.n3581 VDD.n3580 0.152939
R24316 VDD.n3582 VDD.n3581 0.152939
R24317 VDD.n3583 VDD.n3582 0.152939
R24318 VDD.n3583 VDD.n205 0.152939
R24319 VDD.n3599 VDD.n205 0.152939
R24320 VDD.n3600 VDD.n3599 0.152939
R24321 VDD.n3601 VDD.n3600 0.152939
R24322 VDD.n3603 VDD.n3601 0.152939
R24323 VDD.n3603 VDD.n3602 0.152939
R24324 VDD.n3602 VDD.n194 0.152939
R24325 VDD.n194 VDD.n192 0.152939
R24326 VDD.n3623 VDD.n192 0.152939
R24327 VDD.n3624 VDD.n3623 0.152939
R24328 VDD.n3625 VDD.n3624 0.152939
R24329 VDD.n3625 VDD.n190 0.152939
R24330 VDD.n3630 VDD.n190 0.152939
R24331 VDD.n3631 VDD.n3630 0.152939
R24332 VDD.n3632 VDD.n3631 0.152939
R24333 VDD.n3632 VDD.n188 0.152939
R24334 VDD.n3637 VDD.n188 0.152939
R24335 VDD.n3638 VDD.n3637 0.152939
R24336 VDD.n3639 VDD.n3638 0.152939
R24337 VDD.n3639 VDD.n186 0.152939
R24338 VDD.n3644 VDD.n186 0.152939
R24339 VDD.n3645 VDD.n3644 0.152939
R24340 VDD.n3646 VDD.n3645 0.152939
R24341 VDD.n3646 VDD.n184 0.152939
R24342 VDD.n3651 VDD.n184 0.152939
R24343 VDD.n3652 VDD.n3651 0.152939
R24344 VDD.n3653 VDD.n3652 0.152939
R24345 VDD.n3653 VDD.n182 0.152939
R24346 VDD.n3658 VDD.n182 0.152939
R24347 VDD.n122 VDD.n116 0.152939
R24348 VDD.n123 VDD.n122 0.152939
R24349 VDD.n124 VDD.n123 0.152939
R24350 VDD.n124 VDD.n113 0.152939
R24351 VDD.n132 VDD.n113 0.152939
R24352 VDD.n133 VDD.n132 0.152939
R24353 VDD.n134 VDD.n133 0.152939
R24354 VDD.n134 VDD.n111 0.152939
R24355 VDD.n142 VDD.n111 0.152939
R24356 VDD.n143 VDD.n142 0.152939
R24357 VDD.n144 VDD.n143 0.152939
R24358 VDD.n144 VDD.n106 0.152939
R24359 VDD.n151 VDD.n106 0.152939
R24360 VDD.n152 VDD.n151 0.152939
R24361 VDD.n153 VDD.n152 0.152939
R24362 VDD.n153 VDD.n104 0.152939
R24363 VDD.n161 VDD.n104 0.152939
R24364 VDD.n162 VDD.n161 0.152939
R24365 VDD.n163 VDD.n162 0.152939
R24366 VDD.n163 VDD.n102 0.152939
R24367 VDD.n171 VDD.n102 0.152939
R24368 VDD.n172 VDD.n171 0.152939
R24369 VDD.n173 VDD.n172 0.152939
R24370 VDD.n173 VDD.n100 0.152939
R24371 VDD.n180 VDD.n100 0.152939
R24372 VDD.n181 VDD.n180 0.152939
R24373 VDD.n3659 VDD.n181 0.152939
R24374 VDD.n3709 VDD.n20 0.152939
R24375 VDD.n31 VDD.n20 0.152939
R24376 VDD.n32 VDD.n31 0.152939
R24377 VDD.n33 VDD.n32 0.152939
R24378 VDD.n34 VDD.n33 0.152939
R24379 VDD.n42 VDD.n34 0.152939
R24380 VDD.n43 VDD.n42 0.152939
R24381 VDD.n44 VDD.n43 0.152939
R24382 VDD.n45 VDD.n44 0.152939
R24383 VDD.n53 VDD.n45 0.152939
R24384 VDD.n54 VDD.n53 0.152939
R24385 VDD.n55 VDD.n54 0.152939
R24386 VDD.n56 VDD.n55 0.152939
R24387 VDD.n64 VDD.n56 0.152939
R24388 VDD.n65 VDD.n64 0.152939
R24389 VDD.n66 VDD.n65 0.152939
R24390 VDD.n67 VDD.n66 0.152939
R24391 VDD.n75 VDD.n67 0.152939
R24392 VDD.n76 VDD.n75 0.152939
R24393 VDD.n77 VDD.n76 0.152939
R24394 VDD.n78 VDD.n77 0.152939
R24395 VDD.n115 VDD.n78 0.152939
R24396 VDD.n3526 VDD.n3525 0.152939
R24397 VDD.n3526 VDD.n247 0.152939
R24398 VDD.n3540 VDD.n247 0.152939
R24399 VDD.n3541 VDD.n3540 0.152939
R24400 VDD.n3542 VDD.n3541 0.152939
R24401 VDD.n3542 VDD.n235 0.152939
R24402 VDD.n3556 VDD.n235 0.152939
R24403 VDD.n3557 VDD.n3556 0.152939
R24404 VDD.n3558 VDD.n3557 0.152939
R24405 VDD.n3558 VDD.n223 0.152939
R24406 VDD.n3572 VDD.n223 0.152939
R24407 VDD.n3573 VDD.n3572 0.152939
R24408 VDD.n3574 VDD.n3573 0.152939
R24409 VDD.n3574 VDD.n211 0.152939
R24410 VDD.n3590 VDD.n211 0.152939
R24411 VDD.n3591 VDD.n3590 0.152939
R24412 VDD.n3592 VDD.n3591 0.152939
R24413 VDD.n3592 VDD.n199 0.152939
R24414 VDD.n3611 VDD.n199 0.152939
R24415 VDD.n3612 VDD.n3611 0.152939
R24416 VDD.n3613 VDD.n3612 0.152939
R24417 VDD.n3613 VDD.n19 0.152939
R24418 VDD.n292 VDD.n259 0.152939
R24419 VDD.n293 VDD.n259 0.152939
R24420 VDD.n1542 VDD.n1541 0.152939
R24421 VDD.n1543 VDD.n1542 0.152939
R24422 VDD.n1543 VDD.n1255 0.152939
R24423 VDD.n1557 VDD.n1255 0.152939
R24424 VDD.n1558 VDD.n1557 0.152939
R24425 VDD.n1559 VDD.n1558 0.152939
R24426 VDD.n1559 VDD.n1243 0.152939
R24427 VDD.n1573 VDD.n1243 0.152939
R24428 VDD.n1574 VDD.n1573 0.152939
R24429 VDD.n1575 VDD.n1574 0.152939
R24430 VDD.n1575 VDD.n1231 0.152939
R24431 VDD.n1589 VDD.n1231 0.152939
R24432 VDD.n1590 VDD.n1589 0.152939
R24433 VDD.n1591 VDD.n1590 0.152939
R24434 VDD.n1591 VDD.n1218 0.152939
R24435 VDD.n1606 VDD.n1218 0.152939
R24436 VDD.n1607 VDD.n1606 0.152939
R24437 VDD.n1608 VDD.n1607 0.152939
R24438 VDD.n1608 VDD.n1205 0.152939
R24439 VDD.n1627 VDD.n1205 0.152939
R24440 VDD.n1628 VDD.n1627 0.152939
R24441 VDD.n1629 VDD.n1628 0.152939
R24442 VDD.n1695 VDD.n1161 0.152939
R24443 VDD.n1695 VDD.n1694 0.152939
R24444 VDD.n1452 VDD.n1337 0.152939
R24445 VDD.n1453 VDD.n1452 0.152939
R24446 VDD.n1454 VDD.n1453 0.152939
R24447 VDD.n1454 VDD.n1325 0.152939
R24448 VDD.n1468 VDD.n1325 0.152939
R24449 VDD.n1469 VDD.n1468 0.152939
R24450 VDD.n1470 VDD.n1469 0.152939
R24451 VDD.n1470 VDD.n1313 0.152939
R24452 VDD.n1484 VDD.n1313 0.152939
R24453 VDD.n1485 VDD.n1484 0.152939
R24454 VDD.n1486 VDD.n1485 0.152939
R24455 VDD.n1486 VDD.n1301 0.152939
R24456 VDD.n1500 VDD.n1301 0.152939
R24457 VDD.n1501 VDD.n1500 0.152939
R24458 VDD.n1502 VDD.n1501 0.152939
R24459 VDD.n1502 VDD.n1289 0.152939
R24460 VDD.n1516 VDD.n1289 0.152939
R24461 VDD.n1517 VDD.n1516 0.152939
R24462 VDD.n1518 VDD.n1517 0.152939
R24463 VDD.n1518 VDD.n1277 0.152939
R24464 VDD.n1533 VDD.n1277 0.152939
R24465 VDD.n1534 VDD.n1533 0.152939
R24466 VDD.n1535 VDD.n1534 0.152939
R24467 VDD.n1535 VDD.n1261 0.152939
R24468 VDD.n1549 VDD.n1261 0.152939
R24469 VDD.n1550 VDD.n1549 0.152939
R24470 VDD.n1551 VDD.n1550 0.152939
R24471 VDD.n1551 VDD.n1249 0.152939
R24472 VDD.n1565 VDD.n1249 0.152939
R24473 VDD.n1566 VDD.n1565 0.152939
R24474 VDD.n1567 VDD.n1566 0.152939
R24475 VDD.n1567 VDD.n1237 0.152939
R24476 VDD.n1581 VDD.n1237 0.152939
R24477 VDD.n1582 VDD.n1581 0.152939
R24478 VDD.n1583 VDD.n1582 0.152939
R24479 VDD.n1583 VDD.n1225 0.152939
R24480 VDD.n1597 VDD.n1225 0.152939
R24481 VDD.n1598 VDD.n1597 0.152939
R24482 VDD.n1600 VDD.n1598 0.152939
R24483 VDD.n1600 VDD.n1599 0.152939
R24484 VDD.n1599 VDD.n1212 0.152939
R24485 VDD.n1615 VDD.n1212 0.152939
R24486 VDD.n1616 VDD.n1615 0.152939
R24487 VDD.n1620 VDD.n1616 0.152939
R24488 VDD.n1620 VDD.n1619 0.152939
R24489 VDD.n1444 VDD.n1343 0.152939
R24490 VDD.n1437 VDD.n1343 0.152939
R24491 VDD.n1437 VDD.n1436 0.152939
R24492 VDD.n1436 VDD.n1435 0.152939
R24493 VDD.n1435 VDD.n1361 0.152939
R24494 VDD.n1431 VDD.n1361 0.152939
R24495 VDD.n1431 VDD.n1430 0.152939
R24496 VDD.n1430 VDD.n1429 0.152939
R24497 VDD.n1429 VDD.n1367 0.152939
R24498 VDD.n1425 VDD.n1367 0.152939
R24499 VDD.n1425 VDD.n1424 0.152939
R24500 VDD.n1424 VDD.n1423 0.152939
R24501 VDD.n1423 VDD.n1373 0.152939
R24502 VDD.n1415 VDD.n1373 0.152939
R24503 VDD.n1415 VDD.n1414 0.152939
R24504 VDD.n1414 VDD.n1413 0.152939
R24505 VDD.n1413 VDD.n1377 0.152939
R24506 VDD.n1409 VDD.n1377 0.152939
R24507 VDD.n1409 VDD.n1408 0.152939
R24508 VDD.n1408 VDD.n1407 0.152939
R24509 VDD.n1407 VDD.n1383 0.152939
R24510 VDD.n1403 VDD.n1383 0.152939
R24511 VDD.n1403 VDD.n1402 0.152939
R24512 VDD.n1402 VDD.n1401 0.152939
R24513 VDD.n1401 VDD.n1389 0.152939
R24514 VDD.n1394 VDD.n1389 0.152939
R24515 VDD.n1394 VDD.n1393 0.152939
R24516 VDD.n1446 VDD.n1445 0.152939
R24517 VDD.n1446 VDD.n1331 0.152939
R24518 VDD.n1460 VDD.n1331 0.152939
R24519 VDD.n1461 VDD.n1460 0.152939
R24520 VDD.n1462 VDD.n1461 0.152939
R24521 VDD.n1462 VDD.n1319 0.152939
R24522 VDD.n1476 VDD.n1319 0.152939
R24523 VDD.n1477 VDD.n1476 0.152939
R24524 VDD.n1478 VDD.n1477 0.152939
R24525 VDD.n1478 VDD.n1307 0.152939
R24526 VDD.n1492 VDD.n1307 0.152939
R24527 VDD.n1493 VDD.n1492 0.152939
R24528 VDD.n1494 VDD.n1493 0.152939
R24529 VDD.n1494 VDD.n1295 0.152939
R24530 VDD.n1508 VDD.n1295 0.152939
R24531 VDD.n1509 VDD.n1508 0.152939
R24532 VDD.n1510 VDD.n1509 0.152939
R24533 VDD.n1510 VDD.n1283 0.152939
R24534 VDD.n1524 VDD.n1283 0.152939
R24535 VDD.n1525 VDD.n1524 0.152939
R24536 VDD.n1527 VDD.n1525 0.152939
R24537 VDD.n1527 VDD.n1526 0.152939
R24538 VDD.n3710 VDD.n3709 0.0695946
R24539 VDD.n3710 VDD.n19 0.0695946
R24540 VDD.n1541 VDD.n1271 0.0695946
R24541 VDD.n1526 VDD.n1271 0.0695946
R24542 VDD.n3466 VDD.n3465 0.0645244
R24543 VDD.n1618 VDD.n1617 0.0645244
R24544 VDD.n1617 VDD.n1160 0.0158509
R24545 VDD.n3467 VDD.n3466 0.0151199
R24546 VDD VDD.n15 0.00833333
R24547 VDD.n1696 VDD.n1159 0.0070625
R24548 VDD.n3524 VDD.n3523 0.00675
R24549 VP.n208 VP.n207 161.3
R24550 VP.n206 VP.n106 161.3
R24551 VP.n205 VP.n204 161.3
R24552 VP.n203 VP.n107 161.3
R24553 VP.n202 VP.n201 161.3
R24554 VP.n200 VP.n108 161.3
R24555 VP.n199 VP.n198 161.3
R24556 VP.n197 VP.n109 161.3
R24557 VP.n196 VP.n195 161.3
R24558 VP.n194 VP.n110 161.3
R24559 VP.n193 VP.n192 161.3
R24560 VP.n191 VP.n111 161.3
R24561 VP.n190 VP.n189 161.3
R24562 VP.n188 VP.n112 161.3
R24563 VP.n187 VP.n186 161.3
R24564 VP.n185 VP.n114 161.3
R24565 VP.n184 VP.n183 161.3
R24566 VP.n182 VP.n115 161.3
R24567 VP.n181 VP.n180 161.3
R24568 VP.n179 VP.n116 161.3
R24569 VP.n178 VP.n177 161.3
R24570 VP.n176 VP.n117 161.3
R24571 VP.n175 VP.n174 161.3
R24572 VP.n173 VP.n118 161.3
R24573 VP.n172 VP.n171 161.3
R24574 VP.n170 VP.n119 161.3
R24575 VP.n169 VP.n168 161.3
R24576 VP.n167 VP.n121 161.3
R24577 VP.n166 VP.n165 161.3
R24578 VP.n164 VP.n122 161.3
R24579 VP.n163 VP.n162 161.3
R24580 VP.n161 VP.n123 161.3
R24581 VP.n160 VP.n159 161.3
R24582 VP.n158 VP.n124 161.3
R24583 VP.n157 VP.n156 161.3
R24584 VP.n155 VP.n125 161.3
R24585 VP.n154 VP.n153 161.3
R24586 VP.n151 VP.n126 161.3
R24587 VP.n150 VP.n149 161.3
R24588 VP.n148 VP.n127 161.3
R24589 VP.n147 VP.n146 161.3
R24590 VP.n145 VP.n128 161.3
R24591 VP.n144 VP.n143 161.3
R24592 VP.n142 VP.n129 161.3
R24593 VP.n141 VP.n140 161.3
R24594 VP.n139 VP.n130 161.3
R24595 VP.n138 VP.n137 161.3
R24596 VP.n136 VP.n131 161.3
R24597 VP.n135 VP.n134 161.3
R24598 VP.n103 VP.n102 161.3
R24599 VP.n101 VP.n1 161.3
R24600 VP.n100 VP.n99 161.3
R24601 VP.n98 VP.n2 161.3
R24602 VP.n97 VP.n96 161.3
R24603 VP.n95 VP.n3 161.3
R24604 VP.n94 VP.n93 161.3
R24605 VP.n92 VP.n4 161.3
R24606 VP.n91 VP.n90 161.3
R24607 VP.n89 VP.n5 161.3
R24608 VP.n88 VP.n87 161.3
R24609 VP.n86 VP.n6 161.3
R24610 VP.n85 VP.n84 161.3
R24611 VP.n82 VP.n7 161.3
R24612 VP.n81 VP.n80 161.3
R24613 VP.n79 VP.n8 161.3
R24614 VP.n78 VP.n77 161.3
R24615 VP.n76 VP.n9 161.3
R24616 VP.n75 VP.n74 161.3
R24617 VP.n73 VP.n10 161.3
R24618 VP.n72 VP.n71 161.3
R24619 VP.n70 VP.n11 161.3
R24620 VP.n69 VP.n68 161.3
R24621 VP.n67 VP.n12 161.3
R24622 VP.n66 VP.n65 161.3
R24623 VP.n63 VP.n13 161.3
R24624 VP.n62 VP.n61 161.3
R24625 VP.n60 VP.n14 161.3
R24626 VP.n59 VP.n58 161.3
R24627 VP.n57 VP.n15 161.3
R24628 VP.n56 VP.n55 161.3
R24629 VP.n54 VP.n16 161.3
R24630 VP.n53 VP.n52 161.3
R24631 VP.n51 VP.n17 161.3
R24632 VP.n50 VP.n49 161.3
R24633 VP.n48 VP.n18 161.3
R24634 VP.n47 VP.n46 161.3
R24635 VP.n44 VP.n19 161.3
R24636 VP.n43 VP.n42 161.3
R24637 VP.n41 VP.n20 161.3
R24638 VP.n40 VP.n39 161.3
R24639 VP.n38 VP.n21 161.3
R24640 VP.n37 VP.n36 161.3
R24641 VP.n35 VP.n22 161.3
R24642 VP.n34 VP.n33 161.3
R24643 VP.n32 VP.n23 161.3
R24644 VP.n31 VP.n30 161.3
R24645 VP.n29 VP.n24 161.3
R24646 VP.n28 VP.n27 161.3
R24647 VP.n200 VP.n199 72.0595
R24648 VP.n95 VP.n94 72.0595
R24649 VP.n133 VP.n132 70.3045
R24650 VP.n26 VP.n25 70.3045
R24651 VP.n209 VP.n105 69.0311
R24652 VP.n104 VP.n0 69.0311
R24653 VP.n144 VP.n129 64.2894
R24654 VP.n182 VP.n181 64.2894
R24655 VP.n37 VP.n22 64.2894
R24656 VP.n76 VP.n75 64.2894
R24657 VP.n210 VP.n209 57.2702
R24658 VP.n163 VP.n123 56.5193
R24659 VP.n164 VP.n163 56.5193
R24660 VP.n56 VP.n16 56.5193
R24661 VP.n57 VP.n56 56.5193
R24662 VP.n145 VP.n144 48.7492
R24663 VP.n181 VP.n116 48.7492
R24664 VP.n38 VP.n37 48.7492
R24665 VP.n75 VP.n10 48.7492
R24666 VP.n132 VP.t7 46.6433
R24667 VP.n25 VP.t8 46.6433
R24668 VP.n199 VP.n109 40.979
R24669 VP.n94 VP.n4 40.979
R24670 VP.n140 VP.n129 24.4675
R24671 VP.n140 VP.n139 24.4675
R24672 VP.n139 VP.n138 24.4675
R24673 VP.n138 VP.n131 24.4675
R24674 VP.n134 VP.n131 24.4675
R24675 VP.n159 VP.n123 24.4675
R24676 VP.n159 VP.n158 24.4675
R24677 VP.n158 VP.n157 24.4675
R24678 VP.n157 VP.n125 24.4675
R24679 VP.n153 VP.n125 24.4675
R24680 VP.n151 VP.n150 24.4675
R24681 VP.n150 VP.n127 24.4675
R24682 VP.n146 VP.n127 24.4675
R24683 VP.n146 VP.n145 24.4675
R24684 VP.n177 VP.n116 24.4675
R24685 VP.n177 VP.n176 24.4675
R24686 VP.n176 VP.n175 24.4675
R24687 VP.n175 VP.n118 24.4675
R24688 VP.n171 VP.n170 24.4675
R24689 VP.n170 VP.n169 24.4675
R24690 VP.n169 VP.n121 24.4675
R24691 VP.n165 VP.n121 24.4675
R24692 VP.n165 VP.n164 24.4675
R24693 VP.n195 VP.n109 24.4675
R24694 VP.n195 VP.n194 24.4675
R24695 VP.n194 VP.n193 24.4675
R24696 VP.n193 VP.n111 24.4675
R24697 VP.n189 VP.n188 24.4675
R24698 VP.n188 VP.n187 24.4675
R24699 VP.n187 VP.n114 24.4675
R24700 VP.n183 VP.n114 24.4675
R24701 VP.n183 VP.n182 24.4675
R24702 VP.n207 VP.n206 24.4675
R24703 VP.n206 VP.n205 24.4675
R24704 VP.n205 VP.n107 24.4675
R24705 VP.n201 VP.n107 24.4675
R24706 VP.n201 VP.n200 24.4675
R24707 VP.n27 VP.n24 24.4675
R24708 VP.n31 VP.n24 24.4675
R24709 VP.n32 VP.n31 24.4675
R24710 VP.n33 VP.n32 24.4675
R24711 VP.n33 VP.n22 24.4675
R24712 VP.n39 VP.n38 24.4675
R24713 VP.n39 VP.n20 24.4675
R24714 VP.n43 VP.n20 24.4675
R24715 VP.n44 VP.n43 24.4675
R24716 VP.n46 VP.n18 24.4675
R24717 VP.n50 VP.n18 24.4675
R24718 VP.n51 VP.n50 24.4675
R24719 VP.n52 VP.n51 24.4675
R24720 VP.n52 VP.n16 24.4675
R24721 VP.n58 VP.n57 24.4675
R24722 VP.n58 VP.n14 24.4675
R24723 VP.n62 VP.n14 24.4675
R24724 VP.n63 VP.n62 24.4675
R24725 VP.n65 VP.n63 24.4675
R24726 VP.n69 VP.n12 24.4675
R24727 VP.n70 VP.n69 24.4675
R24728 VP.n71 VP.n70 24.4675
R24729 VP.n71 VP.n10 24.4675
R24730 VP.n77 VP.n76 24.4675
R24731 VP.n77 VP.n8 24.4675
R24732 VP.n81 VP.n8 24.4675
R24733 VP.n82 VP.n81 24.4675
R24734 VP.n84 VP.n82 24.4675
R24735 VP.n88 VP.n6 24.4675
R24736 VP.n89 VP.n88 24.4675
R24737 VP.n90 VP.n89 24.4675
R24738 VP.n90 VP.n4 24.4675
R24739 VP.n96 VP.n95 24.4675
R24740 VP.n96 VP.n2 24.4675
R24741 VP.n100 VP.n2 24.4675
R24742 VP.n101 VP.n100 24.4675
R24743 VP.n102 VP.n101 24.4675
R24744 VP.n152 VP.n151 22.5101
R24745 VP.n120 VP.n118 22.5101
R24746 VP.n45 VP.n44 22.5101
R24747 VP.n64 VP.n12 22.5101
R24748 VP.n113 VP.n111 18.5954
R24749 VP.n83 VP.n6 18.5954
R24750 VP VP.n210 13.8377
R24751 VP.n210 VP.n104 13.3686
R24752 VP.n133 VP.t2 12.9398
R24753 VP.n152 VP.t1 12.9398
R24754 VP.n120 VP.t6 12.9398
R24755 VP.n113 VP.t9 12.9398
R24756 VP.n105 VP.t3 12.9398
R24757 VP.n26 VP.t0 12.9398
R24758 VP.n45 VP.t11 12.9398
R24759 VP.n64 VP.t10 12.9398
R24760 VP.n83 VP.t5 12.9398
R24761 VP.n0 VP.t4 12.9398
R24762 VP.n207 VP.n105 9.7873
R24763 VP.n102 VP.n0 9.7873
R24764 VP.n134 VP.n133 5.87258
R24765 VP.n189 VP.n113 5.87258
R24766 VP.n27 VP.n26 5.87258
R24767 VP.n84 VP.n83 5.87258
R24768 VP.n153 VP.n152 1.95786
R24769 VP.n171 VP.n120 1.95786
R24770 VP.n46 VP.n45 1.95786
R24771 VP.n65 VP.n64 1.95786
R24772 VP.n135 VP.n132 0.976621
R24773 VP.n28 VP.n25 0.976621
R24774 VP.n209 VP.n208 0.466196
R24775 VP.n104 VP.n103 0.466196
R24776 VP.n208 VP.n106 0.189894
R24777 VP.n204 VP.n106 0.189894
R24778 VP.n204 VP.n203 0.189894
R24779 VP.n203 VP.n202 0.189894
R24780 VP.n202 VP.n108 0.189894
R24781 VP.n198 VP.n108 0.189894
R24782 VP.n198 VP.n197 0.189894
R24783 VP.n197 VP.n196 0.189894
R24784 VP.n196 VP.n110 0.189894
R24785 VP.n192 VP.n110 0.189894
R24786 VP.n192 VP.n191 0.189894
R24787 VP.n191 VP.n190 0.189894
R24788 VP.n190 VP.n112 0.189894
R24789 VP.n186 VP.n112 0.189894
R24790 VP.n186 VP.n185 0.189894
R24791 VP.n185 VP.n184 0.189894
R24792 VP.n184 VP.n115 0.189894
R24793 VP.n180 VP.n115 0.189894
R24794 VP.n180 VP.n179 0.189894
R24795 VP.n179 VP.n178 0.189894
R24796 VP.n178 VP.n117 0.189894
R24797 VP.n174 VP.n117 0.189894
R24798 VP.n174 VP.n173 0.189894
R24799 VP.n173 VP.n172 0.189894
R24800 VP.n172 VP.n119 0.189894
R24801 VP.n168 VP.n119 0.189894
R24802 VP.n168 VP.n167 0.189894
R24803 VP.n167 VP.n166 0.189894
R24804 VP.n166 VP.n122 0.189894
R24805 VP.n162 VP.n122 0.189894
R24806 VP.n162 VP.n161 0.189894
R24807 VP.n161 VP.n160 0.189894
R24808 VP.n160 VP.n124 0.189894
R24809 VP.n156 VP.n124 0.189894
R24810 VP.n156 VP.n155 0.189894
R24811 VP.n155 VP.n154 0.189894
R24812 VP.n154 VP.n126 0.189894
R24813 VP.n149 VP.n126 0.189894
R24814 VP.n149 VP.n148 0.189894
R24815 VP.n148 VP.n147 0.189894
R24816 VP.n147 VP.n128 0.189894
R24817 VP.n143 VP.n128 0.189894
R24818 VP.n143 VP.n142 0.189894
R24819 VP.n142 VP.n141 0.189894
R24820 VP.n141 VP.n130 0.189894
R24821 VP.n137 VP.n130 0.189894
R24822 VP.n137 VP.n136 0.189894
R24823 VP.n136 VP.n135 0.189894
R24824 VP.n29 VP.n28 0.189894
R24825 VP.n30 VP.n29 0.189894
R24826 VP.n30 VP.n23 0.189894
R24827 VP.n34 VP.n23 0.189894
R24828 VP.n35 VP.n34 0.189894
R24829 VP.n36 VP.n35 0.189894
R24830 VP.n36 VP.n21 0.189894
R24831 VP.n40 VP.n21 0.189894
R24832 VP.n41 VP.n40 0.189894
R24833 VP.n42 VP.n41 0.189894
R24834 VP.n42 VP.n19 0.189894
R24835 VP.n47 VP.n19 0.189894
R24836 VP.n48 VP.n47 0.189894
R24837 VP.n49 VP.n48 0.189894
R24838 VP.n49 VP.n17 0.189894
R24839 VP.n53 VP.n17 0.189894
R24840 VP.n54 VP.n53 0.189894
R24841 VP.n55 VP.n54 0.189894
R24842 VP.n55 VP.n15 0.189894
R24843 VP.n59 VP.n15 0.189894
R24844 VP.n60 VP.n59 0.189894
R24845 VP.n61 VP.n60 0.189894
R24846 VP.n61 VP.n13 0.189894
R24847 VP.n66 VP.n13 0.189894
R24848 VP.n67 VP.n66 0.189894
R24849 VP.n68 VP.n67 0.189894
R24850 VP.n68 VP.n11 0.189894
R24851 VP.n72 VP.n11 0.189894
R24852 VP.n73 VP.n72 0.189894
R24853 VP.n74 VP.n73 0.189894
R24854 VP.n74 VP.n9 0.189894
R24855 VP.n78 VP.n9 0.189894
R24856 VP.n79 VP.n78 0.189894
R24857 VP.n80 VP.n79 0.189894
R24858 VP.n80 VP.n7 0.189894
R24859 VP.n85 VP.n7 0.189894
R24860 VP.n86 VP.n85 0.189894
R24861 VP.n87 VP.n86 0.189894
R24862 VP.n87 VP.n5 0.189894
R24863 VP.n91 VP.n5 0.189894
R24864 VP.n92 VP.n91 0.189894
R24865 VP.n93 VP.n92 0.189894
R24866 VP.n93 VP.n3 0.189894
R24867 VP.n97 VP.n3 0.189894
R24868 VP.n98 VP.n97 0.189894
R24869 VP.n99 VP.n98 0.189894
R24870 VP.n99 VP.n1 0.189894
R24871 VP.n103 VP.n1 0.189894
R24872 VOUT.n8 VOUT.n6 115.419
R24873 VOUT.n2 VOUT.n0 115.419
R24874 VOUT.n2 VOUT.n1 114.382
R24875 VOUT.n8 VOUT.n7 114.382
R24876 VOUT.n30 VOUT.t7 107.871
R24877 VOUT.n25 VOUT.t6 107.871
R24878 VOUT.n20 VOUT.t5 107.871
R24879 VOUT.n15 VOUT.t32 107.871
R24880 VOUT.n11 VOUT.t24 107.871
R24881 VOUT.n57 VOUT.t11 106.037
R24882 VOUT.n52 VOUT.t8 106.037
R24883 VOUT.n47 VOUT.t9 106.037
R24884 VOUT.n42 VOUT.t39 106.037
R24885 VOUT.n38 VOUT.t50 106.037
R24886 VOUT.n56 VOUT.n54 88.8325
R24887 VOUT.n51 VOUT.n49 88.8325
R24888 VOUT.n46 VOUT.n44 88.8325
R24889 VOUT.n41 VOUT.n39 88.8325
R24890 VOUT.n37 VOUT.n35 88.8325
R24891 VOUT.n32 VOUT.n31 86.9991
R24892 VOUT.n30 VOUT.n29 86.9991
R24893 VOUT.n27 VOUT.n26 86.9991
R24894 VOUT.n25 VOUT.n24 86.9991
R24895 VOUT.n22 VOUT.n21 86.9991
R24896 VOUT.n20 VOUT.n19 86.9991
R24897 VOUT.n17 VOUT.n16 86.9991
R24898 VOUT.n15 VOUT.n14 86.9991
R24899 VOUT.n13 VOUT.n12 86.9991
R24900 VOUT.n11 VOUT.n10 86.9991
R24901 VOUT.n56 VOUT.n55 86.9991
R24902 VOUT.n51 VOUT.n50 86.9991
R24903 VOUT.n46 VOUT.n45 86.9991
R24904 VOUT.n41 VOUT.n40 86.9991
R24905 VOUT.n37 VOUT.n36 86.9991
R24906 VOUT.n31 VOUT.t23 19.039
R24907 VOUT.n31 VOUT.t29 19.039
R24908 VOUT.n29 VOUT.t38 19.039
R24909 VOUT.n29 VOUT.t48 19.039
R24910 VOUT.n26 VOUT.t22 19.039
R24911 VOUT.n26 VOUT.t28 19.039
R24912 VOUT.n24 VOUT.t36 19.039
R24913 VOUT.n24 VOUT.t45 19.039
R24914 VOUT.n21 VOUT.t21 19.039
R24915 VOUT.n21 VOUT.t27 19.039
R24916 VOUT.n19 VOUT.t35 19.039
R24917 VOUT.n19 VOUT.t44 19.039
R24918 VOUT.n16 VOUT.t13 19.039
R24919 VOUT.n16 VOUT.t25 19.039
R24920 VOUT.n14 VOUT.t26 19.039
R24921 VOUT.n14 VOUT.t42 19.039
R24922 VOUT.n12 VOUT.t30 19.039
R24923 VOUT.n12 VOUT.t12 19.039
R24924 VOUT.n10 VOUT.t31 19.039
R24925 VOUT.n10 VOUT.t16 19.039
R24926 VOUT.n54 VOUT.t46 19.039
R24927 VOUT.n54 VOUT.t37 19.039
R24928 VOUT.n55 VOUT.t17 19.039
R24929 VOUT.n55 VOUT.t53 19.039
R24930 VOUT.n49 VOUT.t47 19.039
R24931 VOUT.n49 VOUT.t33 19.039
R24932 VOUT.n50 VOUT.t15 19.039
R24933 VOUT.n50 VOUT.t54 19.039
R24934 VOUT.n44 VOUT.t43 19.039
R24935 VOUT.n44 VOUT.t34 19.039
R24936 VOUT.n45 VOUT.t14 19.039
R24937 VOUT.n45 VOUT.t52 19.039
R24938 VOUT.n39 VOUT.t18 19.039
R24939 VOUT.n39 VOUT.t49 19.039
R24940 VOUT.n40 VOUT.t10 19.039
R24941 VOUT.n40 VOUT.t40 19.039
R24942 VOUT.n35 VOUT.t41 19.039
R24943 VOUT.n35 VOUT.t19 19.039
R24944 VOUT.n36 VOUT.t51 19.039
R24945 VOUT.n36 VOUT.t20 19.039
R24946 VOUT.n7 VOUT.t3 17.1535
R24947 VOUT.n7 VOUT.t56 17.1535
R24948 VOUT.n6 VOUT.t0 17.1535
R24949 VOUT.n6 VOUT.t4 17.1535
R24950 VOUT.n1 VOUT.t57 17.1535
R24951 VOUT.n1 VOUT.t1 17.1535
R24952 VOUT.n0 VOUT.t2 17.1535
R24953 VOUT.n0 VOUT.t55 17.1535
R24954 VOUT.n34 VOUT.n9 8.51908
R24955 VOUT.n18 VOUT.n13 6.51846
R24956 VOUT.n59 VOUT.n34 5.75299
R24957 VOUT.n33 VOUT.n32 5.72751
R24958 VOUT.n28 VOUT.n27 5.72751
R24959 VOUT.n23 VOUT.n22 5.72751
R24960 VOUT.n18 VOUT.n17 5.72751
R24961 VOUT.n9 VOUT.n3 5.61637
R24962 VOUT.n43 VOUT.n38 5.60179
R24963 VOUT.n9 VOUT.n8 4.91768
R24964 VOUT.n3 VOUT.n2 4.91768
R24965 VOUT.n58 VOUT.n57 4.81084
R24966 VOUT.n53 VOUT.n52 4.81084
R24967 VOUT.n48 VOUT.n47 4.81084
R24968 VOUT.n43 VOUT.n42 4.81084
R24969 VOUT.n60 VOUT.n3 4.76136
R24970 VOUT.n5 VOUT 4.5219
R24971 VOUT.n34 VOUT.n33 4.24958
R24972 VOUT.n59 VOUT.n58 4.24958
R24973 VOUT.n60 VOUT.n59 3.73872
R24974 VOUT.n32 VOUT.n30 1.83383
R24975 VOUT.n27 VOUT.n25 1.83383
R24976 VOUT.n22 VOUT.n20 1.83383
R24977 VOUT.n17 VOUT.n15 1.83383
R24978 VOUT.n13 VOUT.n11 1.83383
R24979 VOUT.n57 VOUT.n56 1.83383
R24980 VOUT.n52 VOUT.n51 1.83383
R24981 VOUT.n47 VOUT.n46 1.83383
R24982 VOUT.n42 VOUT.n41 1.83383
R24983 VOUT.n38 VOUT.n37 1.83383
R24984 VOUT.n33 VOUT.n28 0.791448
R24985 VOUT.n28 VOUT.n23 0.791448
R24986 VOUT.n23 VOUT.n18 0.791448
R24987 VOUT.n58 VOUT.n53 0.791448
R24988 VOUT.n53 VOUT.n48 0.791448
R24989 VOUT.n48 VOUT.n43 0.791448
R24990 VOUT.n60 VOUT.n5 0.44324
R24991 VOUT.n5 VOUT.n4 0.420369
R24992 VOUT.n4 VOUT.t58 0.122428
R24993 VOUT VOUT.n60 0.0099
R24994 VOUT.n4 VOUT.t59 0.00976471
R24995 a_n7386_8166.n1 a_n7386_8166.t2 180.57
R24996 a_n7386_8166.n2 a_n7386_8166.t9 180.57
R24997 a_n7386_8166.n4 a_n7386_8166.t0 180.57
R24998 a_n7386_8166.n1 a_n7386_8166.t4 178.721
R24999 a_n7386_8166.n2 a_n7386_8166.t10 178.721
R25000 a_n7386_8166.n2 a_n7386_8166.t8 178.721
R25001 a_n7386_8166.n3 a_n7386_8166.t12 178.721
R25002 a_n7386_8166.n4 a_n7386_8166.t3 178.721
R25003 a_n7386_8166.n1 a_n7386_8166.n8 147.466
R25004 a_n7386_8166.n2 a_n7386_8166.n6 147.466
R25005 a_n7386_8166.n3 a_n7386_8166.n7 147.466
R25006 a_n7386_8166.n4 a_n7386_8166.n5 147.466
R25007 a_n7386_8166.n8 a_n7386_8166.t14 31.2553
R25008 a_n7386_8166.n8 a_n7386_8166.t15 31.2553
R25009 a_n7386_8166.n6 a_n7386_8166.t11 31.2553
R25010 a_n7386_8166.n6 a_n7386_8166.t6 31.2553
R25011 a_n7386_8166.n7 a_n7386_8166.t7 31.2553
R25012 a_n7386_8166.n7 a_n7386_8166.t5 31.2553
R25013 a_n7386_8166.n5 a_n7386_8166.t1 31.2553
R25014 a_n7386_8166.n5 a_n7386_8166.t13 31.2553
R25015 a_n7386_8166.n0 a_n7386_8166.n4 28.6915
R25016 a_n7386_8166.t16 a_n7386_8166.n0 11.0065
R25017 a_n7386_8166.n0 a_n7386_8166.n1 10.7713
R25018 a_n7386_8166.n0 a_n7386_8166.n3 9.10512
R25019 a_n7386_8166.n3 a_n7386_8166.n2 5.98829
R25020 a_n17362_8608.n20 a_n17362_8608.n2 168.903
R25021 a_n17362_8608.n5 a_n17362_8608.n3 168.903
R25022 a_n17362_8608.n5 a_n17362_8608.n4 167.054
R25023 a_n17362_8608.n21 a_n17362_8608.n20 167.054
R25024 a_n17362_8608.n1 a_n17362_8608.n6 79.8686
R25025 a_n17362_8608.n11 a_n17362_8608.n10 79.8684
R25026 a_n17362_8608.n11 a_n17362_8608.n8 79.8684
R25027 a_n17362_8608.n1 a_n17362_8608.n12 78.1215
R25028 a_n17362_8608.n1 a_n17362_8608.n7 78.1215
R25029 a_n17362_8608.n11 a_n17362_8608.n9 78.1213
R25030 a_n17362_8608.n14 a_n17362_8608.t27 56.79
R25031 a_n17362_8608.n13 a_n17362_8608.t22 56.79
R25032 a_n17362_8608.n17 a_n17362_8608.t23 56.7896
R25033 a_n17362_8608.n16 a_n17362_8608.t20 56.7896
R25034 a_n17362_8608.n17 a_n17362_8608.t24 55.1548
R25035 a_n17362_8608.n16 a_n17362_8608.t26 55.1548
R25036 a_n17362_8608.n14 a_n17362_8608.t21 55.1548
R25037 a_n17362_8608.n13 a_n17362_8608.t25 55.1548
R25038 a_n17362_8608.n1 a_n17362_8608.n11 36.6551
R25039 a_n17362_8608.n19 a_n17362_8608.n5 35.2333
R25040 a_n17362_8608.n2 a_n17362_8608.t14 31.2553
R25041 a_n17362_8608.n2 a_n17362_8608.t11 31.2553
R25042 a_n17362_8608.n3 a_n17362_8608.t15 31.2553
R25043 a_n17362_8608.n3 a_n17362_8608.t17 31.2553
R25044 a_n17362_8608.n4 a_n17362_8608.t13 31.2553
R25045 a_n17362_8608.n4 a_n17362_8608.t12 31.2553
R25046 a_n17362_8608.n21 a_n17362_8608.t16 31.2553
R25047 a_n17362_8608.t18 a_n17362_8608.n21 31.2553
R25048 a_n17362_8608.n20 a_n17362_8608.n19 23.6288
R25049 a_n17362_8608.n0 a_n17362_8608.n1 14.1734
R25050 a_n17362_8608.n12 a_n17362_8608.t7 13.6087
R25051 a_n17362_8608.n12 a_n17362_8608.t10 13.6087
R25052 a_n17362_8608.n7 a_n17362_8608.t0 13.6087
R25053 a_n17362_8608.n7 a_n17362_8608.t19 13.6087
R25054 a_n17362_8608.n6 a_n17362_8608.t4 13.6087
R25055 a_n17362_8608.n6 a_n17362_8608.t2 13.6087
R25056 a_n17362_8608.n10 a_n17362_8608.t3 13.6087
R25057 a_n17362_8608.n10 a_n17362_8608.t6 13.6087
R25058 a_n17362_8608.n9 a_n17362_8608.t5 13.6087
R25059 a_n17362_8608.n9 a_n17362_8608.t1 13.6087
R25060 a_n17362_8608.n8 a_n17362_8608.t9 13.6087
R25061 a_n17362_8608.n8 a_n17362_8608.t8 13.6087
R25062 a_n17362_8608.n19 a_n17362_8608.n0 11.4887
R25063 a_n17362_8608.n0 a_n17362_8608.n18 11.1777
R25064 a_n17362_8608.n0 a_n17362_8608.n15 8.95524
R25065 a_n17362_8608.n15 a_n17362_8608.n13 8.91593
R25066 a_n17362_8608.n18 a_n17362_8608.n16 8.91593
R25067 a_n17362_8608.n15 a_n17362_8608.n14 6.21896
R25068 a_n17362_8608.n18 a_n17362_8608.n17 6.21896
R25069 VN.n133 VN.n132 161.3
R25070 VN.n134 VN.n129 161.3
R25071 VN.n136 VN.n135 161.3
R25072 VN.n137 VN.n128 161.3
R25073 VN.n139 VN.n138 161.3
R25074 VN.n140 VN.n127 161.3
R25075 VN.n142 VN.n141 161.3
R25076 VN.n143 VN.n126 161.3
R25077 VN.n145 VN.n144 161.3
R25078 VN.n146 VN.n125 161.3
R25079 VN.n148 VN.n147 161.3
R25080 VN.n149 VN.n124 161.3
R25081 VN.n152 VN.n151 161.3
R25082 VN.n153 VN.n123 161.3
R25083 VN.n155 VN.n154 161.3
R25084 VN.n156 VN.n122 161.3
R25085 VN.n158 VN.n157 161.3
R25086 VN.n159 VN.n121 161.3
R25087 VN.n161 VN.n160 161.3
R25088 VN.n162 VN.n120 161.3
R25089 VN.n164 VN.n163 161.3
R25090 VN.n165 VN.n119 161.3
R25091 VN.n167 VN.n166 161.3
R25092 VN.n168 VN.n118 161.3
R25093 VN.n171 VN.n170 161.3
R25094 VN.n172 VN.n117 161.3
R25095 VN.n174 VN.n173 161.3
R25096 VN.n175 VN.n116 161.3
R25097 VN.n177 VN.n176 161.3
R25098 VN.n178 VN.n115 161.3
R25099 VN.n180 VN.n179 161.3
R25100 VN.n181 VN.n114 161.3
R25101 VN.n183 VN.n182 161.3
R25102 VN.n184 VN.n113 161.3
R25103 VN.n186 VN.n185 161.3
R25104 VN.n187 VN.n112 161.3
R25105 VN.n190 VN.n189 161.3
R25106 VN.n191 VN.n111 161.3
R25107 VN.n193 VN.n192 161.3
R25108 VN.n194 VN.n110 161.3
R25109 VN.n196 VN.n195 161.3
R25110 VN.n197 VN.n109 161.3
R25111 VN.n199 VN.n198 161.3
R25112 VN.n200 VN.n108 161.3
R25113 VN.n202 VN.n201 161.3
R25114 VN.n203 VN.n107 161.3
R25115 VN.n205 VN.n204 161.3
R25116 VN.n206 VN.n106 161.3
R25117 VN.n208 VN.n207 161.3
R25118 VN.n30 VN.n29 161.3
R25119 VN.n31 VN.n26 161.3
R25120 VN.n33 VN.n32 161.3
R25121 VN.n34 VN.n25 161.3
R25122 VN.n36 VN.n35 161.3
R25123 VN.n37 VN.n24 161.3
R25124 VN.n39 VN.n38 161.3
R25125 VN.n40 VN.n23 161.3
R25126 VN.n42 VN.n41 161.3
R25127 VN.n43 VN.n22 161.3
R25128 VN.n45 VN.n44 161.3
R25129 VN.n46 VN.n21 161.3
R25130 VN.n49 VN.n48 161.3
R25131 VN.n50 VN.n20 161.3
R25132 VN.n52 VN.n51 161.3
R25133 VN.n53 VN.n19 161.3
R25134 VN.n55 VN.n54 161.3
R25135 VN.n56 VN.n18 161.3
R25136 VN.n58 VN.n57 161.3
R25137 VN.n59 VN.n17 161.3
R25138 VN.n61 VN.n60 161.3
R25139 VN.n62 VN.n16 161.3
R25140 VN.n64 VN.n63 161.3
R25141 VN.n65 VN.n14 161.3
R25142 VN.n67 VN.n66 161.3
R25143 VN.n68 VN.n13 161.3
R25144 VN.n70 VN.n69 161.3
R25145 VN.n71 VN.n12 161.3
R25146 VN.n73 VN.n72 161.3
R25147 VN.n74 VN.n11 161.3
R25148 VN.n76 VN.n75 161.3
R25149 VN.n77 VN.n10 161.3
R25150 VN.n79 VN.n78 161.3
R25151 VN.n80 VN.n9 161.3
R25152 VN.n82 VN.n81 161.3
R25153 VN.n83 VN.n7 161.3
R25154 VN.n85 VN.n84 161.3
R25155 VN.n86 VN.n6 161.3
R25156 VN.n88 VN.n87 161.3
R25157 VN.n89 VN.n5 161.3
R25158 VN.n91 VN.n90 161.3
R25159 VN.n92 VN.n4 161.3
R25160 VN.n94 VN.n93 161.3
R25161 VN.n95 VN.n3 161.3
R25162 VN.n97 VN.n96 161.3
R25163 VN.n98 VN.n2 161.3
R25164 VN.n100 VN.n99 161.3
R25165 VN.n101 VN.n1 161.3
R25166 VN.n103 VN.n102 161.3
R25167 VN.n200 VN.n199 72.0595
R25168 VN.n95 VN.n94 72.0595
R25169 VN.n131 VN.n130 70.3045
R25170 VN.n28 VN.n27 70.3045
R25171 VN.n209 VN.n105 69.0311
R25172 VN.n104 VN.n0 69.0311
R25173 VN.n181 VN.n180 64.2894
R25174 VN.n142 VN.n127 64.2894
R25175 VN.n77 VN.n76 64.2894
R25176 VN.n39 VN.n24 64.2894
R25177 VN.n210 VN.n209 57.0542
R25178 VN.n162 VN.n161 56.5193
R25179 VN.n161 VN.n121 56.5193
R25180 VN.n59 VN.n58 56.5193
R25181 VN.n58 VN.n18 56.5193
R25182 VN.n180 VN.n115 48.7492
R25183 VN.n143 VN.n142 48.7492
R25184 VN.n76 VN.n11 48.7492
R25185 VN.n40 VN.n39 48.7492
R25186 VN.n130 VN.t6 46.6431
R25187 VN.n27 VN.t5 46.6431
R25188 VN.n199 VN.n109 40.979
R25189 VN.n94 VN.n4 40.979
R25190 VN.n201 VN.n200 24.4675
R25191 VN.n201 VN.n107 24.4675
R25192 VN.n205 VN.n107 24.4675
R25193 VN.n206 VN.n205 24.4675
R25194 VN.n207 VN.n206 24.4675
R25195 VN.n182 VN.n181 24.4675
R25196 VN.n182 VN.n113 24.4675
R25197 VN.n186 VN.n113 24.4675
R25198 VN.n187 VN.n186 24.4675
R25199 VN.n189 VN.n187 24.4675
R25200 VN.n193 VN.n111 24.4675
R25201 VN.n194 VN.n193 24.4675
R25202 VN.n195 VN.n194 24.4675
R25203 VN.n195 VN.n109 24.4675
R25204 VN.n163 VN.n162 24.4675
R25205 VN.n163 VN.n119 24.4675
R25206 VN.n167 VN.n119 24.4675
R25207 VN.n168 VN.n167 24.4675
R25208 VN.n170 VN.n168 24.4675
R25209 VN.n174 VN.n117 24.4675
R25210 VN.n175 VN.n174 24.4675
R25211 VN.n176 VN.n175 24.4675
R25212 VN.n176 VN.n115 24.4675
R25213 VN.n144 VN.n143 24.4675
R25214 VN.n144 VN.n125 24.4675
R25215 VN.n148 VN.n125 24.4675
R25216 VN.n149 VN.n148 24.4675
R25217 VN.n151 VN.n123 24.4675
R25218 VN.n155 VN.n123 24.4675
R25219 VN.n156 VN.n155 24.4675
R25220 VN.n157 VN.n156 24.4675
R25221 VN.n157 VN.n121 24.4675
R25222 VN.n132 VN.n129 24.4675
R25223 VN.n136 VN.n129 24.4675
R25224 VN.n137 VN.n136 24.4675
R25225 VN.n138 VN.n137 24.4675
R25226 VN.n138 VN.n127 24.4675
R25227 VN.n102 VN.n101 24.4675
R25228 VN.n101 VN.n100 24.4675
R25229 VN.n100 VN.n2 24.4675
R25230 VN.n96 VN.n2 24.4675
R25231 VN.n96 VN.n95 24.4675
R25232 VN.n90 VN.n4 24.4675
R25233 VN.n90 VN.n89 24.4675
R25234 VN.n89 VN.n88 24.4675
R25235 VN.n88 VN.n6 24.4675
R25236 VN.n84 VN.n83 24.4675
R25237 VN.n83 VN.n82 24.4675
R25238 VN.n82 VN.n9 24.4675
R25239 VN.n78 VN.n9 24.4675
R25240 VN.n78 VN.n77 24.4675
R25241 VN.n72 VN.n11 24.4675
R25242 VN.n72 VN.n71 24.4675
R25243 VN.n71 VN.n70 24.4675
R25244 VN.n70 VN.n13 24.4675
R25245 VN.n66 VN.n65 24.4675
R25246 VN.n65 VN.n64 24.4675
R25247 VN.n64 VN.n16 24.4675
R25248 VN.n60 VN.n16 24.4675
R25249 VN.n60 VN.n59 24.4675
R25250 VN.n54 VN.n18 24.4675
R25251 VN.n54 VN.n53 24.4675
R25252 VN.n53 VN.n52 24.4675
R25253 VN.n52 VN.n20 24.4675
R25254 VN.n48 VN.n20 24.4675
R25255 VN.n46 VN.n45 24.4675
R25256 VN.n45 VN.n22 24.4675
R25257 VN.n41 VN.n22 24.4675
R25258 VN.n41 VN.n40 24.4675
R25259 VN.n35 VN.n24 24.4675
R25260 VN.n35 VN.n34 24.4675
R25261 VN.n34 VN.n33 24.4675
R25262 VN.n33 VN.n26 24.4675
R25263 VN.n29 VN.n26 24.4675
R25264 VN.n169 VN.n117 22.5101
R25265 VN.n150 VN.n149 22.5101
R25266 VN.n15 VN.n13 22.5101
R25267 VN.n47 VN.n46 22.5101
R25268 VN VN.n210 20.9445
R25269 VN.n188 VN.n111 18.5954
R25270 VN.n8 VN.n6 18.5954
R25271 VN.n210 VN.n104 13.1527
R25272 VN.n105 VN.t1 12.9398
R25273 VN.n188 VN.t4 12.9398
R25274 VN.n169 VN.t0 12.9398
R25275 VN.n150 VN.t8 12.9398
R25276 VN.n131 VN.t11 12.9398
R25277 VN.n0 VN.t2 12.9398
R25278 VN.n8 VN.t3 12.9398
R25279 VN.n15 VN.t7 12.9398
R25280 VN.n47 VN.t9 12.9398
R25281 VN.n28 VN.t10 12.9398
R25282 VN.n207 VN.n105 9.7873
R25283 VN.n102 VN.n0 9.7873
R25284 VN.n189 VN.n188 5.87258
R25285 VN.n132 VN.n131 5.87258
R25286 VN.n84 VN.n8 5.87258
R25287 VN.n29 VN.n28 5.87258
R25288 VN.n170 VN.n169 1.95786
R25289 VN.n151 VN.n150 1.95786
R25290 VN.n66 VN.n15 1.95786
R25291 VN.n48 VN.n47 1.95786
R25292 VN.n133 VN.n130 0.976619
R25293 VN.n30 VN.n27 0.976619
R25294 VN.n209 VN.n208 0.466196
R25295 VN.n104 VN.n103 0.466196
R25296 VN.n134 VN.n133 0.189894
R25297 VN.n135 VN.n134 0.189894
R25298 VN.n135 VN.n128 0.189894
R25299 VN.n139 VN.n128 0.189894
R25300 VN.n140 VN.n139 0.189894
R25301 VN.n141 VN.n140 0.189894
R25302 VN.n141 VN.n126 0.189894
R25303 VN.n145 VN.n126 0.189894
R25304 VN.n146 VN.n145 0.189894
R25305 VN.n147 VN.n146 0.189894
R25306 VN.n147 VN.n124 0.189894
R25307 VN.n152 VN.n124 0.189894
R25308 VN.n153 VN.n152 0.189894
R25309 VN.n154 VN.n153 0.189894
R25310 VN.n154 VN.n122 0.189894
R25311 VN.n158 VN.n122 0.189894
R25312 VN.n159 VN.n158 0.189894
R25313 VN.n160 VN.n159 0.189894
R25314 VN.n160 VN.n120 0.189894
R25315 VN.n164 VN.n120 0.189894
R25316 VN.n165 VN.n164 0.189894
R25317 VN.n166 VN.n165 0.189894
R25318 VN.n166 VN.n118 0.189894
R25319 VN.n171 VN.n118 0.189894
R25320 VN.n172 VN.n171 0.189894
R25321 VN.n173 VN.n172 0.189894
R25322 VN.n173 VN.n116 0.189894
R25323 VN.n177 VN.n116 0.189894
R25324 VN.n178 VN.n177 0.189894
R25325 VN.n179 VN.n178 0.189894
R25326 VN.n179 VN.n114 0.189894
R25327 VN.n183 VN.n114 0.189894
R25328 VN.n184 VN.n183 0.189894
R25329 VN.n185 VN.n184 0.189894
R25330 VN.n185 VN.n112 0.189894
R25331 VN.n190 VN.n112 0.189894
R25332 VN.n191 VN.n190 0.189894
R25333 VN.n192 VN.n191 0.189894
R25334 VN.n192 VN.n110 0.189894
R25335 VN.n196 VN.n110 0.189894
R25336 VN.n197 VN.n196 0.189894
R25337 VN.n198 VN.n197 0.189894
R25338 VN.n198 VN.n108 0.189894
R25339 VN.n202 VN.n108 0.189894
R25340 VN.n203 VN.n202 0.189894
R25341 VN.n204 VN.n203 0.189894
R25342 VN.n204 VN.n106 0.189894
R25343 VN.n208 VN.n106 0.189894
R25344 VN.n103 VN.n1 0.189894
R25345 VN.n99 VN.n1 0.189894
R25346 VN.n99 VN.n98 0.189894
R25347 VN.n98 VN.n97 0.189894
R25348 VN.n97 VN.n3 0.189894
R25349 VN.n93 VN.n3 0.189894
R25350 VN.n93 VN.n92 0.189894
R25351 VN.n92 VN.n91 0.189894
R25352 VN.n91 VN.n5 0.189894
R25353 VN.n87 VN.n5 0.189894
R25354 VN.n87 VN.n86 0.189894
R25355 VN.n86 VN.n85 0.189894
R25356 VN.n85 VN.n7 0.189894
R25357 VN.n81 VN.n7 0.189894
R25358 VN.n81 VN.n80 0.189894
R25359 VN.n80 VN.n79 0.189894
R25360 VN.n79 VN.n10 0.189894
R25361 VN.n75 VN.n10 0.189894
R25362 VN.n75 VN.n74 0.189894
R25363 VN.n74 VN.n73 0.189894
R25364 VN.n73 VN.n12 0.189894
R25365 VN.n69 VN.n12 0.189894
R25366 VN.n69 VN.n68 0.189894
R25367 VN.n68 VN.n67 0.189894
R25368 VN.n67 VN.n14 0.189894
R25369 VN.n63 VN.n14 0.189894
R25370 VN.n63 VN.n62 0.189894
R25371 VN.n62 VN.n61 0.189894
R25372 VN.n61 VN.n17 0.189894
R25373 VN.n57 VN.n17 0.189894
R25374 VN.n57 VN.n56 0.189894
R25375 VN.n56 VN.n55 0.189894
R25376 VN.n55 VN.n19 0.189894
R25377 VN.n51 VN.n19 0.189894
R25378 VN.n51 VN.n50 0.189894
R25379 VN.n50 VN.n49 0.189894
R25380 VN.n49 VN.n21 0.189894
R25381 VN.n44 VN.n21 0.189894
R25382 VN.n44 VN.n43 0.189894
R25383 VN.n43 VN.n42 0.189894
R25384 VN.n42 VN.n23 0.189894
R25385 VN.n38 VN.n23 0.189894
R25386 VN.n38 VN.n37 0.189894
R25387 VN.n37 VN.n36 0.189894
R25388 VN.n36 VN.n25 0.189894
R25389 VN.n32 VN.n25 0.189894
R25390 VN.n32 VN.n31 0.189894
R25391 VN.n31 VN.n30 0.189894
C0 VDD VN 0.09836f
C1 VOUT CS_BIAS 42.5062f
C2 a_n13259_9690# VDD 1.88516f
C3 VOUT VN 1.28096f
C4 VOUT VP 3.58819f
C5 CS_BIAS VN 0.315346f
C6 CS_BIAS VP 0.393257f
C7 VN VP 17.4083f
C8 VN DIFFPAIR_BIAS 9.01e-20
C9 VP DIFFPAIR_BIAS 9.01e-20
C10 a_11817_9690# VDD 1.88517f
C11 VDD VOUT 22.471802f
C12 DIFFPAIR_BIAS GND 18.0931f
C13 VP GND 50.19553f
C14 VN GND 65.0381f
C15 CS_BIAS GND 0.229178p
C16 VOUT GND 0.122812p
C17 VDD GND 0.576774p
C18 a_11817_9690# GND 0.738921f
C19 a_n13259_9690# GND 0.738921f
C20 VN.t2 GND 0.512858f
C21 VN.n0 GND 0.260315f
C22 VN.n1 GND 0.013104f
C23 VN.n2 GND 0.024422f
C24 VN.n3 GND 0.013104f
C25 VN.n4 GND 0.025977f
C26 VN.n5 GND 0.013104f
C27 VN.n6 GND 0.021529f
C28 VN.n7 GND 0.013104f
C29 VN.t3 GND 0.512858f
C30 VN.n8 GND 0.205126f
C31 VN.n9 GND 0.024422f
C32 VN.n10 GND 0.013104f
C33 VN.n11 GND 0.024422f
C34 VN.n12 GND 0.013104f
C35 VN.n13 GND 0.023458f
C36 VN.n14 GND 0.013104f
C37 VN.t7 GND 0.512858f
C38 VN.n15 GND 0.205126f
C39 VN.n16 GND 0.024422f
C40 VN.n17 GND 0.013104f
C41 VN.n18 GND 0.022234f
C42 VN.n19 GND 0.013104f
C43 VN.n20 GND 0.024422f
C44 VN.n21 GND 0.013104f
C45 VN.t9 GND 0.512858f
C46 VN.n22 GND 0.024422f
C47 VN.n23 GND 0.013104f
C48 VN.n24 GND 0.019642f
C49 VN.n25 GND 0.013104f
C50 VN.n26 GND 0.024422f
C51 VN.t5 GND 0.748638f
C52 VN.n27 GND 0.39055f
C53 VN.t10 GND 0.512858f
C54 VN.n28 GND 0.254926f
C55 VN.n29 GND 0.015259f
C56 VN.n30 GND 0.154226f
C57 VN.n31 GND 0.013104f
C58 VN.n32 GND 0.013104f
C59 VN.n33 GND 0.024422f
C60 VN.n34 GND 0.024422f
C61 VN.n35 GND 0.024422f
C62 VN.n36 GND 0.013104f
C63 VN.n37 GND 0.013104f
C64 VN.n38 GND 0.013104f
C65 VN.n39 GND 0.008035f
C66 VN.n40 GND 0.024422f
C67 VN.n41 GND 0.024422f
C68 VN.n42 GND 0.013104f
C69 VN.n43 GND 0.013104f
C70 VN.n44 GND 0.013104f
C71 VN.n45 GND 0.024422f
C72 VN.n46 GND 0.023458f
C73 VN.n47 GND 0.205126f
C74 VN.n48 GND 0.01333f
C75 VN.n49 GND 0.013104f
C76 VN.n50 GND 0.013104f
C77 VN.n51 GND 0.013104f
C78 VN.n52 GND 0.024422f
C79 VN.n53 GND 0.024422f
C80 VN.n54 GND 0.024422f
C81 VN.n55 GND 0.013104f
C82 VN.n56 GND 0.013104f
C83 VN.n57 GND 0.013104f
C84 VN.n58 GND 0.007631f
C85 VN.n59 GND 0.022234f
C86 VN.n60 GND 0.024422f
C87 VN.n61 GND 0.013104f
C88 VN.n62 GND 0.013104f
C89 VN.n63 GND 0.013104f
C90 VN.n64 GND 0.024422f
C91 VN.n65 GND 0.024422f
C92 VN.n66 GND 0.01333f
C93 VN.n67 GND 0.013104f
C94 VN.n68 GND 0.013104f
C95 VN.n69 GND 0.013104f
C96 VN.n70 GND 0.024422f
C97 VN.n71 GND 0.024422f
C98 VN.n72 GND 0.024422f
C99 VN.n73 GND 0.013104f
C100 VN.n74 GND 0.013104f
C101 VN.n75 GND 0.013104f
C102 VN.n76 GND 0.008035f
C103 VN.n77 GND 0.019642f
C104 VN.n78 GND 0.024422f
C105 VN.n79 GND 0.013104f
C106 VN.n80 GND 0.013104f
C107 VN.n81 GND 0.013104f
C108 VN.n82 GND 0.024422f
C109 VN.n83 GND 0.024422f
C110 VN.n84 GND 0.015259f
C111 VN.n85 GND 0.013104f
C112 VN.n86 GND 0.013104f
C113 VN.n87 GND 0.013104f
C114 VN.n88 GND 0.024422f
C115 VN.n89 GND 0.024422f
C116 VN.n90 GND 0.024422f
C117 VN.n91 GND 0.013104f
C118 VN.n92 GND 0.013104f
C119 VN.n93 GND 0.013104f
C120 VN.n94 GND 0.009345f
C121 VN.n95 GND 0.016777f
C122 VN.n96 GND 0.024422f
C123 VN.n97 GND 0.013104f
C124 VN.n98 GND 0.013104f
C125 VN.n99 GND 0.013104f
C126 VN.n100 GND 0.024422f
C127 VN.n101 GND 0.024422f
C128 VN.n102 GND 0.017188f
C129 VN.n103 GND 0.027728f
C130 VN.n104 GND 0.290541f
C131 VN.t1 GND 0.512858f
C132 VN.n105 GND 0.260315f
C133 VN.n106 GND 0.013104f
C134 VN.n107 GND 0.024422f
C135 VN.n108 GND 0.013104f
C136 VN.n109 GND 0.025977f
C137 VN.n110 GND 0.013104f
C138 VN.n111 GND 0.021529f
C139 VN.n112 GND 0.013104f
C140 VN.n113 GND 0.024422f
C141 VN.n114 GND 0.013104f
C142 VN.n115 GND 0.024422f
C143 VN.n116 GND 0.013104f
C144 VN.n117 GND 0.023458f
C145 VN.n118 GND 0.013104f
C146 VN.n119 GND 0.024422f
C147 VN.n120 GND 0.013104f
C148 VN.n121 GND 0.022234f
C149 VN.n122 GND 0.013104f
C150 VN.n123 GND 0.024422f
C151 VN.n124 GND 0.013104f
C152 VN.t8 GND 0.512858f
C153 VN.n125 GND 0.024422f
C154 VN.n126 GND 0.013104f
C155 VN.n127 GND 0.019642f
C156 VN.n128 GND 0.013104f
C157 VN.n129 GND 0.024422f
C158 VN.t6 GND 0.748638f
C159 VN.n130 GND 0.39055f
C160 VN.t11 GND 0.512858f
C161 VN.n131 GND 0.254926f
C162 VN.n132 GND 0.015259f
C163 VN.n133 GND 0.154226f
C164 VN.n134 GND 0.013104f
C165 VN.n135 GND 0.013104f
C166 VN.n136 GND 0.024422f
C167 VN.n137 GND 0.024422f
C168 VN.n138 GND 0.024422f
C169 VN.n139 GND 0.013104f
C170 VN.n140 GND 0.013104f
C171 VN.n141 GND 0.013104f
C172 VN.n142 GND 0.008035f
C173 VN.n143 GND 0.024422f
C174 VN.n144 GND 0.024422f
C175 VN.n145 GND 0.013104f
C176 VN.n146 GND 0.013104f
C177 VN.n147 GND 0.013104f
C178 VN.n148 GND 0.024422f
C179 VN.n149 GND 0.023458f
C180 VN.n150 GND 0.205126f
C181 VN.n151 GND 0.01333f
C182 VN.n152 GND 0.013104f
C183 VN.n153 GND 0.013104f
C184 VN.n154 GND 0.013104f
C185 VN.n155 GND 0.024422f
C186 VN.n156 GND 0.024422f
C187 VN.n157 GND 0.024422f
C188 VN.n158 GND 0.013104f
C189 VN.n159 GND 0.013104f
C190 VN.n160 GND 0.013104f
C191 VN.n161 GND 0.007631f
C192 VN.n162 GND 0.022234f
C193 VN.n163 GND 0.024422f
C194 VN.n164 GND 0.013104f
C195 VN.n165 GND 0.013104f
C196 VN.n166 GND 0.013104f
C197 VN.n167 GND 0.024422f
C198 VN.n168 GND 0.024422f
C199 VN.t0 GND 0.512858f
C200 VN.n169 GND 0.205126f
C201 VN.n170 GND 0.01333f
C202 VN.n171 GND 0.013104f
C203 VN.n172 GND 0.013104f
C204 VN.n173 GND 0.013104f
C205 VN.n174 GND 0.024422f
C206 VN.n175 GND 0.024422f
C207 VN.n176 GND 0.024422f
C208 VN.n177 GND 0.013104f
C209 VN.n178 GND 0.013104f
C210 VN.n179 GND 0.013104f
C211 VN.n180 GND 0.008035f
C212 VN.n181 GND 0.019642f
C213 VN.n182 GND 0.024422f
C214 VN.n183 GND 0.013104f
C215 VN.n184 GND 0.013104f
C216 VN.n185 GND 0.013104f
C217 VN.n186 GND 0.024422f
C218 VN.n187 GND 0.024422f
C219 VN.t4 GND 0.512858f
C220 VN.n188 GND 0.205126f
C221 VN.n189 GND 0.015259f
C222 VN.n190 GND 0.013104f
C223 VN.n191 GND 0.013104f
C224 VN.n192 GND 0.013104f
C225 VN.n193 GND 0.024422f
C226 VN.n194 GND 0.024422f
C227 VN.n195 GND 0.024422f
C228 VN.n196 GND 0.013104f
C229 VN.n197 GND 0.013104f
C230 VN.n198 GND 0.013104f
C231 VN.n199 GND 0.009345f
C232 VN.n200 GND 0.016777f
C233 VN.n201 GND 0.024422f
C234 VN.n202 GND 0.013104f
C235 VN.n203 GND 0.013104f
C236 VN.n204 GND 0.013104f
C237 VN.n205 GND 0.024422f
C238 VN.n206 GND 0.024422f
C239 VN.n207 GND 0.017188f
C240 VN.n208 GND 0.027728f
C241 VN.n209 GND 1.0074f
C242 VN.n210 GND 4.85797f
C243 a_n17362_8608.n0 GND 25.4333f
C244 a_n17362_8608.n1 GND 8.35256f
C245 a_n17362_8608.t16 GND 0.039098f
C246 a_n17362_8608.t14 GND 0.039098f
C247 a_n17362_8608.t11 GND 0.039098f
C248 a_n17362_8608.n2 GND 0.179945f
C249 a_n17362_8608.t15 GND 0.039098f
C250 a_n17362_8608.t17 GND 0.039098f
C251 a_n17362_8608.n3 GND 0.179945f
C252 a_n17362_8608.t13 GND 0.039098f
C253 a_n17362_8608.t12 GND 0.039098f
C254 a_n17362_8608.n4 GND 0.162932f
C255 a_n17362_8608.n5 GND 8.00958f
C256 a_n17362_8608.t4 GND 0.054699f
C257 a_n17362_8608.t2 GND 0.054699f
C258 a_n17362_8608.n6 GND 0.384858f
C259 a_n17362_8608.t0 GND 0.054699f
C260 a_n17362_8608.t19 GND 0.054699f
C261 a_n17362_8608.n7 GND 0.353883f
C262 a_n17362_8608.t9 GND 0.054699f
C263 a_n17362_8608.t8 GND 0.054699f
C264 a_n17362_8608.n8 GND 0.384857f
C265 a_n17362_8608.t5 GND 0.054699f
C266 a_n17362_8608.t1 GND 0.054699f
C267 a_n17362_8608.n9 GND 0.353883f
C268 a_n17362_8608.t3 GND 0.054699f
C269 a_n17362_8608.t6 GND 0.054699f
C270 a_n17362_8608.n10 GND 0.384857f
C271 a_n17362_8608.n11 GND 8.41179f
C272 a_n17362_8608.t7 GND 0.054699f
C273 a_n17362_8608.t10 GND 0.054699f
C274 a_n17362_8608.n12 GND 0.353883f
C275 a_n17362_8608.t22 GND 1.66108f
C276 a_n17362_8608.t25 GND 1.63912f
C277 a_n17362_8608.n13 GND 1.528f
C278 a_n17362_8608.t27 GND 1.66108f
C279 a_n17362_8608.t21 GND 1.63912f
C280 a_n17362_8608.n14 GND 1.45383f
C281 a_n17362_8608.n15 GND 3.57481f
C282 a_n17362_8608.t26 GND 1.63912f
C283 a_n17362_8608.t20 GND 1.66108f
C284 a_n17362_8608.n16 GND 1.528f
C285 a_n17362_8608.t24 GND 1.63912f
C286 a_n17362_8608.t23 GND 1.66108f
C287 a_n17362_8608.n17 GND 1.45383f
C288 a_n17362_8608.n18 GND 1.96266f
C289 a_n17362_8608.n19 GND 12.7443f
C290 a_n17362_8608.n20 GND 6.67535f
C291 a_n17362_8608.n21 GND 0.162931f
C292 a_n17362_8608.t18 GND 0.039098f
C293 a_n7386_8166.n0 GND 9.543571f
C294 a_n7386_8166.n1 GND 5.77171f
C295 a_n7386_8166.n2 GND 4.63214f
C296 a_n7386_8166.n3 GND 3.32359f
C297 a_n7386_8166.n4 GND 7.34636f
C298 a_n7386_8166.t16 GND 73.3396f
C299 a_n7386_8166.t0 GND 0.204722f
C300 a_n7386_8166.t1 GND 0.040315f
C301 a_n7386_8166.t13 GND 0.040315f
C302 a_n7386_8166.n5 GND 0.132665f
C303 a_n7386_8166.t3 GND 0.19514f
C304 a_n7386_8166.t9 GND 0.204722f
C305 a_n7386_8166.t11 GND 0.040315f
C306 a_n7386_8166.t6 GND 0.040315f
C307 a_n7386_8166.n6 GND 0.132665f
C308 a_n7386_8166.t10 GND 0.19514f
C309 a_n7386_8166.t8 GND 0.19514f
C310 a_n7386_8166.t7 GND 0.040315f
C311 a_n7386_8166.t5 GND 0.040315f
C312 a_n7386_8166.n7 GND 0.132665f
C313 a_n7386_8166.t12 GND 0.19514f
C314 a_n7386_8166.t2 GND 0.204721f
C315 a_n7386_8166.t14 GND 0.040315f
C316 a_n7386_8166.t15 GND 0.040315f
C317 a_n7386_8166.n8 GND 0.132665f
C318 a_n7386_8166.t4 GND 0.19514f
C319 VOUT.t2 GND 0.030708f
C320 VOUT.t55 GND 0.030708f
C321 VOUT.n0 GND 0.191636f
C322 VOUT.t57 GND 0.030708f
C323 VOUT.t1 GND 0.030708f
C324 VOUT.n1 GND 0.184567f
C325 VOUT.n2 GND 2.00031f
C326 VOUT.n3 GND 8.044491f
C327 VOUT.t58 GND 24.846401f
C328 VOUT.t59 GND 15.075599f
C329 VOUT.n4 GND 14.3873f
C330 VOUT.n5 GND 1.9233f
C331 VOUT.t0 GND 0.030708f
C332 VOUT.t4 GND 0.030708f
C333 VOUT.n6 GND 0.191636f
C334 VOUT.t3 GND 0.030708f
C335 VOUT.t56 GND 0.030708f
C336 VOUT.n7 GND 0.184566f
C337 VOUT.n8 GND 2.00031f
C338 VOUT.n9 GND 9.71271f
C339 VOUT.t24 GND 0.12736f
C340 VOUT.t31 GND 0.016853f
C341 VOUT.t16 GND 0.016853f
C342 VOUT.n10 GND 0.10378f
C343 VOUT.n11 GND 1.00262f
C344 VOUT.t30 GND 0.016853f
C345 VOUT.t12 GND 0.016853f
C346 VOUT.n12 GND 0.10378f
C347 VOUT.n13 GND 0.707146f
C348 VOUT.t32 GND 0.12736f
C349 VOUT.t26 GND 0.016853f
C350 VOUT.t42 GND 0.016853f
C351 VOUT.n14 GND 0.10378f
C352 VOUT.n15 GND 1.00262f
C353 VOUT.t13 GND 0.016853f
C354 VOUT.t25 GND 0.016853f
C355 VOUT.n16 GND 0.10378f
C356 VOUT.n17 GND 0.68678f
C357 VOUT.n18 GND 0.423694f
C358 VOUT.t5 GND 0.12736f
C359 VOUT.t35 GND 0.016853f
C360 VOUT.t44 GND 0.016853f
C361 VOUT.n19 GND 0.10378f
C362 VOUT.n20 GND 1.00262f
C363 VOUT.t21 GND 0.016853f
C364 VOUT.t27 GND 0.016853f
C365 VOUT.n21 GND 0.10378f
C366 VOUT.n22 GND 0.68678f
C367 VOUT.n23 GND 0.276233f
C368 VOUT.t6 GND 0.12736f
C369 VOUT.t36 GND 0.016853f
C370 VOUT.t45 GND 0.016853f
C371 VOUT.n24 GND 0.10378f
C372 VOUT.n25 GND 1.00262f
C373 VOUT.t22 GND 0.016853f
C374 VOUT.t28 GND 0.016853f
C375 VOUT.n26 GND 0.10378f
C376 VOUT.n27 GND 0.68678f
C377 VOUT.n28 GND 0.276233f
C378 VOUT.t7 GND 0.12736f
C379 VOUT.t38 GND 0.016853f
C380 VOUT.t48 GND 0.016853f
C381 VOUT.n29 GND 0.10378f
C382 VOUT.n30 GND 1.00262f
C383 VOUT.t23 GND 0.016853f
C384 VOUT.t29 GND 0.016853f
C385 VOUT.n31 GND 0.10378f
C386 VOUT.n32 GND 0.68678f
C387 VOUT.n33 GND 0.457525f
C388 VOUT.n34 GND 9.70605f
C389 VOUT.t41 GND 0.016853f
C390 VOUT.t19 GND 0.016853f
C391 VOUT.n35 GND 0.116835f
C392 VOUT.t51 GND 0.016853f
C393 VOUT.t20 GND 0.016853f
C394 VOUT.n36 GND 0.10378f
C395 VOUT.n37 GND 1.24588f
C396 VOUT.t50 GND 0.120855f
C397 VOUT.n38 GND 0.492865f
C398 VOUT.t18 GND 0.016853f
C399 VOUT.t49 GND 0.016853f
C400 VOUT.n39 GND 0.116835f
C401 VOUT.t10 GND 0.016853f
C402 VOUT.t40 GND 0.016853f
C403 VOUT.n40 GND 0.10378f
C404 VOUT.n41 GND 1.24588f
C405 VOUT.t39 GND 0.120855f
C406 VOUT.n42 GND 0.474459f
C407 VOUT.n43 GND 0.35069f
C408 VOUT.t43 GND 0.016853f
C409 VOUT.t34 GND 0.016853f
C410 VOUT.n44 GND 0.116835f
C411 VOUT.t14 GND 0.016853f
C412 VOUT.t52 GND 0.016853f
C413 VOUT.n45 GND 0.10378f
C414 VOUT.n46 GND 1.24588f
C415 VOUT.t9 GND 0.120855f
C416 VOUT.n47 GND 0.474459f
C417 VOUT.n48 GND 0.238751f
C418 VOUT.t47 GND 0.016853f
C419 VOUT.t33 GND 0.016853f
C420 VOUT.n49 GND 0.116835f
C421 VOUT.t15 GND 0.016853f
C422 VOUT.t54 GND 0.016853f
C423 VOUT.n50 GND 0.10378f
C424 VOUT.n51 GND 1.24588f
C425 VOUT.t8 GND 0.120855f
C426 VOUT.n52 GND 0.474459f
C427 VOUT.n53 GND 0.238751f
C428 VOUT.t46 GND 0.016853f
C429 VOUT.t37 GND 0.016853f
C430 VOUT.n54 GND 0.116835f
C431 VOUT.t17 GND 0.016853f
C432 VOUT.t53 GND 0.016853f
C433 VOUT.n55 GND 0.10378f
C434 VOUT.n56 GND 1.24588f
C435 VOUT.t11 GND 0.120855f
C436 VOUT.n57 GND 0.474459f
C437 VOUT.n58 GND 0.420043f
C438 VOUT.n59 GND 7.592f
C439 VOUT.n60 GND 3.92026f
C440 VP.t4 GND 0.775277f
C441 VP.n0 GND 0.393512f
C442 VP.n1 GND 0.019809f
C443 VP.n2 GND 0.036919f
C444 VP.n3 GND 0.019809f
C445 VP.n4 GND 0.039269f
C446 VP.n5 GND 0.019809f
C447 VP.n6 GND 0.032544f
C448 VP.n7 GND 0.019809f
C449 VP.n8 GND 0.036919f
C450 VP.n9 GND 0.019809f
C451 VP.n10 GND 0.036919f
C452 VP.n11 GND 0.019809f
C453 VP.n12 GND 0.03546f
C454 VP.n13 GND 0.019809f
C455 VP.n14 GND 0.036919f
C456 VP.n15 GND 0.019809f
C457 VP.n16 GND 0.033611f
C458 VP.n17 GND 0.019809f
C459 VP.n18 GND 0.036919f
C460 VP.n19 GND 0.019809f
C461 VP.t11 GND 0.775277f
C462 VP.n20 GND 0.036919f
C463 VP.n21 GND 0.019809f
C464 VP.n22 GND 0.029693f
C465 VP.n23 GND 0.019809f
C466 VP.n24 GND 0.036919f
C467 VP.t8 GND 1.1317f
C468 VP.n25 GND 0.590385f
C469 VP.t0 GND 0.775277f
C470 VP.n26 GND 0.385367f
C471 VP.n27 GND 0.023066f
C472 VP.n28 GND 0.23314f
C473 VP.n29 GND 0.019809f
C474 VP.n30 GND 0.019809f
C475 VP.n31 GND 0.036919f
C476 VP.n32 GND 0.036919f
C477 VP.n33 GND 0.036919f
C478 VP.n34 GND 0.019809f
C479 VP.n35 GND 0.019809f
C480 VP.n36 GND 0.019809f
C481 VP.n37 GND 0.012146f
C482 VP.n38 GND 0.036919f
C483 VP.n39 GND 0.036919f
C484 VP.n40 GND 0.019809f
C485 VP.n41 GND 0.019809f
C486 VP.n42 GND 0.019809f
C487 VP.n43 GND 0.036919f
C488 VP.n44 GND 0.03546f
C489 VP.n45 GND 0.310084f
C490 VP.n46 GND 0.02015f
C491 VP.n47 GND 0.019809f
C492 VP.n48 GND 0.019809f
C493 VP.n49 GND 0.019809f
C494 VP.n50 GND 0.036919f
C495 VP.n51 GND 0.036919f
C496 VP.n52 GND 0.036919f
C497 VP.n53 GND 0.019809f
C498 VP.n54 GND 0.019809f
C499 VP.n55 GND 0.019809f
C500 VP.n56 GND 0.011536f
C501 VP.n57 GND 0.033611f
C502 VP.n58 GND 0.036919f
C503 VP.n59 GND 0.019809f
C504 VP.n60 GND 0.019809f
C505 VP.n61 GND 0.019809f
C506 VP.n62 GND 0.036919f
C507 VP.n63 GND 0.036919f
C508 VP.t10 GND 0.775277f
C509 VP.n64 GND 0.310084f
C510 VP.n65 GND 0.02015f
C511 VP.n66 GND 0.019809f
C512 VP.n67 GND 0.019809f
C513 VP.n68 GND 0.019809f
C514 VP.n69 GND 0.036919f
C515 VP.n70 GND 0.036919f
C516 VP.n71 GND 0.036919f
C517 VP.n72 GND 0.019809f
C518 VP.n73 GND 0.019809f
C519 VP.n74 GND 0.019809f
C520 VP.n75 GND 0.012146f
C521 VP.n76 GND 0.029693f
C522 VP.n77 GND 0.036919f
C523 VP.n78 GND 0.019809f
C524 VP.n79 GND 0.019809f
C525 VP.n80 GND 0.019809f
C526 VP.n81 GND 0.036919f
C527 VP.n82 GND 0.036919f
C528 VP.t5 GND 0.775277f
C529 VP.n83 GND 0.310084f
C530 VP.n84 GND 0.023066f
C531 VP.n85 GND 0.019809f
C532 VP.n86 GND 0.019809f
C533 VP.n87 GND 0.019809f
C534 VP.n88 GND 0.036919f
C535 VP.n89 GND 0.036919f
C536 VP.n90 GND 0.036919f
C537 VP.n91 GND 0.019809f
C538 VP.n92 GND 0.019809f
C539 VP.n93 GND 0.019809f
C540 VP.n94 GND 0.014127f
C541 VP.n95 GND 0.025362f
C542 VP.n96 GND 0.036919f
C543 VP.n97 GND 0.019809f
C544 VP.n98 GND 0.019809f
C545 VP.n99 GND 0.019809f
C546 VP.n100 GND 0.036919f
C547 VP.n101 GND 0.036919f
C548 VP.n102 GND 0.025983f
C549 VP.n103 GND 0.041916f
C550 VP.n104 GND 0.443801f
C551 VP.t3 GND 0.775277f
C552 VP.n105 GND 0.393512f
C553 VP.n106 GND 0.019809f
C554 VP.n107 GND 0.036919f
C555 VP.n108 GND 0.019809f
C556 VP.n109 GND 0.039269f
C557 VP.n110 GND 0.019809f
C558 VP.n111 GND 0.032544f
C559 VP.n112 GND 0.019809f
C560 VP.t9 GND 0.775277f
C561 VP.n113 GND 0.310084f
C562 VP.n114 GND 0.036919f
C563 VP.n115 GND 0.019809f
C564 VP.n116 GND 0.036919f
C565 VP.n117 GND 0.019809f
C566 VP.n118 GND 0.03546f
C567 VP.n119 GND 0.019809f
C568 VP.t6 GND 0.775277f
C569 VP.n120 GND 0.310084f
C570 VP.n121 GND 0.036919f
C571 VP.n122 GND 0.019809f
C572 VP.n123 GND 0.033611f
C573 VP.n124 GND 0.019809f
C574 VP.n125 GND 0.036919f
C575 VP.n126 GND 0.019809f
C576 VP.t1 GND 0.775277f
C577 VP.n127 GND 0.036919f
C578 VP.n128 GND 0.019809f
C579 VP.n129 GND 0.029693f
C580 VP.n130 GND 0.019809f
C581 VP.n131 GND 0.036919f
C582 VP.t7 GND 1.1317f
C583 VP.n132 GND 0.590385f
C584 VP.t2 GND 0.775277f
C585 VP.n133 GND 0.385367f
C586 VP.n134 GND 0.023066f
C587 VP.n135 GND 0.23314f
C588 VP.n136 GND 0.019809f
C589 VP.n137 GND 0.019809f
C590 VP.n138 GND 0.036919f
C591 VP.n139 GND 0.036919f
C592 VP.n140 GND 0.036919f
C593 VP.n141 GND 0.019809f
C594 VP.n142 GND 0.019809f
C595 VP.n143 GND 0.019809f
C596 VP.n144 GND 0.012146f
C597 VP.n145 GND 0.036919f
C598 VP.n146 GND 0.036919f
C599 VP.n147 GND 0.019809f
C600 VP.n148 GND 0.019809f
C601 VP.n149 GND 0.019809f
C602 VP.n150 GND 0.036919f
C603 VP.n151 GND 0.03546f
C604 VP.n152 GND 0.310084f
C605 VP.n153 GND 0.02015f
C606 VP.n154 GND 0.019809f
C607 VP.n155 GND 0.019809f
C608 VP.n156 GND 0.019809f
C609 VP.n157 GND 0.036919f
C610 VP.n158 GND 0.036919f
C611 VP.n159 GND 0.036919f
C612 VP.n160 GND 0.019809f
C613 VP.n161 GND 0.019809f
C614 VP.n162 GND 0.019809f
C615 VP.n163 GND 0.011536f
C616 VP.n164 GND 0.033611f
C617 VP.n165 GND 0.036919f
C618 VP.n166 GND 0.019809f
C619 VP.n167 GND 0.019809f
C620 VP.n168 GND 0.019809f
C621 VP.n169 GND 0.036919f
C622 VP.n170 GND 0.036919f
C623 VP.n171 GND 0.02015f
C624 VP.n172 GND 0.019809f
C625 VP.n173 GND 0.019809f
C626 VP.n174 GND 0.019809f
C627 VP.n175 GND 0.036919f
C628 VP.n176 GND 0.036919f
C629 VP.n177 GND 0.036919f
C630 VP.n178 GND 0.019809f
C631 VP.n179 GND 0.019809f
C632 VP.n180 GND 0.019809f
C633 VP.n181 GND 0.012146f
C634 VP.n182 GND 0.029693f
C635 VP.n183 GND 0.036919f
C636 VP.n184 GND 0.019809f
C637 VP.n185 GND 0.019809f
C638 VP.n186 GND 0.019809f
C639 VP.n187 GND 0.036919f
C640 VP.n188 GND 0.036919f
C641 VP.n189 GND 0.023066f
C642 VP.n190 GND 0.019809f
C643 VP.n191 GND 0.019809f
C644 VP.n192 GND 0.019809f
C645 VP.n193 GND 0.036919f
C646 VP.n194 GND 0.036919f
C647 VP.n195 GND 0.036919f
C648 VP.n196 GND 0.019809f
C649 VP.n197 GND 0.019809f
C650 VP.n198 GND 0.019809f
C651 VP.n199 GND 0.014127f
C652 VP.n200 GND 0.025362f
C653 VP.n201 GND 0.036919f
C654 VP.n202 GND 0.019809f
C655 VP.n203 GND 0.019809f
C656 VP.n204 GND 0.019809f
C657 VP.n205 GND 0.036919f
C658 VP.n206 GND 0.036919f
C659 VP.n207 GND 0.025983f
C660 VP.n208 GND 0.041916f
C661 VP.n209 GND 1.53053f
C662 VP.n210 GND 3.37409f
C663 VDD.t99 GND 0.011185f
C664 VDD.t77 GND 0.011185f
C665 VDD.n0 GND 0.051477f
C666 VDD.t70 GND 0.011185f
C667 VDD.t80 GND 0.011185f
C668 VDD.n1 GND 0.046609f
C669 VDD.n2 GND 0.924719f
C670 VDD.t85 GND 0.011185f
C671 VDD.t97 GND 0.011185f
C672 VDD.n3 GND 0.046609f
C673 VDD.n4 GND 0.484675f
C674 VDD.t72 GND 0.011185f
C675 VDD.t82 GND 0.011185f
C676 VDD.n5 GND 0.046609f
C677 VDD.n6 GND 0.399546f
C678 VDD.t103 GND 0.011185f
C679 VDD.t87 GND 0.011185f
C680 VDD.n7 GND 0.051477f
C681 VDD.t106 GND 0.011185f
C682 VDD.t89 GND 0.011185f
C683 VDD.n8 GND 0.046609f
C684 VDD.n9 GND 0.924718f
C685 VDD.t75 GND 0.011185f
C686 VDD.t101 GND 0.011185f
C687 VDD.n10 GND 0.046609f
C688 VDD.n11 GND 0.484675f
C689 VDD.t94 GND 0.011185f
C690 VDD.t108 GND 0.011185f
C691 VDD.n12 GND 0.046609f
C692 VDD.n13 GND 0.399546f
C693 VDD.n14 GND 0.299267f
C694 VDD.n15 GND 2.74383f
C695 VDD.t2 GND 0.116461f
C696 VDD.t9 GND 0.113326f
C697 VDD.n16 GND 0.538609f
C698 VDD.t7 GND 0.116461f
C699 VDD.t11 GND 0.113326f
C700 VDD.n17 GND 0.518679f
C701 VDD.n18 GND 0.445762f
C702 VDD.n19 GND 0.005135f
C703 VDD.n20 GND 0.006681f
C704 VDD.n21 GND 0.005377f
C705 VDD.n22 GND 0.006681f
C706 VDD.n23 GND 0.005377f
C707 VDD.n24 GND 0.006681f
C708 VDD.n25 GND 0.391723f
C709 VDD.n26 GND 0.006681f
C710 VDD.n27 GND 0.006681f
C711 VDD.n28 GND 0.006681f
C712 VDD.n29 GND 0.248744f
C713 VDD.n30 GND 0.006681f
C714 VDD.n31 GND 0.006681f
C715 VDD.n32 GND 0.006681f
C716 VDD.n33 GND 0.006681f
C717 VDD.n34 GND 0.006681f
C718 VDD.n35 GND 0.005377f
C719 VDD.n36 GND 0.006681f
C720 VDD.t8 GND 0.195862f
C721 VDD.n37 GND 0.006681f
C722 VDD.n38 GND 0.006681f
C723 VDD.n39 GND 0.006681f
C724 VDD.n40 GND 0.391723f
C725 VDD.n41 GND 0.006681f
C726 VDD.n42 GND 0.006681f
C727 VDD.n43 GND 0.006681f
C728 VDD.n44 GND 0.006681f
C729 VDD.n45 GND 0.006681f
C730 VDD.n46 GND 0.005377f
C731 VDD.n47 GND 0.006681f
C732 VDD.n48 GND 0.006681f
C733 VDD.n49 GND 0.006681f
C734 VDD.n50 GND 0.006681f
C735 VDD.n51 GND 0.391723f
C736 VDD.n52 GND 0.006681f
C737 VDD.n53 GND 0.006681f
C738 VDD.n54 GND 0.006681f
C739 VDD.n55 GND 0.006681f
C740 VDD.n56 GND 0.006681f
C741 VDD.n57 GND 0.005377f
C742 VDD.n58 GND 0.006681f
C743 VDD.n59 GND 0.006681f
C744 VDD.n60 GND 0.006681f
C745 VDD.n61 GND 0.006681f
C746 VDD.n62 GND 0.323172f
C747 VDD.n63 GND 0.006681f
C748 VDD.n64 GND 0.006681f
C749 VDD.n65 GND 0.006681f
C750 VDD.n66 GND 0.006681f
C751 VDD.n67 GND 0.006681f
C752 VDD.n68 GND 0.005377f
C753 VDD.n69 GND 0.006681f
C754 VDD.t13 GND 0.195862f
C755 VDD.n70 GND 0.006681f
C756 VDD.n71 GND 0.006681f
C757 VDD.n72 GND 0.006681f
C758 VDD.n73 GND 0.391723f
C759 VDD.n74 GND 0.006681f
C760 VDD.n75 GND 0.006681f
C761 VDD.n76 GND 0.006681f
C762 VDD.n77 GND 0.006681f
C763 VDD.n78 GND 0.006681f
C764 VDD.n79 GND 0.004463f
C765 VDD.n80 GND 0.014921f
C766 VDD.n81 GND 0.006681f
C767 VDD.n82 GND 0.014921f
C768 VDD.n96 GND 0.006681f
C769 VDD.t57 GND 0.141206f
C770 VDD.t56 GND 0.493991f
C771 VDD.n97 GND 0.092067f
C772 VDD.t58 GND 0.102298f
C773 VDD.n98 GND 0.095951f
C774 VDD.n99 GND 0.010082f
C775 VDD.n100 GND 0.006681f
C776 VDD.n101 GND 0.005377f
C777 VDD.n102 GND 0.006681f
C778 VDD.n103 GND 0.005377f
C779 VDD.n104 GND 0.006681f
C780 VDD.n105 GND 0.005377f
C781 VDD.n106 GND 0.006681f
C782 VDD.t14 GND 0.141206f
C783 VDD.t12 GND 0.493991f
C784 VDD.n107 GND 0.092067f
C785 VDD.t15 GND 0.102298f
C786 VDD.n108 GND 0.095951f
C787 VDD.n109 GND 0.006681f
C788 VDD.n110 GND 0.005377f
C789 VDD.n111 GND 0.006681f
C790 VDD.n112 GND 0.005377f
C791 VDD.n113 GND 0.006681f
C792 VDD.n114 GND 0.005377f
C793 VDD.n115 GND 0.014921f
C794 VDD.n116 GND 0.015143f
C795 VDD.n117 GND 0.015143f
C796 VDD.n118 GND 0.004463f
C797 VDD.n119 GND 0.006681f
C798 VDD.n120 GND 0.006681f
C799 VDD.n121 GND 0.005377f
C800 VDD.n122 GND 0.006681f
C801 VDD.n123 GND 0.006681f
C802 VDD.n124 GND 0.006681f
C803 VDD.n125 GND 0.005377f
C804 VDD.n126 GND 0.006681f
C805 VDD.n127 GND 0.006681f
C806 VDD.n128 GND 0.005377f
C807 VDD.n129 GND 0.006681f
C808 VDD.n130 GND 0.006681f
C809 VDD.n131 GND 0.005377f
C810 VDD.n132 GND 0.006681f
C811 VDD.n133 GND 0.006681f
C812 VDD.n134 GND 0.006681f
C813 VDD.n135 GND 0.005377f
C814 VDD.n136 GND 0.006681f
C815 VDD.n137 GND 0.006681f
C816 VDD.n138 GND 0.005377f
C817 VDD.n139 GND 0.006681f
C818 VDD.n140 GND 0.006681f
C819 VDD.n141 GND 0.005377f
C820 VDD.n142 GND 0.006681f
C821 VDD.n143 GND 0.006681f
C822 VDD.n144 GND 0.006681f
C823 VDD.n145 GND 0.006681f
C824 VDD.n146 GND 0.00406f
C825 VDD.n147 GND 0.010082f
C826 VDD.n148 GND 0.006681f
C827 VDD.n149 GND 0.006681f
C828 VDD.n150 GND 0.00492f
C829 VDD.n151 GND 0.006681f
C830 VDD.n152 GND 0.006681f
C831 VDD.n153 GND 0.006681f
C832 VDD.n154 GND 0.005377f
C833 VDD.n155 GND 0.006681f
C834 VDD.n156 GND 0.006681f
C835 VDD.n157 GND 0.005377f
C836 VDD.n158 GND 0.006681f
C837 VDD.n159 GND 0.006681f
C838 VDD.n160 GND 0.005377f
C839 VDD.n161 GND 0.006681f
C840 VDD.n162 GND 0.006681f
C841 VDD.n163 GND 0.006681f
C842 VDD.n164 GND 0.005377f
C843 VDD.n165 GND 0.006681f
C844 VDD.n166 GND 0.006681f
C845 VDD.n167 GND 0.005377f
C846 VDD.n168 GND 0.006681f
C847 VDD.n169 GND 0.006681f
C848 VDD.n170 GND 0.005377f
C849 VDD.n171 GND 0.006681f
C850 VDD.n172 GND 0.006681f
C851 VDD.n173 GND 0.006681f
C852 VDD.n174 GND 0.005377f
C853 VDD.n175 GND 0.006681f
C854 VDD.n176 GND 0.006681f
C855 VDD.n177 GND 0.005377f
C856 VDD.n178 GND 0.006681f
C857 VDD.n179 GND 0.005243f
C858 VDD.n180 GND 0.006681f
C859 VDD.n181 GND 0.006681f
C860 VDD.n182 GND 0.006681f
C861 VDD.n183 GND 0.005377f
C862 VDD.n184 GND 0.006681f
C863 VDD.n185 GND 0.005377f
C864 VDD.n186 GND 0.006681f
C865 VDD.n187 GND 0.005377f
C866 VDD.n188 GND 0.006681f
C867 VDD.n189 GND 0.005377f
C868 VDD.n190 GND 0.006681f
C869 VDD.n191 GND 0.005377f
C870 VDD.n192 GND 0.006681f
C871 VDD.n193 GND 0.005377f
C872 VDD.n194 GND 0.006681f
C873 VDD.n195 GND 0.006681f
C874 VDD.n196 GND 0.391723f
C875 VDD.n197 GND 0.006681f
C876 VDD.n198 GND 0.005377f
C877 VDD.n199 GND 0.006681f
C878 VDD.n200 GND 0.005377f
C879 VDD.n201 GND 0.006681f
C880 VDD.n202 GND 0.248744f
C881 VDD.n203 GND 0.006681f
C882 VDD.n204 GND 0.005377f
C883 VDD.n205 GND 0.006681f
C884 VDD.n206 GND 0.005377f
C885 VDD.n207 GND 0.006681f
C886 VDD.n208 GND 0.391723f
C887 VDD.t1 GND 0.195862f
C888 VDD.n209 GND 0.006681f
C889 VDD.n210 GND 0.005377f
C890 VDD.n211 GND 0.006681f
C891 VDD.n212 GND 0.005377f
C892 VDD.n213 GND 0.006681f
C893 VDD.n214 GND 0.391723f
C894 VDD.n215 GND 0.006681f
C895 VDD.n216 GND 0.005377f
C896 VDD.n217 GND 0.006681f
C897 VDD.n218 GND 0.005377f
C898 VDD.n219 GND 0.006681f
C899 VDD.n220 GND 0.391723f
C900 VDD.n221 GND 0.006681f
C901 VDD.n222 GND 0.005377f
C902 VDD.n223 GND 0.006681f
C903 VDD.n224 GND 0.005377f
C904 VDD.n225 GND 0.006681f
C905 VDD.n226 GND 0.391723f
C906 VDD.n227 GND 0.006681f
C907 VDD.n228 GND 0.005377f
C908 VDD.n229 GND 0.006681f
C909 VDD.n230 GND 0.005377f
C910 VDD.n231 GND 0.006681f
C911 VDD.n232 GND 0.391723f
C912 VDD.n233 GND 0.006681f
C913 VDD.n234 GND 0.005377f
C914 VDD.n235 GND 0.006681f
C915 VDD.n236 GND 0.005377f
C916 VDD.n237 GND 0.006681f
C917 VDD.n238 GND 0.323172f
C918 VDD.n239 GND 0.006681f
C919 VDD.n240 GND 0.005377f
C920 VDD.n241 GND 0.006681f
C921 VDD.n242 GND 0.005377f
C922 VDD.n243 GND 0.006681f
C923 VDD.n244 GND 0.391723f
C924 VDD.t50 GND 0.195862f
C925 VDD.n245 GND 0.006681f
C926 VDD.n246 GND 0.005377f
C927 VDD.n247 GND 0.006681f
C928 VDD.n248 GND 0.005377f
C929 VDD.n249 GND 0.006681f
C930 VDD.n250 GND 0.391723f
C931 VDD.n251 GND 0.006681f
C932 VDD.n252 GND 0.005377f
C933 VDD.n253 GND 0.007549f
C934 VDD.n254 GND 0.004463f
C935 VDD.n255 GND 0.014921f
C936 VDD.n256 GND 0.522951f
C937 VDD.n257 GND 0.014921f
C938 VDD.n258 GND 0.004463f
C939 VDD.n259 GND 0.051977f
C940 VDD.n260 GND 0.113416f
C941 VDD.n261 GND 0.00334f
C942 VDD.n262 GND 0.005377f
C943 VDD.n263 GND 0.006681f
C944 VDD.t0 GND 6.05017f
C945 VDD.n276 GND 0.015143f
C946 VDD.n277 GND 0.006681f
C947 VDD.n278 GND 0.00334f
C948 VDD.n279 GND 0.00334f
C949 VDD.n280 GND 0.00334f
C950 VDD.n281 GND 0.00334f
C951 VDD.n282 GND 0.00334f
C952 VDD.n283 GND 0.00334f
C953 VDD.n284 GND 0.00334f
C954 VDD.n285 GND 0.00334f
C955 VDD.n286 GND 0.00334f
C956 VDD.n287 GND 0.00334f
C957 VDD.n288 GND 0.006681f
C958 VDD.n289 GND 0.00334f
C959 VDD.t64 GND 0.141206f
C960 VDD.t62 GND 0.493991f
C961 VDD.n290 GND 0.092067f
C962 VDD.t63 GND 0.102298f
C963 VDD.n291 GND 0.095951f
C964 VDD.n292 GND 0.002505f
C965 VDD.n293 GND 0.002505f
C966 VDD.n294 GND 0.00334f
C967 VDD.n295 GND 0.00334f
C968 VDD.n296 GND 0.00334f
C969 VDD.n297 GND 0.00334f
C970 VDD.n298 GND 0.00334f
C971 VDD.n299 GND 0.00334f
C972 VDD.n300 GND 0.00334f
C973 VDD.n301 GND 0.00334f
C974 VDD.n302 GND 0.00334f
C975 VDD.n303 GND 0.00334f
C976 VDD.n304 GND 0.006681f
C977 VDD.t52 GND 0.141206f
C978 VDD.t49 GND 0.493991f
C979 VDD.n305 GND 0.092067f
C980 VDD.t51 GND 0.102298f
C981 VDD.n306 GND 0.095951f
C982 VDD.n307 GND 0.010082f
C983 VDD.n308 GND 0.003407f
C984 VDD.n309 GND 0.004543f
C985 VDD.n310 GND 0.004543f
C986 VDD.t86 GND 5.59381f
C987 VDD.t102 GND 3.64107f
C988 VDD.n311 GND 1.3632f
C989 VDD.n312 GND 0.004543f
C990 VDD.n313 GND 0.004543f
C991 VDD.t41 GND 0.077008f
C992 VDD.t40 GND 0.389773f
C993 VDD.n314 GND 0.080451f
C994 VDD.t42 GND 0.047872f
C995 VDD.n315 GND 0.076995f
C996 VDD.n316 GND 0.004543f
C997 VDD.n318 GND 0.010421f
C998 VDD.n319 GND 0.004543f
C999 VDD.n320 GND 0.004543f
C1000 VDD.n321 GND 0.266372f
C1001 VDD.n322 GND 0.004543f
C1002 VDD.n323 GND 0.374096f
C1003 VDD.n324 GND 0.004543f
C1004 VDD.n325 GND 0.004543f
C1005 VDD.n326 GND 0.010421f
C1006 VDD.n327 GND 0.004543f
C1007 VDD.n328 GND 0.004543f
C1008 VDD.n329 GND 0.004543f
C1009 VDD.n330 GND 0.004543f
C1010 VDD.n331 GND 0.004543f
C1011 VDD.n333 GND 0.003407f
C1012 VDD.n334 GND 0.004543f
C1013 VDD.t22 GND 0.077008f
C1014 VDD.t20 GND 0.389773f
C1015 VDD.n335 GND 0.080451f
C1016 VDD.t23 GND 0.047872f
C1017 VDD.n336 GND 0.076995f
C1018 VDD.n337 GND 0.005605f
C1019 VDD.n339 GND 0.002773f
C1020 VDD.n340 GND 0.004543f
C1021 VDD.n341 GND 0.004543f
C1022 VDD.n342 GND 0.004543f
C1023 VDD.n343 GND 0.266372f
C1024 VDD.n344 GND 0.004543f
C1025 VDD.n345 GND 0.004543f
C1026 VDD.n346 GND 0.004543f
C1027 VDD.n347 GND 0.004543f
C1028 VDD.n348 GND 0.004543f
C1029 VDD.n349 GND 0.266372f
C1030 VDD.n350 GND 0.004543f
C1031 VDD.n351 GND 0.004543f
C1032 VDD.n352 GND 0.004543f
C1033 VDD.n353 GND 0.004543f
C1034 VDD.n354 GND 0.004543f
C1035 VDD.n355 GND 0.004543f
C1036 VDD.n356 GND 0.223282f
C1037 VDD.n357 GND 0.004543f
C1038 VDD.n358 GND 0.004543f
C1039 VDD.n359 GND 0.004543f
C1040 VDD.n360 GND 0.004543f
C1041 VDD.n361 GND 0.004543f
C1042 VDD.n362 GND 0.266372f
C1043 VDD.n363 GND 0.004543f
C1044 VDD.n364 GND 0.004543f
C1045 VDD.t88 GND 0.133186f
C1046 VDD.n365 GND 0.004543f
C1047 VDD.n366 GND 0.004543f
C1048 VDD.n367 GND 0.004543f
C1049 VDD.t21 GND 0.133186f
C1050 VDD.n368 GND 0.004543f
C1051 VDD.n369 GND 0.004543f
C1052 VDD.n370 GND 0.004543f
C1053 VDD.n371 GND 0.004543f
C1054 VDD.n372 GND 0.004543f
C1055 VDD.n373 GND 0.266372f
C1056 VDD.n374 GND 0.004543f
C1057 VDD.n375 GND 0.004543f
C1058 VDD.n376 GND 0.260496f
C1059 VDD.n377 GND 0.004543f
C1060 VDD.n378 GND 0.004543f
C1061 VDD.n379 GND 0.004543f
C1062 VDD.n380 GND 0.266372f
C1063 VDD.n381 GND 0.004543f
C1064 VDD.n382 GND 0.004543f
C1065 VDD.n383 GND 0.004543f
C1066 VDD.n384 GND 0.004543f
C1067 VDD.n385 GND 0.004543f
C1068 VDD.n386 GND 0.266372f
C1069 VDD.n387 GND 0.004543f
C1070 VDD.n388 GND 0.004543f
C1071 VDD.n389 GND 0.004543f
C1072 VDD.n390 GND 0.004543f
C1073 VDD.n391 GND 0.004543f
C1074 VDD.n392 GND 0.266372f
C1075 VDD.n393 GND 0.004543f
C1076 VDD.n394 GND 0.004543f
C1077 VDD.n395 GND 0.004543f
C1078 VDD.n396 GND 0.004543f
C1079 VDD.n397 GND 0.004543f
C1080 VDD.n398 GND 0.266372f
C1081 VDD.n399 GND 0.004543f
C1082 VDD.n400 GND 0.004543f
C1083 VDD.n401 GND 0.004543f
C1084 VDD.n402 GND 0.004543f
C1085 VDD.n403 GND 0.004543f
C1086 VDD.n404 GND 0.266372f
C1087 VDD.n405 GND 0.004543f
C1088 VDD.n406 GND 0.004543f
C1089 VDD.n407 GND 0.004543f
C1090 VDD.n408 GND 0.004543f
C1091 VDD.n409 GND 0.004543f
C1092 VDD.n410 GND 0.266372f
C1093 VDD.n411 GND 0.004543f
C1094 VDD.n412 GND 0.004543f
C1095 VDD.n413 GND 0.004543f
C1096 VDD.n414 GND 0.004543f
C1097 VDD.n415 GND 0.004543f
C1098 VDD.t105 GND 0.133186f
C1099 VDD.n416 GND 0.004543f
C1100 VDD.n417 GND 0.004543f
C1101 VDD.n418 GND 0.004543f
C1102 VDD.n419 GND 0.004543f
C1103 VDD.n420 GND 0.004543f
C1104 VDD.n421 GND 0.266372f
C1105 VDD.n422 GND 0.004543f
C1106 VDD.n423 GND 0.004543f
C1107 VDD.n424 GND 0.188027f
C1108 VDD.n425 GND 0.004543f
C1109 VDD.n426 GND 0.004543f
C1110 VDD.n427 GND 0.004543f
C1111 VDD.n428 GND 0.266372f
C1112 VDD.n429 GND 0.004543f
C1113 VDD.n430 GND 0.004543f
C1114 VDD.n431 GND 0.004543f
C1115 VDD.n432 GND 0.004543f
C1116 VDD.n433 GND 0.004543f
C1117 VDD.n434 GND 0.150813f
C1118 VDD.n435 GND 0.004543f
C1119 VDD.n436 GND 0.004543f
C1120 VDD.n437 GND 0.004543f
C1121 VDD.n438 GND 0.004543f
C1122 VDD.n439 GND 0.004543f
C1123 VDD.n440 GND 0.266372f
C1124 VDD.n441 GND 0.004543f
C1125 VDD.n442 GND 0.004543f
C1126 VDD.t90 GND 0.133186f
C1127 VDD.n443 GND 0.004543f
C1128 VDD.n444 GND 0.004543f
C1129 VDD.n445 GND 0.004543f
C1130 VDD.n446 GND 0.266372f
C1131 VDD.n447 GND 0.004543f
C1132 VDD.n448 GND 0.004543f
C1133 VDD.n449 GND 0.004543f
C1134 VDD.n450 GND 0.004543f
C1135 VDD.n451 GND 0.004543f
C1136 VDD.n452 GND 0.266372f
C1137 VDD.n453 GND 0.004543f
C1138 VDD.n454 GND 0.004543f
C1139 VDD.n455 GND 0.004543f
C1140 VDD.n456 GND 0.004543f
C1141 VDD.n457 GND 0.004543f
C1142 VDD.n458 GND 0.266372f
C1143 VDD.n459 GND 0.004543f
C1144 VDD.n460 GND 0.004543f
C1145 VDD.n461 GND 0.004543f
C1146 VDD.n462 GND 0.004543f
C1147 VDD.n463 GND 0.004543f
C1148 VDD.n464 GND 0.266372f
C1149 VDD.n465 GND 0.004543f
C1150 VDD.n466 GND 0.004543f
C1151 VDD.n467 GND 0.004543f
C1152 VDD.n468 GND 0.004543f
C1153 VDD.n469 GND 0.004543f
C1154 VDD.n470 GND 0.266372f
C1155 VDD.n471 GND 0.004543f
C1156 VDD.n472 GND 0.004543f
C1157 VDD.n473 GND 0.004543f
C1158 VDD.n474 GND 0.004543f
C1159 VDD.n475 GND 0.004543f
C1160 VDD.n476 GND 0.266372f
C1161 VDD.n477 GND 0.004543f
C1162 VDD.n478 GND 0.004543f
C1163 VDD.n479 GND 0.004543f
C1164 VDD.n480 GND 0.004543f
C1165 VDD.n481 GND 0.004543f
C1166 VDD.n482 GND 0.266372f
C1167 VDD.n483 GND 0.004543f
C1168 VDD.n484 GND 0.004543f
C1169 VDD.n485 GND 0.004543f
C1170 VDD.n486 GND 0.004543f
C1171 VDD.n487 GND 0.004543f
C1172 VDD.n488 GND 0.266372f
C1173 VDD.n489 GND 0.004543f
C1174 VDD.n490 GND 0.004543f
C1175 VDD.n491 GND 0.004543f
C1176 VDD.n492 GND 0.004543f
C1177 VDD.n493 GND 0.004543f
C1178 VDD.t91 GND 0.133186f
C1179 VDD.n494 GND 0.004543f
C1180 VDD.n495 GND 0.004543f
C1181 VDD.n496 GND 0.004543f
C1182 VDD.n497 GND 0.004543f
C1183 VDD.n498 GND 0.004543f
C1184 VDD.t100 GND 0.133186f
C1185 VDD.n499 GND 0.004543f
C1186 VDD.n500 GND 0.004543f
C1187 VDD.n501 GND 0.260496f
C1188 VDD.n502 GND 0.004543f
C1189 VDD.n503 GND 0.004543f
C1190 VDD.n504 GND 0.004543f
C1191 VDD.n505 GND 0.266372f
C1192 VDD.n506 GND 0.004543f
C1193 VDD.n507 GND 0.004543f
C1194 VDD.n508 GND 0.186069f
C1195 VDD.n509 GND 0.004543f
C1196 VDD.n510 GND 0.004543f
C1197 VDD.n511 GND 0.004543f
C1198 VDD.n512 GND 0.266372f
C1199 VDD.n513 GND 0.004543f
C1200 VDD.n514 GND 0.004543f
C1201 VDD.n515 GND 0.004543f
C1202 VDD.n516 GND 0.004543f
C1203 VDD.n517 GND 0.004543f
C1204 VDD.n518 GND 0.266372f
C1205 VDD.n519 GND 0.004543f
C1206 VDD.n520 GND 0.004543f
C1207 VDD.n521 GND 0.004543f
C1208 VDD.n522 GND 0.004543f
C1209 VDD.n523 GND 0.004543f
C1210 VDD.n524 GND 0.266372f
C1211 VDD.n525 GND 0.004543f
C1212 VDD.n526 GND 0.004543f
C1213 VDD.n527 GND 0.004543f
C1214 VDD.n528 GND 0.004543f
C1215 VDD.n529 GND 0.004543f
C1216 VDD.n530 GND 0.266372f
C1217 VDD.n531 GND 0.004543f
C1218 VDD.n532 GND 0.004543f
C1219 VDD.n533 GND 0.004543f
C1220 VDD.n534 GND 0.004543f
C1221 VDD.n535 GND 0.004543f
C1222 VDD.n536 GND 0.266372f
C1223 VDD.n537 GND 0.004543f
C1224 VDD.n538 GND 0.004543f
C1225 VDD.n539 GND 0.004543f
C1226 VDD.n540 GND 0.004543f
C1227 VDD.n541 GND 0.004543f
C1228 VDD.n542 GND 0.266372f
C1229 VDD.n543 GND 0.004543f
C1230 VDD.n544 GND 0.004543f
C1231 VDD.n545 GND 0.004543f
C1232 VDD.n546 GND 0.004543f
C1233 VDD.n547 GND 0.004543f
C1234 VDD.t78 GND 0.133186f
C1235 VDD.n548 GND 0.004543f
C1236 VDD.n549 GND 0.004543f
C1237 VDD.n550 GND 0.004543f
C1238 VDD.n551 GND 0.004543f
C1239 VDD.n552 GND 0.004543f
C1240 VDD.n553 GND 0.201738f
C1241 VDD.n554 GND 0.004543f
C1242 VDD.n555 GND 0.004543f
C1243 VDD.n556 GND 0.139062f
C1244 VDD.n557 GND 0.004543f
C1245 VDD.n558 GND 0.004543f
C1246 VDD.n559 GND 0.004543f
C1247 VDD.n560 GND 0.266372f
C1248 VDD.n561 GND 0.004543f
C1249 VDD.n562 GND 0.004543f
C1250 VDD.t74 GND 0.133186f
C1251 VDD.n563 GND 0.004543f
C1252 VDD.n564 GND 0.004543f
C1253 VDD.n565 GND 0.004543f
C1254 VDD.n566 GND 0.266372f
C1255 VDD.n567 GND 0.004543f
C1256 VDD.n568 GND 0.004543f
C1257 VDD.n569 GND 0.004543f
C1258 VDD.n570 GND 0.004543f
C1259 VDD.n571 GND 0.004543f
C1260 VDD.n572 GND 0.266372f
C1261 VDD.n573 GND 0.004543f
C1262 VDD.n574 GND 0.004543f
C1263 VDD.n575 GND 0.004543f
C1264 VDD.n576 GND 0.004543f
C1265 VDD.n577 GND 0.004543f
C1266 VDD.n578 GND 0.266372f
C1267 VDD.n579 GND 0.004543f
C1268 VDD.n580 GND 0.004543f
C1269 VDD.n581 GND 0.004543f
C1270 VDD.n582 GND 0.004543f
C1271 VDD.n583 GND 0.004543f
C1272 VDD.n584 GND 0.266372f
C1273 VDD.n585 GND 0.004543f
C1274 VDD.n586 GND 0.004543f
C1275 VDD.n587 GND 0.004543f
C1276 VDD.n588 GND 0.004543f
C1277 VDD.n589 GND 0.004543f
C1278 VDD.n590 GND 0.266372f
C1279 VDD.n591 GND 0.004543f
C1280 VDD.n592 GND 0.004543f
C1281 VDD.n593 GND 0.004543f
C1282 VDD.n594 GND 0.004543f
C1283 VDD.n595 GND 0.004543f
C1284 VDD.n596 GND 0.266372f
C1285 VDD.n597 GND 0.004543f
C1286 VDD.n598 GND 0.004543f
C1287 VDD.n599 GND 0.004543f
C1288 VDD.n600 GND 0.004543f
C1289 VDD.n601 GND 0.004543f
C1290 VDD.n602 GND 0.248744f
C1291 VDD.n603 GND 0.004543f
C1292 VDD.n604 GND 0.004543f
C1293 VDD.n605 GND 0.004543f
C1294 VDD.n606 GND 0.004543f
C1295 VDD.n607 GND 0.004543f
C1296 VDD.n608 GND 0.266372f
C1297 VDD.n609 GND 0.004543f
C1298 VDD.n610 GND 0.004543f
C1299 VDD.t92 GND 0.133186f
C1300 VDD.n611 GND 0.004543f
C1301 VDD.n612 GND 0.004543f
C1302 VDD.n613 GND 0.004543f
C1303 VDD.t107 GND 0.133186f
C1304 VDD.n614 GND 0.004543f
C1305 VDD.n615 GND 0.004543f
C1306 VDD.n616 GND 0.004543f
C1307 VDD.n617 GND 0.004543f
C1308 VDD.n618 GND 0.004543f
C1309 VDD.n619 GND 0.266372f
C1310 VDD.n620 GND 0.004543f
C1311 VDD.n621 GND 0.004543f
C1312 VDD.n622 GND 0.209572f
C1313 VDD.n623 GND 0.004543f
C1314 VDD.n624 GND 0.004543f
C1315 VDD.n625 GND 0.004543f
C1316 VDD.n626 GND 0.266372f
C1317 VDD.n627 GND 0.004543f
C1318 VDD.n628 GND 0.004543f
C1319 VDD.n629 GND 0.004543f
C1320 VDD.n630 GND 0.004543f
C1321 VDD.n631 GND 0.004543f
C1322 VDD.n632 GND 0.266372f
C1323 VDD.n633 GND 0.004543f
C1324 VDD.n634 GND 0.004543f
C1325 VDD.n635 GND 0.004543f
C1326 VDD.n636 GND 0.004543f
C1327 VDD.n637 GND 0.004543f
C1328 VDD.n638 GND 0.266372f
C1329 VDD.n639 GND 0.004543f
C1330 VDD.n640 GND 0.004543f
C1331 VDD.n641 GND 0.004543f
C1332 VDD.n642 GND 0.004543f
C1333 VDD.n643 GND 0.004543f
C1334 VDD.n644 GND 0.266372f
C1335 VDD.n645 GND 0.004543f
C1336 VDD.n646 GND 0.004543f
C1337 VDD.n647 GND 0.004543f
C1338 VDD.n648 GND 0.004543f
C1339 VDD.n649 GND 0.004543f
C1340 VDD.n650 GND 0.266372f
C1341 VDD.n651 GND 0.004543f
C1342 VDD.n652 GND 0.004543f
C1343 VDD.n653 GND 0.004543f
C1344 VDD.n654 GND 0.004543f
C1345 VDD.n655 GND 0.004543f
C1346 VDD.n656 GND 0.266372f
C1347 VDD.n657 GND 0.004543f
C1348 VDD.n658 GND 0.004543f
C1349 VDD.n659 GND 0.004543f
C1350 VDD.n660 GND 0.004543f
C1351 VDD.n661 GND 0.004543f
C1352 VDD.n662 GND 0.266372f
C1353 VDD.n663 GND 0.004543f
C1354 VDD.n664 GND 0.004543f
C1355 VDD.n665 GND 0.004543f
C1356 VDD.n666 GND 0.004543f
C1357 VDD.n667 GND 0.004543f
C1358 VDD.n668 GND 0.178234f
C1359 VDD.n669 GND 0.004543f
C1360 VDD.n670 GND 0.004543f
C1361 VDD.n671 GND 0.004543f
C1362 VDD.n672 GND 0.004543f
C1363 VDD.n673 GND 0.004543f
C1364 VDD.t33 GND 0.133186f
C1365 VDD.n674 GND 0.004543f
C1366 VDD.n675 GND 0.004543f
C1367 VDD.t93 GND 0.133186f
C1368 VDD.n676 GND 0.004543f
C1369 VDD.n677 GND 0.004543f
C1370 VDD.n678 GND 0.004543f
C1371 VDD.n679 GND 0.266372f
C1372 VDD.n680 GND 0.004543f
C1373 VDD.n681 GND 0.004543f
C1374 VDD.n682 GND 0.139062f
C1375 VDD.n683 GND 0.004543f
C1376 VDD.n684 GND 0.004543f
C1377 VDD.n685 GND 0.004543f
C1378 VDD.n686 GND 0.266372f
C1379 VDD.n687 GND 0.004543f
C1380 VDD.n688 GND 0.004543f
C1381 VDD.n689 GND 0.004543f
C1382 VDD.n690 GND 0.004543f
C1383 VDD.n691 GND 0.004543f
C1384 VDD.n692 GND 0.266372f
C1385 VDD.n693 GND 0.004543f
C1386 VDD.n694 GND 0.004543f
C1387 VDD.n695 GND 0.004543f
C1388 VDD.n696 GND 0.004543f
C1389 VDD.n697 GND 0.004543f
C1390 VDD.n698 GND 0.266372f
C1391 VDD.n699 GND 0.004543f
C1392 VDD.n700 GND 0.004543f
C1393 VDD.n701 GND 0.004543f
C1394 VDD.n702 GND 0.004543f
C1395 VDD.n703 GND 0.004543f
C1396 VDD.n704 GND 0.266372f
C1397 VDD.n705 GND 0.004543f
C1398 VDD.n706 GND 0.004543f
C1399 VDD.n707 GND 0.004543f
C1400 VDD.n708 GND 0.010891f
C1401 VDD.n709 GND 0.010891f
C1402 VDD.n710 GND 0.374096f
C1403 VDD.n726 GND 0.004543f
C1404 VDD.n727 GND 0.010421f
C1405 VDD.n728 GND 0.004543f
C1406 VDD.n729 GND 0.004543f
C1407 VDD.n730 GND 0.004543f
C1408 VDD.n731 GND 0.266372f
C1409 VDD.n732 GND 0.004543f
C1410 VDD.n733 GND 0.004543f
C1411 VDD.n734 GND 0.004543f
C1412 VDD.n735 GND 0.010421f
C1413 VDD.n736 GND 0.004543f
C1414 VDD.t60 GND 0.077008f
C1415 VDD.t59 GND 0.389773f
C1416 VDD.n737 GND 0.080451f
C1417 VDD.t61 GND 0.047872f
C1418 VDD.n738 GND 0.076995f
C1419 VDD.n739 GND 0.005605f
C1420 VDD.n740 GND 0.004543f
C1421 VDD.n741 GND 0.004543f
C1422 VDD.n742 GND 0.266372f
C1423 VDD.n743 GND 0.004543f
C1424 VDD.n744 GND 0.004543f
C1425 VDD.n745 GND 0.004543f
C1426 VDD.n746 GND 0.004543f
C1427 VDD.n747 GND 0.004543f
C1428 VDD.n748 GND 0.266372f
C1429 VDD.n749 GND 0.004543f
C1430 VDD.n750 GND 0.004543f
C1431 VDD.n751 GND 0.004543f
C1432 VDD.n752 GND 0.004543f
C1433 VDD.n753 GND 0.004543f
C1434 VDD.n754 GND 0.004543f
C1435 VDD.n755 GND 0.266372f
C1436 VDD.n756 GND 0.004543f
C1437 VDD.n757 GND 0.004543f
C1438 VDD.n758 GND 0.004543f
C1439 VDD.n759 GND 0.004543f
C1440 VDD.n760 GND 0.004543f
C1441 VDD.n761 GND 0.266372f
C1442 VDD.n762 GND 0.004543f
C1443 VDD.n763 GND 0.004543f
C1444 VDD.n764 GND 0.004543f
C1445 VDD.n765 GND 0.004543f
C1446 VDD.n766 GND 0.004543f
C1447 VDD.t17 GND 0.133186f
C1448 VDD.n767 GND 0.004543f
C1449 VDD.n768 GND 0.004543f
C1450 VDD.n769 GND 0.004543f
C1451 VDD.n770 GND 0.004543f
C1452 VDD.n771 GND 0.004543f
C1453 VDD.n772 GND 0.266372f
C1454 VDD.n773 GND 0.004543f
C1455 VDD.n774 GND 0.004543f
C1456 VDD.t81 GND 0.133186f
C1457 VDD.n775 GND 0.004543f
C1458 VDD.n776 GND 0.004543f
C1459 VDD.n777 GND 0.004543f
C1460 VDD.n778 GND 0.266372f
C1461 VDD.n779 GND 0.004543f
C1462 VDD.n780 GND 0.004543f
C1463 VDD.n781 GND 0.004543f
C1464 VDD.n782 GND 0.004543f
C1465 VDD.n783 GND 0.004543f
C1466 VDD.n784 GND 0.266372f
C1467 VDD.n785 GND 0.004543f
C1468 VDD.n786 GND 0.004543f
C1469 VDD.n787 GND 0.004543f
C1470 VDD.n788 GND 0.004543f
C1471 VDD.n789 GND 0.004543f
C1472 VDD.n790 GND 0.266372f
C1473 VDD.n791 GND 0.004543f
C1474 VDD.n792 GND 0.004543f
C1475 VDD.n793 GND 0.004543f
C1476 VDD.n794 GND 0.004543f
C1477 VDD.n795 GND 0.004543f
C1478 VDD.n796 GND 0.266372f
C1479 VDD.n797 GND 0.004543f
C1480 VDD.n798 GND 0.004543f
C1481 VDD.n799 GND 0.004543f
C1482 VDD.n800 GND 0.004543f
C1483 VDD.n801 GND 0.004543f
C1484 VDD.n802 GND 0.266372f
C1485 VDD.n803 GND 0.004543f
C1486 VDD.n804 GND 0.004543f
C1487 VDD.n805 GND 0.004543f
C1488 VDD.n806 GND 0.004543f
C1489 VDD.n807 GND 0.004543f
C1490 VDD.n808 GND 0.266372f
C1491 VDD.n809 GND 0.004543f
C1492 VDD.n810 GND 0.004543f
C1493 VDD.n811 GND 0.004543f
C1494 VDD.n812 GND 0.004543f
C1495 VDD.n813 GND 0.004543f
C1496 VDD.n814 GND 0.266372f
C1497 VDD.n815 GND 0.004543f
C1498 VDD.n816 GND 0.004543f
C1499 VDD.n817 GND 0.004543f
C1500 VDD.n818 GND 0.004543f
C1501 VDD.n819 GND 0.004543f
C1502 VDD.n820 GND 0.266372f
C1503 VDD.n821 GND 0.004543f
C1504 VDD.n822 GND 0.004543f
C1505 VDD.n823 GND 0.004543f
C1506 VDD.n824 GND 0.004543f
C1507 VDD.n825 GND 0.004543f
C1508 VDD.t71 GND 0.133186f
C1509 VDD.n826 GND 0.004543f
C1510 VDD.n827 GND 0.004543f
C1511 VDD.n828 GND 0.004543f
C1512 VDD.n829 GND 0.004543f
C1513 VDD.n830 GND 0.004543f
C1514 VDD.n831 GND 0.150813f
C1515 VDD.n832 GND 0.004543f
C1516 VDD.n833 GND 0.004543f
C1517 VDD.n834 GND 0.189986f
C1518 VDD.n835 GND 0.004543f
C1519 VDD.n836 GND 0.004543f
C1520 VDD.n837 GND 0.004543f
C1521 VDD.n838 GND 0.266372f
C1522 VDD.n839 GND 0.004543f
C1523 VDD.n840 GND 0.004543f
C1524 VDD.t104 GND 0.133186f
C1525 VDD.n841 GND 0.004543f
C1526 VDD.n842 GND 0.004543f
C1527 VDD.n843 GND 0.004543f
C1528 VDD.n844 GND 0.266372f
C1529 VDD.n845 GND 0.004543f
C1530 VDD.n846 GND 0.004543f
C1531 VDD.n847 GND 0.004543f
C1532 VDD.n848 GND 0.004543f
C1533 VDD.n849 GND 0.004543f
C1534 VDD.n850 GND 0.266372f
C1535 VDD.n851 GND 0.004543f
C1536 VDD.n852 GND 0.004543f
C1537 VDD.n853 GND 0.004543f
C1538 VDD.n854 GND 0.004543f
C1539 VDD.n855 GND 0.004543f
C1540 VDD.n856 GND 0.266372f
C1541 VDD.n857 GND 0.004543f
C1542 VDD.n858 GND 0.004543f
C1543 VDD.n859 GND 0.004543f
C1544 VDD.n860 GND 0.004543f
C1545 VDD.n861 GND 0.004543f
C1546 VDD.n862 GND 0.266372f
C1547 VDD.n863 GND 0.004543f
C1548 VDD.n864 GND 0.004543f
C1549 VDD.n865 GND 0.004543f
C1550 VDD.n866 GND 0.004543f
C1551 VDD.n867 GND 0.004543f
C1552 VDD.n868 GND 0.266372f
C1553 VDD.n869 GND 0.004543f
C1554 VDD.n870 GND 0.004543f
C1555 VDD.n871 GND 0.004543f
C1556 VDD.n872 GND 0.004543f
C1557 VDD.n873 GND 0.004543f
C1558 VDD.n874 GND 0.266372f
C1559 VDD.n875 GND 0.004543f
C1560 VDD.n876 GND 0.004543f
C1561 VDD.n877 GND 0.004543f
C1562 VDD.n878 GND 0.004543f
C1563 VDD.n879 GND 0.004543f
C1564 VDD.n880 GND 0.19782f
C1565 VDD.n881 GND 0.004543f
C1566 VDD.n882 GND 0.004543f
C1567 VDD.n883 GND 0.004543f
C1568 VDD.n884 GND 0.004543f
C1569 VDD.n885 GND 0.004543f
C1570 VDD.n886 GND 0.266372f
C1571 VDD.n887 GND 0.004543f
C1572 VDD.n888 GND 0.004543f
C1573 VDD.t96 GND 0.133186f
C1574 VDD.n889 GND 0.004543f
C1575 VDD.n890 GND 0.004543f
C1576 VDD.n891 GND 0.004543f
C1577 VDD.t95 GND 0.133186f
C1578 VDD.n892 GND 0.004543f
C1579 VDD.n893 GND 0.004543f
C1580 VDD.n894 GND 0.004543f
C1581 VDD.n895 GND 0.004543f
C1582 VDD.n896 GND 0.004543f
C1583 VDD.n897 GND 0.266372f
C1584 VDD.n898 GND 0.004543f
C1585 VDD.n899 GND 0.004543f
C1586 VDD.n900 GND 0.260496f
C1587 VDD.n901 GND 0.004543f
C1588 VDD.n902 GND 0.004543f
C1589 VDD.n903 GND 0.004543f
C1590 VDD.n904 GND 0.266372f
C1591 VDD.n905 GND 0.004543f
C1592 VDD.n906 GND 0.004543f
C1593 VDD.n907 GND 0.004543f
C1594 VDD.n908 GND 0.004543f
C1595 VDD.n909 GND 0.004543f
C1596 VDD.n910 GND 0.266372f
C1597 VDD.n911 GND 0.004543f
C1598 VDD.n912 GND 0.004543f
C1599 VDD.n913 GND 0.004543f
C1600 VDD.n914 GND 0.004543f
C1601 VDD.n915 GND 0.004543f
C1602 VDD.n916 GND 0.266372f
C1603 VDD.n917 GND 0.004543f
C1604 VDD.n918 GND 0.004543f
C1605 VDD.n919 GND 0.004543f
C1606 VDD.n920 GND 0.004543f
C1607 VDD.n921 GND 0.004543f
C1608 VDD.n922 GND 0.266372f
C1609 VDD.n923 GND 0.004543f
C1610 VDD.n924 GND 0.004543f
C1611 VDD.n925 GND 0.004543f
C1612 VDD.n926 GND 0.004543f
C1613 VDD.n927 GND 0.004543f
C1614 VDD.n928 GND 0.266372f
C1615 VDD.n929 GND 0.004543f
C1616 VDD.n930 GND 0.004543f
C1617 VDD.n931 GND 0.004543f
C1618 VDD.n932 GND 0.004543f
C1619 VDD.n933 GND 0.004543f
C1620 VDD.n934 GND 0.266372f
C1621 VDD.n935 GND 0.004543f
C1622 VDD.n936 GND 0.004543f
C1623 VDD.n937 GND 0.004543f
C1624 VDD.n938 GND 0.004543f
C1625 VDD.n939 GND 0.004543f
C1626 VDD.t84 GND 0.133186f
C1627 VDD.n940 GND 0.004543f
C1628 VDD.n941 GND 0.004543f
C1629 VDD.n942 GND 0.004543f
C1630 VDD.n943 GND 0.004543f
C1631 VDD.n944 GND 0.004543f
C1632 VDD.t73 GND 0.133186f
C1633 VDD.n945 GND 0.004543f
C1634 VDD.n946 GND 0.004543f
C1635 VDD.n947 GND 0.213489f
C1636 VDD.n948 GND 0.004543f
C1637 VDD.n949 GND 0.004543f
C1638 VDD.n950 GND 0.004543f
C1639 VDD.n951 GND 0.266372f
C1640 VDD.n952 GND 0.004543f
C1641 VDD.n953 GND 0.004543f
C1642 VDD.n954 GND 0.139062f
C1643 VDD.n955 GND 0.004543f
C1644 VDD.n956 GND 0.004543f
C1645 VDD.n957 GND 0.004543f
C1646 VDD.n958 GND 0.266372f
C1647 VDD.n959 GND 0.004543f
C1648 VDD.n960 GND 0.004543f
C1649 VDD.n961 GND 0.004543f
C1650 VDD.n962 GND 0.004543f
C1651 VDD.n963 GND 0.004543f
C1652 VDD.n964 GND 0.266372f
C1653 VDD.n965 GND 0.004543f
C1654 VDD.n966 GND 0.004543f
C1655 VDD.n967 GND 0.004543f
C1656 VDD.n968 GND 0.004543f
C1657 VDD.n969 GND 0.004543f
C1658 VDD.n970 GND 0.266372f
C1659 VDD.n971 GND 0.004543f
C1660 VDD.n972 GND 0.004543f
C1661 VDD.n973 GND 0.004543f
C1662 VDD.n974 GND 0.004543f
C1663 VDD.n975 GND 0.004543f
C1664 VDD.n976 GND 0.266372f
C1665 VDD.n977 GND 0.004543f
C1666 VDD.n978 GND 0.004543f
C1667 VDD.n979 GND 0.004543f
C1668 VDD.n980 GND 0.004543f
C1669 VDD.n981 GND 0.004543f
C1670 VDD.n982 GND 0.266372f
C1671 VDD.n983 GND 0.004543f
C1672 VDD.n984 GND 0.004543f
C1673 VDD.n985 GND 0.004543f
C1674 VDD.n986 GND 0.004543f
C1675 VDD.n987 GND 0.004543f
C1676 VDD.n988 GND 0.266372f
C1677 VDD.n989 GND 0.004543f
C1678 VDD.n990 GND 0.004543f
C1679 VDD.n991 GND 0.004543f
C1680 VDD.n992 GND 0.004543f
C1681 VDD.n993 GND 0.004543f
C1682 VDD.n994 GND 0.266372f
C1683 VDD.n995 GND 0.004543f
C1684 VDD.n996 GND 0.004543f
C1685 VDD.n997 GND 0.004543f
C1686 VDD.n998 GND 0.004543f
C1687 VDD.n999 GND 0.004543f
C1688 VDD.n1000 GND 0.248744f
C1689 VDD.n1001 GND 0.004543f
C1690 VDD.n1002 GND 0.004543f
C1691 VDD.n1003 GND 0.004543f
C1692 VDD.n1004 GND 0.004543f
C1693 VDD.n1005 GND 0.004543f
C1694 VDD.n1006 GND 0.266372f
C1695 VDD.n1007 GND 0.004543f
C1696 VDD.n1008 GND 0.004543f
C1697 VDD.t83 GND 0.133186f
C1698 VDD.n1009 GND 0.004543f
C1699 VDD.n1010 GND 0.004543f
C1700 VDD.n1011 GND 0.004543f
C1701 VDD.n1012 GND 0.266372f
C1702 VDD.n1013 GND 0.004543f
C1703 VDD.n1014 GND 0.004543f
C1704 VDD.n1015 GND 0.004543f
C1705 VDD.n1016 GND 0.004543f
C1706 VDD.n1017 GND 0.004543f
C1707 VDD.n1018 GND 0.266372f
C1708 VDD.n1019 GND 0.004543f
C1709 VDD.n1020 GND 0.004543f
C1710 VDD.n1021 GND 0.004543f
C1711 VDD.n1022 GND 0.004543f
C1712 VDD.n1023 GND 0.004543f
C1713 VDD.t79 GND 0.133186f
C1714 VDD.n1024 GND 0.004543f
C1715 VDD.n1025 GND 0.004543f
C1716 VDD.n1026 GND 0.004543f
C1717 VDD.n1027 GND 0.004543f
C1718 VDD.n1028 GND 0.004543f
C1719 VDD.n1029 GND 0.266372f
C1720 VDD.n1030 GND 0.004543f
C1721 VDD.n1031 GND 0.004543f
C1722 VDD.n1032 GND 0.211531f
C1723 VDD.n1033 GND 0.004543f
C1724 VDD.n1034 GND 0.004543f
C1725 VDD.n1035 GND 0.004543f
C1726 VDD.n1036 GND 0.266372f
C1727 VDD.n1037 GND 0.004543f
C1728 VDD.n1038 GND 0.004543f
C1729 VDD.n1039 GND 0.004543f
C1730 VDD.n1040 GND 0.004543f
C1731 VDD.n1041 GND 0.004543f
C1732 VDD.n1042 GND 0.266372f
C1733 VDD.n1043 GND 0.004543f
C1734 VDD.n1044 GND 0.004543f
C1735 VDD.n1045 GND 0.004543f
C1736 VDD.n1046 GND 0.004543f
C1737 VDD.n1047 GND 0.004543f
C1738 VDD.n1048 GND 0.266372f
C1739 VDD.n1049 GND 0.004543f
C1740 VDD.n1050 GND 0.004543f
C1741 VDD.n1051 GND 0.004543f
C1742 VDD.n1052 GND 0.004543f
C1743 VDD.n1053 GND 0.004543f
C1744 VDD.n1054 GND 0.266372f
C1745 VDD.n1055 GND 0.004543f
C1746 VDD.n1056 GND 0.004543f
C1747 VDD.n1057 GND 0.004543f
C1748 VDD.n1058 GND 0.004543f
C1749 VDD.n1059 GND 0.004543f
C1750 VDD.n1060 GND 0.266372f
C1751 VDD.n1061 GND 0.004543f
C1752 VDD.n1062 GND 0.004543f
C1753 VDD.n1063 GND 0.004543f
C1754 VDD.n1064 GND 0.004543f
C1755 VDD.n1065 GND 0.004543f
C1756 VDD.n1066 GND 0.266372f
C1757 VDD.n1067 GND 0.004543f
C1758 VDD.n1068 GND 0.004543f
C1759 VDD.n1069 GND 0.004543f
C1760 VDD.n1070 GND 0.004543f
C1761 VDD.n1071 GND 0.004543f
C1762 VDD.t25 GND 0.133186f
C1763 VDD.n1072 GND 0.004543f
C1764 VDD.n1073 GND 0.004543f
C1765 VDD.n1074 GND 0.004543f
C1766 VDD.n1075 GND 0.004543f
C1767 VDD.n1076 GND 0.004543f
C1768 VDD.n1077 GND 0.176275f
C1769 VDD.n1078 GND 0.004543f
C1770 VDD.n1079 GND 0.004543f
C1771 VDD.n1080 GND 0.139062f
C1772 VDD.n1081 GND 0.004543f
C1773 VDD.n1082 GND 0.004543f
C1774 VDD.n1083 GND 0.004543f
C1775 VDD.n1084 GND 0.266372f
C1776 VDD.n1085 GND 0.004543f
C1777 VDD.n1086 GND 0.004543f
C1778 VDD.t69 GND 0.133186f
C1779 VDD.n1087 GND 0.004543f
C1780 VDD.n1088 GND 0.004543f
C1781 VDD.n1089 GND 0.004543f
C1782 VDD.n1090 GND 0.266372f
C1783 VDD.n1091 GND 0.004543f
C1784 VDD.n1092 GND 0.004543f
C1785 VDD.n1093 GND 0.004543f
C1786 VDD.n1094 GND 0.004543f
C1787 VDD.n1095 GND 0.004543f
C1788 VDD.n1096 GND 0.266372f
C1789 VDD.n1097 GND 0.004543f
C1790 VDD.n1098 GND 0.004543f
C1791 VDD.n1099 GND 0.004543f
C1792 VDD.n1100 GND 0.004543f
C1793 VDD.n1101 GND 0.004543f
C1794 VDD.n1102 GND 0.266372f
C1795 VDD.n1103 GND 0.004543f
C1796 VDD.n1104 GND 0.004543f
C1797 VDD.n1105 GND 0.004543f
C1798 VDD.n1106 GND 0.010891f
C1799 VDD.n1107 GND 0.010891f
C1800 VDD.n1108 GND 1.3632f
C1801 VDD.n1109 GND 0.010421f
C1802 VDD.n1110 GND 0.010421f
C1803 VDD.n1111 GND 0.010891f
C1804 VDD.n1112 GND 0.004543f
C1805 VDD.n1113 GND 0.004543f
C1806 VDD.n1114 GND 0.004543f
C1807 VDD.n1115 GND 0.004543f
C1808 VDD.n1116 GND 1.2391f
C1809 VDD.n1117 GND 0.004543f
C1810 VDD.n1118 GND 0.004543f
C1811 VDD.t67 GND 0.077008f
C1812 VDD.t65 GND 0.389773f
C1813 VDD.n1119 GND 0.080451f
C1814 VDD.t66 GND 0.047872f
C1815 VDD.n1120 GND 0.076995f
C1816 VDD.n1121 GND 0.004543f
C1817 VDD.n1122 GND 0.004543f
C1818 VDD.n1123 GND 0.004543f
C1819 VDD.n1124 GND 0.004543f
C1820 VDD.n1125 GND 0.004543f
C1821 VDD.n1126 GND 0.004543f
C1822 VDD.n1127 GND 0.004543f
C1823 VDD.n1128 GND 0.004543f
C1824 VDD.n1129 GND 0.004543f
C1825 VDD.n1130 GND 0.004543f
C1826 VDD.n1131 GND 0.004543f
C1827 VDD.n1132 GND 0.004543f
C1828 VDD.n1133 GND 0.004543f
C1829 VDD.n1134 GND 0.004543f
C1830 VDD.n1135 GND 0.004543f
C1831 VDD.n1136 GND 0.004543f
C1832 VDD.t27 GND 0.077008f
C1833 VDD.t24 GND 0.389773f
C1834 VDD.n1137 GND 0.080451f
C1835 VDD.t26 GND 0.047872f
C1836 VDD.n1138 GND 0.076995f
C1837 VDD.n1139 GND 0.004543f
C1838 VDD.n1140 GND 0.004543f
C1839 VDD.n1141 GND 0.004543f
C1840 VDD.n1142 GND 0.004543f
C1841 VDD.n1143 GND 0.004543f
C1842 VDD.n1144 GND 0.004543f
C1843 VDD.n1146 GND 0.004543f
C1844 VDD.n1147 GND 0.004543f
C1845 VDD.n1149 GND 0.004543f
C1846 VDD.n1150 GND 0.004543f
C1847 VDD.n1151 GND 0.004543f
C1848 VDD.n1152 GND 0.004543f
C1849 VDD.n1153 GND 0.004543f
C1850 VDD.n1155 GND 0.004543f
C1851 VDD.n1157 GND 0.004543f
C1852 VDD.n1158 GND 0.003407f
C1853 VDD.n1159 GND 0.0105f
C1854 VDD.n1160 GND 0.194761f
C1855 VDD.n1161 GND 0.002505f
C1856 VDD.n1162 GND 0.00334f
C1857 VDD.n1163 GND 0.00492f
C1858 VDD.n1164 GND 0.006681f
C1859 VDD.n1165 GND 0.006681f
C1860 VDD.n1166 GND 0.006681f
C1861 VDD.n1167 GND 0.005377f
C1862 VDD.n1168 GND 0.00334f
C1863 VDD.n1169 GND 0.006681f
C1864 VDD.n1170 GND 0.006681f
C1865 VDD.n1171 GND 0.006681f
C1866 VDD.n1172 GND 0.005377f
C1867 VDD.n1173 GND 0.00334f
C1868 VDD.n1174 GND 0.006681f
C1869 VDD.n1175 GND 0.006681f
C1870 VDD.n1176 GND 0.006681f
C1871 VDD.n1177 GND 0.005243f
C1872 VDD.n1178 GND 0.004376f
C1873 VDD.t30 GND 0.141206f
C1874 VDD.t28 GND 0.493991f
C1875 VDD.n1179 GND 0.092067f
C1876 VDD.t31 GND 0.102298f
C1877 VDD.n1180 GND 0.095951f
C1878 VDD.n1181 GND 0.006681f
C1879 VDD.n1182 GND 0.014921f
C1880 VDD.n1183 GND 0.522951f
C1881 VDD.n1190 GND 0.006681f
C1882 VDD.n1191 GND 0.00406f
C1883 VDD.t44 GND 0.141206f
C1884 VDD.t43 GND 0.493991f
C1885 VDD.n1192 GND 0.092067f
C1886 VDD.t45 GND 0.102298f
C1887 VDD.n1193 GND 0.095951f
C1888 VDD.n1194 GND 0.00334f
C1889 VDD.n1195 GND 0.005377f
C1890 VDD.n1196 GND 0.006681f
C1891 VDD.n1197 GND 0.006681f
C1892 VDD.n1198 GND 0.00334f
C1893 VDD.n1199 GND 0.005377f
C1894 VDD.n1200 GND 0.006681f
C1895 VDD.n1201 GND 0.006681f
C1896 VDD.n1202 GND 0.00334f
C1897 VDD.n1203 GND 0.006681f
C1898 VDD.n1204 GND 0.005377f
C1899 VDD.n1205 GND 0.006681f
C1900 VDD.n1206 GND 0.005377f
C1901 VDD.n1207 GND 0.006681f
C1902 VDD.n1208 GND 0.391723f
C1903 VDD.n1209 GND 0.006681f
C1904 VDD.n1210 GND 0.005377f
C1905 VDD.n1211 GND 0.004463f
C1906 VDD.n1212 GND 0.006681f
C1907 VDD.n1213 GND 0.005377f
C1908 VDD.n1214 GND 0.006681f
C1909 VDD.n1215 GND 0.264413f
C1910 VDD.n1216 GND 0.006681f
C1911 VDD.n1217 GND 0.005377f
C1912 VDD.n1218 GND 0.006681f
C1913 VDD.n1219 GND 0.005377f
C1914 VDD.n1220 GND 0.006681f
C1915 VDD.n1221 GND 0.391723f
C1916 VDD.n1222 GND 0.006681f
C1917 VDD.n1223 GND 0.005377f
C1918 VDD.n1224 GND 0.005377f
C1919 VDD.n1225 GND 0.006681f
C1920 VDD.n1226 GND 0.005377f
C1921 VDD.n1227 GND 0.006681f
C1922 VDD.n1228 GND 0.391723f
C1923 VDD.n1229 GND 0.006681f
C1924 VDD.n1230 GND 0.005377f
C1925 VDD.n1231 GND 0.006681f
C1926 VDD.n1232 GND 0.005377f
C1927 VDD.n1233 GND 0.006681f
C1928 VDD.n1234 GND 0.391723f
C1929 VDD.n1235 GND 0.006681f
C1930 VDD.n1236 GND 0.005377f
C1931 VDD.n1237 GND 0.006681f
C1932 VDD.n1238 GND 0.005377f
C1933 VDD.n1239 GND 0.006681f
C1934 VDD.n1240 GND 0.391723f
C1935 VDD.n1241 GND 0.006681f
C1936 VDD.n1242 GND 0.005377f
C1937 VDD.n1243 GND 0.006681f
C1938 VDD.n1244 GND 0.005377f
C1939 VDD.n1245 GND 0.006681f
C1940 VDD.n1246 GND 0.391723f
C1941 VDD.n1247 GND 0.006681f
C1942 VDD.n1248 GND 0.005377f
C1943 VDD.n1249 GND 0.006681f
C1944 VDD.n1250 GND 0.005377f
C1945 VDD.n1251 GND 0.006681f
C1946 VDD.n1252 GND 0.338841f
C1947 VDD.n1253 GND 0.006681f
C1948 VDD.n1254 GND 0.005377f
C1949 VDD.n1255 GND 0.006681f
C1950 VDD.n1256 GND 0.005377f
C1951 VDD.n1257 GND 0.006681f
C1952 VDD.n1258 GND 0.391723f
C1953 VDD.n1259 GND 0.006681f
C1954 VDD.n1260 GND 0.005377f
C1955 VDD.n1261 GND 0.006681f
C1956 VDD.n1262 GND 0.005377f
C1957 VDD.n1263 GND 0.006681f
C1958 VDD.n1264 GND 0.391723f
C1959 VDD.n1265 GND 0.006681f
C1960 VDD.n1266 GND 0.005377f
C1961 VDD.t10 GND 0.116461f
C1962 VDD.t6 GND 0.113326f
C1963 VDD.n1267 GND 0.538609f
C1964 VDD.t4 GND 0.116461f
C1965 VDD.t109 GND 0.113326f
C1966 VDD.n1268 GND 0.518679f
C1967 VDD.n1269 GND 0.445762f
C1968 VDD.n1270 GND 2.84627f
C1969 VDD.n1271 GND 0.40254f
C1970 VDD.n1272 GND 0.005377f
C1971 VDD.n1273 GND 0.006681f
C1972 VDD.n1274 GND 0.391723f
C1973 VDD.n1275 GND 0.006681f
C1974 VDD.n1276 GND 0.005377f
C1975 VDD.n1277 GND 0.006681f
C1976 VDD.n1278 GND 0.005377f
C1977 VDD.n1279 GND 0.006681f
C1978 VDD.n1280 GND 0.391723f
C1979 VDD.n1281 GND 0.006681f
C1980 VDD.n1282 GND 0.005377f
C1981 VDD.n1283 GND 0.006681f
C1982 VDD.n1284 GND 0.005377f
C1983 VDD.n1285 GND 0.006681f
C1984 VDD.n1286 GND 0.248744f
C1985 VDD.n1287 GND 0.006681f
C1986 VDD.n1288 GND 0.005377f
C1987 VDD.n1289 GND 0.006681f
C1988 VDD.n1290 GND 0.005377f
C1989 VDD.n1291 GND 0.006681f
C1990 VDD.n1292 GND 0.391723f
C1991 VDD.t5 GND 0.195862f
C1992 VDD.n1293 GND 0.006681f
C1993 VDD.n1294 GND 0.005377f
C1994 VDD.n1295 GND 0.006681f
C1995 VDD.n1296 GND 0.005377f
C1996 VDD.n1297 GND 0.006681f
C1997 VDD.n1298 GND 0.391723f
C1998 VDD.n1299 GND 0.006681f
C1999 VDD.n1300 GND 0.005377f
C2000 VDD.n1301 GND 0.006681f
C2001 VDD.n1302 GND 0.005377f
C2002 VDD.n1303 GND 0.006681f
C2003 VDD.n1304 GND 0.391723f
C2004 VDD.n1305 GND 0.006681f
C2005 VDD.n1306 GND 0.005377f
C2006 VDD.n1307 GND 0.006681f
C2007 VDD.n1308 GND 0.005377f
C2008 VDD.n1309 GND 0.006681f
C2009 VDD.n1310 GND 0.391723f
C2010 VDD.n1311 GND 0.006681f
C2011 VDD.n1312 GND 0.005377f
C2012 VDD.n1313 GND 0.006681f
C2013 VDD.n1314 GND 0.005377f
C2014 VDD.n1315 GND 0.006681f
C2015 VDD.n1316 GND 0.391723f
C2016 VDD.n1317 GND 0.006681f
C2017 VDD.n1318 GND 0.005377f
C2018 VDD.n1319 GND 0.006681f
C2019 VDD.n1320 GND 0.005377f
C2020 VDD.n1321 GND 0.006681f
C2021 VDD.n1322 GND 0.323172f
C2022 VDD.n1323 GND 0.006681f
C2023 VDD.n1324 GND 0.005377f
C2024 VDD.n1325 GND 0.006681f
C2025 VDD.n1326 GND 0.005377f
C2026 VDD.n1327 GND 0.006681f
C2027 VDD.n1328 GND 0.391723f
C2028 VDD.t37 GND 0.195862f
C2029 VDD.n1329 GND 0.006681f
C2030 VDD.n1330 GND 0.005377f
C2031 VDD.n1331 GND 0.006681f
C2032 VDD.n1332 GND 0.005377f
C2033 VDD.n1333 GND 0.006681f
C2034 VDD.n1334 GND 0.391723f
C2035 VDD.n1335 GND 0.006681f
C2036 VDD.n1336 GND 0.005377f
C2037 VDD.n1337 GND 0.014921f
C2038 VDD.n1338 GND 0.004463f
C2039 VDD.n1339 GND 0.014921f
C2040 VDD.n1340 GND 0.522951f
C2041 VDD.n1341 GND 0.014921f
C2042 VDD.n1342 GND 0.004463f
C2043 VDD.n1343 GND 0.006681f
C2044 VDD.n1344 GND 0.005377f
C2045 VDD.n1345 GND 0.006681f
C2046 VDD.n1358 GND 0.015143f
C2047 VDD.n1359 GND 0.006681f
C2048 VDD.n1360 GND 0.005377f
C2049 VDD.n1361 GND 0.006681f
C2050 VDD.n1362 GND 0.006681f
C2051 VDD.n1363 GND 0.006681f
C2052 VDD.n1364 GND 0.006681f
C2053 VDD.n1365 GND 0.006681f
C2054 VDD.n1366 GND 0.005377f
C2055 VDD.n1367 GND 0.006681f
C2056 VDD.n1368 GND 0.006681f
C2057 VDD.n1369 GND 0.006681f
C2058 VDD.n1370 GND 0.006681f
C2059 VDD.n1371 GND 0.006681f
C2060 VDD.n1372 GND 0.00406f
C2061 VDD.n1373 GND 0.006681f
C2062 VDD.n1374 GND 0.006681f
C2063 VDD.n1375 GND 0.006681f
C2064 VDD.n1376 GND 0.005377f
C2065 VDD.n1377 GND 0.006681f
C2066 VDD.n1378 GND 0.006681f
C2067 VDD.n1379 GND 0.006681f
C2068 VDD.n1380 GND 0.006681f
C2069 VDD.n1381 GND 0.006681f
C2070 VDD.n1382 GND 0.005377f
C2071 VDD.n1383 GND 0.006681f
C2072 VDD.n1384 GND 0.006681f
C2073 VDD.n1385 GND 0.006681f
C2074 VDD.n1386 GND 0.006681f
C2075 VDD.n1387 GND 0.006681f
C2076 VDD.n1388 GND 0.005377f
C2077 VDD.n1389 GND 0.006681f
C2078 VDD.n1390 GND 0.006681f
C2079 VDD.n1391 GND 0.006681f
C2080 VDD.n1392 GND 0.002823f
C2081 VDD.n1393 GND 0.015143f
C2082 VDD.n1394 GND 0.006681f
C2083 VDD.n1395 GND 0.006681f
C2084 VDD.t39 GND 0.141206f
C2085 VDD.t36 GND 0.493991f
C2086 VDD.n1396 GND 0.092067f
C2087 VDD.t38 GND 0.102298f
C2088 VDD.n1397 GND 0.095951f
C2089 VDD.n1398 GND 0.010082f
C2090 VDD.n1399 GND 0.005243f
C2091 VDD.n1400 GND 0.005377f
C2092 VDD.n1401 GND 0.006681f
C2093 VDD.n1402 GND 0.006681f
C2094 VDD.n1403 GND 0.006681f
C2095 VDD.n1404 GND 0.005377f
C2096 VDD.n1405 GND 0.005377f
C2097 VDD.n1406 GND 0.005377f
C2098 VDD.n1407 GND 0.006681f
C2099 VDD.n1408 GND 0.006681f
C2100 VDD.n1409 GND 0.006681f
C2101 VDD.n1410 GND 0.005377f
C2102 VDD.n1411 GND 0.005377f
C2103 VDD.n1412 GND 0.005377f
C2104 VDD.n1413 GND 0.006681f
C2105 VDD.n1414 GND 0.006681f
C2106 VDD.n1415 GND 0.006681f
C2107 VDD.n1416 GND 0.005377f
C2108 VDD.n1417 GND 0.00492f
C2109 VDD.n1418 GND 0.006681f
C2110 VDD.n1419 GND 0.006681f
C2111 VDD.t55 GND 0.141206f
C2112 VDD.t53 GND 0.493991f
C2113 VDD.n1420 GND 0.092067f
C2114 VDD.t54 GND 0.102298f
C2115 VDD.n1421 GND 0.095951f
C2116 VDD.n1422 GND 0.010082f
C2117 VDD.n1423 GND 0.006681f
C2118 VDD.n1424 GND 0.006681f
C2119 VDD.n1425 GND 0.006681f
C2120 VDD.n1426 GND 0.005377f
C2121 VDD.n1427 GND 0.005377f
C2122 VDD.n1428 GND 0.005377f
C2123 VDD.n1429 GND 0.006681f
C2124 VDD.n1430 GND 0.006681f
C2125 VDD.n1431 GND 0.006681f
C2126 VDD.n1432 GND 0.005377f
C2127 VDD.n1433 GND 0.005377f
C2128 VDD.n1434 GND 0.005377f
C2129 VDD.n1435 GND 0.006681f
C2130 VDD.n1436 GND 0.006681f
C2131 VDD.n1437 GND 0.006681f
C2132 VDD.n1438 GND 0.005377f
C2133 VDD.n1439 GND 0.006681f
C2134 VDD.n1440 GND 0.871584f
C2135 VDD.n1442 GND 0.015143f
C2136 VDD.n1443 GND 0.004463f
C2137 VDD.n1444 GND 0.015143f
C2138 VDD.n1445 GND 0.014921f
C2139 VDD.n1446 GND 0.006681f
C2140 VDD.n1447 GND 0.005377f
C2141 VDD.n1448 GND 0.006681f
C2142 VDD.n1449 GND 0.391723f
C2143 VDD.n1450 GND 0.006681f
C2144 VDD.n1451 GND 0.005377f
C2145 VDD.n1452 GND 0.006681f
C2146 VDD.n1453 GND 0.006681f
C2147 VDD.n1454 GND 0.006681f
C2148 VDD.n1455 GND 0.005377f
C2149 VDD.n1456 GND 0.006681f
C2150 VDD.n1457 GND 0.391723f
C2151 VDD.n1458 GND 0.006681f
C2152 VDD.n1459 GND 0.005377f
C2153 VDD.n1460 GND 0.006681f
C2154 VDD.n1461 GND 0.006681f
C2155 VDD.n1462 GND 0.006681f
C2156 VDD.n1463 GND 0.005377f
C2157 VDD.n1464 GND 0.006681f
C2158 VDD.n1465 GND 0.264413f
C2159 VDD.n1466 GND 0.006681f
C2160 VDD.n1467 GND 0.005377f
C2161 VDD.n1468 GND 0.006681f
C2162 VDD.n1469 GND 0.006681f
C2163 VDD.n1470 GND 0.006681f
C2164 VDD.n1471 GND 0.005377f
C2165 VDD.n1472 GND 0.006681f
C2166 VDD.n1473 GND 0.391723f
C2167 VDD.n1474 GND 0.006681f
C2168 VDD.n1475 GND 0.005377f
C2169 VDD.n1476 GND 0.006681f
C2170 VDD.n1477 GND 0.006681f
C2171 VDD.n1478 GND 0.006681f
C2172 VDD.n1479 GND 0.005377f
C2173 VDD.n1480 GND 0.006681f
C2174 VDD.n1481 GND 0.391723f
C2175 VDD.n1482 GND 0.006681f
C2176 VDD.n1483 GND 0.005377f
C2177 VDD.n1484 GND 0.006681f
C2178 VDD.n1485 GND 0.006681f
C2179 VDD.n1486 GND 0.006681f
C2180 VDD.n1487 GND 0.005377f
C2181 VDD.n1488 GND 0.006681f
C2182 VDD.n1489 GND 0.391723f
C2183 VDD.n1490 GND 0.006681f
C2184 VDD.n1491 GND 0.005377f
C2185 VDD.n1492 GND 0.006681f
C2186 VDD.n1493 GND 0.006681f
C2187 VDD.n1494 GND 0.006681f
C2188 VDD.n1495 GND 0.005377f
C2189 VDD.n1496 GND 0.006681f
C2190 VDD.n1497 GND 0.391723f
C2191 VDD.n1498 GND 0.006681f
C2192 VDD.n1499 GND 0.005377f
C2193 VDD.n1500 GND 0.006681f
C2194 VDD.n1501 GND 0.006681f
C2195 VDD.n1502 GND 0.006681f
C2196 VDD.n1503 GND 0.005377f
C2197 VDD.n1504 GND 0.006681f
C2198 VDD.n1505 GND 0.391723f
C2199 VDD.n1506 GND 0.006681f
C2200 VDD.n1507 GND 0.005377f
C2201 VDD.n1508 GND 0.006681f
C2202 VDD.n1509 GND 0.006681f
C2203 VDD.n1510 GND 0.006681f
C2204 VDD.n1511 GND 0.005377f
C2205 VDD.n1512 GND 0.006681f
C2206 VDD.n1513 GND 0.338841f
C2207 VDD.n1514 GND 0.006681f
C2208 VDD.n1515 GND 0.005377f
C2209 VDD.n1516 GND 0.006681f
C2210 VDD.n1517 GND 0.006681f
C2211 VDD.n1518 GND 0.006681f
C2212 VDD.n1519 GND 0.005377f
C2213 VDD.n1520 GND 0.006681f
C2214 VDD.n1521 GND 0.391723f
C2215 VDD.n1522 GND 0.006681f
C2216 VDD.n1523 GND 0.005377f
C2217 VDD.n1524 GND 0.006681f
C2218 VDD.n1525 GND 0.006681f
C2219 VDD.n1526 GND 0.005135f
C2220 VDD.n1527 GND 0.006681f
C2221 VDD.n1528 GND 0.005377f
C2222 VDD.n1529 GND 0.006681f
C2223 VDD.n1530 GND 0.391723f
C2224 VDD.n1531 GND 0.006681f
C2225 VDD.n1532 GND 0.005377f
C2226 VDD.n1533 GND 0.006681f
C2227 VDD.n1534 GND 0.006681f
C2228 VDD.n1535 GND 0.006681f
C2229 VDD.n1536 GND 0.005377f
C2230 VDD.n1537 GND 0.006681f
C2231 VDD.n1538 GND 0.391723f
C2232 VDD.n1539 GND 0.006681f
C2233 VDD.n1540 GND 0.005377f
C2234 VDD.n1541 GND 0.005135f
C2235 VDD.n1542 GND 0.006681f
C2236 VDD.n1543 GND 0.006681f
C2237 VDD.n1544 GND 0.005377f
C2238 VDD.n1545 GND 0.006681f
C2239 VDD.n1546 GND 0.391723f
C2240 VDD.n1547 GND 0.006681f
C2241 VDD.n1548 GND 0.005377f
C2242 VDD.n1549 GND 0.006681f
C2243 VDD.n1550 GND 0.006681f
C2244 VDD.n1551 GND 0.006681f
C2245 VDD.n1552 GND 0.005377f
C2246 VDD.n1553 GND 0.006681f
C2247 VDD.t3 GND 0.195862f
C2248 VDD.n1554 GND 0.248744f
C2249 VDD.n1555 GND 0.006681f
C2250 VDD.n1556 GND 0.005377f
C2251 VDD.n1557 GND 0.006681f
C2252 VDD.n1558 GND 0.006681f
C2253 VDD.n1559 GND 0.006681f
C2254 VDD.n1560 GND 0.005377f
C2255 VDD.n1561 GND 0.006681f
C2256 VDD.n1562 GND 0.391723f
C2257 VDD.n1563 GND 0.006681f
C2258 VDD.n1564 GND 0.005377f
C2259 VDD.n1565 GND 0.006681f
C2260 VDD.n1566 GND 0.006681f
C2261 VDD.n1567 GND 0.006681f
C2262 VDD.n1568 GND 0.005377f
C2263 VDD.n1569 GND 0.006681f
C2264 VDD.n1570 GND 0.391723f
C2265 VDD.n1571 GND 0.006681f
C2266 VDD.n1572 GND 0.005377f
C2267 VDD.n1573 GND 0.006681f
C2268 VDD.n1574 GND 0.006681f
C2269 VDD.n1575 GND 0.006681f
C2270 VDD.n1576 GND 0.005377f
C2271 VDD.n1577 GND 0.006681f
C2272 VDD.n1578 GND 0.391723f
C2273 VDD.n1579 GND 0.006681f
C2274 VDD.n1580 GND 0.005377f
C2275 VDD.n1581 GND 0.006681f
C2276 VDD.n1582 GND 0.006681f
C2277 VDD.n1583 GND 0.006681f
C2278 VDD.n1584 GND 0.005377f
C2279 VDD.n1585 GND 0.006681f
C2280 VDD.n1586 GND 0.391723f
C2281 VDD.n1587 GND 0.006681f
C2282 VDD.n1588 GND 0.005377f
C2283 VDD.n1589 GND 0.006681f
C2284 VDD.n1590 GND 0.006681f
C2285 VDD.n1591 GND 0.006681f
C2286 VDD.n1592 GND 0.005377f
C2287 VDD.n1593 GND 0.006681f
C2288 VDD.n1594 GND 0.391723f
C2289 VDD.n1595 GND 0.006681f
C2290 VDD.n1596 GND 0.005377f
C2291 VDD.n1597 GND 0.006681f
C2292 VDD.n1598 GND 0.006681f
C2293 VDD.n1599 GND 0.006681f
C2294 VDD.n1600 GND 0.006681f
C2295 VDD.n1601 GND 0.005377f
C2296 VDD.n1602 GND 0.006681f
C2297 VDD.t29 GND 0.195862f
C2298 VDD.n1603 GND 0.323172f
C2299 VDD.n1604 GND 0.006681f
C2300 VDD.n1605 GND 0.005377f
C2301 VDD.n1606 GND 0.006681f
C2302 VDD.n1607 GND 0.006681f
C2303 VDD.n1608 GND 0.006681f
C2304 VDD.n1609 GND 0.005377f
C2305 VDD.n1610 GND 0.006681f
C2306 VDD.n1611 GND 0.391723f
C2307 VDD.n1612 GND 0.006681f
C2308 VDD.n1613 GND 0.006681f
C2309 VDD.n1614 GND 0.005377f
C2310 VDD.n1615 GND 0.006681f
C2311 VDD.n1616 GND 0.006681f
C2312 VDD.n1617 GND 0.004519f
C2313 VDD.n1618 GND 0.181867f
C2314 VDD.n1619 GND 0.007549f
C2315 VDD.n1620 GND 0.006681f
C2316 VDD.n1621 GND 0.005377f
C2317 VDD.n1622 GND 0.006681f
C2318 VDD.n1623 GND 0.391723f
C2319 VDD.n1624 GND 0.391723f
C2320 VDD.n1625 GND 0.006681f
C2321 VDD.n1626 GND 0.005377f
C2322 VDD.n1627 GND 0.006681f
C2323 VDD.n1628 GND 0.006681f
C2324 VDD.n1629 GND 0.009656f
C2325 VDD.n1630 GND 0.004463f
C2326 VDD.n1631 GND 0.014921f
C2327 VDD.n1632 GND 0.015143f
C2328 VDD.n1633 GND 0.004176f
C2329 VDD.n1634 GND 0.004463f
C2330 VDD.n1635 GND 0.005377f
C2331 VDD.n1636 GND 0.006681f
C2332 VDD.n1637 GND 0.006681f
C2333 VDD.n1638 GND 0.005377f
C2334 VDD.n1639 GND 0.00334f
C2335 VDD.n1640 GND 0.00334f
C2336 VDD.n1641 GND 0.00334f
C2337 VDD.n1642 GND 0.005377f
C2338 VDD.n1643 GND 0.005377f
C2339 VDD.n1644 GND 0.006681f
C2340 VDD.n1645 GND 0.006681f
C2341 VDD.n1646 GND 0.005377f
C2342 VDD.n1647 GND 0.00334f
C2343 VDD.n1648 GND 0.00334f
C2344 VDD.n1649 GND 0.00334f
C2345 VDD.n1650 GND 0.005377f
C2346 VDD.n1651 GND 0.005377f
C2347 VDD.n1652 GND 0.006681f
C2348 VDD.n1653 GND 0.006681f
C2349 VDD.n1654 GND 0.005377f
C2350 VDD.n1655 GND 0.00334f
C2351 VDD.n1656 GND 0.00334f
C2352 VDD.n1657 GND 0.00334f
C2353 VDD.n1658 GND 0.010082f
C2354 VDD.n1659 GND 0.006681f
C2355 VDD.n1660 GND 0.006681f
C2356 VDD.n1663 GND 0.006681f
C2357 VDD.n1666 GND 0.006681f
C2358 VDD.n1669 GND 0.006681f
C2359 VDD.t76 GND 3.64107f
C2360 VDD.t98 GND 5.59381f
C2361 VDD.t68 GND 6.05017f
C2362 VDD.n1671 GND 3.30223f
C2363 VDD.n1673 GND 0.015143f
C2364 VDD.n1674 GND 0.002823f
C2365 VDD.n1675 GND 0.010082f
C2366 VDD.n1676 GND 0.00334f
C2367 VDD.n1677 GND 0.00334f
C2368 VDD.n1678 GND 0.00334f
C2369 VDD.n1679 GND 0.005377f
C2370 VDD.n1680 GND 0.005377f
C2371 VDD.n1681 GND 0.005377f
C2372 VDD.n1682 GND 0.00334f
C2373 VDD.n1683 GND 0.00334f
C2374 VDD.n1684 GND 0.00334f
C2375 VDD.n1685 GND 0.005377f
C2376 VDD.n1686 GND 0.005377f
C2377 VDD.n1687 GND 0.005377f
C2378 VDD.n1688 GND 0.00334f
C2379 VDD.n1689 GND 0.00334f
C2380 VDD.n1690 GND 0.00334f
C2381 VDD.n1691 GND 0.005377f
C2382 VDD.n1692 GND 0.005377f
C2383 VDD.n1693 GND 0.005377f
C2384 VDD.n1694 GND 0.002505f
C2385 VDD.n1695 GND 0.049304f
C2386 VDD.n1696 GND 1.5061f
C2387 VDD.n1697 GND 0.115728f
C2388 VDD.n1698 GND 0.003407f
C2389 VDD.n1699 GND 0.004543f
C2390 VDD.n1700 GND 0.004543f
C2391 VDD.n1702 GND 0.004543f
C2392 VDD.n1704 GND 0.004543f
C2393 VDD.n1705 GND 0.004042f
C2394 VDD.n1706 GND 0.005605f
C2395 VDD.n1707 GND 0.002773f
C2396 VDD.n1708 GND 0.004543f
C2397 VDD.n1709 GND 0.004543f
C2398 VDD.n1711 GND 0.004543f
C2399 VDD.n1712 GND 0.010891f
C2400 VDD.n1713 GND 0.010891f
C2401 VDD.n1714 GND 0.010421f
C2402 VDD.n1715 GND 0.004543f
C2403 VDD.n1716 GND 0.004543f
C2404 VDD.n1717 GND 0.004543f
C2405 VDD.n1718 GND 0.004543f
C2406 VDD.n1719 GND 0.004543f
C2407 VDD.n1720 GND 0.004543f
C2408 VDD.n1721 GND 0.004543f
C2409 VDD.n1722 GND 0.004543f
C2410 VDD.n1723 GND 0.004543f
C2411 VDD.n1724 GND 0.004543f
C2412 VDD.n1725 GND 0.004543f
C2413 VDD.n1726 GND 0.004543f
C2414 VDD.n1727 GND 0.004543f
C2415 VDD.n1728 GND 0.004543f
C2416 VDD.n1729 GND 0.004543f
C2417 VDD.n1730 GND 0.004543f
C2418 VDD.n1731 GND 0.004543f
C2419 VDD.n1732 GND 0.004543f
C2420 VDD.n1733 GND 0.004543f
C2421 VDD.n1734 GND 0.004543f
C2422 VDD.n1735 GND 0.004543f
C2423 VDD.n1736 GND 0.004543f
C2424 VDD.n1737 GND 0.004543f
C2425 VDD.n1738 GND 0.004543f
C2426 VDD.n1739 GND 0.004543f
C2427 VDD.n1740 GND 0.004543f
C2428 VDD.n1741 GND 0.004543f
C2429 VDD.n1742 GND 0.004543f
C2430 VDD.n1743 GND 0.004543f
C2431 VDD.n1744 GND 0.004543f
C2432 VDD.n1745 GND 0.004543f
C2433 VDD.n1746 GND 0.004543f
C2434 VDD.n1747 GND 0.004543f
C2435 VDD.n1748 GND 0.004543f
C2436 VDD.n1749 GND 0.004543f
C2437 VDD.n1750 GND 0.004543f
C2438 VDD.n1751 GND 0.004543f
C2439 VDD.n1752 GND 0.004543f
C2440 VDD.n1753 GND 0.004543f
C2441 VDD.n1754 GND 0.004543f
C2442 VDD.n1755 GND 0.004543f
C2443 VDD.n1756 GND 0.004543f
C2444 VDD.n1757 GND 0.004543f
C2445 VDD.n1758 GND 0.004543f
C2446 VDD.n1759 GND 0.004543f
C2447 VDD.n1760 GND 0.004543f
C2448 VDD.n1761 GND 0.004543f
C2449 VDD.n1762 GND 0.004543f
C2450 VDD.n1763 GND 0.004543f
C2451 VDD.n1764 GND 0.004543f
C2452 VDD.n1765 GND 0.004543f
C2453 VDD.n1766 GND 0.004543f
C2454 VDD.n1767 GND 0.004543f
C2455 VDD.n1768 GND 0.004543f
C2456 VDD.n1769 GND 0.004543f
C2457 VDD.n1770 GND 0.004543f
C2458 VDD.n1771 GND 0.004543f
C2459 VDD.n1772 GND 0.004543f
C2460 VDD.n1773 GND 0.004543f
C2461 VDD.n1774 GND 0.004543f
C2462 VDD.n1775 GND 0.004543f
C2463 VDD.n1776 GND 0.004543f
C2464 VDD.n1777 GND 0.004543f
C2465 VDD.n1778 GND 0.004543f
C2466 VDD.n1779 GND 0.004543f
C2467 VDD.n1780 GND 0.004543f
C2468 VDD.n1781 GND 0.004543f
C2469 VDD.n1782 GND 0.004543f
C2470 VDD.n1783 GND 0.004543f
C2471 VDD.n1784 GND 0.004543f
C2472 VDD.n1785 GND 0.004543f
C2473 VDD.n1786 GND 0.004543f
C2474 VDD.n1787 GND 0.004543f
C2475 VDD.n1788 GND 0.004543f
C2476 VDD.n1789 GND 0.004543f
C2477 VDD.n1790 GND 0.004543f
C2478 VDD.n1791 GND 0.004543f
C2479 VDD.n1792 GND 0.004543f
C2480 VDD.n1793 GND 0.004543f
C2481 VDD.n1794 GND 0.004543f
C2482 VDD.n1795 GND 0.004543f
C2483 VDD.n1796 GND 0.004543f
C2484 VDD.n1797 GND 0.004543f
C2485 VDD.n1798 GND 0.004543f
C2486 VDD.n1799 GND 0.004543f
C2487 VDD.n1800 GND 0.004543f
C2488 VDD.n1801 GND 0.004543f
C2489 VDD.n1802 GND 0.004543f
C2490 VDD.n1803 GND 0.004543f
C2491 VDD.n1804 GND 0.004543f
C2492 VDD.n1805 GND 0.004543f
C2493 VDD.n1806 GND 0.004543f
C2494 VDD.n1807 GND 0.004543f
C2495 VDD.n1808 GND 0.004543f
C2496 VDD.n1809 GND 0.004543f
C2497 VDD.n1810 GND 0.004543f
C2498 VDD.n1811 GND 0.004543f
C2499 VDD.n1812 GND 0.004543f
C2500 VDD.n1813 GND 0.004543f
C2501 VDD.n1814 GND 0.004543f
C2502 VDD.n1815 GND 0.004543f
C2503 VDD.n1816 GND 0.004543f
C2504 VDD.n1817 GND 0.004543f
C2505 VDD.n1818 GND 0.004543f
C2506 VDD.n1819 GND 0.004543f
C2507 VDD.n1820 GND 0.004543f
C2508 VDD.n1821 GND 0.004543f
C2509 VDD.n1822 GND 0.004543f
C2510 VDD.n1823 GND 0.004543f
C2511 VDD.n1824 GND 0.004543f
C2512 VDD.n1825 GND 0.004543f
C2513 VDD.n1826 GND 0.004543f
C2514 VDD.n1827 GND 0.004543f
C2515 VDD.n1828 GND 0.004543f
C2516 VDD.n1829 GND 0.004543f
C2517 VDD.n1830 GND 0.004543f
C2518 VDD.n1831 GND 0.004543f
C2519 VDD.n1832 GND 0.004543f
C2520 VDD.n1833 GND 0.004543f
C2521 VDD.n1834 GND 0.004543f
C2522 VDD.n1835 GND 0.004543f
C2523 VDD.n1836 GND 0.004543f
C2524 VDD.n1837 GND 0.004543f
C2525 VDD.n1838 GND 0.004543f
C2526 VDD.n1839 GND 0.004543f
C2527 VDD.n1840 GND 0.004543f
C2528 VDD.n1841 GND 0.004543f
C2529 VDD.n1842 GND 0.004543f
C2530 VDD.n1843 GND 0.004543f
C2531 VDD.n1844 GND 0.004543f
C2532 VDD.n1845 GND 0.004543f
C2533 VDD.n1846 GND 0.004543f
C2534 VDD.n1847 GND 0.004543f
C2535 VDD.n1848 GND 0.004543f
C2536 VDD.n1849 GND 0.004543f
C2537 VDD.n1850 GND 0.004543f
C2538 VDD.n1851 GND 0.004543f
C2539 VDD.n1852 GND 0.004543f
C2540 VDD.n1853 GND 0.004543f
C2541 VDD.n1854 GND 0.004543f
C2542 VDD.n1855 GND 0.004543f
C2543 VDD.n1856 GND 0.004543f
C2544 VDD.n1857 GND 0.004543f
C2545 VDD.n1858 GND 0.004543f
C2546 VDD.n1859 GND 0.004543f
C2547 VDD.n1860 GND 0.004543f
C2548 VDD.n1861 GND 0.004543f
C2549 VDD.n1862 GND 0.004543f
C2550 VDD.n1863 GND 0.004543f
C2551 VDD.n1864 GND 0.004543f
C2552 VDD.n1865 GND 0.004543f
C2553 VDD.n1866 GND 0.004543f
C2554 VDD.n1867 GND 0.004543f
C2555 VDD.n1868 GND 0.004543f
C2556 VDD.n1869 GND 0.004543f
C2557 VDD.n1870 GND 0.004543f
C2558 VDD.n1871 GND 0.004543f
C2559 VDD.n1872 GND 0.004543f
C2560 VDD.n1873 GND 0.004543f
C2561 VDD.n1874 GND 0.004543f
C2562 VDD.n1875 GND 0.004543f
C2563 VDD.n1876 GND 0.004543f
C2564 VDD.n1877 GND 0.004543f
C2565 VDD.n1878 GND 0.004543f
C2566 VDD.n1879 GND 0.004543f
C2567 VDD.n1880 GND 0.004543f
C2568 VDD.n1881 GND 0.004543f
C2569 VDD.n1882 GND 0.004543f
C2570 VDD.n1883 GND 0.004543f
C2571 VDD.n1884 GND 0.004543f
C2572 VDD.n1885 GND 0.004543f
C2573 VDD.n1886 GND 0.004543f
C2574 VDD.n1887 GND 0.004543f
C2575 VDD.n1888 GND 0.004543f
C2576 VDD.n1889 GND 0.004543f
C2577 VDD.n1890 GND 0.004543f
C2578 VDD.n1891 GND 0.004543f
C2579 VDD.n1892 GND 0.004543f
C2580 VDD.n1893 GND 0.004543f
C2581 VDD.n1894 GND 0.004543f
C2582 VDD.n1895 GND 0.004543f
C2583 VDD.n1896 GND 0.215448f
C2584 VDD.n1897 GND 0.004543f
C2585 VDD.n1898 GND 0.004543f
C2586 VDD.n1899 GND 0.004543f
C2587 VDD.n1900 GND 0.004543f
C2588 VDD.n1901 GND 0.004543f
C2589 VDD.n1902 GND 0.004543f
C2590 VDD.n1903 GND 0.004543f
C2591 VDD.n1904 GND 0.004543f
C2592 VDD.n1905 GND 0.004543f
C2593 VDD.n1906 GND 0.004543f
C2594 VDD.n1907 GND 0.004543f
C2595 VDD.n1908 GND 0.004543f
C2596 VDD.n1909 GND 0.004543f
C2597 VDD.n1910 GND 0.004543f
C2598 VDD.n1911 GND 0.004543f
C2599 VDD.n1912 GND 0.004543f
C2600 VDD.n1913 GND 0.004543f
C2601 VDD.n1914 GND 0.004543f
C2602 VDD.n1915 GND 0.004543f
C2603 VDD.n1916 GND 0.004543f
C2604 VDD.n1917 GND 0.004543f
C2605 VDD.n1918 GND 0.004543f
C2606 VDD.n1919 GND 0.004543f
C2607 VDD.n1920 GND 0.004543f
C2608 VDD.n1921 GND 0.004543f
C2609 VDD.n1922 GND 0.004543f
C2610 VDD.n1923 GND 0.004543f
C2611 VDD.n1924 GND 0.004543f
C2612 VDD.n1925 GND 0.004543f
C2613 VDD.n1926 GND 0.004543f
C2614 VDD.n1927 GND 0.004543f
C2615 VDD.n1928 GND 0.004543f
C2616 VDD.n1929 GND 0.004543f
C2617 VDD.n1930 GND 0.004543f
C2618 VDD.n1931 GND 0.004543f
C2619 VDD.n1932 GND 0.004543f
C2620 VDD.n1933 GND 0.004543f
C2621 VDD.n1934 GND 0.004543f
C2622 VDD.n1935 GND 0.004543f
C2623 VDD.n1936 GND 0.004543f
C2624 VDD.n1937 GND 0.004543f
C2625 VDD.n1938 GND 0.004543f
C2626 VDD.n1939 GND 0.004543f
C2627 VDD.n1940 GND 0.004543f
C2628 VDD.n1941 GND 0.004543f
C2629 VDD.n1942 GND 0.004543f
C2630 VDD.n1943 GND 0.004543f
C2631 VDD.n1944 GND 0.004543f
C2632 VDD.n1945 GND 0.004543f
C2633 VDD.n1946 GND 0.004543f
C2634 VDD.n1947 GND 0.004543f
C2635 VDD.n1948 GND 0.004543f
C2636 VDD.n1949 GND 0.004543f
C2637 VDD.n1950 GND 0.004543f
C2638 VDD.n1951 GND 0.004543f
C2639 VDD.n1952 GND 0.004543f
C2640 VDD.n1953 GND 0.004543f
C2641 VDD.n1954 GND 0.004543f
C2642 VDD.n1955 GND 0.004543f
C2643 VDD.n1956 GND 0.004543f
C2644 VDD.n1957 GND 0.004543f
C2645 VDD.n1958 GND 0.004543f
C2646 VDD.n1959 GND 0.004543f
C2647 VDD.n1960 GND 0.004543f
C2648 VDD.n1961 GND 0.004543f
C2649 VDD.n1962 GND 0.004543f
C2650 VDD.n1963 GND 0.004543f
C2651 VDD.n1964 GND 0.004543f
C2652 VDD.n1965 GND 0.004543f
C2653 VDD.n1966 GND 0.004543f
C2654 VDD.n1967 GND 0.004543f
C2655 VDD.n1968 GND 0.004543f
C2656 VDD.n1969 GND 0.004543f
C2657 VDD.n1970 GND 0.004543f
C2658 VDD.n1971 GND 0.004543f
C2659 VDD.n1972 GND 0.004543f
C2660 VDD.n1973 GND 0.004543f
C2661 VDD.n1974 GND 0.004543f
C2662 VDD.n1975 GND 0.004543f
C2663 VDD.n1976 GND 0.004543f
C2664 VDD.n1977 GND 0.004543f
C2665 VDD.n1978 GND 0.004543f
C2666 VDD.n1979 GND 0.004543f
C2667 VDD.n1980 GND 0.004543f
C2668 VDD.n1981 GND 0.004543f
C2669 VDD.n1982 GND 0.004543f
C2670 VDD.n1983 GND 0.004543f
C2671 VDD.n1984 GND 0.004543f
C2672 VDD.n1985 GND 0.004543f
C2673 VDD.n1986 GND 0.004543f
C2674 VDD.n1987 GND 0.004543f
C2675 VDD.n1988 GND 0.004543f
C2676 VDD.n1989 GND 0.004543f
C2677 VDD.n1990 GND 0.004543f
C2678 VDD.n1991 GND 0.004543f
C2679 VDD.n1992 GND 0.004543f
C2680 VDD.n1993 GND 0.004543f
C2681 VDD.n1994 GND 0.004543f
C2682 VDD.n1995 GND 0.004543f
C2683 VDD.n1996 GND 0.004543f
C2684 VDD.n1997 GND 0.004543f
C2685 VDD.n1998 GND 0.004543f
C2686 VDD.n1999 GND 0.004543f
C2687 VDD.n2000 GND 0.004543f
C2688 VDD.n2001 GND 0.004543f
C2689 VDD.n2002 GND 0.004543f
C2690 VDD.n2003 GND 0.004543f
C2691 VDD.n2004 GND 0.004543f
C2692 VDD.n2005 GND 0.004543f
C2693 VDD.n2006 GND 0.004543f
C2694 VDD.n2007 GND 0.004543f
C2695 VDD.n2008 GND 0.004543f
C2696 VDD.n2009 GND 0.004543f
C2697 VDD.n2010 GND 0.004543f
C2698 VDD.n2011 GND 0.004543f
C2699 VDD.n2012 GND 0.004543f
C2700 VDD.n2013 GND 0.004543f
C2701 VDD.n2014 GND 0.004543f
C2702 VDD.n2015 GND 0.004543f
C2703 VDD.n2016 GND 0.004543f
C2704 VDD.n2017 GND 0.004543f
C2705 VDD.n2018 GND 0.004543f
C2706 VDD.n2019 GND 0.004543f
C2707 VDD.n2020 GND 0.004543f
C2708 VDD.n2021 GND 0.004543f
C2709 VDD.n2022 GND 0.004543f
C2710 VDD.n2023 GND 0.004543f
C2711 VDD.n2024 GND 0.004543f
C2712 VDD.n2025 GND 0.004543f
C2713 VDD.n2026 GND 0.004543f
C2714 VDD.n2027 GND 0.004543f
C2715 VDD.n2028 GND 0.004543f
C2716 VDD.n2029 GND 0.004543f
C2717 VDD.n2030 GND 0.004543f
C2718 VDD.n2031 GND 0.004543f
C2719 VDD.n2032 GND 0.004543f
C2720 VDD.n2033 GND 0.004543f
C2721 VDD.n2034 GND 0.004543f
C2722 VDD.n2035 GND 0.004543f
C2723 VDD.n2036 GND 0.004543f
C2724 VDD.n2037 GND 0.004543f
C2725 VDD.n2038 GND 0.004543f
C2726 VDD.n2039 GND 0.004543f
C2727 VDD.n2040 GND 0.004543f
C2728 VDD.n2041 GND 0.004543f
C2729 VDD.n2042 GND 0.004543f
C2730 VDD.n2043 GND 0.004543f
C2731 VDD.n2044 GND 0.004543f
C2732 VDD.n2045 GND 0.004543f
C2733 VDD.n2046 GND 0.004543f
C2734 VDD.n2047 GND 0.004543f
C2735 VDD.n2048 GND 0.004543f
C2736 VDD.n2049 GND 0.004543f
C2737 VDD.n2050 GND 0.004543f
C2738 VDD.n2051 GND 0.004543f
C2739 VDD.n2052 GND 0.004543f
C2740 VDD.n2053 GND 0.004543f
C2741 VDD.n2054 GND 0.004543f
C2742 VDD.n2055 GND 0.004543f
C2743 VDD.n2056 GND 0.004543f
C2744 VDD.n2057 GND 0.004543f
C2745 VDD.n2058 GND 0.004543f
C2746 VDD.n2059 GND 0.004543f
C2747 VDD.n2060 GND 0.004543f
C2748 VDD.n2061 GND 0.004543f
C2749 VDD.n2062 GND 0.004543f
C2750 VDD.n2063 GND 0.004543f
C2751 VDD.n2064 GND 0.004543f
C2752 VDD.n2065 GND 0.004543f
C2753 VDD.n2066 GND 0.004543f
C2754 VDD.n2067 GND 0.010421f
C2755 VDD.n2068 GND 0.010891f
C2756 VDD.n2069 GND 0.010891f
C2757 VDD.n2071 GND 0.004543f
C2758 VDD.n2073 GND 0.004543f
C2759 VDD.n2074 GND 0.004543f
C2760 VDD.n2075 GND 0.002773f
C2761 VDD.n2076 GND 0.005605f
C2762 VDD.n2077 GND 0.004042f
C2763 VDD.n2078 GND 0.004543f
C2764 VDD.n2080 GND 0.004543f
C2765 VDD.n2082 GND 0.004543f
C2766 VDD.n2083 GND 0.004543f
C2767 VDD.n2084 GND 0.003407f
C2768 VDD.n2085 GND 0.025144f
C2769 VDD.n2086 GND 0.003407f
C2770 VDD.n2087 GND 0.004543f
C2771 VDD.n2089 GND 0.004543f
C2772 VDD.n2091 GND 0.004543f
C2773 VDD.n2092 GND 0.004543f
C2774 VDD.n2093 GND 0.004543f
C2775 VDD.n2094 GND 0.004543f
C2776 VDD.n2095 GND 0.004543f
C2777 VDD.n2097 GND 0.004543f
C2778 VDD.n2099 GND 0.004543f
C2779 VDD.n2100 GND 0.004543f
C2780 VDD.n2101 GND 0.010891f
C2781 VDD.n2102 GND 0.010421f
C2782 VDD.n2103 GND 0.010421f
C2783 VDD.n2104 GND 0.374096f
C2784 VDD.n2105 GND 0.010421f
C2785 VDD.n2106 GND 0.010421f
C2786 VDD.n2107 GND 0.004543f
C2787 VDD.n2108 GND 0.004543f
C2788 VDD.n2109 GND 0.004543f
C2789 VDD.n2110 GND 0.266372f
C2790 VDD.n2111 GND 0.004543f
C2791 VDD.n2112 GND 0.004543f
C2792 VDD.n2113 GND 0.004543f
C2793 VDD.n2114 GND 0.004543f
C2794 VDD.n2115 GND 0.004543f
C2795 VDD.n2116 GND 0.266372f
C2796 VDD.n2117 GND 0.004543f
C2797 VDD.n2118 GND 0.004543f
C2798 VDD.n2119 GND 0.004543f
C2799 VDD.n2120 GND 0.004543f
C2800 VDD.n2121 GND 0.004543f
C2801 VDD.n2122 GND 0.266372f
C2802 VDD.n2123 GND 0.004543f
C2803 VDD.n2124 GND 0.004543f
C2804 VDD.n2125 GND 0.004543f
C2805 VDD.n2126 GND 0.004543f
C2806 VDD.n2127 GND 0.004543f
C2807 VDD.n2128 GND 0.223282f
C2808 VDD.n2129 GND 0.004543f
C2809 VDD.n2130 GND 0.004543f
C2810 VDD.n2131 GND 0.004543f
C2811 VDD.n2132 GND 0.004543f
C2812 VDD.n2133 GND 0.004543f
C2813 VDD.n2134 GND 0.266372f
C2814 VDD.n2135 GND 0.004543f
C2815 VDD.n2136 GND 0.004543f
C2816 VDD.n2137 GND 0.004543f
C2817 VDD.n2138 GND 0.004543f
C2818 VDD.n2139 GND 0.004543f
C2819 VDD.n2140 GND 0.260496f
C2820 VDD.n2141 GND 0.004543f
C2821 VDD.n2142 GND 0.004543f
C2822 VDD.n2143 GND 0.004543f
C2823 VDD.n2144 GND 0.004543f
C2824 VDD.n2145 GND 0.004543f
C2825 VDD.n2146 GND 0.266372f
C2826 VDD.n2147 GND 0.004543f
C2827 VDD.n2148 GND 0.004543f
C2828 VDD.n2149 GND 0.004543f
C2829 VDD.n2150 GND 0.004543f
C2830 VDD.n2151 GND 0.004543f
C2831 VDD.n2152 GND 0.266372f
C2832 VDD.n2153 GND 0.004543f
C2833 VDD.n2154 GND 0.004543f
C2834 VDD.n2155 GND 0.004543f
C2835 VDD.n2156 GND 0.004543f
C2836 VDD.n2157 GND 0.004543f
C2837 VDD.n2158 GND 0.266372f
C2838 VDD.n2159 GND 0.004543f
C2839 VDD.n2160 GND 0.004543f
C2840 VDD.n2161 GND 0.004543f
C2841 VDD.n2162 GND 0.004543f
C2842 VDD.n2163 GND 0.004543f
C2843 VDD.n2164 GND 0.266372f
C2844 VDD.n2165 GND 0.004543f
C2845 VDD.n2166 GND 0.004543f
C2846 VDD.n2167 GND 0.004543f
C2847 VDD.n2168 GND 0.004543f
C2848 VDD.n2169 GND 0.004543f
C2849 VDD.n2170 GND 0.266372f
C2850 VDD.n2171 GND 0.004543f
C2851 VDD.n2172 GND 0.004543f
C2852 VDD.n2173 GND 0.004543f
C2853 VDD.n2174 GND 0.004543f
C2854 VDD.n2175 GND 0.004543f
C2855 VDD.n2176 GND 0.266372f
C2856 VDD.n2177 GND 0.004543f
C2857 VDD.n2178 GND 0.004543f
C2858 VDD.n2179 GND 0.004543f
C2859 VDD.n2180 GND 0.004543f
C2860 VDD.n2181 GND 0.004543f
C2861 VDD.n2182 GND 0.266372f
C2862 VDD.n2183 GND 0.004543f
C2863 VDD.n2184 GND 0.004543f
C2864 VDD.n2185 GND 0.004543f
C2865 VDD.n2186 GND 0.004543f
C2866 VDD.n2187 GND 0.004543f
C2867 VDD.n2188 GND 0.188027f
C2868 VDD.n2189 GND 0.004543f
C2869 VDD.n2190 GND 0.004543f
C2870 VDD.n2191 GND 0.004543f
C2871 VDD.n2192 GND 0.004543f
C2872 VDD.n2193 GND 0.004543f
C2873 VDD.n2194 GND 0.266372f
C2874 VDD.n2195 GND 0.004543f
C2875 VDD.n2196 GND 0.004543f
C2876 VDD.n2197 GND 0.004543f
C2877 VDD.n2198 GND 0.004543f
C2878 VDD.n2199 GND 0.004543f
C2879 VDD.n2200 GND 0.266372f
C2880 VDD.n2201 GND 0.004543f
C2881 VDD.n2202 GND 0.004543f
C2882 VDD.n2203 GND 0.004543f
C2883 VDD.n2204 GND 0.004543f
C2884 VDD.n2205 GND 0.004543f
C2885 VDD.n2206 GND 0.150813f
C2886 VDD.n2207 GND 0.004543f
C2887 VDD.n2208 GND 0.004543f
C2888 VDD.n2209 GND 0.004543f
C2889 VDD.n2210 GND 0.004543f
C2890 VDD.n2211 GND 0.004543f
C2891 VDD.n2212 GND 0.266372f
C2892 VDD.n2213 GND 0.004543f
C2893 VDD.n2214 GND 0.004543f
C2894 VDD.n2215 GND 0.004543f
C2895 VDD.n2216 GND 0.004543f
C2896 VDD.n2217 GND 0.004543f
C2897 VDD.n2218 GND 0.266372f
C2898 VDD.n2219 GND 0.004543f
C2899 VDD.n2220 GND 0.004543f
C2900 VDD.n2221 GND 0.004543f
C2901 VDD.n2222 GND 0.004543f
C2902 VDD.n2223 GND 0.004543f
C2903 VDD.n2224 GND 0.266372f
C2904 VDD.n2225 GND 0.004543f
C2905 VDD.n2226 GND 0.004543f
C2906 VDD.n2227 GND 0.004543f
C2907 VDD.n2228 GND 0.004543f
C2908 VDD.n2229 GND 0.004543f
C2909 VDD.n2230 GND 0.266372f
C2910 VDD.n2231 GND 0.004543f
C2911 VDD.n2232 GND 0.004543f
C2912 VDD.n2233 GND 0.004543f
C2913 VDD.n2234 GND 0.004543f
C2914 VDD.n2235 GND 0.004543f
C2915 VDD.n2236 GND 0.266372f
C2916 VDD.n2237 GND 0.004543f
C2917 VDD.n2238 GND 0.004543f
C2918 VDD.n2239 GND 0.004543f
C2919 VDD.n2240 GND 0.004543f
C2920 VDD.n2241 GND 0.004543f
C2921 VDD.n2242 GND 0.266372f
C2922 VDD.n2243 GND 0.004543f
C2923 VDD.n2244 GND 0.004543f
C2924 VDD.n2245 GND 0.004543f
C2925 VDD.n2246 GND 0.004543f
C2926 VDD.n2247 GND 0.004543f
C2927 VDD.n2248 GND 0.266372f
C2928 VDD.n2249 GND 0.004543f
C2929 VDD.n2250 GND 0.004543f
C2930 VDD.n2251 GND 0.004543f
C2931 VDD.n2252 GND 0.004543f
C2932 VDD.n2253 GND 0.004543f
C2933 VDD.n2254 GND 0.266372f
C2934 VDD.n2255 GND 0.004543f
C2935 VDD.n2256 GND 0.004543f
C2936 VDD.n2257 GND 0.004543f
C2937 VDD.n2258 GND 0.004543f
C2938 VDD.n2259 GND 0.004543f
C2939 VDD.n2260 GND 0.266372f
C2940 VDD.n2261 GND 0.004543f
C2941 VDD.n2262 GND 0.004543f
C2942 VDD.n2263 GND 0.004543f
C2943 VDD.n2264 GND 0.004543f
C2944 VDD.n2265 GND 0.004543f
C2945 VDD.n2266 GND 0.260496f
C2946 VDD.n2267 GND 0.004543f
C2947 VDD.n2268 GND 0.004543f
C2948 VDD.n2269 GND 0.004543f
C2949 VDD.n2270 GND 0.004543f
C2950 VDD.n2271 GND 0.004543f
C2951 VDD.n2272 GND 0.186069f
C2952 VDD.n2273 GND 0.004543f
C2953 VDD.n2274 GND 0.004543f
C2954 VDD.n2275 GND 0.004543f
C2955 VDD.n2276 GND 0.004543f
C2956 VDD.n2277 GND 0.004543f
C2957 VDD.n2278 GND 0.266372f
C2958 VDD.n2279 GND 0.004543f
C2959 VDD.n2280 GND 0.004543f
C2960 VDD.n2281 GND 0.004543f
C2961 VDD.n2282 GND 0.004543f
C2962 VDD.n2283 GND 0.004543f
C2963 VDD.n2284 GND 0.266372f
C2964 VDD.n2285 GND 0.004543f
C2965 VDD.n2286 GND 0.004543f
C2966 VDD.n2287 GND 0.004543f
C2967 VDD.n2288 GND 0.004543f
C2968 VDD.n2289 GND 0.004543f
C2969 VDD.n2290 GND 0.266372f
C2970 VDD.n2291 GND 0.004543f
C2971 VDD.n2292 GND 0.004543f
C2972 VDD.n2293 GND 0.004543f
C2973 VDD.n2294 GND 0.004543f
C2974 VDD.n2295 GND 0.004543f
C2975 VDD.n2296 GND 0.266372f
C2976 VDD.n2297 GND 0.004543f
C2977 VDD.n2298 GND 0.004543f
C2978 VDD.n2299 GND 0.004543f
C2979 VDD.n2300 GND 0.004543f
C2980 VDD.n2301 GND 0.004543f
C2981 VDD.n2302 GND 0.266372f
C2982 VDD.n2303 GND 0.004543f
C2983 VDD.n2304 GND 0.004543f
C2984 VDD.n2305 GND 0.004543f
C2985 VDD.n2306 GND 0.004543f
C2986 VDD.n2307 GND 0.004543f
C2987 VDD.n2308 GND 0.266372f
C2988 VDD.n2309 GND 0.004543f
C2989 VDD.n2310 GND 0.004543f
C2990 VDD.n2311 GND 0.004543f
C2991 VDD.n2312 GND 0.004543f
C2992 VDD.n2313 GND 0.004543f
C2993 VDD.n2314 GND 0.266372f
C2994 VDD.n2315 GND 0.004543f
C2995 VDD.n2316 GND 0.004543f
C2996 VDD.n2317 GND 0.004543f
C2997 VDD.n2318 GND 0.004543f
C2998 VDD.n2319 GND 0.004543f
C2999 VDD.n2320 GND 0.139062f
C3000 VDD.n2321 GND 0.004543f
C3001 VDD.n2322 GND 0.004543f
C3002 VDD.n2323 GND 0.004543f
C3003 VDD.n2324 GND 0.004543f
C3004 VDD.n2325 GND 0.004543f
C3005 VDD.n2326 GND 0.201738f
C3006 VDD.n2327 GND 0.004543f
C3007 VDD.n2328 GND 0.004543f
C3008 VDD.n2329 GND 0.004543f
C3009 VDD.n2330 GND 0.004543f
C3010 VDD.n2331 GND 0.004543f
C3011 VDD.n2332 GND 0.266372f
C3012 VDD.n2333 GND 0.004543f
C3013 VDD.n2334 GND 0.004543f
C3014 VDD.n2335 GND 0.004543f
C3015 VDD.n2336 GND 0.004543f
C3016 VDD.n2337 GND 0.004543f
C3017 VDD.n2338 GND 0.266372f
C3018 VDD.n2339 GND 0.004543f
C3019 VDD.n2340 GND 0.004543f
C3020 VDD.n2341 GND 0.004543f
C3021 VDD.n2342 GND 0.004543f
C3022 VDD.n2343 GND 0.004543f
C3023 VDD.n2344 GND 0.266372f
C3024 VDD.n2345 GND 0.004543f
C3025 VDD.n2346 GND 0.004543f
C3026 VDD.n2347 GND 0.004543f
C3027 VDD.n2348 GND 0.004543f
C3028 VDD.n2349 GND 0.004543f
C3029 VDD.n2350 GND 0.266372f
C3030 VDD.n2351 GND 0.004543f
C3031 VDD.n2352 GND 0.004543f
C3032 VDD.n2353 GND 0.004543f
C3033 VDD.n2354 GND 0.004543f
C3034 VDD.n2355 GND 0.004543f
C3035 VDD.n2356 GND 0.266372f
C3036 VDD.n2357 GND 0.004543f
C3037 VDD.n2358 GND 0.004543f
C3038 VDD.n2359 GND 0.004543f
C3039 VDD.n2360 GND 0.004543f
C3040 VDD.n2361 GND 0.004543f
C3041 VDD.n2362 GND 0.266372f
C3042 VDD.n2363 GND 0.004543f
C3043 VDD.n2364 GND 0.004543f
C3044 VDD.n2365 GND 0.004543f
C3045 VDD.n2366 GND 0.004543f
C3046 VDD.n2367 GND 0.004543f
C3047 VDD.n2368 GND 0.266372f
C3048 VDD.n2369 GND 0.004543f
C3049 VDD.n2370 GND 0.004543f
C3050 VDD.n2371 GND 0.004543f
C3051 VDD.n2372 GND 0.004543f
C3052 VDD.n2373 GND 0.004543f
C3053 VDD.n2374 GND 0.248744f
C3054 VDD.n2375 GND 0.004543f
C3055 VDD.n2376 GND 0.004543f
C3056 VDD.n2377 GND 0.004543f
C3057 VDD.n2378 GND 0.004543f
C3058 VDD.n2379 GND 0.004543f
C3059 VDD.n2380 GND 0.266372f
C3060 VDD.n2381 GND 0.004543f
C3061 VDD.n2382 GND 0.004543f
C3062 VDD.n2383 GND 0.004543f
C3063 VDD.n2384 GND 0.004543f
C3064 VDD.n2385 GND 0.004543f
C3065 VDD.n2386 GND 0.209572f
C3066 VDD.n2387 GND 0.004543f
C3067 VDD.n2388 GND 0.004543f
C3068 VDD.n2389 GND 0.004543f
C3069 VDD.n2390 GND 0.004543f
C3070 VDD.n2391 GND 0.004543f
C3071 VDD.n2392 GND 0.266372f
C3072 VDD.n2393 GND 0.004543f
C3073 VDD.n2394 GND 0.004543f
C3074 VDD.n2395 GND 0.004543f
C3075 VDD.n2396 GND 0.004543f
C3076 VDD.n2397 GND 0.004543f
C3077 VDD.n2398 GND 0.266372f
C3078 VDD.n2399 GND 0.004543f
C3079 VDD.n2400 GND 0.004543f
C3080 VDD.n2401 GND 0.004543f
C3081 VDD.n2402 GND 0.004543f
C3082 VDD.n2403 GND 0.004543f
C3083 VDD.n2404 GND 0.266372f
C3084 VDD.n2405 GND 0.004543f
C3085 VDD.n2406 GND 0.004543f
C3086 VDD.n2407 GND 0.004543f
C3087 VDD.n2408 GND 0.004543f
C3088 VDD.n2409 GND 0.004543f
C3089 VDD.n2410 GND 0.266372f
C3090 VDD.n2411 GND 0.004543f
C3091 VDD.n2412 GND 0.004543f
C3092 VDD.n2413 GND 0.004543f
C3093 VDD.n2414 GND 0.004543f
C3094 VDD.n2415 GND 0.004543f
C3095 VDD.n2416 GND 0.266372f
C3096 VDD.n2417 GND 0.004543f
C3097 VDD.n2418 GND 0.004543f
C3098 VDD.n2419 GND 0.004543f
C3099 VDD.n2420 GND 0.004543f
C3100 VDD.n2421 GND 0.004543f
C3101 VDD.n2422 GND 0.266372f
C3102 VDD.n2423 GND 0.004543f
C3103 VDD.n2424 GND 0.004543f
C3104 VDD.n2425 GND 0.004543f
C3105 VDD.n2426 GND 0.004543f
C3106 VDD.n2427 GND 0.004543f
C3107 VDD.n2428 GND 0.266372f
C3108 VDD.n2429 GND 0.004543f
C3109 VDD.n2430 GND 0.004543f
C3110 VDD.n2431 GND 0.004543f
C3111 VDD.n2432 GND 0.004543f
C3112 VDD.n2433 GND 0.004543f
C3113 VDD.n2434 GND 0.266372f
C3114 VDD.n2435 GND 0.004543f
C3115 VDD.n2436 GND 0.004543f
C3116 VDD.n2437 GND 0.004543f
C3117 VDD.n2438 GND 0.004543f
C3118 VDD.n2439 GND 0.004543f
C3119 VDD.n2440 GND 0.178234f
C3120 VDD.n2441 GND 0.004543f
C3121 VDD.n2442 GND 0.004543f
C3122 VDD.n2443 GND 0.004543f
C3123 VDD.n2444 GND 0.004543f
C3124 VDD.n2445 GND 0.004543f
C3125 VDD.n2446 GND 0.139062f
C3126 VDD.n2447 GND 0.004543f
C3127 VDD.n2448 GND 0.004543f
C3128 VDD.n2449 GND 0.004543f
C3129 VDD.n2450 GND 0.004543f
C3130 VDD.n2451 GND 0.004543f
C3131 VDD.n2452 GND 0.266372f
C3132 VDD.n2453 GND 0.004543f
C3133 VDD.n2454 GND 0.004543f
C3134 VDD.n2455 GND 0.004543f
C3135 VDD.n2456 GND 0.004543f
C3136 VDD.n2457 GND 0.004543f
C3137 VDD.n2458 GND 0.266372f
C3138 VDD.n2459 GND 0.004543f
C3139 VDD.n2460 GND 0.004543f
C3140 VDD.n2461 GND 0.004543f
C3141 VDD.t18 GND 0.077008f
C3142 VDD.t16 GND 0.389773f
C3143 VDD.n2462 GND 0.080451f
C3144 VDD.t19 GND 0.047872f
C3145 VDD.n2463 GND 0.076995f
C3146 VDD.n2464 GND 0.005605f
C3147 VDD.n2465 GND 0.004543f
C3148 VDD.n2466 GND 0.004543f
C3149 VDD.n2467 GND 0.002773f
C3150 VDD.n2468 GND 0.004543f
C3151 VDD.n2469 GND 0.004543f
C3152 VDD.n2470 GND 0.004042f
C3153 VDD.n2471 GND 0.004543f
C3154 VDD.n2472 GND 0.004543f
C3155 VDD.n2473 GND 0.004543f
C3156 VDD.n2474 GND 0.004543f
C3157 VDD.n2475 GND 0.004543f
C3158 VDD.n2476 GND 0.004543f
C3159 VDD.n2477 GND 0.004543f
C3160 VDD.n2478 GND 0.004543f
C3161 VDD.n2479 GND 0.004543f
C3162 VDD.n2480 GND 0.004543f
C3163 VDD.n2481 GND 0.004543f
C3164 VDD.n2482 GND 0.004543f
C3165 VDD.n2483 GND 0.004543f
C3166 VDD.n2484 GND 0.004543f
C3167 VDD.n2485 GND 0.004543f
C3168 VDD.n2486 GND 0.004543f
C3169 VDD.n2487 GND 0.004543f
C3170 VDD.n2488 GND 0.004543f
C3171 VDD.n2489 GND 0.004543f
C3172 VDD.n2490 GND 0.004543f
C3173 VDD.n2491 GND 0.010891f
C3174 VDD.n2492 GND 0.010891f
C3175 VDD.n2493 GND 0.010421f
C3176 VDD.n2494 GND 0.010421f
C3177 VDD.n2495 GND 0.004543f
C3178 VDD.n2496 GND 0.004543f
C3179 VDD.n2497 GND 0.004543f
C3180 VDD.n2498 GND 0.004543f
C3181 VDD.n2499 GND 0.004543f
C3182 VDD.n2500 GND 0.004543f
C3183 VDD.n2501 GND 0.004543f
C3184 VDD.n2502 GND 0.266372f
C3185 VDD.n2503 GND 0.004543f
C3186 VDD.n2504 GND 0.004543f
C3187 VDD.n2505 GND 0.004543f
C3188 VDD.n2506 GND 0.004543f
C3189 VDD.n2507 GND 0.004543f
C3190 VDD.n2508 GND 0.266372f
C3191 VDD.n2509 GND 0.004543f
C3192 VDD.n2510 GND 0.004543f
C3193 VDD.n2511 GND 0.004543f
C3194 VDD.n2512 GND 0.004543f
C3195 VDD.n2513 GND 0.010956f
C3196 VDD.n2514 GND 0.010421f
C3197 VDD.n2515 GND 0.010891f
C3198 VDD.n2516 GND 0.010356f
C3199 VDD.n2517 GND 0.004543f
C3200 VDD.n2518 GND 0.004543f
C3201 VDD.n2519 GND 0.004543f
C3202 VDD.n2520 GND 0.004543f
C3203 VDD.n2521 GND 0.002773f
C3204 VDD.n2522 GND 0.004543f
C3205 VDD.n2523 GND 0.004543f
C3206 VDD.n2524 GND 0.004042f
C3207 VDD.n2525 GND 0.004543f
C3208 VDD.n2526 GND 0.004543f
C3209 VDD.n2527 GND 0.004543f
C3210 VDD.n2528 GND 0.004543f
C3211 VDD.n2529 GND 0.004543f
C3212 VDD.n2530 GND 0.004543f
C3213 VDD.n2531 GND 0.004543f
C3214 VDD.n2532 GND 0.004543f
C3215 VDD.n2533 GND 0.004543f
C3216 VDD.n2534 GND 0.004543f
C3217 VDD.n2535 GND 0.004543f
C3218 VDD.n2536 GND 0.004543f
C3219 VDD.n2537 GND 0.004543f
C3220 VDD.n2538 GND 0.004543f
C3221 VDD.n2539 GND 0.004543f
C3222 VDD.n2540 GND 0.004543f
C3223 VDD.n2541 GND 0.004543f
C3224 VDD.n2542 GND 0.004543f
C3225 VDD.n2543 GND 0.004543f
C3226 VDD.n2544 GND 0.004543f
C3227 VDD.n2545 GND 0.010891f
C3228 VDD.n2546 GND 0.010891f
C3229 VDD.n2547 GND 0.010421f
C3230 VDD.n2548 GND 0.004543f
C3231 VDD.n2549 GND 0.004543f
C3232 VDD.n2550 GND 0.266372f
C3233 VDD.n2551 GND 0.004543f
C3234 VDD.n2552 GND 0.004543f
C3235 VDD.n2553 GND 0.010956f
C3236 VDD.n2554 GND 0.010356f
C3237 VDD.n2555 GND 0.010891f
C3238 VDD.n2557 GND 1.66287f
C3239 VDD.n2558 GND 1.66287f
C3240 VDD.n2559 GND 0.010891f
C3241 VDD.n2560 GND 0.004543f
C3242 VDD.n2561 GND 0.004543f
C3243 VDD.n2562 GND 0.002773f
C3244 VDD.n2563 GND 0.004543f
C3245 VDD.n2564 GND 0.004543f
C3246 VDD.n2565 GND 0.004543f
C3247 VDD.n2566 GND 0.004543f
C3248 VDD.n2567 GND 0.004543f
C3249 VDD.n2569 GND 0.004543f
C3250 VDD.n2570 GND 0.004543f
C3251 VDD.n2571 GND 0.004543f
C3252 VDD.n2572 GND 0.004543f
C3253 VDD.n2573 GND 0.004543f
C3254 VDD.n2575 GND 0.004543f
C3255 VDD.n2577 GND 0.004543f
C3256 VDD.n2578 GND 0.004543f
C3257 VDD.n2579 GND 0.004543f
C3258 VDD.n2580 GND 0.004543f
C3259 VDD.n2581 GND 0.004543f
C3260 VDD.n2583 GND 0.004543f
C3261 VDD.n2585 GND 0.004543f
C3262 VDD.n2586 GND 0.004543f
C3263 VDD.n2587 GND 0.004543f
C3264 VDD.t48 GND 0.077008f
C3265 VDD.t46 GND 0.389773f
C3266 VDD.n2588 GND 0.080451f
C3267 VDD.t47 GND 0.047872f
C3268 VDD.n2589 GND 0.076995f
C3269 VDD.n2590 GND 0.005605f
C3270 VDD.n2591 GND 0.004042f
C3271 VDD.n2592 GND 0.004543f
C3272 VDD.n2594 GND 0.004543f
C3273 VDD.n2595 GND 0.004543f
C3274 VDD.n2597 GND 0.004543f
C3275 VDD.n2598 GND 0.004543f
C3276 VDD.n2599 GND 0.010891f
C3277 VDD.n2600 GND 0.004543f
C3278 VDD.n2601 GND 0.004543f
C3279 VDD.n2602 GND 0.004543f
C3280 VDD.n2603 GND 0.004543f
C3281 VDD.n2604 GND 0.004543f
C3282 VDD.n2605 GND 0.004543f
C3283 VDD.n2606 GND 0.004543f
C3284 VDD.n2607 GND 0.004543f
C3285 VDD.n2608 GND 0.004543f
C3286 VDD.n2609 GND 0.004543f
C3287 VDD.n2610 GND 0.004543f
C3288 VDD.n2611 GND 0.004543f
C3289 VDD.n2612 GND 0.004543f
C3290 VDD.n2613 GND 0.004543f
C3291 VDD.n2614 GND 0.004543f
C3292 VDD.n2615 GND 0.004543f
C3293 VDD.n2616 GND 0.004543f
C3294 VDD.n2617 GND 0.004543f
C3295 VDD.n2618 GND 0.004543f
C3296 VDD.n2619 GND 0.004543f
C3297 VDD.n2620 GND 0.004543f
C3298 VDD.n2621 GND 0.004543f
C3299 VDD.n2622 GND 0.004543f
C3300 VDD.n2623 GND 0.004543f
C3301 VDD.n2624 GND 0.004543f
C3302 VDD.n2625 GND 0.004543f
C3303 VDD.n2626 GND 0.004543f
C3304 VDD.n2627 GND 0.004543f
C3305 VDD.n2628 GND 0.004543f
C3306 VDD.n2629 GND 0.004543f
C3307 VDD.n2630 GND 0.004543f
C3308 VDD.n2631 GND 0.004543f
C3309 VDD.n2632 GND 0.004543f
C3310 VDD.n2633 GND 0.004543f
C3311 VDD.n2634 GND 0.004543f
C3312 VDD.n2635 GND 0.004543f
C3313 VDD.n2636 GND 0.004543f
C3314 VDD.n2637 GND 0.004543f
C3315 VDD.n2638 GND 0.004543f
C3316 VDD.n2639 GND 0.004543f
C3317 VDD.n2640 GND 0.004543f
C3318 VDD.n2641 GND 0.004543f
C3319 VDD.n2642 GND 0.004543f
C3320 VDD.n2643 GND 0.004543f
C3321 VDD.n2644 GND 0.004543f
C3322 VDD.n2645 GND 0.004543f
C3323 VDD.n2646 GND 0.004543f
C3324 VDD.n2647 GND 0.004543f
C3325 VDD.n2648 GND 0.004543f
C3326 VDD.n2649 GND 0.004543f
C3327 VDD.n2650 GND 0.004543f
C3328 VDD.n2651 GND 0.004543f
C3329 VDD.n2652 GND 0.004543f
C3330 VDD.n2653 GND 0.004543f
C3331 VDD.n2654 GND 0.004543f
C3332 VDD.n2655 GND 0.004543f
C3333 VDD.n2656 GND 0.004543f
C3334 VDD.n2657 GND 0.004543f
C3335 VDD.n2658 GND 0.004543f
C3336 VDD.n2659 GND 0.004543f
C3337 VDD.n2660 GND 0.004543f
C3338 VDD.n2661 GND 0.004543f
C3339 VDD.n2662 GND 0.004543f
C3340 VDD.n2663 GND 0.004543f
C3341 VDD.n2664 GND 0.004543f
C3342 VDD.n2665 GND 0.004543f
C3343 VDD.n2666 GND 0.004543f
C3344 VDD.n2667 GND 0.004543f
C3345 VDD.n2668 GND 0.004543f
C3346 VDD.n2669 GND 0.004543f
C3347 VDD.n2670 GND 0.004543f
C3348 VDD.n2671 GND 0.004543f
C3349 VDD.n2672 GND 0.004543f
C3350 VDD.n2673 GND 0.004543f
C3351 VDD.n2674 GND 0.004543f
C3352 VDD.n2675 GND 0.004543f
C3353 VDD.n2676 GND 0.004543f
C3354 VDD.n2677 GND 0.004543f
C3355 VDD.n2678 GND 0.004543f
C3356 VDD.n2679 GND 0.004543f
C3357 VDD.n2680 GND 0.004543f
C3358 VDD.n2681 GND 0.004543f
C3359 VDD.n2682 GND 0.004543f
C3360 VDD.n2683 GND 0.004543f
C3361 VDD.n2684 GND 0.004543f
C3362 VDD.n2685 GND 0.004543f
C3363 VDD.n2686 GND 0.004543f
C3364 VDD.n2687 GND 0.004543f
C3365 VDD.n2688 GND 0.004543f
C3366 VDD.n2689 GND 0.004543f
C3367 VDD.n2690 GND 0.004543f
C3368 VDD.n2691 GND 0.004543f
C3369 VDD.n2692 GND 0.004543f
C3370 VDD.n2693 GND 0.004543f
C3371 VDD.n2694 GND 0.004543f
C3372 VDD.n2695 GND 0.004543f
C3373 VDD.n2696 GND 0.004543f
C3374 VDD.n2697 GND 0.004543f
C3375 VDD.n2698 GND 0.004543f
C3376 VDD.n2699 GND 0.004543f
C3377 VDD.n2700 GND 0.004543f
C3378 VDD.n2701 GND 0.004543f
C3379 VDD.n2702 GND 0.004543f
C3380 VDD.n2703 GND 0.004543f
C3381 VDD.n2704 GND 0.004543f
C3382 VDD.n2705 GND 0.004543f
C3383 VDD.n2706 GND 0.004543f
C3384 VDD.n2707 GND 0.004543f
C3385 VDD.n2708 GND 0.004543f
C3386 VDD.n2709 GND 0.004543f
C3387 VDD.n2710 GND 0.004543f
C3388 VDD.n2711 GND 0.004543f
C3389 VDD.n2712 GND 0.004543f
C3390 VDD.n2713 GND 0.004543f
C3391 VDD.n2714 GND 0.004543f
C3392 VDD.n2715 GND 0.004543f
C3393 VDD.n2716 GND 0.004543f
C3394 VDD.n2717 GND 0.004543f
C3395 VDD.n2718 GND 0.004543f
C3396 VDD.n2719 GND 0.004543f
C3397 VDD.n2720 GND 0.004543f
C3398 VDD.n2721 GND 0.004543f
C3399 VDD.n2722 GND 0.004543f
C3400 VDD.n2723 GND 0.004543f
C3401 VDD.n2724 GND 0.004543f
C3402 VDD.n2725 GND 0.004543f
C3403 VDD.n2726 GND 0.004543f
C3404 VDD.n2727 GND 0.004543f
C3405 VDD.n2728 GND 0.004543f
C3406 VDD.n2729 GND 0.004543f
C3407 VDD.n2730 GND 0.004543f
C3408 VDD.n2731 GND 0.004543f
C3409 VDD.n2732 GND 0.004543f
C3410 VDD.n2733 GND 0.004543f
C3411 VDD.n2734 GND 0.004543f
C3412 VDD.n2735 GND 0.004543f
C3413 VDD.n2736 GND 0.004543f
C3414 VDD.n2737 GND 0.004543f
C3415 VDD.n2738 GND 0.004543f
C3416 VDD.n2739 GND 0.004543f
C3417 VDD.n2740 GND 0.004543f
C3418 VDD.n2741 GND 0.004543f
C3419 VDD.n2742 GND 0.004543f
C3420 VDD.n2743 GND 0.004543f
C3421 VDD.n2744 GND 0.004543f
C3422 VDD.n2745 GND 0.004543f
C3423 VDD.n2746 GND 0.004543f
C3424 VDD.n2747 GND 0.004543f
C3425 VDD.n2748 GND 0.004543f
C3426 VDD.n2749 GND 0.004543f
C3427 VDD.n2750 GND 0.004543f
C3428 VDD.n2751 GND 0.004543f
C3429 VDD.n2752 GND 0.004543f
C3430 VDD.n2753 GND 0.004543f
C3431 VDD.n2754 GND 0.004543f
C3432 VDD.n2755 GND 0.004543f
C3433 VDD.n2756 GND 0.004543f
C3434 VDD.n2757 GND 0.004543f
C3435 VDD.n2758 GND 0.004543f
C3436 VDD.n2759 GND 0.004543f
C3437 VDD.n2760 GND 0.004543f
C3438 VDD.n2761 GND 0.004543f
C3439 VDD.n2762 GND 0.004543f
C3440 VDD.n2763 GND 0.004543f
C3441 VDD.n2764 GND 0.004543f
C3442 VDD.n2765 GND 0.004543f
C3443 VDD.n2766 GND 0.004543f
C3444 VDD.n2767 GND 0.004543f
C3445 VDD.n2768 GND 0.004543f
C3446 VDD.n2769 GND 0.004543f
C3447 VDD.n2770 GND 0.004543f
C3448 VDD.n2771 GND 0.004543f
C3449 VDD.n2772 GND 0.004543f
C3450 VDD.n2773 GND 0.004543f
C3451 VDD.n2774 GND 0.004543f
C3452 VDD.n2775 GND 0.004543f
C3453 VDD.n2776 GND 0.004543f
C3454 VDD.n2777 GND 0.004543f
C3455 VDD.n2778 GND 0.004543f
C3456 VDD.n2779 GND 0.004543f
C3457 VDD.n2780 GND 0.010421f
C3458 VDD.n2781 GND 0.010421f
C3459 VDD.n2782 GND 0.010421f
C3460 VDD.n2783 GND 0.010891f
C3461 VDD.n2784 GND 0.004543f
C3462 VDD.n2785 GND 0.004543f
C3463 VDD.n2786 GND 0.004543f
C3464 VDD.n2787 GND 0.004543f
C3465 VDD.n2788 GND 0.004543f
C3466 VDD.n2789 GND 0.004543f
C3467 VDD.t35 GND 0.077008f
C3468 VDD.t32 GND 0.389773f
C3469 VDD.n2790 GND 0.080451f
C3470 VDD.t34 GND 0.047872f
C3471 VDD.n2791 GND 0.076995f
C3472 VDD.n2792 GND 0.004543f
C3473 VDD.n2793 GND 0.004543f
C3474 VDD.n2794 GND 0.004543f
C3475 VDD.n2795 GND 0.004543f
C3476 VDD.n2796 GND 0.004543f
C3477 VDD.n2797 GND 0.004543f
C3478 VDD.n2798 GND 0.004543f
C3479 VDD.n2799 GND 0.004543f
C3480 VDD.n2800 GND 0.004543f
C3481 VDD.n2801 GND 0.004543f
C3482 VDD.n2802 GND 0.004543f
C3483 VDD.n2803 GND 0.004543f
C3484 VDD.n2804 GND 0.004543f
C3485 VDD.n2805 GND 0.004543f
C3486 VDD.n2806 GND 0.004543f
C3487 VDD.n2807 GND 0.004543f
C3488 VDD.n2808 GND 0.004543f
C3489 VDD.n2809 GND 0.004543f
C3490 VDD.n2810 GND 0.004543f
C3491 VDD.n2811 GND 0.004543f
C3492 VDD.n2812 GND 0.004543f
C3493 VDD.n2813 GND 0.004543f
C3494 VDD.n2814 GND 0.004543f
C3495 VDD.n2815 GND 0.004543f
C3496 VDD.n2816 GND 0.004543f
C3497 VDD.n2817 GND 0.004543f
C3498 VDD.n2818 GND 0.004543f
C3499 VDD.n2819 GND 0.004543f
C3500 VDD.n2820 GND 0.004543f
C3501 VDD.n2821 GND 0.004543f
C3502 VDD.n2822 GND 0.004543f
C3503 VDD.n2823 GND 0.004543f
C3504 VDD.n2824 GND 0.004543f
C3505 VDD.n2825 GND 0.004543f
C3506 VDD.n2826 GND 0.004543f
C3507 VDD.n2827 GND 0.004543f
C3508 VDD.n2828 GND 0.004543f
C3509 VDD.n2829 GND 0.004543f
C3510 VDD.n2830 GND 0.004543f
C3511 VDD.n2831 GND 0.004543f
C3512 VDD.n2832 GND 0.004543f
C3513 VDD.n2833 GND 0.004543f
C3514 VDD.n2834 GND 0.004543f
C3515 VDD.n2835 GND 0.004543f
C3516 VDD.n2836 GND 0.004543f
C3517 VDD.n2837 GND 0.004543f
C3518 VDD.n2838 GND 0.004543f
C3519 VDD.n2839 GND 0.004543f
C3520 VDD.n2840 GND 0.004543f
C3521 VDD.n2841 GND 0.004543f
C3522 VDD.n2842 GND 0.004543f
C3523 VDD.n2843 GND 0.004543f
C3524 VDD.n2844 GND 0.004543f
C3525 VDD.n2845 GND 0.004543f
C3526 VDD.n2846 GND 0.004543f
C3527 VDD.n2847 GND 0.004543f
C3528 VDD.n2848 GND 0.004543f
C3529 VDD.n2849 GND 0.004543f
C3530 VDD.n2850 GND 0.004543f
C3531 VDD.n2851 GND 0.004543f
C3532 VDD.n2852 GND 0.004543f
C3533 VDD.n2853 GND 0.004543f
C3534 VDD.n2854 GND 0.004543f
C3535 VDD.n2855 GND 0.004543f
C3536 VDD.n2856 GND 0.004543f
C3537 VDD.n2857 GND 0.004543f
C3538 VDD.n2858 GND 0.004543f
C3539 VDD.n2859 GND 0.004543f
C3540 VDD.n2860 GND 0.004543f
C3541 VDD.n2861 GND 0.004543f
C3542 VDD.n2862 GND 0.004543f
C3543 VDD.n2863 GND 0.004543f
C3544 VDD.n2864 GND 0.004543f
C3545 VDD.n2865 GND 0.004543f
C3546 VDD.n2866 GND 0.004543f
C3547 VDD.n2867 GND 0.004543f
C3548 VDD.n2868 GND 0.004543f
C3549 VDD.n2869 GND 0.004543f
C3550 VDD.n2870 GND 0.004543f
C3551 VDD.n2871 GND 0.004543f
C3552 VDD.n2872 GND 0.004543f
C3553 VDD.n2873 GND 0.004543f
C3554 VDD.n2874 GND 0.004543f
C3555 VDD.n2875 GND 0.004543f
C3556 VDD.n2876 GND 0.004543f
C3557 VDD.n2877 GND 0.004543f
C3558 VDD.n2878 GND 0.004543f
C3559 VDD.n2879 GND 0.004543f
C3560 VDD.n2880 GND 0.004543f
C3561 VDD.n2881 GND 0.004543f
C3562 VDD.n2882 GND 0.004543f
C3563 VDD.n2883 GND 0.004543f
C3564 VDD.n2884 GND 0.004543f
C3565 VDD.n2885 GND 0.004543f
C3566 VDD.n2886 GND 0.004543f
C3567 VDD.n2887 GND 0.004543f
C3568 VDD.n2888 GND 0.004543f
C3569 VDD.n2889 GND 0.004543f
C3570 VDD.n2890 GND 0.004543f
C3571 VDD.n2891 GND 0.004543f
C3572 VDD.n2892 GND 0.004543f
C3573 VDD.n2893 GND 0.004543f
C3574 VDD.n2894 GND 0.004543f
C3575 VDD.n2895 GND 0.004543f
C3576 VDD.n2896 GND 0.004543f
C3577 VDD.n2897 GND 0.004543f
C3578 VDD.n2898 GND 0.004543f
C3579 VDD.n2899 GND 0.004543f
C3580 VDD.n2900 GND 0.004543f
C3581 VDD.n2901 GND 0.004543f
C3582 VDD.n2902 GND 0.004543f
C3583 VDD.n2903 GND 0.004543f
C3584 VDD.n2904 GND 0.004543f
C3585 VDD.n2905 GND 0.004543f
C3586 VDD.n2906 GND 0.004543f
C3587 VDD.n2907 GND 0.004543f
C3588 VDD.n2908 GND 0.004543f
C3589 VDD.n2909 GND 0.004543f
C3590 VDD.n2910 GND 0.004543f
C3591 VDD.n2911 GND 0.004543f
C3592 VDD.n2912 GND 0.004543f
C3593 VDD.n2913 GND 0.004543f
C3594 VDD.n2914 GND 0.004543f
C3595 VDD.n2915 GND 0.004543f
C3596 VDD.n2916 GND 0.004543f
C3597 VDD.n2917 GND 0.004543f
C3598 VDD.n2918 GND 0.004543f
C3599 VDD.n2919 GND 0.004543f
C3600 VDD.n2920 GND 0.004543f
C3601 VDD.n2921 GND 0.004543f
C3602 VDD.n2922 GND 0.004543f
C3603 VDD.n2923 GND 0.004543f
C3604 VDD.n2924 GND 0.004543f
C3605 VDD.n2925 GND 0.004543f
C3606 VDD.n2926 GND 0.004543f
C3607 VDD.n2927 GND 0.004543f
C3608 VDD.n2928 GND 0.004543f
C3609 VDD.n2929 GND 0.004543f
C3610 VDD.n2930 GND 0.004543f
C3611 VDD.n2931 GND 0.004543f
C3612 VDD.n2932 GND 0.004543f
C3613 VDD.n2933 GND 0.004543f
C3614 VDD.n2934 GND 0.004543f
C3615 VDD.n2935 GND 0.004543f
C3616 VDD.n2936 GND 0.004543f
C3617 VDD.n2937 GND 0.004543f
C3618 VDD.n2938 GND 0.004543f
C3619 VDD.n2939 GND 0.004543f
C3620 VDD.n2940 GND 0.004543f
C3621 VDD.n2941 GND 0.004543f
C3622 VDD.n2942 GND 0.004543f
C3623 VDD.n2943 GND 0.004543f
C3624 VDD.n2944 GND 0.004543f
C3625 VDD.n2945 GND 0.004543f
C3626 VDD.n2946 GND 0.004543f
C3627 VDD.n2947 GND 0.004543f
C3628 VDD.n2948 GND 0.004543f
C3629 VDD.n2949 GND 0.004543f
C3630 VDD.n2950 GND 0.004543f
C3631 VDD.n2951 GND 0.004543f
C3632 VDD.n2952 GND 0.004543f
C3633 VDD.n2953 GND 0.004543f
C3634 VDD.n2954 GND 0.004543f
C3635 VDD.n2955 GND 0.004543f
C3636 VDD.n2956 GND 0.004543f
C3637 VDD.n2957 GND 0.004543f
C3638 VDD.n2958 GND 0.004543f
C3639 VDD.n2959 GND 0.004543f
C3640 VDD.n2960 GND 0.004543f
C3641 VDD.n2961 GND 0.004543f
C3642 VDD.n2962 GND 0.004543f
C3643 VDD.n2963 GND 0.004543f
C3644 VDD.n2964 GND 0.004543f
C3645 VDD.n2965 GND 0.004543f
C3646 VDD.n2966 GND 0.004543f
C3647 VDD.n2967 GND 0.004543f
C3648 VDD.n2968 GND 0.004543f
C3649 VDD.n2969 GND 0.004543f
C3650 VDD.n2970 GND 0.004543f
C3651 VDD.n2971 GND 0.004543f
C3652 VDD.n2972 GND 0.004543f
C3653 VDD.n2973 GND 0.004543f
C3654 VDD.n2974 GND 0.004543f
C3655 VDD.n2975 GND 0.004543f
C3656 VDD.n2976 GND 0.010421f
C3657 VDD.n2977 GND 0.010891f
C3658 VDD.n2978 GND 0.010891f
C3659 VDD.n2980 GND 0.004543f
C3660 VDD.n2982 GND 0.004543f
C3661 VDD.n2983 GND 0.004543f
C3662 VDD.n2984 GND 0.002773f
C3663 VDD.n2985 GND 0.005605f
C3664 VDD.n2986 GND 0.004042f
C3665 VDD.n2987 GND 0.004543f
C3666 VDD.n2989 GND 0.004543f
C3667 VDD.n2991 GND 0.004543f
C3668 VDD.n2992 GND 0.004543f
C3669 VDD.n2993 GND 0.004543f
C3670 VDD.n2994 GND 0.004543f
C3671 VDD.n2995 GND 0.004543f
C3672 VDD.n2997 GND 0.004543f
C3673 VDD.n2999 GND 0.004543f
C3674 VDD.n3000 GND 0.004543f
C3675 VDD.n3001 GND 0.004543f
C3676 VDD.n3002 GND 0.004543f
C3677 VDD.n3003 GND 0.004543f
C3678 VDD.n3005 GND 0.004543f
C3679 VDD.n3007 GND 0.004543f
C3680 VDD.n3008 GND 0.004543f
C3681 VDD.n3009 GND 0.010891f
C3682 VDD.n3010 GND 0.010421f
C3683 VDD.n3011 GND 0.010421f
C3684 VDD.n3012 GND 0.374096f
C3685 VDD.n3013 GND 0.010421f
C3686 VDD.n3014 GND 0.010421f
C3687 VDD.n3015 GND 0.004543f
C3688 VDD.n3016 GND 0.004543f
C3689 VDD.n3017 GND 0.004543f
C3690 VDD.n3018 GND 0.266372f
C3691 VDD.n3019 GND 0.004543f
C3692 VDD.n3020 GND 0.004543f
C3693 VDD.n3021 GND 0.004543f
C3694 VDD.n3022 GND 0.004543f
C3695 VDD.n3023 GND 0.004543f
C3696 VDD.n3024 GND 0.266372f
C3697 VDD.n3025 GND 0.004543f
C3698 VDD.n3026 GND 0.004543f
C3699 VDD.n3027 GND 0.004543f
C3700 VDD.n3028 GND 0.004543f
C3701 VDD.n3029 GND 0.004543f
C3702 VDD.n3030 GND 0.266372f
C3703 VDD.n3031 GND 0.004543f
C3704 VDD.n3032 GND 0.004543f
C3705 VDD.n3033 GND 0.004543f
C3706 VDD.n3034 GND 0.004543f
C3707 VDD.n3035 GND 0.004543f
C3708 VDD.n3036 GND 0.266372f
C3709 VDD.n3037 GND 0.004543f
C3710 VDD.n3038 GND 0.004543f
C3711 VDD.n3039 GND 0.004543f
C3712 VDD.n3040 GND 0.004543f
C3713 VDD.n3041 GND 0.004543f
C3714 VDD.n3042 GND 0.266372f
C3715 VDD.n3043 GND 0.004543f
C3716 VDD.n3044 GND 0.004543f
C3717 VDD.n3045 GND 0.004543f
C3718 VDD.n3046 GND 0.004543f
C3719 VDD.n3047 GND 0.004543f
C3720 VDD.n3048 GND 0.215448f
C3721 VDD.n3049 GND 0.004543f
C3722 VDD.n3050 GND 0.004543f
C3723 VDD.n3051 GND 0.004543f
C3724 VDD.n3052 GND 0.004543f
C3725 VDD.n3053 GND 0.004543f
C3726 VDD.n3054 GND 0.266372f
C3727 VDD.n3055 GND 0.004543f
C3728 VDD.n3056 GND 0.004543f
C3729 VDD.n3057 GND 0.004543f
C3730 VDD.n3058 GND 0.004543f
C3731 VDD.n3059 GND 0.004543f
C3732 VDD.n3060 GND 0.266372f
C3733 VDD.n3061 GND 0.004543f
C3734 VDD.n3062 GND 0.004543f
C3735 VDD.n3063 GND 0.004543f
C3736 VDD.n3064 GND 0.004543f
C3737 VDD.n3065 GND 0.004543f
C3738 VDD.n3066 GND 0.266372f
C3739 VDD.n3067 GND 0.004543f
C3740 VDD.n3068 GND 0.004543f
C3741 VDD.n3069 GND 0.004543f
C3742 VDD.n3070 GND 0.004543f
C3743 VDD.n3071 GND 0.004543f
C3744 VDD.n3072 GND 0.266372f
C3745 VDD.n3073 GND 0.004543f
C3746 VDD.n3074 GND 0.004543f
C3747 VDD.n3075 GND 0.004543f
C3748 VDD.n3076 GND 0.004543f
C3749 VDD.n3077 GND 0.004543f
C3750 VDD.n3078 GND 0.266372f
C3751 VDD.n3079 GND 0.004543f
C3752 VDD.n3080 GND 0.004543f
C3753 VDD.n3081 GND 0.004543f
C3754 VDD.n3082 GND 0.004543f
C3755 VDD.n3083 GND 0.004543f
C3756 VDD.n3084 GND 0.266372f
C3757 VDD.n3085 GND 0.004543f
C3758 VDD.n3086 GND 0.004543f
C3759 VDD.n3087 GND 0.004543f
C3760 VDD.n3088 GND 0.004543f
C3761 VDD.n3089 GND 0.004543f
C3762 VDD.n3090 GND 0.266372f
C3763 VDD.n3091 GND 0.004543f
C3764 VDD.n3092 GND 0.004543f
C3765 VDD.n3093 GND 0.004543f
C3766 VDD.n3094 GND 0.004543f
C3767 VDD.n3095 GND 0.004543f
C3768 VDD.n3096 GND 0.266372f
C3769 VDD.n3097 GND 0.004543f
C3770 VDD.n3098 GND 0.004543f
C3771 VDD.n3099 GND 0.004543f
C3772 VDD.n3100 GND 0.004543f
C3773 VDD.n3101 GND 0.004543f
C3774 VDD.n3102 GND 0.266372f
C3775 VDD.n3103 GND 0.004543f
C3776 VDD.n3104 GND 0.004543f
C3777 VDD.n3105 GND 0.004543f
C3778 VDD.n3106 GND 0.004543f
C3779 VDD.n3107 GND 0.004543f
C3780 VDD.n3108 GND 0.189986f
C3781 VDD.n3109 GND 0.004543f
C3782 VDD.n3110 GND 0.004543f
C3783 VDD.n3111 GND 0.004543f
C3784 VDD.n3112 GND 0.004543f
C3785 VDD.n3113 GND 0.004543f
C3786 VDD.n3114 GND 0.150813f
C3787 VDD.n3115 GND 0.004543f
C3788 VDD.n3116 GND 0.004543f
C3789 VDD.n3117 GND 0.004543f
C3790 VDD.n3118 GND 0.004543f
C3791 VDD.n3119 GND 0.004543f
C3792 VDD.n3120 GND 0.266372f
C3793 VDD.n3121 GND 0.004543f
C3794 VDD.n3122 GND 0.004543f
C3795 VDD.n3123 GND 0.004543f
C3796 VDD.n3124 GND 0.004543f
C3797 VDD.n3125 GND 0.004543f
C3798 VDD.n3126 GND 0.266372f
C3799 VDD.n3127 GND 0.004543f
C3800 VDD.n3128 GND 0.004543f
C3801 VDD.n3129 GND 0.004543f
C3802 VDD.n3130 GND 0.004543f
C3803 VDD.n3131 GND 0.004543f
C3804 VDD.n3132 GND 0.266372f
C3805 VDD.n3133 GND 0.004543f
C3806 VDD.n3134 GND 0.004543f
C3807 VDD.n3135 GND 0.004543f
C3808 VDD.n3136 GND 0.004543f
C3809 VDD.n3137 GND 0.004543f
C3810 VDD.n3138 GND 0.266372f
C3811 VDD.n3139 GND 0.004543f
C3812 VDD.n3140 GND 0.004543f
C3813 VDD.n3141 GND 0.004543f
C3814 VDD.n3142 GND 0.004543f
C3815 VDD.n3143 GND 0.004543f
C3816 VDD.n3144 GND 0.266372f
C3817 VDD.n3145 GND 0.004543f
C3818 VDD.n3146 GND 0.004543f
C3819 VDD.n3147 GND 0.004543f
C3820 VDD.n3148 GND 0.004543f
C3821 VDD.n3149 GND 0.004543f
C3822 VDD.n3150 GND 0.266372f
C3823 VDD.n3151 GND 0.004543f
C3824 VDD.n3152 GND 0.004543f
C3825 VDD.n3153 GND 0.004543f
C3826 VDD.n3154 GND 0.004543f
C3827 VDD.n3155 GND 0.004543f
C3828 VDD.n3156 GND 0.266372f
C3829 VDD.n3157 GND 0.004543f
C3830 VDD.n3158 GND 0.004543f
C3831 VDD.n3159 GND 0.004543f
C3832 VDD.n3160 GND 0.004543f
C3833 VDD.n3161 GND 0.004543f
C3834 VDD.n3162 GND 0.19782f
C3835 VDD.n3163 GND 0.004543f
C3836 VDD.n3164 GND 0.004543f
C3837 VDD.n3165 GND 0.004543f
C3838 VDD.n3166 GND 0.004543f
C3839 VDD.n3167 GND 0.004543f
C3840 VDD.n3168 GND 0.266372f
C3841 VDD.n3169 GND 0.004543f
C3842 VDD.n3170 GND 0.004543f
C3843 VDD.n3171 GND 0.004543f
C3844 VDD.n3172 GND 0.004543f
C3845 VDD.n3173 GND 0.004543f
C3846 VDD.n3174 GND 0.260496f
C3847 VDD.n3175 GND 0.004543f
C3848 VDD.n3176 GND 0.004543f
C3849 VDD.n3177 GND 0.004543f
C3850 VDD.n3178 GND 0.004543f
C3851 VDD.n3179 GND 0.004543f
C3852 VDD.n3180 GND 0.266372f
C3853 VDD.n3181 GND 0.004543f
C3854 VDD.n3182 GND 0.004543f
C3855 VDD.n3183 GND 0.004543f
C3856 VDD.n3184 GND 0.004543f
C3857 VDD.n3185 GND 0.004543f
C3858 VDD.n3186 GND 0.266372f
C3859 VDD.n3187 GND 0.004543f
C3860 VDD.n3188 GND 0.004543f
C3861 VDD.n3189 GND 0.004543f
C3862 VDD.n3190 GND 0.004543f
C3863 VDD.n3191 GND 0.004543f
C3864 VDD.n3192 GND 0.266372f
C3865 VDD.n3193 GND 0.004543f
C3866 VDD.n3194 GND 0.004543f
C3867 VDD.n3195 GND 0.004543f
C3868 VDD.n3196 GND 0.004543f
C3869 VDD.n3197 GND 0.004543f
C3870 VDD.n3198 GND 0.266372f
C3871 VDD.n3199 GND 0.004543f
C3872 VDD.n3200 GND 0.004543f
C3873 VDD.n3201 GND 0.004543f
C3874 VDD.n3202 GND 0.004543f
C3875 VDD.n3203 GND 0.004543f
C3876 VDD.n3204 GND 0.266372f
C3877 VDD.n3205 GND 0.004543f
C3878 VDD.n3206 GND 0.004543f
C3879 VDD.n3207 GND 0.004543f
C3880 VDD.n3208 GND 0.004543f
C3881 VDD.n3209 GND 0.004543f
C3882 VDD.n3210 GND 0.266372f
C3883 VDD.n3211 GND 0.004543f
C3884 VDD.n3212 GND 0.004543f
C3885 VDD.n3213 GND 0.004543f
C3886 VDD.n3214 GND 0.004543f
C3887 VDD.n3215 GND 0.004543f
C3888 VDD.n3216 GND 0.266372f
C3889 VDD.n3217 GND 0.004543f
C3890 VDD.n3218 GND 0.004543f
C3891 VDD.n3219 GND 0.004543f
C3892 VDD.n3220 GND 0.004543f
C3893 VDD.n3221 GND 0.004543f
C3894 VDD.n3222 GND 0.213489f
C3895 VDD.n3223 GND 0.004543f
C3896 VDD.n3224 GND 0.004543f
C3897 VDD.n3225 GND 0.004543f
C3898 VDD.n3226 GND 0.004543f
C3899 VDD.n3227 GND 0.004543f
C3900 VDD.n3228 GND 0.139062f
C3901 VDD.n3229 GND 0.004543f
C3902 VDD.n3230 GND 0.004543f
C3903 VDD.n3231 GND 0.004543f
C3904 VDD.n3232 GND 0.004543f
C3905 VDD.n3233 GND 0.004543f
C3906 VDD.n3234 GND 0.266372f
C3907 VDD.n3235 GND 0.004543f
C3908 VDD.n3236 GND 0.004543f
C3909 VDD.n3237 GND 0.004543f
C3910 VDD.n3238 GND 0.004543f
C3911 VDD.n3239 GND 0.004543f
C3912 VDD.n3240 GND 0.266372f
C3913 VDD.n3241 GND 0.004543f
C3914 VDD.n3242 GND 0.004543f
C3915 VDD.n3243 GND 0.004543f
C3916 VDD.n3244 GND 0.004543f
C3917 VDD.n3245 GND 0.004543f
C3918 VDD.n3246 GND 0.266372f
C3919 VDD.n3247 GND 0.004543f
C3920 VDD.n3248 GND 0.004543f
C3921 VDD.n3249 GND 0.004543f
C3922 VDD.n3250 GND 0.004543f
C3923 VDD.n3251 GND 0.004543f
C3924 VDD.n3252 GND 0.266372f
C3925 VDD.n3253 GND 0.004543f
C3926 VDD.n3254 GND 0.004543f
C3927 VDD.n3255 GND 0.004543f
C3928 VDD.n3256 GND 0.004543f
C3929 VDD.n3257 GND 0.004543f
C3930 VDD.n3258 GND 0.266372f
C3931 VDD.n3259 GND 0.004543f
C3932 VDD.n3260 GND 0.004543f
C3933 VDD.n3261 GND 0.004543f
C3934 VDD.n3262 GND 0.004543f
C3935 VDD.n3263 GND 0.004543f
C3936 VDD.n3264 GND 0.266372f
C3937 VDD.n3265 GND 0.004543f
C3938 VDD.n3266 GND 0.004543f
C3939 VDD.n3267 GND 0.004543f
C3940 VDD.n3268 GND 0.004543f
C3941 VDD.n3269 GND 0.004543f
C3942 VDD.n3270 GND 0.266372f
C3943 VDD.n3271 GND 0.004543f
C3944 VDD.n3272 GND 0.004543f
C3945 VDD.n3273 GND 0.004543f
C3946 VDD.n3274 GND 0.004543f
C3947 VDD.n3275 GND 0.004543f
C3948 VDD.n3276 GND 0.266372f
C3949 VDD.n3277 GND 0.004543f
C3950 VDD.n3278 GND 0.004543f
C3951 VDD.n3279 GND 0.004543f
C3952 VDD.n3280 GND 0.004543f
C3953 VDD.n3281 GND 0.004543f
C3954 VDD.n3282 GND 0.248744f
C3955 VDD.n3283 GND 0.004543f
C3956 VDD.n3284 GND 0.004543f
C3957 VDD.n3285 GND 0.004543f
C3958 VDD.n3286 GND 0.004543f
C3959 VDD.n3287 GND 0.004543f
C3960 VDD.n3288 GND 0.266372f
C3961 VDD.n3289 GND 0.004543f
C3962 VDD.n3290 GND 0.004543f
C3963 VDD.n3291 GND 0.004543f
C3964 VDD.n3292 GND 0.004543f
C3965 VDD.n3293 GND 0.004543f
C3966 VDD.n3294 GND 0.266372f
C3967 VDD.n3295 GND 0.004543f
C3968 VDD.n3296 GND 0.004543f
C3969 VDD.n3297 GND 0.004543f
C3970 VDD.n3298 GND 0.004543f
C3971 VDD.n3299 GND 0.004543f
C3972 VDD.n3300 GND 0.266372f
C3973 VDD.n3301 GND 0.004543f
C3974 VDD.n3302 GND 0.004543f
C3975 VDD.n3303 GND 0.004543f
C3976 VDD.n3304 GND 0.004543f
C3977 VDD.n3305 GND 0.004543f
C3978 VDD.n3306 GND 0.211531f
C3979 VDD.n3307 GND 0.004543f
C3980 VDD.n3308 GND 0.004543f
C3981 VDD.n3309 GND 0.004543f
C3982 VDD.n3310 GND 0.004543f
C3983 VDD.n3311 GND 0.004543f
C3984 VDD.n3312 GND 0.266372f
C3985 VDD.n3313 GND 0.004543f
C3986 VDD.n3314 GND 0.004543f
C3987 VDD.n3315 GND 0.004543f
C3988 VDD.n3316 GND 0.004543f
C3989 VDD.n3317 GND 0.004543f
C3990 VDD.n3318 GND 0.266372f
C3991 VDD.n3319 GND 0.004543f
C3992 VDD.n3320 GND 0.004543f
C3993 VDD.n3321 GND 0.004543f
C3994 VDD.n3322 GND 0.004543f
C3995 VDD.n3323 GND 0.004543f
C3996 VDD.n3324 GND 0.266372f
C3997 VDD.n3325 GND 0.004543f
C3998 VDD.n3326 GND 0.004543f
C3999 VDD.n3327 GND 0.004543f
C4000 VDD.n3328 GND 0.004543f
C4001 VDD.n3329 GND 0.004543f
C4002 VDD.n3330 GND 0.266372f
C4003 VDD.n3331 GND 0.004543f
C4004 VDD.n3332 GND 0.004543f
C4005 VDD.n3333 GND 0.004543f
C4006 VDD.n3334 GND 0.004543f
C4007 VDD.n3335 GND 0.004543f
C4008 VDD.n3336 GND 0.266372f
C4009 VDD.n3337 GND 0.004543f
C4010 VDD.n3338 GND 0.004543f
C4011 VDD.n3339 GND 0.004543f
C4012 VDD.n3340 GND 0.004543f
C4013 VDD.n3341 GND 0.004543f
C4014 VDD.n3342 GND 0.266372f
C4015 VDD.n3343 GND 0.004543f
C4016 VDD.n3344 GND 0.004543f
C4017 VDD.n3345 GND 0.004543f
C4018 VDD.n3346 GND 0.004543f
C4019 VDD.n3347 GND 0.004543f
C4020 VDD.n3348 GND 0.266372f
C4021 VDD.n3349 GND 0.004543f
C4022 VDD.n3350 GND 0.004543f
C4023 VDD.n3351 GND 0.004543f
C4024 VDD.n3352 GND 0.004543f
C4025 VDD.n3353 GND 0.004543f
C4026 VDD.n3354 GND 0.139062f
C4027 VDD.n3355 GND 0.004543f
C4028 VDD.n3356 GND 0.004543f
C4029 VDD.n3357 GND 0.004543f
C4030 VDD.n3358 GND 0.004543f
C4031 VDD.n3359 GND 0.004543f
C4032 VDD.n3360 GND 0.176275f
C4033 VDD.n3361 GND 0.004543f
C4034 VDD.n3362 GND 0.004543f
C4035 VDD.n3363 GND 0.004543f
C4036 VDD.n3364 GND 0.004543f
C4037 VDD.n3365 GND 0.004543f
C4038 VDD.n3366 GND 0.266372f
C4039 VDD.n3367 GND 0.004543f
C4040 VDD.n3368 GND 0.004543f
C4041 VDD.n3369 GND 0.004543f
C4042 VDD.n3370 GND 0.010891f
C4043 VDD.n3371 GND 0.004543f
C4044 VDD.n3372 GND 0.004543f
C4045 VDD.n3375 GND 0.004543f
C4046 VDD.n3376 GND 0.004543f
C4047 VDD.n3377 GND 0.004543f
C4048 VDD.n3378 GND 0.004543f
C4049 VDD.n3380 GND 0.004543f
C4050 VDD.n3381 GND 0.004543f
C4051 VDD.n3382 GND 0.004543f
C4052 VDD.n3383 GND 0.004543f
C4053 VDD.n3384 GND 0.004543f
C4054 VDD.n3385 GND 0.004543f
C4055 VDD.n3387 GND 0.010891f
C4056 VDD.n3388 GND 0.010421f
C4057 VDD.n3389 GND 0.010421f
C4058 VDD.n3390 GND 0.004543f
C4059 VDD.n3391 GND 0.004543f
C4060 VDD.n3392 GND 0.004543f
C4061 VDD.n3393 GND 0.004543f
C4062 VDD.n3394 GND 0.004543f
C4063 VDD.n3395 GND 0.004543f
C4064 VDD.n3396 GND 0.004543f
C4065 VDD.n3397 GND 0.266372f
C4066 VDD.n3398 GND 0.004543f
C4067 VDD.n3399 GND 0.004543f
C4068 VDD.n3400 GND 0.004543f
C4069 VDD.n3401 GND 0.004543f
C4070 VDD.n3402 GND 0.004543f
C4071 VDD.n3403 GND 0.266372f
C4072 VDD.n3404 GND 0.004543f
C4073 VDD.n3405 GND 0.004543f
C4074 VDD.n3406 GND 0.004543f
C4075 VDD.n3407 GND 0.004543f
C4076 VDD.n3408 GND 0.010956f
C4077 VDD.n3410 GND 0.010421f
C4078 VDD.n3411 GND 0.010891f
C4079 VDD.n3412 GND 0.010356f
C4080 VDD.n3413 GND 0.004543f
C4081 VDD.n3414 GND 0.004543f
C4082 VDD.n3415 GND 0.004543f
C4083 VDD.n3417 GND 0.004543f
C4084 VDD.n3418 GND 0.004543f
C4085 VDD.n3419 GND 0.004042f
C4086 VDD.n3420 GND 0.004543f
C4087 VDD.n3421 GND 0.004543f
C4088 VDD.n3422 GND 0.004543f
C4089 VDD.n3424 GND 0.004543f
C4090 VDD.n3425 GND 0.003407f
C4091 VDD.n3426 GND 0.004543f
C4092 VDD.n3428 GND 0.004543f
C4093 VDD.n3429 GND 0.004543f
C4094 VDD.n3430 GND 0.004543f
C4095 VDD.n3431 GND 0.004543f
C4096 VDD.n3432 GND 0.004543f
C4097 VDD.n3433 GND 0.004543f
C4098 VDD.n3435 GND 0.004543f
C4099 VDD.n3436 GND 0.004543f
C4100 VDD.n3438 GND 0.010891f
C4101 VDD.n3439 GND 0.010891f
C4102 VDD.n3440 GND 0.010421f
C4103 VDD.n3441 GND 0.004543f
C4104 VDD.n3442 GND 0.004543f
C4105 VDD.n3443 GND 0.266372f
C4106 VDD.n3444 GND 0.004543f
C4107 VDD.n3445 GND 0.004543f
C4108 VDD.n3446 GND 0.010956f
C4109 VDD.n3447 GND 0.010356f
C4110 VDD.n3448 GND 0.010891f
C4111 VDD.n3450 GND 0.004543f
C4112 VDD.n3451 GND 0.004543f
C4113 VDD.n3452 GND 0.004543f
C4114 VDD.n3453 GND 0.002773f
C4115 VDD.n3454 GND 0.005605f
C4116 VDD.n3455 GND 0.004042f
C4117 VDD.n3456 GND 0.004543f
C4118 VDD.n3458 GND 0.004543f
C4119 VDD.n3459 GND 0.004543f
C4120 VDD.n3461 GND 0.004543f
C4121 VDD.n3462 GND 0.003407f
C4122 VDD.n3463 GND 0.022417f
C4123 VDD.n3464 GND 1.23929f
C4124 VDD.n3465 GND 0.181794f
C4125 VDD.n3466 GND 0.026997f
C4126 VDD.n3467 GND 0.172144f
C4127 VDD.n3468 GND 0.002823f
C4128 VDD.n3469 GND 0.00294f
C4129 VDD.n3470 GND 0.00334f
C4130 VDD.n3471 GND 0.00334f
C4131 VDD.n3472 GND 0.005243f
C4132 VDD.n3473 GND 0.006681f
C4133 VDD.n3474 GND 0.006681f
C4134 VDD.n3475 GND 0.005377f
C4135 VDD.n3476 GND 0.005377f
C4136 VDD.n3477 GND 0.006681f
C4137 VDD.n3478 GND 0.006681f
C4138 VDD.n3479 GND 0.005377f
C4139 VDD.n3480 GND 0.005377f
C4140 VDD.n3481 GND 0.006681f
C4141 VDD.n3482 GND 0.006681f
C4142 VDD.n3483 GND 0.005377f
C4143 VDD.n3484 GND 0.005377f
C4144 VDD.n3485 GND 0.006681f
C4145 VDD.n3486 GND 0.006681f
C4146 VDD.n3487 GND 0.005377f
C4147 VDD.n3488 GND 0.005377f
C4148 VDD.n3489 GND 0.006681f
C4149 VDD.n3490 GND 0.006681f
C4150 VDD.n3491 GND 0.005377f
C4151 VDD.n3492 GND 0.005377f
C4152 VDD.n3493 GND 0.006681f
C4153 VDD.n3494 GND 0.006681f
C4154 VDD.n3495 GND 0.005377f
C4155 VDD.n3496 GND 0.006681f
C4156 VDD.n3497 GND 0.00492f
C4157 VDD.n3498 GND 0.010082f
C4158 VDD.n3499 GND 0.00406f
C4159 VDD.n3500 GND 0.006681f
C4160 VDD.n3501 GND 0.006681f
C4161 VDD.n3502 GND 0.005377f
C4162 VDD.n3503 GND 0.005377f
C4163 VDD.n3504 GND 0.006681f
C4164 VDD.n3505 GND 0.006681f
C4165 VDD.n3506 GND 0.005377f
C4166 VDD.n3507 GND 0.005377f
C4167 VDD.n3508 GND 0.006681f
C4168 VDD.n3509 GND 0.006681f
C4169 VDD.n3510 GND 0.005377f
C4170 VDD.n3511 GND 0.005377f
C4171 VDD.n3512 GND 0.006681f
C4172 VDD.n3513 GND 0.006681f
C4173 VDD.n3514 GND 0.005377f
C4174 VDD.n3515 GND 0.005377f
C4175 VDD.n3516 GND 0.005377f
C4176 VDD.n3517 GND 0.006681f
C4177 VDD.n3518 GND 3.30223f
C4178 VDD.n3520 GND 0.015143f
C4179 VDD.n3521 GND 0.004463f
C4180 VDD.n3522 GND 0.00294f
C4181 VDD.n3523 GND 1.48602f
C4182 VDD.n3524 GND 0.032885f
C4183 VDD.n3525 GND 0.009656f
C4184 VDD.n3526 GND 0.006681f
C4185 VDD.n3527 GND 0.005377f
C4186 VDD.n3528 GND 0.006681f
C4187 VDD.n3529 GND 0.391723f
C4188 VDD.n3530 GND 0.006681f
C4189 VDD.n3531 GND 0.005377f
C4190 VDD.n3532 GND 0.006681f
C4191 VDD.n3533 GND 0.006681f
C4192 VDD.n3534 GND 0.006681f
C4193 VDD.n3535 GND 0.005377f
C4194 VDD.n3536 GND 0.006681f
C4195 VDD.n3537 GND 0.391723f
C4196 VDD.n3538 GND 0.006681f
C4197 VDD.n3539 GND 0.005377f
C4198 VDD.n3540 GND 0.006681f
C4199 VDD.n3541 GND 0.006681f
C4200 VDD.n3542 GND 0.006681f
C4201 VDD.n3543 GND 0.005377f
C4202 VDD.n3544 GND 0.006681f
C4203 VDD.n3545 GND 0.264413f
C4204 VDD.n3546 GND 0.006681f
C4205 VDD.n3547 GND 0.005377f
C4206 VDD.n3548 GND 0.006681f
C4207 VDD.n3549 GND 0.006681f
C4208 VDD.n3550 GND 0.006681f
C4209 VDD.n3551 GND 0.005377f
C4210 VDD.n3552 GND 0.006681f
C4211 VDD.n3553 GND 0.391723f
C4212 VDD.n3554 GND 0.006681f
C4213 VDD.n3555 GND 0.005377f
C4214 VDD.n3556 GND 0.006681f
C4215 VDD.n3557 GND 0.006681f
C4216 VDD.n3558 GND 0.006681f
C4217 VDD.n3559 GND 0.005377f
C4218 VDD.n3560 GND 0.006681f
C4219 VDD.n3561 GND 0.391723f
C4220 VDD.n3562 GND 0.006681f
C4221 VDD.n3563 GND 0.005377f
C4222 VDD.n3564 GND 0.006681f
C4223 VDD.n3565 GND 0.006681f
C4224 VDD.n3566 GND 0.006681f
C4225 VDD.n3567 GND 0.005377f
C4226 VDD.n3568 GND 0.006681f
C4227 VDD.n3569 GND 0.391723f
C4228 VDD.n3570 GND 0.006681f
C4229 VDD.n3571 GND 0.005377f
C4230 VDD.n3572 GND 0.006681f
C4231 VDD.n3573 GND 0.006681f
C4232 VDD.n3574 GND 0.006681f
C4233 VDD.n3575 GND 0.005377f
C4234 VDD.n3576 GND 0.006681f
C4235 VDD.n3577 GND 0.391723f
C4236 VDD.n3578 GND 0.006681f
C4237 VDD.n3579 GND 0.005377f
C4238 VDD.n3580 GND 0.006681f
C4239 VDD.n3581 GND 0.006681f
C4240 VDD.n3582 GND 0.006681f
C4241 VDD.n3583 GND 0.006681f
C4242 VDD.n3584 GND 0.005377f
C4243 VDD.n3585 GND 0.005377f
C4244 VDD.n3586 GND 0.006681f
C4245 VDD.n3587 GND 0.391723f
C4246 VDD.n3588 GND 0.006681f
C4247 VDD.n3589 GND 0.005377f
C4248 VDD.n3590 GND 0.006681f
C4249 VDD.n3591 GND 0.006681f
C4250 VDD.n3592 GND 0.006681f
C4251 VDD.n3593 GND 0.005377f
C4252 VDD.n3594 GND 0.006681f
C4253 VDD.n3595 GND 0.338841f
C4254 VDD.n3596 GND 0.006681f
C4255 VDD.n3597 GND 0.006681f
C4256 VDD.n3598 GND 0.005377f
C4257 VDD.n3599 GND 0.006681f
C4258 VDD.n3600 GND 0.006681f
C4259 VDD.n3601 GND 0.006681f
C4260 VDD.n3602 GND 0.006681f
C4261 VDD.n3603 GND 0.006681f
C4262 VDD.n3604 GND 0.005377f
C4263 VDD.n3605 GND 0.005377f
C4264 VDD.n3606 GND 0.006681f
C4265 VDD.n3607 GND 0.391723f
C4266 VDD.n3608 GND 0.391723f
C4267 VDD.n3609 GND 0.006681f
C4268 VDD.n3610 GND 0.005377f
C4269 VDD.n3611 GND 0.006681f
C4270 VDD.n3612 GND 0.006681f
C4271 VDD.n3613 GND 0.006681f
C4272 VDD.n3614 GND 0.005377f
C4273 VDD.n3615 GND 0.006681f
C4274 VDD.n3616 GND 0.006681f
C4275 VDD.n3617 GND 0.391723f
C4276 VDD.n3618 GND 0.006681f
C4277 VDD.n3619 GND 0.006681f
C4278 VDD.n3620 GND 0.005377f
C4279 VDD.n3621 GND 0.005377f
C4280 VDD.n3622 GND 0.005377f
C4281 VDD.n3623 GND 0.006681f
C4282 VDD.n3624 GND 0.006681f
C4283 VDD.n3625 GND 0.006681f
C4284 VDD.n3626 GND 0.006681f
C4285 VDD.n3627 GND 0.005377f
C4286 VDD.n3628 GND 0.005377f
C4287 VDD.n3629 GND 0.005377f
C4288 VDD.n3630 GND 0.006681f
C4289 VDD.n3631 GND 0.006681f
C4290 VDD.n3632 GND 0.006681f
C4291 VDD.n3633 GND 0.006681f
C4292 VDD.n3634 GND 0.005377f
C4293 VDD.n3635 GND 0.005377f
C4294 VDD.n3636 GND 0.005377f
C4295 VDD.n3637 GND 0.006681f
C4296 VDD.n3638 GND 0.006681f
C4297 VDD.n3639 GND 0.006681f
C4298 VDD.n3640 GND 0.006681f
C4299 VDD.n3641 GND 0.005377f
C4300 VDD.n3642 GND 0.005377f
C4301 VDD.n3643 GND 0.005377f
C4302 VDD.n3644 GND 0.006681f
C4303 VDD.n3645 GND 0.006681f
C4304 VDD.n3646 GND 0.006681f
C4305 VDD.n3647 GND 0.006681f
C4306 VDD.n3648 GND 0.005377f
C4307 VDD.n3649 GND 0.005377f
C4308 VDD.n3650 GND 0.005377f
C4309 VDD.n3651 GND 0.006681f
C4310 VDD.n3652 GND 0.006681f
C4311 VDD.n3653 GND 0.006681f
C4312 VDD.n3654 GND 0.006681f
C4313 VDD.n3655 GND 0.005377f
C4314 VDD.n3656 GND 0.005377f
C4315 VDD.n3657 GND 0.004463f
C4316 VDD.n3658 GND 0.014921f
C4317 VDD.n3659 GND 0.015143f
C4318 VDD.n3660 GND 0.002823f
C4319 VDD.n3661 GND 0.015143f
C4320 VDD.n3663 GND 0.871584f
C4321 VDD.n3664 GND 0.522951f
C4322 VDD.n3665 GND 0.391723f
C4323 VDD.n3666 GND 0.006681f
C4324 VDD.n3667 GND 0.005377f
C4325 VDD.n3668 GND 0.005377f
C4326 VDD.n3669 GND 0.005377f
C4327 VDD.n3670 GND 0.006681f
C4328 VDD.n3671 GND 0.391723f
C4329 VDD.n3672 GND 0.391723f
C4330 VDD.n3673 GND 0.264413f
C4331 VDD.n3674 GND 0.006681f
C4332 VDD.n3675 GND 0.005377f
C4333 VDD.n3676 GND 0.005377f
C4334 VDD.n3677 GND 0.005377f
C4335 VDD.n3678 GND 0.006681f
C4336 VDD.n3679 GND 0.391723f
C4337 VDD.n3680 GND 0.391723f
C4338 VDD.n3681 GND 0.391723f
C4339 VDD.n3682 GND 0.006681f
C4340 VDD.n3683 GND 0.005377f
C4341 VDD.n3684 GND 0.005377f
C4342 VDD.n3685 GND 0.005377f
C4343 VDD.n3686 GND 0.006681f
C4344 VDD.n3687 GND 0.391723f
C4345 VDD.n3688 GND 0.391723f
C4346 VDD.n3689 GND 0.391723f
C4347 VDD.n3690 GND 0.006681f
C4348 VDD.n3691 GND 0.005377f
C4349 VDD.n3692 GND 0.005377f
C4350 VDD.n3693 GND 0.005377f
C4351 VDD.n3694 GND 0.006681f
C4352 VDD.n3695 GND 0.391723f
C4353 VDD.n3696 GND 0.391723f
C4354 VDD.n3697 GND 0.338841f
C4355 VDD.n3698 GND 0.006681f
C4356 VDD.n3699 GND 0.005377f
C4357 VDD.n3700 GND 0.005377f
C4358 VDD.n3701 GND 0.005377f
C4359 VDD.n3702 GND 0.006681f
C4360 VDD.n3703 GND 0.391723f
C4361 VDD.n3704 GND 0.391723f
C4362 VDD.n3705 GND 0.391723f
C4363 VDD.n3706 GND 0.006681f
C4364 VDD.n3707 GND 0.005377f
C4365 VDD.n3708 GND 0.005377f
C4366 VDD.n3709 GND 0.005135f
C4367 VDD.n3710 GND 0.40254f
C4368 VDD.n3711 GND 2.83965f
C4369 a_n11689_9690.n0 GND 7.92416f
C4370 a_n11689_9690.n1 GND 5.68564f
C4371 a_n11689_9690.t8 GND 0.068966f
C4372 a_n11689_9690.t5 GND 0.068966f
C4373 a_n11689_9690.t4 GND 0.068966f
C4374 a_n11689_9690.n2 GND 0.314677f
C4375 a_n11689_9690.t9 GND 0.068966f
C4376 a_n11689_9690.t10 GND 0.068966f
C4377 a_n11689_9690.n3 GND 0.287401f
C4378 a_n11689_9690.n4 GND 20.4885f
C4379 a_n11689_9690.t15 GND 0.350216f
C4380 a_n11689_9690.t12 GND 0.068966f
C4381 a_n11689_9690.t2 GND 0.068966f
C4382 a_n11689_9690.n5 GND 0.226949f
C4383 a_n11689_9690.t3 GND 0.333824f
C4384 a_n11689_9690.t14 GND 0.333824f
C4385 a_n11689_9690.t0 GND 0.068966f
C4386 a_n11689_9690.t13 GND 0.068966f
C4387 a_n11689_9690.n6 GND 0.226949f
C4388 a_n11689_9690.t1 GND 0.333824f
C4389 a_n11689_9690.n7 GND 6.94725f
C4390 a_n11689_9690.t7 GND 0.068966f
C4391 a_n11689_9690.t6 GND 0.068966f
C4392 a_n11689_9690.n8 GND 0.2874f
C4393 a_n11689_9690.n9 GND 9.61436f
C4394 a_n11689_9690.n10 GND 0.317411f
C4395 a_n11689_9690.t11 GND 0.068966f
C4396 a_n11545_9494.t28 GND 1.94323f
C4397 a_n11545_9494.t49 GND 1.8955f
C4398 a_n11545_9494.n0 GND 22.9935f
C4399 a_n11545_9494.n1 GND 7.96038f
C4400 a_n11545_9494.n2 GND 10.9607f
C4401 a_n11545_9494.t48 GND 1.94323f
C4402 a_n11545_9494.t51 GND 1.8955f
C4403 a_n11545_9494.t41 GND 1.94105f
C4404 a_n11545_9494.t32 GND 1.89583f
C4405 a_n11545_9494.t36 GND 1.94105f
C4406 a_n11545_9494.t50 GND 1.89583f
C4407 a_n11545_9494.n3 GND 5.34125f
C4408 a_n11545_9494.n4 GND 5.48553f
C4409 a_n11545_9494.n5 GND 0.898296f
C4410 a_n11545_9494.n6 GND 0.898296f
C4411 a_n11545_9494.n7 GND 5.46522f
C4412 a_n11545_9494.n8 GND 0.898296f
C4413 a_n11545_9494.t14 GND 1.9019f
C4414 a_n11545_9494.n9 GND 0.74751f
C4415 a_n11545_9494.t12 GND 2.09814f
C4416 a_n11545_9494.n10 GND 7.08247f
C4417 a_n11545_9494.t39 GND 2.09865f
C4418 a_n11545_9494.t24 GND 2.09865f
C4419 a_n11545_9494.t40 GND 2.09865f
C4420 a_n11545_9494.n11 GND 0.555058f
C4421 a_n11545_9494.n12 GND 13.646799f
C4422 a_n11545_9494.t35 GND 2.19451f
C4423 a_n11545_9494.t44 GND 2.19451f
C4424 a_n11545_9494.t38 GND 2.19451f
C4425 a_n11545_9494.t31 GND 2.19451f
C4426 a_n11545_9494.t18 GND 2.09772f
C4427 a_n11545_9494.t47 GND 1.94546f
C4428 a_n11545_9494.t33 GND 1.89517f
C4429 a_n11545_9494.t29 GND 2.11814f
C4430 a_n11545_9494.t25 GND 0.280208f
C4431 a_n11545_9494.t21 GND 0.05518f
C4432 a_n11545_9494.t17 GND 0.05518f
C4433 a_n11545_9494.n13 GND 0.181582f
C4434 a_n11545_9494.t11 GND 0.267092f
C4435 a_n11545_9494.t43 GND 2.11814f
C4436 a_n11545_9494.t34 GND 2.11814f
C4437 a_n11545_9494.t45 GND 2.11814f
C4438 a_n11545_9494.t46 GND 2.11814f
C4439 a_n11545_9494.t42 GND 1.94546f
C4440 a_n11545_9494.t37 GND 1.89517f
C4441 a_n11545_9494.t30 GND 2.11814f
C4442 a_n11545_9494.t20 GND 1.94546f
C4443 a_n11545_9494.t16 GND 1.89517f
C4444 a_n11545_9494.t10 GND 2.11814f
C4445 a_n11545_9494.t22 GND 1.21529f
C4446 a_n11545_9494.n14 GND 0.903114f
C4447 a_n11545_9494.t19 GND 0.280208f
C4448 a_n11545_9494.t15 GND 0.05518f
C4449 a_n11545_9494.t23 GND 0.05518f
C4450 a_n11545_9494.n15 GND 0.181582f
C4451 a_n11545_9494.t13 GND 0.267093f
C4452 a_n11545_9494.t1 GND 0.620358f
C4453 a_n11545_9494.t8 GND 0.077199f
C4454 a_n11545_9494.t3 GND 0.576643f
C4455 a_n11545_9494.t26 GND 0.077199f
C4456 a_n11545_9494.t4 GND 0.576643f
C4457 a_n11545_9494.t6 GND 0.077199f
C4458 a_n11545_9494.t5 GND 0.620358f
C4459 a_n11545_9494.t7 GND 0.077199f
C4460 a_n11545_9494.t9 GND 0.576643f
C4461 a_n11545_9494.t2 GND 0.077199f
C4462 a_n11545_9494.n16 GND 11.843599f
C4463 a_n11545_9494.t27 GND 0.620356f
C4464 a_n11545_9494.t0 GND 0.077199f
C4465 a_n7516_558.n0 GND 4.21682f
C4466 a_n7516_558.n1 GND 4.21682f
C4467 a_n7516_558.n2 GND 2.16822f
C4468 a_n7516_558.n3 GND 2.85011f
C4469 a_n7516_558.n4 GND 2.85011f
C4470 a_n7516_558.n5 GND 2.73908f
C4471 a_n7516_558.n6 GND 2.73908f
C4472 a_n7516_558.n7 GND 9.49142f
C4473 a_n7516_558.t10 GND 0.320083f
C4474 a_n7516_558.t12 GND 0.049842f
C4475 a_n7516_558.t9 GND 0.049842f
C4476 a_n7516_558.n8 GND 0.265103f
C4477 a_n7516_558.t22 GND 0.049842f
C4478 a_n7516_558.t4 GND 0.049842f
C4479 a_n7516_558.n9 GND 0.265103f
C4480 a_n7516_558.t14 GND 0.320083f
C4481 a_n7516_558.t6 GND 0.320083f
C4482 a_n7516_558.t2 GND 0.049842f
C4483 a_n7516_558.t0 GND 0.049842f
C4484 a_n7516_558.n10 GND 0.265103f
C4485 a_n7516_558.t21 GND 0.049842f
C4486 a_n7516_558.t17 GND 0.049842f
C4487 a_n7516_558.n11 GND 0.265103f
C4488 a_n7516_558.t20 GND 0.320082f
C4489 a_n7516_558.t19 GND 0.320082f
C4490 a_n7516_558.t18 GND 0.049842f
C4491 a_n7516_558.t7 GND 0.049842f
C4492 a_n7516_558.n12 GND 0.265102f
C4493 a_n7516_558.t1 GND 0.049842f
C4494 a_n7516_558.t5 GND 0.049842f
C4495 a_n7516_558.n13 GND 0.265102f
C4496 a_n7516_558.t16 GND 0.320082f
C4497 a_n7516_558.t11 GND 0.320082f
C4498 a_n7516_558.t13 GND 0.049842f
C4499 a_n7516_558.t15 GND 0.049842f
C4500 a_n7516_558.n14 GND 0.265102f
C4501 a_n7516_558.t8 GND 0.049842f
C4502 a_n7516_558.t3 GND 0.049842f
C4503 a_n7516_558.n15 GND 0.265102f
C4504 a_n7516_558.t25 GND 0.320082f
C4505 a_n7516_558.n16 GND 2.55745f
C4506 a_n7516_558.t23 GND 0.695968f
C4507 a_n7516_558.t24 GND 0.695968f
C4508 CS_BIAS.t50 GND 0.191402f
C4509 CS_BIAS.n0 GND 0.108818f
C4510 CS_BIAS.n1 GND 0.006836f
C4511 CS_BIAS.n2 GND 0.012677f
C4512 CS_BIAS.n3 GND 0.006836f
C4513 CS_BIAS.n4 GND 0.008132f
C4514 CS_BIAS.n5 GND 0.006836f
C4515 CS_BIAS.n6 GND 0.012677f
C4516 CS_BIAS.n7 GND 0.006836f
C4517 CS_BIAS.t43 GND 0.191402f
C4518 CS_BIAS.n8 GND 0.012677f
C4519 CS_BIAS.n9 GND 0.006836f
C4520 CS_BIAS.n10 GND 0.004099f
C4521 CS_BIAS.n11 GND 0.006836f
C4522 CS_BIAS.n12 GND 0.012677f
C4523 CS_BIAS.n13 GND 0.005972f
C4524 CS_BIAS.t58 GND 0.191402f
C4525 CS_BIAS.n14 GND 0.012677f
C4526 CS_BIAS.t14 GND 0.191402f
C4527 CS_BIAS.n15 GND 0.108818f
C4528 CS_BIAS.n16 GND 0.006836f
C4529 CS_BIAS.n17 GND 0.012677f
C4530 CS_BIAS.n18 GND 0.006836f
C4531 CS_BIAS.n19 GND 0.008132f
C4532 CS_BIAS.n20 GND 0.006836f
C4533 CS_BIAS.n21 GND 0.012677f
C4534 CS_BIAS.n22 GND 0.006836f
C4535 CS_BIAS.t18 GND 0.191402f
C4536 CS_BIAS.n23 GND 0.012677f
C4537 CS_BIAS.n24 GND 0.006836f
C4538 CS_BIAS.n25 GND 0.004099f
C4539 CS_BIAS.n26 GND 0.006836f
C4540 CS_BIAS.n27 GND 0.012677f
C4541 CS_BIAS.n28 GND 0.006836f
C4542 CS_BIAS.t2 GND 0.191402f
C4543 CS_BIAS.n29 GND 0.012677f
C4544 CS_BIAS.n30 GND 0.006836f
C4545 CS_BIAS.n31 GND 0.010554f
C4546 CS_BIAS.n32 GND 0.006836f
C4547 CS_BIAS.n33 GND 0.012677f
C4548 CS_BIAS.n34 GND 0.006836f
C4549 CS_BIAS.t16 GND 0.191402f
C4550 CS_BIAS.n35 GND 0.108333f
C4551 CS_BIAS.t0 GND 0.307989f
C4552 CS_BIAS.n36 GND 0.208121f
C4553 CS_BIAS.n37 GND 0.074665f
C4554 CS_BIAS.n38 GND 0.008046f
C4555 CS_BIAS.n39 GND 0.012677f
C4556 CS_BIAS.n40 GND 0.012677f
C4557 CS_BIAS.n41 GND 0.006836f
C4558 CS_BIAS.n42 GND 0.006836f
C4559 CS_BIAS.n43 GND 0.006836f
C4560 CS_BIAS.n44 GND 0.012677f
C4561 CS_BIAS.n45 GND 0.012419f
C4562 CS_BIAS.n46 GND 0.004099f
C4563 CS_BIAS.n47 GND 0.006836f
C4564 CS_BIAS.n48 GND 0.006836f
C4565 CS_BIAS.n49 GND 0.006836f
C4566 CS_BIAS.n50 GND 0.012677f
C4567 CS_BIAS.n51 GND 0.012677f
C4568 CS_BIAS.n52 GND 0.012677f
C4569 CS_BIAS.n53 GND 0.006836f
C4570 CS_BIAS.n54 GND 0.006836f
C4571 CS_BIAS.n55 GND 0.006836f
C4572 CS_BIAS.n56 GND 0.009548f
C4573 CS_BIAS.n57 GND 0.082235f
C4574 CS_BIAS.n58 GND 0.009548f
C4575 CS_BIAS.n59 GND 0.012677f
C4576 CS_BIAS.n60 GND 0.006836f
C4577 CS_BIAS.n61 GND 0.006836f
C4578 CS_BIAS.n62 GND 0.006836f
C4579 CS_BIAS.n63 GND 0.012677f
C4580 CS_BIAS.n64 GND 0.012677f
C4581 CS_BIAS.n65 GND 0.010554f
C4582 CS_BIAS.n66 GND 0.006836f
C4583 CS_BIAS.n67 GND 0.006836f
C4584 CS_BIAS.n68 GND 0.006836f
C4585 CS_BIAS.n69 GND 0.012419f
C4586 CS_BIAS.n70 GND 0.012677f
C4587 CS_BIAS.n71 GND 0.012677f
C4588 CS_BIAS.n72 GND 0.006836f
C4589 CS_BIAS.n73 GND 0.006836f
C4590 CS_BIAS.n74 GND 0.006836f
C4591 CS_BIAS.n75 GND 0.012677f
C4592 CS_BIAS.n76 GND 0.008046f
C4593 CS_BIAS.n77 GND 0.082235f
C4594 CS_BIAS.n78 GND 0.01105f
C4595 CS_BIAS.n79 GND 0.006836f
C4596 CS_BIAS.n80 GND 0.006836f
C4597 CS_BIAS.n81 GND 0.006836f
C4598 CS_BIAS.n82 GND 0.012677f
C4599 CS_BIAS.n83 GND 0.012677f
C4600 CS_BIAS.n84 GND 0.012904f
C4601 CS_BIAS.n85 GND 0.006836f
C4602 CS_BIAS.n86 GND 0.006836f
C4603 CS_BIAS.n87 GND 0.006836f
C4604 CS_BIAS.n88 GND 0.005106f
C4605 CS_BIAS.n89 GND 0.013606f
C4606 CS_BIAS.n90 GND 0.012677f
C4607 CS_BIAS.n91 GND 0.006836f
C4608 CS_BIAS.n92 GND 0.006836f
C4609 CS_BIAS.n93 GND 0.006836f
C4610 CS_BIAS.n94 GND 0.012677f
C4611 CS_BIAS.n95 GND 0.012677f
C4612 CS_BIAS.n96 GND 0.006544f
C4613 CS_BIAS.n97 GND 0.014459f
C4614 CS_BIAS.n98 GND 0.1106f
C4615 CS_BIAS.t15 GND 0.062866f
C4616 CS_BIAS.n99 GND 0.240076f
C4617 CS_BIAS.t19 GND 0.008767f
C4618 CS_BIAS.t3 GND 0.008767f
C4619 CS_BIAS.n100 GND 0.053984f
C4620 CS_BIAS.n101 GND 0.219488f
C4621 CS_BIAS.t17 GND 0.008767f
C4622 CS_BIAS.t1 GND 0.008767f
C4623 CS_BIAS.n102 GND 0.058552f
C4624 CS_BIAS.n103 GND 0.471682f
C4625 CS_BIAS.n104 GND 0.044243f
C4626 CS_BIAS.n105 GND 0.006836f
C4627 CS_BIAS.n106 GND 0.010554f
C4628 CS_BIAS.n107 GND 0.006836f
C4629 CS_BIAS.n108 GND 0.012677f
C4630 CS_BIAS.n109 GND 0.006836f
C4631 CS_BIAS.t44 GND 0.191402f
C4632 CS_BIAS.n110 GND 0.108333f
C4633 CS_BIAS.t62 GND 0.307989f
C4634 CS_BIAS.n111 GND 0.208121f
C4635 CS_BIAS.n112 GND 0.074665f
C4636 CS_BIAS.n113 GND 0.008046f
C4637 CS_BIAS.n114 GND 0.012677f
C4638 CS_BIAS.n115 GND 0.012677f
C4639 CS_BIAS.n116 GND 0.006836f
C4640 CS_BIAS.n117 GND 0.006836f
C4641 CS_BIAS.n118 GND 0.006836f
C4642 CS_BIAS.n119 GND 0.012677f
C4643 CS_BIAS.n120 GND 0.012419f
C4644 CS_BIAS.n121 GND 0.004099f
C4645 CS_BIAS.n122 GND 0.006836f
C4646 CS_BIAS.n123 GND 0.006836f
C4647 CS_BIAS.n124 GND 0.006836f
C4648 CS_BIAS.n125 GND 0.012677f
C4649 CS_BIAS.n126 GND 0.012677f
C4650 CS_BIAS.n127 GND 0.012677f
C4651 CS_BIAS.n128 GND 0.006836f
C4652 CS_BIAS.n129 GND 0.006836f
C4653 CS_BIAS.n130 GND 0.005972f
C4654 CS_BIAS.n131 GND 0.009548f
C4655 CS_BIAS.n132 GND 0.082235f
C4656 CS_BIAS.n133 GND 0.009548f
C4657 CS_BIAS.n134 GND 0.012677f
C4658 CS_BIAS.n135 GND 0.006836f
C4659 CS_BIAS.n136 GND 0.006836f
C4660 CS_BIAS.n137 GND 0.006836f
C4661 CS_BIAS.n138 GND 0.012677f
C4662 CS_BIAS.n139 GND 0.012677f
C4663 CS_BIAS.n140 GND 0.010554f
C4664 CS_BIAS.n141 GND 0.006836f
C4665 CS_BIAS.n142 GND 0.006836f
C4666 CS_BIAS.n143 GND 0.006836f
C4667 CS_BIAS.n144 GND 0.012419f
C4668 CS_BIAS.n145 GND 0.012677f
C4669 CS_BIAS.n146 GND 0.012677f
C4670 CS_BIAS.n147 GND 0.006836f
C4671 CS_BIAS.n148 GND 0.006836f
C4672 CS_BIAS.n149 GND 0.006836f
C4673 CS_BIAS.n150 GND 0.012677f
C4674 CS_BIAS.n151 GND 0.008046f
C4675 CS_BIAS.n152 GND 0.082235f
C4676 CS_BIAS.n153 GND 0.01105f
C4677 CS_BIAS.n154 GND 0.006836f
C4678 CS_BIAS.n155 GND 0.006836f
C4679 CS_BIAS.n156 GND 0.006836f
C4680 CS_BIAS.n157 GND 0.012677f
C4681 CS_BIAS.n158 GND 0.012677f
C4682 CS_BIAS.n159 GND 0.012904f
C4683 CS_BIAS.n160 GND 0.006836f
C4684 CS_BIAS.n161 GND 0.006836f
C4685 CS_BIAS.n162 GND 0.006836f
C4686 CS_BIAS.n163 GND 0.005106f
C4687 CS_BIAS.n164 GND 0.013606f
C4688 CS_BIAS.n165 GND 0.012677f
C4689 CS_BIAS.n166 GND 0.006836f
C4690 CS_BIAS.n167 GND 0.006836f
C4691 CS_BIAS.n168 GND 0.006836f
C4692 CS_BIAS.n169 GND 0.012677f
C4693 CS_BIAS.n170 GND 0.012677f
C4694 CS_BIAS.n171 GND 0.006544f
C4695 CS_BIAS.n172 GND 0.014459f
C4696 CS_BIAS.n173 GND 0.081113f
C4697 CS_BIAS.t42 GND 0.191402f
C4698 CS_BIAS.n174 GND 0.108818f
C4699 CS_BIAS.n175 GND 0.006836f
C4700 CS_BIAS.n176 GND 0.012677f
C4701 CS_BIAS.n177 GND 0.006836f
C4702 CS_BIAS.n178 GND 0.008132f
C4703 CS_BIAS.n179 GND 0.006836f
C4704 CS_BIAS.n180 GND 0.012677f
C4705 CS_BIAS.n181 GND 0.006836f
C4706 CS_BIAS.t48 GND 0.191402f
C4707 CS_BIAS.n182 GND 0.012677f
C4708 CS_BIAS.n183 GND 0.006836f
C4709 CS_BIAS.n184 GND 0.004099f
C4710 CS_BIAS.n185 GND 0.006836f
C4711 CS_BIAS.n186 GND 0.012677f
C4712 CS_BIAS.n187 GND 0.006836f
C4713 CS_BIAS.t32 GND 0.191402f
C4714 CS_BIAS.n188 GND 0.012677f
C4715 CS_BIAS.n189 GND 0.006836f
C4716 CS_BIAS.n190 GND 0.010554f
C4717 CS_BIAS.n191 GND 0.006836f
C4718 CS_BIAS.n192 GND 0.012677f
C4719 CS_BIAS.n193 GND 0.006836f
C4720 CS_BIAS.t61 GND 0.191402f
C4721 CS_BIAS.n194 GND 0.108333f
C4722 CS_BIAS.t49 GND 0.307989f
C4723 CS_BIAS.n195 GND 0.208121f
C4724 CS_BIAS.n196 GND 0.074665f
C4725 CS_BIAS.n197 GND 0.008046f
C4726 CS_BIAS.n198 GND 0.012677f
C4727 CS_BIAS.n199 GND 0.012677f
C4728 CS_BIAS.n200 GND 0.006836f
C4729 CS_BIAS.n201 GND 0.006836f
C4730 CS_BIAS.n202 GND 0.006836f
C4731 CS_BIAS.n203 GND 0.012677f
C4732 CS_BIAS.n204 GND 0.012419f
C4733 CS_BIAS.n205 GND 0.004099f
C4734 CS_BIAS.n206 GND 0.006836f
C4735 CS_BIAS.n207 GND 0.006836f
C4736 CS_BIAS.n208 GND 0.006836f
C4737 CS_BIAS.n209 GND 0.012677f
C4738 CS_BIAS.n210 GND 0.012677f
C4739 CS_BIAS.n211 GND 0.012677f
C4740 CS_BIAS.n212 GND 0.006836f
C4741 CS_BIAS.n213 GND 0.006836f
C4742 CS_BIAS.n214 GND 0.006836f
C4743 CS_BIAS.n215 GND 0.009548f
C4744 CS_BIAS.n216 GND 0.082235f
C4745 CS_BIAS.n217 GND 0.009548f
C4746 CS_BIAS.n218 GND 0.012677f
C4747 CS_BIAS.n219 GND 0.006836f
C4748 CS_BIAS.n220 GND 0.006836f
C4749 CS_BIAS.n221 GND 0.006836f
C4750 CS_BIAS.n222 GND 0.012677f
C4751 CS_BIAS.n223 GND 0.012677f
C4752 CS_BIAS.n224 GND 0.010554f
C4753 CS_BIAS.n225 GND 0.006836f
C4754 CS_BIAS.n226 GND 0.006836f
C4755 CS_BIAS.n227 GND 0.006836f
C4756 CS_BIAS.n228 GND 0.012419f
C4757 CS_BIAS.n229 GND 0.012677f
C4758 CS_BIAS.n230 GND 0.012677f
C4759 CS_BIAS.n231 GND 0.006836f
C4760 CS_BIAS.n232 GND 0.006836f
C4761 CS_BIAS.n233 GND 0.006836f
C4762 CS_BIAS.n234 GND 0.012677f
C4763 CS_BIAS.n235 GND 0.008046f
C4764 CS_BIAS.n236 GND 0.082235f
C4765 CS_BIAS.n237 GND 0.01105f
C4766 CS_BIAS.n238 GND 0.006836f
C4767 CS_BIAS.n239 GND 0.006836f
C4768 CS_BIAS.n240 GND 0.006836f
C4769 CS_BIAS.n241 GND 0.012677f
C4770 CS_BIAS.n242 GND 0.012677f
C4771 CS_BIAS.n243 GND 0.012904f
C4772 CS_BIAS.n244 GND 0.006836f
C4773 CS_BIAS.n245 GND 0.006836f
C4774 CS_BIAS.n246 GND 0.006836f
C4775 CS_BIAS.n247 GND 0.005106f
C4776 CS_BIAS.n248 GND 0.013606f
C4777 CS_BIAS.n249 GND 0.012677f
C4778 CS_BIAS.n250 GND 0.006836f
C4779 CS_BIAS.n251 GND 0.006836f
C4780 CS_BIAS.n252 GND 0.006836f
C4781 CS_BIAS.n253 GND 0.012677f
C4782 CS_BIAS.n254 GND 0.012677f
C4783 CS_BIAS.n255 GND 0.006544f
C4784 CS_BIAS.n256 GND 0.014459f
C4785 CS_BIAS.n257 GND 0.072784f
C4786 CS_BIAS.n258 GND 0.073774f
C4787 CS_BIAS.t69 GND 0.191402f
C4788 CS_BIAS.n259 GND 0.108818f
C4789 CS_BIAS.n260 GND 0.006836f
C4790 CS_BIAS.n261 GND 0.012677f
C4791 CS_BIAS.n262 GND 0.006836f
C4792 CS_BIAS.n263 GND 0.008132f
C4793 CS_BIAS.n264 GND 0.006836f
C4794 CS_BIAS.n265 GND 0.012677f
C4795 CS_BIAS.n266 GND 0.006836f
C4796 CS_BIAS.t39 GND 0.191402f
C4797 CS_BIAS.n267 GND 0.012677f
C4798 CS_BIAS.n268 GND 0.006836f
C4799 CS_BIAS.n269 GND 0.004099f
C4800 CS_BIAS.n270 GND 0.006836f
C4801 CS_BIAS.n271 GND 0.012677f
C4802 CS_BIAS.n272 GND 0.006836f
C4803 CS_BIAS.t30 GND 0.191402f
C4804 CS_BIAS.n273 GND 0.012677f
C4805 CS_BIAS.n274 GND 0.006836f
C4806 CS_BIAS.n275 GND 0.010554f
C4807 CS_BIAS.n276 GND 0.006836f
C4808 CS_BIAS.n277 GND 0.012677f
C4809 CS_BIAS.n278 GND 0.006836f
C4810 CS_BIAS.t53 GND 0.191402f
C4811 CS_BIAS.n279 GND 0.108333f
C4812 CS_BIAS.t47 GND 0.307989f
C4813 CS_BIAS.n280 GND 0.208121f
C4814 CS_BIAS.n281 GND 0.074665f
C4815 CS_BIAS.n282 GND 0.008046f
C4816 CS_BIAS.n283 GND 0.012677f
C4817 CS_BIAS.n284 GND 0.012677f
C4818 CS_BIAS.n285 GND 0.006836f
C4819 CS_BIAS.n286 GND 0.006836f
C4820 CS_BIAS.n287 GND 0.006836f
C4821 CS_BIAS.n288 GND 0.012677f
C4822 CS_BIAS.n289 GND 0.012419f
C4823 CS_BIAS.n290 GND 0.004099f
C4824 CS_BIAS.n291 GND 0.006836f
C4825 CS_BIAS.n292 GND 0.006836f
C4826 CS_BIAS.n293 GND 0.006836f
C4827 CS_BIAS.n294 GND 0.012677f
C4828 CS_BIAS.n295 GND 0.012677f
C4829 CS_BIAS.n296 GND 0.012677f
C4830 CS_BIAS.n297 GND 0.006836f
C4831 CS_BIAS.n298 GND 0.006836f
C4832 CS_BIAS.n299 GND 0.006836f
C4833 CS_BIAS.n300 GND 0.009548f
C4834 CS_BIAS.n301 GND 0.082235f
C4835 CS_BIAS.n302 GND 0.009548f
C4836 CS_BIAS.n303 GND 0.012677f
C4837 CS_BIAS.n304 GND 0.006836f
C4838 CS_BIAS.n305 GND 0.006836f
C4839 CS_BIAS.n306 GND 0.006836f
C4840 CS_BIAS.n307 GND 0.012677f
C4841 CS_BIAS.n308 GND 0.012677f
C4842 CS_BIAS.n309 GND 0.010554f
C4843 CS_BIAS.n310 GND 0.006836f
C4844 CS_BIAS.n311 GND 0.006836f
C4845 CS_BIAS.n312 GND 0.006836f
C4846 CS_BIAS.n313 GND 0.012419f
C4847 CS_BIAS.n314 GND 0.012677f
C4848 CS_BIAS.n315 GND 0.012677f
C4849 CS_BIAS.n316 GND 0.006836f
C4850 CS_BIAS.n317 GND 0.006836f
C4851 CS_BIAS.n318 GND 0.006836f
C4852 CS_BIAS.n319 GND 0.012677f
C4853 CS_BIAS.n320 GND 0.008046f
C4854 CS_BIAS.n321 GND 0.082235f
C4855 CS_BIAS.n322 GND 0.01105f
C4856 CS_BIAS.n323 GND 0.006836f
C4857 CS_BIAS.n324 GND 0.006836f
C4858 CS_BIAS.n325 GND 0.006836f
C4859 CS_BIAS.n326 GND 0.012677f
C4860 CS_BIAS.n327 GND 0.012677f
C4861 CS_BIAS.n328 GND 0.012904f
C4862 CS_BIAS.n329 GND 0.006836f
C4863 CS_BIAS.n330 GND 0.006836f
C4864 CS_BIAS.n331 GND 0.006836f
C4865 CS_BIAS.n332 GND 0.005106f
C4866 CS_BIAS.n333 GND 0.013606f
C4867 CS_BIAS.n334 GND 0.012677f
C4868 CS_BIAS.n335 GND 0.006836f
C4869 CS_BIAS.n336 GND 0.006836f
C4870 CS_BIAS.n337 GND 0.006836f
C4871 CS_BIAS.n338 GND 0.012677f
C4872 CS_BIAS.n339 GND 0.012677f
C4873 CS_BIAS.n340 GND 0.006544f
C4874 CS_BIAS.n341 GND 0.014459f
C4875 CS_BIAS.n342 GND 0.072784f
C4876 CS_BIAS.n343 GND 0.051747f
C4877 CS_BIAS.t68 GND 0.191402f
C4878 CS_BIAS.n344 GND 0.108818f
C4879 CS_BIAS.n345 GND 0.006836f
C4880 CS_BIAS.n346 GND 0.012677f
C4881 CS_BIAS.n347 GND 0.006836f
C4882 CS_BIAS.n348 GND 0.008132f
C4883 CS_BIAS.n349 GND 0.006836f
C4884 CS_BIAS.n350 GND 0.012677f
C4885 CS_BIAS.n351 GND 0.006836f
C4886 CS_BIAS.t38 GND 0.191402f
C4887 CS_BIAS.n352 GND 0.012677f
C4888 CS_BIAS.n353 GND 0.006836f
C4889 CS_BIAS.n354 GND 0.004099f
C4890 CS_BIAS.n355 GND 0.006836f
C4891 CS_BIAS.n356 GND 0.012677f
C4892 CS_BIAS.n357 GND 0.006836f
C4893 CS_BIAS.t29 GND 0.191402f
C4894 CS_BIAS.n358 GND 0.012677f
C4895 CS_BIAS.n359 GND 0.006836f
C4896 CS_BIAS.n360 GND 0.010554f
C4897 CS_BIAS.n361 GND 0.006836f
C4898 CS_BIAS.n362 GND 0.012677f
C4899 CS_BIAS.n363 GND 0.006836f
C4900 CS_BIAS.t52 GND 0.191402f
C4901 CS_BIAS.n364 GND 0.108333f
C4902 CS_BIAS.t46 GND 0.307989f
C4903 CS_BIAS.n365 GND 0.208121f
C4904 CS_BIAS.n366 GND 0.074665f
C4905 CS_BIAS.n367 GND 0.008046f
C4906 CS_BIAS.n368 GND 0.012677f
C4907 CS_BIAS.n369 GND 0.012677f
C4908 CS_BIAS.n370 GND 0.006836f
C4909 CS_BIAS.n371 GND 0.006836f
C4910 CS_BIAS.n372 GND 0.006836f
C4911 CS_BIAS.n373 GND 0.012677f
C4912 CS_BIAS.n374 GND 0.012419f
C4913 CS_BIAS.n375 GND 0.004099f
C4914 CS_BIAS.n376 GND 0.006836f
C4915 CS_BIAS.n377 GND 0.006836f
C4916 CS_BIAS.n378 GND 0.006836f
C4917 CS_BIAS.n379 GND 0.012677f
C4918 CS_BIAS.n380 GND 0.012677f
C4919 CS_BIAS.n381 GND 0.012677f
C4920 CS_BIAS.n382 GND 0.006836f
C4921 CS_BIAS.n383 GND 0.006836f
C4922 CS_BIAS.n384 GND 0.006836f
C4923 CS_BIAS.n385 GND 0.009548f
C4924 CS_BIAS.n386 GND 0.082235f
C4925 CS_BIAS.n387 GND 0.009548f
C4926 CS_BIAS.n388 GND 0.012677f
C4927 CS_BIAS.n389 GND 0.006836f
C4928 CS_BIAS.n390 GND 0.006836f
C4929 CS_BIAS.n391 GND 0.006836f
C4930 CS_BIAS.n392 GND 0.012677f
C4931 CS_BIAS.n393 GND 0.012677f
C4932 CS_BIAS.n394 GND 0.010554f
C4933 CS_BIAS.n395 GND 0.006836f
C4934 CS_BIAS.n396 GND 0.006836f
C4935 CS_BIAS.n397 GND 0.006836f
C4936 CS_BIAS.n398 GND 0.012419f
C4937 CS_BIAS.n399 GND 0.012677f
C4938 CS_BIAS.n400 GND 0.012677f
C4939 CS_BIAS.n401 GND 0.006836f
C4940 CS_BIAS.n402 GND 0.006836f
C4941 CS_BIAS.n403 GND 0.006836f
C4942 CS_BIAS.n404 GND 0.012677f
C4943 CS_BIAS.n405 GND 0.008046f
C4944 CS_BIAS.n406 GND 0.082235f
C4945 CS_BIAS.n407 GND 0.01105f
C4946 CS_BIAS.n408 GND 0.006836f
C4947 CS_BIAS.n409 GND 0.006836f
C4948 CS_BIAS.n410 GND 0.006836f
C4949 CS_BIAS.n411 GND 0.012677f
C4950 CS_BIAS.n412 GND 0.012677f
C4951 CS_BIAS.n413 GND 0.012904f
C4952 CS_BIAS.n414 GND 0.006836f
C4953 CS_BIAS.n415 GND 0.006836f
C4954 CS_BIAS.n416 GND 0.006836f
C4955 CS_BIAS.n417 GND 0.005106f
C4956 CS_BIAS.n418 GND 0.013606f
C4957 CS_BIAS.n419 GND 0.012677f
C4958 CS_BIAS.n420 GND 0.006836f
C4959 CS_BIAS.n421 GND 0.006836f
C4960 CS_BIAS.n422 GND 0.006836f
C4961 CS_BIAS.n423 GND 0.012677f
C4962 CS_BIAS.n424 GND 0.012677f
C4963 CS_BIAS.n425 GND 0.006544f
C4964 CS_BIAS.n426 GND 0.014459f
C4965 CS_BIAS.n427 GND 0.072784f
C4966 CS_BIAS.n428 GND 0.051747f
C4967 CS_BIAS.t67 GND 0.191402f
C4968 CS_BIAS.n429 GND 0.108818f
C4969 CS_BIAS.n430 GND 0.006836f
C4970 CS_BIAS.n431 GND 0.012677f
C4971 CS_BIAS.n432 GND 0.006836f
C4972 CS_BIAS.n433 GND 0.008132f
C4973 CS_BIAS.n434 GND 0.006836f
C4974 CS_BIAS.n435 GND 0.012677f
C4975 CS_BIAS.n436 GND 0.006836f
C4976 CS_BIAS.t36 GND 0.191402f
C4977 CS_BIAS.n437 GND 0.012677f
C4978 CS_BIAS.n438 GND 0.006836f
C4979 CS_BIAS.n439 GND 0.004099f
C4980 CS_BIAS.n440 GND 0.006836f
C4981 CS_BIAS.n441 GND 0.012677f
C4982 CS_BIAS.n442 GND 0.006836f
C4983 CS_BIAS.t26 GND 0.191402f
C4984 CS_BIAS.n443 GND 0.012677f
C4985 CS_BIAS.n444 GND 0.006836f
C4986 CS_BIAS.n445 GND 0.010554f
C4987 CS_BIAS.n446 GND 0.006836f
C4988 CS_BIAS.n447 GND 0.012677f
C4989 CS_BIAS.n448 GND 0.006836f
C4990 CS_BIAS.t51 GND 0.191402f
C4991 CS_BIAS.n449 GND 0.108333f
C4992 CS_BIAS.t45 GND 0.307989f
C4993 CS_BIAS.n450 GND 0.20812f
C4994 CS_BIAS.n451 GND 0.074665f
C4995 CS_BIAS.n452 GND 0.008046f
C4996 CS_BIAS.n453 GND 0.012677f
C4997 CS_BIAS.n454 GND 0.012677f
C4998 CS_BIAS.n455 GND 0.006836f
C4999 CS_BIAS.n456 GND 0.006836f
C5000 CS_BIAS.n457 GND 0.006836f
C5001 CS_BIAS.n458 GND 0.012677f
C5002 CS_BIAS.n459 GND 0.012419f
C5003 CS_BIAS.n460 GND 0.004099f
C5004 CS_BIAS.n461 GND 0.006836f
C5005 CS_BIAS.n462 GND 0.006836f
C5006 CS_BIAS.n463 GND 0.006836f
C5007 CS_BIAS.n464 GND 0.012677f
C5008 CS_BIAS.n465 GND 0.012677f
C5009 CS_BIAS.n466 GND 0.012677f
C5010 CS_BIAS.n467 GND 0.006836f
C5011 CS_BIAS.n468 GND 0.006836f
C5012 CS_BIAS.n469 GND 0.006836f
C5013 CS_BIAS.n470 GND 0.009548f
C5014 CS_BIAS.n471 GND 0.082235f
C5015 CS_BIAS.n472 GND 0.009548f
C5016 CS_BIAS.n473 GND 0.012677f
C5017 CS_BIAS.n474 GND 0.006836f
C5018 CS_BIAS.n475 GND 0.006836f
C5019 CS_BIAS.n476 GND 0.006836f
C5020 CS_BIAS.n477 GND 0.012677f
C5021 CS_BIAS.n478 GND 0.012677f
C5022 CS_BIAS.n479 GND 0.010554f
C5023 CS_BIAS.n480 GND 0.006836f
C5024 CS_BIAS.n481 GND 0.006836f
C5025 CS_BIAS.n482 GND 0.006836f
C5026 CS_BIAS.n483 GND 0.012419f
C5027 CS_BIAS.n484 GND 0.012677f
C5028 CS_BIAS.n485 GND 0.012677f
C5029 CS_BIAS.n486 GND 0.006836f
C5030 CS_BIAS.n487 GND 0.006836f
C5031 CS_BIAS.n488 GND 0.006836f
C5032 CS_BIAS.n489 GND 0.012677f
C5033 CS_BIAS.n490 GND 0.008046f
C5034 CS_BIAS.n491 GND 0.082235f
C5035 CS_BIAS.n492 GND 0.01105f
C5036 CS_BIAS.n493 GND 0.006836f
C5037 CS_BIAS.n494 GND 0.006836f
C5038 CS_BIAS.n495 GND 0.006836f
C5039 CS_BIAS.n496 GND 0.012677f
C5040 CS_BIAS.n497 GND 0.012677f
C5041 CS_BIAS.n498 GND 0.012904f
C5042 CS_BIAS.n499 GND 0.006836f
C5043 CS_BIAS.n500 GND 0.006836f
C5044 CS_BIAS.n501 GND 0.006836f
C5045 CS_BIAS.n502 GND 0.005106f
C5046 CS_BIAS.n503 GND 0.013606f
C5047 CS_BIAS.n504 GND 0.012677f
C5048 CS_BIAS.n505 GND 0.006836f
C5049 CS_BIAS.n506 GND 0.006836f
C5050 CS_BIAS.n507 GND 0.006836f
C5051 CS_BIAS.n508 GND 0.012677f
C5052 CS_BIAS.n509 GND 0.012677f
C5053 CS_BIAS.n510 GND 0.006544f
C5054 CS_BIAS.n511 GND 0.014459f
C5055 CS_BIAS.n512 GND 0.072784f
C5056 CS_BIAS.n513 GND 0.958771f
C5057 CS_BIAS.t55 GND 0.191402f
C5058 CS_BIAS.n514 GND 0.108818f
C5059 CS_BIAS.n515 GND 0.006836f
C5060 CS_BIAS.n516 GND 0.012677f
C5061 CS_BIAS.n517 GND 0.006836f
C5062 CS_BIAS.n518 GND 0.008132f
C5063 CS_BIAS.n519 GND 0.006836f
C5064 CS_BIAS.n520 GND 0.012677f
C5065 CS_BIAS.n521 GND 0.006836f
C5066 CS_BIAS.t33 GND 0.191402f
C5067 CS_BIAS.n522 GND 0.012677f
C5068 CS_BIAS.n523 GND 0.006836f
C5069 CS_BIAS.n524 GND 0.004099f
C5070 CS_BIAS.n525 GND 0.006836f
C5071 CS_BIAS.n526 GND 0.012677f
C5072 CS_BIAS.n527 GND 0.005972f
C5073 CS_BIAS.t54 GND 0.191402f
C5074 CS_BIAS.n528 GND 0.012677f
C5075 CS_BIAS.n529 GND 0.006836f
C5076 CS_BIAS.n530 GND 0.010554f
C5077 CS_BIAS.n531 GND 0.006836f
C5078 CS_BIAS.n532 GND 0.012677f
C5079 CS_BIAS.n533 GND 0.006836f
C5080 CS_BIAS.t23 GND 0.191402f
C5081 CS_BIAS.n534 GND 0.108333f
C5082 CS_BIAS.t24 GND 0.307989f
C5083 CS_BIAS.n535 GND 0.20812f
C5084 CS_BIAS.n536 GND 0.074665f
C5085 CS_BIAS.n537 GND 0.008046f
C5086 CS_BIAS.n538 GND 0.012677f
C5087 CS_BIAS.n539 GND 0.012677f
C5088 CS_BIAS.n540 GND 0.006836f
C5089 CS_BIAS.n541 GND 0.006836f
C5090 CS_BIAS.n542 GND 0.006836f
C5091 CS_BIAS.n543 GND 0.012677f
C5092 CS_BIAS.n544 GND 0.012419f
C5093 CS_BIAS.n545 GND 0.004099f
C5094 CS_BIAS.n546 GND 0.006836f
C5095 CS_BIAS.n547 GND 0.006836f
C5096 CS_BIAS.n548 GND 0.006836f
C5097 CS_BIAS.n549 GND 0.012677f
C5098 CS_BIAS.n550 GND 0.012677f
C5099 CS_BIAS.n551 GND 0.012677f
C5100 CS_BIAS.n552 GND 0.006836f
C5101 CS_BIAS.n553 GND 0.006836f
C5102 CS_BIAS.t11 GND 0.06625f
C5103 CS_BIAS.t13 GND 0.008767f
C5104 CS_BIAS.t7 GND 0.008767f
C5105 CS_BIAS.n554 GND 0.053984f
C5106 CS_BIAS.n555 GND 0.415208f
C5107 CS_BIAS.t4 GND 0.191402f
C5108 CS_BIAS.n556 GND 0.108818f
C5109 CS_BIAS.n557 GND 0.006836f
C5110 CS_BIAS.n558 GND 0.012677f
C5111 CS_BIAS.n559 GND 0.006836f
C5112 CS_BIAS.n560 GND 0.008132f
C5113 CS_BIAS.n561 GND 0.006836f
C5114 CS_BIAS.n562 GND 0.012677f
C5115 CS_BIAS.n563 GND 0.006836f
C5116 CS_BIAS.t8 GND 0.191402f
C5117 CS_BIAS.n564 GND 0.012677f
C5118 CS_BIAS.n565 GND 0.006836f
C5119 CS_BIAS.n566 GND 0.004099f
C5120 CS_BIAS.n567 GND 0.006836f
C5121 CS_BIAS.n568 GND 0.012677f
C5122 CS_BIAS.n569 GND 0.006836f
C5123 CS_BIAS.t6 GND 0.191402f
C5124 CS_BIAS.n570 GND 0.012677f
C5125 CS_BIAS.n571 GND 0.006836f
C5126 CS_BIAS.n572 GND 0.010554f
C5127 CS_BIAS.n573 GND 0.006836f
C5128 CS_BIAS.n574 GND 0.012677f
C5129 CS_BIAS.n575 GND 0.006836f
C5130 CS_BIAS.t12 GND 0.191402f
C5131 CS_BIAS.n576 GND 0.108333f
C5132 CS_BIAS.t10 GND 0.307989f
C5133 CS_BIAS.n577 GND 0.20812f
C5134 CS_BIAS.n578 GND 0.074665f
C5135 CS_BIAS.n579 GND 0.008046f
C5136 CS_BIAS.n580 GND 0.012677f
C5137 CS_BIAS.n581 GND 0.012677f
C5138 CS_BIAS.n582 GND 0.006836f
C5139 CS_BIAS.n583 GND 0.006836f
C5140 CS_BIAS.n584 GND 0.006836f
C5141 CS_BIAS.n585 GND 0.012677f
C5142 CS_BIAS.n586 GND 0.012419f
C5143 CS_BIAS.n587 GND 0.004099f
C5144 CS_BIAS.n588 GND 0.006836f
C5145 CS_BIAS.n589 GND 0.006836f
C5146 CS_BIAS.n590 GND 0.006836f
C5147 CS_BIAS.n591 GND 0.012677f
C5148 CS_BIAS.n592 GND 0.012677f
C5149 CS_BIAS.n593 GND 0.012677f
C5150 CS_BIAS.n594 GND 0.006836f
C5151 CS_BIAS.n595 GND 0.006836f
C5152 CS_BIAS.n596 GND 0.006836f
C5153 CS_BIAS.n597 GND 0.009548f
C5154 CS_BIAS.n598 GND 0.082235f
C5155 CS_BIAS.n599 GND 0.009548f
C5156 CS_BIAS.n600 GND 0.012677f
C5157 CS_BIAS.n601 GND 0.006836f
C5158 CS_BIAS.n602 GND 0.006836f
C5159 CS_BIAS.n603 GND 0.006836f
C5160 CS_BIAS.n604 GND 0.012677f
C5161 CS_BIAS.n605 GND 0.012677f
C5162 CS_BIAS.n606 GND 0.010554f
C5163 CS_BIAS.n607 GND 0.006836f
C5164 CS_BIAS.n608 GND 0.006836f
C5165 CS_BIAS.n609 GND 0.006836f
C5166 CS_BIAS.n610 GND 0.012419f
C5167 CS_BIAS.n611 GND 0.012677f
C5168 CS_BIAS.n612 GND 0.012677f
C5169 CS_BIAS.n613 GND 0.006836f
C5170 CS_BIAS.n614 GND 0.006836f
C5171 CS_BIAS.n615 GND 0.006836f
C5172 CS_BIAS.n616 GND 0.012677f
C5173 CS_BIAS.n617 GND 0.008046f
C5174 CS_BIAS.n618 GND 0.082235f
C5175 CS_BIAS.n619 GND 0.01105f
C5176 CS_BIAS.n620 GND 0.006836f
C5177 CS_BIAS.n621 GND 0.006836f
C5178 CS_BIAS.n622 GND 0.006836f
C5179 CS_BIAS.n623 GND 0.012677f
C5180 CS_BIAS.n624 GND 0.012677f
C5181 CS_BIAS.n625 GND 0.012904f
C5182 CS_BIAS.n626 GND 0.006836f
C5183 CS_BIAS.n627 GND 0.006836f
C5184 CS_BIAS.n628 GND 0.006836f
C5185 CS_BIAS.n629 GND 0.005106f
C5186 CS_BIAS.n630 GND 0.013606f
C5187 CS_BIAS.n631 GND 0.012677f
C5188 CS_BIAS.n632 GND 0.006836f
C5189 CS_BIAS.n633 GND 0.006836f
C5190 CS_BIAS.n634 GND 0.006836f
C5191 CS_BIAS.n635 GND 0.012677f
C5192 CS_BIAS.n636 GND 0.012677f
C5193 CS_BIAS.n637 GND 0.006544f
C5194 CS_BIAS.n638 GND 0.014459f
C5195 CS_BIAS.n639 GND 0.119149f
C5196 CS_BIAS.t9 GND 0.008767f
C5197 CS_BIAS.t5 GND 0.008767f
C5198 CS_BIAS.n640 GND 0.053984f
C5199 CS_BIAS.n641 GND 0.326024f
C5200 CS_BIAS.n642 GND 0.182649f
C5201 CS_BIAS.n643 GND 0.044243f
C5202 CS_BIAS.n644 GND 0.005972f
C5203 CS_BIAS.n645 GND 0.009548f
C5204 CS_BIAS.n646 GND 0.082235f
C5205 CS_BIAS.n647 GND 0.009548f
C5206 CS_BIAS.n648 GND 0.012677f
C5207 CS_BIAS.n649 GND 0.006836f
C5208 CS_BIAS.n650 GND 0.006836f
C5209 CS_BIAS.n651 GND 0.006836f
C5210 CS_BIAS.n652 GND 0.012677f
C5211 CS_BIAS.n653 GND 0.012677f
C5212 CS_BIAS.n654 GND 0.010554f
C5213 CS_BIAS.n655 GND 0.006836f
C5214 CS_BIAS.n656 GND 0.006836f
C5215 CS_BIAS.n657 GND 0.006836f
C5216 CS_BIAS.n658 GND 0.012419f
C5217 CS_BIAS.n659 GND 0.012677f
C5218 CS_BIAS.n660 GND 0.012677f
C5219 CS_BIAS.n661 GND 0.006836f
C5220 CS_BIAS.n662 GND 0.006836f
C5221 CS_BIAS.n663 GND 0.006836f
C5222 CS_BIAS.n664 GND 0.012677f
C5223 CS_BIAS.n665 GND 0.008046f
C5224 CS_BIAS.n666 GND 0.082235f
C5225 CS_BIAS.n667 GND 0.01105f
C5226 CS_BIAS.n668 GND 0.006836f
C5227 CS_BIAS.n669 GND 0.006836f
C5228 CS_BIAS.n670 GND 0.006836f
C5229 CS_BIAS.n671 GND 0.012677f
C5230 CS_BIAS.n672 GND 0.012677f
C5231 CS_BIAS.n673 GND 0.012904f
C5232 CS_BIAS.n674 GND 0.006836f
C5233 CS_BIAS.n675 GND 0.006836f
C5234 CS_BIAS.n676 GND 0.006836f
C5235 CS_BIAS.n677 GND 0.005106f
C5236 CS_BIAS.n678 GND 0.013606f
C5237 CS_BIAS.n679 GND 0.012677f
C5238 CS_BIAS.n680 GND 0.006836f
C5239 CS_BIAS.n681 GND 0.006836f
C5240 CS_BIAS.n682 GND 0.006836f
C5241 CS_BIAS.n683 GND 0.012677f
C5242 CS_BIAS.n684 GND 0.012677f
C5243 CS_BIAS.n685 GND 0.006544f
C5244 CS_BIAS.n686 GND 0.014459f
C5245 CS_BIAS.n687 GND 0.081113f
C5246 CS_BIAS.t25 GND 0.191402f
C5247 CS_BIAS.n688 GND 0.108818f
C5248 CS_BIAS.n689 GND 0.006836f
C5249 CS_BIAS.n690 GND 0.012677f
C5250 CS_BIAS.n691 GND 0.006836f
C5251 CS_BIAS.n692 GND 0.008132f
C5252 CS_BIAS.n693 GND 0.006836f
C5253 CS_BIAS.n694 GND 0.012677f
C5254 CS_BIAS.n695 GND 0.006836f
C5255 CS_BIAS.t56 GND 0.191402f
C5256 CS_BIAS.n696 GND 0.012677f
C5257 CS_BIAS.n697 GND 0.006836f
C5258 CS_BIAS.n698 GND 0.004099f
C5259 CS_BIAS.n699 GND 0.006836f
C5260 CS_BIAS.n700 GND 0.012677f
C5261 CS_BIAS.n701 GND 0.006836f
C5262 CS_BIAS.t34 GND 0.191402f
C5263 CS_BIAS.n702 GND 0.012677f
C5264 CS_BIAS.n703 GND 0.006836f
C5265 CS_BIAS.n704 GND 0.010554f
C5266 CS_BIAS.n705 GND 0.006836f
C5267 CS_BIAS.n706 GND 0.012677f
C5268 CS_BIAS.n707 GND 0.006836f
C5269 CS_BIAS.t64 GND 0.191402f
C5270 CS_BIAS.n708 GND 0.108333f
C5271 CS_BIAS.t35 GND 0.307989f
C5272 CS_BIAS.n709 GND 0.20812f
C5273 CS_BIAS.n710 GND 0.074665f
C5274 CS_BIAS.n711 GND 0.008046f
C5275 CS_BIAS.n712 GND 0.012677f
C5276 CS_BIAS.n713 GND 0.012677f
C5277 CS_BIAS.n714 GND 0.006836f
C5278 CS_BIAS.n715 GND 0.006836f
C5279 CS_BIAS.n716 GND 0.006836f
C5280 CS_BIAS.n717 GND 0.012677f
C5281 CS_BIAS.n718 GND 0.012419f
C5282 CS_BIAS.n719 GND 0.004099f
C5283 CS_BIAS.n720 GND 0.006836f
C5284 CS_BIAS.n721 GND 0.006836f
C5285 CS_BIAS.n722 GND 0.006836f
C5286 CS_BIAS.n723 GND 0.012677f
C5287 CS_BIAS.n724 GND 0.012677f
C5288 CS_BIAS.n725 GND 0.012677f
C5289 CS_BIAS.n726 GND 0.006836f
C5290 CS_BIAS.n727 GND 0.006836f
C5291 CS_BIAS.n728 GND 0.006836f
C5292 CS_BIAS.n729 GND 0.009548f
C5293 CS_BIAS.n730 GND 0.082235f
C5294 CS_BIAS.n731 GND 0.009548f
C5295 CS_BIAS.n732 GND 0.012677f
C5296 CS_BIAS.n733 GND 0.006836f
C5297 CS_BIAS.n734 GND 0.006836f
C5298 CS_BIAS.n735 GND 0.006836f
C5299 CS_BIAS.n736 GND 0.012677f
C5300 CS_BIAS.n737 GND 0.012677f
C5301 CS_BIAS.n738 GND 0.010554f
C5302 CS_BIAS.n739 GND 0.006836f
C5303 CS_BIAS.n740 GND 0.006836f
C5304 CS_BIAS.n741 GND 0.006836f
C5305 CS_BIAS.n742 GND 0.012419f
C5306 CS_BIAS.n743 GND 0.012677f
C5307 CS_BIAS.n744 GND 0.012677f
C5308 CS_BIAS.n745 GND 0.006836f
C5309 CS_BIAS.n746 GND 0.006836f
C5310 CS_BIAS.n747 GND 0.006836f
C5311 CS_BIAS.n748 GND 0.012677f
C5312 CS_BIAS.n749 GND 0.008046f
C5313 CS_BIAS.n750 GND 0.082235f
C5314 CS_BIAS.n751 GND 0.01105f
C5315 CS_BIAS.n752 GND 0.006836f
C5316 CS_BIAS.n753 GND 0.006836f
C5317 CS_BIAS.n754 GND 0.006836f
C5318 CS_BIAS.n755 GND 0.012677f
C5319 CS_BIAS.n756 GND 0.012677f
C5320 CS_BIAS.n757 GND 0.012904f
C5321 CS_BIAS.n758 GND 0.006836f
C5322 CS_BIAS.n759 GND 0.006836f
C5323 CS_BIAS.n760 GND 0.006836f
C5324 CS_BIAS.n761 GND 0.005106f
C5325 CS_BIAS.n762 GND 0.013606f
C5326 CS_BIAS.n763 GND 0.012677f
C5327 CS_BIAS.n764 GND 0.006836f
C5328 CS_BIAS.n765 GND 0.006836f
C5329 CS_BIAS.n766 GND 0.006836f
C5330 CS_BIAS.n767 GND 0.012677f
C5331 CS_BIAS.n768 GND 0.012677f
C5332 CS_BIAS.n769 GND 0.006544f
C5333 CS_BIAS.n770 GND 0.014459f
C5334 CS_BIAS.n771 GND 0.072784f
C5335 CS_BIAS.n772 GND 0.073774f
C5336 CS_BIAS.t40 GND 0.191402f
C5337 CS_BIAS.n773 GND 0.108818f
C5338 CS_BIAS.n774 GND 0.006836f
C5339 CS_BIAS.n775 GND 0.012677f
C5340 CS_BIAS.n776 GND 0.006836f
C5341 CS_BIAS.n777 GND 0.008132f
C5342 CS_BIAS.n778 GND 0.006836f
C5343 CS_BIAS.n779 GND 0.012677f
C5344 CS_BIAS.n780 GND 0.006836f
C5345 CS_BIAS.t31 GND 0.191402f
C5346 CS_BIAS.n781 GND 0.012677f
C5347 CS_BIAS.n782 GND 0.006836f
C5348 CS_BIAS.n783 GND 0.004099f
C5349 CS_BIAS.n784 GND 0.006836f
C5350 CS_BIAS.n785 GND 0.012677f
C5351 CS_BIAS.n786 GND 0.006836f
C5352 CS_BIAS.t22 GND 0.191402f
C5353 CS_BIAS.n787 GND 0.012677f
C5354 CS_BIAS.n788 GND 0.006836f
C5355 CS_BIAS.n789 GND 0.010554f
C5356 CS_BIAS.n790 GND 0.006836f
C5357 CS_BIAS.n791 GND 0.012677f
C5358 CS_BIAS.n792 GND 0.006836f
C5359 CS_BIAS.t60 GND 0.191402f
C5360 CS_BIAS.n793 GND 0.108333f
C5361 CS_BIAS.t65 GND 0.307989f
C5362 CS_BIAS.n794 GND 0.20812f
C5363 CS_BIAS.n795 GND 0.074665f
C5364 CS_BIAS.n796 GND 0.008046f
C5365 CS_BIAS.n797 GND 0.012677f
C5366 CS_BIAS.n798 GND 0.012677f
C5367 CS_BIAS.n799 GND 0.006836f
C5368 CS_BIAS.n800 GND 0.006836f
C5369 CS_BIAS.n801 GND 0.006836f
C5370 CS_BIAS.n802 GND 0.012677f
C5371 CS_BIAS.n803 GND 0.012419f
C5372 CS_BIAS.n804 GND 0.004099f
C5373 CS_BIAS.n805 GND 0.006836f
C5374 CS_BIAS.n806 GND 0.006836f
C5375 CS_BIAS.n807 GND 0.006836f
C5376 CS_BIAS.n808 GND 0.012677f
C5377 CS_BIAS.n809 GND 0.012677f
C5378 CS_BIAS.n810 GND 0.012677f
C5379 CS_BIAS.n811 GND 0.006836f
C5380 CS_BIAS.n812 GND 0.006836f
C5381 CS_BIAS.n813 GND 0.006836f
C5382 CS_BIAS.n814 GND 0.009548f
C5383 CS_BIAS.n815 GND 0.082235f
C5384 CS_BIAS.n816 GND 0.009548f
C5385 CS_BIAS.n817 GND 0.012677f
C5386 CS_BIAS.n818 GND 0.006836f
C5387 CS_BIAS.n819 GND 0.006836f
C5388 CS_BIAS.n820 GND 0.006836f
C5389 CS_BIAS.n821 GND 0.012677f
C5390 CS_BIAS.n822 GND 0.012677f
C5391 CS_BIAS.n823 GND 0.010554f
C5392 CS_BIAS.n824 GND 0.006836f
C5393 CS_BIAS.n825 GND 0.006836f
C5394 CS_BIAS.n826 GND 0.006836f
C5395 CS_BIAS.n827 GND 0.012419f
C5396 CS_BIAS.n828 GND 0.012677f
C5397 CS_BIAS.n829 GND 0.012677f
C5398 CS_BIAS.n830 GND 0.006836f
C5399 CS_BIAS.n831 GND 0.006836f
C5400 CS_BIAS.n832 GND 0.006836f
C5401 CS_BIAS.n833 GND 0.012677f
C5402 CS_BIAS.n834 GND 0.008046f
C5403 CS_BIAS.n835 GND 0.082235f
C5404 CS_BIAS.n836 GND 0.01105f
C5405 CS_BIAS.n837 GND 0.006836f
C5406 CS_BIAS.n838 GND 0.006836f
C5407 CS_BIAS.n839 GND 0.006836f
C5408 CS_BIAS.n840 GND 0.012677f
C5409 CS_BIAS.n841 GND 0.012677f
C5410 CS_BIAS.n842 GND 0.012904f
C5411 CS_BIAS.n843 GND 0.006836f
C5412 CS_BIAS.n844 GND 0.006836f
C5413 CS_BIAS.n845 GND 0.006836f
C5414 CS_BIAS.n846 GND 0.005106f
C5415 CS_BIAS.n847 GND 0.013606f
C5416 CS_BIAS.n848 GND 0.012677f
C5417 CS_BIAS.n849 GND 0.006836f
C5418 CS_BIAS.n850 GND 0.006836f
C5419 CS_BIAS.n851 GND 0.006836f
C5420 CS_BIAS.n852 GND 0.012677f
C5421 CS_BIAS.n853 GND 0.012677f
C5422 CS_BIAS.n854 GND 0.006544f
C5423 CS_BIAS.n855 GND 0.014459f
C5424 CS_BIAS.n856 GND 0.072784f
C5425 CS_BIAS.n857 GND 0.051747f
C5426 CS_BIAS.t41 GND 0.191402f
C5427 CS_BIAS.n858 GND 0.108818f
C5428 CS_BIAS.n859 GND 0.006836f
C5429 CS_BIAS.n860 GND 0.012677f
C5430 CS_BIAS.n861 GND 0.006836f
C5431 CS_BIAS.n862 GND 0.008132f
C5432 CS_BIAS.n863 GND 0.006836f
C5433 CS_BIAS.n864 GND 0.012677f
C5434 CS_BIAS.n865 GND 0.006836f
C5435 CS_BIAS.t27 GND 0.191402f
C5436 CS_BIAS.n866 GND 0.012677f
C5437 CS_BIAS.n867 GND 0.006836f
C5438 CS_BIAS.n868 GND 0.004099f
C5439 CS_BIAS.n869 GND 0.006836f
C5440 CS_BIAS.n870 GND 0.012677f
C5441 CS_BIAS.n871 GND 0.006836f
C5442 CS_BIAS.t20 GND 0.191402f
C5443 CS_BIAS.n872 GND 0.012677f
C5444 CS_BIAS.n873 GND 0.006836f
C5445 CS_BIAS.n874 GND 0.010554f
C5446 CS_BIAS.n875 GND 0.006836f
C5447 CS_BIAS.n876 GND 0.012677f
C5448 CS_BIAS.n877 GND 0.006836f
C5449 CS_BIAS.t59 GND 0.191402f
C5450 CS_BIAS.n878 GND 0.108333f
C5451 CS_BIAS.t66 GND 0.307989f
C5452 CS_BIAS.n879 GND 0.20812f
C5453 CS_BIAS.n880 GND 0.074665f
C5454 CS_BIAS.n881 GND 0.008046f
C5455 CS_BIAS.n882 GND 0.012677f
C5456 CS_BIAS.n883 GND 0.012677f
C5457 CS_BIAS.n884 GND 0.006836f
C5458 CS_BIAS.n885 GND 0.006836f
C5459 CS_BIAS.n886 GND 0.006836f
C5460 CS_BIAS.n887 GND 0.012677f
C5461 CS_BIAS.n888 GND 0.012419f
C5462 CS_BIAS.n889 GND 0.004099f
C5463 CS_BIAS.n890 GND 0.006836f
C5464 CS_BIAS.n891 GND 0.006836f
C5465 CS_BIAS.n892 GND 0.006836f
C5466 CS_BIAS.n893 GND 0.012677f
C5467 CS_BIAS.n894 GND 0.012677f
C5468 CS_BIAS.n895 GND 0.012677f
C5469 CS_BIAS.n896 GND 0.006836f
C5470 CS_BIAS.n897 GND 0.006836f
C5471 CS_BIAS.n898 GND 0.006836f
C5472 CS_BIAS.n899 GND 0.009548f
C5473 CS_BIAS.n900 GND 0.082235f
C5474 CS_BIAS.n901 GND 0.009548f
C5475 CS_BIAS.n902 GND 0.012677f
C5476 CS_BIAS.n903 GND 0.006836f
C5477 CS_BIAS.n904 GND 0.006836f
C5478 CS_BIAS.n905 GND 0.006836f
C5479 CS_BIAS.n906 GND 0.012677f
C5480 CS_BIAS.n907 GND 0.012677f
C5481 CS_BIAS.n908 GND 0.010554f
C5482 CS_BIAS.n909 GND 0.006836f
C5483 CS_BIAS.n910 GND 0.006836f
C5484 CS_BIAS.n911 GND 0.006836f
C5485 CS_BIAS.n912 GND 0.012419f
C5486 CS_BIAS.n913 GND 0.012677f
C5487 CS_BIAS.n914 GND 0.012677f
C5488 CS_BIAS.n915 GND 0.006836f
C5489 CS_BIAS.n916 GND 0.006836f
C5490 CS_BIAS.n917 GND 0.006836f
C5491 CS_BIAS.n918 GND 0.012677f
C5492 CS_BIAS.n919 GND 0.008046f
C5493 CS_BIAS.n920 GND 0.082235f
C5494 CS_BIAS.n921 GND 0.01105f
C5495 CS_BIAS.n922 GND 0.006836f
C5496 CS_BIAS.n923 GND 0.006836f
C5497 CS_BIAS.n924 GND 0.006836f
C5498 CS_BIAS.n925 GND 0.012677f
C5499 CS_BIAS.n926 GND 0.012677f
C5500 CS_BIAS.n927 GND 0.012904f
C5501 CS_BIAS.n928 GND 0.006836f
C5502 CS_BIAS.n929 GND 0.006836f
C5503 CS_BIAS.n930 GND 0.006836f
C5504 CS_BIAS.n931 GND 0.005106f
C5505 CS_BIAS.n932 GND 0.013606f
C5506 CS_BIAS.n933 GND 0.012677f
C5507 CS_BIAS.n934 GND 0.006836f
C5508 CS_BIAS.n935 GND 0.006836f
C5509 CS_BIAS.n936 GND 0.006836f
C5510 CS_BIAS.n937 GND 0.012677f
C5511 CS_BIAS.n938 GND 0.012677f
C5512 CS_BIAS.n939 GND 0.006544f
C5513 CS_BIAS.n940 GND 0.014459f
C5514 CS_BIAS.n941 GND 0.072784f
C5515 CS_BIAS.n942 GND 0.051747f
C5516 CS_BIAS.t37 GND 0.191402f
C5517 CS_BIAS.n943 GND 0.108818f
C5518 CS_BIAS.n944 GND 0.006836f
C5519 CS_BIAS.n945 GND 0.012677f
C5520 CS_BIAS.n946 GND 0.006836f
C5521 CS_BIAS.n947 GND 0.008132f
C5522 CS_BIAS.n948 GND 0.006836f
C5523 CS_BIAS.n949 GND 0.012677f
C5524 CS_BIAS.n950 GND 0.006836f
C5525 CS_BIAS.t28 GND 0.191402f
C5526 CS_BIAS.n951 GND 0.012677f
C5527 CS_BIAS.n952 GND 0.006836f
C5528 CS_BIAS.n953 GND 0.004099f
C5529 CS_BIAS.n954 GND 0.006836f
C5530 CS_BIAS.n955 GND 0.012677f
C5531 CS_BIAS.n956 GND 0.006836f
C5532 CS_BIAS.t21 GND 0.191402f
C5533 CS_BIAS.n957 GND 0.012677f
C5534 CS_BIAS.n958 GND 0.006836f
C5535 CS_BIAS.n959 GND 0.010554f
C5536 CS_BIAS.n960 GND 0.006836f
C5537 CS_BIAS.n961 GND 0.012677f
C5538 CS_BIAS.n962 GND 0.006836f
C5539 CS_BIAS.t57 GND 0.191402f
C5540 CS_BIAS.n963 GND 0.108333f
C5541 CS_BIAS.t63 GND 0.307989f
C5542 CS_BIAS.n964 GND 0.20812f
C5543 CS_BIAS.n965 GND 0.074665f
C5544 CS_BIAS.n966 GND 0.008046f
C5545 CS_BIAS.n967 GND 0.012677f
C5546 CS_BIAS.n968 GND 0.012677f
C5547 CS_BIAS.n969 GND 0.006836f
C5548 CS_BIAS.n970 GND 0.006836f
C5549 CS_BIAS.n971 GND 0.006836f
C5550 CS_BIAS.n972 GND 0.012677f
C5551 CS_BIAS.n973 GND 0.012419f
C5552 CS_BIAS.n974 GND 0.004099f
C5553 CS_BIAS.n975 GND 0.006836f
C5554 CS_BIAS.n976 GND 0.006836f
C5555 CS_BIAS.n977 GND 0.006836f
C5556 CS_BIAS.n978 GND 0.012677f
C5557 CS_BIAS.n979 GND 0.012677f
C5558 CS_BIAS.n980 GND 0.012677f
C5559 CS_BIAS.n981 GND 0.006836f
C5560 CS_BIAS.n982 GND 0.006836f
C5561 CS_BIAS.n983 GND 0.006836f
C5562 CS_BIAS.n984 GND 0.009548f
C5563 CS_BIAS.n985 GND 0.082235f
C5564 CS_BIAS.n986 GND 0.009548f
C5565 CS_BIAS.n987 GND 0.012677f
C5566 CS_BIAS.n988 GND 0.006836f
C5567 CS_BIAS.n989 GND 0.006836f
C5568 CS_BIAS.n990 GND 0.006836f
C5569 CS_BIAS.n991 GND 0.012677f
C5570 CS_BIAS.n992 GND 0.012677f
C5571 CS_BIAS.n993 GND 0.010554f
C5572 CS_BIAS.n994 GND 0.006836f
C5573 CS_BIAS.n995 GND 0.006836f
C5574 CS_BIAS.n996 GND 0.006836f
C5575 CS_BIAS.n997 GND 0.012419f
C5576 CS_BIAS.n998 GND 0.012677f
C5577 CS_BIAS.n999 GND 0.012677f
C5578 CS_BIAS.n1000 GND 0.006836f
C5579 CS_BIAS.n1001 GND 0.006836f
C5580 CS_BIAS.n1002 GND 0.006836f
C5581 CS_BIAS.n1003 GND 0.012677f
C5582 CS_BIAS.n1004 GND 0.008046f
C5583 CS_BIAS.n1005 GND 0.082235f
C5584 CS_BIAS.n1006 GND 0.01105f
C5585 CS_BIAS.n1007 GND 0.006836f
C5586 CS_BIAS.n1008 GND 0.006836f
C5587 CS_BIAS.n1009 GND 0.006836f
C5588 CS_BIAS.n1010 GND 0.012677f
C5589 CS_BIAS.n1011 GND 0.012677f
C5590 CS_BIAS.n1012 GND 0.012904f
C5591 CS_BIAS.n1013 GND 0.006836f
C5592 CS_BIAS.n1014 GND 0.006836f
C5593 CS_BIAS.n1015 GND 0.006836f
C5594 CS_BIAS.n1016 GND 0.005106f
C5595 CS_BIAS.n1017 GND 0.013606f
C5596 CS_BIAS.n1018 GND 0.012677f
C5597 CS_BIAS.n1019 GND 0.006836f
C5598 CS_BIAS.n1020 GND 0.006836f
C5599 CS_BIAS.n1021 GND 0.006836f
C5600 CS_BIAS.n1022 GND 0.012677f
C5601 CS_BIAS.n1023 GND 0.012677f
C5602 CS_BIAS.n1024 GND 0.006544f
C5603 CS_BIAS.n1025 GND 0.014459f
C5604 CS_BIAS.n1026 GND 0.072784f
C5605 CS_BIAS.n1027 GND 0.107952f
C5606 CS_BIAS.n1028 GND 5.6322f
.ends

