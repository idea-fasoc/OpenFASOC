* NGSPICE file created from diff_pair_sample_1401.ext - technology: sky130A

.subckt diff_pair_sample_1401 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=1.17
X1 B.t8 B.t6 B.t7 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=1.17
X2 B.t5 B.t3 B.t4 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=1.17
X3 VDD2.t1 VN.t0 VTAIL.t2 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.6591 ps=4.16 w=1.69 l=1.17
X4 B.t2 B.t0 B.t1 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0 ps=0 w=1.69 l=1.17
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.6591 ps=4.16 w=1.69 l=1.17
X6 VDD1.t1 VP.t0 VTAIL.t1 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.6591 ps=4.16 w=1.69 l=1.17
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1570_n1306# sky130_fd_pr__pfet_01v8 ad=0.6591 pd=4.16 as=0.6591 ps=4.16 w=1.69 l=1.17
R0 B.n204 B.n203 585
R1 B.n205 B.n30 585
R2 B.n207 B.n206 585
R3 B.n208 B.n29 585
R4 B.n210 B.n209 585
R5 B.n211 B.n28 585
R6 B.n213 B.n212 585
R7 B.n214 B.n27 585
R8 B.n216 B.n215 585
R9 B.n217 B.n26 585
R10 B.n219 B.n218 585
R11 B.n221 B.n23 585
R12 B.n223 B.n222 585
R13 B.n224 B.n22 585
R14 B.n226 B.n225 585
R15 B.n227 B.n21 585
R16 B.n229 B.n228 585
R17 B.n230 B.n20 585
R18 B.n232 B.n231 585
R19 B.n233 B.n19 585
R20 B.n235 B.n234 585
R21 B.n237 B.n236 585
R22 B.n238 B.n15 585
R23 B.n240 B.n239 585
R24 B.n241 B.n14 585
R25 B.n243 B.n242 585
R26 B.n244 B.n13 585
R27 B.n246 B.n245 585
R28 B.n247 B.n12 585
R29 B.n249 B.n248 585
R30 B.n250 B.n11 585
R31 B.n252 B.n251 585
R32 B.n202 B.n31 585
R33 B.n201 B.n200 585
R34 B.n199 B.n32 585
R35 B.n198 B.n197 585
R36 B.n196 B.n33 585
R37 B.n195 B.n194 585
R38 B.n193 B.n34 585
R39 B.n192 B.n191 585
R40 B.n190 B.n35 585
R41 B.n189 B.n188 585
R42 B.n187 B.n36 585
R43 B.n186 B.n185 585
R44 B.n184 B.n37 585
R45 B.n183 B.n182 585
R46 B.n181 B.n38 585
R47 B.n180 B.n179 585
R48 B.n178 B.n39 585
R49 B.n177 B.n176 585
R50 B.n175 B.n40 585
R51 B.n174 B.n173 585
R52 B.n172 B.n41 585
R53 B.n171 B.n170 585
R54 B.n169 B.n42 585
R55 B.n168 B.n167 585
R56 B.n166 B.n43 585
R57 B.n165 B.n164 585
R58 B.n163 B.n44 585
R59 B.n162 B.n161 585
R60 B.n160 B.n45 585
R61 B.n159 B.n158 585
R62 B.n157 B.n46 585
R63 B.n156 B.n155 585
R64 B.n154 B.n47 585
R65 B.n153 B.n152 585
R66 B.n151 B.n48 585
R67 B.n102 B.n101 585
R68 B.n103 B.n68 585
R69 B.n105 B.n104 585
R70 B.n106 B.n67 585
R71 B.n108 B.n107 585
R72 B.n109 B.n66 585
R73 B.n111 B.n110 585
R74 B.n112 B.n65 585
R75 B.n114 B.n113 585
R76 B.n115 B.n64 585
R77 B.n117 B.n116 585
R78 B.n119 B.n61 585
R79 B.n121 B.n120 585
R80 B.n122 B.n60 585
R81 B.n124 B.n123 585
R82 B.n125 B.n59 585
R83 B.n127 B.n126 585
R84 B.n128 B.n58 585
R85 B.n130 B.n129 585
R86 B.n131 B.n57 585
R87 B.n133 B.n132 585
R88 B.n135 B.n134 585
R89 B.n136 B.n53 585
R90 B.n138 B.n137 585
R91 B.n139 B.n52 585
R92 B.n141 B.n140 585
R93 B.n142 B.n51 585
R94 B.n144 B.n143 585
R95 B.n145 B.n50 585
R96 B.n147 B.n146 585
R97 B.n148 B.n49 585
R98 B.n150 B.n149 585
R99 B.n100 B.n69 585
R100 B.n99 B.n98 585
R101 B.n97 B.n70 585
R102 B.n96 B.n95 585
R103 B.n94 B.n71 585
R104 B.n93 B.n92 585
R105 B.n91 B.n72 585
R106 B.n90 B.n89 585
R107 B.n88 B.n73 585
R108 B.n87 B.n86 585
R109 B.n85 B.n74 585
R110 B.n84 B.n83 585
R111 B.n82 B.n75 585
R112 B.n81 B.n80 585
R113 B.n79 B.n76 585
R114 B.n78 B.n77 585
R115 B.n2 B.n0 585
R116 B.n277 B.n1 585
R117 B.n276 B.n275 585
R118 B.n274 B.n3 585
R119 B.n273 B.n272 585
R120 B.n271 B.n4 585
R121 B.n270 B.n269 585
R122 B.n268 B.n5 585
R123 B.n267 B.n266 585
R124 B.n265 B.n6 585
R125 B.n264 B.n263 585
R126 B.n262 B.n7 585
R127 B.n261 B.n260 585
R128 B.n259 B.n8 585
R129 B.n258 B.n257 585
R130 B.n256 B.n9 585
R131 B.n255 B.n254 585
R132 B.n253 B.n10 585
R133 B.n279 B.n278 585
R134 B.n102 B.n69 502.111
R135 B.n253 B.n252 502.111
R136 B.n151 B.n150 502.111
R137 B.n204 B.n31 502.111
R138 B.n54 B.t2 279.788
R139 B.n24 B.t4 279.788
R140 B.n62 B.t11 279.786
R141 B.n16 B.t7 279.786
R142 B.n55 B.t1 250.696
R143 B.n25 B.t5 250.696
R144 B.n63 B.t10 250.696
R145 B.n17 B.t8 250.696
R146 B.n54 B.t0 238.768
R147 B.n62 B.t9 238.768
R148 B.n16 B.t6 238.768
R149 B.n24 B.t3 238.768
R150 B.n98 B.n69 163.367
R151 B.n98 B.n97 163.367
R152 B.n97 B.n96 163.367
R153 B.n96 B.n71 163.367
R154 B.n92 B.n71 163.367
R155 B.n92 B.n91 163.367
R156 B.n91 B.n90 163.367
R157 B.n90 B.n73 163.367
R158 B.n86 B.n73 163.367
R159 B.n86 B.n85 163.367
R160 B.n85 B.n84 163.367
R161 B.n84 B.n75 163.367
R162 B.n80 B.n75 163.367
R163 B.n80 B.n79 163.367
R164 B.n79 B.n78 163.367
R165 B.n78 B.n2 163.367
R166 B.n278 B.n2 163.367
R167 B.n278 B.n277 163.367
R168 B.n277 B.n276 163.367
R169 B.n276 B.n3 163.367
R170 B.n272 B.n3 163.367
R171 B.n272 B.n271 163.367
R172 B.n271 B.n270 163.367
R173 B.n270 B.n5 163.367
R174 B.n266 B.n5 163.367
R175 B.n266 B.n265 163.367
R176 B.n265 B.n264 163.367
R177 B.n264 B.n7 163.367
R178 B.n260 B.n7 163.367
R179 B.n260 B.n259 163.367
R180 B.n259 B.n258 163.367
R181 B.n258 B.n9 163.367
R182 B.n254 B.n9 163.367
R183 B.n254 B.n253 163.367
R184 B.n103 B.n102 163.367
R185 B.n104 B.n103 163.367
R186 B.n104 B.n67 163.367
R187 B.n108 B.n67 163.367
R188 B.n109 B.n108 163.367
R189 B.n110 B.n109 163.367
R190 B.n110 B.n65 163.367
R191 B.n114 B.n65 163.367
R192 B.n115 B.n114 163.367
R193 B.n116 B.n115 163.367
R194 B.n116 B.n61 163.367
R195 B.n121 B.n61 163.367
R196 B.n122 B.n121 163.367
R197 B.n123 B.n122 163.367
R198 B.n123 B.n59 163.367
R199 B.n127 B.n59 163.367
R200 B.n128 B.n127 163.367
R201 B.n129 B.n128 163.367
R202 B.n129 B.n57 163.367
R203 B.n133 B.n57 163.367
R204 B.n134 B.n133 163.367
R205 B.n134 B.n53 163.367
R206 B.n138 B.n53 163.367
R207 B.n139 B.n138 163.367
R208 B.n140 B.n139 163.367
R209 B.n140 B.n51 163.367
R210 B.n144 B.n51 163.367
R211 B.n145 B.n144 163.367
R212 B.n146 B.n145 163.367
R213 B.n146 B.n49 163.367
R214 B.n150 B.n49 163.367
R215 B.n152 B.n151 163.367
R216 B.n152 B.n47 163.367
R217 B.n156 B.n47 163.367
R218 B.n157 B.n156 163.367
R219 B.n158 B.n157 163.367
R220 B.n158 B.n45 163.367
R221 B.n162 B.n45 163.367
R222 B.n163 B.n162 163.367
R223 B.n164 B.n163 163.367
R224 B.n164 B.n43 163.367
R225 B.n168 B.n43 163.367
R226 B.n169 B.n168 163.367
R227 B.n170 B.n169 163.367
R228 B.n170 B.n41 163.367
R229 B.n174 B.n41 163.367
R230 B.n175 B.n174 163.367
R231 B.n176 B.n175 163.367
R232 B.n176 B.n39 163.367
R233 B.n180 B.n39 163.367
R234 B.n181 B.n180 163.367
R235 B.n182 B.n181 163.367
R236 B.n182 B.n37 163.367
R237 B.n186 B.n37 163.367
R238 B.n187 B.n186 163.367
R239 B.n188 B.n187 163.367
R240 B.n188 B.n35 163.367
R241 B.n192 B.n35 163.367
R242 B.n193 B.n192 163.367
R243 B.n194 B.n193 163.367
R244 B.n194 B.n33 163.367
R245 B.n198 B.n33 163.367
R246 B.n199 B.n198 163.367
R247 B.n200 B.n199 163.367
R248 B.n200 B.n31 163.367
R249 B.n252 B.n11 163.367
R250 B.n248 B.n11 163.367
R251 B.n248 B.n247 163.367
R252 B.n247 B.n246 163.367
R253 B.n246 B.n13 163.367
R254 B.n242 B.n13 163.367
R255 B.n242 B.n241 163.367
R256 B.n241 B.n240 163.367
R257 B.n240 B.n15 163.367
R258 B.n236 B.n15 163.367
R259 B.n236 B.n235 163.367
R260 B.n235 B.n19 163.367
R261 B.n231 B.n19 163.367
R262 B.n231 B.n230 163.367
R263 B.n230 B.n229 163.367
R264 B.n229 B.n21 163.367
R265 B.n225 B.n21 163.367
R266 B.n225 B.n224 163.367
R267 B.n224 B.n223 163.367
R268 B.n223 B.n23 163.367
R269 B.n218 B.n23 163.367
R270 B.n218 B.n217 163.367
R271 B.n217 B.n216 163.367
R272 B.n216 B.n27 163.367
R273 B.n212 B.n27 163.367
R274 B.n212 B.n211 163.367
R275 B.n211 B.n210 163.367
R276 B.n210 B.n29 163.367
R277 B.n206 B.n29 163.367
R278 B.n206 B.n205 163.367
R279 B.n205 B.n204 163.367
R280 B.n56 B.n55 59.5399
R281 B.n118 B.n63 59.5399
R282 B.n18 B.n17 59.5399
R283 B.n220 B.n25 59.5399
R284 B.n251 B.n10 32.6249
R285 B.n203 B.n202 32.6249
R286 B.n149 B.n48 32.6249
R287 B.n101 B.n100 32.6249
R288 B.n55 B.n54 29.0914
R289 B.n63 B.n62 29.0914
R290 B.n17 B.n16 29.0914
R291 B.n25 B.n24 29.0914
R292 B B.n279 18.0485
R293 B.n251 B.n250 10.6151
R294 B.n250 B.n249 10.6151
R295 B.n249 B.n12 10.6151
R296 B.n245 B.n12 10.6151
R297 B.n245 B.n244 10.6151
R298 B.n244 B.n243 10.6151
R299 B.n243 B.n14 10.6151
R300 B.n239 B.n14 10.6151
R301 B.n239 B.n238 10.6151
R302 B.n238 B.n237 10.6151
R303 B.n234 B.n233 10.6151
R304 B.n233 B.n232 10.6151
R305 B.n232 B.n20 10.6151
R306 B.n228 B.n20 10.6151
R307 B.n228 B.n227 10.6151
R308 B.n227 B.n226 10.6151
R309 B.n226 B.n22 10.6151
R310 B.n222 B.n22 10.6151
R311 B.n222 B.n221 10.6151
R312 B.n219 B.n26 10.6151
R313 B.n215 B.n26 10.6151
R314 B.n215 B.n214 10.6151
R315 B.n214 B.n213 10.6151
R316 B.n213 B.n28 10.6151
R317 B.n209 B.n28 10.6151
R318 B.n209 B.n208 10.6151
R319 B.n208 B.n207 10.6151
R320 B.n207 B.n30 10.6151
R321 B.n203 B.n30 10.6151
R322 B.n153 B.n48 10.6151
R323 B.n154 B.n153 10.6151
R324 B.n155 B.n154 10.6151
R325 B.n155 B.n46 10.6151
R326 B.n159 B.n46 10.6151
R327 B.n160 B.n159 10.6151
R328 B.n161 B.n160 10.6151
R329 B.n161 B.n44 10.6151
R330 B.n165 B.n44 10.6151
R331 B.n166 B.n165 10.6151
R332 B.n167 B.n166 10.6151
R333 B.n167 B.n42 10.6151
R334 B.n171 B.n42 10.6151
R335 B.n172 B.n171 10.6151
R336 B.n173 B.n172 10.6151
R337 B.n173 B.n40 10.6151
R338 B.n177 B.n40 10.6151
R339 B.n178 B.n177 10.6151
R340 B.n179 B.n178 10.6151
R341 B.n179 B.n38 10.6151
R342 B.n183 B.n38 10.6151
R343 B.n184 B.n183 10.6151
R344 B.n185 B.n184 10.6151
R345 B.n185 B.n36 10.6151
R346 B.n189 B.n36 10.6151
R347 B.n190 B.n189 10.6151
R348 B.n191 B.n190 10.6151
R349 B.n191 B.n34 10.6151
R350 B.n195 B.n34 10.6151
R351 B.n196 B.n195 10.6151
R352 B.n197 B.n196 10.6151
R353 B.n197 B.n32 10.6151
R354 B.n201 B.n32 10.6151
R355 B.n202 B.n201 10.6151
R356 B.n101 B.n68 10.6151
R357 B.n105 B.n68 10.6151
R358 B.n106 B.n105 10.6151
R359 B.n107 B.n106 10.6151
R360 B.n107 B.n66 10.6151
R361 B.n111 B.n66 10.6151
R362 B.n112 B.n111 10.6151
R363 B.n113 B.n112 10.6151
R364 B.n113 B.n64 10.6151
R365 B.n117 B.n64 10.6151
R366 B.n120 B.n119 10.6151
R367 B.n120 B.n60 10.6151
R368 B.n124 B.n60 10.6151
R369 B.n125 B.n124 10.6151
R370 B.n126 B.n125 10.6151
R371 B.n126 B.n58 10.6151
R372 B.n130 B.n58 10.6151
R373 B.n131 B.n130 10.6151
R374 B.n132 B.n131 10.6151
R375 B.n136 B.n135 10.6151
R376 B.n137 B.n136 10.6151
R377 B.n137 B.n52 10.6151
R378 B.n141 B.n52 10.6151
R379 B.n142 B.n141 10.6151
R380 B.n143 B.n142 10.6151
R381 B.n143 B.n50 10.6151
R382 B.n147 B.n50 10.6151
R383 B.n148 B.n147 10.6151
R384 B.n149 B.n148 10.6151
R385 B.n100 B.n99 10.6151
R386 B.n99 B.n70 10.6151
R387 B.n95 B.n70 10.6151
R388 B.n95 B.n94 10.6151
R389 B.n94 B.n93 10.6151
R390 B.n93 B.n72 10.6151
R391 B.n89 B.n72 10.6151
R392 B.n89 B.n88 10.6151
R393 B.n88 B.n87 10.6151
R394 B.n87 B.n74 10.6151
R395 B.n83 B.n74 10.6151
R396 B.n83 B.n82 10.6151
R397 B.n82 B.n81 10.6151
R398 B.n81 B.n76 10.6151
R399 B.n77 B.n76 10.6151
R400 B.n77 B.n0 10.6151
R401 B.n275 B.n1 10.6151
R402 B.n275 B.n274 10.6151
R403 B.n274 B.n273 10.6151
R404 B.n273 B.n4 10.6151
R405 B.n269 B.n4 10.6151
R406 B.n269 B.n268 10.6151
R407 B.n268 B.n267 10.6151
R408 B.n267 B.n6 10.6151
R409 B.n263 B.n6 10.6151
R410 B.n263 B.n262 10.6151
R411 B.n262 B.n261 10.6151
R412 B.n261 B.n8 10.6151
R413 B.n257 B.n8 10.6151
R414 B.n257 B.n256 10.6151
R415 B.n256 B.n255 10.6151
R416 B.n255 B.n10 10.6151
R417 B.n237 B.n18 9.36635
R418 B.n220 B.n219 9.36635
R419 B.n118 B.n117 9.36635
R420 B.n135 B.n56 9.36635
R421 B.n279 B.n0 2.81026
R422 B.n279 B.n1 2.81026
R423 B.n234 B.n18 1.24928
R424 B.n221 B.n220 1.24928
R425 B.n119 B.n118 1.24928
R426 B.n132 B.n56 1.24928
R427 VN VN.t0 182.536
R428 VN VN.t1 149.343
R429 VTAIL.n3 VTAIL.t3 252.861
R430 VTAIL.n0 VTAIL.t0 252.861
R431 VTAIL.n2 VTAIL.t1 252.861
R432 VTAIL.n1 VTAIL.t2 252.861
R433 VTAIL.n1 VTAIL.n0 16.41
R434 VTAIL.n3 VTAIL.n2 15.1169
R435 VTAIL.n2 VTAIL.n1 1.11688
R436 VTAIL VTAIL.n0 0.851793
R437 VTAIL VTAIL.n3 0.265586
R438 VDD2.n0 VDD2.t0 297.241
R439 VDD2.n0 VDD2.t1 269.539
R440 VDD2 VDD2.n0 0.381966
R441 VP.n0 VP.t0 182.25
R442 VP.n0 VP.t1 149.196
R443 VP VP.n0 0.146778
R444 VDD1 VDD1.t0 298.089
R445 VDD1 VDD1.t1 269.921
C0 w_n1570_n1306# VTAIL 1.16717f
C1 w_n1570_n1306# B 4.36515f
C2 VDD1 VDD2 0.507835f
C3 VDD1 VTAIL 1.92282f
C4 VDD1 B 0.720759f
C5 VTAIL VDD2 1.96583f
C6 VDD2 B 0.738908f
C7 VTAIL B 0.917338f
C8 VP VN 2.88582f
C9 VN w_n1570_n1306# 1.81661f
C10 VN VDD1 0.154229f
C11 VN VDD2 0.540058f
C12 VN VTAIL 0.663067f
C13 VN B 0.661279f
C14 VP w_n1570_n1306# 2.00787f
C15 VP VDD1 0.663716f
C16 VP VDD2 0.279447f
C17 VP VTAIL 0.677227f
C18 VP B 0.978383f
C19 w_n1570_n1306# VDD1 0.869763f
C20 w_n1570_n1306# VDD2 0.878301f
C21 VDD2 VSUBS 0.36452f
C22 VDD1 VSUBS 0.537847f
C23 VTAIL VSUBS 0.218403f
C24 VN VSUBS 3.42755f
C25 VP VSUBS 0.789672f
C26 B VSUBS 1.870052f
C27 w_n1570_n1306# VSUBS 26.244099f
C28 VP.t0 VSUBS 0.886231f
C29 VP.t1 VSUBS 0.54743f
C30 VP.n0 VSUBS 3.41339f
C31 VN.t1 VSUBS 0.318317f
C32 VN.t0 VSUBS 0.520474f
C33 B.n0 VSUBS 0.006103f
C34 B.n1 VSUBS 0.006103f
C35 B.n2 VSUBS 0.009651f
C36 B.n3 VSUBS 0.009651f
C37 B.n4 VSUBS 0.009651f
C38 B.n5 VSUBS 0.009651f
C39 B.n6 VSUBS 0.009651f
C40 B.n7 VSUBS 0.009651f
C41 B.n8 VSUBS 0.009651f
C42 B.n9 VSUBS 0.009651f
C43 B.n10 VSUBS 0.022162f
C44 B.n11 VSUBS 0.009651f
C45 B.n12 VSUBS 0.009651f
C46 B.n13 VSUBS 0.009651f
C47 B.n14 VSUBS 0.009651f
C48 B.n15 VSUBS 0.009651f
C49 B.t8 VSUBS 0.048099f
C50 B.t7 VSUBS 0.053733f
C51 B.t6 VSUBS 0.133507f
C52 B.n16 VSUBS 0.076605f
C53 B.n17 VSUBS 0.067951f
C54 B.n18 VSUBS 0.022359f
C55 B.n19 VSUBS 0.009651f
C56 B.n20 VSUBS 0.009651f
C57 B.n21 VSUBS 0.009651f
C58 B.n22 VSUBS 0.009651f
C59 B.n23 VSUBS 0.009651f
C60 B.t5 VSUBS 0.048099f
C61 B.t4 VSUBS 0.053733f
C62 B.t3 VSUBS 0.133507f
C63 B.n24 VSUBS 0.076605f
C64 B.n25 VSUBS 0.067951f
C65 B.n26 VSUBS 0.009651f
C66 B.n27 VSUBS 0.009651f
C67 B.n28 VSUBS 0.009651f
C68 B.n29 VSUBS 0.009651f
C69 B.n30 VSUBS 0.009651f
C70 B.n31 VSUBS 0.022162f
C71 B.n32 VSUBS 0.009651f
C72 B.n33 VSUBS 0.009651f
C73 B.n34 VSUBS 0.009651f
C74 B.n35 VSUBS 0.009651f
C75 B.n36 VSUBS 0.009651f
C76 B.n37 VSUBS 0.009651f
C77 B.n38 VSUBS 0.009651f
C78 B.n39 VSUBS 0.009651f
C79 B.n40 VSUBS 0.009651f
C80 B.n41 VSUBS 0.009651f
C81 B.n42 VSUBS 0.009651f
C82 B.n43 VSUBS 0.009651f
C83 B.n44 VSUBS 0.009651f
C84 B.n45 VSUBS 0.009651f
C85 B.n46 VSUBS 0.009651f
C86 B.n47 VSUBS 0.009651f
C87 B.n48 VSUBS 0.022162f
C88 B.n49 VSUBS 0.009651f
C89 B.n50 VSUBS 0.009651f
C90 B.n51 VSUBS 0.009651f
C91 B.n52 VSUBS 0.009651f
C92 B.n53 VSUBS 0.009651f
C93 B.t1 VSUBS 0.048099f
C94 B.t2 VSUBS 0.053733f
C95 B.t0 VSUBS 0.133507f
C96 B.n54 VSUBS 0.076605f
C97 B.n55 VSUBS 0.067951f
C98 B.n56 VSUBS 0.022359f
C99 B.n57 VSUBS 0.009651f
C100 B.n58 VSUBS 0.009651f
C101 B.n59 VSUBS 0.009651f
C102 B.n60 VSUBS 0.009651f
C103 B.n61 VSUBS 0.009651f
C104 B.t10 VSUBS 0.048099f
C105 B.t11 VSUBS 0.053733f
C106 B.t9 VSUBS 0.133507f
C107 B.n62 VSUBS 0.076605f
C108 B.n63 VSUBS 0.067951f
C109 B.n64 VSUBS 0.009651f
C110 B.n65 VSUBS 0.009651f
C111 B.n66 VSUBS 0.009651f
C112 B.n67 VSUBS 0.009651f
C113 B.n68 VSUBS 0.009651f
C114 B.n69 VSUBS 0.022162f
C115 B.n70 VSUBS 0.009651f
C116 B.n71 VSUBS 0.009651f
C117 B.n72 VSUBS 0.009651f
C118 B.n73 VSUBS 0.009651f
C119 B.n74 VSUBS 0.009651f
C120 B.n75 VSUBS 0.009651f
C121 B.n76 VSUBS 0.009651f
C122 B.n77 VSUBS 0.009651f
C123 B.n78 VSUBS 0.009651f
C124 B.n79 VSUBS 0.009651f
C125 B.n80 VSUBS 0.009651f
C126 B.n81 VSUBS 0.009651f
C127 B.n82 VSUBS 0.009651f
C128 B.n83 VSUBS 0.009651f
C129 B.n84 VSUBS 0.009651f
C130 B.n85 VSUBS 0.009651f
C131 B.n86 VSUBS 0.009651f
C132 B.n87 VSUBS 0.009651f
C133 B.n88 VSUBS 0.009651f
C134 B.n89 VSUBS 0.009651f
C135 B.n90 VSUBS 0.009651f
C136 B.n91 VSUBS 0.009651f
C137 B.n92 VSUBS 0.009651f
C138 B.n93 VSUBS 0.009651f
C139 B.n94 VSUBS 0.009651f
C140 B.n95 VSUBS 0.009651f
C141 B.n96 VSUBS 0.009651f
C142 B.n97 VSUBS 0.009651f
C143 B.n98 VSUBS 0.009651f
C144 B.n99 VSUBS 0.009651f
C145 B.n100 VSUBS 0.022162f
C146 B.n101 VSUBS 0.022969f
C147 B.n102 VSUBS 0.022969f
C148 B.n103 VSUBS 0.009651f
C149 B.n104 VSUBS 0.009651f
C150 B.n105 VSUBS 0.009651f
C151 B.n106 VSUBS 0.009651f
C152 B.n107 VSUBS 0.009651f
C153 B.n108 VSUBS 0.009651f
C154 B.n109 VSUBS 0.009651f
C155 B.n110 VSUBS 0.009651f
C156 B.n111 VSUBS 0.009651f
C157 B.n112 VSUBS 0.009651f
C158 B.n113 VSUBS 0.009651f
C159 B.n114 VSUBS 0.009651f
C160 B.n115 VSUBS 0.009651f
C161 B.n116 VSUBS 0.009651f
C162 B.n117 VSUBS 0.009083f
C163 B.n118 VSUBS 0.022359f
C164 B.n119 VSUBS 0.005393f
C165 B.n120 VSUBS 0.009651f
C166 B.n121 VSUBS 0.009651f
C167 B.n122 VSUBS 0.009651f
C168 B.n123 VSUBS 0.009651f
C169 B.n124 VSUBS 0.009651f
C170 B.n125 VSUBS 0.009651f
C171 B.n126 VSUBS 0.009651f
C172 B.n127 VSUBS 0.009651f
C173 B.n128 VSUBS 0.009651f
C174 B.n129 VSUBS 0.009651f
C175 B.n130 VSUBS 0.009651f
C176 B.n131 VSUBS 0.009651f
C177 B.n132 VSUBS 0.005393f
C178 B.n133 VSUBS 0.009651f
C179 B.n134 VSUBS 0.009651f
C180 B.n135 VSUBS 0.009083f
C181 B.n136 VSUBS 0.009651f
C182 B.n137 VSUBS 0.009651f
C183 B.n138 VSUBS 0.009651f
C184 B.n139 VSUBS 0.009651f
C185 B.n140 VSUBS 0.009651f
C186 B.n141 VSUBS 0.009651f
C187 B.n142 VSUBS 0.009651f
C188 B.n143 VSUBS 0.009651f
C189 B.n144 VSUBS 0.009651f
C190 B.n145 VSUBS 0.009651f
C191 B.n146 VSUBS 0.009651f
C192 B.n147 VSUBS 0.009651f
C193 B.n148 VSUBS 0.009651f
C194 B.n149 VSUBS 0.022969f
C195 B.n150 VSUBS 0.022969f
C196 B.n151 VSUBS 0.022162f
C197 B.n152 VSUBS 0.009651f
C198 B.n153 VSUBS 0.009651f
C199 B.n154 VSUBS 0.009651f
C200 B.n155 VSUBS 0.009651f
C201 B.n156 VSUBS 0.009651f
C202 B.n157 VSUBS 0.009651f
C203 B.n158 VSUBS 0.009651f
C204 B.n159 VSUBS 0.009651f
C205 B.n160 VSUBS 0.009651f
C206 B.n161 VSUBS 0.009651f
C207 B.n162 VSUBS 0.009651f
C208 B.n163 VSUBS 0.009651f
C209 B.n164 VSUBS 0.009651f
C210 B.n165 VSUBS 0.009651f
C211 B.n166 VSUBS 0.009651f
C212 B.n167 VSUBS 0.009651f
C213 B.n168 VSUBS 0.009651f
C214 B.n169 VSUBS 0.009651f
C215 B.n170 VSUBS 0.009651f
C216 B.n171 VSUBS 0.009651f
C217 B.n172 VSUBS 0.009651f
C218 B.n173 VSUBS 0.009651f
C219 B.n174 VSUBS 0.009651f
C220 B.n175 VSUBS 0.009651f
C221 B.n176 VSUBS 0.009651f
C222 B.n177 VSUBS 0.009651f
C223 B.n178 VSUBS 0.009651f
C224 B.n179 VSUBS 0.009651f
C225 B.n180 VSUBS 0.009651f
C226 B.n181 VSUBS 0.009651f
C227 B.n182 VSUBS 0.009651f
C228 B.n183 VSUBS 0.009651f
C229 B.n184 VSUBS 0.009651f
C230 B.n185 VSUBS 0.009651f
C231 B.n186 VSUBS 0.009651f
C232 B.n187 VSUBS 0.009651f
C233 B.n188 VSUBS 0.009651f
C234 B.n189 VSUBS 0.009651f
C235 B.n190 VSUBS 0.009651f
C236 B.n191 VSUBS 0.009651f
C237 B.n192 VSUBS 0.009651f
C238 B.n193 VSUBS 0.009651f
C239 B.n194 VSUBS 0.009651f
C240 B.n195 VSUBS 0.009651f
C241 B.n196 VSUBS 0.009651f
C242 B.n197 VSUBS 0.009651f
C243 B.n198 VSUBS 0.009651f
C244 B.n199 VSUBS 0.009651f
C245 B.n200 VSUBS 0.009651f
C246 B.n201 VSUBS 0.009651f
C247 B.n202 VSUBS 0.023303f
C248 B.n203 VSUBS 0.021827f
C249 B.n204 VSUBS 0.022969f
C250 B.n205 VSUBS 0.009651f
C251 B.n206 VSUBS 0.009651f
C252 B.n207 VSUBS 0.009651f
C253 B.n208 VSUBS 0.009651f
C254 B.n209 VSUBS 0.009651f
C255 B.n210 VSUBS 0.009651f
C256 B.n211 VSUBS 0.009651f
C257 B.n212 VSUBS 0.009651f
C258 B.n213 VSUBS 0.009651f
C259 B.n214 VSUBS 0.009651f
C260 B.n215 VSUBS 0.009651f
C261 B.n216 VSUBS 0.009651f
C262 B.n217 VSUBS 0.009651f
C263 B.n218 VSUBS 0.009651f
C264 B.n219 VSUBS 0.009083f
C265 B.n220 VSUBS 0.022359f
C266 B.n221 VSUBS 0.005393f
C267 B.n222 VSUBS 0.009651f
C268 B.n223 VSUBS 0.009651f
C269 B.n224 VSUBS 0.009651f
C270 B.n225 VSUBS 0.009651f
C271 B.n226 VSUBS 0.009651f
C272 B.n227 VSUBS 0.009651f
C273 B.n228 VSUBS 0.009651f
C274 B.n229 VSUBS 0.009651f
C275 B.n230 VSUBS 0.009651f
C276 B.n231 VSUBS 0.009651f
C277 B.n232 VSUBS 0.009651f
C278 B.n233 VSUBS 0.009651f
C279 B.n234 VSUBS 0.005393f
C280 B.n235 VSUBS 0.009651f
C281 B.n236 VSUBS 0.009651f
C282 B.n237 VSUBS 0.009083f
C283 B.n238 VSUBS 0.009651f
C284 B.n239 VSUBS 0.009651f
C285 B.n240 VSUBS 0.009651f
C286 B.n241 VSUBS 0.009651f
C287 B.n242 VSUBS 0.009651f
C288 B.n243 VSUBS 0.009651f
C289 B.n244 VSUBS 0.009651f
C290 B.n245 VSUBS 0.009651f
C291 B.n246 VSUBS 0.009651f
C292 B.n247 VSUBS 0.009651f
C293 B.n248 VSUBS 0.009651f
C294 B.n249 VSUBS 0.009651f
C295 B.n250 VSUBS 0.009651f
C296 B.n251 VSUBS 0.022969f
C297 B.n252 VSUBS 0.022969f
C298 B.n253 VSUBS 0.022162f
C299 B.n254 VSUBS 0.009651f
C300 B.n255 VSUBS 0.009651f
C301 B.n256 VSUBS 0.009651f
C302 B.n257 VSUBS 0.009651f
C303 B.n258 VSUBS 0.009651f
C304 B.n259 VSUBS 0.009651f
C305 B.n260 VSUBS 0.009651f
C306 B.n261 VSUBS 0.009651f
C307 B.n262 VSUBS 0.009651f
C308 B.n263 VSUBS 0.009651f
C309 B.n264 VSUBS 0.009651f
C310 B.n265 VSUBS 0.009651f
C311 B.n266 VSUBS 0.009651f
C312 B.n267 VSUBS 0.009651f
C313 B.n268 VSUBS 0.009651f
C314 B.n269 VSUBS 0.009651f
C315 B.n270 VSUBS 0.009651f
C316 B.n271 VSUBS 0.009651f
C317 B.n272 VSUBS 0.009651f
C318 B.n273 VSUBS 0.009651f
C319 B.n274 VSUBS 0.009651f
C320 B.n275 VSUBS 0.009651f
C321 B.n276 VSUBS 0.009651f
C322 B.n277 VSUBS 0.009651f
C323 B.n278 VSUBS 0.009651f
C324 B.n279 VSUBS 0.021852f
.ends

