* NGSPICE file created from diff_pair_sample_1315.ext - technology: sky130A

.subckt diff_pair_sample_1315 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t1 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=1.93215 ps=12.04 w=11.71 l=2.83
X1 B.t11 B.t9 B.t10 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=0 ps=0 w=11.71 l=2.83
X2 VDD2.t3 VN.t1 VTAIL.t5 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=1.93215 pd=12.04 as=4.5669 ps=24.2 w=11.71 l=2.83
X3 VDD1.t3 VP.t0 VTAIL.t1 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=1.93215 pd=12.04 as=4.5669 ps=24.2 w=11.71 l=2.83
X4 VTAIL.t4 VN.t2 VDD2.t2 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=1.93215 ps=12.04 w=11.71 l=2.83
X5 VDD1.t2 VP.t1 VTAIL.t7 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=1.93215 pd=12.04 as=4.5669 ps=24.2 w=11.71 l=2.83
X6 VTAIL.t2 VP.t2 VDD1.t1 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=1.93215 ps=12.04 w=11.71 l=2.83
X7 B.t8 B.t6 B.t7 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=0 ps=0 w=11.71 l=2.83
X8 VDD2.t0 VN.t3 VTAIL.t3 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=1.93215 pd=12.04 as=4.5669 ps=24.2 w=11.71 l=2.83
X9 B.t5 B.t3 B.t4 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=0 ps=0 w=11.71 l=2.83
X10 VTAIL.t0 VP.t3 VDD1.t0 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=1.93215 ps=12.04 w=11.71 l=2.83
X11 B.t2 B.t0 B.t1 w_n2866_n3310# sky130_fd_pr__pfet_01v8 ad=4.5669 pd=24.2 as=0 ps=0 w=11.71 l=2.83
R0 VN.n0 VN.t0 134.948
R1 VN.n1 VN.t3 134.948
R2 VN.n0 VN.t1 134.054
R3 VN.n1 VN.t2 134.054
R4 VN VN.n1 50.5371
R5 VN VN.n0 3.46509
R6 VDD2.n2 VDD2.n0 115.308
R7 VDD2.n2 VDD2.n1 73.325
R8 VDD2.n1 VDD2.t2 2.77633
R9 VDD2.n1 VDD2.t0 2.77633
R10 VDD2.n0 VDD2.t1 2.77633
R11 VDD2.n0 VDD2.t3 2.77633
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t0 59.4223
R14 VTAIL.n4 VTAIL.t3 59.4223
R15 VTAIL.n3 VTAIL.t4 59.4223
R16 VTAIL.n7 VTAIL.t5 59.422
R17 VTAIL.n0 VTAIL.t6 59.422
R18 VTAIL.n1 VTAIL.t1 59.422
R19 VTAIL.n2 VTAIL.t2 59.422
R20 VTAIL.n6 VTAIL.t7 59.422
R21 VTAIL.n7 VTAIL.n6 25.1858
R22 VTAIL.n3 VTAIL.n2 25.1858
R23 VTAIL.n4 VTAIL.n3 2.72464
R24 VTAIL.n6 VTAIL.n5 2.72464
R25 VTAIL.n2 VTAIL.n1 2.72464
R26 VTAIL VTAIL.n0 1.42076
R27 VTAIL VTAIL.n7 1.30438
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n475 B.n70 585
R31 B.n477 B.n476 585
R32 B.n478 B.n69 585
R33 B.n480 B.n479 585
R34 B.n481 B.n68 585
R35 B.n483 B.n482 585
R36 B.n484 B.n67 585
R37 B.n486 B.n485 585
R38 B.n487 B.n66 585
R39 B.n489 B.n488 585
R40 B.n490 B.n65 585
R41 B.n492 B.n491 585
R42 B.n493 B.n64 585
R43 B.n495 B.n494 585
R44 B.n496 B.n63 585
R45 B.n498 B.n497 585
R46 B.n499 B.n62 585
R47 B.n501 B.n500 585
R48 B.n502 B.n61 585
R49 B.n504 B.n503 585
R50 B.n505 B.n60 585
R51 B.n507 B.n506 585
R52 B.n508 B.n59 585
R53 B.n510 B.n509 585
R54 B.n511 B.n58 585
R55 B.n513 B.n512 585
R56 B.n514 B.n57 585
R57 B.n516 B.n515 585
R58 B.n517 B.n56 585
R59 B.n519 B.n518 585
R60 B.n520 B.n55 585
R61 B.n522 B.n521 585
R62 B.n523 B.n54 585
R63 B.n525 B.n524 585
R64 B.n526 B.n53 585
R65 B.n528 B.n527 585
R66 B.n529 B.n52 585
R67 B.n531 B.n530 585
R68 B.n532 B.n51 585
R69 B.n534 B.n533 585
R70 B.n535 B.n48 585
R71 B.n538 B.n537 585
R72 B.n539 B.n47 585
R73 B.n541 B.n540 585
R74 B.n542 B.n46 585
R75 B.n544 B.n543 585
R76 B.n545 B.n45 585
R77 B.n547 B.n546 585
R78 B.n548 B.n41 585
R79 B.n550 B.n549 585
R80 B.n551 B.n40 585
R81 B.n553 B.n552 585
R82 B.n554 B.n39 585
R83 B.n556 B.n555 585
R84 B.n557 B.n38 585
R85 B.n559 B.n558 585
R86 B.n560 B.n37 585
R87 B.n562 B.n561 585
R88 B.n563 B.n36 585
R89 B.n565 B.n564 585
R90 B.n566 B.n35 585
R91 B.n568 B.n567 585
R92 B.n569 B.n34 585
R93 B.n571 B.n570 585
R94 B.n572 B.n33 585
R95 B.n574 B.n573 585
R96 B.n575 B.n32 585
R97 B.n577 B.n576 585
R98 B.n578 B.n31 585
R99 B.n580 B.n579 585
R100 B.n581 B.n30 585
R101 B.n583 B.n582 585
R102 B.n584 B.n29 585
R103 B.n586 B.n585 585
R104 B.n587 B.n28 585
R105 B.n589 B.n588 585
R106 B.n590 B.n27 585
R107 B.n592 B.n591 585
R108 B.n593 B.n26 585
R109 B.n595 B.n594 585
R110 B.n596 B.n25 585
R111 B.n598 B.n597 585
R112 B.n599 B.n24 585
R113 B.n601 B.n600 585
R114 B.n602 B.n23 585
R115 B.n604 B.n603 585
R116 B.n605 B.n22 585
R117 B.n607 B.n606 585
R118 B.n608 B.n21 585
R119 B.n610 B.n609 585
R120 B.n611 B.n20 585
R121 B.n474 B.n473 585
R122 B.n472 B.n71 585
R123 B.n471 B.n470 585
R124 B.n469 B.n72 585
R125 B.n468 B.n467 585
R126 B.n466 B.n73 585
R127 B.n465 B.n464 585
R128 B.n463 B.n74 585
R129 B.n462 B.n461 585
R130 B.n460 B.n75 585
R131 B.n459 B.n458 585
R132 B.n457 B.n76 585
R133 B.n456 B.n455 585
R134 B.n454 B.n77 585
R135 B.n453 B.n452 585
R136 B.n451 B.n78 585
R137 B.n450 B.n449 585
R138 B.n448 B.n79 585
R139 B.n447 B.n446 585
R140 B.n445 B.n80 585
R141 B.n444 B.n443 585
R142 B.n442 B.n81 585
R143 B.n441 B.n440 585
R144 B.n439 B.n82 585
R145 B.n438 B.n437 585
R146 B.n436 B.n83 585
R147 B.n435 B.n434 585
R148 B.n433 B.n84 585
R149 B.n432 B.n431 585
R150 B.n430 B.n85 585
R151 B.n429 B.n428 585
R152 B.n427 B.n86 585
R153 B.n426 B.n425 585
R154 B.n424 B.n87 585
R155 B.n423 B.n422 585
R156 B.n421 B.n88 585
R157 B.n420 B.n419 585
R158 B.n418 B.n89 585
R159 B.n417 B.n416 585
R160 B.n415 B.n90 585
R161 B.n414 B.n413 585
R162 B.n412 B.n91 585
R163 B.n411 B.n410 585
R164 B.n409 B.n92 585
R165 B.n408 B.n407 585
R166 B.n406 B.n93 585
R167 B.n405 B.n404 585
R168 B.n403 B.n94 585
R169 B.n402 B.n401 585
R170 B.n400 B.n95 585
R171 B.n399 B.n398 585
R172 B.n397 B.n96 585
R173 B.n396 B.n395 585
R174 B.n394 B.n97 585
R175 B.n393 B.n392 585
R176 B.n391 B.n98 585
R177 B.n390 B.n389 585
R178 B.n388 B.n99 585
R179 B.n387 B.n386 585
R180 B.n385 B.n100 585
R181 B.n384 B.n383 585
R182 B.n382 B.n101 585
R183 B.n381 B.n380 585
R184 B.n379 B.n102 585
R185 B.n378 B.n377 585
R186 B.n376 B.n103 585
R187 B.n375 B.n374 585
R188 B.n373 B.n104 585
R189 B.n372 B.n371 585
R190 B.n370 B.n105 585
R191 B.n369 B.n368 585
R192 B.n367 B.n106 585
R193 B.n366 B.n365 585
R194 B.n225 B.n154 585
R195 B.n227 B.n226 585
R196 B.n228 B.n153 585
R197 B.n230 B.n229 585
R198 B.n231 B.n152 585
R199 B.n233 B.n232 585
R200 B.n234 B.n151 585
R201 B.n236 B.n235 585
R202 B.n237 B.n150 585
R203 B.n239 B.n238 585
R204 B.n240 B.n149 585
R205 B.n242 B.n241 585
R206 B.n243 B.n148 585
R207 B.n245 B.n244 585
R208 B.n246 B.n147 585
R209 B.n248 B.n247 585
R210 B.n249 B.n146 585
R211 B.n251 B.n250 585
R212 B.n252 B.n145 585
R213 B.n254 B.n253 585
R214 B.n255 B.n144 585
R215 B.n257 B.n256 585
R216 B.n258 B.n143 585
R217 B.n260 B.n259 585
R218 B.n261 B.n142 585
R219 B.n263 B.n262 585
R220 B.n264 B.n141 585
R221 B.n266 B.n265 585
R222 B.n267 B.n140 585
R223 B.n269 B.n268 585
R224 B.n270 B.n139 585
R225 B.n272 B.n271 585
R226 B.n273 B.n138 585
R227 B.n275 B.n274 585
R228 B.n276 B.n137 585
R229 B.n278 B.n277 585
R230 B.n279 B.n136 585
R231 B.n281 B.n280 585
R232 B.n282 B.n135 585
R233 B.n284 B.n283 585
R234 B.n285 B.n132 585
R235 B.n288 B.n287 585
R236 B.n289 B.n131 585
R237 B.n291 B.n290 585
R238 B.n292 B.n130 585
R239 B.n294 B.n293 585
R240 B.n295 B.n129 585
R241 B.n297 B.n296 585
R242 B.n298 B.n128 585
R243 B.n303 B.n302 585
R244 B.n304 B.n127 585
R245 B.n306 B.n305 585
R246 B.n307 B.n126 585
R247 B.n309 B.n308 585
R248 B.n310 B.n125 585
R249 B.n312 B.n311 585
R250 B.n313 B.n124 585
R251 B.n315 B.n314 585
R252 B.n316 B.n123 585
R253 B.n318 B.n317 585
R254 B.n319 B.n122 585
R255 B.n321 B.n320 585
R256 B.n322 B.n121 585
R257 B.n324 B.n323 585
R258 B.n325 B.n120 585
R259 B.n327 B.n326 585
R260 B.n328 B.n119 585
R261 B.n330 B.n329 585
R262 B.n331 B.n118 585
R263 B.n333 B.n332 585
R264 B.n334 B.n117 585
R265 B.n336 B.n335 585
R266 B.n337 B.n116 585
R267 B.n339 B.n338 585
R268 B.n340 B.n115 585
R269 B.n342 B.n341 585
R270 B.n343 B.n114 585
R271 B.n345 B.n344 585
R272 B.n346 B.n113 585
R273 B.n348 B.n347 585
R274 B.n349 B.n112 585
R275 B.n351 B.n350 585
R276 B.n352 B.n111 585
R277 B.n354 B.n353 585
R278 B.n355 B.n110 585
R279 B.n357 B.n356 585
R280 B.n358 B.n109 585
R281 B.n360 B.n359 585
R282 B.n361 B.n108 585
R283 B.n363 B.n362 585
R284 B.n364 B.n107 585
R285 B.n224 B.n223 585
R286 B.n222 B.n155 585
R287 B.n221 B.n220 585
R288 B.n219 B.n156 585
R289 B.n218 B.n217 585
R290 B.n216 B.n157 585
R291 B.n215 B.n214 585
R292 B.n213 B.n158 585
R293 B.n212 B.n211 585
R294 B.n210 B.n159 585
R295 B.n209 B.n208 585
R296 B.n207 B.n160 585
R297 B.n206 B.n205 585
R298 B.n204 B.n161 585
R299 B.n203 B.n202 585
R300 B.n201 B.n162 585
R301 B.n200 B.n199 585
R302 B.n198 B.n163 585
R303 B.n197 B.n196 585
R304 B.n195 B.n164 585
R305 B.n194 B.n193 585
R306 B.n192 B.n165 585
R307 B.n191 B.n190 585
R308 B.n189 B.n166 585
R309 B.n188 B.n187 585
R310 B.n186 B.n167 585
R311 B.n185 B.n184 585
R312 B.n183 B.n168 585
R313 B.n182 B.n181 585
R314 B.n180 B.n169 585
R315 B.n179 B.n178 585
R316 B.n177 B.n170 585
R317 B.n176 B.n175 585
R318 B.n174 B.n171 585
R319 B.n173 B.n172 585
R320 B.n2 B.n0 585
R321 B.n665 B.n1 585
R322 B.n664 B.n663 585
R323 B.n662 B.n3 585
R324 B.n661 B.n660 585
R325 B.n659 B.n4 585
R326 B.n658 B.n657 585
R327 B.n656 B.n5 585
R328 B.n655 B.n654 585
R329 B.n653 B.n6 585
R330 B.n652 B.n651 585
R331 B.n650 B.n7 585
R332 B.n649 B.n648 585
R333 B.n647 B.n8 585
R334 B.n646 B.n645 585
R335 B.n644 B.n9 585
R336 B.n643 B.n642 585
R337 B.n641 B.n10 585
R338 B.n640 B.n639 585
R339 B.n638 B.n11 585
R340 B.n637 B.n636 585
R341 B.n635 B.n12 585
R342 B.n634 B.n633 585
R343 B.n632 B.n13 585
R344 B.n631 B.n630 585
R345 B.n629 B.n14 585
R346 B.n628 B.n627 585
R347 B.n626 B.n15 585
R348 B.n625 B.n624 585
R349 B.n623 B.n16 585
R350 B.n622 B.n621 585
R351 B.n620 B.n17 585
R352 B.n619 B.n618 585
R353 B.n617 B.n18 585
R354 B.n616 B.n615 585
R355 B.n614 B.n19 585
R356 B.n613 B.n612 585
R357 B.n667 B.n666 585
R358 B.n223 B.n154 506.916
R359 B.n612 B.n611 506.916
R360 B.n365 B.n364 506.916
R361 B.n473 B.n70 506.916
R362 B.n299 B.t3 308.091
R363 B.n133 B.t0 308.091
R364 B.n42 B.t6 308.091
R365 B.n49 B.t9 308.091
R366 B.n299 B.t5 171.368
R367 B.n49 B.t10 171.368
R368 B.n133 B.t2 171.353
R369 B.n42 B.t7 171.353
R370 B.n223 B.n222 163.367
R371 B.n222 B.n221 163.367
R372 B.n221 B.n156 163.367
R373 B.n217 B.n156 163.367
R374 B.n217 B.n216 163.367
R375 B.n216 B.n215 163.367
R376 B.n215 B.n158 163.367
R377 B.n211 B.n158 163.367
R378 B.n211 B.n210 163.367
R379 B.n210 B.n209 163.367
R380 B.n209 B.n160 163.367
R381 B.n205 B.n160 163.367
R382 B.n205 B.n204 163.367
R383 B.n204 B.n203 163.367
R384 B.n203 B.n162 163.367
R385 B.n199 B.n162 163.367
R386 B.n199 B.n198 163.367
R387 B.n198 B.n197 163.367
R388 B.n197 B.n164 163.367
R389 B.n193 B.n164 163.367
R390 B.n193 B.n192 163.367
R391 B.n192 B.n191 163.367
R392 B.n191 B.n166 163.367
R393 B.n187 B.n166 163.367
R394 B.n187 B.n186 163.367
R395 B.n186 B.n185 163.367
R396 B.n185 B.n168 163.367
R397 B.n181 B.n168 163.367
R398 B.n181 B.n180 163.367
R399 B.n180 B.n179 163.367
R400 B.n179 B.n170 163.367
R401 B.n175 B.n170 163.367
R402 B.n175 B.n174 163.367
R403 B.n174 B.n173 163.367
R404 B.n173 B.n2 163.367
R405 B.n666 B.n2 163.367
R406 B.n666 B.n665 163.367
R407 B.n665 B.n664 163.367
R408 B.n664 B.n3 163.367
R409 B.n660 B.n3 163.367
R410 B.n660 B.n659 163.367
R411 B.n659 B.n658 163.367
R412 B.n658 B.n5 163.367
R413 B.n654 B.n5 163.367
R414 B.n654 B.n653 163.367
R415 B.n653 B.n652 163.367
R416 B.n652 B.n7 163.367
R417 B.n648 B.n7 163.367
R418 B.n648 B.n647 163.367
R419 B.n647 B.n646 163.367
R420 B.n646 B.n9 163.367
R421 B.n642 B.n9 163.367
R422 B.n642 B.n641 163.367
R423 B.n641 B.n640 163.367
R424 B.n640 B.n11 163.367
R425 B.n636 B.n11 163.367
R426 B.n636 B.n635 163.367
R427 B.n635 B.n634 163.367
R428 B.n634 B.n13 163.367
R429 B.n630 B.n13 163.367
R430 B.n630 B.n629 163.367
R431 B.n629 B.n628 163.367
R432 B.n628 B.n15 163.367
R433 B.n624 B.n15 163.367
R434 B.n624 B.n623 163.367
R435 B.n623 B.n622 163.367
R436 B.n622 B.n17 163.367
R437 B.n618 B.n17 163.367
R438 B.n618 B.n617 163.367
R439 B.n617 B.n616 163.367
R440 B.n616 B.n19 163.367
R441 B.n612 B.n19 163.367
R442 B.n227 B.n154 163.367
R443 B.n228 B.n227 163.367
R444 B.n229 B.n228 163.367
R445 B.n229 B.n152 163.367
R446 B.n233 B.n152 163.367
R447 B.n234 B.n233 163.367
R448 B.n235 B.n234 163.367
R449 B.n235 B.n150 163.367
R450 B.n239 B.n150 163.367
R451 B.n240 B.n239 163.367
R452 B.n241 B.n240 163.367
R453 B.n241 B.n148 163.367
R454 B.n245 B.n148 163.367
R455 B.n246 B.n245 163.367
R456 B.n247 B.n246 163.367
R457 B.n247 B.n146 163.367
R458 B.n251 B.n146 163.367
R459 B.n252 B.n251 163.367
R460 B.n253 B.n252 163.367
R461 B.n253 B.n144 163.367
R462 B.n257 B.n144 163.367
R463 B.n258 B.n257 163.367
R464 B.n259 B.n258 163.367
R465 B.n259 B.n142 163.367
R466 B.n263 B.n142 163.367
R467 B.n264 B.n263 163.367
R468 B.n265 B.n264 163.367
R469 B.n265 B.n140 163.367
R470 B.n269 B.n140 163.367
R471 B.n270 B.n269 163.367
R472 B.n271 B.n270 163.367
R473 B.n271 B.n138 163.367
R474 B.n275 B.n138 163.367
R475 B.n276 B.n275 163.367
R476 B.n277 B.n276 163.367
R477 B.n277 B.n136 163.367
R478 B.n281 B.n136 163.367
R479 B.n282 B.n281 163.367
R480 B.n283 B.n282 163.367
R481 B.n283 B.n132 163.367
R482 B.n288 B.n132 163.367
R483 B.n289 B.n288 163.367
R484 B.n290 B.n289 163.367
R485 B.n290 B.n130 163.367
R486 B.n294 B.n130 163.367
R487 B.n295 B.n294 163.367
R488 B.n296 B.n295 163.367
R489 B.n296 B.n128 163.367
R490 B.n303 B.n128 163.367
R491 B.n304 B.n303 163.367
R492 B.n305 B.n304 163.367
R493 B.n305 B.n126 163.367
R494 B.n309 B.n126 163.367
R495 B.n310 B.n309 163.367
R496 B.n311 B.n310 163.367
R497 B.n311 B.n124 163.367
R498 B.n315 B.n124 163.367
R499 B.n316 B.n315 163.367
R500 B.n317 B.n316 163.367
R501 B.n317 B.n122 163.367
R502 B.n321 B.n122 163.367
R503 B.n322 B.n321 163.367
R504 B.n323 B.n322 163.367
R505 B.n323 B.n120 163.367
R506 B.n327 B.n120 163.367
R507 B.n328 B.n327 163.367
R508 B.n329 B.n328 163.367
R509 B.n329 B.n118 163.367
R510 B.n333 B.n118 163.367
R511 B.n334 B.n333 163.367
R512 B.n335 B.n334 163.367
R513 B.n335 B.n116 163.367
R514 B.n339 B.n116 163.367
R515 B.n340 B.n339 163.367
R516 B.n341 B.n340 163.367
R517 B.n341 B.n114 163.367
R518 B.n345 B.n114 163.367
R519 B.n346 B.n345 163.367
R520 B.n347 B.n346 163.367
R521 B.n347 B.n112 163.367
R522 B.n351 B.n112 163.367
R523 B.n352 B.n351 163.367
R524 B.n353 B.n352 163.367
R525 B.n353 B.n110 163.367
R526 B.n357 B.n110 163.367
R527 B.n358 B.n357 163.367
R528 B.n359 B.n358 163.367
R529 B.n359 B.n108 163.367
R530 B.n363 B.n108 163.367
R531 B.n364 B.n363 163.367
R532 B.n365 B.n106 163.367
R533 B.n369 B.n106 163.367
R534 B.n370 B.n369 163.367
R535 B.n371 B.n370 163.367
R536 B.n371 B.n104 163.367
R537 B.n375 B.n104 163.367
R538 B.n376 B.n375 163.367
R539 B.n377 B.n376 163.367
R540 B.n377 B.n102 163.367
R541 B.n381 B.n102 163.367
R542 B.n382 B.n381 163.367
R543 B.n383 B.n382 163.367
R544 B.n383 B.n100 163.367
R545 B.n387 B.n100 163.367
R546 B.n388 B.n387 163.367
R547 B.n389 B.n388 163.367
R548 B.n389 B.n98 163.367
R549 B.n393 B.n98 163.367
R550 B.n394 B.n393 163.367
R551 B.n395 B.n394 163.367
R552 B.n395 B.n96 163.367
R553 B.n399 B.n96 163.367
R554 B.n400 B.n399 163.367
R555 B.n401 B.n400 163.367
R556 B.n401 B.n94 163.367
R557 B.n405 B.n94 163.367
R558 B.n406 B.n405 163.367
R559 B.n407 B.n406 163.367
R560 B.n407 B.n92 163.367
R561 B.n411 B.n92 163.367
R562 B.n412 B.n411 163.367
R563 B.n413 B.n412 163.367
R564 B.n413 B.n90 163.367
R565 B.n417 B.n90 163.367
R566 B.n418 B.n417 163.367
R567 B.n419 B.n418 163.367
R568 B.n419 B.n88 163.367
R569 B.n423 B.n88 163.367
R570 B.n424 B.n423 163.367
R571 B.n425 B.n424 163.367
R572 B.n425 B.n86 163.367
R573 B.n429 B.n86 163.367
R574 B.n430 B.n429 163.367
R575 B.n431 B.n430 163.367
R576 B.n431 B.n84 163.367
R577 B.n435 B.n84 163.367
R578 B.n436 B.n435 163.367
R579 B.n437 B.n436 163.367
R580 B.n437 B.n82 163.367
R581 B.n441 B.n82 163.367
R582 B.n442 B.n441 163.367
R583 B.n443 B.n442 163.367
R584 B.n443 B.n80 163.367
R585 B.n447 B.n80 163.367
R586 B.n448 B.n447 163.367
R587 B.n449 B.n448 163.367
R588 B.n449 B.n78 163.367
R589 B.n453 B.n78 163.367
R590 B.n454 B.n453 163.367
R591 B.n455 B.n454 163.367
R592 B.n455 B.n76 163.367
R593 B.n459 B.n76 163.367
R594 B.n460 B.n459 163.367
R595 B.n461 B.n460 163.367
R596 B.n461 B.n74 163.367
R597 B.n465 B.n74 163.367
R598 B.n466 B.n465 163.367
R599 B.n467 B.n466 163.367
R600 B.n467 B.n72 163.367
R601 B.n471 B.n72 163.367
R602 B.n472 B.n471 163.367
R603 B.n473 B.n472 163.367
R604 B.n611 B.n610 163.367
R605 B.n610 B.n21 163.367
R606 B.n606 B.n21 163.367
R607 B.n606 B.n605 163.367
R608 B.n605 B.n604 163.367
R609 B.n604 B.n23 163.367
R610 B.n600 B.n23 163.367
R611 B.n600 B.n599 163.367
R612 B.n599 B.n598 163.367
R613 B.n598 B.n25 163.367
R614 B.n594 B.n25 163.367
R615 B.n594 B.n593 163.367
R616 B.n593 B.n592 163.367
R617 B.n592 B.n27 163.367
R618 B.n588 B.n27 163.367
R619 B.n588 B.n587 163.367
R620 B.n587 B.n586 163.367
R621 B.n586 B.n29 163.367
R622 B.n582 B.n29 163.367
R623 B.n582 B.n581 163.367
R624 B.n581 B.n580 163.367
R625 B.n580 B.n31 163.367
R626 B.n576 B.n31 163.367
R627 B.n576 B.n575 163.367
R628 B.n575 B.n574 163.367
R629 B.n574 B.n33 163.367
R630 B.n570 B.n33 163.367
R631 B.n570 B.n569 163.367
R632 B.n569 B.n568 163.367
R633 B.n568 B.n35 163.367
R634 B.n564 B.n35 163.367
R635 B.n564 B.n563 163.367
R636 B.n563 B.n562 163.367
R637 B.n562 B.n37 163.367
R638 B.n558 B.n37 163.367
R639 B.n558 B.n557 163.367
R640 B.n557 B.n556 163.367
R641 B.n556 B.n39 163.367
R642 B.n552 B.n39 163.367
R643 B.n552 B.n551 163.367
R644 B.n551 B.n550 163.367
R645 B.n550 B.n41 163.367
R646 B.n546 B.n41 163.367
R647 B.n546 B.n545 163.367
R648 B.n545 B.n544 163.367
R649 B.n544 B.n46 163.367
R650 B.n540 B.n46 163.367
R651 B.n540 B.n539 163.367
R652 B.n539 B.n538 163.367
R653 B.n538 B.n48 163.367
R654 B.n533 B.n48 163.367
R655 B.n533 B.n532 163.367
R656 B.n532 B.n531 163.367
R657 B.n531 B.n52 163.367
R658 B.n527 B.n52 163.367
R659 B.n527 B.n526 163.367
R660 B.n526 B.n525 163.367
R661 B.n525 B.n54 163.367
R662 B.n521 B.n54 163.367
R663 B.n521 B.n520 163.367
R664 B.n520 B.n519 163.367
R665 B.n519 B.n56 163.367
R666 B.n515 B.n56 163.367
R667 B.n515 B.n514 163.367
R668 B.n514 B.n513 163.367
R669 B.n513 B.n58 163.367
R670 B.n509 B.n58 163.367
R671 B.n509 B.n508 163.367
R672 B.n508 B.n507 163.367
R673 B.n507 B.n60 163.367
R674 B.n503 B.n60 163.367
R675 B.n503 B.n502 163.367
R676 B.n502 B.n501 163.367
R677 B.n501 B.n62 163.367
R678 B.n497 B.n62 163.367
R679 B.n497 B.n496 163.367
R680 B.n496 B.n495 163.367
R681 B.n495 B.n64 163.367
R682 B.n491 B.n64 163.367
R683 B.n491 B.n490 163.367
R684 B.n490 B.n489 163.367
R685 B.n489 B.n66 163.367
R686 B.n485 B.n66 163.367
R687 B.n485 B.n484 163.367
R688 B.n484 B.n483 163.367
R689 B.n483 B.n68 163.367
R690 B.n479 B.n68 163.367
R691 B.n479 B.n478 163.367
R692 B.n478 B.n477 163.367
R693 B.n477 B.n70 163.367
R694 B.n300 B.t4 110.082
R695 B.n50 B.t11 110.082
R696 B.n134 B.t1 110.069
R697 B.n43 B.t8 110.069
R698 B.n300 B.n299 61.2853
R699 B.n134 B.n133 61.2853
R700 B.n43 B.n42 61.2853
R701 B.n50 B.n49 61.2853
R702 B.n301 B.n300 59.5399
R703 B.n286 B.n134 59.5399
R704 B.n44 B.n43 59.5399
R705 B.n536 B.n50 59.5399
R706 B.n613 B.n20 32.9371
R707 B.n475 B.n474 32.9371
R708 B.n366 B.n107 32.9371
R709 B.n225 B.n224 32.9371
R710 B B.n667 18.0485
R711 B.n609 B.n20 10.6151
R712 B.n609 B.n608 10.6151
R713 B.n608 B.n607 10.6151
R714 B.n607 B.n22 10.6151
R715 B.n603 B.n22 10.6151
R716 B.n603 B.n602 10.6151
R717 B.n602 B.n601 10.6151
R718 B.n601 B.n24 10.6151
R719 B.n597 B.n24 10.6151
R720 B.n597 B.n596 10.6151
R721 B.n596 B.n595 10.6151
R722 B.n595 B.n26 10.6151
R723 B.n591 B.n26 10.6151
R724 B.n591 B.n590 10.6151
R725 B.n590 B.n589 10.6151
R726 B.n589 B.n28 10.6151
R727 B.n585 B.n28 10.6151
R728 B.n585 B.n584 10.6151
R729 B.n584 B.n583 10.6151
R730 B.n583 B.n30 10.6151
R731 B.n579 B.n30 10.6151
R732 B.n579 B.n578 10.6151
R733 B.n578 B.n577 10.6151
R734 B.n577 B.n32 10.6151
R735 B.n573 B.n32 10.6151
R736 B.n573 B.n572 10.6151
R737 B.n572 B.n571 10.6151
R738 B.n571 B.n34 10.6151
R739 B.n567 B.n34 10.6151
R740 B.n567 B.n566 10.6151
R741 B.n566 B.n565 10.6151
R742 B.n565 B.n36 10.6151
R743 B.n561 B.n36 10.6151
R744 B.n561 B.n560 10.6151
R745 B.n560 B.n559 10.6151
R746 B.n559 B.n38 10.6151
R747 B.n555 B.n38 10.6151
R748 B.n555 B.n554 10.6151
R749 B.n554 B.n553 10.6151
R750 B.n553 B.n40 10.6151
R751 B.n549 B.n548 10.6151
R752 B.n548 B.n547 10.6151
R753 B.n547 B.n45 10.6151
R754 B.n543 B.n45 10.6151
R755 B.n543 B.n542 10.6151
R756 B.n542 B.n541 10.6151
R757 B.n541 B.n47 10.6151
R758 B.n537 B.n47 10.6151
R759 B.n535 B.n534 10.6151
R760 B.n534 B.n51 10.6151
R761 B.n530 B.n51 10.6151
R762 B.n530 B.n529 10.6151
R763 B.n529 B.n528 10.6151
R764 B.n528 B.n53 10.6151
R765 B.n524 B.n53 10.6151
R766 B.n524 B.n523 10.6151
R767 B.n523 B.n522 10.6151
R768 B.n522 B.n55 10.6151
R769 B.n518 B.n55 10.6151
R770 B.n518 B.n517 10.6151
R771 B.n517 B.n516 10.6151
R772 B.n516 B.n57 10.6151
R773 B.n512 B.n57 10.6151
R774 B.n512 B.n511 10.6151
R775 B.n511 B.n510 10.6151
R776 B.n510 B.n59 10.6151
R777 B.n506 B.n59 10.6151
R778 B.n506 B.n505 10.6151
R779 B.n505 B.n504 10.6151
R780 B.n504 B.n61 10.6151
R781 B.n500 B.n61 10.6151
R782 B.n500 B.n499 10.6151
R783 B.n499 B.n498 10.6151
R784 B.n498 B.n63 10.6151
R785 B.n494 B.n63 10.6151
R786 B.n494 B.n493 10.6151
R787 B.n493 B.n492 10.6151
R788 B.n492 B.n65 10.6151
R789 B.n488 B.n65 10.6151
R790 B.n488 B.n487 10.6151
R791 B.n487 B.n486 10.6151
R792 B.n486 B.n67 10.6151
R793 B.n482 B.n67 10.6151
R794 B.n482 B.n481 10.6151
R795 B.n481 B.n480 10.6151
R796 B.n480 B.n69 10.6151
R797 B.n476 B.n69 10.6151
R798 B.n476 B.n475 10.6151
R799 B.n367 B.n366 10.6151
R800 B.n368 B.n367 10.6151
R801 B.n368 B.n105 10.6151
R802 B.n372 B.n105 10.6151
R803 B.n373 B.n372 10.6151
R804 B.n374 B.n373 10.6151
R805 B.n374 B.n103 10.6151
R806 B.n378 B.n103 10.6151
R807 B.n379 B.n378 10.6151
R808 B.n380 B.n379 10.6151
R809 B.n380 B.n101 10.6151
R810 B.n384 B.n101 10.6151
R811 B.n385 B.n384 10.6151
R812 B.n386 B.n385 10.6151
R813 B.n386 B.n99 10.6151
R814 B.n390 B.n99 10.6151
R815 B.n391 B.n390 10.6151
R816 B.n392 B.n391 10.6151
R817 B.n392 B.n97 10.6151
R818 B.n396 B.n97 10.6151
R819 B.n397 B.n396 10.6151
R820 B.n398 B.n397 10.6151
R821 B.n398 B.n95 10.6151
R822 B.n402 B.n95 10.6151
R823 B.n403 B.n402 10.6151
R824 B.n404 B.n403 10.6151
R825 B.n404 B.n93 10.6151
R826 B.n408 B.n93 10.6151
R827 B.n409 B.n408 10.6151
R828 B.n410 B.n409 10.6151
R829 B.n410 B.n91 10.6151
R830 B.n414 B.n91 10.6151
R831 B.n415 B.n414 10.6151
R832 B.n416 B.n415 10.6151
R833 B.n416 B.n89 10.6151
R834 B.n420 B.n89 10.6151
R835 B.n421 B.n420 10.6151
R836 B.n422 B.n421 10.6151
R837 B.n422 B.n87 10.6151
R838 B.n426 B.n87 10.6151
R839 B.n427 B.n426 10.6151
R840 B.n428 B.n427 10.6151
R841 B.n428 B.n85 10.6151
R842 B.n432 B.n85 10.6151
R843 B.n433 B.n432 10.6151
R844 B.n434 B.n433 10.6151
R845 B.n434 B.n83 10.6151
R846 B.n438 B.n83 10.6151
R847 B.n439 B.n438 10.6151
R848 B.n440 B.n439 10.6151
R849 B.n440 B.n81 10.6151
R850 B.n444 B.n81 10.6151
R851 B.n445 B.n444 10.6151
R852 B.n446 B.n445 10.6151
R853 B.n446 B.n79 10.6151
R854 B.n450 B.n79 10.6151
R855 B.n451 B.n450 10.6151
R856 B.n452 B.n451 10.6151
R857 B.n452 B.n77 10.6151
R858 B.n456 B.n77 10.6151
R859 B.n457 B.n456 10.6151
R860 B.n458 B.n457 10.6151
R861 B.n458 B.n75 10.6151
R862 B.n462 B.n75 10.6151
R863 B.n463 B.n462 10.6151
R864 B.n464 B.n463 10.6151
R865 B.n464 B.n73 10.6151
R866 B.n468 B.n73 10.6151
R867 B.n469 B.n468 10.6151
R868 B.n470 B.n469 10.6151
R869 B.n470 B.n71 10.6151
R870 B.n474 B.n71 10.6151
R871 B.n226 B.n225 10.6151
R872 B.n226 B.n153 10.6151
R873 B.n230 B.n153 10.6151
R874 B.n231 B.n230 10.6151
R875 B.n232 B.n231 10.6151
R876 B.n232 B.n151 10.6151
R877 B.n236 B.n151 10.6151
R878 B.n237 B.n236 10.6151
R879 B.n238 B.n237 10.6151
R880 B.n238 B.n149 10.6151
R881 B.n242 B.n149 10.6151
R882 B.n243 B.n242 10.6151
R883 B.n244 B.n243 10.6151
R884 B.n244 B.n147 10.6151
R885 B.n248 B.n147 10.6151
R886 B.n249 B.n248 10.6151
R887 B.n250 B.n249 10.6151
R888 B.n250 B.n145 10.6151
R889 B.n254 B.n145 10.6151
R890 B.n255 B.n254 10.6151
R891 B.n256 B.n255 10.6151
R892 B.n256 B.n143 10.6151
R893 B.n260 B.n143 10.6151
R894 B.n261 B.n260 10.6151
R895 B.n262 B.n261 10.6151
R896 B.n262 B.n141 10.6151
R897 B.n266 B.n141 10.6151
R898 B.n267 B.n266 10.6151
R899 B.n268 B.n267 10.6151
R900 B.n268 B.n139 10.6151
R901 B.n272 B.n139 10.6151
R902 B.n273 B.n272 10.6151
R903 B.n274 B.n273 10.6151
R904 B.n274 B.n137 10.6151
R905 B.n278 B.n137 10.6151
R906 B.n279 B.n278 10.6151
R907 B.n280 B.n279 10.6151
R908 B.n280 B.n135 10.6151
R909 B.n284 B.n135 10.6151
R910 B.n285 B.n284 10.6151
R911 B.n287 B.n131 10.6151
R912 B.n291 B.n131 10.6151
R913 B.n292 B.n291 10.6151
R914 B.n293 B.n292 10.6151
R915 B.n293 B.n129 10.6151
R916 B.n297 B.n129 10.6151
R917 B.n298 B.n297 10.6151
R918 B.n302 B.n298 10.6151
R919 B.n306 B.n127 10.6151
R920 B.n307 B.n306 10.6151
R921 B.n308 B.n307 10.6151
R922 B.n308 B.n125 10.6151
R923 B.n312 B.n125 10.6151
R924 B.n313 B.n312 10.6151
R925 B.n314 B.n313 10.6151
R926 B.n314 B.n123 10.6151
R927 B.n318 B.n123 10.6151
R928 B.n319 B.n318 10.6151
R929 B.n320 B.n319 10.6151
R930 B.n320 B.n121 10.6151
R931 B.n324 B.n121 10.6151
R932 B.n325 B.n324 10.6151
R933 B.n326 B.n325 10.6151
R934 B.n326 B.n119 10.6151
R935 B.n330 B.n119 10.6151
R936 B.n331 B.n330 10.6151
R937 B.n332 B.n331 10.6151
R938 B.n332 B.n117 10.6151
R939 B.n336 B.n117 10.6151
R940 B.n337 B.n336 10.6151
R941 B.n338 B.n337 10.6151
R942 B.n338 B.n115 10.6151
R943 B.n342 B.n115 10.6151
R944 B.n343 B.n342 10.6151
R945 B.n344 B.n343 10.6151
R946 B.n344 B.n113 10.6151
R947 B.n348 B.n113 10.6151
R948 B.n349 B.n348 10.6151
R949 B.n350 B.n349 10.6151
R950 B.n350 B.n111 10.6151
R951 B.n354 B.n111 10.6151
R952 B.n355 B.n354 10.6151
R953 B.n356 B.n355 10.6151
R954 B.n356 B.n109 10.6151
R955 B.n360 B.n109 10.6151
R956 B.n361 B.n360 10.6151
R957 B.n362 B.n361 10.6151
R958 B.n362 B.n107 10.6151
R959 B.n224 B.n155 10.6151
R960 B.n220 B.n155 10.6151
R961 B.n220 B.n219 10.6151
R962 B.n219 B.n218 10.6151
R963 B.n218 B.n157 10.6151
R964 B.n214 B.n157 10.6151
R965 B.n214 B.n213 10.6151
R966 B.n213 B.n212 10.6151
R967 B.n212 B.n159 10.6151
R968 B.n208 B.n159 10.6151
R969 B.n208 B.n207 10.6151
R970 B.n207 B.n206 10.6151
R971 B.n206 B.n161 10.6151
R972 B.n202 B.n161 10.6151
R973 B.n202 B.n201 10.6151
R974 B.n201 B.n200 10.6151
R975 B.n200 B.n163 10.6151
R976 B.n196 B.n163 10.6151
R977 B.n196 B.n195 10.6151
R978 B.n195 B.n194 10.6151
R979 B.n194 B.n165 10.6151
R980 B.n190 B.n165 10.6151
R981 B.n190 B.n189 10.6151
R982 B.n189 B.n188 10.6151
R983 B.n188 B.n167 10.6151
R984 B.n184 B.n167 10.6151
R985 B.n184 B.n183 10.6151
R986 B.n183 B.n182 10.6151
R987 B.n182 B.n169 10.6151
R988 B.n178 B.n169 10.6151
R989 B.n178 B.n177 10.6151
R990 B.n177 B.n176 10.6151
R991 B.n176 B.n171 10.6151
R992 B.n172 B.n171 10.6151
R993 B.n172 B.n0 10.6151
R994 B.n663 B.n1 10.6151
R995 B.n663 B.n662 10.6151
R996 B.n662 B.n661 10.6151
R997 B.n661 B.n4 10.6151
R998 B.n657 B.n4 10.6151
R999 B.n657 B.n656 10.6151
R1000 B.n656 B.n655 10.6151
R1001 B.n655 B.n6 10.6151
R1002 B.n651 B.n6 10.6151
R1003 B.n651 B.n650 10.6151
R1004 B.n650 B.n649 10.6151
R1005 B.n649 B.n8 10.6151
R1006 B.n645 B.n8 10.6151
R1007 B.n645 B.n644 10.6151
R1008 B.n644 B.n643 10.6151
R1009 B.n643 B.n10 10.6151
R1010 B.n639 B.n10 10.6151
R1011 B.n639 B.n638 10.6151
R1012 B.n638 B.n637 10.6151
R1013 B.n637 B.n12 10.6151
R1014 B.n633 B.n12 10.6151
R1015 B.n633 B.n632 10.6151
R1016 B.n632 B.n631 10.6151
R1017 B.n631 B.n14 10.6151
R1018 B.n627 B.n14 10.6151
R1019 B.n627 B.n626 10.6151
R1020 B.n626 B.n625 10.6151
R1021 B.n625 B.n16 10.6151
R1022 B.n621 B.n16 10.6151
R1023 B.n621 B.n620 10.6151
R1024 B.n620 B.n619 10.6151
R1025 B.n619 B.n18 10.6151
R1026 B.n615 B.n18 10.6151
R1027 B.n615 B.n614 10.6151
R1028 B.n614 B.n613 10.6151
R1029 B.n549 B.n44 6.5566
R1030 B.n537 B.n536 6.5566
R1031 B.n287 B.n286 6.5566
R1032 B.n302 B.n301 6.5566
R1033 B.n44 B.n40 4.05904
R1034 B.n536 B.n535 4.05904
R1035 B.n286 B.n285 4.05904
R1036 B.n301 B.n127 4.05904
R1037 B.n667 B.n0 2.81026
R1038 B.n667 B.n1 2.81026
R1039 VP.n16 VP.n0 161.3
R1040 VP.n15 VP.n14 161.3
R1041 VP.n13 VP.n1 161.3
R1042 VP.n12 VP.n11 161.3
R1043 VP.n10 VP.n2 161.3
R1044 VP.n9 VP.n8 161.3
R1045 VP.n7 VP.n3 161.3
R1046 VP.n4 VP.t3 134.948
R1047 VP.n4 VP.t1 134.054
R1048 VP.n6 VP.n5 106.841
R1049 VP.n18 VP.n17 106.841
R1050 VP.n5 VP.t2 99.7217
R1051 VP.n17 VP.t0 99.7217
R1052 VP.n6 VP.n4 50.2582
R1053 VP.n11 VP.n10 40.4934
R1054 VP.n11 VP.n1 40.4934
R1055 VP.n9 VP.n3 24.4675
R1056 VP.n10 VP.n9 24.4675
R1057 VP.n15 VP.n1 24.4675
R1058 VP.n16 VP.n15 24.4675
R1059 VP.n5 VP.n3 3.91522
R1060 VP.n17 VP.n16 3.91522
R1061 VP.n7 VP.n6 0.278367
R1062 VP.n18 VP.n0 0.278367
R1063 VP.n8 VP.n7 0.189894
R1064 VP.n8 VP.n2 0.189894
R1065 VP.n12 VP.n2 0.189894
R1066 VP.n13 VP.n12 0.189894
R1067 VP.n14 VP.n13 0.189894
R1068 VP.n14 VP.n0 0.189894
R1069 VP VP.n18 0.153454
R1070 VDD1 VDD1.n1 115.832
R1071 VDD1 VDD1.n0 73.3832
R1072 VDD1.n0 VDD1.t0 2.77633
R1073 VDD1.n0 VDD1.t2 2.77633
R1074 VDD1.n1 VDD1.t1 2.77633
R1075 VDD1.n1 VDD1.t3 2.77633
C0 VDD1 VN 0.149046f
C1 w_n2866_n3310# VN 4.89041f
C2 B VP 1.7624f
C3 VTAIL VP 4.68323f
C4 VDD2 VDD1 1.07745f
C5 VTAIL B 4.95121f
C6 w_n2866_n3310# VDD2 1.54785f
C7 VP VN 6.30209f
C8 w_n2866_n3310# VDD1 1.48664f
C9 B VN 1.14896f
C10 VTAIL VN 4.66912f
C11 VDD2 VP 0.408779f
C12 B VDD2 1.34987f
C13 VP VDD1 4.97468f
C14 w_n2866_n3310# VP 5.25942f
C15 VTAIL VDD2 5.43886f
C16 B VDD1 1.29391f
C17 B w_n2866_n3310# 9.44755f
C18 VTAIL VDD1 5.38311f
C19 VTAIL w_n2866_n3310# 3.91573f
C20 VDD2 VN 4.71574f
C21 VDD2 VSUBS 0.978996f
C22 VDD1 VSUBS 5.85718f
C23 VTAIL VSUBS 1.228812f
C24 VN VSUBS 5.55728f
C25 VP VSUBS 2.387607f
C26 B VSUBS 4.450267f
C27 w_n2866_n3310# VSUBS 0.11683p
C28 VDD1.t0 VSUBS 0.252925f
C29 VDD1.t2 VSUBS 0.252925f
C30 VDD1.n0 VSUBS 1.96181f
C31 VDD1.t1 VSUBS 0.252925f
C32 VDD1.t3 VSUBS 0.252925f
C33 VDD1.n1 VSUBS 2.7113f
C34 VP.n0 VSUBS 0.043391f
C35 VP.t0 VSUBS 2.96955f
C36 VP.n1 VSUBS 0.065411f
C37 VP.n2 VSUBS 0.032911f
C38 VP.n3 VSUBS 0.035901f
C39 VP.t1 VSUBS 3.29505f
C40 VP.t3 VSUBS 3.30324f
C41 VP.n4 VSUBS 3.90781f
C42 VP.t2 VSUBS 2.96955f
C43 VP.n5 VSUBS 1.15859f
C44 VP.n6 VSUBS 1.83104f
C45 VP.n7 VSUBS 0.043391f
C46 VP.n8 VSUBS 0.032911f
C47 VP.n9 VSUBS 0.061339f
C48 VP.n10 VSUBS 0.065411f
C49 VP.n11 VSUBS 0.026606f
C50 VP.n12 VSUBS 0.032911f
C51 VP.n13 VSUBS 0.032911f
C52 VP.n14 VSUBS 0.032911f
C53 VP.n15 VSUBS 0.061339f
C54 VP.n16 VSUBS 0.035901f
C55 VP.n17 VSUBS 1.15859f
C56 VP.n18 VSUBS 0.061037f
C57 B.n0 VSUBS 0.0042f
C58 B.n1 VSUBS 0.0042f
C59 B.n2 VSUBS 0.006642f
C60 B.n3 VSUBS 0.006642f
C61 B.n4 VSUBS 0.006642f
C62 B.n5 VSUBS 0.006642f
C63 B.n6 VSUBS 0.006642f
C64 B.n7 VSUBS 0.006642f
C65 B.n8 VSUBS 0.006642f
C66 B.n9 VSUBS 0.006642f
C67 B.n10 VSUBS 0.006642f
C68 B.n11 VSUBS 0.006642f
C69 B.n12 VSUBS 0.006642f
C70 B.n13 VSUBS 0.006642f
C71 B.n14 VSUBS 0.006642f
C72 B.n15 VSUBS 0.006642f
C73 B.n16 VSUBS 0.006642f
C74 B.n17 VSUBS 0.006642f
C75 B.n18 VSUBS 0.006642f
C76 B.n19 VSUBS 0.006642f
C77 B.n20 VSUBS 0.01596f
C78 B.n21 VSUBS 0.006642f
C79 B.n22 VSUBS 0.006642f
C80 B.n23 VSUBS 0.006642f
C81 B.n24 VSUBS 0.006642f
C82 B.n25 VSUBS 0.006642f
C83 B.n26 VSUBS 0.006642f
C84 B.n27 VSUBS 0.006642f
C85 B.n28 VSUBS 0.006642f
C86 B.n29 VSUBS 0.006642f
C87 B.n30 VSUBS 0.006642f
C88 B.n31 VSUBS 0.006642f
C89 B.n32 VSUBS 0.006642f
C90 B.n33 VSUBS 0.006642f
C91 B.n34 VSUBS 0.006642f
C92 B.n35 VSUBS 0.006642f
C93 B.n36 VSUBS 0.006642f
C94 B.n37 VSUBS 0.006642f
C95 B.n38 VSUBS 0.006642f
C96 B.n39 VSUBS 0.006642f
C97 B.n40 VSUBS 0.004591f
C98 B.n41 VSUBS 0.006642f
C99 B.t8 VSUBS 0.361127f
C100 B.t7 VSUBS 0.382418f
C101 B.t6 VSUBS 1.44239f
C102 B.n42 VSUBS 0.204816f
C103 B.n43 VSUBS 0.069002f
C104 B.n44 VSUBS 0.015388f
C105 B.n45 VSUBS 0.006642f
C106 B.n46 VSUBS 0.006642f
C107 B.n47 VSUBS 0.006642f
C108 B.n48 VSUBS 0.006642f
C109 B.t11 VSUBS 0.36112f
C110 B.t10 VSUBS 0.382411f
C111 B.t9 VSUBS 1.44239f
C112 B.n49 VSUBS 0.204822f
C113 B.n50 VSUBS 0.069008f
C114 B.n51 VSUBS 0.006642f
C115 B.n52 VSUBS 0.006642f
C116 B.n53 VSUBS 0.006642f
C117 B.n54 VSUBS 0.006642f
C118 B.n55 VSUBS 0.006642f
C119 B.n56 VSUBS 0.006642f
C120 B.n57 VSUBS 0.006642f
C121 B.n58 VSUBS 0.006642f
C122 B.n59 VSUBS 0.006642f
C123 B.n60 VSUBS 0.006642f
C124 B.n61 VSUBS 0.006642f
C125 B.n62 VSUBS 0.006642f
C126 B.n63 VSUBS 0.006642f
C127 B.n64 VSUBS 0.006642f
C128 B.n65 VSUBS 0.006642f
C129 B.n66 VSUBS 0.006642f
C130 B.n67 VSUBS 0.006642f
C131 B.n68 VSUBS 0.006642f
C132 B.n69 VSUBS 0.006642f
C133 B.n70 VSUBS 0.01596f
C134 B.n71 VSUBS 0.006642f
C135 B.n72 VSUBS 0.006642f
C136 B.n73 VSUBS 0.006642f
C137 B.n74 VSUBS 0.006642f
C138 B.n75 VSUBS 0.006642f
C139 B.n76 VSUBS 0.006642f
C140 B.n77 VSUBS 0.006642f
C141 B.n78 VSUBS 0.006642f
C142 B.n79 VSUBS 0.006642f
C143 B.n80 VSUBS 0.006642f
C144 B.n81 VSUBS 0.006642f
C145 B.n82 VSUBS 0.006642f
C146 B.n83 VSUBS 0.006642f
C147 B.n84 VSUBS 0.006642f
C148 B.n85 VSUBS 0.006642f
C149 B.n86 VSUBS 0.006642f
C150 B.n87 VSUBS 0.006642f
C151 B.n88 VSUBS 0.006642f
C152 B.n89 VSUBS 0.006642f
C153 B.n90 VSUBS 0.006642f
C154 B.n91 VSUBS 0.006642f
C155 B.n92 VSUBS 0.006642f
C156 B.n93 VSUBS 0.006642f
C157 B.n94 VSUBS 0.006642f
C158 B.n95 VSUBS 0.006642f
C159 B.n96 VSUBS 0.006642f
C160 B.n97 VSUBS 0.006642f
C161 B.n98 VSUBS 0.006642f
C162 B.n99 VSUBS 0.006642f
C163 B.n100 VSUBS 0.006642f
C164 B.n101 VSUBS 0.006642f
C165 B.n102 VSUBS 0.006642f
C166 B.n103 VSUBS 0.006642f
C167 B.n104 VSUBS 0.006642f
C168 B.n105 VSUBS 0.006642f
C169 B.n106 VSUBS 0.006642f
C170 B.n107 VSUBS 0.01596f
C171 B.n108 VSUBS 0.006642f
C172 B.n109 VSUBS 0.006642f
C173 B.n110 VSUBS 0.006642f
C174 B.n111 VSUBS 0.006642f
C175 B.n112 VSUBS 0.006642f
C176 B.n113 VSUBS 0.006642f
C177 B.n114 VSUBS 0.006642f
C178 B.n115 VSUBS 0.006642f
C179 B.n116 VSUBS 0.006642f
C180 B.n117 VSUBS 0.006642f
C181 B.n118 VSUBS 0.006642f
C182 B.n119 VSUBS 0.006642f
C183 B.n120 VSUBS 0.006642f
C184 B.n121 VSUBS 0.006642f
C185 B.n122 VSUBS 0.006642f
C186 B.n123 VSUBS 0.006642f
C187 B.n124 VSUBS 0.006642f
C188 B.n125 VSUBS 0.006642f
C189 B.n126 VSUBS 0.006642f
C190 B.n127 VSUBS 0.004591f
C191 B.n128 VSUBS 0.006642f
C192 B.n129 VSUBS 0.006642f
C193 B.n130 VSUBS 0.006642f
C194 B.n131 VSUBS 0.006642f
C195 B.n132 VSUBS 0.006642f
C196 B.t1 VSUBS 0.361127f
C197 B.t2 VSUBS 0.382418f
C198 B.t0 VSUBS 1.44239f
C199 B.n133 VSUBS 0.204816f
C200 B.n134 VSUBS 0.069002f
C201 B.n135 VSUBS 0.006642f
C202 B.n136 VSUBS 0.006642f
C203 B.n137 VSUBS 0.006642f
C204 B.n138 VSUBS 0.006642f
C205 B.n139 VSUBS 0.006642f
C206 B.n140 VSUBS 0.006642f
C207 B.n141 VSUBS 0.006642f
C208 B.n142 VSUBS 0.006642f
C209 B.n143 VSUBS 0.006642f
C210 B.n144 VSUBS 0.006642f
C211 B.n145 VSUBS 0.006642f
C212 B.n146 VSUBS 0.006642f
C213 B.n147 VSUBS 0.006642f
C214 B.n148 VSUBS 0.006642f
C215 B.n149 VSUBS 0.006642f
C216 B.n150 VSUBS 0.006642f
C217 B.n151 VSUBS 0.006642f
C218 B.n152 VSUBS 0.006642f
C219 B.n153 VSUBS 0.006642f
C220 B.n154 VSUBS 0.01596f
C221 B.n155 VSUBS 0.006642f
C222 B.n156 VSUBS 0.006642f
C223 B.n157 VSUBS 0.006642f
C224 B.n158 VSUBS 0.006642f
C225 B.n159 VSUBS 0.006642f
C226 B.n160 VSUBS 0.006642f
C227 B.n161 VSUBS 0.006642f
C228 B.n162 VSUBS 0.006642f
C229 B.n163 VSUBS 0.006642f
C230 B.n164 VSUBS 0.006642f
C231 B.n165 VSUBS 0.006642f
C232 B.n166 VSUBS 0.006642f
C233 B.n167 VSUBS 0.006642f
C234 B.n168 VSUBS 0.006642f
C235 B.n169 VSUBS 0.006642f
C236 B.n170 VSUBS 0.006642f
C237 B.n171 VSUBS 0.006642f
C238 B.n172 VSUBS 0.006642f
C239 B.n173 VSUBS 0.006642f
C240 B.n174 VSUBS 0.006642f
C241 B.n175 VSUBS 0.006642f
C242 B.n176 VSUBS 0.006642f
C243 B.n177 VSUBS 0.006642f
C244 B.n178 VSUBS 0.006642f
C245 B.n179 VSUBS 0.006642f
C246 B.n180 VSUBS 0.006642f
C247 B.n181 VSUBS 0.006642f
C248 B.n182 VSUBS 0.006642f
C249 B.n183 VSUBS 0.006642f
C250 B.n184 VSUBS 0.006642f
C251 B.n185 VSUBS 0.006642f
C252 B.n186 VSUBS 0.006642f
C253 B.n187 VSUBS 0.006642f
C254 B.n188 VSUBS 0.006642f
C255 B.n189 VSUBS 0.006642f
C256 B.n190 VSUBS 0.006642f
C257 B.n191 VSUBS 0.006642f
C258 B.n192 VSUBS 0.006642f
C259 B.n193 VSUBS 0.006642f
C260 B.n194 VSUBS 0.006642f
C261 B.n195 VSUBS 0.006642f
C262 B.n196 VSUBS 0.006642f
C263 B.n197 VSUBS 0.006642f
C264 B.n198 VSUBS 0.006642f
C265 B.n199 VSUBS 0.006642f
C266 B.n200 VSUBS 0.006642f
C267 B.n201 VSUBS 0.006642f
C268 B.n202 VSUBS 0.006642f
C269 B.n203 VSUBS 0.006642f
C270 B.n204 VSUBS 0.006642f
C271 B.n205 VSUBS 0.006642f
C272 B.n206 VSUBS 0.006642f
C273 B.n207 VSUBS 0.006642f
C274 B.n208 VSUBS 0.006642f
C275 B.n209 VSUBS 0.006642f
C276 B.n210 VSUBS 0.006642f
C277 B.n211 VSUBS 0.006642f
C278 B.n212 VSUBS 0.006642f
C279 B.n213 VSUBS 0.006642f
C280 B.n214 VSUBS 0.006642f
C281 B.n215 VSUBS 0.006642f
C282 B.n216 VSUBS 0.006642f
C283 B.n217 VSUBS 0.006642f
C284 B.n218 VSUBS 0.006642f
C285 B.n219 VSUBS 0.006642f
C286 B.n220 VSUBS 0.006642f
C287 B.n221 VSUBS 0.006642f
C288 B.n222 VSUBS 0.006642f
C289 B.n223 VSUBS 0.015296f
C290 B.n224 VSUBS 0.015296f
C291 B.n225 VSUBS 0.01596f
C292 B.n226 VSUBS 0.006642f
C293 B.n227 VSUBS 0.006642f
C294 B.n228 VSUBS 0.006642f
C295 B.n229 VSUBS 0.006642f
C296 B.n230 VSUBS 0.006642f
C297 B.n231 VSUBS 0.006642f
C298 B.n232 VSUBS 0.006642f
C299 B.n233 VSUBS 0.006642f
C300 B.n234 VSUBS 0.006642f
C301 B.n235 VSUBS 0.006642f
C302 B.n236 VSUBS 0.006642f
C303 B.n237 VSUBS 0.006642f
C304 B.n238 VSUBS 0.006642f
C305 B.n239 VSUBS 0.006642f
C306 B.n240 VSUBS 0.006642f
C307 B.n241 VSUBS 0.006642f
C308 B.n242 VSUBS 0.006642f
C309 B.n243 VSUBS 0.006642f
C310 B.n244 VSUBS 0.006642f
C311 B.n245 VSUBS 0.006642f
C312 B.n246 VSUBS 0.006642f
C313 B.n247 VSUBS 0.006642f
C314 B.n248 VSUBS 0.006642f
C315 B.n249 VSUBS 0.006642f
C316 B.n250 VSUBS 0.006642f
C317 B.n251 VSUBS 0.006642f
C318 B.n252 VSUBS 0.006642f
C319 B.n253 VSUBS 0.006642f
C320 B.n254 VSUBS 0.006642f
C321 B.n255 VSUBS 0.006642f
C322 B.n256 VSUBS 0.006642f
C323 B.n257 VSUBS 0.006642f
C324 B.n258 VSUBS 0.006642f
C325 B.n259 VSUBS 0.006642f
C326 B.n260 VSUBS 0.006642f
C327 B.n261 VSUBS 0.006642f
C328 B.n262 VSUBS 0.006642f
C329 B.n263 VSUBS 0.006642f
C330 B.n264 VSUBS 0.006642f
C331 B.n265 VSUBS 0.006642f
C332 B.n266 VSUBS 0.006642f
C333 B.n267 VSUBS 0.006642f
C334 B.n268 VSUBS 0.006642f
C335 B.n269 VSUBS 0.006642f
C336 B.n270 VSUBS 0.006642f
C337 B.n271 VSUBS 0.006642f
C338 B.n272 VSUBS 0.006642f
C339 B.n273 VSUBS 0.006642f
C340 B.n274 VSUBS 0.006642f
C341 B.n275 VSUBS 0.006642f
C342 B.n276 VSUBS 0.006642f
C343 B.n277 VSUBS 0.006642f
C344 B.n278 VSUBS 0.006642f
C345 B.n279 VSUBS 0.006642f
C346 B.n280 VSUBS 0.006642f
C347 B.n281 VSUBS 0.006642f
C348 B.n282 VSUBS 0.006642f
C349 B.n283 VSUBS 0.006642f
C350 B.n284 VSUBS 0.006642f
C351 B.n285 VSUBS 0.004591f
C352 B.n286 VSUBS 0.015388f
C353 B.n287 VSUBS 0.005372f
C354 B.n288 VSUBS 0.006642f
C355 B.n289 VSUBS 0.006642f
C356 B.n290 VSUBS 0.006642f
C357 B.n291 VSUBS 0.006642f
C358 B.n292 VSUBS 0.006642f
C359 B.n293 VSUBS 0.006642f
C360 B.n294 VSUBS 0.006642f
C361 B.n295 VSUBS 0.006642f
C362 B.n296 VSUBS 0.006642f
C363 B.n297 VSUBS 0.006642f
C364 B.n298 VSUBS 0.006642f
C365 B.t4 VSUBS 0.36112f
C366 B.t5 VSUBS 0.382411f
C367 B.t3 VSUBS 1.44239f
C368 B.n299 VSUBS 0.204822f
C369 B.n300 VSUBS 0.069008f
C370 B.n301 VSUBS 0.015388f
C371 B.n302 VSUBS 0.005372f
C372 B.n303 VSUBS 0.006642f
C373 B.n304 VSUBS 0.006642f
C374 B.n305 VSUBS 0.006642f
C375 B.n306 VSUBS 0.006642f
C376 B.n307 VSUBS 0.006642f
C377 B.n308 VSUBS 0.006642f
C378 B.n309 VSUBS 0.006642f
C379 B.n310 VSUBS 0.006642f
C380 B.n311 VSUBS 0.006642f
C381 B.n312 VSUBS 0.006642f
C382 B.n313 VSUBS 0.006642f
C383 B.n314 VSUBS 0.006642f
C384 B.n315 VSUBS 0.006642f
C385 B.n316 VSUBS 0.006642f
C386 B.n317 VSUBS 0.006642f
C387 B.n318 VSUBS 0.006642f
C388 B.n319 VSUBS 0.006642f
C389 B.n320 VSUBS 0.006642f
C390 B.n321 VSUBS 0.006642f
C391 B.n322 VSUBS 0.006642f
C392 B.n323 VSUBS 0.006642f
C393 B.n324 VSUBS 0.006642f
C394 B.n325 VSUBS 0.006642f
C395 B.n326 VSUBS 0.006642f
C396 B.n327 VSUBS 0.006642f
C397 B.n328 VSUBS 0.006642f
C398 B.n329 VSUBS 0.006642f
C399 B.n330 VSUBS 0.006642f
C400 B.n331 VSUBS 0.006642f
C401 B.n332 VSUBS 0.006642f
C402 B.n333 VSUBS 0.006642f
C403 B.n334 VSUBS 0.006642f
C404 B.n335 VSUBS 0.006642f
C405 B.n336 VSUBS 0.006642f
C406 B.n337 VSUBS 0.006642f
C407 B.n338 VSUBS 0.006642f
C408 B.n339 VSUBS 0.006642f
C409 B.n340 VSUBS 0.006642f
C410 B.n341 VSUBS 0.006642f
C411 B.n342 VSUBS 0.006642f
C412 B.n343 VSUBS 0.006642f
C413 B.n344 VSUBS 0.006642f
C414 B.n345 VSUBS 0.006642f
C415 B.n346 VSUBS 0.006642f
C416 B.n347 VSUBS 0.006642f
C417 B.n348 VSUBS 0.006642f
C418 B.n349 VSUBS 0.006642f
C419 B.n350 VSUBS 0.006642f
C420 B.n351 VSUBS 0.006642f
C421 B.n352 VSUBS 0.006642f
C422 B.n353 VSUBS 0.006642f
C423 B.n354 VSUBS 0.006642f
C424 B.n355 VSUBS 0.006642f
C425 B.n356 VSUBS 0.006642f
C426 B.n357 VSUBS 0.006642f
C427 B.n358 VSUBS 0.006642f
C428 B.n359 VSUBS 0.006642f
C429 B.n360 VSUBS 0.006642f
C430 B.n361 VSUBS 0.006642f
C431 B.n362 VSUBS 0.006642f
C432 B.n363 VSUBS 0.006642f
C433 B.n364 VSUBS 0.01596f
C434 B.n365 VSUBS 0.015296f
C435 B.n366 VSUBS 0.015296f
C436 B.n367 VSUBS 0.006642f
C437 B.n368 VSUBS 0.006642f
C438 B.n369 VSUBS 0.006642f
C439 B.n370 VSUBS 0.006642f
C440 B.n371 VSUBS 0.006642f
C441 B.n372 VSUBS 0.006642f
C442 B.n373 VSUBS 0.006642f
C443 B.n374 VSUBS 0.006642f
C444 B.n375 VSUBS 0.006642f
C445 B.n376 VSUBS 0.006642f
C446 B.n377 VSUBS 0.006642f
C447 B.n378 VSUBS 0.006642f
C448 B.n379 VSUBS 0.006642f
C449 B.n380 VSUBS 0.006642f
C450 B.n381 VSUBS 0.006642f
C451 B.n382 VSUBS 0.006642f
C452 B.n383 VSUBS 0.006642f
C453 B.n384 VSUBS 0.006642f
C454 B.n385 VSUBS 0.006642f
C455 B.n386 VSUBS 0.006642f
C456 B.n387 VSUBS 0.006642f
C457 B.n388 VSUBS 0.006642f
C458 B.n389 VSUBS 0.006642f
C459 B.n390 VSUBS 0.006642f
C460 B.n391 VSUBS 0.006642f
C461 B.n392 VSUBS 0.006642f
C462 B.n393 VSUBS 0.006642f
C463 B.n394 VSUBS 0.006642f
C464 B.n395 VSUBS 0.006642f
C465 B.n396 VSUBS 0.006642f
C466 B.n397 VSUBS 0.006642f
C467 B.n398 VSUBS 0.006642f
C468 B.n399 VSUBS 0.006642f
C469 B.n400 VSUBS 0.006642f
C470 B.n401 VSUBS 0.006642f
C471 B.n402 VSUBS 0.006642f
C472 B.n403 VSUBS 0.006642f
C473 B.n404 VSUBS 0.006642f
C474 B.n405 VSUBS 0.006642f
C475 B.n406 VSUBS 0.006642f
C476 B.n407 VSUBS 0.006642f
C477 B.n408 VSUBS 0.006642f
C478 B.n409 VSUBS 0.006642f
C479 B.n410 VSUBS 0.006642f
C480 B.n411 VSUBS 0.006642f
C481 B.n412 VSUBS 0.006642f
C482 B.n413 VSUBS 0.006642f
C483 B.n414 VSUBS 0.006642f
C484 B.n415 VSUBS 0.006642f
C485 B.n416 VSUBS 0.006642f
C486 B.n417 VSUBS 0.006642f
C487 B.n418 VSUBS 0.006642f
C488 B.n419 VSUBS 0.006642f
C489 B.n420 VSUBS 0.006642f
C490 B.n421 VSUBS 0.006642f
C491 B.n422 VSUBS 0.006642f
C492 B.n423 VSUBS 0.006642f
C493 B.n424 VSUBS 0.006642f
C494 B.n425 VSUBS 0.006642f
C495 B.n426 VSUBS 0.006642f
C496 B.n427 VSUBS 0.006642f
C497 B.n428 VSUBS 0.006642f
C498 B.n429 VSUBS 0.006642f
C499 B.n430 VSUBS 0.006642f
C500 B.n431 VSUBS 0.006642f
C501 B.n432 VSUBS 0.006642f
C502 B.n433 VSUBS 0.006642f
C503 B.n434 VSUBS 0.006642f
C504 B.n435 VSUBS 0.006642f
C505 B.n436 VSUBS 0.006642f
C506 B.n437 VSUBS 0.006642f
C507 B.n438 VSUBS 0.006642f
C508 B.n439 VSUBS 0.006642f
C509 B.n440 VSUBS 0.006642f
C510 B.n441 VSUBS 0.006642f
C511 B.n442 VSUBS 0.006642f
C512 B.n443 VSUBS 0.006642f
C513 B.n444 VSUBS 0.006642f
C514 B.n445 VSUBS 0.006642f
C515 B.n446 VSUBS 0.006642f
C516 B.n447 VSUBS 0.006642f
C517 B.n448 VSUBS 0.006642f
C518 B.n449 VSUBS 0.006642f
C519 B.n450 VSUBS 0.006642f
C520 B.n451 VSUBS 0.006642f
C521 B.n452 VSUBS 0.006642f
C522 B.n453 VSUBS 0.006642f
C523 B.n454 VSUBS 0.006642f
C524 B.n455 VSUBS 0.006642f
C525 B.n456 VSUBS 0.006642f
C526 B.n457 VSUBS 0.006642f
C527 B.n458 VSUBS 0.006642f
C528 B.n459 VSUBS 0.006642f
C529 B.n460 VSUBS 0.006642f
C530 B.n461 VSUBS 0.006642f
C531 B.n462 VSUBS 0.006642f
C532 B.n463 VSUBS 0.006642f
C533 B.n464 VSUBS 0.006642f
C534 B.n465 VSUBS 0.006642f
C535 B.n466 VSUBS 0.006642f
C536 B.n467 VSUBS 0.006642f
C537 B.n468 VSUBS 0.006642f
C538 B.n469 VSUBS 0.006642f
C539 B.n470 VSUBS 0.006642f
C540 B.n471 VSUBS 0.006642f
C541 B.n472 VSUBS 0.006642f
C542 B.n473 VSUBS 0.015296f
C543 B.n474 VSUBS 0.016074f
C544 B.n475 VSUBS 0.015182f
C545 B.n476 VSUBS 0.006642f
C546 B.n477 VSUBS 0.006642f
C547 B.n478 VSUBS 0.006642f
C548 B.n479 VSUBS 0.006642f
C549 B.n480 VSUBS 0.006642f
C550 B.n481 VSUBS 0.006642f
C551 B.n482 VSUBS 0.006642f
C552 B.n483 VSUBS 0.006642f
C553 B.n484 VSUBS 0.006642f
C554 B.n485 VSUBS 0.006642f
C555 B.n486 VSUBS 0.006642f
C556 B.n487 VSUBS 0.006642f
C557 B.n488 VSUBS 0.006642f
C558 B.n489 VSUBS 0.006642f
C559 B.n490 VSUBS 0.006642f
C560 B.n491 VSUBS 0.006642f
C561 B.n492 VSUBS 0.006642f
C562 B.n493 VSUBS 0.006642f
C563 B.n494 VSUBS 0.006642f
C564 B.n495 VSUBS 0.006642f
C565 B.n496 VSUBS 0.006642f
C566 B.n497 VSUBS 0.006642f
C567 B.n498 VSUBS 0.006642f
C568 B.n499 VSUBS 0.006642f
C569 B.n500 VSUBS 0.006642f
C570 B.n501 VSUBS 0.006642f
C571 B.n502 VSUBS 0.006642f
C572 B.n503 VSUBS 0.006642f
C573 B.n504 VSUBS 0.006642f
C574 B.n505 VSUBS 0.006642f
C575 B.n506 VSUBS 0.006642f
C576 B.n507 VSUBS 0.006642f
C577 B.n508 VSUBS 0.006642f
C578 B.n509 VSUBS 0.006642f
C579 B.n510 VSUBS 0.006642f
C580 B.n511 VSUBS 0.006642f
C581 B.n512 VSUBS 0.006642f
C582 B.n513 VSUBS 0.006642f
C583 B.n514 VSUBS 0.006642f
C584 B.n515 VSUBS 0.006642f
C585 B.n516 VSUBS 0.006642f
C586 B.n517 VSUBS 0.006642f
C587 B.n518 VSUBS 0.006642f
C588 B.n519 VSUBS 0.006642f
C589 B.n520 VSUBS 0.006642f
C590 B.n521 VSUBS 0.006642f
C591 B.n522 VSUBS 0.006642f
C592 B.n523 VSUBS 0.006642f
C593 B.n524 VSUBS 0.006642f
C594 B.n525 VSUBS 0.006642f
C595 B.n526 VSUBS 0.006642f
C596 B.n527 VSUBS 0.006642f
C597 B.n528 VSUBS 0.006642f
C598 B.n529 VSUBS 0.006642f
C599 B.n530 VSUBS 0.006642f
C600 B.n531 VSUBS 0.006642f
C601 B.n532 VSUBS 0.006642f
C602 B.n533 VSUBS 0.006642f
C603 B.n534 VSUBS 0.006642f
C604 B.n535 VSUBS 0.004591f
C605 B.n536 VSUBS 0.015388f
C606 B.n537 VSUBS 0.005372f
C607 B.n538 VSUBS 0.006642f
C608 B.n539 VSUBS 0.006642f
C609 B.n540 VSUBS 0.006642f
C610 B.n541 VSUBS 0.006642f
C611 B.n542 VSUBS 0.006642f
C612 B.n543 VSUBS 0.006642f
C613 B.n544 VSUBS 0.006642f
C614 B.n545 VSUBS 0.006642f
C615 B.n546 VSUBS 0.006642f
C616 B.n547 VSUBS 0.006642f
C617 B.n548 VSUBS 0.006642f
C618 B.n549 VSUBS 0.005372f
C619 B.n550 VSUBS 0.006642f
C620 B.n551 VSUBS 0.006642f
C621 B.n552 VSUBS 0.006642f
C622 B.n553 VSUBS 0.006642f
C623 B.n554 VSUBS 0.006642f
C624 B.n555 VSUBS 0.006642f
C625 B.n556 VSUBS 0.006642f
C626 B.n557 VSUBS 0.006642f
C627 B.n558 VSUBS 0.006642f
C628 B.n559 VSUBS 0.006642f
C629 B.n560 VSUBS 0.006642f
C630 B.n561 VSUBS 0.006642f
C631 B.n562 VSUBS 0.006642f
C632 B.n563 VSUBS 0.006642f
C633 B.n564 VSUBS 0.006642f
C634 B.n565 VSUBS 0.006642f
C635 B.n566 VSUBS 0.006642f
C636 B.n567 VSUBS 0.006642f
C637 B.n568 VSUBS 0.006642f
C638 B.n569 VSUBS 0.006642f
C639 B.n570 VSUBS 0.006642f
C640 B.n571 VSUBS 0.006642f
C641 B.n572 VSUBS 0.006642f
C642 B.n573 VSUBS 0.006642f
C643 B.n574 VSUBS 0.006642f
C644 B.n575 VSUBS 0.006642f
C645 B.n576 VSUBS 0.006642f
C646 B.n577 VSUBS 0.006642f
C647 B.n578 VSUBS 0.006642f
C648 B.n579 VSUBS 0.006642f
C649 B.n580 VSUBS 0.006642f
C650 B.n581 VSUBS 0.006642f
C651 B.n582 VSUBS 0.006642f
C652 B.n583 VSUBS 0.006642f
C653 B.n584 VSUBS 0.006642f
C654 B.n585 VSUBS 0.006642f
C655 B.n586 VSUBS 0.006642f
C656 B.n587 VSUBS 0.006642f
C657 B.n588 VSUBS 0.006642f
C658 B.n589 VSUBS 0.006642f
C659 B.n590 VSUBS 0.006642f
C660 B.n591 VSUBS 0.006642f
C661 B.n592 VSUBS 0.006642f
C662 B.n593 VSUBS 0.006642f
C663 B.n594 VSUBS 0.006642f
C664 B.n595 VSUBS 0.006642f
C665 B.n596 VSUBS 0.006642f
C666 B.n597 VSUBS 0.006642f
C667 B.n598 VSUBS 0.006642f
C668 B.n599 VSUBS 0.006642f
C669 B.n600 VSUBS 0.006642f
C670 B.n601 VSUBS 0.006642f
C671 B.n602 VSUBS 0.006642f
C672 B.n603 VSUBS 0.006642f
C673 B.n604 VSUBS 0.006642f
C674 B.n605 VSUBS 0.006642f
C675 B.n606 VSUBS 0.006642f
C676 B.n607 VSUBS 0.006642f
C677 B.n608 VSUBS 0.006642f
C678 B.n609 VSUBS 0.006642f
C679 B.n610 VSUBS 0.006642f
C680 B.n611 VSUBS 0.01596f
C681 B.n612 VSUBS 0.015296f
C682 B.n613 VSUBS 0.015296f
C683 B.n614 VSUBS 0.006642f
C684 B.n615 VSUBS 0.006642f
C685 B.n616 VSUBS 0.006642f
C686 B.n617 VSUBS 0.006642f
C687 B.n618 VSUBS 0.006642f
C688 B.n619 VSUBS 0.006642f
C689 B.n620 VSUBS 0.006642f
C690 B.n621 VSUBS 0.006642f
C691 B.n622 VSUBS 0.006642f
C692 B.n623 VSUBS 0.006642f
C693 B.n624 VSUBS 0.006642f
C694 B.n625 VSUBS 0.006642f
C695 B.n626 VSUBS 0.006642f
C696 B.n627 VSUBS 0.006642f
C697 B.n628 VSUBS 0.006642f
C698 B.n629 VSUBS 0.006642f
C699 B.n630 VSUBS 0.006642f
C700 B.n631 VSUBS 0.006642f
C701 B.n632 VSUBS 0.006642f
C702 B.n633 VSUBS 0.006642f
C703 B.n634 VSUBS 0.006642f
C704 B.n635 VSUBS 0.006642f
C705 B.n636 VSUBS 0.006642f
C706 B.n637 VSUBS 0.006642f
C707 B.n638 VSUBS 0.006642f
C708 B.n639 VSUBS 0.006642f
C709 B.n640 VSUBS 0.006642f
C710 B.n641 VSUBS 0.006642f
C711 B.n642 VSUBS 0.006642f
C712 B.n643 VSUBS 0.006642f
C713 B.n644 VSUBS 0.006642f
C714 B.n645 VSUBS 0.006642f
C715 B.n646 VSUBS 0.006642f
C716 B.n647 VSUBS 0.006642f
C717 B.n648 VSUBS 0.006642f
C718 B.n649 VSUBS 0.006642f
C719 B.n650 VSUBS 0.006642f
C720 B.n651 VSUBS 0.006642f
C721 B.n652 VSUBS 0.006642f
C722 B.n653 VSUBS 0.006642f
C723 B.n654 VSUBS 0.006642f
C724 B.n655 VSUBS 0.006642f
C725 B.n656 VSUBS 0.006642f
C726 B.n657 VSUBS 0.006642f
C727 B.n658 VSUBS 0.006642f
C728 B.n659 VSUBS 0.006642f
C729 B.n660 VSUBS 0.006642f
C730 B.n661 VSUBS 0.006642f
C731 B.n662 VSUBS 0.006642f
C732 B.n663 VSUBS 0.006642f
C733 B.n664 VSUBS 0.006642f
C734 B.n665 VSUBS 0.006642f
C735 B.n666 VSUBS 0.006642f
C736 B.n667 VSUBS 0.015039f
C737 VTAIL.t6 VSUBS 2.1053f
C738 VTAIL.n0 VSUBS 0.790312f
C739 VTAIL.t1 VSUBS 2.1053f
C740 VTAIL.n1 VSUBS 0.89122f
C741 VTAIL.t2 VSUBS 2.1053f
C742 VTAIL.n2 VSUBS 2.17317f
C743 VTAIL.t4 VSUBS 2.10531f
C744 VTAIL.n3 VSUBS 2.17317f
C745 VTAIL.t3 VSUBS 2.10531f
C746 VTAIL.n4 VSUBS 0.891213f
C747 VTAIL.t0 VSUBS 2.10531f
C748 VTAIL.n5 VSUBS 0.891213f
C749 VTAIL.t7 VSUBS 2.1053f
C750 VTAIL.n6 VSUBS 2.17317f
C751 VTAIL.t5 VSUBS 2.1053f
C752 VTAIL.n7 VSUBS 2.06326f
C753 VDD2.t1 VSUBS 0.248037f
C754 VDD2.t3 VSUBS 0.248037f
C755 VDD2.n0 VSUBS 2.63374f
C756 VDD2.t2 VSUBS 0.248037f
C757 VDD2.t0 VSUBS 0.248037f
C758 VDD2.n1 VSUBS 1.92329f
C759 VDD2.n2 VSUBS 4.30976f
C760 VN.t0 VSUBS 3.18776f
C761 VN.t1 VSUBS 3.17985f
C762 VN.n0 VSUBS 1.99104f
C763 VN.t3 VSUBS 3.18776f
C764 VN.t2 VSUBS 3.17985f
C765 VN.n1 VSUBS 3.788f
.ends

