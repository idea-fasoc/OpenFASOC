* NGSPICE file created from diff_pair_sample_0391.ext - technology: sky130A

.subckt diff_pair_sample_0391 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=0 ps=0 w=11.8 l=3.01
X1 VTAIL.t15 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=1.947 ps=12.13 w=11.8 l=3.01
X2 VDD2.t7 VN.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=4.602 ps=24.38 w=11.8 l=3.01
X3 VDD1.t6 VP.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=4.602 ps=24.38 w=11.8 l=3.01
X4 VDD2.t6 VN.t1 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
X5 VTAIL.t13 VP.t2 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
X6 VTAIL.t1 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=1.947 ps=12.13 w=11.8 l=3.01
X7 VDD1.t1 VP.t3 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
X8 VTAIL.t3 VN.t3 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=1.947 ps=12.13 w=11.8 l=3.01
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=0 ps=0 w=11.8 l=3.01
X10 VDD1.t0 VP.t4 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
X11 VTAIL.t6 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
X12 VDD1.t7 VP.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=4.602 ps=24.38 w=11.8 l=3.01
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=0 ps=0 w=11.8 l=3.01
X14 VDD2.t2 VN.t5 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=4.602 ps=24.38 w=11.8 l=3.01
X15 VTAIL.t9 VP.t6 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=1.947 ps=12.13 w=11.8 l=3.01
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.602 pd=24.38 as=0 ps=0 w=11.8 l=3.01
X17 VTAIL.t8 VP.t7 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
X18 VDD2.t1 VN.t6 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
X19 VTAIL.t5 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.947 pd=12.13 as=1.947 ps=12.13 w=11.8 l=3.01
R0 B.n929 B.n928 585
R1 B.n337 B.n150 585
R2 B.n336 B.n335 585
R3 B.n334 B.n333 585
R4 B.n332 B.n331 585
R5 B.n330 B.n329 585
R6 B.n328 B.n327 585
R7 B.n326 B.n325 585
R8 B.n324 B.n323 585
R9 B.n322 B.n321 585
R10 B.n320 B.n319 585
R11 B.n318 B.n317 585
R12 B.n316 B.n315 585
R13 B.n314 B.n313 585
R14 B.n312 B.n311 585
R15 B.n310 B.n309 585
R16 B.n308 B.n307 585
R17 B.n306 B.n305 585
R18 B.n304 B.n303 585
R19 B.n302 B.n301 585
R20 B.n300 B.n299 585
R21 B.n298 B.n297 585
R22 B.n296 B.n295 585
R23 B.n294 B.n293 585
R24 B.n292 B.n291 585
R25 B.n290 B.n289 585
R26 B.n288 B.n287 585
R27 B.n286 B.n285 585
R28 B.n284 B.n283 585
R29 B.n282 B.n281 585
R30 B.n280 B.n279 585
R31 B.n278 B.n277 585
R32 B.n276 B.n275 585
R33 B.n274 B.n273 585
R34 B.n272 B.n271 585
R35 B.n270 B.n269 585
R36 B.n268 B.n267 585
R37 B.n266 B.n265 585
R38 B.n264 B.n263 585
R39 B.n262 B.n261 585
R40 B.n260 B.n259 585
R41 B.n257 B.n256 585
R42 B.n255 B.n254 585
R43 B.n253 B.n252 585
R44 B.n251 B.n250 585
R45 B.n249 B.n248 585
R46 B.n247 B.n246 585
R47 B.n245 B.n244 585
R48 B.n243 B.n242 585
R49 B.n241 B.n240 585
R50 B.n239 B.n238 585
R51 B.n236 B.n235 585
R52 B.n234 B.n233 585
R53 B.n232 B.n231 585
R54 B.n230 B.n229 585
R55 B.n228 B.n227 585
R56 B.n226 B.n225 585
R57 B.n224 B.n223 585
R58 B.n222 B.n221 585
R59 B.n220 B.n219 585
R60 B.n218 B.n217 585
R61 B.n216 B.n215 585
R62 B.n214 B.n213 585
R63 B.n212 B.n211 585
R64 B.n210 B.n209 585
R65 B.n208 B.n207 585
R66 B.n206 B.n205 585
R67 B.n204 B.n203 585
R68 B.n202 B.n201 585
R69 B.n200 B.n199 585
R70 B.n198 B.n197 585
R71 B.n196 B.n195 585
R72 B.n194 B.n193 585
R73 B.n192 B.n191 585
R74 B.n190 B.n189 585
R75 B.n188 B.n187 585
R76 B.n186 B.n185 585
R77 B.n184 B.n183 585
R78 B.n182 B.n181 585
R79 B.n180 B.n179 585
R80 B.n178 B.n177 585
R81 B.n176 B.n175 585
R82 B.n174 B.n173 585
R83 B.n172 B.n171 585
R84 B.n170 B.n169 585
R85 B.n168 B.n167 585
R86 B.n166 B.n165 585
R87 B.n164 B.n163 585
R88 B.n162 B.n161 585
R89 B.n160 B.n159 585
R90 B.n158 B.n157 585
R91 B.n156 B.n155 585
R92 B.n927 B.n104 585
R93 B.n932 B.n104 585
R94 B.n926 B.n103 585
R95 B.n933 B.n103 585
R96 B.n925 B.n924 585
R97 B.n924 B.n99 585
R98 B.n923 B.n98 585
R99 B.n939 B.n98 585
R100 B.n922 B.n97 585
R101 B.n940 B.n97 585
R102 B.n921 B.n96 585
R103 B.n941 B.n96 585
R104 B.n920 B.n919 585
R105 B.n919 B.n92 585
R106 B.n918 B.n91 585
R107 B.n947 B.n91 585
R108 B.n917 B.n90 585
R109 B.n948 B.n90 585
R110 B.n916 B.n89 585
R111 B.n949 B.n89 585
R112 B.n915 B.n914 585
R113 B.n914 B.n85 585
R114 B.n913 B.n84 585
R115 B.n955 B.n84 585
R116 B.n912 B.n83 585
R117 B.n956 B.n83 585
R118 B.n911 B.n82 585
R119 B.n957 B.n82 585
R120 B.n910 B.n909 585
R121 B.n909 B.n78 585
R122 B.n908 B.n77 585
R123 B.n963 B.n77 585
R124 B.n907 B.n76 585
R125 B.n964 B.n76 585
R126 B.n906 B.n75 585
R127 B.n965 B.n75 585
R128 B.n905 B.n904 585
R129 B.n904 B.n71 585
R130 B.n903 B.n70 585
R131 B.n971 B.n70 585
R132 B.n902 B.n69 585
R133 B.n972 B.n69 585
R134 B.n901 B.n68 585
R135 B.n973 B.n68 585
R136 B.n900 B.n899 585
R137 B.n899 B.n64 585
R138 B.n898 B.n63 585
R139 B.n979 B.n63 585
R140 B.n897 B.n62 585
R141 B.n980 B.n62 585
R142 B.n896 B.n61 585
R143 B.n981 B.n61 585
R144 B.n895 B.n894 585
R145 B.n894 B.n57 585
R146 B.n893 B.n56 585
R147 B.n987 B.n56 585
R148 B.n892 B.n55 585
R149 B.n988 B.n55 585
R150 B.n891 B.n54 585
R151 B.n989 B.n54 585
R152 B.n890 B.n889 585
R153 B.n889 B.n53 585
R154 B.n888 B.n49 585
R155 B.n995 B.n49 585
R156 B.n887 B.n48 585
R157 B.n996 B.n48 585
R158 B.n886 B.n47 585
R159 B.n997 B.n47 585
R160 B.n885 B.n884 585
R161 B.n884 B.n43 585
R162 B.n883 B.n42 585
R163 B.n1003 B.n42 585
R164 B.n882 B.n41 585
R165 B.n1004 B.n41 585
R166 B.n881 B.n40 585
R167 B.n1005 B.n40 585
R168 B.n880 B.n879 585
R169 B.n879 B.n36 585
R170 B.n878 B.n35 585
R171 B.n1011 B.n35 585
R172 B.n877 B.n34 585
R173 B.n1012 B.n34 585
R174 B.n876 B.n33 585
R175 B.n1013 B.n33 585
R176 B.n875 B.n874 585
R177 B.n874 B.n29 585
R178 B.n873 B.n28 585
R179 B.n1019 B.n28 585
R180 B.n872 B.n27 585
R181 B.n1020 B.n27 585
R182 B.n871 B.n26 585
R183 B.n1021 B.n26 585
R184 B.n870 B.n869 585
R185 B.n869 B.n22 585
R186 B.n868 B.n21 585
R187 B.n1027 B.n21 585
R188 B.n867 B.n20 585
R189 B.n1028 B.n20 585
R190 B.n866 B.n19 585
R191 B.n1029 B.n19 585
R192 B.n865 B.n864 585
R193 B.n864 B.n18 585
R194 B.n863 B.n14 585
R195 B.n1035 B.n14 585
R196 B.n862 B.n13 585
R197 B.n1036 B.n13 585
R198 B.n861 B.n12 585
R199 B.n1037 B.n12 585
R200 B.n860 B.n859 585
R201 B.n859 B.n8 585
R202 B.n858 B.n7 585
R203 B.n1043 B.n7 585
R204 B.n857 B.n6 585
R205 B.n1044 B.n6 585
R206 B.n856 B.n5 585
R207 B.n1045 B.n5 585
R208 B.n855 B.n854 585
R209 B.n854 B.n4 585
R210 B.n853 B.n338 585
R211 B.n853 B.n852 585
R212 B.n843 B.n339 585
R213 B.n340 B.n339 585
R214 B.n845 B.n844 585
R215 B.n846 B.n845 585
R216 B.n842 B.n345 585
R217 B.n345 B.n344 585
R218 B.n841 B.n840 585
R219 B.n840 B.n839 585
R220 B.n347 B.n346 585
R221 B.n832 B.n347 585
R222 B.n831 B.n830 585
R223 B.n833 B.n831 585
R224 B.n829 B.n352 585
R225 B.n352 B.n351 585
R226 B.n828 B.n827 585
R227 B.n827 B.n826 585
R228 B.n354 B.n353 585
R229 B.n355 B.n354 585
R230 B.n819 B.n818 585
R231 B.n820 B.n819 585
R232 B.n817 B.n360 585
R233 B.n360 B.n359 585
R234 B.n816 B.n815 585
R235 B.n815 B.n814 585
R236 B.n362 B.n361 585
R237 B.n363 B.n362 585
R238 B.n807 B.n806 585
R239 B.n808 B.n807 585
R240 B.n805 B.n367 585
R241 B.n371 B.n367 585
R242 B.n804 B.n803 585
R243 B.n803 B.n802 585
R244 B.n369 B.n368 585
R245 B.n370 B.n369 585
R246 B.n795 B.n794 585
R247 B.n796 B.n795 585
R248 B.n793 B.n376 585
R249 B.n376 B.n375 585
R250 B.n792 B.n791 585
R251 B.n791 B.n790 585
R252 B.n378 B.n377 585
R253 B.n379 B.n378 585
R254 B.n783 B.n782 585
R255 B.n784 B.n783 585
R256 B.n781 B.n384 585
R257 B.n384 B.n383 585
R258 B.n780 B.n779 585
R259 B.n779 B.n778 585
R260 B.n386 B.n385 585
R261 B.n771 B.n386 585
R262 B.n770 B.n769 585
R263 B.n772 B.n770 585
R264 B.n768 B.n391 585
R265 B.n391 B.n390 585
R266 B.n767 B.n766 585
R267 B.n766 B.n765 585
R268 B.n393 B.n392 585
R269 B.n394 B.n393 585
R270 B.n758 B.n757 585
R271 B.n759 B.n758 585
R272 B.n756 B.n399 585
R273 B.n399 B.n398 585
R274 B.n755 B.n754 585
R275 B.n754 B.n753 585
R276 B.n401 B.n400 585
R277 B.n402 B.n401 585
R278 B.n746 B.n745 585
R279 B.n747 B.n746 585
R280 B.n744 B.n407 585
R281 B.n407 B.n406 585
R282 B.n743 B.n742 585
R283 B.n742 B.n741 585
R284 B.n409 B.n408 585
R285 B.n410 B.n409 585
R286 B.n734 B.n733 585
R287 B.n735 B.n734 585
R288 B.n732 B.n415 585
R289 B.n415 B.n414 585
R290 B.n731 B.n730 585
R291 B.n730 B.n729 585
R292 B.n417 B.n416 585
R293 B.n418 B.n417 585
R294 B.n722 B.n721 585
R295 B.n723 B.n722 585
R296 B.n720 B.n423 585
R297 B.n423 B.n422 585
R298 B.n719 B.n718 585
R299 B.n718 B.n717 585
R300 B.n425 B.n424 585
R301 B.n426 B.n425 585
R302 B.n710 B.n709 585
R303 B.n711 B.n710 585
R304 B.n708 B.n431 585
R305 B.n431 B.n430 585
R306 B.n707 B.n706 585
R307 B.n706 B.n705 585
R308 B.n433 B.n432 585
R309 B.n434 B.n433 585
R310 B.n698 B.n697 585
R311 B.n699 B.n698 585
R312 B.n696 B.n439 585
R313 B.n439 B.n438 585
R314 B.n695 B.n694 585
R315 B.n694 B.n693 585
R316 B.n441 B.n440 585
R317 B.n442 B.n441 585
R318 B.n686 B.n685 585
R319 B.n687 B.n686 585
R320 B.n684 B.n447 585
R321 B.n447 B.n446 585
R322 B.n679 B.n678 585
R323 B.n677 B.n495 585
R324 B.n676 B.n494 585
R325 B.n681 B.n494 585
R326 B.n675 B.n674 585
R327 B.n673 B.n672 585
R328 B.n671 B.n670 585
R329 B.n669 B.n668 585
R330 B.n667 B.n666 585
R331 B.n665 B.n664 585
R332 B.n663 B.n662 585
R333 B.n661 B.n660 585
R334 B.n659 B.n658 585
R335 B.n657 B.n656 585
R336 B.n655 B.n654 585
R337 B.n653 B.n652 585
R338 B.n651 B.n650 585
R339 B.n649 B.n648 585
R340 B.n647 B.n646 585
R341 B.n645 B.n644 585
R342 B.n643 B.n642 585
R343 B.n641 B.n640 585
R344 B.n639 B.n638 585
R345 B.n637 B.n636 585
R346 B.n635 B.n634 585
R347 B.n633 B.n632 585
R348 B.n631 B.n630 585
R349 B.n629 B.n628 585
R350 B.n627 B.n626 585
R351 B.n625 B.n624 585
R352 B.n623 B.n622 585
R353 B.n621 B.n620 585
R354 B.n619 B.n618 585
R355 B.n617 B.n616 585
R356 B.n615 B.n614 585
R357 B.n613 B.n612 585
R358 B.n611 B.n610 585
R359 B.n609 B.n608 585
R360 B.n607 B.n606 585
R361 B.n605 B.n604 585
R362 B.n603 B.n602 585
R363 B.n601 B.n600 585
R364 B.n599 B.n598 585
R365 B.n597 B.n596 585
R366 B.n595 B.n594 585
R367 B.n593 B.n592 585
R368 B.n591 B.n590 585
R369 B.n589 B.n588 585
R370 B.n587 B.n586 585
R371 B.n585 B.n584 585
R372 B.n583 B.n582 585
R373 B.n581 B.n580 585
R374 B.n579 B.n578 585
R375 B.n577 B.n576 585
R376 B.n575 B.n574 585
R377 B.n573 B.n572 585
R378 B.n571 B.n570 585
R379 B.n569 B.n568 585
R380 B.n567 B.n566 585
R381 B.n565 B.n564 585
R382 B.n563 B.n562 585
R383 B.n561 B.n560 585
R384 B.n559 B.n558 585
R385 B.n557 B.n556 585
R386 B.n555 B.n554 585
R387 B.n553 B.n552 585
R388 B.n551 B.n550 585
R389 B.n549 B.n548 585
R390 B.n547 B.n546 585
R391 B.n545 B.n544 585
R392 B.n543 B.n542 585
R393 B.n541 B.n540 585
R394 B.n539 B.n538 585
R395 B.n537 B.n536 585
R396 B.n535 B.n534 585
R397 B.n533 B.n532 585
R398 B.n531 B.n530 585
R399 B.n529 B.n528 585
R400 B.n527 B.n526 585
R401 B.n525 B.n524 585
R402 B.n523 B.n522 585
R403 B.n521 B.n520 585
R404 B.n519 B.n518 585
R405 B.n517 B.n516 585
R406 B.n515 B.n514 585
R407 B.n513 B.n512 585
R408 B.n511 B.n510 585
R409 B.n509 B.n508 585
R410 B.n507 B.n506 585
R411 B.n505 B.n504 585
R412 B.n503 B.n502 585
R413 B.n449 B.n448 585
R414 B.n683 B.n682 585
R415 B.n682 B.n681 585
R416 B.n445 B.n444 585
R417 B.n446 B.n445 585
R418 B.n689 B.n688 585
R419 B.n688 B.n687 585
R420 B.n690 B.n443 585
R421 B.n443 B.n442 585
R422 B.n692 B.n691 585
R423 B.n693 B.n692 585
R424 B.n437 B.n436 585
R425 B.n438 B.n437 585
R426 B.n701 B.n700 585
R427 B.n700 B.n699 585
R428 B.n702 B.n435 585
R429 B.n435 B.n434 585
R430 B.n704 B.n703 585
R431 B.n705 B.n704 585
R432 B.n429 B.n428 585
R433 B.n430 B.n429 585
R434 B.n713 B.n712 585
R435 B.n712 B.n711 585
R436 B.n714 B.n427 585
R437 B.n427 B.n426 585
R438 B.n716 B.n715 585
R439 B.n717 B.n716 585
R440 B.n421 B.n420 585
R441 B.n422 B.n421 585
R442 B.n725 B.n724 585
R443 B.n724 B.n723 585
R444 B.n726 B.n419 585
R445 B.n419 B.n418 585
R446 B.n728 B.n727 585
R447 B.n729 B.n728 585
R448 B.n413 B.n412 585
R449 B.n414 B.n413 585
R450 B.n737 B.n736 585
R451 B.n736 B.n735 585
R452 B.n738 B.n411 585
R453 B.n411 B.n410 585
R454 B.n740 B.n739 585
R455 B.n741 B.n740 585
R456 B.n405 B.n404 585
R457 B.n406 B.n405 585
R458 B.n749 B.n748 585
R459 B.n748 B.n747 585
R460 B.n750 B.n403 585
R461 B.n403 B.n402 585
R462 B.n752 B.n751 585
R463 B.n753 B.n752 585
R464 B.n397 B.n396 585
R465 B.n398 B.n397 585
R466 B.n761 B.n760 585
R467 B.n760 B.n759 585
R468 B.n762 B.n395 585
R469 B.n395 B.n394 585
R470 B.n764 B.n763 585
R471 B.n765 B.n764 585
R472 B.n389 B.n388 585
R473 B.n390 B.n389 585
R474 B.n774 B.n773 585
R475 B.n773 B.n772 585
R476 B.n775 B.n387 585
R477 B.n771 B.n387 585
R478 B.n777 B.n776 585
R479 B.n778 B.n777 585
R480 B.n382 B.n381 585
R481 B.n383 B.n382 585
R482 B.n786 B.n785 585
R483 B.n785 B.n784 585
R484 B.n787 B.n380 585
R485 B.n380 B.n379 585
R486 B.n789 B.n788 585
R487 B.n790 B.n789 585
R488 B.n374 B.n373 585
R489 B.n375 B.n374 585
R490 B.n798 B.n797 585
R491 B.n797 B.n796 585
R492 B.n799 B.n372 585
R493 B.n372 B.n370 585
R494 B.n801 B.n800 585
R495 B.n802 B.n801 585
R496 B.n366 B.n365 585
R497 B.n371 B.n366 585
R498 B.n810 B.n809 585
R499 B.n809 B.n808 585
R500 B.n811 B.n364 585
R501 B.n364 B.n363 585
R502 B.n813 B.n812 585
R503 B.n814 B.n813 585
R504 B.n358 B.n357 585
R505 B.n359 B.n358 585
R506 B.n822 B.n821 585
R507 B.n821 B.n820 585
R508 B.n823 B.n356 585
R509 B.n356 B.n355 585
R510 B.n825 B.n824 585
R511 B.n826 B.n825 585
R512 B.n350 B.n349 585
R513 B.n351 B.n350 585
R514 B.n835 B.n834 585
R515 B.n834 B.n833 585
R516 B.n836 B.n348 585
R517 B.n832 B.n348 585
R518 B.n838 B.n837 585
R519 B.n839 B.n838 585
R520 B.n343 B.n342 585
R521 B.n344 B.n343 585
R522 B.n848 B.n847 585
R523 B.n847 B.n846 585
R524 B.n849 B.n341 585
R525 B.n341 B.n340 585
R526 B.n851 B.n850 585
R527 B.n852 B.n851 585
R528 B.n2 B.n0 585
R529 B.n4 B.n2 585
R530 B.n3 B.n1 585
R531 B.n1044 B.n3 585
R532 B.n1042 B.n1041 585
R533 B.n1043 B.n1042 585
R534 B.n1040 B.n9 585
R535 B.n9 B.n8 585
R536 B.n1039 B.n1038 585
R537 B.n1038 B.n1037 585
R538 B.n11 B.n10 585
R539 B.n1036 B.n11 585
R540 B.n1034 B.n1033 585
R541 B.n1035 B.n1034 585
R542 B.n1032 B.n15 585
R543 B.n18 B.n15 585
R544 B.n1031 B.n1030 585
R545 B.n1030 B.n1029 585
R546 B.n17 B.n16 585
R547 B.n1028 B.n17 585
R548 B.n1026 B.n1025 585
R549 B.n1027 B.n1026 585
R550 B.n1024 B.n23 585
R551 B.n23 B.n22 585
R552 B.n1023 B.n1022 585
R553 B.n1022 B.n1021 585
R554 B.n25 B.n24 585
R555 B.n1020 B.n25 585
R556 B.n1018 B.n1017 585
R557 B.n1019 B.n1018 585
R558 B.n1016 B.n30 585
R559 B.n30 B.n29 585
R560 B.n1015 B.n1014 585
R561 B.n1014 B.n1013 585
R562 B.n32 B.n31 585
R563 B.n1012 B.n32 585
R564 B.n1010 B.n1009 585
R565 B.n1011 B.n1010 585
R566 B.n1008 B.n37 585
R567 B.n37 B.n36 585
R568 B.n1007 B.n1006 585
R569 B.n1006 B.n1005 585
R570 B.n39 B.n38 585
R571 B.n1004 B.n39 585
R572 B.n1002 B.n1001 585
R573 B.n1003 B.n1002 585
R574 B.n1000 B.n44 585
R575 B.n44 B.n43 585
R576 B.n999 B.n998 585
R577 B.n998 B.n997 585
R578 B.n46 B.n45 585
R579 B.n996 B.n46 585
R580 B.n994 B.n993 585
R581 B.n995 B.n994 585
R582 B.n992 B.n50 585
R583 B.n53 B.n50 585
R584 B.n991 B.n990 585
R585 B.n990 B.n989 585
R586 B.n52 B.n51 585
R587 B.n988 B.n52 585
R588 B.n986 B.n985 585
R589 B.n987 B.n986 585
R590 B.n984 B.n58 585
R591 B.n58 B.n57 585
R592 B.n983 B.n982 585
R593 B.n982 B.n981 585
R594 B.n60 B.n59 585
R595 B.n980 B.n60 585
R596 B.n978 B.n977 585
R597 B.n979 B.n978 585
R598 B.n976 B.n65 585
R599 B.n65 B.n64 585
R600 B.n975 B.n974 585
R601 B.n974 B.n973 585
R602 B.n67 B.n66 585
R603 B.n972 B.n67 585
R604 B.n970 B.n969 585
R605 B.n971 B.n970 585
R606 B.n968 B.n72 585
R607 B.n72 B.n71 585
R608 B.n967 B.n966 585
R609 B.n966 B.n965 585
R610 B.n74 B.n73 585
R611 B.n964 B.n74 585
R612 B.n962 B.n961 585
R613 B.n963 B.n962 585
R614 B.n960 B.n79 585
R615 B.n79 B.n78 585
R616 B.n959 B.n958 585
R617 B.n958 B.n957 585
R618 B.n81 B.n80 585
R619 B.n956 B.n81 585
R620 B.n954 B.n953 585
R621 B.n955 B.n954 585
R622 B.n952 B.n86 585
R623 B.n86 B.n85 585
R624 B.n951 B.n950 585
R625 B.n950 B.n949 585
R626 B.n88 B.n87 585
R627 B.n948 B.n88 585
R628 B.n946 B.n945 585
R629 B.n947 B.n946 585
R630 B.n944 B.n93 585
R631 B.n93 B.n92 585
R632 B.n943 B.n942 585
R633 B.n942 B.n941 585
R634 B.n95 B.n94 585
R635 B.n940 B.n95 585
R636 B.n938 B.n937 585
R637 B.n939 B.n938 585
R638 B.n936 B.n100 585
R639 B.n100 B.n99 585
R640 B.n935 B.n934 585
R641 B.n934 B.n933 585
R642 B.n102 B.n101 585
R643 B.n932 B.n102 585
R644 B.n1047 B.n1046 585
R645 B.n1046 B.n1045 585
R646 B.n679 B.n445 506.916
R647 B.n155 B.n102 506.916
R648 B.n682 B.n447 506.916
R649 B.n929 B.n104 506.916
R650 B.n499 B.t16 303.07
R651 B.n496 B.t8 303.07
R652 B.n153 B.t19 303.07
R653 B.n151 B.t12 303.07
R654 B.n931 B.n930 256.663
R655 B.n931 B.n149 256.663
R656 B.n931 B.n148 256.663
R657 B.n931 B.n147 256.663
R658 B.n931 B.n146 256.663
R659 B.n931 B.n145 256.663
R660 B.n931 B.n144 256.663
R661 B.n931 B.n143 256.663
R662 B.n931 B.n142 256.663
R663 B.n931 B.n141 256.663
R664 B.n931 B.n140 256.663
R665 B.n931 B.n139 256.663
R666 B.n931 B.n138 256.663
R667 B.n931 B.n137 256.663
R668 B.n931 B.n136 256.663
R669 B.n931 B.n135 256.663
R670 B.n931 B.n134 256.663
R671 B.n931 B.n133 256.663
R672 B.n931 B.n132 256.663
R673 B.n931 B.n131 256.663
R674 B.n931 B.n130 256.663
R675 B.n931 B.n129 256.663
R676 B.n931 B.n128 256.663
R677 B.n931 B.n127 256.663
R678 B.n931 B.n126 256.663
R679 B.n931 B.n125 256.663
R680 B.n931 B.n124 256.663
R681 B.n931 B.n123 256.663
R682 B.n931 B.n122 256.663
R683 B.n931 B.n121 256.663
R684 B.n931 B.n120 256.663
R685 B.n931 B.n119 256.663
R686 B.n931 B.n118 256.663
R687 B.n931 B.n117 256.663
R688 B.n931 B.n116 256.663
R689 B.n931 B.n115 256.663
R690 B.n931 B.n114 256.663
R691 B.n931 B.n113 256.663
R692 B.n931 B.n112 256.663
R693 B.n931 B.n111 256.663
R694 B.n931 B.n110 256.663
R695 B.n931 B.n109 256.663
R696 B.n931 B.n108 256.663
R697 B.n931 B.n107 256.663
R698 B.n931 B.n106 256.663
R699 B.n931 B.n105 256.663
R700 B.n681 B.n680 256.663
R701 B.n681 B.n450 256.663
R702 B.n681 B.n451 256.663
R703 B.n681 B.n452 256.663
R704 B.n681 B.n453 256.663
R705 B.n681 B.n454 256.663
R706 B.n681 B.n455 256.663
R707 B.n681 B.n456 256.663
R708 B.n681 B.n457 256.663
R709 B.n681 B.n458 256.663
R710 B.n681 B.n459 256.663
R711 B.n681 B.n460 256.663
R712 B.n681 B.n461 256.663
R713 B.n681 B.n462 256.663
R714 B.n681 B.n463 256.663
R715 B.n681 B.n464 256.663
R716 B.n681 B.n465 256.663
R717 B.n681 B.n466 256.663
R718 B.n681 B.n467 256.663
R719 B.n681 B.n468 256.663
R720 B.n681 B.n469 256.663
R721 B.n681 B.n470 256.663
R722 B.n681 B.n471 256.663
R723 B.n681 B.n472 256.663
R724 B.n681 B.n473 256.663
R725 B.n681 B.n474 256.663
R726 B.n681 B.n475 256.663
R727 B.n681 B.n476 256.663
R728 B.n681 B.n477 256.663
R729 B.n681 B.n478 256.663
R730 B.n681 B.n479 256.663
R731 B.n681 B.n480 256.663
R732 B.n681 B.n481 256.663
R733 B.n681 B.n482 256.663
R734 B.n681 B.n483 256.663
R735 B.n681 B.n484 256.663
R736 B.n681 B.n485 256.663
R737 B.n681 B.n486 256.663
R738 B.n681 B.n487 256.663
R739 B.n681 B.n488 256.663
R740 B.n681 B.n489 256.663
R741 B.n681 B.n490 256.663
R742 B.n681 B.n491 256.663
R743 B.n681 B.n492 256.663
R744 B.n681 B.n493 256.663
R745 B.n688 B.n445 163.367
R746 B.n688 B.n443 163.367
R747 B.n692 B.n443 163.367
R748 B.n692 B.n437 163.367
R749 B.n700 B.n437 163.367
R750 B.n700 B.n435 163.367
R751 B.n704 B.n435 163.367
R752 B.n704 B.n429 163.367
R753 B.n712 B.n429 163.367
R754 B.n712 B.n427 163.367
R755 B.n716 B.n427 163.367
R756 B.n716 B.n421 163.367
R757 B.n724 B.n421 163.367
R758 B.n724 B.n419 163.367
R759 B.n728 B.n419 163.367
R760 B.n728 B.n413 163.367
R761 B.n736 B.n413 163.367
R762 B.n736 B.n411 163.367
R763 B.n740 B.n411 163.367
R764 B.n740 B.n405 163.367
R765 B.n748 B.n405 163.367
R766 B.n748 B.n403 163.367
R767 B.n752 B.n403 163.367
R768 B.n752 B.n397 163.367
R769 B.n760 B.n397 163.367
R770 B.n760 B.n395 163.367
R771 B.n764 B.n395 163.367
R772 B.n764 B.n389 163.367
R773 B.n773 B.n389 163.367
R774 B.n773 B.n387 163.367
R775 B.n777 B.n387 163.367
R776 B.n777 B.n382 163.367
R777 B.n785 B.n382 163.367
R778 B.n785 B.n380 163.367
R779 B.n789 B.n380 163.367
R780 B.n789 B.n374 163.367
R781 B.n797 B.n374 163.367
R782 B.n797 B.n372 163.367
R783 B.n801 B.n372 163.367
R784 B.n801 B.n366 163.367
R785 B.n809 B.n366 163.367
R786 B.n809 B.n364 163.367
R787 B.n813 B.n364 163.367
R788 B.n813 B.n358 163.367
R789 B.n821 B.n358 163.367
R790 B.n821 B.n356 163.367
R791 B.n825 B.n356 163.367
R792 B.n825 B.n350 163.367
R793 B.n834 B.n350 163.367
R794 B.n834 B.n348 163.367
R795 B.n838 B.n348 163.367
R796 B.n838 B.n343 163.367
R797 B.n847 B.n343 163.367
R798 B.n847 B.n341 163.367
R799 B.n851 B.n341 163.367
R800 B.n851 B.n2 163.367
R801 B.n1046 B.n2 163.367
R802 B.n1046 B.n3 163.367
R803 B.n1042 B.n3 163.367
R804 B.n1042 B.n9 163.367
R805 B.n1038 B.n9 163.367
R806 B.n1038 B.n11 163.367
R807 B.n1034 B.n11 163.367
R808 B.n1034 B.n15 163.367
R809 B.n1030 B.n15 163.367
R810 B.n1030 B.n17 163.367
R811 B.n1026 B.n17 163.367
R812 B.n1026 B.n23 163.367
R813 B.n1022 B.n23 163.367
R814 B.n1022 B.n25 163.367
R815 B.n1018 B.n25 163.367
R816 B.n1018 B.n30 163.367
R817 B.n1014 B.n30 163.367
R818 B.n1014 B.n32 163.367
R819 B.n1010 B.n32 163.367
R820 B.n1010 B.n37 163.367
R821 B.n1006 B.n37 163.367
R822 B.n1006 B.n39 163.367
R823 B.n1002 B.n39 163.367
R824 B.n1002 B.n44 163.367
R825 B.n998 B.n44 163.367
R826 B.n998 B.n46 163.367
R827 B.n994 B.n46 163.367
R828 B.n994 B.n50 163.367
R829 B.n990 B.n50 163.367
R830 B.n990 B.n52 163.367
R831 B.n986 B.n52 163.367
R832 B.n986 B.n58 163.367
R833 B.n982 B.n58 163.367
R834 B.n982 B.n60 163.367
R835 B.n978 B.n60 163.367
R836 B.n978 B.n65 163.367
R837 B.n974 B.n65 163.367
R838 B.n974 B.n67 163.367
R839 B.n970 B.n67 163.367
R840 B.n970 B.n72 163.367
R841 B.n966 B.n72 163.367
R842 B.n966 B.n74 163.367
R843 B.n962 B.n74 163.367
R844 B.n962 B.n79 163.367
R845 B.n958 B.n79 163.367
R846 B.n958 B.n81 163.367
R847 B.n954 B.n81 163.367
R848 B.n954 B.n86 163.367
R849 B.n950 B.n86 163.367
R850 B.n950 B.n88 163.367
R851 B.n946 B.n88 163.367
R852 B.n946 B.n93 163.367
R853 B.n942 B.n93 163.367
R854 B.n942 B.n95 163.367
R855 B.n938 B.n95 163.367
R856 B.n938 B.n100 163.367
R857 B.n934 B.n100 163.367
R858 B.n934 B.n102 163.367
R859 B.n495 B.n494 163.367
R860 B.n674 B.n494 163.367
R861 B.n672 B.n671 163.367
R862 B.n668 B.n667 163.367
R863 B.n664 B.n663 163.367
R864 B.n660 B.n659 163.367
R865 B.n656 B.n655 163.367
R866 B.n652 B.n651 163.367
R867 B.n648 B.n647 163.367
R868 B.n644 B.n643 163.367
R869 B.n640 B.n639 163.367
R870 B.n636 B.n635 163.367
R871 B.n632 B.n631 163.367
R872 B.n628 B.n627 163.367
R873 B.n624 B.n623 163.367
R874 B.n620 B.n619 163.367
R875 B.n616 B.n615 163.367
R876 B.n612 B.n611 163.367
R877 B.n608 B.n607 163.367
R878 B.n604 B.n603 163.367
R879 B.n600 B.n599 163.367
R880 B.n596 B.n595 163.367
R881 B.n592 B.n591 163.367
R882 B.n588 B.n587 163.367
R883 B.n584 B.n583 163.367
R884 B.n580 B.n579 163.367
R885 B.n576 B.n575 163.367
R886 B.n572 B.n571 163.367
R887 B.n568 B.n567 163.367
R888 B.n564 B.n563 163.367
R889 B.n560 B.n559 163.367
R890 B.n556 B.n555 163.367
R891 B.n552 B.n551 163.367
R892 B.n548 B.n547 163.367
R893 B.n544 B.n543 163.367
R894 B.n540 B.n539 163.367
R895 B.n536 B.n535 163.367
R896 B.n532 B.n531 163.367
R897 B.n528 B.n527 163.367
R898 B.n524 B.n523 163.367
R899 B.n520 B.n519 163.367
R900 B.n516 B.n515 163.367
R901 B.n512 B.n511 163.367
R902 B.n508 B.n507 163.367
R903 B.n504 B.n503 163.367
R904 B.n682 B.n449 163.367
R905 B.n686 B.n447 163.367
R906 B.n686 B.n441 163.367
R907 B.n694 B.n441 163.367
R908 B.n694 B.n439 163.367
R909 B.n698 B.n439 163.367
R910 B.n698 B.n433 163.367
R911 B.n706 B.n433 163.367
R912 B.n706 B.n431 163.367
R913 B.n710 B.n431 163.367
R914 B.n710 B.n425 163.367
R915 B.n718 B.n425 163.367
R916 B.n718 B.n423 163.367
R917 B.n722 B.n423 163.367
R918 B.n722 B.n417 163.367
R919 B.n730 B.n417 163.367
R920 B.n730 B.n415 163.367
R921 B.n734 B.n415 163.367
R922 B.n734 B.n409 163.367
R923 B.n742 B.n409 163.367
R924 B.n742 B.n407 163.367
R925 B.n746 B.n407 163.367
R926 B.n746 B.n401 163.367
R927 B.n754 B.n401 163.367
R928 B.n754 B.n399 163.367
R929 B.n758 B.n399 163.367
R930 B.n758 B.n393 163.367
R931 B.n766 B.n393 163.367
R932 B.n766 B.n391 163.367
R933 B.n770 B.n391 163.367
R934 B.n770 B.n386 163.367
R935 B.n779 B.n386 163.367
R936 B.n779 B.n384 163.367
R937 B.n783 B.n384 163.367
R938 B.n783 B.n378 163.367
R939 B.n791 B.n378 163.367
R940 B.n791 B.n376 163.367
R941 B.n795 B.n376 163.367
R942 B.n795 B.n369 163.367
R943 B.n803 B.n369 163.367
R944 B.n803 B.n367 163.367
R945 B.n807 B.n367 163.367
R946 B.n807 B.n362 163.367
R947 B.n815 B.n362 163.367
R948 B.n815 B.n360 163.367
R949 B.n819 B.n360 163.367
R950 B.n819 B.n354 163.367
R951 B.n827 B.n354 163.367
R952 B.n827 B.n352 163.367
R953 B.n831 B.n352 163.367
R954 B.n831 B.n347 163.367
R955 B.n840 B.n347 163.367
R956 B.n840 B.n345 163.367
R957 B.n845 B.n345 163.367
R958 B.n845 B.n339 163.367
R959 B.n853 B.n339 163.367
R960 B.n854 B.n853 163.367
R961 B.n854 B.n5 163.367
R962 B.n6 B.n5 163.367
R963 B.n7 B.n6 163.367
R964 B.n859 B.n7 163.367
R965 B.n859 B.n12 163.367
R966 B.n13 B.n12 163.367
R967 B.n14 B.n13 163.367
R968 B.n864 B.n14 163.367
R969 B.n864 B.n19 163.367
R970 B.n20 B.n19 163.367
R971 B.n21 B.n20 163.367
R972 B.n869 B.n21 163.367
R973 B.n869 B.n26 163.367
R974 B.n27 B.n26 163.367
R975 B.n28 B.n27 163.367
R976 B.n874 B.n28 163.367
R977 B.n874 B.n33 163.367
R978 B.n34 B.n33 163.367
R979 B.n35 B.n34 163.367
R980 B.n879 B.n35 163.367
R981 B.n879 B.n40 163.367
R982 B.n41 B.n40 163.367
R983 B.n42 B.n41 163.367
R984 B.n884 B.n42 163.367
R985 B.n884 B.n47 163.367
R986 B.n48 B.n47 163.367
R987 B.n49 B.n48 163.367
R988 B.n889 B.n49 163.367
R989 B.n889 B.n54 163.367
R990 B.n55 B.n54 163.367
R991 B.n56 B.n55 163.367
R992 B.n894 B.n56 163.367
R993 B.n894 B.n61 163.367
R994 B.n62 B.n61 163.367
R995 B.n63 B.n62 163.367
R996 B.n899 B.n63 163.367
R997 B.n899 B.n68 163.367
R998 B.n69 B.n68 163.367
R999 B.n70 B.n69 163.367
R1000 B.n904 B.n70 163.367
R1001 B.n904 B.n75 163.367
R1002 B.n76 B.n75 163.367
R1003 B.n77 B.n76 163.367
R1004 B.n909 B.n77 163.367
R1005 B.n909 B.n82 163.367
R1006 B.n83 B.n82 163.367
R1007 B.n84 B.n83 163.367
R1008 B.n914 B.n84 163.367
R1009 B.n914 B.n89 163.367
R1010 B.n90 B.n89 163.367
R1011 B.n91 B.n90 163.367
R1012 B.n919 B.n91 163.367
R1013 B.n919 B.n96 163.367
R1014 B.n97 B.n96 163.367
R1015 B.n98 B.n97 163.367
R1016 B.n924 B.n98 163.367
R1017 B.n924 B.n103 163.367
R1018 B.n104 B.n103 163.367
R1019 B.n159 B.n158 163.367
R1020 B.n163 B.n162 163.367
R1021 B.n167 B.n166 163.367
R1022 B.n171 B.n170 163.367
R1023 B.n175 B.n174 163.367
R1024 B.n179 B.n178 163.367
R1025 B.n183 B.n182 163.367
R1026 B.n187 B.n186 163.367
R1027 B.n191 B.n190 163.367
R1028 B.n195 B.n194 163.367
R1029 B.n199 B.n198 163.367
R1030 B.n203 B.n202 163.367
R1031 B.n207 B.n206 163.367
R1032 B.n211 B.n210 163.367
R1033 B.n215 B.n214 163.367
R1034 B.n219 B.n218 163.367
R1035 B.n223 B.n222 163.367
R1036 B.n227 B.n226 163.367
R1037 B.n231 B.n230 163.367
R1038 B.n235 B.n234 163.367
R1039 B.n240 B.n239 163.367
R1040 B.n244 B.n243 163.367
R1041 B.n248 B.n247 163.367
R1042 B.n252 B.n251 163.367
R1043 B.n256 B.n255 163.367
R1044 B.n261 B.n260 163.367
R1045 B.n265 B.n264 163.367
R1046 B.n269 B.n268 163.367
R1047 B.n273 B.n272 163.367
R1048 B.n277 B.n276 163.367
R1049 B.n281 B.n280 163.367
R1050 B.n285 B.n284 163.367
R1051 B.n289 B.n288 163.367
R1052 B.n293 B.n292 163.367
R1053 B.n297 B.n296 163.367
R1054 B.n301 B.n300 163.367
R1055 B.n305 B.n304 163.367
R1056 B.n309 B.n308 163.367
R1057 B.n313 B.n312 163.367
R1058 B.n317 B.n316 163.367
R1059 B.n321 B.n320 163.367
R1060 B.n325 B.n324 163.367
R1061 B.n329 B.n328 163.367
R1062 B.n333 B.n332 163.367
R1063 B.n335 B.n150 163.367
R1064 B.n499 B.t18 137.248
R1065 B.n151 B.t14 137.248
R1066 B.n496 B.t11 137.232
R1067 B.n153 B.t20 137.232
R1068 B.n681 B.n446 89.5466
R1069 B.n932 B.n931 89.5466
R1070 B.n500 B.t17 72.4719
R1071 B.n152 B.t15 72.4719
R1072 B.n497 B.t10 72.4572
R1073 B.n154 B.t21 72.4572
R1074 B.n680 B.n679 71.676
R1075 B.n674 B.n450 71.676
R1076 B.n671 B.n451 71.676
R1077 B.n667 B.n452 71.676
R1078 B.n663 B.n453 71.676
R1079 B.n659 B.n454 71.676
R1080 B.n655 B.n455 71.676
R1081 B.n651 B.n456 71.676
R1082 B.n647 B.n457 71.676
R1083 B.n643 B.n458 71.676
R1084 B.n639 B.n459 71.676
R1085 B.n635 B.n460 71.676
R1086 B.n631 B.n461 71.676
R1087 B.n627 B.n462 71.676
R1088 B.n623 B.n463 71.676
R1089 B.n619 B.n464 71.676
R1090 B.n615 B.n465 71.676
R1091 B.n611 B.n466 71.676
R1092 B.n607 B.n467 71.676
R1093 B.n603 B.n468 71.676
R1094 B.n599 B.n469 71.676
R1095 B.n595 B.n470 71.676
R1096 B.n591 B.n471 71.676
R1097 B.n587 B.n472 71.676
R1098 B.n583 B.n473 71.676
R1099 B.n579 B.n474 71.676
R1100 B.n575 B.n475 71.676
R1101 B.n571 B.n476 71.676
R1102 B.n567 B.n477 71.676
R1103 B.n563 B.n478 71.676
R1104 B.n559 B.n479 71.676
R1105 B.n555 B.n480 71.676
R1106 B.n551 B.n481 71.676
R1107 B.n547 B.n482 71.676
R1108 B.n543 B.n483 71.676
R1109 B.n539 B.n484 71.676
R1110 B.n535 B.n485 71.676
R1111 B.n531 B.n486 71.676
R1112 B.n527 B.n487 71.676
R1113 B.n523 B.n488 71.676
R1114 B.n519 B.n489 71.676
R1115 B.n515 B.n490 71.676
R1116 B.n511 B.n491 71.676
R1117 B.n507 B.n492 71.676
R1118 B.n503 B.n493 71.676
R1119 B.n155 B.n105 71.676
R1120 B.n159 B.n106 71.676
R1121 B.n163 B.n107 71.676
R1122 B.n167 B.n108 71.676
R1123 B.n171 B.n109 71.676
R1124 B.n175 B.n110 71.676
R1125 B.n179 B.n111 71.676
R1126 B.n183 B.n112 71.676
R1127 B.n187 B.n113 71.676
R1128 B.n191 B.n114 71.676
R1129 B.n195 B.n115 71.676
R1130 B.n199 B.n116 71.676
R1131 B.n203 B.n117 71.676
R1132 B.n207 B.n118 71.676
R1133 B.n211 B.n119 71.676
R1134 B.n215 B.n120 71.676
R1135 B.n219 B.n121 71.676
R1136 B.n223 B.n122 71.676
R1137 B.n227 B.n123 71.676
R1138 B.n231 B.n124 71.676
R1139 B.n235 B.n125 71.676
R1140 B.n240 B.n126 71.676
R1141 B.n244 B.n127 71.676
R1142 B.n248 B.n128 71.676
R1143 B.n252 B.n129 71.676
R1144 B.n256 B.n130 71.676
R1145 B.n261 B.n131 71.676
R1146 B.n265 B.n132 71.676
R1147 B.n269 B.n133 71.676
R1148 B.n273 B.n134 71.676
R1149 B.n277 B.n135 71.676
R1150 B.n281 B.n136 71.676
R1151 B.n285 B.n137 71.676
R1152 B.n289 B.n138 71.676
R1153 B.n293 B.n139 71.676
R1154 B.n297 B.n140 71.676
R1155 B.n301 B.n141 71.676
R1156 B.n305 B.n142 71.676
R1157 B.n309 B.n143 71.676
R1158 B.n313 B.n144 71.676
R1159 B.n317 B.n145 71.676
R1160 B.n321 B.n146 71.676
R1161 B.n325 B.n147 71.676
R1162 B.n329 B.n148 71.676
R1163 B.n333 B.n149 71.676
R1164 B.n930 B.n150 71.676
R1165 B.n930 B.n929 71.676
R1166 B.n335 B.n149 71.676
R1167 B.n332 B.n148 71.676
R1168 B.n328 B.n147 71.676
R1169 B.n324 B.n146 71.676
R1170 B.n320 B.n145 71.676
R1171 B.n316 B.n144 71.676
R1172 B.n312 B.n143 71.676
R1173 B.n308 B.n142 71.676
R1174 B.n304 B.n141 71.676
R1175 B.n300 B.n140 71.676
R1176 B.n296 B.n139 71.676
R1177 B.n292 B.n138 71.676
R1178 B.n288 B.n137 71.676
R1179 B.n284 B.n136 71.676
R1180 B.n280 B.n135 71.676
R1181 B.n276 B.n134 71.676
R1182 B.n272 B.n133 71.676
R1183 B.n268 B.n132 71.676
R1184 B.n264 B.n131 71.676
R1185 B.n260 B.n130 71.676
R1186 B.n255 B.n129 71.676
R1187 B.n251 B.n128 71.676
R1188 B.n247 B.n127 71.676
R1189 B.n243 B.n126 71.676
R1190 B.n239 B.n125 71.676
R1191 B.n234 B.n124 71.676
R1192 B.n230 B.n123 71.676
R1193 B.n226 B.n122 71.676
R1194 B.n222 B.n121 71.676
R1195 B.n218 B.n120 71.676
R1196 B.n214 B.n119 71.676
R1197 B.n210 B.n118 71.676
R1198 B.n206 B.n117 71.676
R1199 B.n202 B.n116 71.676
R1200 B.n198 B.n115 71.676
R1201 B.n194 B.n114 71.676
R1202 B.n190 B.n113 71.676
R1203 B.n186 B.n112 71.676
R1204 B.n182 B.n111 71.676
R1205 B.n178 B.n110 71.676
R1206 B.n174 B.n109 71.676
R1207 B.n170 B.n108 71.676
R1208 B.n166 B.n107 71.676
R1209 B.n162 B.n106 71.676
R1210 B.n158 B.n105 71.676
R1211 B.n680 B.n495 71.676
R1212 B.n672 B.n450 71.676
R1213 B.n668 B.n451 71.676
R1214 B.n664 B.n452 71.676
R1215 B.n660 B.n453 71.676
R1216 B.n656 B.n454 71.676
R1217 B.n652 B.n455 71.676
R1218 B.n648 B.n456 71.676
R1219 B.n644 B.n457 71.676
R1220 B.n640 B.n458 71.676
R1221 B.n636 B.n459 71.676
R1222 B.n632 B.n460 71.676
R1223 B.n628 B.n461 71.676
R1224 B.n624 B.n462 71.676
R1225 B.n620 B.n463 71.676
R1226 B.n616 B.n464 71.676
R1227 B.n612 B.n465 71.676
R1228 B.n608 B.n466 71.676
R1229 B.n604 B.n467 71.676
R1230 B.n600 B.n468 71.676
R1231 B.n596 B.n469 71.676
R1232 B.n592 B.n470 71.676
R1233 B.n588 B.n471 71.676
R1234 B.n584 B.n472 71.676
R1235 B.n580 B.n473 71.676
R1236 B.n576 B.n474 71.676
R1237 B.n572 B.n475 71.676
R1238 B.n568 B.n476 71.676
R1239 B.n564 B.n477 71.676
R1240 B.n560 B.n478 71.676
R1241 B.n556 B.n479 71.676
R1242 B.n552 B.n480 71.676
R1243 B.n548 B.n481 71.676
R1244 B.n544 B.n482 71.676
R1245 B.n540 B.n483 71.676
R1246 B.n536 B.n484 71.676
R1247 B.n532 B.n485 71.676
R1248 B.n528 B.n486 71.676
R1249 B.n524 B.n487 71.676
R1250 B.n520 B.n488 71.676
R1251 B.n516 B.n489 71.676
R1252 B.n512 B.n490 71.676
R1253 B.n508 B.n491 71.676
R1254 B.n504 B.n492 71.676
R1255 B.n493 B.n449 71.676
R1256 B.n500 B.n499 64.7763
R1257 B.n497 B.n496 64.7763
R1258 B.n154 B.n153 64.7763
R1259 B.n152 B.n151 64.7763
R1260 B.n501 B.n500 59.5399
R1261 B.n498 B.n497 59.5399
R1262 B.n237 B.n154 59.5399
R1263 B.n258 B.n152 59.5399
R1264 B.n687 B.n446 43.8072
R1265 B.n687 B.n442 43.8072
R1266 B.n693 B.n442 43.8072
R1267 B.n693 B.n438 43.8072
R1268 B.n699 B.n438 43.8072
R1269 B.n699 B.n434 43.8072
R1270 B.n705 B.n434 43.8072
R1271 B.n711 B.n430 43.8072
R1272 B.n711 B.n426 43.8072
R1273 B.n717 B.n426 43.8072
R1274 B.n717 B.n422 43.8072
R1275 B.n723 B.n422 43.8072
R1276 B.n723 B.n418 43.8072
R1277 B.n729 B.n418 43.8072
R1278 B.n729 B.n414 43.8072
R1279 B.n735 B.n414 43.8072
R1280 B.n735 B.n410 43.8072
R1281 B.n741 B.n410 43.8072
R1282 B.n741 B.n406 43.8072
R1283 B.n747 B.n406 43.8072
R1284 B.n753 B.n402 43.8072
R1285 B.n753 B.n398 43.8072
R1286 B.n759 B.n398 43.8072
R1287 B.n759 B.n394 43.8072
R1288 B.n765 B.n394 43.8072
R1289 B.n765 B.n390 43.8072
R1290 B.n772 B.n390 43.8072
R1291 B.n772 B.n771 43.8072
R1292 B.n778 B.n383 43.8072
R1293 B.n784 B.n383 43.8072
R1294 B.n784 B.n379 43.8072
R1295 B.n790 B.n379 43.8072
R1296 B.n790 B.n375 43.8072
R1297 B.n796 B.n375 43.8072
R1298 B.n796 B.n370 43.8072
R1299 B.n802 B.n370 43.8072
R1300 B.n802 B.n371 43.8072
R1301 B.n808 B.n363 43.8072
R1302 B.n814 B.n363 43.8072
R1303 B.n814 B.n359 43.8072
R1304 B.n820 B.n359 43.8072
R1305 B.n820 B.n355 43.8072
R1306 B.n826 B.n355 43.8072
R1307 B.n826 B.n351 43.8072
R1308 B.n833 B.n351 43.8072
R1309 B.n833 B.n832 43.8072
R1310 B.n839 B.n344 43.8072
R1311 B.n846 B.n344 43.8072
R1312 B.n846 B.n340 43.8072
R1313 B.n852 B.n340 43.8072
R1314 B.n852 B.n4 43.8072
R1315 B.n1045 B.n4 43.8072
R1316 B.n1045 B.n1044 43.8072
R1317 B.n1044 B.n1043 43.8072
R1318 B.n1043 B.n8 43.8072
R1319 B.n1037 B.n8 43.8072
R1320 B.n1037 B.n1036 43.8072
R1321 B.n1036 B.n1035 43.8072
R1322 B.n1029 B.n18 43.8072
R1323 B.n1029 B.n1028 43.8072
R1324 B.n1028 B.n1027 43.8072
R1325 B.n1027 B.n22 43.8072
R1326 B.n1021 B.n22 43.8072
R1327 B.n1021 B.n1020 43.8072
R1328 B.n1020 B.n1019 43.8072
R1329 B.n1019 B.n29 43.8072
R1330 B.n1013 B.n29 43.8072
R1331 B.n1012 B.n1011 43.8072
R1332 B.n1011 B.n36 43.8072
R1333 B.n1005 B.n36 43.8072
R1334 B.n1005 B.n1004 43.8072
R1335 B.n1004 B.n1003 43.8072
R1336 B.n1003 B.n43 43.8072
R1337 B.n997 B.n43 43.8072
R1338 B.n997 B.n996 43.8072
R1339 B.n996 B.n995 43.8072
R1340 B.n989 B.n53 43.8072
R1341 B.n989 B.n988 43.8072
R1342 B.n988 B.n987 43.8072
R1343 B.n987 B.n57 43.8072
R1344 B.n981 B.n57 43.8072
R1345 B.n981 B.n980 43.8072
R1346 B.n980 B.n979 43.8072
R1347 B.n979 B.n64 43.8072
R1348 B.n973 B.n972 43.8072
R1349 B.n972 B.n971 43.8072
R1350 B.n971 B.n71 43.8072
R1351 B.n965 B.n71 43.8072
R1352 B.n965 B.n964 43.8072
R1353 B.n964 B.n963 43.8072
R1354 B.n963 B.n78 43.8072
R1355 B.n957 B.n78 43.8072
R1356 B.n957 B.n956 43.8072
R1357 B.n956 B.n955 43.8072
R1358 B.n955 B.n85 43.8072
R1359 B.n949 B.n85 43.8072
R1360 B.n949 B.n948 43.8072
R1361 B.n947 B.n92 43.8072
R1362 B.n941 B.n92 43.8072
R1363 B.n941 B.n940 43.8072
R1364 B.n940 B.n939 43.8072
R1365 B.n939 B.n99 43.8072
R1366 B.n933 B.n99 43.8072
R1367 B.n933 B.n932 43.8072
R1368 B.n705 B.t9 43.163
R1369 B.t2 B.n402 43.163
R1370 B.t0 B.n64 43.163
R1371 B.t13 B.n947 43.163
R1372 B.n771 B.t6 36.7209
R1373 B.n53 B.t7 36.7209
R1374 B.n156 B.n101 32.9371
R1375 B.n928 B.n927 32.9371
R1376 B.n684 B.n683 32.9371
R1377 B.n678 B.n444 32.9371
R1378 B.n371 B.t4 28.9903
R1379 B.t3 B.n1012 28.9903
R1380 B.n839 B.t1 22.5481
R1381 B.n1035 B.t5 22.5481
R1382 B.n832 B.t1 21.2596
R1383 B.n18 B.t5 21.2596
R1384 B B.n1047 18.0485
R1385 B.n808 B.t4 14.8175
R1386 B.n1013 B.t3 14.8175
R1387 B.n157 B.n156 10.6151
R1388 B.n160 B.n157 10.6151
R1389 B.n161 B.n160 10.6151
R1390 B.n164 B.n161 10.6151
R1391 B.n165 B.n164 10.6151
R1392 B.n168 B.n165 10.6151
R1393 B.n169 B.n168 10.6151
R1394 B.n172 B.n169 10.6151
R1395 B.n173 B.n172 10.6151
R1396 B.n176 B.n173 10.6151
R1397 B.n177 B.n176 10.6151
R1398 B.n180 B.n177 10.6151
R1399 B.n181 B.n180 10.6151
R1400 B.n184 B.n181 10.6151
R1401 B.n185 B.n184 10.6151
R1402 B.n188 B.n185 10.6151
R1403 B.n189 B.n188 10.6151
R1404 B.n192 B.n189 10.6151
R1405 B.n193 B.n192 10.6151
R1406 B.n196 B.n193 10.6151
R1407 B.n197 B.n196 10.6151
R1408 B.n200 B.n197 10.6151
R1409 B.n201 B.n200 10.6151
R1410 B.n204 B.n201 10.6151
R1411 B.n205 B.n204 10.6151
R1412 B.n208 B.n205 10.6151
R1413 B.n209 B.n208 10.6151
R1414 B.n212 B.n209 10.6151
R1415 B.n213 B.n212 10.6151
R1416 B.n216 B.n213 10.6151
R1417 B.n217 B.n216 10.6151
R1418 B.n220 B.n217 10.6151
R1419 B.n221 B.n220 10.6151
R1420 B.n224 B.n221 10.6151
R1421 B.n225 B.n224 10.6151
R1422 B.n228 B.n225 10.6151
R1423 B.n229 B.n228 10.6151
R1424 B.n232 B.n229 10.6151
R1425 B.n233 B.n232 10.6151
R1426 B.n236 B.n233 10.6151
R1427 B.n241 B.n238 10.6151
R1428 B.n242 B.n241 10.6151
R1429 B.n245 B.n242 10.6151
R1430 B.n246 B.n245 10.6151
R1431 B.n249 B.n246 10.6151
R1432 B.n250 B.n249 10.6151
R1433 B.n253 B.n250 10.6151
R1434 B.n254 B.n253 10.6151
R1435 B.n257 B.n254 10.6151
R1436 B.n262 B.n259 10.6151
R1437 B.n263 B.n262 10.6151
R1438 B.n266 B.n263 10.6151
R1439 B.n267 B.n266 10.6151
R1440 B.n270 B.n267 10.6151
R1441 B.n271 B.n270 10.6151
R1442 B.n274 B.n271 10.6151
R1443 B.n275 B.n274 10.6151
R1444 B.n278 B.n275 10.6151
R1445 B.n279 B.n278 10.6151
R1446 B.n282 B.n279 10.6151
R1447 B.n283 B.n282 10.6151
R1448 B.n286 B.n283 10.6151
R1449 B.n287 B.n286 10.6151
R1450 B.n290 B.n287 10.6151
R1451 B.n291 B.n290 10.6151
R1452 B.n294 B.n291 10.6151
R1453 B.n295 B.n294 10.6151
R1454 B.n298 B.n295 10.6151
R1455 B.n299 B.n298 10.6151
R1456 B.n302 B.n299 10.6151
R1457 B.n303 B.n302 10.6151
R1458 B.n306 B.n303 10.6151
R1459 B.n307 B.n306 10.6151
R1460 B.n310 B.n307 10.6151
R1461 B.n311 B.n310 10.6151
R1462 B.n314 B.n311 10.6151
R1463 B.n315 B.n314 10.6151
R1464 B.n318 B.n315 10.6151
R1465 B.n319 B.n318 10.6151
R1466 B.n322 B.n319 10.6151
R1467 B.n323 B.n322 10.6151
R1468 B.n326 B.n323 10.6151
R1469 B.n327 B.n326 10.6151
R1470 B.n330 B.n327 10.6151
R1471 B.n331 B.n330 10.6151
R1472 B.n334 B.n331 10.6151
R1473 B.n336 B.n334 10.6151
R1474 B.n337 B.n336 10.6151
R1475 B.n928 B.n337 10.6151
R1476 B.n685 B.n684 10.6151
R1477 B.n685 B.n440 10.6151
R1478 B.n695 B.n440 10.6151
R1479 B.n696 B.n695 10.6151
R1480 B.n697 B.n696 10.6151
R1481 B.n697 B.n432 10.6151
R1482 B.n707 B.n432 10.6151
R1483 B.n708 B.n707 10.6151
R1484 B.n709 B.n708 10.6151
R1485 B.n709 B.n424 10.6151
R1486 B.n719 B.n424 10.6151
R1487 B.n720 B.n719 10.6151
R1488 B.n721 B.n720 10.6151
R1489 B.n721 B.n416 10.6151
R1490 B.n731 B.n416 10.6151
R1491 B.n732 B.n731 10.6151
R1492 B.n733 B.n732 10.6151
R1493 B.n733 B.n408 10.6151
R1494 B.n743 B.n408 10.6151
R1495 B.n744 B.n743 10.6151
R1496 B.n745 B.n744 10.6151
R1497 B.n745 B.n400 10.6151
R1498 B.n755 B.n400 10.6151
R1499 B.n756 B.n755 10.6151
R1500 B.n757 B.n756 10.6151
R1501 B.n757 B.n392 10.6151
R1502 B.n767 B.n392 10.6151
R1503 B.n768 B.n767 10.6151
R1504 B.n769 B.n768 10.6151
R1505 B.n769 B.n385 10.6151
R1506 B.n780 B.n385 10.6151
R1507 B.n781 B.n780 10.6151
R1508 B.n782 B.n781 10.6151
R1509 B.n782 B.n377 10.6151
R1510 B.n792 B.n377 10.6151
R1511 B.n793 B.n792 10.6151
R1512 B.n794 B.n793 10.6151
R1513 B.n794 B.n368 10.6151
R1514 B.n804 B.n368 10.6151
R1515 B.n805 B.n804 10.6151
R1516 B.n806 B.n805 10.6151
R1517 B.n806 B.n361 10.6151
R1518 B.n816 B.n361 10.6151
R1519 B.n817 B.n816 10.6151
R1520 B.n818 B.n817 10.6151
R1521 B.n818 B.n353 10.6151
R1522 B.n828 B.n353 10.6151
R1523 B.n829 B.n828 10.6151
R1524 B.n830 B.n829 10.6151
R1525 B.n830 B.n346 10.6151
R1526 B.n841 B.n346 10.6151
R1527 B.n842 B.n841 10.6151
R1528 B.n844 B.n842 10.6151
R1529 B.n844 B.n843 10.6151
R1530 B.n843 B.n338 10.6151
R1531 B.n855 B.n338 10.6151
R1532 B.n856 B.n855 10.6151
R1533 B.n857 B.n856 10.6151
R1534 B.n858 B.n857 10.6151
R1535 B.n860 B.n858 10.6151
R1536 B.n861 B.n860 10.6151
R1537 B.n862 B.n861 10.6151
R1538 B.n863 B.n862 10.6151
R1539 B.n865 B.n863 10.6151
R1540 B.n866 B.n865 10.6151
R1541 B.n867 B.n866 10.6151
R1542 B.n868 B.n867 10.6151
R1543 B.n870 B.n868 10.6151
R1544 B.n871 B.n870 10.6151
R1545 B.n872 B.n871 10.6151
R1546 B.n873 B.n872 10.6151
R1547 B.n875 B.n873 10.6151
R1548 B.n876 B.n875 10.6151
R1549 B.n877 B.n876 10.6151
R1550 B.n878 B.n877 10.6151
R1551 B.n880 B.n878 10.6151
R1552 B.n881 B.n880 10.6151
R1553 B.n882 B.n881 10.6151
R1554 B.n883 B.n882 10.6151
R1555 B.n885 B.n883 10.6151
R1556 B.n886 B.n885 10.6151
R1557 B.n887 B.n886 10.6151
R1558 B.n888 B.n887 10.6151
R1559 B.n890 B.n888 10.6151
R1560 B.n891 B.n890 10.6151
R1561 B.n892 B.n891 10.6151
R1562 B.n893 B.n892 10.6151
R1563 B.n895 B.n893 10.6151
R1564 B.n896 B.n895 10.6151
R1565 B.n897 B.n896 10.6151
R1566 B.n898 B.n897 10.6151
R1567 B.n900 B.n898 10.6151
R1568 B.n901 B.n900 10.6151
R1569 B.n902 B.n901 10.6151
R1570 B.n903 B.n902 10.6151
R1571 B.n905 B.n903 10.6151
R1572 B.n906 B.n905 10.6151
R1573 B.n907 B.n906 10.6151
R1574 B.n908 B.n907 10.6151
R1575 B.n910 B.n908 10.6151
R1576 B.n911 B.n910 10.6151
R1577 B.n912 B.n911 10.6151
R1578 B.n913 B.n912 10.6151
R1579 B.n915 B.n913 10.6151
R1580 B.n916 B.n915 10.6151
R1581 B.n917 B.n916 10.6151
R1582 B.n918 B.n917 10.6151
R1583 B.n920 B.n918 10.6151
R1584 B.n921 B.n920 10.6151
R1585 B.n922 B.n921 10.6151
R1586 B.n923 B.n922 10.6151
R1587 B.n925 B.n923 10.6151
R1588 B.n926 B.n925 10.6151
R1589 B.n927 B.n926 10.6151
R1590 B.n678 B.n677 10.6151
R1591 B.n677 B.n676 10.6151
R1592 B.n676 B.n675 10.6151
R1593 B.n675 B.n673 10.6151
R1594 B.n673 B.n670 10.6151
R1595 B.n670 B.n669 10.6151
R1596 B.n669 B.n666 10.6151
R1597 B.n666 B.n665 10.6151
R1598 B.n665 B.n662 10.6151
R1599 B.n662 B.n661 10.6151
R1600 B.n661 B.n658 10.6151
R1601 B.n658 B.n657 10.6151
R1602 B.n657 B.n654 10.6151
R1603 B.n654 B.n653 10.6151
R1604 B.n653 B.n650 10.6151
R1605 B.n650 B.n649 10.6151
R1606 B.n649 B.n646 10.6151
R1607 B.n646 B.n645 10.6151
R1608 B.n645 B.n642 10.6151
R1609 B.n642 B.n641 10.6151
R1610 B.n641 B.n638 10.6151
R1611 B.n638 B.n637 10.6151
R1612 B.n637 B.n634 10.6151
R1613 B.n634 B.n633 10.6151
R1614 B.n633 B.n630 10.6151
R1615 B.n630 B.n629 10.6151
R1616 B.n629 B.n626 10.6151
R1617 B.n626 B.n625 10.6151
R1618 B.n625 B.n622 10.6151
R1619 B.n622 B.n621 10.6151
R1620 B.n621 B.n618 10.6151
R1621 B.n618 B.n617 10.6151
R1622 B.n617 B.n614 10.6151
R1623 B.n614 B.n613 10.6151
R1624 B.n613 B.n610 10.6151
R1625 B.n610 B.n609 10.6151
R1626 B.n609 B.n606 10.6151
R1627 B.n606 B.n605 10.6151
R1628 B.n605 B.n602 10.6151
R1629 B.n602 B.n601 10.6151
R1630 B.n598 B.n597 10.6151
R1631 B.n597 B.n594 10.6151
R1632 B.n594 B.n593 10.6151
R1633 B.n593 B.n590 10.6151
R1634 B.n590 B.n589 10.6151
R1635 B.n589 B.n586 10.6151
R1636 B.n586 B.n585 10.6151
R1637 B.n585 B.n582 10.6151
R1638 B.n582 B.n581 10.6151
R1639 B.n578 B.n577 10.6151
R1640 B.n577 B.n574 10.6151
R1641 B.n574 B.n573 10.6151
R1642 B.n573 B.n570 10.6151
R1643 B.n570 B.n569 10.6151
R1644 B.n569 B.n566 10.6151
R1645 B.n566 B.n565 10.6151
R1646 B.n565 B.n562 10.6151
R1647 B.n562 B.n561 10.6151
R1648 B.n561 B.n558 10.6151
R1649 B.n558 B.n557 10.6151
R1650 B.n557 B.n554 10.6151
R1651 B.n554 B.n553 10.6151
R1652 B.n553 B.n550 10.6151
R1653 B.n550 B.n549 10.6151
R1654 B.n549 B.n546 10.6151
R1655 B.n546 B.n545 10.6151
R1656 B.n545 B.n542 10.6151
R1657 B.n542 B.n541 10.6151
R1658 B.n541 B.n538 10.6151
R1659 B.n538 B.n537 10.6151
R1660 B.n537 B.n534 10.6151
R1661 B.n534 B.n533 10.6151
R1662 B.n533 B.n530 10.6151
R1663 B.n530 B.n529 10.6151
R1664 B.n529 B.n526 10.6151
R1665 B.n526 B.n525 10.6151
R1666 B.n525 B.n522 10.6151
R1667 B.n522 B.n521 10.6151
R1668 B.n521 B.n518 10.6151
R1669 B.n518 B.n517 10.6151
R1670 B.n517 B.n514 10.6151
R1671 B.n514 B.n513 10.6151
R1672 B.n513 B.n510 10.6151
R1673 B.n510 B.n509 10.6151
R1674 B.n509 B.n506 10.6151
R1675 B.n506 B.n505 10.6151
R1676 B.n505 B.n502 10.6151
R1677 B.n502 B.n448 10.6151
R1678 B.n683 B.n448 10.6151
R1679 B.n689 B.n444 10.6151
R1680 B.n690 B.n689 10.6151
R1681 B.n691 B.n690 10.6151
R1682 B.n691 B.n436 10.6151
R1683 B.n701 B.n436 10.6151
R1684 B.n702 B.n701 10.6151
R1685 B.n703 B.n702 10.6151
R1686 B.n703 B.n428 10.6151
R1687 B.n713 B.n428 10.6151
R1688 B.n714 B.n713 10.6151
R1689 B.n715 B.n714 10.6151
R1690 B.n715 B.n420 10.6151
R1691 B.n725 B.n420 10.6151
R1692 B.n726 B.n725 10.6151
R1693 B.n727 B.n726 10.6151
R1694 B.n727 B.n412 10.6151
R1695 B.n737 B.n412 10.6151
R1696 B.n738 B.n737 10.6151
R1697 B.n739 B.n738 10.6151
R1698 B.n739 B.n404 10.6151
R1699 B.n749 B.n404 10.6151
R1700 B.n750 B.n749 10.6151
R1701 B.n751 B.n750 10.6151
R1702 B.n751 B.n396 10.6151
R1703 B.n761 B.n396 10.6151
R1704 B.n762 B.n761 10.6151
R1705 B.n763 B.n762 10.6151
R1706 B.n763 B.n388 10.6151
R1707 B.n774 B.n388 10.6151
R1708 B.n775 B.n774 10.6151
R1709 B.n776 B.n775 10.6151
R1710 B.n776 B.n381 10.6151
R1711 B.n786 B.n381 10.6151
R1712 B.n787 B.n786 10.6151
R1713 B.n788 B.n787 10.6151
R1714 B.n788 B.n373 10.6151
R1715 B.n798 B.n373 10.6151
R1716 B.n799 B.n798 10.6151
R1717 B.n800 B.n799 10.6151
R1718 B.n800 B.n365 10.6151
R1719 B.n810 B.n365 10.6151
R1720 B.n811 B.n810 10.6151
R1721 B.n812 B.n811 10.6151
R1722 B.n812 B.n357 10.6151
R1723 B.n822 B.n357 10.6151
R1724 B.n823 B.n822 10.6151
R1725 B.n824 B.n823 10.6151
R1726 B.n824 B.n349 10.6151
R1727 B.n835 B.n349 10.6151
R1728 B.n836 B.n835 10.6151
R1729 B.n837 B.n836 10.6151
R1730 B.n837 B.n342 10.6151
R1731 B.n848 B.n342 10.6151
R1732 B.n849 B.n848 10.6151
R1733 B.n850 B.n849 10.6151
R1734 B.n850 B.n0 10.6151
R1735 B.n1041 B.n1 10.6151
R1736 B.n1041 B.n1040 10.6151
R1737 B.n1040 B.n1039 10.6151
R1738 B.n1039 B.n10 10.6151
R1739 B.n1033 B.n10 10.6151
R1740 B.n1033 B.n1032 10.6151
R1741 B.n1032 B.n1031 10.6151
R1742 B.n1031 B.n16 10.6151
R1743 B.n1025 B.n16 10.6151
R1744 B.n1025 B.n1024 10.6151
R1745 B.n1024 B.n1023 10.6151
R1746 B.n1023 B.n24 10.6151
R1747 B.n1017 B.n24 10.6151
R1748 B.n1017 B.n1016 10.6151
R1749 B.n1016 B.n1015 10.6151
R1750 B.n1015 B.n31 10.6151
R1751 B.n1009 B.n31 10.6151
R1752 B.n1009 B.n1008 10.6151
R1753 B.n1008 B.n1007 10.6151
R1754 B.n1007 B.n38 10.6151
R1755 B.n1001 B.n38 10.6151
R1756 B.n1001 B.n1000 10.6151
R1757 B.n1000 B.n999 10.6151
R1758 B.n999 B.n45 10.6151
R1759 B.n993 B.n45 10.6151
R1760 B.n993 B.n992 10.6151
R1761 B.n992 B.n991 10.6151
R1762 B.n991 B.n51 10.6151
R1763 B.n985 B.n51 10.6151
R1764 B.n985 B.n984 10.6151
R1765 B.n984 B.n983 10.6151
R1766 B.n983 B.n59 10.6151
R1767 B.n977 B.n59 10.6151
R1768 B.n977 B.n976 10.6151
R1769 B.n976 B.n975 10.6151
R1770 B.n975 B.n66 10.6151
R1771 B.n969 B.n66 10.6151
R1772 B.n969 B.n968 10.6151
R1773 B.n968 B.n967 10.6151
R1774 B.n967 B.n73 10.6151
R1775 B.n961 B.n73 10.6151
R1776 B.n961 B.n960 10.6151
R1777 B.n960 B.n959 10.6151
R1778 B.n959 B.n80 10.6151
R1779 B.n953 B.n80 10.6151
R1780 B.n953 B.n952 10.6151
R1781 B.n952 B.n951 10.6151
R1782 B.n951 B.n87 10.6151
R1783 B.n945 B.n87 10.6151
R1784 B.n945 B.n944 10.6151
R1785 B.n944 B.n943 10.6151
R1786 B.n943 B.n94 10.6151
R1787 B.n937 B.n94 10.6151
R1788 B.n937 B.n936 10.6151
R1789 B.n936 B.n935 10.6151
R1790 B.n935 B.n101 10.6151
R1791 B.n237 B.n236 9.36635
R1792 B.n259 B.n258 9.36635
R1793 B.n601 B.n498 9.36635
R1794 B.n578 B.n501 9.36635
R1795 B.n778 B.t6 7.08688
R1796 B.n995 B.t7 7.08688
R1797 B.n1047 B.n0 2.81026
R1798 B.n1047 B.n1 2.81026
R1799 B.n238 B.n237 1.24928
R1800 B.n258 B.n257 1.24928
R1801 B.n598 B.n498 1.24928
R1802 B.n581 B.n501 1.24928
R1803 B.t9 B.n430 0.644717
R1804 B.n747 B.t2 0.644717
R1805 B.n973 B.t0 0.644717
R1806 B.n948 B.t13 0.644717
R1807 VP.n22 VP.n21 161.3
R1808 VP.n23 VP.n18 161.3
R1809 VP.n25 VP.n24 161.3
R1810 VP.n26 VP.n17 161.3
R1811 VP.n28 VP.n27 161.3
R1812 VP.n29 VP.n16 161.3
R1813 VP.n32 VP.n31 161.3
R1814 VP.n33 VP.n15 161.3
R1815 VP.n35 VP.n34 161.3
R1816 VP.n36 VP.n14 161.3
R1817 VP.n38 VP.n37 161.3
R1818 VP.n39 VP.n13 161.3
R1819 VP.n41 VP.n40 161.3
R1820 VP.n42 VP.n12 161.3
R1821 VP.n78 VP.n0 161.3
R1822 VP.n77 VP.n76 161.3
R1823 VP.n75 VP.n1 161.3
R1824 VP.n74 VP.n73 161.3
R1825 VP.n72 VP.n2 161.3
R1826 VP.n71 VP.n70 161.3
R1827 VP.n69 VP.n3 161.3
R1828 VP.n68 VP.n67 161.3
R1829 VP.n65 VP.n4 161.3
R1830 VP.n64 VP.n63 161.3
R1831 VP.n62 VP.n5 161.3
R1832 VP.n61 VP.n60 161.3
R1833 VP.n59 VP.n6 161.3
R1834 VP.n58 VP.n57 161.3
R1835 VP.n56 VP.n55 161.3
R1836 VP.n54 VP.n8 161.3
R1837 VP.n53 VP.n52 161.3
R1838 VP.n51 VP.n9 161.3
R1839 VP.n50 VP.n49 161.3
R1840 VP.n48 VP.n10 161.3
R1841 VP.n47 VP.n46 161.3
R1842 VP.n20 VP.t0 126.361
R1843 VP.n45 VP.n11 110.12
R1844 VP.n80 VP.n79 110.12
R1845 VP.n44 VP.n43 110.12
R1846 VP.n11 VP.t6 94.4789
R1847 VP.n7 VP.t3 94.4789
R1848 VP.n66 VP.t7 94.4789
R1849 VP.n79 VP.t1 94.4789
R1850 VP.n43 VP.t5 94.4789
R1851 VP.n30 VP.t2 94.4789
R1852 VP.n19 VP.t4 94.4789
R1853 VP.n20 VP.n19 65.4799
R1854 VP.n53 VP.n9 55.9904
R1855 VP.n73 VP.n72 55.9904
R1856 VP.n37 VP.n36 55.9904
R1857 VP.n45 VP.n44 52.6359
R1858 VP.n60 VP.n5 40.4106
R1859 VP.n64 VP.n5 40.4106
R1860 VP.n28 VP.n17 40.4106
R1861 VP.n24 VP.n17 40.4106
R1862 VP.n49 VP.n9 24.8308
R1863 VP.n73 VP.n1 24.8308
R1864 VP.n37 VP.n13 24.8308
R1865 VP.n48 VP.n47 24.3439
R1866 VP.n49 VP.n48 24.3439
R1867 VP.n54 VP.n53 24.3439
R1868 VP.n55 VP.n54 24.3439
R1869 VP.n59 VP.n58 24.3439
R1870 VP.n60 VP.n59 24.3439
R1871 VP.n65 VP.n64 24.3439
R1872 VP.n67 VP.n65 24.3439
R1873 VP.n71 VP.n3 24.3439
R1874 VP.n72 VP.n71 24.3439
R1875 VP.n77 VP.n1 24.3439
R1876 VP.n78 VP.n77 24.3439
R1877 VP.n41 VP.n13 24.3439
R1878 VP.n42 VP.n41 24.3439
R1879 VP.n29 VP.n28 24.3439
R1880 VP.n31 VP.n29 24.3439
R1881 VP.n35 VP.n15 24.3439
R1882 VP.n36 VP.n35 24.3439
R1883 VP.n23 VP.n22 24.3439
R1884 VP.n24 VP.n23 24.3439
R1885 VP.n55 VP.n7 16.0672
R1886 VP.n66 VP.n3 16.0672
R1887 VP.n30 VP.n15 16.0672
R1888 VP.n58 VP.n7 8.27727
R1889 VP.n67 VP.n66 8.27727
R1890 VP.n31 VP.n30 8.27727
R1891 VP.n22 VP.n19 8.27727
R1892 VP.n21 VP.n20 5.22731
R1893 VP.n47 VP.n11 0.487369
R1894 VP.n79 VP.n78 0.487369
R1895 VP.n43 VP.n42 0.487369
R1896 VP.n44 VP.n12 0.278398
R1897 VP.n46 VP.n45 0.278398
R1898 VP.n80 VP.n0 0.278398
R1899 VP.n21 VP.n18 0.189894
R1900 VP.n25 VP.n18 0.189894
R1901 VP.n26 VP.n25 0.189894
R1902 VP.n27 VP.n26 0.189894
R1903 VP.n27 VP.n16 0.189894
R1904 VP.n32 VP.n16 0.189894
R1905 VP.n33 VP.n32 0.189894
R1906 VP.n34 VP.n33 0.189894
R1907 VP.n34 VP.n14 0.189894
R1908 VP.n38 VP.n14 0.189894
R1909 VP.n39 VP.n38 0.189894
R1910 VP.n40 VP.n39 0.189894
R1911 VP.n40 VP.n12 0.189894
R1912 VP.n46 VP.n10 0.189894
R1913 VP.n50 VP.n10 0.189894
R1914 VP.n51 VP.n50 0.189894
R1915 VP.n52 VP.n51 0.189894
R1916 VP.n52 VP.n8 0.189894
R1917 VP.n56 VP.n8 0.189894
R1918 VP.n57 VP.n56 0.189894
R1919 VP.n57 VP.n6 0.189894
R1920 VP.n61 VP.n6 0.189894
R1921 VP.n62 VP.n61 0.189894
R1922 VP.n63 VP.n62 0.189894
R1923 VP.n63 VP.n4 0.189894
R1924 VP.n68 VP.n4 0.189894
R1925 VP.n69 VP.n68 0.189894
R1926 VP.n70 VP.n69 0.189894
R1927 VP.n70 VP.n2 0.189894
R1928 VP.n74 VP.n2 0.189894
R1929 VP.n75 VP.n74 0.189894
R1930 VP.n76 VP.n75 0.189894
R1931 VP.n76 VP.n0 0.189894
R1932 VP VP.n80 0.153422
R1933 VDD1 VDD1.n0 64.2536
R1934 VDD1.n3 VDD1.n2 64.1399
R1935 VDD1.n3 VDD1.n1 64.1399
R1936 VDD1.n5 VDD1.n4 62.7556
R1937 VDD1.n5 VDD1.n3 47.4276
R1938 VDD1.n4 VDD1.t2 1.67847
R1939 VDD1.n4 VDD1.t7 1.67847
R1940 VDD1.n0 VDD1.t5 1.67847
R1941 VDD1.n0 VDD1.t0 1.67847
R1942 VDD1.n2 VDD1.t3 1.67847
R1943 VDD1.n2 VDD1.t6 1.67847
R1944 VDD1.n1 VDD1.t4 1.67847
R1945 VDD1.n1 VDD1.t1 1.67847
R1946 VDD1 VDD1.n5 1.38197
R1947 VTAIL.n11 VTAIL.t15 47.755
R1948 VTAIL.n10 VTAIL.t0 47.755
R1949 VTAIL.n7 VTAIL.t1 47.755
R1950 VTAIL.n15 VTAIL.t7 47.7547
R1951 VTAIL.n2 VTAIL.t3 47.7547
R1952 VTAIL.n3 VTAIL.t14 47.7547
R1953 VTAIL.n6 VTAIL.t9 47.7547
R1954 VTAIL.n14 VTAIL.t10 47.7547
R1955 VTAIL.n13 VTAIL.n12 46.077
R1956 VTAIL.n9 VTAIL.n8 46.077
R1957 VTAIL.n1 VTAIL.n0 46.0768
R1958 VTAIL.n5 VTAIL.n4 46.0768
R1959 VTAIL.n15 VTAIL.n14 25.4186
R1960 VTAIL.n7 VTAIL.n6 25.4186
R1961 VTAIL.n9 VTAIL.n7 2.87981
R1962 VTAIL.n10 VTAIL.n9 2.87981
R1963 VTAIL.n13 VTAIL.n11 2.87981
R1964 VTAIL.n14 VTAIL.n13 2.87981
R1965 VTAIL.n6 VTAIL.n5 2.87981
R1966 VTAIL.n5 VTAIL.n3 2.87981
R1967 VTAIL.n2 VTAIL.n1 2.87981
R1968 VTAIL VTAIL.n15 2.82162
R1969 VTAIL.n0 VTAIL.t2 1.67847
R1970 VTAIL.n0 VTAIL.t6 1.67847
R1971 VTAIL.n4 VTAIL.t12 1.67847
R1972 VTAIL.n4 VTAIL.t8 1.67847
R1973 VTAIL.n12 VTAIL.t11 1.67847
R1974 VTAIL.n12 VTAIL.t13 1.67847
R1975 VTAIL.n8 VTAIL.t4 1.67847
R1976 VTAIL.n8 VTAIL.t5 1.67847
R1977 VTAIL.n11 VTAIL.n10 0.470328
R1978 VTAIL.n3 VTAIL.n2 0.470328
R1979 VTAIL VTAIL.n1 0.0586897
R1980 VN.n63 VN.n33 161.3
R1981 VN.n62 VN.n61 161.3
R1982 VN.n60 VN.n34 161.3
R1983 VN.n59 VN.n58 161.3
R1984 VN.n57 VN.n35 161.3
R1985 VN.n56 VN.n55 161.3
R1986 VN.n54 VN.n36 161.3
R1987 VN.n53 VN.n52 161.3
R1988 VN.n51 VN.n37 161.3
R1989 VN.n50 VN.n49 161.3
R1990 VN.n48 VN.n39 161.3
R1991 VN.n47 VN.n46 161.3
R1992 VN.n45 VN.n40 161.3
R1993 VN.n44 VN.n43 161.3
R1994 VN.n30 VN.n0 161.3
R1995 VN.n29 VN.n28 161.3
R1996 VN.n27 VN.n1 161.3
R1997 VN.n26 VN.n25 161.3
R1998 VN.n24 VN.n2 161.3
R1999 VN.n23 VN.n22 161.3
R2000 VN.n21 VN.n3 161.3
R2001 VN.n20 VN.n19 161.3
R2002 VN.n17 VN.n4 161.3
R2003 VN.n16 VN.n15 161.3
R2004 VN.n14 VN.n5 161.3
R2005 VN.n13 VN.n12 161.3
R2006 VN.n11 VN.n6 161.3
R2007 VN.n10 VN.n9 161.3
R2008 VN.n8 VN.t3 126.361
R2009 VN.n42 VN.t5 126.361
R2010 VN.n32 VN.n31 110.12
R2011 VN.n65 VN.n64 110.12
R2012 VN.n7 VN.t6 94.4789
R2013 VN.n18 VN.t4 94.4789
R2014 VN.n31 VN.t0 94.4789
R2015 VN.n41 VN.t7 94.4789
R2016 VN.n38 VN.t1 94.4789
R2017 VN.n64 VN.t2 94.4789
R2018 VN.n8 VN.n7 65.4799
R2019 VN.n42 VN.n41 65.4799
R2020 VN.n25 VN.n24 55.9904
R2021 VN.n58 VN.n57 55.9904
R2022 VN VN.n65 52.9148
R2023 VN.n12 VN.n5 40.4106
R2024 VN.n16 VN.n5 40.4106
R2025 VN.n46 VN.n39 40.4106
R2026 VN.n50 VN.n39 40.4106
R2027 VN.n25 VN.n1 24.8308
R2028 VN.n58 VN.n34 24.8308
R2029 VN.n11 VN.n10 24.3439
R2030 VN.n12 VN.n11 24.3439
R2031 VN.n17 VN.n16 24.3439
R2032 VN.n19 VN.n17 24.3439
R2033 VN.n23 VN.n3 24.3439
R2034 VN.n24 VN.n23 24.3439
R2035 VN.n29 VN.n1 24.3439
R2036 VN.n30 VN.n29 24.3439
R2037 VN.n46 VN.n45 24.3439
R2038 VN.n45 VN.n44 24.3439
R2039 VN.n57 VN.n56 24.3439
R2040 VN.n56 VN.n36 24.3439
R2041 VN.n52 VN.n51 24.3439
R2042 VN.n51 VN.n50 24.3439
R2043 VN.n63 VN.n62 24.3439
R2044 VN.n62 VN.n34 24.3439
R2045 VN.n18 VN.n3 16.0672
R2046 VN.n38 VN.n36 16.0672
R2047 VN.n10 VN.n7 8.27727
R2048 VN.n19 VN.n18 8.27727
R2049 VN.n44 VN.n41 8.27727
R2050 VN.n52 VN.n38 8.27727
R2051 VN.n43 VN.n42 5.22731
R2052 VN.n9 VN.n8 5.22731
R2053 VN.n31 VN.n30 0.487369
R2054 VN.n64 VN.n63 0.487369
R2055 VN.n65 VN.n33 0.278398
R2056 VN.n32 VN.n0 0.278398
R2057 VN.n61 VN.n33 0.189894
R2058 VN.n61 VN.n60 0.189894
R2059 VN.n60 VN.n59 0.189894
R2060 VN.n59 VN.n35 0.189894
R2061 VN.n55 VN.n35 0.189894
R2062 VN.n55 VN.n54 0.189894
R2063 VN.n54 VN.n53 0.189894
R2064 VN.n53 VN.n37 0.189894
R2065 VN.n49 VN.n37 0.189894
R2066 VN.n49 VN.n48 0.189894
R2067 VN.n48 VN.n47 0.189894
R2068 VN.n47 VN.n40 0.189894
R2069 VN.n43 VN.n40 0.189894
R2070 VN.n9 VN.n6 0.189894
R2071 VN.n13 VN.n6 0.189894
R2072 VN.n14 VN.n13 0.189894
R2073 VN.n15 VN.n14 0.189894
R2074 VN.n15 VN.n4 0.189894
R2075 VN.n20 VN.n4 0.189894
R2076 VN.n21 VN.n20 0.189894
R2077 VN.n22 VN.n21 0.189894
R2078 VN.n22 VN.n2 0.189894
R2079 VN.n26 VN.n2 0.189894
R2080 VN.n27 VN.n26 0.189894
R2081 VN.n28 VN.n27 0.189894
R2082 VN.n28 VN.n0 0.189894
R2083 VN VN.n32 0.153422
R2084 VDD2.n2 VDD2.n1 64.1399
R2085 VDD2.n2 VDD2.n0 64.1399
R2086 VDD2 VDD2.n5 64.1371
R2087 VDD2.n4 VDD2.n3 62.7558
R2088 VDD2.n4 VDD2.n2 46.8446
R2089 VDD2.n5 VDD2.t0 1.67847
R2090 VDD2.n5 VDD2.t2 1.67847
R2091 VDD2.n3 VDD2.t5 1.67847
R2092 VDD2.n3 VDD2.t6 1.67847
R2093 VDD2.n1 VDD2.t3 1.67847
R2094 VDD2.n1 VDD2.t7 1.67847
R2095 VDD2.n0 VDD2.t4 1.67847
R2096 VDD2.n0 VDD2.t1 1.67847
R2097 VDD2 VDD2.n4 1.49834
C0 VDD2 VP 0.563051f
C1 VN VDD2 8.78471f
C2 VN VP 8.13227f
C3 VTAIL VDD1 8.13451f
C4 VDD2 VDD1 1.99156f
C5 VDD1 VP 9.19393f
C6 VDD2 VTAIL 8.19168f
C7 VN VDD1 0.152221f
C8 VTAIL VP 9.351269f
C9 VN VTAIL 9.33716f
C10 VDD2 B 5.723052f
C11 VDD1 B 6.202721f
C12 VTAIL B 10.640762f
C13 VN B 17.054472f
C14 VP B 15.683986f
C15 VDD2.t4 B 0.225632f
C16 VDD2.t1 B 0.225632f
C17 VDD2.n0 B 2.0208f
C18 VDD2.t3 B 0.225632f
C19 VDD2.t7 B 0.225632f
C20 VDD2.n1 B 2.0208f
C21 VDD2.n2 B 3.39073f
C22 VDD2.t5 B 0.225632f
C23 VDD2.t6 B 0.225632f
C24 VDD2.n3 B 2.0091f
C25 VDD2.n4 B 2.97857f
C26 VDD2.t0 B 0.225632f
C27 VDD2.t2 B 0.225632f
C28 VDD2.n5 B 2.02076f
C29 VN.n0 B 0.026585f
C30 VN.t0 B 1.95036f
C31 VN.n1 B 0.038127f
C32 VN.n2 B 0.020164f
C33 VN.n3 B 0.031428f
C34 VN.n4 B 0.020164f
C35 VN.n5 B 0.016317f
C36 VN.n6 B 0.020164f
C37 VN.t6 B 1.95036f
C38 VN.n7 B 0.749575f
C39 VN.t3 B 2.15934f
C40 VN.n8 B 0.726808f
C41 VN.n9 B 0.216475f
C42 VN.n10 B 0.025461f
C43 VN.n11 B 0.037768f
C44 VN.n12 B 0.040289f
C45 VN.n13 B 0.020164f
C46 VN.n14 B 0.020164f
C47 VN.n15 B 0.020164f
C48 VN.n16 B 0.040289f
C49 VN.n17 B 0.037768f
C50 VN.t4 B 1.95036f
C51 VN.n18 B 0.687665f
C52 VN.n19 B 0.025461f
C53 VN.n20 B 0.020164f
C54 VN.n21 B 0.020164f
C55 VN.n22 B 0.020164f
C56 VN.n23 B 0.037768f
C57 VN.n24 B 0.034606f
C58 VN.n25 B 0.024162f
C59 VN.n26 B 0.020164f
C60 VN.n27 B 0.020164f
C61 VN.n28 B 0.020164f
C62 VN.n29 B 0.037768f
C63 VN.n30 B 0.019494f
C64 VN.n31 B 0.756119f
C65 VN.n32 B 0.040422f
C66 VN.n33 B 0.026585f
C67 VN.t2 B 1.95036f
C68 VN.n34 B 0.038127f
C69 VN.n35 B 0.020164f
C70 VN.n36 B 0.031428f
C71 VN.n37 B 0.020164f
C72 VN.t1 B 1.95036f
C73 VN.n38 B 0.687665f
C74 VN.n39 B 0.016317f
C75 VN.n40 B 0.020164f
C76 VN.t7 B 1.95036f
C77 VN.n41 B 0.749575f
C78 VN.t5 B 2.15934f
C79 VN.n42 B 0.726808f
C80 VN.n43 B 0.216475f
C81 VN.n44 B 0.025461f
C82 VN.n45 B 0.037768f
C83 VN.n46 B 0.040289f
C84 VN.n47 B 0.020164f
C85 VN.n48 B 0.020164f
C86 VN.n49 B 0.020164f
C87 VN.n50 B 0.040289f
C88 VN.n51 B 0.037768f
C89 VN.n52 B 0.025461f
C90 VN.n53 B 0.020164f
C91 VN.n54 B 0.020164f
C92 VN.n55 B 0.020164f
C93 VN.n56 B 0.037768f
C94 VN.n57 B 0.034606f
C95 VN.n58 B 0.024162f
C96 VN.n59 B 0.020164f
C97 VN.n60 B 0.020164f
C98 VN.n61 B 0.020164f
C99 VN.n62 B 0.037768f
C100 VN.n63 B 0.019494f
C101 VN.n64 B 0.756119f
C102 VN.n65 B 1.22741f
C103 VTAIL.t2 B 0.188211f
C104 VTAIL.t6 B 0.188211f
C105 VTAIL.n0 B 1.61707f
C106 VTAIL.n1 B 0.388758f
C107 VTAIL.t3 B 2.06213f
C108 VTAIL.n2 B 0.483773f
C109 VTAIL.t14 B 2.06213f
C110 VTAIL.n3 B 0.483773f
C111 VTAIL.t12 B 0.188211f
C112 VTAIL.t8 B 0.188211f
C113 VTAIL.n4 B 1.61707f
C114 VTAIL.n5 B 0.572237f
C115 VTAIL.t9 B 2.06213f
C116 VTAIL.n6 B 1.57625f
C117 VTAIL.t1 B 2.06213f
C118 VTAIL.n7 B 1.57624f
C119 VTAIL.t4 B 0.188211f
C120 VTAIL.t5 B 0.188211f
C121 VTAIL.n8 B 1.61707f
C122 VTAIL.n9 B 0.572232f
C123 VTAIL.t0 B 2.06213f
C124 VTAIL.n10 B 0.483768f
C125 VTAIL.t15 B 2.06213f
C126 VTAIL.n11 B 0.483768f
C127 VTAIL.t11 B 0.188211f
C128 VTAIL.t13 B 0.188211f
C129 VTAIL.n12 B 1.61707f
C130 VTAIL.n13 B 0.572232f
C131 VTAIL.t10 B 2.06213f
C132 VTAIL.n14 B 1.57625f
C133 VTAIL.t7 B 2.06213f
C134 VTAIL.n15 B 1.57246f
C135 VDD1.t5 B 0.228413f
C136 VDD1.t0 B 0.228413f
C137 VDD1.n0 B 2.04685f
C138 VDD1.t4 B 0.228413f
C139 VDD1.t1 B 0.228413f
C140 VDD1.n1 B 2.0457f
C141 VDD1.t3 B 0.228413f
C142 VDD1.t6 B 0.228413f
C143 VDD1.n2 B 2.0457f
C144 VDD1.n3 B 3.48333f
C145 VDD1.t2 B 0.228413f
C146 VDD1.t7 B 0.228413f
C147 VDD1.n4 B 2.03386f
C148 VDD1.n5 B 3.04577f
C149 VP.n0 B 0.027122f
C150 VP.t1 B 1.98973f
C151 VP.n1 B 0.038896f
C152 VP.n2 B 0.020571f
C153 VP.n3 B 0.032063f
C154 VP.n4 B 0.020571f
C155 VP.n5 B 0.016646f
C156 VP.n6 B 0.020571f
C157 VP.t3 B 1.98973f
C158 VP.n7 B 0.701547f
C159 VP.n8 B 0.020571f
C160 VP.n9 B 0.02465f
C161 VP.n10 B 0.020571f
C162 VP.t6 B 1.98973f
C163 VP.n11 B 0.771383f
C164 VP.n12 B 0.027122f
C165 VP.t5 B 1.98973f
C166 VP.n13 B 0.038896f
C167 VP.n14 B 0.020571f
C168 VP.n15 B 0.032063f
C169 VP.n16 B 0.020571f
C170 VP.n17 B 0.016646f
C171 VP.n18 B 0.020571f
C172 VP.t4 B 1.98973f
C173 VP.n19 B 0.764707f
C174 VP.t0 B 2.20293f
C175 VP.n20 B 0.74148f
C176 VP.n21 B 0.220845f
C177 VP.n22 B 0.025975f
C178 VP.n23 B 0.038531f
C179 VP.n24 B 0.041103f
C180 VP.n25 B 0.020571f
C181 VP.n26 B 0.020571f
C182 VP.n27 B 0.020571f
C183 VP.n28 B 0.041103f
C184 VP.n29 B 0.038531f
C185 VP.t2 B 1.98973f
C186 VP.n30 B 0.701547f
C187 VP.n31 B 0.025975f
C188 VP.n32 B 0.020571f
C189 VP.n33 B 0.020571f
C190 VP.n34 B 0.020571f
C191 VP.n35 B 0.038531f
C192 VP.n36 B 0.035305f
C193 VP.n37 B 0.02465f
C194 VP.n38 B 0.020571f
C195 VP.n39 B 0.020571f
C196 VP.n40 B 0.020571f
C197 VP.n41 B 0.038531f
C198 VP.n42 B 0.019887f
C199 VP.n43 B 0.771383f
C200 VP.n44 B 1.24122f
C201 VP.n45 B 1.25523f
C202 VP.n46 B 0.027122f
C203 VP.n47 B 0.019887f
C204 VP.n48 B 0.038531f
C205 VP.n49 B 0.038896f
C206 VP.n50 B 0.020571f
C207 VP.n51 B 0.020571f
C208 VP.n52 B 0.020571f
C209 VP.n53 B 0.035305f
C210 VP.n54 B 0.038531f
C211 VP.n55 B 0.032063f
C212 VP.n56 B 0.020571f
C213 VP.n57 B 0.020571f
C214 VP.n58 B 0.025975f
C215 VP.n59 B 0.038531f
C216 VP.n60 B 0.041103f
C217 VP.n61 B 0.020571f
C218 VP.n62 B 0.020571f
C219 VP.n63 B 0.020571f
C220 VP.n64 B 0.041103f
C221 VP.n65 B 0.038531f
C222 VP.t7 B 1.98973f
C223 VP.n66 B 0.701547f
C224 VP.n67 B 0.025975f
C225 VP.n68 B 0.020571f
C226 VP.n69 B 0.020571f
C227 VP.n70 B 0.020571f
C228 VP.n71 B 0.038531f
C229 VP.n72 B 0.035305f
C230 VP.n73 B 0.02465f
C231 VP.n74 B 0.020571f
C232 VP.n75 B 0.020571f
C233 VP.n76 B 0.020571f
C234 VP.n77 B 0.038531f
C235 VP.n78 B 0.019887f
C236 VP.n79 B 0.771383f
C237 VP.n80 B 0.041238f
.ends

