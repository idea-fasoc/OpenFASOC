* NGSPICE file created from diff_pair_sample_1632.ext - technology: sky130A

.subckt diff_pair_sample_1632 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=1.86
X1 VDD1.t9 VP.t0 VTAIL.t13 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X2 VTAIL.t8 VN.t0 VDD2.t9 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X3 VDD1.t8 VP.t1 VTAIL.t11 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X4 B.t8 B.t6 B.t7 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=1.86
X5 VDD1.t7 VP.t2 VTAIL.t15 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=1.86
X6 VDD2.t8 VN.t1 VTAIL.t1 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=1.86
X7 VDD1.t6 VP.t3 VTAIL.t16 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=1.86
X8 B.t5 B.t3 B.t4 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=1.86
X9 VTAIL.t14 VP.t4 VDD1.t5 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X10 VDD2.t7 VN.t2 VTAIL.t7 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=1.86
X11 VTAIL.t12 VP.t5 VDD1.t4 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X12 B.t2 B.t0 B.t1 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=1.86
X13 VTAIL.t4 VN.t3 VDD2.t6 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X14 VDD2.t5 VN.t4 VTAIL.t3 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=1.86
X15 VTAIL.t6 VN.t5 VDD2.t4 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X16 VDD1.t3 VP.t6 VTAIL.t17 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=1.86
X17 VTAIL.t10 VP.t7 VDD1.t2 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X18 VDD2.t3 VN.t6 VTAIL.t9 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X19 VTAIL.t19 VP.t8 VDD1.t1 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X20 VDD2.t2 VN.t7 VTAIL.t5 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=1.86
X21 VTAIL.t0 VN.t8 VDD2.t1 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
X22 VDD1.t0 VP.t9 VTAIL.t18 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=1.86
X23 VDD2.t0 VN.t9 VTAIL.t2 w_n3598_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=1.86
R0 B.n387 B.n386 585
R1 B.n385 B.n120 585
R2 B.n384 B.n383 585
R3 B.n382 B.n121 585
R4 B.n381 B.n380 585
R5 B.n379 B.n122 585
R6 B.n378 B.n377 585
R7 B.n376 B.n123 585
R8 B.n375 B.n374 585
R9 B.n373 B.n124 585
R10 B.n372 B.n371 585
R11 B.n370 B.n125 585
R12 B.n369 B.n368 585
R13 B.n367 B.n126 585
R14 B.n366 B.n365 585
R15 B.n364 B.n127 585
R16 B.n363 B.n362 585
R17 B.n361 B.n128 585
R18 B.n360 B.n359 585
R19 B.n358 B.n129 585
R20 B.n357 B.n356 585
R21 B.n355 B.n130 585
R22 B.n354 B.n353 585
R23 B.n352 B.n131 585
R24 B.n351 B.n350 585
R25 B.n349 B.n132 585
R26 B.n348 B.n347 585
R27 B.n346 B.n133 585
R28 B.n345 B.n344 585
R29 B.n343 B.n134 585
R30 B.n342 B.n341 585
R31 B.n340 B.n135 585
R32 B.n339 B.n338 585
R33 B.n337 B.n136 585
R34 B.n336 B.n335 585
R35 B.n334 B.n137 585
R36 B.n333 B.n332 585
R37 B.n331 B.n138 585
R38 B.n330 B.n329 585
R39 B.n325 B.n139 585
R40 B.n324 B.n323 585
R41 B.n322 B.n140 585
R42 B.n321 B.n320 585
R43 B.n319 B.n141 585
R44 B.n318 B.n317 585
R45 B.n316 B.n142 585
R46 B.n315 B.n314 585
R47 B.n313 B.n143 585
R48 B.n311 B.n310 585
R49 B.n309 B.n146 585
R50 B.n308 B.n307 585
R51 B.n306 B.n147 585
R52 B.n305 B.n304 585
R53 B.n303 B.n148 585
R54 B.n302 B.n301 585
R55 B.n300 B.n149 585
R56 B.n299 B.n298 585
R57 B.n297 B.n150 585
R58 B.n296 B.n295 585
R59 B.n294 B.n151 585
R60 B.n293 B.n292 585
R61 B.n291 B.n152 585
R62 B.n290 B.n289 585
R63 B.n288 B.n153 585
R64 B.n287 B.n286 585
R65 B.n285 B.n154 585
R66 B.n284 B.n283 585
R67 B.n282 B.n155 585
R68 B.n281 B.n280 585
R69 B.n279 B.n156 585
R70 B.n278 B.n277 585
R71 B.n276 B.n157 585
R72 B.n275 B.n274 585
R73 B.n273 B.n158 585
R74 B.n272 B.n271 585
R75 B.n270 B.n159 585
R76 B.n269 B.n268 585
R77 B.n267 B.n160 585
R78 B.n266 B.n265 585
R79 B.n264 B.n161 585
R80 B.n263 B.n262 585
R81 B.n261 B.n162 585
R82 B.n260 B.n259 585
R83 B.n258 B.n163 585
R84 B.n257 B.n256 585
R85 B.n255 B.n164 585
R86 B.n388 B.n119 585
R87 B.n390 B.n389 585
R88 B.n391 B.n118 585
R89 B.n393 B.n392 585
R90 B.n394 B.n117 585
R91 B.n396 B.n395 585
R92 B.n397 B.n116 585
R93 B.n399 B.n398 585
R94 B.n400 B.n115 585
R95 B.n402 B.n401 585
R96 B.n403 B.n114 585
R97 B.n405 B.n404 585
R98 B.n406 B.n113 585
R99 B.n408 B.n407 585
R100 B.n409 B.n112 585
R101 B.n411 B.n410 585
R102 B.n412 B.n111 585
R103 B.n414 B.n413 585
R104 B.n415 B.n110 585
R105 B.n417 B.n416 585
R106 B.n418 B.n109 585
R107 B.n420 B.n419 585
R108 B.n421 B.n108 585
R109 B.n423 B.n422 585
R110 B.n424 B.n107 585
R111 B.n426 B.n425 585
R112 B.n427 B.n106 585
R113 B.n429 B.n428 585
R114 B.n430 B.n105 585
R115 B.n432 B.n431 585
R116 B.n433 B.n104 585
R117 B.n435 B.n434 585
R118 B.n436 B.n103 585
R119 B.n438 B.n437 585
R120 B.n439 B.n102 585
R121 B.n441 B.n440 585
R122 B.n442 B.n101 585
R123 B.n444 B.n443 585
R124 B.n445 B.n100 585
R125 B.n447 B.n446 585
R126 B.n448 B.n99 585
R127 B.n450 B.n449 585
R128 B.n451 B.n98 585
R129 B.n453 B.n452 585
R130 B.n454 B.n97 585
R131 B.n456 B.n455 585
R132 B.n457 B.n96 585
R133 B.n459 B.n458 585
R134 B.n460 B.n95 585
R135 B.n462 B.n461 585
R136 B.n463 B.n94 585
R137 B.n465 B.n464 585
R138 B.n466 B.n93 585
R139 B.n468 B.n467 585
R140 B.n469 B.n92 585
R141 B.n471 B.n470 585
R142 B.n472 B.n91 585
R143 B.n474 B.n473 585
R144 B.n475 B.n90 585
R145 B.n477 B.n476 585
R146 B.n478 B.n89 585
R147 B.n480 B.n479 585
R148 B.n481 B.n88 585
R149 B.n483 B.n482 585
R150 B.n484 B.n87 585
R151 B.n486 B.n485 585
R152 B.n487 B.n86 585
R153 B.n489 B.n488 585
R154 B.n490 B.n85 585
R155 B.n492 B.n491 585
R156 B.n493 B.n84 585
R157 B.n495 B.n494 585
R158 B.n496 B.n83 585
R159 B.n498 B.n497 585
R160 B.n499 B.n82 585
R161 B.n501 B.n500 585
R162 B.n502 B.n81 585
R163 B.n504 B.n503 585
R164 B.n505 B.n80 585
R165 B.n507 B.n506 585
R166 B.n508 B.n79 585
R167 B.n510 B.n509 585
R168 B.n511 B.n78 585
R169 B.n513 B.n512 585
R170 B.n514 B.n77 585
R171 B.n516 B.n515 585
R172 B.n517 B.n76 585
R173 B.n519 B.n518 585
R174 B.n520 B.n75 585
R175 B.n522 B.n521 585
R176 B.n523 B.n74 585
R177 B.n525 B.n524 585
R178 B.n526 B.n73 585
R179 B.n528 B.n527 585
R180 B.n658 B.n25 585
R181 B.n657 B.n656 585
R182 B.n655 B.n26 585
R183 B.n654 B.n653 585
R184 B.n652 B.n27 585
R185 B.n651 B.n650 585
R186 B.n649 B.n28 585
R187 B.n648 B.n647 585
R188 B.n646 B.n29 585
R189 B.n645 B.n644 585
R190 B.n643 B.n30 585
R191 B.n642 B.n641 585
R192 B.n640 B.n31 585
R193 B.n639 B.n638 585
R194 B.n637 B.n32 585
R195 B.n636 B.n635 585
R196 B.n634 B.n33 585
R197 B.n633 B.n632 585
R198 B.n631 B.n34 585
R199 B.n630 B.n629 585
R200 B.n628 B.n35 585
R201 B.n627 B.n626 585
R202 B.n625 B.n36 585
R203 B.n624 B.n623 585
R204 B.n622 B.n37 585
R205 B.n621 B.n620 585
R206 B.n619 B.n38 585
R207 B.n618 B.n617 585
R208 B.n616 B.n39 585
R209 B.n615 B.n614 585
R210 B.n613 B.n40 585
R211 B.n612 B.n611 585
R212 B.n610 B.n41 585
R213 B.n609 B.n608 585
R214 B.n607 B.n42 585
R215 B.n606 B.n605 585
R216 B.n604 B.n43 585
R217 B.n603 B.n602 585
R218 B.n601 B.n600 585
R219 B.n599 B.n47 585
R220 B.n598 B.n597 585
R221 B.n596 B.n48 585
R222 B.n595 B.n594 585
R223 B.n593 B.n49 585
R224 B.n592 B.n591 585
R225 B.n590 B.n50 585
R226 B.n589 B.n588 585
R227 B.n587 B.n51 585
R228 B.n585 B.n584 585
R229 B.n583 B.n54 585
R230 B.n582 B.n581 585
R231 B.n580 B.n55 585
R232 B.n579 B.n578 585
R233 B.n577 B.n56 585
R234 B.n576 B.n575 585
R235 B.n574 B.n57 585
R236 B.n573 B.n572 585
R237 B.n571 B.n58 585
R238 B.n570 B.n569 585
R239 B.n568 B.n59 585
R240 B.n567 B.n566 585
R241 B.n565 B.n60 585
R242 B.n564 B.n563 585
R243 B.n562 B.n61 585
R244 B.n561 B.n560 585
R245 B.n559 B.n62 585
R246 B.n558 B.n557 585
R247 B.n556 B.n63 585
R248 B.n555 B.n554 585
R249 B.n553 B.n64 585
R250 B.n552 B.n551 585
R251 B.n550 B.n65 585
R252 B.n549 B.n548 585
R253 B.n547 B.n66 585
R254 B.n546 B.n545 585
R255 B.n544 B.n67 585
R256 B.n543 B.n542 585
R257 B.n541 B.n68 585
R258 B.n540 B.n539 585
R259 B.n538 B.n69 585
R260 B.n537 B.n536 585
R261 B.n535 B.n70 585
R262 B.n534 B.n533 585
R263 B.n532 B.n71 585
R264 B.n531 B.n530 585
R265 B.n529 B.n72 585
R266 B.n660 B.n659 585
R267 B.n661 B.n24 585
R268 B.n663 B.n662 585
R269 B.n664 B.n23 585
R270 B.n666 B.n665 585
R271 B.n667 B.n22 585
R272 B.n669 B.n668 585
R273 B.n670 B.n21 585
R274 B.n672 B.n671 585
R275 B.n673 B.n20 585
R276 B.n675 B.n674 585
R277 B.n676 B.n19 585
R278 B.n678 B.n677 585
R279 B.n679 B.n18 585
R280 B.n681 B.n680 585
R281 B.n682 B.n17 585
R282 B.n684 B.n683 585
R283 B.n685 B.n16 585
R284 B.n687 B.n686 585
R285 B.n688 B.n15 585
R286 B.n690 B.n689 585
R287 B.n691 B.n14 585
R288 B.n693 B.n692 585
R289 B.n694 B.n13 585
R290 B.n696 B.n695 585
R291 B.n697 B.n12 585
R292 B.n699 B.n698 585
R293 B.n700 B.n11 585
R294 B.n702 B.n701 585
R295 B.n703 B.n10 585
R296 B.n705 B.n704 585
R297 B.n706 B.n9 585
R298 B.n708 B.n707 585
R299 B.n709 B.n8 585
R300 B.n711 B.n710 585
R301 B.n712 B.n7 585
R302 B.n714 B.n713 585
R303 B.n715 B.n6 585
R304 B.n717 B.n716 585
R305 B.n718 B.n5 585
R306 B.n720 B.n719 585
R307 B.n721 B.n4 585
R308 B.n723 B.n722 585
R309 B.n724 B.n3 585
R310 B.n726 B.n725 585
R311 B.n727 B.n0 585
R312 B.n2 B.n1 585
R313 B.n188 B.n187 585
R314 B.n189 B.n186 585
R315 B.n191 B.n190 585
R316 B.n192 B.n185 585
R317 B.n194 B.n193 585
R318 B.n195 B.n184 585
R319 B.n197 B.n196 585
R320 B.n198 B.n183 585
R321 B.n200 B.n199 585
R322 B.n201 B.n182 585
R323 B.n203 B.n202 585
R324 B.n204 B.n181 585
R325 B.n206 B.n205 585
R326 B.n207 B.n180 585
R327 B.n209 B.n208 585
R328 B.n210 B.n179 585
R329 B.n212 B.n211 585
R330 B.n213 B.n178 585
R331 B.n215 B.n214 585
R332 B.n216 B.n177 585
R333 B.n218 B.n217 585
R334 B.n219 B.n176 585
R335 B.n221 B.n220 585
R336 B.n222 B.n175 585
R337 B.n224 B.n223 585
R338 B.n225 B.n174 585
R339 B.n227 B.n226 585
R340 B.n228 B.n173 585
R341 B.n230 B.n229 585
R342 B.n231 B.n172 585
R343 B.n233 B.n232 585
R344 B.n234 B.n171 585
R345 B.n236 B.n235 585
R346 B.n237 B.n170 585
R347 B.n239 B.n238 585
R348 B.n240 B.n169 585
R349 B.n242 B.n241 585
R350 B.n243 B.n168 585
R351 B.n245 B.n244 585
R352 B.n246 B.n167 585
R353 B.n248 B.n247 585
R354 B.n249 B.n166 585
R355 B.n251 B.n250 585
R356 B.n252 B.n165 585
R357 B.n254 B.n253 585
R358 B.n255 B.n254 530.939
R359 B.n386 B.n119 530.939
R360 B.n529 B.n528 530.939
R361 B.n660 B.n25 530.939
R362 B.n326 B.t4 397.005
R363 B.n52 B.t11 397.005
R364 B.n144 B.t7 397.005
R365 B.n44 B.t2 397.005
R366 B.n327 B.t5 354.531
R367 B.n53 B.t10 354.531
R368 B.n145 B.t8 354.531
R369 B.n45 B.t1 354.531
R370 B.n144 B.t6 346.764
R371 B.n326 B.t3 346.764
R372 B.n52 B.t9 346.764
R373 B.n44 B.t0 346.764
R374 B.n729 B.n728 256.663
R375 B.n728 B.n727 235.042
R376 B.n728 B.n2 235.042
R377 B.n256 B.n255 163.367
R378 B.n256 B.n163 163.367
R379 B.n260 B.n163 163.367
R380 B.n261 B.n260 163.367
R381 B.n262 B.n261 163.367
R382 B.n262 B.n161 163.367
R383 B.n266 B.n161 163.367
R384 B.n267 B.n266 163.367
R385 B.n268 B.n267 163.367
R386 B.n268 B.n159 163.367
R387 B.n272 B.n159 163.367
R388 B.n273 B.n272 163.367
R389 B.n274 B.n273 163.367
R390 B.n274 B.n157 163.367
R391 B.n278 B.n157 163.367
R392 B.n279 B.n278 163.367
R393 B.n280 B.n279 163.367
R394 B.n280 B.n155 163.367
R395 B.n284 B.n155 163.367
R396 B.n285 B.n284 163.367
R397 B.n286 B.n285 163.367
R398 B.n286 B.n153 163.367
R399 B.n290 B.n153 163.367
R400 B.n291 B.n290 163.367
R401 B.n292 B.n291 163.367
R402 B.n292 B.n151 163.367
R403 B.n296 B.n151 163.367
R404 B.n297 B.n296 163.367
R405 B.n298 B.n297 163.367
R406 B.n298 B.n149 163.367
R407 B.n302 B.n149 163.367
R408 B.n303 B.n302 163.367
R409 B.n304 B.n303 163.367
R410 B.n304 B.n147 163.367
R411 B.n308 B.n147 163.367
R412 B.n309 B.n308 163.367
R413 B.n310 B.n309 163.367
R414 B.n310 B.n143 163.367
R415 B.n315 B.n143 163.367
R416 B.n316 B.n315 163.367
R417 B.n317 B.n316 163.367
R418 B.n317 B.n141 163.367
R419 B.n321 B.n141 163.367
R420 B.n322 B.n321 163.367
R421 B.n323 B.n322 163.367
R422 B.n323 B.n139 163.367
R423 B.n330 B.n139 163.367
R424 B.n331 B.n330 163.367
R425 B.n332 B.n331 163.367
R426 B.n332 B.n137 163.367
R427 B.n336 B.n137 163.367
R428 B.n337 B.n336 163.367
R429 B.n338 B.n337 163.367
R430 B.n338 B.n135 163.367
R431 B.n342 B.n135 163.367
R432 B.n343 B.n342 163.367
R433 B.n344 B.n343 163.367
R434 B.n344 B.n133 163.367
R435 B.n348 B.n133 163.367
R436 B.n349 B.n348 163.367
R437 B.n350 B.n349 163.367
R438 B.n350 B.n131 163.367
R439 B.n354 B.n131 163.367
R440 B.n355 B.n354 163.367
R441 B.n356 B.n355 163.367
R442 B.n356 B.n129 163.367
R443 B.n360 B.n129 163.367
R444 B.n361 B.n360 163.367
R445 B.n362 B.n361 163.367
R446 B.n362 B.n127 163.367
R447 B.n366 B.n127 163.367
R448 B.n367 B.n366 163.367
R449 B.n368 B.n367 163.367
R450 B.n368 B.n125 163.367
R451 B.n372 B.n125 163.367
R452 B.n373 B.n372 163.367
R453 B.n374 B.n373 163.367
R454 B.n374 B.n123 163.367
R455 B.n378 B.n123 163.367
R456 B.n379 B.n378 163.367
R457 B.n380 B.n379 163.367
R458 B.n380 B.n121 163.367
R459 B.n384 B.n121 163.367
R460 B.n385 B.n384 163.367
R461 B.n386 B.n385 163.367
R462 B.n528 B.n73 163.367
R463 B.n524 B.n73 163.367
R464 B.n524 B.n523 163.367
R465 B.n523 B.n522 163.367
R466 B.n522 B.n75 163.367
R467 B.n518 B.n75 163.367
R468 B.n518 B.n517 163.367
R469 B.n517 B.n516 163.367
R470 B.n516 B.n77 163.367
R471 B.n512 B.n77 163.367
R472 B.n512 B.n511 163.367
R473 B.n511 B.n510 163.367
R474 B.n510 B.n79 163.367
R475 B.n506 B.n79 163.367
R476 B.n506 B.n505 163.367
R477 B.n505 B.n504 163.367
R478 B.n504 B.n81 163.367
R479 B.n500 B.n81 163.367
R480 B.n500 B.n499 163.367
R481 B.n499 B.n498 163.367
R482 B.n498 B.n83 163.367
R483 B.n494 B.n83 163.367
R484 B.n494 B.n493 163.367
R485 B.n493 B.n492 163.367
R486 B.n492 B.n85 163.367
R487 B.n488 B.n85 163.367
R488 B.n488 B.n487 163.367
R489 B.n487 B.n486 163.367
R490 B.n486 B.n87 163.367
R491 B.n482 B.n87 163.367
R492 B.n482 B.n481 163.367
R493 B.n481 B.n480 163.367
R494 B.n480 B.n89 163.367
R495 B.n476 B.n89 163.367
R496 B.n476 B.n475 163.367
R497 B.n475 B.n474 163.367
R498 B.n474 B.n91 163.367
R499 B.n470 B.n91 163.367
R500 B.n470 B.n469 163.367
R501 B.n469 B.n468 163.367
R502 B.n468 B.n93 163.367
R503 B.n464 B.n93 163.367
R504 B.n464 B.n463 163.367
R505 B.n463 B.n462 163.367
R506 B.n462 B.n95 163.367
R507 B.n458 B.n95 163.367
R508 B.n458 B.n457 163.367
R509 B.n457 B.n456 163.367
R510 B.n456 B.n97 163.367
R511 B.n452 B.n97 163.367
R512 B.n452 B.n451 163.367
R513 B.n451 B.n450 163.367
R514 B.n450 B.n99 163.367
R515 B.n446 B.n99 163.367
R516 B.n446 B.n445 163.367
R517 B.n445 B.n444 163.367
R518 B.n444 B.n101 163.367
R519 B.n440 B.n101 163.367
R520 B.n440 B.n439 163.367
R521 B.n439 B.n438 163.367
R522 B.n438 B.n103 163.367
R523 B.n434 B.n103 163.367
R524 B.n434 B.n433 163.367
R525 B.n433 B.n432 163.367
R526 B.n432 B.n105 163.367
R527 B.n428 B.n105 163.367
R528 B.n428 B.n427 163.367
R529 B.n427 B.n426 163.367
R530 B.n426 B.n107 163.367
R531 B.n422 B.n107 163.367
R532 B.n422 B.n421 163.367
R533 B.n421 B.n420 163.367
R534 B.n420 B.n109 163.367
R535 B.n416 B.n109 163.367
R536 B.n416 B.n415 163.367
R537 B.n415 B.n414 163.367
R538 B.n414 B.n111 163.367
R539 B.n410 B.n111 163.367
R540 B.n410 B.n409 163.367
R541 B.n409 B.n408 163.367
R542 B.n408 B.n113 163.367
R543 B.n404 B.n113 163.367
R544 B.n404 B.n403 163.367
R545 B.n403 B.n402 163.367
R546 B.n402 B.n115 163.367
R547 B.n398 B.n115 163.367
R548 B.n398 B.n397 163.367
R549 B.n397 B.n396 163.367
R550 B.n396 B.n117 163.367
R551 B.n392 B.n117 163.367
R552 B.n392 B.n391 163.367
R553 B.n391 B.n390 163.367
R554 B.n390 B.n119 163.367
R555 B.n656 B.n25 163.367
R556 B.n656 B.n655 163.367
R557 B.n655 B.n654 163.367
R558 B.n654 B.n27 163.367
R559 B.n650 B.n27 163.367
R560 B.n650 B.n649 163.367
R561 B.n649 B.n648 163.367
R562 B.n648 B.n29 163.367
R563 B.n644 B.n29 163.367
R564 B.n644 B.n643 163.367
R565 B.n643 B.n642 163.367
R566 B.n642 B.n31 163.367
R567 B.n638 B.n31 163.367
R568 B.n638 B.n637 163.367
R569 B.n637 B.n636 163.367
R570 B.n636 B.n33 163.367
R571 B.n632 B.n33 163.367
R572 B.n632 B.n631 163.367
R573 B.n631 B.n630 163.367
R574 B.n630 B.n35 163.367
R575 B.n626 B.n35 163.367
R576 B.n626 B.n625 163.367
R577 B.n625 B.n624 163.367
R578 B.n624 B.n37 163.367
R579 B.n620 B.n37 163.367
R580 B.n620 B.n619 163.367
R581 B.n619 B.n618 163.367
R582 B.n618 B.n39 163.367
R583 B.n614 B.n39 163.367
R584 B.n614 B.n613 163.367
R585 B.n613 B.n612 163.367
R586 B.n612 B.n41 163.367
R587 B.n608 B.n41 163.367
R588 B.n608 B.n607 163.367
R589 B.n607 B.n606 163.367
R590 B.n606 B.n43 163.367
R591 B.n602 B.n43 163.367
R592 B.n602 B.n601 163.367
R593 B.n601 B.n47 163.367
R594 B.n597 B.n47 163.367
R595 B.n597 B.n596 163.367
R596 B.n596 B.n595 163.367
R597 B.n595 B.n49 163.367
R598 B.n591 B.n49 163.367
R599 B.n591 B.n590 163.367
R600 B.n590 B.n589 163.367
R601 B.n589 B.n51 163.367
R602 B.n584 B.n51 163.367
R603 B.n584 B.n583 163.367
R604 B.n583 B.n582 163.367
R605 B.n582 B.n55 163.367
R606 B.n578 B.n55 163.367
R607 B.n578 B.n577 163.367
R608 B.n577 B.n576 163.367
R609 B.n576 B.n57 163.367
R610 B.n572 B.n57 163.367
R611 B.n572 B.n571 163.367
R612 B.n571 B.n570 163.367
R613 B.n570 B.n59 163.367
R614 B.n566 B.n59 163.367
R615 B.n566 B.n565 163.367
R616 B.n565 B.n564 163.367
R617 B.n564 B.n61 163.367
R618 B.n560 B.n61 163.367
R619 B.n560 B.n559 163.367
R620 B.n559 B.n558 163.367
R621 B.n558 B.n63 163.367
R622 B.n554 B.n63 163.367
R623 B.n554 B.n553 163.367
R624 B.n553 B.n552 163.367
R625 B.n552 B.n65 163.367
R626 B.n548 B.n65 163.367
R627 B.n548 B.n547 163.367
R628 B.n547 B.n546 163.367
R629 B.n546 B.n67 163.367
R630 B.n542 B.n67 163.367
R631 B.n542 B.n541 163.367
R632 B.n541 B.n540 163.367
R633 B.n540 B.n69 163.367
R634 B.n536 B.n69 163.367
R635 B.n536 B.n535 163.367
R636 B.n535 B.n534 163.367
R637 B.n534 B.n71 163.367
R638 B.n530 B.n71 163.367
R639 B.n530 B.n529 163.367
R640 B.n661 B.n660 163.367
R641 B.n662 B.n661 163.367
R642 B.n662 B.n23 163.367
R643 B.n666 B.n23 163.367
R644 B.n667 B.n666 163.367
R645 B.n668 B.n667 163.367
R646 B.n668 B.n21 163.367
R647 B.n672 B.n21 163.367
R648 B.n673 B.n672 163.367
R649 B.n674 B.n673 163.367
R650 B.n674 B.n19 163.367
R651 B.n678 B.n19 163.367
R652 B.n679 B.n678 163.367
R653 B.n680 B.n679 163.367
R654 B.n680 B.n17 163.367
R655 B.n684 B.n17 163.367
R656 B.n685 B.n684 163.367
R657 B.n686 B.n685 163.367
R658 B.n686 B.n15 163.367
R659 B.n690 B.n15 163.367
R660 B.n691 B.n690 163.367
R661 B.n692 B.n691 163.367
R662 B.n692 B.n13 163.367
R663 B.n696 B.n13 163.367
R664 B.n697 B.n696 163.367
R665 B.n698 B.n697 163.367
R666 B.n698 B.n11 163.367
R667 B.n702 B.n11 163.367
R668 B.n703 B.n702 163.367
R669 B.n704 B.n703 163.367
R670 B.n704 B.n9 163.367
R671 B.n708 B.n9 163.367
R672 B.n709 B.n708 163.367
R673 B.n710 B.n709 163.367
R674 B.n710 B.n7 163.367
R675 B.n714 B.n7 163.367
R676 B.n715 B.n714 163.367
R677 B.n716 B.n715 163.367
R678 B.n716 B.n5 163.367
R679 B.n720 B.n5 163.367
R680 B.n721 B.n720 163.367
R681 B.n722 B.n721 163.367
R682 B.n722 B.n3 163.367
R683 B.n726 B.n3 163.367
R684 B.n727 B.n726 163.367
R685 B.n188 B.n2 163.367
R686 B.n189 B.n188 163.367
R687 B.n190 B.n189 163.367
R688 B.n190 B.n185 163.367
R689 B.n194 B.n185 163.367
R690 B.n195 B.n194 163.367
R691 B.n196 B.n195 163.367
R692 B.n196 B.n183 163.367
R693 B.n200 B.n183 163.367
R694 B.n201 B.n200 163.367
R695 B.n202 B.n201 163.367
R696 B.n202 B.n181 163.367
R697 B.n206 B.n181 163.367
R698 B.n207 B.n206 163.367
R699 B.n208 B.n207 163.367
R700 B.n208 B.n179 163.367
R701 B.n212 B.n179 163.367
R702 B.n213 B.n212 163.367
R703 B.n214 B.n213 163.367
R704 B.n214 B.n177 163.367
R705 B.n218 B.n177 163.367
R706 B.n219 B.n218 163.367
R707 B.n220 B.n219 163.367
R708 B.n220 B.n175 163.367
R709 B.n224 B.n175 163.367
R710 B.n225 B.n224 163.367
R711 B.n226 B.n225 163.367
R712 B.n226 B.n173 163.367
R713 B.n230 B.n173 163.367
R714 B.n231 B.n230 163.367
R715 B.n232 B.n231 163.367
R716 B.n232 B.n171 163.367
R717 B.n236 B.n171 163.367
R718 B.n237 B.n236 163.367
R719 B.n238 B.n237 163.367
R720 B.n238 B.n169 163.367
R721 B.n242 B.n169 163.367
R722 B.n243 B.n242 163.367
R723 B.n244 B.n243 163.367
R724 B.n244 B.n167 163.367
R725 B.n248 B.n167 163.367
R726 B.n249 B.n248 163.367
R727 B.n250 B.n249 163.367
R728 B.n250 B.n165 163.367
R729 B.n254 B.n165 163.367
R730 B.n312 B.n145 59.5399
R731 B.n328 B.n327 59.5399
R732 B.n586 B.n53 59.5399
R733 B.n46 B.n45 59.5399
R734 B.n145 B.n144 42.4732
R735 B.n327 B.n326 42.4732
R736 B.n53 B.n52 42.4732
R737 B.n45 B.n44 42.4732
R738 B.n659 B.n658 34.4981
R739 B.n527 B.n72 34.4981
R740 B.n388 B.n387 34.4981
R741 B.n253 B.n164 34.4981
R742 B B.n729 18.0485
R743 B.n659 B.n24 10.6151
R744 B.n663 B.n24 10.6151
R745 B.n664 B.n663 10.6151
R746 B.n665 B.n664 10.6151
R747 B.n665 B.n22 10.6151
R748 B.n669 B.n22 10.6151
R749 B.n670 B.n669 10.6151
R750 B.n671 B.n670 10.6151
R751 B.n671 B.n20 10.6151
R752 B.n675 B.n20 10.6151
R753 B.n676 B.n675 10.6151
R754 B.n677 B.n676 10.6151
R755 B.n677 B.n18 10.6151
R756 B.n681 B.n18 10.6151
R757 B.n682 B.n681 10.6151
R758 B.n683 B.n682 10.6151
R759 B.n683 B.n16 10.6151
R760 B.n687 B.n16 10.6151
R761 B.n688 B.n687 10.6151
R762 B.n689 B.n688 10.6151
R763 B.n689 B.n14 10.6151
R764 B.n693 B.n14 10.6151
R765 B.n694 B.n693 10.6151
R766 B.n695 B.n694 10.6151
R767 B.n695 B.n12 10.6151
R768 B.n699 B.n12 10.6151
R769 B.n700 B.n699 10.6151
R770 B.n701 B.n700 10.6151
R771 B.n701 B.n10 10.6151
R772 B.n705 B.n10 10.6151
R773 B.n706 B.n705 10.6151
R774 B.n707 B.n706 10.6151
R775 B.n707 B.n8 10.6151
R776 B.n711 B.n8 10.6151
R777 B.n712 B.n711 10.6151
R778 B.n713 B.n712 10.6151
R779 B.n713 B.n6 10.6151
R780 B.n717 B.n6 10.6151
R781 B.n718 B.n717 10.6151
R782 B.n719 B.n718 10.6151
R783 B.n719 B.n4 10.6151
R784 B.n723 B.n4 10.6151
R785 B.n724 B.n723 10.6151
R786 B.n725 B.n724 10.6151
R787 B.n725 B.n0 10.6151
R788 B.n658 B.n657 10.6151
R789 B.n657 B.n26 10.6151
R790 B.n653 B.n26 10.6151
R791 B.n653 B.n652 10.6151
R792 B.n652 B.n651 10.6151
R793 B.n651 B.n28 10.6151
R794 B.n647 B.n28 10.6151
R795 B.n647 B.n646 10.6151
R796 B.n646 B.n645 10.6151
R797 B.n645 B.n30 10.6151
R798 B.n641 B.n30 10.6151
R799 B.n641 B.n640 10.6151
R800 B.n640 B.n639 10.6151
R801 B.n639 B.n32 10.6151
R802 B.n635 B.n32 10.6151
R803 B.n635 B.n634 10.6151
R804 B.n634 B.n633 10.6151
R805 B.n633 B.n34 10.6151
R806 B.n629 B.n34 10.6151
R807 B.n629 B.n628 10.6151
R808 B.n628 B.n627 10.6151
R809 B.n627 B.n36 10.6151
R810 B.n623 B.n36 10.6151
R811 B.n623 B.n622 10.6151
R812 B.n622 B.n621 10.6151
R813 B.n621 B.n38 10.6151
R814 B.n617 B.n38 10.6151
R815 B.n617 B.n616 10.6151
R816 B.n616 B.n615 10.6151
R817 B.n615 B.n40 10.6151
R818 B.n611 B.n40 10.6151
R819 B.n611 B.n610 10.6151
R820 B.n610 B.n609 10.6151
R821 B.n609 B.n42 10.6151
R822 B.n605 B.n42 10.6151
R823 B.n605 B.n604 10.6151
R824 B.n604 B.n603 10.6151
R825 B.n600 B.n599 10.6151
R826 B.n599 B.n598 10.6151
R827 B.n598 B.n48 10.6151
R828 B.n594 B.n48 10.6151
R829 B.n594 B.n593 10.6151
R830 B.n593 B.n592 10.6151
R831 B.n592 B.n50 10.6151
R832 B.n588 B.n50 10.6151
R833 B.n588 B.n587 10.6151
R834 B.n585 B.n54 10.6151
R835 B.n581 B.n54 10.6151
R836 B.n581 B.n580 10.6151
R837 B.n580 B.n579 10.6151
R838 B.n579 B.n56 10.6151
R839 B.n575 B.n56 10.6151
R840 B.n575 B.n574 10.6151
R841 B.n574 B.n573 10.6151
R842 B.n573 B.n58 10.6151
R843 B.n569 B.n58 10.6151
R844 B.n569 B.n568 10.6151
R845 B.n568 B.n567 10.6151
R846 B.n567 B.n60 10.6151
R847 B.n563 B.n60 10.6151
R848 B.n563 B.n562 10.6151
R849 B.n562 B.n561 10.6151
R850 B.n561 B.n62 10.6151
R851 B.n557 B.n62 10.6151
R852 B.n557 B.n556 10.6151
R853 B.n556 B.n555 10.6151
R854 B.n555 B.n64 10.6151
R855 B.n551 B.n64 10.6151
R856 B.n551 B.n550 10.6151
R857 B.n550 B.n549 10.6151
R858 B.n549 B.n66 10.6151
R859 B.n545 B.n66 10.6151
R860 B.n545 B.n544 10.6151
R861 B.n544 B.n543 10.6151
R862 B.n543 B.n68 10.6151
R863 B.n539 B.n68 10.6151
R864 B.n539 B.n538 10.6151
R865 B.n538 B.n537 10.6151
R866 B.n537 B.n70 10.6151
R867 B.n533 B.n70 10.6151
R868 B.n533 B.n532 10.6151
R869 B.n532 B.n531 10.6151
R870 B.n531 B.n72 10.6151
R871 B.n527 B.n526 10.6151
R872 B.n526 B.n525 10.6151
R873 B.n525 B.n74 10.6151
R874 B.n521 B.n74 10.6151
R875 B.n521 B.n520 10.6151
R876 B.n520 B.n519 10.6151
R877 B.n519 B.n76 10.6151
R878 B.n515 B.n76 10.6151
R879 B.n515 B.n514 10.6151
R880 B.n514 B.n513 10.6151
R881 B.n513 B.n78 10.6151
R882 B.n509 B.n78 10.6151
R883 B.n509 B.n508 10.6151
R884 B.n508 B.n507 10.6151
R885 B.n507 B.n80 10.6151
R886 B.n503 B.n80 10.6151
R887 B.n503 B.n502 10.6151
R888 B.n502 B.n501 10.6151
R889 B.n501 B.n82 10.6151
R890 B.n497 B.n82 10.6151
R891 B.n497 B.n496 10.6151
R892 B.n496 B.n495 10.6151
R893 B.n495 B.n84 10.6151
R894 B.n491 B.n84 10.6151
R895 B.n491 B.n490 10.6151
R896 B.n490 B.n489 10.6151
R897 B.n489 B.n86 10.6151
R898 B.n485 B.n86 10.6151
R899 B.n485 B.n484 10.6151
R900 B.n484 B.n483 10.6151
R901 B.n483 B.n88 10.6151
R902 B.n479 B.n88 10.6151
R903 B.n479 B.n478 10.6151
R904 B.n478 B.n477 10.6151
R905 B.n477 B.n90 10.6151
R906 B.n473 B.n90 10.6151
R907 B.n473 B.n472 10.6151
R908 B.n472 B.n471 10.6151
R909 B.n471 B.n92 10.6151
R910 B.n467 B.n92 10.6151
R911 B.n467 B.n466 10.6151
R912 B.n466 B.n465 10.6151
R913 B.n465 B.n94 10.6151
R914 B.n461 B.n94 10.6151
R915 B.n461 B.n460 10.6151
R916 B.n460 B.n459 10.6151
R917 B.n459 B.n96 10.6151
R918 B.n455 B.n96 10.6151
R919 B.n455 B.n454 10.6151
R920 B.n454 B.n453 10.6151
R921 B.n453 B.n98 10.6151
R922 B.n449 B.n98 10.6151
R923 B.n449 B.n448 10.6151
R924 B.n448 B.n447 10.6151
R925 B.n447 B.n100 10.6151
R926 B.n443 B.n100 10.6151
R927 B.n443 B.n442 10.6151
R928 B.n442 B.n441 10.6151
R929 B.n441 B.n102 10.6151
R930 B.n437 B.n102 10.6151
R931 B.n437 B.n436 10.6151
R932 B.n436 B.n435 10.6151
R933 B.n435 B.n104 10.6151
R934 B.n431 B.n104 10.6151
R935 B.n431 B.n430 10.6151
R936 B.n430 B.n429 10.6151
R937 B.n429 B.n106 10.6151
R938 B.n425 B.n106 10.6151
R939 B.n425 B.n424 10.6151
R940 B.n424 B.n423 10.6151
R941 B.n423 B.n108 10.6151
R942 B.n419 B.n108 10.6151
R943 B.n419 B.n418 10.6151
R944 B.n418 B.n417 10.6151
R945 B.n417 B.n110 10.6151
R946 B.n413 B.n110 10.6151
R947 B.n413 B.n412 10.6151
R948 B.n412 B.n411 10.6151
R949 B.n411 B.n112 10.6151
R950 B.n407 B.n112 10.6151
R951 B.n407 B.n406 10.6151
R952 B.n406 B.n405 10.6151
R953 B.n405 B.n114 10.6151
R954 B.n401 B.n114 10.6151
R955 B.n401 B.n400 10.6151
R956 B.n400 B.n399 10.6151
R957 B.n399 B.n116 10.6151
R958 B.n395 B.n116 10.6151
R959 B.n395 B.n394 10.6151
R960 B.n394 B.n393 10.6151
R961 B.n393 B.n118 10.6151
R962 B.n389 B.n118 10.6151
R963 B.n389 B.n388 10.6151
R964 B.n187 B.n1 10.6151
R965 B.n187 B.n186 10.6151
R966 B.n191 B.n186 10.6151
R967 B.n192 B.n191 10.6151
R968 B.n193 B.n192 10.6151
R969 B.n193 B.n184 10.6151
R970 B.n197 B.n184 10.6151
R971 B.n198 B.n197 10.6151
R972 B.n199 B.n198 10.6151
R973 B.n199 B.n182 10.6151
R974 B.n203 B.n182 10.6151
R975 B.n204 B.n203 10.6151
R976 B.n205 B.n204 10.6151
R977 B.n205 B.n180 10.6151
R978 B.n209 B.n180 10.6151
R979 B.n210 B.n209 10.6151
R980 B.n211 B.n210 10.6151
R981 B.n211 B.n178 10.6151
R982 B.n215 B.n178 10.6151
R983 B.n216 B.n215 10.6151
R984 B.n217 B.n216 10.6151
R985 B.n217 B.n176 10.6151
R986 B.n221 B.n176 10.6151
R987 B.n222 B.n221 10.6151
R988 B.n223 B.n222 10.6151
R989 B.n223 B.n174 10.6151
R990 B.n227 B.n174 10.6151
R991 B.n228 B.n227 10.6151
R992 B.n229 B.n228 10.6151
R993 B.n229 B.n172 10.6151
R994 B.n233 B.n172 10.6151
R995 B.n234 B.n233 10.6151
R996 B.n235 B.n234 10.6151
R997 B.n235 B.n170 10.6151
R998 B.n239 B.n170 10.6151
R999 B.n240 B.n239 10.6151
R1000 B.n241 B.n240 10.6151
R1001 B.n241 B.n168 10.6151
R1002 B.n245 B.n168 10.6151
R1003 B.n246 B.n245 10.6151
R1004 B.n247 B.n246 10.6151
R1005 B.n247 B.n166 10.6151
R1006 B.n251 B.n166 10.6151
R1007 B.n252 B.n251 10.6151
R1008 B.n253 B.n252 10.6151
R1009 B.n257 B.n164 10.6151
R1010 B.n258 B.n257 10.6151
R1011 B.n259 B.n258 10.6151
R1012 B.n259 B.n162 10.6151
R1013 B.n263 B.n162 10.6151
R1014 B.n264 B.n263 10.6151
R1015 B.n265 B.n264 10.6151
R1016 B.n265 B.n160 10.6151
R1017 B.n269 B.n160 10.6151
R1018 B.n270 B.n269 10.6151
R1019 B.n271 B.n270 10.6151
R1020 B.n271 B.n158 10.6151
R1021 B.n275 B.n158 10.6151
R1022 B.n276 B.n275 10.6151
R1023 B.n277 B.n276 10.6151
R1024 B.n277 B.n156 10.6151
R1025 B.n281 B.n156 10.6151
R1026 B.n282 B.n281 10.6151
R1027 B.n283 B.n282 10.6151
R1028 B.n283 B.n154 10.6151
R1029 B.n287 B.n154 10.6151
R1030 B.n288 B.n287 10.6151
R1031 B.n289 B.n288 10.6151
R1032 B.n289 B.n152 10.6151
R1033 B.n293 B.n152 10.6151
R1034 B.n294 B.n293 10.6151
R1035 B.n295 B.n294 10.6151
R1036 B.n295 B.n150 10.6151
R1037 B.n299 B.n150 10.6151
R1038 B.n300 B.n299 10.6151
R1039 B.n301 B.n300 10.6151
R1040 B.n301 B.n148 10.6151
R1041 B.n305 B.n148 10.6151
R1042 B.n306 B.n305 10.6151
R1043 B.n307 B.n306 10.6151
R1044 B.n307 B.n146 10.6151
R1045 B.n311 B.n146 10.6151
R1046 B.n314 B.n313 10.6151
R1047 B.n314 B.n142 10.6151
R1048 B.n318 B.n142 10.6151
R1049 B.n319 B.n318 10.6151
R1050 B.n320 B.n319 10.6151
R1051 B.n320 B.n140 10.6151
R1052 B.n324 B.n140 10.6151
R1053 B.n325 B.n324 10.6151
R1054 B.n329 B.n325 10.6151
R1055 B.n333 B.n138 10.6151
R1056 B.n334 B.n333 10.6151
R1057 B.n335 B.n334 10.6151
R1058 B.n335 B.n136 10.6151
R1059 B.n339 B.n136 10.6151
R1060 B.n340 B.n339 10.6151
R1061 B.n341 B.n340 10.6151
R1062 B.n341 B.n134 10.6151
R1063 B.n345 B.n134 10.6151
R1064 B.n346 B.n345 10.6151
R1065 B.n347 B.n346 10.6151
R1066 B.n347 B.n132 10.6151
R1067 B.n351 B.n132 10.6151
R1068 B.n352 B.n351 10.6151
R1069 B.n353 B.n352 10.6151
R1070 B.n353 B.n130 10.6151
R1071 B.n357 B.n130 10.6151
R1072 B.n358 B.n357 10.6151
R1073 B.n359 B.n358 10.6151
R1074 B.n359 B.n128 10.6151
R1075 B.n363 B.n128 10.6151
R1076 B.n364 B.n363 10.6151
R1077 B.n365 B.n364 10.6151
R1078 B.n365 B.n126 10.6151
R1079 B.n369 B.n126 10.6151
R1080 B.n370 B.n369 10.6151
R1081 B.n371 B.n370 10.6151
R1082 B.n371 B.n124 10.6151
R1083 B.n375 B.n124 10.6151
R1084 B.n376 B.n375 10.6151
R1085 B.n377 B.n376 10.6151
R1086 B.n377 B.n122 10.6151
R1087 B.n381 B.n122 10.6151
R1088 B.n382 B.n381 10.6151
R1089 B.n383 B.n382 10.6151
R1090 B.n383 B.n120 10.6151
R1091 B.n387 B.n120 10.6151
R1092 B.n603 B.n46 9.36635
R1093 B.n586 B.n585 9.36635
R1094 B.n312 B.n311 9.36635
R1095 B.n328 B.n138 9.36635
R1096 B.n729 B.n0 8.11757
R1097 B.n729 B.n1 8.11757
R1098 B.n600 B.n46 1.24928
R1099 B.n587 B.n586 1.24928
R1100 B.n313 B.n312 1.24928
R1101 B.n329 B.n328 1.24928
R1102 VP.n16 VP.t3 170.185
R1103 VP.n18 VP.n15 161.3
R1104 VP.n20 VP.n19 161.3
R1105 VP.n21 VP.n14 161.3
R1106 VP.n23 VP.n22 161.3
R1107 VP.n24 VP.n13 161.3
R1108 VP.n26 VP.n25 161.3
R1109 VP.n27 VP.n12 161.3
R1110 VP.n29 VP.n28 161.3
R1111 VP.n30 VP.n11 161.3
R1112 VP.n33 VP.n32 161.3
R1113 VP.n34 VP.n10 161.3
R1114 VP.n36 VP.n35 161.3
R1115 VP.n37 VP.n9 161.3
R1116 VP.n68 VP.n0 161.3
R1117 VP.n67 VP.n66 161.3
R1118 VP.n65 VP.n1 161.3
R1119 VP.n64 VP.n63 161.3
R1120 VP.n61 VP.n2 161.3
R1121 VP.n60 VP.n59 161.3
R1122 VP.n58 VP.n3 161.3
R1123 VP.n57 VP.n56 161.3
R1124 VP.n55 VP.n4 161.3
R1125 VP.n54 VP.n53 161.3
R1126 VP.n52 VP.n5 161.3
R1127 VP.n51 VP.n50 161.3
R1128 VP.n49 VP.n6 161.3
R1129 VP.n47 VP.n46 161.3
R1130 VP.n45 VP.n7 161.3
R1131 VP.n44 VP.n43 161.3
R1132 VP.n42 VP.n8 161.3
R1133 VP.n55 VP.t1 140.196
R1134 VP.n41 VP.t6 140.196
R1135 VP.n48 VP.t4 140.196
R1136 VP.n62 VP.t5 140.196
R1137 VP.n69 VP.t2 140.196
R1138 VP.n24 VP.t0 140.196
R1139 VP.n38 VP.t9 140.196
R1140 VP.n31 VP.t8 140.196
R1141 VP.n17 VP.t7 140.196
R1142 VP.n41 VP.n40 92.1052
R1143 VP.n70 VP.n69 92.1052
R1144 VP.n39 VP.n38 92.1052
R1145 VP.n17 VP.n16 60.1448
R1146 VP.n43 VP.n7 56.4773
R1147 VP.n67 VP.n1 56.4773
R1148 VP.n36 VP.n10 56.4773
R1149 VP.n50 VP.n5 49.6611
R1150 VP.n60 VP.n3 49.6611
R1151 VP.n29 VP.n12 49.6611
R1152 VP.n19 VP.n14 49.6611
R1153 VP.n40 VP.n39 48.17
R1154 VP.n54 VP.n5 31.1601
R1155 VP.n56 VP.n3 31.1601
R1156 VP.n25 VP.n12 31.1601
R1157 VP.n23 VP.n14 31.1601
R1158 VP.n43 VP.n42 24.3439
R1159 VP.n47 VP.n7 24.3439
R1160 VP.n50 VP.n49 24.3439
R1161 VP.n55 VP.n54 24.3439
R1162 VP.n56 VP.n55 24.3439
R1163 VP.n61 VP.n60 24.3439
R1164 VP.n63 VP.n1 24.3439
R1165 VP.n68 VP.n67 24.3439
R1166 VP.n37 VP.n36 24.3439
R1167 VP.n30 VP.n29 24.3439
R1168 VP.n32 VP.n10 24.3439
R1169 VP.n24 VP.n23 24.3439
R1170 VP.n25 VP.n24 24.3439
R1171 VP.n19 VP.n18 24.3439
R1172 VP.n42 VP.n41 18.5015
R1173 VP.n69 VP.n68 18.5015
R1174 VP.n38 VP.n37 18.5015
R1175 VP.n48 VP.n47 15.0934
R1176 VP.n63 VP.n62 15.0934
R1177 VP.n32 VP.n31 15.0934
R1178 VP.n16 VP.n15 13.5258
R1179 VP.n49 VP.n48 9.251
R1180 VP.n62 VP.n61 9.251
R1181 VP.n31 VP.n30 9.251
R1182 VP.n18 VP.n17 9.251
R1183 VP.n39 VP.n9 0.278398
R1184 VP.n40 VP.n8 0.278398
R1185 VP.n70 VP.n0 0.278398
R1186 VP.n20 VP.n15 0.189894
R1187 VP.n21 VP.n20 0.189894
R1188 VP.n22 VP.n21 0.189894
R1189 VP.n22 VP.n13 0.189894
R1190 VP.n26 VP.n13 0.189894
R1191 VP.n27 VP.n26 0.189894
R1192 VP.n28 VP.n27 0.189894
R1193 VP.n28 VP.n11 0.189894
R1194 VP.n33 VP.n11 0.189894
R1195 VP.n34 VP.n33 0.189894
R1196 VP.n35 VP.n34 0.189894
R1197 VP.n35 VP.n9 0.189894
R1198 VP.n44 VP.n8 0.189894
R1199 VP.n45 VP.n44 0.189894
R1200 VP.n46 VP.n45 0.189894
R1201 VP.n46 VP.n6 0.189894
R1202 VP.n51 VP.n6 0.189894
R1203 VP.n52 VP.n51 0.189894
R1204 VP.n53 VP.n52 0.189894
R1205 VP.n53 VP.n4 0.189894
R1206 VP.n57 VP.n4 0.189894
R1207 VP.n58 VP.n57 0.189894
R1208 VP.n59 VP.n58 0.189894
R1209 VP.n59 VP.n2 0.189894
R1210 VP.n64 VP.n2 0.189894
R1211 VP.n65 VP.n64 0.189894
R1212 VP.n66 VP.n65 0.189894
R1213 VP.n66 VP.n0 0.189894
R1214 VP VP.n70 0.153422
R1215 VTAIL.n240 VTAIL.n188 756.745
R1216 VTAIL.n54 VTAIL.n2 756.745
R1217 VTAIL.n182 VTAIL.n130 756.745
R1218 VTAIL.n120 VTAIL.n68 756.745
R1219 VTAIL.n207 VTAIL.n206 585
R1220 VTAIL.n204 VTAIL.n203 585
R1221 VTAIL.n213 VTAIL.n212 585
R1222 VTAIL.n215 VTAIL.n214 585
R1223 VTAIL.n200 VTAIL.n199 585
R1224 VTAIL.n221 VTAIL.n220 585
R1225 VTAIL.n224 VTAIL.n223 585
R1226 VTAIL.n222 VTAIL.n196 585
R1227 VTAIL.n229 VTAIL.n195 585
R1228 VTAIL.n231 VTAIL.n230 585
R1229 VTAIL.n233 VTAIL.n232 585
R1230 VTAIL.n192 VTAIL.n191 585
R1231 VTAIL.n239 VTAIL.n238 585
R1232 VTAIL.n241 VTAIL.n240 585
R1233 VTAIL.n21 VTAIL.n20 585
R1234 VTAIL.n18 VTAIL.n17 585
R1235 VTAIL.n27 VTAIL.n26 585
R1236 VTAIL.n29 VTAIL.n28 585
R1237 VTAIL.n14 VTAIL.n13 585
R1238 VTAIL.n35 VTAIL.n34 585
R1239 VTAIL.n38 VTAIL.n37 585
R1240 VTAIL.n36 VTAIL.n10 585
R1241 VTAIL.n43 VTAIL.n9 585
R1242 VTAIL.n45 VTAIL.n44 585
R1243 VTAIL.n47 VTAIL.n46 585
R1244 VTAIL.n6 VTAIL.n5 585
R1245 VTAIL.n53 VTAIL.n52 585
R1246 VTAIL.n55 VTAIL.n54 585
R1247 VTAIL.n183 VTAIL.n182 585
R1248 VTAIL.n181 VTAIL.n180 585
R1249 VTAIL.n134 VTAIL.n133 585
R1250 VTAIL.n175 VTAIL.n174 585
R1251 VTAIL.n173 VTAIL.n172 585
R1252 VTAIL.n171 VTAIL.n137 585
R1253 VTAIL.n141 VTAIL.n138 585
R1254 VTAIL.n166 VTAIL.n165 585
R1255 VTAIL.n164 VTAIL.n163 585
R1256 VTAIL.n143 VTAIL.n142 585
R1257 VTAIL.n158 VTAIL.n157 585
R1258 VTAIL.n156 VTAIL.n155 585
R1259 VTAIL.n147 VTAIL.n146 585
R1260 VTAIL.n150 VTAIL.n149 585
R1261 VTAIL.n121 VTAIL.n120 585
R1262 VTAIL.n119 VTAIL.n118 585
R1263 VTAIL.n72 VTAIL.n71 585
R1264 VTAIL.n113 VTAIL.n112 585
R1265 VTAIL.n111 VTAIL.n110 585
R1266 VTAIL.n109 VTAIL.n75 585
R1267 VTAIL.n79 VTAIL.n76 585
R1268 VTAIL.n104 VTAIL.n103 585
R1269 VTAIL.n102 VTAIL.n101 585
R1270 VTAIL.n81 VTAIL.n80 585
R1271 VTAIL.n96 VTAIL.n95 585
R1272 VTAIL.n94 VTAIL.n93 585
R1273 VTAIL.n85 VTAIL.n84 585
R1274 VTAIL.n88 VTAIL.n87 585
R1275 VTAIL.t18 VTAIL.n148 329.038
R1276 VTAIL.t7 VTAIL.n86 329.038
R1277 VTAIL.t5 VTAIL.n205 329.038
R1278 VTAIL.t15 VTAIL.n19 329.038
R1279 VTAIL.n206 VTAIL.n203 171.744
R1280 VTAIL.n213 VTAIL.n203 171.744
R1281 VTAIL.n214 VTAIL.n213 171.744
R1282 VTAIL.n214 VTAIL.n199 171.744
R1283 VTAIL.n221 VTAIL.n199 171.744
R1284 VTAIL.n223 VTAIL.n221 171.744
R1285 VTAIL.n223 VTAIL.n222 171.744
R1286 VTAIL.n222 VTAIL.n195 171.744
R1287 VTAIL.n231 VTAIL.n195 171.744
R1288 VTAIL.n232 VTAIL.n231 171.744
R1289 VTAIL.n232 VTAIL.n191 171.744
R1290 VTAIL.n239 VTAIL.n191 171.744
R1291 VTAIL.n240 VTAIL.n239 171.744
R1292 VTAIL.n20 VTAIL.n17 171.744
R1293 VTAIL.n27 VTAIL.n17 171.744
R1294 VTAIL.n28 VTAIL.n27 171.744
R1295 VTAIL.n28 VTAIL.n13 171.744
R1296 VTAIL.n35 VTAIL.n13 171.744
R1297 VTAIL.n37 VTAIL.n35 171.744
R1298 VTAIL.n37 VTAIL.n36 171.744
R1299 VTAIL.n36 VTAIL.n9 171.744
R1300 VTAIL.n45 VTAIL.n9 171.744
R1301 VTAIL.n46 VTAIL.n45 171.744
R1302 VTAIL.n46 VTAIL.n5 171.744
R1303 VTAIL.n53 VTAIL.n5 171.744
R1304 VTAIL.n54 VTAIL.n53 171.744
R1305 VTAIL.n182 VTAIL.n181 171.744
R1306 VTAIL.n181 VTAIL.n133 171.744
R1307 VTAIL.n174 VTAIL.n133 171.744
R1308 VTAIL.n174 VTAIL.n173 171.744
R1309 VTAIL.n173 VTAIL.n137 171.744
R1310 VTAIL.n141 VTAIL.n137 171.744
R1311 VTAIL.n165 VTAIL.n141 171.744
R1312 VTAIL.n165 VTAIL.n164 171.744
R1313 VTAIL.n164 VTAIL.n142 171.744
R1314 VTAIL.n157 VTAIL.n142 171.744
R1315 VTAIL.n157 VTAIL.n156 171.744
R1316 VTAIL.n156 VTAIL.n146 171.744
R1317 VTAIL.n149 VTAIL.n146 171.744
R1318 VTAIL.n120 VTAIL.n119 171.744
R1319 VTAIL.n119 VTAIL.n71 171.744
R1320 VTAIL.n112 VTAIL.n71 171.744
R1321 VTAIL.n112 VTAIL.n111 171.744
R1322 VTAIL.n111 VTAIL.n75 171.744
R1323 VTAIL.n79 VTAIL.n75 171.744
R1324 VTAIL.n103 VTAIL.n79 171.744
R1325 VTAIL.n103 VTAIL.n102 171.744
R1326 VTAIL.n102 VTAIL.n80 171.744
R1327 VTAIL.n95 VTAIL.n80 171.744
R1328 VTAIL.n95 VTAIL.n94 171.744
R1329 VTAIL.n94 VTAIL.n84 171.744
R1330 VTAIL.n87 VTAIL.n84 171.744
R1331 VTAIL.n206 VTAIL.t5 85.8723
R1332 VTAIL.n20 VTAIL.t15 85.8723
R1333 VTAIL.n149 VTAIL.t18 85.8723
R1334 VTAIL.n87 VTAIL.t7 85.8723
R1335 VTAIL.n129 VTAIL.n128 61.9025
R1336 VTAIL.n127 VTAIL.n126 61.9025
R1337 VTAIL.n67 VTAIL.n66 61.9025
R1338 VTAIL.n65 VTAIL.n64 61.9025
R1339 VTAIL.n247 VTAIL.n246 61.9023
R1340 VTAIL.n1 VTAIL.n0 61.9023
R1341 VTAIL.n61 VTAIL.n60 61.9023
R1342 VTAIL.n63 VTAIL.n62 61.9023
R1343 VTAIL.n245 VTAIL.n244 34.9005
R1344 VTAIL.n59 VTAIL.n58 34.9005
R1345 VTAIL.n187 VTAIL.n186 34.9005
R1346 VTAIL.n125 VTAIL.n124 34.9005
R1347 VTAIL.n65 VTAIL.n63 25.4703
R1348 VTAIL.n245 VTAIL.n187 23.5824
R1349 VTAIL.n230 VTAIL.n229 13.1884
R1350 VTAIL.n44 VTAIL.n43 13.1884
R1351 VTAIL.n172 VTAIL.n171 13.1884
R1352 VTAIL.n110 VTAIL.n109 13.1884
R1353 VTAIL.n228 VTAIL.n196 12.8005
R1354 VTAIL.n233 VTAIL.n194 12.8005
R1355 VTAIL.n42 VTAIL.n10 12.8005
R1356 VTAIL.n47 VTAIL.n8 12.8005
R1357 VTAIL.n175 VTAIL.n136 12.8005
R1358 VTAIL.n170 VTAIL.n138 12.8005
R1359 VTAIL.n113 VTAIL.n74 12.8005
R1360 VTAIL.n108 VTAIL.n76 12.8005
R1361 VTAIL.n225 VTAIL.n224 12.0247
R1362 VTAIL.n234 VTAIL.n192 12.0247
R1363 VTAIL.n39 VTAIL.n38 12.0247
R1364 VTAIL.n48 VTAIL.n6 12.0247
R1365 VTAIL.n176 VTAIL.n134 12.0247
R1366 VTAIL.n167 VTAIL.n166 12.0247
R1367 VTAIL.n114 VTAIL.n72 12.0247
R1368 VTAIL.n105 VTAIL.n104 12.0247
R1369 VTAIL.n220 VTAIL.n198 11.249
R1370 VTAIL.n238 VTAIL.n237 11.249
R1371 VTAIL.n34 VTAIL.n12 11.249
R1372 VTAIL.n52 VTAIL.n51 11.249
R1373 VTAIL.n180 VTAIL.n179 11.249
R1374 VTAIL.n163 VTAIL.n140 11.249
R1375 VTAIL.n118 VTAIL.n117 11.249
R1376 VTAIL.n101 VTAIL.n78 11.249
R1377 VTAIL.n207 VTAIL.n205 10.7239
R1378 VTAIL.n21 VTAIL.n19 10.7239
R1379 VTAIL.n150 VTAIL.n148 10.7239
R1380 VTAIL.n88 VTAIL.n86 10.7239
R1381 VTAIL.n219 VTAIL.n200 10.4732
R1382 VTAIL.n241 VTAIL.n190 10.4732
R1383 VTAIL.n33 VTAIL.n14 10.4732
R1384 VTAIL.n55 VTAIL.n4 10.4732
R1385 VTAIL.n183 VTAIL.n132 10.4732
R1386 VTAIL.n162 VTAIL.n143 10.4732
R1387 VTAIL.n121 VTAIL.n70 10.4732
R1388 VTAIL.n100 VTAIL.n81 10.4732
R1389 VTAIL.n216 VTAIL.n215 9.69747
R1390 VTAIL.n242 VTAIL.n188 9.69747
R1391 VTAIL.n30 VTAIL.n29 9.69747
R1392 VTAIL.n56 VTAIL.n2 9.69747
R1393 VTAIL.n184 VTAIL.n130 9.69747
R1394 VTAIL.n159 VTAIL.n158 9.69747
R1395 VTAIL.n122 VTAIL.n68 9.69747
R1396 VTAIL.n97 VTAIL.n96 9.69747
R1397 VTAIL.n244 VTAIL.n243 9.45567
R1398 VTAIL.n58 VTAIL.n57 9.45567
R1399 VTAIL.n186 VTAIL.n185 9.45567
R1400 VTAIL.n124 VTAIL.n123 9.45567
R1401 VTAIL.n243 VTAIL.n242 9.3005
R1402 VTAIL.n190 VTAIL.n189 9.3005
R1403 VTAIL.n237 VTAIL.n236 9.3005
R1404 VTAIL.n235 VTAIL.n234 9.3005
R1405 VTAIL.n194 VTAIL.n193 9.3005
R1406 VTAIL.n209 VTAIL.n208 9.3005
R1407 VTAIL.n211 VTAIL.n210 9.3005
R1408 VTAIL.n202 VTAIL.n201 9.3005
R1409 VTAIL.n217 VTAIL.n216 9.3005
R1410 VTAIL.n219 VTAIL.n218 9.3005
R1411 VTAIL.n198 VTAIL.n197 9.3005
R1412 VTAIL.n226 VTAIL.n225 9.3005
R1413 VTAIL.n228 VTAIL.n227 9.3005
R1414 VTAIL.n57 VTAIL.n56 9.3005
R1415 VTAIL.n4 VTAIL.n3 9.3005
R1416 VTAIL.n51 VTAIL.n50 9.3005
R1417 VTAIL.n49 VTAIL.n48 9.3005
R1418 VTAIL.n8 VTAIL.n7 9.3005
R1419 VTAIL.n23 VTAIL.n22 9.3005
R1420 VTAIL.n25 VTAIL.n24 9.3005
R1421 VTAIL.n16 VTAIL.n15 9.3005
R1422 VTAIL.n31 VTAIL.n30 9.3005
R1423 VTAIL.n33 VTAIL.n32 9.3005
R1424 VTAIL.n12 VTAIL.n11 9.3005
R1425 VTAIL.n40 VTAIL.n39 9.3005
R1426 VTAIL.n42 VTAIL.n41 9.3005
R1427 VTAIL.n152 VTAIL.n151 9.3005
R1428 VTAIL.n154 VTAIL.n153 9.3005
R1429 VTAIL.n145 VTAIL.n144 9.3005
R1430 VTAIL.n160 VTAIL.n159 9.3005
R1431 VTAIL.n162 VTAIL.n161 9.3005
R1432 VTAIL.n140 VTAIL.n139 9.3005
R1433 VTAIL.n168 VTAIL.n167 9.3005
R1434 VTAIL.n170 VTAIL.n169 9.3005
R1435 VTAIL.n185 VTAIL.n184 9.3005
R1436 VTAIL.n132 VTAIL.n131 9.3005
R1437 VTAIL.n179 VTAIL.n178 9.3005
R1438 VTAIL.n177 VTAIL.n176 9.3005
R1439 VTAIL.n136 VTAIL.n135 9.3005
R1440 VTAIL.n90 VTAIL.n89 9.3005
R1441 VTAIL.n92 VTAIL.n91 9.3005
R1442 VTAIL.n83 VTAIL.n82 9.3005
R1443 VTAIL.n98 VTAIL.n97 9.3005
R1444 VTAIL.n100 VTAIL.n99 9.3005
R1445 VTAIL.n78 VTAIL.n77 9.3005
R1446 VTAIL.n106 VTAIL.n105 9.3005
R1447 VTAIL.n108 VTAIL.n107 9.3005
R1448 VTAIL.n123 VTAIL.n122 9.3005
R1449 VTAIL.n70 VTAIL.n69 9.3005
R1450 VTAIL.n117 VTAIL.n116 9.3005
R1451 VTAIL.n115 VTAIL.n114 9.3005
R1452 VTAIL.n74 VTAIL.n73 9.3005
R1453 VTAIL.n212 VTAIL.n202 8.92171
R1454 VTAIL.n26 VTAIL.n16 8.92171
R1455 VTAIL.n155 VTAIL.n145 8.92171
R1456 VTAIL.n93 VTAIL.n83 8.92171
R1457 VTAIL.n211 VTAIL.n204 8.14595
R1458 VTAIL.n25 VTAIL.n18 8.14595
R1459 VTAIL.n154 VTAIL.n147 8.14595
R1460 VTAIL.n92 VTAIL.n85 8.14595
R1461 VTAIL.n208 VTAIL.n207 7.3702
R1462 VTAIL.n22 VTAIL.n21 7.3702
R1463 VTAIL.n151 VTAIL.n150 7.3702
R1464 VTAIL.n89 VTAIL.n88 7.3702
R1465 VTAIL.n208 VTAIL.n204 5.81868
R1466 VTAIL.n22 VTAIL.n18 5.81868
R1467 VTAIL.n151 VTAIL.n147 5.81868
R1468 VTAIL.n89 VTAIL.n85 5.81868
R1469 VTAIL.n212 VTAIL.n211 5.04292
R1470 VTAIL.n26 VTAIL.n25 5.04292
R1471 VTAIL.n155 VTAIL.n154 5.04292
R1472 VTAIL.n93 VTAIL.n92 5.04292
R1473 VTAIL.n215 VTAIL.n202 4.26717
R1474 VTAIL.n244 VTAIL.n188 4.26717
R1475 VTAIL.n29 VTAIL.n16 4.26717
R1476 VTAIL.n58 VTAIL.n2 4.26717
R1477 VTAIL.n186 VTAIL.n130 4.26717
R1478 VTAIL.n158 VTAIL.n145 4.26717
R1479 VTAIL.n124 VTAIL.n68 4.26717
R1480 VTAIL.n96 VTAIL.n83 4.26717
R1481 VTAIL.n216 VTAIL.n200 3.49141
R1482 VTAIL.n242 VTAIL.n241 3.49141
R1483 VTAIL.n30 VTAIL.n14 3.49141
R1484 VTAIL.n56 VTAIL.n55 3.49141
R1485 VTAIL.n184 VTAIL.n183 3.49141
R1486 VTAIL.n159 VTAIL.n143 3.49141
R1487 VTAIL.n122 VTAIL.n121 3.49141
R1488 VTAIL.n97 VTAIL.n81 3.49141
R1489 VTAIL.n246 VTAIL.t2 3.00466
R1490 VTAIL.n246 VTAIL.t6 3.00466
R1491 VTAIL.n0 VTAIL.t1 3.00466
R1492 VTAIL.n0 VTAIL.t4 3.00466
R1493 VTAIL.n60 VTAIL.t11 3.00466
R1494 VTAIL.n60 VTAIL.t12 3.00466
R1495 VTAIL.n62 VTAIL.t17 3.00466
R1496 VTAIL.n62 VTAIL.t14 3.00466
R1497 VTAIL.n128 VTAIL.t13 3.00466
R1498 VTAIL.n128 VTAIL.t19 3.00466
R1499 VTAIL.n126 VTAIL.t16 3.00466
R1500 VTAIL.n126 VTAIL.t10 3.00466
R1501 VTAIL.n66 VTAIL.t9 3.00466
R1502 VTAIL.n66 VTAIL.t0 3.00466
R1503 VTAIL.n64 VTAIL.t3 3.00466
R1504 VTAIL.n64 VTAIL.t8 3.00466
R1505 VTAIL.n220 VTAIL.n219 2.71565
R1506 VTAIL.n238 VTAIL.n190 2.71565
R1507 VTAIL.n34 VTAIL.n33 2.71565
R1508 VTAIL.n52 VTAIL.n4 2.71565
R1509 VTAIL.n180 VTAIL.n132 2.71565
R1510 VTAIL.n163 VTAIL.n162 2.71565
R1511 VTAIL.n118 VTAIL.n70 2.71565
R1512 VTAIL.n101 VTAIL.n100 2.71565
R1513 VTAIL.n209 VTAIL.n205 2.41282
R1514 VTAIL.n23 VTAIL.n19 2.41282
R1515 VTAIL.n152 VTAIL.n148 2.41282
R1516 VTAIL.n90 VTAIL.n86 2.41282
R1517 VTAIL.n224 VTAIL.n198 1.93989
R1518 VTAIL.n237 VTAIL.n192 1.93989
R1519 VTAIL.n38 VTAIL.n12 1.93989
R1520 VTAIL.n51 VTAIL.n6 1.93989
R1521 VTAIL.n179 VTAIL.n134 1.93989
R1522 VTAIL.n166 VTAIL.n140 1.93989
R1523 VTAIL.n117 VTAIL.n72 1.93989
R1524 VTAIL.n104 VTAIL.n78 1.93989
R1525 VTAIL.n67 VTAIL.n65 1.88843
R1526 VTAIL.n125 VTAIL.n67 1.88843
R1527 VTAIL.n129 VTAIL.n127 1.88843
R1528 VTAIL.n187 VTAIL.n129 1.88843
R1529 VTAIL.n63 VTAIL.n61 1.88843
R1530 VTAIL.n61 VTAIL.n59 1.88843
R1531 VTAIL.n247 VTAIL.n245 1.88843
R1532 VTAIL VTAIL.n1 1.47464
R1533 VTAIL.n127 VTAIL.n125 1.41429
R1534 VTAIL.n59 VTAIL.n1 1.41429
R1535 VTAIL.n225 VTAIL.n196 1.16414
R1536 VTAIL.n234 VTAIL.n233 1.16414
R1537 VTAIL.n39 VTAIL.n10 1.16414
R1538 VTAIL.n48 VTAIL.n47 1.16414
R1539 VTAIL.n176 VTAIL.n175 1.16414
R1540 VTAIL.n167 VTAIL.n138 1.16414
R1541 VTAIL.n114 VTAIL.n113 1.16414
R1542 VTAIL.n105 VTAIL.n76 1.16414
R1543 VTAIL VTAIL.n247 0.414293
R1544 VTAIL.n229 VTAIL.n228 0.388379
R1545 VTAIL.n230 VTAIL.n194 0.388379
R1546 VTAIL.n43 VTAIL.n42 0.388379
R1547 VTAIL.n44 VTAIL.n8 0.388379
R1548 VTAIL.n172 VTAIL.n136 0.388379
R1549 VTAIL.n171 VTAIL.n170 0.388379
R1550 VTAIL.n110 VTAIL.n74 0.388379
R1551 VTAIL.n109 VTAIL.n108 0.388379
R1552 VTAIL.n210 VTAIL.n209 0.155672
R1553 VTAIL.n210 VTAIL.n201 0.155672
R1554 VTAIL.n217 VTAIL.n201 0.155672
R1555 VTAIL.n218 VTAIL.n217 0.155672
R1556 VTAIL.n218 VTAIL.n197 0.155672
R1557 VTAIL.n226 VTAIL.n197 0.155672
R1558 VTAIL.n227 VTAIL.n226 0.155672
R1559 VTAIL.n227 VTAIL.n193 0.155672
R1560 VTAIL.n235 VTAIL.n193 0.155672
R1561 VTAIL.n236 VTAIL.n235 0.155672
R1562 VTAIL.n236 VTAIL.n189 0.155672
R1563 VTAIL.n243 VTAIL.n189 0.155672
R1564 VTAIL.n24 VTAIL.n23 0.155672
R1565 VTAIL.n24 VTAIL.n15 0.155672
R1566 VTAIL.n31 VTAIL.n15 0.155672
R1567 VTAIL.n32 VTAIL.n31 0.155672
R1568 VTAIL.n32 VTAIL.n11 0.155672
R1569 VTAIL.n40 VTAIL.n11 0.155672
R1570 VTAIL.n41 VTAIL.n40 0.155672
R1571 VTAIL.n41 VTAIL.n7 0.155672
R1572 VTAIL.n49 VTAIL.n7 0.155672
R1573 VTAIL.n50 VTAIL.n49 0.155672
R1574 VTAIL.n50 VTAIL.n3 0.155672
R1575 VTAIL.n57 VTAIL.n3 0.155672
R1576 VTAIL.n185 VTAIL.n131 0.155672
R1577 VTAIL.n178 VTAIL.n131 0.155672
R1578 VTAIL.n178 VTAIL.n177 0.155672
R1579 VTAIL.n177 VTAIL.n135 0.155672
R1580 VTAIL.n169 VTAIL.n135 0.155672
R1581 VTAIL.n169 VTAIL.n168 0.155672
R1582 VTAIL.n168 VTAIL.n139 0.155672
R1583 VTAIL.n161 VTAIL.n139 0.155672
R1584 VTAIL.n161 VTAIL.n160 0.155672
R1585 VTAIL.n160 VTAIL.n144 0.155672
R1586 VTAIL.n153 VTAIL.n144 0.155672
R1587 VTAIL.n153 VTAIL.n152 0.155672
R1588 VTAIL.n123 VTAIL.n69 0.155672
R1589 VTAIL.n116 VTAIL.n69 0.155672
R1590 VTAIL.n116 VTAIL.n115 0.155672
R1591 VTAIL.n115 VTAIL.n73 0.155672
R1592 VTAIL.n107 VTAIL.n73 0.155672
R1593 VTAIL.n107 VTAIL.n106 0.155672
R1594 VTAIL.n106 VTAIL.n77 0.155672
R1595 VTAIL.n99 VTAIL.n77 0.155672
R1596 VTAIL.n99 VTAIL.n98 0.155672
R1597 VTAIL.n98 VTAIL.n82 0.155672
R1598 VTAIL.n91 VTAIL.n82 0.155672
R1599 VTAIL.n91 VTAIL.n90 0.155672
R1600 VDD1.n52 VDD1.n0 756.745
R1601 VDD1.n111 VDD1.n59 756.745
R1602 VDD1.n53 VDD1.n52 585
R1603 VDD1.n51 VDD1.n50 585
R1604 VDD1.n4 VDD1.n3 585
R1605 VDD1.n45 VDD1.n44 585
R1606 VDD1.n43 VDD1.n42 585
R1607 VDD1.n41 VDD1.n7 585
R1608 VDD1.n11 VDD1.n8 585
R1609 VDD1.n36 VDD1.n35 585
R1610 VDD1.n34 VDD1.n33 585
R1611 VDD1.n13 VDD1.n12 585
R1612 VDD1.n28 VDD1.n27 585
R1613 VDD1.n26 VDD1.n25 585
R1614 VDD1.n17 VDD1.n16 585
R1615 VDD1.n20 VDD1.n19 585
R1616 VDD1.n78 VDD1.n77 585
R1617 VDD1.n75 VDD1.n74 585
R1618 VDD1.n84 VDD1.n83 585
R1619 VDD1.n86 VDD1.n85 585
R1620 VDD1.n71 VDD1.n70 585
R1621 VDD1.n92 VDD1.n91 585
R1622 VDD1.n95 VDD1.n94 585
R1623 VDD1.n93 VDD1.n67 585
R1624 VDD1.n100 VDD1.n66 585
R1625 VDD1.n102 VDD1.n101 585
R1626 VDD1.n104 VDD1.n103 585
R1627 VDD1.n63 VDD1.n62 585
R1628 VDD1.n110 VDD1.n109 585
R1629 VDD1.n112 VDD1.n111 585
R1630 VDD1.t6 VDD1.n18 329.038
R1631 VDD1.t3 VDD1.n76 329.038
R1632 VDD1.n52 VDD1.n51 171.744
R1633 VDD1.n51 VDD1.n3 171.744
R1634 VDD1.n44 VDD1.n3 171.744
R1635 VDD1.n44 VDD1.n43 171.744
R1636 VDD1.n43 VDD1.n7 171.744
R1637 VDD1.n11 VDD1.n7 171.744
R1638 VDD1.n35 VDD1.n11 171.744
R1639 VDD1.n35 VDD1.n34 171.744
R1640 VDD1.n34 VDD1.n12 171.744
R1641 VDD1.n27 VDD1.n12 171.744
R1642 VDD1.n27 VDD1.n26 171.744
R1643 VDD1.n26 VDD1.n16 171.744
R1644 VDD1.n19 VDD1.n16 171.744
R1645 VDD1.n77 VDD1.n74 171.744
R1646 VDD1.n84 VDD1.n74 171.744
R1647 VDD1.n85 VDD1.n84 171.744
R1648 VDD1.n85 VDD1.n70 171.744
R1649 VDD1.n92 VDD1.n70 171.744
R1650 VDD1.n94 VDD1.n92 171.744
R1651 VDD1.n94 VDD1.n93 171.744
R1652 VDD1.n93 VDD1.n66 171.744
R1653 VDD1.n102 VDD1.n66 171.744
R1654 VDD1.n103 VDD1.n102 171.744
R1655 VDD1.n103 VDD1.n62 171.744
R1656 VDD1.n110 VDD1.n62 171.744
R1657 VDD1.n111 VDD1.n110 171.744
R1658 VDD1.n19 VDD1.t6 85.8723
R1659 VDD1.n77 VDD1.t3 85.8723
R1660 VDD1.n119 VDD1.n118 79.9417
R1661 VDD1.n58 VDD1.n57 78.5813
R1662 VDD1.n121 VDD1.n120 78.5811
R1663 VDD1.n117 VDD1.n116 78.5811
R1664 VDD1.n58 VDD1.n56 53.4672
R1665 VDD1.n117 VDD1.n115 53.4672
R1666 VDD1.n121 VDD1.n119 43.5375
R1667 VDD1.n42 VDD1.n41 13.1884
R1668 VDD1.n101 VDD1.n100 13.1884
R1669 VDD1.n45 VDD1.n6 12.8005
R1670 VDD1.n40 VDD1.n8 12.8005
R1671 VDD1.n99 VDD1.n67 12.8005
R1672 VDD1.n104 VDD1.n65 12.8005
R1673 VDD1.n46 VDD1.n4 12.0247
R1674 VDD1.n37 VDD1.n36 12.0247
R1675 VDD1.n96 VDD1.n95 12.0247
R1676 VDD1.n105 VDD1.n63 12.0247
R1677 VDD1.n50 VDD1.n49 11.249
R1678 VDD1.n33 VDD1.n10 11.249
R1679 VDD1.n91 VDD1.n69 11.249
R1680 VDD1.n109 VDD1.n108 11.249
R1681 VDD1.n20 VDD1.n18 10.7239
R1682 VDD1.n78 VDD1.n76 10.7239
R1683 VDD1.n53 VDD1.n2 10.4732
R1684 VDD1.n32 VDD1.n13 10.4732
R1685 VDD1.n90 VDD1.n71 10.4732
R1686 VDD1.n112 VDD1.n61 10.4732
R1687 VDD1.n54 VDD1.n0 9.69747
R1688 VDD1.n29 VDD1.n28 9.69747
R1689 VDD1.n87 VDD1.n86 9.69747
R1690 VDD1.n113 VDD1.n59 9.69747
R1691 VDD1.n56 VDD1.n55 9.45567
R1692 VDD1.n115 VDD1.n114 9.45567
R1693 VDD1.n22 VDD1.n21 9.3005
R1694 VDD1.n24 VDD1.n23 9.3005
R1695 VDD1.n15 VDD1.n14 9.3005
R1696 VDD1.n30 VDD1.n29 9.3005
R1697 VDD1.n32 VDD1.n31 9.3005
R1698 VDD1.n10 VDD1.n9 9.3005
R1699 VDD1.n38 VDD1.n37 9.3005
R1700 VDD1.n40 VDD1.n39 9.3005
R1701 VDD1.n55 VDD1.n54 9.3005
R1702 VDD1.n2 VDD1.n1 9.3005
R1703 VDD1.n49 VDD1.n48 9.3005
R1704 VDD1.n47 VDD1.n46 9.3005
R1705 VDD1.n6 VDD1.n5 9.3005
R1706 VDD1.n114 VDD1.n113 9.3005
R1707 VDD1.n61 VDD1.n60 9.3005
R1708 VDD1.n108 VDD1.n107 9.3005
R1709 VDD1.n106 VDD1.n105 9.3005
R1710 VDD1.n65 VDD1.n64 9.3005
R1711 VDD1.n80 VDD1.n79 9.3005
R1712 VDD1.n82 VDD1.n81 9.3005
R1713 VDD1.n73 VDD1.n72 9.3005
R1714 VDD1.n88 VDD1.n87 9.3005
R1715 VDD1.n90 VDD1.n89 9.3005
R1716 VDD1.n69 VDD1.n68 9.3005
R1717 VDD1.n97 VDD1.n96 9.3005
R1718 VDD1.n99 VDD1.n98 9.3005
R1719 VDD1.n25 VDD1.n15 8.92171
R1720 VDD1.n83 VDD1.n73 8.92171
R1721 VDD1.n24 VDD1.n17 8.14595
R1722 VDD1.n82 VDD1.n75 8.14595
R1723 VDD1.n21 VDD1.n20 7.3702
R1724 VDD1.n79 VDD1.n78 7.3702
R1725 VDD1.n21 VDD1.n17 5.81868
R1726 VDD1.n79 VDD1.n75 5.81868
R1727 VDD1.n25 VDD1.n24 5.04292
R1728 VDD1.n83 VDD1.n82 5.04292
R1729 VDD1.n56 VDD1.n0 4.26717
R1730 VDD1.n28 VDD1.n15 4.26717
R1731 VDD1.n86 VDD1.n73 4.26717
R1732 VDD1.n115 VDD1.n59 4.26717
R1733 VDD1.n54 VDD1.n53 3.49141
R1734 VDD1.n29 VDD1.n13 3.49141
R1735 VDD1.n87 VDD1.n71 3.49141
R1736 VDD1.n113 VDD1.n112 3.49141
R1737 VDD1.n120 VDD1.t1 3.00466
R1738 VDD1.n120 VDD1.t0 3.00466
R1739 VDD1.n57 VDD1.t2 3.00466
R1740 VDD1.n57 VDD1.t9 3.00466
R1741 VDD1.n118 VDD1.t4 3.00466
R1742 VDD1.n118 VDD1.t7 3.00466
R1743 VDD1.n116 VDD1.t5 3.00466
R1744 VDD1.n116 VDD1.t8 3.00466
R1745 VDD1.n50 VDD1.n2 2.71565
R1746 VDD1.n33 VDD1.n32 2.71565
R1747 VDD1.n91 VDD1.n90 2.71565
R1748 VDD1.n109 VDD1.n61 2.71565
R1749 VDD1.n22 VDD1.n18 2.41282
R1750 VDD1.n80 VDD1.n76 2.41282
R1751 VDD1.n49 VDD1.n4 1.93989
R1752 VDD1.n36 VDD1.n10 1.93989
R1753 VDD1.n95 VDD1.n69 1.93989
R1754 VDD1.n108 VDD1.n63 1.93989
R1755 VDD1 VDD1.n121 1.35826
R1756 VDD1.n46 VDD1.n45 1.16414
R1757 VDD1.n37 VDD1.n8 1.16414
R1758 VDD1.n96 VDD1.n67 1.16414
R1759 VDD1.n105 VDD1.n104 1.16414
R1760 VDD1 VDD1.n58 0.530672
R1761 VDD1.n119 VDD1.n117 0.417137
R1762 VDD1.n42 VDD1.n6 0.388379
R1763 VDD1.n41 VDD1.n40 0.388379
R1764 VDD1.n100 VDD1.n99 0.388379
R1765 VDD1.n101 VDD1.n65 0.388379
R1766 VDD1.n55 VDD1.n1 0.155672
R1767 VDD1.n48 VDD1.n1 0.155672
R1768 VDD1.n48 VDD1.n47 0.155672
R1769 VDD1.n47 VDD1.n5 0.155672
R1770 VDD1.n39 VDD1.n5 0.155672
R1771 VDD1.n39 VDD1.n38 0.155672
R1772 VDD1.n38 VDD1.n9 0.155672
R1773 VDD1.n31 VDD1.n9 0.155672
R1774 VDD1.n31 VDD1.n30 0.155672
R1775 VDD1.n30 VDD1.n14 0.155672
R1776 VDD1.n23 VDD1.n14 0.155672
R1777 VDD1.n23 VDD1.n22 0.155672
R1778 VDD1.n81 VDD1.n80 0.155672
R1779 VDD1.n81 VDD1.n72 0.155672
R1780 VDD1.n88 VDD1.n72 0.155672
R1781 VDD1.n89 VDD1.n88 0.155672
R1782 VDD1.n89 VDD1.n68 0.155672
R1783 VDD1.n97 VDD1.n68 0.155672
R1784 VDD1.n98 VDD1.n97 0.155672
R1785 VDD1.n98 VDD1.n64 0.155672
R1786 VDD1.n106 VDD1.n64 0.155672
R1787 VDD1.n107 VDD1.n106 0.155672
R1788 VDD1.n107 VDD1.n60 0.155672
R1789 VDD1.n114 VDD1.n60 0.155672
R1790 VN.n7 VN.t1 170.185
R1791 VN.n38 VN.t2 170.185
R1792 VN.n59 VN.n31 161.3
R1793 VN.n58 VN.n57 161.3
R1794 VN.n56 VN.n32 161.3
R1795 VN.n55 VN.n54 161.3
R1796 VN.n52 VN.n33 161.3
R1797 VN.n51 VN.n50 161.3
R1798 VN.n49 VN.n34 161.3
R1799 VN.n48 VN.n47 161.3
R1800 VN.n46 VN.n35 161.3
R1801 VN.n45 VN.n44 161.3
R1802 VN.n43 VN.n36 161.3
R1803 VN.n42 VN.n41 161.3
R1804 VN.n40 VN.n37 161.3
R1805 VN.n28 VN.n0 161.3
R1806 VN.n27 VN.n26 161.3
R1807 VN.n25 VN.n1 161.3
R1808 VN.n24 VN.n23 161.3
R1809 VN.n21 VN.n2 161.3
R1810 VN.n20 VN.n19 161.3
R1811 VN.n18 VN.n3 161.3
R1812 VN.n17 VN.n16 161.3
R1813 VN.n15 VN.n4 161.3
R1814 VN.n14 VN.n13 161.3
R1815 VN.n12 VN.n5 161.3
R1816 VN.n11 VN.n10 161.3
R1817 VN.n9 VN.n6 161.3
R1818 VN.n15 VN.t9 140.196
R1819 VN.n8 VN.t3 140.196
R1820 VN.n22 VN.t5 140.196
R1821 VN.n29 VN.t7 140.196
R1822 VN.n46 VN.t6 140.196
R1823 VN.n39 VN.t8 140.196
R1824 VN.n53 VN.t0 140.196
R1825 VN.n60 VN.t4 140.196
R1826 VN.n30 VN.n29 92.1052
R1827 VN.n61 VN.n60 92.1052
R1828 VN.n8 VN.n7 60.1448
R1829 VN.n39 VN.n38 60.1448
R1830 VN.n27 VN.n1 56.4773
R1831 VN.n58 VN.n32 56.4773
R1832 VN.n10 VN.n5 49.6611
R1833 VN.n20 VN.n3 49.6611
R1834 VN.n41 VN.n36 49.6611
R1835 VN.n51 VN.n34 49.6611
R1836 VN VN.n61 48.4489
R1837 VN.n14 VN.n5 31.1601
R1838 VN.n16 VN.n3 31.1601
R1839 VN.n45 VN.n36 31.1601
R1840 VN.n47 VN.n34 31.1601
R1841 VN.n10 VN.n9 24.3439
R1842 VN.n15 VN.n14 24.3439
R1843 VN.n16 VN.n15 24.3439
R1844 VN.n21 VN.n20 24.3439
R1845 VN.n23 VN.n1 24.3439
R1846 VN.n28 VN.n27 24.3439
R1847 VN.n41 VN.n40 24.3439
R1848 VN.n47 VN.n46 24.3439
R1849 VN.n46 VN.n45 24.3439
R1850 VN.n54 VN.n32 24.3439
R1851 VN.n52 VN.n51 24.3439
R1852 VN.n59 VN.n58 24.3439
R1853 VN.n29 VN.n28 18.5015
R1854 VN.n60 VN.n59 18.5015
R1855 VN.n23 VN.n22 15.0934
R1856 VN.n54 VN.n53 15.0934
R1857 VN.n38 VN.n37 13.5258
R1858 VN.n7 VN.n6 13.5258
R1859 VN.n9 VN.n8 9.251
R1860 VN.n22 VN.n21 9.251
R1861 VN.n40 VN.n39 9.251
R1862 VN.n53 VN.n52 9.251
R1863 VN.n61 VN.n31 0.278398
R1864 VN.n30 VN.n0 0.278398
R1865 VN.n57 VN.n31 0.189894
R1866 VN.n57 VN.n56 0.189894
R1867 VN.n56 VN.n55 0.189894
R1868 VN.n55 VN.n33 0.189894
R1869 VN.n50 VN.n33 0.189894
R1870 VN.n50 VN.n49 0.189894
R1871 VN.n49 VN.n48 0.189894
R1872 VN.n48 VN.n35 0.189894
R1873 VN.n44 VN.n35 0.189894
R1874 VN.n44 VN.n43 0.189894
R1875 VN.n43 VN.n42 0.189894
R1876 VN.n42 VN.n37 0.189894
R1877 VN.n11 VN.n6 0.189894
R1878 VN.n12 VN.n11 0.189894
R1879 VN.n13 VN.n12 0.189894
R1880 VN.n13 VN.n4 0.189894
R1881 VN.n17 VN.n4 0.189894
R1882 VN.n18 VN.n17 0.189894
R1883 VN.n19 VN.n18 0.189894
R1884 VN.n19 VN.n2 0.189894
R1885 VN.n24 VN.n2 0.189894
R1886 VN.n25 VN.n24 0.189894
R1887 VN.n26 VN.n25 0.189894
R1888 VN.n26 VN.n0 0.189894
R1889 VN VN.n30 0.153422
R1890 VDD2.n113 VDD2.n61 756.745
R1891 VDD2.n52 VDD2.n0 756.745
R1892 VDD2.n114 VDD2.n113 585
R1893 VDD2.n112 VDD2.n111 585
R1894 VDD2.n65 VDD2.n64 585
R1895 VDD2.n106 VDD2.n105 585
R1896 VDD2.n104 VDD2.n103 585
R1897 VDD2.n102 VDD2.n68 585
R1898 VDD2.n72 VDD2.n69 585
R1899 VDD2.n97 VDD2.n96 585
R1900 VDD2.n95 VDD2.n94 585
R1901 VDD2.n74 VDD2.n73 585
R1902 VDD2.n89 VDD2.n88 585
R1903 VDD2.n87 VDD2.n86 585
R1904 VDD2.n78 VDD2.n77 585
R1905 VDD2.n81 VDD2.n80 585
R1906 VDD2.n19 VDD2.n18 585
R1907 VDD2.n16 VDD2.n15 585
R1908 VDD2.n25 VDD2.n24 585
R1909 VDD2.n27 VDD2.n26 585
R1910 VDD2.n12 VDD2.n11 585
R1911 VDD2.n33 VDD2.n32 585
R1912 VDD2.n36 VDD2.n35 585
R1913 VDD2.n34 VDD2.n8 585
R1914 VDD2.n41 VDD2.n7 585
R1915 VDD2.n43 VDD2.n42 585
R1916 VDD2.n45 VDD2.n44 585
R1917 VDD2.n4 VDD2.n3 585
R1918 VDD2.n51 VDD2.n50 585
R1919 VDD2.n53 VDD2.n52 585
R1920 VDD2.t5 VDD2.n79 329.038
R1921 VDD2.t8 VDD2.n17 329.038
R1922 VDD2.n113 VDD2.n112 171.744
R1923 VDD2.n112 VDD2.n64 171.744
R1924 VDD2.n105 VDD2.n64 171.744
R1925 VDD2.n105 VDD2.n104 171.744
R1926 VDD2.n104 VDD2.n68 171.744
R1927 VDD2.n72 VDD2.n68 171.744
R1928 VDD2.n96 VDD2.n72 171.744
R1929 VDD2.n96 VDD2.n95 171.744
R1930 VDD2.n95 VDD2.n73 171.744
R1931 VDD2.n88 VDD2.n73 171.744
R1932 VDD2.n88 VDD2.n87 171.744
R1933 VDD2.n87 VDD2.n77 171.744
R1934 VDD2.n80 VDD2.n77 171.744
R1935 VDD2.n18 VDD2.n15 171.744
R1936 VDD2.n25 VDD2.n15 171.744
R1937 VDD2.n26 VDD2.n25 171.744
R1938 VDD2.n26 VDD2.n11 171.744
R1939 VDD2.n33 VDD2.n11 171.744
R1940 VDD2.n35 VDD2.n33 171.744
R1941 VDD2.n35 VDD2.n34 171.744
R1942 VDD2.n34 VDD2.n7 171.744
R1943 VDD2.n43 VDD2.n7 171.744
R1944 VDD2.n44 VDD2.n43 171.744
R1945 VDD2.n44 VDD2.n3 171.744
R1946 VDD2.n51 VDD2.n3 171.744
R1947 VDD2.n52 VDD2.n51 171.744
R1948 VDD2.n80 VDD2.t5 85.8723
R1949 VDD2.n18 VDD2.t8 85.8723
R1950 VDD2.n60 VDD2.n59 79.9417
R1951 VDD2 VDD2.n121 79.9389
R1952 VDD2.n120 VDD2.n119 78.5813
R1953 VDD2.n58 VDD2.n57 78.5811
R1954 VDD2.n58 VDD2.n56 53.4672
R1955 VDD2.n118 VDD2.n117 51.5793
R1956 VDD2.n118 VDD2.n60 42.0106
R1957 VDD2.n103 VDD2.n102 13.1884
R1958 VDD2.n42 VDD2.n41 13.1884
R1959 VDD2.n106 VDD2.n67 12.8005
R1960 VDD2.n101 VDD2.n69 12.8005
R1961 VDD2.n40 VDD2.n8 12.8005
R1962 VDD2.n45 VDD2.n6 12.8005
R1963 VDD2.n107 VDD2.n65 12.0247
R1964 VDD2.n98 VDD2.n97 12.0247
R1965 VDD2.n37 VDD2.n36 12.0247
R1966 VDD2.n46 VDD2.n4 12.0247
R1967 VDD2.n111 VDD2.n110 11.249
R1968 VDD2.n94 VDD2.n71 11.249
R1969 VDD2.n32 VDD2.n10 11.249
R1970 VDD2.n50 VDD2.n49 11.249
R1971 VDD2.n81 VDD2.n79 10.7239
R1972 VDD2.n19 VDD2.n17 10.7239
R1973 VDD2.n114 VDD2.n63 10.4732
R1974 VDD2.n93 VDD2.n74 10.4732
R1975 VDD2.n31 VDD2.n12 10.4732
R1976 VDD2.n53 VDD2.n2 10.4732
R1977 VDD2.n115 VDD2.n61 9.69747
R1978 VDD2.n90 VDD2.n89 9.69747
R1979 VDD2.n28 VDD2.n27 9.69747
R1980 VDD2.n54 VDD2.n0 9.69747
R1981 VDD2.n117 VDD2.n116 9.45567
R1982 VDD2.n56 VDD2.n55 9.45567
R1983 VDD2.n83 VDD2.n82 9.3005
R1984 VDD2.n85 VDD2.n84 9.3005
R1985 VDD2.n76 VDD2.n75 9.3005
R1986 VDD2.n91 VDD2.n90 9.3005
R1987 VDD2.n93 VDD2.n92 9.3005
R1988 VDD2.n71 VDD2.n70 9.3005
R1989 VDD2.n99 VDD2.n98 9.3005
R1990 VDD2.n101 VDD2.n100 9.3005
R1991 VDD2.n116 VDD2.n115 9.3005
R1992 VDD2.n63 VDD2.n62 9.3005
R1993 VDD2.n110 VDD2.n109 9.3005
R1994 VDD2.n108 VDD2.n107 9.3005
R1995 VDD2.n67 VDD2.n66 9.3005
R1996 VDD2.n55 VDD2.n54 9.3005
R1997 VDD2.n2 VDD2.n1 9.3005
R1998 VDD2.n49 VDD2.n48 9.3005
R1999 VDD2.n47 VDD2.n46 9.3005
R2000 VDD2.n6 VDD2.n5 9.3005
R2001 VDD2.n21 VDD2.n20 9.3005
R2002 VDD2.n23 VDD2.n22 9.3005
R2003 VDD2.n14 VDD2.n13 9.3005
R2004 VDD2.n29 VDD2.n28 9.3005
R2005 VDD2.n31 VDD2.n30 9.3005
R2006 VDD2.n10 VDD2.n9 9.3005
R2007 VDD2.n38 VDD2.n37 9.3005
R2008 VDD2.n40 VDD2.n39 9.3005
R2009 VDD2.n86 VDD2.n76 8.92171
R2010 VDD2.n24 VDD2.n14 8.92171
R2011 VDD2.n85 VDD2.n78 8.14595
R2012 VDD2.n23 VDD2.n16 8.14595
R2013 VDD2.n82 VDD2.n81 7.3702
R2014 VDD2.n20 VDD2.n19 7.3702
R2015 VDD2.n82 VDD2.n78 5.81868
R2016 VDD2.n20 VDD2.n16 5.81868
R2017 VDD2.n86 VDD2.n85 5.04292
R2018 VDD2.n24 VDD2.n23 5.04292
R2019 VDD2.n117 VDD2.n61 4.26717
R2020 VDD2.n89 VDD2.n76 4.26717
R2021 VDD2.n27 VDD2.n14 4.26717
R2022 VDD2.n56 VDD2.n0 4.26717
R2023 VDD2.n115 VDD2.n114 3.49141
R2024 VDD2.n90 VDD2.n74 3.49141
R2025 VDD2.n28 VDD2.n12 3.49141
R2026 VDD2.n54 VDD2.n53 3.49141
R2027 VDD2.n121 VDD2.t1 3.00466
R2028 VDD2.n121 VDD2.t7 3.00466
R2029 VDD2.n119 VDD2.t9 3.00466
R2030 VDD2.n119 VDD2.t3 3.00466
R2031 VDD2.n59 VDD2.t4 3.00466
R2032 VDD2.n59 VDD2.t2 3.00466
R2033 VDD2.n57 VDD2.t6 3.00466
R2034 VDD2.n57 VDD2.t0 3.00466
R2035 VDD2.n111 VDD2.n63 2.71565
R2036 VDD2.n94 VDD2.n93 2.71565
R2037 VDD2.n32 VDD2.n31 2.71565
R2038 VDD2.n50 VDD2.n2 2.71565
R2039 VDD2.n83 VDD2.n79 2.41282
R2040 VDD2.n21 VDD2.n17 2.41282
R2041 VDD2.n110 VDD2.n65 1.93989
R2042 VDD2.n97 VDD2.n71 1.93989
R2043 VDD2.n36 VDD2.n10 1.93989
R2044 VDD2.n49 VDD2.n4 1.93989
R2045 VDD2.n120 VDD2.n118 1.88843
R2046 VDD2.n107 VDD2.n106 1.16414
R2047 VDD2.n98 VDD2.n69 1.16414
R2048 VDD2.n37 VDD2.n8 1.16414
R2049 VDD2.n46 VDD2.n45 1.16414
R2050 VDD2 VDD2.n120 0.530672
R2051 VDD2.n60 VDD2.n58 0.417137
R2052 VDD2.n103 VDD2.n67 0.388379
R2053 VDD2.n102 VDD2.n101 0.388379
R2054 VDD2.n41 VDD2.n40 0.388379
R2055 VDD2.n42 VDD2.n6 0.388379
R2056 VDD2.n116 VDD2.n62 0.155672
R2057 VDD2.n109 VDD2.n62 0.155672
R2058 VDD2.n109 VDD2.n108 0.155672
R2059 VDD2.n108 VDD2.n66 0.155672
R2060 VDD2.n100 VDD2.n66 0.155672
R2061 VDD2.n100 VDD2.n99 0.155672
R2062 VDD2.n99 VDD2.n70 0.155672
R2063 VDD2.n92 VDD2.n70 0.155672
R2064 VDD2.n92 VDD2.n91 0.155672
R2065 VDD2.n91 VDD2.n75 0.155672
R2066 VDD2.n84 VDD2.n75 0.155672
R2067 VDD2.n84 VDD2.n83 0.155672
R2068 VDD2.n22 VDD2.n21 0.155672
R2069 VDD2.n22 VDD2.n13 0.155672
R2070 VDD2.n29 VDD2.n13 0.155672
R2071 VDD2.n30 VDD2.n29 0.155672
R2072 VDD2.n30 VDD2.n9 0.155672
R2073 VDD2.n38 VDD2.n9 0.155672
R2074 VDD2.n39 VDD2.n38 0.155672
R2075 VDD2.n39 VDD2.n5 0.155672
R2076 VDD2.n47 VDD2.n5 0.155672
R2077 VDD2.n48 VDD2.n47 0.155672
R2078 VDD2.n48 VDD2.n1 0.155672
R2079 VDD2.n55 VDD2.n1 0.155672
C0 VN VDD2 8.94099f
C1 VDD1 VDD2 1.69297f
C2 VTAIL VN 9.32573f
C3 VDD1 VTAIL 9.87772f
C4 B VDD2 2.18533f
C5 B VTAIL 3.15002f
C6 VDD2 VP 0.488796f
C7 VTAIL VP 9.340071f
C8 VDD1 VN 0.15135f
C9 VDD2 w_n3598_n3132# 2.52933f
C10 VTAIL w_n3598_n3132# 2.94888f
C11 B VN 1.07802f
C12 B VDD1 2.09623f
C13 VN VP 7.0993f
C14 VDD1 VP 9.27475f
C15 B VP 1.85781f
C16 VN w_n3598_n3132# 7.46846f
C17 VDD1 w_n3598_n3132# 2.42414f
C18 VTAIL VDD2 9.923079f
C19 B w_n3598_n3132# 8.97159f
C20 VP w_n3598_n3132# 7.93462f
C21 VDD2 VSUBS 1.81002f
C22 VDD1 VSUBS 1.614016f
C23 VTAIL VSUBS 1.086049f
C24 VN VSUBS 6.44494f
C25 VP VSUBS 3.255373f
C26 B VSUBS 4.348561f
C27 w_n3598_n3132# VSUBS 0.138984p
C28 VDD2.n0 VSUBS 0.03111f
C29 VDD2.n1 VSUBS 0.027776f
C30 VDD2.n2 VSUBS 0.014925f
C31 VDD2.n3 VSUBS 0.035278f
C32 VDD2.n4 VSUBS 0.015803f
C33 VDD2.n5 VSUBS 0.027776f
C34 VDD2.n6 VSUBS 0.014925f
C35 VDD2.n7 VSUBS 0.035278f
C36 VDD2.n8 VSUBS 0.015803f
C37 VDD2.n9 VSUBS 0.027776f
C38 VDD2.n10 VSUBS 0.014925f
C39 VDD2.n11 VSUBS 0.035278f
C40 VDD2.n12 VSUBS 0.015803f
C41 VDD2.n13 VSUBS 0.027776f
C42 VDD2.n14 VSUBS 0.014925f
C43 VDD2.n15 VSUBS 0.035278f
C44 VDD2.n16 VSUBS 0.015803f
C45 VDD2.n17 VSUBS 0.203942f
C46 VDD2.t8 VSUBS 0.075924f
C47 VDD2.n18 VSUBS 0.026459f
C48 VDD2.n19 VSUBS 0.026538f
C49 VDD2.n20 VSUBS 0.014925f
C50 VDD2.n21 VSUBS 1.22107f
C51 VDD2.n22 VSUBS 0.027776f
C52 VDD2.n23 VSUBS 0.014925f
C53 VDD2.n24 VSUBS 0.015803f
C54 VDD2.n25 VSUBS 0.035278f
C55 VDD2.n26 VSUBS 0.035278f
C56 VDD2.n27 VSUBS 0.015803f
C57 VDD2.n28 VSUBS 0.014925f
C58 VDD2.n29 VSUBS 0.027776f
C59 VDD2.n30 VSUBS 0.027776f
C60 VDD2.n31 VSUBS 0.014925f
C61 VDD2.n32 VSUBS 0.015803f
C62 VDD2.n33 VSUBS 0.035278f
C63 VDD2.n34 VSUBS 0.035278f
C64 VDD2.n35 VSUBS 0.035278f
C65 VDD2.n36 VSUBS 0.015803f
C66 VDD2.n37 VSUBS 0.014925f
C67 VDD2.n38 VSUBS 0.027776f
C68 VDD2.n39 VSUBS 0.027776f
C69 VDD2.n40 VSUBS 0.014925f
C70 VDD2.n41 VSUBS 0.015364f
C71 VDD2.n42 VSUBS 0.015364f
C72 VDD2.n43 VSUBS 0.035278f
C73 VDD2.n44 VSUBS 0.035278f
C74 VDD2.n45 VSUBS 0.015803f
C75 VDD2.n46 VSUBS 0.014925f
C76 VDD2.n47 VSUBS 0.027776f
C77 VDD2.n48 VSUBS 0.027776f
C78 VDD2.n49 VSUBS 0.014925f
C79 VDD2.n50 VSUBS 0.015803f
C80 VDD2.n51 VSUBS 0.035278f
C81 VDD2.n52 VSUBS 0.087415f
C82 VDD2.n53 VSUBS 0.015803f
C83 VDD2.n54 VSUBS 0.014925f
C84 VDD2.n55 VSUBS 0.069514f
C85 VDD2.n56 VSUBS 0.07131f
C86 VDD2.t6 VSUBS 0.237489f
C87 VDD2.t0 VSUBS 0.237489f
C88 VDD2.n57 VSUBS 1.82871f
C89 VDD2.n58 VSUBS 0.927049f
C90 VDD2.t4 VSUBS 0.237489f
C91 VDD2.t2 VSUBS 0.237489f
C92 VDD2.n59 VSUBS 1.84239f
C93 VDD2.n60 VSUBS 2.98749f
C94 VDD2.n61 VSUBS 0.03111f
C95 VDD2.n62 VSUBS 0.027776f
C96 VDD2.n63 VSUBS 0.014925f
C97 VDD2.n64 VSUBS 0.035278f
C98 VDD2.n65 VSUBS 0.015803f
C99 VDD2.n66 VSUBS 0.027776f
C100 VDD2.n67 VSUBS 0.014925f
C101 VDD2.n68 VSUBS 0.035278f
C102 VDD2.n69 VSUBS 0.015803f
C103 VDD2.n70 VSUBS 0.027776f
C104 VDD2.n71 VSUBS 0.014925f
C105 VDD2.n72 VSUBS 0.035278f
C106 VDD2.n73 VSUBS 0.035278f
C107 VDD2.n74 VSUBS 0.015803f
C108 VDD2.n75 VSUBS 0.027776f
C109 VDD2.n76 VSUBS 0.014925f
C110 VDD2.n77 VSUBS 0.035278f
C111 VDD2.n78 VSUBS 0.015803f
C112 VDD2.n79 VSUBS 0.203942f
C113 VDD2.t5 VSUBS 0.075924f
C114 VDD2.n80 VSUBS 0.026459f
C115 VDD2.n81 VSUBS 0.026538f
C116 VDD2.n82 VSUBS 0.014925f
C117 VDD2.n83 VSUBS 1.22107f
C118 VDD2.n84 VSUBS 0.027776f
C119 VDD2.n85 VSUBS 0.014925f
C120 VDD2.n86 VSUBS 0.015803f
C121 VDD2.n87 VSUBS 0.035278f
C122 VDD2.n88 VSUBS 0.035278f
C123 VDD2.n89 VSUBS 0.015803f
C124 VDD2.n90 VSUBS 0.014925f
C125 VDD2.n91 VSUBS 0.027776f
C126 VDD2.n92 VSUBS 0.027776f
C127 VDD2.n93 VSUBS 0.014925f
C128 VDD2.n94 VSUBS 0.015803f
C129 VDD2.n95 VSUBS 0.035278f
C130 VDD2.n96 VSUBS 0.035278f
C131 VDD2.n97 VSUBS 0.015803f
C132 VDD2.n98 VSUBS 0.014925f
C133 VDD2.n99 VSUBS 0.027776f
C134 VDD2.n100 VSUBS 0.027776f
C135 VDD2.n101 VSUBS 0.014925f
C136 VDD2.n102 VSUBS 0.015364f
C137 VDD2.n103 VSUBS 0.015364f
C138 VDD2.n104 VSUBS 0.035278f
C139 VDD2.n105 VSUBS 0.035278f
C140 VDD2.n106 VSUBS 0.015803f
C141 VDD2.n107 VSUBS 0.014925f
C142 VDD2.n108 VSUBS 0.027776f
C143 VDD2.n109 VSUBS 0.027776f
C144 VDD2.n110 VSUBS 0.014925f
C145 VDD2.n111 VSUBS 0.015803f
C146 VDD2.n112 VSUBS 0.035278f
C147 VDD2.n113 VSUBS 0.087415f
C148 VDD2.n114 VSUBS 0.015803f
C149 VDD2.n115 VSUBS 0.014925f
C150 VDD2.n116 VSUBS 0.069514f
C151 VDD2.n117 VSUBS 0.063347f
C152 VDD2.n118 VSUBS 2.79301f
C153 VDD2.t9 VSUBS 0.237489f
C154 VDD2.t3 VSUBS 0.237489f
C155 VDD2.n119 VSUBS 1.82872f
C156 VDD2.n120 VSUBS 0.718124f
C157 VDD2.t1 VSUBS 0.237489f
C158 VDD2.t7 VSUBS 0.237489f
C159 VDD2.n121 VSUBS 1.84235f
C160 VN.n0 VSUBS 0.045424f
C161 VN.t7 VSUBS 1.88322f
C162 VN.n1 VSUBS 0.053896f
C163 VN.n2 VSUBS 0.034452f
C164 VN.t5 VSUBS 1.88322f
C165 VN.n3 VSUBS 0.032124f
C166 VN.n4 VSUBS 0.034452f
C167 VN.t9 VSUBS 1.88322f
C168 VN.n5 VSUBS 0.032124f
C169 VN.n6 VSUBS 0.253403f
C170 VN.t3 VSUBS 1.88322f
C171 VN.t1 VSUBS 2.03087f
C172 VN.n7 VSUBS 0.770209f
C173 VN.n8 VSUBS 0.754375f
C174 VN.n9 VSUBS 0.044777f
C175 VN.n10 VSUBS 0.063881f
C176 VN.n11 VSUBS 0.034452f
C177 VN.n12 VSUBS 0.034452f
C178 VN.n13 VSUBS 0.034452f
C179 VN.n14 VSUBS 0.069549f
C180 VN.n15 VSUBS 0.712223f
C181 VN.n16 VSUBS 0.069549f
C182 VN.n17 VSUBS 0.034452f
C183 VN.n18 VSUBS 0.034452f
C184 VN.n19 VSUBS 0.034452f
C185 VN.n20 VSUBS 0.063881f
C186 VN.n21 VSUBS 0.044777f
C187 VN.n22 VSUBS 0.679554f
C188 VN.n23 VSUBS 0.052424f
C189 VN.n24 VSUBS 0.034452f
C190 VN.n25 VSUBS 0.034452f
C191 VN.n26 VSUBS 0.034452f
C192 VN.n27 VSUBS 0.047128f
C193 VN.n28 VSUBS 0.056884f
C194 VN.n29 VSUBS 0.776048f
C195 VN.n30 VSUBS 0.042108f
C196 VN.n31 VSUBS 0.045424f
C197 VN.t4 VSUBS 1.88322f
C198 VN.n32 VSUBS 0.053896f
C199 VN.n33 VSUBS 0.034452f
C200 VN.t0 VSUBS 1.88322f
C201 VN.n34 VSUBS 0.032124f
C202 VN.n35 VSUBS 0.034452f
C203 VN.t6 VSUBS 1.88322f
C204 VN.n36 VSUBS 0.032124f
C205 VN.n37 VSUBS 0.253403f
C206 VN.t8 VSUBS 1.88322f
C207 VN.t2 VSUBS 2.03087f
C208 VN.n38 VSUBS 0.770209f
C209 VN.n39 VSUBS 0.754375f
C210 VN.n40 VSUBS 0.044777f
C211 VN.n41 VSUBS 0.063881f
C212 VN.n42 VSUBS 0.034452f
C213 VN.n43 VSUBS 0.034452f
C214 VN.n44 VSUBS 0.034452f
C215 VN.n45 VSUBS 0.069549f
C216 VN.n46 VSUBS 0.712223f
C217 VN.n47 VSUBS 0.069549f
C218 VN.n48 VSUBS 0.034452f
C219 VN.n49 VSUBS 0.034452f
C220 VN.n50 VSUBS 0.034452f
C221 VN.n51 VSUBS 0.063881f
C222 VN.n52 VSUBS 0.044777f
C223 VN.n53 VSUBS 0.679554f
C224 VN.n54 VSUBS 0.052424f
C225 VN.n55 VSUBS 0.034452f
C226 VN.n56 VSUBS 0.034452f
C227 VN.n57 VSUBS 0.034452f
C228 VN.n58 VSUBS 0.047128f
C229 VN.n59 VSUBS 0.056884f
C230 VN.n60 VSUBS 0.776048f
C231 VN.n61 VSUBS 1.81666f
C232 VDD1.n0 VSUBS 0.031238f
C233 VDD1.n1 VSUBS 0.02789f
C234 VDD1.n2 VSUBS 0.014987f
C235 VDD1.n3 VSUBS 0.035424f
C236 VDD1.n4 VSUBS 0.015869f
C237 VDD1.n5 VSUBS 0.02789f
C238 VDD1.n6 VSUBS 0.014987f
C239 VDD1.n7 VSUBS 0.035424f
C240 VDD1.n8 VSUBS 0.015869f
C241 VDD1.n9 VSUBS 0.02789f
C242 VDD1.n10 VSUBS 0.014987f
C243 VDD1.n11 VSUBS 0.035424f
C244 VDD1.n12 VSUBS 0.035424f
C245 VDD1.n13 VSUBS 0.015869f
C246 VDD1.n14 VSUBS 0.02789f
C247 VDD1.n15 VSUBS 0.014987f
C248 VDD1.n16 VSUBS 0.035424f
C249 VDD1.n17 VSUBS 0.015869f
C250 VDD1.n18 VSUBS 0.204784f
C251 VDD1.t6 VSUBS 0.076238f
C252 VDD1.n19 VSUBS 0.026568f
C253 VDD1.n20 VSUBS 0.026648f
C254 VDD1.n21 VSUBS 0.014987f
C255 VDD1.n22 VSUBS 1.22611f
C256 VDD1.n23 VSUBS 0.02789f
C257 VDD1.n24 VSUBS 0.014987f
C258 VDD1.n25 VSUBS 0.015869f
C259 VDD1.n26 VSUBS 0.035424f
C260 VDD1.n27 VSUBS 0.035424f
C261 VDD1.n28 VSUBS 0.015869f
C262 VDD1.n29 VSUBS 0.014987f
C263 VDD1.n30 VSUBS 0.02789f
C264 VDD1.n31 VSUBS 0.02789f
C265 VDD1.n32 VSUBS 0.014987f
C266 VDD1.n33 VSUBS 0.015869f
C267 VDD1.n34 VSUBS 0.035424f
C268 VDD1.n35 VSUBS 0.035424f
C269 VDD1.n36 VSUBS 0.015869f
C270 VDD1.n37 VSUBS 0.014987f
C271 VDD1.n38 VSUBS 0.02789f
C272 VDD1.n39 VSUBS 0.02789f
C273 VDD1.n40 VSUBS 0.014987f
C274 VDD1.n41 VSUBS 0.015428f
C275 VDD1.n42 VSUBS 0.015428f
C276 VDD1.n43 VSUBS 0.035424f
C277 VDD1.n44 VSUBS 0.035424f
C278 VDD1.n45 VSUBS 0.015869f
C279 VDD1.n46 VSUBS 0.014987f
C280 VDD1.n47 VSUBS 0.02789f
C281 VDD1.n48 VSUBS 0.02789f
C282 VDD1.n49 VSUBS 0.014987f
C283 VDD1.n50 VSUBS 0.015869f
C284 VDD1.n51 VSUBS 0.035424f
C285 VDD1.n52 VSUBS 0.087776f
C286 VDD1.n53 VSUBS 0.015869f
C287 VDD1.n54 VSUBS 0.014987f
C288 VDD1.n55 VSUBS 0.069801f
C289 VDD1.n56 VSUBS 0.071604f
C290 VDD1.t2 VSUBS 0.238469f
C291 VDD1.t9 VSUBS 0.238469f
C292 VDD1.n57 VSUBS 1.83626f
C293 VDD1.n58 VSUBS 0.939518f
C294 VDD1.n59 VSUBS 0.031238f
C295 VDD1.n60 VSUBS 0.02789f
C296 VDD1.n61 VSUBS 0.014987f
C297 VDD1.n62 VSUBS 0.035424f
C298 VDD1.n63 VSUBS 0.015869f
C299 VDD1.n64 VSUBS 0.02789f
C300 VDD1.n65 VSUBS 0.014987f
C301 VDD1.n66 VSUBS 0.035424f
C302 VDD1.n67 VSUBS 0.015869f
C303 VDD1.n68 VSUBS 0.02789f
C304 VDD1.n69 VSUBS 0.014987f
C305 VDD1.n70 VSUBS 0.035424f
C306 VDD1.n71 VSUBS 0.015869f
C307 VDD1.n72 VSUBS 0.02789f
C308 VDD1.n73 VSUBS 0.014987f
C309 VDD1.n74 VSUBS 0.035424f
C310 VDD1.n75 VSUBS 0.015869f
C311 VDD1.n76 VSUBS 0.204784f
C312 VDD1.t3 VSUBS 0.076238f
C313 VDD1.n77 VSUBS 0.026568f
C314 VDD1.n78 VSUBS 0.026648f
C315 VDD1.n79 VSUBS 0.014987f
C316 VDD1.n80 VSUBS 1.22611f
C317 VDD1.n81 VSUBS 0.02789f
C318 VDD1.n82 VSUBS 0.014987f
C319 VDD1.n83 VSUBS 0.015869f
C320 VDD1.n84 VSUBS 0.035424f
C321 VDD1.n85 VSUBS 0.035424f
C322 VDD1.n86 VSUBS 0.015869f
C323 VDD1.n87 VSUBS 0.014987f
C324 VDD1.n88 VSUBS 0.02789f
C325 VDD1.n89 VSUBS 0.02789f
C326 VDD1.n90 VSUBS 0.014987f
C327 VDD1.n91 VSUBS 0.015869f
C328 VDD1.n92 VSUBS 0.035424f
C329 VDD1.n93 VSUBS 0.035424f
C330 VDD1.n94 VSUBS 0.035424f
C331 VDD1.n95 VSUBS 0.015869f
C332 VDD1.n96 VSUBS 0.014987f
C333 VDD1.n97 VSUBS 0.02789f
C334 VDD1.n98 VSUBS 0.02789f
C335 VDD1.n99 VSUBS 0.014987f
C336 VDD1.n100 VSUBS 0.015428f
C337 VDD1.n101 VSUBS 0.015428f
C338 VDD1.n102 VSUBS 0.035424f
C339 VDD1.n103 VSUBS 0.035424f
C340 VDD1.n104 VSUBS 0.015869f
C341 VDD1.n105 VSUBS 0.014987f
C342 VDD1.n106 VSUBS 0.02789f
C343 VDD1.n107 VSUBS 0.02789f
C344 VDD1.n108 VSUBS 0.014987f
C345 VDD1.n109 VSUBS 0.015869f
C346 VDD1.n110 VSUBS 0.035424f
C347 VDD1.n111 VSUBS 0.087776f
C348 VDD1.n112 VSUBS 0.015869f
C349 VDD1.n113 VSUBS 0.014987f
C350 VDD1.n114 VSUBS 0.069801f
C351 VDD1.n115 VSUBS 0.071604f
C352 VDD1.t5 VSUBS 0.238469f
C353 VDD1.t8 VSUBS 0.238469f
C354 VDD1.n116 VSUBS 1.83626f
C355 VDD1.n117 VSUBS 0.930875f
C356 VDD1.t4 VSUBS 0.238469f
C357 VDD1.t7 VSUBS 0.238469f
C358 VDD1.n118 VSUBS 1.85f
C359 VDD1.n119 VSUBS 3.11683f
C360 VDD1.t1 VSUBS 0.238469f
C361 VDD1.t0 VSUBS 0.238469f
C362 VDD1.n120 VSUBS 1.83626f
C363 VDD1.n121 VSUBS 3.37082f
C364 VTAIL.t1 VSUBS 0.245919f
C365 VTAIL.t4 VSUBS 0.245919f
C366 VTAIL.n0 VSUBS 1.75512f
C367 VTAIL.n1 VSUBS 0.886578f
C368 VTAIL.n2 VSUBS 0.032214f
C369 VTAIL.n3 VSUBS 0.028762f
C370 VTAIL.n4 VSUBS 0.015455f
C371 VTAIL.n5 VSUBS 0.03653f
C372 VTAIL.n6 VSUBS 0.016364f
C373 VTAIL.n7 VSUBS 0.028762f
C374 VTAIL.n8 VSUBS 0.015455f
C375 VTAIL.n9 VSUBS 0.03653f
C376 VTAIL.n10 VSUBS 0.016364f
C377 VTAIL.n11 VSUBS 0.028762f
C378 VTAIL.n12 VSUBS 0.015455f
C379 VTAIL.n13 VSUBS 0.03653f
C380 VTAIL.n14 VSUBS 0.016364f
C381 VTAIL.n15 VSUBS 0.028762f
C382 VTAIL.n16 VSUBS 0.015455f
C383 VTAIL.n17 VSUBS 0.03653f
C384 VTAIL.n18 VSUBS 0.016364f
C385 VTAIL.n19 VSUBS 0.211181f
C386 VTAIL.t15 VSUBS 0.07862f
C387 VTAIL.n20 VSUBS 0.027398f
C388 VTAIL.n21 VSUBS 0.02748f
C389 VTAIL.n22 VSUBS 0.015455f
C390 VTAIL.n23 VSUBS 1.26441f
C391 VTAIL.n24 VSUBS 0.028762f
C392 VTAIL.n25 VSUBS 0.015455f
C393 VTAIL.n26 VSUBS 0.016364f
C394 VTAIL.n27 VSUBS 0.03653f
C395 VTAIL.n28 VSUBS 0.03653f
C396 VTAIL.n29 VSUBS 0.016364f
C397 VTAIL.n30 VSUBS 0.015455f
C398 VTAIL.n31 VSUBS 0.028762f
C399 VTAIL.n32 VSUBS 0.028762f
C400 VTAIL.n33 VSUBS 0.015455f
C401 VTAIL.n34 VSUBS 0.016364f
C402 VTAIL.n35 VSUBS 0.03653f
C403 VTAIL.n36 VSUBS 0.03653f
C404 VTAIL.n37 VSUBS 0.03653f
C405 VTAIL.n38 VSUBS 0.016364f
C406 VTAIL.n39 VSUBS 0.015455f
C407 VTAIL.n40 VSUBS 0.028762f
C408 VTAIL.n41 VSUBS 0.028762f
C409 VTAIL.n42 VSUBS 0.015455f
C410 VTAIL.n43 VSUBS 0.01591f
C411 VTAIL.n44 VSUBS 0.01591f
C412 VTAIL.n45 VSUBS 0.03653f
C413 VTAIL.n46 VSUBS 0.03653f
C414 VTAIL.n47 VSUBS 0.016364f
C415 VTAIL.n48 VSUBS 0.015455f
C416 VTAIL.n49 VSUBS 0.028762f
C417 VTAIL.n50 VSUBS 0.028762f
C418 VTAIL.n51 VSUBS 0.015455f
C419 VTAIL.n52 VSUBS 0.016364f
C420 VTAIL.n53 VSUBS 0.03653f
C421 VTAIL.n54 VSUBS 0.090518f
C422 VTAIL.n55 VSUBS 0.016364f
C423 VTAIL.n56 VSUBS 0.015455f
C424 VTAIL.n57 VSUBS 0.071982f
C425 VTAIL.n58 VSUBS 0.045776f
C426 VTAIL.n59 VSUBS 0.333666f
C427 VTAIL.t11 VSUBS 0.245919f
C428 VTAIL.t12 VSUBS 0.245919f
C429 VTAIL.n60 VSUBS 1.75512f
C430 VTAIL.n61 VSUBS 0.968868f
C431 VTAIL.t17 VSUBS 0.245919f
C432 VTAIL.t14 VSUBS 0.245919f
C433 VTAIL.n62 VSUBS 1.75512f
C434 VTAIL.n63 VSUBS 2.39897f
C435 VTAIL.t3 VSUBS 0.245919f
C436 VTAIL.t8 VSUBS 0.245919f
C437 VTAIL.n64 VSUBS 1.75513f
C438 VTAIL.n65 VSUBS 2.39896f
C439 VTAIL.t9 VSUBS 0.245919f
C440 VTAIL.t0 VSUBS 0.245919f
C441 VTAIL.n66 VSUBS 1.75513f
C442 VTAIL.n67 VSUBS 0.968857f
C443 VTAIL.n68 VSUBS 0.032214f
C444 VTAIL.n69 VSUBS 0.028762f
C445 VTAIL.n70 VSUBS 0.015455f
C446 VTAIL.n71 VSUBS 0.03653f
C447 VTAIL.n72 VSUBS 0.016364f
C448 VTAIL.n73 VSUBS 0.028762f
C449 VTAIL.n74 VSUBS 0.015455f
C450 VTAIL.n75 VSUBS 0.03653f
C451 VTAIL.n76 VSUBS 0.016364f
C452 VTAIL.n77 VSUBS 0.028762f
C453 VTAIL.n78 VSUBS 0.015455f
C454 VTAIL.n79 VSUBS 0.03653f
C455 VTAIL.n80 VSUBS 0.03653f
C456 VTAIL.n81 VSUBS 0.016364f
C457 VTAIL.n82 VSUBS 0.028762f
C458 VTAIL.n83 VSUBS 0.015455f
C459 VTAIL.n84 VSUBS 0.03653f
C460 VTAIL.n85 VSUBS 0.016364f
C461 VTAIL.n86 VSUBS 0.211181f
C462 VTAIL.t7 VSUBS 0.07862f
C463 VTAIL.n87 VSUBS 0.027398f
C464 VTAIL.n88 VSUBS 0.02748f
C465 VTAIL.n89 VSUBS 0.015455f
C466 VTAIL.n90 VSUBS 1.26441f
C467 VTAIL.n91 VSUBS 0.028762f
C468 VTAIL.n92 VSUBS 0.015455f
C469 VTAIL.n93 VSUBS 0.016364f
C470 VTAIL.n94 VSUBS 0.03653f
C471 VTAIL.n95 VSUBS 0.03653f
C472 VTAIL.n96 VSUBS 0.016364f
C473 VTAIL.n97 VSUBS 0.015455f
C474 VTAIL.n98 VSUBS 0.028762f
C475 VTAIL.n99 VSUBS 0.028762f
C476 VTAIL.n100 VSUBS 0.015455f
C477 VTAIL.n101 VSUBS 0.016364f
C478 VTAIL.n102 VSUBS 0.03653f
C479 VTAIL.n103 VSUBS 0.03653f
C480 VTAIL.n104 VSUBS 0.016364f
C481 VTAIL.n105 VSUBS 0.015455f
C482 VTAIL.n106 VSUBS 0.028762f
C483 VTAIL.n107 VSUBS 0.028762f
C484 VTAIL.n108 VSUBS 0.015455f
C485 VTAIL.n109 VSUBS 0.01591f
C486 VTAIL.n110 VSUBS 0.01591f
C487 VTAIL.n111 VSUBS 0.03653f
C488 VTAIL.n112 VSUBS 0.03653f
C489 VTAIL.n113 VSUBS 0.016364f
C490 VTAIL.n114 VSUBS 0.015455f
C491 VTAIL.n115 VSUBS 0.028762f
C492 VTAIL.n116 VSUBS 0.028762f
C493 VTAIL.n117 VSUBS 0.015455f
C494 VTAIL.n118 VSUBS 0.016364f
C495 VTAIL.n119 VSUBS 0.03653f
C496 VTAIL.n120 VSUBS 0.090518f
C497 VTAIL.n121 VSUBS 0.016364f
C498 VTAIL.n122 VSUBS 0.015455f
C499 VTAIL.n123 VSUBS 0.071982f
C500 VTAIL.n124 VSUBS 0.045776f
C501 VTAIL.n125 VSUBS 0.333666f
C502 VTAIL.t16 VSUBS 0.245919f
C503 VTAIL.t10 VSUBS 0.245919f
C504 VTAIL.n126 VSUBS 1.75513f
C505 VTAIL.n127 VSUBS 0.924916f
C506 VTAIL.t13 VSUBS 0.245919f
C507 VTAIL.t19 VSUBS 0.245919f
C508 VTAIL.n128 VSUBS 1.75513f
C509 VTAIL.n129 VSUBS 0.968857f
C510 VTAIL.n130 VSUBS 0.032214f
C511 VTAIL.n131 VSUBS 0.028762f
C512 VTAIL.n132 VSUBS 0.015455f
C513 VTAIL.n133 VSUBS 0.03653f
C514 VTAIL.n134 VSUBS 0.016364f
C515 VTAIL.n135 VSUBS 0.028762f
C516 VTAIL.n136 VSUBS 0.015455f
C517 VTAIL.n137 VSUBS 0.03653f
C518 VTAIL.n138 VSUBS 0.016364f
C519 VTAIL.n139 VSUBS 0.028762f
C520 VTAIL.n140 VSUBS 0.015455f
C521 VTAIL.n141 VSUBS 0.03653f
C522 VTAIL.n142 VSUBS 0.03653f
C523 VTAIL.n143 VSUBS 0.016364f
C524 VTAIL.n144 VSUBS 0.028762f
C525 VTAIL.n145 VSUBS 0.015455f
C526 VTAIL.n146 VSUBS 0.03653f
C527 VTAIL.n147 VSUBS 0.016364f
C528 VTAIL.n148 VSUBS 0.211181f
C529 VTAIL.t18 VSUBS 0.07862f
C530 VTAIL.n149 VSUBS 0.027398f
C531 VTAIL.n150 VSUBS 0.02748f
C532 VTAIL.n151 VSUBS 0.015455f
C533 VTAIL.n152 VSUBS 1.26441f
C534 VTAIL.n153 VSUBS 0.028762f
C535 VTAIL.n154 VSUBS 0.015455f
C536 VTAIL.n155 VSUBS 0.016364f
C537 VTAIL.n156 VSUBS 0.03653f
C538 VTAIL.n157 VSUBS 0.03653f
C539 VTAIL.n158 VSUBS 0.016364f
C540 VTAIL.n159 VSUBS 0.015455f
C541 VTAIL.n160 VSUBS 0.028762f
C542 VTAIL.n161 VSUBS 0.028762f
C543 VTAIL.n162 VSUBS 0.015455f
C544 VTAIL.n163 VSUBS 0.016364f
C545 VTAIL.n164 VSUBS 0.03653f
C546 VTAIL.n165 VSUBS 0.03653f
C547 VTAIL.n166 VSUBS 0.016364f
C548 VTAIL.n167 VSUBS 0.015455f
C549 VTAIL.n168 VSUBS 0.028762f
C550 VTAIL.n169 VSUBS 0.028762f
C551 VTAIL.n170 VSUBS 0.015455f
C552 VTAIL.n171 VSUBS 0.01591f
C553 VTAIL.n172 VSUBS 0.01591f
C554 VTAIL.n173 VSUBS 0.03653f
C555 VTAIL.n174 VSUBS 0.03653f
C556 VTAIL.n175 VSUBS 0.016364f
C557 VTAIL.n176 VSUBS 0.015455f
C558 VTAIL.n177 VSUBS 0.028762f
C559 VTAIL.n178 VSUBS 0.028762f
C560 VTAIL.n179 VSUBS 0.015455f
C561 VTAIL.n180 VSUBS 0.016364f
C562 VTAIL.n181 VSUBS 0.03653f
C563 VTAIL.n182 VSUBS 0.090518f
C564 VTAIL.n183 VSUBS 0.016364f
C565 VTAIL.n184 VSUBS 0.015455f
C566 VTAIL.n185 VSUBS 0.071982f
C567 VTAIL.n186 VSUBS 0.045776f
C568 VTAIL.n187 VSUBS 1.63274f
C569 VTAIL.n188 VSUBS 0.032214f
C570 VTAIL.n189 VSUBS 0.028762f
C571 VTAIL.n190 VSUBS 0.015455f
C572 VTAIL.n191 VSUBS 0.03653f
C573 VTAIL.n192 VSUBS 0.016364f
C574 VTAIL.n193 VSUBS 0.028762f
C575 VTAIL.n194 VSUBS 0.015455f
C576 VTAIL.n195 VSUBS 0.03653f
C577 VTAIL.n196 VSUBS 0.016364f
C578 VTAIL.n197 VSUBS 0.028762f
C579 VTAIL.n198 VSUBS 0.015455f
C580 VTAIL.n199 VSUBS 0.03653f
C581 VTAIL.n200 VSUBS 0.016364f
C582 VTAIL.n201 VSUBS 0.028762f
C583 VTAIL.n202 VSUBS 0.015455f
C584 VTAIL.n203 VSUBS 0.03653f
C585 VTAIL.n204 VSUBS 0.016364f
C586 VTAIL.n205 VSUBS 0.211181f
C587 VTAIL.t5 VSUBS 0.07862f
C588 VTAIL.n206 VSUBS 0.027398f
C589 VTAIL.n207 VSUBS 0.02748f
C590 VTAIL.n208 VSUBS 0.015455f
C591 VTAIL.n209 VSUBS 1.26441f
C592 VTAIL.n210 VSUBS 0.028762f
C593 VTAIL.n211 VSUBS 0.015455f
C594 VTAIL.n212 VSUBS 0.016364f
C595 VTAIL.n213 VSUBS 0.03653f
C596 VTAIL.n214 VSUBS 0.03653f
C597 VTAIL.n215 VSUBS 0.016364f
C598 VTAIL.n216 VSUBS 0.015455f
C599 VTAIL.n217 VSUBS 0.028762f
C600 VTAIL.n218 VSUBS 0.028762f
C601 VTAIL.n219 VSUBS 0.015455f
C602 VTAIL.n220 VSUBS 0.016364f
C603 VTAIL.n221 VSUBS 0.03653f
C604 VTAIL.n222 VSUBS 0.03653f
C605 VTAIL.n223 VSUBS 0.03653f
C606 VTAIL.n224 VSUBS 0.016364f
C607 VTAIL.n225 VSUBS 0.015455f
C608 VTAIL.n226 VSUBS 0.028762f
C609 VTAIL.n227 VSUBS 0.028762f
C610 VTAIL.n228 VSUBS 0.015455f
C611 VTAIL.n229 VSUBS 0.01591f
C612 VTAIL.n230 VSUBS 0.01591f
C613 VTAIL.n231 VSUBS 0.03653f
C614 VTAIL.n232 VSUBS 0.03653f
C615 VTAIL.n233 VSUBS 0.016364f
C616 VTAIL.n234 VSUBS 0.015455f
C617 VTAIL.n235 VSUBS 0.028762f
C618 VTAIL.n236 VSUBS 0.028762f
C619 VTAIL.n237 VSUBS 0.015455f
C620 VTAIL.n238 VSUBS 0.016364f
C621 VTAIL.n239 VSUBS 0.03653f
C622 VTAIL.n240 VSUBS 0.090518f
C623 VTAIL.n241 VSUBS 0.016364f
C624 VTAIL.n242 VSUBS 0.015455f
C625 VTAIL.n243 VSUBS 0.071982f
C626 VTAIL.n244 VSUBS 0.045776f
C627 VTAIL.n245 VSUBS 1.63274f
C628 VTAIL.t2 VSUBS 0.245919f
C629 VTAIL.t6 VSUBS 0.245919f
C630 VTAIL.n246 VSUBS 1.75512f
C631 VTAIL.n247 VSUBS 0.832251f
C632 VP.n0 VSUBS 0.0466f
C633 VP.t2 VSUBS 1.932f
C634 VP.n1 VSUBS 0.055292f
C635 VP.n2 VSUBS 0.035344f
C636 VP.t5 VSUBS 1.932f
C637 VP.n3 VSUBS 0.032957f
C638 VP.n4 VSUBS 0.035344f
C639 VP.t1 VSUBS 1.932f
C640 VP.n5 VSUBS 0.032957f
C641 VP.n6 VSUBS 0.035344f
C642 VP.t4 VSUBS 1.932f
C643 VP.n7 VSUBS 0.055292f
C644 VP.n8 VSUBS 0.0466f
C645 VP.t6 VSUBS 1.932f
C646 VP.n9 VSUBS 0.0466f
C647 VP.t9 VSUBS 1.932f
C648 VP.n10 VSUBS 0.055292f
C649 VP.n11 VSUBS 0.035344f
C650 VP.t8 VSUBS 1.932f
C651 VP.n12 VSUBS 0.032957f
C652 VP.n13 VSUBS 0.035344f
C653 VP.t0 VSUBS 1.932f
C654 VP.n14 VSUBS 0.032957f
C655 VP.n15 VSUBS 0.259967f
C656 VP.t7 VSUBS 1.932f
C657 VP.t3 VSUBS 2.08348f
C658 VP.n16 VSUBS 0.790161f
C659 VP.n17 VSUBS 0.773917f
C660 VP.n18 VSUBS 0.045937f
C661 VP.n19 VSUBS 0.065536f
C662 VP.n20 VSUBS 0.035344f
C663 VP.n21 VSUBS 0.035344f
C664 VP.n22 VSUBS 0.035344f
C665 VP.n23 VSUBS 0.071351f
C666 VP.n24 VSUBS 0.730673f
C667 VP.n25 VSUBS 0.071351f
C668 VP.n26 VSUBS 0.035344f
C669 VP.n27 VSUBS 0.035344f
C670 VP.n28 VSUBS 0.035344f
C671 VP.n29 VSUBS 0.065536f
C672 VP.n30 VSUBS 0.045937f
C673 VP.n31 VSUBS 0.697157f
C674 VP.n32 VSUBS 0.053782f
C675 VP.n33 VSUBS 0.035344f
C676 VP.n34 VSUBS 0.035344f
C677 VP.n35 VSUBS 0.035344f
C678 VP.n36 VSUBS 0.048349f
C679 VP.n37 VSUBS 0.058358f
C680 VP.n38 VSUBS 0.796151f
C681 VP.n39 VSUBS 1.84461f
C682 VP.n40 VSUBS 1.87091f
C683 VP.n41 VSUBS 0.796151f
C684 VP.n42 VSUBS 0.058358f
C685 VP.n43 VSUBS 0.048349f
C686 VP.n44 VSUBS 0.035344f
C687 VP.n45 VSUBS 0.035344f
C688 VP.n46 VSUBS 0.035344f
C689 VP.n47 VSUBS 0.053782f
C690 VP.n48 VSUBS 0.697157f
C691 VP.n49 VSUBS 0.045937f
C692 VP.n50 VSUBS 0.065536f
C693 VP.n51 VSUBS 0.035344f
C694 VP.n52 VSUBS 0.035344f
C695 VP.n53 VSUBS 0.035344f
C696 VP.n54 VSUBS 0.071351f
C697 VP.n55 VSUBS 0.730673f
C698 VP.n56 VSUBS 0.071351f
C699 VP.n57 VSUBS 0.035344f
C700 VP.n58 VSUBS 0.035344f
C701 VP.n59 VSUBS 0.035344f
C702 VP.n60 VSUBS 0.065536f
C703 VP.n61 VSUBS 0.045937f
C704 VP.n62 VSUBS 0.697157f
C705 VP.n63 VSUBS 0.053782f
C706 VP.n64 VSUBS 0.035344f
C707 VP.n65 VSUBS 0.035344f
C708 VP.n66 VSUBS 0.035344f
C709 VP.n67 VSUBS 0.048349f
C710 VP.n68 VSUBS 0.058358f
C711 VP.n69 VSUBS 0.796151f
C712 VP.n70 VSUBS 0.043198f
C713 B.n0 VSUBS 0.008026f
C714 B.n1 VSUBS 0.008026f
C715 B.n2 VSUBS 0.01187f
C716 B.n3 VSUBS 0.009097f
C717 B.n4 VSUBS 0.009097f
C718 B.n5 VSUBS 0.009097f
C719 B.n6 VSUBS 0.009097f
C720 B.n7 VSUBS 0.009097f
C721 B.n8 VSUBS 0.009097f
C722 B.n9 VSUBS 0.009097f
C723 B.n10 VSUBS 0.009097f
C724 B.n11 VSUBS 0.009097f
C725 B.n12 VSUBS 0.009097f
C726 B.n13 VSUBS 0.009097f
C727 B.n14 VSUBS 0.009097f
C728 B.n15 VSUBS 0.009097f
C729 B.n16 VSUBS 0.009097f
C730 B.n17 VSUBS 0.009097f
C731 B.n18 VSUBS 0.009097f
C732 B.n19 VSUBS 0.009097f
C733 B.n20 VSUBS 0.009097f
C734 B.n21 VSUBS 0.009097f
C735 B.n22 VSUBS 0.009097f
C736 B.n23 VSUBS 0.009097f
C737 B.n24 VSUBS 0.009097f
C738 B.n25 VSUBS 0.022829f
C739 B.n26 VSUBS 0.009097f
C740 B.n27 VSUBS 0.009097f
C741 B.n28 VSUBS 0.009097f
C742 B.n29 VSUBS 0.009097f
C743 B.n30 VSUBS 0.009097f
C744 B.n31 VSUBS 0.009097f
C745 B.n32 VSUBS 0.009097f
C746 B.n33 VSUBS 0.009097f
C747 B.n34 VSUBS 0.009097f
C748 B.n35 VSUBS 0.009097f
C749 B.n36 VSUBS 0.009097f
C750 B.n37 VSUBS 0.009097f
C751 B.n38 VSUBS 0.009097f
C752 B.n39 VSUBS 0.009097f
C753 B.n40 VSUBS 0.009097f
C754 B.n41 VSUBS 0.009097f
C755 B.n42 VSUBS 0.009097f
C756 B.n43 VSUBS 0.009097f
C757 B.t1 VSUBS 0.240773f
C758 B.t2 VSUBS 0.271618f
C759 B.t0 VSUBS 1.17107f
C760 B.n44 VSUBS 0.430357f
C761 B.n45 VSUBS 0.301291f
C762 B.n46 VSUBS 0.021076f
C763 B.n47 VSUBS 0.009097f
C764 B.n48 VSUBS 0.009097f
C765 B.n49 VSUBS 0.009097f
C766 B.n50 VSUBS 0.009097f
C767 B.n51 VSUBS 0.009097f
C768 B.t10 VSUBS 0.240777f
C769 B.t11 VSUBS 0.271621f
C770 B.t9 VSUBS 1.17107f
C771 B.n52 VSUBS 0.430354f
C772 B.n53 VSUBS 0.301287f
C773 B.n54 VSUBS 0.009097f
C774 B.n55 VSUBS 0.009097f
C775 B.n56 VSUBS 0.009097f
C776 B.n57 VSUBS 0.009097f
C777 B.n58 VSUBS 0.009097f
C778 B.n59 VSUBS 0.009097f
C779 B.n60 VSUBS 0.009097f
C780 B.n61 VSUBS 0.009097f
C781 B.n62 VSUBS 0.009097f
C782 B.n63 VSUBS 0.009097f
C783 B.n64 VSUBS 0.009097f
C784 B.n65 VSUBS 0.009097f
C785 B.n66 VSUBS 0.009097f
C786 B.n67 VSUBS 0.009097f
C787 B.n68 VSUBS 0.009097f
C788 B.n69 VSUBS 0.009097f
C789 B.n70 VSUBS 0.009097f
C790 B.n71 VSUBS 0.009097f
C791 B.n72 VSUBS 0.022829f
C792 B.n73 VSUBS 0.009097f
C793 B.n74 VSUBS 0.009097f
C794 B.n75 VSUBS 0.009097f
C795 B.n76 VSUBS 0.009097f
C796 B.n77 VSUBS 0.009097f
C797 B.n78 VSUBS 0.009097f
C798 B.n79 VSUBS 0.009097f
C799 B.n80 VSUBS 0.009097f
C800 B.n81 VSUBS 0.009097f
C801 B.n82 VSUBS 0.009097f
C802 B.n83 VSUBS 0.009097f
C803 B.n84 VSUBS 0.009097f
C804 B.n85 VSUBS 0.009097f
C805 B.n86 VSUBS 0.009097f
C806 B.n87 VSUBS 0.009097f
C807 B.n88 VSUBS 0.009097f
C808 B.n89 VSUBS 0.009097f
C809 B.n90 VSUBS 0.009097f
C810 B.n91 VSUBS 0.009097f
C811 B.n92 VSUBS 0.009097f
C812 B.n93 VSUBS 0.009097f
C813 B.n94 VSUBS 0.009097f
C814 B.n95 VSUBS 0.009097f
C815 B.n96 VSUBS 0.009097f
C816 B.n97 VSUBS 0.009097f
C817 B.n98 VSUBS 0.009097f
C818 B.n99 VSUBS 0.009097f
C819 B.n100 VSUBS 0.009097f
C820 B.n101 VSUBS 0.009097f
C821 B.n102 VSUBS 0.009097f
C822 B.n103 VSUBS 0.009097f
C823 B.n104 VSUBS 0.009097f
C824 B.n105 VSUBS 0.009097f
C825 B.n106 VSUBS 0.009097f
C826 B.n107 VSUBS 0.009097f
C827 B.n108 VSUBS 0.009097f
C828 B.n109 VSUBS 0.009097f
C829 B.n110 VSUBS 0.009097f
C830 B.n111 VSUBS 0.009097f
C831 B.n112 VSUBS 0.009097f
C832 B.n113 VSUBS 0.009097f
C833 B.n114 VSUBS 0.009097f
C834 B.n115 VSUBS 0.009097f
C835 B.n116 VSUBS 0.009097f
C836 B.n117 VSUBS 0.009097f
C837 B.n118 VSUBS 0.009097f
C838 B.n119 VSUBS 0.021316f
C839 B.n120 VSUBS 0.009097f
C840 B.n121 VSUBS 0.009097f
C841 B.n122 VSUBS 0.009097f
C842 B.n123 VSUBS 0.009097f
C843 B.n124 VSUBS 0.009097f
C844 B.n125 VSUBS 0.009097f
C845 B.n126 VSUBS 0.009097f
C846 B.n127 VSUBS 0.009097f
C847 B.n128 VSUBS 0.009097f
C848 B.n129 VSUBS 0.009097f
C849 B.n130 VSUBS 0.009097f
C850 B.n131 VSUBS 0.009097f
C851 B.n132 VSUBS 0.009097f
C852 B.n133 VSUBS 0.009097f
C853 B.n134 VSUBS 0.009097f
C854 B.n135 VSUBS 0.009097f
C855 B.n136 VSUBS 0.009097f
C856 B.n137 VSUBS 0.009097f
C857 B.n138 VSUBS 0.008561f
C858 B.n139 VSUBS 0.009097f
C859 B.n140 VSUBS 0.009097f
C860 B.n141 VSUBS 0.009097f
C861 B.n142 VSUBS 0.009097f
C862 B.n143 VSUBS 0.009097f
C863 B.t8 VSUBS 0.240773f
C864 B.t7 VSUBS 0.271618f
C865 B.t6 VSUBS 1.17107f
C866 B.n144 VSUBS 0.430357f
C867 B.n145 VSUBS 0.301291f
C868 B.n146 VSUBS 0.009097f
C869 B.n147 VSUBS 0.009097f
C870 B.n148 VSUBS 0.009097f
C871 B.n149 VSUBS 0.009097f
C872 B.n150 VSUBS 0.009097f
C873 B.n151 VSUBS 0.009097f
C874 B.n152 VSUBS 0.009097f
C875 B.n153 VSUBS 0.009097f
C876 B.n154 VSUBS 0.009097f
C877 B.n155 VSUBS 0.009097f
C878 B.n156 VSUBS 0.009097f
C879 B.n157 VSUBS 0.009097f
C880 B.n158 VSUBS 0.009097f
C881 B.n159 VSUBS 0.009097f
C882 B.n160 VSUBS 0.009097f
C883 B.n161 VSUBS 0.009097f
C884 B.n162 VSUBS 0.009097f
C885 B.n163 VSUBS 0.009097f
C886 B.n164 VSUBS 0.022829f
C887 B.n165 VSUBS 0.009097f
C888 B.n166 VSUBS 0.009097f
C889 B.n167 VSUBS 0.009097f
C890 B.n168 VSUBS 0.009097f
C891 B.n169 VSUBS 0.009097f
C892 B.n170 VSUBS 0.009097f
C893 B.n171 VSUBS 0.009097f
C894 B.n172 VSUBS 0.009097f
C895 B.n173 VSUBS 0.009097f
C896 B.n174 VSUBS 0.009097f
C897 B.n175 VSUBS 0.009097f
C898 B.n176 VSUBS 0.009097f
C899 B.n177 VSUBS 0.009097f
C900 B.n178 VSUBS 0.009097f
C901 B.n179 VSUBS 0.009097f
C902 B.n180 VSUBS 0.009097f
C903 B.n181 VSUBS 0.009097f
C904 B.n182 VSUBS 0.009097f
C905 B.n183 VSUBS 0.009097f
C906 B.n184 VSUBS 0.009097f
C907 B.n185 VSUBS 0.009097f
C908 B.n186 VSUBS 0.009097f
C909 B.n187 VSUBS 0.009097f
C910 B.n188 VSUBS 0.009097f
C911 B.n189 VSUBS 0.009097f
C912 B.n190 VSUBS 0.009097f
C913 B.n191 VSUBS 0.009097f
C914 B.n192 VSUBS 0.009097f
C915 B.n193 VSUBS 0.009097f
C916 B.n194 VSUBS 0.009097f
C917 B.n195 VSUBS 0.009097f
C918 B.n196 VSUBS 0.009097f
C919 B.n197 VSUBS 0.009097f
C920 B.n198 VSUBS 0.009097f
C921 B.n199 VSUBS 0.009097f
C922 B.n200 VSUBS 0.009097f
C923 B.n201 VSUBS 0.009097f
C924 B.n202 VSUBS 0.009097f
C925 B.n203 VSUBS 0.009097f
C926 B.n204 VSUBS 0.009097f
C927 B.n205 VSUBS 0.009097f
C928 B.n206 VSUBS 0.009097f
C929 B.n207 VSUBS 0.009097f
C930 B.n208 VSUBS 0.009097f
C931 B.n209 VSUBS 0.009097f
C932 B.n210 VSUBS 0.009097f
C933 B.n211 VSUBS 0.009097f
C934 B.n212 VSUBS 0.009097f
C935 B.n213 VSUBS 0.009097f
C936 B.n214 VSUBS 0.009097f
C937 B.n215 VSUBS 0.009097f
C938 B.n216 VSUBS 0.009097f
C939 B.n217 VSUBS 0.009097f
C940 B.n218 VSUBS 0.009097f
C941 B.n219 VSUBS 0.009097f
C942 B.n220 VSUBS 0.009097f
C943 B.n221 VSUBS 0.009097f
C944 B.n222 VSUBS 0.009097f
C945 B.n223 VSUBS 0.009097f
C946 B.n224 VSUBS 0.009097f
C947 B.n225 VSUBS 0.009097f
C948 B.n226 VSUBS 0.009097f
C949 B.n227 VSUBS 0.009097f
C950 B.n228 VSUBS 0.009097f
C951 B.n229 VSUBS 0.009097f
C952 B.n230 VSUBS 0.009097f
C953 B.n231 VSUBS 0.009097f
C954 B.n232 VSUBS 0.009097f
C955 B.n233 VSUBS 0.009097f
C956 B.n234 VSUBS 0.009097f
C957 B.n235 VSUBS 0.009097f
C958 B.n236 VSUBS 0.009097f
C959 B.n237 VSUBS 0.009097f
C960 B.n238 VSUBS 0.009097f
C961 B.n239 VSUBS 0.009097f
C962 B.n240 VSUBS 0.009097f
C963 B.n241 VSUBS 0.009097f
C964 B.n242 VSUBS 0.009097f
C965 B.n243 VSUBS 0.009097f
C966 B.n244 VSUBS 0.009097f
C967 B.n245 VSUBS 0.009097f
C968 B.n246 VSUBS 0.009097f
C969 B.n247 VSUBS 0.009097f
C970 B.n248 VSUBS 0.009097f
C971 B.n249 VSUBS 0.009097f
C972 B.n250 VSUBS 0.009097f
C973 B.n251 VSUBS 0.009097f
C974 B.n252 VSUBS 0.009097f
C975 B.n253 VSUBS 0.021316f
C976 B.n254 VSUBS 0.021316f
C977 B.n255 VSUBS 0.022829f
C978 B.n256 VSUBS 0.009097f
C979 B.n257 VSUBS 0.009097f
C980 B.n258 VSUBS 0.009097f
C981 B.n259 VSUBS 0.009097f
C982 B.n260 VSUBS 0.009097f
C983 B.n261 VSUBS 0.009097f
C984 B.n262 VSUBS 0.009097f
C985 B.n263 VSUBS 0.009097f
C986 B.n264 VSUBS 0.009097f
C987 B.n265 VSUBS 0.009097f
C988 B.n266 VSUBS 0.009097f
C989 B.n267 VSUBS 0.009097f
C990 B.n268 VSUBS 0.009097f
C991 B.n269 VSUBS 0.009097f
C992 B.n270 VSUBS 0.009097f
C993 B.n271 VSUBS 0.009097f
C994 B.n272 VSUBS 0.009097f
C995 B.n273 VSUBS 0.009097f
C996 B.n274 VSUBS 0.009097f
C997 B.n275 VSUBS 0.009097f
C998 B.n276 VSUBS 0.009097f
C999 B.n277 VSUBS 0.009097f
C1000 B.n278 VSUBS 0.009097f
C1001 B.n279 VSUBS 0.009097f
C1002 B.n280 VSUBS 0.009097f
C1003 B.n281 VSUBS 0.009097f
C1004 B.n282 VSUBS 0.009097f
C1005 B.n283 VSUBS 0.009097f
C1006 B.n284 VSUBS 0.009097f
C1007 B.n285 VSUBS 0.009097f
C1008 B.n286 VSUBS 0.009097f
C1009 B.n287 VSUBS 0.009097f
C1010 B.n288 VSUBS 0.009097f
C1011 B.n289 VSUBS 0.009097f
C1012 B.n290 VSUBS 0.009097f
C1013 B.n291 VSUBS 0.009097f
C1014 B.n292 VSUBS 0.009097f
C1015 B.n293 VSUBS 0.009097f
C1016 B.n294 VSUBS 0.009097f
C1017 B.n295 VSUBS 0.009097f
C1018 B.n296 VSUBS 0.009097f
C1019 B.n297 VSUBS 0.009097f
C1020 B.n298 VSUBS 0.009097f
C1021 B.n299 VSUBS 0.009097f
C1022 B.n300 VSUBS 0.009097f
C1023 B.n301 VSUBS 0.009097f
C1024 B.n302 VSUBS 0.009097f
C1025 B.n303 VSUBS 0.009097f
C1026 B.n304 VSUBS 0.009097f
C1027 B.n305 VSUBS 0.009097f
C1028 B.n306 VSUBS 0.009097f
C1029 B.n307 VSUBS 0.009097f
C1030 B.n308 VSUBS 0.009097f
C1031 B.n309 VSUBS 0.009097f
C1032 B.n310 VSUBS 0.009097f
C1033 B.n311 VSUBS 0.008561f
C1034 B.n312 VSUBS 0.021076f
C1035 B.n313 VSUBS 0.005083f
C1036 B.n314 VSUBS 0.009097f
C1037 B.n315 VSUBS 0.009097f
C1038 B.n316 VSUBS 0.009097f
C1039 B.n317 VSUBS 0.009097f
C1040 B.n318 VSUBS 0.009097f
C1041 B.n319 VSUBS 0.009097f
C1042 B.n320 VSUBS 0.009097f
C1043 B.n321 VSUBS 0.009097f
C1044 B.n322 VSUBS 0.009097f
C1045 B.n323 VSUBS 0.009097f
C1046 B.n324 VSUBS 0.009097f
C1047 B.n325 VSUBS 0.009097f
C1048 B.t5 VSUBS 0.240777f
C1049 B.t4 VSUBS 0.271621f
C1050 B.t3 VSUBS 1.17107f
C1051 B.n326 VSUBS 0.430354f
C1052 B.n327 VSUBS 0.301287f
C1053 B.n328 VSUBS 0.021076f
C1054 B.n329 VSUBS 0.005083f
C1055 B.n330 VSUBS 0.009097f
C1056 B.n331 VSUBS 0.009097f
C1057 B.n332 VSUBS 0.009097f
C1058 B.n333 VSUBS 0.009097f
C1059 B.n334 VSUBS 0.009097f
C1060 B.n335 VSUBS 0.009097f
C1061 B.n336 VSUBS 0.009097f
C1062 B.n337 VSUBS 0.009097f
C1063 B.n338 VSUBS 0.009097f
C1064 B.n339 VSUBS 0.009097f
C1065 B.n340 VSUBS 0.009097f
C1066 B.n341 VSUBS 0.009097f
C1067 B.n342 VSUBS 0.009097f
C1068 B.n343 VSUBS 0.009097f
C1069 B.n344 VSUBS 0.009097f
C1070 B.n345 VSUBS 0.009097f
C1071 B.n346 VSUBS 0.009097f
C1072 B.n347 VSUBS 0.009097f
C1073 B.n348 VSUBS 0.009097f
C1074 B.n349 VSUBS 0.009097f
C1075 B.n350 VSUBS 0.009097f
C1076 B.n351 VSUBS 0.009097f
C1077 B.n352 VSUBS 0.009097f
C1078 B.n353 VSUBS 0.009097f
C1079 B.n354 VSUBS 0.009097f
C1080 B.n355 VSUBS 0.009097f
C1081 B.n356 VSUBS 0.009097f
C1082 B.n357 VSUBS 0.009097f
C1083 B.n358 VSUBS 0.009097f
C1084 B.n359 VSUBS 0.009097f
C1085 B.n360 VSUBS 0.009097f
C1086 B.n361 VSUBS 0.009097f
C1087 B.n362 VSUBS 0.009097f
C1088 B.n363 VSUBS 0.009097f
C1089 B.n364 VSUBS 0.009097f
C1090 B.n365 VSUBS 0.009097f
C1091 B.n366 VSUBS 0.009097f
C1092 B.n367 VSUBS 0.009097f
C1093 B.n368 VSUBS 0.009097f
C1094 B.n369 VSUBS 0.009097f
C1095 B.n370 VSUBS 0.009097f
C1096 B.n371 VSUBS 0.009097f
C1097 B.n372 VSUBS 0.009097f
C1098 B.n373 VSUBS 0.009097f
C1099 B.n374 VSUBS 0.009097f
C1100 B.n375 VSUBS 0.009097f
C1101 B.n376 VSUBS 0.009097f
C1102 B.n377 VSUBS 0.009097f
C1103 B.n378 VSUBS 0.009097f
C1104 B.n379 VSUBS 0.009097f
C1105 B.n380 VSUBS 0.009097f
C1106 B.n381 VSUBS 0.009097f
C1107 B.n382 VSUBS 0.009097f
C1108 B.n383 VSUBS 0.009097f
C1109 B.n384 VSUBS 0.009097f
C1110 B.n385 VSUBS 0.009097f
C1111 B.n386 VSUBS 0.022829f
C1112 B.n387 VSUBS 0.021812f
C1113 B.n388 VSUBS 0.022333f
C1114 B.n389 VSUBS 0.009097f
C1115 B.n390 VSUBS 0.009097f
C1116 B.n391 VSUBS 0.009097f
C1117 B.n392 VSUBS 0.009097f
C1118 B.n393 VSUBS 0.009097f
C1119 B.n394 VSUBS 0.009097f
C1120 B.n395 VSUBS 0.009097f
C1121 B.n396 VSUBS 0.009097f
C1122 B.n397 VSUBS 0.009097f
C1123 B.n398 VSUBS 0.009097f
C1124 B.n399 VSUBS 0.009097f
C1125 B.n400 VSUBS 0.009097f
C1126 B.n401 VSUBS 0.009097f
C1127 B.n402 VSUBS 0.009097f
C1128 B.n403 VSUBS 0.009097f
C1129 B.n404 VSUBS 0.009097f
C1130 B.n405 VSUBS 0.009097f
C1131 B.n406 VSUBS 0.009097f
C1132 B.n407 VSUBS 0.009097f
C1133 B.n408 VSUBS 0.009097f
C1134 B.n409 VSUBS 0.009097f
C1135 B.n410 VSUBS 0.009097f
C1136 B.n411 VSUBS 0.009097f
C1137 B.n412 VSUBS 0.009097f
C1138 B.n413 VSUBS 0.009097f
C1139 B.n414 VSUBS 0.009097f
C1140 B.n415 VSUBS 0.009097f
C1141 B.n416 VSUBS 0.009097f
C1142 B.n417 VSUBS 0.009097f
C1143 B.n418 VSUBS 0.009097f
C1144 B.n419 VSUBS 0.009097f
C1145 B.n420 VSUBS 0.009097f
C1146 B.n421 VSUBS 0.009097f
C1147 B.n422 VSUBS 0.009097f
C1148 B.n423 VSUBS 0.009097f
C1149 B.n424 VSUBS 0.009097f
C1150 B.n425 VSUBS 0.009097f
C1151 B.n426 VSUBS 0.009097f
C1152 B.n427 VSUBS 0.009097f
C1153 B.n428 VSUBS 0.009097f
C1154 B.n429 VSUBS 0.009097f
C1155 B.n430 VSUBS 0.009097f
C1156 B.n431 VSUBS 0.009097f
C1157 B.n432 VSUBS 0.009097f
C1158 B.n433 VSUBS 0.009097f
C1159 B.n434 VSUBS 0.009097f
C1160 B.n435 VSUBS 0.009097f
C1161 B.n436 VSUBS 0.009097f
C1162 B.n437 VSUBS 0.009097f
C1163 B.n438 VSUBS 0.009097f
C1164 B.n439 VSUBS 0.009097f
C1165 B.n440 VSUBS 0.009097f
C1166 B.n441 VSUBS 0.009097f
C1167 B.n442 VSUBS 0.009097f
C1168 B.n443 VSUBS 0.009097f
C1169 B.n444 VSUBS 0.009097f
C1170 B.n445 VSUBS 0.009097f
C1171 B.n446 VSUBS 0.009097f
C1172 B.n447 VSUBS 0.009097f
C1173 B.n448 VSUBS 0.009097f
C1174 B.n449 VSUBS 0.009097f
C1175 B.n450 VSUBS 0.009097f
C1176 B.n451 VSUBS 0.009097f
C1177 B.n452 VSUBS 0.009097f
C1178 B.n453 VSUBS 0.009097f
C1179 B.n454 VSUBS 0.009097f
C1180 B.n455 VSUBS 0.009097f
C1181 B.n456 VSUBS 0.009097f
C1182 B.n457 VSUBS 0.009097f
C1183 B.n458 VSUBS 0.009097f
C1184 B.n459 VSUBS 0.009097f
C1185 B.n460 VSUBS 0.009097f
C1186 B.n461 VSUBS 0.009097f
C1187 B.n462 VSUBS 0.009097f
C1188 B.n463 VSUBS 0.009097f
C1189 B.n464 VSUBS 0.009097f
C1190 B.n465 VSUBS 0.009097f
C1191 B.n466 VSUBS 0.009097f
C1192 B.n467 VSUBS 0.009097f
C1193 B.n468 VSUBS 0.009097f
C1194 B.n469 VSUBS 0.009097f
C1195 B.n470 VSUBS 0.009097f
C1196 B.n471 VSUBS 0.009097f
C1197 B.n472 VSUBS 0.009097f
C1198 B.n473 VSUBS 0.009097f
C1199 B.n474 VSUBS 0.009097f
C1200 B.n475 VSUBS 0.009097f
C1201 B.n476 VSUBS 0.009097f
C1202 B.n477 VSUBS 0.009097f
C1203 B.n478 VSUBS 0.009097f
C1204 B.n479 VSUBS 0.009097f
C1205 B.n480 VSUBS 0.009097f
C1206 B.n481 VSUBS 0.009097f
C1207 B.n482 VSUBS 0.009097f
C1208 B.n483 VSUBS 0.009097f
C1209 B.n484 VSUBS 0.009097f
C1210 B.n485 VSUBS 0.009097f
C1211 B.n486 VSUBS 0.009097f
C1212 B.n487 VSUBS 0.009097f
C1213 B.n488 VSUBS 0.009097f
C1214 B.n489 VSUBS 0.009097f
C1215 B.n490 VSUBS 0.009097f
C1216 B.n491 VSUBS 0.009097f
C1217 B.n492 VSUBS 0.009097f
C1218 B.n493 VSUBS 0.009097f
C1219 B.n494 VSUBS 0.009097f
C1220 B.n495 VSUBS 0.009097f
C1221 B.n496 VSUBS 0.009097f
C1222 B.n497 VSUBS 0.009097f
C1223 B.n498 VSUBS 0.009097f
C1224 B.n499 VSUBS 0.009097f
C1225 B.n500 VSUBS 0.009097f
C1226 B.n501 VSUBS 0.009097f
C1227 B.n502 VSUBS 0.009097f
C1228 B.n503 VSUBS 0.009097f
C1229 B.n504 VSUBS 0.009097f
C1230 B.n505 VSUBS 0.009097f
C1231 B.n506 VSUBS 0.009097f
C1232 B.n507 VSUBS 0.009097f
C1233 B.n508 VSUBS 0.009097f
C1234 B.n509 VSUBS 0.009097f
C1235 B.n510 VSUBS 0.009097f
C1236 B.n511 VSUBS 0.009097f
C1237 B.n512 VSUBS 0.009097f
C1238 B.n513 VSUBS 0.009097f
C1239 B.n514 VSUBS 0.009097f
C1240 B.n515 VSUBS 0.009097f
C1241 B.n516 VSUBS 0.009097f
C1242 B.n517 VSUBS 0.009097f
C1243 B.n518 VSUBS 0.009097f
C1244 B.n519 VSUBS 0.009097f
C1245 B.n520 VSUBS 0.009097f
C1246 B.n521 VSUBS 0.009097f
C1247 B.n522 VSUBS 0.009097f
C1248 B.n523 VSUBS 0.009097f
C1249 B.n524 VSUBS 0.009097f
C1250 B.n525 VSUBS 0.009097f
C1251 B.n526 VSUBS 0.009097f
C1252 B.n527 VSUBS 0.021316f
C1253 B.n528 VSUBS 0.021316f
C1254 B.n529 VSUBS 0.022829f
C1255 B.n530 VSUBS 0.009097f
C1256 B.n531 VSUBS 0.009097f
C1257 B.n532 VSUBS 0.009097f
C1258 B.n533 VSUBS 0.009097f
C1259 B.n534 VSUBS 0.009097f
C1260 B.n535 VSUBS 0.009097f
C1261 B.n536 VSUBS 0.009097f
C1262 B.n537 VSUBS 0.009097f
C1263 B.n538 VSUBS 0.009097f
C1264 B.n539 VSUBS 0.009097f
C1265 B.n540 VSUBS 0.009097f
C1266 B.n541 VSUBS 0.009097f
C1267 B.n542 VSUBS 0.009097f
C1268 B.n543 VSUBS 0.009097f
C1269 B.n544 VSUBS 0.009097f
C1270 B.n545 VSUBS 0.009097f
C1271 B.n546 VSUBS 0.009097f
C1272 B.n547 VSUBS 0.009097f
C1273 B.n548 VSUBS 0.009097f
C1274 B.n549 VSUBS 0.009097f
C1275 B.n550 VSUBS 0.009097f
C1276 B.n551 VSUBS 0.009097f
C1277 B.n552 VSUBS 0.009097f
C1278 B.n553 VSUBS 0.009097f
C1279 B.n554 VSUBS 0.009097f
C1280 B.n555 VSUBS 0.009097f
C1281 B.n556 VSUBS 0.009097f
C1282 B.n557 VSUBS 0.009097f
C1283 B.n558 VSUBS 0.009097f
C1284 B.n559 VSUBS 0.009097f
C1285 B.n560 VSUBS 0.009097f
C1286 B.n561 VSUBS 0.009097f
C1287 B.n562 VSUBS 0.009097f
C1288 B.n563 VSUBS 0.009097f
C1289 B.n564 VSUBS 0.009097f
C1290 B.n565 VSUBS 0.009097f
C1291 B.n566 VSUBS 0.009097f
C1292 B.n567 VSUBS 0.009097f
C1293 B.n568 VSUBS 0.009097f
C1294 B.n569 VSUBS 0.009097f
C1295 B.n570 VSUBS 0.009097f
C1296 B.n571 VSUBS 0.009097f
C1297 B.n572 VSUBS 0.009097f
C1298 B.n573 VSUBS 0.009097f
C1299 B.n574 VSUBS 0.009097f
C1300 B.n575 VSUBS 0.009097f
C1301 B.n576 VSUBS 0.009097f
C1302 B.n577 VSUBS 0.009097f
C1303 B.n578 VSUBS 0.009097f
C1304 B.n579 VSUBS 0.009097f
C1305 B.n580 VSUBS 0.009097f
C1306 B.n581 VSUBS 0.009097f
C1307 B.n582 VSUBS 0.009097f
C1308 B.n583 VSUBS 0.009097f
C1309 B.n584 VSUBS 0.009097f
C1310 B.n585 VSUBS 0.008561f
C1311 B.n586 VSUBS 0.021076f
C1312 B.n587 VSUBS 0.005083f
C1313 B.n588 VSUBS 0.009097f
C1314 B.n589 VSUBS 0.009097f
C1315 B.n590 VSUBS 0.009097f
C1316 B.n591 VSUBS 0.009097f
C1317 B.n592 VSUBS 0.009097f
C1318 B.n593 VSUBS 0.009097f
C1319 B.n594 VSUBS 0.009097f
C1320 B.n595 VSUBS 0.009097f
C1321 B.n596 VSUBS 0.009097f
C1322 B.n597 VSUBS 0.009097f
C1323 B.n598 VSUBS 0.009097f
C1324 B.n599 VSUBS 0.009097f
C1325 B.n600 VSUBS 0.005083f
C1326 B.n601 VSUBS 0.009097f
C1327 B.n602 VSUBS 0.009097f
C1328 B.n603 VSUBS 0.008561f
C1329 B.n604 VSUBS 0.009097f
C1330 B.n605 VSUBS 0.009097f
C1331 B.n606 VSUBS 0.009097f
C1332 B.n607 VSUBS 0.009097f
C1333 B.n608 VSUBS 0.009097f
C1334 B.n609 VSUBS 0.009097f
C1335 B.n610 VSUBS 0.009097f
C1336 B.n611 VSUBS 0.009097f
C1337 B.n612 VSUBS 0.009097f
C1338 B.n613 VSUBS 0.009097f
C1339 B.n614 VSUBS 0.009097f
C1340 B.n615 VSUBS 0.009097f
C1341 B.n616 VSUBS 0.009097f
C1342 B.n617 VSUBS 0.009097f
C1343 B.n618 VSUBS 0.009097f
C1344 B.n619 VSUBS 0.009097f
C1345 B.n620 VSUBS 0.009097f
C1346 B.n621 VSUBS 0.009097f
C1347 B.n622 VSUBS 0.009097f
C1348 B.n623 VSUBS 0.009097f
C1349 B.n624 VSUBS 0.009097f
C1350 B.n625 VSUBS 0.009097f
C1351 B.n626 VSUBS 0.009097f
C1352 B.n627 VSUBS 0.009097f
C1353 B.n628 VSUBS 0.009097f
C1354 B.n629 VSUBS 0.009097f
C1355 B.n630 VSUBS 0.009097f
C1356 B.n631 VSUBS 0.009097f
C1357 B.n632 VSUBS 0.009097f
C1358 B.n633 VSUBS 0.009097f
C1359 B.n634 VSUBS 0.009097f
C1360 B.n635 VSUBS 0.009097f
C1361 B.n636 VSUBS 0.009097f
C1362 B.n637 VSUBS 0.009097f
C1363 B.n638 VSUBS 0.009097f
C1364 B.n639 VSUBS 0.009097f
C1365 B.n640 VSUBS 0.009097f
C1366 B.n641 VSUBS 0.009097f
C1367 B.n642 VSUBS 0.009097f
C1368 B.n643 VSUBS 0.009097f
C1369 B.n644 VSUBS 0.009097f
C1370 B.n645 VSUBS 0.009097f
C1371 B.n646 VSUBS 0.009097f
C1372 B.n647 VSUBS 0.009097f
C1373 B.n648 VSUBS 0.009097f
C1374 B.n649 VSUBS 0.009097f
C1375 B.n650 VSUBS 0.009097f
C1376 B.n651 VSUBS 0.009097f
C1377 B.n652 VSUBS 0.009097f
C1378 B.n653 VSUBS 0.009097f
C1379 B.n654 VSUBS 0.009097f
C1380 B.n655 VSUBS 0.009097f
C1381 B.n656 VSUBS 0.009097f
C1382 B.n657 VSUBS 0.009097f
C1383 B.n658 VSUBS 0.022829f
C1384 B.n659 VSUBS 0.021316f
C1385 B.n660 VSUBS 0.021316f
C1386 B.n661 VSUBS 0.009097f
C1387 B.n662 VSUBS 0.009097f
C1388 B.n663 VSUBS 0.009097f
C1389 B.n664 VSUBS 0.009097f
C1390 B.n665 VSUBS 0.009097f
C1391 B.n666 VSUBS 0.009097f
C1392 B.n667 VSUBS 0.009097f
C1393 B.n668 VSUBS 0.009097f
C1394 B.n669 VSUBS 0.009097f
C1395 B.n670 VSUBS 0.009097f
C1396 B.n671 VSUBS 0.009097f
C1397 B.n672 VSUBS 0.009097f
C1398 B.n673 VSUBS 0.009097f
C1399 B.n674 VSUBS 0.009097f
C1400 B.n675 VSUBS 0.009097f
C1401 B.n676 VSUBS 0.009097f
C1402 B.n677 VSUBS 0.009097f
C1403 B.n678 VSUBS 0.009097f
C1404 B.n679 VSUBS 0.009097f
C1405 B.n680 VSUBS 0.009097f
C1406 B.n681 VSUBS 0.009097f
C1407 B.n682 VSUBS 0.009097f
C1408 B.n683 VSUBS 0.009097f
C1409 B.n684 VSUBS 0.009097f
C1410 B.n685 VSUBS 0.009097f
C1411 B.n686 VSUBS 0.009097f
C1412 B.n687 VSUBS 0.009097f
C1413 B.n688 VSUBS 0.009097f
C1414 B.n689 VSUBS 0.009097f
C1415 B.n690 VSUBS 0.009097f
C1416 B.n691 VSUBS 0.009097f
C1417 B.n692 VSUBS 0.009097f
C1418 B.n693 VSUBS 0.009097f
C1419 B.n694 VSUBS 0.009097f
C1420 B.n695 VSUBS 0.009097f
C1421 B.n696 VSUBS 0.009097f
C1422 B.n697 VSUBS 0.009097f
C1423 B.n698 VSUBS 0.009097f
C1424 B.n699 VSUBS 0.009097f
C1425 B.n700 VSUBS 0.009097f
C1426 B.n701 VSUBS 0.009097f
C1427 B.n702 VSUBS 0.009097f
C1428 B.n703 VSUBS 0.009097f
C1429 B.n704 VSUBS 0.009097f
C1430 B.n705 VSUBS 0.009097f
C1431 B.n706 VSUBS 0.009097f
C1432 B.n707 VSUBS 0.009097f
C1433 B.n708 VSUBS 0.009097f
C1434 B.n709 VSUBS 0.009097f
C1435 B.n710 VSUBS 0.009097f
C1436 B.n711 VSUBS 0.009097f
C1437 B.n712 VSUBS 0.009097f
C1438 B.n713 VSUBS 0.009097f
C1439 B.n714 VSUBS 0.009097f
C1440 B.n715 VSUBS 0.009097f
C1441 B.n716 VSUBS 0.009097f
C1442 B.n717 VSUBS 0.009097f
C1443 B.n718 VSUBS 0.009097f
C1444 B.n719 VSUBS 0.009097f
C1445 B.n720 VSUBS 0.009097f
C1446 B.n721 VSUBS 0.009097f
C1447 B.n722 VSUBS 0.009097f
C1448 B.n723 VSUBS 0.009097f
C1449 B.n724 VSUBS 0.009097f
C1450 B.n725 VSUBS 0.009097f
C1451 B.n726 VSUBS 0.009097f
C1452 B.n727 VSUBS 0.01187f
C1453 B.n728 VSUBS 0.012645f
C1454 B.n729 VSUBS 0.025146f
.ends

