* NGSPICE file created from diff_pair_sample_1056.ext - technology: sky130A

.subckt diff_pair_sample_1056 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=2.45025 ps=15.18 w=14.85 l=1.45
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=0 ps=0 w=14.85 l=1.45
X2 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=0 ps=0 w=14.85 l=1.45
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=0 ps=0 w=14.85 l=1.45
X4 VTAIL.t11 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=2.45025 ps=15.18 w=14.85 l=1.45
X5 VDD1.t5 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=2.45025 ps=15.18 w=14.85 l=1.45
X6 VDD2.t3 VN.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=5.7915 ps=30.48 w=14.85 l=1.45
X7 VDD2.t2 VN.t3 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=2.45025 ps=15.18 w=14.85 l=1.45
X8 VTAIL.t1 VP.t1 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=2.45025 ps=15.18 w=14.85 l=1.45
X9 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=0 ps=0 w=14.85 l=1.45
X10 VDD2.t1 VN.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=5.7915 ps=30.48 w=14.85 l=1.45
X11 VTAIL.t5 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=2.45025 ps=15.18 w=14.85 l=1.45
X12 VDD1.t2 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=5.7915 ps=30.48 w=14.85 l=1.45
X13 VDD1.t1 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7915 pd=30.48 as=2.45025 ps=15.18 w=14.85 l=1.45
X14 VTAIL.t9 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=2.45025 ps=15.18 w=14.85 l=1.45
X15 VDD1.t0 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.45025 pd=15.18 as=5.7915 ps=30.48 w=14.85 l=1.45
R0 VN.n3 VN.t0 283.149
R1 VN.n13 VN.t2 283.149
R2 VN.n2 VN.t5 246.817
R3 VN.n8 VN.t4 246.817
R4 VN.n12 VN.t1 246.817
R5 VN.n18 VN.t3 246.817
R6 VN.n9 VN.n8 172.065
R7 VN.n19 VN.n18 172.065
R8 VN.n17 VN.n10 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n11 161.3
R11 VN.n7 VN.n0 161.3
R12 VN.n6 VN.n5 161.3
R13 VN.n4 VN.n1 161.3
R14 VN.n6 VN.n1 51.1773
R15 VN.n16 VN.n11 51.1773
R16 VN VN.n19 46.6766
R17 VN.n3 VN.n2 41.8525
R18 VN.n13 VN.n12 41.8525
R19 VN.n7 VN.n6 29.8095
R20 VN.n17 VN.n16 29.8095
R21 VN.n2 VN.n1 24.4675
R22 VN.n12 VN.n11 24.4675
R23 VN.n14 VN.n13 17.3787
R24 VN.n4 VN.n3 17.3787
R25 VN.n8 VN.n7 13.702
R26 VN.n18 VN.n17 13.702
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VTAIL.n330 VTAIL.n254 289.615
R35 VTAIL.n78 VTAIL.n2 289.615
R36 VTAIL.n248 VTAIL.n172 289.615
R37 VTAIL.n164 VTAIL.n88 289.615
R38 VTAIL.n281 VTAIL.n280 185
R39 VTAIL.n278 VTAIL.n277 185
R40 VTAIL.n287 VTAIL.n286 185
R41 VTAIL.n289 VTAIL.n288 185
R42 VTAIL.n274 VTAIL.n273 185
R43 VTAIL.n295 VTAIL.n294 185
R44 VTAIL.n297 VTAIL.n296 185
R45 VTAIL.n270 VTAIL.n269 185
R46 VTAIL.n303 VTAIL.n302 185
R47 VTAIL.n305 VTAIL.n304 185
R48 VTAIL.n266 VTAIL.n265 185
R49 VTAIL.n311 VTAIL.n310 185
R50 VTAIL.n313 VTAIL.n312 185
R51 VTAIL.n262 VTAIL.n261 185
R52 VTAIL.n319 VTAIL.n318 185
R53 VTAIL.n322 VTAIL.n321 185
R54 VTAIL.n320 VTAIL.n258 185
R55 VTAIL.n327 VTAIL.n257 185
R56 VTAIL.n329 VTAIL.n328 185
R57 VTAIL.n331 VTAIL.n330 185
R58 VTAIL.n29 VTAIL.n28 185
R59 VTAIL.n26 VTAIL.n25 185
R60 VTAIL.n35 VTAIL.n34 185
R61 VTAIL.n37 VTAIL.n36 185
R62 VTAIL.n22 VTAIL.n21 185
R63 VTAIL.n43 VTAIL.n42 185
R64 VTAIL.n45 VTAIL.n44 185
R65 VTAIL.n18 VTAIL.n17 185
R66 VTAIL.n51 VTAIL.n50 185
R67 VTAIL.n53 VTAIL.n52 185
R68 VTAIL.n14 VTAIL.n13 185
R69 VTAIL.n59 VTAIL.n58 185
R70 VTAIL.n61 VTAIL.n60 185
R71 VTAIL.n10 VTAIL.n9 185
R72 VTAIL.n67 VTAIL.n66 185
R73 VTAIL.n70 VTAIL.n69 185
R74 VTAIL.n68 VTAIL.n6 185
R75 VTAIL.n75 VTAIL.n5 185
R76 VTAIL.n77 VTAIL.n76 185
R77 VTAIL.n79 VTAIL.n78 185
R78 VTAIL.n249 VTAIL.n248 185
R79 VTAIL.n247 VTAIL.n246 185
R80 VTAIL.n245 VTAIL.n175 185
R81 VTAIL.n179 VTAIL.n176 185
R82 VTAIL.n240 VTAIL.n239 185
R83 VTAIL.n238 VTAIL.n237 185
R84 VTAIL.n181 VTAIL.n180 185
R85 VTAIL.n232 VTAIL.n231 185
R86 VTAIL.n230 VTAIL.n229 185
R87 VTAIL.n185 VTAIL.n184 185
R88 VTAIL.n224 VTAIL.n223 185
R89 VTAIL.n222 VTAIL.n221 185
R90 VTAIL.n189 VTAIL.n188 185
R91 VTAIL.n216 VTAIL.n215 185
R92 VTAIL.n214 VTAIL.n213 185
R93 VTAIL.n193 VTAIL.n192 185
R94 VTAIL.n208 VTAIL.n207 185
R95 VTAIL.n206 VTAIL.n205 185
R96 VTAIL.n197 VTAIL.n196 185
R97 VTAIL.n200 VTAIL.n199 185
R98 VTAIL.n165 VTAIL.n164 185
R99 VTAIL.n163 VTAIL.n162 185
R100 VTAIL.n161 VTAIL.n91 185
R101 VTAIL.n95 VTAIL.n92 185
R102 VTAIL.n156 VTAIL.n155 185
R103 VTAIL.n154 VTAIL.n153 185
R104 VTAIL.n97 VTAIL.n96 185
R105 VTAIL.n148 VTAIL.n147 185
R106 VTAIL.n146 VTAIL.n145 185
R107 VTAIL.n101 VTAIL.n100 185
R108 VTAIL.n140 VTAIL.n139 185
R109 VTAIL.n138 VTAIL.n137 185
R110 VTAIL.n105 VTAIL.n104 185
R111 VTAIL.n132 VTAIL.n131 185
R112 VTAIL.n130 VTAIL.n129 185
R113 VTAIL.n109 VTAIL.n108 185
R114 VTAIL.n124 VTAIL.n123 185
R115 VTAIL.n122 VTAIL.n121 185
R116 VTAIL.n113 VTAIL.n112 185
R117 VTAIL.n116 VTAIL.n115 185
R118 VTAIL.t2 VTAIL.n198 147.659
R119 VTAIL.t10 VTAIL.n114 147.659
R120 VTAIL.t7 VTAIL.n279 147.659
R121 VTAIL.t4 VTAIL.n27 147.659
R122 VTAIL.n280 VTAIL.n277 104.615
R123 VTAIL.n287 VTAIL.n277 104.615
R124 VTAIL.n288 VTAIL.n287 104.615
R125 VTAIL.n288 VTAIL.n273 104.615
R126 VTAIL.n295 VTAIL.n273 104.615
R127 VTAIL.n296 VTAIL.n295 104.615
R128 VTAIL.n296 VTAIL.n269 104.615
R129 VTAIL.n303 VTAIL.n269 104.615
R130 VTAIL.n304 VTAIL.n303 104.615
R131 VTAIL.n304 VTAIL.n265 104.615
R132 VTAIL.n311 VTAIL.n265 104.615
R133 VTAIL.n312 VTAIL.n311 104.615
R134 VTAIL.n312 VTAIL.n261 104.615
R135 VTAIL.n319 VTAIL.n261 104.615
R136 VTAIL.n321 VTAIL.n319 104.615
R137 VTAIL.n321 VTAIL.n320 104.615
R138 VTAIL.n320 VTAIL.n257 104.615
R139 VTAIL.n329 VTAIL.n257 104.615
R140 VTAIL.n330 VTAIL.n329 104.615
R141 VTAIL.n28 VTAIL.n25 104.615
R142 VTAIL.n35 VTAIL.n25 104.615
R143 VTAIL.n36 VTAIL.n35 104.615
R144 VTAIL.n36 VTAIL.n21 104.615
R145 VTAIL.n43 VTAIL.n21 104.615
R146 VTAIL.n44 VTAIL.n43 104.615
R147 VTAIL.n44 VTAIL.n17 104.615
R148 VTAIL.n51 VTAIL.n17 104.615
R149 VTAIL.n52 VTAIL.n51 104.615
R150 VTAIL.n52 VTAIL.n13 104.615
R151 VTAIL.n59 VTAIL.n13 104.615
R152 VTAIL.n60 VTAIL.n59 104.615
R153 VTAIL.n60 VTAIL.n9 104.615
R154 VTAIL.n67 VTAIL.n9 104.615
R155 VTAIL.n69 VTAIL.n67 104.615
R156 VTAIL.n69 VTAIL.n68 104.615
R157 VTAIL.n68 VTAIL.n5 104.615
R158 VTAIL.n77 VTAIL.n5 104.615
R159 VTAIL.n78 VTAIL.n77 104.615
R160 VTAIL.n248 VTAIL.n247 104.615
R161 VTAIL.n247 VTAIL.n175 104.615
R162 VTAIL.n179 VTAIL.n175 104.615
R163 VTAIL.n239 VTAIL.n179 104.615
R164 VTAIL.n239 VTAIL.n238 104.615
R165 VTAIL.n238 VTAIL.n180 104.615
R166 VTAIL.n231 VTAIL.n180 104.615
R167 VTAIL.n231 VTAIL.n230 104.615
R168 VTAIL.n230 VTAIL.n184 104.615
R169 VTAIL.n223 VTAIL.n184 104.615
R170 VTAIL.n223 VTAIL.n222 104.615
R171 VTAIL.n222 VTAIL.n188 104.615
R172 VTAIL.n215 VTAIL.n188 104.615
R173 VTAIL.n215 VTAIL.n214 104.615
R174 VTAIL.n214 VTAIL.n192 104.615
R175 VTAIL.n207 VTAIL.n192 104.615
R176 VTAIL.n207 VTAIL.n206 104.615
R177 VTAIL.n206 VTAIL.n196 104.615
R178 VTAIL.n199 VTAIL.n196 104.615
R179 VTAIL.n164 VTAIL.n163 104.615
R180 VTAIL.n163 VTAIL.n91 104.615
R181 VTAIL.n95 VTAIL.n91 104.615
R182 VTAIL.n155 VTAIL.n95 104.615
R183 VTAIL.n155 VTAIL.n154 104.615
R184 VTAIL.n154 VTAIL.n96 104.615
R185 VTAIL.n147 VTAIL.n96 104.615
R186 VTAIL.n147 VTAIL.n146 104.615
R187 VTAIL.n146 VTAIL.n100 104.615
R188 VTAIL.n139 VTAIL.n100 104.615
R189 VTAIL.n139 VTAIL.n138 104.615
R190 VTAIL.n138 VTAIL.n104 104.615
R191 VTAIL.n131 VTAIL.n104 104.615
R192 VTAIL.n131 VTAIL.n130 104.615
R193 VTAIL.n130 VTAIL.n108 104.615
R194 VTAIL.n123 VTAIL.n108 104.615
R195 VTAIL.n123 VTAIL.n122 104.615
R196 VTAIL.n122 VTAIL.n112 104.615
R197 VTAIL.n115 VTAIL.n112 104.615
R198 VTAIL.n280 VTAIL.t7 52.3082
R199 VTAIL.n28 VTAIL.t4 52.3082
R200 VTAIL.n199 VTAIL.t2 52.3082
R201 VTAIL.n115 VTAIL.t10 52.3082
R202 VTAIL.n171 VTAIL.n170 48.315
R203 VTAIL.n87 VTAIL.n86 48.315
R204 VTAIL.n1 VTAIL.n0 48.3149
R205 VTAIL.n85 VTAIL.n84 48.3149
R206 VTAIL.n335 VTAIL.n334 36.2581
R207 VTAIL.n83 VTAIL.n82 36.2581
R208 VTAIL.n253 VTAIL.n252 36.2581
R209 VTAIL.n169 VTAIL.n168 36.2581
R210 VTAIL.n87 VTAIL.n85 28.2376
R211 VTAIL.n335 VTAIL.n253 26.7031
R212 VTAIL.n281 VTAIL.n279 15.6677
R213 VTAIL.n29 VTAIL.n27 15.6677
R214 VTAIL.n200 VTAIL.n198 15.6677
R215 VTAIL.n116 VTAIL.n114 15.6677
R216 VTAIL.n328 VTAIL.n327 13.1884
R217 VTAIL.n76 VTAIL.n75 13.1884
R218 VTAIL.n246 VTAIL.n245 13.1884
R219 VTAIL.n162 VTAIL.n161 13.1884
R220 VTAIL.n282 VTAIL.n278 12.8005
R221 VTAIL.n326 VTAIL.n258 12.8005
R222 VTAIL.n331 VTAIL.n256 12.8005
R223 VTAIL.n30 VTAIL.n26 12.8005
R224 VTAIL.n74 VTAIL.n6 12.8005
R225 VTAIL.n79 VTAIL.n4 12.8005
R226 VTAIL.n249 VTAIL.n174 12.8005
R227 VTAIL.n244 VTAIL.n176 12.8005
R228 VTAIL.n201 VTAIL.n197 12.8005
R229 VTAIL.n165 VTAIL.n90 12.8005
R230 VTAIL.n160 VTAIL.n92 12.8005
R231 VTAIL.n117 VTAIL.n113 12.8005
R232 VTAIL.n286 VTAIL.n285 12.0247
R233 VTAIL.n323 VTAIL.n322 12.0247
R234 VTAIL.n332 VTAIL.n254 12.0247
R235 VTAIL.n34 VTAIL.n33 12.0247
R236 VTAIL.n71 VTAIL.n70 12.0247
R237 VTAIL.n80 VTAIL.n2 12.0247
R238 VTAIL.n250 VTAIL.n172 12.0247
R239 VTAIL.n241 VTAIL.n240 12.0247
R240 VTAIL.n205 VTAIL.n204 12.0247
R241 VTAIL.n166 VTAIL.n88 12.0247
R242 VTAIL.n157 VTAIL.n156 12.0247
R243 VTAIL.n121 VTAIL.n120 12.0247
R244 VTAIL.n289 VTAIL.n276 11.249
R245 VTAIL.n318 VTAIL.n260 11.249
R246 VTAIL.n37 VTAIL.n24 11.249
R247 VTAIL.n66 VTAIL.n8 11.249
R248 VTAIL.n237 VTAIL.n178 11.249
R249 VTAIL.n208 VTAIL.n195 11.249
R250 VTAIL.n153 VTAIL.n94 11.249
R251 VTAIL.n124 VTAIL.n111 11.249
R252 VTAIL.n290 VTAIL.n274 10.4732
R253 VTAIL.n317 VTAIL.n262 10.4732
R254 VTAIL.n38 VTAIL.n22 10.4732
R255 VTAIL.n65 VTAIL.n10 10.4732
R256 VTAIL.n236 VTAIL.n181 10.4732
R257 VTAIL.n209 VTAIL.n193 10.4732
R258 VTAIL.n152 VTAIL.n97 10.4732
R259 VTAIL.n125 VTAIL.n109 10.4732
R260 VTAIL.n294 VTAIL.n293 9.69747
R261 VTAIL.n314 VTAIL.n313 9.69747
R262 VTAIL.n42 VTAIL.n41 9.69747
R263 VTAIL.n62 VTAIL.n61 9.69747
R264 VTAIL.n233 VTAIL.n232 9.69747
R265 VTAIL.n213 VTAIL.n212 9.69747
R266 VTAIL.n149 VTAIL.n148 9.69747
R267 VTAIL.n129 VTAIL.n128 9.69747
R268 VTAIL.n334 VTAIL.n333 9.45567
R269 VTAIL.n82 VTAIL.n81 9.45567
R270 VTAIL.n252 VTAIL.n251 9.45567
R271 VTAIL.n168 VTAIL.n167 9.45567
R272 VTAIL.n333 VTAIL.n332 9.3005
R273 VTAIL.n256 VTAIL.n255 9.3005
R274 VTAIL.n301 VTAIL.n300 9.3005
R275 VTAIL.n299 VTAIL.n298 9.3005
R276 VTAIL.n272 VTAIL.n271 9.3005
R277 VTAIL.n293 VTAIL.n292 9.3005
R278 VTAIL.n291 VTAIL.n290 9.3005
R279 VTAIL.n276 VTAIL.n275 9.3005
R280 VTAIL.n285 VTAIL.n284 9.3005
R281 VTAIL.n283 VTAIL.n282 9.3005
R282 VTAIL.n268 VTAIL.n267 9.3005
R283 VTAIL.n307 VTAIL.n306 9.3005
R284 VTAIL.n309 VTAIL.n308 9.3005
R285 VTAIL.n264 VTAIL.n263 9.3005
R286 VTAIL.n315 VTAIL.n314 9.3005
R287 VTAIL.n317 VTAIL.n316 9.3005
R288 VTAIL.n260 VTAIL.n259 9.3005
R289 VTAIL.n324 VTAIL.n323 9.3005
R290 VTAIL.n326 VTAIL.n325 9.3005
R291 VTAIL.n81 VTAIL.n80 9.3005
R292 VTAIL.n4 VTAIL.n3 9.3005
R293 VTAIL.n49 VTAIL.n48 9.3005
R294 VTAIL.n47 VTAIL.n46 9.3005
R295 VTAIL.n20 VTAIL.n19 9.3005
R296 VTAIL.n41 VTAIL.n40 9.3005
R297 VTAIL.n39 VTAIL.n38 9.3005
R298 VTAIL.n24 VTAIL.n23 9.3005
R299 VTAIL.n33 VTAIL.n32 9.3005
R300 VTAIL.n31 VTAIL.n30 9.3005
R301 VTAIL.n16 VTAIL.n15 9.3005
R302 VTAIL.n55 VTAIL.n54 9.3005
R303 VTAIL.n57 VTAIL.n56 9.3005
R304 VTAIL.n12 VTAIL.n11 9.3005
R305 VTAIL.n63 VTAIL.n62 9.3005
R306 VTAIL.n65 VTAIL.n64 9.3005
R307 VTAIL.n8 VTAIL.n7 9.3005
R308 VTAIL.n72 VTAIL.n71 9.3005
R309 VTAIL.n74 VTAIL.n73 9.3005
R310 VTAIL.n226 VTAIL.n225 9.3005
R311 VTAIL.n228 VTAIL.n227 9.3005
R312 VTAIL.n183 VTAIL.n182 9.3005
R313 VTAIL.n234 VTAIL.n233 9.3005
R314 VTAIL.n236 VTAIL.n235 9.3005
R315 VTAIL.n178 VTAIL.n177 9.3005
R316 VTAIL.n242 VTAIL.n241 9.3005
R317 VTAIL.n244 VTAIL.n243 9.3005
R318 VTAIL.n251 VTAIL.n250 9.3005
R319 VTAIL.n174 VTAIL.n173 9.3005
R320 VTAIL.n187 VTAIL.n186 9.3005
R321 VTAIL.n220 VTAIL.n219 9.3005
R322 VTAIL.n218 VTAIL.n217 9.3005
R323 VTAIL.n191 VTAIL.n190 9.3005
R324 VTAIL.n212 VTAIL.n211 9.3005
R325 VTAIL.n210 VTAIL.n209 9.3005
R326 VTAIL.n195 VTAIL.n194 9.3005
R327 VTAIL.n204 VTAIL.n203 9.3005
R328 VTAIL.n202 VTAIL.n201 9.3005
R329 VTAIL.n142 VTAIL.n141 9.3005
R330 VTAIL.n144 VTAIL.n143 9.3005
R331 VTAIL.n99 VTAIL.n98 9.3005
R332 VTAIL.n150 VTAIL.n149 9.3005
R333 VTAIL.n152 VTAIL.n151 9.3005
R334 VTAIL.n94 VTAIL.n93 9.3005
R335 VTAIL.n158 VTAIL.n157 9.3005
R336 VTAIL.n160 VTAIL.n159 9.3005
R337 VTAIL.n167 VTAIL.n166 9.3005
R338 VTAIL.n90 VTAIL.n89 9.3005
R339 VTAIL.n103 VTAIL.n102 9.3005
R340 VTAIL.n136 VTAIL.n135 9.3005
R341 VTAIL.n134 VTAIL.n133 9.3005
R342 VTAIL.n107 VTAIL.n106 9.3005
R343 VTAIL.n128 VTAIL.n127 9.3005
R344 VTAIL.n126 VTAIL.n125 9.3005
R345 VTAIL.n111 VTAIL.n110 9.3005
R346 VTAIL.n120 VTAIL.n119 9.3005
R347 VTAIL.n118 VTAIL.n117 9.3005
R348 VTAIL.n297 VTAIL.n272 8.92171
R349 VTAIL.n310 VTAIL.n264 8.92171
R350 VTAIL.n45 VTAIL.n20 8.92171
R351 VTAIL.n58 VTAIL.n12 8.92171
R352 VTAIL.n229 VTAIL.n183 8.92171
R353 VTAIL.n216 VTAIL.n191 8.92171
R354 VTAIL.n145 VTAIL.n99 8.92171
R355 VTAIL.n132 VTAIL.n107 8.92171
R356 VTAIL.n298 VTAIL.n270 8.14595
R357 VTAIL.n309 VTAIL.n266 8.14595
R358 VTAIL.n46 VTAIL.n18 8.14595
R359 VTAIL.n57 VTAIL.n14 8.14595
R360 VTAIL.n228 VTAIL.n185 8.14595
R361 VTAIL.n217 VTAIL.n189 8.14595
R362 VTAIL.n144 VTAIL.n101 8.14595
R363 VTAIL.n133 VTAIL.n105 8.14595
R364 VTAIL.n302 VTAIL.n301 7.3702
R365 VTAIL.n306 VTAIL.n305 7.3702
R366 VTAIL.n50 VTAIL.n49 7.3702
R367 VTAIL.n54 VTAIL.n53 7.3702
R368 VTAIL.n225 VTAIL.n224 7.3702
R369 VTAIL.n221 VTAIL.n220 7.3702
R370 VTAIL.n141 VTAIL.n140 7.3702
R371 VTAIL.n137 VTAIL.n136 7.3702
R372 VTAIL.n302 VTAIL.n268 6.59444
R373 VTAIL.n305 VTAIL.n268 6.59444
R374 VTAIL.n50 VTAIL.n16 6.59444
R375 VTAIL.n53 VTAIL.n16 6.59444
R376 VTAIL.n224 VTAIL.n187 6.59444
R377 VTAIL.n221 VTAIL.n187 6.59444
R378 VTAIL.n140 VTAIL.n103 6.59444
R379 VTAIL.n137 VTAIL.n103 6.59444
R380 VTAIL.n301 VTAIL.n270 5.81868
R381 VTAIL.n306 VTAIL.n266 5.81868
R382 VTAIL.n49 VTAIL.n18 5.81868
R383 VTAIL.n54 VTAIL.n14 5.81868
R384 VTAIL.n225 VTAIL.n185 5.81868
R385 VTAIL.n220 VTAIL.n189 5.81868
R386 VTAIL.n141 VTAIL.n101 5.81868
R387 VTAIL.n136 VTAIL.n105 5.81868
R388 VTAIL.n298 VTAIL.n297 5.04292
R389 VTAIL.n310 VTAIL.n309 5.04292
R390 VTAIL.n46 VTAIL.n45 5.04292
R391 VTAIL.n58 VTAIL.n57 5.04292
R392 VTAIL.n229 VTAIL.n228 5.04292
R393 VTAIL.n217 VTAIL.n216 5.04292
R394 VTAIL.n145 VTAIL.n144 5.04292
R395 VTAIL.n133 VTAIL.n132 5.04292
R396 VTAIL.n202 VTAIL.n198 4.38563
R397 VTAIL.n118 VTAIL.n114 4.38563
R398 VTAIL.n283 VTAIL.n279 4.38563
R399 VTAIL.n31 VTAIL.n27 4.38563
R400 VTAIL.n294 VTAIL.n272 4.26717
R401 VTAIL.n313 VTAIL.n264 4.26717
R402 VTAIL.n42 VTAIL.n20 4.26717
R403 VTAIL.n61 VTAIL.n12 4.26717
R404 VTAIL.n232 VTAIL.n183 4.26717
R405 VTAIL.n213 VTAIL.n191 4.26717
R406 VTAIL.n148 VTAIL.n99 4.26717
R407 VTAIL.n129 VTAIL.n107 4.26717
R408 VTAIL.n293 VTAIL.n274 3.49141
R409 VTAIL.n314 VTAIL.n262 3.49141
R410 VTAIL.n41 VTAIL.n22 3.49141
R411 VTAIL.n62 VTAIL.n10 3.49141
R412 VTAIL.n233 VTAIL.n181 3.49141
R413 VTAIL.n212 VTAIL.n193 3.49141
R414 VTAIL.n149 VTAIL.n97 3.49141
R415 VTAIL.n128 VTAIL.n109 3.49141
R416 VTAIL.n290 VTAIL.n289 2.71565
R417 VTAIL.n318 VTAIL.n317 2.71565
R418 VTAIL.n38 VTAIL.n37 2.71565
R419 VTAIL.n66 VTAIL.n65 2.71565
R420 VTAIL.n237 VTAIL.n236 2.71565
R421 VTAIL.n209 VTAIL.n208 2.71565
R422 VTAIL.n153 VTAIL.n152 2.71565
R423 VTAIL.n125 VTAIL.n124 2.71565
R424 VTAIL.n286 VTAIL.n276 1.93989
R425 VTAIL.n322 VTAIL.n260 1.93989
R426 VTAIL.n334 VTAIL.n254 1.93989
R427 VTAIL.n34 VTAIL.n24 1.93989
R428 VTAIL.n70 VTAIL.n8 1.93989
R429 VTAIL.n82 VTAIL.n2 1.93989
R430 VTAIL.n252 VTAIL.n172 1.93989
R431 VTAIL.n240 VTAIL.n178 1.93989
R432 VTAIL.n205 VTAIL.n195 1.93989
R433 VTAIL.n168 VTAIL.n88 1.93989
R434 VTAIL.n156 VTAIL.n94 1.93989
R435 VTAIL.n121 VTAIL.n111 1.93989
R436 VTAIL.n169 VTAIL.n87 1.53498
R437 VTAIL.n253 VTAIL.n171 1.53498
R438 VTAIL.n85 VTAIL.n83 1.53498
R439 VTAIL.n0 VTAIL.t6 1.33383
R440 VTAIL.n0 VTAIL.t9 1.33383
R441 VTAIL.n84 VTAIL.t3 1.33383
R442 VTAIL.n84 VTAIL.t1 1.33383
R443 VTAIL.n170 VTAIL.t0 1.33383
R444 VTAIL.n170 VTAIL.t5 1.33383
R445 VTAIL.n86 VTAIL.t8 1.33383
R446 VTAIL.n86 VTAIL.t11 1.33383
R447 VTAIL.n171 VTAIL.n169 1.23757
R448 VTAIL.n83 VTAIL.n1 1.23757
R449 VTAIL.n285 VTAIL.n278 1.16414
R450 VTAIL.n323 VTAIL.n258 1.16414
R451 VTAIL.n332 VTAIL.n331 1.16414
R452 VTAIL.n33 VTAIL.n26 1.16414
R453 VTAIL.n71 VTAIL.n6 1.16414
R454 VTAIL.n80 VTAIL.n79 1.16414
R455 VTAIL.n250 VTAIL.n249 1.16414
R456 VTAIL.n241 VTAIL.n176 1.16414
R457 VTAIL.n204 VTAIL.n197 1.16414
R458 VTAIL.n166 VTAIL.n165 1.16414
R459 VTAIL.n157 VTAIL.n92 1.16414
R460 VTAIL.n120 VTAIL.n113 1.16414
R461 VTAIL VTAIL.n335 1.09317
R462 VTAIL VTAIL.n1 0.44231
R463 VTAIL.n282 VTAIL.n281 0.388379
R464 VTAIL.n327 VTAIL.n326 0.388379
R465 VTAIL.n328 VTAIL.n256 0.388379
R466 VTAIL.n30 VTAIL.n29 0.388379
R467 VTAIL.n75 VTAIL.n74 0.388379
R468 VTAIL.n76 VTAIL.n4 0.388379
R469 VTAIL.n246 VTAIL.n174 0.388379
R470 VTAIL.n245 VTAIL.n244 0.388379
R471 VTAIL.n201 VTAIL.n200 0.388379
R472 VTAIL.n162 VTAIL.n90 0.388379
R473 VTAIL.n161 VTAIL.n160 0.388379
R474 VTAIL.n117 VTAIL.n116 0.388379
R475 VTAIL.n284 VTAIL.n283 0.155672
R476 VTAIL.n284 VTAIL.n275 0.155672
R477 VTAIL.n291 VTAIL.n275 0.155672
R478 VTAIL.n292 VTAIL.n291 0.155672
R479 VTAIL.n292 VTAIL.n271 0.155672
R480 VTAIL.n299 VTAIL.n271 0.155672
R481 VTAIL.n300 VTAIL.n299 0.155672
R482 VTAIL.n300 VTAIL.n267 0.155672
R483 VTAIL.n307 VTAIL.n267 0.155672
R484 VTAIL.n308 VTAIL.n307 0.155672
R485 VTAIL.n308 VTAIL.n263 0.155672
R486 VTAIL.n315 VTAIL.n263 0.155672
R487 VTAIL.n316 VTAIL.n315 0.155672
R488 VTAIL.n316 VTAIL.n259 0.155672
R489 VTAIL.n324 VTAIL.n259 0.155672
R490 VTAIL.n325 VTAIL.n324 0.155672
R491 VTAIL.n325 VTAIL.n255 0.155672
R492 VTAIL.n333 VTAIL.n255 0.155672
R493 VTAIL.n32 VTAIL.n31 0.155672
R494 VTAIL.n32 VTAIL.n23 0.155672
R495 VTAIL.n39 VTAIL.n23 0.155672
R496 VTAIL.n40 VTAIL.n39 0.155672
R497 VTAIL.n40 VTAIL.n19 0.155672
R498 VTAIL.n47 VTAIL.n19 0.155672
R499 VTAIL.n48 VTAIL.n47 0.155672
R500 VTAIL.n48 VTAIL.n15 0.155672
R501 VTAIL.n55 VTAIL.n15 0.155672
R502 VTAIL.n56 VTAIL.n55 0.155672
R503 VTAIL.n56 VTAIL.n11 0.155672
R504 VTAIL.n63 VTAIL.n11 0.155672
R505 VTAIL.n64 VTAIL.n63 0.155672
R506 VTAIL.n64 VTAIL.n7 0.155672
R507 VTAIL.n72 VTAIL.n7 0.155672
R508 VTAIL.n73 VTAIL.n72 0.155672
R509 VTAIL.n73 VTAIL.n3 0.155672
R510 VTAIL.n81 VTAIL.n3 0.155672
R511 VTAIL.n251 VTAIL.n173 0.155672
R512 VTAIL.n243 VTAIL.n173 0.155672
R513 VTAIL.n243 VTAIL.n242 0.155672
R514 VTAIL.n242 VTAIL.n177 0.155672
R515 VTAIL.n235 VTAIL.n177 0.155672
R516 VTAIL.n235 VTAIL.n234 0.155672
R517 VTAIL.n234 VTAIL.n182 0.155672
R518 VTAIL.n227 VTAIL.n182 0.155672
R519 VTAIL.n227 VTAIL.n226 0.155672
R520 VTAIL.n226 VTAIL.n186 0.155672
R521 VTAIL.n219 VTAIL.n186 0.155672
R522 VTAIL.n219 VTAIL.n218 0.155672
R523 VTAIL.n218 VTAIL.n190 0.155672
R524 VTAIL.n211 VTAIL.n190 0.155672
R525 VTAIL.n211 VTAIL.n210 0.155672
R526 VTAIL.n210 VTAIL.n194 0.155672
R527 VTAIL.n203 VTAIL.n194 0.155672
R528 VTAIL.n203 VTAIL.n202 0.155672
R529 VTAIL.n167 VTAIL.n89 0.155672
R530 VTAIL.n159 VTAIL.n89 0.155672
R531 VTAIL.n159 VTAIL.n158 0.155672
R532 VTAIL.n158 VTAIL.n93 0.155672
R533 VTAIL.n151 VTAIL.n93 0.155672
R534 VTAIL.n151 VTAIL.n150 0.155672
R535 VTAIL.n150 VTAIL.n98 0.155672
R536 VTAIL.n143 VTAIL.n98 0.155672
R537 VTAIL.n143 VTAIL.n142 0.155672
R538 VTAIL.n142 VTAIL.n102 0.155672
R539 VTAIL.n135 VTAIL.n102 0.155672
R540 VTAIL.n135 VTAIL.n134 0.155672
R541 VTAIL.n134 VTAIL.n106 0.155672
R542 VTAIL.n127 VTAIL.n106 0.155672
R543 VTAIL.n127 VTAIL.n126 0.155672
R544 VTAIL.n126 VTAIL.n110 0.155672
R545 VTAIL.n119 VTAIL.n110 0.155672
R546 VTAIL.n119 VTAIL.n118 0.155672
R547 VDD2.n159 VDD2.n83 289.615
R548 VDD2.n76 VDD2.n0 289.615
R549 VDD2.n160 VDD2.n159 185
R550 VDD2.n158 VDD2.n157 185
R551 VDD2.n156 VDD2.n86 185
R552 VDD2.n90 VDD2.n87 185
R553 VDD2.n151 VDD2.n150 185
R554 VDD2.n149 VDD2.n148 185
R555 VDD2.n92 VDD2.n91 185
R556 VDD2.n143 VDD2.n142 185
R557 VDD2.n141 VDD2.n140 185
R558 VDD2.n96 VDD2.n95 185
R559 VDD2.n135 VDD2.n134 185
R560 VDD2.n133 VDD2.n132 185
R561 VDD2.n100 VDD2.n99 185
R562 VDD2.n127 VDD2.n126 185
R563 VDD2.n125 VDD2.n124 185
R564 VDD2.n104 VDD2.n103 185
R565 VDD2.n119 VDD2.n118 185
R566 VDD2.n117 VDD2.n116 185
R567 VDD2.n108 VDD2.n107 185
R568 VDD2.n111 VDD2.n110 185
R569 VDD2.n27 VDD2.n26 185
R570 VDD2.n24 VDD2.n23 185
R571 VDD2.n33 VDD2.n32 185
R572 VDD2.n35 VDD2.n34 185
R573 VDD2.n20 VDD2.n19 185
R574 VDD2.n41 VDD2.n40 185
R575 VDD2.n43 VDD2.n42 185
R576 VDD2.n16 VDD2.n15 185
R577 VDD2.n49 VDD2.n48 185
R578 VDD2.n51 VDD2.n50 185
R579 VDD2.n12 VDD2.n11 185
R580 VDD2.n57 VDD2.n56 185
R581 VDD2.n59 VDD2.n58 185
R582 VDD2.n8 VDD2.n7 185
R583 VDD2.n65 VDD2.n64 185
R584 VDD2.n68 VDD2.n67 185
R585 VDD2.n66 VDD2.n4 185
R586 VDD2.n73 VDD2.n3 185
R587 VDD2.n75 VDD2.n74 185
R588 VDD2.n77 VDD2.n76 185
R589 VDD2.t2 VDD2.n109 147.659
R590 VDD2.t5 VDD2.n25 147.659
R591 VDD2.n159 VDD2.n158 104.615
R592 VDD2.n158 VDD2.n86 104.615
R593 VDD2.n90 VDD2.n86 104.615
R594 VDD2.n150 VDD2.n90 104.615
R595 VDD2.n150 VDD2.n149 104.615
R596 VDD2.n149 VDD2.n91 104.615
R597 VDD2.n142 VDD2.n91 104.615
R598 VDD2.n142 VDD2.n141 104.615
R599 VDD2.n141 VDD2.n95 104.615
R600 VDD2.n134 VDD2.n95 104.615
R601 VDD2.n134 VDD2.n133 104.615
R602 VDD2.n133 VDD2.n99 104.615
R603 VDD2.n126 VDD2.n99 104.615
R604 VDD2.n126 VDD2.n125 104.615
R605 VDD2.n125 VDD2.n103 104.615
R606 VDD2.n118 VDD2.n103 104.615
R607 VDD2.n118 VDD2.n117 104.615
R608 VDD2.n117 VDD2.n107 104.615
R609 VDD2.n110 VDD2.n107 104.615
R610 VDD2.n26 VDD2.n23 104.615
R611 VDD2.n33 VDD2.n23 104.615
R612 VDD2.n34 VDD2.n33 104.615
R613 VDD2.n34 VDD2.n19 104.615
R614 VDD2.n41 VDD2.n19 104.615
R615 VDD2.n42 VDD2.n41 104.615
R616 VDD2.n42 VDD2.n15 104.615
R617 VDD2.n49 VDD2.n15 104.615
R618 VDD2.n50 VDD2.n49 104.615
R619 VDD2.n50 VDD2.n11 104.615
R620 VDD2.n57 VDD2.n11 104.615
R621 VDD2.n58 VDD2.n57 104.615
R622 VDD2.n58 VDD2.n7 104.615
R623 VDD2.n65 VDD2.n7 104.615
R624 VDD2.n67 VDD2.n65 104.615
R625 VDD2.n67 VDD2.n66 104.615
R626 VDD2.n66 VDD2.n3 104.615
R627 VDD2.n75 VDD2.n3 104.615
R628 VDD2.n76 VDD2.n75 104.615
R629 VDD2.n82 VDD2.n81 65.3219
R630 VDD2 VDD2.n165 65.3191
R631 VDD2.n82 VDD2.n80 54.0324
R632 VDD2.n164 VDD2.n163 52.9369
R633 VDD2.n110 VDD2.t2 52.3082
R634 VDD2.n26 VDD2.t5 52.3082
R635 VDD2.n164 VDD2.n82 41.5041
R636 VDD2.n111 VDD2.n109 15.6677
R637 VDD2.n27 VDD2.n25 15.6677
R638 VDD2.n157 VDD2.n156 13.1884
R639 VDD2.n74 VDD2.n73 13.1884
R640 VDD2.n160 VDD2.n85 12.8005
R641 VDD2.n155 VDD2.n87 12.8005
R642 VDD2.n112 VDD2.n108 12.8005
R643 VDD2.n28 VDD2.n24 12.8005
R644 VDD2.n72 VDD2.n4 12.8005
R645 VDD2.n77 VDD2.n2 12.8005
R646 VDD2.n161 VDD2.n83 12.0247
R647 VDD2.n152 VDD2.n151 12.0247
R648 VDD2.n116 VDD2.n115 12.0247
R649 VDD2.n32 VDD2.n31 12.0247
R650 VDD2.n69 VDD2.n68 12.0247
R651 VDD2.n78 VDD2.n0 12.0247
R652 VDD2.n148 VDD2.n89 11.249
R653 VDD2.n119 VDD2.n106 11.249
R654 VDD2.n35 VDD2.n22 11.249
R655 VDD2.n64 VDD2.n6 11.249
R656 VDD2.n147 VDD2.n92 10.4732
R657 VDD2.n120 VDD2.n104 10.4732
R658 VDD2.n36 VDD2.n20 10.4732
R659 VDD2.n63 VDD2.n8 10.4732
R660 VDD2.n144 VDD2.n143 9.69747
R661 VDD2.n124 VDD2.n123 9.69747
R662 VDD2.n40 VDD2.n39 9.69747
R663 VDD2.n60 VDD2.n59 9.69747
R664 VDD2.n163 VDD2.n162 9.45567
R665 VDD2.n80 VDD2.n79 9.45567
R666 VDD2.n137 VDD2.n136 9.3005
R667 VDD2.n139 VDD2.n138 9.3005
R668 VDD2.n94 VDD2.n93 9.3005
R669 VDD2.n145 VDD2.n144 9.3005
R670 VDD2.n147 VDD2.n146 9.3005
R671 VDD2.n89 VDD2.n88 9.3005
R672 VDD2.n153 VDD2.n152 9.3005
R673 VDD2.n155 VDD2.n154 9.3005
R674 VDD2.n162 VDD2.n161 9.3005
R675 VDD2.n85 VDD2.n84 9.3005
R676 VDD2.n98 VDD2.n97 9.3005
R677 VDD2.n131 VDD2.n130 9.3005
R678 VDD2.n129 VDD2.n128 9.3005
R679 VDD2.n102 VDD2.n101 9.3005
R680 VDD2.n123 VDD2.n122 9.3005
R681 VDD2.n121 VDD2.n120 9.3005
R682 VDD2.n106 VDD2.n105 9.3005
R683 VDD2.n115 VDD2.n114 9.3005
R684 VDD2.n113 VDD2.n112 9.3005
R685 VDD2.n79 VDD2.n78 9.3005
R686 VDD2.n2 VDD2.n1 9.3005
R687 VDD2.n47 VDD2.n46 9.3005
R688 VDD2.n45 VDD2.n44 9.3005
R689 VDD2.n18 VDD2.n17 9.3005
R690 VDD2.n39 VDD2.n38 9.3005
R691 VDD2.n37 VDD2.n36 9.3005
R692 VDD2.n22 VDD2.n21 9.3005
R693 VDD2.n31 VDD2.n30 9.3005
R694 VDD2.n29 VDD2.n28 9.3005
R695 VDD2.n14 VDD2.n13 9.3005
R696 VDD2.n53 VDD2.n52 9.3005
R697 VDD2.n55 VDD2.n54 9.3005
R698 VDD2.n10 VDD2.n9 9.3005
R699 VDD2.n61 VDD2.n60 9.3005
R700 VDD2.n63 VDD2.n62 9.3005
R701 VDD2.n6 VDD2.n5 9.3005
R702 VDD2.n70 VDD2.n69 9.3005
R703 VDD2.n72 VDD2.n71 9.3005
R704 VDD2.n140 VDD2.n94 8.92171
R705 VDD2.n127 VDD2.n102 8.92171
R706 VDD2.n43 VDD2.n18 8.92171
R707 VDD2.n56 VDD2.n10 8.92171
R708 VDD2.n139 VDD2.n96 8.14595
R709 VDD2.n128 VDD2.n100 8.14595
R710 VDD2.n44 VDD2.n16 8.14595
R711 VDD2.n55 VDD2.n12 8.14595
R712 VDD2.n136 VDD2.n135 7.3702
R713 VDD2.n132 VDD2.n131 7.3702
R714 VDD2.n48 VDD2.n47 7.3702
R715 VDD2.n52 VDD2.n51 7.3702
R716 VDD2.n135 VDD2.n98 6.59444
R717 VDD2.n132 VDD2.n98 6.59444
R718 VDD2.n48 VDD2.n14 6.59444
R719 VDD2.n51 VDD2.n14 6.59444
R720 VDD2.n136 VDD2.n96 5.81868
R721 VDD2.n131 VDD2.n100 5.81868
R722 VDD2.n47 VDD2.n16 5.81868
R723 VDD2.n52 VDD2.n12 5.81868
R724 VDD2.n140 VDD2.n139 5.04292
R725 VDD2.n128 VDD2.n127 5.04292
R726 VDD2.n44 VDD2.n43 5.04292
R727 VDD2.n56 VDD2.n55 5.04292
R728 VDD2.n113 VDD2.n109 4.38563
R729 VDD2.n29 VDD2.n25 4.38563
R730 VDD2.n143 VDD2.n94 4.26717
R731 VDD2.n124 VDD2.n102 4.26717
R732 VDD2.n40 VDD2.n18 4.26717
R733 VDD2.n59 VDD2.n10 4.26717
R734 VDD2.n144 VDD2.n92 3.49141
R735 VDD2.n123 VDD2.n104 3.49141
R736 VDD2.n39 VDD2.n20 3.49141
R737 VDD2.n60 VDD2.n8 3.49141
R738 VDD2.n148 VDD2.n147 2.71565
R739 VDD2.n120 VDD2.n119 2.71565
R740 VDD2.n36 VDD2.n35 2.71565
R741 VDD2.n64 VDD2.n63 2.71565
R742 VDD2.n163 VDD2.n83 1.93989
R743 VDD2.n151 VDD2.n89 1.93989
R744 VDD2.n116 VDD2.n106 1.93989
R745 VDD2.n32 VDD2.n22 1.93989
R746 VDD2.n68 VDD2.n6 1.93989
R747 VDD2.n80 VDD2.n0 1.93989
R748 VDD2.n165 VDD2.t4 1.33383
R749 VDD2.n165 VDD2.t3 1.33383
R750 VDD2.n81 VDD2.t0 1.33383
R751 VDD2.n81 VDD2.t1 1.33383
R752 VDD2 VDD2.n164 1.20955
R753 VDD2.n161 VDD2.n160 1.16414
R754 VDD2.n152 VDD2.n87 1.16414
R755 VDD2.n115 VDD2.n108 1.16414
R756 VDD2.n31 VDD2.n24 1.16414
R757 VDD2.n69 VDD2.n4 1.16414
R758 VDD2.n78 VDD2.n77 1.16414
R759 VDD2.n157 VDD2.n85 0.388379
R760 VDD2.n156 VDD2.n155 0.388379
R761 VDD2.n112 VDD2.n111 0.388379
R762 VDD2.n28 VDD2.n27 0.388379
R763 VDD2.n73 VDD2.n72 0.388379
R764 VDD2.n74 VDD2.n2 0.388379
R765 VDD2.n162 VDD2.n84 0.155672
R766 VDD2.n154 VDD2.n84 0.155672
R767 VDD2.n154 VDD2.n153 0.155672
R768 VDD2.n153 VDD2.n88 0.155672
R769 VDD2.n146 VDD2.n88 0.155672
R770 VDD2.n146 VDD2.n145 0.155672
R771 VDD2.n145 VDD2.n93 0.155672
R772 VDD2.n138 VDD2.n93 0.155672
R773 VDD2.n138 VDD2.n137 0.155672
R774 VDD2.n137 VDD2.n97 0.155672
R775 VDD2.n130 VDD2.n97 0.155672
R776 VDD2.n130 VDD2.n129 0.155672
R777 VDD2.n129 VDD2.n101 0.155672
R778 VDD2.n122 VDD2.n101 0.155672
R779 VDD2.n122 VDD2.n121 0.155672
R780 VDD2.n121 VDD2.n105 0.155672
R781 VDD2.n114 VDD2.n105 0.155672
R782 VDD2.n114 VDD2.n113 0.155672
R783 VDD2.n30 VDD2.n29 0.155672
R784 VDD2.n30 VDD2.n21 0.155672
R785 VDD2.n37 VDD2.n21 0.155672
R786 VDD2.n38 VDD2.n37 0.155672
R787 VDD2.n38 VDD2.n17 0.155672
R788 VDD2.n45 VDD2.n17 0.155672
R789 VDD2.n46 VDD2.n45 0.155672
R790 VDD2.n46 VDD2.n13 0.155672
R791 VDD2.n53 VDD2.n13 0.155672
R792 VDD2.n54 VDD2.n53 0.155672
R793 VDD2.n54 VDD2.n9 0.155672
R794 VDD2.n61 VDD2.n9 0.155672
R795 VDD2.n62 VDD2.n61 0.155672
R796 VDD2.n62 VDD2.n5 0.155672
R797 VDD2.n70 VDD2.n5 0.155672
R798 VDD2.n71 VDD2.n70 0.155672
R799 VDD2.n71 VDD2.n1 0.155672
R800 VDD2.n79 VDD2.n1 0.155672
R801 B.n795 B.n794 585
R802 B.n333 B.n110 585
R803 B.n332 B.n331 585
R804 B.n330 B.n329 585
R805 B.n328 B.n327 585
R806 B.n326 B.n325 585
R807 B.n324 B.n323 585
R808 B.n322 B.n321 585
R809 B.n320 B.n319 585
R810 B.n318 B.n317 585
R811 B.n316 B.n315 585
R812 B.n314 B.n313 585
R813 B.n312 B.n311 585
R814 B.n310 B.n309 585
R815 B.n308 B.n307 585
R816 B.n306 B.n305 585
R817 B.n304 B.n303 585
R818 B.n302 B.n301 585
R819 B.n300 B.n299 585
R820 B.n298 B.n297 585
R821 B.n296 B.n295 585
R822 B.n294 B.n293 585
R823 B.n292 B.n291 585
R824 B.n290 B.n289 585
R825 B.n288 B.n287 585
R826 B.n286 B.n285 585
R827 B.n284 B.n283 585
R828 B.n282 B.n281 585
R829 B.n280 B.n279 585
R830 B.n278 B.n277 585
R831 B.n276 B.n275 585
R832 B.n274 B.n273 585
R833 B.n272 B.n271 585
R834 B.n270 B.n269 585
R835 B.n268 B.n267 585
R836 B.n266 B.n265 585
R837 B.n264 B.n263 585
R838 B.n262 B.n261 585
R839 B.n260 B.n259 585
R840 B.n258 B.n257 585
R841 B.n256 B.n255 585
R842 B.n254 B.n253 585
R843 B.n252 B.n251 585
R844 B.n250 B.n249 585
R845 B.n248 B.n247 585
R846 B.n246 B.n245 585
R847 B.n244 B.n243 585
R848 B.n242 B.n241 585
R849 B.n240 B.n239 585
R850 B.n238 B.n237 585
R851 B.n236 B.n235 585
R852 B.n234 B.n233 585
R853 B.n232 B.n231 585
R854 B.n230 B.n229 585
R855 B.n228 B.n227 585
R856 B.n226 B.n225 585
R857 B.n224 B.n223 585
R858 B.n222 B.n221 585
R859 B.n220 B.n219 585
R860 B.n218 B.n217 585
R861 B.n216 B.n215 585
R862 B.n214 B.n213 585
R863 B.n212 B.n211 585
R864 B.n210 B.n209 585
R865 B.n208 B.n207 585
R866 B.n206 B.n205 585
R867 B.n204 B.n203 585
R868 B.n202 B.n201 585
R869 B.n200 B.n199 585
R870 B.n198 B.n197 585
R871 B.n196 B.n195 585
R872 B.n194 B.n193 585
R873 B.n192 B.n191 585
R874 B.n190 B.n189 585
R875 B.n188 B.n187 585
R876 B.n186 B.n185 585
R877 B.n184 B.n183 585
R878 B.n182 B.n181 585
R879 B.n180 B.n179 585
R880 B.n178 B.n177 585
R881 B.n176 B.n175 585
R882 B.n174 B.n173 585
R883 B.n172 B.n171 585
R884 B.n170 B.n169 585
R885 B.n168 B.n167 585
R886 B.n166 B.n165 585
R887 B.n164 B.n163 585
R888 B.n162 B.n161 585
R889 B.n160 B.n159 585
R890 B.n158 B.n157 585
R891 B.n156 B.n155 585
R892 B.n154 B.n153 585
R893 B.n152 B.n151 585
R894 B.n150 B.n149 585
R895 B.n148 B.n147 585
R896 B.n146 B.n145 585
R897 B.n144 B.n143 585
R898 B.n142 B.n141 585
R899 B.n140 B.n139 585
R900 B.n138 B.n137 585
R901 B.n136 B.n135 585
R902 B.n134 B.n133 585
R903 B.n132 B.n131 585
R904 B.n130 B.n129 585
R905 B.n128 B.n127 585
R906 B.n126 B.n125 585
R907 B.n124 B.n123 585
R908 B.n122 B.n121 585
R909 B.n120 B.n119 585
R910 B.n118 B.n117 585
R911 B.n793 B.n55 585
R912 B.n798 B.n55 585
R913 B.n792 B.n54 585
R914 B.n799 B.n54 585
R915 B.n791 B.n790 585
R916 B.n790 B.n50 585
R917 B.n789 B.n49 585
R918 B.n805 B.n49 585
R919 B.n788 B.n48 585
R920 B.n806 B.n48 585
R921 B.n787 B.n47 585
R922 B.n807 B.n47 585
R923 B.n786 B.n785 585
R924 B.n785 B.n43 585
R925 B.n784 B.n42 585
R926 B.n813 B.n42 585
R927 B.n783 B.n41 585
R928 B.n814 B.n41 585
R929 B.n782 B.n40 585
R930 B.n815 B.n40 585
R931 B.n781 B.n780 585
R932 B.n780 B.n36 585
R933 B.n779 B.n35 585
R934 B.n821 B.n35 585
R935 B.n778 B.n34 585
R936 B.n822 B.n34 585
R937 B.n777 B.n33 585
R938 B.n823 B.n33 585
R939 B.n776 B.n775 585
R940 B.n775 B.n32 585
R941 B.n774 B.n28 585
R942 B.n829 B.n28 585
R943 B.n773 B.n27 585
R944 B.n830 B.n27 585
R945 B.n772 B.n26 585
R946 B.n831 B.n26 585
R947 B.n771 B.n770 585
R948 B.n770 B.n22 585
R949 B.n769 B.n21 585
R950 B.n837 B.n21 585
R951 B.n768 B.n20 585
R952 B.n838 B.n20 585
R953 B.n767 B.n19 585
R954 B.n839 B.n19 585
R955 B.n766 B.n765 585
R956 B.n765 B.n15 585
R957 B.n764 B.n14 585
R958 B.n845 B.n14 585
R959 B.n763 B.n13 585
R960 B.n846 B.n13 585
R961 B.n762 B.n12 585
R962 B.n847 B.n12 585
R963 B.n761 B.n760 585
R964 B.n760 B.n8 585
R965 B.n759 B.n7 585
R966 B.n853 B.n7 585
R967 B.n758 B.n6 585
R968 B.n854 B.n6 585
R969 B.n757 B.n5 585
R970 B.n855 B.n5 585
R971 B.n756 B.n755 585
R972 B.n755 B.n4 585
R973 B.n754 B.n334 585
R974 B.n754 B.n753 585
R975 B.n744 B.n335 585
R976 B.n336 B.n335 585
R977 B.n746 B.n745 585
R978 B.n747 B.n746 585
R979 B.n743 B.n340 585
R980 B.n344 B.n340 585
R981 B.n742 B.n741 585
R982 B.n741 B.n740 585
R983 B.n342 B.n341 585
R984 B.n343 B.n342 585
R985 B.n733 B.n732 585
R986 B.n734 B.n733 585
R987 B.n731 B.n349 585
R988 B.n349 B.n348 585
R989 B.n730 B.n729 585
R990 B.n729 B.n728 585
R991 B.n351 B.n350 585
R992 B.n352 B.n351 585
R993 B.n721 B.n720 585
R994 B.n722 B.n721 585
R995 B.n719 B.n357 585
R996 B.n357 B.n356 585
R997 B.n718 B.n717 585
R998 B.n717 B.n716 585
R999 B.n359 B.n358 585
R1000 B.n709 B.n359 585
R1001 B.n708 B.n707 585
R1002 B.n710 B.n708 585
R1003 B.n706 B.n364 585
R1004 B.n364 B.n363 585
R1005 B.n705 B.n704 585
R1006 B.n704 B.n703 585
R1007 B.n366 B.n365 585
R1008 B.n367 B.n366 585
R1009 B.n696 B.n695 585
R1010 B.n697 B.n696 585
R1011 B.n694 B.n372 585
R1012 B.n372 B.n371 585
R1013 B.n693 B.n692 585
R1014 B.n692 B.n691 585
R1015 B.n374 B.n373 585
R1016 B.n375 B.n374 585
R1017 B.n684 B.n683 585
R1018 B.n685 B.n684 585
R1019 B.n682 B.n380 585
R1020 B.n380 B.n379 585
R1021 B.n681 B.n680 585
R1022 B.n680 B.n679 585
R1023 B.n382 B.n381 585
R1024 B.n383 B.n382 585
R1025 B.n672 B.n671 585
R1026 B.n673 B.n672 585
R1027 B.n670 B.n388 585
R1028 B.n388 B.n387 585
R1029 B.n665 B.n664 585
R1030 B.n663 B.n445 585
R1031 B.n662 B.n444 585
R1032 B.n667 B.n444 585
R1033 B.n661 B.n660 585
R1034 B.n659 B.n658 585
R1035 B.n657 B.n656 585
R1036 B.n655 B.n654 585
R1037 B.n653 B.n652 585
R1038 B.n651 B.n650 585
R1039 B.n649 B.n648 585
R1040 B.n647 B.n646 585
R1041 B.n645 B.n644 585
R1042 B.n643 B.n642 585
R1043 B.n641 B.n640 585
R1044 B.n639 B.n638 585
R1045 B.n637 B.n636 585
R1046 B.n635 B.n634 585
R1047 B.n633 B.n632 585
R1048 B.n631 B.n630 585
R1049 B.n629 B.n628 585
R1050 B.n627 B.n626 585
R1051 B.n625 B.n624 585
R1052 B.n623 B.n622 585
R1053 B.n621 B.n620 585
R1054 B.n619 B.n618 585
R1055 B.n617 B.n616 585
R1056 B.n615 B.n614 585
R1057 B.n613 B.n612 585
R1058 B.n611 B.n610 585
R1059 B.n609 B.n608 585
R1060 B.n607 B.n606 585
R1061 B.n605 B.n604 585
R1062 B.n603 B.n602 585
R1063 B.n601 B.n600 585
R1064 B.n599 B.n598 585
R1065 B.n597 B.n596 585
R1066 B.n595 B.n594 585
R1067 B.n593 B.n592 585
R1068 B.n591 B.n590 585
R1069 B.n589 B.n588 585
R1070 B.n587 B.n586 585
R1071 B.n585 B.n584 585
R1072 B.n583 B.n582 585
R1073 B.n581 B.n580 585
R1074 B.n579 B.n578 585
R1075 B.n577 B.n576 585
R1076 B.n575 B.n574 585
R1077 B.n573 B.n572 585
R1078 B.n571 B.n570 585
R1079 B.n569 B.n568 585
R1080 B.n566 B.n565 585
R1081 B.n564 B.n563 585
R1082 B.n562 B.n561 585
R1083 B.n560 B.n559 585
R1084 B.n558 B.n557 585
R1085 B.n556 B.n555 585
R1086 B.n554 B.n553 585
R1087 B.n552 B.n551 585
R1088 B.n550 B.n549 585
R1089 B.n548 B.n547 585
R1090 B.n545 B.n544 585
R1091 B.n543 B.n542 585
R1092 B.n541 B.n540 585
R1093 B.n539 B.n538 585
R1094 B.n537 B.n536 585
R1095 B.n535 B.n534 585
R1096 B.n533 B.n532 585
R1097 B.n531 B.n530 585
R1098 B.n529 B.n528 585
R1099 B.n527 B.n526 585
R1100 B.n525 B.n524 585
R1101 B.n523 B.n522 585
R1102 B.n521 B.n520 585
R1103 B.n519 B.n518 585
R1104 B.n517 B.n516 585
R1105 B.n515 B.n514 585
R1106 B.n513 B.n512 585
R1107 B.n511 B.n510 585
R1108 B.n509 B.n508 585
R1109 B.n507 B.n506 585
R1110 B.n505 B.n504 585
R1111 B.n503 B.n502 585
R1112 B.n501 B.n500 585
R1113 B.n499 B.n498 585
R1114 B.n497 B.n496 585
R1115 B.n495 B.n494 585
R1116 B.n493 B.n492 585
R1117 B.n491 B.n490 585
R1118 B.n489 B.n488 585
R1119 B.n487 B.n486 585
R1120 B.n485 B.n484 585
R1121 B.n483 B.n482 585
R1122 B.n481 B.n480 585
R1123 B.n479 B.n478 585
R1124 B.n477 B.n476 585
R1125 B.n475 B.n474 585
R1126 B.n473 B.n472 585
R1127 B.n471 B.n470 585
R1128 B.n469 B.n468 585
R1129 B.n467 B.n466 585
R1130 B.n465 B.n464 585
R1131 B.n463 B.n462 585
R1132 B.n461 B.n460 585
R1133 B.n459 B.n458 585
R1134 B.n457 B.n456 585
R1135 B.n455 B.n454 585
R1136 B.n453 B.n452 585
R1137 B.n451 B.n450 585
R1138 B.n390 B.n389 585
R1139 B.n669 B.n668 585
R1140 B.n668 B.n667 585
R1141 B.n386 B.n385 585
R1142 B.n387 B.n386 585
R1143 B.n675 B.n674 585
R1144 B.n674 B.n673 585
R1145 B.n676 B.n384 585
R1146 B.n384 B.n383 585
R1147 B.n678 B.n677 585
R1148 B.n679 B.n678 585
R1149 B.n378 B.n377 585
R1150 B.n379 B.n378 585
R1151 B.n687 B.n686 585
R1152 B.n686 B.n685 585
R1153 B.n688 B.n376 585
R1154 B.n376 B.n375 585
R1155 B.n690 B.n689 585
R1156 B.n691 B.n690 585
R1157 B.n370 B.n369 585
R1158 B.n371 B.n370 585
R1159 B.n699 B.n698 585
R1160 B.n698 B.n697 585
R1161 B.n700 B.n368 585
R1162 B.n368 B.n367 585
R1163 B.n702 B.n701 585
R1164 B.n703 B.n702 585
R1165 B.n362 B.n361 585
R1166 B.n363 B.n362 585
R1167 B.n712 B.n711 585
R1168 B.n711 B.n710 585
R1169 B.n713 B.n360 585
R1170 B.n709 B.n360 585
R1171 B.n715 B.n714 585
R1172 B.n716 B.n715 585
R1173 B.n355 B.n354 585
R1174 B.n356 B.n355 585
R1175 B.n724 B.n723 585
R1176 B.n723 B.n722 585
R1177 B.n725 B.n353 585
R1178 B.n353 B.n352 585
R1179 B.n727 B.n726 585
R1180 B.n728 B.n727 585
R1181 B.n347 B.n346 585
R1182 B.n348 B.n347 585
R1183 B.n736 B.n735 585
R1184 B.n735 B.n734 585
R1185 B.n737 B.n345 585
R1186 B.n345 B.n343 585
R1187 B.n739 B.n738 585
R1188 B.n740 B.n739 585
R1189 B.n339 B.n338 585
R1190 B.n344 B.n339 585
R1191 B.n749 B.n748 585
R1192 B.n748 B.n747 585
R1193 B.n750 B.n337 585
R1194 B.n337 B.n336 585
R1195 B.n752 B.n751 585
R1196 B.n753 B.n752 585
R1197 B.n2 B.n0 585
R1198 B.n4 B.n2 585
R1199 B.n3 B.n1 585
R1200 B.n854 B.n3 585
R1201 B.n852 B.n851 585
R1202 B.n853 B.n852 585
R1203 B.n850 B.n9 585
R1204 B.n9 B.n8 585
R1205 B.n849 B.n848 585
R1206 B.n848 B.n847 585
R1207 B.n11 B.n10 585
R1208 B.n846 B.n11 585
R1209 B.n844 B.n843 585
R1210 B.n845 B.n844 585
R1211 B.n842 B.n16 585
R1212 B.n16 B.n15 585
R1213 B.n841 B.n840 585
R1214 B.n840 B.n839 585
R1215 B.n18 B.n17 585
R1216 B.n838 B.n18 585
R1217 B.n836 B.n835 585
R1218 B.n837 B.n836 585
R1219 B.n834 B.n23 585
R1220 B.n23 B.n22 585
R1221 B.n833 B.n832 585
R1222 B.n832 B.n831 585
R1223 B.n25 B.n24 585
R1224 B.n830 B.n25 585
R1225 B.n828 B.n827 585
R1226 B.n829 B.n828 585
R1227 B.n826 B.n29 585
R1228 B.n32 B.n29 585
R1229 B.n825 B.n824 585
R1230 B.n824 B.n823 585
R1231 B.n31 B.n30 585
R1232 B.n822 B.n31 585
R1233 B.n820 B.n819 585
R1234 B.n821 B.n820 585
R1235 B.n818 B.n37 585
R1236 B.n37 B.n36 585
R1237 B.n817 B.n816 585
R1238 B.n816 B.n815 585
R1239 B.n39 B.n38 585
R1240 B.n814 B.n39 585
R1241 B.n812 B.n811 585
R1242 B.n813 B.n812 585
R1243 B.n810 B.n44 585
R1244 B.n44 B.n43 585
R1245 B.n809 B.n808 585
R1246 B.n808 B.n807 585
R1247 B.n46 B.n45 585
R1248 B.n806 B.n46 585
R1249 B.n804 B.n803 585
R1250 B.n805 B.n804 585
R1251 B.n802 B.n51 585
R1252 B.n51 B.n50 585
R1253 B.n801 B.n800 585
R1254 B.n800 B.n799 585
R1255 B.n53 B.n52 585
R1256 B.n798 B.n53 585
R1257 B.n857 B.n856 585
R1258 B.n856 B.n855 585
R1259 B.n665 B.n386 473.281
R1260 B.n117 B.n53 473.281
R1261 B.n668 B.n388 473.281
R1262 B.n795 B.n55 473.281
R1263 B.n448 B.t17 452.067
R1264 B.n446 B.t13 452.067
R1265 B.n114 B.t10 452.067
R1266 B.n111 B.t6 452.067
R1267 B.n448 B.t19 365.901
R1268 B.n446 B.t16 365.901
R1269 B.n114 B.t11 365.901
R1270 B.n111 B.t8 365.901
R1271 B.n449 B.t18 331.38
R1272 B.n112 B.t9 331.38
R1273 B.n447 B.t15 331.378
R1274 B.n115 B.t12 331.378
R1275 B.n797 B.n796 256.663
R1276 B.n797 B.n109 256.663
R1277 B.n797 B.n108 256.663
R1278 B.n797 B.n107 256.663
R1279 B.n797 B.n106 256.663
R1280 B.n797 B.n105 256.663
R1281 B.n797 B.n104 256.663
R1282 B.n797 B.n103 256.663
R1283 B.n797 B.n102 256.663
R1284 B.n797 B.n101 256.663
R1285 B.n797 B.n100 256.663
R1286 B.n797 B.n99 256.663
R1287 B.n797 B.n98 256.663
R1288 B.n797 B.n97 256.663
R1289 B.n797 B.n96 256.663
R1290 B.n797 B.n95 256.663
R1291 B.n797 B.n94 256.663
R1292 B.n797 B.n93 256.663
R1293 B.n797 B.n92 256.663
R1294 B.n797 B.n91 256.663
R1295 B.n797 B.n90 256.663
R1296 B.n797 B.n89 256.663
R1297 B.n797 B.n88 256.663
R1298 B.n797 B.n87 256.663
R1299 B.n797 B.n86 256.663
R1300 B.n797 B.n85 256.663
R1301 B.n797 B.n84 256.663
R1302 B.n797 B.n83 256.663
R1303 B.n797 B.n82 256.663
R1304 B.n797 B.n81 256.663
R1305 B.n797 B.n80 256.663
R1306 B.n797 B.n79 256.663
R1307 B.n797 B.n78 256.663
R1308 B.n797 B.n77 256.663
R1309 B.n797 B.n76 256.663
R1310 B.n797 B.n75 256.663
R1311 B.n797 B.n74 256.663
R1312 B.n797 B.n73 256.663
R1313 B.n797 B.n72 256.663
R1314 B.n797 B.n71 256.663
R1315 B.n797 B.n70 256.663
R1316 B.n797 B.n69 256.663
R1317 B.n797 B.n68 256.663
R1318 B.n797 B.n67 256.663
R1319 B.n797 B.n66 256.663
R1320 B.n797 B.n65 256.663
R1321 B.n797 B.n64 256.663
R1322 B.n797 B.n63 256.663
R1323 B.n797 B.n62 256.663
R1324 B.n797 B.n61 256.663
R1325 B.n797 B.n60 256.663
R1326 B.n797 B.n59 256.663
R1327 B.n797 B.n58 256.663
R1328 B.n797 B.n57 256.663
R1329 B.n797 B.n56 256.663
R1330 B.n667 B.n666 256.663
R1331 B.n667 B.n391 256.663
R1332 B.n667 B.n392 256.663
R1333 B.n667 B.n393 256.663
R1334 B.n667 B.n394 256.663
R1335 B.n667 B.n395 256.663
R1336 B.n667 B.n396 256.663
R1337 B.n667 B.n397 256.663
R1338 B.n667 B.n398 256.663
R1339 B.n667 B.n399 256.663
R1340 B.n667 B.n400 256.663
R1341 B.n667 B.n401 256.663
R1342 B.n667 B.n402 256.663
R1343 B.n667 B.n403 256.663
R1344 B.n667 B.n404 256.663
R1345 B.n667 B.n405 256.663
R1346 B.n667 B.n406 256.663
R1347 B.n667 B.n407 256.663
R1348 B.n667 B.n408 256.663
R1349 B.n667 B.n409 256.663
R1350 B.n667 B.n410 256.663
R1351 B.n667 B.n411 256.663
R1352 B.n667 B.n412 256.663
R1353 B.n667 B.n413 256.663
R1354 B.n667 B.n414 256.663
R1355 B.n667 B.n415 256.663
R1356 B.n667 B.n416 256.663
R1357 B.n667 B.n417 256.663
R1358 B.n667 B.n418 256.663
R1359 B.n667 B.n419 256.663
R1360 B.n667 B.n420 256.663
R1361 B.n667 B.n421 256.663
R1362 B.n667 B.n422 256.663
R1363 B.n667 B.n423 256.663
R1364 B.n667 B.n424 256.663
R1365 B.n667 B.n425 256.663
R1366 B.n667 B.n426 256.663
R1367 B.n667 B.n427 256.663
R1368 B.n667 B.n428 256.663
R1369 B.n667 B.n429 256.663
R1370 B.n667 B.n430 256.663
R1371 B.n667 B.n431 256.663
R1372 B.n667 B.n432 256.663
R1373 B.n667 B.n433 256.663
R1374 B.n667 B.n434 256.663
R1375 B.n667 B.n435 256.663
R1376 B.n667 B.n436 256.663
R1377 B.n667 B.n437 256.663
R1378 B.n667 B.n438 256.663
R1379 B.n667 B.n439 256.663
R1380 B.n667 B.n440 256.663
R1381 B.n667 B.n441 256.663
R1382 B.n667 B.n442 256.663
R1383 B.n667 B.n443 256.663
R1384 B.n674 B.n386 163.367
R1385 B.n674 B.n384 163.367
R1386 B.n678 B.n384 163.367
R1387 B.n678 B.n378 163.367
R1388 B.n686 B.n378 163.367
R1389 B.n686 B.n376 163.367
R1390 B.n690 B.n376 163.367
R1391 B.n690 B.n370 163.367
R1392 B.n698 B.n370 163.367
R1393 B.n698 B.n368 163.367
R1394 B.n702 B.n368 163.367
R1395 B.n702 B.n362 163.367
R1396 B.n711 B.n362 163.367
R1397 B.n711 B.n360 163.367
R1398 B.n715 B.n360 163.367
R1399 B.n715 B.n355 163.367
R1400 B.n723 B.n355 163.367
R1401 B.n723 B.n353 163.367
R1402 B.n727 B.n353 163.367
R1403 B.n727 B.n347 163.367
R1404 B.n735 B.n347 163.367
R1405 B.n735 B.n345 163.367
R1406 B.n739 B.n345 163.367
R1407 B.n739 B.n339 163.367
R1408 B.n748 B.n339 163.367
R1409 B.n748 B.n337 163.367
R1410 B.n752 B.n337 163.367
R1411 B.n752 B.n2 163.367
R1412 B.n856 B.n2 163.367
R1413 B.n856 B.n3 163.367
R1414 B.n852 B.n3 163.367
R1415 B.n852 B.n9 163.367
R1416 B.n848 B.n9 163.367
R1417 B.n848 B.n11 163.367
R1418 B.n844 B.n11 163.367
R1419 B.n844 B.n16 163.367
R1420 B.n840 B.n16 163.367
R1421 B.n840 B.n18 163.367
R1422 B.n836 B.n18 163.367
R1423 B.n836 B.n23 163.367
R1424 B.n832 B.n23 163.367
R1425 B.n832 B.n25 163.367
R1426 B.n828 B.n25 163.367
R1427 B.n828 B.n29 163.367
R1428 B.n824 B.n29 163.367
R1429 B.n824 B.n31 163.367
R1430 B.n820 B.n31 163.367
R1431 B.n820 B.n37 163.367
R1432 B.n816 B.n37 163.367
R1433 B.n816 B.n39 163.367
R1434 B.n812 B.n39 163.367
R1435 B.n812 B.n44 163.367
R1436 B.n808 B.n44 163.367
R1437 B.n808 B.n46 163.367
R1438 B.n804 B.n46 163.367
R1439 B.n804 B.n51 163.367
R1440 B.n800 B.n51 163.367
R1441 B.n800 B.n53 163.367
R1442 B.n445 B.n444 163.367
R1443 B.n660 B.n444 163.367
R1444 B.n658 B.n657 163.367
R1445 B.n654 B.n653 163.367
R1446 B.n650 B.n649 163.367
R1447 B.n646 B.n645 163.367
R1448 B.n642 B.n641 163.367
R1449 B.n638 B.n637 163.367
R1450 B.n634 B.n633 163.367
R1451 B.n630 B.n629 163.367
R1452 B.n626 B.n625 163.367
R1453 B.n622 B.n621 163.367
R1454 B.n618 B.n617 163.367
R1455 B.n614 B.n613 163.367
R1456 B.n610 B.n609 163.367
R1457 B.n606 B.n605 163.367
R1458 B.n602 B.n601 163.367
R1459 B.n598 B.n597 163.367
R1460 B.n594 B.n593 163.367
R1461 B.n590 B.n589 163.367
R1462 B.n586 B.n585 163.367
R1463 B.n582 B.n581 163.367
R1464 B.n578 B.n577 163.367
R1465 B.n574 B.n573 163.367
R1466 B.n570 B.n569 163.367
R1467 B.n565 B.n564 163.367
R1468 B.n561 B.n560 163.367
R1469 B.n557 B.n556 163.367
R1470 B.n553 B.n552 163.367
R1471 B.n549 B.n548 163.367
R1472 B.n544 B.n543 163.367
R1473 B.n540 B.n539 163.367
R1474 B.n536 B.n535 163.367
R1475 B.n532 B.n531 163.367
R1476 B.n528 B.n527 163.367
R1477 B.n524 B.n523 163.367
R1478 B.n520 B.n519 163.367
R1479 B.n516 B.n515 163.367
R1480 B.n512 B.n511 163.367
R1481 B.n508 B.n507 163.367
R1482 B.n504 B.n503 163.367
R1483 B.n500 B.n499 163.367
R1484 B.n496 B.n495 163.367
R1485 B.n492 B.n491 163.367
R1486 B.n488 B.n487 163.367
R1487 B.n484 B.n483 163.367
R1488 B.n480 B.n479 163.367
R1489 B.n476 B.n475 163.367
R1490 B.n472 B.n471 163.367
R1491 B.n468 B.n467 163.367
R1492 B.n464 B.n463 163.367
R1493 B.n460 B.n459 163.367
R1494 B.n456 B.n455 163.367
R1495 B.n452 B.n451 163.367
R1496 B.n668 B.n390 163.367
R1497 B.n672 B.n388 163.367
R1498 B.n672 B.n382 163.367
R1499 B.n680 B.n382 163.367
R1500 B.n680 B.n380 163.367
R1501 B.n684 B.n380 163.367
R1502 B.n684 B.n374 163.367
R1503 B.n692 B.n374 163.367
R1504 B.n692 B.n372 163.367
R1505 B.n696 B.n372 163.367
R1506 B.n696 B.n366 163.367
R1507 B.n704 B.n366 163.367
R1508 B.n704 B.n364 163.367
R1509 B.n708 B.n364 163.367
R1510 B.n708 B.n359 163.367
R1511 B.n717 B.n359 163.367
R1512 B.n717 B.n357 163.367
R1513 B.n721 B.n357 163.367
R1514 B.n721 B.n351 163.367
R1515 B.n729 B.n351 163.367
R1516 B.n729 B.n349 163.367
R1517 B.n733 B.n349 163.367
R1518 B.n733 B.n342 163.367
R1519 B.n741 B.n342 163.367
R1520 B.n741 B.n340 163.367
R1521 B.n746 B.n340 163.367
R1522 B.n746 B.n335 163.367
R1523 B.n754 B.n335 163.367
R1524 B.n755 B.n754 163.367
R1525 B.n755 B.n5 163.367
R1526 B.n6 B.n5 163.367
R1527 B.n7 B.n6 163.367
R1528 B.n760 B.n7 163.367
R1529 B.n760 B.n12 163.367
R1530 B.n13 B.n12 163.367
R1531 B.n14 B.n13 163.367
R1532 B.n765 B.n14 163.367
R1533 B.n765 B.n19 163.367
R1534 B.n20 B.n19 163.367
R1535 B.n21 B.n20 163.367
R1536 B.n770 B.n21 163.367
R1537 B.n770 B.n26 163.367
R1538 B.n27 B.n26 163.367
R1539 B.n28 B.n27 163.367
R1540 B.n775 B.n28 163.367
R1541 B.n775 B.n33 163.367
R1542 B.n34 B.n33 163.367
R1543 B.n35 B.n34 163.367
R1544 B.n780 B.n35 163.367
R1545 B.n780 B.n40 163.367
R1546 B.n41 B.n40 163.367
R1547 B.n42 B.n41 163.367
R1548 B.n785 B.n42 163.367
R1549 B.n785 B.n47 163.367
R1550 B.n48 B.n47 163.367
R1551 B.n49 B.n48 163.367
R1552 B.n790 B.n49 163.367
R1553 B.n790 B.n54 163.367
R1554 B.n55 B.n54 163.367
R1555 B.n121 B.n120 163.367
R1556 B.n125 B.n124 163.367
R1557 B.n129 B.n128 163.367
R1558 B.n133 B.n132 163.367
R1559 B.n137 B.n136 163.367
R1560 B.n141 B.n140 163.367
R1561 B.n145 B.n144 163.367
R1562 B.n149 B.n148 163.367
R1563 B.n153 B.n152 163.367
R1564 B.n157 B.n156 163.367
R1565 B.n161 B.n160 163.367
R1566 B.n165 B.n164 163.367
R1567 B.n169 B.n168 163.367
R1568 B.n173 B.n172 163.367
R1569 B.n177 B.n176 163.367
R1570 B.n181 B.n180 163.367
R1571 B.n185 B.n184 163.367
R1572 B.n189 B.n188 163.367
R1573 B.n193 B.n192 163.367
R1574 B.n197 B.n196 163.367
R1575 B.n201 B.n200 163.367
R1576 B.n205 B.n204 163.367
R1577 B.n209 B.n208 163.367
R1578 B.n213 B.n212 163.367
R1579 B.n217 B.n216 163.367
R1580 B.n221 B.n220 163.367
R1581 B.n225 B.n224 163.367
R1582 B.n229 B.n228 163.367
R1583 B.n233 B.n232 163.367
R1584 B.n237 B.n236 163.367
R1585 B.n241 B.n240 163.367
R1586 B.n245 B.n244 163.367
R1587 B.n249 B.n248 163.367
R1588 B.n253 B.n252 163.367
R1589 B.n257 B.n256 163.367
R1590 B.n261 B.n260 163.367
R1591 B.n265 B.n264 163.367
R1592 B.n269 B.n268 163.367
R1593 B.n273 B.n272 163.367
R1594 B.n277 B.n276 163.367
R1595 B.n281 B.n280 163.367
R1596 B.n285 B.n284 163.367
R1597 B.n289 B.n288 163.367
R1598 B.n293 B.n292 163.367
R1599 B.n297 B.n296 163.367
R1600 B.n301 B.n300 163.367
R1601 B.n305 B.n304 163.367
R1602 B.n309 B.n308 163.367
R1603 B.n313 B.n312 163.367
R1604 B.n317 B.n316 163.367
R1605 B.n321 B.n320 163.367
R1606 B.n325 B.n324 163.367
R1607 B.n329 B.n328 163.367
R1608 B.n331 B.n110 163.367
R1609 B.n666 B.n665 71.676
R1610 B.n660 B.n391 71.676
R1611 B.n657 B.n392 71.676
R1612 B.n653 B.n393 71.676
R1613 B.n649 B.n394 71.676
R1614 B.n645 B.n395 71.676
R1615 B.n641 B.n396 71.676
R1616 B.n637 B.n397 71.676
R1617 B.n633 B.n398 71.676
R1618 B.n629 B.n399 71.676
R1619 B.n625 B.n400 71.676
R1620 B.n621 B.n401 71.676
R1621 B.n617 B.n402 71.676
R1622 B.n613 B.n403 71.676
R1623 B.n609 B.n404 71.676
R1624 B.n605 B.n405 71.676
R1625 B.n601 B.n406 71.676
R1626 B.n597 B.n407 71.676
R1627 B.n593 B.n408 71.676
R1628 B.n589 B.n409 71.676
R1629 B.n585 B.n410 71.676
R1630 B.n581 B.n411 71.676
R1631 B.n577 B.n412 71.676
R1632 B.n573 B.n413 71.676
R1633 B.n569 B.n414 71.676
R1634 B.n564 B.n415 71.676
R1635 B.n560 B.n416 71.676
R1636 B.n556 B.n417 71.676
R1637 B.n552 B.n418 71.676
R1638 B.n548 B.n419 71.676
R1639 B.n543 B.n420 71.676
R1640 B.n539 B.n421 71.676
R1641 B.n535 B.n422 71.676
R1642 B.n531 B.n423 71.676
R1643 B.n527 B.n424 71.676
R1644 B.n523 B.n425 71.676
R1645 B.n519 B.n426 71.676
R1646 B.n515 B.n427 71.676
R1647 B.n511 B.n428 71.676
R1648 B.n507 B.n429 71.676
R1649 B.n503 B.n430 71.676
R1650 B.n499 B.n431 71.676
R1651 B.n495 B.n432 71.676
R1652 B.n491 B.n433 71.676
R1653 B.n487 B.n434 71.676
R1654 B.n483 B.n435 71.676
R1655 B.n479 B.n436 71.676
R1656 B.n475 B.n437 71.676
R1657 B.n471 B.n438 71.676
R1658 B.n467 B.n439 71.676
R1659 B.n463 B.n440 71.676
R1660 B.n459 B.n441 71.676
R1661 B.n455 B.n442 71.676
R1662 B.n451 B.n443 71.676
R1663 B.n117 B.n56 71.676
R1664 B.n121 B.n57 71.676
R1665 B.n125 B.n58 71.676
R1666 B.n129 B.n59 71.676
R1667 B.n133 B.n60 71.676
R1668 B.n137 B.n61 71.676
R1669 B.n141 B.n62 71.676
R1670 B.n145 B.n63 71.676
R1671 B.n149 B.n64 71.676
R1672 B.n153 B.n65 71.676
R1673 B.n157 B.n66 71.676
R1674 B.n161 B.n67 71.676
R1675 B.n165 B.n68 71.676
R1676 B.n169 B.n69 71.676
R1677 B.n173 B.n70 71.676
R1678 B.n177 B.n71 71.676
R1679 B.n181 B.n72 71.676
R1680 B.n185 B.n73 71.676
R1681 B.n189 B.n74 71.676
R1682 B.n193 B.n75 71.676
R1683 B.n197 B.n76 71.676
R1684 B.n201 B.n77 71.676
R1685 B.n205 B.n78 71.676
R1686 B.n209 B.n79 71.676
R1687 B.n213 B.n80 71.676
R1688 B.n217 B.n81 71.676
R1689 B.n221 B.n82 71.676
R1690 B.n225 B.n83 71.676
R1691 B.n229 B.n84 71.676
R1692 B.n233 B.n85 71.676
R1693 B.n237 B.n86 71.676
R1694 B.n241 B.n87 71.676
R1695 B.n245 B.n88 71.676
R1696 B.n249 B.n89 71.676
R1697 B.n253 B.n90 71.676
R1698 B.n257 B.n91 71.676
R1699 B.n261 B.n92 71.676
R1700 B.n265 B.n93 71.676
R1701 B.n269 B.n94 71.676
R1702 B.n273 B.n95 71.676
R1703 B.n277 B.n96 71.676
R1704 B.n281 B.n97 71.676
R1705 B.n285 B.n98 71.676
R1706 B.n289 B.n99 71.676
R1707 B.n293 B.n100 71.676
R1708 B.n297 B.n101 71.676
R1709 B.n301 B.n102 71.676
R1710 B.n305 B.n103 71.676
R1711 B.n309 B.n104 71.676
R1712 B.n313 B.n105 71.676
R1713 B.n317 B.n106 71.676
R1714 B.n321 B.n107 71.676
R1715 B.n325 B.n108 71.676
R1716 B.n329 B.n109 71.676
R1717 B.n796 B.n110 71.676
R1718 B.n796 B.n795 71.676
R1719 B.n331 B.n109 71.676
R1720 B.n328 B.n108 71.676
R1721 B.n324 B.n107 71.676
R1722 B.n320 B.n106 71.676
R1723 B.n316 B.n105 71.676
R1724 B.n312 B.n104 71.676
R1725 B.n308 B.n103 71.676
R1726 B.n304 B.n102 71.676
R1727 B.n300 B.n101 71.676
R1728 B.n296 B.n100 71.676
R1729 B.n292 B.n99 71.676
R1730 B.n288 B.n98 71.676
R1731 B.n284 B.n97 71.676
R1732 B.n280 B.n96 71.676
R1733 B.n276 B.n95 71.676
R1734 B.n272 B.n94 71.676
R1735 B.n268 B.n93 71.676
R1736 B.n264 B.n92 71.676
R1737 B.n260 B.n91 71.676
R1738 B.n256 B.n90 71.676
R1739 B.n252 B.n89 71.676
R1740 B.n248 B.n88 71.676
R1741 B.n244 B.n87 71.676
R1742 B.n240 B.n86 71.676
R1743 B.n236 B.n85 71.676
R1744 B.n232 B.n84 71.676
R1745 B.n228 B.n83 71.676
R1746 B.n224 B.n82 71.676
R1747 B.n220 B.n81 71.676
R1748 B.n216 B.n80 71.676
R1749 B.n212 B.n79 71.676
R1750 B.n208 B.n78 71.676
R1751 B.n204 B.n77 71.676
R1752 B.n200 B.n76 71.676
R1753 B.n196 B.n75 71.676
R1754 B.n192 B.n74 71.676
R1755 B.n188 B.n73 71.676
R1756 B.n184 B.n72 71.676
R1757 B.n180 B.n71 71.676
R1758 B.n176 B.n70 71.676
R1759 B.n172 B.n69 71.676
R1760 B.n168 B.n68 71.676
R1761 B.n164 B.n67 71.676
R1762 B.n160 B.n66 71.676
R1763 B.n156 B.n65 71.676
R1764 B.n152 B.n64 71.676
R1765 B.n148 B.n63 71.676
R1766 B.n144 B.n62 71.676
R1767 B.n140 B.n61 71.676
R1768 B.n136 B.n60 71.676
R1769 B.n132 B.n59 71.676
R1770 B.n128 B.n58 71.676
R1771 B.n124 B.n57 71.676
R1772 B.n120 B.n56 71.676
R1773 B.n666 B.n445 71.676
R1774 B.n658 B.n391 71.676
R1775 B.n654 B.n392 71.676
R1776 B.n650 B.n393 71.676
R1777 B.n646 B.n394 71.676
R1778 B.n642 B.n395 71.676
R1779 B.n638 B.n396 71.676
R1780 B.n634 B.n397 71.676
R1781 B.n630 B.n398 71.676
R1782 B.n626 B.n399 71.676
R1783 B.n622 B.n400 71.676
R1784 B.n618 B.n401 71.676
R1785 B.n614 B.n402 71.676
R1786 B.n610 B.n403 71.676
R1787 B.n606 B.n404 71.676
R1788 B.n602 B.n405 71.676
R1789 B.n598 B.n406 71.676
R1790 B.n594 B.n407 71.676
R1791 B.n590 B.n408 71.676
R1792 B.n586 B.n409 71.676
R1793 B.n582 B.n410 71.676
R1794 B.n578 B.n411 71.676
R1795 B.n574 B.n412 71.676
R1796 B.n570 B.n413 71.676
R1797 B.n565 B.n414 71.676
R1798 B.n561 B.n415 71.676
R1799 B.n557 B.n416 71.676
R1800 B.n553 B.n417 71.676
R1801 B.n549 B.n418 71.676
R1802 B.n544 B.n419 71.676
R1803 B.n540 B.n420 71.676
R1804 B.n536 B.n421 71.676
R1805 B.n532 B.n422 71.676
R1806 B.n528 B.n423 71.676
R1807 B.n524 B.n424 71.676
R1808 B.n520 B.n425 71.676
R1809 B.n516 B.n426 71.676
R1810 B.n512 B.n427 71.676
R1811 B.n508 B.n428 71.676
R1812 B.n504 B.n429 71.676
R1813 B.n500 B.n430 71.676
R1814 B.n496 B.n431 71.676
R1815 B.n492 B.n432 71.676
R1816 B.n488 B.n433 71.676
R1817 B.n484 B.n434 71.676
R1818 B.n480 B.n435 71.676
R1819 B.n476 B.n436 71.676
R1820 B.n472 B.n437 71.676
R1821 B.n468 B.n438 71.676
R1822 B.n464 B.n439 71.676
R1823 B.n460 B.n440 71.676
R1824 B.n456 B.n441 71.676
R1825 B.n452 B.n442 71.676
R1826 B.n443 B.n390 71.676
R1827 B.n667 B.n387 69.4166
R1828 B.n798 B.n797 69.4166
R1829 B.n546 B.n449 59.5399
R1830 B.n567 B.n447 59.5399
R1831 B.n116 B.n115 59.5399
R1832 B.n113 B.n112 59.5399
R1833 B.n673 B.n387 37.1682
R1834 B.n673 B.n383 37.1682
R1835 B.n679 B.n383 37.1682
R1836 B.n679 B.n379 37.1682
R1837 B.n685 B.n379 37.1682
R1838 B.n691 B.n375 37.1682
R1839 B.n691 B.n371 37.1682
R1840 B.n697 B.n371 37.1682
R1841 B.n697 B.n367 37.1682
R1842 B.n703 B.n367 37.1682
R1843 B.n703 B.n363 37.1682
R1844 B.n710 B.n363 37.1682
R1845 B.n710 B.n709 37.1682
R1846 B.n716 B.n356 37.1682
R1847 B.n722 B.n356 37.1682
R1848 B.n722 B.n352 37.1682
R1849 B.n728 B.n352 37.1682
R1850 B.n734 B.n348 37.1682
R1851 B.n734 B.n343 37.1682
R1852 B.n740 B.n343 37.1682
R1853 B.n740 B.n344 37.1682
R1854 B.n747 B.n336 37.1682
R1855 B.n753 B.n336 37.1682
R1856 B.n753 B.n4 37.1682
R1857 B.n855 B.n4 37.1682
R1858 B.n855 B.n854 37.1682
R1859 B.n854 B.n853 37.1682
R1860 B.n853 B.n8 37.1682
R1861 B.n847 B.n8 37.1682
R1862 B.n846 B.n845 37.1682
R1863 B.n845 B.n15 37.1682
R1864 B.n839 B.n15 37.1682
R1865 B.n839 B.n838 37.1682
R1866 B.n837 B.n22 37.1682
R1867 B.n831 B.n22 37.1682
R1868 B.n831 B.n830 37.1682
R1869 B.n830 B.n829 37.1682
R1870 B.n823 B.n32 37.1682
R1871 B.n823 B.n822 37.1682
R1872 B.n822 B.n821 37.1682
R1873 B.n821 B.n36 37.1682
R1874 B.n815 B.n36 37.1682
R1875 B.n815 B.n814 37.1682
R1876 B.n814 B.n813 37.1682
R1877 B.n813 B.n43 37.1682
R1878 B.n807 B.n806 37.1682
R1879 B.n806 B.n805 37.1682
R1880 B.n805 B.n50 37.1682
R1881 B.n799 B.n50 37.1682
R1882 B.n799 B.n798 37.1682
R1883 B.n449 B.n448 34.5217
R1884 B.n447 B.n446 34.5217
R1885 B.n115 B.n114 34.5217
R1886 B.n112 B.n111 34.5217
R1887 B.n685 B.t14 32.2489
R1888 B.n807 B.t7 32.2489
R1889 B.n794 B.n793 30.7517
R1890 B.n118 B.n52 30.7517
R1891 B.n670 B.n669 30.7517
R1892 B.n664 B.n385 30.7517
R1893 B.n344 B.t4 28.9694
R1894 B.t0 B.n846 28.9694
R1895 B.n716 B.t3 25.6899
R1896 B.n829 B.t2 25.6899
R1897 B.n728 B.t1 20.2241
R1898 B.t5 B.n837 20.2241
R1899 B B.n857 18.0485
R1900 B.t1 B.n348 16.9446
R1901 B.n838 B.t5 16.9446
R1902 B.n709 B.t3 11.4788
R1903 B.n32 B.t2 11.4788
R1904 B.n119 B.n118 10.6151
R1905 B.n122 B.n119 10.6151
R1906 B.n123 B.n122 10.6151
R1907 B.n126 B.n123 10.6151
R1908 B.n127 B.n126 10.6151
R1909 B.n130 B.n127 10.6151
R1910 B.n131 B.n130 10.6151
R1911 B.n134 B.n131 10.6151
R1912 B.n135 B.n134 10.6151
R1913 B.n138 B.n135 10.6151
R1914 B.n139 B.n138 10.6151
R1915 B.n142 B.n139 10.6151
R1916 B.n143 B.n142 10.6151
R1917 B.n146 B.n143 10.6151
R1918 B.n147 B.n146 10.6151
R1919 B.n150 B.n147 10.6151
R1920 B.n151 B.n150 10.6151
R1921 B.n154 B.n151 10.6151
R1922 B.n155 B.n154 10.6151
R1923 B.n158 B.n155 10.6151
R1924 B.n159 B.n158 10.6151
R1925 B.n162 B.n159 10.6151
R1926 B.n163 B.n162 10.6151
R1927 B.n166 B.n163 10.6151
R1928 B.n167 B.n166 10.6151
R1929 B.n170 B.n167 10.6151
R1930 B.n171 B.n170 10.6151
R1931 B.n174 B.n171 10.6151
R1932 B.n175 B.n174 10.6151
R1933 B.n178 B.n175 10.6151
R1934 B.n179 B.n178 10.6151
R1935 B.n182 B.n179 10.6151
R1936 B.n183 B.n182 10.6151
R1937 B.n186 B.n183 10.6151
R1938 B.n187 B.n186 10.6151
R1939 B.n190 B.n187 10.6151
R1940 B.n191 B.n190 10.6151
R1941 B.n194 B.n191 10.6151
R1942 B.n195 B.n194 10.6151
R1943 B.n198 B.n195 10.6151
R1944 B.n199 B.n198 10.6151
R1945 B.n202 B.n199 10.6151
R1946 B.n203 B.n202 10.6151
R1947 B.n206 B.n203 10.6151
R1948 B.n207 B.n206 10.6151
R1949 B.n210 B.n207 10.6151
R1950 B.n211 B.n210 10.6151
R1951 B.n214 B.n211 10.6151
R1952 B.n215 B.n214 10.6151
R1953 B.n219 B.n218 10.6151
R1954 B.n222 B.n219 10.6151
R1955 B.n223 B.n222 10.6151
R1956 B.n226 B.n223 10.6151
R1957 B.n227 B.n226 10.6151
R1958 B.n230 B.n227 10.6151
R1959 B.n231 B.n230 10.6151
R1960 B.n234 B.n231 10.6151
R1961 B.n235 B.n234 10.6151
R1962 B.n239 B.n238 10.6151
R1963 B.n242 B.n239 10.6151
R1964 B.n243 B.n242 10.6151
R1965 B.n246 B.n243 10.6151
R1966 B.n247 B.n246 10.6151
R1967 B.n250 B.n247 10.6151
R1968 B.n251 B.n250 10.6151
R1969 B.n254 B.n251 10.6151
R1970 B.n255 B.n254 10.6151
R1971 B.n258 B.n255 10.6151
R1972 B.n259 B.n258 10.6151
R1973 B.n262 B.n259 10.6151
R1974 B.n263 B.n262 10.6151
R1975 B.n266 B.n263 10.6151
R1976 B.n267 B.n266 10.6151
R1977 B.n270 B.n267 10.6151
R1978 B.n271 B.n270 10.6151
R1979 B.n274 B.n271 10.6151
R1980 B.n275 B.n274 10.6151
R1981 B.n278 B.n275 10.6151
R1982 B.n279 B.n278 10.6151
R1983 B.n282 B.n279 10.6151
R1984 B.n283 B.n282 10.6151
R1985 B.n286 B.n283 10.6151
R1986 B.n287 B.n286 10.6151
R1987 B.n290 B.n287 10.6151
R1988 B.n291 B.n290 10.6151
R1989 B.n294 B.n291 10.6151
R1990 B.n295 B.n294 10.6151
R1991 B.n298 B.n295 10.6151
R1992 B.n299 B.n298 10.6151
R1993 B.n302 B.n299 10.6151
R1994 B.n303 B.n302 10.6151
R1995 B.n306 B.n303 10.6151
R1996 B.n307 B.n306 10.6151
R1997 B.n310 B.n307 10.6151
R1998 B.n311 B.n310 10.6151
R1999 B.n314 B.n311 10.6151
R2000 B.n315 B.n314 10.6151
R2001 B.n318 B.n315 10.6151
R2002 B.n319 B.n318 10.6151
R2003 B.n322 B.n319 10.6151
R2004 B.n323 B.n322 10.6151
R2005 B.n326 B.n323 10.6151
R2006 B.n327 B.n326 10.6151
R2007 B.n330 B.n327 10.6151
R2008 B.n332 B.n330 10.6151
R2009 B.n333 B.n332 10.6151
R2010 B.n794 B.n333 10.6151
R2011 B.n671 B.n670 10.6151
R2012 B.n671 B.n381 10.6151
R2013 B.n681 B.n381 10.6151
R2014 B.n682 B.n681 10.6151
R2015 B.n683 B.n682 10.6151
R2016 B.n683 B.n373 10.6151
R2017 B.n693 B.n373 10.6151
R2018 B.n694 B.n693 10.6151
R2019 B.n695 B.n694 10.6151
R2020 B.n695 B.n365 10.6151
R2021 B.n705 B.n365 10.6151
R2022 B.n706 B.n705 10.6151
R2023 B.n707 B.n706 10.6151
R2024 B.n707 B.n358 10.6151
R2025 B.n718 B.n358 10.6151
R2026 B.n719 B.n718 10.6151
R2027 B.n720 B.n719 10.6151
R2028 B.n720 B.n350 10.6151
R2029 B.n730 B.n350 10.6151
R2030 B.n731 B.n730 10.6151
R2031 B.n732 B.n731 10.6151
R2032 B.n732 B.n341 10.6151
R2033 B.n742 B.n341 10.6151
R2034 B.n743 B.n742 10.6151
R2035 B.n745 B.n743 10.6151
R2036 B.n745 B.n744 10.6151
R2037 B.n744 B.n334 10.6151
R2038 B.n756 B.n334 10.6151
R2039 B.n757 B.n756 10.6151
R2040 B.n758 B.n757 10.6151
R2041 B.n759 B.n758 10.6151
R2042 B.n761 B.n759 10.6151
R2043 B.n762 B.n761 10.6151
R2044 B.n763 B.n762 10.6151
R2045 B.n764 B.n763 10.6151
R2046 B.n766 B.n764 10.6151
R2047 B.n767 B.n766 10.6151
R2048 B.n768 B.n767 10.6151
R2049 B.n769 B.n768 10.6151
R2050 B.n771 B.n769 10.6151
R2051 B.n772 B.n771 10.6151
R2052 B.n773 B.n772 10.6151
R2053 B.n774 B.n773 10.6151
R2054 B.n776 B.n774 10.6151
R2055 B.n777 B.n776 10.6151
R2056 B.n778 B.n777 10.6151
R2057 B.n779 B.n778 10.6151
R2058 B.n781 B.n779 10.6151
R2059 B.n782 B.n781 10.6151
R2060 B.n783 B.n782 10.6151
R2061 B.n784 B.n783 10.6151
R2062 B.n786 B.n784 10.6151
R2063 B.n787 B.n786 10.6151
R2064 B.n788 B.n787 10.6151
R2065 B.n789 B.n788 10.6151
R2066 B.n791 B.n789 10.6151
R2067 B.n792 B.n791 10.6151
R2068 B.n793 B.n792 10.6151
R2069 B.n664 B.n663 10.6151
R2070 B.n663 B.n662 10.6151
R2071 B.n662 B.n661 10.6151
R2072 B.n661 B.n659 10.6151
R2073 B.n659 B.n656 10.6151
R2074 B.n656 B.n655 10.6151
R2075 B.n655 B.n652 10.6151
R2076 B.n652 B.n651 10.6151
R2077 B.n651 B.n648 10.6151
R2078 B.n648 B.n647 10.6151
R2079 B.n647 B.n644 10.6151
R2080 B.n644 B.n643 10.6151
R2081 B.n643 B.n640 10.6151
R2082 B.n640 B.n639 10.6151
R2083 B.n639 B.n636 10.6151
R2084 B.n636 B.n635 10.6151
R2085 B.n635 B.n632 10.6151
R2086 B.n632 B.n631 10.6151
R2087 B.n631 B.n628 10.6151
R2088 B.n628 B.n627 10.6151
R2089 B.n627 B.n624 10.6151
R2090 B.n624 B.n623 10.6151
R2091 B.n623 B.n620 10.6151
R2092 B.n620 B.n619 10.6151
R2093 B.n619 B.n616 10.6151
R2094 B.n616 B.n615 10.6151
R2095 B.n615 B.n612 10.6151
R2096 B.n612 B.n611 10.6151
R2097 B.n611 B.n608 10.6151
R2098 B.n608 B.n607 10.6151
R2099 B.n607 B.n604 10.6151
R2100 B.n604 B.n603 10.6151
R2101 B.n603 B.n600 10.6151
R2102 B.n600 B.n599 10.6151
R2103 B.n599 B.n596 10.6151
R2104 B.n596 B.n595 10.6151
R2105 B.n595 B.n592 10.6151
R2106 B.n592 B.n591 10.6151
R2107 B.n591 B.n588 10.6151
R2108 B.n588 B.n587 10.6151
R2109 B.n587 B.n584 10.6151
R2110 B.n584 B.n583 10.6151
R2111 B.n583 B.n580 10.6151
R2112 B.n580 B.n579 10.6151
R2113 B.n579 B.n576 10.6151
R2114 B.n576 B.n575 10.6151
R2115 B.n575 B.n572 10.6151
R2116 B.n572 B.n571 10.6151
R2117 B.n571 B.n568 10.6151
R2118 B.n566 B.n563 10.6151
R2119 B.n563 B.n562 10.6151
R2120 B.n562 B.n559 10.6151
R2121 B.n559 B.n558 10.6151
R2122 B.n558 B.n555 10.6151
R2123 B.n555 B.n554 10.6151
R2124 B.n554 B.n551 10.6151
R2125 B.n551 B.n550 10.6151
R2126 B.n550 B.n547 10.6151
R2127 B.n545 B.n542 10.6151
R2128 B.n542 B.n541 10.6151
R2129 B.n541 B.n538 10.6151
R2130 B.n538 B.n537 10.6151
R2131 B.n537 B.n534 10.6151
R2132 B.n534 B.n533 10.6151
R2133 B.n533 B.n530 10.6151
R2134 B.n530 B.n529 10.6151
R2135 B.n529 B.n526 10.6151
R2136 B.n526 B.n525 10.6151
R2137 B.n525 B.n522 10.6151
R2138 B.n522 B.n521 10.6151
R2139 B.n521 B.n518 10.6151
R2140 B.n518 B.n517 10.6151
R2141 B.n517 B.n514 10.6151
R2142 B.n514 B.n513 10.6151
R2143 B.n513 B.n510 10.6151
R2144 B.n510 B.n509 10.6151
R2145 B.n509 B.n506 10.6151
R2146 B.n506 B.n505 10.6151
R2147 B.n505 B.n502 10.6151
R2148 B.n502 B.n501 10.6151
R2149 B.n501 B.n498 10.6151
R2150 B.n498 B.n497 10.6151
R2151 B.n497 B.n494 10.6151
R2152 B.n494 B.n493 10.6151
R2153 B.n493 B.n490 10.6151
R2154 B.n490 B.n489 10.6151
R2155 B.n489 B.n486 10.6151
R2156 B.n486 B.n485 10.6151
R2157 B.n485 B.n482 10.6151
R2158 B.n482 B.n481 10.6151
R2159 B.n481 B.n478 10.6151
R2160 B.n478 B.n477 10.6151
R2161 B.n477 B.n474 10.6151
R2162 B.n474 B.n473 10.6151
R2163 B.n473 B.n470 10.6151
R2164 B.n470 B.n469 10.6151
R2165 B.n469 B.n466 10.6151
R2166 B.n466 B.n465 10.6151
R2167 B.n465 B.n462 10.6151
R2168 B.n462 B.n461 10.6151
R2169 B.n461 B.n458 10.6151
R2170 B.n458 B.n457 10.6151
R2171 B.n457 B.n454 10.6151
R2172 B.n454 B.n453 10.6151
R2173 B.n453 B.n450 10.6151
R2174 B.n450 B.n389 10.6151
R2175 B.n669 B.n389 10.6151
R2176 B.n675 B.n385 10.6151
R2177 B.n676 B.n675 10.6151
R2178 B.n677 B.n676 10.6151
R2179 B.n677 B.n377 10.6151
R2180 B.n687 B.n377 10.6151
R2181 B.n688 B.n687 10.6151
R2182 B.n689 B.n688 10.6151
R2183 B.n689 B.n369 10.6151
R2184 B.n699 B.n369 10.6151
R2185 B.n700 B.n699 10.6151
R2186 B.n701 B.n700 10.6151
R2187 B.n701 B.n361 10.6151
R2188 B.n712 B.n361 10.6151
R2189 B.n713 B.n712 10.6151
R2190 B.n714 B.n713 10.6151
R2191 B.n714 B.n354 10.6151
R2192 B.n724 B.n354 10.6151
R2193 B.n725 B.n724 10.6151
R2194 B.n726 B.n725 10.6151
R2195 B.n726 B.n346 10.6151
R2196 B.n736 B.n346 10.6151
R2197 B.n737 B.n736 10.6151
R2198 B.n738 B.n737 10.6151
R2199 B.n738 B.n338 10.6151
R2200 B.n749 B.n338 10.6151
R2201 B.n750 B.n749 10.6151
R2202 B.n751 B.n750 10.6151
R2203 B.n751 B.n0 10.6151
R2204 B.n851 B.n1 10.6151
R2205 B.n851 B.n850 10.6151
R2206 B.n850 B.n849 10.6151
R2207 B.n849 B.n10 10.6151
R2208 B.n843 B.n10 10.6151
R2209 B.n843 B.n842 10.6151
R2210 B.n842 B.n841 10.6151
R2211 B.n841 B.n17 10.6151
R2212 B.n835 B.n17 10.6151
R2213 B.n835 B.n834 10.6151
R2214 B.n834 B.n833 10.6151
R2215 B.n833 B.n24 10.6151
R2216 B.n827 B.n24 10.6151
R2217 B.n827 B.n826 10.6151
R2218 B.n826 B.n825 10.6151
R2219 B.n825 B.n30 10.6151
R2220 B.n819 B.n30 10.6151
R2221 B.n819 B.n818 10.6151
R2222 B.n818 B.n817 10.6151
R2223 B.n817 B.n38 10.6151
R2224 B.n811 B.n38 10.6151
R2225 B.n811 B.n810 10.6151
R2226 B.n810 B.n809 10.6151
R2227 B.n809 B.n45 10.6151
R2228 B.n803 B.n45 10.6151
R2229 B.n803 B.n802 10.6151
R2230 B.n802 B.n801 10.6151
R2231 B.n801 B.n52 10.6151
R2232 B.n215 B.n116 9.36635
R2233 B.n238 B.n113 9.36635
R2234 B.n568 B.n567 9.36635
R2235 B.n546 B.n545 9.36635
R2236 B.n747 B.t4 8.19926
R2237 B.n847 B.t0 8.19926
R2238 B.t14 B.n375 4.91975
R2239 B.t7 B.n43 4.91975
R2240 B.n857 B.n0 2.81026
R2241 B.n857 B.n1 2.81026
R2242 B.n218 B.n116 1.24928
R2243 B.n235 B.n113 1.24928
R2244 B.n567 B.n566 1.24928
R2245 B.n547 B.n546 1.24928
R2246 VP.n7 VP.t4 283.149
R2247 VP.n20 VP.t1 246.817
R2248 VP.n14 VP.t0 246.817
R2249 VP.n26 VP.t5 246.817
R2250 VP.n6 VP.t2 246.817
R2251 VP.n12 VP.t3 246.817
R2252 VP.n15 VP.n14 172.065
R2253 VP.n27 VP.n26 172.065
R2254 VP.n13 VP.n12 172.065
R2255 VP.n8 VP.n5 161.3
R2256 VP.n10 VP.n9 161.3
R2257 VP.n11 VP.n4 161.3
R2258 VP.n25 VP.n0 161.3
R2259 VP.n24 VP.n23 161.3
R2260 VP.n22 VP.n1 161.3
R2261 VP.n21 VP.n20 161.3
R2262 VP.n19 VP.n2 161.3
R2263 VP.n18 VP.n17 161.3
R2264 VP.n16 VP.n3 161.3
R2265 VP.n19 VP.n18 51.1773
R2266 VP.n24 VP.n1 51.1773
R2267 VP.n10 VP.n5 51.1773
R2268 VP.n15 VP.n13 46.296
R2269 VP.n7 VP.n6 41.8525
R2270 VP.n18 VP.n3 29.8095
R2271 VP.n25 VP.n24 29.8095
R2272 VP.n11 VP.n10 29.8095
R2273 VP.n20 VP.n19 24.4675
R2274 VP.n20 VP.n1 24.4675
R2275 VP.n6 VP.n5 24.4675
R2276 VP.n8 VP.n7 17.3787
R2277 VP.n14 VP.n3 13.702
R2278 VP.n26 VP.n25 13.702
R2279 VP.n12 VP.n11 13.702
R2280 VP.n9 VP.n8 0.189894
R2281 VP.n9 VP.n4 0.189894
R2282 VP.n13 VP.n4 0.189894
R2283 VP.n16 VP.n15 0.189894
R2284 VP.n17 VP.n16 0.189894
R2285 VP.n17 VP.n2 0.189894
R2286 VP.n21 VP.n2 0.189894
R2287 VP.n22 VP.n21 0.189894
R2288 VP.n23 VP.n22 0.189894
R2289 VP.n23 VP.n0 0.189894
R2290 VP.n27 VP.n0 0.189894
R2291 VP VP.n27 0.0516364
R2292 VDD1.n76 VDD1.n0 289.615
R2293 VDD1.n157 VDD1.n81 289.615
R2294 VDD1.n77 VDD1.n76 185
R2295 VDD1.n75 VDD1.n74 185
R2296 VDD1.n73 VDD1.n3 185
R2297 VDD1.n7 VDD1.n4 185
R2298 VDD1.n68 VDD1.n67 185
R2299 VDD1.n66 VDD1.n65 185
R2300 VDD1.n9 VDD1.n8 185
R2301 VDD1.n60 VDD1.n59 185
R2302 VDD1.n58 VDD1.n57 185
R2303 VDD1.n13 VDD1.n12 185
R2304 VDD1.n52 VDD1.n51 185
R2305 VDD1.n50 VDD1.n49 185
R2306 VDD1.n17 VDD1.n16 185
R2307 VDD1.n44 VDD1.n43 185
R2308 VDD1.n42 VDD1.n41 185
R2309 VDD1.n21 VDD1.n20 185
R2310 VDD1.n36 VDD1.n35 185
R2311 VDD1.n34 VDD1.n33 185
R2312 VDD1.n25 VDD1.n24 185
R2313 VDD1.n28 VDD1.n27 185
R2314 VDD1.n108 VDD1.n107 185
R2315 VDD1.n105 VDD1.n104 185
R2316 VDD1.n114 VDD1.n113 185
R2317 VDD1.n116 VDD1.n115 185
R2318 VDD1.n101 VDD1.n100 185
R2319 VDD1.n122 VDD1.n121 185
R2320 VDD1.n124 VDD1.n123 185
R2321 VDD1.n97 VDD1.n96 185
R2322 VDD1.n130 VDD1.n129 185
R2323 VDD1.n132 VDD1.n131 185
R2324 VDD1.n93 VDD1.n92 185
R2325 VDD1.n138 VDD1.n137 185
R2326 VDD1.n140 VDD1.n139 185
R2327 VDD1.n89 VDD1.n88 185
R2328 VDD1.n146 VDD1.n145 185
R2329 VDD1.n149 VDD1.n148 185
R2330 VDD1.n147 VDD1.n85 185
R2331 VDD1.n154 VDD1.n84 185
R2332 VDD1.n156 VDD1.n155 185
R2333 VDD1.n158 VDD1.n157 185
R2334 VDD1.t1 VDD1.n26 147.659
R2335 VDD1.t5 VDD1.n106 147.659
R2336 VDD1.n76 VDD1.n75 104.615
R2337 VDD1.n75 VDD1.n3 104.615
R2338 VDD1.n7 VDD1.n3 104.615
R2339 VDD1.n67 VDD1.n7 104.615
R2340 VDD1.n67 VDD1.n66 104.615
R2341 VDD1.n66 VDD1.n8 104.615
R2342 VDD1.n59 VDD1.n8 104.615
R2343 VDD1.n59 VDD1.n58 104.615
R2344 VDD1.n58 VDD1.n12 104.615
R2345 VDD1.n51 VDD1.n12 104.615
R2346 VDD1.n51 VDD1.n50 104.615
R2347 VDD1.n50 VDD1.n16 104.615
R2348 VDD1.n43 VDD1.n16 104.615
R2349 VDD1.n43 VDD1.n42 104.615
R2350 VDD1.n42 VDD1.n20 104.615
R2351 VDD1.n35 VDD1.n20 104.615
R2352 VDD1.n35 VDD1.n34 104.615
R2353 VDD1.n34 VDD1.n24 104.615
R2354 VDD1.n27 VDD1.n24 104.615
R2355 VDD1.n107 VDD1.n104 104.615
R2356 VDD1.n114 VDD1.n104 104.615
R2357 VDD1.n115 VDD1.n114 104.615
R2358 VDD1.n115 VDD1.n100 104.615
R2359 VDD1.n122 VDD1.n100 104.615
R2360 VDD1.n123 VDD1.n122 104.615
R2361 VDD1.n123 VDD1.n96 104.615
R2362 VDD1.n130 VDD1.n96 104.615
R2363 VDD1.n131 VDD1.n130 104.615
R2364 VDD1.n131 VDD1.n92 104.615
R2365 VDD1.n138 VDD1.n92 104.615
R2366 VDD1.n139 VDD1.n138 104.615
R2367 VDD1.n139 VDD1.n88 104.615
R2368 VDD1.n146 VDD1.n88 104.615
R2369 VDD1.n148 VDD1.n146 104.615
R2370 VDD1.n148 VDD1.n147 104.615
R2371 VDD1.n147 VDD1.n84 104.615
R2372 VDD1.n156 VDD1.n84 104.615
R2373 VDD1.n157 VDD1.n156 104.615
R2374 VDD1.n163 VDD1.n162 65.3219
R2375 VDD1.n165 VDD1.n164 64.9936
R2376 VDD1 VDD1.n80 54.1459
R2377 VDD1.n163 VDD1.n161 54.0324
R2378 VDD1.n27 VDD1.t1 52.3082
R2379 VDD1.n107 VDD1.t5 52.3082
R2380 VDD1.n165 VDD1.n163 42.8543
R2381 VDD1.n28 VDD1.n26 15.6677
R2382 VDD1.n108 VDD1.n106 15.6677
R2383 VDD1.n74 VDD1.n73 13.1884
R2384 VDD1.n155 VDD1.n154 13.1884
R2385 VDD1.n77 VDD1.n2 12.8005
R2386 VDD1.n72 VDD1.n4 12.8005
R2387 VDD1.n29 VDD1.n25 12.8005
R2388 VDD1.n109 VDD1.n105 12.8005
R2389 VDD1.n153 VDD1.n85 12.8005
R2390 VDD1.n158 VDD1.n83 12.8005
R2391 VDD1.n78 VDD1.n0 12.0247
R2392 VDD1.n69 VDD1.n68 12.0247
R2393 VDD1.n33 VDD1.n32 12.0247
R2394 VDD1.n113 VDD1.n112 12.0247
R2395 VDD1.n150 VDD1.n149 12.0247
R2396 VDD1.n159 VDD1.n81 12.0247
R2397 VDD1.n65 VDD1.n6 11.249
R2398 VDD1.n36 VDD1.n23 11.249
R2399 VDD1.n116 VDD1.n103 11.249
R2400 VDD1.n145 VDD1.n87 11.249
R2401 VDD1.n64 VDD1.n9 10.4732
R2402 VDD1.n37 VDD1.n21 10.4732
R2403 VDD1.n117 VDD1.n101 10.4732
R2404 VDD1.n144 VDD1.n89 10.4732
R2405 VDD1.n61 VDD1.n60 9.69747
R2406 VDD1.n41 VDD1.n40 9.69747
R2407 VDD1.n121 VDD1.n120 9.69747
R2408 VDD1.n141 VDD1.n140 9.69747
R2409 VDD1.n80 VDD1.n79 9.45567
R2410 VDD1.n161 VDD1.n160 9.45567
R2411 VDD1.n54 VDD1.n53 9.3005
R2412 VDD1.n56 VDD1.n55 9.3005
R2413 VDD1.n11 VDD1.n10 9.3005
R2414 VDD1.n62 VDD1.n61 9.3005
R2415 VDD1.n64 VDD1.n63 9.3005
R2416 VDD1.n6 VDD1.n5 9.3005
R2417 VDD1.n70 VDD1.n69 9.3005
R2418 VDD1.n72 VDD1.n71 9.3005
R2419 VDD1.n79 VDD1.n78 9.3005
R2420 VDD1.n2 VDD1.n1 9.3005
R2421 VDD1.n15 VDD1.n14 9.3005
R2422 VDD1.n48 VDD1.n47 9.3005
R2423 VDD1.n46 VDD1.n45 9.3005
R2424 VDD1.n19 VDD1.n18 9.3005
R2425 VDD1.n40 VDD1.n39 9.3005
R2426 VDD1.n38 VDD1.n37 9.3005
R2427 VDD1.n23 VDD1.n22 9.3005
R2428 VDD1.n32 VDD1.n31 9.3005
R2429 VDD1.n30 VDD1.n29 9.3005
R2430 VDD1.n160 VDD1.n159 9.3005
R2431 VDD1.n83 VDD1.n82 9.3005
R2432 VDD1.n128 VDD1.n127 9.3005
R2433 VDD1.n126 VDD1.n125 9.3005
R2434 VDD1.n99 VDD1.n98 9.3005
R2435 VDD1.n120 VDD1.n119 9.3005
R2436 VDD1.n118 VDD1.n117 9.3005
R2437 VDD1.n103 VDD1.n102 9.3005
R2438 VDD1.n112 VDD1.n111 9.3005
R2439 VDD1.n110 VDD1.n109 9.3005
R2440 VDD1.n95 VDD1.n94 9.3005
R2441 VDD1.n134 VDD1.n133 9.3005
R2442 VDD1.n136 VDD1.n135 9.3005
R2443 VDD1.n91 VDD1.n90 9.3005
R2444 VDD1.n142 VDD1.n141 9.3005
R2445 VDD1.n144 VDD1.n143 9.3005
R2446 VDD1.n87 VDD1.n86 9.3005
R2447 VDD1.n151 VDD1.n150 9.3005
R2448 VDD1.n153 VDD1.n152 9.3005
R2449 VDD1.n57 VDD1.n11 8.92171
R2450 VDD1.n44 VDD1.n19 8.92171
R2451 VDD1.n124 VDD1.n99 8.92171
R2452 VDD1.n137 VDD1.n91 8.92171
R2453 VDD1.n56 VDD1.n13 8.14595
R2454 VDD1.n45 VDD1.n17 8.14595
R2455 VDD1.n125 VDD1.n97 8.14595
R2456 VDD1.n136 VDD1.n93 8.14595
R2457 VDD1.n53 VDD1.n52 7.3702
R2458 VDD1.n49 VDD1.n48 7.3702
R2459 VDD1.n129 VDD1.n128 7.3702
R2460 VDD1.n133 VDD1.n132 7.3702
R2461 VDD1.n52 VDD1.n15 6.59444
R2462 VDD1.n49 VDD1.n15 6.59444
R2463 VDD1.n129 VDD1.n95 6.59444
R2464 VDD1.n132 VDD1.n95 6.59444
R2465 VDD1.n53 VDD1.n13 5.81868
R2466 VDD1.n48 VDD1.n17 5.81868
R2467 VDD1.n128 VDD1.n97 5.81868
R2468 VDD1.n133 VDD1.n93 5.81868
R2469 VDD1.n57 VDD1.n56 5.04292
R2470 VDD1.n45 VDD1.n44 5.04292
R2471 VDD1.n125 VDD1.n124 5.04292
R2472 VDD1.n137 VDD1.n136 5.04292
R2473 VDD1.n30 VDD1.n26 4.38563
R2474 VDD1.n110 VDD1.n106 4.38563
R2475 VDD1.n60 VDD1.n11 4.26717
R2476 VDD1.n41 VDD1.n19 4.26717
R2477 VDD1.n121 VDD1.n99 4.26717
R2478 VDD1.n140 VDD1.n91 4.26717
R2479 VDD1.n61 VDD1.n9 3.49141
R2480 VDD1.n40 VDD1.n21 3.49141
R2481 VDD1.n120 VDD1.n101 3.49141
R2482 VDD1.n141 VDD1.n89 3.49141
R2483 VDD1.n65 VDD1.n64 2.71565
R2484 VDD1.n37 VDD1.n36 2.71565
R2485 VDD1.n117 VDD1.n116 2.71565
R2486 VDD1.n145 VDD1.n144 2.71565
R2487 VDD1.n80 VDD1.n0 1.93989
R2488 VDD1.n68 VDD1.n6 1.93989
R2489 VDD1.n33 VDD1.n23 1.93989
R2490 VDD1.n113 VDD1.n103 1.93989
R2491 VDD1.n149 VDD1.n87 1.93989
R2492 VDD1.n161 VDD1.n81 1.93989
R2493 VDD1.n164 VDD1.t3 1.33383
R2494 VDD1.n164 VDD1.t2 1.33383
R2495 VDD1.n162 VDD1.t4 1.33383
R2496 VDD1.n162 VDD1.t0 1.33383
R2497 VDD1.n78 VDD1.n77 1.16414
R2498 VDD1.n69 VDD1.n4 1.16414
R2499 VDD1.n32 VDD1.n25 1.16414
R2500 VDD1.n112 VDD1.n105 1.16414
R2501 VDD1.n150 VDD1.n85 1.16414
R2502 VDD1.n159 VDD1.n158 1.16414
R2503 VDD1.n74 VDD1.n2 0.388379
R2504 VDD1.n73 VDD1.n72 0.388379
R2505 VDD1.n29 VDD1.n28 0.388379
R2506 VDD1.n109 VDD1.n108 0.388379
R2507 VDD1.n154 VDD1.n153 0.388379
R2508 VDD1.n155 VDD1.n83 0.388379
R2509 VDD1 VDD1.n165 0.325931
R2510 VDD1.n79 VDD1.n1 0.155672
R2511 VDD1.n71 VDD1.n1 0.155672
R2512 VDD1.n71 VDD1.n70 0.155672
R2513 VDD1.n70 VDD1.n5 0.155672
R2514 VDD1.n63 VDD1.n5 0.155672
R2515 VDD1.n63 VDD1.n62 0.155672
R2516 VDD1.n62 VDD1.n10 0.155672
R2517 VDD1.n55 VDD1.n10 0.155672
R2518 VDD1.n55 VDD1.n54 0.155672
R2519 VDD1.n54 VDD1.n14 0.155672
R2520 VDD1.n47 VDD1.n14 0.155672
R2521 VDD1.n47 VDD1.n46 0.155672
R2522 VDD1.n46 VDD1.n18 0.155672
R2523 VDD1.n39 VDD1.n18 0.155672
R2524 VDD1.n39 VDD1.n38 0.155672
R2525 VDD1.n38 VDD1.n22 0.155672
R2526 VDD1.n31 VDD1.n22 0.155672
R2527 VDD1.n31 VDD1.n30 0.155672
R2528 VDD1.n111 VDD1.n110 0.155672
R2529 VDD1.n111 VDD1.n102 0.155672
R2530 VDD1.n118 VDD1.n102 0.155672
R2531 VDD1.n119 VDD1.n118 0.155672
R2532 VDD1.n119 VDD1.n98 0.155672
R2533 VDD1.n126 VDD1.n98 0.155672
R2534 VDD1.n127 VDD1.n126 0.155672
R2535 VDD1.n127 VDD1.n94 0.155672
R2536 VDD1.n134 VDD1.n94 0.155672
R2537 VDD1.n135 VDD1.n134 0.155672
R2538 VDD1.n135 VDD1.n90 0.155672
R2539 VDD1.n142 VDD1.n90 0.155672
R2540 VDD1.n143 VDD1.n142 0.155672
R2541 VDD1.n143 VDD1.n86 0.155672
R2542 VDD1.n151 VDD1.n86 0.155672
R2543 VDD1.n152 VDD1.n151 0.155672
R2544 VDD1.n152 VDD1.n82 0.155672
R2545 VDD1.n160 VDD1.n82 0.155672
C0 VDD2 VP 0.361243f
C1 VTAIL VDD1 9.367781f
C2 VDD2 VN 7.11328f
C3 VDD2 VTAIL 9.408031f
C4 VP VN 6.33497f
C5 VDD2 VDD1 0.988568f
C6 VTAIL VP 6.90602f
C7 VDD1 VP 7.32093f
C8 VTAIL VN 6.89152f
C9 VDD1 VN 0.149127f
C10 VDD2 B 5.57866f
C11 VDD1 B 5.654479f
C12 VTAIL B 8.092096f
C13 VN B 9.92062f
C14 VP B 8.213449f
C15 VDD1.n0 B 0.030846f
C16 VDD1.n1 B 0.02184f
C17 VDD1.n2 B 0.011736f
C18 VDD1.n3 B 0.02774f
C19 VDD1.n4 B 0.012426f
C20 VDD1.n5 B 0.02184f
C21 VDD1.n6 B 0.011736f
C22 VDD1.n7 B 0.02774f
C23 VDD1.n8 B 0.02774f
C24 VDD1.n9 B 0.012426f
C25 VDD1.n10 B 0.02184f
C26 VDD1.n11 B 0.011736f
C27 VDD1.n12 B 0.02774f
C28 VDD1.n13 B 0.012426f
C29 VDD1.n14 B 0.02184f
C30 VDD1.n15 B 0.011736f
C31 VDD1.n16 B 0.02774f
C32 VDD1.n17 B 0.012426f
C33 VDD1.n18 B 0.02184f
C34 VDD1.n19 B 0.011736f
C35 VDD1.n20 B 0.02774f
C36 VDD1.n21 B 0.012426f
C37 VDD1.n22 B 0.02184f
C38 VDD1.n23 B 0.011736f
C39 VDD1.n24 B 0.02774f
C40 VDD1.n25 B 0.012426f
C41 VDD1.n26 B 0.141625f
C42 VDD1.t1 B 0.045728f
C43 VDD1.n27 B 0.020805f
C44 VDD1.n28 B 0.016387f
C45 VDD1.n29 B 0.011736f
C46 VDD1.n30 B 1.40594f
C47 VDD1.n31 B 0.02184f
C48 VDD1.n32 B 0.011736f
C49 VDD1.n33 B 0.012426f
C50 VDD1.n34 B 0.02774f
C51 VDD1.n35 B 0.02774f
C52 VDD1.n36 B 0.012426f
C53 VDD1.n37 B 0.011736f
C54 VDD1.n38 B 0.02184f
C55 VDD1.n39 B 0.02184f
C56 VDD1.n40 B 0.011736f
C57 VDD1.n41 B 0.012426f
C58 VDD1.n42 B 0.02774f
C59 VDD1.n43 B 0.02774f
C60 VDD1.n44 B 0.012426f
C61 VDD1.n45 B 0.011736f
C62 VDD1.n46 B 0.02184f
C63 VDD1.n47 B 0.02184f
C64 VDD1.n48 B 0.011736f
C65 VDD1.n49 B 0.012426f
C66 VDD1.n50 B 0.02774f
C67 VDD1.n51 B 0.02774f
C68 VDD1.n52 B 0.012426f
C69 VDD1.n53 B 0.011736f
C70 VDD1.n54 B 0.02184f
C71 VDD1.n55 B 0.02184f
C72 VDD1.n56 B 0.011736f
C73 VDD1.n57 B 0.012426f
C74 VDD1.n58 B 0.02774f
C75 VDD1.n59 B 0.02774f
C76 VDD1.n60 B 0.012426f
C77 VDD1.n61 B 0.011736f
C78 VDD1.n62 B 0.02184f
C79 VDD1.n63 B 0.02184f
C80 VDD1.n64 B 0.011736f
C81 VDD1.n65 B 0.012426f
C82 VDD1.n66 B 0.02774f
C83 VDD1.n67 B 0.02774f
C84 VDD1.n68 B 0.012426f
C85 VDD1.n69 B 0.011736f
C86 VDD1.n70 B 0.02184f
C87 VDD1.n71 B 0.02184f
C88 VDD1.n72 B 0.011736f
C89 VDD1.n73 B 0.012081f
C90 VDD1.n74 B 0.012081f
C91 VDD1.n75 B 0.02774f
C92 VDD1.n76 B 0.060312f
C93 VDD1.n77 B 0.012426f
C94 VDD1.n78 B 0.011736f
C95 VDD1.n79 B 0.056748f
C96 VDD1.n80 B 0.051913f
C97 VDD1.n81 B 0.030846f
C98 VDD1.n82 B 0.02184f
C99 VDD1.n83 B 0.011736f
C100 VDD1.n84 B 0.02774f
C101 VDD1.n85 B 0.012426f
C102 VDD1.n86 B 0.02184f
C103 VDD1.n87 B 0.011736f
C104 VDD1.n88 B 0.02774f
C105 VDD1.n89 B 0.012426f
C106 VDD1.n90 B 0.02184f
C107 VDD1.n91 B 0.011736f
C108 VDD1.n92 B 0.02774f
C109 VDD1.n93 B 0.012426f
C110 VDD1.n94 B 0.02184f
C111 VDD1.n95 B 0.011736f
C112 VDD1.n96 B 0.02774f
C113 VDD1.n97 B 0.012426f
C114 VDD1.n98 B 0.02184f
C115 VDD1.n99 B 0.011736f
C116 VDD1.n100 B 0.02774f
C117 VDD1.n101 B 0.012426f
C118 VDD1.n102 B 0.02184f
C119 VDD1.n103 B 0.011736f
C120 VDD1.n104 B 0.02774f
C121 VDD1.n105 B 0.012426f
C122 VDD1.n106 B 0.141625f
C123 VDD1.t5 B 0.045728f
C124 VDD1.n107 B 0.020805f
C125 VDD1.n108 B 0.016387f
C126 VDD1.n109 B 0.011736f
C127 VDD1.n110 B 1.40594f
C128 VDD1.n111 B 0.02184f
C129 VDD1.n112 B 0.011736f
C130 VDD1.n113 B 0.012426f
C131 VDD1.n114 B 0.02774f
C132 VDD1.n115 B 0.02774f
C133 VDD1.n116 B 0.012426f
C134 VDD1.n117 B 0.011736f
C135 VDD1.n118 B 0.02184f
C136 VDD1.n119 B 0.02184f
C137 VDD1.n120 B 0.011736f
C138 VDD1.n121 B 0.012426f
C139 VDD1.n122 B 0.02774f
C140 VDD1.n123 B 0.02774f
C141 VDD1.n124 B 0.012426f
C142 VDD1.n125 B 0.011736f
C143 VDD1.n126 B 0.02184f
C144 VDD1.n127 B 0.02184f
C145 VDD1.n128 B 0.011736f
C146 VDD1.n129 B 0.012426f
C147 VDD1.n130 B 0.02774f
C148 VDD1.n131 B 0.02774f
C149 VDD1.n132 B 0.012426f
C150 VDD1.n133 B 0.011736f
C151 VDD1.n134 B 0.02184f
C152 VDD1.n135 B 0.02184f
C153 VDD1.n136 B 0.011736f
C154 VDD1.n137 B 0.012426f
C155 VDD1.n138 B 0.02774f
C156 VDD1.n139 B 0.02774f
C157 VDD1.n140 B 0.012426f
C158 VDD1.n141 B 0.011736f
C159 VDD1.n142 B 0.02184f
C160 VDD1.n143 B 0.02184f
C161 VDD1.n144 B 0.011736f
C162 VDD1.n145 B 0.012426f
C163 VDD1.n146 B 0.02774f
C164 VDD1.n147 B 0.02774f
C165 VDD1.n148 B 0.02774f
C166 VDD1.n149 B 0.012426f
C167 VDD1.n150 B 0.011736f
C168 VDD1.n151 B 0.02184f
C169 VDD1.n152 B 0.02184f
C170 VDD1.n153 B 0.011736f
C171 VDD1.n154 B 0.012081f
C172 VDD1.n155 B 0.012081f
C173 VDD1.n156 B 0.02774f
C174 VDD1.n157 B 0.060312f
C175 VDD1.n158 B 0.012426f
C176 VDD1.n159 B 0.011736f
C177 VDD1.n160 B 0.056748f
C178 VDD1.n161 B 0.051492f
C179 VDD1.t4 B 0.256294f
C180 VDD1.t0 B 0.256294f
C181 VDD1.n162 B 2.3208f
C182 VDD1.n163 B 2.14066f
C183 VDD1.t3 B 0.256294f
C184 VDD1.t2 B 0.256294f
C185 VDD1.n164 B 2.31921f
C186 VDD1.n165 B 2.34018f
C187 VP.n0 B 0.03292f
C188 VP.t5 B 1.94194f
C189 VP.n1 B 0.059771f
C190 VP.n2 B 0.03292f
C191 VP.t1 B 1.94194f
C192 VP.n3 B 0.052259f
C193 VP.n4 B 0.03292f
C194 VP.t3 B 1.94194f
C195 VP.n5 B 0.059771f
C196 VP.t4 B 2.04706f
C197 VP.t2 B 1.94194f
C198 VP.n6 B 0.768719f
C199 VP.n7 B 0.760552f
C200 VP.n8 B 0.20892f
C201 VP.n9 B 0.03292f
C202 VP.n10 B 0.032111f
C203 VP.n11 B 0.052259f
C204 VP.n12 B 0.763048f
C205 VP.n13 B 1.59505f
C206 VP.t0 B 1.94194f
C207 VP.n14 B 0.763048f
C208 VP.n15 B 1.62061f
C209 VP.n16 B 0.03292f
C210 VP.n17 B 0.03292f
C211 VP.n18 B 0.032111f
C212 VP.n19 B 0.059771f
C213 VP.n20 B 0.723534f
C214 VP.n21 B 0.03292f
C215 VP.n22 B 0.03292f
C216 VP.n23 B 0.03292f
C217 VP.n24 B 0.032111f
C218 VP.n25 B 0.052259f
C219 VP.n26 B 0.763048f
C220 VP.n27 B 0.030222f
C221 VDD2.n0 B 0.030624f
C222 VDD2.n1 B 0.021683f
C223 VDD2.n2 B 0.011652f
C224 VDD2.n3 B 0.027541f
C225 VDD2.n4 B 0.012337f
C226 VDD2.n5 B 0.021683f
C227 VDD2.n6 B 0.011652f
C228 VDD2.n7 B 0.027541f
C229 VDD2.n8 B 0.012337f
C230 VDD2.n9 B 0.021683f
C231 VDD2.n10 B 0.011652f
C232 VDD2.n11 B 0.027541f
C233 VDD2.n12 B 0.012337f
C234 VDD2.n13 B 0.021683f
C235 VDD2.n14 B 0.011652f
C236 VDD2.n15 B 0.027541f
C237 VDD2.n16 B 0.012337f
C238 VDD2.n17 B 0.021683f
C239 VDD2.n18 B 0.011652f
C240 VDD2.n19 B 0.027541f
C241 VDD2.n20 B 0.012337f
C242 VDD2.n21 B 0.021683f
C243 VDD2.n22 B 0.011652f
C244 VDD2.n23 B 0.027541f
C245 VDD2.n24 B 0.012337f
C246 VDD2.n25 B 0.140608f
C247 VDD2.t5 B 0.0454f
C248 VDD2.n26 B 0.020655f
C249 VDD2.n27 B 0.016269f
C250 VDD2.n28 B 0.011652f
C251 VDD2.n29 B 1.39585f
C252 VDD2.n30 B 0.021683f
C253 VDD2.n31 B 0.011652f
C254 VDD2.n32 B 0.012337f
C255 VDD2.n33 B 0.027541f
C256 VDD2.n34 B 0.027541f
C257 VDD2.n35 B 0.012337f
C258 VDD2.n36 B 0.011652f
C259 VDD2.n37 B 0.021683f
C260 VDD2.n38 B 0.021683f
C261 VDD2.n39 B 0.011652f
C262 VDD2.n40 B 0.012337f
C263 VDD2.n41 B 0.027541f
C264 VDD2.n42 B 0.027541f
C265 VDD2.n43 B 0.012337f
C266 VDD2.n44 B 0.011652f
C267 VDD2.n45 B 0.021683f
C268 VDD2.n46 B 0.021683f
C269 VDD2.n47 B 0.011652f
C270 VDD2.n48 B 0.012337f
C271 VDD2.n49 B 0.027541f
C272 VDD2.n50 B 0.027541f
C273 VDD2.n51 B 0.012337f
C274 VDD2.n52 B 0.011652f
C275 VDD2.n53 B 0.021683f
C276 VDD2.n54 B 0.021683f
C277 VDD2.n55 B 0.011652f
C278 VDD2.n56 B 0.012337f
C279 VDD2.n57 B 0.027541f
C280 VDD2.n58 B 0.027541f
C281 VDD2.n59 B 0.012337f
C282 VDD2.n60 B 0.011652f
C283 VDD2.n61 B 0.021683f
C284 VDD2.n62 B 0.021683f
C285 VDD2.n63 B 0.011652f
C286 VDD2.n64 B 0.012337f
C287 VDD2.n65 B 0.027541f
C288 VDD2.n66 B 0.027541f
C289 VDD2.n67 B 0.027541f
C290 VDD2.n68 B 0.012337f
C291 VDD2.n69 B 0.011652f
C292 VDD2.n70 B 0.021683f
C293 VDD2.n71 B 0.021683f
C294 VDD2.n72 B 0.011652f
C295 VDD2.n73 B 0.011994f
C296 VDD2.n74 B 0.011994f
C297 VDD2.n75 B 0.027541f
C298 VDD2.n76 B 0.059879f
C299 VDD2.n77 B 0.012337f
C300 VDD2.n78 B 0.011652f
C301 VDD2.n79 B 0.056341f
C302 VDD2.n80 B 0.051122f
C303 VDD2.t0 B 0.254453f
C304 VDD2.t1 B 0.254453f
C305 VDD2.n81 B 2.30414f
C306 VDD2.n82 B 2.04166f
C307 VDD2.n83 B 0.030624f
C308 VDD2.n84 B 0.021683f
C309 VDD2.n85 B 0.011652f
C310 VDD2.n86 B 0.027541f
C311 VDD2.n87 B 0.012337f
C312 VDD2.n88 B 0.021683f
C313 VDD2.n89 B 0.011652f
C314 VDD2.n90 B 0.027541f
C315 VDD2.n91 B 0.027541f
C316 VDD2.n92 B 0.012337f
C317 VDD2.n93 B 0.021683f
C318 VDD2.n94 B 0.011652f
C319 VDD2.n95 B 0.027541f
C320 VDD2.n96 B 0.012337f
C321 VDD2.n97 B 0.021683f
C322 VDD2.n98 B 0.011652f
C323 VDD2.n99 B 0.027541f
C324 VDD2.n100 B 0.012337f
C325 VDD2.n101 B 0.021683f
C326 VDD2.n102 B 0.011652f
C327 VDD2.n103 B 0.027541f
C328 VDD2.n104 B 0.012337f
C329 VDD2.n105 B 0.021683f
C330 VDD2.n106 B 0.011652f
C331 VDD2.n107 B 0.027541f
C332 VDD2.n108 B 0.012337f
C333 VDD2.n109 B 0.140608f
C334 VDD2.t2 B 0.0454f
C335 VDD2.n110 B 0.020655f
C336 VDD2.n111 B 0.016269f
C337 VDD2.n112 B 0.011652f
C338 VDD2.n113 B 1.39585f
C339 VDD2.n114 B 0.021683f
C340 VDD2.n115 B 0.011652f
C341 VDD2.n116 B 0.012337f
C342 VDD2.n117 B 0.027541f
C343 VDD2.n118 B 0.027541f
C344 VDD2.n119 B 0.012337f
C345 VDD2.n120 B 0.011652f
C346 VDD2.n121 B 0.021683f
C347 VDD2.n122 B 0.021683f
C348 VDD2.n123 B 0.011652f
C349 VDD2.n124 B 0.012337f
C350 VDD2.n125 B 0.027541f
C351 VDD2.n126 B 0.027541f
C352 VDD2.n127 B 0.012337f
C353 VDD2.n128 B 0.011652f
C354 VDD2.n129 B 0.021683f
C355 VDD2.n130 B 0.021683f
C356 VDD2.n131 B 0.011652f
C357 VDD2.n132 B 0.012337f
C358 VDD2.n133 B 0.027541f
C359 VDD2.n134 B 0.027541f
C360 VDD2.n135 B 0.012337f
C361 VDD2.n136 B 0.011652f
C362 VDD2.n137 B 0.021683f
C363 VDD2.n138 B 0.021683f
C364 VDD2.n139 B 0.011652f
C365 VDD2.n140 B 0.012337f
C366 VDD2.n141 B 0.027541f
C367 VDD2.n142 B 0.027541f
C368 VDD2.n143 B 0.012337f
C369 VDD2.n144 B 0.011652f
C370 VDD2.n145 B 0.021683f
C371 VDD2.n146 B 0.021683f
C372 VDD2.n147 B 0.011652f
C373 VDD2.n148 B 0.012337f
C374 VDD2.n149 B 0.027541f
C375 VDD2.n150 B 0.027541f
C376 VDD2.n151 B 0.012337f
C377 VDD2.n152 B 0.011652f
C378 VDD2.n153 B 0.021683f
C379 VDD2.n154 B 0.021683f
C380 VDD2.n155 B 0.011652f
C381 VDD2.n156 B 0.011994f
C382 VDD2.n157 B 0.011994f
C383 VDD2.n158 B 0.027541f
C384 VDD2.n159 B 0.059879f
C385 VDD2.n160 B 0.012337f
C386 VDD2.n161 B 0.011652f
C387 VDD2.n162 B 0.056341f
C388 VDD2.n163 B 0.048642f
C389 VDD2.n164 B 2.14425f
C390 VDD2.t4 B 0.254453f
C391 VDD2.t3 B 0.254453f
C392 VDD2.n165 B 2.30411f
C393 VTAIL.t6 B 0.267681f
C394 VTAIL.t9 B 0.267681f
C395 VTAIL.n0 B 2.36064f
C396 VTAIL.n1 B 0.33682f
C397 VTAIL.n2 B 0.032216f
C398 VTAIL.n3 B 0.022811f
C399 VTAIL.n4 B 0.012257f
C400 VTAIL.n5 B 0.028972f
C401 VTAIL.n6 B 0.012978f
C402 VTAIL.n7 B 0.022811f
C403 VTAIL.n8 B 0.012257f
C404 VTAIL.n9 B 0.028972f
C405 VTAIL.n10 B 0.012978f
C406 VTAIL.n11 B 0.022811f
C407 VTAIL.n12 B 0.012257f
C408 VTAIL.n13 B 0.028972f
C409 VTAIL.n14 B 0.012978f
C410 VTAIL.n15 B 0.022811f
C411 VTAIL.n16 B 0.012257f
C412 VTAIL.n17 B 0.028972f
C413 VTAIL.n18 B 0.012978f
C414 VTAIL.n19 B 0.022811f
C415 VTAIL.n20 B 0.012257f
C416 VTAIL.n21 B 0.028972f
C417 VTAIL.n22 B 0.012978f
C418 VTAIL.n23 B 0.022811f
C419 VTAIL.n24 B 0.012257f
C420 VTAIL.n25 B 0.028972f
C421 VTAIL.n26 B 0.012978f
C422 VTAIL.n27 B 0.147918f
C423 VTAIL.t4 B 0.04776f
C424 VTAIL.n28 B 0.021729f
C425 VTAIL.n29 B 0.017115f
C426 VTAIL.n30 B 0.012257f
C427 VTAIL.n31 B 1.46841f
C428 VTAIL.n32 B 0.022811f
C429 VTAIL.n33 B 0.012257f
C430 VTAIL.n34 B 0.012978f
C431 VTAIL.n35 B 0.028972f
C432 VTAIL.n36 B 0.028972f
C433 VTAIL.n37 B 0.012978f
C434 VTAIL.n38 B 0.012257f
C435 VTAIL.n39 B 0.022811f
C436 VTAIL.n40 B 0.022811f
C437 VTAIL.n41 B 0.012257f
C438 VTAIL.n42 B 0.012978f
C439 VTAIL.n43 B 0.028972f
C440 VTAIL.n44 B 0.028972f
C441 VTAIL.n45 B 0.012978f
C442 VTAIL.n46 B 0.012257f
C443 VTAIL.n47 B 0.022811f
C444 VTAIL.n48 B 0.022811f
C445 VTAIL.n49 B 0.012257f
C446 VTAIL.n50 B 0.012978f
C447 VTAIL.n51 B 0.028972f
C448 VTAIL.n52 B 0.028972f
C449 VTAIL.n53 B 0.012978f
C450 VTAIL.n54 B 0.012257f
C451 VTAIL.n55 B 0.022811f
C452 VTAIL.n56 B 0.022811f
C453 VTAIL.n57 B 0.012257f
C454 VTAIL.n58 B 0.012978f
C455 VTAIL.n59 B 0.028972f
C456 VTAIL.n60 B 0.028972f
C457 VTAIL.n61 B 0.012978f
C458 VTAIL.n62 B 0.012257f
C459 VTAIL.n63 B 0.022811f
C460 VTAIL.n64 B 0.022811f
C461 VTAIL.n65 B 0.012257f
C462 VTAIL.n66 B 0.012978f
C463 VTAIL.n67 B 0.028972f
C464 VTAIL.n68 B 0.028972f
C465 VTAIL.n69 B 0.028972f
C466 VTAIL.n70 B 0.012978f
C467 VTAIL.n71 B 0.012257f
C468 VTAIL.n72 B 0.022811f
C469 VTAIL.n73 B 0.022811f
C470 VTAIL.n74 B 0.012257f
C471 VTAIL.n75 B 0.012618f
C472 VTAIL.n76 B 0.012618f
C473 VTAIL.n77 B 0.028972f
C474 VTAIL.n78 B 0.062992f
C475 VTAIL.n79 B 0.012978f
C476 VTAIL.n80 B 0.012257f
C477 VTAIL.n81 B 0.05927f
C478 VTAIL.n82 B 0.035465f
C479 VTAIL.n83 B 0.226897f
C480 VTAIL.t3 B 0.267681f
C481 VTAIL.t1 B 0.267681f
C482 VTAIL.n84 B 2.36064f
C483 VTAIL.n85 B 1.80257f
C484 VTAIL.t8 B 0.267681f
C485 VTAIL.t11 B 0.267681f
C486 VTAIL.n86 B 2.36065f
C487 VTAIL.n87 B 1.80256f
C488 VTAIL.n88 B 0.032216f
C489 VTAIL.n89 B 0.022811f
C490 VTAIL.n90 B 0.012257f
C491 VTAIL.n91 B 0.028972f
C492 VTAIL.n92 B 0.012978f
C493 VTAIL.n93 B 0.022811f
C494 VTAIL.n94 B 0.012257f
C495 VTAIL.n95 B 0.028972f
C496 VTAIL.n96 B 0.028972f
C497 VTAIL.n97 B 0.012978f
C498 VTAIL.n98 B 0.022811f
C499 VTAIL.n99 B 0.012257f
C500 VTAIL.n100 B 0.028972f
C501 VTAIL.n101 B 0.012978f
C502 VTAIL.n102 B 0.022811f
C503 VTAIL.n103 B 0.012257f
C504 VTAIL.n104 B 0.028972f
C505 VTAIL.n105 B 0.012978f
C506 VTAIL.n106 B 0.022811f
C507 VTAIL.n107 B 0.012257f
C508 VTAIL.n108 B 0.028972f
C509 VTAIL.n109 B 0.012978f
C510 VTAIL.n110 B 0.022811f
C511 VTAIL.n111 B 0.012257f
C512 VTAIL.n112 B 0.028972f
C513 VTAIL.n113 B 0.012978f
C514 VTAIL.n114 B 0.147918f
C515 VTAIL.t10 B 0.04776f
C516 VTAIL.n115 B 0.021729f
C517 VTAIL.n116 B 0.017115f
C518 VTAIL.n117 B 0.012257f
C519 VTAIL.n118 B 1.46841f
C520 VTAIL.n119 B 0.022811f
C521 VTAIL.n120 B 0.012257f
C522 VTAIL.n121 B 0.012978f
C523 VTAIL.n122 B 0.028972f
C524 VTAIL.n123 B 0.028972f
C525 VTAIL.n124 B 0.012978f
C526 VTAIL.n125 B 0.012257f
C527 VTAIL.n126 B 0.022811f
C528 VTAIL.n127 B 0.022811f
C529 VTAIL.n128 B 0.012257f
C530 VTAIL.n129 B 0.012978f
C531 VTAIL.n130 B 0.028972f
C532 VTAIL.n131 B 0.028972f
C533 VTAIL.n132 B 0.012978f
C534 VTAIL.n133 B 0.012257f
C535 VTAIL.n134 B 0.022811f
C536 VTAIL.n135 B 0.022811f
C537 VTAIL.n136 B 0.012257f
C538 VTAIL.n137 B 0.012978f
C539 VTAIL.n138 B 0.028972f
C540 VTAIL.n139 B 0.028972f
C541 VTAIL.n140 B 0.012978f
C542 VTAIL.n141 B 0.012257f
C543 VTAIL.n142 B 0.022811f
C544 VTAIL.n143 B 0.022811f
C545 VTAIL.n144 B 0.012257f
C546 VTAIL.n145 B 0.012978f
C547 VTAIL.n146 B 0.028972f
C548 VTAIL.n147 B 0.028972f
C549 VTAIL.n148 B 0.012978f
C550 VTAIL.n149 B 0.012257f
C551 VTAIL.n150 B 0.022811f
C552 VTAIL.n151 B 0.022811f
C553 VTAIL.n152 B 0.012257f
C554 VTAIL.n153 B 0.012978f
C555 VTAIL.n154 B 0.028972f
C556 VTAIL.n155 B 0.028972f
C557 VTAIL.n156 B 0.012978f
C558 VTAIL.n157 B 0.012257f
C559 VTAIL.n158 B 0.022811f
C560 VTAIL.n159 B 0.022811f
C561 VTAIL.n160 B 0.012257f
C562 VTAIL.n161 B 0.012618f
C563 VTAIL.n162 B 0.012618f
C564 VTAIL.n163 B 0.028972f
C565 VTAIL.n164 B 0.062992f
C566 VTAIL.n165 B 0.012978f
C567 VTAIL.n166 B 0.012257f
C568 VTAIL.n167 B 0.05927f
C569 VTAIL.n168 B 0.035465f
C570 VTAIL.n169 B 0.226897f
C571 VTAIL.t0 B 0.267681f
C572 VTAIL.t5 B 0.267681f
C573 VTAIL.n170 B 2.36065f
C574 VTAIL.n171 B 0.417122f
C575 VTAIL.n172 B 0.032216f
C576 VTAIL.n173 B 0.022811f
C577 VTAIL.n174 B 0.012257f
C578 VTAIL.n175 B 0.028972f
C579 VTAIL.n176 B 0.012978f
C580 VTAIL.n177 B 0.022811f
C581 VTAIL.n178 B 0.012257f
C582 VTAIL.n179 B 0.028972f
C583 VTAIL.n180 B 0.028972f
C584 VTAIL.n181 B 0.012978f
C585 VTAIL.n182 B 0.022811f
C586 VTAIL.n183 B 0.012257f
C587 VTAIL.n184 B 0.028972f
C588 VTAIL.n185 B 0.012978f
C589 VTAIL.n186 B 0.022811f
C590 VTAIL.n187 B 0.012257f
C591 VTAIL.n188 B 0.028972f
C592 VTAIL.n189 B 0.012978f
C593 VTAIL.n190 B 0.022811f
C594 VTAIL.n191 B 0.012257f
C595 VTAIL.n192 B 0.028972f
C596 VTAIL.n193 B 0.012978f
C597 VTAIL.n194 B 0.022811f
C598 VTAIL.n195 B 0.012257f
C599 VTAIL.n196 B 0.028972f
C600 VTAIL.n197 B 0.012978f
C601 VTAIL.n198 B 0.147918f
C602 VTAIL.t2 B 0.04776f
C603 VTAIL.n199 B 0.021729f
C604 VTAIL.n200 B 0.017115f
C605 VTAIL.n201 B 0.012257f
C606 VTAIL.n202 B 1.46841f
C607 VTAIL.n203 B 0.022811f
C608 VTAIL.n204 B 0.012257f
C609 VTAIL.n205 B 0.012978f
C610 VTAIL.n206 B 0.028972f
C611 VTAIL.n207 B 0.028972f
C612 VTAIL.n208 B 0.012978f
C613 VTAIL.n209 B 0.012257f
C614 VTAIL.n210 B 0.022811f
C615 VTAIL.n211 B 0.022811f
C616 VTAIL.n212 B 0.012257f
C617 VTAIL.n213 B 0.012978f
C618 VTAIL.n214 B 0.028972f
C619 VTAIL.n215 B 0.028972f
C620 VTAIL.n216 B 0.012978f
C621 VTAIL.n217 B 0.012257f
C622 VTAIL.n218 B 0.022811f
C623 VTAIL.n219 B 0.022811f
C624 VTAIL.n220 B 0.012257f
C625 VTAIL.n221 B 0.012978f
C626 VTAIL.n222 B 0.028972f
C627 VTAIL.n223 B 0.028972f
C628 VTAIL.n224 B 0.012978f
C629 VTAIL.n225 B 0.012257f
C630 VTAIL.n226 B 0.022811f
C631 VTAIL.n227 B 0.022811f
C632 VTAIL.n228 B 0.012257f
C633 VTAIL.n229 B 0.012978f
C634 VTAIL.n230 B 0.028972f
C635 VTAIL.n231 B 0.028972f
C636 VTAIL.n232 B 0.012978f
C637 VTAIL.n233 B 0.012257f
C638 VTAIL.n234 B 0.022811f
C639 VTAIL.n235 B 0.022811f
C640 VTAIL.n236 B 0.012257f
C641 VTAIL.n237 B 0.012978f
C642 VTAIL.n238 B 0.028972f
C643 VTAIL.n239 B 0.028972f
C644 VTAIL.n240 B 0.012978f
C645 VTAIL.n241 B 0.012257f
C646 VTAIL.n242 B 0.022811f
C647 VTAIL.n243 B 0.022811f
C648 VTAIL.n244 B 0.012257f
C649 VTAIL.n245 B 0.012618f
C650 VTAIL.n246 B 0.012618f
C651 VTAIL.n247 B 0.028972f
C652 VTAIL.n248 B 0.062992f
C653 VTAIL.n249 B 0.012978f
C654 VTAIL.n250 B 0.012257f
C655 VTAIL.n251 B 0.05927f
C656 VTAIL.n252 B 0.035465f
C657 VTAIL.n253 B 1.49955f
C658 VTAIL.n254 B 0.032216f
C659 VTAIL.n255 B 0.022811f
C660 VTAIL.n256 B 0.012257f
C661 VTAIL.n257 B 0.028972f
C662 VTAIL.n258 B 0.012978f
C663 VTAIL.n259 B 0.022811f
C664 VTAIL.n260 B 0.012257f
C665 VTAIL.n261 B 0.028972f
C666 VTAIL.n262 B 0.012978f
C667 VTAIL.n263 B 0.022811f
C668 VTAIL.n264 B 0.012257f
C669 VTAIL.n265 B 0.028972f
C670 VTAIL.n266 B 0.012978f
C671 VTAIL.n267 B 0.022811f
C672 VTAIL.n268 B 0.012257f
C673 VTAIL.n269 B 0.028972f
C674 VTAIL.n270 B 0.012978f
C675 VTAIL.n271 B 0.022811f
C676 VTAIL.n272 B 0.012257f
C677 VTAIL.n273 B 0.028972f
C678 VTAIL.n274 B 0.012978f
C679 VTAIL.n275 B 0.022811f
C680 VTAIL.n276 B 0.012257f
C681 VTAIL.n277 B 0.028972f
C682 VTAIL.n278 B 0.012978f
C683 VTAIL.n279 B 0.147918f
C684 VTAIL.t7 B 0.04776f
C685 VTAIL.n280 B 0.021729f
C686 VTAIL.n281 B 0.017115f
C687 VTAIL.n282 B 0.012257f
C688 VTAIL.n283 B 1.46841f
C689 VTAIL.n284 B 0.022811f
C690 VTAIL.n285 B 0.012257f
C691 VTAIL.n286 B 0.012978f
C692 VTAIL.n287 B 0.028972f
C693 VTAIL.n288 B 0.028972f
C694 VTAIL.n289 B 0.012978f
C695 VTAIL.n290 B 0.012257f
C696 VTAIL.n291 B 0.022811f
C697 VTAIL.n292 B 0.022811f
C698 VTAIL.n293 B 0.012257f
C699 VTAIL.n294 B 0.012978f
C700 VTAIL.n295 B 0.028972f
C701 VTAIL.n296 B 0.028972f
C702 VTAIL.n297 B 0.012978f
C703 VTAIL.n298 B 0.012257f
C704 VTAIL.n299 B 0.022811f
C705 VTAIL.n300 B 0.022811f
C706 VTAIL.n301 B 0.012257f
C707 VTAIL.n302 B 0.012978f
C708 VTAIL.n303 B 0.028972f
C709 VTAIL.n304 B 0.028972f
C710 VTAIL.n305 B 0.012978f
C711 VTAIL.n306 B 0.012257f
C712 VTAIL.n307 B 0.022811f
C713 VTAIL.n308 B 0.022811f
C714 VTAIL.n309 B 0.012257f
C715 VTAIL.n310 B 0.012978f
C716 VTAIL.n311 B 0.028972f
C717 VTAIL.n312 B 0.028972f
C718 VTAIL.n313 B 0.012978f
C719 VTAIL.n314 B 0.012257f
C720 VTAIL.n315 B 0.022811f
C721 VTAIL.n316 B 0.022811f
C722 VTAIL.n317 B 0.012257f
C723 VTAIL.n318 B 0.012978f
C724 VTAIL.n319 B 0.028972f
C725 VTAIL.n320 B 0.028972f
C726 VTAIL.n321 B 0.028972f
C727 VTAIL.n322 B 0.012978f
C728 VTAIL.n323 B 0.012257f
C729 VTAIL.n324 B 0.022811f
C730 VTAIL.n325 B 0.022811f
C731 VTAIL.n326 B 0.012257f
C732 VTAIL.n327 B 0.012618f
C733 VTAIL.n328 B 0.012618f
C734 VTAIL.n329 B 0.028972f
C735 VTAIL.n330 B 0.062992f
C736 VTAIL.n331 B 0.012978f
C737 VTAIL.n332 B 0.012257f
C738 VTAIL.n333 B 0.05927f
C739 VTAIL.n334 B 0.035465f
C740 VTAIL.n335 B 1.46708f
C741 VN.n0 B 0.032526f
C742 VN.t4 B 1.91867f
C743 VN.n1 B 0.059055f
C744 VN.t0 B 2.02252f
C745 VN.t5 B 1.91867f
C746 VN.n2 B 0.759505f
C747 VN.n3 B 0.751435f
C748 VN.n4 B 0.206415f
C749 VN.n5 B 0.032526f
C750 VN.n6 B 0.031727f
C751 VN.n7 B 0.051633f
C752 VN.n8 B 0.753902f
C753 VN.n9 B 0.02986f
C754 VN.n10 B 0.032526f
C755 VN.t3 B 1.91867f
C756 VN.n11 B 0.059055f
C757 VN.t2 B 2.02252f
C758 VN.t1 B 1.91867f
C759 VN.n12 B 0.759505f
C760 VN.n13 B 0.751435f
C761 VN.n14 B 0.206415f
C762 VN.n15 B 0.032526f
C763 VN.n16 B 0.031727f
C764 VN.n17 B 0.051633f
C765 VN.n18 B 0.753902f
C766 VN.n19 B 1.59716f
.ends

