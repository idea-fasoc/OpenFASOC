* NGSPICE file created from diff_pair_sample_0615.ext - technology: sky130A

.subckt diff_pair_sample_0615 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=2.6928 ps=16.65 w=16.32 l=0.94
X1 B.t11 B.t9 B.t10 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=0 ps=0 w=16.32 l=0.94
X2 B.t8 B.t6 B.t7 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=0 ps=0 w=16.32 l=0.94
X3 VTAIL.t7 VN.t1 VDD2.t4 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=2.6928 ps=16.65 w=16.32 l=0.94
X4 B.t5 B.t3 B.t4 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=0 ps=0 w=16.32 l=0.94
X5 VTAIL.t1 VP.t0 VDD1.t5 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=2.6928 ps=16.65 w=16.32 l=0.94
X6 VTAIL.t10 VN.t2 VDD2.t3 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=2.6928 ps=16.65 w=16.32 l=0.94
X7 VDD2.t2 VN.t3 VTAIL.t11 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=2.6928 ps=16.65 w=16.32 l=0.94
X8 VDD2.t1 VN.t4 VTAIL.t9 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=6.3648 ps=33.42 w=16.32 l=0.94
X9 VTAIL.t0 VP.t1 VDD1.t4 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=2.6928 ps=16.65 w=16.32 l=0.94
X10 VDD1.t3 VP.t2 VTAIL.t4 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=6.3648 ps=33.42 w=16.32 l=0.94
X11 B.t2 B.t0 B.t1 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=0 ps=0 w=16.32 l=0.94
X12 VDD1.t2 VP.t3 VTAIL.t2 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=2.6928 ps=16.65 w=16.32 l=0.94
X13 VDD1.t1 VP.t4 VTAIL.t3 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=6.3648 pd=33.42 as=2.6928 ps=16.65 w=16.32 l=0.94
X14 VDD1.t0 VP.t5 VTAIL.t5 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=6.3648 ps=33.42 w=16.32 l=0.94
X15 VDD2.t0 VN.t5 VTAIL.t6 w_n1986_n4232# sky130_fd_pr__pfet_01v8 ad=2.6928 pd=16.65 as=6.3648 ps=33.42 w=16.32 l=0.94
R0 VN.n2 VN.t0 478.572
R1 VN.n10 VN.t4 478.572
R2 VN.n6 VN.t5 460.207
R3 VN.n14 VN.t3 460.207
R4 VN.n1 VN.t1 418.418
R5 VN.n9 VN.t2 418.418
R6 VN.n7 VN.n6 161.3
R7 VN.n15 VN.n14 161.3
R8 VN.n13 VN.n8 161.3
R9 VN.n12 VN.n11 161.3
R10 VN.n5 VN.n0 161.3
R11 VN.n4 VN.n3 161.3
R12 VN.n5 VN.n4 51.7179
R13 VN.n13 VN.n12 51.7179
R14 VN VN.n15 45.8471
R15 VN.n11 VN.n10 43.341
R16 VN.n3 VN.n2 43.341
R17 VN.n2 VN.n1 42.4561
R18 VN.n10 VN.n9 42.4561
R19 VN.n4 VN.n1 12.2964
R20 VN.n12 VN.n9 12.2964
R21 VN.n6 VN.n5 7.30353
R22 VN.n14 VN.n13 7.30353
R23 VN.n15 VN.n8 0.189894
R24 VN.n11 VN.n8 0.189894
R25 VN.n3 VN.n0 0.189894
R26 VN.n7 VN.n0 0.189894
R27 VN VN.n7 0.0516364
R28 VTAIL.n7 VTAIL.t9 52.5771
R29 VTAIL.n11 VTAIL.t6 52.5769
R30 VTAIL.n2 VTAIL.t5 52.5769
R31 VTAIL.n10 VTAIL.t4 52.5769
R32 VTAIL.n9 VTAIL.n8 50.5854
R33 VTAIL.n6 VTAIL.n5 50.5854
R34 VTAIL.n1 VTAIL.n0 50.5852
R35 VTAIL.n4 VTAIL.n3 50.5852
R36 VTAIL.n6 VTAIL.n4 28.6255
R37 VTAIL.n11 VTAIL.n10 27.5307
R38 VTAIL.n0 VTAIL.t8 1.99223
R39 VTAIL.n0 VTAIL.t7 1.99223
R40 VTAIL.n3 VTAIL.t3 1.99223
R41 VTAIL.n3 VTAIL.t1 1.99223
R42 VTAIL.n8 VTAIL.t2 1.99223
R43 VTAIL.n8 VTAIL.t0 1.99223
R44 VTAIL.n5 VTAIL.t11 1.99223
R45 VTAIL.n5 VTAIL.t10 1.99223
R46 VTAIL.n7 VTAIL.n6 1.09533
R47 VTAIL.n10 VTAIL.n9 1.09533
R48 VTAIL.n4 VTAIL.n2 1.09533
R49 VTAIL.n9 VTAIL.n7 1.01774
R50 VTAIL.n2 VTAIL.n1 1.01774
R51 VTAIL VTAIL.n11 0.763431
R52 VTAIL VTAIL.n1 0.332397
R53 VDD2.n1 VDD2.t5 70.0214
R54 VDD2.n2 VDD2.t2 69.2559
R55 VDD2.n1 VDD2.n0 67.4823
R56 VDD2 VDD2.n3 67.4795
R57 VDD2.n2 VDD2.n1 41.3424
R58 VDD2.n3 VDD2.t3 1.99223
R59 VDD2.n3 VDD2.t1 1.99223
R60 VDD2.n0 VDD2.t4 1.99223
R61 VDD2.n0 VDD2.t0 1.99223
R62 VDD2 VDD2.n2 0.87981
R63 B.n129 B.t3 620.918
R64 B.n135 B.t9 620.918
R65 B.n42 B.t6 620.918
R66 B.n49 B.t0 620.918
R67 B.n458 B.n77 585
R68 B.n460 B.n459 585
R69 B.n461 B.n76 585
R70 B.n463 B.n462 585
R71 B.n464 B.n75 585
R72 B.n466 B.n465 585
R73 B.n467 B.n74 585
R74 B.n469 B.n468 585
R75 B.n470 B.n73 585
R76 B.n472 B.n471 585
R77 B.n473 B.n72 585
R78 B.n475 B.n474 585
R79 B.n476 B.n71 585
R80 B.n478 B.n477 585
R81 B.n479 B.n70 585
R82 B.n481 B.n480 585
R83 B.n482 B.n69 585
R84 B.n484 B.n483 585
R85 B.n485 B.n68 585
R86 B.n487 B.n486 585
R87 B.n488 B.n67 585
R88 B.n490 B.n489 585
R89 B.n491 B.n66 585
R90 B.n493 B.n492 585
R91 B.n494 B.n65 585
R92 B.n496 B.n495 585
R93 B.n497 B.n64 585
R94 B.n499 B.n498 585
R95 B.n500 B.n63 585
R96 B.n502 B.n501 585
R97 B.n503 B.n62 585
R98 B.n505 B.n504 585
R99 B.n506 B.n61 585
R100 B.n508 B.n507 585
R101 B.n509 B.n60 585
R102 B.n511 B.n510 585
R103 B.n512 B.n59 585
R104 B.n514 B.n513 585
R105 B.n515 B.n58 585
R106 B.n517 B.n516 585
R107 B.n518 B.n57 585
R108 B.n520 B.n519 585
R109 B.n521 B.n56 585
R110 B.n523 B.n522 585
R111 B.n524 B.n55 585
R112 B.n526 B.n525 585
R113 B.n527 B.n54 585
R114 B.n529 B.n528 585
R115 B.n530 B.n53 585
R116 B.n532 B.n531 585
R117 B.n533 B.n52 585
R118 B.n535 B.n534 585
R119 B.n536 B.n51 585
R120 B.n538 B.n537 585
R121 B.n540 B.n48 585
R122 B.n542 B.n541 585
R123 B.n543 B.n47 585
R124 B.n545 B.n544 585
R125 B.n546 B.n46 585
R126 B.n548 B.n547 585
R127 B.n549 B.n45 585
R128 B.n551 B.n550 585
R129 B.n552 B.n41 585
R130 B.n554 B.n553 585
R131 B.n555 B.n40 585
R132 B.n557 B.n556 585
R133 B.n558 B.n39 585
R134 B.n560 B.n559 585
R135 B.n561 B.n38 585
R136 B.n563 B.n562 585
R137 B.n564 B.n37 585
R138 B.n566 B.n565 585
R139 B.n567 B.n36 585
R140 B.n569 B.n568 585
R141 B.n570 B.n35 585
R142 B.n572 B.n571 585
R143 B.n573 B.n34 585
R144 B.n575 B.n574 585
R145 B.n576 B.n33 585
R146 B.n578 B.n577 585
R147 B.n579 B.n32 585
R148 B.n581 B.n580 585
R149 B.n582 B.n31 585
R150 B.n584 B.n583 585
R151 B.n585 B.n30 585
R152 B.n587 B.n586 585
R153 B.n588 B.n29 585
R154 B.n590 B.n589 585
R155 B.n591 B.n28 585
R156 B.n593 B.n592 585
R157 B.n594 B.n27 585
R158 B.n596 B.n595 585
R159 B.n597 B.n26 585
R160 B.n599 B.n598 585
R161 B.n600 B.n25 585
R162 B.n602 B.n601 585
R163 B.n603 B.n24 585
R164 B.n605 B.n604 585
R165 B.n606 B.n23 585
R166 B.n608 B.n607 585
R167 B.n609 B.n22 585
R168 B.n611 B.n610 585
R169 B.n612 B.n21 585
R170 B.n614 B.n613 585
R171 B.n615 B.n20 585
R172 B.n617 B.n616 585
R173 B.n618 B.n19 585
R174 B.n620 B.n619 585
R175 B.n621 B.n18 585
R176 B.n623 B.n622 585
R177 B.n624 B.n17 585
R178 B.n626 B.n625 585
R179 B.n627 B.n16 585
R180 B.n629 B.n628 585
R181 B.n630 B.n15 585
R182 B.n632 B.n631 585
R183 B.n633 B.n14 585
R184 B.n635 B.n634 585
R185 B.n457 B.n456 585
R186 B.n455 B.n78 585
R187 B.n454 B.n453 585
R188 B.n452 B.n79 585
R189 B.n451 B.n450 585
R190 B.n449 B.n80 585
R191 B.n448 B.n447 585
R192 B.n446 B.n81 585
R193 B.n445 B.n444 585
R194 B.n443 B.n82 585
R195 B.n442 B.n441 585
R196 B.n440 B.n83 585
R197 B.n439 B.n438 585
R198 B.n437 B.n84 585
R199 B.n436 B.n435 585
R200 B.n434 B.n85 585
R201 B.n433 B.n432 585
R202 B.n431 B.n86 585
R203 B.n430 B.n429 585
R204 B.n428 B.n87 585
R205 B.n427 B.n426 585
R206 B.n425 B.n88 585
R207 B.n424 B.n423 585
R208 B.n422 B.n89 585
R209 B.n421 B.n420 585
R210 B.n419 B.n90 585
R211 B.n418 B.n417 585
R212 B.n416 B.n91 585
R213 B.n415 B.n414 585
R214 B.n413 B.n92 585
R215 B.n412 B.n411 585
R216 B.n410 B.n93 585
R217 B.n409 B.n408 585
R218 B.n407 B.n94 585
R219 B.n406 B.n405 585
R220 B.n404 B.n95 585
R221 B.n403 B.n402 585
R222 B.n401 B.n96 585
R223 B.n400 B.n399 585
R224 B.n398 B.n97 585
R225 B.n397 B.n396 585
R226 B.n395 B.n98 585
R227 B.n394 B.n393 585
R228 B.n392 B.n99 585
R229 B.n391 B.n390 585
R230 B.n389 B.n100 585
R231 B.n388 B.n387 585
R232 B.n209 B.n164 585
R233 B.n211 B.n210 585
R234 B.n212 B.n163 585
R235 B.n214 B.n213 585
R236 B.n215 B.n162 585
R237 B.n217 B.n216 585
R238 B.n218 B.n161 585
R239 B.n220 B.n219 585
R240 B.n221 B.n160 585
R241 B.n223 B.n222 585
R242 B.n224 B.n159 585
R243 B.n226 B.n225 585
R244 B.n227 B.n158 585
R245 B.n229 B.n228 585
R246 B.n230 B.n157 585
R247 B.n232 B.n231 585
R248 B.n233 B.n156 585
R249 B.n235 B.n234 585
R250 B.n236 B.n155 585
R251 B.n238 B.n237 585
R252 B.n239 B.n154 585
R253 B.n241 B.n240 585
R254 B.n242 B.n153 585
R255 B.n244 B.n243 585
R256 B.n245 B.n152 585
R257 B.n247 B.n246 585
R258 B.n248 B.n151 585
R259 B.n250 B.n249 585
R260 B.n251 B.n150 585
R261 B.n253 B.n252 585
R262 B.n254 B.n149 585
R263 B.n256 B.n255 585
R264 B.n257 B.n148 585
R265 B.n259 B.n258 585
R266 B.n260 B.n147 585
R267 B.n262 B.n261 585
R268 B.n263 B.n146 585
R269 B.n265 B.n264 585
R270 B.n266 B.n145 585
R271 B.n268 B.n267 585
R272 B.n269 B.n144 585
R273 B.n271 B.n270 585
R274 B.n272 B.n143 585
R275 B.n274 B.n273 585
R276 B.n275 B.n142 585
R277 B.n277 B.n276 585
R278 B.n278 B.n141 585
R279 B.n280 B.n279 585
R280 B.n281 B.n140 585
R281 B.n283 B.n282 585
R282 B.n284 B.n139 585
R283 B.n286 B.n285 585
R284 B.n287 B.n138 585
R285 B.n289 B.n288 585
R286 B.n291 B.n290 585
R287 B.n292 B.n134 585
R288 B.n294 B.n293 585
R289 B.n295 B.n133 585
R290 B.n297 B.n296 585
R291 B.n298 B.n132 585
R292 B.n300 B.n299 585
R293 B.n301 B.n131 585
R294 B.n303 B.n302 585
R295 B.n304 B.n128 585
R296 B.n307 B.n306 585
R297 B.n308 B.n127 585
R298 B.n310 B.n309 585
R299 B.n311 B.n126 585
R300 B.n313 B.n312 585
R301 B.n314 B.n125 585
R302 B.n316 B.n315 585
R303 B.n317 B.n124 585
R304 B.n319 B.n318 585
R305 B.n320 B.n123 585
R306 B.n322 B.n321 585
R307 B.n323 B.n122 585
R308 B.n325 B.n324 585
R309 B.n326 B.n121 585
R310 B.n328 B.n327 585
R311 B.n329 B.n120 585
R312 B.n331 B.n330 585
R313 B.n332 B.n119 585
R314 B.n334 B.n333 585
R315 B.n335 B.n118 585
R316 B.n337 B.n336 585
R317 B.n338 B.n117 585
R318 B.n340 B.n339 585
R319 B.n341 B.n116 585
R320 B.n343 B.n342 585
R321 B.n344 B.n115 585
R322 B.n346 B.n345 585
R323 B.n347 B.n114 585
R324 B.n349 B.n348 585
R325 B.n350 B.n113 585
R326 B.n352 B.n351 585
R327 B.n353 B.n112 585
R328 B.n355 B.n354 585
R329 B.n356 B.n111 585
R330 B.n358 B.n357 585
R331 B.n359 B.n110 585
R332 B.n361 B.n360 585
R333 B.n362 B.n109 585
R334 B.n364 B.n363 585
R335 B.n365 B.n108 585
R336 B.n367 B.n366 585
R337 B.n368 B.n107 585
R338 B.n370 B.n369 585
R339 B.n371 B.n106 585
R340 B.n373 B.n372 585
R341 B.n374 B.n105 585
R342 B.n376 B.n375 585
R343 B.n377 B.n104 585
R344 B.n379 B.n378 585
R345 B.n380 B.n103 585
R346 B.n382 B.n381 585
R347 B.n383 B.n102 585
R348 B.n385 B.n384 585
R349 B.n386 B.n101 585
R350 B.n208 B.n207 585
R351 B.n206 B.n165 585
R352 B.n205 B.n204 585
R353 B.n203 B.n166 585
R354 B.n202 B.n201 585
R355 B.n200 B.n167 585
R356 B.n199 B.n198 585
R357 B.n197 B.n168 585
R358 B.n196 B.n195 585
R359 B.n194 B.n169 585
R360 B.n193 B.n192 585
R361 B.n191 B.n170 585
R362 B.n190 B.n189 585
R363 B.n188 B.n171 585
R364 B.n187 B.n186 585
R365 B.n185 B.n172 585
R366 B.n184 B.n183 585
R367 B.n182 B.n173 585
R368 B.n181 B.n180 585
R369 B.n179 B.n174 585
R370 B.n178 B.n177 585
R371 B.n176 B.n175 585
R372 B.n2 B.n0 585
R373 B.n669 B.n1 585
R374 B.n668 B.n667 585
R375 B.n666 B.n3 585
R376 B.n665 B.n664 585
R377 B.n663 B.n4 585
R378 B.n662 B.n661 585
R379 B.n660 B.n5 585
R380 B.n659 B.n658 585
R381 B.n657 B.n6 585
R382 B.n656 B.n655 585
R383 B.n654 B.n7 585
R384 B.n653 B.n652 585
R385 B.n651 B.n8 585
R386 B.n650 B.n649 585
R387 B.n648 B.n9 585
R388 B.n647 B.n646 585
R389 B.n645 B.n10 585
R390 B.n644 B.n643 585
R391 B.n642 B.n11 585
R392 B.n641 B.n640 585
R393 B.n639 B.n12 585
R394 B.n638 B.n637 585
R395 B.n636 B.n13 585
R396 B.n671 B.n670 585
R397 B.n207 B.n164 526.135
R398 B.n634 B.n13 526.135
R399 B.n387 B.n386 526.135
R400 B.n458 B.n457 526.135
R401 B.n207 B.n206 163.367
R402 B.n206 B.n205 163.367
R403 B.n205 B.n166 163.367
R404 B.n201 B.n166 163.367
R405 B.n201 B.n200 163.367
R406 B.n200 B.n199 163.367
R407 B.n199 B.n168 163.367
R408 B.n195 B.n168 163.367
R409 B.n195 B.n194 163.367
R410 B.n194 B.n193 163.367
R411 B.n193 B.n170 163.367
R412 B.n189 B.n170 163.367
R413 B.n189 B.n188 163.367
R414 B.n188 B.n187 163.367
R415 B.n187 B.n172 163.367
R416 B.n183 B.n172 163.367
R417 B.n183 B.n182 163.367
R418 B.n182 B.n181 163.367
R419 B.n181 B.n174 163.367
R420 B.n177 B.n174 163.367
R421 B.n177 B.n176 163.367
R422 B.n176 B.n2 163.367
R423 B.n670 B.n2 163.367
R424 B.n670 B.n669 163.367
R425 B.n669 B.n668 163.367
R426 B.n668 B.n3 163.367
R427 B.n664 B.n3 163.367
R428 B.n664 B.n663 163.367
R429 B.n663 B.n662 163.367
R430 B.n662 B.n5 163.367
R431 B.n658 B.n5 163.367
R432 B.n658 B.n657 163.367
R433 B.n657 B.n656 163.367
R434 B.n656 B.n7 163.367
R435 B.n652 B.n7 163.367
R436 B.n652 B.n651 163.367
R437 B.n651 B.n650 163.367
R438 B.n650 B.n9 163.367
R439 B.n646 B.n9 163.367
R440 B.n646 B.n645 163.367
R441 B.n645 B.n644 163.367
R442 B.n644 B.n11 163.367
R443 B.n640 B.n11 163.367
R444 B.n640 B.n639 163.367
R445 B.n639 B.n638 163.367
R446 B.n638 B.n13 163.367
R447 B.n211 B.n164 163.367
R448 B.n212 B.n211 163.367
R449 B.n213 B.n212 163.367
R450 B.n213 B.n162 163.367
R451 B.n217 B.n162 163.367
R452 B.n218 B.n217 163.367
R453 B.n219 B.n218 163.367
R454 B.n219 B.n160 163.367
R455 B.n223 B.n160 163.367
R456 B.n224 B.n223 163.367
R457 B.n225 B.n224 163.367
R458 B.n225 B.n158 163.367
R459 B.n229 B.n158 163.367
R460 B.n230 B.n229 163.367
R461 B.n231 B.n230 163.367
R462 B.n231 B.n156 163.367
R463 B.n235 B.n156 163.367
R464 B.n236 B.n235 163.367
R465 B.n237 B.n236 163.367
R466 B.n237 B.n154 163.367
R467 B.n241 B.n154 163.367
R468 B.n242 B.n241 163.367
R469 B.n243 B.n242 163.367
R470 B.n243 B.n152 163.367
R471 B.n247 B.n152 163.367
R472 B.n248 B.n247 163.367
R473 B.n249 B.n248 163.367
R474 B.n249 B.n150 163.367
R475 B.n253 B.n150 163.367
R476 B.n254 B.n253 163.367
R477 B.n255 B.n254 163.367
R478 B.n255 B.n148 163.367
R479 B.n259 B.n148 163.367
R480 B.n260 B.n259 163.367
R481 B.n261 B.n260 163.367
R482 B.n261 B.n146 163.367
R483 B.n265 B.n146 163.367
R484 B.n266 B.n265 163.367
R485 B.n267 B.n266 163.367
R486 B.n267 B.n144 163.367
R487 B.n271 B.n144 163.367
R488 B.n272 B.n271 163.367
R489 B.n273 B.n272 163.367
R490 B.n273 B.n142 163.367
R491 B.n277 B.n142 163.367
R492 B.n278 B.n277 163.367
R493 B.n279 B.n278 163.367
R494 B.n279 B.n140 163.367
R495 B.n283 B.n140 163.367
R496 B.n284 B.n283 163.367
R497 B.n285 B.n284 163.367
R498 B.n285 B.n138 163.367
R499 B.n289 B.n138 163.367
R500 B.n290 B.n289 163.367
R501 B.n290 B.n134 163.367
R502 B.n294 B.n134 163.367
R503 B.n295 B.n294 163.367
R504 B.n296 B.n295 163.367
R505 B.n296 B.n132 163.367
R506 B.n300 B.n132 163.367
R507 B.n301 B.n300 163.367
R508 B.n302 B.n301 163.367
R509 B.n302 B.n128 163.367
R510 B.n307 B.n128 163.367
R511 B.n308 B.n307 163.367
R512 B.n309 B.n308 163.367
R513 B.n309 B.n126 163.367
R514 B.n313 B.n126 163.367
R515 B.n314 B.n313 163.367
R516 B.n315 B.n314 163.367
R517 B.n315 B.n124 163.367
R518 B.n319 B.n124 163.367
R519 B.n320 B.n319 163.367
R520 B.n321 B.n320 163.367
R521 B.n321 B.n122 163.367
R522 B.n325 B.n122 163.367
R523 B.n326 B.n325 163.367
R524 B.n327 B.n326 163.367
R525 B.n327 B.n120 163.367
R526 B.n331 B.n120 163.367
R527 B.n332 B.n331 163.367
R528 B.n333 B.n332 163.367
R529 B.n333 B.n118 163.367
R530 B.n337 B.n118 163.367
R531 B.n338 B.n337 163.367
R532 B.n339 B.n338 163.367
R533 B.n339 B.n116 163.367
R534 B.n343 B.n116 163.367
R535 B.n344 B.n343 163.367
R536 B.n345 B.n344 163.367
R537 B.n345 B.n114 163.367
R538 B.n349 B.n114 163.367
R539 B.n350 B.n349 163.367
R540 B.n351 B.n350 163.367
R541 B.n351 B.n112 163.367
R542 B.n355 B.n112 163.367
R543 B.n356 B.n355 163.367
R544 B.n357 B.n356 163.367
R545 B.n357 B.n110 163.367
R546 B.n361 B.n110 163.367
R547 B.n362 B.n361 163.367
R548 B.n363 B.n362 163.367
R549 B.n363 B.n108 163.367
R550 B.n367 B.n108 163.367
R551 B.n368 B.n367 163.367
R552 B.n369 B.n368 163.367
R553 B.n369 B.n106 163.367
R554 B.n373 B.n106 163.367
R555 B.n374 B.n373 163.367
R556 B.n375 B.n374 163.367
R557 B.n375 B.n104 163.367
R558 B.n379 B.n104 163.367
R559 B.n380 B.n379 163.367
R560 B.n381 B.n380 163.367
R561 B.n381 B.n102 163.367
R562 B.n385 B.n102 163.367
R563 B.n386 B.n385 163.367
R564 B.n387 B.n100 163.367
R565 B.n391 B.n100 163.367
R566 B.n392 B.n391 163.367
R567 B.n393 B.n392 163.367
R568 B.n393 B.n98 163.367
R569 B.n397 B.n98 163.367
R570 B.n398 B.n397 163.367
R571 B.n399 B.n398 163.367
R572 B.n399 B.n96 163.367
R573 B.n403 B.n96 163.367
R574 B.n404 B.n403 163.367
R575 B.n405 B.n404 163.367
R576 B.n405 B.n94 163.367
R577 B.n409 B.n94 163.367
R578 B.n410 B.n409 163.367
R579 B.n411 B.n410 163.367
R580 B.n411 B.n92 163.367
R581 B.n415 B.n92 163.367
R582 B.n416 B.n415 163.367
R583 B.n417 B.n416 163.367
R584 B.n417 B.n90 163.367
R585 B.n421 B.n90 163.367
R586 B.n422 B.n421 163.367
R587 B.n423 B.n422 163.367
R588 B.n423 B.n88 163.367
R589 B.n427 B.n88 163.367
R590 B.n428 B.n427 163.367
R591 B.n429 B.n428 163.367
R592 B.n429 B.n86 163.367
R593 B.n433 B.n86 163.367
R594 B.n434 B.n433 163.367
R595 B.n435 B.n434 163.367
R596 B.n435 B.n84 163.367
R597 B.n439 B.n84 163.367
R598 B.n440 B.n439 163.367
R599 B.n441 B.n440 163.367
R600 B.n441 B.n82 163.367
R601 B.n445 B.n82 163.367
R602 B.n446 B.n445 163.367
R603 B.n447 B.n446 163.367
R604 B.n447 B.n80 163.367
R605 B.n451 B.n80 163.367
R606 B.n452 B.n451 163.367
R607 B.n453 B.n452 163.367
R608 B.n453 B.n78 163.367
R609 B.n457 B.n78 163.367
R610 B.n634 B.n633 163.367
R611 B.n633 B.n632 163.367
R612 B.n632 B.n15 163.367
R613 B.n628 B.n15 163.367
R614 B.n628 B.n627 163.367
R615 B.n627 B.n626 163.367
R616 B.n626 B.n17 163.367
R617 B.n622 B.n17 163.367
R618 B.n622 B.n621 163.367
R619 B.n621 B.n620 163.367
R620 B.n620 B.n19 163.367
R621 B.n616 B.n19 163.367
R622 B.n616 B.n615 163.367
R623 B.n615 B.n614 163.367
R624 B.n614 B.n21 163.367
R625 B.n610 B.n21 163.367
R626 B.n610 B.n609 163.367
R627 B.n609 B.n608 163.367
R628 B.n608 B.n23 163.367
R629 B.n604 B.n23 163.367
R630 B.n604 B.n603 163.367
R631 B.n603 B.n602 163.367
R632 B.n602 B.n25 163.367
R633 B.n598 B.n25 163.367
R634 B.n598 B.n597 163.367
R635 B.n597 B.n596 163.367
R636 B.n596 B.n27 163.367
R637 B.n592 B.n27 163.367
R638 B.n592 B.n591 163.367
R639 B.n591 B.n590 163.367
R640 B.n590 B.n29 163.367
R641 B.n586 B.n29 163.367
R642 B.n586 B.n585 163.367
R643 B.n585 B.n584 163.367
R644 B.n584 B.n31 163.367
R645 B.n580 B.n31 163.367
R646 B.n580 B.n579 163.367
R647 B.n579 B.n578 163.367
R648 B.n578 B.n33 163.367
R649 B.n574 B.n33 163.367
R650 B.n574 B.n573 163.367
R651 B.n573 B.n572 163.367
R652 B.n572 B.n35 163.367
R653 B.n568 B.n35 163.367
R654 B.n568 B.n567 163.367
R655 B.n567 B.n566 163.367
R656 B.n566 B.n37 163.367
R657 B.n562 B.n37 163.367
R658 B.n562 B.n561 163.367
R659 B.n561 B.n560 163.367
R660 B.n560 B.n39 163.367
R661 B.n556 B.n39 163.367
R662 B.n556 B.n555 163.367
R663 B.n555 B.n554 163.367
R664 B.n554 B.n41 163.367
R665 B.n550 B.n41 163.367
R666 B.n550 B.n549 163.367
R667 B.n549 B.n548 163.367
R668 B.n548 B.n46 163.367
R669 B.n544 B.n46 163.367
R670 B.n544 B.n543 163.367
R671 B.n543 B.n542 163.367
R672 B.n542 B.n48 163.367
R673 B.n537 B.n48 163.367
R674 B.n537 B.n536 163.367
R675 B.n536 B.n535 163.367
R676 B.n535 B.n52 163.367
R677 B.n531 B.n52 163.367
R678 B.n531 B.n530 163.367
R679 B.n530 B.n529 163.367
R680 B.n529 B.n54 163.367
R681 B.n525 B.n54 163.367
R682 B.n525 B.n524 163.367
R683 B.n524 B.n523 163.367
R684 B.n523 B.n56 163.367
R685 B.n519 B.n56 163.367
R686 B.n519 B.n518 163.367
R687 B.n518 B.n517 163.367
R688 B.n517 B.n58 163.367
R689 B.n513 B.n58 163.367
R690 B.n513 B.n512 163.367
R691 B.n512 B.n511 163.367
R692 B.n511 B.n60 163.367
R693 B.n507 B.n60 163.367
R694 B.n507 B.n506 163.367
R695 B.n506 B.n505 163.367
R696 B.n505 B.n62 163.367
R697 B.n501 B.n62 163.367
R698 B.n501 B.n500 163.367
R699 B.n500 B.n499 163.367
R700 B.n499 B.n64 163.367
R701 B.n495 B.n64 163.367
R702 B.n495 B.n494 163.367
R703 B.n494 B.n493 163.367
R704 B.n493 B.n66 163.367
R705 B.n489 B.n66 163.367
R706 B.n489 B.n488 163.367
R707 B.n488 B.n487 163.367
R708 B.n487 B.n68 163.367
R709 B.n483 B.n68 163.367
R710 B.n483 B.n482 163.367
R711 B.n482 B.n481 163.367
R712 B.n481 B.n70 163.367
R713 B.n477 B.n70 163.367
R714 B.n477 B.n476 163.367
R715 B.n476 B.n475 163.367
R716 B.n475 B.n72 163.367
R717 B.n471 B.n72 163.367
R718 B.n471 B.n470 163.367
R719 B.n470 B.n469 163.367
R720 B.n469 B.n74 163.367
R721 B.n465 B.n74 163.367
R722 B.n465 B.n464 163.367
R723 B.n464 B.n463 163.367
R724 B.n463 B.n76 163.367
R725 B.n459 B.n76 163.367
R726 B.n459 B.n458 163.367
R727 B.n129 B.t5 131.018
R728 B.n49 B.t1 131.018
R729 B.n135 B.t11 130.998
R730 B.n42 B.t7 130.998
R731 B.n130 B.t4 106.388
R732 B.n50 B.t2 106.388
R733 B.n136 B.t10 106.367
R734 B.n43 B.t8 106.367
R735 B.n305 B.n130 59.5399
R736 B.n137 B.n136 59.5399
R737 B.n44 B.n43 59.5399
R738 B.n539 B.n50 59.5399
R739 B.n636 B.n635 34.1859
R740 B.n456 B.n77 34.1859
R741 B.n388 B.n101 34.1859
R742 B.n209 B.n208 34.1859
R743 B.n130 B.n129 24.6308
R744 B.n136 B.n135 24.6308
R745 B.n43 B.n42 24.6308
R746 B.n50 B.n49 24.6308
R747 B B.n671 18.0485
R748 B.n635 B.n14 10.6151
R749 B.n631 B.n14 10.6151
R750 B.n631 B.n630 10.6151
R751 B.n630 B.n629 10.6151
R752 B.n629 B.n16 10.6151
R753 B.n625 B.n16 10.6151
R754 B.n625 B.n624 10.6151
R755 B.n624 B.n623 10.6151
R756 B.n623 B.n18 10.6151
R757 B.n619 B.n18 10.6151
R758 B.n619 B.n618 10.6151
R759 B.n618 B.n617 10.6151
R760 B.n617 B.n20 10.6151
R761 B.n613 B.n20 10.6151
R762 B.n613 B.n612 10.6151
R763 B.n612 B.n611 10.6151
R764 B.n611 B.n22 10.6151
R765 B.n607 B.n22 10.6151
R766 B.n607 B.n606 10.6151
R767 B.n606 B.n605 10.6151
R768 B.n605 B.n24 10.6151
R769 B.n601 B.n24 10.6151
R770 B.n601 B.n600 10.6151
R771 B.n600 B.n599 10.6151
R772 B.n599 B.n26 10.6151
R773 B.n595 B.n26 10.6151
R774 B.n595 B.n594 10.6151
R775 B.n594 B.n593 10.6151
R776 B.n593 B.n28 10.6151
R777 B.n589 B.n28 10.6151
R778 B.n589 B.n588 10.6151
R779 B.n588 B.n587 10.6151
R780 B.n587 B.n30 10.6151
R781 B.n583 B.n30 10.6151
R782 B.n583 B.n582 10.6151
R783 B.n582 B.n581 10.6151
R784 B.n581 B.n32 10.6151
R785 B.n577 B.n32 10.6151
R786 B.n577 B.n576 10.6151
R787 B.n576 B.n575 10.6151
R788 B.n575 B.n34 10.6151
R789 B.n571 B.n34 10.6151
R790 B.n571 B.n570 10.6151
R791 B.n570 B.n569 10.6151
R792 B.n569 B.n36 10.6151
R793 B.n565 B.n36 10.6151
R794 B.n565 B.n564 10.6151
R795 B.n564 B.n563 10.6151
R796 B.n563 B.n38 10.6151
R797 B.n559 B.n38 10.6151
R798 B.n559 B.n558 10.6151
R799 B.n558 B.n557 10.6151
R800 B.n557 B.n40 10.6151
R801 B.n553 B.n552 10.6151
R802 B.n552 B.n551 10.6151
R803 B.n551 B.n45 10.6151
R804 B.n547 B.n45 10.6151
R805 B.n547 B.n546 10.6151
R806 B.n546 B.n545 10.6151
R807 B.n545 B.n47 10.6151
R808 B.n541 B.n47 10.6151
R809 B.n541 B.n540 10.6151
R810 B.n538 B.n51 10.6151
R811 B.n534 B.n51 10.6151
R812 B.n534 B.n533 10.6151
R813 B.n533 B.n532 10.6151
R814 B.n532 B.n53 10.6151
R815 B.n528 B.n53 10.6151
R816 B.n528 B.n527 10.6151
R817 B.n527 B.n526 10.6151
R818 B.n526 B.n55 10.6151
R819 B.n522 B.n55 10.6151
R820 B.n522 B.n521 10.6151
R821 B.n521 B.n520 10.6151
R822 B.n520 B.n57 10.6151
R823 B.n516 B.n57 10.6151
R824 B.n516 B.n515 10.6151
R825 B.n515 B.n514 10.6151
R826 B.n514 B.n59 10.6151
R827 B.n510 B.n59 10.6151
R828 B.n510 B.n509 10.6151
R829 B.n509 B.n508 10.6151
R830 B.n508 B.n61 10.6151
R831 B.n504 B.n61 10.6151
R832 B.n504 B.n503 10.6151
R833 B.n503 B.n502 10.6151
R834 B.n502 B.n63 10.6151
R835 B.n498 B.n63 10.6151
R836 B.n498 B.n497 10.6151
R837 B.n497 B.n496 10.6151
R838 B.n496 B.n65 10.6151
R839 B.n492 B.n65 10.6151
R840 B.n492 B.n491 10.6151
R841 B.n491 B.n490 10.6151
R842 B.n490 B.n67 10.6151
R843 B.n486 B.n67 10.6151
R844 B.n486 B.n485 10.6151
R845 B.n485 B.n484 10.6151
R846 B.n484 B.n69 10.6151
R847 B.n480 B.n69 10.6151
R848 B.n480 B.n479 10.6151
R849 B.n479 B.n478 10.6151
R850 B.n478 B.n71 10.6151
R851 B.n474 B.n71 10.6151
R852 B.n474 B.n473 10.6151
R853 B.n473 B.n472 10.6151
R854 B.n472 B.n73 10.6151
R855 B.n468 B.n73 10.6151
R856 B.n468 B.n467 10.6151
R857 B.n467 B.n466 10.6151
R858 B.n466 B.n75 10.6151
R859 B.n462 B.n75 10.6151
R860 B.n462 B.n461 10.6151
R861 B.n461 B.n460 10.6151
R862 B.n460 B.n77 10.6151
R863 B.n389 B.n388 10.6151
R864 B.n390 B.n389 10.6151
R865 B.n390 B.n99 10.6151
R866 B.n394 B.n99 10.6151
R867 B.n395 B.n394 10.6151
R868 B.n396 B.n395 10.6151
R869 B.n396 B.n97 10.6151
R870 B.n400 B.n97 10.6151
R871 B.n401 B.n400 10.6151
R872 B.n402 B.n401 10.6151
R873 B.n402 B.n95 10.6151
R874 B.n406 B.n95 10.6151
R875 B.n407 B.n406 10.6151
R876 B.n408 B.n407 10.6151
R877 B.n408 B.n93 10.6151
R878 B.n412 B.n93 10.6151
R879 B.n413 B.n412 10.6151
R880 B.n414 B.n413 10.6151
R881 B.n414 B.n91 10.6151
R882 B.n418 B.n91 10.6151
R883 B.n419 B.n418 10.6151
R884 B.n420 B.n419 10.6151
R885 B.n420 B.n89 10.6151
R886 B.n424 B.n89 10.6151
R887 B.n425 B.n424 10.6151
R888 B.n426 B.n425 10.6151
R889 B.n426 B.n87 10.6151
R890 B.n430 B.n87 10.6151
R891 B.n431 B.n430 10.6151
R892 B.n432 B.n431 10.6151
R893 B.n432 B.n85 10.6151
R894 B.n436 B.n85 10.6151
R895 B.n437 B.n436 10.6151
R896 B.n438 B.n437 10.6151
R897 B.n438 B.n83 10.6151
R898 B.n442 B.n83 10.6151
R899 B.n443 B.n442 10.6151
R900 B.n444 B.n443 10.6151
R901 B.n444 B.n81 10.6151
R902 B.n448 B.n81 10.6151
R903 B.n449 B.n448 10.6151
R904 B.n450 B.n449 10.6151
R905 B.n450 B.n79 10.6151
R906 B.n454 B.n79 10.6151
R907 B.n455 B.n454 10.6151
R908 B.n456 B.n455 10.6151
R909 B.n210 B.n209 10.6151
R910 B.n210 B.n163 10.6151
R911 B.n214 B.n163 10.6151
R912 B.n215 B.n214 10.6151
R913 B.n216 B.n215 10.6151
R914 B.n216 B.n161 10.6151
R915 B.n220 B.n161 10.6151
R916 B.n221 B.n220 10.6151
R917 B.n222 B.n221 10.6151
R918 B.n222 B.n159 10.6151
R919 B.n226 B.n159 10.6151
R920 B.n227 B.n226 10.6151
R921 B.n228 B.n227 10.6151
R922 B.n228 B.n157 10.6151
R923 B.n232 B.n157 10.6151
R924 B.n233 B.n232 10.6151
R925 B.n234 B.n233 10.6151
R926 B.n234 B.n155 10.6151
R927 B.n238 B.n155 10.6151
R928 B.n239 B.n238 10.6151
R929 B.n240 B.n239 10.6151
R930 B.n240 B.n153 10.6151
R931 B.n244 B.n153 10.6151
R932 B.n245 B.n244 10.6151
R933 B.n246 B.n245 10.6151
R934 B.n246 B.n151 10.6151
R935 B.n250 B.n151 10.6151
R936 B.n251 B.n250 10.6151
R937 B.n252 B.n251 10.6151
R938 B.n252 B.n149 10.6151
R939 B.n256 B.n149 10.6151
R940 B.n257 B.n256 10.6151
R941 B.n258 B.n257 10.6151
R942 B.n258 B.n147 10.6151
R943 B.n262 B.n147 10.6151
R944 B.n263 B.n262 10.6151
R945 B.n264 B.n263 10.6151
R946 B.n264 B.n145 10.6151
R947 B.n268 B.n145 10.6151
R948 B.n269 B.n268 10.6151
R949 B.n270 B.n269 10.6151
R950 B.n270 B.n143 10.6151
R951 B.n274 B.n143 10.6151
R952 B.n275 B.n274 10.6151
R953 B.n276 B.n275 10.6151
R954 B.n276 B.n141 10.6151
R955 B.n280 B.n141 10.6151
R956 B.n281 B.n280 10.6151
R957 B.n282 B.n281 10.6151
R958 B.n282 B.n139 10.6151
R959 B.n286 B.n139 10.6151
R960 B.n287 B.n286 10.6151
R961 B.n288 B.n287 10.6151
R962 B.n292 B.n291 10.6151
R963 B.n293 B.n292 10.6151
R964 B.n293 B.n133 10.6151
R965 B.n297 B.n133 10.6151
R966 B.n298 B.n297 10.6151
R967 B.n299 B.n298 10.6151
R968 B.n299 B.n131 10.6151
R969 B.n303 B.n131 10.6151
R970 B.n304 B.n303 10.6151
R971 B.n306 B.n127 10.6151
R972 B.n310 B.n127 10.6151
R973 B.n311 B.n310 10.6151
R974 B.n312 B.n311 10.6151
R975 B.n312 B.n125 10.6151
R976 B.n316 B.n125 10.6151
R977 B.n317 B.n316 10.6151
R978 B.n318 B.n317 10.6151
R979 B.n318 B.n123 10.6151
R980 B.n322 B.n123 10.6151
R981 B.n323 B.n322 10.6151
R982 B.n324 B.n323 10.6151
R983 B.n324 B.n121 10.6151
R984 B.n328 B.n121 10.6151
R985 B.n329 B.n328 10.6151
R986 B.n330 B.n329 10.6151
R987 B.n330 B.n119 10.6151
R988 B.n334 B.n119 10.6151
R989 B.n335 B.n334 10.6151
R990 B.n336 B.n335 10.6151
R991 B.n336 B.n117 10.6151
R992 B.n340 B.n117 10.6151
R993 B.n341 B.n340 10.6151
R994 B.n342 B.n341 10.6151
R995 B.n342 B.n115 10.6151
R996 B.n346 B.n115 10.6151
R997 B.n347 B.n346 10.6151
R998 B.n348 B.n347 10.6151
R999 B.n348 B.n113 10.6151
R1000 B.n352 B.n113 10.6151
R1001 B.n353 B.n352 10.6151
R1002 B.n354 B.n353 10.6151
R1003 B.n354 B.n111 10.6151
R1004 B.n358 B.n111 10.6151
R1005 B.n359 B.n358 10.6151
R1006 B.n360 B.n359 10.6151
R1007 B.n360 B.n109 10.6151
R1008 B.n364 B.n109 10.6151
R1009 B.n365 B.n364 10.6151
R1010 B.n366 B.n365 10.6151
R1011 B.n366 B.n107 10.6151
R1012 B.n370 B.n107 10.6151
R1013 B.n371 B.n370 10.6151
R1014 B.n372 B.n371 10.6151
R1015 B.n372 B.n105 10.6151
R1016 B.n376 B.n105 10.6151
R1017 B.n377 B.n376 10.6151
R1018 B.n378 B.n377 10.6151
R1019 B.n378 B.n103 10.6151
R1020 B.n382 B.n103 10.6151
R1021 B.n383 B.n382 10.6151
R1022 B.n384 B.n383 10.6151
R1023 B.n384 B.n101 10.6151
R1024 B.n208 B.n165 10.6151
R1025 B.n204 B.n165 10.6151
R1026 B.n204 B.n203 10.6151
R1027 B.n203 B.n202 10.6151
R1028 B.n202 B.n167 10.6151
R1029 B.n198 B.n167 10.6151
R1030 B.n198 B.n197 10.6151
R1031 B.n197 B.n196 10.6151
R1032 B.n196 B.n169 10.6151
R1033 B.n192 B.n169 10.6151
R1034 B.n192 B.n191 10.6151
R1035 B.n191 B.n190 10.6151
R1036 B.n190 B.n171 10.6151
R1037 B.n186 B.n171 10.6151
R1038 B.n186 B.n185 10.6151
R1039 B.n185 B.n184 10.6151
R1040 B.n184 B.n173 10.6151
R1041 B.n180 B.n173 10.6151
R1042 B.n180 B.n179 10.6151
R1043 B.n179 B.n178 10.6151
R1044 B.n178 B.n175 10.6151
R1045 B.n175 B.n0 10.6151
R1046 B.n667 B.n1 10.6151
R1047 B.n667 B.n666 10.6151
R1048 B.n666 B.n665 10.6151
R1049 B.n665 B.n4 10.6151
R1050 B.n661 B.n4 10.6151
R1051 B.n661 B.n660 10.6151
R1052 B.n660 B.n659 10.6151
R1053 B.n659 B.n6 10.6151
R1054 B.n655 B.n6 10.6151
R1055 B.n655 B.n654 10.6151
R1056 B.n654 B.n653 10.6151
R1057 B.n653 B.n8 10.6151
R1058 B.n649 B.n8 10.6151
R1059 B.n649 B.n648 10.6151
R1060 B.n648 B.n647 10.6151
R1061 B.n647 B.n10 10.6151
R1062 B.n643 B.n10 10.6151
R1063 B.n643 B.n642 10.6151
R1064 B.n642 B.n641 10.6151
R1065 B.n641 B.n12 10.6151
R1066 B.n637 B.n12 10.6151
R1067 B.n637 B.n636 10.6151
R1068 B.n44 B.n40 9.36635
R1069 B.n539 B.n538 9.36635
R1070 B.n288 B.n137 9.36635
R1071 B.n306 B.n305 9.36635
R1072 B.n671 B.n0 2.81026
R1073 B.n671 B.n1 2.81026
R1074 B.n553 B.n44 1.24928
R1075 B.n540 B.n539 1.24928
R1076 B.n291 B.n137 1.24928
R1077 B.n305 B.n304 1.24928
R1078 VP.n5 VP.t3 478.572
R1079 VP.n12 VP.t4 460.207
R1080 VP.n19 VP.t5 460.207
R1081 VP.n9 VP.t2 460.207
R1082 VP.n1 VP.t0 418.418
R1083 VP.n4 VP.t1 418.418
R1084 VP.n20 VP.n19 161.3
R1085 VP.n7 VP.n6 161.3
R1086 VP.n8 VP.n3 161.3
R1087 VP.n10 VP.n9 161.3
R1088 VP.n18 VP.n0 161.3
R1089 VP.n17 VP.n16 161.3
R1090 VP.n15 VP.n14 161.3
R1091 VP.n13 VP.n2 161.3
R1092 VP.n12 VP.n11 161.3
R1093 VP.n14 VP.n13 51.7179
R1094 VP.n18 VP.n17 51.7179
R1095 VP.n8 VP.n7 51.7179
R1096 VP.n11 VP.n10 45.4664
R1097 VP.n6 VP.n5 43.341
R1098 VP.n5 VP.n4 42.4561
R1099 VP.n14 VP.n1 12.2964
R1100 VP.n17 VP.n1 12.2964
R1101 VP.n7 VP.n4 12.2964
R1102 VP.n13 VP.n12 7.30353
R1103 VP.n19 VP.n18 7.30353
R1104 VP.n9 VP.n8 7.30353
R1105 VP.n6 VP.n3 0.189894
R1106 VP.n10 VP.n3 0.189894
R1107 VP.n11 VP.n2 0.189894
R1108 VP.n15 VP.n2 0.189894
R1109 VP.n16 VP.n15 0.189894
R1110 VP.n16 VP.n0 0.189894
R1111 VP.n20 VP.n0 0.189894
R1112 VP VP.n20 0.0516364
R1113 VDD1 VDD1.t2 70.1352
R1114 VDD1.n1 VDD1.t1 70.0214
R1115 VDD1.n1 VDD1.n0 67.4823
R1116 VDD1.n3 VDD1.n2 67.264
R1117 VDD1.n3 VDD1.n1 42.4729
R1118 VDD1.n2 VDD1.t4 1.99223
R1119 VDD1.n2 VDD1.t3 1.99223
R1120 VDD1.n0 VDD1.t5 1.99223
R1121 VDD1.n0 VDD1.t0 1.99223
R1122 VDD1 VDD1.n3 0.216017
C0 VDD2 VDD1 0.799095f
C1 VP VN 6.10871f
C2 VTAIL VDD1 11.4656f
C3 VP B 1.28128f
C4 VN VDD2 6.62499f
C5 w_n1986_n4232# VDD1 2.19022f
C6 VDD2 B 1.98672f
C7 VTAIL VN 6.20225f
C8 VTAIL B 3.66846f
C9 w_n1986_n4232# VN 3.43297f
C10 w_n1986_n4232# B 8.59558f
C11 VP VDD2 0.318765f
C12 VTAIL VP 6.21694f
C13 w_n1986_n4232# VP 3.6851f
C14 VTAIL VDD2 11.5f
C15 w_n1986_n4232# VDD2 2.22199f
C16 VN VDD1 0.148765f
C17 w_n1986_n4232# VTAIL 3.59891f
C18 VDD1 B 1.95211f
C19 VN B 0.868666f
C20 VP VDD1 6.78942f
C21 VDD2 VSUBS 1.579185f
C22 VDD1 VSUBS 1.918735f
C23 VTAIL VSUBS 0.966055f
C24 VN VSUBS 4.8427f
C25 VP VSUBS 1.812962f
C26 B VSUBS 3.363195f
C27 w_n1986_n4232# VSUBS 0.10293p
C28 VDD1.t2 VSUBS 3.47144f
C29 VDD1.t1 VSUBS 3.47026f
C30 VDD1.t5 VSUBS 0.326275f
C31 VDD1.t0 VSUBS 0.326275f
C32 VDD1.n0 VSUBS 2.66799f
C33 VDD1.n1 VSUBS 3.18091f
C34 VDD1.t4 VSUBS 0.326275f
C35 VDD1.t3 VSUBS 0.326275f
C36 VDD1.n2 VSUBS 2.66597f
C37 VDD1.n3 VSUBS 2.97988f
C38 VP.n0 VSUBS 0.048873f
C39 VP.t0 VSUBS 2.05823f
C40 VP.n1 VSUBS 0.745124f
C41 VP.n2 VSUBS 0.048873f
C42 VP.n3 VSUBS 0.048873f
C43 VP.t2 VSUBS 2.12818f
C44 VP.t1 VSUBS 2.05823f
C45 VP.n4 VSUBS 0.792393f
C46 VP.t3 VSUBS 2.15943f
C47 VP.n5 VSUBS 0.806257f
C48 VP.n6 VSUBS 0.20891f
C49 VP.n7 VSUBS 0.065443f
C50 VP.n8 VSUBS 0.016974f
C51 VP.n9 VSUBS 0.801313f
C52 VP.n10 VSUBS 2.29461f
C53 VP.n11 VSUBS 2.33336f
C54 VP.t4 VSUBS 2.12818f
C55 VP.n12 VSUBS 0.801313f
C56 VP.n13 VSUBS 0.016974f
C57 VP.n14 VSUBS 0.065443f
C58 VP.n15 VSUBS 0.048873f
C59 VP.n16 VSUBS 0.048873f
C60 VP.n17 VSUBS 0.065443f
C61 VP.n18 VSUBS 0.016974f
C62 VP.t5 VSUBS 2.12818f
C63 VP.n19 VSUBS 0.801313f
C64 VP.n20 VSUBS 0.037875f
C65 B.n0 VSUBS 0.004239f
C66 B.n1 VSUBS 0.004239f
C67 B.n2 VSUBS 0.006703f
C68 B.n3 VSUBS 0.006703f
C69 B.n4 VSUBS 0.006703f
C70 B.n5 VSUBS 0.006703f
C71 B.n6 VSUBS 0.006703f
C72 B.n7 VSUBS 0.006703f
C73 B.n8 VSUBS 0.006703f
C74 B.n9 VSUBS 0.006703f
C75 B.n10 VSUBS 0.006703f
C76 B.n11 VSUBS 0.006703f
C77 B.n12 VSUBS 0.006703f
C78 B.n13 VSUBS 0.015844f
C79 B.n14 VSUBS 0.006703f
C80 B.n15 VSUBS 0.006703f
C81 B.n16 VSUBS 0.006703f
C82 B.n17 VSUBS 0.006703f
C83 B.n18 VSUBS 0.006703f
C84 B.n19 VSUBS 0.006703f
C85 B.n20 VSUBS 0.006703f
C86 B.n21 VSUBS 0.006703f
C87 B.n22 VSUBS 0.006703f
C88 B.n23 VSUBS 0.006703f
C89 B.n24 VSUBS 0.006703f
C90 B.n25 VSUBS 0.006703f
C91 B.n26 VSUBS 0.006703f
C92 B.n27 VSUBS 0.006703f
C93 B.n28 VSUBS 0.006703f
C94 B.n29 VSUBS 0.006703f
C95 B.n30 VSUBS 0.006703f
C96 B.n31 VSUBS 0.006703f
C97 B.n32 VSUBS 0.006703f
C98 B.n33 VSUBS 0.006703f
C99 B.n34 VSUBS 0.006703f
C100 B.n35 VSUBS 0.006703f
C101 B.n36 VSUBS 0.006703f
C102 B.n37 VSUBS 0.006703f
C103 B.n38 VSUBS 0.006703f
C104 B.n39 VSUBS 0.006703f
C105 B.n40 VSUBS 0.006309f
C106 B.n41 VSUBS 0.006703f
C107 B.t8 VSUBS 0.523778f
C108 B.t7 VSUBS 0.533722f
C109 B.t6 VSUBS 0.607044f
C110 B.n42 VSUBS 0.188911f
C111 B.n43 VSUBS 0.062451f
C112 B.n44 VSUBS 0.015531f
C113 B.n45 VSUBS 0.006703f
C114 B.n46 VSUBS 0.006703f
C115 B.n47 VSUBS 0.006703f
C116 B.n48 VSUBS 0.006703f
C117 B.t2 VSUBS 0.52376f
C118 B.t1 VSUBS 0.533706f
C119 B.t0 VSUBS 0.607044f
C120 B.n49 VSUBS 0.188927f
C121 B.n50 VSUBS 0.062469f
C122 B.n51 VSUBS 0.006703f
C123 B.n52 VSUBS 0.006703f
C124 B.n53 VSUBS 0.006703f
C125 B.n54 VSUBS 0.006703f
C126 B.n55 VSUBS 0.006703f
C127 B.n56 VSUBS 0.006703f
C128 B.n57 VSUBS 0.006703f
C129 B.n58 VSUBS 0.006703f
C130 B.n59 VSUBS 0.006703f
C131 B.n60 VSUBS 0.006703f
C132 B.n61 VSUBS 0.006703f
C133 B.n62 VSUBS 0.006703f
C134 B.n63 VSUBS 0.006703f
C135 B.n64 VSUBS 0.006703f
C136 B.n65 VSUBS 0.006703f
C137 B.n66 VSUBS 0.006703f
C138 B.n67 VSUBS 0.006703f
C139 B.n68 VSUBS 0.006703f
C140 B.n69 VSUBS 0.006703f
C141 B.n70 VSUBS 0.006703f
C142 B.n71 VSUBS 0.006703f
C143 B.n72 VSUBS 0.006703f
C144 B.n73 VSUBS 0.006703f
C145 B.n74 VSUBS 0.006703f
C146 B.n75 VSUBS 0.006703f
C147 B.n76 VSUBS 0.006703f
C148 B.n77 VSUBS 0.015733f
C149 B.n78 VSUBS 0.006703f
C150 B.n79 VSUBS 0.006703f
C151 B.n80 VSUBS 0.006703f
C152 B.n81 VSUBS 0.006703f
C153 B.n82 VSUBS 0.006703f
C154 B.n83 VSUBS 0.006703f
C155 B.n84 VSUBS 0.006703f
C156 B.n85 VSUBS 0.006703f
C157 B.n86 VSUBS 0.006703f
C158 B.n87 VSUBS 0.006703f
C159 B.n88 VSUBS 0.006703f
C160 B.n89 VSUBS 0.006703f
C161 B.n90 VSUBS 0.006703f
C162 B.n91 VSUBS 0.006703f
C163 B.n92 VSUBS 0.006703f
C164 B.n93 VSUBS 0.006703f
C165 B.n94 VSUBS 0.006703f
C166 B.n95 VSUBS 0.006703f
C167 B.n96 VSUBS 0.006703f
C168 B.n97 VSUBS 0.006703f
C169 B.n98 VSUBS 0.006703f
C170 B.n99 VSUBS 0.006703f
C171 B.n100 VSUBS 0.006703f
C172 B.n101 VSUBS 0.01649f
C173 B.n102 VSUBS 0.006703f
C174 B.n103 VSUBS 0.006703f
C175 B.n104 VSUBS 0.006703f
C176 B.n105 VSUBS 0.006703f
C177 B.n106 VSUBS 0.006703f
C178 B.n107 VSUBS 0.006703f
C179 B.n108 VSUBS 0.006703f
C180 B.n109 VSUBS 0.006703f
C181 B.n110 VSUBS 0.006703f
C182 B.n111 VSUBS 0.006703f
C183 B.n112 VSUBS 0.006703f
C184 B.n113 VSUBS 0.006703f
C185 B.n114 VSUBS 0.006703f
C186 B.n115 VSUBS 0.006703f
C187 B.n116 VSUBS 0.006703f
C188 B.n117 VSUBS 0.006703f
C189 B.n118 VSUBS 0.006703f
C190 B.n119 VSUBS 0.006703f
C191 B.n120 VSUBS 0.006703f
C192 B.n121 VSUBS 0.006703f
C193 B.n122 VSUBS 0.006703f
C194 B.n123 VSUBS 0.006703f
C195 B.n124 VSUBS 0.006703f
C196 B.n125 VSUBS 0.006703f
C197 B.n126 VSUBS 0.006703f
C198 B.n127 VSUBS 0.006703f
C199 B.n128 VSUBS 0.006703f
C200 B.t4 VSUBS 0.52376f
C201 B.t5 VSUBS 0.533706f
C202 B.t3 VSUBS 0.607044f
C203 B.n129 VSUBS 0.188927f
C204 B.n130 VSUBS 0.062469f
C205 B.n131 VSUBS 0.006703f
C206 B.n132 VSUBS 0.006703f
C207 B.n133 VSUBS 0.006703f
C208 B.n134 VSUBS 0.006703f
C209 B.t10 VSUBS 0.523778f
C210 B.t11 VSUBS 0.533722f
C211 B.t9 VSUBS 0.607044f
C212 B.n135 VSUBS 0.188911f
C213 B.n136 VSUBS 0.062451f
C214 B.n137 VSUBS 0.015531f
C215 B.n138 VSUBS 0.006703f
C216 B.n139 VSUBS 0.006703f
C217 B.n140 VSUBS 0.006703f
C218 B.n141 VSUBS 0.006703f
C219 B.n142 VSUBS 0.006703f
C220 B.n143 VSUBS 0.006703f
C221 B.n144 VSUBS 0.006703f
C222 B.n145 VSUBS 0.006703f
C223 B.n146 VSUBS 0.006703f
C224 B.n147 VSUBS 0.006703f
C225 B.n148 VSUBS 0.006703f
C226 B.n149 VSUBS 0.006703f
C227 B.n150 VSUBS 0.006703f
C228 B.n151 VSUBS 0.006703f
C229 B.n152 VSUBS 0.006703f
C230 B.n153 VSUBS 0.006703f
C231 B.n154 VSUBS 0.006703f
C232 B.n155 VSUBS 0.006703f
C233 B.n156 VSUBS 0.006703f
C234 B.n157 VSUBS 0.006703f
C235 B.n158 VSUBS 0.006703f
C236 B.n159 VSUBS 0.006703f
C237 B.n160 VSUBS 0.006703f
C238 B.n161 VSUBS 0.006703f
C239 B.n162 VSUBS 0.006703f
C240 B.n163 VSUBS 0.006703f
C241 B.n164 VSUBS 0.01649f
C242 B.n165 VSUBS 0.006703f
C243 B.n166 VSUBS 0.006703f
C244 B.n167 VSUBS 0.006703f
C245 B.n168 VSUBS 0.006703f
C246 B.n169 VSUBS 0.006703f
C247 B.n170 VSUBS 0.006703f
C248 B.n171 VSUBS 0.006703f
C249 B.n172 VSUBS 0.006703f
C250 B.n173 VSUBS 0.006703f
C251 B.n174 VSUBS 0.006703f
C252 B.n175 VSUBS 0.006703f
C253 B.n176 VSUBS 0.006703f
C254 B.n177 VSUBS 0.006703f
C255 B.n178 VSUBS 0.006703f
C256 B.n179 VSUBS 0.006703f
C257 B.n180 VSUBS 0.006703f
C258 B.n181 VSUBS 0.006703f
C259 B.n182 VSUBS 0.006703f
C260 B.n183 VSUBS 0.006703f
C261 B.n184 VSUBS 0.006703f
C262 B.n185 VSUBS 0.006703f
C263 B.n186 VSUBS 0.006703f
C264 B.n187 VSUBS 0.006703f
C265 B.n188 VSUBS 0.006703f
C266 B.n189 VSUBS 0.006703f
C267 B.n190 VSUBS 0.006703f
C268 B.n191 VSUBS 0.006703f
C269 B.n192 VSUBS 0.006703f
C270 B.n193 VSUBS 0.006703f
C271 B.n194 VSUBS 0.006703f
C272 B.n195 VSUBS 0.006703f
C273 B.n196 VSUBS 0.006703f
C274 B.n197 VSUBS 0.006703f
C275 B.n198 VSUBS 0.006703f
C276 B.n199 VSUBS 0.006703f
C277 B.n200 VSUBS 0.006703f
C278 B.n201 VSUBS 0.006703f
C279 B.n202 VSUBS 0.006703f
C280 B.n203 VSUBS 0.006703f
C281 B.n204 VSUBS 0.006703f
C282 B.n205 VSUBS 0.006703f
C283 B.n206 VSUBS 0.006703f
C284 B.n207 VSUBS 0.015844f
C285 B.n208 VSUBS 0.015844f
C286 B.n209 VSUBS 0.01649f
C287 B.n210 VSUBS 0.006703f
C288 B.n211 VSUBS 0.006703f
C289 B.n212 VSUBS 0.006703f
C290 B.n213 VSUBS 0.006703f
C291 B.n214 VSUBS 0.006703f
C292 B.n215 VSUBS 0.006703f
C293 B.n216 VSUBS 0.006703f
C294 B.n217 VSUBS 0.006703f
C295 B.n218 VSUBS 0.006703f
C296 B.n219 VSUBS 0.006703f
C297 B.n220 VSUBS 0.006703f
C298 B.n221 VSUBS 0.006703f
C299 B.n222 VSUBS 0.006703f
C300 B.n223 VSUBS 0.006703f
C301 B.n224 VSUBS 0.006703f
C302 B.n225 VSUBS 0.006703f
C303 B.n226 VSUBS 0.006703f
C304 B.n227 VSUBS 0.006703f
C305 B.n228 VSUBS 0.006703f
C306 B.n229 VSUBS 0.006703f
C307 B.n230 VSUBS 0.006703f
C308 B.n231 VSUBS 0.006703f
C309 B.n232 VSUBS 0.006703f
C310 B.n233 VSUBS 0.006703f
C311 B.n234 VSUBS 0.006703f
C312 B.n235 VSUBS 0.006703f
C313 B.n236 VSUBS 0.006703f
C314 B.n237 VSUBS 0.006703f
C315 B.n238 VSUBS 0.006703f
C316 B.n239 VSUBS 0.006703f
C317 B.n240 VSUBS 0.006703f
C318 B.n241 VSUBS 0.006703f
C319 B.n242 VSUBS 0.006703f
C320 B.n243 VSUBS 0.006703f
C321 B.n244 VSUBS 0.006703f
C322 B.n245 VSUBS 0.006703f
C323 B.n246 VSUBS 0.006703f
C324 B.n247 VSUBS 0.006703f
C325 B.n248 VSUBS 0.006703f
C326 B.n249 VSUBS 0.006703f
C327 B.n250 VSUBS 0.006703f
C328 B.n251 VSUBS 0.006703f
C329 B.n252 VSUBS 0.006703f
C330 B.n253 VSUBS 0.006703f
C331 B.n254 VSUBS 0.006703f
C332 B.n255 VSUBS 0.006703f
C333 B.n256 VSUBS 0.006703f
C334 B.n257 VSUBS 0.006703f
C335 B.n258 VSUBS 0.006703f
C336 B.n259 VSUBS 0.006703f
C337 B.n260 VSUBS 0.006703f
C338 B.n261 VSUBS 0.006703f
C339 B.n262 VSUBS 0.006703f
C340 B.n263 VSUBS 0.006703f
C341 B.n264 VSUBS 0.006703f
C342 B.n265 VSUBS 0.006703f
C343 B.n266 VSUBS 0.006703f
C344 B.n267 VSUBS 0.006703f
C345 B.n268 VSUBS 0.006703f
C346 B.n269 VSUBS 0.006703f
C347 B.n270 VSUBS 0.006703f
C348 B.n271 VSUBS 0.006703f
C349 B.n272 VSUBS 0.006703f
C350 B.n273 VSUBS 0.006703f
C351 B.n274 VSUBS 0.006703f
C352 B.n275 VSUBS 0.006703f
C353 B.n276 VSUBS 0.006703f
C354 B.n277 VSUBS 0.006703f
C355 B.n278 VSUBS 0.006703f
C356 B.n279 VSUBS 0.006703f
C357 B.n280 VSUBS 0.006703f
C358 B.n281 VSUBS 0.006703f
C359 B.n282 VSUBS 0.006703f
C360 B.n283 VSUBS 0.006703f
C361 B.n284 VSUBS 0.006703f
C362 B.n285 VSUBS 0.006703f
C363 B.n286 VSUBS 0.006703f
C364 B.n287 VSUBS 0.006703f
C365 B.n288 VSUBS 0.006309f
C366 B.n289 VSUBS 0.006703f
C367 B.n290 VSUBS 0.006703f
C368 B.n291 VSUBS 0.003746f
C369 B.n292 VSUBS 0.006703f
C370 B.n293 VSUBS 0.006703f
C371 B.n294 VSUBS 0.006703f
C372 B.n295 VSUBS 0.006703f
C373 B.n296 VSUBS 0.006703f
C374 B.n297 VSUBS 0.006703f
C375 B.n298 VSUBS 0.006703f
C376 B.n299 VSUBS 0.006703f
C377 B.n300 VSUBS 0.006703f
C378 B.n301 VSUBS 0.006703f
C379 B.n302 VSUBS 0.006703f
C380 B.n303 VSUBS 0.006703f
C381 B.n304 VSUBS 0.003746f
C382 B.n305 VSUBS 0.015531f
C383 B.n306 VSUBS 0.006309f
C384 B.n307 VSUBS 0.006703f
C385 B.n308 VSUBS 0.006703f
C386 B.n309 VSUBS 0.006703f
C387 B.n310 VSUBS 0.006703f
C388 B.n311 VSUBS 0.006703f
C389 B.n312 VSUBS 0.006703f
C390 B.n313 VSUBS 0.006703f
C391 B.n314 VSUBS 0.006703f
C392 B.n315 VSUBS 0.006703f
C393 B.n316 VSUBS 0.006703f
C394 B.n317 VSUBS 0.006703f
C395 B.n318 VSUBS 0.006703f
C396 B.n319 VSUBS 0.006703f
C397 B.n320 VSUBS 0.006703f
C398 B.n321 VSUBS 0.006703f
C399 B.n322 VSUBS 0.006703f
C400 B.n323 VSUBS 0.006703f
C401 B.n324 VSUBS 0.006703f
C402 B.n325 VSUBS 0.006703f
C403 B.n326 VSUBS 0.006703f
C404 B.n327 VSUBS 0.006703f
C405 B.n328 VSUBS 0.006703f
C406 B.n329 VSUBS 0.006703f
C407 B.n330 VSUBS 0.006703f
C408 B.n331 VSUBS 0.006703f
C409 B.n332 VSUBS 0.006703f
C410 B.n333 VSUBS 0.006703f
C411 B.n334 VSUBS 0.006703f
C412 B.n335 VSUBS 0.006703f
C413 B.n336 VSUBS 0.006703f
C414 B.n337 VSUBS 0.006703f
C415 B.n338 VSUBS 0.006703f
C416 B.n339 VSUBS 0.006703f
C417 B.n340 VSUBS 0.006703f
C418 B.n341 VSUBS 0.006703f
C419 B.n342 VSUBS 0.006703f
C420 B.n343 VSUBS 0.006703f
C421 B.n344 VSUBS 0.006703f
C422 B.n345 VSUBS 0.006703f
C423 B.n346 VSUBS 0.006703f
C424 B.n347 VSUBS 0.006703f
C425 B.n348 VSUBS 0.006703f
C426 B.n349 VSUBS 0.006703f
C427 B.n350 VSUBS 0.006703f
C428 B.n351 VSUBS 0.006703f
C429 B.n352 VSUBS 0.006703f
C430 B.n353 VSUBS 0.006703f
C431 B.n354 VSUBS 0.006703f
C432 B.n355 VSUBS 0.006703f
C433 B.n356 VSUBS 0.006703f
C434 B.n357 VSUBS 0.006703f
C435 B.n358 VSUBS 0.006703f
C436 B.n359 VSUBS 0.006703f
C437 B.n360 VSUBS 0.006703f
C438 B.n361 VSUBS 0.006703f
C439 B.n362 VSUBS 0.006703f
C440 B.n363 VSUBS 0.006703f
C441 B.n364 VSUBS 0.006703f
C442 B.n365 VSUBS 0.006703f
C443 B.n366 VSUBS 0.006703f
C444 B.n367 VSUBS 0.006703f
C445 B.n368 VSUBS 0.006703f
C446 B.n369 VSUBS 0.006703f
C447 B.n370 VSUBS 0.006703f
C448 B.n371 VSUBS 0.006703f
C449 B.n372 VSUBS 0.006703f
C450 B.n373 VSUBS 0.006703f
C451 B.n374 VSUBS 0.006703f
C452 B.n375 VSUBS 0.006703f
C453 B.n376 VSUBS 0.006703f
C454 B.n377 VSUBS 0.006703f
C455 B.n378 VSUBS 0.006703f
C456 B.n379 VSUBS 0.006703f
C457 B.n380 VSUBS 0.006703f
C458 B.n381 VSUBS 0.006703f
C459 B.n382 VSUBS 0.006703f
C460 B.n383 VSUBS 0.006703f
C461 B.n384 VSUBS 0.006703f
C462 B.n385 VSUBS 0.006703f
C463 B.n386 VSUBS 0.01649f
C464 B.n387 VSUBS 0.015844f
C465 B.n388 VSUBS 0.015844f
C466 B.n389 VSUBS 0.006703f
C467 B.n390 VSUBS 0.006703f
C468 B.n391 VSUBS 0.006703f
C469 B.n392 VSUBS 0.006703f
C470 B.n393 VSUBS 0.006703f
C471 B.n394 VSUBS 0.006703f
C472 B.n395 VSUBS 0.006703f
C473 B.n396 VSUBS 0.006703f
C474 B.n397 VSUBS 0.006703f
C475 B.n398 VSUBS 0.006703f
C476 B.n399 VSUBS 0.006703f
C477 B.n400 VSUBS 0.006703f
C478 B.n401 VSUBS 0.006703f
C479 B.n402 VSUBS 0.006703f
C480 B.n403 VSUBS 0.006703f
C481 B.n404 VSUBS 0.006703f
C482 B.n405 VSUBS 0.006703f
C483 B.n406 VSUBS 0.006703f
C484 B.n407 VSUBS 0.006703f
C485 B.n408 VSUBS 0.006703f
C486 B.n409 VSUBS 0.006703f
C487 B.n410 VSUBS 0.006703f
C488 B.n411 VSUBS 0.006703f
C489 B.n412 VSUBS 0.006703f
C490 B.n413 VSUBS 0.006703f
C491 B.n414 VSUBS 0.006703f
C492 B.n415 VSUBS 0.006703f
C493 B.n416 VSUBS 0.006703f
C494 B.n417 VSUBS 0.006703f
C495 B.n418 VSUBS 0.006703f
C496 B.n419 VSUBS 0.006703f
C497 B.n420 VSUBS 0.006703f
C498 B.n421 VSUBS 0.006703f
C499 B.n422 VSUBS 0.006703f
C500 B.n423 VSUBS 0.006703f
C501 B.n424 VSUBS 0.006703f
C502 B.n425 VSUBS 0.006703f
C503 B.n426 VSUBS 0.006703f
C504 B.n427 VSUBS 0.006703f
C505 B.n428 VSUBS 0.006703f
C506 B.n429 VSUBS 0.006703f
C507 B.n430 VSUBS 0.006703f
C508 B.n431 VSUBS 0.006703f
C509 B.n432 VSUBS 0.006703f
C510 B.n433 VSUBS 0.006703f
C511 B.n434 VSUBS 0.006703f
C512 B.n435 VSUBS 0.006703f
C513 B.n436 VSUBS 0.006703f
C514 B.n437 VSUBS 0.006703f
C515 B.n438 VSUBS 0.006703f
C516 B.n439 VSUBS 0.006703f
C517 B.n440 VSUBS 0.006703f
C518 B.n441 VSUBS 0.006703f
C519 B.n442 VSUBS 0.006703f
C520 B.n443 VSUBS 0.006703f
C521 B.n444 VSUBS 0.006703f
C522 B.n445 VSUBS 0.006703f
C523 B.n446 VSUBS 0.006703f
C524 B.n447 VSUBS 0.006703f
C525 B.n448 VSUBS 0.006703f
C526 B.n449 VSUBS 0.006703f
C527 B.n450 VSUBS 0.006703f
C528 B.n451 VSUBS 0.006703f
C529 B.n452 VSUBS 0.006703f
C530 B.n453 VSUBS 0.006703f
C531 B.n454 VSUBS 0.006703f
C532 B.n455 VSUBS 0.006703f
C533 B.n456 VSUBS 0.016601f
C534 B.n457 VSUBS 0.015844f
C535 B.n458 VSUBS 0.01649f
C536 B.n459 VSUBS 0.006703f
C537 B.n460 VSUBS 0.006703f
C538 B.n461 VSUBS 0.006703f
C539 B.n462 VSUBS 0.006703f
C540 B.n463 VSUBS 0.006703f
C541 B.n464 VSUBS 0.006703f
C542 B.n465 VSUBS 0.006703f
C543 B.n466 VSUBS 0.006703f
C544 B.n467 VSUBS 0.006703f
C545 B.n468 VSUBS 0.006703f
C546 B.n469 VSUBS 0.006703f
C547 B.n470 VSUBS 0.006703f
C548 B.n471 VSUBS 0.006703f
C549 B.n472 VSUBS 0.006703f
C550 B.n473 VSUBS 0.006703f
C551 B.n474 VSUBS 0.006703f
C552 B.n475 VSUBS 0.006703f
C553 B.n476 VSUBS 0.006703f
C554 B.n477 VSUBS 0.006703f
C555 B.n478 VSUBS 0.006703f
C556 B.n479 VSUBS 0.006703f
C557 B.n480 VSUBS 0.006703f
C558 B.n481 VSUBS 0.006703f
C559 B.n482 VSUBS 0.006703f
C560 B.n483 VSUBS 0.006703f
C561 B.n484 VSUBS 0.006703f
C562 B.n485 VSUBS 0.006703f
C563 B.n486 VSUBS 0.006703f
C564 B.n487 VSUBS 0.006703f
C565 B.n488 VSUBS 0.006703f
C566 B.n489 VSUBS 0.006703f
C567 B.n490 VSUBS 0.006703f
C568 B.n491 VSUBS 0.006703f
C569 B.n492 VSUBS 0.006703f
C570 B.n493 VSUBS 0.006703f
C571 B.n494 VSUBS 0.006703f
C572 B.n495 VSUBS 0.006703f
C573 B.n496 VSUBS 0.006703f
C574 B.n497 VSUBS 0.006703f
C575 B.n498 VSUBS 0.006703f
C576 B.n499 VSUBS 0.006703f
C577 B.n500 VSUBS 0.006703f
C578 B.n501 VSUBS 0.006703f
C579 B.n502 VSUBS 0.006703f
C580 B.n503 VSUBS 0.006703f
C581 B.n504 VSUBS 0.006703f
C582 B.n505 VSUBS 0.006703f
C583 B.n506 VSUBS 0.006703f
C584 B.n507 VSUBS 0.006703f
C585 B.n508 VSUBS 0.006703f
C586 B.n509 VSUBS 0.006703f
C587 B.n510 VSUBS 0.006703f
C588 B.n511 VSUBS 0.006703f
C589 B.n512 VSUBS 0.006703f
C590 B.n513 VSUBS 0.006703f
C591 B.n514 VSUBS 0.006703f
C592 B.n515 VSUBS 0.006703f
C593 B.n516 VSUBS 0.006703f
C594 B.n517 VSUBS 0.006703f
C595 B.n518 VSUBS 0.006703f
C596 B.n519 VSUBS 0.006703f
C597 B.n520 VSUBS 0.006703f
C598 B.n521 VSUBS 0.006703f
C599 B.n522 VSUBS 0.006703f
C600 B.n523 VSUBS 0.006703f
C601 B.n524 VSUBS 0.006703f
C602 B.n525 VSUBS 0.006703f
C603 B.n526 VSUBS 0.006703f
C604 B.n527 VSUBS 0.006703f
C605 B.n528 VSUBS 0.006703f
C606 B.n529 VSUBS 0.006703f
C607 B.n530 VSUBS 0.006703f
C608 B.n531 VSUBS 0.006703f
C609 B.n532 VSUBS 0.006703f
C610 B.n533 VSUBS 0.006703f
C611 B.n534 VSUBS 0.006703f
C612 B.n535 VSUBS 0.006703f
C613 B.n536 VSUBS 0.006703f
C614 B.n537 VSUBS 0.006703f
C615 B.n538 VSUBS 0.006309f
C616 B.n539 VSUBS 0.015531f
C617 B.n540 VSUBS 0.003746f
C618 B.n541 VSUBS 0.006703f
C619 B.n542 VSUBS 0.006703f
C620 B.n543 VSUBS 0.006703f
C621 B.n544 VSUBS 0.006703f
C622 B.n545 VSUBS 0.006703f
C623 B.n546 VSUBS 0.006703f
C624 B.n547 VSUBS 0.006703f
C625 B.n548 VSUBS 0.006703f
C626 B.n549 VSUBS 0.006703f
C627 B.n550 VSUBS 0.006703f
C628 B.n551 VSUBS 0.006703f
C629 B.n552 VSUBS 0.006703f
C630 B.n553 VSUBS 0.003746f
C631 B.n554 VSUBS 0.006703f
C632 B.n555 VSUBS 0.006703f
C633 B.n556 VSUBS 0.006703f
C634 B.n557 VSUBS 0.006703f
C635 B.n558 VSUBS 0.006703f
C636 B.n559 VSUBS 0.006703f
C637 B.n560 VSUBS 0.006703f
C638 B.n561 VSUBS 0.006703f
C639 B.n562 VSUBS 0.006703f
C640 B.n563 VSUBS 0.006703f
C641 B.n564 VSUBS 0.006703f
C642 B.n565 VSUBS 0.006703f
C643 B.n566 VSUBS 0.006703f
C644 B.n567 VSUBS 0.006703f
C645 B.n568 VSUBS 0.006703f
C646 B.n569 VSUBS 0.006703f
C647 B.n570 VSUBS 0.006703f
C648 B.n571 VSUBS 0.006703f
C649 B.n572 VSUBS 0.006703f
C650 B.n573 VSUBS 0.006703f
C651 B.n574 VSUBS 0.006703f
C652 B.n575 VSUBS 0.006703f
C653 B.n576 VSUBS 0.006703f
C654 B.n577 VSUBS 0.006703f
C655 B.n578 VSUBS 0.006703f
C656 B.n579 VSUBS 0.006703f
C657 B.n580 VSUBS 0.006703f
C658 B.n581 VSUBS 0.006703f
C659 B.n582 VSUBS 0.006703f
C660 B.n583 VSUBS 0.006703f
C661 B.n584 VSUBS 0.006703f
C662 B.n585 VSUBS 0.006703f
C663 B.n586 VSUBS 0.006703f
C664 B.n587 VSUBS 0.006703f
C665 B.n588 VSUBS 0.006703f
C666 B.n589 VSUBS 0.006703f
C667 B.n590 VSUBS 0.006703f
C668 B.n591 VSUBS 0.006703f
C669 B.n592 VSUBS 0.006703f
C670 B.n593 VSUBS 0.006703f
C671 B.n594 VSUBS 0.006703f
C672 B.n595 VSUBS 0.006703f
C673 B.n596 VSUBS 0.006703f
C674 B.n597 VSUBS 0.006703f
C675 B.n598 VSUBS 0.006703f
C676 B.n599 VSUBS 0.006703f
C677 B.n600 VSUBS 0.006703f
C678 B.n601 VSUBS 0.006703f
C679 B.n602 VSUBS 0.006703f
C680 B.n603 VSUBS 0.006703f
C681 B.n604 VSUBS 0.006703f
C682 B.n605 VSUBS 0.006703f
C683 B.n606 VSUBS 0.006703f
C684 B.n607 VSUBS 0.006703f
C685 B.n608 VSUBS 0.006703f
C686 B.n609 VSUBS 0.006703f
C687 B.n610 VSUBS 0.006703f
C688 B.n611 VSUBS 0.006703f
C689 B.n612 VSUBS 0.006703f
C690 B.n613 VSUBS 0.006703f
C691 B.n614 VSUBS 0.006703f
C692 B.n615 VSUBS 0.006703f
C693 B.n616 VSUBS 0.006703f
C694 B.n617 VSUBS 0.006703f
C695 B.n618 VSUBS 0.006703f
C696 B.n619 VSUBS 0.006703f
C697 B.n620 VSUBS 0.006703f
C698 B.n621 VSUBS 0.006703f
C699 B.n622 VSUBS 0.006703f
C700 B.n623 VSUBS 0.006703f
C701 B.n624 VSUBS 0.006703f
C702 B.n625 VSUBS 0.006703f
C703 B.n626 VSUBS 0.006703f
C704 B.n627 VSUBS 0.006703f
C705 B.n628 VSUBS 0.006703f
C706 B.n629 VSUBS 0.006703f
C707 B.n630 VSUBS 0.006703f
C708 B.n631 VSUBS 0.006703f
C709 B.n632 VSUBS 0.006703f
C710 B.n633 VSUBS 0.006703f
C711 B.n634 VSUBS 0.01649f
C712 B.n635 VSUBS 0.01649f
C713 B.n636 VSUBS 0.015844f
C714 B.n637 VSUBS 0.006703f
C715 B.n638 VSUBS 0.006703f
C716 B.n639 VSUBS 0.006703f
C717 B.n640 VSUBS 0.006703f
C718 B.n641 VSUBS 0.006703f
C719 B.n642 VSUBS 0.006703f
C720 B.n643 VSUBS 0.006703f
C721 B.n644 VSUBS 0.006703f
C722 B.n645 VSUBS 0.006703f
C723 B.n646 VSUBS 0.006703f
C724 B.n647 VSUBS 0.006703f
C725 B.n648 VSUBS 0.006703f
C726 B.n649 VSUBS 0.006703f
C727 B.n650 VSUBS 0.006703f
C728 B.n651 VSUBS 0.006703f
C729 B.n652 VSUBS 0.006703f
C730 B.n653 VSUBS 0.006703f
C731 B.n654 VSUBS 0.006703f
C732 B.n655 VSUBS 0.006703f
C733 B.n656 VSUBS 0.006703f
C734 B.n657 VSUBS 0.006703f
C735 B.n658 VSUBS 0.006703f
C736 B.n659 VSUBS 0.006703f
C737 B.n660 VSUBS 0.006703f
C738 B.n661 VSUBS 0.006703f
C739 B.n662 VSUBS 0.006703f
C740 B.n663 VSUBS 0.006703f
C741 B.n664 VSUBS 0.006703f
C742 B.n665 VSUBS 0.006703f
C743 B.n666 VSUBS 0.006703f
C744 B.n667 VSUBS 0.006703f
C745 B.n668 VSUBS 0.006703f
C746 B.n669 VSUBS 0.006703f
C747 B.n670 VSUBS 0.006703f
C748 B.n671 VSUBS 0.015179f
C749 VDD2.t5 VSUBS 3.45213f
C750 VDD2.t4 VSUBS 0.324571f
C751 VDD2.t0 VSUBS 0.324571f
C752 VDD2.n0 VSUBS 2.65406f
C753 VDD2.n1 VSUBS 3.07951f
C754 VDD2.t2 VSUBS 3.44486f
C755 VDD2.n2 VSUBS 3.01359f
C756 VDD2.t3 VSUBS 0.324571f
C757 VDD2.t1 VSUBS 0.324571f
C758 VDD2.n3 VSUBS 2.65402f
C759 VTAIL.t8 VSUBS 0.359169f
C760 VTAIL.t7 VSUBS 0.359169f
C761 VTAIL.n0 VSUBS 2.75395f
C762 VTAIL.n1 VSUBS 0.817681f
C763 VTAIL.t5 VSUBS 3.60567f
C764 VTAIL.n2 VSUBS 1.01397f
C765 VTAIL.t3 VSUBS 0.359169f
C766 VTAIL.t1 VSUBS 0.359169f
C767 VTAIL.n3 VSUBS 2.75395f
C768 VTAIL.n4 VSUBS 2.6322f
C769 VTAIL.t11 VSUBS 0.359169f
C770 VTAIL.t10 VSUBS 0.359169f
C771 VTAIL.n5 VSUBS 2.75395f
C772 VTAIL.n6 VSUBS 2.63219f
C773 VTAIL.t9 VSUBS 3.60568f
C774 VTAIL.n7 VSUBS 1.01397f
C775 VTAIL.t2 VSUBS 0.359169f
C776 VTAIL.t0 VSUBS 0.359169f
C777 VTAIL.n8 VSUBS 2.75395f
C778 VTAIL.n9 VSUBS 0.88614f
C779 VTAIL.t4 VSUBS 3.60567f
C780 VTAIL.n10 VSUBS 2.66178f
C781 VTAIL.t6 VSUBS 3.60567f
C782 VTAIL.n11 VSUBS 2.63199f
C783 VN.n0 VSUBS 0.047658f
C784 VN.t1 VSUBS 2.00705f
C785 VN.n1 VSUBS 0.772687f
C786 VN.t0 VSUBS 2.10573f
C787 VN.n2 VSUBS 0.786207f
C788 VN.n3 VSUBS 0.203715f
C789 VN.n4 VSUBS 0.063816f
C790 VN.n5 VSUBS 0.016552f
C791 VN.t5 VSUBS 2.07526f
C792 VN.n6 VSUBS 0.781386f
C793 VN.n7 VSUBS 0.036933f
C794 VN.n8 VSUBS 0.047658f
C795 VN.t2 VSUBS 2.00705f
C796 VN.n9 VSUBS 0.772687f
C797 VN.t4 VSUBS 2.10573f
C798 VN.n10 VSUBS 0.786207f
C799 VN.n11 VSUBS 0.203715f
C800 VN.n12 VSUBS 0.063816f
C801 VN.n13 VSUBS 0.016552f
C802 VN.t3 VSUBS 2.07526f
C803 VN.n14 VSUBS 0.781386f
C804 VN.n15 VSUBS 2.26869f
.ends

