* NGSPICE file created from diff_pair_sample_0599.ext - technology: sky130A

.subckt diff_pair_sample_0599 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=3.77
X1 VTAIL.t19 VP.t0 VDD1.t6 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X2 B.t8 B.t6 B.t7 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=3.77
X3 VTAIL.t18 VP.t1 VDD1.t5 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X4 B.t5 B.t3 B.t4 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=3.77
X5 B.t2 B.t0 B.t1 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=3.77
X6 VDD2.t9 VN.t0 VTAIL.t4 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=3.77
X7 VDD2.t8 VN.t1 VTAIL.t1 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=3.77
X8 VTAIL.t3 VN.t2 VDD2.t7 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X9 VDD1.t3 VP.t2 VTAIL.t17 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=3.77
X10 VTAIL.t5 VN.t3 VDD2.t6 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X11 VDD1.t0 VP.t3 VTAIL.t16 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X12 VDD2.t5 VN.t4 VTAIL.t7 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=3.77
X13 VTAIL.t15 VP.t4 VDD1.t4 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X14 VDD1.t1 VP.t5 VTAIL.t14 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=3.77
X15 VDD2.t4 VN.t5 VTAIL.t8 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=3.77
X16 VDD2.t3 VN.t6 VTAIL.t0 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X17 VDD1.t2 VP.t6 VTAIL.t13 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=3.77
X18 VDD2.t2 VN.t7 VTAIL.t9 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X19 VDD1.t9 VP.t7 VTAIL.t12 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X20 VTAIL.t2 VN.t8 VDD2.t1 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X21 VTAIL.t6 VN.t9 VDD2.t0 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
X22 VDD1.t7 VP.t8 VTAIL.t11 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=3.77
X23 VTAIL.t10 VP.t9 VDD1.t8 w_n5890_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=3.77
R0 B.n388 B.n147 585
R1 B.n387 B.n386 585
R2 B.n385 B.n148 585
R3 B.n384 B.n383 585
R4 B.n382 B.n149 585
R5 B.n381 B.n380 585
R6 B.n379 B.n150 585
R7 B.n378 B.n377 585
R8 B.n376 B.n151 585
R9 B.n375 B.n374 585
R10 B.n373 B.n152 585
R11 B.n372 B.n371 585
R12 B.n370 B.n153 585
R13 B.n369 B.n368 585
R14 B.n367 B.n154 585
R15 B.n366 B.n365 585
R16 B.n361 B.n155 585
R17 B.n360 B.n359 585
R18 B.n358 B.n156 585
R19 B.n357 B.n356 585
R20 B.n355 B.n157 585
R21 B.n354 B.n353 585
R22 B.n352 B.n158 585
R23 B.n351 B.n350 585
R24 B.n348 B.n159 585
R25 B.n347 B.n346 585
R26 B.n345 B.n162 585
R27 B.n344 B.n343 585
R28 B.n342 B.n163 585
R29 B.n341 B.n340 585
R30 B.n339 B.n164 585
R31 B.n338 B.n337 585
R32 B.n336 B.n165 585
R33 B.n335 B.n334 585
R34 B.n333 B.n166 585
R35 B.n332 B.n331 585
R36 B.n330 B.n167 585
R37 B.n329 B.n328 585
R38 B.n327 B.n168 585
R39 B.n390 B.n389 585
R40 B.n391 B.n146 585
R41 B.n393 B.n392 585
R42 B.n394 B.n145 585
R43 B.n396 B.n395 585
R44 B.n397 B.n144 585
R45 B.n399 B.n398 585
R46 B.n400 B.n143 585
R47 B.n402 B.n401 585
R48 B.n403 B.n142 585
R49 B.n405 B.n404 585
R50 B.n406 B.n141 585
R51 B.n408 B.n407 585
R52 B.n409 B.n140 585
R53 B.n411 B.n410 585
R54 B.n412 B.n139 585
R55 B.n414 B.n413 585
R56 B.n415 B.n138 585
R57 B.n417 B.n416 585
R58 B.n418 B.n137 585
R59 B.n420 B.n419 585
R60 B.n421 B.n136 585
R61 B.n423 B.n422 585
R62 B.n424 B.n135 585
R63 B.n426 B.n425 585
R64 B.n427 B.n134 585
R65 B.n429 B.n428 585
R66 B.n430 B.n133 585
R67 B.n432 B.n431 585
R68 B.n433 B.n132 585
R69 B.n435 B.n434 585
R70 B.n436 B.n131 585
R71 B.n438 B.n437 585
R72 B.n439 B.n130 585
R73 B.n441 B.n440 585
R74 B.n442 B.n129 585
R75 B.n444 B.n443 585
R76 B.n445 B.n128 585
R77 B.n447 B.n446 585
R78 B.n448 B.n127 585
R79 B.n450 B.n449 585
R80 B.n451 B.n126 585
R81 B.n453 B.n452 585
R82 B.n454 B.n125 585
R83 B.n456 B.n455 585
R84 B.n457 B.n124 585
R85 B.n459 B.n458 585
R86 B.n460 B.n123 585
R87 B.n462 B.n461 585
R88 B.n463 B.n122 585
R89 B.n465 B.n464 585
R90 B.n466 B.n121 585
R91 B.n468 B.n467 585
R92 B.n469 B.n120 585
R93 B.n471 B.n470 585
R94 B.n472 B.n119 585
R95 B.n474 B.n473 585
R96 B.n475 B.n118 585
R97 B.n477 B.n476 585
R98 B.n478 B.n117 585
R99 B.n480 B.n479 585
R100 B.n481 B.n116 585
R101 B.n483 B.n482 585
R102 B.n484 B.n115 585
R103 B.n486 B.n485 585
R104 B.n487 B.n114 585
R105 B.n489 B.n488 585
R106 B.n490 B.n113 585
R107 B.n492 B.n491 585
R108 B.n493 B.n112 585
R109 B.n495 B.n494 585
R110 B.n496 B.n111 585
R111 B.n498 B.n497 585
R112 B.n499 B.n110 585
R113 B.n501 B.n500 585
R114 B.n502 B.n109 585
R115 B.n504 B.n503 585
R116 B.n505 B.n108 585
R117 B.n507 B.n506 585
R118 B.n508 B.n107 585
R119 B.n510 B.n509 585
R120 B.n511 B.n106 585
R121 B.n513 B.n512 585
R122 B.n514 B.n105 585
R123 B.n516 B.n515 585
R124 B.n517 B.n104 585
R125 B.n519 B.n518 585
R126 B.n520 B.n103 585
R127 B.n522 B.n521 585
R128 B.n523 B.n102 585
R129 B.n525 B.n524 585
R130 B.n526 B.n101 585
R131 B.n528 B.n527 585
R132 B.n529 B.n100 585
R133 B.n531 B.n530 585
R134 B.n532 B.n99 585
R135 B.n534 B.n533 585
R136 B.n535 B.n98 585
R137 B.n537 B.n536 585
R138 B.n538 B.n97 585
R139 B.n540 B.n539 585
R140 B.n541 B.n96 585
R141 B.n543 B.n542 585
R142 B.n544 B.n95 585
R143 B.n546 B.n545 585
R144 B.n547 B.n94 585
R145 B.n549 B.n548 585
R146 B.n550 B.n93 585
R147 B.n552 B.n551 585
R148 B.n553 B.n92 585
R149 B.n555 B.n554 585
R150 B.n556 B.n91 585
R151 B.n558 B.n557 585
R152 B.n559 B.n90 585
R153 B.n561 B.n560 585
R154 B.n562 B.n89 585
R155 B.n564 B.n563 585
R156 B.n565 B.n88 585
R157 B.n567 B.n566 585
R158 B.n568 B.n87 585
R159 B.n570 B.n569 585
R160 B.n571 B.n86 585
R161 B.n573 B.n572 585
R162 B.n574 B.n85 585
R163 B.n576 B.n575 585
R164 B.n577 B.n84 585
R165 B.n579 B.n578 585
R166 B.n580 B.n83 585
R167 B.n582 B.n581 585
R168 B.n583 B.n82 585
R169 B.n585 B.n584 585
R170 B.n586 B.n81 585
R171 B.n588 B.n587 585
R172 B.n589 B.n80 585
R173 B.n591 B.n590 585
R174 B.n592 B.n79 585
R175 B.n594 B.n593 585
R176 B.n595 B.n78 585
R177 B.n597 B.n596 585
R178 B.n598 B.n77 585
R179 B.n600 B.n599 585
R180 B.n601 B.n76 585
R181 B.n603 B.n602 585
R182 B.n604 B.n75 585
R183 B.n606 B.n605 585
R184 B.n607 B.n74 585
R185 B.n609 B.n608 585
R186 B.n610 B.n73 585
R187 B.n612 B.n611 585
R188 B.n613 B.n72 585
R189 B.n615 B.n614 585
R190 B.n616 B.n71 585
R191 B.n618 B.n617 585
R192 B.n619 B.n70 585
R193 B.n621 B.n620 585
R194 B.n622 B.n69 585
R195 B.n624 B.n623 585
R196 B.n625 B.n68 585
R197 B.n627 B.n626 585
R198 B.n628 B.n67 585
R199 B.n630 B.n629 585
R200 B.n631 B.n66 585
R201 B.n691 B.n42 585
R202 B.n690 B.n689 585
R203 B.n688 B.n43 585
R204 B.n687 B.n686 585
R205 B.n685 B.n44 585
R206 B.n684 B.n683 585
R207 B.n682 B.n45 585
R208 B.n681 B.n680 585
R209 B.n679 B.n46 585
R210 B.n678 B.n677 585
R211 B.n676 B.n47 585
R212 B.n675 B.n674 585
R213 B.n673 B.n48 585
R214 B.n672 B.n671 585
R215 B.n670 B.n49 585
R216 B.n668 B.n667 585
R217 B.n666 B.n52 585
R218 B.n665 B.n664 585
R219 B.n663 B.n53 585
R220 B.n662 B.n661 585
R221 B.n660 B.n54 585
R222 B.n659 B.n658 585
R223 B.n657 B.n55 585
R224 B.n656 B.n655 585
R225 B.n654 B.n653 585
R226 B.n652 B.n59 585
R227 B.n651 B.n650 585
R228 B.n649 B.n60 585
R229 B.n648 B.n647 585
R230 B.n646 B.n61 585
R231 B.n645 B.n644 585
R232 B.n643 B.n62 585
R233 B.n642 B.n641 585
R234 B.n640 B.n63 585
R235 B.n639 B.n638 585
R236 B.n637 B.n64 585
R237 B.n636 B.n635 585
R238 B.n634 B.n65 585
R239 B.n633 B.n632 585
R240 B.n693 B.n692 585
R241 B.n694 B.n41 585
R242 B.n696 B.n695 585
R243 B.n697 B.n40 585
R244 B.n699 B.n698 585
R245 B.n700 B.n39 585
R246 B.n702 B.n701 585
R247 B.n703 B.n38 585
R248 B.n705 B.n704 585
R249 B.n706 B.n37 585
R250 B.n708 B.n707 585
R251 B.n709 B.n36 585
R252 B.n711 B.n710 585
R253 B.n712 B.n35 585
R254 B.n714 B.n713 585
R255 B.n715 B.n34 585
R256 B.n717 B.n716 585
R257 B.n718 B.n33 585
R258 B.n720 B.n719 585
R259 B.n721 B.n32 585
R260 B.n723 B.n722 585
R261 B.n724 B.n31 585
R262 B.n726 B.n725 585
R263 B.n727 B.n30 585
R264 B.n729 B.n728 585
R265 B.n730 B.n29 585
R266 B.n732 B.n731 585
R267 B.n733 B.n28 585
R268 B.n735 B.n734 585
R269 B.n736 B.n27 585
R270 B.n738 B.n737 585
R271 B.n739 B.n26 585
R272 B.n741 B.n740 585
R273 B.n742 B.n25 585
R274 B.n744 B.n743 585
R275 B.n745 B.n24 585
R276 B.n747 B.n746 585
R277 B.n748 B.n23 585
R278 B.n750 B.n749 585
R279 B.n751 B.n22 585
R280 B.n753 B.n752 585
R281 B.n754 B.n21 585
R282 B.n756 B.n755 585
R283 B.n757 B.n20 585
R284 B.n759 B.n758 585
R285 B.n760 B.n19 585
R286 B.n762 B.n761 585
R287 B.n763 B.n18 585
R288 B.n765 B.n764 585
R289 B.n766 B.n17 585
R290 B.n768 B.n767 585
R291 B.n769 B.n16 585
R292 B.n771 B.n770 585
R293 B.n772 B.n15 585
R294 B.n774 B.n773 585
R295 B.n775 B.n14 585
R296 B.n777 B.n776 585
R297 B.n778 B.n13 585
R298 B.n780 B.n779 585
R299 B.n781 B.n12 585
R300 B.n783 B.n782 585
R301 B.n784 B.n11 585
R302 B.n786 B.n785 585
R303 B.n787 B.n10 585
R304 B.n789 B.n788 585
R305 B.n790 B.n9 585
R306 B.n792 B.n791 585
R307 B.n793 B.n8 585
R308 B.n795 B.n794 585
R309 B.n796 B.n7 585
R310 B.n798 B.n797 585
R311 B.n799 B.n6 585
R312 B.n801 B.n800 585
R313 B.n802 B.n5 585
R314 B.n804 B.n803 585
R315 B.n805 B.n4 585
R316 B.n807 B.n806 585
R317 B.n808 B.n3 585
R318 B.n810 B.n809 585
R319 B.n811 B.n0 585
R320 B.n2 B.n1 585
R321 B.n209 B.n208 585
R322 B.n210 B.n207 585
R323 B.n212 B.n211 585
R324 B.n213 B.n206 585
R325 B.n215 B.n214 585
R326 B.n216 B.n205 585
R327 B.n218 B.n217 585
R328 B.n219 B.n204 585
R329 B.n221 B.n220 585
R330 B.n222 B.n203 585
R331 B.n224 B.n223 585
R332 B.n225 B.n202 585
R333 B.n227 B.n226 585
R334 B.n228 B.n201 585
R335 B.n230 B.n229 585
R336 B.n231 B.n200 585
R337 B.n233 B.n232 585
R338 B.n234 B.n199 585
R339 B.n236 B.n235 585
R340 B.n237 B.n198 585
R341 B.n239 B.n238 585
R342 B.n240 B.n197 585
R343 B.n242 B.n241 585
R344 B.n243 B.n196 585
R345 B.n245 B.n244 585
R346 B.n246 B.n195 585
R347 B.n248 B.n247 585
R348 B.n249 B.n194 585
R349 B.n251 B.n250 585
R350 B.n252 B.n193 585
R351 B.n254 B.n253 585
R352 B.n255 B.n192 585
R353 B.n257 B.n256 585
R354 B.n258 B.n191 585
R355 B.n260 B.n259 585
R356 B.n261 B.n190 585
R357 B.n263 B.n262 585
R358 B.n264 B.n189 585
R359 B.n266 B.n265 585
R360 B.n267 B.n188 585
R361 B.n269 B.n268 585
R362 B.n270 B.n187 585
R363 B.n272 B.n271 585
R364 B.n273 B.n186 585
R365 B.n275 B.n274 585
R366 B.n276 B.n185 585
R367 B.n278 B.n277 585
R368 B.n279 B.n184 585
R369 B.n281 B.n280 585
R370 B.n282 B.n183 585
R371 B.n284 B.n283 585
R372 B.n285 B.n182 585
R373 B.n287 B.n286 585
R374 B.n288 B.n181 585
R375 B.n290 B.n289 585
R376 B.n291 B.n180 585
R377 B.n293 B.n292 585
R378 B.n294 B.n179 585
R379 B.n296 B.n295 585
R380 B.n297 B.n178 585
R381 B.n299 B.n298 585
R382 B.n300 B.n177 585
R383 B.n302 B.n301 585
R384 B.n303 B.n176 585
R385 B.n305 B.n304 585
R386 B.n306 B.n175 585
R387 B.n308 B.n307 585
R388 B.n309 B.n174 585
R389 B.n311 B.n310 585
R390 B.n312 B.n173 585
R391 B.n314 B.n313 585
R392 B.n315 B.n172 585
R393 B.n317 B.n316 585
R394 B.n318 B.n171 585
R395 B.n320 B.n319 585
R396 B.n321 B.n170 585
R397 B.n323 B.n322 585
R398 B.n324 B.n169 585
R399 B.n326 B.n325 585
R400 B.n327 B.n326 463.671
R401 B.n390 B.n147 463.671
R402 B.n632 B.n631 463.671
R403 B.n692 B.n691 463.671
R404 B.n813 B.n812 256.663
R405 B.n812 B.n811 235.042
R406 B.n812 B.n2 235.042
R407 B.n160 B.t6 227.155
R408 B.n362 B.t0 227.155
R409 B.n56 B.t3 227.155
R410 B.n50 B.t9 227.155
R411 B.n362 B.t1 221.481
R412 B.n56 B.t5 221.481
R413 B.n160 B.t7 221.48
R414 B.n50 B.t11 221.48
R415 B.n328 B.n327 163.367
R416 B.n328 B.n167 163.367
R417 B.n332 B.n167 163.367
R418 B.n333 B.n332 163.367
R419 B.n334 B.n333 163.367
R420 B.n334 B.n165 163.367
R421 B.n338 B.n165 163.367
R422 B.n339 B.n338 163.367
R423 B.n340 B.n339 163.367
R424 B.n340 B.n163 163.367
R425 B.n344 B.n163 163.367
R426 B.n345 B.n344 163.367
R427 B.n346 B.n345 163.367
R428 B.n346 B.n159 163.367
R429 B.n351 B.n159 163.367
R430 B.n352 B.n351 163.367
R431 B.n353 B.n352 163.367
R432 B.n353 B.n157 163.367
R433 B.n357 B.n157 163.367
R434 B.n358 B.n357 163.367
R435 B.n359 B.n358 163.367
R436 B.n359 B.n155 163.367
R437 B.n366 B.n155 163.367
R438 B.n367 B.n366 163.367
R439 B.n368 B.n367 163.367
R440 B.n368 B.n153 163.367
R441 B.n372 B.n153 163.367
R442 B.n373 B.n372 163.367
R443 B.n374 B.n373 163.367
R444 B.n374 B.n151 163.367
R445 B.n378 B.n151 163.367
R446 B.n379 B.n378 163.367
R447 B.n380 B.n379 163.367
R448 B.n380 B.n149 163.367
R449 B.n384 B.n149 163.367
R450 B.n385 B.n384 163.367
R451 B.n386 B.n385 163.367
R452 B.n386 B.n147 163.367
R453 B.n631 B.n630 163.367
R454 B.n630 B.n67 163.367
R455 B.n626 B.n67 163.367
R456 B.n626 B.n625 163.367
R457 B.n625 B.n624 163.367
R458 B.n624 B.n69 163.367
R459 B.n620 B.n69 163.367
R460 B.n620 B.n619 163.367
R461 B.n619 B.n618 163.367
R462 B.n618 B.n71 163.367
R463 B.n614 B.n71 163.367
R464 B.n614 B.n613 163.367
R465 B.n613 B.n612 163.367
R466 B.n612 B.n73 163.367
R467 B.n608 B.n73 163.367
R468 B.n608 B.n607 163.367
R469 B.n607 B.n606 163.367
R470 B.n606 B.n75 163.367
R471 B.n602 B.n75 163.367
R472 B.n602 B.n601 163.367
R473 B.n601 B.n600 163.367
R474 B.n600 B.n77 163.367
R475 B.n596 B.n77 163.367
R476 B.n596 B.n595 163.367
R477 B.n595 B.n594 163.367
R478 B.n594 B.n79 163.367
R479 B.n590 B.n79 163.367
R480 B.n590 B.n589 163.367
R481 B.n589 B.n588 163.367
R482 B.n588 B.n81 163.367
R483 B.n584 B.n81 163.367
R484 B.n584 B.n583 163.367
R485 B.n583 B.n582 163.367
R486 B.n582 B.n83 163.367
R487 B.n578 B.n83 163.367
R488 B.n578 B.n577 163.367
R489 B.n577 B.n576 163.367
R490 B.n576 B.n85 163.367
R491 B.n572 B.n85 163.367
R492 B.n572 B.n571 163.367
R493 B.n571 B.n570 163.367
R494 B.n570 B.n87 163.367
R495 B.n566 B.n87 163.367
R496 B.n566 B.n565 163.367
R497 B.n565 B.n564 163.367
R498 B.n564 B.n89 163.367
R499 B.n560 B.n89 163.367
R500 B.n560 B.n559 163.367
R501 B.n559 B.n558 163.367
R502 B.n558 B.n91 163.367
R503 B.n554 B.n91 163.367
R504 B.n554 B.n553 163.367
R505 B.n553 B.n552 163.367
R506 B.n552 B.n93 163.367
R507 B.n548 B.n93 163.367
R508 B.n548 B.n547 163.367
R509 B.n547 B.n546 163.367
R510 B.n546 B.n95 163.367
R511 B.n542 B.n95 163.367
R512 B.n542 B.n541 163.367
R513 B.n541 B.n540 163.367
R514 B.n540 B.n97 163.367
R515 B.n536 B.n97 163.367
R516 B.n536 B.n535 163.367
R517 B.n535 B.n534 163.367
R518 B.n534 B.n99 163.367
R519 B.n530 B.n99 163.367
R520 B.n530 B.n529 163.367
R521 B.n529 B.n528 163.367
R522 B.n528 B.n101 163.367
R523 B.n524 B.n101 163.367
R524 B.n524 B.n523 163.367
R525 B.n523 B.n522 163.367
R526 B.n522 B.n103 163.367
R527 B.n518 B.n103 163.367
R528 B.n518 B.n517 163.367
R529 B.n517 B.n516 163.367
R530 B.n516 B.n105 163.367
R531 B.n512 B.n105 163.367
R532 B.n512 B.n511 163.367
R533 B.n511 B.n510 163.367
R534 B.n510 B.n107 163.367
R535 B.n506 B.n107 163.367
R536 B.n506 B.n505 163.367
R537 B.n505 B.n504 163.367
R538 B.n504 B.n109 163.367
R539 B.n500 B.n109 163.367
R540 B.n500 B.n499 163.367
R541 B.n499 B.n498 163.367
R542 B.n498 B.n111 163.367
R543 B.n494 B.n111 163.367
R544 B.n494 B.n493 163.367
R545 B.n493 B.n492 163.367
R546 B.n492 B.n113 163.367
R547 B.n488 B.n113 163.367
R548 B.n488 B.n487 163.367
R549 B.n487 B.n486 163.367
R550 B.n486 B.n115 163.367
R551 B.n482 B.n115 163.367
R552 B.n482 B.n481 163.367
R553 B.n481 B.n480 163.367
R554 B.n480 B.n117 163.367
R555 B.n476 B.n117 163.367
R556 B.n476 B.n475 163.367
R557 B.n475 B.n474 163.367
R558 B.n474 B.n119 163.367
R559 B.n470 B.n119 163.367
R560 B.n470 B.n469 163.367
R561 B.n469 B.n468 163.367
R562 B.n468 B.n121 163.367
R563 B.n464 B.n121 163.367
R564 B.n464 B.n463 163.367
R565 B.n463 B.n462 163.367
R566 B.n462 B.n123 163.367
R567 B.n458 B.n123 163.367
R568 B.n458 B.n457 163.367
R569 B.n457 B.n456 163.367
R570 B.n456 B.n125 163.367
R571 B.n452 B.n125 163.367
R572 B.n452 B.n451 163.367
R573 B.n451 B.n450 163.367
R574 B.n450 B.n127 163.367
R575 B.n446 B.n127 163.367
R576 B.n446 B.n445 163.367
R577 B.n445 B.n444 163.367
R578 B.n444 B.n129 163.367
R579 B.n440 B.n129 163.367
R580 B.n440 B.n439 163.367
R581 B.n439 B.n438 163.367
R582 B.n438 B.n131 163.367
R583 B.n434 B.n131 163.367
R584 B.n434 B.n433 163.367
R585 B.n433 B.n432 163.367
R586 B.n432 B.n133 163.367
R587 B.n428 B.n133 163.367
R588 B.n428 B.n427 163.367
R589 B.n427 B.n426 163.367
R590 B.n426 B.n135 163.367
R591 B.n422 B.n135 163.367
R592 B.n422 B.n421 163.367
R593 B.n421 B.n420 163.367
R594 B.n420 B.n137 163.367
R595 B.n416 B.n137 163.367
R596 B.n416 B.n415 163.367
R597 B.n415 B.n414 163.367
R598 B.n414 B.n139 163.367
R599 B.n410 B.n139 163.367
R600 B.n410 B.n409 163.367
R601 B.n409 B.n408 163.367
R602 B.n408 B.n141 163.367
R603 B.n404 B.n141 163.367
R604 B.n404 B.n403 163.367
R605 B.n403 B.n402 163.367
R606 B.n402 B.n143 163.367
R607 B.n398 B.n143 163.367
R608 B.n398 B.n397 163.367
R609 B.n397 B.n396 163.367
R610 B.n396 B.n145 163.367
R611 B.n392 B.n145 163.367
R612 B.n392 B.n391 163.367
R613 B.n391 B.n390 163.367
R614 B.n691 B.n690 163.367
R615 B.n690 B.n43 163.367
R616 B.n686 B.n43 163.367
R617 B.n686 B.n685 163.367
R618 B.n685 B.n684 163.367
R619 B.n684 B.n45 163.367
R620 B.n680 B.n45 163.367
R621 B.n680 B.n679 163.367
R622 B.n679 B.n678 163.367
R623 B.n678 B.n47 163.367
R624 B.n674 B.n47 163.367
R625 B.n674 B.n673 163.367
R626 B.n673 B.n672 163.367
R627 B.n672 B.n49 163.367
R628 B.n667 B.n49 163.367
R629 B.n667 B.n666 163.367
R630 B.n666 B.n665 163.367
R631 B.n665 B.n53 163.367
R632 B.n661 B.n53 163.367
R633 B.n661 B.n660 163.367
R634 B.n660 B.n659 163.367
R635 B.n659 B.n55 163.367
R636 B.n655 B.n55 163.367
R637 B.n655 B.n654 163.367
R638 B.n654 B.n59 163.367
R639 B.n650 B.n59 163.367
R640 B.n650 B.n649 163.367
R641 B.n649 B.n648 163.367
R642 B.n648 B.n61 163.367
R643 B.n644 B.n61 163.367
R644 B.n644 B.n643 163.367
R645 B.n643 B.n642 163.367
R646 B.n642 B.n63 163.367
R647 B.n638 B.n63 163.367
R648 B.n638 B.n637 163.367
R649 B.n637 B.n636 163.367
R650 B.n636 B.n65 163.367
R651 B.n632 B.n65 163.367
R652 B.n692 B.n41 163.367
R653 B.n696 B.n41 163.367
R654 B.n697 B.n696 163.367
R655 B.n698 B.n697 163.367
R656 B.n698 B.n39 163.367
R657 B.n702 B.n39 163.367
R658 B.n703 B.n702 163.367
R659 B.n704 B.n703 163.367
R660 B.n704 B.n37 163.367
R661 B.n708 B.n37 163.367
R662 B.n709 B.n708 163.367
R663 B.n710 B.n709 163.367
R664 B.n710 B.n35 163.367
R665 B.n714 B.n35 163.367
R666 B.n715 B.n714 163.367
R667 B.n716 B.n715 163.367
R668 B.n716 B.n33 163.367
R669 B.n720 B.n33 163.367
R670 B.n721 B.n720 163.367
R671 B.n722 B.n721 163.367
R672 B.n722 B.n31 163.367
R673 B.n726 B.n31 163.367
R674 B.n727 B.n726 163.367
R675 B.n728 B.n727 163.367
R676 B.n728 B.n29 163.367
R677 B.n732 B.n29 163.367
R678 B.n733 B.n732 163.367
R679 B.n734 B.n733 163.367
R680 B.n734 B.n27 163.367
R681 B.n738 B.n27 163.367
R682 B.n739 B.n738 163.367
R683 B.n740 B.n739 163.367
R684 B.n740 B.n25 163.367
R685 B.n744 B.n25 163.367
R686 B.n745 B.n744 163.367
R687 B.n746 B.n745 163.367
R688 B.n746 B.n23 163.367
R689 B.n750 B.n23 163.367
R690 B.n751 B.n750 163.367
R691 B.n752 B.n751 163.367
R692 B.n752 B.n21 163.367
R693 B.n756 B.n21 163.367
R694 B.n757 B.n756 163.367
R695 B.n758 B.n757 163.367
R696 B.n758 B.n19 163.367
R697 B.n762 B.n19 163.367
R698 B.n763 B.n762 163.367
R699 B.n764 B.n763 163.367
R700 B.n764 B.n17 163.367
R701 B.n768 B.n17 163.367
R702 B.n769 B.n768 163.367
R703 B.n770 B.n769 163.367
R704 B.n770 B.n15 163.367
R705 B.n774 B.n15 163.367
R706 B.n775 B.n774 163.367
R707 B.n776 B.n775 163.367
R708 B.n776 B.n13 163.367
R709 B.n780 B.n13 163.367
R710 B.n781 B.n780 163.367
R711 B.n782 B.n781 163.367
R712 B.n782 B.n11 163.367
R713 B.n786 B.n11 163.367
R714 B.n787 B.n786 163.367
R715 B.n788 B.n787 163.367
R716 B.n788 B.n9 163.367
R717 B.n792 B.n9 163.367
R718 B.n793 B.n792 163.367
R719 B.n794 B.n793 163.367
R720 B.n794 B.n7 163.367
R721 B.n798 B.n7 163.367
R722 B.n799 B.n798 163.367
R723 B.n800 B.n799 163.367
R724 B.n800 B.n5 163.367
R725 B.n804 B.n5 163.367
R726 B.n805 B.n804 163.367
R727 B.n806 B.n805 163.367
R728 B.n806 B.n3 163.367
R729 B.n810 B.n3 163.367
R730 B.n811 B.n810 163.367
R731 B.n208 B.n2 163.367
R732 B.n208 B.n207 163.367
R733 B.n212 B.n207 163.367
R734 B.n213 B.n212 163.367
R735 B.n214 B.n213 163.367
R736 B.n214 B.n205 163.367
R737 B.n218 B.n205 163.367
R738 B.n219 B.n218 163.367
R739 B.n220 B.n219 163.367
R740 B.n220 B.n203 163.367
R741 B.n224 B.n203 163.367
R742 B.n225 B.n224 163.367
R743 B.n226 B.n225 163.367
R744 B.n226 B.n201 163.367
R745 B.n230 B.n201 163.367
R746 B.n231 B.n230 163.367
R747 B.n232 B.n231 163.367
R748 B.n232 B.n199 163.367
R749 B.n236 B.n199 163.367
R750 B.n237 B.n236 163.367
R751 B.n238 B.n237 163.367
R752 B.n238 B.n197 163.367
R753 B.n242 B.n197 163.367
R754 B.n243 B.n242 163.367
R755 B.n244 B.n243 163.367
R756 B.n244 B.n195 163.367
R757 B.n248 B.n195 163.367
R758 B.n249 B.n248 163.367
R759 B.n250 B.n249 163.367
R760 B.n250 B.n193 163.367
R761 B.n254 B.n193 163.367
R762 B.n255 B.n254 163.367
R763 B.n256 B.n255 163.367
R764 B.n256 B.n191 163.367
R765 B.n260 B.n191 163.367
R766 B.n261 B.n260 163.367
R767 B.n262 B.n261 163.367
R768 B.n262 B.n189 163.367
R769 B.n266 B.n189 163.367
R770 B.n267 B.n266 163.367
R771 B.n268 B.n267 163.367
R772 B.n268 B.n187 163.367
R773 B.n272 B.n187 163.367
R774 B.n273 B.n272 163.367
R775 B.n274 B.n273 163.367
R776 B.n274 B.n185 163.367
R777 B.n278 B.n185 163.367
R778 B.n279 B.n278 163.367
R779 B.n280 B.n279 163.367
R780 B.n280 B.n183 163.367
R781 B.n284 B.n183 163.367
R782 B.n285 B.n284 163.367
R783 B.n286 B.n285 163.367
R784 B.n286 B.n181 163.367
R785 B.n290 B.n181 163.367
R786 B.n291 B.n290 163.367
R787 B.n292 B.n291 163.367
R788 B.n292 B.n179 163.367
R789 B.n296 B.n179 163.367
R790 B.n297 B.n296 163.367
R791 B.n298 B.n297 163.367
R792 B.n298 B.n177 163.367
R793 B.n302 B.n177 163.367
R794 B.n303 B.n302 163.367
R795 B.n304 B.n303 163.367
R796 B.n304 B.n175 163.367
R797 B.n308 B.n175 163.367
R798 B.n309 B.n308 163.367
R799 B.n310 B.n309 163.367
R800 B.n310 B.n173 163.367
R801 B.n314 B.n173 163.367
R802 B.n315 B.n314 163.367
R803 B.n316 B.n315 163.367
R804 B.n316 B.n171 163.367
R805 B.n320 B.n171 163.367
R806 B.n321 B.n320 163.367
R807 B.n322 B.n321 163.367
R808 B.n322 B.n169 163.367
R809 B.n326 B.n169 163.367
R810 B.n363 B.t2 141.965
R811 B.n57 B.t4 141.965
R812 B.n161 B.t8 141.964
R813 B.n51 B.t10 141.964
R814 B.n161 B.n160 79.5157
R815 B.n363 B.n362 79.5157
R816 B.n57 B.n56 79.5157
R817 B.n51 B.n50 79.5157
R818 B.n349 B.n161 59.5399
R819 B.n364 B.n363 59.5399
R820 B.n58 B.n57 59.5399
R821 B.n669 B.n51 59.5399
R822 B.n693 B.n42 30.1273
R823 B.n633 B.n66 30.1273
R824 B.n389 B.n388 30.1273
R825 B.n325 B.n168 30.1273
R826 B B.n813 18.0485
R827 B.n694 B.n693 10.6151
R828 B.n695 B.n694 10.6151
R829 B.n695 B.n40 10.6151
R830 B.n699 B.n40 10.6151
R831 B.n700 B.n699 10.6151
R832 B.n701 B.n700 10.6151
R833 B.n701 B.n38 10.6151
R834 B.n705 B.n38 10.6151
R835 B.n706 B.n705 10.6151
R836 B.n707 B.n706 10.6151
R837 B.n707 B.n36 10.6151
R838 B.n711 B.n36 10.6151
R839 B.n712 B.n711 10.6151
R840 B.n713 B.n712 10.6151
R841 B.n713 B.n34 10.6151
R842 B.n717 B.n34 10.6151
R843 B.n718 B.n717 10.6151
R844 B.n719 B.n718 10.6151
R845 B.n719 B.n32 10.6151
R846 B.n723 B.n32 10.6151
R847 B.n724 B.n723 10.6151
R848 B.n725 B.n724 10.6151
R849 B.n725 B.n30 10.6151
R850 B.n729 B.n30 10.6151
R851 B.n730 B.n729 10.6151
R852 B.n731 B.n730 10.6151
R853 B.n731 B.n28 10.6151
R854 B.n735 B.n28 10.6151
R855 B.n736 B.n735 10.6151
R856 B.n737 B.n736 10.6151
R857 B.n737 B.n26 10.6151
R858 B.n741 B.n26 10.6151
R859 B.n742 B.n741 10.6151
R860 B.n743 B.n742 10.6151
R861 B.n743 B.n24 10.6151
R862 B.n747 B.n24 10.6151
R863 B.n748 B.n747 10.6151
R864 B.n749 B.n748 10.6151
R865 B.n749 B.n22 10.6151
R866 B.n753 B.n22 10.6151
R867 B.n754 B.n753 10.6151
R868 B.n755 B.n754 10.6151
R869 B.n755 B.n20 10.6151
R870 B.n759 B.n20 10.6151
R871 B.n760 B.n759 10.6151
R872 B.n761 B.n760 10.6151
R873 B.n761 B.n18 10.6151
R874 B.n765 B.n18 10.6151
R875 B.n766 B.n765 10.6151
R876 B.n767 B.n766 10.6151
R877 B.n767 B.n16 10.6151
R878 B.n771 B.n16 10.6151
R879 B.n772 B.n771 10.6151
R880 B.n773 B.n772 10.6151
R881 B.n773 B.n14 10.6151
R882 B.n777 B.n14 10.6151
R883 B.n778 B.n777 10.6151
R884 B.n779 B.n778 10.6151
R885 B.n779 B.n12 10.6151
R886 B.n783 B.n12 10.6151
R887 B.n784 B.n783 10.6151
R888 B.n785 B.n784 10.6151
R889 B.n785 B.n10 10.6151
R890 B.n789 B.n10 10.6151
R891 B.n790 B.n789 10.6151
R892 B.n791 B.n790 10.6151
R893 B.n791 B.n8 10.6151
R894 B.n795 B.n8 10.6151
R895 B.n796 B.n795 10.6151
R896 B.n797 B.n796 10.6151
R897 B.n797 B.n6 10.6151
R898 B.n801 B.n6 10.6151
R899 B.n802 B.n801 10.6151
R900 B.n803 B.n802 10.6151
R901 B.n803 B.n4 10.6151
R902 B.n807 B.n4 10.6151
R903 B.n808 B.n807 10.6151
R904 B.n809 B.n808 10.6151
R905 B.n809 B.n0 10.6151
R906 B.n689 B.n42 10.6151
R907 B.n689 B.n688 10.6151
R908 B.n688 B.n687 10.6151
R909 B.n687 B.n44 10.6151
R910 B.n683 B.n44 10.6151
R911 B.n683 B.n682 10.6151
R912 B.n682 B.n681 10.6151
R913 B.n681 B.n46 10.6151
R914 B.n677 B.n46 10.6151
R915 B.n677 B.n676 10.6151
R916 B.n676 B.n675 10.6151
R917 B.n675 B.n48 10.6151
R918 B.n671 B.n48 10.6151
R919 B.n671 B.n670 10.6151
R920 B.n668 B.n52 10.6151
R921 B.n664 B.n52 10.6151
R922 B.n664 B.n663 10.6151
R923 B.n663 B.n662 10.6151
R924 B.n662 B.n54 10.6151
R925 B.n658 B.n54 10.6151
R926 B.n658 B.n657 10.6151
R927 B.n657 B.n656 10.6151
R928 B.n653 B.n652 10.6151
R929 B.n652 B.n651 10.6151
R930 B.n651 B.n60 10.6151
R931 B.n647 B.n60 10.6151
R932 B.n647 B.n646 10.6151
R933 B.n646 B.n645 10.6151
R934 B.n645 B.n62 10.6151
R935 B.n641 B.n62 10.6151
R936 B.n641 B.n640 10.6151
R937 B.n640 B.n639 10.6151
R938 B.n639 B.n64 10.6151
R939 B.n635 B.n64 10.6151
R940 B.n635 B.n634 10.6151
R941 B.n634 B.n633 10.6151
R942 B.n629 B.n66 10.6151
R943 B.n629 B.n628 10.6151
R944 B.n628 B.n627 10.6151
R945 B.n627 B.n68 10.6151
R946 B.n623 B.n68 10.6151
R947 B.n623 B.n622 10.6151
R948 B.n622 B.n621 10.6151
R949 B.n621 B.n70 10.6151
R950 B.n617 B.n70 10.6151
R951 B.n617 B.n616 10.6151
R952 B.n616 B.n615 10.6151
R953 B.n615 B.n72 10.6151
R954 B.n611 B.n72 10.6151
R955 B.n611 B.n610 10.6151
R956 B.n610 B.n609 10.6151
R957 B.n609 B.n74 10.6151
R958 B.n605 B.n74 10.6151
R959 B.n605 B.n604 10.6151
R960 B.n604 B.n603 10.6151
R961 B.n603 B.n76 10.6151
R962 B.n599 B.n76 10.6151
R963 B.n599 B.n598 10.6151
R964 B.n598 B.n597 10.6151
R965 B.n597 B.n78 10.6151
R966 B.n593 B.n78 10.6151
R967 B.n593 B.n592 10.6151
R968 B.n592 B.n591 10.6151
R969 B.n591 B.n80 10.6151
R970 B.n587 B.n80 10.6151
R971 B.n587 B.n586 10.6151
R972 B.n586 B.n585 10.6151
R973 B.n585 B.n82 10.6151
R974 B.n581 B.n82 10.6151
R975 B.n581 B.n580 10.6151
R976 B.n580 B.n579 10.6151
R977 B.n579 B.n84 10.6151
R978 B.n575 B.n84 10.6151
R979 B.n575 B.n574 10.6151
R980 B.n574 B.n573 10.6151
R981 B.n573 B.n86 10.6151
R982 B.n569 B.n86 10.6151
R983 B.n569 B.n568 10.6151
R984 B.n568 B.n567 10.6151
R985 B.n567 B.n88 10.6151
R986 B.n563 B.n88 10.6151
R987 B.n563 B.n562 10.6151
R988 B.n562 B.n561 10.6151
R989 B.n561 B.n90 10.6151
R990 B.n557 B.n90 10.6151
R991 B.n557 B.n556 10.6151
R992 B.n556 B.n555 10.6151
R993 B.n555 B.n92 10.6151
R994 B.n551 B.n92 10.6151
R995 B.n551 B.n550 10.6151
R996 B.n550 B.n549 10.6151
R997 B.n549 B.n94 10.6151
R998 B.n545 B.n94 10.6151
R999 B.n545 B.n544 10.6151
R1000 B.n544 B.n543 10.6151
R1001 B.n543 B.n96 10.6151
R1002 B.n539 B.n96 10.6151
R1003 B.n539 B.n538 10.6151
R1004 B.n538 B.n537 10.6151
R1005 B.n537 B.n98 10.6151
R1006 B.n533 B.n98 10.6151
R1007 B.n533 B.n532 10.6151
R1008 B.n532 B.n531 10.6151
R1009 B.n531 B.n100 10.6151
R1010 B.n527 B.n100 10.6151
R1011 B.n527 B.n526 10.6151
R1012 B.n526 B.n525 10.6151
R1013 B.n525 B.n102 10.6151
R1014 B.n521 B.n102 10.6151
R1015 B.n521 B.n520 10.6151
R1016 B.n520 B.n519 10.6151
R1017 B.n519 B.n104 10.6151
R1018 B.n515 B.n104 10.6151
R1019 B.n515 B.n514 10.6151
R1020 B.n514 B.n513 10.6151
R1021 B.n513 B.n106 10.6151
R1022 B.n509 B.n106 10.6151
R1023 B.n509 B.n508 10.6151
R1024 B.n508 B.n507 10.6151
R1025 B.n507 B.n108 10.6151
R1026 B.n503 B.n108 10.6151
R1027 B.n503 B.n502 10.6151
R1028 B.n502 B.n501 10.6151
R1029 B.n501 B.n110 10.6151
R1030 B.n497 B.n110 10.6151
R1031 B.n497 B.n496 10.6151
R1032 B.n496 B.n495 10.6151
R1033 B.n495 B.n112 10.6151
R1034 B.n491 B.n112 10.6151
R1035 B.n491 B.n490 10.6151
R1036 B.n490 B.n489 10.6151
R1037 B.n489 B.n114 10.6151
R1038 B.n485 B.n114 10.6151
R1039 B.n485 B.n484 10.6151
R1040 B.n484 B.n483 10.6151
R1041 B.n483 B.n116 10.6151
R1042 B.n479 B.n116 10.6151
R1043 B.n479 B.n478 10.6151
R1044 B.n478 B.n477 10.6151
R1045 B.n477 B.n118 10.6151
R1046 B.n473 B.n118 10.6151
R1047 B.n473 B.n472 10.6151
R1048 B.n472 B.n471 10.6151
R1049 B.n471 B.n120 10.6151
R1050 B.n467 B.n120 10.6151
R1051 B.n467 B.n466 10.6151
R1052 B.n466 B.n465 10.6151
R1053 B.n465 B.n122 10.6151
R1054 B.n461 B.n122 10.6151
R1055 B.n461 B.n460 10.6151
R1056 B.n460 B.n459 10.6151
R1057 B.n459 B.n124 10.6151
R1058 B.n455 B.n124 10.6151
R1059 B.n455 B.n454 10.6151
R1060 B.n454 B.n453 10.6151
R1061 B.n453 B.n126 10.6151
R1062 B.n449 B.n126 10.6151
R1063 B.n449 B.n448 10.6151
R1064 B.n448 B.n447 10.6151
R1065 B.n447 B.n128 10.6151
R1066 B.n443 B.n128 10.6151
R1067 B.n443 B.n442 10.6151
R1068 B.n442 B.n441 10.6151
R1069 B.n441 B.n130 10.6151
R1070 B.n437 B.n130 10.6151
R1071 B.n437 B.n436 10.6151
R1072 B.n436 B.n435 10.6151
R1073 B.n435 B.n132 10.6151
R1074 B.n431 B.n132 10.6151
R1075 B.n431 B.n430 10.6151
R1076 B.n430 B.n429 10.6151
R1077 B.n429 B.n134 10.6151
R1078 B.n425 B.n134 10.6151
R1079 B.n425 B.n424 10.6151
R1080 B.n424 B.n423 10.6151
R1081 B.n423 B.n136 10.6151
R1082 B.n419 B.n136 10.6151
R1083 B.n419 B.n418 10.6151
R1084 B.n418 B.n417 10.6151
R1085 B.n417 B.n138 10.6151
R1086 B.n413 B.n138 10.6151
R1087 B.n413 B.n412 10.6151
R1088 B.n412 B.n411 10.6151
R1089 B.n411 B.n140 10.6151
R1090 B.n407 B.n140 10.6151
R1091 B.n407 B.n406 10.6151
R1092 B.n406 B.n405 10.6151
R1093 B.n405 B.n142 10.6151
R1094 B.n401 B.n142 10.6151
R1095 B.n401 B.n400 10.6151
R1096 B.n400 B.n399 10.6151
R1097 B.n399 B.n144 10.6151
R1098 B.n395 B.n144 10.6151
R1099 B.n395 B.n394 10.6151
R1100 B.n394 B.n393 10.6151
R1101 B.n393 B.n146 10.6151
R1102 B.n389 B.n146 10.6151
R1103 B.n209 B.n1 10.6151
R1104 B.n210 B.n209 10.6151
R1105 B.n211 B.n210 10.6151
R1106 B.n211 B.n206 10.6151
R1107 B.n215 B.n206 10.6151
R1108 B.n216 B.n215 10.6151
R1109 B.n217 B.n216 10.6151
R1110 B.n217 B.n204 10.6151
R1111 B.n221 B.n204 10.6151
R1112 B.n222 B.n221 10.6151
R1113 B.n223 B.n222 10.6151
R1114 B.n223 B.n202 10.6151
R1115 B.n227 B.n202 10.6151
R1116 B.n228 B.n227 10.6151
R1117 B.n229 B.n228 10.6151
R1118 B.n229 B.n200 10.6151
R1119 B.n233 B.n200 10.6151
R1120 B.n234 B.n233 10.6151
R1121 B.n235 B.n234 10.6151
R1122 B.n235 B.n198 10.6151
R1123 B.n239 B.n198 10.6151
R1124 B.n240 B.n239 10.6151
R1125 B.n241 B.n240 10.6151
R1126 B.n241 B.n196 10.6151
R1127 B.n245 B.n196 10.6151
R1128 B.n246 B.n245 10.6151
R1129 B.n247 B.n246 10.6151
R1130 B.n247 B.n194 10.6151
R1131 B.n251 B.n194 10.6151
R1132 B.n252 B.n251 10.6151
R1133 B.n253 B.n252 10.6151
R1134 B.n253 B.n192 10.6151
R1135 B.n257 B.n192 10.6151
R1136 B.n258 B.n257 10.6151
R1137 B.n259 B.n258 10.6151
R1138 B.n259 B.n190 10.6151
R1139 B.n263 B.n190 10.6151
R1140 B.n264 B.n263 10.6151
R1141 B.n265 B.n264 10.6151
R1142 B.n265 B.n188 10.6151
R1143 B.n269 B.n188 10.6151
R1144 B.n270 B.n269 10.6151
R1145 B.n271 B.n270 10.6151
R1146 B.n271 B.n186 10.6151
R1147 B.n275 B.n186 10.6151
R1148 B.n276 B.n275 10.6151
R1149 B.n277 B.n276 10.6151
R1150 B.n277 B.n184 10.6151
R1151 B.n281 B.n184 10.6151
R1152 B.n282 B.n281 10.6151
R1153 B.n283 B.n282 10.6151
R1154 B.n283 B.n182 10.6151
R1155 B.n287 B.n182 10.6151
R1156 B.n288 B.n287 10.6151
R1157 B.n289 B.n288 10.6151
R1158 B.n289 B.n180 10.6151
R1159 B.n293 B.n180 10.6151
R1160 B.n294 B.n293 10.6151
R1161 B.n295 B.n294 10.6151
R1162 B.n295 B.n178 10.6151
R1163 B.n299 B.n178 10.6151
R1164 B.n300 B.n299 10.6151
R1165 B.n301 B.n300 10.6151
R1166 B.n301 B.n176 10.6151
R1167 B.n305 B.n176 10.6151
R1168 B.n306 B.n305 10.6151
R1169 B.n307 B.n306 10.6151
R1170 B.n307 B.n174 10.6151
R1171 B.n311 B.n174 10.6151
R1172 B.n312 B.n311 10.6151
R1173 B.n313 B.n312 10.6151
R1174 B.n313 B.n172 10.6151
R1175 B.n317 B.n172 10.6151
R1176 B.n318 B.n317 10.6151
R1177 B.n319 B.n318 10.6151
R1178 B.n319 B.n170 10.6151
R1179 B.n323 B.n170 10.6151
R1180 B.n324 B.n323 10.6151
R1181 B.n325 B.n324 10.6151
R1182 B.n329 B.n168 10.6151
R1183 B.n330 B.n329 10.6151
R1184 B.n331 B.n330 10.6151
R1185 B.n331 B.n166 10.6151
R1186 B.n335 B.n166 10.6151
R1187 B.n336 B.n335 10.6151
R1188 B.n337 B.n336 10.6151
R1189 B.n337 B.n164 10.6151
R1190 B.n341 B.n164 10.6151
R1191 B.n342 B.n341 10.6151
R1192 B.n343 B.n342 10.6151
R1193 B.n343 B.n162 10.6151
R1194 B.n347 B.n162 10.6151
R1195 B.n348 B.n347 10.6151
R1196 B.n350 B.n158 10.6151
R1197 B.n354 B.n158 10.6151
R1198 B.n355 B.n354 10.6151
R1199 B.n356 B.n355 10.6151
R1200 B.n356 B.n156 10.6151
R1201 B.n360 B.n156 10.6151
R1202 B.n361 B.n360 10.6151
R1203 B.n365 B.n361 10.6151
R1204 B.n369 B.n154 10.6151
R1205 B.n370 B.n369 10.6151
R1206 B.n371 B.n370 10.6151
R1207 B.n371 B.n152 10.6151
R1208 B.n375 B.n152 10.6151
R1209 B.n376 B.n375 10.6151
R1210 B.n377 B.n376 10.6151
R1211 B.n377 B.n150 10.6151
R1212 B.n381 B.n150 10.6151
R1213 B.n382 B.n381 10.6151
R1214 B.n383 B.n382 10.6151
R1215 B.n383 B.n148 10.6151
R1216 B.n387 B.n148 10.6151
R1217 B.n388 B.n387 10.6151
R1218 B.n813 B.n0 8.11757
R1219 B.n813 B.n1 8.11757
R1220 B.n669 B.n668 6.5566
R1221 B.n656 B.n58 6.5566
R1222 B.n350 B.n349 6.5566
R1223 B.n365 B.n364 6.5566
R1224 B.n670 B.n669 4.05904
R1225 B.n653 B.n58 4.05904
R1226 B.n349 B.n348 4.05904
R1227 B.n364 B.n154 4.05904
R1228 VP.n31 VP.n30 161.3
R1229 VP.n32 VP.n27 161.3
R1230 VP.n34 VP.n33 161.3
R1231 VP.n35 VP.n26 161.3
R1232 VP.n37 VP.n36 161.3
R1233 VP.n38 VP.n25 161.3
R1234 VP.n40 VP.n39 161.3
R1235 VP.n41 VP.n24 161.3
R1236 VP.n44 VP.n43 161.3
R1237 VP.n45 VP.n23 161.3
R1238 VP.n47 VP.n46 161.3
R1239 VP.n48 VP.n22 161.3
R1240 VP.n50 VP.n49 161.3
R1241 VP.n51 VP.n21 161.3
R1242 VP.n53 VP.n52 161.3
R1243 VP.n54 VP.n20 161.3
R1244 VP.n57 VP.n56 161.3
R1245 VP.n58 VP.n19 161.3
R1246 VP.n60 VP.n59 161.3
R1247 VP.n61 VP.n18 161.3
R1248 VP.n63 VP.n62 161.3
R1249 VP.n64 VP.n17 161.3
R1250 VP.n66 VP.n65 161.3
R1251 VP.n67 VP.n16 161.3
R1252 VP.n122 VP.n0 161.3
R1253 VP.n121 VP.n120 161.3
R1254 VP.n119 VP.n1 161.3
R1255 VP.n118 VP.n117 161.3
R1256 VP.n116 VP.n2 161.3
R1257 VP.n115 VP.n114 161.3
R1258 VP.n113 VP.n3 161.3
R1259 VP.n112 VP.n111 161.3
R1260 VP.n109 VP.n4 161.3
R1261 VP.n108 VP.n107 161.3
R1262 VP.n106 VP.n5 161.3
R1263 VP.n105 VP.n104 161.3
R1264 VP.n103 VP.n6 161.3
R1265 VP.n102 VP.n101 161.3
R1266 VP.n100 VP.n7 161.3
R1267 VP.n99 VP.n98 161.3
R1268 VP.n96 VP.n8 161.3
R1269 VP.n95 VP.n94 161.3
R1270 VP.n93 VP.n9 161.3
R1271 VP.n92 VP.n91 161.3
R1272 VP.n90 VP.n10 161.3
R1273 VP.n89 VP.n88 161.3
R1274 VP.n87 VP.n11 161.3
R1275 VP.n86 VP.n85 161.3
R1276 VP.n83 VP.n12 161.3
R1277 VP.n82 VP.n81 161.3
R1278 VP.n80 VP.n13 161.3
R1279 VP.n79 VP.n78 161.3
R1280 VP.n77 VP.n14 161.3
R1281 VP.n76 VP.n75 161.3
R1282 VP.n74 VP.n15 161.3
R1283 VP.n73 VP.n72 161.3
R1284 VP.n71 VP.n70 60.1615
R1285 VP.n124 VP.n123 60.1615
R1286 VP.n69 VP.n68 60.1615
R1287 VP.n29 VP.n28 57.9068
R1288 VP.n91 VP.n90 56.5193
R1289 VP.n104 VP.n103 56.5193
R1290 VP.n49 VP.n48 56.5193
R1291 VP.n36 VP.n35 56.5193
R1292 VP.n70 VP.n69 52.7161
R1293 VP.n78 VP.n77 50.2061
R1294 VP.n117 VP.n116 50.2061
R1295 VP.n62 VP.n61 50.2061
R1296 VP.n28 VP.t5 50.0736
R1297 VP.n77 VP.n76 30.7807
R1298 VP.n117 VP.n1 30.7807
R1299 VP.n62 VP.n17 30.7807
R1300 VP.n72 VP.n15 24.4675
R1301 VP.n76 VP.n15 24.4675
R1302 VP.n78 VP.n13 24.4675
R1303 VP.n82 VP.n13 24.4675
R1304 VP.n83 VP.n82 24.4675
R1305 VP.n85 VP.n11 24.4675
R1306 VP.n89 VP.n11 24.4675
R1307 VP.n90 VP.n89 24.4675
R1308 VP.n91 VP.n9 24.4675
R1309 VP.n95 VP.n9 24.4675
R1310 VP.n96 VP.n95 24.4675
R1311 VP.n98 VP.n7 24.4675
R1312 VP.n102 VP.n7 24.4675
R1313 VP.n103 VP.n102 24.4675
R1314 VP.n104 VP.n5 24.4675
R1315 VP.n108 VP.n5 24.4675
R1316 VP.n109 VP.n108 24.4675
R1317 VP.n111 VP.n3 24.4675
R1318 VP.n115 VP.n3 24.4675
R1319 VP.n116 VP.n115 24.4675
R1320 VP.n121 VP.n1 24.4675
R1321 VP.n122 VP.n121 24.4675
R1322 VP.n66 VP.n17 24.4675
R1323 VP.n67 VP.n66 24.4675
R1324 VP.n49 VP.n21 24.4675
R1325 VP.n53 VP.n21 24.4675
R1326 VP.n54 VP.n53 24.4675
R1327 VP.n56 VP.n19 24.4675
R1328 VP.n60 VP.n19 24.4675
R1329 VP.n61 VP.n60 24.4675
R1330 VP.n36 VP.n25 24.4675
R1331 VP.n40 VP.n25 24.4675
R1332 VP.n41 VP.n40 24.4675
R1333 VP.n43 VP.n23 24.4675
R1334 VP.n47 VP.n23 24.4675
R1335 VP.n48 VP.n47 24.4675
R1336 VP.n30 VP.n27 24.4675
R1337 VP.n34 VP.n27 24.4675
R1338 VP.n35 VP.n34 24.4675
R1339 VP.n72 VP.n71 22.0208
R1340 VP.n123 VP.n122 22.0208
R1341 VP.n68 VP.n67 22.0208
R1342 VP.n71 VP.t8 17.8358
R1343 VP.n84 VP.t0 17.8358
R1344 VP.n97 VP.t3 17.8358
R1345 VP.n110 VP.t1 17.8358
R1346 VP.n123 VP.t6 17.8358
R1347 VP.n68 VP.t2 17.8358
R1348 VP.n55 VP.t4 17.8358
R1349 VP.n42 VP.t7 17.8358
R1350 VP.n29 VP.t9 17.8358
R1351 VP.n85 VP.n84 17.1274
R1352 VP.n110 VP.n109 17.1274
R1353 VP.n55 VP.n54 17.1274
R1354 VP.n30 VP.n29 17.1274
R1355 VP.n97 VP.n96 12.234
R1356 VP.n98 VP.n97 12.234
R1357 VP.n42 VP.n41 12.234
R1358 VP.n43 VP.n42 12.234
R1359 VP.n84 VP.n83 7.3406
R1360 VP.n111 VP.n110 7.3406
R1361 VP.n56 VP.n55 7.3406
R1362 VP.n31 VP.n28 2.61532
R1363 VP.n69 VP.n16 0.417535
R1364 VP.n73 VP.n70 0.417535
R1365 VP.n124 VP.n0 0.417535
R1366 VP VP.n124 0.394291
R1367 VP.n32 VP.n31 0.189894
R1368 VP.n33 VP.n32 0.189894
R1369 VP.n33 VP.n26 0.189894
R1370 VP.n37 VP.n26 0.189894
R1371 VP.n38 VP.n37 0.189894
R1372 VP.n39 VP.n38 0.189894
R1373 VP.n39 VP.n24 0.189894
R1374 VP.n44 VP.n24 0.189894
R1375 VP.n45 VP.n44 0.189894
R1376 VP.n46 VP.n45 0.189894
R1377 VP.n46 VP.n22 0.189894
R1378 VP.n50 VP.n22 0.189894
R1379 VP.n51 VP.n50 0.189894
R1380 VP.n52 VP.n51 0.189894
R1381 VP.n52 VP.n20 0.189894
R1382 VP.n57 VP.n20 0.189894
R1383 VP.n58 VP.n57 0.189894
R1384 VP.n59 VP.n58 0.189894
R1385 VP.n59 VP.n18 0.189894
R1386 VP.n63 VP.n18 0.189894
R1387 VP.n64 VP.n63 0.189894
R1388 VP.n65 VP.n64 0.189894
R1389 VP.n65 VP.n16 0.189894
R1390 VP.n74 VP.n73 0.189894
R1391 VP.n75 VP.n74 0.189894
R1392 VP.n75 VP.n14 0.189894
R1393 VP.n79 VP.n14 0.189894
R1394 VP.n80 VP.n79 0.189894
R1395 VP.n81 VP.n80 0.189894
R1396 VP.n81 VP.n12 0.189894
R1397 VP.n86 VP.n12 0.189894
R1398 VP.n87 VP.n86 0.189894
R1399 VP.n88 VP.n87 0.189894
R1400 VP.n88 VP.n10 0.189894
R1401 VP.n92 VP.n10 0.189894
R1402 VP.n93 VP.n92 0.189894
R1403 VP.n94 VP.n93 0.189894
R1404 VP.n94 VP.n8 0.189894
R1405 VP.n99 VP.n8 0.189894
R1406 VP.n100 VP.n99 0.189894
R1407 VP.n101 VP.n100 0.189894
R1408 VP.n101 VP.n6 0.189894
R1409 VP.n105 VP.n6 0.189894
R1410 VP.n106 VP.n105 0.189894
R1411 VP.n107 VP.n106 0.189894
R1412 VP.n107 VP.n4 0.189894
R1413 VP.n112 VP.n4 0.189894
R1414 VP.n113 VP.n112 0.189894
R1415 VP.n114 VP.n113 0.189894
R1416 VP.n114 VP.n2 0.189894
R1417 VP.n118 VP.n2 0.189894
R1418 VP.n119 VP.n118 0.189894
R1419 VP.n120 VP.n119 0.189894
R1420 VP.n120 VP.n0 0.189894
R1421 VDD1.n1 VDD1.t1 153.838
R1422 VDD1.n3 VDD1.t7 153.837
R1423 VDD1.n5 VDD1.n4 141.248
R1424 VDD1.n1 VDD1.n0 138.653
R1425 VDD1.n7 VDD1.n6 138.651
R1426 VDD1.n3 VDD1.n2 138.651
R1427 VDD1.n7 VDD1.n5 45.2595
R1428 VDD1.n6 VDD1.t4 11.651
R1429 VDD1.n6 VDD1.t3 11.651
R1430 VDD1.n0 VDD1.t8 11.651
R1431 VDD1.n0 VDD1.t9 11.651
R1432 VDD1.n4 VDD1.t5 11.651
R1433 VDD1.n4 VDD1.t2 11.651
R1434 VDD1.n2 VDD1.t6 11.651
R1435 VDD1.n2 VDD1.t0 11.651
R1436 VDD1 VDD1.n7 2.59317
R1437 VDD1 VDD1.n1 0.94231
R1438 VDD1.n5 VDD1.n3 0.828775
R1439 VTAIL.n11 VTAIL.t1 133.624
R1440 VTAIL.n17 VTAIL.t4 133.624
R1441 VTAIL.n2 VTAIL.t13 133.624
R1442 VTAIL.n16 VTAIL.t17 133.624
R1443 VTAIL.n15 VTAIL.n14 121.974
R1444 VTAIL.n13 VTAIL.n12 121.974
R1445 VTAIL.n10 VTAIL.n9 121.974
R1446 VTAIL.n8 VTAIL.n7 121.974
R1447 VTAIL.n19 VTAIL.n18 121.972
R1448 VTAIL.n1 VTAIL.n0 121.972
R1449 VTAIL.n4 VTAIL.n3 121.972
R1450 VTAIL.n6 VTAIL.n5 121.972
R1451 VTAIL.n8 VTAIL.n6 21.841
R1452 VTAIL.n17 VTAIL.n16 18.3065
R1453 VTAIL.n18 VTAIL.t0 11.651
R1454 VTAIL.n18 VTAIL.t3 11.651
R1455 VTAIL.n0 VTAIL.t7 11.651
R1456 VTAIL.n0 VTAIL.t6 11.651
R1457 VTAIL.n3 VTAIL.t16 11.651
R1458 VTAIL.n3 VTAIL.t18 11.651
R1459 VTAIL.n5 VTAIL.t11 11.651
R1460 VTAIL.n5 VTAIL.t19 11.651
R1461 VTAIL.n14 VTAIL.t12 11.651
R1462 VTAIL.n14 VTAIL.t15 11.651
R1463 VTAIL.n12 VTAIL.t14 11.651
R1464 VTAIL.n12 VTAIL.t10 11.651
R1465 VTAIL.n9 VTAIL.t9 11.651
R1466 VTAIL.n9 VTAIL.t5 11.651
R1467 VTAIL.n7 VTAIL.t8 11.651
R1468 VTAIL.n7 VTAIL.t2 11.651
R1469 VTAIL.n10 VTAIL.n8 3.53498
R1470 VTAIL.n11 VTAIL.n10 3.53498
R1471 VTAIL.n15 VTAIL.n13 3.53498
R1472 VTAIL.n16 VTAIL.n15 3.53498
R1473 VTAIL.n6 VTAIL.n4 3.53498
R1474 VTAIL.n4 VTAIL.n2 3.53498
R1475 VTAIL.n19 VTAIL.n17 3.53498
R1476 VTAIL VTAIL.n1 2.70955
R1477 VTAIL.n13 VTAIL.n11 2.23757
R1478 VTAIL.n2 VTAIL.n1 2.23757
R1479 VTAIL VTAIL.n19 0.825931
R1480 VN.n105 VN.n54 161.3
R1481 VN.n104 VN.n103 161.3
R1482 VN.n102 VN.n55 161.3
R1483 VN.n101 VN.n100 161.3
R1484 VN.n99 VN.n56 161.3
R1485 VN.n98 VN.n97 161.3
R1486 VN.n96 VN.n57 161.3
R1487 VN.n95 VN.n94 161.3
R1488 VN.n92 VN.n58 161.3
R1489 VN.n91 VN.n90 161.3
R1490 VN.n89 VN.n59 161.3
R1491 VN.n88 VN.n87 161.3
R1492 VN.n86 VN.n60 161.3
R1493 VN.n85 VN.n84 161.3
R1494 VN.n83 VN.n61 161.3
R1495 VN.n82 VN.n81 161.3
R1496 VN.n79 VN.n62 161.3
R1497 VN.n78 VN.n77 161.3
R1498 VN.n76 VN.n63 161.3
R1499 VN.n75 VN.n74 161.3
R1500 VN.n73 VN.n64 161.3
R1501 VN.n72 VN.n71 161.3
R1502 VN.n70 VN.n65 161.3
R1503 VN.n69 VN.n68 161.3
R1504 VN.n51 VN.n0 161.3
R1505 VN.n50 VN.n49 161.3
R1506 VN.n48 VN.n1 161.3
R1507 VN.n47 VN.n46 161.3
R1508 VN.n45 VN.n2 161.3
R1509 VN.n44 VN.n43 161.3
R1510 VN.n42 VN.n3 161.3
R1511 VN.n41 VN.n40 161.3
R1512 VN.n38 VN.n4 161.3
R1513 VN.n37 VN.n36 161.3
R1514 VN.n35 VN.n5 161.3
R1515 VN.n34 VN.n33 161.3
R1516 VN.n32 VN.n6 161.3
R1517 VN.n31 VN.n30 161.3
R1518 VN.n29 VN.n7 161.3
R1519 VN.n28 VN.n27 161.3
R1520 VN.n25 VN.n8 161.3
R1521 VN.n24 VN.n23 161.3
R1522 VN.n22 VN.n9 161.3
R1523 VN.n21 VN.n20 161.3
R1524 VN.n19 VN.n10 161.3
R1525 VN.n18 VN.n17 161.3
R1526 VN.n16 VN.n11 161.3
R1527 VN.n15 VN.n14 161.3
R1528 VN.n53 VN.n52 60.1615
R1529 VN.n107 VN.n106 60.1615
R1530 VN.n13 VN.n12 57.9067
R1531 VN.n67 VN.n66 57.9067
R1532 VN.n20 VN.n19 56.5193
R1533 VN.n33 VN.n32 56.5193
R1534 VN.n74 VN.n73 56.5193
R1535 VN.n87 VN.n86 56.5193
R1536 VN VN.n107 52.7541
R1537 VN.n46 VN.n45 50.2061
R1538 VN.n100 VN.n99 50.2061
R1539 VN.n12 VN.t4 50.074
R1540 VN.n66 VN.t1 50.074
R1541 VN.n46 VN.n1 30.7807
R1542 VN.n100 VN.n55 30.7807
R1543 VN.n14 VN.n11 24.4675
R1544 VN.n18 VN.n11 24.4675
R1545 VN.n19 VN.n18 24.4675
R1546 VN.n20 VN.n9 24.4675
R1547 VN.n24 VN.n9 24.4675
R1548 VN.n25 VN.n24 24.4675
R1549 VN.n27 VN.n7 24.4675
R1550 VN.n31 VN.n7 24.4675
R1551 VN.n32 VN.n31 24.4675
R1552 VN.n33 VN.n5 24.4675
R1553 VN.n37 VN.n5 24.4675
R1554 VN.n38 VN.n37 24.4675
R1555 VN.n40 VN.n3 24.4675
R1556 VN.n44 VN.n3 24.4675
R1557 VN.n45 VN.n44 24.4675
R1558 VN.n50 VN.n1 24.4675
R1559 VN.n51 VN.n50 24.4675
R1560 VN.n73 VN.n72 24.4675
R1561 VN.n72 VN.n65 24.4675
R1562 VN.n68 VN.n65 24.4675
R1563 VN.n86 VN.n85 24.4675
R1564 VN.n85 VN.n61 24.4675
R1565 VN.n81 VN.n61 24.4675
R1566 VN.n79 VN.n78 24.4675
R1567 VN.n78 VN.n63 24.4675
R1568 VN.n74 VN.n63 24.4675
R1569 VN.n99 VN.n98 24.4675
R1570 VN.n98 VN.n57 24.4675
R1571 VN.n94 VN.n57 24.4675
R1572 VN.n92 VN.n91 24.4675
R1573 VN.n91 VN.n59 24.4675
R1574 VN.n87 VN.n59 24.4675
R1575 VN.n105 VN.n104 24.4675
R1576 VN.n104 VN.n55 24.4675
R1577 VN.n52 VN.n51 22.0208
R1578 VN.n106 VN.n105 22.0208
R1579 VN.n13 VN.t9 17.8358
R1580 VN.n26 VN.t6 17.8358
R1581 VN.n39 VN.t2 17.8358
R1582 VN.n52 VN.t0 17.8358
R1583 VN.n67 VN.t3 17.8358
R1584 VN.n80 VN.t7 17.8358
R1585 VN.n93 VN.t8 17.8358
R1586 VN.n106 VN.t5 17.8358
R1587 VN.n14 VN.n13 17.1274
R1588 VN.n39 VN.n38 17.1274
R1589 VN.n68 VN.n67 17.1274
R1590 VN.n93 VN.n92 17.1274
R1591 VN.n26 VN.n25 12.234
R1592 VN.n27 VN.n26 12.234
R1593 VN.n81 VN.n80 12.234
R1594 VN.n80 VN.n79 12.234
R1595 VN.n40 VN.n39 7.3406
R1596 VN.n94 VN.n93 7.3406
R1597 VN.n69 VN.n66 2.61535
R1598 VN.n15 VN.n12 2.61535
R1599 VN.n107 VN.n54 0.417535
R1600 VN.n53 VN.n0 0.417535
R1601 VN VN.n53 0.394291
R1602 VN.n103 VN.n54 0.189894
R1603 VN.n103 VN.n102 0.189894
R1604 VN.n102 VN.n101 0.189894
R1605 VN.n101 VN.n56 0.189894
R1606 VN.n97 VN.n56 0.189894
R1607 VN.n97 VN.n96 0.189894
R1608 VN.n96 VN.n95 0.189894
R1609 VN.n95 VN.n58 0.189894
R1610 VN.n90 VN.n58 0.189894
R1611 VN.n90 VN.n89 0.189894
R1612 VN.n89 VN.n88 0.189894
R1613 VN.n88 VN.n60 0.189894
R1614 VN.n84 VN.n60 0.189894
R1615 VN.n84 VN.n83 0.189894
R1616 VN.n83 VN.n82 0.189894
R1617 VN.n82 VN.n62 0.189894
R1618 VN.n77 VN.n62 0.189894
R1619 VN.n77 VN.n76 0.189894
R1620 VN.n76 VN.n75 0.189894
R1621 VN.n75 VN.n64 0.189894
R1622 VN.n71 VN.n64 0.189894
R1623 VN.n71 VN.n70 0.189894
R1624 VN.n70 VN.n69 0.189894
R1625 VN.n16 VN.n15 0.189894
R1626 VN.n17 VN.n16 0.189894
R1627 VN.n17 VN.n10 0.189894
R1628 VN.n21 VN.n10 0.189894
R1629 VN.n22 VN.n21 0.189894
R1630 VN.n23 VN.n22 0.189894
R1631 VN.n23 VN.n8 0.189894
R1632 VN.n28 VN.n8 0.189894
R1633 VN.n29 VN.n28 0.189894
R1634 VN.n30 VN.n29 0.189894
R1635 VN.n30 VN.n6 0.189894
R1636 VN.n34 VN.n6 0.189894
R1637 VN.n35 VN.n34 0.189894
R1638 VN.n36 VN.n35 0.189894
R1639 VN.n36 VN.n4 0.189894
R1640 VN.n41 VN.n4 0.189894
R1641 VN.n42 VN.n41 0.189894
R1642 VN.n43 VN.n42 0.189894
R1643 VN.n43 VN.n2 0.189894
R1644 VN.n47 VN.n2 0.189894
R1645 VN.n48 VN.n47 0.189894
R1646 VN.n49 VN.n48 0.189894
R1647 VN.n49 VN.n0 0.189894
R1648 VDD2.n1 VDD2.t5 153.837
R1649 VDD2.n4 VDD2.t4 150.303
R1650 VDD2.n3 VDD2.n2 141.248
R1651 VDD2 VDD2.n7 141.244
R1652 VDD2.n6 VDD2.n5 138.653
R1653 VDD2.n1 VDD2.n0 138.651
R1654 VDD2.n4 VDD2.n3 42.9093
R1655 VDD2.n7 VDD2.t6 11.651
R1656 VDD2.n7 VDD2.t8 11.651
R1657 VDD2.n5 VDD2.t1 11.651
R1658 VDD2.n5 VDD2.t2 11.651
R1659 VDD2.n2 VDD2.t7 11.651
R1660 VDD2.n2 VDD2.t9 11.651
R1661 VDD2.n0 VDD2.t0 11.651
R1662 VDD2.n0 VDD2.t3 11.651
R1663 VDD2.n6 VDD2.n4 3.53498
R1664 VDD2 VDD2.n6 0.94231
R1665 VDD2.n3 VDD2.n1 0.828775
C0 B VDD1 2.19002f
C1 VN VDD1 0.161515f
C2 w_n5890_n1526# VTAIL 2.10981f
C3 VN B 1.51065f
C4 VDD2 VTAIL 7.47035f
C5 VTAIL VP 5.05144f
C6 VTAIL VDD1 7.40918f
C7 B VTAIL 1.88255f
C8 VN VTAIL 5.03721f
C9 w_n5890_n1526# VDD2 2.80427f
C10 w_n5890_n1526# VP 13.6013f
C11 VDD2 VP 0.738956f
C12 w_n5890_n1526# VDD1 2.60047f
C13 VDD2 VDD1 2.93636f
C14 VP VDD1 3.64014f
C15 B w_n5890_n1526# 9.99831f
C16 B VDD2 2.35381f
C17 VN w_n5890_n1526# 12.8335f
C18 B VP 2.81219f
C19 VN VDD2 3.06708f
C20 VN VP 8.42968f
C21 VDD2 VSUBS 2.575436f
C22 VDD1 VSUBS 2.283281f
C23 VTAIL VSUBS 0.738709f
C24 VN VSUBS 9.79093f
C25 VP VSUBS 5.028906f
C26 B VSUBS 5.648806f
C27 w_n5890_n1526# VSUBS 0.114007p
C28 VDD2.t5 VSUBS 0.683906f
C29 VDD2.t0 VSUBS 0.090164f
C30 VDD2.t3 VSUBS 0.090164f
C31 VDD2.n0 VSUBS 0.462246f
C32 VDD2.n1 VSUBS 2.08198f
C33 VDD2.t7 VSUBS 0.090164f
C34 VDD2.t9 VSUBS 0.090164f
C35 VDD2.n2 VSUBS 0.486582f
C36 VDD2.n3 VSUBS 5.01234f
C37 VDD2.t4 VSUBS 0.660246f
C38 VDD2.n4 VSUBS 4.787951f
C39 VDD2.t1 VSUBS 0.090164f
C40 VDD2.t2 VSUBS 0.090164f
C41 VDD2.n5 VSUBS 0.462247f
C42 VDD2.n6 VSUBS 1.08959f
C43 VDD2.t6 VSUBS 0.090164f
C44 VDD2.t8 VSUBS 0.090164f
C45 VDD2.n7 VSUBS 0.486541f
C46 VN.n0 VSUBS 0.079029f
C47 VN.t0 VSUBS 1.0905f
C48 VN.n1 VSUBS 0.08417f
C49 VN.n2 VSUBS 0.042014f
C50 VN.n3 VSUBS 0.078304f
C51 VN.n4 VSUBS 0.042014f
C52 VN.t2 VSUBS 1.0905f
C53 VN.n5 VSUBS 0.078304f
C54 VN.n6 VSUBS 0.042014f
C55 VN.n7 VSUBS 0.078304f
C56 VN.n8 VSUBS 0.042014f
C57 VN.t6 VSUBS 1.0905f
C58 VN.n9 VSUBS 0.078304f
C59 VN.n10 VSUBS 0.042014f
C60 VN.n11 VSUBS 0.078304f
C61 VN.t4 VSUBS 1.59164f
C62 VN.n12 VSUBS 0.649749f
C63 VN.t9 VSUBS 1.0905f
C64 VN.n13 VSUBS 0.609885f
C65 VN.n14 VSUBS 0.066707f
C66 VN.n15 VSUBS 0.545926f
C67 VN.n16 VSUBS 0.042014f
C68 VN.n17 VSUBS 0.042014f
C69 VN.n18 VSUBS 0.078304f
C70 VN.n19 VSUBS 0.05548f
C71 VN.n20 VSUBS 0.067188f
C72 VN.n21 VSUBS 0.042014f
C73 VN.n22 VSUBS 0.042014f
C74 VN.n23 VSUBS 0.042014f
C75 VN.n24 VSUBS 0.078304f
C76 VN.n25 VSUBS 0.058975f
C77 VN.n26 VSUBS 0.451482f
C78 VN.n27 VSUBS 0.058975f
C79 VN.n28 VSUBS 0.042014f
C80 VN.n29 VSUBS 0.042014f
C81 VN.n30 VSUBS 0.042014f
C82 VN.n31 VSUBS 0.078304f
C83 VN.n32 VSUBS 0.067188f
C84 VN.n33 VSUBS 0.05548f
C85 VN.n34 VSUBS 0.042014f
C86 VN.n35 VSUBS 0.042014f
C87 VN.n36 VSUBS 0.042014f
C88 VN.n37 VSUBS 0.078304f
C89 VN.n38 VSUBS 0.066707f
C90 VN.n39 VSUBS 0.451482f
C91 VN.n40 VSUBS 0.051243f
C92 VN.n41 VSUBS 0.042014f
C93 VN.n42 VSUBS 0.042014f
C94 VN.n43 VSUBS 0.042014f
C95 VN.n44 VSUBS 0.078304f
C96 VN.n45 VSUBS 0.077112f
C97 VN.n46 VSUBS 0.03969f
C98 VN.n47 VSUBS 0.042014f
C99 VN.n48 VSUBS 0.042014f
C100 VN.n49 VSUBS 0.042014f
C101 VN.n50 VSUBS 0.078304f
C102 VN.n51 VSUBS 0.074438f
C103 VN.n52 VSUBS 0.633789f
C104 VN.n53 VSUBS 0.125976f
C105 VN.n54 VSUBS 0.079029f
C106 VN.t5 VSUBS 1.0905f
C107 VN.n55 VSUBS 0.08417f
C108 VN.n56 VSUBS 0.042014f
C109 VN.n57 VSUBS 0.078304f
C110 VN.n58 VSUBS 0.042014f
C111 VN.t8 VSUBS 1.0905f
C112 VN.n59 VSUBS 0.078304f
C113 VN.n60 VSUBS 0.042014f
C114 VN.n61 VSUBS 0.078304f
C115 VN.n62 VSUBS 0.042014f
C116 VN.t7 VSUBS 1.0905f
C117 VN.n63 VSUBS 0.078304f
C118 VN.n64 VSUBS 0.042014f
C119 VN.n65 VSUBS 0.078304f
C120 VN.t1 VSUBS 1.59164f
C121 VN.n66 VSUBS 0.649749f
C122 VN.t3 VSUBS 1.0905f
C123 VN.n67 VSUBS 0.609885f
C124 VN.n68 VSUBS 0.066707f
C125 VN.n69 VSUBS 0.545926f
C126 VN.n70 VSUBS 0.042014f
C127 VN.n71 VSUBS 0.042014f
C128 VN.n72 VSUBS 0.078304f
C129 VN.n73 VSUBS 0.05548f
C130 VN.n74 VSUBS 0.067188f
C131 VN.n75 VSUBS 0.042014f
C132 VN.n76 VSUBS 0.042014f
C133 VN.n77 VSUBS 0.042014f
C134 VN.n78 VSUBS 0.078304f
C135 VN.n79 VSUBS 0.058975f
C136 VN.n80 VSUBS 0.451482f
C137 VN.n81 VSUBS 0.058975f
C138 VN.n82 VSUBS 0.042014f
C139 VN.n83 VSUBS 0.042014f
C140 VN.n84 VSUBS 0.042014f
C141 VN.n85 VSUBS 0.078304f
C142 VN.n86 VSUBS 0.067188f
C143 VN.n87 VSUBS 0.05548f
C144 VN.n88 VSUBS 0.042014f
C145 VN.n89 VSUBS 0.042014f
C146 VN.n90 VSUBS 0.042014f
C147 VN.n91 VSUBS 0.078304f
C148 VN.n92 VSUBS 0.066707f
C149 VN.n93 VSUBS 0.451482f
C150 VN.n94 VSUBS 0.051243f
C151 VN.n95 VSUBS 0.042014f
C152 VN.n96 VSUBS 0.042014f
C153 VN.n97 VSUBS 0.042014f
C154 VN.n98 VSUBS 0.078304f
C155 VN.n99 VSUBS 0.077112f
C156 VN.n100 VSUBS 0.03969f
C157 VN.n101 VSUBS 0.042014f
C158 VN.n102 VSUBS 0.042014f
C159 VN.n103 VSUBS 0.042014f
C160 VN.n104 VSUBS 0.078304f
C161 VN.n105 VSUBS 0.074438f
C162 VN.n106 VSUBS 0.633789f
C163 VN.n107 VSUBS 2.63272f
C164 VTAIL.t7 VSUBS 0.08659f
C165 VTAIL.t6 VSUBS 0.08659f
C166 VTAIL.n0 VSUBS 0.37932f
C167 VTAIL.n1 VSUBS 1.11709f
C168 VTAIL.t13 VSUBS 0.569361f
C169 VTAIL.n2 VSUBS 1.26766f
C170 VTAIL.t16 VSUBS 0.08659f
C171 VTAIL.t18 VSUBS 0.08659f
C172 VTAIL.n3 VSUBS 0.37932f
C173 VTAIL.n4 VSUBS 1.38573f
C174 VTAIL.t11 VSUBS 0.08659f
C175 VTAIL.t19 VSUBS 0.08659f
C176 VTAIL.n5 VSUBS 0.37932f
C177 VTAIL.n6 VSUBS 2.6709f
C178 VTAIL.t8 VSUBS 0.08659f
C179 VTAIL.t2 VSUBS 0.08659f
C180 VTAIL.n7 VSUBS 0.379321f
C181 VTAIL.n8 VSUBS 2.67089f
C182 VTAIL.t9 VSUBS 0.08659f
C183 VTAIL.t5 VSUBS 0.08659f
C184 VTAIL.n9 VSUBS 0.379321f
C185 VTAIL.n10 VSUBS 1.38573f
C186 VTAIL.t1 VSUBS 0.569362f
C187 VTAIL.n11 VSUBS 1.26766f
C188 VTAIL.t14 VSUBS 0.08659f
C189 VTAIL.t10 VSUBS 0.08659f
C190 VTAIL.n12 VSUBS 0.379321f
C191 VTAIL.n13 VSUBS 1.22154f
C192 VTAIL.t12 VSUBS 0.08659f
C193 VTAIL.t15 VSUBS 0.08659f
C194 VTAIL.n14 VSUBS 0.379321f
C195 VTAIL.n15 VSUBS 1.38573f
C196 VTAIL.t17 VSUBS 0.569361f
C197 VTAIL.n16 VSUBS 2.26972f
C198 VTAIL.t4 VSUBS 0.569361f
C199 VTAIL.n17 VSUBS 2.26972f
C200 VTAIL.t0 VSUBS 0.08659f
C201 VTAIL.t3 VSUBS 0.08659f
C202 VTAIL.n18 VSUBS 0.37932f
C203 VTAIL.n19 VSUBS 1.0429f
C204 VDD1.t1 VSUBS 0.678428f
C205 VDD1.t8 VSUBS 0.089441f
C206 VDD1.t9 VSUBS 0.089441f
C207 VDD1.n0 VSUBS 0.458544f
C208 VDD1.n1 VSUBS 2.079f
C209 VDD1.t7 VSUBS 0.678426f
C210 VDD1.t6 VSUBS 0.089441f
C211 VDD1.t0 VSUBS 0.089441f
C212 VDD1.n2 VSUBS 0.458542f
C213 VDD1.n3 VSUBS 2.0653f
C214 VDD1.t5 VSUBS 0.089441f
C215 VDD1.t2 VSUBS 0.089441f
C216 VDD1.n4 VSUBS 0.482683f
C217 VDD1.n5 VSUBS 5.21239f
C218 VDD1.t4 VSUBS 0.089441f
C219 VDD1.t3 VSUBS 0.089441f
C220 VDD1.n6 VSUBS 0.458541f
C221 VDD1.n7 VSUBS 4.9506f
C222 VP.n0 VSUBS 0.09054f
C223 VP.t6 VSUBS 1.24934f
C224 VP.n1 VSUBS 0.096429f
C225 VP.n2 VSUBS 0.048134f
C226 VP.n3 VSUBS 0.08971f
C227 VP.n4 VSUBS 0.048134f
C228 VP.t1 VSUBS 1.24934f
C229 VP.n5 VSUBS 0.08971f
C230 VP.n6 VSUBS 0.048134f
C231 VP.n7 VSUBS 0.08971f
C232 VP.n8 VSUBS 0.048134f
C233 VP.t3 VSUBS 1.24934f
C234 VP.n9 VSUBS 0.08971f
C235 VP.n10 VSUBS 0.048134f
C236 VP.n11 VSUBS 0.08971f
C237 VP.n12 VSUBS 0.048134f
C238 VP.t0 VSUBS 1.24934f
C239 VP.n13 VSUBS 0.08971f
C240 VP.n14 VSUBS 0.048134f
C241 VP.n15 VSUBS 0.08971f
C242 VP.n16 VSUBS 0.09054f
C243 VP.t2 VSUBS 1.24934f
C244 VP.n17 VSUBS 0.096429f
C245 VP.n18 VSUBS 0.048134f
C246 VP.n19 VSUBS 0.08971f
C247 VP.n20 VSUBS 0.048134f
C248 VP.t4 VSUBS 1.24934f
C249 VP.n21 VSUBS 0.08971f
C250 VP.n22 VSUBS 0.048134f
C251 VP.n23 VSUBS 0.08971f
C252 VP.n24 VSUBS 0.048134f
C253 VP.t7 VSUBS 1.24934f
C254 VP.n25 VSUBS 0.08971f
C255 VP.n26 VSUBS 0.048134f
C256 VP.n27 VSUBS 0.08971f
C257 VP.t5 VSUBS 1.82346f
C258 VP.n28 VSUBS 0.744391f
C259 VP.t9 VSUBS 1.24934f
C260 VP.n29 VSUBS 0.698718f
C261 VP.n30 VSUBS 0.076423f
C262 VP.n31 VSUBS 0.625443f
C263 VP.n32 VSUBS 0.048134f
C264 VP.n33 VSUBS 0.048134f
C265 VP.n34 VSUBS 0.08971f
C266 VP.n35 VSUBS 0.063561f
C267 VP.n36 VSUBS 0.076974f
C268 VP.n37 VSUBS 0.048134f
C269 VP.n38 VSUBS 0.048134f
C270 VP.n39 VSUBS 0.048134f
C271 VP.n40 VSUBS 0.08971f
C272 VP.n41 VSUBS 0.067565f
C273 VP.n42 VSUBS 0.517242f
C274 VP.n43 VSUBS 0.067565f
C275 VP.n44 VSUBS 0.048134f
C276 VP.n45 VSUBS 0.048134f
C277 VP.n46 VSUBS 0.048134f
C278 VP.n47 VSUBS 0.08971f
C279 VP.n48 VSUBS 0.076974f
C280 VP.n49 VSUBS 0.063561f
C281 VP.n50 VSUBS 0.048134f
C282 VP.n51 VSUBS 0.048134f
C283 VP.n52 VSUBS 0.048134f
C284 VP.n53 VSUBS 0.08971f
C285 VP.n54 VSUBS 0.076423f
C286 VP.n55 VSUBS 0.517242f
C287 VP.n56 VSUBS 0.058707f
C288 VP.n57 VSUBS 0.048134f
C289 VP.n58 VSUBS 0.048134f
C290 VP.n59 VSUBS 0.048134f
C291 VP.n60 VSUBS 0.08971f
C292 VP.n61 VSUBS 0.088343f
C293 VP.n62 VSUBS 0.045471f
C294 VP.n63 VSUBS 0.048134f
C295 VP.n64 VSUBS 0.048134f
C296 VP.n65 VSUBS 0.048134f
C297 VP.n66 VSUBS 0.08971f
C298 VP.n67 VSUBS 0.085281f
C299 VP.n68 VSUBS 0.726103f
C300 VP.n69 VSUBS 3.00406f
C301 VP.n70 VSUBS 3.03688f
C302 VP.t8 VSUBS 1.24934f
C303 VP.n71 VSUBS 0.726103f
C304 VP.n72 VSUBS 0.085281f
C305 VP.n73 VSUBS 0.09054f
C306 VP.n74 VSUBS 0.048134f
C307 VP.n75 VSUBS 0.048134f
C308 VP.n76 VSUBS 0.096429f
C309 VP.n77 VSUBS 0.045471f
C310 VP.n78 VSUBS 0.088343f
C311 VP.n79 VSUBS 0.048134f
C312 VP.n80 VSUBS 0.048134f
C313 VP.n81 VSUBS 0.048134f
C314 VP.n82 VSUBS 0.08971f
C315 VP.n83 VSUBS 0.058707f
C316 VP.n84 VSUBS 0.517242f
C317 VP.n85 VSUBS 0.076423f
C318 VP.n86 VSUBS 0.048134f
C319 VP.n87 VSUBS 0.048134f
C320 VP.n88 VSUBS 0.048134f
C321 VP.n89 VSUBS 0.08971f
C322 VP.n90 VSUBS 0.063561f
C323 VP.n91 VSUBS 0.076974f
C324 VP.n92 VSUBS 0.048134f
C325 VP.n93 VSUBS 0.048134f
C326 VP.n94 VSUBS 0.048134f
C327 VP.n95 VSUBS 0.08971f
C328 VP.n96 VSUBS 0.067565f
C329 VP.n97 VSUBS 0.517242f
C330 VP.n98 VSUBS 0.067565f
C331 VP.n99 VSUBS 0.048134f
C332 VP.n100 VSUBS 0.048134f
C333 VP.n101 VSUBS 0.048134f
C334 VP.n102 VSUBS 0.08971f
C335 VP.n103 VSUBS 0.076974f
C336 VP.n104 VSUBS 0.063561f
C337 VP.n105 VSUBS 0.048134f
C338 VP.n106 VSUBS 0.048134f
C339 VP.n107 VSUBS 0.048134f
C340 VP.n108 VSUBS 0.08971f
C341 VP.n109 VSUBS 0.076423f
C342 VP.n110 VSUBS 0.517242f
C343 VP.n111 VSUBS 0.058707f
C344 VP.n112 VSUBS 0.048134f
C345 VP.n113 VSUBS 0.048134f
C346 VP.n114 VSUBS 0.048134f
C347 VP.n115 VSUBS 0.08971f
C348 VP.n116 VSUBS 0.088343f
C349 VP.n117 VSUBS 0.045471f
C350 VP.n118 VSUBS 0.048134f
C351 VP.n119 VSUBS 0.048134f
C352 VP.n120 VSUBS 0.048134f
C353 VP.n121 VSUBS 0.08971f
C354 VP.n122 VSUBS 0.085281f
C355 VP.n123 VSUBS 0.726103f
C356 VP.n124 VSUBS 0.144325f
C357 B.n0 VSUBS 0.011763f
C358 B.n1 VSUBS 0.011763f
C359 B.n2 VSUBS 0.017397f
C360 B.n3 VSUBS 0.013331f
C361 B.n4 VSUBS 0.013331f
C362 B.n5 VSUBS 0.013331f
C363 B.n6 VSUBS 0.013331f
C364 B.n7 VSUBS 0.013331f
C365 B.n8 VSUBS 0.013331f
C366 B.n9 VSUBS 0.013331f
C367 B.n10 VSUBS 0.013331f
C368 B.n11 VSUBS 0.013331f
C369 B.n12 VSUBS 0.013331f
C370 B.n13 VSUBS 0.013331f
C371 B.n14 VSUBS 0.013331f
C372 B.n15 VSUBS 0.013331f
C373 B.n16 VSUBS 0.013331f
C374 B.n17 VSUBS 0.013331f
C375 B.n18 VSUBS 0.013331f
C376 B.n19 VSUBS 0.013331f
C377 B.n20 VSUBS 0.013331f
C378 B.n21 VSUBS 0.013331f
C379 B.n22 VSUBS 0.013331f
C380 B.n23 VSUBS 0.013331f
C381 B.n24 VSUBS 0.013331f
C382 B.n25 VSUBS 0.013331f
C383 B.n26 VSUBS 0.013331f
C384 B.n27 VSUBS 0.013331f
C385 B.n28 VSUBS 0.013331f
C386 B.n29 VSUBS 0.013331f
C387 B.n30 VSUBS 0.013331f
C388 B.n31 VSUBS 0.013331f
C389 B.n32 VSUBS 0.013331f
C390 B.n33 VSUBS 0.013331f
C391 B.n34 VSUBS 0.013331f
C392 B.n35 VSUBS 0.013331f
C393 B.n36 VSUBS 0.013331f
C394 B.n37 VSUBS 0.013331f
C395 B.n38 VSUBS 0.013331f
C396 B.n39 VSUBS 0.013331f
C397 B.n40 VSUBS 0.013331f
C398 B.n41 VSUBS 0.013331f
C399 B.n42 VSUBS 0.030624f
C400 B.n43 VSUBS 0.013331f
C401 B.n44 VSUBS 0.013331f
C402 B.n45 VSUBS 0.013331f
C403 B.n46 VSUBS 0.013331f
C404 B.n47 VSUBS 0.013331f
C405 B.n48 VSUBS 0.013331f
C406 B.n49 VSUBS 0.013331f
C407 B.t10 VSUBS 0.12556f
C408 B.t11 VSUBS 0.165768f
C409 B.t9 VSUBS 0.984419f
C410 B.n50 VSUBS 0.168375f
C411 B.n51 VSUBS 0.131007f
C412 B.n52 VSUBS 0.013331f
C413 B.n53 VSUBS 0.013331f
C414 B.n54 VSUBS 0.013331f
C415 B.n55 VSUBS 0.013331f
C416 B.t4 VSUBS 0.12556f
C417 B.t5 VSUBS 0.165768f
C418 B.t3 VSUBS 0.984419f
C419 B.n56 VSUBS 0.168375f
C420 B.n57 VSUBS 0.131007f
C421 B.n58 VSUBS 0.030887f
C422 B.n59 VSUBS 0.013331f
C423 B.n60 VSUBS 0.013331f
C424 B.n61 VSUBS 0.013331f
C425 B.n62 VSUBS 0.013331f
C426 B.n63 VSUBS 0.013331f
C427 B.n64 VSUBS 0.013331f
C428 B.n65 VSUBS 0.013331f
C429 B.n66 VSUBS 0.028583f
C430 B.n67 VSUBS 0.013331f
C431 B.n68 VSUBS 0.013331f
C432 B.n69 VSUBS 0.013331f
C433 B.n70 VSUBS 0.013331f
C434 B.n71 VSUBS 0.013331f
C435 B.n72 VSUBS 0.013331f
C436 B.n73 VSUBS 0.013331f
C437 B.n74 VSUBS 0.013331f
C438 B.n75 VSUBS 0.013331f
C439 B.n76 VSUBS 0.013331f
C440 B.n77 VSUBS 0.013331f
C441 B.n78 VSUBS 0.013331f
C442 B.n79 VSUBS 0.013331f
C443 B.n80 VSUBS 0.013331f
C444 B.n81 VSUBS 0.013331f
C445 B.n82 VSUBS 0.013331f
C446 B.n83 VSUBS 0.013331f
C447 B.n84 VSUBS 0.013331f
C448 B.n85 VSUBS 0.013331f
C449 B.n86 VSUBS 0.013331f
C450 B.n87 VSUBS 0.013331f
C451 B.n88 VSUBS 0.013331f
C452 B.n89 VSUBS 0.013331f
C453 B.n90 VSUBS 0.013331f
C454 B.n91 VSUBS 0.013331f
C455 B.n92 VSUBS 0.013331f
C456 B.n93 VSUBS 0.013331f
C457 B.n94 VSUBS 0.013331f
C458 B.n95 VSUBS 0.013331f
C459 B.n96 VSUBS 0.013331f
C460 B.n97 VSUBS 0.013331f
C461 B.n98 VSUBS 0.013331f
C462 B.n99 VSUBS 0.013331f
C463 B.n100 VSUBS 0.013331f
C464 B.n101 VSUBS 0.013331f
C465 B.n102 VSUBS 0.013331f
C466 B.n103 VSUBS 0.013331f
C467 B.n104 VSUBS 0.013331f
C468 B.n105 VSUBS 0.013331f
C469 B.n106 VSUBS 0.013331f
C470 B.n107 VSUBS 0.013331f
C471 B.n108 VSUBS 0.013331f
C472 B.n109 VSUBS 0.013331f
C473 B.n110 VSUBS 0.013331f
C474 B.n111 VSUBS 0.013331f
C475 B.n112 VSUBS 0.013331f
C476 B.n113 VSUBS 0.013331f
C477 B.n114 VSUBS 0.013331f
C478 B.n115 VSUBS 0.013331f
C479 B.n116 VSUBS 0.013331f
C480 B.n117 VSUBS 0.013331f
C481 B.n118 VSUBS 0.013331f
C482 B.n119 VSUBS 0.013331f
C483 B.n120 VSUBS 0.013331f
C484 B.n121 VSUBS 0.013331f
C485 B.n122 VSUBS 0.013331f
C486 B.n123 VSUBS 0.013331f
C487 B.n124 VSUBS 0.013331f
C488 B.n125 VSUBS 0.013331f
C489 B.n126 VSUBS 0.013331f
C490 B.n127 VSUBS 0.013331f
C491 B.n128 VSUBS 0.013331f
C492 B.n129 VSUBS 0.013331f
C493 B.n130 VSUBS 0.013331f
C494 B.n131 VSUBS 0.013331f
C495 B.n132 VSUBS 0.013331f
C496 B.n133 VSUBS 0.013331f
C497 B.n134 VSUBS 0.013331f
C498 B.n135 VSUBS 0.013331f
C499 B.n136 VSUBS 0.013331f
C500 B.n137 VSUBS 0.013331f
C501 B.n138 VSUBS 0.013331f
C502 B.n139 VSUBS 0.013331f
C503 B.n140 VSUBS 0.013331f
C504 B.n141 VSUBS 0.013331f
C505 B.n142 VSUBS 0.013331f
C506 B.n143 VSUBS 0.013331f
C507 B.n144 VSUBS 0.013331f
C508 B.n145 VSUBS 0.013331f
C509 B.n146 VSUBS 0.013331f
C510 B.n147 VSUBS 0.030624f
C511 B.n148 VSUBS 0.013331f
C512 B.n149 VSUBS 0.013331f
C513 B.n150 VSUBS 0.013331f
C514 B.n151 VSUBS 0.013331f
C515 B.n152 VSUBS 0.013331f
C516 B.n153 VSUBS 0.013331f
C517 B.n154 VSUBS 0.009214f
C518 B.n155 VSUBS 0.013331f
C519 B.n156 VSUBS 0.013331f
C520 B.n157 VSUBS 0.013331f
C521 B.n158 VSUBS 0.013331f
C522 B.n159 VSUBS 0.013331f
C523 B.t8 VSUBS 0.12556f
C524 B.t7 VSUBS 0.165768f
C525 B.t6 VSUBS 0.984419f
C526 B.n160 VSUBS 0.168375f
C527 B.n161 VSUBS 0.131007f
C528 B.n162 VSUBS 0.013331f
C529 B.n163 VSUBS 0.013331f
C530 B.n164 VSUBS 0.013331f
C531 B.n165 VSUBS 0.013331f
C532 B.n166 VSUBS 0.013331f
C533 B.n167 VSUBS 0.013331f
C534 B.n168 VSUBS 0.030624f
C535 B.n169 VSUBS 0.013331f
C536 B.n170 VSUBS 0.013331f
C537 B.n171 VSUBS 0.013331f
C538 B.n172 VSUBS 0.013331f
C539 B.n173 VSUBS 0.013331f
C540 B.n174 VSUBS 0.013331f
C541 B.n175 VSUBS 0.013331f
C542 B.n176 VSUBS 0.013331f
C543 B.n177 VSUBS 0.013331f
C544 B.n178 VSUBS 0.013331f
C545 B.n179 VSUBS 0.013331f
C546 B.n180 VSUBS 0.013331f
C547 B.n181 VSUBS 0.013331f
C548 B.n182 VSUBS 0.013331f
C549 B.n183 VSUBS 0.013331f
C550 B.n184 VSUBS 0.013331f
C551 B.n185 VSUBS 0.013331f
C552 B.n186 VSUBS 0.013331f
C553 B.n187 VSUBS 0.013331f
C554 B.n188 VSUBS 0.013331f
C555 B.n189 VSUBS 0.013331f
C556 B.n190 VSUBS 0.013331f
C557 B.n191 VSUBS 0.013331f
C558 B.n192 VSUBS 0.013331f
C559 B.n193 VSUBS 0.013331f
C560 B.n194 VSUBS 0.013331f
C561 B.n195 VSUBS 0.013331f
C562 B.n196 VSUBS 0.013331f
C563 B.n197 VSUBS 0.013331f
C564 B.n198 VSUBS 0.013331f
C565 B.n199 VSUBS 0.013331f
C566 B.n200 VSUBS 0.013331f
C567 B.n201 VSUBS 0.013331f
C568 B.n202 VSUBS 0.013331f
C569 B.n203 VSUBS 0.013331f
C570 B.n204 VSUBS 0.013331f
C571 B.n205 VSUBS 0.013331f
C572 B.n206 VSUBS 0.013331f
C573 B.n207 VSUBS 0.013331f
C574 B.n208 VSUBS 0.013331f
C575 B.n209 VSUBS 0.013331f
C576 B.n210 VSUBS 0.013331f
C577 B.n211 VSUBS 0.013331f
C578 B.n212 VSUBS 0.013331f
C579 B.n213 VSUBS 0.013331f
C580 B.n214 VSUBS 0.013331f
C581 B.n215 VSUBS 0.013331f
C582 B.n216 VSUBS 0.013331f
C583 B.n217 VSUBS 0.013331f
C584 B.n218 VSUBS 0.013331f
C585 B.n219 VSUBS 0.013331f
C586 B.n220 VSUBS 0.013331f
C587 B.n221 VSUBS 0.013331f
C588 B.n222 VSUBS 0.013331f
C589 B.n223 VSUBS 0.013331f
C590 B.n224 VSUBS 0.013331f
C591 B.n225 VSUBS 0.013331f
C592 B.n226 VSUBS 0.013331f
C593 B.n227 VSUBS 0.013331f
C594 B.n228 VSUBS 0.013331f
C595 B.n229 VSUBS 0.013331f
C596 B.n230 VSUBS 0.013331f
C597 B.n231 VSUBS 0.013331f
C598 B.n232 VSUBS 0.013331f
C599 B.n233 VSUBS 0.013331f
C600 B.n234 VSUBS 0.013331f
C601 B.n235 VSUBS 0.013331f
C602 B.n236 VSUBS 0.013331f
C603 B.n237 VSUBS 0.013331f
C604 B.n238 VSUBS 0.013331f
C605 B.n239 VSUBS 0.013331f
C606 B.n240 VSUBS 0.013331f
C607 B.n241 VSUBS 0.013331f
C608 B.n242 VSUBS 0.013331f
C609 B.n243 VSUBS 0.013331f
C610 B.n244 VSUBS 0.013331f
C611 B.n245 VSUBS 0.013331f
C612 B.n246 VSUBS 0.013331f
C613 B.n247 VSUBS 0.013331f
C614 B.n248 VSUBS 0.013331f
C615 B.n249 VSUBS 0.013331f
C616 B.n250 VSUBS 0.013331f
C617 B.n251 VSUBS 0.013331f
C618 B.n252 VSUBS 0.013331f
C619 B.n253 VSUBS 0.013331f
C620 B.n254 VSUBS 0.013331f
C621 B.n255 VSUBS 0.013331f
C622 B.n256 VSUBS 0.013331f
C623 B.n257 VSUBS 0.013331f
C624 B.n258 VSUBS 0.013331f
C625 B.n259 VSUBS 0.013331f
C626 B.n260 VSUBS 0.013331f
C627 B.n261 VSUBS 0.013331f
C628 B.n262 VSUBS 0.013331f
C629 B.n263 VSUBS 0.013331f
C630 B.n264 VSUBS 0.013331f
C631 B.n265 VSUBS 0.013331f
C632 B.n266 VSUBS 0.013331f
C633 B.n267 VSUBS 0.013331f
C634 B.n268 VSUBS 0.013331f
C635 B.n269 VSUBS 0.013331f
C636 B.n270 VSUBS 0.013331f
C637 B.n271 VSUBS 0.013331f
C638 B.n272 VSUBS 0.013331f
C639 B.n273 VSUBS 0.013331f
C640 B.n274 VSUBS 0.013331f
C641 B.n275 VSUBS 0.013331f
C642 B.n276 VSUBS 0.013331f
C643 B.n277 VSUBS 0.013331f
C644 B.n278 VSUBS 0.013331f
C645 B.n279 VSUBS 0.013331f
C646 B.n280 VSUBS 0.013331f
C647 B.n281 VSUBS 0.013331f
C648 B.n282 VSUBS 0.013331f
C649 B.n283 VSUBS 0.013331f
C650 B.n284 VSUBS 0.013331f
C651 B.n285 VSUBS 0.013331f
C652 B.n286 VSUBS 0.013331f
C653 B.n287 VSUBS 0.013331f
C654 B.n288 VSUBS 0.013331f
C655 B.n289 VSUBS 0.013331f
C656 B.n290 VSUBS 0.013331f
C657 B.n291 VSUBS 0.013331f
C658 B.n292 VSUBS 0.013331f
C659 B.n293 VSUBS 0.013331f
C660 B.n294 VSUBS 0.013331f
C661 B.n295 VSUBS 0.013331f
C662 B.n296 VSUBS 0.013331f
C663 B.n297 VSUBS 0.013331f
C664 B.n298 VSUBS 0.013331f
C665 B.n299 VSUBS 0.013331f
C666 B.n300 VSUBS 0.013331f
C667 B.n301 VSUBS 0.013331f
C668 B.n302 VSUBS 0.013331f
C669 B.n303 VSUBS 0.013331f
C670 B.n304 VSUBS 0.013331f
C671 B.n305 VSUBS 0.013331f
C672 B.n306 VSUBS 0.013331f
C673 B.n307 VSUBS 0.013331f
C674 B.n308 VSUBS 0.013331f
C675 B.n309 VSUBS 0.013331f
C676 B.n310 VSUBS 0.013331f
C677 B.n311 VSUBS 0.013331f
C678 B.n312 VSUBS 0.013331f
C679 B.n313 VSUBS 0.013331f
C680 B.n314 VSUBS 0.013331f
C681 B.n315 VSUBS 0.013331f
C682 B.n316 VSUBS 0.013331f
C683 B.n317 VSUBS 0.013331f
C684 B.n318 VSUBS 0.013331f
C685 B.n319 VSUBS 0.013331f
C686 B.n320 VSUBS 0.013331f
C687 B.n321 VSUBS 0.013331f
C688 B.n322 VSUBS 0.013331f
C689 B.n323 VSUBS 0.013331f
C690 B.n324 VSUBS 0.013331f
C691 B.n325 VSUBS 0.028583f
C692 B.n326 VSUBS 0.028583f
C693 B.n327 VSUBS 0.030624f
C694 B.n328 VSUBS 0.013331f
C695 B.n329 VSUBS 0.013331f
C696 B.n330 VSUBS 0.013331f
C697 B.n331 VSUBS 0.013331f
C698 B.n332 VSUBS 0.013331f
C699 B.n333 VSUBS 0.013331f
C700 B.n334 VSUBS 0.013331f
C701 B.n335 VSUBS 0.013331f
C702 B.n336 VSUBS 0.013331f
C703 B.n337 VSUBS 0.013331f
C704 B.n338 VSUBS 0.013331f
C705 B.n339 VSUBS 0.013331f
C706 B.n340 VSUBS 0.013331f
C707 B.n341 VSUBS 0.013331f
C708 B.n342 VSUBS 0.013331f
C709 B.n343 VSUBS 0.013331f
C710 B.n344 VSUBS 0.013331f
C711 B.n345 VSUBS 0.013331f
C712 B.n346 VSUBS 0.013331f
C713 B.n347 VSUBS 0.013331f
C714 B.n348 VSUBS 0.009214f
C715 B.n349 VSUBS 0.030887f
C716 B.n350 VSUBS 0.010783f
C717 B.n351 VSUBS 0.013331f
C718 B.n352 VSUBS 0.013331f
C719 B.n353 VSUBS 0.013331f
C720 B.n354 VSUBS 0.013331f
C721 B.n355 VSUBS 0.013331f
C722 B.n356 VSUBS 0.013331f
C723 B.n357 VSUBS 0.013331f
C724 B.n358 VSUBS 0.013331f
C725 B.n359 VSUBS 0.013331f
C726 B.n360 VSUBS 0.013331f
C727 B.n361 VSUBS 0.013331f
C728 B.t2 VSUBS 0.12556f
C729 B.t1 VSUBS 0.165768f
C730 B.t0 VSUBS 0.984419f
C731 B.n362 VSUBS 0.168375f
C732 B.n363 VSUBS 0.131007f
C733 B.n364 VSUBS 0.030887f
C734 B.n365 VSUBS 0.010783f
C735 B.n366 VSUBS 0.013331f
C736 B.n367 VSUBS 0.013331f
C737 B.n368 VSUBS 0.013331f
C738 B.n369 VSUBS 0.013331f
C739 B.n370 VSUBS 0.013331f
C740 B.n371 VSUBS 0.013331f
C741 B.n372 VSUBS 0.013331f
C742 B.n373 VSUBS 0.013331f
C743 B.n374 VSUBS 0.013331f
C744 B.n375 VSUBS 0.013331f
C745 B.n376 VSUBS 0.013331f
C746 B.n377 VSUBS 0.013331f
C747 B.n378 VSUBS 0.013331f
C748 B.n379 VSUBS 0.013331f
C749 B.n380 VSUBS 0.013331f
C750 B.n381 VSUBS 0.013331f
C751 B.n382 VSUBS 0.013331f
C752 B.n383 VSUBS 0.013331f
C753 B.n384 VSUBS 0.013331f
C754 B.n385 VSUBS 0.013331f
C755 B.n386 VSUBS 0.013331f
C756 B.n387 VSUBS 0.013331f
C757 B.n388 VSUBS 0.028916f
C758 B.n389 VSUBS 0.03029f
C759 B.n390 VSUBS 0.028583f
C760 B.n391 VSUBS 0.013331f
C761 B.n392 VSUBS 0.013331f
C762 B.n393 VSUBS 0.013331f
C763 B.n394 VSUBS 0.013331f
C764 B.n395 VSUBS 0.013331f
C765 B.n396 VSUBS 0.013331f
C766 B.n397 VSUBS 0.013331f
C767 B.n398 VSUBS 0.013331f
C768 B.n399 VSUBS 0.013331f
C769 B.n400 VSUBS 0.013331f
C770 B.n401 VSUBS 0.013331f
C771 B.n402 VSUBS 0.013331f
C772 B.n403 VSUBS 0.013331f
C773 B.n404 VSUBS 0.013331f
C774 B.n405 VSUBS 0.013331f
C775 B.n406 VSUBS 0.013331f
C776 B.n407 VSUBS 0.013331f
C777 B.n408 VSUBS 0.013331f
C778 B.n409 VSUBS 0.013331f
C779 B.n410 VSUBS 0.013331f
C780 B.n411 VSUBS 0.013331f
C781 B.n412 VSUBS 0.013331f
C782 B.n413 VSUBS 0.013331f
C783 B.n414 VSUBS 0.013331f
C784 B.n415 VSUBS 0.013331f
C785 B.n416 VSUBS 0.013331f
C786 B.n417 VSUBS 0.013331f
C787 B.n418 VSUBS 0.013331f
C788 B.n419 VSUBS 0.013331f
C789 B.n420 VSUBS 0.013331f
C790 B.n421 VSUBS 0.013331f
C791 B.n422 VSUBS 0.013331f
C792 B.n423 VSUBS 0.013331f
C793 B.n424 VSUBS 0.013331f
C794 B.n425 VSUBS 0.013331f
C795 B.n426 VSUBS 0.013331f
C796 B.n427 VSUBS 0.013331f
C797 B.n428 VSUBS 0.013331f
C798 B.n429 VSUBS 0.013331f
C799 B.n430 VSUBS 0.013331f
C800 B.n431 VSUBS 0.013331f
C801 B.n432 VSUBS 0.013331f
C802 B.n433 VSUBS 0.013331f
C803 B.n434 VSUBS 0.013331f
C804 B.n435 VSUBS 0.013331f
C805 B.n436 VSUBS 0.013331f
C806 B.n437 VSUBS 0.013331f
C807 B.n438 VSUBS 0.013331f
C808 B.n439 VSUBS 0.013331f
C809 B.n440 VSUBS 0.013331f
C810 B.n441 VSUBS 0.013331f
C811 B.n442 VSUBS 0.013331f
C812 B.n443 VSUBS 0.013331f
C813 B.n444 VSUBS 0.013331f
C814 B.n445 VSUBS 0.013331f
C815 B.n446 VSUBS 0.013331f
C816 B.n447 VSUBS 0.013331f
C817 B.n448 VSUBS 0.013331f
C818 B.n449 VSUBS 0.013331f
C819 B.n450 VSUBS 0.013331f
C820 B.n451 VSUBS 0.013331f
C821 B.n452 VSUBS 0.013331f
C822 B.n453 VSUBS 0.013331f
C823 B.n454 VSUBS 0.013331f
C824 B.n455 VSUBS 0.013331f
C825 B.n456 VSUBS 0.013331f
C826 B.n457 VSUBS 0.013331f
C827 B.n458 VSUBS 0.013331f
C828 B.n459 VSUBS 0.013331f
C829 B.n460 VSUBS 0.013331f
C830 B.n461 VSUBS 0.013331f
C831 B.n462 VSUBS 0.013331f
C832 B.n463 VSUBS 0.013331f
C833 B.n464 VSUBS 0.013331f
C834 B.n465 VSUBS 0.013331f
C835 B.n466 VSUBS 0.013331f
C836 B.n467 VSUBS 0.013331f
C837 B.n468 VSUBS 0.013331f
C838 B.n469 VSUBS 0.013331f
C839 B.n470 VSUBS 0.013331f
C840 B.n471 VSUBS 0.013331f
C841 B.n472 VSUBS 0.013331f
C842 B.n473 VSUBS 0.013331f
C843 B.n474 VSUBS 0.013331f
C844 B.n475 VSUBS 0.013331f
C845 B.n476 VSUBS 0.013331f
C846 B.n477 VSUBS 0.013331f
C847 B.n478 VSUBS 0.013331f
C848 B.n479 VSUBS 0.013331f
C849 B.n480 VSUBS 0.013331f
C850 B.n481 VSUBS 0.013331f
C851 B.n482 VSUBS 0.013331f
C852 B.n483 VSUBS 0.013331f
C853 B.n484 VSUBS 0.013331f
C854 B.n485 VSUBS 0.013331f
C855 B.n486 VSUBS 0.013331f
C856 B.n487 VSUBS 0.013331f
C857 B.n488 VSUBS 0.013331f
C858 B.n489 VSUBS 0.013331f
C859 B.n490 VSUBS 0.013331f
C860 B.n491 VSUBS 0.013331f
C861 B.n492 VSUBS 0.013331f
C862 B.n493 VSUBS 0.013331f
C863 B.n494 VSUBS 0.013331f
C864 B.n495 VSUBS 0.013331f
C865 B.n496 VSUBS 0.013331f
C866 B.n497 VSUBS 0.013331f
C867 B.n498 VSUBS 0.013331f
C868 B.n499 VSUBS 0.013331f
C869 B.n500 VSUBS 0.013331f
C870 B.n501 VSUBS 0.013331f
C871 B.n502 VSUBS 0.013331f
C872 B.n503 VSUBS 0.013331f
C873 B.n504 VSUBS 0.013331f
C874 B.n505 VSUBS 0.013331f
C875 B.n506 VSUBS 0.013331f
C876 B.n507 VSUBS 0.013331f
C877 B.n508 VSUBS 0.013331f
C878 B.n509 VSUBS 0.013331f
C879 B.n510 VSUBS 0.013331f
C880 B.n511 VSUBS 0.013331f
C881 B.n512 VSUBS 0.013331f
C882 B.n513 VSUBS 0.013331f
C883 B.n514 VSUBS 0.013331f
C884 B.n515 VSUBS 0.013331f
C885 B.n516 VSUBS 0.013331f
C886 B.n517 VSUBS 0.013331f
C887 B.n518 VSUBS 0.013331f
C888 B.n519 VSUBS 0.013331f
C889 B.n520 VSUBS 0.013331f
C890 B.n521 VSUBS 0.013331f
C891 B.n522 VSUBS 0.013331f
C892 B.n523 VSUBS 0.013331f
C893 B.n524 VSUBS 0.013331f
C894 B.n525 VSUBS 0.013331f
C895 B.n526 VSUBS 0.013331f
C896 B.n527 VSUBS 0.013331f
C897 B.n528 VSUBS 0.013331f
C898 B.n529 VSUBS 0.013331f
C899 B.n530 VSUBS 0.013331f
C900 B.n531 VSUBS 0.013331f
C901 B.n532 VSUBS 0.013331f
C902 B.n533 VSUBS 0.013331f
C903 B.n534 VSUBS 0.013331f
C904 B.n535 VSUBS 0.013331f
C905 B.n536 VSUBS 0.013331f
C906 B.n537 VSUBS 0.013331f
C907 B.n538 VSUBS 0.013331f
C908 B.n539 VSUBS 0.013331f
C909 B.n540 VSUBS 0.013331f
C910 B.n541 VSUBS 0.013331f
C911 B.n542 VSUBS 0.013331f
C912 B.n543 VSUBS 0.013331f
C913 B.n544 VSUBS 0.013331f
C914 B.n545 VSUBS 0.013331f
C915 B.n546 VSUBS 0.013331f
C916 B.n547 VSUBS 0.013331f
C917 B.n548 VSUBS 0.013331f
C918 B.n549 VSUBS 0.013331f
C919 B.n550 VSUBS 0.013331f
C920 B.n551 VSUBS 0.013331f
C921 B.n552 VSUBS 0.013331f
C922 B.n553 VSUBS 0.013331f
C923 B.n554 VSUBS 0.013331f
C924 B.n555 VSUBS 0.013331f
C925 B.n556 VSUBS 0.013331f
C926 B.n557 VSUBS 0.013331f
C927 B.n558 VSUBS 0.013331f
C928 B.n559 VSUBS 0.013331f
C929 B.n560 VSUBS 0.013331f
C930 B.n561 VSUBS 0.013331f
C931 B.n562 VSUBS 0.013331f
C932 B.n563 VSUBS 0.013331f
C933 B.n564 VSUBS 0.013331f
C934 B.n565 VSUBS 0.013331f
C935 B.n566 VSUBS 0.013331f
C936 B.n567 VSUBS 0.013331f
C937 B.n568 VSUBS 0.013331f
C938 B.n569 VSUBS 0.013331f
C939 B.n570 VSUBS 0.013331f
C940 B.n571 VSUBS 0.013331f
C941 B.n572 VSUBS 0.013331f
C942 B.n573 VSUBS 0.013331f
C943 B.n574 VSUBS 0.013331f
C944 B.n575 VSUBS 0.013331f
C945 B.n576 VSUBS 0.013331f
C946 B.n577 VSUBS 0.013331f
C947 B.n578 VSUBS 0.013331f
C948 B.n579 VSUBS 0.013331f
C949 B.n580 VSUBS 0.013331f
C950 B.n581 VSUBS 0.013331f
C951 B.n582 VSUBS 0.013331f
C952 B.n583 VSUBS 0.013331f
C953 B.n584 VSUBS 0.013331f
C954 B.n585 VSUBS 0.013331f
C955 B.n586 VSUBS 0.013331f
C956 B.n587 VSUBS 0.013331f
C957 B.n588 VSUBS 0.013331f
C958 B.n589 VSUBS 0.013331f
C959 B.n590 VSUBS 0.013331f
C960 B.n591 VSUBS 0.013331f
C961 B.n592 VSUBS 0.013331f
C962 B.n593 VSUBS 0.013331f
C963 B.n594 VSUBS 0.013331f
C964 B.n595 VSUBS 0.013331f
C965 B.n596 VSUBS 0.013331f
C966 B.n597 VSUBS 0.013331f
C967 B.n598 VSUBS 0.013331f
C968 B.n599 VSUBS 0.013331f
C969 B.n600 VSUBS 0.013331f
C970 B.n601 VSUBS 0.013331f
C971 B.n602 VSUBS 0.013331f
C972 B.n603 VSUBS 0.013331f
C973 B.n604 VSUBS 0.013331f
C974 B.n605 VSUBS 0.013331f
C975 B.n606 VSUBS 0.013331f
C976 B.n607 VSUBS 0.013331f
C977 B.n608 VSUBS 0.013331f
C978 B.n609 VSUBS 0.013331f
C979 B.n610 VSUBS 0.013331f
C980 B.n611 VSUBS 0.013331f
C981 B.n612 VSUBS 0.013331f
C982 B.n613 VSUBS 0.013331f
C983 B.n614 VSUBS 0.013331f
C984 B.n615 VSUBS 0.013331f
C985 B.n616 VSUBS 0.013331f
C986 B.n617 VSUBS 0.013331f
C987 B.n618 VSUBS 0.013331f
C988 B.n619 VSUBS 0.013331f
C989 B.n620 VSUBS 0.013331f
C990 B.n621 VSUBS 0.013331f
C991 B.n622 VSUBS 0.013331f
C992 B.n623 VSUBS 0.013331f
C993 B.n624 VSUBS 0.013331f
C994 B.n625 VSUBS 0.013331f
C995 B.n626 VSUBS 0.013331f
C996 B.n627 VSUBS 0.013331f
C997 B.n628 VSUBS 0.013331f
C998 B.n629 VSUBS 0.013331f
C999 B.n630 VSUBS 0.013331f
C1000 B.n631 VSUBS 0.028583f
C1001 B.n632 VSUBS 0.030624f
C1002 B.n633 VSUBS 0.030624f
C1003 B.n634 VSUBS 0.013331f
C1004 B.n635 VSUBS 0.013331f
C1005 B.n636 VSUBS 0.013331f
C1006 B.n637 VSUBS 0.013331f
C1007 B.n638 VSUBS 0.013331f
C1008 B.n639 VSUBS 0.013331f
C1009 B.n640 VSUBS 0.013331f
C1010 B.n641 VSUBS 0.013331f
C1011 B.n642 VSUBS 0.013331f
C1012 B.n643 VSUBS 0.013331f
C1013 B.n644 VSUBS 0.013331f
C1014 B.n645 VSUBS 0.013331f
C1015 B.n646 VSUBS 0.013331f
C1016 B.n647 VSUBS 0.013331f
C1017 B.n648 VSUBS 0.013331f
C1018 B.n649 VSUBS 0.013331f
C1019 B.n650 VSUBS 0.013331f
C1020 B.n651 VSUBS 0.013331f
C1021 B.n652 VSUBS 0.013331f
C1022 B.n653 VSUBS 0.009214f
C1023 B.n654 VSUBS 0.013331f
C1024 B.n655 VSUBS 0.013331f
C1025 B.n656 VSUBS 0.010783f
C1026 B.n657 VSUBS 0.013331f
C1027 B.n658 VSUBS 0.013331f
C1028 B.n659 VSUBS 0.013331f
C1029 B.n660 VSUBS 0.013331f
C1030 B.n661 VSUBS 0.013331f
C1031 B.n662 VSUBS 0.013331f
C1032 B.n663 VSUBS 0.013331f
C1033 B.n664 VSUBS 0.013331f
C1034 B.n665 VSUBS 0.013331f
C1035 B.n666 VSUBS 0.013331f
C1036 B.n667 VSUBS 0.013331f
C1037 B.n668 VSUBS 0.010783f
C1038 B.n669 VSUBS 0.030887f
C1039 B.n670 VSUBS 0.009214f
C1040 B.n671 VSUBS 0.013331f
C1041 B.n672 VSUBS 0.013331f
C1042 B.n673 VSUBS 0.013331f
C1043 B.n674 VSUBS 0.013331f
C1044 B.n675 VSUBS 0.013331f
C1045 B.n676 VSUBS 0.013331f
C1046 B.n677 VSUBS 0.013331f
C1047 B.n678 VSUBS 0.013331f
C1048 B.n679 VSUBS 0.013331f
C1049 B.n680 VSUBS 0.013331f
C1050 B.n681 VSUBS 0.013331f
C1051 B.n682 VSUBS 0.013331f
C1052 B.n683 VSUBS 0.013331f
C1053 B.n684 VSUBS 0.013331f
C1054 B.n685 VSUBS 0.013331f
C1055 B.n686 VSUBS 0.013331f
C1056 B.n687 VSUBS 0.013331f
C1057 B.n688 VSUBS 0.013331f
C1058 B.n689 VSUBS 0.013331f
C1059 B.n690 VSUBS 0.013331f
C1060 B.n691 VSUBS 0.030624f
C1061 B.n692 VSUBS 0.028583f
C1062 B.n693 VSUBS 0.028583f
C1063 B.n694 VSUBS 0.013331f
C1064 B.n695 VSUBS 0.013331f
C1065 B.n696 VSUBS 0.013331f
C1066 B.n697 VSUBS 0.013331f
C1067 B.n698 VSUBS 0.013331f
C1068 B.n699 VSUBS 0.013331f
C1069 B.n700 VSUBS 0.013331f
C1070 B.n701 VSUBS 0.013331f
C1071 B.n702 VSUBS 0.013331f
C1072 B.n703 VSUBS 0.013331f
C1073 B.n704 VSUBS 0.013331f
C1074 B.n705 VSUBS 0.013331f
C1075 B.n706 VSUBS 0.013331f
C1076 B.n707 VSUBS 0.013331f
C1077 B.n708 VSUBS 0.013331f
C1078 B.n709 VSUBS 0.013331f
C1079 B.n710 VSUBS 0.013331f
C1080 B.n711 VSUBS 0.013331f
C1081 B.n712 VSUBS 0.013331f
C1082 B.n713 VSUBS 0.013331f
C1083 B.n714 VSUBS 0.013331f
C1084 B.n715 VSUBS 0.013331f
C1085 B.n716 VSUBS 0.013331f
C1086 B.n717 VSUBS 0.013331f
C1087 B.n718 VSUBS 0.013331f
C1088 B.n719 VSUBS 0.013331f
C1089 B.n720 VSUBS 0.013331f
C1090 B.n721 VSUBS 0.013331f
C1091 B.n722 VSUBS 0.013331f
C1092 B.n723 VSUBS 0.013331f
C1093 B.n724 VSUBS 0.013331f
C1094 B.n725 VSUBS 0.013331f
C1095 B.n726 VSUBS 0.013331f
C1096 B.n727 VSUBS 0.013331f
C1097 B.n728 VSUBS 0.013331f
C1098 B.n729 VSUBS 0.013331f
C1099 B.n730 VSUBS 0.013331f
C1100 B.n731 VSUBS 0.013331f
C1101 B.n732 VSUBS 0.013331f
C1102 B.n733 VSUBS 0.013331f
C1103 B.n734 VSUBS 0.013331f
C1104 B.n735 VSUBS 0.013331f
C1105 B.n736 VSUBS 0.013331f
C1106 B.n737 VSUBS 0.013331f
C1107 B.n738 VSUBS 0.013331f
C1108 B.n739 VSUBS 0.013331f
C1109 B.n740 VSUBS 0.013331f
C1110 B.n741 VSUBS 0.013331f
C1111 B.n742 VSUBS 0.013331f
C1112 B.n743 VSUBS 0.013331f
C1113 B.n744 VSUBS 0.013331f
C1114 B.n745 VSUBS 0.013331f
C1115 B.n746 VSUBS 0.013331f
C1116 B.n747 VSUBS 0.013331f
C1117 B.n748 VSUBS 0.013331f
C1118 B.n749 VSUBS 0.013331f
C1119 B.n750 VSUBS 0.013331f
C1120 B.n751 VSUBS 0.013331f
C1121 B.n752 VSUBS 0.013331f
C1122 B.n753 VSUBS 0.013331f
C1123 B.n754 VSUBS 0.013331f
C1124 B.n755 VSUBS 0.013331f
C1125 B.n756 VSUBS 0.013331f
C1126 B.n757 VSUBS 0.013331f
C1127 B.n758 VSUBS 0.013331f
C1128 B.n759 VSUBS 0.013331f
C1129 B.n760 VSUBS 0.013331f
C1130 B.n761 VSUBS 0.013331f
C1131 B.n762 VSUBS 0.013331f
C1132 B.n763 VSUBS 0.013331f
C1133 B.n764 VSUBS 0.013331f
C1134 B.n765 VSUBS 0.013331f
C1135 B.n766 VSUBS 0.013331f
C1136 B.n767 VSUBS 0.013331f
C1137 B.n768 VSUBS 0.013331f
C1138 B.n769 VSUBS 0.013331f
C1139 B.n770 VSUBS 0.013331f
C1140 B.n771 VSUBS 0.013331f
C1141 B.n772 VSUBS 0.013331f
C1142 B.n773 VSUBS 0.013331f
C1143 B.n774 VSUBS 0.013331f
C1144 B.n775 VSUBS 0.013331f
C1145 B.n776 VSUBS 0.013331f
C1146 B.n777 VSUBS 0.013331f
C1147 B.n778 VSUBS 0.013331f
C1148 B.n779 VSUBS 0.013331f
C1149 B.n780 VSUBS 0.013331f
C1150 B.n781 VSUBS 0.013331f
C1151 B.n782 VSUBS 0.013331f
C1152 B.n783 VSUBS 0.013331f
C1153 B.n784 VSUBS 0.013331f
C1154 B.n785 VSUBS 0.013331f
C1155 B.n786 VSUBS 0.013331f
C1156 B.n787 VSUBS 0.013331f
C1157 B.n788 VSUBS 0.013331f
C1158 B.n789 VSUBS 0.013331f
C1159 B.n790 VSUBS 0.013331f
C1160 B.n791 VSUBS 0.013331f
C1161 B.n792 VSUBS 0.013331f
C1162 B.n793 VSUBS 0.013331f
C1163 B.n794 VSUBS 0.013331f
C1164 B.n795 VSUBS 0.013331f
C1165 B.n796 VSUBS 0.013331f
C1166 B.n797 VSUBS 0.013331f
C1167 B.n798 VSUBS 0.013331f
C1168 B.n799 VSUBS 0.013331f
C1169 B.n800 VSUBS 0.013331f
C1170 B.n801 VSUBS 0.013331f
C1171 B.n802 VSUBS 0.013331f
C1172 B.n803 VSUBS 0.013331f
C1173 B.n804 VSUBS 0.013331f
C1174 B.n805 VSUBS 0.013331f
C1175 B.n806 VSUBS 0.013331f
C1176 B.n807 VSUBS 0.013331f
C1177 B.n808 VSUBS 0.013331f
C1178 B.n809 VSUBS 0.013331f
C1179 B.n810 VSUBS 0.013331f
C1180 B.n811 VSUBS 0.017397f
C1181 B.n812 VSUBS 0.018532f
C1182 B.n813 VSUBS 0.036852f
.ends

