* NGSPICE file created from diff_pair_sample_1755.ext - technology: sky130A

.subckt diff_pair_sample_1755 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.871 pd=17.73 as=6.786 ps=35.58 w=17.4 l=1.94
X1 VTAIL.t4 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=2.871 ps=17.73 w=17.4 l=1.94
X2 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.871 pd=17.73 as=6.786 ps=35.58 w=17.4 l=1.94
X3 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=2.871 ps=17.73 w=17.4 l=1.94
X4 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=2.871 ps=17.73 w=17.4 l=1.94
X5 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=0 ps=0 w=17.4 l=1.94
X6 VDD1.t0 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.871 pd=17.73 as=6.786 ps=35.58 w=17.4 l=1.94
X7 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=0 ps=0 w=17.4 l=1.94
X8 VDD2.t1 VN.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.871 pd=17.73 as=6.786 ps=35.58 w=17.4 l=1.94
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=0 ps=0 w=17.4 l=1.94
X10 VTAIL.t5 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=2.871 ps=17.73 w=17.4 l=1.94
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.786 pd=35.58 as=0 ps=0 w=17.4 l=1.94
R0 VN.n0 VN.t1 251.471
R1 VN.n1 VN.t2 251.471
R2 VN.n0 VN.t0 250.948
R3 VN.n1 VN.t3 250.948
R4 VN VN.n1 56.0682
R5 VN VN.n0 7.48867
R6 VTAIL.n766 VTAIL.n765 289.615
R7 VTAIL.n94 VTAIL.n93 289.615
R8 VTAIL.n190 VTAIL.n189 289.615
R9 VTAIL.n286 VTAIL.n285 289.615
R10 VTAIL.n670 VTAIL.n669 289.615
R11 VTAIL.n574 VTAIL.n573 289.615
R12 VTAIL.n478 VTAIL.n477 289.615
R13 VTAIL.n382 VTAIL.n381 289.615
R14 VTAIL.n702 VTAIL.n701 185
R15 VTAIL.n707 VTAIL.n706 185
R16 VTAIL.n709 VTAIL.n708 185
R17 VTAIL.n698 VTAIL.n697 185
R18 VTAIL.n715 VTAIL.n714 185
R19 VTAIL.n717 VTAIL.n716 185
R20 VTAIL.n694 VTAIL.n693 185
R21 VTAIL.n724 VTAIL.n723 185
R22 VTAIL.n725 VTAIL.n692 185
R23 VTAIL.n727 VTAIL.n726 185
R24 VTAIL.n690 VTAIL.n689 185
R25 VTAIL.n733 VTAIL.n732 185
R26 VTAIL.n735 VTAIL.n734 185
R27 VTAIL.n686 VTAIL.n685 185
R28 VTAIL.n741 VTAIL.n740 185
R29 VTAIL.n743 VTAIL.n742 185
R30 VTAIL.n682 VTAIL.n681 185
R31 VTAIL.n749 VTAIL.n748 185
R32 VTAIL.n751 VTAIL.n750 185
R33 VTAIL.n678 VTAIL.n677 185
R34 VTAIL.n757 VTAIL.n756 185
R35 VTAIL.n759 VTAIL.n758 185
R36 VTAIL.n674 VTAIL.n673 185
R37 VTAIL.n765 VTAIL.n764 185
R38 VTAIL.n30 VTAIL.n29 185
R39 VTAIL.n35 VTAIL.n34 185
R40 VTAIL.n37 VTAIL.n36 185
R41 VTAIL.n26 VTAIL.n25 185
R42 VTAIL.n43 VTAIL.n42 185
R43 VTAIL.n45 VTAIL.n44 185
R44 VTAIL.n22 VTAIL.n21 185
R45 VTAIL.n52 VTAIL.n51 185
R46 VTAIL.n53 VTAIL.n20 185
R47 VTAIL.n55 VTAIL.n54 185
R48 VTAIL.n18 VTAIL.n17 185
R49 VTAIL.n61 VTAIL.n60 185
R50 VTAIL.n63 VTAIL.n62 185
R51 VTAIL.n14 VTAIL.n13 185
R52 VTAIL.n69 VTAIL.n68 185
R53 VTAIL.n71 VTAIL.n70 185
R54 VTAIL.n10 VTAIL.n9 185
R55 VTAIL.n77 VTAIL.n76 185
R56 VTAIL.n79 VTAIL.n78 185
R57 VTAIL.n6 VTAIL.n5 185
R58 VTAIL.n85 VTAIL.n84 185
R59 VTAIL.n87 VTAIL.n86 185
R60 VTAIL.n2 VTAIL.n1 185
R61 VTAIL.n93 VTAIL.n92 185
R62 VTAIL.n126 VTAIL.n125 185
R63 VTAIL.n131 VTAIL.n130 185
R64 VTAIL.n133 VTAIL.n132 185
R65 VTAIL.n122 VTAIL.n121 185
R66 VTAIL.n139 VTAIL.n138 185
R67 VTAIL.n141 VTAIL.n140 185
R68 VTAIL.n118 VTAIL.n117 185
R69 VTAIL.n148 VTAIL.n147 185
R70 VTAIL.n149 VTAIL.n116 185
R71 VTAIL.n151 VTAIL.n150 185
R72 VTAIL.n114 VTAIL.n113 185
R73 VTAIL.n157 VTAIL.n156 185
R74 VTAIL.n159 VTAIL.n158 185
R75 VTAIL.n110 VTAIL.n109 185
R76 VTAIL.n165 VTAIL.n164 185
R77 VTAIL.n167 VTAIL.n166 185
R78 VTAIL.n106 VTAIL.n105 185
R79 VTAIL.n173 VTAIL.n172 185
R80 VTAIL.n175 VTAIL.n174 185
R81 VTAIL.n102 VTAIL.n101 185
R82 VTAIL.n181 VTAIL.n180 185
R83 VTAIL.n183 VTAIL.n182 185
R84 VTAIL.n98 VTAIL.n97 185
R85 VTAIL.n189 VTAIL.n188 185
R86 VTAIL.n222 VTAIL.n221 185
R87 VTAIL.n227 VTAIL.n226 185
R88 VTAIL.n229 VTAIL.n228 185
R89 VTAIL.n218 VTAIL.n217 185
R90 VTAIL.n235 VTAIL.n234 185
R91 VTAIL.n237 VTAIL.n236 185
R92 VTAIL.n214 VTAIL.n213 185
R93 VTAIL.n244 VTAIL.n243 185
R94 VTAIL.n245 VTAIL.n212 185
R95 VTAIL.n247 VTAIL.n246 185
R96 VTAIL.n210 VTAIL.n209 185
R97 VTAIL.n253 VTAIL.n252 185
R98 VTAIL.n255 VTAIL.n254 185
R99 VTAIL.n206 VTAIL.n205 185
R100 VTAIL.n261 VTAIL.n260 185
R101 VTAIL.n263 VTAIL.n262 185
R102 VTAIL.n202 VTAIL.n201 185
R103 VTAIL.n269 VTAIL.n268 185
R104 VTAIL.n271 VTAIL.n270 185
R105 VTAIL.n198 VTAIL.n197 185
R106 VTAIL.n277 VTAIL.n276 185
R107 VTAIL.n279 VTAIL.n278 185
R108 VTAIL.n194 VTAIL.n193 185
R109 VTAIL.n285 VTAIL.n284 185
R110 VTAIL.n669 VTAIL.n668 185
R111 VTAIL.n578 VTAIL.n577 185
R112 VTAIL.n663 VTAIL.n662 185
R113 VTAIL.n661 VTAIL.n660 185
R114 VTAIL.n582 VTAIL.n581 185
R115 VTAIL.n655 VTAIL.n654 185
R116 VTAIL.n653 VTAIL.n652 185
R117 VTAIL.n586 VTAIL.n585 185
R118 VTAIL.n647 VTAIL.n646 185
R119 VTAIL.n645 VTAIL.n644 185
R120 VTAIL.n590 VTAIL.n589 185
R121 VTAIL.n639 VTAIL.n638 185
R122 VTAIL.n637 VTAIL.n636 185
R123 VTAIL.n594 VTAIL.n593 185
R124 VTAIL.n631 VTAIL.n630 185
R125 VTAIL.n629 VTAIL.n596 185
R126 VTAIL.n628 VTAIL.n627 185
R127 VTAIL.n599 VTAIL.n597 185
R128 VTAIL.n622 VTAIL.n621 185
R129 VTAIL.n620 VTAIL.n619 185
R130 VTAIL.n603 VTAIL.n602 185
R131 VTAIL.n614 VTAIL.n613 185
R132 VTAIL.n612 VTAIL.n611 185
R133 VTAIL.n607 VTAIL.n606 185
R134 VTAIL.n573 VTAIL.n572 185
R135 VTAIL.n482 VTAIL.n481 185
R136 VTAIL.n567 VTAIL.n566 185
R137 VTAIL.n565 VTAIL.n564 185
R138 VTAIL.n486 VTAIL.n485 185
R139 VTAIL.n559 VTAIL.n558 185
R140 VTAIL.n557 VTAIL.n556 185
R141 VTAIL.n490 VTAIL.n489 185
R142 VTAIL.n551 VTAIL.n550 185
R143 VTAIL.n549 VTAIL.n548 185
R144 VTAIL.n494 VTAIL.n493 185
R145 VTAIL.n543 VTAIL.n542 185
R146 VTAIL.n541 VTAIL.n540 185
R147 VTAIL.n498 VTAIL.n497 185
R148 VTAIL.n535 VTAIL.n534 185
R149 VTAIL.n533 VTAIL.n500 185
R150 VTAIL.n532 VTAIL.n531 185
R151 VTAIL.n503 VTAIL.n501 185
R152 VTAIL.n526 VTAIL.n525 185
R153 VTAIL.n524 VTAIL.n523 185
R154 VTAIL.n507 VTAIL.n506 185
R155 VTAIL.n518 VTAIL.n517 185
R156 VTAIL.n516 VTAIL.n515 185
R157 VTAIL.n511 VTAIL.n510 185
R158 VTAIL.n477 VTAIL.n476 185
R159 VTAIL.n386 VTAIL.n385 185
R160 VTAIL.n471 VTAIL.n470 185
R161 VTAIL.n469 VTAIL.n468 185
R162 VTAIL.n390 VTAIL.n389 185
R163 VTAIL.n463 VTAIL.n462 185
R164 VTAIL.n461 VTAIL.n460 185
R165 VTAIL.n394 VTAIL.n393 185
R166 VTAIL.n455 VTAIL.n454 185
R167 VTAIL.n453 VTAIL.n452 185
R168 VTAIL.n398 VTAIL.n397 185
R169 VTAIL.n447 VTAIL.n446 185
R170 VTAIL.n445 VTAIL.n444 185
R171 VTAIL.n402 VTAIL.n401 185
R172 VTAIL.n439 VTAIL.n438 185
R173 VTAIL.n437 VTAIL.n404 185
R174 VTAIL.n436 VTAIL.n435 185
R175 VTAIL.n407 VTAIL.n405 185
R176 VTAIL.n430 VTAIL.n429 185
R177 VTAIL.n428 VTAIL.n427 185
R178 VTAIL.n411 VTAIL.n410 185
R179 VTAIL.n422 VTAIL.n421 185
R180 VTAIL.n420 VTAIL.n419 185
R181 VTAIL.n415 VTAIL.n414 185
R182 VTAIL.n381 VTAIL.n380 185
R183 VTAIL.n290 VTAIL.n289 185
R184 VTAIL.n375 VTAIL.n374 185
R185 VTAIL.n373 VTAIL.n372 185
R186 VTAIL.n294 VTAIL.n293 185
R187 VTAIL.n367 VTAIL.n366 185
R188 VTAIL.n365 VTAIL.n364 185
R189 VTAIL.n298 VTAIL.n297 185
R190 VTAIL.n359 VTAIL.n358 185
R191 VTAIL.n357 VTAIL.n356 185
R192 VTAIL.n302 VTAIL.n301 185
R193 VTAIL.n351 VTAIL.n350 185
R194 VTAIL.n349 VTAIL.n348 185
R195 VTAIL.n306 VTAIL.n305 185
R196 VTAIL.n343 VTAIL.n342 185
R197 VTAIL.n341 VTAIL.n308 185
R198 VTAIL.n340 VTAIL.n339 185
R199 VTAIL.n311 VTAIL.n309 185
R200 VTAIL.n334 VTAIL.n333 185
R201 VTAIL.n332 VTAIL.n331 185
R202 VTAIL.n315 VTAIL.n314 185
R203 VTAIL.n326 VTAIL.n325 185
R204 VTAIL.n324 VTAIL.n323 185
R205 VTAIL.n319 VTAIL.n318 185
R206 VTAIL.n703 VTAIL.t7 149.524
R207 VTAIL.n31 VTAIL.t4 149.524
R208 VTAIL.n127 VTAIL.t1 149.524
R209 VTAIL.n223 VTAIL.t0 149.524
R210 VTAIL.n608 VTAIL.t3 149.524
R211 VTAIL.n512 VTAIL.t2 149.524
R212 VTAIL.n416 VTAIL.t6 149.524
R213 VTAIL.n320 VTAIL.t5 149.524
R214 VTAIL.n707 VTAIL.n701 104.615
R215 VTAIL.n708 VTAIL.n707 104.615
R216 VTAIL.n708 VTAIL.n697 104.615
R217 VTAIL.n715 VTAIL.n697 104.615
R218 VTAIL.n716 VTAIL.n715 104.615
R219 VTAIL.n716 VTAIL.n693 104.615
R220 VTAIL.n724 VTAIL.n693 104.615
R221 VTAIL.n725 VTAIL.n724 104.615
R222 VTAIL.n726 VTAIL.n725 104.615
R223 VTAIL.n726 VTAIL.n689 104.615
R224 VTAIL.n733 VTAIL.n689 104.615
R225 VTAIL.n734 VTAIL.n733 104.615
R226 VTAIL.n734 VTAIL.n685 104.615
R227 VTAIL.n741 VTAIL.n685 104.615
R228 VTAIL.n742 VTAIL.n741 104.615
R229 VTAIL.n742 VTAIL.n681 104.615
R230 VTAIL.n749 VTAIL.n681 104.615
R231 VTAIL.n750 VTAIL.n749 104.615
R232 VTAIL.n750 VTAIL.n677 104.615
R233 VTAIL.n757 VTAIL.n677 104.615
R234 VTAIL.n758 VTAIL.n757 104.615
R235 VTAIL.n758 VTAIL.n673 104.615
R236 VTAIL.n765 VTAIL.n673 104.615
R237 VTAIL.n35 VTAIL.n29 104.615
R238 VTAIL.n36 VTAIL.n35 104.615
R239 VTAIL.n36 VTAIL.n25 104.615
R240 VTAIL.n43 VTAIL.n25 104.615
R241 VTAIL.n44 VTAIL.n43 104.615
R242 VTAIL.n44 VTAIL.n21 104.615
R243 VTAIL.n52 VTAIL.n21 104.615
R244 VTAIL.n53 VTAIL.n52 104.615
R245 VTAIL.n54 VTAIL.n53 104.615
R246 VTAIL.n54 VTAIL.n17 104.615
R247 VTAIL.n61 VTAIL.n17 104.615
R248 VTAIL.n62 VTAIL.n61 104.615
R249 VTAIL.n62 VTAIL.n13 104.615
R250 VTAIL.n69 VTAIL.n13 104.615
R251 VTAIL.n70 VTAIL.n69 104.615
R252 VTAIL.n70 VTAIL.n9 104.615
R253 VTAIL.n77 VTAIL.n9 104.615
R254 VTAIL.n78 VTAIL.n77 104.615
R255 VTAIL.n78 VTAIL.n5 104.615
R256 VTAIL.n85 VTAIL.n5 104.615
R257 VTAIL.n86 VTAIL.n85 104.615
R258 VTAIL.n86 VTAIL.n1 104.615
R259 VTAIL.n93 VTAIL.n1 104.615
R260 VTAIL.n131 VTAIL.n125 104.615
R261 VTAIL.n132 VTAIL.n131 104.615
R262 VTAIL.n132 VTAIL.n121 104.615
R263 VTAIL.n139 VTAIL.n121 104.615
R264 VTAIL.n140 VTAIL.n139 104.615
R265 VTAIL.n140 VTAIL.n117 104.615
R266 VTAIL.n148 VTAIL.n117 104.615
R267 VTAIL.n149 VTAIL.n148 104.615
R268 VTAIL.n150 VTAIL.n149 104.615
R269 VTAIL.n150 VTAIL.n113 104.615
R270 VTAIL.n157 VTAIL.n113 104.615
R271 VTAIL.n158 VTAIL.n157 104.615
R272 VTAIL.n158 VTAIL.n109 104.615
R273 VTAIL.n165 VTAIL.n109 104.615
R274 VTAIL.n166 VTAIL.n165 104.615
R275 VTAIL.n166 VTAIL.n105 104.615
R276 VTAIL.n173 VTAIL.n105 104.615
R277 VTAIL.n174 VTAIL.n173 104.615
R278 VTAIL.n174 VTAIL.n101 104.615
R279 VTAIL.n181 VTAIL.n101 104.615
R280 VTAIL.n182 VTAIL.n181 104.615
R281 VTAIL.n182 VTAIL.n97 104.615
R282 VTAIL.n189 VTAIL.n97 104.615
R283 VTAIL.n227 VTAIL.n221 104.615
R284 VTAIL.n228 VTAIL.n227 104.615
R285 VTAIL.n228 VTAIL.n217 104.615
R286 VTAIL.n235 VTAIL.n217 104.615
R287 VTAIL.n236 VTAIL.n235 104.615
R288 VTAIL.n236 VTAIL.n213 104.615
R289 VTAIL.n244 VTAIL.n213 104.615
R290 VTAIL.n245 VTAIL.n244 104.615
R291 VTAIL.n246 VTAIL.n245 104.615
R292 VTAIL.n246 VTAIL.n209 104.615
R293 VTAIL.n253 VTAIL.n209 104.615
R294 VTAIL.n254 VTAIL.n253 104.615
R295 VTAIL.n254 VTAIL.n205 104.615
R296 VTAIL.n261 VTAIL.n205 104.615
R297 VTAIL.n262 VTAIL.n261 104.615
R298 VTAIL.n262 VTAIL.n201 104.615
R299 VTAIL.n269 VTAIL.n201 104.615
R300 VTAIL.n270 VTAIL.n269 104.615
R301 VTAIL.n270 VTAIL.n197 104.615
R302 VTAIL.n277 VTAIL.n197 104.615
R303 VTAIL.n278 VTAIL.n277 104.615
R304 VTAIL.n278 VTAIL.n193 104.615
R305 VTAIL.n285 VTAIL.n193 104.615
R306 VTAIL.n669 VTAIL.n577 104.615
R307 VTAIL.n662 VTAIL.n577 104.615
R308 VTAIL.n662 VTAIL.n661 104.615
R309 VTAIL.n661 VTAIL.n581 104.615
R310 VTAIL.n654 VTAIL.n581 104.615
R311 VTAIL.n654 VTAIL.n653 104.615
R312 VTAIL.n653 VTAIL.n585 104.615
R313 VTAIL.n646 VTAIL.n585 104.615
R314 VTAIL.n646 VTAIL.n645 104.615
R315 VTAIL.n645 VTAIL.n589 104.615
R316 VTAIL.n638 VTAIL.n589 104.615
R317 VTAIL.n638 VTAIL.n637 104.615
R318 VTAIL.n637 VTAIL.n593 104.615
R319 VTAIL.n630 VTAIL.n593 104.615
R320 VTAIL.n630 VTAIL.n629 104.615
R321 VTAIL.n629 VTAIL.n628 104.615
R322 VTAIL.n628 VTAIL.n597 104.615
R323 VTAIL.n621 VTAIL.n597 104.615
R324 VTAIL.n621 VTAIL.n620 104.615
R325 VTAIL.n620 VTAIL.n602 104.615
R326 VTAIL.n613 VTAIL.n602 104.615
R327 VTAIL.n613 VTAIL.n612 104.615
R328 VTAIL.n612 VTAIL.n606 104.615
R329 VTAIL.n573 VTAIL.n481 104.615
R330 VTAIL.n566 VTAIL.n481 104.615
R331 VTAIL.n566 VTAIL.n565 104.615
R332 VTAIL.n565 VTAIL.n485 104.615
R333 VTAIL.n558 VTAIL.n485 104.615
R334 VTAIL.n558 VTAIL.n557 104.615
R335 VTAIL.n557 VTAIL.n489 104.615
R336 VTAIL.n550 VTAIL.n489 104.615
R337 VTAIL.n550 VTAIL.n549 104.615
R338 VTAIL.n549 VTAIL.n493 104.615
R339 VTAIL.n542 VTAIL.n493 104.615
R340 VTAIL.n542 VTAIL.n541 104.615
R341 VTAIL.n541 VTAIL.n497 104.615
R342 VTAIL.n534 VTAIL.n497 104.615
R343 VTAIL.n534 VTAIL.n533 104.615
R344 VTAIL.n533 VTAIL.n532 104.615
R345 VTAIL.n532 VTAIL.n501 104.615
R346 VTAIL.n525 VTAIL.n501 104.615
R347 VTAIL.n525 VTAIL.n524 104.615
R348 VTAIL.n524 VTAIL.n506 104.615
R349 VTAIL.n517 VTAIL.n506 104.615
R350 VTAIL.n517 VTAIL.n516 104.615
R351 VTAIL.n516 VTAIL.n510 104.615
R352 VTAIL.n477 VTAIL.n385 104.615
R353 VTAIL.n470 VTAIL.n385 104.615
R354 VTAIL.n470 VTAIL.n469 104.615
R355 VTAIL.n469 VTAIL.n389 104.615
R356 VTAIL.n462 VTAIL.n389 104.615
R357 VTAIL.n462 VTAIL.n461 104.615
R358 VTAIL.n461 VTAIL.n393 104.615
R359 VTAIL.n454 VTAIL.n393 104.615
R360 VTAIL.n454 VTAIL.n453 104.615
R361 VTAIL.n453 VTAIL.n397 104.615
R362 VTAIL.n446 VTAIL.n397 104.615
R363 VTAIL.n446 VTAIL.n445 104.615
R364 VTAIL.n445 VTAIL.n401 104.615
R365 VTAIL.n438 VTAIL.n401 104.615
R366 VTAIL.n438 VTAIL.n437 104.615
R367 VTAIL.n437 VTAIL.n436 104.615
R368 VTAIL.n436 VTAIL.n405 104.615
R369 VTAIL.n429 VTAIL.n405 104.615
R370 VTAIL.n429 VTAIL.n428 104.615
R371 VTAIL.n428 VTAIL.n410 104.615
R372 VTAIL.n421 VTAIL.n410 104.615
R373 VTAIL.n421 VTAIL.n420 104.615
R374 VTAIL.n420 VTAIL.n414 104.615
R375 VTAIL.n381 VTAIL.n289 104.615
R376 VTAIL.n374 VTAIL.n289 104.615
R377 VTAIL.n374 VTAIL.n373 104.615
R378 VTAIL.n373 VTAIL.n293 104.615
R379 VTAIL.n366 VTAIL.n293 104.615
R380 VTAIL.n366 VTAIL.n365 104.615
R381 VTAIL.n365 VTAIL.n297 104.615
R382 VTAIL.n358 VTAIL.n297 104.615
R383 VTAIL.n358 VTAIL.n357 104.615
R384 VTAIL.n357 VTAIL.n301 104.615
R385 VTAIL.n350 VTAIL.n301 104.615
R386 VTAIL.n350 VTAIL.n349 104.615
R387 VTAIL.n349 VTAIL.n305 104.615
R388 VTAIL.n342 VTAIL.n305 104.615
R389 VTAIL.n342 VTAIL.n341 104.615
R390 VTAIL.n341 VTAIL.n340 104.615
R391 VTAIL.n340 VTAIL.n309 104.615
R392 VTAIL.n333 VTAIL.n309 104.615
R393 VTAIL.n333 VTAIL.n332 104.615
R394 VTAIL.n332 VTAIL.n314 104.615
R395 VTAIL.n325 VTAIL.n314 104.615
R396 VTAIL.n325 VTAIL.n324 104.615
R397 VTAIL.n324 VTAIL.n318 104.615
R398 VTAIL.t7 VTAIL.n701 52.3082
R399 VTAIL.t4 VTAIL.n29 52.3082
R400 VTAIL.t1 VTAIL.n125 52.3082
R401 VTAIL.t0 VTAIL.n221 52.3082
R402 VTAIL.t3 VTAIL.n606 52.3082
R403 VTAIL.t2 VTAIL.n510 52.3082
R404 VTAIL.t6 VTAIL.n414 52.3082
R405 VTAIL.t5 VTAIL.n318 52.3082
R406 VTAIL.n767 VTAIL.n766 34.9005
R407 VTAIL.n95 VTAIL.n94 34.9005
R408 VTAIL.n191 VTAIL.n190 34.9005
R409 VTAIL.n287 VTAIL.n286 34.9005
R410 VTAIL.n671 VTAIL.n670 34.9005
R411 VTAIL.n575 VTAIL.n574 34.9005
R412 VTAIL.n479 VTAIL.n478 34.9005
R413 VTAIL.n383 VTAIL.n382 34.9005
R414 VTAIL.n767 VTAIL.n671 29.3238
R415 VTAIL.n383 VTAIL.n287 29.3238
R416 VTAIL.n727 VTAIL.n692 13.1884
R417 VTAIL.n55 VTAIL.n20 13.1884
R418 VTAIL.n151 VTAIL.n116 13.1884
R419 VTAIL.n247 VTAIL.n212 13.1884
R420 VTAIL.n631 VTAIL.n596 13.1884
R421 VTAIL.n535 VTAIL.n500 13.1884
R422 VTAIL.n439 VTAIL.n404 13.1884
R423 VTAIL.n343 VTAIL.n308 13.1884
R424 VTAIL.n723 VTAIL.n722 12.8005
R425 VTAIL.n728 VTAIL.n690 12.8005
R426 VTAIL.n51 VTAIL.n50 12.8005
R427 VTAIL.n56 VTAIL.n18 12.8005
R428 VTAIL.n147 VTAIL.n146 12.8005
R429 VTAIL.n152 VTAIL.n114 12.8005
R430 VTAIL.n243 VTAIL.n242 12.8005
R431 VTAIL.n248 VTAIL.n210 12.8005
R432 VTAIL.n632 VTAIL.n594 12.8005
R433 VTAIL.n627 VTAIL.n598 12.8005
R434 VTAIL.n536 VTAIL.n498 12.8005
R435 VTAIL.n531 VTAIL.n502 12.8005
R436 VTAIL.n440 VTAIL.n402 12.8005
R437 VTAIL.n435 VTAIL.n406 12.8005
R438 VTAIL.n344 VTAIL.n306 12.8005
R439 VTAIL.n339 VTAIL.n310 12.8005
R440 VTAIL.n721 VTAIL.n694 12.0247
R441 VTAIL.n732 VTAIL.n731 12.0247
R442 VTAIL.n49 VTAIL.n22 12.0247
R443 VTAIL.n60 VTAIL.n59 12.0247
R444 VTAIL.n145 VTAIL.n118 12.0247
R445 VTAIL.n156 VTAIL.n155 12.0247
R446 VTAIL.n241 VTAIL.n214 12.0247
R447 VTAIL.n252 VTAIL.n251 12.0247
R448 VTAIL.n636 VTAIL.n635 12.0247
R449 VTAIL.n626 VTAIL.n599 12.0247
R450 VTAIL.n540 VTAIL.n539 12.0247
R451 VTAIL.n530 VTAIL.n503 12.0247
R452 VTAIL.n444 VTAIL.n443 12.0247
R453 VTAIL.n434 VTAIL.n407 12.0247
R454 VTAIL.n348 VTAIL.n347 12.0247
R455 VTAIL.n338 VTAIL.n311 12.0247
R456 VTAIL.n718 VTAIL.n717 11.249
R457 VTAIL.n735 VTAIL.n688 11.249
R458 VTAIL.n764 VTAIL.n672 11.249
R459 VTAIL.n46 VTAIL.n45 11.249
R460 VTAIL.n63 VTAIL.n16 11.249
R461 VTAIL.n92 VTAIL.n0 11.249
R462 VTAIL.n142 VTAIL.n141 11.249
R463 VTAIL.n159 VTAIL.n112 11.249
R464 VTAIL.n188 VTAIL.n96 11.249
R465 VTAIL.n238 VTAIL.n237 11.249
R466 VTAIL.n255 VTAIL.n208 11.249
R467 VTAIL.n284 VTAIL.n192 11.249
R468 VTAIL.n668 VTAIL.n576 11.249
R469 VTAIL.n639 VTAIL.n592 11.249
R470 VTAIL.n623 VTAIL.n622 11.249
R471 VTAIL.n572 VTAIL.n480 11.249
R472 VTAIL.n543 VTAIL.n496 11.249
R473 VTAIL.n527 VTAIL.n526 11.249
R474 VTAIL.n476 VTAIL.n384 11.249
R475 VTAIL.n447 VTAIL.n400 11.249
R476 VTAIL.n431 VTAIL.n430 11.249
R477 VTAIL.n380 VTAIL.n288 11.249
R478 VTAIL.n351 VTAIL.n304 11.249
R479 VTAIL.n335 VTAIL.n334 11.249
R480 VTAIL.n714 VTAIL.n696 10.4732
R481 VTAIL.n736 VTAIL.n686 10.4732
R482 VTAIL.n763 VTAIL.n674 10.4732
R483 VTAIL.n42 VTAIL.n24 10.4732
R484 VTAIL.n64 VTAIL.n14 10.4732
R485 VTAIL.n91 VTAIL.n2 10.4732
R486 VTAIL.n138 VTAIL.n120 10.4732
R487 VTAIL.n160 VTAIL.n110 10.4732
R488 VTAIL.n187 VTAIL.n98 10.4732
R489 VTAIL.n234 VTAIL.n216 10.4732
R490 VTAIL.n256 VTAIL.n206 10.4732
R491 VTAIL.n283 VTAIL.n194 10.4732
R492 VTAIL.n667 VTAIL.n578 10.4732
R493 VTAIL.n640 VTAIL.n590 10.4732
R494 VTAIL.n619 VTAIL.n601 10.4732
R495 VTAIL.n571 VTAIL.n482 10.4732
R496 VTAIL.n544 VTAIL.n494 10.4732
R497 VTAIL.n523 VTAIL.n505 10.4732
R498 VTAIL.n475 VTAIL.n386 10.4732
R499 VTAIL.n448 VTAIL.n398 10.4732
R500 VTAIL.n427 VTAIL.n409 10.4732
R501 VTAIL.n379 VTAIL.n290 10.4732
R502 VTAIL.n352 VTAIL.n302 10.4732
R503 VTAIL.n331 VTAIL.n313 10.4732
R504 VTAIL.n703 VTAIL.n702 10.2747
R505 VTAIL.n31 VTAIL.n30 10.2747
R506 VTAIL.n127 VTAIL.n126 10.2747
R507 VTAIL.n223 VTAIL.n222 10.2747
R508 VTAIL.n608 VTAIL.n607 10.2747
R509 VTAIL.n512 VTAIL.n511 10.2747
R510 VTAIL.n416 VTAIL.n415 10.2747
R511 VTAIL.n320 VTAIL.n319 10.2747
R512 VTAIL.n713 VTAIL.n698 9.69747
R513 VTAIL.n740 VTAIL.n739 9.69747
R514 VTAIL.n760 VTAIL.n759 9.69747
R515 VTAIL.n41 VTAIL.n26 9.69747
R516 VTAIL.n68 VTAIL.n67 9.69747
R517 VTAIL.n88 VTAIL.n87 9.69747
R518 VTAIL.n137 VTAIL.n122 9.69747
R519 VTAIL.n164 VTAIL.n163 9.69747
R520 VTAIL.n184 VTAIL.n183 9.69747
R521 VTAIL.n233 VTAIL.n218 9.69747
R522 VTAIL.n260 VTAIL.n259 9.69747
R523 VTAIL.n280 VTAIL.n279 9.69747
R524 VTAIL.n664 VTAIL.n663 9.69747
R525 VTAIL.n644 VTAIL.n643 9.69747
R526 VTAIL.n618 VTAIL.n603 9.69747
R527 VTAIL.n568 VTAIL.n567 9.69747
R528 VTAIL.n548 VTAIL.n547 9.69747
R529 VTAIL.n522 VTAIL.n507 9.69747
R530 VTAIL.n472 VTAIL.n471 9.69747
R531 VTAIL.n452 VTAIL.n451 9.69747
R532 VTAIL.n426 VTAIL.n411 9.69747
R533 VTAIL.n376 VTAIL.n375 9.69747
R534 VTAIL.n356 VTAIL.n355 9.69747
R535 VTAIL.n330 VTAIL.n315 9.69747
R536 VTAIL.n762 VTAIL.n672 9.45567
R537 VTAIL.n90 VTAIL.n0 9.45567
R538 VTAIL.n186 VTAIL.n96 9.45567
R539 VTAIL.n282 VTAIL.n192 9.45567
R540 VTAIL.n666 VTAIL.n576 9.45567
R541 VTAIL.n570 VTAIL.n480 9.45567
R542 VTAIL.n474 VTAIL.n384 9.45567
R543 VTAIL.n378 VTAIL.n288 9.45567
R544 VTAIL.n680 VTAIL.n679 9.3005
R545 VTAIL.n753 VTAIL.n752 9.3005
R546 VTAIL.n755 VTAIL.n754 9.3005
R547 VTAIL.n676 VTAIL.n675 9.3005
R548 VTAIL.n761 VTAIL.n760 9.3005
R549 VTAIL.n763 VTAIL.n762 9.3005
R550 VTAIL.n745 VTAIL.n744 9.3005
R551 VTAIL.n684 VTAIL.n683 9.3005
R552 VTAIL.n739 VTAIL.n738 9.3005
R553 VTAIL.n737 VTAIL.n736 9.3005
R554 VTAIL.n688 VTAIL.n687 9.3005
R555 VTAIL.n731 VTAIL.n730 9.3005
R556 VTAIL.n729 VTAIL.n728 9.3005
R557 VTAIL.n705 VTAIL.n704 9.3005
R558 VTAIL.n700 VTAIL.n699 9.3005
R559 VTAIL.n711 VTAIL.n710 9.3005
R560 VTAIL.n713 VTAIL.n712 9.3005
R561 VTAIL.n696 VTAIL.n695 9.3005
R562 VTAIL.n719 VTAIL.n718 9.3005
R563 VTAIL.n721 VTAIL.n720 9.3005
R564 VTAIL.n722 VTAIL.n691 9.3005
R565 VTAIL.n747 VTAIL.n746 9.3005
R566 VTAIL.n8 VTAIL.n7 9.3005
R567 VTAIL.n81 VTAIL.n80 9.3005
R568 VTAIL.n83 VTAIL.n82 9.3005
R569 VTAIL.n4 VTAIL.n3 9.3005
R570 VTAIL.n89 VTAIL.n88 9.3005
R571 VTAIL.n91 VTAIL.n90 9.3005
R572 VTAIL.n73 VTAIL.n72 9.3005
R573 VTAIL.n12 VTAIL.n11 9.3005
R574 VTAIL.n67 VTAIL.n66 9.3005
R575 VTAIL.n65 VTAIL.n64 9.3005
R576 VTAIL.n16 VTAIL.n15 9.3005
R577 VTAIL.n59 VTAIL.n58 9.3005
R578 VTAIL.n57 VTAIL.n56 9.3005
R579 VTAIL.n33 VTAIL.n32 9.3005
R580 VTAIL.n28 VTAIL.n27 9.3005
R581 VTAIL.n39 VTAIL.n38 9.3005
R582 VTAIL.n41 VTAIL.n40 9.3005
R583 VTAIL.n24 VTAIL.n23 9.3005
R584 VTAIL.n47 VTAIL.n46 9.3005
R585 VTAIL.n49 VTAIL.n48 9.3005
R586 VTAIL.n50 VTAIL.n19 9.3005
R587 VTAIL.n75 VTAIL.n74 9.3005
R588 VTAIL.n104 VTAIL.n103 9.3005
R589 VTAIL.n177 VTAIL.n176 9.3005
R590 VTAIL.n179 VTAIL.n178 9.3005
R591 VTAIL.n100 VTAIL.n99 9.3005
R592 VTAIL.n185 VTAIL.n184 9.3005
R593 VTAIL.n187 VTAIL.n186 9.3005
R594 VTAIL.n169 VTAIL.n168 9.3005
R595 VTAIL.n108 VTAIL.n107 9.3005
R596 VTAIL.n163 VTAIL.n162 9.3005
R597 VTAIL.n161 VTAIL.n160 9.3005
R598 VTAIL.n112 VTAIL.n111 9.3005
R599 VTAIL.n155 VTAIL.n154 9.3005
R600 VTAIL.n153 VTAIL.n152 9.3005
R601 VTAIL.n129 VTAIL.n128 9.3005
R602 VTAIL.n124 VTAIL.n123 9.3005
R603 VTAIL.n135 VTAIL.n134 9.3005
R604 VTAIL.n137 VTAIL.n136 9.3005
R605 VTAIL.n120 VTAIL.n119 9.3005
R606 VTAIL.n143 VTAIL.n142 9.3005
R607 VTAIL.n145 VTAIL.n144 9.3005
R608 VTAIL.n146 VTAIL.n115 9.3005
R609 VTAIL.n171 VTAIL.n170 9.3005
R610 VTAIL.n200 VTAIL.n199 9.3005
R611 VTAIL.n273 VTAIL.n272 9.3005
R612 VTAIL.n275 VTAIL.n274 9.3005
R613 VTAIL.n196 VTAIL.n195 9.3005
R614 VTAIL.n281 VTAIL.n280 9.3005
R615 VTAIL.n283 VTAIL.n282 9.3005
R616 VTAIL.n265 VTAIL.n264 9.3005
R617 VTAIL.n204 VTAIL.n203 9.3005
R618 VTAIL.n259 VTAIL.n258 9.3005
R619 VTAIL.n257 VTAIL.n256 9.3005
R620 VTAIL.n208 VTAIL.n207 9.3005
R621 VTAIL.n251 VTAIL.n250 9.3005
R622 VTAIL.n249 VTAIL.n248 9.3005
R623 VTAIL.n225 VTAIL.n224 9.3005
R624 VTAIL.n220 VTAIL.n219 9.3005
R625 VTAIL.n231 VTAIL.n230 9.3005
R626 VTAIL.n233 VTAIL.n232 9.3005
R627 VTAIL.n216 VTAIL.n215 9.3005
R628 VTAIL.n239 VTAIL.n238 9.3005
R629 VTAIL.n241 VTAIL.n240 9.3005
R630 VTAIL.n242 VTAIL.n211 9.3005
R631 VTAIL.n267 VTAIL.n266 9.3005
R632 VTAIL.n667 VTAIL.n666 9.3005
R633 VTAIL.n665 VTAIL.n664 9.3005
R634 VTAIL.n580 VTAIL.n579 9.3005
R635 VTAIL.n659 VTAIL.n658 9.3005
R636 VTAIL.n657 VTAIL.n656 9.3005
R637 VTAIL.n584 VTAIL.n583 9.3005
R638 VTAIL.n651 VTAIL.n650 9.3005
R639 VTAIL.n649 VTAIL.n648 9.3005
R640 VTAIL.n588 VTAIL.n587 9.3005
R641 VTAIL.n643 VTAIL.n642 9.3005
R642 VTAIL.n641 VTAIL.n640 9.3005
R643 VTAIL.n592 VTAIL.n591 9.3005
R644 VTAIL.n635 VTAIL.n634 9.3005
R645 VTAIL.n633 VTAIL.n632 9.3005
R646 VTAIL.n598 VTAIL.n595 9.3005
R647 VTAIL.n626 VTAIL.n625 9.3005
R648 VTAIL.n624 VTAIL.n623 9.3005
R649 VTAIL.n601 VTAIL.n600 9.3005
R650 VTAIL.n618 VTAIL.n617 9.3005
R651 VTAIL.n616 VTAIL.n615 9.3005
R652 VTAIL.n605 VTAIL.n604 9.3005
R653 VTAIL.n610 VTAIL.n609 9.3005
R654 VTAIL.n514 VTAIL.n513 9.3005
R655 VTAIL.n509 VTAIL.n508 9.3005
R656 VTAIL.n520 VTAIL.n519 9.3005
R657 VTAIL.n522 VTAIL.n521 9.3005
R658 VTAIL.n505 VTAIL.n504 9.3005
R659 VTAIL.n528 VTAIL.n527 9.3005
R660 VTAIL.n530 VTAIL.n529 9.3005
R661 VTAIL.n502 VTAIL.n499 9.3005
R662 VTAIL.n561 VTAIL.n560 9.3005
R663 VTAIL.n563 VTAIL.n562 9.3005
R664 VTAIL.n484 VTAIL.n483 9.3005
R665 VTAIL.n569 VTAIL.n568 9.3005
R666 VTAIL.n571 VTAIL.n570 9.3005
R667 VTAIL.n488 VTAIL.n487 9.3005
R668 VTAIL.n555 VTAIL.n554 9.3005
R669 VTAIL.n553 VTAIL.n552 9.3005
R670 VTAIL.n492 VTAIL.n491 9.3005
R671 VTAIL.n547 VTAIL.n546 9.3005
R672 VTAIL.n545 VTAIL.n544 9.3005
R673 VTAIL.n496 VTAIL.n495 9.3005
R674 VTAIL.n539 VTAIL.n538 9.3005
R675 VTAIL.n537 VTAIL.n536 9.3005
R676 VTAIL.n418 VTAIL.n417 9.3005
R677 VTAIL.n413 VTAIL.n412 9.3005
R678 VTAIL.n424 VTAIL.n423 9.3005
R679 VTAIL.n426 VTAIL.n425 9.3005
R680 VTAIL.n409 VTAIL.n408 9.3005
R681 VTAIL.n432 VTAIL.n431 9.3005
R682 VTAIL.n434 VTAIL.n433 9.3005
R683 VTAIL.n406 VTAIL.n403 9.3005
R684 VTAIL.n465 VTAIL.n464 9.3005
R685 VTAIL.n467 VTAIL.n466 9.3005
R686 VTAIL.n388 VTAIL.n387 9.3005
R687 VTAIL.n473 VTAIL.n472 9.3005
R688 VTAIL.n475 VTAIL.n474 9.3005
R689 VTAIL.n392 VTAIL.n391 9.3005
R690 VTAIL.n459 VTAIL.n458 9.3005
R691 VTAIL.n457 VTAIL.n456 9.3005
R692 VTAIL.n396 VTAIL.n395 9.3005
R693 VTAIL.n451 VTAIL.n450 9.3005
R694 VTAIL.n449 VTAIL.n448 9.3005
R695 VTAIL.n400 VTAIL.n399 9.3005
R696 VTAIL.n443 VTAIL.n442 9.3005
R697 VTAIL.n441 VTAIL.n440 9.3005
R698 VTAIL.n322 VTAIL.n321 9.3005
R699 VTAIL.n317 VTAIL.n316 9.3005
R700 VTAIL.n328 VTAIL.n327 9.3005
R701 VTAIL.n330 VTAIL.n329 9.3005
R702 VTAIL.n313 VTAIL.n312 9.3005
R703 VTAIL.n336 VTAIL.n335 9.3005
R704 VTAIL.n338 VTAIL.n337 9.3005
R705 VTAIL.n310 VTAIL.n307 9.3005
R706 VTAIL.n369 VTAIL.n368 9.3005
R707 VTAIL.n371 VTAIL.n370 9.3005
R708 VTAIL.n292 VTAIL.n291 9.3005
R709 VTAIL.n377 VTAIL.n376 9.3005
R710 VTAIL.n379 VTAIL.n378 9.3005
R711 VTAIL.n296 VTAIL.n295 9.3005
R712 VTAIL.n363 VTAIL.n362 9.3005
R713 VTAIL.n361 VTAIL.n360 9.3005
R714 VTAIL.n300 VTAIL.n299 9.3005
R715 VTAIL.n355 VTAIL.n354 9.3005
R716 VTAIL.n353 VTAIL.n352 9.3005
R717 VTAIL.n304 VTAIL.n303 9.3005
R718 VTAIL.n347 VTAIL.n346 9.3005
R719 VTAIL.n345 VTAIL.n344 9.3005
R720 VTAIL.n710 VTAIL.n709 8.92171
R721 VTAIL.n743 VTAIL.n684 8.92171
R722 VTAIL.n756 VTAIL.n676 8.92171
R723 VTAIL.n38 VTAIL.n37 8.92171
R724 VTAIL.n71 VTAIL.n12 8.92171
R725 VTAIL.n84 VTAIL.n4 8.92171
R726 VTAIL.n134 VTAIL.n133 8.92171
R727 VTAIL.n167 VTAIL.n108 8.92171
R728 VTAIL.n180 VTAIL.n100 8.92171
R729 VTAIL.n230 VTAIL.n229 8.92171
R730 VTAIL.n263 VTAIL.n204 8.92171
R731 VTAIL.n276 VTAIL.n196 8.92171
R732 VTAIL.n660 VTAIL.n580 8.92171
R733 VTAIL.n647 VTAIL.n588 8.92171
R734 VTAIL.n615 VTAIL.n614 8.92171
R735 VTAIL.n564 VTAIL.n484 8.92171
R736 VTAIL.n551 VTAIL.n492 8.92171
R737 VTAIL.n519 VTAIL.n518 8.92171
R738 VTAIL.n468 VTAIL.n388 8.92171
R739 VTAIL.n455 VTAIL.n396 8.92171
R740 VTAIL.n423 VTAIL.n422 8.92171
R741 VTAIL.n372 VTAIL.n292 8.92171
R742 VTAIL.n359 VTAIL.n300 8.92171
R743 VTAIL.n327 VTAIL.n326 8.92171
R744 VTAIL.n706 VTAIL.n700 8.14595
R745 VTAIL.n744 VTAIL.n682 8.14595
R746 VTAIL.n755 VTAIL.n678 8.14595
R747 VTAIL.n34 VTAIL.n28 8.14595
R748 VTAIL.n72 VTAIL.n10 8.14595
R749 VTAIL.n83 VTAIL.n6 8.14595
R750 VTAIL.n130 VTAIL.n124 8.14595
R751 VTAIL.n168 VTAIL.n106 8.14595
R752 VTAIL.n179 VTAIL.n102 8.14595
R753 VTAIL.n226 VTAIL.n220 8.14595
R754 VTAIL.n264 VTAIL.n202 8.14595
R755 VTAIL.n275 VTAIL.n198 8.14595
R756 VTAIL.n659 VTAIL.n582 8.14595
R757 VTAIL.n648 VTAIL.n586 8.14595
R758 VTAIL.n611 VTAIL.n605 8.14595
R759 VTAIL.n563 VTAIL.n486 8.14595
R760 VTAIL.n552 VTAIL.n490 8.14595
R761 VTAIL.n515 VTAIL.n509 8.14595
R762 VTAIL.n467 VTAIL.n390 8.14595
R763 VTAIL.n456 VTAIL.n394 8.14595
R764 VTAIL.n419 VTAIL.n413 8.14595
R765 VTAIL.n371 VTAIL.n294 8.14595
R766 VTAIL.n360 VTAIL.n298 8.14595
R767 VTAIL.n323 VTAIL.n317 8.14595
R768 VTAIL.n705 VTAIL.n702 7.3702
R769 VTAIL.n748 VTAIL.n747 7.3702
R770 VTAIL.n752 VTAIL.n751 7.3702
R771 VTAIL.n33 VTAIL.n30 7.3702
R772 VTAIL.n76 VTAIL.n75 7.3702
R773 VTAIL.n80 VTAIL.n79 7.3702
R774 VTAIL.n129 VTAIL.n126 7.3702
R775 VTAIL.n172 VTAIL.n171 7.3702
R776 VTAIL.n176 VTAIL.n175 7.3702
R777 VTAIL.n225 VTAIL.n222 7.3702
R778 VTAIL.n268 VTAIL.n267 7.3702
R779 VTAIL.n272 VTAIL.n271 7.3702
R780 VTAIL.n656 VTAIL.n655 7.3702
R781 VTAIL.n652 VTAIL.n651 7.3702
R782 VTAIL.n610 VTAIL.n607 7.3702
R783 VTAIL.n560 VTAIL.n559 7.3702
R784 VTAIL.n556 VTAIL.n555 7.3702
R785 VTAIL.n514 VTAIL.n511 7.3702
R786 VTAIL.n464 VTAIL.n463 7.3702
R787 VTAIL.n460 VTAIL.n459 7.3702
R788 VTAIL.n418 VTAIL.n415 7.3702
R789 VTAIL.n368 VTAIL.n367 7.3702
R790 VTAIL.n364 VTAIL.n363 7.3702
R791 VTAIL.n322 VTAIL.n319 7.3702
R792 VTAIL.n748 VTAIL.n680 6.59444
R793 VTAIL.n751 VTAIL.n680 6.59444
R794 VTAIL.n76 VTAIL.n8 6.59444
R795 VTAIL.n79 VTAIL.n8 6.59444
R796 VTAIL.n172 VTAIL.n104 6.59444
R797 VTAIL.n175 VTAIL.n104 6.59444
R798 VTAIL.n268 VTAIL.n200 6.59444
R799 VTAIL.n271 VTAIL.n200 6.59444
R800 VTAIL.n655 VTAIL.n584 6.59444
R801 VTAIL.n652 VTAIL.n584 6.59444
R802 VTAIL.n559 VTAIL.n488 6.59444
R803 VTAIL.n556 VTAIL.n488 6.59444
R804 VTAIL.n463 VTAIL.n392 6.59444
R805 VTAIL.n460 VTAIL.n392 6.59444
R806 VTAIL.n367 VTAIL.n296 6.59444
R807 VTAIL.n364 VTAIL.n296 6.59444
R808 VTAIL.n706 VTAIL.n705 5.81868
R809 VTAIL.n747 VTAIL.n682 5.81868
R810 VTAIL.n752 VTAIL.n678 5.81868
R811 VTAIL.n34 VTAIL.n33 5.81868
R812 VTAIL.n75 VTAIL.n10 5.81868
R813 VTAIL.n80 VTAIL.n6 5.81868
R814 VTAIL.n130 VTAIL.n129 5.81868
R815 VTAIL.n171 VTAIL.n106 5.81868
R816 VTAIL.n176 VTAIL.n102 5.81868
R817 VTAIL.n226 VTAIL.n225 5.81868
R818 VTAIL.n267 VTAIL.n202 5.81868
R819 VTAIL.n272 VTAIL.n198 5.81868
R820 VTAIL.n656 VTAIL.n582 5.81868
R821 VTAIL.n651 VTAIL.n586 5.81868
R822 VTAIL.n611 VTAIL.n610 5.81868
R823 VTAIL.n560 VTAIL.n486 5.81868
R824 VTAIL.n555 VTAIL.n490 5.81868
R825 VTAIL.n515 VTAIL.n514 5.81868
R826 VTAIL.n464 VTAIL.n390 5.81868
R827 VTAIL.n459 VTAIL.n394 5.81868
R828 VTAIL.n419 VTAIL.n418 5.81868
R829 VTAIL.n368 VTAIL.n294 5.81868
R830 VTAIL.n363 VTAIL.n298 5.81868
R831 VTAIL.n323 VTAIL.n322 5.81868
R832 VTAIL.n709 VTAIL.n700 5.04292
R833 VTAIL.n744 VTAIL.n743 5.04292
R834 VTAIL.n756 VTAIL.n755 5.04292
R835 VTAIL.n37 VTAIL.n28 5.04292
R836 VTAIL.n72 VTAIL.n71 5.04292
R837 VTAIL.n84 VTAIL.n83 5.04292
R838 VTAIL.n133 VTAIL.n124 5.04292
R839 VTAIL.n168 VTAIL.n167 5.04292
R840 VTAIL.n180 VTAIL.n179 5.04292
R841 VTAIL.n229 VTAIL.n220 5.04292
R842 VTAIL.n264 VTAIL.n263 5.04292
R843 VTAIL.n276 VTAIL.n275 5.04292
R844 VTAIL.n660 VTAIL.n659 5.04292
R845 VTAIL.n648 VTAIL.n647 5.04292
R846 VTAIL.n614 VTAIL.n605 5.04292
R847 VTAIL.n564 VTAIL.n563 5.04292
R848 VTAIL.n552 VTAIL.n551 5.04292
R849 VTAIL.n518 VTAIL.n509 5.04292
R850 VTAIL.n468 VTAIL.n467 5.04292
R851 VTAIL.n456 VTAIL.n455 5.04292
R852 VTAIL.n422 VTAIL.n413 5.04292
R853 VTAIL.n372 VTAIL.n371 5.04292
R854 VTAIL.n360 VTAIL.n359 5.04292
R855 VTAIL.n326 VTAIL.n317 5.04292
R856 VTAIL.n710 VTAIL.n698 4.26717
R857 VTAIL.n740 VTAIL.n684 4.26717
R858 VTAIL.n759 VTAIL.n676 4.26717
R859 VTAIL.n38 VTAIL.n26 4.26717
R860 VTAIL.n68 VTAIL.n12 4.26717
R861 VTAIL.n87 VTAIL.n4 4.26717
R862 VTAIL.n134 VTAIL.n122 4.26717
R863 VTAIL.n164 VTAIL.n108 4.26717
R864 VTAIL.n183 VTAIL.n100 4.26717
R865 VTAIL.n230 VTAIL.n218 4.26717
R866 VTAIL.n260 VTAIL.n204 4.26717
R867 VTAIL.n279 VTAIL.n196 4.26717
R868 VTAIL.n663 VTAIL.n580 4.26717
R869 VTAIL.n644 VTAIL.n588 4.26717
R870 VTAIL.n615 VTAIL.n603 4.26717
R871 VTAIL.n567 VTAIL.n484 4.26717
R872 VTAIL.n548 VTAIL.n492 4.26717
R873 VTAIL.n519 VTAIL.n507 4.26717
R874 VTAIL.n471 VTAIL.n388 4.26717
R875 VTAIL.n452 VTAIL.n396 4.26717
R876 VTAIL.n423 VTAIL.n411 4.26717
R877 VTAIL.n375 VTAIL.n292 4.26717
R878 VTAIL.n356 VTAIL.n300 4.26717
R879 VTAIL.n327 VTAIL.n315 4.26717
R880 VTAIL.n714 VTAIL.n713 3.49141
R881 VTAIL.n739 VTAIL.n686 3.49141
R882 VTAIL.n760 VTAIL.n674 3.49141
R883 VTAIL.n42 VTAIL.n41 3.49141
R884 VTAIL.n67 VTAIL.n14 3.49141
R885 VTAIL.n88 VTAIL.n2 3.49141
R886 VTAIL.n138 VTAIL.n137 3.49141
R887 VTAIL.n163 VTAIL.n110 3.49141
R888 VTAIL.n184 VTAIL.n98 3.49141
R889 VTAIL.n234 VTAIL.n233 3.49141
R890 VTAIL.n259 VTAIL.n206 3.49141
R891 VTAIL.n280 VTAIL.n194 3.49141
R892 VTAIL.n664 VTAIL.n578 3.49141
R893 VTAIL.n643 VTAIL.n590 3.49141
R894 VTAIL.n619 VTAIL.n618 3.49141
R895 VTAIL.n568 VTAIL.n482 3.49141
R896 VTAIL.n547 VTAIL.n494 3.49141
R897 VTAIL.n523 VTAIL.n522 3.49141
R898 VTAIL.n472 VTAIL.n386 3.49141
R899 VTAIL.n451 VTAIL.n398 3.49141
R900 VTAIL.n427 VTAIL.n426 3.49141
R901 VTAIL.n376 VTAIL.n290 3.49141
R902 VTAIL.n355 VTAIL.n302 3.49141
R903 VTAIL.n331 VTAIL.n330 3.49141
R904 VTAIL.n704 VTAIL.n703 2.84303
R905 VTAIL.n32 VTAIL.n31 2.84303
R906 VTAIL.n128 VTAIL.n127 2.84303
R907 VTAIL.n224 VTAIL.n223 2.84303
R908 VTAIL.n609 VTAIL.n608 2.84303
R909 VTAIL.n513 VTAIL.n512 2.84303
R910 VTAIL.n417 VTAIL.n416 2.84303
R911 VTAIL.n321 VTAIL.n320 2.84303
R912 VTAIL.n717 VTAIL.n696 2.71565
R913 VTAIL.n736 VTAIL.n735 2.71565
R914 VTAIL.n764 VTAIL.n763 2.71565
R915 VTAIL.n45 VTAIL.n24 2.71565
R916 VTAIL.n64 VTAIL.n63 2.71565
R917 VTAIL.n92 VTAIL.n91 2.71565
R918 VTAIL.n141 VTAIL.n120 2.71565
R919 VTAIL.n160 VTAIL.n159 2.71565
R920 VTAIL.n188 VTAIL.n187 2.71565
R921 VTAIL.n237 VTAIL.n216 2.71565
R922 VTAIL.n256 VTAIL.n255 2.71565
R923 VTAIL.n284 VTAIL.n283 2.71565
R924 VTAIL.n668 VTAIL.n667 2.71565
R925 VTAIL.n640 VTAIL.n639 2.71565
R926 VTAIL.n622 VTAIL.n601 2.71565
R927 VTAIL.n572 VTAIL.n571 2.71565
R928 VTAIL.n544 VTAIL.n543 2.71565
R929 VTAIL.n526 VTAIL.n505 2.71565
R930 VTAIL.n476 VTAIL.n475 2.71565
R931 VTAIL.n448 VTAIL.n447 2.71565
R932 VTAIL.n430 VTAIL.n409 2.71565
R933 VTAIL.n380 VTAIL.n379 2.71565
R934 VTAIL.n352 VTAIL.n351 2.71565
R935 VTAIL.n334 VTAIL.n313 2.71565
R936 VTAIL.n479 VTAIL.n383 1.9574
R937 VTAIL.n671 VTAIL.n575 1.9574
R938 VTAIL.n287 VTAIL.n191 1.9574
R939 VTAIL.n718 VTAIL.n694 1.93989
R940 VTAIL.n732 VTAIL.n688 1.93989
R941 VTAIL.n766 VTAIL.n672 1.93989
R942 VTAIL.n46 VTAIL.n22 1.93989
R943 VTAIL.n60 VTAIL.n16 1.93989
R944 VTAIL.n94 VTAIL.n0 1.93989
R945 VTAIL.n142 VTAIL.n118 1.93989
R946 VTAIL.n156 VTAIL.n112 1.93989
R947 VTAIL.n190 VTAIL.n96 1.93989
R948 VTAIL.n238 VTAIL.n214 1.93989
R949 VTAIL.n252 VTAIL.n208 1.93989
R950 VTAIL.n286 VTAIL.n192 1.93989
R951 VTAIL.n670 VTAIL.n576 1.93989
R952 VTAIL.n636 VTAIL.n592 1.93989
R953 VTAIL.n623 VTAIL.n599 1.93989
R954 VTAIL.n574 VTAIL.n480 1.93989
R955 VTAIL.n540 VTAIL.n496 1.93989
R956 VTAIL.n527 VTAIL.n503 1.93989
R957 VTAIL.n478 VTAIL.n384 1.93989
R958 VTAIL.n444 VTAIL.n400 1.93989
R959 VTAIL.n431 VTAIL.n407 1.93989
R960 VTAIL.n382 VTAIL.n288 1.93989
R961 VTAIL.n348 VTAIL.n304 1.93989
R962 VTAIL.n335 VTAIL.n311 1.93989
R963 VTAIL.n723 VTAIL.n721 1.16414
R964 VTAIL.n731 VTAIL.n690 1.16414
R965 VTAIL.n51 VTAIL.n49 1.16414
R966 VTAIL.n59 VTAIL.n18 1.16414
R967 VTAIL.n147 VTAIL.n145 1.16414
R968 VTAIL.n155 VTAIL.n114 1.16414
R969 VTAIL.n243 VTAIL.n241 1.16414
R970 VTAIL.n251 VTAIL.n210 1.16414
R971 VTAIL.n635 VTAIL.n594 1.16414
R972 VTAIL.n627 VTAIL.n626 1.16414
R973 VTAIL.n539 VTAIL.n498 1.16414
R974 VTAIL.n531 VTAIL.n530 1.16414
R975 VTAIL.n443 VTAIL.n402 1.16414
R976 VTAIL.n435 VTAIL.n434 1.16414
R977 VTAIL.n347 VTAIL.n306 1.16414
R978 VTAIL.n339 VTAIL.n338 1.16414
R979 VTAIL VTAIL.n95 1.03714
R980 VTAIL VTAIL.n767 0.920759
R981 VTAIL.n575 VTAIL.n479 0.470328
R982 VTAIL.n191 VTAIL.n95 0.470328
R983 VTAIL.n722 VTAIL.n692 0.388379
R984 VTAIL.n728 VTAIL.n727 0.388379
R985 VTAIL.n50 VTAIL.n20 0.388379
R986 VTAIL.n56 VTAIL.n55 0.388379
R987 VTAIL.n146 VTAIL.n116 0.388379
R988 VTAIL.n152 VTAIL.n151 0.388379
R989 VTAIL.n242 VTAIL.n212 0.388379
R990 VTAIL.n248 VTAIL.n247 0.388379
R991 VTAIL.n632 VTAIL.n631 0.388379
R992 VTAIL.n598 VTAIL.n596 0.388379
R993 VTAIL.n536 VTAIL.n535 0.388379
R994 VTAIL.n502 VTAIL.n500 0.388379
R995 VTAIL.n440 VTAIL.n439 0.388379
R996 VTAIL.n406 VTAIL.n404 0.388379
R997 VTAIL.n344 VTAIL.n343 0.388379
R998 VTAIL.n310 VTAIL.n308 0.388379
R999 VTAIL.n704 VTAIL.n699 0.155672
R1000 VTAIL.n711 VTAIL.n699 0.155672
R1001 VTAIL.n712 VTAIL.n711 0.155672
R1002 VTAIL.n712 VTAIL.n695 0.155672
R1003 VTAIL.n719 VTAIL.n695 0.155672
R1004 VTAIL.n720 VTAIL.n719 0.155672
R1005 VTAIL.n720 VTAIL.n691 0.155672
R1006 VTAIL.n729 VTAIL.n691 0.155672
R1007 VTAIL.n730 VTAIL.n729 0.155672
R1008 VTAIL.n730 VTAIL.n687 0.155672
R1009 VTAIL.n737 VTAIL.n687 0.155672
R1010 VTAIL.n738 VTAIL.n737 0.155672
R1011 VTAIL.n738 VTAIL.n683 0.155672
R1012 VTAIL.n745 VTAIL.n683 0.155672
R1013 VTAIL.n746 VTAIL.n745 0.155672
R1014 VTAIL.n746 VTAIL.n679 0.155672
R1015 VTAIL.n753 VTAIL.n679 0.155672
R1016 VTAIL.n754 VTAIL.n753 0.155672
R1017 VTAIL.n754 VTAIL.n675 0.155672
R1018 VTAIL.n761 VTAIL.n675 0.155672
R1019 VTAIL.n762 VTAIL.n761 0.155672
R1020 VTAIL.n32 VTAIL.n27 0.155672
R1021 VTAIL.n39 VTAIL.n27 0.155672
R1022 VTAIL.n40 VTAIL.n39 0.155672
R1023 VTAIL.n40 VTAIL.n23 0.155672
R1024 VTAIL.n47 VTAIL.n23 0.155672
R1025 VTAIL.n48 VTAIL.n47 0.155672
R1026 VTAIL.n48 VTAIL.n19 0.155672
R1027 VTAIL.n57 VTAIL.n19 0.155672
R1028 VTAIL.n58 VTAIL.n57 0.155672
R1029 VTAIL.n58 VTAIL.n15 0.155672
R1030 VTAIL.n65 VTAIL.n15 0.155672
R1031 VTAIL.n66 VTAIL.n65 0.155672
R1032 VTAIL.n66 VTAIL.n11 0.155672
R1033 VTAIL.n73 VTAIL.n11 0.155672
R1034 VTAIL.n74 VTAIL.n73 0.155672
R1035 VTAIL.n74 VTAIL.n7 0.155672
R1036 VTAIL.n81 VTAIL.n7 0.155672
R1037 VTAIL.n82 VTAIL.n81 0.155672
R1038 VTAIL.n82 VTAIL.n3 0.155672
R1039 VTAIL.n89 VTAIL.n3 0.155672
R1040 VTAIL.n90 VTAIL.n89 0.155672
R1041 VTAIL.n128 VTAIL.n123 0.155672
R1042 VTAIL.n135 VTAIL.n123 0.155672
R1043 VTAIL.n136 VTAIL.n135 0.155672
R1044 VTAIL.n136 VTAIL.n119 0.155672
R1045 VTAIL.n143 VTAIL.n119 0.155672
R1046 VTAIL.n144 VTAIL.n143 0.155672
R1047 VTAIL.n144 VTAIL.n115 0.155672
R1048 VTAIL.n153 VTAIL.n115 0.155672
R1049 VTAIL.n154 VTAIL.n153 0.155672
R1050 VTAIL.n154 VTAIL.n111 0.155672
R1051 VTAIL.n161 VTAIL.n111 0.155672
R1052 VTAIL.n162 VTAIL.n161 0.155672
R1053 VTAIL.n162 VTAIL.n107 0.155672
R1054 VTAIL.n169 VTAIL.n107 0.155672
R1055 VTAIL.n170 VTAIL.n169 0.155672
R1056 VTAIL.n170 VTAIL.n103 0.155672
R1057 VTAIL.n177 VTAIL.n103 0.155672
R1058 VTAIL.n178 VTAIL.n177 0.155672
R1059 VTAIL.n178 VTAIL.n99 0.155672
R1060 VTAIL.n185 VTAIL.n99 0.155672
R1061 VTAIL.n186 VTAIL.n185 0.155672
R1062 VTAIL.n224 VTAIL.n219 0.155672
R1063 VTAIL.n231 VTAIL.n219 0.155672
R1064 VTAIL.n232 VTAIL.n231 0.155672
R1065 VTAIL.n232 VTAIL.n215 0.155672
R1066 VTAIL.n239 VTAIL.n215 0.155672
R1067 VTAIL.n240 VTAIL.n239 0.155672
R1068 VTAIL.n240 VTAIL.n211 0.155672
R1069 VTAIL.n249 VTAIL.n211 0.155672
R1070 VTAIL.n250 VTAIL.n249 0.155672
R1071 VTAIL.n250 VTAIL.n207 0.155672
R1072 VTAIL.n257 VTAIL.n207 0.155672
R1073 VTAIL.n258 VTAIL.n257 0.155672
R1074 VTAIL.n258 VTAIL.n203 0.155672
R1075 VTAIL.n265 VTAIL.n203 0.155672
R1076 VTAIL.n266 VTAIL.n265 0.155672
R1077 VTAIL.n266 VTAIL.n199 0.155672
R1078 VTAIL.n273 VTAIL.n199 0.155672
R1079 VTAIL.n274 VTAIL.n273 0.155672
R1080 VTAIL.n274 VTAIL.n195 0.155672
R1081 VTAIL.n281 VTAIL.n195 0.155672
R1082 VTAIL.n282 VTAIL.n281 0.155672
R1083 VTAIL.n666 VTAIL.n665 0.155672
R1084 VTAIL.n665 VTAIL.n579 0.155672
R1085 VTAIL.n658 VTAIL.n579 0.155672
R1086 VTAIL.n658 VTAIL.n657 0.155672
R1087 VTAIL.n657 VTAIL.n583 0.155672
R1088 VTAIL.n650 VTAIL.n583 0.155672
R1089 VTAIL.n650 VTAIL.n649 0.155672
R1090 VTAIL.n649 VTAIL.n587 0.155672
R1091 VTAIL.n642 VTAIL.n587 0.155672
R1092 VTAIL.n642 VTAIL.n641 0.155672
R1093 VTAIL.n641 VTAIL.n591 0.155672
R1094 VTAIL.n634 VTAIL.n591 0.155672
R1095 VTAIL.n634 VTAIL.n633 0.155672
R1096 VTAIL.n633 VTAIL.n595 0.155672
R1097 VTAIL.n625 VTAIL.n595 0.155672
R1098 VTAIL.n625 VTAIL.n624 0.155672
R1099 VTAIL.n624 VTAIL.n600 0.155672
R1100 VTAIL.n617 VTAIL.n600 0.155672
R1101 VTAIL.n617 VTAIL.n616 0.155672
R1102 VTAIL.n616 VTAIL.n604 0.155672
R1103 VTAIL.n609 VTAIL.n604 0.155672
R1104 VTAIL.n570 VTAIL.n569 0.155672
R1105 VTAIL.n569 VTAIL.n483 0.155672
R1106 VTAIL.n562 VTAIL.n483 0.155672
R1107 VTAIL.n562 VTAIL.n561 0.155672
R1108 VTAIL.n561 VTAIL.n487 0.155672
R1109 VTAIL.n554 VTAIL.n487 0.155672
R1110 VTAIL.n554 VTAIL.n553 0.155672
R1111 VTAIL.n553 VTAIL.n491 0.155672
R1112 VTAIL.n546 VTAIL.n491 0.155672
R1113 VTAIL.n546 VTAIL.n545 0.155672
R1114 VTAIL.n545 VTAIL.n495 0.155672
R1115 VTAIL.n538 VTAIL.n495 0.155672
R1116 VTAIL.n538 VTAIL.n537 0.155672
R1117 VTAIL.n537 VTAIL.n499 0.155672
R1118 VTAIL.n529 VTAIL.n499 0.155672
R1119 VTAIL.n529 VTAIL.n528 0.155672
R1120 VTAIL.n528 VTAIL.n504 0.155672
R1121 VTAIL.n521 VTAIL.n504 0.155672
R1122 VTAIL.n521 VTAIL.n520 0.155672
R1123 VTAIL.n520 VTAIL.n508 0.155672
R1124 VTAIL.n513 VTAIL.n508 0.155672
R1125 VTAIL.n474 VTAIL.n473 0.155672
R1126 VTAIL.n473 VTAIL.n387 0.155672
R1127 VTAIL.n466 VTAIL.n387 0.155672
R1128 VTAIL.n466 VTAIL.n465 0.155672
R1129 VTAIL.n465 VTAIL.n391 0.155672
R1130 VTAIL.n458 VTAIL.n391 0.155672
R1131 VTAIL.n458 VTAIL.n457 0.155672
R1132 VTAIL.n457 VTAIL.n395 0.155672
R1133 VTAIL.n450 VTAIL.n395 0.155672
R1134 VTAIL.n450 VTAIL.n449 0.155672
R1135 VTAIL.n449 VTAIL.n399 0.155672
R1136 VTAIL.n442 VTAIL.n399 0.155672
R1137 VTAIL.n442 VTAIL.n441 0.155672
R1138 VTAIL.n441 VTAIL.n403 0.155672
R1139 VTAIL.n433 VTAIL.n403 0.155672
R1140 VTAIL.n433 VTAIL.n432 0.155672
R1141 VTAIL.n432 VTAIL.n408 0.155672
R1142 VTAIL.n425 VTAIL.n408 0.155672
R1143 VTAIL.n425 VTAIL.n424 0.155672
R1144 VTAIL.n424 VTAIL.n412 0.155672
R1145 VTAIL.n417 VTAIL.n412 0.155672
R1146 VTAIL.n378 VTAIL.n377 0.155672
R1147 VTAIL.n377 VTAIL.n291 0.155672
R1148 VTAIL.n370 VTAIL.n291 0.155672
R1149 VTAIL.n370 VTAIL.n369 0.155672
R1150 VTAIL.n369 VTAIL.n295 0.155672
R1151 VTAIL.n362 VTAIL.n295 0.155672
R1152 VTAIL.n362 VTAIL.n361 0.155672
R1153 VTAIL.n361 VTAIL.n299 0.155672
R1154 VTAIL.n354 VTAIL.n299 0.155672
R1155 VTAIL.n354 VTAIL.n353 0.155672
R1156 VTAIL.n353 VTAIL.n303 0.155672
R1157 VTAIL.n346 VTAIL.n303 0.155672
R1158 VTAIL.n346 VTAIL.n345 0.155672
R1159 VTAIL.n345 VTAIL.n307 0.155672
R1160 VTAIL.n337 VTAIL.n307 0.155672
R1161 VTAIL.n337 VTAIL.n336 0.155672
R1162 VTAIL.n336 VTAIL.n312 0.155672
R1163 VTAIL.n329 VTAIL.n312 0.155672
R1164 VTAIL.n329 VTAIL.n328 0.155672
R1165 VTAIL.n328 VTAIL.n316 0.155672
R1166 VTAIL.n321 VTAIL.n316 0.155672
R1167 VDD2.n2 VDD2.n0 109.285
R1168 VDD2.n2 VDD2.n1 64.6994
R1169 VDD2.n1 VDD2.t0 1.13843
R1170 VDD2.n1 VDD2.t1 1.13843
R1171 VDD2.n0 VDD2.t2 1.13843
R1172 VDD2.n0 VDD2.t3 1.13843
R1173 VDD2 VDD2.n2 0.0586897
R1174 B.n862 B.n861 585
R1175 B.n863 B.n862 585
R1176 B.n368 B.n117 585
R1177 B.n367 B.n366 585
R1178 B.n365 B.n364 585
R1179 B.n363 B.n362 585
R1180 B.n361 B.n360 585
R1181 B.n359 B.n358 585
R1182 B.n357 B.n356 585
R1183 B.n355 B.n354 585
R1184 B.n353 B.n352 585
R1185 B.n351 B.n350 585
R1186 B.n349 B.n348 585
R1187 B.n347 B.n346 585
R1188 B.n345 B.n344 585
R1189 B.n343 B.n342 585
R1190 B.n341 B.n340 585
R1191 B.n339 B.n338 585
R1192 B.n337 B.n336 585
R1193 B.n335 B.n334 585
R1194 B.n333 B.n332 585
R1195 B.n331 B.n330 585
R1196 B.n329 B.n328 585
R1197 B.n327 B.n326 585
R1198 B.n325 B.n324 585
R1199 B.n323 B.n322 585
R1200 B.n321 B.n320 585
R1201 B.n319 B.n318 585
R1202 B.n317 B.n316 585
R1203 B.n315 B.n314 585
R1204 B.n313 B.n312 585
R1205 B.n311 B.n310 585
R1206 B.n309 B.n308 585
R1207 B.n307 B.n306 585
R1208 B.n305 B.n304 585
R1209 B.n303 B.n302 585
R1210 B.n301 B.n300 585
R1211 B.n299 B.n298 585
R1212 B.n297 B.n296 585
R1213 B.n295 B.n294 585
R1214 B.n293 B.n292 585
R1215 B.n291 B.n290 585
R1216 B.n289 B.n288 585
R1217 B.n287 B.n286 585
R1218 B.n285 B.n284 585
R1219 B.n283 B.n282 585
R1220 B.n281 B.n280 585
R1221 B.n279 B.n278 585
R1222 B.n277 B.n276 585
R1223 B.n275 B.n274 585
R1224 B.n273 B.n272 585
R1225 B.n271 B.n270 585
R1226 B.n269 B.n268 585
R1227 B.n267 B.n266 585
R1228 B.n265 B.n264 585
R1229 B.n263 B.n262 585
R1230 B.n261 B.n260 585
R1231 B.n259 B.n258 585
R1232 B.n257 B.n256 585
R1233 B.n254 B.n253 585
R1234 B.n252 B.n251 585
R1235 B.n250 B.n249 585
R1236 B.n248 B.n247 585
R1237 B.n246 B.n245 585
R1238 B.n244 B.n243 585
R1239 B.n242 B.n241 585
R1240 B.n240 B.n239 585
R1241 B.n238 B.n237 585
R1242 B.n236 B.n235 585
R1243 B.n234 B.n233 585
R1244 B.n232 B.n231 585
R1245 B.n230 B.n229 585
R1246 B.n228 B.n227 585
R1247 B.n226 B.n225 585
R1248 B.n224 B.n223 585
R1249 B.n222 B.n221 585
R1250 B.n220 B.n219 585
R1251 B.n218 B.n217 585
R1252 B.n216 B.n215 585
R1253 B.n214 B.n213 585
R1254 B.n212 B.n211 585
R1255 B.n210 B.n209 585
R1256 B.n208 B.n207 585
R1257 B.n206 B.n205 585
R1258 B.n204 B.n203 585
R1259 B.n202 B.n201 585
R1260 B.n200 B.n199 585
R1261 B.n198 B.n197 585
R1262 B.n196 B.n195 585
R1263 B.n194 B.n193 585
R1264 B.n192 B.n191 585
R1265 B.n190 B.n189 585
R1266 B.n188 B.n187 585
R1267 B.n186 B.n185 585
R1268 B.n184 B.n183 585
R1269 B.n182 B.n181 585
R1270 B.n180 B.n179 585
R1271 B.n178 B.n177 585
R1272 B.n176 B.n175 585
R1273 B.n174 B.n173 585
R1274 B.n172 B.n171 585
R1275 B.n170 B.n169 585
R1276 B.n168 B.n167 585
R1277 B.n166 B.n165 585
R1278 B.n164 B.n163 585
R1279 B.n162 B.n161 585
R1280 B.n160 B.n159 585
R1281 B.n158 B.n157 585
R1282 B.n156 B.n155 585
R1283 B.n154 B.n153 585
R1284 B.n152 B.n151 585
R1285 B.n150 B.n149 585
R1286 B.n148 B.n147 585
R1287 B.n146 B.n145 585
R1288 B.n144 B.n143 585
R1289 B.n142 B.n141 585
R1290 B.n140 B.n139 585
R1291 B.n138 B.n137 585
R1292 B.n136 B.n135 585
R1293 B.n134 B.n133 585
R1294 B.n132 B.n131 585
R1295 B.n130 B.n129 585
R1296 B.n128 B.n127 585
R1297 B.n126 B.n125 585
R1298 B.n124 B.n123 585
R1299 B.n53 B.n52 585
R1300 B.n860 B.n54 585
R1301 B.n864 B.n54 585
R1302 B.n859 B.n858 585
R1303 B.n858 B.n50 585
R1304 B.n857 B.n49 585
R1305 B.n870 B.n49 585
R1306 B.n856 B.n48 585
R1307 B.n871 B.n48 585
R1308 B.n855 B.n47 585
R1309 B.n872 B.n47 585
R1310 B.n854 B.n853 585
R1311 B.n853 B.n43 585
R1312 B.n852 B.n42 585
R1313 B.n878 B.n42 585
R1314 B.n851 B.n41 585
R1315 B.n879 B.n41 585
R1316 B.n850 B.n40 585
R1317 B.n880 B.n40 585
R1318 B.n849 B.n848 585
R1319 B.n848 B.n36 585
R1320 B.n847 B.n35 585
R1321 B.n886 B.n35 585
R1322 B.n846 B.n34 585
R1323 B.n887 B.n34 585
R1324 B.n845 B.n33 585
R1325 B.n888 B.n33 585
R1326 B.n844 B.n843 585
R1327 B.n843 B.n29 585
R1328 B.n842 B.n28 585
R1329 B.n894 B.n28 585
R1330 B.n841 B.n27 585
R1331 B.n895 B.n27 585
R1332 B.n840 B.n26 585
R1333 B.n896 B.n26 585
R1334 B.n839 B.n838 585
R1335 B.n838 B.n22 585
R1336 B.n837 B.n21 585
R1337 B.n902 B.n21 585
R1338 B.n836 B.n20 585
R1339 B.n903 B.n20 585
R1340 B.n835 B.n19 585
R1341 B.n904 B.n19 585
R1342 B.n834 B.n833 585
R1343 B.n833 B.n15 585
R1344 B.n832 B.n14 585
R1345 B.n910 B.n14 585
R1346 B.n831 B.n13 585
R1347 B.n911 B.n13 585
R1348 B.n830 B.n12 585
R1349 B.n912 B.n12 585
R1350 B.n829 B.n828 585
R1351 B.n828 B.n8 585
R1352 B.n827 B.n7 585
R1353 B.n918 B.n7 585
R1354 B.n826 B.n6 585
R1355 B.n919 B.n6 585
R1356 B.n825 B.n5 585
R1357 B.n920 B.n5 585
R1358 B.n824 B.n823 585
R1359 B.n823 B.n4 585
R1360 B.n822 B.n369 585
R1361 B.n822 B.n821 585
R1362 B.n812 B.n370 585
R1363 B.n371 B.n370 585
R1364 B.n814 B.n813 585
R1365 B.n815 B.n814 585
R1366 B.n811 B.n375 585
R1367 B.n379 B.n375 585
R1368 B.n810 B.n809 585
R1369 B.n809 B.n808 585
R1370 B.n377 B.n376 585
R1371 B.n378 B.n377 585
R1372 B.n801 B.n800 585
R1373 B.n802 B.n801 585
R1374 B.n799 B.n384 585
R1375 B.n384 B.n383 585
R1376 B.n798 B.n797 585
R1377 B.n797 B.n796 585
R1378 B.n386 B.n385 585
R1379 B.n387 B.n386 585
R1380 B.n789 B.n788 585
R1381 B.n790 B.n789 585
R1382 B.n787 B.n392 585
R1383 B.n392 B.n391 585
R1384 B.n786 B.n785 585
R1385 B.n785 B.n784 585
R1386 B.n394 B.n393 585
R1387 B.n395 B.n394 585
R1388 B.n777 B.n776 585
R1389 B.n778 B.n777 585
R1390 B.n775 B.n400 585
R1391 B.n400 B.n399 585
R1392 B.n774 B.n773 585
R1393 B.n773 B.n772 585
R1394 B.n402 B.n401 585
R1395 B.n403 B.n402 585
R1396 B.n765 B.n764 585
R1397 B.n766 B.n765 585
R1398 B.n763 B.n408 585
R1399 B.n408 B.n407 585
R1400 B.n762 B.n761 585
R1401 B.n761 B.n760 585
R1402 B.n410 B.n409 585
R1403 B.n411 B.n410 585
R1404 B.n753 B.n752 585
R1405 B.n754 B.n753 585
R1406 B.n751 B.n416 585
R1407 B.n416 B.n415 585
R1408 B.n750 B.n749 585
R1409 B.n749 B.n748 585
R1410 B.n418 B.n417 585
R1411 B.n419 B.n418 585
R1412 B.n741 B.n740 585
R1413 B.n742 B.n741 585
R1414 B.n422 B.n421 585
R1415 B.n491 B.n489 585
R1416 B.n492 B.n488 585
R1417 B.n492 B.n423 585
R1418 B.n495 B.n494 585
R1419 B.n496 B.n487 585
R1420 B.n498 B.n497 585
R1421 B.n500 B.n486 585
R1422 B.n503 B.n502 585
R1423 B.n504 B.n485 585
R1424 B.n506 B.n505 585
R1425 B.n508 B.n484 585
R1426 B.n511 B.n510 585
R1427 B.n512 B.n483 585
R1428 B.n514 B.n513 585
R1429 B.n516 B.n482 585
R1430 B.n519 B.n518 585
R1431 B.n520 B.n481 585
R1432 B.n522 B.n521 585
R1433 B.n524 B.n480 585
R1434 B.n527 B.n526 585
R1435 B.n528 B.n479 585
R1436 B.n530 B.n529 585
R1437 B.n532 B.n478 585
R1438 B.n535 B.n534 585
R1439 B.n536 B.n477 585
R1440 B.n538 B.n537 585
R1441 B.n540 B.n476 585
R1442 B.n543 B.n542 585
R1443 B.n544 B.n475 585
R1444 B.n546 B.n545 585
R1445 B.n548 B.n474 585
R1446 B.n551 B.n550 585
R1447 B.n552 B.n473 585
R1448 B.n554 B.n553 585
R1449 B.n556 B.n472 585
R1450 B.n559 B.n558 585
R1451 B.n560 B.n471 585
R1452 B.n562 B.n561 585
R1453 B.n564 B.n470 585
R1454 B.n567 B.n566 585
R1455 B.n568 B.n469 585
R1456 B.n570 B.n569 585
R1457 B.n572 B.n468 585
R1458 B.n575 B.n574 585
R1459 B.n576 B.n467 585
R1460 B.n578 B.n577 585
R1461 B.n580 B.n466 585
R1462 B.n583 B.n582 585
R1463 B.n584 B.n465 585
R1464 B.n586 B.n585 585
R1465 B.n588 B.n464 585
R1466 B.n591 B.n590 585
R1467 B.n592 B.n463 585
R1468 B.n594 B.n593 585
R1469 B.n596 B.n462 585
R1470 B.n599 B.n598 585
R1471 B.n600 B.n461 585
R1472 B.n605 B.n604 585
R1473 B.n607 B.n460 585
R1474 B.n610 B.n609 585
R1475 B.n611 B.n459 585
R1476 B.n613 B.n612 585
R1477 B.n615 B.n458 585
R1478 B.n618 B.n617 585
R1479 B.n619 B.n457 585
R1480 B.n621 B.n620 585
R1481 B.n623 B.n456 585
R1482 B.n626 B.n625 585
R1483 B.n627 B.n452 585
R1484 B.n629 B.n628 585
R1485 B.n631 B.n451 585
R1486 B.n634 B.n633 585
R1487 B.n635 B.n450 585
R1488 B.n637 B.n636 585
R1489 B.n639 B.n449 585
R1490 B.n642 B.n641 585
R1491 B.n643 B.n448 585
R1492 B.n645 B.n644 585
R1493 B.n647 B.n447 585
R1494 B.n650 B.n649 585
R1495 B.n651 B.n446 585
R1496 B.n653 B.n652 585
R1497 B.n655 B.n445 585
R1498 B.n658 B.n657 585
R1499 B.n659 B.n444 585
R1500 B.n661 B.n660 585
R1501 B.n663 B.n443 585
R1502 B.n666 B.n665 585
R1503 B.n667 B.n442 585
R1504 B.n669 B.n668 585
R1505 B.n671 B.n441 585
R1506 B.n674 B.n673 585
R1507 B.n675 B.n440 585
R1508 B.n677 B.n676 585
R1509 B.n679 B.n439 585
R1510 B.n682 B.n681 585
R1511 B.n683 B.n438 585
R1512 B.n685 B.n684 585
R1513 B.n687 B.n437 585
R1514 B.n690 B.n689 585
R1515 B.n691 B.n436 585
R1516 B.n693 B.n692 585
R1517 B.n695 B.n435 585
R1518 B.n698 B.n697 585
R1519 B.n699 B.n434 585
R1520 B.n701 B.n700 585
R1521 B.n703 B.n433 585
R1522 B.n706 B.n705 585
R1523 B.n707 B.n432 585
R1524 B.n709 B.n708 585
R1525 B.n711 B.n431 585
R1526 B.n714 B.n713 585
R1527 B.n715 B.n430 585
R1528 B.n717 B.n716 585
R1529 B.n719 B.n429 585
R1530 B.n722 B.n721 585
R1531 B.n723 B.n428 585
R1532 B.n725 B.n724 585
R1533 B.n727 B.n427 585
R1534 B.n730 B.n729 585
R1535 B.n731 B.n426 585
R1536 B.n733 B.n732 585
R1537 B.n735 B.n425 585
R1538 B.n738 B.n737 585
R1539 B.n739 B.n424 585
R1540 B.n744 B.n743 585
R1541 B.n743 B.n742 585
R1542 B.n745 B.n420 585
R1543 B.n420 B.n419 585
R1544 B.n747 B.n746 585
R1545 B.n748 B.n747 585
R1546 B.n414 B.n413 585
R1547 B.n415 B.n414 585
R1548 B.n756 B.n755 585
R1549 B.n755 B.n754 585
R1550 B.n757 B.n412 585
R1551 B.n412 B.n411 585
R1552 B.n759 B.n758 585
R1553 B.n760 B.n759 585
R1554 B.n406 B.n405 585
R1555 B.n407 B.n406 585
R1556 B.n768 B.n767 585
R1557 B.n767 B.n766 585
R1558 B.n769 B.n404 585
R1559 B.n404 B.n403 585
R1560 B.n771 B.n770 585
R1561 B.n772 B.n771 585
R1562 B.n398 B.n397 585
R1563 B.n399 B.n398 585
R1564 B.n780 B.n779 585
R1565 B.n779 B.n778 585
R1566 B.n781 B.n396 585
R1567 B.n396 B.n395 585
R1568 B.n783 B.n782 585
R1569 B.n784 B.n783 585
R1570 B.n390 B.n389 585
R1571 B.n391 B.n390 585
R1572 B.n792 B.n791 585
R1573 B.n791 B.n790 585
R1574 B.n793 B.n388 585
R1575 B.n388 B.n387 585
R1576 B.n795 B.n794 585
R1577 B.n796 B.n795 585
R1578 B.n382 B.n381 585
R1579 B.n383 B.n382 585
R1580 B.n804 B.n803 585
R1581 B.n803 B.n802 585
R1582 B.n805 B.n380 585
R1583 B.n380 B.n378 585
R1584 B.n807 B.n806 585
R1585 B.n808 B.n807 585
R1586 B.n374 B.n373 585
R1587 B.n379 B.n374 585
R1588 B.n817 B.n816 585
R1589 B.n816 B.n815 585
R1590 B.n818 B.n372 585
R1591 B.n372 B.n371 585
R1592 B.n820 B.n819 585
R1593 B.n821 B.n820 585
R1594 B.n2 B.n0 585
R1595 B.n4 B.n2 585
R1596 B.n3 B.n1 585
R1597 B.n919 B.n3 585
R1598 B.n917 B.n916 585
R1599 B.n918 B.n917 585
R1600 B.n915 B.n9 585
R1601 B.n9 B.n8 585
R1602 B.n914 B.n913 585
R1603 B.n913 B.n912 585
R1604 B.n11 B.n10 585
R1605 B.n911 B.n11 585
R1606 B.n909 B.n908 585
R1607 B.n910 B.n909 585
R1608 B.n907 B.n16 585
R1609 B.n16 B.n15 585
R1610 B.n906 B.n905 585
R1611 B.n905 B.n904 585
R1612 B.n18 B.n17 585
R1613 B.n903 B.n18 585
R1614 B.n901 B.n900 585
R1615 B.n902 B.n901 585
R1616 B.n899 B.n23 585
R1617 B.n23 B.n22 585
R1618 B.n898 B.n897 585
R1619 B.n897 B.n896 585
R1620 B.n25 B.n24 585
R1621 B.n895 B.n25 585
R1622 B.n893 B.n892 585
R1623 B.n894 B.n893 585
R1624 B.n891 B.n30 585
R1625 B.n30 B.n29 585
R1626 B.n890 B.n889 585
R1627 B.n889 B.n888 585
R1628 B.n32 B.n31 585
R1629 B.n887 B.n32 585
R1630 B.n885 B.n884 585
R1631 B.n886 B.n885 585
R1632 B.n883 B.n37 585
R1633 B.n37 B.n36 585
R1634 B.n882 B.n881 585
R1635 B.n881 B.n880 585
R1636 B.n39 B.n38 585
R1637 B.n879 B.n39 585
R1638 B.n877 B.n876 585
R1639 B.n878 B.n877 585
R1640 B.n875 B.n44 585
R1641 B.n44 B.n43 585
R1642 B.n874 B.n873 585
R1643 B.n873 B.n872 585
R1644 B.n46 B.n45 585
R1645 B.n871 B.n46 585
R1646 B.n869 B.n868 585
R1647 B.n870 B.n869 585
R1648 B.n867 B.n51 585
R1649 B.n51 B.n50 585
R1650 B.n866 B.n865 585
R1651 B.n865 B.n864 585
R1652 B.n922 B.n921 585
R1653 B.n921 B.n920 585
R1654 B.n743 B.n422 487.695
R1655 B.n865 B.n53 487.695
R1656 B.n741 B.n424 487.695
R1657 B.n862 B.n54 487.695
R1658 B.n453 B.t8 422.928
R1659 B.n601 B.t4 422.928
R1660 B.n120 B.t15 422.928
R1661 B.n118 B.t11 422.928
R1662 B.n453 B.t10 418.955
R1663 B.n601 B.t7 418.955
R1664 B.n120 B.t16 418.955
R1665 B.n118 B.t13 418.955
R1666 B.n454 B.t9 374.932
R1667 B.n119 B.t14 374.932
R1668 B.n602 B.t6 374.932
R1669 B.n121 B.t17 374.932
R1670 B.n863 B.n116 256.663
R1671 B.n863 B.n115 256.663
R1672 B.n863 B.n114 256.663
R1673 B.n863 B.n113 256.663
R1674 B.n863 B.n112 256.663
R1675 B.n863 B.n111 256.663
R1676 B.n863 B.n110 256.663
R1677 B.n863 B.n109 256.663
R1678 B.n863 B.n108 256.663
R1679 B.n863 B.n107 256.663
R1680 B.n863 B.n106 256.663
R1681 B.n863 B.n105 256.663
R1682 B.n863 B.n104 256.663
R1683 B.n863 B.n103 256.663
R1684 B.n863 B.n102 256.663
R1685 B.n863 B.n101 256.663
R1686 B.n863 B.n100 256.663
R1687 B.n863 B.n99 256.663
R1688 B.n863 B.n98 256.663
R1689 B.n863 B.n97 256.663
R1690 B.n863 B.n96 256.663
R1691 B.n863 B.n95 256.663
R1692 B.n863 B.n94 256.663
R1693 B.n863 B.n93 256.663
R1694 B.n863 B.n92 256.663
R1695 B.n863 B.n91 256.663
R1696 B.n863 B.n90 256.663
R1697 B.n863 B.n89 256.663
R1698 B.n863 B.n88 256.663
R1699 B.n863 B.n87 256.663
R1700 B.n863 B.n86 256.663
R1701 B.n863 B.n85 256.663
R1702 B.n863 B.n84 256.663
R1703 B.n863 B.n83 256.663
R1704 B.n863 B.n82 256.663
R1705 B.n863 B.n81 256.663
R1706 B.n863 B.n80 256.663
R1707 B.n863 B.n79 256.663
R1708 B.n863 B.n78 256.663
R1709 B.n863 B.n77 256.663
R1710 B.n863 B.n76 256.663
R1711 B.n863 B.n75 256.663
R1712 B.n863 B.n74 256.663
R1713 B.n863 B.n73 256.663
R1714 B.n863 B.n72 256.663
R1715 B.n863 B.n71 256.663
R1716 B.n863 B.n70 256.663
R1717 B.n863 B.n69 256.663
R1718 B.n863 B.n68 256.663
R1719 B.n863 B.n67 256.663
R1720 B.n863 B.n66 256.663
R1721 B.n863 B.n65 256.663
R1722 B.n863 B.n64 256.663
R1723 B.n863 B.n63 256.663
R1724 B.n863 B.n62 256.663
R1725 B.n863 B.n61 256.663
R1726 B.n863 B.n60 256.663
R1727 B.n863 B.n59 256.663
R1728 B.n863 B.n58 256.663
R1729 B.n863 B.n57 256.663
R1730 B.n863 B.n56 256.663
R1731 B.n863 B.n55 256.663
R1732 B.n490 B.n423 256.663
R1733 B.n493 B.n423 256.663
R1734 B.n499 B.n423 256.663
R1735 B.n501 B.n423 256.663
R1736 B.n507 B.n423 256.663
R1737 B.n509 B.n423 256.663
R1738 B.n515 B.n423 256.663
R1739 B.n517 B.n423 256.663
R1740 B.n523 B.n423 256.663
R1741 B.n525 B.n423 256.663
R1742 B.n531 B.n423 256.663
R1743 B.n533 B.n423 256.663
R1744 B.n539 B.n423 256.663
R1745 B.n541 B.n423 256.663
R1746 B.n547 B.n423 256.663
R1747 B.n549 B.n423 256.663
R1748 B.n555 B.n423 256.663
R1749 B.n557 B.n423 256.663
R1750 B.n563 B.n423 256.663
R1751 B.n565 B.n423 256.663
R1752 B.n571 B.n423 256.663
R1753 B.n573 B.n423 256.663
R1754 B.n579 B.n423 256.663
R1755 B.n581 B.n423 256.663
R1756 B.n587 B.n423 256.663
R1757 B.n589 B.n423 256.663
R1758 B.n595 B.n423 256.663
R1759 B.n597 B.n423 256.663
R1760 B.n606 B.n423 256.663
R1761 B.n608 B.n423 256.663
R1762 B.n614 B.n423 256.663
R1763 B.n616 B.n423 256.663
R1764 B.n622 B.n423 256.663
R1765 B.n624 B.n423 256.663
R1766 B.n630 B.n423 256.663
R1767 B.n632 B.n423 256.663
R1768 B.n638 B.n423 256.663
R1769 B.n640 B.n423 256.663
R1770 B.n646 B.n423 256.663
R1771 B.n648 B.n423 256.663
R1772 B.n654 B.n423 256.663
R1773 B.n656 B.n423 256.663
R1774 B.n662 B.n423 256.663
R1775 B.n664 B.n423 256.663
R1776 B.n670 B.n423 256.663
R1777 B.n672 B.n423 256.663
R1778 B.n678 B.n423 256.663
R1779 B.n680 B.n423 256.663
R1780 B.n686 B.n423 256.663
R1781 B.n688 B.n423 256.663
R1782 B.n694 B.n423 256.663
R1783 B.n696 B.n423 256.663
R1784 B.n702 B.n423 256.663
R1785 B.n704 B.n423 256.663
R1786 B.n710 B.n423 256.663
R1787 B.n712 B.n423 256.663
R1788 B.n718 B.n423 256.663
R1789 B.n720 B.n423 256.663
R1790 B.n726 B.n423 256.663
R1791 B.n728 B.n423 256.663
R1792 B.n734 B.n423 256.663
R1793 B.n736 B.n423 256.663
R1794 B.n743 B.n420 163.367
R1795 B.n747 B.n420 163.367
R1796 B.n747 B.n414 163.367
R1797 B.n755 B.n414 163.367
R1798 B.n755 B.n412 163.367
R1799 B.n759 B.n412 163.367
R1800 B.n759 B.n406 163.367
R1801 B.n767 B.n406 163.367
R1802 B.n767 B.n404 163.367
R1803 B.n771 B.n404 163.367
R1804 B.n771 B.n398 163.367
R1805 B.n779 B.n398 163.367
R1806 B.n779 B.n396 163.367
R1807 B.n783 B.n396 163.367
R1808 B.n783 B.n390 163.367
R1809 B.n791 B.n390 163.367
R1810 B.n791 B.n388 163.367
R1811 B.n795 B.n388 163.367
R1812 B.n795 B.n382 163.367
R1813 B.n803 B.n382 163.367
R1814 B.n803 B.n380 163.367
R1815 B.n807 B.n380 163.367
R1816 B.n807 B.n374 163.367
R1817 B.n816 B.n374 163.367
R1818 B.n816 B.n372 163.367
R1819 B.n820 B.n372 163.367
R1820 B.n820 B.n2 163.367
R1821 B.n921 B.n2 163.367
R1822 B.n921 B.n3 163.367
R1823 B.n917 B.n3 163.367
R1824 B.n917 B.n9 163.367
R1825 B.n913 B.n9 163.367
R1826 B.n913 B.n11 163.367
R1827 B.n909 B.n11 163.367
R1828 B.n909 B.n16 163.367
R1829 B.n905 B.n16 163.367
R1830 B.n905 B.n18 163.367
R1831 B.n901 B.n18 163.367
R1832 B.n901 B.n23 163.367
R1833 B.n897 B.n23 163.367
R1834 B.n897 B.n25 163.367
R1835 B.n893 B.n25 163.367
R1836 B.n893 B.n30 163.367
R1837 B.n889 B.n30 163.367
R1838 B.n889 B.n32 163.367
R1839 B.n885 B.n32 163.367
R1840 B.n885 B.n37 163.367
R1841 B.n881 B.n37 163.367
R1842 B.n881 B.n39 163.367
R1843 B.n877 B.n39 163.367
R1844 B.n877 B.n44 163.367
R1845 B.n873 B.n44 163.367
R1846 B.n873 B.n46 163.367
R1847 B.n869 B.n46 163.367
R1848 B.n869 B.n51 163.367
R1849 B.n865 B.n51 163.367
R1850 B.n492 B.n491 163.367
R1851 B.n494 B.n492 163.367
R1852 B.n498 B.n487 163.367
R1853 B.n502 B.n500 163.367
R1854 B.n506 B.n485 163.367
R1855 B.n510 B.n508 163.367
R1856 B.n514 B.n483 163.367
R1857 B.n518 B.n516 163.367
R1858 B.n522 B.n481 163.367
R1859 B.n526 B.n524 163.367
R1860 B.n530 B.n479 163.367
R1861 B.n534 B.n532 163.367
R1862 B.n538 B.n477 163.367
R1863 B.n542 B.n540 163.367
R1864 B.n546 B.n475 163.367
R1865 B.n550 B.n548 163.367
R1866 B.n554 B.n473 163.367
R1867 B.n558 B.n556 163.367
R1868 B.n562 B.n471 163.367
R1869 B.n566 B.n564 163.367
R1870 B.n570 B.n469 163.367
R1871 B.n574 B.n572 163.367
R1872 B.n578 B.n467 163.367
R1873 B.n582 B.n580 163.367
R1874 B.n586 B.n465 163.367
R1875 B.n590 B.n588 163.367
R1876 B.n594 B.n463 163.367
R1877 B.n598 B.n596 163.367
R1878 B.n605 B.n461 163.367
R1879 B.n609 B.n607 163.367
R1880 B.n613 B.n459 163.367
R1881 B.n617 B.n615 163.367
R1882 B.n621 B.n457 163.367
R1883 B.n625 B.n623 163.367
R1884 B.n629 B.n452 163.367
R1885 B.n633 B.n631 163.367
R1886 B.n637 B.n450 163.367
R1887 B.n641 B.n639 163.367
R1888 B.n645 B.n448 163.367
R1889 B.n649 B.n647 163.367
R1890 B.n653 B.n446 163.367
R1891 B.n657 B.n655 163.367
R1892 B.n661 B.n444 163.367
R1893 B.n665 B.n663 163.367
R1894 B.n669 B.n442 163.367
R1895 B.n673 B.n671 163.367
R1896 B.n677 B.n440 163.367
R1897 B.n681 B.n679 163.367
R1898 B.n685 B.n438 163.367
R1899 B.n689 B.n687 163.367
R1900 B.n693 B.n436 163.367
R1901 B.n697 B.n695 163.367
R1902 B.n701 B.n434 163.367
R1903 B.n705 B.n703 163.367
R1904 B.n709 B.n432 163.367
R1905 B.n713 B.n711 163.367
R1906 B.n717 B.n430 163.367
R1907 B.n721 B.n719 163.367
R1908 B.n725 B.n428 163.367
R1909 B.n729 B.n727 163.367
R1910 B.n733 B.n426 163.367
R1911 B.n737 B.n735 163.367
R1912 B.n741 B.n418 163.367
R1913 B.n749 B.n418 163.367
R1914 B.n749 B.n416 163.367
R1915 B.n753 B.n416 163.367
R1916 B.n753 B.n410 163.367
R1917 B.n761 B.n410 163.367
R1918 B.n761 B.n408 163.367
R1919 B.n765 B.n408 163.367
R1920 B.n765 B.n402 163.367
R1921 B.n773 B.n402 163.367
R1922 B.n773 B.n400 163.367
R1923 B.n777 B.n400 163.367
R1924 B.n777 B.n394 163.367
R1925 B.n785 B.n394 163.367
R1926 B.n785 B.n392 163.367
R1927 B.n789 B.n392 163.367
R1928 B.n789 B.n386 163.367
R1929 B.n797 B.n386 163.367
R1930 B.n797 B.n384 163.367
R1931 B.n801 B.n384 163.367
R1932 B.n801 B.n377 163.367
R1933 B.n809 B.n377 163.367
R1934 B.n809 B.n375 163.367
R1935 B.n814 B.n375 163.367
R1936 B.n814 B.n370 163.367
R1937 B.n822 B.n370 163.367
R1938 B.n823 B.n822 163.367
R1939 B.n823 B.n5 163.367
R1940 B.n6 B.n5 163.367
R1941 B.n7 B.n6 163.367
R1942 B.n828 B.n7 163.367
R1943 B.n828 B.n12 163.367
R1944 B.n13 B.n12 163.367
R1945 B.n14 B.n13 163.367
R1946 B.n833 B.n14 163.367
R1947 B.n833 B.n19 163.367
R1948 B.n20 B.n19 163.367
R1949 B.n21 B.n20 163.367
R1950 B.n838 B.n21 163.367
R1951 B.n838 B.n26 163.367
R1952 B.n27 B.n26 163.367
R1953 B.n28 B.n27 163.367
R1954 B.n843 B.n28 163.367
R1955 B.n843 B.n33 163.367
R1956 B.n34 B.n33 163.367
R1957 B.n35 B.n34 163.367
R1958 B.n848 B.n35 163.367
R1959 B.n848 B.n40 163.367
R1960 B.n41 B.n40 163.367
R1961 B.n42 B.n41 163.367
R1962 B.n853 B.n42 163.367
R1963 B.n853 B.n47 163.367
R1964 B.n48 B.n47 163.367
R1965 B.n49 B.n48 163.367
R1966 B.n858 B.n49 163.367
R1967 B.n858 B.n54 163.367
R1968 B.n125 B.n124 163.367
R1969 B.n129 B.n128 163.367
R1970 B.n133 B.n132 163.367
R1971 B.n137 B.n136 163.367
R1972 B.n141 B.n140 163.367
R1973 B.n145 B.n144 163.367
R1974 B.n149 B.n148 163.367
R1975 B.n153 B.n152 163.367
R1976 B.n157 B.n156 163.367
R1977 B.n161 B.n160 163.367
R1978 B.n165 B.n164 163.367
R1979 B.n169 B.n168 163.367
R1980 B.n173 B.n172 163.367
R1981 B.n177 B.n176 163.367
R1982 B.n181 B.n180 163.367
R1983 B.n185 B.n184 163.367
R1984 B.n189 B.n188 163.367
R1985 B.n193 B.n192 163.367
R1986 B.n197 B.n196 163.367
R1987 B.n201 B.n200 163.367
R1988 B.n205 B.n204 163.367
R1989 B.n209 B.n208 163.367
R1990 B.n213 B.n212 163.367
R1991 B.n217 B.n216 163.367
R1992 B.n221 B.n220 163.367
R1993 B.n225 B.n224 163.367
R1994 B.n229 B.n228 163.367
R1995 B.n233 B.n232 163.367
R1996 B.n237 B.n236 163.367
R1997 B.n241 B.n240 163.367
R1998 B.n245 B.n244 163.367
R1999 B.n249 B.n248 163.367
R2000 B.n253 B.n252 163.367
R2001 B.n258 B.n257 163.367
R2002 B.n262 B.n261 163.367
R2003 B.n266 B.n265 163.367
R2004 B.n270 B.n269 163.367
R2005 B.n274 B.n273 163.367
R2006 B.n278 B.n277 163.367
R2007 B.n282 B.n281 163.367
R2008 B.n286 B.n285 163.367
R2009 B.n290 B.n289 163.367
R2010 B.n294 B.n293 163.367
R2011 B.n298 B.n297 163.367
R2012 B.n302 B.n301 163.367
R2013 B.n306 B.n305 163.367
R2014 B.n310 B.n309 163.367
R2015 B.n314 B.n313 163.367
R2016 B.n318 B.n317 163.367
R2017 B.n322 B.n321 163.367
R2018 B.n326 B.n325 163.367
R2019 B.n330 B.n329 163.367
R2020 B.n334 B.n333 163.367
R2021 B.n338 B.n337 163.367
R2022 B.n342 B.n341 163.367
R2023 B.n346 B.n345 163.367
R2024 B.n350 B.n349 163.367
R2025 B.n354 B.n353 163.367
R2026 B.n358 B.n357 163.367
R2027 B.n362 B.n361 163.367
R2028 B.n366 B.n365 163.367
R2029 B.n862 B.n117 163.367
R2030 B.n490 B.n422 71.676
R2031 B.n494 B.n493 71.676
R2032 B.n499 B.n498 71.676
R2033 B.n502 B.n501 71.676
R2034 B.n507 B.n506 71.676
R2035 B.n510 B.n509 71.676
R2036 B.n515 B.n514 71.676
R2037 B.n518 B.n517 71.676
R2038 B.n523 B.n522 71.676
R2039 B.n526 B.n525 71.676
R2040 B.n531 B.n530 71.676
R2041 B.n534 B.n533 71.676
R2042 B.n539 B.n538 71.676
R2043 B.n542 B.n541 71.676
R2044 B.n547 B.n546 71.676
R2045 B.n550 B.n549 71.676
R2046 B.n555 B.n554 71.676
R2047 B.n558 B.n557 71.676
R2048 B.n563 B.n562 71.676
R2049 B.n566 B.n565 71.676
R2050 B.n571 B.n570 71.676
R2051 B.n574 B.n573 71.676
R2052 B.n579 B.n578 71.676
R2053 B.n582 B.n581 71.676
R2054 B.n587 B.n586 71.676
R2055 B.n590 B.n589 71.676
R2056 B.n595 B.n594 71.676
R2057 B.n598 B.n597 71.676
R2058 B.n606 B.n605 71.676
R2059 B.n609 B.n608 71.676
R2060 B.n614 B.n613 71.676
R2061 B.n617 B.n616 71.676
R2062 B.n622 B.n621 71.676
R2063 B.n625 B.n624 71.676
R2064 B.n630 B.n629 71.676
R2065 B.n633 B.n632 71.676
R2066 B.n638 B.n637 71.676
R2067 B.n641 B.n640 71.676
R2068 B.n646 B.n645 71.676
R2069 B.n649 B.n648 71.676
R2070 B.n654 B.n653 71.676
R2071 B.n657 B.n656 71.676
R2072 B.n662 B.n661 71.676
R2073 B.n665 B.n664 71.676
R2074 B.n670 B.n669 71.676
R2075 B.n673 B.n672 71.676
R2076 B.n678 B.n677 71.676
R2077 B.n681 B.n680 71.676
R2078 B.n686 B.n685 71.676
R2079 B.n689 B.n688 71.676
R2080 B.n694 B.n693 71.676
R2081 B.n697 B.n696 71.676
R2082 B.n702 B.n701 71.676
R2083 B.n705 B.n704 71.676
R2084 B.n710 B.n709 71.676
R2085 B.n713 B.n712 71.676
R2086 B.n718 B.n717 71.676
R2087 B.n721 B.n720 71.676
R2088 B.n726 B.n725 71.676
R2089 B.n729 B.n728 71.676
R2090 B.n734 B.n733 71.676
R2091 B.n737 B.n736 71.676
R2092 B.n55 B.n53 71.676
R2093 B.n125 B.n56 71.676
R2094 B.n129 B.n57 71.676
R2095 B.n133 B.n58 71.676
R2096 B.n137 B.n59 71.676
R2097 B.n141 B.n60 71.676
R2098 B.n145 B.n61 71.676
R2099 B.n149 B.n62 71.676
R2100 B.n153 B.n63 71.676
R2101 B.n157 B.n64 71.676
R2102 B.n161 B.n65 71.676
R2103 B.n165 B.n66 71.676
R2104 B.n169 B.n67 71.676
R2105 B.n173 B.n68 71.676
R2106 B.n177 B.n69 71.676
R2107 B.n181 B.n70 71.676
R2108 B.n185 B.n71 71.676
R2109 B.n189 B.n72 71.676
R2110 B.n193 B.n73 71.676
R2111 B.n197 B.n74 71.676
R2112 B.n201 B.n75 71.676
R2113 B.n205 B.n76 71.676
R2114 B.n209 B.n77 71.676
R2115 B.n213 B.n78 71.676
R2116 B.n217 B.n79 71.676
R2117 B.n221 B.n80 71.676
R2118 B.n225 B.n81 71.676
R2119 B.n229 B.n82 71.676
R2120 B.n233 B.n83 71.676
R2121 B.n237 B.n84 71.676
R2122 B.n241 B.n85 71.676
R2123 B.n245 B.n86 71.676
R2124 B.n249 B.n87 71.676
R2125 B.n253 B.n88 71.676
R2126 B.n258 B.n89 71.676
R2127 B.n262 B.n90 71.676
R2128 B.n266 B.n91 71.676
R2129 B.n270 B.n92 71.676
R2130 B.n274 B.n93 71.676
R2131 B.n278 B.n94 71.676
R2132 B.n282 B.n95 71.676
R2133 B.n286 B.n96 71.676
R2134 B.n290 B.n97 71.676
R2135 B.n294 B.n98 71.676
R2136 B.n298 B.n99 71.676
R2137 B.n302 B.n100 71.676
R2138 B.n306 B.n101 71.676
R2139 B.n310 B.n102 71.676
R2140 B.n314 B.n103 71.676
R2141 B.n318 B.n104 71.676
R2142 B.n322 B.n105 71.676
R2143 B.n326 B.n106 71.676
R2144 B.n330 B.n107 71.676
R2145 B.n334 B.n108 71.676
R2146 B.n338 B.n109 71.676
R2147 B.n342 B.n110 71.676
R2148 B.n346 B.n111 71.676
R2149 B.n350 B.n112 71.676
R2150 B.n354 B.n113 71.676
R2151 B.n358 B.n114 71.676
R2152 B.n362 B.n115 71.676
R2153 B.n366 B.n116 71.676
R2154 B.n117 B.n116 71.676
R2155 B.n365 B.n115 71.676
R2156 B.n361 B.n114 71.676
R2157 B.n357 B.n113 71.676
R2158 B.n353 B.n112 71.676
R2159 B.n349 B.n111 71.676
R2160 B.n345 B.n110 71.676
R2161 B.n341 B.n109 71.676
R2162 B.n337 B.n108 71.676
R2163 B.n333 B.n107 71.676
R2164 B.n329 B.n106 71.676
R2165 B.n325 B.n105 71.676
R2166 B.n321 B.n104 71.676
R2167 B.n317 B.n103 71.676
R2168 B.n313 B.n102 71.676
R2169 B.n309 B.n101 71.676
R2170 B.n305 B.n100 71.676
R2171 B.n301 B.n99 71.676
R2172 B.n297 B.n98 71.676
R2173 B.n293 B.n97 71.676
R2174 B.n289 B.n96 71.676
R2175 B.n285 B.n95 71.676
R2176 B.n281 B.n94 71.676
R2177 B.n277 B.n93 71.676
R2178 B.n273 B.n92 71.676
R2179 B.n269 B.n91 71.676
R2180 B.n265 B.n90 71.676
R2181 B.n261 B.n89 71.676
R2182 B.n257 B.n88 71.676
R2183 B.n252 B.n87 71.676
R2184 B.n248 B.n86 71.676
R2185 B.n244 B.n85 71.676
R2186 B.n240 B.n84 71.676
R2187 B.n236 B.n83 71.676
R2188 B.n232 B.n82 71.676
R2189 B.n228 B.n81 71.676
R2190 B.n224 B.n80 71.676
R2191 B.n220 B.n79 71.676
R2192 B.n216 B.n78 71.676
R2193 B.n212 B.n77 71.676
R2194 B.n208 B.n76 71.676
R2195 B.n204 B.n75 71.676
R2196 B.n200 B.n74 71.676
R2197 B.n196 B.n73 71.676
R2198 B.n192 B.n72 71.676
R2199 B.n188 B.n71 71.676
R2200 B.n184 B.n70 71.676
R2201 B.n180 B.n69 71.676
R2202 B.n176 B.n68 71.676
R2203 B.n172 B.n67 71.676
R2204 B.n168 B.n66 71.676
R2205 B.n164 B.n65 71.676
R2206 B.n160 B.n64 71.676
R2207 B.n156 B.n63 71.676
R2208 B.n152 B.n62 71.676
R2209 B.n148 B.n61 71.676
R2210 B.n144 B.n60 71.676
R2211 B.n140 B.n59 71.676
R2212 B.n136 B.n58 71.676
R2213 B.n132 B.n57 71.676
R2214 B.n128 B.n56 71.676
R2215 B.n124 B.n55 71.676
R2216 B.n491 B.n490 71.676
R2217 B.n493 B.n487 71.676
R2218 B.n500 B.n499 71.676
R2219 B.n501 B.n485 71.676
R2220 B.n508 B.n507 71.676
R2221 B.n509 B.n483 71.676
R2222 B.n516 B.n515 71.676
R2223 B.n517 B.n481 71.676
R2224 B.n524 B.n523 71.676
R2225 B.n525 B.n479 71.676
R2226 B.n532 B.n531 71.676
R2227 B.n533 B.n477 71.676
R2228 B.n540 B.n539 71.676
R2229 B.n541 B.n475 71.676
R2230 B.n548 B.n547 71.676
R2231 B.n549 B.n473 71.676
R2232 B.n556 B.n555 71.676
R2233 B.n557 B.n471 71.676
R2234 B.n564 B.n563 71.676
R2235 B.n565 B.n469 71.676
R2236 B.n572 B.n571 71.676
R2237 B.n573 B.n467 71.676
R2238 B.n580 B.n579 71.676
R2239 B.n581 B.n465 71.676
R2240 B.n588 B.n587 71.676
R2241 B.n589 B.n463 71.676
R2242 B.n596 B.n595 71.676
R2243 B.n597 B.n461 71.676
R2244 B.n607 B.n606 71.676
R2245 B.n608 B.n459 71.676
R2246 B.n615 B.n614 71.676
R2247 B.n616 B.n457 71.676
R2248 B.n623 B.n622 71.676
R2249 B.n624 B.n452 71.676
R2250 B.n631 B.n630 71.676
R2251 B.n632 B.n450 71.676
R2252 B.n639 B.n638 71.676
R2253 B.n640 B.n448 71.676
R2254 B.n647 B.n646 71.676
R2255 B.n648 B.n446 71.676
R2256 B.n655 B.n654 71.676
R2257 B.n656 B.n444 71.676
R2258 B.n663 B.n662 71.676
R2259 B.n664 B.n442 71.676
R2260 B.n671 B.n670 71.676
R2261 B.n672 B.n440 71.676
R2262 B.n679 B.n678 71.676
R2263 B.n680 B.n438 71.676
R2264 B.n687 B.n686 71.676
R2265 B.n688 B.n436 71.676
R2266 B.n695 B.n694 71.676
R2267 B.n696 B.n434 71.676
R2268 B.n703 B.n702 71.676
R2269 B.n704 B.n432 71.676
R2270 B.n711 B.n710 71.676
R2271 B.n712 B.n430 71.676
R2272 B.n719 B.n718 71.676
R2273 B.n720 B.n428 71.676
R2274 B.n727 B.n726 71.676
R2275 B.n728 B.n426 71.676
R2276 B.n735 B.n734 71.676
R2277 B.n736 B.n424 71.676
R2278 B.n742 B.n423 64.5209
R2279 B.n864 B.n863 64.5209
R2280 B.n455 B.n454 59.5399
R2281 B.n603 B.n602 59.5399
R2282 B.n122 B.n121 59.5399
R2283 B.n255 B.n119 59.5399
R2284 B.n454 B.n453 44.0247
R2285 B.n602 B.n601 44.0247
R2286 B.n121 B.n120 44.0247
R2287 B.n119 B.n118 44.0247
R2288 B.n742 B.n419 32.9884
R2289 B.n748 B.n419 32.9884
R2290 B.n748 B.n415 32.9884
R2291 B.n754 B.n415 32.9884
R2292 B.n754 B.n411 32.9884
R2293 B.n760 B.n411 32.9884
R2294 B.n766 B.n407 32.9884
R2295 B.n766 B.n403 32.9884
R2296 B.n772 B.n403 32.9884
R2297 B.n772 B.n399 32.9884
R2298 B.n778 B.n399 32.9884
R2299 B.n778 B.n395 32.9884
R2300 B.n784 B.n395 32.9884
R2301 B.n784 B.n391 32.9884
R2302 B.n790 B.n391 32.9884
R2303 B.n796 B.n387 32.9884
R2304 B.n796 B.n383 32.9884
R2305 B.n802 B.n383 32.9884
R2306 B.n802 B.n378 32.9884
R2307 B.n808 B.n378 32.9884
R2308 B.n808 B.n379 32.9884
R2309 B.n815 B.n371 32.9884
R2310 B.n821 B.n371 32.9884
R2311 B.n821 B.n4 32.9884
R2312 B.n920 B.n4 32.9884
R2313 B.n920 B.n919 32.9884
R2314 B.n919 B.n918 32.9884
R2315 B.n918 B.n8 32.9884
R2316 B.n912 B.n8 32.9884
R2317 B.n911 B.n910 32.9884
R2318 B.n910 B.n15 32.9884
R2319 B.n904 B.n15 32.9884
R2320 B.n904 B.n903 32.9884
R2321 B.n903 B.n902 32.9884
R2322 B.n902 B.n22 32.9884
R2323 B.n896 B.n895 32.9884
R2324 B.n895 B.n894 32.9884
R2325 B.n894 B.n29 32.9884
R2326 B.n888 B.n29 32.9884
R2327 B.n888 B.n887 32.9884
R2328 B.n887 B.n886 32.9884
R2329 B.n886 B.n36 32.9884
R2330 B.n880 B.n36 32.9884
R2331 B.n880 B.n879 32.9884
R2332 B.n878 B.n43 32.9884
R2333 B.n872 B.n43 32.9884
R2334 B.n872 B.n871 32.9884
R2335 B.n871 B.n870 32.9884
R2336 B.n870 B.n50 32.9884
R2337 B.n864 B.n50 32.9884
R2338 B.n866 B.n52 31.6883
R2339 B.n861 B.n860 31.6883
R2340 B.n740 B.n739 31.6883
R2341 B.n744 B.n421 31.6883
R2342 B.n815 B.t1 31.0479
R2343 B.n912 B.t2 31.0479
R2344 B.t0 B.n387 20.3754
R2345 B.t3 B.n22 20.3754
R2346 B B.n922 18.0485
R2347 B.n760 B.t5 16.4944
R2348 B.t5 B.n407 16.4944
R2349 B.n879 B.t12 16.4944
R2350 B.t12 B.n878 16.4944
R2351 B.n790 B.t0 12.6135
R2352 B.n896 B.t3 12.6135
R2353 B.n123 B.n52 10.6151
R2354 B.n126 B.n123 10.6151
R2355 B.n127 B.n126 10.6151
R2356 B.n130 B.n127 10.6151
R2357 B.n131 B.n130 10.6151
R2358 B.n134 B.n131 10.6151
R2359 B.n135 B.n134 10.6151
R2360 B.n138 B.n135 10.6151
R2361 B.n139 B.n138 10.6151
R2362 B.n142 B.n139 10.6151
R2363 B.n143 B.n142 10.6151
R2364 B.n146 B.n143 10.6151
R2365 B.n147 B.n146 10.6151
R2366 B.n150 B.n147 10.6151
R2367 B.n151 B.n150 10.6151
R2368 B.n154 B.n151 10.6151
R2369 B.n155 B.n154 10.6151
R2370 B.n158 B.n155 10.6151
R2371 B.n159 B.n158 10.6151
R2372 B.n162 B.n159 10.6151
R2373 B.n163 B.n162 10.6151
R2374 B.n166 B.n163 10.6151
R2375 B.n167 B.n166 10.6151
R2376 B.n170 B.n167 10.6151
R2377 B.n171 B.n170 10.6151
R2378 B.n174 B.n171 10.6151
R2379 B.n175 B.n174 10.6151
R2380 B.n178 B.n175 10.6151
R2381 B.n179 B.n178 10.6151
R2382 B.n182 B.n179 10.6151
R2383 B.n183 B.n182 10.6151
R2384 B.n186 B.n183 10.6151
R2385 B.n187 B.n186 10.6151
R2386 B.n190 B.n187 10.6151
R2387 B.n191 B.n190 10.6151
R2388 B.n194 B.n191 10.6151
R2389 B.n195 B.n194 10.6151
R2390 B.n198 B.n195 10.6151
R2391 B.n199 B.n198 10.6151
R2392 B.n202 B.n199 10.6151
R2393 B.n203 B.n202 10.6151
R2394 B.n206 B.n203 10.6151
R2395 B.n207 B.n206 10.6151
R2396 B.n210 B.n207 10.6151
R2397 B.n211 B.n210 10.6151
R2398 B.n214 B.n211 10.6151
R2399 B.n215 B.n214 10.6151
R2400 B.n218 B.n215 10.6151
R2401 B.n219 B.n218 10.6151
R2402 B.n222 B.n219 10.6151
R2403 B.n223 B.n222 10.6151
R2404 B.n226 B.n223 10.6151
R2405 B.n227 B.n226 10.6151
R2406 B.n230 B.n227 10.6151
R2407 B.n231 B.n230 10.6151
R2408 B.n234 B.n231 10.6151
R2409 B.n235 B.n234 10.6151
R2410 B.n239 B.n238 10.6151
R2411 B.n242 B.n239 10.6151
R2412 B.n243 B.n242 10.6151
R2413 B.n246 B.n243 10.6151
R2414 B.n247 B.n246 10.6151
R2415 B.n250 B.n247 10.6151
R2416 B.n251 B.n250 10.6151
R2417 B.n254 B.n251 10.6151
R2418 B.n259 B.n256 10.6151
R2419 B.n260 B.n259 10.6151
R2420 B.n263 B.n260 10.6151
R2421 B.n264 B.n263 10.6151
R2422 B.n267 B.n264 10.6151
R2423 B.n268 B.n267 10.6151
R2424 B.n271 B.n268 10.6151
R2425 B.n272 B.n271 10.6151
R2426 B.n275 B.n272 10.6151
R2427 B.n276 B.n275 10.6151
R2428 B.n279 B.n276 10.6151
R2429 B.n280 B.n279 10.6151
R2430 B.n283 B.n280 10.6151
R2431 B.n284 B.n283 10.6151
R2432 B.n287 B.n284 10.6151
R2433 B.n288 B.n287 10.6151
R2434 B.n291 B.n288 10.6151
R2435 B.n292 B.n291 10.6151
R2436 B.n295 B.n292 10.6151
R2437 B.n296 B.n295 10.6151
R2438 B.n299 B.n296 10.6151
R2439 B.n300 B.n299 10.6151
R2440 B.n303 B.n300 10.6151
R2441 B.n304 B.n303 10.6151
R2442 B.n307 B.n304 10.6151
R2443 B.n308 B.n307 10.6151
R2444 B.n311 B.n308 10.6151
R2445 B.n312 B.n311 10.6151
R2446 B.n315 B.n312 10.6151
R2447 B.n316 B.n315 10.6151
R2448 B.n319 B.n316 10.6151
R2449 B.n320 B.n319 10.6151
R2450 B.n323 B.n320 10.6151
R2451 B.n324 B.n323 10.6151
R2452 B.n327 B.n324 10.6151
R2453 B.n328 B.n327 10.6151
R2454 B.n331 B.n328 10.6151
R2455 B.n332 B.n331 10.6151
R2456 B.n335 B.n332 10.6151
R2457 B.n336 B.n335 10.6151
R2458 B.n339 B.n336 10.6151
R2459 B.n340 B.n339 10.6151
R2460 B.n343 B.n340 10.6151
R2461 B.n344 B.n343 10.6151
R2462 B.n347 B.n344 10.6151
R2463 B.n348 B.n347 10.6151
R2464 B.n351 B.n348 10.6151
R2465 B.n352 B.n351 10.6151
R2466 B.n355 B.n352 10.6151
R2467 B.n356 B.n355 10.6151
R2468 B.n359 B.n356 10.6151
R2469 B.n360 B.n359 10.6151
R2470 B.n363 B.n360 10.6151
R2471 B.n364 B.n363 10.6151
R2472 B.n367 B.n364 10.6151
R2473 B.n368 B.n367 10.6151
R2474 B.n861 B.n368 10.6151
R2475 B.n740 B.n417 10.6151
R2476 B.n750 B.n417 10.6151
R2477 B.n751 B.n750 10.6151
R2478 B.n752 B.n751 10.6151
R2479 B.n752 B.n409 10.6151
R2480 B.n762 B.n409 10.6151
R2481 B.n763 B.n762 10.6151
R2482 B.n764 B.n763 10.6151
R2483 B.n764 B.n401 10.6151
R2484 B.n774 B.n401 10.6151
R2485 B.n775 B.n774 10.6151
R2486 B.n776 B.n775 10.6151
R2487 B.n776 B.n393 10.6151
R2488 B.n786 B.n393 10.6151
R2489 B.n787 B.n786 10.6151
R2490 B.n788 B.n787 10.6151
R2491 B.n788 B.n385 10.6151
R2492 B.n798 B.n385 10.6151
R2493 B.n799 B.n798 10.6151
R2494 B.n800 B.n799 10.6151
R2495 B.n800 B.n376 10.6151
R2496 B.n810 B.n376 10.6151
R2497 B.n811 B.n810 10.6151
R2498 B.n813 B.n811 10.6151
R2499 B.n813 B.n812 10.6151
R2500 B.n812 B.n369 10.6151
R2501 B.n824 B.n369 10.6151
R2502 B.n825 B.n824 10.6151
R2503 B.n826 B.n825 10.6151
R2504 B.n827 B.n826 10.6151
R2505 B.n829 B.n827 10.6151
R2506 B.n830 B.n829 10.6151
R2507 B.n831 B.n830 10.6151
R2508 B.n832 B.n831 10.6151
R2509 B.n834 B.n832 10.6151
R2510 B.n835 B.n834 10.6151
R2511 B.n836 B.n835 10.6151
R2512 B.n837 B.n836 10.6151
R2513 B.n839 B.n837 10.6151
R2514 B.n840 B.n839 10.6151
R2515 B.n841 B.n840 10.6151
R2516 B.n842 B.n841 10.6151
R2517 B.n844 B.n842 10.6151
R2518 B.n845 B.n844 10.6151
R2519 B.n846 B.n845 10.6151
R2520 B.n847 B.n846 10.6151
R2521 B.n849 B.n847 10.6151
R2522 B.n850 B.n849 10.6151
R2523 B.n851 B.n850 10.6151
R2524 B.n852 B.n851 10.6151
R2525 B.n854 B.n852 10.6151
R2526 B.n855 B.n854 10.6151
R2527 B.n856 B.n855 10.6151
R2528 B.n857 B.n856 10.6151
R2529 B.n859 B.n857 10.6151
R2530 B.n860 B.n859 10.6151
R2531 B.n489 B.n421 10.6151
R2532 B.n489 B.n488 10.6151
R2533 B.n495 B.n488 10.6151
R2534 B.n496 B.n495 10.6151
R2535 B.n497 B.n496 10.6151
R2536 B.n497 B.n486 10.6151
R2537 B.n503 B.n486 10.6151
R2538 B.n504 B.n503 10.6151
R2539 B.n505 B.n504 10.6151
R2540 B.n505 B.n484 10.6151
R2541 B.n511 B.n484 10.6151
R2542 B.n512 B.n511 10.6151
R2543 B.n513 B.n512 10.6151
R2544 B.n513 B.n482 10.6151
R2545 B.n519 B.n482 10.6151
R2546 B.n520 B.n519 10.6151
R2547 B.n521 B.n520 10.6151
R2548 B.n521 B.n480 10.6151
R2549 B.n527 B.n480 10.6151
R2550 B.n528 B.n527 10.6151
R2551 B.n529 B.n528 10.6151
R2552 B.n529 B.n478 10.6151
R2553 B.n535 B.n478 10.6151
R2554 B.n536 B.n535 10.6151
R2555 B.n537 B.n536 10.6151
R2556 B.n537 B.n476 10.6151
R2557 B.n543 B.n476 10.6151
R2558 B.n544 B.n543 10.6151
R2559 B.n545 B.n544 10.6151
R2560 B.n545 B.n474 10.6151
R2561 B.n551 B.n474 10.6151
R2562 B.n552 B.n551 10.6151
R2563 B.n553 B.n552 10.6151
R2564 B.n553 B.n472 10.6151
R2565 B.n559 B.n472 10.6151
R2566 B.n560 B.n559 10.6151
R2567 B.n561 B.n560 10.6151
R2568 B.n561 B.n470 10.6151
R2569 B.n567 B.n470 10.6151
R2570 B.n568 B.n567 10.6151
R2571 B.n569 B.n568 10.6151
R2572 B.n569 B.n468 10.6151
R2573 B.n575 B.n468 10.6151
R2574 B.n576 B.n575 10.6151
R2575 B.n577 B.n576 10.6151
R2576 B.n577 B.n466 10.6151
R2577 B.n583 B.n466 10.6151
R2578 B.n584 B.n583 10.6151
R2579 B.n585 B.n584 10.6151
R2580 B.n585 B.n464 10.6151
R2581 B.n591 B.n464 10.6151
R2582 B.n592 B.n591 10.6151
R2583 B.n593 B.n592 10.6151
R2584 B.n593 B.n462 10.6151
R2585 B.n599 B.n462 10.6151
R2586 B.n600 B.n599 10.6151
R2587 B.n604 B.n600 10.6151
R2588 B.n610 B.n460 10.6151
R2589 B.n611 B.n610 10.6151
R2590 B.n612 B.n611 10.6151
R2591 B.n612 B.n458 10.6151
R2592 B.n618 B.n458 10.6151
R2593 B.n619 B.n618 10.6151
R2594 B.n620 B.n619 10.6151
R2595 B.n620 B.n456 10.6151
R2596 B.n627 B.n626 10.6151
R2597 B.n628 B.n627 10.6151
R2598 B.n628 B.n451 10.6151
R2599 B.n634 B.n451 10.6151
R2600 B.n635 B.n634 10.6151
R2601 B.n636 B.n635 10.6151
R2602 B.n636 B.n449 10.6151
R2603 B.n642 B.n449 10.6151
R2604 B.n643 B.n642 10.6151
R2605 B.n644 B.n643 10.6151
R2606 B.n644 B.n447 10.6151
R2607 B.n650 B.n447 10.6151
R2608 B.n651 B.n650 10.6151
R2609 B.n652 B.n651 10.6151
R2610 B.n652 B.n445 10.6151
R2611 B.n658 B.n445 10.6151
R2612 B.n659 B.n658 10.6151
R2613 B.n660 B.n659 10.6151
R2614 B.n660 B.n443 10.6151
R2615 B.n666 B.n443 10.6151
R2616 B.n667 B.n666 10.6151
R2617 B.n668 B.n667 10.6151
R2618 B.n668 B.n441 10.6151
R2619 B.n674 B.n441 10.6151
R2620 B.n675 B.n674 10.6151
R2621 B.n676 B.n675 10.6151
R2622 B.n676 B.n439 10.6151
R2623 B.n682 B.n439 10.6151
R2624 B.n683 B.n682 10.6151
R2625 B.n684 B.n683 10.6151
R2626 B.n684 B.n437 10.6151
R2627 B.n690 B.n437 10.6151
R2628 B.n691 B.n690 10.6151
R2629 B.n692 B.n691 10.6151
R2630 B.n692 B.n435 10.6151
R2631 B.n698 B.n435 10.6151
R2632 B.n699 B.n698 10.6151
R2633 B.n700 B.n699 10.6151
R2634 B.n700 B.n433 10.6151
R2635 B.n706 B.n433 10.6151
R2636 B.n707 B.n706 10.6151
R2637 B.n708 B.n707 10.6151
R2638 B.n708 B.n431 10.6151
R2639 B.n714 B.n431 10.6151
R2640 B.n715 B.n714 10.6151
R2641 B.n716 B.n715 10.6151
R2642 B.n716 B.n429 10.6151
R2643 B.n722 B.n429 10.6151
R2644 B.n723 B.n722 10.6151
R2645 B.n724 B.n723 10.6151
R2646 B.n724 B.n427 10.6151
R2647 B.n730 B.n427 10.6151
R2648 B.n731 B.n730 10.6151
R2649 B.n732 B.n731 10.6151
R2650 B.n732 B.n425 10.6151
R2651 B.n738 B.n425 10.6151
R2652 B.n739 B.n738 10.6151
R2653 B.n745 B.n744 10.6151
R2654 B.n746 B.n745 10.6151
R2655 B.n746 B.n413 10.6151
R2656 B.n756 B.n413 10.6151
R2657 B.n757 B.n756 10.6151
R2658 B.n758 B.n757 10.6151
R2659 B.n758 B.n405 10.6151
R2660 B.n768 B.n405 10.6151
R2661 B.n769 B.n768 10.6151
R2662 B.n770 B.n769 10.6151
R2663 B.n770 B.n397 10.6151
R2664 B.n780 B.n397 10.6151
R2665 B.n781 B.n780 10.6151
R2666 B.n782 B.n781 10.6151
R2667 B.n782 B.n389 10.6151
R2668 B.n792 B.n389 10.6151
R2669 B.n793 B.n792 10.6151
R2670 B.n794 B.n793 10.6151
R2671 B.n794 B.n381 10.6151
R2672 B.n804 B.n381 10.6151
R2673 B.n805 B.n804 10.6151
R2674 B.n806 B.n805 10.6151
R2675 B.n806 B.n373 10.6151
R2676 B.n817 B.n373 10.6151
R2677 B.n818 B.n817 10.6151
R2678 B.n819 B.n818 10.6151
R2679 B.n819 B.n0 10.6151
R2680 B.n916 B.n1 10.6151
R2681 B.n916 B.n915 10.6151
R2682 B.n915 B.n914 10.6151
R2683 B.n914 B.n10 10.6151
R2684 B.n908 B.n10 10.6151
R2685 B.n908 B.n907 10.6151
R2686 B.n907 B.n906 10.6151
R2687 B.n906 B.n17 10.6151
R2688 B.n900 B.n17 10.6151
R2689 B.n900 B.n899 10.6151
R2690 B.n899 B.n898 10.6151
R2691 B.n898 B.n24 10.6151
R2692 B.n892 B.n24 10.6151
R2693 B.n892 B.n891 10.6151
R2694 B.n891 B.n890 10.6151
R2695 B.n890 B.n31 10.6151
R2696 B.n884 B.n31 10.6151
R2697 B.n884 B.n883 10.6151
R2698 B.n883 B.n882 10.6151
R2699 B.n882 B.n38 10.6151
R2700 B.n876 B.n38 10.6151
R2701 B.n876 B.n875 10.6151
R2702 B.n875 B.n874 10.6151
R2703 B.n874 B.n45 10.6151
R2704 B.n868 B.n45 10.6151
R2705 B.n868 B.n867 10.6151
R2706 B.n867 B.n866 10.6151
R2707 B.n238 B.n122 6.5566
R2708 B.n255 B.n254 6.5566
R2709 B.n603 B.n460 6.5566
R2710 B.n456 B.n455 6.5566
R2711 B.n235 B.n122 4.05904
R2712 B.n256 B.n255 4.05904
R2713 B.n604 B.n603 4.05904
R2714 B.n626 B.n455 4.05904
R2715 B.n922 B.n0 2.81026
R2716 B.n922 B.n1 2.81026
R2717 B.n379 B.t1 1.94096
R2718 B.t2 B.n911 1.94096
R2719 VP.n2 VP.t1 251.471
R2720 VP.n2 VP.t3 250.948
R2721 VP.n4 VP.t2 216.155
R2722 VP.n11 VP.t0 216.155
R2723 VP.n10 VP.n0 161.3
R2724 VP.n9 VP.n8 161.3
R2725 VP.n7 VP.n1 161.3
R2726 VP.n6 VP.n5 161.3
R2727 VP.n4 VP.n3 91.9725
R2728 VP.n12 VP.n11 91.9725
R2729 VP.n9 VP.n1 56.5617
R2730 VP.n3 VP.n2 55.7894
R2731 VP.n5 VP.n1 24.5923
R2732 VP.n10 VP.n9 24.5923
R2733 VP.n5 VP.n4 18.9362
R2734 VP.n11 VP.n10 18.9362
R2735 VP.n6 VP.n3 0.278335
R2736 VP.n12 VP.n0 0.278335
R2737 VP.n7 VP.n6 0.189894
R2738 VP.n8 VP.n7 0.189894
R2739 VP.n8 VP.n0 0.189894
R2740 VP VP.n12 0.153485
R2741 VDD1 VDD1.n1 109.809
R2742 VDD1 VDD1.n0 64.7576
R2743 VDD1.n0 VDD1.t2 1.13843
R2744 VDD1.n0 VDD1.t0 1.13843
R2745 VDD1.n1 VDD1.t1 1.13843
R2746 VDD1.n1 VDD1.t3 1.13843
C0 VN VP 6.71509f
C1 VDD2 VP 0.352766f
C2 VTAIL VP 5.95941f
C3 VDD1 VN 0.148862f
C4 VDD1 VDD2 0.86879f
C5 VDD1 VTAIL 6.83662f
C6 VDD2 VN 6.34588f
C7 VN VTAIL 5.9453f
C8 VDD2 VTAIL 6.8864f
C9 VDD1 VP 6.54922f
C10 VDD2 B 3.814895f
C11 VDD1 B 8.270161f
C12 VTAIL B 12.893569f
C13 VN B 10.010799f
C14 VP B 7.907845f
C15 VDD1.t2 B 0.363351f
C16 VDD1.t0 B 0.363351f
C17 VDD1.n0 B 3.3177f
C18 VDD1.t1 B 0.363351f
C19 VDD1.t3 B 0.363351f
C20 VDD1.n1 B 4.14097f
C21 VP.n0 B 0.039249f
C22 VP.t0 B 2.76246f
C23 VP.n1 B 0.043278f
C24 VP.t3 B 2.91701f
C25 VP.t1 B 2.91935f
C26 VP.n2 B 3.52015f
C27 VP.n3 B 1.82278f
C28 VP.t2 B 2.76246f
C29 VP.n4 B 1.05246f
C30 VP.n5 B 0.04894f
C31 VP.n6 B 0.039249f
C32 VP.n7 B 0.029772f
C33 VP.n8 B 0.029772f
C34 VP.n9 B 0.043278f
C35 VP.n10 B 0.04894f
C36 VP.n11 B 1.05246f
C37 VP.n12 B 0.036616f
C38 VDD2.t2 B 0.363285f
C39 VDD2.t3 B 0.363285f
C40 VDD2.n0 B 4.11321f
C41 VDD2.t0 B 0.363285f
C42 VDD2.t1 B 0.363285f
C43 VDD2.n1 B 3.31674f
C44 VDD2.n2 B 4.14462f
C45 VTAIL.n0 B 0.008577f
C46 VTAIL.n1 B 0.019291f
C47 VTAIL.n2 B 0.008641f
C48 VTAIL.n3 B 0.015188f
C49 VTAIL.n4 B 0.008161f
C50 VTAIL.n5 B 0.019291f
C51 VTAIL.n6 B 0.008641f
C52 VTAIL.n7 B 0.015188f
C53 VTAIL.n8 B 0.008161f
C54 VTAIL.n9 B 0.019291f
C55 VTAIL.n10 B 0.008641f
C56 VTAIL.n11 B 0.015188f
C57 VTAIL.n12 B 0.008161f
C58 VTAIL.n13 B 0.019291f
C59 VTAIL.n14 B 0.008641f
C60 VTAIL.n15 B 0.015188f
C61 VTAIL.n16 B 0.008161f
C62 VTAIL.n17 B 0.019291f
C63 VTAIL.n18 B 0.008641f
C64 VTAIL.n19 B 0.015188f
C65 VTAIL.n20 B 0.008401f
C66 VTAIL.n21 B 0.019291f
C67 VTAIL.n22 B 0.008641f
C68 VTAIL.n23 B 0.015188f
C69 VTAIL.n24 B 0.008161f
C70 VTAIL.n25 B 0.019291f
C71 VTAIL.n26 B 0.008641f
C72 VTAIL.n27 B 0.015188f
C73 VTAIL.n28 B 0.008161f
C74 VTAIL.n29 B 0.014468f
C75 VTAIL.n30 B 0.013637f
C76 VTAIL.t4 B 0.033022f
C77 VTAIL.n31 B 0.140991f
C78 VTAIL.n32 B 1.131f
C79 VTAIL.n33 B 0.008161f
C80 VTAIL.n34 B 0.008641f
C81 VTAIL.n35 B 0.019291f
C82 VTAIL.n36 B 0.019291f
C83 VTAIL.n37 B 0.008641f
C84 VTAIL.n38 B 0.008161f
C85 VTAIL.n39 B 0.015188f
C86 VTAIL.n40 B 0.015188f
C87 VTAIL.n41 B 0.008161f
C88 VTAIL.n42 B 0.008641f
C89 VTAIL.n43 B 0.019291f
C90 VTAIL.n44 B 0.019291f
C91 VTAIL.n45 B 0.008641f
C92 VTAIL.n46 B 0.008161f
C93 VTAIL.n47 B 0.015188f
C94 VTAIL.n48 B 0.015188f
C95 VTAIL.n49 B 0.008161f
C96 VTAIL.n50 B 0.008161f
C97 VTAIL.n51 B 0.008641f
C98 VTAIL.n52 B 0.019291f
C99 VTAIL.n53 B 0.019291f
C100 VTAIL.n54 B 0.019291f
C101 VTAIL.n55 B 0.008401f
C102 VTAIL.n56 B 0.008161f
C103 VTAIL.n57 B 0.015188f
C104 VTAIL.n58 B 0.015188f
C105 VTAIL.n59 B 0.008161f
C106 VTAIL.n60 B 0.008641f
C107 VTAIL.n61 B 0.019291f
C108 VTAIL.n62 B 0.019291f
C109 VTAIL.n63 B 0.008641f
C110 VTAIL.n64 B 0.008161f
C111 VTAIL.n65 B 0.015188f
C112 VTAIL.n66 B 0.015188f
C113 VTAIL.n67 B 0.008161f
C114 VTAIL.n68 B 0.008641f
C115 VTAIL.n69 B 0.019291f
C116 VTAIL.n70 B 0.019291f
C117 VTAIL.n71 B 0.008641f
C118 VTAIL.n72 B 0.008161f
C119 VTAIL.n73 B 0.015188f
C120 VTAIL.n74 B 0.015188f
C121 VTAIL.n75 B 0.008161f
C122 VTAIL.n76 B 0.008641f
C123 VTAIL.n77 B 0.019291f
C124 VTAIL.n78 B 0.019291f
C125 VTAIL.n79 B 0.008641f
C126 VTAIL.n80 B 0.008161f
C127 VTAIL.n81 B 0.015188f
C128 VTAIL.n82 B 0.015188f
C129 VTAIL.n83 B 0.008161f
C130 VTAIL.n84 B 0.008641f
C131 VTAIL.n85 B 0.019291f
C132 VTAIL.n86 B 0.019291f
C133 VTAIL.n87 B 0.008641f
C134 VTAIL.n88 B 0.008161f
C135 VTAIL.n89 B 0.015188f
C136 VTAIL.n90 B 0.040086f
C137 VTAIL.n91 B 0.008161f
C138 VTAIL.n92 B 0.008641f
C139 VTAIL.n93 B 0.038861f
C140 VTAIL.n94 B 0.033419f
C141 VTAIL.n95 B 0.088339f
C142 VTAIL.n96 B 0.008577f
C143 VTAIL.n97 B 0.019291f
C144 VTAIL.n98 B 0.008641f
C145 VTAIL.n99 B 0.015188f
C146 VTAIL.n100 B 0.008161f
C147 VTAIL.n101 B 0.019291f
C148 VTAIL.n102 B 0.008641f
C149 VTAIL.n103 B 0.015188f
C150 VTAIL.n104 B 0.008161f
C151 VTAIL.n105 B 0.019291f
C152 VTAIL.n106 B 0.008641f
C153 VTAIL.n107 B 0.015188f
C154 VTAIL.n108 B 0.008161f
C155 VTAIL.n109 B 0.019291f
C156 VTAIL.n110 B 0.008641f
C157 VTAIL.n111 B 0.015188f
C158 VTAIL.n112 B 0.008161f
C159 VTAIL.n113 B 0.019291f
C160 VTAIL.n114 B 0.008641f
C161 VTAIL.n115 B 0.015188f
C162 VTAIL.n116 B 0.008401f
C163 VTAIL.n117 B 0.019291f
C164 VTAIL.n118 B 0.008641f
C165 VTAIL.n119 B 0.015188f
C166 VTAIL.n120 B 0.008161f
C167 VTAIL.n121 B 0.019291f
C168 VTAIL.n122 B 0.008641f
C169 VTAIL.n123 B 0.015188f
C170 VTAIL.n124 B 0.008161f
C171 VTAIL.n125 B 0.014468f
C172 VTAIL.n126 B 0.013637f
C173 VTAIL.t1 B 0.033022f
C174 VTAIL.n127 B 0.140991f
C175 VTAIL.n128 B 1.131f
C176 VTAIL.n129 B 0.008161f
C177 VTAIL.n130 B 0.008641f
C178 VTAIL.n131 B 0.019291f
C179 VTAIL.n132 B 0.019291f
C180 VTAIL.n133 B 0.008641f
C181 VTAIL.n134 B 0.008161f
C182 VTAIL.n135 B 0.015188f
C183 VTAIL.n136 B 0.015188f
C184 VTAIL.n137 B 0.008161f
C185 VTAIL.n138 B 0.008641f
C186 VTAIL.n139 B 0.019291f
C187 VTAIL.n140 B 0.019291f
C188 VTAIL.n141 B 0.008641f
C189 VTAIL.n142 B 0.008161f
C190 VTAIL.n143 B 0.015188f
C191 VTAIL.n144 B 0.015188f
C192 VTAIL.n145 B 0.008161f
C193 VTAIL.n146 B 0.008161f
C194 VTAIL.n147 B 0.008641f
C195 VTAIL.n148 B 0.019291f
C196 VTAIL.n149 B 0.019291f
C197 VTAIL.n150 B 0.019291f
C198 VTAIL.n151 B 0.008401f
C199 VTAIL.n152 B 0.008161f
C200 VTAIL.n153 B 0.015188f
C201 VTAIL.n154 B 0.015188f
C202 VTAIL.n155 B 0.008161f
C203 VTAIL.n156 B 0.008641f
C204 VTAIL.n157 B 0.019291f
C205 VTAIL.n158 B 0.019291f
C206 VTAIL.n159 B 0.008641f
C207 VTAIL.n160 B 0.008161f
C208 VTAIL.n161 B 0.015188f
C209 VTAIL.n162 B 0.015188f
C210 VTAIL.n163 B 0.008161f
C211 VTAIL.n164 B 0.008641f
C212 VTAIL.n165 B 0.019291f
C213 VTAIL.n166 B 0.019291f
C214 VTAIL.n167 B 0.008641f
C215 VTAIL.n168 B 0.008161f
C216 VTAIL.n169 B 0.015188f
C217 VTAIL.n170 B 0.015188f
C218 VTAIL.n171 B 0.008161f
C219 VTAIL.n172 B 0.008641f
C220 VTAIL.n173 B 0.019291f
C221 VTAIL.n174 B 0.019291f
C222 VTAIL.n175 B 0.008641f
C223 VTAIL.n176 B 0.008161f
C224 VTAIL.n177 B 0.015188f
C225 VTAIL.n178 B 0.015188f
C226 VTAIL.n179 B 0.008161f
C227 VTAIL.n180 B 0.008641f
C228 VTAIL.n181 B 0.019291f
C229 VTAIL.n182 B 0.019291f
C230 VTAIL.n183 B 0.008641f
C231 VTAIL.n184 B 0.008161f
C232 VTAIL.n185 B 0.015188f
C233 VTAIL.n186 B 0.040086f
C234 VTAIL.n187 B 0.008161f
C235 VTAIL.n188 B 0.008641f
C236 VTAIL.n189 B 0.038861f
C237 VTAIL.n190 B 0.033419f
C238 VTAIL.n191 B 0.133376f
C239 VTAIL.n192 B 0.008577f
C240 VTAIL.n193 B 0.019291f
C241 VTAIL.n194 B 0.008641f
C242 VTAIL.n195 B 0.015188f
C243 VTAIL.n196 B 0.008161f
C244 VTAIL.n197 B 0.019291f
C245 VTAIL.n198 B 0.008641f
C246 VTAIL.n199 B 0.015188f
C247 VTAIL.n200 B 0.008161f
C248 VTAIL.n201 B 0.019291f
C249 VTAIL.n202 B 0.008641f
C250 VTAIL.n203 B 0.015188f
C251 VTAIL.n204 B 0.008161f
C252 VTAIL.n205 B 0.019291f
C253 VTAIL.n206 B 0.008641f
C254 VTAIL.n207 B 0.015188f
C255 VTAIL.n208 B 0.008161f
C256 VTAIL.n209 B 0.019291f
C257 VTAIL.n210 B 0.008641f
C258 VTAIL.n211 B 0.015188f
C259 VTAIL.n212 B 0.008401f
C260 VTAIL.n213 B 0.019291f
C261 VTAIL.n214 B 0.008641f
C262 VTAIL.n215 B 0.015188f
C263 VTAIL.n216 B 0.008161f
C264 VTAIL.n217 B 0.019291f
C265 VTAIL.n218 B 0.008641f
C266 VTAIL.n219 B 0.015188f
C267 VTAIL.n220 B 0.008161f
C268 VTAIL.n221 B 0.014468f
C269 VTAIL.n222 B 0.013637f
C270 VTAIL.t0 B 0.033022f
C271 VTAIL.n223 B 0.140991f
C272 VTAIL.n224 B 1.131f
C273 VTAIL.n225 B 0.008161f
C274 VTAIL.n226 B 0.008641f
C275 VTAIL.n227 B 0.019291f
C276 VTAIL.n228 B 0.019291f
C277 VTAIL.n229 B 0.008641f
C278 VTAIL.n230 B 0.008161f
C279 VTAIL.n231 B 0.015188f
C280 VTAIL.n232 B 0.015188f
C281 VTAIL.n233 B 0.008161f
C282 VTAIL.n234 B 0.008641f
C283 VTAIL.n235 B 0.019291f
C284 VTAIL.n236 B 0.019291f
C285 VTAIL.n237 B 0.008641f
C286 VTAIL.n238 B 0.008161f
C287 VTAIL.n239 B 0.015188f
C288 VTAIL.n240 B 0.015188f
C289 VTAIL.n241 B 0.008161f
C290 VTAIL.n242 B 0.008161f
C291 VTAIL.n243 B 0.008641f
C292 VTAIL.n244 B 0.019291f
C293 VTAIL.n245 B 0.019291f
C294 VTAIL.n246 B 0.019291f
C295 VTAIL.n247 B 0.008401f
C296 VTAIL.n248 B 0.008161f
C297 VTAIL.n249 B 0.015188f
C298 VTAIL.n250 B 0.015188f
C299 VTAIL.n251 B 0.008161f
C300 VTAIL.n252 B 0.008641f
C301 VTAIL.n253 B 0.019291f
C302 VTAIL.n254 B 0.019291f
C303 VTAIL.n255 B 0.008641f
C304 VTAIL.n256 B 0.008161f
C305 VTAIL.n257 B 0.015188f
C306 VTAIL.n258 B 0.015188f
C307 VTAIL.n259 B 0.008161f
C308 VTAIL.n260 B 0.008641f
C309 VTAIL.n261 B 0.019291f
C310 VTAIL.n262 B 0.019291f
C311 VTAIL.n263 B 0.008641f
C312 VTAIL.n264 B 0.008161f
C313 VTAIL.n265 B 0.015188f
C314 VTAIL.n266 B 0.015188f
C315 VTAIL.n267 B 0.008161f
C316 VTAIL.n268 B 0.008641f
C317 VTAIL.n269 B 0.019291f
C318 VTAIL.n270 B 0.019291f
C319 VTAIL.n271 B 0.008641f
C320 VTAIL.n272 B 0.008161f
C321 VTAIL.n273 B 0.015188f
C322 VTAIL.n274 B 0.015188f
C323 VTAIL.n275 B 0.008161f
C324 VTAIL.n276 B 0.008641f
C325 VTAIL.n277 B 0.019291f
C326 VTAIL.n278 B 0.019291f
C327 VTAIL.n279 B 0.008641f
C328 VTAIL.n280 B 0.008161f
C329 VTAIL.n281 B 0.015188f
C330 VTAIL.n282 B 0.040086f
C331 VTAIL.n283 B 0.008161f
C332 VTAIL.n284 B 0.008641f
C333 VTAIL.n285 B 0.038861f
C334 VTAIL.n286 B 0.033419f
C335 VTAIL.n287 B 1.14655f
C336 VTAIL.n288 B 0.008577f
C337 VTAIL.n289 B 0.019291f
C338 VTAIL.n290 B 0.008641f
C339 VTAIL.n291 B 0.015188f
C340 VTAIL.n292 B 0.008161f
C341 VTAIL.n293 B 0.019291f
C342 VTAIL.n294 B 0.008641f
C343 VTAIL.n295 B 0.015188f
C344 VTAIL.n296 B 0.008161f
C345 VTAIL.n297 B 0.019291f
C346 VTAIL.n298 B 0.008641f
C347 VTAIL.n299 B 0.015188f
C348 VTAIL.n300 B 0.008161f
C349 VTAIL.n301 B 0.019291f
C350 VTAIL.n302 B 0.008641f
C351 VTAIL.n303 B 0.015188f
C352 VTAIL.n304 B 0.008161f
C353 VTAIL.n305 B 0.019291f
C354 VTAIL.n306 B 0.008641f
C355 VTAIL.n307 B 0.015188f
C356 VTAIL.n308 B 0.008401f
C357 VTAIL.n309 B 0.019291f
C358 VTAIL.n310 B 0.008161f
C359 VTAIL.n311 B 0.008641f
C360 VTAIL.n312 B 0.015188f
C361 VTAIL.n313 B 0.008161f
C362 VTAIL.n314 B 0.019291f
C363 VTAIL.n315 B 0.008641f
C364 VTAIL.n316 B 0.015188f
C365 VTAIL.n317 B 0.008161f
C366 VTAIL.n318 B 0.014468f
C367 VTAIL.n319 B 0.013637f
C368 VTAIL.t5 B 0.033022f
C369 VTAIL.n320 B 0.140991f
C370 VTAIL.n321 B 1.131f
C371 VTAIL.n322 B 0.008161f
C372 VTAIL.n323 B 0.008641f
C373 VTAIL.n324 B 0.019291f
C374 VTAIL.n325 B 0.019291f
C375 VTAIL.n326 B 0.008641f
C376 VTAIL.n327 B 0.008161f
C377 VTAIL.n328 B 0.015188f
C378 VTAIL.n329 B 0.015188f
C379 VTAIL.n330 B 0.008161f
C380 VTAIL.n331 B 0.008641f
C381 VTAIL.n332 B 0.019291f
C382 VTAIL.n333 B 0.019291f
C383 VTAIL.n334 B 0.008641f
C384 VTAIL.n335 B 0.008161f
C385 VTAIL.n336 B 0.015188f
C386 VTAIL.n337 B 0.015188f
C387 VTAIL.n338 B 0.008161f
C388 VTAIL.n339 B 0.008641f
C389 VTAIL.n340 B 0.019291f
C390 VTAIL.n341 B 0.019291f
C391 VTAIL.n342 B 0.019291f
C392 VTAIL.n343 B 0.008401f
C393 VTAIL.n344 B 0.008161f
C394 VTAIL.n345 B 0.015188f
C395 VTAIL.n346 B 0.015188f
C396 VTAIL.n347 B 0.008161f
C397 VTAIL.n348 B 0.008641f
C398 VTAIL.n349 B 0.019291f
C399 VTAIL.n350 B 0.019291f
C400 VTAIL.n351 B 0.008641f
C401 VTAIL.n352 B 0.008161f
C402 VTAIL.n353 B 0.015188f
C403 VTAIL.n354 B 0.015188f
C404 VTAIL.n355 B 0.008161f
C405 VTAIL.n356 B 0.008641f
C406 VTAIL.n357 B 0.019291f
C407 VTAIL.n358 B 0.019291f
C408 VTAIL.n359 B 0.008641f
C409 VTAIL.n360 B 0.008161f
C410 VTAIL.n361 B 0.015188f
C411 VTAIL.n362 B 0.015188f
C412 VTAIL.n363 B 0.008161f
C413 VTAIL.n364 B 0.008641f
C414 VTAIL.n365 B 0.019291f
C415 VTAIL.n366 B 0.019291f
C416 VTAIL.n367 B 0.008641f
C417 VTAIL.n368 B 0.008161f
C418 VTAIL.n369 B 0.015188f
C419 VTAIL.n370 B 0.015188f
C420 VTAIL.n371 B 0.008161f
C421 VTAIL.n372 B 0.008641f
C422 VTAIL.n373 B 0.019291f
C423 VTAIL.n374 B 0.019291f
C424 VTAIL.n375 B 0.008641f
C425 VTAIL.n376 B 0.008161f
C426 VTAIL.n377 B 0.015188f
C427 VTAIL.n378 B 0.040086f
C428 VTAIL.n379 B 0.008161f
C429 VTAIL.n380 B 0.008641f
C430 VTAIL.n381 B 0.038861f
C431 VTAIL.n382 B 0.033419f
C432 VTAIL.n383 B 1.14655f
C433 VTAIL.n384 B 0.008577f
C434 VTAIL.n385 B 0.019291f
C435 VTAIL.n386 B 0.008641f
C436 VTAIL.n387 B 0.015188f
C437 VTAIL.n388 B 0.008161f
C438 VTAIL.n389 B 0.019291f
C439 VTAIL.n390 B 0.008641f
C440 VTAIL.n391 B 0.015188f
C441 VTAIL.n392 B 0.008161f
C442 VTAIL.n393 B 0.019291f
C443 VTAIL.n394 B 0.008641f
C444 VTAIL.n395 B 0.015188f
C445 VTAIL.n396 B 0.008161f
C446 VTAIL.n397 B 0.019291f
C447 VTAIL.n398 B 0.008641f
C448 VTAIL.n399 B 0.015188f
C449 VTAIL.n400 B 0.008161f
C450 VTAIL.n401 B 0.019291f
C451 VTAIL.n402 B 0.008641f
C452 VTAIL.n403 B 0.015188f
C453 VTAIL.n404 B 0.008401f
C454 VTAIL.n405 B 0.019291f
C455 VTAIL.n406 B 0.008161f
C456 VTAIL.n407 B 0.008641f
C457 VTAIL.n408 B 0.015188f
C458 VTAIL.n409 B 0.008161f
C459 VTAIL.n410 B 0.019291f
C460 VTAIL.n411 B 0.008641f
C461 VTAIL.n412 B 0.015188f
C462 VTAIL.n413 B 0.008161f
C463 VTAIL.n414 B 0.014468f
C464 VTAIL.n415 B 0.013637f
C465 VTAIL.t6 B 0.033022f
C466 VTAIL.n416 B 0.140991f
C467 VTAIL.n417 B 1.131f
C468 VTAIL.n418 B 0.008161f
C469 VTAIL.n419 B 0.008641f
C470 VTAIL.n420 B 0.019291f
C471 VTAIL.n421 B 0.019291f
C472 VTAIL.n422 B 0.008641f
C473 VTAIL.n423 B 0.008161f
C474 VTAIL.n424 B 0.015188f
C475 VTAIL.n425 B 0.015188f
C476 VTAIL.n426 B 0.008161f
C477 VTAIL.n427 B 0.008641f
C478 VTAIL.n428 B 0.019291f
C479 VTAIL.n429 B 0.019291f
C480 VTAIL.n430 B 0.008641f
C481 VTAIL.n431 B 0.008161f
C482 VTAIL.n432 B 0.015188f
C483 VTAIL.n433 B 0.015188f
C484 VTAIL.n434 B 0.008161f
C485 VTAIL.n435 B 0.008641f
C486 VTAIL.n436 B 0.019291f
C487 VTAIL.n437 B 0.019291f
C488 VTAIL.n438 B 0.019291f
C489 VTAIL.n439 B 0.008401f
C490 VTAIL.n440 B 0.008161f
C491 VTAIL.n441 B 0.015188f
C492 VTAIL.n442 B 0.015188f
C493 VTAIL.n443 B 0.008161f
C494 VTAIL.n444 B 0.008641f
C495 VTAIL.n445 B 0.019291f
C496 VTAIL.n446 B 0.019291f
C497 VTAIL.n447 B 0.008641f
C498 VTAIL.n448 B 0.008161f
C499 VTAIL.n449 B 0.015188f
C500 VTAIL.n450 B 0.015188f
C501 VTAIL.n451 B 0.008161f
C502 VTAIL.n452 B 0.008641f
C503 VTAIL.n453 B 0.019291f
C504 VTAIL.n454 B 0.019291f
C505 VTAIL.n455 B 0.008641f
C506 VTAIL.n456 B 0.008161f
C507 VTAIL.n457 B 0.015188f
C508 VTAIL.n458 B 0.015188f
C509 VTAIL.n459 B 0.008161f
C510 VTAIL.n460 B 0.008641f
C511 VTAIL.n461 B 0.019291f
C512 VTAIL.n462 B 0.019291f
C513 VTAIL.n463 B 0.008641f
C514 VTAIL.n464 B 0.008161f
C515 VTAIL.n465 B 0.015188f
C516 VTAIL.n466 B 0.015188f
C517 VTAIL.n467 B 0.008161f
C518 VTAIL.n468 B 0.008641f
C519 VTAIL.n469 B 0.019291f
C520 VTAIL.n470 B 0.019291f
C521 VTAIL.n471 B 0.008641f
C522 VTAIL.n472 B 0.008161f
C523 VTAIL.n473 B 0.015188f
C524 VTAIL.n474 B 0.040086f
C525 VTAIL.n475 B 0.008161f
C526 VTAIL.n476 B 0.008641f
C527 VTAIL.n477 B 0.038861f
C528 VTAIL.n478 B 0.033419f
C529 VTAIL.n479 B 0.133376f
C530 VTAIL.n480 B 0.008577f
C531 VTAIL.n481 B 0.019291f
C532 VTAIL.n482 B 0.008641f
C533 VTAIL.n483 B 0.015188f
C534 VTAIL.n484 B 0.008161f
C535 VTAIL.n485 B 0.019291f
C536 VTAIL.n486 B 0.008641f
C537 VTAIL.n487 B 0.015188f
C538 VTAIL.n488 B 0.008161f
C539 VTAIL.n489 B 0.019291f
C540 VTAIL.n490 B 0.008641f
C541 VTAIL.n491 B 0.015188f
C542 VTAIL.n492 B 0.008161f
C543 VTAIL.n493 B 0.019291f
C544 VTAIL.n494 B 0.008641f
C545 VTAIL.n495 B 0.015188f
C546 VTAIL.n496 B 0.008161f
C547 VTAIL.n497 B 0.019291f
C548 VTAIL.n498 B 0.008641f
C549 VTAIL.n499 B 0.015188f
C550 VTAIL.n500 B 0.008401f
C551 VTAIL.n501 B 0.019291f
C552 VTAIL.n502 B 0.008161f
C553 VTAIL.n503 B 0.008641f
C554 VTAIL.n504 B 0.015188f
C555 VTAIL.n505 B 0.008161f
C556 VTAIL.n506 B 0.019291f
C557 VTAIL.n507 B 0.008641f
C558 VTAIL.n508 B 0.015188f
C559 VTAIL.n509 B 0.008161f
C560 VTAIL.n510 B 0.014468f
C561 VTAIL.n511 B 0.013637f
C562 VTAIL.t2 B 0.033022f
C563 VTAIL.n512 B 0.140991f
C564 VTAIL.n513 B 1.131f
C565 VTAIL.n514 B 0.008161f
C566 VTAIL.n515 B 0.008641f
C567 VTAIL.n516 B 0.019291f
C568 VTAIL.n517 B 0.019291f
C569 VTAIL.n518 B 0.008641f
C570 VTAIL.n519 B 0.008161f
C571 VTAIL.n520 B 0.015188f
C572 VTAIL.n521 B 0.015188f
C573 VTAIL.n522 B 0.008161f
C574 VTAIL.n523 B 0.008641f
C575 VTAIL.n524 B 0.019291f
C576 VTAIL.n525 B 0.019291f
C577 VTAIL.n526 B 0.008641f
C578 VTAIL.n527 B 0.008161f
C579 VTAIL.n528 B 0.015188f
C580 VTAIL.n529 B 0.015188f
C581 VTAIL.n530 B 0.008161f
C582 VTAIL.n531 B 0.008641f
C583 VTAIL.n532 B 0.019291f
C584 VTAIL.n533 B 0.019291f
C585 VTAIL.n534 B 0.019291f
C586 VTAIL.n535 B 0.008401f
C587 VTAIL.n536 B 0.008161f
C588 VTAIL.n537 B 0.015188f
C589 VTAIL.n538 B 0.015188f
C590 VTAIL.n539 B 0.008161f
C591 VTAIL.n540 B 0.008641f
C592 VTAIL.n541 B 0.019291f
C593 VTAIL.n542 B 0.019291f
C594 VTAIL.n543 B 0.008641f
C595 VTAIL.n544 B 0.008161f
C596 VTAIL.n545 B 0.015188f
C597 VTAIL.n546 B 0.015188f
C598 VTAIL.n547 B 0.008161f
C599 VTAIL.n548 B 0.008641f
C600 VTAIL.n549 B 0.019291f
C601 VTAIL.n550 B 0.019291f
C602 VTAIL.n551 B 0.008641f
C603 VTAIL.n552 B 0.008161f
C604 VTAIL.n553 B 0.015188f
C605 VTAIL.n554 B 0.015188f
C606 VTAIL.n555 B 0.008161f
C607 VTAIL.n556 B 0.008641f
C608 VTAIL.n557 B 0.019291f
C609 VTAIL.n558 B 0.019291f
C610 VTAIL.n559 B 0.008641f
C611 VTAIL.n560 B 0.008161f
C612 VTAIL.n561 B 0.015188f
C613 VTAIL.n562 B 0.015188f
C614 VTAIL.n563 B 0.008161f
C615 VTAIL.n564 B 0.008641f
C616 VTAIL.n565 B 0.019291f
C617 VTAIL.n566 B 0.019291f
C618 VTAIL.n567 B 0.008641f
C619 VTAIL.n568 B 0.008161f
C620 VTAIL.n569 B 0.015188f
C621 VTAIL.n570 B 0.040086f
C622 VTAIL.n571 B 0.008161f
C623 VTAIL.n572 B 0.008641f
C624 VTAIL.n573 B 0.038861f
C625 VTAIL.n574 B 0.033419f
C626 VTAIL.n575 B 0.133376f
C627 VTAIL.n576 B 0.008577f
C628 VTAIL.n577 B 0.019291f
C629 VTAIL.n578 B 0.008641f
C630 VTAIL.n579 B 0.015188f
C631 VTAIL.n580 B 0.008161f
C632 VTAIL.n581 B 0.019291f
C633 VTAIL.n582 B 0.008641f
C634 VTAIL.n583 B 0.015188f
C635 VTAIL.n584 B 0.008161f
C636 VTAIL.n585 B 0.019291f
C637 VTAIL.n586 B 0.008641f
C638 VTAIL.n587 B 0.015188f
C639 VTAIL.n588 B 0.008161f
C640 VTAIL.n589 B 0.019291f
C641 VTAIL.n590 B 0.008641f
C642 VTAIL.n591 B 0.015188f
C643 VTAIL.n592 B 0.008161f
C644 VTAIL.n593 B 0.019291f
C645 VTAIL.n594 B 0.008641f
C646 VTAIL.n595 B 0.015188f
C647 VTAIL.n596 B 0.008401f
C648 VTAIL.n597 B 0.019291f
C649 VTAIL.n598 B 0.008161f
C650 VTAIL.n599 B 0.008641f
C651 VTAIL.n600 B 0.015188f
C652 VTAIL.n601 B 0.008161f
C653 VTAIL.n602 B 0.019291f
C654 VTAIL.n603 B 0.008641f
C655 VTAIL.n604 B 0.015188f
C656 VTAIL.n605 B 0.008161f
C657 VTAIL.n606 B 0.014468f
C658 VTAIL.n607 B 0.013637f
C659 VTAIL.t3 B 0.033022f
C660 VTAIL.n608 B 0.140991f
C661 VTAIL.n609 B 1.131f
C662 VTAIL.n610 B 0.008161f
C663 VTAIL.n611 B 0.008641f
C664 VTAIL.n612 B 0.019291f
C665 VTAIL.n613 B 0.019291f
C666 VTAIL.n614 B 0.008641f
C667 VTAIL.n615 B 0.008161f
C668 VTAIL.n616 B 0.015188f
C669 VTAIL.n617 B 0.015188f
C670 VTAIL.n618 B 0.008161f
C671 VTAIL.n619 B 0.008641f
C672 VTAIL.n620 B 0.019291f
C673 VTAIL.n621 B 0.019291f
C674 VTAIL.n622 B 0.008641f
C675 VTAIL.n623 B 0.008161f
C676 VTAIL.n624 B 0.015188f
C677 VTAIL.n625 B 0.015188f
C678 VTAIL.n626 B 0.008161f
C679 VTAIL.n627 B 0.008641f
C680 VTAIL.n628 B 0.019291f
C681 VTAIL.n629 B 0.019291f
C682 VTAIL.n630 B 0.019291f
C683 VTAIL.n631 B 0.008401f
C684 VTAIL.n632 B 0.008161f
C685 VTAIL.n633 B 0.015188f
C686 VTAIL.n634 B 0.015188f
C687 VTAIL.n635 B 0.008161f
C688 VTAIL.n636 B 0.008641f
C689 VTAIL.n637 B 0.019291f
C690 VTAIL.n638 B 0.019291f
C691 VTAIL.n639 B 0.008641f
C692 VTAIL.n640 B 0.008161f
C693 VTAIL.n641 B 0.015188f
C694 VTAIL.n642 B 0.015188f
C695 VTAIL.n643 B 0.008161f
C696 VTAIL.n644 B 0.008641f
C697 VTAIL.n645 B 0.019291f
C698 VTAIL.n646 B 0.019291f
C699 VTAIL.n647 B 0.008641f
C700 VTAIL.n648 B 0.008161f
C701 VTAIL.n649 B 0.015188f
C702 VTAIL.n650 B 0.015188f
C703 VTAIL.n651 B 0.008161f
C704 VTAIL.n652 B 0.008641f
C705 VTAIL.n653 B 0.019291f
C706 VTAIL.n654 B 0.019291f
C707 VTAIL.n655 B 0.008641f
C708 VTAIL.n656 B 0.008161f
C709 VTAIL.n657 B 0.015188f
C710 VTAIL.n658 B 0.015188f
C711 VTAIL.n659 B 0.008161f
C712 VTAIL.n660 B 0.008641f
C713 VTAIL.n661 B 0.019291f
C714 VTAIL.n662 B 0.019291f
C715 VTAIL.n663 B 0.008641f
C716 VTAIL.n664 B 0.008161f
C717 VTAIL.n665 B 0.015188f
C718 VTAIL.n666 B 0.040086f
C719 VTAIL.n667 B 0.008161f
C720 VTAIL.n668 B 0.008641f
C721 VTAIL.n669 B 0.038861f
C722 VTAIL.n670 B 0.033419f
C723 VTAIL.n671 B 1.14655f
C724 VTAIL.n672 B 0.008577f
C725 VTAIL.n673 B 0.019291f
C726 VTAIL.n674 B 0.008641f
C727 VTAIL.n675 B 0.015188f
C728 VTAIL.n676 B 0.008161f
C729 VTAIL.n677 B 0.019291f
C730 VTAIL.n678 B 0.008641f
C731 VTAIL.n679 B 0.015188f
C732 VTAIL.n680 B 0.008161f
C733 VTAIL.n681 B 0.019291f
C734 VTAIL.n682 B 0.008641f
C735 VTAIL.n683 B 0.015188f
C736 VTAIL.n684 B 0.008161f
C737 VTAIL.n685 B 0.019291f
C738 VTAIL.n686 B 0.008641f
C739 VTAIL.n687 B 0.015188f
C740 VTAIL.n688 B 0.008161f
C741 VTAIL.n689 B 0.019291f
C742 VTAIL.n690 B 0.008641f
C743 VTAIL.n691 B 0.015188f
C744 VTAIL.n692 B 0.008401f
C745 VTAIL.n693 B 0.019291f
C746 VTAIL.n694 B 0.008641f
C747 VTAIL.n695 B 0.015188f
C748 VTAIL.n696 B 0.008161f
C749 VTAIL.n697 B 0.019291f
C750 VTAIL.n698 B 0.008641f
C751 VTAIL.n699 B 0.015188f
C752 VTAIL.n700 B 0.008161f
C753 VTAIL.n701 B 0.014468f
C754 VTAIL.n702 B 0.013637f
C755 VTAIL.t7 B 0.033022f
C756 VTAIL.n703 B 0.140991f
C757 VTAIL.n704 B 1.131f
C758 VTAIL.n705 B 0.008161f
C759 VTAIL.n706 B 0.008641f
C760 VTAIL.n707 B 0.019291f
C761 VTAIL.n708 B 0.019291f
C762 VTAIL.n709 B 0.008641f
C763 VTAIL.n710 B 0.008161f
C764 VTAIL.n711 B 0.015188f
C765 VTAIL.n712 B 0.015188f
C766 VTAIL.n713 B 0.008161f
C767 VTAIL.n714 B 0.008641f
C768 VTAIL.n715 B 0.019291f
C769 VTAIL.n716 B 0.019291f
C770 VTAIL.n717 B 0.008641f
C771 VTAIL.n718 B 0.008161f
C772 VTAIL.n719 B 0.015188f
C773 VTAIL.n720 B 0.015188f
C774 VTAIL.n721 B 0.008161f
C775 VTAIL.n722 B 0.008161f
C776 VTAIL.n723 B 0.008641f
C777 VTAIL.n724 B 0.019291f
C778 VTAIL.n725 B 0.019291f
C779 VTAIL.n726 B 0.019291f
C780 VTAIL.n727 B 0.008401f
C781 VTAIL.n728 B 0.008161f
C782 VTAIL.n729 B 0.015188f
C783 VTAIL.n730 B 0.015188f
C784 VTAIL.n731 B 0.008161f
C785 VTAIL.n732 B 0.008641f
C786 VTAIL.n733 B 0.019291f
C787 VTAIL.n734 B 0.019291f
C788 VTAIL.n735 B 0.008641f
C789 VTAIL.n736 B 0.008161f
C790 VTAIL.n737 B 0.015188f
C791 VTAIL.n738 B 0.015188f
C792 VTAIL.n739 B 0.008161f
C793 VTAIL.n740 B 0.008641f
C794 VTAIL.n741 B 0.019291f
C795 VTAIL.n742 B 0.019291f
C796 VTAIL.n743 B 0.008641f
C797 VTAIL.n744 B 0.008161f
C798 VTAIL.n745 B 0.015188f
C799 VTAIL.n746 B 0.015188f
C800 VTAIL.n747 B 0.008161f
C801 VTAIL.n748 B 0.008641f
C802 VTAIL.n749 B 0.019291f
C803 VTAIL.n750 B 0.019291f
C804 VTAIL.n751 B 0.008641f
C805 VTAIL.n752 B 0.008161f
C806 VTAIL.n753 B 0.015188f
C807 VTAIL.n754 B 0.015188f
C808 VTAIL.n755 B 0.008161f
C809 VTAIL.n756 B 0.008641f
C810 VTAIL.n757 B 0.019291f
C811 VTAIL.n758 B 0.019291f
C812 VTAIL.n759 B 0.008641f
C813 VTAIL.n760 B 0.008161f
C814 VTAIL.n761 B 0.015188f
C815 VTAIL.n762 B 0.040086f
C816 VTAIL.n763 B 0.008161f
C817 VTAIL.n764 B 0.008641f
C818 VTAIL.n765 B 0.038861f
C819 VTAIL.n766 B 0.033419f
C820 VTAIL.n767 B 1.09582f
C821 VN.t1 B 2.86749f
C822 VN.t0 B 2.86519f
C823 VN.n0 B 1.95438f
C824 VN.t2 B 2.86749f
C825 VN.t3 B 2.86519f
C826 VN.n1 B 3.47247f
.ends

