* NGSPICE file created from diff_pair_sample_1451.ext - technology: sky130A

.subckt diff_pair_sample_1451 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t3 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=2.145 pd=13.33 as=5.07 ps=26.78 w=13 l=0.29
X1 VTAIL.t7 VN.t0 VDD2.t3 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=2.145 ps=13.33 w=13 l=0.29
X2 B.t11 B.t9 B.t10 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=0 ps=0 w=13 l=0.29
X3 B.t8 B.t6 B.t7 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=0 ps=0 w=13 l=0.29
X4 B.t5 B.t3 B.t4 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=0 ps=0 w=13 l=0.29
X5 VDD2.t2 VN.t1 VTAIL.t2 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=2.145 pd=13.33 as=5.07 ps=26.78 w=13 l=0.29
X6 VDD1.t2 VP.t1 VTAIL.t4 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=2.145 pd=13.33 as=5.07 ps=26.78 w=13 l=0.29
X7 B.t2 B.t0 B.t1 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=0 ps=0 w=13 l=0.29
X8 VTAIL.t5 VP.t2 VDD1.t1 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=2.145 ps=13.33 w=13 l=0.29
X9 VTAIL.t1 VN.t2 VDD2.t1 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=2.145 ps=13.33 w=13 l=0.29
X10 VDD2.t0 VN.t3 VTAIL.t0 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=2.145 pd=13.33 as=5.07 ps=26.78 w=13 l=0.29
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n1342_n3572# sky130_fd_pr__pfet_01v8 ad=5.07 pd=26.78 as=2.145 ps=13.33 w=13 l=0.29
R0 VP.n1 VP.t1 1233.66
R1 VP.n1 VP.t2 1233.66
R2 VP.n0 VP.t3 1233.66
R3 VP.n0 VP.t0 1233.66
R4 VP.n2 VP.n0 201.309
R5 VP.n2 VP.n1 161.3
R6 VP VP.n2 0.0516364
R7 VTAIL.n5 VTAIL.t6 61.2344
R8 VTAIL.n4 VTAIL.t0 61.2344
R9 VTAIL.n3 VTAIL.t1 61.2344
R10 VTAIL.n7 VTAIL.t2 61.2332
R11 VTAIL.n0 VTAIL.t7 61.2332
R12 VTAIL.n1 VTAIL.t4 61.2332
R13 VTAIL.n2 VTAIL.t5 61.2332
R14 VTAIL.n6 VTAIL.t3 61.2332
R15 VTAIL.n7 VTAIL.n6 24.1255
R16 VTAIL.n3 VTAIL.n2 24.1255
R17 VTAIL.n4 VTAIL.n3 0.534983
R18 VTAIL.n6 VTAIL.n5 0.534983
R19 VTAIL.n2 VTAIL.n1 0.534983
R20 VTAIL.n5 VTAIL.n4 0.470328
R21 VTAIL.n1 VTAIL.n0 0.470328
R22 VTAIL VTAIL.n0 0.325931
R23 VTAIL VTAIL.n7 0.209552
R24 VDD1 VDD1.n1 112.478
R25 VDD1 VDD1.n0 75.4698
R26 VDD1.n0 VDD1.t0 2.50088
R27 VDD1.n0 VDD1.t3 2.50088
R28 VDD1.n1 VDD1.t1 2.50088
R29 VDD1.n1 VDD1.t2 2.50088
R30 VN.n0 VN.t1 1233.66
R31 VN.n0 VN.t0 1233.66
R32 VN.n1 VN.t2 1233.66
R33 VN.n1 VN.t3 1233.66
R34 VN VN.n1 201.689
R35 VN VN.n0 161.351
R36 VDD2.n2 VDD2.n0 111.954
R37 VDD2.n2 VDD2.n1 75.4117
R38 VDD2.n1 VDD2.t1 2.50088
R39 VDD2.n1 VDD2.t0 2.50088
R40 VDD2.n0 VDD2.t3 2.50088
R41 VDD2.n0 VDD2.t2 2.50088
R42 VDD2 VDD2.n2 0.0586897
R43 B.n104 B.t6 1298
R44 B.n232 B.t0 1298
R45 B.n38 B.t9 1298
R46 B.n32 B.t3 1298
R47 B.n303 B.n76 585
R48 B.n302 B.n301 585
R49 B.n300 B.n77 585
R50 B.n299 B.n298 585
R51 B.n297 B.n78 585
R52 B.n296 B.n295 585
R53 B.n294 B.n79 585
R54 B.n293 B.n292 585
R55 B.n291 B.n80 585
R56 B.n290 B.n289 585
R57 B.n288 B.n81 585
R58 B.n287 B.n286 585
R59 B.n285 B.n82 585
R60 B.n284 B.n283 585
R61 B.n282 B.n83 585
R62 B.n281 B.n280 585
R63 B.n279 B.n84 585
R64 B.n278 B.n277 585
R65 B.n276 B.n85 585
R66 B.n275 B.n274 585
R67 B.n273 B.n86 585
R68 B.n272 B.n271 585
R69 B.n270 B.n87 585
R70 B.n269 B.n268 585
R71 B.n267 B.n88 585
R72 B.n266 B.n265 585
R73 B.n264 B.n89 585
R74 B.n263 B.n262 585
R75 B.n261 B.n90 585
R76 B.n260 B.n259 585
R77 B.n258 B.n91 585
R78 B.n257 B.n256 585
R79 B.n255 B.n92 585
R80 B.n254 B.n253 585
R81 B.n252 B.n93 585
R82 B.n251 B.n250 585
R83 B.n249 B.n94 585
R84 B.n248 B.n247 585
R85 B.n246 B.n95 585
R86 B.n245 B.n244 585
R87 B.n243 B.n96 585
R88 B.n242 B.n241 585
R89 B.n240 B.n97 585
R90 B.n239 B.n238 585
R91 B.n237 B.n98 585
R92 B.n236 B.n235 585
R93 B.n231 B.n99 585
R94 B.n230 B.n229 585
R95 B.n228 B.n100 585
R96 B.n227 B.n226 585
R97 B.n225 B.n101 585
R98 B.n224 B.n223 585
R99 B.n222 B.n102 585
R100 B.n221 B.n220 585
R101 B.n218 B.n103 585
R102 B.n217 B.n216 585
R103 B.n215 B.n106 585
R104 B.n214 B.n213 585
R105 B.n212 B.n107 585
R106 B.n211 B.n210 585
R107 B.n209 B.n108 585
R108 B.n208 B.n207 585
R109 B.n206 B.n109 585
R110 B.n205 B.n204 585
R111 B.n203 B.n110 585
R112 B.n202 B.n201 585
R113 B.n200 B.n111 585
R114 B.n199 B.n198 585
R115 B.n197 B.n112 585
R116 B.n196 B.n195 585
R117 B.n194 B.n113 585
R118 B.n193 B.n192 585
R119 B.n191 B.n114 585
R120 B.n190 B.n189 585
R121 B.n188 B.n115 585
R122 B.n187 B.n186 585
R123 B.n185 B.n116 585
R124 B.n184 B.n183 585
R125 B.n182 B.n117 585
R126 B.n181 B.n180 585
R127 B.n179 B.n118 585
R128 B.n178 B.n177 585
R129 B.n176 B.n119 585
R130 B.n175 B.n174 585
R131 B.n173 B.n120 585
R132 B.n172 B.n171 585
R133 B.n170 B.n121 585
R134 B.n169 B.n168 585
R135 B.n167 B.n122 585
R136 B.n166 B.n165 585
R137 B.n164 B.n123 585
R138 B.n163 B.n162 585
R139 B.n161 B.n124 585
R140 B.n160 B.n159 585
R141 B.n158 B.n125 585
R142 B.n157 B.n156 585
R143 B.n155 B.n126 585
R144 B.n154 B.n153 585
R145 B.n152 B.n127 585
R146 B.n305 B.n304 585
R147 B.n306 B.n75 585
R148 B.n308 B.n307 585
R149 B.n309 B.n74 585
R150 B.n311 B.n310 585
R151 B.n312 B.n73 585
R152 B.n314 B.n313 585
R153 B.n315 B.n72 585
R154 B.n317 B.n316 585
R155 B.n318 B.n71 585
R156 B.n320 B.n319 585
R157 B.n321 B.n70 585
R158 B.n323 B.n322 585
R159 B.n324 B.n69 585
R160 B.n326 B.n325 585
R161 B.n327 B.n68 585
R162 B.n329 B.n328 585
R163 B.n330 B.n67 585
R164 B.n332 B.n331 585
R165 B.n333 B.n66 585
R166 B.n335 B.n334 585
R167 B.n336 B.n65 585
R168 B.n338 B.n337 585
R169 B.n339 B.n64 585
R170 B.n341 B.n340 585
R171 B.n342 B.n63 585
R172 B.n344 B.n343 585
R173 B.n345 B.n62 585
R174 B.n496 B.n495 585
R175 B.n494 B.n9 585
R176 B.n493 B.n492 585
R177 B.n491 B.n10 585
R178 B.n490 B.n489 585
R179 B.n488 B.n11 585
R180 B.n487 B.n486 585
R181 B.n485 B.n12 585
R182 B.n484 B.n483 585
R183 B.n482 B.n13 585
R184 B.n481 B.n480 585
R185 B.n479 B.n14 585
R186 B.n478 B.n477 585
R187 B.n476 B.n15 585
R188 B.n475 B.n474 585
R189 B.n473 B.n16 585
R190 B.n472 B.n471 585
R191 B.n470 B.n17 585
R192 B.n469 B.n468 585
R193 B.n467 B.n18 585
R194 B.n466 B.n465 585
R195 B.n464 B.n19 585
R196 B.n463 B.n462 585
R197 B.n461 B.n20 585
R198 B.n460 B.n459 585
R199 B.n458 B.n21 585
R200 B.n457 B.n456 585
R201 B.n455 B.n22 585
R202 B.n454 B.n453 585
R203 B.n452 B.n23 585
R204 B.n451 B.n450 585
R205 B.n449 B.n24 585
R206 B.n448 B.n447 585
R207 B.n446 B.n25 585
R208 B.n445 B.n444 585
R209 B.n443 B.n26 585
R210 B.n442 B.n441 585
R211 B.n440 B.n27 585
R212 B.n439 B.n438 585
R213 B.n437 B.n28 585
R214 B.n436 B.n435 585
R215 B.n434 B.n29 585
R216 B.n433 B.n432 585
R217 B.n431 B.n30 585
R218 B.n430 B.n429 585
R219 B.n427 B.n31 585
R220 B.n426 B.n425 585
R221 B.n424 B.n34 585
R222 B.n423 B.n422 585
R223 B.n421 B.n35 585
R224 B.n420 B.n419 585
R225 B.n418 B.n36 585
R226 B.n417 B.n416 585
R227 B.n415 B.n37 585
R228 B.n413 B.n412 585
R229 B.n411 B.n40 585
R230 B.n410 B.n409 585
R231 B.n408 B.n41 585
R232 B.n407 B.n406 585
R233 B.n405 B.n42 585
R234 B.n404 B.n403 585
R235 B.n402 B.n43 585
R236 B.n401 B.n400 585
R237 B.n399 B.n44 585
R238 B.n398 B.n397 585
R239 B.n396 B.n45 585
R240 B.n395 B.n394 585
R241 B.n393 B.n46 585
R242 B.n392 B.n391 585
R243 B.n390 B.n47 585
R244 B.n389 B.n388 585
R245 B.n387 B.n48 585
R246 B.n386 B.n385 585
R247 B.n384 B.n49 585
R248 B.n383 B.n382 585
R249 B.n381 B.n50 585
R250 B.n380 B.n379 585
R251 B.n378 B.n51 585
R252 B.n377 B.n376 585
R253 B.n375 B.n52 585
R254 B.n374 B.n373 585
R255 B.n372 B.n53 585
R256 B.n371 B.n370 585
R257 B.n369 B.n54 585
R258 B.n368 B.n367 585
R259 B.n366 B.n55 585
R260 B.n365 B.n364 585
R261 B.n363 B.n56 585
R262 B.n362 B.n361 585
R263 B.n360 B.n57 585
R264 B.n359 B.n358 585
R265 B.n357 B.n58 585
R266 B.n356 B.n355 585
R267 B.n354 B.n59 585
R268 B.n353 B.n352 585
R269 B.n351 B.n60 585
R270 B.n350 B.n349 585
R271 B.n348 B.n61 585
R272 B.n347 B.n346 585
R273 B.n497 B.n8 585
R274 B.n499 B.n498 585
R275 B.n500 B.n7 585
R276 B.n502 B.n501 585
R277 B.n503 B.n6 585
R278 B.n505 B.n504 585
R279 B.n506 B.n5 585
R280 B.n508 B.n507 585
R281 B.n509 B.n4 585
R282 B.n511 B.n510 585
R283 B.n512 B.n3 585
R284 B.n514 B.n513 585
R285 B.n515 B.n0 585
R286 B.n2 B.n1 585
R287 B.n134 B.n133 585
R288 B.n136 B.n135 585
R289 B.n137 B.n132 585
R290 B.n139 B.n138 585
R291 B.n140 B.n131 585
R292 B.n142 B.n141 585
R293 B.n143 B.n130 585
R294 B.n145 B.n144 585
R295 B.n146 B.n129 585
R296 B.n148 B.n147 585
R297 B.n149 B.n128 585
R298 B.n151 B.n150 585
R299 B.n150 B.n127 497.305
R300 B.n304 B.n303 497.305
R301 B.n346 B.n345 497.305
R302 B.n497 B.n496 497.305
R303 B.n517 B.n516 256.663
R304 B.n516 B.n515 235.042
R305 B.n516 B.n2 235.042
R306 B.n154 B.n127 163.367
R307 B.n155 B.n154 163.367
R308 B.n156 B.n155 163.367
R309 B.n156 B.n125 163.367
R310 B.n160 B.n125 163.367
R311 B.n161 B.n160 163.367
R312 B.n162 B.n161 163.367
R313 B.n162 B.n123 163.367
R314 B.n166 B.n123 163.367
R315 B.n167 B.n166 163.367
R316 B.n168 B.n167 163.367
R317 B.n168 B.n121 163.367
R318 B.n172 B.n121 163.367
R319 B.n173 B.n172 163.367
R320 B.n174 B.n173 163.367
R321 B.n174 B.n119 163.367
R322 B.n178 B.n119 163.367
R323 B.n179 B.n178 163.367
R324 B.n180 B.n179 163.367
R325 B.n180 B.n117 163.367
R326 B.n184 B.n117 163.367
R327 B.n185 B.n184 163.367
R328 B.n186 B.n185 163.367
R329 B.n186 B.n115 163.367
R330 B.n190 B.n115 163.367
R331 B.n191 B.n190 163.367
R332 B.n192 B.n191 163.367
R333 B.n192 B.n113 163.367
R334 B.n196 B.n113 163.367
R335 B.n197 B.n196 163.367
R336 B.n198 B.n197 163.367
R337 B.n198 B.n111 163.367
R338 B.n202 B.n111 163.367
R339 B.n203 B.n202 163.367
R340 B.n204 B.n203 163.367
R341 B.n204 B.n109 163.367
R342 B.n208 B.n109 163.367
R343 B.n209 B.n208 163.367
R344 B.n210 B.n209 163.367
R345 B.n210 B.n107 163.367
R346 B.n214 B.n107 163.367
R347 B.n215 B.n214 163.367
R348 B.n216 B.n215 163.367
R349 B.n216 B.n103 163.367
R350 B.n221 B.n103 163.367
R351 B.n222 B.n221 163.367
R352 B.n223 B.n222 163.367
R353 B.n223 B.n101 163.367
R354 B.n227 B.n101 163.367
R355 B.n228 B.n227 163.367
R356 B.n229 B.n228 163.367
R357 B.n229 B.n99 163.367
R358 B.n236 B.n99 163.367
R359 B.n237 B.n236 163.367
R360 B.n238 B.n237 163.367
R361 B.n238 B.n97 163.367
R362 B.n242 B.n97 163.367
R363 B.n243 B.n242 163.367
R364 B.n244 B.n243 163.367
R365 B.n244 B.n95 163.367
R366 B.n248 B.n95 163.367
R367 B.n249 B.n248 163.367
R368 B.n250 B.n249 163.367
R369 B.n250 B.n93 163.367
R370 B.n254 B.n93 163.367
R371 B.n255 B.n254 163.367
R372 B.n256 B.n255 163.367
R373 B.n256 B.n91 163.367
R374 B.n260 B.n91 163.367
R375 B.n261 B.n260 163.367
R376 B.n262 B.n261 163.367
R377 B.n262 B.n89 163.367
R378 B.n266 B.n89 163.367
R379 B.n267 B.n266 163.367
R380 B.n268 B.n267 163.367
R381 B.n268 B.n87 163.367
R382 B.n272 B.n87 163.367
R383 B.n273 B.n272 163.367
R384 B.n274 B.n273 163.367
R385 B.n274 B.n85 163.367
R386 B.n278 B.n85 163.367
R387 B.n279 B.n278 163.367
R388 B.n280 B.n279 163.367
R389 B.n280 B.n83 163.367
R390 B.n284 B.n83 163.367
R391 B.n285 B.n284 163.367
R392 B.n286 B.n285 163.367
R393 B.n286 B.n81 163.367
R394 B.n290 B.n81 163.367
R395 B.n291 B.n290 163.367
R396 B.n292 B.n291 163.367
R397 B.n292 B.n79 163.367
R398 B.n296 B.n79 163.367
R399 B.n297 B.n296 163.367
R400 B.n298 B.n297 163.367
R401 B.n298 B.n77 163.367
R402 B.n302 B.n77 163.367
R403 B.n303 B.n302 163.367
R404 B.n345 B.n344 163.367
R405 B.n344 B.n63 163.367
R406 B.n340 B.n63 163.367
R407 B.n340 B.n339 163.367
R408 B.n339 B.n338 163.367
R409 B.n338 B.n65 163.367
R410 B.n334 B.n65 163.367
R411 B.n334 B.n333 163.367
R412 B.n333 B.n332 163.367
R413 B.n332 B.n67 163.367
R414 B.n328 B.n67 163.367
R415 B.n328 B.n327 163.367
R416 B.n327 B.n326 163.367
R417 B.n326 B.n69 163.367
R418 B.n322 B.n69 163.367
R419 B.n322 B.n321 163.367
R420 B.n321 B.n320 163.367
R421 B.n320 B.n71 163.367
R422 B.n316 B.n71 163.367
R423 B.n316 B.n315 163.367
R424 B.n315 B.n314 163.367
R425 B.n314 B.n73 163.367
R426 B.n310 B.n73 163.367
R427 B.n310 B.n309 163.367
R428 B.n309 B.n308 163.367
R429 B.n308 B.n75 163.367
R430 B.n304 B.n75 163.367
R431 B.n496 B.n9 163.367
R432 B.n492 B.n9 163.367
R433 B.n492 B.n491 163.367
R434 B.n491 B.n490 163.367
R435 B.n490 B.n11 163.367
R436 B.n486 B.n11 163.367
R437 B.n486 B.n485 163.367
R438 B.n485 B.n484 163.367
R439 B.n484 B.n13 163.367
R440 B.n480 B.n13 163.367
R441 B.n480 B.n479 163.367
R442 B.n479 B.n478 163.367
R443 B.n478 B.n15 163.367
R444 B.n474 B.n15 163.367
R445 B.n474 B.n473 163.367
R446 B.n473 B.n472 163.367
R447 B.n472 B.n17 163.367
R448 B.n468 B.n17 163.367
R449 B.n468 B.n467 163.367
R450 B.n467 B.n466 163.367
R451 B.n466 B.n19 163.367
R452 B.n462 B.n19 163.367
R453 B.n462 B.n461 163.367
R454 B.n461 B.n460 163.367
R455 B.n460 B.n21 163.367
R456 B.n456 B.n21 163.367
R457 B.n456 B.n455 163.367
R458 B.n455 B.n454 163.367
R459 B.n454 B.n23 163.367
R460 B.n450 B.n23 163.367
R461 B.n450 B.n449 163.367
R462 B.n449 B.n448 163.367
R463 B.n448 B.n25 163.367
R464 B.n444 B.n25 163.367
R465 B.n444 B.n443 163.367
R466 B.n443 B.n442 163.367
R467 B.n442 B.n27 163.367
R468 B.n438 B.n27 163.367
R469 B.n438 B.n437 163.367
R470 B.n437 B.n436 163.367
R471 B.n436 B.n29 163.367
R472 B.n432 B.n29 163.367
R473 B.n432 B.n431 163.367
R474 B.n431 B.n430 163.367
R475 B.n430 B.n31 163.367
R476 B.n425 B.n31 163.367
R477 B.n425 B.n424 163.367
R478 B.n424 B.n423 163.367
R479 B.n423 B.n35 163.367
R480 B.n419 B.n35 163.367
R481 B.n419 B.n418 163.367
R482 B.n418 B.n417 163.367
R483 B.n417 B.n37 163.367
R484 B.n412 B.n37 163.367
R485 B.n412 B.n411 163.367
R486 B.n411 B.n410 163.367
R487 B.n410 B.n41 163.367
R488 B.n406 B.n41 163.367
R489 B.n406 B.n405 163.367
R490 B.n405 B.n404 163.367
R491 B.n404 B.n43 163.367
R492 B.n400 B.n43 163.367
R493 B.n400 B.n399 163.367
R494 B.n399 B.n398 163.367
R495 B.n398 B.n45 163.367
R496 B.n394 B.n45 163.367
R497 B.n394 B.n393 163.367
R498 B.n393 B.n392 163.367
R499 B.n392 B.n47 163.367
R500 B.n388 B.n47 163.367
R501 B.n388 B.n387 163.367
R502 B.n387 B.n386 163.367
R503 B.n386 B.n49 163.367
R504 B.n382 B.n49 163.367
R505 B.n382 B.n381 163.367
R506 B.n381 B.n380 163.367
R507 B.n380 B.n51 163.367
R508 B.n376 B.n51 163.367
R509 B.n376 B.n375 163.367
R510 B.n375 B.n374 163.367
R511 B.n374 B.n53 163.367
R512 B.n370 B.n53 163.367
R513 B.n370 B.n369 163.367
R514 B.n369 B.n368 163.367
R515 B.n368 B.n55 163.367
R516 B.n364 B.n55 163.367
R517 B.n364 B.n363 163.367
R518 B.n363 B.n362 163.367
R519 B.n362 B.n57 163.367
R520 B.n358 B.n57 163.367
R521 B.n358 B.n357 163.367
R522 B.n357 B.n356 163.367
R523 B.n356 B.n59 163.367
R524 B.n352 B.n59 163.367
R525 B.n352 B.n351 163.367
R526 B.n351 B.n350 163.367
R527 B.n350 B.n61 163.367
R528 B.n346 B.n61 163.367
R529 B.n498 B.n497 163.367
R530 B.n498 B.n7 163.367
R531 B.n502 B.n7 163.367
R532 B.n503 B.n502 163.367
R533 B.n504 B.n503 163.367
R534 B.n504 B.n5 163.367
R535 B.n508 B.n5 163.367
R536 B.n509 B.n508 163.367
R537 B.n510 B.n509 163.367
R538 B.n510 B.n3 163.367
R539 B.n514 B.n3 163.367
R540 B.n515 B.n514 163.367
R541 B.n133 B.n2 163.367
R542 B.n136 B.n133 163.367
R543 B.n137 B.n136 163.367
R544 B.n138 B.n137 163.367
R545 B.n138 B.n131 163.367
R546 B.n142 B.n131 163.367
R547 B.n143 B.n142 163.367
R548 B.n144 B.n143 163.367
R549 B.n144 B.n129 163.367
R550 B.n148 B.n129 163.367
R551 B.n149 B.n148 163.367
R552 B.n150 B.n149 163.367
R553 B.n232 B.t1 120.469
R554 B.n38 B.t11 120.469
R555 B.n104 B.t7 120.454
R556 B.n32 B.t5 120.454
R557 B.n233 B.t2 108.445
R558 B.n39 B.t10 108.445
R559 B.n105 B.t8 108.43
R560 B.n33 B.t4 108.43
R561 B.n219 B.n105 59.5399
R562 B.n234 B.n233 59.5399
R563 B.n414 B.n39 59.5399
R564 B.n428 B.n33 59.5399
R565 B.n495 B.n8 32.3127
R566 B.n347 B.n62 32.3127
R567 B.n305 B.n76 32.3127
R568 B.n152 B.n151 32.3127
R569 B B.n517 18.0485
R570 B.n105 B.n104 12.0247
R571 B.n233 B.n232 12.0247
R572 B.n39 B.n38 12.0247
R573 B.n33 B.n32 12.0247
R574 B.n499 B.n8 10.6151
R575 B.n500 B.n499 10.6151
R576 B.n501 B.n500 10.6151
R577 B.n501 B.n6 10.6151
R578 B.n505 B.n6 10.6151
R579 B.n506 B.n505 10.6151
R580 B.n507 B.n506 10.6151
R581 B.n507 B.n4 10.6151
R582 B.n511 B.n4 10.6151
R583 B.n512 B.n511 10.6151
R584 B.n513 B.n512 10.6151
R585 B.n513 B.n0 10.6151
R586 B.n495 B.n494 10.6151
R587 B.n494 B.n493 10.6151
R588 B.n493 B.n10 10.6151
R589 B.n489 B.n10 10.6151
R590 B.n489 B.n488 10.6151
R591 B.n488 B.n487 10.6151
R592 B.n487 B.n12 10.6151
R593 B.n483 B.n12 10.6151
R594 B.n483 B.n482 10.6151
R595 B.n482 B.n481 10.6151
R596 B.n481 B.n14 10.6151
R597 B.n477 B.n14 10.6151
R598 B.n477 B.n476 10.6151
R599 B.n476 B.n475 10.6151
R600 B.n475 B.n16 10.6151
R601 B.n471 B.n16 10.6151
R602 B.n471 B.n470 10.6151
R603 B.n470 B.n469 10.6151
R604 B.n469 B.n18 10.6151
R605 B.n465 B.n18 10.6151
R606 B.n465 B.n464 10.6151
R607 B.n464 B.n463 10.6151
R608 B.n463 B.n20 10.6151
R609 B.n459 B.n20 10.6151
R610 B.n459 B.n458 10.6151
R611 B.n458 B.n457 10.6151
R612 B.n457 B.n22 10.6151
R613 B.n453 B.n22 10.6151
R614 B.n453 B.n452 10.6151
R615 B.n452 B.n451 10.6151
R616 B.n451 B.n24 10.6151
R617 B.n447 B.n24 10.6151
R618 B.n447 B.n446 10.6151
R619 B.n446 B.n445 10.6151
R620 B.n445 B.n26 10.6151
R621 B.n441 B.n26 10.6151
R622 B.n441 B.n440 10.6151
R623 B.n440 B.n439 10.6151
R624 B.n439 B.n28 10.6151
R625 B.n435 B.n28 10.6151
R626 B.n435 B.n434 10.6151
R627 B.n434 B.n433 10.6151
R628 B.n433 B.n30 10.6151
R629 B.n429 B.n30 10.6151
R630 B.n427 B.n426 10.6151
R631 B.n426 B.n34 10.6151
R632 B.n422 B.n34 10.6151
R633 B.n422 B.n421 10.6151
R634 B.n421 B.n420 10.6151
R635 B.n420 B.n36 10.6151
R636 B.n416 B.n36 10.6151
R637 B.n416 B.n415 10.6151
R638 B.n413 B.n40 10.6151
R639 B.n409 B.n40 10.6151
R640 B.n409 B.n408 10.6151
R641 B.n408 B.n407 10.6151
R642 B.n407 B.n42 10.6151
R643 B.n403 B.n42 10.6151
R644 B.n403 B.n402 10.6151
R645 B.n402 B.n401 10.6151
R646 B.n401 B.n44 10.6151
R647 B.n397 B.n44 10.6151
R648 B.n397 B.n396 10.6151
R649 B.n396 B.n395 10.6151
R650 B.n395 B.n46 10.6151
R651 B.n391 B.n46 10.6151
R652 B.n391 B.n390 10.6151
R653 B.n390 B.n389 10.6151
R654 B.n389 B.n48 10.6151
R655 B.n385 B.n48 10.6151
R656 B.n385 B.n384 10.6151
R657 B.n384 B.n383 10.6151
R658 B.n383 B.n50 10.6151
R659 B.n379 B.n50 10.6151
R660 B.n379 B.n378 10.6151
R661 B.n378 B.n377 10.6151
R662 B.n377 B.n52 10.6151
R663 B.n373 B.n52 10.6151
R664 B.n373 B.n372 10.6151
R665 B.n372 B.n371 10.6151
R666 B.n371 B.n54 10.6151
R667 B.n367 B.n54 10.6151
R668 B.n367 B.n366 10.6151
R669 B.n366 B.n365 10.6151
R670 B.n365 B.n56 10.6151
R671 B.n361 B.n56 10.6151
R672 B.n361 B.n360 10.6151
R673 B.n360 B.n359 10.6151
R674 B.n359 B.n58 10.6151
R675 B.n355 B.n58 10.6151
R676 B.n355 B.n354 10.6151
R677 B.n354 B.n353 10.6151
R678 B.n353 B.n60 10.6151
R679 B.n349 B.n60 10.6151
R680 B.n349 B.n348 10.6151
R681 B.n348 B.n347 10.6151
R682 B.n343 B.n62 10.6151
R683 B.n343 B.n342 10.6151
R684 B.n342 B.n341 10.6151
R685 B.n341 B.n64 10.6151
R686 B.n337 B.n64 10.6151
R687 B.n337 B.n336 10.6151
R688 B.n336 B.n335 10.6151
R689 B.n335 B.n66 10.6151
R690 B.n331 B.n66 10.6151
R691 B.n331 B.n330 10.6151
R692 B.n330 B.n329 10.6151
R693 B.n329 B.n68 10.6151
R694 B.n325 B.n68 10.6151
R695 B.n325 B.n324 10.6151
R696 B.n324 B.n323 10.6151
R697 B.n323 B.n70 10.6151
R698 B.n319 B.n70 10.6151
R699 B.n319 B.n318 10.6151
R700 B.n318 B.n317 10.6151
R701 B.n317 B.n72 10.6151
R702 B.n313 B.n72 10.6151
R703 B.n313 B.n312 10.6151
R704 B.n312 B.n311 10.6151
R705 B.n311 B.n74 10.6151
R706 B.n307 B.n74 10.6151
R707 B.n307 B.n306 10.6151
R708 B.n306 B.n305 10.6151
R709 B.n134 B.n1 10.6151
R710 B.n135 B.n134 10.6151
R711 B.n135 B.n132 10.6151
R712 B.n139 B.n132 10.6151
R713 B.n140 B.n139 10.6151
R714 B.n141 B.n140 10.6151
R715 B.n141 B.n130 10.6151
R716 B.n145 B.n130 10.6151
R717 B.n146 B.n145 10.6151
R718 B.n147 B.n146 10.6151
R719 B.n147 B.n128 10.6151
R720 B.n151 B.n128 10.6151
R721 B.n153 B.n152 10.6151
R722 B.n153 B.n126 10.6151
R723 B.n157 B.n126 10.6151
R724 B.n158 B.n157 10.6151
R725 B.n159 B.n158 10.6151
R726 B.n159 B.n124 10.6151
R727 B.n163 B.n124 10.6151
R728 B.n164 B.n163 10.6151
R729 B.n165 B.n164 10.6151
R730 B.n165 B.n122 10.6151
R731 B.n169 B.n122 10.6151
R732 B.n170 B.n169 10.6151
R733 B.n171 B.n170 10.6151
R734 B.n171 B.n120 10.6151
R735 B.n175 B.n120 10.6151
R736 B.n176 B.n175 10.6151
R737 B.n177 B.n176 10.6151
R738 B.n177 B.n118 10.6151
R739 B.n181 B.n118 10.6151
R740 B.n182 B.n181 10.6151
R741 B.n183 B.n182 10.6151
R742 B.n183 B.n116 10.6151
R743 B.n187 B.n116 10.6151
R744 B.n188 B.n187 10.6151
R745 B.n189 B.n188 10.6151
R746 B.n189 B.n114 10.6151
R747 B.n193 B.n114 10.6151
R748 B.n194 B.n193 10.6151
R749 B.n195 B.n194 10.6151
R750 B.n195 B.n112 10.6151
R751 B.n199 B.n112 10.6151
R752 B.n200 B.n199 10.6151
R753 B.n201 B.n200 10.6151
R754 B.n201 B.n110 10.6151
R755 B.n205 B.n110 10.6151
R756 B.n206 B.n205 10.6151
R757 B.n207 B.n206 10.6151
R758 B.n207 B.n108 10.6151
R759 B.n211 B.n108 10.6151
R760 B.n212 B.n211 10.6151
R761 B.n213 B.n212 10.6151
R762 B.n213 B.n106 10.6151
R763 B.n217 B.n106 10.6151
R764 B.n218 B.n217 10.6151
R765 B.n220 B.n102 10.6151
R766 B.n224 B.n102 10.6151
R767 B.n225 B.n224 10.6151
R768 B.n226 B.n225 10.6151
R769 B.n226 B.n100 10.6151
R770 B.n230 B.n100 10.6151
R771 B.n231 B.n230 10.6151
R772 B.n235 B.n231 10.6151
R773 B.n239 B.n98 10.6151
R774 B.n240 B.n239 10.6151
R775 B.n241 B.n240 10.6151
R776 B.n241 B.n96 10.6151
R777 B.n245 B.n96 10.6151
R778 B.n246 B.n245 10.6151
R779 B.n247 B.n246 10.6151
R780 B.n247 B.n94 10.6151
R781 B.n251 B.n94 10.6151
R782 B.n252 B.n251 10.6151
R783 B.n253 B.n252 10.6151
R784 B.n253 B.n92 10.6151
R785 B.n257 B.n92 10.6151
R786 B.n258 B.n257 10.6151
R787 B.n259 B.n258 10.6151
R788 B.n259 B.n90 10.6151
R789 B.n263 B.n90 10.6151
R790 B.n264 B.n263 10.6151
R791 B.n265 B.n264 10.6151
R792 B.n265 B.n88 10.6151
R793 B.n269 B.n88 10.6151
R794 B.n270 B.n269 10.6151
R795 B.n271 B.n270 10.6151
R796 B.n271 B.n86 10.6151
R797 B.n275 B.n86 10.6151
R798 B.n276 B.n275 10.6151
R799 B.n277 B.n276 10.6151
R800 B.n277 B.n84 10.6151
R801 B.n281 B.n84 10.6151
R802 B.n282 B.n281 10.6151
R803 B.n283 B.n282 10.6151
R804 B.n283 B.n82 10.6151
R805 B.n287 B.n82 10.6151
R806 B.n288 B.n287 10.6151
R807 B.n289 B.n288 10.6151
R808 B.n289 B.n80 10.6151
R809 B.n293 B.n80 10.6151
R810 B.n294 B.n293 10.6151
R811 B.n295 B.n294 10.6151
R812 B.n295 B.n78 10.6151
R813 B.n299 B.n78 10.6151
R814 B.n300 B.n299 10.6151
R815 B.n301 B.n300 10.6151
R816 B.n301 B.n76 10.6151
R817 B.n517 B.n0 8.11757
R818 B.n517 B.n1 8.11757
R819 B.n428 B.n427 7.18099
R820 B.n415 B.n414 7.18099
R821 B.n220 B.n219 7.18099
R822 B.n235 B.n234 7.18099
R823 B.n429 B.n428 3.43465
R824 B.n414 B.n413 3.43465
R825 B.n219 B.n218 3.43465
R826 B.n234 B.n98 3.43465
C0 VDD2 VDD1 0.476453f
C1 VN VTAIL 1.61723f
C2 VTAIL VDD2 10.2891f
C3 VN w_n1342_n3572# 1.86538f
C4 B VP 0.945365f
C5 w_n1342_n3572# VDD2 0.999054f
C6 VP VDD1 2.293f
C7 B VDD1 0.88026f
C8 VTAIL VP 1.63133f
C9 VN VDD2 2.19275f
C10 VTAIL B 3.75822f
C11 w_n1342_n3572# VP 2.03205f
C12 VTAIL VDD1 10.250299f
C13 w_n1342_n3572# B 6.70722f
C14 w_n1342_n3572# VDD1 0.992438f
C15 VN VP 4.70433f
C16 VP VDD2 0.248789f
C17 VTAIL w_n1342_n3572# 4.54196f
C18 VN B 0.679522f
C19 B VDD2 0.896141f
C20 VN VDD1 0.148385f
C21 VDD2 VSUBS 0.654157f
C22 VDD1 VSUBS 5.680971f
C23 VTAIL VSUBS 0.774858f
C24 VN VSUBS 5.14405f
C25 VP VSUBS 1.125757f
C26 B VSUBS 2.355407f
C27 w_n1342_n3572# VSUBS 58.924496f
C28 B.n0 VSUBS 0.007681f
C29 B.n1 VSUBS 0.007681f
C30 B.n2 VSUBS 0.01136f
C31 B.n3 VSUBS 0.008705f
C32 B.n4 VSUBS 0.008705f
C33 B.n5 VSUBS 0.008705f
C34 B.n6 VSUBS 0.008705f
C35 B.n7 VSUBS 0.008705f
C36 B.n8 VSUBS 0.019581f
C37 B.n9 VSUBS 0.008705f
C38 B.n10 VSUBS 0.008705f
C39 B.n11 VSUBS 0.008705f
C40 B.n12 VSUBS 0.008705f
C41 B.n13 VSUBS 0.008705f
C42 B.n14 VSUBS 0.008705f
C43 B.n15 VSUBS 0.008705f
C44 B.n16 VSUBS 0.008705f
C45 B.n17 VSUBS 0.008705f
C46 B.n18 VSUBS 0.008705f
C47 B.n19 VSUBS 0.008705f
C48 B.n20 VSUBS 0.008705f
C49 B.n21 VSUBS 0.008705f
C50 B.n22 VSUBS 0.008705f
C51 B.n23 VSUBS 0.008705f
C52 B.n24 VSUBS 0.008705f
C53 B.n25 VSUBS 0.008705f
C54 B.n26 VSUBS 0.008705f
C55 B.n27 VSUBS 0.008705f
C56 B.n28 VSUBS 0.008705f
C57 B.n29 VSUBS 0.008705f
C58 B.n30 VSUBS 0.008705f
C59 B.n31 VSUBS 0.008705f
C60 B.t4 VSUBS 0.531209f
C61 B.t5 VSUBS 0.537704f
C62 B.t3 VSUBS 0.183433f
C63 B.n32 VSUBS 0.123763f
C64 B.n33 VSUBS 0.077484f
C65 B.n34 VSUBS 0.008705f
C66 B.n35 VSUBS 0.008705f
C67 B.n36 VSUBS 0.008705f
C68 B.n37 VSUBS 0.008705f
C69 B.t10 VSUBS 0.531197f
C70 B.t11 VSUBS 0.537693f
C71 B.t9 VSUBS 0.183433f
C72 B.n38 VSUBS 0.123775f
C73 B.n39 VSUBS 0.077496f
C74 B.n40 VSUBS 0.008705f
C75 B.n41 VSUBS 0.008705f
C76 B.n42 VSUBS 0.008705f
C77 B.n43 VSUBS 0.008705f
C78 B.n44 VSUBS 0.008705f
C79 B.n45 VSUBS 0.008705f
C80 B.n46 VSUBS 0.008705f
C81 B.n47 VSUBS 0.008705f
C82 B.n48 VSUBS 0.008705f
C83 B.n49 VSUBS 0.008705f
C84 B.n50 VSUBS 0.008705f
C85 B.n51 VSUBS 0.008705f
C86 B.n52 VSUBS 0.008705f
C87 B.n53 VSUBS 0.008705f
C88 B.n54 VSUBS 0.008705f
C89 B.n55 VSUBS 0.008705f
C90 B.n56 VSUBS 0.008705f
C91 B.n57 VSUBS 0.008705f
C92 B.n58 VSUBS 0.008705f
C93 B.n59 VSUBS 0.008705f
C94 B.n60 VSUBS 0.008705f
C95 B.n61 VSUBS 0.008705f
C96 B.n62 VSUBS 0.019581f
C97 B.n63 VSUBS 0.008705f
C98 B.n64 VSUBS 0.008705f
C99 B.n65 VSUBS 0.008705f
C100 B.n66 VSUBS 0.008705f
C101 B.n67 VSUBS 0.008705f
C102 B.n68 VSUBS 0.008705f
C103 B.n69 VSUBS 0.008705f
C104 B.n70 VSUBS 0.008705f
C105 B.n71 VSUBS 0.008705f
C106 B.n72 VSUBS 0.008705f
C107 B.n73 VSUBS 0.008705f
C108 B.n74 VSUBS 0.008705f
C109 B.n75 VSUBS 0.008705f
C110 B.n76 VSUBS 0.019834f
C111 B.n77 VSUBS 0.008705f
C112 B.n78 VSUBS 0.008705f
C113 B.n79 VSUBS 0.008705f
C114 B.n80 VSUBS 0.008705f
C115 B.n81 VSUBS 0.008705f
C116 B.n82 VSUBS 0.008705f
C117 B.n83 VSUBS 0.008705f
C118 B.n84 VSUBS 0.008705f
C119 B.n85 VSUBS 0.008705f
C120 B.n86 VSUBS 0.008705f
C121 B.n87 VSUBS 0.008705f
C122 B.n88 VSUBS 0.008705f
C123 B.n89 VSUBS 0.008705f
C124 B.n90 VSUBS 0.008705f
C125 B.n91 VSUBS 0.008705f
C126 B.n92 VSUBS 0.008705f
C127 B.n93 VSUBS 0.008705f
C128 B.n94 VSUBS 0.008705f
C129 B.n95 VSUBS 0.008705f
C130 B.n96 VSUBS 0.008705f
C131 B.n97 VSUBS 0.008705f
C132 B.n98 VSUBS 0.005761f
C133 B.n99 VSUBS 0.008705f
C134 B.n100 VSUBS 0.008705f
C135 B.n101 VSUBS 0.008705f
C136 B.n102 VSUBS 0.008705f
C137 B.n103 VSUBS 0.008705f
C138 B.t8 VSUBS 0.531209f
C139 B.t7 VSUBS 0.537704f
C140 B.t6 VSUBS 0.183433f
C141 B.n104 VSUBS 0.123763f
C142 B.n105 VSUBS 0.077484f
C143 B.n106 VSUBS 0.008705f
C144 B.n107 VSUBS 0.008705f
C145 B.n108 VSUBS 0.008705f
C146 B.n109 VSUBS 0.008705f
C147 B.n110 VSUBS 0.008705f
C148 B.n111 VSUBS 0.008705f
C149 B.n112 VSUBS 0.008705f
C150 B.n113 VSUBS 0.008705f
C151 B.n114 VSUBS 0.008705f
C152 B.n115 VSUBS 0.008705f
C153 B.n116 VSUBS 0.008705f
C154 B.n117 VSUBS 0.008705f
C155 B.n118 VSUBS 0.008705f
C156 B.n119 VSUBS 0.008705f
C157 B.n120 VSUBS 0.008705f
C158 B.n121 VSUBS 0.008705f
C159 B.n122 VSUBS 0.008705f
C160 B.n123 VSUBS 0.008705f
C161 B.n124 VSUBS 0.008705f
C162 B.n125 VSUBS 0.008705f
C163 B.n126 VSUBS 0.008705f
C164 B.n127 VSUBS 0.020874f
C165 B.n128 VSUBS 0.008705f
C166 B.n129 VSUBS 0.008705f
C167 B.n130 VSUBS 0.008705f
C168 B.n131 VSUBS 0.008705f
C169 B.n132 VSUBS 0.008705f
C170 B.n133 VSUBS 0.008705f
C171 B.n134 VSUBS 0.008705f
C172 B.n135 VSUBS 0.008705f
C173 B.n136 VSUBS 0.008705f
C174 B.n137 VSUBS 0.008705f
C175 B.n138 VSUBS 0.008705f
C176 B.n139 VSUBS 0.008705f
C177 B.n140 VSUBS 0.008705f
C178 B.n141 VSUBS 0.008705f
C179 B.n142 VSUBS 0.008705f
C180 B.n143 VSUBS 0.008705f
C181 B.n144 VSUBS 0.008705f
C182 B.n145 VSUBS 0.008705f
C183 B.n146 VSUBS 0.008705f
C184 B.n147 VSUBS 0.008705f
C185 B.n148 VSUBS 0.008705f
C186 B.n149 VSUBS 0.008705f
C187 B.n150 VSUBS 0.019581f
C188 B.n151 VSUBS 0.019581f
C189 B.n152 VSUBS 0.020874f
C190 B.n153 VSUBS 0.008705f
C191 B.n154 VSUBS 0.008705f
C192 B.n155 VSUBS 0.008705f
C193 B.n156 VSUBS 0.008705f
C194 B.n157 VSUBS 0.008705f
C195 B.n158 VSUBS 0.008705f
C196 B.n159 VSUBS 0.008705f
C197 B.n160 VSUBS 0.008705f
C198 B.n161 VSUBS 0.008705f
C199 B.n162 VSUBS 0.008705f
C200 B.n163 VSUBS 0.008705f
C201 B.n164 VSUBS 0.008705f
C202 B.n165 VSUBS 0.008705f
C203 B.n166 VSUBS 0.008705f
C204 B.n167 VSUBS 0.008705f
C205 B.n168 VSUBS 0.008705f
C206 B.n169 VSUBS 0.008705f
C207 B.n170 VSUBS 0.008705f
C208 B.n171 VSUBS 0.008705f
C209 B.n172 VSUBS 0.008705f
C210 B.n173 VSUBS 0.008705f
C211 B.n174 VSUBS 0.008705f
C212 B.n175 VSUBS 0.008705f
C213 B.n176 VSUBS 0.008705f
C214 B.n177 VSUBS 0.008705f
C215 B.n178 VSUBS 0.008705f
C216 B.n179 VSUBS 0.008705f
C217 B.n180 VSUBS 0.008705f
C218 B.n181 VSUBS 0.008705f
C219 B.n182 VSUBS 0.008705f
C220 B.n183 VSUBS 0.008705f
C221 B.n184 VSUBS 0.008705f
C222 B.n185 VSUBS 0.008705f
C223 B.n186 VSUBS 0.008705f
C224 B.n187 VSUBS 0.008705f
C225 B.n188 VSUBS 0.008705f
C226 B.n189 VSUBS 0.008705f
C227 B.n190 VSUBS 0.008705f
C228 B.n191 VSUBS 0.008705f
C229 B.n192 VSUBS 0.008705f
C230 B.n193 VSUBS 0.008705f
C231 B.n194 VSUBS 0.008705f
C232 B.n195 VSUBS 0.008705f
C233 B.n196 VSUBS 0.008705f
C234 B.n197 VSUBS 0.008705f
C235 B.n198 VSUBS 0.008705f
C236 B.n199 VSUBS 0.008705f
C237 B.n200 VSUBS 0.008705f
C238 B.n201 VSUBS 0.008705f
C239 B.n202 VSUBS 0.008705f
C240 B.n203 VSUBS 0.008705f
C241 B.n204 VSUBS 0.008705f
C242 B.n205 VSUBS 0.008705f
C243 B.n206 VSUBS 0.008705f
C244 B.n207 VSUBS 0.008705f
C245 B.n208 VSUBS 0.008705f
C246 B.n209 VSUBS 0.008705f
C247 B.n210 VSUBS 0.008705f
C248 B.n211 VSUBS 0.008705f
C249 B.n212 VSUBS 0.008705f
C250 B.n213 VSUBS 0.008705f
C251 B.n214 VSUBS 0.008705f
C252 B.n215 VSUBS 0.008705f
C253 B.n216 VSUBS 0.008705f
C254 B.n217 VSUBS 0.008705f
C255 B.n218 VSUBS 0.005761f
C256 B.n219 VSUBS 0.02017f
C257 B.n220 VSUBS 0.007297f
C258 B.n221 VSUBS 0.008705f
C259 B.n222 VSUBS 0.008705f
C260 B.n223 VSUBS 0.008705f
C261 B.n224 VSUBS 0.008705f
C262 B.n225 VSUBS 0.008705f
C263 B.n226 VSUBS 0.008705f
C264 B.n227 VSUBS 0.008705f
C265 B.n228 VSUBS 0.008705f
C266 B.n229 VSUBS 0.008705f
C267 B.n230 VSUBS 0.008705f
C268 B.n231 VSUBS 0.008705f
C269 B.t2 VSUBS 0.531197f
C270 B.t1 VSUBS 0.537693f
C271 B.t0 VSUBS 0.183433f
C272 B.n232 VSUBS 0.123775f
C273 B.n233 VSUBS 0.077496f
C274 B.n234 VSUBS 0.02017f
C275 B.n235 VSUBS 0.007297f
C276 B.n236 VSUBS 0.008705f
C277 B.n237 VSUBS 0.008705f
C278 B.n238 VSUBS 0.008705f
C279 B.n239 VSUBS 0.008705f
C280 B.n240 VSUBS 0.008705f
C281 B.n241 VSUBS 0.008705f
C282 B.n242 VSUBS 0.008705f
C283 B.n243 VSUBS 0.008705f
C284 B.n244 VSUBS 0.008705f
C285 B.n245 VSUBS 0.008705f
C286 B.n246 VSUBS 0.008705f
C287 B.n247 VSUBS 0.008705f
C288 B.n248 VSUBS 0.008705f
C289 B.n249 VSUBS 0.008705f
C290 B.n250 VSUBS 0.008705f
C291 B.n251 VSUBS 0.008705f
C292 B.n252 VSUBS 0.008705f
C293 B.n253 VSUBS 0.008705f
C294 B.n254 VSUBS 0.008705f
C295 B.n255 VSUBS 0.008705f
C296 B.n256 VSUBS 0.008705f
C297 B.n257 VSUBS 0.008705f
C298 B.n258 VSUBS 0.008705f
C299 B.n259 VSUBS 0.008705f
C300 B.n260 VSUBS 0.008705f
C301 B.n261 VSUBS 0.008705f
C302 B.n262 VSUBS 0.008705f
C303 B.n263 VSUBS 0.008705f
C304 B.n264 VSUBS 0.008705f
C305 B.n265 VSUBS 0.008705f
C306 B.n266 VSUBS 0.008705f
C307 B.n267 VSUBS 0.008705f
C308 B.n268 VSUBS 0.008705f
C309 B.n269 VSUBS 0.008705f
C310 B.n270 VSUBS 0.008705f
C311 B.n271 VSUBS 0.008705f
C312 B.n272 VSUBS 0.008705f
C313 B.n273 VSUBS 0.008705f
C314 B.n274 VSUBS 0.008705f
C315 B.n275 VSUBS 0.008705f
C316 B.n276 VSUBS 0.008705f
C317 B.n277 VSUBS 0.008705f
C318 B.n278 VSUBS 0.008705f
C319 B.n279 VSUBS 0.008705f
C320 B.n280 VSUBS 0.008705f
C321 B.n281 VSUBS 0.008705f
C322 B.n282 VSUBS 0.008705f
C323 B.n283 VSUBS 0.008705f
C324 B.n284 VSUBS 0.008705f
C325 B.n285 VSUBS 0.008705f
C326 B.n286 VSUBS 0.008705f
C327 B.n287 VSUBS 0.008705f
C328 B.n288 VSUBS 0.008705f
C329 B.n289 VSUBS 0.008705f
C330 B.n290 VSUBS 0.008705f
C331 B.n291 VSUBS 0.008705f
C332 B.n292 VSUBS 0.008705f
C333 B.n293 VSUBS 0.008705f
C334 B.n294 VSUBS 0.008705f
C335 B.n295 VSUBS 0.008705f
C336 B.n296 VSUBS 0.008705f
C337 B.n297 VSUBS 0.008705f
C338 B.n298 VSUBS 0.008705f
C339 B.n299 VSUBS 0.008705f
C340 B.n300 VSUBS 0.008705f
C341 B.n301 VSUBS 0.008705f
C342 B.n302 VSUBS 0.008705f
C343 B.n303 VSUBS 0.020874f
C344 B.n304 VSUBS 0.019581f
C345 B.n305 VSUBS 0.020621f
C346 B.n306 VSUBS 0.008705f
C347 B.n307 VSUBS 0.008705f
C348 B.n308 VSUBS 0.008705f
C349 B.n309 VSUBS 0.008705f
C350 B.n310 VSUBS 0.008705f
C351 B.n311 VSUBS 0.008705f
C352 B.n312 VSUBS 0.008705f
C353 B.n313 VSUBS 0.008705f
C354 B.n314 VSUBS 0.008705f
C355 B.n315 VSUBS 0.008705f
C356 B.n316 VSUBS 0.008705f
C357 B.n317 VSUBS 0.008705f
C358 B.n318 VSUBS 0.008705f
C359 B.n319 VSUBS 0.008705f
C360 B.n320 VSUBS 0.008705f
C361 B.n321 VSUBS 0.008705f
C362 B.n322 VSUBS 0.008705f
C363 B.n323 VSUBS 0.008705f
C364 B.n324 VSUBS 0.008705f
C365 B.n325 VSUBS 0.008705f
C366 B.n326 VSUBS 0.008705f
C367 B.n327 VSUBS 0.008705f
C368 B.n328 VSUBS 0.008705f
C369 B.n329 VSUBS 0.008705f
C370 B.n330 VSUBS 0.008705f
C371 B.n331 VSUBS 0.008705f
C372 B.n332 VSUBS 0.008705f
C373 B.n333 VSUBS 0.008705f
C374 B.n334 VSUBS 0.008705f
C375 B.n335 VSUBS 0.008705f
C376 B.n336 VSUBS 0.008705f
C377 B.n337 VSUBS 0.008705f
C378 B.n338 VSUBS 0.008705f
C379 B.n339 VSUBS 0.008705f
C380 B.n340 VSUBS 0.008705f
C381 B.n341 VSUBS 0.008705f
C382 B.n342 VSUBS 0.008705f
C383 B.n343 VSUBS 0.008705f
C384 B.n344 VSUBS 0.008705f
C385 B.n345 VSUBS 0.019581f
C386 B.n346 VSUBS 0.020874f
C387 B.n347 VSUBS 0.020874f
C388 B.n348 VSUBS 0.008705f
C389 B.n349 VSUBS 0.008705f
C390 B.n350 VSUBS 0.008705f
C391 B.n351 VSUBS 0.008705f
C392 B.n352 VSUBS 0.008705f
C393 B.n353 VSUBS 0.008705f
C394 B.n354 VSUBS 0.008705f
C395 B.n355 VSUBS 0.008705f
C396 B.n356 VSUBS 0.008705f
C397 B.n357 VSUBS 0.008705f
C398 B.n358 VSUBS 0.008705f
C399 B.n359 VSUBS 0.008705f
C400 B.n360 VSUBS 0.008705f
C401 B.n361 VSUBS 0.008705f
C402 B.n362 VSUBS 0.008705f
C403 B.n363 VSUBS 0.008705f
C404 B.n364 VSUBS 0.008705f
C405 B.n365 VSUBS 0.008705f
C406 B.n366 VSUBS 0.008705f
C407 B.n367 VSUBS 0.008705f
C408 B.n368 VSUBS 0.008705f
C409 B.n369 VSUBS 0.008705f
C410 B.n370 VSUBS 0.008705f
C411 B.n371 VSUBS 0.008705f
C412 B.n372 VSUBS 0.008705f
C413 B.n373 VSUBS 0.008705f
C414 B.n374 VSUBS 0.008705f
C415 B.n375 VSUBS 0.008705f
C416 B.n376 VSUBS 0.008705f
C417 B.n377 VSUBS 0.008705f
C418 B.n378 VSUBS 0.008705f
C419 B.n379 VSUBS 0.008705f
C420 B.n380 VSUBS 0.008705f
C421 B.n381 VSUBS 0.008705f
C422 B.n382 VSUBS 0.008705f
C423 B.n383 VSUBS 0.008705f
C424 B.n384 VSUBS 0.008705f
C425 B.n385 VSUBS 0.008705f
C426 B.n386 VSUBS 0.008705f
C427 B.n387 VSUBS 0.008705f
C428 B.n388 VSUBS 0.008705f
C429 B.n389 VSUBS 0.008705f
C430 B.n390 VSUBS 0.008705f
C431 B.n391 VSUBS 0.008705f
C432 B.n392 VSUBS 0.008705f
C433 B.n393 VSUBS 0.008705f
C434 B.n394 VSUBS 0.008705f
C435 B.n395 VSUBS 0.008705f
C436 B.n396 VSUBS 0.008705f
C437 B.n397 VSUBS 0.008705f
C438 B.n398 VSUBS 0.008705f
C439 B.n399 VSUBS 0.008705f
C440 B.n400 VSUBS 0.008705f
C441 B.n401 VSUBS 0.008705f
C442 B.n402 VSUBS 0.008705f
C443 B.n403 VSUBS 0.008705f
C444 B.n404 VSUBS 0.008705f
C445 B.n405 VSUBS 0.008705f
C446 B.n406 VSUBS 0.008705f
C447 B.n407 VSUBS 0.008705f
C448 B.n408 VSUBS 0.008705f
C449 B.n409 VSUBS 0.008705f
C450 B.n410 VSUBS 0.008705f
C451 B.n411 VSUBS 0.008705f
C452 B.n412 VSUBS 0.008705f
C453 B.n413 VSUBS 0.005761f
C454 B.n414 VSUBS 0.02017f
C455 B.n415 VSUBS 0.007297f
C456 B.n416 VSUBS 0.008705f
C457 B.n417 VSUBS 0.008705f
C458 B.n418 VSUBS 0.008705f
C459 B.n419 VSUBS 0.008705f
C460 B.n420 VSUBS 0.008705f
C461 B.n421 VSUBS 0.008705f
C462 B.n422 VSUBS 0.008705f
C463 B.n423 VSUBS 0.008705f
C464 B.n424 VSUBS 0.008705f
C465 B.n425 VSUBS 0.008705f
C466 B.n426 VSUBS 0.008705f
C467 B.n427 VSUBS 0.007297f
C468 B.n428 VSUBS 0.02017f
C469 B.n429 VSUBS 0.005761f
C470 B.n430 VSUBS 0.008705f
C471 B.n431 VSUBS 0.008705f
C472 B.n432 VSUBS 0.008705f
C473 B.n433 VSUBS 0.008705f
C474 B.n434 VSUBS 0.008705f
C475 B.n435 VSUBS 0.008705f
C476 B.n436 VSUBS 0.008705f
C477 B.n437 VSUBS 0.008705f
C478 B.n438 VSUBS 0.008705f
C479 B.n439 VSUBS 0.008705f
C480 B.n440 VSUBS 0.008705f
C481 B.n441 VSUBS 0.008705f
C482 B.n442 VSUBS 0.008705f
C483 B.n443 VSUBS 0.008705f
C484 B.n444 VSUBS 0.008705f
C485 B.n445 VSUBS 0.008705f
C486 B.n446 VSUBS 0.008705f
C487 B.n447 VSUBS 0.008705f
C488 B.n448 VSUBS 0.008705f
C489 B.n449 VSUBS 0.008705f
C490 B.n450 VSUBS 0.008705f
C491 B.n451 VSUBS 0.008705f
C492 B.n452 VSUBS 0.008705f
C493 B.n453 VSUBS 0.008705f
C494 B.n454 VSUBS 0.008705f
C495 B.n455 VSUBS 0.008705f
C496 B.n456 VSUBS 0.008705f
C497 B.n457 VSUBS 0.008705f
C498 B.n458 VSUBS 0.008705f
C499 B.n459 VSUBS 0.008705f
C500 B.n460 VSUBS 0.008705f
C501 B.n461 VSUBS 0.008705f
C502 B.n462 VSUBS 0.008705f
C503 B.n463 VSUBS 0.008705f
C504 B.n464 VSUBS 0.008705f
C505 B.n465 VSUBS 0.008705f
C506 B.n466 VSUBS 0.008705f
C507 B.n467 VSUBS 0.008705f
C508 B.n468 VSUBS 0.008705f
C509 B.n469 VSUBS 0.008705f
C510 B.n470 VSUBS 0.008705f
C511 B.n471 VSUBS 0.008705f
C512 B.n472 VSUBS 0.008705f
C513 B.n473 VSUBS 0.008705f
C514 B.n474 VSUBS 0.008705f
C515 B.n475 VSUBS 0.008705f
C516 B.n476 VSUBS 0.008705f
C517 B.n477 VSUBS 0.008705f
C518 B.n478 VSUBS 0.008705f
C519 B.n479 VSUBS 0.008705f
C520 B.n480 VSUBS 0.008705f
C521 B.n481 VSUBS 0.008705f
C522 B.n482 VSUBS 0.008705f
C523 B.n483 VSUBS 0.008705f
C524 B.n484 VSUBS 0.008705f
C525 B.n485 VSUBS 0.008705f
C526 B.n486 VSUBS 0.008705f
C527 B.n487 VSUBS 0.008705f
C528 B.n488 VSUBS 0.008705f
C529 B.n489 VSUBS 0.008705f
C530 B.n490 VSUBS 0.008705f
C531 B.n491 VSUBS 0.008705f
C532 B.n492 VSUBS 0.008705f
C533 B.n493 VSUBS 0.008705f
C534 B.n494 VSUBS 0.008705f
C535 B.n495 VSUBS 0.020874f
C536 B.n496 VSUBS 0.020874f
C537 B.n497 VSUBS 0.019581f
C538 B.n498 VSUBS 0.008705f
C539 B.n499 VSUBS 0.008705f
C540 B.n500 VSUBS 0.008705f
C541 B.n501 VSUBS 0.008705f
C542 B.n502 VSUBS 0.008705f
C543 B.n503 VSUBS 0.008705f
C544 B.n504 VSUBS 0.008705f
C545 B.n505 VSUBS 0.008705f
C546 B.n506 VSUBS 0.008705f
C547 B.n507 VSUBS 0.008705f
C548 B.n508 VSUBS 0.008705f
C549 B.n509 VSUBS 0.008705f
C550 B.n510 VSUBS 0.008705f
C551 B.n511 VSUBS 0.008705f
C552 B.n512 VSUBS 0.008705f
C553 B.n513 VSUBS 0.008705f
C554 B.n514 VSUBS 0.008705f
C555 B.n515 VSUBS 0.01136f
C556 B.n516 VSUBS 0.012101f
C557 B.n517 VSUBS 0.024065f
C558 VDD2.t3 VSUBS 0.344934f
C559 VDD2.t2 VSUBS 0.344934f
C560 VDD2.n0 VSUBS 3.51386f
C561 VDD2.t1 VSUBS 0.344934f
C562 VDD2.t0 VSUBS 0.344934f
C563 VDD2.n1 VSUBS 2.75524f
C564 VDD2.n2 VSUBS 4.78611f
C565 VN.t0 VSUBS 0.535423f
C566 VN.t1 VSUBS 0.535423f
C567 VN.n0 VSUBS 0.425384f
C568 VN.t2 VSUBS 0.535423f
C569 VN.t3 VSUBS 0.535423f
C570 VN.n1 VSUBS 0.811652f
C571 VDD1.t0 VSUBS 0.344278f
C572 VDD1.t3 VSUBS 0.344278f
C573 VDD1.n0 VSUBS 2.75053f
C574 VDD1.t1 VSUBS 0.344278f
C575 VDD1.t2 VSUBS 0.344278f
C576 VDD1.n1 VSUBS 3.53691f
C577 VTAIL.t7 VSUBS 2.35338f
C578 VTAIL.n0 VSUBS 0.661881f
C579 VTAIL.t4 VSUBS 2.35338f
C580 VTAIL.n1 VSUBS 0.677564f
C581 VTAIL.t5 VSUBS 2.35338f
C582 VTAIL.n2 VSUBS 1.84067f
C583 VTAIL.t1 VSUBS 2.3534f
C584 VTAIL.n3 VSUBS 1.84065f
C585 VTAIL.t0 VSUBS 2.3534f
C586 VTAIL.n4 VSUBS 0.677544f
C587 VTAIL.t6 VSUBS 2.3534f
C588 VTAIL.n5 VSUBS 0.677544f
C589 VTAIL.t3 VSUBS 2.35338f
C590 VTAIL.n6 VSUBS 1.84067f
C591 VTAIL.t2 VSUBS 2.35338f
C592 VTAIL.n7 VSUBS 1.81626f
C593 VP.t3 VSUBS 0.705502f
C594 VP.t0 VSUBS 0.705502f
C595 VP.n0 VSUBS 1.05708f
C596 VP.t2 VSUBS 0.705502f
C597 VP.t1 VSUBS 0.705502f
C598 VP.n1 VSUBS 0.560487f
C599 VP.n2 VSUBS 4.52921f
.ends

