* NGSPICE file created from diff_pair_sample_1240.ext - technology: sky130A

.subckt diff_pair_sample_1240 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=6.3726 ps=33.46 w=16.34 l=2.8
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=0 ps=0 w=16.34 l=2.8
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=6.3726 ps=33.46 w=16.34 l=2.8
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=0 ps=0 w=16.34 l=2.8
X4 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=6.3726 ps=33.46 w=16.34 l=2.8
X5 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=6.3726 ps=33.46 w=16.34 l=2.8
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=0 ps=0 w=16.34 l=2.8
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.3726 pd=33.46 as=0 ps=0 w=16.34 l=2.8
R0 VN VN.t1 230.256
R1 VN VN.t0 182.21
R2 VTAIL.n1 VTAIL.t2 43.3432
R3 VTAIL.n3 VTAIL.t3 43.343
R4 VTAIL.n0 VTAIL.t1 43.343
R5 VTAIL.n2 VTAIL.t0 43.343
R6 VTAIL.n1 VTAIL.n0 31.8496
R7 VTAIL.n3 VTAIL.n2 29.1514
R8 VTAIL.n2 VTAIL.n1 1.81947
R9 VTAIL VTAIL.n0 1.20309
R10 VTAIL VTAIL.n3 0.616879
R11 VDD2.n0 VDD2.t1 103.163
R12 VDD2.n0 VDD2.t0 60.0218
R13 VDD2 VDD2.n0 0.733259
R14 B.n582 B.n581 585
R15 B.n583 B.n116 585
R16 B.n585 B.n584 585
R17 B.n587 B.n115 585
R18 B.n590 B.n589 585
R19 B.n591 B.n114 585
R20 B.n593 B.n592 585
R21 B.n595 B.n113 585
R22 B.n598 B.n597 585
R23 B.n599 B.n112 585
R24 B.n601 B.n600 585
R25 B.n603 B.n111 585
R26 B.n606 B.n605 585
R27 B.n607 B.n110 585
R28 B.n609 B.n608 585
R29 B.n611 B.n109 585
R30 B.n614 B.n613 585
R31 B.n615 B.n108 585
R32 B.n617 B.n616 585
R33 B.n619 B.n107 585
R34 B.n622 B.n621 585
R35 B.n623 B.n106 585
R36 B.n625 B.n624 585
R37 B.n627 B.n105 585
R38 B.n630 B.n629 585
R39 B.n631 B.n104 585
R40 B.n633 B.n632 585
R41 B.n635 B.n103 585
R42 B.n638 B.n637 585
R43 B.n639 B.n102 585
R44 B.n641 B.n640 585
R45 B.n643 B.n101 585
R46 B.n646 B.n645 585
R47 B.n647 B.n100 585
R48 B.n649 B.n648 585
R49 B.n651 B.n99 585
R50 B.n654 B.n653 585
R51 B.n655 B.n98 585
R52 B.n657 B.n656 585
R53 B.n659 B.n97 585
R54 B.n662 B.n661 585
R55 B.n663 B.n96 585
R56 B.n665 B.n664 585
R57 B.n667 B.n95 585
R58 B.n670 B.n669 585
R59 B.n671 B.n94 585
R60 B.n673 B.n672 585
R61 B.n675 B.n93 585
R62 B.n678 B.n677 585
R63 B.n679 B.n92 585
R64 B.n681 B.n680 585
R65 B.n683 B.n91 585
R66 B.n685 B.n684 585
R67 B.n687 B.n686 585
R68 B.n690 B.n689 585
R69 B.n691 B.n86 585
R70 B.n693 B.n692 585
R71 B.n695 B.n85 585
R72 B.n698 B.n697 585
R73 B.n699 B.n84 585
R74 B.n701 B.n700 585
R75 B.n703 B.n83 585
R76 B.n705 B.n704 585
R77 B.n707 B.n706 585
R78 B.n710 B.n709 585
R79 B.n711 B.n78 585
R80 B.n713 B.n712 585
R81 B.n715 B.n77 585
R82 B.n718 B.n717 585
R83 B.n719 B.n76 585
R84 B.n721 B.n720 585
R85 B.n723 B.n75 585
R86 B.n726 B.n725 585
R87 B.n727 B.n74 585
R88 B.n729 B.n728 585
R89 B.n731 B.n73 585
R90 B.n734 B.n733 585
R91 B.n735 B.n72 585
R92 B.n737 B.n736 585
R93 B.n739 B.n71 585
R94 B.n742 B.n741 585
R95 B.n743 B.n70 585
R96 B.n745 B.n744 585
R97 B.n747 B.n69 585
R98 B.n750 B.n749 585
R99 B.n751 B.n68 585
R100 B.n753 B.n752 585
R101 B.n755 B.n67 585
R102 B.n758 B.n757 585
R103 B.n759 B.n66 585
R104 B.n761 B.n760 585
R105 B.n763 B.n65 585
R106 B.n766 B.n765 585
R107 B.n767 B.n64 585
R108 B.n769 B.n768 585
R109 B.n771 B.n63 585
R110 B.n774 B.n773 585
R111 B.n775 B.n62 585
R112 B.n777 B.n776 585
R113 B.n779 B.n61 585
R114 B.n782 B.n781 585
R115 B.n783 B.n60 585
R116 B.n785 B.n784 585
R117 B.n787 B.n59 585
R118 B.n790 B.n789 585
R119 B.n791 B.n58 585
R120 B.n793 B.n792 585
R121 B.n795 B.n57 585
R122 B.n798 B.n797 585
R123 B.n799 B.n56 585
R124 B.n801 B.n800 585
R125 B.n803 B.n55 585
R126 B.n806 B.n805 585
R127 B.n807 B.n54 585
R128 B.n809 B.n808 585
R129 B.n811 B.n53 585
R130 B.n814 B.n813 585
R131 B.n815 B.n52 585
R132 B.n579 B.n50 585
R133 B.n818 B.n50 585
R134 B.n578 B.n49 585
R135 B.n819 B.n49 585
R136 B.n577 B.n48 585
R137 B.n820 B.n48 585
R138 B.n576 B.n575 585
R139 B.n575 B.n44 585
R140 B.n574 B.n43 585
R141 B.n826 B.n43 585
R142 B.n573 B.n42 585
R143 B.n827 B.n42 585
R144 B.n572 B.n41 585
R145 B.n828 B.n41 585
R146 B.n571 B.n570 585
R147 B.n570 B.n40 585
R148 B.n569 B.n36 585
R149 B.n834 B.n36 585
R150 B.n568 B.n35 585
R151 B.n835 B.n35 585
R152 B.n567 B.n34 585
R153 B.n836 B.n34 585
R154 B.n566 B.n565 585
R155 B.n565 B.n30 585
R156 B.n564 B.n29 585
R157 B.n842 B.n29 585
R158 B.n563 B.n28 585
R159 B.n843 B.n28 585
R160 B.n562 B.n27 585
R161 B.n844 B.n27 585
R162 B.n561 B.n560 585
R163 B.n560 B.n23 585
R164 B.n559 B.n22 585
R165 B.n850 B.n22 585
R166 B.n558 B.n21 585
R167 B.n851 B.n21 585
R168 B.n557 B.n20 585
R169 B.n852 B.n20 585
R170 B.n556 B.n555 585
R171 B.n555 B.n16 585
R172 B.n554 B.n15 585
R173 B.n858 B.n15 585
R174 B.n553 B.n14 585
R175 B.n859 B.n14 585
R176 B.n552 B.n13 585
R177 B.n860 B.n13 585
R178 B.n551 B.n550 585
R179 B.n550 B.n12 585
R180 B.n549 B.n548 585
R181 B.n549 B.n8 585
R182 B.n547 B.n7 585
R183 B.n867 B.n7 585
R184 B.n546 B.n6 585
R185 B.n868 B.n6 585
R186 B.n545 B.n5 585
R187 B.n869 B.n5 585
R188 B.n544 B.n543 585
R189 B.n543 B.n4 585
R190 B.n542 B.n117 585
R191 B.n542 B.n541 585
R192 B.n532 B.n118 585
R193 B.n119 B.n118 585
R194 B.n534 B.n533 585
R195 B.n535 B.n534 585
R196 B.n531 B.n124 585
R197 B.n124 B.n123 585
R198 B.n530 B.n529 585
R199 B.n529 B.n528 585
R200 B.n126 B.n125 585
R201 B.n127 B.n126 585
R202 B.n521 B.n520 585
R203 B.n522 B.n521 585
R204 B.n519 B.n132 585
R205 B.n132 B.n131 585
R206 B.n518 B.n517 585
R207 B.n517 B.n516 585
R208 B.n134 B.n133 585
R209 B.n135 B.n134 585
R210 B.n509 B.n508 585
R211 B.n510 B.n509 585
R212 B.n507 B.n140 585
R213 B.n140 B.n139 585
R214 B.n506 B.n505 585
R215 B.n505 B.n504 585
R216 B.n142 B.n141 585
R217 B.n143 B.n142 585
R218 B.n497 B.n496 585
R219 B.n498 B.n497 585
R220 B.n495 B.n148 585
R221 B.n148 B.n147 585
R222 B.n494 B.n493 585
R223 B.n493 B.n492 585
R224 B.n150 B.n149 585
R225 B.n485 B.n150 585
R226 B.n484 B.n483 585
R227 B.n486 B.n484 585
R228 B.n482 B.n155 585
R229 B.n155 B.n154 585
R230 B.n481 B.n480 585
R231 B.n480 B.n479 585
R232 B.n157 B.n156 585
R233 B.n158 B.n157 585
R234 B.n472 B.n471 585
R235 B.n473 B.n472 585
R236 B.n470 B.n163 585
R237 B.n163 B.n162 585
R238 B.n469 B.n468 585
R239 B.n468 B.n467 585
R240 B.n464 B.n167 585
R241 B.n463 B.n462 585
R242 B.n460 B.n168 585
R243 B.n460 B.n166 585
R244 B.n459 B.n458 585
R245 B.n457 B.n456 585
R246 B.n455 B.n170 585
R247 B.n453 B.n452 585
R248 B.n451 B.n171 585
R249 B.n450 B.n449 585
R250 B.n447 B.n172 585
R251 B.n445 B.n444 585
R252 B.n443 B.n173 585
R253 B.n442 B.n441 585
R254 B.n439 B.n174 585
R255 B.n437 B.n436 585
R256 B.n435 B.n175 585
R257 B.n434 B.n433 585
R258 B.n431 B.n176 585
R259 B.n429 B.n428 585
R260 B.n427 B.n177 585
R261 B.n426 B.n425 585
R262 B.n423 B.n178 585
R263 B.n421 B.n420 585
R264 B.n419 B.n179 585
R265 B.n418 B.n417 585
R266 B.n415 B.n180 585
R267 B.n413 B.n412 585
R268 B.n411 B.n181 585
R269 B.n410 B.n409 585
R270 B.n407 B.n182 585
R271 B.n405 B.n404 585
R272 B.n403 B.n183 585
R273 B.n402 B.n401 585
R274 B.n399 B.n184 585
R275 B.n397 B.n396 585
R276 B.n395 B.n185 585
R277 B.n394 B.n393 585
R278 B.n391 B.n186 585
R279 B.n389 B.n388 585
R280 B.n387 B.n187 585
R281 B.n386 B.n385 585
R282 B.n383 B.n188 585
R283 B.n381 B.n380 585
R284 B.n379 B.n189 585
R285 B.n378 B.n377 585
R286 B.n375 B.n190 585
R287 B.n373 B.n372 585
R288 B.n371 B.n191 585
R289 B.n370 B.n369 585
R290 B.n367 B.n192 585
R291 B.n365 B.n364 585
R292 B.n363 B.n193 585
R293 B.n362 B.n361 585
R294 B.n359 B.n194 585
R295 B.n357 B.n356 585
R296 B.n355 B.n195 585
R297 B.n354 B.n353 585
R298 B.n351 B.n199 585
R299 B.n349 B.n348 585
R300 B.n347 B.n200 585
R301 B.n346 B.n345 585
R302 B.n343 B.n201 585
R303 B.n341 B.n340 585
R304 B.n339 B.n202 585
R305 B.n337 B.n336 585
R306 B.n334 B.n205 585
R307 B.n332 B.n331 585
R308 B.n330 B.n206 585
R309 B.n329 B.n328 585
R310 B.n326 B.n207 585
R311 B.n324 B.n323 585
R312 B.n322 B.n208 585
R313 B.n321 B.n320 585
R314 B.n318 B.n209 585
R315 B.n316 B.n315 585
R316 B.n314 B.n210 585
R317 B.n313 B.n312 585
R318 B.n310 B.n211 585
R319 B.n308 B.n307 585
R320 B.n306 B.n212 585
R321 B.n305 B.n304 585
R322 B.n302 B.n213 585
R323 B.n300 B.n299 585
R324 B.n298 B.n214 585
R325 B.n297 B.n296 585
R326 B.n294 B.n215 585
R327 B.n292 B.n291 585
R328 B.n290 B.n216 585
R329 B.n289 B.n288 585
R330 B.n286 B.n217 585
R331 B.n284 B.n283 585
R332 B.n282 B.n218 585
R333 B.n281 B.n280 585
R334 B.n278 B.n219 585
R335 B.n276 B.n275 585
R336 B.n274 B.n220 585
R337 B.n273 B.n272 585
R338 B.n270 B.n221 585
R339 B.n268 B.n267 585
R340 B.n266 B.n222 585
R341 B.n265 B.n264 585
R342 B.n262 B.n223 585
R343 B.n260 B.n259 585
R344 B.n258 B.n224 585
R345 B.n257 B.n256 585
R346 B.n254 B.n225 585
R347 B.n252 B.n251 585
R348 B.n250 B.n226 585
R349 B.n249 B.n248 585
R350 B.n246 B.n227 585
R351 B.n244 B.n243 585
R352 B.n242 B.n228 585
R353 B.n241 B.n240 585
R354 B.n238 B.n229 585
R355 B.n236 B.n235 585
R356 B.n234 B.n230 585
R357 B.n233 B.n232 585
R358 B.n165 B.n164 585
R359 B.n166 B.n165 585
R360 B.n466 B.n465 585
R361 B.n467 B.n466 585
R362 B.n161 B.n160 585
R363 B.n162 B.n161 585
R364 B.n475 B.n474 585
R365 B.n474 B.n473 585
R366 B.n476 B.n159 585
R367 B.n159 B.n158 585
R368 B.n478 B.n477 585
R369 B.n479 B.n478 585
R370 B.n153 B.n152 585
R371 B.n154 B.n153 585
R372 B.n488 B.n487 585
R373 B.n487 B.n486 585
R374 B.n489 B.n151 585
R375 B.n485 B.n151 585
R376 B.n491 B.n490 585
R377 B.n492 B.n491 585
R378 B.n146 B.n145 585
R379 B.n147 B.n146 585
R380 B.n500 B.n499 585
R381 B.n499 B.n498 585
R382 B.n501 B.n144 585
R383 B.n144 B.n143 585
R384 B.n503 B.n502 585
R385 B.n504 B.n503 585
R386 B.n138 B.n137 585
R387 B.n139 B.n138 585
R388 B.n512 B.n511 585
R389 B.n511 B.n510 585
R390 B.n513 B.n136 585
R391 B.n136 B.n135 585
R392 B.n515 B.n514 585
R393 B.n516 B.n515 585
R394 B.n130 B.n129 585
R395 B.n131 B.n130 585
R396 B.n524 B.n523 585
R397 B.n523 B.n522 585
R398 B.n525 B.n128 585
R399 B.n128 B.n127 585
R400 B.n527 B.n526 585
R401 B.n528 B.n527 585
R402 B.n122 B.n121 585
R403 B.n123 B.n122 585
R404 B.n537 B.n536 585
R405 B.n536 B.n535 585
R406 B.n538 B.n120 585
R407 B.n120 B.n119 585
R408 B.n540 B.n539 585
R409 B.n541 B.n540 585
R410 B.n3 B.n0 585
R411 B.n4 B.n3 585
R412 B.n866 B.n1 585
R413 B.n867 B.n866 585
R414 B.n865 B.n864 585
R415 B.n865 B.n8 585
R416 B.n863 B.n9 585
R417 B.n12 B.n9 585
R418 B.n862 B.n861 585
R419 B.n861 B.n860 585
R420 B.n11 B.n10 585
R421 B.n859 B.n11 585
R422 B.n857 B.n856 585
R423 B.n858 B.n857 585
R424 B.n855 B.n17 585
R425 B.n17 B.n16 585
R426 B.n854 B.n853 585
R427 B.n853 B.n852 585
R428 B.n19 B.n18 585
R429 B.n851 B.n19 585
R430 B.n849 B.n848 585
R431 B.n850 B.n849 585
R432 B.n847 B.n24 585
R433 B.n24 B.n23 585
R434 B.n846 B.n845 585
R435 B.n845 B.n844 585
R436 B.n26 B.n25 585
R437 B.n843 B.n26 585
R438 B.n841 B.n840 585
R439 B.n842 B.n841 585
R440 B.n839 B.n31 585
R441 B.n31 B.n30 585
R442 B.n838 B.n837 585
R443 B.n837 B.n836 585
R444 B.n33 B.n32 585
R445 B.n835 B.n33 585
R446 B.n833 B.n832 585
R447 B.n834 B.n833 585
R448 B.n831 B.n37 585
R449 B.n40 B.n37 585
R450 B.n830 B.n829 585
R451 B.n829 B.n828 585
R452 B.n39 B.n38 585
R453 B.n827 B.n39 585
R454 B.n825 B.n824 585
R455 B.n826 B.n825 585
R456 B.n823 B.n45 585
R457 B.n45 B.n44 585
R458 B.n822 B.n821 585
R459 B.n821 B.n820 585
R460 B.n47 B.n46 585
R461 B.n819 B.n47 585
R462 B.n817 B.n816 585
R463 B.n818 B.n817 585
R464 B.n870 B.n869 585
R465 B.n868 B.n2 585
R466 B.n817 B.n52 530.939
R467 B.n581 B.n50 530.939
R468 B.n468 B.n165 530.939
R469 B.n466 B.n167 530.939
R470 B.n79 B.t2 348.971
R471 B.n87 B.t13 348.971
R472 B.n203 B.t10 348.971
R473 B.n196 B.t6 348.971
R474 B.n580 B.n51 256.663
R475 B.n586 B.n51 256.663
R476 B.n588 B.n51 256.663
R477 B.n594 B.n51 256.663
R478 B.n596 B.n51 256.663
R479 B.n602 B.n51 256.663
R480 B.n604 B.n51 256.663
R481 B.n610 B.n51 256.663
R482 B.n612 B.n51 256.663
R483 B.n618 B.n51 256.663
R484 B.n620 B.n51 256.663
R485 B.n626 B.n51 256.663
R486 B.n628 B.n51 256.663
R487 B.n634 B.n51 256.663
R488 B.n636 B.n51 256.663
R489 B.n642 B.n51 256.663
R490 B.n644 B.n51 256.663
R491 B.n650 B.n51 256.663
R492 B.n652 B.n51 256.663
R493 B.n658 B.n51 256.663
R494 B.n660 B.n51 256.663
R495 B.n666 B.n51 256.663
R496 B.n668 B.n51 256.663
R497 B.n674 B.n51 256.663
R498 B.n676 B.n51 256.663
R499 B.n682 B.n51 256.663
R500 B.n90 B.n51 256.663
R501 B.n688 B.n51 256.663
R502 B.n694 B.n51 256.663
R503 B.n696 B.n51 256.663
R504 B.n702 B.n51 256.663
R505 B.n82 B.n51 256.663
R506 B.n708 B.n51 256.663
R507 B.n714 B.n51 256.663
R508 B.n716 B.n51 256.663
R509 B.n722 B.n51 256.663
R510 B.n724 B.n51 256.663
R511 B.n730 B.n51 256.663
R512 B.n732 B.n51 256.663
R513 B.n738 B.n51 256.663
R514 B.n740 B.n51 256.663
R515 B.n746 B.n51 256.663
R516 B.n748 B.n51 256.663
R517 B.n754 B.n51 256.663
R518 B.n756 B.n51 256.663
R519 B.n762 B.n51 256.663
R520 B.n764 B.n51 256.663
R521 B.n770 B.n51 256.663
R522 B.n772 B.n51 256.663
R523 B.n778 B.n51 256.663
R524 B.n780 B.n51 256.663
R525 B.n786 B.n51 256.663
R526 B.n788 B.n51 256.663
R527 B.n794 B.n51 256.663
R528 B.n796 B.n51 256.663
R529 B.n802 B.n51 256.663
R530 B.n804 B.n51 256.663
R531 B.n810 B.n51 256.663
R532 B.n812 B.n51 256.663
R533 B.n461 B.n166 256.663
R534 B.n169 B.n166 256.663
R535 B.n454 B.n166 256.663
R536 B.n448 B.n166 256.663
R537 B.n446 B.n166 256.663
R538 B.n440 B.n166 256.663
R539 B.n438 B.n166 256.663
R540 B.n432 B.n166 256.663
R541 B.n430 B.n166 256.663
R542 B.n424 B.n166 256.663
R543 B.n422 B.n166 256.663
R544 B.n416 B.n166 256.663
R545 B.n414 B.n166 256.663
R546 B.n408 B.n166 256.663
R547 B.n406 B.n166 256.663
R548 B.n400 B.n166 256.663
R549 B.n398 B.n166 256.663
R550 B.n392 B.n166 256.663
R551 B.n390 B.n166 256.663
R552 B.n384 B.n166 256.663
R553 B.n382 B.n166 256.663
R554 B.n376 B.n166 256.663
R555 B.n374 B.n166 256.663
R556 B.n368 B.n166 256.663
R557 B.n366 B.n166 256.663
R558 B.n360 B.n166 256.663
R559 B.n358 B.n166 256.663
R560 B.n352 B.n166 256.663
R561 B.n350 B.n166 256.663
R562 B.n344 B.n166 256.663
R563 B.n342 B.n166 256.663
R564 B.n335 B.n166 256.663
R565 B.n333 B.n166 256.663
R566 B.n327 B.n166 256.663
R567 B.n325 B.n166 256.663
R568 B.n319 B.n166 256.663
R569 B.n317 B.n166 256.663
R570 B.n311 B.n166 256.663
R571 B.n309 B.n166 256.663
R572 B.n303 B.n166 256.663
R573 B.n301 B.n166 256.663
R574 B.n295 B.n166 256.663
R575 B.n293 B.n166 256.663
R576 B.n287 B.n166 256.663
R577 B.n285 B.n166 256.663
R578 B.n279 B.n166 256.663
R579 B.n277 B.n166 256.663
R580 B.n271 B.n166 256.663
R581 B.n269 B.n166 256.663
R582 B.n263 B.n166 256.663
R583 B.n261 B.n166 256.663
R584 B.n255 B.n166 256.663
R585 B.n253 B.n166 256.663
R586 B.n247 B.n166 256.663
R587 B.n245 B.n166 256.663
R588 B.n239 B.n166 256.663
R589 B.n237 B.n166 256.663
R590 B.n231 B.n166 256.663
R591 B.n872 B.n871 256.663
R592 B.n813 B.n811 163.367
R593 B.n809 B.n54 163.367
R594 B.n805 B.n803 163.367
R595 B.n801 B.n56 163.367
R596 B.n797 B.n795 163.367
R597 B.n793 B.n58 163.367
R598 B.n789 B.n787 163.367
R599 B.n785 B.n60 163.367
R600 B.n781 B.n779 163.367
R601 B.n777 B.n62 163.367
R602 B.n773 B.n771 163.367
R603 B.n769 B.n64 163.367
R604 B.n765 B.n763 163.367
R605 B.n761 B.n66 163.367
R606 B.n757 B.n755 163.367
R607 B.n753 B.n68 163.367
R608 B.n749 B.n747 163.367
R609 B.n745 B.n70 163.367
R610 B.n741 B.n739 163.367
R611 B.n737 B.n72 163.367
R612 B.n733 B.n731 163.367
R613 B.n729 B.n74 163.367
R614 B.n725 B.n723 163.367
R615 B.n721 B.n76 163.367
R616 B.n717 B.n715 163.367
R617 B.n713 B.n78 163.367
R618 B.n709 B.n707 163.367
R619 B.n704 B.n703 163.367
R620 B.n701 B.n84 163.367
R621 B.n697 B.n695 163.367
R622 B.n693 B.n86 163.367
R623 B.n689 B.n687 163.367
R624 B.n684 B.n683 163.367
R625 B.n681 B.n92 163.367
R626 B.n677 B.n675 163.367
R627 B.n673 B.n94 163.367
R628 B.n669 B.n667 163.367
R629 B.n665 B.n96 163.367
R630 B.n661 B.n659 163.367
R631 B.n657 B.n98 163.367
R632 B.n653 B.n651 163.367
R633 B.n649 B.n100 163.367
R634 B.n645 B.n643 163.367
R635 B.n641 B.n102 163.367
R636 B.n637 B.n635 163.367
R637 B.n633 B.n104 163.367
R638 B.n629 B.n627 163.367
R639 B.n625 B.n106 163.367
R640 B.n621 B.n619 163.367
R641 B.n617 B.n108 163.367
R642 B.n613 B.n611 163.367
R643 B.n609 B.n110 163.367
R644 B.n605 B.n603 163.367
R645 B.n601 B.n112 163.367
R646 B.n597 B.n595 163.367
R647 B.n593 B.n114 163.367
R648 B.n589 B.n587 163.367
R649 B.n585 B.n116 163.367
R650 B.n468 B.n163 163.367
R651 B.n472 B.n163 163.367
R652 B.n472 B.n157 163.367
R653 B.n480 B.n157 163.367
R654 B.n480 B.n155 163.367
R655 B.n484 B.n155 163.367
R656 B.n484 B.n150 163.367
R657 B.n493 B.n150 163.367
R658 B.n493 B.n148 163.367
R659 B.n497 B.n148 163.367
R660 B.n497 B.n142 163.367
R661 B.n505 B.n142 163.367
R662 B.n505 B.n140 163.367
R663 B.n509 B.n140 163.367
R664 B.n509 B.n134 163.367
R665 B.n517 B.n134 163.367
R666 B.n517 B.n132 163.367
R667 B.n521 B.n132 163.367
R668 B.n521 B.n126 163.367
R669 B.n529 B.n126 163.367
R670 B.n529 B.n124 163.367
R671 B.n534 B.n124 163.367
R672 B.n534 B.n118 163.367
R673 B.n542 B.n118 163.367
R674 B.n543 B.n542 163.367
R675 B.n543 B.n5 163.367
R676 B.n6 B.n5 163.367
R677 B.n7 B.n6 163.367
R678 B.n549 B.n7 163.367
R679 B.n550 B.n549 163.367
R680 B.n550 B.n13 163.367
R681 B.n14 B.n13 163.367
R682 B.n15 B.n14 163.367
R683 B.n555 B.n15 163.367
R684 B.n555 B.n20 163.367
R685 B.n21 B.n20 163.367
R686 B.n22 B.n21 163.367
R687 B.n560 B.n22 163.367
R688 B.n560 B.n27 163.367
R689 B.n28 B.n27 163.367
R690 B.n29 B.n28 163.367
R691 B.n565 B.n29 163.367
R692 B.n565 B.n34 163.367
R693 B.n35 B.n34 163.367
R694 B.n36 B.n35 163.367
R695 B.n570 B.n36 163.367
R696 B.n570 B.n41 163.367
R697 B.n42 B.n41 163.367
R698 B.n43 B.n42 163.367
R699 B.n575 B.n43 163.367
R700 B.n575 B.n48 163.367
R701 B.n49 B.n48 163.367
R702 B.n50 B.n49 163.367
R703 B.n462 B.n460 163.367
R704 B.n460 B.n459 163.367
R705 B.n456 B.n455 163.367
R706 B.n453 B.n171 163.367
R707 B.n449 B.n447 163.367
R708 B.n445 B.n173 163.367
R709 B.n441 B.n439 163.367
R710 B.n437 B.n175 163.367
R711 B.n433 B.n431 163.367
R712 B.n429 B.n177 163.367
R713 B.n425 B.n423 163.367
R714 B.n421 B.n179 163.367
R715 B.n417 B.n415 163.367
R716 B.n413 B.n181 163.367
R717 B.n409 B.n407 163.367
R718 B.n405 B.n183 163.367
R719 B.n401 B.n399 163.367
R720 B.n397 B.n185 163.367
R721 B.n393 B.n391 163.367
R722 B.n389 B.n187 163.367
R723 B.n385 B.n383 163.367
R724 B.n381 B.n189 163.367
R725 B.n377 B.n375 163.367
R726 B.n373 B.n191 163.367
R727 B.n369 B.n367 163.367
R728 B.n365 B.n193 163.367
R729 B.n361 B.n359 163.367
R730 B.n357 B.n195 163.367
R731 B.n353 B.n351 163.367
R732 B.n349 B.n200 163.367
R733 B.n345 B.n343 163.367
R734 B.n341 B.n202 163.367
R735 B.n336 B.n334 163.367
R736 B.n332 B.n206 163.367
R737 B.n328 B.n326 163.367
R738 B.n324 B.n208 163.367
R739 B.n320 B.n318 163.367
R740 B.n316 B.n210 163.367
R741 B.n312 B.n310 163.367
R742 B.n308 B.n212 163.367
R743 B.n304 B.n302 163.367
R744 B.n300 B.n214 163.367
R745 B.n296 B.n294 163.367
R746 B.n292 B.n216 163.367
R747 B.n288 B.n286 163.367
R748 B.n284 B.n218 163.367
R749 B.n280 B.n278 163.367
R750 B.n276 B.n220 163.367
R751 B.n272 B.n270 163.367
R752 B.n268 B.n222 163.367
R753 B.n264 B.n262 163.367
R754 B.n260 B.n224 163.367
R755 B.n256 B.n254 163.367
R756 B.n252 B.n226 163.367
R757 B.n248 B.n246 163.367
R758 B.n244 B.n228 163.367
R759 B.n240 B.n238 163.367
R760 B.n236 B.n230 163.367
R761 B.n232 B.n165 163.367
R762 B.n466 B.n161 163.367
R763 B.n474 B.n161 163.367
R764 B.n474 B.n159 163.367
R765 B.n478 B.n159 163.367
R766 B.n478 B.n153 163.367
R767 B.n487 B.n153 163.367
R768 B.n487 B.n151 163.367
R769 B.n491 B.n151 163.367
R770 B.n491 B.n146 163.367
R771 B.n499 B.n146 163.367
R772 B.n499 B.n144 163.367
R773 B.n503 B.n144 163.367
R774 B.n503 B.n138 163.367
R775 B.n511 B.n138 163.367
R776 B.n511 B.n136 163.367
R777 B.n515 B.n136 163.367
R778 B.n515 B.n130 163.367
R779 B.n523 B.n130 163.367
R780 B.n523 B.n128 163.367
R781 B.n527 B.n128 163.367
R782 B.n527 B.n122 163.367
R783 B.n536 B.n122 163.367
R784 B.n536 B.n120 163.367
R785 B.n540 B.n120 163.367
R786 B.n540 B.n3 163.367
R787 B.n870 B.n3 163.367
R788 B.n866 B.n2 163.367
R789 B.n866 B.n865 163.367
R790 B.n865 B.n9 163.367
R791 B.n861 B.n9 163.367
R792 B.n861 B.n11 163.367
R793 B.n857 B.n11 163.367
R794 B.n857 B.n17 163.367
R795 B.n853 B.n17 163.367
R796 B.n853 B.n19 163.367
R797 B.n849 B.n19 163.367
R798 B.n849 B.n24 163.367
R799 B.n845 B.n24 163.367
R800 B.n845 B.n26 163.367
R801 B.n841 B.n26 163.367
R802 B.n841 B.n31 163.367
R803 B.n837 B.n31 163.367
R804 B.n837 B.n33 163.367
R805 B.n833 B.n33 163.367
R806 B.n833 B.n37 163.367
R807 B.n829 B.n37 163.367
R808 B.n829 B.n39 163.367
R809 B.n825 B.n39 163.367
R810 B.n825 B.n45 163.367
R811 B.n821 B.n45 163.367
R812 B.n821 B.n47 163.367
R813 B.n817 B.n47 163.367
R814 B.n87 B.t14 128.45
R815 B.n203 B.t12 128.45
R816 B.n79 B.t4 128.428
R817 B.n196 B.t9 128.428
R818 B.n812 B.n52 71.676
R819 B.n811 B.n810 71.676
R820 B.n804 B.n54 71.676
R821 B.n803 B.n802 71.676
R822 B.n796 B.n56 71.676
R823 B.n795 B.n794 71.676
R824 B.n788 B.n58 71.676
R825 B.n787 B.n786 71.676
R826 B.n780 B.n60 71.676
R827 B.n779 B.n778 71.676
R828 B.n772 B.n62 71.676
R829 B.n771 B.n770 71.676
R830 B.n764 B.n64 71.676
R831 B.n763 B.n762 71.676
R832 B.n756 B.n66 71.676
R833 B.n755 B.n754 71.676
R834 B.n748 B.n68 71.676
R835 B.n747 B.n746 71.676
R836 B.n740 B.n70 71.676
R837 B.n739 B.n738 71.676
R838 B.n732 B.n72 71.676
R839 B.n731 B.n730 71.676
R840 B.n724 B.n74 71.676
R841 B.n723 B.n722 71.676
R842 B.n716 B.n76 71.676
R843 B.n715 B.n714 71.676
R844 B.n708 B.n78 71.676
R845 B.n707 B.n82 71.676
R846 B.n703 B.n702 71.676
R847 B.n696 B.n84 71.676
R848 B.n695 B.n694 71.676
R849 B.n688 B.n86 71.676
R850 B.n687 B.n90 71.676
R851 B.n683 B.n682 71.676
R852 B.n676 B.n92 71.676
R853 B.n675 B.n674 71.676
R854 B.n668 B.n94 71.676
R855 B.n667 B.n666 71.676
R856 B.n660 B.n96 71.676
R857 B.n659 B.n658 71.676
R858 B.n652 B.n98 71.676
R859 B.n651 B.n650 71.676
R860 B.n644 B.n100 71.676
R861 B.n643 B.n642 71.676
R862 B.n636 B.n102 71.676
R863 B.n635 B.n634 71.676
R864 B.n628 B.n104 71.676
R865 B.n627 B.n626 71.676
R866 B.n620 B.n106 71.676
R867 B.n619 B.n618 71.676
R868 B.n612 B.n108 71.676
R869 B.n611 B.n610 71.676
R870 B.n604 B.n110 71.676
R871 B.n603 B.n602 71.676
R872 B.n596 B.n112 71.676
R873 B.n595 B.n594 71.676
R874 B.n588 B.n114 71.676
R875 B.n587 B.n586 71.676
R876 B.n580 B.n116 71.676
R877 B.n581 B.n580 71.676
R878 B.n586 B.n585 71.676
R879 B.n589 B.n588 71.676
R880 B.n594 B.n593 71.676
R881 B.n597 B.n596 71.676
R882 B.n602 B.n601 71.676
R883 B.n605 B.n604 71.676
R884 B.n610 B.n609 71.676
R885 B.n613 B.n612 71.676
R886 B.n618 B.n617 71.676
R887 B.n621 B.n620 71.676
R888 B.n626 B.n625 71.676
R889 B.n629 B.n628 71.676
R890 B.n634 B.n633 71.676
R891 B.n637 B.n636 71.676
R892 B.n642 B.n641 71.676
R893 B.n645 B.n644 71.676
R894 B.n650 B.n649 71.676
R895 B.n653 B.n652 71.676
R896 B.n658 B.n657 71.676
R897 B.n661 B.n660 71.676
R898 B.n666 B.n665 71.676
R899 B.n669 B.n668 71.676
R900 B.n674 B.n673 71.676
R901 B.n677 B.n676 71.676
R902 B.n682 B.n681 71.676
R903 B.n684 B.n90 71.676
R904 B.n689 B.n688 71.676
R905 B.n694 B.n693 71.676
R906 B.n697 B.n696 71.676
R907 B.n702 B.n701 71.676
R908 B.n704 B.n82 71.676
R909 B.n709 B.n708 71.676
R910 B.n714 B.n713 71.676
R911 B.n717 B.n716 71.676
R912 B.n722 B.n721 71.676
R913 B.n725 B.n724 71.676
R914 B.n730 B.n729 71.676
R915 B.n733 B.n732 71.676
R916 B.n738 B.n737 71.676
R917 B.n741 B.n740 71.676
R918 B.n746 B.n745 71.676
R919 B.n749 B.n748 71.676
R920 B.n754 B.n753 71.676
R921 B.n757 B.n756 71.676
R922 B.n762 B.n761 71.676
R923 B.n765 B.n764 71.676
R924 B.n770 B.n769 71.676
R925 B.n773 B.n772 71.676
R926 B.n778 B.n777 71.676
R927 B.n781 B.n780 71.676
R928 B.n786 B.n785 71.676
R929 B.n789 B.n788 71.676
R930 B.n794 B.n793 71.676
R931 B.n797 B.n796 71.676
R932 B.n802 B.n801 71.676
R933 B.n805 B.n804 71.676
R934 B.n810 B.n809 71.676
R935 B.n813 B.n812 71.676
R936 B.n461 B.n167 71.676
R937 B.n459 B.n169 71.676
R938 B.n455 B.n454 71.676
R939 B.n448 B.n171 71.676
R940 B.n447 B.n446 71.676
R941 B.n440 B.n173 71.676
R942 B.n439 B.n438 71.676
R943 B.n432 B.n175 71.676
R944 B.n431 B.n430 71.676
R945 B.n424 B.n177 71.676
R946 B.n423 B.n422 71.676
R947 B.n416 B.n179 71.676
R948 B.n415 B.n414 71.676
R949 B.n408 B.n181 71.676
R950 B.n407 B.n406 71.676
R951 B.n400 B.n183 71.676
R952 B.n399 B.n398 71.676
R953 B.n392 B.n185 71.676
R954 B.n391 B.n390 71.676
R955 B.n384 B.n187 71.676
R956 B.n383 B.n382 71.676
R957 B.n376 B.n189 71.676
R958 B.n375 B.n374 71.676
R959 B.n368 B.n191 71.676
R960 B.n367 B.n366 71.676
R961 B.n360 B.n193 71.676
R962 B.n359 B.n358 71.676
R963 B.n352 B.n195 71.676
R964 B.n351 B.n350 71.676
R965 B.n344 B.n200 71.676
R966 B.n343 B.n342 71.676
R967 B.n335 B.n202 71.676
R968 B.n334 B.n333 71.676
R969 B.n327 B.n206 71.676
R970 B.n326 B.n325 71.676
R971 B.n319 B.n208 71.676
R972 B.n318 B.n317 71.676
R973 B.n311 B.n210 71.676
R974 B.n310 B.n309 71.676
R975 B.n303 B.n212 71.676
R976 B.n302 B.n301 71.676
R977 B.n295 B.n214 71.676
R978 B.n294 B.n293 71.676
R979 B.n287 B.n216 71.676
R980 B.n286 B.n285 71.676
R981 B.n279 B.n218 71.676
R982 B.n278 B.n277 71.676
R983 B.n271 B.n220 71.676
R984 B.n270 B.n269 71.676
R985 B.n263 B.n222 71.676
R986 B.n262 B.n261 71.676
R987 B.n255 B.n224 71.676
R988 B.n254 B.n253 71.676
R989 B.n247 B.n226 71.676
R990 B.n246 B.n245 71.676
R991 B.n239 B.n228 71.676
R992 B.n238 B.n237 71.676
R993 B.n231 B.n230 71.676
R994 B.n462 B.n461 71.676
R995 B.n456 B.n169 71.676
R996 B.n454 B.n453 71.676
R997 B.n449 B.n448 71.676
R998 B.n446 B.n445 71.676
R999 B.n441 B.n440 71.676
R1000 B.n438 B.n437 71.676
R1001 B.n433 B.n432 71.676
R1002 B.n430 B.n429 71.676
R1003 B.n425 B.n424 71.676
R1004 B.n422 B.n421 71.676
R1005 B.n417 B.n416 71.676
R1006 B.n414 B.n413 71.676
R1007 B.n409 B.n408 71.676
R1008 B.n406 B.n405 71.676
R1009 B.n401 B.n400 71.676
R1010 B.n398 B.n397 71.676
R1011 B.n393 B.n392 71.676
R1012 B.n390 B.n389 71.676
R1013 B.n385 B.n384 71.676
R1014 B.n382 B.n381 71.676
R1015 B.n377 B.n376 71.676
R1016 B.n374 B.n373 71.676
R1017 B.n369 B.n368 71.676
R1018 B.n366 B.n365 71.676
R1019 B.n361 B.n360 71.676
R1020 B.n358 B.n357 71.676
R1021 B.n353 B.n352 71.676
R1022 B.n350 B.n349 71.676
R1023 B.n345 B.n344 71.676
R1024 B.n342 B.n341 71.676
R1025 B.n336 B.n335 71.676
R1026 B.n333 B.n332 71.676
R1027 B.n328 B.n327 71.676
R1028 B.n325 B.n324 71.676
R1029 B.n320 B.n319 71.676
R1030 B.n317 B.n316 71.676
R1031 B.n312 B.n311 71.676
R1032 B.n309 B.n308 71.676
R1033 B.n304 B.n303 71.676
R1034 B.n301 B.n300 71.676
R1035 B.n296 B.n295 71.676
R1036 B.n293 B.n292 71.676
R1037 B.n288 B.n287 71.676
R1038 B.n285 B.n284 71.676
R1039 B.n280 B.n279 71.676
R1040 B.n277 B.n276 71.676
R1041 B.n272 B.n271 71.676
R1042 B.n269 B.n268 71.676
R1043 B.n264 B.n263 71.676
R1044 B.n261 B.n260 71.676
R1045 B.n256 B.n255 71.676
R1046 B.n253 B.n252 71.676
R1047 B.n248 B.n247 71.676
R1048 B.n245 B.n244 71.676
R1049 B.n240 B.n239 71.676
R1050 B.n237 B.n236 71.676
R1051 B.n232 B.n231 71.676
R1052 B.n871 B.n870 71.676
R1053 B.n871 B.n2 71.676
R1054 B.n88 B.t15 67.746
R1055 B.n204 B.t11 67.746
R1056 B.n80 B.t5 67.7243
R1057 B.n197 B.t8 67.7243
R1058 B.n467 B.n166 63.6137
R1059 B.n818 B.n51 63.6137
R1060 B.n80 B.n79 60.7035
R1061 B.n88 B.n87 60.7035
R1062 B.n204 B.n203 60.7035
R1063 B.n197 B.n196 60.7035
R1064 B.n81 B.n80 59.5399
R1065 B.n89 B.n88 59.5399
R1066 B.n338 B.n204 59.5399
R1067 B.n198 B.n197 59.5399
R1068 B.n467 B.n162 34.6061
R1069 B.n473 B.n162 34.6061
R1070 B.n473 B.n158 34.6061
R1071 B.n479 B.n158 34.6061
R1072 B.n479 B.n154 34.6061
R1073 B.n486 B.n154 34.6061
R1074 B.n486 B.n485 34.6061
R1075 B.n492 B.n147 34.6061
R1076 B.n498 B.n147 34.6061
R1077 B.n498 B.n143 34.6061
R1078 B.n504 B.n143 34.6061
R1079 B.n504 B.n139 34.6061
R1080 B.n510 B.n139 34.6061
R1081 B.n510 B.n135 34.6061
R1082 B.n516 B.n135 34.6061
R1083 B.n516 B.n131 34.6061
R1084 B.n522 B.n131 34.6061
R1085 B.n522 B.n127 34.6061
R1086 B.n528 B.n127 34.6061
R1087 B.n535 B.n123 34.6061
R1088 B.n535 B.n119 34.6061
R1089 B.n541 B.n119 34.6061
R1090 B.n541 B.n4 34.6061
R1091 B.n869 B.n4 34.6061
R1092 B.n869 B.n868 34.6061
R1093 B.n868 B.n867 34.6061
R1094 B.n867 B.n8 34.6061
R1095 B.n12 B.n8 34.6061
R1096 B.n860 B.n12 34.6061
R1097 B.n860 B.n859 34.6061
R1098 B.n858 B.n16 34.6061
R1099 B.n852 B.n16 34.6061
R1100 B.n852 B.n851 34.6061
R1101 B.n851 B.n850 34.6061
R1102 B.n850 B.n23 34.6061
R1103 B.n844 B.n23 34.6061
R1104 B.n844 B.n843 34.6061
R1105 B.n843 B.n842 34.6061
R1106 B.n842 B.n30 34.6061
R1107 B.n836 B.n30 34.6061
R1108 B.n836 B.n835 34.6061
R1109 B.n835 B.n834 34.6061
R1110 B.n828 B.n40 34.6061
R1111 B.n828 B.n827 34.6061
R1112 B.n827 B.n826 34.6061
R1113 B.n826 B.n44 34.6061
R1114 B.n820 B.n44 34.6061
R1115 B.n820 B.n819 34.6061
R1116 B.n819 B.n818 34.6061
R1117 B.n465 B.n464 34.4981
R1118 B.n469 B.n164 34.4981
R1119 B.n582 B.n579 34.4981
R1120 B.n816 B.n815 34.4981
R1121 B.n485 B.t7 30.5349
R1122 B.n40 B.t3 30.5349
R1123 B.t1 B.n123 24.428
R1124 B.n859 B.t0 24.428
R1125 B B.n872 18.0485
R1126 B.n465 B.n160 10.6151
R1127 B.n475 B.n160 10.6151
R1128 B.n476 B.n475 10.6151
R1129 B.n477 B.n476 10.6151
R1130 B.n477 B.n152 10.6151
R1131 B.n488 B.n152 10.6151
R1132 B.n489 B.n488 10.6151
R1133 B.n490 B.n489 10.6151
R1134 B.n490 B.n145 10.6151
R1135 B.n500 B.n145 10.6151
R1136 B.n501 B.n500 10.6151
R1137 B.n502 B.n501 10.6151
R1138 B.n502 B.n137 10.6151
R1139 B.n512 B.n137 10.6151
R1140 B.n513 B.n512 10.6151
R1141 B.n514 B.n513 10.6151
R1142 B.n514 B.n129 10.6151
R1143 B.n524 B.n129 10.6151
R1144 B.n525 B.n524 10.6151
R1145 B.n526 B.n525 10.6151
R1146 B.n526 B.n121 10.6151
R1147 B.n537 B.n121 10.6151
R1148 B.n538 B.n537 10.6151
R1149 B.n539 B.n538 10.6151
R1150 B.n539 B.n0 10.6151
R1151 B.n464 B.n463 10.6151
R1152 B.n463 B.n168 10.6151
R1153 B.n458 B.n168 10.6151
R1154 B.n458 B.n457 10.6151
R1155 B.n457 B.n170 10.6151
R1156 B.n452 B.n170 10.6151
R1157 B.n452 B.n451 10.6151
R1158 B.n451 B.n450 10.6151
R1159 B.n450 B.n172 10.6151
R1160 B.n444 B.n172 10.6151
R1161 B.n444 B.n443 10.6151
R1162 B.n443 B.n442 10.6151
R1163 B.n442 B.n174 10.6151
R1164 B.n436 B.n174 10.6151
R1165 B.n436 B.n435 10.6151
R1166 B.n435 B.n434 10.6151
R1167 B.n434 B.n176 10.6151
R1168 B.n428 B.n176 10.6151
R1169 B.n428 B.n427 10.6151
R1170 B.n427 B.n426 10.6151
R1171 B.n426 B.n178 10.6151
R1172 B.n420 B.n178 10.6151
R1173 B.n420 B.n419 10.6151
R1174 B.n419 B.n418 10.6151
R1175 B.n418 B.n180 10.6151
R1176 B.n412 B.n180 10.6151
R1177 B.n412 B.n411 10.6151
R1178 B.n411 B.n410 10.6151
R1179 B.n410 B.n182 10.6151
R1180 B.n404 B.n182 10.6151
R1181 B.n404 B.n403 10.6151
R1182 B.n403 B.n402 10.6151
R1183 B.n402 B.n184 10.6151
R1184 B.n396 B.n184 10.6151
R1185 B.n396 B.n395 10.6151
R1186 B.n395 B.n394 10.6151
R1187 B.n394 B.n186 10.6151
R1188 B.n388 B.n186 10.6151
R1189 B.n388 B.n387 10.6151
R1190 B.n387 B.n386 10.6151
R1191 B.n386 B.n188 10.6151
R1192 B.n380 B.n188 10.6151
R1193 B.n380 B.n379 10.6151
R1194 B.n379 B.n378 10.6151
R1195 B.n378 B.n190 10.6151
R1196 B.n372 B.n190 10.6151
R1197 B.n372 B.n371 10.6151
R1198 B.n371 B.n370 10.6151
R1199 B.n370 B.n192 10.6151
R1200 B.n364 B.n192 10.6151
R1201 B.n364 B.n363 10.6151
R1202 B.n363 B.n362 10.6151
R1203 B.n362 B.n194 10.6151
R1204 B.n356 B.n355 10.6151
R1205 B.n355 B.n354 10.6151
R1206 B.n354 B.n199 10.6151
R1207 B.n348 B.n199 10.6151
R1208 B.n348 B.n347 10.6151
R1209 B.n347 B.n346 10.6151
R1210 B.n346 B.n201 10.6151
R1211 B.n340 B.n201 10.6151
R1212 B.n340 B.n339 10.6151
R1213 B.n337 B.n205 10.6151
R1214 B.n331 B.n205 10.6151
R1215 B.n331 B.n330 10.6151
R1216 B.n330 B.n329 10.6151
R1217 B.n329 B.n207 10.6151
R1218 B.n323 B.n207 10.6151
R1219 B.n323 B.n322 10.6151
R1220 B.n322 B.n321 10.6151
R1221 B.n321 B.n209 10.6151
R1222 B.n315 B.n209 10.6151
R1223 B.n315 B.n314 10.6151
R1224 B.n314 B.n313 10.6151
R1225 B.n313 B.n211 10.6151
R1226 B.n307 B.n211 10.6151
R1227 B.n307 B.n306 10.6151
R1228 B.n306 B.n305 10.6151
R1229 B.n305 B.n213 10.6151
R1230 B.n299 B.n213 10.6151
R1231 B.n299 B.n298 10.6151
R1232 B.n298 B.n297 10.6151
R1233 B.n297 B.n215 10.6151
R1234 B.n291 B.n215 10.6151
R1235 B.n291 B.n290 10.6151
R1236 B.n290 B.n289 10.6151
R1237 B.n289 B.n217 10.6151
R1238 B.n283 B.n217 10.6151
R1239 B.n283 B.n282 10.6151
R1240 B.n282 B.n281 10.6151
R1241 B.n281 B.n219 10.6151
R1242 B.n275 B.n219 10.6151
R1243 B.n275 B.n274 10.6151
R1244 B.n274 B.n273 10.6151
R1245 B.n273 B.n221 10.6151
R1246 B.n267 B.n221 10.6151
R1247 B.n267 B.n266 10.6151
R1248 B.n266 B.n265 10.6151
R1249 B.n265 B.n223 10.6151
R1250 B.n259 B.n223 10.6151
R1251 B.n259 B.n258 10.6151
R1252 B.n258 B.n257 10.6151
R1253 B.n257 B.n225 10.6151
R1254 B.n251 B.n225 10.6151
R1255 B.n251 B.n250 10.6151
R1256 B.n250 B.n249 10.6151
R1257 B.n249 B.n227 10.6151
R1258 B.n243 B.n227 10.6151
R1259 B.n243 B.n242 10.6151
R1260 B.n242 B.n241 10.6151
R1261 B.n241 B.n229 10.6151
R1262 B.n235 B.n229 10.6151
R1263 B.n235 B.n234 10.6151
R1264 B.n234 B.n233 10.6151
R1265 B.n233 B.n164 10.6151
R1266 B.n470 B.n469 10.6151
R1267 B.n471 B.n470 10.6151
R1268 B.n471 B.n156 10.6151
R1269 B.n481 B.n156 10.6151
R1270 B.n482 B.n481 10.6151
R1271 B.n483 B.n482 10.6151
R1272 B.n483 B.n149 10.6151
R1273 B.n494 B.n149 10.6151
R1274 B.n495 B.n494 10.6151
R1275 B.n496 B.n495 10.6151
R1276 B.n496 B.n141 10.6151
R1277 B.n506 B.n141 10.6151
R1278 B.n507 B.n506 10.6151
R1279 B.n508 B.n507 10.6151
R1280 B.n508 B.n133 10.6151
R1281 B.n518 B.n133 10.6151
R1282 B.n519 B.n518 10.6151
R1283 B.n520 B.n519 10.6151
R1284 B.n520 B.n125 10.6151
R1285 B.n530 B.n125 10.6151
R1286 B.n531 B.n530 10.6151
R1287 B.n533 B.n531 10.6151
R1288 B.n533 B.n532 10.6151
R1289 B.n532 B.n117 10.6151
R1290 B.n544 B.n117 10.6151
R1291 B.n545 B.n544 10.6151
R1292 B.n546 B.n545 10.6151
R1293 B.n547 B.n546 10.6151
R1294 B.n548 B.n547 10.6151
R1295 B.n551 B.n548 10.6151
R1296 B.n552 B.n551 10.6151
R1297 B.n553 B.n552 10.6151
R1298 B.n554 B.n553 10.6151
R1299 B.n556 B.n554 10.6151
R1300 B.n557 B.n556 10.6151
R1301 B.n558 B.n557 10.6151
R1302 B.n559 B.n558 10.6151
R1303 B.n561 B.n559 10.6151
R1304 B.n562 B.n561 10.6151
R1305 B.n563 B.n562 10.6151
R1306 B.n564 B.n563 10.6151
R1307 B.n566 B.n564 10.6151
R1308 B.n567 B.n566 10.6151
R1309 B.n568 B.n567 10.6151
R1310 B.n569 B.n568 10.6151
R1311 B.n571 B.n569 10.6151
R1312 B.n572 B.n571 10.6151
R1313 B.n573 B.n572 10.6151
R1314 B.n574 B.n573 10.6151
R1315 B.n576 B.n574 10.6151
R1316 B.n577 B.n576 10.6151
R1317 B.n578 B.n577 10.6151
R1318 B.n579 B.n578 10.6151
R1319 B.n864 B.n1 10.6151
R1320 B.n864 B.n863 10.6151
R1321 B.n863 B.n862 10.6151
R1322 B.n862 B.n10 10.6151
R1323 B.n856 B.n10 10.6151
R1324 B.n856 B.n855 10.6151
R1325 B.n855 B.n854 10.6151
R1326 B.n854 B.n18 10.6151
R1327 B.n848 B.n18 10.6151
R1328 B.n848 B.n847 10.6151
R1329 B.n847 B.n846 10.6151
R1330 B.n846 B.n25 10.6151
R1331 B.n840 B.n25 10.6151
R1332 B.n840 B.n839 10.6151
R1333 B.n839 B.n838 10.6151
R1334 B.n838 B.n32 10.6151
R1335 B.n832 B.n32 10.6151
R1336 B.n832 B.n831 10.6151
R1337 B.n831 B.n830 10.6151
R1338 B.n830 B.n38 10.6151
R1339 B.n824 B.n38 10.6151
R1340 B.n824 B.n823 10.6151
R1341 B.n823 B.n822 10.6151
R1342 B.n822 B.n46 10.6151
R1343 B.n816 B.n46 10.6151
R1344 B.n815 B.n814 10.6151
R1345 B.n814 B.n53 10.6151
R1346 B.n808 B.n53 10.6151
R1347 B.n808 B.n807 10.6151
R1348 B.n807 B.n806 10.6151
R1349 B.n806 B.n55 10.6151
R1350 B.n800 B.n55 10.6151
R1351 B.n800 B.n799 10.6151
R1352 B.n799 B.n798 10.6151
R1353 B.n798 B.n57 10.6151
R1354 B.n792 B.n57 10.6151
R1355 B.n792 B.n791 10.6151
R1356 B.n791 B.n790 10.6151
R1357 B.n790 B.n59 10.6151
R1358 B.n784 B.n59 10.6151
R1359 B.n784 B.n783 10.6151
R1360 B.n783 B.n782 10.6151
R1361 B.n782 B.n61 10.6151
R1362 B.n776 B.n61 10.6151
R1363 B.n776 B.n775 10.6151
R1364 B.n775 B.n774 10.6151
R1365 B.n774 B.n63 10.6151
R1366 B.n768 B.n63 10.6151
R1367 B.n768 B.n767 10.6151
R1368 B.n767 B.n766 10.6151
R1369 B.n766 B.n65 10.6151
R1370 B.n760 B.n65 10.6151
R1371 B.n760 B.n759 10.6151
R1372 B.n759 B.n758 10.6151
R1373 B.n758 B.n67 10.6151
R1374 B.n752 B.n67 10.6151
R1375 B.n752 B.n751 10.6151
R1376 B.n751 B.n750 10.6151
R1377 B.n750 B.n69 10.6151
R1378 B.n744 B.n69 10.6151
R1379 B.n744 B.n743 10.6151
R1380 B.n743 B.n742 10.6151
R1381 B.n742 B.n71 10.6151
R1382 B.n736 B.n71 10.6151
R1383 B.n736 B.n735 10.6151
R1384 B.n735 B.n734 10.6151
R1385 B.n734 B.n73 10.6151
R1386 B.n728 B.n73 10.6151
R1387 B.n728 B.n727 10.6151
R1388 B.n727 B.n726 10.6151
R1389 B.n726 B.n75 10.6151
R1390 B.n720 B.n75 10.6151
R1391 B.n720 B.n719 10.6151
R1392 B.n719 B.n718 10.6151
R1393 B.n718 B.n77 10.6151
R1394 B.n712 B.n77 10.6151
R1395 B.n712 B.n711 10.6151
R1396 B.n711 B.n710 10.6151
R1397 B.n706 B.n705 10.6151
R1398 B.n705 B.n83 10.6151
R1399 B.n700 B.n83 10.6151
R1400 B.n700 B.n699 10.6151
R1401 B.n699 B.n698 10.6151
R1402 B.n698 B.n85 10.6151
R1403 B.n692 B.n85 10.6151
R1404 B.n692 B.n691 10.6151
R1405 B.n691 B.n690 10.6151
R1406 B.n686 B.n685 10.6151
R1407 B.n685 B.n91 10.6151
R1408 B.n680 B.n91 10.6151
R1409 B.n680 B.n679 10.6151
R1410 B.n679 B.n678 10.6151
R1411 B.n678 B.n93 10.6151
R1412 B.n672 B.n93 10.6151
R1413 B.n672 B.n671 10.6151
R1414 B.n671 B.n670 10.6151
R1415 B.n670 B.n95 10.6151
R1416 B.n664 B.n95 10.6151
R1417 B.n664 B.n663 10.6151
R1418 B.n663 B.n662 10.6151
R1419 B.n662 B.n97 10.6151
R1420 B.n656 B.n97 10.6151
R1421 B.n656 B.n655 10.6151
R1422 B.n655 B.n654 10.6151
R1423 B.n654 B.n99 10.6151
R1424 B.n648 B.n99 10.6151
R1425 B.n648 B.n647 10.6151
R1426 B.n647 B.n646 10.6151
R1427 B.n646 B.n101 10.6151
R1428 B.n640 B.n101 10.6151
R1429 B.n640 B.n639 10.6151
R1430 B.n639 B.n638 10.6151
R1431 B.n638 B.n103 10.6151
R1432 B.n632 B.n103 10.6151
R1433 B.n632 B.n631 10.6151
R1434 B.n631 B.n630 10.6151
R1435 B.n630 B.n105 10.6151
R1436 B.n624 B.n105 10.6151
R1437 B.n624 B.n623 10.6151
R1438 B.n623 B.n622 10.6151
R1439 B.n622 B.n107 10.6151
R1440 B.n616 B.n107 10.6151
R1441 B.n616 B.n615 10.6151
R1442 B.n615 B.n614 10.6151
R1443 B.n614 B.n109 10.6151
R1444 B.n608 B.n109 10.6151
R1445 B.n608 B.n607 10.6151
R1446 B.n607 B.n606 10.6151
R1447 B.n606 B.n111 10.6151
R1448 B.n600 B.n111 10.6151
R1449 B.n600 B.n599 10.6151
R1450 B.n599 B.n598 10.6151
R1451 B.n598 B.n113 10.6151
R1452 B.n592 B.n113 10.6151
R1453 B.n592 B.n591 10.6151
R1454 B.n591 B.n590 10.6151
R1455 B.n590 B.n115 10.6151
R1456 B.n584 B.n115 10.6151
R1457 B.n584 B.n583 10.6151
R1458 B.n583 B.n582 10.6151
R1459 B.n528 B.t1 10.1786
R1460 B.t0 B.n858 10.1786
R1461 B.n198 B.n194 9.36635
R1462 B.n338 B.n337 9.36635
R1463 B.n710 B.n81 9.36635
R1464 B.n686 B.n89 9.36635
R1465 B.n872 B.n0 8.11757
R1466 B.n872 B.n1 8.11757
R1467 B.n492 B.t7 4.07175
R1468 B.n834 B.t3 4.07175
R1469 B.n356 B.n198 1.24928
R1470 B.n339 B.n338 1.24928
R1471 B.n706 B.n81 1.24928
R1472 B.n690 B.n89 1.24928
R1473 VP.n0 VP.t1 230.255
R1474 VP.n0 VP.t0 181.779
R1475 VP VP.n0 0.431812
R1476 VDD1 VDD1.t1 104.364
R1477 VDD1 VDD1.t0 60.7545
C0 VN VDD2 3.73688f
C1 VDD2 VDD1 0.699257f
C2 VP VN 6.35171f
C3 VDD2 VTAIL 6.28008f
C4 VP VDD1 3.92731f
C5 VP VTAIL 3.239f
C6 VN VDD1 0.148548f
C7 VN VTAIL 3.22466f
C8 VP VDD2 0.342124f
C9 VDD1 VTAIL 6.22886f
C10 VDD2 B 5.27813f
C11 VDD1 B 8.72845f
C12 VTAIL B 9.212254f
C13 VN B 11.93742f
C14 VP B 6.945214f
C15 VDD1.t0 B 2.99776f
C16 VDD1.t1 B 3.7261f
C17 VP.t0 B 3.95588f
C18 VP.t1 B 4.54187f
C19 VP.n0 B 4.92234f
C20 VDD2.t1 B 3.67545f
C21 VDD2.t0 B 2.98663f
C22 VDD2.n0 B 3.20331f
C23 VTAIL.t1 B 2.89375f
C24 VTAIL.n0 B 1.8783f
C25 VTAIL.t2 B 2.89375f
C26 VTAIL.n1 B 1.91787f
C27 VTAIL.t0 B 2.89375f
C28 VTAIL.n2 B 1.74464f
C29 VTAIL.t3 B 2.89375f
C30 VTAIL.n3 B 1.66743f
C31 VN.t0 B 3.88856f
C32 VN.t1 B 4.46255f
.ends

