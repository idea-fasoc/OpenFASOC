* NGSPICE file created from diff_pair_sample_0703.ext - technology: sky130A

.subckt diff_pair_sample_0703 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t4 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=0.62535 ps=4.12 w=3.79 l=2.36
X1 VDD2.t5 VN.t0 VTAIL.t0 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0.62535 ps=4.12 w=3.79 l=2.36
X2 VDD2.t4 VN.t1 VTAIL.t2 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0.62535 ps=4.12 w=3.79 l=2.36
X3 VDD1.t5 VP.t1 VTAIL.t10 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=1.4781 ps=8.36 w=3.79 l=2.36
X4 VDD1.t3 VP.t2 VTAIL.t9 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=1.4781 ps=8.36 w=3.79 l=2.36
X5 VTAIL.t3 VN.t2 VDD2.t3 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=0.62535 ps=4.12 w=3.79 l=2.36
X6 VTAIL.t8 VP.t3 VDD1.t2 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=0.62535 ps=4.12 w=3.79 l=2.36
X7 VDD2.t2 VN.t3 VTAIL.t4 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=1.4781 ps=8.36 w=3.79 l=2.36
X8 VTAIL.t5 VN.t4 VDD2.t1 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=0.62535 ps=4.12 w=3.79 l=2.36
X9 VDD2.t0 VN.t5 VTAIL.t1 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=0.62535 pd=4.12 as=1.4781 ps=8.36 w=3.79 l=2.36
X10 B.t11 B.t9 B.t10 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0 ps=0 w=3.79 l=2.36
X11 B.t8 B.t6 B.t7 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0 ps=0 w=3.79 l=2.36
X12 VDD1.t1 VP.t4 VTAIL.t7 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0.62535 ps=4.12 w=3.79 l=2.36
X13 VDD1.t0 VP.t5 VTAIL.t6 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0.62535 ps=4.12 w=3.79 l=2.36
X14 B.t5 B.t3 B.t4 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0 ps=0 w=3.79 l=2.36
X15 B.t2 B.t0 B.t1 w_n3122_n1726# sky130_fd_pr__pfet_01v8 ad=1.4781 pd=8.36 as=0 ps=0 w=3.79 l=2.36
R0 VP.n11 VP.n8 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n7 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n6 161.3
R5 VP.n37 VP.n0 161.3
R6 VP.n36 VP.n35 161.3
R7 VP.n34 VP.n1 161.3
R8 VP.n33 VP.n32 161.3
R9 VP.n31 VP.n2 161.3
R10 VP.n30 VP.n29 161.3
R11 VP.n28 VP.n3 161.3
R12 VP.n27 VP.n26 161.3
R13 VP.n25 VP.n4 161.3
R14 VP.n24 VP.n23 161.3
R15 VP.n22 VP.n5 161.3
R16 VP.n21 VP.n20 101.459
R17 VP.n39 VP.n38 101.459
R18 VP.n19 VP.n18 101.459
R19 VP.n9 VP.t5 72.1577
R20 VP.n26 VP.n25 55.548
R21 VP.n32 VP.n1 55.548
R22 VP.n12 VP.n7 55.548
R23 VP.n10 VP.n9 47.9127
R24 VP.n21 VP.n19 41.4655
R25 VP.n30 VP.t3 38.7035
R26 VP.n20 VP.t4 38.7035
R27 VP.n38 VP.t1 38.7035
R28 VP.n10 VP.t0 38.7035
R29 VP.n18 VP.t2 38.7035
R30 VP.n25 VP.n24 25.4388
R31 VP.n36 VP.n1 25.4388
R32 VP.n16 VP.n7 25.4388
R33 VP.n24 VP.n5 24.4675
R34 VP.n26 VP.n3 24.4675
R35 VP.n30 VP.n3 24.4675
R36 VP.n31 VP.n30 24.4675
R37 VP.n32 VP.n31 24.4675
R38 VP.n37 VP.n36 24.4675
R39 VP.n17 VP.n16 24.4675
R40 VP.n11 VP.n10 24.4675
R41 VP.n12 VP.n11 24.4675
R42 VP.n20 VP.n5 9.29796
R43 VP.n38 VP.n37 9.29796
R44 VP.n18 VP.n17 9.29796
R45 VP.n9 VP.n8 6.8888
R46 VP.n19 VP.n6 0.278367
R47 VP.n22 VP.n21 0.278367
R48 VP.n39 VP.n0 0.278367
R49 VP.n13 VP.n8 0.189894
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n6 0.189894
R53 VP.n23 VP.n22 0.189894
R54 VP.n23 VP.n4 0.189894
R55 VP.n27 VP.n4 0.189894
R56 VP.n28 VP.n27 0.189894
R57 VP.n29 VP.n28 0.189894
R58 VP.n29 VP.n2 0.189894
R59 VP.n33 VP.n2 0.189894
R60 VP.n34 VP.n33 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n35 VP.n0 0.189894
R63 VP VP.n39 0.153454
R64 VDD1.n14 VDD1.n0 756.745
R65 VDD1.n33 VDD1.n19 756.745
R66 VDD1.n15 VDD1.n14 585
R67 VDD1.n13 VDD1.n12 585
R68 VDD1.n4 VDD1.n3 585
R69 VDD1.n7 VDD1.n6 585
R70 VDD1.n26 VDD1.n25 585
R71 VDD1.n23 VDD1.n22 585
R72 VDD1.n32 VDD1.n31 585
R73 VDD1.n34 VDD1.n33 585
R74 VDD1.t0 VDD1.n5 330.707
R75 VDD1.t1 VDD1.n24 330.707
R76 VDD1.n14 VDD1.n13 171.744
R77 VDD1.n13 VDD1.n3 171.744
R78 VDD1.n6 VDD1.n3 171.744
R79 VDD1.n25 VDD1.n22 171.744
R80 VDD1.n32 VDD1.n22 171.744
R81 VDD1.n33 VDD1.n32 171.744
R82 VDD1.n39 VDD1.n38 113.123
R83 VDD1.n41 VDD1.n40 112.599
R84 VDD1.n6 VDD1.t0 85.8723
R85 VDD1.n25 VDD1.t1 85.8723
R86 VDD1 VDD1.n18 49.6919
R87 VDD1.n39 VDD1.n37 49.5783
R88 VDD1.n41 VDD1.n39 36.2617
R89 VDD1.n7 VDD1.n5 16.3201
R90 VDD1.n26 VDD1.n24 16.3201
R91 VDD1.n8 VDD1.n4 12.8005
R92 VDD1.n27 VDD1.n23 12.8005
R93 VDD1.n12 VDD1.n11 12.0247
R94 VDD1.n31 VDD1.n30 12.0247
R95 VDD1.n15 VDD1.n2 11.249
R96 VDD1.n34 VDD1.n21 11.249
R97 VDD1.n16 VDD1.n0 10.4732
R98 VDD1.n35 VDD1.n19 10.4732
R99 VDD1.n18 VDD1.n17 9.45567
R100 VDD1.n37 VDD1.n36 9.45567
R101 VDD1.n17 VDD1.n16 9.3005
R102 VDD1.n2 VDD1.n1 9.3005
R103 VDD1.n11 VDD1.n10 9.3005
R104 VDD1.n9 VDD1.n8 9.3005
R105 VDD1.n36 VDD1.n35 9.3005
R106 VDD1.n21 VDD1.n20 9.3005
R107 VDD1.n30 VDD1.n29 9.3005
R108 VDD1.n28 VDD1.n27 9.3005
R109 VDD1.n40 VDD1.t4 8.57702
R110 VDD1.n40 VDD1.t3 8.57702
R111 VDD1.n38 VDD1.t2 8.57702
R112 VDD1.n38 VDD1.t5 8.57702
R113 VDD1.n9 VDD1.n5 3.78097
R114 VDD1.n28 VDD1.n24 3.78097
R115 VDD1.n18 VDD1.n0 3.49141
R116 VDD1.n37 VDD1.n19 3.49141
R117 VDD1.n16 VDD1.n15 2.71565
R118 VDD1.n35 VDD1.n34 2.71565
R119 VDD1.n12 VDD1.n2 1.93989
R120 VDD1.n31 VDD1.n21 1.93989
R121 VDD1.n11 VDD1.n4 1.16414
R122 VDD1.n30 VDD1.n23 1.16414
R123 VDD1 VDD1.n41 0.522052
R124 VDD1.n8 VDD1.n7 0.388379
R125 VDD1.n27 VDD1.n26 0.388379
R126 VDD1.n17 VDD1.n1 0.155672
R127 VDD1.n10 VDD1.n1 0.155672
R128 VDD1.n10 VDD1.n9 0.155672
R129 VDD1.n29 VDD1.n28 0.155672
R130 VDD1.n29 VDD1.n20 0.155672
R131 VDD1.n36 VDD1.n20 0.155672
R132 VTAIL.n82 VTAIL.n68 756.745
R133 VTAIL.n16 VTAIL.n2 756.745
R134 VTAIL.n62 VTAIL.n48 756.745
R135 VTAIL.n40 VTAIL.n26 756.745
R136 VTAIL.n75 VTAIL.n74 585
R137 VTAIL.n72 VTAIL.n71 585
R138 VTAIL.n81 VTAIL.n80 585
R139 VTAIL.n83 VTAIL.n82 585
R140 VTAIL.n9 VTAIL.n8 585
R141 VTAIL.n6 VTAIL.n5 585
R142 VTAIL.n15 VTAIL.n14 585
R143 VTAIL.n17 VTAIL.n16 585
R144 VTAIL.n63 VTAIL.n62 585
R145 VTAIL.n61 VTAIL.n60 585
R146 VTAIL.n52 VTAIL.n51 585
R147 VTAIL.n55 VTAIL.n54 585
R148 VTAIL.n41 VTAIL.n40 585
R149 VTAIL.n39 VTAIL.n38 585
R150 VTAIL.n30 VTAIL.n29 585
R151 VTAIL.n33 VTAIL.n32 585
R152 VTAIL.t1 VTAIL.n73 330.707
R153 VTAIL.t10 VTAIL.n7 330.707
R154 VTAIL.t9 VTAIL.n53 330.707
R155 VTAIL.t4 VTAIL.n31 330.707
R156 VTAIL.n74 VTAIL.n71 171.744
R157 VTAIL.n81 VTAIL.n71 171.744
R158 VTAIL.n82 VTAIL.n81 171.744
R159 VTAIL.n8 VTAIL.n5 171.744
R160 VTAIL.n15 VTAIL.n5 171.744
R161 VTAIL.n16 VTAIL.n15 171.744
R162 VTAIL.n62 VTAIL.n61 171.744
R163 VTAIL.n61 VTAIL.n51 171.744
R164 VTAIL.n54 VTAIL.n51 171.744
R165 VTAIL.n40 VTAIL.n39 171.744
R166 VTAIL.n39 VTAIL.n29 171.744
R167 VTAIL.n32 VTAIL.n29 171.744
R168 VTAIL.n47 VTAIL.n46 95.9198
R169 VTAIL.n25 VTAIL.n24 95.9198
R170 VTAIL.n1 VTAIL.n0 95.9197
R171 VTAIL.n23 VTAIL.n22 95.9197
R172 VTAIL.n74 VTAIL.t1 85.8723
R173 VTAIL.n8 VTAIL.t10 85.8723
R174 VTAIL.n54 VTAIL.t9 85.8723
R175 VTAIL.n32 VTAIL.t4 85.8723
R176 VTAIL.n87 VTAIL.n86 31.2157
R177 VTAIL.n21 VTAIL.n20 31.2157
R178 VTAIL.n67 VTAIL.n66 31.2157
R179 VTAIL.n45 VTAIL.n44 31.2157
R180 VTAIL.n25 VTAIL.n23 20.2721
R181 VTAIL.n87 VTAIL.n67 17.9531
R182 VTAIL.n75 VTAIL.n73 16.3201
R183 VTAIL.n9 VTAIL.n7 16.3201
R184 VTAIL.n55 VTAIL.n53 16.3201
R185 VTAIL.n33 VTAIL.n31 16.3201
R186 VTAIL.n76 VTAIL.n72 12.8005
R187 VTAIL.n10 VTAIL.n6 12.8005
R188 VTAIL.n56 VTAIL.n52 12.8005
R189 VTAIL.n34 VTAIL.n30 12.8005
R190 VTAIL.n80 VTAIL.n79 12.0247
R191 VTAIL.n14 VTAIL.n13 12.0247
R192 VTAIL.n60 VTAIL.n59 12.0247
R193 VTAIL.n38 VTAIL.n37 12.0247
R194 VTAIL.n83 VTAIL.n70 11.249
R195 VTAIL.n17 VTAIL.n4 11.249
R196 VTAIL.n63 VTAIL.n50 11.249
R197 VTAIL.n41 VTAIL.n28 11.249
R198 VTAIL.n84 VTAIL.n68 10.4732
R199 VTAIL.n18 VTAIL.n2 10.4732
R200 VTAIL.n64 VTAIL.n48 10.4732
R201 VTAIL.n42 VTAIL.n26 10.4732
R202 VTAIL.n86 VTAIL.n85 9.45567
R203 VTAIL.n20 VTAIL.n19 9.45567
R204 VTAIL.n66 VTAIL.n65 9.45567
R205 VTAIL.n44 VTAIL.n43 9.45567
R206 VTAIL.n85 VTAIL.n84 9.3005
R207 VTAIL.n70 VTAIL.n69 9.3005
R208 VTAIL.n79 VTAIL.n78 9.3005
R209 VTAIL.n77 VTAIL.n76 9.3005
R210 VTAIL.n19 VTAIL.n18 9.3005
R211 VTAIL.n4 VTAIL.n3 9.3005
R212 VTAIL.n13 VTAIL.n12 9.3005
R213 VTAIL.n11 VTAIL.n10 9.3005
R214 VTAIL.n65 VTAIL.n64 9.3005
R215 VTAIL.n50 VTAIL.n49 9.3005
R216 VTAIL.n59 VTAIL.n58 9.3005
R217 VTAIL.n57 VTAIL.n56 9.3005
R218 VTAIL.n43 VTAIL.n42 9.3005
R219 VTAIL.n28 VTAIL.n27 9.3005
R220 VTAIL.n37 VTAIL.n36 9.3005
R221 VTAIL.n35 VTAIL.n34 9.3005
R222 VTAIL.n0 VTAIL.t2 8.57702
R223 VTAIL.n0 VTAIL.t3 8.57702
R224 VTAIL.n22 VTAIL.t7 8.57702
R225 VTAIL.n22 VTAIL.t8 8.57702
R226 VTAIL.n46 VTAIL.t6 8.57702
R227 VTAIL.n46 VTAIL.t11 8.57702
R228 VTAIL.n24 VTAIL.t0 8.57702
R229 VTAIL.n24 VTAIL.t5 8.57702
R230 VTAIL.n77 VTAIL.n73 3.78097
R231 VTAIL.n11 VTAIL.n7 3.78097
R232 VTAIL.n57 VTAIL.n53 3.78097
R233 VTAIL.n35 VTAIL.n31 3.78097
R234 VTAIL.n86 VTAIL.n68 3.49141
R235 VTAIL.n20 VTAIL.n2 3.49141
R236 VTAIL.n66 VTAIL.n48 3.49141
R237 VTAIL.n44 VTAIL.n26 3.49141
R238 VTAIL.n84 VTAIL.n83 2.71565
R239 VTAIL.n18 VTAIL.n17 2.71565
R240 VTAIL.n64 VTAIL.n63 2.71565
R241 VTAIL.n42 VTAIL.n41 2.71565
R242 VTAIL.n45 VTAIL.n25 2.31947
R243 VTAIL.n67 VTAIL.n47 2.31947
R244 VTAIL.n23 VTAIL.n21 2.31947
R245 VTAIL.n80 VTAIL.n70 1.93989
R246 VTAIL.n14 VTAIL.n4 1.93989
R247 VTAIL.n60 VTAIL.n50 1.93989
R248 VTAIL.n38 VTAIL.n28 1.93989
R249 VTAIL VTAIL.n87 1.68153
R250 VTAIL.n47 VTAIL.n45 1.62981
R251 VTAIL.n21 VTAIL.n1 1.62981
R252 VTAIL.n79 VTAIL.n72 1.16414
R253 VTAIL.n13 VTAIL.n6 1.16414
R254 VTAIL.n59 VTAIL.n52 1.16414
R255 VTAIL.n37 VTAIL.n30 1.16414
R256 VTAIL VTAIL.n1 0.638431
R257 VTAIL.n76 VTAIL.n75 0.388379
R258 VTAIL.n10 VTAIL.n9 0.388379
R259 VTAIL.n56 VTAIL.n55 0.388379
R260 VTAIL.n34 VTAIL.n33 0.388379
R261 VTAIL.n78 VTAIL.n77 0.155672
R262 VTAIL.n78 VTAIL.n69 0.155672
R263 VTAIL.n85 VTAIL.n69 0.155672
R264 VTAIL.n12 VTAIL.n11 0.155672
R265 VTAIL.n12 VTAIL.n3 0.155672
R266 VTAIL.n19 VTAIL.n3 0.155672
R267 VTAIL.n65 VTAIL.n49 0.155672
R268 VTAIL.n58 VTAIL.n49 0.155672
R269 VTAIL.n58 VTAIL.n57 0.155672
R270 VTAIL.n43 VTAIL.n27 0.155672
R271 VTAIL.n36 VTAIL.n27 0.155672
R272 VTAIL.n36 VTAIL.n35 0.155672
R273 VN.n25 VN.n14 161.3
R274 VN.n24 VN.n23 161.3
R275 VN.n22 VN.n15 161.3
R276 VN.n21 VN.n20 161.3
R277 VN.n19 VN.n16 161.3
R278 VN.n11 VN.n0 161.3
R279 VN.n10 VN.n9 161.3
R280 VN.n8 VN.n1 161.3
R281 VN.n7 VN.n6 161.3
R282 VN.n5 VN.n2 161.3
R283 VN.n13 VN.n12 101.459
R284 VN.n27 VN.n26 101.459
R285 VN.n3 VN.t1 72.1577
R286 VN.n17 VN.t3 72.1577
R287 VN.n6 VN.n1 55.548
R288 VN.n20 VN.n15 55.548
R289 VN.n4 VN.n3 47.9127
R290 VN.n18 VN.n17 47.9127
R291 VN VN.n27 41.7444
R292 VN.n4 VN.t2 38.7035
R293 VN.n12 VN.t5 38.7035
R294 VN.n18 VN.t4 38.7035
R295 VN.n26 VN.t0 38.7035
R296 VN.n10 VN.n1 25.4388
R297 VN.n24 VN.n15 25.4388
R298 VN.n5 VN.n4 24.4675
R299 VN.n6 VN.n5 24.4675
R300 VN.n11 VN.n10 24.4675
R301 VN.n20 VN.n19 24.4675
R302 VN.n19 VN.n18 24.4675
R303 VN.n25 VN.n24 24.4675
R304 VN.n12 VN.n11 9.29796
R305 VN.n26 VN.n25 9.29796
R306 VN.n17 VN.n16 6.8888
R307 VN.n3 VN.n2 6.8888
R308 VN.n27 VN.n14 0.278367
R309 VN.n13 VN.n0 0.278367
R310 VN.n23 VN.n14 0.189894
R311 VN.n23 VN.n22 0.189894
R312 VN.n22 VN.n21 0.189894
R313 VN.n21 VN.n16 0.189894
R314 VN.n7 VN.n2 0.189894
R315 VN.n8 VN.n7 0.189894
R316 VN.n9 VN.n8 0.189894
R317 VN.n9 VN.n0 0.189894
R318 VN VN.n13 0.153454
R319 VDD2.n35 VDD2.n21 756.745
R320 VDD2.n14 VDD2.n0 756.745
R321 VDD2.n36 VDD2.n35 585
R322 VDD2.n34 VDD2.n33 585
R323 VDD2.n25 VDD2.n24 585
R324 VDD2.n28 VDD2.n27 585
R325 VDD2.n7 VDD2.n6 585
R326 VDD2.n4 VDD2.n3 585
R327 VDD2.n13 VDD2.n12 585
R328 VDD2.n15 VDD2.n14 585
R329 VDD2.t5 VDD2.n26 330.707
R330 VDD2.t4 VDD2.n5 330.707
R331 VDD2.n35 VDD2.n34 171.744
R332 VDD2.n34 VDD2.n24 171.744
R333 VDD2.n27 VDD2.n24 171.744
R334 VDD2.n6 VDD2.n3 171.744
R335 VDD2.n13 VDD2.n3 171.744
R336 VDD2.n14 VDD2.n13 171.744
R337 VDD2.n20 VDD2.n19 113.123
R338 VDD2 VDD2.n41 113.121
R339 VDD2.n27 VDD2.t5 85.8723
R340 VDD2.n6 VDD2.t4 85.8723
R341 VDD2.n20 VDD2.n18 49.5783
R342 VDD2.n40 VDD2.n39 47.8944
R343 VDD2.n40 VDD2.n20 34.5192
R344 VDD2.n28 VDD2.n26 16.3201
R345 VDD2.n7 VDD2.n5 16.3201
R346 VDD2.n29 VDD2.n25 12.8005
R347 VDD2.n8 VDD2.n4 12.8005
R348 VDD2.n33 VDD2.n32 12.0247
R349 VDD2.n12 VDD2.n11 12.0247
R350 VDD2.n36 VDD2.n23 11.249
R351 VDD2.n15 VDD2.n2 11.249
R352 VDD2.n37 VDD2.n21 10.4732
R353 VDD2.n16 VDD2.n0 10.4732
R354 VDD2.n39 VDD2.n38 9.45567
R355 VDD2.n18 VDD2.n17 9.45567
R356 VDD2.n38 VDD2.n37 9.3005
R357 VDD2.n23 VDD2.n22 9.3005
R358 VDD2.n32 VDD2.n31 9.3005
R359 VDD2.n30 VDD2.n29 9.3005
R360 VDD2.n17 VDD2.n16 9.3005
R361 VDD2.n2 VDD2.n1 9.3005
R362 VDD2.n11 VDD2.n10 9.3005
R363 VDD2.n9 VDD2.n8 9.3005
R364 VDD2.n41 VDD2.t1 8.57702
R365 VDD2.n41 VDD2.t2 8.57702
R366 VDD2.n19 VDD2.t3 8.57702
R367 VDD2.n19 VDD2.t0 8.57702
R368 VDD2.n30 VDD2.n26 3.78097
R369 VDD2.n9 VDD2.n5 3.78097
R370 VDD2.n39 VDD2.n21 3.49141
R371 VDD2.n18 VDD2.n0 3.49141
R372 VDD2.n37 VDD2.n36 2.71565
R373 VDD2.n16 VDD2.n15 2.71565
R374 VDD2.n33 VDD2.n23 1.93989
R375 VDD2.n12 VDD2.n2 1.93989
R376 VDD2 VDD2.n40 1.79791
R377 VDD2.n32 VDD2.n25 1.16414
R378 VDD2.n11 VDD2.n4 1.16414
R379 VDD2.n29 VDD2.n28 0.388379
R380 VDD2.n8 VDD2.n7 0.388379
R381 VDD2.n38 VDD2.n22 0.155672
R382 VDD2.n31 VDD2.n22 0.155672
R383 VDD2.n31 VDD2.n30 0.155672
R384 VDD2.n10 VDD2.n9 0.155672
R385 VDD2.n10 VDD2.n1 0.155672
R386 VDD2.n17 VDD2.n1 0.155672
R387 B.n260 B.n89 585
R388 B.n259 B.n258 585
R389 B.n257 B.n90 585
R390 B.n256 B.n255 585
R391 B.n254 B.n91 585
R392 B.n253 B.n252 585
R393 B.n251 B.n92 585
R394 B.n250 B.n249 585
R395 B.n248 B.n93 585
R396 B.n247 B.n246 585
R397 B.n245 B.n94 585
R398 B.n244 B.n243 585
R399 B.n242 B.n95 585
R400 B.n241 B.n240 585
R401 B.n239 B.n96 585
R402 B.n238 B.n237 585
R403 B.n236 B.n97 585
R404 B.n235 B.n234 585
R405 B.n232 B.n98 585
R406 B.n231 B.n230 585
R407 B.n229 B.n101 585
R408 B.n228 B.n227 585
R409 B.n226 B.n102 585
R410 B.n225 B.n224 585
R411 B.n223 B.n103 585
R412 B.n222 B.n221 585
R413 B.n220 B.n104 585
R414 B.n218 B.n217 585
R415 B.n216 B.n107 585
R416 B.n215 B.n214 585
R417 B.n213 B.n108 585
R418 B.n212 B.n211 585
R419 B.n210 B.n109 585
R420 B.n209 B.n208 585
R421 B.n207 B.n110 585
R422 B.n206 B.n205 585
R423 B.n204 B.n111 585
R424 B.n203 B.n202 585
R425 B.n201 B.n112 585
R426 B.n200 B.n199 585
R427 B.n198 B.n113 585
R428 B.n197 B.n196 585
R429 B.n195 B.n114 585
R430 B.n194 B.n193 585
R431 B.n192 B.n115 585
R432 B.n262 B.n261 585
R433 B.n263 B.n88 585
R434 B.n265 B.n264 585
R435 B.n266 B.n87 585
R436 B.n268 B.n267 585
R437 B.n269 B.n86 585
R438 B.n271 B.n270 585
R439 B.n272 B.n85 585
R440 B.n274 B.n273 585
R441 B.n275 B.n84 585
R442 B.n277 B.n276 585
R443 B.n278 B.n83 585
R444 B.n280 B.n279 585
R445 B.n281 B.n82 585
R446 B.n283 B.n282 585
R447 B.n284 B.n81 585
R448 B.n286 B.n285 585
R449 B.n287 B.n80 585
R450 B.n289 B.n288 585
R451 B.n290 B.n79 585
R452 B.n292 B.n291 585
R453 B.n293 B.n78 585
R454 B.n295 B.n294 585
R455 B.n296 B.n77 585
R456 B.n298 B.n297 585
R457 B.n299 B.n76 585
R458 B.n301 B.n300 585
R459 B.n302 B.n75 585
R460 B.n304 B.n303 585
R461 B.n305 B.n74 585
R462 B.n307 B.n306 585
R463 B.n308 B.n73 585
R464 B.n310 B.n309 585
R465 B.n311 B.n72 585
R466 B.n313 B.n312 585
R467 B.n314 B.n71 585
R468 B.n316 B.n315 585
R469 B.n317 B.n70 585
R470 B.n319 B.n318 585
R471 B.n320 B.n69 585
R472 B.n322 B.n321 585
R473 B.n323 B.n68 585
R474 B.n325 B.n324 585
R475 B.n326 B.n67 585
R476 B.n328 B.n327 585
R477 B.n329 B.n66 585
R478 B.n331 B.n330 585
R479 B.n332 B.n65 585
R480 B.n334 B.n333 585
R481 B.n335 B.n64 585
R482 B.n337 B.n336 585
R483 B.n338 B.n63 585
R484 B.n340 B.n339 585
R485 B.n341 B.n62 585
R486 B.n343 B.n342 585
R487 B.n344 B.n61 585
R488 B.n346 B.n345 585
R489 B.n347 B.n60 585
R490 B.n349 B.n348 585
R491 B.n350 B.n59 585
R492 B.n352 B.n351 585
R493 B.n353 B.n58 585
R494 B.n355 B.n354 585
R495 B.n356 B.n57 585
R496 B.n358 B.n357 585
R497 B.n359 B.n56 585
R498 B.n361 B.n360 585
R499 B.n362 B.n55 585
R500 B.n364 B.n363 585
R501 B.n365 B.n54 585
R502 B.n367 B.n366 585
R503 B.n368 B.n53 585
R504 B.n370 B.n369 585
R505 B.n371 B.n52 585
R506 B.n373 B.n372 585
R507 B.n374 B.n51 585
R508 B.n376 B.n375 585
R509 B.n377 B.n50 585
R510 B.n379 B.n378 585
R511 B.n380 B.n49 585
R512 B.n449 B.n448 585
R513 B.n447 B.n22 585
R514 B.n446 B.n445 585
R515 B.n444 B.n23 585
R516 B.n443 B.n442 585
R517 B.n441 B.n24 585
R518 B.n440 B.n439 585
R519 B.n438 B.n25 585
R520 B.n437 B.n436 585
R521 B.n435 B.n26 585
R522 B.n434 B.n433 585
R523 B.n432 B.n27 585
R524 B.n431 B.n430 585
R525 B.n429 B.n28 585
R526 B.n428 B.n427 585
R527 B.n426 B.n29 585
R528 B.n425 B.n424 585
R529 B.n423 B.n30 585
R530 B.n422 B.n421 585
R531 B.n420 B.n31 585
R532 B.n419 B.n418 585
R533 B.n417 B.n35 585
R534 B.n416 B.n415 585
R535 B.n414 B.n36 585
R536 B.n413 B.n412 585
R537 B.n411 B.n37 585
R538 B.n410 B.n409 585
R539 B.n407 B.n38 585
R540 B.n406 B.n405 585
R541 B.n404 B.n41 585
R542 B.n403 B.n402 585
R543 B.n401 B.n42 585
R544 B.n400 B.n399 585
R545 B.n398 B.n43 585
R546 B.n397 B.n396 585
R547 B.n395 B.n44 585
R548 B.n394 B.n393 585
R549 B.n392 B.n45 585
R550 B.n391 B.n390 585
R551 B.n389 B.n46 585
R552 B.n388 B.n387 585
R553 B.n386 B.n47 585
R554 B.n385 B.n384 585
R555 B.n383 B.n48 585
R556 B.n382 B.n381 585
R557 B.n450 B.n21 585
R558 B.n452 B.n451 585
R559 B.n453 B.n20 585
R560 B.n455 B.n454 585
R561 B.n456 B.n19 585
R562 B.n458 B.n457 585
R563 B.n459 B.n18 585
R564 B.n461 B.n460 585
R565 B.n462 B.n17 585
R566 B.n464 B.n463 585
R567 B.n465 B.n16 585
R568 B.n467 B.n466 585
R569 B.n468 B.n15 585
R570 B.n470 B.n469 585
R571 B.n471 B.n14 585
R572 B.n473 B.n472 585
R573 B.n474 B.n13 585
R574 B.n476 B.n475 585
R575 B.n477 B.n12 585
R576 B.n479 B.n478 585
R577 B.n480 B.n11 585
R578 B.n482 B.n481 585
R579 B.n483 B.n10 585
R580 B.n485 B.n484 585
R581 B.n486 B.n9 585
R582 B.n488 B.n487 585
R583 B.n489 B.n8 585
R584 B.n491 B.n490 585
R585 B.n492 B.n7 585
R586 B.n494 B.n493 585
R587 B.n495 B.n6 585
R588 B.n497 B.n496 585
R589 B.n498 B.n5 585
R590 B.n500 B.n499 585
R591 B.n501 B.n4 585
R592 B.n503 B.n502 585
R593 B.n504 B.n3 585
R594 B.n506 B.n505 585
R595 B.n507 B.n0 585
R596 B.n2 B.n1 585
R597 B.n135 B.n134 585
R598 B.n137 B.n136 585
R599 B.n138 B.n133 585
R600 B.n140 B.n139 585
R601 B.n141 B.n132 585
R602 B.n143 B.n142 585
R603 B.n144 B.n131 585
R604 B.n146 B.n145 585
R605 B.n147 B.n130 585
R606 B.n149 B.n148 585
R607 B.n150 B.n129 585
R608 B.n152 B.n151 585
R609 B.n153 B.n128 585
R610 B.n155 B.n154 585
R611 B.n156 B.n127 585
R612 B.n158 B.n157 585
R613 B.n159 B.n126 585
R614 B.n161 B.n160 585
R615 B.n162 B.n125 585
R616 B.n164 B.n163 585
R617 B.n165 B.n124 585
R618 B.n167 B.n166 585
R619 B.n168 B.n123 585
R620 B.n170 B.n169 585
R621 B.n171 B.n122 585
R622 B.n173 B.n172 585
R623 B.n174 B.n121 585
R624 B.n176 B.n175 585
R625 B.n177 B.n120 585
R626 B.n179 B.n178 585
R627 B.n180 B.n119 585
R628 B.n182 B.n181 585
R629 B.n183 B.n118 585
R630 B.n185 B.n184 585
R631 B.n186 B.n117 585
R632 B.n188 B.n187 585
R633 B.n189 B.n116 585
R634 B.n191 B.n190 585
R635 B.n192 B.n191 502.111
R636 B.n261 B.n260 502.111
R637 B.n381 B.n380 502.111
R638 B.n448 B.n21 502.111
R639 B.n99 B.t1 283.726
R640 B.n39 B.t5 283.726
R641 B.n105 B.t7 283.726
R642 B.n32 B.t11 283.726
R643 B.n509 B.n508 256.663
R644 B.n105 B.t6 246.357
R645 B.n99 B.t0 246.357
R646 B.n39 B.t3 246.357
R647 B.n32 B.t9 246.357
R648 B.n508 B.n507 235.042
R649 B.n508 B.n2 235.042
R650 B.n100 B.t2 231.556
R651 B.n40 B.t4 231.556
R652 B.n106 B.t8 231.556
R653 B.n33 B.t10 231.556
R654 B.n193 B.n192 163.367
R655 B.n193 B.n114 163.367
R656 B.n197 B.n114 163.367
R657 B.n198 B.n197 163.367
R658 B.n199 B.n198 163.367
R659 B.n199 B.n112 163.367
R660 B.n203 B.n112 163.367
R661 B.n204 B.n203 163.367
R662 B.n205 B.n204 163.367
R663 B.n205 B.n110 163.367
R664 B.n209 B.n110 163.367
R665 B.n210 B.n209 163.367
R666 B.n211 B.n210 163.367
R667 B.n211 B.n108 163.367
R668 B.n215 B.n108 163.367
R669 B.n216 B.n215 163.367
R670 B.n217 B.n216 163.367
R671 B.n217 B.n104 163.367
R672 B.n222 B.n104 163.367
R673 B.n223 B.n222 163.367
R674 B.n224 B.n223 163.367
R675 B.n224 B.n102 163.367
R676 B.n228 B.n102 163.367
R677 B.n229 B.n228 163.367
R678 B.n230 B.n229 163.367
R679 B.n230 B.n98 163.367
R680 B.n235 B.n98 163.367
R681 B.n236 B.n235 163.367
R682 B.n237 B.n236 163.367
R683 B.n237 B.n96 163.367
R684 B.n241 B.n96 163.367
R685 B.n242 B.n241 163.367
R686 B.n243 B.n242 163.367
R687 B.n243 B.n94 163.367
R688 B.n247 B.n94 163.367
R689 B.n248 B.n247 163.367
R690 B.n249 B.n248 163.367
R691 B.n249 B.n92 163.367
R692 B.n253 B.n92 163.367
R693 B.n254 B.n253 163.367
R694 B.n255 B.n254 163.367
R695 B.n255 B.n90 163.367
R696 B.n259 B.n90 163.367
R697 B.n260 B.n259 163.367
R698 B.n380 B.n379 163.367
R699 B.n379 B.n50 163.367
R700 B.n375 B.n50 163.367
R701 B.n375 B.n374 163.367
R702 B.n374 B.n373 163.367
R703 B.n373 B.n52 163.367
R704 B.n369 B.n52 163.367
R705 B.n369 B.n368 163.367
R706 B.n368 B.n367 163.367
R707 B.n367 B.n54 163.367
R708 B.n363 B.n54 163.367
R709 B.n363 B.n362 163.367
R710 B.n362 B.n361 163.367
R711 B.n361 B.n56 163.367
R712 B.n357 B.n56 163.367
R713 B.n357 B.n356 163.367
R714 B.n356 B.n355 163.367
R715 B.n355 B.n58 163.367
R716 B.n351 B.n58 163.367
R717 B.n351 B.n350 163.367
R718 B.n350 B.n349 163.367
R719 B.n349 B.n60 163.367
R720 B.n345 B.n60 163.367
R721 B.n345 B.n344 163.367
R722 B.n344 B.n343 163.367
R723 B.n343 B.n62 163.367
R724 B.n339 B.n62 163.367
R725 B.n339 B.n338 163.367
R726 B.n338 B.n337 163.367
R727 B.n337 B.n64 163.367
R728 B.n333 B.n64 163.367
R729 B.n333 B.n332 163.367
R730 B.n332 B.n331 163.367
R731 B.n331 B.n66 163.367
R732 B.n327 B.n66 163.367
R733 B.n327 B.n326 163.367
R734 B.n326 B.n325 163.367
R735 B.n325 B.n68 163.367
R736 B.n321 B.n68 163.367
R737 B.n321 B.n320 163.367
R738 B.n320 B.n319 163.367
R739 B.n319 B.n70 163.367
R740 B.n315 B.n70 163.367
R741 B.n315 B.n314 163.367
R742 B.n314 B.n313 163.367
R743 B.n313 B.n72 163.367
R744 B.n309 B.n72 163.367
R745 B.n309 B.n308 163.367
R746 B.n308 B.n307 163.367
R747 B.n307 B.n74 163.367
R748 B.n303 B.n74 163.367
R749 B.n303 B.n302 163.367
R750 B.n302 B.n301 163.367
R751 B.n301 B.n76 163.367
R752 B.n297 B.n76 163.367
R753 B.n297 B.n296 163.367
R754 B.n296 B.n295 163.367
R755 B.n295 B.n78 163.367
R756 B.n291 B.n78 163.367
R757 B.n291 B.n290 163.367
R758 B.n290 B.n289 163.367
R759 B.n289 B.n80 163.367
R760 B.n285 B.n80 163.367
R761 B.n285 B.n284 163.367
R762 B.n284 B.n283 163.367
R763 B.n283 B.n82 163.367
R764 B.n279 B.n82 163.367
R765 B.n279 B.n278 163.367
R766 B.n278 B.n277 163.367
R767 B.n277 B.n84 163.367
R768 B.n273 B.n84 163.367
R769 B.n273 B.n272 163.367
R770 B.n272 B.n271 163.367
R771 B.n271 B.n86 163.367
R772 B.n267 B.n86 163.367
R773 B.n267 B.n266 163.367
R774 B.n266 B.n265 163.367
R775 B.n265 B.n88 163.367
R776 B.n261 B.n88 163.367
R777 B.n448 B.n447 163.367
R778 B.n447 B.n446 163.367
R779 B.n446 B.n23 163.367
R780 B.n442 B.n23 163.367
R781 B.n442 B.n441 163.367
R782 B.n441 B.n440 163.367
R783 B.n440 B.n25 163.367
R784 B.n436 B.n25 163.367
R785 B.n436 B.n435 163.367
R786 B.n435 B.n434 163.367
R787 B.n434 B.n27 163.367
R788 B.n430 B.n27 163.367
R789 B.n430 B.n429 163.367
R790 B.n429 B.n428 163.367
R791 B.n428 B.n29 163.367
R792 B.n424 B.n29 163.367
R793 B.n424 B.n423 163.367
R794 B.n423 B.n422 163.367
R795 B.n422 B.n31 163.367
R796 B.n418 B.n31 163.367
R797 B.n418 B.n417 163.367
R798 B.n417 B.n416 163.367
R799 B.n416 B.n36 163.367
R800 B.n412 B.n36 163.367
R801 B.n412 B.n411 163.367
R802 B.n411 B.n410 163.367
R803 B.n410 B.n38 163.367
R804 B.n405 B.n38 163.367
R805 B.n405 B.n404 163.367
R806 B.n404 B.n403 163.367
R807 B.n403 B.n42 163.367
R808 B.n399 B.n42 163.367
R809 B.n399 B.n398 163.367
R810 B.n398 B.n397 163.367
R811 B.n397 B.n44 163.367
R812 B.n393 B.n44 163.367
R813 B.n393 B.n392 163.367
R814 B.n392 B.n391 163.367
R815 B.n391 B.n46 163.367
R816 B.n387 B.n46 163.367
R817 B.n387 B.n386 163.367
R818 B.n386 B.n385 163.367
R819 B.n385 B.n48 163.367
R820 B.n381 B.n48 163.367
R821 B.n452 B.n21 163.367
R822 B.n453 B.n452 163.367
R823 B.n454 B.n453 163.367
R824 B.n454 B.n19 163.367
R825 B.n458 B.n19 163.367
R826 B.n459 B.n458 163.367
R827 B.n460 B.n459 163.367
R828 B.n460 B.n17 163.367
R829 B.n464 B.n17 163.367
R830 B.n465 B.n464 163.367
R831 B.n466 B.n465 163.367
R832 B.n466 B.n15 163.367
R833 B.n470 B.n15 163.367
R834 B.n471 B.n470 163.367
R835 B.n472 B.n471 163.367
R836 B.n472 B.n13 163.367
R837 B.n476 B.n13 163.367
R838 B.n477 B.n476 163.367
R839 B.n478 B.n477 163.367
R840 B.n478 B.n11 163.367
R841 B.n482 B.n11 163.367
R842 B.n483 B.n482 163.367
R843 B.n484 B.n483 163.367
R844 B.n484 B.n9 163.367
R845 B.n488 B.n9 163.367
R846 B.n489 B.n488 163.367
R847 B.n490 B.n489 163.367
R848 B.n490 B.n7 163.367
R849 B.n494 B.n7 163.367
R850 B.n495 B.n494 163.367
R851 B.n496 B.n495 163.367
R852 B.n496 B.n5 163.367
R853 B.n500 B.n5 163.367
R854 B.n501 B.n500 163.367
R855 B.n502 B.n501 163.367
R856 B.n502 B.n3 163.367
R857 B.n506 B.n3 163.367
R858 B.n507 B.n506 163.367
R859 B.n134 B.n2 163.367
R860 B.n137 B.n134 163.367
R861 B.n138 B.n137 163.367
R862 B.n139 B.n138 163.367
R863 B.n139 B.n132 163.367
R864 B.n143 B.n132 163.367
R865 B.n144 B.n143 163.367
R866 B.n145 B.n144 163.367
R867 B.n145 B.n130 163.367
R868 B.n149 B.n130 163.367
R869 B.n150 B.n149 163.367
R870 B.n151 B.n150 163.367
R871 B.n151 B.n128 163.367
R872 B.n155 B.n128 163.367
R873 B.n156 B.n155 163.367
R874 B.n157 B.n156 163.367
R875 B.n157 B.n126 163.367
R876 B.n161 B.n126 163.367
R877 B.n162 B.n161 163.367
R878 B.n163 B.n162 163.367
R879 B.n163 B.n124 163.367
R880 B.n167 B.n124 163.367
R881 B.n168 B.n167 163.367
R882 B.n169 B.n168 163.367
R883 B.n169 B.n122 163.367
R884 B.n173 B.n122 163.367
R885 B.n174 B.n173 163.367
R886 B.n175 B.n174 163.367
R887 B.n175 B.n120 163.367
R888 B.n179 B.n120 163.367
R889 B.n180 B.n179 163.367
R890 B.n181 B.n180 163.367
R891 B.n181 B.n118 163.367
R892 B.n185 B.n118 163.367
R893 B.n186 B.n185 163.367
R894 B.n187 B.n186 163.367
R895 B.n187 B.n116 163.367
R896 B.n191 B.n116 163.367
R897 B.n219 B.n106 59.5399
R898 B.n233 B.n100 59.5399
R899 B.n408 B.n40 59.5399
R900 B.n34 B.n33 59.5399
R901 B.n106 B.n105 52.1702
R902 B.n100 B.n99 52.1702
R903 B.n40 B.n39 52.1702
R904 B.n33 B.n32 52.1702
R905 B.n450 B.n449 32.6249
R906 B.n382 B.n49 32.6249
R907 B.n262 B.n89 32.6249
R908 B.n190 B.n115 32.6249
R909 B B.n509 18.0485
R910 B.n451 B.n450 10.6151
R911 B.n451 B.n20 10.6151
R912 B.n455 B.n20 10.6151
R913 B.n456 B.n455 10.6151
R914 B.n457 B.n456 10.6151
R915 B.n457 B.n18 10.6151
R916 B.n461 B.n18 10.6151
R917 B.n462 B.n461 10.6151
R918 B.n463 B.n462 10.6151
R919 B.n463 B.n16 10.6151
R920 B.n467 B.n16 10.6151
R921 B.n468 B.n467 10.6151
R922 B.n469 B.n468 10.6151
R923 B.n469 B.n14 10.6151
R924 B.n473 B.n14 10.6151
R925 B.n474 B.n473 10.6151
R926 B.n475 B.n474 10.6151
R927 B.n475 B.n12 10.6151
R928 B.n479 B.n12 10.6151
R929 B.n480 B.n479 10.6151
R930 B.n481 B.n480 10.6151
R931 B.n481 B.n10 10.6151
R932 B.n485 B.n10 10.6151
R933 B.n486 B.n485 10.6151
R934 B.n487 B.n486 10.6151
R935 B.n487 B.n8 10.6151
R936 B.n491 B.n8 10.6151
R937 B.n492 B.n491 10.6151
R938 B.n493 B.n492 10.6151
R939 B.n493 B.n6 10.6151
R940 B.n497 B.n6 10.6151
R941 B.n498 B.n497 10.6151
R942 B.n499 B.n498 10.6151
R943 B.n499 B.n4 10.6151
R944 B.n503 B.n4 10.6151
R945 B.n504 B.n503 10.6151
R946 B.n505 B.n504 10.6151
R947 B.n505 B.n0 10.6151
R948 B.n449 B.n22 10.6151
R949 B.n445 B.n22 10.6151
R950 B.n445 B.n444 10.6151
R951 B.n444 B.n443 10.6151
R952 B.n443 B.n24 10.6151
R953 B.n439 B.n24 10.6151
R954 B.n439 B.n438 10.6151
R955 B.n438 B.n437 10.6151
R956 B.n437 B.n26 10.6151
R957 B.n433 B.n26 10.6151
R958 B.n433 B.n432 10.6151
R959 B.n432 B.n431 10.6151
R960 B.n431 B.n28 10.6151
R961 B.n427 B.n28 10.6151
R962 B.n427 B.n426 10.6151
R963 B.n426 B.n425 10.6151
R964 B.n425 B.n30 10.6151
R965 B.n421 B.n420 10.6151
R966 B.n420 B.n419 10.6151
R967 B.n419 B.n35 10.6151
R968 B.n415 B.n35 10.6151
R969 B.n415 B.n414 10.6151
R970 B.n414 B.n413 10.6151
R971 B.n413 B.n37 10.6151
R972 B.n409 B.n37 10.6151
R973 B.n407 B.n406 10.6151
R974 B.n406 B.n41 10.6151
R975 B.n402 B.n41 10.6151
R976 B.n402 B.n401 10.6151
R977 B.n401 B.n400 10.6151
R978 B.n400 B.n43 10.6151
R979 B.n396 B.n43 10.6151
R980 B.n396 B.n395 10.6151
R981 B.n395 B.n394 10.6151
R982 B.n394 B.n45 10.6151
R983 B.n390 B.n45 10.6151
R984 B.n390 B.n389 10.6151
R985 B.n389 B.n388 10.6151
R986 B.n388 B.n47 10.6151
R987 B.n384 B.n47 10.6151
R988 B.n384 B.n383 10.6151
R989 B.n383 B.n382 10.6151
R990 B.n378 B.n49 10.6151
R991 B.n378 B.n377 10.6151
R992 B.n377 B.n376 10.6151
R993 B.n376 B.n51 10.6151
R994 B.n372 B.n51 10.6151
R995 B.n372 B.n371 10.6151
R996 B.n371 B.n370 10.6151
R997 B.n370 B.n53 10.6151
R998 B.n366 B.n53 10.6151
R999 B.n366 B.n365 10.6151
R1000 B.n365 B.n364 10.6151
R1001 B.n364 B.n55 10.6151
R1002 B.n360 B.n55 10.6151
R1003 B.n360 B.n359 10.6151
R1004 B.n359 B.n358 10.6151
R1005 B.n358 B.n57 10.6151
R1006 B.n354 B.n57 10.6151
R1007 B.n354 B.n353 10.6151
R1008 B.n353 B.n352 10.6151
R1009 B.n352 B.n59 10.6151
R1010 B.n348 B.n59 10.6151
R1011 B.n348 B.n347 10.6151
R1012 B.n347 B.n346 10.6151
R1013 B.n346 B.n61 10.6151
R1014 B.n342 B.n61 10.6151
R1015 B.n342 B.n341 10.6151
R1016 B.n341 B.n340 10.6151
R1017 B.n340 B.n63 10.6151
R1018 B.n336 B.n63 10.6151
R1019 B.n336 B.n335 10.6151
R1020 B.n335 B.n334 10.6151
R1021 B.n334 B.n65 10.6151
R1022 B.n330 B.n65 10.6151
R1023 B.n330 B.n329 10.6151
R1024 B.n329 B.n328 10.6151
R1025 B.n328 B.n67 10.6151
R1026 B.n324 B.n67 10.6151
R1027 B.n324 B.n323 10.6151
R1028 B.n323 B.n322 10.6151
R1029 B.n322 B.n69 10.6151
R1030 B.n318 B.n69 10.6151
R1031 B.n318 B.n317 10.6151
R1032 B.n317 B.n316 10.6151
R1033 B.n316 B.n71 10.6151
R1034 B.n312 B.n71 10.6151
R1035 B.n312 B.n311 10.6151
R1036 B.n311 B.n310 10.6151
R1037 B.n310 B.n73 10.6151
R1038 B.n306 B.n73 10.6151
R1039 B.n306 B.n305 10.6151
R1040 B.n305 B.n304 10.6151
R1041 B.n304 B.n75 10.6151
R1042 B.n300 B.n75 10.6151
R1043 B.n300 B.n299 10.6151
R1044 B.n299 B.n298 10.6151
R1045 B.n298 B.n77 10.6151
R1046 B.n294 B.n77 10.6151
R1047 B.n294 B.n293 10.6151
R1048 B.n293 B.n292 10.6151
R1049 B.n292 B.n79 10.6151
R1050 B.n288 B.n79 10.6151
R1051 B.n288 B.n287 10.6151
R1052 B.n287 B.n286 10.6151
R1053 B.n286 B.n81 10.6151
R1054 B.n282 B.n81 10.6151
R1055 B.n282 B.n281 10.6151
R1056 B.n281 B.n280 10.6151
R1057 B.n280 B.n83 10.6151
R1058 B.n276 B.n83 10.6151
R1059 B.n276 B.n275 10.6151
R1060 B.n275 B.n274 10.6151
R1061 B.n274 B.n85 10.6151
R1062 B.n270 B.n85 10.6151
R1063 B.n270 B.n269 10.6151
R1064 B.n269 B.n268 10.6151
R1065 B.n268 B.n87 10.6151
R1066 B.n264 B.n87 10.6151
R1067 B.n264 B.n263 10.6151
R1068 B.n263 B.n262 10.6151
R1069 B.n135 B.n1 10.6151
R1070 B.n136 B.n135 10.6151
R1071 B.n136 B.n133 10.6151
R1072 B.n140 B.n133 10.6151
R1073 B.n141 B.n140 10.6151
R1074 B.n142 B.n141 10.6151
R1075 B.n142 B.n131 10.6151
R1076 B.n146 B.n131 10.6151
R1077 B.n147 B.n146 10.6151
R1078 B.n148 B.n147 10.6151
R1079 B.n148 B.n129 10.6151
R1080 B.n152 B.n129 10.6151
R1081 B.n153 B.n152 10.6151
R1082 B.n154 B.n153 10.6151
R1083 B.n154 B.n127 10.6151
R1084 B.n158 B.n127 10.6151
R1085 B.n159 B.n158 10.6151
R1086 B.n160 B.n159 10.6151
R1087 B.n160 B.n125 10.6151
R1088 B.n164 B.n125 10.6151
R1089 B.n165 B.n164 10.6151
R1090 B.n166 B.n165 10.6151
R1091 B.n166 B.n123 10.6151
R1092 B.n170 B.n123 10.6151
R1093 B.n171 B.n170 10.6151
R1094 B.n172 B.n171 10.6151
R1095 B.n172 B.n121 10.6151
R1096 B.n176 B.n121 10.6151
R1097 B.n177 B.n176 10.6151
R1098 B.n178 B.n177 10.6151
R1099 B.n178 B.n119 10.6151
R1100 B.n182 B.n119 10.6151
R1101 B.n183 B.n182 10.6151
R1102 B.n184 B.n183 10.6151
R1103 B.n184 B.n117 10.6151
R1104 B.n188 B.n117 10.6151
R1105 B.n189 B.n188 10.6151
R1106 B.n190 B.n189 10.6151
R1107 B.n194 B.n115 10.6151
R1108 B.n195 B.n194 10.6151
R1109 B.n196 B.n195 10.6151
R1110 B.n196 B.n113 10.6151
R1111 B.n200 B.n113 10.6151
R1112 B.n201 B.n200 10.6151
R1113 B.n202 B.n201 10.6151
R1114 B.n202 B.n111 10.6151
R1115 B.n206 B.n111 10.6151
R1116 B.n207 B.n206 10.6151
R1117 B.n208 B.n207 10.6151
R1118 B.n208 B.n109 10.6151
R1119 B.n212 B.n109 10.6151
R1120 B.n213 B.n212 10.6151
R1121 B.n214 B.n213 10.6151
R1122 B.n214 B.n107 10.6151
R1123 B.n218 B.n107 10.6151
R1124 B.n221 B.n220 10.6151
R1125 B.n221 B.n103 10.6151
R1126 B.n225 B.n103 10.6151
R1127 B.n226 B.n225 10.6151
R1128 B.n227 B.n226 10.6151
R1129 B.n227 B.n101 10.6151
R1130 B.n231 B.n101 10.6151
R1131 B.n232 B.n231 10.6151
R1132 B.n234 B.n97 10.6151
R1133 B.n238 B.n97 10.6151
R1134 B.n239 B.n238 10.6151
R1135 B.n240 B.n239 10.6151
R1136 B.n240 B.n95 10.6151
R1137 B.n244 B.n95 10.6151
R1138 B.n245 B.n244 10.6151
R1139 B.n246 B.n245 10.6151
R1140 B.n246 B.n93 10.6151
R1141 B.n250 B.n93 10.6151
R1142 B.n251 B.n250 10.6151
R1143 B.n252 B.n251 10.6151
R1144 B.n252 B.n91 10.6151
R1145 B.n256 B.n91 10.6151
R1146 B.n257 B.n256 10.6151
R1147 B.n258 B.n257 10.6151
R1148 B.n258 B.n89 10.6151
R1149 B.n509 B.n0 8.11757
R1150 B.n509 B.n1 8.11757
R1151 B.n421 B.n34 6.5566
R1152 B.n409 B.n408 6.5566
R1153 B.n220 B.n219 6.5566
R1154 B.n233 B.n232 6.5566
R1155 B.n34 B.n30 4.05904
R1156 B.n408 B.n407 4.05904
R1157 B.n219 B.n218 4.05904
R1158 B.n234 B.n233 4.05904
C0 B VN 1.03207f
C1 VDD2 VN 2.34363f
C2 VDD2 B 1.45346f
C3 w_n3122_n1726# VP 6.11271f
C4 VDD1 w_n3122_n1726# 1.65909f
C5 w_n3122_n1726# VTAIL 1.78234f
C6 VP VN 5.18198f
C7 B VP 1.70341f
C8 VDD1 VN 0.154877f
C9 VTAIL VN 2.97056f
C10 VDD1 B 1.38497f
C11 B VTAIL 1.74846f
C12 VDD2 VP 0.442288f
C13 VDD1 VDD2 1.31285f
C14 VDD2 VTAIL 4.66219f
C15 VDD1 VP 2.6287f
C16 VTAIL VP 2.98473f
C17 VDD1 VTAIL 4.61115f
C18 w_n3122_n1726# VN 5.71091f
C19 B w_n3122_n1726# 7.05908f
C20 VDD2 w_n3122_n1726# 1.73614f
C21 VDD2 VSUBS 1.281737f
C22 VDD1 VSUBS 1.409532f
C23 VTAIL VSUBS 0.545587f
C24 VN VSUBS 5.34925f
C25 VP VSUBS 2.245112f
C26 B VSUBS 3.493625f
C27 w_n3122_n1726# VSUBS 67.9222f
C28 B.n0 VSUBS 0.006354f
C29 B.n1 VSUBS 0.006354f
C30 B.n2 VSUBS 0.009398f
C31 B.n3 VSUBS 0.007202f
C32 B.n4 VSUBS 0.007202f
C33 B.n5 VSUBS 0.007202f
C34 B.n6 VSUBS 0.007202f
C35 B.n7 VSUBS 0.007202f
C36 B.n8 VSUBS 0.007202f
C37 B.n9 VSUBS 0.007202f
C38 B.n10 VSUBS 0.007202f
C39 B.n11 VSUBS 0.007202f
C40 B.n12 VSUBS 0.007202f
C41 B.n13 VSUBS 0.007202f
C42 B.n14 VSUBS 0.007202f
C43 B.n15 VSUBS 0.007202f
C44 B.n16 VSUBS 0.007202f
C45 B.n17 VSUBS 0.007202f
C46 B.n18 VSUBS 0.007202f
C47 B.n19 VSUBS 0.007202f
C48 B.n20 VSUBS 0.007202f
C49 B.n21 VSUBS 0.016081f
C50 B.n22 VSUBS 0.007202f
C51 B.n23 VSUBS 0.007202f
C52 B.n24 VSUBS 0.007202f
C53 B.n25 VSUBS 0.007202f
C54 B.n26 VSUBS 0.007202f
C55 B.n27 VSUBS 0.007202f
C56 B.n28 VSUBS 0.007202f
C57 B.n29 VSUBS 0.007202f
C58 B.n30 VSUBS 0.004978f
C59 B.n31 VSUBS 0.007202f
C60 B.t10 VSUBS 0.056035f
C61 B.t11 VSUBS 0.075062f
C62 B.t9 VSUBS 0.442147f
C63 B.n32 VSUBS 0.132941f
C64 B.n33 VSUBS 0.113751f
C65 B.n34 VSUBS 0.016685f
C66 B.n35 VSUBS 0.007202f
C67 B.n36 VSUBS 0.007202f
C68 B.n37 VSUBS 0.007202f
C69 B.n38 VSUBS 0.007202f
C70 B.t4 VSUBS 0.056036f
C71 B.t5 VSUBS 0.075063f
C72 B.t3 VSUBS 0.442147f
C73 B.n39 VSUBS 0.13294f
C74 B.n40 VSUBS 0.11375f
C75 B.n41 VSUBS 0.007202f
C76 B.n42 VSUBS 0.007202f
C77 B.n43 VSUBS 0.007202f
C78 B.n44 VSUBS 0.007202f
C79 B.n45 VSUBS 0.007202f
C80 B.n46 VSUBS 0.007202f
C81 B.n47 VSUBS 0.007202f
C82 B.n48 VSUBS 0.007202f
C83 B.n49 VSUBS 0.016081f
C84 B.n50 VSUBS 0.007202f
C85 B.n51 VSUBS 0.007202f
C86 B.n52 VSUBS 0.007202f
C87 B.n53 VSUBS 0.007202f
C88 B.n54 VSUBS 0.007202f
C89 B.n55 VSUBS 0.007202f
C90 B.n56 VSUBS 0.007202f
C91 B.n57 VSUBS 0.007202f
C92 B.n58 VSUBS 0.007202f
C93 B.n59 VSUBS 0.007202f
C94 B.n60 VSUBS 0.007202f
C95 B.n61 VSUBS 0.007202f
C96 B.n62 VSUBS 0.007202f
C97 B.n63 VSUBS 0.007202f
C98 B.n64 VSUBS 0.007202f
C99 B.n65 VSUBS 0.007202f
C100 B.n66 VSUBS 0.007202f
C101 B.n67 VSUBS 0.007202f
C102 B.n68 VSUBS 0.007202f
C103 B.n69 VSUBS 0.007202f
C104 B.n70 VSUBS 0.007202f
C105 B.n71 VSUBS 0.007202f
C106 B.n72 VSUBS 0.007202f
C107 B.n73 VSUBS 0.007202f
C108 B.n74 VSUBS 0.007202f
C109 B.n75 VSUBS 0.007202f
C110 B.n76 VSUBS 0.007202f
C111 B.n77 VSUBS 0.007202f
C112 B.n78 VSUBS 0.007202f
C113 B.n79 VSUBS 0.007202f
C114 B.n80 VSUBS 0.007202f
C115 B.n81 VSUBS 0.007202f
C116 B.n82 VSUBS 0.007202f
C117 B.n83 VSUBS 0.007202f
C118 B.n84 VSUBS 0.007202f
C119 B.n85 VSUBS 0.007202f
C120 B.n86 VSUBS 0.007202f
C121 B.n87 VSUBS 0.007202f
C122 B.n88 VSUBS 0.007202f
C123 B.n89 VSUBS 0.016746f
C124 B.n90 VSUBS 0.007202f
C125 B.n91 VSUBS 0.007202f
C126 B.n92 VSUBS 0.007202f
C127 B.n93 VSUBS 0.007202f
C128 B.n94 VSUBS 0.007202f
C129 B.n95 VSUBS 0.007202f
C130 B.n96 VSUBS 0.007202f
C131 B.n97 VSUBS 0.007202f
C132 B.n98 VSUBS 0.007202f
C133 B.t2 VSUBS 0.056036f
C134 B.t1 VSUBS 0.075063f
C135 B.t0 VSUBS 0.442147f
C136 B.n99 VSUBS 0.13294f
C137 B.n100 VSUBS 0.11375f
C138 B.n101 VSUBS 0.007202f
C139 B.n102 VSUBS 0.007202f
C140 B.n103 VSUBS 0.007202f
C141 B.n104 VSUBS 0.007202f
C142 B.t8 VSUBS 0.056035f
C143 B.t7 VSUBS 0.075062f
C144 B.t6 VSUBS 0.442147f
C145 B.n105 VSUBS 0.132941f
C146 B.n106 VSUBS 0.113751f
C147 B.n107 VSUBS 0.007202f
C148 B.n108 VSUBS 0.007202f
C149 B.n109 VSUBS 0.007202f
C150 B.n110 VSUBS 0.007202f
C151 B.n111 VSUBS 0.007202f
C152 B.n112 VSUBS 0.007202f
C153 B.n113 VSUBS 0.007202f
C154 B.n114 VSUBS 0.007202f
C155 B.n115 VSUBS 0.017597f
C156 B.n116 VSUBS 0.007202f
C157 B.n117 VSUBS 0.007202f
C158 B.n118 VSUBS 0.007202f
C159 B.n119 VSUBS 0.007202f
C160 B.n120 VSUBS 0.007202f
C161 B.n121 VSUBS 0.007202f
C162 B.n122 VSUBS 0.007202f
C163 B.n123 VSUBS 0.007202f
C164 B.n124 VSUBS 0.007202f
C165 B.n125 VSUBS 0.007202f
C166 B.n126 VSUBS 0.007202f
C167 B.n127 VSUBS 0.007202f
C168 B.n128 VSUBS 0.007202f
C169 B.n129 VSUBS 0.007202f
C170 B.n130 VSUBS 0.007202f
C171 B.n131 VSUBS 0.007202f
C172 B.n132 VSUBS 0.007202f
C173 B.n133 VSUBS 0.007202f
C174 B.n134 VSUBS 0.007202f
C175 B.n135 VSUBS 0.007202f
C176 B.n136 VSUBS 0.007202f
C177 B.n137 VSUBS 0.007202f
C178 B.n138 VSUBS 0.007202f
C179 B.n139 VSUBS 0.007202f
C180 B.n140 VSUBS 0.007202f
C181 B.n141 VSUBS 0.007202f
C182 B.n142 VSUBS 0.007202f
C183 B.n143 VSUBS 0.007202f
C184 B.n144 VSUBS 0.007202f
C185 B.n145 VSUBS 0.007202f
C186 B.n146 VSUBS 0.007202f
C187 B.n147 VSUBS 0.007202f
C188 B.n148 VSUBS 0.007202f
C189 B.n149 VSUBS 0.007202f
C190 B.n150 VSUBS 0.007202f
C191 B.n151 VSUBS 0.007202f
C192 B.n152 VSUBS 0.007202f
C193 B.n153 VSUBS 0.007202f
C194 B.n154 VSUBS 0.007202f
C195 B.n155 VSUBS 0.007202f
C196 B.n156 VSUBS 0.007202f
C197 B.n157 VSUBS 0.007202f
C198 B.n158 VSUBS 0.007202f
C199 B.n159 VSUBS 0.007202f
C200 B.n160 VSUBS 0.007202f
C201 B.n161 VSUBS 0.007202f
C202 B.n162 VSUBS 0.007202f
C203 B.n163 VSUBS 0.007202f
C204 B.n164 VSUBS 0.007202f
C205 B.n165 VSUBS 0.007202f
C206 B.n166 VSUBS 0.007202f
C207 B.n167 VSUBS 0.007202f
C208 B.n168 VSUBS 0.007202f
C209 B.n169 VSUBS 0.007202f
C210 B.n170 VSUBS 0.007202f
C211 B.n171 VSUBS 0.007202f
C212 B.n172 VSUBS 0.007202f
C213 B.n173 VSUBS 0.007202f
C214 B.n174 VSUBS 0.007202f
C215 B.n175 VSUBS 0.007202f
C216 B.n176 VSUBS 0.007202f
C217 B.n177 VSUBS 0.007202f
C218 B.n178 VSUBS 0.007202f
C219 B.n179 VSUBS 0.007202f
C220 B.n180 VSUBS 0.007202f
C221 B.n181 VSUBS 0.007202f
C222 B.n182 VSUBS 0.007202f
C223 B.n183 VSUBS 0.007202f
C224 B.n184 VSUBS 0.007202f
C225 B.n185 VSUBS 0.007202f
C226 B.n186 VSUBS 0.007202f
C227 B.n187 VSUBS 0.007202f
C228 B.n188 VSUBS 0.007202f
C229 B.n189 VSUBS 0.007202f
C230 B.n190 VSUBS 0.016081f
C231 B.n191 VSUBS 0.016081f
C232 B.n192 VSUBS 0.017597f
C233 B.n193 VSUBS 0.007202f
C234 B.n194 VSUBS 0.007202f
C235 B.n195 VSUBS 0.007202f
C236 B.n196 VSUBS 0.007202f
C237 B.n197 VSUBS 0.007202f
C238 B.n198 VSUBS 0.007202f
C239 B.n199 VSUBS 0.007202f
C240 B.n200 VSUBS 0.007202f
C241 B.n201 VSUBS 0.007202f
C242 B.n202 VSUBS 0.007202f
C243 B.n203 VSUBS 0.007202f
C244 B.n204 VSUBS 0.007202f
C245 B.n205 VSUBS 0.007202f
C246 B.n206 VSUBS 0.007202f
C247 B.n207 VSUBS 0.007202f
C248 B.n208 VSUBS 0.007202f
C249 B.n209 VSUBS 0.007202f
C250 B.n210 VSUBS 0.007202f
C251 B.n211 VSUBS 0.007202f
C252 B.n212 VSUBS 0.007202f
C253 B.n213 VSUBS 0.007202f
C254 B.n214 VSUBS 0.007202f
C255 B.n215 VSUBS 0.007202f
C256 B.n216 VSUBS 0.007202f
C257 B.n217 VSUBS 0.007202f
C258 B.n218 VSUBS 0.004978f
C259 B.n219 VSUBS 0.016685f
C260 B.n220 VSUBS 0.005825f
C261 B.n221 VSUBS 0.007202f
C262 B.n222 VSUBS 0.007202f
C263 B.n223 VSUBS 0.007202f
C264 B.n224 VSUBS 0.007202f
C265 B.n225 VSUBS 0.007202f
C266 B.n226 VSUBS 0.007202f
C267 B.n227 VSUBS 0.007202f
C268 B.n228 VSUBS 0.007202f
C269 B.n229 VSUBS 0.007202f
C270 B.n230 VSUBS 0.007202f
C271 B.n231 VSUBS 0.007202f
C272 B.n232 VSUBS 0.005825f
C273 B.n233 VSUBS 0.016685f
C274 B.n234 VSUBS 0.004978f
C275 B.n235 VSUBS 0.007202f
C276 B.n236 VSUBS 0.007202f
C277 B.n237 VSUBS 0.007202f
C278 B.n238 VSUBS 0.007202f
C279 B.n239 VSUBS 0.007202f
C280 B.n240 VSUBS 0.007202f
C281 B.n241 VSUBS 0.007202f
C282 B.n242 VSUBS 0.007202f
C283 B.n243 VSUBS 0.007202f
C284 B.n244 VSUBS 0.007202f
C285 B.n245 VSUBS 0.007202f
C286 B.n246 VSUBS 0.007202f
C287 B.n247 VSUBS 0.007202f
C288 B.n248 VSUBS 0.007202f
C289 B.n249 VSUBS 0.007202f
C290 B.n250 VSUBS 0.007202f
C291 B.n251 VSUBS 0.007202f
C292 B.n252 VSUBS 0.007202f
C293 B.n253 VSUBS 0.007202f
C294 B.n254 VSUBS 0.007202f
C295 B.n255 VSUBS 0.007202f
C296 B.n256 VSUBS 0.007202f
C297 B.n257 VSUBS 0.007202f
C298 B.n258 VSUBS 0.007202f
C299 B.n259 VSUBS 0.007202f
C300 B.n260 VSUBS 0.017597f
C301 B.n261 VSUBS 0.016081f
C302 B.n262 VSUBS 0.016933f
C303 B.n263 VSUBS 0.007202f
C304 B.n264 VSUBS 0.007202f
C305 B.n265 VSUBS 0.007202f
C306 B.n266 VSUBS 0.007202f
C307 B.n267 VSUBS 0.007202f
C308 B.n268 VSUBS 0.007202f
C309 B.n269 VSUBS 0.007202f
C310 B.n270 VSUBS 0.007202f
C311 B.n271 VSUBS 0.007202f
C312 B.n272 VSUBS 0.007202f
C313 B.n273 VSUBS 0.007202f
C314 B.n274 VSUBS 0.007202f
C315 B.n275 VSUBS 0.007202f
C316 B.n276 VSUBS 0.007202f
C317 B.n277 VSUBS 0.007202f
C318 B.n278 VSUBS 0.007202f
C319 B.n279 VSUBS 0.007202f
C320 B.n280 VSUBS 0.007202f
C321 B.n281 VSUBS 0.007202f
C322 B.n282 VSUBS 0.007202f
C323 B.n283 VSUBS 0.007202f
C324 B.n284 VSUBS 0.007202f
C325 B.n285 VSUBS 0.007202f
C326 B.n286 VSUBS 0.007202f
C327 B.n287 VSUBS 0.007202f
C328 B.n288 VSUBS 0.007202f
C329 B.n289 VSUBS 0.007202f
C330 B.n290 VSUBS 0.007202f
C331 B.n291 VSUBS 0.007202f
C332 B.n292 VSUBS 0.007202f
C333 B.n293 VSUBS 0.007202f
C334 B.n294 VSUBS 0.007202f
C335 B.n295 VSUBS 0.007202f
C336 B.n296 VSUBS 0.007202f
C337 B.n297 VSUBS 0.007202f
C338 B.n298 VSUBS 0.007202f
C339 B.n299 VSUBS 0.007202f
C340 B.n300 VSUBS 0.007202f
C341 B.n301 VSUBS 0.007202f
C342 B.n302 VSUBS 0.007202f
C343 B.n303 VSUBS 0.007202f
C344 B.n304 VSUBS 0.007202f
C345 B.n305 VSUBS 0.007202f
C346 B.n306 VSUBS 0.007202f
C347 B.n307 VSUBS 0.007202f
C348 B.n308 VSUBS 0.007202f
C349 B.n309 VSUBS 0.007202f
C350 B.n310 VSUBS 0.007202f
C351 B.n311 VSUBS 0.007202f
C352 B.n312 VSUBS 0.007202f
C353 B.n313 VSUBS 0.007202f
C354 B.n314 VSUBS 0.007202f
C355 B.n315 VSUBS 0.007202f
C356 B.n316 VSUBS 0.007202f
C357 B.n317 VSUBS 0.007202f
C358 B.n318 VSUBS 0.007202f
C359 B.n319 VSUBS 0.007202f
C360 B.n320 VSUBS 0.007202f
C361 B.n321 VSUBS 0.007202f
C362 B.n322 VSUBS 0.007202f
C363 B.n323 VSUBS 0.007202f
C364 B.n324 VSUBS 0.007202f
C365 B.n325 VSUBS 0.007202f
C366 B.n326 VSUBS 0.007202f
C367 B.n327 VSUBS 0.007202f
C368 B.n328 VSUBS 0.007202f
C369 B.n329 VSUBS 0.007202f
C370 B.n330 VSUBS 0.007202f
C371 B.n331 VSUBS 0.007202f
C372 B.n332 VSUBS 0.007202f
C373 B.n333 VSUBS 0.007202f
C374 B.n334 VSUBS 0.007202f
C375 B.n335 VSUBS 0.007202f
C376 B.n336 VSUBS 0.007202f
C377 B.n337 VSUBS 0.007202f
C378 B.n338 VSUBS 0.007202f
C379 B.n339 VSUBS 0.007202f
C380 B.n340 VSUBS 0.007202f
C381 B.n341 VSUBS 0.007202f
C382 B.n342 VSUBS 0.007202f
C383 B.n343 VSUBS 0.007202f
C384 B.n344 VSUBS 0.007202f
C385 B.n345 VSUBS 0.007202f
C386 B.n346 VSUBS 0.007202f
C387 B.n347 VSUBS 0.007202f
C388 B.n348 VSUBS 0.007202f
C389 B.n349 VSUBS 0.007202f
C390 B.n350 VSUBS 0.007202f
C391 B.n351 VSUBS 0.007202f
C392 B.n352 VSUBS 0.007202f
C393 B.n353 VSUBS 0.007202f
C394 B.n354 VSUBS 0.007202f
C395 B.n355 VSUBS 0.007202f
C396 B.n356 VSUBS 0.007202f
C397 B.n357 VSUBS 0.007202f
C398 B.n358 VSUBS 0.007202f
C399 B.n359 VSUBS 0.007202f
C400 B.n360 VSUBS 0.007202f
C401 B.n361 VSUBS 0.007202f
C402 B.n362 VSUBS 0.007202f
C403 B.n363 VSUBS 0.007202f
C404 B.n364 VSUBS 0.007202f
C405 B.n365 VSUBS 0.007202f
C406 B.n366 VSUBS 0.007202f
C407 B.n367 VSUBS 0.007202f
C408 B.n368 VSUBS 0.007202f
C409 B.n369 VSUBS 0.007202f
C410 B.n370 VSUBS 0.007202f
C411 B.n371 VSUBS 0.007202f
C412 B.n372 VSUBS 0.007202f
C413 B.n373 VSUBS 0.007202f
C414 B.n374 VSUBS 0.007202f
C415 B.n375 VSUBS 0.007202f
C416 B.n376 VSUBS 0.007202f
C417 B.n377 VSUBS 0.007202f
C418 B.n378 VSUBS 0.007202f
C419 B.n379 VSUBS 0.007202f
C420 B.n380 VSUBS 0.016081f
C421 B.n381 VSUBS 0.017597f
C422 B.n382 VSUBS 0.017597f
C423 B.n383 VSUBS 0.007202f
C424 B.n384 VSUBS 0.007202f
C425 B.n385 VSUBS 0.007202f
C426 B.n386 VSUBS 0.007202f
C427 B.n387 VSUBS 0.007202f
C428 B.n388 VSUBS 0.007202f
C429 B.n389 VSUBS 0.007202f
C430 B.n390 VSUBS 0.007202f
C431 B.n391 VSUBS 0.007202f
C432 B.n392 VSUBS 0.007202f
C433 B.n393 VSUBS 0.007202f
C434 B.n394 VSUBS 0.007202f
C435 B.n395 VSUBS 0.007202f
C436 B.n396 VSUBS 0.007202f
C437 B.n397 VSUBS 0.007202f
C438 B.n398 VSUBS 0.007202f
C439 B.n399 VSUBS 0.007202f
C440 B.n400 VSUBS 0.007202f
C441 B.n401 VSUBS 0.007202f
C442 B.n402 VSUBS 0.007202f
C443 B.n403 VSUBS 0.007202f
C444 B.n404 VSUBS 0.007202f
C445 B.n405 VSUBS 0.007202f
C446 B.n406 VSUBS 0.007202f
C447 B.n407 VSUBS 0.004978f
C448 B.n408 VSUBS 0.016685f
C449 B.n409 VSUBS 0.005825f
C450 B.n410 VSUBS 0.007202f
C451 B.n411 VSUBS 0.007202f
C452 B.n412 VSUBS 0.007202f
C453 B.n413 VSUBS 0.007202f
C454 B.n414 VSUBS 0.007202f
C455 B.n415 VSUBS 0.007202f
C456 B.n416 VSUBS 0.007202f
C457 B.n417 VSUBS 0.007202f
C458 B.n418 VSUBS 0.007202f
C459 B.n419 VSUBS 0.007202f
C460 B.n420 VSUBS 0.007202f
C461 B.n421 VSUBS 0.005825f
C462 B.n422 VSUBS 0.007202f
C463 B.n423 VSUBS 0.007202f
C464 B.n424 VSUBS 0.007202f
C465 B.n425 VSUBS 0.007202f
C466 B.n426 VSUBS 0.007202f
C467 B.n427 VSUBS 0.007202f
C468 B.n428 VSUBS 0.007202f
C469 B.n429 VSUBS 0.007202f
C470 B.n430 VSUBS 0.007202f
C471 B.n431 VSUBS 0.007202f
C472 B.n432 VSUBS 0.007202f
C473 B.n433 VSUBS 0.007202f
C474 B.n434 VSUBS 0.007202f
C475 B.n435 VSUBS 0.007202f
C476 B.n436 VSUBS 0.007202f
C477 B.n437 VSUBS 0.007202f
C478 B.n438 VSUBS 0.007202f
C479 B.n439 VSUBS 0.007202f
C480 B.n440 VSUBS 0.007202f
C481 B.n441 VSUBS 0.007202f
C482 B.n442 VSUBS 0.007202f
C483 B.n443 VSUBS 0.007202f
C484 B.n444 VSUBS 0.007202f
C485 B.n445 VSUBS 0.007202f
C486 B.n446 VSUBS 0.007202f
C487 B.n447 VSUBS 0.007202f
C488 B.n448 VSUBS 0.017597f
C489 B.n449 VSUBS 0.017597f
C490 B.n450 VSUBS 0.016081f
C491 B.n451 VSUBS 0.007202f
C492 B.n452 VSUBS 0.007202f
C493 B.n453 VSUBS 0.007202f
C494 B.n454 VSUBS 0.007202f
C495 B.n455 VSUBS 0.007202f
C496 B.n456 VSUBS 0.007202f
C497 B.n457 VSUBS 0.007202f
C498 B.n458 VSUBS 0.007202f
C499 B.n459 VSUBS 0.007202f
C500 B.n460 VSUBS 0.007202f
C501 B.n461 VSUBS 0.007202f
C502 B.n462 VSUBS 0.007202f
C503 B.n463 VSUBS 0.007202f
C504 B.n464 VSUBS 0.007202f
C505 B.n465 VSUBS 0.007202f
C506 B.n466 VSUBS 0.007202f
C507 B.n467 VSUBS 0.007202f
C508 B.n468 VSUBS 0.007202f
C509 B.n469 VSUBS 0.007202f
C510 B.n470 VSUBS 0.007202f
C511 B.n471 VSUBS 0.007202f
C512 B.n472 VSUBS 0.007202f
C513 B.n473 VSUBS 0.007202f
C514 B.n474 VSUBS 0.007202f
C515 B.n475 VSUBS 0.007202f
C516 B.n476 VSUBS 0.007202f
C517 B.n477 VSUBS 0.007202f
C518 B.n478 VSUBS 0.007202f
C519 B.n479 VSUBS 0.007202f
C520 B.n480 VSUBS 0.007202f
C521 B.n481 VSUBS 0.007202f
C522 B.n482 VSUBS 0.007202f
C523 B.n483 VSUBS 0.007202f
C524 B.n484 VSUBS 0.007202f
C525 B.n485 VSUBS 0.007202f
C526 B.n486 VSUBS 0.007202f
C527 B.n487 VSUBS 0.007202f
C528 B.n488 VSUBS 0.007202f
C529 B.n489 VSUBS 0.007202f
C530 B.n490 VSUBS 0.007202f
C531 B.n491 VSUBS 0.007202f
C532 B.n492 VSUBS 0.007202f
C533 B.n493 VSUBS 0.007202f
C534 B.n494 VSUBS 0.007202f
C535 B.n495 VSUBS 0.007202f
C536 B.n496 VSUBS 0.007202f
C537 B.n497 VSUBS 0.007202f
C538 B.n498 VSUBS 0.007202f
C539 B.n499 VSUBS 0.007202f
C540 B.n500 VSUBS 0.007202f
C541 B.n501 VSUBS 0.007202f
C542 B.n502 VSUBS 0.007202f
C543 B.n503 VSUBS 0.007202f
C544 B.n504 VSUBS 0.007202f
C545 B.n505 VSUBS 0.007202f
C546 B.n506 VSUBS 0.007202f
C547 B.n507 VSUBS 0.009398f
C548 B.n508 VSUBS 0.010011f
C549 B.n509 VSUBS 0.019908f
C550 VDD2.n0 VSUBS 0.022664f
C551 VDD2.n1 VSUBS 0.022164f
C552 VDD2.n2 VSUBS 0.01191f
C553 VDD2.n3 VSUBS 0.028151f
C554 VDD2.n4 VSUBS 0.012611f
C555 VDD2.n5 VSUBS 0.083981f
C556 VDD2.t4 VSUBS 0.061351f
C557 VDD2.n6 VSUBS 0.021113f
C558 VDD2.n7 VSUBS 0.017707f
C559 VDD2.n8 VSUBS 0.01191f
C560 VDD2.n9 VSUBS 0.28476f
C561 VDD2.n10 VSUBS 0.022164f
C562 VDD2.n11 VSUBS 0.01191f
C563 VDD2.n12 VSUBS 0.012611f
C564 VDD2.n13 VSUBS 0.028151f
C565 VDD2.n14 VSUBS 0.062395f
C566 VDD2.n15 VSUBS 0.012611f
C567 VDD2.n16 VSUBS 0.01191f
C568 VDD2.n17 VSUBS 0.049718f
C569 VDD2.n18 VSUBS 0.051907f
C570 VDD2.t3 VSUBS 0.066382f
C571 VDD2.t0 VSUBS 0.066382f
C572 VDD2.n19 VSUBS 0.383324f
C573 VDD2.n20 VSUBS 1.97066f
C574 VDD2.n21 VSUBS 0.022664f
C575 VDD2.n22 VSUBS 0.022164f
C576 VDD2.n23 VSUBS 0.01191f
C577 VDD2.n24 VSUBS 0.028151f
C578 VDD2.n25 VSUBS 0.012611f
C579 VDD2.n26 VSUBS 0.083981f
C580 VDD2.t5 VSUBS 0.061351f
C581 VDD2.n27 VSUBS 0.021113f
C582 VDD2.n28 VSUBS 0.017707f
C583 VDD2.n29 VSUBS 0.01191f
C584 VDD2.n30 VSUBS 0.28476f
C585 VDD2.n31 VSUBS 0.022164f
C586 VDD2.n32 VSUBS 0.01191f
C587 VDD2.n33 VSUBS 0.012611f
C588 VDD2.n34 VSUBS 0.028151f
C589 VDD2.n35 VSUBS 0.062395f
C590 VDD2.n36 VSUBS 0.012611f
C591 VDD2.n37 VSUBS 0.01191f
C592 VDD2.n38 VSUBS 0.049718f
C593 VDD2.n39 VSUBS 0.046392f
C594 VDD2.n40 VSUBS 1.63717f
C595 VDD2.t1 VSUBS 0.066382f
C596 VDD2.t2 VSUBS 0.066382f
C597 VDD2.n41 VSUBS 0.383305f
C598 VN.n0 VSUBS 0.060597f
C599 VN.t5 VSUBS 1.05079f
C600 VN.n1 VSUBS 0.053616f
C601 VN.n2 VSUBS 0.433046f
C602 VN.t2 VSUBS 1.05079f
C603 VN.t1 VSUBS 1.37161f
C604 VN.n3 VSUBS 0.52671f
C605 VN.n4 VSUBS 0.576443f
C606 VN.n5 VSUBS 0.085663f
C607 VN.n6 VSUBS 0.079037f
C608 VN.n7 VSUBS 0.045963f
C609 VN.n8 VSUBS 0.045963f
C610 VN.n9 VSUBS 0.045963f
C611 VN.n10 VSUBS 0.087213f
C612 VN.n11 VSUBS 0.059442f
C613 VN.n12 VSUBS 0.563768f
C614 VN.n13 VSUBS 0.072064f
C615 VN.n14 VSUBS 0.060597f
C616 VN.t0 VSUBS 1.05079f
C617 VN.n15 VSUBS 0.053616f
C618 VN.n16 VSUBS 0.433046f
C619 VN.t4 VSUBS 1.05079f
C620 VN.t3 VSUBS 1.37161f
C621 VN.n17 VSUBS 0.52671f
C622 VN.n18 VSUBS 0.576443f
C623 VN.n19 VSUBS 0.085663f
C624 VN.n20 VSUBS 0.079037f
C625 VN.n21 VSUBS 0.045963f
C626 VN.n22 VSUBS 0.045963f
C627 VN.n23 VSUBS 0.045963f
C628 VN.n24 VSUBS 0.087213f
C629 VN.n25 VSUBS 0.059442f
C630 VN.n26 VSUBS 0.563768f
C631 VN.n27 VSUBS 1.93667f
C632 VTAIL.t2 VSUBS 0.088778f
C633 VTAIL.t3 VSUBS 0.088778f
C634 VTAIL.n0 VSUBS 0.438989f
C635 VTAIL.n1 VSUBS 0.657437f
C636 VTAIL.n2 VSUBS 0.03031f
C637 VTAIL.n3 VSUBS 0.029642f
C638 VTAIL.n4 VSUBS 0.015929f
C639 VTAIL.n5 VSUBS 0.037649f
C640 VTAIL.n6 VSUBS 0.016865f
C641 VTAIL.n7 VSUBS 0.112316f
C642 VTAIL.t10 VSUBS 0.08205f
C643 VTAIL.n8 VSUBS 0.028237f
C644 VTAIL.n9 VSUBS 0.023681f
C645 VTAIL.n10 VSUBS 0.015929f
C646 VTAIL.n11 VSUBS 0.380834f
C647 VTAIL.n12 VSUBS 0.029642f
C648 VTAIL.n13 VSUBS 0.015929f
C649 VTAIL.n14 VSUBS 0.016865f
C650 VTAIL.n15 VSUBS 0.037649f
C651 VTAIL.n16 VSUBS 0.083446f
C652 VTAIL.n17 VSUBS 0.016865f
C653 VTAIL.n18 VSUBS 0.015929f
C654 VTAIL.n19 VSUBS 0.066492f
C655 VTAIL.n20 VSUBS 0.04156f
C656 VTAIL.n21 VSUBS 0.401291f
C657 VTAIL.t7 VSUBS 0.088778f
C658 VTAIL.t8 VSUBS 0.088778f
C659 VTAIL.n22 VSUBS 0.438989f
C660 VTAIL.n23 VSUBS 1.82009f
C661 VTAIL.t0 VSUBS 0.088778f
C662 VTAIL.t5 VSUBS 0.088778f
C663 VTAIL.n24 VSUBS 0.438993f
C664 VTAIL.n25 VSUBS 1.82009f
C665 VTAIL.n26 VSUBS 0.03031f
C666 VTAIL.n27 VSUBS 0.029642f
C667 VTAIL.n28 VSUBS 0.015929f
C668 VTAIL.n29 VSUBS 0.037649f
C669 VTAIL.n30 VSUBS 0.016865f
C670 VTAIL.n31 VSUBS 0.112316f
C671 VTAIL.t4 VSUBS 0.08205f
C672 VTAIL.n32 VSUBS 0.028237f
C673 VTAIL.n33 VSUBS 0.023681f
C674 VTAIL.n34 VSUBS 0.015929f
C675 VTAIL.n35 VSUBS 0.380834f
C676 VTAIL.n36 VSUBS 0.029642f
C677 VTAIL.n37 VSUBS 0.015929f
C678 VTAIL.n38 VSUBS 0.016865f
C679 VTAIL.n39 VSUBS 0.037649f
C680 VTAIL.n40 VSUBS 0.083446f
C681 VTAIL.n41 VSUBS 0.016865f
C682 VTAIL.n42 VSUBS 0.015929f
C683 VTAIL.n43 VSUBS 0.066492f
C684 VTAIL.n44 VSUBS 0.04156f
C685 VTAIL.n45 VSUBS 0.401291f
C686 VTAIL.t6 VSUBS 0.088778f
C687 VTAIL.t11 VSUBS 0.088778f
C688 VTAIL.n46 VSUBS 0.438993f
C689 VTAIL.n47 VSUBS 0.817997f
C690 VTAIL.n48 VSUBS 0.03031f
C691 VTAIL.n49 VSUBS 0.029642f
C692 VTAIL.n50 VSUBS 0.015929f
C693 VTAIL.n51 VSUBS 0.037649f
C694 VTAIL.n52 VSUBS 0.016865f
C695 VTAIL.n53 VSUBS 0.112316f
C696 VTAIL.t9 VSUBS 0.08205f
C697 VTAIL.n54 VSUBS 0.028237f
C698 VTAIL.n55 VSUBS 0.023681f
C699 VTAIL.n56 VSUBS 0.015929f
C700 VTAIL.n57 VSUBS 0.380834f
C701 VTAIL.n58 VSUBS 0.029642f
C702 VTAIL.n59 VSUBS 0.015929f
C703 VTAIL.n60 VSUBS 0.016865f
C704 VTAIL.n61 VSUBS 0.037649f
C705 VTAIL.n62 VSUBS 0.083446f
C706 VTAIL.n63 VSUBS 0.016865f
C707 VTAIL.n64 VSUBS 0.015929f
C708 VTAIL.n65 VSUBS 0.066492f
C709 VTAIL.n66 VSUBS 0.04156f
C710 VTAIL.n67 VSUBS 1.18189f
C711 VTAIL.n68 VSUBS 0.03031f
C712 VTAIL.n69 VSUBS 0.029642f
C713 VTAIL.n70 VSUBS 0.015929f
C714 VTAIL.n71 VSUBS 0.037649f
C715 VTAIL.n72 VSUBS 0.016865f
C716 VTAIL.n73 VSUBS 0.112316f
C717 VTAIL.t1 VSUBS 0.08205f
C718 VTAIL.n74 VSUBS 0.028237f
C719 VTAIL.n75 VSUBS 0.023681f
C720 VTAIL.n76 VSUBS 0.015929f
C721 VTAIL.n77 VSUBS 0.380834f
C722 VTAIL.n78 VSUBS 0.029642f
C723 VTAIL.n79 VSUBS 0.015929f
C724 VTAIL.n80 VSUBS 0.016865f
C725 VTAIL.n81 VSUBS 0.037649f
C726 VTAIL.n82 VSUBS 0.083446f
C727 VTAIL.n83 VSUBS 0.016865f
C728 VTAIL.n84 VSUBS 0.015929f
C729 VTAIL.n85 VSUBS 0.066492f
C730 VTAIL.n86 VSUBS 0.04156f
C731 VTAIL.n87 VSUBS 1.12096f
C732 VDD1.n0 VSUBS 0.023042f
C733 VDD1.n1 VSUBS 0.022534f
C734 VDD1.n2 VSUBS 0.012109f
C735 VDD1.n3 VSUBS 0.028621f
C736 VDD1.n4 VSUBS 0.012821f
C737 VDD1.n5 VSUBS 0.085382f
C738 VDD1.t0 VSUBS 0.062374f
C739 VDD1.n6 VSUBS 0.021466f
C740 VDD1.n7 VSUBS 0.018002f
C741 VDD1.n8 VSUBS 0.012109f
C742 VDD1.n9 VSUBS 0.28951f
C743 VDD1.n10 VSUBS 0.022534f
C744 VDD1.n11 VSUBS 0.012109f
C745 VDD1.n12 VSUBS 0.012821f
C746 VDD1.n13 VSUBS 0.028621f
C747 VDD1.n14 VSUBS 0.063436f
C748 VDD1.n15 VSUBS 0.012821f
C749 VDD1.n16 VSUBS 0.012109f
C750 VDD1.n17 VSUBS 0.050547f
C751 VDD1.n18 VSUBS 0.053424f
C752 VDD1.n19 VSUBS 0.023042f
C753 VDD1.n20 VSUBS 0.022534f
C754 VDD1.n21 VSUBS 0.012109f
C755 VDD1.n22 VSUBS 0.028621f
C756 VDD1.n23 VSUBS 0.012821f
C757 VDD1.n24 VSUBS 0.085382f
C758 VDD1.t1 VSUBS 0.062374f
C759 VDD1.n25 VSUBS 0.021466f
C760 VDD1.n26 VSUBS 0.018002f
C761 VDD1.n27 VSUBS 0.012109f
C762 VDD1.n28 VSUBS 0.28951f
C763 VDD1.n29 VSUBS 0.022534f
C764 VDD1.n30 VSUBS 0.012109f
C765 VDD1.n31 VSUBS 0.012821f
C766 VDD1.n32 VSUBS 0.028621f
C767 VDD1.n33 VSUBS 0.063436f
C768 VDD1.n34 VSUBS 0.012821f
C769 VDD1.n35 VSUBS 0.012109f
C770 VDD1.n36 VSUBS 0.050547f
C771 VDD1.n37 VSUBS 0.052772f
C772 VDD1.t2 VSUBS 0.067489f
C773 VDD1.t5 VSUBS 0.067489f
C774 VDD1.n38 VSUBS 0.389718f
C775 VDD1.n39 VSUBS 2.10275f
C776 VDD1.t4 VSUBS 0.067489f
C777 VDD1.t3 VSUBS 0.067489f
C778 VDD1.n40 VSUBS 0.387267f
C779 VDD1.n41 VSUBS 2.00304f
C780 VP.n0 VSUBS 0.063469f
C781 VP.t1 VSUBS 1.10058f
C782 VP.n1 VSUBS 0.056157f
C783 VP.n2 VSUBS 0.048141f
C784 VP.t3 VSUBS 1.10058f
C785 VP.n3 VSUBS 0.089722f
C786 VP.n4 VSUBS 0.048141f
C787 VP.n5 VSUBS 0.062258f
C788 VP.n6 VSUBS 0.063469f
C789 VP.t2 VSUBS 1.10058f
C790 VP.n7 VSUBS 0.056157f
C791 VP.n8 VSUBS 0.453567f
C792 VP.t0 VSUBS 1.10058f
C793 VP.t5 VSUBS 1.43661f
C794 VP.n9 VSUBS 0.551669f
C795 VP.n10 VSUBS 0.603759f
C796 VP.n11 VSUBS 0.089722f
C797 VP.n12 VSUBS 0.082782f
C798 VP.n13 VSUBS 0.048141f
C799 VP.n14 VSUBS 0.048141f
C800 VP.n15 VSUBS 0.048141f
C801 VP.n16 VSUBS 0.091346f
C802 VP.n17 VSUBS 0.062258f
C803 VP.n18 VSUBS 0.590484f
C804 VP.n19 VSUBS 2.00173f
C805 VP.t4 VSUBS 1.10058f
C806 VP.n20 VSUBS 0.590484f
C807 VP.n21 VSUBS 2.04346f
C808 VP.n22 VSUBS 0.063469f
C809 VP.n23 VSUBS 0.048141f
C810 VP.n24 VSUBS 0.091346f
C811 VP.n25 VSUBS 0.056157f
C812 VP.n26 VSUBS 0.082782f
C813 VP.n27 VSUBS 0.048141f
C814 VP.n28 VSUBS 0.048141f
C815 VP.n29 VSUBS 0.048141f
C816 VP.n30 VSUBS 0.49196f
C817 VP.n31 VSUBS 0.089722f
C818 VP.n32 VSUBS 0.082782f
C819 VP.n33 VSUBS 0.048141f
C820 VP.n34 VSUBS 0.048141f
C821 VP.n35 VSUBS 0.048141f
C822 VP.n36 VSUBS 0.091346f
C823 VP.n37 VSUBS 0.062258f
C824 VP.n38 VSUBS 0.590484f
C825 VP.n39 VSUBS 0.075479f
.ends

