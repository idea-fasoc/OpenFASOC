* NGSPICE file created from diff_pair_sample_0172.ext - technology: sky130A

.subckt diff_pair_sample_0172 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=0.7491 pd=4.87 as=1.7706 ps=9.86 w=4.54 l=2.84
X1 VDD1.t2 VP.t1 VTAIL.t6 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=0.7491 pd=4.87 as=1.7706 ps=9.86 w=4.54 l=2.84
X2 B.t11 B.t9 B.t10 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0 ps=0 w=4.54 l=2.84
X3 VTAIL.t2 VN.t0 VDD2.t3 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0.7491 ps=4.87 w=4.54 l=2.84
X4 VDD2.t2 VN.t1 VTAIL.t3 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=0.7491 pd=4.87 as=1.7706 ps=9.86 w=4.54 l=2.84
X5 B.t8 B.t6 B.t7 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0 ps=0 w=4.54 l=2.84
X6 VTAIL.t4 VP.t2 VDD1.t1 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0.7491 ps=4.87 w=4.54 l=2.84
X7 VTAIL.t0 VN.t2 VDD2.t1 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0.7491 ps=4.87 w=4.54 l=2.84
X8 B.t5 B.t3 B.t4 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0 ps=0 w=4.54 l=2.84
X9 VDD2.t0 VN.t3 VTAIL.t1 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=0.7491 pd=4.87 as=1.7706 ps=9.86 w=4.54 l=2.84
X10 B.t2 B.t0 B.t1 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0 ps=0 w=4.54 l=2.84
X11 VTAIL.t5 VP.t3 VDD1.t0 w_n2872_n1876# sky130_fd_pr__pfet_01v8 ad=1.7706 pd=9.86 as=0.7491 ps=4.87 w=4.54 l=2.84
R0 VP.n16 VP.n0 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n13 VP.n1 161.3
R3 VP.n12 VP.n11 161.3
R4 VP.n10 VP.n2 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n3 161.3
R7 VP.n6 VP.n5 106.728
R8 VP.n18 VP.n17 106.728
R9 VP.n4 VP.t3 73.9162
R10 VP.n4 VP.t0 73.0193
R11 VP.n6 VP.n4 44.8383
R12 VP.n11 VP.n10 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n5 VP.t2 38.5266
R15 VP.n17 VP.t1 38.5266
R16 VP.n9 VP.n3 24.5923
R17 VP.n10 VP.n9 24.5923
R18 VP.n15 VP.n1 24.5923
R19 VP.n16 VP.n15 24.5923
R20 VP.n5 VP.n3 4.18111
R21 VP.n17 VP.n16 4.18111
R22 VP.n7 VP.n6 0.278335
R23 VP.n18 VP.n0 0.278335
R24 VP.n8 VP.n7 0.189894
R25 VP.n8 VP.n2 0.189894
R26 VP.n12 VP.n2 0.189894
R27 VP.n13 VP.n12 0.189894
R28 VP.n14 VP.n13 0.189894
R29 VP.n14 VP.n0 0.189894
R30 VP VP.n18 0.153485
R31 VTAIL.n186 VTAIL.n168 756.745
R32 VTAIL.n18 VTAIL.n0 756.745
R33 VTAIL.n42 VTAIL.n24 756.745
R34 VTAIL.n66 VTAIL.n48 756.745
R35 VTAIL.n162 VTAIL.n144 756.745
R36 VTAIL.n138 VTAIL.n120 756.745
R37 VTAIL.n114 VTAIL.n96 756.745
R38 VTAIL.n90 VTAIL.n72 756.745
R39 VTAIL.n177 VTAIL.n176 585
R40 VTAIL.n179 VTAIL.n178 585
R41 VTAIL.n172 VTAIL.n171 585
R42 VTAIL.n185 VTAIL.n184 585
R43 VTAIL.n187 VTAIL.n186 585
R44 VTAIL.n9 VTAIL.n8 585
R45 VTAIL.n11 VTAIL.n10 585
R46 VTAIL.n4 VTAIL.n3 585
R47 VTAIL.n17 VTAIL.n16 585
R48 VTAIL.n19 VTAIL.n18 585
R49 VTAIL.n33 VTAIL.n32 585
R50 VTAIL.n35 VTAIL.n34 585
R51 VTAIL.n28 VTAIL.n27 585
R52 VTAIL.n41 VTAIL.n40 585
R53 VTAIL.n43 VTAIL.n42 585
R54 VTAIL.n57 VTAIL.n56 585
R55 VTAIL.n59 VTAIL.n58 585
R56 VTAIL.n52 VTAIL.n51 585
R57 VTAIL.n65 VTAIL.n64 585
R58 VTAIL.n67 VTAIL.n66 585
R59 VTAIL.n163 VTAIL.n162 585
R60 VTAIL.n161 VTAIL.n160 585
R61 VTAIL.n148 VTAIL.n147 585
R62 VTAIL.n155 VTAIL.n154 585
R63 VTAIL.n153 VTAIL.n152 585
R64 VTAIL.n139 VTAIL.n138 585
R65 VTAIL.n137 VTAIL.n136 585
R66 VTAIL.n124 VTAIL.n123 585
R67 VTAIL.n131 VTAIL.n130 585
R68 VTAIL.n129 VTAIL.n128 585
R69 VTAIL.n115 VTAIL.n114 585
R70 VTAIL.n113 VTAIL.n112 585
R71 VTAIL.n100 VTAIL.n99 585
R72 VTAIL.n107 VTAIL.n106 585
R73 VTAIL.n105 VTAIL.n104 585
R74 VTAIL.n91 VTAIL.n90 585
R75 VTAIL.n89 VTAIL.n88 585
R76 VTAIL.n76 VTAIL.n75 585
R77 VTAIL.n83 VTAIL.n82 585
R78 VTAIL.n81 VTAIL.n80 585
R79 VTAIL.n175 VTAIL.t1 328.587
R80 VTAIL.n7 VTAIL.t2 328.587
R81 VTAIL.n31 VTAIL.t6 328.587
R82 VTAIL.n55 VTAIL.t4 328.587
R83 VTAIL.n151 VTAIL.t7 328.587
R84 VTAIL.n127 VTAIL.t5 328.587
R85 VTAIL.n103 VTAIL.t3 328.587
R86 VTAIL.n79 VTAIL.t0 328.587
R87 VTAIL.n178 VTAIL.n177 171.744
R88 VTAIL.n178 VTAIL.n171 171.744
R89 VTAIL.n185 VTAIL.n171 171.744
R90 VTAIL.n186 VTAIL.n185 171.744
R91 VTAIL.n10 VTAIL.n9 171.744
R92 VTAIL.n10 VTAIL.n3 171.744
R93 VTAIL.n17 VTAIL.n3 171.744
R94 VTAIL.n18 VTAIL.n17 171.744
R95 VTAIL.n34 VTAIL.n33 171.744
R96 VTAIL.n34 VTAIL.n27 171.744
R97 VTAIL.n41 VTAIL.n27 171.744
R98 VTAIL.n42 VTAIL.n41 171.744
R99 VTAIL.n58 VTAIL.n57 171.744
R100 VTAIL.n58 VTAIL.n51 171.744
R101 VTAIL.n65 VTAIL.n51 171.744
R102 VTAIL.n66 VTAIL.n65 171.744
R103 VTAIL.n162 VTAIL.n161 171.744
R104 VTAIL.n161 VTAIL.n147 171.744
R105 VTAIL.n154 VTAIL.n147 171.744
R106 VTAIL.n154 VTAIL.n153 171.744
R107 VTAIL.n138 VTAIL.n137 171.744
R108 VTAIL.n137 VTAIL.n123 171.744
R109 VTAIL.n130 VTAIL.n123 171.744
R110 VTAIL.n130 VTAIL.n129 171.744
R111 VTAIL.n114 VTAIL.n113 171.744
R112 VTAIL.n113 VTAIL.n99 171.744
R113 VTAIL.n106 VTAIL.n99 171.744
R114 VTAIL.n106 VTAIL.n105 171.744
R115 VTAIL.n90 VTAIL.n89 171.744
R116 VTAIL.n89 VTAIL.n75 171.744
R117 VTAIL.n82 VTAIL.n75 171.744
R118 VTAIL.n82 VTAIL.n81 171.744
R119 VTAIL.n177 VTAIL.t1 85.8723
R120 VTAIL.n9 VTAIL.t2 85.8723
R121 VTAIL.n33 VTAIL.t6 85.8723
R122 VTAIL.n57 VTAIL.t4 85.8723
R123 VTAIL.n153 VTAIL.t7 85.8723
R124 VTAIL.n129 VTAIL.t5 85.8723
R125 VTAIL.n105 VTAIL.t3 85.8723
R126 VTAIL.n81 VTAIL.t0 85.8723
R127 VTAIL.n191 VTAIL.n190 31.7975
R128 VTAIL.n23 VTAIL.n22 31.7975
R129 VTAIL.n47 VTAIL.n46 31.7975
R130 VTAIL.n71 VTAIL.n70 31.7975
R131 VTAIL.n167 VTAIL.n166 31.7975
R132 VTAIL.n143 VTAIL.n142 31.7975
R133 VTAIL.n119 VTAIL.n118 31.7975
R134 VTAIL.n95 VTAIL.n94 31.7975
R135 VTAIL.n191 VTAIL.n167 19.0134
R136 VTAIL.n95 VTAIL.n71 19.0134
R137 VTAIL.n176 VTAIL.n175 16.3651
R138 VTAIL.n8 VTAIL.n7 16.3651
R139 VTAIL.n32 VTAIL.n31 16.3651
R140 VTAIL.n56 VTAIL.n55 16.3651
R141 VTAIL.n152 VTAIL.n151 16.3651
R142 VTAIL.n128 VTAIL.n127 16.3651
R143 VTAIL.n104 VTAIL.n103 16.3651
R144 VTAIL.n80 VTAIL.n79 16.3651
R145 VTAIL.n179 VTAIL.n174 12.8005
R146 VTAIL.n11 VTAIL.n6 12.8005
R147 VTAIL.n35 VTAIL.n30 12.8005
R148 VTAIL.n59 VTAIL.n54 12.8005
R149 VTAIL.n155 VTAIL.n150 12.8005
R150 VTAIL.n131 VTAIL.n126 12.8005
R151 VTAIL.n107 VTAIL.n102 12.8005
R152 VTAIL.n83 VTAIL.n78 12.8005
R153 VTAIL.n180 VTAIL.n172 12.0247
R154 VTAIL.n12 VTAIL.n4 12.0247
R155 VTAIL.n36 VTAIL.n28 12.0247
R156 VTAIL.n60 VTAIL.n52 12.0247
R157 VTAIL.n156 VTAIL.n148 12.0247
R158 VTAIL.n132 VTAIL.n124 12.0247
R159 VTAIL.n108 VTAIL.n100 12.0247
R160 VTAIL.n84 VTAIL.n76 12.0247
R161 VTAIL.n184 VTAIL.n183 11.249
R162 VTAIL.n16 VTAIL.n15 11.249
R163 VTAIL.n40 VTAIL.n39 11.249
R164 VTAIL.n64 VTAIL.n63 11.249
R165 VTAIL.n160 VTAIL.n159 11.249
R166 VTAIL.n136 VTAIL.n135 11.249
R167 VTAIL.n112 VTAIL.n111 11.249
R168 VTAIL.n88 VTAIL.n87 11.249
R169 VTAIL.n187 VTAIL.n170 10.4732
R170 VTAIL.n19 VTAIL.n2 10.4732
R171 VTAIL.n43 VTAIL.n26 10.4732
R172 VTAIL.n67 VTAIL.n50 10.4732
R173 VTAIL.n163 VTAIL.n146 10.4732
R174 VTAIL.n139 VTAIL.n122 10.4732
R175 VTAIL.n115 VTAIL.n98 10.4732
R176 VTAIL.n91 VTAIL.n74 10.4732
R177 VTAIL.n188 VTAIL.n168 9.69747
R178 VTAIL.n20 VTAIL.n0 9.69747
R179 VTAIL.n44 VTAIL.n24 9.69747
R180 VTAIL.n68 VTAIL.n48 9.69747
R181 VTAIL.n164 VTAIL.n144 9.69747
R182 VTAIL.n140 VTAIL.n120 9.69747
R183 VTAIL.n116 VTAIL.n96 9.69747
R184 VTAIL.n92 VTAIL.n72 9.69747
R185 VTAIL.n190 VTAIL.n189 9.45567
R186 VTAIL.n22 VTAIL.n21 9.45567
R187 VTAIL.n46 VTAIL.n45 9.45567
R188 VTAIL.n70 VTAIL.n69 9.45567
R189 VTAIL.n166 VTAIL.n165 9.45567
R190 VTAIL.n142 VTAIL.n141 9.45567
R191 VTAIL.n118 VTAIL.n117 9.45567
R192 VTAIL.n94 VTAIL.n93 9.45567
R193 VTAIL.n189 VTAIL.n188 9.3005
R194 VTAIL.n170 VTAIL.n169 9.3005
R195 VTAIL.n183 VTAIL.n182 9.3005
R196 VTAIL.n181 VTAIL.n180 9.3005
R197 VTAIL.n174 VTAIL.n173 9.3005
R198 VTAIL.n21 VTAIL.n20 9.3005
R199 VTAIL.n2 VTAIL.n1 9.3005
R200 VTAIL.n15 VTAIL.n14 9.3005
R201 VTAIL.n13 VTAIL.n12 9.3005
R202 VTAIL.n6 VTAIL.n5 9.3005
R203 VTAIL.n45 VTAIL.n44 9.3005
R204 VTAIL.n26 VTAIL.n25 9.3005
R205 VTAIL.n39 VTAIL.n38 9.3005
R206 VTAIL.n37 VTAIL.n36 9.3005
R207 VTAIL.n30 VTAIL.n29 9.3005
R208 VTAIL.n69 VTAIL.n68 9.3005
R209 VTAIL.n50 VTAIL.n49 9.3005
R210 VTAIL.n63 VTAIL.n62 9.3005
R211 VTAIL.n61 VTAIL.n60 9.3005
R212 VTAIL.n54 VTAIL.n53 9.3005
R213 VTAIL.n165 VTAIL.n164 9.3005
R214 VTAIL.n146 VTAIL.n145 9.3005
R215 VTAIL.n159 VTAIL.n158 9.3005
R216 VTAIL.n157 VTAIL.n156 9.3005
R217 VTAIL.n150 VTAIL.n149 9.3005
R218 VTAIL.n141 VTAIL.n140 9.3005
R219 VTAIL.n122 VTAIL.n121 9.3005
R220 VTAIL.n135 VTAIL.n134 9.3005
R221 VTAIL.n133 VTAIL.n132 9.3005
R222 VTAIL.n126 VTAIL.n125 9.3005
R223 VTAIL.n117 VTAIL.n116 9.3005
R224 VTAIL.n98 VTAIL.n97 9.3005
R225 VTAIL.n111 VTAIL.n110 9.3005
R226 VTAIL.n109 VTAIL.n108 9.3005
R227 VTAIL.n102 VTAIL.n101 9.3005
R228 VTAIL.n93 VTAIL.n92 9.3005
R229 VTAIL.n74 VTAIL.n73 9.3005
R230 VTAIL.n87 VTAIL.n86 9.3005
R231 VTAIL.n85 VTAIL.n84 9.3005
R232 VTAIL.n78 VTAIL.n77 9.3005
R233 VTAIL.n190 VTAIL.n168 4.26717
R234 VTAIL.n22 VTAIL.n0 4.26717
R235 VTAIL.n46 VTAIL.n24 4.26717
R236 VTAIL.n70 VTAIL.n48 4.26717
R237 VTAIL.n166 VTAIL.n144 4.26717
R238 VTAIL.n142 VTAIL.n120 4.26717
R239 VTAIL.n118 VTAIL.n96 4.26717
R240 VTAIL.n94 VTAIL.n72 4.26717
R241 VTAIL.n175 VTAIL.n173 3.73474
R242 VTAIL.n7 VTAIL.n5 3.73474
R243 VTAIL.n31 VTAIL.n29 3.73474
R244 VTAIL.n55 VTAIL.n53 3.73474
R245 VTAIL.n151 VTAIL.n149 3.73474
R246 VTAIL.n127 VTAIL.n125 3.73474
R247 VTAIL.n103 VTAIL.n101 3.73474
R248 VTAIL.n79 VTAIL.n77 3.73474
R249 VTAIL.n188 VTAIL.n187 3.49141
R250 VTAIL.n20 VTAIL.n19 3.49141
R251 VTAIL.n44 VTAIL.n43 3.49141
R252 VTAIL.n68 VTAIL.n67 3.49141
R253 VTAIL.n164 VTAIL.n163 3.49141
R254 VTAIL.n140 VTAIL.n139 3.49141
R255 VTAIL.n116 VTAIL.n115 3.49141
R256 VTAIL.n92 VTAIL.n91 3.49141
R257 VTAIL.n119 VTAIL.n95 2.73326
R258 VTAIL.n167 VTAIL.n143 2.73326
R259 VTAIL.n71 VTAIL.n47 2.73326
R260 VTAIL.n184 VTAIL.n170 2.71565
R261 VTAIL.n16 VTAIL.n2 2.71565
R262 VTAIL.n40 VTAIL.n26 2.71565
R263 VTAIL.n64 VTAIL.n50 2.71565
R264 VTAIL.n160 VTAIL.n146 2.71565
R265 VTAIL.n136 VTAIL.n122 2.71565
R266 VTAIL.n112 VTAIL.n98 2.71565
R267 VTAIL.n88 VTAIL.n74 2.71565
R268 VTAIL.n183 VTAIL.n172 1.93989
R269 VTAIL.n15 VTAIL.n4 1.93989
R270 VTAIL.n39 VTAIL.n28 1.93989
R271 VTAIL.n63 VTAIL.n52 1.93989
R272 VTAIL.n159 VTAIL.n148 1.93989
R273 VTAIL.n135 VTAIL.n124 1.93989
R274 VTAIL.n111 VTAIL.n100 1.93989
R275 VTAIL.n87 VTAIL.n76 1.93989
R276 VTAIL VTAIL.n23 1.42507
R277 VTAIL VTAIL.n191 1.30869
R278 VTAIL.n180 VTAIL.n179 1.16414
R279 VTAIL.n12 VTAIL.n11 1.16414
R280 VTAIL.n36 VTAIL.n35 1.16414
R281 VTAIL.n60 VTAIL.n59 1.16414
R282 VTAIL.n156 VTAIL.n155 1.16414
R283 VTAIL.n132 VTAIL.n131 1.16414
R284 VTAIL.n108 VTAIL.n107 1.16414
R285 VTAIL.n84 VTAIL.n83 1.16414
R286 VTAIL.n143 VTAIL.n119 0.470328
R287 VTAIL.n47 VTAIL.n23 0.470328
R288 VTAIL.n176 VTAIL.n174 0.388379
R289 VTAIL.n8 VTAIL.n6 0.388379
R290 VTAIL.n32 VTAIL.n30 0.388379
R291 VTAIL.n56 VTAIL.n54 0.388379
R292 VTAIL.n152 VTAIL.n150 0.388379
R293 VTAIL.n128 VTAIL.n126 0.388379
R294 VTAIL.n104 VTAIL.n102 0.388379
R295 VTAIL.n80 VTAIL.n78 0.388379
R296 VTAIL.n181 VTAIL.n173 0.155672
R297 VTAIL.n182 VTAIL.n181 0.155672
R298 VTAIL.n182 VTAIL.n169 0.155672
R299 VTAIL.n189 VTAIL.n169 0.155672
R300 VTAIL.n13 VTAIL.n5 0.155672
R301 VTAIL.n14 VTAIL.n13 0.155672
R302 VTAIL.n14 VTAIL.n1 0.155672
R303 VTAIL.n21 VTAIL.n1 0.155672
R304 VTAIL.n37 VTAIL.n29 0.155672
R305 VTAIL.n38 VTAIL.n37 0.155672
R306 VTAIL.n38 VTAIL.n25 0.155672
R307 VTAIL.n45 VTAIL.n25 0.155672
R308 VTAIL.n61 VTAIL.n53 0.155672
R309 VTAIL.n62 VTAIL.n61 0.155672
R310 VTAIL.n62 VTAIL.n49 0.155672
R311 VTAIL.n69 VTAIL.n49 0.155672
R312 VTAIL.n165 VTAIL.n145 0.155672
R313 VTAIL.n158 VTAIL.n145 0.155672
R314 VTAIL.n158 VTAIL.n157 0.155672
R315 VTAIL.n157 VTAIL.n149 0.155672
R316 VTAIL.n141 VTAIL.n121 0.155672
R317 VTAIL.n134 VTAIL.n121 0.155672
R318 VTAIL.n134 VTAIL.n133 0.155672
R319 VTAIL.n133 VTAIL.n125 0.155672
R320 VTAIL.n117 VTAIL.n97 0.155672
R321 VTAIL.n110 VTAIL.n97 0.155672
R322 VTAIL.n110 VTAIL.n109 0.155672
R323 VTAIL.n109 VTAIL.n101 0.155672
R324 VTAIL.n93 VTAIL.n73 0.155672
R325 VTAIL.n86 VTAIL.n73 0.155672
R326 VTAIL.n86 VTAIL.n85 0.155672
R327 VTAIL.n85 VTAIL.n77 0.155672
R328 VDD1 VDD1.n1 140.043
R329 VDD1 VDD1.n0 103.749
R330 VDD1.n0 VDD1.t0 7.16019
R331 VDD1.n0 VDD1.t3 7.16019
R332 VDD1.n1 VDD1.t1 7.16019
R333 VDD1.n1 VDD1.t2 7.16019
R334 B.n370 B.n369 585
R335 B.n371 B.n48 585
R336 B.n373 B.n372 585
R337 B.n374 B.n47 585
R338 B.n376 B.n375 585
R339 B.n377 B.n46 585
R340 B.n379 B.n378 585
R341 B.n380 B.n45 585
R342 B.n382 B.n381 585
R343 B.n383 B.n44 585
R344 B.n385 B.n384 585
R345 B.n386 B.n43 585
R346 B.n388 B.n387 585
R347 B.n389 B.n42 585
R348 B.n391 B.n390 585
R349 B.n392 B.n41 585
R350 B.n394 B.n393 585
R351 B.n395 B.n40 585
R352 B.n397 B.n396 585
R353 B.n398 B.n37 585
R354 B.n401 B.n400 585
R355 B.n402 B.n36 585
R356 B.n404 B.n403 585
R357 B.n405 B.n35 585
R358 B.n407 B.n406 585
R359 B.n408 B.n34 585
R360 B.n410 B.n409 585
R361 B.n411 B.n33 585
R362 B.n413 B.n412 585
R363 B.n415 B.n414 585
R364 B.n416 B.n29 585
R365 B.n418 B.n417 585
R366 B.n419 B.n28 585
R367 B.n421 B.n420 585
R368 B.n422 B.n27 585
R369 B.n424 B.n423 585
R370 B.n425 B.n26 585
R371 B.n427 B.n426 585
R372 B.n428 B.n25 585
R373 B.n430 B.n429 585
R374 B.n431 B.n24 585
R375 B.n433 B.n432 585
R376 B.n434 B.n23 585
R377 B.n436 B.n435 585
R378 B.n437 B.n22 585
R379 B.n439 B.n438 585
R380 B.n440 B.n21 585
R381 B.n442 B.n441 585
R382 B.n443 B.n20 585
R383 B.n368 B.n49 585
R384 B.n367 B.n366 585
R385 B.n365 B.n50 585
R386 B.n364 B.n363 585
R387 B.n362 B.n51 585
R388 B.n361 B.n360 585
R389 B.n359 B.n52 585
R390 B.n358 B.n357 585
R391 B.n356 B.n53 585
R392 B.n355 B.n354 585
R393 B.n353 B.n54 585
R394 B.n352 B.n351 585
R395 B.n350 B.n55 585
R396 B.n349 B.n348 585
R397 B.n347 B.n56 585
R398 B.n346 B.n345 585
R399 B.n344 B.n57 585
R400 B.n343 B.n342 585
R401 B.n341 B.n58 585
R402 B.n340 B.n339 585
R403 B.n338 B.n59 585
R404 B.n337 B.n336 585
R405 B.n335 B.n60 585
R406 B.n334 B.n333 585
R407 B.n332 B.n61 585
R408 B.n331 B.n330 585
R409 B.n329 B.n62 585
R410 B.n328 B.n327 585
R411 B.n326 B.n63 585
R412 B.n325 B.n324 585
R413 B.n323 B.n64 585
R414 B.n322 B.n321 585
R415 B.n320 B.n65 585
R416 B.n319 B.n318 585
R417 B.n317 B.n66 585
R418 B.n316 B.n315 585
R419 B.n314 B.n67 585
R420 B.n313 B.n312 585
R421 B.n311 B.n68 585
R422 B.n310 B.n309 585
R423 B.n308 B.n69 585
R424 B.n307 B.n306 585
R425 B.n305 B.n70 585
R426 B.n304 B.n303 585
R427 B.n302 B.n71 585
R428 B.n301 B.n300 585
R429 B.n299 B.n72 585
R430 B.n298 B.n297 585
R431 B.n296 B.n73 585
R432 B.n295 B.n294 585
R433 B.n293 B.n74 585
R434 B.n292 B.n291 585
R435 B.n290 B.n75 585
R436 B.n289 B.n288 585
R437 B.n287 B.n76 585
R438 B.n286 B.n285 585
R439 B.n284 B.n77 585
R440 B.n283 B.n282 585
R441 B.n281 B.n78 585
R442 B.n280 B.n279 585
R443 B.n278 B.n79 585
R444 B.n277 B.n276 585
R445 B.n275 B.n80 585
R446 B.n274 B.n273 585
R447 B.n272 B.n81 585
R448 B.n271 B.n270 585
R449 B.n269 B.n82 585
R450 B.n268 B.n267 585
R451 B.n266 B.n83 585
R452 B.n265 B.n264 585
R453 B.n263 B.n84 585
R454 B.n262 B.n261 585
R455 B.n260 B.n85 585
R456 B.n185 B.n114 585
R457 B.n187 B.n186 585
R458 B.n188 B.n113 585
R459 B.n190 B.n189 585
R460 B.n191 B.n112 585
R461 B.n193 B.n192 585
R462 B.n194 B.n111 585
R463 B.n196 B.n195 585
R464 B.n197 B.n110 585
R465 B.n199 B.n198 585
R466 B.n200 B.n109 585
R467 B.n202 B.n201 585
R468 B.n203 B.n108 585
R469 B.n205 B.n204 585
R470 B.n206 B.n107 585
R471 B.n208 B.n207 585
R472 B.n209 B.n106 585
R473 B.n211 B.n210 585
R474 B.n212 B.n105 585
R475 B.n214 B.n213 585
R476 B.n216 B.n215 585
R477 B.n217 B.n101 585
R478 B.n219 B.n218 585
R479 B.n220 B.n100 585
R480 B.n222 B.n221 585
R481 B.n223 B.n99 585
R482 B.n225 B.n224 585
R483 B.n226 B.n98 585
R484 B.n228 B.n227 585
R485 B.n230 B.n95 585
R486 B.n232 B.n231 585
R487 B.n233 B.n94 585
R488 B.n235 B.n234 585
R489 B.n236 B.n93 585
R490 B.n238 B.n237 585
R491 B.n239 B.n92 585
R492 B.n241 B.n240 585
R493 B.n242 B.n91 585
R494 B.n244 B.n243 585
R495 B.n245 B.n90 585
R496 B.n247 B.n246 585
R497 B.n248 B.n89 585
R498 B.n250 B.n249 585
R499 B.n251 B.n88 585
R500 B.n253 B.n252 585
R501 B.n254 B.n87 585
R502 B.n256 B.n255 585
R503 B.n257 B.n86 585
R504 B.n259 B.n258 585
R505 B.n184 B.n183 585
R506 B.n182 B.n115 585
R507 B.n181 B.n180 585
R508 B.n179 B.n116 585
R509 B.n178 B.n177 585
R510 B.n176 B.n117 585
R511 B.n175 B.n174 585
R512 B.n173 B.n118 585
R513 B.n172 B.n171 585
R514 B.n170 B.n119 585
R515 B.n169 B.n168 585
R516 B.n167 B.n120 585
R517 B.n166 B.n165 585
R518 B.n164 B.n121 585
R519 B.n163 B.n162 585
R520 B.n161 B.n122 585
R521 B.n160 B.n159 585
R522 B.n158 B.n123 585
R523 B.n157 B.n156 585
R524 B.n155 B.n124 585
R525 B.n154 B.n153 585
R526 B.n152 B.n125 585
R527 B.n151 B.n150 585
R528 B.n149 B.n126 585
R529 B.n148 B.n147 585
R530 B.n146 B.n127 585
R531 B.n145 B.n144 585
R532 B.n143 B.n128 585
R533 B.n142 B.n141 585
R534 B.n140 B.n129 585
R535 B.n139 B.n138 585
R536 B.n137 B.n130 585
R537 B.n136 B.n135 585
R538 B.n134 B.n131 585
R539 B.n133 B.n132 585
R540 B.n2 B.n0 585
R541 B.n497 B.n1 585
R542 B.n496 B.n495 585
R543 B.n494 B.n3 585
R544 B.n493 B.n492 585
R545 B.n491 B.n4 585
R546 B.n490 B.n489 585
R547 B.n488 B.n5 585
R548 B.n487 B.n486 585
R549 B.n485 B.n6 585
R550 B.n484 B.n483 585
R551 B.n482 B.n7 585
R552 B.n481 B.n480 585
R553 B.n479 B.n8 585
R554 B.n478 B.n477 585
R555 B.n476 B.n9 585
R556 B.n475 B.n474 585
R557 B.n473 B.n10 585
R558 B.n472 B.n471 585
R559 B.n470 B.n11 585
R560 B.n469 B.n468 585
R561 B.n467 B.n12 585
R562 B.n466 B.n465 585
R563 B.n464 B.n13 585
R564 B.n463 B.n462 585
R565 B.n461 B.n14 585
R566 B.n460 B.n459 585
R567 B.n458 B.n15 585
R568 B.n457 B.n456 585
R569 B.n455 B.n16 585
R570 B.n454 B.n453 585
R571 B.n452 B.n17 585
R572 B.n451 B.n450 585
R573 B.n449 B.n18 585
R574 B.n448 B.n447 585
R575 B.n446 B.n19 585
R576 B.n445 B.n444 585
R577 B.n499 B.n498 585
R578 B.n185 B.n184 506.916
R579 B.n444 B.n443 506.916
R580 B.n258 B.n85 506.916
R581 B.n370 B.n49 506.916
R582 B.n96 B.t11 304.659
R583 B.n38 B.t1 304.659
R584 B.n102 B.t5 304.659
R585 B.n30 B.t7 304.659
R586 B.n96 B.t9 246.909
R587 B.n102 B.t3 246.909
R588 B.n30 B.t6 246.909
R589 B.n38 B.t0 246.909
R590 B.n97 B.t10 243.181
R591 B.n39 B.t2 243.181
R592 B.n103 B.t4 243.18
R593 B.n31 B.t8 243.18
R594 B.n184 B.n115 163.367
R595 B.n180 B.n115 163.367
R596 B.n180 B.n179 163.367
R597 B.n179 B.n178 163.367
R598 B.n178 B.n117 163.367
R599 B.n174 B.n117 163.367
R600 B.n174 B.n173 163.367
R601 B.n173 B.n172 163.367
R602 B.n172 B.n119 163.367
R603 B.n168 B.n119 163.367
R604 B.n168 B.n167 163.367
R605 B.n167 B.n166 163.367
R606 B.n166 B.n121 163.367
R607 B.n162 B.n121 163.367
R608 B.n162 B.n161 163.367
R609 B.n161 B.n160 163.367
R610 B.n160 B.n123 163.367
R611 B.n156 B.n123 163.367
R612 B.n156 B.n155 163.367
R613 B.n155 B.n154 163.367
R614 B.n154 B.n125 163.367
R615 B.n150 B.n125 163.367
R616 B.n150 B.n149 163.367
R617 B.n149 B.n148 163.367
R618 B.n148 B.n127 163.367
R619 B.n144 B.n127 163.367
R620 B.n144 B.n143 163.367
R621 B.n143 B.n142 163.367
R622 B.n142 B.n129 163.367
R623 B.n138 B.n129 163.367
R624 B.n138 B.n137 163.367
R625 B.n137 B.n136 163.367
R626 B.n136 B.n131 163.367
R627 B.n132 B.n131 163.367
R628 B.n132 B.n2 163.367
R629 B.n498 B.n2 163.367
R630 B.n498 B.n497 163.367
R631 B.n497 B.n496 163.367
R632 B.n496 B.n3 163.367
R633 B.n492 B.n3 163.367
R634 B.n492 B.n491 163.367
R635 B.n491 B.n490 163.367
R636 B.n490 B.n5 163.367
R637 B.n486 B.n5 163.367
R638 B.n486 B.n485 163.367
R639 B.n485 B.n484 163.367
R640 B.n484 B.n7 163.367
R641 B.n480 B.n7 163.367
R642 B.n480 B.n479 163.367
R643 B.n479 B.n478 163.367
R644 B.n478 B.n9 163.367
R645 B.n474 B.n9 163.367
R646 B.n474 B.n473 163.367
R647 B.n473 B.n472 163.367
R648 B.n472 B.n11 163.367
R649 B.n468 B.n11 163.367
R650 B.n468 B.n467 163.367
R651 B.n467 B.n466 163.367
R652 B.n466 B.n13 163.367
R653 B.n462 B.n13 163.367
R654 B.n462 B.n461 163.367
R655 B.n461 B.n460 163.367
R656 B.n460 B.n15 163.367
R657 B.n456 B.n15 163.367
R658 B.n456 B.n455 163.367
R659 B.n455 B.n454 163.367
R660 B.n454 B.n17 163.367
R661 B.n450 B.n17 163.367
R662 B.n450 B.n449 163.367
R663 B.n449 B.n448 163.367
R664 B.n448 B.n19 163.367
R665 B.n444 B.n19 163.367
R666 B.n186 B.n185 163.367
R667 B.n186 B.n113 163.367
R668 B.n190 B.n113 163.367
R669 B.n191 B.n190 163.367
R670 B.n192 B.n191 163.367
R671 B.n192 B.n111 163.367
R672 B.n196 B.n111 163.367
R673 B.n197 B.n196 163.367
R674 B.n198 B.n197 163.367
R675 B.n198 B.n109 163.367
R676 B.n202 B.n109 163.367
R677 B.n203 B.n202 163.367
R678 B.n204 B.n203 163.367
R679 B.n204 B.n107 163.367
R680 B.n208 B.n107 163.367
R681 B.n209 B.n208 163.367
R682 B.n210 B.n209 163.367
R683 B.n210 B.n105 163.367
R684 B.n214 B.n105 163.367
R685 B.n215 B.n214 163.367
R686 B.n215 B.n101 163.367
R687 B.n219 B.n101 163.367
R688 B.n220 B.n219 163.367
R689 B.n221 B.n220 163.367
R690 B.n221 B.n99 163.367
R691 B.n225 B.n99 163.367
R692 B.n226 B.n225 163.367
R693 B.n227 B.n226 163.367
R694 B.n227 B.n95 163.367
R695 B.n232 B.n95 163.367
R696 B.n233 B.n232 163.367
R697 B.n234 B.n233 163.367
R698 B.n234 B.n93 163.367
R699 B.n238 B.n93 163.367
R700 B.n239 B.n238 163.367
R701 B.n240 B.n239 163.367
R702 B.n240 B.n91 163.367
R703 B.n244 B.n91 163.367
R704 B.n245 B.n244 163.367
R705 B.n246 B.n245 163.367
R706 B.n246 B.n89 163.367
R707 B.n250 B.n89 163.367
R708 B.n251 B.n250 163.367
R709 B.n252 B.n251 163.367
R710 B.n252 B.n87 163.367
R711 B.n256 B.n87 163.367
R712 B.n257 B.n256 163.367
R713 B.n258 B.n257 163.367
R714 B.n262 B.n85 163.367
R715 B.n263 B.n262 163.367
R716 B.n264 B.n263 163.367
R717 B.n264 B.n83 163.367
R718 B.n268 B.n83 163.367
R719 B.n269 B.n268 163.367
R720 B.n270 B.n269 163.367
R721 B.n270 B.n81 163.367
R722 B.n274 B.n81 163.367
R723 B.n275 B.n274 163.367
R724 B.n276 B.n275 163.367
R725 B.n276 B.n79 163.367
R726 B.n280 B.n79 163.367
R727 B.n281 B.n280 163.367
R728 B.n282 B.n281 163.367
R729 B.n282 B.n77 163.367
R730 B.n286 B.n77 163.367
R731 B.n287 B.n286 163.367
R732 B.n288 B.n287 163.367
R733 B.n288 B.n75 163.367
R734 B.n292 B.n75 163.367
R735 B.n293 B.n292 163.367
R736 B.n294 B.n293 163.367
R737 B.n294 B.n73 163.367
R738 B.n298 B.n73 163.367
R739 B.n299 B.n298 163.367
R740 B.n300 B.n299 163.367
R741 B.n300 B.n71 163.367
R742 B.n304 B.n71 163.367
R743 B.n305 B.n304 163.367
R744 B.n306 B.n305 163.367
R745 B.n306 B.n69 163.367
R746 B.n310 B.n69 163.367
R747 B.n311 B.n310 163.367
R748 B.n312 B.n311 163.367
R749 B.n312 B.n67 163.367
R750 B.n316 B.n67 163.367
R751 B.n317 B.n316 163.367
R752 B.n318 B.n317 163.367
R753 B.n318 B.n65 163.367
R754 B.n322 B.n65 163.367
R755 B.n323 B.n322 163.367
R756 B.n324 B.n323 163.367
R757 B.n324 B.n63 163.367
R758 B.n328 B.n63 163.367
R759 B.n329 B.n328 163.367
R760 B.n330 B.n329 163.367
R761 B.n330 B.n61 163.367
R762 B.n334 B.n61 163.367
R763 B.n335 B.n334 163.367
R764 B.n336 B.n335 163.367
R765 B.n336 B.n59 163.367
R766 B.n340 B.n59 163.367
R767 B.n341 B.n340 163.367
R768 B.n342 B.n341 163.367
R769 B.n342 B.n57 163.367
R770 B.n346 B.n57 163.367
R771 B.n347 B.n346 163.367
R772 B.n348 B.n347 163.367
R773 B.n348 B.n55 163.367
R774 B.n352 B.n55 163.367
R775 B.n353 B.n352 163.367
R776 B.n354 B.n353 163.367
R777 B.n354 B.n53 163.367
R778 B.n358 B.n53 163.367
R779 B.n359 B.n358 163.367
R780 B.n360 B.n359 163.367
R781 B.n360 B.n51 163.367
R782 B.n364 B.n51 163.367
R783 B.n365 B.n364 163.367
R784 B.n366 B.n365 163.367
R785 B.n366 B.n49 163.367
R786 B.n443 B.n442 163.367
R787 B.n442 B.n21 163.367
R788 B.n438 B.n21 163.367
R789 B.n438 B.n437 163.367
R790 B.n437 B.n436 163.367
R791 B.n436 B.n23 163.367
R792 B.n432 B.n23 163.367
R793 B.n432 B.n431 163.367
R794 B.n431 B.n430 163.367
R795 B.n430 B.n25 163.367
R796 B.n426 B.n25 163.367
R797 B.n426 B.n425 163.367
R798 B.n425 B.n424 163.367
R799 B.n424 B.n27 163.367
R800 B.n420 B.n27 163.367
R801 B.n420 B.n419 163.367
R802 B.n419 B.n418 163.367
R803 B.n418 B.n29 163.367
R804 B.n414 B.n29 163.367
R805 B.n414 B.n413 163.367
R806 B.n413 B.n33 163.367
R807 B.n409 B.n33 163.367
R808 B.n409 B.n408 163.367
R809 B.n408 B.n407 163.367
R810 B.n407 B.n35 163.367
R811 B.n403 B.n35 163.367
R812 B.n403 B.n402 163.367
R813 B.n402 B.n401 163.367
R814 B.n401 B.n37 163.367
R815 B.n396 B.n37 163.367
R816 B.n396 B.n395 163.367
R817 B.n395 B.n394 163.367
R818 B.n394 B.n41 163.367
R819 B.n390 B.n41 163.367
R820 B.n390 B.n389 163.367
R821 B.n389 B.n388 163.367
R822 B.n388 B.n43 163.367
R823 B.n384 B.n43 163.367
R824 B.n384 B.n383 163.367
R825 B.n383 B.n382 163.367
R826 B.n382 B.n45 163.367
R827 B.n378 B.n45 163.367
R828 B.n378 B.n377 163.367
R829 B.n377 B.n376 163.367
R830 B.n376 B.n47 163.367
R831 B.n372 B.n47 163.367
R832 B.n372 B.n371 163.367
R833 B.n371 B.n370 163.367
R834 B.n97 B.n96 61.4793
R835 B.n103 B.n102 61.4793
R836 B.n31 B.n30 61.4793
R837 B.n39 B.n38 61.4793
R838 B.n229 B.n97 59.5399
R839 B.n104 B.n103 59.5399
R840 B.n32 B.n31 59.5399
R841 B.n399 B.n39 59.5399
R842 B.n445 B.n20 32.9371
R843 B.n369 B.n368 32.9371
R844 B.n260 B.n259 32.9371
R845 B.n183 B.n114 32.9371
R846 B B.n499 18.0485
R847 B.n441 B.n20 10.6151
R848 B.n441 B.n440 10.6151
R849 B.n440 B.n439 10.6151
R850 B.n439 B.n22 10.6151
R851 B.n435 B.n22 10.6151
R852 B.n435 B.n434 10.6151
R853 B.n434 B.n433 10.6151
R854 B.n433 B.n24 10.6151
R855 B.n429 B.n24 10.6151
R856 B.n429 B.n428 10.6151
R857 B.n428 B.n427 10.6151
R858 B.n427 B.n26 10.6151
R859 B.n423 B.n26 10.6151
R860 B.n423 B.n422 10.6151
R861 B.n422 B.n421 10.6151
R862 B.n421 B.n28 10.6151
R863 B.n417 B.n28 10.6151
R864 B.n417 B.n416 10.6151
R865 B.n416 B.n415 10.6151
R866 B.n412 B.n411 10.6151
R867 B.n411 B.n410 10.6151
R868 B.n410 B.n34 10.6151
R869 B.n406 B.n34 10.6151
R870 B.n406 B.n405 10.6151
R871 B.n405 B.n404 10.6151
R872 B.n404 B.n36 10.6151
R873 B.n400 B.n36 10.6151
R874 B.n398 B.n397 10.6151
R875 B.n397 B.n40 10.6151
R876 B.n393 B.n40 10.6151
R877 B.n393 B.n392 10.6151
R878 B.n392 B.n391 10.6151
R879 B.n391 B.n42 10.6151
R880 B.n387 B.n42 10.6151
R881 B.n387 B.n386 10.6151
R882 B.n386 B.n385 10.6151
R883 B.n385 B.n44 10.6151
R884 B.n381 B.n44 10.6151
R885 B.n381 B.n380 10.6151
R886 B.n380 B.n379 10.6151
R887 B.n379 B.n46 10.6151
R888 B.n375 B.n46 10.6151
R889 B.n375 B.n374 10.6151
R890 B.n374 B.n373 10.6151
R891 B.n373 B.n48 10.6151
R892 B.n369 B.n48 10.6151
R893 B.n261 B.n260 10.6151
R894 B.n261 B.n84 10.6151
R895 B.n265 B.n84 10.6151
R896 B.n266 B.n265 10.6151
R897 B.n267 B.n266 10.6151
R898 B.n267 B.n82 10.6151
R899 B.n271 B.n82 10.6151
R900 B.n272 B.n271 10.6151
R901 B.n273 B.n272 10.6151
R902 B.n273 B.n80 10.6151
R903 B.n277 B.n80 10.6151
R904 B.n278 B.n277 10.6151
R905 B.n279 B.n278 10.6151
R906 B.n279 B.n78 10.6151
R907 B.n283 B.n78 10.6151
R908 B.n284 B.n283 10.6151
R909 B.n285 B.n284 10.6151
R910 B.n285 B.n76 10.6151
R911 B.n289 B.n76 10.6151
R912 B.n290 B.n289 10.6151
R913 B.n291 B.n290 10.6151
R914 B.n291 B.n74 10.6151
R915 B.n295 B.n74 10.6151
R916 B.n296 B.n295 10.6151
R917 B.n297 B.n296 10.6151
R918 B.n297 B.n72 10.6151
R919 B.n301 B.n72 10.6151
R920 B.n302 B.n301 10.6151
R921 B.n303 B.n302 10.6151
R922 B.n303 B.n70 10.6151
R923 B.n307 B.n70 10.6151
R924 B.n308 B.n307 10.6151
R925 B.n309 B.n308 10.6151
R926 B.n309 B.n68 10.6151
R927 B.n313 B.n68 10.6151
R928 B.n314 B.n313 10.6151
R929 B.n315 B.n314 10.6151
R930 B.n315 B.n66 10.6151
R931 B.n319 B.n66 10.6151
R932 B.n320 B.n319 10.6151
R933 B.n321 B.n320 10.6151
R934 B.n321 B.n64 10.6151
R935 B.n325 B.n64 10.6151
R936 B.n326 B.n325 10.6151
R937 B.n327 B.n326 10.6151
R938 B.n327 B.n62 10.6151
R939 B.n331 B.n62 10.6151
R940 B.n332 B.n331 10.6151
R941 B.n333 B.n332 10.6151
R942 B.n333 B.n60 10.6151
R943 B.n337 B.n60 10.6151
R944 B.n338 B.n337 10.6151
R945 B.n339 B.n338 10.6151
R946 B.n339 B.n58 10.6151
R947 B.n343 B.n58 10.6151
R948 B.n344 B.n343 10.6151
R949 B.n345 B.n344 10.6151
R950 B.n345 B.n56 10.6151
R951 B.n349 B.n56 10.6151
R952 B.n350 B.n349 10.6151
R953 B.n351 B.n350 10.6151
R954 B.n351 B.n54 10.6151
R955 B.n355 B.n54 10.6151
R956 B.n356 B.n355 10.6151
R957 B.n357 B.n356 10.6151
R958 B.n357 B.n52 10.6151
R959 B.n361 B.n52 10.6151
R960 B.n362 B.n361 10.6151
R961 B.n363 B.n362 10.6151
R962 B.n363 B.n50 10.6151
R963 B.n367 B.n50 10.6151
R964 B.n368 B.n367 10.6151
R965 B.n187 B.n114 10.6151
R966 B.n188 B.n187 10.6151
R967 B.n189 B.n188 10.6151
R968 B.n189 B.n112 10.6151
R969 B.n193 B.n112 10.6151
R970 B.n194 B.n193 10.6151
R971 B.n195 B.n194 10.6151
R972 B.n195 B.n110 10.6151
R973 B.n199 B.n110 10.6151
R974 B.n200 B.n199 10.6151
R975 B.n201 B.n200 10.6151
R976 B.n201 B.n108 10.6151
R977 B.n205 B.n108 10.6151
R978 B.n206 B.n205 10.6151
R979 B.n207 B.n206 10.6151
R980 B.n207 B.n106 10.6151
R981 B.n211 B.n106 10.6151
R982 B.n212 B.n211 10.6151
R983 B.n213 B.n212 10.6151
R984 B.n217 B.n216 10.6151
R985 B.n218 B.n217 10.6151
R986 B.n218 B.n100 10.6151
R987 B.n222 B.n100 10.6151
R988 B.n223 B.n222 10.6151
R989 B.n224 B.n223 10.6151
R990 B.n224 B.n98 10.6151
R991 B.n228 B.n98 10.6151
R992 B.n231 B.n230 10.6151
R993 B.n231 B.n94 10.6151
R994 B.n235 B.n94 10.6151
R995 B.n236 B.n235 10.6151
R996 B.n237 B.n236 10.6151
R997 B.n237 B.n92 10.6151
R998 B.n241 B.n92 10.6151
R999 B.n242 B.n241 10.6151
R1000 B.n243 B.n242 10.6151
R1001 B.n243 B.n90 10.6151
R1002 B.n247 B.n90 10.6151
R1003 B.n248 B.n247 10.6151
R1004 B.n249 B.n248 10.6151
R1005 B.n249 B.n88 10.6151
R1006 B.n253 B.n88 10.6151
R1007 B.n254 B.n253 10.6151
R1008 B.n255 B.n254 10.6151
R1009 B.n255 B.n86 10.6151
R1010 B.n259 B.n86 10.6151
R1011 B.n183 B.n182 10.6151
R1012 B.n182 B.n181 10.6151
R1013 B.n181 B.n116 10.6151
R1014 B.n177 B.n116 10.6151
R1015 B.n177 B.n176 10.6151
R1016 B.n176 B.n175 10.6151
R1017 B.n175 B.n118 10.6151
R1018 B.n171 B.n118 10.6151
R1019 B.n171 B.n170 10.6151
R1020 B.n170 B.n169 10.6151
R1021 B.n169 B.n120 10.6151
R1022 B.n165 B.n120 10.6151
R1023 B.n165 B.n164 10.6151
R1024 B.n164 B.n163 10.6151
R1025 B.n163 B.n122 10.6151
R1026 B.n159 B.n122 10.6151
R1027 B.n159 B.n158 10.6151
R1028 B.n158 B.n157 10.6151
R1029 B.n157 B.n124 10.6151
R1030 B.n153 B.n124 10.6151
R1031 B.n153 B.n152 10.6151
R1032 B.n152 B.n151 10.6151
R1033 B.n151 B.n126 10.6151
R1034 B.n147 B.n126 10.6151
R1035 B.n147 B.n146 10.6151
R1036 B.n146 B.n145 10.6151
R1037 B.n145 B.n128 10.6151
R1038 B.n141 B.n128 10.6151
R1039 B.n141 B.n140 10.6151
R1040 B.n140 B.n139 10.6151
R1041 B.n139 B.n130 10.6151
R1042 B.n135 B.n130 10.6151
R1043 B.n135 B.n134 10.6151
R1044 B.n134 B.n133 10.6151
R1045 B.n133 B.n0 10.6151
R1046 B.n495 B.n1 10.6151
R1047 B.n495 B.n494 10.6151
R1048 B.n494 B.n493 10.6151
R1049 B.n493 B.n4 10.6151
R1050 B.n489 B.n4 10.6151
R1051 B.n489 B.n488 10.6151
R1052 B.n488 B.n487 10.6151
R1053 B.n487 B.n6 10.6151
R1054 B.n483 B.n6 10.6151
R1055 B.n483 B.n482 10.6151
R1056 B.n482 B.n481 10.6151
R1057 B.n481 B.n8 10.6151
R1058 B.n477 B.n8 10.6151
R1059 B.n477 B.n476 10.6151
R1060 B.n476 B.n475 10.6151
R1061 B.n475 B.n10 10.6151
R1062 B.n471 B.n10 10.6151
R1063 B.n471 B.n470 10.6151
R1064 B.n470 B.n469 10.6151
R1065 B.n469 B.n12 10.6151
R1066 B.n465 B.n12 10.6151
R1067 B.n465 B.n464 10.6151
R1068 B.n464 B.n463 10.6151
R1069 B.n463 B.n14 10.6151
R1070 B.n459 B.n14 10.6151
R1071 B.n459 B.n458 10.6151
R1072 B.n458 B.n457 10.6151
R1073 B.n457 B.n16 10.6151
R1074 B.n453 B.n16 10.6151
R1075 B.n453 B.n452 10.6151
R1076 B.n452 B.n451 10.6151
R1077 B.n451 B.n18 10.6151
R1078 B.n447 B.n18 10.6151
R1079 B.n447 B.n446 10.6151
R1080 B.n446 B.n445 10.6151
R1081 B.n412 B.n32 6.5566
R1082 B.n400 B.n399 6.5566
R1083 B.n216 B.n104 6.5566
R1084 B.n229 B.n228 6.5566
R1085 B.n415 B.n32 4.05904
R1086 B.n399 B.n398 4.05904
R1087 B.n213 B.n104 4.05904
R1088 B.n230 B.n229 4.05904
R1089 B.n499 B.n0 2.81026
R1090 B.n499 B.n1 2.81026
R1091 VN.n0 VN.t0 73.9162
R1092 VN.n1 VN.t1 73.9162
R1093 VN.n0 VN.t3 73.0193
R1094 VN.n1 VN.t2 73.0193
R1095 VN VN.n1 45.1171
R1096 VN VN.n0 3.4391
R1097 VDD2.n2 VDD2.n0 139.518
R1098 VDD2.n2 VDD2.n1 103.692
R1099 VDD2.n1 VDD2.t1 7.16019
R1100 VDD2.n1 VDD2.t2 7.16019
R1101 VDD2.n0 VDD2.t3 7.16019
R1102 VDD2.n0 VDD2.t0 7.16019
R1103 VDD2 VDD2.n2 0.0586897
C0 VTAIL B 2.54045f
C1 B VDD2 1.15873f
C2 VTAIL VN 2.45148f
C3 VP B 1.69283f
C4 w_n2872_n1876# B 7.46527f
C5 VDD2 VN 2.03131f
C6 VP VN 4.98222f
C7 w_n2872_n1876# VN 4.76283f
C8 VTAIL VDD2 3.79222f
C9 VP VTAIL 2.46559f
C10 VDD1 B 1.10246f
C11 w_n2872_n1876# VTAIL 2.30298f
C12 VP VDD2 0.414123f
C13 VDD1 VN 0.153369f
C14 w_n2872_n1876# VDD2 1.35624f
C15 VP w_n2872_n1876# 5.13245f
C16 VDD1 VTAIL 3.7364f
C17 VDD1 VDD2 1.08002f
C18 VDD1 VP 2.29082f
C19 VDD1 w_n2872_n1876# 1.29512f
C20 B VN 1.07812f
C21 VDD2 VSUBS 0.810359f
C22 VDD1 VSUBS 4.911074f
C23 VTAIL VSUBS 0.665056f
C24 VN VSUBS 5.50595f
C25 VP VSUBS 1.952238f
C26 B VSUBS 3.651549f
C27 w_n2872_n1876# VSUBS 67.6528f
C28 VDD2.t3 VSUBS 0.100708f
C29 VDD2.t0 VSUBS 0.100708f
C30 VDD2.n0 VSUBS 0.982741f
C31 VDD2.t1 VSUBS 0.100708f
C32 VDD2.t2 VSUBS 0.100708f
C33 VDD2.n1 VSUBS 0.613472f
C34 VDD2.n2 VSUBS 3.54773f
C35 VN.t0 VSUBS 1.87309f
C36 VN.t3 VSUBS 1.86292f
C37 VN.n0 VSUBS 1.1343f
C38 VN.t1 VSUBS 1.87309f
C39 VN.t2 VSUBS 1.86292f
C40 VN.n1 VSUBS 3.22284f
C41 B.n0 VSUBS 0.005631f
C42 B.n1 VSUBS 0.005631f
C43 B.n2 VSUBS 0.008905f
C44 B.n3 VSUBS 0.008905f
C45 B.n4 VSUBS 0.008905f
C46 B.n5 VSUBS 0.008905f
C47 B.n6 VSUBS 0.008905f
C48 B.n7 VSUBS 0.008905f
C49 B.n8 VSUBS 0.008905f
C50 B.n9 VSUBS 0.008905f
C51 B.n10 VSUBS 0.008905f
C52 B.n11 VSUBS 0.008905f
C53 B.n12 VSUBS 0.008905f
C54 B.n13 VSUBS 0.008905f
C55 B.n14 VSUBS 0.008905f
C56 B.n15 VSUBS 0.008905f
C57 B.n16 VSUBS 0.008905f
C58 B.n17 VSUBS 0.008905f
C59 B.n18 VSUBS 0.008905f
C60 B.n19 VSUBS 0.008905f
C61 B.n20 VSUBS 0.021551f
C62 B.n21 VSUBS 0.008905f
C63 B.n22 VSUBS 0.008905f
C64 B.n23 VSUBS 0.008905f
C65 B.n24 VSUBS 0.008905f
C66 B.n25 VSUBS 0.008905f
C67 B.n26 VSUBS 0.008905f
C68 B.n27 VSUBS 0.008905f
C69 B.n28 VSUBS 0.008905f
C70 B.n29 VSUBS 0.008905f
C71 B.t8 VSUBS 0.083276f
C72 B.t7 VSUBS 0.113745f
C73 B.t6 VSUBS 0.787998f
C74 B.n30 VSUBS 0.196534f
C75 B.n31 VSUBS 0.16369f
C76 B.n32 VSUBS 0.020632f
C77 B.n33 VSUBS 0.008905f
C78 B.n34 VSUBS 0.008905f
C79 B.n35 VSUBS 0.008905f
C80 B.n36 VSUBS 0.008905f
C81 B.n37 VSUBS 0.008905f
C82 B.t2 VSUBS 0.083278f
C83 B.t1 VSUBS 0.113747f
C84 B.t0 VSUBS 0.787998f
C85 B.n38 VSUBS 0.196533f
C86 B.n39 VSUBS 0.163688f
C87 B.n40 VSUBS 0.008905f
C88 B.n41 VSUBS 0.008905f
C89 B.n42 VSUBS 0.008905f
C90 B.n43 VSUBS 0.008905f
C91 B.n44 VSUBS 0.008905f
C92 B.n45 VSUBS 0.008905f
C93 B.n46 VSUBS 0.008905f
C94 B.n47 VSUBS 0.008905f
C95 B.n48 VSUBS 0.008905f
C96 B.n49 VSUBS 0.020355f
C97 B.n50 VSUBS 0.008905f
C98 B.n51 VSUBS 0.008905f
C99 B.n52 VSUBS 0.008905f
C100 B.n53 VSUBS 0.008905f
C101 B.n54 VSUBS 0.008905f
C102 B.n55 VSUBS 0.008905f
C103 B.n56 VSUBS 0.008905f
C104 B.n57 VSUBS 0.008905f
C105 B.n58 VSUBS 0.008905f
C106 B.n59 VSUBS 0.008905f
C107 B.n60 VSUBS 0.008905f
C108 B.n61 VSUBS 0.008905f
C109 B.n62 VSUBS 0.008905f
C110 B.n63 VSUBS 0.008905f
C111 B.n64 VSUBS 0.008905f
C112 B.n65 VSUBS 0.008905f
C113 B.n66 VSUBS 0.008905f
C114 B.n67 VSUBS 0.008905f
C115 B.n68 VSUBS 0.008905f
C116 B.n69 VSUBS 0.008905f
C117 B.n70 VSUBS 0.008905f
C118 B.n71 VSUBS 0.008905f
C119 B.n72 VSUBS 0.008905f
C120 B.n73 VSUBS 0.008905f
C121 B.n74 VSUBS 0.008905f
C122 B.n75 VSUBS 0.008905f
C123 B.n76 VSUBS 0.008905f
C124 B.n77 VSUBS 0.008905f
C125 B.n78 VSUBS 0.008905f
C126 B.n79 VSUBS 0.008905f
C127 B.n80 VSUBS 0.008905f
C128 B.n81 VSUBS 0.008905f
C129 B.n82 VSUBS 0.008905f
C130 B.n83 VSUBS 0.008905f
C131 B.n84 VSUBS 0.008905f
C132 B.n85 VSUBS 0.020355f
C133 B.n86 VSUBS 0.008905f
C134 B.n87 VSUBS 0.008905f
C135 B.n88 VSUBS 0.008905f
C136 B.n89 VSUBS 0.008905f
C137 B.n90 VSUBS 0.008905f
C138 B.n91 VSUBS 0.008905f
C139 B.n92 VSUBS 0.008905f
C140 B.n93 VSUBS 0.008905f
C141 B.n94 VSUBS 0.008905f
C142 B.n95 VSUBS 0.008905f
C143 B.t10 VSUBS 0.083278f
C144 B.t11 VSUBS 0.113747f
C145 B.t9 VSUBS 0.787998f
C146 B.n96 VSUBS 0.196533f
C147 B.n97 VSUBS 0.163688f
C148 B.n98 VSUBS 0.008905f
C149 B.n99 VSUBS 0.008905f
C150 B.n100 VSUBS 0.008905f
C151 B.n101 VSUBS 0.008905f
C152 B.t4 VSUBS 0.083276f
C153 B.t5 VSUBS 0.113745f
C154 B.t3 VSUBS 0.787998f
C155 B.n102 VSUBS 0.196534f
C156 B.n103 VSUBS 0.16369f
C157 B.n104 VSUBS 0.020632f
C158 B.n105 VSUBS 0.008905f
C159 B.n106 VSUBS 0.008905f
C160 B.n107 VSUBS 0.008905f
C161 B.n108 VSUBS 0.008905f
C162 B.n109 VSUBS 0.008905f
C163 B.n110 VSUBS 0.008905f
C164 B.n111 VSUBS 0.008905f
C165 B.n112 VSUBS 0.008905f
C166 B.n113 VSUBS 0.008905f
C167 B.n114 VSUBS 0.021551f
C168 B.n115 VSUBS 0.008905f
C169 B.n116 VSUBS 0.008905f
C170 B.n117 VSUBS 0.008905f
C171 B.n118 VSUBS 0.008905f
C172 B.n119 VSUBS 0.008905f
C173 B.n120 VSUBS 0.008905f
C174 B.n121 VSUBS 0.008905f
C175 B.n122 VSUBS 0.008905f
C176 B.n123 VSUBS 0.008905f
C177 B.n124 VSUBS 0.008905f
C178 B.n125 VSUBS 0.008905f
C179 B.n126 VSUBS 0.008905f
C180 B.n127 VSUBS 0.008905f
C181 B.n128 VSUBS 0.008905f
C182 B.n129 VSUBS 0.008905f
C183 B.n130 VSUBS 0.008905f
C184 B.n131 VSUBS 0.008905f
C185 B.n132 VSUBS 0.008905f
C186 B.n133 VSUBS 0.008905f
C187 B.n134 VSUBS 0.008905f
C188 B.n135 VSUBS 0.008905f
C189 B.n136 VSUBS 0.008905f
C190 B.n137 VSUBS 0.008905f
C191 B.n138 VSUBS 0.008905f
C192 B.n139 VSUBS 0.008905f
C193 B.n140 VSUBS 0.008905f
C194 B.n141 VSUBS 0.008905f
C195 B.n142 VSUBS 0.008905f
C196 B.n143 VSUBS 0.008905f
C197 B.n144 VSUBS 0.008905f
C198 B.n145 VSUBS 0.008905f
C199 B.n146 VSUBS 0.008905f
C200 B.n147 VSUBS 0.008905f
C201 B.n148 VSUBS 0.008905f
C202 B.n149 VSUBS 0.008905f
C203 B.n150 VSUBS 0.008905f
C204 B.n151 VSUBS 0.008905f
C205 B.n152 VSUBS 0.008905f
C206 B.n153 VSUBS 0.008905f
C207 B.n154 VSUBS 0.008905f
C208 B.n155 VSUBS 0.008905f
C209 B.n156 VSUBS 0.008905f
C210 B.n157 VSUBS 0.008905f
C211 B.n158 VSUBS 0.008905f
C212 B.n159 VSUBS 0.008905f
C213 B.n160 VSUBS 0.008905f
C214 B.n161 VSUBS 0.008905f
C215 B.n162 VSUBS 0.008905f
C216 B.n163 VSUBS 0.008905f
C217 B.n164 VSUBS 0.008905f
C218 B.n165 VSUBS 0.008905f
C219 B.n166 VSUBS 0.008905f
C220 B.n167 VSUBS 0.008905f
C221 B.n168 VSUBS 0.008905f
C222 B.n169 VSUBS 0.008905f
C223 B.n170 VSUBS 0.008905f
C224 B.n171 VSUBS 0.008905f
C225 B.n172 VSUBS 0.008905f
C226 B.n173 VSUBS 0.008905f
C227 B.n174 VSUBS 0.008905f
C228 B.n175 VSUBS 0.008905f
C229 B.n176 VSUBS 0.008905f
C230 B.n177 VSUBS 0.008905f
C231 B.n178 VSUBS 0.008905f
C232 B.n179 VSUBS 0.008905f
C233 B.n180 VSUBS 0.008905f
C234 B.n181 VSUBS 0.008905f
C235 B.n182 VSUBS 0.008905f
C236 B.n183 VSUBS 0.020355f
C237 B.n184 VSUBS 0.020355f
C238 B.n185 VSUBS 0.021551f
C239 B.n186 VSUBS 0.008905f
C240 B.n187 VSUBS 0.008905f
C241 B.n188 VSUBS 0.008905f
C242 B.n189 VSUBS 0.008905f
C243 B.n190 VSUBS 0.008905f
C244 B.n191 VSUBS 0.008905f
C245 B.n192 VSUBS 0.008905f
C246 B.n193 VSUBS 0.008905f
C247 B.n194 VSUBS 0.008905f
C248 B.n195 VSUBS 0.008905f
C249 B.n196 VSUBS 0.008905f
C250 B.n197 VSUBS 0.008905f
C251 B.n198 VSUBS 0.008905f
C252 B.n199 VSUBS 0.008905f
C253 B.n200 VSUBS 0.008905f
C254 B.n201 VSUBS 0.008905f
C255 B.n202 VSUBS 0.008905f
C256 B.n203 VSUBS 0.008905f
C257 B.n204 VSUBS 0.008905f
C258 B.n205 VSUBS 0.008905f
C259 B.n206 VSUBS 0.008905f
C260 B.n207 VSUBS 0.008905f
C261 B.n208 VSUBS 0.008905f
C262 B.n209 VSUBS 0.008905f
C263 B.n210 VSUBS 0.008905f
C264 B.n211 VSUBS 0.008905f
C265 B.n212 VSUBS 0.008905f
C266 B.n213 VSUBS 0.006155f
C267 B.n214 VSUBS 0.008905f
C268 B.n215 VSUBS 0.008905f
C269 B.n216 VSUBS 0.007202f
C270 B.n217 VSUBS 0.008905f
C271 B.n218 VSUBS 0.008905f
C272 B.n219 VSUBS 0.008905f
C273 B.n220 VSUBS 0.008905f
C274 B.n221 VSUBS 0.008905f
C275 B.n222 VSUBS 0.008905f
C276 B.n223 VSUBS 0.008905f
C277 B.n224 VSUBS 0.008905f
C278 B.n225 VSUBS 0.008905f
C279 B.n226 VSUBS 0.008905f
C280 B.n227 VSUBS 0.008905f
C281 B.n228 VSUBS 0.007202f
C282 B.n229 VSUBS 0.020632f
C283 B.n230 VSUBS 0.006155f
C284 B.n231 VSUBS 0.008905f
C285 B.n232 VSUBS 0.008905f
C286 B.n233 VSUBS 0.008905f
C287 B.n234 VSUBS 0.008905f
C288 B.n235 VSUBS 0.008905f
C289 B.n236 VSUBS 0.008905f
C290 B.n237 VSUBS 0.008905f
C291 B.n238 VSUBS 0.008905f
C292 B.n239 VSUBS 0.008905f
C293 B.n240 VSUBS 0.008905f
C294 B.n241 VSUBS 0.008905f
C295 B.n242 VSUBS 0.008905f
C296 B.n243 VSUBS 0.008905f
C297 B.n244 VSUBS 0.008905f
C298 B.n245 VSUBS 0.008905f
C299 B.n246 VSUBS 0.008905f
C300 B.n247 VSUBS 0.008905f
C301 B.n248 VSUBS 0.008905f
C302 B.n249 VSUBS 0.008905f
C303 B.n250 VSUBS 0.008905f
C304 B.n251 VSUBS 0.008905f
C305 B.n252 VSUBS 0.008905f
C306 B.n253 VSUBS 0.008905f
C307 B.n254 VSUBS 0.008905f
C308 B.n255 VSUBS 0.008905f
C309 B.n256 VSUBS 0.008905f
C310 B.n257 VSUBS 0.008905f
C311 B.n258 VSUBS 0.021551f
C312 B.n259 VSUBS 0.021551f
C313 B.n260 VSUBS 0.020355f
C314 B.n261 VSUBS 0.008905f
C315 B.n262 VSUBS 0.008905f
C316 B.n263 VSUBS 0.008905f
C317 B.n264 VSUBS 0.008905f
C318 B.n265 VSUBS 0.008905f
C319 B.n266 VSUBS 0.008905f
C320 B.n267 VSUBS 0.008905f
C321 B.n268 VSUBS 0.008905f
C322 B.n269 VSUBS 0.008905f
C323 B.n270 VSUBS 0.008905f
C324 B.n271 VSUBS 0.008905f
C325 B.n272 VSUBS 0.008905f
C326 B.n273 VSUBS 0.008905f
C327 B.n274 VSUBS 0.008905f
C328 B.n275 VSUBS 0.008905f
C329 B.n276 VSUBS 0.008905f
C330 B.n277 VSUBS 0.008905f
C331 B.n278 VSUBS 0.008905f
C332 B.n279 VSUBS 0.008905f
C333 B.n280 VSUBS 0.008905f
C334 B.n281 VSUBS 0.008905f
C335 B.n282 VSUBS 0.008905f
C336 B.n283 VSUBS 0.008905f
C337 B.n284 VSUBS 0.008905f
C338 B.n285 VSUBS 0.008905f
C339 B.n286 VSUBS 0.008905f
C340 B.n287 VSUBS 0.008905f
C341 B.n288 VSUBS 0.008905f
C342 B.n289 VSUBS 0.008905f
C343 B.n290 VSUBS 0.008905f
C344 B.n291 VSUBS 0.008905f
C345 B.n292 VSUBS 0.008905f
C346 B.n293 VSUBS 0.008905f
C347 B.n294 VSUBS 0.008905f
C348 B.n295 VSUBS 0.008905f
C349 B.n296 VSUBS 0.008905f
C350 B.n297 VSUBS 0.008905f
C351 B.n298 VSUBS 0.008905f
C352 B.n299 VSUBS 0.008905f
C353 B.n300 VSUBS 0.008905f
C354 B.n301 VSUBS 0.008905f
C355 B.n302 VSUBS 0.008905f
C356 B.n303 VSUBS 0.008905f
C357 B.n304 VSUBS 0.008905f
C358 B.n305 VSUBS 0.008905f
C359 B.n306 VSUBS 0.008905f
C360 B.n307 VSUBS 0.008905f
C361 B.n308 VSUBS 0.008905f
C362 B.n309 VSUBS 0.008905f
C363 B.n310 VSUBS 0.008905f
C364 B.n311 VSUBS 0.008905f
C365 B.n312 VSUBS 0.008905f
C366 B.n313 VSUBS 0.008905f
C367 B.n314 VSUBS 0.008905f
C368 B.n315 VSUBS 0.008905f
C369 B.n316 VSUBS 0.008905f
C370 B.n317 VSUBS 0.008905f
C371 B.n318 VSUBS 0.008905f
C372 B.n319 VSUBS 0.008905f
C373 B.n320 VSUBS 0.008905f
C374 B.n321 VSUBS 0.008905f
C375 B.n322 VSUBS 0.008905f
C376 B.n323 VSUBS 0.008905f
C377 B.n324 VSUBS 0.008905f
C378 B.n325 VSUBS 0.008905f
C379 B.n326 VSUBS 0.008905f
C380 B.n327 VSUBS 0.008905f
C381 B.n328 VSUBS 0.008905f
C382 B.n329 VSUBS 0.008905f
C383 B.n330 VSUBS 0.008905f
C384 B.n331 VSUBS 0.008905f
C385 B.n332 VSUBS 0.008905f
C386 B.n333 VSUBS 0.008905f
C387 B.n334 VSUBS 0.008905f
C388 B.n335 VSUBS 0.008905f
C389 B.n336 VSUBS 0.008905f
C390 B.n337 VSUBS 0.008905f
C391 B.n338 VSUBS 0.008905f
C392 B.n339 VSUBS 0.008905f
C393 B.n340 VSUBS 0.008905f
C394 B.n341 VSUBS 0.008905f
C395 B.n342 VSUBS 0.008905f
C396 B.n343 VSUBS 0.008905f
C397 B.n344 VSUBS 0.008905f
C398 B.n345 VSUBS 0.008905f
C399 B.n346 VSUBS 0.008905f
C400 B.n347 VSUBS 0.008905f
C401 B.n348 VSUBS 0.008905f
C402 B.n349 VSUBS 0.008905f
C403 B.n350 VSUBS 0.008905f
C404 B.n351 VSUBS 0.008905f
C405 B.n352 VSUBS 0.008905f
C406 B.n353 VSUBS 0.008905f
C407 B.n354 VSUBS 0.008905f
C408 B.n355 VSUBS 0.008905f
C409 B.n356 VSUBS 0.008905f
C410 B.n357 VSUBS 0.008905f
C411 B.n358 VSUBS 0.008905f
C412 B.n359 VSUBS 0.008905f
C413 B.n360 VSUBS 0.008905f
C414 B.n361 VSUBS 0.008905f
C415 B.n362 VSUBS 0.008905f
C416 B.n363 VSUBS 0.008905f
C417 B.n364 VSUBS 0.008905f
C418 B.n365 VSUBS 0.008905f
C419 B.n366 VSUBS 0.008905f
C420 B.n367 VSUBS 0.008905f
C421 B.n368 VSUBS 0.021398f
C422 B.n369 VSUBS 0.020507f
C423 B.n370 VSUBS 0.021551f
C424 B.n371 VSUBS 0.008905f
C425 B.n372 VSUBS 0.008905f
C426 B.n373 VSUBS 0.008905f
C427 B.n374 VSUBS 0.008905f
C428 B.n375 VSUBS 0.008905f
C429 B.n376 VSUBS 0.008905f
C430 B.n377 VSUBS 0.008905f
C431 B.n378 VSUBS 0.008905f
C432 B.n379 VSUBS 0.008905f
C433 B.n380 VSUBS 0.008905f
C434 B.n381 VSUBS 0.008905f
C435 B.n382 VSUBS 0.008905f
C436 B.n383 VSUBS 0.008905f
C437 B.n384 VSUBS 0.008905f
C438 B.n385 VSUBS 0.008905f
C439 B.n386 VSUBS 0.008905f
C440 B.n387 VSUBS 0.008905f
C441 B.n388 VSUBS 0.008905f
C442 B.n389 VSUBS 0.008905f
C443 B.n390 VSUBS 0.008905f
C444 B.n391 VSUBS 0.008905f
C445 B.n392 VSUBS 0.008905f
C446 B.n393 VSUBS 0.008905f
C447 B.n394 VSUBS 0.008905f
C448 B.n395 VSUBS 0.008905f
C449 B.n396 VSUBS 0.008905f
C450 B.n397 VSUBS 0.008905f
C451 B.n398 VSUBS 0.006155f
C452 B.n399 VSUBS 0.020632f
C453 B.n400 VSUBS 0.007202f
C454 B.n401 VSUBS 0.008905f
C455 B.n402 VSUBS 0.008905f
C456 B.n403 VSUBS 0.008905f
C457 B.n404 VSUBS 0.008905f
C458 B.n405 VSUBS 0.008905f
C459 B.n406 VSUBS 0.008905f
C460 B.n407 VSUBS 0.008905f
C461 B.n408 VSUBS 0.008905f
C462 B.n409 VSUBS 0.008905f
C463 B.n410 VSUBS 0.008905f
C464 B.n411 VSUBS 0.008905f
C465 B.n412 VSUBS 0.007202f
C466 B.n413 VSUBS 0.008905f
C467 B.n414 VSUBS 0.008905f
C468 B.n415 VSUBS 0.006155f
C469 B.n416 VSUBS 0.008905f
C470 B.n417 VSUBS 0.008905f
C471 B.n418 VSUBS 0.008905f
C472 B.n419 VSUBS 0.008905f
C473 B.n420 VSUBS 0.008905f
C474 B.n421 VSUBS 0.008905f
C475 B.n422 VSUBS 0.008905f
C476 B.n423 VSUBS 0.008905f
C477 B.n424 VSUBS 0.008905f
C478 B.n425 VSUBS 0.008905f
C479 B.n426 VSUBS 0.008905f
C480 B.n427 VSUBS 0.008905f
C481 B.n428 VSUBS 0.008905f
C482 B.n429 VSUBS 0.008905f
C483 B.n430 VSUBS 0.008905f
C484 B.n431 VSUBS 0.008905f
C485 B.n432 VSUBS 0.008905f
C486 B.n433 VSUBS 0.008905f
C487 B.n434 VSUBS 0.008905f
C488 B.n435 VSUBS 0.008905f
C489 B.n436 VSUBS 0.008905f
C490 B.n437 VSUBS 0.008905f
C491 B.n438 VSUBS 0.008905f
C492 B.n439 VSUBS 0.008905f
C493 B.n440 VSUBS 0.008905f
C494 B.n441 VSUBS 0.008905f
C495 B.n442 VSUBS 0.008905f
C496 B.n443 VSUBS 0.021551f
C497 B.n444 VSUBS 0.020355f
C498 B.n445 VSUBS 0.020355f
C499 B.n446 VSUBS 0.008905f
C500 B.n447 VSUBS 0.008905f
C501 B.n448 VSUBS 0.008905f
C502 B.n449 VSUBS 0.008905f
C503 B.n450 VSUBS 0.008905f
C504 B.n451 VSUBS 0.008905f
C505 B.n452 VSUBS 0.008905f
C506 B.n453 VSUBS 0.008905f
C507 B.n454 VSUBS 0.008905f
C508 B.n455 VSUBS 0.008905f
C509 B.n456 VSUBS 0.008905f
C510 B.n457 VSUBS 0.008905f
C511 B.n458 VSUBS 0.008905f
C512 B.n459 VSUBS 0.008905f
C513 B.n460 VSUBS 0.008905f
C514 B.n461 VSUBS 0.008905f
C515 B.n462 VSUBS 0.008905f
C516 B.n463 VSUBS 0.008905f
C517 B.n464 VSUBS 0.008905f
C518 B.n465 VSUBS 0.008905f
C519 B.n466 VSUBS 0.008905f
C520 B.n467 VSUBS 0.008905f
C521 B.n468 VSUBS 0.008905f
C522 B.n469 VSUBS 0.008905f
C523 B.n470 VSUBS 0.008905f
C524 B.n471 VSUBS 0.008905f
C525 B.n472 VSUBS 0.008905f
C526 B.n473 VSUBS 0.008905f
C527 B.n474 VSUBS 0.008905f
C528 B.n475 VSUBS 0.008905f
C529 B.n476 VSUBS 0.008905f
C530 B.n477 VSUBS 0.008905f
C531 B.n478 VSUBS 0.008905f
C532 B.n479 VSUBS 0.008905f
C533 B.n480 VSUBS 0.008905f
C534 B.n481 VSUBS 0.008905f
C535 B.n482 VSUBS 0.008905f
C536 B.n483 VSUBS 0.008905f
C537 B.n484 VSUBS 0.008905f
C538 B.n485 VSUBS 0.008905f
C539 B.n486 VSUBS 0.008905f
C540 B.n487 VSUBS 0.008905f
C541 B.n488 VSUBS 0.008905f
C542 B.n489 VSUBS 0.008905f
C543 B.n490 VSUBS 0.008905f
C544 B.n491 VSUBS 0.008905f
C545 B.n492 VSUBS 0.008905f
C546 B.n493 VSUBS 0.008905f
C547 B.n494 VSUBS 0.008905f
C548 B.n495 VSUBS 0.008905f
C549 B.n496 VSUBS 0.008905f
C550 B.n497 VSUBS 0.008905f
C551 B.n498 VSUBS 0.008905f
C552 B.n499 VSUBS 0.020164f
C553 VDD1.t0 VSUBS 0.102351f
C554 VDD1.t3 VSUBS 0.102351f
C555 VDD1.n0 VSUBS 0.623868f
C556 VDD1.t1 VSUBS 0.102351f
C557 VDD1.t2 VSUBS 0.102351f
C558 VDD1.n1 VSUBS 1.01776f
C559 VTAIL.n0 VSUBS 0.031529f
C560 VTAIL.n1 VSUBS 0.029964f
C561 VTAIL.n2 VSUBS 0.016101f
C562 VTAIL.n3 VSUBS 0.038058f
C563 VTAIL.n4 VSUBS 0.017049f
C564 VTAIL.n5 VSUBS 0.487157f
C565 VTAIL.n6 VSUBS 0.016101f
C566 VTAIL.t2 VSUBS 0.082547f
C567 VTAIL.n7 VSUBS 0.120274f
C568 VTAIL.n8 VSUBS 0.02411f
C569 VTAIL.n9 VSUBS 0.028543f
C570 VTAIL.n10 VSUBS 0.038058f
C571 VTAIL.n11 VSUBS 0.017049f
C572 VTAIL.n12 VSUBS 0.016101f
C573 VTAIL.n13 VSUBS 0.029964f
C574 VTAIL.n14 VSUBS 0.029964f
C575 VTAIL.n15 VSUBS 0.016101f
C576 VTAIL.n16 VSUBS 0.017049f
C577 VTAIL.n17 VSUBS 0.038058f
C578 VTAIL.n18 VSUBS 0.087381f
C579 VTAIL.n19 VSUBS 0.017049f
C580 VTAIL.n20 VSUBS 0.016101f
C581 VTAIL.n21 VSUBS 0.068442f
C582 VTAIL.n22 VSUBS 0.043707f
C583 VTAIL.n23 VSUBS 0.208036f
C584 VTAIL.n24 VSUBS 0.031529f
C585 VTAIL.n25 VSUBS 0.029964f
C586 VTAIL.n26 VSUBS 0.016101f
C587 VTAIL.n27 VSUBS 0.038058f
C588 VTAIL.n28 VSUBS 0.017049f
C589 VTAIL.n29 VSUBS 0.487157f
C590 VTAIL.n30 VSUBS 0.016101f
C591 VTAIL.t6 VSUBS 0.082547f
C592 VTAIL.n31 VSUBS 0.120274f
C593 VTAIL.n32 VSUBS 0.02411f
C594 VTAIL.n33 VSUBS 0.028543f
C595 VTAIL.n34 VSUBS 0.038058f
C596 VTAIL.n35 VSUBS 0.017049f
C597 VTAIL.n36 VSUBS 0.016101f
C598 VTAIL.n37 VSUBS 0.029964f
C599 VTAIL.n38 VSUBS 0.029964f
C600 VTAIL.n39 VSUBS 0.016101f
C601 VTAIL.n40 VSUBS 0.017049f
C602 VTAIL.n41 VSUBS 0.038058f
C603 VTAIL.n42 VSUBS 0.087381f
C604 VTAIL.n43 VSUBS 0.017049f
C605 VTAIL.n44 VSUBS 0.016101f
C606 VTAIL.n45 VSUBS 0.068442f
C607 VTAIL.n46 VSUBS 0.043707f
C608 VTAIL.n47 VSUBS 0.334343f
C609 VTAIL.n48 VSUBS 0.031529f
C610 VTAIL.n49 VSUBS 0.029964f
C611 VTAIL.n50 VSUBS 0.016101f
C612 VTAIL.n51 VSUBS 0.038058f
C613 VTAIL.n52 VSUBS 0.017049f
C614 VTAIL.n53 VSUBS 0.487157f
C615 VTAIL.n54 VSUBS 0.016101f
C616 VTAIL.t4 VSUBS 0.082547f
C617 VTAIL.n55 VSUBS 0.120274f
C618 VTAIL.n56 VSUBS 0.02411f
C619 VTAIL.n57 VSUBS 0.028543f
C620 VTAIL.n58 VSUBS 0.038058f
C621 VTAIL.n59 VSUBS 0.017049f
C622 VTAIL.n60 VSUBS 0.016101f
C623 VTAIL.n61 VSUBS 0.029964f
C624 VTAIL.n62 VSUBS 0.029964f
C625 VTAIL.n63 VSUBS 0.016101f
C626 VTAIL.n64 VSUBS 0.017049f
C627 VTAIL.n65 VSUBS 0.038058f
C628 VTAIL.n66 VSUBS 0.087381f
C629 VTAIL.n67 VSUBS 0.017049f
C630 VTAIL.n68 VSUBS 0.016101f
C631 VTAIL.n69 VSUBS 0.068442f
C632 VTAIL.n70 VSUBS 0.043707f
C633 VTAIL.n71 VSUBS 1.33774f
C634 VTAIL.n72 VSUBS 0.031529f
C635 VTAIL.n73 VSUBS 0.029964f
C636 VTAIL.n74 VSUBS 0.016101f
C637 VTAIL.n75 VSUBS 0.038058f
C638 VTAIL.n76 VSUBS 0.017049f
C639 VTAIL.n77 VSUBS 0.487157f
C640 VTAIL.n78 VSUBS 0.016101f
C641 VTAIL.t0 VSUBS 0.082547f
C642 VTAIL.n79 VSUBS 0.120274f
C643 VTAIL.n80 VSUBS 0.02411f
C644 VTAIL.n81 VSUBS 0.028543f
C645 VTAIL.n82 VSUBS 0.038058f
C646 VTAIL.n83 VSUBS 0.017049f
C647 VTAIL.n84 VSUBS 0.016101f
C648 VTAIL.n85 VSUBS 0.029964f
C649 VTAIL.n86 VSUBS 0.029964f
C650 VTAIL.n87 VSUBS 0.016101f
C651 VTAIL.n88 VSUBS 0.017049f
C652 VTAIL.n89 VSUBS 0.038058f
C653 VTAIL.n90 VSUBS 0.087381f
C654 VTAIL.n91 VSUBS 0.017049f
C655 VTAIL.n92 VSUBS 0.016101f
C656 VTAIL.n93 VSUBS 0.068442f
C657 VTAIL.n94 VSUBS 0.043707f
C658 VTAIL.n95 VSUBS 1.33774f
C659 VTAIL.n96 VSUBS 0.031529f
C660 VTAIL.n97 VSUBS 0.029964f
C661 VTAIL.n98 VSUBS 0.016101f
C662 VTAIL.n99 VSUBS 0.038058f
C663 VTAIL.n100 VSUBS 0.017049f
C664 VTAIL.n101 VSUBS 0.487157f
C665 VTAIL.n102 VSUBS 0.016101f
C666 VTAIL.t3 VSUBS 0.082547f
C667 VTAIL.n103 VSUBS 0.120274f
C668 VTAIL.n104 VSUBS 0.02411f
C669 VTAIL.n105 VSUBS 0.028543f
C670 VTAIL.n106 VSUBS 0.038058f
C671 VTAIL.n107 VSUBS 0.017049f
C672 VTAIL.n108 VSUBS 0.016101f
C673 VTAIL.n109 VSUBS 0.029964f
C674 VTAIL.n110 VSUBS 0.029964f
C675 VTAIL.n111 VSUBS 0.016101f
C676 VTAIL.n112 VSUBS 0.017049f
C677 VTAIL.n113 VSUBS 0.038058f
C678 VTAIL.n114 VSUBS 0.087381f
C679 VTAIL.n115 VSUBS 0.017049f
C680 VTAIL.n116 VSUBS 0.016101f
C681 VTAIL.n117 VSUBS 0.068442f
C682 VTAIL.n118 VSUBS 0.043707f
C683 VTAIL.n119 VSUBS 0.334343f
C684 VTAIL.n120 VSUBS 0.031529f
C685 VTAIL.n121 VSUBS 0.029964f
C686 VTAIL.n122 VSUBS 0.016101f
C687 VTAIL.n123 VSUBS 0.038058f
C688 VTAIL.n124 VSUBS 0.017049f
C689 VTAIL.n125 VSUBS 0.487157f
C690 VTAIL.n126 VSUBS 0.016101f
C691 VTAIL.t5 VSUBS 0.082547f
C692 VTAIL.n127 VSUBS 0.120274f
C693 VTAIL.n128 VSUBS 0.02411f
C694 VTAIL.n129 VSUBS 0.028543f
C695 VTAIL.n130 VSUBS 0.038058f
C696 VTAIL.n131 VSUBS 0.017049f
C697 VTAIL.n132 VSUBS 0.016101f
C698 VTAIL.n133 VSUBS 0.029964f
C699 VTAIL.n134 VSUBS 0.029964f
C700 VTAIL.n135 VSUBS 0.016101f
C701 VTAIL.n136 VSUBS 0.017049f
C702 VTAIL.n137 VSUBS 0.038058f
C703 VTAIL.n138 VSUBS 0.087381f
C704 VTAIL.n139 VSUBS 0.017049f
C705 VTAIL.n140 VSUBS 0.016101f
C706 VTAIL.n141 VSUBS 0.068442f
C707 VTAIL.n142 VSUBS 0.043707f
C708 VTAIL.n143 VSUBS 0.334343f
C709 VTAIL.n144 VSUBS 0.031529f
C710 VTAIL.n145 VSUBS 0.029964f
C711 VTAIL.n146 VSUBS 0.016101f
C712 VTAIL.n147 VSUBS 0.038058f
C713 VTAIL.n148 VSUBS 0.017049f
C714 VTAIL.n149 VSUBS 0.487157f
C715 VTAIL.n150 VSUBS 0.016101f
C716 VTAIL.t7 VSUBS 0.082547f
C717 VTAIL.n151 VSUBS 0.120274f
C718 VTAIL.n152 VSUBS 0.02411f
C719 VTAIL.n153 VSUBS 0.028543f
C720 VTAIL.n154 VSUBS 0.038058f
C721 VTAIL.n155 VSUBS 0.017049f
C722 VTAIL.n156 VSUBS 0.016101f
C723 VTAIL.n157 VSUBS 0.029964f
C724 VTAIL.n158 VSUBS 0.029964f
C725 VTAIL.n159 VSUBS 0.016101f
C726 VTAIL.n160 VSUBS 0.017049f
C727 VTAIL.n161 VSUBS 0.038058f
C728 VTAIL.n162 VSUBS 0.087381f
C729 VTAIL.n163 VSUBS 0.017049f
C730 VTAIL.n164 VSUBS 0.016101f
C731 VTAIL.n165 VSUBS 0.068442f
C732 VTAIL.n166 VSUBS 0.043707f
C733 VTAIL.n167 VSUBS 1.33774f
C734 VTAIL.n168 VSUBS 0.031529f
C735 VTAIL.n169 VSUBS 0.029964f
C736 VTAIL.n170 VSUBS 0.016101f
C737 VTAIL.n171 VSUBS 0.038058f
C738 VTAIL.n172 VSUBS 0.017049f
C739 VTAIL.n173 VSUBS 0.487157f
C740 VTAIL.n174 VSUBS 0.016101f
C741 VTAIL.t1 VSUBS 0.082547f
C742 VTAIL.n175 VSUBS 0.120274f
C743 VTAIL.n176 VSUBS 0.02411f
C744 VTAIL.n177 VSUBS 0.028543f
C745 VTAIL.n178 VSUBS 0.038058f
C746 VTAIL.n179 VSUBS 0.017049f
C747 VTAIL.n180 VSUBS 0.016101f
C748 VTAIL.n181 VSUBS 0.029964f
C749 VTAIL.n182 VSUBS 0.029964f
C750 VTAIL.n183 VSUBS 0.016101f
C751 VTAIL.n184 VSUBS 0.017049f
C752 VTAIL.n185 VSUBS 0.038058f
C753 VTAIL.n186 VSUBS 0.087381f
C754 VTAIL.n187 VSUBS 0.017049f
C755 VTAIL.n188 VSUBS 0.016101f
C756 VTAIL.n189 VSUBS 0.068442f
C757 VTAIL.n190 VSUBS 0.043707f
C758 VTAIL.n191 VSUBS 1.2002f
C759 VP.n0 VSUBS 0.060079f
C760 VP.t1 VSUBS 1.52581f
C761 VP.n1 VSUBS 0.090098f
C762 VP.n2 VSUBS 0.045573f
C763 VP.n3 VSUBS 0.049882f
C764 VP.t0 VSUBS 1.94943f
C765 VP.t3 VSUBS 1.96007f
C766 VP.n4 VSUBS 3.34801f
C767 VP.t2 VSUBS 1.52581f
C768 VP.n5 VSUBS 0.742408f
C769 VP.n6 VSUBS 2.12857f
C770 VP.n7 VSUBS 0.060079f
C771 VP.n8 VSUBS 0.045573f
C772 VP.n9 VSUBS 0.08451f
C773 VP.n10 VSUBS 0.090098f
C774 VP.n11 VSUBS 0.036807f
C775 VP.n12 VSUBS 0.045573f
C776 VP.n13 VSUBS 0.045573f
C777 VP.n14 VSUBS 0.045573f
C778 VP.n15 VSUBS 0.08451f
C779 VP.n16 VSUBS 0.049882f
C780 VP.n17 VSUBS 0.742408f
C781 VP.n18 VSUBS 0.084381f
.ends

