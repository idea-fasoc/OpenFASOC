* NGSPICE file created from diff_pair_sample_0232.ext - technology: sky130A

.subckt diff_pair_sample_0232 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0 ps=0 w=0.81 l=0.44
X1 VDD2.t5 VN.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0.13365 ps=1.14 w=0.81 l=0.44
X2 VDD1.t5 VP.t0 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0.13365 ps=1.14 w=0.81 l=0.44
X3 VTAIL.t4 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.13365 ps=1.14 w=0.81 l=0.44
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0 ps=0 w=0.81 l=0.44
X5 VDD2.t4 VN.t1 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.3159 ps=2.4 w=0.81 l=0.44
X6 VTAIL.t8 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.13365 ps=1.14 w=0.81 l=0.44
X7 VDD1.t3 VP.t2 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.3159 ps=2.4 w=0.81 l=0.44
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0 ps=0 w=0.81 l=0.44
X9 VDD1.t2 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.3159 ps=2.4 w=0.81 l=0.44
X10 VDD2.t2 VN.t3 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.3159 ps=2.4 w=0.81 l=0.44
X11 VTAIL.t5 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.13365 ps=1.14 w=0.81 l=0.44
X12 VTAIL.t10 VN.t4 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.13365 pd=1.14 as=0.13365 ps=1.14 w=0.81 l=0.44
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0 ps=0 w=0.81 l=0.44
X14 VDD2.t0 VN.t5 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0.13365 ps=1.14 w=0.81 l=0.44
X15 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3159 pd=2.4 as=0.13365 ps=1.14 w=0.81 l=0.44
R0 B.n284 B.n283 585
R1 B.n285 B.n284 585
R2 B.n105 B.n48 585
R3 B.n104 B.n103 585
R4 B.n102 B.n101 585
R5 B.n100 B.n99 585
R6 B.n98 B.n97 585
R7 B.n96 B.n95 585
R8 B.n94 B.n93 585
R9 B.n92 B.n91 585
R10 B.n90 B.n89 585
R11 B.n88 B.n87 585
R12 B.n86 B.n85 585
R13 B.n84 B.n83 585
R14 B.n82 B.n81 585
R15 B.n80 B.n79 585
R16 B.n78 B.n77 585
R17 B.n76 B.n75 585
R18 B.n74 B.n73 585
R19 B.n71 B.n70 585
R20 B.n69 B.n68 585
R21 B.n67 B.n66 585
R22 B.n65 B.n64 585
R23 B.n63 B.n62 585
R24 B.n61 B.n60 585
R25 B.n59 B.n58 585
R26 B.n57 B.n56 585
R27 B.n55 B.n54 585
R28 B.n282 B.n34 585
R29 B.n286 B.n34 585
R30 B.n281 B.n33 585
R31 B.n287 B.n33 585
R32 B.n280 B.n279 585
R33 B.n279 B.n29 585
R34 B.n278 B.n28 585
R35 B.n293 B.n28 585
R36 B.n277 B.n27 585
R37 B.n294 B.n27 585
R38 B.n276 B.n26 585
R39 B.n295 B.n26 585
R40 B.n275 B.n274 585
R41 B.n274 B.n22 585
R42 B.n273 B.n21 585
R43 B.n301 B.n21 585
R44 B.n272 B.n20 585
R45 B.n302 B.n20 585
R46 B.n271 B.n19 585
R47 B.n303 B.n19 585
R48 B.n270 B.n269 585
R49 B.n269 B.n15 585
R50 B.n268 B.n14 585
R51 B.n309 B.n14 585
R52 B.n267 B.n13 585
R53 B.t4 B.n13 585
R54 B.n266 B.n12 585
R55 B.n310 B.n12 585
R56 B.n265 B.n264 585
R57 B.n264 B.n11 585
R58 B.n263 B.n7 585
R59 B.n316 B.n7 585
R60 B.n262 B.n6 585
R61 B.n317 B.n6 585
R62 B.n261 B.n5 585
R63 B.n318 B.n5 585
R64 B.n260 B.n259 585
R65 B.n259 B.n4 585
R66 B.n258 B.n106 585
R67 B.n258 B.n257 585
R68 B.n247 B.n107 585
R69 B.n250 B.n107 585
R70 B.n249 B.n248 585
R71 B.n251 B.n249 585
R72 B.n246 B.n111 585
R73 B.n111 B.t2 585
R74 B.n245 B.n244 585
R75 B.n244 B.n243 585
R76 B.n113 B.n112 585
R77 B.n114 B.n113 585
R78 B.n236 B.n235 585
R79 B.n237 B.n236 585
R80 B.n234 B.n119 585
R81 B.n119 B.n118 585
R82 B.n233 B.n232 585
R83 B.n232 B.n231 585
R84 B.n121 B.n120 585
R85 B.n122 B.n121 585
R86 B.n224 B.n223 585
R87 B.n225 B.n224 585
R88 B.n222 B.n126 585
R89 B.n130 B.n126 585
R90 B.n221 B.n220 585
R91 B.n220 B.n219 585
R92 B.n128 B.n127 585
R93 B.n129 B.n128 585
R94 B.n212 B.n211 585
R95 B.n213 B.n212 585
R96 B.n210 B.n135 585
R97 B.n135 B.n134 585
R98 B.n204 B.n203 585
R99 B.n202 B.n150 585
R100 B.n201 B.n149 585
R101 B.n206 B.n149 585
R102 B.n200 B.n199 585
R103 B.n198 B.n197 585
R104 B.n196 B.n195 585
R105 B.n194 B.n193 585
R106 B.n192 B.n191 585
R107 B.n190 B.n189 585
R108 B.n188 B.n187 585
R109 B.n186 B.n185 585
R110 B.n184 B.n183 585
R111 B.n182 B.n181 585
R112 B.n180 B.n179 585
R113 B.n178 B.n177 585
R114 B.n176 B.n175 585
R115 B.n174 B.n173 585
R116 B.n172 B.n171 585
R117 B.n169 B.n168 585
R118 B.n167 B.n166 585
R119 B.n165 B.n164 585
R120 B.n163 B.n162 585
R121 B.n161 B.n160 585
R122 B.n159 B.n158 585
R123 B.n157 B.n156 585
R124 B.n137 B.n136 585
R125 B.n209 B.n208 585
R126 B.n133 B.n132 585
R127 B.n134 B.n133 585
R128 B.n215 B.n214 585
R129 B.n214 B.n213 585
R130 B.n216 B.n131 585
R131 B.n131 B.n129 585
R132 B.n218 B.n217 585
R133 B.n219 B.n218 585
R134 B.n125 B.n124 585
R135 B.n130 B.n125 585
R136 B.n227 B.n226 585
R137 B.n226 B.n225 585
R138 B.n228 B.n123 585
R139 B.n123 B.n122 585
R140 B.n230 B.n229 585
R141 B.n231 B.n230 585
R142 B.n117 B.n116 585
R143 B.n118 B.n117 585
R144 B.n239 B.n238 585
R145 B.n238 B.n237 585
R146 B.n240 B.n115 585
R147 B.n115 B.n114 585
R148 B.n242 B.n241 585
R149 B.n243 B.n242 585
R150 B.n110 B.n109 585
R151 B.t2 B.n110 585
R152 B.n253 B.n252 585
R153 B.n252 B.n251 585
R154 B.n254 B.n108 585
R155 B.n250 B.n108 585
R156 B.n256 B.n255 585
R157 B.n257 B.n256 585
R158 B.n2 B.n0 585
R159 B.n4 B.n2 585
R160 B.n3 B.n1 585
R161 B.n317 B.n3 585
R162 B.n315 B.n314 585
R163 B.n316 B.n315 585
R164 B.n313 B.n8 585
R165 B.n11 B.n8 585
R166 B.n312 B.n311 585
R167 B.n311 B.n310 585
R168 B.n10 B.n9 585
R169 B.t4 B.n10 585
R170 B.n308 B.n307 585
R171 B.n309 B.n308 585
R172 B.n306 B.n16 585
R173 B.n16 B.n15 585
R174 B.n305 B.n304 585
R175 B.n304 B.n303 585
R176 B.n18 B.n17 585
R177 B.n302 B.n18 585
R178 B.n300 B.n299 585
R179 B.n301 B.n300 585
R180 B.n298 B.n23 585
R181 B.n23 B.n22 585
R182 B.n297 B.n296 585
R183 B.n296 B.n295 585
R184 B.n25 B.n24 585
R185 B.n294 B.n25 585
R186 B.n292 B.n291 585
R187 B.n293 B.n292 585
R188 B.n290 B.n30 585
R189 B.n30 B.n29 585
R190 B.n289 B.n288 585
R191 B.n288 B.n287 585
R192 B.n32 B.n31 585
R193 B.n286 B.n32 585
R194 B.n320 B.n319 585
R195 B.n319 B.n318 585
R196 B.n204 B.n133 526.135
R197 B.n54 B.n32 526.135
R198 B.n208 B.n135 526.135
R199 B.n284 B.n34 526.135
R200 B.n285 B.n47 256.663
R201 B.n285 B.n46 256.663
R202 B.n285 B.n45 256.663
R203 B.n285 B.n44 256.663
R204 B.n285 B.n43 256.663
R205 B.n285 B.n42 256.663
R206 B.n285 B.n41 256.663
R207 B.n285 B.n40 256.663
R208 B.n285 B.n39 256.663
R209 B.n285 B.n38 256.663
R210 B.n285 B.n37 256.663
R211 B.n285 B.n36 256.663
R212 B.n285 B.n35 256.663
R213 B.n206 B.n205 256.663
R214 B.n206 B.n138 256.663
R215 B.n206 B.n139 256.663
R216 B.n206 B.n140 256.663
R217 B.n206 B.n141 256.663
R218 B.n206 B.n142 256.663
R219 B.n206 B.n143 256.663
R220 B.n206 B.n144 256.663
R221 B.n206 B.n145 256.663
R222 B.n206 B.n146 256.663
R223 B.n206 B.n147 256.663
R224 B.n206 B.n148 256.663
R225 B.n207 B.n206 256.663
R226 B.n154 B.t13 252.417
R227 B.n151 B.t17 252.417
R228 B.n52 B.t10 252.417
R229 B.n49 B.t6 252.417
R230 B.n154 B.t16 249.785
R231 B.n151 B.t19 249.785
R232 B.n52 B.t11 249.785
R233 B.n49 B.t8 249.785
R234 B.n206 B.n134 244.043
R235 B.n286 B.n285 244.043
R236 B.n155 B.t15 234.851
R237 B.n152 B.t18 234.851
R238 B.n53 B.t12 234.851
R239 B.n50 B.t9 234.851
R240 B.n214 B.n133 163.367
R241 B.n214 B.n131 163.367
R242 B.n218 B.n131 163.367
R243 B.n218 B.n125 163.367
R244 B.n226 B.n125 163.367
R245 B.n226 B.n123 163.367
R246 B.n230 B.n123 163.367
R247 B.n230 B.n117 163.367
R248 B.n238 B.n117 163.367
R249 B.n238 B.n115 163.367
R250 B.n242 B.n115 163.367
R251 B.n242 B.n110 163.367
R252 B.n252 B.n110 163.367
R253 B.n252 B.n108 163.367
R254 B.n256 B.n108 163.367
R255 B.n256 B.n2 163.367
R256 B.n319 B.n2 163.367
R257 B.n319 B.n3 163.367
R258 B.n315 B.n3 163.367
R259 B.n315 B.n8 163.367
R260 B.n311 B.n8 163.367
R261 B.n311 B.n10 163.367
R262 B.n308 B.n10 163.367
R263 B.n308 B.n16 163.367
R264 B.n304 B.n16 163.367
R265 B.n304 B.n18 163.367
R266 B.n300 B.n18 163.367
R267 B.n300 B.n23 163.367
R268 B.n296 B.n23 163.367
R269 B.n296 B.n25 163.367
R270 B.n292 B.n25 163.367
R271 B.n292 B.n30 163.367
R272 B.n288 B.n30 163.367
R273 B.n288 B.n32 163.367
R274 B.n150 B.n149 163.367
R275 B.n199 B.n149 163.367
R276 B.n197 B.n196 163.367
R277 B.n193 B.n192 163.367
R278 B.n189 B.n188 163.367
R279 B.n185 B.n184 163.367
R280 B.n181 B.n180 163.367
R281 B.n177 B.n176 163.367
R282 B.n173 B.n172 163.367
R283 B.n168 B.n167 163.367
R284 B.n164 B.n163 163.367
R285 B.n160 B.n159 163.367
R286 B.n156 B.n137 163.367
R287 B.n212 B.n135 163.367
R288 B.n212 B.n128 163.367
R289 B.n220 B.n128 163.367
R290 B.n220 B.n126 163.367
R291 B.n224 B.n126 163.367
R292 B.n224 B.n121 163.367
R293 B.n232 B.n121 163.367
R294 B.n232 B.n119 163.367
R295 B.n236 B.n119 163.367
R296 B.n236 B.n113 163.367
R297 B.n244 B.n113 163.367
R298 B.n244 B.n111 163.367
R299 B.n249 B.n111 163.367
R300 B.n249 B.n107 163.367
R301 B.n258 B.n107 163.367
R302 B.n259 B.n258 163.367
R303 B.n259 B.n5 163.367
R304 B.n6 B.n5 163.367
R305 B.n7 B.n6 163.367
R306 B.n264 B.n7 163.367
R307 B.n264 B.n12 163.367
R308 B.n13 B.n12 163.367
R309 B.n14 B.n13 163.367
R310 B.n269 B.n14 163.367
R311 B.n269 B.n19 163.367
R312 B.n20 B.n19 163.367
R313 B.n21 B.n20 163.367
R314 B.n274 B.n21 163.367
R315 B.n274 B.n26 163.367
R316 B.n27 B.n26 163.367
R317 B.n28 B.n27 163.367
R318 B.n279 B.n28 163.367
R319 B.n279 B.n33 163.367
R320 B.n34 B.n33 163.367
R321 B.n58 B.n57 163.367
R322 B.n62 B.n61 163.367
R323 B.n66 B.n65 163.367
R324 B.n70 B.n69 163.367
R325 B.n75 B.n74 163.367
R326 B.n79 B.n78 163.367
R327 B.n83 B.n82 163.367
R328 B.n87 B.n86 163.367
R329 B.n91 B.n90 163.367
R330 B.n95 B.n94 163.367
R331 B.n99 B.n98 163.367
R332 B.n103 B.n102 163.367
R333 B.n284 B.n48 163.367
R334 B.n213 B.n134 122.925
R335 B.n213 B.n129 122.925
R336 B.n219 B.n129 122.925
R337 B.n219 B.n130 122.925
R338 B.n225 B.n122 122.925
R339 B.n231 B.n122 122.925
R340 B.n231 B.n118 122.925
R341 B.n237 B.n118 122.925
R342 B.n243 B.n114 122.925
R343 B.n243 B.t2 122.925
R344 B.n251 B.t2 122.925
R345 B.n251 B.n250 122.925
R346 B.n257 B.n4 122.925
R347 B.n318 B.n4 122.925
R348 B.n318 B.n317 122.925
R349 B.n317 B.n316 122.925
R350 B.n310 B.n11 122.925
R351 B.n310 B.t4 122.925
R352 B.t4 B.n309 122.925
R353 B.n309 B.n15 122.925
R354 B.n303 B.n302 122.925
R355 B.n302 B.n301 122.925
R356 B.n301 B.n22 122.925
R357 B.n295 B.n22 122.925
R358 B.n294 B.n293 122.925
R359 B.n293 B.n29 122.925
R360 B.n287 B.n29 122.925
R361 B.n287 B.n286 122.925
R362 B.n225 B.t14 90.3867
R363 B.n237 B.t1 90.3867
R364 B.n257 B.t5 90.3867
R365 B.n316 B.t3 90.3867
R366 B.n303 B.t0 90.3867
R367 B.n295 B.t7 90.3867
R368 B.n205 B.n204 71.676
R369 B.n199 B.n138 71.676
R370 B.n196 B.n139 71.676
R371 B.n192 B.n140 71.676
R372 B.n188 B.n141 71.676
R373 B.n184 B.n142 71.676
R374 B.n180 B.n143 71.676
R375 B.n176 B.n144 71.676
R376 B.n172 B.n145 71.676
R377 B.n167 B.n146 71.676
R378 B.n163 B.n147 71.676
R379 B.n159 B.n148 71.676
R380 B.n207 B.n137 71.676
R381 B.n54 B.n35 71.676
R382 B.n58 B.n36 71.676
R383 B.n62 B.n37 71.676
R384 B.n66 B.n38 71.676
R385 B.n70 B.n39 71.676
R386 B.n75 B.n40 71.676
R387 B.n79 B.n41 71.676
R388 B.n83 B.n42 71.676
R389 B.n87 B.n43 71.676
R390 B.n91 B.n44 71.676
R391 B.n95 B.n45 71.676
R392 B.n99 B.n46 71.676
R393 B.n103 B.n47 71.676
R394 B.n48 B.n47 71.676
R395 B.n102 B.n46 71.676
R396 B.n98 B.n45 71.676
R397 B.n94 B.n44 71.676
R398 B.n90 B.n43 71.676
R399 B.n86 B.n42 71.676
R400 B.n82 B.n41 71.676
R401 B.n78 B.n40 71.676
R402 B.n74 B.n39 71.676
R403 B.n69 B.n38 71.676
R404 B.n65 B.n37 71.676
R405 B.n61 B.n36 71.676
R406 B.n57 B.n35 71.676
R407 B.n205 B.n150 71.676
R408 B.n197 B.n138 71.676
R409 B.n193 B.n139 71.676
R410 B.n189 B.n140 71.676
R411 B.n185 B.n141 71.676
R412 B.n181 B.n142 71.676
R413 B.n177 B.n143 71.676
R414 B.n173 B.n144 71.676
R415 B.n168 B.n145 71.676
R416 B.n164 B.n146 71.676
R417 B.n160 B.n147 71.676
R418 B.n156 B.n148 71.676
R419 B.n208 B.n207 71.676
R420 B.n170 B.n155 59.5399
R421 B.n153 B.n152 59.5399
R422 B.n72 B.n53 59.5399
R423 B.n51 B.n50 59.5399
R424 B.n55 B.n31 34.1859
R425 B.n283 B.n282 34.1859
R426 B.n210 B.n209 34.1859
R427 B.n203 B.n132 34.1859
R428 B.n130 B.t14 32.5395
R429 B.t1 B.n114 32.5395
R430 B.n250 B.t5 32.5395
R431 B.n11 B.t3 32.5395
R432 B.t0 B.n15 32.5395
R433 B.t7 B.n294 32.5395
R434 B B.n320 18.0485
R435 B.n155 B.n154 14.9338
R436 B.n152 B.n151 14.9338
R437 B.n53 B.n52 14.9338
R438 B.n50 B.n49 14.9338
R439 B.n56 B.n55 10.6151
R440 B.n59 B.n56 10.6151
R441 B.n60 B.n59 10.6151
R442 B.n63 B.n60 10.6151
R443 B.n64 B.n63 10.6151
R444 B.n67 B.n64 10.6151
R445 B.n68 B.n67 10.6151
R446 B.n71 B.n68 10.6151
R447 B.n76 B.n73 10.6151
R448 B.n77 B.n76 10.6151
R449 B.n80 B.n77 10.6151
R450 B.n81 B.n80 10.6151
R451 B.n84 B.n81 10.6151
R452 B.n85 B.n84 10.6151
R453 B.n88 B.n85 10.6151
R454 B.n89 B.n88 10.6151
R455 B.n93 B.n92 10.6151
R456 B.n96 B.n93 10.6151
R457 B.n97 B.n96 10.6151
R458 B.n100 B.n97 10.6151
R459 B.n101 B.n100 10.6151
R460 B.n104 B.n101 10.6151
R461 B.n105 B.n104 10.6151
R462 B.n283 B.n105 10.6151
R463 B.n211 B.n210 10.6151
R464 B.n211 B.n127 10.6151
R465 B.n221 B.n127 10.6151
R466 B.n222 B.n221 10.6151
R467 B.n223 B.n222 10.6151
R468 B.n223 B.n120 10.6151
R469 B.n233 B.n120 10.6151
R470 B.n234 B.n233 10.6151
R471 B.n235 B.n234 10.6151
R472 B.n235 B.n112 10.6151
R473 B.n245 B.n112 10.6151
R474 B.n246 B.n245 10.6151
R475 B.n248 B.n246 10.6151
R476 B.n248 B.n247 10.6151
R477 B.n247 B.n106 10.6151
R478 B.n260 B.n106 10.6151
R479 B.n261 B.n260 10.6151
R480 B.n262 B.n261 10.6151
R481 B.n263 B.n262 10.6151
R482 B.n265 B.n263 10.6151
R483 B.n266 B.n265 10.6151
R484 B.n267 B.n266 10.6151
R485 B.n268 B.n267 10.6151
R486 B.n270 B.n268 10.6151
R487 B.n271 B.n270 10.6151
R488 B.n272 B.n271 10.6151
R489 B.n273 B.n272 10.6151
R490 B.n275 B.n273 10.6151
R491 B.n276 B.n275 10.6151
R492 B.n277 B.n276 10.6151
R493 B.n278 B.n277 10.6151
R494 B.n280 B.n278 10.6151
R495 B.n281 B.n280 10.6151
R496 B.n282 B.n281 10.6151
R497 B.n203 B.n202 10.6151
R498 B.n202 B.n201 10.6151
R499 B.n201 B.n200 10.6151
R500 B.n200 B.n198 10.6151
R501 B.n198 B.n195 10.6151
R502 B.n195 B.n194 10.6151
R503 B.n194 B.n191 10.6151
R504 B.n191 B.n190 10.6151
R505 B.n187 B.n186 10.6151
R506 B.n186 B.n183 10.6151
R507 B.n183 B.n182 10.6151
R508 B.n182 B.n179 10.6151
R509 B.n179 B.n178 10.6151
R510 B.n178 B.n175 10.6151
R511 B.n175 B.n174 10.6151
R512 B.n174 B.n171 10.6151
R513 B.n169 B.n166 10.6151
R514 B.n166 B.n165 10.6151
R515 B.n165 B.n162 10.6151
R516 B.n162 B.n161 10.6151
R517 B.n161 B.n158 10.6151
R518 B.n158 B.n157 10.6151
R519 B.n157 B.n136 10.6151
R520 B.n209 B.n136 10.6151
R521 B.n215 B.n132 10.6151
R522 B.n216 B.n215 10.6151
R523 B.n217 B.n216 10.6151
R524 B.n217 B.n124 10.6151
R525 B.n227 B.n124 10.6151
R526 B.n228 B.n227 10.6151
R527 B.n229 B.n228 10.6151
R528 B.n229 B.n116 10.6151
R529 B.n239 B.n116 10.6151
R530 B.n240 B.n239 10.6151
R531 B.n241 B.n240 10.6151
R532 B.n241 B.n109 10.6151
R533 B.n253 B.n109 10.6151
R534 B.n254 B.n253 10.6151
R535 B.n255 B.n254 10.6151
R536 B.n255 B.n0 10.6151
R537 B.n314 B.n1 10.6151
R538 B.n314 B.n313 10.6151
R539 B.n313 B.n312 10.6151
R540 B.n312 B.n9 10.6151
R541 B.n307 B.n9 10.6151
R542 B.n307 B.n306 10.6151
R543 B.n306 B.n305 10.6151
R544 B.n305 B.n17 10.6151
R545 B.n299 B.n17 10.6151
R546 B.n299 B.n298 10.6151
R547 B.n298 B.n297 10.6151
R548 B.n297 B.n24 10.6151
R549 B.n291 B.n24 10.6151
R550 B.n291 B.n290 10.6151
R551 B.n290 B.n289 10.6151
R552 B.n289 B.n31 10.6151
R553 B.n73 B.n72 6.5566
R554 B.n89 B.n51 6.5566
R555 B.n187 B.n153 6.5566
R556 B.n171 B.n170 6.5566
R557 B.n72 B.n71 4.05904
R558 B.n92 B.n51 4.05904
R559 B.n190 B.n153 4.05904
R560 B.n170 B.n169 4.05904
R561 B.n320 B.n0 2.81026
R562 B.n320 B.n1 2.81026
R563 VN.n3 VN.n2 161.3
R564 VN.n7 VN.n6 161.3
R565 VN.n0 VN.t5 159.656
R566 VN.n4 VN.t3 159.656
R567 VN.n2 VN.t1 141.496
R568 VN.n6 VN.t0 141.496
R569 VN.n1 VN.t2 134.194
R570 VN.n5 VN.t4 134.194
R571 VN.n7 VN.n4 71.8132
R572 VN.n3 VN.n0 71.8132
R573 VN.n2 VN.n1 40.8975
R574 VN.n6 VN.n5 40.8975
R575 VN VN.n7 32.2032
R576 VN.n5 VN.n4 18.1394
R577 VN.n1 VN.n0 18.1394
R578 VN VN.n3 0.0516364
R579 VTAIL.n11 VTAIL.t9 245.702
R580 VTAIL.n2 VTAIL.t3 245.702
R581 VTAIL.n10 VTAIL.t0 245.702
R582 VTAIL.n7 VTAIL.t7 245.702
R583 VTAIL.n1 VTAIL.n0 221.258
R584 VTAIL.n4 VTAIL.n3 221.258
R585 VTAIL.n9 VTAIL.n8 221.258
R586 VTAIL.n6 VTAIL.n5 221.258
R587 VTAIL.n0 VTAIL.t11 24.4449
R588 VTAIL.n0 VTAIL.t8 24.4449
R589 VTAIL.n3 VTAIL.t1 24.4449
R590 VTAIL.n3 VTAIL.t5 24.4449
R591 VTAIL.n8 VTAIL.t2 24.4449
R592 VTAIL.n8 VTAIL.t4 24.4449
R593 VTAIL.n5 VTAIL.t6 24.4449
R594 VTAIL.n5 VTAIL.t10 24.4449
R595 VTAIL.n6 VTAIL.n4 14.3927
R596 VTAIL.n11 VTAIL.n10 13.7289
R597 VTAIL.n9 VTAIL.n7 0.802224
R598 VTAIL.n2 VTAIL.n1 0.802224
R599 VTAIL.n7 VTAIL.n6 0.664293
R600 VTAIL.n10 VTAIL.n9 0.664293
R601 VTAIL.n4 VTAIL.n2 0.664293
R602 VTAIL VTAIL.n11 0.440155
R603 VTAIL VTAIL.n1 0.224638
R604 VDD2.n1 VDD2.t0 262.824
R605 VDD2.n2 VDD2.t5 262.382
R606 VDD2.n1 VDD2.n0 238.048
R607 VDD2 VDD2.n3 238.044
R608 VDD2.n2 VDD2.n1 26.5709
R609 VDD2.n3 VDD2.t1 24.4449
R610 VDD2.n3 VDD2.t2 24.4449
R611 VDD2.n0 VDD2.t3 24.4449
R612 VDD2.n0 VDD2.t4 24.4449
R613 VDD2 VDD2.n2 0.556535
R614 VP.n9 VP.n8 161.3
R615 VP.n4 VP.n3 161.3
R616 VP.n7 VP.n0 161.3
R617 VP.n6 VP.n5 161.3
R618 VP.n1 VP.t0 159.656
R619 VP.n8 VP.t2 141.496
R620 VP.n6 VP.t5 141.496
R621 VP.n3 VP.t3 141.496
R622 VP.n7 VP.t4 134.194
R623 VP.n2 VP.t1 134.194
R624 VP.n4 VP.n1 71.8132
R625 VP.n7 VP.n6 40.8975
R626 VP.n8 VP.n7 40.8975
R627 VP.n3 VP.n2 40.8975
R628 VP.n5 VP.n4 31.8225
R629 VP.n2 VP.n1 18.1394
R630 VP.n5 VP.n0 0.189894
R631 VP.n9 VP.n0 0.189894
R632 VP VP.n9 0.0516364
R633 VDD1 VDD1.t5 262.938
R634 VDD1.n1 VDD1.t0 262.824
R635 VDD1.n1 VDD1.n0 238.048
R636 VDD1.n3 VDD1.n2 237.936
R637 VDD1.n3 VDD1.n1 27.4858
R638 VDD1.n2 VDD1.t4 24.4449
R639 VDD1.n2 VDD1.t2 24.4449
R640 VDD1.n0 VDD1.t1 24.4449
R641 VDD1.n0 VDD1.t3 24.4449
R642 VDD1 VDD1.n3 0.108259
C0 VP VN 2.76277f
C1 VN VDD2 0.528754f
C2 VP VDD1 0.654193f
C3 VDD1 VDD2 0.61472f
C4 VP VDD2 0.28308f
C5 VN VTAIL 0.733115f
C6 VTAIL VDD1 2.37405f
C7 VP VTAIL 0.747261f
C8 VTAIL VDD2 2.41251f
C9 VN VDD1 0.155874f
C10 VDD2 B 2.114578f
C11 VDD1 B 2.262258f
C12 VTAIL B 1.895108f
C13 VN B 5.116458f
C14 VP B 4.030944f
C15 VDD1.t5 B 0.068793f
C16 VDD1.t0 B 0.068732f
C17 VDD1.t1 B 0.014438f
C18 VDD1.t3 B 0.014438f
C19 VDD1.n0 B 0.034796f
C20 VDD1.n1 B 0.952147f
C21 VDD1.t4 B 0.014438f
C22 VDD1.t2 B 0.014438f
C23 VDD1.n2 B 0.034736f
C24 VDD1.n3 B 1.02145f
C25 VP.n0 B 0.038954f
C26 VP.t5 B 0.051787f
C27 VP.t0 B 0.0583f
C28 VP.n1 B 0.050985f
C29 VP.t1 B 0.049155f
C30 VP.n2 B 0.064158f
C31 VP.t3 B 0.051787f
C32 VP.n3 B 0.057203f
C33 VP.n4 B 1.04641f
C34 VP.n5 B 1.00127f
C35 VP.n6 B 0.057203f
C36 VP.t4 B 0.049155f
C37 VP.n7 B 0.064158f
C38 VP.t2 B 0.051787f
C39 VP.n8 B 0.057203f
C40 VP.n9 B 0.030188f
C41 VDD2.t0 B 0.071204f
C42 VDD2.t3 B 0.014957f
C43 VDD2.t4 B 0.014957f
C44 VDD2.n0 B 0.036047f
C45 VDD2.n1 B 0.924386f
C46 VDD2.t5 B 0.071018f
C47 VDD2.n2 B 1.02341f
C48 VDD2.t1 B 0.014957f
C49 VDD2.t2 B 0.014957f
C50 VDD2.n3 B 0.036043f
C51 VTAIL.t11 B 0.022276f
C52 VTAIL.t8 B 0.022276f
C53 VTAIL.n0 B 0.047286f
C54 VTAIL.n1 B 0.164359f
C55 VTAIL.t3 B 0.099507f
C56 VTAIL.n2 B 0.222195f
C57 VTAIL.t1 B 0.022276f
C58 VTAIL.t5 B 0.022276f
C59 VTAIL.n3 B 0.047286f
C60 VTAIL.n4 B 0.823679f
C61 VTAIL.t6 B 0.022276f
C62 VTAIL.t10 B 0.022276f
C63 VTAIL.n5 B 0.047286f
C64 VTAIL.n6 B 0.823679f
C65 VTAIL.t7 B 0.099507f
C66 VTAIL.n7 B 0.222195f
C67 VTAIL.t2 B 0.022276f
C68 VTAIL.t4 B 0.022276f
C69 VTAIL.n8 B 0.047286f
C70 VTAIL.n9 B 0.213662f
C71 VTAIL.t0 B 0.099507f
C72 VTAIL.n10 B 0.757774f
C73 VTAIL.t9 B 0.099507f
C74 VTAIL.n11 B 0.73264f
C75 VN.t5 B 0.057182f
C76 VN.n0 B 0.050007f
C77 VN.t2 B 0.048212f
C78 VN.n1 B 0.062928f
C79 VN.t1 B 0.050793f
C80 VN.n2 B 0.056106f
C81 VN.n3 B 0.11704f
C82 VN.t3 B 0.057182f
C83 VN.n4 B 0.050007f
C84 VN.t0 B 0.050793f
C85 VN.t4 B 0.048212f
C86 VN.n5 B 0.062928f
C87 VN.n6 B 0.056106f
C88 VN.n7 B 1.05193f
.ends

