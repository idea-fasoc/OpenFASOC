* NGSPICE file created from diff_pair_sample_1278.ext - technology: sky130A

.subckt diff_pair_sample_1278 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=1.75395 pd=10.96 as=4.1457 ps=22.04 w=10.63 l=3.96
X1 B.t11 B.t9 B.t10 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=0 ps=0 w=10.63 l=3.96
X2 VDD1.t2 VP.t1 VTAIL.t3 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=1.75395 pd=10.96 as=4.1457 ps=22.04 w=10.63 l=3.96
X3 VTAIL.t1 VN.t0 VDD2.t3 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=1.75395 ps=10.96 w=10.63 l=3.96
X4 VDD2.t2 VN.t1 VTAIL.t7 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=1.75395 pd=10.96 as=4.1457 ps=22.04 w=10.63 l=3.96
X5 B.t8 B.t6 B.t7 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=0 ps=0 w=10.63 l=3.96
X6 VTAIL.t2 VN.t2 VDD2.t1 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=1.75395 ps=10.96 w=10.63 l=3.96
X7 B.t5 B.t3 B.t4 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=0 ps=0 w=10.63 l=3.96
X8 VTAIL.t6 VP.t2 VDD1.t1 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=1.75395 ps=10.96 w=10.63 l=3.96
X9 B.t2 B.t0 B.t1 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=0 ps=0 w=10.63 l=3.96
X10 VTAIL.t5 VP.t3 VDD1.t0 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=4.1457 pd=22.04 as=1.75395 ps=10.96 w=10.63 l=3.96
X11 VDD2.t0 VN.t3 VTAIL.t0 w_n3544_n3094# sky130_fd_pr__pfet_01v8 ad=1.75395 pd=10.96 as=4.1457 ps=22.04 w=10.63 l=3.96
R0 VP.n18 VP.n0 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n15 VP.n1 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n12 VP.n2 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n3 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n4 VP.t2 98.5048
R9 VP.n4 VP.t1 97.0695
R10 VP.n6 VP.t3 64.6932
R11 VP.n19 VP.t0 64.6932
R12 VP.n6 VP.n5 62.8529
R13 VP.n20 VP.n19 62.8529
R14 VP.n13 VP.n12 56.5193
R15 VP.n5 VP.n4 51.3077
R16 VP.n7 VP.n3 24.4675
R17 VP.n11 VP.n3 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n13 VP.n1 24.4675
R20 VP.n17 VP.n1 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n7 VP.n6 19.3294
R23 VP.n19 VP.n18 19.3294
R24 VP.n8 VP.n5 0.417535
R25 VP.n20 VP.n0 0.417535
R26 VP VP.n20 0.394291
R27 VP.n9 VP.n8 0.189894
R28 VP.n10 VP.n9 0.189894
R29 VP.n10 VP.n2 0.189894
R30 VP.n14 VP.n2 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VTAIL.n458 VTAIL.n406 756.745
R35 VTAIL.n52 VTAIL.n0 756.745
R36 VTAIL.n110 VTAIL.n58 756.745
R37 VTAIL.n168 VTAIL.n116 756.745
R38 VTAIL.n400 VTAIL.n348 756.745
R39 VTAIL.n342 VTAIL.n290 756.745
R40 VTAIL.n284 VTAIL.n232 756.745
R41 VTAIL.n226 VTAIL.n174 756.745
R42 VTAIL.n425 VTAIL.n424 585
R43 VTAIL.n422 VTAIL.n421 585
R44 VTAIL.n431 VTAIL.n430 585
R45 VTAIL.n433 VTAIL.n432 585
R46 VTAIL.n418 VTAIL.n417 585
R47 VTAIL.n439 VTAIL.n438 585
R48 VTAIL.n442 VTAIL.n441 585
R49 VTAIL.n440 VTAIL.n414 585
R50 VTAIL.n447 VTAIL.n413 585
R51 VTAIL.n449 VTAIL.n448 585
R52 VTAIL.n451 VTAIL.n450 585
R53 VTAIL.n410 VTAIL.n409 585
R54 VTAIL.n457 VTAIL.n456 585
R55 VTAIL.n459 VTAIL.n458 585
R56 VTAIL.n19 VTAIL.n18 585
R57 VTAIL.n16 VTAIL.n15 585
R58 VTAIL.n25 VTAIL.n24 585
R59 VTAIL.n27 VTAIL.n26 585
R60 VTAIL.n12 VTAIL.n11 585
R61 VTAIL.n33 VTAIL.n32 585
R62 VTAIL.n36 VTAIL.n35 585
R63 VTAIL.n34 VTAIL.n8 585
R64 VTAIL.n41 VTAIL.n7 585
R65 VTAIL.n43 VTAIL.n42 585
R66 VTAIL.n45 VTAIL.n44 585
R67 VTAIL.n4 VTAIL.n3 585
R68 VTAIL.n51 VTAIL.n50 585
R69 VTAIL.n53 VTAIL.n52 585
R70 VTAIL.n77 VTAIL.n76 585
R71 VTAIL.n74 VTAIL.n73 585
R72 VTAIL.n83 VTAIL.n82 585
R73 VTAIL.n85 VTAIL.n84 585
R74 VTAIL.n70 VTAIL.n69 585
R75 VTAIL.n91 VTAIL.n90 585
R76 VTAIL.n94 VTAIL.n93 585
R77 VTAIL.n92 VTAIL.n66 585
R78 VTAIL.n99 VTAIL.n65 585
R79 VTAIL.n101 VTAIL.n100 585
R80 VTAIL.n103 VTAIL.n102 585
R81 VTAIL.n62 VTAIL.n61 585
R82 VTAIL.n109 VTAIL.n108 585
R83 VTAIL.n111 VTAIL.n110 585
R84 VTAIL.n135 VTAIL.n134 585
R85 VTAIL.n132 VTAIL.n131 585
R86 VTAIL.n141 VTAIL.n140 585
R87 VTAIL.n143 VTAIL.n142 585
R88 VTAIL.n128 VTAIL.n127 585
R89 VTAIL.n149 VTAIL.n148 585
R90 VTAIL.n152 VTAIL.n151 585
R91 VTAIL.n150 VTAIL.n124 585
R92 VTAIL.n157 VTAIL.n123 585
R93 VTAIL.n159 VTAIL.n158 585
R94 VTAIL.n161 VTAIL.n160 585
R95 VTAIL.n120 VTAIL.n119 585
R96 VTAIL.n167 VTAIL.n166 585
R97 VTAIL.n169 VTAIL.n168 585
R98 VTAIL.n401 VTAIL.n400 585
R99 VTAIL.n399 VTAIL.n398 585
R100 VTAIL.n352 VTAIL.n351 585
R101 VTAIL.n393 VTAIL.n392 585
R102 VTAIL.n391 VTAIL.n390 585
R103 VTAIL.n389 VTAIL.n355 585
R104 VTAIL.n359 VTAIL.n356 585
R105 VTAIL.n384 VTAIL.n383 585
R106 VTAIL.n382 VTAIL.n381 585
R107 VTAIL.n361 VTAIL.n360 585
R108 VTAIL.n376 VTAIL.n375 585
R109 VTAIL.n374 VTAIL.n373 585
R110 VTAIL.n365 VTAIL.n364 585
R111 VTAIL.n368 VTAIL.n367 585
R112 VTAIL.n343 VTAIL.n342 585
R113 VTAIL.n341 VTAIL.n340 585
R114 VTAIL.n294 VTAIL.n293 585
R115 VTAIL.n335 VTAIL.n334 585
R116 VTAIL.n333 VTAIL.n332 585
R117 VTAIL.n331 VTAIL.n297 585
R118 VTAIL.n301 VTAIL.n298 585
R119 VTAIL.n326 VTAIL.n325 585
R120 VTAIL.n324 VTAIL.n323 585
R121 VTAIL.n303 VTAIL.n302 585
R122 VTAIL.n318 VTAIL.n317 585
R123 VTAIL.n316 VTAIL.n315 585
R124 VTAIL.n307 VTAIL.n306 585
R125 VTAIL.n310 VTAIL.n309 585
R126 VTAIL.n285 VTAIL.n284 585
R127 VTAIL.n283 VTAIL.n282 585
R128 VTAIL.n236 VTAIL.n235 585
R129 VTAIL.n277 VTAIL.n276 585
R130 VTAIL.n275 VTAIL.n274 585
R131 VTAIL.n273 VTAIL.n239 585
R132 VTAIL.n243 VTAIL.n240 585
R133 VTAIL.n268 VTAIL.n267 585
R134 VTAIL.n266 VTAIL.n265 585
R135 VTAIL.n245 VTAIL.n244 585
R136 VTAIL.n260 VTAIL.n259 585
R137 VTAIL.n258 VTAIL.n257 585
R138 VTAIL.n249 VTAIL.n248 585
R139 VTAIL.n252 VTAIL.n251 585
R140 VTAIL.n227 VTAIL.n226 585
R141 VTAIL.n225 VTAIL.n224 585
R142 VTAIL.n178 VTAIL.n177 585
R143 VTAIL.n219 VTAIL.n218 585
R144 VTAIL.n217 VTAIL.n216 585
R145 VTAIL.n215 VTAIL.n181 585
R146 VTAIL.n185 VTAIL.n182 585
R147 VTAIL.n210 VTAIL.n209 585
R148 VTAIL.n208 VTAIL.n207 585
R149 VTAIL.n187 VTAIL.n186 585
R150 VTAIL.n202 VTAIL.n201 585
R151 VTAIL.n200 VTAIL.n199 585
R152 VTAIL.n191 VTAIL.n190 585
R153 VTAIL.n194 VTAIL.n193 585
R154 VTAIL.t3 VTAIL.n366 329.038
R155 VTAIL.t6 VTAIL.n308 329.038
R156 VTAIL.t7 VTAIL.n250 329.038
R157 VTAIL.t2 VTAIL.n192 329.038
R158 VTAIL.t0 VTAIL.n423 329.038
R159 VTAIL.t1 VTAIL.n17 329.038
R160 VTAIL.t4 VTAIL.n75 329.038
R161 VTAIL.t5 VTAIL.n133 329.038
R162 VTAIL.n424 VTAIL.n421 171.744
R163 VTAIL.n431 VTAIL.n421 171.744
R164 VTAIL.n432 VTAIL.n431 171.744
R165 VTAIL.n432 VTAIL.n417 171.744
R166 VTAIL.n439 VTAIL.n417 171.744
R167 VTAIL.n441 VTAIL.n439 171.744
R168 VTAIL.n441 VTAIL.n440 171.744
R169 VTAIL.n440 VTAIL.n413 171.744
R170 VTAIL.n449 VTAIL.n413 171.744
R171 VTAIL.n450 VTAIL.n449 171.744
R172 VTAIL.n450 VTAIL.n409 171.744
R173 VTAIL.n457 VTAIL.n409 171.744
R174 VTAIL.n458 VTAIL.n457 171.744
R175 VTAIL.n18 VTAIL.n15 171.744
R176 VTAIL.n25 VTAIL.n15 171.744
R177 VTAIL.n26 VTAIL.n25 171.744
R178 VTAIL.n26 VTAIL.n11 171.744
R179 VTAIL.n33 VTAIL.n11 171.744
R180 VTAIL.n35 VTAIL.n33 171.744
R181 VTAIL.n35 VTAIL.n34 171.744
R182 VTAIL.n34 VTAIL.n7 171.744
R183 VTAIL.n43 VTAIL.n7 171.744
R184 VTAIL.n44 VTAIL.n43 171.744
R185 VTAIL.n44 VTAIL.n3 171.744
R186 VTAIL.n51 VTAIL.n3 171.744
R187 VTAIL.n52 VTAIL.n51 171.744
R188 VTAIL.n76 VTAIL.n73 171.744
R189 VTAIL.n83 VTAIL.n73 171.744
R190 VTAIL.n84 VTAIL.n83 171.744
R191 VTAIL.n84 VTAIL.n69 171.744
R192 VTAIL.n91 VTAIL.n69 171.744
R193 VTAIL.n93 VTAIL.n91 171.744
R194 VTAIL.n93 VTAIL.n92 171.744
R195 VTAIL.n92 VTAIL.n65 171.744
R196 VTAIL.n101 VTAIL.n65 171.744
R197 VTAIL.n102 VTAIL.n101 171.744
R198 VTAIL.n102 VTAIL.n61 171.744
R199 VTAIL.n109 VTAIL.n61 171.744
R200 VTAIL.n110 VTAIL.n109 171.744
R201 VTAIL.n134 VTAIL.n131 171.744
R202 VTAIL.n141 VTAIL.n131 171.744
R203 VTAIL.n142 VTAIL.n141 171.744
R204 VTAIL.n142 VTAIL.n127 171.744
R205 VTAIL.n149 VTAIL.n127 171.744
R206 VTAIL.n151 VTAIL.n149 171.744
R207 VTAIL.n151 VTAIL.n150 171.744
R208 VTAIL.n150 VTAIL.n123 171.744
R209 VTAIL.n159 VTAIL.n123 171.744
R210 VTAIL.n160 VTAIL.n159 171.744
R211 VTAIL.n160 VTAIL.n119 171.744
R212 VTAIL.n167 VTAIL.n119 171.744
R213 VTAIL.n168 VTAIL.n167 171.744
R214 VTAIL.n400 VTAIL.n399 171.744
R215 VTAIL.n399 VTAIL.n351 171.744
R216 VTAIL.n392 VTAIL.n351 171.744
R217 VTAIL.n392 VTAIL.n391 171.744
R218 VTAIL.n391 VTAIL.n355 171.744
R219 VTAIL.n359 VTAIL.n355 171.744
R220 VTAIL.n383 VTAIL.n359 171.744
R221 VTAIL.n383 VTAIL.n382 171.744
R222 VTAIL.n382 VTAIL.n360 171.744
R223 VTAIL.n375 VTAIL.n360 171.744
R224 VTAIL.n375 VTAIL.n374 171.744
R225 VTAIL.n374 VTAIL.n364 171.744
R226 VTAIL.n367 VTAIL.n364 171.744
R227 VTAIL.n342 VTAIL.n341 171.744
R228 VTAIL.n341 VTAIL.n293 171.744
R229 VTAIL.n334 VTAIL.n293 171.744
R230 VTAIL.n334 VTAIL.n333 171.744
R231 VTAIL.n333 VTAIL.n297 171.744
R232 VTAIL.n301 VTAIL.n297 171.744
R233 VTAIL.n325 VTAIL.n301 171.744
R234 VTAIL.n325 VTAIL.n324 171.744
R235 VTAIL.n324 VTAIL.n302 171.744
R236 VTAIL.n317 VTAIL.n302 171.744
R237 VTAIL.n317 VTAIL.n316 171.744
R238 VTAIL.n316 VTAIL.n306 171.744
R239 VTAIL.n309 VTAIL.n306 171.744
R240 VTAIL.n284 VTAIL.n283 171.744
R241 VTAIL.n283 VTAIL.n235 171.744
R242 VTAIL.n276 VTAIL.n235 171.744
R243 VTAIL.n276 VTAIL.n275 171.744
R244 VTAIL.n275 VTAIL.n239 171.744
R245 VTAIL.n243 VTAIL.n239 171.744
R246 VTAIL.n267 VTAIL.n243 171.744
R247 VTAIL.n267 VTAIL.n266 171.744
R248 VTAIL.n266 VTAIL.n244 171.744
R249 VTAIL.n259 VTAIL.n244 171.744
R250 VTAIL.n259 VTAIL.n258 171.744
R251 VTAIL.n258 VTAIL.n248 171.744
R252 VTAIL.n251 VTAIL.n248 171.744
R253 VTAIL.n226 VTAIL.n225 171.744
R254 VTAIL.n225 VTAIL.n177 171.744
R255 VTAIL.n218 VTAIL.n177 171.744
R256 VTAIL.n218 VTAIL.n217 171.744
R257 VTAIL.n217 VTAIL.n181 171.744
R258 VTAIL.n185 VTAIL.n181 171.744
R259 VTAIL.n209 VTAIL.n185 171.744
R260 VTAIL.n209 VTAIL.n208 171.744
R261 VTAIL.n208 VTAIL.n186 171.744
R262 VTAIL.n201 VTAIL.n186 171.744
R263 VTAIL.n201 VTAIL.n200 171.744
R264 VTAIL.n200 VTAIL.n190 171.744
R265 VTAIL.n193 VTAIL.n190 171.744
R266 VTAIL.n424 VTAIL.t0 85.8723
R267 VTAIL.n18 VTAIL.t1 85.8723
R268 VTAIL.n76 VTAIL.t4 85.8723
R269 VTAIL.n134 VTAIL.t5 85.8723
R270 VTAIL.n367 VTAIL.t3 85.8723
R271 VTAIL.n309 VTAIL.t6 85.8723
R272 VTAIL.n251 VTAIL.t7 85.8723
R273 VTAIL.n193 VTAIL.t2 85.8723
R274 VTAIL.n463 VTAIL.n462 31.2157
R275 VTAIL.n57 VTAIL.n56 31.2157
R276 VTAIL.n115 VTAIL.n114 31.2157
R277 VTAIL.n173 VTAIL.n172 31.2157
R278 VTAIL.n405 VTAIL.n404 31.2157
R279 VTAIL.n347 VTAIL.n346 31.2157
R280 VTAIL.n289 VTAIL.n288 31.2157
R281 VTAIL.n231 VTAIL.n230 31.2157
R282 VTAIL.n463 VTAIL.n405 25.2289
R283 VTAIL.n231 VTAIL.n173 25.2289
R284 VTAIL.n448 VTAIL.n447 13.1884
R285 VTAIL.n42 VTAIL.n41 13.1884
R286 VTAIL.n100 VTAIL.n99 13.1884
R287 VTAIL.n158 VTAIL.n157 13.1884
R288 VTAIL.n390 VTAIL.n389 13.1884
R289 VTAIL.n332 VTAIL.n331 13.1884
R290 VTAIL.n274 VTAIL.n273 13.1884
R291 VTAIL.n216 VTAIL.n215 13.1884
R292 VTAIL.n446 VTAIL.n414 12.8005
R293 VTAIL.n451 VTAIL.n412 12.8005
R294 VTAIL.n40 VTAIL.n8 12.8005
R295 VTAIL.n45 VTAIL.n6 12.8005
R296 VTAIL.n98 VTAIL.n66 12.8005
R297 VTAIL.n103 VTAIL.n64 12.8005
R298 VTAIL.n156 VTAIL.n124 12.8005
R299 VTAIL.n161 VTAIL.n122 12.8005
R300 VTAIL.n393 VTAIL.n354 12.8005
R301 VTAIL.n388 VTAIL.n356 12.8005
R302 VTAIL.n335 VTAIL.n296 12.8005
R303 VTAIL.n330 VTAIL.n298 12.8005
R304 VTAIL.n277 VTAIL.n238 12.8005
R305 VTAIL.n272 VTAIL.n240 12.8005
R306 VTAIL.n219 VTAIL.n180 12.8005
R307 VTAIL.n214 VTAIL.n182 12.8005
R308 VTAIL.n443 VTAIL.n442 12.0247
R309 VTAIL.n452 VTAIL.n410 12.0247
R310 VTAIL.n37 VTAIL.n36 12.0247
R311 VTAIL.n46 VTAIL.n4 12.0247
R312 VTAIL.n95 VTAIL.n94 12.0247
R313 VTAIL.n104 VTAIL.n62 12.0247
R314 VTAIL.n153 VTAIL.n152 12.0247
R315 VTAIL.n162 VTAIL.n120 12.0247
R316 VTAIL.n394 VTAIL.n352 12.0247
R317 VTAIL.n385 VTAIL.n384 12.0247
R318 VTAIL.n336 VTAIL.n294 12.0247
R319 VTAIL.n327 VTAIL.n326 12.0247
R320 VTAIL.n278 VTAIL.n236 12.0247
R321 VTAIL.n269 VTAIL.n268 12.0247
R322 VTAIL.n220 VTAIL.n178 12.0247
R323 VTAIL.n211 VTAIL.n210 12.0247
R324 VTAIL.n438 VTAIL.n416 11.249
R325 VTAIL.n456 VTAIL.n455 11.249
R326 VTAIL.n32 VTAIL.n10 11.249
R327 VTAIL.n50 VTAIL.n49 11.249
R328 VTAIL.n90 VTAIL.n68 11.249
R329 VTAIL.n108 VTAIL.n107 11.249
R330 VTAIL.n148 VTAIL.n126 11.249
R331 VTAIL.n166 VTAIL.n165 11.249
R332 VTAIL.n398 VTAIL.n397 11.249
R333 VTAIL.n381 VTAIL.n358 11.249
R334 VTAIL.n340 VTAIL.n339 11.249
R335 VTAIL.n323 VTAIL.n300 11.249
R336 VTAIL.n282 VTAIL.n281 11.249
R337 VTAIL.n265 VTAIL.n242 11.249
R338 VTAIL.n224 VTAIL.n223 11.249
R339 VTAIL.n207 VTAIL.n184 11.249
R340 VTAIL.n425 VTAIL.n423 10.7239
R341 VTAIL.n19 VTAIL.n17 10.7239
R342 VTAIL.n77 VTAIL.n75 10.7239
R343 VTAIL.n135 VTAIL.n133 10.7239
R344 VTAIL.n368 VTAIL.n366 10.7239
R345 VTAIL.n310 VTAIL.n308 10.7239
R346 VTAIL.n252 VTAIL.n250 10.7239
R347 VTAIL.n194 VTAIL.n192 10.7239
R348 VTAIL.n437 VTAIL.n418 10.4732
R349 VTAIL.n459 VTAIL.n408 10.4732
R350 VTAIL.n31 VTAIL.n12 10.4732
R351 VTAIL.n53 VTAIL.n2 10.4732
R352 VTAIL.n89 VTAIL.n70 10.4732
R353 VTAIL.n111 VTAIL.n60 10.4732
R354 VTAIL.n147 VTAIL.n128 10.4732
R355 VTAIL.n169 VTAIL.n118 10.4732
R356 VTAIL.n401 VTAIL.n350 10.4732
R357 VTAIL.n380 VTAIL.n361 10.4732
R358 VTAIL.n343 VTAIL.n292 10.4732
R359 VTAIL.n322 VTAIL.n303 10.4732
R360 VTAIL.n285 VTAIL.n234 10.4732
R361 VTAIL.n264 VTAIL.n245 10.4732
R362 VTAIL.n227 VTAIL.n176 10.4732
R363 VTAIL.n206 VTAIL.n187 10.4732
R364 VTAIL.n434 VTAIL.n433 9.69747
R365 VTAIL.n460 VTAIL.n406 9.69747
R366 VTAIL.n28 VTAIL.n27 9.69747
R367 VTAIL.n54 VTAIL.n0 9.69747
R368 VTAIL.n86 VTAIL.n85 9.69747
R369 VTAIL.n112 VTAIL.n58 9.69747
R370 VTAIL.n144 VTAIL.n143 9.69747
R371 VTAIL.n170 VTAIL.n116 9.69747
R372 VTAIL.n402 VTAIL.n348 9.69747
R373 VTAIL.n377 VTAIL.n376 9.69747
R374 VTAIL.n344 VTAIL.n290 9.69747
R375 VTAIL.n319 VTAIL.n318 9.69747
R376 VTAIL.n286 VTAIL.n232 9.69747
R377 VTAIL.n261 VTAIL.n260 9.69747
R378 VTAIL.n228 VTAIL.n174 9.69747
R379 VTAIL.n203 VTAIL.n202 9.69747
R380 VTAIL.n462 VTAIL.n461 9.45567
R381 VTAIL.n56 VTAIL.n55 9.45567
R382 VTAIL.n114 VTAIL.n113 9.45567
R383 VTAIL.n172 VTAIL.n171 9.45567
R384 VTAIL.n404 VTAIL.n403 9.45567
R385 VTAIL.n346 VTAIL.n345 9.45567
R386 VTAIL.n288 VTAIL.n287 9.45567
R387 VTAIL.n230 VTAIL.n229 9.45567
R388 VTAIL.n461 VTAIL.n460 9.3005
R389 VTAIL.n408 VTAIL.n407 9.3005
R390 VTAIL.n455 VTAIL.n454 9.3005
R391 VTAIL.n453 VTAIL.n452 9.3005
R392 VTAIL.n412 VTAIL.n411 9.3005
R393 VTAIL.n427 VTAIL.n426 9.3005
R394 VTAIL.n429 VTAIL.n428 9.3005
R395 VTAIL.n420 VTAIL.n419 9.3005
R396 VTAIL.n435 VTAIL.n434 9.3005
R397 VTAIL.n437 VTAIL.n436 9.3005
R398 VTAIL.n416 VTAIL.n415 9.3005
R399 VTAIL.n444 VTAIL.n443 9.3005
R400 VTAIL.n446 VTAIL.n445 9.3005
R401 VTAIL.n55 VTAIL.n54 9.3005
R402 VTAIL.n2 VTAIL.n1 9.3005
R403 VTAIL.n49 VTAIL.n48 9.3005
R404 VTAIL.n47 VTAIL.n46 9.3005
R405 VTAIL.n6 VTAIL.n5 9.3005
R406 VTAIL.n21 VTAIL.n20 9.3005
R407 VTAIL.n23 VTAIL.n22 9.3005
R408 VTAIL.n14 VTAIL.n13 9.3005
R409 VTAIL.n29 VTAIL.n28 9.3005
R410 VTAIL.n31 VTAIL.n30 9.3005
R411 VTAIL.n10 VTAIL.n9 9.3005
R412 VTAIL.n38 VTAIL.n37 9.3005
R413 VTAIL.n40 VTAIL.n39 9.3005
R414 VTAIL.n113 VTAIL.n112 9.3005
R415 VTAIL.n60 VTAIL.n59 9.3005
R416 VTAIL.n107 VTAIL.n106 9.3005
R417 VTAIL.n105 VTAIL.n104 9.3005
R418 VTAIL.n64 VTAIL.n63 9.3005
R419 VTAIL.n79 VTAIL.n78 9.3005
R420 VTAIL.n81 VTAIL.n80 9.3005
R421 VTAIL.n72 VTAIL.n71 9.3005
R422 VTAIL.n87 VTAIL.n86 9.3005
R423 VTAIL.n89 VTAIL.n88 9.3005
R424 VTAIL.n68 VTAIL.n67 9.3005
R425 VTAIL.n96 VTAIL.n95 9.3005
R426 VTAIL.n98 VTAIL.n97 9.3005
R427 VTAIL.n171 VTAIL.n170 9.3005
R428 VTAIL.n118 VTAIL.n117 9.3005
R429 VTAIL.n165 VTAIL.n164 9.3005
R430 VTAIL.n163 VTAIL.n162 9.3005
R431 VTAIL.n122 VTAIL.n121 9.3005
R432 VTAIL.n137 VTAIL.n136 9.3005
R433 VTAIL.n139 VTAIL.n138 9.3005
R434 VTAIL.n130 VTAIL.n129 9.3005
R435 VTAIL.n145 VTAIL.n144 9.3005
R436 VTAIL.n147 VTAIL.n146 9.3005
R437 VTAIL.n126 VTAIL.n125 9.3005
R438 VTAIL.n154 VTAIL.n153 9.3005
R439 VTAIL.n156 VTAIL.n155 9.3005
R440 VTAIL.n370 VTAIL.n369 9.3005
R441 VTAIL.n372 VTAIL.n371 9.3005
R442 VTAIL.n363 VTAIL.n362 9.3005
R443 VTAIL.n378 VTAIL.n377 9.3005
R444 VTAIL.n380 VTAIL.n379 9.3005
R445 VTAIL.n358 VTAIL.n357 9.3005
R446 VTAIL.n386 VTAIL.n385 9.3005
R447 VTAIL.n388 VTAIL.n387 9.3005
R448 VTAIL.n403 VTAIL.n402 9.3005
R449 VTAIL.n350 VTAIL.n349 9.3005
R450 VTAIL.n397 VTAIL.n396 9.3005
R451 VTAIL.n395 VTAIL.n394 9.3005
R452 VTAIL.n354 VTAIL.n353 9.3005
R453 VTAIL.n312 VTAIL.n311 9.3005
R454 VTAIL.n314 VTAIL.n313 9.3005
R455 VTAIL.n305 VTAIL.n304 9.3005
R456 VTAIL.n320 VTAIL.n319 9.3005
R457 VTAIL.n322 VTAIL.n321 9.3005
R458 VTAIL.n300 VTAIL.n299 9.3005
R459 VTAIL.n328 VTAIL.n327 9.3005
R460 VTAIL.n330 VTAIL.n329 9.3005
R461 VTAIL.n345 VTAIL.n344 9.3005
R462 VTAIL.n292 VTAIL.n291 9.3005
R463 VTAIL.n339 VTAIL.n338 9.3005
R464 VTAIL.n337 VTAIL.n336 9.3005
R465 VTAIL.n296 VTAIL.n295 9.3005
R466 VTAIL.n254 VTAIL.n253 9.3005
R467 VTAIL.n256 VTAIL.n255 9.3005
R468 VTAIL.n247 VTAIL.n246 9.3005
R469 VTAIL.n262 VTAIL.n261 9.3005
R470 VTAIL.n264 VTAIL.n263 9.3005
R471 VTAIL.n242 VTAIL.n241 9.3005
R472 VTAIL.n270 VTAIL.n269 9.3005
R473 VTAIL.n272 VTAIL.n271 9.3005
R474 VTAIL.n287 VTAIL.n286 9.3005
R475 VTAIL.n234 VTAIL.n233 9.3005
R476 VTAIL.n281 VTAIL.n280 9.3005
R477 VTAIL.n279 VTAIL.n278 9.3005
R478 VTAIL.n238 VTAIL.n237 9.3005
R479 VTAIL.n196 VTAIL.n195 9.3005
R480 VTAIL.n198 VTAIL.n197 9.3005
R481 VTAIL.n189 VTAIL.n188 9.3005
R482 VTAIL.n204 VTAIL.n203 9.3005
R483 VTAIL.n206 VTAIL.n205 9.3005
R484 VTAIL.n184 VTAIL.n183 9.3005
R485 VTAIL.n212 VTAIL.n211 9.3005
R486 VTAIL.n214 VTAIL.n213 9.3005
R487 VTAIL.n229 VTAIL.n228 9.3005
R488 VTAIL.n176 VTAIL.n175 9.3005
R489 VTAIL.n223 VTAIL.n222 9.3005
R490 VTAIL.n221 VTAIL.n220 9.3005
R491 VTAIL.n180 VTAIL.n179 9.3005
R492 VTAIL.n430 VTAIL.n420 8.92171
R493 VTAIL.n24 VTAIL.n14 8.92171
R494 VTAIL.n82 VTAIL.n72 8.92171
R495 VTAIL.n140 VTAIL.n130 8.92171
R496 VTAIL.n373 VTAIL.n363 8.92171
R497 VTAIL.n315 VTAIL.n305 8.92171
R498 VTAIL.n257 VTAIL.n247 8.92171
R499 VTAIL.n199 VTAIL.n189 8.92171
R500 VTAIL.n429 VTAIL.n422 8.14595
R501 VTAIL.n23 VTAIL.n16 8.14595
R502 VTAIL.n81 VTAIL.n74 8.14595
R503 VTAIL.n139 VTAIL.n132 8.14595
R504 VTAIL.n372 VTAIL.n365 8.14595
R505 VTAIL.n314 VTAIL.n307 8.14595
R506 VTAIL.n256 VTAIL.n249 8.14595
R507 VTAIL.n198 VTAIL.n191 8.14595
R508 VTAIL.n426 VTAIL.n425 7.3702
R509 VTAIL.n20 VTAIL.n19 7.3702
R510 VTAIL.n78 VTAIL.n77 7.3702
R511 VTAIL.n136 VTAIL.n135 7.3702
R512 VTAIL.n369 VTAIL.n368 7.3702
R513 VTAIL.n311 VTAIL.n310 7.3702
R514 VTAIL.n253 VTAIL.n252 7.3702
R515 VTAIL.n195 VTAIL.n194 7.3702
R516 VTAIL.n426 VTAIL.n422 5.81868
R517 VTAIL.n20 VTAIL.n16 5.81868
R518 VTAIL.n78 VTAIL.n74 5.81868
R519 VTAIL.n136 VTAIL.n132 5.81868
R520 VTAIL.n369 VTAIL.n365 5.81868
R521 VTAIL.n311 VTAIL.n307 5.81868
R522 VTAIL.n253 VTAIL.n249 5.81868
R523 VTAIL.n195 VTAIL.n191 5.81868
R524 VTAIL.n430 VTAIL.n429 5.04292
R525 VTAIL.n24 VTAIL.n23 5.04292
R526 VTAIL.n82 VTAIL.n81 5.04292
R527 VTAIL.n140 VTAIL.n139 5.04292
R528 VTAIL.n373 VTAIL.n372 5.04292
R529 VTAIL.n315 VTAIL.n314 5.04292
R530 VTAIL.n257 VTAIL.n256 5.04292
R531 VTAIL.n199 VTAIL.n198 5.04292
R532 VTAIL.n433 VTAIL.n420 4.26717
R533 VTAIL.n462 VTAIL.n406 4.26717
R534 VTAIL.n27 VTAIL.n14 4.26717
R535 VTAIL.n56 VTAIL.n0 4.26717
R536 VTAIL.n85 VTAIL.n72 4.26717
R537 VTAIL.n114 VTAIL.n58 4.26717
R538 VTAIL.n143 VTAIL.n130 4.26717
R539 VTAIL.n172 VTAIL.n116 4.26717
R540 VTAIL.n404 VTAIL.n348 4.26717
R541 VTAIL.n376 VTAIL.n363 4.26717
R542 VTAIL.n346 VTAIL.n290 4.26717
R543 VTAIL.n318 VTAIL.n305 4.26717
R544 VTAIL.n288 VTAIL.n232 4.26717
R545 VTAIL.n260 VTAIL.n247 4.26717
R546 VTAIL.n230 VTAIL.n174 4.26717
R547 VTAIL.n202 VTAIL.n189 4.26717
R548 VTAIL.n289 VTAIL.n231 3.69878
R549 VTAIL.n405 VTAIL.n347 3.69878
R550 VTAIL.n173 VTAIL.n115 3.69878
R551 VTAIL.n434 VTAIL.n418 3.49141
R552 VTAIL.n460 VTAIL.n459 3.49141
R553 VTAIL.n28 VTAIL.n12 3.49141
R554 VTAIL.n54 VTAIL.n53 3.49141
R555 VTAIL.n86 VTAIL.n70 3.49141
R556 VTAIL.n112 VTAIL.n111 3.49141
R557 VTAIL.n144 VTAIL.n128 3.49141
R558 VTAIL.n170 VTAIL.n169 3.49141
R559 VTAIL.n402 VTAIL.n401 3.49141
R560 VTAIL.n377 VTAIL.n361 3.49141
R561 VTAIL.n344 VTAIL.n343 3.49141
R562 VTAIL.n319 VTAIL.n303 3.49141
R563 VTAIL.n286 VTAIL.n285 3.49141
R564 VTAIL.n261 VTAIL.n245 3.49141
R565 VTAIL.n228 VTAIL.n227 3.49141
R566 VTAIL.n203 VTAIL.n187 3.49141
R567 VTAIL.n438 VTAIL.n437 2.71565
R568 VTAIL.n456 VTAIL.n408 2.71565
R569 VTAIL.n32 VTAIL.n31 2.71565
R570 VTAIL.n50 VTAIL.n2 2.71565
R571 VTAIL.n90 VTAIL.n89 2.71565
R572 VTAIL.n108 VTAIL.n60 2.71565
R573 VTAIL.n148 VTAIL.n147 2.71565
R574 VTAIL.n166 VTAIL.n118 2.71565
R575 VTAIL.n398 VTAIL.n350 2.71565
R576 VTAIL.n381 VTAIL.n380 2.71565
R577 VTAIL.n340 VTAIL.n292 2.71565
R578 VTAIL.n323 VTAIL.n322 2.71565
R579 VTAIL.n282 VTAIL.n234 2.71565
R580 VTAIL.n265 VTAIL.n264 2.71565
R581 VTAIL.n224 VTAIL.n176 2.71565
R582 VTAIL.n207 VTAIL.n206 2.71565
R583 VTAIL.n427 VTAIL.n423 2.41282
R584 VTAIL.n21 VTAIL.n17 2.41282
R585 VTAIL.n79 VTAIL.n75 2.41282
R586 VTAIL.n137 VTAIL.n133 2.41282
R587 VTAIL.n370 VTAIL.n366 2.41282
R588 VTAIL.n312 VTAIL.n308 2.41282
R589 VTAIL.n254 VTAIL.n250 2.41282
R590 VTAIL.n196 VTAIL.n192 2.41282
R591 VTAIL.n442 VTAIL.n416 1.93989
R592 VTAIL.n455 VTAIL.n410 1.93989
R593 VTAIL.n36 VTAIL.n10 1.93989
R594 VTAIL.n49 VTAIL.n4 1.93989
R595 VTAIL.n94 VTAIL.n68 1.93989
R596 VTAIL.n107 VTAIL.n62 1.93989
R597 VTAIL.n152 VTAIL.n126 1.93989
R598 VTAIL.n165 VTAIL.n120 1.93989
R599 VTAIL.n397 VTAIL.n352 1.93989
R600 VTAIL.n384 VTAIL.n358 1.93989
R601 VTAIL.n339 VTAIL.n294 1.93989
R602 VTAIL.n326 VTAIL.n300 1.93989
R603 VTAIL.n281 VTAIL.n236 1.93989
R604 VTAIL.n268 VTAIL.n242 1.93989
R605 VTAIL.n223 VTAIL.n178 1.93989
R606 VTAIL.n210 VTAIL.n184 1.93989
R607 VTAIL VTAIL.n57 1.90783
R608 VTAIL VTAIL.n463 1.79145
R609 VTAIL.n443 VTAIL.n414 1.16414
R610 VTAIL.n452 VTAIL.n451 1.16414
R611 VTAIL.n37 VTAIL.n8 1.16414
R612 VTAIL.n46 VTAIL.n45 1.16414
R613 VTAIL.n95 VTAIL.n66 1.16414
R614 VTAIL.n104 VTAIL.n103 1.16414
R615 VTAIL.n153 VTAIL.n124 1.16414
R616 VTAIL.n162 VTAIL.n161 1.16414
R617 VTAIL.n394 VTAIL.n393 1.16414
R618 VTAIL.n385 VTAIL.n356 1.16414
R619 VTAIL.n336 VTAIL.n335 1.16414
R620 VTAIL.n327 VTAIL.n298 1.16414
R621 VTAIL.n278 VTAIL.n277 1.16414
R622 VTAIL.n269 VTAIL.n240 1.16414
R623 VTAIL.n220 VTAIL.n219 1.16414
R624 VTAIL.n211 VTAIL.n182 1.16414
R625 VTAIL.n347 VTAIL.n289 0.470328
R626 VTAIL.n115 VTAIL.n57 0.470328
R627 VTAIL.n447 VTAIL.n446 0.388379
R628 VTAIL.n448 VTAIL.n412 0.388379
R629 VTAIL.n41 VTAIL.n40 0.388379
R630 VTAIL.n42 VTAIL.n6 0.388379
R631 VTAIL.n99 VTAIL.n98 0.388379
R632 VTAIL.n100 VTAIL.n64 0.388379
R633 VTAIL.n157 VTAIL.n156 0.388379
R634 VTAIL.n158 VTAIL.n122 0.388379
R635 VTAIL.n390 VTAIL.n354 0.388379
R636 VTAIL.n389 VTAIL.n388 0.388379
R637 VTAIL.n332 VTAIL.n296 0.388379
R638 VTAIL.n331 VTAIL.n330 0.388379
R639 VTAIL.n274 VTAIL.n238 0.388379
R640 VTAIL.n273 VTAIL.n272 0.388379
R641 VTAIL.n216 VTAIL.n180 0.388379
R642 VTAIL.n215 VTAIL.n214 0.388379
R643 VTAIL.n428 VTAIL.n427 0.155672
R644 VTAIL.n428 VTAIL.n419 0.155672
R645 VTAIL.n435 VTAIL.n419 0.155672
R646 VTAIL.n436 VTAIL.n435 0.155672
R647 VTAIL.n436 VTAIL.n415 0.155672
R648 VTAIL.n444 VTAIL.n415 0.155672
R649 VTAIL.n445 VTAIL.n444 0.155672
R650 VTAIL.n445 VTAIL.n411 0.155672
R651 VTAIL.n453 VTAIL.n411 0.155672
R652 VTAIL.n454 VTAIL.n453 0.155672
R653 VTAIL.n454 VTAIL.n407 0.155672
R654 VTAIL.n461 VTAIL.n407 0.155672
R655 VTAIL.n22 VTAIL.n21 0.155672
R656 VTAIL.n22 VTAIL.n13 0.155672
R657 VTAIL.n29 VTAIL.n13 0.155672
R658 VTAIL.n30 VTAIL.n29 0.155672
R659 VTAIL.n30 VTAIL.n9 0.155672
R660 VTAIL.n38 VTAIL.n9 0.155672
R661 VTAIL.n39 VTAIL.n38 0.155672
R662 VTAIL.n39 VTAIL.n5 0.155672
R663 VTAIL.n47 VTAIL.n5 0.155672
R664 VTAIL.n48 VTAIL.n47 0.155672
R665 VTAIL.n48 VTAIL.n1 0.155672
R666 VTAIL.n55 VTAIL.n1 0.155672
R667 VTAIL.n80 VTAIL.n79 0.155672
R668 VTAIL.n80 VTAIL.n71 0.155672
R669 VTAIL.n87 VTAIL.n71 0.155672
R670 VTAIL.n88 VTAIL.n87 0.155672
R671 VTAIL.n88 VTAIL.n67 0.155672
R672 VTAIL.n96 VTAIL.n67 0.155672
R673 VTAIL.n97 VTAIL.n96 0.155672
R674 VTAIL.n97 VTAIL.n63 0.155672
R675 VTAIL.n105 VTAIL.n63 0.155672
R676 VTAIL.n106 VTAIL.n105 0.155672
R677 VTAIL.n106 VTAIL.n59 0.155672
R678 VTAIL.n113 VTAIL.n59 0.155672
R679 VTAIL.n138 VTAIL.n137 0.155672
R680 VTAIL.n138 VTAIL.n129 0.155672
R681 VTAIL.n145 VTAIL.n129 0.155672
R682 VTAIL.n146 VTAIL.n145 0.155672
R683 VTAIL.n146 VTAIL.n125 0.155672
R684 VTAIL.n154 VTAIL.n125 0.155672
R685 VTAIL.n155 VTAIL.n154 0.155672
R686 VTAIL.n155 VTAIL.n121 0.155672
R687 VTAIL.n163 VTAIL.n121 0.155672
R688 VTAIL.n164 VTAIL.n163 0.155672
R689 VTAIL.n164 VTAIL.n117 0.155672
R690 VTAIL.n171 VTAIL.n117 0.155672
R691 VTAIL.n403 VTAIL.n349 0.155672
R692 VTAIL.n396 VTAIL.n349 0.155672
R693 VTAIL.n396 VTAIL.n395 0.155672
R694 VTAIL.n395 VTAIL.n353 0.155672
R695 VTAIL.n387 VTAIL.n353 0.155672
R696 VTAIL.n387 VTAIL.n386 0.155672
R697 VTAIL.n386 VTAIL.n357 0.155672
R698 VTAIL.n379 VTAIL.n357 0.155672
R699 VTAIL.n379 VTAIL.n378 0.155672
R700 VTAIL.n378 VTAIL.n362 0.155672
R701 VTAIL.n371 VTAIL.n362 0.155672
R702 VTAIL.n371 VTAIL.n370 0.155672
R703 VTAIL.n345 VTAIL.n291 0.155672
R704 VTAIL.n338 VTAIL.n291 0.155672
R705 VTAIL.n338 VTAIL.n337 0.155672
R706 VTAIL.n337 VTAIL.n295 0.155672
R707 VTAIL.n329 VTAIL.n295 0.155672
R708 VTAIL.n329 VTAIL.n328 0.155672
R709 VTAIL.n328 VTAIL.n299 0.155672
R710 VTAIL.n321 VTAIL.n299 0.155672
R711 VTAIL.n321 VTAIL.n320 0.155672
R712 VTAIL.n320 VTAIL.n304 0.155672
R713 VTAIL.n313 VTAIL.n304 0.155672
R714 VTAIL.n313 VTAIL.n312 0.155672
R715 VTAIL.n287 VTAIL.n233 0.155672
R716 VTAIL.n280 VTAIL.n233 0.155672
R717 VTAIL.n280 VTAIL.n279 0.155672
R718 VTAIL.n279 VTAIL.n237 0.155672
R719 VTAIL.n271 VTAIL.n237 0.155672
R720 VTAIL.n271 VTAIL.n270 0.155672
R721 VTAIL.n270 VTAIL.n241 0.155672
R722 VTAIL.n263 VTAIL.n241 0.155672
R723 VTAIL.n263 VTAIL.n262 0.155672
R724 VTAIL.n262 VTAIL.n246 0.155672
R725 VTAIL.n255 VTAIL.n246 0.155672
R726 VTAIL.n255 VTAIL.n254 0.155672
R727 VTAIL.n229 VTAIL.n175 0.155672
R728 VTAIL.n222 VTAIL.n175 0.155672
R729 VTAIL.n222 VTAIL.n221 0.155672
R730 VTAIL.n221 VTAIL.n179 0.155672
R731 VTAIL.n213 VTAIL.n179 0.155672
R732 VTAIL.n213 VTAIL.n212 0.155672
R733 VTAIL.n212 VTAIL.n183 0.155672
R734 VTAIL.n205 VTAIL.n183 0.155672
R735 VTAIL.n205 VTAIL.n204 0.155672
R736 VTAIL.n204 VTAIL.n188 0.155672
R737 VTAIL.n197 VTAIL.n188 0.155672
R738 VTAIL.n197 VTAIL.n196 0.155672
R739 VDD1 VDD1.n1 119.394
R740 VDD1 VDD1.n0 74.9545
R741 VDD1.n0 VDD1.t1 3.05836
R742 VDD1.n0 VDD1.t2 3.05836
R743 VDD1.n1 VDD1.t0 3.05836
R744 VDD1.n1 VDD1.t3 3.05836
R745 B.n525 B.n524 585
R746 B.n526 B.n71 585
R747 B.n528 B.n527 585
R748 B.n529 B.n70 585
R749 B.n531 B.n530 585
R750 B.n532 B.n69 585
R751 B.n534 B.n533 585
R752 B.n535 B.n68 585
R753 B.n537 B.n536 585
R754 B.n538 B.n67 585
R755 B.n540 B.n539 585
R756 B.n541 B.n66 585
R757 B.n543 B.n542 585
R758 B.n544 B.n65 585
R759 B.n546 B.n545 585
R760 B.n547 B.n64 585
R761 B.n549 B.n548 585
R762 B.n550 B.n63 585
R763 B.n552 B.n551 585
R764 B.n553 B.n62 585
R765 B.n555 B.n554 585
R766 B.n556 B.n61 585
R767 B.n558 B.n557 585
R768 B.n559 B.n60 585
R769 B.n561 B.n560 585
R770 B.n562 B.n59 585
R771 B.n564 B.n563 585
R772 B.n565 B.n58 585
R773 B.n567 B.n566 585
R774 B.n568 B.n57 585
R775 B.n570 B.n569 585
R776 B.n571 B.n56 585
R777 B.n573 B.n572 585
R778 B.n574 B.n55 585
R779 B.n576 B.n575 585
R780 B.n577 B.n54 585
R781 B.n579 B.n578 585
R782 B.n580 B.n51 585
R783 B.n583 B.n582 585
R784 B.n584 B.n50 585
R785 B.n586 B.n585 585
R786 B.n587 B.n49 585
R787 B.n589 B.n588 585
R788 B.n590 B.n48 585
R789 B.n592 B.n591 585
R790 B.n593 B.n47 585
R791 B.n595 B.n594 585
R792 B.n597 B.n596 585
R793 B.n598 B.n43 585
R794 B.n600 B.n599 585
R795 B.n601 B.n42 585
R796 B.n603 B.n602 585
R797 B.n604 B.n41 585
R798 B.n606 B.n605 585
R799 B.n607 B.n40 585
R800 B.n609 B.n608 585
R801 B.n610 B.n39 585
R802 B.n612 B.n611 585
R803 B.n613 B.n38 585
R804 B.n615 B.n614 585
R805 B.n616 B.n37 585
R806 B.n618 B.n617 585
R807 B.n619 B.n36 585
R808 B.n621 B.n620 585
R809 B.n622 B.n35 585
R810 B.n624 B.n623 585
R811 B.n625 B.n34 585
R812 B.n627 B.n626 585
R813 B.n628 B.n33 585
R814 B.n630 B.n629 585
R815 B.n631 B.n32 585
R816 B.n633 B.n632 585
R817 B.n634 B.n31 585
R818 B.n636 B.n635 585
R819 B.n637 B.n30 585
R820 B.n639 B.n638 585
R821 B.n640 B.n29 585
R822 B.n642 B.n641 585
R823 B.n643 B.n28 585
R824 B.n645 B.n644 585
R825 B.n646 B.n27 585
R826 B.n648 B.n647 585
R827 B.n649 B.n26 585
R828 B.n651 B.n650 585
R829 B.n652 B.n25 585
R830 B.n523 B.n72 585
R831 B.n522 B.n521 585
R832 B.n520 B.n73 585
R833 B.n519 B.n518 585
R834 B.n517 B.n74 585
R835 B.n516 B.n515 585
R836 B.n514 B.n75 585
R837 B.n513 B.n512 585
R838 B.n511 B.n76 585
R839 B.n510 B.n509 585
R840 B.n508 B.n77 585
R841 B.n507 B.n506 585
R842 B.n505 B.n78 585
R843 B.n504 B.n503 585
R844 B.n502 B.n79 585
R845 B.n501 B.n500 585
R846 B.n499 B.n80 585
R847 B.n498 B.n497 585
R848 B.n496 B.n81 585
R849 B.n495 B.n494 585
R850 B.n493 B.n82 585
R851 B.n492 B.n491 585
R852 B.n490 B.n83 585
R853 B.n489 B.n488 585
R854 B.n487 B.n84 585
R855 B.n486 B.n485 585
R856 B.n484 B.n85 585
R857 B.n483 B.n482 585
R858 B.n481 B.n86 585
R859 B.n480 B.n479 585
R860 B.n478 B.n87 585
R861 B.n477 B.n476 585
R862 B.n475 B.n88 585
R863 B.n474 B.n473 585
R864 B.n472 B.n89 585
R865 B.n471 B.n470 585
R866 B.n469 B.n90 585
R867 B.n468 B.n467 585
R868 B.n466 B.n91 585
R869 B.n465 B.n464 585
R870 B.n463 B.n92 585
R871 B.n462 B.n461 585
R872 B.n460 B.n93 585
R873 B.n459 B.n458 585
R874 B.n457 B.n94 585
R875 B.n456 B.n455 585
R876 B.n454 B.n95 585
R877 B.n453 B.n452 585
R878 B.n451 B.n96 585
R879 B.n450 B.n449 585
R880 B.n448 B.n97 585
R881 B.n447 B.n446 585
R882 B.n445 B.n98 585
R883 B.n444 B.n443 585
R884 B.n442 B.n99 585
R885 B.n441 B.n440 585
R886 B.n439 B.n100 585
R887 B.n438 B.n437 585
R888 B.n436 B.n101 585
R889 B.n435 B.n434 585
R890 B.n433 B.n102 585
R891 B.n432 B.n431 585
R892 B.n430 B.n103 585
R893 B.n429 B.n428 585
R894 B.n427 B.n104 585
R895 B.n426 B.n425 585
R896 B.n424 B.n105 585
R897 B.n423 B.n422 585
R898 B.n421 B.n106 585
R899 B.n420 B.n419 585
R900 B.n418 B.n107 585
R901 B.n417 B.n416 585
R902 B.n415 B.n108 585
R903 B.n414 B.n413 585
R904 B.n412 B.n109 585
R905 B.n411 B.n410 585
R906 B.n409 B.n110 585
R907 B.n408 B.n407 585
R908 B.n406 B.n111 585
R909 B.n405 B.n404 585
R910 B.n403 B.n112 585
R911 B.n402 B.n401 585
R912 B.n400 B.n113 585
R913 B.n399 B.n398 585
R914 B.n397 B.n114 585
R915 B.n396 B.n395 585
R916 B.n394 B.n115 585
R917 B.n393 B.n392 585
R918 B.n391 B.n116 585
R919 B.n390 B.n389 585
R920 B.n388 B.n117 585
R921 B.n387 B.n386 585
R922 B.n385 B.n118 585
R923 B.n256 B.n165 585
R924 B.n258 B.n257 585
R925 B.n259 B.n164 585
R926 B.n261 B.n260 585
R927 B.n262 B.n163 585
R928 B.n264 B.n263 585
R929 B.n265 B.n162 585
R930 B.n267 B.n266 585
R931 B.n268 B.n161 585
R932 B.n270 B.n269 585
R933 B.n271 B.n160 585
R934 B.n273 B.n272 585
R935 B.n274 B.n159 585
R936 B.n276 B.n275 585
R937 B.n277 B.n158 585
R938 B.n279 B.n278 585
R939 B.n280 B.n157 585
R940 B.n282 B.n281 585
R941 B.n283 B.n156 585
R942 B.n285 B.n284 585
R943 B.n286 B.n155 585
R944 B.n288 B.n287 585
R945 B.n289 B.n154 585
R946 B.n291 B.n290 585
R947 B.n292 B.n153 585
R948 B.n294 B.n293 585
R949 B.n295 B.n152 585
R950 B.n297 B.n296 585
R951 B.n298 B.n151 585
R952 B.n300 B.n299 585
R953 B.n301 B.n150 585
R954 B.n303 B.n302 585
R955 B.n304 B.n149 585
R956 B.n306 B.n305 585
R957 B.n307 B.n148 585
R958 B.n309 B.n308 585
R959 B.n310 B.n147 585
R960 B.n312 B.n311 585
R961 B.n314 B.n313 585
R962 B.n315 B.n143 585
R963 B.n317 B.n316 585
R964 B.n318 B.n142 585
R965 B.n320 B.n319 585
R966 B.n321 B.n141 585
R967 B.n323 B.n322 585
R968 B.n324 B.n140 585
R969 B.n326 B.n325 585
R970 B.n328 B.n137 585
R971 B.n330 B.n329 585
R972 B.n331 B.n136 585
R973 B.n333 B.n332 585
R974 B.n334 B.n135 585
R975 B.n336 B.n335 585
R976 B.n337 B.n134 585
R977 B.n339 B.n338 585
R978 B.n340 B.n133 585
R979 B.n342 B.n341 585
R980 B.n343 B.n132 585
R981 B.n345 B.n344 585
R982 B.n346 B.n131 585
R983 B.n348 B.n347 585
R984 B.n349 B.n130 585
R985 B.n351 B.n350 585
R986 B.n352 B.n129 585
R987 B.n354 B.n353 585
R988 B.n355 B.n128 585
R989 B.n357 B.n356 585
R990 B.n358 B.n127 585
R991 B.n360 B.n359 585
R992 B.n361 B.n126 585
R993 B.n363 B.n362 585
R994 B.n364 B.n125 585
R995 B.n366 B.n365 585
R996 B.n367 B.n124 585
R997 B.n369 B.n368 585
R998 B.n370 B.n123 585
R999 B.n372 B.n371 585
R1000 B.n373 B.n122 585
R1001 B.n375 B.n374 585
R1002 B.n376 B.n121 585
R1003 B.n378 B.n377 585
R1004 B.n379 B.n120 585
R1005 B.n381 B.n380 585
R1006 B.n382 B.n119 585
R1007 B.n384 B.n383 585
R1008 B.n255 B.n254 585
R1009 B.n253 B.n166 585
R1010 B.n252 B.n251 585
R1011 B.n250 B.n167 585
R1012 B.n249 B.n248 585
R1013 B.n247 B.n168 585
R1014 B.n246 B.n245 585
R1015 B.n244 B.n169 585
R1016 B.n243 B.n242 585
R1017 B.n241 B.n170 585
R1018 B.n240 B.n239 585
R1019 B.n238 B.n171 585
R1020 B.n237 B.n236 585
R1021 B.n235 B.n172 585
R1022 B.n234 B.n233 585
R1023 B.n232 B.n173 585
R1024 B.n231 B.n230 585
R1025 B.n229 B.n174 585
R1026 B.n228 B.n227 585
R1027 B.n226 B.n175 585
R1028 B.n225 B.n224 585
R1029 B.n223 B.n176 585
R1030 B.n222 B.n221 585
R1031 B.n220 B.n177 585
R1032 B.n219 B.n218 585
R1033 B.n217 B.n178 585
R1034 B.n216 B.n215 585
R1035 B.n214 B.n179 585
R1036 B.n213 B.n212 585
R1037 B.n211 B.n180 585
R1038 B.n210 B.n209 585
R1039 B.n208 B.n181 585
R1040 B.n207 B.n206 585
R1041 B.n205 B.n182 585
R1042 B.n204 B.n203 585
R1043 B.n202 B.n183 585
R1044 B.n201 B.n200 585
R1045 B.n199 B.n184 585
R1046 B.n198 B.n197 585
R1047 B.n196 B.n185 585
R1048 B.n195 B.n194 585
R1049 B.n193 B.n186 585
R1050 B.n192 B.n191 585
R1051 B.n190 B.n187 585
R1052 B.n189 B.n188 585
R1053 B.n2 B.n0 585
R1054 B.n721 B.n1 585
R1055 B.n720 B.n719 585
R1056 B.n718 B.n3 585
R1057 B.n717 B.n716 585
R1058 B.n715 B.n4 585
R1059 B.n714 B.n713 585
R1060 B.n712 B.n5 585
R1061 B.n711 B.n710 585
R1062 B.n709 B.n6 585
R1063 B.n708 B.n707 585
R1064 B.n706 B.n7 585
R1065 B.n705 B.n704 585
R1066 B.n703 B.n8 585
R1067 B.n702 B.n701 585
R1068 B.n700 B.n9 585
R1069 B.n699 B.n698 585
R1070 B.n697 B.n10 585
R1071 B.n696 B.n695 585
R1072 B.n694 B.n11 585
R1073 B.n693 B.n692 585
R1074 B.n691 B.n12 585
R1075 B.n690 B.n689 585
R1076 B.n688 B.n13 585
R1077 B.n687 B.n686 585
R1078 B.n685 B.n14 585
R1079 B.n684 B.n683 585
R1080 B.n682 B.n15 585
R1081 B.n681 B.n680 585
R1082 B.n679 B.n16 585
R1083 B.n678 B.n677 585
R1084 B.n676 B.n17 585
R1085 B.n675 B.n674 585
R1086 B.n673 B.n18 585
R1087 B.n672 B.n671 585
R1088 B.n670 B.n19 585
R1089 B.n669 B.n668 585
R1090 B.n667 B.n20 585
R1091 B.n666 B.n665 585
R1092 B.n664 B.n21 585
R1093 B.n663 B.n662 585
R1094 B.n661 B.n22 585
R1095 B.n660 B.n659 585
R1096 B.n658 B.n23 585
R1097 B.n657 B.n656 585
R1098 B.n655 B.n24 585
R1099 B.n654 B.n653 585
R1100 B.n723 B.n722 585
R1101 B.n254 B.n165 473.281
R1102 B.n654 B.n25 473.281
R1103 B.n385 B.n384 473.281
R1104 B.n524 B.n523 473.281
R1105 B.n138 B.t11 434.046
R1106 B.n52 B.t4 434.046
R1107 B.n144 B.t2 434.046
R1108 B.n44 B.t7 434.046
R1109 B.n139 B.t10 350.846
R1110 B.n53 B.t5 350.846
R1111 B.n145 B.t1 350.846
R1112 B.n45 B.t8 350.846
R1113 B.n138 B.t9 274.156
R1114 B.n144 B.t0 274.156
R1115 B.n44 B.t6 274.156
R1116 B.n52 B.t3 274.156
R1117 B.n254 B.n253 163.367
R1118 B.n253 B.n252 163.367
R1119 B.n252 B.n167 163.367
R1120 B.n248 B.n167 163.367
R1121 B.n248 B.n247 163.367
R1122 B.n247 B.n246 163.367
R1123 B.n246 B.n169 163.367
R1124 B.n242 B.n169 163.367
R1125 B.n242 B.n241 163.367
R1126 B.n241 B.n240 163.367
R1127 B.n240 B.n171 163.367
R1128 B.n236 B.n171 163.367
R1129 B.n236 B.n235 163.367
R1130 B.n235 B.n234 163.367
R1131 B.n234 B.n173 163.367
R1132 B.n230 B.n173 163.367
R1133 B.n230 B.n229 163.367
R1134 B.n229 B.n228 163.367
R1135 B.n228 B.n175 163.367
R1136 B.n224 B.n175 163.367
R1137 B.n224 B.n223 163.367
R1138 B.n223 B.n222 163.367
R1139 B.n222 B.n177 163.367
R1140 B.n218 B.n177 163.367
R1141 B.n218 B.n217 163.367
R1142 B.n217 B.n216 163.367
R1143 B.n216 B.n179 163.367
R1144 B.n212 B.n179 163.367
R1145 B.n212 B.n211 163.367
R1146 B.n211 B.n210 163.367
R1147 B.n210 B.n181 163.367
R1148 B.n206 B.n181 163.367
R1149 B.n206 B.n205 163.367
R1150 B.n205 B.n204 163.367
R1151 B.n204 B.n183 163.367
R1152 B.n200 B.n183 163.367
R1153 B.n200 B.n199 163.367
R1154 B.n199 B.n198 163.367
R1155 B.n198 B.n185 163.367
R1156 B.n194 B.n185 163.367
R1157 B.n194 B.n193 163.367
R1158 B.n193 B.n192 163.367
R1159 B.n192 B.n187 163.367
R1160 B.n188 B.n187 163.367
R1161 B.n188 B.n2 163.367
R1162 B.n722 B.n2 163.367
R1163 B.n722 B.n721 163.367
R1164 B.n721 B.n720 163.367
R1165 B.n720 B.n3 163.367
R1166 B.n716 B.n3 163.367
R1167 B.n716 B.n715 163.367
R1168 B.n715 B.n714 163.367
R1169 B.n714 B.n5 163.367
R1170 B.n710 B.n5 163.367
R1171 B.n710 B.n709 163.367
R1172 B.n709 B.n708 163.367
R1173 B.n708 B.n7 163.367
R1174 B.n704 B.n7 163.367
R1175 B.n704 B.n703 163.367
R1176 B.n703 B.n702 163.367
R1177 B.n702 B.n9 163.367
R1178 B.n698 B.n9 163.367
R1179 B.n698 B.n697 163.367
R1180 B.n697 B.n696 163.367
R1181 B.n696 B.n11 163.367
R1182 B.n692 B.n11 163.367
R1183 B.n692 B.n691 163.367
R1184 B.n691 B.n690 163.367
R1185 B.n690 B.n13 163.367
R1186 B.n686 B.n13 163.367
R1187 B.n686 B.n685 163.367
R1188 B.n685 B.n684 163.367
R1189 B.n684 B.n15 163.367
R1190 B.n680 B.n15 163.367
R1191 B.n680 B.n679 163.367
R1192 B.n679 B.n678 163.367
R1193 B.n678 B.n17 163.367
R1194 B.n674 B.n17 163.367
R1195 B.n674 B.n673 163.367
R1196 B.n673 B.n672 163.367
R1197 B.n672 B.n19 163.367
R1198 B.n668 B.n19 163.367
R1199 B.n668 B.n667 163.367
R1200 B.n667 B.n666 163.367
R1201 B.n666 B.n21 163.367
R1202 B.n662 B.n21 163.367
R1203 B.n662 B.n661 163.367
R1204 B.n661 B.n660 163.367
R1205 B.n660 B.n23 163.367
R1206 B.n656 B.n23 163.367
R1207 B.n656 B.n655 163.367
R1208 B.n655 B.n654 163.367
R1209 B.n258 B.n165 163.367
R1210 B.n259 B.n258 163.367
R1211 B.n260 B.n259 163.367
R1212 B.n260 B.n163 163.367
R1213 B.n264 B.n163 163.367
R1214 B.n265 B.n264 163.367
R1215 B.n266 B.n265 163.367
R1216 B.n266 B.n161 163.367
R1217 B.n270 B.n161 163.367
R1218 B.n271 B.n270 163.367
R1219 B.n272 B.n271 163.367
R1220 B.n272 B.n159 163.367
R1221 B.n276 B.n159 163.367
R1222 B.n277 B.n276 163.367
R1223 B.n278 B.n277 163.367
R1224 B.n278 B.n157 163.367
R1225 B.n282 B.n157 163.367
R1226 B.n283 B.n282 163.367
R1227 B.n284 B.n283 163.367
R1228 B.n284 B.n155 163.367
R1229 B.n288 B.n155 163.367
R1230 B.n289 B.n288 163.367
R1231 B.n290 B.n289 163.367
R1232 B.n290 B.n153 163.367
R1233 B.n294 B.n153 163.367
R1234 B.n295 B.n294 163.367
R1235 B.n296 B.n295 163.367
R1236 B.n296 B.n151 163.367
R1237 B.n300 B.n151 163.367
R1238 B.n301 B.n300 163.367
R1239 B.n302 B.n301 163.367
R1240 B.n302 B.n149 163.367
R1241 B.n306 B.n149 163.367
R1242 B.n307 B.n306 163.367
R1243 B.n308 B.n307 163.367
R1244 B.n308 B.n147 163.367
R1245 B.n312 B.n147 163.367
R1246 B.n313 B.n312 163.367
R1247 B.n313 B.n143 163.367
R1248 B.n317 B.n143 163.367
R1249 B.n318 B.n317 163.367
R1250 B.n319 B.n318 163.367
R1251 B.n319 B.n141 163.367
R1252 B.n323 B.n141 163.367
R1253 B.n324 B.n323 163.367
R1254 B.n325 B.n324 163.367
R1255 B.n325 B.n137 163.367
R1256 B.n330 B.n137 163.367
R1257 B.n331 B.n330 163.367
R1258 B.n332 B.n331 163.367
R1259 B.n332 B.n135 163.367
R1260 B.n336 B.n135 163.367
R1261 B.n337 B.n336 163.367
R1262 B.n338 B.n337 163.367
R1263 B.n338 B.n133 163.367
R1264 B.n342 B.n133 163.367
R1265 B.n343 B.n342 163.367
R1266 B.n344 B.n343 163.367
R1267 B.n344 B.n131 163.367
R1268 B.n348 B.n131 163.367
R1269 B.n349 B.n348 163.367
R1270 B.n350 B.n349 163.367
R1271 B.n350 B.n129 163.367
R1272 B.n354 B.n129 163.367
R1273 B.n355 B.n354 163.367
R1274 B.n356 B.n355 163.367
R1275 B.n356 B.n127 163.367
R1276 B.n360 B.n127 163.367
R1277 B.n361 B.n360 163.367
R1278 B.n362 B.n361 163.367
R1279 B.n362 B.n125 163.367
R1280 B.n366 B.n125 163.367
R1281 B.n367 B.n366 163.367
R1282 B.n368 B.n367 163.367
R1283 B.n368 B.n123 163.367
R1284 B.n372 B.n123 163.367
R1285 B.n373 B.n372 163.367
R1286 B.n374 B.n373 163.367
R1287 B.n374 B.n121 163.367
R1288 B.n378 B.n121 163.367
R1289 B.n379 B.n378 163.367
R1290 B.n380 B.n379 163.367
R1291 B.n380 B.n119 163.367
R1292 B.n384 B.n119 163.367
R1293 B.n386 B.n385 163.367
R1294 B.n386 B.n117 163.367
R1295 B.n390 B.n117 163.367
R1296 B.n391 B.n390 163.367
R1297 B.n392 B.n391 163.367
R1298 B.n392 B.n115 163.367
R1299 B.n396 B.n115 163.367
R1300 B.n397 B.n396 163.367
R1301 B.n398 B.n397 163.367
R1302 B.n398 B.n113 163.367
R1303 B.n402 B.n113 163.367
R1304 B.n403 B.n402 163.367
R1305 B.n404 B.n403 163.367
R1306 B.n404 B.n111 163.367
R1307 B.n408 B.n111 163.367
R1308 B.n409 B.n408 163.367
R1309 B.n410 B.n409 163.367
R1310 B.n410 B.n109 163.367
R1311 B.n414 B.n109 163.367
R1312 B.n415 B.n414 163.367
R1313 B.n416 B.n415 163.367
R1314 B.n416 B.n107 163.367
R1315 B.n420 B.n107 163.367
R1316 B.n421 B.n420 163.367
R1317 B.n422 B.n421 163.367
R1318 B.n422 B.n105 163.367
R1319 B.n426 B.n105 163.367
R1320 B.n427 B.n426 163.367
R1321 B.n428 B.n427 163.367
R1322 B.n428 B.n103 163.367
R1323 B.n432 B.n103 163.367
R1324 B.n433 B.n432 163.367
R1325 B.n434 B.n433 163.367
R1326 B.n434 B.n101 163.367
R1327 B.n438 B.n101 163.367
R1328 B.n439 B.n438 163.367
R1329 B.n440 B.n439 163.367
R1330 B.n440 B.n99 163.367
R1331 B.n444 B.n99 163.367
R1332 B.n445 B.n444 163.367
R1333 B.n446 B.n445 163.367
R1334 B.n446 B.n97 163.367
R1335 B.n450 B.n97 163.367
R1336 B.n451 B.n450 163.367
R1337 B.n452 B.n451 163.367
R1338 B.n452 B.n95 163.367
R1339 B.n456 B.n95 163.367
R1340 B.n457 B.n456 163.367
R1341 B.n458 B.n457 163.367
R1342 B.n458 B.n93 163.367
R1343 B.n462 B.n93 163.367
R1344 B.n463 B.n462 163.367
R1345 B.n464 B.n463 163.367
R1346 B.n464 B.n91 163.367
R1347 B.n468 B.n91 163.367
R1348 B.n469 B.n468 163.367
R1349 B.n470 B.n469 163.367
R1350 B.n470 B.n89 163.367
R1351 B.n474 B.n89 163.367
R1352 B.n475 B.n474 163.367
R1353 B.n476 B.n475 163.367
R1354 B.n476 B.n87 163.367
R1355 B.n480 B.n87 163.367
R1356 B.n481 B.n480 163.367
R1357 B.n482 B.n481 163.367
R1358 B.n482 B.n85 163.367
R1359 B.n486 B.n85 163.367
R1360 B.n487 B.n486 163.367
R1361 B.n488 B.n487 163.367
R1362 B.n488 B.n83 163.367
R1363 B.n492 B.n83 163.367
R1364 B.n493 B.n492 163.367
R1365 B.n494 B.n493 163.367
R1366 B.n494 B.n81 163.367
R1367 B.n498 B.n81 163.367
R1368 B.n499 B.n498 163.367
R1369 B.n500 B.n499 163.367
R1370 B.n500 B.n79 163.367
R1371 B.n504 B.n79 163.367
R1372 B.n505 B.n504 163.367
R1373 B.n506 B.n505 163.367
R1374 B.n506 B.n77 163.367
R1375 B.n510 B.n77 163.367
R1376 B.n511 B.n510 163.367
R1377 B.n512 B.n511 163.367
R1378 B.n512 B.n75 163.367
R1379 B.n516 B.n75 163.367
R1380 B.n517 B.n516 163.367
R1381 B.n518 B.n517 163.367
R1382 B.n518 B.n73 163.367
R1383 B.n522 B.n73 163.367
R1384 B.n523 B.n522 163.367
R1385 B.n650 B.n25 163.367
R1386 B.n650 B.n649 163.367
R1387 B.n649 B.n648 163.367
R1388 B.n648 B.n27 163.367
R1389 B.n644 B.n27 163.367
R1390 B.n644 B.n643 163.367
R1391 B.n643 B.n642 163.367
R1392 B.n642 B.n29 163.367
R1393 B.n638 B.n29 163.367
R1394 B.n638 B.n637 163.367
R1395 B.n637 B.n636 163.367
R1396 B.n636 B.n31 163.367
R1397 B.n632 B.n31 163.367
R1398 B.n632 B.n631 163.367
R1399 B.n631 B.n630 163.367
R1400 B.n630 B.n33 163.367
R1401 B.n626 B.n33 163.367
R1402 B.n626 B.n625 163.367
R1403 B.n625 B.n624 163.367
R1404 B.n624 B.n35 163.367
R1405 B.n620 B.n35 163.367
R1406 B.n620 B.n619 163.367
R1407 B.n619 B.n618 163.367
R1408 B.n618 B.n37 163.367
R1409 B.n614 B.n37 163.367
R1410 B.n614 B.n613 163.367
R1411 B.n613 B.n612 163.367
R1412 B.n612 B.n39 163.367
R1413 B.n608 B.n39 163.367
R1414 B.n608 B.n607 163.367
R1415 B.n607 B.n606 163.367
R1416 B.n606 B.n41 163.367
R1417 B.n602 B.n41 163.367
R1418 B.n602 B.n601 163.367
R1419 B.n601 B.n600 163.367
R1420 B.n600 B.n43 163.367
R1421 B.n596 B.n43 163.367
R1422 B.n596 B.n595 163.367
R1423 B.n595 B.n47 163.367
R1424 B.n591 B.n47 163.367
R1425 B.n591 B.n590 163.367
R1426 B.n590 B.n589 163.367
R1427 B.n589 B.n49 163.367
R1428 B.n585 B.n49 163.367
R1429 B.n585 B.n584 163.367
R1430 B.n584 B.n583 163.367
R1431 B.n583 B.n51 163.367
R1432 B.n578 B.n51 163.367
R1433 B.n578 B.n577 163.367
R1434 B.n577 B.n576 163.367
R1435 B.n576 B.n55 163.367
R1436 B.n572 B.n55 163.367
R1437 B.n572 B.n571 163.367
R1438 B.n571 B.n570 163.367
R1439 B.n570 B.n57 163.367
R1440 B.n566 B.n57 163.367
R1441 B.n566 B.n565 163.367
R1442 B.n565 B.n564 163.367
R1443 B.n564 B.n59 163.367
R1444 B.n560 B.n59 163.367
R1445 B.n560 B.n559 163.367
R1446 B.n559 B.n558 163.367
R1447 B.n558 B.n61 163.367
R1448 B.n554 B.n61 163.367
R1449 B.n554 B.n553 163.367
R1450 B.n553 B.n552 163.367
R1451 B.n552 B.n63 163.367
R1452 B.n548 B.n63 163.367
R1453 B.n548 B.n547 163.367
R1454 B.n547 B.n546 163.367
R1455 B.n546 B.n65 163.367
R1456 B.n542 B.n65 163.367
R1457 B.n542 B.n541 163.367
R1458 B.n541 B.n540 163.367
R1459 B.n540 B.n67 163.367
R1460 B.n536 B.n67 163.367
R1461 B.n536 B.n535 163.367
R1462 B.n535 B.n534 163.367
R1463 B.n534 B.n69 163.367
R1464 B.n530 B.n69 163.367
R1465 B.n530 B.n529 163.367
R1466 B.n529 B.n528 163.367
R1467 B.n528 B.n71 163.367
R1468 B.n524 B.n71 163.367
R1469 B.n139 B.n138 83.2005
R1470 B.n145 B.n144 83.2005
R1471 B.n45 B.n44 83.2005
R1472 B.n53 B.n52 83.2005
R1473 B.n327 B.n139 59.5399
R1474 B.n146 B.n145 59.5399
R1475 B.n46 B.n45 59.5399
R1476 B.n581 B.n53 59.5399
R1477 B.n653 B.n652 30.7517
R1478 B.n525 B.n72 30.7517
R1479 B.n383 B.n118 30.7517
R1480 B.n256 B.n255 30.7517
R1481 B B.n723 18.0485
R1482 B.n652 B.n651 10.6151
R1483 B.n651 B.n26 10.6151
R1484 B.n647 B.n26 10.6151
R1485 B.n647 B.n646 10.6151
R1486 B.n646 B.n645 10.6151
R1487 B.n645 B.n28 10.6151
R1488 B.n641 B.n28 10.6151
R1489 B.n641 B.n640 10.6151
R1490 B.n640 B.n639 10.6151
R1491 B.n639 B.n30 10.6151
R1492 B.n635 B.n30 10.6151
R1493 B.n635 B.n634 10.6151
R1494 B.n634 B.n633 10.6151
R1495 B.n633 B.n32 10.6151
R1496 B.n629 B.n32 10.6151
R1497 B.n629 B.n628 10.6151
R1498 B.n628 B.n627 10.6151
R1499 B.n627 B.n34 10.6151
R1500 B.n623 B.n34 10.6151
R1501 B.n623 B.n622 10.6151
R1502 B.n622 B.n621 10.6151
R1503 B.n621 B.n36 10.6151
R1504 B.n617 B.n36 10.6151
R1505 B.n617 B.n616 10.6151
R1506 B.n616 B.n615 10.6151
R1507 B.n615 B.n38 10.6151
R1508 B.n611 B.n38 10.6151
R1509 B.n611 B.n610 10.6151
R1510 B.n610 B.n609 10.6151
R1511 B.n609 B.n40 10.6151
R1512 B.n605 B.n40 10.6151
R1513 B.n605 B.n604 10.6151
R1514 B.n604 B.n603 10.6151
R1515 B.n603 B.n42 10.6151
R1516 B.n599 B.n42 10.6151
R1517 B.n599 B.n598 10.6151
R1518 B.n598 B.n597 10.6151
R1519 B.n594 B.n593 10.6151
R1520 B.n593 B.n592 10.6151
R1521 B.n592 B.n48 10.6151
R1522 B.n588 B.n48 10.6151
R1523 B.n588 B.n587 10.6151
R1524 B.n587 B.n586 10.6151
R1525 B.n586 B.n50 10.6151
R1526 B.n582 B.n50 10.6151
R1527 B.n580 B.n579 10.6151
R1528 B.n579 B.n54 10.6151
R1529 B.n575 B.n54 10.6151
R1530 B.n575 B.n574 10.6151
R1531 B.n574 B.n573 10.6151
R1532 B.n573 B.n56 10.6151
R1533 B.n569 B.n56 10.6151
R1534 B.n569 B.n568 10.6151
R1535 B.n568 B.n567 10.6151
R1536 B.n567 B.n58 10.6151
R1537 B.n563 B.n58 10.6151
R1538 B.n563 B.n562 10.6151
R1539 B.n562 B.n561 10.6151
R1540 B.n561 B.n60 10.6151
R1541 B.n557 B.n60 10.6151
R1542 B.n557 B.n556 10.6151
R1543 B.n556 B.n555 10.6151
R1544 B.n555 B.n62 10.6151
R1545 B.n551 B.n62 10.6151
R1546 B.n551 B.n550 10.6151
R1547 B.n550 B.n549 10.6151
R1548 B.n549 B.n64 10.6151
R1549 B.n545 B.n64 10.6151
R1550 B.n545 B.n544 10.6151
R1551 B.n544 B.n543 10.6151
R1552 B.n543 B.n66 10.6151
R1553 B.n539 B.n66 10.6151
R1554 B.n539 B.n538 10.6151
R1555 B.n538 B.n537 10.6151
R1556 B.n537 B.n68 10.6151
R1557 B.n533 B.n68 10.6151
R1558 B.n533 B.n532 10.6151
R1559 B.n532 B.n531 10.6151
R1560 B.n531 B.n70 10.6151
R1561 B.n527 B.n70 10.6151
R1562 B.n527 B.n526 10.6151
R1563 B.n526 B.n525 10.6151
R1564 B.n387 B.n118 10.6151
R1565 B.n388 B.n387 10.6151
R1566 B.n389 B.n388 10.6151
R1567 B.n389 B.n116 10.6151
R1568 B.n393 B.n116 10.6151
R1569 B.n394 B.n393 10.6151
R1570 B.n395 B.n394 10.6151
R1571 B.n395 B.n114 10.6151
R1572 B.n399 B.n114 10.6151
R1573 B.n400 B.n399 10.6151
R1574 B.n401 B.n400 10.6151
R1575 B.n401 B.n112 10.6151
R1576 B.n405 B.n112 10.6151
R1577 B.n406 B.n405 10.6151
R1578 B.n407 B.n406 10.6151
R1579 B.n407 B.n110 10.6151
R1580 B.n411 B.n110 10.6151
R1581 B.n412 B.n411 10.6151
R1582 B.n413 B.n412 10.6151
R1583 B.n413 B.n108 10.6151
R1584 B.n417 B.n108 10.6151
R1585 B.n418 B.n417 10.6151
R1586 B.n419 B.n418 10.6151
R1587 B.n419 B.n106 10.6151
R1588 B.n423 B.n106 10.6151
R1589 B.n424 B.n423 10.6151
R1590 B.n425 B.n424 10.6151
R1591 B.n425 B.n104 10.6151
R1592 B.n429 B.n104 10.6151
R1593 B.n430 B.n429 10.6151
R1594 B.n431 B.n430 10.6151
R1595 B.n431 B.n102 10.6151
R1596 B.n435 B.n102 10.6151
R1597 B.n436 B.n435 10.6151
R1598 B.n437 B.n436 10.6151
R1599 B.n437 B.n100 10.6151
R1600 B.n441 B.n100 10.6151
R1601 B.n442 B.n441 10.6151
R1602 B.n443 B.n442 10.6151
R1603 B.n443 B.n98 10.6151
R1604 B.n447 B.n98 10.6151
R1605 B.n448 B.n447 10.6151
R1606 B.n449 B.n448 10.6151
R1607 B.n449 B.n96 10.6151
R1608 B.n453 B.n96 10.6151
R1609 B.n454 B.n453 10.6151
R1610 B.n455 B.n454 10.6151
R1611 B.n455 B.n94 10.6151
R1612 B.n459 B.n94 10.6151
R1613 B.n460 B.n459 10.6151
R1614 B.n461 B.n460 10.6151
R1615 B.n461 B.n92 10.6151
R1616 B.n465 B.n92 10.6151
R1617 B.n466 B.n465 10.6151
R1618 B.n467 B.n466 10.6151
R1619 B.n467 B.n90 10.6151
R1620 B.n471 B.n90 10.6151
R1621 B.n472 B.n471 10.6151
R1622 B.n473 B.n472 10.6151
R1623 B.n473 B.n88 10.6151
R1624 B.n477 B.n88 10.6151
R1625 B.n478 B.n477 10.6151
R1626 B.n479 B.n478 10.6151
R1627 B.n479 B.n86 10.6151
R1628 B.n483 B.n86 10.6151
R1629 B.n484 B.n483 10.6151
R1630 B.n485 B.n484 10.6151
R1631 B.n485 B.n84 10.6151
R1632 B.n489 B.n84 10.6151
R1633 B.n490 B.n489 10.6151
R1634 B.n491 B.n490 10.6151
R1635 B.n491 B.n82 10.6151
R1636 B.n495 B.n82 10.6151
R1637 B.n496 B.n495 10.6151
R1638 B.n497 B.n496 10.6151
R1639 B.n497 B.n80 10.6151
R1640 B.n501 B.n80 10.6151
R1641 B.n502 B.n501 10.6151
R1642 B.n503 B.n502 10.6151
R1643 B.n503 B.n78 10.6151
R1644 B.n507 B.n78 10.6151
R1645 B.n508 B.n507 10.6151
R1646 B.n509 B.n508 10.6151
R1647 B.n509 B.n76 10.6151
R1648 B.n513 B.n76 10.6151
R1649 B.n514 B.n513 10.6151
R1650 B.n515 B.n514 10.6151
R1651 B.n515 B.n74 10.6151
R1652 B.n519 B.n74 10.6151
R1653 B.n520 B.n519 10.6151
R1654 B.n521 B.n520 10.6151
R1655 B.n521 B.n72 10.6151
R1656 B.n257 B.n256 10.6151
R1657 B.n257 B.n164 10.6151
R1658 B.n261 B.n164 10.6151
R1659 B.n262 B.n261 10.6151
R1660 B.n263 B.n262 10.6151
R1661 B.n263 B.n162 10.6151
R1662 B.n267 B.n162 10.6151
R1663 B.n268 B.n267 10.6151
R1664 B.n269 B.n268 10.6151
R1665 B.n269 B.n160 10.6151
R1666 B.n273 B.n160 10.6151
R1667 B.n274 B.n273 10.6151
R1668 B.n275 B.n274 10.6151
R1669 B.n275 B.n158 10.6151
R1670 B.n279 B.n158 10.6151
R1671 B.n280 B.n279 10.6151
R1672 B.n281 B.n280 10.6151
R1673 B.n281 B.n156 10.6151
R1674 B.n285 B.n156 10.6151
R1675 B.n286 B.n285 10.6151
R1676 B.n287 B.n286 10.6151
R1677 B.n287 B.n154 10.6151
R1678 B.n291 B.n154 10.6151
R1679 B.n292 B.n291 10.6151
R1680 B.n293 B.n292 10.6151
R1681 B.n293 B.n152 10.6151
R1682 B.n297 B.n152 10.6151
R1683 B.n298 B.n297 10.6151
R1684 B.n299 B.n298 10.6151
R1685 B.n299 B.n150 10.6151
R1686 B.n303 B.n150 10.6151
R1687 B.n304 B.n303 10.6151
R1688 B.n305 B.n304 10.6151
R1689 B.n305 B.n148 10.6151
R1690 B.n309 B.n148 10.6151
R1691 B.n310 B.n309 10.6151
R1692 B.n311 B.n310 10.6151
R1693 B.n315 B.n314 10.6151
R1694 B.n316 B.n315 10.6151
R1695 B.n316 B.n142 10.6151
R1696 B.n320 B.n142 10.6151
R1697 B.n321 B.n320 10.6151
R1698 B.n322 B.n321 10.6151
R1699 B.n322 B.n140 10.6151
R1700 B.n326 B.n140 10.6151
R1701 B.n329 B.n328 10.6151
R1702 B.n329 B.n136 10.6151
R1703 B.n333 B.n136 10.6151
R1704 B.n334 B.n333 10.6151
R1705 B.n335 B.n334 10.6151
R1706 B.n335 B.n134 10.6151
R1707 B.n339 B.n134 10.6151
R1708 B.n340 B.n339 10.6151
R1709 B.n341 B.n340 10.6151
R1710 B.n341 B.n132 10.6151
R1711 B.n345 B.n132 10.6151
R1712 B.n346 B.n345 10.6151
R1713 B.n347 B.n346 10.6151
R1714 B.n347 B.n130 10.6151
R1715 B.n351 B.n130 10.6151
R1716 B.n352 B.n351 10.6151
R1717 B.n353 B.n352 10.6151
R1718 B.n353 B.n128 10.6151
R1719 B.n357 B.n128 10.6151
R1720 B.n358 B.n357 10.6151
R1721 B.n359 B.n358 10.6151
R1722 B.n359 B.n126 10.6151
R1723 B.n363 B.n126 10.6151
R1724 B.n364 B.n363 10.6151
R1725 B.n365 B.n364 10.6151
R1726 B.n365 B.n124 10.6151
R1727 B.n369 B.n124 10.6151
R1728 B.n370 B.n369 10.6151
R1729 B.n371 B.n370 10.6151
R1730 B.n371 B.n122 10.6151
R1731 B.n375 B.n122 10.6151
R1732 B.n376 B.n375 10.6151
R1733 B.n377 B.n376 10.6151
R1734 B.n377 B.n120 10.6151
R1735 B.n381 B.n120 10.6151
R1736 B.n382 B.n381 10.6151
R1737 B.n383 B.n382 10.6151
R1738 B.n255 B.n166 10.6151
R1739 B.n251 B.n166 10.6151
R1740 B.n251 B.n250 10.6151
R1741 B.n250 B.n249 10.6151
R1742 B.n249 B.n168 10.6151
R1743 B.n245 B.n168 10.6151
R1744 B.n245 B.n244 10.6151
R1745 B.n244 B.n243 10.6151
R1746 B.n243 B.n170 10.6151
R1747 B.n239 B.n170 10.6151
R1748 B.n239 B.n238 10.6151
R1749 B.n238 B.n237 10.6151
R1750 B.n237 B.n172 10.6151
R1751 B.n233 B.n172 10.6151
R1752 B.n233 B.n232 10.6151
R1753 B.n232 B.n231 10.6151
R1754 B.n231 B.n174 10.6151
R1755 B.n227 B.n174 10.6151
R1756 B.n227 B.n226 10.6151
R1757 B.n226 B.n225 10.6151
R1758 B.n225 B.n176 10.6151
R1759 B.n221 B.n176 10.6151
R1760 B.n221 B.n220 10.6151
R1761 B.n220 B.n219 10.6151
R1762 B.n219 B.n178 10.6151
R1763 B.n215 B.n178 10.6151
R1764 B.n215 B.n214 10.6151
R1765 B.n214 B.n213 10.6151
R1766 B.n213 B.n180 10.6151
R1767 B.n209 B.n180 10.6151
R1768 B.n209 B.n208 10.6151
R1769 B.n208 B.n207 10.6151
R1770 B.n207 B.n182 10.6151
R1771 B.n203 B.n182 10.6151
R1772 B.n203 B.n202 10.6151
R1773 B.n202 B.n201 10.6151
R1774 B.n201 B.n184 10.6151
R1775 B.n197 B.n184 10.6151
R1776 B.n197 B.n196 10.6151
R1777 B.n196 B.n195 10.6151
R1778 B.n195 B.n186 10.6151
R1779 B.n191 B.n186 10.6151
R1780 B.n191 B.n190 10.6151
R1781 B.n190 B.n189 10.6151
R1782 B.n189 B.n0 10.6151
R1783 B.n719 B.n1 10.6151
R1784 B.n719 B.n718 10.6151
R1785 B.n718 B.n717 10.6151
R1786 B.n717 B.n4 10.6151
R1787 B.n713 B.n4 10.6151
R1788 B.n713 B.n712 10.6151
R1789 B.n712 B.n711 10.6151
R1790 B.n711 B.n6 10.6151
R1791 B.n707 B.n6 10.6151
R1792 B.n707 B.n706 10.6151
R1793 B.n706 B.n705 10.6151
R1794 B.n705 B.n8 10.6151
R1795 B.n701 B.n8 10.6151
R1796 B.n701 B.n700 10.6151
R1797 B.n700 B.n699 10.6151
R1798 B.n699 B.n10 10.6151
R1799 B.n695 B.n10 10.6151
R1800 B.n695 B.n694 10.6151
R1801 B.n694 B.n693 10.6151
R1802 B.n693 B.n12 10.6151
R1803 B.n689 B.n12 10.6151
R1804 B.n689 B.n688 10.6151
R1805 B.n688 B.n687 10.6151
R1806 B.n687 B.n14 10.6151
R1807 B.n683 B.n14 10.6151
R1808 B.n683 B.n682 10.6151
R1809 B.n682 B.n681 10.6151
R1810 B.n681 B.n16 10.6151
R1811 B.n677 B.n16 10.6151
R1812 B.n677 B.n676 10.6151
R1813 B.n676 B.n675 10.6151
R1814 B.n675 B.n18 10.6151
R1815 B.n671 B.n18 10.6151
R1816 B.n671 B.n670 10.6151
R1817 B.n670 B.n669 10.6151
R1818 B.n669 B.n20 10.6151
R1819 B.n665 B.n20 10.6151
R1820 B.n665 B.n664 10.6151
R1821 B.n664 B.n663 10.6151
R1822 B.n663 B.n22 10.6151
R1823 B.n659 B.n22 10.6151
R1824 B.n659 B.n658 10.6151
R1825 B.n658 B.n657 10.6151
R1826 B.n657 B.n24 10.6151
R1827 B.n653 B.n24 10.6151
R1828 B.n594 B.n46 6.5566
R1829 B.n582 B.n581 6.5566
R1830 B.n314 B.n146 6.5566
R1831 B.n327 B.n326 6.5566
R1832 B.n597 B.n46 4.05904
R1833 B.n581 B.n580 4.05904
R1834 B.n311 B.n146 4.05904
R1835 B.n328 B.n327 4.05904
R1836 B.n723 B.n0 2.81026
R1837 B.n723 B.n1 2.81026
R1838 VN.n0 VN.t0 98.5052
R1839 VN.n1 VN.t1 98.5052
R1840 VN.n0 VN.t3 97.0695
R1841 VN.n1 VN.t2 97.0695
R1842 VN VN.n1 51.3457
R1843 VN VN.n0 1.75857
R1844 VDD2.n2 VDD2.n0 118.87
R1845 VDD2.n2 VDD2.n1 74.8963
R1846 VDD2.n1 VDD2.t1 3.05836
R1847 VDD2.n1 VDD2.t2 3.05836
R1848 VDD2.n0 VDD2.t3 3.05836
R1849 VDD2.n0 VDD2.t0 3.05836
R1850 VDD2 VDD2.n2 0.0586897
C0 w_n3544_n3094# VTAIL 3.72085f
C1 VTAIL VDD2 5.59132f
C2 VDD1 VP 4.84479f
C3 VDD1 VTAIL 5.528f
C4 w_n3544_n3094# VDD2 1.75825f
C5 VN B 1.35052f
C6 VDD1 w_n3544_n3094# 1.67217f
C7 VDD1 VDD2 1.36149f
C8 VP B 2.1186f
C9 VN VP 6.92095f
C10 VTAIL B 5.00698f
C11 VTAIL VN 4.69723f
C12 w_n3544_n3094# B 10.5342f
C13 VDD2 B 1.54071f
C14 w_n3544_n3094# VN 6.23366f
C15 VN VDD2 4.51526f
C16 VTAIL VP 4.71134f
C17 VDD1 B 1.46607f
C18 VDD1 VN 0.150387f
C19 w_n3544_n3094# VP 6.6927f
C20 VDD2 VP 0.481003f
C21 VDD2 VSUBS 1.131649f
C22 VDD1 VSUBS 6.33983f
C23 VTAIL VSUBS 1.342622f
C24 VN VSUBS 6.21588f
C25 VP VSUBS 2.977541f
C26 B VSUBS 5.330939f
C27 w_n3544_n3094# VSUBS 0.135282p
C28 VDD2.t3 VSUBS 0.231275f
C29 VDD2.t0 VSUBS 0.231275f
C30 VDD2.n0 VSUBS 2.50121f
C31 VDD2.t1 VSUBS 0.231275f
C32 VDD2.t2 VSUBS 0.231275f
C33 VDD2.n1 VSUBS 1.76263f
C34 VDD2.n2 VSUBS 4.57704f
C35 VN.t0 VSUBS 3.59159f
C36 VN.t3 VSUBS 3.57304f
C37 VN.n0 VSUBS 2.1221f
C38 VN.t1 VSUBS 3.59159f
C39 VN.t2 VSUBS 3.57304f
C40 VN.n1 VSUBS 3.91196f
C41 B.n0 VSUBS 0.004551f
C42 B.n1 VSUBS 0.004551f
C43 B.n2 VSUBS 0.007197f
C44 B.n3 VSUBS 0.007197f
C45 B.n4 VSUBS 0.007197f
C46 B.n5 VSUBS 0.007197f
C47 B.n6 VSUBS 0.007197f
C48 B.n7 VSUBS 0.007197f
C49 B.n8 VSUBS 0.007197f
C50 B.n9 VSUBS 0.007197f
C51 B.n10 VSUBS 0.007197f
C52 B.n11 VSUBS 0.007197f
C53 B.n12 VSUBS 0.007197f
C54 B.n13 VSUBS 0.007197f
C55 B.n14 VSUBS 0.007197f
C56 B.n15 VSUBS 0.007197f
C57 B.n16 VSUBS 0.007197f
C58 B.n17 VSUBS 0.007197f
C59 B.n18 VSUBS 0.007197f
C60 B.n19 VSUBS 0.007197f
C61 B.n20 VSUBS 0.007197f
C62 B.n21 VSUBS 0.007197f
C63 B.n22 VSUBS 0.007197f
C64 B.n23 VSUBS 0.007197f
C65 B.n24 VSUBS 0.007197f
C66 B.n25 VSUBS 0.016689f
C67 B.n26 VSUBS 0.007197f
C68 B.n27 VSUBS 0.007197f
C69 B.n28 VSUBS 0.007197f
C70 B.n29 VSUBS 0.007197f
C71 B.n30 VSUBS 0.007197f
C72 B.n31 VSUBS 0.007197f
C73 B.n32 VSUBS 0.007197f
C74 B.n33 VSUBS 0.007197f
C75 B.n34 VSUBS 0.007197f
C76 B.n35 VSUBS 0.007197f
C77 B.n36 VSUBS 0.007197f
C78 B.n37 VSUBS 0.007197f
C79 B.n38 VSUBS 0.007197f
C80 B.n39 VSUBS 0.007197f
C81 B.n40 VSUBS 0.007197f
C82 B.n41 VSUBS 0.007197f
C83 B.n42 VSUBS 0.007197f
C84 B.n43 VSUBS 0.007197f
C85 B.t8 VSUBS 0.185952f
C86 B.t7 VSUBS 0.230908f
C87 B.t6 VSUBS 2.03534f
C88 B.n44 VSUBS 0.36966f
C89 B.n45 VSUBS 0.244794f
C90 B.n46 VSUBS 0.016674f
C91 B.n47 VSUBS 0.007197f
C92 B.n48 VSUBS 0.007197f
C93 B.n49 VSUBS 0.007197f
C94 B.n50 VSUBS 0.007197f
C95 B.n51 VSUBS 0.007197f
C96 B.t5 VSUBS 0.185955f
C97 B.t4 VSUBS 0.23091f
C98 B.t3 VSUBS 2.03534f
C99 B.n52 VSUBS 0.369658f
C100 B.n53 VSUBS 0.244791f
C101 B.n54 VSUBS 0.007197f
C102 B.n55 VSUBS 0.007197f
C103 B.n56 VSUBS 0.007197f
C104 B.n57 VSUBS 0.007197f
C105 B.n58 VSUBS 0.007197f
C106 B.n59 VSUBS 0.007197f
C107 B.n60 VSUBS 0.007197f
C108 B.n61 VSUBS 0.007197f
C109 B.n62 VSUBS 0.007197f
C110 B.n63 VSUBS 0.007197f
C111 B.n64 VSUBS 0.007197f
C112 B.n65 VSUBS 0.007197f
C113 B.n66 VSUBS 0.007197f
C114 B.n67 VSUBS 0.007197f
C115 B.n68 VSUBS 0.007197f
C116 B.n69 VSUBS 0.007197f
C117 B.n70 VSUBS 0.007197f
C118 B.n71 VSUBS 0.007197f
C119 B.n72 VSUBS 0.016601f
C120 B.n73 VSUBS 0.007197f
C121 B.n74 VSUBS 0.007197f
C122 B.n75 VSUBS 0.007197f
C123 B.n76 VSUBS 0.007197f
C124 B.n77 VSUBS 0.007197f
C125 B.n78 VSUBS 0.007197f
C126 B.n79 VSUBS 0.007197f
C127 B.n80 VSUBS 0.007197f
C128 B.n81 VSUBS 0.007197f
C129 B.n82 VSUBS 0.007197f
C130 B.n83 VSUBS 0.007197f
C131 B.n84 VSUBS 0.007197f
C132 B.n85 VSUBS 0.007197f
C133 B.n86 VSUBS 0.007197f
C134 B.n87 VSUBS 0.007197f
C135 B.n88 VSUBS 0.007197f
C136 B.n89 VSUBS 0.007197f
C137 B.n90 VSUBS 0.007197f
C138 B.n91 VSUBS 0.007197f
C139 B.n92 VSUBS 0.007197f
C140 B.n93 VSUBS 0.007197f
C141 B.n94 VSUBS 0.007197f
C142 B.n95 VSUBS 0.007197f
C143 B.n96 VSUBS 0.007197f
C144 B.n97 VSUBS 0.007197f
C145 B.n98 VSUBS 0.007197f
C146 B.n99 VSUBS 0.007197f
C147 B.n100 VSUBS 0.007197f
C148 B.n101 VSUBS 0.007197f
C149 B.n102 VSUBS 0.007197f
C150 B.n103 VSUBS 0.007197f
C151 B.n104 VSUBS 0.007197f
C152 B.n105 VSUBS 0.007197f
C153 B.n106 VSUBS 0.007197f
C154 B.n107 VSUBS 0.007197f
C155 B.n108 VSUBS 0.007197f
C156 B.n109 VSUBS 0.007197f
C157 B.n110 VSUBS 0.007197f
C158 B.n111 VSUBS 0.007197f
C159 B.n112 VSUBS 0.007197f
C160 B.n113 VSUBS 0.007197f
C161 B.n114 VSUBS 0.007197f
C162 B.n115 VSUBS 0.007197f
C163 B.n116 VSUBS 0.007197f
C164 B.n117 VSUBS 0.007197f
C165 B.n118 VSUBS 0.015698f
C166 B.n119 VSUBS 0.007197f
C167 B.n120 VSUBS 0.007197f
C168 B.n121 VSUBS 0.007197f
C169 B.n122 VSUBS 0.007197f
C170 B.n123 VSUBS 0.007197f
C171 B.n124 VSUBS 0.007197f
C172 B.n125 VSUBS 0.007197f
C173 B.n126 VSUBS 0.007197f
C174 B.n127 VSUBS 0.007197f
C175 B.n128 VSUBS 0.007197f
C176 B.n129 VSUBS 0.007197f
C177 B.n130 VSUBS 0.007197f
C178 B.n131 VSUBS 0.007197f
C179 B.n132 VSUBS 0.007197f
C180 B.n133 VSUBS 0.007197f
C181 B.n134 VSUBS 0.007197f
C182 B.n135 VSUBS 0.007197f
C183 B.n136 VSUBS 0.007197f
C184 B.n137 VSUBS 0.007197f
C185 B.t10 VSUBS 0.185955f
C186 B.t11 VSUBS 0.23091f
C187 B.t9 VSUBS 2.03534f
C188 B.n138 VSUBS 0.369658f
C189 B.n139 VSUBS 0.244791f
C190 B.n140 VSUBS 0.007197f
C191 B.n141 VSUBS 0.007197f
C192 B.n142 VSUBS 0.007197f
C193 B.n143 VSUBS 0.007197f
C194 B.t1 VSUBS 0.185952f
C195 B.t2 VSUBS 0.230908f
C196 B.t0 VSUBS 2.03534f
C197 B.n144 VSUBS 0.36966f
C198 B.n145 VSUBS 0.244794f
C199 B.n146 VSUBS 0.016674f
C200 B.n147 VSUBS 0.007197f
C201 B.n148 VSUBS 0.007197f
C202 B.n149 VSUBS 0.007197f
C203 B.n150 VSUBS 0.007197f
C204 B.n151 VSUBS 0.007197f
C205 B.n152 VSUBS 0.007197f
C206 B.n153 VSUBS 0.007197f
C207 B.n154 VSUBS 0.007197f
C208 B.n155 VSUBS 0.007197f
C209 B.n156 VSUBS 0.007197f
C210 B.n157 VSUBS 0.007197f
C211 B.n158 VSUBS 0.007197f
C212 B.n159 VSUBS 0.007197f
C213 B.n160 VSUBS 0.007197f
C214 B.n161 VSUBS 0.007197f
C215 B.n162 VSUBS 0.007197f
C216 B.n163 VSUBS 0.007197f
C217 B.n164 VSUBS 0.007197f
C218 B.n165 VSUBS 0.016689f
C219 B.n166 VSUBS 0.007197f
C220 B.n167 VSUBS 0.007197f
C221 B.n168 VSUBS 0.007197f
C222 B.n169 VSUBS 0.007197f
C223 B.n170 VSUBS 0.007197f
C224 B.n171 VSUBS 0.007197f
C225 B.n172 VSUBS 0.007197f
C226 B.n173 VSUBS 0.007197f
C227 B.n174 VSUBS 0.007197f
C228 B.n175 VSUBS 0.007197f
C229 B.n176 VSUBS 0.007197f
C230 B.n177 VSUBS 0.007197f
C231 B.n178 VSUBS 0.007197f
C232 B.n179 VSUBS 0.007197f
C233 B.n180 VSUBS 0.007197f
C234 B.n181 VSUBS 0.007197f
C235 B.n182 VSUBS 0.007197f
C236 B.n183 VSUBS 0.007197f
C237 B.n184 VSUBS 0.007197f
C238 B.n185 VSUBS 0.007197f
C239 B.n186 VSUBS 0.007197f
C240 B.n187 VSUBS 0.007197f
C241 B.n188 VSUBS 0.007197f
C242 B.n189 VSUBS 0.007197f
C243 B.n190 VSUBS 0.007197f
C244 B.n191 VSUBS 0.007197f
C245 B.n192 VSUBS 0.007197f
C246 B.n193 VSUBS 0.007197f
C247 B.n194 VSUBS 0.007197f
C248 B.n195 VSUBS 0.007197f
C249 B.n196 VSUBS 0.007197f
C250 B.n197 VSUBS 0.007197f
C251 B.n198 VSUBS 0.007197f
C252 B.n199 VSUBS 0.007197f
C253 B.n200 VSUBS 0.007197f
C254 B.n201 VSUBS 0.007197f
C255 B.n202 VSUBS 0.007197f
C256 B.n203 VSUBS 0.007197f
C257 B.n204 VSUBS 0.007197f
C258 B.n205 VSUBS 0.007197f
C259 B.n206 VSUBS 0.007197f
C260 B.n207 VSUBS 0.007197f
C261 B.n208 VSUBS 0.007197f
C262 B.n209 VSUBS 0.007197f
C263 B.n210 VSUBS 0.007197f
C264 B.n211 VSUBS 0.007197f
C265 B.n212 VSUBS 0.007197f
C266 B.n213 VSUBS 0.007197f
C267 B.n214 VSUBS 0.007197f
C268 B.n215 VSUBS 0.007197f
C269 B.n216 VSUBS 0.007197f
C270 B.n217 VSUBS 0.007197f
C271 B.n218 VSUBS 0.007197f
C272 B.n219 VSUBS 0.007197f
C273 B.n220 VSUBS 0.007197f
C274 B.n221 VSUBS 0.007197f
C275 B.n222 VSUBS 0.007197f
C276 B.n223 VSUBS 0.007197f
C277 B.n224 VSUBS 0.007197f
C278 B.n225 VSUBS 0.007197f
C279 B.n226 VSUBS 0.007197f
C280 B.n227 VSUBS 0.007197f
C281 B.n228 VSUBS 0.007197f
C282 B.n229 VSUBS 0.007197f
C283 B.n230 VSUBS 0.007197f
C284 B.n231 VSUBS 0.007197f
C285 B.n232 VSUBS 0.007197f
C286 B.n233 VSUBS 0.007197f
C287 B.n234 VSUBS 0.007197f
C288 B.n235 VSUBS 0.007197f
C289 B.n236 VSUBS 0.007197f
C290 B.n237 VSUBS 0.007197f
C291 B.n238 VSUBS 0.007197f
C292 B.n239 VSUBS 0.007197f
C293 B.n240 VSUBS 0.007197f
C294 B.n241 VSUBS 0.007197f
C295 B.n242 VSUBS 0.007197f
C296 B.n243 VSUBS 0.007197f
C297 B.n244 VSUBS 0.007197f
C298 B.n245 VSUBS 0.007197f
C299 B.n246 VSUBS 0.007197f
C300 B.n247 VSUBS 0.007197f
C301 B.n248 VSUBS 0.007197f
C302 B.n249 VSUBS 0.007197f
C303 B.n250 VSUBS 0.007197f
C304 B.n251 VSUBS 0.007197f
C305 B.n252 VSUBS 0.007197f
C306 B.n253 VSUBS 0.007197f
C307 B.n254 VSUBS 0.015698f
C308 B.n255 VSUBS 0.015698f
C309 B.n256 VSUBS 0.016689f
C310 B.n257 VSUBS 0.007197f
C311 B.n258 VSUBS 0.007197f
C312 B.n259 VSUBS 0.007197f
C313 B.n260 VSUBS 0.007197f
C314 B.n261 VSUBS 0.007197f
C315 B.n262 VSUBS 0.007197f
C316 B.n263 VSUBS 0.007197f
C317 B.n264 VSUBS 0.007197f
C318 B.n265 VSUBS 0.007197f
C319 B.n266 VSUBS 0.007197f
C320 B.n267 VSUBS 0.007197f
C321 B.n268 VSUBS 0.007197f
C322 B.n269 VSUBS 0.007197f
C323 B.n270 VSUBS 0.007197f
C324 B.n271 VSUBS 0.007197f
C325 B.n272 VSUBS 0.007197f
C326 B.n273 VSUBS 0.007197f
C327 B.n274 VSUBS 0.007197f
C328 B.n275 VSUBS 0.007197f
C329 B.n276 VSUBS 0.007197f
C330 B.n277 VSUBS 0.007197f
C331 B.n278 VSUBS 0.007197f
C332 B.n279 VSUBS 0.007197f
C333 B.n280 VSUBS 0.007197f
C334 B.n281 VSUBS 0.007197f
C335 B.n282 VSUBS 0.007197f
C336 B.n283 VSUBS 0.007197f
C337 B.n284 VSUBS 0.007197f
C338 B.n285 VSUBS 0.007197f
C339 B.n286 VSUBS 0.007197f
C340 B.n287 VSUBS 0.007197f
C341 B.n288 VSUBS 0.007197f
C342 B.n289 VSUBS 0.007197f
C343 B.n290 VSUBS 0.007197f
C344 B.n291 VSUBS 0.007197f
C345 B.n292 VSUBS 0.007197f
C346 B.n293 VSUBS 0.007197f
C347 B.n294 VSUBS 0.007197f
C348 B.n295 VSUBS 0.007197f
C349 B.n296 VSUBS 0.007197f
C350 B.n297 VSUBS 0.007197f
C351 B.n298 VSUBS 0.007197f
C352 B.n299 VSUBS 0.007197f
C353 B.n300 VSUBS 0.007197f
C354 B.n301 VSUBS 0.007197f
C355 B.n302 VSUBS 0.007197f
C356 B.n303 VSUBS 0.007197f
C357 B.n304 VSUBS 0.007197f
C358 B.n305 VSUBS 0.007197f
C359 B.n306 VSUBS 0.007197f
C360 B.n307 VSUBS 0.007197f
C361 B.n308 VSUBS 0.007197f
C362 B.n309 VSUBS 0.007197f
C363 B.n310 VSUBS 0.007197f
C364 B.n311 VSUBS 0.004974f
C365 B.n312 VSUBS 0.007197f
C366 B.n313 VSUBS 0.007197f
C367 B.n314 VSUBS 0.005821f
C368 B.n315 VSUBS 0.007197f
C369 B.n316 VSUBS 0.007197f
C370 B.n317 VSUBS 0.007197f
C371 B.n318 VSUBS 0.007197f
C372 B.n319 VSUBS 0.007197f
C373 B.n320 VSUBS 0.007197f
C374 B.n321 VSUBS 0.007197f
C375 B.n322 VSUBS 0.007197f
C376 B.n323 VSUBS 0.007197f
C377 B.n324 VSUBS 0.007197f
C378 B.n325 VSUBS 0.007197f
C379 B.n326 VSUBS 0.005821f
C380 B.n327 VSUBS 0.016674f
C381 B.n328 VSUBS 0.004974f
C382 B.n329 VSUBS 0.007197f
C383 B.n330 VSUBS 0.007197f
C384 B.n331 VSUBS 0.007197f
C385 B.n332 VSUBS 0.007197f
C386 B.n333 VSUBS 0.007197f
C387 B.n334 VSUBS 0.007197f
C388 B.n335 VSUBS 0.007197f
C389 B.n336 VSUBS 0.007197f
C390 B.n337 VSUBS 0.007197f
C391 B.n338 VSUBS 0.007197f
C392 B.n339 VSUBS 0.007197f
C393 B.n340 VSUBS 0.007197f
C394 B.n341 VSUBS 0.007197f
C395 B.n342 VSUBS 0.007197f
C396 B.n343 VSUBS 0.007197f
C397 B.n344 VSUBS 0.007197f
C398 B.n345 VSUBS 0.007197f
C399 B.n346 VSUBS 0.007197f
C400 B.n347 VSUBS 0.007197f
C401 B.n348 VSUBS 0.007197f
C402 B.n349 VSUBS 0.007197f
C403 B.n350 VSUBS 0.007197f
C404 B.n351 VSUBS 0.007197f
C405 B.n352 VSUBS 0.007197f
C406 B.n353 VSUBS 0.007197f
C407 B.n354 VSUBS 0.007197f
C408 B.n355 VSUBS 0.007197f
C409 B.n356 VSUBS 0.007197f
C410 B.n357 VSUBS 0.007197f
C411 B.n358 VSUBS 0.007197f
C412 B.n359 VSUBS 0.007197f
C413 B.n360 VSUBS 0.007197f
C414 B.n361 VSUBS 0.007197f
C415 B.n362 VSUBS 0.007197f
C416 B.n363 VSUBS 0.007197f
C417 B.n364 VSUBS 0.007197f
C418 B.n365 VSUBS 0.007197f
C419 B.n366 VSUBS 0.007197f
C420 B.n367 VSUBS 0.007197f
C421 B.n368 VSUBS 0.007197f
C422 B.n369 VSUBS 0.007197f
C423 B.n370 VSUBS 0.007197f
C424 B.n371 VSUBS 0.007197f
C425 B.n372 VSUBS 0.007197f
C426 B.n373 VSUBS 0.007197f
C427 B.n374 VSUBS 0.007197f
C428 B.n375 VSUBS 0.007197f
C429 B.n376 VSUBS 0.007197f
C430 B.n377 VSUBS 0.007197f
C431 B.n378 VSUBS 0.007197f
C432 B.n379 VSUBS 0.007197f
C433 B.n380 VSUBS 0.007197f
C434 B.n381 VSUBS 0.007197f
C435 B.n382 VSUBS 0.007197f
C436 B.n383 VSUBS 0.016689f
C437 B.n384 VSUBS 0.016689f
C438 B.n385 VSUBS 0.015698f
C439 B.n386 VSUBS 0.007197f
C440 B.n387 VSUBS 0.007197f
C441 B.n388 VSUBS 0.007197f
C442 B.n389 VSUBS 0.007197f
C443 B.n390 VSUBS 0.007197f
C444 B.n391 VSUBS 0.007197f
C445 B.n392 VSUBS 0.007197f
C446 B.n393 VSUBS 0.007197f
C447 B.n394 VSUBS 0.007197f
C448 B.n395 VSUBS 0.007197f
C449 B.n396 VSUBS 0.007197f
C450 B.n397 VSUBS 0.007197f
C451 B.n398 VSUBS 0.007197f
C452 B.n399 VSUBS 0.007197f
C453 B.n400 VSUBS 0.007197f
C454 B.n401 VSUBS 0.007197f
C455 B.n402 VSUBS 0.007197f
C456 B.n403 VSUBS 0.007197f
C457 B.n404 VSUBS 0.007197f
C458 B.n405 VSUBS 0.007197f
C459 B.n406 VSUBS 0.007197f
C460 B.n407 VSUBS 0.007197f
C461 B.n408 VSUBS 0.007197f
C462 B.n409 VSUBS 0.007197f
C463 B.n410 VSUBS 0.007197f
C464 B.n411 VSUBS 0.007197f
C465 B.n412 VSUBS 0.007197f
C466 B.n413 VSUBS 0.007197f
C467 B.n414 VSUBS 0.007197f
C468 B.n415 VSUBS 0.007197f
C469 B.n416 VSUBS 0.007197f
C470 B.n417 VSUBS 0.007197f
C471 B.n418 VSUBS 0.007197f
C472 B.n419 VSUBS 0.007197f
C473 B.n420 VSUBS 0.007197f
C474 B.n421 VSUBS 0.007197f
C475 B.n422 VSUBS 0.007197f
C476 B.n423 VSUBS 0.007197f
C477 B.n424 VSUBS 0.007197f
C478 B.n425 VSUBS 0.007197f
C479 B.n426 VSUBS 0.007197f
C480 B.n427 VSUBS 0.007197f
C481 B.n428 VSUBS 0.007197f
C482 B.n429 VSUBS 0.007197f
C483 B.n430 VSUBS 0.007197f
C484 B.n431 VSUBS 0.007197f
C485 B.n432 VSUBS 0.007197f
C486 B.n433 VSUBS 0.007197f
C487 B.n434 VSUBS 0.007197f
C488 B.n435 VSUBS 0.007197f
C489 B.n436 VSUBS 0.007197f
C490 B.n437 VSUBS 0.007197f
C491 B.n438 VSUBS 0.007197f
C492 B.n439 VSUBS 0.007197f
C493 B.n440 VSUBS 0.007197f
C494 B.n441 VSUBS 0.007197f
C495 B.n442 VSUBS 0.007197f
C496 B.n443 VSUBS 0.007197f
C497 B.n444 VSUBS 0.007197f
C498 B.n445 VSUBS 0.007197f
C499 B.n446 VSUBS 0.007197f
C500 B.n447 VSUBS 0.007197f
C501 B.n448 VSUBS 0.007197f
C502 B.n449 VSUBS 0.007197f
C503 B.n450 VSUBS 0.007197f
C504 B.n451 VSUBS 0.007197f
C505 B.n452 VSUBS 0.007197f
C506 B.n453 VSUBS 0.007197f
C507 B.n454 VSUBS 0.007197f
C508 B.n455 VSUBS 0.007197f
C509 B.n456 VSUBS 0.007197f
C510 B.n457 VSUBS 0.007197f
C511 B.n458 VSUBS 0.007197f
C512 B.n459 VSUBS 0.007197f
C513 B.n460 VSUBS 0.007197f
C514 B.n461 VSUBS 0.007197f
C515 B.n462 VSUBS 0.007197f
C516 B.n463 VSUBS 0.007197f
C517 B.n464 VSUBS 0.007197f
C518 B.n465 VSUBS 0.007197f
C519 B.n466 VSUBS 0.007197f
C520 B.n467 VSUBS 0.007197f
C521 B.n468 VSUBS 0.007197f
C522 B.n469 VSUBS 0.007197f
C523 B.n470 VSUBS 0.007197f
C524 B.n471 VSUBS 0.007197f
C525 B.n472 VSUBS 0.007197f
C526 B.n473 VSUBS 0.007197f
C527 B.n474 VSUBS 0.007197f
C528 B.n475 VSUBS 0.007197f
C529 B.n476 VSUBS 0.007197f
C530 B.n477 VSUBS 0.007197f
C531 B.n478 VSUBS 0.007197f
C532 B.n479 VSUBS 0.007197f
C533 B.n480 VSUBS 0.007197f
C534 B.n481 VSUBS 0.007197f
C535 B.n482 VSUBS 0.007197f
C536 B.n483 VSUBS 0.007197f
C537 B.n484 VSUBS 0.007197f
C538 B.n485 VSUBS 0.007197f
C539 B.n486 VSUBS 0.007197f
C540 B.n487 VSUBS 0.007197f
C541 B.n488 VSUBS 0.007197f
C542 B.n489 VSUBS 0.007197f
C543 B.n490 VSUBS 0.007197f
C544 B.n491 VSUBS 0.007197f
C545 B.n492 VSUBS 0.007197f
C546 B.n493 VSUBS 0.007197f
C547 B.n494 VSUBS 0.007197f
C548 B.n495 VSUBS 0.007197f
C549 B.n496 VSUBS 0.007197f
C550 B.n497 VSUBS 0.007197f
C551 B.n498 VSUBS 0.007197f
C552 B.n499 VSUBS 0.007197f
C553 B.n500 VSUBS 0.007197f
C554 B.n501 VSUBS 0.007197f
C555 B.n502 VSUBS 0.007197f
C556 B.n503 VSUBS 0.007197f
C557 B.n504 VSUBS 0.007197f
C558 B.n505 VSUBS 0.007197f
C559 B.n506 VSUBS 0.007197f
C560 B.n507 VSUBS 0.007197f
C561 B.n508 VSUBS 0.007197f
C562 B.n509 VSUBS 0.007197f
C563 B.n510 VSUBS 0.007197f
C564 B.n511 VSUBS 0.007197f
C565 B.n512 VSUBS 0.007197f
C566 B.n513 VSUBS 0.007197f
C567 B.n514 VSUBS 0.007197f
C568 B.n515 VSUBS 0.007197f
C569 B.n516 VSUBS 0.007197f
C570 B.n517 VSUBS 0.007197f
C571 B.n518 VSUBS 0.007197f
C572 B.n519 VSUBS 0.007197f
C573 B.n520 VSUBS 0.007197f
C574 B.n521 VSUBS 0.007197f
C575 B.n522 VSUBS 0.007197f
C576 B.n523 VSUBS 0.015698f
C577 B.n524 VSUBS 0.016689f
C578 B.n525 VSUBS 0.015786f
C579 B.n526 VSUBS 0.007197f
C580 B.n527 VSUBS 0.007197f
C581 B.n528 VSUBS 0.007197f
C582 B.n529 VSUBS 0.007197f
C583 B.n530 VSUBS 0.007197f
C584 B.n531 VSUBS 0.007197f
C585 B.n532 VSUBS 0.007197f
C586 B.n533 VSUBS 0.007197f
C587 B.n534 VSUBS 0.007197f
C588 B.n535 VSUBS 0.007197f
C589 B.n536 VSUBS 0.007197f
C590 B.n537 VSUBS 0.007197f
C591 B.n538 VSUBS 0.007197f
C592 B.n539 VSUBS 0.007197f
C593 B.n540 VSUBS 0.007197f
C594 B.n541 VSUBS 0.007197f
C595 B.n542 VSUBS 0.007197f
C596 B.n543 VSUBS 0.007197f
C597 B.n544 VSUBS 0.007197f
C598 B.n545 VSUBS 0.007197f
C599 B.n546 VSUBS 0.007197f
C600 B.n547 VSUBS 0.007197f
C601 B.n548 VSUBS 0.007197f
C602 B.n549 VSUBS 0.007197f
C603 B.n550 VSUBS 0.007197f
C604 B.n551 VSUBS 0.007197f
C605 B.n552 VSUBS 0.007197f
C606 B.n553 VSUBS 0.007197f
C607 B.n554 VSUBS 0.007197f
C608 B.n555 VSUBS 0.007197f
C609 B.n556 VSUBS 0.007197f
C610 B.n557 VSUBS 0.007197f
C611 B.n558 VSUBS 0.007197f
C612 B.n559 VSUBS 0.007197f
C613 B.n560 VSUBS 0.007197f
C614 B.n561 VSUBS 0.007197f
C615 B.n562 VSUBS 0.007197f
C616 B.n563 VSUBS 0.007197f
C617 B.n564 VSUBS 0.007197f
C618 B.n565 VSUBS 0.007197f
C619 B.n566 VSUBS 0.007197f
C620 B.n567 VSUBS 0.007197f
C621 B.n568 VSUBS 0.007197f
C622 B.n569 VSUBS 0.007197f
C623 B.n570 VSUBS 0.007197f
C624 B.n571 VSUBS 0.007197f
C625 B.n572 VSUBS 0.007197f
C626 B.n573 VSUBS 0.007197f
C627 B.n574 VSUBS 0.007197f
C628 B.n575 VSUBS 0.007197f
C629 B.n576 VSUBS 0.007197f
C630 B.n577 VSUBS 0.007197f
C631 B.n578 VSUBS 0.007197f
C632 B.n579 VSUBS 0.007197f
C633 B.n580 VSUBS 0.004974f
C634 B.n581 VSUBS 0.016674f
C635 B.n582 VSUBS 0.005821f
C636 B.n583 VSUBS 0.007197f
C637 B.n584 VSUBS 0.007197f
C638 B.n585 VSUBS 0.007197f
C639 B.n586 VSUBS 0.007197f
C640 B.n587 VSUBS 0.007197f
C641 B.n588 VSUBS 0.007197f
C642 B.n589 VSUBS 0.007197f
C643 B.n590 VSUBS 0.007197f
C644 B.n591 VSUBS 0.007197f
C645 B.n592 VSUBS 0.007197f
C646 B.n593 VSUBS 0.007197f
C647 B.n594 VSUBS 0.005821f
C648 B.n595 VSUBS 0.007197f
C649 B.n596 VSUBS 0.007197f
C650 B.n597 VSUBS 0.004974f
C651 B.n598 VSUBS 0.007197f
C652 B.n599 VSUBS 0.007197f
C653 B.n600 VSUBS 0.007197f
C654 B.n601 VSUBS 0.007197f
C655 B.n602 VSUBS 0.007197f
C656 B.n603 VSUBS 0.007197f
C657 B.n604 VSUBS 0.007197f
C658 B.n605 VSUBS 0.007197f
C659 B.n606 VSUBS 0.007197f
C660 B.n607 VSUBS 0.007197f
C661 B.n608 VSUBS 0.007197f
C662 B.n609 VSUBS 0.007197f
C663 B.n610 VSUBS 0.007197f
C664 B.n611 VSUBS 0.007197f
C665 B.n612 VSUBS 0.007197f
C666 B.n613 VSUBS 0.007197f
C667 B.n614 VSUBS 0.007197f
C668 B.n615 VSUBS 0.007197f
C669 B.n616 VSUBS 0.007197f
C670 B.n617 VSUBS 0.007197f
C671 B.n618 VSUBS 0.007197f
C672 B.n619 VSUBS 0.007197f
C673 B.n620 VSUBS 0.007197f
C674 B.n621 VSUBS 0.007197f
C675 B.n622 VSUBS 0.007197f
C676 B.n623 VSUBS 0.007197f
C677 B.n624 VSUBS 0.007197f
C678 B.n625 VSUBS 0.007197f
C679 B.n626 VSUBS 0.007197f
C680 B.n627 VSUBS 0.007197f
C681 B.n628 VSUBS 0.007197f
C682 B.n629 VSUBS 0.007197f
C683 B.n630 VSUBS 0.007197f
C684 B.n631 VSUBS 0.007197f
C685 B.n632 VSUBS 0.007197f
C686 B.n633 VSUBS 0.007197f
C687 B.n634 VSUBS 0.007197f
C688 B.n635 VSUBS 0.007197f
C689 B.n636 VSUBS 0.007197f
C690 B.n637 VSUBS 0.007197f
C691 B.n638 VSUBS 0.007197f
C692 B.n639 VSUBS 0.007197f
C693 B.n640 VSUBS 0.007197f
C694 B.n641 VSUBS 0.007197f
C695 B.n642 VSUBS 0.007197f
C696 B.n643 VSUBS 0.007197f
C697 B.n644 VSUBS 0.007197f
C698 B.n645 VSUBS 0.007197f
C699 B.n646 VSUBS 0.007197f
C700 B.n647 VSUBS 0.007197f
C701 B.n648 VSUBS 0.007197f
C702 B.n649 VSUBS 0.007197f
C703 B.n650 VSUBS 0.007197f
C704 B.n651 VSUBS 0.007197f
C705 B.n652 VSUBS 0.016689f
C706 B.n653 VSUBS 0.015698f
C707 B.n654 VSUBS 0.015698f
C708 B.n655 VSUBS 0.007197f
C709 B.n656 VSUBS 0.007197f
C710 B.n657 VSUBS 0.007197f
C711 B.n658 VSUBS 0.007197f
C712 B.n659 VSUBS 0.007197f
C713 B.n660 VSUBS 0.007197f
C714 B.n661 VSUBS 0.007197f
C715 B.n662 VSUBS 0.007197f
C716 B.n663 VSUBS 0.007197f
C717 B.n664 VSUBS 0.007197f
C718 B.n665 VSUBS 0.007197f
C719 B.n666 VSUBS 0.007197f
C720 B.n667 VSUBS 0.007197f
C721 B.n668 VSUBS 0.007197f
C722 B.n669 VSUBS 0.007197f
C723 B.n670 VSUBS 0.007197f
C724 B.n671 VSUBS 0.007197f
C725 B.n672 VSUBS 0.007197f
C726 B.n673 VSUBS 0.007197f
C727 B.n674 VSUBS 0.007197f
C728 B.n675 VSUBS 0.007197f
C729 B.n676 VSUBS 0.007197f
C730 B.n677 VSUBS 0.007197f
C731 B.n678 VSUBS 0.007197f
C732 B.n679 VSUBS 0.007197f
C733 B.n680 VSUBS 0.007197f
C734 B.n681 VSUBS 0.007197f
C735 B.n682 VSUBS 0.007197f
C736 B.n683 VSUBS 0.007197f
C737 B.n684 VSUBS 0.007197f
C738 B.n685 VSUBS 0.007197f
C739 B.n686 VSUBS 0.007197f
C740 B.n687 VSUBS 0.007197f
C741 B.n688 VSUBS 0.007197f
C742 B.n689 VSUBS 0.007197f
C743 B.n690 VSUBS 0.007197f
C744 B.n691 VSUBS 0.007197f
C745 B.n692 VSUBS 0.007197f
C746 B.n693 VSUBS 0.007197f
C747 B.n694 VSUBS 0.007197f
C748 B.n695 VSUBS 0.007197f
C749 B.n696 VSUBS 0.007197f
C750 B.n697 VSUBS 0.007197f
C751 B.n698 VSUBS 0.007197f
C752 B.n699 VSUBS 0.007197f
C753 B.n700 VSUBS 0.007197f
C754 B.n701 VSUBS 0.007197f
C755 B.n702 VSUBS 0.007197f
C756 B.n703 VSUBS 0.007197f
C757 B.n704 VSUBS 0.007197f
C758 B.n705 VSUBS 0.007197f
C759 B.n706 VSUBS 0.007197f
C760 B.n707 VSUBS 0.007197f
C761 B.n708 VSUBS 0.007197f
C762 B.n709 VSUBS 0.007197f
C763 B.n710 VSUBS 0.007197f
C764 B.n711 VSUBS 0.007197f
C765 B.n712 VSUBS 0.007197f
C766 B.n713 VSUBS 0.007197f
C767 B.n714 VSUBS 0.007197f
C768 B.n715 VSUBS 0.007197f
C769 B.n716 VSUBS 0.007197f
C770 B.n717 VSUBS 0.007197f
C771 B.n718 VSUBS 0.007197f
C772 B.n719 VSUBS 0.007197f
C773 B.n720 VSUBS 0.007197f
C774 B.n721 VSUBS 0.007197f
C775 B.n722 VSUBS 0.007197f
C776 B.n723 VSUBS 0.016296f
C777 VDD1.t1 VSUBS 0.233503f
C778 VDD1.t2 VSUBS 0.233503f
C779 VDD1.n0 VSUBS 1.78029f
C780 VDD1.t0 VSUBS 0.233503f
C781 VDD1.t3 VSUBS 0.233503f
C782 VDD1.n1 VSUBS 2.55131f
C783 VTAIL.n0 VSUBS 0.02631f
C784 VTAIL.n1 VSUBS 0.02531f
C785 VTAIL.n2 VSUBS 0.013601f
C786 VTAIL.n3 VSUBS 0.032147f
C787 VTAIL.n4 VSUBS 0.014401f
C788 VTAIL.n5 VSUBS 0.02531f
C789 VTAIL.n6 VSUBS 0.013601f
C790 VTAIL.n7 VSUBS 0.032147f
C791 VTAIL.n8 VSUBS 0.014401f
C792 VTAIL.n9 VSUBS 0.02531f
C793 VTAIL.n10 VSUBS 0.013601f
C794 VTAIL.n11 VSUBS 0.032147f
C795 VTAIL.n12 VSUBS 0.014401f
C796 VTAIL.n13 VSUBS 0.02531f
C797 VTAIL.n14 VSUBS 0.013601f
C798 VTAIL.n15 VSUBS 0.032147f
C799 VTAIL.n16 VSUBS 0.014401f
C800 VTAIL.n17 VSUBS 0.183659f
C801 VTAIL.t1 VSUBS 0.069162f
C802 VTAIL.n18 VSUBS 0.02411f
C803 VTAIL.n19 VSUBS 0.024183f
C804 VTAIL.n20 VSUBS 0.013601f
C805 VTAIL.n21 VSUBS 1.09162f
C806 VTAIL.n22 VSUBS 0.02531f
C807 VTAIL.n23 VSUBS 0.013601f
C808 VTAIL.n24 VSUBS 0.014401f
C809 VTAIL.n25 VSUBS 0.032147f
C810 VTAIL.n26 VSUBS 0.032147f
C811 VTAIL.n27 VSUBS 0.014401f
C812 VTAIL.n28 VSUBS 0.013601f
C813 VTAIL.n29 VSUBS 0.02531f
C814 VTAIL.n30 VSUBS 0.02531f
C815 VTAIL.n31 VSUBS 0.013601f
C816 VTAIL.n32 VSUBS 0.014401f
C817 VTAIL.n33 VSUBS 0.032147f
C818 VTAIL.n34 VSUBS 0.032147f
C819 VTAIL.n35 VSUBS 0.032147f
C820 VTAIL.n36 VSUBS 0.014401f
C821 VTAIL.n37 VSUBS 0.013601f
C822 VTAIL.n38 VSUBS 0.02531f
C823 VTAIL.n39 VSUBS 0.02531f
C824 VTAIL.n40 VSUBS 0.013601f
C825 VTAIL.n41 VSUBS 0.014001f
C826 VTAIL.n42 VSUBS 0.014001f
C827 VTAIL.n43 VSUBS 0.032147f
C828 VTAIL.n44 VSUBS 0.032147f
C829 VTAIL.n45 VSUBS 0.014401f
C830 VTAIL.n46 VSUBS 0.013601f
C831 VTAIL.n47 VSUBS 0.02531f
C832 VTAIL.n48 VSUBS 0.02531f
C833 VTAIL.n49 VSUBS 0.013601f
C834 VTAIL.n50 VSUBS 0.014401f
C835 VTAIL.n51 VSUBS 0.032147f
C836 VTAIL.n52 VSUBS 0.072712f
C837 VTAIL.n53 VSUBS 0.014401f
C838 VTAIL.n54 VSUBS 0.013601f
C839 VTAIL.n55 VSUBS 0.056774f
C840 VTAIL.n56 VSUBS 0.036286f
C841 VTAIL.n57 VSUBS 0.21451f
C842 VTAIL.n58 VSUBS 0.02631f
C843 VTAIL.n59 VSUBS 0.02531f
C844 VTAIL.n60 VSUBS 0.013601f
C845 VTAIL.n61 VSUBS 0.032147f
C846 VTAIL.n62 VSUBS 0.014401f
C847 VTAIL.n63 VSUBS 0.02531f
C848 VTAIL.n64 VSUBS 0.013601f
C849 VTAIL.n65 VSUBS 0.032147f
C850 VTAIL.n66 VSUBS 0.014401f
C851 VTAIL.n67 VSUBS 0.02531f
C852 VTAIL.n68 VSUBS 0.013601f
C853 VTAIL.n69 VSUBS 0.032147f
C854 VTAIL.n70 VSUBS 0.014401f
C855 VTAIL.n71 VSUBS 0.02531f
C856 VTAIL.n72 VSUBS 0.013601f
C857 VTAIL.n73 VSUBS 0.032147f
C858 VTAIL.n74 VSUBS 0.014401f
C859 VTAIL.n75 VSUBS 0.183659f
C860 VTAIL.t4 VSUBS 0.069162f
C861 VTAIL.n76 VSUBS 0.02411f
C862 VTAIL.n77 VSUBS 0.024183f
C863 VTAIL.n78 VSUBS 0.013601f
C864 VTAIL.n79 VSUBS 1.09162f
C865 VTAIL.n80 VSUBS 0.02531f
C866 VTAIL.n81 VSUBS 0.013601f
C867 VTAIL.n82 VSUBS 0.014401f
C868 VTAIL.n83 VSUBS 0.032147f
C869 VTAIL.n84 VSUBS 0.032147f
C870 VTAIL.n85 VSUBS 0.014401f
C871 VTAIL.n86 VSUBS 0.013601f
C872 VTAIL.n87 VSUBS 0.02531f
C873 VTAIL.n88 VSUBS 0.02531f
C874 VTAIL.n89 VSUBS 0.013601f
C875 VTAIL.n90 VSUBS 0.014401f
C876 VTAIL.n91 VSUBS 0.032147f
C877 VTAIL.n92 VSUBS 0.032147f
C878 VTAIL.n93 VSUBS 0.032147f
C879 VTAIL.n94 VSUBS 0.014401f
C880 VTAIL.n95 VSUBS 0.013601f
C881 VTAIL.n96 VSUBS 0.02531f
C882 VTAIL.n97 VSUBS 0.02531f
C883 VTAIL.n98 VSUBS 0.013601f
C884 VTAIL.n99 VSUBS 0.014001f
C885 VTAIL.n100 VSUBS 0.014001f
C886 VTAIL.n101 VSUBS 0.032147f
C887 VTAIL.n102 VSUBS 0.032147f
C888 VTAIL.n103 VSUBS 0.014401f
C889 VTAIL.n104 VSUBS 0.013601f
C890 VTAIL.n105 VSUBS 0.02531f
C891 VTAIL.n106 VSUBS 0.02531f
C892 VTAIL.n107 VSUBS 0.013601f
C893 VTAIL.n108 VSUBS 0.014401f
C894 VTAIL.n109 VSUBS 0.032147f
C895 VTAIL.n110 VSUBS 0.072712f
C896 VTAIL.n111 VSUBS 0.014401f
C897 VTAIL.n112 VSUBS 0.013601f
C898 VTAIL.n113 VSUBS 0.056774f
C899 VTAIL.n114 VSUBS 0.036286f
C900 VTAIL.n115 VSUBS 0.36057f
C901 VTAIL.n116 VSUBS 0.02631f
C902 VTAIL.n117 VSUBS 0.02531f
C903 VTAIL.n118 VSUBS 0.013601f
C904 VTAIL.n119 VSUBS 0.032147f
C905 VTAIL.n120 VSUBS 0.014401f
C906 VTAIL.n121 VSUBS 0.02531f
C907 VTAIL.n122 VSUBS 0.013601f
C908 VTAIL.n123 VSUBS 0.032147f
C909 VTAIL.n124 VSUBS 0.014401f
C910 VTAIL.n125 VSUBS 0.02531f
C911 VTAIL.n126 VSUBS 0.013601f
C912 VTAIL.n127 VSUBS 0.032147f
C913 VTAIL.n128 VSUBS 0.014401f
C914 VTAIL.n129 VSUBS 0.02531f
C915 VTAIL.n130 VSUBS 0.013601f
C916 VTAIL.n131 VSUBS 0.032147f
C917 VTAIL.n132 VSUBS 0.014401f
C918 VTAIL.n133 VSUBS 0.183659f
C919 VTAIL.t5 VSUBS 0.069162f
C920 VTAIL.n134 VSUBS 0.02411f
C921 VTAIL.n135 VSUBS 0.024183f
C922 VTAIL.n136 VSUBS 0.013601f
C923 VTAIL.n137 VSUBS 1.09162f
C924 VTAIL.n138 VSUBS 0.02531f
C925 VTAIL.n139 VSUBS 0.013601f
C926 VTAIL.n140 VSUBS 0.014401f
C927 VTAIL.n141 VSUBS 0.032147f
C928 VTAIL.n142 VSUBS 0.032147f
C929 VTAIL.n143 VSUBS 0.014401f
C930 VTAIL.n144 VSUBS 0.013601f
C931 VTAIL.n145 VSUBS 0.02531f
C932 VTAIL.n146 VSUBS 0.02531f
C933 VTAIL.n147 VSUBS 0.013601f
C934 VTAIL.n148 VSUBS 0.014401f
C935 VTAIL.n149 VSUBS 0.032147f
C936 VTAIL.n150 VSUBS 0.032147f
C937 VTAIL.n151 VSUBS 0.032147f
C938 VTAIL.n152 VSUBS 0.014401f
C939 VTAIL.n153 VSUBS 0.013601f
C940 VTAIL.n154 VSUBS 0.02531f
C941 VTAIL.n155 VSUBS 0.02531f
C942 VTAIL.n156 VSUBS 0.013601f
C943 VTAIL.n157 VSUBS 0.014001f
C944 VTAIL.n158 VSUBS 0.014001f
C945 VTAIL.n159 VSUBS 0.032147f
C946 VTAIL.n160 VSUBS 0.032147f
C947 VTAIL.n161 VSUBS 0.014401f
C948 VTAIL.n162 VSUBS 0.013601f
C949 VTAIL.n163 VSUBS 0.02531f
C950 VTAIL.n164 VSUBS 0.02531f
C951 VTAIL.n165 VSUBS 0.013601f
C952 VTAIL.n166 VSUBS 0.014401f
C953 VTAIL.n167 VSUBS 0.032147f
C954 VTAIL.n168 VSUBS 0.072712f
C955 VTAIL.n169 VSUBS 0.014401f
C956 VTAIL.n170 VSUBS 0.013601f
C957 VTAIL.n171 VSUBS 0.056774f
C958 VTAIL.n172 VSUBS 0.036286f
C959 VTAIL.n173 VSUBS 1.71502f
C960 VTAIL.n174 VSUBS 0.02631f
C961 VTAIL.n175 VSUBS 0.02531f
C962 VTAIL.n176 VSUBS 0.013601f
C963 VTAIL.n177 VSUBS 0.032147f
C964 VTAIL.n178 VSUBS 0.014401f
C965 VTAIL.n179 VSUBS 0.02531f
C966 VTAIL.n180 VSUBS 0.013601f
C967 VTAIL.n181 VSUBS 0.032147f
C968 VTAIL.n182 VSUBS 0.014401f
C969 VTAIL.n183 VSUBS 0.02531f
C970 VTAIL.n184 VSUBS 0.013601f
C971 VTAIL.n185 VSUBS 0.032147f
C972 VTAIL.n186 VSUBS 0.032147f
C973 VTAIL.n187 VSUBS 0.014401f
C974 VTAIL.n188 VSUBS 0.02531f
C975 VTAIL.n189 VSUBS 0.013601f
C976 VTAIL.n190 VSUBS 0.032147f
C977 VTAIL.n191 VSUBS 0.014401f
C978 VTAIL.n192 VSUBS 0.183659f
C979 VTAIL.t2 VSUBS 0.069162f
C980 VTAIL.n193 VSUBS 0.02411f
C981 VTAIL.n194 VSUBS 0.024183f
C982 VTAIL.n195 VSUBS 0.013601f
C983 VTAIL.n196 VSUBS 1.09162f
C984 VTAIL.n197 VSUBS 0.02531f
C985 VTAIL.n198 VSUBS 0.013601f
C986 VTAIL.n199 VSUBS 0.014401f
C987 VTAIL.n200 VSUBS 0.032147f
C988 VTAIL.n201 VSUBS 0.032147f
C989 VTAIL.n202 VSUBS 0.014401f
C990 VTAIL.n203 VSUBS 0.013601f
C991 VTAIL.n204 VSUBS 0.02531f
C992 VTAIL.n205 VSUBS 0.02531f
C993 VTAIL.n206 VSUBS 0.013601f
C994 VTAIL.n207 VSUBS 0.014401f
C995 VTAIL.n208 VSUBS 0.032147f
C996 VTAIL.n209 VSUBS 0.032147f
C997 VTAIL.n210 VSUBS 0.014401f
C998 VTAIL.n211 VSUBS 0.013601f
C999 VTAIL.n212 VSUBS 0.02531f
C1000 VTAIL.n213 VSUBS 0.02531f
C1001 VTAIL.n214 VSUBS 0.013601f
C1002 VTAIL.n215 VSUBS 0.014001f
C1003 VTAIL.n216 VSUBS 0.014001f
C1004 VTAIL.n217 VSUBS 0.032147f
C1005 VTAIL.n218 VSUBS 0.032147f
C1006 VTAIL.n219 VSUBS 0.014401f
C1007 VTAIL.n220 VSUBS 0.013601f
C1008 VTAIL.n221 VSUBS 0.02531f
C1009 VTAIL.n222 VSUBS 0.02531f
C1010 VTAIL.n223 VSUBS 0.013601f
C1011 VTAIL.n224 VSUBS 0.014401f
C1012 VTAIL.n225 VSUBS 0.032147f
C1013 VTAIL.n226 VSUBS 0.072712f
C1014 VTAIL.n227 VSUBS 0.014401f
C1015 VTAIL.n228 VSUBS 0.013601f
C1016 VTAIL.n229 VSUBS 0.056774f
C1017 VTAIL.n230 VSUBS 0.036286f
C1018 VTAIL.n231 VSUBS 1.71502f
C1019 VTAIL.n232 VSUBS 0.02631f
C1020 VTAIL.n233 VSUBS 0.02531f
C1021 VTAIL.n234 VSUBS 0.013601f
C1022 VTAIL.n235 VSUBS 0.032147f
C1023 VTAIL.n236 VSUBS 0.014401f
C1024 VTAIL.n237 VSUBS 0.02531f
C1025 VTAIL.n238 VSUBS 0.013601f
C1026 VTAIL.n239 VSUBS 0.032147f
C1027 VTAIL.n240 VSUBS 0.014401f
C1028 VTAIL.n241 VSUBS 0.02531f
C1029 VTAIL.n242 VSUBS 0.013601f
C1030 VTAIL.n243 VSUBS 0.032147f
C1031 VTAIL.n244 VSUBS 0.032147f
C1032 VTAIL.n245 VSUBS 0.014401f
C1033 VTAIL.n246 VSUBS 0.02531f
C1034 VTAIL.n247 VSUBS 0.013601f
C1035 VTAIL.n248 VSUBS 0.032147f
C1036 VTAIL.n249 VSUBS 0.014401f
C1037 VTAIL.n250 VSUBS 0.183659f
C1038 VTAIL.t7 VSUBS 0.069162f
C1039 VTAIL.n251 VSUBS 0.02411f
C1040 VTAIL.n252 VSUBS 0.024183f
C1041 VTAIL.n253 VSUBS 0.013601f
C1042 VTAIL.n254 VSUBS 1.09162f
C1043 VTAIL.n255 VSUBS 0.02531f
C1044 VTAIL.n256 VSUBS 0.013601f
C1045 VTAIL.n257 VSUBS 0.014401f
C1046 VTAIL.n258 VSUBS 0.032147f
C1047 VTAIL.n259 VSUBS 0.032147f
C1048 VTAIL.n260 VSUBS 0.014401f
C1049 VTAIL.n261 VSUBS 0.013601f
C1050 VTAIL.n262 VSUBS 0.02531f
C1051 VTAIL.n263 VSUBS 0.02531f
C1052 VTAIL.n264 VSUBS 0.013601f
C1053 VTAIL.n265 VSUBS 0.014401f
C1054 VTAIL.n266 VSUBS 0.032147f
C1055 VTAIL.n267 VSUBS 0.032147f
C1056 VTAIL.n268 VSUBS 0.014401f
C1057 VTAIL.n269 VSUBS 0.013601f
C1058 VTAIL.n270 VSUBS 0.02531f
C1059 VTAIL.n271 VSUBS 0.02531f
C1060 VTAIL.n272 VSUBS 0.013601f
C1061 VTAIL.n273 VSUBS 0.014001f
C1062 VTAIL.n274 VSUBS 0.014001f
C1063 VTAIL.n275 VSUBS 0.032147f
C1064 VTAIL.n276 VSUBS 0.032147f
C1065 VTAIL.n277 VSUBS 0.014401f
C1066 VTAIL.n278 VSUBS 0.013601f
C1067 VTAIL.n279 VSUBS 0.02531f
C1068 VTAIL.n280 VSUBS 0.02531f
C1069 VTAIL.n281 VSUBS 0.013601f
C1070 VTAIL.n282 VSUBS 0.014401f
C1071 VTAIL.n283 VSUBS 0.032147f
C1072 VTAIL.n284 VSUBS 0.072712f
C1073 VTAIL.n285 VSUBS 0.014401f
C1074 VTAIL.n286 VSUBS 0.013601f
C1075 VTAIL.n287 VSUBS 0.056774f
C1076 VTAIL.n288 VSUBS 0.036286f
C1077 VTAIL.n289 VSUBS 0.36057f
C1078 VTAIL.n290 VSUBS 0.02631f
C1079 VTAIL.n291 VSUBS 0.02531f
C1080 VTAIL.n292 VSUBS 0.013601f
C1081 VTAIL.n293 VSUBS 0.032147f
C1082 VTAIL.n294 VSUBS 0.014401f
C1083 VTAIL.n295 VSUBS 0.02531f
C1084 VTAIL.n296 VSUBS 0.013601f
C1085 VTAIL.n297 VSUBS 0.032147f
C1086 VTAIL.n298 VSUBS 0.014401f
C1087 VTAIL.n299 VSUBS 0.02531f
C1088 VTAIL.n300 VSUBS 0.013601f
C1089 VTAIL.n301 VSUBS 0.032147f
C1090 VTAIL.n302 VSUBS 0.032147f
C1091 VTAIL.n303 VSUBS 0.014401f
C1092 VTAIL.n304 VSUBS 0.02531f
C1093 VTAIL.n305 VSUBS 0.013601f
C1094 VTAIL.n306 VSUBS 0.032147f
C1095 VTAIL.n307 VSUBS 0.014401f
C1096 VTAIL.n308 VSUBS 0.183659f
C1097 VTAIL.t6 VSUBS 0.069162f
C1098 VTAIL.n309 VSUBS 0.02411f
C1099 VTAIL.n310 VSUBS 0.024183f
C1100 VTAIL.n311 VSUBS 0.013601f
C1101 VTAIL.n312 VSUBS 1.09162f
C1102 VTAIL.n313 VSUBS 0.02531f
C1103 VTAIL.n314 VSUBS 0.013601f
C1104 VTAIL.n315 VSUBS 0.014401f
C1105 VTAIL.n316 VSUBS 0.032147f
C1106 VTAIL.n317 VSUBS 0.032147f
C1107 VTAIL.n318 VSUBS 0.014401f
C1108 VTAIL.n319 VSUBS 0.013601f
C1109 VTAIL.n320 VSUBS 0.02531f
C1110 VTAIL.n321 VSUBS 0.02531f
C1111 VTAIL.n322 VSUBS 0.013601f
C1112 VTAIL.n323 VSUBS 0.014401f
C1113 VTAIL.n324 VSUBS 0.032147f
C1114 VTAIL.n325 VSUBS 0.032147f
C1115 VTAIL.n326 VSUBS 0.014401f
C1116 VTAIL.n327 VSUBS 0.013601f
C1117 VTAIL.n328 VSUBS 0.02531f
C1118 VTAIL.n329 VSUBS 0.02531f
C1119 VTAIL.n330 VSUBS 0.013601f
C1120 VTAIL.n331 VSUBS 0.014001f
C1121 VTAIL.n332 VSUBS 0.014001f
C1122 VTAIL.n333 VSUBS 0.032147f
C1123 VTAIL.n334 VSUBS 0.032147f
C1124 VTAIL.n335 VSUBS 0.014401f
C1125 VTAIL.n336 VSUBS 0.013601f
C1126 VTAIL.n337 VSUBS 0.02531f
C1127 VTAIL.n338 VSUBS 0.02531f
C1128 VTAIL.n339 VSUBS 0.013601f
C1129 VTAIL.n340 VSUBS 0.014401f
C1130 VTAIL.n341 VSUBS 0.032147f
C1131 VTAIL.n342 VSUBS 0.072712f
C1132 VTAIL.n343 VSUBS 0.014401f
C1133 VTAIL.n344 VSUBS 0.013601f
C1134 VTAIL.n345 VSUBS 0.056774f
C1135 VTAIL.n346 VSUBS 0.036286f
C1136 VTAIL.n347 VSUBS 0.36057f
C1137 VTAIL.n348 VSUBS 0.02631f
C1138 VTAIL.n349 VSUBS 0.02531f
C1139 VTAIL.n350 VSUBS 0.013601f
C1140 VTAIL.n351 VSUBS 0.032147f
C1141 VTAIL.n352 VSUBS 0.014401f
C1142 VTAIL.n353 VSUBS 0.02531f
C1143 VTAIL.n354 VSUBS 0.013601f
C1144 VTAIL.n355 VSUBS 0.032147f
C1145 VTAIL.n356 VSUBS 0.014401f
C1146 VTAIL.n357 VSUBS 0.02531f
C1147 VTAIL.n358 VSUBS 0.013601f
C1148 VTAIL.n359 VSUBS 0.032147f
C1149 VTAIL.n360 VSUBS 0.032147f
C1150 VTAIL.n361 VSUBS 0.014401f
C1151 VTAIL.n362 VSUBS 0.02531f
C1152 VTAIL.n363 VSUBS 0.013601f
C1153 VTAIL.n364 VSUBS 0.032147f
C1154 VTAIL.n365 VSUBS 0.014401f
C1155 VTAIL.n366 VSUBS 0.183659f
C1156 VTAIL.t3 VSUBS 0.069162f
C1157 VTAIL.n367 VSUBS 0.02411f
C1158 VTAIL.n368 VSUBS 0.024183f
C1159 VTAIL.n369 VSUBS 0.013601f
C1160 VTAIL.n370 VSUBS 1.09162f
C1161 VTAIL.n371 VSUBS 0.02531f
C1162 VTAIL.n372 VSUBS 0.013601f
C1163 VTAIL.n373 VSUBS 0.014401f
C1164 VTAIL.n374 VSUBS 0.032147f
C1165 VTAIL.n375 VSUBS 0.032147f
C1166 VTAIL.n376 VSUBS 0.014401f
C1167 VTAIL.n377 VSUBS 0.013601f
C1168 VTAIL.n378 VSUBS 0.02531f
C1169 VTAIL.n379 VSUBS 0.02531f
C1170 VTAIL.n380 VSUBS 0.013601f
C1171 VTAIL.n381 VSUBS 0.014401f
C1172 VTAIL.n382 VSUBS 0.032147f
C1173 VTAIL.n383 VSUBS 0.032147f
C1174 VTAIL.n384 VSUBS 0.014401f
C1175 VTAIL.n385 VSUBS 0.013601f
C1176 VTAIL.n386 VSUBS 0.02531f
C1177 VTAIL.n387 VSUBS 0.02531f
C1178 VTAIL.n388 VSUBS 0.013601f
C1179 VTAIL.n389 VSUBS 0.014001f
C1180 VTAIL.n390 VSUBS 0.014001f
C1181 VTAIL.n391 VSUBS 0.032147f
C1182 VTAIL.n392 VSUBS 0.032147f
C1183 VTAIL.n393 VSUBS 0.014401f
C1184 VTAIL.n394 VSUBS 0.013601f
C1185 VTAIL.n395 VSUBS 0.02531f
C1186 VTAIL.n396 VSUBS 0.02531f
C1187 VTAIL.n397 VSUBS 0.013601f
C1188 VTAIL.n398 VSUBS 0.014401f
C1189 VTAIL.n399 VSUBS 0.032147f
C1190 VTAIL.n400 VSUBS 0.072712f
C1191 VTAIL.n401 VSUBS 0.014401f
C1192 VTAIL.n402 VSUBS 0.013601f
C1193 VTAIL.n403 VSUBS 0.056774f
C1194 VTAIL.n404 VSUBS 0.036286f
C1195 VTAIL.n405 VSUBS 1.71502f
C1196 VTAIL.n406 VSUBS 0.02631f
C1197 VTAIL.n407 VSUBS 0.02531f
C1198 VTAIL.n408 VSUBS 0.013601f
C1199 VTAIL.n409 VSUBS 0.032147f
C1200 VTAIL.n410 VSUBS 0.014401f
C1201 VTAIL.n411 VSUBS 0.02531f
C1202 VTAIL.n412 VSUBS 0.013601f
C1203 VTAIL.n413 VSUBS 0.032147f
C1204 VTAIL.n414 VSUBS 0.014401f
C1205 VTAIL.n415 VSUBS 0.02531f
C1206 VTAIL.n416 VSUBS 0.013601f
C1207 VTAIL.n417 VSUBS 0.032147f
C1208 VTAIL.n418 VSUBS 0.014401f
C1209 VTAIL.n419 VSUBS 0.02531f
C1210 VTAIL.n420 VSUBS 0.013601f
C1211 VTAIL.n421 VSUBS 0.032147f
C1212 VTAIL.n422 VSUBS 0.014401f
C1213 VTAIL.n423 VSUBS 0.183659f
C1214 VTAIL.t0 VSUBS 0.069162f
C1215 VTAIL.n424 VSUBS 0.02411f
C1216 VTAIL.n425 VSUBS 0.024183f
C1217 VTAIL.n426 VSUBS 0.013601f
C1218 VTAIL.n427 VSUBS 1.09162f
C1219 VTAIL.n428 VSUBS 0.02531f
C1220 VTAIL.n429 VSUBS 0.013601f
C1221 VTAIL.n430 VSUBS 0.014401f
C1222 VTAIL.n431 VSUBS 0.032147f
C1223 VTAIL.n432 VSUBS 0.032147f
C1224 VTAIL.n433 VSUBS 0.014401f
C1225 VTAIL.n434 VSUBS 0.013601f
C1226 VTAIL.n435 VSUBS 0.02531f
C1227 VTAIL.n436 VSUBS 0.02531f
C1228 VTAIL.n437 VSUBS 0.013601f
C1229 VTAIL.n438 VSUBS 0.014401f
C1230 VTAIL.n439 VSUBS 0.032147f
C1231 VTAIL.n440 VSUBS 0.032147f
C1232 VTAIL.n441 VSUBS 0.032147f
C1233 VTAIL.n442 VSUBS 0.014401f
C1234 VTAIL.n443 VSUBS 0.013601f
C1235 VTAIL.n444 VSUBS 0.02531f
C1236 VTAIL.n445 VSUBS 0.02531f
C1237 VTAIL.n446 VSUBS 0.013601f
C1238 VTAIL.n447 VSUBS 0.014001f
C1239 VTAIL.n448 VSUBS 0.014001f
C1240 VTAIL.n449 VSUBS 0.032147f
C1241 VTAIL.n450 VSUBS 0.032147f
C1242 VTAIL.n451 VSUBS 0.014401f
C1243 VTAIL.n452 VSUBS 0.013601f
C1244 VTAIL.n453 VSUBS 0.02531f
C1245 VTAIL.n454 VSUBS 0.02531f
C1246 VTAIL.n455 VSUBS 0.013601f
C1247 VTAIL.n456 VSUBS 0.014401f
C1248 VTAIL.n457 VSUBS 0.032147f
C1249 VTAIL.n458 VSUBS 0.072712f
C1250 VTAIL.n459 VSUBS 0.014401f
C1251 VTAIL.n460 VSUBS 0.013601f
C1252 VTAIL.n461 VSUBS 0.056774f
C1253 VTAIL.n462 VSUBS 0.036286f
C1254 VTAIL.n463 VSUBS 1.55947f
C1255 VP.n0 VSUBS 0.058406f
C1256 VP.t0 VSUBS 3.54814f
C1257 VP.n1 VSUBS 0.05787f
C1258 VP.n2 VSUBS 0.031051f
C1259 VP.n3 VSUBS 0.05787f
C1260 VP.t1 VSUBS 4.04469f
C1261 VP.t2 VSUBS 4.06569f
C1262 VP.n4 VSUBS 4.42039f
C1263 VP.n5 VSUBS 1.88608f
C1264 VP.t3 VSUBS 3.54814f
C1265 VP.n6 VSUBS 1.38348f
C1266 VP.n7 VSUBS 0.051869f
C1267 VP.n8 VSUBS 0.058406f
C1268 VP.n9 VSUBS 0.031051f
C1269 VP.n10 VSUBS 0.031051f
C1270 VP.n11 VSUBS 0.05787f
C1271 VP.n12 VSUBS 0.045328f
C1272 VP.n13 VSUBS 0.045328f
C1273 VP.n14 VSUBS 0.031051f
C1274 VP.n15 VSUBS 0.031051f
C1275 VP.n16 VSUBS 0.031051f
C1276 VP.n17 VSUBS 0.05787f
C1277 VP.n18 VSUBS 0.051869f
C1278 VP.n19 VSUBS 1.38348f
C1279 VP.n20 VSUBS 0.100299f
.ends

