* NGSPICE file created from diff_pair_sample_0998.ext - technology: sky130A

.subckt diff_pair_sample_0998 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=0 ps=0 w=12.85 l=2.65
X1 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=0 ps=0 w=12.85 l=2.65
X2 VTAIL.t15 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X3 VDD2.t7 VN.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X4 VTAIL.t2 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X5 VDD1.t4 VP.t1 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=5.0115 ps=26.48 w=12.85 l=2.65
X6 VTAIL.t13 VP.t2 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=2.12025 ps=13.18 w=12.85 l=2.65
X7 VTAIL.t12 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X8 VTAIL.t5 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=2.12025 ps=13.18 w=12.85 l=2.65
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=0 ps=0 w=12.85 l=2.65
X10 VTAIL.t11 VP.t4 VDD1.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=2.12025 ps=13.18 w=12.85 l=2.65
X11 VTAIL.t6 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=2.12025 ps=13.18 w=12.85 l=2.65
X12 VDD1.t6 VP.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=5.0115 ps=26.48 w=12.85 l=2.65
X13 VDD1.t5 VP.t6 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X14 VDD2.t3 VN.t4 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=5.0115 ps=26.48 w=12.85 l=2.65
X15 VDD2.t2 VN.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=5.0115 ps=26.48 w=12.85 l=2.65
X16 VDD1.t2 VP.t7 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X17 VDD2.t1 VN.t6 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X18 VTAIL.t0 VN.t7 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.12025 pd=13.18 as=2.12025 ps=13.18 w=12.85 l=2.65
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0115 pd=26.48 as=0 ps=0 w=12.85 l=2.65
R0 B.n918 B.n917 585
R1 B.n342 B.n145 585
R2 B.n341 B.n340 585
R3 B.n339 B.n338 585
R4 B.n337 B.n336 585
R5 B.n335 B.n334 585
R6 B.n333 B.n332 585
R7 B.n331 B.n330 585
R8 B.n329 B.n328 585
R9 B.n327 B.n326 585
R10 B.n325 B.n324 585
R11 B.n323 B.n322 585
R12 B.n321 B.n320 585
R13 B.n319 B.n318 585
R14 B.n317 B.n316 585
R15 B.n315 B.n314 585
R16 B.n313 B.n312 585
R17 B.n311 B.n310 585
R18 B.n309 B.n308 585
R19 B.n307 B.n306 585
R20 B.n305 B.n304 585
R21 B.n303 B.n302 585
R22 B.n301 B.n300 585
R23 B.n299 B.n298 585
R24 B.n297 B.n296 585
R25 B.n295 B.n294 585
R26 B.n293 B.n292 585
R27 B.n291 B.n290 585
R28 B.n289 B.n288 585
R29 B.n287 B.n286 585
R30 B.n285 B.n284 585
R31 B.n283 B.n282 585
R32 B.n281 B.n280 585
R33 B.n279 B.n278 585
R34 B.n277 B.n276 585
R35 B.n275 B.n274 585
R36 B.n273 B.n272 585
R37 B.n271 B.n270 585
R38 B.n269 B.n268 585
R39 B.n267 B.n266 585
R40 B.n265 B.n264 585
R41 B.n263 B.n262 585
R42 B.n261 B.n260 585
R43 B.n259 B.n258 585
R44 B.n257 B.n256 585
R45 B.n255 B.n254 585
R46 B.n253 B.n252 585
R47 B.n251 B.n250 585
R48 B.n249 B.n248 585
R49 B.n247 B.n246 585
R50 B.n245 B.n244 585
R51 B.n243 B.n242 585
R52 B.n241 B.n240 585
R53 B.n239 B.n238 585
R54 B.n237 B.n236 585
R55 B.n235 B.n234 585
R56 B.n233 B.n232 585
R57 B.n231 B.n230 585
R58 B.n229 B.n228 585
R59 B.n227 B.n226 585
R60 B.n225 B.n224 585
R61 B.n223 B.n222 585
R62 B.n221 B.n220 585
R63 B.n219 B.n218 585
R64 B.n217 B.n216 585
R65 B.n215 B.n214 585
R66 B.n213 B.n212 585
R67 B.n211 B.n210 585
R68 B.n209 B.n208 585
R69 B.n207 B.n206 585
R70 B.n205 B.n204 585
R71 B.n203 B.n202 585
R72 B.n201 B.n200 585
R73 B.n199 B.n198 585
R74 B.n197 B.n196 585
R75 B.n195 B.n194 585
R76 B.n193 B.n192 585
R77 B.n191 B.n190 585
R78 B.n189 B.n188 585
R79 B.n187 B.n186 585
R80 B.n185 B.n184 585
R81 B.n183 B.n182 585
R82 B.n181 B.n180 585
R83 B.n179 B.n178 585
R84 B.n177 B.n176 585
R85 B.n175 B.n174 585
R86 B.n173 B.n172 585
R87 B.n171 B.n170 585
R88 B.n169 B.n168 585
R89 B.n167 B.n166 585
R90 B.n165 B.n164 585
R91 B.n163 B.n162 585
R92 B.n161 B.n160 585
R93 B.n159 B.n158 585
R94 B.n157 B.n156 585
R95 B.n155 B.n154 585
R96 B.n153 B.n152 585
R97 B.n95 B.n94 585
R98 B.n916 B.n96 585
R99 B.n921 B.n96 585
R100 B.n915 B.n914 585
R101 B.n914 B.n92 585
R102 B.n913 B.n91 585
R103 B.n927 B.n91 585
R104 B.n912 B.n90 585
R105 B.n928 B.n90 585
R106 B.n911 B.n89 585
R107 B.n929 B.n89 585
R108 B.n910 B.n909 585
R109 B.n909 B.n85 585
R110 B.n908 B.n84 585
R111 B.n935 B.n84 585
R112 B.n907 B.n83 585
R113 B.n936 B.n83 585
R114 B.n906 B.n82 585
R115 B.n937 B.n82 585
R116 B.n905 B.n904 585
R117 B.n904 B.n78 585
R118 B.n903 B.n77 585
R119 B.n943 B.n77 585
R120 B.n902 B.n76 585
R121 B.n944 B.n76 585
R122 B.n901 B.n75 585
R123 B.n945 B.n75 585
R124 B.n900 B.n899 585
R125 B.n899 B.n71 585
R126 B.n898 B.n70 585
R127 B.n951 B.n70 585
R128 B.n897 B.n69 585
R129 B.n952 B.n69 585
R130 B.n896 B.n68 585
R131 B.n953 B.n68 585
R132 B.n895 B.n894 585
R133 B.n894 B.n64 585
R134 B.n893 B.n63 585
R135 B.n959 B.n63 585
R136 B.n892 B.n62 585
R137 B.n960 B.n62 585
R138 B.n891 B.n61 585
R139 B.n961 B.n61 585
R140 B.n890 B.n889 585
R141 B.n889 B.n57 585
R142 B.n888 B.n56 585
R143 B.n967 B.n56 585
R144 B.n887 B.n55 585
R145 B.n968 B.n55 585
R146 B.n886 B.n54 585
R147 B.n969 B.n54 585
R148 B.n885 B.n884 585
R149 B.n884 B.n50 585
R150 B.n883 B.n49 585
R151 B.n975 B.n49 585
R152 B.n882 B.n48 585
R153 B.n976 B.n48 585
R154 B.n881 B.n47 585
R155 B.n977 B.n47 585
R156 B.n880 B.n879 585
R157 B.n879 B.n43 585
R158 B.n878 B.n42 585
R159 B.n983 B.n42 585
R160 B.n877 B.n41 585
R161 B.n984 B.n41 585
R162 B.n876 B.n40 585
R163 B.n985 B.n40 585
R164 B.n875 B.n874 585
R165 B.n874 B.n36 585
R166 B.n873 B.n35 585
R167 B.n991 B.n35 585
R168 B.n872 B.n34 585
R169 B.n992 B.n34 585
R170 B.n871 B.n33 585
R171 B.n993 B.n33 585
R172 B.n870 B.n869 585
R173 B.n869 B.n32 585
R174 B.n868 B.n28 585
R175 B.n999 B.n28 585
R176 B.n867 B.n27 585
R177 B.n1000 B.n27 585
R178 B.n866 B.n26 585
R179 B.n1001 B.n26 585
R180 B.n865 B.n864 585
R181 B.n864 B.n22 585
R182 B.n863 B.n21 585
R183 B.n1007 B.n21 585
R184 B.n862 B.n20 585
R185 B.n1008 B.n20 585
R186 B.n861 B.n19 585
R187 B.n1009 B.n19 585
R188 B.n860 B.n859 585
R189 B.n859 B.n15 585
R190 B.n858 B.n14 585
R191 B.n1015 B.n14 585
R192 B.n857 B.n13 585
R193 B.n1016 B.n13 585
R194 B.n856 B.n12 585
R195 B.n1017 B.n12 585
R196 B.n855 B.n854 585
R197 B.n854 B.n8 585
R198 B.n853 B.n7 585
R199 B.n1023 B.n7 585
R200 B.n852 B.n6 585
R201 B.n1024 B.n6 585
R202 B.n851 B.n5 585
R203 B.n1025 B.n5 585
R204 B.n850 B.n849 585
R205 B.n849 B.n4 585
R206 B.n848 B.n343 585
R207 B.n848 B.n847 585
R208 B.n838 B.n344 585
R209 B.n345 B.n344 585
R210 B.n840 B.n839 585
R211 B.n841 B.n840 585
R212 B.n837 B.n350 585
R213 B.n350 B.n349 585
R214 B.n836 B.n835 585
R215 B.n835 B.n834 585
R216 B.n352 B.n351 585
R217 B.n353 B.n352 585
R218 B.n827 B.n826 585
R219 B.n828 B.n827 585
R220 B.n825 B.n358 585
R221 B.n358 B.n357 585
R222 B.n824 B.n823 585
R223 B.n823 B.n822 585
R224 B.n360 B.n359 585
R225 B.n361 B.n360 585
R226 B.n815 B.n814 585
R227 B.n816 B.n815 585
R228 B.n813 B.n366 585
R229 B.n366 B.n365 585
R230 B.n812 B.n811 585
R231 B.n811 B.n810 585
R232 B.n368 B.n367 585
R233 B.n803 B.n368 585
R234 B.n802 B.n801 585
R235 B.n804 B.n802 585
R236 B.n800 B.n373 585
R237 B.n373 B.n372 585
R238 B.n799 B.n798 585
R239 B.n798 B.n797 585
R240 B.n375 B.n374 585
R241 B.n376 B.n375 585
R242 B.n790 B.n789 585
R243 B.n791 B.n790 585
R244 B.n788 B.n381 585
R245 B.n381 B.n380 585
R246 B.n787 B.n786 585
R247 B.n786 B.n785 585
R248 B.n383 B.n382 585
R249 B.n384 B.n383 585
R250 B.n778 B.n777 585
R251 B.n779 B.n778 585
R252 B.n776 B.n389 585
R253 B.n389 B.n388 585
R254 B.n775 B.n774 585
R255 B.n774 B.n773 585
R256 B.n391 B.n390 585
R257 B.n392 B.n391 585
R258 B.n766 B.n765 585
R259 B.n767 B.n766 585
R260 B.n764 B.n397 585
R261 B.n397 B.n396 585
R262 B.n763 B.n762 585
R263 B.n762 B.n761 585
R264 B.n399 B.n398 585
R265 B.n400 B.n399 585
R266 B.n754 B.n753 585
R267 B.n755 B.n754 585
R268 B.n752 B.n404 585
R269 B.n408 B.n404 585
R270 B.n751 B.n750 585
R271 B.n750 B.n749 585
R272 B.n406 B.n405 585
R273 B.n407 B.n406 585
R274 B.n742 B.n741 585
R275 B.n743 B.n742 585
R276 B.n740 B.n413 585
R277 B.n413 B.n412 585
R278 B.n739 B.n738 585
R279 B.n738 B.n737 585
R280 B.n415 B.n414 585
R281 B.n416 B.n415 585
R282 B.n730 B.n729 585
R283 B.n731 B.n730 585
R284 B.n728 B.n421 585
R285 B.n421 B.n420 585
R286 B.n727 B.n726 585
R287 B.n726 B.n725 585
R288 B.n423 B.n422 585
R289 B.n424 B.n423 585
R290 B.n718 B.n717 585
R291 B.n719 B.n718 585
R292 B.n716 B.n428 585
R293 B.n432 B.n428 585
R294 B.n715 B.n714 585
R295 B.n714 B.n713 585
R296 B.n430 B.n429 585
R297 B.n431 B.n430 585
R298 B.n706 B.n705 585
R299 B.n707 B.n706 585
R300 B.n704 B.n437 585
R301 B.n437 B.n436 585
R302 B.n703 B.n702 585
R303 B.n702 B.n701 585
R304 B.n439 B.n438 585
R305 B.n440 B.n439 585
R306 B.n694 B.n693 585
R307 B.n695 B.n694 585
R308 B.n443 B.n442 585
R309 B.n498 B.n496 585
R310 B.n499 B.n495 585
R311 B.n499 B.n444 585
R312 B.n502 B.n501 585
R313 B.n503 B.n494 585
R314 B.n505 B.n504 585
R315 B.n507 B.n493 585
R316 B.n510 B.n509 585
R317 B.n511 B.n492 585
R318 B.n513 B.n512 585
R319 B.n515 B.n491 585
R320 B.n518 B.n517 585
R321 B.n519 B.n490 585
R322 B.n521 B.n520 585
R323 B.n523 B.n489 585
R324 B.n526 B.n525 585
R325 B.n527 B.n488 585
R326 B.n529 B.n528 585
R327 B.n531 B.n487 585
R328 B.n534 B.n533 585
R329 B.n535 B.n486 585
R330 B.n537 B.n536 585
R331 B.n539 B.n485 585
R332 B.n542 B.n541 585
R333 B.n543 B.n484 585
R334 B.n545 B.n544 585
R335 B.n547 B.n483 585
R336 B.n550 B.n549 585
R337 B.n551 B.n482 585
R338 B.n553 B.n552 585
R339 B.n555 B.n481 585
R340 B.n558 B.n557 585
R341 B.n559 B.n480 585
R342 B.n561 B.n560 585
R343 B.n563 B.n479 585
R344 B.n566 B.n565 585
R345 B.n567 B.n478 585
R346 B.n569 B.n568 585
R347 B.n571 B.n477 585
R348 B.n574 B.n573 585
R349 B.n575 B.n476 585
R350 B.n577 B.n576 585
R351 B.n579 B.n475 585
R352 B.n582 B.n581 585
R353 B.n584 B.n472 585
R354 B.n586 B.n585 585
R355 B.n588 B.n471 585
R356 B.n591 B.n590 585
R357 B.n592 B.n470 585
R358 B.n594 B.n593 585
R359 B.n596 B.n469 585
R360 B.n599 B.n598 585
R361 B.n600 B.n468 585
R362 B.n605 B.n604 585
R363 B.n607 B.n467 585
R364 B.n610 B.n609 585
R365 B.n611 B.n466 585
R366 B.n613 B.n612 585
R367 B.n615 B.n465 585
R368 B.n618 B.n617 585
R369 B.n619 B.n464 585
R370 B.n621 B.n620 585
R371 B.n623 B.n463 585
R372 B.n626 B.n625 585
R373 B.n627 B.n462 585
R374 B.n629 B.n628 585
R375 B.n631 B.n461 585
R376 B.n634 B.n633 585
R377 B.n635 B.n460 585
R378 B.n637 B.n636 585
R379 B.n639 B.n459 585
R380 B.n642 B.n641 585
R381 B.n643 B.n458 585
R382 B.n645 B.n644 585
R383 B.n647 B.n457 585
R384 B.n650 B.n649 585
R385 B.n651 B.n456 585
R386 B.n653 B.n652 585
R387 B.n655 B.n455 585
R388 B.n658 B.n657 585
R389 B.n659 B.n454 585
R390 B.n661 B.n660 585
R391 B.n663 B.n453 585
R392 B.n666 B.n665 585
R393 B.n667 B.n452 585
R394 B.n669 B.n668 585
R395 B.n671 B.n451 585
R396 B.n674 B.n673 585
R397 B.n675 B.n450 585
R398 B.n677 B.n676 585
R399 B.n679 B.n449 585
R400 B.n682 B.n681 585
R401 B.n683 B.n448 585
R402 B.n685 B.n684 585
R403 B.n687 B.n447 585
R404 B.n688 B.n446 585
R405 B.n691 B.n690 585
R406 B.n692 B.n445 585
R407 B.n445 B.n444 585
R408 B.n697 B.n696 585
R409 B.n696 B.n695 585
R410 B.n698 B.n441 585
R411 B.n441 B.n440 585
R412 B.n700 B.n699 585
R413 B.n701 B.n700 585
R414 B.n435 B.n434 585
R415 B.n436 B.n435 585
R416 B.n709 B.n708 585
R417 B.n708 B.n707 585
R418 B.n710 B.n433 585
R419 B.n433 B.n431 585
R420 B.n712 B.n711 585
R421 B.n713 B.n712 585
R422 B.n427 B.n426 585
R423 B.n432 B.n427 585
R424 B.n721 B.n720 585
R425 B.n720 B.n719 585
R426 B.n722 B.n425 585
R427 B.n425 B.n424 585
R428 B.n724 B.n723 585
R429 B.n725 B.n724 585
R430 B.n419 B.n418 585
R431 B.n420 B.n419 585
R432 B.n733 B.n732 585
R433 B.n732 B.n731 585
R434 B.n734 B.n417 585
R435 B.n417 B.n416 585
R436 B.n736 B.n735 585
R437 B.n737 B.n736 585
R438 B.n411 B.n410 585
R439 B.n412 B.n411 585
R440 B.n745 B.n744 585
R441 B.n744 B.n743 585
R442 B.n746 B.n409 585
R443 B.n409 B.n407 585
R444 B.n748 B.n747 585
R445 B.n749 B.n748 585
R446 B.n403 B.n402 585
R447 B.n408 B.n403 585
R448 B.n757 B.n756 585
R449 B.n756 B.n755 585
R450 B.n758 B.n401 585
R451 B.n401 B.n400 585
R452 B.n760 B.n759 585
R453 B.n761 B.n760 585
R454 B.n395 B.n394 585
R455 B.n396 B.n395 585
R456 B.n769 B.n768 585
R457 B.n768 B.n767 585
R458 B.n770 B.n393 585
R459 B.n393 B.n392 585
R460 B.n772 B.n771 585
R461 B.n773 B.n772 585
R462 B.n387 B.n386 585
R463 B.n388 B.n387 585
R464 B.n781 B.n780 585
R465 B.n780 B.n779 585
R466 B.n782 B.n385 585
R467 B.n385 B.n384 585
R468 B.n784 B.n783 585
R469 B.n785 B.n784 585
R470 B.n379 B.n378 585
R471 B.n380 B.n379 585
R472 B.n793 B.n792 585
R473 B.n792 B.n791 585
R474 B.n794 B.n377 585
R475 B.n377 B.n376 585
R476 B.n796 B.n795 585
R477 B.n797 B.n796 585
R478 B.n371 B.n370 585
R479 B.n372 B.n371 585
R480 B.n806 B.n805 585
R481 B.n805 B.n804 585
R482 B.n807 B.n369 585
R483 B.n803 B.n369 585
R484 B.n809 B.n808 585
R485 B.n810 B.n809 585
R486 B.n364 B.n363 585
R487 B.n365 B.n364 585
R488 B.n818 B.n817 585
R489 B.n817 B.n816 585
R490 B.n819 B.n362 585
R491 B.n362 B.n361 585
R492 B.n821 B.n820 585
R493 B.n822 B.n821 585
R494 B.n356 B.n355 585
R495 B.n357 B.n356 585
R496 B.n830 B.n829 585
R497 B.n829 B.n828 585
R498 B.n831 B.n354 585
R499 B.n354 B.n353 585
R500 B.n833 B.n832 585
R501 B.n834 B.n833 585
R502 B.n348 B.n347 585
R503 B.n349 B.n348 585
R504 B.n843 B.n842 585
R505 B.n842 B.n841 585
R506 B.n844 B.n346 585
R507 B.n346 B.n345 585
R508 B.n846 B.n845 585
R509 B.n847 B.n846 585
R510 B.n2 B.n0 585
R511 B.n4 B.n2 585
R512 B.n3 B.n1 585
R513 B.n1024 B.n3 585
R514 B.n1022 B.n1021 585
R515 B.n1023 B.n1022 585
R516 B.n1020 B.n9 585
R517 B.n9 B.n8 585
R518 B.n1019 B.n1018 585
R519 B.n1018 B.n1017 585
R520 B.n11 B.n10 585
R521 B.n1016 B.n11 585
R522 B.n1014 B.n1013 585
R523 B.n1015 B.n1014 585
R524 B.n1012 B.n16 585
R525 B.n16 B.n15 585
R526 B.n1011 B.n1010 585
R527 B.n1010 B.n1009 585
R528 B.n18 B.n17 585
R529 B.n1008 B.n18 585
R530 B.n1006 B.n1005 585
R531 B.n1007 B.n1006 585
R532 B.n1004 B.n23 585
R533 B.n23 B.n22 585
R534 B.n1003 B.n1002 585
R535 B.n1002 B.n1001 585
R536 B.n25 B.n24 585
R537 B.n1000 B.n25 585
R538 B.n998 B.n997 585
R539 B.n999 B.n998 585
R540 B.n996 B.n29 585
R541 B.n32 B.n29 585
R542 B.n995 B.n994 585
R543 B.n994 B.n993 585
R544 B.n31 B.n30 585
R545 B.n992 B.n31 585
R546 B.n990 B.n989 585
R547 B.n991 B.n990 585
R548 B.n988 B.n37 585
R549 B.n37 B.n36 585
R550 B.n987 B.n986 585
R551 B.n986 B.n985 585
R552 B.n39 B.n38 585
R553 B.n984 B.n39 585
R554 B.n982 B.n981 585
R555 B.n983 B.n982 585
R556 B.n980 B.n44 585
R557 B.n44 B.n43 585
R558 B.n979 B.n978 585
R559 B.n978 B.n977 585
R560 B.n46 B.n45 585
R561 B.n976 B.n46 585
R562 B.n974 B.n973 585
R563 B.n975 B.n974 585
R564 B.n972 B.n51 585
R565 B.n51 B.n50 585
R566 B.n971 B.n970 585
R567 B.n970 B.n969 585
R568 B.n53 B.n52 585
R569 B.n968 B.n53 585
R570 B.n966 B.n965 585
R571 B.n967 B.n966 585
R572 B.n964 B.n58 585
R573 B.n58 B.n57 585
R574 B.n963 B.n962 585
R575 B.n962 B.n961 585
R576 B.n60 B.n59 585
R577 B.n960 B.n60 585
R578 B.n958 B.n957 585
R579 B.n959 B.n958 585
R580 B.n956 B.n65 585
R581 B.n65 B.n64 585
R582 B.n955 B.n954 585
R583 B.n954 B.n953 585
R584 B.n67 B.n66 585
R585 B.n952 B.n67 585
R586 B.n950 B.n949 585
R587 B.n951 B.n950 585
R588 B.n948 B.n72 585
R589 B.n72 B.n71 585
R590 B.n947 B.n946 585
R591 B.n946 B.n945 585
R592 B.n74 B.n73 585
R593 B.n944 B.n74 585
R594 B.n942 B.n941 585
R595 B.n943 B.n942 585
R596 B.n940 B.n79 585
R597 B.n79 B.n78 585
R598 B.n939 B.n938 585
R599 B.n938 B.n937 585
R600 B.n81 B.n80 585
R601 B.n936 B.n81 585
R602 B.n934 B.n933 585
R603 B.n935 B.n934 585
R604 B.n932 B.n86 585
R605 B.n86 B.n85 585
R606 B.n931 B.n930 585
R607 B.n930 B.n929 585
R608 B.n88 B.n87 585
R609 B.n928 B.n88 585
R610 B.n926 B.n925 585
R611 B.n927 B.n926 585
R612 B.n924 B.n93 585
R613 B.n93 B.n92 585
R614 B.n923 B.n922 585
R615 B.n922 B.n921 585
R616 B.n1027 B.n1026 585
R617 B.n1026 B.n1025 585
R618 B.n696 B.n443 473.281
R619 B.n922 B.n95 473.281
R620 B.n694 B.n445 473.281
R621 B.n918 B.n96 473.281
R622 B.n601 B.t11 354.812
R623 B.n146 B.t17 354.812
R624 B.n473 B.t21 354.812
R625 B.n149 B.t14 354.812
R626 B.n601 B.t8 324.983
R627 B.n473 B.t19 324.983
R628 B.n149 B.t12 324.983
R629 B.n146 B.t16 324.983
R630 B.n602 B.t10 297.017
R631 B.n147 B.t18 297.017
R632 B.n474 B.t20 297.017
R633 B.n150 B.t15 297.017
R634 B.n920 B.n919 256.663
R635 B.n920 B.n144 256.663
R636 B.n920 B.n143 256.663
R637 B.n920 B.n142 256.663
R638 B.n920 B.n141 256.663
R639 B.n920 B.n140 256.663
R640 B.n920 B.n139 256.663
R641 B.n920 B.n138 256.663
R642 B.n920 B.n137 256.663
R643 B.n920 B.n136 256.663
R644 B.n920 B.n135 256.663
R645 B.n920 B.n134 256.663
R646 B.n920 B.n133 256.663
R647 B.n920 B.n132 256.663
R648 B.n920 B.n131 256.663
R649 B.n920 B.n130 256.663
R650 B.n920 B.n129 256.663
R651 B.n920 B.n128 256.663
R652 B.n920 B.n127 256.663
R653 B.n920 B.n126 256.663
R654 B.n920 B.n125 256.663
R655 B.n920 B.n124 256.663
R656 B.n920 B.n123 256.663
R657 B.n920 B.n122 256.663
R658 B.n920 B.n121 256.663
R659 B.n920 B.n120 256.663
R660 B.n920 B.n119 256.663
R661 B.n920 B.n118 256.663
R662 B.n920 B.n117 256.663
R663 B.n920 B.n116 256.663
R664 B.n920 B.n115 256.663
R665 B.n920 B.n114 256.663
R666 B.n920 B.n113 256.663
R667 B.n920 B.n112 256.663
R668 B.n920 B.n111 256.663
R669 B.n920 B.n110 256.663
R670 B.n920 B.n109 256.663
R671 B.n920 B.n108 256.663
R672 B.n920 B.n107 256.663
R673 B.n920 B.n106 256.663
R674 B.n920 B.n105 256.663
R675 B.n920 B.n104 256.663
R676 B.n920 B.n103 256.663
R677 B.n920 B.n102 256.663
R678 B.n920 B.n101 256.663
R679 B.n920 B.n100 256.663
R680 B.n920 B.n99 256.663
R681 B.n920 B.n98 256.663
R682 B.n920 B.n97 256.663
R683 B.n497 B.n444 256.663
R684 B.n500 B.n444 256.663
R685 B.n506 B.n444 256.663
R686 B.n508 B.n444 256.663
R687 B.n514 B.n444 256.663
R688 B.n516 B.n444 256.663
R689 B.n522 B.n444 256.663
R690 B.n524 B.n444 256.663
R691 B.n530 B.n444 256.663
R692 B.n532 B.n444 256.663
R693 B.n538 B.n444 256.663
R694 B.n540 B.n444 256.663
R695 B.n546 B.n444 256.663
R696 B.n548 B.n444 256.663
R697 B.n554 B.n444 256.663
R698 B.n556 B.n444 256.663
R699 B.n562 B.n444 256.663
R700 B.n564 B.n444 256.663
R701 B.n570 B.n444 256.663
R702 B.n572 B.n444 256.663
R703 B.n578 B.n444 256.663
R704 B.n580 B.n444 256.663
R705 B.n587 B.n444 256.663
R706 B.n589 B.n444 256.663
R707 B.n595 B.n444 256.663
R708 B.n597 B.n444 256.663
R709 B.n606 B.n444 256.663
R710 B.n608 B.n444 256.663
R711 B.n614 B.n444 256.663
R712 B.n616 B.n444 256.663
R713 B.n622 B.n444 256.663
R714 B.n624 B.n444 256.663
R715 B.n630 B.n444 256.663
R716 B.n632 B.n444 256.663
R717 B.n638 B.n444 256.663
R718 B.n640 B.n444 256.663
R719 B.n646 B.n444 256.663
R720 B.n648 B.n444 256.663
R721 B.n654 B.n444 256.663
R722 B.n656 B.n444 256.663
R723 B.n662 B.n444 256.663
R724 B.n664 B.n444 256.663
R725 B.n670 B.n444 256.663
R726 B.n672 B.n444 256.663
R727 B.n678 B.n444 256.663
R728 B.n680 B.n444 256.663
R729 B.n686 B.n444 256.663
R730 B.n689 B.n444 256.663
R731 B.n696 B.n441 163.367
R732 B.n700 B.n441 163.367
R733 B.n700 B.n435 163.367
R734 B.n708 B.n435 163.367
R735 B.n708 B.n433 163.367
R736 B.n712 B.n433 163.367
R737 B.n712 B.n427 163.367
R738 B.n720 B.n427 163.367
R739 B.n720 B.n425 163.367
R740 B.n724 B.n425 163.367
R741 B.n724 B.n419 163.367
R742 B.n732 B.n419 163.367
R743 B.n732 B.n417 163.367
R744 B.n736 B.n417 163.367
R745 B.n736 B.n411 163.367
R746 B.n744 B.n411 163.367
R747 B.n744 B.n409 163.367
R748 B.n748 B.n409 163.367
R749 B.n748 B.n403 163.367
R750 B.n756 B.n403 163.367
R751 B.n756 B.n401 163.367
R752 B.n760 B.n401 163.367
R753 B.n760 B.n395 163.367
R754 B.n768 B.n395 163.367
R755 B.n768 B.n393 163.367
R756 B.n772 B.n393 163.367
R757 B.n772 B.n387 163.367
R758 B.n780 B.n387 163.367
R759 B.n780 B.n385 163.367
R760 B.n784 B.n385 163.367
R761 B.n784 B.n379 163.367
R762 B.n792 B.n379 163.367
R763 B.n792 B.n377 163.367
R764 B.n796 B.n377 163.367
R765 B.n796 B.n371 163.367
R766 B.n805 B.n371 163.367
R767 B.n805 B.n369 163.367
R768 B.n809 B.n369 163.367
R769 B.n809 B.n364 163.367
R770 B.n817 B.n364 163.367
R771 B.n817 B.n362 163.367
R772 B.n821 B.n362 163.367
R773 B.n821 B.n356 163.367
R774 B.n829 B.n356 163.367
R775 B.n829 B.n354 163.367
R776 B.n833 B.n354 163.367
R777 B.n833 B.n348 163.367
R778 B.n842 B.n348 163.367
R779 B.n842 B.n346 163.367
R780 B.n846 B.n346 163.367
R781 B.n846 B.n2 163.367
R782 B.n1026 B.n2 163.367
R783 B.n1026 B.n3 163.367
R784 B.n1022 B.n3 163.367
R785 B.n1022 B.n9 163.367
R786 B.n1018 B.n9 163.367
R787 B.n1018 B.n11 163.367
R788 B.n1014 B.n11 163.367
R789 B.n1014 B.n16 163.367
R790 B.n1010 B.n16 163.367
R791 B.n1010 B.n18 163.367
R792 B.n1006 B.n18 163.367
R793 B.n1006 B.n23 163.367
R794 B.n1002 B.n23 163.367
R795 B.n1002 B.n25 163.367
R796 B.n998 B.n25 163.367
R797 B.n998 B.n29 163.367
R798 B.n994 B.n29 163.367
R799 B.n994 B.n31 163.367
R800 B.n990 B.n31 163.367
R801 B.n990 B.n37 163.367
R802 B.n986 B.n37 163.367
R803 B.n986 B.n39 163.367
R804 B.n982 B.n39 163.367
R805 B.n982 B.n44 163.367
R806 B.n978 B.n44 163.367
R807 B.n978 B.n46 163.367
R808 B.n974 B.n46 163.367
R809 B.n974 B.n51 163.367
R810 B.n970 B.n51 163.367
R811 B.n970 B.n53 163.367
R812 B.n966 B.n53 163.367
R813 B.n966 B.n58 163.367
R814 B.n962 B.n58 163.367
R815 B.n962 B.n60 163.367
R816 B.n958 B.n60 163.367
R817 B.n958 B.n65 163.367
R818 B.n954 B.n65 163.367
R819 B.n954 B.n67 163.367
R820 B.n950 B.n67 163.367
R821 B.n950 B.n72 163.367
R822 B.n946 B.n72 163.367
R823 B.n946 B.n74 163.367
R824 B.n942 B.n74 163.367
R825 B.n942 B.n79 163.367
R826 B.n938 B.n79 163.367
R827 B.n938 B.n81 163.367
R828 B.n934 B.n81 163.367
R829 B.n934 B.n86 163.367
R830 B.n930 B.n86 163.367
R831 B.n930 B.n88 163.367
R832 B.n926 B.n88 163.367
R833 B.n926 B.n93 163.367
R834 B.n922 B.n93 163.367
R835 B.n499 B.n498 163.367
R836 B.n501 B.n499 163.367
R837 B.n505 B.n494 163.367
R838 B.n509 B.n507 163.367
R839 B.n513 B.n492 163.367
R840 B.n517 B.n515 163.367
R841 B.n521 B.n490 163.367
R842 B.n525 B.n523 163.367
R843 B.n529 B.n488 163.367
R844 B.n533 B.n531 163.367
R845 B.n537 B.n486 163.367
R846 B.n541 B.n539 163.367
R847 B.n545 B.n484 163.367
R848 B.n549 B.n547 163.367
R849 B.n553 B.n482 163.367
R850 B.n557 B.n555 163.367
R851 B.n561 B.n480 163.367
R852 B.n565 B.n563 163.367
R853 B.n569 B.n478 163.367
R854 B.n573 B.n571 163.367
R855 B.n577 B.n476 163.367
R856 B.n581 B.n579 163.367
R857 B.n586 B.n472 163.367
R858 B.n590 B.n588 163.367
R859 B.n594 B.n470 163.367
R860 B.n598 B.n596 163.367
R861 B.n605 B.n468 163.367
R862 B.n609 B.n607 163.367
R863 B.n613 B.n466 163.367
R864 B.n617 B.n615 163.367
R865 B.n621 B.n464 163.367
R866 B.n625 B.n623 163.367
R867 B.n629 B.n462 163.367
R868 B.n633 B.n631 163.367
R869 B.n637 B.n460 163.367
R870 B.n641 B.n639 163.367
R871 B.n645 B.n458 163.367
R872 B.n649 B.n647 163.367
R873 B.n653 B.n456 163.367
R874 B.n657 B.n655 163.367
R875 B.n661 B.n454 163.367
R876 B.n665 B.n663 163.367
R877 B.n669 B.n452 163.367
R878 B.n673 B.n671 163.367
R879 B.n677 B.n450 163.367
R880 B.n681 B.n679 163.367
R881 B.n685 B.n448 163.367
R882 B.n688 B.n687 163.367
R883 B.n690 B.n445 163.367
R884 B.n694 B.n439 163.367
R885 B.n702 B.n439 163.367
R886 B.n702 B.n437 163.367
R887 B.n706 B.n437 163.367
R888 B.n706 B.n430 163.367
R889 B.n714 B.n430 163.367
R890 B.n714 B.n428 163.367
R891 B.n718 B.n428 163.367
R892 B.n718 B.n423 163.367
R893 B.n726 B.n423 163.367
R894 B.n726 B.n421 163.367
R895 B.n730 B.n421 163.367
R896 B.n730 B.n415 163.367
R897 B.n738 B.n415 163.367
R898 B.n738 B.n413 163.367
R899 B.n742 B.n413 163.367
R900 B.n742 B.n406 163.367
R901 B.n750 B.n406 163.367
R902 B.n750 B.n404 163.367
R903 B.n754 B.n404 163.367
R904 B.n754 B.n399 163.367
R905 B.n762 B.n399 163.367
R906 B.n762 B.n397 163.367
R907 B.n766 B.n397 163.367
R908 B.n766 B.n391 163.367
R909 B.n774 B.n391 163.367
R910 B.n774 B.n389 163.367
R911 B.n778 B.n389 163.367
R912 B.n778 B.n383 163.367
R913 B.n786 B.n383 163.367
R914 B.n786 B.n381 163.367
R915 B.n790 B.n381 163.367
R916 B.n790 B.n375 163.367
R917 B.n798 B.n375 163.367
R918 B.n798 B.n373 163.367
R919 B.n802 B.n373 163.367
R920 B.n802 B.n368 163.367
R921 B.n811 B.n368 163.367
R922 B.n811 B.n366 163.367
R923 B.n815 B.n366 163.367
R924 B.n815 B.n360 163.367
R925 B.n823 B.n360 163.367
R926 B.n823 B.n358 163.367
R927 B.n827 B.n358 163.367
R928 B.n827 B.n352 163.367
R929 B.n835 B.n352 163.367
R930 B.n835 B.n350 163.367
R931 B.n840 B.n350 163.367
R932 B.n840 B.n344 163.367
R933 B.n848 B.n344 163.367
R934 B.n849 B.n848 163.367
R935 B.n849 B.n5 163.367
R936 B.n6 B.n5 163.367
R937 B.n7 B.n6 163.367
R938 B.n854 B.n7 163.367
R939 B.n854 B.n12 163.367
R940 B.n13 B.n12 163.367
R941 B.n14 B.n13 163.367
R942 B.n859 B.n14 163.367
R943 B.n859 B.n19 163.367
R944 B.n20 B.n19 163.367
R945 B.n21 B.n20 163.367
R946 B.n864 B.n21 163.367
R947 B.n864 B.n26 163.367
R948 B.n27 B.n26 163.367
R949 B.n28 B.n27 163.367
R950 B.n869 B.n28 163.367
R951 B.n869 B.n33 163.367
R952 B.n34 B.n33 163.367
R953 B.n35 B.n34 163.367
R954 B.n874 B.n35 163.367
R955 B.n874 B.n40 163.367
R956 B.n41 B.n40 163.367
R957 B.n42 B.n41 163.367
R958 B.n879 B.n42 163.367
R959 B.n879 B.n47 163.367
R960 B.n48 B.n47 163.367
R961 B.n49 B.n48 163.367
R962 B.n884 B.n49 163.367
R963 B.n884 B.n54 163.367
R964 B.n55 B.n54 163.367
R965 B.n56 B.n55 163.367
R966 B.n889 B.n56 163.367
R967 B.n889 B.n61 163.367
R968 B.n62 B.n61 163.367
R969 B.n63 B.n62 163.367
R970 B.n894 B.n63 163.367
R971 B.n894 B.n68 163.367
R972 B.n69 B.n68 163.367
R973 B.n70 B.n69 163.367
R974 B.n899 B.n70 163.367
R975 B.n899 B.n75 163.367
R976 B.n76 B.n75 163.367
R977 B.n77 B.n76 163.367
R978 B.n904 B.n77 163.367
R979 B.n904 B.n82 163.367
R980 B.n83 B.n82 163.367
R981 B.n84 B.n83 163.367
R982 B.n909 B.n84 163.367
R983 B.n909 B.n89 163.367
R984 B.n90 B.n89 163.367
R985 B.n91 B.n90 163.367
R986 B.n914 B.n91 163.367
R987 B.n914 B.n96 163.367
R988 B.n154 B.n153 163.367
R989 B.n158 B.n157 163.367
R990 B.n162 B.n161 163.367
R991 B.n166 B.n165 163.367
R992 B.n170 B.n169 163.367
R993 B.n174 B.n173 163.367
R994 B.n178 B.n177 163.367
R995 B.n182 B.n181 163.367
R996 B.n186 B.n185 163.367
R997 B.n190 B.n189 163.367
R998 B.n194 B.n193 163.367
R999 B.n198 B.n197 163.367
R1000 B.n202 B.n201 163.367
R1001 B.n206 B.n205 163.367
R1002 B.n210 B.n209 163.367
R1003 B.n214 B.n213 163.367
R1004 B.n218 B.n217 163.367
R1005 B.n222 B.n221 163.367
R1006 B.n226 B.n225 163.367
R1007 B.n230 B.n229 163.367
R1008 B.n234 B.n233 163.367
R1009 B.n238 B.n237 163.367
R1010 B.n242 B.n241 163.367
R1011 B.n246 B.n245 163.367
R1012 B.n250 B.n249 163.367
R1013 B.n254 B.n253 163.367
R1014 B.n258 B.n257 163.367
R1015 B.n262 B.n261 163.367
R1016 B.n266 B.n265 163.367
R1017 B.n270 B.n269 163.367
R1018 B.n274 B.n273 163.367
R1019 B.n278 B.n277 163.367
R1020 B.n282 B.n281 163.367
R1021 B.n286 B.n285 163.367
R1022 B.n290 B.n289 163.367
R1023 B.n294 B.n293 163.367
R1024 B.n298 B.n297 163.367
R1025 B.n302 B.n301 163.367
R1026 B.n306 B.n305 163.367
R1027 B.n310 B.n309 163.367
R1028 B.n314 B.n313 163.367
R1029 B.n318 B.n317 163.367
R1030 B.n322 B.n321 163.367
R1031 B.n326 B.n325 163.367
R1032 B.n330 B.n329 163.367
R1033 B.n334 B.n333 163.367
R1034 B.n338 B.n337 163.367
R1035 B.n340 B.n145 163.367
R1036 B.n695 B.n444 72.2212
R1037 B.n921 B.n920 72.2212
R1038 B.n497 B.n443 71.676
R1039 B.n501 B.n500 71.676
R1040 B.n506 B.n505 71.676
R1041 B.n509 B.n508 71.676
R1042 B.n514 B.n513 71.676
R1043 B.n517 B.n516 71.676
R1044 B.n522 B.n521 71.676
R1045 B.n525 B.n524 71.676
R1046 B.n530 B.n529 71.676
R1047 B.n533 B.n532 71.676
R1048 B.n538 B.n537 71.676
R1049 B.n541 B.n540 71.676
R1050 B.n546 B.n545 71.676
R1051 B.n549 B.n548 71.676
R1052 B.n554 B.n553 71.676
R1053 B.n557 B.n556 71.676
R1054 B.n562 B.n561 71.676
R1055 B.n565 B.n564 71.676
R1056 B.n570 B.n569 71.676
R1057 B.n573 B.n572 71.676
R1058 B.n578 B.n577 71.676
R1059 B.n581 B.n580 71.676
R1060 B.n587 B.n586 71.676
R1061 B.n590 B.n589 71.676
R1062 B.n595 B.n594 71.676
R1063 B.n598 B.n597 71.676
R1064 B.n606 B.n605 71.676
R1065 B.n609 B.n608 71.676
R1066 B.n614 B.n613 71.676
R1067 B.n617 B.n616 71.676
R1068 B.n622 B.n621 71.676
R1069 B.n625 B.n624 71.676
R1070 B.n630 B.n629 71.676
R1071 B.n633 B.n632 71.676
R1072 B.n638 B.n637 71.676
R1073 B.n641 B.n640 71.676
R1074 B.n646 B.n645 71.676
R1075 B.n649 B.n648 71.676
R1076 B.n654 B.n653 71.676
R1077 B.n657 B.n656 71.676
R1078 B.n662 B.n661 71.676
R1079 B.n665 B.n664 71.676
R1080 B.n670 B.n669 71.676
R1081 B.n673 B.n672 71.676
R1082 B.n678 B.n677 71.676
R1083 B.n681 B.n680 71.676
R1084 B.n686 B.n685 71.676
R1085 B.n689 B.n688 71.676
R1086 B.n97 B.n95 71.676
R1087 B.n154 B.n98 71.676
R1088 B.n158 B.n99 71.676
R1089 B.n162 B.n100 71.676
R1090 B.n166 B.n101 71.676
R1091 B.n170 B.n102 71.676
R1092 B.n174 B.n103 71.676
R1093 B.n178 B.n104 71.676
R1094 B.n182 B.n105 71.676
R1095 B.n186 B.n106 71.676
R1096 B.n190 B.n107 71.676
R1097 B.n194 B.n108 71.676
R1098 B.n198 B.n109 71.676
R1099 B.n202 B.n110 71.676
R1100 B.n206 B.n111 71.676
R1101 B.n210 B.n112 71.676
R1102 B.n214 B.n113 71.676
R1103 B.n218 B.n114 71.676
R1104 B.n222 B.n115 71.676
R1105 B.n226 B.n116 71.676
R1106 B.n230 B.n117 71.676
R1107 B.n234 B.n118 71.676
R1108 B.n238 B.n119 71.676
R1109 B.n242 B.n120 71.676
R1110 B.n246 B.n121 71.676
R1111 B.n250 B.n122 71.676
R1112 B.n254 B.n123 71.676
R1113 B.n258 B.n124 71.676
R1114 B.n262 B.n125 71.676
R1115 B.n266 B.n126 71.676
R1116 B.n270 B.n127 71.676
R1117 B.n274 B.n128 71.676
R1118 B.n278 B.n129 71.676
R1119 B.n282 B.n130 71.676
R1120 B.n286 B.n131 71.676
R1121 B.n290 B.n132 71.676
R1122 B.n294 B.n133 71.676
R1123 B.n298 B.n134 71.676
R1124 B.n302 B.n135 71.676
R1125 B.n306 B.n136 71.676
R1126 B.n310 B.n137 71.676
R1127 B.n314 B.n138 71.676
R1128 B.n318 B.n139 71.676
R1129 B.n322 B.n140 71.676
R1130 B.n326 B.n141 71.676
R1131 B.n330 B.n142 71.676
R1132 B.n334 B.n143 71.676
R1133 B.n338 B.n144 71.676
R1134 B.n919 B.n145 71.676
R1135 B.n919 B.n918 71.676
R1136 B.n340 B.n144 71.676
R1137 B.n337 B.n143 71.676
R1138 B.n333 B.n142 71.676
R1139 B.n329 B.n141 71.676
R1140 B.n325 B.n140 71.676
R1141 B.n321 B.n139 71.676
R1142 B.n317 B.n138 71.676
R1143 B.n313 B.n137 71.676
R1144 B.n309 B.n136 71.676
R1145 B.n305 B.n135 71.676
R1146 B.n301 B.n134 71.676
R1147 B.n297 B.n133 71.676
R1148 B.n293 B.n132 71.676
R1149 B.n289 B.n131 71.676
R1150 B.n285 B.n130 71.676
R1151 B.n281 B.n129 71.676
R1152 B.n277 B.n128 71.676
R1153 B.n273 B.n127 71.676
R1154 B.n269 B.n126 71.676
R1155 B.n265 B.n125 71.676
R1156 B.n261 B.n124 71.676
R1157 B.n257 B.n123 71.676
R1158 B.n253 B.n122 71.676
R1159 B.n249 B.n121 71.676
R1160 B.n245 B.n120 71.676
R1161 B.n241 B.n119 71.676
R1162 B.n237 B.n118 71.676
R1163 B.n233 B.n117 71.676
R1164 B.n229 B.n116 71.676
R1165 B.n225 B.n115 71.676
R1166 B.n221 B.n114 71.676
R1167 B.n217 B.n113 71.676
R1168 B.n213 B.n112 71.676
R1169 B.n209 B.n111 71.676
R1170 B.n205 B.n110 71.676
R1171 B.n201 B.n109 71.676
R1172 B.n197 B.n108 71.676
R1173 B.n193 B.n107 71.676
R1174 B.n189 B.n106 71.676
R1175 B.n185 B.n105 71.676
R1176 B.n181 B.n104 71.676
R1177 B.n177 B.n103 71.676
R1178 B.n173 B.n102 71.676
R1179 B.n169 B.n101 71.676
R1180 B.n165 B.n100 71.676
R1181 B.n161 B.n99 71.676
R1182 B.n157 B.n98 71.676
R1183 B.n153 B.n97 71.676
R1184 B.n498 B.n497 71.676
R1185 B.n500 B.n494 71.676
R1186 B.n507 B.n506 71.676
R1187 B.n508 B.n492 71.676
R1188 B.n515 B.n514 71.676
R1189 B.n516 B.n490 71.676
R1190 B.n523 B.n522 71.676
R1191 B.n524 B.n488 71.676
R1192 B.n531 B.n530 71.676
R1193 B.n532 B.n486 71.676
R1194 B.n539 B.n538 71.676
R1195 B.n540 B.n484 71.676
R1196 B.n547 B.n546 71.676
R1197 B.n548 B.n482 71.676
R1198 B.n555 B.n554 71.676
R1199 B.n556 B.n480 71.676
R1200 B.n563 B.n562 71.676
R1201 B.n564 B.n478 71.676
R1202 B.n571 B.n570 71.676
R1203 B.n572 B.n476 71.676
R1204 B.n579 B.n578 71.676
R1205 B.n580 B.n472 71.676
R1206 B.n588 B.n587 71.676
R1207 B.n589 B.n470 71.676
R1208 B.n596 B.n595 71.676
R1209 B.n597 B.n468 71.676
R1210 B.n607 B.n606 71.676
R1211 B.n608 B.n466 71.676
R1212 B.n615 B.n614 71.676
R1213 B.n616 B.n464 71.676
R1214 B.n623 B.n622 71.676
R1215 B.n624 B.n462 71.676
R1216 B.n631 B.n630 71.676
R1217 B.n632 B.n460 71.676
R1218 B.n639 B.n638 71.676
R1219 B.n640 B.n458 71.676
R1220 B.n647 B.n646 71.676
R1221 B.n648 B.n456 71.676
R1222 B.n655 B.n654 71.676
R1223 B.n656 B.n454 71.676
R1224 B.n663 B.n662 71.676
R1225 B.n664 B.n452 71.676
R1226 B.n671 B.n670 71.676
R1227 B.n672 B.n450 71.676
R1228 B.n679 B.n678 71.676
R1229 B.n680 B.n448 71.676
R1230 B.n687 B.n686 71.676
R1231 B.n690 B.n689 71.676
R1232 B.n603 B.n602 59.5399
R1233 B.n583 B.n474 59.5399
R1234 B.n151 B.n150 59.5399
R1235 B.n148 B.n147 59.5399
R1236 B.n602 B.n601 57.7944
R1237 B.n474 B.n473 57.7944
R1238 B.n150 B.n149 57.7944
R1239 B.n147 B.n146 57.7944
R1240 B.n695 B.n440 41.2695
R1241 B.n701 B.n440 41.2695
R1242 B.n701 B.n436 41.2695
R1243 B.n707 B.n436 41.2695
R1244 B.n707 B.n431 41.2695
R1245 B.n713 B.n431 41.2695
R1246 B.n713 B.n432 41.2695
R1247 B.n719 B.n424 41.2695
R1248 B.n725 B.n424 41.2695
R1249 B.n725 B.n420 41.2695
R1250 B.n731 B.n420 41.2695
R1251 B.n731 B.n416 41.2695
R1252 B.n737 B.n416 41.2695
R1253 B.n737 B.n412 41.2695
R1254 B.n743 B.n412 41.2695
R1255 B.n743 B.n407 41.2695
R1256 B.n749 B.n407 41.2695
R1257 B.n749 B.n408 41.2695
R1258 B.n755 B.n400 41.2695
R1259 B.n761 B.n400 41.2695
R1260 B.n761 B.n396 41.2695
R1261 B.n767 B.n396 41.2695
R1262 B.n767 B.n392 41.2695
R1263 B.n773 B.n392 41.2695
R1264 B.n773 B.n388 41.2695
R1265 B.n779 B.n388 41.2695
R1266 B.n785 B.n384 41.2695
R1267 B.n785 B.n380 41.2695
R1268 B.n791 B.n380 41.2695
R1269 B.n791 B.n376 41.2695
R1270 B.n797 B.n376 41.2695
R1271 B.n797 B.n372 41.2695
R1272 B.n804 B.n372 41.2695
R1273 B.n804 B.n803 41.2695
R1274 B.n810 B.n365 41.2695
R1275 B.n816 B.n365 41.2695
R1276 B.n816 B.n361 41.2695
R1277 B.n822 B.n361 41.2695
R1278 B.n822 B.n357 41.2695
R1279 B.n828 B.n357 41.2695
R1280 B.n828 B.n353 41.2695
R1281 B.n834 B.n353 41.2695
R1282 B.n841 B.n349 41.2695
R1283 B.n841 B.n345 41.2695
R1284 B.n847 B.n345 41.2695
R1285 B.n847 B.n4 41.2695
R1286 B.n1025 B.n4 41.2695
R1287 B.n1025 B.n1024 41.2695
R1288 B.n1024 B.n1023 41.2695
R1289 B.n1023 B.n8 41.2695
R1290 B.n1017 B.n8 41.2695
R1291 B.n1017 B.n1016 41.2695
R1292 B.n1015 B.n15 41.2695
R1293 B.n1009 B.n15 41.2695
R1294 B.n1009 B.n1008 41.2695
R1295 B.n1008 B.n1007 41.2695
R1296 B.n1007 B.n22 41.2695
R1297 B.n1001 B.n22 41.2695
R1298 B.n1001 B.n1000 41.2695
R1299 B.n1000 B.n999 41.2695
R1300 B.n993 B.n32 41.2695
R1301 B.n993 B.n992 41.2695
R1302 B.n992 B.n991 41.2695
R1303 B.n991 B.n36 41.2695
R1304 B.n985 B.n36 41.2695
R1305 B.n985 B.n984 41.2695
R1306 B.n984 B.n983 41.2695
R1307 B.n983 B.n43 41.2695
R1308 B.n977 B.n976 41.2695
R1309 B.n976 B.n975 41.2695
R1310 B.n975 B.n50 41.2695
R1311 B.n969 B.n50 41.2695
R1312 B.n969 B.n968 41.2695
R1313 B.n968 B.n967 41.2695
R1314 B.n967 B.n57 41.2695
R1315 B.n961 B.n57 41.2695
R1316 B.n960 B.n959 41.2695
R1317 B.n959 B.n64 41.2695
R1318 B.n953 B.n64 41.2695
R1319 B.n953 B.n952 41.2695
R1320 B.n952 B.n951 41.2695
R1321 B.n951 B.n71 41.2695
R1322 B.n945 B.n71 41.2695
R1323 B.n945 B.n944 41.2695
R1324 B.n944 B.n943 41.2695
R1325 B.n943 B.n78 41.2695
R1326 B.n937 B.n78 41.2695
R1327 B.n936 B.n935 41.2695
R1328 B.n935 B.n85 41.2695
R1329 B.n929 B.n85 41.2695
R1330 B.n929 B.n928 41.2695
R1331 B.n928 B.n927 41.2695
R1332 B.n927 B.n92 41.2695
R1333 B.n921 B.n92 41.2695
R1334 B.t7 B.n349 40.6626
R1335 B.n1016 B.t6 40.6626
R1336 B.n432 B.t9 30.9522
R1337 B.n810 B.t3 30.9522
R1338 B.n999 B.t0 30.9522
R1339 B.t13 B.n936 30.9522
R1340 B.n923 B.n94 30.7517
R1341 B.n917 B.n916 30.7517
R1342 B.n693 B.n692 30.7517
R1343 B.n697 B.n442 30.7517
R1344 B.n408 B.t5 29.7384
R1345 B.t2 B.n960 29.7384
R1346 B.t4 B.n384 21.2419
R1347 B.t1 B.n43 21.2419
R1348 B.n779 B.t4 20.0281
R1349 B.n977 B.t1 20.0281
R1350 B B.n1027 18.0485
R1351 B.n755 B.t5 11.5315
R1352 B.n961 B.t2 11.5315
R1353 B.n152 B.n94 10.6151
R1354 B.n155 B.n152 10.6151
R1355 B.n156 B.n155 10.6151
R1356 B.n159 B.n156 10.6151
R1357 B.n160 B.n159 10.6151
R1358 B.n163 B.n160 10.6151
R1359 B.n164 B.n163 10.6151
R1360 B.n167 B.n164 10.6151
R1361 B.n168 B.n167 10.6151
R1362 B.n171 B.n168 10.6151
R1363 B.n172 B.n171 10.6151
R1364 B.n175 B.n172 10.6151
R1365 B.n176 B.n175 10.6151
R1366 B.n179 B.n176 10.6151
R1367 B.n180 B.n179 10.6151
R1368 B.n183 B.n180 10.6151
R1369 B.n184 B.n183 10.6151
R1370 B.n187 B.n184 10.6151
R1371 B.n188 B.n187 10.6151
R1372 B.n191 B.n188 10.6151
R1373 B.n192 B.n191 10.6151
R1374 B.n195 B.n192 10.6151
R1375 B.n196 B.n195 10.6151
R1376 B.n199 B.n196 10.6151
R1377 B.n200 B.n199 10.6151
R1378 B.n203 B.n200 10.6151
R1379 B.n204 B.n203 10.6151
R1380 B.n207 B.n204 10.6151
R1381 B.n208 B.n207 10.6151
R1382 B.n211 B.n208 10.6151
R1383 B.n212 B.n211 10.6151
R1384 B.n215 B.n212 10.6151
R1385 B.n216 B.n215 10.6151
R1386 B.n219 B.n216 10.6151
R1387 B.n220 B.n219 10.6151
R1388 B.n223 B.n220 10.6151
R1389 B.n224 B.n223 10.6151
R1390 B.n227 B.n224 10.6151
R1391 B.n228 B.n227 10.6151
R1392 B.n231 B.n228 10.6151
R1393 B.n232 B.n231 10.6151
R1394 B.n235 B.n232 10.6151
R1395 B.n236 B.n235 10.6151
R1396 B.n240 B.n239 10.6151
R1397 B.n243 B.n240 10.6151
R1398 B.n244 B.n243 10.6151
R1399 B.n247 B.n244 10.6151
R1400 B.n248 B.n247 10.6151
R1401 B.n251 B.n248 10.6151
R1402 B.n252 B.n251 10.6151
R1403 B.n255 B.n252 10.6151
R1404 B.n256 B.n255 10.6151
R1405 B.n260 B.n259 10.6151
R1406 B.n263 B.n260 10.6151
R1407 B.n264 B.n263 10.6151
R1408 B.n267 B.n264 10.6151
R1409 B.n268 B.n267 10.6151
R1410 B.n271 B.n268 10.6151
R1411 B.n272 B.n271 10.6151
R1412 B.n275 B.n272 10.6151
R1413 B.n276 B.n275 10.6151
R1414 B.n279 B.n276 10.6151
R1415 B.n280 B.n279 10.6151
R1416 B.n283 B.n280 10.6151
R1417 B.n284 B.n283 10.6151
R1418 B.n287 B.n284 10.6151
R1419 B.n288 B.n287 10.6151
R1420 B.n291 B.n288 10.6151
R1421 B.n292 B.n291 10.6151
R1422 B.n295 B.n292 10.6151
R1423 B.n296 B.n295 10.6151
R1424 B.n299 B.n296 10.6151
R1425 B.n300 B.n299 10.6151
R1426 B.n303 B.n300 10.6151
R1427 B.n304 B.n303 10.6151
R1428 B.n307 B.n304 10.6151
R1429 B.n308 B.n307 10.6151
R1430 B.n311 B.n308 10.6151
R1431 B.n312 B.n311 10.6151
R1432 B.n315 B.n312 10.6151
R1433 B.n316 B.n315 10.6151
R1434 B.n319 B.n316 10.6151
R1435 B.n320 B.n319 10.6151
R1436 B.n323 B.n320 10.6151
R1437 B.n324 B.n323 10.6151
R1438 B.n327 B.n324 10.6151
R1439 B.n328 B.n327 10.6151
R1440 B.n331 B.n328 10.6151
R1441 B.n332 B.n331 10.6151
R1442 B.n335 B.n332 10.6151
R1443 B.n336 B.n335 10.6151
R1444 B.n339 B.n336 10.6151
R1445 B.n341 B.n339 10.6151
R1446 B.n342 B.n341 10.6151
R1447 B.n917 B.n342 10.6151
R1448 B.n693 B.n438 10.6151
R1449 B.n703 B.n438 10.6151
R1450 B.n704 B.n703 10.6151
R1451 B.n705 B.n704 10.6151
R1452 B.n705 B.n429 10.6151
R1453 B.n715 B.n429 10.6151
R1454 B.n716 B.n715 10.6151
R1455 B.n717 B.n716 10.6151
R1456 B.n717 B.n422 10.6151
R1457 B.n727 B.n422 10.6151
R1458 B.n728 B.n727 10.6151
R1459 B.n729 B.n728 10.6151
R1460 B.n729 B.n414 10.6151
R1461 B.n739 B.n414 10.6151
R1462 B.n740 B.n739 10.6151
R1463 B.n741 B.n740 10.6151
R1464 B.n741 B.n405 10.6151
R1465 B.n751 B.n405 10.6151
R1466 B.n752 B.n751 10.6151
R1467 B.n753 B.n752 10.6151
R1468 B.n753 B.n398 10.6151
R1469 B.n763 B.n398 10.6151
R1470 B.n764 B.n763 10.6151
R1471 B.n765 B.n764 10.6151
R1472 B.n765 B.n390 10.6151
R1473 B.n775 B.n390 10.6151
R1474 B.n776 B.n775 10.6151
R1475 B.n777 B.n776 10.6151
R1476 B.n777 B.n382 10.6151
R1477 B.n787 B.n382 10.6151
R1478 B.n788 B.n787 10.6151
R1479 B.n789 B.n788 10.6151
R1480 B.n789 B.n374 10.6151
R1481 B.n799 B.n374 10.6151
R1482 B.n800 B.n799 10.6151
R1483 B.n801 B.n800 10.6151
R1484 B.n801 B.n367 10.6151
R1485 B.n812 B.n367 10.6151
R1486 B.n813 B.n812 10.6151
R1487 B.n814 B.n813 10.6151
R1488 B.n814 B.n359 10.6151
R1489 B.n824 B.n359 10.6151
R1490 B.n825 B.n824 10.6151
R1491 B.n826 B.n825 10.6151
R1492 B.n826 B.n351 10.6151
R1493 B.n836 B.n351 10.6151
R1494 B.n837 B.n836 10.6151
R1495 B.n839 B.n837 10.6151
R1496 B.n839 B.n838 10.6151
R1497 B.n838 B.n343 10.6151
R1498 B.n850 B.n343 10.6151
R1499 B.n851 B.n850 10.6151
R1500 B.n852 B.n851 10.6151
R1501 B.n853 B.n852 10.6151
R1502 B.n855 B.n853 10.6151
R1503 B.n856 B.n855 10.6151
R1504 B.n857 B.n856 10.6151
R1505 B.n858 B.n857 10.6151
R1506 B.n860 B.n858 10.6151
R1507 B.n861 B.n860 10.6151
R1508 B.n862 B.n861 10.6151
R1509 B.n863 B.n862 10.6151
R1510 B.n865 B.n863 10.6151
R1511 B.n866 B.n865 10.6151
R1512 B.n867 B.n866 10.6151
R1513 B.n868 B.n867 10.6151
R1514 B.n870 B.n868 10.6151
R1515 B.n871 B.n870 10.6151
R1516 B.n872 B.n871 10.6151
R1517 B.n873 B.n872 10.6151
R1518 B.n875 B.n873 10.6151
R1519 B.n876 B.n875 10.6151
R1520 B.n877 B.n876 10.6151
R1521 B.n878 B.n877 10.6151
R1522 B.n880 B.n878 10.6151
R1523 B.n881 B.n880 10.6151
R1524 B.n882 B.n881 10.6151
R1525 B.n883 B.n882 10.6151
R1526 B.n885 B.n883 10.6151
R1527 B.n886 B.n885 10.6151
R1528 B.n887 B.n886 10.6151
R1529 B.n888 B.n887 10.6151
R1530 B.n890 B.n888 10.6151
R1531 B.n891 B.n890 10.6151
R1532 B.n892 B.n891 10.6151
R1533 B.n893 B.n892 10.6151
R1534 B.n895 B.n893 10.6151
R1535 B.n896 B.n895 10.6151
R1536 B.n897 B.n896 10.6151
R1537 B.n898 B.n897 10.6151
R1538 B.n900 B.n898 10.6151
R1539 B.n901 B.n900 10.6151
R1540 B.n902 B.n901 10.6151
R1541 B.n903 B.n902 10.6151
R1542 B.n905 B.n903 10.6151
R1543 B.n906 B.n905 10.6151
R1544 B.n907 B.n906 10.6151
R1545 B.n908 B.n907 10.6151
R1546 B.n910 B.n908 10.6151
R1547 B.n911 B.n910 10.6151
R1548 B.n912 B.n911 10.6151
R1549 B.n913 B.n912 10.6151
R1550 B.n915 B.n913 10.6151
R1551 B.n916 B.n915 10.6151
R1552 B.n496 B.n442 10.6151
R1553 B.n496 B.n495 10.6151
R1554 B.n502 B.n495 10.6151
R1555 B.n503 B.n502 10.6151
R1556 B.n504 B.n503 10.6151
R1557 B.n504 B.n493 10.6151
R1558 B.n510 B.n493 10.6151
R1559 B.n511 B.n510 10.6151
R1560 B.n512 B.n511 10.6151
R1561 B.n512 B.n491 10.6151
R1562 B.n518 B.n491 10.6151
R1563 B.n519 B.n518 10.6151
R1564 B.n520 B.n519 10.6151
R1565 B.n520 B.n489 10.6151
R1566 B.n526 B.n489 10.6151
R1567 B.n527 B.n526 10.6151
R1568 B.n528 B.n527 10.6151
R1569 B.n528 B.n487 10.6151
R1570 B.n534 B.n487 10.6151
R1571 B.n535 B.n534 10.6151
R1572 B.n536 B.n535 10.6151
R1573 B.n536 B.n485 10.6151
R1574 B.n542 B.n485 10.6151
R1575 B.n543 B.n542 10.6151
R1576 B.n544 B.n543 10.6151
R1577 B.n544 B.n483 10.6151
R1578 B.n550 B.n483 10.6151
R1579 B.n551 B.n550 10.6151
R1580 B.n552 B.n551 10.6151
R1581 B.n552 B.n481 10.6151
R1582 B.n558 B.n481 10.6151
R1583 B.n559 B.n558 10.6151
R1584 B.n560 B.n559 10.6151
R1585 B.n560 B.n479 10.6151
R1586 B.n566 B.n479 10.6151
R1587 B.n567 B.n566 10.6151
R1588 B.n568 B.n567 10.6151
R1589 B.n568 B.n477 10.6151
R1590 B.n574 B.n477 10.6151
R1591 B.n575 B.n574 10.6151
R1592 B.n576 B.n575 10.6151
R1593 B.n576 B.n475 10.6151
R1594 B.n582 B.n475 10.6151
R1595 B.n585 B.n584 10.6151
R1596 B.n585 B.n471 10.6151
R1597 B.n591 B.n471 10.6151
R1598 B.n592 B.n591 10.6151
R1599 B.n593 B.n592 10.6151
R1600 B.n593 B.n469 10.6151
R1601 B.n599 B.n469 10.6151
R1602 B.n600 B.n599 10.6151
R1603 B.n604 B.n600 10.6151
R1604 B.n610 B.n467 10.6151
R1605 B.n611 B.n610 10.6151
R1606 B.n612 B.n611 10.6151
R1607 B.n612 B.n465 10.6151
R1608 B.n618 B.n465 10.6151
R1609 B.n619 B.n618 10.6151
R1610 B.n620 B.n619 10.6151
R1611 B.n620 B.n463 10.6151
R1612 B.n626 B.n463 10.6151
R1613 B.n627 B.n626 10.6151
R1614 B.n628 B.n627 10.6151
R1615 B.n628 B.n461 10.6151
R1616 B.n634 B.n461 10.6151
R1617 B.n635 B.n634 10.6151
R1618 B.n636 B.n635 10.6151
R1619 B.n636 B.n459 10.6151
R1620 B.n642 B.n459 10.6151
R1621 B.n643 B.n642 10.6151
R1622 B.n644 B.n643 10.6151
R1623 B.n644 B.n457 10.6151
R1624 B.n650 B.n457 10.6151
R1625 B.n651 B.n650 10.6151
R1626 B.n652 B.n651 10.6151
R1627 B.n652 B.n455 10.6151
R1628 B.n658 B.n455 10.6151
R1629 B.n659 B.n658 10.6151
R1630 B.n660 B.n659 10.6151
R1631 B.n660 B.n453 10.6151
R1632 B.n666 B.n453 10.6151
R1633 B.n667 B.n666 10.6151
R1634 B.n668 B.n667 10.6151
R1635 B.n668 B.n451 10.6151
R1636 B.n674 B.n451 10.6151
R1637 B.n675 B.n674 10.6151
R1638 B.n676 B.n675 10.6151
R1639 B.n676 B.n449 10.6151
R1640 B.n682 B.n449 10.6151
R1641 B.n683 B.n682 10.6151
R1642 B.n684 B.n683 10.6151
R1643 B.n684 B.n447 10.6151
R1644 B.n447 B.n446 10.6151
R1645 B.n691 B.n446 10.6151
R1646 B.n692 B.n691 10.6151
R1647 B.n698 B.n697 10.6151
R1648 B.n699 B.n698 10.6151
R1649 B.n699 B.n434 10.6151
R1650 B.n709 B.n434 10.6151
R1651 B.n710 B.n709 10.6151
R1652 B.n711 B.n710 10.6151
R1653 B.n711 B.n426 10.6151
R1654 B.n721 B.n426 10.6151
R1655 B.n722 B.n721 10.6151
R1656 B.n723 B.n722 10.6151
R1657 B.n723 B.n418 10.6151
R1658 B.n733 B.n418 10.6151
R1659 B.n734 B.n733 10.6151
R1660 B.n735 B.n734 10.6151
R1661 B.n735 B.n410 10.6151
R1662 B.n745 B.n410 10.6151
R1663 B.n746 B.n745 10.6151
R1664 B.n747 B.n746 10.6151
R1665 B.n747 B.n402 10.6151
R1666 B.n757 B.n402 10.6151
R1667 B.n758 B.n757 10.6151
R1668 B.n759 B.n758 10.6151
R1669 B.n759 B.n394 10.6151
R1670 B.n769 B.n394 10.6151
R1671 B.n770 B.n769 10.6151
R1672 B.n771 B.n770 10.6151
R1673 B.n771 B.n386 10.6151
R1674 B.n781 B.n386 10.6151
R1675 B.n782 B.n781 10.6151
R1676 B.n783 B.n782 10.6151
R1677 B.n783 B.n378 10.6151
R1678 B.n793 B.n378 10.6151
R1679 B.n794 B.n793 10.6151
R1680 B.n795 B.n794 10.6151
R1681 B.n795 B.n370 10.6151
R1682 B.n806 B.n370 10.6151
R1683 B.n807 B.n806 10.6151
R1684 B.n808 B.n807 10.6151
R1685 B.n808 B.n363 10.6151
R1686 B.n818 B.n363 10.6151
R1687 B.n819 B.n818 10.6151
R1688 B.n820 B.n819 10.6151
R1689 B.n820 B.n355 10.6151
R1690 B.n830 B.n355 10.6151
R1691 B.n831 B.n830 10.6151
R1692 B.n832 B.n831 10.6151
R1693 B.n832 B.n347 10.6151
R1694 B.n843 B.n347 10.6151
R1695 B.n844 B.n843 10.6151
R1696 B.n845 B.n844 10.6151
R1697 B.n845 B.n0 10.6151
R1698 B.n1021 B.n1 10.6151
R1699 B.n1021 B.n1020 10.6151
R1700 B.n1020 B.n1019 10.6151
R1701 B.n1019 B.n10 10.6151
R1702 B.n1013 B.n10 10.6151
R1703 B.n1013 B.n1012 10.6151
R1704 B.n1012 B.n1011 10.6151
R1705 B.n1011 B.n17 10.6151
R1706 B.n1005 B.n17 10.6151
R1707 B.n1005 B.n1004 10.6151
R1708 B.n1004 B.n1003 10.6151
R1709 B.n1003 B.n24 10.6151
R1710 B.n997 B.n24 10.6151
R1711 B.n997 B.n996 10.6151
R1712 B.n996 B.n995 10.6151
R1713 B.n995 B.n30 10.6151
R1714 B.n989 B.n30 10.6151
R1715 B.n989 B.n988 10.6151
R1716 B.n988 B.n987 10.6151
R1717 B.n987 B.n38 10.6151
R1718 B.n981 B.n38 10.6151
R1719 B.n981 B.n980 10.6151
R1720 B.n980 B.n979 10.6151
R1721 B.n979 B.n45 10.6151
R1722 B.n973 B.n45 10.6151
R1723 B.n973 B.n972 10.6151
R1724 B.n972 B.n971 10.6151
R1725 B.n971 B.n52 10.6151
R1726 B.n965 B.n52 10.6151
R1727 B.n965 B.n964 10.6151
R1728 B.n964 B.n963 10.6151
R1729 B.n963 B.n59 10.6151
R1730 B.n957 B.n59 10.6151
R1731 B.n957 B.n956 10.6151
R1732 B.n956 B.n955 10.6151
R1733 B.n955 B.n66 10.6151
R1734 B.n949 B.n66 10.6151
R1735 B.n949 B.n948 10.6151
R1736 B.n948 B.n947 10.6151
R1737 B.n947 B.n73 10.6151
R1738 B.n941 B.n73 10.6151
R1739 B.n941 B.n940 10.6151
R1740 B.n940 B.n939 10.6151
R1741 B.n939 B.n80 10.6151
R1742 B.n933 B.n80 10.6151
R1743 B.n933 B.n932 10.6151
R1744 B.n932 B.n931 10.6151
R1745 B.n931 B.n87 10.6151
R1746 B.n925 B.n87 10.6151
R1747 B.n925 B.n924 10.6151
R1748 B.n924 B.n923 10.6151
R1749 B.n719 B.t9 10.3177
R1750 B.n803 B.t3 10.3177
R1751 B.n32 B.t0 10.3177
R1752 B.n937 B.t13 10.3177
R1753 B.n236 B.n151 9.36635
R1754 B.n259 B.n148 9.36635
R1755 B.n583 B.n582 9.36635
R1756 B.n603 B.n467 9.36635
R1757 B.n1027 B.n0 2.81026
R1758 B.n1027 B.n1 2.81026
R1759 B.n239 B.n151 1.24928
R1760 B.n256 B.n148 1.24928
R1761 B.n584 B.n583 1.24928
R1762 B.n604 B.n603 1.24928
R1763 B.n834 B.t7 0.607397
R1764 B.t6 B.n1015 0.607397
R1765 VP.n19 VP.n16 161.3
R1766 VP.n21 VP.n20 161.3
R1767 VP.n22 VP.n15 161.3
R1768 VP.n24 VP.n23 161.3
R1769 VP.n25 VP.n14 161.3
R1770 VP.n27 VP.n26 161.3
R1771 VP.n29 VP.n28 161.3
R1772 VP.n30 VP.n12 161.3
R1773 VP.n32 VP.n31 161.3
R1774 VP.n33 VP.n11 161.3
R1775 VP.n35 VP.n34 161.3
R1776 VP.n36 VP.n10 161.3
R1777 VP.n68 VP.n0 161.3
R1778 VP.n67 VP.n66 161.3
R1779 VP.n65 VP.n1 161.3
R1780 VP.n64 VP.n63 161.3
R1781 VP.n62 VP.n2 161.3
R1782 VP.n61 VP.n60 161.3
R1783 VP.n59 VP.n58 161.3
R1784 VP.n57 VP.n4 161.3
R1785 VP.n56 VP.n55 161.3
R1786 VP.n54 VP.n5 161.3
R1787 VP.n53 VP.n52 161.3
R1788 VP.n51 VP.n6 161.3
R1789 VP.n49 VP.n48 161.3
R1790 VP.n47 VP.n7 161.3
R1791 VP.n46 VP.n45 161.3
R1792 VP.n44 VP.n8 161.3
R1793 VP.n43 VP.n42 161.3
R1794 VP.n41 VP.n9 161.3
R1795 VP.n17 VP.t4 150.681
R1796 VP.n39 VP.t2 116.862
R1797 VP.n50 VP.t6 116.862
R1798 VP.n3 VP.t0 116.862
R1799 VP.n69 VP.t1 116.862
R1800 VP.n37 VP.t5 116.862
R1801 VP.n13 VP.t3 116.862
R1802 VP.n18 VP.t7 116.862
R1803 VP.n40 VP.n39 99.991
R1804 VP.n70 VP.n69 99.991
R1805 VP.n38 VP.n37 99.991
R1806 VP.n18 VP.n17 60.757
R1807 VP.n45 VP.n44 56.5193
R1808 VP.n56 VP.n5 56.5193
R1809 VP.n63 VP.n1 56.5193
R1810 VP.n31 VP.n11 56.5193
R1811 VP.n24 VP.n15 56.5193
R1812 VP.n40 VP.n38 51.8178
R1813 VP.n43 VP.n9 24.4675
R1814 VP.n44 VP.n43 24.4675
R1815 VP.n45 VP.n7 24.4675
R1816 VP.n49 VP.n7 24.4675
R1817 VP.n52 VP.n51 24.4675
R1818 VP.n52 VP.n5 24.4675
R1819 VP.n57 VP.n56 24.4675
R1820 VP.n58 VP.n57 24.4675
R1821 VP.n62 VP.n61 24.4675
R1822 VP.n63 VP.n62 24.4675
R1823 VP.n67 VP.n1 24.4675
R1824 VP.n68 VP.n67 24.4675
R1825 VP.n35 VP.n11 24.4675
R1826 VP.n36 VP.n35 24.4675
R1827 VP.n25 VP.n24 24.4675
R1828 VP.n26 VP.n25 24.4675
R1829 VP.n30 VP.n29 24.4675
R1830 VP.n31 VP.n30 24.4675
R1831 VP.n20 VP.n19 24.4675
R1832 VP.n20 VP.n15 24.4675
R1833 VP.n50 VP.n49 12.7233
R1834 VP.n61 VP.n3 12.7233
R1835 VP.n29 VP.n13 12.7233
R1836 VP.n51 VP.n50 11.7447
R1837 VP.n58 VP.n3 11.7447
R1838 VP.n26 VP.n13 11.7447
R1839 VP.n19 VP.n18 11.7447
R1840 VP.n39 VP.n9 10.766
R1841 VP.n69 VP.n68 10.766
R1842 VP.n37 VP.n36 10.766
R1843 VP.n17 VP.n16 6.80183
R1844 VP.n38 VP.n10 0.278367
R1845 VP.n41 VP.n40 0.278367
R1846 VP.n70 VP.n0 0.278367
R1847 VP.n21 VP.n16 0.189894
R1848 VP.n22 VP.n21 0.189894
R1849 VP.n23 VP.n22 0.189894
R1850 VP.n23 VP.n14 0.189894
R1851 VP.n27 VP.n14 0.189894
R1852 VP.n28 VP.n27 0.189894
R1853 VP.n28 VP.n12 0.189894
R1854 VP.n32 VP.n12 0.189894
R1855 VP.n33 VP.n32 0.189894
R1856 VP.n34 VP.n33 0.189894
R1857 VP.n34 VP.n10 0.189894
R1858 VP.n42 VP.n41 0.189894
R1859 VP.n42 VP.n8 0.189894
R1860 VP.n46 VP.n8 0.189894
R1861 VP.n47 VP.n46 0.189894
R1862 VP.n48 VP.n47 0.189894
R1863 VP.n48 VP.n6 0.189894
R1864 VP.n53 VP.n6 0.189894
R1865 VP.n54 VP.n53 0.189894
R1866 VP.n55 VP.n54 0.189894
R1867 VP.n55 VP.n4 0.189894
R1868 VP.n59 VP.n4 0.189894
R1869 VP.n60 VP.n59 0.189894
R1870 VP.n60 VP.n2 0.189894
R1871 VP.n64 VP.n2 0.189894
R1872 VP.n65 VP.n64 0.189894
R1873 VP.n66 VP.n65 0.189894
R1874 VP.n66 VP.n0 0.189894
R1875 VP VP.n70 0.153454
R1876 VDD1 VDD1.n0 63.2399
R1877 VDD1.n3 VDD1.n2 63.1263
R1878 VDD1.n3 VDD1.n1 63.1263
R1879 VDD1.n5 VDD1.n4 61.897
R1880 VDD1.n5 VDD1.n3 46.9362
R1881 VDD1.n4 VDD1.t0 1.54136
R1882 VDD1.n4 VDD1.t6 1.54136
R1883 VDD1.n0 VDD1.t7 1.54136
R1884 VDD1.n0 VDD1.t2 1.54136
R1885 VDD1.n2 VDD1.t3 1.54136
R1886 VDD1.n2 VDD1.t4 1.54136
R1887 VDD1.n1 VDD1.t1 1.54136
R1888 VDD1.n1 VDD1.t5 1.54136
R1889 VDD1 VDD1.n5 1.22679
R1890 VTAIL.n562 VTAIL.n498 289.615
R1891 VTAIL.n66 VTAIL.n2 289.615
R1892 VTAIL.n136 VTAIL.n72 289.615
R1893 VTAIL.n208 VTAIL.n144 289.615
R1894 VTAIL.n492 VTAIL.n428 289.615
R1895 VTAIL.n420 VTAIL.n356 289.615
R1896 VTAIL.n350 VTAIL.n286 289.615
R1897 VTAIL.n278 VTAIL.n214 289.615
R1898 VTAIL.n521 VTAIL.n520 185
R1899 VTAIL.n518 VTAIL.n517 185
R1900 VTAIL.n527 VTAIL.n526 185
R1901 VTAIL.n529 VTAIL.n528 185
R1902 VTAIL.n514 VTAIL.n513 185
R1903 VTAIL.n535 VTAIL.n534 185
R1904 VTAIL.n538 VTAIL.n537 185
R1905 VTAIL.n536 VTAIL.n510 185
R1906 VTAIL.n543 VTAIL.n509 185
R1907 VTAIL.n545 VTAIL.n544 185
R1908 VTAIL.n547 VTAIL.n546 185
R1909 VTAIL.n506 VTAIL.n505 185
R1910 VTAIL.n553 VTAIL.n552 185
R1911 VTAIL.n555 VTAIL.n554 185
R1912 VTAIL.n502 VTAIL.n501 185
R1913 VTAIL.n561 VTAIL.n560 185
R1914 VTAIL.n563 VTAIL.n562 185
R1915 VTAIL.n25 VTAIL.n24 185
R1916 VTAIL.n22 VTAIL.n21 185
R1917 VTAIL.n31 VTAIL.n30 185
R1918 VTAIL.n33 VTAIL.n32 185
R1919 VTAIL.n18 VTAIL.n17 185
R1920 VTAIL.n39 VTAIL.n38 185
R1921 VTAIL.n42 VTAIL.n41 185
R1922 VTAIL.n40 VTAIL.n14 185
R1923 VTAIL.n47 VTAIL.n13 185
R1924 VTAIL.n49 VTAIL.n48 185
R1925 VTAIL.n51 VTAIL.n50 185
R1926 VTAIL.n10 VTAIL.n9 185
R1927 VTAIL.n57 VTAIL.n56 185
R1928 VTAIL.n59 VTAIL.n58 185
R1929 VTAIL.n6 VTAIL.n5 185
R1930 VTAIL.n65 VTAIL.n64 185
R1931 VTAIL.n67 VTAIL.n66 185
R1932 VTAIL.n95 VTAIL.n94 185
R1933 VTAIL.n92 VTAIL.n91 185
R1934 VTAIL.n101 VTAIL.n100 185
R1935 VTAIL.n103 VTAIL.n102 185
R1936 VTAIL.n88 VTAIL.n87 185
R1937 VTAIL.n109 VTAIL.n108 185
R1938 VTAIL.n112 VTAIL.n111 185
R1939 VTAIL.n110 VTAIL.n84 185
R1940 VTAIL.n117 VTAIL.n83 185
R1941 VTAIL.n119 VTAIL.n118 185
R1942 VTAIL.n121 VTAIL.n120 185
R1943 VTAIL.n80 VTAIL.n79 185
R1944 VTAIL.n127 VTAIL.n126 185
R1945 VTAIL.n129 VTAIL.n128 185
R1946 VTAIL.n76 VTAIL.n75 185
R1947 VTAIL.n135 VTAIL.n134 185
R1948 VTAIL.n137 VTAIL.n136 185
R1949 VTAIL.n167 VTAIL.n166 185
R1950 VTAIL.n164 VTAIL.n163 185
R1951 VTAIL.n173 VTAIL.n172 185
R1952 VTAIL.n175 VTAIL.n174 185
R1953 VTAIL.n160 VTAIL.n159 185
R1954 VTAIL.n181 VTAIL.n180 185
R1955 VTAIL.n184 VTAIL.n183 185
R1956 VTAIL.n182 VTAIL.n156 185
R1957 VTAIL.n189 VTAIL.n155 185
R1958 VTAIL.n191 VTAIL.n190 185
R1959 VTAIL.n193 VTAIL.n192 185
R1960 VTAIL.n152 VTAIL.n151 185
R1961 VTAIL.n199 VTAIL.n198 185
R1962 VTAIL.n201 VTAIL.n200 185
R1963 VTAIL.n148 VTAIL.n147 185
R1964 VTAIL.n207 VTAIL.n206 185
R1965 VTAIL.n209 VTAIL.n208 185
R1966 VTAIL.n493 VTAIL.n492 185
R1967 VTAIL.n491 VTAIL.n490 185
R1968 VTAIL.n432 VTAIL.n431 185
R1969 VTAIL.n485 VTAIL.n484 185
R1970 VTAIL.n483 VTAIL.n482 185
R1971 VTAIL.n436 VTAIL.n435 185
R1972 VTAIL.n477 VTAIL.n476 185
R1973 VTAIL.n475 VTAIL.n474 185
R1974 VTAIL.n473 VTAIL.n439 185
R1975 VTAIL.n443 VTAIL.n440 185
R1976 VTAIL.n468 VTAIL.n467 185
R1977 VTAIL.n466 VTAIL.n465 185
R1978 VTAIL.n445 VTAIL.n444 185
R1979 VTAIL.n460 VTAIL.n459 185
R1980 VTAIL.n458 VTAIL.n457 185
R1981 VTAIL.n449 VTAIL.n448 185
R1982 VTAIL.n452 VTAIL.n451 185
R1983 VTAIL.n421 VTAIL.n420 185
R1984 VTAIL.n419 VTAIL.n418 185
R1985 VTAIL.n360 VTAIL.n359 185
R1986 VTAIL.n413 VTAIL.n412 185
R1987 VTAIL.n411 VTAIL.n410 185
R1988 VTAIL.n364 VTAIL.n363 185
R1989 VTAIL.n405 VTAIL.n404 185
R1990 VTAIL.n403 VTAIL.n402 185
R1991 VTAIL.n401 VTAIL.n367 185
R1992 VTAIL.n371 VTAIL.n368 185
R1993 VTAIL.n396 VTAIL.n395 185
R1994 VTAIL.n394 VTAIL.n393 185
R1995 VTAIL.n373 VTAIL.n372 185
R1996 VTAIL.n388 VTAIL.n387 185
R1997 VTAIL.n386 VTAIL.n385 185
R1998 VTAIL.n377 VTAIL.n376 185
R1999 VTAIL.n380 VTAIL.n379 185
R2000 VTAIL.n351 VTAIL.n350 185
R2001 VTAIL.n349 VTAIL.n348 185
R2002 VTAIL.n290 VTAIL.n289 185
R2003 VTAIL.n343 VTAIL.n342 185
R2004 VTAIL.n341 VTAIL.n340 185
R2005 VTAIL.n294 VTAIL.n293 185
R2006 VTAIL.n335 VTAIL.n334 185
R2007 VTAIL.n333 VTAIL.n332 185
R2008 VTAIL.n331 VTAIL.n297 185
R2009 VTAIL.n301 VTAIL.n298 185
R2010 VTAIL.n326 VTAIL.n325 185
R2011 VTAIL.n324 VTAIL.n323 185
R2012 VTAIL.n303 VTAIL.n302 185
R2013 VTAIL.n318 VTAIL.n317 185
R2014 VTAIL.n316 VTAIL.n315 185
R2015 VTAIL.n307 VTAIL.n306 185
R2016 VTAIL.n310 VTAIL.n309 185
R2017 VTAIL.n279 VTAIL.n278 185
R2018 VTAIL.n277 VTAIL.n276 185
R2019 VTAIL.n218 VTAIL.n217 185
R2020 VTAIL.n271 VTAIL.n270 185
R2021 VTAIL.n269 VTAIL.n268 185
R2022 VTAIL.n222 VTAIL.n221 185
R2023 VTAIL.n263 VTAIL.n262 185
R2024 VTAIL.n261 VTAIL.n260 185
R2025 VTAIL.n259 VTAIL.n225 185
R2026 VTAIL.n229 VTAIL.n226 185
R2027 VTAIL.n254 VTAIL.n253 185
R2028 VTAIL.n252 VTAIL.n251 185
R2029 VTAIL.n231 VTAIL.n230 185
R2030 VTAIL.n246 VTAIL.n245 185
R2031 VTAIL.n244 VTAIL.n243 185
R2032 VTAIL.n235 VTAIL.n234 185
R2033 VTAIL.n238 VTAIL.n237 185
R2034 VTAIL.t1 VTAIL.n519 149.524
R2035 VTAIL.t6 VTAIL.n23 149.524
R2036 VTAIL.t14 VTAIL.n93 149.524
R2037 VTAIL.t13 VTAIL.n165 149.524
R2038 VTAIL.t10 VTAIL.n450 149.524
R2039 VTAIL.t11 VTAIL.n378 149.524
R2040 VTAIL.t7 VTAIL.n308 149.524
R2041 VTAIL.t5 VTAIL.n236 149.524
R2042 VTAIL.n520 VTAIL.n517 104.615
R2043 VTAIL.n527 VTAIL.n517 104.615
R2044 VTAIL.n528 VTAIL.n527 104.615
R2045 VTAIL.n528 VTAIL.n513 104.615
R2046 VTAIL.n535 VTAIL.n513 104.615
R2047 VTAIL.n537 VTAIL.n535 104.615
R2048 VTAIL.n537 VTAIL.n536 104.615
R2049 VTAIL.n536 VTAIL.n509 104.615
R2050 VTAIL.n545 VTAIL.n509 104.615
R2051 VTAIL.n546 VTAIL.n545 104.615
R2052 VTAIL.n546 VTAIL.n505 104.615
R2053 VTAIL.n553 VTAIL.n505 104.615
R2054 VTAIL.n554 VTAIL.n553 104.615
R2055 VTAIL.n554 VTAIL.n501 104.615
R2056 VTAIL.n561 VTAIL.n501 104.615
R2057 VTAIL.n562 VTAIL.n561 104.615
R2058 VTAIL.n24 VTAIL.n21 104.615
R2059 VTAIL.n31 VTAIL.n21 104.615
R2060 VTAIL.n32 VTAIL.n31 104.615
R2061 VTAIL.n32 VTAIL.n17 104.615
R2062 VTAIL.n39 VTAIL.n17 104.615
R2063 VTAIL.n41 VTAIL.n39 104.615
R2064 VTAIL.n41 VTAIL.n40 104.615
R2065 VTAIL.n40 VTAIL.n13 104.615
R2066 VTAIL.n49 VTAIL.n13 104.615
R2067 VTAIL.n50 VTAIL.n49 104.615
R2068 VTAIL.n50 VTAIL.n9 104.615
R2069 VTAIL.n57 VTAIL.n9 104.615
R2070 VTAIL.n58 VTAIL.n57 104.615
R2071 VTAIL.n58 VTAIL.n5 104.615
R2072 VTAIL.n65 VTAIL.n5 104.615
R2073 VTAIL.n66 VTAIL.n65 104.615
R2074 VTAIL.n94 VTAIL.n91 104.615
R2075 VTAIL.n101 VTAIL.n91 104.615
R2076 VTAIL.n102 VTAIL.n101 104.615
R2077 VTAIL.n102 VTAIL.n87 104.615
R2078 VTAIL.n109 VTAIL.n87 104.615
R2079 VTAIL.n111 VTAIL.n109 104.615
R2080 VTAIL.n111 VTAIL.n110 104.615
R2081 VTAIL.n110 VTAIL.n83 104.615
R2082 VTAIL.n119 VTAIL.n83 104.615
R2083 VTAIL.n120 VTAIL.n119 104.615
R2084 VTAIL.n120 VTAIL.n79 104.615
R2085 VTAIL.n127 VTAIL.n79 104.615
R2086 VTAIL.n128 VTAIL.n127 104.615
R2087 VTAIL.n128 VTAIL.n75 104.615
R2088 VTAIL.n135 VTAIL.n75 104.615
R2089 VTAIL.n136 VTAIL.n135 104.615
R2090 VTAIL.n166 VTAIL.n163 104.615
R2091 VTAIL.n173 VTAIL.n163 104.615
R2092 VTAIL.n174 VTAIL.n173 104.615
R2093 VTAIL.n174 VTAIL.n159 104.615
R2094 VTAIL.n181 VTAIL.n159 104.615
R2095 VTAIL.n183 VTAIL.n181 104.615
R2096 VTAIL.n183 VTAIL.n182 104.615
R2097 VTAIL.n182 VTAIL.n155 104.615
R2098 VTAIL.n191 VTAIL.n155 104.615
R2099 VTAIL.n192 VTAIL.n191 104.615
R2100 VTAIL.n192 VTAIL.n151 104.615
R2101 VTAIL.n199 VTAIL.n151 104.615
R2102 VTAIL.n200 VTAIL.n199 104.615
R2103 VTAIL.n200 VTAIL.n147 104.615
R2104 VTAIL.n207 VTAIL.n147 104.615
R2105 VTAIL.n208 VTAIL.n207 104.615
R2106 VTAIL.n492 VTAIL.n491 104.615
R2107 VTAIL.n491 VTAIL.n431 104.615
R2108 VTAIL.n484 VTAIL.n431 104.615
R2109 VTAIL.n484 VTAIL.n483 104.615
R2110 VTAIL.n483 VTAIL.n435 104.615
R2111 VTAIL.n476 VTAIL.n435 104.615
R2112 VTAIL.n476 VTAIL.n475 104.615
R2113 VTAIL.n475 VTAIL.n439 104.615
R2114 VTAIL.n443 VTAIL.n439 104.615
R2115 VTAIL.n467 VTAIL.n443 104.615
R2116 VTAIL.n467 VTAIL.n466 104.615
R2117 VTAIL.n466 VTAIL.n444 104.615
R2118 VTAIL.n459 VTAIL.n444 104.615
R2119 VTAIL.n459 VTAIL.n458 104.615
R2120 VTAIL.n458 VTAIL.n448 104.615
R2121 VTAIL.n451 VTAIL.n448 104.615
R2122 VTAIL.n420 VTAIL.n419 104.615
R2123 VTAIL.n419 VTAIL.n359 104.615
R2124 VTAIL.n412 VTAIL.n359 104.615
R2125 VTAIL.n412 VTAIL.n411 104.615
R2126 VTAIL.n411 VTAIL.n363 104.615
R2127 VTAIL.n404 VTAIL.n363 104.615
R2128 VTAIL.n404 VTAIL.n403 104.615
R2129 VTAIL.n403 VTAIL.n367 104.615
R2130 VTAIL.n371 VTAIL.n367 104.615
R2131 VTAIL.n395 VTAIL.n371 104.615
R2132 VTAIL.n395 VTAIL.n394 104.615
R2133 VTAIL.n394 VTAIL.n372 104.615
R2134 VTAIL.n387 VTAIL.n372 104.615
R2135 VTAIL.n387 VTAIL.n386 104.615
R2136 VTAIL.n386 VTAIL.n376 104.615
R2137 VTAIL.n379 VTAIL.n376 104.615
R2138 VTAIL.n350 VTAIL.n349 104.615
R2139 VTAIL.n349 VTAIL.n289 104.615
R2140 VTAIL.n342 VTAIL.n289 104.615
R2141 VTAIL.n342 VTAIL.n341 104.615
R2142 VTAIL.n341 VTAIL.n293 104.615
R2143 VTAIL.n334 VTAIL.n293 104.615
R2144 VTAIL.n334 VTAIL.n333 104.615
R2145 VTAIL.n333 VTAIL.n297 104.615
R2146 VTAIL.n301 VTAIL.n297 104.615
R2147 VTAIL.n325 VTAIL.n301 104.615
R2148 VTAIL.n325 VTAIL.n324 104.615
R2149 VTAIL.n324 VTAIL.n302 104.615
R2150 VTAIL.n317 VTAIL.n302 104.615
R2151 VTAIL.n317 VTAIL.n316 104.615
R2152 VTAIL.n316 VTAIL.n306 104.615
R2153 VTAIL.n309 VTAIL.n306 104.615
R2154 VTAIL.n278 VTAIL.n277 104.615
R2155 VTAIL.n277 VTAIL.n217 104.615
R2156 VTAIL.n270 VTAIL.n217 104.615
R2157 VTAIL.n270 VTAIL.n269 104.615
R2158 VTAIL.n269 VTAIL.n221 104.615
R2159 VTAIL.n262 VTAIL.n221 104.615
R2160 VTAIL.n262 VTAIL.n261 104.615
R2161 VTAIL.n261 VTAIL.n225 104.615
R2162 VTAIL.n229 VTAIL.n225 104.615
R2163 VTAIL.n253 VTAIL.n229 104.615
R2164 VTAIL.n253 VTAIL.n252 104.615
R2165 VTAIL.n252 VTAIL.n230 104.615
R2166 VTAIL.n245 VTAIL.n230 104.615
R2167 VTAIL.n245 VTAIL.n244 104.615
R2168 VTAIL.n244 VTAIL.n234 104.615
R2169 VTAIL.n237 VTAIL.n234 104.615
R2170 VTAIL.n520 VTAIL.t1 52.3082
R2171 VTAIL.n24 VTAIL.t6 52.3082
R2172 VTAIL.n94 VTAIL.t14 52.3082
R2173 VTAIL.n166 VTAIL.t13 52.3082
R2174 VTAIL.n451 VTAIL.t10 52.3082
R2175 VTAIL.n379 VTAIL.t11 52.3082
R2176 VTAIL.n309 VTAIL.t7 52.3082
R2177 VTAIL.n237 VTAIL.t5 52.3082
R2178 VTAIL.n427 VTAIL.n426 45.2184
R2179 VTAIL.n285 VTAIL.n284 45.2184
R2180 VTAIL.n1 VTAIL.n0 45.2184
R2181 VTAIL.n143 VTAIL.n142 45.2184
R2182 VTAIL.n567 VTAIL.n566 32.3793
R2183 VTAIL.n71 VTAIL.n70 32.3793
R2184 VTAIL.n141 VTAIL.n140 32.3793
R2185 VTAIL.n213 VTAIL.n212 32.3793
R2186 VTAIL.n497 VTAIL.n496 32.3793
R2187 VTAIL.n425 VTAIL.n424 32.3793
R2188 VTAIL.n355 VTAIL.n354 32.3793
R2189 VTAIL.n283 VTAIL.n282 32.3793
R2190 VTAIL.n567 VTAIL.n497 26.0134
R2191 VTAIL.n283 VTAIL.n213 26.0134
R2192 VTAIL.n544 VTAIL.n543 13.1884
R2193 VTAIL.n48 VTAIL.n47 13.1884
R2194 VTAIL.n118 VTAIL.n117 13.1884
R2195 VTAIL.n190 VTAIL.n189 13.1884
R2196 VTAIL.n474 VTAIL.n473 13.1884
R2197 VTAIL.n402 VTAIL.n401 13.1884
R2198 VTAIL.n332 VTAIL.n331 13.1884
R2199 VTAIL.n260 VTAIL.n259 13.1884
R2200 VTAIL.n542 VTAIL.n510 12.8005
R2201 VTAIL.n547 VTAIL.n508 12.8005
R2202 VTAIL.n46 VTAIL.n14 12.8005
R2203 VTAIL.n51 VTAIL.n12 12.8005
R2204 VTAIL.n116 VTAIL.n84 12.8005
R2205 VTAIL.n121 VTAIL.n82 12.8005
R2206 VTAIL.n188 VTAIL.n156 12.8005
R2207 VTAIL.n193 VTAIL.n154 12.8005
R2208 VTAIL.n477 VTAIL.n438 12.8005
R2209 VTAIL.n472 VTAIL.n440 12.8005
R2210 VTAIL.n405 VTAIL.n366 12.8005
R2211 VTAIL.n400 VTAIL.n368 12.8005
R2212 VTAIL.n335 VTAIL.n296 12.8005
R2213 VTAIL.n330 VTAIL.n298 12.8005
R2214 VTAIL.n263 VTAIL.n224 12.8005
R2215 VTAIL.n258 VTAIL.n226 12.8005
R2216 VTAIL.n539 VTAIL.n538 12.0247
R2217 VTAIL.n548 VTAIL.n506 12.0247
R2218 VTAIL.n43 VTAIL.n42 12.0247
R2219 VTAIL.n52 VTAIL.n10 12.0247
R2220 VTAIL.n113 VTAIL.n112 12.0247
R2221 VTAIL.n122 VTAIL.n80 12.0247
R2222 VTAIL.n185 VTAIL.n184 12.0247
R2223 VTAIL.n194 VTAIL.n152 12.0247
R2224 VTAIL.n478 VTAIL.n436 12.0247
R2225 VTAIL.n469 VTAIL.n468 12.0247
R2226 VTAIL.n406 VTAIL.n364 12.0247
R2227 VTAIL.n397 VTAIL.n396 12.0247
R2228 VTAIL.n336 VTAIL.n294 12.0247
R2229 VTAIL.n327 VTAIL.n326 12.0247
R2230 VTAIL.n264 VTAIL.n222 12.0247
R2231 VTAIL.n255 VTAIL.n254 12.0247
R2232 VTAIL.n534 VTAIL.n512 11.249
R2233 VTAIL.n552 VTAIL.n551 11.249
R2234 VTAIL.n38 VTAIL.n16 11.249
R2235 VTAIL.n56 VTAIL.n55 11.249
R2236 VTAIL.n108 VTAIL.n86 11.249
R2237 VTAIL.n126 VTAIL.n125 11.249
R2238 VTAIL.n180 VTAIL.n158 11.249
R2239 VTAIL.n198 VTAIL.n197 11.249
R2240 VTAIL.n482 VTAIL.n481 11.249
R2241 VTAIL.n465 VTAIL.n442 11.249
R2242 VTAIL.n410 VTAIL.n409 11.249
R2243 VTAIL.n393 VTAIL.n370 11.249
R2244 VTAIL.n340 VTAIL.n339 11.249
R2245 VTAIL.n323 VTAIL.n300 11.249
R2246 VTAIL.n268 VTAIL.n267 11.249
R2247 VTAIL.n251 VTAIL.n228 11.249
R2248 VTAIL.n533 VTAIL.n514 10.4732
R2249 VTAIL.n555 VTAIL.n504 10.4732
R2250 VTAIL.n37 VTAIL.n18 10.4732
R2251 VTAIL.n59 VTAIL.n8 10.4732
R2252 VTAIL.n107 VTAIL.n88 10.4732
R2253 VTAIL.n129 VTAIL.n78 10.4732
R2254 VTAIL.n179 VTAIL.n160 10.4732
R2255 VTAIL.n201 VTAIL.n150 10.4732
R2256 VTAIL.n485 VTAIL.n434 10.4732
R2257 VTAIL.n464 VTAIL.n445 10.4732
R2258 VTAIL.n413 VTAIL.n362 10.4732
R2259 VTAIL.n392 VTAIL.n373 10.4732
R2260 VTAIL.n343 VTAIL.n292 10.4732
R2261 VTAIL.n322 VTAIL.n303 10.4732
R2262 VTAIL.n271 VTAIL.n220 10.4732
R2263 VTAIL.n250 VTAIL.n231 10.4732
R2264 VTAIL.n521 VTAIL.n519 10.2747
R2265 VTAIL.n25 VTAIL.n23 10.2747
R2266 VTAIL.n95 VTAIL.n93 10.2747
R2267 VTAIL.n167 VTAIL.n165 10.2747
R2268 VTAIL.n452 VTAIL.n450 10.2747
R2269 VTAIL.n380 VTAIL.n378 10.2747
R2270 VTAIL.n310 VTAIL.n308 10.2747
R2271 VTAIL.n238 VTAIL.n236 10.2747
R2272 VTAIL.n530 VTAIL.n529 9.69747
R2273 VTAIL.n556 VTAIL.n502 9.69747
R2274 VTAIL.n34 VTAIL.n33 9.69747
R2275 VTAIL.n60 VTAIL.n6 9.69747
R2276 VTAIL.n104 VTAIL.n103 9.69747
R2277 VTAIL.n130 VTAIL.n76 9.69747
R2278 VTAIL.n176 VTAIL.n175 9.69747
R2279 VTAIL.n202 VTAIL.n148 9.69747
R2280 VTAIL.n486 VTAIL.n432 9.69747
R2281 VTAIL.n461 VTAIL.n460 9.69747
R2282 VTAIL.n414 VTAIL.n360 9.69747
R2283 VTAIL.n389 VTAIL.n388 9.69747
R2284 VTAIL.n344 VTAIL.n290 9.69747
R2285 VTAIL.n319 VTAIL.n318 9.69747
R2286 VTAIL.n272 VTAIL.n218 9.69747
R2287 VTAIL.n247 VTAIL.n246 9.69747
R2288 VTAIL.n566 VTAIL.n565 9.45567
R2289 VTAIL.n70 VTAIL.n69 9.45567
R2290 VTAIL.n140 VTAIL.n139 9.45567
R2291 VTAIL.n212 VTAIL.n211 9.45567
R2292 VTAIL.n496 VTAIL.n495 9.45567
R2293 VTAIL.n424 VTAIL.n423 9.45567
R2294 VTAIL.n354 VTAIL.n353 9.45567
R2295 VTAIL.n282 VTAIL.n281 9.45567
R2296 VTAIL.n500 VTAIL.n499 9.3005
R2297 VTAIL.n559 VTAIL.n558 9.3005
R2298 VTAIL.n557 VTAIL.n556 9.3005
R2299 VTAIL.n504 VTAIL.n503 9.3005
R2300 VTAIL.n551 VTAIL.n550 9.3005
R2301 VTAIL.n549 VTAIL.n548 9.3005
R2302 VTAIL.n508 VTAIL.n507 9.3005
R2303 VTAIL.n523 VTAIL.n522 9.3005
R2304 VTAIL.n525 VTAIL.n524 9.3005
R2305 VTAIL.n516 VTAIL.n515 9.3005
R2306 VTAIL.n531 VTAIL.n530 9.3005
R2307 VTAIL.n533 VTAIL.n532 9.3005
R2308 VTAIL.n512 VTAIL.n511 9.3005
R2309 VTAIL.n540 VTAIL.n539 9.3005
R2310 VTAIL.n542 VTAIL.n541 9.3005
R2311 VTAIL.n565 VTAIL.n564 9.3005
R2312 VTAIL.n4 VTAIL.n3 9.3005
R2313 VTAIL.n63 VTAIL.n62 9.3005
R2314 VTAIL.n61 VTAIL.n60 9.3005
R2315 VTAIL.n8 VTAIL.n7 9.3005
R2316 VTAIL.n55 VTAIL.n54 9.3005
R2317 VTAIL.n53 VTAIL.n52 9.3005
R2318 VTAIL.n12 VTAIL.n11 9.3005
R2319 VTAIL.n27 VTAIL.n26 9.3005
R2320 VTAIL.n29 VTAIL.n28 9.3005
R2321 VTAIL.n20 VTAIL.n19 9.3005
R2322 VTAIL.n35 VTAIL.n34 9.3005
R2323 VTAIL.n37 VTAIL.n36 9.3005
R2324 VTAIL.n16 VTAIL.n15 9.3005
R2325 VTAIL.n44 VTAIL.n43 9.3005
R2326 VTAIL.n46 VTAIL.n45 9.3005
R2327 VTAIL.n69 VTAIL.n68 9.3005
R2328 VTAIL.n74 VTAIL.n73 9.3005
R2329 VTAIL.n133 VTAIL.n132 9.3005
R2330 VTAIL.n131 VTAIL.n130 9.3005
R2331 VTAIL.n78 VTAIL.n77 9.3005
R2332 VTAIL.n125 VTAIL.n124 9.3005
R2333 VTAIL.n123 VTAIL.n122 9.3005
R2334 VTAIL.n82 VTAIL.n81 9.3005
R2335 VTAIL.n97 VTAIL.n96 9.3005
R2336 VTAIL.n99 VTAIL.n98 9.3005
R2337 VTAIL.n90 VTAIL.n89 9.3005
R2338 VTAIL.n105 VTAIL.n104 9.3005
R2339 VTAIL.n107 VTAIL.n106 9.3005
R2340 VTAIL.n86 VTAIL.n85 9.3005
R2341 VTAIL.n114 VTAIL.n113 9.3005
R2342 VTAIL.n116 VTAIL.n115 9.3005
R2343 VTAIL.n139 VTAIL.n138 9.3005
R2344 VTAIL.n146 VTAIL.n145 9.3005
R2345 VTAIL.n205 VTAIL.n204 9.3005
R2346 VTAIL.n203 VTAIL.n202 9.3005
R2347 VTAIL.n150 VTAIL.n149 9.3005
R2348 VTAIL.n197 VTAIL.n196 9.3005
R2349 VTAIL.n195 VTAIL.n194 9.3005
R2350 VTAIL.n154 VTAIL.n153 9.3005
R2351 VTAIL.n169 VTAIL.n168 9.3005
R2352 VTAIL.n171 VTAIL.n170 9.3005
R2353 VTAIL.n162 VTAIL.n161 9.3005
R2354 VTAIL.n177 VTAIL.n176 9.3005
R2355 VTAIL.n179 VTAIL.n178 9.3005
R2356 VTAIL.n158 VTAIL.n157 9.3005
R2357 VTAIL.n186 VTAIL.n185 9.3005
R2358 VTAIL.n188 VTAIL.n187 9.3005
R2359 VTAIL.n211 VTAIL.n210 9.3005
R2360 VTAIL.n454 VTAIL.n453 9.3005
R2361 VTAIL.n456 VTAIL.n455 9.3005
R2362 VTAIL.n447 VTAIL.n446 9.3005
R2363 VTAIL.n462 VTAIL.n461 9.3005
R2364 VTAIL.n464 VTAIL.n463 9.3005
R2365 VTAIL.n442 VTAIL.n441 9.3005
R2366 VTAIL.n470 VTAIL.n469 9.3005
R2367 VTAIL.n472 VTAIL.n471 9.3005
R2368 VTAIL.n495 VTAIL.n494 9.3005
R2369 VTAIL.n430 VTAIL.n429 9.3005
R2370 VTAIL.n489 VTAIL.n488 9.3005
R2371 VTAIL.n487 VTAIL.n486 9.3005
R2372 VTAIL.n434 VTAIL.n433 9.3005
R2373 VTAIL.n481 VTAIL.n480 9.3005
R2374 VTAIL.n479 VTAIL.n478 9.3005
R2375 VTAIL.n438 VTAIL.n437 9.3005
R2376 VTAIL.n382 VTAIL.n381 9.3005
R2377 VTAIL.n384 VTAIL.n383 9.3005
R2378 VTAIL.n375 VTAIL.n374 9.3005
R2379 VTAIL.n390 VTAIL.n389 9.3005
R2380 VTAIL.n392 VTAIL.n391 9.3005
R2381 VTAIL.n370 VTAIL.n369 9.3005
R2382 VTAIL.n398 VTAIL.n397 9.3005
R2383 VTAIL.n400 VTAIL.n399 9.3005
R2384 VTAIL.n423 VTAIL.n422 9.3005
R2385 VTAIL.n358 VTAIL.n357 9.3005
R2386 VTAIL.n417 VTAIL.n416 9.3005
R2387 VTAIL.n415 VTAIL.n414 9.3005
R2388 VTAIL.n362 VTAIL.n361 9.3005
R2389 VTAIL.n409 VTAIL.n408 9.3005
R2390 VTAIL.n407 VTAIL.n406 9.3005
R2391 VTAIL.n366 VTAIL.n365 9.3005
R2392 VTAIL.n312 VTAIL.n311 9.3005
R2393 VTAIL.n314 VTAIL.n313 9.3005
R2394 VTAIL.n305 VTAIL.n304 9.3005
R2395 VTAIL.n320 VTAIL.n319 9.3005
R2396 VTAIL.n322 VTAIL.n321 9.3005
R2397 VTAIL.n300 VTAIL.n299 9.3005
R2398 VTAIL.n328 VTAIL.n327 9.3005
R2399 VTAIL.n330 VTAIL.n329 9.3005
R2400 VTAIL.n353 VTAIL.n352 9.3005
R2401 VTAIL.n288 VTAIL.n287 9.3005
R2402 VTAIL.n347 VTAIL.n346 9.3005
R2403 VTAIL.n345 VTAIL.n344 9.3005
R2404 VTAIL.n292 VTAIL.n291 9.3005
R2405 VTAIL.n339 VTAIL.n338 9.3005
R2406 VTAIL.n337 VTAIL.n336 9.3005
R2407 VTAIL.n296 VTAIL.n295 9.3005
R2408 VTAIL.n240 VTAIL.n239 9.3005
R2409 VTAIL.n242 VTAIL.n241 9.3005
R2410 VTAIL.n233 VTAIL.n232 9.3005
R2411 VTAIL.n248 VTAIL.n247 9.3005
R2412 VTAIL.n250 VTAIL.n249 9.3005
R2413 VTAIL.n228 VTAIL.n227 9.3005
R2414 VTAIL.n256 VTAIL.n255 9.3005
R2415 VTAIL.n258 VTAIL.n257 9.3005
R2416 VTAIL.n281 VTAIL.n280 9.3005
R2417 VTAIL.n216 VTAIL.n215 9.3005
R2418 VTAIL.n275 VTAIL.n274 9.3005
R2419 VTAIL.n273 VTAIL.n272 9.3005
R2420 VTAIL.n220 VTAIL.n219 9.3005
R2421 VTAIL.n267 VTAIL.n266 9.3005
R2422 VTAIL.n265 VTAIL.n264 9.3005
R2423 VTAIL.n224 VTAIL.n223 9.3005
R2424 VTAIL.n526 VTAIL.n516 8.92171
R2425 VTAIL.n560 VTAIL.n559 8.92171
R2426 VTAIL.n30 VTAIL.n20 8.92171
R2427 VTAIL.n64 VTAIL.n63 8.92171
R2428 VTAIL.n100 VTAIL.n90 8.92171
R2429 VTAIL.n134 VTAIL.n133 8.92171
R2430 VTAIL.n172 VTAIL.n162 8.92171
R2431 VTAIL.n206 VTAIL.n205 8.92171
R2432 VTAIL.n490 VTAIL.n489 8.92171
R2433 VTAIL.n457 VTAIL.n447 8.92171
R2434 VTAIL.n418 VTAIL.n417 8.92171
R2435 VTAIL.n385 VTAIL.n375 8.92171
R2436 VTAIL.n348 VTAIL.n347 8.92171
R2437 VTAIL.n315 VTAIL.n305 8.92171
R2438 VTAIL.n276 VTAIL.n275 8.92171
R2439 VTAIL.n243 VTAIL.n233 8.92171
R2440 VTAIL.n525 VTAIL.n518 8.14595
R2441 VTAIL.n563 VTAIL.n500 8.14595
R2442 VTAIL.n29 VTAIL.n22 8.14595
R2443 VTAIL.n67 VTAIL.n4 8.14595
R2444 VTAIL.n99 VTAIL.n92 8.14595
R2445 VTAIL.n137 VTAIL.n74 8.14595
R2446 VTAIL.n171 VTAIL.n164 8.14595
R2447 VTAIL.n209 VTAIL.n146 8.14595
R2448 VTAIL.n493 VTAIL.n430 8.14595
R2449 VTAIL.n456 VTAIL.n449 8.14595
R2450 VTAIL.n421 VTAIL.n358 8.14595
R2451 VTAIL.n384 VTAIL.n377 8.14595
R2452 VTAIL.n351 VTAIL.n288 8.14595
R2453 VTAIL.n314 VTAIL.n307 8.14595
R2454 VTAIL.n279 VTAIL.n216 8.14595
R2455 VTAIL.n242 VTAIL.n235 8.14595
R2456 VTAIL.n522 VTAIL.n521 7.3702
R2457 VTAIL.n564 VTAIL.n498 7.3702
R2458 VTAIL.n26 VTAIL.n25 7.3702
R2459 VTAIL.n68 VTAIL.n2 7.3702
R2460 VTAIL.n96 VTAIL.n95 7.3702
R2461 VTAIL.n138 VTAIL.n72 7.3702
R2462 VTAIL.n168 VTAIL.n167 7.3702
R2463 VTAIL.n210 VTAIL.n144 7.3702
R2464 VTAIL.n494 VTAIL.n428 7.3702
R2465 VTAIL.n453 VTAIL.n452 7.3702
R2466 VTAIL.n422 VTAIL.n356 7.3702
R2467 VTAIL.n381 VTAIL.n380 7.3702
R2468 VTAIL.n352 VTAIL.n286 7.3702
R2469 VTAIL.n311 VTAIL.n310 7.3702
R2470 VTAIL.n280 VTAIL.n214 7.3702
R2471 VTAIL.n239 VTAIL.n238 7.3702
R2472 VTAIL.n566 VTAIL.n498 6.59444
R2473 VTAIL.n70 VTAIL.n2 6.59444
R2474 VTAIL.n140 VTAIL.n72 6.59444
R2475 VTAIL.n212 VTAIL.n144 6.59444
R2476 VTAIL.n496 VTAIL.n428 6.59444
R2477 VTAIL.n424 VTAIL.n356 6.59444
R2478 VTAIL.n354 VTAIL.n286 6.59444
R2479 VTAIL.n282 VTAIL.n214 6.59444
R2480 VTAIL.n522 VTAIL.n518 5.81868
R2481 VTAIL.n564 VTAIL.n563 5.81868
R2482 VTAIL.n26 VTAIL.n22 5.81868
R2483 VTAIL.n68 VTAIL.n67 5.81868
R2484 VTAIL.n96 VTAIL.n92 5.81868
R2485 VTAIL.n138 VTAIL.n137 5.81868
R2486 VTAIL.n168 VTAIL.n164 5.81868
R2487 VTAIL.n210 VTAIL.n209 5.81868
R2488 VTAIL.n494 VTAIL.n493 5.81868
R2489 VTAIL.n453 VTAIL.n449 5.81868
R2490 VTAIL.n422 VTAIL.n421 5.81868
R2491 VTAIL.n381 VTAIL.n377 5.81868
R2492 VTAIL.n352 VTAIL.n351 5.81868
R2493 VTAIL.n311 VTAIL.n307 5.81868
R2494 VTAIL.n280 VTAIL.n279 5.81868
R2495 VTAIL.n239 VTAIL.n235 5.81868
R2496 VTAIL.n526 VTAIL.n525 5.04292
R2497 VTAIL.n560 VTAIL.n500 5.04292
R2498 VTAIL.n30 VTAIL.n29 5.04292
R2499 VTAIL.n64 VTAIL.n4 5.04292
R2500 VTAIL.n100 VTAIL.n99 5.04292
R2501 VTAIL.n134 VTAIL.n74 5.04292
R2502 VTAIL.n172 VTAIL.n171 5.04292
R2503 VTAIL.n206 VTAIL.n146 5.04292
R2504 VTAIL.n490 VTAIL.n430 5.04292
R2505 VTAIL.n457 VTAIL.n456 5.04292
R2506 VTAIL.n418 VTAIL.n358 5.04292
R2507 VTAIL.n385 VTAIL.n384 5.04292
R2508 VTAIL.n348 VTAIL.n288 5.04292
R2509 VTAIL.n315 VTAIL.n314 5.04292
R2510 VTAIL.n276 VTAIL.n216 5.04292
R2511 VTAIL.n243 VTAIL.n242 5.04292
R2512 VTAIL.n529 VTAIL.n516 4.26717
R2513 VTAIL.n559 VTAIL.n502 4.26717
R2514 VTAIL.n33 VTAIL.n20 4.26717
R2515 VTAIL.n63 VTAIL.n6 4.26717
R2516 VTAIL.n103 VTAIL.n90 4.26717
R2517 VTAIL.n133 VTAIL.n76 4.26717
R2518 VTAIL.n175 VTAIL.n162 4.26717
R2519 VTAIL.n205 VTAIL.n148 4.26717
R2520 VTAIL.n489 VTAIL.n432 4.26717
R2521 VTAIL.n460 VTAIL.n447 4.26717
R2522 VTAIL.n417 VTAIL.n360 4.26717
R2523 VTAIL.n388 VTAIL.n375 4.26717
R2524 VTAIL.n347 VTAIL.n290 4.26717
R2525 VTAIL.n318 VTAIL.n305 4.26717
R2526 VTAIL.n275 VTAIL.n218 4.26717
R2527 VTAIL.n246 VTAIL.n233 4.26717
R2528 VTAIL.n530 VTAIL.n514 3.49141
R2529 VTAIL.n556 VTAIL.n555 3.49141
R2530 VTAIL.n34 VTAIL.n18 3.49141
R2531 VTAIL.n60 VTAIL.n59 3.49141
R2532 VTAIL.n104 VTAIL.n88 3.49141
R2533 VTAIL.n130 VTAIL.n129 3.49141
R2534 VTAIL.n176 VTAIL.n160 3.49141
R2535 VTAIL.n202 VTAIL.n201 3.49141
R2536 VTAIL.n486 VTAIL.n485 3.49141
R2537 VTAIL.n461 VTAIL.n445 3.49141
R2538 VTAIL.n414 VTAIL.n413 3.49141
R2539 VTAIL.n389 VTAIL.n373 3.49141
R2540 VTAIL.n344 VTAIL.n343 3.49141
R2541 VTAIL.n319 VTAIL.n303 3.49141
R2542 VTAIL.n272 VTAIL.n271 3.49141
R2543 VTAIL.n247 VTAIL.n231 3.49141
R2544 VTAIL.n523 VTAIL.n519 2.84303
R2545 VTAIL.n27 VTAIL.n23 2.84303
R2546 VTAIL.n97 VTAIL.n93 2.84303
R2547 VTAIL.n169 VTAIL.n165 2.84303
R2548 VTAIL.n454 VTAIL.n450 2.84303
R2549 VTAIL.n382 VTAIL.n378 2.84303
R2550 VTAIL.n312 VTAIL.n308 2.84303
R2551 VTAIL.n240 VTAIL.n236 2.84303
R2552 VTAIL.n534 VTAIL.n533 2.71565
R2553 VTAIL.n552 VTAIL.n504 2.71565
R2554 VTAIL.n38 VTAIL.n37 2.71565
R2555 VTAIL.n56 VTAIL.n8 2.71565
R2556 VTAIL.n108 VTAIL.n107 2.71565
R2557 VTAIL.n126 VTAIL.n78 2.71565
R2558 VTAIL.n180 VTAIL.n179 2.71565
R2559 VTAIL.n198 VTAIL.n150 2.71565
R2560 VTAIL.n482 VTAIL.n434 2.71565
R2561 VTAIL.n465 VTAIL.n464 2.71565
R2562 VTAIL.n410 VTAIL.n362 2.71565
R2563 VTAIL.n393 VTAIL.n392 2.71565
R2564 VTAIL.n340 VTAIL.n292 2.71565
R2565 VTAIL.n323 VTAIL.n322 2.71565
R2566 VTAIL.n268 VTAIL.n220 2.71565
R2567 VTAIL.n251 VTAIL.n250 2.71565
R2568 VTAIL.n285 VTAIL.n283 2.56947
R2569 VTAIL.n355 VTAIL.n285 2.56947
R2570 VTAIL.n427 VTAIL.n425 2.56947
R2571 VTAIL.n497 VTAIL.n427 2.56947
R2572 VTAIL.n213 VTAIL.n143 2.56947
R2573 VTAIL.n143 VTAIL.n141 2.56947
R2574 VTAIL.n71 VTAIL.n1 2.56947
R2575 VTAIL VTAIL.n567 2.51128
R2576 VTAIL.n538 VTAIL.n512 1.93989
R2577 VTAIL.n551 VTAIL.n506 1.93989
R2578 VTAIL.n42 VTAIL.n16 1.93989
R2579 VTAIL.n55 VTAIL.n10 1.93989
R2580 VTAIL.n112 VTAIL.n86 1.93989
R2581 VTAIL.n125 VTAIL.n80 1.93989
R2582 VTAIL.n184 VTAIL.n158 1.93989
R2583 VTAIL.n197 VTAIL.n152 1.93989
R2584 VTAIL.n481 VTAIL.n436 1.93989
R2585 VTAIL.n468 VTAIL.n442 1.93989
R2586 VTAIL.n409 VTAIL.n364 1.93989
R2587 VTAIL.n396 VTAIL.n370 1.93989
R2588 VTAIL.n339 VTAIL.n294 1.93989
R2589 VTAIL.n326 VTAIL.n300 1.93989
R2590 VTAIL.n267 VTAIL.n222 1.93989
R2591 VTAIL.n254 VTAIL.n228 1.93989
R2592 VTAIL.n0 VTAIL.t4 1.54136
R2593 VTAIL.n0 VTAIL.t0 1.54136
R2594 VTAIL.n142 VTAIL.t9 1.54136
R2595 VTAIL.n142 VTAIL.t15 1.54136
R2596 VTAIL.n426 VTAIL.t8 1.54136
R2597 VTAIL.n426 VTAIL.t12 1.54136
R2598 VTAIL.n284 VTAIL.t3 1.54136
R2599 VTAIL.n284 VTAIL.t2 1.54136
R2600 VTAIL.n539 VTAIL.n510 1.16414
R2601 VTAIL.n548 VTAIL.n547 1.16414
R2602 VTAIL.n43 VTAIL.n14 1.16414
R2603 VTAIL.n52 VTAIL.n51 1.16414
R2604 VTAIL.n113 VTAIL.n84 1.16414
R2605 VTAIL.n122 VTAIL.n121 1.16414
R2606 VTAIL.n185 VTAIL.n156 1.16414
R2607 VTAIL.n194 VTAIL.n193 1.16414
R2608 VTAIL.n478 VTAIL.n477 1.16414
R2609 VTAIL.n469 VTAIL.n440 1.16414
R2610 VTAIL.n406 VTAIL.n405 1.16414
R2611 VTAIL.n397 VTAIL.n368 1.16414
R2612 VTAIL.n336 VTAIL.n335 1.16414
R2613 VTAIL.n327 VTAIL.n298 1.16414
R2614 VTAIL.n264 VTAIL.n263 1.16414
R2615 VTAIL.n255 VTAIL.n226 1.16414
R2616 VTAIL.n425 VTAIL.n355 0.470328
R2617 VTAIL.n141 VTAIL.n71 0.470328
R2618 VTAIL.n543 VTAIL.n542 0.388379
R2619 VTAIL.n544 VTAIL.n508 0.388379
R2620 VTAIL.n47 VTAIL.n46 0.388379
R2621 VTAIL.n48 VTAIL.n12 0.388379
R2622 VTAIL.n117 VTAIL.n116 0.388379
R2623 VTAIL.n118 VTAIL.n82 0.388379
R2624 VTAIL.n189 VTAIL.n188 0.388379
R2625 VTAIL.n190 VTAIL.n154 0.388379
R2626 VTAIL.n474 VTAIL.n438 0.388379
R2627 VTAIL.n473 VTAIL.n472 0.388379
R2628 VTAIL.n402 VTAIL.n366 0.388379
R2629 VTAIL.n401 VTAIL.n400 0.388379
R2630 VTAIL.n332 VTAIL.n296 0.388379
R2631 VTAIL.n331 VTAIL.n330 0.388379
R2632 VTAIL.n260 VTAIL.n224 0.388379
R2633 VTAIL.n259 VTAIL.n258 0.388379
R2634 VTAIL.n524 VTAIL.n523 0.155672
R2635 VTAIL.n524 VTAIL.n515 0.155672
R2636 VTAIL.n531 VTAIL.n515 0.155672
R2637 VTAIL.n532 VTAIL.n531 0.155672
R2638 VTAIL.n532 VTAIL.n511 0.155672
R2639 VTAIL.n540 VTAIL.n511 0.155672
R2640 VTAIL.n541 VTAIL.n540 0.155672
R2641 VTAIL.n541 VTAIL.n507 0.155672
R2642 VTAIL.n549 VTAIL.n507 0.155672
R2643 VTAIL.n550 VTAIL.n549 0.155672
R2644 VTAIL.n550 VTAIL.n503 0.155672
R2645 VTAIL.n557 VTAIL.n503 0.155672
R2646 VTAIL.n558 VTAIL.n557 0.155672
R2647 VTAIL.n558 VTAIL.n499 0.155672
R2648 VTAIL.n565 VTAIL.n499 0.155672
R2649 VTAIL.n28 VTAIL.n27 0.155672
R2650 VTAIL.n28 VTAIL.n19 0.155672
R2651 VTAIL.n35 VTAIL.n19 0.155672
R2652 VTAIL.n36 VTAIL.n35 0.155672
R2653 VTAIL.n36 VTAIL.n15 0.155672
R2654 VTAIL.n44 VTAIL.n15 0.155672
R2655 VTAIL.n45 VTAIL.n44 0.155672
R2656 VTAIL.n45 VTAIL.n11 0.155672
R2657 VTAIL.n53 VTAIL.n11 0.155672
R2658 VTAIL.n54 VTAIL.n53 0.155672
R2659 VTAIL.n54 VTAIL.n7 0.155672
R2660 VTAIL.n61 VTAIL.n7 0.155672
R2661 VTAIL.n62 VTAIL.n61 0.155672
R2662 VTAIL.n62 VTAIL.n3 0.155672
R2663 VTAIL.n69 VTAIL.n3 0.155672
R2664 VTAIL.n98 VTAIL.n97 0.155672
R2665 VTAIL.n98 VTAIL.n89 0.155672
R2666 VTAIL.n105 VTAIL.n89 0.155672
R2667 VTAIL.n106 VTAIL.n105 0.155672
R2668 VTAIL.n106 VTAIL.n85 0.155672
R2669 VTAIL.n114 VTAIL.n85 0.155672
R2670 VTAIL.n115 VTAIL.n114 0.155672
R2671 VTAIL.n115 VTAIL.n81 0.155672
R2672 VTAIL.n123 VTAIL.n81 0.155672
R2673 VTAIL.n124 VTAIL.n123 0.155672
R2674 VTAIL.n124 VTAIL.n77 0.155672
R2675 VTAIL.n131 VTAIL.n77 0.155672
R2676 VTAIL.n132 VTAIL.n131 0.155672
R2677 VTAIL.n132 VTAIL.n73 0.155672
R2678 VTAIL.n139 VTAIL.n73 0.155672
R2679 VTAIL.n170 VTAIL.n169 0.155672
R2680 VTAIL.n170 VTAIL.n161 0.155672
R2681 VTAIL.n177 VTAIL.n161 0.155672
R2682 VTAIL.n178 VTAIL.n177 0.155672
R2683 VTAIL.n178 VTAIL.n157 0.155672
R2684 VTAIL.n186 VTAIL.n157 0.155672
R2685 VTAIL.n187 VTAIL.n186 0.155672
R2686 VTAIL.n187 VTAIL.n153 0.155672
R2687 VTAIL.n195 VTAIL.n153 0.155672
R2688 VTAIL.n196 VTAIL.n195 0.155672
R2689 VTAIL.n196 VTAIL.n149 0.155672
R2690 VTAIL.n203 VTAIL.n149 0.155672
R2691 VTAIL.n204 VTAIL.n203 0.155672
R2692 VTAIL.n204 VTAIL.n145 0.155672
R2693 VTAIL.n211 VTAIL.n145 0.155672
R2694 VTAIL.n495 VTAIL.n429 0.155672
R2695 VTAIL.n488 VTAIL.n429 0.155672
R2696 VTAIL.n488 VTAIL.n487 0.155672
R2697 VTAIL.n487 VTAIL.n433 0.155672
R2698 VTAIL.n480 VTAIL.n433 0.155672
R2699 VTAIL.n480 VTAIL.n479 0.155672
R2700 VTAIL.n479 VTAIL.n437 0.155672
R2701 VTAIL.n471 VTAIL.n437 0.155672
R2702 VTAIL.n471 VTAIL.n470 0.155672
R2703 VTAIL.n470 VTAIL.n441 0.155672
R2704 VTAIL.n463 VTAIL.n441 0.155672
R2705 VTAIL.n463 VTAIL.n462 0.155672
R2706 VTAIL.n462 VTAIL.n446 0.155672
R2707 VTAIL.n455 VTAIL.n446 0.155672
R2708 VTAIL.n455 VTAIL.n454 0.155672
R2709 VTAIL.n423 VTAIL.n357 0.155672
R2710 VTAIL.n416 VTAIL.n357 0.155672
R2711 VTAIL.n416 VTAIL.n415 0.155672
R2712 VTAIL.n415 VTAIL.n361 0.155672
R2713 VTAIL.n408 VTAIL.n361 0.155672
R2714 VTAIL.n408 VTAIL.n407 0.155672
R2715 VTAIL.n407 VTAIL.n365 0.155672
R2716 VTAIL.n399 VTAIL.n365 0.155672
R2717 VTAIL.n399 VTAIL.n398 0.155672
R2718 VTAIL.n398 VTAIL.n369 0.155672
R2719 VTAIL.n391 VTAIL.n369 0.155672
R2720 VTAIL.n391 VTAIL.n390 0.155672
R2721 VTAIL.n390 VTAIL.n374 0.155672
R2722 VTAIL.n383 VTAIL.n374 0.155672
R2723 VTAIL.n383 VTAIL.n382 0.155672
R2724 VTAIL.n353 VTAIL.n287 0.155672
R2725 VTAIL.n346 VTAIL.n287 0.155672
R2726 VTAIL.n346 VTAIL.n345 0.155672
R2727 VTAIL.n345 VTAIL.n291 0.155672
R2728 VTAIL.n338 VTAIL.n291 0.155672
R2729 VTAIL.n338 VTAIL.n337 0.155672
R2730 VTAIL.n337 VTAIL.n295 0.155672
R2731 VTAIL.n329 VTAIL.n295 0.155672
R2732 VTAIL.n329 VTAIL.n328 0.155672
R2733 VTAIL.n328 VTAIL.n299 0.155672
R2734 VTAIL.n321 VTAIL.n299 0.155672
R2735 VTAIL.n321 VTAIL.n320 0.155672
R2736 VTAIL.n320 VTAIL.n304 0.155672
R2737 VTAIL.n313 VTAIL.n304 0.155672
R2738 VTAIL.n313 VTAIL.n312 0.155672
R2739 VTAIL.n281 VTAIL.n215 0.155672
R2740 VTAIL.n274 VTAIL.n215 0.155672
R2741 VTAIL.n274 VTAIL.n273 0.155672
R2742 VTAIL.n273 VTAIL.n219 0.155672
R2743 VTAIL.n266 VTAIL.n219 0.155672
R2744 VTAIL.n266 VTAIL.n265 0.155672
R2745 VTAIL.n265 VTAIL.n223 0.155672
R2746 VTAIL.n257 VTAIL.n223 0.155672
R2747 VTAIL.n257 VTAIL.n256 0.155672
R2748 VTAIL.n256 VTAIL.n227 0.155672
R2749 VTAIL.n249 VTAIL.n227 0.155672
R2750 VTAIL.n249 VTAIL.n248 0.155672
R2751 VTAIL.n248 VTAIL.n232 0.155672
R2752 VTAIL.n241 VTAIL.n232 0.155672
R2753 VTAIL.n241 VTAIL.n240 0.155672
R2754 VTAIL VTAIL.n1 0.0586897
R2755 VN.n55 VN.n29 161.3
R2756 VN.n54 VN.n53 161.3
R2757 VN.n52 VN.n30 161.3
R2758 VN.n51 VN.n50 161.3
R2759 VN.n49 VN.n31 161.3
R2760 VN.n48 VN.n47 161.3
R2761 VN.n46 VN.n45 161.3
R2762 VN.n44 VN.n33 161.3
R2763 VN.n43 VN.n42 161.3
R2764 VN.n41 VN.n34 161.3
R2765 VN.n40 VN.n39 161.3
R2766 VN.n38 VN.n35 161.3
R2767 VN.n26 VN.n0 161.3
R2768 VN.n25 VN.n24 161.3
R2769 VN.n23 VN.n1 161.3
R2770 VN.n22 VN.n21 161.3
R2771 VN.n20 VN.n2 161.3
R2772 VN.n19 VN.n18 161.3
R2773 VN.n17 VN.n16 161.3
R2774 VN.n15 VN.n4 161.3
R2775 VN.n14 VN.n13 161.3
R2776 VN.n12 VN.n5 161.3
R2777 VN.n11 VN.n10 161.3
R2778 VN.n9 VN.n6 161.3
R2779 VN.n7 VN.t3 150.681
R2780 VN.n36 VN.t5 150.681
R2781 VN.n8 VN.t0 116.862
R2782 VN.n3 VN.t7 116.862
R2783 VN.n27 VN.t4 116.862
R2784 VN.n37 VN.t1 116.862
R2785 VN.n32 VN.t6 116.862
R2786 VN.n56 VN.t2 116.862
R2787 VN.n28 VN.n27 99.991
R2788 VN.n57 VN.n56 99.991
R2789 VN.n8 VN.n7 60.757
R2790 VN.n37 VN.n36 60.757
R2791 VN.n14 VN.n5 56.5193
R2792 VN.n21 VN.n1 56.5193
R2793 VN.n43 VN.n34 56.5193
R2794 VN.n50 VN.n30 56.5193
R2795 VN VN.n57 52.0966
R2796 VN.n10 VN.n9 24.4675
R2797 VN.n10 VN.n5 24.4675
R2798 VN.n15 VN.n14 24.4675
R2799 VN.n16 VN.n15 24.4675
R2800 VN.n20 VN.n19 24.4675
R2801 VN.n21 VN.n20 24.4675
R2802 VN.n25 VN.n1 24.4675
R2803 VN.n26 VN.n25 24.4675
R2804 VN.n39 VN.n34 24.4675
R2805 VN.n39 VN.n38 24.4675
R2806 VN.n50 VN.n49 24.4675
R2807 VN.n49 VN.n48 24.4675
R2808 VN.n45 VN.n44 24.4675
R2809 VN.n44 VN.n43 24.4675
R2810 VN.n55 VN.n54 24.4675
R2811 VN.n54 VN.n30 24.4675
R2812 VN.n19 VN.n3 12.7233
R2813 VN.n48 VN.n32 12.7233
R2814 VN.n9 VN.n8 11.7447
R2815 VN.n16 VN.n3 11.7447
R2816 VN.n38 VN.n37 11.7447
R2817 VN.n45 VN.n32 11.7447
R2818 VN.n27 VN.n26 10.766
R2819 VN.n56 VN.n55 10.766
R2820 VN.n36 VN.n35 6.80183
R2821 VN.n7 VN.n6 6.80183
R2822 VN.n57 VN.n29 0.278367
R2823 VN.n28 VN.n0 0.278367
R2824 VN.n53 VN.n29 0.189894
R2825 VN.n53 VN.n52 0.189894
R2826 VN.n52 VN.n51 0.189894
R2827 VN.n51 VN.n31 0.189894
R2828 VN.n47 VN.n31 0.189894
R2829 VN.n47 VN.n46 0.189894
R2830 VN.n46 VN.n33 0.189894
R2831 VN.n42 VN.n33 0.189894
R2832 VN.n42 VN.n41 0.189894
R2833 VN.n41 VN.n40 0.189894
R2834 VN.n40 VN.n35 0.189894
R2835 VN.n11 VN.n6 0.189894
R2836 VN.n12 VN.n11 0.189894
R2837 VN.n13 VN.n12 0.189894
R2838 VN.n13 VN.n4 0.189894
R2839 VN.n17 VN.n4 0.189894
R2840 VN.n18 VN.n17 0.189894
R2841 VN.n18 VN.n2 0.189894
R2842 VN.n22 VN.n2 0.189894
R2843 VN.n23 VN.n22 0.189894
R2844 VN.n24 VN.n23 0.189894
R2845 VN.n24 VN.n0 0.189894
R2846 VN VN.n28 0.153454
R2847 VDD2.n2 VDD2.n1 63.1263
R2848 VDD2.n2 VDD2.n0 63.1263
R2849 VDD2 VDD2.n5 63.1233
R2850 VDD2.n4 VDD2.n3 61.8972
R2851 VDD2.n4 VDD2.n2 46.3532
R2852 VDD2.n5 VDD2.t6 1.54136
R2853 VDD2.n5 VDD2.t2 1.54136
R2854 VDD2.n3 VDD2.t5 1.54136
R2855 VDD2.n3 VDD2.t1 1.54136
R2856 VDD2.n1 VDD2.t0 1.54136
R2857 VDD2.n1 VDD2.t3 1.54136
R2858 VDD2.n0 VDD2.t4 1.54136
R2859 VDD2.n0 VDD2.t7 1.54136
R2860 VDD2 VDD2.n4 1.34317
C0 VN VTAIL 9.68213f
C1 VDD2 VN 9.307099f
C2 VDD2 VTAIL 8.425961f
C3 VDD1 VN 0.151926f
C4 VDD1 VTAIL 8.371201f
C5 VDD1 VDD2 1.80416f
C6 VN VP 7.87862f
C7 VTAIL VP 9.69624f
C8 VDD2 VP 0.525099f
C9 VDD1 VP 9.67885f
C10 VDD2 B 5.46155f
C11 VDD1 B 5.907126f
C12 VTAIL B 11.034698f
C13 VN B 15.754689f
C14 VP B 14.334085f
C15 VDD2.t4 B 0.246005f
C16 VDD2.t7 B 0.246005f
C17 VDD2.n0 B 2.21072f
C18 VDD2.t0 B 0.246005f
C19 VDD2.t3 B 0.246005f
C20 VDD2.n1 B 2.21072f
C21 VDD2.n2 B 3.2602f
C22 VDD2.t5 B 0.246005f
C23 VDD2.t1 B 0.246005f
C24 VDD2.n3 B 2.20082f
C25 VDD2.n4 B 2.94053f
C26 VDD2.t6 B 0.246005f
C27 VDD2.t2 B 0.246005f
C28 VDD2.n5 B 2.21067f
C29 VN.n0 B 0.028636f
C30 VN.t4 B 2.01903f
C31 VN.n1 B 0.032918f
C32 VN.n2 B 0.02172f
C33 VN.t7 B 2.01903f
C34 VN.n3 B 0.710919f
C35 VN.n4 B 0.02172f
C36 VN.n5 B 0.031708f
C37 VN.n6 B 0.211038f
C38 VN.t0 B 2.01903f
C39 VN.t3 B 2.20935f
C40 VN.n7 B 0.750337f
C41 VN.n8 B 0.773832f
C42 VN.n9 B 0.030089f
C43 VN.n10 B 0.040481f
C44 VN.n11 B 0.02172f
C45 VN.n12 B 0.02172f
C46 VN.n13 B 0.02172f
C47 VN.n14 B 0.031708f
C48 VN.n15 B 0.040481f
C49 VN.n16 B 0.030089f
C50 VN.n17 B 0.02172f
C51 VN.n18 B 0.02172f
C52 VN.n19 B 0.030888f
C53 VN.n20 B 0.040481f
C54 VN.n21 B 0.030497f
C55 VN.n22 B 0.02172f
C56 VN.n23 B 0.02172f
C57 VN.n24 B 0.02172f
C58 VN.n25 B 0.040481f
C59 VN.n26 B 0.029289f
C60 VN.n27 B 0.786269f
C61 VN.n28 B 0.035218f
C62 VN.n29 B 0.028636f
C63 VN.t2 B 2.01903f
C64 VN.n30 B 0.032918f
C65 VN.n31 B 0.02172f
C66 VN.t6 B 2.01903f
C67 VN.n32 B 0.710919f
C68 VN.n33 B 0.02172f
C69 VN.n34 B 0.031708f
C70 VN.n35 B 0.211038f
C71 VN.t1 B 2.01903f
C72 VN.t5 B 2.20935f
C73 VN.n36 B 0.750337f
C74 VN.n37 B 0.773832f
C75 VN.n38 B 0.030089f
C76 VN.n39 B 0.040481f
C77 VN.n40 B 0.02172f
C78 VN.n41 B 0.02172f
C79 VN.n42 B 0.02172f
C80 VN.n43 B 0.031708f
C81 VN.n44 B 0.040481f
C82 VN.n45 B 0.030089f
C83 VN.n46 B 0.02172f
C84 VN.n47 B 0.02172f
C85 VN.n48 B 0.030888f
C86 VN.n49 B 0.040481f
C87 VN.n50 B 0.030497f
C88 VN.n51 B 0.02172f
C89 VN.n52 B 0.02172f
C90 VN.n53 B 0.02172f
C91 VN.n54 B 0.040481f
C92 VN.n55 B 0.029289f
C93 VN.n56 B 0.786269f
C94 VN.n57 B 1.28502f
C95 VTAIL.t4 B 0.199216f
C96 VTAIL.t0 B 0.199216f
C97 VTAIL.n0 B 1.72339f
C98 VTAIL.n1 B 0.361508f
C99 VTAIL.n2 B 0.028237f
C100 VTAIL.n3 B 0.019619f
C101 VTAIL.n4 B 0.010542f
C102 VTAIL.n5 B 0.024918f
C103 VTAIL.n6 B 0.011162f
C104 VTAIL.n7 B 0.019619f
C105 VTAIL.n8 B 0.010542f
C106 VTAIL.n9 B 0.024918f
C107 VTAIL.n10 B 0.011162f
C108 VTAIL.n11 B 0.019619f
C109 VTAIL.n12 B 0.010542f
C110 VTAIL.n13 B 0.024918f
C111 VTAIL.n14 B 0.011162f
C112 VTAIL.n15 B 0.019619f
C113 VTAIL.n16 B 0.010542f
C114 VTAIL.n17 B 0.024918f
C115 VTAIL.n18 B 0.011162f
C116 VTAIL.n19 B 0.019619f
C117 VTAIL.n20 B 0.010542f
C118 VTAIL.n21 B 0.024918f
C119 VTAIL.n22 B 0.011162f
C120 VTAIL.n23 B 0.14785f
C121 VTAIL.t6 B 0.042174f
C122 VTAIL.n24 B 0.018688f
C123 VTAIL.n25 B 0.017615f
C124 VTAIL.n26 B 0.010542f
C125 VTAIL.n27 B 1.0639f
C126 VTAIL.n28 B 0.019619f
C127 VTAIL.n29 B 0.010542f
C128 VTAIL.n30 B 0.011162f
C129 VTAIL.n31 B 0.024918f
C130 VTAIL.n32 B 0.024918f
C131 VTAIL.n33 B 0.011162f
C132 VTAIL.n34 B 0.010542f
C133 VTAIL.n35 B 0.019619f
C134 VTAIL.n36 B 0.019619f
C135 VTAIL.n37 B 0.010542f
C136 VTAIL.n38 B 0.011162f
C137 VTAIL.n39 B 0.024918f
C138 VTAIL.n40 B 0.024918f
C139 VTAIL.n41 B 0.024918f
C140 VTAIL.n42 B 0.011162f
C141 VTAIL.n43 B 0.010542f
C142 VTAIL.n44 B 0.019619f
C143 VTAIL.n45 B 0.019619f
C144 VTAIL.n46 B 0.010542f
C145 VTAIL.n47 B 0.010852f
C146 VTAIL.n48 B 0.010852f
C147 VTAIL.n49 B 0.024918f
C148 VTAIL.n50 B 0.024918f
C149 VTAIL.n51 B 0.011162f
C150 VTAIL.n52 B 0.010542f
C151 VTAIL.n53 B 0.019619f
C152 VTAIL.n54 B 0.019619f
C153 VTAIL.n55 B 0.010542f
C154 VTAIL.n56 B 0.011162f
C155 VTAIL.n57 B 0.024918f
C156 VTAIL.n58 B 0.024918f
C157 VTAIL.n59 B 0.011162f
C158 VTAIL.n60 B 0.010542f
C159 VTAIL.n61 B 0.019619f
C160 VTAIL.n62 B 0.019619f
C161 VTAIL.n63 B 0.010542f
C162 VTAIL.n64 B 0.011162f
C163 VTAIL.n65 B 0.024918f
C164 VTAIL.n66 B 0.055113f
C165 VTAIL.n67 B 0.011162f
C166 VTAIL.n68 B 0.010542f
C167 VTAIL.n69 B 0.045615f
C168 VTAIL.n70 B 0.030967f
C169 VTAIL.n71 B 0.209006f
C170 VTAIL.n72 B 0.028237f
C171 VTAIL.n73 B 0.019619f
C172 VTAIL.n74 B 0.010542f
C173 VTAIL.n75 B 0.024918f
C174 VTAIL.n76 B 0.011162f
C175 VTAIL.n77 B 0.019619f
C176 VTAIL.n78 B 0.010542f
C177 VTAIL.n79 B 0.024918f
C178 VTAIL.n80 B 0.011162f
C179 VTAIL.n81 B 0.019619f
C180 VTAIL.n82 B 0.010542f
C181 VTAIL.n83 B 0.024918f
C182 VTAIL.n84 B 0.011162f
C183 VTAIL.n85 B 0.019619f
C184 VTAIL.n86 B 0.010542f
C185 VTAIL.n87 B 0.024918f
C186 VTAIL.n88 B 0.011162f
C187 VTAIL.n89 B 0.019619f
C188 VTAIL.n90 B 0.010542f
C189 VTAIL.n91 B 0.024918f
C190 VTAIL.n92 B 0.011162f
C191 VTAIL.n93 B 0.14785f
C192 VTAIL.t14 B 0.042174f
C193 VTAIL.n94 B 0.018688f
C194 VTAIL.n95 B 0.017615f
C195 VTAIL.n96 B 0.010542f
C196 VTAIL.n97 B 1.0639f
C197 VTAIL.n98 B 0.019619f
C198 VTAIL.n99 B 0.010542f
C199 VTAIL.n100 B 0.011162f
C200 VTAIL.n101 B 0.024918f
C201 VTAIL.n102 B 0.024918f
C202 VTAIL.n103 B 0.011162f
C203 VTAIL.n104 B 0.010542f
C204 VTAIL.n105 B 0.019619f
C205 VTAIL.n106 B 0.019619f
C206 VTAIL.n107 B 0.010542f
C207 VTAIL.n108 B 0.011162f
C208 VTAIL.n109 B 0.024918f
C209 VTAIL.n110 B 0.024918f
C210 VTAIL.n111 B 0.024918f
C211 VTAIL.n112 B 0.011162f
C212 VTAIL.n113 B 0.010542f
C213 VTAIL.n114 B 0.019619f
C214 VTAIL.n115 B 0.019619f
C215 VTAIL.n116 B 0.010542f
C216 VTAIL.n117 B 0.010852f
C217 VTAIL.n118 B 0.010852f
C218 VTAIL.n119 B 0.024918f
C219 VTAIL.n120 B 0.024918f
C220 VTAIL.n121 B 0.011162f
C221 VTAIL.n122 B 0.010542f
C222 VTAIL.n123 B 0.019619f
C223 VTAIL.n124 B 0.019619f
C224 VTAIL.n125 B 0.010542f
C225 VTAIL.n126 B 0.011162f
C226 VTAIL.n127 B 0.024918f
C227 VTAIL.n128 B 0.024918f
C228 VTAIL.n129 B 0.011162f
C229 VTAIL.n130 B 0.010542f
C230 VTAIL.n131 B 0.019619f
C231 VTAIL.n132 B 0.019619f
C232 VTAIL.n133 B 0.010542f
C233 VTAIL.n134 B 0.011162f
C234 VTAIL.n135 B 0.024918f
C235 VTAIL.n136 B 0.055113f
C236 VTAIL.n137 B 0.011162f
C237 VTAIL.n138 B 0.010542f
C238 VTAIL.n139 B 0.045615f
C239 VTAIL.n140 B 0.030967f
C240 VTAIL.n141 B 0.209006f
C241 VTAIL.t9 B 0.199216f
C242 VTAIL.t15 B 0.199216f
C243 VTAIL.n142 B 1.72339f
C244 VTAIL.n143 B 0.520228f
C245 VTAIL.n144 B 0.028237f
C246 VTAIL.n145 B 0.019619f
C247 VTAIL.n146 B 0.010542f
C248 VTAIL.n147 B 0.024918f
C249 VTAIL.n148 B 0.011162f
C250 VTAIL.n149 B 0.019619f
C251 VTAIL.n150 B 0.010542f
C252 VTAIL.n151 B 0.024918f
C253 VTAIL.n152 B 0.011162f
C254 VTAIL.n153 B 0.019619f
C255 VTAIL.n154 B 0.010542f
C256 VTAIL.n155 B 0.024918f
C257 VTAIL.n156 B 0.011162f
C258 VTAIL.n157 B 0.019619f
C259 VTAIL.n158 B 0.010542f
C260 VTAIL.n159 B 0.024918f
C261 VTAIL.n160 B 0.011162f
C262 VTAIL.n161 B 0.019619f
C263 VTAIL.n162 B 0.010542f
C264 VTAIL.n163 B 0.024918f
C265 VTAIL.n164 B 0.011162f
C266 VTAIL.n165 B 0.14785f
C267 VTAIL.t13 B 0.042174f
C268 VTAIL.n166 B 0.018688f
C269 VTAIL.n167 B 0.017615f
C270 VTAIL.n168 B 0.010542f
C271 VTAIL.n169 B 1.0639f
C272 VTAIL.n170 B 0.019619f
C273 VTAIL.n171 B 0.010542f
C274 VTAIL.n172 B 0.011162f
C275 VTAIL.n173 B 0.024918f
C276 VTAIL.n174 B 0.024918f
C277 VTAIL.n175 B 0.011162f
C278 VTAIL.n176 B 0.010542f
C279 VTAIL.n177 B 0.019619f
C280 VTAIL.n178 B 0.019619f
C281 VTAIL.n179 B 0.010542f
C282 VTAIL.n180 B 0.011162f
C283 VTAIL.n181 B 0.024918f
C284 VTAIL.n182 B 0.024918f
C285 VTAIL.n183 B 0.024918f
C286 VTAIL.n184 B 0.011162f
C287 VTAIL.n185 B 0.010542f
C288 VTAIL.n186 B 0.019619f
C289 VTAIL.n187 B 0.019619f
C290 VTAIL.n188 B 0.010542f
C291 VTAIL.n189 B 0.010852f
C292 VTAIL.n190 B 0.010852f
C293 VTAIL.n191 B 0.024918f
C294 VTAIL.n192 B 0.024918f
C295 VTAIL.n193 B 0.011162f
C296 VTAIL.n194 B 0.010542f
C297 VTAIL.n195 B 0.019619f
C298 VTAIL.n196 B 0.019619f
C299 VTAIL.n197 B 0.010542f
C300 VTAIL.n198 B 0.011162f
C301 VTAIL.n199 B 0.024918f
C302 VTAIL.n200 B 0.024918f
C303 VTAIL.n201 B 0.011162f
C304 VTAIL.n202 B 0.010542f
C305 VTAIL.n203 B 0.019619f
C306 VTAIL.n204 B 0.019619f
C307 VTAIL.n205 B 0.010542f
C308 VTAIL.n206 B 0.011162f
C309 VTAIL.n207 B 0.024918f
C310 VTAIL.n208 B 0.055113f
C311 VTAIL.n209 B 0.011162f
C312 VTAIL.n210 B 0.010542f
C313 VTAIL.n211 B 0.045615f
C314 VTAIL.n212 B 0.030967f
C315 VTAIL.n213 B 1.30847f
C316 VTAIL.n214 B 0.028237f
C317 VTAIL.n215 B 0.019619f
C318 VTAIL.n216 B 0.010542f
C319 VTAIL.n217 B 0.024918f
C320 VTAIL.n218 B 0.011162f
C321 VTAIL.n219 B 0.019619f
C322 VTAIL.n220 B 0.010542f
C323 VTAIL.n221 B 0.024918f
C324 VTAIL.n222 B 0.011162f
C325 VTAIL.n223 B 0.019619f
C326 VTAIL.n224 B 0.010542f
C327 VTAIL.n225 B 0.024918f
C328 VTAIL.n226 B 0.011162f
C329 VTAIL.n227 B 0.019619f
C330 VTAIL.n228 B 0.010542f
C331 VTAIL.n229 B 0.024918f
C332 VTAIL.n230 B 0.024918f
C333 VTAIL.n231 B 0.011162f
C334 VTAIL.n232 B 0.019619f
C335 VTAIL.n233 B 0.010542f
C336 VTAIL.n234 B 0.024918f
C337 VTAIL.n235 B 0.011162f
C338 VTAIL.n236 B 0.14785f
C339 VTAIL.t5 B 0.042174f
C340 VTAIL.n237 B 0.018688f
C341 VTAIL.n238 B 0.017615f
C342 VTAIL.n239 B 0.010542f
C343 VTAIL.n240 B 1.0639f
C344 VTAIL.n241 B 0.019619f
C345 VTAIL.n242 B 0.010542f
C346 VTAIL.n243 B 0.011162f
C347 VTAIL.n244 B 0.024918f
C348 VTAIL.n245 B 0.024918f
C349 VTAIL.n246 B 0.011162f
C350 VTAIL.n247 B 0.010542f
C351 VTAIL.n248 B 0.019619f
C352 VTAIL.n249 B 0.019619f
C353 VTAIL.n250 B 0.010542f
C354 VTAIL.n251 B 0.011162f
C355 VTAIL.n252 B 0.024918f
C356 VTAIL.n253 B 0.024918f
C357 VTAIL.n254 B 0.011162f
C358 VTAIL.n255 B 0.010542f
C359 VTAIL.n256 B 0.019619f
C360 VTAIL.n257 B 0.019619f
C361 VTAIL.n258 B 0.010542f
C362 VTAIL.n259 B 0.010852f
C363 VTAIL.n260 B 0.010852f
C364 VTAIL.n261 B 0.024918f
C365 VTAIL.n262 B 0.024918f
C366 VTAIL.n263 B 0.011162f
C367 VTAIL.n264 B 0.010542f
C368 VTAIL.n265 B 0.019619f
C369 VTAIL.n266 B 0.019619f
C370 VTAIL.n267 B 0.010542f
C371 VTAIL.n268 B 0.011162f
C372 VTAIL.n269 B 0.024918f
C373 VTAIL.n270 B 0.024918f
C374 VTAIL.n271 B 0.011162f
C375 VTAIL.n272 B 0.010542f
C376 VTAIL.n273 B 0.019619f
C377 VTAIL.n274 B 0.019619f
C378 VTAIL.n275 B 0.010542f
C379 VTAIL.n276 B 0.011162f
C380 VTAIL.n277 B 0.024918f
C381 VTAIL.n278 B 0.055113f
C382 VTAIL.n279 B 0.011162f
C383 VTAIL.n280 B 0.010542f
C384 VTAIL.n281 B 0.045615f
C385 VTAIL.n282 B 0.030967f
C386 VTAIL.n283 B 1.30847f
C387 VTAIL.t3 B 0.199216f
C388 VTAIL.t2 B 0.199216f
C389 VTAIL.n284 B 1.7234f
C390 VTAIL.n285 B 0.520226f
C391 VTAIL.n286 B 0.028237f
C392 VTAIL.n287 B 0.019619f
C393 VTAIL.n288 B 0.010542f
C394 VTAIL.n289 B 0.024918f
C395 VTAIL.n290 B 0.011162f
C396 VTAIL.n291 B 0.019619f
C397 VTAIL.n292 B 0.010542f
C398 VTAIL.n293 B 0.024918f
C399 VTAIL.n294 B 0.011162f
C400 VTAIL.n295 B 0.019619f
C401 VTAIL.n296 B 0.010542f
C402 VTAIL.n297 B 0.024918f
C403 VTAIL.n298 B 0.011162f
C404 VTAIL.n299 B 0.019619f
C405 VTAIL.n300 B 0.010542f
C406 VTAIL.n301 B 0.024918f
C407 VTAIL.n302 B 0.024918f
C408 VTAIL.n303 B 0.011162f
C409 VTAIL.n304 B 0.019619f
C410 VTAIL.n305 B 0.010542f
C411 VTAIL.n306 B 0.024918f
C412 VTAIL.n307 B 0.011162f
C413 VTAIL.n308 B 0.14785f
C414 VTAIL.t7 B 0.042174f
C415 VTAIL.n309 B 0.018688f
C416 VTAIL.n310 B 0.017615f
C417 VTAIL.n311 B 0.010542f
C418 VTAIL.n312 B 1.0639f
C419 VTAIL.n313 B 0.019619f
C420 VTAIL.n314 B 0.010542f
C421 VTAIL.n315 B 0.011162f
C422 VTAIL.n316 B 0.024918f
C423 VTAIL.n317 B 0.024918f
C424 VTAIL.n318 B 0.011162f
C425 VTAIL.n319 B 0.010542f
C426 VTAIL.n320 B 0.019619f
C427 VTAIL.n321 B 0.019619f
C428 VTAIL.n322 B 0.010542f
C429 VTAIL.n323 B 0.011162f
C430 VTAIL.n324 B 0.024918f
C431 VTAIL.n325 B 0.024918f
C432 VTAIL.n326 B 0.011162f
C433 VTAIL.n327 B 0.010542f
C434 VTAIL.n328 B 0.019619f
C435 VTAIL.n329 B 0.019619f
C436 VTAIL.n330 B 0.010542f
C437 VTAIL.n331 B 0.010852f
C438 VTAIL.n332 B 0.010852f
C439 VTAIL.n333 B 0.024918f
C440 VTAIL.n334 B 0.024918f
C441 VTAIL.n335 B 0.011162f
C442 VTAIL.n336 B 0.010542f
C443 VTAIL.n337 B 0.019619f
C444 VTAIL.n338 B 0.019619f
C445 VTAIL.n339 B 0.010542f
C446 VTAIL.n340 B 0.011162f
C447 VTAIL.n341 B 0.024918f
C448 VTAIL.n342 B 0.024918f
C449 VTAIL.n343 B 0.011162f
C450 VTAIL.n344 B 0.010542f
C451 VTAIL.n345 B 0.019619f
C452 VTAIL.n346 B 0.019619f
C453 VTAIL.n347 B 0.010542f
C454 VTAIL.n348 B 0.011162f
C455 VTAIL.n349 B 0.024918f
C456 VTAIL.n350 B 0.055113f
C457 VTAIL.n351 B 0.011162f
C458 VTAIL.n352 B 0.010542f
C459 VTAIL.n353 B 0.045615f
C460 VTAIL.n354 B 0.030967f
C461 VTAIL.n355 B 0.209006f
C462 VTAIL.n356 B 0.028237f
C463 VTAIL.n357 B 0.019619f
C464 VTAIL.n358 B 0.010542f
C465 VTAIL.n359 B 0.024918f
C466 VTAIL.n360 B 0.011162f
C467 VTAIL.n361 B 0.019619f
C468 VTAIL.n362 B 0.010542f
C469 VTAIL.n363 B 0.024918f
C470 VTAIL.n364 B 0.011162f
C471 VTAIL.n365 B 0.019619f
C472 VTAIL.n366 B 0.010542f
C473 VTAIL.n367 B 0.024918f
C474 VTAIL.n368 B 0.011162f
C475 VTAIL.n369 B 0.019619f
C476 VTAIL.n370 B 0.010542f
C477 VTAIL.n371 B 0.024918f
C478 VTAIL.n372 B 0.024918f
C479 VTAIL.n373 B 0.011162f
C480 VTAIL.n374 B 0.019619f
C481 VTAIL.n375 B 0.010542f
C482 VTAIL.n376 B 0.024918f
C483 VTAIL.n377 B 0.011162f
C484 VTAIL.n378 B 0.14785f
C485 VTAIL.t11 B 0.042174f
C486 VTAIL.n379 B 0.018688f
C487 VTAIL.n380 B 0.017615f
C488 VTAIL.n381 B 0.010542f
C489 VTAIL.n382 B 1.0639f
C490 VTAIL.n383 B 0.019619f
C491 VTAIL.n384 B 0.010542f
C492 VTAIL.n385 B 0.011162f
C493 VTAIL.n386 B 0.024918f
C494 VTAIL.n387 B 0.024918f
C495 VTAIL.n388 B 0.011162f
C496 VTAIL.n389 B 0.010542f
C497 VTAIL.n390 B 0.019619f
C498 VTAIL.n391 B 0.019619f
C499 VTAIL.n392 B 0.010542f
C500 VTAIL.n393 B 0.011162f
C501 VTAIL.n394 B 0.024918f
C502 VTAIL.n395 B 0.024918f
C503 VTAIL.n396 B 0.011162f
C504 VTAIL.n397 B 0.010542f
C505 VTAIL.n398 B 0.019619f
C506 VTAIL.n399 B 0.019619f
C507 VTAIL.n400 B 0.010542f
C508 VTAIL.n401 B 0.010852f
C509 VTAIL.n402 B 0.010852f
C510 VTAIL.n403 B 0.024918f
C511 VTAIL.n404 B 0.024918f
C512 VTAIL.n405 B 0.011162f
C513 VTAIL.n406 B 0.010542f
C514 VTAIL.n407 B 0.019619f
C515 VTAIL.n408 B 0.019619f
C516 VTAIL.n409 B 0.010542f
C517 VTAIL.n410 B 0.011162f
C518 VTAIL.n411 B 0.024918f
C519 VTAIL.n412 B 0.024918f
C520 VTAIL.n413 B 0.011162f
C521 VTAIL.n414 B 0.010542f
C522 VTAIL.n415 B 0.019619f
C523 VTAIL.n416 B 0.019619f
C524 VTAIL.n417 B 0.010542f
C525 VTAIL.n418 B 0.011162f
C526 VTAIL.n419 B 0.024918f
C527 VTAIL.n420 B 0.055113f
C528 VTAIL.n421 B 0.011162f
C529 VTAIL.n422 B 0.010542f
C530 VTAIL.n423 B 0.045615f
C531 VTAIL.n424 B 0.030967f
C532 VTAIL.n425 B 0.209006f
C533 VTAIL.t8 B 0.199216f
C534 VTAIL.t12 B 0.199216f
C535 VTAIL.n426 B 1.7234f
C536 VTAIL.n427 B 0.520226f
C537 VTAIL.n428 B 0.028237f
C538 VTAIL.n429 B 0.019619f
C539 VTAIL.n430 B 0.010542f
C540 VTAIL.n431 B 0.024918f
C541 VTAIL.n432 B 0.011162f
C542 VTAIL.n433 B 0.019619f
C543 VTAIL.n434 B 0.010542f
C544 VTAIL.n435 B 0.024918f
C545 VTAIL.n436 B 0.011162f
C546 VTAIL.n437 B 0.019619f
C547 VTAIL.n438 B 0.010542f
C548 VTAIL.n439 B 0.024918f
C549 VTAIL.n440 B 0.011162f
C550 VTAIL.n441 B 0.019619f
C551 VTAIL.n442 B 0.010542f
C552 VTAIL.n443 B 0.024918f
C553 VTAIL.n444 B 0.024918f
C554 VTAIL.n445 B 0.011162f
C555 VTAIL.n446 B 0.019619f
C556 VTAIL.n447 B 0.010542f
C557 VTAIL.n448 B 0.024918f
C558 VTAIL.n449 B 0.011162f
C559 VTAIL.n450 B 0.14785f
C560 VTAIL.t10 B 0.042174f
C561 VTAIL.n451 B 0.018688f
C562 VTAIL.n452 B 0.017615f
C563 VTAIL.n453 B 0.010542f
C564 VTAIL.n454 B 1.0639f
C565 VTAIL.n455 B 0.019619f
C566 VTAIL.n456 B 0.010542f
C567 VTAIL.n457 B 0.011162f
C568 VTAIL.n458 B 0.024918f
C569 VTAIL.n459 B 0.024918f
C570 VTAIL.n460 B 0.011162f
C571 VTAIL.n461 B 0.010542f
C572 VTAIL.n462 B 0.019619f
C573 VTAIL.n463 B 0.019619f
C574 VTAIL.n464 B 0.010542f
C575 VTAIL.n465 B 0.011162f
C576 VTAIL.n466 B 0.024918f
C577 VTAIL.n467 B 0.024918f
C578 VTAIL.n468 B 0.011162f
C579 VTAIL.n469 B 0.010542f
C580 VTAIL.n470 B 0.019619f
C581 VTAIL.n471 B 0.019619f
C582 VTAIL.n472 B 0.010542f
C583 VTAIL.n473 B 0.010852f
C584 VTAIL.n474 B 0.010852f
C585 VTAIL.n475 B 0.024918f
C586 VTAIL.n476 B 0.024918f
C587 VTAIL.n477 B 0.011162f
C588 VTAIL.n478 B 0.010542f
C589 VTAIL.n479 B 0.019619f
C590 VTAIL.n480 B 0.019619f
C591 VTAIL.n481 B 0.010542f
C592 VTAIL.n482 B 0.011162f
C593 VTAIL.n483 B 0.024918f
C594 VTAIL.n484 B 0.024918f
C595 VTAIL.n485 B 0.011162f
C596 VTAIL.n486 B 0.010542f
C597 VTAIL.n487 B 0.019619f
C598 VTAIL.n488 B 0.019619f
C599 VTAIL.n489 B 0.010542f
C600 VTAIL.n490 B 0.011162f
C601 VTAIL.n491 B 0.024918f
C602 VTAIL.n492 B 0.055113f
C603 VTAIL.n493 B 0.011162f
C604 VTAIL.n494 B 0.010542f
C605 VTAIL.n495 B 0.045615f
C606 VTAIL.n496 B 0.030967f
C607 VTAIL.n497 B 1.30847f
C608 VTAIL.n498 B 0.028237f
C609 VTAIL.n499 B 0.019619f
C610 VTAIL.n500 B 0.010542f
C611 VTAIL.n501 B 0.024918f
C612 VTAIL.n502 B 0.011162f
C613 VTAIL.n503 B 0.019619f
C614 VTAIL.n504 B 0.010542f
C615 VTAIL.n505 B 0.024918f
C616 VTAIL.n506 B 0.011162f
C617 VTAIL.n507 B 0.019619f
C618 VTAIL.n508 B 0.010542f
C619 VTAIL.n509 B 0.024918f
C620 VTAIL.n510 B 0.011162f
C621 VTAIL.n511 B 0.019619f
C622 VTAIL.n512 B 0.010542f
C623 VTAIL.n513 B 0.024918f
C624 VTAIL.n514 B 0.011162f
C625 VTAIL.n515 B 0.019619f
C626 VTAIL.n516 B 0.010542f
C627 VTAIL.n517 B 0.024918f
C628 VTAIL.n518 B 0.011162f
C629 VTAIL.n519 B 0.14785f
C630 VTAIL.t1 B 0.042174f
C631 VTAIL.n520 B 0.018688f
C632 VTAIL.n521 B 0.017615f
C633 VTAIL.n522 B 0.010542f
C634 VTAIL.n523 B 1.0639f
C635 VTAIL.n524 B 0.019619f
C636 VTAIL.n525 B 0.010542f
C637 VTAIL.n526 B 0.011162f
C638 VTAIL.n527 B 0.024918f
C639 VTAIL.n528 B 0.024918f
C640 VTAIL.n529 B 0.011162f
C641 VTAIL.n530 B 0.010542f
C642 VTAIL.n531 B 0.019619f
C643 VTAIL.n532 B 0.019619f
C644 VTAIL.n533 B 0.010542f
C645 VTAIL.n534 B 0.011162f
C646 VTAIL.n535 B 0.024918f
C647 VTAIL.n536 B 0.024918f
C648 VTAIL.n537 B 0.024918f
C649 VTAIL.n538 B 0.011162f
C650 VTAIL.n539 B 0.010542f
C651 VTAIL.n540 B 0.019619f
C652 VTAIL.n541 B 0.019619f
C653 VTAIL.n542 B 0.010542f
C654 VTAIL.n543 B 0.010852f
C655 VTAIL.n544 B 0.010852f
C656 VTAIL.n545 B 0.024918f
C657 VTAIL.n546 B 0.024918f
C658 VTAIL.n547 B 0.011162f
C659 VTAIL.n548 B 0.010542f
C660 VTAIL.n549 B 0.019619f
C661 VTAIL.n550 B 0.019619f
C662 VTAIL.n551 B 0.010542f
C663 VTAIL.n552 B 0.011162f
C664 VTAIL.n553 B 0.024918f
C665 VTAIL.n554 B 0.024918f
C666 VTAIL.n555 B 0.011162f
C667 VTAIL.n556 B 0.010542f
C668 VTAIL.n557 B 0.019619f
C669 VTAIL.n558 B 0.019619f
C670 VTAIL.n559 B 0.010542f
C671 VTAIL.n560 B 0.011162f
C672 VTAIL.n561 B 0.024918f
C673 VTAIL.n562 B 0.055113f
C674 VTAIL.n563 B 0.011162f
C675 VTAIL.n564 B 0.010542f
C676 VTAIL.n565 B 0.045615f
C677 VTAIL.n566 B 0.030967f
C678 VTAIL.n567 B 1.30479f
C679 VDD1.t7 B 0.250299f
C680 VDD1.t2 B 0.250299f
C681 VDD1.n0 B 2.2504f
C682 VDD1.t1 B 0.250299f
C683 VDD1.t5 B 0.250299f
C684 VDD1.n1 B 2.2493f
C685 VDD1.t3 B 0.250299f
C686 VDD1.t4 B 0.250299f
C687 VDD1.n2 B 2.2493f
C688 VDD1.n3 B 3.36839f
C689 VDD1.t0 B 0.250299f
C690 VDD1.t6 B 0.250299f
C691 VDD1.n4 B 2.23923f
C692 VDD1.n5 B 3.02238f
C693 VP.n0 B 0.029095f
C694 VP.t1 B 2.05138f
C695 VP.n1 B 0.033446f
C696 VP.n2 B 0.022068f
C697 VP.t0 B 2.05138f
C698 VP.n3 B 0.72231f
C699 VP.n4 B 0.022068f
C700 VP.n5 B 0.032216f
C701 VP.n6 B 0.022068f
C702 VP.t6 B 2.05138f
C703 VP.n7 B 0.04113f
C704 VP.n8 B 0.022068f
C705 VP.n9 B 0.029759f
C706 VP.n10 B 0.029095f
C707 VP.t5 B 2.05138f
C708 VP.n11 B 0.033446f
C709 VP.n12 B 0.022068f
C710 VP.t3 B 2.05138f
C711 VP.n13 B 0.72231f
C712 VP.n14 B 0.022068f
C713 VP.n15 B 0.032216f
C714 VP.n16 B 0.214419f
C715 VP.t7 B 2.05138f
C716 VP.t4 B 2.24475f
C717 VP.n17 B 0.762359f
C718 VP.n18 B 0.786232f
C719 VP.n19 B 0.030571f
C720 VP.n20 B 0.04113f
C721 VP.n21 B 0.022068f
C722 VP.n22 B 0.022068f
C723 VP.n23 B 0.022068f
C724 VP.n24 B 0.032216f
C725 VP.n25 B 0.04113f
C726 VP.n26 B 0.030571f
C727 VP.n27 B 0.022068f
C728 VP.n28 B 0.022068f
C729 VP.n29 B 0.031383f
C730 VP.n30 B 0.04113f
C731 VP.n31 B 0.030986f
C732 VP.n32 B 0.022068f
C733 VP.n33 B 0.022068f
C734 VP.n34 B 0.022068f
C735 VP.n35 B 0.04113f
C736 VP.n36 B 0.029759f
C737 VP.n37 B 0.798867f
C738 VP.n38 B 1.29382f
C739 VP.t2 B 2.05138f
C740 VP.n39 B 0.798867f
C741 VP.n40 B 1.30913f
C742 VP.n41 B 0.029095f
C743 VP.n42 B 0.022068f
C744 VP.n43 B 0.04113f
C745 VP.n44 B 0.033446f
C746 VP.n45 B 0.030986f
C747 VP.n46 B 0.022068f
C748 VP.n47 B 0.022068f
C749 VP.n48 B 0.022068f
C750 VP.n49 B 0.031383f
C751 VP.n50 B 0.72231f
C752 VP.n51 B 0.030571f
C753 VP.n52 B 0.04113f
C754 VP.n53 B 0.022068f
C755 VP.n54 B 0.022068f
C756 VP.n55 B 0.022068f
C757 VP.n56 B 0.032216f
C758 VP.n57 B 0.04113f
C759 VP.n58 B 0.030571f
C760 VP.n59 B 0.022068f
C761 VP.n60 B 0.022068f
C762 VP.n61 B 0.031383f
C763 VP.n62 B 0.04113f
C764 VP.n63 B 0.030986f
C765 VP.n64 B 0.022068f
C766 VP.n65 B 0.022068f
C767 VP.n66 B 0.022068f
C768 VP.n67 B 0.04113f
C769 VP.n68 B 0.029759f
C770 VP.n69 B 0.798867f
C771 VP.n70 B 0.035782f
.ends

