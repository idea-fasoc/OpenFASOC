* NGSPICE file created from diff_pair_sample_0032.ext - technology: sky130A

.subckt diff_pair_sample_0032 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0.32505 ps=2.3 w=1.97 l=1.72
X1 VDD2.t7 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.7683 ps=4.72 w=1.97 l=1.72
X2 VTAIL.t7 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0.32505 ps=2.3 w=1.97 l=1.72
X3 VDD1.t6 VP.t1 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.7683 ps=4.72 w=1.97 l=1.72
X4 VTAIL.t1 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X5 VTAIL.t13 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0.32505 ps=2.3 w=1.97 l=1.72
X6 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=1.72
X7 VDD1.t3 VP.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X8 VTAIL.t3 VN.t3 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0.32505 ps=2.3 w=1.97 l=1.72
X9 VTAIL.t0 VN.t4 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X10 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=1.72
X11 VTAIL.t11 VP.t4 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X12 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=1.72
X13 VTAIL.t10 VP.t5 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X14 VDD2.t2 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.7683 ps=4.72 w=1.97 l=1.72
X15 VDD2.t1 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X16 VDD2.t0 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X17 VDD1.t1 VP.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.32505 ps=2.3 w=1.97 l=1.72
X18 VDD1.t7 VP.t7 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.32505 pd=2.3 as=0.7683 ps=4.72 w=1.97 l=1.72
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7683 pd=4.72 as=0 ps=0 w=1.97 l=1.72
R0 VP.n31 VP.n30 182.097
R1 VP.n54 VP.n53 182.097
R2 VP.n29 VP.n28 182.097
R3 VP.n14 VP.n11 161.3
R4 VP.n16 VP.n15 161.3
R5 VP.n17 VP.n10 161.3
R6 VP.n19 VP.n18 161.3
R7 VP.n20 VP.n9 161.3
R8 VP.n23 VP.n22 161.3
R9 VP.n24 VP.n8 161.3
R10 VP.n26 VP.n25 161.3
R11 VP.n27 VP.n7 161.3
R12 VP.n52 VP.n0 161.3
R13 VP.n51 VP.n50 161.3
R14 VP.n49 VP.n1 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n45 VP.n2 161.3
R17 VP.n44 VP.n43 161.3
R18 VP.n42 VP.n3 161.3
R19 VP.n41 VP.n40 161.3
R20 VP.n39 VP.n4 161.3
R21 VP.n37 VP.n36 161.3
R22 VP.n35 VP.n5 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n6 161.3
R25 VP.n13 VP.n12 67.1862
R26 VP.n12 VP.t2 57.1338
R27 VP.n33 VP.n5 45.3497
R28 VP.n51 VP.n1 45.3497
R29 VP.n26 VP.n8 45.3497
R30 VP.n40 VP.n3 40.4934
R31 VP.n44 VP.n3 40.4934
R32 VP.n19 VP.n10 40.4934
R33 VP.n15 VP.n10 40.4934
R34 VP.n30 VP.n29 39.0611
R35 VP.n37 VP.n5 35.6371
R36 VP.n47 VP.n1 35.6371
R37 VP.n22 VP.n8 35.6371
R38 VP.n31 VP.t0 27.6034
R39 VP.n38 VP.t3 27.6034
R40 VP.n46 VP.t5 27.6034
R41 VP.n53 VP.t7 27.6034
R42 VP.n28 VP.t1 27.6034
R43 VP.n21 VP.t4 27.6034
R44 VP.n13 VP.t6 27.6034
R45 VP.n33 VP.n32 24.4675
R46 VP.n40 VP.n39 24.4675
R47 VP.n45 VP.n44 24.4675
R48 VP.n52 VP.n51 24.4675
R49 VP.n27 VP.n26 24.4675
R50 VP.n20 VP.n19 24.4675
R51 VP.n15 VP.n14 24.4675
R52 VP.n38 VP.n37 23.2442
R53 VP.n47 VP.n46 23.2442
R54 VP.n22 VP.n21 23.2442
R55 VP.n12 VP.n11 18.6168
R56 VP.n32 VP.n31 3.67055
R57 VP.n53 VP.n52 3.67055
R58 VP.n28 VP.n27 3.67055
R59 VP.n39 VP.n38 1.22385
R60 VP.n46 VP.n45 1.22385
R61 VP.n21 VP.n20 1.22385
R62 VP.n14 VP.n13 1.22385
R63 VP.n16 VP.n11 0.189894
R64 VP.n17 VP.n16 0.189894
R65 VP.n18 VP.n17 0.189894
R66 VP.n18 VP.n9 0.189894
R67 VP.n23 VP.n9 0.189894
R68 VP.n24 VP.n23 0.189894
R69 VP.n25 VP.n24 0.189894
R70 VP.n25 VP.n7 0.189894
R71 VP.n29 VP.n7 0.189894
R72 VP.n30 VP.n6 0.189894
R73 VP.n34 VP.n6 0.189894
R74 VP.n35 VP.n34 0.189894
R75 VP.n36 VP.n35 0.189894
R76 VP.n36 VP.n4 0.189894
R77 VP.n41 VP.n4 0.189894
R78 VP.n42 VP.n41 0.189894
R79 VP.n43 VP.n42 0.189894
R80 VP.n43 VP.n2 0.189894
R81 VP.n48 VP.n2 0.189894
R82 VP.n49 VP.n48 0.189894
R83 VP.n50 VP.n49 0.189894
R84 VP.n50 VP.n0 0.189894
R85 VP.n54 VP.n0 0.189894
R86 VP VP.n54 0.0516364
R87 VDD1 VDD1.n0 101.156
R88 VDD1.n3 VDD1.n2 101.043
R89 VDD1.n3 VDD1.n1 101.043
R90 VDD1.n5 VDD1.n4 100.213
R91 VDD1.n5 VDD1.n3 33.9492
R92 VDD1.n4 VDD1.t2 10.0513
R93 VDD1.n4 VDD1.t6 10.0513
R94 VDD1.n0 VDD1.t5 10.0513
R95 VDD1.n0 VDD1.t1 10.0513
R96 VDD1.n2 VDD1.t4 10.0513
R97 VDD1.n2 VDD1.t7 10.0513
R98 VDD1.n1 VDD1.t0 10.0513
R99 VDD1.n1 VDD1.t3 10.0513
R100 VDD1 VDD1.n5 0.825931
R101 VTAIL.n66 VTAIL.n64 289.615
R102 VTAIL.n4 VTAIL.n2 289.615
R103 VTAIL.n12 VTAIL.n10 289.615
R104 VTAIL.n22 VTAIL.n20 289.615
R105 VTAIL.n58 VTAIL.n56 289.615
R106 VTAIL.n48 VTAIL.n46 289.615
R107 VTAIL.n40 VTAIL.n38 289.615
R108 VTAIL.n30 VTAIL.n28 289.615
R109 VTAIL.n67 VTAIL.n66 185
R110 VTAIL.n5 VTAIL.n4 185
R111 VTAIL.n13 VTAIL.n12 185
R112 VTAIL.n23 VTAIL.n22 185
R113 VTAIL.n59 VTAIL.n58 185
R114 VTAIL.n49 VTAIL.n48 185
R115 VTAIL.n41 VTAIL.n40 185
R116 VTAIL.n31 VTAIL.n30 185
R117 VTAIL.t6 VTAIL.n65 167.117
R118 VTAIL.t7 VTAIL.n3 167.117
R119 VTAIL.t8 VTAIL.n11 167.117
R120 VTAIL.t15 VTAIL.n21 167.117
R121 VTAIL.t14 VTAIL.n57 167.117
R122 VTAIL.t13 VTAIL.n47 167.117
R123 VTAIL.t2 VTAIL.n39 167.117
R124 VTAIL.t3 VTAIL.n29 167.117
R125 VTAIL.n55 VTAIL.n54 83.535
R126 VTAIL.n37 VTAIL.n36 83.535
R127 VTAIL.n1 VTAIL.n0 83.535
R128 VTAIL.n19 VTAIL.n18 83.535
R129 VTAIL.n66 VTAIL.t6 52.3082
R130 VTAIL.n4 VTAIL.t7 52.3082
R131 VTAIL.n12 VTAIL.t8 52.3082
R132 VTAIL.n22 VTAIL.t15 52.3082
R133 VTAIL.n58 VTAIL.t14 52.3082
R134 VTAIL.n48 VTAIL.t13 52.3082
R135 VTAIL.n40 VTAIL.t2 52.3082
R136 VTAIL.n30 VTAIL.t3 52.3082
R137 VTAIL.n71 VTAIL.n70 30.8278
R138 VTAIL.n9 VTAIL.n8 30.8278
R139 VTAIL.n17 VTAIL.n16 30.8278
R140 VTAIL.n27 VTAIL.n26 30.8278
R141 VTAIL.n63 VTAIL.n62 30.8278
R142 VTAIL.n53 VTAIL.n52 30.8278
R143 VTAIL.n45 VTAIL.n44 30.8278
R144 VTAIL.n35 VTAIL.n34 30.8278
R145 VTAIL.n71 VTAIL.n63 15.8324
R146 VTAIL.n35 VTAIL.n27 15.8324
R147 VTAIL.n0 VTAIL.t5 10.0513
R148 VTAIL.n0 VTAIL.t0 10.0513
R149 VTAIL.n18 VTAIL.t12 10.0513
R150 VTAIL.n18 VTAIL.t10 10.0513
R151 VTAIL.n54 VTAIL.t9 10.0513
R152 VTAIL.n54 VTAIL.t11 10.0513
R153 VTAIL.n36 VTAIL.t4 10.0513
R154 VTAIL.n36 VTAIL.t1 10.0513
R155 VTAIL.n67 VTAIL.n65 9.71174
R156 VTAIL.n5 VTAIL.n3 9.71174
R157 VTAIL.n13 VTAIL.n11 9.71174
R158 VTAIL.n23 VTAIL.n21 9.71174
R159 VTAIL.n59 VTAIL.n57 9.71174
R160 VTAIL.n49 VTAIL.n47 9.71174
R161 VTAIL.n41 VTAIL.n39 9.71174
R162 VTAIL.n31 VTAIL.n29 9.71174
R163 VTAIL.n70 VTAIL.n69 9.45567
R164 VTAIL.n8 VTAIL.n7 9.45567
R165 VTAIL.n16 VTAIL.n15 9.45567
R166 VTAIL.n26 VTAIL.n25 9.45567
R167 VTAIL.n62 VTAIL.n61 9.45567
R168 VTAIL.n52 VTAIL.n51 9.45567
R169 VTAIL.n44 VTAIL.n43 9.45567
R170 VTAIL.n34 VTAIL.n33 9.45567
R171 VTAIL.n69 VTAIL.n68 9.3005
R172 VTAIL.n7 VTAIL.n6 9.3005
R173 VTAIL.n15 VTAIL.n14 9.3005
R174 VTAIL.n25 VTAIL.n24 9.3005
R175 VTAIL.n61 VTAIL.n60 9.3005
R176 VTAIL.n51 VTAIL.n50 9.3005
R177 VTAIL.n43 VTAIL.n42 9.3005
R178 VTAIL.n33 VTAIL.n32 9.3005
R179 VTAIL.n70 VTAIL.n64 8.14595
R180 VTAIL.n8 VTAIL.n2 8.14595
R181 VTAIL.n16 VTAIL.n10 8.14595
R182 VTAIL.n26 VTAIL.n20 8.14595
R183 VTAIL.n62 VTAIL.n56 8.14595
R184 VTAIL.n52 VTAIL.n46 8.14595
R185 VTAIL.n44 VTAIL.n38 8.14595
R186 VTAIL.n34 VTAIL.n28 8.14595
R187 VTAIL.n68 VTAIL.n67 7.3702
R188 VTAIL.n6 VTAIL.n5 7.3702
R189 VTAIL.n14 VTAIL.n13 7.3702
R190 VTAIL.n24 VTAIL.n23 7.3702
R191 VTAIL.n60 VTAIL.n59 7.3702
R192 VTAIL.n50 VTAIL.n49 7.3702
R193 VTAIL.n42 VTAIL.n41 7.3702
R194 VTAIL.n32 VTAIL.n31 7.3702
R195 VTAIL.n68 VTAIL.n64 5.81868
R196 VTAIL.n6 VTAIL.n2 5.81868
R197 VTAIL.n14 VTAIL.n10 5.81868
R198 VTAIL.n24 VTAIL.n20 5.81868
R199 VTAIL.n60 VTAIL.n56 5.81868
R200 VTAIL.n50 VTAIL.n46 5.81868
R201 VTAIL.n42 VTAIL.n38 5.81868
R202 VTAIL.n32 VTAIL.n28 5.81868
R203 VTAIL.n69 VTAIL.n65 3.44771
R204 VTAIL.n7 VTAIL.n3 3.44771
R205 VTAIL.n15 VTAIL.n11 3.44771
R206 VTAIL.n25 VTAIL.n21 3.44771
R207 VTAIL.n61 VTAIL.n57 3.44771
R208 VTAIL.n51 VTAIL.n47 3.44771
R209 VTAIL.n43 VTAIL.n39 3.44771
R210 VTAIL.n33 VTAIL.n29 3.44771
R211 VTAIL.n37 VTAIL.n35 1.76774
R212 VTAIL.n45 VTAIL.n37 1.76774
R213 VTAIL.n55 VTAIL.n53 1.76774
R214 VTAIL.n63 VTAIL.n55 1.76774
R215 VTAIL.n27 VTAIL.n19 1.76774
R216 VTAIL.n19 VTAIL.n17 1.76774
R217 VTAIL.n9 VTAIL.n1 1.76774
R218 VTAIL VTAIL.n71 1.70955
R219 VTAIL.n53 VTAIL.n45 0.470328
R220 VTAIL.n17 VTAIL.n9 0.470328
R221 VTAIL VTAIL.n1 0.0586897
R222 B.n421 B.n420 585
R223 B.n423 B.n93 585
R224 B.n426 B.n425 585
R225 B.n427 B.n92 585
R226 B.n429 B.n428 585
R227 B.n431 B.n91 585
R228 B.n434 B.n433 585
R229 B.n435 B.n90 585
R230 B.n437 B.n436 585
R231 B.n439 B.n89 585
R232 B.n441 B.n440 585
R233 B.n443 B.n442 585
R234 B.n446 B.n445 585
R235 B.n447 B.n84 585
R236 B.n449 B.n448 585
R237 B.n451 B.n83 585
R238 B.n454 B.n453 585
R239 B.n455 B.n82 585
R240 B.n457 B.n456 585
R241 B.n459 B.n81 585
R242 B.n462 B.n461 585
R243 B.n463 B.n78 585
R244 B.n466 B.n465 585
R245 B.n468 B.n77 585
R246 B.n471 B.n470 585
R247 B.n472 B.n76 585
R248 B.n474 B.n473 585
R249 B.n476 B.n75 585
R250 B.n479 B.n478 585
R251 B.n480 B.n74 585
R252 B.n482 B.n481 585
R253 B.n484 B.n73 585
R254 B.n487 B.n486 585
R255 B.n488 B.n72 585
R256 B.n419 B.n70 585
R257 B.n491 B.n70 585
R258 B.n418 B.n69 585
R259 B.n492 B.n69 585
R260 B.n417 B.n68 585
R261 B.n493 B.n68 585
R262 B.n416 B.n415 585
R263 B.n415 B.n64 585
R264 B.n414 B.n63 585
R265 B.n499 B.n63 585
R266 B.n413 B.n62 585
R267 B.n500 B.n62 585
R268 B.n412 B.n61 585
R269 B.n501 B.n61 585
R270 B.n411 B.n410 585
R271 B.n410 B.n57 585
R272 B.n409 B.n56 585
R273 B.n507 B.n56 585
R274 B.n408 B.n55 585
R275 B.n508 B.n55 585
R276 B.n407 B.n54 585
R277 B.n509 B.n54 585
R278 B.n406 B.n405 585
R279 B.n405 B.n50 585
R280 B.n404 B.n49 585
R281 B.n515 B.n49 585
R282 B.n403 B.n48 585
R283 B.n516 B.n48 585
R284 B.n402 B.n47 585
R285 B.n517 B.n47 585
R286 B.n401 B.n400 585
R287 B.n400 B.n46 585
R288 B.n399 B.n42 585
R289 B.n523 B.n42 585
R290 B.n398 B.n41 585
R291 B.n524 B.n41 585
R292 B.n397 B.n40 585
R293 B.n525 B.n40 585
R294 B.n396 B.n395 585
R295 B.n395 B.n36 585
R296 B.n394 B.n35 585
R297 B.n531 B.n35 585
R298 B.n393 B.n34 585
R299 B.n532 B.n34 585
R300 B.n392 B.n33 585
R301 B.n533 B.n33 585
R302 B.n391 B.n390 585
R303 B.n390 B.n29 585
R304 B.n389 B.n28 585
R305 B.n539 B.n28 585
R306 B.n388 B.n27 585
R307 B.n540 B.n27 585
R308 B.n387 B.n26 585
R309 B.n541 B.n26 585
R310 B.n386 B.n385 585
R311 B.n385 B.n25 585
R312 B.n384 B.n21 585
R313 B.n547 B.n21 585
R314 B.n383 B.n20 585
R315 B.n548 B.n20 585
R316 B.n382 B.n19 585
R317 B.n549 B.n19 585
R318 B.n381 B.n380 585
R319 B.n380 B.n15 585
R320 B.n379 B.n14 585
R321 B.n555 B.n14 585
R322 B.n378 B.n13 585
R323 B.n556 B.n13 585
R324 B.n377 B.n12 585
R325 B.n557 B.n12 585
R326 B.n376 B.n375 585
R327 B.n375 B.n8 585
R328 B.n374 B.n7 585
R329 B.n563 B.n7 585
R330 B.n373 B.n6 585
R331 B.n564 B.n6 585
R332 B.n372 B.n5 585
R333 B.n565 B.n5 585
R334 B.n371 B.n370 585
R335 B.n370 B.n4 585
R336 B.n369 B.n94 585
R337 B.n369 B.n368 585
R338 B.n359 B.n95 585
R339 B.n96 B.n95 585
R340 B.n361 B.n360 585
R341 B.n362 B.n361 585
R342 B.n358 B.n100 585
R343 B.n104 B.n100 585
R344 B.n357 B.n356 585
R345 B.n356 B.n355 585
R346 B.n102 B.n101 585
R347 B.n103 B.n102 585
R348 B.n348 B.n347 585
R349 B.n349 B.n348 585
R350 B.n346 B.n109 585
R351 B.n109 B.n108 585
R352 B.n345 B.n344 585
R353 B.n344 B.n343 585
R354 B.n111 B.n110 585
R355 B.n336 B.n111 585
R356 B.n335 B.n334 585
R357 B.n337 B.n335 585
R358 B.n333 B.n116 585
R359 B.n116 B.n115 585
R360 B.n332 B.n331 585
R361 B.n331 B.n330 585
R362 B.n118 B.n117 585
R363 B.n119 B.n118 585
R364 B.n323 B.n322 585
R365 B.n324 B.n323 585
R366 B.n321 B.n123 585
R367 B.n127 B.n123 585
R368 B.n320 B.n319 585
R369 B.n319 B.n318 585
R370 B.n125 B.n124 585
R371 B.n126 B.n125 585
R372 B.n311 B.n310 585
R373 B.n312 B.n311 585
R374 B.n309 B.n132 585
R375 B.n132 B.n131 585
R376 B.n308 B.n307 585
R377 B.n307 B.n306 585
R378 B.n134 B.n133 585
R379 B.n299 B.n134 585
R380 B.n298 B.n297 585
R381 B.n300 B.n298 585
R382 B.n296 B.n139 585
R383 B.n139 B.n138 585
R384 B.n295 B.n294 585
R385 B.n294 B.n293 585
R386 B.n141 B.n140 585
R387 B.n142 B.n141 585
R388 B.n286 B.n285 585
R389 B.n287 B.n286 585
R390 B.n284 B.n147 585
R391 B.n147 B.n146 585
R392 B.n283 B.n282 585
R393 B.n282 B.n281 585
R394 B.n149 B.n148 585
R395 B.n150 B.n149 585
R396 B.n274 B.n273 585
R397 B.n275 B.n274 585
R398 B.n272 B.n155 585
R399 B.n155 B.n154 585
R400 B.n271 B.n270 585
R401 B.n270 B.n269 585
R402 B.n157 B.n156 585
R403 B.n158 B.n157 585
R404 B.n262 B.n261 585
R405 B.n263 B.n262 585
R406 B.n260 B.n163 585
R407 B.n163 B.n162 585
R408 B.n259 B.n258 585
R409 B.n258 B.n257 585
R410 B.n254 B.n167 585
R411 B.n253 B.n252 585
R412 B.n250 B.n168 585
R413 B.n250 B.n166 585
R414 B.n249 B.n248 585
R415 B.n247 B.n246 585
R416 B.n245 B.n170 585
R417 B.n243 B.n242 585
R418 B.n241 B.n171 585
R419 B.n240 B.n239 585
R420 B.n237 B.n172 585
R421 B.n235 B.n234 585
R422 B.n233 B.n173 585
R423 B.n231 B.n230 585
R424 B.n228 B.n176 585
R425 B.n226 B.n225 585
R426 B.n224 B.n177 585
R427 B.n223 B.n222 585
R428 B.n220 B.n178 585
R429 B.n218 B.n217 585
R430 B.n216 B.n179 585
R431 B.n215 B.n214 585
R432 B.n212 B.n180 585
R433 B.n210 B.n209 585
R434 B.n208 B.n181 585
R435 B.n207 B.n206 585
R436 B.n204 B.n185 585
R437 B.n202 B.n201 585
R438 B.n200 B.n186 585
R439 B.n199 B.n198 585
R440 B.n196 B.n187 585
R441 B.n194 B.n193 585
R442 B.n192 B.n188 585
R443 B.n191 B.n190 585
R444 B.n165 B.n164 585
R445 B.n166 B.n165 585
R446 B.n256 B.n255 585
R447 B.n257 B.n256 585
R448 B.n161 B.n160 585
R449 B.n162 B.n161 585
R450 B.n265 B.n264 585
R451 B.n264 B.n263 585
R452 B.n266 B.n159 585
R453 B.n159 B.n158 585
R454 B.n268 B.n267 585
R455 B.n269 B.n268 585
R456 B.n153 B.n152 585
R457 B.n154 B.n153 585
R458 B.n277 B.n276 585
R459 B.n276 B.n275 585
R460 B.n278 B.n151 585
R461 B.n151 B.n150 585
R462 B.n280 B.n279 585
R463 B.n281 B.n280 585
R464 B.n145 B.n144 585
R465 B.n146 B.n145 585
R466 B.n289 B.n288 585
R467 B.n288 B.n287 585
R468 B.n290 B.n143 585
R469 B.n143 B.n142 585
R470 B.n292 B.n291 585
R471 B.n293 B.n292 585
R472 B.n137 B.n136 585
R473 B.n138 B.n137 585
R474 B.n302 B.n301 585
R475 B.n301 B.n300 585
R476 B.n303 B.n135 585
R477 B.n299 B.n135 585
R478 B.n305 B.n304 585
R479 B.n306 B.n305 585
R480 B.n130 B.n129 585
R481 B.n131 B.n130 585
R482 B.n314 B.n313 585
R483 B.n313 B.n312 585
R484 B.n315 B.n128 585
R485 B.n128 B.n126 585
R486 B.n317 B.n316 585
R487 B.n318 B.n317 585
R488 B.n122 B.n121 585
R489 B.n127 B.n122 585
R490 B.n326 B.n325 585
R491 B.n325 B.n324 585
R492 B.n327 B.n120 585
R493 B.n120 B.n119 585
R494 B.n329 B.n328 585
R495 B.n330 B.n329 585
R496 B.n114 B.n113 585
R497 B.n115 B.n114 585
R498 B.n339 B.n338 585
R499 B.n338 B.n337 585
R500 B.n340 B.n112 585
R501 B.n336 B.n112 585
R502 B.n342 B.n341 585
R503 B.n343 B.n342 585
R504 B.n107 B.n106 585
R505 B.n108 B.n107 585
R506 B.n351 B.n350 585
R507 B.n350 B.n349 585
R508 B.n352 B.n105 585
R509 B.n105 B.n103 585
R510 B.n354 B.n353 585
R511 B.n355 B.n354 585
R512 B.n99 B.n98 585
R513 B.n104 B.n99 585
R514 B.n364 B.n363 585
R515 B.n363 B.n362 585
R516 B.n365 B.n97 585
R517 B.n97 B.n96 585
R518 B.n367 B.n366 585
R519 B.n368 B.n367 585
R520 B.n2 B.n0 585
R521 B.n4 B.n2 585
R522 B.n3 B.n1 585
R523 B.n564 B.n3 585
R524 B.n562 B.n561 585
R525 B.n563 B.n562 585
R526 B.n560 B.n9 585
R527 B.n9 B.n8 585
R528 B.n559 B.n558 585
R529 B.n558 B.n557 585
R530 B.n11 B.n10 585
R531 B.n556 B.n11 585
R532 B.n554 B.n553 585
R533 B.n555 B.n554 585
R534 B.n552 B.n16 585
R535 B.n16 B.n15 585
R536 B.n551 B.n550 585
R537 B.n550 B.n549 585
R538 B.n18 B.n17 585
R539 B.n548 B.n18 585
R540 B.n546 B.n545 585
R541 B.n547 B.n546 585
R542 B.n544 B.n22 585
R543 B.n25 B.n22 585
R544 B.n543 B.n542 585
R545 B.n542 B.n541 585
R546 B.n24 B.n23 585
R547 B.n540 B.n24 585
R548 B.n538 B.n537 585
R549 B.n539 B.n538 585
R550 B.n536 B.n30 585
R551 B.n30 B.n29 585
R552 B.n535 B.n534 585
R553 B.n534 B.n533 585
R554 B.n32 B.n31 585
R555 B.n532 B.n32 585
R556 B.n530 B.n529 585
R557 B.n531 B.n530 585
R558 B.n528 B.n37 585
R559 B.n37 B.n36 585
R560 B.n527 B.n526 585
R561 B.n526 B.n525 585
R562 B.n39 B.n38 585
R563 B.n524 B.n39 585
R564 B.n522 B.n521 585
R565 B.n523 B.n522 585
R566 B.n520 B.n43 585
R567 B.n46 B.n43 585
R568 B.n519 B.n518 585
R569 B.n518 B.n517 585
R570 B.n45 B.n44 585
R571 B.n516 B.n45 585
R572 B.n514 B.n513 585
R573 B.n515 B.n514 585
R574 B.n512 B.n51 585
R575 B.n51 B.n50 585
R576 B.n511 B.n510 585
R577 B.n510 B.n509 585
R578 B.n53 B.n52 585
R579 B.n508 B.n53 585
R580 B.n506 B.n505 585
R581 B.n507 B.n506 585
R582 B.n504 B.n58 585
R583 B.n58 B.n57 585
R584 B.n503 B.n502 585
R585 B.n502 B.n501 585
R586 B.n60 B.n59 585
R587 B.n500 B.n60 585
R588 B.n498 B.n497 585
R589 B.n499 B.n498 585
R590 B.n496 B.n65 585
R591 B.n65 B.n64 585
R592 B.n495 B.n494 585
R593 B.n494 B.n493 585
R594 B.n67 B.n66 585
R595 B.n492 B.n67 585
R596 B.n490 B.n489 585
R597 B.n491 B.n490 585
R598 B.n567 B.n566 585
R599 B.n566 B.n565 585
R600 B.n256 B.n167 526.135
R601 B.n490 B.n72 526.135
R602 B.n258 B.n165 526.135
R603 B.n421 B.n70 526.135
R604 B.n422 B.n71 256.663
R605 B.n424 B.n71 256.663
R606 B.n430 B.n71 256.663
R607 B.n432 B.n71 256.663
R608 B.n438 B.n71 256.663
R609 B.n88 B.n71 256.663
R610 B.n444 B.n71 256.663
R611 B.n450 B.n71 256.663
R612 B.n452 B.n71 256.663
R613 B.n458 B.n71 256.663
R614 B.n460 B.n71 256.663
R615 B.n467 B.n71 256.663
R616 B.n469 B.n71 256.663
R617 B.n475 B.n71 256.663
R618 B.n477 B.n71 256.663
R619 B.n483 B.n71 256.663
R620 B.n485 B.n71 256.663
R621 B.n251 B.n166 256.663
R622 B.n169 B.n166 256.663
R623 B.n244 B.n166 256.663
R624 B.n238 B.n166 256.663
R625 B.n236 B.n166 256.663
R626 B.n229 B.n166 256.663
R627 B.n227 B.n166 256.663
R628 B.n221 B.n166 256.663
R629 B.n219 B.n166 256.663
R630 B.n213 B.n166 256.663
R631 B.n211 B.n166 256.663
R632 B.n205 B.n166 256.663
R633 B.n203 B.n166 256.663
R634 B.n197 B.n166 256.663
R635 B.n195 B.n166 256.663
R636 B.n189 B.n166 256.663
R637 B.n182 B.t19 233.778
R638 B.n174 B.t15 233.778
R639 B.n79 B.t8 233.778
R640 B.n85 B.t12 233.778
R641 B.n257 B.n166 214.079
R642 B.n491 B.n71 214.079
R643 B.n256 B.n161 163.367
R644 B.n264 B.n161 163.367
R645 B.n264 B.n159 163.367
R646 B.n268 B.n159 163.367
R647 B.n268 B.n153 163.367
R648 B.n276 B.n153 163.367
R649 B.n276 B.n151 163.367
R650 B.n280 B.n151 163.367
R651 B.n280 B.n145 163.367
R652 B.n288 B.n145 163.367
R653 B.n288 B.n143 163.367
R654 B.n292 B.n143 163.367
R655 B.n292 B.n137 163.367
R656 B.n301 B.n137 163.367
R657 B.n301 B.n135 163.367
R658 B.n305 B.n135 163.367
R659 B.n305 B.n130 163.367
R660 B.n313 B.n130 163.367
R661 B.n313 B.n128 163.367
R662 B.n317 B.n128 163.367
R663 B.n317 B.n122 163.367
R664 B.n325 B.n122 163.367
R665 B.n325 B.n120 163.367
R666 B.n329 B.n120 163.367
R667 B.n329 B.n114 163.367
R668 B.n338 B.n114 163.367
R669 B.n338 B.n112 163.367
R670 B.n342 B.n112 163.367
R671 B.n342 B.n107 163.367
R672 B.n350 B.n107 163.367
R673 B.n350 B.n105 163.367
R674 B.n354 B.n105 163.367
R675 B.n354 B.n99 163.367
R676 B.n363 B.n99 163.367
R677 B.n363 B.n97 163.367
R678 B.n367 B.n97 163.367
R679 B.n367 B.n2 163.367
R680 B.n566 B.n2 163.367
R681 B.n566 B.n3 163.367
R682 B.n562 B.n3 163.367
R683 B.n562 B.n9 163.367
R684 B.n558 B.n9 163.367
R685 B.n558 B.n11 163.367
R686 B.n554 B.n11 163.367
R687 B.n554 B.n16 163.367
R688 B.n550 B.n16 163.367
R689 B.n550 B.n18 163.367
R690 B.n546 B.n18 163.367
R691 B.n546 B.n22 163.367
R692 B.n542 B.n22 163.367
R693 B.n542 B.n24 163.367
R694 B.n538 B.n24 163.367
R695 B.n538 B.n30 163.367
R696 B.n534 B.n30 163.367
R697 B.n534 B.n32 163.367
R698 B.n530 B.n32 163.367
R699 B.n530 B.n37 163.367
R700 B.n526 B.n37 163.367
R701 B.n526 B.n39 163.367
R702 B.n522 B.n39 163.367
R703 B.n522 B.n43 163.367
R704 B.n518 B.n43 163.367
R705 B.n518 B.n45 163.367
R706 B.n514 B.n45 163.367
R707 B.n514 B.n51 163.367
R708 B.n510 B.n51 163.367
R709 B.n510 B.n53 163.367
R710 B.n506 B.n53 163.367
R711 B.n506 B.n58 163.367
R712 B.n502 B.n58 163.367
R713 B.n502 B.n60 163.367
R714 B.n498 B.n60 163.367
R715 B.n498 B.n65 163.367
R716 B.n494 B.n65 163.367
R717 B.n494 B.n67 163.367
R718 B.n490 B.n67 163.367
R719 B.n252 B.n250 163.367
R720 B.n250 B.n249 163.367
R721 B.n246 B.n245 163.367
R722 B.n243 B.n171 163.367
R723 B.n239 B.n237 163.367
R724 B.n235 B.n173 163.367
R725 B.n230 B.n228 163.367
R726 B.n226 B.n177 163.367
R727 B.n222 B.n220 163.367
R728 B.n218 B.n179 163.367
R729 B.n214 B.n212 163.367
R730 B.n210 B.n181 163.367
R731 B.n206 B.n204 163.367
R732 B.n202 B.n186 163.367
R733 B.n198 B.n196 163.367
R734 B.n194 B.n188 163.367
R735 B.n190 B.n165 163.367
R736 B.n258 B.n163 163.367
R737 B.n262 B.n163 163.367
R738 B.n262 B.n157 163.367
R739 B.n270 B.n157 163.367
R740 B.n270 B.n155 163.367
R741 B.n274 B.n155 163.367
R742 B.n274 B.n149 163.367
R743 B.n282 B.n149 163.367
R744 B.n282 B.n147 163.367
R745 B.n286 B.n147 163.367
R746 B.n286 B.n141 163.367
R747 B.n294 B.n141 163.367
R748 B.n294 B.n139 163.367
R749 B.n298 B.n139 163.367
R750 B.n298 B.n134 163.367
R751 B.n307 B.n134 163.367
R752 B.n307 B.n132 163.367
R753 B.n311 B.n132 163.367
R754 B.n311 B.n125 163.367
R755 B.n319 B.n125 163.367
R756 B.n319 B.n123 163.367
R757 B.n323 B.n123 163.367
R758 B.n323 B.n118 163.367
R759 B.n331 B.n118 163.367
R760 B.n331 B.n116 163.367
R761 B.n335 B.n116 163.367
R762 B.n335 B.n111 163.367
R763 B.n344 B.n111 163.367
R764 B.n344 B.n109 163.367
R765 B.n348 B.n109 163.367
R766 B.n348 B.n102 163.367
R767 B.n356 B.n102 163.367
R768 B.n356 B.n100 163.367
R769 B.n361 B.n100 163.367
R770 B.n361 B.n95 163.367
R771 B.n369 B.n95 163.367
R772 B.n370 B.n369 163.367
R773 B.n370 B.n5 163.367
R774 B.n6 B.n5 163.367
R775 B.n7 B.n6 163.367
R776 B.n375 B.n7 163.367
R777 B.n375 B.n12 163.367
R778 B.n13 B.n12 163.367
R779 B.n14 B.n13 163.367
R780 B.n380 B.n14 163.367
R781 B.n380 B.n19 163.367
R782 B.n20 B.n19 163.367
R783 B.n21 B.n20 163.367
R784 B.n385 B.n21 163.367
R785 B.n385 B.n26 163.367
R786 B.n27 B.n26 163.367
R787 B.n28 B.n27 163.367
R788 B.n390 B.n28 163.367
R789 B.n390 B.n33 163.367
R790 B.n34 B.n33 163.367
R791 B.n35 B.n34 163.367
R792 B.n395 B.n35 163.367
R793 B.n395 B.n40 163.367
R794 B.n41 B.n40 163.367
R795 B.n42 B.n41 163.367
R796 B.n400 B.n42 163.367
R797 B.n400 B.n47 163.367
R798 B.n48 B.n47 163.367
R799 B.n49 B.n48 163.367
R800 B.n405 B.n49 163.367
R801 B.n405 B.n54 163.367
R802 B.n55 B.n54 163.367
R803 B.n56 B.n55 163.367
R804 B.n410 B.n56 163.367
R805 B.n410 B.n61 163.367
R806 B.n62 B.n61 163.367
R807 B.n63 B.n62 163.367
R808 B.n415 B.n63 163.367
R809 B.n415 B.n68 163.367
R810 B.n69 B.n68 163.367
R811 B.n70 B.n69 163.367
R812 B.n486 B.n484 163.367
R813 B.n482 B.n74 163.367
R814 B.n478 B.n476 163.367
R815 B.n474 B.n76 163.367
R816 B.n470 B.n468 163.367
R817 B.n466 B.n78 163.367
R818 B.n461 B.n459 163.367
R819 B.n457 B.n82 163.367
R820 B.n453 B.n451 163.367
R821 B.n449 B.n84 163.367
R822 B.n445 B.n443 163.367
R823 B.n440 B.n439 163.367
R824 B.n437 B.n90 163.367
R825 B.n433 B.n431 163.367
R826 B.n429 B.n92 163.367
R827 B.n425 B.n423 163.367
R828 B.n182 B.t21 162.195
R829 B.n85 B.t13 162.195
R830 B.n174 B.t18 162.195
R831 B.n79 B.t10 162.195
R832 B.n183 B.t20 122.436
R833 B.n86 B.t14 122.436
R834 B.n175 B.t17 122.436
R835 B.n80 B.t11 122.436
R836 B.n257 B.n162 103.245
R837 B.n263 B.n162 103.245
R838 B.n263 B.n158 103.245
R839 B.n269 B.n158 103.245
R840 B.n269 B.n154 103.245
R841 B.n275 B.n154 103.245
R842 B.n281 B.n150 103.245
R843 B.n281 B.n146 103.245
R844 B.n287 B.n146 103.245
R845 B.n287 B.n142 103.245
R846 B.n293 B.n142 103.245
R847 B.n293 B.n138 103.245
R848 B.n300 B.n138 103.245
R849 B.n300 B.n299 103.245
R850 B.n306 B.n131 103.245
R851 B.n312 B.n131 103.245
R852 B.n312 B.n126 103.245
R853 B.n318 B.n126 103.245
R854 B.n318 B.n127 103.245
R855 B.n324 B.n119 103.245
R856 B.n330 B.n119 103.245
R857 B.n330 B.n115 103.245
R858 B.n337 B.n115 103.245
R859 B.n337 B.n336 103.245
R860 B.n343 B.n108 103.245
R861 B.n349 B.n108 103.245
R862 B.n349 B.n103 103.245
R863 B.n355 B.n103 103.245
R864 B.n355 B.n104 103.245
R865 B.n362 B.n96 103.245
R866 B.n368 B.n96 103.245
R867 B.n368 B.n4 103.245
R868 B.n565 B.n4 103.245
R869 B.n565 B.n564 103.245
R870 B.n564 B.n563 103.245
R871 B.n563 B.n8 103.245
R872 B.n557 B.n8 103.245
R873 B.n556 B.n555 103.245
R874 B.n555 B.n15 103.245
R875 B.n549 B.n15 103.245
R876 B.n549 B.n548 103.245
R877 B.n548 B.n547 103.245
R878 B.n541 B.n25 103.245
R879 B.n541 B.n540 103.245
R880 B.n540 B.n539 103.245
R881 B.n539 B.n29 103.245
R882 B.n533 B.n29 103.245
R883 B.n532 B.n531 103.245
R884 B.n531 B.n36 103.245
R885 B.n525 B.n36 103.245
R886 B.n525 B.n524 103.245
R887 B.n524 B.n523 103.245
R888 B.n517 B.n46 103.245
R889 B.n517 B.n516 103.245
R890 B.n516 B.n515 103.245
R891 B.n515 B.n50 103.245
R892 B.n509 B.n50 103.245
R893 B.n509 B.n508 103.245
R894 B.n508 B.n507 103.245
R895 B.n507 B.n57 103.245
R896 B.n501 B.n500 103.245
R897 B.n500 B.n499 103.245
R898 B.n499 B.n64 103.245
R899 B.n493 B.n64 103.245
R900 B.n493 B.n492 103.245
R901 B.n492 B.n491 103.245
R902 B.t16 B.n150 97.171
R903 B.t9 B.n57 97.171
R904 B.n306 B.t3 72.8783
R905 B.n523 B.t6 72.8783
R906 B.n251 B.n167 71.676
R907 B.n249 B.n169 71.676
R908 B.n245 B.n244 71.676
R909 B.n238 B.n171 71.676
R910 B.n237 B.n236 71.676
R911 B.n229 B.n173 71.676
R912 B.n228 B.n227 71.676
R913 B.n221 B.n177 71.676
R914 B.n220 B.n219 71.676
R915 B.n213 B.n179 71.676
R916 B.n212 B.n211 71.676
R917 B.n205 B.n181 71.676
R918 B.n204 B.n203 71.676
R919 B.n197 B.n186 71.676
R920 B.n196 B.n195 71.676
R921 B.n189 B.n188 71.676
R922 B.n485 B.n72 71.676
R923 B.n484 B.n483 71.676
R924 B.n477 B.n74 71.676
R925 B.n476 B.n475 71.676
R926 B.n469 B.n76 71.676
R927 B.n468 B.n467 71.676
R928 B.n460 B.n78 71.676
R929 B.n459 B.n458 71.676
R930 B.n452 B.n82 71.676
R931 B.n451 B.n450 71.676
R932 B.n444 B.n84 71.676
R933 B.n443 B.n88 71.676
R934 B.n439 B.n438 71.676
R935 B.n432 B.n90 71.676
R936 B.n431 B.n430 71.676
R937 B.n424 B.n92 71.676
R938 B.n423 B.n422 71.676
R939 B.n422 B.n421 71.676
R940 B.n425 B.n424 71.676
R941 B.n430 B.n429 71.676
R942 B.n433 B.n432 71.676
R943 B.n438 B.n437 71.676
R944 B.n440 B.n88 71.676
R945 B.n445 B.n444 71.676
R946 B.n450 B.n449 71.676
R947 B.n453 B.n452 71.676
R948 B.n458 B.n457 71.676
R949 B.n461 B.n460 71.676
R950 B.n467 B.n466 71.676
R951 B.n470 B.n469 71.676
R952 B.n475 B.n474 71.676
R953 B.n478 B.n477 71.676
R954 B.n483 B.n482 71.676
R955 B.n486 B.n485 71.676
R956 B.n252 B.n251 71.676
R957 B.n246 B.n169 71.676
R958 B.n244 B.n243 71.676
R959 B.n239 B.n238 71.676
R960 B.n236 B.n235 71.676
R961 B.n230 B.n229 71.676
R962 B.n227 B.n226 71.676
R963 B.n222 B.n221 71.676
R964 B.n219 B.n218 71.676
R965 B.n214 B.n213 71.676
R966 B.n211 B.n210 71.676
R967 B.n206 B.n205 71.676
R968 B.n203 B.n202 71.676
R969 B.n198 B.n197 71.676
R970 B.n195 B.n194 71.676
R971 B.n190 B.n189 71.676
R972 B.n324 B.t4 69.8418
R973 B.n533 B.t0 69.8418
R974 B.n343 B.t1 66.8052
R975 B.n547 B.t5 66.8052
R976 B.n362 B.t2 63.7686
R977 B.n557 B.t7 63.7686
R978 B.n184 B.n183 59.5399
R979 B.n232 B.n175 59.5399
R980 B.n464 B.n80 59.5399
R981 B.n87 B.n86 59.5399
R982 B.n183 B.n182 39.7581
R983 B.n175 B.n174 39.7581
R984 B.n80 B.n79 39.7581
R985 B.n86 B.n85 39.7581
R986 B.n104 B.t2 39.476
R987 B.t7 B.n556 39.476
R988 B.n336 B.t1 36.4394
R989 B.n25 B.t5 36.4394
R990 B.n489 B.n488 34.1859
R991 B.n420 B.n419 34.1859
R992 B.n259 B.n164 34.1859
R993 B.n255 B.n254 34.1859
R994 B.n127 B.t4 33.4028
R995 B.t0 B.n532 33.4028
R996 B.n299 B.t3 30.3663
R997 B.n46 B.t6 30.3663
R998 B B.n567 18.0485
R999 B.n488 B.n487 10.6151
R1000 B.n487 B.n73 10.6151
R1001 B.n481 B.n73 10.6151
R1002 B.n481 B.n480 10.6151
R1003 B.n480 B.n479 10.6151
R1004 B.n479 B.n75 10.6151
R1005 B.n473 B.n75 10.6151
R1006 B.n473 B.n472 10.6151
R1007 B.n472 B.n471 10.6151
R1008 B.n471 B.n77 10.6151
R1009 B.n465 B.n77 10.6151
R1010 B.n463 B.n462 10.6151
R1011 B.n462 B.n81 10.6151
R1012 B.n456 B.n81 10.6151
R1013 B.n456 B.n455 10.6151
R1014 B.n455 B.n454 10.6151
R1015 B.n454 B.n83 10.6151
R1016 B.n448 B.n83 10.6151
R1017 B.n448 B.n447 10.6151
R1018 B.n447 B.n446 10.6151
R1019 B.n442 B.n441 10.6151
R1020 B.n441 B.n89 10.6151
R1021 B.n436 B.n89 10.6151
R1022 B.n436 B.n435 10.6151
R1023 B.n435 B.n434 10.6151
R1024 B.n434 B.n91 10.6151
R1025 B.n428 B.n91 10.6151
R1026 B.n428 B.n427 10.6151
R1027 B.n427 B.n426 10.6151
R1028 B.n426 B.n93 10.6151
R1029 B.n420 B.n93 10.6151
R1030 B.n260 B.n259 10.6151
R1031 B.n261 B.n260 10.6151
R1032 B.n261 B.n156 10.6151
R1033 B.n271 B.n156 10.6151
R1034 B.n272 B.n271 10.6151
R1035 B.n273 B.n272 10.6151
R1036 B.n273 B.n148 10.6151
R1037 B.n283 B.n148 10.6151
R1038 B.n284 B.n283 10.6151
R1039 B.n285 B.n284 10.6151
R1040 B.n285 B.n140 10.6151
R1041 B.n295 B.n140 10.6151
R1042 B.n296 B.n295 10.6151
R1043 B.n297 B.n296 10.6151
R1044 B.n297 B.n133 10.6151
R1045 B.n308 B.n133 10.6151
R1046 B.n309 B.n308 10.6151
R1047 B.n310 B.n309 10.6151
R1048 B.n310 B.n124 10.6151
R1049 B.n320 B.n124 10.6151
R1050 B.n321 B.n320 10.6151
R1051 B.n322 B.n321 10.6151
R1052 B.n322 B.n117 10.6151
R1053 B.n332 B.n117 10.6151
R1054 B.n333 B.n332 10.6151
R1055 B.n334 B.n333 10.6151
R1056 B.n334 B.n110 10.6151
R1057 B.n345 B.n110 10.6151
R1058 B.n346 B.n345 10.6151
R1059 B.n347 B.n346 10.6151
R1060 B.n347 B.n101 10.6151
R1061 B.n357 B.n101 10.6151
R1062 B.n358 B.n357 10.6151
R1063 B.n360 B.n358 10.6151
R1064 B.n360 B.n359 10.6151
R1065 B.n359 B.n94 10.6151
R1066 B.n371 B.n94 10.6151
R1067 B.n372 B.n371 10.6151
R1068 B.n373 B.n372 10.6151
R1069 B.n374 B.n373 10.6151
R1070 B.n376 B.n374 10.6151
R1071 B.n377 B.n376 10.6151
R1072 B.n378 B.n377 10.6151
R1073 B.n379 B.n378 10.6151
R1074 B.n381 B.n379 10.6151
R1075 B.n382 B.n381 10.6151
R1076 B.n383 B.n382 10.6151
R1077 B.n384 B.n383 10.6151
R1078 B.n386 B.n384 10.6151
R1079 B.n387 B.n386 10.6151
R1080 B.n388 B.n387 10.6151
R1081 B.n389 B.n388 10.6151
R1082 B.n391 B.n389 10.6151
R1083 B.n392 B.n391 10.6151
R1084 B.n393 B.n392 10.6151
R1085 B.n394 B.n393 10.6151
R1086 B.n396 B.n394 10.6151
R1087 B.n397 B.n396 10.6151
R1088 B.n398 B.n397 10.6151
R1089 B.n399 B.n398 10.6151
R1090 B.n401 B.n399 10.6151
R1091 B.n402 B.n401 10.6151
R1092 B.n403 B.n402 10.6151
R1093 B.n404 B.n403 10.6151
R1094 B.n406 B.n404 10.6151
R1095 B.n407 B.n406 10.6151
R1096 B.n408 B.n407 10.6151
R1097 B.n409 B.n408 10.6151
R1098 B.n411 B.n409 10.6151
R1099 B.n412 B.n411 10.6151
R1100 B.n413 B.n412 10.6151
R1101 B.n414 B.n413 10.6151
R1102 B.n416 B.n414 10.6151
R1103 B.n417 B.n416 10.6151
R1104 B.n418 B.n417 10.6151
R1105 B.n419 B.n418 10.6151
R1106 B.n254 B.n253 10.6151
R1107 B.n253 B.n168 10.6151
R1108 B.n248 B.n168 10.6151
R1109 B.n248 B.n247 10.6151
R1110 B.n247 B.n170 10.6151
R1111 B.n242 B.n170 10.6151
R1112 B.n242 B.n241 10.6151
R1113 B.n241 B.n240 10.6151
R1114 B.n240 B.n172 10.6151
R1115 B.n234 B.n172 10.6151
R1116 B.n234 B.n233 10.6151
R1117 B.n231 B.n176 10.6151
R1118 B.n225 B.n176 10.6151
R1119 B.n225 B.n224 10.6151
R1120 B.n224 B.n223 10.6151
R1121 B.n223 B.n178 10.6151
R1122 B.n217 B.n178 10.6151
R1123 B.n217 B.n216 10.6151
R1124 B.n216 B.n215 10.6151
R1125 B.n215 B.n180 10.6151
R1126 B.n209 B.n208 10.6151
R1127 B.n208 B.n207 10.6151
R1128 B.n207 B.n185 10.6151
R1129 B.n201 B.n185 10.6151
R1130 B.n201 B.n200 10.6151
R1131 B.n200 B.n199 10.6151
R1132 B.n199 B.n187 10.6151
R1133 B.n193 B.n187 10.6151
R1134 B.n193 B.n192 10.6151
R1135 B.n192 B.n191 10.6151
R1136 B.n191 B.n164 10.6151
R1137 B.n255 B.n160 10.6151
R1138 B.n265 B.n160 10.6151
R1139 B.n266 B.n265 10.6151
R1140 B.n267 B.n266 10.6151
R1141 B.n267 B.n152 10.6151
R1142 B.n277 B.n152 10.6151
R1143 B.n278 B.n277 10.6151
R1144 B.n279 B.n278 10.6151
R1145 B.n279 B.n144 10.6151
R1146 B.n289 B.n144 10.6151
R1147 B.n290 B.n289 10.6151
R1148 B.n291 B.n290 10.6151
R1149 B.n291 B.n136 10.6151
R1150 B.n302 B.n136 10.6151
R1151 B.n303 B.n302 10.6151
R1152 B.n304 B.n303 10.6151
R1153 B.n304 B.n129 10.6151
R1154 B.n314 B.n129 10.6151
R1155 B.n315 B.n314 10.6151
R1156 B.n316 B.n315 10.6151
R1157 B.n316 B.n121 10.6151
R1158 B.n326 B.n121 10.6151
R1159 B.n327 B.n326 10.6151
R1160 B.n328 B.n327 10.6151
R1161 B.n328 B.n113 10.6151
R1162 B.n339 B.n113 10.6151
R1163 B.n340 B.n339 10.6151
R1164 B.n341 B.n340 10.6151
R1165 B.n341 B.n106 10.6151
R1166 B.n351 B.n106 10.6151
R1167 B.n352 B.n351 10.6151
R1168 B.n353 B.n352 10.6151
R1169 B.n353 B.n98 10.6151
R1170 B.n364 B.n98 10.6151
R1171 B.n365 B.n364 10.6151
R1172 B.n366 B.n365 10.6151
R1173 B.n366 B.n0 10.6151
R1174 B.n561 B.n1 10.6151
R1175 B.n561 B.n560 10.6151
R1176 B.n560 B.n559 10.6151
R1177 B.n559 B.n10 10.6151
R1178 B.n553 B.n10 10.6151
R1179 B.n553 B.n552 10.6151
R1180 B.n552 B.n551 10.6151
R1181 B.n551 B.n17 10.6151
R1182 B.n545 B.n17 10.6151
R1183 B.n545 B.n544 10.6151
R1184 B.n544 B.n543 10.6151
R1185 B.n543 B.n23 10.6151
R1186 B.n537 B.n23 10.6151
R1187 B.n537 B.n536 10.6151
R1188 B.n536 B.n535 10.6151
R1189 B.n535 B.n31 10.6151
R1190 B.n529 B.n31 10.6151
R1191 B.n529 B.n528 10.6151
R1192 B.n528 B.n527 10.6151
R1193 B.n527 B.n38 10.6151
R1194 B.n521 B.n38 10.6151
R1195 B.n521 B.n520 10.6151
R1196 B.n520 B.n519 10.6151
R1197 B.n519 B.n44 10.6151
R1198 B.n513 B.n44 10.6151
R1199 B.n513 B.n512 10.6151
R1200 B.n512 B.n511 10.6151
R1201 B.n511 B.n52 10.6151
R1202 B.n505 B.n52 10.6151
R1203 B.n505 B.n504 10.6151
R1204 B.n504 B.n503 10.6151
R1205 B.n503 B.n59 10.6151
R1206 B.n497 B.n59 10.6151
R1207 B.n497 B.n496 10.6151
R1208 B.n496 B.n495 10.6151
R1209 B.n495 B.n66 10.6151
R1210 B.n489 B.n66 10.6151
R1211 B.n465 B.n464 9.36635
R1212 B.n442 B.n87 9.36635
R1213 B.n233 B.n232 9.36635
R1214 B.n209 B.n184 9.36635
R1215 B.n275 B.t16 6.07365
R1216 B.n501 B.t9 6.07365
R1217 B.n567 B.n0 2.81026
R1218 B.n567 B.n1 2.81026
R1219 B.n464 B.n463 1.24928
R1220 B.n446 B.n87 1.24928
R1221 B.n232 B.n231 1.24928
R1222 B.n184 B.n180 1.24928
R1223 VN.n22 VN.n21 182.097
R1224 VN.n45 VN.n44 182.097
R1225 VN.n43 VN.n23 161.3
R1226 VN.n42 VN.n41 161.3
R1227 VN.n40 VN.n24 161.3
R1228 VN.n39 VN.n38 161.3
R1229 VN.n36 VN.n25 161.3
R1230 VN.n35 VN.n34 161.3
R1231 VN.n33 VN.n26 161.3
R1232 VN.n32 VN.n31 161.3
R1233 VN.n30 VN.n27 161.3
R1234 VN.n20 VN.n0 161.3
R1235 VN.n19 VN.n18 161.3
R1236 VN.n17 VN.n1 161.3
R1237 VN.n16 VN.n15 161.3
R1238 VN.n13 VN.n2 161.3
R1239 VN.n12 VN.n11 161.3
R1240 VN.n10 VN.n3 161.3
R1241 VN.n9 VN.n8 161.3
R1242 VN.n7 VN.n4 161.3
R1243 VN.n6 VN.n5 67.1862
R1244 VN.n29 VN.n28 67.1862
R1245 VN.n5 VN.t1 57.1338
R1246 VN.n28 VN.t5 57.1338
R1247 VN.n19 VN.n1 45.3497
R1248 VN.n42 VN.n24 45.3497
R1249 VN.n8 VN.n3 40.4934
R1250 VN.n12 VN.n3 40.4934
R1251 VN.n31 VN.n26 40.4934
R1252 VN.n35 VN.n26 40.4934
R1253 VN VN.n45 39.4418
R1254 VN.n15 VN.n1 35.6371
R1255 VN.n38 VN.n24 35.6371
R1256 VN.n6 VN.t7 27.6034
R1257 VN.n14 VN.t4 27.6034
R1258 VN.n21 VN.t0 27.6034
R1259 VN.n29 VN.t2 27.6034
R1260 VN.n37 VN.t6 27.6034
R1261 VN.n44 VN.t3 27.6034
R1262 VN.n8 VN.n7 24.4675
R1263 VN.n13 VN.n12 24.4675
R1264 VN.n20 VN.n19 24.4675
R1265 VN.n31 VN.n30 24.4675
R1266 VN.n36 VN.n35 24.4675
R1267 VN.n43 VN.n42 24.4675
R1268 VN.n15 VN.n14 23.2442
R1269 VN.n38 VN.n37 23.2442
R1270 VN.n28 VN.n27 18.6168
R1271 VN.n5 VN.n4 18.6168
R1272 VN.n21 VN.n20 3.67055
R1273 VN.n44 VN.n43 3.67055
R1274 VN.n7 VN.n6 1.22385
R1275 VN.n14 VN.n13 1.22385
R1276 VN.n30 VN.n29 1.22385
R1277 VN.n37 VN.n36 1.22385
R1278 VN.n45 VN.n23 0.189894
R1279 VN.n41 VN.n23 0.189894
R1280 VN.n41 VN.n40 0.189894
R1281 VN.n40 VN.n39 0.189894
R1282 VN.n39 VN.n25 0.189894
R1283 VN.n34 VN.n25 0.189894
R1284 VN.n34 VN.n33 0.189894
R1285 VN.n33 VN.n32 0.189894
R1286 VN.n32 VN.n27 0.189894
R1287 VN.n9 VN.n4 0.189894
R1288 VN.n10 VN.n9 0.189894
R1289 VN.n11 VN.n10 0.189894
R1290 VN.n11 VN.n2 0.189894
R1291 VN.n16 VN.n2 0.189894
R1292 VN.n17 VN.n16 0.189894
R1293 VN.n18 VN.n17 0.189894
R1294 VN.n18 VN.n0 0.189894
R1295 VN.n22 VN.n0 0.189894
R1296 VN VN.n22 0.0516364
R1297 VDD2.n2 VDD2.n1 101.043
R1298 VDD2.n2 VDD2.n0 101.043
R1299 VDD2 VDD2.n5 101.04
R1300 VDD2.n4 VDD2.n3 100.213
R1301 VDD2.n4 VDD2.n2 33.3662
R1302 VDD2.n5 VDD2.t5 10.0513
R1303 VDD2.n5 VDD2.t2 10.0513
R1304 VDD2.n3 VDD2.t4 10.0513
R1305 VDD2.n3 VDD2.t1 10.0513
R1306 VDD2.n1 VDD2.t3 10.0513
R1307 VDD2.n1 VDD2.t7 10.0513
R1308 VDD2.n0 VDD2.t6 10.0513
R1309 VDD2.n0 VDD2.t0 10.0513
R1310 VDD2 VDD2.n4 0.94231
C0 VN VDD1 0.155646f
C1 VP VDD1 1.93505f
C2 VTAIL VDD2 4.02665f
C3 VN VDD2 1.66026f
C4 VTAIL VN 2.39105f
C5 VDD2 VP 0.432519f
C6 VTAIL VP 2.40516f
C7 VDD2 VDD1 1.31716f
C8 VN VP 4.73709f
C9 VTAIL VDD1 3.97813f
C10 VDD2 B 3.531549f
C11 VDD1 B 3.861558f
C12 VTAIL B 3.591138f
C13 VN B 10.96921f
C14 VP B 9.728958f
C15 VDD2.t6 B 0.026746f
C16 VDD2.t0 B 0.026746f
C17 VDD2.n0 B 0.170082f
C18 VDD2.t3 B 0.026746f
C19 VDD2.t7 B 0.026746f
C20 VDD2.n1 B 0.170082f
C21 VDD2.n2 B 1.46888f
C22 VDD2.t4 B 0.026746f
C23 VDD2.t1 B 0.026746f
C24 VDD2.n3 B 0.167775f
C25 VDD2.n4 B 1.26271f
C26 VDD2.t5 B 0.026746f
C27 VDD2.t2 B 0.026746f
C28 VDD2.n5 B 0.17007f
C29 VN.n0 B 0.02887f
C30 VN.t0 B 0.227762f
C31 VN.n1 B 0.024279f
C32 VN.n2 B 0.02887f
C33 VN.t4 B 0.227762f
C34 VN.n3 B 0.023339f
C35 VN.n4 B 0.18474f
C36 VN.t7 B 0.227762f
C37 VN.t1 B 0.352358f
C38 VN.n5 B 0.175827f
C39 VN.n6 B 0.168007f
C40 VN.n7 B 0.028569f
C41 VN.n8 B 0.057379f
C42 VN.n9 B 0.02887f
C43 VN.n10 B 0.02887f
C44 VN.n11 B 0.02887f
C45 VN.n12 B 0.057379f
C46 VN.n13 B 0.028569f
C47 VN.n14 B 0.117945f
C48 VN.n15 B 0.056972f
C49 VN.n16 B 0.02887f
C50 VN.n17 B 0.02887f
C51 VN.n18 B 0.02887f
C52 VN.n19 B 0.055517f
C53 VN.n20 B 0.031225f
C54 VN.n21 B 0.179489f
C55 VN.n22 B 0.030308f
C56 VN.n23 B 0.02887f
C57 VN.t3 B 0.227762f
C58 VN.n24 B 0.024279f
C59 VN.n25 B 0.02887f
C60 VN.t6 B 0.227762f
C61 VN.n26 B 0.023339f
C62 VN.n27 B 0.18474f
C63 VN.t2 B 0.227762f
C64 VN.t5 B 0.352358f
C65 VN.n28 B 0.175827f
C66 VN.n29 B 0.168007f
C67 VN.n30 B 0.028569f
C68 VN.n31 B 0.057379f
C69 VN.n32 B 0.02887f
C70 VN.n33 B 0.02887f
C71 VN.n34 B 0.02887f
C72 VN.n35 B 0.057379f
C73 VN.n36 B 0.028569f
C74 VN.n37 B 0.117945f
C75 VN.n38 B 0.056972f
C76 VN.n39 B 0.02887f
C77 VN.n40 B 0.02887f
C78 VN.n41 B 0.02887f
C79 VN.n42 B 0.055517f
C80 VN.n43 B 0.031225f
C81 VN.n44 B 0.179489f
C82 VN.n45 B 1.07962f
C83 VTAIL.t5 B 0.045854f
C84 VTAIL.t0 B 0.045854f
C85 VTAIL.n0 B 0.244102f
C86 VTAIL.n1 B 0.400368f
C87 VTAIL.n2 B 0.042395f
C88 VTAIL.n3 B 0.094008f
C89 VTAIL.t7 B 0.070636f
C90 VTAIL.n4 B 0.073393f
C91 VTAIL.n5 B 0.023999f
C92 VTAIL.n6 B 0.015828f
C93 VTAIL.n7 B 0.206057f
C94 VTAIL.n8 B 0.046392f
C95 VTAIL.n9 B 0.235888f
C96 VTAIL.n10 B 0.042395f
C97 VTAIL.n11 B 0.094008f
C98 VTAIL.t8 B 0.070636f
C99 VTAIL.n12 B 0.073393f
C100 VTAIL.n13 B 0.023999f
C101 VTAIL.n14 B 0.015828f
C102 VTAIL.n15 B 0.206057f
C103 VTAIL.n16 B 0.046392f
C104 VTAIL.n17 B 0.235888f
C105 VTAIL.t12 B 0.045854f
C106 VTAIL.t10 B 0.045854f
C107 VTAIL.n18 B 0.244102f
C108 VTAIL.n19 B 0.562573f
C109 VTAIL.n20 B 0.042395f
C110 VTAIL.n21 B 0.094008f
C111 VTAIL.t15 B 0.070636f
C112 VTAIL.n22 B 0.073393f
C113 VTAIL.n23 B 0.023999f
C114 VTAIL.n24 B 0.015828f
C115 VTAIL.n25 B 0.206057f
C116 VTAIL.n26 B 0.046392f
C117 VTAIL.n27 B 0.920315f
C118 VTAIL.n28 B 0.042395f
C119 VTAIL.n29 B 0.094008f
C120 VTAIL.t3 B 0.070636f
C121 VTAIL.n30 B 0.073393f
C122 VTAIL.n31 B 0.023999f
C123 VTAIL.n32 B 0.015828f
C124 VTAIL.n33 B 0.206057f
C125 VTAIL.n34 B 0.046392f
C126 VTAIL.n35 B 0.920315f
C127 VTAIL.t4 B 0.045854f
C128 VTAIL.t1 B 0.045854f
C129 VTAIL.n36 B 0.244104f
C130 VTAIL.n37 B 0.562572f
C131 VTAIL.n38 B 0.042395f
C132 VTAIL.n39 B 0.094008f
C133 VTAIL.t2 B 0.070636f
C134 VTAIL.n40 B 0.073393f
C135 VTAIL.n41 B 0.023999f
C136 VTAIL.n42 B 0.015828f
C137 VTAIL.n43 B 0.206057f
C138 VTAIL.n44 B 0.046392f
C139 VTAIL.n45 B 0.235888f
C140 VTAIL.n46 B 0.042395f
C141 VTAIL.n47 B 0.094008f
C142 VTAIL.t13 B 0.070636f
C143 VTAIL.n48 B 0.073393f
C144 VTAIL.n49 B 0.023999f
C145 VTAIL.n50 B 0.015828f
C146 VTAIL.n51 B 0.206057f
C147 VTAIL.n52 B 0.046392f
C148 VTAIL.n53 B 0.235888f
C149 VTAIL.t9 B 0.045854f
C150 VTAIL.t11 B 0.045854f
C151 VTAIL.n54 B 0.244104f
C152 VTAIL.n55 B 0.562572f
C153 VTAIL.n56 B 0.042395f
C154 VTAIL.n57 B 0.094008f
C155 VTAIL.t14 B 0.070636f
C156 VTAIL.n58 B 0.073393f
C157 VTAIL.n59 B 0.023999f
C158 VTAIL.n60 B 0.015828f
C159 VTAIL.n61 B 0.206057f
C160 VTAIL.n62 B 0.046392f
C161 VTAIL.n63 B 0.920315f
C162 VTAIL.n64 B 0.042395f
C163 VTAIL.n65 B 0.094008f
C164 VTAIL.t6 B 0.070636f
C165 VTAIL.n66 B 0.073393f
C166 VTAIL.n67 B 0.023999f
C167 VTAIL.n68 B 0.015828f
C168 VTAIL.n69 B 0.206057f
C169 VTAIL.n70 B 0.046392f
C170 VTAIL.n71 B 0.914792f
C171 VDD1.t5 B 0.026329f
C172 VDD1.t1 B 0.026329f
C173 VDD1.n0 B 0.167788f
C174 VDD1.t0 B 0.026329f
C175 VDD1.t3 B 0.026329f
C176 VDD1.n1 B 0.167426f
C177 VDD1.t4 B 0.026329f
C178 VDD1.t7 B 0.026329f
C179 VDD1.n2 B 0.167426f
C180 VDD1.n3 B 1.48168f
C181 VDD1.t2 B 0.026329f
C182 VDD1.t6 B 0.026329f
C183 VDD1.n4 B 0.165155f
C184 VDD1.n5 B 1.26338f
C185 VP.n0 B 0.029036f
C186 VP.t7 B 0.229071f
C187 VP.n1 B 0.024419f
C188 VP.n2 B 0.029036f
C189 VP.t5 B 0.229071f
C190 VP.n3 B 0.023473f
C191 VP.n4 B 0.029036f
C192 VP.t3 B 0.229071f
C193 VP.n5 B 0.024419f
C194 VP.n6 B 0.029036f
C195 VP.t0 B 0.229071f
C196 VP.n7 B 0.029036f
C197 VP.t1 B 0.229071f
C198 VP.n8 B 0.024419f
C199 VP.n9 B 0.029036f
C200 VP.t4 B 0.229071f
C201 VP.n10 B 0.023473f
C202 VP.n11 B 0.185802f
C203 VP.t6 B 0.229071f
C204 VP.t2 B 0.354384f
C205 VP.n12 B 0.176838f
C206 VP.n13 B 0.168973f
C207 VP.n14 B 0.028733f
C208 VP.n15 B 0.057709f
C209 VP.n16 B 0.029036f
C210 VP.n17 B 0.029036f
C211 VP.n18 B 0.029036f
C212 VP.n19 B 0.057709f
C213 VP.n20 B 0.028733f
C214 VP.n21 B 0.118623f
C215 VP.n22 B 0.057299f
C216 VP.n23 B 0.029036f
C217 VP.n24 B 0.029036f
C218 VP.n25 B 0.029036f
C219 VP.n26 B 0.055836f
C220 VP.n27 B 0.031405f
C221 VP.n28 B 0.180521f
C222 VP.n29 B 1.06668f
C223 VP.n30 B 1.0934f
C224 VP.n31 B 0.180521f
C225 VP.n32 B 0.031405f
C226 VP.n33 B 0.055836f
C227 VP.n34 B 0.029036f
C228 VP.n35 B 0.029036f
C229 VP.n36 B 0.029036f
C230 VP.n37 B 0.057299f
C231 VP.n38 B 0.118623f
C232 VP.n39 B 0.028733f
C233 VP.n40 B 0.057709f
C234 VP.n41 B 0.029036f
C235 VP.n42 B 0.029036f
C236 VP.n43 B 0.029036f
C237 VP.n44 B 0.057709f
C238 VP.n45 B 0.028733f
C239 VP.n46 B 0.118623f
C240 VP.n47 B 0.057299f
C241 VP.n48 B 0.029036f
C242 VP.n49 B 0.029036f
C243 VP.n50 B 0.029036f
C244 VP.n51 B 0.055836f
C245 VP.n52 B 0.031405f
C246 VP.n53 B 0.180521f
C247 VP.n54 B 0.030483f
.ends

