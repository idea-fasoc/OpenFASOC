* NGSPICE file created from diff_pair_sample_0233.ext - technology: sky130A

.subckt diff_pair_sample_0233 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=6.6339 ps=34.8 w=17.01 l=1.01
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=6.6339 ps=34.8 w=17.01 l=1.01
X2 B.t11 B.t9 B.t10 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=0 ps=0 w=17.01 l=1.01
X3 B.t8 B.t6 B.t7 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=0 ps=0 w=17.01 l=1.01
X4 VDD1.t0 VP.t1 VTAIL.t0 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=6.6339 ps=34.8 w=17.01 l=1.01
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=6.6339 ps=34.8 w=17.01 l=1.01
X6 B.t5 B.t3 B.t4 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=0 ps=0 w=17.01 l=1.01
X7 B.t2 B.t0 B.t1 w_n1506_n4374# sky130_fd_pr__pfet_01v8 ad=6.6339 pd=34.8 as=0 ps=0 w=17.01 l=1.01
R0 VN VN.t1 650.946
R1 VN VN.t0 606.366
R2 VTAIL.n1 VTAIL.t3 58.073
R3 VTAIL.n3 VTAIL.t2 58.072
R4 VTAIL.n0 VTAIL.t0 58.072
R5 VTAIL.n2 VTAIL.t1 58.0719
R6 VTAIL.n1 VTAIL.n0 29.3583
R7 VTAIL.n3 VTAIL.n2 28.2031
R8 VTAIL.n2 VTAIL.n1 1.04791
R9 VTAIL VTAIL.n0 0.81731
R10 VTAIL VTAIL.n3 0.231103
R11 VDD2.n0 VDD2.t1 115.401
R12 VDD2.n0 VDD2.t0 74.7506
R13 VDD2 VDD2.n0 0.347483
R14 VP.n0 VP.t0 650.566
R15 VP.n0 VP.t1 606.316
R16 VP VP.n0 0.0516364
R17 VDD1 VDD1.t0 116.216
R18 VDD1 VDD1.t1 75.0976
R19 B.n120 B.t0 608.876
R20 B.n128 B.t3 608.876
R21 B.n38 B.t6 608.876
R22 B.n46 B.t9 608.876
R23 B.n422 B.n75 585
R24 B.n424 B.n423 585
R25 B.n425 B.n74 585
R26 B.n427 B.n426 585
R27 B.n428 B.n73 585
R28 B.n430 B.n429 585
R29 B.n431 B.n72 585
R30 B.n433 B.n432 585
R31 B.n434 B.n71 585
R32 B.n436 B.n435 585
R33 B.n437 B.n70 585
R34 B.n439 B.n438 585
R35 B.n440 B.n69 585
R36 B.n442 B.n441 585
R37 B.n443 B.n68 585
R38 B.n445 B.n444 585
R39 B.n446 B.n67 585
R40 B.n448 B.n447 585
R41 B.n449 B.n66 585
R42 B.n451 B.n450 585
R43 B.n452 B.n65 585
R44 B.n454 B.n453 585
R45 B.n455 B.n64 585
R46 B.n457 B.n456 585
R47 B.n458 B.n63 585
R48 B.n460 B.n459 585
R49 B.n461 B.n62 585
R50 B.n463 B.n462 585
R51 B.n464 B.n61 585
R52 B.n466 B.n465 585
R53 B.n467 B.n60 585
R54 B.n469 B.n468 585
R55 B.n470 B.n59 585
R56 B.n472 B.n471 585
R57 B.n473 B.n58 585
R58 B.n475 B.n474 585
R59 B.n476 B.n57 585
R60 B.n478 B.n477 585
R61 B.n479 B.n56 585
R62 B.n481 B.n480 585
R63 B.n482 B.n55 585
R64 B.n484 B.n483 585
R65 B.n485 B.n54 585
R66 B.n487 B.n486 585
R67 B.n488 B.n53 585
R68 B.n490 B.n489 585
R69 B.n491 B.n52 585
R70 B.n493 B.n492 585
R71 B.n494 B.n51 585
R72 B.n496 B.n495 585
R73 B.n497 B.n50 585
R74 B.n499 B.n498 585
R75 B.n500 B.n49 585
R76 B.n502 B.n501 585
R77 B.n503 B.n48 585
R78 B.n505 B.n504 585
R79 B.n507 B.n45 585
R80 B.n509 B.n508 585
R81 B.n510 B.n44 585
R82 B.n512 B.n511 585
R83 B.n513 B.n43 585
R84 B.n515 B.n514 585
R85 B.n516 B.n42 585
R86 B.n518 B.n517 585
R87 B.n519 B.n41 585
R88 B.n521 B.n520 585
R89 B.n523 B.n522 585
R90 B.n524 B.n37 585
R91 B.n526 B.n525 585
R92 B.n527 B.n36 585
R93 B.n529 B.n528 585
R94 B.n530 B.n35 585
R95 B.n532 B.n531 585
R96 B.n533 B.n34 585
R97 B.n535 B.n534 585
R98 B.n536 B.n33 585
R99 B.n538 B.n537 585
R100 B.n539 B.n32 585
R101 B.n541 B.n540 585
R102 B.n542 B.n31 585
R103 B.n544 B.n543 585
R104 B.n545 B.n30 585
R105 B.n547 B.n546 585
R106 B.n548 B.n29 585
R107 B.n550 B.n549 585
R108 B.n551 B.n28 585
R109 B.n553 B.n552 585
R110 B.n554 B.n27 585
R111 B.n556 B.n555 585
R112 B.n557 B.n26 585
R113 B.n559 B.n558 585
R114 B.n560 B.n25 585
R115 B.n562 B.n561 585
R116 B.n563 B.n24 585
R117 B.n565 B.n564 585
R118 B.n566 B.n23 585
R119 B.n568 B.n567 585
R120 B.n569 B.n22 585
R121 B.n571 B.n570 585
R122 B.n572 B.n21 585
R123 B.n574 B.n573 585
R124 B.n575 B.n20 585
R125 B.n577 B.n576 585
R126 B.n578 B.n19 585
R127 B.n580 B.n579 585
R128 B.n581 B.n18 585
R129 B.n583 B.n582 585
R130 B.n584 B.n17 585
R131 B.n586 B.n585 585
R132 B.n587 B.n16 585
R133 B.n589 B.n588 585
R134 B.n590 B.n15 585
R135 B.n592 B.n591 585
R136 B.n593 B.n14 585
R137 B.n595 B.n594 585
R138 B.n596 B.n13 585
R139 B.n598 B.n597 585
R140 B.n599 B.n12 585
R141 B.n601 B.n600 585
R142 B.n602 B.n11 585
R143 B.n604 B.n603 585
R144 B.n605 B.n10 585
R145 B.n421 B.n420 585
R146 B.n419 B.n76 585
R147 B.n418 B.n417 585
R148 B.n416 B.n77 585
R149 B.n415 B.n414 585
R150 B.n413 B.n78 585
R151 B.n412 B.n411 585
R152 B.n410 B.n79 585
R153 B.n409 B.n408 585
R154 B.n407 B.n80 585
R155 B.n406 B.n405 585
R156 B.n404 B.n81 585
R157 B.n403 B.n402 585
R158 B.n401 B.n82 585
R159 B.n400 B.n399 585
R160 B.n398 B.n83 585
R161 B.n397 B.n396 585
R162 B.n395 B.n84 585
R163 B.n394 B.n393 585
R164 B.n392 B.n85 585
R165 B.n391 B.n390 585
R166 B.n389 B.n86 585
R167 B.n388 B.n387 585
R168 B.n386 B.n87 585
R169 B.n385 B.n384 585
R170 B.n383 B.n88 585
R171 B.n382 B.n381 585
R172 B.n380 B.n89 585
R173 B.n379 B.n378 585
R174 B.n377 B.n90 585
R175 B.n376 B.n375 585
R176 B.n374 B.n91 585
R177 B.n373 B.n372 585
R178 B.n188 B.n157 585
R179 B.n190 B.n189 585
R180 B.n191 B.n156 585
R181 B.n193 B.n192 585
R182 B.n194 B.n155 585
R183 B.n196 B.n195 585
R184 B.n197 B.n154 585
R185 B.n199 B.n198 585
R186 B.n200 B.n153 585
R187 B.n202 B.n201 585
R188 B.n203 B.n152 585
R189 B.n205 B.n204 585
R190 B.n206 B.n151 585
R191 B.n208 B.n207 585
R192 B.n209 B.n150 585
R193 B.n211 B.n210 585
R194 B.n212 B.n149 585
R195 B.n214 B.n213 585
R196 B.n215 B.n148 585
R197 B.n217 B.n216 585
R198 B.n218 B.n147 585
R199 B.n220 B.n219 585
R200 B.n221 B.n146 585
R201 B.n223 B.n222 585
R202 B.n224 B.n145 585
R203 B.n226 B.n225 585
R204 B.n227 B.n144 585
R205 B.n229 B.n228 585
R206 B.n230 B.n143 585
R207 B.n232 B.n231 585
R208 B.n233 B.n142 585
R209 B.n235 B.n234 585
R210 B.n236 B.n141 585
R211 B.n238 B.n237 585
R212 B.n239 B.n140 585
R213 B.n241 B.n240 585
R214 B.n242 B.n139 585
R215 B.n244 B.n243 585
R216 B.n245 B.n138 585
R217 B.n247 B.n246 585
R218 B.n248 B.n137 585
R219 B.n250 B.n249 585
R220 B.n251 B.n136 585
R221 B.n253 B.n252 585
R222 B.n254 B.n135 585
R223 B.n256 B.n255 585
R224 B.n257 B.n134 585
R225 B.n259 B.n258 585
R226 B.n260 B.n133 585
R227 B.n262 B.n261 585
R228 B.n263 B.n132 585
R229 B.n265 B.n264 585
R230 B.n266 B.n131 585
R231 B.n268 B.n267 585
R232 B.n269 B.n130 585
R233 B.n271 B.n270 585
R234 B.n273 B.n127 585
R235 B.n275 B.n274 585
R236 B.n276 B.n126 585
R237 B.n278 B.n277 585
R238 B.n279 B.n125 585
R239 B.n281 B.n280 585
R240 B.n282 B.n124 585
R241 B.n284 B.n283 585
R242 B.n285 B.n123 585
R243 B.n287 B.n286 585
R244 B.n289 B.n288 585
R245 B.n290 B.n119 585
R246 B.n292 B.n291 585
R247 B.n293 B.n118 585
R248 B.n295 B.n294 585
R249 B.n296 B.n117 585
R250 B.n298 B.n297 585
R251 B.n299 B.n116 585
R252 B.n301 B.n300 585
R253 B.n302 B.n115 585
R254 B.n304 B.n303 585
R255 B.n305 B.n114 585
R256 B.n307 B.n306 585
R257 B.n308 B.n113 585
R258 B.n310 B.n309 585
R259 B.n311 B.n112 585
R260 B.n313 B.n312 585
R261 B.n314 B.n111 585
R262 B.n316 B.n315 585
R263 B.n317 B.n110 585
R264 B.n319 B.n318 585
R265 B.n320 B.n109 585
R266 B.n322 B.n321 585
R267 B.n323 B.n108 585
R268 B.n325 B.n324 585
R269 B.n326 B.n107 585
R270 B.n328 B.n327 585
R271 B.n329 B.n106 585
R272 B.n331 B.n330 585
R273 B.n332 B.n105 585
R274 B.n334 B.n333 585
R275 B.n335 B.n104 585
R276 B.n337 B.n336 585
R277 B.n338 B.n103 585
R278 B.n340 B.n339 585
R279 B.n341 B.n102 585
R280 B.n343 B.n342 585
R281 B.n344 B.n101 585
R282 B.n346 B.n345 585
R283 B.n347 B.n100 585
R284 B.n349 B.n348 585
R285 B.n350 B.n99 585
R286 B.n352 B.n351 585
R287 B.n353 B.n98 585
R288 B.n355 B.n354 585
R289 B.n356 B.n97 585
R290 B.n358 B.n357 585
R291 B.n359 B.n96 585
R292 B.n361 B.n360 585
R293 B.n362 B.n95 585
R294 B.n364 B.n363 585
R295 B.n365 B.n94 585
R296 B.n367 B.n366 585
R297 B.n368 B.n93 585
R298 B.n370 B.n369 585
R299 B.n371 B.n92 585
R300 B.n187 B.n186 585
R301 B.n185 B.n158 585
R302 B.n184 B.n183 585
R303 B.n182 B.n159 585
R304 B.n181 B.n180 585
R305 B.n179 B.n160 585
R306 B.n178 B.n177 585
R307 B.n176 B.n161 585
R308 B.n175 B.n174 585
R309 B.n173 B.n162 585
R310 B.n172 B.n171 585
R311 B.n170 B.n163 585
R312 B.n169 B.n168 585
R313 B.n167 B.n164 585
R314 B.n166 B.n165 585
R315 B.n2 B.n0 585
R316 B.n629 B.n1 585
R317 B.n628 B.n627 585
R318 B.n626 B.n3 585
R319 B.n625 B.n624 585
R320 B.n623 B.n4 585
R321 B.n622 B.n621 585
R322 B.n620 B.n5 585
R323 B.n619 B.n618 585
R324 B.n617 B.n6 585
R325 B.n616 B.n615 585
R326 B.n614 B.n7 585
R327 B.n613 B.n612 585
R328 B.n611 B.n8 585
R329 B.n610 B.n609 585
R330 B.n608 B.n9 585
R331 B.n607 B.n606 585
R332 B.n631 B.n630 585
R333 B.n186 B.n157 530.939
R334 B.n606 B.n605 530.939
R335 B.n372 B.n371 530.939
R336 B.n420 B.n75 530.939
R337 B.n186 B.n185 163.367
R338 B.n185 B.n184 163.367
R339 B.n184 B.n159 163.367
R340 B.n180 B.n159 163.367
R341 B.n180 B.n179 163.367
R342 B.n179 B.n178 163.367
R343 B.n178 B.n161 163.367
R344 B.n174 B.n161 163.367
R345 B.n174 B.n173 163.367
R346 B.n173 B.n172 163.367
R347 B.n172 B.n163 163.367
R348 B.n168 B.n163 163.367
R349 B.n168 B.n167 163.367
R350 B.n167 B.n166 163.367
R351 B.n166 B.n2 163.367
R352 B.n630 B.n2 163.367
R353 B.n630 B.n629 163.367
R354 B.n629 B.n628 163.367
R355 B.n628 B.n3 163.367
R356 B.n624 B.n3 163.367
R357 B.n624 B.n623 163.367
R358 B.n623 B.n622 163.367
R359 B.n622 B.n5 163.367
R360 B.n618 B.n5 163.367
R361 B.n618 B.n617 163.367
R362 B.n617 B.n616 163.367
R363 B.n616 B.n7 163.367
R364 B.n612 B.n7 163.367
R365 B.n612 B.n611 163.367
R366 B.n611 B.n610 163.367
R367 B.n610 B.n9 163.367
R368 B.n606 B.n9 163.367
R369 B.n190 B.n157 163.367
R370 B.n191 B.n190 163.367
R371 B.n192 B.n191 163.367
R372 B.n192 B.n155 163.367
R373 B.n196 B.n155 163.367
R374 B.n197 B.n196 163.367
R375 B.n198 B.n197 163.367
R376 B.n198 B.n153 163.367
R377 B.n202 B.n153 163.367
R378 B.n203 B.n202 163.367
R379 B.n204 B.n203 163.367
R380 B.n204 B.n151 163.367
R381 B.n208 B.n151 163.367
R382 B.n209 B.n208 163.367
R383 B.n210 B.n209 163.367
R384 B.n210 B.n149 163.367
R385 B.n214 B.n149 163.367
R386 B.n215 B.n214 163.367
R387 B.n216 B.n215 163.367
R388 B.n216 B.n147 163.367
R389 B.n220 B.n147 163.367
R390 B.n221 B.n220 163.367
R391 B.n222 B.n221 163.367
R392 B.n222 B.n145 163.367
R393 B.n226 B.n145 163.367
R394 B.n227 B.n226 163.367
R395 B.n228 B.n227 163.367
R396 B.n228 B.n143 163.367
R397 B.n232 B.n143 163.367
R398 B.n233 B.n232 163.367
R399 B.n234 B.n233 163.367
R400 B.n234 B.n141 163.367
R401 B.n238 B.n141 163.367
R402 B.n239 B.n238 163.367
R403 B.n240 B.n239 163.367
R404 B.n240 B.n139 163.367
R405 B.n244 B.n139 163.367
R406 B.n245 B.n244 163.367
R407 B.n246 B.n245 163.367
R408 B.n246 B.n137 163.367
R409 B.n250 B.n137 163.367
R410 B.n251 B.n250 163.367
R411 B.n252 B.n251 163.367
R412 B.n252 B.n135 163.367
R413 B.n256 B.n135 163.367
R414 B.n257 B.n256 163.367
R415 B.n258 B.n257 163.367
R416 B.n258 B.n133 163.367
R417 B.n262 B.n133 163.367
R418 B.n263 B.n262 163.367
R419 B.n264 B.n263 163.367
R420 B.n264 B.n131 163.367
R421 B.n268 B.n131 163.367
R422 B.n269 B.n268 163.367
R423 B.n270 B.n269 163.367
R424 B.n270 B.n127 163.367
R425 B.n275 B.n127 163.367
R426 B.n276 B.n275 163.367
R427 B.n277 B.n276 163.367
R428 B.n277 B.n125 163.367
R429 B.n281 B.n125 163.367
R430 B.n282 B.n281 163.367
R431 B.n283 B.n282 163.367
R432 B.n283 B.n123 163.367
R433 B.n287 B.n123 163.367
R434 B.n288 B.n287 163.367
R435 B.n288 B.n119 163.367
R436 B.n292 B.n119 163.367
R437 B.n293 B.n292 163.367
R438 B.n294 B.n293 163.367
R439 B.n294 B.n117 163.367
R440 B.n298 B.n117 163.367
R441 B.n299 B.n298 163.367
R442 B.n300 B.n299 163.367
R443 B.n300 B.n115 163.367
R444 B.n304 B.n115 163.367
R445 B.n305 B.n304 163.367
R446 B.n306 B.n305 163.367
R447 B.n306 B.n113 163.367
R448 B.n310 B.n113 163.367
R449 B.n311 B.n310 163.367
R450 B.n312 B.n311 163.367
R451 B.n312 B.n111 163.367
R452 B.n316 B.n111 163.367
R453 B.n317 B.n316 163.367
R454 B.n318 B.n317 163.367
R455 B.n318 B.n109 163.367
R456 B.n322 B.n109 163.367
R457 B.n323 B.n322 163.367
R458 B.n324 B.n323 163.367
R459 B.n324 B.n107 163.367
R460 B.n328 B.n107 163.367
R461 B.n329 B.n328 163.367
R462 B.n330 B.n329 163.367
R463 B.n330 B.n105 163.367
R464 B.n334 B.n105 163.367
R465 B.n335 B.n334 163.367
R466 B.n336 B.n335 163.367
R467 B.n336 B.n103 163.367
R468 B.n340 B.n103 163.367
R469 B.n341 B.n340 163.367
R470 B.n342 B.n341 163.367
R471 B.n342 B.n101 163.367
R472 B.n346 B.n101 163.367
R473 B.n347 B.n346 163.367
R474 B.n348 B.n347 163.367
R475 B.n348 B.n99 163.367
R476 B.n352 B.n99 163.367
R477 B.n353 B.n352 163.367
R478 B.n354 B.n353 163.367
R479 B.n354 B.n97 163.367
R480 B.n358 B.n97 163.367
R481 B.n359 B.n358 163.367
R482 B.n360 B.n359 163.367
R483 B.n360 B.n95 163.367
R484 B.n364 B.n95 163.367
R485 B.n365 B.n364 163.367
R486 B.n366 B.n365 163.367
R487 B.n366 B.n93 163.367
R488 B.n370 B.n93 163.367
R489 B.n371 B.n370 163.367
R490 B.n372 B.n91 163.367
R491 B.n376 B.n91 163.367
R492 B.n377 B.n376 163.367
R493 B.n378 B.n377 163.367
R494 B.n378 B.n89 163.367
R495 B.n382 B.n89 163.367
R496 B.n383 B.n382 163.367
R497 B.n384 B.n383 163.367
R498 B.n384 B.n87 163.367
R499 B.n388 B.n87 163.367
R500 B.n389 B.n388 163.367
R501 B.n390 B.n389 163.367
R502 B.n390 B.n85 163.367
R503 B.n394 B.n85 163.367
R504 B.n395 B.n394 163.367
R505 B.n396 B.n395 163.367
R506 B.n396 B.n83 163.367
R507 B.n400 B.n83 163.367
R508 B.n401 B.n400 163.367
R509 B.n402 B.n401 163.367
R510 B.n402 B.n81 163.367
R511 B.n406 B.n81 163.367
R512 B.n407 B.n406 163.367
R513 B.n408 B.n407 163.367
R514 B.n408 B.n79 163.367
R515 B.n412 B.n79 163.367
R516 B.n413 B.n412 163.367
R517 B.n414 B.n413 163.367
R518 B.n414 B.n77 163.367
R519 B.n418 B.n77 163.367
R520 B.n419 B.n418 163.367
R521 B.n420 B.n419 163.367
R522 B.n605 B.n604 163.367
R523 B.n604 B.n11 163.367
R524 B.n600 B.n11 163.367
R525 B.n600 B.n599 163.367
R526 B.n599 B.n598 163.367
R527 B.n598 B.n13 163.367
R528 B.n594 B.n13 163.367
R529 B.n594 B.n593 163.367
R530 B.n593 B.n592 163.367
R531 B.n592 B.n15 163.367
R532 B.n588 B.n15 163.367
R533 B.n588 B.n587 163.367
R534 B.n587 B.n586 163.367
R535 B.n586 B.n17 163.367
R536 B.n582 B.n17 163.367
R537 B.n582 B.n581 163.367
R538 B.n581 B.n580 163.367
R539 B.n580 B.n19 163.367
R540 B.n576 B.n19 163.367
R541 B.n576 B.n575 163.367
R542 B.n575 B.n574 163.367
R543 B.n574 B.n21 163.367
R544 B.n570 B.n21 163.367
R545 B.n570 B.n569 163.367
R546 B.n569 B.n568 163.367
R547 B.n568 B.n23 163.367
R548 B.n564 B.n23 163.367
R549 B.n564 B.n563 163.367
R550 B.n563 B.n562 163.367
R551 B.n562 B.n25 163.367
R552 B.n558 B.n25 163.367
R553 B.n558 B.n557 163.367
R554 B.n557 B.n556 163.367
R555 B.n556 B.n27 163.367
R556 B.n552 B.n27 163.367
R557 B.n552 B.n551 163.367
R558 B.n551 B.n550 163.367
R559 B.n550 B.n29 163.367
R560 B.n546 B.n29 163.367
R561 B.n546 B.n545 163.367
R562 B.n545 B.n544 163.367
R563 B.n544 B.n31 163.367
R564 B.n540 B.n31 163.367
R565 B.n540 B.n539 163.367
R566 B.n539 B.n538 163.367
R567 B.n538 B.n33 163.367
R568 B.n534 B.n33 163.367
R569 B.n534 B.n533 163.367
R570 B.n533 B.n532 163.367
R571 B.n532 B.n35 163.367
R572 B.n528 B.n35 163.367
R573 B.n528 B.n527 163.367
R574 B.n527 B.n526 163.367
R575 B.n526 B.n37 163.367
R576 B.n522 B.n37 163.367
R577 B.n522 B.n521 163.367
R578 B.n521 B.n41 163.367
R579 B.n517 B.n41 163.367
R580 B.n517 B.n516 163.367
R581 B.n516 B.n515 163.367
R582 B.n515 B.n43 163.367
R583 B.n511 B.n43 163.367
R584 B.n511 B.n510 163.367
R585 B.n510 B.n509 163.367
R586 B.n509 B.n45 163.367
R587 B.n504 B.n45 163.367
R588 B.n504 B.n503 163.367
R589 B.n503 B.n502 163.367
R590 B.n502 B.n49 163.367
R591 B.n498 B.n49 163.367
R592 B.n498 B.n497 163.367
R593 B.n497 B.n496 163.367
R594 B.n496 B.n51 163.367
R595 B.n492 B.n51 163.367
R596 B.n492 B.n491 163.367
R597 B.n491 B.n490 163.367
R598 B.n490 B.n53 163.367
R599 B.n486 B.n53 163.367
R600 B.n486 B.n485 163.367
R601 B.n485 B.n484 163.367
R602 B.n484 B.n55 163.367
R603 B.n480 B.n55 163.367
R604 B.n480 B.n479 163.367
R605 B.n479 B.n478 163.367
R606 B.n478 B.n57 163.367
R607 B.n474 B.n57 163.367
R608 B.n474 B.n473 163.367
R609 B.n473 B.n472 163.367
R610 B.n472 B.n59 163.367
R611 B.n468 B.n59 163.367
R612 B.n468 B.n467 163.367
R613 B.n467 B.n466 163.367
R614 B.n466 B.n61 163.367
R615 B.n462 B.n61 163.367
R616 B.n462 B.n461 163.367
R617 B.n461 B.n460 163.367
R618 B.n460 B.n63 163.367
R619 B.n456 B.n63 163.367
R620 B.n456 B.n455 163.367
R621 B.n455 B.n454 163.367
R622 B.n454 B.n65 163.367
R623 B.n450 B.n65 163.367
R624 B.n450 B.n449 163.367
R625 B.n449 B.n448 163.367
R626 B.n448 B.n67 163.367
R627 B.n444 B.n67 163.367
R628 B.n444 B.n443 163.367
R629 B.n443 B.n442 163.367
R630 B.n442 B.n69 163.367
R631 B.n438 B.n69 163.367
R632 B.n438 B.n437 163.367
R633 B.n437 B.n436 163.367
R634 B.n436 B.n71 163.367
R635 B.n432 B.n71 163.367
R636 B.n432 B.n431 163.367
R637 B.n431 B.n430 163.367
R638 B.n430 B.n73 163.367
R639 B.n426 B.n73 163.367
R640 B.n426 B.n425 163.367
R641 B.n425 B.n424 163.367
R642 B.n424 B.n75 163.367
R643 B.n120 B.t2 132.489
R644 B.n46 B.t10 132.489
R645 B.n128 B.t5 132.468
R646 B.n38 B.t7 132.468
R647 B.n121 B.t1 106.501
R648 B.n47 B.t11 106.501
R649 B.n129 B.t4 106.48
R650 B.n39 B.t8 106.48
R651 B.n122 B.n121 59.5399
R652 B.n272 B.n129 59.5399
R653 B.n40 B.n39 59.5399
R654 B.n506 B.n47 59.5399
R655 B.n607 B.n10 34.4981
R656 B.n422 B.n421 34.4981
R657 B.n373 B.n92 34.4981
R658 B.n188 B.n187 34.4981
R659 B.n121 B.n120 25.9884
R660 B.n129 B.n128 25.9884
R661 B.n39 B.n38 25.9884
R662 B.n47 B.n46 25.9884
R663 B B.n631 18.0485
R664 B.n603 B.n10 10.6151
R665 B.n603 B.n602 10.6151
R666 B.n602 B.n601 10.6151
R667 B.n601 B.n12 10.6151
R668 B.n597 B.n12 10.6151
R669 B.n597 B.n596 10.6151
R670 B.n596 B.n595 10.6151
R671 B.n595 B.n14 10.6151
R672 B.n591 B.n14 10.6151
R673 B.n591 B.n590 10.6151
R674 B.n590 B.n589 10.6151
R675 B.n589 B.n16 10.6151
R676 B.n585 B.n16 10.6151
R677 B.n585 B.n584 10.6151
R678 B.n584 B.n583 10.6151
R679 B.n583 B.n18 10.6151
R680 B.n579 B.n18 10.6151
R681 B.n579 B.n578 10.6151
R682 B.n578 B.n577 10.6151
R683 B.n577 B.n20 10.6151
R684 B.n573 B.n20 10.6151
R685 B.n573 B.n572 10.6151
R686 B.n572 B.n571 10.6151
R687 B.n571 B.n22 10.6151
R688 B.n567 B.n22 10.6151
R689 B.n567 B.n566 10.6151
R690 B.n566 B.n565 10.6151
R691 B.n565 B.n24 10.6151
R692 B.n561 B.n24 10.6151
R693 B.n561 B.n560 10.6151
R694 B.n560 B.n559 10.6151
R695 B.n559 B.n26 10.6151
R696 B.n555 B.n26 10.6151
R697 B.n555 B.n554 10.6151
R698 B.n554 B.n553 10.6151
R699 B.n553 B.n28 10.6151
R700 B.n549 B.n28 10.6151
R701 B.n549 B.n548 10.6151
R702 B.n548 B.n547 10.6151
R703 B.n547 B.n30 10.6151
R704 B.n543 B.n30 10.6151
R705 B.n543 B.n542 10.6151
R706 B.n542 B.n541 10.6151
R707 B.n541 B.n32 10.6151
R708 B.n537 B.n32 10.6151
R709 B.n537 B.n536 10.6151
R710 B.n536 B.n535 10.6151
R711 B.n535 B.n34 10.6151
R712 B.n531 B.n34 10.6151
R713 B.n531 B.n530 10.6151
R714 B.n530 B.n529 10.6151
R715 B.n529 B.n36 10.6151
R716 B.n525 B.n36 10.6151
R717 B.n525 B.n524 10.6151
R718 B.n524 B.n523 10.6151
R719 B.n520 B.n519 10.6151
R720 B.n519 B.n518 10.6151
R721 B.n518 B.n42 10.6151
R722 B.n514 B.n42 10.6151
R723 B.n514 B.n513 10.6151
R724 B.n513 B.n512 10.6151
R725 B.n512 B.n44 10.6151
R726 B.n508 B.n44 10.6151
R727 B.n508 B.n507 10.6151
R728 B.n505 B.n48 10.6151
R729 B.n501 B.n48 10.6151
R730 B.n501 B.n500 10.6151
R731 B.n500 B.n499 10.6151
R732 B.n499 B.n50 10.6151
R733 B.n495 B.n50 10.6151
R734 B.n495 B.n494 10.6151
R735 B.n494 B.n493 10.6151
R736 B.n493 B.n52 10.6151
R737 B.n489 B.n52 10.6151
R738 B.n489 B.n488 10.6151
R739 B.n488 B.n487 10.6151
R740 B.n487 B.n54 10.6151
R741 B.n483 B.n54 10.6151
R742 B.n483 B.n482 10.6151
R743 B.n482 B.n481 10.6151
R744 B.n481 B.n56 10.6151
R745 B.n477 B.n56 10.6151
R746 B.n477 B.n476 10.6151
R747 B.n476 B.n475 10.6151
R748 B.n475 B.n58 10.6151
R749 B.n471 B.n58 10.6151
R750 B.n471 B.n470 10.6151
R751 B.n470 B.n469 10.6151
R752 B.n469 B.n60 10.6151
R753 B.n465 B.n60 10.6151
R754 B.n465 B.n464 10.6151
R755 B.n464 B.n463 10.6151
R756 B.n463 B.n62 10.6151
R757 B.n459 B.n62 10.6151
R758 B.n459 B.n458 10.6151
R759 B.n458 B.n457 10.6151
R760 B.n457 B.n64 10.6151
R761 B.n453 B.n64 10.6151
R762 B.n453 B.n452 10.6151
R763 B.n452 B.n451 10.6151
R764 B.n451 B.n66 10.6151
R765 B.n447 B.n66 10.6151
R766 B.n447 B.n446 10.6151
R767 B.n446 B.n445 10.6151
R768 B.n445 B.n68 10.6151
R769 B.n441 B.n68 10.6151
R770 B.n441 B.n440 10.6151
R771 B.n440 B.n439 10.6151
R772 B.n439 B.n70 10.6151
R773 B.n435 B.n70 10.6151
R774 B.n435 B.n434 10.6151
R775 B.n434 B.n433 10.6151
R776 B.n433 B.n72 10.6151
R777 B.n429 B.n72 10.6151
R778 B.n429 B.n428 10.6151
R779 B.n428 B.n427 10.6151
R780 B.n427 B.n74 10.6151
R781 B.n423 B.n74 10.6151
R782 B.n423 B.n422 10.6151
R783 B.n374 B.n373 10.6151
R784 B.n375 B.n374 10.6151
R785 B.n375 B.n90 10.6151
R786 B.n379 B.n90 10.6151
R787 B.n380 B.n379 10.6151
R788 B.n381 B.n380 10.6151
R789 B.n381 B.n88 10.6151
R790 B.n385 B.n88 10.6151
R791 B.n386 B.n385 10.6151
R792 B.n387 B.n386 10.6151
R793 B.n387 B.n86 10.6151
R794 B.n391 B.n86 10.6151
R795 B.n392 B.n391 10.6151
R796 B.n393 B.n392 10.6151
R797 B.n393 B.n84 10.6151
R798 B.n397 B.n84 10.6151
R799 B.n398 B.n397 10.6151
R800 B.n399 B.n398 10.6151
R801 B.n399 B.n82 10.6151
R802 B.n403 B.n82 10.6151
R803 B.n404 B.n403 10.6151
R804 B.n405 B.n404 10.6151
R805 B.n405 B.n80 10.6151
R806 B.n409 B.n80 10.6151
R807 B.n410 B.n409 10.6151
R808 B.n411 B.n410 10.6151
R809 B.n411 B.n78 10.6151
R810 B.n415 B.n78 10.6151
R811 B.n416 B.n415 10.6151
R812 B.n417 B.n416 10.6151
R813 B.n417 B.n76 10.6151
R814 B.n421 B.n76 10.6151
R815 B.n189 B.n188 10.6151
R816 B.n189 B.n156 10.6151
R817 B.n193 B.n156 10.6151
R818 B.n194 B.n193 10.6151
R819 B.n195 B.n194 10.6151
R820 B.n195 B.n154 10.6151
R821 B.n199 B.n154 10.6151
R822 B.n200 B.n199 10.6151
R823 B.n201 B.n200 10.6151
R824 B.n201 B.n152 10.6151
R825 B.n205 B.n152 10.6151
R826 B.n206 B.n205 10.6151
R827 B.n207 B.n206 10.6151
R828 B.n207 B.n150 10.6151
R829 B.n211 B.n150 10.6151
R830 B.n212 B.n211 10.6151
R831 B.n213 B.n212 10.6151
R832 B.n213 B.n148 10.6151
R833 B.n217 B.n148 10.6151
R834 B.n218 B.n217 10.6151
R835 B.n219 B.n218 10.6151
R836 B.n219 B.n146 10.6151
R837 B.n223 B.n146 10.6151
R838 B.n224 B.n223 10.6151
R839 B.n225 B.n224 10.6151
R840 B.n225 B.n144 10.6151
R841 B.n229 B.n144 10.6151
R842 B.n230 B.n229 10.6151
R843 B.n231 B.n230 10.6151
R844 B.n231 B.n142 10.6151
R845 B.n235 B.n142 10.6151
R846 B.n236 B.n235 10.6151
R847 B.n237 B.n236 10.6151
R848 B.n237 B.n140 10.6151
R849 B.n241 B.n140 10.6151
R850 B.n242 B.n241 10.6151
R851 B.n243 B.n242 10.6151
R852 B.n243 B.n138 10.6151
R853 B.n247 B.n138 10.6151
R854 B.n248 B.n247 10.6151
R855 B.n249 B.n248 10.6151
R856 B.n249 B.n136 10.6151
R857 B.n253 B.n136 10.6151
R858 B.n254 B.n253 10.6151
R859 B.n255 B.n254 10.6151
R860 B.n255 B.n134 10.6151
R861 B.n259 B.n134 10.6151
R862 B.n260 B.n259 10.6151
R863 B.n261 B.n260 10.6151
R864 B.n261 B.n132 10.6151
R865 B.n265 B.n132 10.6151
R866 B.n266 B.n265 10.6151
R867 B.n267 B.n266 10.6151
R868 B.n267 B.n130 10.6151
R869 B.n271 B.n130 10.6151
R870 B.n274 B.n273 10.6151
R871 B.n274 B.n126 10.6151
R872 B.n278 B.n126 10.6151
R873 B.n279 B.n278 10.6151
R874 B.n280 B.n279 10.6151
R875 B.n280 B.n124 10.6151
R876 B.n284 B.n124 10.6151
R877 B.n285 B.n284 10.6151
R878 B.n286 B.n285 10.6151
R879 B.n290 B.n289 10.6151
R880 B.n291 B.n290 10.6151
R881 B.n291 B.n118 10.6151
R882 B.n295 B.n118 10.6151
R883 B.n296 B.n295 10.6151
R884 B.n297 B.n296 10.6151
R885 B.n297 B.n116 10.6151
R886 B.n301 B.n116 10.6151
R887 B.n302 B.n301 10.6151
R888 B.n303 B.n302 10.6151
R889 B.n303 B.n114 10.6151
R890 B.n307 B.n114 10.6151
R891 B.n308 B.n307 10.6151
R892 B.n309 B.n308 10.6151
R893 B.n309 B.n112 10.6151
R894 B.n313 B.n112 10.6151
R895 B.n314 B.n313 10.6151
R896 B.n315 B.n314 10.6151
R897 B.n315 B.n110 10.6151
R898 B.n319 B.n110 10.6151
R899 B.n320 B.n319 10.6151
R900 B.n321 B.n320 10.6151
R901 B.n321 B.n108 10.6151
R902 B.n325 B.n108 10.6151
R903 B.n326 B.n325 10.6151
R904 B.n327 B.n326 10.6151
R905 B.n327 B.n106 10.6151
R906 B.n331 B.n106 10.6151
R907 B.n332 B.n331 10.6151
R908 B.n333 B.n332 10.6151
R909 B.n333 B.n104 10.6151
R910 B.n337 B.n104 10.6151
R911 B.n338 B.n337 10.6151
R912 B.n339 B.n338 10.6151
R913 B.n339 B.n102 10.6151
R914 B.n343 B.n102 10.6151
R915 B.n344 B.n343 10.6151
R916 B.n345 B.n344 10.6151
R917 B.n345 B.n100 10.6151
R918 B.n349 B.n100 10.6151
R919 B.n350 B.n349 10.6151
R920 B.n351 B.n350 10.6151
R921 B.n351 B.n98 10.6151
R922 B.n355 B.n98 10.6151
R923 B.n356 B.n355 10.6151
R924 B.n357 B.n356 10.6151
R925 B.n357 B.n96 10.6151
R926 B.n361 B.n96 10.6151
R927 B.n362 B.n361 10.6151
R928 B.n363 B.n362 10.6151
R929 B.n363 B.n94 10.6151
R930 B.n367 B.n94 10.6151
R931 B.n368 B.n367 10.6151
R932 B.n369 B.n368 10.6151
R933 B.n369 B.n92 10.6151
R934 B.n187 B.n158 10.6151
R935 B.n183 B.n158 10.6151
R936 B.n183 B.n182 10.6151
R937 B.n182 B.n181 10.6151
R938 B.n181 B.n160 10.6151
R939 B.n177 B.n160 10.6151
R940 B.n177 B.n176 10.6151
R941 B.n176 B.n175 10.6151
R942 B.n175 B.n162 10.6151
R943 B.n171 B.n162 10.6151
R944 B.n171 B.n170 10.6151
R945 B.n170 B.n169 10.6151
R946 B.n169 B.n164 10.6151
R947 B.n165 B.n164 10.6151
R948 B.n165 B.n0 10.6151
R949 B.n627 B.n1 10.6151
R950 B.n627 B.n626 10.6151
R951 B.n626 B.n625 10.6151
R952 B.n625 B.n4 10.6151
R953 B.n621 B.n4 10.6151
R954 B.n621 B.n620 10.6151
R955 B.n620 B.n619 10.6151
R956 B.n619 B.n6 10.6151
R957 B.n615 B.n6 10.6151
R958 B.n615 B.n614 10.6151
R959 B.n614 B.n613 10.6151
R960 B.n613 B.n8 10.6151
R961 B.n609 B.n8 10.6151
R962 B.n609 B.n608 10.6151
R963 B.n608 B.n607 10.6151
R964 B.n523 B.n40 8.74196
R965 B.n506 B.n505 8.74196
R966 B.n272 B.n271 8.74196
R967 B.n289 B.n122 8.74196
R968 B.n631 B.n0 2.81026
R969 B.n631 B.n1 2.81026
R970 B.n520 B.n40 1.87367
R971 B.n507 B.n506 1.87367
R972 B.n273 B.n272 1.87367
R973 B.n286 B.n122 1.87367
C0 w_n1506_n4374# VDD2 1.97724f
C1 VP VDD1 3.19514f
C2 B VTAIL 3.84128f
C3 VN VTAIL 2.40233f
C4 VDD1 VDD2 0.494323f
C5 VN B 0.839568f
C6 w_n1506_n4374# VTAIL 3.66659f
C7 VP VDD2 0.268563f
C8 B w_n1506_n4374# 8.50012f
C9 VDD1 VTAIL 6.94602f
C10 VN w_n1506_n4374# 2.0287f
C11 B VDD1 1.84221f
C12 VP VTAIL 2.41702f
C13 VN VDD1 0.14873f
C14 VTAIL VDD2 6.98067f
C15 B VP 1.14294f
C16 w_n1506_n4374# VDD1 1.96948f
C17 VN VP 5.62952f
C18 B VDD2 1.85893f
C19 VN VDD2 3.08071f
C20 VP w_n1506_n4374# 2.21711f
C21 VDD2 VSUBS 0.935122f
C22 VDD1 VSUBS 4.60897f
C23 VTAIL VSUBS 0.989685f
C24 VN VSUBS 8.62283f
C25 VP VSUBS 1.390829f
C26 B VSUBS 3.147035f
C27 w_n1506_n4374# VSUBS 80.6192f
C28 B.n0 VSUBS 0.004144f
C29 B.n1 VSUBS 0.004144f
C30 B.n2 VSUBS 0.006553f
C31 B.n3 VSUBS 0.006553f
C32 B.n4 VSUBS 0.006553f
C33 B.n5 VSUBS 0.006553f
C34 B.n6 VSUBS 0.006553f
C35 B.n7 VSUBS 0.006553f
C36 B.n8 VSUBS 0.006553f
C37 B.n9 VSUBS 0.006553f
C38 B.n10 VSUBS 0.016123f
C39 B.n11 VSUBS 0.006553f
C40 B.n12 VSUBS 0.006553f
C41 B.n13 VSUBS 0.006553f
C42 B.n14 VSUBS 0.006553f
C43 B.n15 VSUBS 0.006553f
C44 B.n16 VSUBS 0.006553f
C45 B.n17 VSUBS 0.006553f
C46 B.n18 VSUBS 0.006553f
C47 B.n19 VSUBS 0.006553f
C48 B.n20 VSUBS 0.006553f
C49 B.n21 VSUBS 0.006553f
C50 B.n22 VSUBS 0.006553f
C51 B.n23 VSUBS 0.006553f
C52 B.n24 VSUBS 0.006553f
C53 B.n25 VSUBS 0.006553f
C54 B.n26 VSUBS 0.006553f
C55 B.n27 VSUBS 0.006553f
C56 B.n28 VSUBS 0.006553f
C57 B.n29 VSUBS 0.006553f
C58 B.n30 VSUBS 0.006553f
C59 B.n31 VSUBS 0.006553f
C60 B.n32 VSUBS 0.006553f
C61 B.n33 VSUBS 0.006553f
C62 B.n34 VSUBS 0.006553f
C63 B.n35 VSUBS 0.006553f
C64 B.n36 VSUBS 0.006553f
C65 B.n37 VSUBS 0.006553f
C66 B.t8 VSUBS 0.535333f
C67 B.t7 VSUBS 0.545535f
C68 B.t6 VSUBS 0.66631f
C69 B.n38 VSUBS 0.198576f
C70 B.n39 VSUBS 0.061345f
C71 B.n40 VSUBS 0.015182f
C72 B.n41 VSUBS 0.006553f
C73 B.n42 VSUBS 0.006553f
C74 B.n43 VSUBS 0.006553f
C75 B.n44 VSUBS 0.006553f
C76 B.n45 VSUBS 0.006553f
C77 B.t11 VSUBS 0.535315f
C78 B.t10 VSUBS 0.545518f
C79 B.t9 VSUBS 0.66631f
C80 B.n46 VSUBS 0.198593f
C81 B.n47 VSUBS 0.061363f
C82 B.n48 VSUBS 0.006553f
C83 B.n49 VSUBS 0.006553f
C84 B.n50 VSUBS 0.006553f
C85 B.n51 VSUBS 0.006553f
C86 B.n52 VSUBS 0.006553f
C87 B.n53 VSUBS 0.006553f
C88 B.n54 VSUBS 0.006553f
C89 B.n55 VSUBS 0.006553f
C90 B.n56 VSUBS 0.006553f
C91 B.n57 VSUBS 0.006553f
C92 B.n58 VSUBS 0.006553f
C93 B.n59 VSUBS 0.006553f
C94 B.n60 VSUBS 0.006553f
C95 B.n61 VSUBS 0.006553f
C96 B.n62 VSUBS 0.006553f
C97 B.n63 VSUBS 0.006553f
C98 B.n64 VSUBS 0.006553f
C99 B.n65 VSUBS 0.006553f
C100 B.n66 VSUBS 0.006553f
C101 B.n67 VSUBS 0.006553f
C102 B.n68 VSUBS 0.006553f
C103 B.n69 VSUBS 0.006553f
C104 B.n70 VSUBS 0.006553f
C105 B.n71 VSUBS 0.006553f
C106 B.n72 VSUBS 0.006553f
C107 B.n73 VSUBS 0.006553f
C108 B.n74 VSUBS 0.006553f
C109 B.n75 VSUBS 0.016123f
C110 B.n76 VSUBS 0.006553f
C111 B.n77 VSUBS 0.006553f
C112 B.n78 VSUBS 0.006553f
C113 B.n79 VSUBS 0.006553f
C114 B.n80 VSUBS 0.006553f
C115 B.n81 VSUBS 0.006553f
C116 B.n82 VSUBS 0.006553f
C117 B.n83 VSUBS 0.006553f
C118 B.n84 VSUBS 0.006553f
C119 B.n85 VSUBS 0.006553f
C120 B.n86 VSUBS 0.006553f
C121 B.n87 VSUBS 0.006553f
C122 B.n88 VSUBS 0.006553f
C123 B.n89 VSUBS 0.006553f
C124 B.n90 VSUBS 0.006553f
C125 B.n91 VSUBS 0.006553f
C126 B.n92 VSUBS 0.016123f
C127 B.n93 VSUBS 0.006553f
C128 B.n94 VSUBS 0.006553f
C129 B.n95 VSUBS 0.006553f
C130 B.n96 VSUBS 0.006553f
C131 B.n97 VSUBS 0.006553f
C132 B.n98 VSUBS 0.006553f
C133 B.n99 VSUBS 0.006553f
C134 B.n100 VSUBS 0.006553f
C135 B.n101 VSUBS 0.006553f
C136 B.n102 VSUBS 0.006553f
C137 B.n103 VSUBS 0.006553f
C138 B.n104 VSUBS 0.006553f
C139 B.n105 VSUBS 0.006553f
C140 B.n106 VSUBS 0.006553f
C141 B.n107 VSUBS 0.006553f
C142 B.n108 VSUBS 0.006553f
C143 B.n109 VSUBS 0.006553f
C144 B.n110 VSUBS 0.006553f
C145 B.n111 VSUBS 0.006553f
C146 B.n112 VSUBS 0.006553f
C147 B.n113 VSUBS 0.006553f
C148 B.n114 VSUBS 0.006553f
C149 B.n115 VSUBS 0.006553f
C150 B.n116 VSUBS 0.006553f
C151 B.n117 VSUBS 0.006553f
C152 B.n118 VSUBS 0.006553f
C153 B.n119 VSUBS 0.006553f
C154 B.t1 VSUBS 0.535315f
C155 B.t2 VSUBS 0.545518f
C156 B.t0 VSUBS 0.66631f
C157 B.n120 VSUBS 0.198593f
C158 B.n121 VSUBS 0.061363f
C159 B.n122 VSUBS 0.015182f
C160 B.n123 VSUBS 0.006553f
C161 B.n124 VSUBS 0.006553f
C162 B.n125 VSUBS 0.006553f
C163 B.n126 VSUBS 0.006553f
C164 B.n127 VSUBS 0.006553f
C165 B.t4 VSUBS 0.535333f
C166 B.t5 VSUBS 0.545535f
C167 B.t3 VSUBS 0.66631f
C168 B.n128 VSUBS 0.198576f
C169 B.n129 VSUBS 0.061345f
C170 B.n130 VSUBS 0.006553f
C171 B.n131 VSUBS 0.006553f
C172 B.n132 VSUBS 0.006553f
C173 B.n133 VSUBS 0.006553f
C174 B.n134 VSUBS 0.006553f
C175 B.n135 VSUBS 0.006553f
C176 B.n136 VSUBS 0.006553f
C177 B.n137 VSUBS 0.006553f
C178 B.n138 VSUBS 0.006553f
C179 B.n139 VSUBS 0.006553f
C180 B.n140 VSUBS 0.006553f
C181 B.n141 VSUBS 0.006553f
C182 B.n142 VSUBS 0.006553f
C183 B.n143 VSUBS 0.006553f
C184 B.n144 VSUBS 0.006553f
C185 B.n145 VSUBS 0.006553f
C186 B.n146 VSUBS 0.006553f
C187 B.n147 VSUBS 0.006553f
C188 B.n148 VSUBS 0.006553f
C189 B.n149 VSUBS 0.006553f
C190 B.n150 VSUBS 0.006553f
C191 B.n151 VSUBS 0.006553f
C192 B.n152 VSUBS 0.006553f
C193 B.n153 VSUBS 0.006553f
C194 B.n154 VSUBS 0.006553f
C195 B.n155 VSUBS 0.006553f
C196 B.n156 VSUBS 0.006553f
C197 B.n157 VSUBS 0.016123f
C198 B.n158 VSUBS 0.006553f
C199 B.n159 VSUBS 0.006553f
C200 B.n160 VSUBS 0.006553f
C201 B.n161 VSUBS 0.006553f
C202 B.n162 VSUBS 0.006553f
C203 B.n163 VSUBS 0.006553f
C204 B.n164 VSUBS 0.006553f
C205 B.n165 VSUBS 0.006553f
C206 B.n166 VSUBS 0.006553f
C207 B.n167 VSUBS 0.006553f
C208 B.n168 VSUBS 0.006553f
C209 B.n169 VSUBS 0.006553f
C210 B.n170 VSUBS 0.006553f
C211 B.n171 VSUBS 0.006553f
C212 B.n172 VSUBS 0.006553f
C213 B.n173 VSUBS 0.006553f
C214 B.n174 VSUBS 0.006553f
C215 B.n175 VSUBS 0.006553f
C216 B.n176 VSUBS 0.006553f
C217 B.n177 VSUBS 0.006553f
C218 B.n178 VSUBS 0.006553f
C219 B.n179 VSUBS 0.006553f
C220 B.n180 VSUBS 0.006553f
C221 B.n181 VSUBS 0.006553f
C222 B.n182 VSUBS 0.006553f
C223 B.n183 VSUBS 0.006553f
C224 B.n184 VSUBS 0.006553f
C225 B.n185 VSUBS 0.006553f
C226 B.n186 VSUBS 0.015677f
C227 B.n187 VSUBS 0.015677f
C228 B.n188 VSUBS 0.016123f
C229 B.n189 VSUBS 0.006553f
C230 B.n190 VSUBS 0.006553f
C231 B.n191 VSUBS 0.006553f
C232 B.n192 VSUBS 0.006553f
C233 B.n193 VSUBS 0.006553f
C234 B.n194 VSUBS 0.006553f
C235 B.n195 VSUBS 0.006553f
C236 B.n196 VSUBS 0.006553f
C237 B.n197 VSUBS 0.006553f
C238 B.n198 VSUBS 0.006553f
C239 B.n199 VSUBS 0.006553f
C240 B.n200 VSUBS 0.006553f
C241 B.n201 VSUBS 0.006553f
C242 B.n202 VSUBS 0.006553f
C243 B.n203 VSUBS 0.006553f
C244 B.n204 VSUBS 0.006553f
C245 B.n205 VSUBS 0.006553f
C246 B.n206 VSUBS 0.006553f
C247 B.n207 VSUBS 0.006553f
C248 B.n208 VSUBS 0.006553f
C249 B.n209 VSUBS 0.006553f
C250 B.n210 VSUBS 0.006553f
C251 B.n211 VSUBS 0.006553f
C252 B.n212 VSUBS 0.006553f
C253 B.n213 VSUBS 0.006553f
C254 B.n214 VSUBS 0.006553f
C255 B.n215 VSUBS 0.006553f
C256 B.n216 VSUBS 0.006553f
C257 B.n217 VSUBS 0.006553f
C258 B.n218 VSUBS 0.006553f
C259 B.n219 VSUBS 0.006553f
C260 B.n220 VSUBS 0.006553f
C261 B.n221 VSUBS 0.006553f
C262 B.n222 VSUBS 0.006553f
C263 B.n223 VSUBS 0.006553f
C264 B.n224 VSUBS 0.006553f
C265 B.n225 VSUBS 0.006553f
C266 B.n226 VSUBS 0.006553f
C267 B.n227 VSUBS 0.006553f
C268 B.n228 VSUBS 0.006553f
C269 B.n229 VSUBS 0.006553f
C270 B.n230 VSUBS 0.006553f
C271 B.n231 VSUBS 0.006553f
C272 B.n232 VSUBS 0.006553f
C273 B.n233 VSUBS 0.006553f
C274 B.n234 VSUBS 0.006553f
C275 B.n235 VSUBS 0.006553f
C276 B.n236 VSUBS 0.006553f
C277 B.n237 VSUBS 0.006553f
C278 B.n238 VSUBS 0.006553f
C279 B.n239 VSUBS 0.006553f
C280 B.n240 VSUBS 0.006553f
C281 B.n241 VSUBS 0.006553f
C282 B.n242 VSUBS 0.006553f
C283 B.n243 VSUBS 0.006553f
C284 B.n244 VSUBS 0.006553f
C285 B.n245 VSUBS 0.006553f
C286 B.n246 VSUBS 0.006553f
C287 B.n247 VSUBS 0.006553f
C288 B.n248 VSUBS 0.006553f
C289 B.n249 VSUBS 0.006553f
C290 B.n250 VSUBS 0.006553f
C291 B.n251 VSUBS 0.006553f
C292 B.n252 VSUBS 0.006553f
C293 B.n253 VSUBS 0.006553f
C294 B.n254 VSUBS 0.006553f
C295 B.n255 VSUBS 0.006553f
C296 B.n256 VSUBS 0.006553f
C297 B.n257 VSUBS 0.006553f
C298 B.n258 VSUBS 0.006553f
C299 B.n259 VSUBS 0.006553f
C300 B.n260 VSUBS 0.006553f
C301 B.n261 VSUBS 0.006553f
C302 B.n262 VSUBS 0.006553f
C303 B.n263 VSUBS 0.006553f
C304 B.n264 VSUBS 0.006553f
C305 B.n265 VSUBS 0.006553f
C306 B.n266 VSUBS 0.006553f
C307 B.n267 VSUBS 0.006553f
C308 B.n268 VSUBS 0.006553f
C309 B.n269 VSUBS 0.006553f
C310 B.n270 VSUBS 0.006553f
C311 B.n271 VSUBS 0.005975f
C312 B.n272 VSUBS 0.015182f
C313 B.n273 VSUBS 0.003855f
C314 B.n274 VSUBS 0.006553f
C315 B.n275 VSUBS 0.006553f
C316 B.n276 VSUBS 0.006553f
C317 B.n277 VSUBS 0.006553f
C318 B.n278 VSUBS 0.006553f
C319 B.n279 VSUBS 0.006553f
C320 B.n280 VSUBS 0.006553f
C321 B.n281 VSUBS 0.006553f
C322 B.n282 VSUBS 0.006553f
C323 B.n283 VSUBS 0.006553f
C324 B.n284 VSUBS 0.006553f
C325 B.n285 VSUBS 0.006553f
C326 B.n286 VSUBS 0.003855f
C327 B.n287 VSUBS 0.006553f
C328 B.n288 VSUBS 0.006553f
C329 B.n289 VSUBS 0.005975f
C330 B.n290 VSUBS 0.006553f
C331 B.n291 VSUBS 0.006553f
C332 B.n292 VSUBS 0.006553f
C333 B.n293 VSUBS 0.006553f
C334 B.n294 VSUBS 0.006553f
C335 B.n295 VSUBS 0.006553f
C336 B.n296 VSUBS 0.006553f
C337 B.n297 VSUBS 0.006553f
C338 B.n298 VSUBS 0.006553f
C339 B.n299 VSUBS 0.006553f
C340 B.n300 VSUBS 0.006553f
C341 B.n301 VSUBS 0.006553f
C342 B.n302 VSUBS 0.006553f
C343 B.n303 VSUBS 0.006553f
C344 B.n304 VSUBS 0.006553f
C345 B.n305 VSUBS 0.006553f
C346 B.n306 VSUBS 0.006553f
C347 B.n307 VSUBS 0.006553f
C348 B.n308 VSUBS 0.006553f
C349 B.n309 VSUBS 0.006553f
C350 B.n310 VSUBS 0.006553f
C351 B.n311 VSUBS 0.006553f
C352 B.n312 VSUBS 0.006553f
C353 B.n313 VSUBS 0.006553f
C354 B.n314 VSUBS 0.006553f
C355 B.n315 VSUBS 0.006553f
C356 B.n316 VSUBS 0.006553f
C357 B.n317 VSUBS 0.006553f
C358 B.n318 VSUBS 0.006553f
C359 B.n319 VSUBS 0.006553f
C360 B.n320 VSUBS 0.006553f
C361 B.n321 VSUBS 0.006553f
C362 B.n322 VSUBS 0.006553f
C363 B.n323 VSUBS 0.006553f
C364 B.n324 VSUBS 0.006553f
C365 B.n325 VSUBS 0.006553f
C366 B.n326 VSUBS 0.006553f
C367 B.n327 VSUBS 0.006553f
C368 B.n328 VSUBS 0.006553f
C369 B.n329 VSUBS 0.006553f
C370 B.n330 VSUBS 0.006553f
C371 B.n331 VSUBS 0.006553f
C372 B.n332 VSUBS 0.006553f
C373 B.n333 VSUBS 0.006553f
C374 B.n334 VSUBS 0.006553f
C375 B.n335 VSUBS 0.006553f
C376 B.n336 VSUBS 0.006553f
C377 B.n337 VSUBS 0.006553f
C378 B.n338 VSUBS 0.006553f
C379 B.n339 VSUBS 0.006553f
C380 B.n340 VSUBS 0.006553f
C381 B.n341 VSUBS 0.006553f
C382 B.n342 VSUBS 0.006553f
C383 B.n343 VSUBS 0.006553f
C384 B.n344 VSUBS 0.006553f
C385 B.n345 VSUBS 0.006553f
C386 B.n346 VSUBS 0.006553f
C387 B.n347 VSUBS 0.006553f
C388 B.n348 VSUBS 0.006553f
C389 B.n349 VSUBS 0.006553f
C390 B.n350 VSUBS 0.006553f
C391 B.n351 VSUBS 0.006553f
C392 B.n352 VSUBS 0.006553f
C393 B.n353 VSUBS 0.006553f
C394 B.n354 VSUBS 0.006553f
C395 B.n355 VSUBS 0.006553f
C396 B.n356 VSUBS 0.006553f
C397 B.n357 VSUBS 0.006553f
C398 B.n358 VSUBS 0.006553f
C399 B.n359 VSUBS 0.006553f
C400 B.n360 VSUBS 0.006553f
C401 B.n361 VSUBS 0.006553f
C402 B.n362 VSUBS 0.006553f
C403 B.n363 VSUBS 0.006553f
C404 B.n364 VSUBS 0.006553f
C405 B.n365 VSUBS 0.006553f
C406 B.n366 VSUBS 0.006553f
C407 B.n367 VSUBS 0.006553f
C408 B.n368 VSUBS 0.006553f
C409 B.n369 VSUBS 0.006553f
C410 B.n370 VSUBS 0.006553f
C411 B.n371 VSUBS 0.016123f
C412 B.n372 VSUBS 0.015677f
C413 B.n373 VSUBS 0.015677f
C414 B.n374 VSUBS 0.006553f
C415 B.n375 VSUBS 0.006553f
C416 B.n376 VSUBS 0.006553f
C417 B.n377 VSUBS 0.006553f
C418 B.n378 VSUBS 0.006553f
C419 B.n379 VSUBS 0.006553f
C420 B.n380 VSUBS 0.006553f
C421 B.n381 VSUBS 0.006553f
C422 B.n382 VSUBS 0.006553f
C423 B.n383 VSUBS 0.006553f
C424 B.n384 VSUBS 0.006553f
C425 B.n385 VSUBS 0.006553f
C426 B.n386 VSUBS 0.006553f
C427 B.n387 VSUBS 0.006553f
C428 B.n388 VSUBS 0.006553f
C429 B.n389 VSUBS 0.006553f
C430 B.n390 VSUBS 0.006553f
C431 B.n391 VSUBS 0.006553f
C432 B.n392 VSUBS 0.006553f
C433 B.n393 VSUBS 0.006553f
C434 B.n394 VSUBS 0.006553f
C435 B.n395 VSUBS 0.006553f
C436 B.n396 VSUBS 0.006553f
C437 B.n397 VSUBS 0.006553f
C438 B.n398 VSUBS 0.006553f
C439 B.n399 VSUBS 0.006553f
C440 B.n400 VSUBS 0.006553f
C441 B.n401 VSUBS 0.006553f
C442 B.n402 VSUBS 0.006553f
C443 B.n403 VSUBS 0.006553f
C444 B.n404 VSUBS 0.006553f
C445 B.n405 VSUBS 0.006553f
C446 B.n406 VSUBS 0.006553f
C447 B.n407 VSUBS 0.006553f
C448 B.n408 VSUBS 0.006553f
C449 B.n409 VSUBS 0.006553f
C450 B.n410 VSUBS 0.006553f
C451 B.n411 VSUBS 0.006553f
C452 B.n412 VSUBS 0.006553f
C453 B.n413 VSUBS 0.006553f
C454 B.n414 VSUBS 0.006553f
C455 B.n415 VSUBS 0.006553f
C456 B.n416 VSUBS 0.006553f
C457 B.n417 VSUBS 0.006553f
C458 B.n418 VSUBS 0.006553f
C459 B.n419 VSUBS 0.006553f
C460 B.n420 VSUBS 0.015677f
C461 B.n421 VSUBS 0.016409f
C462 B.n422 VSUBS 0.01539f
C463 B.n423 VSUBS 0.006553f
C464 B.n424 VSUBS 0.006553f
C465 B.n425 VSUBS 0.006553f
C466 B.n426 VSUBS 0.006553f
C467 B.n427 VSUBS 0.006553f
C468 B.n428 VSUBS 0.006553f
C469 B.n429 VSUBS 0.006553f
C470 B.n430 VSUBS 0.006553f
C471 B.n431 VSUBS 0.006553f
C472 B.n432 VSUBS 0.006553f
C473 B.n433 VSUBS 0.006553f
C474 B.n434 VSUBS 0.006553f
C475 B.n435 VSUBS 0.006553f
C476 B.n436 VSUBS 0.006553f
C477 B.n437 VSUBS 0.006553f
C478 B.n438 VSUBS 0.006553f
C479 B.n439 VSUBS 0.006553f
C480 B.n440 VSUBS 0.006553f
C481 B.n441 VSUBS 0.006553f
C482 B.n442 VSUBS 0.006553f
C483 B.n443 VSUBS 0.006553f
C484 B.n444 VSUBS 0.006553f
C485 B.n445 VSUBS 0.006553f
C486 B.n446 VSUBS 0.006553f
C487 B.n447 VSUBS 0.006553f
C488 B.n448 VSUBS 0.006553f
C489 B.n449 VSUBS 0.006553f
C490 B.n450 VSUBS 0.006553f
C491 B.n451 VSUBS 0.006553f
C492 B.n452 VSUBS 0.006553f
C493 B.n453 VSUBS 0.006553f
C494 B.n454 VSUBS 0.006553f
C495 B.n455 VSUBS 0.006553f
C496 B.n456 VSUBS 0.006553f
C497 B.n457 VSUBS 0.006553f
C498 B.n458 VSUBS 0.006553f
C499 B.n459 VSUBS 0.006553f
C500 B.n460 VSUBS 0.006553f
C501 B.n461 VSUBS 0.006553f
C502 B.n462 VSUBS 0.006553f
C503 B.n463 VSUBS 0.006553f
C504 B.n464 VSUBS 0.006553f
C505 B.n465 VSUBS 0.006553f
C506 B.n466 VSUBS 0.006553f
C507 B.n467 VSUBS 0.006553f
C508 B.n468 VSUBS 0.006553f
C509 B.n469 VSUBS 0.006553f
C510 B.n470 VSUBS 0.006553f
C511 B.n471 VSUBS 0.006553f
C512 B.n472 VSUBS 0.006553f
C513 B.n473 VSUBS 0.006553f
C514 B.n474 VSUBS 0.006553f
C515 B.n475 VSUBS 0.006553f
C516 B.n476 VSUBS 0.006553f
C517 B.n477 VSUBS 0.006553f
C518 B.n478 VSUBS 0.006553f
C519 B.n479 VSUBS 0.006553f
C520 B.n480 VSUBS 0.006553f
C521 B.n481 VSUBS 0.006553f
C522 B.n482 VSUBS 0.006553f
C523 B.n483 VSUBS 0.006553f
C524 B.n484 VSUBS 0.006553f
C525 B.n485 VSUBS 0.006553f
C526 B.n486 VSUBS 0.006553f
C527 B.n487 VSUBS 0.006553f
C528 B.n488 VSUBS 0.006553f
C529 B.n489 VSUBS 0.006553f
C530 B.n490 VSUBS 0.006553f
C531 B.n491 VSUBS 0.006553f
C532 B.n492 VSUBS 0.006553f
C533 B.n493 VSUBS 0.006553f
C534 B.n494 VSUBS 0.006553f
C535 B.n495 VSUBS 0.006553f
C536 B.n496 VSUBS 0.006553f
C537 B.n497 VSUBS 0.006553f
C538 B.n498 VSUBS 0.006553f
C539 B.n499 VSUBS 0.006553f
C540 B.n500 VSUBS 0.006553f
C541 B.n501 VSUBS 0.006553f
C542 B.n502 VSUBS 0.006553f
C543 B.n503 VSUBS 0.006553f
C544 B.n504 VSUBS 0.006553f
C545 B.n505 VSUBS 0.005975f
C546 B.n506 VSUBS 0.015182f
C547 B.n507 VSUBS 0.003855f
C548 B.n508 VSUBS 0.006553f
C549 B.n509 VSUBS 0.006553f
C550 B.n510 VSUBS 0.006553f
C551 B.n511 VSUBS 0.006553f
C552 B.n512 VSUBS 0.006553f
C553 B.n513 VSUBS 0.006553f
C554 B.n514 VSUBS 0.006553f
C555 B.n515 VSUBS 0.006553f
C556 B.n516 VSUBS 0.006553f
C557 B.n517 VSUBS 0.006553f
C558 B.n518 VSUBS 0.006553f
C559 B.n519 VSUBS 0.006553f
C560 B.n520 VSUBS 0.003855f
C561 B.n521 VSUBS 0.006553f
C562 B.n522 VSUBS 0.006553f
C563 B.n523 VSUBS 0.005975f
C564 B.n524 VSUBS 0.006553f
C565 B.n525 VSUBS 0.006553f
C566 B.n526 VSUBS 0.006553f
C567 B.n527 VSUBS 0.006553f
C568 B.n528 VSUBS 0.006553f
C569 B.n529 VSUBS 0.006553f
C570 B.n530 VSUBS 0.006553f
C571 B.n531 VSUBS 0.006553f
C572 B.n532 VSUBS 0.006553f
C573 B.n533 VSUBS 0.006553f
C574 B.n534 VSUBS 0.006553f
C575 B.n535 VSUBS 0.006553f
C576 B.n536 VSUBS 0.006553f
C577 B.n537 VSUBS 0.006553f
C578 B.n538 VSUBS 0.006553f
C579 B.n539 VSUBS 0.006553f
C580 B.n540 VSUBS 0.006553f
C581 B.n541 VSUBS 0.006553f
C582 B.n542 VSUBS 0.006553f
C583 B.n543 VSUBS 0.006553f
C584 B.n544 VSUBS 0.006553f
C585 B.n545 VSUBS 0.006553f
C586 B.n546 VSUBS 0.006553f
C587 B.n547 VSUBS 0.006553f
C588 B.n548 VSUBS 0.006553f
C589 B.n549 VSUBS 0.006553f
C590 B.n550 VSUBS 0.006553f
C591 B.n551 VSUBS 0.006553f
C592 B.n552 VSUBS 0.006553f
C593 B.n553 VSUBS 0.006553f
C594 B.n554 VSUBS 0.006553f
C595 B.n555 VSUBS 0.006553f
C596 B.n556 VSUBS 0.006553f
C597 B.n557 VSUBS 0.006553f
C598 B.n558 VSUBS 0.006553f
C599 B.n559 VSUBS 0.006553f
C600 B.n560 VSUBS 0.006553f
C601 B.n561 VSUBS 0.006553f
C602 B.n562 VSUBS 0.006553f
C603 B.n563 VSUBS 0.006553f
C604 B.n564 VSUBS 0.006553f
C605 B.n565 VSUBS 0.006553f
C606 B.n566 VSUBS 0.006553f
C607 B.n567 VSUBS 0.006553f
C608 B.n568 VSUBS 0.006553f
C609 B.n569 VSUBS 0.006553f
C610 B.n570 VSUBS 0.006553f
C611 B.n571 VSUBS 0.006553f
C612 B.n572 VSUBS 0.006553f
C613 B.n573 VSUBS 0.006553f
C614 B.n574 VSUBS 0.006553f
C615 B.n575 VSUBS 0.006553f
C616 B.n576 VSUBS 0.006553f
C617 B.n577 VSUBS 0.006553f
C618 B.n578 VSUBS 0.006553f
C619 B.n579 VSUBS 0.006553f
C620 B.n580 VSUBS 0.006553f
C621 B.n581 VSUBS 0.006553f
C622 B.n582 VSUBS 0.006553f
C623 B.n583 VSUBS 0.006553f
C624 B.n584 VSUBS 0.006553f
C625 B.n585 VSUBS 0.006553f
C626 B.n586 VSUBS 0.006553f
C627 B.n587 VSUBS 0.006553f
C628 B.n588 VSUBS 0.006553f
C629 B.n589 VSUBS 0.006553f
C630 B.n590 VSUBS 0.006553f
C631 B.n591 VSUBS 0.006553f
C632 B.n592 VSUBS 0.006553f
C633 B.n593 VSUBS 0.006553f
C634 B.n594 VSUBS 0.006553f
C635 B.n595 VSUBS 0.006553f
C636 B.n596 VSUBS 0.006553f
C637 B.n597 VSUBS 0.006553f
C638 B.n598 VSUBS 0.006553f
C639 B.n599 VSUBS 0.006553f
C640 B.n600 VSUBS 0.006553f
C641 B.n601 VSUBS 0.006553f
C642 B.n602 VSUBS 0.006553f
C643 B.n603 VSUBS 0.006553f
C644 B.n604 VSUBS 0.006553f
C645 B.n605 VSUBS 0.016123f
C646 B.n606 VSUBS 0.015677f
C647 B.n607 VSUBS 0.015677f
C648 B.n608 VSUBS 0.006553f
C649 B.n609 VSUBS 0.006553f
C650 B.n610 VSUBS 0.006553f
C651 B.n611 VSUBS 0.006553f
C652 B.n612 VSUBS 0.006553f
C653 B.n613 VSUBS 0.006553f
C654 B.n614 VSUBS 0.006553f
C655 B.n615 VSUBS 0.006553f
C656 B.n616 VSUBS 0.006553f
C657 B.n617 VSUBS 0.006553f
C658 B.n618 VSUBS 0.006553f
C659 B.n619 VSUBS 0.006553f
C660 B.n620 VSUBS 0.006553f
C661 B.n621 VSUBS 0.006553f
C662 B.n622 VSUBS 0.006553f
C663 B.n623 VSUBS 0.006553f
C664 B.n624 VSUBS 0.006553f
C665 B.n625 VSUBS 0.006553f
C666 B.n626 VSUBS 0.006553f
C667 B.n627 VSUBS 0.006553f
C668 B.n628 VSUBS 0.006553f
C669 B.n629 VSUBS 0.006553f
C670 B.n630 VSUBS 0.006553f
C671 B.n631 VSUBS 0.014838f
C672 VDD1.t1 VSUBS 2.94214f
C673 VDD1.t0 VSUBS 3.58815f
C674 VP.t0 VSUBS 3.42468f
C675 VP.t1 VSUBS 3.18743f
C676 VP.n0 VSUBS 6.75581f
C677 VDD2.t1 VSUBS 3.58755f
C678 VDD2.t0 VSUBS 2.96188f
C679 VDD2.n0 VSUBS 3.4892f
C680 VTAIL.t0 VSUBS 3.86042f
C681 VTAIL.n0 VSUBS 2.72066f
C682 VTAIL.t3 VSUBS 3.86042f
C683 VTAIL.n1 VSUBS 2.74132f
C684 VTAIL.t1 VSUBS 3.86041f
C685 VTAIL.n2 VSUBS 2.63785f
C686 VTAIL.t2 VSUBS 3.86042f
C687 VTAIL.n3 VSUBS 2.56466f
C688 VN.t0 VSUBS 3.09682f
C689 VN.t1 VSUBS 3.33169f
.ends

