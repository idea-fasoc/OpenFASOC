* NGSPICE file created from diff_pair_sample_0728.ext - technology: sky130A

.subckt diff_pair_sample_0728 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t3 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X1 VDD1.t2 VP.t1 VTAIL.t18 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X2 VDD1.t6 VP.t2 VTAIL.t17 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0.77385 ps=5.02 w=4.69 l=3.16
X3 VDD1.t4 VP.t3 VTAIL.t16 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=1.8291 ps=10.16 w=4.69 l=3.16
X4 B.t11 B.t9 B.t10 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0 ps=0 w=4.69 l=3.16
X5 B.t8 B.t6 B.t7 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0 ps=0 w=4.69 l=3.16
X6 VDD2.t9 VN.t0 VTAIL.t2 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=1.8291 ps=10.16 w=4.69 l=3.16
X7 VDD2.t8 VN.t1 VTAIL.t8 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=1.8291 ps=10.16 w=4.69 l=3.16
X8 VTAIL.t6 VN.t2 VDD2.t7 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X9 VTAIL.t15 VP.t4 VDD1.t0 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X10 VDD2.t6 VN.t3 VTAIL.t7 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0.77385 ps=5.02 w=4.69 l=3.16
X11 VTAIL.t4 VN.t4 VDD2.t5 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X12 VDD2.t4 VN.t5 VTAIL.t9 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0.77385 ps=5.02 w=4.69 l=3.16
X13 VDD2.t3 VN.t6 VTAIL.t5 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X14 VTAIL.t14 VP.t5 VDD1.t7 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X15 B.t5 B.t3 B.t4 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0 ps=0 w=4.69 l=3.16
X16 VDD2.t2 VN.t7 VTAIL.t3 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X17 B.t2 B.t0 B.t1 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0 ps=0 w=4.69 l=3.16
X18 VDD1.t9 VP.t6 VTAIL.t13 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=1.8291 ps=10.16 w=4.69 l=3.16
X19 VDD1.t8 VP.t7 VTAIL.t12 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=1.8291 pd=10.16 as=0.77385 ps=5.02 w=4.69 l=3.16
X20 VDD1.t5 VP.t8 VTAIL.t11 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X21 VTAIL.t0 VN.t8 VDD2.t1 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X22 VTAIL.t10 VP.t9 VDD1.t1 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
X23 VTAIL.t1 VN.t9 VDD2.t0 w_n5158_n1906# sky130_fd_pr__pfet_01v8 ad=0.77385 pd=5.02 as=0.77385 ps=5.02 w=4.69 l=3.16
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n20 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n19 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n18 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n109 VP.n108 161.3
R22 VP.n107 VP.n1 161.3
R23 VP.n106 VP.n105 161.3
R24 VP.n104 VP.n2 161.3
R25 VP.n103 VP.n102 161.3
R26 VP.n101 VP.n3 161.3
R27 VP.n100 VP.n99 161.3
R28 VP.n98 VP.n97 161.3
R29 VP.n96 VP.n5 161.3
R30 VP.n95 VP.n94 161.3
R31 VP.n93 VP.n6 161.3
R32 VP.n92 VP.n91 161.3
R33 VP.n90 VP.n7 161.3
R34 VP.n89 VP.n88 161.3
R35 VP.n87 VP.n86 161.3
R36 VP.n85 VP.n9 161.3
R37 VP.n84 VP.n83 161.3
R38 VP.n82 VP.n10 161.3
R39 VP.n81 VP.n80 161.3
R40 VP.n79 VP.n11 161.3
R41 VP.n78 VP.n77 161.3
R42 VP.n76 VP.n75 161.3
R43 VP.n74 VP.n13 161.3
R44 VP.n73 VP.n72 161.3
R45 VP.n71 VP.n14 161.3
R46 VP.n70 VP.n69 161.3
R47 VP.n68 VP.n15 161.3
R48 VP.n67 VP.n66 161.3
R49 VP.n65 VP.n16 78.8126
R50 VP.n110 VP.n0 78.8126
R51 VP.n64 VP.n17 78.8126
R52 VP.n30 VP.t2 68.2467
R53 VP.n30 VP.n29 62.5352
R54 VP.n65 VP.n64 50.6471
R55 VP.n73 VP.n14 41.9503
R56 VP.n102 VP.n2 41.9503
R57 VP.n56 VP.n19 41.9503
R58 VP.n84 VP.n10 40.979
R59 VP.n91 VP.n6 40.979
R60 VP.n45 VP.n23 40.979
R61 VP.n38 VP.n27 40.979
R62 VP.n80 VP.n10 40.0078
R63 VP.n95 VP.n6 40.0078
R64 VP.n49 VP.n23 40.0078
R65 VP.n34 VP.n27 40.0078
R66 VP.n69 VP.n14 39.0365
R67 VP.n106 VP.n2 39.0365
R68 VP.n60 VP.n19 39.0365
R69 VP.n16 VP.t7 35.7692
R70 VP.n12 VP.t9 35.7692
R71 VP.n8 VP.t1 35.7692
R72 VP.n4 VP.t0 35.7692
R73 VP.n0 VP.t3 35.7692
R74 VP.n17 VP.t6 35.7692
R75 VP.n21 VP.t4 35.7692
R76 VP.n25 VP.t8 35.7692
R77 VP.n29 VP.t5 35.7692
R78 VP.n68 VP.n67 24.4675
R79 VP.n69 VP.n68 24.4675
R80 VP.n74 VP.n73 24.4675
R81 VP.n75 VP.n74 24.4675
R82 VP.n79 VP.n78 24.4675
R83 VP.n80 VP.n79 24.4675
R84 VP.n85 VP.n84 24.4675
R85 VP.n86 VP.n85 24.4675
R86 VP.n90 VP.n89 24.4675
R87 VP.n91 VP.n90 24.4675
R88 VP.n96 VP.n95 24.4675
R89 VP.n97 VP.n96 24.4675
R90 VP.n101 VP.n100 24.4675
R91 VP.n102 VP.n101 24.4675
R92 VP.n107 VP.n106 24.4675
R93 VP.n108 VP.n107 24.4675
R94 VP.n61 VP.n60 24.4675
R95 VP.n62 VP.n61 24.4675
R96 VP.n50 VP.n49 24.4675
R97 VP.n51 VP.n50 24.4675
R98 VP.n55 VP.n54 24.4675
R99 VP.n56 VP.n55 24.4675
R100 VP.n39 VP.n38 24.4675
R101 VP.n40 VP.n39 24.4675
R102 VP.n44 VP.n43 24.4675
R103 VP.n45 VP.n44 24.4675
R104 VP.n33 VP.n32 24.4675
R105 VP.n34 VP.n33 24.4675
R106 VP.n75 VP.n12 12.7233
R107 VP.n100 VP.n4 12.7233
R108 VP.n54 VP.n21 12.7233
R109 VP.n86 VP.n8 12.234
R110 VP.n89 VP.n8 12.234
R111 VP.n40 VP.n25 12.234
R112 VP.n43 VP.n25 12.234
R113 VP.n78 VP.n12 11.7447
R114 VP.n97 VP.n4 11.7447
R115 VP.n51 VP.n21 11.7447
R116 VP.n32 VP.n29 11.7447
R117 VP.n67 VP.n16 11.2553
R118 VP.n108 VP.n0 11.2553
R119 VP.n62 VP.n17 11.2553
R120 VP.n31 VP.n30 4.32599
R121 VP.n64 VP.n63 0.354971
R122 VP.n66 VP.n65 0.354971
R123 VP.n110 VP.n109 0.354971
R124 VP VP.n110 0.26696
R125 VP.n31 VP.n28 0.189894
R126 VP.n35 VP.n28 0.189894
R127 VP.n36 VP.n35 0.189894
R128 VP.n37 VP.n36 0.189894
R129 VP.n37 VP.n26 0.189894
R130 VP.n41 VP.n26 0.189894
R131 VP.n42 VP.n41 0.189894
R132 VP.n42 VP.n24 0.189894
R133 VP.n46 VP.n24 0.189894
R134 VP.n47 VP.n46 0.189894
R135 VP.n48 VP.n47 0.189894
R136 VP.n48 VP.n22 0.189894
R137 VP.n52 VP.n22 0.189894
R138 VP.n53 VP.n52 0.189894
R139 VP.n53 VP.n20 0.189894
R140 VP.n57 VP.n20 0.189894
R141 VP.n58 VP.n57 0.189894
R142 VP.n59 VP.n58 0.189894
R143 VP.n59 VP.n18 0.189894
R144 VP.n63 VP.n18 0.189894
R145 VP.n66 VP.n15 0.189894
R146 VP.n70 VP.n15 0.189894
R147 VP.n71 VP.n70 0.189894
R148 VP.n72 VP.n71 0.189894
R149 VP.n72 VP.n13 0.189894
R150 VP.n76 VP.n13 0.189894
R151 VP.n77 VP.n76 0.189894
R152 VP.n77 VP.n11 0.189894
R153 VP.n81 VP.n11 0.189894
R154 VP.n82 VP.n81 0.189894
R155 VP.n83 VP.n82 0.189894
R156 VP.n83 VP.n9 0.189894
R157 VP.n87 VP.n9 0.189894
R158 VP.n88 VP.n87 0.189894
R159 VP.n88 VP.n7 0.189894
R160 VP.n92 VP.n7 0.189894
R161 VP.n93 VP.n92 0.189894
R162 VP.n94 VP.n93 0.189894
R163 VP.n94 VP.n5 0.189894
R164 VP.n98 VP.n5 0.189894
R165 VP.n99 VP.n98 0.189894
R166 VP.n99 VP.n3 0.189894
R167 VP.n103 VP.n3 0.189894
R168 VP.n104 VP.n103 0.189894
R169 VP.n105 VP.n104 0.189894
R170 VP.n105 VP.n1 0.189894
R171 VP.n109 VP.n1 0.189894
R172 VDD1.n18 VDD1.n0 756.745
R173 VDD1.n43 VDD1.n25 756.745
R174 VDD1.n19 VDD1.n18 585
R175 VDD1.n17 VDD1.n16 585
R176 VDD1.n4 VDD1.n3 585
R177 VDD1.n11 VDD1.n10 585
R178 VDD1.n9 VDD1.n8 585
R179 VDD1.n34 VDD1.n33 585
R180 VDD1.n36 VDD1.n35 585
R181 VDD1.n29 VDD1.n28 585
R182 VDD1.n42 VDD1.n41 585
R183 VDD1.n44 VDD1.n43 585
R184 VDD1.n7 VDD1.t6 328.587
R185 VDD1.n32 VDD1.t8 328.587
R186 VDD1.n18 VDD1.n17 171.744
R187 VDD1.n17 VDD1.n3 171.744
R188 VDD1.n10 VDD1.n3 171.744
R189 VDD1.n10 VDD1.n9 171.744
R190 VDD1.n35 VDD1.n34 171.744
R191 VDD1.n35 VDD1.n28 171.744
R192 VDD1.n42 VDD1.n28 171.744
R193 VDD1.n43 VDD1.n42 171.744
R194 VDD1.n51 VDD1.n50 108.802
R195 VDD1.n24 VDD1.n23 106.602
R196 VDD1.n53 VDD1.n52 106.6
R197 VDD1.n49 VDD1.n48 106.6
R198 VDD1.n9 VDD1.t6 85.8723
R199 VDD1.n34 VDD1.t8 85.8723
R200 VDD1.n24 VDD1.n22 54.394
R201 VDD1.n49 VDD1.n47 54.394
R202 VDD1.n53 VDD1.n51 44.1367
R203 VDD1.n8 VDD1.n7 16.3651
R204 VDD1.n33 VDD1.n32 16.3651
R205 VDD1.n11 VDD1.n6 12.8005
R206 VDD1.n36 VDD1.n31 12.8005
R207 VDD1.n12 VDD1.n4 12.0247
R208 VDD1.n37 VDD1.n29 12.0247
R209 VDD1.n16 VDD1.n15 11.249
R210 VDD1.n41 VDD1.n40 11.249
R211 VDD1.n19 VDD1.n2 10.4732
R212 VDD1.n44 VDD1.n27 10.4732
R213 VDD1.n20 VDD1.n0 9.69747
R214 VDD1.n45 VDD1.n25 9.69747
R215 VDD1.n22 VDD1.n21 9.45567
R216 VDD1.n47 VDD1.n46 9.45567
R217 VDD1.n21 VDD1.n20 9.3005
R218 VDD1.n2 VDD1.n1 9.3005
R219 VDD1.n15 VDD1.n14 9.3005
R220 VDD1.n13 VDD1.n12 9.3005
R221 VDD1.n6 VDD1.n5 9.3005
R222 VDD1.n46 VDD1.n45 9.3005
R223 VDD1.n27 VDD1.n26 9.3005
R224 VDD1.n40 VDD1.n39 9.3005
R225 VDD1.n38 VDD1.n37 9.3005
R226 VDD1.n31 VDD1.n30 9.3005
R227 VDD1.n52 VDD1.t0 6.9312
R228 VDD1.n52 VDD1.t9 6.9312
R229 VDD1.n23 VDD1.t7 6.9312
R230 VDD1.n23 VDD1.t5 6.9312
R231 VDD1.n50 VDD1.t3 6.9312
R232 VDD1.n50 VDD1.t4 6.9312
R233 VDD1.n48 VDD1.t1 6.9312
R234 VDD1.n48 VDD1.t2 6.9312
R235 VDD1.n22 VDD1.n0 4.26717
R236 VDD1.n47 VDD1.n25 4.26717
R237 VDD1.n7 VDD1.n5 3.73474
R238 VDD1.n32 VDD1.n30 3.73474
R239 VDD1.n20 VDD1.n19 3.49141
R240 VDD1.n45 VDD1.n44 3.49141
R241 VDD1.n16 VDD1.n2 2.71565
R242 VDD1.n41 VDD1.n27 2.71565
R243 VDD1 VDD1.n53 2.19878
R244 VDD1.n15 VDD1.n4 1.93989
R245 VDD1.n40 VDD1.n29 1.93989
R246 VDD1.n12 VDD1.n11 1.16414
R247 VDD1.n37 VDD1.n36 1.16414
R248 VDD1 VDD1.n24 0.810845
R249 VDD1.n51 VDD1.n49 0.697309
R250 VDD1.n8 VDD1.n6 0.388379
R251 VDD1.n33 VDD1.n31 0.388379
R252 VDD1.n21 VDD1.n1 0.155672
R253 VDD1.n14 VDD1.n1 0.155672
R254 VDD1.n14 VDD1.n13 0.155672
R255 VDD1.n13 VDD1.n5 0.155672
R256 VDD1.n38 VDD1.n30 0.155672
R257 VDD1.n39 VDD1.n38 0.155672
R258 VDD1.n39 VDD1.n26 0.155672
R259 VDD1.n46 VDD1.n26 0.155672
R260 VTAIL.n104 VTAIL.n86 756.745
R261 VTAIL.n20 VTAIL.n2 756.745
R262 VTAIL.n80 VTAIL.n62 756.745
R263 VTAIL.n52 VTAIL.n34 756.745
R264 VTAIL.n95 VTAIL.n94 585
R265 VTAIL.n97 VTAIL.n96 585
R266 VTAIL.n90 VTAIL.n89 585
R267 VTAIL.n103 VTAIL.n102 585
R268 VTAIL.n105 VTAIL.n104 585
R269 VTAIL.n11 VTAIL.n10 585
R270 VTAIL.n13 VTAIL.n12 585
R271 VTAIL.n6 VTAIL.n5 585
R272 VTAIL.n19 VTAIL.n18 585
R273 VTAIL.n21 VTAIL.n20 585
R274 VTAIL.n81 VTAIL.n80 585
R275 VTAIL.n79 VTAIL.n78 585
R276 VTAIL.n66 VTAIL.n65 585
R277 VTAIL.n73 VTAIL.n72 585
R278 VTAIL.n71 VTAIL.n70 585
R279 VTAIL.n53 VTAIL.n52 585
R280 VTAIL.n51 VTAIL.n50 585
R281 VTAIL.n38 VTAIL.n37 585
R282 VTAIL.n45 VTAIL.n44 585
R283 VTAIL.n43 VTAIL.n42 585
R284 VTAIL.n93 VTAIL.t2 328.587
R285 VTAIL.n9 VTAIL.t16 328.587
R286 VTAIL.n69 VTAIL.t13 328.587
R287 VTAIL.n41 VTAIL.t8 328.587
R288 VTAIL.n96 VTAIL.n95 171.744
R289 VTAIL.n96 VTAIL.n89 171.744
R290 VTAIL.n103 VTAIL.n89 171.744
R291 VTAIL.n104 VTAIL.n103 171.744
R292 VTAIL.n12 VTAIL.n11 171.744
R293 VTAIL.n12 VTAIL.n5 171.744
R294 VTAIL.n19 VTAIL.n5 171.744
R295 VTAIL.n20 VTAIL.n19 171.744
R296 VTAIL.n80 VTAIL.n79 171.744
R297 VTAIL.n79 VTAIL.n65 171.744
R298 VTAIL.n72 VTAIL.n65 171.744
R299 VTAIL.n72 VTAIL.n71 171.744
R300 VTAIL.n52 VTAIL.n51 171.744
R301 VTAIL.n51 VTAIL.n37 171.744
R302 VTAIL.n44 VTAIL.n37 171.744
R303 VTAIL.n44 VTAIL.n43 171.744
R304 VTAIL.n61 VTAIL.n60 89.9223
R305 VTAIL.n59 VTAIL.n58 89.9223
R306 VTAIL.n33 VTAIL.n32 89.9223
R307 VTAIL.n31 VTAIL.n30 89.9223
R308 VTAIL.n111 VTAIL.n110 89.9221
R309 VTAIL.n1 VTAIL.n0 89.9221
R310 VTAIL.n27 VTAIL.n26 89.9221
R311 VTAIL.n29 VTAIL.n28 89.9221
R312 VTAIL.n95 VTAIL.t2 85.8723
R313 VTAIL.n11 VTAIL.t16 85.8723
R314 VTAIL.n71 VTAIL.t13 85.8723
R315 VTAIL.n43 VTAIL.t8 85.8723
R316 VTAIL.n109 VTAIL.n108 34.7066
R317 VTAIL.n25 VTAIL.n24 34.7066
R318 VTAIL.n85 VTAIL.n84 34.7066
R319 VTAIL.n57 VTAIL.n56 34.7066
R320 VTAIL.n31 VTAIL.n29 22.4272
R321 VTAIL.n109 VTAIL.n85 19.4186
R322 VTAIL.n94 VTAIL.n93 16.3651
R323 VTAIL.n10 VTAIL.n9 16.3651
R324 VTAIL.n70 VTAIL.n69 16.3651
R325 VTAIL.n42 VTAIL.n41 16.3651
R326 VTAIL.n97 VTAIL.n92 12.8005
R327 VTAIL.n13 VTAIL.n8 12.8005
R328 VTAIL.n73 VTAIL.n68 12.8005
R329 VTAIL.n45 VTAIL.n40 12.8005
R330 VTAIL.n98 VTAIL.n90 12.0247
R331 VTAIL.n14 VTAIL.n6 12.0247
R332 VTAIL.n74 VTAIL.n66 12.0247
R333 VTAIL.n46 VTAIL.n38 12.0247
R334 VTAIL.n102 VTAIL.n101 11.249
R335 VTAIL.n18 VTAIL.n17 11.249
R336 VTAIL.n78 VTAIL.n77 11.249
R337 VTAIL.n50 VTAIL.n49 11.249
R338 VTAIL.n105 VTAIL.n88 10.4732
R339 VTAIL.n21 VTAIL.n4 10.4732
R340 VTAIL.n81 VTAIL.n64 10.4732
R341 VTAIL.n53 VTAIL.n36 10.4732
R342 VTAIL.n106 VTAIL.n86 9.69747
R343 VTAIL.n22 VTAIL.n2 9.69747
R344 VTAIL.n82 VTAIL.n62 9.69747
R345 VTAIL.n54 VTAIL.n34 9.69747
R346 VTAIL.n108 VTAIL.n107 9.45567
R347 VTAIL.n24 VTAIL.n23 9.45567
R348 VTAIL.n84 VTAIL.n83 9.45567
R349 VTAIL.n56 VTAIL.n55 9.45567
R350 VTAIL.n107 VTAIL.n106 9.3005
R351 VTAIL.n88 VTAIL.n87 9.3005
R352 VTAIL.n101 VTAIL.n100 9.3005
R353 VTAIL.n99 VTAIL.n98 9.3005
R354 VTAIL.n92 VTAIL.n91 9.3005
R355 VTAIL.n23 VTAIL.n22 9.3005
R356 VTAIL.n4 VTAIL.n3 9.3005
R357 VTAIL.n17 VTAIL.n16 9.3005
R358 VTAIL.n15 VTAIL.n14 9.3005
R359 VTAIL.n8 VTAIL.n7 9.3005
R360 VTAIL.n83 VTAIL.n82 9.3005
R361 VTAIL.n64 VTAIL.n63 9.3005
R362 VTAIL.n77 VTAIL.n76 9.3005
R363 VTAIL.n75 VTAIL.n74 9.3005
R364 VTAIL.n68 VTAIL.n67 9.3005
R365 VTAIL.n55 VTAIL.n54 9.3005
R366 VTAIL.n36 VTAIL.n35 9.3005
R367 VTAIL.n49 VTAIL.n48 9.3005
R368 VTAIL.n47 VTAIL.n46 9.3005
R369 VTAIL.n40 VTAIL.n39 9.3005
R370 VTAIL.n110 VTAIL.t5 6.9312
R371 VTAIL.n110 VTAIL.t4 6.9312
R372 VTAIL.n0 VTAIL.t9 6.9312
R373 VTAIL.n0 VTAIL.t6 6.9312
R374 VTAIL.n26 VTAIL.t18 6.9312
R375 VTAIL.n26 VTAIL.t19 6.9312
R376 VTAIL.n28 VTAIL.t12 6.9312
R377 VTAIL.n28 VTAIL.t10 6.9312
R378 VTAIL.n60 VTAIL.t11 6.9312
R379 VTAIL.n60 VTAIL.t15 6.9312
R380 VTAIL.n58 VTAIL.t17 6.9312
R381 VTAIL.n58 VTAIL.t14 6.9312
R382 VTAIL.n32 VTAIL.t3 6.9312
R383 VTAIL.n32 VTAIL.t1 6.9312
R384 VTAIL.n30 VTAIL.t7 6.9312
R385 VTAIL.n30 VTAIL.t0 6.9312
R386 VTAIL.n108 VTAIL.n86 4.26717
R387 VTAIL.n24 VTAIL.n2 4.26717
R388 VTAIL.n84 VTAIL.n62 4.26717
R389 VTAIL.n56 VTAIL.n34 4.26717
R390 VTAIL.n93 VTAIL.n91 3.73474
R391 VTAIL.n9 VTAIL.n7 3.73474
R392 VTAIL.n69 VTAIL.n67 3.73474
R393 VTAIL.n41 VTAIL.n39 3.73474
R394 VTAIL.n106 VTAIL.n105 3.49141
R395 VTAIL.n22 VTAIL.n21 3.49141
R396 VTAIL.n82 VTAIL.n81 3.49141
R397 VTAIL.n54 VTAIL.n53 3.49141
R398 VTAIL.n33 VTAIL.n31 3.00912
R399 VTAIL.n57 VTAIL.n33 3.00912
R400 VTAIL.n61 VTAIL.n59 3.00912
R401 VTAIL.n85 VTAIL.n61 3.00912
R402 VTAIL.n29 VTAIL.n27 3.00912
R403 VTAIL.n27 VTAIL.n25 3.00912
R404 VTAIL.n111 VTAIL.n109 3.00912
R405 VTAIL.n102 VTAIL.n88 2.71565
R406 VTAIL.n18 VTAIL.n4 2.71565
R407 VTAIL.n78 VTAIL.n64 2.71565
R408 VTAIL.n50 VTAIL.n36 2.71565
R409 VTAIL VTAIL.n1 2.31516
R410 VTAIL.n59 VTAIL.n57 1.97464
R411 VTAIL.n25 VTAIL.n1 1.97464
R412 VTAIL.n101 VTAIL.n90 1.93989
R413 VTAIL.n17 VTAIL.n6 1.93989
R414 VTAIL.n77 VTAIL.n66 1.93989
R415 VTAIL.n49 VTAIL.n38 1.93989
R416 VTAIL.n98 VTAIL.n97 1.16414
R417 VTAIL.n14 VTAIL.n13 1.16414
R418 VTAIL.n74 VTAIL.n73 1.16414
R419 VTAIL.n46 VTAIL.n45 1.16414
R420 VTAIL VTAIL.n111 0.694465
R421 VTAIL.n94 VTAIL.n92 0.388379
R422 VTAIL.n10 VTAIL.n8 0.388379
R423 VTAIL.n70 VTAIL.n68 0.388379
R424 VTAIL.n42 VTAIL.n40 0.388379
R425 VTAIL.n99 VTAIL.n91 0.155672
R426 VTAIL.n100 VTAIL.n99 0.155672
R427 VTAIL.n100 VTAIL.n87 0.155672
R428 VTAIL.n107 VTAIL.n87 0.155672
R429 VTAIL.n15 VTAIL.n7 0.155672
R430 VTAIL.n16 VTAIL.n15 0.155672
R431 VTAIL.n16 VTAIL.n3 0.155672
R432 VTAIL.n23 VTAIL.n3 0.155672
R433 VTAIL.n83 VTAIL.n63 0.155672
R434 VTAIL.n76 VTAIL.n63 0.155672
R435 VTAIL.n76 VTAIL.n75 0.155672
R436 VTAIL.n75 VTAIL.n67 0.155672
R437 VTAIL.n55 VTAIL.n35 0.155672
R438 VTAIL.n48 VTAIL.n35 0.155672
R439 VTAIL.n48 VTAIL.n47 0.155672
R440 VTAIL.n47 VTAIL.n39 0.155672
R441 B.n378 B.n377 585
R442 B.n376 B.n137 585
R443 B.n375 B.n374 585
R444 B.n373 B.n138 585
R445 B.n372 B.n371 585
R446 B.n370 B.n139 585
R447 B.n369 B.n368 585
R448 B.n367 B.n140 585
R449 B.n366 B.n365 585
R450 B.n364 B.n141 585
R451 B.n363 B.n362 585
R452 B.n361 B.n142 585
R453 B.n360 B.n359 585
R454 B.n358 B.n143 585
R455 B.n357 B.n356 585
R456 B.n355 B.n144 585
R457 B.n354 B.n353 585
R458 B.n352 B.n145 585
R459 B.n351 B.n350 585
R460 B.n349 B.n146 585
R461 B.n347 B.n346 585
R462 B.n345 B.n149 585
R463 B.n344 B.n343 585
R464 B.n342 B.n150 585
R465 B.n341 B.n340 585
R466 B.n339 B.n151 585
R467 B.n338 B.n337 585
R468 B.n336 B.n152 585
R469 B.n335 B.n334 585
R470 B.n333 B.n153 585
R471 B.n332 B.n331 585
R472 B.n327 B.n154 585
R473 B.n326 B.n325 585
R474 B.n324 B.n155 585
R475 B.n323 B.n322 585
R476 B.n321 B.n156 585
R477 B.n320 B.n319 585
R478 B.n318 B.n157 585
R479 B.n317 B.n316 585
R480 B.n315 B.n158 585
R481 B.n314 B.n313 585
R482 B.n312 B.n159 585
R483 B.n311 B.n310 585
R484 B.n309 B.n160 585
R485 B.n308 B.n307 585
R486 B.n306 B.n161 585
R487 B.n305 B.n304 585
R488 B.n303 B.n162 585
R489 B.n302 B.n301 585
R490 B.n300 B.n163 585
R491 B.n379 B.n136 585
R492 B.n381 B.n380 585
R493 B.n382 B.n135 585
R494 B.n384 B.n383 585
R495 B.n385 B.n134 585
R496 B.n387 B.n386 585
R497 B.n388 B.n133 585
R498 B.n390 B.n389 585
R499 B.n391 B.n132 585
R500 B.n393 B.n392 585
R501 B.n394 B.n131 585
R502 B.n396 B.n395 585
R503 B.n397 B.n130 585
R504 B.n399 B.n398 585
R505 B.n400 B.n129 585
R506 B.n402 B.n401 585
R507 B.n403 B.n128 585
R508 B.n405 B.n404 585
R509 B.n406 B.n127 585
R510 B.n408 B.n407 585
R511 B.n409 B.n126 585
R512 B.n411 B.n410 585
R513 B.n412 B.n125 585
R514 B.n414 B.n413 585
R515 B.n415 B.n124 585
R516 B.n417 B.n416 585
R517 B.n418 B.n123 585
R518 B.n420 B.n419 585
R519 B.n421 B.n122 585
R520 B.n423 B.n422 585
R521 B.n424 B.n121 585
R522 B.n426 B.n425 585
R523 B.n427 B.n120 585
R524 B.n429 B.n428 585
R525 B.n430 B.n119 585
R526 B.n432 B.n431 585
R527 B.n433 B.n118 585
R528 B.n435 B.n434 585
R529 B.n436 B.n117 585
R530 B.n438 B.n437 585
R531 B.n439 B.n116 585
R532 B.n441 B.n440 585
R533 B.n442 B.n115 585
R534 B.n444 B.n443 585
R535 B.n445 B.n114 585
R536 B.n447 B.n446 585
R537 B.n448 B.n113 585
R538 B.n450 B.n449 585
R539 B.n451 B.n112 585
R540 B.n453 B.n452 585
R541 B.n454 B.n111 585
R542 B.n456 B.n455 585
R543 B.n457 B.n110 585
R544 B.n459 B.n458 585
R545 B.n460 B.n109 585
R546 B.n462 B.n461 585
R547 B.n463 B.n108 585
R548 B.n465 B.n464 585
R549 B.n466 B.n107 585
R550 B.n468 B.n467 585
R551 B.n469 B.n106 585
R552 B.n471 B.n470 585
R553 B.n472 B.n105 585
R554 B.n474 B.n473 585
R555 B.n475 B.n104 585
R556 B.n477 B.n476 585
R557 B.n478 B.n103 585
R558 B.n480 B.n479 585
R559 B.n481 B.n102 585
R560 B.n483 B.n482 585
R561 B.n484 B.n101 585
R562 B.n486 B.n485 585
R563 B.n487 B.n100 585
R564 B.n489 B.n488 585
R565 B.n490 B.n99 585
R566 B.n492 B.n491 585
R567 B.n493 B.n98 585
R568 B.n495 B.n494 585
R569 B.n496 B.n97 585
R570 B.n498 B.n497 585
R571 B.n499 B.n96 585
R572 B.n501 B.n500 585
R573 B.n502 B.n95 585
R574 B.n504 B.n503 585
R575 B.n505 B.n94 585
R576 B.n507 B.n506 585
R577 B.n508 B.n93 585
R578 B.n510 B.n509 585
R579 B.n511 B.n92 585
R580 B.n513 B.n512 585
R581 B.n514 B.n91 585
R582 B.n516 B.n515 585
R583 B.n517 B.n90 585
R584 B.n519 B.n518 585
R585 B.n520 B.n89 585
R586 B.n522 B.n521 585
R587 B.n523 B.n88 585
R588 B.n525 B.n524 585
R589 B.n526 B.n87 585
R590 B.n528 B.n527 585
R591 B.n529 B.n86 585
R592 B.n531 B.n530 585
R593 B.n532 B.n85 585
R594 B.n534 B.n533 585
R595 B.n535 B.n84 585
R596 B.n537 B.n536 585
R597 B.n538 B.n83 585
R598 B.n540 B.n539 585
R599 B.n541 B.n82 585
R600 B.n543 B.n542 585
R601 B.n544 B.n81 585
R602 B.n546 B.n545 585
R603 B.n547 B.n80 585
R604 B.n549 B.n548 585
R605 B.n550 B.n79 585
R606 B.n552 B.n551 585
R607 B.n553 B.n78 585
R608 B.n555 B.n554 585
R609 B.n556 B.n77 585
R610 B.n558 B.n557 585
R611 B.n559 B.n76 585
R612 B.n561 B.n560 585
R613 B.n562 B.n75 585
R614 B.n564 B.n563 585
R615 B.n565 B.n74 585
R616 B.n567 B.n566 585
R617 B.n568 B.n73 585
R618 B.n570 B.n569 585
R619 B.n571 B.n72 585
R620 B.n573 B.n572 585
R621 B.n574 B.n71 585
R622 B.n576 B.n575 585
R623 B.n577 B.n70 585
R624 B.n579 B.n578 585
R625 B.n580 B.n69 585
R626 B.n582 B.n581 585
R627 B.n583 B.n68 585
R628 B.n585 B.n584 585
R629 B.n586 B.n67 585
R630 B.n588 B.n587 585
R631 B.n664 B.n663 585
R632 B.n662 B.n37 585
R633 B.n661 B.n660 585
R634 B.n659 B.n38 585
R635 B.n658 B.n657 585
R636 B.n656 B.n39 585
R637 B.n655 B.n654 585
R638 B.n653 B.n40 585
R639 B.n652 B.n651 585
R640 B.n650 B.n41 585
R641 B.n649 B.n648 585
R642 B.n647 B.n42 585
R643 B.n646 B.n645 585
R644 B.n644 B.n43 585
R645 B.n643 B.n642 585
R646 B.n641 B.n44 585
R647 B.n640 B.n639 585
R648 B.n638 B.n45 585
R649 B.n637 B.n636 585
R650 B.n635 B.n46 585
R651 B.n634 B.n633 585
R652 B.n632 B.n47 585
R653 B.n631 B.n630 585
R654 B.n629 B.n51 585
R655 B.n628 B.n627 585
R656 B.n626 B.n52 585
R657 B.n625 B.n624 585
R658 B.n623 B.n53 585
R659 B.n622 B.n621 585
R660 B.n620 B.n54 585
R661 B.n618 B.n617 585
R662 B.n616 B.n57 585
R663 B.n615 B.n614 585
R664 B.n613 B.n58 585
R665 B.n612 B.n611 585
R666 B.n610 B.n59 585
R667 B.n609 B.n608 585
R668 B.n607 B.n60 585
R669 B.n606 B.n605 585
R670 B.n604 B.n61 585
R671 B.n603 B.n602 585
R672 B.n601 B.n62 585
R673 B.n600 B.n599 585
R674 B.n598 B.n63 585
R675 B.n597 B.n596 585
R676 B.n595 B.n64 585
R677 B.n594 B.n593 585
R678 B.n592 B.n65 585
R679 B.n591 B.n590 585
R680 B.n589 B.n66 585
R681 B.n665 B.n36 585
R682 B.n667 B.n666 585
R683 B.n668 B.n35 585
R684 B.n670 B.n669 585
R685 B.n671 B.n34 585
R686 B.n673 B.n672 585
R687 B.n674 B.n33 585
R688 B.n676 B.n675 585
R689 B.n677 B.n32 585
R690 B.n679 B.n678 585
R691 B.n680 B.n31 585
R692 B.n682 B.n681 585
R693 B.n683 B.n30 585
R694 B.n685 B.n684 585
R695 B.n686 B.n29 585
R696 B.n688 B.n687 585
R697 B.n689 B.n28 585
R698 B.n691 B.n690 585
R699 B.n692 B.n27 585
R700 B.n694 B.n693 585
R701 B.n695 B.n26 585
R702 B.n697 B.n696 585
R703 B.n698 B.n25 585
R704 B.n700 B.n699 585
R705 B.n701 B.n24 585
R706 B.n703 B.n702 585
R707 B.n704 B.n23 585
R708 B.n706 B.n705 585
R709 B.n707 B.n22 585
R710 B.n709 B.n708 585
R711 B.n710 B.n21 585
R712 B.n712 B.n711 585
R713 B.n713 B.n20 585
R714 B.n715 B.n714 585
R715 B.n716 B.n19 585
R716 B.n718 B.n717 585
R717 B.n719 B.n18 585
R718 B.n721 B.n720 585
R719 B.n722 B.n17 585
R720 B.n724 B.n723 585
R721 B.n725 B.n16 585
R722 B.n727 B.n726 585
R723 B.n728 B.n15 585
R724 B.n730 B.n729 585
R725 B.n731 B.n14 585
R726 B.n733 B.n732 585
R727 B.n734 B.n13 585
R728 B.n736 B.n735 585
R729 B.n737 B.n12 585
R730 B.n739 B.n738 585
R731 B.n740 B.n11 585
R732 B.n742 B.n741 585
R733 B.n743 B.n10 585
R734 B.n745 B.n744 585
R735 B.n746 B.n9 585
R736 B.n748 B.n747 585
R737 B.n749 B.n8 585
R738 B.n751 B.n750 585
R739 B.n752 B.n7 585
R740 B.n754 B.n753 585
R741 B.n755 B.n6 585
R742 B.n757 B.n756 585
R743 B.n758 B.n5 585
R744 B.n760 B.n759 585
R745 B.n761 B.n4 585
R746 B.n763 B.n762 585
R747 B.n764 B.n3 585
R748 B.n766 B.n765 585
R749 B.n767 B.n0 585
R750 B.n2 B.n1 585
R751 B.n198 B.n197 585
R752 B.n200 B.n199 585
R753 B.n201 B.n196 585
R754 B.n203 B.n202 585
R755 B.n204 B.n195 585
R756 B.n206 B.n205 585
R757 B.n207 B.n194 585
R758 B.n209 B.n208 585
R759 B.n210 B.n193 585
R760 B.n212 B.n211 585
R761 B.n213 B.n192 585
R762 B.n215 B.n214 585
R763 B.n216 B.n191 585
R764 B.n218 B.n217 585
R765 B.n219 B.n190 585
R766 B.n221 B.n220 585
R767 B.n222 B.n189 585
R768 B.n224 B.n223 585
R769 B.n225 B.n188 585
R770 B.n227 B.n226 585
R771 B.n228 B.n187 585
R772 B.n230 B.n229 585
R773 B.n231 B.n186 585
R774 B.n233 B.n232 585
R775 B.n234 B.n185 585
R776 B.n236 B.n235 585
R777 B.n237 B.n184 585
R778 B.n239 B.n238 585
R779 B.n240 B.n183 585
R780 B.n242 B.n241 585
R781 B.n243 B.n182 585
R782 B.n245 B.n244 585
R783 B.n246 B.n181 585
R784 B.n248 B.n247 585
R785 B.n249 B.n180 585
R786 B.n251 B.n250 585
R787 B.n252 B.n179 585
R788 B.n254 B.n253 585
R789 B.n255 B.n178 585
R790 B.n257 B.n256 585
R791 B.n258 B.n177 585
R792 B.n260 B.n259 585
R793 B.n261 B.n176 585
R794 B.n263 B.n262 585
R795 B.n264 B.n175 585
R796 B.n266 B.n265 585
R797 B.n267 B.n174 585
R798 B.n269 B.n268 585
R799 B.n270 B.n173 585
R800 B.n272 B.n271 585
R801 B.n273 B.n172 585
R802 B.n275 B.n274 585
R803 B.n276 B.n171 585
R804 B.n278 B.n277 585
R805 B.n279 B.n170 585
R806 B.n281 B.n280 585
R807 B.n282 B.n169 585
R808 B.n284 B.n283 585
R809 B.n285 B.n168 585
R810 B.n287 B.n286 585
R811 B.n288 B.n167 585
R812 B.n290 B.n289 585
R813 B.n291 B.n166 585
R814 B.n293 B.n292 585
R815 B.n294 B.n165 585
R816 B.n296 B.n295 585
R817 B.n297 B.n164 585
R818 B.n299 B.n298 585
R819 B.n300 B.n299 516.524
R820 B.n377 B.n136 516.524
R821 B.n587 B.n66 516.524
R822 B.n665 B.n664 516.524
R823 B.n147 B.t10 313.774
R824 B.n55 B.t2 313.774
R825 B.n328 B.t4 313.774
R826 B.n48 B.t8 313.774
R827 B.n769 B.n768 256.663
R828 B.n148 B.t11 246.09
R829 B.n56 B.t1 246.09
R830 B.n329 B.t5 246.089
R831 B.n49 B.t7 246.089
R832 B.n328 B.t3 244.529
R833 B.n147 B.t9 244.529
R834 B.n55 B.t0 244.529
R835 B.n48 B.t6 244.529
R836 B.n768 B.n767 235.042
R837 B.n768 B.n2 235.042
R838 B.n301 B.n300 163.367
R839 B.n301 B.n162 163.367
R840 B.n305 B.n162 163.367
R841 B.n306 B.n305 163.367
R842 B.n307 B.n306 163.367
R843 B.n307 B.n160 163.367
R844 B.n311 B.n160 163.367
R845 B.n312 B.n311 163.367
R846 B.n313 B.n312 163.367
R847 B.n313 B.n158 163.367
R848 B.n317 B.n158 163.367
R849 B.n318 B.n317 163.367
R850 B.n319 B.n318 163.367
R851 B.n319 B.n156 163.367
R852 B.n323 B.n156 163.367
R853 B.n324 B.n323 163.367
R854 B.n325 B.n324 163.367
R855 B.n325 B.n154 163.367
R856 B.n332 B.n154 163.367
R857 B.n333 B.n332 163.367
R858 B.n334 B.n333 163.367
R859 B.n334 B.n152 163.367
R860 B.n338 B.n152 163.367
R861 B.n339 B.n338 163.367
R862 B.n340 B.n339 163.367
R863 B.n340 B.n150 163.367
R864 B.n344 B.n150 163.367
R865 B.n345 B.n344 163.367
R866 B.n346 B.n345 163.367
R867 B.n346 B.n146 163.367
R868 B.n351 B.n146 163.367
R869 B.n352 B.n351 163.367
R870 B.n353 B.n352 163.367
R871 B.n353 B.n144 163.367
R872 B.n357 B.n144 163.367
R873 B.n358 B.n357 163.367
R874 B.n359 B.n358 163.367
R875 B.n359 B.n142 163.367
R876 B.n363 B.n142 163.367
R877 B.n364 B.n363 163.367
R878 B.n365 B.n364 163.367
R879 B.n365 B.n140 163.367
R880 B.n369 B.n140 163.367
R881 B.n370 B.n369 163.367
R882 B.n371 B.n370 163.367
R883 B.n371 B.n138 163.367
R884 B.n375 B.n138 163.367
R885 B.n376 B.n375 163.367
R886 B.n377 B.n376 163.367
R887 B.n587 B.n586 163.367
R888 B.n586 B.n585 163.367
R889 B.n585 B.n68 163.367
R890 B.n581 B.n68 163.367
R891 B.n581 B.n580 163.367
R892 B.n580 B.n579 163.367
R893 B.n579 B.n70 163.367
R894 B.n575 B.n70 163.367
R895 B.n575 B.n574 163.367
R896 B.n574 B.n573 163.367
R897 B.n573 B.n72 163.367
R898 B.n569 B.n72 163.367
R899 B.n569 B.n568 163.367
R900 B.n568 B.n567 163.367
R901 B.n567 B.n74 163.367
R902 B.n563 B.n74 163.367
R903 B.n563 B.n562 163.367
R904 B.n562 B.n561 163.367
R905 B.n561 B.n76 163.367
R906 B.n557 B.n76 163.367
R907 B.n557 B.n556 163.367
R908 B.n556 B.n555 163.367
R909 B.n555 B.n78 163.367
R910 B.n551 B.n78 163.367
R911 B.n551 B.n550 163.367
R912 B.n550 B.n549 163.367
R913 B.n549 B.n80 163.367
R914 B.n545 B.n80 163.367
R915 B.n545 B.n544 163.367
R916 B.n544 B.n543 163.367
R917 B.n543 B.n82 163.367
R918 B.n539 B.n82 163.367
R919 B.n539 B.n538 163.367
R920 B.n538 B.n537 163.367
R921 B.n537 B.n84 163.367
R922 B.n533 B.n84 163.367
R923 B.n533 B.n532 163.367
R924 B.n532 B.n531 163.367
R925 B.n531 B.n86 163.367
R926 B.n527 B.n86 163.367
R927 B.n527 B.n526 163.367
R928 B.n526 B.n525 163.367
R929 B.n525 B.n88 163.367
R930 B.n521 B.n88 163.367
R931 B.n521 B.n520 163.367
R932 B.n520 B.n519 163.367
R933 B.n519 B.n90 163.367
R934 B.n515 B.n90 163.367
R935 B.n515 B.n514 163.367
R936 B.n514 B.n513 163.367
R937 B.n513 B.n92 163.367
R938 B.n509 B.n92 163.367
R939 B.n509 B.n508 163.367
R940 B.n508 B.n507 163.367
R941 B.n507 B.n94 163.367
R942 B.n503 B.n94 163.367
R943 B.n503 B.n502 163.367
R944 B.n502 B.n501 163.367
R945 B.n501 B.n96 163.367
R946 B.n497 B.n96 163.367
R947 B.n497 B.n496 163.367
R948 B.n496 B.n495 163.367
R949 B.n495 B.n98 163.367
R950 B.n491 B.n98 163.367
R951 B.n491 B.n490 163.367
R952 B.n490 B.n489 163.367
R953 B.n489 B.n100 163.367
R954 B.n485 B.n100 163.367
R955 B.n485 B.n484 163.367
R956 B.n484 B.n483 163.367
R957 B.n483 B.n102 163.367
R958 B.n479 B.n102 163.367
R959 B.n479 B.n478 163.367
R960 B.n478 B.n477 163.367
R961 B.n477 B.n104 163.367
R962 B.n473 B.n104 163.367
R963 B.n473 B.n472 163.367
R964 B.n472 B.n471 163.367
R965 B.n471 B.n106 163.367
R966 B.n467 B.n106 163.367
R967 B.n467 B.n466 163.367
R968 B.n466 B.n465 163.367
R969 B.n465 B.n108 163.367
R970 B.n461 B.n108 163.367
R971 B.n461 B.n460 163.367
R972 B.n460 B.n459 163.367
R973 B.n459 B.n110 163.367
R974 B.n455 B.n110 163.367
R975 B.n455 B.n454 163.367
R976 B.n454 B.n453 163.367
R977 B.n453 B.n112 163.367
R978 B.n449 B.n112 163.367
R979 B.n449 B.n448 163.367
R980 B.n448 B.n447 163.367
R981 B.n447 B.n114 163.367
R982 B.n443 B.n114 163.367
R983 B.n443 B.n442 163.367
R984 B.n442 B.n441 163.367
R985 B.n441 B.n116 163.367
R986 B.n437 B.n116 163.367
R987 B.n437 B.n436 163.367
R988 B.n436 B.n435 163.367
R989 B.n435 B.n118 163.367
R990 B.n431 B.n118 163.367
R991 B.n431 B.n430 163.367
R992 B.n430 B.n429 163.367
R993 B.n429 B.n120 163.367
R994 B.n425 B.n120 163.367
R995 B.n425 B.n424 163.367
R996 B.n424 B.n423 163.367
R997 B.n423 B.n122 163.367
R998 B.n419 B.n122 163.367
R999 B.n419 B.n418 163.367
R1000 B.n418 B.n417 163.367
R1001 B.n417 B.n124 163.367
R1002 B.n413 B.n124 163.367
R1003 B.n413 B.n412 163.367
R1004 B.n412 B.n411 163.367
R1005 B.n411 B.n126 163.367
R1006 B.n407 B.n126 163.367
R1007 B.n407 B.n406 163.367
R1008 B.n406 B.n405 163.367
R1009 B.n405 B.n128 163.367
R1010 B.n401 B.n128 163.367
R1011 B.n401 B.n400 163.367
R1012 B.n400 B.n399 163.367
R1013 B.n399 B.n130 163.367
R1014 B.n395 B.n130 163.367
R1015 B.n395 B.n394 163.367
R1016 B.n394 B.n393 163.367
R1017 B.n393 B.n132 163.367
R1018 B.n389 B.n132 163.367
R1019 B.n389 B.n388 163.367
R1020 B.n388 B.n387 163.367
R1021 B.n387 B.n134 163.367
R1022 B.n383 B.n134 163.367
R1023 B.n383 B.n382 163.367
R1024 B.n382 B.n381 163.367
R1025 B.n381 B.n136 163.367
R1026 B.n664 B.n37 163.367
R1027 B.n660 B.n37 163.367
R1028 B.n660 B.n659 163.367
R1029 B.n659 B.n658 163.367
R1030 B.n658 B.n39 163.367
R1031 B.n654 B.n39 163.367
R1032 B.n654 B.n653 163.367
R1033 B.n653 B.n652 163.367
R1034 B.n652 B.n41 163.367
R1035 B.n648 B.n41 163.367
R1036 B.n648 B.n647 163.367
R1037 B.n647 B.n646 163.367
R1038 B.n646 B.n43 163.367
R1039 B.n642 B.n43 163.367
R1040 B.n642 B.n641 163.367
R1041 B.n641 B.n640 163.367
R1042 B.n640 B.n45 163.367
R1043 B.n636 B.n45 163.367
R1044 B.n636 B.n635 163.367
R1045 B.n635 B.n634 163.367
R1046 B.n634 B.n47 163.367
R1047 B.n630 B.n47 163.367
R1048 B.n630 B.n629 163.367
R1049 B.n629 B.n628 163.367
R1050 B.n628 B.n52 163.367
R1051 B.n624 B.n52 163.367
R1052 B.n624 B.n623 163.367
R1053 B.n623 B.n622 163.367
R1054 B.n622 B.n54 163.367
R1055 B.n617 B.n54 163.367
R1056 B.n617 B.n616 163.367
R1057 B.n616 B.n615 163.367
R1058 B.n615 B.n58 163.367
R1059 B.n611 B.n58 163.367
R1060 B.n611 B.n610 163.367
R1061 B.n610 B.n609 163.367
R1062 B.n609 B.n60 163.367
R1063 B.n605 B.n60 163.367
R1064 B.n605 B.n604 163.367
R1065 B.n604 B.n603 163.367
R1066 B.n603 B.n62 163.367
R1067 B.n599 B.n62 163.367
R1068 B.n599 B.n598 163.367
R1069 B.n598 B.n597 163.367
R1070 B.n597 B.n64 163.367
R1071 B.n593 B.n64 163.367
R1072 B.n593 B.n592 163.367
R1073 B.n592 B.n591 163.367
R1074 B.n591 B.n66 163.367
R1075 B.n666 B.n665 163.367
R1076 B.n666 B.n35 163.367
R1077 B.n670 B.n35 163.367
R1078 B.n671 B.n670 163.367
R1079 B.n672 B.n671 163.367
R1080 B.n672 B.n33 163.367
R1081 B.n676 B.n33 163.367
R1082 B.n677 B.n676 163.367
R1083 B.n678 B.n677 163.367
R1084 B.n678 B.n31 163.367
R1085 B.n682 B.n31 163.367
R1086 B.n683 B.n682 163.367
R1087 B.n684 B.n683 163.367
R1088 B.n684 B.n29 163.367
R1089 B.n688 B.n29 163.367
R1090 B.n689 B.n688 163.367
R1091 B.n690 B.n689 163.367
R1092 B.n690 B.n27 163.367
R1093 B.n694 B.n27 163.367
R1094 B.n695 B.n694 163.367
R1095 B.n696 B.n695 163.367
R1096 B.n696 B.n25 163.367
R1097 B.n700 B.n25 163.367
R1098 B.n701 B.n700 163.367
R1099 B.n702 B.n701 163.367
R1100 B.n702 B.n23 163.367
R1101 B.n706 B.n23 163.367
R1102 B.n707 B.n706 163.367
R1103 B.n708 B.n707 163.367
R1104 B.n708 B.n21 163.367
R1105 B.n712 B.n21 163.367
R1106 B.n713 B.n712 163.367
R1107 B.n714 B.n713 163.367
R1108 B.n714 B.n19 163.367
R1109 B.n718 B.n19 163.367
R1110 B.n719 B.n718 163.367
R1111 B.n720 B.n719 163.367
R1112 B.n720 B.n17 163.367
R1113 B.n724 B.n17 163.367
R1114 B.n725 B.n724 163.367
R1115 B.n726 B.n725 163.367
R1116 B.n726 B.n15 163.367
R1117 B.n730 B.n15 163.367
R1118 B.n731 B.n730 163.367
R1119 B.n732 B.n731 163.367
R1120 B.n732 B.n13 163.367
R1121 B.n736 B.n13 163.367
R1122 B.n737 B.n736 163.367
R1123 B.n738 B.n737 163.367
R1124 B.n738 B.n11 163.367
R1125 B.n742 B.n11 163.367
R1126 B.n743 B.n742 163.367
R1127 B.n744 B.n743 163.367
R1128 B.n744 B.n9 163.367
R1129 B.n748 B.n9 163.367
R1130 B.n749 B.n748 163.367
R1131 B.n750 B.n749 163.367
R1132 B.n750 B.n7 163.367
R1133 B.n754 B.n7 163.367
R1134 B.n755 B.n754 163.367
R1135 B.n756 B.n755 163.367
R1136 B.n756 B.n5 163.367
R1137 B.n760 B.n5 163.367
R1138 B.n761 B.n760 163.367
R1139 B.n762 B.n761 163.367
R1140 B.n762 B.n3 163.367
R1141 B.n766 B.n3 163.367
R1142 B.n767 B.n766 163.367
R1143 B.n198 B.n2 163.367
R1144 B.n199 B.n198 163.367
R1145 B.n199 B.n196 163.367
R1146 B.n203 B.n196 163.367
R1147 B.n204 B.n203 163.367
R1148 B.n205 B.n204 163.367
R1149 B.n205 B.n194 163.367
R1150 B.n209 B.n194 163.367
R1151 B.n210 B.n209 163.367
R1152 B.n211 B.n210 163.367
R1153 B.n211 B.n192 163.367
R1154 B.n215 B.n192 163.367
R1155 B.n216 B.n215 163.367
R1156 B.n217 B.n216 163.367
R1157 B.n217 B.n190 163.367
R1158 B.n221 B.n190 163.367
R1159 B.n222 B.n221 163.367
R1160 B.n223 B.n222 163.367
R1161 B.n223 B.n188 163.367
R1162 B.n227 B.n188 163.367
R1163 B.n228 B.n227 163.367
R1164 B.n229 B.n228 163.367
R1165 B.n229 B.n186 163.367
R1166 B.n233 B.n186 163.367
R1167 B.n234 B.n233 163.367
R1168 B.n235 B.n234 163.367
R1169 B.n235 B.n184 163.367
R1170 B.n239 B.n184 163.367
R1171 B.n240 B.n239 163.367
R1172 B.n241 B.n240 163.367
R1173 B.n241 B.n182 163.367
R1174 B.n245 B.n182 163.367
R1175 B.n246 B.n245 163.367
R1176 B.n247 B.n246 163.367
R1177 B.n247 B.n180 163.367
R1178 B.n251 B.n180 163.367
R1179 B.n252 B.n251 163.367
R1180 B.n253 B.n252 163.367
R1181 B.n253 B.n178 163.367
R1182 B.n257 B.n178 163.367
R1183 B.n258 B.n257 163.367
R1184 B.n259 B.n258 163.367
R1185 B.n259 B.n176 163.367
R1186 B.n263 B.n176 163.367
R1187 B.n264 B.n263 163.367
R1188 B.n265 B.n264 163.367
R1189 B.n265 B.n174 163.367
R1190 B.n269 B.n174 163.367
R1191 B.n270 B.n269 163.367
R1192 B.n271 B.n270 163.367
R1193 B.n271 B.n172 163.367
R1194 B.n275 B.n172 163.367
R1195 B.n276 B.n275 163.367
R1196 B.n277 B.n276 163.367
R1197 B.n277 B.n170 163.367
R1198 B.n281 B.n170 163.367
R1199 B.n282 B.n281 163.367
R1200 B.n283 B.n282 163.367
R1201 B.n283 B.n168 163.367
R1202 B.n287 B.n168 163.367
R1203 B.n288 B.n287 163.367
R1204 B.n289 B.n288 163.367
R1205 B.n289 B.n166 163.367
R1206 B.n293 B.n166 163.367
R1207 B.n294 B.n293 163.367
R1208 B.n295 B.n294 163.367
R1209 B.n295 B.n164 163.367
R1210 B.n299 B.n164 163.367
R1211 B.n329 B.n328 67.6854
R1212 B.n148 B.n147 67.6854
R1213 B.n56 B.n55 67.6854
R1214 B.n49 B.n48 67.6854
R1215 B.n330 B.n329 59.5399
R1216 B.n348 B.n148 59.5399
R1217 B.n619 B.n56 59.5399
R1218 B.n50 B.n49 59.5399
R1219 B.n663 B.n36 33.5615
R1220 B.n589 B.n588 33.5615
R1221 B.n379 B.n378 33.5615
R1222 B.n298 B.n163 33.5615
R1223 B B.n769 18.0485
R1224 B.n667 B.n36 10.6151
R1225 B.n668 B.n667 10.6151
R1226 B.n669 B.n668 10.6151
R1227 B.n669 B.n34 10.6151
R1228 B.n673 B.n34 10.6151
R1229 B.n674 B.n673 10.6151
R1230 B.n675 B.n674 10.6151
R1231 B.n675 B.n32 10.6151
R1232 B.n679 B.n32 10.6151
R1233 B.n680 B.n679 10.6151
R1234 B.n681 B.n680 10.6151
R1235 B.n681 B.n30 10.6151
R1236 B.n685 B.n30 10.6151
R1237 B.n686 B.n685 10.6151
R1238 B.n687 B.n686 10.6151
R1239 B.n687 B.n28 10.6151
R1240 B.n691 B.n28 10.6151
R1241 B.n692 B.n691 10.6151
R1242 B.n693 B.n692 10.6151
R1243 B.n693 B.n26 10.6151
R1244 B.n697 B.n26 10.6151
R1245 B.n698 B.n697 10.6151
R1246 B.n699 B.n698 10.6151
R1247 B.n699 B.n24 10.6151
R1248 B.n703 B.n24 10.6151
R1249 B.n704 B.n703 10.6151
R1250 B.n705 B.n704 10.6151
R1251 B.n705 B.n22 10.6151
R1252 B.n709 B.n22 10.6151
R1253 B.n710 B.n709 10.6151
R1254 B.n711 B.n710 10.6151
R1255 B.n711 B.n20 10.6151
R1256 B.n715 B.n20 10.6151
R1257 B.n716 B.n715 10.6151
R1258 B.n717 B.n716 10.6151
R1259 B.n717 B.n18 10.6151
R1260 B.n721 B.n18 10.6151
R1261 B.n722 B.n721 10.6151
R1262 B.n723 B.n722 10.6151
R1263 B.n723 B.n16 10.6151
R1264 B.n727 B.n16 10.6151
R1265 B.n728 B.n727 10.6151
R1266 B.n729 B.n728 10.6151
R1267 B.n729 B.n14 10.6151
R1268 B.n733 B.n14 10.6151
R1269 B.n734 B.n733 10.6151
R1270 B.n735 B.n734 10.6151
R1271 B.n735 B.n12 10.6151
R1272 B.n739 B.n12 10.6151
R1273 B.n740 B.n739 10.6151
R1274 B.n741 B.n740 10.6151
R1275 B.n741 B.n10 10.6151
R1276 B.n745 B.n10 10.6151
R1277 B.n746 B.n745 10.6151
R1278 B.n747 B.n746 10.6151
R1279 B.n747 B.n8 10.6151
R1280 B.n751 B.n8 10.6151
R1281 B.n752 B.n751 10.6151
R1282 B.n753 B.n752 10.6151
R1283 B.n753 B.n6 10.6151
R1284 B.n757 B.n6 10.6151
R1285 B.n758 B.n757 10.6151
R1286 B.n759 B.n758 10.6151
R1287 B.n759 B.n4 10.6151
R1288 B.n763 B.n4 10.6151
R1289 B.n764 B.n763 10.6151
R1290 B.n765 B.n764 10.6151
R1291 B.n765 B.n0 10.6151
R1292 B.n663 B.n662 10.6151
R1293 B.n662 B.n661 10.6151
R1294 B.n661 B.n38 10.6151
R1295 B.n657 B.n38 10.6151
R1296 B.n657 B.n656 10.6151
R1297 B.n656 B.n655 10.6151
R1298 B.n655 B.n40 10.6151
R1299 B.n651 B.n40 10.6151
R1300 B.n651 B.n650 10.6151
R1301 B.n650 B.n649 10.6151
R1302 B.n649 B.n42 10.6151
R1303 B.n645 B.n42 10.6151
R1304 B.n645 B.n644 10.6151
R1305 B.n644 B.n643 10.6151
R1306 B.n643 B.n44 10.6151
R1307 B.n639 B.n44 10.6151
R1308 B.n639 B.n638 10.6151
R1309 B.n638 B.n637 10.6151
R1310 B.n637 B.n46 10.6151
R1311 B.n633 B.n632 10.6151
R1312 B.n632 B.n631 10.6151
R1313 B.n631 B.n51 10.6151
R1314 B.n627 B.n51 10.6151
R1315 B.n627 B.n626 10.6151
R1316 B.n626 B.n625 10.6151
R1317 B.n625 B.n53 10.6151
R1318 B.n621 B.n53 10.6151
R1319 B.n621 B.n620 10.6151
R1320 B.n618 B.n57 10.6151
R1321 B.n614 B.n57 10.6151
R1322 B.n614 B.n613 10.6151
R1323 B.n613 B.n612 10.6151
R1324 B.n612 B.n59 10.6151
R1325 B.n608 B.n59 10.6151
R1326 B.n608 B.n607 10.6151
R1327 B.n607 B.n606 10.6151
R1328 B.n606 B.n61 10.6151
R1329 B.n602 B.n61 10.6151
R1330 B.n602 B.n601 10.6151
R1331 B.n601 B.n600 10.6151
R1332 B.n600 B.n63 10.6151
R1333 B.n596 B.n63 10.6151
R1334 B.n596 B.n595 10.6151
R1335 B.n595 B.n594 10.6151
R1336 B.n594 B.n65 10.6151
R1337 B.n590 B.n65 10.6151
R1338 B.n590 B.n589 10.6151
R1339 B.n588 B.n67 10.6151
R1340 B.n584 B.n67 10.6151
R1341 B.n584 B.n583 10.6151
R1342 B.n583 B.n582 10.6151
R1343 B.n582 B.n69 10.6151
R1344 B.n578 B.n69 10.6151
R1345 B.n578 B.n577 10.6151
R1346 B.n577 B.n576 10.6151
R1347 B.n576 B.n71 10.6151
R1348 B.n572 B.n71 10.6151
R1349 B.n572 B.n571 10.6151
R1350 B.n571 B.n570 10.6151
R1351 B.n570 B.n73 10.6151
R1352 B.n566 B.n73 10.6151
R1353 B.n566 B.n565 10.6151
R1354 B.n565 B.n564 10.6151
R1355 B.n564 B.n75 10.6151
R1356 B.n560 B.n75 10.6151
R1357 B.n560 B.n559 10.6151
R1358 B.n559 B.n558 10.6151
R1359 B.n558 B.n77 10.6151
R1360 B.n554 B.n77 10.6151
R1361 B.n554 B.n553 10.6151
R1362 B.n553 B.n552 10.6151
R1363 B.n552 B.n79 10.6151
R1364 B.n548 B.n79 10.6151
R1365 B.n548 B.n547 10.6151
R1366 B.n547 B.n546 10.6151
R1367 B.n546 B.n81 10.6151
R1368 B.n542 B.n81 10.6151
R1369 B.n542 B.n541 10.6151
R1370 B.n541 B.n540 10.6151
R1371 B.n540 B.n83 10.6151
R1372 B.n536 B.n83 10.6151
R1373 B.n536 B.n535 10.6151
R1374 B.n535 B.n534 10.6151
R1375 B.n534 B.n85 10.6151
R1376 B.n530 B.n85 10.6151
R1377 B.n530 B.n529 10.6151
R1378 B.n529 B.n528 10.6151
R1379 B.n528 B.n87 10.6151
R1380 B.n524 B.n87 10.6151
R1381 B.n524 B.n523 10.6151
R1382 B.n523 B.n522 10.6151
R1383 B.n522 B.n89 10.6151
R1384 B.n518 B.n89 10.6151
R1385 B.n518 B.n517 10.6151
R1386 B.n517 B.n516 10.6151
R1387 B.n516 B.n91 10.6151
R1388 B.n512 B.n91 10.6151
R1389 B.n512 B.n511 10.6151
R1390 B.n511 B.n510 10.6151
R1391 B.n510 B.n93 10.6151
R1392 B.n506 B.n93 10.6151
R1393 B.n506 B.n505 10.6151
R1394 B.n505 B.n504 10.6151
R1395 B.n504 B.n95 10.6151
R1396 B.n500 B.n95 10.6151
R1397 B.n500 B.n499 10.6151
R1398 B.n499 B.n498 10.6151
R1399 B.n498 B.n97 10.6151
R1400 B.n494 B.n97 10.6151
R1401 B.n494 B.n493 10.6151
R1402 B.n493 B.n492 10.6151
R1403 B.n492 B.n99 10.6151
R1404 B.n488 B.n99 10.6151
R1405 B.n488 B.n487 10.6151
R1406 B.n487 B.n486 10.6151
R1407 B.n486 B.n101 10.6151
R1408 B.n482 B.n101 10.6151
R1409 B.n482 B.n481 10.6151
R1410 B.n481 B.n480 10.6151
R1411 B.n480 B.n103 10.6151
R1412 B.n476 B.n103 10.6151
R1413 B.n476 B.n475 10.6151
R1414 B.n475 B.n474 10.6151
R1415 B.n474 B.n105 10.6151
R1416 B.n470 B.n105 10.6151
R1417 B.n470 B.n469 10.6151
R1418 B.n469 B.n468 10.6151
R1419 B.n468 B.n107 10.6151
R1420 B.n464 B.n107 10.6151
R1421 B.n464 B.n463 10.6151
R1422 B.n463 B.n462 10.6151
R1423 B.n462 B.n109 10.6151
R1424 B.n458 B.n109 10.6151
R1425 B.n458 B.n457 10.6151
R1426 B.n457 B.n456 10.6151
R1427 B.n456 B.n111 10.6151
R1428 B.n452 B.n111 10.6151
R1429 B.n452 B.n451 10.6151
R1430 B.n451 B.n450 10.6151
R1431 B.n450 B.n113 10.6151
R1432 B.n446 B.n113 10.6151
R1433 B.n446 B.n445 10.6151
R1434 B.n445 B.n444 10.6151
R1435 B.n444 B.n115 10.6151
R1436 B.n440 B.n115 10.6151
R1437 B.n440 B.n439 10.6151
R1438 B.n439 B.n438 10.6151
R1439 B.n438 B.n117 10.6151
R1440 B.n434 B.n117 10.6151
R1441 B.n434 B.n433 10.6151
R1442 B.n433 B.n432 10.6151
R1443 B.n432 B.n119 10.6151
R1444 B.n428 B.n119 10.6151
R1445 B.n428 B.n427 10.6151
R1446 B.n427 B.n426 10.6151
R1447 B.n426 B.n121 10.6151
R1448 B.n422 B.n121 10.6151
R1449 B.n422 B.n421 10.6151
R1450 B.n421 B.n420 10.6151
R1451 B.n420 B.n123 10.6151
R1452 B.n416 B.n123 10.6151
R1453 B.n416 B.n415 10.6151
R1454 B.n415 B.n414 10.6151
R1455 B.n414 B.n125 10.6151
R1456 B.n410 B.n125 10.6151
R1457 B.n410 B.n409 10.6151
R1458 B.n409 B.n408 10.6151
R1459 B.n408 B.n127 10.6151
R1460 B.n404 B.n127 10.6151
R1461 B.n404 B.n403 10.6151
R1462 B.n403 B.n402 10.6151
R1463 B.n402 B.n129 10.6151
R1464 B.n398 B.n129 10.6151
R1465 B.n398 B.n397 10.6151
R1466 B.n397 B.n396 10.6151
R1467 B.n396 B.n131 10.6151
R1468 B.n392 B.n131 10.6151
R1469 B.n392 B.n391 10.6151
R1470 B.n391 B.n390 10.6151
R1471 B.n390 B.n133 10.6151
R1472 B.n386 B.n133 10.6151
R1473 B.n386 B.n385 10.6151
R1474 B.n385 B.n384 10.6151
R1475 B.n384 B.n135 10.6151
R1476 B.n380 B.n135 10.6151
R1477 B.n380 B.n379 10.6151
R1478 B.n197 B.n1 10.6151
R1479 B.n200 B.n197 10.6151
R1480 B.n201 B.n200 10.6151
R1481 B.n202 B.n201 10.6151
R1482 B.n202 B.n195 10.6151
R1483 B.n206 B.n195 10.6151
R1484 B.n207 B.n206 10.6151
R1485 B.n208 B.n207 10.6151
R1486 B.n208 B.n193 10.6151
R1487 B.n212 B.n193 10.6151
R1488 B.n213 B.n212 10.6151
R1489 B.n214 B.n213 10.6151
R1490 B.n214 B.n191 10.6151
R1491 B.n218 B.n191 10.6151
R1492 B.n219 B.n218 10.6151
R1493 B.n220 B.n219 10.6151
R1494 B.n220 B.n189 10.6151
R1495 B.n224 B.n189 10.6151
R1496 B.n225 B.n224 10.6151
R1497 B.n226 B.n225 10.6151
R1498 B.n226 B.n187 10.6151
R1499 B.n230 B.n187 10.6151
R1500 B.n231 B.n230 10.6151
R1501 B.n232 B.n231 10.6151
R1502 B.n232 B.n185 10.6151
R1503 B.n236 B.n185 10.6151
R1504 B.n237 B.n236 10.6151
R1505 B.n238 B.n237 10.6151
R1506 B.n238 B.n183 10.6151
R1507 B.n242 B.n183 10.6151
R1508 B.n243 B.n242 10.6151
R1509 B.n244 B.n243 10.6151
R1510 B.n244 B.n181 10.6151
R1511 B.n248 B.n181 10.6151
R1512 B.n249 B.n248 10.6151
R1513 B.n250 B.n249 10.6151
R1514 B.n250 B.n179 10.6151
R1515 B.n254 B.n179 10.6151
R1516 B.n255 B.n254 10.6151
R1517 B.n256 B.n255 10.6151
R1518 B.n256 B.n177 10.6151
R1519 B.n260 B.n177 10.6151
R1520 B.n261 B.n260 10.6151
R1521 B.n262 B.n261 10.6151
R1522 B.n262 B.n175 10.6151
R1523 B.n266 B.n175 10.6151
R1524 B.n267 B.n266 10.6151
R1525 B.n268 B.n267 10.6151
R1526 B.n268 B.n173 10.6151
R1527 B.n272 B.n173 10.6151
R1528 B.n273 B.n272 10.6151
R1529 B.n274 B.n273 10.6151
R1530 B.n274 B.n171 10.6151
R1531 B.n278 B.n171 10.6151
R1532 B.n279 B.n278 10.6151
R1533 B.n280 B.n279 10.6151
R1534 B.n280 B.n169 10.6151
R1535 B.n284 B.n169 10.6151
R1536 B.n285 B.n284 10.6151
R1537 B.n286 B.n285 10.6151
R1538 B.n286 B.n167 10.6151
R1539 B.n290 B.n167 10.6151
R1540 B.n291 B.n290 10.6151
R1541 B.n292 B.n291 10.6151
R1542 B.n292 B.n165 10.6151
R1543 B.n296 B.n165 10.6151
R1544 B.n297 B.n296 10.6151
R1545 B.n298 B.n297 10.6151
R1546 B.n302 B.n163 10.6151
R1547 B.n303 B.n302 10.6151
R1548 B.n304 B.n303 10.6151
R1549 B.n304 B.n161 10.6151
R1550 B.n308 B.n161 10.6151
R1551 B.n309 B.n308 10.6151
R1552 B.n310 B.n309 10.6151
R1553 B.n310 B.n159 10.6151
R1554 B.n314 B.n159 10.6151
R1555 B.n315 B.n314 10.6151
R1556 B.n316 B.n315 10.6151
R1557 B.n316 B.n157 10.6151
R1558 B.n320 B.n157 10.6151
R1559 B.n321 B.n320 10.6151
R1560 B.n322 B.n321 10.6151
R1561 B.n322 B.n155 10.6151
R1562 B.n326 B.n155 10.6151
R1563 B.n327 B.n326 10.6151
R1564 B.n331 B.n327 10.6151
R1565 B.n335 B.n153 10.6151
R1566 B.n336 B.n335 10.6151
R1567 B.n337 B.n336 10.6151
R1568 B.n337 B.n151 10.6151
R1569 B.n341 B.n151 10.6151
R1570 B.n342 B.n341 10.6151
R1571 B.n343 B.n342 10.6151
R1572 B.n343 B.n149 10.6151
R1573 B.n347 B.n149 10.6151
R1574 B.n350 B.n349 10.6151
R1575 B.n350 B.n145 10.6151
R1576 B.n354 B.n145 10.6151
R1577 B.n355 B.n354 10.6151
R1578 B.n356 B.n355 10.6151
R1579 B.n356 B.n143 10.6151
R1580 B.n360 B.n143 10.6151
R1581 B.n361 B.n360 10.6151
R1582 B.n362 B.n361 10.6151
R1583 B.n362 B.n141 10.6151
R1584 B.n366 B.n141 10.6151
R1585 B.n367 B.n366 10.6151
R1586 B.n368 B.n367 10.6151
R1587 B.n368 B.n139 10.6151
R1588 B.n372 B.n139 10.6151
R1589 B.n373 B.n372 10.6151
R1590 B.n374 B.n373 10.6151
R1591 B.n374 B.n137 10.6151
R1592 B.n378 B.n137 10.6151
R1593 B.n50 B.n46 9.36635
R1594 B.n619 B.n618 9.36635
R1595 B.n331 B.n330 9.36635
R1596 B.n349 B.n348 9.36635
R1597 B.n769 B.n0 8.11757
R1598 B.n769 B.n1 8.11757
R1599 B.n633 B.n50 1.24928
R1600 B.n620 B.n619 1.24928
R1601 B.n330 B.n153 1.24928
R1602 B.n348 B.n347 1.24928
R1603 VN.n94 VN.n93 161.3
R1604 VN.n92 VN.n49 161.3
R1605 VN.n91 VN.n90 161.3
R1606 VN.n89 VN.n50 161.3
R1607 VN.n88 VN.n87 161.3
R1608 VN.n86 VN.n51 161.3
R1609 VN.n85 VN.n84 161.3
R1610 VN.n83 VN.n82 161.3
R1611 VN.n81 VN.n53 161.3
R1612 VN.n80 VN.n79 161.3
R1613 VN.n78 VN.n54 161.3
R1614 VN.n77 VN.n76 161.3
R1615 VN.n75 VN.n55 161.3
R1616 VN.n74 VN.n73 161.3
R1617 VN.n72 VN.n71 161.3
R1618 VN.n70 VN.n57 161.3
R1619 VN.n69 VN.n68 161.3
R1620 VN.n67 VN.n58 161.3
R1621 VN.n66 VN.n65 161.3
R1622 VN.n64 VN.n59 161.3
R1623 VN.n63 VN.n62 161.3
R1624 VN.n46 VN.n45 161.3
R1625 VN.n44 VN.n1 161.3
R1626 VN.n43 VN.n42 161.3
R1627 VN.n41 VN.n2 161.3
R1628 VN.n40 VN.n39 161.3
R1629 VN.n38 VN.n3 161.3
R1630 VN.n37 VN.n36 161.3
R1631 VN.n35 VN.n34 161.3
R1632 VN.n33 VN.n5 161.3
R1633 VN.n32 VN.n31 161.3
R1634 VN.n30 VN.n6 161.3
R1635 VN.n29 VN.n28 161.3
R1636 VN.n27 VN.n7 161.3
R1637 VN.n26 VN.n25 161.3
R1638 VN.n24 VN.n23 161.3
R1639 VN.n22 VN.n9 161.3
R1640 VN.n21 VN.n20 161.3
R1641 VN.n19 VN.n10 161.3
R1642 VN.n18 VN.n17 161.3
R1643 VN.n16 VN.n11 161.3
R1644 VN.n15 VN.n14 161.3
R1645 VN.n47 VN.n0 78.8126
R1646 VN.n95 VN.n48 78.8126
R1647 VN.n61 VN.t1 68.2469
R1648 VN.n13 VN.t5 68.2469
R1649 VN.n13 VN.n12 62.5352
R1650 VN.n61 VN.n60 62.5352
R1651 VN VN.n95 50.8124
R1652 VN.n39 VN.n2 41.9503
R1653 VN.n87 VN.n50 41.9503
R1654 VN.n21 VN.n10 40.979
R1655 VN.n28 VN.n6 40.979
R1656 VN.n69 VN.n58 40.979
R1657 VN.n76 VN.n54 40.979
R1658 VN.n17 VN.n10 40.0078
R1659 VN.n32 VN.n6 40.0078
R1660 VN.n65 VN.n58 40.0078
R1661 VN.n80 VN.n54 40.0078
R1662 VN.n43 VN.n2 39.0365
R1663 VN.n91 VN.n50 39.0365
R1664 VN.n12 VN.t2 35.7692
R1665 VN.n8 VN.t6 35.7692
R1666 VN.n4 VN.t4 35.7692
R1667 VN.n0 VN.t0 35.7692
R1668 VN.n60 VN.t9 35.7692
R1669 VN.n56 VN.t7 35.7692
R1670 VN.n52 VN.t8 35.7692
R1671 VN.n48 VN.t3 35.7692
R1672 VN.n16 VN.n15 24.4675
R1673 VN.n17 VN.n16 24.4675
R1674 VN.n22 VN.n21 24.4675
R1675 VN.n23 VN.n22 24.4675
R1676 VN.n27 VN.n26 24.4675
R1677 VN.n28 VN.n27 24.4675
R1678 VN.n33 VN.n32 24.4675
R1679 VN.n34 VN.n33 24.4675
R1680 VN.n38 VN.n37 24.4675
R1681 VN.n39 VN.n38 24.4675
R1682 VN.n44 VN.n43 24.4675
R1683 VN.n45 VN.n44 24.4675
R1684 VN.n65 VN.n64 24.4675
R1685 VN.n64 VN.n63 24.4675
R1686 VN.n76 VN.n75 24.4675
R1687 VN.n75 VN.n74 24.4675
R1688 VN.n71 VN.n70 24.4675
R1689 VN.n70 VN.n69 24.4675
R1690 VN.n87 VN.n86 24.4675
R1691 VN.n86 VN.n85 24.4675
R1692 VN.n82 VN.n81 24.4675
R1693 VN.n81 VN.n80 24.4675
R1694 VN.n93 VN.n92 24.4675
R1695 VN.n92 VN.n91 24.4675
R1696 VN.n37 VN.n4 12.7233
R1697 VN.n85 VN.n52 12.7233
R1698 VN.n23 VN.n8 12.234
R1699 VN.n26 VN.n8 12.234
R1700 VN.n74 VN.n56 12.234
R1701 VN.n71 VN.n56 12.234
R1702 VN.n15 VN.n12 11.7447
R1703 VN.n34 VN.n4 11.7447
R1704 VN.n63 VN.n60 11.7447
R1705 VN.n82 VN.n52 11.7447
R1706 VN.n45 VN.n0 11.2553
R1707 VN.n93 VN.n48 11.2553
R1708 VN.n14 VN.n13 4.32602
R1709 VN.n62 VN.n61 4.32602
R1710 VN.n95 VN.n94 0.354971
R1711 VN.n47 VN.n46 0.354971
R1712 VN VN.n47 0.26696
R1713 VN.n94 VN.n49 0.189894
R1714 VN.n90 VN.n49 0.189894
R1715 VN.n90 VN.n89 0.189894
R1716 VN.n89 VN.n88 0.189894
R1717 VN.n88 VN.n51 0.189894
R1718 VN.n84 VN.n51 0.189894
R1719 VN.n84 VN.n83 0.189894
R1720 VN.n83 VN.n53 0.189894
R1721 VN.n79 VN.n53 0.189894
R1722 VN.n79 VN.n78 0.189894
R1723 VN.n78 VN.n77 0.189894
R1724 VN.n77 VN.n55 0.189894
R1725 VN.n73 VN.n55 0.189894
R1726 VN.n73 VN.n72 0.189894
R1727 VN.n72 VN.n57 0.189894
R1728 VN.n68 VN.n57 0.189894
R1729 VN.n68 VN.n67 0.189894
R1730 VN.n67 VN.n66 0.189894
R1731 VN.n66 VN.n59 0.189894
R1732 VN.n62 VN.n59 0.189894
R1733 VN.n14 VN.n11 0.189894
R1734 VN.n18 VN.n11 0.189894
R1735 VN.n19 VN.n18 0.189894
R1736 VN.n20 VN.n19 0.189894
R1737 VN.n20 VN.n9 0.189894
R1738 VN.n24 VN.n9 0.189894
R1739 VN.n25 VN.n24 0.189894
R1740 VN.n25 VN.n7 0.189894
R1741 VN.n29 VN.n7 0.189894
R1742 VN.n30 VN.n29 0.189894
R1743 VN.n31 VN.n30 0.189894
R1744 VN.n31 VN.n5 0.189894
R1745 VN.n35 VN.n5 0.189894
R1746 VN.n36 VN.n35 0.189894
R1747 VN.n36 VN.n3 0.189894
R1748 VN.n40 VN.n3 0.189894
R1749 VN.n41 VN.n40 0.189894
R1750 VN.n42 VN.n41 0.189894
R1751 VN.n42 VN.n1 0.189894
R1752 VN.n46 VN.n1 0.189894
R1753 VDD2.n45 VDD2.n27 756.745
R1754 VDD2.n18 VDD2.n0 756.745
R1755 VDD2.n46 VDD2.n45 585
R1756 VDD2.n44 VDD2.n43 585
R1757 VDD2.n31 VDD2.n30 585
R1758 VDD2.n38 VDD2.n37 585
R1759 VDD2.n36 VDD2.n35 585
R1760 VDD2.n9 VDD2.n8 585
R1761 VDD2.n11 VDD2.n10 585
R1762 VDD2.n4 VDD2.n3 585
R1763 VDD2.n17 VDD2.n16 585
R1764 VDD2.n19 VDD2.n18 585
R1765 VDD2.n34 VDD2.t6 328.587
R1766 VDD2.n7 VDD2.t4 328.587
R1767 VDD2.n45 VDD2.n44 171.744
R1768 VDD2.n44 VDD2.n30 171.744
R1769 VDD2.n37 VDD2.n30 171.744
R1770 VDD2.n37 VDD2.n36 171.744
R1771 VDD2.n10 VDD2.n9 171.744
R1772 VDD2.n10 VDD2.n3 171.744
R1773 VDD2.n17 VDD2.n3 171.744
R1774 VDD2.n18 VDD2.n17 171.744
R1775 VDD2.n26 VDD2.n25 108.802
R1776 VDD2 VDD2.n53 108.799
R1777 VDD2.n52 VDD2.n51 106.602
R1778 VDD2.n24 VDD2.n23 106.6
R1779 VDD2.n36 VDD2.t6 85.8723
R1780 VDD2.n9 VDD2.t4 85.8723
R1781 VDD2.n24 VDD2.n22 54.394
R1782 VDD2.n50 VDD2.n49 51.3853
R1783 VDD2.n50 VDD2.n26 42.0493
R1784 VDD2.n35 VDD2.n34 16.3651
R1785 VDD2.n8 VDD2.n7 16.3651
R1786 VDD2.n38 VDD2.n33 12.8005
R1787 VDD2.n11 VDD2.n6 12.8005
R1788 VDD2.n39 VDD2.n31 12.0247
R1789 VDD2.n12 VDD2.n4 12.0247
R1790 VDD2.n43 VDD2.n42 11.249
R1791 VDD2.n16 VDD2.n15 11.249
R1792 VDD2.n46 VDD2.n29 10.4732
R1793 VDD2.n19 VDD2.n2 10.4732
R1794 VDD2.n47 VDD2.n27 9.69747
R1795 VDD2.n20 VDD2.n0 9.69747
R1796 VDD2.n49 VDD2.n48 9.45567
R1797 VDD2.n22 VDD2.n21 9.45567
R1798 VDD2.n48 VDD2.n47 9.3005
R1799 VDD2.n29 VDD2.n28 9.3005
R1800 VDD2.n42 VDD2.n41 9.3005
R1801 VDD2.n40 VDD2.n39 9.3005
R1802 VDD2.n33 VDD2.n32 9.3005
R1803 VDD2.n21 VDD2.n20 9.3005
R1804 VDD2.n2 VDD2.n1 9.3005
R1805 VDD2.n15 VDD2.n14 9.3005
R1806 VDD2.n13 VDD2.n12 9.3005
R1807 VDD2.n6 VDD2.n5 9.3005
R1808 VDD2.n53 VDD2.t0 6.9312
R1809 VDD2.n53 VDD2.t8 6.9312
R1810 VDD2.n51 VDD2.t1 6.9312
R1811 VDD2.n51 VDD2.t2 6.9312
R1812 VDD2.n25 VDD2.t5 6.9312
R1813 VDD2.n25 VDD2.t9 6.9312
R1814 VDD2.n23 VDD2.t7 6.9312
R1815 VDD2.n23 VDD2.t3 6.9312
R1816 VDD2.n49 VDD2.n27 4.26717
R1817 VDD2.n22 VDD2.n0 4.26717
R1818 VDD2.n34 VDD2.n32 3.73474
R1819 VDD2.n7 VDD2.n5 3.73474
R1820 VDD2.n47 VDD2.n46 3.49141
R1821 VDD2.n20 VDD2.n19 3.49141
R1822 VDD2.n52 VDD2.n50 3.00912
R1823 VDD2.n43 VDD2.n29 2.71565
R1824 VDD2.n16 VDD2.n2 2.71565
R1825 VDD2.n42 VDD2.n31 1.93989
R1826 VDD2.n15 VDD2.n4 1.93989
R1827 VDD2.n39 VDD2.n38 1.16414
R1828 VDD2.n12 VDD2.n11 1.16414
R1829 VDD2 VDD2.n52 0.810845
R1830 VDD2.n26 VDD2.n24 0.697309
R1831 VDD2.n35 VDD2.n33 0.388379
R1832 VDD2.n8 VDD2.n6 0.388379
R1833 VDD2.n48 VDD2.n28 0.155672
R1834 VDD2.n41 VDD2.n28 0.155672
R1835 VDD2.n41 VDD2.n40 0.155672
R1836 VDD2.n40 VDD2.n32 0.155672
R1837 VDD2.n13 VDD2.n5 0.155672
R1838 VDD2.n14 VDD2.n13 0.155672
R1839 VDD2.n14 VDD2.n1 0.155672
R1840 VDD2.n21 VDD2.n1 0.155672
C0 VTAIL VN 6.14238f
C1 VDD1 VTAIL 7.53054f
C2 w_n5158_n1906# VN 11.109599f
C3 VDD1 w_n5158_n1906# 2.49086f
C4 B VP 2.52515f
C5 VDD2 VN 4.65806f
C6 VDD1 VDD2 2.53565f
C7 VTAIL VP 6.15654f
C8 w_n5158_n1906# VP 11.7828f
C9 VDD1 VN 0.158184f
C10 B VTAIL 2.22724f
C11 VDD2 VP 0.658685f
C12 w_n5158_n1906# B 9.45819f
C13 w_n5158_n1906# VTAIL 2.26323f
C14 B VDD2 2.25424f
C15 VP VN 7.87592f
C16 VDD1 VP 5.15497f
C17 VDD2 VTAIL 7.587161f
C18 w_n5158_n1906# VDD2 2.66321f
C19 B VN 1.39f
C20 VDD1 B 2.11438f
C21 VDD2 VSUBS 2.305893f
C22 VDD1 VSUBS 2.028396f
C23 VTAIL VSUBS 0.710142f
C24 VN VSUBS 8.365241f
C25 VP VSUBS 4.343874f
C26 B VSUBS 5.117818f
C27 w_n5158_n1906# VSUBS 0.123359p
C28 VDD2.n0 VSUBS 0.04086f
C29 VDD2.n1 VSUBS 0.036619f
C30 VDD2.n2 VSUBS 0.019678f
C31 VDD2.n3 VSUBS 0.046511f
C32 VDD2.n4 VSUBS 0.020835f
C33 VDD2.n5 VSUBS 0.618588f
C34 VDD2.n6 VSUBS 0.019678f
C35 VDD2.t4 VSUBS 0.101746f
C36 VDD2.n7 VSUBS 0.149461f
C37 VDD2.n8 VSUBS 0.029465f
C38 VDD2.n9 VSUBS 0.034883f
C39 VDD2.n10 VSUBS 0.046511f
C40 VDD2.n11 VSUBS 0.020835f
C41 VDD2.n12 VSUBS 0.019678f
C42 VDD2.n13 VSUBS 0.036619f
C43 VDD2.n14 VSUBS 0.036619f
C44 VDD2.n15 VSUBS 0.019678f
C45 VDD2.n16 VSUBS 0.020835f
C46 VDD2.n17 VSUBS 0.046511f
C47 VDD2.n18 VSUBS 0.11472f
C48 VDD2.n19 VSUBS 0.020835f
C49 VDD2.n20 VSUBS 0.019678f
C50 VDD2.n21 VSUBS 0.091147f
C51 VDD2.n22 VSUBS 0.106959f
C52 VDD2.t7 VSUBS 0.135718f
C53 VDD2.t3 VSUBS 0.135718f
C54 VDD2.n23 VSUBS 0.837381f
C55 VDD2.n24 VSUBS 1.39112f
C56 VDD2.t5 VSUBS 0.135718f
C57 VDD2.t9 VSUBS 0.135718f
C58 VDD2.n25 VSUBS 0.861193f
C59 VDD2.n26 VSUBS 4.28327f
C60 VDD2.n27 VSUBS 0.04086f
C61 VDD2.n28 VSUBS 0.036619f
C62 VDD2.n29 VSUBS 0.019678f
C63 VDD2.n30 VSUBS 0.046511f
C64 VDD2.n31 VSUBS 0.020835f
C65 VDD2.n32 VSUBS 0.618588f
C66 VDD2.n33 VSUBS 0.019678f
C67 VDD2.t6 VSUBS 0.101746f
C68 VDD2.n34 VSUBS 0.149461f
C69 VDD2.n35 VSUBS 0.029465f
C70 VDD2.n36 VSUBS 0.034883f
C71 VDD2.n37 VSUBS 0.046511f
C72 VDD2.n38 VSUBS 0.020835f
C73 VDD2.n39 VSUBS 0.019678f
C74 VDD2.n40 VSUBS 0.036619f
C75 VDD2.n41 VSUBS 0.036619f
C76 VDD2.n42 VSUBS 0.019678f
C77 VDD2.n43 VSUBS 0.020835f
C78 VDD2.n44 VSUBS 0.046511f
C79 VDD2.n45 VSUBS 0.11472f
C80 VDD2.n46 VSUBS 0.020835f
C81 VDD2.n47 VSUBS 0.019678f
C82 VDD2.n48 VSUBS 0.091147f
C83 VDD2.n49 VSUBS 0.083217f
C84 VDD2.n50 VSUBS 3.72327f
C85 VDD2.t1 VSUBS 0.135718f
C86 VDD2.t2 VSUBS 0.135718f
C87 VDD2.n51 VSUBS 0.837385f
C88 VDD2.n52 VSUBS 0.997792f
C89 VDD2.t0 VSUBS 0.135718f
C90 VDD2.t8 VSUBS 0.135718f
C91 VDD2.n53 VSUBS 0.861148f
C92 VN.t0 VSUBS 1.39678f
C93 VN.n0 VSUBS 0.664188f
C94 VN.n1 VSUBS 0.036203f
C95 VN.n2 VSUBS 0.029373f
C96 VN.n3 VSUBS 0.036203f
C97 VN.t4 VSUBS 1.39678f
C98 VN.n4 VSUBS 0.53453f
C99 VN.n5 VSUBS 0.036203f
C100 VN.n6 VSUBS 0.02928f
C101 VN.n7 VSUBS 0.036203f
C102 VN.t6 VSUBS 1.39678f
C103 VN.n8 VSUBS 0.53453f
C104 VN.n9 VSUBS 0.036203f
C105 VN.n10 VSUBS 0.02928f
C106 VN.n11 VSUBS 0.036203f
C107 VN.t2 VSUBS 1.39678f
C108 VN.n12 VSUBS 0.652385f
C109 VN.t5 VSUBS 1.76937f
C110 VN.n13 VSUBS 0.628358f
C111 VN.n14 VSUBS 0.420838f
C112 VN.n15 VSUBS 0.050151f
C113 VN.n16 VSUBS 0.067474f
C114 VN.n17 VSUBS 0.072132f
C115 VN.n18 VSUBS 0.036203f
C116 VN.n19 VSUBS 0.036203f
C117 VN.n20 VSUBS 0.036203f
C118 VN.n21 VSUBS 0.071769f
C119 VN.n22 VSUBS 0.067474f
C120 VN.n23 VSUBS 0.050818f
C121 VN.n24 VSUBS 0.036203f
C122 VN.n25 VSUBS 0.036203f
C123 VN.n26 VSUBS 0.050818f
C124 VN.n27 VSUBS 0.067474f
C125 VN.n28 VSUBS 0.071769f
C126 VN.n29 VSUBS 0.036203f
C127 VN.n30 VSUBS 0.036203f
C128 VN.n31 VSUBS 0.036203f
C129 VN.n32 VSUBS 0.072132f
C130 VN.n33 VSUBS 0.067474f
C131 VN.n34 VSUBS 0.050151f
C132 VN.n35 VSUBS 0.036203f
C133 VN.n36 VSUBS 0.036203f
C134 VN.n37 VSUBS 0.051484f
C135 VN.n38 VSUBS 0.067474f
C136 VN.n39 VSUBS 0.071361f
C137 VN.n40 VSUBS 0.036203f
C138 VN.n41 VSUBS 0.036203f
C139 VN.n42 VSUBS 0.036203f
C140 VN.n43 VSUBS 0.072447f
C141 VN.n44 VSUBS 0.067474f
C142 VN.n45 VSUBS 0.049485f
C143 VN.n46 VSUBS 0.058431f
C144 VN.n47 VSUBS 0.089938f
C145 VN.t3 VSUBS 1.39678f
C146 VN.n48 VSUBS 0.664188f
C147 VN.n49 VSUBS 0.036203f
C148 VN.n50 VSUBS 0.029373f
C149 VN.n51 VSUBS 0.036203f
C150 VN.t8 VSUBS 1.39678f
C151 VN.n52 VSUBS 0.53453f
C152 VN.n53 VSUBS 0.036203f
C153 VN.n54 VSUBS 0.02928f
C154 VN.n55 VSUBS 0.036203f
C155 VN.t7 VSUBS 1.39678f
C156 VN.n56 VSUBS 0.53453f
C157 VN.n57 VSUBS 0.036203f
C158 VN.n58 VSUBS 0.02928f
C159 VN.n59 VSUBS 0.036203f
C160 VN.t9 VSUBS 1.39678f
C161 VN.n60 VSUBS 0.652385f
C162 VN.t1 VSUBS 1.76937f
C163 VN.n61 VSUBS 0.628358f
C164 VN.n62 VSUBS 0.420838f
C165 VN.n63 VSUBS 0.050151f
C166 VN.n64 VSUBS 0.067474f
C167 VN.n65 VSUBS 0.072132f
C168 VN.n66 VSUBS 0.036203f
C169 VN.n67 VSUBS 0.036203f
C170 VN.n68 VSUBS 0.036203f
C171 VN.n69 VSUBS 0.071769f
C172 VN.n70 VSUBS 0.067474f
C173 VN.n71 VSUBS 0.050818f
C174 VN.n72 VSUBS 0.036203f
C175 VN.n73 VSUBS 0.036203f
C176 VN.n74 VSUBS 0.050818f
C177 VN.n75 VSUBS 0.067474f
C178 VN.n76 VSUBS 0.071769f
C179 VN.n77 VSUBS 0.036203f
C180 VN.n78 VSUBS 0.036203f
C181 VN.n79 VSUBS 0.036203f
C182 VN.n80 VSUBS 0.072132f
C183 VN.n81 VSUBS 0.067474f
C184 VN.n82 VSUBS 0.050151f
C185 VN.n83 VSUBS 0.036203f
C186 VN.n84 VSUBS 0.036203f
C187 VN.n85 VSUBS 0.051484f
C188 VN.n86 VSUBS 0.067474f
C189 VN.n87 VSUBS 0.071361f
C190 VN.n88 VSUBS 0.036203f
C191 VN.n89 VSUBS 0.036203f
C192 VN.n90 VSUBS 0.036203f
C193 VN.n91 VSUBS 0.072447f
C194 VN.n92 VSUBS 0.067474f
C195 VN.n93 VSUBS 0.049485f
C196 VN.n94 VSUBS 0.058431f
C197 VN.n95 VSUBS 2.11155f
C198 B.n0 VSUBS 0.011241f
C199 B.n1 VSUBS 0.011241f
C200 B.n2 VSUBS 0.016625f
C201 B.n3 VSUBS 0.01274f
C202 B.n4 VSUBS 0.01274f
C203 B.n5 VSUBS 0.01274f
C204 B.n6 VSUBS 0.01274f
C205 B.n7 VSUBS 0.01274f
C206 B.n8 VSUBS 0.01274f
C207 B.n9 VSUBS 0.01274f
C208 B.n10 VSUBS 0.01274f
C209 B.n11 VSUBS 0.01274f
C210 B.n12 VSUBS 0.01274f
C211 B.n13 VSUBS 0.01274f
C212 B.n14 VSUBS 0.01274f
C213 B.n15 VSUBS 0.01274f
C214 B.n16 VSUBS 0.01274f
C215 B.n17 VSUBS 0.01274f
C216 B.n18 VSUBS 0.01274f
C217 B.n19 VSUBS 0.01274f
C218 B.n20 VSUBS 0.01274f
C219 B.n21 VSUBS 0.01274f
C220 B.n22 VSUBS 0.01274f
C221 B.n23 VSUBS 0.01274f
C222 B.n24 VSUBS 0.01274f
C223 B.n25 VSUBS 0.01274f
C224 B.n26 VSUBS 0.01274f
C225 B.n27 VSUBS 0.01274f
C226 B.n28 VSUBS 0.01274f
C227 B.n29 VSUBS 0.01274f
C228 B.n30 VSUBS 0.01274f
C229 B.n31 VSUBS 0.01274f
C230 B.n32 VSUBS 0.01274f
C231 B.n33 VSUBS 0.01274f
C232 B.n34 VSUBS 0.01274f
C233 B.n35 VSUBS 0.01274f
C234 B.n36 VSUBS 0.029297f
C235 B.n37 VSUBS 0.01274f
C236 B.n38 VSUBS 0.01274f
C237 B.n39 VSUBS 0.01274f
C238 B.n40 VSUBS 0.01274f
C239 B.n41 VSUBS 0.01274f
C240 B.n42 VSUBS 0.01274f
C241 B.n43 VSUBS 0.01274f
C242 B.n44 VSUBS 0.01274f
C243 B.n45 VSUBS 0.01274f
C244 B.n46 VSUBS 0.011991f
C245 B.n47 VSUBS 0.01274f
C246 B.t7 VSUBS 0.124054f
C247 B.t8 VSUBS 0.172241f
C248 B.t6 VSUBS 1.29937f
C249 B.n48 VSUBS 0.292867f
C250 B.n49 VSUBS 0.241559f
C251 B.n50 VSUBS 0.029517f
C252 B.n51 VSUBS 0.01274f
C253 B.n52 VSUBS 0.01274f
C254 B.n53 VSUBS 0.01274f
C255 B.n54 VSUBS 0.01274f
C256 B.t1 VSUBS 0.124056f
C257 B.t2 VSUBS 0.172243f
C258 B.t0 VSUBS 1.29937f
C259 B.n55 VSUBS 0.292866f
C260 B.n56 VSUBS 0.241557f
C261 B.n57 VSUBS 0.01274f
C262 B.n58 VSUBS 0.01274f
C263 B.n59 VSUBS 0.01274f
C264 B.n60 VSUBS 0.01274f
C265 B.n61 VSUBS 0.01274f
C266 B.n62 VSUBS 0.01274f
C267 B.n63 VSUBS 0.01274f
C268 B.n64 VSUBS 0.01274f
C269 B.n65 VSUBS 0.01274f
C270 B.n66 VSUBS 0.031405f
C271 B.n67 VSUBS 0.01274f
C272 B.n68 VSUBS 0.01274f
C273 B.n69 VSUBS 0.01274f
C274 B.n70 VSUBS 0.01274f
C275 B.n71 VSUBS 0.01274f
C276 B.n72 VSUBS 0.01274f
C277 B.n73 VSUBS 0.01274f
C278 B.n74 VSUBS 0.01274f
C279 B.n75 VSUBS 0.01274f
C280 B.n76 VSUBS 0.01274f
C281 B.n77 VSUBS 0.01274f
C282 B.n78 VSUBS 0.01274f
C283 B.n79 VSUBS 0.01274f
C284 B.n80 VSUBS 0.01274f
C285 B.n81 VSUBS 0.01274f
C286 B.n82 VSUBS 0.01274f
C287 B.n83 VSUBS 0.01274f
C288 B.n84 VSUBS 0.01274f
C289 B.n85 VSUBS 0.01274f
C290 B.n86 VSUBS 0.01274f
C291 B.n87 VSUBS 0.01274f
C292 B.n88 VSUBS 0.01274f
C293 B.n89 VSUBS 0.01274f
C294 B.n90 VSUBS 0.01274f
C295 B.n91 VSUBS 0.01274f
C296 B.n92 VSUBS 0.01274f
C297 B.n93 VSUBS 0.01274f
C298 B.n94 VSUBS 0.01274f
C299 B.n95 VSUBS 0.01274f
C300 B.n96 VSUBS 0.01274f
C301 B.n97 VSUBS 0.01274f
C302 B.n98 VSUBS 0.01274f
C303 B.n99 VSUBS 0.01274f
C304 B.n100 VSUBS 0.01274f
C305 B.n101 VSUBS 0.01274f
C306 B.n102 VSUBS 0.01274f
C307 B.n103 VSUBS 0.01274f
C308 B.n104 VSUBS 0.01274f
C309 B.n105 VSUBS 0.01274f
C310 B.n106 VSUBS 0.01274f
C311 B.n107 VSUBS 0.01274f
C312 B.n108 VSUBS 0.01274f
C313 B.n109 VSUBS 0.01274f
C314 B.n110 VSUBS 0.01274f
C315 B.n111 VSUBS 0.01274f
C316 B.n112 VSUBS 0.01274f
C317 B.n113 VSUBS 0.01274f
C318 B.n114 VSUBS 0.01274f
C319 B.n115 VSUBS 0.01274f
C320 B.n116 VSUBS 0.01274f
C321 B.n117 VSUBS 0.01274f
C322 B.n118 VSUBS 0.01274f
C323 B.n119 VSUBS 0.01274f
C324 B.n120 VSUBS 0.01274f
C325 B.n121 VSUBS 0.01274f
C326 B.n122 VSUBS 0.01274f
C327 B.n123 VSUBS 0.01274f
C328 B.n124 VSUBS 0.01274f
C329 B.n125 VSUBS 0.01274f
C330 B.n126 VSUBS 0.01274f
C331 B.n127 VSUBS 0.01274f
C332 B.n128 VSUBS 0.01274f
C333 B.n129 VSUBS 0.01274f
C334 B.n130 VSUBS 0.01274f
C335 B.n131 VSUBS 0.01274f
C336 B.n132 VSUBS 0.01274f
C337 B.n133 VSUBS 0.01274f
C338 B.n134 VSUBS 0.01274f
C339 B.n135 VSUBS 0.01274f
C340 B.n136 VSUBS 0.029297f
C341 B.n137 VSUBS 0.01274f
C342 B.n138 VSUBS 0.01274f
C343 B.n139 VSUBS 0.01274f
C344 B.n140 VSUBS 0.01274f
C345 B.n141 VSUBS 0.01274f
C346 B.n142 VSUBS 0.01274f
C347 B.n143 VSUBS 0.01274f
C348 B.n144 VSUBS 0.01274f
C349 B.n145 VSUBS 0.01274f
C350 B.n146 VSUBS 0.01274f
C351 B.t11 VSUBS 0.124056f
C352 B.t10 VSUBS 0.172243f
C353 B.t9 VSUBS 1.29937f
C354 B.n147 VSUBS 0.292866f
C355 B.n148 VSUBS 0.241557f
C356 B.n149 VSUBS 0.01274f
C357 B.n150 VSUBS 0.01274f
C358 B.n151 VSUBS 0.01274f
C359 B.n152 VSUBS 0.01274f
C360 B.n153 VSUBS 0.007119f
C361 B.n154 VSUBS 0.01274f
C362 B.n155 VSUBS 0.01274f
C363 B.n156 VSUBS 0.01274f
C364 B.n157 VSUBS 0.01274f
C365 B.n158 VSUBS 0.01274f
C366 B.n159 VSUBS 0.01274f
C367 B.n160 VSUBS 0.01274f
C368 B.n161 VSUBS 0.01274f
C369 B.n162 VSUBS 0.01274f
C370 B.n163 VSUBS 0.031405f
C371 B.n164 VSUBS 0.01274f
C372 B.n165 VSUBS 0.01274f
C373 B.n166 VSUBS 0.01274f
C374 B.n167 VSUBS 0.01274f
C375 B.n168 VSUBS 0.01274f
C376 B.n169 VSUBS 0.01274f
C377 B.n170 VSUBS 0.01274f
C378 B.n171 VSUBS 0.01274f
C379 B.n172 VSUBS 0.01274f
C380 B.n173 VSUBS 0.01274f
C381 B.n174 VSUBS 0.01274f
C382 B.n175 VSUBS 0.01274f
C383 B.n176 VSUBS 0.01274f
C384 B.n177 VSUBS 0.01274f
C385 B.n178 VSUBS 0.01274f
C386 B.n179 VSUBS 0.01274f
C387 B.n180 VSUBS 0.01274f
C388 B.n181 VSUBS 0.01274f
C389 B.n182 VSUBS 0.01274f
C390 B.n183 VSUBS 0.01274f
C391 B.n184 VSUBS 0.01274f
C392 B.n185 VSUBS 0.01274f
C393 B.n186 VSUBS 0.01274f
C394 B.n187 VSUBS 0.01274f
C395 B.n188 VSUBS 0.01274f
C396 B.n189 VSUBS 0.01274f
C397 B.n190 VSUBS 0.01274f
C398 B.n191 VSUBS 0.01274f
C399 B.n192 VSUBS 0.01274f
C400 B.n193 VSUBS 0.01274f
C401 B.n194 VSUBS 0.01274f
C402 B.n195 VSUBS 0.01274f
C403 B.n196 VSUBS 0.01274f
C404 B.n197 VSUBS 0.01274f
C405 B.n198 VSUBS 0.01274f
C406 B.n199 VSUBS 0.01274f
C407 B.n200 VSUBS 0.01274f
C408 B.n201 VSUBS 0.01274f
C409 B.n202 VSUBS 0.01274f
C410 B.n203 VSUBS 0.01274f
C411 B.n204 VSUBS 0.01274f
C412 B.n205 VSUBS 0.01274f
C413 B.n206 VSUBS 0.01274f
C414 B.n207 VSUBS 0.01274f
C415 B.n208 VSUBS 0.01274f
C416 B.n209 VSUBS 0.01274f
C417 B.n210 VSUBS 0.01274f
C418 B.n211 VSUBS 0.01274f
C419 B.n212 VSUBS 0.01274f
C420 B.n213 VSUBS 0.01274f
C421 B.n214 VSUBS 0.01274f
C422 B.n215 VSUBS 0.01274f
C423 B.n216 VSUBS 0.01274f
C424 B.n217 VSUBS 0.01274f
C425 B.n218 VSUBS 0.01274f
C426 B.n219 VSUBS 0.01274f
C427 B.n220 VSUBS 0.01274f
C428 B.n221 VSUBS 0.01274f
C429 B.n222 VSUBS 0.01274f
C430 B.n223 VSUBS 0.01274f
C431 B.n224 VSUBS 0.01274f
C432 B.n225 VSUBS 0.01274f
C433 B.n226 VSUBS 0.01274f
C434 B.n227 VSUBS 0.01274f
C435 B.n228 VSUBS 0.01274f
C436 B.n229 VSUBS 0.01274f
C437 B.n230 VSUBS 0.01274f
C438 B.n231 VSUBS 0.01274f
C439 B.n232 VSUBS 0.01274f
C440 B.n233 VSUBS 0.01274f
C441 B.n234 VSUBS 0.01274f
C442 B.n235 VSUBS 0.01274f
C443 B.n236 VSUBS 0.01274f
C444 B.n237 VSUBS 0.01274f
C445 B.n238 VSUBS 0.01274f
C446 B.n239 VSUBS 0.01274f
C447 B.n240 VSUBS 0.01274f
C448 B.n241 VSUBS 0.01274f
C449 B.n242 VSUBS 0.01274f
C450 B.n243 VSUBS 0.01274f
C451 B.n244 VSUBS 0.01274f
C452 B.n245 VSUBS 0.01274f
C453 B.n246 VSUBS 0.01274f
C454 B.n247 VSUBS 0.01274f
C455 B.n248 VSUBS 0.01274f
C456 B.n249 VSUBS 0.01274f
C457 B.n250 VSUBS 0.01274f
C458 B.n251 VSUBS 0.01274f
C459 B.n252 VSUBS 0.01274f
C460 B.n253 VSUBS 0.01274f
C461 B.n254 VSUBS 0.01274f
C462 B.n255 VSUBS 0.01274f
C463 B.n256 VSUBS 0.01274f
C464 B.n257 VSUBS 0.01274f
C465 B.n258 VSUBS 0.01274f
C466 B.n259 VSUBS 0.01274f
C467 B.n260 VSUBS 0.01274f
C468 B.n261 VSUBS 0.01274f
C469 B.n262 VSUBS 0.01274f
C470 B.n263 VSUBS 0.01274f
C471 B.n264 VSUBS 0.01274f
C472 B.n265 VSUBS 0.01274f
C473 B.n266 VSUBS 0.01274f
C474 B.n267 VSUBS 0.01274f
C475 B.n268 VSUBS 0.01274f
C476 B.n269 VSUBS 0.01274f
C477 B.n270 VSUBS 0.01274f
C478 B.n271 VSUBS 0.01274f
C479 B.n272 VSUBS 0.01274f
C480 B.n273 VSUBS 0.01274f
C481 B.n274 VSUBS 0.01274f
C482 B.n275 VSUBS 0.01274f
C483 B.n276 VSUBS 0.01274f
C484 B.n277 VSUBS 0.01274f
C485 B.n278 VSUBS 0.01274f
C486 B.n279 VSUBS 0.01274f
C487 B.n280 VSUBS 0.01274f
C488 B.n281 VSUBS 0.01274f
C489 B.n282 VSUBS 0.01274f
C490 B.n283 VSUBS 0.01274f
C491 B.n284 VSUBS 0.01274f
C492 B.n285 VSUBS 0.01274f
C493 B.n286 VSUBS 0.01274f
C494 B.n287 VSUBS 0.01274f
C495 B.n288 VSUBS 0.01274f
C496 B.n289 VSUBS 0.01274f
C497 B.n290 VSUBS 0.01274f
C498 B.n291 VSUBS 0.01274f
C499 B.n292 VSUBS 0.01274f
C500 B.n293 VSUBS 0.01274f
C501 B.n294 VSUBS 0.01274f
C502 B.n295 VSUBS 0.01274f
C503 B.n296 VSUBS 0.01274f
C504 B.n297 VSUBS 0.01274f
C505 B.n298 VSUBS 0.029297f
C506 B.n299 VSUBS 0.029297f
C507 B.n300 VSUBS 0.031405f
C508 B.n301 VSUBS 0.01274f
C509 B.n302 VSUBS 0.01274f
C510 B.n303 VSUBS 0.01274f
C511 B.n304 VSUBS 0.01274f
C512 B.n305 VSUBS 0.01274f
C513 B.n306 VSUBS 0.01274f
C514 B.n307 VSUBS 0.01274f
C515 B.n308 VSUBS 0.01274f
C516 B.n309 VSUBS 0.01274f
C517 B.n310 VSUBS 0.01274f
C518 B.n311 VSUBS 0.01274f
C519 B.n312 VSUBS 0.01274f
C520 B.n313 VSUBS 0.01274f
C521 B.n314 VSUBS 0.01274f
C522 B.n315 VSUBS 0.01274f
C523 B.n316 VSUBS 0.01274f
C524 B.n317 VSUBS 0.01274f
C525 B.n318 VSUBS 0.01274f
C526 B.n319 VSUBS 0.01274f
C527 B.n320 VSUBS 0.01274f
C528 B.n321 VSUBS 0.01274f
C529 B.n322 VSUBS 0.01274f
C530 B.n323 VSUBS 0.01274f
C531 B.n324 VSUBS 0.01274f
C532 B.n325 VSUBS 0.01274f
C533 B.n326 VSUBS 0.01274f
C534 B.n327 VSUBS 0.01274f
C535 B.t5 VSUBS 0.124054f
C536 B.t4 VSUBS 0.172241f
C537 B.t3 VSUBS 1.29937f
C538 B.n328 VSUBS 0.292867f
C539 B.n329 VSUBS 0.241559f
C540 B.n330 VSUBS 0.029517f
C541 B.n331 VSUBS 0.011991f
C542 B.n332 VSUBS 0.01274f
C543 B.n333 VSUBS 0.01274f
C544 B.n334 VSUBS 0.01274f
C545 B.n335 VSUBS 0.01274f
C546 B.n336 VSUBS 0.01274f
C547 B.n337 VSUBS 0.01274f
C548 B.n338 VSUBS 0.01274f
C549 B.n339 VSUBS 0.01274f
C550 B.n340 VSUBS 0.01274f
C551 B.n341 VSUBS 0.01274f
C552 B.n342 VSUBS 0.01274f
C553 B.n343 VSUBS 0.01274f
C554 B.n344 VSUBS 0.01274f
C555 B.n345 VSUBS 0.01274f
C556 B.n346 VSUBS 0.01274f
C557 B.n347 VSUBS 0.007119f
C558 B.n348 VSUBS 0.029517f
C559 B.n349 VSUBS 0.011991f
C560 B.n350 VSUBS 0.01274f
C561 B.n351 VSUBS 0.01274f
C562 B.n352 VSUBS 0.01274f
C563 B.n353 VSUBS 0.01274f
C564 B.n354 VSUBS 0.01274f
C565 B.n355 VSUBS 0.01274f
C566 B.n356 VSUBS 0.01274f
C567 B.n357 VSUBS 0.01274f
C568 B.n358 VSUBS 0.01274f
C569 B.n359 VSUBS 0.01274f
C570 B.n360 VSUBS 0.01274f
C571 B.n361 VSUBS 0.01274f
C572 B.n362 VSUBS 0.01274f
C573 B.n363 VSUBS 0.01274f
C574 B.n364 VSUBS 0.01274f
C575 B.n365 VSUBS 0.01274f
C576 B.n366 VSUBS 0.01274f
C577 B.n367 VSUBS 0.01274f
C578 B.n368 VSUBS 0.01274f
C579 B.n369 VSUBS 0.01274f
C580 B.n370 VSUBS 0.01274f
C581 B.n371 VSUBS 0.01274f
C582 B.n372 VSUBS 0.01274f
C583 B.n373 VSUBS 0.01274f
C584 B.n374 VSUBS 0.01274f
C585 B.n375 VSUBS 0.01274f
C586 B.n376 VSUBS 0.01274f
C587 B.n377 VSUBS 0.031405f
C588 B.n378 VSUBS 0.02994f
C589 B.n379 VSUBS 0.030762f
C590 B.n380 VSUBS 0.01274f
C591 B.n381 VSUBS 0.01274f
C592 B.n382 VSUBS 0.01274f
C593 B.n383 VSUBS 0.01274f
C594 B.n384 VSUBS 0.01274f
C595 B.n385 VSUBS 0.01274f
C596 B.n386 VSUBS 0.01274f
C597 B.n387 VSUBS 0.01274f
C598 B.n388 VSUBS 0.01274f
C599 B.n389 VSUBS 0.01274f
C600 B.n390 VSUBS 0.01274f
C601 B.n391 VSUBS 0.01274f
C602 B.n392 VSUBS 0.01274f
C603 B.n393 VSUBS 0.01274f
C604 B.n394 VSUBS 0.01274f
C605 B.n395 VSUBS 0.01274f
C606 B.n396 VSUBS 0.01274f
C607 B.n397 VSUBS 0.01274f
C608 B.n398 VSUBS 0.01274f
C609 B.n399 VSUBS 0.01274f
C610 B.n400 VSUBS 0.01274f
C611 B.n401 VSUBS 0.01274f
C612 B.n402 VSUBS 0.01274f
C613 B.n403 VSUBS 0.01274f
C614 B.n404 VSUBS 0.01274f
C615 B.n405 VSUBS 0.01274f
C616 B.n406 VSUBS 0.01274f
C617 B.n407 VSUBS 0.01274f
C618 B.n408 VSUBS 0.01274f
C619 B.n409 VSUBS 0.01274f
C620 B.n410 VSUBS 0.01274f
C621 B.n411 VSUBS 0.01274f
C622 B.n412 VSUBS 0.01274f
C623 B.n413 VSUBS 0.01274f
C624 B.n414 VSUBS 0.01274f
C625 B.n415 VSUBS 0.01274f
C626 B.n416 VSUBS 0.01274f
C627 B.n417 VSUBS 0.01274f
C628 B.n418 VSUBS 0.01274f
C629 B.n419 VSUBS 0.01274f
C630 B.n420 VSUBS 0.01274f
C631 B.n421 VSUBS 0.01274f
C632 B.n422 VSUBS 0.01274f
C633 B.n423 VSUBS 0.01274f
C634 B.n424 VSUBS 0.01274f
C635 B.n425 VSUBS 0.01274f
C636 B.n426 VSUBS 0.01274f
C637 B.n427 VSUBS 0.01274f
C638 B.n428 VSUBS 0.01274f
C639 B.n429 VSUBS 0.01274f
C640 B.n430 VSUBS 0.01274f
C641 B.n431 VSUBS 0.01274f
C642 B.n432 VSUBS 0.01274f
C643 B.n433 VSUBS 0.01274f
C644 B.n434 VSUBS 0.01274f
C645 B.n435 VSUBS 0.01274f
C646 B.n436 VSUBS 0.01274f
C647 B.n437 VSUBS 0.01274f
C648 B.n438 VSUBS 0.01274f
C649 B.n439 VSUBS 0.01274f
C650 B.n440 VSUBS 0.01274f
C651 B.n441 VSUBS 0.01274f
C652 B.n442 VSUBS 0.01274f
C653 B.n443 VSUBS 0.01274f
C654 B.n444 VSUBS 0.01274f
C655 B.n445 VSUBS 0.01274f
C656 B.n446 VSUBS 0.01274f
C657 B.n447 VSUBS 0.01274f
C658 B.n448 VSUBS 0.01274f
C659 B.n449 VSUBS 0.01274f
C660 B.n450 VSUBS 0.01274f
C661 B.n451 VSUBS 0.01274f
C662 B.n452 VSUBS 0.01274f
C663 B.n453 VSUBS 0.01274f
C664 B.n454 VSUBS 0.01274f
C665 B.n455 VSUBS 0.01274f
C666 B.n456 VSUBS 0.01274f
C667 B.n457 VSUBS 0.01274f
C668 B.n458 VSUBS 0.01274f
C669 B.n459 VSUBS 0.01274f
C670 B.n460 VSUBS 0.01274f
C671 B.n461 VSUBS 0.01274f
C672 B.n462 VSUBS 0.01274f
C673 B.n463 VSUBS 0.01274f
C674 B.n464 VSUBS 0.01274f
C675 B.n465 VSUBS 0.01274f
C676 B.n466 VSUBS 0.01274f
C677 B.n467 VSUBS 0.01274f
C678 B.n468 VSUBS 0.01274f
C679 B.n469 VSUBS 0.01274f
C680 B.n470 VSUBS 0.01274f
C681 B.n471 VSUBS 0.01274f
C682 B.n472 VSUBS 0.01274f
C683 B.n473 VSUBS 0.01274f
C684 B.n474 VSUBS 0.01274f
C685 B.n475 VSUBS 0.01274f
C686 B.n476 VSUBS 0.01274f
C687 B.n477 VSUBS 0.01274f
C688 B.n478 VSUBS 0.01274f
C689 B.n479 VSUBS 0.01274f
C690 B.n480 VSUBS 0.01274f
C691 B.n481 VSUBS 0.01274f
C692 B.n482 VSUBS 0.01274f
C693 B.n483 VSUBS 0.01274f
C694 B.n484 VSUBS 0.01274f
C695 B.n485 VSUBS 0.01274f
C696 B.n486 VSUBS 0.01274f
C697 B.n487 VSUBS 0.01274f
C698 B.n488 VSUBS 0.01274f
C699 B.n489 VSUBS 0.01274f
C700 B.n490 VSUBS 0.01274f
C701 B.n491 VSUBS 0.01274f
C702 B.n492 VSUBS 0.01274f
C703 B.n493 VSUBS 0.01274f
C704 B.n494 VSUBS 0.01274f
C705 B.n495 VSUBS 0.01274f
C706 B.n496 VSUBS 0.01274f
C707 B.n497 VSUBS 0.01274f
C708 B.n498 VSUBS 0.01274f
C709 B.n499 VSUBS 0.01274f
C710 B.n500 VSUBS 0.01274f
C711 B.n501 VSUBS 0.01274f
C712 B.n502 VSUBS 0.01274f
C713 B.n503 VSUBS 0.01274f
C714 B.n504 VSUBS 0.01274f
C715 B.n505 VSUBS 0.01274f
C716 B.n506 VSUBS 0.01274f
C717 B.n507 VSUBS 0.01274f
C718 B.n508 VSUBS 0.01274f
C719 B.n509 VSUBS 0.01274f
C720 B.n510 VSUBS 0.01274f
C721 B.n511 VSUBS 0.01274f
C722 B.n512 VSUBS 0.01274f
C723 B.n513 VSUBS 0.01274f
C724 B.n514 VSUBS 0.01274f
C725 B.n515 VSUBS 0.01274f
C726 B.n516 VSUBS 0.01274f
C727 B.n517 VSUBS 0.01274f
C728 B.n518 VSUBS 0.01274f
C729 B.n519 VSUBS 0.01274f
C730 B.n520 VSUBS 0.01274f
C731 B.n521 VSUBS 0.01274f
C732 B.n522 VSUBS 0.01274f
C733 B.n523 VSUBS 0.01274f
C734 B.n524 VSUBS 0.01274f
C735 B.n525 VSUBS 0.01274f
C736 B.n526 VSUBS 0.01274f
C737 B.n527 VSUBS 0.01274f
C738 B.n528 VSUBS 0.01274f
C739 B.n529 VSUBS 0.01274f
C740 B.n530 VSUBS 0.01274f
C741 B.n531 VSUBS 0.01274f
C742 B.n532 VSUBS 0.01274f
C743 B.n533 VSUBS 0.01274f
C744 B.n534 VSUBS 0.01274f
C745 B.n535 VSUBS 0.01274f
C746 B.n536 VSUBS 0.01274f
C747 B.n537 VSUBS 0.01274f
C748 B.n538 VSUBS 0.01274f
C749 B.n539 VSUBS 0.01274f
C750 B.n540 VSUBS 0.01274f
C751 B.n541 VSUBS 0.01274f
C752 B.n542 VSUBS 0.01274f
C753 B.n543 VSUBS 0.01274f
C754 B.n544 VSUBS 0.01274f
C755 B.n545 VSUBS 0.01274f
C756 B.n546 VSUBS 0.01274f
C757 B.n547 VSUBS 0.01274f
C758 B.n548 VSUBS 0.01274f
C759 B.n549 VSUBS 0.01274f
C760 B.n550 VSUBS 0.01274f
C761 B.n551 VSUBS 0.01274f
C762 B.n552 VSUBS 0.01274f
C763 B.n553 VSUBS 0.01274f
C764 B.n554 VSUBS 0.01274f
C765 B.n555 VSUBS 0.01274f
C766 B.n556 VSUBS 0.01274f
C767 B.n557 VSUBS 0.01274f
C768 B.n558 VSUBS 0.01274f
C769 B.n559 VSUBS 0.01274f
C770 B.n560 VSUBS 0.01274f
C771 B.n561 VSUBS 0.01274f
C772 B.n562 VSUBS 0.01274f
C773 B.n563 VSUBS 0.01274f
C774 B.n564 VSUBS 0.01274f
C775 B.n565 VSUBS 0.01274f
C776 B.n566 VSUBS 0.01274f
C777 B.n567 VSUBS 0.01274f
C778 B.n568 VSUBS 0.01274f
C779 B.n569 VSUBS 0.01274f
C780 B.n570 VSUBS 0.01274f
C781 B.n571 VSUBS 0.01274f
C782 B.n572 VSUBS 0.01274f
C783 B.n573 VSUBS 0.01274f
C784 B.n574 VSUBS 0.01274f
C785 B.n575 VSUBS 0.01274f
C786 B.n576 VSUBS 0.01274f
C787 B.n577 VSUBS 0.01274f
C788 B.n578 VSUBS 0.01274f
C789 B.n579 VSUBS 0.01274f
C790 B.n580 VSUBS 0.01274f
C791 B.n581 VSUBS 0.01274f
C792 B.n582 VSUBS 0.01274f
C793 B.n583 VSUBS 0.01274f
C794 B.n584 VSUBS 0.01274f
C795 B.n585 VSUBS 0.01274f
C796 B.n586 VSUBS 0.01274f
C797 B.n587 VSUBS 0.029297f
C798 B.n588 VSUBS 0.029297f
C799 B.n589 VSUBS 0.031405f
C800 B.n590 VSUBS 0.01274f
C801 B.n591 VSUBS 0.01274f
C802 B.n592 VSUBS 0.01274f
C803 B.n593 VSUBS 0.01274f
C804 B.n594 VSUBS 0.01274f
C805 B.n595 VSUBS 0.01274f
C806 B.n596 VSUBS 0.01274f
C807 B.n597 VSUBS 0.01274f
C808 B.n598 VSUBS 0.01274f
C809 B.n599 VSUBS 0.01274f
C810 B.n600 VSUBS 0.01274f
C811 B.n601 VSUBS 0.01274f
C812 B.n602 VSUBS 0.01274f
C813 B.n603 VSUBS 0.01274f
C814 B.n604 VSUBS 0.01274f
C815 B.n605 VSUBS 0.01274f
C816 B.n606 VSUBS 0.01274f
C817 B.n607 VSUBS 0.01274f
C818 B.n608 VSUBS 0.01274f
C819 B.n609 VSUBS 0.01274f
C820 B.n610 VSUBS 0.01274f
C821 B.n611 VSUBS 0.01274f
C822 B.n612 VSUBS 0.01274f
C823 B.n613 VSUBS 0.01274f
C824 B.n614 VSUBS 0.01274f
C825 B.n615 VSUBS 0.01274f
C826 B.n616 VSUBS 0.01274f
C827 B.n617 VSUBS 0.01274f
C828 B.n618 VSUBS 0.011991f
C829 B.n619 VSUBS 0.029517f
C830 B.n620 VSUBS 0.007119f
C831 B.n621 VSUBS 0.01274f
C832 B.n622 VSUBS 0.01274f
C833 B.n623 VSUBS 0.01274f
C834 B.n624 VSUBS 0.01274f
C835 B.n625 VSUBS 0.01274f
C836 B.n626 VSUBS 0.01274f
C837 B.n627 VSUBS 0.01274f
C838 B.n628 VSUBS 0.01274f
C839 B.n629 VSUBS 0.01274f
C840 B.n630 VSUBS 0.01274f
C841 B.n631 VSUBS 0.01274f
C842 B.n632 VSUBS 0.01274f
C843 B.n633 VSUBS 0.007119f
C844 B.n634 VSUBS 0.01274f
C845 B.n635 VSUBS 0.01274f
C846 B.n636 VSUBS 0.01274f
C847 B.n637 VSUBS 0.01274f
C848 B.n638 VSUBS 0.01274f
C849 B.n639 VSUBS 0.01274f
C850 B.n640 VSUBS 0.01274f
C851 B.n641 VSUBS 0.01274f
C852 B.n642 VSUBS 0.01274f
C853 B.n643 VSUBS 0.01274f
C854 B.n644 VSUBS 0.01274f
C855 B.n645 VSUBS 0.01274f
C856 B.n646 VSUBS 0.01274f
C857 B.n647 VSUBS 0.01274f
C858 B.n648 VSUBS 0.01274f
C859 B.n649 VSUBS 0.01274f
C860 B.n650 VSUBS 0.01274f
C861 B.n651 VSUBS 0.01274f
C862 B.n652 VSUBS 0.01274f
C863 B.n653 VSUBS 0.01274f
C864 B.n654 VSUBS 0.01274f
C865 B.n655 VSUBS 0.01274f
C866 B.n656 VSUBS 0.01274f
C867 B.n657 VSUBS 0.01274f
C868 B.n658 VSUBS 0.01274f
C869 B.n659 VSUBS 0.01274f
C870 B.n660 VSUBS 0.01274f
C871 B.n661 VSUBS 0.01274f
C872 B.n662 VSUBS 0.01274f
C873 B.n663 VSUBS 0.031405f
C874 B.n664 VSUBS 0.031405f
C875 B.n665 VSUBS 0.029297f
C876 B.n666 VSUBS 0.01274f
C877 B.n667 VSUBS 0.01274f
C878 B.n668 VSUBS 0.01274f
C879 B.n669 VSUBS 0.01274f
C880 B.n670 VSUBS 0.01274f
C881 B.n671 VSUBS 0.01274f
C882 B.n672 VSUBS 0.01274f
C883 B.n673 VSUBS 0.01274f
C884 B.n674 VSUBS 0.01274f
C885 B.n675 VSUBS 0.01274f
C886 B.n676 VSUBS 0.01274f
C887 B.n677 VSUBS 0.01274f
C888 B.n678 VSUBS 0.01274f
C889 B.n679 VSUBS 0.01274f
C890 B.n680 VSUBS 0.01274f
C891 B.n681 VSUBS 0.01274f
C892 B.n682 VSUBS 0.01274f
C893 B.n683 VSUBS 0.01274f
C894 B.n684 VSUBS 0.01274f
C895 B.n685 VSUBS 0.01274f
C896 B.n686 VSUBS 0.01274f
C897 B.n687 VSUBS 0.01274f
C898 B.n688 VSUBS 0.01274f
C899 B.n689 VSUBS 0.01274f
C900 B.n690 VSUBS 0.01274f
C901 B.n691 VSUBS 0.01274f
C902 B.n692 VSUBS 0.01274f
C903 B.n693 VSUBS 0.01274f
C904 B.n694 VSUBS 0.01274f
C905 B.n695 VSUBS 0.01274f
C906 B.n696 VSUBS 0.01274f
C907 B.n697 VSUBS 0.01274f
C908 B.n698 VSUBS 0.01274f
C909 B.n699 VSUBS 0.01274f
C910 B.n700 VSUBS 0.01274f
C911 B.n701 VSUBS 0.01274f
C912 B.n702 VSUBS 0.01274f
C913 B.n703 VSUBS 0.01274f
C914 B.n704 VSUBS 0.01274f
C915 B.n705 VSUBS 0.01274f
C916 B.n706 VSUBS 0.01274f
C917 B.n707 VSUBS 0.01274f
C918 B.n708 VSUBS 0.01274f
C919 B.n709 VSUBS 0.01274f
C920 B.n710 VSUBS 0.01274f
C921 B.n711 VSUBS 0.01274f
C922 B.n712 VSUBS 0.01274f
C923 B.n713 VSUBS 0.01274f
C924 B.n714 VSUBS 0.01274f
C925 B.n715 VSUBS 0.01274f
C926 B.n716 VSUBS 0.01274f
C927 B.n717 VSUBS 0.01274f
C928 B.n718 VSUBS 0.01274f
C929 B.n719 VSUBS 0.01274f
C930 B.n720 VSUBS 0.01274f
C931 B.n721 VSUBS 0.01274f
C932 B.n722 VSUBS 0.01274f
C933 B.n723 VSUBS 0.01274f
C934 B.n724 VSUBS 0.01274f
C935 B.n725 VSUBS 0.01274f
C936 B.n726 VSUBS 0.01274f
C937 B.n727 VSUBS 0.01274f
C938 B.n728 VSUBS 0.01274f
C939 B.n729 VSUBS 0.01274f
C940 B.n730 VSUBS 0.01274f
C941 B.n731 VSUBS 0.01274f
C942 B.n732 VSUBS 0.01274f
C943 B.n733 VSUBS 0.01274f
C944 B.n734 VSUBS 0.01274f
C945 B.n735 VSUBS 0.01274f
C946 B.n736 VSUBS 0.01274f
C947 B.n737 VSUBS 0.01274f
C948 B.n738 VSUBS 0.01274f
C949 B.n739 VSUBS 0.01274f
C950 B.n740 VSUBS 0.01274f
C951 B.n741 VSUBS 0.01274f
C952 B.n742 VSUBS 0.01274f
C953 B.n743 VSUBS 0.01274f
C954 B.n744 VSUBS 0.01274f
C955 B.n745 VSUBS 0.01274f
C956 B.n746 VSUBS 0.01274f
C957 B.n747 VSUBS 0.01274f
C958 B.n748 VSUBS 0.01274f
C959 B.n749 VSUBS 0.01274f
C960 B.n750 VSUBS 0.01274f
C961 B.n751 VSUBS 0.01274f
C962 B.n752 VSUBS 0.01274f
C963 B.n753 VSUBS 0.01274f
C964 B.n754 VSUBS 0.01274f
C965 B.n755 VSUBS 0.01274f
C966 B.n756 VSUBS 0.01274f
C967 B.n757 VSUBS 0.01274f
C968 B.n758 VSUBS 0.01274f
C969 B.n759 VSUBS 0.01274f
C970 B.n760 VSUBS 0.01274f
C971 B.n761 VSUBS 0.01274f
C972 B.n762 VSUBS 0.01274f
C973 B.n763 VSUBS 0.01274f
C974 B.n764 VSUBS 0.01274f
C975 B.n765 VSUBS 0.01274f
C976 B.n766 VSUBS 0.01274f
C977 B.n767 VSUBS 0.016625f
C978 B.n768 VSUBS 0.01771f
C979 B.n769 VSUBS 0.035218f
C980 VTAIL.t9 VSUBS 0.133999f
C981 VTAIL.t6 VSUBS 0.133999f
C982 VTAIL.n0 VSUBS 0.727845f
C983 VTAIL.n1 VSUBS 1.08968f
C984 VTAIL.n2 VSUBS 0.040342f
C985 VTAIL.n3 VSUBS 0.036155f
C986 VTAIL.n4 VSUBS 0.019428f
C987 VTAIL.n5 VSUBS 0.045922f
C988 VTAIL.n6 VSUBS 0.020571f
C989 VTAIL.n7 VSUBS 0.610752f
C990 VTAIL.n8 VSUBS 0.019428f
C991 VTAIL.t16 VSUBS 0.100458f
C992 VTAIL.n9 VSUBS 0.147568f
C993 VTAIL.n10 VSUBS 0.029092f
C994 VTAIL.n11 VSUBS 0.034441f
C995 VTAIL.n12 VSUBS 0.045922f
C996 VTAIL.n13 VSUBS 0.020571f
C997 VTAIL.n14 VSUBS 0.019428f
C998 VTAIL.n15 VSUBS 0.036155f
C999 VTAIL.n16 VSUBS 0.036155f
C1000 VTAIL.n17 VSUBS 0.019428f
C1001 VTAIL.n18 VSUBS 0.020571f
C1002 VTAIL.n19 VSUBS 0.045922f
C1003 VTAIL.n20 VSUBS 0.113267f
C1004 VTAIL.n21 VSUBS 0.020571f
C1005 VTAIL.n22 VSUBS 0.019428f
C1006 VTAIL.n23 VSUBS 0.089993f
C1007 VTAIL.n24 VSUBS 0.057245f
C1008 VTAIL.n25 VSUBS 0.615006f
C1009 VTAIL.t18 VSUBS 0.133999f
C1010 VTAIL.t19 VSUBS 0.133999f
C1011 VTAIL.n26 VSUBS 0.727845f
C1012 VTAIL.n27 VSUBS 1.29104f
C1013 VTAIL.t12 VSUBS 0.133999f
C1014 VTAIL.t10 VSUBS 0.133999f
C1015 VTAIL.n28 VSUBS 0.727845f
C1016 VTAIL.n29 VSUBS 2.60371f
C1017 VTAIL.t7 VSUBS 0.133999f
C1018 VTAIL.t0 VSUBS 0.133999f
C1019 VTAIL.n30 VSUBS 0.72785f
C1020 VTAIL.n31 VSUBS 2.6037f
C1021 VTAIL.t3 VSUBS 0.133999f
C1022 VTAIL.t1 VSUBS 0.133999f
C1023 VTAIL.n32 VSUBS 0.72785f
C1024 VTAIL.n33 VSUBS 1.29104f
C1025 VTAIL.n34 VSUBS 0.040342f
C1026 VTAIL.n35 VSUBS 0.036155f
C1027 VTAIL.n36 VSUBS 0.019428f
C1028 VTAIL.n37 VSUBS 0.045922f
C1029 VTAIL.n38 VSUBS 0.020571f
C1030 VTAIL.n39 VSUBS 0.610752f
C1031 VTAIL.n40 VSUBS 0.019428f
C1032 VTAIL.t8 VSUBS 0.100458f
C1033 VTAIL.n41 VSUBS 0.147568f
C1034 VTAIL.n42 VSUBS 0.029092f
C1035 VTAIL.n43 VSUBS 0.034441f
C1036 VTAIL.n44 VSUBS 0.045922f
C1037 VTAIL.n45 VSUBS 0.020571f
C1038 VTAIL.n46 VSUBS 0.019428f
C1039 VTAIL.n47 VSUBS 0.036155f
C1040 VTAIL.n48 VSUBS 0.036155f
C1041 VTAIL.n49 VSUBS 0.019428f
C1042 VTAIL.n50 VSUBS 0.020571f
C1043 VTAIL.n51 VSUBS 0.045922f
C1044 VTAIL.n52 VSUBS 0.113267f
C1045 VTAIL.n53 VSUBS 0.020571f
C1046 VTAIL.n54 VSUBS 0.019428f
C1047 VTAIL.n55 VSUBS 0.089993f
C1048 VTAIL.n56 VSUBS 0.057245f
C1049 VTAIL.n57 VSUBS 0.615006f
C1050 VTAIL.t17 VSUBS 0.133999f
C1051 VTAIL.t14 VSUBS 0.133999f
C1052 VTAIL.n58 VSUBS 0.72785f
C1053 VTAIL.n59 VSUBS 1.17052f
C1054 VTAIL.t11 VSUBS 0.133999f
C1055 VTAIL.t15 VSUBS 0.133999f
C1056 VTAIL.n60 VSUBS 0.72785f
C1057 VTAIL.n61 VSUBS 1.29104f
C1058 VTAIL.n62 VSUBS 0.040342f
C1059 VTAIL.n63 VSUBS 0.036155f
C1060 VTAIL.n64 VSUBS 0.019428f
C1061 VTAIL.n65 VSUBS 0.045922f
C1062 VTAIL.n66 VSUBS 0.020571f
C1063 VTAIL.n67 VSUBS 0.610752f
C1064 VTAIL.n68 VSUBS 0.019428f
C1065 VTAIL.t13 VSUBS 0.100458f
C1066 VTAIL.n69 VSUBS 0.147568f
C1067 VTAIL.n70 VSUBS 0.029092f
C1068 VTAIL.n71 VSUBS 0.034441f
C1069 VTAIL.n72 VSUBS 0.045922f
C1070 VTAIL.n73 VSUBS 0.020571f
C1071 VTAIL.n74 VSUBS 0.019428f
C1072 VTAIL.n75 VSUBS 0.036155f
C1073 VTAIL.n76 VSUBS 0.036155f
C1074 VTAIL.n77 VSUBS 0.019428f
C1075 VTAIL.n78 VSUBS 0.020571f
C1076 VTAIL.n79 VSUBS 0.045922f
C1077 VTAIL.n80 VSUBS 0.113267f
C1078 VTAIL.n81 VSUBS 0.020571f
C1079 VTAIL.n82 VSUBS 0.019428f
C1080 VTAIL.n83 VSUBS 0.089993f
C1081 VTAIL.n84 VSUBS 0.057245f
C1082 VTAIL.n85 VSUBS 1.69768f
C1083 VTAIL.n86 VSUBS 0.040342f
C1084 VTAIL.n87 VSUBS 0.036155f
C1085 VTAIL.n88 VSUBS 0.019428f
C1086 VTAIL.n89 VSUBS 0.045922f
C1087 VTAIL.n90 VSUBS 0.020571f
C1088 VTAIL.n91 VSUBS 0.610752f
C1089 VTAIL.n92 VSUBS 0.019428f
C1090 VTAIL.t2 VSUBS 0.100458f
C1091 VTAIL.n93 VSUBS 0.147568f
C1092 VTAIL.n94 VSUBS 0.029092f
C1093 VTAIL.n95 VSUBS 0.034441f
C1094 VTAIL.n96 VSUBS 0.045922f
C1095 VTAIL.n97 VSUBS 0.020571f
C1096 VTAIL.n98 VSUBS 0.019428f
C1097 VTAIL.n99 VSUBS 0.036155f
C1098 VTAIL.n100 VSUBS 0.036155f
C1099 VTAIL.n101 VSUBS 0.019428f
C1100 VTAIL.n102 VSUBS 0.020571f
C1101 VTAIL.n103 VSUBS 0.045922f
C1102 VTAIL.n104 VSUBS 0.113267f
C1103 VTAIL.n105 VSUBS 0.020571f
C1104 VTAIL.n106 VSUBS 0.019428f
C1105 VTAIL.n107 VSUBS 0.089993f
C1106 VTAIL.n108 VSUBS 0.057245f
C1107 VTAIL.n109 VSUBS 1.69768f
C1108 VTAIL.t5 VSUBS 0.133999f
C1109 VTAIL.t4 VSUBS 0.133999f
C1110 VTAIL.n110 VSUBS 0.727845f
C1111 VTAIL.n111 VSUBS 1.02138f
C1112 VDD1.n0 VSUBS 0.040583f
C1113 VDD1.n1 VSUBS 0.036371f
C1114 VDD1.n2 VSUBS 0.019544f
C1115 VDD1.n3 VSUBS 0.046195f
C1116 VDD1.n4 VSUBS 0.020694f
C1117 VDD1.n5 VSUBS 0.614391f
C1118 VDD1.n6 VSUBS 0.019544f
C1119 VDD1.t6 VSUBS 0.101056f
C1120 VDD1.n7 VSUBS 0.148447f
C1121 VDD1.n8 VSUBS 0.029265f
C1122 VDD1.n9 VSUBS 0.034646f
C1123 VDD1.n10 VSUBS 0.046195f
C1124 VDD1.n11 VSUBS 0.020694f
C1125 VDD1.n12 VSUBS 0.019544f
C1126 VDD1.n13 VSUBS 0.036371f
C1127 VDD1.n14 VSUBS 0.036371f
C1128 VDD1.n15 VSUBS 0.019544f
C1129 VDD1.n16 VSUBS 0.020694f
C1130 VDD1.n17 VSUBS 0.046195f
C1131 VDD1.n18 VSUBS 0.113941f
C1132 VDD1.n19 VSUBS 0.020694f
C1133 VDD1.n20 VSUBS 0.019544f
C1134 VDD1.n21 VSUBS 0.090529f
C1135 VDD1.n22 VSUBS 0.106233f
C1136 VDD1.t7 VSUBS 0.134797f
C1137 VDD1.t5 VSUBS 0.134797f
C1138 VDD1.n23 VSUBS 0.831703f
C1139 VDD1.n24 VSUBS 1.39377f
C1140 VDD1.n25 VSUBS 0.040583f
C1141 VDD1.n26 VSUBS 0.036371f
C1142 VDD1.n27 VSUBS 0.019544f
C1143 VDD1.n28 VSUBS 0.046195f
C1144 VDD1.n29 VSUBS 0.020694f
C1145 VDD1.n30 VSUBS 0.614391f
C1146 VDD1.n31 VSUBS 0.019544f
C1147 VDD1.t8 VSUBS 0.101056f
C1148 VDD1.n32 VSUBS 0.148447f
C1149 VDD1.n33 VSUBS 0.029265f
C1150 VDD1.n34 VSUBS 0.034646f
C1151 VDD1.n35 VSUBS 0.046195f
C1152 VDD1.n36 VSUBS 0.020694f
C1153 VDD1.n37 VSUBS 0.019544f
C1154 VDD1.n38 VSUBS 0.036371f
C1155 VDD1.n39 VSUBS 0.036371f
C1156 VDD1.n40 VSUBS 0.019544f
C1157 VDD1.n41 VSUBS 0.020694f
C1158 VDD1.n42 VSUBS 0.046195f
C1159 VDD1.n43 VSUBS 0.113941f
C1160 VDD1.n44 VSUBS 0.020694f
C1161 VDD1.n45 VSUBS 0.019544f
C1162 VDD1.n46 VSUBS 0.090529f
C1163 VDD1.n47 VSUBS 0.106233f
C1164 VDD1.t1 VSUBS 0.134797f
C1165 VDD1.t2 VSUBS 0.134797f
C1166 VDD1.n48 VSUBS 0.831699f
C1167 VDD1.n49 VSUBS 1.38168f
C1168 VDD1.t3 VSUBS 0.134797f
C1169 VDD1.t4 VSUBS 0.134797f
C1170 VDD1.n50 VSUBS 0.85535f
C1171 VDD1.n51 VSUBS 4.44867f
C1172 VDD1.t0 VSUBS 0.134797f
C1173 VDD1.t9 VSUBS 0.134797f
C1174 VDD1.n52 VSUBS 0.831699f
C1175 VDD1.n53 VSUBS 4.37988f
C1176 VP.t3 VSUBS 1.57759f
C1177 VP.n0 VSUBS 0.750164f
C1178 VP.n1 VSUBS 0.04089f
C1179 VP.n2 VSUBS 0.033175f
C1180 VP.n3 VSUBS 0.04089f
C1181 VP.t0 VSUBS 1.57759f
C1182 VP.n4 VSUBS 0.603723f
C1183 VP.n5 VSUBS 0.04089f
C1184 VP.n6 VSUBS 0.03307f
C1185 VP.n7 VSUBS 0.04089f
C1186 VP.t1 VSUBS 1.57759f
C1187 VP.n8 VSUBS 0.603723f
C1188 VP.n9 VSUBS 0.04089f
C1189 VP.n10 VSUBS 0.03307f
C1190 VP.n11 VSUBS 0.04089f
C1191 VP.t9 VSUBS 1.57759f
C1192 VP.n12 VSUBS 0.603723f
C1193 VP.n13 VSUBS 0.04089f
C1194 VP.n14 VSUBS 0.033175f
C1195 VP.n15 VSUBS 0.04089f
C1196 VP.t7 VSUBS 1.57759f
C1197 VP.n16 VSUBS 0.750164f
C1198 VP.t6 VSUBS 1.57759f
C1199 VP.n17 VSUBS 0.750164f
C1200 VP.n18 VSUBS 0.04089f
C1201 VP.n19 VSUBS 0.033175f
C1202 VP.n20 VSUBS 0.04089f
C1203 VP.t4 VSUBS 1.57759f
C1204 VP.n21 VSUBS 0.603723f
C1205 VP.n22 VSUBS 0.04089f
C1206 VP.n23 VSUBS 0.03307f
C1207 VP.n24 VSUBS 0.04089f
C1208 VP.t8 VSUBS 1.57759f
C1209 VP.n25 VSUBS 0.603723f
C1210 VP.n26 VSUBS 0.04089f
C1211 VP.n27 VSUBS 0.03307f
C1212 VP.n28 VSUBS 0.04089f
C1213 VP.t5 VSUBS 1.57759f
C1214 VP.n29 VSUBS 0.736834f
C1215 VP.t2 VSUBS 1.9984f
C1216 VP.n30 VSUBS 0.709697f
C1217 VP.n31 VSUBS 0.475315f
C1218 VP.n32 VSUBS 0.056643f
C1219 VP.n33 VSUBS 0.076208f
C1220 VP.n34 VSUBS 0.081469f
C1221 VP.n35 VSUBS 0.04089f
C1222 VP.n36 VSUBS 0.04089f
C1223 VP.n37 VSUBS 0.04089f
C1224 VP.n38 VSUBS 0.081059f
C1225 VP.n39 VSUBS 0.076208f
C1226 VP.n40 VSUBS 0.057396f
C1227 VP.n41 VSUBS 0.04089f
C1228 VP.n42 VSUBS 0.04089f
C1229 VP.n43 VSUBS 0.057396f
C1230 VP.n44 VSUBS 0.076208f
C1231 VP.n45 VSUBS 0.081059f
C1232 VP.n46 VSUBS 0.04089f
C1233 VP.n47 VSUBS 0.04089f
C1234 VP.n48 VSUBS 0.04089f
C1235 VP.n49 VSUBS 0.081469f
C1236 VP.n50 VSUBS 0.076208f
C1237 VP.n51 VSUBS 0.056643f
C1238 VP.n52 VSUBS 0.04089f
C1239 VP.n53 VSUBS 0.04089f
C1240 VP.n54 VSUBS 0.058148f
C1241 VP.n55 VSUBS 0.076208f
C1242 VP.n56 VSUBS 0.080598f
C1243 VP.n57 VSUBS 0.04089f
C1244 VP.n58 VSUBS 0.04089f
C1245 VP.n59 VSUBS 0.04089f
C1246 VP.n60 VSUBS 0.081825f
C1247 VP.n61 VSUBS 0.076208f
C1248 VP.n62 VSUBS 0.055891f
C1249 VP.n63 VSUBS 0.065995f
C1250 VP.n64 VSUBS 2.3682f
C1251 VP.n65 VSUBS 2.39723f
C1252 VP.n66 VSUBS 0.065995f
C1253 VP.n67 VSUBS 0.055891f
C1254 VP.n68 VSUBS 0.076208f
C1255 VP.n69 VSUBS 0.081825f
C1256 VP.n70 VSUBS 0.04089f
C1257 VP.n71 VSUBS 0.04089f
C1258 VP.n72 VSUBS 0.04089f
C1259 VP.n73 VSUBS 0.080598f
C1260 VP.n74 VSUBS 0.076208f
C1261 VP.n75 VSUBS 0.058148f
C1262 VP.n76 VSUBS 0.04089f
C1263 VP.n77 VSUBS 0.04089f
C1264 VP.n78 VSUBS 0.056643f
C1265 VP.n79 VSUBS 0.076208f
C1266 VP.n80 VSUBS 0.081469f
C1267 VP.n81 VSUBS 0.04089f
C1268 VP.n82 VSUBS 0.04089f
C1269 VP.n83 VSUBS 0.04089f
C1270 VP.n84 VSUBS 0.081059f
C1271 VP.n85 VSUBS 0.076208f
C1272 VP.n86 VSUBS 0.057396f
C1273 VP.n87 VSUBS 0.04089f
C1274 VP.n88 VSUBS 0.04089f
C1275 VP.n89 VSUBS 0.057396f
C1276 VP.n90 VSUBS 0.076208f
C1277 VP.n91 VSUBS 0.081059f
C1278 VP.n92 VSUBS 0.04089f
C1279 VP.n93 VSUBS 0.04089f
C1280 VP.n94 VSUBS 0.04089f
C1281 VP.n95 VSUBS 0.081469f
C1282 VP.n96 VSUBS 0.076208f
C1283 VP.n97 VSUBS 0.056643f
C1284 VP.n98 VSUBS 0.04089f
C1285 VP.n99 VSUBS 0.04089f
C1286 VP.n100 VSUBS 0.058148f
C1287 VP.n101 VSUBS 0.076208f
C1288 VP.n102 VSUBS 0.080598f
C1289 VP.n103 VSUBS 0.04089f
C1290 VP.n104 VSUBS 0.04089f
C1291 VP.n105 VSUBS 0.04089f
C1292 VP.n106 VSUBS 0.081825f
C1293 VP.n107 VSUBS 0.076208f
C1294 VP.n108 VSUBS 0.055891f
C1295 VP.n109 VSUBS 0.065995f
C1296 VP.n110 VSUBS 0.10158f
.ends

