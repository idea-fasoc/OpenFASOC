* NGSPICE file created from diff_pair_sample_0515.ext - technology: sky130A

.subckt diff_pair_sample_0515 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=0 ps=0 w=15.08 l=2.15
X1 VTAIL.t19 VP.t0 VDD1.t4 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X2 VDD2.t9 VN.t0 VTAIL.t8 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X3 VDD2.t8 VN.t1 VTAIL.t7 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=5.8812 ps=30.94 w=15.08 l=2.15
X4 VDD1.t3 VP.t1 VTAIL.t18 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X5 VDD1.t8 VP.t2 VTAIL.t17 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=5.8812 ps=30.94 w=15.08 l=2.15
X6 VTAIL.t1 VN.t2 VDD2.t7 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X7 VDD1.t0 VP.t3 VTAIL.t16 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=2.4882 ps=15.41 w=15.08 l=2.15
X8 B.t8 B.t6 B.t7 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=0 ps=0 w=15.08 l=2.15
X9 VDD2.t6 VN.t3 VTAIL.t6 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=5.8812 ps=30.94 w=15.08 l=2.15
X10 VTAIL.t5 VN.t4 VDD2.t5 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X11 VTAIL.t15 VP.t4 VDD1.t1 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X12 B.t5 B.t3 B.t4 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=0 ps=0 w=15.08 l=2.15
X13 VDD2.t4 VN.t5 VTAIL.t4 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=2.4882 ps=15.41 w=15.08 l=2.15
X14 VDD2.t3 VN.t6 VTAIL.t3 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X15 VTAIL.t14 VP.t5 VDD1.t5 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X16 VDD1.t2 VP.t6 VTAIL.t13 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=5.8812 ps=30.94 w=15.08 l=2.15
X17 B.t2 B.t0 B.t1 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=0 ps=0 w=15.08 l=2.15
X18 VTAIL.t9 VN.t7 VDD2.t2 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X19 VDD1.t6 VP.t7 VTAIL.t12 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=2.4882 ps=15.41 w=15.08 l=2.15
X20 VDD2.t1 VN.t8 VTAIL.t2 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=5.8812 pd=30.94 as=2.4882 ps=15.41 w=15.08 l=2.15
X21 VDD1.t9 VP.t8 VTAIL.t11 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X22 VTAIL.t0 VN.t9 VDD2.t0 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
X23 VTAIL.t10 VP.t9 VDD1.t7 w_n3946_n3984# sky130_fd_pr__pfet_01v8 ad=2.4882 pd=15.41 as=2.4882 ps=15.41 w=15.08 l=2.15
R0 B.n629 B.n628 585
R1 B.n630 B.n87 585
R2 B.n632 B.n631 585
R3 B.n633 B.n86 585
R4 B.n635 B.n634 585
R5 B.n636 B.n85 585
R6 B.n638 B.n637 585
R7 B.n639 B.n84 585
R8 B.n641 B.n640 585
R9 B.n642 B.n83 585
R10 B.n644 B.n643 585
R11 B.n645 B.n82 585
R12 B.n647 B.n646 585
R13 B.n648 B.n81 585
R14 B.n650 B.n649 585
R15 B.n651 B.n80 585
R16 B.n653 B.n652 585
R17 B.n654 B.n79 585
R18 B.n656 B.n655 585
R19 B.n657 B.n78 585
R20 B.n659 B.n658 585
R21 B.n660 B.n77 585
R22 B.n662 B.n661 585
R23 B.n663 B.n76 585
R24 B.n665 B.n664 585
R25 B.n666 B.n75 585
R26 B.n668 B.n667 585
R27 B.n669 B.n74 585
R28 B.n671 B.n670 585
R29 B.n672 B.n73 585
R30 B.n674 B.n673 585
R31 B.n675 B.n72 585
R32 B.n677 B.n676 585
R33 B.n678 B.n71 585
R34 B.n680 B.n679 585
R35 B.n681 B.n70 585
R36 B.n683 B.n682 585
R37 B.n684 B.n69 585
R38 B.n686 B.n685 585
R39 B.n687 B.n68 585
R40 B.n689 B.n688 585
R41 B.n690 B.n67 585
R42 B.n692 B.n691 585
R43 B.n693 B.n66 585
R44 B.n695 B.n694 585
R45 B.n696 B.n65 585
R46 B.n698 B.n697 585
R47 B.n699 B.n64 585
R48 B.n701 B.n700 585
R49 B.n702 B.n63 585
R50 B.n704 B.n703 585
R51 B.n706 B.n705 585
R52 B.n707 B.n59 585
R53 B.n709 B.n708 585
R54 B.n710 B.n58 585
R55 B.n712 B.n711 585
R56 B.n713 B.n57 585
R57 B.n715 B.n714 585
R58 B.n716 B.n56 585
R59 B.n718 B.n717 585
R60 B.n720 B.n53 585
R61 B.n722 B.n721 585
R62 B.n723 B.n52 585
R63 B.n725 B.n724 585
R64 B.n726 B.n51 585
R65 B.n728 B.n727 585
R66 B.n729 B.n50 585
R67 B.n731 B.n730 585
R68 B.n732 B.n49 585
R69 B.n734 B.n733 585
R70 B.n735 B.n48 585
R71 B.n737 B.n736 585
R72 B.n738 B.n47 585
R73 B.n740 B.n739 585
R74 B.n741 B.n46 585
R75 B.n743 B.n742 585
R76 B.n744 B.n45 585
R77 B.n746 B.n745 585
R78 B.n747 B.n44 585
R79 B.n749 B.n748 585
R80 B.n750 B.n43 585
R81 B.n752 B.n751 585
R82 B.n753 B.n42 585
R83 B.n755 B.n754 585
R84 B.n756 B.n41 585
R85 B.n758 B.n757 585
R86 B.n759 B.n40 585
R87 B.n761 B.n760 585
R88 B.n762 B.n39 585
R89 B.n764 B.n763 585
R90 B.n765 B.n38 585
R91 B.n767 B.n766 585
R92 B.n768 B.n37 585
R93 B.n770 B.n769 585
R94 B.n771 B.n36 585
R95 B.n773 B.n772 585
R96 B.n774 B.n35 585
R97 B.n776 B.n775 585
R98 B.n777 B.n34 585
R99 B.n779 B.n778 585
R100 B.n780 B.n33 585
R101 B.n782 B.n781 585
R102 B.n783 B.n32 585
R103 B.n785 B.n784 585
R104 B.n786 B.n31 585
R105 B.n788 B.n787 585
R106 B.n789 B.n30 585
R107 B.n791 B.n790 585
R108 B.n792 B.n29 585
R109 B.n794 B.n793 585
R110 B.n795 B.n28 585
R111 B.n627 B.n88 585
R112 B.n626 B.n625 585
R113 B.n624 B.n89 585
R114 B.n623 B.n622 585
R115 B.n621 B.n90 585
R116 B.n620 B.n619 585
R117 B.n618 B.n91 585
R118 B.n617 B.n616 585
R119 B.n615 B.n92 585
R120 B.n614 B.n613 585
R121 B.n612 B.n93 585
R122 B.n611 B.n610 585
R123 B.n609 B.n94 585
R124 B.n608 B.n607 585
R125 B.n606 B.n95 585
R126 B.n605 B.n604 585
R127 B.n603 B.n96 585
R128 B.n602 B.n601 585
R129 B.n600 B.n97 585
R130 B.n599 B.n598 585
R131 B.n597 B.n98 585
R132 B.n596 B.n595 585
R133 B.n594 B.n99 585
R134 B.n593 B.n592 585
R135 B.n591 B.n100 585
R136 B.n590 B.n589 585
R137 B.n588 B.n101 585
R138 B.n587 B.n586 585
R139 B.n585 B.n102 585
R140 B.n584 B.n583 585
R141 B.n582 B.n103 585
R142 B.n581 B.n580 585
R143 B.n579 B.n104 585
R144 B.n578 B.n577 585
R145 B.n576 B.n105 585
R146 B.n575 B.n574 585
R147 B.n573 B.n106 585
R148 B.n572 B.n571 585
R149 B.n570 B.n107 585
R150 B.n569 B.n568 585
R151 B.n567 B.n108 585
R152 B.n566 B.n565 585
R153 B.n564 B.n109 585
R154 B.n563 B.n562 585
R155 B.n561 B.n110 585
R156 B.n560 B.n559 585
R157 B.n558 B.n111 585
R158 B.n557 B.n556 585
R159 B.n555 B.n112 585
R160 B.n554 B.n553 585
R161 B.n552 B.n113 585
R162 B.n551 B.n550 585
R163 B.n549 B.n114 585
R164 B.n548 B.n547 585
R165 B.n546 B.n115 585
R166 B.n545 B.n544 585
R167 B.n543 B.n116 585
R168 B.n542 B.n541 585
R169 B.n540 B.n117 585
R170 B.n539 B.n538 585
R171 B.n537 B.n118 585
R172 B.n536 B.n535 585
R173 B.n534 B.n119 585
R174 B.n533 B.n532 585
R175 B.n531 B.n120 585
R176 B.n530 B.n529 585
R177 B.n528 B.n121 585
R178 B.n527 B.n526 585
R179 B.n525 B.n122 585
R180 B.n524 B.n523 585
R181 B.n522 B.n123 585
R182 B.n521 B.n520 585
R183 B.n519 B.n124 585
R184 B.n518 B.n517 585
R185 B.n516 B.n125 585
R186 B.n515 B.n514 585
R187 B.n513 B.n126 585
R188 B.n512 B.n511 585
R189 B.n510 B.n127 585
R190 B.n509 B.n508 585
R191 B.n507 B.n128 585
R192 B.n506 B.n505 585
R193 B.n504 B.n129 585
R194 B.n503 B.n502 585
R195 B.n501 B.n130 585
R196 B.n500 B.n499 585
R197 B.n498 B.n131 585
R198 B.n497 B.n496 585
R199 B.n495 B.n132 585
R200 B.n494 B.n493 585
R201 B.n492 B.n133 585
R202 B.n491 B.n490 585
R203 B.n489 B.n134 585
R204 B.n488 B.n487 585
R205 B.n486 B.n135 585
R206 B.n485 B.n484 585
R207 B.n483 B.n136 585
R208 B.n482 B.n481 585
R209 B.n480 B.n137 585
R210 B.n479 B.n478 585
R211 B.n477 B.n138 585
R212 B.n476 B.n475 585
R213 B.n474 B.n139 585
R214 B.n473 B.n472 585
R215 B.n471 B.n140 585
R216 B.n303 B.n200 585
R217 B.n305 B.n304 585
R218 B.n306 B.n199 585
R219 B.n308 B.n307 585
R220 B.n309 B.n198 585
R221 B.n311 B.n310 585
R222 B.n312 B.n197 585
R223 B.n314 B.n313 585
R224 B.n315 B.n196 585
R225 B.n317 B.n316 585
R226 B.n318 B.n195 585
R227 B.n320 B.n319 585
R228 B.n321 B.n194 585
R229 B.n323 B.n322 585
R230 B.n324 B.n193 585
R231 B.n326 B.n325 585
R232 B.n327 B.n192 585
R233 B.n329 B.n328 585
R234 B.n330 B.n191 585
R235 B.n332 B.n331 585
R236 B.n333 B.n190 585
R237 B.n335 B.n334 585
R238 B.n336 B.n189 585
R239 B.n338 B.n337 585
R240 B.n339 B.n188 585
R241 B.n341 B.n340 585
R242 B.n342 B.n187 585
R243 B.n344 B.n343 585
R244 B.n345 B.n186 585
R245 B.n347 B.n346 585
R246 B.n348 B.n185 585
R247 B.n350 B.n349 585
R248 B.n351 B.n184 585
R249 B.n353 B.n352 585
R250 B.n354 B.n183 585
R251 B.n356 B.n355 585
R252 B.n357 B.n182 585
R253 B.n359 B.n358 585
R254 B.n360 B.n181 585
R255 B.n362 B.n361 585
R256 B.n363 B.n180 585
R257 B.n365 B.n364 585
R258 B.n366 B.n179 585
R259 B.n368 B.n367 585
R260 B.n369 B.n178 585
R261 B.n371 B.n370 585
R262 B.n372 B.n177 585
R263 B.n374 B.n373 585
R264 B.n375 B.n176 585
R265 B.n377 B.n376 585
R266 B.n378 B.n173 585
R267 B.n381 B.n380 585
R268 B.n382 B.n172 585
R269 B.n384 B.n383 585
R270 B.n385 B.n171 585
R271 B.n387 B.n386 585
R272 B.n388 B.n170 585
R273 B.n390 B.n389 585
R274 B.n391 B.n169 585
R275 B.n393 B.n392 585
R276 B.n395 B.n394 585
R277 B.n396 B.n165 585
R278 B.n398 B.n397 585
R279 B.n399 B.n164 585
R280 B.n401 B.n400 585
R281 B.n402 B.n163 585
R282 B.n404 B.n403 585
R283 B.n405 B.n162 585
R284 B.n407 B.n406 585
R285 B.n408 B.n161 585
R286 B.n410 B.n409 585
R287 B.n411 B.n160 585
R288 B.n413 B.n412 585
R289 B.n414 B.n159 585
R290 B.n416 B.n415 585
R291 B.n417 B.n158 585
R292 B.n419 B.n418 585
R293 B.n420 B.n157 585
R294 B.n422 B.n421 585
R295 B.n423 B.n156 585
R296 B.n425 B.n424 585
R297 B.n426 B.n155 585
R298 B.n428 B.n427 585
R299 B.n429 B.n154 585
R300 B.n431 B.n430 585
R301 B.n432 B.n153 585
R302 B.n434 B.n433 585
R303 B.n435 B.n152 585
R304 B.n437 B.n436 585
R305 B.n438 B.n151 585
R306 B.n440 B.n439 585
R307 B.n441 B.n150 585
R308 B.n443 B.n442 585
R309 B.n444 B.n149 585
R310 B.n446 B.n445 585
R311 B.n447 B.n148 585
R312 B.n449 B.n448 585
R313 B.n450 B.n147 585
R314 B.n452 B.n451 585
R315 B.n453 B.n146 585
R316 B.n455 B.n454 585
R317 B.n456 B.n145 585
R318 B.n458 B.n457 585
R319 B.n459 B.n144 585
R320 B.n461 B.n460 585
R321 B.n462 B.n143 585
R322 B.n464 B.n463 585
R323 B.n465 B.n142 585
R324 B.n467 B.n466 585
R325 B.n468 B.n141 585
R326 B.n470 B.n469 585
R327 B.n302 B.n301 585
R328 B.n300 B.n201 585
R329 B.n299 B.n298 585
R330 B.n297 B.n202 585
R331 B.n296 B.n295 585
R332 B.n294 B.n203 585
R333 B.n293 B.n292 585
R334 B.n291 B.n204 585
R335 B.n290 B.n289 585
R336 B.n288 B.n205 585
R337 B.n287 B.n286 585
R338 B.n285 B.n206 585
R339 B.n284 B.n283 585
R340 B.n282 B.n207 585
R341 B.n281 B.n280 585
R342 B.n279 B.n208 585
R343 B.n278 B.n277 585
R344 B.n276 B.n209 585
R345 B.n275 B.n274 585
R346 B.n273 B.n210 585
R347 B.n272 B.n271 585
R348 B.n270 B.n211 585
R349 B.n269 B.n268 585
R350 B.n267 B.n212 585
R351 B.n266 B.n265 585
R352 B.n264 B.n213 585
R353 B.n263 B.n262 585
R354 B.n261 B.n214 585
R355 B.n260 B.n259 585
R356 B.n258 B.n215 585
R357 B.n257 B.n256 585
R358 B.n255 B.n216 585
R359 B.n254 B.n253 585
R360 B.n252 B.n217 585
R361 B.n251 B.n250 585
R362 B.n249 B.n218 585
R363 B.n248 B.n247 585
R364 B.n246 B.n219 585
R365 B.n245 B.n244 585
R366 B.n243 B.n220 585
R367 B.n242 B.n241 585
R368 B.n240 B.n221 585
R369 B.n239 B.n238 585
R370 B.n237 B.n222 585
R371 B.n236 B.n235 585
R372 B.n234 B.n223 585
R373 B.n233 B.n232 585
R374 B.n231 B.n224 585
R375 B.n230 B.n229 585
R376 B.n228 B.n225 585
R377 B.n227 B.n226 585
R378 B.n2 B.n0 585
R379 B.n873 B.n1 585
R380 B.n872 B.n871 585
R381 B.n870 B.n3 585
R382 B.n869 B.n868 585
R383 B.n867 B.n4 585
R384 B.n866 B.n865 585
R385 B.n864 B.n5 585
R386 B.n863 B.n862 585
R387 B.n861 B.n6 585
R388 B.n860 B.n859 585
R389 B.n858 B.n7 585
R390 B.n857 B.n856 585
R391 B.n855 B.n8 585
R392 B.n854 B.n853 585
R393 B.n852 B.n9 585
R394 B.n851 B.n850 585
R395 B.n849 B.n10 585
R396 B.n848 B.n847 585
R397 B.n846 B.n11 585
R398 B.n845 B.n844 585
R399 B.n843 B.n12 585
R400 B.n842 B.n841 585
R401 B.n840 B.n13 585
R402 B.n839 B.n838 585
R403 B.n837 B.n14 585
R404 B.n836 B.n835 585
R405 B.n834 B.n15 585
R406 B.n833 B.n832 585
R407 B.n831 B.n16 585
R408 B.n830 B.n829 585
R409 B.n828 B.n17 585
R410 B.n827 B.n826 585
R411 B.n825 B.n18 585
R412 B.n824 B.n823 585
R413 B.n822 B.n19 585
R414 B.n821 B.n820 585
R415 B.n819 B.n20 585
R416 B.n818 B.n817 585
R417 B.n816 B.n21 585
R418 B.n815 B.n814 585
R419 B.n813 B.n22 585
R420 B.n812 B.n811 585
R421 B.n810 B.n23 585
R422 B.n809 B.n808 585
R423 B.n807 B.n24 585
R424 B.n806 B.n805 585
R425 B.n804 B.n25 585
R426 B.n803 B.n802 585
R427 B.n801 B.n26 585
R428 B.n800 B.n799 585
R429 B.n798 B.n27 585
R430 B.n797 B.n796 585
R431 B.n875 B.n874 585
R432 B.n303 B.n302 473.281
R433 B.n796 B.n795 473.281
R434 B.n471 B.n470 473.281
R435 B.n628 B.n627 473.281
R436 B.n166 B.t3 376.286
R437 B.n174 B.t0 376.286
R438 B.n54 B.t6 376.286
R439 B.n60 B.t9 376.286
R440 B.n302 B.n201 163.367
R441 B.n298 B.n201 163.367
R442 B.n298 B.n297 163.367
R443 B.n297 B.n296 163.367
R444 B.n296 B.n203 163.367
R445 B.n292 B.n203 163.367
R446 B.n292 B.n291 163.367
R447 B.n291 B.n290 163.367
R448 B.n290 B.n205 163.367
R449 B.n286 B.n205 163.367
R450 B.n286 B.n285 163.367
R451 B.n285 B.n284 163.367
R452 B.n284 B.n207 163.367
R453 B.n280 B.n207 163.367
R454 B.n280 B.n279 163.367
R455 B.n279 B.n278 163.367
R456 B.n278 B.n209 163.367
R457 B.n274 B.n209 163.367
R458 B.n274 B.n273 163.367
R459 B.n273 B.n272 163.367
R460 B.n272 B.n211 163.367
R461 B.n268 B.n211 163.367
R462 B.n268 B.n267 163.367
R463 B.n267 B.n266 163.367
R464 B.n266 B.n213 163.367
R465 B.n262 B.n213 163.367
R466 B.n262 B.n261 163.367
R467 B.n261 B.n260 163.367
R468 B.n260 B.n215 163.367
R469 B.n256 B.n215 163.367
R470 B.n256 B.n255 163.367
R471 B.n255 B.n254 163.367
R472 B.n254 B.n217 163.367
R473 B.n250 B.n217 163.367
R474 B.n250 B.n249 163.367
R475 B.n249 B.n248 163.367
R476 B.n248 B.n219 163.367
R477 B.n244 B.n219 163.367
R478 B.n244 B.n243 163.367
R479 B.n243 B.n242 163.367
R480 B.n242 B.n221 163.367
R481 B.n238 B.n221 163.367
R482 B.n238 B.n237 163.367
R483 B.n237 B.n236 163.367
R484 B.n236 B.n223 163.367
R485 B.n232 B.n223 163.367
R486 B.n232 B.n231 163.367
R487 B.n231 B.n230 163.367
R488 B.n230 B.n225 163.367
R489 B.n226 B.n225 163.367
R490 B.n226 B.n2 163.367
R491 B.n874 B.n2 163.367
R492 B.n874 B.n873 163.367
R493 B.n873 B.n872 163.367
R494 B.n872 B.n3 163.367
R495 B.n868 B.n3 163.367
R496 B.n868 B.n867 163.367
R497 B.n867 B.n866 163.367
R498 B.n866 B.n5 163.367
R499 B.n862 B.n5 163.367
R500 B.n862 B.n861 163.367
R501 B.n861 B.n860 163.367
R502 B.n860 B.n7 163.367
R503 B.n856 B.n7 163.367
R504 B.n856 B.n855 163.367
R505 B.n855 B.n854 163.367
R506 B.n854 B.n9 163.367
R507 B.n850 B.n9 163.367
R508 B.n850 B.n849 163.367
R509 B.n849 B.n848 163.367
R510 B.n848 B.n11 163.367
R511 B.n844 B.n11 163.367
R512 B.n844 B.n843 163.367
R513 B.n843 B.n842 163.367
R514 B.n842 B.n13 163.367
R515 B.n838 B.n13 163.367
R516 B.n838 B.n837 163.367
R517 B.n837 B.n836 163.367
R518 B.n836 B.n15 163.367
R519 B.n832 B.n15 163.367
R520 B.n832 B.n831 163.367
R521 B.n831 B.n830 163.367
R522 B.n830 B.n17 163.367
R523 B.n826 B.n17 163.367
R524 B.n826 B.n825 163.367
R525 B.n825 B.n824 163.367
R526 B.n824 B.n19 163.367
R527 B.n820 B.n19 163.367
R528 B.n820 B.n819 163.367
R529 B.n819 B.n818 163.367
R530 B.n818 B.n21 163.367
R531 B.n814 B.n21 163.367
R532 B.n814 B.n813 163.367
R533 B.n813 B.n812 163.367
R534 B.n812 B.n23 163.367
R535 B.n808 B.n23 163.367
R536 B.n808 B.n807 163.367
R537 B.n807 B.n806 163.367
R538 B.n806 B.n25 163.367
R539 B.n802 B.n25 163.367
R540 B.n802 B.n801 163.367
R541 B.n801 B.n800 163.367
R542 B.n800 B.n27 163.367
R543 B.n796 B.n27 163.367
R544 B.n304 B.n303 163.367
R545 B.n304 B.n199 163.367
R546 B.n308 B.n199 163.367
R547 B.n309 B.n308 163.367
R548 B.n310 B.n309 163.367
R549 B.n310 B.n197 163.367
R550 B.n314 B.n197 163.367
R551 B.n315 B.n314 163.367
R552 B.n316 B.n315 163.367
R553 B.n316 B.n195 163.367
R554 B.n320 B.n195 163.367
R555 B.n321 B.n320 163.367
R556 B.n322 B.n321 163.367
R557 B.n322 B.n193 163.367
R558 B.n326 B.n193 163.367
R559 B.n327 B.n326 163.367
R560 B.n328 B.n327 163.367
R561 B.n328 B.n191 163.367
R562 B.n332 B.n191 163.367
R563 B.n333 B.n332 163.367
R564 B.n334 B.n333 163.367
R565 B.n334 B.n189 163.367
R566 B.n338 B.n189 163.367
R567 B.n339 B.n338 163.367
R568 B.n340 B.n339 163.367
R569 B.n340 B.n187 163.367
R570 B.n344 B.n187 163.367
R571 B.n345 B.n344 163.367
R572 B.n346 B.n345 163.367
R573 B.n346 B.n185 163.367
R574 B.n350 B.n185 163.367
R575 B.n351 B.n350 163.367
R576 B.n352 B.n351 163.367
R577 B.n352 B.n183 163.367
R578 B.n356 B.n183 163.367
R579 B.n357 B.n356 163.367
R580 B.n358 B.n357 163.367
R581 B.n358 B.n181 163.367
R582 B.n362 B.n181 163.367
R583 B.n363 B.n362 163.367
R584 B.n364 B.n363 163.367
R585 B.n364 B.n179 163.367
R586 B.n368 B.n179 163.367
R587 B.n369 B.n368 163.367
R588 B.n370 B.n369 163.367
R589 B.n370 B.n177 163.367
R590 B.n374 B.n177 163.367
R591 B.n375 B.n374 163.367
R592 B.n376 B.n375 163.367
R593 B.n376 B.n173 163.367
R594 B.n381 B.n173 163.367
R595 B.n382 B.n381 163.367
R596 B.n383 B.n382 163.367
R597 B.n383 B.n171 163.367
R598 B.n387 B.n171 163.367
R599 B.n388 B.n387 163.367
R600 B.n389 B.n388 163.367
R601 B.n389 B.n169 163.367
R602 B.n393 B.n169 163.367
R603 B.n394 B.n393 163.367
R604 B.n394 B.n165 163.367
R605 B.n398 B.n165 163.367
R606 B.n399 B.n398 163.367
R607 B.n400 B.n399 163.367
R608 B.n400 B.n163 163.367
R609 B.n404 B.n163 163.367
R610 B.n405 B.n404 163.367
R611 B.n406 B.n405 163.367
R612 B.n406 B.n161 163.367
R613 B.n410 B.n161 163.367
R614 B.n411 B.n410 163.367
R615 B.n412 B.n411 163.367
R616 B.n412 B.n159 163.367
R617 B.n416 B.n159 163.367
R618 B.n417 B.n416 163.367
R619 B.n418 B.n417 163.367
R620 B.n418 B.n157 163.367
R621 B.n422 B.n157 163.367
R622 B.n423 B.n422 163.367
R623 B.n424 B.n423 163.367
R624 B.n424 B.n155 163.367
R625 B.n428 B.n155 163.367
R626 B.n429 B.n428 163.367
R627 B.n430 B.n429 163.367
R628 B.n430 B.n153 163.367
R629 B.n434 B.n153 163.367
R630 B.n435 B.n434 163.367
R631 B.n436 B.n435 163.367
R632 B.n436 B.n151 163.367
R633 B.n440 B.n151 163.367
R634 B.n441 B.n440 163.367
R635 B.n442 B.n441 163.367
R636 B.n442 B.n149 163.367
R637 B.n446 B.n149 163.367
R638 B.n447 B.n446 163.367
R639 B.n448 B.n447 163.367
R640 B.n448 B.n147 163.367
R641 B.n452 B.n147 163.367
R642 B.n453 B.n452 163.367
R643 B.n454 B.n453 163.367
R644 B.n454 B.n145 163.367
R645 B.n458 B.n145 163.367
R646 B.n459 B.n458 163.367
R647 B.n460 B.n459 163.367
R648 B.n460 B.n143 163.367
R649 B.n464 B.n143 163.367
R650 B.n465 B.n464 163.367
R651 B.n466 B.n465 163.367
R652 B.n466 B.n141 163.367
R653 B.n470 B.n141 163.367
R654 B.n472 B.n471 163.367
R655 B.n472 B.n139 163.367
R656 B.n476 B.n139 163.367
R657 B.n477 B.n476 163.367
R658 B.n478 B.n477 163.367
R659 B.n478 B.n137 163.367
R660 B.n482 B.n137 163.367
R661 B.n483 B.n482 163.367
R662 B.n484 B.n483 163.367
R663 B.n484 B.n135 163.367
R664 B.n488 B.n135 163.367
R665 B.n489 B.n488 163.367
R666 B.n490 B.n489 163.367
R667 B.n490 B.n133 163.367
R668 B.n494 B.n133 163.367
R669 B.n495 B.n494 163.367
R670 B.n496 B.n495 163.367
R671 B.n496 B.n131 163.367
R672 B.n500 B.n131 163.367
R673 B.n501 B.n500 163.367
R674 B.n502 B.n501 163.367
R675 B.n502 B.n129 163.367
R676 B.n506 B.n129 163.367
R677 B.n507 B.n506 163.367
R678 B.n508 B.n507 163.367
R679 B.n508 B.n127 163.367
R680 B.n512 B.n127 163.367
R681 B.n513 B.n512 163.367
R682 B.n514 B.n513 163.367
R683 B.n514 B.n125 163.367
R684 B.n518 B.n125 163.367
R685 B.n519 B.n518 163.367
R686 B.n520 B.n519 163.367
R687 B.n520 B.n123 163.367
R688 B.n524 B.n123 163.367
R689 B.n525 B.n524 163.367
R690 B.n526 B.n525 163.367
R691 B.n526 B.n121 163.367
R692 B.n530 B.n121 163.367
R693 B.n531 B.n530 163.367
R694 B.n532 B.n531 163.367
R695 B.n532 B.n119 163.367
R696 B.n536 B.n119 163.367
R697 B.n537 B.n536 163.367
R698 B.n538 B.n537 163.367
R699 B.n538 B.n117 163.367
R700 B.n542 B.n117 163.367
R701 B.n543 B.n542 163.367
R702 B.n544 B.n543 163.367
R703 B.n544 B.n115 163.367
R704 B.n548 B.n115 163.367
R705 B.n549 B.n548 163.367
R706 B.n550 B.n549 163.367
R707 B.n550 B.n113 163.367
R708 B.n554 B.n113 163.367
R709 B.n555 B.n554 163.367
R710 B.n556 B.n555 163.367
R711 B.n556 B.n111 163.367
R712 B.n560 B.n111 163.367
R713 B.n561 B.n560 163.367
R714 B.n562 B.n561 163.367
R715 B.n562 B.n109 163.367
R716 B.n566 B.n109 163.367
R717 B.n567 B.n566 163.367
R718 B.n568 B.n567 163.367
R719 B.n568 B.n107 163.367
R720 B.n572 B.n107 163.367
R721 B.n573 B.n572 163.367
R722 B.n574 B.n573 163.367
R723 B.n574 B.n105 163.367
R724 B.n578 B.n105 163.367
R725 B.n579 B.n578 163.367
R726 B.n580 B.n579 163.367
R727 B.n580 B.n103 163.367
R728 B.n584 B.n103 163.367
R729 B.n585 B.n584 163.367
R730 B.n586 B.n585 163.367
R731 B.n586 B.n101 163.367
R732 B.n590 B.n101 163.367
R733 B.n591 B.n590 163.367
R734 B.n592 B.n591 163.367
R735 B.n592 B.n99 163.367
R736 B.n596 B.n99 163.367
R737 B.n597 B.n596 163.367
R738 B.n598 B.n597 163.367
R739 B.n598 B.n97 163.367
R740 B.n602 B.n97 163.367
R741 B.n603 B.n602 163.367
R742 B.n604 B.n603 163.367
R743 B.n604 B.n95 163.367
R744 B.n608 B.n95 163.367
R745 B.n609 B.n608 163.367
R746 B.n610 B.n609 163.367
R747 B.n610 B.n93 163.367
R748 B.n614 B.n93 163.367
R749 B.n615 B.n614 163.367
R750 B.n616 B.n615 163.367
R751 B.n616 B.n91 163.367
R752 B.n620 B.n91 163.367
R753 B.n621 B.n620 163.367
R754 B.n622 B.n621 163.367
R755 B.n622 B.n89 163.367
R756 B.n626 B.n89 163.367
R757 B.n627 B.n626 163.367
R758 B.n795 B.n794 163.367
R759 B.n794 B.n29 163.367
R760 B.n790 B.n29 163.367
R761 B.n790 B.n789 163.367
R762 B.n789 B.n788 163.367
R763 B.n788 B.n31 163.367
R764 B.n784 B.n31 163.367
R765 B.n784 B.n783 163.367
R766 B.n783 B.n782 163.367
R767 B.n782 B.n33 163.367
R768 B.n778 B.n33 163.367
R769 B.n778 B.n777 163.367
R770 B.n777 B.n776 163.367
R771 B.n776 B.n35 163.367
R772 B.n772 B.n35 163.367
R773 B.n772 B.n771 163.367
R774 B.n771 B.n770 163.367
R775 B.n770 B.n37 163.367
R776 B.n766 B.n37 163.367
R777 B.n766 B.n765 163.367
R778 B.n765 B.n764 163.367
R779 B.n764 B.n39 163.367
R780 B.n760 B.n39 163.367
R781 B.n760 B.n759 163.367
R782 B.n759 B.n758 163.367
R783 B.n758 B.n41 163.367
R784 B.n754 B.n41 163.367
R785 B.n754 B.n753 163.367
R786 B.n753 B.n752 163.367
R787 B.n752 B.n43 163.367
R788 B.n748 B.n43 163.367
R789 B.n748 B.n747 163.367
R790 B.n747 B.n746 163.367
R791 B.n746 B.n45 163.367
R792 B.n742 B.n45 163.367
R793 B.n742 B.n741 163.367
R794 B.n741 B.n740 163.367
R795 B.n740 B.n47 163.367
R796 B.n736 B.n47 163.367
R797 B.n736 B.n735 163.367
R798 B.n735 B.n734 163.367
R799 B.n734 B.n49 163.367
R800 B.n730 B.n49 163.367
R801 B.n730 B.n729 163.367
R802 B.n729 B.n728 163.367
R803 B.n728 B.n51 163.367
R804 B.n724 B.n51 163.367
R805 B.n724 B.n723 163.367
R806 B.n723 B.n722 163.367
R807 B.n722 B.n53 163.367
R808 B.n717 B.n53 163.367
R809 B.n717 B.n716 163.367
R810 B.n716 B.n715 163.367
R811 B.n715 B.n57 163.367
R812 B.n711 B.n57 163.367
R813 B.n711 B.n710 163.367
R814 B.n710 B.n709 163.367
R815 B.n709 B.n59 163.367
R816 B.n705 B.n59 163.367
R817 B.n705 B.n704 163.367
R818 B.n704 B.n63 163.367
R819 B.n700 B.n63 163.367
R820 B.n700 B.n699 163.367
R821 B.n699 B.n698 163.367
R822 B.n698 B.n65 163.367
R823 B.n694 B.n65 163.367
R824 B.n694 B.n693 163.367
R825 B.n693 B.n692 163.367
R826 B.n692 B.n67 163.367
R827 B.n688 B.n67 163.367
R828 B.n688 B.n687 163.367
R829 B.n687 B.n686 163.367
R830 B.n686 B.n69 163.367
R831 B.n682 B.n69 163.367
R832 B.n682 B.n681 163.367
R833 B.n681 B.n680 163.367
R834 B.n680 B.n71 163.367
R835 B.n676 B.n71 163.367
R836 B.n676 B.n675 163.367
R837 B.n675 B.n674 163.367
R838 B.n674 B.n73 163.367
R839 B.n670 B.n73 163.367
R840 B.n670 B.n669 163.367
R841 B.n669 B.n668 163.367
R842 B.n668 B.n75 163.367
R843 B.n664 B.n75 163.367
R844 B.n664 B.n663 163.367
R845 B.n663 B.n662 163.367
R846 B.n662 B.n77 163.367
R847 B.n658 B.n77 163.367
R848 B.n658 B.n657 163.367
R849 B.n657 B.n656 163.367
R850 B.n656 B.n79 163.367
R851 B.n652 B.n79 163.367
R852 B.n652 B.n651 163.367
R853 B.n651 B.n650 163.367
R854 B.n650 B.n81 163.367
R855 B.n646 B.n81 163.367
R856 B.n646 B.n645 163.367
R857 B.n645 B.n644 163.367
R858 B.n644 B.n83 163.367
R859 B.n640 B.n83 163.367
R860 B.n640 B.n639 163.367
R861 B.n639 B.n638 163.367
R862 B.n638 B.n85 163.367
R863 B.n634 B.n85 163.367
R864 B.n634 B.n633 163.367
R865 B.n633 B.n632 163.367
R866 B.n632 B.n87 163.367
R867 B.n628 B.n87 163.367
R868 B.n166 B.t5 156.975
R869 B.n60 B.t10 156.975
R870 B.n174 B.t2 156.956
R871 B.n54 B.t7 156.956
R872 B.n167 B.t4 108.877
R873 B.n61 B.t11 108.877
R874 B.n175 B.t1 108.859
R875 B.n55 B.t8 108.859
R876 B.n168 B.n167 59.5399
R877 B.n379 B.n175 59.5399
R878 B.n719 B.n55 59.5399
R879 B.n62 B.n61 59.5399
R880 B.n167 B.n166 48.0975
R881 B.n175 B.n174 48.0975
R882 B.n55 B.n54 48.0975
R883 B.n61 B.n60 48.0975
R884 B.n797 B.n28 30.7517
R885 B.n629 B.n88 30.7517
R886 B.n469 B.n140 30.7517
R887 B.n301 B.n200 30.7517
R888 B B.n875 18.0485
R889 B.n793 B.n28 10.6151
R890 B.n793 B.n792 10.6151
R891 B.n792 B.n791 10.6151
R892 B.n791 B.n30 10.6151
R893 B.n787 B.n30 10.6151
R894 B.n787 B.n786 10.6151
R895 B.n786 B.n785 10.6151
R896 B.n785 B.n32 10.6151
R897 B.n781 B.n32 10.6151
R898 B.n781 B.n780 10.6151
R899 B.n780 B.n779 10.6151
R900 B.n779 B.n34 10.6151
R901 B.n775 B.n34 10.6151
R902 B.n775 B.n774 10.6151
R903 B.n774 B.n773 10.6151
R904 B.n773 B.n36 10.6151
R905 B.n769 B.n36 10.6151
R906 B.n769 B.n768 10.6151
R907 B.n768 B.n767 10.6151
R908 B.n767 B.n38 10.6151
R909 B.n763 B.n38 10.6151
R910 B.n763 B.n762 10.6151
R911 B.n762 B.n761 10.6151
R912 B.n761 B.n40 10.6151
R913 B.n757 B.n40 10.6151
R914 B.n757 B.n756 10.6151
R915 B.n756 B.n755 10.6151
R916 B.n755 B.n42 10.6151
R917 B.n751 B.n42 10.6151
R918 B.n751 B.n750 10.6151
R919 B.n750 B.n749 10.6151
R920 B.n749 B.n44 10.6151
R921 B.n745 B.n44 10.6151
R922 B.n745 B.n744 10.6151
R923 B.n744 B.n743 10.6151
R924 B.n743 B.n46 10.6151
R925 B.n739 B.n46 10.6151
R926 B.n739 B.n738 10.6151
R927 B.n738 B.n737 10.6151
R928 B.n737 B.n48 10.6151
R929 B.n733 B.n48 10.6151
R930 B.n733 B.n732 10.6151
R931 B.n732 B.n731 10.6151
R932 B.n731 B.n50 10.6151
R933 B.n727 B.n50 10.6151
R934 B.n727 B.n726 10.6151
R935 B.n726 B.n725 10.6151
R936 B.n725 B.n52 10.6151
R937 B.n721 B.n52 10.6151
R938 B.n721 B.n720 10.6151
R939 B.n718 B.n56 10.6151
R940 B.n714 B.n56 10.6151
R941 B.n714 B.n713 10.6151
R942 B.n713 B.n712 10.6151
R943 B.n712 B.n58 10.6151
R944 B.n708 B.n58 10.6151
R945 B.n708 B.n707 10.6151
R946 B.n707 B.n706 10.6151
R947 B.n703 B.n702 10.6151
R948 B.n702 B.n701 10.6151
R949 B.n701 B.n64 10.6151
R950 B.n697 B.n64 10.6151
R951 B.n697 B.n696 10.6151
R952 B.n696 B.n695 10.6151
R953 B.n695 B.n66 10.6151
R954 B.n691 B.n66 10.6151
R955 B.n691 B.n690 10.6151
R956 B.n690 B.n689 10.6151
R957 B.n689 B.n68 10.6151
R958 B.n685 B.n68 10.6151
R959 B.n685 B.n684 10.6151
R960 B.n684 B.n683 10.6151
R961 B.n683 B.n70 10.6151
R962 B.n679 B.n70 10.6151
R963 B.n679 B.n678 10.6151
R964 B.n678 B.n677 10.6151
R965 B.n677 B.n72 10.6151
R966 B.n673 B.n72 10.6151
R967 B.n673 B.n672 10.6151
R968 B.n672 B.n671 10.6151
R969 B.n671 B.n74 10.6151
R970 B.n667 B.n74 10.6151
R971 B.n667 B.n666 10.6151
R972 B.n666 B.n665 10.6151
R973 B.n665 B.n76 10.6151
R974 B.n661 B.n76 10.6151
R975 B.n661 B.n660 10.6151
R976 B.n660 B.n659 10.6151
R977 B.n659 B.n78 10.6151
R978 B.n655 B.n78 10.6151
R979 B.n655 B.n654 10.6151
R980 B.n654 B.n653 10.6151
R981 B.n653 B.n80 10.6151
R982 B.n649 B.n80 10.6151
R983 B.n649 B.n648 10.6151
R984 B.n648 B.n647 10.6151
R985 B.n647 B.n82 10.6151
R986 B.n643 B.n82 10.6151
R987 B.n643 B.n642 10.6151
R988 B.n642 B.n641 10.6151
R989 B.n641 B.n84 10.6151
R990 B.n637 B.n84 10.6151
R991 B.n637 B.n636 10.6151
R992 B.n636 B.n635 10.6151
R993 B.n635 B.n86 10.6151
R994 B.n631 B.n86 10.6151
R995 B.n631 B.n630 10.6151
R996 B.n630 B.n629 10.6151
R997 B.n473 B.n140 10.6151
R998 B.n474 B.n473 10.6151
R999 B.n475 B.n474 10.6151
R1000 B.n475 B.n138 10.6151
R1001 B.n479 B.n138 10.6151
R1002 B.n480 B.n479 10.6151
R1003 B.n481 B.n480 10.6151
R1004 B.n481 B.n136 10.6151
R1005 B.n485 B.n136 10.6151
R1006 B.n486 B.n485 10.6151
R1007 B.n487 B.n486 10.6151
R1008 B.n487 B.n134 10.6151
R1009 B.n491 B.n134 10.6151
R1010 B.n492 B.n491 10.6151
R1011 B.n493 B.n492 10.6151
R1012 B.n493 B.n132 10.6151
R1013 B.n497 B.n132 10.6151
R1014 B.n498 B.n497 10.6151
R1015 B.n499 B.n498 10.6151
R1016 B.n499 B.n130 10.6151
R1017 B.n503 B.n130 10.6151
R1018 B.n504 B.n503 10.6151
R1019 B.n505 B.n504 10.6151
R1020 B.n505 B.n128 10.6151
R1021 B.n509 B.n128 10.6151
R1022 B.n510 B.n509 10.6151
R1023 B.n511 B.n510 10.6151
R1024 B.n511 B.n126 10.6151
R1025 B.n515 B.n126 10.6151
R1026 B.n516 B.n515 10.6151
R1027 B.n517 B.n516 10.6151
R1028 B.n517 B.n124 10.6151
R1029 B.n521 B.n124 10.6151
R1030 B.n522 B.n521 10.6151
R1031 B.n523 B.n522 10.6151
R1032 B.n523 B.n122 10.6151
R1033 B.n527 B.n122 10.6151
R1034 B.n528 B.n527 10.6151
R1035 B.n529 B.n528 10.6151
R1036 B.n529 B.n120 10.6151
R1037 B.n533 B.n120 10.6151
R1038 B.n534 B.n533 10.6151
R1039 B.n535 B.n534 10.6151
R1040 B.n535 B.n118 10.6151
R1041 B.n539 B.n118 10.6151
R1042 B.n540 B.n539 10.6151
R1043 B.n541 B.n540 10.6151
R1044 B.n541 B.n116 10.6151
R1045 B.n545 B.n116 10.6151
R1046 B.n546 B.n545 10.6151
R1047 B.n547 B.n546 10.6151
R1048 B.n547 B.n114 10.6151
R1049 B.n551 B.n114 10.6151
R1050 B.n552 B.n551 10.6151
R1051 B.n553 B.n552 10.6151
R1052 B.n553 B.n112 10.6151
R1053 B.n557 B.n112 10.6151
R1054 B.n558 B.n557 10.6151
R1055 B.n559 B.n558 10.6151
R1056 B.n559 B.n110 10.6151
R1057 B.n563 B.n110 10.6151
R1058 B.n564 B.n563 10.6151
R1059 B.n565 B.n564 10.6151
R1060 B.n565 B.n108 10.6151
R1061 B.n569 B.n108 10.6151
R1062 B.n570 B.n569 10.6151
R1063 B.n571 B.n570 10.6151
R1064 B.n571 B.n106 10.6151
R1065 B.n575 B.n106 10.6151
R1066 B.n576 B.n575 10.6151
R1067 B.n577 B.n576 10.6151
R1068 B.n577 B.n104 10.6151
R1069 B.n581 B.n104 10.6151
R1070 B.n582 B.n581 10.6151
R1071 B.n583 B.n582 10.6151
R1072 B.n583 B.n102 10.6151
R1073 B.n587 B.n102 10.6151
R1074 B.n588 B.n587 10.6151
R1075 B.n589 B.n588 10.6151
R1076 B.n589 B.n100 10.6151
R1077 B.n593 B.n100 10.6151
R1078 B.n594 B.n593 10.6151
R1079 B.n595 B.n594 10.6151
R1080 B.n595 B.n98 10.6151
R1081 B.n599 B.n98 10.6151
R1082 B.n600 B.n599 10.6151
R1083 B.n601 B.n600 10.6151
R1084 B.n601 B.n96 10.6151
R1085 B.n605 B.n96 10.6151
R1086 B.n606 B.n605 10.6151
R1087 B.n607 B.n606 10.6151
R1088 B.n607 B.n94 10.6151
R1089 B.n611 B.n94 10.6151
R1090 B.n612 B.n611 10.6151
R1091 B.n613 B.n612 10.6151
R1092 B.n613 B.n92 10.6151
R1093 B.n617 B.n92 10.6151
R1094 B.n618 B.n617 10.6151
R1095 B.n619 B.n618 10.6151
R1096 B.n619 B.n90 10.6151
R1097 B.n623 B.n90 10.6151
R1098 B.n624 B.n623 10.6151
R1099 B.n625 B.n624 10.6151
R1100 B.n625 B.n88 10.6151
R1101 B.n305 B.n200 10.6151
R1102 B.n306 B.n305 10.6151
R1103 B.n307 B.n306 10.6151
R1104 B.n307 B.n198 10.6151
R1105 B.n311 B.n198 10.6151
R1106 B.n312 B.n311 10.6151
R1107 B.n313 B.n312 10.6151
R1108 B.n313 B.n196 10.6151
R1109 B.n317 B.n196 10.6151
R1110 B.n318 B.n317 10.6151
R1111 B.n319 B.n318 10.6151
R1112 B.n319 B.n194 10.6151
R1113 B.n323 B.n194 10.6151
R1114 B.n324 B.n323 10.6151
R1115 B.n325 B.n324 10.6151
R1116 B.n325 B.n192 10.6151
R1117 B.n329 B.n192 10.6151
R1118 B.n330 B.n329 10.6151
R1119 B.n331 B.n330 10.6151
R1120 B.n331 B.n190 10.6151
R1121 B.n335 B.n190 10.6151
R1122 B.n336 B.n335 10.6151
R1123 B.n337 B.n336 10.6151
R1124 B.n337 B.n188 10.6151
R1125 B.n341 B.n188 10.6151
R1126 B.n342 B.n341 10.6151
R1127 B.n343 B.n342 10.6151
R1128 B.n343 B.n186 10.6151
R1129 B.n347 B.n186 10.6151
R1130 B.n348 B.n347 10.6151
R1131 B.n349 B.n348 10.6151
R1132 B.n349 B.n184 10.6151
R1133 B.n353 B.n184 10.6151
R1134 B.n354 B.n353 10.6151
R1135 B.n355 B.n354 10.6151
R1136 B.n355 B.n182 10.6151
R1137 B.n359 B.n182 10.6151
R1138 B.n360 B.n359 10.6151
R1139 B.n361 B.n360 10.6151
R1140 B.n361 B.n180 10.6151
R1141 B.n365 B.n180 10.6151
R1142 B.n366 B.n365 10.6151
R1143 B.n367 B.n366 10.6151
R1144 B.n367 B.n178 10.6151
R1145 B.n371 B.n178 10.6151
R1146 B.n372 B.n371 10.6151
R1147 B.n373 B.n372 10.6151
R1148 B.n373 B.n176 10.6151
R1149 B.n377 B.n176 10.6151
R1150 B.n378 B.n377 10.6151
R1151 B.n380 B.n172 10.6151
R1152 B.n384 B.n172 10.6151
R1153 B.n385 B.n384 10.6151
R1154 B.n386 B.n385 10.6151
R1155 B.n386 B.n170 10.6151
R1156 B.n390 B.n170 10.6151
R1157 B.n391 B.n390 10.6151
R1158 B.n392 B.n391 10.6151
R1159 B.n396 B.n395 10.6151
R1160 B.n397 B.n396 10.6151
R1161 B.n397 B.n164 10.6151
R1162 B.n401 B.n164 10.6151
R1163 B.n402 B.n401 10.6151
R1164 B.n403 B.n402 10.6151
R1165 B.n403 B.n162 10.6151
R1166 B.n407 B.n162 10.6151
R1167 B.n408 B.n407 10.6151
R1168 B.n409 B.n408 10.6151
R1169 B.n409 B.n160 10.6151
R1170 B.n413 B.n160 10.6151
R1171 B.n414 B.n413 10.6151
R1172 B.n415 B.n414 10.6151
R1173 B.n415 B.n158 10.6151
R1174 B.n419 B.n158 10.6151
R1175 B.n420 B.n419 10.6151
R1176 B.n421 B.n420 10.6151
R1177 B.n421 B.n156 10.6151
R1178 B.n425 B.n156 10.6151
R1179 B.n426 B.n425 10.6151
R1180 B.n427 B.n426 10.6151
R1181 B.n427 B.n154 10.6151
R1182 B.n431 B.n154 10.6151
R1183 B.n432 B.n431 10.6151
R1184 B.n433 B.n432 10.6151
R1185 B.n433 B.n152 10.6151
R1186 B.n437 B.n152 10.6151
R1187 B.n438 B.n437 10.6151
R1188 B.n439 B.n438 10.6151
R1189 B.n439 B.n150 10.6151
R1190 B.n443 B.n150 10.6151
R1191 B.n444 B.n443 10.6151
R1192 B.n445 B.n444 10.6151
R1193 B.n445 B.n148 10.6151
R1194 B.n449 B.n148 10.6151
R1195 B.n450 B.n449 10.6151
R1196 B.n451 B.n450 10.6151
R1197 B.n451 B.n146 10.6151
R1198 B.n455 B.n146 10.6151
R1199 B.n456 B.n455 10.6151
R1200 B.n457 B.n456 10.6151
R1201 B.n457 B.n144 10.6151
R1202 B.n461 B.n144 10.6151
R1203 B.n462 B.n461 10.6151
R1204 B.n463 B.n462 10.6151
R1205 B.n463 B.n142 10.6151
R1206 B.n467 B.n142 10.6151
R1207 B.n468 B.n467 10.6151
R1208 B.n469 B.n468 10.6151
R1209 B.n301 B.n300 10.6151
R1210 B.n300 B.n299 10.6151
R1211 B.n299 B.n202 10.6151
R1212 B.n295 B.n202 10.6151
R1213 B.n295 B.n294 10.6151
R1214 B.n294 B.n293 10.6151
R1215 B.n293 B.n204 10.6151
R1216 B.n289 B.n204 10.6151
R1217 B.n289 B.n288 10.6151
R1218 B.n288 B.n287 10.6151
R1219 B.n287 B.n206 10.6151
R1220 B.n283 B.n206 10.6151
R1221 B.n283 B.n282 10.6151
R1222 B.n282 B.n281 10.6151
R1223 B.n281 B.n208 10.6151
R1224 B.n277 B.n208 10.6151
R1225 B.n277 B.n276 10.6151
R1226 B.n276 B.n275 10.6151
R1227 B.n275 B.n210 10.6151
R1228 B.n271 B.n210 10.6151
R1229 B.n271 B.n270 10.6151
R1230 B.n270 B.n269 10.6151
R1231 B.n269 B.n212 10.6151
R1232 B.n265 B.n212 10.6151
R1233 B.n265 B.n264 10.6151
R1234 B.n264 B.n263 10.6151
R1235 B.n263 B.n214 10.6151
R1236 B.n259 B.n214 10.6151
R1237 B.n259 B.n258 10.6151
R1238 B.n258 B.n257 10.6151
R1239 B.n257 B.n216 10.6151
R1240 B.n253 B.n216 10.6151
R1241 B.n253 B.n252 10.6151
R1242 B.n252 B.n251 10.6151
R1243 B.n251 B.n218 10.6151
R1244 B.n247 B.n218 10.6151
R1245 B.n247 B.n246 10.6151
R1246 B.n246 B.n245 10.6151
R1247 B.n245 B.n220 10.6151
R1248 B.n241 B.n220 10.6151
R1249 B.n241 B.n240 10.6151
R1250 B.n240 B.n239 10.6151
R1251 B.n239 B.n222 10.6151
R1252 B.n235 B.n222 10.6151
R1253 B.n235 B.n234 10.6151
R1254 B.n234 B.n233 10.6151
R1255 B.n233 B.n224 10.6151
R1256 B.n229 B.n224 10.6151
R1257 B.n229 B.n228 10.6151
R1258 B.n228 B.n227 10.6151
R1259 B.n227 B.n0 10.6151
R1260 B.n871 B.n1 10.6151
R1261 B.n871 B.n870 10.6151
R1262 B.n870 B.n869 10.6151
R1263 B.n869 B.n4 10.6151
R1264 B.n865 B.n4 10.6151
R1265 B.n865 B.n864 10.6151
R1266 B.n864 B.n863 10.6151
R1267 B.n863 B.n6 10.6151
R1268 B.n859 B.n6 10.6151
R1269 B.n859 B.n858 10.6151
R1270 B.n858 B.n857 10.6151
R1271 B.n857 B.n8 10.6151
R1272 B.n853 B.n8 10.6151
R1273 B.n853 B.n852 10.6151
R1274 B.n852 B.n851 10.6151
R1275 B.n851 B.n10 10.6151
R1276 B.n847 B.n10 10.6151
R1277 B.n847 B.n846 10.6151
R1278 B.n846 B.n845 10.6151
R1279 B.n845 B.n12 10.6151
R1280 B.n841 B.n12 10.6151
R1281 B.n841 B.n840 10.6151
R1282 B.n840 B.n839 10.6151
R1283 B.n839 B.n14 10.6151
R1284 B.n835 B.n14 10.6151
R1285 B.n835 B.n834 10.6151
R1286 B.n834 B.n833 10.6151
R1287 B.n833 B.n16 10.6151
R1288 B.n829 B.n16 10.6151
R1289 B.n829 B.n828 10.6151
R1290 B.n828 B.n827 10.6151
R1291 B.n827 B.n18 10.6151
R1292 B.n823 B.n18 10.6151
R1293 B.n823 B.n822 10.6151
R1294 B.n822 B.n821 10.6151
R1295 B.n821 B.n20 10.6151
R1296 B.n817 B.n20 10.6151
R1297 B.n817 B.n816 10.6151
R1298 B.n816 B.n815 10.6151
R1299 B.n815 B.n22 10.6151
R1300 B.n811 B.n22 10.6151
R1301 B.n811 B.n810 10.6151
R1302 B.n810 B.n809 10.6151
R1303 B.n809 B.n24 10.6151
R1304 B.n805 B.n24 10.6151
R1305 B.n805 B.n804 10.6151
R1306 B.n804 B.n803 10.6151
R1307 B.n803 B.n26 10.6151
R1308 B.n799 B.n26 10.6151
R1309 B.n799 B.n798 10.6151
R1310 B.n798 B.n797 10.6151
R1311 B.n719 B.n718 6.5566
R1312 B.n706 B.n62 6.5566
R1313 B.n380 B.n379 6.5566
R1314 B.n392 B.n168 6.5566
R1315 B.n720 B.n719 4.05904
R1316 B.n703 B.n62 4.05904
R1317 B.n379 B.n378 4.05904
R1318 B.n395 B.n168 4.05904
R1319 B.n875 B.n0 2.81026
R1320 B.n875 B.n1 2.81026
R1321 VP.n18 VP.t3 203.644
R1322 VP.n60 VP.t1 169.036
R1323 VP.n44 VP.t7 169.036
R1324 VP.n7 VP.t9 169.036
R1325 VP.n67 VP.t5 169.036
R1326 VP.n75 VP.t6 169.036
R1327 VP.n26 VP.t8 169.036
R1328 VP.n41 VP.t2 169.036
R1329 VP.n33 VP.t4 169.036
R1330 VP.n17 VP.t0 169.036
R1331 VP.n20 VP.n19 161.3
R1332 VP.n21 VP.n16 161.3
R1333 VP.n23 VP.n22 161.3
R1334 VP.n24 VP.n15 161.3
R1335 VP.n26 VP.n25 161.3
R1336 VP.n27 VP.n14 161.3
R1337 VP.n29 VP.n28 161.3
R1338 VP.n30 VP.n13 161.3
R1339 VP.n32 VP.n31 161.3
R1340 VP.n34 VP.n12 161.3
R1341 VP.n36 VP.n35 161.3
R1342 VP.n37 VP.n11 161.3
R1343 VP.n39 VP.n38 161.3
R1344 VP.n40 VP.n10 161.3
R1345 VP.n74 VP.n0 161.3
R1346 VP.n73 VP.n72 161.3
R1347 VP.n71 VP.n1 161.3
R1348 VP.n70 VP.n69 161.3
R1349 VP.n68 VP.n2 161.3
R1350 VP.n66 VP.n65 161.3
R1351 VP.n64 VP.n3 161.3
R1352 VP.n63 VP.n62 161.3
R1353 VP.n61 VP.n4 161.3
R1354 VP.n60 VP.n59 161.3
R1355 VP.n58 VP.n5 161.3
R1356 VP.n57 VP.n56 161.3
R1357 VP.n55 VP.n6 161.3
R1358 VP.n54 VP.n53 161.3
R1359 VP.n52 VP.n51 161.3
R1360 VP.n50 VP.n8 161.3
R1361 VP.n49 VP.n48 161.3
R1362 VP.n47 VP.n9 161.3
R1363 VP.n46 VP.n45 161.3
R1364 VP.n44 VP.n43 88.2837
R1365 VP.n76 VP.n75 88.2837
R1366 VP.n42 VP.n41 88.2837
R1367 VP.n62 VP.n3 56.5617
R1368 VP.n22 VP.n21 56.5617
R1369 VP.n49 VP.n9 56.5617
R1370 VP.n56 VP.n55 56.5617
R1371 VP.n73 VP.n1 56.5617
R1372 VP.n39 VP.n11 56.5617
R1373 VP.n28 VP.n13 56.5617
R1374 VP.n43 VP.n42 53.1057
R1375 VP.n18 VP.n17 47.3938
R1376 VP.n45 VP.n9 24.5923
R1377 VP.n50 VP.n49 24.5923
R1378 VP.n51 VP.n50 24.5923
R1379 VP.n55 VP.n54 24.5923
R1380 VP.n56 VP.n5 24.5923
R1381 VP.n60 VP.n5 24.5923
R1382 VP.n61 VP.n60 24.5923
R1383 VP.n62 VP.n61 24.5923
R1384 VP.n66 VP.n3 24.5923
R1385 VP.n69 VP.n68 24.5923
R1386 VP.n69 VP.n1 24.5923
R1387 VP.n74 VP.n73 24.5923
R1388 VP.n40 VP.n39 24.5923
R1389 VP.n32 VP.n13 24.5923
R1390 VP.n35 VP.n34 24.5923
R1391 VP.n35 VP.n11 24.5923
R1392 VP.n22 VP.n15 24.5923
R1393 VP.n26 VP.n15 24.5923
R1394 VP.n27 VP.n26 24.5923
R1395 VP.n28 VP.n27 24.5923
R1396 VP.n21 VP.n20 24.5923
R1397 VP.n54 VP.n7 23.6087
R1398 VP.n67 VP.n66 23.6087
R1399 VP.n33 VP.n32 23.6087
R1400 VP.n20 VP.n17 23.6087
R1401 VP.n45 VP.n44 22.625
R1402 VP.n75 VP.n74 22.625
R1403 VP.n41 VP.n40 22.625
R1404 VP.n19 VP.n18 8.71357
R1405 VP.n51 VP.n7 0.984173
R1406 VP.n68 VP.n67 0.984173
R1407 VP.n34 VP.n33 0.984173
R1408 VP.n42 VP.n10 0.278335
R1409 VP.n46 VP.n43 0.278335
R1410 VP.n76 VP.n0 0.278335
R1411 VP.n19 VP.n16 0.189894
R1412 VP.n23 VP.n16 0.189894
R1413 VP.n24 VP.n23 0.189894
R1414 VP.n25 VP.n24 0.189894
R1415 VP.n25 VP.n14 0.189894
R1416 VP.n29 VP.n14 0.189894
R1417 VP.n30 VP.n29 0.189894
R1418 VP.n31 VP.n30 0.189894
R1419 VP.n31 VP.n12 0.189894
R1420 VP.n36 VP.n12 0.189894
R1421 VP.n37 VP.n36 0.189894
R1422 VP.n38 VP.n37 0.189894
R1423 VP.n38 VP.n10 0.189894
R1424 VP.n47 VP.n46 0.189894
R1425 VP.n48 VP.n47 0.189894
R1426 VP.n48 VP.n8 0.189894
R1427 VP.n52 VP.n8 0.189894
R1428 VP.n53 VP.n52 0.189894
R1429 VP.n53 VP.n6 0.189894
R1430 VP.n57 VP.n6 0.189894
R1431 VP.n58 VP.n57 0.189894
R1432 VP.n59 VP.n58 0.189894
R1433 VP.n59 VP.n4 0.189894
R1434 VP.n63 VP.n4 0.189894
R1435 VP.n64 VP.n63 0.189894
R1436 VP.n65 VP.n64 0.189894
R1437 VP.n65 VP.n2 0.189894
R1438 VP.n70 VP.n2 0.189894
R1439 VP.n71 VP.n70 0.189894
R1440 VP.n72 VP.n71 0.189894
R1441 VP.n72 VP.n0 0.189894
R1442 VP VP.n76 0.153485
R1443 VDD1.n1 VDD1.t0 76.3501
R1444 VDD1.n3 VDD1.t6 76.3499
R1445 VDD1.n5 VDD1.n4 73.6045
R1446 VDD1.n1 VDD1.n0 72.0567
R1447 VDD1.n7 VDD1.n6 72.0565
R1448 VDD1.n3 VDD1.n2 72.0564
R1449 VDD1.n7 VDD1.n5 48.5224
R1450 VDD1.n6 VDD1.t1 2.156
R1451 VDD1.n6 VDD1.t8 2.156
R1452 VDD1.n0 VDD1.t4 2.156
R1453 VDD1.n0 VDD1.t9 2.156
R1454 VDD1.n4 VDD1.t5 2.156
R1455 VDD1.n4 VDD1.t2 2.156
R1456 VDD1.n2 VDD1.t7 2.156
R1457 VDD1.n2 VDD1.t3 2.156
R1458 VDD1 VDD1.n7 1.54576
R1459 VDD1 VDD1.n1 0.593172
R1460 VDD1.n5 VDD1.n3 0.479637
R1461 VTAIL.n11 VTAIL.t6 57.5334
R1462 VTAIL.n17 VTAIL.t7 57.5331
R1463 VTAIL.n2 VTAIL.t13 57.5331
R1464 VTAIL.n16 VTAIL.t17 57.5331
R1465 VTAIL.n15 VTAIL.n14 55.3779
R1466 VTAIL.n13 VTAIL.n12 55.3779
R1467 VTAIL.n10 VTAIL.n9 55.3779
R1468 VTAIL.n8 VTAIL.n7 55.3779
R1469 VTAIL.n19 VTAIL.n18 55.3776
R1470 VTAIL.n1 VTAIL.n0 55.3776
R1471 VTAIL.n4 VTAIL.n3 55.3776
R1472 VTAIL.n6 VTAIL.n5 55.3776
R1473 VTAIL.n8 VTAIL.n6 29.6427
R1474 VTAIL.n17 VTAIL.n16 27.5048
R1475 VTAIL.n18 VTAIL.t3 2.156
R1476 VTAIL.n18 VTAIL.t5 2.156
R1477 VTAIL.n0 VTAIL.t2 2.156
R1478 VTAIL.n0 VTAIL.t9 2.156
R1479 VTAIL.n3 VTAIL.t18 2.156
R1480 VTAIL.n3 VTAIL.t14 2.156
R1481 VTAIL.n5 VTAIL.t12 2.156
R1482 VTAIL.n5 VTAIL.t10 2.156
R1483 VTAIL.n14 VTAIL.t11 2.156
R1484 VTAIL.n14 VTAIL.t15 2.156
R1485 VTAIL.n12 VTAIL.t16 2.156
R1486 VTAIL.n12 VTAIL.t19 2.156
R1487 VTAIL.n9 VTAIL.t8 2.156
R1488 VTAIL.n9 VTAIL.t1 2.156
R1489 VTAIL.n7 VTAIL.t4 2.156
R1490 VTAIL.n7 VTAIL.t0 2.156
R1491 VTAIL.n10 VTAIL.n8 2.13843
R1492 VTAIL.n11 VTAIL.n10 2.13843
R1493 VTAIL.n15 VTAIL.n13 2.13843
R1494 VTAIL.n16 VTAIL.n15 2.13843
R1495 VTAIL.n6 VTAIL.n4 2.13843
R1496 VTAIL.n4 VTAIL.n2 2.13843
R1497 VTAIL.n19 VTAIL.n17 2.13843
R1498 VTAIL VTAIL.n1 1.66214
R1499 VTAIL.n13 VTAIL.n11 1.53929
R1500 VTAIL.n2 VTAIL.n1 1.53929
R1501 VTAIL VTAIL.n19 0.476793
R1502 VN.n8 VN.t8 203.644
R1503 VN.n41 VN.t3 203.644
R1504 VN.n16 VN.t6 169.036
R1505 VN.n7 VN.t7 169.036
R1506 VN.n23 VN.t4 169.036
R1507 VN.n31 VN.t1 169.036
R1508 VN.n49 VN.t0 169.036
R1509 VN.n40 VN.t2 169.036
R1510 VN.n56 VN.t9 169.036
R1511 VN.n64 VN.t5 169.036
R1512 VN.n63 VN.n33 161.3
R1513 VN.n62 VN.n61 161.3
R1514 VN.n60 VN.n34 161.3
R1515 VN.n59 VN.n58 161.3
R1516 VN.n57 VN.n35 161.3
R1517 VN.n55 VN.n54 161.3
R1518 VN.n53 VN.n36 161.3
R1519 VN.n52 VN.n51 161.3
R1520 VN.n50 VN.n37 161.3
R1521 VN.n49 VN.n48 161.3
R1522 VN.n47 VN.n38 161.3
R1523 VN.n46 VN.n45 161.3
R1524 VN.n44 VN.n39 161.3
R1525 VN.n43 VN.n42 161.3
R1526 VN.n30 VN.n0 161.3
R1527 VN.n29 VN.n28 161.3
R1528 VN.n27 VN.n1 161.3
R1529 VN.n26 VN.n25 161.3
R1530 VN.n24 VN.n2 161.3
R1531 VN.n22 VN.n21 161.3
R1532 VN.n20 VN.n3 161.3
R1533 VN.n19 VN.n18 161.3
R1534 VN.n17 VN.n4 161.3
R1535 VN.n16 VN.n15 161.3
R1536 VN.n14 VN.n5 161.3
R1537 VN.n13 VN.n12 161.3
R1538 VN.n11 VN.n6 161.3
R1539 VN.n10 VN.n9 161.3
R1540 VN.n32 VN.n31 88.2837
R1541 VN.n65 VN.n64 88.2837
R1542 VN.n18 VN.n3 56.5617
R1543 VN.n51 VN.n36 56.5617
R1544 VN.n12 VN.n11 56.5617
R1545 VN.n29 VN.n1 56.5617
R1546 VN.n45 VN.n44 56.5617
R1547 VN.n62 VN.n34 56.5617
R1548 VN VN.n65 53.3845
R1549 VN.n8 VN.n7 47.3938
R1550 VN.n41 VN.n40 47.3938
R1551 VN.n11 VN.n10 24.5923
R1552 VN.n12 VN.n5 24.5923
R1553 VN.n16 VN.n5 24.5923
R1554 VN.n17 VN.n16 24.5923
R1555 VN.n18 VN.n17 24.5923
R1556 VN.n22 VN.n3 24.5923
R1557 VN.n25 VN.n24 24.5923
R1558 VN.n25 VN.n1 24.5923
R1559 VN.n30 VN.n29 24.5923
R1560 VN.n44 VN.n43 24.5923
R1561 VN.n51 VN.n50 24.5923
R1562 VN.n50 VN.n49 24.5923
R1563 VN.n49 VN.n38 24.5923
R1564 VN.n45 VN.n38 24.5923
R1565 VN.n58 VN.n34 24.5923
R1566 VN.n58 VN.n57 24.5923
R1567 VN.n55 VN.n36 24.5923
R1568 VN.n63 VN.n62 24.5923
R1569 VN.n10 VN.n7 23.6087
R1570 VN.n23 VN.n22 23.6087
R1571 VN.n43 VN.n40 23.6087
R1572 VN.n56 VN.n55 23.6087
R1573 VN.n31 VN.n30 22.625
R1574 VN.n64 VN.n63 22.625
R1575 VN.n42 VN.n41 8.71357
R1576 VN.n9 VN.n8 8.71357
R1577 VN.n24 VN.n23 0.984173
R1578 VN.n57 VN.n56 0.984173
R1579 VN.n65 VN.n33 0.278335
R1580 VN.n32 VN.n0 0.278335
R1581 VN.n61 VN.n33 0.189894
R1582 VN.n61 VN.n60 0.189894
R1583 VN.n60 VN.n59 0.189894
R1584 VN.n59 VN.n35 0.189894
R1585 VN.n54 VN.n35 0.189894
R1586 VN.n54 VN.n53 0.189894
R1587 VN.n53 VN.n52 0.189894
R1588 VN.n52 VN.n37 0.189894
R1589 VN.n48 VN.n37 0.189894
R1590 VN.n48 VN.n47 0.189894
R1591 VN.n47 VN.n46 0.189894
R1592 VN.n46 VN.n39 0.189894
R1593 VN.n42 VN.n39 0.189894
R1594 VN.n9 VN.n6 0.189894
R1595 VN.n13 VN.n6 0.189894
R1596 VN.n14 VN.n13 0.189894
R1597 VN.n15 VN.n14 0.189894
R1598 VN.n15 VN.n4 0.189894
R1599 VN.n19 VN.n4 0.189894
R1600 VN.n20 VN.n19 0.189894
R1601 VN.n21 VN.n20 0.189894
R1602 VN.n21 VN.n2 0.189894
R1603 VN.n26 VN.n2 0.189894
R1604 VN.n27 VN.n26 0.189894
R1605 VN.n28 VN.n27 0.189894
R1606 VN.n28 VN.n0 0.189894
R1607 VN VN.n32 0.153485
R1608 VDD2.n1 VDD2.t1 76.3499
R1609 VDD2.n4 VDD2.t4 74.2122
R1610 VDD2.n3 VDD2.n2 73.6045
R1611 VDD2 VDD2.n7 73.6017
R1612 VDD2.n6 VDD2.n5 72.0567
R1613 VDD2.n1 VDD2.n0 72.0564
R1614 VDD2.n4 VDD2.n3 46.8705
R1615 VDD2.n7 VDD2.t7 2.156
R1616 VDD2.n7 VDD2.t6 2.156
R1617 VDD2.n5 VDD2.t0 2.156
R1618 VDD2.n5 VDD2.t9 2.156
R1619 VDD2.n2 VDD2.t5 2.156
R1620 VDD2.n2 VDD2.t8 2.156
R1621 VDD2.n0 VDD2.t2 2.156
R1622 VDD2.n0 VDD2.t3 2.156
R1623 VDD2.n6 VDD2.n4 2.13843
R1624 VDD2 VDD2.n6 0.593172
R1625 VDD2.n3 VDD2.n1 0.479637
C0 VN VDD1 0.152815f
C1 VP VTAIL 13.065599f
C2 B w_n3946_n3984# 10.653599f
C3 VDD1 w_n3946_n3984# 2.8363f
C4 VN VDD2 12.728701f
C5 B VTAIL 4.20183f
C6 VP B 2.06756f
C7 VDD1 VTAIL 11.9593f
C8 VP VDD1 13.0983f
C9 VDD2 w_n3946_n3984# 2.95655f
C10 VN w_n3946_n3984# 8.338039f
C11 VDD2 VTAIL 12.0058f
C12 VP VDD2 0.526961f
C13 B VDD1 2.54407f
C14 VN VTAIL 13.0513f
C15 VP VN 8.296849f
C16 VDD2 B 2.64446f
C17 w_n3946_n3984# VTAIL 3.59481f
C18 VP w_n3946_n3984# 8.850401f
C19 VDD2 VDD1 1.8831f
C20 VN B 1.20848f
C21 VDD2 VSUBS 2.01609f
C22 VDD1 VSUBS 1.847866f
C23 VTAIL VSUBS 1.299601f
C24 VN VSUBS 7.08113f
C25 VP VSUBS 3.787038f
C26 B VSUBS 5.067826f
C27 w_n3946_n3984# VSUBS 0.19277p
C28 VDD2.t1 VSUBS 3.42418f
C29 VDD2.t2 VSUBS 0.321549f
C30 VDD2.t3 VSUBS 0.321549f
C31 VDD2.n0 VSUBS 2.61697f
C32 VDD2.n1 VSUBS 1.51789f
C33 VDD2.t5 VSUBS 0.321549f
C34 VDD2.t8 VSUBS 0.321549f
C35 VDD2.n2 VSUBS 2.6347f
C36 VDD2.n3 VSUBS 3.37289f
C37 VDD2.t4 VSUBS 3.40178f
C38 VDD2.n4 VSUBS 3.7483f
C39 VDD2.t0 VSUBS 0.321549f
C40 VDD2.t9 VSUBS 0.321549f
C41 VDD2.n5 VSUBS 2.61697f
C42 VDD2.n6 VSUBS 0.748686f
C43 VDD2.t7 VSUBS 0.321549f
C44 VDD2.t6 VSUBS 0.321549f
C45 VDD2.n7 VSUBS 2.63465f
C46 VN.n0 VSUBS 0.038831f
C47 VN.t1 VSUBS 2.61718f
C48 VN.n1 VSUBS 0.040373f
C49 VN.n2 VSUBS 0.029455f
C50 VN.t4 VSUBS 2.61718f
C51 VN.n3 VSUBS 0.043632f
C52 VN.n4 VSUBS 0.029455f
C53 VN.t6 VSUBS 2.61718f
C54 VN.n5 VSUBS 0.054622f
C55 VN.n6 VSUBS 0.029455f
C56 VN.t7 VSUBS 2.61718f
C57 VN.n7 VSUBS 1.00697f
C58 VN.t8 VSUBS 2.80124f
C59 VN.n8 VSUBS 0.980957f
C60 VN.n9 VSUBS 0.248798f
C61 VN.n10 VSUBS 0.053543f
C62 VN.n11 VSUBS 0.043632f
C63 VN.n12 VSUBS 0.042003f
C64 VN.n13 VSUBS 0.029455f
C65 VN.n14 VSUBS 0.029455f
C66 VN.n15 VSUBS 0.029455f
C67 VN.n16 VSUBS 0.946736f
C68 VN.n17 VSUBS 0.054622f
C69 VN.n18 VSUBS 0.042003f
C70 VN.n19 VSUBS 0.029455f
C71 VN.n20 VSUBS 0.029455f
C72 VN.n21 VSUBS 0.029455f
C73 VN.n22 VSUBS 0.053543f
C74 VN.n23 VSUBS 0.919079f
C75 VN.n24 VSUBS 0.028735f
C76 VN.n25 VSUBS 0.054622f
C77 VN.n26 VSUBS 0.029455f
C78 VN.n27 VSUBS 0.029455f
C79 VN.n28 VSUBS 0.029455f
C80 VN.n29 VSUBS 0.045262f
C81 VN.n30 VSUBS 0.052465f
C82 VN.n31 VSUBS 1.02065f
C83 VN.n32 VSUBS 0.033798f
C84 VN.n33 VSUBS 0.038831f
C85 VN.t5 VSUBS 2.61718f
C86 VN.n34 VSUBS 0.040373f
C87 VN.n35 VSUBS 0.029455f
C88 VN.t9 VSUBS 2.61718f
C89 VN.n36 VSUBS 0.043632f
C90 VN.n37 VSUBS 0.029455f
C91 VN.t0 VSUBS 2.61718f
C92 VN.n38 VSUBS 0.054622f
C93 VN.n39 VSUBS 0.029455f
C94 VN.t2 VSUBS 2.61718f
C95 VN.n40 VSUBS 1.00697f
C96 VN.t3 VSUBS 2.80124f
C97 VN.n41 VSUBS 0.980957f
C98 VN.n42 VSUBS 0.248798f
C99 VN.n43 VSUBS 0.053543f
C100 VN.n44 VSUBS 0.043632f
C101 VN.n45 VSUBS 0.042003f
C102 VN.n46 VSUBS 0.029455f
C103 VN.n47 VSUBS 0.029455f
C104 VN.n48 VSUBS 0.029455f
C105 VN.n49 VSUBS 0.946736f
C106 VN.n50 VSUBS 0.054622f
C107 VN.n51 VSUBS 0.042003f
C108 VN.n52 VSUBS 0.029455f
C109 VN.n53 VSUBS 0.029455f
C110 VN.n54 VSUBS 0.029455f
C111 VN.n55 VSUBS 0.053543f
C112 VN.n56 VSUBS 0.919079f
C113 VN.n57 VSUBS 0.028735f
C114 VN.n58 VSUBS 0.054622f
C115 VN.n59 VSUBS 0.029455f
C116 VN.n60 VSUBS 0.029455f
C117 VN.n61 VSUBS 0.029455f
C118 VN.n62 VSUBS 0.045262f
C119 VN.n63 VSUBS 0.052465f
C120 VN.n64 VSUBS 1.02065f
C121 VN.n65 VSUBS 1.79047f
C122 VTAIL.t2 VSUBS 0.330886f
C123 VTAIL.t9 VSUBS 0.330886f
C124 VTAIL.n0 VSUBS 2.53609f
C125 VTAIL.n1 VSUBS 0.931592f
C126 VTAIL.t13 VSUBS 3.32208f
C127 VTAIL.n2 VSUBS 1.09064f
C128 VTAIL.t18 VSUBS 0.330886f
C129 VTAIL.t14 VSUBS 0.330886f
C130 VTAIL.n3 VSUBS 2.53609f
C131 VTAIL.n4 VSUBS 1.02781f
C132 VTAIL.t12 VSUBS 0.330886f
C133 VTAIL.t10 VSUBS 0.330886f
C134 VTAIL.n5 VSUBS 2.53609f
C135 VTAIL.n6 VSUBS 2.75938f
C136 VTAIL.t4 VSUBS 0.330886f
C137 VTAIL.t0 VSUBS 0.330886f
C138 VTAIL.n7 VSUBS 2.5361f
C139 VTAIL.n8 VSUBS 2.75938f
C140 VTAIL.t8 VSUBS 0.330886f
C141 VTAIL.t1 VSUBS 0.330886f
C142 VTAIL.n9 VSUBS 2.5361f
C143 VTAIL.n10 VSUBS 1.02781f
C144 VTAIL.t6 VSUBS 3.32209f
C145 VTAIL.n11 VSUBS 1.09063f
C146 VTAIL.t16 VSUBS 0.330886f
C147 VTAIL.t19 VSUBS 0.330886f
C148 VTAIL.n12 VSUBS 2.5361f
C149 VTAIL.n13 VSUBS 0.974201f
C150 VTAIL.t11 VSUBS 0.330886f
C151 VTAIL.t15 VSUBS 0.330886f
C152 VTAIL.n14 VSUBS 2.5361f
C153 VTAIL.n15 VSUBS 1.02781f
C154 VTAIL.t17 VSUBS 3.32208f
C155 VTAIL.n16 VSUBS 2.68453f
C156 VTAIL.t7 VSUBS 3.32208f
C157 VTAIL.n17 VSUBS 2.68453f
C158 VTAIL.t3 VSUBS 0.330886f
C159 VTAIL.t5 VSUBS 0.330886f
C160 VTAIL.n18 VSUBS 2.53609f
C161 VTAIL.n19 VSUBS 0.879144f
C162 VDD1.t0 VSUBS 3.42423f
C163 VDD1.t4 VSUBS 0.321552f
C164 VDD1.t9 VSUBS 0.321552f
C165 VDD1.n0 VSUBS 2.617f
C166 VDD1.n1 VSUBS 1.52646f
C167 VDD1.t6 VSUBS 3.42422f
C168 VDD1.t7 VSUBS 0.321552f
C169 VDD1.t3 VSUBS 0.321552f
C170 VDD1.n2 VSUBS 2.617f
C171 VDD1.n3 VSUBS 1.5179f
C172 VDD1.t5 VSUBS 0.321552f
C173 VDD1.t2 VSUBS 0.321552f
C174 VDD1.n4 VSUBS 2.63473f
C175 VDD1.n5 VSUBS 3.49694f
C176 VDD1.t1 VSUBS 0.321552f
C177 VDD1.t8 VSUBS 0.321552f
C178 VDD1.n6 VSUBS 2.61699f
C179 VDD1.n7 VSUBS 3.76621f
C180 VP.n0 VSUBS 0.041711f
C181 VP.t6 VSUBS 2.81128f
C182 VP.n1 VSUBS 0.043367f
C183 VP.n2 VSUBS 0.03164f
C184 VP.t5 VSUBS 2.81128f
C185 VP.n3 VSUBS 0.046868f
C186 VP.n4 VSUBS 0.03164f
C187 VP.t1 VSUBS 2.81128f
C188 VP.n5 VSUBS 0.058673f
C189 VP.n6 VSUBS 0.03164f
C190 VP.t9 VSUBS 2.81128f
C191 VP.n7 VSUBS 0.98724f
C192 VP.n8 VSUBS 0.03164f
C193 VP.n9 VSUBS 0.048619f
C194 VP.n10 VSUBS 0.041711f
C195 VP.t2 VSUBS 2.81128f
C196 VP.n11 VSUBS 0.043367f
C197 VP.n12 VSUBS 0.03164f
C198 VP.t4 VSUBS 2.81128f
C199 VP.n13 VSUBS 0.046868f
C200 VP.n14 VSUBS 0.03164f
C201 VP.t8 VSUBS 2.81128f
C202 VP.n15 VSUBS 0.058673f
C203 VP.n16 VSUBS 0.03164f
C204 VP.t0 VSUBS 2.81128f
C205 VP.n17 VSUBS 1.08165f
C206 VP.t3 VSUBS 3.00899f
C207 VP.n18 VSUBS 1.05371f
C208 VP.n19 VSUBS 0.267249f
C209 VP.n20 VSUBS 0.057514f
C210 VP.n21 VSUBS 0.046868f
C211 VP.n22 VSUBS 0.045118f
C212 VP.n23 VSUBS 0.03164f
C213 VP.n24 VSUBS 0.03164f
C214 VP.n25 VSUBS 0.03164f
C215 VP.n26 VSUBS 1.01695f
C216 VP.n27 VSUBS 0.058673f
C217 VP.n28 VSUBS 0.045118f
C218 VP.n29 VSUBS 0.03164f
C219 VP.n30 VSUBS 0.03164f
C220 VP.n31 VSUBS 0.03164f
C221 VP.n32 VSUBS 0.057514f
C222 VP.n33 VSUBS 0.98724f
C223 VP.n34 VSUBS 0.030866f
C224 VP.n35 VSUBS 0.058673f
C225 VP.n36 VSUBS 0.03164f
C226 VP.n37 VSUBS 0.03164f
C227 VP.n38 VSUBS 0.03164f
C228 VP.n39 VSUBS 0.048619f
C229 VP.n40 VSUBS 0.056355f
C230 VP.n41 VSUBS 1.09634f
C231 VP.n42 VSUBS 1.90641f
C232 VP.n43 VSUBS 1.92789f
C233 VP.t7 VSUBS 2.81128f
C234 VP.n44 VSUBS 1.09634f
C235 VP.n45 VSUBS 0.056355f
C236 VP.n46 VSUBS 0.041711f
C237 VP.n47 VSUBS 0.03164f
C238 VP.n48 VSUBS 0.03164f
C239 VP.n49 VSUBS 0.043367f
C240 VP.n50 VSUBS 0.058673f
C241 VP.n51 VSUBS 0.030866f
C242 VP.n52 VSUBS 0.03164f
C243 VP.n53 VSUBS 0.03164f
C244 VP.n54 VSUBS 0.057514f
C245 VP.n55 VSUBS 0.046868f
C246 VP.n56 VSUBS 0.045118f
C247 VP.n57 VSUBS 0.03164f
C248 VP.n58 VSUBS 0.03164f
C249 VP.n59 VSUBS 0.03164f
C250 VP.n60 VSUBS 1.01695f
C251 VP.n61 VSUBS 0.058673f
C252 VP.n62 VSUBS 0.045118f
C253 VP.n63 VSUBS 0.03164f
C254 VP.n64 VSUBS 0.03164f
C255 VP.n65 VSUBS 0.03164f
C256 VP.n66 VSUBS 0.057514f
C257 VP.n67 VSUBS 0.98724f
C258 VP.n68 VSUBS 0.030866f
C259 VP.n69 VSUBS 0.058673f
C260 VP.n70 VSUBS 0.03164f
C261 VP.n71 VSUBS 0.03164f
C262 VP.n72 VSUBS 0.03164f
C263 VP.n73 VSUBS 0.048619f
C264 VP.n74 VSUBS 0.056355f
C265 VP.n75 VSUBS 1.09634f
C266 VP.n76 VSUBS 0.036305f
C267 B.n0 VSUBS 0.00562f
C268 B.n1 VSUBS 0.00562f
C269 B.n2 VSUBS 0.008887f
C270 B.n3 VSUBS 0.008887f
C271 B.n4 VSUBS 0.008887f
C272 B.n5 VSUBS 0.008887f
C273 B.n6 VSUBS 0.008887f
C274 B.n7 VSUBS 0.008887f
C275 B.n8 VSUBS 0.008887f
C276 B.n9 VSUBS 0.008887f
C277 B.n10 VSUBS 0.008887f
C278 B.n11 VSUBS 0.008887f
C279 B.n12 VSUBS 0.008887f
C280 B.n13 VSUBS 0.008887f
C281 B.n14 VSUBS 0.008887f
C282 B.n15 VSUBS 0.008887f
C283 B.n16 VSUBS 0.008887f
C284 B.n17 VSUBS 0.008887f
C285 B.n18 VSUBS 0.008887f
C286 B.n19 VSUBS 0.008887f
C287 B.n20 VSUBS 0.008887f
C288 B.n21 VSUBS 0.008887f
C289 B.n22 VSUBS 0.008887f
C290 B.n23 VSUBS 0.008887f
C291 B.n24 VSUBS 0.008887f
C292 B.n25 VSUBS 0.008887f
C293 B.n26 VSUBS 0.008887f
C294 B.n27 VSUBS 0.008887f
C295 B.n28 VSUBS 0.020445f
C296 B.n29 VSUBS 0.008887f
C297 B.n30 VSUBS 0.008887f
C298 B.n31 VSUBS 0.008887f
C299 B.n32 VSUBS 0.008887f
C300 B.n33 VSUBS 0.008887f
C301 B.n34 VSUBS 0.008887f
C302 B.n35 VSUBS 0.008887f
C303 B.n36 VSUBS 0.008887f
C304 B.n37 VSUBS 0.008887f
C305 B.n38 VSUBS 0.008887f
C306 B.n39 VSUBS 0.008887f
C307 B.n40 VSUBS 0.008887f
C308 B.n41 VSUBS 0.008887f
C309 B.n42 VSUBS 0.008887f
C310 B.n43 VSUBS 0.008887f
C311 B.n44 VSUBS 0.008887f
C312 B.n45 VSUBS 0.008887f
C313 B.n46 VSUBS 0.008887f
C314 B.n47 VSUBS 0.008887f
C315 B.n48 VSUBS 0.008887f
C316 B.n49 VSUBS 0.008887f
C317 B.n50 VSUBS 0.008887f
C318 B.n51 VSUBS 0.008887f
C319 B.n52 VSUBS 0.008887f
C320 B.n53 VSUBS 0.008887f
C321 B.t8 VSUBS 0.637644f
C322 B.t7 VSUBS 0.661042f
C323 B.t6 VSUBS 1.82198f
C324 B.n54 VSUBS 0.331055f
C325 B.n55 VSUBS 0.08903f
C326 B.n56 VSUBS 0.008887f
C327 B.n57 VSUBS 0.008887f
C328 B.n58 VSUBS 0.008887f
C329 B.n59 VSUBS 0.008887f
C330 B.t11 VSUBS 0.637626f
C331 B.t10 VSUBS 0.661026f
C332 B.t9 VSUBS 1.82198f
C333 B.n60 VSUBS 0.33107f
C334 B.n61 VSUBS 0.089048f
C335 B.n62 VSUBS 0.020591f
C336 B.n63 VSUBS 0.008887f
C337 B.n64 VSUBS 0.008887f
C338 B.n65 VSUBS 0.008887f
C339 B.n66 VSUBS 0.008887f
C340 B.n67 VSUBS 0.008887f
C341 B.n68 VSUBS 0.008887f
C342 B.n69 VSUBS 0.008887f
C343 B.n70 VSUBS 0.008887f
C344 B.n71 VSUBS 0.008887f
C345 B.n72 VSUBS 0.008887f
C346 B.n73 VSUBS 0.008887f
C347 B.n74 VSUBS 0.008887f
C348 B.n75 VSUBS 0.008887f
C349 B.n76 VSUBS 0.008887f
C350 B.n77 VSUBS 0.008887f
C351 B.n78 VSUBS 0.008887f
C352 B.n79 VSUBS 0.008887f
C353 B.n80 VSUBS 0.008887f
C354 B.n81 VSUBS 0.008887f
C355 B.n82 VSUBS 0.008887f
C356 B.n83 VSUBS 0.008887f
C357 B.n84 VSUBS 0.008887f
C358 B.n85 VSUBS 0.008887f
C359 B.n86 VSUBS 0.008887f
C360 B.n87 VSUBS 0.008887f
C361 B.n88 VSUBS 0.020663f
C362 B.n89 VSUBS 0.008887f
C363 B.n90 VSUBS 0.008887f
C364 B.n91 VSUBS 0.008887f
C365 B.n92 VSUBS 0.008887f
C366 B.n93 VSUBS 0.008887f
C367 B.n94 VSUBS 0.008887f
C368 B.n95 VSUBS 0.008887f
C369 B.n96 VSUBS 0.008887f
C370 B.n97 VSUBS 0.008887f
C371 B.n98 VSUBS 0.008887f
C372 B.n99 VSUBS 0.008887f
C373 B.n100 VSUBS 0.008887f
C374 B.n101 VSUBS 0.008887f
C375 B.n102 VSUBS 0.008887f
C376 B.n103 VSUBS 0.008887f
C377 B.n104 VSUBS 0.008887f
C378 B.n105 VSUBS 0.008887f
C379 B.n106 VSUBS 0.008887f
C380 B.n107 VSUBS 0.008887f
C381 B.n108 VSUBS 0.008887f
C382 B.n109 VSUBS 0.008887f
C383 B.n110 VSUBS 0.008887f
C384 B.n111 VSUBS 0.008887f
C385 B.n112 VSUBS 0.008887f
C386 B.n113 VSUBS 0.008887f
C387 B.n114 VSUBS 0.008887f
C388 B.n115 VSUBS 0.008887f
C389 B.n116 VSUBS 0.008887f
C390 B.n117 VSUBS 0.008887f
C391 B.n118 VSUBS 0.008887f
C392 B.n119 VSUBS 0.008887f
C393 B.n120 VSUBS 0.008887f
C394 B.n121 VSUBS 0.008887f
C395 B.n122 VSUBS 0.008887f
C396 B.n123 VSUBS 0.008887f
C397 B.n124 VSUBS 0.008887f
C398 B.n125 VSUBS 0.008887f
C399 B.n126 VSUBS 0.008887f
C400 B.n127 VSUBS 0.008887f
C401 B.n128 VSUBS 0.008887f
C402 B.n129 VSUBS 0.008887f
C403 B.n130 VSUBS 0.008887f
C404 B.n131 VSUBS 0.008887f
C405 B.n132 VSUBS 0.008887f
C406 B.n133 VSUBS 0.008887f
C407 B.n134 VSUBS 0.008887f
C408 B.n135 VSUBS 0.008887f
C409 B.n136 VSUBS 0.008887f
C410 B.n137 VSUBS 0.008887f
C411 B.n138 VSUBS 0.008887f
C412 B.n139 VSUBS 0.008887f
C413 B.n140 VSUBS 0.019548f
C414 B.n141 VSUBS 0.008887f
C415 B.n142 VSUBS 0.008887f
C416 B.n143 VSUBS 0.008887f
C417 B.n144 VSUBS 0.008887f
C418 B.n145 VSUBS 0.008887f
C419 B.n146 VSUBS 0.008887f
C420 B.n147 VSUBS 0.008887f
C421 B.n148 VSUBS 0.008887f
C422 B.n149 VSUBS 0.008887f
C423 B.n150 VSUBS 0.008887f
C424 B.n151 VSUBS 0.008887f
C425 B.n152 VSUBS 0.008887f
C426 B.n153 VSUBS 0.008887f
C427 B.n154 VSUBS 0.008887f
C428 B.n155 VSUBS 0.008887f
C429 B.n156 VSUBS 0.008887f
C430 B.n157 VSUBS 0.008887f
C431 B.n158 VSUBS 0.008887f
C432 B.n159 VSUBS 0.008887f
C433 B.n160 VSUBS 0.008887f
C434 B.n161 VSUBS 0.008887f
C435 B.n162 VSUBS 0.008887f
C436 B.n163 VSUBS 0.008887f
C437 B.n164 VSUBS 0.008887f
C438 B.n165 VSUBS 0.008887f
C439 B.t4 VSUBS 0.637626f
C440 B.t5 VSUBS 0.661026f
C441 B.t3 VSUBS 1.82198f
C442 B.n166 VSUBS 0.33107f
C443 B.n167 VSUBS 0.089048f
C444 B.n168 VSUBS 0.020591f
C445 B.n169 VSUBS 0.008887f
C446 B.n170 VSUBS 0.008887f
C447 B.n171 VSUBS 0.008887f
C448 B.n172 VSUBS 0.008887f
C449 B.n173 VSUBS 0.008887f
C450 B.t1 VSUBS 0.637644f
C451 B.t2 VSUBS 0.661042f
C452 B.t0 VSUBS 1.82198f
C453 B.n174 VSUBS 0.331055f
C454 B.n175 VSUBS 0.08903f
C455 B.n176 VSUBS 0.008887f
C456 B.n177 VSUBS 0.008887f
C457 B.n178 VSUBS 0.008887f
C458 B.n179 VSUBS 0.008887f
C459 B.n180 VSUBS 0.008887f
C460 B.n181 VSUBS 0.008887f
C461 B.n182 VSUBS 0.008887f
C462 B.n183 VSUBS 0.008887f
C463 B.n184 VSUBS 0.008887f
C464 B.n185 VSUBS 0.008887f
C465 B.n186 VSUBS 0.008887f
C466 B.n187 VSUBS 0.008887f
C467 B.n188 VSUBS 0.008887f
C468 B.n189 VSUBS 0.008887f
C469 B.n190 VSUBS 0.008887f
C470 B.n191 VSUBS 0.008887f
C471 B.n192 VSUBS 0.008887f
C472 B.n193 VSUBS 0.008887f
C473 B.n194 VSUBS 0.008887f
C474 B.n195 VSUBS 0.008887f
C475 B.n196 VSUBS 0.008887f
C476 B.n197 VSUBS 0.008887f
C477 B.n198 VSUBS 0.008887f
C478 B.n199 VSUBS 0.008887f
C479 B.n200 VSUBS 0.020445f
C480 B.n201 VSUBS 0.008887f
C481 B.n202 VSUBS 0.008887f
C482 B.n203 VSUBS 0.008887f
C483 B.n204 VSUBS 0.008887f
C484 B.n205 VSUBS 0.008887f
C485 B.n206 VSUBS 0.008887f
C486 B.n207 VSUBS 0.008887f
C487 B.n208 VSUBS 0.008887f
C488 B.n209 VSUBS 0.008887f
C489 B.n210 VSUBS 0.008887f
C490 B.n211 VSUBS 0.008887f
C491 B.n212 VSUBS 0.008887f
C492 B.n213 VSUBS 0.008887f
C493 B.n214 VSUBS 0.008887f
C494 B.n215 VSUBS 0.008887f
C495 B.n216 VSUBS 0.008887f
C496 B.n217 VSUBS 0.008887f
C497 B.n218 VSUBS 0.008887f
C498 B.n219 VSUBS 0.008887f
C499 B.n220 VSUBS 0.008887f
C500 B.n221 VSUBS 0.008887f
C501 B.n222 VSUBS 0.008887f
C502 B.n223 VSUBS 0.008887f
C503 B.n224 VSUBS 0.008887f
C504 B.n225 VSUBS 0.008887f
C505 B.n226 VSUBS 0.008887f
C506 B.n227 VSUBS 0.008887f
C507 B.n228 VSUBS 0.008887f
C508 B.n229 VSUBS 0.008887f
C509 B.n230 VSUBS 0.008887f
C510 B.n231 VSUBS 0.008887f
C511 B.n232 VSUBS 0.008887f
C512 B.n233 VSUBS 0.008887f
C513 B.n234 VSUBS 0.008887f
C514 B.n235 VSUBS 0.008887f
C515 B.n236 VSUBS 0.008887f
C516 B.n237 VSUBS 0.008887f
C517 B.n238 VSUBS 0.008887f
C518 B.n239 VSUBS 0.008887f
C519 B.n240 VSUBS 0.008887f
C520 B.n241 VSUBS 0.008887f
C521 B.n242 VSUBS 0.008887f
C522 B.n243 VSUBS 0.008887f
C523 B.n244 VSUBS 0.008887f
C524 B.n245 VSUBS 0.008887f
C525 B.n246 VSUBS 0.008887f
C526 B.n247 VSUBS 0.008887f
C527 B.n248 VSUBS 0.008887f
C528 B.n249 VSUBS 0.008887f
C529 B.n250 VSUBS 0.008887f
C530 B.n251 VSUBS 0.008887f
C531 B.n252 VSUBS 0.008887f
C532 B.n253 VSUBS 0.008887f
C533 B.n254 VSUBS 0.008887f
C534 B.n255 VSUBS 0.008887f
C535 B.n256 VSUBS 0.008887f
C536 B.n257 VSUBS 0.008887f
C537 B.n258 VSUBS 0.008887f
C538 B.n259 VSUBS 0.008887f
C539 B.n260 VSUBS 0.008887f
C540 B.n261 VSUBS 0.008887f
C541 B.n262 VSUBS 0.008887f
C542 B.n263 VSUBS 0.008887f
C543 B.n264 VSUBS 0.008887f
C544 B.n265 VSUBS 0.008887f
C545 B.n266 VSUBS 0.008887f
C546 B.n267 VSUBS 0.008887f
C547 B.n268 VSUBS 0.008887f
C548 B.n269 VSUBS 0.008887f
C549 B.n270 VSUBS 0.008887f
C550 B.n271 VSUBS 0.008887f
C551 B.n272 VSUBS 0.008887f
C552 B.n273 VSUBS 0.008887f
C553 B.n274 VSUBS 0.008887f
C554 B.n275 VSUBS 0.008887f
C555 B.n276 VSUBS 0.008887f
C556 B.n277 VSUBS 0.008887f
C557 B.n278 VSUBS 0.008887f
C558 B.n279 VSUBS 0.008887f
C559 B.n280 VSUBS 0.008887f
C560 B.n281 VSUBS 0.008887f
C561 B.n282 VSUBS 0.008887f
C562 B.n283 VSUBS 0.008887f
C563 B.n284 VSUBS 0.008887f
C564 B.n285 VSUBS 0.008887f
C565 B.n286 VSUBS 0.008887f
C566 B.n287 VSUBS 0.008887f
C567 B.n288 VSUBS 0.008887f
C568 B.n289 VSUBS 0.008887f
C569 B.n290 VSUBS 0.008887f
C570 B.n291 VSUBS 0.008887f
C571 B.n292 VSUBS 0.008887f
C572 B.n293 VSUBS 0.008887f
C573 B.n294 VSUBS 0.008887f
C574 B.n295 VSUBS 0.008887f
C575 B.n296 VSUBS 0.008887f
C576 B.n297 VSUBS 0.008887f
C577 B.n298 VSUBS 0.008887f
C578 B.n299 VSUBS 0.008887f
C579 B.n300 VSUBS 0.008887f
C580 B.n301 VSUBS 0.019548f
C581 B.n302 VSUBS 0.019548f
C582 B.n303 VSUBS 0.020445f
C583 B.n304 VSUBS 0.008887f
C584 B.n305 VSUBS 0.008887f
C585 B.n306 VSUBS 0.008887f
C586 B.n307 VSUBS 0.008887f
C587 B.n308 VSUBS 0.008887f
C588 B.n309 VSUBS 0.008887f
C589 B.n310 VSUBS 0.008887f
C590 B.n311 VSUBS 0.008887f
C591 B.n312 VSUBS 0.008887f
C592 B.n313 VSUBS 0.008887f
C593 B.n314 VSUBS 0.008887f
C594 B.n315 VSUBS 0.008887f
C595 B.n316 VSUBS 0.008887f
C596 B.n317 VSUBS 0.008887f
C597 B.n318 VSUBS 0.008887f
C598 B.n319 VSUBS 0.008887f
C599 B.n320 VSUBS 0.008887f
C600 B.n321 VSUBS 0.008887f
C601 B.n322 VSUBS 0.008887f
C602 B.n323 VSUBS 0.008887f
C603 B.n324 VSUBS 0.008887f
C604 B.n325 VSUBS 0.008887f
C605 B.n326 VSUBS 0.008887f
C606 B.n327 VSUBS 0.008887f
C607 B.n328 VSUBS 0.008887f
C608 B.n329 VSUBS 0.008887f
C609 B.n330 VSUBS 0.008887f
C610 B.n331 VSUBS 0.008887f
C611 B.n332 VSUBS 0.008887f
C612 B.n333 VSUBS 0.008887f
C613 B.n334 VSUBS 0.008887f
C614 B.n335 VSUBS 0.008887f
C615 B.n336 VSUBS 0.008887f
C616 B.n337 VSUBS 0.008887f
C617 B.n338 VSUBS 0.008887f
C618 B.n339 VSUBS 0.008887f
C619 B.n340 VSUBS 0.008887f
C620 B.n341 VSUBS 0.008887f
C621 B.n342 VSUBS 0.008887f
C622 B.n343 VSUBS 0.008887f
C623 B.n344 VSUBS 0.008887f
C624 B.n345 VSUBS 0.008887f
C625 B.n346 VSUBS 0.008887f
C626 B.n347 VSUBS 0.008887f
C627 B.n348 VSUBS 0.008887f
C628 B.n349 VSUBS 0.008887f
C629 B.n350 VSUBS 0.008887f
C630 B.n351 VSUBS 0.008887f
C631 B.n352 VSUBS 0.008887f
C632 B.n353 VSUBS 0.008887f
C633 B.n354 VSUBS 0.008887f
C634 B.n355 VSUBS 0.008887f
C635 B.n356 VSUBS 0.008887f
C636 B.n357 VSUBS 0.008887f
C637 B.n358 VSUBS 0.008887f
C638 B.n359 VSUBS 0.008887f
C639 B.n360 VSUBS 0.008887f
C640 B.n361 VSUBS 0.008887f
C641 B.n362 VSUBS 0.008887f
C642 B.n363 VSUBS 0.008887f
C643 B.n364 VSUBS 0.008887f
C644 B.n365 VSUBS 0.008887f
C645 B.n366 VSUBS 0.008887f
C646 B.n367 VSUBS 0.008887f
C647 B.n368 VSUBS 0.008887f
C648 B.n369 VSUBS 0.008887f
C649 B.n370 VSUBS 0.008887f
C650 B.n371 VSUBS 0.008887f
C651 B.n372 VSUBS 0.008887f
C652 B.n373 VSUBS 0.008887f
C653 B.n374 VSUBS 0.008887f
C654 B.n375 VSUBS 0.008887f
C655 B.n376 VSUBS 0.008887f
C656 B.n377 VSUBS 0.008887f
C657 B.n378 VSUBS 0.006143f
C658 B.n379 VSUBS 0.020591f
C659 B.n380 VSUBS 0.007188f
C660 B.n381 VSUBS 0.008887f
C661 B.n382 VSUBS 0.008887f
C662 B.n383 VSUBS 0.008887f
C663 B.n384 VSUBS 0.008887f
C664 B.n385 VSUBS 0.008887f
C665 B.n386 VSUBS 0.008887f
C666 B.n387 VSUBS 0.008887f
C667 B.n388 VSUBS 0.008887f
C668 B.n389 VSUBS 0.008887f
C669 B.n390 VSUBS 0.008887f
C670 B.n391 VSUBS 0.008887f
C671 B.n392 VSUBS 0.007188f
C672 B.n393 VSUBS 0.008887f
C673 B.n394 VSUBS 0.008887f
C674 B.n395 VSUBS 0.006143f
C675 B.n396 VSUBS 0.008887f
C676 B.n397 VSUBS 0.008887f
C677 B.n398 VSUBS 0.008887f
C678 B.n399 VSUBS 0.008887f
C679 B.n400 VSUBS 0.008887f
C680 B.n401 VSUBS 0.008887f
C681 B.n402 VSUBS 0.008887f
C682 B.n403 VSUBS 0.008887f
C683 B.n404 VSUBS 0.008887f
C684 B.n405 VSUBS 0.008887f
C685 B.n406 VSUBS 0.008887f
C686 B.n407 VSUBS 0.008887f
C687 B.n408 VSUBS 0.008887f
C688 B.n409 VSUBS 0.008887f
C689 B.n410 VSUBS 0.008887f
C690 B.n411 VSUBS 0.008887f
C691 B.n412 VSUBS 0.008887f
C692 B.n413 VSUBS 0.008887f
C693 B.n414 VSUBS 0.008887f
C694 B.n415 VSUBS 0.008887f
C695 B.n416 VSUBS 0.008887f
C696 B.n417 VSUBS 0.008887f
C697 B.n418 VSUBS 0.008887f
C698 B.n419 VSUBS 0.008887f
C699 B.n420 VSUBS 0.008887f
C700 B.n421 VSUBS 0.008887f
C701 B.n422 VSUBS 0.008887f
C702 B.n423 VSUBS 0.008887f
C703 B.n424 VSUBS 0.008887f
C704 B.n425 VSUBS 0.008887f
C705 B.n426 VSUBS 0.008887f
C706 B.n427 VSUBS 0.008887f
C707 B.n428 VSUBS 0.008887f
C708 B.n429 VSUBS 0.008887f
C709 B.n430 VSUBS 0.008887f
C710 B.n431 VSUBS 0.008887f
C711 B.n432 VSUBS 0.008887f
C712 B.n433 VSUBS 0.008887f
C713 B.n434 VSUBS 0.008887f
C714 B.n435 VSUBS 0.008887f
C715 B.n436 VSUBS 0.008887f
C716 B.n437 VSUBS 0.008887f
C717 B.n438 VSUBS 0.008887f
C718 B.n439 VSUBS 0.008887f
C719 B.n440 VSUBS 0.008887f
C720 B.n441 VSUBS 0.008887f
C721 B.n442 VSUBS 0.008887f
C722 B.n443 VSUBS 0.008887f
C723 B.n444 VSUBS 0.008887f
C724 B.n445 VSUBS 0.008887f
C725 B.n446 VSUBS 0.008887f
C726 B.n447 VSUBS 0.008887f
C727 B.n448 VSUBS 0.008887f
C728 B.n449 VSUBS 0.008887f
C729 B.n450 VSUBS 0.008887f
C730 B.n451 VSUBS 0.008887f
C731 B.n452 VSUBS 0.008887f
C732 B.n453 VSUBS 0.008887f
C733 B.n454 VSUBS 0.008887f
C734 B.n455 VSUBS 0.008887f
C735 B.n456 VSUBS 0.008887f
C736 B.n457 VSUBS 0.008887f
C737 B.n458 VSUBS 0.008887f
C738 B.n459 VSUBS 0.008887f
C739 B.n460 VSUBS 0.008887f
C740 B.n461 VSUBS 0.008887f
C741 B.n462 VSUBS 0.008887f
C742 B.n463 VSUBS 0.008887f
C743 B.n464 VSUBS 0.008887f
C744 B.n465 VSUBS 0.008887f
C745 B.n466 VSUBS 0.008887f
C746 B.n467 VSUBS 0.008887f
C747 B.n468 VSUBS 0.008887f
C748 B.n469 VSUBS 0.020445f
C749 B.n470 VSUBS 0.020445f
C750 B.n471 VSUBS 0.019548f
C751 B.n472 VSUBS 0.008887f
C752 B.n473 VSUBS 0.008887f
C753 B.n474 VSUBS 0.008887f
C754 B.n475 VSUBS 0.008887f
C755 B.n476 VSUBS 0.008887f
C756 B.n477 VSUBS 0.008887f
C757 B.n478 VSUBS 0.008887f
C758 B.n479 VSUBS 0.008887f
C759 B.n480 VSUBS 0.008887f
C760 B.n481 VSUBS 0.008887f
C761 B.n482 VSUBS 0.008887f
C762 B.n483 VSUBS 0.008887f
C763 B.n484 VSUBS 0.008887f
C764 B.n485 VSUBS 0.008887f
C765 B.n486 VSUBS 0.008887f
C766 B.n487 VSUBS 0.008887f
C767 B.n488 VSUBS 0.008887f
C768 B.n489 VSUBS 0.008887f
C769 B.n490 VSUBS 0.008887f
C770 B.n491 VSUBS 0.008887f
C771 B.n492 VSUBS 0.008887f
C772 B.n493 VSUBS 0.008887f
C773 B.n494 VSUBS 0.008887f
C774 B.n495 VSUBS 0.008887f
C775 B.n496 VSUBS 0.008887f
C776 B.n497 VSUBS 0.008887f
C777 B.n498 VSUBS 0.008887f
C778 B.n499 VSUBS 0.008887f
C779 B.n500 VSUBS 0.008887f
C780 B.n501 VSUBS 0.008887f
C781 B.n502 VSUBS 0.008887f
C782 B.n503 VSUBS 0.008887f
C783 B.n504 VSUBS 0.008887f
C784 B.n505 VSUBS 0.008887f
C785 B.n506 VSUBS 0.008887f
C786 B.n507 VSUBS 0.008887f
C787 B.n508 VSUBS 0.008887f
C788 B.n509 VSUBS 0.008887f
C789 B.n510 VSUBS 0.008887f
C790 B.n511 VSUBS 0.008887f
C791 B.n512 VSUBS 0.008887f
C792 B.n513 VSUBS 0.008887f
C793 B.n514 VSUBS 0.008887f
C794 B.n515 VSUBS 0.008887f
C795 B.n516 VSUBS 0.008887f
C796 B.n517 VSUBS 0.008887f
C797 B.n518 VSUBS 0.008887f
C798 B.n519 VSUBS 0.008887f
C799 B.n520 VSUBS 0.008887f
C800 B.n521 VSUBS 0.008887f
C801 B.n522 VSUBS 0.008887f
C802 B.n523 VSUBS 0.008887f
C803 B.n524 VSUBS 0.008887f
C804 B.n525 VSUBS 0.008887f
C805 B.n526 VSUBS 0.008887f
C806 B.n527 VSUBS 0.008887f
C807 B.n528 VSUBS 0.008887f
C808 B.n529 VSUBS 0.008887f
C809 B.n530 VSUBS 0.008887f
C810 B.n531 VSUBS 0.008887f
C811 B.n532 VSUBS 0.008887f
C812 B.n533 VSUBS 0.008887f
C813 B.n534 VSUBS 0.008887f
C814 B.n535 VSUBS 0.008887f
C815 B.n536 VSUBS 0.008887f
C816 B.n537 VSUBS 0.008887f
C817 B.n538 VSUBS 0.008887f
C818 B.n539 VSUBS 0.008887f
C819 B.n540 VSUBS 0.008887f
C820 B.n541 VSUBS 0.008887f
C821 B.n542 VSUBS 0.008887f
C822 B.n543 VSUBS 0.008887f
C823 B.n544 VSUBS 0.008887f
C824 B.n545 VSUBS 0.008887f
C825 B.n546 VSUBS 0.008887f
C826 B.n547 VSUBS 0.008887f
C827 B.n548 VSUBS 0.008887f
C828 B.n549 VSUBS 0.008887f
C829 B.n550 VSUBS 0.008887f
C830 B.n551 VSUBS 0.008887f
C831 B.n552 VSUBS 0.008887f
C832 B.n553 VSUBS 0.008887f
C833 B.n554 VSUBS 0.008887f
C834 B.n555 VSUBS 0.008887f
C835 B.n556 VSUBS 0.008887f
C836 B.n557 VSUBS 0.008887f
C837 B.n558 VSUBS 0.008887f
C838 B.n559 VSUBS 0.008887f
C839 B.n560 VSUBS 0.008887f
C840 B.n561 VSUBS 0.008887f
C841 B.n562 VSUBS 0.008887f
C842 B.n563 VSUBS 0.008887f
C843 B.n564 VSUBS 0.008887f
C844 B.n565 VSUBS 0.008887f
C845 B.n566 VSUBS 0.008887f
C846 B.n567 VSUBS 0.008887f
C847 B.n568 VSUBS 0.008887f
C848 B.n569 VSUBS 0.008887f
C849 B.n570 VSUBS 0.008887f
C850 B.n571 VSUBS 0.008887f
C851 B.n572 VSUBS 0.008887f
C852 B.n573 VSUBS 0.008887f
C853 B.n574 VSUBS 0.008887f
C854 B.n575 VSUBS 0.008887f
C855 B.n576 VSUBS 0.008887f
C856 B.n577 VSUBS 0.008887f
C857 B.n578 VSUBS 0.008887f
C858 B.n579 VSUBS 0.008887f
C859 B.n580 VSUBS 0.008887f
C860 B.n581 VSUBS 0.008887f
C861 B.n582 VSUBS 0.008887f
C862 B.n583 VSUBS 0.008887f
C863 B.n584 VSUBS 0.008887f
C864 B.n585 VSUBS 0.008887f
C865 B.n586 VSUBS 0.008887f
C866 B.n587 VSUBS 0.008887f
C867 B.n588 VSUBS 0.008887f
C868 B.n589 VSUBS 0.008887f
C869 B.n590 VSUBS 0.008887f
C870 B.n591 VSUBS 0.008887f
C871 B.n592 VSUBS 0.008887f
C872 B.n593 VSUBS 0.008887f
C873 B.n594 VSUBS 0.008887f
C874 B.n595 VSUBS 0.008887f
C875 B.n596 VSUBS 0.008887f
C876 B.n597 VSUBS 0.008887f
C877 B.n598 VSUBS 0.008887f
C878 B.n599 VSUBS 0.008887f
C879 B.n600 VSUBS 0.008887f
C880 B.n601 VSUBS 0.008887f
C881 B.n602 VSUBS 0.008887f
C882 B.n603 VSUBS 0.008887f
C883 B.n604 VSUBS 0.008887f
C884 B.n605 VSUBS 0.008887f
C885 B.n606 VSUBS 0.008887f
C886 B.n607 VSUBS 0.008887f
C887 B.n608 VSUBS 0.008887f
C888 B.n609 VSUBS 0.008887f
C889 B.n610 VSUBS 0.008887f
C890 B.n611 VSUBS 0.008887f
C891 B.n612 VSUBS 0.008887f
C892 B.n613 VSUBS 0.008887f
C893 B.n614 VSUBS 0.008887f
C894 B.n615 VSUBS 0.008887f
C895 B.n616 VSUBS 0.008887f
C896 B.n617 VSUBS 0.008887f
C897 B.n618 VSUBS 0.008887f
C898 B.n619 VSUBS 0.008887f
C899 B.n620 VSUBS 0.008887f
C900 B.n621 VSUBS 0.008887f
C901 B.n622 VSUBS 0.008887f
C902 B.n623 VSUBS 0.008887f
C903 B.n624 VSUBS 0.008887f
C904 B.n625 VSUBS 0.008887f
C905 B.n626 VSUBS 0.008887f
C906 B.n627 VSUBS 0.019548f
C907 B.n628 VSUBS 0.020445f
C908 B.n629 VSUBS 0.01933f
C909 B.n630 VSUBS 0.008887f
C910 B.n631 VSUBS 0.008887f
C911 B.n632 VSUBS 0.008887f
C912 B.n633 VSUBS 0.008887f
C913 B.n634 VSUBS 0.008887f
C914 B.n635 VSUBS 0.008887f
C915 B.n636 VSUBS 0.008887f
C916 B.n637 VSUBS 0.008887f
C917 B.n638 VSUBS 0.008887f
C918 B.n639 VSUBS 0.008887f
C919 B.n640 VSUBS 0.008887f
C920 B.n641 VSUBS 0.008887f
C921 B.n642 VSUBS 0.008887f
C922 B.n643 VSUBS 0.008887f
C923 B.n644 VSUBS 0.008887f
C924 B.n645 VSUBS 0.008887f
C925 B.n646 VSUBS 0.008887f
C926 B.n647 VSUBS 0.008887f
C927 B.n648 VSUBS 0.008887f
C928 B.n649 VSUBS 0.008887f
C929 B.n650 VSUBS 0.008887f
C930 B.n651 VSUBS 0.008887f
C931 B.n652 VSUBS 0.008887f
C932 B.n653 VSUBS 0.008887f
C933 B.n654 VSUBS 0.008887f
C934 B.n655 VSUBS 0.008887f
C935 B.n656 VSUBS 0.008887f
C936 B.n657 VSUBS 0.008887f
C937 B.n658 VSUBS 0.008887f
C938 B.n659 VSUBS 0.008887f
C939 B.n660 VSUBS 0.008887f
C940 B.n661 VSUBS 0.008887f
C941 B.n662 VSUBS 0.008887f
C942 B.n663 VSUBS 0.008887f
C943 B.n664 VSUBS 0.008887f
C944 B.n665 VSUBS 0.008887f
C945 B.n666 VSUBS 0.008887f
C946 B.n667 VSUBS 0.008887f
C947 B.n668 VSUBS 0.008887f
C948 B.n669 VSUBS 0.008887f
C949 B.n670 VSUBS 0.008887f
C950 B.n671 VSUBS 0.008887f
C951 B.n672 VSUBS 0.008887f
C952 B.n673 VSUBS 0.008887f
C953 B.n674 VSUBS 0.008887f
C954 B.n675 VSUBS 0.008887f
C955 B.n676 VSUBS 0.008887f
C956 B.n677 VSUBS 0.008887f
C957 B.n678 VSUBS 0.008887f
C958 B.n679 VSUBS 0.008887f
C959 B.n680 VSUBS 0.008887f
C960 B.n681 VSUBS 0.008887f
C961 B.n682 VSUBS 0.008887f
C962 B.n683 VSUBS 0.008887f
C963 B.n684 VSUBS 0.008887f
C964 B.n685 VSUBS 0.008887f
C965 B.n686 VSUBS 0.008887f
C966 B.n687 VSUBS 0.008887f
C967 B.n688 VSUBS 0.008887f
C968 B.n689 VSUBS 0.008887f
C969 B.n690 VSUBS 0.008887f
C970 B.n691 VSUBS 0.008887f
C971 B.n692 VSUBS 0.008887f
C972 B.n693 VSUBS 0.008887f
C973 B.n694 VSUBS 0.008887f
C974 B.n695 VSUBS 0.008887f
C975 B.n696 VSUBS 0.008887f
C976 B.n697 VSUBS 0.008887f
C977 B.n698 VSUBS 0.008887f
C978 B.n699 VSUBS 0.008887f
C979 B.n700 VSUBS 0.008887f
C980 B.n701 VSUBS 0.008887f
C981 B.n702 VSUBS 0.008887f
C982 B.n703 VSUBS 0.006143f
C983 B.n704 VSUBS 0.008887f
C984 B.n705 VSUBS 0.008887f
C985 B.n706 VSUBS 0.007188f
C986 B.n707 VSUBS 0.008887f
C987 B.n708 VSUBS 0.008887f
C988 B.n709 VSUBS 0.008887f
C989 B.n710 VSUBS 0.008887f
C990 B.n711 VSUBS 0.008887f
C991 B.n712 VSUBS 0.008887f
C992 B.n713 VSUBS 0.008887f
C993 B.n714 VSUBS 0.008887f
C994 B.n715 VSUBS 0.008887f
C995 B.n716 VSUBS 0.008887f
C996 B.n717 VSUBS 0.008887f
C997 B.n718 VSUBS 0.007188f
C998 B.n719 VSUBS 0.020591f
C999 B.n720 VSUBS 0.006143f
C1000 B.n721 VSUBS 0.008887f
C1001 B.n722 VSUBS 0.008887f
C1002 B.n723 VSUBS 0.008887f
C1003 B.n724 VSUBS 0.008887f
C1004 B.n725 VSUBS 0.008887f
C1005 B.n726 VSUBS 0.008887f
C1006 B.n727 VSUBS 0.008887f
C1007 B.n728 VSUBS 0.008887f
C1008 B.n729 VSUBS 0.008887f
C1009 B.n730 VSUBS 0.008887f
C1010 B.n731 VSUBS 0.008887f
C1011 B.n732 VSUBS 0.008887f
C1012 B.n733 VSUBS 0.008887f
C1013 B.n734 VSUBS 0.008887f
C1014 B.n735 VSUBS 0.008887f
C1015 B.n736 VSUBS 0.008887f
C1016 B.n737 VSUBS 0.008887f
C1017 B.n738 VSUBS 0.008887f
C1018 B.n739 VSUBS 0.008887f
C1019 B.n740 VSUBS 0.008887f
C1020 B.n741 VSUBS 0.008887f
C1021 B.n742 VSUBS 0.008887f
C1022 B.n743 VSUBS 0.008887f
C1023 B.n744 VSUBS 0.008887f
C1024 B.n745 VSUBS 0.008887f
C1025 B.n746 VSUBS 0.008887f
C1026 B.n747 VSUBS 0.008887f
C1027 B.n748 VSUBS 0.008887f
C1028 B.n749 VSUBS 0.008887f
C1029 B.n750 VSUBS 0.008887f
C1030 B.n751 VSUBS 0.008887f
C1031 B.n752 VSUBS 0.008887f
C1032 B.n753 VSUBS 0.008887f
C1033 B.n754 VSUBS 0.008887f
C1034 B.n755 VSUBS 0.008887f
C1035 B.n756 VSUBS 0.008887f
C1036 B.n757 VSUBS 0.008887f
C1037 B.n758 VSUBS 0.008887f
C1038 B.n759 VSUBS 0.008887f
C1039 B.n760 VSUBS 0.008887f
C1040 B.n761 VSUBS 0.008887f
C1041 B.n762 VSUBS 0.008887f
C1042 B.n763 VSUBS 0.008887f
C1043 B.n764 VSUBS 0.008887f
C1044 B.n765 VSUBS 0.008887f
C1045 B.n766 VSUBS 0.008887f
C1046 B.n767 VSUBS 0.008887f
C1047 B.n768 VSUBS 0.008887f
C1048 B.n769 VSUBS 0.008887f
C1049 B.n770 VSUBS 0.008887f
C1050 B.n771 VSUBS 0.008887f
C1051 B.n772 VSUBS 0.008887f
C1052 B.n773 VSUBS 0.008887f
C1053 B.n774 VSUBS 0.008887f
C1054 B.n775 VSUBS 0.008887f
C1055 B.n776 VSUBS 0.008887f
C1056 B.n777 VSUBS 0.008887f
C1057 B.n778 VSUBS 0.008887f
C1058 B.n779 VSUBS 0.008887f
C1059 B.n780 VSUBS 0.008887f
C1060 B.n781 VSUBS 0.008887f
C1061 B.n782 VSUBS 0.008887f
C1062 B.n783 VSUBS 0.008887f
C1063 B.n784 VSUBS 0.008887f
C1064 B.n785 VSUBS 0.008887f
C1065 B.n786 VSUBS 0.008887f
C1066 B.n787 VSUBS 0.008887f
C1067 B.n788 VSUBS 0.008887f
C1068 B.n789 VSUBS 0.008887f
C1069 B.n790 VSUBS 0.008887f
C1070 B.n791 VSUBS 0.008887f
C1071 B.n792 VSUBS 0.008887f
C1072 B.n793 VSUBS 0.008887f
C1073 B.n794 VSUBS 0.008887f
C1074 B.n795 VSUBS 0.020445f
C1075 B.n796 VSUBS 0.019548f
C1076 B.n797 VSUBS 0.019548f
C1077 B.n798 VSUBS 0.008887f
C1078 B.n799 VSUBS 0.008887f
C1079 B.n800 VSUBS 0.008887f
C1080 B.n801 VSUBS 0.008887f
C1081 B.n802 VSUBS 0.008887f
C1082 B.n803 VSUBS 0.008887f
C1083 B.n804 VSUBS 0.008887f
C1084 B.n805 VSUBS 0.008887f
C1085 B.n806 VSUBS 0.008887f
C1086 B.n807 VSUBS 0.008887f
C1087 B.n808 VSUBS 0.008887f
C1088 B.n809 VSUBS 0.008887f
C1089 B.n810 VSUBS 0.008887f
C1090 B.n811 VSUBS 0.008887f
C1091 B.n812 VSUBS 0.008887f
C1092 B.n813 VSUBS 0.008887f
C1093 B.n814 VSUBS 0.008887f
C1094 B.n815 VSUBS 0.008887f
C1095 B.n816 VSUBS 0.008887f
C1096 B.n817 VSUBS 0.008887f
C1097 B.n818 VSUBS 0.008887f
C1098 B.n819 VSUBS 0.008887f
C1099 B.n820 VSUBS 0.008887f
C1100 B.n821 VSUBS 0.008887f
C1101 B.n822 VSUBS 0.008887f
C1102 B.n823 VSUBS 0.008887f
C1103 B.n824 VSUBS 0.008887f
C1104 B.n825 VSUBS 0.008887f
C1105 B.n826 VSUBS 0.008887f
C1106 B.n827 VSUBS 0.008887f
C1107 B.n828 VSUBS 0.008887f
C1108 B.n829 VSUBS 0.008887f
C1109 B.n830 VSUBS 0.008887f
C1110 B.n831 VSUBS 0.008887f
C1111 B.n832 VSUBS 0.008887f
C1112 B.n833 VSUBS 0.008887f
C1113 B.n834 VSUBS 0.008887f
C1114 B.n835 VSUBS 0.008887f
C1115 B.n836 VSUBS 0.008887f
C1116 B.n837 VSUBS 0.008887f
C1117 B.n838 VSUBS 0.008887f
C1118 B.n839 VSUBS 0.008887f
C1119 B.n840 VSUBS 0.008887f
C1120 B.n841 VSUBS 0.008887f
C1121 B.n842 VSUBS 0.008887f
C1122 B.n843 VSUBS 0.008887f
C1123 B.n844 VSUBS 0.008887f
C1124 B.n845 VSUBS 0.008887f
C1125 B.n846 VSUBS 0.008887f
C1126 B.n847 VSUBS 0.008887f
C1127 B.n848 VSUBS 0.008887f
C1128 B.n849 VSUBS 0.008887f
C1129 B.n850 VSUBS 0.008887f
C1130 B.n851 VSUBS 0.008887f
C1131 B.n852 VSUBS 0.008887f
C1132 B.n853 VSUBS 0.008887f
C1133 B.n854 VSUBS 0.008887f
C1134 B.n855 VSUBS 0.008887f
C1135 B.n856 VSUBS 0.008887f
C1136 B.n857 VSUBS 0.008887f
C1137 B.n858 VSUBS 0.008887f
C1138 B.n859 VSUBS 0.008887f
C1139 B.n860 VSUBS 0.008887f
C1140 B.n861 VSUBS 0.008887f
C1141 B.n862 VSUBS 0.008887f
C1142 B.n863 VSUBS 0.008887f
C1143 B.n864 VSUBS 0.008887f
C1144 B.n865 VSUBS 0.008887f
C1145 B.n866 VSUBS 0.008887f
C1146 B.n867 VSUBS 0.008887f
C1147 B.n868 VSUBS 0.008887f
C1148 B.n869 VSUBS 0.008887f
C1149 B.n870 VSUBS 0.008887f
C1150 B.n871 VSUBS 0.008887f
C1151 B.n872 VSUBS 0.008887f
C1152 B.n873 VSUBS 0.008887f
C1153 B.n874 VSUBS 0.008887f
C1154 B.n875 VSUBS 0.020124f
.ends

