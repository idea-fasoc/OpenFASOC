* NGSPICE file created from diff_pair_sample_1359.ext - technology: sky130A

.subckt diff_pair_sample_1359 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=0 ps=0 w=13.59 l=1.32
X1 VTAIL.t19 VN.t0 VDD2.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X2 VDD2.t6 VN.t1 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X3 VTAIL.t17 VN.t2 VDD2.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X4 VDD2.t3 VN.t3 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=2.24235 ps=13.92 w=13.59 l=1.32
X5 VTAIL.t9 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X6 VDD2.t0 VN.t4 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=2.24235 ps=13.92 w=13.59 l=1.32
X7 VDD1.t8 VP.t1 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=2.24235 ps=13.92 w=13.59 l=1.32
X8 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=0 ps=0 w=13.59 l=1.32
X9 VDD1.t7 VP.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=5.3001 ps=27.96 w=13.59 l=1.32
X10 VTAIL.t0 VP.t3 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X11 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=0 ps=0 w=13.59 l=1.32
X12 VDD2.t5 VN.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X13 VDD2.t4 VN.t6 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=5.3001 ps=27.96 w=13.59 l=1.32
X14 VTAIL.t6 VP.t4 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X15 VDD1.t4 VP.t5 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=2.24235 ps=13.92 w=13.59 l=1.32
X16 VDD2.t1 VN.t7 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=5.3001 ps=27.96 w=13.59 l=1.32
X17 VTAIL.t3 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3001 pd=27.96 as=0 ps=0 w=13.59 l=1.32
X19 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X20 VDD1.t1 VP.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=5.3001 ps=27.96 w=13.59 l=1.32
X21 VDD1.t0 VP.t9 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X22 VTAIL.t11 VN.t8 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
X23 VTAIL.t10 VN.t9 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.24235 pd=13.92 as=2.24235 ps=13.92 w=13.59 l=1.32
R0 B.n819 B.n818 585
R1 B.n327 B.n120 585
R2 B.n326 B.n325 585
R3 B.n324 B.n323 585
R4 B.n322 B.n321 585
R5 B.n320 B.n319 585
R6 B.n318 B.n317 585
R7 B.n316 B.n315 585
R8 B.n314 B.n313 585
R9 B.n312 B.n311 585
R10 B.n310 B.n309 585
R11 B.n308 B.n307 585
R12 B.n306 B.n305 585
R13 B.n304 B.n303 585
R14 B.n302 B.n301 585
R15 B.n300 B.n299 585
R16 B.n298 B.n297 585
R17 B.n296 B.n295 585
R18 B.n294 B.n293 585
R19 B.n292 B.n291 585
R20 B.n290 B.n289 585
R21 B.n288 B.n287 585
R22 B.n286 B.n285 585
R23 B.n284 B.n283 585
R24 B.n282 B.n281 585
R25 B.n280 B.n279 585
R26 B.n278 B.n277 585
R27 B.n276 B.n275 585
R28 B.n274 B.n273 585
R29 B.n272 B.n271 585
R30 B.n270 B.n269 585
R31 B.n268 B.n267 585
R32 B.n266 B.n265 585
R33 B.n264 B.n263 585
R34 B.n262 B.n261 585
R35 B.n260 B.n259 585
R36 B.n258 B.n257 585
R37 B.n256 B.n255 585
R38 B.n254 B.n253 585
R39 B.n252 B.n251 585
R40 B.n250 B.n249 585
R41 B.n248 B.n247 585
R42 B.n246 B.n245 585
R43 B.n244 B.n243 585
R44 B.n242 B.n241 585
R45 B.n240 B.n239 585
R46 B.n238 B.n237 585
R47 B.n236 B.n235 585
R48 B.n234 B.n233 585
R49 B.n232 B.n231 585
R50 B.n230 B.n229 585
R51 B.n228 B.n227 585
R52 B.n226 B.n225 585
R53 B.n224 B.n223 585
R54 B.n222 B.n221 585
R55 B.n220 B.n219 585
R56 B.n218 B.n217 585
R57 B.n216 B.n215 585
R58 B.n214 B.n213 585
R59 B.n212 B.n211 585
R60 B.n210 B.n209 585
R61 B.n208 B.n207 585
R62 B.n206 B.n205 585
R63 B.n204 B.n203 585
R64 B.n202 B.n201 585
R65 B.n200 B.n199 585
R66 B.n198 B.n197 585
R67 B.n196 B.n195 585
R68 B.n194 B.n193 585
R69 B.n192 B.n191 585
R70 B.n190 B.n189 585
R71 B.n188 B.n187 585
R72 B.n186 B.n185 585
R73 B.n184 B.n183 585
R74 B.n182 B.n181 585
R75 B.n180 B.n179 585
R76 B.n178 B.n177 585
R77 B.n176 B.n175 585
R78 B.n174 B.n173 585
R79 B.n172 B.n171 585
R80 B.n170 B.n169 585
R81 B.n168 B.n167 585
R82 B.n166 B.n165 585
R83 B.n164 B.n163 585
R84 B.n162 B.n161 585
R85 B.n160 B.n159 585
R86 B.n158 B.n157 585
R87 B.n156 B.n155 585
R88 B.n154 B.n153 585
R89 B.n152 B.n151 585
R90 B.n150 B.n149 585
R91 B.n148 B.n147 585
R92 B.n146 B.n145 585
R93 B.n144 B.n143 585
R94 B.n142 B.n141 585
R95 B.n140 B.n139 585
R96 B.n138 B.n137 585
R97 B.n136 B.n135 585
R98 B.n134 B.n133 585
R99 B.n132 B.n131 585
R100 B.n130 B.n129 585
R101 B.n128 B.n127 585
R102 B.n817 B.n69 585
R103 B.n822 B.n69 585
R104 B.n816 B.n68 585
R105 B.n823 B.n68 585
R106 B.n815 B.n814 585
R107 B.n814 B.n64 585
R108 B.n813 B.n63 585
R109 B.n829 B.n63 585
R110 B.n812 B.n62 585
R111 B.n830 B.n62 585
R112 B.n811 B.n61 585
R113 B.n831 B.n61 585
R114 B.n810 B.n809 585
R115 B.n809 B.n57 585
R116 B.n808 B.n56 585
R117 B.n837 B.n56 585
R118 B.n807 B.n55 585
R119 B.n838 B.n55 585
R120 B.n806 B.n54 585
R121 B.n839 B.n54 585
R122 B.n805 B.n804 585
R123 B.n804 B.n50 585
R124 B.n803 B.n49 585
R125 B.n845 B.n49 585
R126 B.n802 B.n48 585
R127 B.n846 B.n48 585
R128 B.n801 B.n47 585
R129 B.n847 B.n47 585
R130 B.n800 B.n799 585
R131 B.n799 B.n43 585
R132 B.n798 B.n42 585
R133 B.n853 B.n42 585
R134 B.n797 B.n41 585
R135 B.n854 B.n41 585
R136 B.n796 B.n40 585
R137 B.n855 B.n40 585
R138 B.n795 B.n794 585
R139 B.n794 B.n39 585
R140 B.n793 B.n35 585
R141 B.n861 B.n35 585
R142 B.n792 B.n34 585
R143 B.n862 B.n34 585
R144 B.n791 B.n33 585
R145 B.n863 B.n33 585
R146 B.n790 B.n789 585
R147 B.n789 B.n29 585
R148 B.n788 B.n28 585
R149 B.n869 B.n28 585
R150 B.n787 B.n27 585
R151 B.n870 B.n27 585
R152 B.n786 B.n26 585
R153 B.n871 B.n26 585
R154 B.n785 B.n784 585
R155 B.n784 B.n22 585
R156 B.n783 B.n21 585
R157 B.n877 B.n21 585
R158 B.n782 B.n20 585
R159 B.n878 B.n20 585
R160 B.n781 B.n19 585
R161 B.n879 B.n19 585
R162 B.n780 B.n779 585
R163 B.n779 B.n15 585
R164 B.n778 B.n14 585
R165 B.n885 B.n14 585
R166 B.n777 B.n13 585
R167 B.n886 B.n13 585
R168 B.n776 B.n12 585
R169 B.n887 B.n12 585
R170 B.n775 B.n774 585
R171 B.n774 B.n8 585
R172 B.n773 B.n7 585
R173 B.n893 B.n7 585
R174 B.n772 B.n6 585
R175 B.n894 B.n6 585
R176 B.n771 B.n5 585
R177 B.n895 B.n5 585
R178 B.n770 B.n769 585
R179 B.n769 B.n4 585
R180 B.n768 B.n328 585
R181 B.n768 B.n767 585
R182 B.n758 B.n329 585
R183 B.n330 B.n329 585
R184 B.n760 B.n759 585
R185 B.n761 B.n760 585
R186 B.n757 B.n334 585
R187 B.n338 B.n334 585
R188 B.n756 B.n755 585
R189 B.n755 B.n754 585
R190 B.n336 B.n335 585
R191 B.n337 B.n336 585
R192 B.n747 B.n746 585
R193 B.n748 B.n747 585
R194 B.n745 B.n342 585
R195 B.n346 B.n342 585
R196 B.n744 B.n743 585
R197 B.n743 B.n742 585
R198 B.n344 B.n343 585
R199 B.n345 B.n344 585
R200 B.n735 B.n734 585
R201 B.n736 B.n735 585
R202 B.n733 B.n351 585
R203 B.n351 B.n350 585
R204 B.n732 B.n731 585
R205 B.n731 B.n730 585
R206 B.n353 B.n352 585
R207 B.n354 B.n353 585
R208 B.n723 B.n722 585
R209 B.n724 B.n723 585
R210 B.n721 B.n359 585
R211 B.n359 B.n358 585
R212 B.n720 B.n719 585
R213 B.n719 B.n718 585
R214 B.n361 B.n360 585
R215 B.n711 B.n361 585
R216 B.n710 B.n709 585
R217 B.n712 B.n710 585
R218 B.n708 B.n366 585
R219 B.n366 B.n365 585
R220 B.n707 B.n706 585
R221 B.n706 B.n705 585
R222 B.n368 B.n367 585
R223 B.n369 B.n368 585
R224 B.n698 B.n697 585
R225 B.n699 B.n698 585
R226 B.n696 B.n374 585
R227 B.n374 B.n373 585
R228 B.n695 B.n694 585
R229 B.n694 B.n693 585
R230 B.n376 B.n375 585
R231 B.n377 B.n376 585
R232 B.n686 B.n685 585
R233 B.n687 B.n686 585
R234 B.n684 B.n382 585
R235 B.n382 B.n381 585
R236 B.n683 B.n682 585
R237 B.n682 B.n681 585
R238 B.n384 B.n383 585
R239 B.n385 B.n384 585
R240 B.n674 B.n673 585
R241 B.n675 B.n674 585
R242 B.n672 B.n390 585
R243 B.n390 B.n389 585
R244 B.n671 B.n670 585
R245 B.n670 B.n669 585
R246 B.n392 B.n391 585
R247 B.n393 B.n392 585
R248 B.n662 B.n661 585
R249 B.n663 B.n662 585
R250 B.n660 B.n398 585
R251 B.n398 B.n397 585
R252 B.n655 B.n654 585
R253 B.n653 B.n451 585
R254 B.n652 B.n450 585
R255 B.n657 B.n450 585
R256 B.n651 B.n650 585
R257 B.n649 B.n648 585
R258 B.n647 B.n646 585
R259 B.n645 B.n644 585
R260 B.n643 B.n642 585
R261 B.n641 B.n640 585
R262 B.n639 B.n638 585
R263 B.n637 B.n636 585
R264 B.n635 B.n634 585
R265 B.n633 B.n632 585
R266 B.n631 B.n630 585
R267 B.n629 B.n628 585
R268 B.n627 B.n626 585
R269 B.n625 B.n624 585
R270 B.n623 B.n622 585
R271 B.n621 B.n620 585
R272 B.n619 B.n618 585
R273 B.n617 B.n616 585
R274 B.n615 B.n614 585
R275 B.n613 B.n612 585
R276 B.n611 B.n610 585
R277 B.n609 B.n608 585
R278 B.n607 B.n606 585
R279 B.n605 B.n604 585
R280 B.n603 B.n602 585
R281 B.n601 B.n600 585
R282 B.n599 B.n598 585
R283 B.n597 B.n596 585
R284 B.n595 B.n594 585
R285 B.n593 B.n592 585
R286 B.n591 B.n590 585
R287 B.n589 B.n588 585
R288 B.n587 B.n586 585
R289 B.n585 B.n584 585
R290 B.n583 B.n582 585
R291 B.n581 B.n580 585
R292 B.n579 B.n578 585
R293 B.n577 B.n576 585
R294 B.n575 B.n574 585
R295 B.n573 B.n572 585
R296 B.n571 B.n570 585
R297 B.n569 B.n568 585
R298 B.n567 B.n566 585
R299 B.n564 B.n563 585
R300 B.n562 B.n561 585
R301 B.n560 B.n559 585
R302 B.n558 B.n557 585
R303 B.n556 B.n555 585
R304 B.n554 B.n553 585
R305 B.n552 B.n551 585
R306 B.n550 B.n549 585
R307 B.n548 B.n547 585
R308 B.n546 B.n545 585
R309 B.n543 B.n542 585
R310 B.n541 B.n540 585
R311 B.n539 B.n538 585
R312 B.n537 B.n536 585
R313 B.n535 B.n534 585
R314 B.n533 B.n532 585
R315 B.n531 B.n530 585
R316 B.n529 B.n528 585
R317 B.n527 B.n526 585
R318 B.n525 B.n524 585
R319 B.n523 B.n522 585
R320 B.n521 B.n520 585
R321 B.n519 B.n518 585
R322 B.n517 B.n516 585
R323 B.n515 B.n514 585
R324 B.n513 B.n512 585
R325 B.n511 B.n510 585
R326 B.n509 B.n508 585
R327 B.n507 B.n506 585
R328 B.n505 B.n504 585
R329 B.n503 B.n502 585
R330 B.n501 B.n500 585
R331 B.n499 B.n498 585
R332 B.n497 B.n496 585
R333 B.n495 B.n494 585
R334 B.n493 B.n492 585
R335 B.n491 B.n490 585
R336 B.n489 B.n488 585
R337 B.n487 B.n486 585
R338 B.n485 B.n484 585
R339 B.n483 B.n482 585
R340 B.n481 B.n480 585
R341 B.n479 B.n478 585
R342 B.n477 B.n476 585
R343 B.n475 B.n474 585
R344 B.n473 B.n472 585
R345 B.n471 B.n470 585
R346 B.n469 B.n468 585
R347 B.n467 B.n466 585
R348 B.n465 B.n464 585
R349 B.n463 B.n462 585
R350 B.n461 B.n460 585
R351 B.n459 B.n458 585
R352 B.n457 B.n456 585
R353 B.n400 B.n399 585
R354 B.n659 B.n658 585
R355 B.n658 B.n657 585
R356 B.n396 B.n395 585
R357 B.n397 B.n396 585
R358 B.n665 B.n664 585
R359 B.n664 B.n663 585
R360 B.n666 B.n394 585
R361 B.n394 B.n393 585
R362 B.n668 B.n667 585
R363 B.n669 B.n668 585
R364 B.n388 B.n387 585
R365 B.n389 B.n388 585
R366 B.n677 B.n676 585
R367 B.n676 B.n675 585
R368 B.n678 B.n386 585
R369 B.n386 B.n385 585
R370 B.n680 B.n679 585
R371 B.n681 B.n680 585
R372 B.n380 B.n379 585
R373 B.n381 B.n380 585
R374 B.n689 B.n688 585
R375 B.n688 B.n687 585
R376 B.n690 B.n378 585
R377 B.n378 B.n377 585
R378 B.n692 B.n691 585
R379 B.n693 B.n692 585
R380 B.n372 B.n371 585
R381 B.n373 B.n372 585
R382 B.n701 B.n700 585
R383 B.n700 B.n699 585
R384 B.n702 B.n370 585
R385 B.n370 B.n369 585
R386 B.n704 B.n703 585
R387 B.n705 B.n704 585
R388 B.n364 B.n363 585
R389 B.n365 B.n364 585
R390 B.n714 B.n713 585
R391 B.n713 B.n712 585
R392 B.n715 B.n362 585
R393 B.n711 B.n362 585
R394 B.n717 B.n716 585
R395 B.n718 B.n717 585
R396 B.n357 B.n356 585
R397 B.n358 B.n357 585
R398 B.n726 B.n725 585
R399 B.n725 B.n724 585
R400 B.n727 B.n355 585
R401 B.n355 B.n354 585
R402 B.n729 B.n728 585
R403 B.n730 B.n729 585
R404 B.n349 B.n348 585
R405 B.n350 B.n349 585
R406 B.n738 B.n737 585
R407 B.n737 B.n736 585
R408 B.n739 B.n347 585
R409 B.n347 B.n345 585
R410 B.n741 B.n740 585
R411 B.n742 B.n741 585
R412 B.n341 B.n340 585
R413 B.n346 B.n341 585
R414 B.n750 B.n749 585
R415 B.n749 B.n748 585
R416 B.n751 B.n339 585
R417 B.n339 B.n337 585
R418 B.n753 B.n752 585
R419 B.n754 B.n753 585
R420 B.n333 B.n332 585
R421 B.n338 B.n333 585
R422 B.n763 B.n762 585
R423 B.n762 B.n761 585
R424 B.n764 B.n331 585
R425 B.n331 B.n330 585
R426 B.n766 B.n765 585
R427 B.n767 B.n766 585
R428 B.n2 B.n0 585
R429 B.n4 B.n2 585
R430 B.n3 B.n1 585
R431 B.n894 B.n3 585
R432 B.n892 B.n891 585
R433 B.n893 B.n892 585
R434 B.n890 B.n9 585
R435 B.n9 B.n8 585
R436 B.n889 B.n888 585
R437 B.n888 B.n887 585
R438 B.n11 B.n10 585
R439 B.n886 B.n11 585
R440 B.n884 B.n883 585
R441 B.n885 B.n884 585
R442 B.n882 B.n16 585
R443 B.n16 B.n15 585
R444 B.n881 B.n880 585
R445 B.n880 B.n879 585
R446 B.n18 B.n17 585
R447 B.n878 B.n18 585
R448 B.n876 B.n875 585
R449 B.n877 B.n876 585
R450 B.n874 B.n23 585
R451 B.n23 B.n22 585
R452 B.n873 B.n872 585
R453 B.n872 B.n871 585
R454 B.n25 B.n24 585
R455 B.n870 B.n25 585
R456 B.n868 B.n867 585
R457 B.n869 B.n868 585
R458 B.n866 B.n30 585
R459 B.n30 B.n29 585
R460 B.n865 B.n864 585
R461 B.n864 B.n863 585
R462 B.n32 B.n31 585
R463 B.n862 B.n32 585
R464 B.n860 B.n859 585
R465 B.n861 B.n860 585
R466 B.n858 B.n36 585
R467 B.n39 B.n36 585
R468 B.n857 B.n856 585
R469 B.n856 B.n855 585
R470 B.n38 B.n37 585
R471 B.n854 B.n38 585
R472 B.n852 B.n851 585
R473 B.n853 B.n852 585
R474 B.n850 B.n44 585
R475 B.n44 B.n43 585
R476 B.n849 B.n848 585
R477 B.n848 B.n847 585
R478 B.n46 B.n45 585
R479 B.n846 B.n46 585
R480 B.n844 B.n843 585
R481 B.n845 B.n844 585
R482 B.n842 B.n51 585
R483 B.n51 B.n50 585
R484 B.n841 B.n840 585
R485 B.n840 B.n839 585
R486 B.n53 B.n52 585
R487 B.n838 B.n53 585
R488 B.n836 B.n835 585
R489 B.n837 B.n836 585
R490 B.n834 B.n58 585
R491 B.n58 B.n57 585
R492 B.n833 B.n832 585
R493 B.n832 B.n831 585
R494 B.n60 B.n59 585
R495 B.n830 B.n60 585
R496 B.n828 B.n827 585
R497 B.n829 B.n828 585
R498 B.n826 B.n65 585
R499 B.n65 B.n64 585
R500 B.n825 B.n824 585
R501 B.n824 B.n823 585
R502 B.n67 B.n66 585
R503 B.n822 B.n67 585
R504 B.n897 B.n896 585
R505 B.n896 B.n895 585
R506 B.n655 B.n396 550.159
R507 B.n127 B.n67 550.159
R508 B.n658 B.n398 550.159
R509 B.n819 B.n69 550.159
R510 B.n454 B.t10 452.82
R511 B.n452 B.t21 452.82
R512 B.n124 B.t14 452.82
R513 B.n121 B.t18 452.82
R514 B.n454 B.t13 341.894
R515 B.n452 B.t23 341.894
R516 B.n124 B.t16 341.894
R517 B.n121 B.t19 341.894
R518 B.n455 B.t12 309.894
R519 B.n122 B.t20 309.894
R520 B.n453 B.t22 309.894
R521 B.n125 B.t17 309.894
R522 B.n821 B.n820 256.663
R523 B.n821 B.n119 256.663
R524 B.n821 B.n118 256.663
R525 B.n821 B.n117 256.663
R526 B.n821 B.n116 256.663
R527 B.n821 B.n115 256.663
R528 B.n821 B.n114 256.663
R529 B.n821 B.n113 256.663
R530 B.n821 B.n112 256.663
R531 B.n821 B.n111 256.663
R532 B.n821 B.n110 256.663
R533 B.n821 B.n109 256.663
R534 B.n821 B.n108 256.663
R535 B.n821 B.n107 256.663
R536 B.n821 B.n106 256.663
R537 B.n821 B.n105 256.663
R538 B.n821 B.n104 256.663
R539 B.n821 B.n103 256.663
R540 B.n821 B.n102 256.663
R541 B.n821 B.n101 256.663
R542 B.n821 B.n100 256.663
R543 B.n821 B.n99 256.663
R544 B.n821 B.n98 256.663
R545 B.n821 B.n97 256.663
R546 B.n821 B.n96 256.663
R547 B.n821 B.n95 256.663
R548 B.n821 B.n94 256.663
R549 B.n821 B.n93 256.663
R550 B.n821 B.n92 256.663
R551 B.n821 B.n91 256.663
R552 B.n821 B.n90 256.663
R553 B.n821 B.n89 256.663
R554 B.n821 B.n88 256.663
R555 B.n821 B.n87 256.663
R556 B.n821 B.n86 256.663
R557 B.n821 B.n85 256.663
R558 B.n821 B.n84 256.663
R559 B.n821 B.n83 256.663
R560 B.n821 B.n82 256.663
R561 B.n821 B.n81 256.663
R562 B.n821 B.n80 256.663
R563 B.n821 B.n79 256.663
R564 B.n821 B.n78 256.663
R565 B.n821 B.n77 256.663
R566 B.n821 B.n76 256.663
R567 B.n821 B.n75 256.663
R568 B.n821 B.n74 256.663
R569 B.n821 B.n73 256.663
R570 B.n821 B.n72 256.663
R571 B.n821 B.n71 256.663
R572 B.n821 B.n70 256.663
R573 B.n657 B.n656 256.663
R574 B.n657 B.n401 256.663
R575 B.n657 B.n402 256.663
R576 B.n657 B.n403 256.663
R577 B.n657 B.n404 256.663
R578 B.n657 B.n405 256.663
R579 B.n657 B.n406 256.663
R580 B.n657 B.n407 256.663
R581 B.n657 B.n408 256.663
R582 B.n657 B.n409 256.663
R583 B.n657 B.n410 256.663
R584 B.n657 B.n411 256.663
R585 B.n657 B.n412 256.663
R586 B.n657 B.n413 256.663
R587 B.n657 B.n414 256.663
R588 B.n657 B.n415 256.663
R589 B.n657 B.n416 256.663
R590 B.n657 B.n417 256.663
R591 B.n657 B.n418 256.663
R592 B.n657 B.n419 256.663
R593 B.n657 B.n420 256.663
R594 B.n657 B.n421 256.663
R595 B.n657 B.n422 256.663
R596 B.n657 B.n423 256.663
R597 B.n657 B.n424 256.663
R598 B.n657 B.n425 256.663
R599 B.n657 B.n426 256.663
R600 B.n657 B.n427 256.663
R601 B.n657 B.n428 256.663
R602 B.n657 B.n429 256.663
R603 B.n657 B.n430 256.663
R604 B.n657 B.n431 256.663
R605 B.n657 B.n432 256.663
R606 B.n657 B.n433 256.663
R607 B.n657 B.n434 256.663
R608 B.n657 B.n435 256.663
R609 B.n657 B.n436 256.663
R610 B.n657 B.n437 256.663
R611 B.n657 B.n438 256.663
R612 B.n657 B.n439 256.663
R613 B.n657 B.n440 256.663
R614 B.n657 B.n441 256.663
R615 B.n657 B.n442 256.663
R616 B.n657 B.n443 256.663
R617 B.n657 B.n444 256.663
R618 B.n657 B.n445 256.663
R619 B.n657 B.n446 256.663
R620 B.n657 B.n447 256.663
R621 B.n657 B.n448 256.663
R622 B.n657 B.n449 256.663
R623 B.n664 B.n396 163.367
R624 B.n664 B.n394 163.367
R625 B.n668 B.n394 163.367
R626 B.n668 B.n388 163.367
R627 B.n676 B.n388 163.367
R628 B.n676 B.n386 163.367
R629 B.n680 B.n386 163.367
R630 B.n680 B.n380 163.367
R631 B.n688 B.n380 163.367
R632 B.n688 B.n378 163.367
R633 B.n692 B.n378 163.367
R634 B.n692 B.n372 163.367
R635 B.n700 B.n372 163.367
R636 B.n700 B.n370 163.367
R637 B.n704 B.n370 163.367
R638 B.n704 B.n364 163.367
R639 B.n713 B.n364 163.367
R640 B.n713 B.n362 163.367
R641 B.n717 B.n362 163.367
R642 B.n717 B.n357 163.367
R643 B.n725 B.n357 163.367
R644 B.n725 B.n355 163.367
R645 B.n729 B.n355 163.367
R646 B.n729 B.n349 163.367
R647 B.n737 B.n349 163.367
R648 B.n737 B.n347 163.367
R649 B.n741 B.n347 163.367
R650 B.n741 B.n341 163.367
R651 B.n749 B.n341 163.367
R652 B.n749 B.n339 163.367
R653 B.n753 B.n339 163.367
R654 B.n753 B.n333 163.367
R655 B.n762 B.n333 163.367
R656 B.n762 B.n331 163.367
R657 B.n766 B.n331 163.367
R658 B.n766 B.n2 163.367
R659 B.n896 B.n2 163.367
R660 B.n896 B.n3 163.367
R661 B.n892 B.n3 163.367
R662 B.n892 B.n9 163.367
R663 B.n888 B.n9 163.367
R664 B.n888 B.n11 163.367
R665 B.n884 B.n11 163.367
R666 B.n884 B.n16 163.367
R667 B.n880 B.n16 163.367
R668 B.n880 B.n18 163.367
R669 B.n876 B.n18 163.367
R670 B.n876 B.n23 163.367
R671 B.n872 B.n23 163.367
R672 B.n872 B.n25 163.367
R673 B.n868 B.n25 163.367
R674 B.n868 B.n30 163.367
R675 B.n864 B.n30 163.367
R676 B.n864 B.n32 163.367
R677 B.n860 B.n32 163.367
R678 B.n860 B.n36 163.367
R679 B.n856 B.n36 163.367
R680 B.n856 B.n38 163.367
R681 B.n852 B.n38 163.367
R682 B.n852 B.n44 163.367
R683 B.n848 B.n44 163.367
R684 B.n848 B.n46 163.367
R685 B.n844 B.n46 163.367
R686 B.n844 B.n51 163.367
R687 B.n840 B.n51 163.367
R688 B.n840 B.n53 163.367
R689 B.n836 B.n53 163.367
R690 B.n836 B.n58 163.367
R691 B.n832 B.n58 163.367
R692 B.n832 B.n60 163.367
R693 B.n828 B.n60 163.367
R694 B.n828 B.n65 163.367
R695 B.n824 B.n65 163.367
R696 B.n824 B.n67 163.367
R697 B.n451 B.n450 163.367
R698 B.n650 B.n450 163.367
R699 B.n648 B.n647 163.367
R700 B.n644 B.n643 163.367
R701 B.n640 B.n639 163.367
R702 B.n636 B.n635 163.367
R703 B.n632 B.n631 163.367
R704 B.n628 B.n627 163.367
R705 B.n624 B.n623 163.367
R706 B.n620 B.n619 163.367
R707 B.n616 B.n615 163.367
R708 B.n612 B.n611 163.367
R709 B.n608 B.n607 163.367
R710 B.n604 B.n603 163.367
R711 B.n600 B.n599 163.367
R712 B.n596 B.n595 163.367
R713 B.n592 B.n591 163.367
R714 B.n588 B.n587 163.367
R715 B.n584 B.n583 163.367
R716 B.n580 B.n579 163.367
R717 B.n576 B.n575 163.367
R718 B.n572 B.n571 163.367
R719 B.n568 B.n567 163.367
R720 B.n563 B.n562 163.367
R721 B.n559 B.n558 163.367
R722 B.n555 B.n554 163.367
R723 B.n551 B.n550 163.367
R724 B.n547 B.n546 163.367
R725 B.n542 B.n541 163.367
R726 B.n538 B.n537 163.367
R727 B.n534 B.n533 163.367
R728 B.n530 B.n529 163.367
R729 B.n526 B.n525 163.367
R730 B.n522 B.n521 163.367
R731 B.n518 B.n517 163.367
R732 B.n514 B.n513 163.367
R733 B.n510 B.n509 163.367
R734 B.n506 B.n505 163.367
R735 B.n502 B.n501 163.367
R736 B.n498 B.n497 163.367
R737 B.n494 B.n493 163.367
R738 B.n490 B.n489 163.367
R739 B.n486 B.n485 163.367
R740 B.n482 B.n481 163.367
R741 B.n478 B.n477 163.367
R742 B.n474 B.n473 163.367
R743 B.n470 B.n469 163.367
R744 B.n466 B.n465 163.367
R745 B.n462 B.n461 163.367
R746 B.n458 B.n457 163.367
R747 B.n658 B.n400 163.367
R748 B.n662 B.n398 163.367
R749 B.n662 B.n392 163.367
R750 B.n670 B.n392 163.367
R751 B.n670 B.n390 163.367
R752 B.n674 B.n390 163.367
R753 B.n674 B.n384 163.367
R754 B.n682 B.n384 163.367
R755 B.n682 B.n382 163.367
R756 B.n686 B.n382 163.367
R757 B.n686 B.n376 163.367
R758 B.n694 B.n376 163.367
R759 B.n694 B.n374 163.367
R760 B.n698 B.n374 163.367
R761 B.n698 B.n368 163.367
R762 B.n706 B.n368 163.367
R763 B.n706 B.n366 163.367
R764 B.n710 B.n366 163.367
R765 B.n710 B.n361 163.367
R766 B.n719 B.n361 163.367
R767 B.n719 B.n359 163.367
R768 B.n723 B.n359 163.367
R769 B.n723 B.n353 163.367
R770 B.n731 B.n353 163.367
R771 B.n731 B.n351 163.367
R772 B.n735 B.n351 163.367
R773 B.n735 B.n344 163.367
R774 B.n743 B.n344 163.367
R775 B.n743 B.n342 163.367
R776 B.n747 B.n342 163.367
R777 B.n747 B.n336 163.367
R778 B.n755 B.n336 163.367
R779 B.n755 B.n334 163.367
R780 B.n760 B.n334 163.367
R781 B.n760 B.n329 163.367
R782 B.n768 B.n329 163.367
R783 B.n769 B.n768 163.367
R784 B.n769 B.n5 163.367
R785 B.n6 B.n5 163.367
R786 B.n7 B.n6 163.367
R787 B.n774 B.n7 163.367
R788 B.n774 B.n12 163.367
R789 B.n13 B.n12 163.367
R790 B.n14 B.n13 163.367
R791 B.n779 B.n14 163.367
R792 B.n779 B.n19 163.367
R793 B.n20 B.n19 163.367
R794 B.n21 B.n20 163.367
R795 B.n784 B.n21 163.367
R796 B.n784 B.n26 163.367
R797 B.n27 B.n26 163.367
R798 B.n28 B.n27 163.367
R799 B.n789 B.n28 163.367
R800 B.n789 B.n33 163.367
R801 B.n34 B.n33 163.367
R802 B.n35 B.n34 163.367
R803 B.n794 B.n35 163.367
R804 B.n794 B.n40 163.367
R805 B.n41 B.n40 163.367
R806 B.n42 B.n41 163.367
R807 B.n799 B.n42 163.367
R808 B.n799 B.n47 163.367
R809 B.n48 B.n47 163.367
R810 B.n49 B.n48 163.367
R811 B.n804 B.n49 163.367
R812 B.n804 B.n54 163.367
R813 B.n55 B.n54 163.367
R814 B.n56 B.n55 163.367
R815 B.n809 B.n56 163.367
R816 B.n809 B.n61 163.367
R817 B.n62 B.n61 163.367
R818 B.n63 B.n62 163.367
R819 B.n814 B.n63 163.367
R820 B.n814 B.n68 163.367
R821 B.n69 B.n68 163.367
R822 B.n131 B.n130 163.367
R823 B.n135 B.n134 163.367
R824 B.n139 B.n138 163.367
R825 B.n143 B.n142 163.367
R826 B.n147 B.n146 163.367
R827 B.n151 B.n150 163.367
R828 B.n155 B.n154 163.367
R829 B.n159 B.n158 163.367
R830 B.n163 B.n162 163.367
R831 B.n167 B.n166 163.367
R832 B.n171 B.n170 163.367
R833 B.n175 B.n174 163.367
R834 B.n179 B.n178 163.367
R835 B.n183 B.n182 163.367
R836 B.n187 B.n186 163.367
R837 B.n191 B.n190 163.367
R838 B.n195 B.n194 163.367
R839 B.n199 B.n198 163.367
R840 B.n203 B.n202 163.367
R841 B.n207 B.n206 163.367
R842 B.n211 B.n210 163.367
R843 B.n215 B.n214 163.367
R844 B.n219 B.n218 163.367
R845 B.n223 B.n222 163.367
R846 B.n227 B.n226 163.367
R847 B.n231 B.n230 163.367
R848 B.n235 B.n234 163.367
R849 B.n239 B.n238 163.367
R850 B.n243 B.n242 163.367
R851 B.n247 B.n246 163.367
R852 B.n251 B.n250 163.367
R853 B.n255 B.n254 163.367
R854 B.n259 B.n258 163.367
R855 B.n263 B.n262 163.367
R856 B.n267 B.n266 163.367
R857 B.n271 B.n270 163.367
R858 B.n275 B.n274 163.367
R859 B.n279 B.n278 163.367
R860 B.n283 B.n282 163.367
R861 B.n287 B.n286 163.367
R862 B.n291 B.n290 163.367
R863 B.n295 B.n294 163.367
R864 B.n299 B.n298 163.367
R865 B.n303 B.n302 163.367
R866 B.n307 B.n306 163.367
R867 B.n311 B.n310 163.367
R868 B.n315 B.n314 163.367
R869 B.n319 B.n318 163.367
R870 B.n323 B.n322 163.367
R871 B.n325 B.n120 163.367
R872 B.n657 B.n397 81.0501
R873 B.n822 B.n821 81.0501
R874 B.n656 B.n655 71.676
R875 B.n650 B.n401 71.676
R876 B.n647 B.n402 71.676
R877 B.n643 B.n403 71.676
R878 B.n639 B.n404 71.676
R879 B.n635 B.n405 71.676
R880 B.n631 B.n406 71.676
R881 B.n627 B.n407 71.676
R882 B.n623 B.n408 71.676
R883 B.n619 B.n409 71.676
R884 B.n615 B.n410 71.676
R885 B.n611 B.n411 71.676
R886 B.n607 B.n412 71.676
R887 B.n603 B.n413 71.676
R888 B.n599 B.n414 71.676
R889 B.n595 B.n415 71.676
R890 B.n591 B.n416 71.676
R891 B.n587 B.n417 71.676
R892 B.n583 B.n418 71.676
R893 B.n579 B.n419 71.676
R894 B.n575 B.n420 71.676
R895 B.n571 B.n421 71.676
R896 B.n567 B.n422 71.676
R897 B.n562 B.n423 71.676
R898 B.n558 B.n424 71.676
R899 B.n554 B.n425 71.676
R900 B.n550 B.n426 71.676
R901 B.n546 B.n427 71.676
R902 B.n541 B.n428 71.676
R903 B.n537 B.n429 71.676
R904 B.n533 B.n430 71.676
R905 B.n529 B.n431 71.676
R906 B.n525 B.n432 71.676
R907 B.n521 B.n433 71.676
R908 B.n517 B.n434 71.676
R909 B.n513 B.n435 71.676
R910 B.n509 B.n436 71.676
R911 B.n505 B.n437 71.676
R912 B.n501 B.n438 71.676
R913 B.n497 B.n439 71.676
R914 B.n493 B.n440 71.676
R915 B.n489 B.n441 71.676
R916 B.n485 B.n442 71.676
R917 B.n481 B.n443 71.676
R918 B.n477 B.n444 71.676
R919 B.n473 B.n445 71.676
R920 B.n469 B.n446 71.676
R921 B.n465 B.n447 71.676
R922 B.n461 B.n448 71.676
R923 B.n457 B.n449 71.676
R924 B.n127 B.n70 71.676
R925 B.n131 B.n71 71.676
R926 B.n135 B.n72 71.676
R927 B.n139 B.n73 71.676
R928 B.n143 B.n74 71.676
R929 B.n147 B.n75 71.676
R930 B.n151 B.n76 71.676
R931 B.n155 B.n77 71.676
R932 B.n159 B.n78 71.676
R933 B.n163 B.n79 71.676
R934 B.n167 B.n80 71.676
R935 B.n171 B.n81 71.676
R936 B.n175 B.n82 71.676
R937 B.n179 B.n83 71.676
R938 B.n183 B.n84 71.676
R939 B.n187 B.n85 71.676
R940 B.n191 B.n86 71.676
R941 B.n195 B.n87 71.676
R942 B.n199 B.n88 71.676
R943 B.n203 B.n89 71.676
R944 B.n207 B.n90 71.676
R945 B.n211 B.n91 71.676
R946 B.n215 B.n92 71.676
R947 B.n219 B.n93 71.676
R948 B.n223 B.n94 71.676
R949 B.n227 B.n95 71.676
R950 B.n231 B.n96 71.676
R951 B.n235 B.n97 71.676
R952 B.n239 B.n98 71.676
R953 B.n243 B.n99 71.676
R954 B.n247 B.n100 71.676
R955 B.n251 B.n101 71.676
R956 B.n255 B.n102 71.676
R957 B.n259 B.n103 71.676
R958 B.n263 B.n104 71.676
R959 B.n267 B.n105 71.676
R960 B.n271 B.n106 71.676
R961 B.n275 B.n107 71.676
R962 B.n279 B.n108 71.676
R963 B.n283 B.n109 71.676
R964 B.n287 B.n110 71.676
R965 B.n291 B.n111 71.676
R966 B.n295 B.n112 71.676
R967 B.n299 B.n113 71.676
R968 B.n303 B.n114 71.676
R969 B.n307 B.n115 71.676
R970 B.n311 B.n116 71.676
R971 B.n315 B.n117 71.676
R972 B.n319 B.n118 71.676
R973 B.n323 B.n119 71.676
R974 B.n820 B.n120 71.676
R975 B.n820 B.n819 71.676
R976 B.n325 B.n119 71.676
R977 B.n322 B.n118 71.676
R978 B.n318 B.n117 71.676
R979 B.n314 B.n116 71.676
R980 B.n310 B.n115 71.676
R981 B.n306 B.n114 71.676
R982 B.n302 B.n113 71.676
R983 B.n298 B.n112 71.676
R984 B.n294 B.n111 71.676
R985 B.n290 B.n110 71.676
R986 B.n286 B.n109 71.676
R987 B.n282 B.n108 71.676
R988 B.n278 B.n107 71.676
R989 B.n274 B.n106 71.676
R990 B.n270 B.n105 71.676
R991 B.n266 B.n104 71.676
R992 B.n262 B.n103 71.676
R993 B.n258 B.n102 71.676
R994 B.n254 B.n101 71.676
R995 B.n250 B.n100 71.676
R996 B.n246 B.n99 71.676
R997 B.n242 B.n98 71.676
R998 B.n238 B.n97 71.676
R999 B.n234 B.n96 71.676
R1000 B.n230 B.n95 71.676
R1001 B.n226 B.n94 71.676
R1002 B.n222 B.n93 71.676
R1003 B.n218 B.n92 71.676
R1004 B.n214 B.n91 71.676
R1005 B.n210 B.n90 71.676
R1006 B.n206 B.n89 71.676
R1007 B.n202 B.n88 71.676
R1008 B.n198 B.n87 71.676
R1009 B.n194 B.n86 71.676
R1010 B.n190 B.n85 71.676
R1011 B.n186 B.n84 71.676
R1012 B.n182 B.n83 71.676
R1013 B.n178 B.n82 71.676
R1014 B.n174 B.n81 71.676
R1015 B.n170 B.n80 71.676
R1016 B.n166 B.n79 71.676
R1017 B.n162 B.n78 71.676
R1018 B.n158 B.n77 71.676
R1019 B.n154 B.n76 71.676
R1020 B.n150 B.n75 71.676
R1021 B.n146 B.n74 71.676
R1022 B.n142 B.n73 71.676
R1023 B.n138 B.n72 71.676
R1024 B.n134 B.n71 71.676
R1025 B.n130 B.n70 71.676
R1026 B.n656 B.n451 71.676
R1027 B.n648 B.n401 71.676
R1028 B.n644 B.n402 71.676
R1029 B.n640 B.n403 71.676
R1030 B.n636 B.n404 71.676
R1031 B.n632 B.n405 71.676
R1032 B.n628 B.n406 71.676
R1033 B.n624 B.n407 71.676
R1034 B.n620 B.n408 71.676
R1035 B.n616 B.n409 71.676
R1036 B.n612 B.n410 71.676
R1037 B.n608 B.n411 71.676
R1038 B.n604 B.n412 71.676
R1039 B.n600 B.n413 71.676
R1040 B.n596 B.n414 71.676
R1041 B.n592 B.n415 71.676
R1042 B.n588 B.n416 71.676
R1043 B.n584 B.n417 71.676
R1044 B.n580 B.n418 71.676
R1045 B.n576 B.n419 71.676
R1046 B.n572 B.n420 71.676
R1047 B.n568 B.n421 71.676
R1048 B.n563 B.n422 71.676
R1049 B.n559 B.n423 71.676
R1050 B.n555 B.n424 71.676
R1051 B.n551 B.n425 71.676
R1052 B.n547 B.n426 71.676
R1053 B.n542 B.n427 71.676
R1054 B.n538 B.n428 71.676
R1055 B.n534 B.n429 71.676
R1056 B.n530 B.n430 71.676
R1057 B.n526 B.n431 71.676
R1058 B.n522 B.n432 71.676
R1059 B.n518 B.n433 71.676
R1060 B.n514 B.n434 71.676
R1061 B.n510 B.n435 71.676
R1062 B.n506 B.n436 71.676
R1063 B.n502 B.n437 71.676
R1064 B.n498 B.n438 71.676
R1065 B.n494 B.n439 71.676
R1066 B.n490 B.n440 71.676
R1067 B.n486 B.n441 71.676
R1068 B.n482 B.n442 71.676
R1069 B.n478 B.n443 71.676
R1070 B.n474 B.n444 71.676
R1071 B.n470 B.n445 71.676
R1072 B.n466 B.n446 71.676
R1073 B.n462 B.n447 71.676
R1074 B.n458 B.n448 71.676
R1075 B.n449 B.n400 71.676
R1076 B.n544 B.n455 59.5399
R1077 B.n565 B.n453 59.5399
R1078 B.n126 B.n125 59.5399
R1079 B.n123 B.n122 59.5399
R1080 B.n663 B.n397 39.6506
R1081 B.n663 B.n393 39.6506
R1082 B.n669 B.n393 39.6506
R1083 B.n669 B.n389 39.6506
R1084 B.n675 B.n389 39.6506
R1085 B.n681 B.n385 39.6506
R1086 B.n681 B.n381 39.6506
R1087 B.n687 B.n381 39.6506
R1088 B.n687 B.n377 39.6506
R1089 B.n693 B.n377 39.6506
R1090 B.n693 B.n373 39.6506
R1091 B.n699 B.n373 39.6506
R1092 B.n705 B.n369 39.6506
R1093 B.n705 B.n365 39.6506
R1094 B.n712 B.n365 39.6506
R1095 B.n712 B.n711 39.6506
R1096 B.n718 B.n358 39.6506
R1097 B.n724 B.n358 39.6506
R1098 B.n724 B.n354 39.6506
R1099 B.n730 B.n354 39.6506
R1100 B.n736 B.n350 39.6506
R1101 B.n736 B.n345 39.6506
R1102 B.n742 B.n345 39.6506
R1103 B.n742 B.n346 39.6506
R1104 B.n748 B.n337 39.6506
R1105 B.n754 B.n337 39.6506
R1106 B.n754 B.n338 39.6506
R1107 B.n761 B.n330 39.6506
R1108 B.n767 B.n330 39.6506
R1109 B.n767 B.n4 39.6506
R1110 B.n895 B.n4 39.6506
R1111 B.n895 B.n894 39.6506
R1112 B.n894 B.n893 39.6506
R1113 B.n893 B.n8 39.6506
R1114 B.n887 B.n8 39.6506
R1115 B.n886 B.n885 39.6506
R1116 B.n885 B.n15 39.6506
R1117 B.n879 B.n15 39.6506
R1118 B.n878 B.n877 39.6506
R1119 B.n877 B.n22 39.6506
R1120 B.n871 B.n22 39.6506
R1121 B.n871 B.n870 39.6506
R1122 B.n869 B.n29 39.6506
R1123 B.n863 B.n29 39.6506
R1124 B.n863 B.n862 39.6506
R1125 B.n862 B.n861 39.6506
R1126 B.n855 B.n39 39.6506
R1127 B.n855 B.n854 39.6506
R1128 B.n854 B.n853 39.6506
R1129 B.n853 B.n43 39.6506
R1130 B.n847 B.n846 39.6506
R1131 B.n846 B.n845 39.6506
R1132 B.n845 B.n50 39.6506
R1133 B.n839 B.n50 39.6506
R1134 B.n839 B.n838 39.6506
R1135 B.n838 B.n837 39.6506
R1136 B.n837 B.n57 39.6506
R1137 B.n831 B.n830 39.6506
R1138 B.n830 B.n829 39.6506
R1139 B.n829 B.n64 39.6506
R1140 B.n823 B.n64 39.6506
R1141 B.n823 B.n822 39.6506
R1142 B.n338 B.t8 38.4845
R1143 B.t7 B.n886 38.4845
R1144 B.n818 B.n817 35.7468
R1145 B.n128 B.n66 35.7468
R1146 B.n660 B.n659 35.7468
R1147 B.n654 B.n395 35.7468
R1148 B.n748 B.t0 34.9859
R1149 B.n879 B.t3 34.9859
R1150 B.n455 B.n454 32.0005
R1151 B.n453 B.n452 32.0005
R1152 B.n125 B.n124 32.0005
R1153 B.n122 B.n121 32.0005
R1154 B.t1 B.n350 29.155
R1155 B.n870 B.t5 29.155
R1156 B.n718 B.t4 23.3241
R1157 B.n861 B.t9 23.3241
R1158 B.n699 B.t6 22.1579
R1159 B.n847 B.t2 22.1579
R1160 B.n675 B.t11 19.8256
R1161 B.t11 B.n385 19.8256
R1162 B.t15 B.n57 19.8256
R1163 B.n831 B.t15 19.8256
R1164 B B.n897 18.0485
R1165 B.t6 B.n369 17.4932
R1166 B.t2 B.n43 17.4932
R1167 B.n711 B.t4 16.327
R1168 B.n39 B.t9 16.327
R1169 B.n129 B.n128 10.6151
R1170 B.n132 B.n129 10.6151
R1171 B.n133 B.n132 10.6151
R1172 B.n136 B.n133 10.6151
R1173 B.n137 B.n136 10.6151
R1174 B.n140 B.n137 10.6151
R1175 B.n141 B.n140 10.6151
R1176 B.n144 B.n141 10.6151
R1177 B.n145 B.n144 10.6151
R1178 B.n148 B.n145 10.6151
R1179 B.n149 B.n148 10.6151
R1180 B.n152 B.n149 10.6151
R1181 B.n153 B.n152 10.6151
R1182 B.n156 B.n153 10.6151
R1183 B.n157 B.n156 10.6151
R1184 B.n160 B.n157 10.6151
R1185 B.n161 B.n160 10.6151
R1186 B.n164 B.n161 10.6151
R1187 B.n165 B.n164 10.6151
R1188 B.n168 B.n165 10.6151
R1189 B.n169 B.n168 10.6151
R1190 B.n172 B.n169 10.6151
R1191 B.n173 B.n172 10.6151
R1192 B.n176 B.n173 10.6151
R1193 B.n177 B.n176 10.6151
R1194 B.n180 B.n177 10.6151
R1195 B.n181 B.n180 10.6151
R1196 B.n184 B.n181 10.6151
R1197 B.n185 B.n184 10.6151
R1198 B.n188 B.n185 10.6151
R1199 B.n189 B.n188 10.6151
R1200 B.n192 B.n189 10.6151
R1201 B.n193 B.n192 10.6151
R1202 B.n196 B.n193 10.6151
R1203 B.n197 B.n196 10.6151
R1204 B.n200 B.n197 10.6151
R1205 B.n201 B.n200 10.6151
R1206 B.n204 B.n201 10.6151
R1207 B.n205 B.n204 10.6151
R1208 B.n208 B.n205 10.6151
R1209 B.n209 B.n208 10.6151
R1210 B.n212 B.n209 10.6151
R1211 B.n213 B.n212 10.6151
R1212 B.n216 B.n213 10.6151
R1213 B.n217 B.n216 10.6151
R1214 B.n221 B.n220 10.6151
R1215 B.n224 B.n221 10.6151
R1216 B.n225 B.n224 10.6151
R1217 B.n228 B.n225 10.6151
R1218 B.n229 B.n228 10.6151
R1219 B.n232 B.n229 10.6151
R1220 B.n233 B.n232 10.6151
R1221 B.n236 B.n233 10.6151
R1222 B.n237 B.n236 10.6151
R1223 B.n241 B.n240 10.6151
R1224 B.n244 B.n241 10.6151
R1225 B.n245 B.n244 10.6151
R1226 B.n248 B.n245 10.6151
R1227 B.n249 B.n248 10.6151
R1228 B.n252 B.n249 10.6151
R1229 B.n253 B.n252 10.6151
R1230 B.n256 B.n253 10.6151
R1231 B.n257 B.n256 10.6151
R1232 B.n260 B.n257 10.6151
R1233 B.n261 B.n260 10.6151
R1234 B.n264 B.n261 10.6151
R1235 B.n265 B.n264 10.6151
R1236 B.n268 B.n265 10.6151
R1237 B.n269 B.n268 10.6151
R1238 B.n272 B.n269 10.6151
R1239 B.n273 B.n272 10.6151
R1240 B.n276 B.n273 10.6151
R1241 B.n277 B.n276 10.6151
R1242 B.n280 B.n277 10.6151
R1243 B.n281 B.n280 10.6151
R1244 B.n284 B.n281 10.6151
R1245 B.n285 B.n284 10.6151
R1246 B.n288 B.n285 10.6151
R1247 B.n289 B.n288 10.6151
R1248 B.n292 B.n289 10.6151
R1249 B.n293 B.n292 10.6151
R1250 B.n296 B.n293 10.6151
R1251 B.n297 B.n296 10.6151
R1252 B.n300 B.n297 10.6151
R1253 B.n301 B.n300 10.6151
R1254 B.n304 B.n301 10.6151
R1255 B.n305 B.n304 10.6151
R1256 B.n308 B.n305 10.6151
R1257 B.n309 B.n308 10.6151
R1258 B.n312 B.n309 10.6151
R1259 B.n313 B.n312 10.6151
R1260 B.n316 B.n313 10.6151
R1261 B.n317 B.n316 10.6151
R1262 B.n320 B.n317 10.6151
R1263 B.n321 B.n320 10.6151
R1264 B.n324 B.n321 10.6151
R1265 B.n326 B.n324 10.6151
R1266 B.n327 B.n326 10.6151
R1267 B.n818 B.n327 10.6151
R1268 B.n661 B.n660 10.6151
R1269 B.n661 B.n391 10.6151
R1270 B.n671 B.n391 10.6151
R1271 B.n672 B.n671 10.6151
R1272 B.n673 B.n672 10.6151
R1273 B.n673 B.n383 10.6151
R1274 B.n683 B.n383 10.6151
R1275 B.n684 B.n683 10.6151
R1276 B.n685 B.n684 10.6151
R1277 B.n685 B.n375 10.6151
R1278 B.n695 B.n375 10.6151
R1279 B.n696 B.n695 10.6151
R1280 B.n697 B.n696 10.6151
R1281 B.n697 B.n367 10.6151
R1282 B.n707 B.n367 10.6151
R1283 B.n708 B.n707 10.6151
R1284 B.n709 B.n708 10.6151
R1285 B.n709 B.n360 10.6151
R1286 B.n720 B.n360 10.6151
R1287 B.n721 B.n720 10.6151
R1288 B.n722 B.n721 10.6151
R1289 B.n722 B.n352 10.6151
R1290 B.n732 B.n352 10.6151
R1291 B.n733 B.n732 10.6151
R1292 B.n734 B.n733 10.6151
R1293 B.n734 B.n343 10.6151
R1294 B.n744 B.n343 10.6151
R1295 B.n745 B.n744 10.6151
R1296 B.n746 B.n745 10.6151
R1297 B.n746 B.n335 10.6151
R1298 B.n756 B.n335 10.6151
R1299 B.n757 B.n756 10.6151
R1300 B.n759 B.n757 10.6151
R1301 B.n759 B.n758 10.6151
R1302 B.n758 B.n328 10.6151
R1303 B.n770 B.n328 10.6151
R1304 B.n771 B.n770 10.6151
R1305 B.n772 B.n771 10.6151
R1306 B.n773 B.n772 10.6151
R1307 B.n775 B.n773 10.6151
R1308 B.n776 B.n775 10.6151
R1309 B.n777 B.n776 10.6151
R1310 B.n778 B.n777 10.6151
R1311 B.n780 B.n778 10.6151
R1312 B.n781 B.n780 10.6151
R1313 B.n782 B.n781 10.6151
R1314 B.n783 B.n782 10.6151
R1315 B.n785 B.n783 10.6151
R1316 B.n786 B.n785 10.6151
R1317 B.n787 B.n786 10.6151
R1318 B.n788 B.n787 10.6151
R1319 B.n790 B.n788 10.6151
R1320 B.n791 B.n790 10.6151
R1321 B.n792 B.n791 10.6151
R1322 B.n793 B.n792 10.6151
R1323 B.n795 B.n793 10.6151
R1324 B.n796 B.n795 10.6151
R1325 B.n797 B.n796 10.6151
R1326 B.n798 B.n797 10.6151
R1327 B.n800 B.n798 10.6151
R1328 B.n801 B.n800 10.6151
R1329 B.n802 B.n801 10.6151
R1330 B.n803 B.n802 10.6151
R1331 B.n805 B.n803 10.6151
R1332 B.n806 B.n805 10.6151
R1333 B.n807 B.n806 10.6151
R1334 B.n808 B.n807 10.6151
R1335 B.n810 B.n808 10.6151
R1336 B.n811 B.n810 10.6151
R1337 B.n812 B.n811 10.6151
R1338 B.n813 B.n812 10.6151
R1339 B.n815 B.n813 10.6151
R1340 B.n816 B.n815 10.6151
R1341 B.n817 B.n816 10.6151
R1342 B.n654 B.n653 10.6151
R1343 B.n653 B.n652 10.6151
R1344 B.n652 B.n651 10.6151
R1345 B.n651 B.n649 10.6151
R1346 B.n649 B.n646 10.6151
R1347 B.n646 B.n645 10.6151
R1348 B.n645 B.n642 10.6151
R1349 B.n642 B.n641 10.6151
R1350 B.n641 B.n638 10.6151
R1351 B.n638 B.n637 10.6151
R1352 B.n637 B.n634 10.6151
R1353 B.n634 B.n633 10.6151
R1354 B.n633 B.n630 10.6151
R1355 B.n630 B.n629 10.6151
R1356 B.n629 B.n626 10.6151
R1357 B.n626 B.n625 10.6151
R1358 B.n625 B.n622 10.6151
R1359 B.n622 B.n621 10.6151
R1360 B.n621 B.n618 10.6151
R1361 B.n618 B.n617 10.6151
R1362 B.n617 B.n614 10.6151
R1363 B.n614 B.n613 10.6151
R1364 B.n613 B.n610 10.6151
R1365 B.n610 B.n609 10.6151
R1366 B.n609 B.n606 10.6151
R1367 B.n606 B.n605 10.6151
R1368 B.n605 B.n602 10.6151
R1369 B.n602 B.n601 10.6151
R1370 B.n601 B.n598 10.6151
R1371 B.n598 B.n597 10.6151
R1372 B.n597 B.n594 10.6151
R1373 B.n594 B.n593 10.6151
R1374 B.n593 B.n590 10.6151
R1375 B.n590 B.n589 10.6151
R1376 B.n589 B.n586 10.6151
R1377 B.n586 B.n585 10.6151
R1378 B.n585 B.n582 10.6151
R1379 B.n582 B.n581 10.6151
R1380 B.n581 B.n578 10.6151
R1381 B.n578 B.n577 10.6151
R1382 B.n577 B.n574 10.6151
R1383 B.n574 B.n573 10.6151
R1384 B.n573 B.n570 10.6151
R1385 B.n570 B.n569 10.6151
R1386 B.n569 B.n566 10.6151
R1387 B.n564 B.n561 10.6151
R1388 B.n561 B.n560 10.6151
R1389 B.n560 B.n557 10.6151
R1390 B.n557 B.n556 10.6151
R1391 B.n556 B.n553 10.6151
R1392 B.n553 B.n552 10.6151
R1393 B.n552 B.n549 10.6151
R1394 B.n549 B.n548 10.6151
R1395 B.n548 B.n545 10.6151
R1396 B.n543 B.n540 10.6151
R1397 B.n540 B.n539 10.6151
R1398 B.n539 B.n536 10.6151
R1399 B.n536 B.n535 10.6151
R1400 B.n535 B.n532 10.6151
R1401 B.n532 B.n531 10.6151
R1402 B.n531 B.n528 10.6151
R1403 B.n528 B.n527 10.6151
R1404 B.n527 B.n524 10.6151
R1405 B.n524 B.n523 10.6151
R1406 B.n523 B.n520 10.6151
R1407 B.n520 B.n519 10.6151
R1408 B.n519 B.n516 10.6151
R1409 B.n516 B.n515 10.6151
R1410 B.n515 B.n512 10.6151
R1411 B.n512 B.n511 10.6151
R1412 B.n511 B.n508 10.6151
R1413 B.n508 B.n507 10.6151
R1414 B.n507 B.n504 10.6151
R1415 B.n504 B.n503 10.6151
R1416 B.n503 B.n500 10.6151
R1417 B.n500 B.n499 10.6151
R1418 B.n499 B.n496 10.6151
R1419 B.n496 B.n495 10.6151
R1420 B.n495 B.n492 10.6151
R1421 B.n492 B.n491 10.6151
R1422 B.n491 B.n488 10.6151
R1423 B.n488 B.n487 10.6151
R1424 B.n487 B.n484 10.6151
R1425 B.n484 B.n483 10.6151
R1426 B.n483 B.n480 10.6151
R1427 B.n480 B.n479 10.6151
R1428 B.n479 B.n476 10.6151
R1429 B.n476 B.n475 10.6151
R1430 B.n475 B.n472 10.6151
R1431 B.n472 B.n471 10.6151
R1432 B.n471 B.n468 10.6151
R1433 B.n468 B.n467 10.6151
R1434 B.n467 B.n464 10.6151
R1435 B.n464 B.n463 10.6151
R1436 B.n463 B.n460 10.6151
R1437 B.n460 B.n459 10.6151
R1438 B.n459 B.n456 10.6151
R1439 B.n456 B.n399 10.6151
R1440 B.n659 B.n399 10.6151
R1441 B.n665 B.n395 10.6151
R1442 B.n666 B.n665 10.6151
R1443 B.n667 B.n666 10.6151
R1444 B.n667 B.n387 10.6151
R1445 B.n677 B.n387 10.6151
R1446 B.n678 B.n677 10.6151
R1447 B.n679 B.n678 10.6151
R1448 B.n679 B.n379 10.6151
R1449 B.n689 B.n379 10.6151
R1450 B.n690 B.n689 10.6151
R1451 B.n691 B.n690 10.6151
R1452 B.n691 B.n371 10.6151
R1453 B.n701 B.n371 10.6151
R1454 B.n702 B.n701 10.6151
R1455 B.n703 B.n702 10.6151
R1456 B.n703 B.n363 10.6151
R1457 B.n714 B.n363 10.6151
R1458 B.n715 B.n714 10.6151
R1459 B.n716 B.n715 10.6151
R1460 B.n716 B.n356 10.6151
R1461 B.n726 B.n356 10.6151
R1462 B.n727 B.n726 10.6151
R1463 B.n728 B.n727 10.6151
R1464 B.n728 B.n348 10.6151
R1465 B.n738 B.n348 10.6151
R1466 B.n739 B.n738 10.6151
R1467 B.n740 B.n739 10.6151
R1468 B.n740 B.n340 10.6151
R1469 B.n750 B.n340 10.6151
R1470 B.n751 B.n750 10.6151
R1471 B.n752 B.n751 10.6151
R1472 B.n752 B.n332 10.6151
R1473 B.n763 B.n332 10.6151
R1474 B.n764 B.n763 10.6151
R1475 B.n765 B.n764 10.6151
R1476 B.n765 B.n0 10.6151
R1477 B.n891 B.n1 10.6151
R1478 B.n891 B.n890 10.6151
R1479 B.n890 B.n889 10.6151
R1480 B.n889 B.n10 10.6151
R1481 B.n883 B.n10 10.6151
R1482 B.n883 B.n882 10.6151
R1483 B.n882 B.n881 10.6151
R1484 B.n881 B.n17 10.6151
R1485 B.n875 B.n17 10.6151
R1486 B.n875 B.n874 10.6151
R1487 B.n874 B.n873 10.6151
R1488 B.n873 B.n24 10.6151
R1489 B.n867 B.n24 10.6151
R1490 B.n867 B.n866 10.6151
R1491 B.n866 B.n865 10.6151
R1492 B.n865 B.n31 10.6151
R1493 B.n859 B.n31 10.6151
R1494 B.n859 B.n858 10.6151
R1495 B.n858 B.n857 10.6151
R1496 B.n857 B.n37 10.6151
R1497 B.n851 B.n37 10.6151
R1498 B.n851 B.n850 10.6151
R1499 B.n850 B.n849 10.6151
R1500 B.n849 B.n45 10.6151
R1501 B.n843 B.n45 10.6151
R1502 B.n843 B.n842 10.6151
R1503 B.n842 B.n841 10.6151
R1504 B.n841 B.n52 10.6151
R1505 B.n835 B.n52 10.6151
R1506 B.n835 B.n834 10.6151
R1507 B.n834 B.n833 10.6151
R1508 B.n833 B.n59 10.6151
R1509 B.n827 B.n59 10.6151
R1510 B.n827 B.n826 10.6151
R1511 B.n826 B.n825 10.6151
R1512 B.n825 B.n66 10.6151
R1513 B.n730 B.t1 10.4961
R1514 B.t5 B.n869 10.4961
R1515 B.n217 B.n126 9.36635
R1516 B.n240 B.n123 9.36635
R1517 B.n566 B.n565 9.36635
R1518 B.n544 B.n543 9.36635
R1519 B.n346 B.t0 4.66522
R1520 B.t3 B.n878 4.66522
R1521 B.n897 B.n0 2.81026
R1522 B.n897 B.n1 2.81026
R1523 B.n220 B.n126 1.24928
R1524 B.n237 B.n123 1.24928
R1525 B.n565 B.n564 1.24928
R1526 B.n545 B.n544 1.24928
R1527 B.n761 B.t8 1.16668
R1528 B.n887 B.t7 1.16668
R1529 VN.n6 VN.t3 279.103
R1530 VN.n32 VN.t7 279.103
R1531 VN.n3 VN.t1 248.12
R1532 VN.n5 VN.t2 248.12
R1533 VN.n16 VN.t0 248.12
R1534 VN.n23 VN.t6 248.12
R1535 VN.n29 VN.t5 248.12
R1536 VN.n31 VN.t8 248.12
R1537 VN.n28 VN.t9 248.12
R1538 VN.n48 VN.t4 248.12
R1539 VN.n24 VN.n23 171.088
R1540 VN.n49 VN.n48 171.088
R1541 VN.n47 VN.n25 161.3
R1542 VN.n46 VN.n45 161.3
R1543 VN.n44 VN.n26 161.3
R1544 VN.n43 VN.n42 161.3
R1545 VN.n41 VN.n27 161.3
R1546 VN.n40 VN.n39 161.3
R1547 VN.n38 VN.n29 161.3
R1548 VN.n37 VN.n36 161.3
R1549 VN.n35 VN.n30 161.3
R1550 VN.n34 VN.n33 161.3
R1551 VN.n22 VN.n0 161.3
R1552 VN.n21 VN.n20 161.3
R1553 VN.n19 VN.n1 161.3
R1554 VN.n18 VN.n17 161.3
R1555 VN.n15 VN.n2 161.3
R1556 VN.n14 VN.n13 161.3
R1557 VN.n12 VN.n3 161.3
R1558 VN.n11 VN.n10 161.3
R1559 VN.n9 VN.n4 161.3
R1560 VN.n8 VN.n7 161.3
R1561 VN.n6 VN.n5 57.1957
R1562 VN.n32 VN.n31 57.1957
R1563 VN.n10 VN.n9 56.5193
R1564 VN.n15 VN.n14 56.5193
R1565 VN.n36 VN.n35 56.5193
R1566 VN.n41 VN.n40 56.5193
R1567 VN VN.n49 47.6956
R1568 VN.n21 VN.n1 42.9216
R1569 VN.n46 VN.n26 42.9216
R1570 VN.n22 VN.n21 38.0652
R1571 VN.n47 VN.n46 38.0652
R1572 VN.n33 VN.n32 26.7159
R1573 VN.n7 VN.n6 26.7159
R1574 VN.n9 VN.n8 24.4675
R1575 VN.n10 VN.n3 24.4675
R1576 VN.n14 VN.n3 24.4675
R1577 VN.n17 VN.n15 24.4675
R1578 VN.n35 VN.n34 24.4675
R1579 VN.n40 VN.n29 24.4675
R1580 VN.n36 VN.n29 24.4675
R1581 VN.n42 VN.n41 24.4675
R1582 VN.n16 VN.n1 17.1274
R1583 VN.n28 VN.n26 17.1274
R1584 VN.n23 VN.n22 14.6807
R1585 VN.n48 VN.n47 14.6807
R1586 VN.n8 VN.n5 7.3406
R1587 VN.n17 VN.n16 7.3406
R1588 VN.n34 VN.n31 7.3406
R1589 VN.n42 VN.n28 7.3406
R1590 VN.n49 VN.n25 0.189894
R1591 VN.n45 VN.n25 0.189894
R1592 VN.n45 VN.n44 0.189894
R1593 VN.n44 VN.n43 0.189894
R1594 VN.n43 VN.n27 0.189894
R1595 VN.n39 VN.n27 0.189894
R1596 VN.n39 VN.n38 0.189894
R1597 VN.n38 VN.n37 0.189894
R1598 VN.n37 VN.n30 0.189894
R1599 VN.n33 VN.n30 0.189894
R1600 VN.n7 VN.n4 0.189894
R1601 VN.n11 VN.n4 0.189894
R1602 VN.n12 VN.n11 0.189894
R1603 VN.n13 VN.n12 0.189894
R1604 VN.n13 VN.n2 0.189894
R1605 VN.n18 VN.n2 0.189894
R1606 VN.n19 VN.n18 0.189894
R1607 VN.n20 VN.n19 0.189894
R1608 VN.n20 VN.n0 0.189894
R1609 VN.n24 VN.n0 0.189894
R1610 VN VN.n24 0.0516364
R1611 VDD2.n145 VDD2.n77 289.615
R1612 VDD2.n68 VDD2.n0 289.615
R1613 VDD2.n146 VDD2.n145 185
R1614 VDD2.n144 VDD2.n143 185
R1615 VDD2.n81 VDD2.n80 185
R1616 VDD2.n138 VDD2.n137 185
R1617 VDD2.n136 VDD2.n135 185
R1618 VDD2.n85 VDD2.n84 185
R1619 VDD2.n130 VDD2.n129 185
R1620 VDD2.n128 VDD2.n127 185
R1621 VDD2.n89 VDD2.n88 185
R1622 VDD2.n93 VDD2.n91 185
R1623 VDD2.n122 VDD2.n121 185
R1624 VDD2.n120 VDD2.n119 185
R1625 VDD2.n95 VDD2.n94 185
R1626 VDD2.n114 VDD2.n113 185
R1627 VDD2.n112 VDD2.n111 185
R1628 VDD2.n99 VDD2.n98 185
R1629 VDD2.n106 VDD2.n105 185
R1630 VDD2.n104 VDD2.n103 185
R1631 VDD2.n25 VDD2.n24 185
R1632 VDD2.n27 VDD2.n26 185
R1633 VDD2.n20 VDD2.n19 185
R1634 VDD2.n33 VDD2.n32 185
R1635 VDD2.n35 VDD2.n34 185
R1636 VDD2.n16 VDD2.n15 185
R1637 VDD2.n42 VDD2.n41 185
R1638 VDD2.n43 VDD2.n14 185
R1639 VDD2.n45 VDD2.n44 185
R1640 VDD2.n12 VDD2.n11 185
R1641 VDD2.n51 VDD2.n50 185
R1642 VDD2.n53 VDD2.n52 185
R1643 VDD2.n8 VDD2.n7 185
R1644 VDD2.n59 VDD2.n58 185
R1645 VDD2.n61 VDD2.n60 185
R1646 VDD2.n4 VDD2.n3 185
R1647 VDD2.n67 VDD2.n66 185
R1648 VDD2.n69 VDD2.n68 185
R1649 VDD2.n102 VDD2.t0 149.524
R1650 VDD2.n23 VDD2.t3 149.524
R1651 VDD2.n145 VDD2.n144 104.615
R1652 VDD2.n144 VDD2.n80 104.615
R1653 VDD2.n137 VDD2.n80 104.615
R1654 VDD2.n137 VDD2.n136 104.615
R1655 VDD2.n136 VDD2.n84 104.615
R1656 VDD2.n129 VDD2.n84 104.615
R1657 VDD2.n129 VDD2.n128 104.615
R1658 VDD2.n128 VDD2.n88 104.615
R1659 VDD2.n93 VDD2.n88 104.615
R1660 VDD2.n121 VDD2.n93 104.615
R1661 VDD2.n121 VDD2.n120 104.615
R1662 VDD2.n120 VDD2.n94 104.615
R1663 VDD2.n113 VDD2.n94 104.615
R1664 VDD2.n113 VDD2.n112 104.615
R1665 VDD2.n112 VDD2.n98 104.615
R1666 VDD2.n105 VDD2.n98 104.615
R1667 VDD2.n105 VDD2.n104 104.615
R1668 VDD2.n26 VDD2.n25 104.615
R1669 VDD2.n26 VDD2.n19 104.615
R1670 VDD2.n33 VDD2.n19 104.615
R1671 VDD2.n34 VDD2.n33 104.615
R1672 VDD2.n34 VDD2.n15 104.615
R1673 VDD2.n42 VDD2.n15 104.615
R1674 VDD2.n43 VDD2.n42 104.615
R1675 VDD2.n44 VDD2.n43 104.615
R1676 VDD2.n44 VDD2.n11 104.615
R1677 VDD2.n51 VDD2.n11 104.615
R1678 VDD2.n52 VDD2.n51 104.615
R1679 VDD2.n52 VDD2.n7 104.615
R1680 VDD2.n59 VDD2.n7 104.615
R1681 VDD2.n60 VDD2.n59 104.615
R1682 VDD2.n60 VDD2.n3 104.615
R1683 VDD2.n67 VDD2.n3 104.615
R1684 VDD2.n68 VDD2.n67 104.615
R1685 VDD2.n76 VDD2.n75 63.1473
R1686 VDD2 VDD2.n153 63.1444
R1687 VDD2.n152 VDD2.n151 62.136
R1688 VDD2.n74 VDD2.n73 62.1358
R1689 VDD2.n104 VDD2.t0 52.3082
R1690 VDD2.n25 VDD2.t3 52.3082
R1691 VDD2.n74 VDD2.n72 50.8684
R1692 VDD2.n150 VDD2.n149 49.446
R1693 VDD2.n150 VDD2.n76 42.1873
R1694 VDD2.n91 VDD2.n89 13.1884
R1695 VDD2.n45 VDD2.n12 13.1884
R1696 VDD2.n127 VDD2.n126 12.8005
R1697 VDD2.n123 VDD2.n122 12.8005
R1698 VDD2.n46 VDD2.n14 12.8005
R1699 VDD2.n50 VDD2.n49 12.8005
R1700 VDD2.n130 VDD2.n87 12.0247
R1701 VDD2.n119 VDD2.n92 12.0247
R1702 VDD2.n41 VDD2.n40 12.0247
R1703 VDD2.n53 VDD2.n10 12.0247
R1704 VDD2.n131 VDD2.n85 11.249
R1705 VDD2.n118 VDD2.n95 11.249
R1706 VDD2.n39 VDD2.n16 11.249
R1707 VDD2.n54 VDD2.n8 11.249
R1708 VDD2.n135 VDD2.n134 10.4732
R1709 VDD2.n115 VDD2.n114 10.4732
R1710 VDD2.n36 VDD2.n35 10.4732
R1711 VDD2.n58 VDD2.n57 10.4732
R1712 VDD2.n103 VDD2.n102 10.2747
R1713 VDD2.n24 VDD2.n23 10.2747
R1714 VDD2.n138 VDD2.n83 9.69747
R1715 VDD2.n111 VDD2.n97 9.69747
R1716 VDD2.n32 VDD2.n18 9.69747
R1717 VDD2.n61 VDD2.n6 9.69747
R1718 VDD2.n149 VDD2.n148 9.45567
R1719 VDD2.n72 VDD2.n71 9.45567
R1720 VDD2.n101 VDD2.n100 9.3005
R1721 VDD2.n108 VDD2.n107 9.3005
R1722 VDD2.n110 VDD2.n109 9.3005
R1723 VDD2.n97 VDD2.n96 9.3005
R1724 VDD2.n116 VDD2.n115 9.3005
R1725 VDD2.n118 VDD2.n117 9.3005
R1726 VDD2.n92 VDD2.n90 9.3005
R1727 VDD2.n124 VDD2.n123 9.3005
R1728 VDD2.n148 VDD2.n147 9.3005
R1729 VDD2.n79 VDD2.n78 9.3005
R1730 VDD2.n142 VDD2.n141 9.3005
R1731 VDD2.n140 VDD2.n139 9.3005
R1732 VDD2.n83 VDD2.n82 9.3005
R1733 VDD2.n134 VDD2.n133 9.3005
R1734 VDD2.n132 VDD2.n131 9.3005
R1735 VDD2.n87 VDD2.n86 9.3005
R1736 VDD2.n126 VDD2.n125 9.3005
R1737 VDD2.n71 VDD2.n70 9.3005
R1738 VDD2.n65 VDD2.n64 9.3005
R1739 VDD2.n63 VDD2.n62 9.3005
R1740 VDD2.n6 VDD2.n5 9.3005
R1741 VDD2.n57 VDD2.n56 9.3005
R1742 VDD2.n55 VDD2.n54 9.3005
R1743 VDD2.n10 VDD2.n9 9.3005
R1744 VDD2.n49 VDD2.n48 9.3005
R1745 VDD2.n22 VDD2.n21 9.3005
R1746 VDD2.n29 VDD2.n28 9.3005
R1747 VDD2.n31 VDD2.n30 9.3005
R1748 VDD2.n18 VDD2.n17 9.3005
R1749 VDD2.n37 VDD2.n36 9.3005
R1750 VDD2.n39 VDD2.n38 9.3005
R1751 VDD2.n40 VDD2.n13 9.3005
R1752 VDD2.n47 VDD2.n46 9.3005
R1753 VDD2.n2 VDD2.n1 9.3005
R1754 VDD2.n139 VDD2.n81 8.92171
R1755 VDD2.n110 VDD2.n99 8.92171
R1756 VDD2.n31 VDD2.n20 8.92171
R1757 VDD2.n62 VDD2.n4 8.92171
R1758 VDD2.n143 VDD2.n142 8.14595
R1759 VDD2.n107 VDD2.n106 8.14595
R1760 VDD2.n28 VDD2.n27 8.14595
R1761 VDD2.n66 VDD2.n65 8.14595
R1762 VDD2.n149 VDD2.n77 7.3702
R1763 VDD2.n146 VDD2.n79 7.3702
R1764 VDD2.n103 VDD2.n101 7.3702
R1765 VDD2.n24 VDD2.n22 7.3702
R1766 VDD2.n69 VDD2.n2 7.3702
R1767 VDD2.n72 VDD2.n0 7.3702
R1768 VDD2.n147 VDD2.n77 6.59444
R1769 VDD2.n147 VDD2.n146 6.59444
R1770 VDD2.n70 VDD2.n69 6.59444
R1771 VDD2.n70 VDD2.n0 6.59444
R1772 VDD2.n143 VDD2.n79 5.81868
R1773 VDD2.n106 VDD2.n101 5.81868
R1774 VDD2.n27 VDD2.n22 5.81868
R1775 VDD2.n66 VDD2.n2 5.81868
R1776 VDD2.n142 VDD2.n81 5.04292
R1777 VDD2.n107 VDD2.n99 5.04292
R1778 VDD2.n28 VDD2.n20 5.04292
R1779 VDD2.n65 VDD2.n4 5.04292
R1780 VDD2.n139 VDD2.n138 4.26717
R1781 VDD2.n111 VDD2.n110 4.26717
R1782 VDD2.n32 VDD2.n31 4.26717
R1783 VDD2.n62 VDD2.n61 4.26717
R1784 VDD2.n135 VDD2.n83 3.49141
R1785 VDD2.n114 VDD2.n97 3.49141
R1786 VDD2.n35 VDD2.n18 3.49141
R1787 VDD2.n58 VDD2.n6 3.49141
R1788 VDD2.n102 VDD2.n100 2.84303
R1789 VDD2.n23 VDD2.n21 2.84303
R1790 VDD2.n134 VDD2.n85 2.71565
R1791 VDD2.n115 VDD2.n95 2.71565
R1792 VDD2.n36 VDD2.n16 2.71565
R1793 VDD2.n57 VDD2.n8 2.71565
R1794 VDD2.n131 VDD2.n130 1.93989
R1795 VDD2.n119 VDD2.n118 1.93989
R1796 VDD2.n41 VDD2.n39 1.93989
R1797 VDD2.n54 VDD2.n53 1.93989
R1798 VDD2.n153 VDD2.t8 1.45745
R1799 VDD2.n153 VDD2.t1 1.45745
R1800 VDD2.n151 VDD2.t7 1.45745
R1801 VDD2.n151 VDD2.t5 1.45745
R1802 VDD2.n75 VDD2.t2 1.45745
R1803 VDD2.n75 VDD2.t4 1.45745
R1804 VDD2.n73 VDD2.t9 1.45745
R1805 VDD2.n73 VDD2.t6 1.45745
R1806 VDD2.n152 VDD2.n150 1.42291
R1807 VDD2.n127 VDD2.n87 1.16414
R1808 VDD2.n122 VDD2.n92 1.16414
R1809 VDD2.n40 VDD2.n14 1.16414
R1810 VDD2.n50 VDD2.n10 1.16414
R1811 VDD2 VDD2.n152 0.414293
R1812 VDD2.n126 VDD2.n89 0.388379
R1813 VDD2.n123 VDD2.n91 0.388379
R1814 VDD2.n46 VDD2.n45 0.388379
R1815 VDD2.n49 VDD2.n12 0.388379
R1816 VDD2.n76 VDD2.n74 0.300757
R1817 VDD2.n148 VDD2.n78 0.155672
R1818 VDD2.n141 VDD2.n78 0.155672
R1819 VDD2.n141 VDD2.n140 0.155672
R1820 VDD2.n140 VDD2.n82 0.155672
R1821 VDD2.n133 VDD2.n82 0.155672
R1822 VDD2.n133 VDD2.n132 0.155672
R1823 VDD2.n132 VDD2.n86 0.155672
R1824 VDD2.n125 VDD2.n86 0.155672
R1825 VDD2.n125 VDD2.n124 0.155672
R1826 VDD2.n124 VDD2.n90 0.155672
R1827 VDD2.n117 VDD2.n90 0.155672
R1828 VDD2.n117 VDD2.n116 0.155672
R1829 VDD2.n116 VDD2.n96 0.155672
R1830 VDD2.n109 VDD2.n96 0.155672
R1831 VDD2.n109 VDD2.n108 0.155672
R1832 VDD2.n108 VDD2.n100 0.155672
R1833 VDD2.n29 VDD2.n21 0.155672
R1834 VDD2.n30 VDD2.n29 0.155672
R1835 VDD2.n30 VDD2.n17 0.155672
R1836 VDD2.n37 VDD2.n17 0.155672
R1837 VDD2.n38 VDD2.n37 0.155672
R1838 VDD2.n38 VDD2.n13 0.155672
R1839 VDD2.n47 VDD2.n13 0.155672
R1840 VDD2.n48 VDD2.n47 0.155672
R1841 VDD2.n48 VDD2.n9 0.155672
R1842 VDD2.n55 VDD2.n9 0.155672
R1843 VDD2.n56 VDD2.n55 0.155672
R1844 VDD2.n56 VDD2.n5 0.155672
R1845 VDD2.n63 VDD2.n5 0.155672
R1846 VDD2.n64 VDD2.n63 0.155672
R1847 VDD2.n64 VDD2.n1 0.155672
R1848 VDD2.n71 VDD2.n1 0.155672
R1849 VTAIL.n304 VTAIL.n236 289.615
R1850 VTAIL.n70 VTAIL.n2 289.615
R1851 VTAIL.n230 VTAIL.n162 289.615
R1852 VTAIL.n152 VTAIL.n84 289.615
R1853 VTAIL.n261 VTAIL.n260 185
R1854 VTAIL.n263 VTAIL.n262 185
R1855 VTAIL.n256 VTAIL.n255 185
R1856 VTAIL.n269 VTAIL.n268 185
R1857 VTAIL.n271 VTAIL.n270 185
R1858 VTAIL.n252 VTAIL.n251 185
R1859 VTAIL.n278 VTAIL.n277 185
R1860 VTAIL.n279 VTAIL.n250 185
R1861 VTAIL.n281 VTAIL.n280 185
R1862 VTAIL.n248 VTAIL.n247 185
R1863 VTAIL.n287 VTAIL.n286 185
R1864 VTAIL.n289 VTAIL.n288 185
R1865 VTAIL.n244 VTAIL.n243 185
R1866 VTAIL.n295 VTAIL.n294 185
R1867 VTAIL.n297 VTAIL.n296 185
R1868 VTAIL.n240 VTAIL.n239 185
R1869 VTAIL.n303 VTAIL.n302 185
R1870 VTAIL.n305 VTAIL.n304 185
R1871 VTAIL.n27 VTAIL.n26 185
R1872 VTAIL.n29 VTAIL.n28 185
R1873 VTAIL.n22 VTAIL.n21 185
R1874 VTAIL.n35 VTAIL.n34 185
R1875 VTAIL.n37 VTAIL.n36 185
R1876 VTAIL.n18 VTAIL.n17 185
R1877 VTAIL.n44 VTAIL.n43 185
R1878 VTAIL.n45 VTAIL.n16 185
R1879 VTAIL.n47 VTAIL.n46 185
R1880 VTAIL.n14 VTAIL.n13 185
R1881 VTAIL.n53 VTAIL.n52 185
R1882 VTAIL.n55 VTAIL.n54 185
R1883 VTAIL.n10 VTAIL.n9 185
R1884 VTAIL.n61 VTAIL.n60 185
R1885 VTAIL.n63 VTAIL.n62 185
R1886 VTAIL.n6 VTAIL.n5 185
R1887 VTAIL.n69 VTAIL.n68 185
R1888 VTAIL.n71 VTAIL.n70 185
R1889 VTAIL.n231 VTAIL.n230 185
R1890 VTAIL.n229 VTAIL.n228 185
R1891 VTAIL.n166 VTAIL.n165 185
R1892 VTAIL.n223 VTAIL.n222 185
R1893 VTAIL.n221 VTAIL.n220 185
R1894 VTAIL.n170 VTAIL.n169 185
R1895 VTAIL.n215 VTAIL.n214 185
R1896 VTAIL.n213 VTAIL.n212 185
R1897 VTAIL.n174 VTAIL.n173 185
R1898 VTAIL.n178 VTAIL.n176 185
R1899 VTAIL.n207 VTAIL.n206 185
R1900 VTAIL.n205 VTAIL.n204 185
R1901 VTAIL.n180 VTAIL.n179 185
R1902 VTAIL.n199 VTAIL.n198 185
R1903 VTAIL.n197 VTAIL.n196 185
R1904 VTAIL.n184 VTAIL.n183 185
R1905 VTAIL.n191 VTAIL.n190 185
R1906 VTAIL.n189 VTAIL.n188 185
R1907 VTAIL.n153 VTAIL.n152 185
R1908 VTAIL.n151 VTAIL.n150 185
R1909 VTAIL.n88 VTAIL.n87 185
R1910 VTAIL.n145 VTAIL.n144 185
R1911 VTAIL.n143 VTAIL.n142 185
R1912 VTAIL.n92 VTAIL.n91 185
R1913 VTAIL.n137 VTAIL.n136 185
R1914 VTAIL.n135 VTAIL.n134 185
R1915 VTAIL.n96 VTAIL.n95 185
R1916 VTAIL.n100 VTAIL.n98 185
R1917 VTAIL.n129 VTAIL.n128 185
R1918 VTAIL.n127 VTAIL.n126 185
R1919 VTAIL.n102 VTAIL.n101 185
R1920 VTAIL.n121 VTAIL.n120 185
R1921 VTAIL.n119 VTAIL.n118 185
R1922 VTAIL.n106 VTAIL.n105 185
R1923 VTAIL.n113 VTAIL.n112 185
R1924 VTAIL.n111 VTAIL.n110 185
R1925 VTAIL.n259 VTAIL.t13 149.524
R1926 VTAIL.n25 VTAIL.t8 149.524
R1927 VTAIL.n187 VTAIL.t2 149.524
R1928 VTAIL.n109 VTAIL.t12 149.524
R1929 VTAIL.n262 VTAIL.n261 104.615
R1930 VTAIL.n262 VTAIL.n255 104.615
R1931 VTAIL.n269 VTAIL.n255 104.615
R1932 VTAIL.n270 VTAIL.n269 104.615
R1933 VTAIL.n270 VTAIL.n251 104.615
R1934 VTAIL.n278 VTAIL.n251 104.615
R1935 VTAIL.n279 VTAIL.n278 104.615
R1936 VTAIL.n280 VTAIL.n279 104.615
R1937 VTAIL.n280 VTAIL.n247 104.615
R1938 VTAIL.n287 VTAIL.n247 104.615
R1939 VTAIL.n288 VTAIL.n287 104.615
R1940 VTAIL.n288 VTAIL.n243 104.615
R1941 VTAIL.n295 VTAIL.n243 104.615
R1942 VTAIL.n296 VTAIL.n295 104.615
R1943 VTAIL.n296 VTAIL.n239 104.615
R1944 VTAIL.n303 VTAIL.n239 104.615
R1945 VTAIL.n304 VTAIL.n303 104.615
R1946 VTAIL.n28 VTAIL.n27 104.615
R1947 VTAIL.n28 VTAIL.n21 104.615
R1948 VTAIL.n35 VTAIL.n21 104.615
R1949 VTAIL.n36 VTAIL.n35 104.615
R1950 VTAIL.n36 VTAIL.n17 104.615
R1951 VTAIL.n44 VTAIL.n17 104.615
R1952 VTAIL.n45 VTAIL.n44 104.615
R1953 VTAIL.n46 VTAIL.n45 104.615
R1954 VTAIL.n46 VTAIL.n13 104.615
R1955 VTAIL.n53 VTAIL.n13 104.615
R1956 VTAIL.n54 VTAIL.n53 104.615
R1957 VTAIL.n54 VTAIL.n9 104.615
R1958 VTAIL.n61 VTAIL.n9 104.615
R1959 VTAIL.n62 VTAIL.n61 104.615
R1960 VTAIL.n62 VTAIL.n5 104.615
R1961 VTAIL.n69 VTAIL.n5 104.615
R1962 VTAIL.n70 VTAIL.n69 104.615
R1963 VTAIL.n230 VTAIL.n229 104.615
R1964 VTAIL.n229 VTAIL.n165 104.615
R1965 VTAIL.n222 VTAIL.n165 104.615
R1966 VTAIL.n222 VTAIL.n221 104.615
R1967 VTAIL.n221 VTAIL.n169 104.615
R1968 VTAIL.n214 VTAIL.n169 104.615
R1969 VTAIL.n214 VTAIL.n213 104.615
R1970 VTAIL.n213 VTAIL.n173 104.615
R1971 VTAIL.n178 VTAIL.n173 104.615
R1972 VTAIL.n206 VTAIL.n178 104.615
R1973 VTAIL.n206 VTAIL.n205 104.615
R1974 VTAIL.n205 VTAIL.n179 104.615
R1975 VTAIL.n198 VTAIL.n179 104.615
R1976 VTAIL.n198 VTAIL.n197 104.615
R1977 VTAIL.n197 VTAIL.n183 104.615
R1978 VTAIL.n190 VTAIL.n183 104.615
R1979 VTAIL.n190 VTAIL.n189 104.615
R1980 VTAIL.n152 VTAIL.n151 104.615
R1981 VTAIL.n151 VTAIL.n87 104.615
R1982 VTAIL.n144 VTAIL.n87 104.615
R1983 VTAIL.n144 VTAIL.n143 104.615
R1984 VTAIL.n143 VTAIL.n91 104.615
R1985 VTAIL.n136 VTAIL.n91 104.615
R1986 VTAIL.n136 VTAIL.n135 104.615
R1987 VTAIL.n135 VTAIL.n95 104.615
R1988 VTAIL.n100 VTAIL.n95 104.615
R1989 VTAIL.n128 VTAIL.n100 104.615
R1990 VTAIL.n128 VTAIL.n127 104.615
R1991 VTAIL.n127 VTAIL.n101 104.615
R1992 VTAIL.n120 VTAIL.n101 104.615
R1993 VTAIL.n120 VTAIL.n119 104.615
R1994 VTAIL.n119 VTAIL.n105 104.615
R1995 VTAIL.n112 VTAIL.n105 104.615
R1996 VTAIL.n112 VTAIL.n111 104.615
R1997 VTAIL.n261 VTAIL.t13 52.3082
R1998 VTAIL.n27 VTAIL.t8 52.3082
R1999 VTAIL.n189 VTAIL.t2 52.3082
R2000 VTAIL.n111 VTAIL.t12 52.3082
R2001 VTAIL.n161 VTAIL.n160 45.4572
R2002 VTAIL.n159 VTAIL.n158 45.4572
R2003 VTAIL.n83 VTAIL.n82 45.4572
R2004 VTAIL.n81 VTAIL.n80 45.4572
R2005 VTAIL.n311 VTAIL.n310 45.457
R2006 VTAIL.n1 VTAIL.n0 45.457
R2007 VTAIL.n77 VTAIL.n76 45.457
R2008 VTAIL.n79 VTAIL.n78 45.457
R2009 VTAIL.n309 VTAIL.n308 32.7672
R2010 VTAIL.n75 VTAIL.n74 32.7672
R2011 VTAIL.n235 VTAIL.n234 32.7672
R2012 VTAIL.n157 VTAIL.n156 32.7672
R2013 VTAIL.n81 VTAIL.n79 26.9272
R2014 VTAIL.n309 VTAIL.n235 25.5048
R2015 VTAIL.n281 VTAIL.n248 13.1884
R2016 VTAIL.n47 VTAIL.n14 13.1884
R2017 VTAIL.n176 VTAIL.n174 13.1884
R2018 VTAIL.n98 VTAIL.n96 13.1884
R2019 VTAIL.n282 VTAIL.n250 12.8005
R2020 VTAIL.n286 VTAIL.n285 12.8005
R2021 VTAIL.n48 VTAIL.n16 12.8005
R2022 VTAIL.n52 VTAIL.n51 12.8005
R2023 VTAIL.n212 VTAIL.n211 12.8005
R2024 VTAIL.n208 VTAIL.n207 12.8005
R2025 VTAIL.n134 VTAIL.n133 12.8005
R2026 VTAIL.n130 VTAIL.n129 12.8005
R2027 VTAIL.n277 VTAIL.n276 12.0247
R2028 VTAIL.n289 VTAIL.n246 12.0247
R2029 VTAIL.n43 VTAIL.n42 12.0247
R2030 VTAIL.n55 VTAIL.n12 12.0247
R2031 VTAIL.n215 VTAIL.n172 12.0247
R2032 VTAIL.n204 VTAIL.n177 12.0247
R2033 VTAIL.n137 VTAIL.n94 12.0247
R2034 VTAIL.n126 VTAIL.n99 12.0247
R2035 VTAIL.n275 VTAIL.n252 11.249
R2036 VTAIL.n290 VTAIL.n244 11.249
R2037 VTAIL.n41 VTAIL.n18 11.249
R2038 VTAIL.n56 VTAIL.n10 11.249
R2039 VTAIL.n216 VTAIL.n170 11.249
R2040 VTAIL.n203 VTAIL.n180 11.249
R2041 VTAIL.n138 VTAIL.n92 11.249
R2042 VTAIL.n125 VTAIL.n102 11.249
R2043 VTAIL.n272 VTAIL.n271 10.4732
R2044 VTAIL.n294 VTAIL.n293 10.4732
R2045 VTAIL.n38 VTAIL.n37 10.4732
R2046 VTAIL.n60 VTAIL.n59 10.4732
R2047 VTAIL.n220 VTAIL.n219 10.4732
R2048 VTAIL.n200 VTAIL.n199 10.4732
R2049 VTAIL.n142 VTAIL.n141 10.4732
R2050 VTAIL.n122 VTAIL.n121 10.4732
R2051 VTAIL.n260 VTAIL.n259 10.2747
R2052 VTAIL.n26 VTAIL.n25 10.2747
R2053 VTAIL.n188 VTAIL.n187 10.2747
R2054 VTAIL.n110 VTAIL.n109 10.2747
R2055 VTAIL.n268 VTAIL.n254 9.69747
R2056 VTAIL.n297 VTAIL.n242 9.69747
R2057 VTAIL.n34 VTAIL.n20 9.69747
R2058 VTAIL.n63 VTAIL.n8 9.69747
R2059 VTAIL.n223 VTAIL.n168 9.69747
R2060 VTAIL.n196 VTAIL.n182 9.69747
R2061 VTAIL.n145 VTAIL.n90 9.69747
R2062 VTAIL.n118 VTAIL.n104 9.69747
R2063 VTAIL.n308 VTAIL.n307 9.45567
R2064 VTAIL.n74 VTAIL.n73 9.45567
R2065 VTAIL.n234 VTAIL.n233 9.45567
R2066 VTAIL.n156 VTAIL.n155 9.45567
R2067 VTAIL.n307 VTAIL.n306 9.3005
R2068 VTAIL.n301 VTAIL.n300 9.3005
R2069 VTAIL.n299 VTAIL.n298 9.3005
R2070 VTAIL.n242 VTAIL.n241 9.3005
R2071 VTAIL.n293 VTAIL.n292 9.3005
R2072 VTAIL.n291 VTAIL.n290 9.3005
R2073 VTAIL.n246 VTAIL.n245 9.3005
R2074 VTAIL.n285 VTAIL.n284 9.3005
R2075 VTAIL.n258 VTAIL.n257 9.3005
R2076 VTAIL.n265 VTAIL.n264 9.3005
R2077 VTAIL.n267 VTAIL.n266 9.3005
R2078 VTAIL.n254 VTAIL.n253 9.3005
R2079 VTAIL.n273 VTAIL.n272 9.3005
R2080 VTAIL.n275 VTAIL.n274 9.3005
R2081 VTAIL.n276 VTAIL.n249 9.3005
R2082 VTAIL.n283 VTAIL.n282 9.3005
R2083 VTAIL.n238 VTAIL.n237 9.3005
R2084 VTAIL.n73 VTAIL.n72 9.3005
R2085 VTAIL.n67 VTAIL.n66 9.3005
R2086 VTAIL.n65 VTAIL.n64 9.3005
R2087 VTAIL.n8 VTAIL.n7 9.3005
R2088 VTAIL.n59 VTAIL.n58 9.3005
R2089 VTAIL.n57 VTAIL.n56 9.3005
R2090 VTAIL.n12 VTAIL.n11 9.3005
R2091 VTAIL.n51 VTAIL.n50 9.3005
R2092 VTAIL.n24 VTAIL.n23 9.3005
R2093 VTAIL.n31 VTAIL.n30 9.3005
R2094 VTAIL.n33 VTAIL.n32 9.3005
R2095 VTAIL.n20 VTAIL.n19 9.3005
R2096 VTAIL.n39 VTAIL.n38 9.3005
R2097 VTAIL.n41 VTAIL.n40 9.3005
R2098 VTAIL.n42 VTAIL.n15 9.3005
R2099 VTAIL.n49 VTAIL.n48 9.3005
R2100 VTAIL.n4 VTAIL.n3 9.3005
R2101 VTAIL.n186 VTAIL.n185 9.3005
R2102 VTAIL.n193 VTAIL.n192 9.3005
R2103 VTAIL.n195 VTAIL.n194 9.3005
R2104 VTAIL.n182 VTAIL.n181 9.3005
R2105 VTAIL.n201 VTAIL.n200 9.3005
R2106 VTAIL.n203 VTAIL.n202 9.3005
R2107 VTAIL.n177 VTAIL.n175 9.3005
R2108 VTAIL.n209 VTAIL.n208 9.3005
R2109 VTAIL.n233 VTAIL.n232 9.3005
R2110 VTAIL.n164 VTAIL.n163 9.3005
R2111 VTAIL.n227 VTAIL.n226 9.3005
R2112 VTAIL.n225 VTAIL.n224 9.3005
R2113 VTAIL.n168 VTAIL.n167 9.3005
R2114 VTAIL.n219 VTAIL.n218 9.3005
R2115 VTAIL.n217 VTAIL.n216 9.3005
R2116 VTAIL.n172 VTAIL.n171 9.3005
R2117 VTAIL.n211 VTAIL.n210 9.3005
R2118 VTAIL.n108 VTAIL.n107 9.3005
R2119 VTAIL.n115 VTAIL.n114 9.3005
R2120 VTAIL.n117 VTAIL.n116 9.3005
R2121 VTAIL.n104 VTAIL.n103 9.3005
R2122 VTAIL.n123 VTAIL.n122 9.3005
R2123 VTAIL.n125 VTAIL.n124 9.3005
R2124 VTAIL.n99 VTAIL.n97 9.3005
R2125 VTAIL.n131 VTAIL.n130 9.3005
R2126 VTAIL.n155 VTAIL.n154 9.3005
R2127 VTAIL.n86 VTAIL.n85 9.3005
R2128 VTAIL.n149 VTAIL.n148 9.3005
R2129 VTAIL.n147 VTAIL.n146 9.3005
R2130 VTAIL.n90 VTAIL.n89 9.3005
R2131 VTAIL.n141 VTAIL.n140 9.3005
R2132 VTAIL.n139 VTAIL.n138 9.3005
R2133 VTAIL.n94 VTAIL.n93 9.3005
R2134 VTAIL.n133 VTAIL.n132 9.3005
R2135 VTAIL.n267 VTAIL.n256 8.92171
R2136 VTAIL.n298 VTAIL.n240 8.92171
R2137 VTAIL.n33 VTAIL.n22 8.92171
R2138 VTAIL.n64 VTAIL.n6 8.92171
R2139 VTAIL.n224 VTAIL.n166 8.92171
R2140 VTAIL.n195 VTAIL.n184 8.92171
R2141 VTAIL.n146 VTAIL.n88 8.92171
R2142 VTAIL.n117 VTAIL.n106 8.92171
R2143 VTAIL.n264 VTAIL.n263 8.14595
R2144 VTAIL.n302 VTAIL.n301 8.14595
R2145 VTAIL.n30 VTAIL.n29 8.14595
R2146 VTAIL.n68 VTAIL.n67 8.14595
R2147 VTAIL.n228 VTAIL.n227 8.14595
R2148 VTAIL.n192 VTAIL.n191 8.14595
R2149 VTAIL.n150 VTAIL.n149 8.14595
R2150 VTAIL.n114 VTAIL.n113 8.14595
R2151 VTAIL.n260 VTAIL.n258 7.3702
R2152 VTAIL.n305 VTAIL.n238 7.3702
R2153 VTAIL.n308 VTAIL.n236 7.3702
R2154 VTAIL.n26 VTAIL.n24 7.3702
R2155 VTAIL.n71 VTAIL.n4 7.3702
R2156 VTAIL.n74 VTAIL.n2 7.3702
R2157 VTAIL.n234 VTAIL.n162 7.3702
R2158 VTAIL.n231 VTAIL.n164 7.3702
R2159 VTAIL.n188 VTAIL.n186 7.3702
R2160 VTAIL.n156 VTAIL.n84 7.3702
R2161 VTAIL.n153 VTAIL.n86 7.3702
R2162 VTAIL.n110 VTAIL.n108 7.3702
R2163 VTAIL.n306 VTAIL.n305 6.59444
R2164 VTAIL.n306 VTAIL.n236 6.59444
R2165 VTAIL.n72 VTAIL.n71 6.59444
R2166 VTAIL.n72 VTAIL.n2 6.59444
R2167 VTAIL.n232 VTAIL.n162 6.59444
R2168 VTAIL.n232 VTAIL.n231 6.59444
R2169 VTAIL.n154 VTAIL.n84 6.59444
R2170 VTAIL.n154 VTAIL.n153 6.59444
R2171 VTAIL.n263 VTAIL.n258 5.81868
R2172 VTAIL.n302 VTAIL.n238 5.81868
R2173 VTAIL.n29 VTAIL.n24 5.81868
R2174 VTAIL.n68 VTAIL.n4 5.81868
R2175 VTAIL.n228 VTAIL.n164 5.81868
R2176 VTAIL.n191 VTAIL.n186 5.81868
R2177 VTAIL.n150 VTAIL.n86 5.81868
R2178 VTAIL.n113 VTAIL.n108 5.81868
R2179 VTAIL.n264 VTAIL.n256 5.04292
R2180 VTAIL.n301 VTAIL.n240 5.04292
R2181 VTAIL.n30 VTAIL.n22 5.04292
R2182 VTAIL.n67 VTAIL.n6 5.04292
R2183 VTAIL.n227 VTAIL.n166 5.04292
R2184 VTAIL.n192 VTAIL.n184 5.04292
R2185 VTAIL.n149 VTAIL.n88 5.04292
R2186 VTAIL.n114 VTAIL.n106 5.04292
R2187 VTAIL.n268 VTAIL.n267 4.26717
R2188 VTAIL.n298 VTAIL.n297 4.26717
R2189 VTAIL.n34 VTAIL.n33 4.26717
R2190 VTAIL.n64 VTAIL.n63 4.26717
R2191 VTAIL.n224 VTAIL.n223 4.26717
R2192 VTAIL.n196 VTAIL.n195 4.26717
R2193 VTAIL.n146 VTAIL.n145 4.26717
R2194 VTAIL.n118 VTAIL.n117 4.26717
R2195 VTAIL.n271 VTAIL.n254 3.49141
R2196 VTAIL.n294 VTAIL.n242 3.49141
R2197 VTAIL.n37 VTAIL.n20 3.49141
R2198 VTAIL.n60 VTAIL.n8 3.49141
R2199 VTAIL.n220 VTAIL.n168 3.49141
R2200 VTAIL.n199 VTAIL.n182 3.49141
R2201 VTAIL.n142 VTAIL.n90 3.49141
R2202 VTAIL.n121 VTAIL.n104 3.49141
R2203 VTAIL.n259 VTAIL.n257 2.84303
R2204 VTAIL.n25 VTAIL.n23 2.84303
R2205 VTAIL.n187 VTAIL.n185 2.84303
R2206 VTAIL.n109 VTAIL.n107 2.84303
R2207 VTAIL.n272 VTAIL.n252 2.71565
R2208 VTAIL.n293 VTAIL.n244 2.71565
R2209 VTAIL.n38 VTAIL.n18 2.71565
R2210 VTAIL.n59 VTAIL.n10 2.71565
R2211 VTAIL.n219 VTAIL.n170 2.71565
R2212 VTAIL.n200 VTAIL.n180 2.71565
R2213 VTAIL.n141 VTAIL.n92 2.71565
R2214 VTAIL.n122 VTAIL.n102 2.71565
R2215 VTAIL.n277 VTAIL.n275 1.93989
R2216 VTAIL.n290 VTAIL.n289 1.93989
R2217 VTAIL.n43 VTAIL.n41 1.93989
R2218 VTAIL.n56 VTAIL.n55 1.93989
R2219 VTAIL.n216 VTAIL.n215 1.93989
R2220 VTAIL.n204 VTAIL.n203 1.93989
R2221 VTAIL.n138 VTAIL.n137 1.93989
R2222 VTAIL.n126 VTAIL.n125 1.93989
R2223 VTAIL.n310 VTAIL.t18 1.45745
R2224 VTAIL.n310 VTAIL.t19 1.45745
R2225 VTAIL.n0 VTAIL.t16 1.45745
R2226 VTAIL.n0 VTAIL.t17 1.45745
R2227 VTAIL.n76 VTAIL.t1 1.45745
R2228 VTAIL.n76 VTAIL.t0 1.45745
R2229 VTAIL.n78 VTAIL.t5 1.45745
R2230 VTAIL.n78 VTAIL.t6 1.45745
R2231 VTAIL.n160 VTAIL.t7 1.45745
R2232 VTAIL.n160 VTAIL.t9 1.45745
R2233 VTAIL.n158 VTAIL.t4 1.45745
R2234 VTAIL.n158 VTAIL.t3 1.45745
R2235 VTAIL.n82 VTAIL.t14 1.45745
R2236 VTAIL.n82 VTAIL.t11 1.45745
R2237 VTAIL.n80 VTAIL.t15 1.45745
R2238 VTAIL.n80 VTAIL.t10 1.45745
R2239 VTAIL.n83 VTAIL.n81 1.42291
R2240 VTAIL.n157 VTAIL.n83 1.42291
R2241 VTAIL.n161 VTAIL.n159 1.42291
R2242 VTAIL.n235 VTAIL.n161 1.42291
R2243 VTAIL.n79 VTAIL.n77 1.42291
R2244 VTAIL.n77 VTAIL.n75 1.42291
R2245 VTAIL.n311 VTAIL.n309 1.42291
R2246 VTAIL.n159 VTAIL.n157 1.18153
R2247 VTAIL.n75 VTAIL.n1 1.18153
R2248 VTAIL.n276 VTAIL.n250 1.16414
R2249 VTAIL.n286 VTAIL.n246 1.16414
R2250 VTAIL.n42 VTAIL.n16 1.16414
R2251 VTAIL.n52 VTAIL.n12 1.16414
R2252 VTAIL.n212 VTAIL.n172 1.16414
R2253 VTAIL.n207 VTAIL.n177 1.16414
R2254 VTAIL.n134 VTAIL.n94 1.16414
R2255 VTAIL.n129 VTAIL.n99 1.16414
R2256 VTAIL VTAIL.n1 1.1255
R2257 VTAIL.n282 VTAIL.n281 0.388379
R2258 VTAIL.n285 VTAIL.n248 0.388379
R2259 VTAIL.n48 VTAIL.n47 0.388379
R2260 VTAIL.n51 VTAIL.n14 0.388379
R2261 VTAIL.n211 VTAIL.n174 0.388379
R2262 VTAIL.n208 VTAIL.n176 0.388379
R2263 VTAIL.n133 VTAIL.n96 0.388379
R2264 VTAIL.n130 VTAIL.n98 0.388379
R2265 VTAIL VTAIL.n311 0.297914
R2266 VTAIL.n265 VTAIL.n257 0.155672
R2267 VTAIL.n266 VTAIL.n265 0.155672
R2268 VTAIL.n266 VTAIL.n253 0.155672
R2269 VTAIL.n273 VTAIL.n253 0.155672
R2270 VTAIL.n274 VTAIL.n273 0.155672
R2271 VTAIL.n274 VTAIL.n249 0.155672
R2272 VTAIL.n283 VTAIL.n249 0.155672
R2273 VTAIL.n284 VTAIL.n283 0.155672
R2274 VTAIL.n284 VTAIL.n245 0.155672
R2275 VTAIL.n291 VTAIL.n245 0.155672
R2276 VTAIL.n292 VTAIL.n291 0.155672
R2277 VTAIL.n292 VTAIL.n241 0.155672
R2278 VTAIL.n299 VTAIL.n241 0.155672
R2279 VTAIL.n300 VTAIL.n299 0.155672
R2280 VTAIL.n300 VTAIL.n237 0.155672
R2281 VTAIL.n307 VTAIL.n237 0.155672
R2282 VTAIL.n31 VTAIL.n23 0.155672
R2283 VTAIL.n32 VTAIL.n31 0.155672
R2284 VTAIL.n32 VTAIL.n19 0.155672
R2285 VTAIL.n39 VTAIL.n19 0.155672
R2286 VTAIL.n40 VTAIL.n39 0.155672
R2287 VTAIL.n40 VTAIL.n15 0.155672
R2288 VTAIL.n49 VTAIL.n15 0.155672
R2289 VTAIL.n50 VTAIL.n49 0.155672
R2290 VTAIL.n50 VTAIL.n11 0.155672
R2291 VTAIL.n57 VTAIL.n11 0.155672
R2292 VTAIL.n58 VTAIL.n57 0.155672
R2293 VTAIL.n58 VTAIL.n7 0.155672
R2294 VTAIL.n65 VTAIL.n7 0.155672
R2295 VTAIL.n66 VTAIL.n65 0.155672
R2296 VTAIL.n66 VTAIL.n3 0.155672
R2297 VTAIL.n73 VTAIL.n3 0.155672
R2298 VTAIL.n233 VTAIL.n163 0.155672
R2299 VTAIL.n226 VTAIL.n163 0.155672
R2300 VTAIL.n226 VTAIL.n225 0.155672
R2301 VTAIL.n225 VTAIL.n167 0.155672
R2302 VTAIL.n218 VTAIL.n167 0.155672
R2303 VTAIL.n218 VTAIL.n217 0.155672
R2304 VTAIL.n217 VTAIL.n171 0.155672
R2305 VTAIL.n210 VTAIL.n171 0.155672
R2306 VTAIL.n210 VTAIL.n209 0.155672
R2307 VTAIL.n209 VTAIL.n175 0.155672
R2308 VTAIL.n202 VTAIL.n175 0.155672
R2309 VTAIL.n202 VTAIL.n201 0.155672
R2310 VTAIL.n201 VTAIL.n181 0.155672
R2311 VTAIL.n194 VTAIL.n181 0.155672
R2312 VTAIL.n194 VTAIL.n193 0.155672
R2313 VTAIL.n193 VTAIL.n185 0.155672
R2314 VTAIL.n155 VTAIL.n85 0.155672
R2315 VTAIL.n148 VTAIL.n85 0.155672
R2316 VTAIL.n148 VTAIL.n147 0.155672
R2317 VTAIL.n147 VTAIL.n89 0.155672
R2318 VTAIL.n140 VTAIL.n89 0.155672
R2319 VTAIL.n140 VTAIL.n139 0.155672
R2320 VTAIL.n139 VTAIL.n93 0.155672
R2321 VTAIL.n132 VTAIL.n93 0.155672
R2322 VTAIL.n132 VTAIL.n131 0.155672
R2323 VTAIL.n131 VTAIL.n97 0.155672
R2324 VTAIL.n124 VTAIL.n97 0.155672
R2325 VTAIL.n124 VTAIL.n123 0.155672
R2326 VTAIL.n123 VTAIL.n103 0.155672
R2327 VTAIL.n116 VTAIL.n103 0.155672
R2328 VTAIL.n116 VTAIL.n115 0.155672
R2329 VTAIL.n115 VTAIL.n107 0.155672
R2330 VP.n14 VP.t1 279.103
R2331 VP.n3 VP.t7 248.12
R2332 VP.n7 VP.t5 248.12
R2333 VP.n5 VP.t4 248.12
R2334 VP.n48 VP.t3 248.12
R2335 VP.n55 VP.t2 248.12
R2336 VP.n11 VP.t9 248.12
R2337 VP.n31 VP.t8 248.12
R2338 VP.n24 VP.t0 248.12
R2339 VP.n13 VP.t6 248.12
R2340 VP.n33 VP.n7 171.088
R2341 VP.n56 VP.n55 171.088
R2342 VP.n32 VP.n31 171.088
R2343 VP.n16 VP.n15 161.3
R2344 VP.n17 VP.n12 161.3
R2345 VP.n19 VP.n18 161.3
R2346 VP.n20 VP.n11 161.3
R2347 VP.n22 VP.n21 161.3
R2348 VP.n23 VP.n10 161.3
R2349 VP.n26 VP.n25 161.3
R2350 VP.n27 VP.n9 161.3
R2351 VP.n29 VP.n28 161.3
R2352 VP.n30 VP.n8 161.3
R2353 VP.n54 VP.n0 161.3
R2354 VP.n53 VP.n52 161.3
R2355 VP.n51 VP.n1 161.3
R2356 VP.n50 VP.n49 161.3
R2357 VP.n47 VP.n2 161.3
R2358 VP.n46 VP.n45 161.3
R2359 VP.n44 VP.n3 161.3
R2360 VP.n43 VP.n42 161.3
R2361 VP.n41 VP.n4 161.3
R2362 VP.n40 VP.n39 161.3
R2363 VP.n38 VP.n37 161.3
R2364 VP.n36 VP.n6 161.3
R2365 VP.n35 VP.n34 161.3
R2366 VP.n14 VP.n13 57.1957
R2367 VP.n42 VP.n41 56.5193
R2368 VP.n47 VP.n46 56.5193
R2369 VP.n23 VP.n22 56.5193
R2370 VP.n18 VP.n17 56.5193
R2371 VP.n33 VP.n32 47.3149
R2372 VP.n37 VP.n36 42.9216
R2373 VP.n53 VP.n1 42.9216
R2374 VP.n29 VP.n9 42.9216
R2375 VP.n36 VP.n35 38.0652
R2376 VP.n54 VP.n53 38.0652
R2377 VP.n30 VP.n29 38.0652
R2378 VP.n15 VP.n14 26.7159
R2379 VP.n41 VP.n40 24.4675
R2380 VP.n42 VP.n3 24.4675
R2381 VP.n46 VP.n3 24.4675
R2382 VP.n49 VP.n47 24.4675
R2383 VP.n25 VP.n23 24.4675
R2384 VP.n18 VP.n11 24.4675
R2385 VP.n22 VP.n11 24.4675
R2386 VP.n17 VP.n16 24.4675
R2387 VP.n37 VP.n5 17.1274
R2388 VP.n48 VP.n1 17.1274
R2389 VP.n24 VP.n9 17.1274
R2390 VP.n35 VP.n7 14.6807
R2391 VP.n55 VP.n54 14.6807
R2392 VP.n31 VP.n30 14.6807
R2393 VP.n40 VP.n5 7.3406
R2394 VP.n49 VP.n48 7.3406
R2395 VP.n25 VP.n24 7.3406
R2396 VP.n16 VP.n13 7.3406
R2397 VP.n15 VP.n12 0.189894
R2398 VP.n19 VP.n12 0.189894
R2399 VP.n20 VP.n19 0.189894
R2400 VP.n21 VP.n20 0.189894
R2401 VP.n21 VP.n10 0.189894
R2402 VP.n26 VP.n10 0.189894
R2403 VP.n27 VP.n26 0.189894
R2404 VP.n28 VP.n27 0.189894
R2405 VP.n28 VP.n8 0.189894
R2406 VP.n32 VP.n8 0.189894
R2407 VP.n34 VP.n33 0.189894
R2408 VP.n34 VP.n6 0.189894
R2409 VP.n38 VP.n6 0.189894
R2410 VP.n39 VP.n38 0.189894
R2411 VP.n39 VP.n4 0.189894
R2412 VP.n43 VP.n4 0.189894
R2413 VP.n44 VP.n43 0.189894
R2414 VP.n45 VP.n44 0.189894
R2415 VP.n45 VP.n2 0.189894
R2416 VP.n50 VP.n2 0.189894
R2417 VP.n51 VP.n50 0.189894
R2418 VP.n52 VP.n51 0.189894
R2419 VP.n52 VP.n0 0.189894
R2420 VP.n56 VP.n0 0.189894
R2421 VP VP.n56 0.0516364
R2422 VDD1.n68 VDD1.n0 289.615
R2423 VDD1.n143 VDD1.n75 289.615
R2424 VDD1.n69 VDD1.n68 185
R2425 VDD1.n67 VDD1.n66 185
R2426 VDD1.n4 VDD1.n3 185
R2427 VDD1.n61 VDD1.n60 185
R2428 VDD1.n59 VDD1.n58 185
R2429 VDD1.n8 VDD1.n7 185
R2430 VDD1.n53 VDD1.n52 185
R2431 VDD1.n51 VDD1.n50 185
R2432 VDD1.n12 VDD1.n11 185
R2433 VDD1.n16 VDD1.n14 185
R2434 VDD1.n45 VDD1.n44 185
R2435 VDD1.n43 VDD1.n42 185
R2436 VDD1.n18 VDD1.n17 185
R2437 VDD1.n37 VDD1.n36 185
R2438 VDD1.n35 VDD1.n34 185
R2439 VDD1.n22 VDD1.n21 185
R2440 VDD1.n29 VDD1.n28 185
R2441 VDD1.n27 VDD1.n26 185
R2442 VDD1.n100 VDD1.n99 185
R2443 VDD1.n102 VDD1.n101 185
R2444 VDD1.n95 VDD1.n94 185
R2445 VDD1.n108 VDD1.n107 185
R2446 VDD1.n110 VDD1.n109 185
R2447 VDD1.n91 VDD1.n90 185
R2448 VDD1.n117 VDD1.n116 185
R2449 VDD1.n118 VDD1.n89 185
R2450 VDD1.n120 VDD1.n119 185
R2451 VDD1.n87 VDD1.n86 185
R2452 VDD1.n126 VDD1.n125 185
R2453 VDD1.n128 VDD1.n127 185
R2454 VDD1.n83 VDD1.n82 185
R2455 VDD1.n134 VDD1.n133 185
R2456 VDD1.n136 VDD1.n135 185
R2457 VDD1.n79 VDD1.n78 185
R2458 VDD1.n142 VDD1.n141 185
R2459 VDD1.n144 VDD1.n143 185
R2460 VDD1.n25 VDD1.t8 149.524
R2461 VDD1.n98 VDD1.t4 149.524
R2462 VDD1.n68 VDD1.n67 104.615
R2463 VDD1.n67 VDD1.n3 104.615
R2464 VDD1.n60 VDD1.n3 104.615
R2465 VDD1.n60 VDD1.n59 104.615
R2466 VDD1.n59 VDD1.n7 104.615
R2467 VDD1.n52 VDD1.n7 104.615
R2468 VDD1.n52 VDD1.n51 104.615
R2469 VDD1.n51 VDD1.n11 104.615
R2470 VDD1.n16 VDD1.n11 104.615
R2471 VDD1.n44 VDD1.n16 104.615
R2472 VDD1.n44 VDD1.n43 104.615
R2473 VDD1.n43 VDD1.n17 104.615
R2474 VDD1.n36 VDD1.n17 104.615
R2475 VDD1.n36 VDD1.n35 104.615
R2476 VDD1.n35 VDD1.n21 104.615
R2477 VDD1.n28 VDD1.n21 104.615
R2478 VDD1.n28 VDD1.n27 104.615
R2479 VDD1.n101 VDD1.n100 104.615
R2480 VDD1.n101 VDD1.n94 104.615
R2481 VDD1.n108 VDD1.n94 104.615
R2482 VDD1.n109 VDD1.n108 104.615
R2483 VDD1.n109 VDD1.n90 104.615
R2484 VDD1.n117 VDD1.n90 104.615
R2485 VDD1.n118 VDD1.n117 104.615
R2486 VDD1.n119 VDD1.n118 104.615
R2487 VDD1.n119 VDD1.n86 104.615
R2488 VDD1.n126 VDD1.n86 104.615
R2489 VDD1.n127 VDD1.n126 104.615
R2490 VDD1.n127 VDD1.n82 104.615
R2491 VDD1.n134 VDD1.n82 104.615
R2492 VDD1.n135 VDD1.n134 104.615
R2493 VDD1.n135 VDD1.n78 104.615
R2494 VDD1.n142 VDD1.n78 104.615
R2495 VDD1.n143 VDD1.n142 104.615
R2496 VDD1.n151 VDD1.n150 63.1473
R2497 VDD1.n74 VDD1.n73 62.136
R2498 VDD1.n153 VDD1.n152 62.1358
R2499 VDD1.n149 VDD1.n148 62.1358
R2500 VDD1.n27 VDD1.t8 52.3082
R2501 VDD1.n100 VDD1.t4 52.3082
R2502 VDD1.n74 VDD1.n72 50.8684
R2503 VDD1.n149 VDD1.n147 50.8684
R2504 VDD1.n153 VDD1.n151 43.4815
R2505 VDD1.n14 VDD1.n12 13.1884
R2506 VDD1.n120 VDD1.n87 13.1884
R2507 VDD1.n50 VDD1.n49 12.8005
R2508 VDD1.n46 VDD1.n45 12.8005
R2509 VDD1.n121 VDD1.n89 12.8005
R2510 VDD1.n125 VDD1.n124 12.8005
R2511 VDD1.n53 VDD1.n10 12.0247
R2512 VDD1.n42 VDD1.n15 12.0247
R2513 VDD1.n116 VDD1.n115 12.0247
R2514 VDD1.n128 VDD1.n85 12.0247
R2515 VDD1.n54 VDD1.n8 11.249
R2516 VDD1.n41 VDD1.n18 11.249
R2517 VDD1.n114 VDD1.n91 11.249
R2518 VDD1.n129 VDD1.n83 11.249
R2519 VDD1.n58 VDD1.n57 10.4732
R2520 VDD1.n38 VDD1.n37 10.4732
R2521 VDD1.n111 VDD1.n110 10.4732
R2522 VDD1.n133 VDD1.n132 10.4732
R2523 VDD1.n26 VDD1.n25 10.2747
R2524 VDD1.n99 VDD1.n98 10.2747
R2525 VDD1.n61 VDD1.n6 9.69747
R2526 VDD1.n34 VDD1.n20 9.69747
R2527 VDD1.n107 VDD1.n93 9.69747
R2528 VDD1.n136 VDD1.n81 9.69747
R2529 VDD1.n72 VDD1.n71 9.45567
R2530 VDD1.n147 VDD1.n146 9.45567
R2531 VDD1.n24 VDD1.n23 9.3005
R2532 VDD1.n31 VDD1.n30 9.3005
R2533 VDD1.n33 VDD1.n32 9.3005
R2534 VDD1.n20 VDD1.n19 9.3005
R2535 VDD1.n39 VDD1.n38 9.3005
R2536 VDD1.n41 VDD1.n40 9.3005
R2537 VDD1.n15 VDD1.n13 9.3005
R2538 VDD1.n47 VDD1.n46 9.3005
R2539 VDD1.n71 VDD1.n70 9.3005
R2540 VDD1.n2 VDD1.n1 9.3005
R2541 VDD1.n65 VDD1.n64 9.3005
R2542 VDD1.n63 VDD1.n62 9.3005
R2543 VDD1.n6 VDD1.n5 9.3005
R2544 VDD1.n57 VDD1.n56 9.3005
R2545 VDD1.n55 VDD1.n54 9.3005
R2546 VDD1.n10 VDD1.n9 9.3005
R2547 VDD1.n49 VDD1.n48 9.3005
R2548 VDD1.n146 VDD1.n145 9.3005
R2549 VDD1.n140 VDD1.n139 9.3005
R2550 VDD1.n138 VDD1.n137 9.3005
R2551 VDD1.n81 VDD1.n80 9.3005
R2552 VDD1.n132 VDD1.n131 9.3005
R2553 VDD1.n130 VDD1.n129 9.3005
R2554 VDD1.n85 VDD1.n84 9.3005
R2555 VDD1.n124 VDD1.n123 9.3005
R2556 VDD1.n97 VDD1.n96 9.3005
R2557 VDD1.n104 VDD1.n103 9.3005
R2558 VDD1.n106 VDD1.n105 9.3005
R2559 VDD1.n93 VDD1.n92 9.3005
R2560 VDD1.n112 VDD1.n111 9.3005
R2561 VDD1.n114 VDD1.n113 9.3005
R2562 VDD1.n115 VDD1.n88 9.3005
R2563 VDD1.n122 VDD1.n121 9.3005
R2564 VDD1.n77 VDD1.n76 9.3005
R2565 VDD1.n62 VDD1.n4 8.92171
R2566 VDD1.n33 VDD1.n22 8.92171
R2567 VDD1.n106 VDD1.n95 8.92171
R2568 VDD1.n137 VDD1.n79 8.92171
R2569 VDD1.n66 VDD1.n65 8.14595
R2570 VDD1.n30 VDD1.n29 8.14595
R2571 VDD1.n103 VDD1.n102 8.14595
R2572 VDD1.n141 VDD1.n140 8.14595
R2573 VDD1.n72 VDD1.n0 7.3702
R2574 VDD1.n69 VDD1.n2 7.3702
R2575 VDD1.n26 VDD1.n24 7.3702
R2576 VDD1.n99 VDD1.n97 7.3702
R2577 VDD1.n144 VDD1.n77 7.3702
R2578 VDD1.n147 VDD1.n75 7.3702
R2579 VDD1.n70 VDD1.n0 6.59444
R2580 VDD1.n70 VDD1.n69 6.59444
R2581 VDD1.n145 VDD1.n144 6.59444
R2582 VDD1.n145 VDD1.n75 6.59444
R2583 VDD1.n66 VDD1.n2 5.81868
R2584 VDD1.n29 VDD1.n24 5.81868
R2585 VDD1.n102 VDD1.n97 5.81868
R2586 VDD1.n141 VDD1.n77 5.81868
R2587 VDD1.n65 VDD1.n4 5.04292
R2588 VDD1.n30 VDD1.n22 5.04292
R2589 VDD1.n103 VDD1.n95 5.04292
R2590 VDD1.n140 VDD1.n79 5.04292
R2591 VDD1.n62 VDD1.n61 4.26717
R2592 VDD1.n34 VDD1.n33 4.26717
R2593 VDD1.n107 VDD1.n106 4.26717
R2594 VDD1.n137 VDD1.n136 4.26717
R2595 VDD1.n58 VDD1.n6 3.49141
R2596 VDD1.n37 VDD1.n20 3.49141
R2597 VDD1.n110 VDD1.n93 3.49141
R2598 VDD1.n133 VDD1.n81 3.49141
R2599 VDD1.n25 VDD1.n23 2.84303
R2600 VDD1.n98 VDD1.n96 2.84303
R2601 VDD1.n57 VDD1.n8 2.71565
R2602 VDD1.n38 VDD1.n18 2.71565
R2603 VDD1.n111 VDD1.n91 2.71565
R2604 VDD1.n132 VDD1.n83 2.71565
R2605 VDD1.n54 VDD1.n53 1.93989
R2606 VDD1.n42 VDD1.n41 1.93989
R2607 VDD1.n116 VDD1.n114 1.93989
R2608 VDD1.n129 VDD1.n128 1.93989
R2609 VDD1.n152 VDD1.t9 1.45745
R2610 VDD1.n152 VDD1.t1 1.45745
R2611 VDD1.n73 VDD1.t3 1.45745
R2612 VDD1.n73 VDD1.t0 1.45745
R2613 VDD1.n150 VDD1.t6 1.45745
R2614 VDD1.n150 VDD1.t7 1.45745
R2615 VDD1.n148 VDD1.t5 1.45745
R2616 VDD1.n148 VDD1.t2 1.45745
R2617 VDD1.n50 VDD1.n10 1.16414
R2618 VDD1.n45 VDD1.n15 1.16414
R2619 VDD1.n115 VDD1.n89 1.16414
R2620 VDD1.n125 VDD1.n85 1.16414
R2621 VDD1 VDD1.n153 1.00912
R2622 VDD1 VDD1.n74 0.414293
R2623 VDD1.n49 VDD1.n12 0.388379
R2624 VDD1.n46 VDD1.n14 0.388379
R2625 VDD1.n121 VDD1.n120 0.388379
R2626 VDD1.n124 VDD1.n87 0.388379
R2627 VDD1.n151 VDD1.n149 0.300757
R2628 VDD1.n71 VDD1.n1 0.155672
R2629 VDD1.n64 VDD1.n1 0.155672
R2630 VDD1.n64 VDD1.n63 0.155672
R2631 VDD1.n63 VDD1.n5 0.155672
R2632 VDD1.n56 VDD1.n5 0.155672
R2633 VDD1.n56 VDD1.n55 0.155672
R2634 VDD1.n55 VDD1.n9 0.155672
R2635 VDD1.n48 VDD1.n9 0.155672
R2636 VDD1.n48 VDD1.n47 0.155672
R2637 VDD1.n47 VDD1.n13 0.155672
R2638 VDD1.n40 VDD1.n13 0.155672
R2639 VDD1.n40 VDD1.n39 0.155672
R2640 VDD1.n39 VDD1.n19 0.155672
R2641 VDD1.n32 VDD1.n19 0.155672
R2642 VDD1.n32 VDD1.n31 0.155672
R2643 VDD1.n31 VDD1.n23 0.155672
R2644 VDD1.n104 VDD1.n96 0.155672
R2645 VDD1.n105 VDD1.n104 0.155672
R2646 VDD1.n105 VDD1.n92 0.155672
R2647 VDD1.n112 VDD1.n92 0.155672
R2648 VDD1.n113 VDD1.n112 0.155672
R2649 VDD1.n113 VDD1.n88 0.155672
R2650 VDD1.n122 VDD1.n88 0.155672
R2651 VDD1.n123 VDD1.n122 0.155672
R2652 VDD1.n123 VDD1.n84 0.155672
R2653 VDD1.n130 VDD1.n84 0.155672
R2654 VDD1.n131 VDD1.n130 0.155672
R2655 VDD1.n131 VDD1.n80 0.155672
R2656 VDD1.n138 VDD1.n80 0.155672
R2657 VDD1.n139 VDD1.n138 0.155672
R2658 VDD1.n139 VDD1.n76 0.155672
R2659 VDD1.n146 VDD1.n76 0.155672
C0 VDD2 VP 0.420521f
C1 VDD2 VTAIL 12.3726f
C2 VP VN 6.8053f
C3 VN VTAIL 10.025701f
C4 VP VTAIL 10.0402f
C5 VDD1 VDD2 1.3446f
C6 VDD1 VN 0.150315f
C7 VDD1 VP 10.243401f
C8 VDD1 VTAIL 12.332999f
C9 VDD2 VN 9.97776f
C10 VDD2 B 5.997463f
C11 VDD1 B 5.957073f
C12 VTAIL B 7.740934f
C13 VN B 12.340211f
C14 VP B 10.593061f
C15 VDD1.n0 B 0.033621f
C16 VDD1.n1 B 0.02272f
C17 VDD1.n2 B 0.012209f
C18 VDD1.n3 B 0.028857f
C19 VDD1.n4 B 0.012927f
C20 VDD1.n5 B 0.02272f
C21 VDD1.n6 B 0.012209f
C22 VDD1.n7 B 0.028857f
C23 VDD1.n8 B 0.012927f
C24 VDD1.n9 B 0.02272f
C25 VDD1.n10 B 0.012209f
C26 VDD1.n11 B 0.028857f
C27 VDD1.n12 B 0.012568f
C28 VDD1.n13 B 0.02272f
C29 VDD1.n14 B 0.012568f
C30 VDD1.n15 B 0.012209f
C31 VDD1.n16 B 0.028857f
C32 VDD1.n17 B 0.028857f
C33 VDD1.n18 B 0.012927f
C34 VDD1.n19 B 0.02272f
C35 VDD1.n20 B 0.012209f
C36 VDD1.n21 B 0.028857f
C37 VDD1.n22 B 0.012927f
C38 VDD1.n23 B 1.30686f
C39 VDD1.n24 B 0.012209f
C40 VDD1.t8 B 0.048932f
C41 VDD1.n25 B 0.177677f
C42 VDD1.n26 B 0.0204f
C43 VDD1.n27 B 0.021643f
C44 VDD1.n28 B 0.028857f
C45 VDD1.n29 B 0.012927f
C46 VDD1.n30 B 0.012209f
C47 VDD1.n31 B 0.02272f
C48 VDD1.n32 B 0.02272f
C49 VDD1.n33 B 0.012209f
C50 VDD1.n34 B 0.012927f
C51 VDD1.n35 B 0.028857f
C52 VDD1.n36 B 0.028857f
C53 VDD1.n37 B 0.012927f
C54 VDD1.n38 B 0.012209f
C55 VDD1.n39 B 0.02272f
C56 VDD1.n40 B 0.02272f
C57 VDD1.n41 B 0.012209f
C58 VDD1.n42 B 0.012927f
C59 VDD1.n43 B 0.028857f
C60 VDD1.n44 B 0.028857f
C61 VDD1.n45 B 0.012927f
C62 VDD1.n46 B 0.012209f
C63 VDD1.n47 B 0.02272f
C64 VDD1.n48 B 0.02272f
C65 VDD1.n49 B 0.012209f
C66 VDD1.n50 B 0.012927f
C67 VDD1.n51 B 0.028857f
C68 VDD1.n52 B 0.028857f
C69 VDD1.n53 B 0.012927f
C70 VDD1.n54 B 0.012209f
C71 VDD1.n55 B 0.02272f
C72 VDD1.n56 B 0.02272f
C73 VDD1.n57 B 0.012209f
C74 VDD1.n58 B 0.012927f
C75 VDD1.n59 B 0.028857f
C76 VDD1.n60 B 0.028857f
C77 VDD1.n61 B 0.012927f
C78 VDD1.n62 B 0.012209f
C79 VDD1.n63 B 0.02272f
C80 VDD1.n64 B 0.02272f
C81 VDD1.n65 B 0.012209f
C82 VDD1.n66 B 0.012927f
C83 VDD1.n67 B 0.028857f
C84 VDD1.n68 B 0.065452f
C85 VDD1.n69 B 0.012927f
C86 VDD1.n70 B 0.012209f
C87 VDD1.n71 B 0.053447f
C88 VDD1.n72 B 0.056788f
C89 VDD1.t3 B 0.243995f
C90 VDD1.t0 B 0.243995f
C91 VDD1.n73 B 2.18997f
C92 VDD1.n74 B 0.468186f
C93 VDD1.n75 B 0.033621f
C94 VDD1.n76 B 0.02272f
C95 VDD1.n77 B 0.012209f
C96 VDD1.n78 B 0.028857f
C97 VDD1.n79 B 0.012927f
C98 VDD1.n80 B 0.02272f
C99 VDD1.n81 B 0.012209f
C100 VDD1.n82 B 0.028857f
C101 VDD1.n83 B 0.012927f
C102 VDD1.n84 B 0.02272f
C103 VDD1.n85 B 0.012209f
C104 VDD1.n86 B 0.028857f
C105 VDD1.n87 B 0.012568f
C106 VDD1.n88 B 0.02272f
C107 VDD1.n89 B 0.012927f
C108 VDD1.n90 B 0.028857f
C109 VDD1.n91 B 0.012927f
C110 VDD1.n92 B 0.02272f
C111 VDD1.n93 B 0.012209f
C112 VDD1.n94 B 0.028857f
C113 VDD1.n95 B 0.012927f
C114 VDD1.n96 B 1.30686f
C115 VDD1.n97 B 0.012209f
C116 VDD1.t4 B 0.048932f
C117 VDD1.n98 B 0.177677f
C118 VDD1.n99 B 0.0204f
C119 VDD1.n100 B 0.021643f
C120 VDD1.n101 B 0.028857f
C121 VDD1.n102 B 0.012927f
C122 VDD1.n103 B 0.012209f
C123 VDD1.n104 B 0.02272f
C124 VDD1.n105 B 0.02272f
C125 VDD1.n106 B 0.012209f
C126 VDD1.n107 B 0.012927f
C127 VDD1.n108 B 0.028857f
C128 VDD1.n109 B 0.028857f
C129 VDD1.n110 B 0.012927f
C130 VDD1.n111 B 0.012209f
C131 VDD1.n112 B 0.02272f
C132 VDD1.n113 B 0.02272f
C133 VDD1.n114 B 0.012209f
C134 VDD1.n115 B 0.012209f
C135 VDD1.n116 B 0.012927f
C136 VDD1.n117 B 0.028857f
C137 VDD1.n118 B 0.028857f
C138 VDD1.n119 B 0.028857f
C139 VDD1.n120 B 0.012568f
C140 VDD1.n121 B 0.012209f
C141 VDD1.n122 B 0.02272f
C142 VDD1.n123 B 0.02272f
C143 VDD1.n124 B 0.012209f
C144 VDD1.n125 B 0.012927f
C145 VDD1.n126 B 0.028857f
C146 VDD1.n127 B 0.028857f
C147 VDD1.n128 B 0.012927f
C148 VDD1.n129 B 0.012209f
C149 VDD1.n130 B 0.02272f
C150 VDD1.n131 B 0.02272f
C151 VDD1.n132 B 0.012209f
C152 VDD1.n133 B 0.012927f
C153 VDD1.n134 B 0.028857f
C154 VDD1.n135 B 0.028857f
C155 VDD1.n136 B 0.012927f
C156 VDD1.n137 B 0.012209f
C157 VDD1.n138 B 0.02272f
C158 VDD1.n139 B 0.02272f
C159 VDD1.n140 B 0.012209f
C160 VDD1.n141 B 0.012927f
C161 VDD1.n142 B 0.028857f
C162 VDD1.n143 B 0.065452f
C163 VDD1.n144 B 0.012927f
C164 VDD1.n145 B 0.012209f
C165 VDD1.n146 B 0.053447f
C166 VDD1.n147 B 0.056788f
C167 VDD1.t5 B 0.243995f
C168 VDD1.t2 B 0.243995f
C169 VDD1.n148 B 2.18996f
C170 VDD1.n149 B 0.461636f
C171 VDD1.t6 B 0.243995f
C172 VDD1.t7 B 0.243995f
C173 VDD1.n150 B 2.196f
C174 VDD1.n151 B 2.20467f
C175 VDD1.t9 B 0.243995f
C176 VDD1.t1 B 0.243995f
C177 VDD1.n152 B 2.18996f
C178 VDD1.n153 B 2.51569f
C179 VP.n0 B 0.032153f
C180 VP.t2 B 1.57676f
C181 VP.n1 B 0.054102f
C182 VP.n2 B 0.032153f
C183 VP.t7 B 1.57676f
C184 VP.n3 B 0.598725f
C185 VP.n4 B 0.032153f
C186 VP.t4 B 1.57676f
C187 VP.n5 B 0.568386f
C188 VP.n6 B 0.032153f
C189 VP.t5 B 1.57676f
C190 VP.n7 B 0.631576f
C191 VP.n8 B 0.032153f
C192 VP.t8 B 1.57676f
C193 VP.n9 B 0.054102f
C194 VP.n10 B 0.032153f
C195 VP.t9 B 1.57676f
C196 VP.n11 B 0.598725f
C197 VP.n12 B 0.032153f
C198 VP.t6 B 1.57676f
C199 VP.n13 B 0.615194f
C200 VP.t1 B 1.65158f
C201 VP.n14 B 0.64472f
C202 VP.n15 B 0.171245f
C203 VP.n16 B 0.039215f
C204 VP.n17 B 0.04022f
C205 VP.n18 B 0.05366f
C206 VP.n19 B 0.032153f
C207 VP.n20 B 0.032153f
C208 VP.n21 B 0.032153f
C209 VP.n22 B 0.05366f
C210 VP.n23 B 0.04022f
C211 VP.t0 B 1.57676f
C212 VP.n24 B 0.568386f
C213 VP.n25 B 0.039215f
C214 VP.n26 B 0.032153f
C215 VP.n27 B 0.032153f
C216 VP.n28 B 0.032153f
C217 VP.n29 B 0.026253f
C218 VP.n30 B 0.05274f
C219 VP.n31 B 0.631576f
C220 VP.n32 B 1.61069f
C221 VP.n33 B 1.63511f
C222 VP.n34 B 0.032153f
C223 VP.n35 B 0.05274f
C224 VP.n36 B 0.026253f
C225 VP.n37 B 0.054102f
C226 VP.n38 B 0.032153f
C227 VP.n39 B 0.032153f
C228 VP.n40 B 0.039215f
C229 VP.n41 B 0.04022f
C230 VP.n42 B 0.05366f
C231 VP.n43 B 0.032153f
C232 VP.n44 B 0.032153f
C233 VP.n45 B 0.032153f
C234 VP.n46 B 0.05366f
C235 VP.n47 B 0.04022f
C236 VP.t3 B 1.57676f
C237 VP.n48 B 0.568386f
C238 VP.n49 B 0.039215f
C239 VP.n50 B 0.032153f
C240 VP.n51 B 0.032153f
C241 VP.n52 B 0.032153f
C242 VP.n53 B 0.026253f
C243 VP.n54 B 0.05274f
C244 VP.n55 B 0.631576f
C245 VP.n56 B 0.028751f
C246 VTAIL.t16 B 0.259368f
C247 VTAIL.t17 B 0.259368f
C248 VTAIL.n0 B 2.25571f
C249 VTAIL.n1 B 0.420299f
C250 VTAIL.n2 B 0.035739f
C251 VTAIL.n3 B 0.024151f
C252 VTAIL.n4 B 0.012978f
C253 VTAIL.n5 B 0.030675f
C254 VTAIL.n6 B 0.013741f
C255 VTAIL.n7 B 0.024151f
C256 VTAIL.n8 B 0.012978f
C257 VTAIL.n9 B 0.030675f
C258 VTAIL.n10 B 0.013741f
C259 VTAIL.n11 B 0.024151f
C260 VTAIL.n12 B 0.012978f
C261 VTAIL.n13 B 0.030675f
C262 VTAIL.n14 B 0.01336f
C263 VTAIL.n15 B 0.024151f
C264 VTAIL.n16 B 0.013741f
C265 VTAIL.n17 B 0.030675f
C266 VTAIL.n18 B 0.013741f
C267 VTAIL.n19 B 0.024151f
C268 VTAIL.n20 B 0.012978f
C269 VTAIL.n21 B 0.030675f
C270 VTAIL.n22 B 0.013741f
C271 VTAIL.n23 B 1.3892f
C272 VTAIL.n24 B 0.012978f
C273 VTAIL.t8 B 0.052015f
C274 VTAIL.n25 B 0.188872f
C275 VTAIL.n26 B 0.021685f
C276 VTAIL.n27 B 0.023006f
C277 VTAIL.n28 B 0.030675f
C278 VTAIL.n29 B 0.013741f
C279 VTAIL.n30 B 0.012978f
C280 VTAIL.n31 B 0.024151f
C281 VTAIL.n32 B 0.024151f
C282 VTAIL.n33 B 0.012978f
C283 VTAIL.n34 B 0.013741f
C284 VTAIL.n35 B 0.030675f
C285 VTAIL.n36 B 0.030675f
C286 VTAIL.n37 B 0.013741f
C287 VTAIL.n38 B 0.012978f
C288 VTAIL.n39 B 0.024151f
C289 VTAIL.n40 B 0.024151f
C290 VTAIL.n41 B 0.012978f
C291 VTAIL.n42 B 0.012978f
C292 VTAIL.n43 B 0.013741f
C293 VTAIL.n44 B 0.030675f
C294 VTAIL.n45 B 0.030675f
C295 VTAIL.n46 B 0.030675f
C296 VTAIL.n47 B 0.01336f
C297 VTAIL.n48 B 0.012978f
C298 VTAIL.n49 B 0.024151f
C299 VTAIL.n50 B 0.024151f
C300 VTAIL.n51 B 0.012978f
C301 VTAIL.n52 B 0.013741f
C302 VTAIL.n53 B 0.030675f
C303 VTAIL.n54 B 0.030675f
C304 VTAIL.n55 B 0.013741f
C305 VTAIL.n56 B 0.012978f
C306 VTAIL.n57 B 0.024151f
C307 VTAIL.n58 B 0.024151f
C308 VTAIL.n59 B 0.012978f
C309 VTAIL.n60 B 0.013741f
C310 VTAIL.n61 B 0.030675f
C311 VTAIL.n62 B 0.030675f
C312 VTAIL.n63 B 0.013741f
C313 VTAIL.n64 B 0.012978f
C314 VTAIL.n65 B 0.024151f
C315 VTAIL.n66 B 0.024151f
C316 VTAIL.n67 B 0.012978f
C317 VTAIL.n68 B 0.013741f
C318 VTAIL.n69 B 0.030675f
C319 VTAIL.n70 B 0.069576f
C320 VTAIL.n71 B 0.013741f
C321 VTAIL.n72 B 0.012978f
C322 VTAIL.n73 B 0.056815f
C323 VTAIL.n74 B 0.039287f
C324 VTAIL.n75 B 0.22379f
C325 VTAIL.t1 B 0.259368f
C326 VTAIL.t0 B 0.259368f
C327 VTAIL.n76 B 2.25571f
C328 VTAIL.n77 B 0.462229f
C329 VTAIL.t5 B 0.259368f
C330 VTAIL.t6 B 0.259368f
C331 VTAIL.n78 B 2.25571f
C332 VTAIL.n79 B 1.81271f
C333 VTAIL.t15 B 0.259368f
C334 VTAIL.t10 B 0.259368f
C335 VTAIL.n80 B 2.25572f
C336 VTAIL.n81 B 1.8127f
C337 VTAIL.t14 B 0.259368f
C338 VTAIL.t11 B 0.259368f
C339 VTAIL.n82 B 2.25572f
C340 VTAIL.n83 B 0.462217f
C341 VTAIL.n84 B 0.035739f
C342 VTAIL.n85 B 0.024151f
C343 VTAIL.n86 B 0.012978f
C344 VTAIL.n87 B 0.030675f
C345 VTAIL.n88 B 0.013741f
C346 VTAIL.n89 B 0.024151f
C347 VTAIL.n90 B 0.012978f
C348 VTAIL.n91 B 0.030675f
C349 VTAIL.n92 B 0.013741f
C350 VTAIL.n93 B 0.024151f
C351 VTAIL.n94 B 0.012978f
C352 VTAIL.n95 B 0.030675f
C353 VTAIL.n96 B 0.01336f
C354 VTAIL.n97 B 0.024151f
C355 VTAIL.n98 B 0.01336f
C356 VTAIL.n99 B 0.012978f
C357 VTAIL.n100 B 0.030675f
C358 VTAIL.n101 B 0.030675f
C359 VTAIL.n102 B 0.013741f
C360 VTAIL.n103 B 0.024151f
C361 VTAIL.n104 B 0.012978f
C362 VTAIL.n105 B 0.030675f
C363 VTAIL.n106 B 0.013741f
C364 VTAIL.n107 B 1.3892f
C365 VTAIL.n108 B 0.012978f
C366 VTAIL.t12 B 0.052015f
C367 VTAIL.n109 B 0.188871f
C368 VTAIL.n110 B 0.021685f
C369 VTAIL.n111 B 0.023006f
C370 VTAIL.n112 B 0.030675f
C371 VTAIL.n113 B 0.013741f
C372 VTAIL.n114 B 0.012978f
C373 VTAIL.n115 B 0.024151f
C374 VTAIL.n116 B 0.024151f
C375 VTAIL.n117 B 0.012978f
C376 VTAIL.n118 B 0.013741f
C377 VTAIL.n119 B 0.030675f
C378 VTAIL.n120 B 0.030675f
C379 VTAIL.n121 B 0.013741f
C380 VTAIL.n122 B 0.012978f
C381 VTAIL.n123 B 0.024151f
C382 VTAIL.n124 B 0.024151f
C383 VTAIL.n125 B 0.012978f
C384 VTAIL.n126 B 0.013741f
C385 VTAIL.n127 B 0.030675f
C386 VTAIL.n128 B 0.030675f
C387 VTAIL.n129 B 0.013741f
C388 VTAIL.n130 B 0.012978f
C389 VTAIL.n131 B 0.024151f
C390 VTAIL.n132 B 0.024151f
C391 VTAIL.n133 B 0.012978f
C392 VTAIL.n134 B 0.013741f
C393 VTAIL.n135 B 0.030675f
C394 VTAIL.n136 B 0.030675f
C395 VTAIL.n137 B 0.013741f
C396 VTAIL.n138 B 0.012978f
C397 VTAIL.n139 B 0.024151f
C398 VTAIL.n140 B 0.024151f
C399 VTAIL.n141 B 0.012978f
C400 VTAIL.n142 B 0.013741f
C401 VTAIL.n143 B 0.030675f
C402 VTAIL.n144 B 0.030675f
C403 VTAIL.n145 B 0.013741f
C404 VTAIL.n146 B 0.012978f
C405 VTAIL.n147 B 0.024151f
C406 VTAIL.n148 B 0.024151f
C407 VTAIL.n149 B 0.012978f
C408 VTAIL.n150 B 0.013741f
C409 VTAIL.n151 B 0.030675f
C410 VTAIL.n152 B 0.069576f
C411 VTAIL.n153 B 0.013741f
C412 VTAIL.n154 B 0.012978f
C413 VTAIL.n155 B 0.056815f
C414 VTAIL.n156 B 0.039287f
C415 VTAIL.n157 B 0.22379f
C416 VTAIL.t4 B 0.259368f
C417 VTAIL.t3 B 0.259368f
C418 VTAIL.n158 B 2.25572f
C419 VTAIL.n159 B 0.443432f
C420 VTAIL.t7 B 0.259368f
C421 VTAIL.t9 B 0.259368f
C422 VTAIL.n160 B 2.25572f
C423 VTAIL.n161 B 0.462217f
C424 VTAIL.n162 B 0.035739f
C425 VTAIL.n163 B 0.024151f
C426 VTAIL.n164 B 0.012978f
C427 VTAIL.n165 B 0.030675f
C428 VTAIL.n166 B 0.013741f
C429 VTAIL.n167 B 0.024151f
C430 VTAIL.n168 B 0.012978f
C431 VTAIL.n169 B 0.030675f
C432 VTAIL.n170 B 0.013741f
C433 VTAIL.n171 B 0.024151f
C434 VTAIL.n172 B 0.012978f
C435 VTAIL.n173 B 0.030675f
C436 VTAIL.n174 B 0.01336f
C437 VTAIL.n175 B 0.024151f
C438 VTAIL.n176 B 0.01336f
C439 VTAIL.n177 B 0.012978f
C440 VTAIL.n178 B 0.030675f
C441 VTAIL.n179 B 0.030675f
C442 VTAIL.n180 B 0.013741f
C443 VTAIL.n181 B 0.024151f
C444 VTAIL.n182 B 0.012978f
C445 VTAIL.n183 B 0.030675f
C446 VTAIL.n184 B 0.013741f
C447 VTAIL.n185 B 1.3892f
C448 VTAIL.n186 B 0.012978f
C449 VTAIL.t2 B 0.052015f
C450 VTAIL.n187 B 0.188871f
C451 VTAIL.n188 B 0.021685f
C452 VTAIL.n189 B 0.023006f
C453 VTAIL.n190 B 0.030675f
C454 VTAIL.n191 B 0.013741f
C455 VTAIL.n192 B 0.012978f
C456 VTAIL.n193 B 0.024151f
C457 VTAIL.n194 B 0.024151f
C458 VTAIL.n195 B 0.012978f
C459 VTAIL.n196 B 0.013741f
C460 VTAIL.n197 B 0.030675f
C461 VTAIL.n198 B 0.030675f
C462 VTAIL.n199 B 0.013741f
C463 VTAIL.n200 B 0.012978f
C464 VTAIL.n201 B 0.024151f
C465 VTAIL.n202 B 0.024151f
C466 VTAIL.n203 B 0.012978f
C467 VTAIL.n204 B 0.013741f
C468 VTAIL.n205 B 0.030675f
C469 VTAIL.n206 B 0.030675f
C470 VTAIL.n207 B 0.013741f
C471 VTAIL.n208 B 0.012978f
C472 VTAIL.n209 B 0.024151f
C473 VTAIL.n210 B 0.024151f
C474 VTAIL.n211 B 0.012978f
C475 VTAIL.n212 B 0.013741f
C476 VTAIL.n213 B 0.030675f
C477 VTAIL.n214 B 0.030675f
C478 VTAIL.n215 B 0.013741f
C479 VTAIL.n216 B 0.012978f
C480 VTAIL.n217 B 0.024151f
C481 VTAIL.n218 B 0.024151f
C482 VTAIL.n219 B 0.012978f
C483 VTAIL.n220 B 0.013741f
C484 VTAIL.n221 B 0.030675f
C485 VTAIL.n222 B 0.030675f
C486 VTAIL.n223 B 0.013741f
C487 VTAIL.n224 B 0.012978f
C488 VTAIL.n225 B 0.024151f
C489 VTAIL.n226 B 0.024151f
C490 VTAIL.n227 B 0.012978f
C491 VTAIL.n228 B 0.013741f
C492 VTAIL.n229 B 0.030675f
C493 VTAIL.n230 B 0.069576f
C494 VTAIL.n231 B 0.013741f
C495 VTAIL.n232 B 0.012978f
C496 VTAIL.n233 B 0.056815f
C497 VTAIL.n234 B 0.039287f
C498 VTAIL.n235 B 1.48236f
C499 VTAIL.n236 B 0.035739f
C500 VTAIL.n237 B 0.024151f
C501 VTAIL.n238 B 0.012978f
C502 VTAIL.n239 B 0.030675f
C503 VTAIL.n240 B 0.013741f
C504 VTAIL.n241 B 0.024151f
C505 VTAIL.n242 B 0.012978f
C506 VTAIL.n243 B 0.030675f
C507 VTAIL.n244 B 0.013741f
C508 VTAIL.n245 B 0.024151f
C509 VTAIL.n246 B 0.012978f
C510 VTAIL.n247 B 0.030675f
C511 VTAIL.n248 B 0.01336f
C512 VTAIL.n249 B 0.024151f
C513 VTAIL.n250 B 0.013741f
C514 VTAIL.n251 B 0.030675f
C515 VTAIL.n252 B 0.013741f
C516 VTAIL.n253 B 0.024151f
C517 VTAIL.n254 B 0.012978f
C518 VTAIL.n255 B 0.030675f
C519 VTAIL.n256 B 0.013741f
C520 VTAIL.n257 B 1.3892f
C521 VTAIL.n258 B 0.012978f
C522 VTAIL.t13 B 0.052015f
C523 VTAIL.n259 B 0.188872f
C524 VTAIL.n260 B 0.021685f
C525 VTAIL.n261 B 0.023006f
C526 VTAIL.n262 B 0.030675f
C527 VTAIL.n263 B 0.013741f
C528 VTAIL.n264 B 0.012978f
C529 VTAIL.n265 B 0.024151f
C530 VTAIL.n266 B 0.024151f
C531 VTAIL.n267 B 0.012978f
C532 VTAIL.n268 B 0.013741f
C533 VTAIL.n269 B 0.030675f
C534 VTAIL.n270 B 0.030675f
C535 VTAIL.n271 B 0.013741f
C536 VTAIL.n272 B 0.012978f
C537 VTAIL.n273 B 0.024151f
C538 VTAIL.n274 B 0.024151f
C539 VTAIL.n275 B 0.012978f
C540 VTAIL.n276 B 0.012978f
C541 VTAIL.n277 B 0.013741f
C542 VTAIL.n278 B 0.030675f
C543 VTAIL.n279 B 0.030675f
C544 VTAIL.n280 B 0.030675f
C545 VTAIL.n281 B 0.01336f
C546 VTAIL.n282 B 0.012978f
C547 VTAIL.n283 B 0.024151f
C548 VTAIL.n284 B 0.024151f
C549 VTAIL.n285 B 0.012978f
C550 VTAIL.n286 B 0.013741f
C551 VTAIL.n287 B 0.030675f
C552 VTAIL.n288 B 0.030675f
C553 VTAIL.n289 B 0.013741f
C554 VTAIL.n290 B 0.012978f
C555 VTAIL.n291 B 0.024151f
C556 VTAIL.n292 B 0.024151f
C557 VTAIL.n293 B 0.012978f
C558 VTAIL.n294 B 0.013741f
C559 VTAIL.n295 B 0.030675f
C560 VTAIL.n296 B 0.030675f
C561 VTAIL.n297 B 0.013741f
C562 VTAIL.n298 B 0.012978f
C563 VTAIL.n299 B 0.024151f
C564 VTAIL.n300 B 0.024151f
C565 VTAIL.n301 B 0.012978f
C566 VTAIL.n302 B 0.013741f
C567 VTAIL.n303 B 0.030675f
C568 VTAIL.n304 B 0.069576f
C569 VTAIL.n305 B 0.013741f
C570 VTAIL.n306 B 0.012978f
C571 VTAIL.n307 B 0.056815f
C572 VTAIL.n308 B 0.039287f
C573 VTAIL.n309 B 1.48236f
C574 VTAIL.t18 B 0.259368f
C575 VTAIL.t19 B 0.259368f
C576 VTAIL.n310 B 2.25571f
C577 VTAIL.n311 B 0.37468f
C578 VDD2.n0 B 0.033597f
C579 VDD2.n1 B 0.022704f
C580 VDD2.n2 B 0.0122f
C581 VDD2.n3 B 0.028836f
C582 VDD2.n4 B 0.012918f
C583 VDD2.n5 B 0.022704f
C584 VDD2.n6 B 0.0122f
C585 VDD2.n7 B 0.028836f
C586 VDD2.n8 B 0.012918f
C587 VDD2.n9 B 0.022704f
C588 VDD2.n10 B 0.0122f
C589 VDD2.n11 B 0.028836f
C590 VDD2.n12 B 0.012559f
C591 VDD2.n13 B 0.022704f
C592 VDD2.n14 B 0.012918f
C593 VDD2.n15 B 0.028836f
C594 VDD2.n16 B 0.012918f
C595 VDD2.n17 B 0.022704f
C596 VDD2.n18 B 0.0122f
C597 VDD2.n19 B 0.028836f
C598 VDD2.n20 B 0.012918f
C599 VDD2.n21 B 1.30592f
C600 VDD2.n22 B 0.0122f
C601 VDD2.t3 B 0.048897f
C602 VDD2.n23 B 0.177549f
C603 VDD2.n24 B 0.020385f
C604 VDD2.n25 B 0.021627f
C605 VDD2.n26 B 0.028836f
C606 VDD2.n27 B 0.012918f
C607 VDD2.n28 B 0.0122f
C608 VDD2.n29 B 0.022704f
C609 VDD2.n30 B 0.022704f
C610 VDD2.n31 B 0.0122f
C611 VDD2.n32 B 0.012918f
C612 VDD2.n33 B 0.028836f
C613 VDD2.n34 B 0.028836f
C614 VDD2.n35 B 0.012918f
C615 VDD2.n36 B 0.0122f
C616 VDD2.n37 B 0.022704f
C617 VDD2.n38 B 0.022704f
C618 VDD2.n39 B 0.0122f
C619 VDD2.n40 B 0.0122f
C620 VDD2.n41 B 0.012918f
C621 VDD2.n42 B 0.028836f
C622 VDD2.n43 B 0.028836f
C623 VDD2.n44 B 0.028836f
C624 VDD2.n45 B 0.012559f
C625 VDD2.n46 B 0.0122f
C626 VDD2.n47 B 0.022704f
C627 VDD2.n48 B 0.022704f
C628 VDD2.n49 B 0.0122f
C629 VDD2.n50 B 0.012918f
C630 VDD2.n51 B 0.028836f
C631 VDD2.n52 B 0.028836f
C632 VDD2.n53 B 0.012918f
C633 VDD2.n54 B 0.0122f
C634 VDD2.n55 B 0.022704f
C635 VDD2.n56 B 0.022704f
C636 VDD2.n57 B 0.0122f
C637 VDD2.n58 B 0.012918f
C638 VDD2.n59 B 0.028836f
C639 VDD2.n60 B 0.028836f
C640 VDD2.n61 B 0.012918f
C641 VDD2.n62 B 0.0122f
C642 VDD2.n63 B 0.022704f
C643 VDD2.n64 B 0.022704f
C644 VDD2.n65 B 0.0122f
C645 VDD2.n66 B 0.012918f
C646 VDD2.n67 B 0.028836f
C647 VDD2.n68 B 0.065405f
C648 VDD2.n69 B 0.012918f
C649 VDD2.n70 B 0.0122f
C650 VDD2.n71 B 0.053409f
C651 VDD2.n72 B 0.056748f
C652 VDD2.t9 B 0.24382f
C653 VDD2.t6 B 0.24382f
C654 VDD2.n73 B 2.18839f
C655 VDD2.n74 B 0.461305f
C656 VDD2.t2 B 0.24382f
C657 VDD2.t4 B 0.24382f
C658 VDD2.n75 B 2.19443f
C659 VDD2.n76 B 2.11894f
C660 VDD2.n77 B 0.033597f
C661 VDD2.n78 B 0.022704f
C662 VDD2.n79 B 0.0122f
C663 VDD2.n80 B 0.028836f
C664 VDD2.n81 B 0.012918f
C665 VDD2.n82 B 0.022704f
C666 VDD2.n83 B 0.0122f
C667 VDD2.n84 B 0.028836f
C668 VDD2.n85 B 0.012918f
C669 VDD2.n86 B 0.022704f
C670 VDD2.n87 B 0.0122f
C671 VDD2.n88 B 0.028836f
C672 VDD2.n89 B 0.012559f
C673 VDD2.n90 B 0.022704f
C674 VDD2.n91 B 0.012559f
C675 VDD2.n92 B 0.0122f
C676 VDD2.n93 B 0.028836f
C677 VDD2.n94 B 0.028836f
C678 VDD2.n95 B 0.012918f
C679 VDD2.n96 B 0.022704f
C680 VDD2.n97 B 0.0122f
C681 VDD2.n98 B 0.028836f
C682 VDD2.n99 B 0.012918f
C683 VDD2.n100 B 1.30592f
C684 VDD2.n101 B 0.0122f
C685 VDD2.t0 B 0.048897f
C686 VDD2.n102 B 0.177549f
C687 VDD2.n103 B 0.020385f
C688 VDD2.n104 B 0.021627f
C689 VDD2.n105 B 0.028836f
C690 VDD2.n106 B 0.012918f
C691 VDD2.n107 B 0.0122f
C692 VDD2.n108 B 0.022704f
C693 VDD2.n109 B 0.022704f
C694 VDD2.n110 B 0.0122f
C695 VDD2.n111 B 0.012918f
C696 VDD2.n112 B 0.028836f
C697 VDD2.n113 B 0.028836f
C698 VDD2.n114 B 0.012918f
C699 VDD2.n115 B 0.0122f
C700 VDD2.n116 B 0.022704f
C701 VDD2.n117 B 0.022704f
C702 VDD2.n118 B 0.0122f
C703 VDD2.n119 B 0.012918f
C704 VDD2.n120 B 0.028836f
C705 VDD2.n121 B 0.028836f
C706 VDD2.n122 B 0.012918f
C707 VDD2.n123 B 0.0122f
C708 VDD2.n124 B 0.022704f
C709 VDD2.n125 B 0.022704f
C710 VDD2.n126 B 0.0122f
C711 VDD2.n127 B 0.012918f
C712 VDD2.n128 B 0.028836f
C713 VDD2.n129 B 0.028836f
C714 VDD2.n130 B 0.012918f
C715 VDD2.n131 B 0.0122f
C716 VDD2.n132 B 0.022704f
C717 VDD2.n133 B 0.022704f
C718 VDD2.n134 B 0.0122f
C719 VDD2.n135 B 0.012918f
C720 VDD2.n136 B 0.028836f
C721 VDD2.n137 B 0.028836f
C722 VDD2.n138 B 0.012918f
C723 VDD2.n139 B 0.0122f
C724 VDD2.n140 B 0.022704f
C725 VDD2.n141 B 0.022704f
C726 VDD2.n142 B 0.0122f
C727 VDD2.n143 B 0.012918f
C728 VDD2.n144 B 0.028836f
C729 VDD2.n145 B 0.065405f
C730 VDD2.n146 B 0.012918f
C731 VDD2.n147 B 0.0122f
C732 VDD2.n148 B 0.053409f
C733 VDD2.n149 B 0.0526f
C734 VDD2.n150 B 2.28614f
C735 VDD2.t7 B 0.24382f
C736 VDD2.t5 B 0.24382f
C737 VDD2.n151 B 2.18839f
C738 VDD2.n152 B 0.323688f
C739 VDD2.t8 B 0.24382f
C740 VDD2.t1 B 0.24382f
C741 VDD2.n153 B 2.1944f
C742 VN.n0 B 0.031861f
C743 VN.t6 B 1.56246f
C744 VN.n1 B 0.053611f
C745 VN.n2 B 0.031861f
C746 VN.t1 B 1.56246f
C747 VN.n3 B 0.593297f
C748 VN.n4 B 0.031861f
C749 VN.t2 B 1.56246f
C750 VN.n5 B 0.609616f
C751 VN.t3 B 1.6366f
C752 VN.n6 B 0.638875f
C753 VN.n7 B 0.169692f
C754 VN.n8 B 0.038859f
C755 VN.n9 B 0.039856f
C756 VN.n10 B 0.053173f
C757 VN.n11 B 0.031861f
C758 VN.n12 B 0.031861f
C759 VN.n13 B 0.031861f
C760 VN.n14 B 0.053173f
C761 VN.n15 B 0.039856f
C762 VN.t0 B 1.56246f
C763 VN.n16 B 0.563233f
C764 VN.n17 B 0.038859f
C765 VN.n18 B 0.031861f
C766 VN.n19 B 0.031861f
C767 VN.n20 B 0.031861f
C768 VN.n21 B 0.026015f
C769 VN.n22 B 0.052262f
C770 VN.n23 B 0.62585f
C771 VN.n24 B 0.02849f
C772 VN.n25 B 0.031861f
C773 VN.t4 B 1.56246f
C774 VN.n26 B 0.053611f
C775 VN.n27 B 0.031861f
C776 VN.t9 B 1.56246f
C777 VN.n28 B 0.563233f
C778 VN.t5 B 1.56246f
C779 VN.n29 B 0.593297f
C780 VN.n30 B 0.031861f
C781 VN.t8 B 1.56246f
C782 VN.n31 B 0.609616f
C783 VN.t7 B 1.6366f
C784 VN.n32 B 0.638875f
C785 VN.n33 B 0.169692f
C786 VN.n34 B 0.038859f
C787 VN.n35 B 0.039856f
C788 VN.n36 B 0.053173f
C789 VN.n37 B 0.031861f
C790 VN.n38 B 0.031861f
C791 VN.n39 B 0.031861f
C792 VN.n40 B 0.053173f
C793 VN.n41 B 0.039856f
C794 VN.n42 B 0.038859f
C795 VN.n43 B 0.031861f
C796 VN.n44 B 0.031861f
C797 VN.n45 B 0.031861f
C798 VN.n46 B 0.026015f
C799 VN.n47 B 0.052262f
C800 VN.n48 B 0.62585f
C801 VN.n49 B 1.61686f
.ends

