* NGSPICE file created from diff_pair_sample_1034.ext - technology: sky130A

.subckt diff_pair_sample_1034 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=2.1645 ps=11.88 w=5.55 l=0.97
X1 B.t11 B.t9 B.t10 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0 ps=0 w=5.55 l=0.97
X2 VDD1.t6 VP.t1 VTAIL.t9 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X3 VTAIL.t2 VN.t0 VDD2.t7 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X4 B.t8 B.t6 B.t7 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0 ps=0 w=5.55 l=0.97
X5 B.t5 B.t3 B.t4 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0 ps=0 w=5.55 l=0.97
X6 VTAIL.t15 VN.t1 VDD2.t6 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X7 B.t2 B.t0 B.t1 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0 ps=0 w=5.55 l=0.97
X8 VDD2.t5 VN.t2 VTAIL.t4 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=2.1645 ps=11.88 w=5.55 l=0.97
X9 VDD2.t4 VN.t3 VTAIL.t1 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X10 VDD1.t5 VP.t2 VTAIL.t14 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X11 VTAIL.t0 VN.t4 VDD2.t3 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X12 VTAIL.t5 VN.t5 VDD2.t2 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X13 VDD2.t1 VN.t6 VTAIL.t6 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X14 VTAIL.t11 VP.t3 VDD1.t4 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X15 VTAIL.t8 VP.t4 VDD1.t3 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X16 VDD1.t2 VP.t5 VTAIL.t10 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=2.1645 ps=11.88 w=5.55 l=0.97
X17 VTAIL.t7 VP.t6 VDD1.t1 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X18 VTAIL.t13 VP.t7 VDD1.t0 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=2.1645 pd=11.88 as=0.91575 ps=5.88 w=5.55 l=0.97
X19 VDD2.t0 VN.t7 VTAIL.t3 w_n2270_n2078# sky130_fd_pr__pfet_01v8 ad=0.91575 pd=5.88 as=2.1645 ps=11.88 w=5.55 l=0.97
R0 VP.n5 VP.t4 193.565
R1 VP.n17 VP.t7 178.638
R2 VP.n27 VP.t0 178.638
R3 VP.n14 VP.t5 178.638
R4 VP.n8 VP.n7 161.3
R5 VP.n9 VP.n4 161.3
R6 VP.n11 VP.n10 161.3
R7 VP.n13 VP.n3 161.3
R8 VP.n26 VP.n0 161.3
R9 VP.n24 VP.n23 161.3
R10 VP.n22 VP.n1 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n18 VP.n2 161.3
R13 VP.n19 VP.t1 137.893
R14 VP.n25 VP.t6 137.893
R15 VP.n12 VP.t3 137.893
R16 VP.n6 VP.t2 137.893
R17 VP.n15 VP.n14 80.6037
R18 VP.n28 VP.n27 80.6037
R19 VP.n17 VP.n16 80.6037
R20 VP.n18 VP.n17 54.8066
R21 VP.n27 VP.n26 54.8066
R22 VP.n14 VP.n13 54.8066
R23 VP.n6 VP.n5 46.8936
R24 VP.n8 VP.n5 44.1212
R25 VP.n20 VP.n1 40.4934
R26 VP.n24 VP.n1 40.4934
R27 VP.n11 VP.n4 40.4934
R28 VP.n7 VP.n4 40.4934
R29 VP.n16 VP.n15 38.5544
R30 VP.n19 VP.n18 17.1274
R31 VP.n26 VP.n25 17.1274
R32 VP.n13 VP.n12 17.1274
R33 VP.n20 VP.n19 7.3406
R34 VP.n25 VP.n24 7.3406
R35 VP.n12 VP.n11 7.3406
R36 VP.n7 VP.n6 7.3406
R37 VP.n15 VP.n3 0.285035
R38 VP.n16 VP.n2 0.285035
R39 VP.n28 VP.n0 0.285035
R40 VP.n9 VP.n8 0.189894
R41 VP.n10 VP.n9 0.189894
R42 VP.n10 VP.n3 0.189894
R43 VP.n21 VP.n2 0.189894
R44 VP.n22 VP.n21 0.189894
R45 VP.n23 VP.n22 0.189894
R46 VP.n23 VP.n0 0.189894
R47 VP VP.n28 0.146778
R48 VTAIL.n11 VTAIL.t8 82.073
R49 VTAIL.n10 VTAIL.t4 82.073
R50 VTAIL.n7 VTAIL.t5 82.073
R51 VTAIL.n15 VTAIL.t3 82.0728
R52 VTAIL.n2 VTAIL.t2 82.0728
R53 VTAIL.n3 VTAIL.t12 82.0728
R54 VTAIL.n6 VTAIL.t13 82.0728
R55 VTAIL.n14 VTAIL.t10 82.0728
R56 VTAIL.n13 VTAIL.n12 76.2163
R57 VTAIL.n9 VTAIL.n8 76.2163
R58 VTAIL.n1 VTAIL.n0 76.216
R59 VTAIL.n5 VTAIL.n4 76.216
R60 VTAIL.n15 VTAIL.n14 18.2721
R61 VTAIL.n7 VTAIL.n6 18.2721
R62 VTAIL.n0 VTAIL.t6 5.85726
R63 VTAIL.n0 VTAIL.t15 5.85726
R64 VTAIL.n4 VTAIL.t9 5.85726
R65 VTAIL.n4 VTAIL.t7 5.85726
R66 VTAIL.n12 VTAIL.t14 5.85726
R67 VTAIL.n12 VTAIL.t11 5.85726
R68 VTAIL.n8 VTAIL.t1 5.85726
R69 VTAIL.n8 VTAIL.t0 5.85726
R70 VTAIL.n9 VTAIL.n7 1.12119
R71 VTAIL.n10 VTAIL.n9 1.12119
R72 VTAIL.n13 VTAIL.n11 1.12119
R73 VTAIL.n14 VTAIL.n13 1.12119
R74 VTAIL.n6 VTAIL.n5 1.12119
R75 VTAIL.n5 VTAIL.n3 1.12119
R76 VTAIL.n2 VTAIL.n1 1.12119
R77 VTAIL VTAIL.n15 1.063
R78 VTAIL.n11 VTAIL.n10 0.470328
R79 VTAIL.n3 VTAIL.n2 0.470328
R80 VTAIL VTAIL.n1 0.0586897
R81 VDD1 VDD1.n0 93.5136
R82 VDD1.n3 VDD1.n2 93.3998
R83 VDD1.n3 VDD1.n1 93.3998
R84 VDD1.n5 VDD1.n4 92.8949
R85 VDD1.n5 VDD1.n3 34.1259
R86 VDD1.n4 VDD1.t4 5.85726
R87 VDD1.n4 VDD1.t2 5.85726
R88 VDD1.n0 VDD1.t3 5.85726
R89 VDD1.n0 VDD1.t5 5.85726
R90 VDD1.n2 VDD1.t1 5.85726
R91 VDD1.n2 VDD1.t7 5.85726
R92 VDD1.n1 VDD1.t0 5.85726
R93 VDD1.n1 VDD1.t6 5.85726
R94 VDD1 VDD1.n5 0.502655
R95 B.n326 B.n325 585
R96 B.n327 B.n46 585
R97 B.n329 B.n328 585
R98 B.n330 B.n45 585
R99 B.n332 B.n331 585
R100 B.n333 B.n44 585
R101 B.n335 B.n334 585
R102 B.n336 B.n43 585
R103 B.n338 B.n337 585
R104 B.n339 B.n42 585
R105 B.n341 B.n340 585
R106 B.n342 B.n41 585
R107 B.n344 B.n343 585
R108 B.n345 B.n40 585
R109 B.n347 B.n346 585
R110 B.n348 B.n39 585
R111 B.n350 B.n349 585
R112 B.n351 B.n38 585
R113 B.n353 B.n352 585
R114 B.n354 B.n37 585
R115 B.n356 B.n355 585
R116 B.n357 B.n36 585
R117 B.n359 B.n358 585
R118 B.n361 B.n33 585
R119 B.n363 B.n362 585
R120 B.n364 B.n32 585
R121 B.n366 B.n365 585
R122 B.n367 B.n31 585
R123 B.n369 B.n368 585
R124 B.n370 B.n30 585
R125 B.n372 B.n371 585
R126 B.n373 B.n27 585
R127 B.n376 B.n375 585
R128 B.n377 B.n26 585
R129 B.n379 B.n378 585
R130 B.n380 B.n25 585
R131 B.n382 B.n381 585
R132 B.n383 B.n24 585
R133 B.n385 B.n384 585
R134 B.n386 B.n23 585
R135 B.n388 B.n387 585
R136 B.n389 B.n22 585
R137 B.n391 B.n390 585
R138 B.n392 B.n21 585
R139 B.n394 B.n393 585
R140 B.n395 B.n20 585
R141 B.n397 B.n396 585
R142 B.n398 B.n19 585
R143 B.n400 B.n399 585
R144 B.n401 B.n18 585
R145 B.n403 B.n402 585
R146 B.n404 B.n17 585
R147 B.n406 B.n405 585
R148 B.n407 B.n16 585
R149 B.n409 B.n408 585
R150 B.n324 B.n47 585
R151 B.n323 B.n322 585
R152 B.n321 B.n48 585
R153 B.n320 B.n319 585
R154 B.n318 B.n49 585
R155 B.n317 B.n316 585
R156 B.n315 B.n50 585
R157 B.n314 B.n313 585
R158 B.n312 B.n51 585
R159 B.n311 B.n310 585
R160 B.n309 B.n52 585
R161 B.n308 B.n307 585
R162 B.n306 B.n53 585
R163 B.n305 B.n304 585
R164 B.n303 B.n54 585
R165 B.n302 B.n301 585
R166 B.n300 B.n55 585
R167 B.n299 B.n298 585
R168 B.n297 B.n56 585
R169 B.n296 B.n295 585
R170 B.n294 B.n57 585
R171 B.n293 B.n292 585
R172 B.n291 B.n58 585
R173 B.n290 B.n289 585
R174 B.n288 B.n59 585
R175 B.n287 B.n286 585
R176 B.n285 B.n60 585
R177 B.n284 B.n283 585
R178 B.n282 B.n61 585
R179 B.n281 B.n280 585
R180 B.n279 B.n62 585
R181 B.n278 B.n277 585
R182 B.n276 B.n63 585
R183 B.n275 B.n274 585
R184 B.n273 B.n64 585
R185 B.n272 B.n271 585
R186 B.n270 B.n65 585
R187 B.n269 B.n268 585
R188 B.n267 B.n66 585
R189 B.n266 B.n265 585
R190 B.n264 B.n67 585
R191 B.n263 B.n262 585
R192 B.n261 B.n68 585
R193 B.n260 B.n259 585
R194 B.n258 B.n69 585
R195 B.n257 B.n256 585
R196 B.n255 B.n70 585
R197 B.n254 B.n253 585
R198 B.n252 B.n71 585
R199 B.n251 B.n250 585
R200 B.n249 B.n72 585
R201 B.n248 B.n247 585
R202 B.n246 B.n73 585
R203 B.n245 B.n244 585
R204 B.n243 B.n74 585
R205 B.n159 B.n106 585
R206 B.n161 B.n160 585
R207 B.n162 B.n105 585
R208 B.n164 B.n163 585
R209 B.n165 B.n104 585
R210 B.n167 B.n166 585
R211 B.n168 B.n103 585
R212 B.n170 B.n169 585
R213 B.n171 B.n102 585
R214 B.n173 B.n172 585
R215 B.n174 B.n101 585
R216 B.n176 B.n175 585
R217 B.n177 B.n100 585
R218 B.n179 B.n178 585
R219 B.n180 B.n99 585
R220 B.n182 B.n181 585
R221 B.n183 B.n98 585
R222 B.n185 B.n184 585
R223 B.n186 B.n97 585
R224 B.n188 B.n187 585
R225 B.n189 B.n96 585
R226 B.n191 B.n190 585
R227 B.n192 B.n93 585
R228 B.n195 B.n194 585
R229 B.n196 B.n92 585
R230 B.n198 B.n197 585
R231 B.n199 B.n91 585
R232 B.n201 B.n200 585
R233 B.n202 B.n90 585
R234 B.n204 B.n203 585
R235 B.n205 B.n89 585
R236 B.n207 B.n206 585
R237 B.n209 B.n208 585
R238 B.n210 B.n85 585
R239 B.n212 B.n211 585
R240 B.n213 B.n84 585
R241 B.n215 B.n214 585
R242 B.n216 B.n83 585
R243 B.n218 B.n217 585
R244 B.n219 B.n82 585
R245 B.n221 B.n220 585
R246 B.n222 B.n81 585
R247 B.n224 B.n223 585
R248 B.n225 B.n80 585
R249 B.n227 B.n226 585
R250 B.n228 B.n79 585
R251 B.n230 B.n229 585
R252 B.n231 B.n78 585
R253 B.n233 B.n232 585
R254 B.n234 B.n77 585
R255 B.n236 B.n235 585
R256 B.n237 B.n76 585
R257 B.n239 B.n238 585
R258 B.n240 B.n75 585
R259 B.n242 B.n241 585
R260 B.n158 B.n157 585
R261 B.n156 B.n107 585
R262 B.n155 B.n154 585
R263 B.n153 B.n108 585
R264 B.n152 B.n151 585
R265 B.n150 B.n109 585
R266 B.n149 B.n148 585
R267 B.n147 B.n110 585
R268 B.n146 B.n145 585
R269 B.n144 B.n111 585
R270 B.n143 B.n142 585
R271 B.n141 B.n112 585
R272 B.n140 B.n139 585
R273 B.n138 B.n113 585
R274 B.n137 B.n136 585
R275 B.n135 B.n114 585
R276 B.n134 B.n133 585
R277 B.n132 B.n115 585
R278 B.n131 B.n130 585
R279 B.n129 B.n116 585
R280 B.n128 B.n127 585
R281 B.n126 B.n117 585
R282 B.n125 B.n124 585
R283 B.n123 B.n118 585
R284 B.n122 B.n121 585
R285 B.n120 B.n119 585
R286 B.n2 B.n0 585
R287 B.n449 B.n1 585
R288 B.n448 B.n447 585
R289 B.n446 B.n3 585
R290 B.n445 B.n444 585
R291 B.n443 B.n4 585
R292 B.n442 B.n441 585
R293 B.n440 B.n5 585
R294 B.n439 B.n438 585
R295 B.n437 B.n6 585
R296 B.n436 B.n435 585
R297 B.n434 B.n7 585
R298 B.n433 B.n432 585
R299 B.n431 B.n8 585
R300 B.n430 B.n429 585
R301 B.n428 B.n9 585
R302 B.n427 B.n426 585
R303 B.n425 B.n10 585
R304 B.n424 B.n423 585
R305 B.n422 B.n11 585
R306 B.n421 B.n420 585
R307 B.n419 B.n12 585
R308 B.n418 B.n417 585
R309 B.n416 B.n13 585
R310 B.n415 B.n414 585
R311 B.n413 B.n14 585
R312 B.n412 B.n411 585
R313 B.n410 B.n15 585
R314 B.n451 B.n450 585
R315 B.n159 B.n158 526.135
R316 B.n408 B.n15 526.135
R317 B.n243 B.n242 526.135
R318 B.n326 B.n47 526.135
R319 B.n86 B.t0 340.611
R320 B.n94 B.t3 340.611
R321 B.n28 B.t9 340.611
R322 B.n34 B.t6 340.611
R323 B.n158 B.n107 163.367
R324 B.n154 B.n107 163.367
R325 B.n154 B.n153 163.367
R326 B.n153 B.n152 163.367
R327 B.n152 B.n109 163.367
R328 B.n148 B.n109 163.367
R329 B.n148 B.n147 163.367
R330 B.n147 B.n146 163.367
R331 B.n146 B.n111 163.367
R332 B.n142 B.n111 163.367
R333 B.n142 B.n141 163.367
R334 B.n141 B.n140 163.367
R335 B.n140 B.n113 163.367
R336 B.n136 B.n113 163.367
R337 B.n136 B.n135 163.367
R338 B.n135 B.n134 163.367
R339 B.n134 B.n115 163.367
R340 B.n130 B.n115 163.367
R341 B.n130 B.n129 163.367
R342 B.n129 B.n128 163.367
R343 B.n128 B.n117 163.367
R344 B.n124 B.n117 163.367
R345 B.n124 B.n123 163.367
R346 B.n123 B.n122 163.367
R347 B.n122 B.n119 163.367
R348 B.n119 B.n2 163.367
R349 B.n450 B.n2 163.367
R350 B.n450 B.n449 163.367
R351 B.n449 B.n448 163.367
R352 B.n448 B.n3 163.367
R353 B.n444 B.n3 163.367
R354 B.n444 B.n443 163.367
R355 B.n443 B.n442 163.367
R356 B.n442 B.n5 163.367
R357 B.n438 B.n5 163.367
R358 B.n438 B.n437 163.367
R359 B.n437 B.n436 163.367
R360 B.n436 B.n7 163.367
R361 B.n432 B.n7 163.367
R362 B.n432 B.n431 163.367
R363 B.n431 B.n430 163.367
R364 B.n430 B.n9 163.367
R365 B.n426 B.n9 163.367
R366 B.n426 B.n425 163.367
R367 B.n425 B.n424 163.367
R368 B.n424 B.n11 163.367
R369 B.n420 B.n11 163.367
R370 B.n420 B.n419 163.367
R371 B.n419 B.n418 163.367
R372 B.n418 B.n13 163.367
R373 B.n414 B.n13 163.367
R374 B.n414 B.n413 163.367
R375 B.n413 B.n412 163.367
R376 B.n412 B.n15 163.367
R377 B.n160 B.n159 163.367
R378 B.n160 B.n105 163.367
R379 B.n164 B.n105 163.367
R380 B.n165 B.n164 163.367
R381 B.n166 B.n165 163.367
R382 B.n166 B.n103 163.367
R383 B.n170 B.n103 163.367
R384 B.n171 B.n170 163.367
R385 B.n172 B.n171 163.367
R386 B.n172 B.n101 163.367
R387 B.n176 B.n101 163.367
R388 B.n177 B.n176 163.367
R389 B.n178 B.n177 163.367
R390 B.n178 B.n99 163.367
R391 B.n182 B.n99 163.367
R392 B.n183 B.n182 163.367
R393 B.n184 B.n183 163.367
R394 B.n184 B.n97 163.367
R395 B.n188 B.n97 163.367
R396 B.n189 B.n188 163.367
R397 B.n190 B.n189 163.367
R398 B.n190 B.n93 163.367
R399 B.n195 B.n93 163.367
R400 B.n196 B.n195 163.367
R401 B.n197 B.n196 163.367
R402 B.n197 B.n91 163.367
R403 B.n201 B.n91 163.367
R404 B.n202 B.n201 163.367
R405 B.n203 B.n202 163.367
R406 B.n203 B.n89 163.367
R407 B.n207 B.n89 163.367
R408 B.n208 B.n207 163.367
R409 B.n208 B.n85 163.367
R410 B.n212 B.n85 163.367
R411 B.n213 B.n212 163.367
R412 B.n214 B.n213 163.367
R413 B.n214 B.n83 163.367
R414 B.n218 B.n83 163.367
R415 B.n219 B.n218 163.367
R416 B.n220 B.n219 163.367
R417 B.n220 B.n81 163.367
R418 B.n224 B.n81 163.367
R419 B.n225 B.n224 163.367
R420 B.n226 B.n225 163.367
R421 B.n226 B.n79 163.367
R422 B.n230 B.n79 163.367
R423 B.n231 B.n230 163.367
R424 B.n232 B.n231 163.367
R425 B.n232 B.n77 163.367
R426 B.n236 B.n77 163.367
R427 B.n237 B.n236 163.367
R428 B.n238 B.n237 163.367
R429 B.n238 B.n75 163.367
R430 B.n242 B.n75 163.367
R431 B.n244 B.n243 163.367
R432 B.n244 B.n73 163.367
R433 B.n248 B.n73 163.367
R434 B.n249 B.n248 163.367
R435 B.n250 B.n249 163.367
R436 B.n250 B.n71 163.367
R437 B.n254 B.n71 163.367
R438 B.n255 B.n254 163.367
R439 B.n256 B.n255 163.367
R440 B.n256 B.n69 163.367
R441 B.n260 B.n69 163.367
R442 B.n261 B.n260 163.367
R443 B.n262 B.n261 163.367
R444 B.n262 B.n67 163.367
R445 B.n266 B.n67 163.367
R446 B.n267 B.n266 163.367
R447 B.n268 B.n267 163.367
R448 B.n268 B.n65 163.367
R449 B.n272 B.n65 163.367
R450 B.n273 B.n272 163.367
R451 B.n274 B.n273 163.367
R452 B.n274 B.n63 163.367
R453 B.n278 B.n63 163.367
R454 B.n279 B.n278 163.367
R455 B.n280 B.n279 163.367
R456 B.n280 B.n61 163.367
R457 B.n284 B.n61 163.367
R458 B.n285 B.n284 163.367
R459 B.n286 B.n285 163.367
R460 B.n286 B.n59 163.367
R461 B.n290 B.n59 163.367
R462 B.n291 B.n290 163.367
R463 B.n292 B.n291 163.367
R464 B.n292 B.n57 163.367
R465 B.n296 B.n57 163.367
R466 B.n297 B.n296 163.367
R467 B.n298 B.n297 163.367
R468 B.n298 B.n55 163.367
R469 B.n302 B.n55 163.367
R470 B.n303 B.n302 163.367
R471 B.n304 B.n303 163.367
R472 B.n304 B.n53 163.367
R473 B.n308 B.n53 163.367
R474 B.n309 B.n308 163.367
R475 B.n310 B.n309 163.367
R476 B.n310 B.n51 163.367
R477 B.n314 B.n51 163.367
R478 B.n315 B.n314 163.367
R479 B.n316 B.n315 163.367
R480 B.n316 B.n49 163.367
R481 B.n320 B.n49 163.367
R482 B.n321 B.n320 163.367
R483 B.n322 B.n321 163.367
R484 B.n322 B.n47 163.367
R485 B.n408 B.n407 163.367
R486 B.n407 B.n406 163.367
R487 B.n406 B.n17 163.367
R488 B.n402 B.n17 163.367
R489 B.n402 B.n401 163.367
R490 B.n401 B.n400 163.367
R491 B.n400 B.n19 163.367
R492 B.n396 B.n19 163.367
R493 B.n396 B.n395 163.367
R494 B.n395 B.n394 163.367
R495 B.n394 B.n21 163.367
R496 B.n390 B.n21 163.367
R497 B.n390 B.n389 163.367
R498 B.n389 B.n388 163.367
R499 B.n388 B.n23 163.367
R500 B.n384 B.n23 163.367
R501 B.n384 B.n383 163.367
R502 B.n383 B.n382 163.367
R503 B.n382 B.n25 163.367
R504 B.n378 B.n25 163.367
R505 B.n378 B.n377 163.367
R506 B.n377 B.n376 163.367
R507 B.n376 B.n27 163.367
R508 B.n371 B.n27 163.367
R509 B.n371 B.n370 163.367
R510 B.n370 B.n369 163.367
R511 B.n369 B.n31 163.367
R512 B.n365 B.n31 163.367
R513 B.n365 B.n364 163.367
R514 B.n364 B.n363 163.367
R515 B.n363 B.n33 163.367
R516 B.n358 B.n33 163.367
R517 B.n358 B.n357 163.367
R518 B.n357 B.n356 163.367
R519 B.n356 B.n37 163.367
R520 B.n352 B.n37 163.367
R521 B.n352 B.n351 163.367
R522 B.n351 B.n350 163.367
R523 B.n350 B.n39 163.367
R524 B.n346 B.n39 163.367
R525 B.n346 B.n345 163.367
R526 B.n345 B.n344 163.367
R527 B.n344 B.n41 163.367
R528 B.n340 B.n41 163.367
R529 B.n340 B.n339 163.367
R530 B.n339 B.n338 163.367
R531 B.n338 B.n43 163.367
R532 B.n334 B.n43 163.367
R533 B.n334 B.n333 163.367
R534 B.n333 B.n332 163.367
R535 B.n332 B.n45 163.367
R536 B.n328 B.n45 163.367
R537 B.n328 B.n327 163.367
R538 B.n327 B.n326 163.367
R539 B.n86 B.t2 139.561
R540 B.n34 B.t7 139.561
R541 B.n94 B.t5 139.555
R542 B.n28 B.t10 139.555
R543 B.n87 B.t1 114.35
R544 B.n35 B.t8 114.35
R545 B.n95 B.t4 114.344
R546 B.n29 B.t11 114.344
R547 B.n88 B.n87 59.5399
R548 B.n193 B.n95 59.5399
R549 B.n374 B.n29 59.5399
R550 B.n360 B.n35 59.5399
R551 B.n410 B.n409 34.1859
R552 B.n325 B.n324 34.1859
R553 B.n241 B.n74 34.1859
R554 B.n157 B.n106 34.1859
R555 B.n87 B.n86 25.2126
R556 B.n95 B.n94 25.2126
R557 B.n29 B.n28 25.2126
R558 B.n35 B.n34 25.2126
R559 B B.n451 18.0485
R560 B.n409 B.n16 10.6151
R561 B.n405 B.n16 10.6151
R562 B.n405 B.n404 10.6151
R563 B.n404 B.n403 10.6151
R564 B.n403 B.n18 10.6151
R565 B.n399 B.n18 10.6151
R566 B.n399 B.n398 10.6151
R567 B.n398 B.n397 10.6151
R568 B.n397 B.n20 10.6151
R569 B.n393 B.n20 10.6151
R570 B.n393 B.n392 10.6151
R571 B.n392 B.n391 10.6151
R572 B.n391 B.n22 10.6151
R573 B.n387 B.n22 10.6151
R574 B.n387 B.n386 10.6151
R575 B.n386 B.n385 10.6151
R576 B.n385 B.n24 10.6151
R577 B.n381 B.n24 10.6151
R578 B.n381 B.n380 10.6151
R579 B.n380 B.n379 10.6151
R580 B.n379 B.n26 10.6151
R581 B.n375 B.n26 10.6151
R582 B.n373 B.n372 10.6151
R583 B.n372 B.n30 10.6151
R584 B.n368 B.n30 10.6151
R585 B.n368 B.n367 10.6151
R586 B.n367 B.n366 10.6151
R587 B.n366 B.n32 10.6151
R588 B.n362 B.n32 10.6151
R589 B.n362 B.n361 10.6151
R590 B.n359 B.n36 10.6151
R591 B.n355 B.n36 10.6151
R592 B.n355 B.n354 10.6151
R593 B.n354 B.n353 10.6151
R594 B.n353 B.n38 10.6151
R595 B.n349 B.n38 10.6151
R596 B.n349 B.n348 10.6151
R597 B.n348 B.n347 10.6151
R598 B.n347 B.n40 10.6151
R599 B.n343 B.n40 10.6151
R600 B.n343 B.n342 10.6151
R601 B.n342 B.n341 10.6151
R602 B.n341 B.n42 10.6151
R603 B.n337 B.n42 10.6151
R604 B.n337 B.n336 10.6151
R605 B.n336 B.n335 10.6151
R606 B.n335 B.n44 10.6151
R607 B.n331 B.n44 10.6151
R608 B.n331 B.n330 10.6151
R609 B.n330 B.n329 10.6151
R610 B.n329 B.n46 10.6151
R611 B.n325 B.n46 10.6151
R612 B.n245 B.n74 10.6151
R613 B.n246 B.n245 10.6151
R614 B.n247 B.n246 10.6151
R615 B.n247 B.n72 10.6151
R616 B.n251 B.n72 10.6151
R617 B.n252 B.n251 10.6151
R618 B.n253 B.n252 10.6151
R619 B.n253 B.n70 10.6151
R620 B.n257 B.n70 10.6151
R621 B.n258 B.n257 10.6151
R622 B.n259 B.n258 10.6151
R623 B.n259 B.n68 10.6151
R624 B.n263 B.n68 10.6151
R625 B.n264 B.n263 10.6151
R626 B.n265 B.n264 10.6151
R627 B.n265 B.n66 10.6151
R628 B.n269 B.n66 10.6151
R629 B.n270 B.n269 10.6151
R630 B.n271 B.n270 10.6151
R631 B.n271 B.n64 10.6151
R632 B.n275 B.n64 10.6151
R633 B.n276 B.n275 10.6151
R634 B.n277 B.n276 10.6151
R635 B.n277 B.n62 10.6151
R636 B.n281 B.n62 10.6151
R637 B.n282 B.n281 10.6151
R638 B.n283 B.n282 10.6151
R639 B.n283 B.n60 10.6151
R640 B.n287 B.n60 10.6151
R641 B.n288 B.n287 10.6151
R642 B.n289 B.n288 10.6151
R643 B.n289 B.n58 10.6151
R644 B.n293 B.n58 10.6151
R645 B.n294 B.n293 10.6151
R646 B.n295 B.n294 10.6151
R647 B.n295 B.n56 10.6151
R648 B.n299 B.n56 10.6151
R649 B.n300 B.n299 10.6151
R650 B.n301 B.n300 10.6151
R651 B.n301 B.n54 10.6151
R652 B.n305 B.n54 10.6151
R653 B.n306 B.n305 10.6151
R654 B.n307 B.n306 10.6151
R655 B.n307 B.n52 10.6151
R656 B.n311 B.n52 10.6151
R657 B.n312 B.n311 10.6151
R658 B.n313 B.n312 10.6151
R659 B.n313 B.n50 10.6151
R660 B.n317 B.n50 10.6151
R661 B.n318 B.n317 10.6151
R662 B.n319 B.n318 10.6151
R663 B.n319 B.n48 10.6151
R664 B.n323 B.n48 10.6151
R665 B.n324 B.n323 10.6151
R666 B.n161 B.n106 10.6151
R667 B.n162 B.n161 10.6151
R668 B.n163 B.n162 10.6151
R669 B.n163 B.n104 10.6151
R670 B.n167 B.n104 10.6151
R671 B.n168 B.n167 10.6151
R672 B.n169 B.n168 10.6151
R673 B.n169 B.n102 10.6151
R674 B.n173 B.n102 10.6151
R675 B.n174 B.n173 10.6151
R676 B.n175 B.n174 10.6151
R677 B.n175 B.n100 10.6151
R678 B.n179 B.n100 10.6151
R679 B.n180 B.n179 10.6151
R680 B.n181 B.n180 10.6151
R681 B.n181 B.n98 10.6151
R682 B.n185 B.n98 10.6151
R683 B.n186 B.n185 10.6151
R684 B.n187 B.n186 10.6151
R685 B.n187 B.n96 10.6151
R686 B.n191 B.n96 10.6151
R687 B.n192 B.n191 10.6151
R688 B.n194 B.n92 10.6151
R689 B.n198 B.n92 10.6151
R690 B.n199 B.n198 10.6151
R691 B.n200 B.n199 10.6151
R692 B.n200 B.n90 10.6151
R693 B.n204 B.n90 10.6151
R694 B.n205 B.n204 10.6151
R695 B.n206 B.n205 10.6151
R696 B.n210 B.n209 10.6151
R697 B.n211 B.n210 10.6151
R698 B.n211 B.n84 10.6151
R699 B.n215 B.n84 10.6151
R700 B.n216 B.n215 10.6151
R701 B.n217 B.n216 10.6151
R702 B.n217 B.n82 10.6151
R703 B.n221 B.n82 10.6151
R704 B.n222 B.n221 10.6151
R705 B.n223 B.n222 10.6151
R706 B.n223 B.n80 10.6151
R707 B.n227 B.n80 10.6151
R708 B.n228 B.n227 10.6151
R709 B.n229 B.n228 10.6151
R710 B.n229 B.n78 10.6151
R711 B.n233 B.n78 10.6151
R712 B.n234 B.n233 10.6151
R713 B.n235 B.n234 10.6151
R714 B.n235 B.n76 10.6151
R715 B.n239 B.n76 10.6151
R716 B.n240 B.n239 10.6151
R717 B.n241 B.n240 10.6151
R718 B.n157 B.n156 10.6151
R719 B.n156 B.n155 10.6151
R720 B.n155 B.n108 10.6151
R721 B.n151 B.n108 10.6151
R722 B.n151 B.n150 10.6151
R723 B.n150 B.n149 10.6151
R724 B.n149 B.n110 10.6151
R725 B.n145 B.n110 10.6151
R726 B.n145 B.n144 10.6151
R727 B.n144 B.n143 10.6151
R728 B.n143 B.n112 10.6151
R729 B.n139 B.n112 10.6151
R730 B.n139 B.n138 10.6151
R731 B.n138 B.n137 10.6151
R732 B.n137 B.n114 10.6151
R733 B.n133 B.n114 10.6151
R734 B.n133 B.n132 10.6151
R735 B.n132 B.n131 10.6151
R736 B.n131 B.n116 10.6151
R737 B.n127 B.n116 10.6151
R738 B.n127 B.n126 10.6151
R739 B.n126 B.n125 10.6151
R740 B.n125 B.n118 10.6151
R741 B.n121 B.n118 10.6151
R742 B.n121 B.n120 10.6151
R743 B.n120 B.n0 10.6151
R744 B.n447 B.n1 10.6151
R745 B.n447 B.n446 10.6151
R746 B.n446 B.n445 10.6151
R747 B.n445 B.n4 10.6151
R748 B.n441 B.n4 10.6151
R749 B.n441 B.n440 10.6151
R750 B.n440 B.n439 10.6151
R751 B.n439 B.n6 10.6151
R752 B.n435 B.n6 10.6151
R753 B.n435 B.n434 10.6151
R754 B.n434 B.n433 10.6151
R755 B.n433 B.n8 10.6151
R756 B.n429 B.n8 10.6151
R757 B.n429 B.n428 10.6151
R758 B.n428 B.n427 10.6151
R759 B.n427 B.n10 10.6151
R760 B.n423 B.n10 10.6151
R761 B.n423 B.n422 10.6151
R762 B.n422 B.n421 10.6151
R763 B.n421 B.n12 10.6151
R764 B.n417 B.n12 10.6151
R765 B.n417 B.n416 10.6151
R766 B.n416 B.n415 10.6151
R767 B.n415 B.n14 10.6151
R768 B.n411 B.n14 10.6151
R769 B.n411 B.n410 10.6151
R770 B.n374 B.n373 6.5566
R771 B.n361 B.n360 6.5566
R772 B.n194 B.n193 6.5566
R773 B.n206 B.n88 6.5566
R774 B.n375 B.n374 4.05904
R775 B.n360 B.n359 4.05904
R776 B.n193 B.n192 4.05904
R777 B.n209 B.n88 4.05904
R778 B.n451 B.n0 2.81026
R779 B.n451 B.n1 2.81026
R780 VN.n2 VN.t0 193.565
R781 VN.n15 VN.t2 193.565
R782 VN.n11 VN.t7 178.638
R783 VN.n24 VN.t5 178.638
R784 VN.n23 VN.n13 161.3
R785 VN.n21 VN.n20 161.3
R786 VN.n19 VN.n14 161.3
R787 VN.n18 VN.n17 161.3
R788 VN.n10 VN.n0 161.3
R789 VN.n8 VN.n7 161.3
R790 VN.n6 VN.n1 161.3
R791 VN.n5 VN.n4 161.3
R792 VN.n3 VN.t6 137.893
R793 VN.n9 VN.t1 137.893
R794 VN.n16 VN.t4 137.893
R795 VN.n22 VN.t3 137.893
R796 VN.n25 VN.n24 80.6037
R797 VN.n12 VN.n11 80.6037
R798 VN.n11 VN.n10 54.8066
R799 VN.n24 VN.n23 54.8066
R800 VN.n3 VN.n2 46.8936
R801 VN.n16 VN.n15 46.8936
R802 VN.n18 VN.n15 44.1212
R803 VN.n5 VN.n2 44.1212
R804 VN.n4 VN.n1 40.4934
R805 VN.n8 VN.n1 40.4934
R806 VN.n17 VN.n14 40.4934
R807 VN.n21 VN.n14 40.4934
R808 VN VN.n25 38.84
R809 VN.n10 VN.n9 17.1274
R810 VN.n23 VN.n22 17.1274
R811 VN.n4 VN.n3 7.3406
R812 VN.n9 VN.n8 7.3406
R813 VN.n17 VN.n16 7.3406
R814 VN.n22 VN.n21 7.3406
R815 VN.n25 VN.n13 0.285035
R816 VN.n12 VN.n0 0.285035
R817 VN.n20 VN.n13 0.189894
R818 VN.n20 VN.n19 0.189894
R819 VN.n19 VN.n18 0.189894
R820 VN.n6 VN.n5 0.189894
R821 VN.n7 VN.n6 0.189894
R822 VN.n7 VN.n0 0.189894
R823 VN VN.n12 0.146778
R824 VDD2.n2 VDD2.n1 93.3998
R825 VDD2.n2 VDD2.n0 93.3998
R826 VDD2 VDD2.n5 93.397
R827 VDD2.n4 VDD2.n3 92.8951
R828 VDD2.n4 VDD2.n2 33.5429
R829 VDD2.n5 VDD2.t3 5.85726
R830 VDD2.n5 VDD2.t5 5.85726
R831 VDD2.n3 VDD2.t2 5.85726
R832 VDD2.n3 VDD2.t4 5.85726
R833 VDD2.n1 VDD2.t6 5.85726
R834 VDD2.n1 VDD2.t0 5.85726
R835 VDD2.n0 VDD2.t7 5.85726
R836 VDD2.n0 VDD2.t1 5.85726
R837 VDD2 VDD2.n4 0.619035
C0 VN VP 4.47467f
C1 VDD2 VDD1 0.961138f
C2 VN B 0.765986f
C3 VTAIL VDD2 5.80205f
C4 VP VDD2 0.346273f
C5 VN w_n2270_n2078# 4.04411f
C6 VDD2 B 1.02391f
C7 VTAIL VDD1 5.75856f
C8 VP VDD1 3.38116f
C9 VDD1 B 0.978771f
C10 VDD2 w_n2270_n2078# 1.27669f
C11 VTAIL VP 3.40675f
C12 VTAIL B 2.22378f
C13 VDD1 w_n2270_n2078# 1.2308f
C14 VP B 1.24325f
C15 VN VDD2 3.18429f
C16 VTAIL w_n2270_n2078# 2.57517f
C17 VP w_n2270_n2078# 4.334f
C18 VN VDD1 0.148833f
C19 w_n2270_n2078# B 5.81681f
C20 VTAIL VN 3.39264f
C21 VDD2 VSUBS 1.143521f
C22 VDD1 VSUBS 1.503229f
C23 VTAIL VSUBS 0.542784f
C24 VN VSUBS 4.47736f
C25 VP VSUBS 1.614631f
C26 B VSUBS 2.561316f
C27 w_n2270_n2078# VSUBS 58.9746f
C28 VDD2.t7 VSUBS 0.11288f
C29 VDD2.t1 VSUBS 0.11288f
C30 VDD2.n0 VSUBS 0.732229f
C31 VDD2.t6 VSUBS 0.11288f
C32 VDD2.t0 VSUBS 0.11288f
C33 VDD2.n1 VSUBS 0.732229f
C34 VDD2.n2 VSUBS 2.39636f
C35 VDD2.t2 VSUBS 0.11288f
C36 VDD2.t4 VSUBS 0.11288f
C37 VDD2.n3 VSUBS 0.729222f
C38 VDD2.n4 VSUBS 2.12946f
C39 VDD2.t3 VSUBS 0.11288f
C40 VDD2.t5 VSUBS 0.11288f
C41 VDD2.n5 VSUBS 0.732204f
C42 VN.n0 VSUBS 0.073392f
C43 VN.t1 VSUBS 0.779968f
C44 VN.n1 VSUBS 0.044463f
C45 VN.t0 VSUBS 0.893195f
C46 VN.n2 VSUBS 0.404015f
C47 VN.t6 VSUBS 0.779968f
C48 VN.n3 VSUBS 0.373064f
C49 VN.n4 VSUBS 0.073888f
C50 VN.n5 VSUBS 0.231424f
C51 VN.n6 VSUBS 0.055001f
C52 VN.n7 VSUBS 0.055001f
C53 VN.n8 VSUBS 0.073888f
C54 VN.n9 VSUBS 0.327211f
C55 VN.n10 VSUBS 0.072235f
C56 VN.t7 VSUBS 0.861703f
C57 VN.n11 VSUBS 0.407997f
C58 VN.n12 VSUBS 0.051511f
C59 VN.n13 VSUBS 0.073392f
C60 VN.t3 VSUBS 0.779968f
C61 VN.n14 VSUBS 0.044463f
C62 VN.t2 VSUBS 0.893195f
C63 VN.n15 VSUBS 0.404015f
C64 VN.t4 VSUBS 0.779968f
C65 VN.n16 VSUBS 0.373064f
C66 VN.n17 VSUBS 0.073888f
C67 VN.n18 VSUBS 0.231424f
C68 VN.n19 VSUBS 0.055001f
C69 VN.n20 VSUBS 0.055001f
C70 VN.n21 VSUBS 0.073888f
C71 VN.n22 VSUBS 0.327211f
C72 VN.n23 VSUBS 0.072235f
C73 VN.t5 VSUBS 0.861703f
C74 VN.n24 VSUBS 0.407997f
C75 VN.n25 VSUBS 2.01063f
C76 B.n0 VSUBS 0.00572f
C77 B.n1 VSUBS 0.00572f
C78 B.n2 VSUBS 0.009045f
C79 B.n3 VSUBS 0.009045f
C80 B.n4 VSUBS 0.009045f
C81 B.n5 VSUBS 0.009045f
C82 B.n6 VSUBS 0.009045f
C83 B.n7 VSUBS 0.009045f
C84 B.n8 VSUBS 0.009045f
C85 B.n9 VSUBS 0.009045f
C86 B.n10 VSUBS 0.009045f
C87 B.n11 VSUBS 0.009045f
C88 B.n12 VSUBS 0.009045f
C89 B.n13 VSUBS 0.009045f
C90 B.n14 VSUBS 0.009045f
C91 B.n15 VSUBS 0.02108f
C92 B.n16 VSUBS 0.009045f
C93 B.n17 VSUBS 0.009045f
C94 B.n18 VSUBS 0.009045f
C95 B.n19 VSUBS 0.009045f
C96 B.n20 VSUBS 0.009045f
C97 B.n21 VSUBS 0.009045f
C98 B.n22 VSUBS 0.009045f
C99 B.n23 VSUBS 0.009045f
C100 B.n24 VSUBS 0.009045f
C101 B.n25 VSUBS 0.009045f
C102 B.n26 VSUBS 0.009045f
C103 B.n27 VSUBS 0.009045f
C104 B.t11 VSUBS 0.205632f
C105 B.t10 VSUBS 0.218188f
C106 B.t9 VSUBS 0.310636f
C107 B.n28 VSUBS 0.116608f
C108 B.n29 VSUBS 0.0824f
C109 B.n30 VSUBS 0.009045f
C110 B.n31 VSUBS 0.009045f
C111 B.n32 VSUBS 0.009045f
C112 B.n33 VSUBS 0.009045f
C113 B.t8 VSUBS 0.205632f
C114 B.t7 VSUBS 0.218187f
C115 B.t6 VSUBS 0.310636f
C116 B.n34 VSUBS 0.116608f
C117 B.n35 VSUBS 0.082401f
C118 B.n36 VSUBS 0.009045f
C119 B.n37 VSUBS 0.009045f
C120 B.n38 VSUBS 0.009045f
C121 B.n39 VSUBS 0.009045f
C122 B.n40 VSUBS 0.009045f
C123 B.n41 VSUBS 0.009045f
C124 B.n42 VSUBS 0.009045f
C125 B.n43 VSUBS 0.009045f
C126 B.n44 VSUBS 0.009045f
C127 B.n45 VSUBS 0.009045f
C128 B.n46 VSUBS 0.009045f
C129 B.n47 VSUBS 0.02108f
C130 B.n48 VSUBS 0.009045f
C131 B.n49 VSUBS 0.009045f
C132 B.n50 VSUBS 0.009045f
C133 B.n51 VSUBS 0.009045f
C134 B.n52 VSUBS 0.009045f
C135 B.n53 VSUBS 0.009045f
C136 B.n54 VSUBS 0.009045f
C137 B.n55 VSUBS 0.009045f
C138 B.n56 VSUBS 0.009045f
C139 B.n57 VSUBS 0.009045f
C140 B.n58 VSUBS 0.009045f
C141 B.n59 VSUBS 0.009045f
C142 B.n60 VSUBS 0.009045f
C143 B.n61 VSUBS 0.009045f
C144 B.n62 VSUBS 0.009045f
C145 B.n63 VSUBS 0.009045f
C146 B.n64 VSUBS 0.009045f
C147 B.n65 VSUBS 0.009045f
C148 B.n66 VSUBS 0.009045f
C149 B.n67 VSUBS 0.009045f
C150 B.n68 VSUBS 0.009045f
C151 B.n69 VSUBS 0.009045f
C152 B.n70 VSUBS 0.009045f
C153 B.n71 VSUBS 0.009045f
C154 B.n72 VSUBS 0.009045f
C155 B.n73 VSUBS 0.009045f
C156 B.n74 VSUBS 0.02108f
C157 B.n75 VSUBS 0.009045f
C158 B.n76 VSUBS 0.009045f
C159 B.n77 VSUBS 0.009045f
C160 B.n78 VSUBS 0.009045f
C161 B.n79 VSUBS 0.009045f
C162 B.n80 VSUBS 0.009045f
C163 B.n81 VSUBS 0.009045f
C164 B.n82 VSUBS 0.009045f
C165 B.n83 VSUBS 0.009045f
C166 B.n84 VSUBS 0.009045f
C167 B.n85 VSUBS 0.009045f
C168 B.t1 VSUBS 0.205632f
C169 B.t2 VSUBS 0.218187f
C170 B.t0 VSUBS 0.310636f
C171 B.n86 VSUBS 0.116608f
C172 B.n87 VSUBS 0.082401f
C173 B.n88 VSUBS 0.020957f
C174 B.n89 VSUBS 0.009045f
C175 B.n90 VSUBS 0.009045f
C176 B.n91 VSUBS 0.009045f
C177 B.n92 VSUBS 0.009045f
C178 B.n93 VSUBS 0.009045f
C179 B.t4 VSUBS 0.205632f
C180 B.t5 VSUBS 0.218188f
C181 B.t3 VSUBS 0.310636f
C182 B.n94 VSUBS 0.116608f
C183 B.n95 VSUBS 0.0824f
C184 B.n96 VSUBS 0.009045f
C185 B.n97 VSUBS 0.009045f
C186 B.n98 VSUBS 0.009045f
C187 B.n99 VSUBS 0.009045f
C188 B.n100 VSUBS 0.009045f
C189 B.n101 VSUBS 0.009045f
C190 B.n102 VSUBS 0.009045f
C191 B.n103 VSUBS 0.009045f
C192 B.n104 VSUBS 0.009045f
C193 B.n105 VSUBS 0.009045f
C194 B.n106 VSUBS 0.022549f
C195 B.n107 VSUBS 0.009045f
C196 B.n108 VSUBS 0.009045f
C197 B.n109 VSUBS 0.009045f
C198 B.n110 VSUBS 0.009045f
C199 B.n111 VSUBS 0.009045f
C200 B.n112 VSUBS 0.009045f
C201 B.n113 VSUBS 0.009045f
C202 B.n114 VSUBS 0.009045f
C203 B.n115 VSUBS 0.009045f
C204 B.n116 VSUBS 0.009045f
C205 B.n117 VSUBS 0.009045f
C206 B.n118 VSUBS 0.009045f
C207 B.n119 VSUBS 0.009045f
C208 B.n120 VSUBS 0.009045f
C209 B.n121 VSUBS 0.009045f
C210 B.n122 VSUBS 0.009045f
C211 B.n123 VSUBS 0.009045f
C212 B.n124 VSUBS 0.009045f
C213 B.n125 VSUBS 0.009045f
C214 B.n126 VSUBS 0.009045f
C215 B.n127 VSUBS 0.009045f
C216 B.n128 VSUBS 0.009045f
C217 B.n129 VSUBS 0.009045f
C218 B.n130 VSUBS 0.009045f
C219 B.n131 VSUBS 0.009045f
C220 B.n132 VSUBS 0.009045f
C221 B.n133 VSUBS 0.009045f
C222 B.n134 VSUBS 0.009045f
C223 B.n135 VSUBS 0.009045f
C224 B.n136 VSUBS 0.009045f
C225 B.n137 VSUBS 0.009045f
C226 B.n138 VSUBS 0.009045f
C227 B.n139 VSUBS 0.009045f
C228 B.n140 VSUBS 0.009045f
C229 B.n141 VSUBS 0.009045f
C230 B.n142 VSUBS 0.009045f
C231 B.n143 VSUBS 0.009045f
C232 B.n144 VSUBS 0.009045f
C233 B.n145 VSUBS 0.009045f
C234 B.n146 VSUBS 0.009045f
C235 B.n147 VSUBS 0.009045f
C236 B.n148 VSUBS 0.009045f
C237 B.n149 VSUBS 0.009045f
C238 B.n150 VSUBS 0.009045f
C239 B.n151 VSUBS 0.009045f
C240 B.n152 VSUBS 0.009045f
C241 B.n153 VSUBS 0.009045f
C242 B.n154 VSUBS 0.009045f
C243 B.n155 VSUBS 0.009045f
C244 B.n156 VSUBS 0.009045f
C245 B.n157 VSUBS 0.02108f
C246 B.n158 VSUBS 0.02108f
C247 B.n159 VSUBS 0.022549f
C248 B.n160 VSUBS 0.009045f
C249 B.n161 VSUBS 0.009045f
C250 B.n162 VSUBS 0.009045f
C251 B.n163 VSUBS 0.009045f
C252 B.n164 VSUBS 0.009045f
C253 B.n165 VSUBS 0.009045f
C254 B.n166 VSUBS 0.009045f
C255 B.n167 VSUBS 0.009045f
C256 B.n168 VSUBS 0.009045f
C257 B.n169 VSUBS 0.009045f
C258 B.n170 VSUBS 0.009045f
C259 B.n171 VSUBS 0.009045f
C260 B.n172 VSUBS 0.009045f
C261 B.n173 VSUBS 0.009045f
C262 B.n174 VSUBS 0.009045f
C263 B.n175 VSUBS 0.009045f
C264 B.n176 VSUBS 0.009045f
C265 B.n177 VSUBS 0.009045f
C266 B.n178 VSUBS 0.009045f
C267 B.n179 VSUBS 0.009045f
C268 B.n180 VSUBS 0.009045f
C269 B.n181 VSUBS 0.009045f
C270 B.n182 VSUBS 0.009045f
C271 B.n183 VSUBS 0.009045f
C272 B.n184 VSUBS 0.009045f
C273 B.n185 VSUBS 0.009045f
C274 B.n186 VSUBS 0.009045f
C275 B.n187 VSUBS 0.009045f
C276 B.n188 VSUBS 0.009045f
C277 B.n189 VSUBS 0.009045f
C278 B.n190 VSUBS 0.009045f
C279 B.n191 VSUBS 0.009045f
C280 B.n192 VSUBS 0.006252f
C281 B.n193 VSUBS 0.020957f
C282 B.n194 VSUBS 0.007316f
C283 B.n195 VSUBS 0.009045f
C284 B.n196 VSUBS 0.009045f
C285 B.n197 VSUBS 0.009045f
C286 B.n198 VSUBS 0.009045f
C287 B.n199 VSUBS 0.009045f
C288 B.n200 VSUBS 0.009045f
C289 B.n201 VSUBS 0.009045f
C290 B.n202 VSUBS 0.009045f
C291 B.n203 VSUBS 0.009045f
C292 B.n204 VSUBS 0.009045f
C293 B.n205 VSUBS 0.009045f
C294 B.n206 VSUBS 0.007316f
C295 B.n207 VSUBS 0.009045f
C296 B.n208 VSUBS 0.009045f
C297 B.n209 VSUBS 0.006252f
C298 B.n210 VSUBS 0.009045f
C299 B.n211 VSUBS 0.009045f
C300 B.n212 VSUBS 0.009045f
C301 B.n213 VSUBS 0.009045f
C302 B.n214 VSUBS 0.009045f
C303 B.n215 VSUBS 0.009045f
C304 B.n216 VSUBS 0.009045f
C305 B.n217 VSUBS 0.009045f
C306 B.n218 VSUBS 0.009045f
C307 B.n219 VSUBS 0.009045f
C308 B.n220 VSUBS 0.009045f
C309 B.n221 VSUBS 0.009045f
C310 B.n222 VSUBS 0.009045f
C311 B.n223 VSUBS 0.009045f
C312 B.n224 VSUBS 0.009045f
C313 B.n225 VSUBS 0.009045f
C314 B.n226 VSUBS 0.009045f
C315 B.n227 VSUBS 0.009045f
C316 B.n228 VSUBS 0.009045f
C317 B.n229 VSUBS 0.009045f
C318 B.n230 VSUBS 0.009045f
C319 B.n231 VSUBS 0.009045f
C320 B.n232 VSUBS 0.009045f
C321 B.n233 VSUBS 0.009045f
C322 B.n234 VSUBS 0.009045f
C323 B.n235 VSUBS 0.009045f
C324 B.n236 VSUBS 0.009045f
C325 B.n237 VSUBS 0.009045f
C326 B.n238 VSUBS 0.009045f
C327 B.n239 VSUBS 0.009045f
C328 B.n240 VSUBS 0.009045f
C329 B.n241 VSUBS 0.022549f
C330 B.n242 VSUBS 0.022549f
C331 B.n243 VSUBS 0.02108f
C332 B.n244 VSUBS 0.009045f
C333 B.n245 VSUBS 0.009045f
C334 B.n246 VSUBS 0.009045f
C335 B.n247 VSUBS 0.009045f
C336 B.n248 VSUBS 0.009045f
C337 B.n249 VSUBS 0.009045f
C338 B.n250 VSUBS 0.009045f
C339 B.n251 VSUBS 0.009045f
C340 B.n252 VSUBS 0.009045f
C341 B.n253 VSUBS 0.009045f
C342 B.n254 VSUBS 0.009045f
C343 B.n255 VSUBS 0.009045f
C344 B.n256 VSUBS 0.009045f
C345 B.n257 VSUBS 0.009045f
C346 B.n258 VSUBS 0.009045f
C347 B.n259 VSUBS 0.009045f
C348 B.n260 VSUBS 0.009045f
C349 B.n261 VSUBS 0.009045f
C350 B.n262 VSUBS 0.009045f
C351 B.n263 VSUBS 0.009045f
C352 B.n264 VSUBS 0.009045f
C353 B.n265 VSUBS 0.009045f
C354 B.n266 VSUBS 0.009045f
C355 B.n267 VSUBS 0.009045f
C356 B.n268 VSUBS 0.009045f
C357 B.n269 VSUBS 0.009045f
C358 B.n270 VSUBS 0.009045f
C359 B.n271 VSUBS 0.009045f
C360 B.n272 VSUBS 0.009045f
C361 B.n273 VSUBS 0.009045f
C362 B.n274 VSUBS 0.009045f
C363 B.n275 VSUBS 0.009045f
C364 B.n276 VSUBS 0.009045f
C365 B.n277 VSUBS 0.009045f
C366 B.n278 VSUBS 0.009045f
C367 B.n279 VSUBS 0.009045f
C368 B.n280 VSUBS 0.009045f
C369 B.n281 VSUBS 0.009045f
C370 B.n282 VSUBS 0.009045f
C371 B.n283 VSUBS 0.009045f
C372 B.n284 VSUBS 0.009045f
C373 B.n285 VSUBS 0.009045f
C374 B.n286 VSUBS 0.009045f
C375 B.n287 VSUBS 0.009045f
C376 B.n288 VSUBS 0.009045f
C377 B.n289 VSUBS 0.009045f
C378 B.n290 VSUBS 0.009045f
C379 B.n291 VSUBS 0.009045f
C380 B.n292 VSUBS 0.009045f
C381 B.n293 VSUBS 0.009045f
C382 B.n294 VSUBS 0.009045f
C383 B.n295 VSUBS 0.009045f
C384 B.n296 VSUBS 0.009045f
C385 B.n297 VSUBS 0.009045f
C386 B.n298 VSUBS 0.009045f
C387 B.n299 VSUBS 0.009045f
C388 B.n300 VSUBS 0.009045f
C389 B.n301 VSUBS 0.009045f
C390 B.n302 VSUBS 0.009045f
C391 B.n303 VSUBS 0.009045f
C392 B.n304 VSUBS 0.009045f
C393 B.n305 VSUBS 0.009045f
C394 B.n306 VSUBS 0.009045f
C395 B.n307 VSUBS 0.009045f
C396 B.n308 VSUBS 0.009045f
C397 B.n309 VSUBS 0.009045f
C398 B.n310 VSUBS 0.009045f
C399 B.n311 VSUBS 0.009045f
C400 B.n312 VSUBS 0.009045f
C401 B.n313 VSUBS 0.009045f
C402 B.n314 VSUBS 0.009045f
C403 B.n315 VSUBS 0.009045f
C404 B.n316 VSUBS 0.009045f
C405 B.n317 VSUBS 0.009045f
C406 B.n318 VSUBS 0.009045f
C407 B.n319 VSUBS 0.009045f
C408 B.n320 VSUBS 0.009045f
C409 B.n321 VSUBS 0.009045f
C410 B.n322 VSUBS 0.009045f
C411 B.n323 VSUBS 0.009045f
C412 B.n324 VSUBS 0.022101f
C413 B.n325 VSUBS 0.021528f
C414 B.n326 VSUBS 0.022549f
C415 B.n327 VSUBS 0.009045f
C416 B.n328 VSUBS 0.009045f
C417 B.n329 VSUBS 0.009045f
C418 B.n330 VSUBS 0.009045f
C419 B.n331 VSUBS 0.009045f
C420 B.n332 VSUBS 0.009045f
C421 B.n333 VSUBS 0.009045f
C422 B.n334 VSUBS 0.009045f
C423 B.n335 VSUBS 0.009045f
C424 B.n336 VSUBS 0.009045f
C425 B.n337 VSUBS 0.009045f
C426 B.n338 VSUBS 0.009045f
C427 B.n339 VSUBS 0.009045f
C428 B.n340 VSUBS 0.009045f
C429 B.n341 VSUBS 0.009045f
C430 B.n342 VSUBS 0.009045f
C431 B.n343 VSUBS 0.009045f
C432 B.n344 VSUBS 0.009045f
C433 B.n345 VSUBS 0.009045f
C434 B.n346 VSUBS 0.009045f
C435 B.n347 VSUBS 0.009045f
C436 B.n348 VSUBS 0.009045f
C437 B.n349 VSUBS 0.009045f
C438 B.n350 VSUBS 0.009045f
C439 B.n351 VSUBS 0.009045f
C440 B.n352 VSUBS 0.009045f
C441 B.n353 VSUBS 0.009045f
C442 B.n354 VSUBS 0.009045f
C443 B.n355 VSUBS 0.009045f
C444 B.n356 VSUBS 0.009045f
C445 B.n357 VSUBS 0.009045f
C446 B.n358 VSUBS 0.009045f
C447 B.n359 VSUBS 0.006252f
C448 B.n360 VSUBS 0.020957f
C449 B.n361 VSUBS 0.007316f
C450 B.n362 VSUBS 0.009045f
C451 B.n363 VSUBS 0.009045f
C452 B.n364 VSUBS 0.009045f
C453 B.n365 VSUBS 0.009045f
C454 B.n366 VSUBS 0.009045f
C455 B.n367 VSUBS 0.009045f
C456 B.n368 VSUBS 0.009045f
C457 B.n369 VSUBS 0.009045f
C458 B.n370 VSUBS 0.009045f
C459 B.n371 VSUBS 0.009045f
C460 B.n372 VSUBS 0.009045f
C461 B.n373 VSUBS 0.007316f
C462 B.n374 VSUBS 0.020957f
C463 B.n375 VSUBS 0.006252f
C464 B.n376 VSUBS 0.009045f
C465 B.n377 VSUBS 0.009045f
C466 B.n378 VSUBS 0.009045f
C467 B.n379 VSUBS 0.009045f
C468 B.n380 VSUBS 0.009045f
C469 B.n381 VSUBS 0.009045f
C470 B.n382 VSUBS 0.009045f
C471 B.n383 VSUBS 0.009045f
C472 B.n384 VSUBS 0.009045f
C473 B.n385 VSUBS 0.009045f
C474 B.n386 VSUBS 0.009045f
C475 B.n387 VSUBS 0.009045f
C476 B.n388 VSUBS 0.009045f
C477 B.n389 VSUBS 0.009045f
C478 B.n390 VSUBS 0.009045f
C479 B.n391 VSUBS 0.009045f
C480 B.n392 VSUBS 0.009045f
C481 B.n393 VSUBS 0.009045f
C482 B.n394 VSUBS 0.009045f
C483 B.n395 VSUBS 0.009045f
C484 B.n396 VSUBS 0.009045f
C485 B.n397 VSUBS 0.009045f
C486 B.n398 VSUBS 0.009045f
C487 B.n399 VSUBS 0.009045f
C488 B.n400 VSUBS 0.009045f
C489 B.n401 VSUBS 0.009045f
C490 B.n402 VSUBS 0.009045f
C491 B.n403 VSUBS 0.009045f
C492 B.n404 VSUBS 0.009045f
C493 B.n405 VSUBS 0.009045f
C494 B.n406 VSUBS 0.009045f
C495 B.n407 VSUBS 0.009045f
C496 B.n408 VSUBS 0.022549f
C497 B.n409 VSUBS 0.022549f
C498 B.n410 VSUBS 0.02108f
C499 B.n411 VSUBS 0.009045f
C500 B.n412 VSUBS 0.009045f
C501 B.n413 VSUBS 0.009045f
C502 B.n414 VSUBS 0.009045f
C503 B.n415 VSUBS 0.009045f
C504 B.n416 VSUBS 0.009045f
C505 B.n417 VSUBS 0.009045f
C506 B.n418 VSUBS 0.009045f
C507 B.n419 VSUBS 0.009045f
C508 B.n420 VSUBS 0.009045f
C509 B.n421 VSUBS 0.009045f
C510 B.n422 VSUBS 0.009045f
C511 B.n423 VSUBS 0.009045f
C512 B.n424 VSUBS 0.009045f
C513 B.n425 VSUBS 0.009045f
C514 B.n426 VSUBS 0.009045f
C515 B.n427 VSUBS 0.009045f
C516 B.n428 VSUBS 0.009045f
C517 B.n429 VSUBS 0.009045f
C518 B.n430 VSUBS 0.009045f
C519 B.n431 VSUBS 0.009045f
C520 B.n432 VSUBS 0.009045f
C521 B.n433 VSUBS 0.009045f
C522 B.n434 VSUBS 0.009045f
C523 B.n435 VSUBS 0.009045f
C524 B.n436 VSUBS 0.009045f
C525 B.n437 VSUBS 0.009045f
C526 B.n438 VSUBS 0.009045f
C527 B.n439 VSUBS 0.009045f
C528 B.n440 VSUBS 0.009045f
C529 B.n441 VSUBS 0.009045f
C530 B.n442 VSUBS 0.009045f
C531 B.n443 VSUBS 0.009045f
C532 B.n444 VSUBS 0.009045f
C533 B.n445 VSUBS 0.009045f
C534 B.n446 VSUBS 0.009045f
C535 B.n447 VSUBS 0.009045f
C536 B.n448 VSUBS 0.009045f
C537 B.n449 VSUBS 0.009045f
C538 B.n450 VSUBS 0.009045f
C539 B.n451 VSUBS 0.020481f
C540 VDD1.t3 VSUBS 0.114183f
C541 VDD1.t5 VSUBS 0.114183f
C542 VDD1.n0 VSUBS 0.741415f
C543 VDD1.t0 VSUBS 0.114183f
C544 VDD1.t6 VSUBS 0.114183f
C545 VDD1.n1 VSUBS 0.740677f
C546 VDD1.t1 VSUBS 0.114183f
C547 VDD1.t7 VSUBS 0.114183f
C548 VDD1.n2 VSUBS 0.740677f
C549 VDD1.n3 VSUBS 2.47958f
C550 VDD1.t4 VSUBS 0.114183f
C551 VDD1.t2 VSUBS 0.114183f
C552 VDD1.n4 VSUBS 0.737632f
C553 VDD1.n5 VSUBS 2.18485f
C554 VTAIL.t6 VSUBS 0.121123f
C555 VTAIL.t15 VSUBS 0.121123f
C556 VTAIL.n0 VSUBS 0.687262f
C557 VTAIL.n1 VSUBS 0.602885f
C558 VTAIL.t2 VSUBS 0.953624f
C559 VTAIL.n2 VSUBS 0.703489f
C560 VTAIL.t12 VSUBS 0.953624f
C561 VTAIL.n3 VSUBS 0.703489f
C562 VTAIL.t9 VSUBS 0.121123f
C563 VTAIL.t7 VSUBS 0.121123f
C564 VTAIL.n4 VSUBS 0.687262f
C565 VTAIL.n5 VSUBS 0.697435f
C566 VTAIL.t13 VSUBS 0.953624f
C567 VTAIL.n6 VSUBS 1.56232f
C568 VTAIL.t5 VSUBS 0.953628f
C569 VTAIL.n7 VSUBS 1.56232f
C570 VTAIL.t1 VSUBS 0.121123f
C571 VTAIL.t0 VSUBS 0.121123f
C572 VTAIL.n8 VSUBS 0.687266f
C573 VTAIL.n9 VSUBS 0.697431f
C574 VTAIL.t4 VSUBS 0.953628f
C575 VTAIL.n10 VSUBS 0.703485f
C576 VTAIL.t8 VSUBS 0.953628f
C577 VTAIL.n11 VSUBS 0.703485f
C578 VTAIL.t14 VSUBS 0.121123f
C579 VTAIL.t11 VSUBS 0.121123f
C580 VTAIL.n12 VSUBS 0.687266f
C581 VTAIL.n13 VSUBS 0.697431f
C582 VTAIL.t10 VSUBS 0.953624f
C583 VTAIL.n14 VSUBS 1.56232f
C584 VTAIL.t3 VSUBS 0.953624f
C585 VTAIL.n15 VSUBS 1.55714f
C586 VP.n0 VSUBS 0.076213f
C587 VP.t6 VSUBS 0.809942f
C588 VP.n1 VSUBS 0.046172f
C589 VP.n2 VSUBS 0.076213f
C590 VP.t1 VSUBS 0.809942f
C591 VP.n3 VSUBS 0.076213f
C592 VP.t5 VSUBS 0.894818f
C593 VP.t3 VSUBS 0.809942f
C594 VP.n4 VSUBS 0.046172f
C595 VP.t4 VSUBS 0.92752f
C596 VP.n5 VSUBS 0.419541f
C597 VP.t2 VSUBS 0.809942f
C598 VP.n6 VSUBS 0.3874f
C599 VP.n7 VSUBS 0.076728f
C600 VP.n8 VSUBS 0.240318f
C601 VP.n9 VSUBS 0.057115f
C602 VP.n10 VSUBS 0.057115f
C603 VP.n11 VSUBS 0.076728f
C604 VP.n12 VSUBS 0.339786f
C605 VP.n13 VSUBS 0.075011f
C606 VP.n14 VSUBS 0.423676f
C607 VP.n15 VSUBS 2.05535f
C608 VP.n16 VSUBS 2.1086f
C609 VP.t7 VSUBS 0.894818f
C610 VP.n17 VSUBS 0.423676f
C611 VP.n18 VSUBS 0.075011f
C612 VP.n19 VSUBS 0.339786f
C613 VP.n20 VSUBS 0.076728f
C614 VP.n21 VSUBS 0.057115f
C615 VP.n22 VSUBS 0.057115f
C616 VP.n23 VSUBS 0.057115f
C617 VP.n24 VSUBS 0.076728f
C618 VP.n25 VSUBS 0.339786f
C619 VP.n26 VSUBS 0.075011f
C620 VP.t0 VSUBS 0.894818f
C621 VP.n27 VSUBS 0.423676f
C622 VP.n28 VSUBS 0.05349f
.ends

