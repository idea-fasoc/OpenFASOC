* NGSPICE file created from diff_pair_sample_1480.ext - technology: sky130A

.subckt diff_pair_sample_1480 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=1.521 ps=8.58 w=3.9 l=1.26
X1 B.t11 B.t9 B.t10 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=0 ps=0 w=3.9 l=1.26
X2 B.t8 B.t6 B.t7 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=0 ps=0 w=3.9 l=1.26
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=1.521 ps=8.58 w=3.9 l=1.26
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=1.521 ps=8.58 w=3.9 l=1.26
X5 VDD1.t0 VP.t1 VTAIL.t2 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=1.521 ps=8.58 w=3.9 l=1.26
X6 B.t5 B.t3 B.t4 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=0 ps=0 w=3.9 l=1.26
X7 B.t2 B.t0 B.t1 w_n1606_n1748# sky130_fd_pr__pfet_01v8 ad=1.521 pd=8.58 as=0 ps=0 w=3.9 l=1.26
R0 VP.n0 VP.t1 221.343
R1 VP.n0 VP.t0 186.375
R2 VP VP.n0 0.146778
R3 VTAIL.n74 VTAIL.n60 756.745
R4 VTAIL.n14 VTAIL.n0 756.745
R5 VTAIL.n54 VTAIL.n40 756.745
R6 VTAIL.n34 VTAIL.n20 756.745
R7 VTAIL.n67 VTAIL.n66 585
R8 VTAIL.n64 VTAIL.n63 585
R9 VTAIL.n73 VTAIL.n72 585
R10 VTAIL.n75 VTAIL.n74 585
R11 VTAIL.n7 VTAIL.n6 585
R12 VTAIL.n4 VTAIL.n3 585
R13 VTAIL.n13 VTAIL.n12 585
R14 VTAIL.n15 VTAIL.n14 585
R15 VTAIL.n55 VTAIL.n54 585
R16 VTAIL.n53 VTAIL.n52 585
R17 VTAIL.n44 VTAIL.n43 585
R18 VTAIL.n47 VTAIL.n46 585
R19 VTAIL.n35 VTAIL.n34 585
R20 VTAIL.n33 VTAIL.n32 585
R21 VTAIL.n24 VTAIL.n23 585
R22 VTAIL.n27 VTAIL.n26 585
R23 VTAIL.t0 VTAIL.n65 330.707
R24 VTAIL.t3 VTAIL.n5 330.707
R25 VTAIL.t2 VTAIL.n45 330.707
R26 VTAIL.t1 VTAIL.n25 330.707
R27 VTAIL.n66 VTAIL.n63 171.744
R28 VTAIL.n73 VTAIL.n63 171.744
R29 VTAIL.n74 VTAIL.n73 171.744
R30 VTAIL.n6 VTAIL.n3 171.744
R31 VTAIL.n13 VTAIL.n3 171.744
R32 VTAIL.n14 VTAIL.n13 171.744
R33 VTAIL.n54 VTAIL.n53 171.744
R34 VTAIL.n53 VTAIL.n43 171.744
R35 VTAIL.n46 VTAIL.n43 171.744
R36 VTAIL.n34 VTAIL.n33 171.744
R37 VTAIL.n33 VTAIL.n23 171.744
R38 VTAIL.n26 VTAIL.n23 171.744
R39 VTAIL.n66 VTAIL.t0 85.8723
R40 VTAIL.n6 VTAIL.t3 85.8723
R41 VTAIL.n46 VTAIL.t2 85.8723
R42 VTAIL.n26 VTAIL.t1 85.8723
R43 VTAIL.n79 VTAIL.n78 33.349
R44 VTAIL.n19 VTAIL.n18 33.349
R45 VTAIL.n59 VTAIL.n58 33.349
R46 VTAIL.n39 VTAIL.n38 33.349
R47 VTAIL.n39 VTAIL.n19 18.4703
R48 VTAIL.n79 VTAIL.n59 17.0996
R49 VTAIL.n67 VTAIL.n65 16.3201
R50 VTAIL.n7 VTAIL.n5 16.3201
R51 VTAIL.n47 VTAIL.n45 16.3201
R52 VTAIL.n27 VTAIL.n25 16.3201
R53 VTAIL.n68 VTAIL.n64 12.8005
R54 VTAIL.n8 VTAIL.n4 12.8005
R55 VTAIL.n48 VTAIL.n44 12.8005
R56 VTAIL.n28 VTAIL.n24 12.8005
R57 VTAIL.n72 VTAIL.n71 12.0247
R58 VTAIL.n12 VTAIL.n11 12.0247
R59 VTAIL.n52 VTAIL.n51 12.0247
R60 VTAIL.n32 VTAIL.n31 12.0247
R61 VTAIL.n75 VTAIL.n62 11.249
R62 VTAIL.n15 VTAIL.n2 11.249
R63 VTAIL.n55 VTAIL.n42 11.249
R64 VTAIL.n35 VTAIL.n22 11.249
R65 VTAIL.n76 VTAIL.n60 10.4732
R66 VTAIL.n16 VTAIL.n0 10.4732
R67 VTAIL.n56 VTAIL.n40 10.4732
R68 VTAIL.n36 VTAIL.n20 10.4732
R69 VTAIL.n78 VTAIL.n77 9.45567
R70 VTAIL.n18 VTAIL.n17 9.45567
R71 VTAIL.n58 VTAIL.n57 9.45567
R72 VTAIL.n38 VTAIL.n37 9.45567
R73 VTAIL.n77 VTAIL.n76 9.3005
R74 VTAIL.n62 VTAIL.n61 9.3005
R75 VTAIL.n71 VTAIL.n70 9.3005
R76 VTAIL.n69 VTAIL.n68 9.3005
R77 VTAIL.n17 VTAIL.n16 9.3005
R78 VTAIL.n2 VTAIL.n1 9.3005
R79 VTAIL.n11 VTAIL.n10 9.3005
R80 VTAIL.n9 VTAIL.n8 9.3005
R81 VTAIL.n57 VTAIL.n56 9.3005
R82 VTAIL.n42 VTAIL.n41 9.3005
R83 VTAIL.n51 VTAIL.n50 9.3005
R84 VTAIL.n49 VTAIL.n48 9.3005
R85 VTAIL.n37 VTAIL.n36 9.3005
R86 VTAIL.n22 VTAIL.n21 9.3005
R87 VTAIL.n31 VTAIL.n30 9.3005
R88 VTAIL.n29 VTAIL.n28 9.3005
R89 VTAIL.n69 VTAIL.n65 3.78097
R90 VTAIL.n9 VTAIL.n5 3.78097
R91 VTAIL.n49 VTAIL.n45 3.78097
R92 VTAIL.n29 VTAIL.n25 3.78097
R93 VTAIL.n78 VTAIL.n60 3.49141
R94 VTAIL.n18 VTAIL.n0 3.49141
R95 VTAIL.n58 VTAIL.n40 3.49141
R96 VTAIL.n38 VTAIL.n20 3.49141
R97 VTAIL.n76 VTAIL.n75 2.71565
R98 VTAIL.n16 VTAIL.n15 2.71565
R99 VTAIL.n56 VTAIL.n55 2.71565
R100 VTAIL.n36 VTAIL.n35 2.71565
R101 VTAIL.n72 VTAIL.n62 1.93989
R102 VTAIL.n12 VTAIL.n2 1.93989
R103 VTAIL.n52 VTAIL.n42 1.93989
R104 VTAIL.n32 VTAIL.n22 1.93989
R105 VTAIL.n71 VTAIL.n64 1.16414
R106 VTAIL.n11 VTAIL.n4 1.16414
R107 VTAIL.n51 VTAIL.n44 1.16414
R108 VTAIL.n31 VTAIL.n24 1.16414
R109 VTAIL.n59 VTAIL.n39 1.15567
R110 VTAIL VTAIL.n19 0.87119
R111 VTAIL.n68 VTAIL.n67 0.388379
R112 VTAIL.n8 VTAIL.n7 0.388379
R113 VTAIL.n48 VTAIL.n47 0.388379
R114 VTAIL.n28 VTAIL.n27 0.388379
R115 VTAIL VTAIL.n79 0.284983
R116 VTAIL.n70 VTAIL.n69 0.155672
R117 VTAIL.n70 VTAIL.n61 0.155672
R118 VTAIL.n77 VTAIL.n61 0.155672
R119 VTAIL.n10 VTAIL.n9 0.155672
R120 VTAIL.n10 VTAIL.n1 0.155672
R121 VTAIL.n17 VTAIL.n1 0.155672
R122 VTAIL.n57 VTAIL.n41 0.155672
R123 VTAIL.n50 VTAIL.n41 0.155672
R124 VTAIL.n50 VTAIL.n49 0.155672
R125 VTAIL.n37 VTAIL.n21 0.155672
R126 VTAIL.n30 VTAIL.n21 0.155672
R127 VTAIL.n30 VTAIL.n29 0.155672
R128 VDD1.n14 VDD1.n0 756.745
R129 VDD1.n33 VDD1.n19 756.745
R130 VDD1.n15 VDD1.n14 585
R131 VDD1.n13 VDD1.n12 585
R132 VDD1.n4 VDD1.n3 585
R133 VDD1.n7 VDD1.n6 585
R134 VDD1.n26 VDD1.n25 585
R135 VDD1.n23 VDD1.n22 585
R136 VDD1.n32 VDD1.n31 585
R137 VDD1.n34 VDD1.n33 585
R138 VDD1.t0 VDD1.n5 330.707
R139 VDD1.t1 VDD1.n24 330.707
R140 VDD1.n14 VDD1.n13 171.744
R141 VDD1.n13 VDD1.n3 171.744
R142 VDD1.n6 VDD1.n3 171.744
R143 VDD1.n25 VDD1.n22 171.744
R144 VDD1.n32 VDD1.n22 171.744
R145 VDD1.n33 VDD1.n32 171.744
R146 VDD1.n6 VDD1.t0 85.8723
R147 VDD1.n25 VDD1.t1 85.8723
R148 VDD1 VDD1.n37 80.6582
R149 VDD1 VDD1.n18 50.4286
R150 VDD1.n7 VDD1.n5 16.3201
R151 VDD1.n26 VDD1.n24 16.3201
R152 VDD1.n8 VDD1.n4 12.8005
R153 VDD1.n27 VDD1.n23 12.8005
R154 VDD1.n12 VDD1.n11 12.0247
R155 VDD1.n31 VDD1.n30 12.0247
R156 VDD1.n15 VDD1.n2 11.249
R157 VDD1.n34 VDD1.n21 11.249
R158 VDD1.n16 VDD1.n0 10.4732
R159 VDD1.n35 VDD1.n19 10.4732
R160 VDD1.n18 VDD1.n17 9.45567
R161 VDD1.n37 VDD1.n36 9.45567
R162 VDD1.n17 VDD1.n16 9.3005
R163 VDD1.n2 VDD1.n1 9.3005
R164 VDD1.n11 VDD1.n10 9.3005
R165 VDD1.n9 VDD1.n8 9.3005
R166 VDD1.n36 VDD1.n35 9.3005
R167 VDD1.n21 VDD1.n20 9.3005
R168 VDD1.n30 VDD1.n29 9.3005
R169 VDD1.n28 VDD1.n27 9.3005
R170 VDD1.n9 VDD1.n5 3.78097
R171 VDD1.n28 VDD1.n24 3.78097
R172 VDD1.n18 VDD1.n0 3.49141
R173 VDD1.n37 VDD1.n19 3.49141
R174 VDD1.n16 VDD1.n15 2.71565
R175 VDD1.n35 VDD1.n34 2.71565
R176 VDD1.n12 VDD1.n2 1.93989
R177 VDD1.n31 VDD1.n21 1.93989
R178 VDD1.n11 VDD1.n4 1.16414
R179 VDD1.n30 VDD1.n23 1.16414
R180 VDD1.n8 VDD1.n7 0.388379
R181 VDD1.n27 VDD1.n26 0.388379
R182 VDD1.n17 VDD1.n1 0.155672
R183 VDD1.n10 VDD1.n1 0.155672
R184 VDD1.n10 VDD1.n9 0.155672
R185 VDD1.n29 VDD1.n28 0.155672
R186 VDD1.n29 VDD1.n20 0.155672
R187 VDD1.n36 VDD1.n20 0.155672
R188 B.n183 B.n182 585
R189 B.n181 B.n56 585
R190 B.n180 B.n179 585
R191 B.n178 B.n57 585
R192 B.n177 B.n176 585
R193 B.n175 B.n58 585
R194 B.n174 B.n173 585
R195 B.n172 B.n59 585
R196 B.n171 B.n170 585
R197 B.n169 B.n60 585
R198 B.n168 B.n167 585
R199 B.n166 B.n61 585
R200 B.n165 B.n164 585
R201 B.n163 B.n62 585
R202 B.n162 B.n161 585
R203 B.n160 B.n63 585
R204 B.n159 B.n158 585
R205 B.n157 B.n64 585
R206 B.n156 B.n155 585
R207 B.n151 B.n65 585
R208 B.n150 B.n149 585
R209 B.n148 B.n66 585
R210 B.n147 B.n146 585
R211 B.n145 B.n67 585
R212 B.n144 B.n143 585
R213 B.n142 B.n68 585
R214 B.n141 B.n140 585
R215 B.n138 B.n69 585
R216 B.n137 B.n136 585
R217 B.n135 B.n72 585
R218 B.n134 B.n133 585
R219 B.n132 B.n73 585
R220 B.n131 B.n130 585
R221 B.n129 B.n74 585
R222 B.n128 B.n127 585
R223 B.n126 B.n75 585
R224 B.n125 B.n124 585
R225 B.n123 B.n76 585
R226 B.n122 B.n121 585
R227 B.n120 B.n77 585
R228 B.n119 B.n118 585
R229 B.n117 B.n78 585
R230 B.n116 B.n115 585
R231 B.n114 B.n79 585
R232 B.n113 B.n112 585
R233 B.n184 B.n55 585
R234 B.n186 B.n185 585
R235 B.n187 B.n54 585
R236 B.n189 B.n188 585
R237 B.n190 B.n53 585
R238 B.n192 B.n191 585
R239 B.n193 B.n52 585
R240 B.n195 B.n194 585
R241 B.n196 B.n51 585
R242 B.n198 B.n197 585
R243 B.n199 B.n50 585
R244 B.n201 B.n200 585
R245 B.n202 B.n49 585
R246 B.n204 B.n203 585
R247 B.n205 B.n48 585
R248 B.n207 B.n206 585
R249 B.n208 B.n47 585
R250 B.n210 B.n209 585
R251 B.n211 B.n46 585
R252 B.n213 B.n212 585
R253 B.n214 B.n45 585
R254 B.n216 B.n215 585
R255 B.n217 B.n44 585
R256 B.n219 B.n218 585
R257 B.n220 B.n43 585
R258 B.n222 B.n221 585
R259 B.n223 B.n42 585
R260 B.n225 B.n224 585
R261 B.n226 B.n41 585
R262 B.n228 B.n227 585
R263 B.n229 B.n40 585
R264 B.n231 B.n230 585
R265 B.n232 B.n39 585
R266 B.n234 B.n233 585
R267 B.n235 B.n38 585
R268 B.n237 B.n236 585
R269 B.n306 B.n305 585
R270 B.n304 B.n11 585
R271 B.n303 B.n302 585
R272 B.n301 B.n12 585
R273 B.n300 B.n299 585
R274 B.n298 B.n13 585
R275 B.n297 B.n296 585
R276 B.n295 B.n14 585
R277 B.n294 B.n293 585
R278 B.n292 B.n15 585
R279 B.n291 B.n290 585
R280 B.n289 B.n16 585
R281 B.n288 B.n287 585
R282 B.n286 B.n17 585
R283 B.n285 B.n284 585
R284 B.n283 B.n18 585
R285 B.n282 B.n281 585
R286 B.n280 B.n19 585
R287 B.n278 B.n277 585
R288 B.n276 B.n22 585
R289 B.n275 B.n274 585
R290 B.n273 B.n23 585
R291 B.n272 B.n271 585
R292 B.n270 B.n24 585
R293 B.n269 B.n268 585
R294 B.n267 B.n25 585
R295 B.n266 B.n265 585
R296 B.n264 B.n263 585
R297 B.n262 B.n29 585
R298 B.n261 B.n260 585
R299 B.n259 B.n30 585
R300 B.n258 B.n257 585
R301 B.n256 B.n31 585
R302 B.n255 B.n254 585
R303 B.n253 B.n32 585
R304 B.n252 B.n251 585
R305 B.n250 B.n33 585
R306 B.n249 B.n248 585
R307 B.n247 B.n34 585
R308 B.n246 B.n245 585
R309 B.n244 B.n35 585
R310 B.n243 B.n242 585
R311 B.n241 B.n36 585
R312 B.n240 B.n239 585
R313 B.n238 B.n37 585
R314 B.n307 B.n10 585
R315 B.n309 B.n308 585
R316 B.n310 B.n9 585
R317 B.n312 B.n311 585
R318 B.n313 B.n8 585
R319 B.n315 B.n314 585
R320 B.n316 B.n7 585
R321 B.n318 B.n317 585
R322 B.n319 B.n6 585
R323 B.n321 B.n320 585
R324 B.n322 B.n5 585
R325 B.n324 B.n323 585
R326 B.n325 B.n4 585
R327 B.n327 B.n326 585
R328 B.n328 B.n3 585
R329 B.n330 B.n329 585
R330 B.n331 B.n0 585
R331 B.n2 B.n1 585
R332 B.n89 B.n88 585
R333 B.n90 B.n87 585
R334 B.n92 B.n91 585
R335 B.n93 B.n86 585
R336 B.n95 B.n94 585
R337 B.n96 B.n85 585
R338 B.n98 B.n97 585
R339 B.n99 B.n84 585
R340 B.n101 B.n100 585
R341 B.n102 B.n83 585
R342 B.n104 B.n103 585
R343 B.n105 B.n82 585
R344 B.n107 B.n106 585
R345 B.n108 B.n81 585
R346 B.n110 B.n109 585
R347 B.n111 B.n80 585
R348 B.n112 B.n111 506.916
R349 B.n182 B.n55 506.916
R350 B.n236 B.n37 506.916
R351 B.n307 B.n306 506.916
R352 B.n70 B.t0 279.014
R353 B.n152 B.t3 279.014
R354 B.n26 B.t9 279.014
R355 B.n20 B.t6 279.014
R356 B.n152 B.t4 264.526
R357 B.n26 B.t11 264.526
R358 B.n70 B.t1 264.526
R359 B.n20 B.t8 264.526
R360 B.n333 B.n332 256.663
R361 B.n332 B.n331 235.042
R362 B.n332 B.n2 235.042
R363 B.n153 B.t5 233.69
R364 B.n27 B.t10 233.69
R365 B.n71 B.t2 233.69
R366 B.n21 B.t7 233.69
R367 B.n112 B.n79 163.367
R368 B.n116 B.n79 163.367
R369 B.n117 B.n116 163.367
R370 B.n118 B.n117 163.367
R371 B.n118 B.n77 163.367
R372 B.n122 B.n77 163.367
R373 B.n123 B.n122 163.367
R374 B.n124 B.n123 163.367
R375 B.n124 B.n75 163.367
R376 B.n128 B.n75 163.367
R377 B.n129 B.n128 163.367
R378 B.n130 B.n129 163.367
R379 B.n130 B.n73 163.367
R380 B.n134 B.n73 163.367
R381 B.n135 B.n134 163.367
R382 B.n136 B.n135 163.367
R383 B.n136 B.n69 163.367
R384 B.n141 B.n69 163.367
R385 B.n142 B.n141 163.367
R386 B.n143 B.n142 163.367
R387 B.n143 B.n67 163.367
R388 B.n147 B.n67 163.367
R389 B.n148 B.n147 163.367
R390 B.n149 B.n148 163.367
R391 B.n149 B.n65 163.367
R392 B.n156 B.n65 163.367
R393 B.n157 B.n156 163.367
R394 B.n158 B.n157 163.367
R395 B.n158 B.n63 163.367
R396 B.n162 B.n63 163.367
R397 B.n163 B.n162 163.367
R398 B.n164 B.n163 163.367
R399 B.n164 B.n61 163.367
R400 B.n168 B.n61 163.367
R401 B.n169 B.n168 163.367
R402 B.n170 B.n169 163.367
R403 B.n170 B.n59 163.367
R404 B.n174 B.n59 163.367
R405 B.n175 B.n174 163.367
R406 B.n176 B.n175 163.367
R407 B.n176 B.n57 163.367
R408 B.n180 B.n57 163.367
R409 B.n181 B.n180 163.367
R410 B.n182 B.n181 163.367
R411 B.n236 B.n235 163.367
R412 B.n235 B.n234 163.367
R413 B.n234 B.n39 163.367
R414 B.n230 B.n39 163.367
R415 B.n230 B.n229 163.367
R416 B.n229 B.n228 163.367
R417 B.n228 B.n41 163.367
R418 B.n224 B.n41 163.367
R419 B.n224 B.n223 163.367
R420 B.n223 B.n222 163.367
R421 B.n222 B.n43 163.367
R422 B.n218 B.n43 163.367
R423 B.n218 B.n217 163.367
R424 B.n217 B.n216 163.367
R425 B.n216 B.n45 163.367
R426 B.n212 B.n45 163.367
R427 B.n212 B.n211 163.367
R428 B.n211 B.n210 163.367
R429 B.n210 B.n47 163.367
R430 B.n206 B.n47 163.367
R431 B.n206 B.n205 163.367
R432 B.n205 B.n204 163.367
R433 B.n204 B.n49 163.367
R434 B.n200 B.n49 163.367
R435 B.n200 B.n199 163.367
R436 B.n199 B.n198 163.367
R437 B.n198 B.n51 163.367
R438 B.n194 B.n51 163.367
R439 B.n194 B.n193 163.367
R440 B.n193 B.n192 163.367
R441 B.n192 B.n53 163.367
R442 B.n188 B.n53 163.367
R443 B.n188 B.n187 163.367
R444 B.n187 B.n186 163.367
R445 B.n186 B.n55 163.367
R446 B.n306 B.n11 163.367
R447 B.n302 B.n11 163.367
R448 B.n302 B.n301 163.367
R449 B.n301 B.n300 163.367
R450 B.n300 B.n13 163.367
R451 B.n296 B.n13 163.367
R452 B.n296 B.n295 163.367
R453 B.n295 B.n294 163.367
R454 B.n294 B.n15 163.367
R455 B.n290 B.n15 163.367
R456 B.n290 B.n289 163.367
R457 B.n289 B.n288 163.367
R458 B.n288 B.n17 163.367
R459 B.n284 B.n17 163.367
R460 B.n284 B.n283 163.367
R461 B.n283 B.n282 163.367
R462 B.n282 B.n19 163.367
R463 B.n277 B.n19 163.367
R464 B.n277 B.n276 163.367
R465 B.n276 B.n275 163.367
R466 B.n275 B.n23 163.367
R467 B.n271 B.n23 163.367
R468 B.n271 B.n270 163.367
R469 B.n270 B.n269 163.367
R470 B.n269 B.n25 163.367
R471 B.n265 B.n25 163.367
R472 B.n265 B.n264 163.367
R473 B.n264 B.n29 163.367
R474 B.n260 B.n29 163.367
R475 B.n260 B.n259 163.367
R476 B.n259 B.n258 163.367
R477 B.n258 B.n31 163.367
R478 B.n254 B.n31 163.367
R479 B.n254 B.n253 163.367
R480 B.n253 B.n252 163.367
R481 B.n252 B.n33 163.367
R482 B.n248 B.n33 163.367
R483 B.n248 B.n247 163.367
R484 B.n247 B.n246 163.367
R485 B.n246 B.n35 163.367
R486 B.n242 B.n35 163.367
R487 B.n242 B.n241 163.367
R488 B.n241 B.n240 163.367
R489 B.n240 B.n37 163.367
R490 B.n308 B.n307 163.367
R491 B.n308 B.n9 163.367
R492 B.n312 B.n9 163.367
R493 B.n313 B.n312 163.367
R494 B.n314 B.n313 163.367
R495 B.n314 B.n7 163.367
R496 B.n318 B.n7 163.367
R497 B.n319 B.n318 163.367
R498 B.n320 B.n319 163.367
R499 B.n320 B.n5 163.367
R500 B.n324 B.n5 163.367
R501 B.n325 B.n324 163.367
R502 B.n326 B.n325 163.367
R503 B.n326 B.n3 163.367
R504 B.n330 B.n3 163.367
R505 B.n331 B.n330 163.367
R506 B.n88 B.n2 163.367
R507 B.n88 B.n87 163.367
R508 B.n92 B.n87 163.367
R509 B.n93 B.n92 163.367
R510 B.n94 B.n93 163.367
R511 B.n94 B.n85 163.367
R512 B.n98 B.n85 163.367
R513 B.n99 B.n98 163.367
R514 B.n100 B.n99 163.367
R515 B.n100 B.n83 163.367
R516 B.n104 B.n83 163.367
R517 B.n105 B.n104 163.367
R518 B.n106 B.n105 163.367
R519 B.n106 B.n81 163.367
R520 B.n110 B.n81 163.367
R521 B.n111 B.n110 163.367
R522 B.n139 B.n71 59.5399
R523 B.n154 B.n153 59.5399
R524 B.n28 B.n27 59.5399
R525 B.n279 B.n21 59.5399
R526 B.n305 B.n10 32.9371
R527 B.n238 B.n237 32.9371
R528 B.n184 B.n183 32.9371
R529 B.n113 B.n80 32.9371
R530 B.n71 B.n70 30.8369
R531 B.n153 B.n152 30.8369
R532 B.n27 B.n26 30.8369
R533 B.n21 B.n20 30.8369
R534 B B.n333 18.0485
R535 B.n309 B.n10 10.6151
R536 B.n310 B.n309 10.6151
R537 B.n311 B.n310 10.6151
R538 B.n311 B.n8 10.6151
R539 B.n315 B.n8 10.6151
R540 B.n316 B.n315 10.6151
R541 B.n317 B.n316 10.6151
R542 B.n317 B.n6 10.6151
R543 B.n321 B.n6 10.6151
R544 B.n322 B.n321 10.6151
R545 B.n323 B.n322 10.6151
R546 B.n323 B.n4 10.6151
R547 B.n327 B.n4 10.6151
R548 B.n328 B.n327 10.6151
R549 B.n329 B.n328 10.6151
R550 B.n329 B.n0 10.6151
R551 B.n305 B.n304 10.6151
R552 B.n304 B.n303 10.6151
R553 B.n303 B.n12 10.6151
R554 B.n299 B.n12 10.6151
R555 B.n299 B.n298 10.6151
R556 B.n298 B.n297 10.6151
R557 B.n297 B.n14 10.6151
R558 B.n293 B.n14 10.6151
R559 B.n293 B.n292 10.6151
R560 B.n292 B.n291 10.6151
R561 B.n291 B.n16 10.6151
R562 B.n287 B.n16 10.6151
R563 B.n287 B.n286 10.6151
R564 B.n286 B.n285 10.6151
R565 B.n285 B.n18 10.6151
R566 B.n281 B.n18 10.6151
R567 B.n281 B.n280 10.6151
R568 B.n278 B.n22 10.6151
R569 B.n274 B.n22 10.6151
R570 B.n274 B.n273 10.6151
R571 B.n273 B.n272 10.6151
R572 B.n272 B.n24 10.6151
R573 B.n268 B.n24 10.6151
R574 B.n268 B.n267 10.6151
R575 B.n267 B.n266 10.6151
R576 B.n263 B.n262 10.6151
R577 B.n262 B.n261 10.6151
R578 B.n261 B.n30 10.6151
R579 B.n257 B.n30 10.6151
R580 B.n257 B.n256 10.6151
R581 B.n256 B.n255 10.6151
R582 B.n255 B.n32 10.6151
R583 B.n251 B.n32 10.6151
R584 B.n251 B.n250 10.6151
R585 B.n250 B.n249 10.6151
R586 B.n249 B.n34 10.6151
R587 B.n245 B.n34 10.6151
R588 B.n245 B.n244 10.6151
R589 B.n244 B.n243 10.6151
R590 B.n243 B.n36 10.6151
R591 B.n239 B.n36 10.6151
R592 B.n239 B.n238 10.6151
R593 B.n237 B.n38 10.6151
R594 B.n233 B.n38 10.6151
R595 B.n233 B.n232 10.6151
R596 B.n232 B.n231 10.6151
R597 B.n231 B.n40 10.6151
R598 B.n227 B.n40 10.6151
R599 B.n227 B.n226 10.6151
R600 B.n226 B.n225 10.6151
R601 B.n225 B.n42 10.6151
R602 B.n221 B.n42 10.6151
R603 B.n221 B.n220 10.6151
R604 B.n220 B.n219 10.6151
R605 B.n219 B.n44 10.6151
R606 B.n215 B.n44 10.6151
R607 B.n215 B.n214 10.6151
R608 B.n214 B.n213 10.6151
R609 B.n213 B.n46 10.6151
R610 B.n209 B.n46 10.6151
R611 B.n209 B.n208 10.6151
R612 B.n208 B.n207 10.6151
R613 B.n207 B.n48 10.6151
R614 B.n203 B.n48 10.6151
R615 B.n203 B.n202 10.6151
R616 B.n202 B.n201 10.6151
R617 B.n201 B.n50 10.6151
R618 B.n197 B.n50 10.6151
R619 B.n197 B.n196 10.6151
R620 B.n196 B.n195 10.6151
R621 B.n195 B.n52 10.6151
R622 B.n191 B.n52 10.6151
R623 B.n191 B.n190 10.6151
R624 B.n190 B.n189 10.6151
R625 B.n189 B.n54 10.6151
R626 B.n185 B.n54 10.6151
R627 B.n185 B.n184 10.6151
R628 B.n89 B.n1 10.6151
R629 B.n90 B.n89 10.6151
R630 B.n91 B.n90 10.6151
R631 B.n91 B.n86 10.6151
R632 B.n95 B.n86 10.6151
R633 B.n96 B.n95 10.6151
R634 B.n97 B.n96 10.6151
R635 B.n97 B.n84 10.6151
R636 B.n101 B.n84 10.6151
R637 B.n102 B.n101 10.6151
R638 B.n103 B.n102 10.6151
R639 B.n103 B.n82 10.6151
R640 B.n107 B.n82 10.6151
R641 B.n108 B.n107 10.6151
R642 B.n109 B.n108 10.6151
R643 B.n109 B.n80 10.6151
R644 B.n114 B.n113 10.6151
R645 B.n115 B.n114 10.6151
R646 B.n115 B.n78 10.6151
R647 B.n119 B.n78 10.6151
R648 B.n120 B.n119 10.6151
R649 B.n121 B.n120 10.6151
R650 B.n121 B.n76 10.6151
R651 B.n125 B.n76 10.6151
R652 B.n126 B.n125 10.6151
R653 B.n127 B.n126 10.6151
R654 B.n127 B.n74 10.6151
R655 B.n131 B.n74 10.6151
R656 B.n132 B.n131 10.6151
R657 B.n133 B.n132 10.6151
R658 B.n133 B.n72 10.6151
R659 B.n137 B.n72 10.6151
R660 B.n138 B.n137 10.6151
R661 B.n140 B.n68 10.6151
R662 B.n144 B.n68 10.6151
R663 B.n145 B.n144 10.6151
R664 B.n146 B.n145 10.6151
R665 B.n146 B.n66 10.6151
R666 B.n150 B.n66 10.6151
R667 B.n151 B.n150 10.6151
R668 B.n155 B.n151 10.6151
R669 B.n159 B.n64 10.6151
R670 B.n160 B.n159 10.6151
R671 B.n161 B.n160 10.6151
R672 B.n161 B.n62 10.6151
R673 B.n165 B.n62 10.6151
R674 B.n166 B.n165 10.6151
R675 B.n167 B.n166 10.6151
R676 B.n167 B.n60 10.6151
R677 B.n171 B.n60 10.6151
R678 B.n172 B.n171 10.6151
R679 B.n173 B.n172 10.6151
R680 B.n173 B.n58 10.6151
R681 B.n177 B.n58 10.6151
R682 B.n178 B.n177 10.6151
R683 B.n179 B.n178 10.6151
R684 B.n179 B.n56 10.6151
R685 B.n183 B.n56 10.6151
R686 B.n333 B.n0 8.11757
R687 B.n333 B.n1 8.11757
R688 B.n279 B.n278 6.5566
R689 B.n266 B.n28 6.5566
R690 B.n140 B.n139 6.5566
R691 B.n155 B.n154 6.5566
R692 B.n280 B.n279 4.05904
R693 B.n263 B.n28 4.05904
R694 B.n139 B.n138 4.05904
R695 B.n154 B.n64 4.05904
R696 VN VN.t0 221.629
R697 VN VN.t1 186.523
R698 VDD2.n33 VDD2.n19 756.745
R699 VDD2.n14 VDD2.n0 756.745
R700 VDD2.n34 VDD2.n33 585
R701 VDD2.n32 VDD2.n31 585
R702 VDD2.n23 VDD2.n22 585
R703 VDD2.n26 VDD2.n25 585
R704 VDD2.n7 VDD2.n6 585
R705 VDD2.n4 VDD2.n3 585
R706 VDD2.n13 VDD2.n12 585
R707 VDD2.n15 VDD2.n14 585
R708 VDD2.t1 VDD2.n24 330.707
R709 VDD2.t0 VDD2.n5 330.707
R710 VDD2.n33 VDD2.n32 171.744
R711 VDD2.n32 VDD2.n22 171.744
R712 VDD2.n25 VDD2.n22 171.744
R713 VDD2.n6 VDD2.n3 171.744
R714 VDD2.n13 VDD2.n3 171.744
R715 VDD2.n14 VDD2.n13 171.744
R716 VDD2.n25 VDD2.t1 85.8723
R717 VDD2.n6 VDD2.t0 85.8723
R718 VDD2.n38 VDD2.n18 79.7907
R719 VDD2.n38 VDD2.n37 50.0278
R720 VDD2.n26 VDD2.n24 16.3201
R721 VDD2.n7 VDD2.n5 16.3201
R722 VDD2.n27 VDD2.n23 12.8005
R723 VDD2.n8 VDD2.n4 12.8005
R724 VDD2.n31 VDD2.n30 12.0247
R725 VDD2.n12 VDD2.n11 12.0247
R726 VDD2.n34 VDD2.n21 11.249
R727 VDD2.n15 VDD2.n2 11.249
R728 VDD2.n35 VDD2.n19 10.4732
R729 VDD2.n16 VDD2.n0 10.4732
R730 VDD2.n37 VDD2.n36 9.45567
R731 VDD2.n18 VDD2.n17 9.45567
R732 VDD2.n36 VDD2.n35 9.3005
R733 VDD2.n21 VDD2.n20 9.3005
R734 VDD2.n30 VDD2.n29 9.3005
R735 VDD2.n28 VDD2.n27 9.3005
R736 VDD2.n17 VDD2.n16 9.3005
R737 VDD2.n2 VDD2.n1 9.3005
R738 VDD2.n11 VDD2.n10 9.3005
R739 VDD2.n9 VDD2.n8 9.3005
R740 VDD2.n28 VDD2.n24 3.78097
R741 VDD2.n9 VDD2.n5 3.78097
R742 VDD2.n37 VDD2.n19 3.49141
R743 VDD2.n18 VDD2.n0 3.49141
R744 VDD2.n35 VDD2.n34 2.71565
R745 VDD2.n16 VDD2.n15 2.71565
R746 VDD2.n31 VDD2.n21 1.93989
R747 VDD2.n12 VDD2.n2 1.93989
R748 VDD2.n30 VDD2.n23 1.16414
R749 VDD2.n11 VDD2.n4 1.16414
R750 VDD2 VDD2.n38 0.401362
R751 VDD2.n27 VDD2.n26 0.388379
R752 VDD2.n8 VDD2.n7 0.388379
R753 VDD2.n36 VDD2.n20 0.155672
R754 VDD2.n29 VDD2.n20 0.155672
R755 VDD2.n29 VDD2.n28 0.155672
R756 VDD2.n10 VDD2.n9 0.155672
R757 VDD2.n10 VDD2.n1 0.155672
R758 VDD2.n17 VDD2.n1 0.155672
C0 VN VP 3.33137f
C1 B VN 0.724506f
C2 VDD1 VN 0.152148f
C3 w_n1606_n1748# VN 1.93826f
C4 VTAIL VN 0.931975f
C5 B VP 1.05049f
C6 VDD1 VP 1.06906f
C7 VDD1 B 0.899559f
C8 w_n1606_n1748# VP 2.13892f
C9 VDD2 VN 0.941953f
C10 VTAIL VP 0.946197f
C11 B w_n1606_n1748# 5.09015f
C12 VDD1 w_n1606_n1748# 1.04658f
C13 VTAIL B 1.41598f
C14 VDD1 VTAIL 2.6307f
C15 VTAIL w_n1606_n1748# 1.54835f
C16 VDD2 VP 0.280974f
C17 B VDD2 0.918242f
C18 VDD1 VDD2 0.518067f
C19 w_n1606_n1748# VDD2 1.05643f
C20 VTAIL VDD2 2.67343f
C21 VDD2 VSUBS 0.496252f
C22 VDD1 VSUBS 1.848567f
C23 VTAIL VSUBS 0.381675f
C24 VN VSUBS 3.52636f
C25 VP VSUBS 0.888548f
C26 B VSUBS 2.117114f
C27 w_n1606_n1748# VSUBS 35.3641f
C28 VDD2.n0 VSUBS 0.016846f
C29 VDD2.n1 VSUBS 0.015756f
C30 VDD2.n2 VSUBS 0.008467f
C31 VDD2.n3 VSUBS 0.020012f
C32 VDD2.n4 VSUBS 0.008965f
C33 VDD2.n5 VSUBS 0.06067f
C34 VDD2.t0 VSUBS 0.044072f
C35 VDD2.n6 VSUBS 0.015009f
C36 VDD2.n7 VSUBS 0.012588f
C37 VDD2.n8 VSUBS 0.008467f
C38 VDD2.n9 VSUBS 0.209389f
C39 VDD2.n10 VSUBS 0.015756f
C40 VDD2.n11 VSUBS 0.008467f
C41 VDD2.n12 VSUBS 0.008965f
C42 VDD2.n13 VSUBS 0.020012f
C43 VDD2.n14 VSUBS 0.046859f
C44 VDD2.n15 VSUBS 0.008965f
C45 VDD2.n16 VSUBS 0.008467f
C46 VDD2.n17 VSUBS 0.037712f
C47 VDD2.n18 VSUBS 0.247789f
C48 VDD2.n19 VSUBS 0.016846f
C49 VDD2.n20 VSUBS 0.015756f
C50 VDD2.n21 VSUBS 0.008467f
C51 VDD2.n22 VSUBS 0.020012f
C52 VDD2.n23 VSUBS 0.008965f
C53 VDD2.n24 VSUBS 0.06067f
C54 VDD2.t1 VSUBS 0.044072f
C55 VDD2.n25 VSUBS 0.015009f
C56 VDD2.n26 VSUBS 0.012588f
C57 VDD2.n27 VSUBS 0.008467f
C58 VDD2.n28 VSUBS 0.209389f
C59 VDD2.n29 VSUBS 0.015756f
C60 VDD2.n30 VSUBS 0.008467f
C61 VDD2.n31 VSUBS 0.008965f
C62 VDD2.n32 VSUBS 0.020012f
C63 VDD2.n33 VSUBS 0.046859f
C64 VDD2.n34 VSUBS 0.008965f
C65 VDD2.n35 VSUBS 0.008467f
C66 VDD2.n36 VSUBS 0.037712f
C67 VDD2.n37 VSUBS 0.034403f
C68 VDD2.n38 VSUBS 1.21133f
C69 VN.t1 VSUBS 0.543937f
C70 VN.t0 VSUBS 0.716638f
C71 B.n0 VSUBS 0.006535f
C72 B.n1 VSUBS 0.006535f
C73 B.n2 VSUBS 0.009665f
C74 B.n3 VSUBS 0.007406f
C75 B.n4 VSUBS 0.007406f
C76 B.n5 VSUBS 0.007406f
C77 B.n6 VSUBS 0.007406f
C78 B.n7 VSUBS 0.007406f
C79 B.n8 VSUBS 0.007406f
C80 B.n9 VSUBS 0.007406f
C81 B.n10 VSUBS 0.017098f
C82 B.n11 VSUBS 0.007406f
C83 B.n12 VSUBS 0.007406f
C84 B.n13 VSUBS 0.007406f
C85 B.n14 VSUBS 0.007406f
C86 B.n15 VSUBS 0.007406f
C87 B.n16 VSUBS 0.007406f
C88 B.n17 VSUBS 0.007406f
C89 B.n18 VSUBS 0.007406f
C90 B.n19 VSUBS 0.007406f
C91 B.t7 VSUBS 0.059619f
C92 B.t8 VSUBS 0.07172f
C93 B.t6 VSUBS 0.24213f
C94 B.n20 VSUBS 0.130386f
C95 B.n21 VSUBS 0.114378f
C96 B.n22 VSUBS 0.007406f
C97 B.n23 VSUBS 0.007406f
C98 B.n24 VSUBS 0.007406f
C99 B.n25 VSUBS 0.007406f
C100 B.t10 VSUBS 0.05962f
C101 B.t11 VSUBS 0.071721f
C102 B.t9 VSUBS 0.24213f
C103 B.n26 VSUBS 0.130386f
C104 B.n27 VSUBS 0.114377f
C105 B.n28 VSUBS 0.017159f
C106 B.n29 VSUBS 0.007406f
C107 B.n30 VSUBS 0.007406f
C108 B.n31 VSUBS 0.007406f
C109 B.n32 VSUBS 0.007406f
C110 B.n33 VSUBS 0.007406f
C111 B.n34 VSUBS 0.007406f
C112 B.n35 VSUBS 0.007406f
C113 B.n36 VSUBS 0.007406f
C114 B.n37 VSUBS 0.017755f
C115 B.n38 VSUBS 0.007406f
C116 B.n39 VSUBS 0.007406f
C117 B.n40 VSUBS 0.007406f
C118 B.n41 VSUBS 0.007406f
C119 B.n42 VSUBS 0.007406f
C120 B.n43 VSUBS 0.007406f
C121 B.n44 VSUBS 0.007406f
C122 B.n45 VSUBS 0.007406f
C123 B.n46 VSUBS 0.007406f
C124 B.n47 VSUBS 0.007406f
C125 B.n48 VSUBS 0.007406f
C126 B.n49 VSUBS 0.007406f
C127 B.n50 VSUBS 0.007406f
C128 B.n51 VSUBS 0.007406f
C129 B.n52 VSUBS 0.007406f
C130 B.n53 VSUBS 0.007406f
C131 B.n54 VSUBS 0.007406f
C132 B.n55 VSUBS 0.017098f
C133 B.n56 VSUBS 0.007406f
C134 B.n57 VSUBS 0.007406f
C135 B.n58 VSUBS 0.007406f
C136 B.n59 VSUBS 0.007406f
C137 B.n60 VSUBS 0.007406f
C138 B.n61 VSUBS 0.007406f
C139 B.n62 VSUBS 0.007406f
C140 B.n63 VSUBS 0.007406f
C141 B.n64 VSUBS 0.005119f
C142 B.n65 VSUBS 0.007406f
C143 B.n66 VSUBS 0.007406f
C144 B.n67 VSUBS 0.007406f
C145 B.n68 VSUBS 0.007406f
C146 B.n69 VSUBS 0.007406f
C147 B.t2 VSUBS 0.059619f
C148 B.t1 VSUBS 0.07172f
C149 B.t0 VSUBS 0.24213f
C150 B.n70 VSUBS 0.130386f
C151 B.n71 VSUBS 0.114378f
C152 B.n72 VSUBS 0.007406f
C153 B.n73 VSUBS 0.007406f
C154 B.n74 VSUBS 0.007406f
C155 B.n75 VSUBS 0.007406f
C156 B.n76 VSUBS 0.007406f
C157 B.n77 VSUBS 0.007406f
C158 B.n78 VSUBS 0.007406f
C159 B.n79 VSUBS 0.007406f
C160 B.n80 VSUBS 0.017098f
C161 B.n81 VSUBS 0.007406f
C162 B.n82 VSUBS 0.007406f
C163 B.n83 VSUBS 0.007406f
C164 B.n84 VSUBS 0.007406f
C165 B.n85 VSUBS 0.007406f
C166 B.n86 VSUBS 0.007406f
C167 B.n87 VSUBS 0.007406f
C168 B.n88 VSUBS 0.007406f
C169 B.n89 VSUBS 0.007406f
C170 B.n90 VSUBS 0.007406f
C171 B.n91 VSUBS 0.007406f
C172 B.n92 VSUBS 0.007406f
C173 B.n93 VSUBS 0.007406f
C174 B.n94 VSUBS 0.007406f
C175 B.n95 VSUBS 0.007406f
C176 B.n96 VSUBS 0.007406f
C177 B.n97 VSUBS 0.007406f
C178 B.n98 VSUBS 0.007406f
C179 B.n99 VSUBS 0.007406f
C180 B.n100 VSUBS 0.007406f
C181 B.n101 VSUBS 0.007406f
C182 B.n102 VSUBS 0.007406f
C183 B.n103 VSUBS 0.007406f
C184 B.n104 VSUBS 0.007406f
C185 B.n105 VSUBS 0.007406f
C186 B.n106 VSUBS 0.007406f
C187 B.n107 VSUBS 0.007406f
C188 B.n108 VSUBS 0.007406f
C189 B.n109 VSUBS 0.007406f
C190 B.n110 VSUBS 0.007406f
C191 B.n111 VSUBS 0.017098f
C192 B.n112 VSUBS 0.017755f
C193 B.n113 VSUBS 0.017755f
C194 B.n114 VSUBS 0.007406f
C195 B.n115 VSUBS 0.007406f
C196 B.n116 VSUBS 0.007406f
C197 B.n117 VSUBS 0.007406f
C198 B.n118 VSUBS 0.007406f
C199 B.n119 VSUBS 0.007406f
C200 B.n120 VSUBS 0.007406f
C201 B.n121 VSUBS 0.007406f
C202 B.n122 VSUBS 0.007406f
C203 B.n123 VSUBS 0.007406f
C204 B.n124 VSUBS 0.007406f
C205 B.n125 VSUBS 0.007406f
C206 B.n126 VSUBS 0.007406f
C207 B.n127 VSUBS 0.007406f
C208 B.n128 VSUBS 0.007406f
C209 B.n129 VSUBS 0.007406f
C210 B.n130 VSUBS 0.007406f
C211 B.n131 VSUBS 0.007406f
C212 B.n132 VSUBS 0.007406f
C213 B.n133 VSUBS 0.007406f
C214 B.n134 VSUBS 0.007406f
C215 B.n135 VSUBS 0.007406f
C216 B.n136 VSUBS 0.007406f
C217 B.n137 VSUBS 0.007406f
C218 B.n138 VSUBS 0.005119f
C219 B.n139 VSUBS 0.017159f
C220 B.n140 VSUBS 0.00599f
C221 B.n141 VSUBS 0.007406f
C222 B.n142 VSUBS 0.007406f
C223 B.n143 VSUBS 0.007406f
C224 B.n144 VSUBS 0.007406f
C225 B.n145 VSUBS 0.007406f
C226 B.n146 VSUBS 0.007406f
C227 B.n147 VSUBS 0.007406f
C228 B.n148 VSUBS 0.007406f
C229 B.n149 VSUBS 0.007406f
C230 B.n150 VSUBS 0.007406f
C231 B.n151 VSUBS 0.007406f
C232 B.t5 VSUBS 0.05962f
C233 B.t4 VSUBS 0.071721f
C234 B.t3 VSUBS 0.24213f
C235 B.n152 VSUBS 0.130386f
C236 B.n153 VSUBS 0.114377f
C237 B.n154 VSUBS 0.017159f
C238 B.n155 VSUBS 0.00599f
C239 B.n156 VSUBS 0.007406f
C240 B.n157 VSUBS 0.007406f
C241 B.n158 VSUBS 0.007406f
C242 B.n159 VSUBS 0.007406f
C243 B.n160 VSUBS 0.007406f
C244 B.n161 VSUBS 0.007406f
C245 B.n162 VSUBS 0.007406f
C246 B.n163 VSUBS 0.007406f
C247 B.n164 VSUBS 0.007406f
C248 B.n165 VSUBS 0.007406f
C249 B.n166 VSUBS 0.007406f
C250 B.n167 VSUBS 0.007406f
C251 B.n168 VSUBS 0.007406f
C252 B.n169 VSUBS 0.007406f
C253 B.n170 VSUBS 0.007406f
C254 B.n171 VSUBS 0.007406f
C255 B.n172 VSUBS 0.007406f
C256 B.n173 VSUBS 0.007406f
C257 B.n174 VSUBS 0.007406f
C258 B.n175 VSUBS 0.007406f
C259 B.n176 VSUBS 0.007406f
C260 B.n177 VSUBS 0.007406f
C261 B.n178 VSUBS 0.007406f
C262 B.n179 VSUBS 0.007406f
C263 B.n180 VSUBS 0.007406f
C264 B.n181 VSUBS 0.007406f
C265 B.n182 VSUBS 0.017755f
C266 B.n183 VSUBS 0.016887f
C267 B.n184 VSUBS 0.017966f
C268 B.n185 VSUBS 0.007406f
C269 B.n186 VSUBS 0.007406f
C270 B.n187 VSUBS 0.007406f
C271 B.n188 VSUBS 0.007406f
C272 B.n189 VSUBS 0.007406f
C273 B.n190 VSUBS 0.007406f
C274 B.n191 VSUBS 0.007406f
C275 B.n192 VSUBS 0.007406f
C276 B.n193 VSUBS 0.007406f
C277 B.n194 VSUBS 0.007406f
C278 B.n195 VSUBS 0.007406f
C279 B.n196 VSUBS 0.007406f
C280 B.n197 VSUBS 0.007406f
C281 B.n198 VSUBS 0.007406f
C282 B.n199 VSUBS 0.007406f
C283 B.n200 VSUBS 0.007406f
C284 B.n201 VSUBS 0.007406f
C285 B.n202 VSUBS 0.007406f
C286 B.n203 VSUBS 0.007406f
C287 B.n204 VSUBS 0.007406f
C288 B.n205 VSUBS 0.007406f
C289 B.n206 VSUBS 0.007406f
C290 B.n207 VSUBS 0.007406f
C291 B.n208 VSUBS 0.007406f
C292 B.n209 VSUBS 0.007406f
C293 B.n210 VSUBS 0.007406f
C294 B.n211 VSUBS 0.007406f
C295 B.n212 VSUBS 0.007406f
C296 B.n213 VSUBS 0.007406f
C297 B.n214 VSUBS 0.007406f
C298 B.n215 VSUBS 0.007406f
C299 B.n216 VSUBS 0.007406f
C300 B.n217 VSUBS 0.007406f
C301 B.n218 VSUBS 0.007406f
C302 B.n219 VSUBS 0.007406f
C303 B.n220 VSUBS 0.007406f
C304 B.n221 VSUBS 0.007406f
C305 B.n222 VSUBS 0.007406f
C306 B.n223 VSUBS 0.007406f
C307 B.n224 VSUBS 0.007406f
C308 B.n225 VSUBS 0.007406f
C309 B.n226 VSUBS 0.007406f
C310 B.n227 VSUBS 0.007406f
C311 B.n228 VSUBS 0.007406f
C312 B.n229 VSUBS 0.007406f
C313 B.n230 VSUBS 0.007406f
C314 B.n231 VSUBS 0.007406f
C315 B.n232 VSUBS 0.007406f
C316 B.n233 VSUBS 0.007406f
C317 B.n234 VSUBS 0.007406f
C318 B.n235 VSUBS 0.007406f
C319 B.n236 VSUBS 0.017098f
C320 B.n237 VSUBS 0.017098f
C321 B.n238 VSUBS 0.017755f
C322 B.n239 VSUBS 0.007406f
C323 B.n240 VSUBS 0.007406f
C324 B.n241 VSUBS 0.007406f
C325 B.n242 VSUBS 0.007406f
C326 B.n243 VSUBS 0.007406f
C327 B.n244 VSUBS 0.007406f
C328 B.n245 VSUBS 0.007406f
C329 B.n246 VSUBS 0.007406f
C330 B.n247 VSUBS 0.007406f
C331 B.n248 VSUBS 0.007406f
C332 B.n249 VSUBS 0.007406f
C333 B.n250 VSUBS 0.007406f
C334 B.n251 VSUBS 0.007406f
C335 B.n252 VSUBS 0.007406f
C336 B.n253 VSUBS 0.007406f
C337 B.n254 VSUBS 0.007406f
C338 B.n255 VSUBS 0.007406f
C339 B.n256 VSUBS 0.007406f
C340 B.n257 VSUBS 0.007406f
C341 B.n258 VSUBS 0.007406f
C342 B.n259 VSUBS 0.007406f
C343 B.n260 VSUBS 0.007406f
C344 B.n261 VSUBS 0.007406f
C345 B.n262 VSUBS 0.007406f
C346 B.n263 VSUBS 0.005119f
C347 B.n264 VSUBS 0.007406f
C348 B.n265 VSUBS 0.007406f
C349 B.n266 VSUBS 0.00599f
C350 B.n267 VSUBS 0.007406f
C351 B.n268 VSUBS 0.007406f
C352 B.n269 VSUBS 0.007406f
C353 B.n270 VSUBS 0.007406f
C354 B.n271 VSUBS 0.007406f
C355 B.n272 VSUBS 0.007406f
C356 B.n273 VSUBS 0.007406f
C357 B.n274 VSUBS 0.007406f
C358 B.n275 VSUBS 0.007406f
C359 B.n276 VSUBS 0.007406f
C360 B.n277 VSUBS 0.007406f
C361 B.n278 VSUBS 0.00599f
C362 B.n279 VSUBS 0.017159f
C363 B.n280 VSUBS 0.005119f
C364 B.n281 VSUBS 0.007406f
C365 B.n282 VSUBS 0.007406f
C366 B.n283 VSUBS 0.007406f
C367 B.n284 VSUBS 0.007406f
C368 B.n285 VSUBS 0.007406f
C369 B.n286 VSUBS 0.007406f
C370 B.n287 VSUBS 0.007406f
C371 B.n288 VSUBS 0.007406f
C372 B.n289 VSUBS 0.007406f
C373 B.n290 VSUBS 0.007406f
C374 B.n291 VSUBS 0.007406f
C375 B.n292 VSUBS 0.007406f
C376 B.n293 VSUBS 0.007406f
C377 B.n294 VSUBS 0.007406f
C378 B.n295 VSUBS 0.007406f
C379 B.n296 VSUBS 0.007406f
C380 B.n297 VSUBS 0.007406f
C381 B.n298 VSUBS 0.007406f
C382 B.n299 VSUBS 0.007406f
C383 B.n300 VSUBS 0.007406f
C384 B.n301 VSUBS 0.007406f
C385 B.n302 VSUBS 0.007406f
C386 B.n303 VSUBS 0.007406f
C387 B.n304 VSUBS 0.007406f
C388 B.n305 VSUBS 0.017755f
C389 B.n306 VSUBS 0.017755f
C390 B.n307 VSUBS 0.017098f
C391 B.n308 VSUBS 0.007406f
C392 B.n309 VSUBS 0.007406f
C393 B.n310 VSUBS 0.007406f
C394 B.n311 VSUBS 0.007406f
C395 B.n312 VSUBS 0.007406f
C396 B.n313 VSUBS 0.007406f
C397 B.n314 VSUBS 0.007406f
C398 B.n315 VSUBS 0.007406f
C399 B.n316 VSUBS 0.007406f
C400 B.n317 VSUBS 0.007406f
C401 B.n318 VSUBS 0.007406f
C402 B.n319 VSUBS 0.007406f
C403 B.n320 VSUBS 0.007406f
C404 B.n321 VSUBS 0.007406f
C405 B.n322 VSUBS 0.007406f
C406 B.n323 VSUBS 0.007406f
C407 B.n324 VSUBS 0.007406f
C408 B.n325 VSUBS 0.007406f
C409 B.n326 VSUBS 0.007406f
C410 B.n327 VSUBS 0.007406f
C411 B.n328 VSUBS 0.007406f
C412 B.n329 VSUBS 0.007406f
C413 B.n330 VSUBS 0.007406f
C414 B.n331 VSUBS 0.009665f
C415 B.n332 VSUBS 0.010296f
C416 B.n333 VSUBS 0.020473f
C417 VDD1.n0 VSUBS 0.01588f
C418 VDD1.n1 VSUBS 0.014853f
C419 VDD1.n2 VSUBS 0.007981f
C420 VDD1.n3 VSUBS 0.018865f
C421 VDD1.n4 VSUBS 0.008451f
C422 VDD1.n5 VSUBS 0.057191f
C423 VDD1.t0 VSUBS 0.041545f
C424 VDD1.n6 VSUBS 0.014149f
C425 VDD1.n7 VSUBS 0.011866f
C426 VDD1.n8 VSUBS 0.007981f
C427 VDD1.n9 VSUBS 0.19738f
C428 VDD1.n10 VSUBS 0.014853f
C429 VDD1.n11 VSUBS 0.007981f
C430 VDD1.n12 VSUBS 0.008451f
C431 VDD1.n13 VSUBS 0.018865f
C432 VDD1.n14 VSUBS 0.044171f
C433 VDD1.n15 VSUBS 0.008451f
C434 VDD1.n16 VSUBS 0.007981f
C435 VDD1.n17 VSUBS 0.035549f
C436 VDD1.n18 VSUBS 0.032815f
C437 VDD1.n19 VSUBS 0.01588f
C438 VDD1.n20 VSUBS 0.014853f
C439 VDD1.n21 VSUBS 0.007981f
C440 VDD1.n22 VSUBS 0.018865f
C441 VDD1.n23 VSUBS 0.008451f
C442 VDD1.n24 VSUBS 0.057191f
C443 VDD1.t1 VSUBS 0.041545f
C444 VDD1.n25 VSUBS 0.014149f
C445 VDD1.n26 VSUBS 0.011866f
C446 VDD1.n27 VSUBS 0.007981f
C447 VDD1.n28 VSUBS 0.19738f
C448 VDD1.n29 VSUBS 0.014853f
C449 VDD1.n30 VSUBS 0.007981f
C450 VDD1.n31 VSUBS 0.008451f
C451 VDD1.n32 VSUBS 0.018865f
C452 VDD1.n33 VSUBS 0.044171f
C453 VDD1.n34 VSUBS 0.008451f
C454 VDD1.n35 VSUBS 0.007981f
C455 VDD1.n36 VSUBS 0.035549f
C456 VDD1.n37 VSUBS 0.252148f
C457 VTAIL.n0 VSUBS 0.019227f
C458 VTAIL.n1 VSUBS 0.017983f
C459 VTAIL.n2 VSUBS 0.009663f
C460 VTAIL.n3 VSUBS 0.022841f
C461 VTAIL.n4 VSUBS 0.010232f
C462 VTAIL.n5 VSUBS 0.069245f
C463 VTAIL.t3 VSUBS 0.050301f
C464 VTAIL.n6 VSUBS 0.017131f
C465 VTAIL.n7 VSUBS 0.014366f
C466 VTAIL.n8 VSUBS 0.009663f
C467 VTAIL.n9 VSUBS 0.238982f
C468 VTAIL.n10 VSUBS 0.017983f
C469 VTAIL.n11 VSUBS 0.009663f
C470 VTAIL.n12 VSUBS 0.010232f
C471 VTAIL.n13 VSUBS 0.022841f
C472 VTAIL.n14 VSUBS 0.053481f
C473 VTAIL.n15 VSUBS 0.010232f
C474 VTAIL.n16 VSUBS 0.009663f
C475 VTAIL.n17 VSUBS 0.043042f
C476 VTAIL.n18 VSUBS 0.026859f
C477 VTAIL.n19 VSUBS 0.664597f
C478 VTAIL.n20 VSUBS 0.019227f
C479 VTAIL.n21 VSUBS 0.017983f
C480 VTAIL.n22 VSUBS 0.009663f
C481 VTAIL.n23 VSUBS 0.022841f
C482 VTAIL.n24 VSUBS 0.010232f
C483 VTAIL.n25 VSUBS 0.069245f
C484 VTAIL.t1 VSUBS 0.050301f
C485 VTAIL.n26 VSUBS 0.017131f
C486 VTAIL.n27 VSUBS 0.014366f
C487 VTAIL.n28 VSUBS 0.009663f
C488 VTAIL.n29 VSUBS 0.238982f
C489 VTAIL.n30 VSUBS 0.017983f
C490 VTAIL.n31 VSUBS 0.009663f
C491 VTAIL.n32 VSUBS 0.010232f
C492 VTAIL.n33 VSUBS 0.022841f
C493 VTAIL.n34 VSUBS 0.053481f
C494 VTAIL.n35 VSUBS 0.010232f
C495 VTAIL.n36 VSUBS 0.009663f
C496 VTAIL.n37 VSUBS 0.043042f
C497 VTAIL.n38 VSUBS 0.026859f
C498 VTAIL.n39 VSUBS 0.681082f
C499 VTAIL.n40 VSUBS 0.019227f
C500 VTAIL.n41 VSUBS 0.017983f
C501 VTAIL.n42 VSUBS 0.009663f
C502 VTAIL.n43 VSUBS 0.022841f
C503 VTAIL.n44 VSUBS 0.010232f
C504 VTAIL.n45 VSUBS 0.069245f
C505 VTAIL.t2 VSUBS 0.050301f
C506 VTAIL.n46 VSUBS 0.017131f
C507 VTAIL.n47 VSUBS 0.014366f
C508 VTAIL.n48 VSUBS 0.009663f
C509 VTAIL.n49 VSUBS 0.238982f
C510 VTAIL.n50 VSUBS 0.017983f
C511 VTAIL.n51 VSUBS 0.009663f
C512 VTAIL.n52 VSUBS 0.010232f
C513 VTAIL.n53 VSUBS 0.022841f
C514 VTAIL.n54 VSUBS 0.053481f
C515 VTAIL.n55 VSUBS 0.010232f
C516 VTAIL.n56 VSUBS 0.009663f
C517 VTAIL.n57 VSUBS 0.043042f
C518 VTAIL.n58 VSUBS 0.026859f
C519 VTAIL.n59 VSUBS 0.601656f
C520 VTAIL.n60 VSUBS 0.019227f
C521 VTAIL.n61 VSUBS 0.017983f
C522 VTAIL.n62 VSUBS 0.009663f
C523 VTAIL.n63 VSUBS 0.022841f
C524 VTAIL.n64 VSUBS 0.010232f
C525 VTAIL.n65 VSUBS 0.069245f
C526 VTAIL.t0 VSUBS 0.050301f
C527 VTAIL.n66 VSUBS 0.017131f
C528 VTAIL.n67 VSUBS 0.014366f
C529 VTAIL.n68 VSUBS 0.009663f
C530 VTAIL.n69 VSUBS 0.238982f
C531 VTAIL.n70 VSUBS 0.017983f
C532 VTAIL.n71 VSUBS 0.009663f
C533 VTAIL.n72 VSUBS 0.010232f
C534 VTAIL.n73 VSUBS 0.022841f
C535 VTAIL.n74 VSUBS 0.053481f
C536 VTAIL.n75 VSUBS 0.010232f
C537 VTAIL.n76 VSUBS 0.009663f
C538 VTAIL.n77 VSUBS 0.043042f
C539 VTAIL.n78 VSUBS 0.026859f
C540 VTAIL.n79 VSUBS 0.551203f
C541 VP.t1 VSUBS 1.18161f
C542 VP.t0 VSUBS 0.90167f
C543 VP.n0 VSUBS 3.27137f
.ends

