* NGSPICE file created from diff_pair_sample_0334.ext - technology: sky130A

.subckt diff_pair_sample_0334 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=5.5653 ps=29.32 w=14.27 l=3.99
X1 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X2 VTAIL.t8 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X3 VTAIL.t7 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=2.35455 ps=14.6 w=14.27 l=3.99
X4 VTAIL.t11 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=0 ps=0 w=14.27 l=3.99
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=0 ps=0 w=14.27 l=3.99
X7 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=0 ps=0 w=14.27 l=3.99
X9 VTAIL.t13 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=2.35455 ps=14.6 w=14.27 l=3.99
X10 VDD1.t3 VP.t4 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=5.5653 ps=29.32 w=14.27 l=3.99
X11 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=0 ps=0 w=14.27 l=3.99
X12 VDD2.t4 VN.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=5.5653 ps=29.32 w=14.27 l=3.99
X13 VDD2.t3 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X14 VDD1.t2 VP.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X15 VDD1.t1 VP.t6 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X16 VTAIL.t4 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=2.35455 ps=14.6 w=14.27 l=3.99
X17 VDD2.t1 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.35455 pd=14.6 as=5.5653 ps=29.32 w=14.27 l=3.99
X18 VTAIL.t12 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=2.35455 ps=14.6 w=14.27 l=3.99
X19 VTAIL.t0 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5653 pd=29.32 as=2.35455 ps=14.6 w=14.27 l=3.99
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n13 161.3
R17 VP.n92 VP.n0 161.3
R18 VP.n91 VP.n90 161.3
R19 VP.n89 VP.n1 161.3
R20 VP.n88 VP.n87 161.3
R21 VP.n86 VP.n2 161.3
R22 VP.n85 VP.n84 161.3
R23 VP.n83 VP.n3 161.3
R24 VP.n82 VP.n81 161.3
R25 VP.n79 VP.n4 161.3
R26 VP.n78 VP.n77 161.3
R27 VP.n76 VP.n5 161.3
R28 VP.n75 VP.n74 161.3
R29 VP.n73 VP.n6 161.3
R30 VP.n72 VP.n71 161.3
R31 VP.n70 VP.n7 161.3
R32 VP.n69 VP.n68 161.3
R33 VP.n67 VP.n8 161.3
R34 VP.n65 VP.n64 161.3
R35 VP.n63 VP.n9 161.3
R36 VP.n62 VP.n61 161.3
R37 VP.n60 VP.n10 161.3
R38 VP.n59 VP.n58 161.3
R39 VP.n57 VP.n11 161.3
R40 VP.n56 VP.n55 161.3
R41 VP.n54 VP.n12 161.3
R42 VP.n22 VP.t7 118.239
R43 VP.n53 VP.t3 86.1927
R44 VP.n66 VP.t5 86.1927
R45 VP.n80 VP.t2 86.1927
R46 VP.n93 VP.t4 86.1927
R47 VP.n50 VP.t0 86.1927
R48 VP.n37 VP.t1 86.1927
R49 VP.n23 VP.t6 86.1927
R50 VP.n23 VP.n22 67.3497
R51 VP.n52 VP.n51 59.4131
R52 VP.n53 VP.n52 58.6935
R53 VP.n94 VP.n93 58.6935
R54 VP.n51 VP.n50 58.6935
R55 VP.n60 VP.n59 56.5193
R56 VP.n44 VP.n43 56.5193
R57 VP.n87 VP.n86 56.5193
R58 VP.n73 VP.n72 40.4934
R59 VP.n74 VP.n73 40.4934
R60 VP.n31 VP.n30 40.4934
R61 VP.n30 VP.n29 40.4934
R62 VP.n55 VP.n54 24.4675
R63 VP.n55 VP.n11 24.4675
R64 VP.n59 VP.n11 24.4675
R65 VP.n61 VP.n60 24.4675
R66 VP.n61 VP.n9 24.4675
R67 VP.n65 VP.n9 24.4675
R68 VP.n68 VP.n67 24.4675
R69 VP.n68 VP.n7 24.4675
R70 VP.n72 VP.n7 24.4675
R71 VP.n74 VP.n5 24.4675
R72 VP.n78 VP.n5 24.4675
R73 VP.n79 VP.n78 24.4675
R74 VP.n81 VP.n3 24.4675
R75 VP.n85 VP.n3 24.4675
R76 VP.n86 VP.n85 24.4675
R77 VP.n87 VP.n1 24.4675
R78 VP.n91 VP.n1 24.4675
R79 VP.n92 VP.n91 24.4675
R80 VP.n44 VP.n14 24.4675
R81 VP.n48 VP.n14 24.4675
R82 VP.n49 VP.n48 24.4675
R83 VP.n31 VP.n18 24.4675
R84 VP.n35 VP.n18 24.4675
R85 VP.n36 VP.n35 24.4675
R86 VP.n38 VP.n16 24.4675
R87 VP.n42 VP.n16 24.4675
R88 VP.n43 VP.n42 24.4675
R89 VP.n25 VP.n24 24.4675
R90 VP.n25 VP.n20 24.4675
R91 VP.n29 VP.n20 24.4675
R92 VP.n54 VP.n53 23.4888
R93 VP.n93 VP.n92 23.4888
R94 VP.n50 VP.n49 23.4888
R95 VP.n66 VP.n65 16.6381
R96 VP.n81 VP.n80 16.6381
R97 VP.n38 VP.n37 16.6381
R98 VP.n67 VP.n66 7.82994
R99 VP.n80 VP.n79 7.82994
R100 VP.n37 VP.n36 7.82994
R101 VP.n24 VP.n23 7.82994
R102 VP.n22 VP.n21 2.57369
R103 VP.n51 VP.n13 0.417535
R104 VP.n52 VP.n12 0.417535
R105 VP.n94 VP.n0 0.417535
R106 VP VP.n94 0.394291
R107 VP.n26 VP.n21 0.189894
R108 VP.n27 VP.n26 0.189894
R109 VP.n28 VP.n27 0.189894
R110 VP.n28 VP.n19 0.189894
R111 VP.n32 VP.n19 0.189894
R112 VP.n33 VP.n32 0.189894
R113 VP.n34 VP.n33 0.189894
R114 VP.n34 VP.n17 0.189894
R115 VP.n39 VP.n17 0.189894
R116 VP.n40 VP.n39 0.189894
R117 VP.n41 VP.n40 0.189894
R118 VP.n41 VP.n15 0.189894
R119 VP.n45 VP.n15 0.189894
R120 VP.n46 VP.n45 0.189894
R121 VP.n47 VP.n46 0.189894
R122 VP.n47 VP.n13 0.189894
R123 VP.n56 VP.n12 0.189894
R124 VP.n57 VP.n56 0.189894
R125 VP.n58 VP.n57 0.189894
R126 VP.n58 VP.n10 0.189894
R127 VP.n62 VP.n10 0.189894
R128 VP.n63 VP.n62 0.189894
R129 VP.n64 VP.n63 0.189894
R130 VP.n64 VP.n8 0.189894
R131 VP.n69 VP.n8 0.189894
R132 VP.n70 VP.n69 0.189894
R133 VP.n71 VP.n70 0.189894
R134 VP.n71 VP.n6 0.189894
R135 VP.n75 VP.n6 0.189894
R136 VP.n76 VP.n75 0.189894
R137 VP.n77 VP.n76 0.189894
R138 VP.n77 VP.n4 0.189894
R139 VP.n82 VP.n4 0.189894
R140 VP.n83 VP.n82 0.189894
R141 VP.n84 VP.n83 0.189894
R142 VP.n84 VP.n2 0.189894
R143 VP.n88 VP.n2 0.189894
R144 VP.n89 VP.n88 0.189894
R145 VP.n90 VP.n89 0.189894
R146 VP.n90 VP.n0 0.189894
R147 VTAIL.n626 VTAIL.n554 289.615
R148 VTAIL.n74 VTAIL.n2 289.615
R149 VTAIL.n152 VTAIL.n80 289.615
R150 VTAIL.n232 VTAIL.n160 289.615
R151 VTAIL.n548 VTAIL.n476 289.615
R152 VTAIL.n468 VTAIL.n396 289.615
R153 VTAIL.n390 VTAIL.n318 289.615
R154 VTAIL.n310 VTAIL.n238 289.615
R155 VTAIL.n578 VTAIL.n577 185
R156 VTAIL.n583 VTAIL.n582 185
R157 VTAIL.n585 VTAIL.n584 185
R158 VTAIL.n574 VTAIL.n573 185
R159 VTAIL.n591 VTAIL.n590 185
R160 VTAIL.n593 VTAIL.n592 185
R161 VTAIL.n570 VTAIL.n569 185
R162 VTAIL.n600 VTAIL.n599 185
R163 VTAIL.n601 VTAIL.n568 185
R164 VTAIL.n603 VTAIL.n602 185
R165 VTAIL.n566 VTAIL.n565 185
R166 VTAIL.n609 VTAIL.n608 185
R167 VTAIL.n611 VTAIL.n610 185
R168 VTAIL.n562 VTAIL.n561 185
R169 VTAIL.n617 VTAIL.n616 185
R170 VTAIL.n619 VTAIL.n618 185
R171 VTAIL.n558 VTAIL.n557 185
R172 VTAIL.n625 VTAIL.n624 185
R173 VTAIL.n627 VTAIL.n626 185
R174 VTAIL.n26 VTAIL.n25 185
R175 VTAIL.n31 VTAIL.n30 185
R176 VTAIL.n33 VTAIL.n32 185
R177 VTAIL.n22 VTAIL.n21 185
R178 VTAIL.n39 VTAIL.n38 185
R179 VTAIL.n41 VTAIL.n40 185
R180 VTAIL.n18 VTAIL.n17 185
R181 VTAIL.n48 VTAIL.n47 185
R182 VTAIL.n49 VTAIL.n16 185
R183 VTAIL.n51 VTAIL.n50 185
R184 VTAIL.n14 VTAIL.n13 185
R185 VTAIL.n57 VTAIL.n56 185
R186 VTAIL.n59 VTAIL.n58 185
R187 VTAIL.n10 VTAIL.n9 185
R188 VTAIL.n65 VTAIL.n64 185
R189 VTAIL.n67 VTAIL.n66 185
R190 VTAIL.n6 VTAIL.n5 185
R191 VTAIL.n73 VTAIL.n72 185
R192 VTAIL.n75 VTAIL.n74 185
R193 VTAIL.n104 VTAIL.n103 185
R194 VTAIL.n109 VTAIL.n108 185
R195 VTAIL.n111 VTAIL.n110 185
R196 VTAIL.n100 VTAIL.n99 185
R197 VTAIL.n117 VTAIL.n116 185
R198 VTAIL.n119 VTAIL.n118 185
R199 VTAIL.n96 VTAIL.n95 185
R200 VTAIL.n126 VTAIL.n125 185
R201 VTAIL.n127 VTAIL.n94 185
R202 VTAIL.n129 VTAIL.n128 185
R203 VTAIL.n92 VTAIL.n91 185
R204 VTAIL.n135 VTAIL.n134 185
R205 VTAIL.n137 VTAIL.n136 185
R206 VTAIL.n88 VTAIL.n87 185
R207 VTAIL.n143 VTAIL.n142 185
R208 VTAIL.n145 VTAIL.n144 185
R209 VTAIL.n84 VTAIL.n83 185
R210 VTAIL.n151 VTAIL.n150 185
R211 VTAIL.n153 VTAIL.n152 185
R212 VTAIL.n184 VTAIL.n183 185
R213 VTAIL.n189 VTAIL.n188 185
R214 VTAIL.n191 VTAIL.n190 185
R215 VTAIL.n180 VTAIL.n179 185
R216 VTAIL.n197 VTAIL.n196 185
R217 VTAIL.n199 VTAIL.n198 185
R218 VTAIL.n176 VTAIL.n175 185
R219 VTAIL.n206 VTAIL.n205 185
R220 VTAIL.n207 VTAIL.n174 185
R221 VTAIL.n209 VTAIL.n208 185
R222 VTAIL.n172 VTAIL.n171 185
R223 VTAIL.n215 VTAIL.n214 185
R224 VTAIL.n217 VTAIL.n216 185
R225 VTAIL.n168 VTAIL.n167 185
R226 VTAIL.n223 VTAIL.n222 185
R227 VTAIL.n225 VTAIL.n224 185
R228 VTAIL.n164 VTAIL.n163 185
R229 VTAIL.n231 VTAIL.n230 185
R230 VTAIL.n233 VTAIL.n232 185
R231 VTAIL.n549 VTAIL.n548 185
R232 VTAIL.n547 VTAIL.n546 185
R233 VTAIL.n480 VTAIL.n479 185
R234 VTAIL.n541 VTAIL.n540 185
R235 VTAIL.n539 VTAIL.n538 185
R236 VTAIL.n484 VTAIL.n483 185
R237 VTAIL.n533 VTAIL.n532 185
R238 VTAIL.n531 VTAIL.n530 185
R239 VTAIL.n488 VTAIL.n487 185
R240 VTAIL.n525 VTAIL.n524 185
R241 VTAIL.n523 VTAIL.n490 185
R242 VTAIL.n522 VTAIL.n521 185
R243 VTAIL.n493 VTAIL.n491 185
R244 VTAIL.n516 VTAIL.n515 185
R245 VTAIL.n514 VTAIL.n513 185
R246 VTAIL.n497 VTAIL.n496 185
R247 VTAIL.n508 VTAIL.n507 185
R248 VTAIL.n506 VTAIL.n505 185
R249 VTAIL.n501 VTAIL.n500 185
R250 VTAIL.n469 VTAIL.n468 185
R251 VTAIL.n467 VTAIL.n466 185
R252 VTAIL.n400 VTAIL.n399 185
R253 VTAIL.n461 VTAIL.n460 185
R254 VTAIL.n459 VTAIL.n458 185
R255 VTAIL.n404 VTAIL.n403 185
R256 VTAIL.n453 VTAIL.n452 185
R257 VTAIL.n451 VTAIL.n450 185
R258 VTAIL.n408 VTAIL.n407 185
R259 VTAIL.n445 VTAIL.n444 185
R260 VTAIL.n443 VTAIL.n410 185
R261 VTAIL.n442 VTAIL.n441 185
R262 VTAIL.n413 VTAIL.n411 185
R263 VTAIL.n436 VTAIL.n435 185
R264 VTAIL.n434 VTAIL.n433 185
R265 VTAIL.n417 VTAIL.n416 185
R266 VTAIL.n428 VTAIL.n427 185
R267 VTAIL.n426 VTAIL.n425 185
R268 VTAIL.n421 VTAIL.n420 185
R269 VTAIL.n391 VTAIL.n390 185
R270 VTAIL.n389 VTAIL.n388 185
R271 VTAIL.n322 VTAIL.n321 185
R272 VTAIL.n383 VTAIL.n382 185
R273 VTAIL.n381 VTAIL.n380 185
R274 VTAIL.n326 VTAIL.n325 185
R275 VTAIL.n375 VTAIL.n374 185
R276 VTAIL.n373 VTAIL.n372 185
R277 VTAIL.n330 VTAIL.n329 185
R278 VTAIL.n367 VTAIL.n366 185
R279 VTAIL.n365 VTAIL.n332 185
R280 VTAIL.n364 VTAIL.n363 185
R281 VTAIL.n335 VTAIL.n333 185
R282 VTAIL.n358 VTAIL.n357 185
R283 VTAIL.n356 VTAIL.n355 185
R284 VTAIL.n339 VTAIL.n338 185
R285 VTAIL.n350 VTAIL.n349 185
R286 VTAIL.n348 VTAIL.n347 185
R287 VTAIL.n343 VTAIL.n342 185
R288 VTAIL.n311 VTAIL.n310 185
R289 VTAIL.n309 VTAIL.n308 185
R290 VTAIL.n242 VTAIL.n241 185
R291 VTAIL.n303 VTAIL.n302 185
R292 VTAIL.n301 VTAIL.n300 185
R293 VTAIL.n246 VTAIL.n245 185
R294 VTAIL.n295 VTAIL.n294 185
R295 VTAIL.n293 VTAIL.n292 185
R296 VTAIL.n250 VTAIL.n249 185
R297 VTAIL.n287 VTAIL.n286 185
R298 VTAIL.n285 VTAIL.n252 185
R299 VTAIL.n284 VTAIL.n283 185
R300 VTAIL.n255 VTAIL.n253 185
R301 VTAIL.n278 VTAIL.n277 185
R302 VTAIL.n276 VTAIL.n275 185
R303 VTAIL.n259 VTAIL.n258 185
R304 VTAIL.n270 VTAIL.n269 185
R305 VTAIL.n268 VTAIL.n267 185
R306 VTAIL.n263 VTAIL.n262 185
R307 VTAIL.n579 VTAIL.t2 149.524
R308 VTAIL.n27 VTAIL.t0 149.524
R309 VTAIL.n105 VTAIL.t15 149.524
R310 VTAIL.n185 VTAIL.t13 149.524
R311 VTAIL.n502 VTAIL.t9 149.524
R312 VTAIL.n422 VTAIL.t12 149.524
R313 VTAIL.n344 VTAIL.t5 149.524
R314 VTAIL.n264 VTAIL.t7 149.524
R315 VTAIL.n583 VTAIL.n577 104.615
R316 VTAIL.n584 VTAIL.n583 104.615
R317 VTAIL.n584 VTAIL.n573 104.615
R318 VTAIL.n591 VTAIL.n573 104.615
R319 VTAIL.n592 VTAIL.n591 104.615
R320 VTAIL.n592 VTAIL.n569 104.615
R321 VTAIL.n600 VTAIL.n569 104.615
R322 VTAIL.n601 VTAIL.n600 104.615
R323 VTAIL.n602 VTAIL.n601 104.615
R324 VTAIL.n602 VTAIL.n565 104.615
R325 VTAIL.n609 VTAIL.n565 104.615
R326 VTAIL.n610 VTAIL.n609 104.615
R327 VTAIL.n610 VTAIL.n561 104.615
R328 VTAIL.n617 VTAIL.n561 104.615
R329 VTAIL.n618 VTAIL.n617 104.615
R330 VTAIL.n618 VTAIL.n557 104.615
R331 VTAIL.n625 VTAIL.n557 104.615
R332 VTAIL.n626 VTAIL.n625 104.615
R333 VTAIL.n31 VTAIL.n25 104.615
R334 VTAIL.n32 VTAIL.n31 104.615
R335 VTAIL.n32 VTAIL.n21 104.615
R336 VTAIL.n39 VTAIL.n21 104.615
R337 VTAIL.n40 VTAIL.n39 104.615
R338 VTAIL.n40 VTAIL.n17 104.615
R339 VTAIL.n48 VTAIL.n17 104.615
R340 VTAIL.n49 VTAIL.n48 104.615
R341 VTAIL.n50 VTAIL.n49 104.615
R342 VTAIL.n50 VTAIL.n13 104.615
R343 VTAIL.n57 VTAIL.n13 104.615
R344 VTAIL.n58 VTAIL.n57 104.615
R345 VTAIL.n58 VTAIL.n9 104.615
R346 VTAIL.n65 VTAIL.n9 104.615
R347 VTAIL.n66 VTAIL.n65 104.615
R348 VTAIL.n66 VTAIL.n5 104.615
R349 VTAIL.n73 VTAIL.n5 104.615
R350 VTAIL.n74 VTAIL.n73 104.615
R351 VTAIL.n109 VTAIL.n103 104.615
R352 VTAIL.n110 VTAIL.n109 104.615
R353 VTAIL.n110 VTAIL.n99 104.615
R354 VTAIL.n117 VTAIL.n99 104.615
R355 VTAIL.n118 VTAIL.n117 104.615
R356 VTAIL.n118 VTAIL.n95 104.615
R357 VTAIL.n126 VTAIL.n95 104.615
R358 VTAIL.n127 VTAIL.n126 104.615
R359 VTAIL.n128 VTAIL.n127 104.615
R360 VTAIL.n128 VTAIL.n91 104.615
R361 VTAIL.n135 VTAIL.n91 104.615
R362 VTAIL.n136 VTAIL.n135 104.615
R363 VTAIL.n136 VTAIL.n87 104.615
R364 VTAIL.n143 VTAIL.n87 104.615
R365 VTAIL.n144 VTAIL.n143 104.615
R366 VTAIL.n144 VTAIL.n83 104.615
R367 VTAIL.n151 VTAIL.n83 104.615
R368 VTAIL.n152 VTAIL.n151 104.615
R369 VTAIL.n189 VTAIL.n183 104.615
R370 VTAIL.n190 VTAIL.n189 104.615
R371 VTAIL.n190 VTAIL.n179 104.615
R372 VTAIL.n197 VTAIL.n179 104.615
R373 VTAIL.n198 VTAIL.n197 104.615
R374 VTAIL.n198 VTAIL.n175 104.615
R375 VTAIL.n206 VTAIL.n175 104.615
R376 VTAIL.n207 VTAIL.n206 104.615
R377 VTAIL.n208 VTAIL.n207 104.615
R378 VTAIL.n208 VTAIL.n171 104.615
R379 VTAIL.n215 VTAIL.n171 104.615
R380 VTAIL.n216 VTAIL.n215 104.615
R381 VTAIL.n216 VTAIL.n167 104.615
R382 VTAIL.n223 VTAIL.n167 104.615
R383 VTAIL.n224 VTAIL.n223 104.615
R384 VTAIL.n224 VTAIL.n163 104.615
R385 VTAIL.n231 VTAIL.n163 104.615
R386 VTAIL.n232 VTAIL.n231 104.615
R387 VTAIL.n548 VTAIL.n547 104.615
R388 VTAIL.n547 VTAIL.n479 104.615
R389 VTAIL.n540 VTAIL.n479 104.615
R390 VTAIL.n540 VTAIL.n539 104.615
R391 VTAIL.n539 VTAIL.n483 104.615
R392 VTAIL.n532 VTAIL.n483 104.615
R393 VTAIL.n532 VTAIL.n531 104.615
R394 VTAIL.n531 VTAIL.n487 104.615
R395 VTAIL.n524 VTAIL.n487 104.615
R396 VTAIL.n524 VTAIL.n523 104.615
R397 VTAIL.n523 VTAIL.n522 104.615
R398 VTAIL.n522 VTAIL.n491 104.615
R399 VTAIL.n515 VTAIL.n491 104.615
R400 VTAIL.n515 VTAIL.n514 104.615
R401 VTAIL.n514 VTAIL.n496 104.615
R402 VTAIL.n507 VTAIL.n496 104.615
R403 VTAIL.n507 VTAIL.n506 104.615
R404 VTAIL.n506 VTAIL.n500 104.615
R405 VTAIL.n468 VTAIL.n467 104.615
R406 VTAIL.n467 VTAIL.n399 104.615
R407 VTAIL.n460 VTAIL.n399 104.615
R408 VTAIL.n460 VTAIL.n459 104.615
R409 VTAIL.n459 VTAIL.n403 104.615
R410 VTAIL.n452 VTAIL.n403 104.615
R411 VTAIL.n452 VTAIL.n451 104.615
R412 VTAIL.n451 VTAIL.n407 104.615
R413 VTAIL.n444 VTAIL.n407 104.615
R414 VTAIL.n444 VTAIL.n443 104.615
R415 VTAIL.n443 VTAIL.n442 104.615
R416 VTAIL.n442 VTAIL.n411 104.615
R417 VTAIL.n435 VTAIL.n411 104.615
R418 VTAIL.n435 VTAIL.n434 104.615
R419 VTAIL.n434 VTAIL.n416 104.615
R420 VTAIL.n427 VTAIL.n416 104.615
R421 VTAIL.n427 VTAIL.n426 104.615
R422 VTAIL.n426 VTAIL.n420 104.615
R423 VTAIL.n390 VTAIL.n389 104.615
R424 VTAIL.n389 VTAIL.n321 104.615
R425 VTAIL.n382 VTAIL.n321 104.615
R426 VTAIL.n382 VTAIL.n381 104.615
R427 VTAIL.n381 VTAIL.n325 104.615
R428 VTAIL.n374 VTAIL.n325 104.615
R429 VTAIL.n374 VTAIL.n373 104.615
R430 VTAIL.n373 VTAIL.n329 104.615
R431 VTAIL.n366 VTAIL.n329 104.615
R432 VTAIL.n366 VTAIL.n365 104.615
R433 VTAIL.n365 VTAIL.n364 104.615
R434 VTAIL.n364 VTAIL.n333 104.615
R435 VTAIL.n357 VTAIL.n333 104.615
R436 VTAIL.n357 VTAIL.n356 104.615
R437 VTAIL.n356 VTAIL.n338 104.615
R438 VTAIL.n349 VTAIL.n338 104.615
R439 VTAIL.n349 VTAIL.n348 104.615
R440 VTAIL.n348 VTAIL.n342 104.615
R441 VTAIL.n310 VTAIL.n309 104.615
R442 VTAIL.n309 VTAIL.n241 104.615
R443 VTAIL.n302 VTAIL.n241 104.615
R444 VTAIL.n302 VTAIL.n301 104.615
R445 VTAIL.n301 VTAIL.n245 104.615
R446 VTAIL.n294 VTAIL.n245 104.615
R447 VTAIL.n294 VTAIL.n293 104.615
R448 VTAIL.n293 VTAIL.n249 104.615
R449 VTAIL.n286 VTAIL.n249 104.615
R450 VTAIL.n286 VTAIL.n285 104.615
R451 VTAIL.n285 VTAIL.n284 104.615
R452 VTAIL.n284 VTAIL.n253 104.615
R453 VTAIL.n277 VTAIL.n253 104.615
R454 VTAIL.n277 VTAIL.n276 104.615
R455 VTAIL.n276 VTAIL.n258 104.615
R456 VTAIL.n269 VTAIL.n258 104.615
R457 VTAIL.n269 VTAIL.n268 104.615
R458 VTAIL.n268 VTAIL.n262 104.615
R459 VTAIL.t2 VTAIL.n577 52.3082
R460 VTAIL.t0 VTAIL.n25 52.3082
R461 VTAIL.t15 VTAIL.n103 52.3082
R462 VTAIL.t13 VTAIL.n183 52.3082
R463 VTAIL.t9 VTAIL.n500 52.3082
R464 VTAIL.t12 VTAIL.n420 52.3082
R465 VTAIL.t5 VTAIL.n342 52.3082
R466 VTAIL.t7 VTAIL.n262 52.3082
R467 VTAIL.n1 VTAIL.n0 44.5555
R468 VTAIL.n159 VTAIL.n158 44.5555
R469 VTAIL.n475 VTAIL.n474 44.5555
R470 VTAIL.n317 VTAIL.n316 44.5555
R471 VTAIL.n631 VTAIL.n630 31.9914
R472 VTAIL.n79 VTAIL.n78 31.9914
R473 VTAIL.n157 VTAIL.n156 31.9914
R474 VTAIL.n237 VTAIL.n236 31.9914
R475 VTAIL.n553 VTAIL.n552 31.9914
R476 VTAIL.n473 VTAIL.n472 31.9914
R477 VTAIL.n395 VTAIL.n394 31.9914
R478 VTAIL.n315 VTAIL.n314 31.9914
R479 VTAIL.n631 VTAIL.n553 28.3927
R480 VTAIL.n315 VTAIL.n237 28.3927
R481 VTAIL.n603 VTAIL.n568 13.1884
R482 VTAIL.n51 VTAIL.n16 13.1884
R483 VTAIL.n129 VTAIL.n94 13.1884
R484 VTAIL.n209 VTAIL.n174 13.1884
R485 VTAIL.n525 VTAIL.n490 13.1884
R486 VTAIL.n445 VTAIL.n410 13.1884
R487 VTAIL.n367 VTAIL.n332 13.1884
R488 VTAIL.n287 VTAIL.n252 13.1884
R489 VTAIL.n599 VTAIL.n598 12.8005
R490 VTAIL.n604 VTAIL.n566 12.8005
R491 VTAIL.n47 VTAIL.n46 12.8005
R492 VTAIL.n52 VTAIL.n14 12.8005
R493 VTAIL.n125 VTAIL.n124 12.8005
R494 VTAIL.n130 VTAIL.n92 12.8005
R495 VTAIL.n205 VTAIL.n204 12.8005
R496 VTAIL.n210 VTAIL.n172 12.8005
R497 VTAIL.n526 VTAIL.n488 12.8005
R498 VTAIL.n521 VTAIL.n492 12.8005
R499 VTAIL.n446 VTAIL.n408 12.8005
R500 VTAIL.n441 VTAIL.n412 12.8005
R501 VTAIL.n368 VTAIL.n330 12.8005
R502 VTAIL.n363 VTAIL.n334 12.8005
R503 VTAIL.n288 VTAIL.n250 12.8005
R504 VTAIL.n283 VTAIL.n254 12.8005
R505 VTAIL.n597 VTAIL.n570 12.0247
R506 VTAIL.n608 VTAIL.n607 12.0247
R507 VTAIL.n45 VTAIL.n18 12.0247
R508 VTAIL.n56 VTAIL.n55 12.0247
R509 VTAIL.n123 VTAIL.n96 12.0247
R510 VTAIL.n134 VTAIL.n133 12.0247
R511 VTAIL.n203 VTAIL.n176 12.0247
R512 VTAIL.n214 VTAIL.n213 12.0247
R513 VTAIL.n530 VTAIL.n529 12.0247
R514 VTAIL.n520 VTAIL.n493 12.0247
R515 VTAIL.n450 VTAIL.n449 12.0247
R516 VTAIL.n440 VTAIL.n413 12.0247
R517 VTAIL.n372 VTAIL.n371 12.0247
R518 VTAIL.n362 VTAIL.n335 12.0247
R519 VTAIL.n292 VTAIL.n291 12.0247
R520 VTAIL.n282 VTAIL.n255 12.0247
R521 VTAIL.n594 VTAIL.n593 11.249
R522 VTAIL.n611 VTAIL.n564 11.249
R523 VTAIL.n42 VTAIL.n41 11.249
R524 VTAIL.n59 VTAIL.n12 11.249
R525 VTAIL.n120 VTAIL.n119 11.249
R526 VTAIL.n137 VTAIL.n90 11.249
R527 VTAIL.n200 VTAIL.n199 11.249
R528 VTAIL.n217 VTAIL.n170 11.249
R529 VTAIL.n533 VTAIL.n486 11.249
R530 VTAIL.n517 VTAIL.n516 11.249
R531 VTAIL.n453 VTAIL.n406 11.249
R532 VTAIL.n437 VTAIL.n436 11.249
R533 VTAIL.n375 VTAIL.n328 11.249
R534 VTAIL.n359 VTAIL.n358 11.249
R535 VTAIL.n295 VTAIL.n248 11.249
R536 VTAIL.n279 VTAIL.n278 11.249
R537 VTAIL.n590 VTAIL.n572 10.4732
R538 VTAIL.n612 VTAIL.n562 10.4732
R539 VTAIL.n38 VTAIL.n20 10.4732
R540 VTAIL.n60 VTAIL.n10 10.4732
R541 VTAIL.n116 VTAIL.n98 10.4732
R542 VTAIL.n138 VTAIL.n88 10.4732
R543 VTAIL.n196 VTAIL.n178 10.4732
R544 VTAIL.n218 VTAIL.n168 10.4732
R545 VTAIL.n534 VTAIL.n484 10.4732
R546 VTAIL.n513 VTAIL.n495 10.4732
R547 VTAIL.n454 VTAIL.n404 10.4732
R548 VTAIL.n433 VTAIL.n415 10.4732
R549 VTAIL.n376 VTAIL.n326 10.4732
R550 VTAIL.n355 VTAIL.n337 10.4732
R551 VTAIL.n296 VTAIL.n246 10.4732
R552 VTAIL.n275 VTAIL.n257 10.4732
R553 VTAIL.n579 VTAIL.n578 10.2747
R554 VTAIL.n27 VTAIL.n26 10.2747
R555 VTAIL.n105 VTAIL.n104 10.2747
R556 VTAIL.n185 VTAIL.n184 10.2747
R557 VTAIL.n502 VTAIL.n501 10.2747
R558 VTAIL.n422 VTAIL.n421 10.2747
R559 VTAIL.n344 VTAIL.n343 10.2747
R560 VTAIL.n264 VTAIL.n263 10.2747
R561 VTAIL.n589 VTAIL.n574 9.69747
R562 VTAIL.n616 VTAIL.n615 9.69747
R563 VTAIL.n37 VTAIL.n22 9.69747
R564 VTAIL.n64 VTAIL.n63 9.69747
R565 VTAIL.n115 VTAIL.n100 9.69747
R566 VTAIL.n142 VTAIL.n141 9.69747
R567 VTAIL.n195 VTAIL.n180 9.69747
R568 VTAIL.n222 VTAIL.n221 9.69747
R569 VTAIL.n538 VTAIL.n537 9.69747
R570 VTAIL.n512 VTAIL.n497 9.69747
R571 VTAIL.n458 VTAIL.n457 9.69747
R572 VTAIL.n432 VTAIL.n417 9.69747
R573 VTAIL.n380 VTAIL.n379 9.69747
R574 VTAIL.n354 VTAIL.n339 9.69747
R575 VTAIL.n300 VTAIL.n299 9.69747
R576 VTAIL.n274 VTAIL.n259 9.69747
R577 VTAIL.n630 VTAIL.n629 9.45567
R578 VTAIL.n78 VTAIL.n77 9.45567
R579 VTAIL.n156 VTAIL.n155 9.45567
R580 VTAIL.n236 VTAIL.n235 9.45567
R581 VTAIL.n552 VTAIL.n551 9.45567
R582 VTAIL.n472 VTAIL.n471 9.45567
R583 VTAIL.n394 VTAIL.n393 9.45567
R584 VTAIL.n314 VTAIL.n313 9.45567
R585 VTAIL.n556 VTAIL.n555 9.3005
R586 VTAIL.n629 VTAIL.n628 9.3005
R587 VTAIL.n621 VTAIL.n620 9.3005
R588 VTAIL.n560 VTAIL.n559 9.3005
R589 VTAIL.n615 VTAIL.n614 9.3005
R590 VTAIL.n613 VTAIL.n612 9.3005
R591 VTAIL.n564 VTAIL.n563 9.3005
R592 VTAIL.n607 VTAIL.n606 9.3005
R593 VTAIL.n605 VTAIL.n604 9.3005
R594 VTAIL.n581 VTAIL.n580 9.3005
R595 VTAIL.n576 VTAIL.n575 9.3005
R596 VTAIL.n587 VTAIL.n586 9.3005
R597 VTAIL.n589 VTAIL.n588 9.3005
R598 VTAIL.n572 VTAIL.n571 9.3005
R599 VTAIL.n595 VTAIL.n594 9.3005
R600 VTAIL.n597 VTAIL.n596 9.3005
R601 VTAIL.n598 VTAIL.n567 9.3005
R602 VTAIL.n623 VTAIL.n622 9.3005
R603 VTAIL.n4 VTAIL.n3 9.3005
R604 VTAIL.n77 VTAIL.n76 9.3005
R605 VTAIL.n69 VTAIL.n68 9.3005
R606 VTAIL.n8 VTAIL.n7 9.3005
R607 VTAIL.n63 VTAIL.n62 9.3005
R608 VTAIL.n61 VTAIL.n60 9.3005
R609 VTAIL.n12 VTAIL.n11 9.3005
R610 VTAIL.n55 VTAIL.n54 9.3005
R611 VTAIL.n53 VTAIL.n52 9.3005
R612 VTAIL.n29 VTAIL.n28 9.3005
R613 VTAIL.n24 VTAIL.n23 9.3005
R614 VTAIL.n35 VTAIL.n34 9.3005
R615 VTAIL.n37 VTAIL.n36 9.3005
R616 VTAIL.n20 VTAIL.n19 9.3005
R617 VTAIL.n43 VTAIL.n42 9.3005
R618 VTAIL.n45 VTAIL.n44 9.3005
R619 VTAIL.n46 VTAIL.n15 9.3005
R620 VTAIL.n71 VTAIL.n70 9.3005
R621 VTAIL.n82 VTAIL.n81 9.3005
R622 VTAIL.n155 VTAIL.n154 9.3005
R623 VTAIL.n147 VTAIL.n146 9.3005
R624 VTAIL.n86 VTAIL.n85 9.3005
R625 VTAIL.n141 VTAIL.n140 9.3005
R626 VTAIL.n139 VTAIL.n138 9.3005
R627 VTAIL.n90 VTAIL.n89 9.3005
R628 VTAIL.n133 VTAIL.n132 9.3005
R629 VTAIL.n131 VTAIL.n130 9.3005
R630 VTAIL.n107 VTAIL.n106 9.3005
R631 VTAIL.n102 VTAIL.n101 9.3005
R632 VTAIL.n113 VTAIL.n112 9.3005
R633 VTAIL.n115 VTAIL.n114 9.3005
R634 VTAIL.n98 VTAIL.n97 9.3005
R635 VTAIL.n121 VTAIL.n120 9.3005
R636 VTAIL.n123 VTAIL.n122 9.3005
R637 VTAIL.n124 VTAIL.n93 9.3005
R638 VTAIL.n149 VTAIL.n148 9.3005
R639 VTAIL.n162 VTAIL.n161 9.3005
R640 VTAIL.n235 VTAIL.n234 9.3005
R641 VTAIL.n227 VTAIL.n226 9.3005
R642 VTAIL.n166 VTAIL.n165 9.3005
R643 VTAIL.n221 VTAIL.n220 9.3005
R644 VTAIL.n219 VTAIL.n218 9.3005
R645 VTAIL.n170 VTAIL.n169 9.3005
R646 VTAIL.n213 VTAIL.n212 9.3005
R647 VTAIL.n211 VTAIL.n210 9.3005
R648 VTAIL.n187 VTAIL.n186 9.3005
R649 VTAIL.n182 VTAIL.n181 9.3005
R650 VTAIL.n193 VTAIL.n192 9.3005
R651 VTAIL.n195 VTAIL.n194 9.3005
R652 VTAIL.n178 VTAIL.n177 9.3005
R653 VTAIL.n201 VTAIL.n200 9.3005
R654 VTAIL.n203 VTAIL.n202 9.3005
R655 VTAIL.n204 VTAIL.n173 9.3005
R656 VTAIL.n229 VTAIL.n228 9.3005
R657 VTAIL.n478 VTAIL.n477 9.3005
R658 VTAIL.n545 VTAIL.n544 9.3005
R659 VTAIL.n543 VTAIL.n542 9.3005
R660 VTAIL.n482 VTAIL.n481 9.3005
R661 VTAIL.n537 VTAIL.n536 9.3005
R662 VTAIL.n535 VTAIL.n534 9.3005
R663 VTAIL.n486 VTAIL.n485 9.3005
R664 VTAIL.n529 VTAIL.n528 9.3005
R665 VTAIL.n527 VTAIL.n526 9.3005
R666 VTAIL.n492 VTAIL.n489 9.3005
R667 VTAIL.n520 VTAIL.n519 9.3005
R668 VTAIL.n518 VTAIL.n517 9.3005
R669 VTAIL.n495 VTAIL.n494 9.3005
R670 VTAIL.n512 VTAIL.n511 9.3005
R671 VTAIL.n510 VTAIL.n509 9.3005
R672 VTAIL.n499 VTAIL.n498 9.3005
R673 VTAIL.n504 VTAIL.n503 9.3005
R674 VTAIL.n551 VTAIL.n550 9.3005
R675 VTAIL.n424 VTAIL.n423 9.3005
R676 VTAIL.n419 VTAIL.n418 9.3005
R677 VTAIL.n430 VTAIL.n429 9.3005
R678 VTAIL.n432 VTAIL.n431 9.3005
R679 VTAIL.n415 VTAIL.n414 9.3005
R680 VTAIL.n438 VTAIL.n437 9.3005
R681 VTAIL.n440 VTAIL.n439 9.3005
R682 VTAIL.n412 VTAIL.n409 9.3005
R683 VTAIL.n471 VTAIL.n470 9.3005
R684 VTAIL.n398 VTAIL.n397 9.3005
R685 VTAIL.n465 VTAIL.n464 9.3005
R686 VTAIL.n463 VTAIL.n462 9.3005
R687 VTAIL.n402 VTAIL.n401 9.3005
R688 VTAIL.n457 VTAIL.n456 9.3005
R689 VTAIL.n455 VTAIL.n454 9.3005
R690 VTAIL.n406 VTAIL.n405 9.3005
R691 VTAIL.n449 VTAIL.n448 9.3005
R692 VTAIL.n447 VTAIL.n446 9.3005
R693 VTAIL.n346 VTAIL.n345 9.3005
R694 VTAIL.n341 VTAIL.n340 9.3005
R695 VTAIL.n352 VTAIL.n351 9.3005
R696 VTAIL.n354 VTAIL.n353 9.3005
R697 VTAIL.n337 VTAIL.n336 9.3005
R698 VTAIL.n360 VTAIL.n359 9.3005
R699 VTAIL.n362 VTAIL.n361 9.3005
R700 VTAIL.n334 VTAIL.n331 9.3005
R701 VTAIL.n393 VTAIL.n392 9.3005
R702 VTAIL.n320 VTAIL.n319 9.3005
R703 VTAIL.n387 VTAIL.n386 9.3005
R704 VTAIL.n385 VTAIL.n384 9.3005
R705 VTAIL.n324 VTAIL.n323 9.3005
R706 VTAIL.n379 VTAIL.n378 9.3005
R707 VTAIL.n377 VTAIL.n376 9.3005
R708 VTAIL.n328 VTAIL.n327 9.3005
R709 VTAIL.n371 VTAIL.n370 9.3005
R710 VTAIL.n369 VTAIL.n368 9.3005
R711 VTAIL.n266 VTAIL.n265 9.3005
R712 VTAIL.n261 VTAIL.n260 9.3005
R713 VTAIL.n272 VTAIL.n271 9.3005
R714 VTAIL.n274 VTAIL.n273 9.3005
R715 VTAIL.n257 VTAIL.n256 9.3005
R716 VTAIL.n280 VTAIL.n279 9.3005
R717 VTAIL.n282 VTAIL.n281 9.3005
R718 VTAIL.n254 VTAIL.n251 9.3005
R719 VTAIL.n313 VTAIL.n312 9.3005
R720 VTAIL.n240 VTAIL.n239 9.3005
R721 VTAIL.n307 VTAIL.n306 9.3005
R722 VTAIL.n305 VTAIL.n304 9.3005
R723 VTAIL.n244 VTAIL.n243 9.3005
R724 VTAIL.n299 VTAIL.n298 9.3005
R725 VTAIL.n297 VTAIL.n296 9.3005
R726 VTAIL.n248 VTAIL.n247 9.3005
R727 VTAIL.n291 VTAIL.n290 9.3005
R728 VTAIL.n289 VTAIL.n288 9.3005
R729 VTAIL.n586 VTAIL.n585 8.92171
R730 VTAIL.n619 VTAIL.n560 8.92171
R731 VTAIL.n34 VTAIL.n33 8.92171
R732 VTAIL.n67 VTAIL.n8 8.92171
R733 VTAIL.n112 VTAIL.n111 8.92171
R734 VTAIL.n145 VTAIL.n86 8.92171
R735 VTAIL.n192 VTAIL.n191 8.92171
R736 VTAIL.n225 VTAIL.n166 8.92171
R737 VTAIL.n541 VTAIL.n482 8.92171
R738 VTAIL.n509 VTAIL.n508 8.92171
R739 VTAIL.n461 VTAIL.n402 8.92171
R740 VTAIL.n429 VTAIL.n428 8.92171
R741 VTAIL.n383 VTAIL.n324 8.92171
R742 VTAIL.n351 VTAIL.n350 8.92171
R743 VTAIL.n303 VTAIL.n244 8.92171
R744 VTAIL.n271 VTAIL.n270 8.92171
R745 VTAIL.n582 VTAIL.n576 8.14595
R746 VTAIL.n620 VTAIL.n558 8.14595
R747 VTAIL.n630 VTAIL.n554 8.14595
R748 VTAIL.n30 VTAIL.n24 8.14595
R749 VTAIL.n68 VTAIL.n6 8.14595
R750 VTAIL.n78 VTAIL.n2 8.14595
R751 VTAIL.n108 VTAIL.n102 8.14595
R752 VTAIL.n146 VTAIL.n84 8.14595
R753 VTAIL.n156 VTAIL.n80 8.14595
R754 VTAIL.n188 VTAIL.n182 8.14595
R755 VTAIL.n226 VTAIL.n164 8.14595
R756 VTAIL.n236 VTAIL.n160 8.14595
R757 VTAIL.n552 VTAIL.n476 8.14595
R758 VTAIL.n542 VTAIL.n480 8.14595
R759 VTAIL.n505 VTAIL.n499 8.14595
R760 VTAIL.n472 VTAIL.n396 8.14595
R761 VTAIL.n462 VTAIL.n400 8.14595
R762 VTAIL.n425 VTAIL.n419 8.14595
R763 VTAIL.n394 VTAIL.n318 8.14595
R764 VTAIL.n384 VTAIL.n322 8.14595
R765 VTAIL.n347 VTAIL.n341 8.14595
R766 VTAIL.n314 VTAIL.n238 8.14595
R767 VTAIL.n304 VTAIL.n242 8.14595
R768 VTAIL.n267 VTAIL.n261 8.14595
R769 VTAIL.n581 VTAIL.n578 7.3702
R770 VTAIL.n624 VTAIL.n623 7.3702
R771 VTAIL.n628 VTAIL.n627 7.3702
R772 VTAIL.n29 VTAIL.n26 7.3702
R773 VTAIL.n72 VTAIL.n71 7.3702
R774 VTAIL.n76 VTAIL.n75 7.3702
R775 VTAIL.n107 VTAIL.n104 7.3702
R776 VTAIL.n150 VTAIL.n149 7.3702
R777 VTAIL.n154 VTAIL.n153 7.3702
R778 VTAIL.n187 VTAIL.n184 7.3702
R779 VTAIL.n230 VTAIL.n229 7.3702
R780 VTAIL.n234 VTAIL.n233 7.3702
R781 VTAIL.n550 VTAIL.n549 7.3702
R782 VTAIL.n546 VTAIL.n545 7.3702
R783 VTAIL.n504 VTAIL.n501 7.3702
R784 VTAIL.n470 VTAIL.n469 7.3702
R785 VTAIL.n466 VTAIL.n465 7.3702
R786 VTAIL.n424 VTAIL.n421 7.3702
R787 VTAIL.n392 VTAIL.n391 7.3702
R788 VTAIL.n388 VTAIL.n387 7.3702
R789 VTAIL.n346 VTAIL.n343 7.3702
R790 VTAIL.n312 VTAIL.n311 7.3702
R791 VTAIL.n308 VTAIL.n307 7.3702
R792 VTAIL.n266 VTAIL.n263 7.3702
R793 VTAIL.n624 VTAIL.n556 6.59444
R794 VTAIL.n627 VTAIL.n556 6.59444
R795 VTAIL.n72 VTAIL.n4 6.59444
R796 VTAIL.n75 VTAIL.n4 6.59444
R797 VTAIL.n150 VTAIL.n82 6.59444
R798 VTAIL.n153 VTAIL.n82 6.59444
R799 VTAIL.n230 VTAIL.n162 6.59444
R800 VTAIL.n233 VTAIL.n162 6.59444
R801 VTAIL.n549 VTAIL.n478 6.59444
R802 VTAIL.n546 VTAIL.n478 6.59444
R803 VTAIL.n469 VTAIL.n398 6.59444
R804 VTAIL.n466 VTAIL.n398 6.59444
R805 VTAIL.n391 VTAIL.n320 6.59444
R806 VTAIL.n388 VTAIL.n320 6.59444
R807 VTAIL.n311 VTAIL.n240 6.59444
R808 VTAIL.n308 VTAIL.n240 6.59444
R809 VTAIL.n582 VTAIL.n581 5.81868
R810 VTAIL.n623 VTAIL.n558 5.81868
R811 VTAIL.n628 VTAIL.n554 5.81868
R812 VTAIL.n30 VTAIL.n29 5.81868
R813 VTAIL.n71 VTAIL.n6 5.81868
R814 VTAIL.n76 VTAIL.n2 5.81868
R815 VTAIL.n108 VTAIL.n107 5.81868
R816 VTAIL.n149 VTAIL.n84 5.81868
R817 VTAIL.n154 VTAIL.n80 5.81868
R818 VTAIL.n188 VTAIL.n187 5.81868
R819 VTAIL.n229 VTAIL.n164 5.81868
R820 VTAIL.n234 VTAIL.n160 5.81868
R821 VTAIL.n550 VTAIL.n476 5.81868
R822 VTAIL.n545 VTAIL.n480 5.81868
R823 VTAIL.n505 VTAIL.n504 5.81868
R824 VTAIL.n470 VTAIL.n396 5.81868
R825 VTAIL.n465 VTAIL.n400 5.81868
R826 VTAIL.n425 VTAIL.n424 5.81868
R827 VTAIL.n392 VTAIL.n318 5.81868
R828 VTAIL.n387 VTAIL.n322 5.81868
R829 VTAIL.n347 VTAIL.n346 5.81868
R830 VTAIL.n312 VTAIL.n238 5.81868
R831 VTAIL.n307 VTAIL.n242 5.81868
R832 VTAIL.n267 VTAIL.n266 5.81868
R833 VTAIL.n585 VTAIL.n576 5.04292
R834 VTAIL.n620 VTAIL.n619 5.04292
R835 VTAIL.n33 VTAIL.n24 5.04292
R836 VTAIL.n68 VTAIL.n67 5.04292
R837 VTAIL.n111 VTAIL.n102 5.04292
R838 VTAIL.n146 VTAIL.n145 5.04292
R839 VTAIL.n191 VTAIL.n182 5.04292
R840 VTAIL.n226 VTAIL.n225 5.04292
R841 VTAIL.n542 VTAIL.n541 5.04292
R842 VTAIL.n508 VTAIL.n499 5.04292
R843 VTAIL.n462 VTAIL.n461 5.04292
R844 VTAIL.n428 VTAIL.n419 5.04292
R845 VTAIL.n384 VTAIL.n383 5.04292
R846 VTAIL.n350 VTAIL.n341 5.04292
R847 VTAIL.n304 VTAIL.n303 5.04292
R848 VTAIL.n270 VTAIL.n261 5.04292
R849 VTAIL.n586 VTAIL.n574 4.26717
R850 VTAIL.n616 VTAIL.n560 4.26717
R851 VTAIL.n34 VTAIL.n22 4.26717
R852 VTAIL.n64 VTAIL.n8 4.26717
R853 VTAIL.n112 VTAIL.n100 4.26717
R854 VTAIL.n142 VTAIL.n86 4.26717
R855 VTAIL.n192 VTAIL.n180 4.26717
R856 VTAIL.n222 VTAIL.n166 4.26717
R857 VTAIL.n538 VTAIL.n482 4.26717
R858 VTAIL.n509 VTAIL.n497 4.26717
R859 VTAIL.n458 VTAIL.n402 4.26717
R860 VTAIL.n429 VTAIL.n417 4.26717
R861 VTAIL.n380 VTAIL.n324 4.26717
R862 VTAIL.n351 VTAIL.n339 4.26717
R863 VTAIL.n300 VTAIL.n244 4.26717
R864 VTAIL.n271 VTAIL.n259 4.26717
R865 VTAIL.n317 VTAIL.n315 3.72464
R866 VTAIL.n395 VTAIL.n317 3.72464
R867 VTAIL.n475 VTAIL.n473 3.72464
R868 VTAIL.n553 VTAIL.n475 3.72464
R869 VTAIL.n237 VTAIL.n159 3.72464
R870 VTAIL.n159 VTAIL.n157 3.72464
R871 VTAIL.n79 VTAIL.n1 3.72464
R872 VTAIL VTAIL.n631 3.66645
R873 VTAIL.n590 VTAIL.n589 3.49141
R874 VTAIL.n615 VTAIL.n562 3.49141
R875 VTAIL.n38 VTAIL.n37 3.49141
R876 VTAIL.n63 VTAIL.n10 3.49141
R877 VTAIL.n116 VTAIL.n115 3.49141
R878 VTAIL.n141 VTAIL.n88 3.49141
R879 VTAIL.n196 VTAIL.n195 3.49141
R880 VTAIL.n221 VTAIL.n168 3.49141
R881 VTAIL.n537 VTAIL.n484 3.49141
R882 VTAIL.n513 VTAIL.n512 3.49141
R883 VTAIL.n457 VTAIL.n404 3.49141
R884 VTAIL.n433 VTAIL.n432 3.49141
R885 VTAIL.n379 VTAIL.n326 3.49141
R886 VTAIL.n355 VTAIL.n354 3.49141
R887 VTAIL.n299 VTAIL.n246 3.49141
R888 VTAIL.n275 VTAIL.n274 3.49141
R889 VTAIL.n580 VTAIL.n579 2.84303
R890 VTAIL.n28 VTAIL.n27 2.84303
R891 VTAIL.n106 VTAIL.n105 2.84303
R892 VTAIL.n186 VTAIL.n185 2.84303
R893 VTAIL.n423 VTAIL.n422 2.84303
R894 VTAIL.n345 VTAIL.n344 2.84303
R895 VTAIL.n265 VTAIL.n264 2.84303
R896 VTAIL.n503 VTAIL.n502 2.84303
R897 VTAIL.n593 VTAIL.n572 2.71565
R898 VTAIL.n612 VTAIL.n611 2.71565
R899 VTAIL.n41 VTAIL.n20 2.71565
R900 VTAIL.n60 VTAIL.n59 2.71565
R901 VTAIL.n119 VTAIL.n98 2.71565
R902 VTAIL.n138 VTAIL.n137 2.71565
R903 VTAIL.n199 VTAIL.n178 2.71565
R904 VTAIL.n218 VTAIL.n217 2.71565
R905 VTAIL.n534 VTAIL.n533 2.71565
R906 VTAIL.n516 VTAIL.n495 2.71565
R907 VTAIL.n454 VTAIL.n453 2.71565
R908 VTAIL.n436 VTAIL.n415 2.71565
R909 VTAIL.n376 VTAIL.n375 2.71565
R910 VTAIL.n358 VTAIL.n337 2.71565
R911 VTAIL.n296 VTAIL.n295 2.71565
R912 VTAIL.n278 VTAIL.n257 2.71565
R913 VTAIL.n594 VTAIL.n570 1.93989
R914 VTAIL.n608 VTAIL.n564 1.93989
R915 VTAIL.n42 VTAIL.n18 1.93989
R916 VTAIL.n56 VTAIL.n12 1.93989
R917 VTAIL.n120 VTAIL.n96 1.93989
R918 VTAIL.n134 VTAIL.n90 1.93989
R919 VTAIL.n200 VTAIL.n176 1.93989
R920 VTAIL.n214 VTAIL.n170 1.93989
R921 VTAIL.n530 VTAIL.n486 1.93989
R922 VTAIL.n517 VTAIL.n493 1.93989
R923 VTAIL.n450 VTAIL.n406 1.93989
R924 VTAIL.n437 VTAIL.n413 1.93989
R925 VTAIL.n372 VTAIL.n328 1.93989
R926 VTAIL.n359 VTAIL.n335 1.93989
R927 VTAIL.n292 VTAIL.n248 1.93989
R928 VTAIL.n279 VTAIL.n255 1.93989
R929 VTAIL.n0 VTAIL.t6 1.38803
R930 VTAIL.n0 VTAIL.t3 1.38803
R931 VTAIL.n158 VTAIL.t10 1.38803
R932 VTAIL.n158 VTAIL.t11 1.38803
R933 VTAIL.n474 VTAIL.t14 1.38803
R934 VTAIL.n474 VTAIL.t8 1.38803
R935 VTAIL.n316 VTAIL.t1 1.38803
R936 VTAIL.n316 VTAIL.t4 1.38803
R937 VTAIL.n599 VTAIL.n597 1.16414
R938 VTAIL.n607 VTAIL.n566 1.16414
R939 VTAIL.n47 VTAIL.n45 1.16414
R940 VTAIL.n55 VTAIL.n14 1.16414
R941 VTAIL.n125 VTAIL.n123 1.16414
R942 VTAIL.n133 VTAIL.n92 1.16414
R943 VTAIL.n205 VTAIL.n203 1.16414
R944 VTAIL.n213 VTAIL.n172 1.16414
R945 VTAIL.n529 VTAIL.n488 1.16414
R946 VTAIL.n521 VTAIL.n520 1.16414
R947 VTAIL.n449 VTAIL.n408 1.16414
R948 VTAIL.n441 VTAIL.n440 1.16414
R949 VTAIL.n371 VTAIL.n330 1.16414
R950 VTAIL.n363 VTAIL.n362 1.16414
R951 VTAIL.n291 VTAIL.n250 1.16414
R952 VTAIL.n283 VTAIL.n282 1.16414
R953 VTAIL.n473 VTAIL.n395 0.470328
R954 VTAIL.n157 VTAIL.n79 0.470328
R955 VTAIL.n598 VTAIL.n568 0.388379
R956 VTAIL.n604 VTAIL.n603 0.388379
R957 VTAIL.n46 VTAIL.n16 0.388379
R958 VTAIL.n52 VTAIL.n51 0.388379
R959 VTAIL.n124 VTAIL.n94 0.388379
R960 VTAIL.n130 VTAIL.n129 0.388379
R961 VTAIL.n204 VTAIL.n174 0.388379
R962 VTAIL.n210 VTAIL.n209 0.388379
R963 VTAIL.n526 VTAIL.n525 0.388379
R964 VTAIL.n492 VTAIL.n490 0.388379
R965 VTAIL.n446 VTAIL.n445 0.388379
R966 VTAIL.n412 VTAIL.n410 0.388379
R967 VTAIL.n368 VTAIL.n367 0.388379
R968 VTAIL.n334 VTAIL.n332 0.388379
R969 VTAIL.n288 VTAIL.n287 0.388379
R970 VTAIL.n254 VTAIL.n252 0.388379
R971 VTAIL.n580 VTAIL.n575 0.155672
R972 VTAIL.n587 VTAIL.n575 0.155672
R973 VTAIL.n588 VTAIL.n587 0.155672
R974 VTAIL.n588 VTAIL.n571 0.155672
R975 VTAIL.n595 VTAIL.n571 0.155672
R976 VTAIL.n596 VTAIL.n595 0.155672
R977 VTAIL.n596 VTAIL.n567 0.155672
R978 VTAIL.n605 VTAIL.n567 0.155672
R979 VTAIL.n606 VTAIL.n605 0.155672
R980 VTAIL.n606 VTAIL.n563 0.155672
R981 VTAIL.n613 VTAIL.n563 0.155672
R982 VTAIL.n614 VTAIL.n613 0.155672
R983 VTAIL.n614 VTAIL.n559 0.155672
R984 VTAIL.n621 VTAIL.n559 0.155672
R985 VTAIL.n622 VTAIL.n621 0.155672
R986 VTAIL.n622 VTAIL.n555 0.155672
R987 VTAIL.n629 VTAIL.n555 0.155672
R988 VTAIL.n28 VTAIL.n23 0.155672
R989 VTAIL.n35 VTAIL.n23 0.155672
R990 VTAIL.n36 VTAIL.n35 0.155672
R991 VTAIL.n36 VTAIL.n19 0.155672
R992 VTAIL.n43 VTAIL.n19 0.155672
R993 VTAIL.n44 VTAIL.n43 0.155672
R994 VTAIL.n44 VTAIL.n15 0.155672
R995 VTAIL.n53 VTAIL.n15 0.155672
R996 VTAIL.n54 VTAIL.n53 0.155672
R997 VTAIL.n54 VTAIL.n11 0.155672
R998 VTAIL.n61 VTAIL.n11 0.155672
R999 VTAIL.n62 VTAIL.n61 0.155672
R1000 VTAIL.n62 VTAIL.n7 0.155672
R1001 VTAIL.n69 VTAIL.n7 0.155672
R1002 VTAIL.n70 VTAIL.n69 0.155672
R1003 VTAIL.n70 VTAIL.n3 0.155672
R1004 VTAIL.n77 VTAIL.n3 0.155672
R1005 VTAIL.n106 VTAIL.n101 0.155672
R1006 VTAIL.n113 VTAIL.n101 0.155672
R1007 VTAIL.n114 VTAIL.n113 0.155672
R1008 VTAIL.n114 VTAIL.n97 0.155672
R1009 VTAIL.n121 VTAIL.n97 0.155672
R1010 VTAIL.n122 VTAIL.n121 0.155672
R1011 VTAIL.n122 VTAIL.n93 0.155672
R1012 VTAIL.n131 VTAIL.n93 0.155672
R1013 VTAIL.n132 VTAIL.n131 0.155672
R1014 VTAIL.n132 VTAIL.n89 0.155672
R1015 VTAIL.n139 VTAIL.n89 0.155672
R1016 VTAIL.n140 VTAIL.n139 0.155672
R1017 VTAIL.n140 VTAIL.n85 0.155672
R1018 VTAIL.n147 VTAIL.n85 0.155672
R1019 VTAIL.n148 VTAIL.n147 0.155672
R1020 VTAIL.n148 VTAIL.n81 0.155672
R1021 VTAIL.n155 VTAIL.n81 0.155672
R1022 VTAIL.n186 VTAIL.n181 0.155672
R1023 VTAIL.n193 VTAIL.n181 0.155672
R1024 VTAIL.n194 VTAIL.n193 0.155672
R1025 VTAIL.n194 VTAIL.n177 0.155672
R1026 VTAIL.n201 VTAIL.n177 0.155672
R1027 VTAIL.n202 VTAIL.n201 0.155672
R1028 VTAIL.n202 VTAIL.n173 0.155672
R1029 VTAIL.n211 VTAIL.n173 0.155672
R1030 VTAIL.n212 VTAIL.n211 0.155672
R1031 VTAIL.n212 VTAIL.n169 0.155672
R1032 VTAIL.n219 VTAIL.n169 0.155672
R1033 VTAIL.n220 VTAIL.n219 0.155672
R1034 VTAIL.n220 VTAIL.n165 0.155672
R1035 VTAIL.n227 VTAIL.n165 0.155672
R1036 VTAIL.n228 VTAIL.n227 0.155672
R1037 VTAIL.n228 VTAIL.n161 0.155672
R1038 VTAIL.n235 VTAIL.n161 0.155672
R1039 VTAIL.n551 VTAIL.n477 0.155672
R1040 VTAIL.n544 VTAIL.n477 0.155672
R1041 VTAIL.n544 VTAIL.n543 0.155672
R1042 VTAIL.n543 VTAIL.n481 0.155672
R1043 VTAIL.n536 VTAIL.n481 0.155672
R1044 VTAIL.n536 VTAIL.n535 0.155672
R1045 VTAIL.n535 VTAIL.n485 0.155672
R1046 VTAIL.n528 VTAIL.n485 0.155672
R1047 VTAIL.n528 VTAIL.n527 0.155672
R1048 VTAIL.n527 VTAIL.n489 0.155672
R1049 VTAIL.n519 VTAIL.n489 0.155672
R1050 VTAIL.n519 VTAIL.n518 0.155672
R1051 VTAIL.n518 VTAIL.n494 0.155672
R1052 VTAIL.n511 VTAIL.n494 0.155672
R1053 VTAIL.n511 VTAIL.n510 0.155672
R1054 VTAIL.n510 VTAIL.n498 0.155672
R1055 VTAIL.n503 VTAIL.n498 0.155672
R1056 VTAIL.n471 VTAIL.n397 0.155672
R1057 VTAIL.n464 VTAIL.n397 0.155672
R1058 VTAIL.n464 VTAIL.n463 0.155672
R1059 VTAIL.n463 VTAIL.n401 0.155672
R1060 VTAIL.n456 VTAIL.n401 0.155672
R1061 VTAIL.n456 VTAIL.n455 0.155672
R1062 VTAIL.n455 VTAIL.n405 0.155672
R1063 VTAIL.n448 VTAIL.n405 0.155672
R1064 VTAIL.n448 VTAIL.n447 0.155672
R1065 VTAIL.n447 VTAIL.n409 0.155672
R1066 VTAIL.n439 VTAIL.n409 0.155672
R1067 VTAIL.n439 VTAIL.n438 0.155672
R1068 VTAIL.n438 VTAIL.n414 0.155672
R1069 VTAIL.n431 VTAIL.n414 0.155672
R1070 VTAIL.n431 VTAIL.n430 0.155672
R1071 VTAIL.n430 VTAIL.n418 0.155672
R1072 VTAIL.n423 VTAIL.n418 0.155672
R1073 VTAIL.n393 VTAIL.n319 0.155672
R1074 VTAIL.n386 VTAIL.n319 0.155672
R1075 VTAIL.n386 VTAIL.n385 0.155672
R1076 VTAIL.n385 VTAIL.n323 0.155672
R1077 VTAIL.n378 VTAIL.n323 0.155672
R1078 VTAIL.n378 VTAIL.n377 0.155672
R1079 VTAIL.n377 VTAIL.n327 0.155672
R1080 VTAIL.n370 VTAIL.n327 0.155672
R1081 VTAIL.n370 VTAIL.n369 0.155672
R1082 VTAIL.n369 VTAIL.n331 0.155672
R1083 VTAIL.n361 VTAIL.n331 0.155672
R1084 VTAIL.n361 VTAIL.n360 0.155672
R1085 VTAIL.n360 VTAIL.n336 0.155672
R1086 VTAIL.n353 VTAIL.n336 0.155672
R1087 VTAIL.n353 VTAIL.n352 0.155672
R1088 VTAIL.n352 VTAIL.n340 0.155672
R1089 VTAIL.n345 VTAIL.n340 0.155672
R1090 VTAIL.n313 VTAIL.n239 0.155672
R1091 VTAIL.n306 VTAIL.n239 0.155672
R1092 VTAIL.n306 VTAIL.n305 0.155672
R1093 VTAIL.n305 VTAIL.n243 0.155672
R1094 VTAIL.n298 VTAIL.n243 0.155672
R1095 VTAIL.n298 VTAIL.n297 0.155672
R1096 VTAIL.n297 VTAIL.n247 0.155672
R1097 VTAIL.n290 VTAIL.n247 0.155672
R1098 VTAIL.n290 VTAIL.n289 0.155672
R1099 VTAIL.n289 VTAIL.n251 0.155672
R1100 VTAIL.n281 VTAIL.n251 0.155672
R1101 VTAIL.n281 VTAIL.n280 0.155672
R1102 VTAIL.n280 VTAIL.n256 0.155672
R1103 VTAIL.n273 VTAIL.n256 0.155672
R1104 VTAIL.n273 VTAIL.n272 0.155672
R1105 VTAIL.n272 VTAIL.n260 0.155672
R1106 VTAIL.n265 VTAIL.n260 0.155672
R1107 VTAIL VTAIL.n1 0.0586897
R1108 VDD1 VDD1.n0 63.1545
R1109 VDD1.n3 VDD1.n2 63.041
R1110 VDD1.n3 VDD1.n1 63.041
R1111 VDD1.n5 VDD1.n4 61.2342
R1112 VDD1.n5 VDD1.n3 53.3587
R1113 VDD1 VDD1.n5 1.80438
R1114 VDD1.n4 VDD1.t6 1.38803
R1115 VDD1.n4 VDD1.t7 1.38803
R1116 VDD1.n0 VDD1.t0 1.38803
R1117 VDD1.n0 VDD1.t1 1.38803
R1118 VDD1.n2 VDD1.t5 1.38803
R1119 VDD1.n2 VDD1.t3 1.38803
R1120 VDD1.n1 VDD1.t4 1.38803
R1121 VDD1.n1 VDD1.t2 1.38803
R1122 B.n1111 B.n1110 585
R1123 B.n395 B.n183 585
R1124 B.n394 B.n393 585
R1125 B.n392 B.n391 585
R1126 B.n390 B.n389 585
R1127 B.n388 B.n387 585
R1128 B.n386 B.n385 585
R1129 B.n384 B.n383 585
R1130 B.n382 B.n381 585
R1131 B.n380 B.n379 585
R1132 B.n378 B.n377 585
R1133 B.n376 B.n375 585
R1134 B.n374 B.n373 585
R1135 B.n372 B.n371 585
R1136 B.n370 B.n369 585
R1137 B.n368 B.n367 585
R1138 B.n366 B.n365 585
R1139 B.n364 B.n363 585
R1140 B.n362 B.n361 585
R1141 B.n360 B.n359 585
R1142 B.n358 B.n357 585
R1143 B.n356 B.n355 585
R1144 B.n354 B.n353 585
R1145 B.n352 B.n351 585
R1146 B.n350 B.n349 585
R1147 B.n348 B.n347 585
R1148 B.n346 B.n345 585
R1149 B.n344 B.n343 585
R1150 B.n342 B.n341 585
R1151 B.n340 B.n339 585
R1152 B.n338 B.n337 585
R1153 B.n336 B.n335 585
R1154 B.n334 B.n333 585
R1155 B.n332 B.n331 585
R1156 B.n330 B.n329 585
R1157 B.n328 B.n327 585
R1158 B.n326 B.n325 585
R1159 B.n324 B.n323 585
R1160 B.n322 B.n321 585
R1161 B.n320 B.n319 585
R1162 B.n318 B.n317 585
R1163 B.n316 B.n315 585
R1164 B.n314 B.n313 585
R1165 B.n312 B.n311 585
R1166 B.n310 B.n309 585
R1167 B.n308 B.n307 585
R1168 B.n306 B.n305 585
R1169 B.n304 B.n303 585
R1170 B.n302 B.n301 585
R1171 B.n300 B.n299 585
R1172 B.n298 B.n297 585
R1173 B.n296 B.n295 585
R1174 B.n294 B.n293 585
R1175 B.n292 B.n291 585
R1176 B.n290 B.n289 585
R1177 B.n288 B.n287 585
R1178 B.n286 B.n285 585
R1179 B.n284 B.n283 585
R1180 B.n282 B.n281 585
R1181 B.n280 B.n279 585
R1182 B.n278 B.n277 585
R1183 B.n276 B.n275 585
R1184 B.n274 B.n273 585
R1185 B.n272 B.n271 585
R1186 B.n270 B.n269 585
R1187 B.n268 B.n267 585
R1188 B.n266 B.n265 585
R1189 B.n264 B.n263 585
R1190 B.n262 B.n261 585
R1191 B.n260 B.n259 585
R1192 B.n258 B.n257 585
R1193 B.n256 B.n255 585
R1194 B.n254 B.n253 585
R1195 B.n252 B.n251 585
R1196 B.n250 B.n249 585
R1197 B.n248 B.n247 585
R1198 B.n246 B.n245 585
R1199 B.n244 B.n243 585
R1200 B.n242 B.n241 585
R1201 B.n240 B.n239 585
R1202 B.n238 B.n237 585
R1203 B.n236 B.n235 585
R1204 B.n234 B.n233 585
R1205 B.n232 B.n231 585
R1206 B.n230 B.n229 585
R1207 B.n228 B.n227 585
R1208 B.n226 B.n225 585
R1209 B.n224 B.n223 585
R1210 B.n222 B.n221 585
R1211 B.n220 B.n219 585
R1212 B.n218 B.n217 585
R1213 B.n216 B.n215 585
R1214 B.n214 B.n213 585
R1215 B.n212 B.n211 585
R1216 B.n210 B.n209 585
R1217 B.n208 B.n207 585
R1218 B.n206 B.n205 585
R1219 B.n204 B.n203 585
R1220 B.n202 B.n201 585
R1221 B.n200 B.n199 585
R1222 B.n198 B.n197 585
R1223 B.n196 B.n195 585
R1224 B.n194 B.n193 585
R1225 B.n192 B.n191 585
R1226 B.n131 B.n130 585
R1227 B.n1116 B.n1115 585
R1228 B.n1109 B.n184 585
R1229 B.n184 B.n128 585
R1230 B.n1108 B.n127 585
R1231 B.n1120 B.n127 585
R1232 B.n1107 B.n126 585
R1233 B.n1121 B.n126 585
R1234 B.n1106 B.n125 585
R1235 B.n1122 B.n125 585
R1236 B.n1105 B.n1104 585
R1237 B.n1104 B.n121 585
R1238 B.n1103 B.n120 585
R1239 B.n1128 B.n120 585
R1240 B.n1102 B.n119 585
R1241 B.n1129 B.n119 585
R1242 B.n1101 B.n118 585
R1243 B.n1130 B.n118 585
R1244 B.n1100 B.n1099 585
R1245 B.n1099 B.n114 585
R1246 B.n1098 B.n113 585
R1247 B.n1136 B.n113 585
R1248 B.n1097 B.n112 585
R1249 B.n1137 B.n112 585
R1250 B.n1096 B.n111 585
R1251 B.n1138 B.n111 585
R1252 B.n1095 B.n1094 585
R1253 B.n1094 B.n107 585
R1254 B.n1093 B.n106 585
R1255 B.n1144 B.n106 585
R1256 B.n1092 B.n105 585
R1257 B.n1145 B.n105 585
R1258 B.n1091 B.n104 585
R1259 B.n1146 B.n104 585
R1260 B.n1090 B.n1089 585
R1261 B.n1089 B.n100 585
R1262 B.n1088 B.n99 585
R1263 B.n1152 B.n99 585
R1264 B.n1087 B.n98 585
R1265 B.n1153 B.n98 585
R1266 B.n1086 B.n97 585
R1267 B.n1154 B.n97 585
R1268 B.n1085 B.n1084 585
R1269 B.n1084 B.n93 585
R1270 B.n1083 B.n92 585
R1271 B.n1160 B.n92 585
R1272 B.n1082 B.n91 585
R1273 B.n1161 B.n91 585
R1274 B.n1081 B.n90 585
R1275 B.n1162 B.n90 585
R1276 B.n1080 B.n1079 585
R1277 B.n1079 B.n86 585
R1278 B.n1078 B.n85 585
R1279 B.n1168 B.n85 585
R1280 B.n1077 B.n84 585
R1281 B.n1169 B.n84 585
R1282 B.n1076 B.n83 585
R1283 B.n1170 B.n83 585
R1284 B.n1075 B.n1074 585
R1285 B.n1074 B.n79 585
R1286 B.n1073 B.n78 585
R1287 B.n1176 B.n78 585
R1288 B.n1072 B.n77 585
R1289 B.n1177 B.n77 585
R1290 B.n1071 B.n76 585
R1291 B.n1178 B.n76 585
R1292 B.n1070 B.n1069 585
R1293 B.n1069 B.n72 585
R1294 B.n1068 B.n71 585
R1295 B.n1184 B.n71 585
R1296 B.n1067 B.n70 585
R1297 B.n1185 B.n70 585
R1298 B.n1066 B.n69 585
R1299 B.n1186 B.n69 585
R1300 B.n1065 B.n1064 585
R1301 B.n1064 B.n65 585
R1302 B.n1063 B.n64 585
R1303 B.n1192 B.n64 585
R1304 B.n1062 B.n63 585
R1305 B.n1193 B.n63 585
R1306 B.n1061 B.n62 585
R1307 B.n1194 B.n62 585
R1308 B.n1060 B.n1059 585
R1309 B.n1059 B.n58 585
R1310 B.n1058 B.n57 585
R1311 B.n1200 B.n57 585
R1312 B.n1057 B.n56 585
R1313 B.n1201 B.n56 585
R1314 B.n1056 B.n55 585
R1315 B.n1202 B.n55 585
R1316 B.n1055 B.n1054 585
R1317 B.n1054 B.n51 585
R1318 B.n1053 B.n50 585
R1319 B.n1208 B.n50 585
R1320 B.n1052 B.n49 585
R1321 B.n1209 B.n49 585
R1322 B.n1051 B.n48 585
R1323 B.n1210 B.n48 585
R1324 B.n1050 B.n1049 585
R1325 B.n1049 B.n44 585
R1326 B.n1048 B.n43 585
R1327 B.n1216 B.n43 585
R1328 B.n1047 B.n42 585
R1329 B.n1217 B.n42 585
R1330 B.n1046 B.n41 585
R1331 B.n1218 B.n41 585
R1332 B.n1045 B.n1044 585
R1333 B.n1044 B.n37 585
R1334 B.n1043 B.n36 585
R1335 B.n1224 B.n36 585
R1336 B.n1042 B.n35 585
R1337 B.n1225 B.n35 585
R1338 B.n1041 B.n34 585
R1339 B.n1226 B.n34 585
R1340 B.n1040 B.n1039 585
R1341 B.n1039 B.n30 585
R1342 B.n1038 B.n29 585
R1343 B.n1232 B.n29 585
R1344 B.n1037 B.n28 585
R1345 B.n1233 B.n28 585
R1346 B.n1036 B.n27 585
R1347 B.n1234 B.n27 585
R1348 B.n1035 B.n1034 585
R1349 B.n1034 B.n23 585
R1350 B.n1033 B.n22 585
R1351 B.n1240 B.n22 585
R1352 B.n1032 B.n21 585
R1353 B.n1241 B.n21 585
R1354 B.n1031 B.n20 585
R1355 B.n1242 B.n20 585
R1356 B.n1030 B.n1029 585
R1357 B.n1029 B.n16 585
R1358 B.n1028 B.n15 585
R1359 B.n1248 B.n15 585
R1360 B.n1027 B.n14 585
R1361 B.n1249 B.n14 585
R1362 B.n1026 B.n13 585
R1363 B.n1250 B.n13 585
R1364 B.n1025 B.n1024 585
R1365 B.n1024 B.n12 585
R1366 B.n1023 B.n1022 585
R1367 B.n1023 B.n8 585
R1368 B.n1021 B.n7 585
R1369 B.n1257 B.n7 585
R1370 B.n1020 B.n6 585
R1371 B.n1258 B.n6 585
R1372 B.n1019 B.n5 585
R1373 B.n1259 B.n5 585
R1374 B.n1018 B.n1017 585
R1375 B.n1017 B.n4 585
R1376 B.n1016 B.n396 585
R1377 B.n1016 B.n1015 585
R1378 B.n1006 B.n397 585
R1379 B.n398 B.n397 585
R1380 B.n1008 B.n1007 585
R1381 B.n1009 B.n1008 585
R1382 B.n1005 B.n403 585
R1383 B.n403 B.n402 585
R1384 B.n1004 B.n1003 585
R1385 B.n1003 B.n1002 585
R1386 B.n405 B.n404 585
R1387 B.n406 B.n405 585
R1388 B.n995 B.n994 585
R1389 B.n996 B.n995 585
R1390 B.n993 B.n411 585
R1391 B.n411 B.n410 585
R1392 B.n992 B.n991 585
R1393 B.n991 B.n990 585
R1394 B.n413 B.n412 585
R1395 B.n414 B.n413 585
R1396 B.n983 B.n982 585
R1397 B.n984 B.n983 585
R1398 B.n981 B.n419 585
R1399 B.n419 B.n418 585
R1400 B.n980 B.n979 585
R1401 B.n979 B.n978 585
R1402 B.n421 B.n420 585
R1403 B.n422 B.n421 585
R1404 B.n971 B.n970 585
R1405 B.n972 B.n971 585
R1406 B.n969 B.n427 585
R1407 B.n427 B.n426 585
R1408 B.n968 B.n967 585
R1409 B.n967 B.n966 585
R1410 B.n429 B.n428 585
R1411 B.n430 B.n429 585
R1412 B.n959 B.n958 585
R1413 B.n960 B.n959 585
R1414 B.n957 B.n434 585
R1415 B.n438 B.n434 585
R1416 B.n956 B.n955 585
R1417 B.n955 B.n954 585
R1418 B.n436 B.n435 585
R1419 B.n437 B.n436 585
R1420 B.n947 B.n946 585
R1421 B.n948 B.n947 585
R1422 B.n945 B.n443 585
R1423 B.n443 B.n442 585
R1424 B.n944 B.n943 585
R1425 B.n943 B.n942 585
R1426 B.n445 B.n444 585
R1427 B.n446 B.n445 585
R1428 B.n935 B.n934 585
R1429 B.n936 B.n935 585
R1430 B.n933 B.n451 585
R1431 B.n451 B.n450 585
R1432 B.n932 B.n931 585
R1433 B.n931 B.n930 585
R1434 B.n453 B.n452 585
R1435 B.n454 B.n453 585
R1436 B.n923 B.n922 585
R1437 B.n924 B.n923 585
R1438 B.n921 B.n458 585
R1439 B.n462 B.n458 585
R1440 B.n920 B.n919 585
R1441 B.n919 B.n918 585
R1442 B.n460 B.n459 585
R1443 B.n461 B.n460 585
R1444 B.n911 B.n910 585
R1445 B.n912 B.n911 585
R1446 B.n909 B.n467 585
R1447 B.n467 B.n466 585
R1448 B.n908 B.n907 585
R1449 B.n907 B.n906 585
R1450 B.n469 B.n468 585
R1451 B.n470 B.n469 585
R1452 B.n899 B.n898 585
R1453 B.n900 B.n899 585
R1454 B.n897 B.n475 585
R1455 B.n475 B.n474 585
R1456 B.n896 B.n895 585
R1457 B.n895 B.n894 585
R1458 B.n477 B.n476 585
R1459 B.n478 B.n477 585
R1460 B.n887 B.n886 585
R1461 B.n888 B.n887 585
R1462 B.n885 B.n483 585
R1463 B.n483 B.n482 585
R1464 B.n884 B.n883 585
R1465 B.n883 B.n882 585
R1466 B.n485 B.n484 585
R1467 B.n486 B.n485 585
R1468 B.n875 B.n874 585
R1469 B.n876 B.n875 585
R1470 B.n873 B.n491 585
R1471 B.n491 B.n490 585
R1472 B.n872 B.n871 585
R1473 B.n871 B.n870 585
R1474 B.n493 B.n492 585
R1475 B.n494 B.n493 585
R1476 B.n863 B.n862 585
R1477 B.n864 B.n863 585
R1478 B.n861 B.n499 585
R1479 B.n499 B.n498 585
R1480 B.n860 B.n859 585
R1481 B.n859 B.n858 585
R1482 B.n501 B.n500 585
R1483 B.n502 B.n501 585
R1484 B.n851 B.n850 585
R1485 B.n852 B.n851 585
R1486 B.n849 B.n507 585
R1487 B.n507 B.n506 585
R1488 B.n848 B.n847 585
R1489 B.n847 B.n846 585
R1490 B.n509 B.n508 585
R1491 B.n510 B.n509 585
R1492 B.n839 B.n838 585
R1493 B.n840 B.n839 585
R1494 B.n837 B.n515 585
R1495 B.n515 B.n514 585
R1496 B.n836 B.n835 585
R1497 B.n835 B.n834 585
R1498 B.n517 B.n516 585
R1499 B.n518 B.n517 585
R1500 B.n827 B.n826 585
R1501 B.n828 B.n827 585
R1502 B.n825 B.n523 585
R1503 B.n523 B.n522 585
R1504 B.n824 B.n823 585
R1505 B.n823 B.n822 585
R1506 B.n525 B.n524 585
R1507 B.n526 B.n525 585
R1508 B.n815 B.n814 585
R1509 B.n816 B.n815 585
R1510 B.n813 B.n531 585
R1511 B.n531 B.n530 585
R1512 B.n812 B.n811 585
R1513 B.n811 B.n810 585
R1514 B.n533 B.n532 585
R1515 B.n534 B.n533 585
R1516 B.n806 B.n805 585
R1517 B.n537 B.n536 585
R1518 B.n802 B.n801 585
R1519 B.n803 B.n802 585
R1520 B.n800 B.n590 585
R1521 B.n799 B.n798 585
R1522 B.n797 B.n796 585
R1523 B.n795 B.n794 585
R1524 B.n793 B.n792 585
R1525 B.n791 B.n790 585
R1526 B.n789 B.n788 585
R1527 B.n787 B.n786 585
R1528 B.n785 B.n784 585
R1529 B.n783 B.n782 585
R1530 B.n781 B.n780 585
R1531 B.n779 B.n778 585
R1532 B.n777 B.n776 585
R1533 B.n775 B.n774 585
R1534 B.n773 B.n772 585
R1535 B.n771 B.n770 585
R1536 B.n769 B.n768 585
R1537 B.n767 B.n766 585
R1538 B.n765 B.n764 585
R1539 B.n763 B.n762 585
R1540 B.n761 B.n760 585
R1541 B.n759 B.n758 585
R1542 B.n757 B.n756 585
R1543 B.n755 B.n754 585
R1544 B.n753 B.n752 585
R1545 B.n751 B.n750 585
R1546 B.n749 B.n748 585
R1547 B.n747 B.n746 585
R1548 B.n745 B.n744 585
R1549 B.n743 B.n742 585
R1550 B.n741 B.n740 585
R1551 B.n739 B.n738 585
R1552 B.n737 B.n736 585
R1553 B.n735 B.n734 585
R1554 B.n733 B.n732 585
R1555 B.n731 B.n730 585
R1556 B.n729 B.n728 585
R1557 B.n727 B.n726 585
R1558 B.n725 B.n724 585
R1559 B.n723 B.n722 585
R1560 B.n721 B.n720 585
R1561 B.n719 B.n718 585
R1562 B.n717 B.n716 585
R1563 B.n715 B.n714 585
R1564 B.n713 B.n712 585
R1565 B.n710 B.n709 585
R1566 B.n708 B.n707 585
R1567 B.n706 B.n705 585
R1568 B.n704 B.n703 585
R1569 B.n702 B.n701 585
R1570 B.n700 B.n699 585
R1571 B.n698 B.n697 585
R1572 B.n696 B.n695 585
R1573 B.n694 B.n693 585
R1574 B.n692 B.n691 585
R1575 B.n689 B.n688 585
R1576 B.n687 B.n686 585
R1577 B.n685 B.n684 585
R1578 B.n683 B.n682 585
R1579 B.n681 B.n680 585
R1580 B.n679 B.n678 585
R1581 B.n677 B.n676 585
R1582 B.n675 B.n674 585
R1583 B.n673 B.n672 585
R1584 B.n671 B.n670 585
R1585 B.n669 B.n668 585
R1586 B.n667 B.n666 585
R1587 B.n665 B.n664 585
R1588 B.n663 B.n662 585
R1589 B.n661 B.n660 585
R1590 B.n659 B.n658 585
R1591 B.n657 B.n656 585
R1592 B.n655 B.n654 585
R1593 B.n653 B.n652 585
R1594 B.n651 B.n650 585
R1595 B.n649 B.n648 585
R1596 B.n647 B.n646 585
R1597 B.n645 B.n644 585
R1598 B.n643 B.n642 585
R1599 B.n641 B.n640 585
R1600 B.n639 B.n638 585
R1601 B.n637 B.n636 585
R1602 B.n635 B.n634 585
R1603 B.n633 B.n632 585
R1604 B.n631 B.n630 585
R1605 B.n629 B.n628 585
R1606 B.n627 B.n626 585
R1607 B.n625 B.n624 585
R1608 B.n623 B.n622 585
R1609 B.n621 B.n620 585
R1610 B.n619 B.n618 585
R1611 B.n617 B.n616 585
R1612 B.n615 B.n614 585
R1613 B.n613 B.n612 585
R1614 B.n611 B.n610 585
R1615 B.n609 B.n608 585
R1616 B.n607 B.n606 585
R1617 B.n605 B.n604 585
R1618 B.n603 B.n602 585
R1619 B.n601 B.n600 585
R1620 B.n599 B.n598 585
R1621 B.n597 B.n596 585
R1622 B.n595 B.n589 585
R1623 B.n803 B.n589 585
R1624 B.n807 B.n535 585
R1625 B.n535 B.n534 585
R1626 B.n809 B.n808 585
R1627 B.n810 B.n809 585
R1628 B.n529 B.n528 585
R1629 B.n530 B.n529 585
R1630 B.n818 B.n817 585
R1631 B.n817 B.n816 585
R1632 B.n819 B.n527 585
R1633 B.n527 B.n526 585
R1634 B.n821 B.n820 585
R1635 B.n822 B.n821 585
R1636 B.n521 B.n520 585
R1637 B.n522 B.n521 585
R1638 B.n830 B.n829 585
R1639 B.n829 B.n828 585
R1640 B.n831 B.n519 585
R1641 B.n519 B.n518 585
R1642 B.n833 B.n832 585
R1643 B.n834 B.n833 585
R1644 B.n513 B.n512 585
R1645 B.n514 B.n513 585
R1646 B.n842 B.n841 585
R1647 B.n841 B.n840 585
R1648 B.n843 B.n511 585
R1649 B.n511 B.n510 585
R1650 B.n845 B.n844 585
R1651 B.n846 B.n845 585
R1652 B.n505 B.n504 585
R1653 B.n506 B.n505 585
R1654 B.n854 B.n853 585
R1655 B.n853 B.n852 585
R1656 B.n855 B.n503 585
R1657 B.n503 B.n502 585
R1658 B.n857 B.n856 585
R1659 B.n858 B.n857 585
R1660 B.n497 B.n496 585
R1661 B.n498 B.n497 585
R1662 B.n866 B.n865 585
R1663 B.n865 B.n864 585
R1664 B.n867 B.n495 585
R1665 B.n495 B.n494 585
R1666 B.n869 B.n868 585
R1667 B.n870 B.n869 585
R1668 B.n489 B.n488 585
R1669 B.n490 B.n489 585
R1670 B.n878 B.n877 585
R1671 B.n877 B.n876 585
R1672 B.n879 B.n487 585
R1673 B.n487 B.n486 585
R1674 B.n881 B.n880 585
R1675 B.n882 B.n881 585
R1676 B.n481 B.n480 585
R1677 B.n482 B.n481 585
R1678 B.n890 B.n889 585
R1679 B.n889 B.n888 585
R1680 B.n891 B.n479 585
R1681 B.n479 B.n478 585
R1682 B.n893 B.n892 585
R1683 B.n894 B.n893 585
R1684 B.n473 B.n472 585
R1685 B.n474 B.n473 585
R1686 B.n902 B.n901 585
R1687 B.n901 B.n900 585
R1688 B.n903 B.n471 585
R1689 B.n471 B.n470 585
R1690 B.n905 B.n904 585
R1691 B.n906 B.n905 585
R1692 B.n465 B.n464 585
R1693 B.n466 B.n465 585
R1694 B.n914 B.n913 585
R1695 B.n913 B.n912 585
R1696 B.n915 B.n463 585
R1697 B.n463 B.n461 585
R1698 B.n917 B.n916 585
R1699 B.n918 B.n917 585
R1700 B.n457 B.n456 585
R1701 B.n462 B.n457 585
R1702 B.n926 B.n925 585
R1703 B.n925 B.n924 585
R1704 B.n927 B.n455 585
R1705 B.n455 B.n454 585
R1706 B.n929 B.n928 585
R1707 B.n930 B.n929 585
R1708 B.n449 B.n448 585
R1709 B.n450 B.n449 585
R1710 B.n938 B.n937 585
R1711 B.n937 B.n936 585
R1712 B.n939 B.n447 585
R1713 B.n447 B.n446 585
R1714 B.n941 B.n940 585
R1715 B.n942 B.n941 585
R1716 B.n441 B.n440 585
R1717 B.n442 B.n441 585
R1718 B.n950 B.n949 585
R1719 B.n949 B.n948 585
R1720 B.n951 B.n439 585
R1721 B.n439 B.n437 585
R1722 B.n953 B.n952 585
R1723 B.n954 B.n953 585
R1724 B.n433 B.n432 585
R1725 B.n438 B.n433 585
R1726 B.n962 B.n961 585
R1727 B.n961 B.n960 585
R1728 B.n963 B.n431 585
R1729 B.n431 B.n430 585
R1730 B.n965 B.n964 585
R1731 B.n966 B.n965 585
R1732 B.n425 B.n424 585
R1733 B.n426 B.n425 585
R1734 B.n974 B.n973 585
R1735 B.n973 B.n972 585
R1736 B.n975 B.n423 585
R1737 B.n423 B.n422 585
R1738 B.n977 B.n976 585
R1739 B.n978 B.n977 585
R1740 B.n417 B.n416 585
R1741 B.n418 B.n417 585
R1742 B.n986 B.n985 585
R1743 B.n985 B.n984 585
R1744 B.n987 B.n415 585
R1745 B.n415 B.n414 585
R1746 B.n989 B.n988 585
R1747 B.n990 B.n989 585
R1748 B.n409 B.n408 585
R1749 B.n410 B.n409 585
R1750 B.n998 B.n997 585
R1751 B.n997 B.n996 585
R1752 B.n999 B.n407 585
R1753 B.n407 B.n406 585
R1754 B.n1001 B.n1000 585
R1755 B.n1002 B.n1001 585
R1756 B.n401 B.n400 585
R1757 B.n402 B.n401 585
R1758 B.n1011 B.n1010 585
R1759 B.n1010 B.n1009 585
R1760 B.n1012 B.n399 585
R1761 B.n399 B.n398 585
R1762 B.n1014 B.n1013 585
R1763 B.n1015 B.n1014 585
R1764 B.n3 B.n0 585
R1765 B.n4 B.n3 585
R1766 B.n1256 B.n1 585
R1767 B.n1257 B.n1256 585
R1768 B.n1255 B.n1254 585
R1769 B.n1255 B.n8 585
R1770 B.n1253 B.n9 585
R1771 B.n12 B.n9 585
R1772 B.n1252 B.n1251 585
R1773 B.n1251 B.n1250 585
R1774 B.n11 B.n10 585
R1775 B.n1249 B.n11 585
R1776 B.n1247 B.n1246 585
R1777 B.n1248 B.n1247 585
R1778 B.n1245 B.n17 585
R1779 B.n17 B.n16 585
R1780 B.n1244 B.n1243 585
R1781 B.n1243 B.n1242 585
R1782 B.n19 B.n18 585
R1783 B.n1241 B.n19 585
R1784 B.n1239 B.n1238 585
R1785 B.n1240 B.n1239 585
R1786 B.n1237 B.n24 585
R1787 B.n24 B.n23 585
R1788 B.n1236 B.n1235 585
R1789 B.n1235 B.n1234 585
R1790 B.n26 B.n25 585
R1791 B.n1233 B.n26 585
R1792 B.n1231 B.n1230 585
R1793 B.n1232 B.n1231 585
R1794 B.n1229 B.n31 585
R1795 B.n31 B.n30 585
R1796 B.n1228 B.n1227 585
R1797 B.n1227 B.n1226 585
R1798 B.n33 B.n32 585
R1799 B.n1225 B.n33 585
R1800 B.n1223 B.n1222 585
R1801 B.n1224 B.n1223 585
R1802 B.n1221 B.n38 585
R1803 B.n38 B.n37 585
R1804 B.n1220 B.n1219 585
R1805 B.n1219 B.n1218 585
R1806 B.n40 B.n39 585
R1807 B.n1217 B.n40 585
R1808 B.n1215 B.n1214 585
R1809 B.n1216 B.n1215 585
R1810 B.n1213 B.n45 585
R1811 B.n45 B.n44 585
R1812 B.n1212 B.n1211 585
R1813 B.n1211 B.n1210 585
R1814 B.n47 B.n46 585
R1815 B.n1209 B.n47 585
R1816 B.n1207 B.n1206 585
R1817 B.n1208 B.n1207 585
R1818 B.n1205 B.n52 585
R1819 B.n52 B.n51 585
R1820 B.n1204 B.n1203 585
R1821 B.n1203 B.n1202 585
R1822 B.n54 B.n53 585
R1823 B.n1201 B.n54 585
R1824 B.n1199 B.n1198 585
R1825 B.n1200 B.n1199 585
R1826 B.n1197 B.n59 585
R1827 B.n59 B.n58 585
R1828 B.n1196 B.n1195 585
R1829 B.n1195 B.n1194 585
R1830 B.n61 B.n60 585
R1831 B.n1193 B.n61 585
R1832 B.n1191 B.n1190 585
R1833 B.n1192 B.n1191 585
R1834 B.n1189 B.n66 585
R1835 B.n66 B.n65 585
R1836 B.n1188 B.n1187 585
R1837 B.n1187 B.n1186 585
R1838 B.n68 B.n67 585
R1839 B.n1185 B.n68 585
R1840 B.n1183 B.n1182 585
R1841 B.n1184 B.n1183 585
R1842 B.n1181 B.n73 585
R1843 B.n73 B.n72 585
R1844 B.n1180 B.n1179 585
R1845 B.n1179 B.n1178 585
R1846 B.n75 B.n74 585
R1847 B.n1177 B.n75 585
R1848 B.n1175 B.n1174 585
R1849 B.n1176 B.n1175 585
R1850 B.n1173 B.n80 585
R1851 B.n80 B.n79 585
R1852 B.n1172 B.n1171 585
R1853 B.n1171 B.n1170 585
R1854 B.n82 B.n81 585
R1855 B.n1169 B.n82 585
R1856 B.n1167 B.n1166 585
R1857 B.n1168 B.n1167 585
R1858 B.n1165 B.n87 585
R1859 B.n87 B.n86 585
R1860 B.n1164 B.n1163 585
R1861 B.n1163 B.n1162 585
R1862 B.n89 B.n88 585
R1863 B.n1161 B.n89 585
R1864 B.n1159 B.n1158 585
R1865 B.n1160 B.n1159 585
R1866 B.n1157 B.n94 585
R1867 B.n94 B.n93 585
R1868 B.n1156 B.n1155 585
R1869 B.n1155 B.n1154 585
R1870 B.n96 B.n95 585
R1871 B.n1153 B.n96 585
R1872 B.n1151 B.n1150 585
R1873 B.n1152 B.n1151 585
R1874 B.n1149 B.n101 585
R1875 B.n101 B.n100 585
R1876 B.n1148 B.n1147 585
R1877 B.n1147 B.n1146 585
R1878 B.n103 B.n102 585
R1879 B.n1145 B.n103 585
R1880 B.n1143 B.n1142 585
R1881 B.n1144 B.n1143 585
R1882 B.n1141 B.n108 585
R1883 B.n108 B.n107 585
R1884 B.n1140 B.n1139 585
R1885 B.n1139 B.n1138 585
R1886 B.n110 B.n109 585
R1887 B.n1137 B.n110 585
R1888 B.n1135 B.n1134 585
R1889 B.n1136 B.n1135 585
R1890 B.n1133 B.n115 585
R1891 B.n115 B.n114 585
R1892 B.n1132 B.n1131 585
R1893 B.n1131 B.n1130 585
R1894 B.n117 B.n116 585
R1895 B.n1129 B.n117 585
R1896 B.n1127 B.n1126 585
R1897 B.n1128 B.n1127 585
R1898 B.n1125 B.n122 585
R1899 B.n122 B.n121 585
R1900 B.n1124 B.n1123 585
R1901 B.n1123 B.n1122 585
R1902 B.n124 B.n123 585
R1903 B.n1121 B.n124 585
R1904 B.n1119 B.n1118 585
R1905 B.n1120 B.n1119 585
R1906 B.n1117 B.n129 585
R1907 B.n129 B.n128 585
R1908 B.n1260 B.n1259 585
R1909 B.n1258 B.n2 585
R1910 B.n1115 B.n129 535.745
R1911 B.n1111 B.n184 535.745
R1912 B.n589 B.n533 535.745
R1913 B.n805 B.n535 535.745
R1914 B.n185 B.t14 405.387
R1915 B.n593 B.t21 405.387
R1916 B.n188 B.t17 405.387
R1917 B.n591 B.t11 405.387
R1918 B.n186 B.t15 321.606
R1919 B.n594 B.t20 321.606
R1920 B.n189 B.t18 321.606
R1921 B.n592 B.t10 321.606
R1922 B.n188 B.t16 295.676
R1923 B.n185 B.t12 295.676
R1924 B.n593 B.t19 295.676
R1925 B.n591 B.t8 295.676
R1926 B.n1113 B.n1112 256.663
R1927 B.n1113 B.n182 256.663
R1928 B.n1113 B.n181 256.663
R1929 B.n1113 B.n180 256.663
R1930 B.n1113 B.n179 256.663
R1931 B.n1113 B.n178 256.663
R1932 B.n1113 B.n177 256.663
R1933 B.n1113 B.n176 256.663
R1934 B.n1113 B.n175 256.663
R1935 B.n1113 B.n174 256.663
R1936 B.n1113 B.n173 256.663
R1937 B.n1113 B.n172 256.663
R1938 B.n1113 B.n171 256.663
R1939 B.n1113 B.n170 256.663
R1940 B.n1113 B.n169 256.663
R1941 B.n1113 B.n168 256.663
R1942 B.n1113 B.n167 256.663
R1943 B.n1113 B.n166 256.663
R1944 B.n1113 B.n165 256.663
R1945 B.n1113 B.n164 256.663
R1946 B.n1113 B.n163 256.663
R1947 B.n1113 B.n162 256.663
R1948 B.n1113 B.n161 256.663
R1949 B.n1113 B.n160 256.663
R1950 B.n1113 B.n159 256.663
R1951 B.n1113 B.n158 256.663
R1952 B.n1113 B.n157 256.663
R1953 B.n1113 B.n156 256.663
R1954 B.n1113 B.n155 256.663
R1955 B.n1113 B.n154 256.663
R1956 B.n1113 B.n153 256.663
R1957 B.n1113 B.n152 256.663
R1958 B.n1113 B.n151 256.663
R1959 B.n1113 B.n150 256.663
R1960 B.n1113 B.n149 256.663
R1961 B.n1113 B.n148 256.663
R1962 B.n1113 B.n147 256.663
R1963 B.n1113 B.n146 256.663
R1964 B.n1113 B.n145 256.663
R1965 B.n1113 B.n144 256.663
R1966 B.n1113 B.n143 256.663
R1967 B.n1113 B.n142 256.663
R1968 B.n1113 B.n141 256.663
R1969 B.n1113 B.n140 256.663
R1970 B.n1113 B.n139 256.663
R1971 B.n1113 B.n138 256.663
R1972 B.n1113 B.n137 256.663
R1973 B.n1113 B.n136 256.663
R1974 B.n1113 B.n135 256.663
R1975 B.n1113 B.n134 256.663
R1976 B.n1113 B.n133 256.663
R1977 B.n1113 B.n132 256.663
R1978 B.n1114 B.n1113 256.663
R1979 B.n804 B.n803 256.663
R1980 B.n803 B.n538 256.663
R1981 B.n803 B.n539 256.663
R1982 B.n803 B.n540 256.663
R1983 B.n803 B.n541 256.663
R1984 B.n803 B.n542 256.663
R1985 B.n803 B.n543 256.663
R1986 B.n803 B.n544 256.663
R1987 B.n803 B.n545 256.663
R1988 B.n803 B.n546 256.663
R1989 B.n803 B.n547 256.663
R1990 B.n803 B.n548 256.663
R1991 B.n803 B.n549 256.663
R1992 B.n803 B.n550 256.663
R1993 B.n803 B.n551 256.663
R1994 B.n803 B.n552 256.663
R1995 B.n803 B.n553 256.663
R1996 B.n803 B.n554 256.663
R1997 B.n803 B.n555 256.663
R1998 B.n803 B.n556 256.663
R1999 B.n803 B.n557 256.663
R2000 B.n803 B.n558 256.663
R2001 B.n803 B.n559 256.663
R2002 B.n803 B.n560 256.663
R2003 B.n803 B.n561 256.663
R2004 B.n803 B.n562 256.663
R2005 B.n803 B.n563 256.663
R2006 B.n803 B.n564 256.663
R2007 B.n803 B.n565 256.663
R2008 B.n803 B.n566 256.663
R2009 B.n803 B.n567 256.663
R2010 B.n803 B.n568 256.663
R2011 B.n803 B.n569 256.663
R2012 B.n803 B.n570 256.663
R2013 B.n803 B.n571 256.663
R2014 B.n803 B.n572 256.663
R2015 B.n803 B.n573 256.663
R2016 B.n803 B.n574 256.663
R2017 B.n803 B.n575 256.663
R2018 B.n803 B.n576 256.663
R2019 B.n803 B.n577 256.663
R2020 B.n803 B.n578 256.663
R2021 B.n803 B.n579 256.663
R2022 B.n803 B.n580 256.663
R2023 B.n803 B.n581 256.663
R2024 B.n803 B.n582 256.663
R2025 B.n803 B.n583 256.663
R2026 B.n803 B.n584 256.663
R2027 B.n803 B.n585 256.663
R2028 B.n803 B.n586 256.663
R2029 B.n803 B.n587 256.663
R2030 B.n803 B.n588 256.663
R2031 B.n1262 B.n1261 256.663
R2032 B.n191 B.n131 163.367
R2033 B.n195 B.n194 163.367
R2034 B.n199 B.n198 163.367
R2035 B.n203 B.n202 163.367
R2036 B.n207 B.n206 163.367
R2037 B.n211 B.n210 163.367
R2038 B.n215 B.n214 163.367
R2039 B.n219 B.n218 163.367
R2040 B.n223 B.n222 163.367
R2041 B.n227 B.n226 163.367
R2042 B.n231 B.n230 163.367
R2043 B.n235 B.n234 163.367
R2044 B.n239 B.n238 163.367
R2045 B.n243 B.n242 163.367
R2046 B.n247 B.n246 163.367
R2047 B.n251 B.n250 163.367
R2048 B.n255 B.n254 163.367
R2049 B.n259 B.n258 163.367
R2050 B.n263 B.n262 163.367
R2051 B.n267 B.n266 163.367
R2052 B.n271 B.n270 163.367
R2053 B.n275 B.n274 163.367
R2054 B.n279 B.n278 163.367
R2055 B.n283 B.n282 163.367
R2056 B.n287 B.n286 163.367
R2057 B.n291 B.n290 163.367
R2058 B.n295 B.n294 163.367
R2059 B.n299 B.n298 163.367
R2060 B.n303 B.n302 163.367
R2061 B.n307 B.n306 163.367
R2062 B.n311 B.n310 163.367
R2063 B.n315 B.n314 163.367
R2064 B.n319 B.n318 163.367
R2065 B.n323 B.n322 163.367
R2066 B.n327 B.n326 163.367
R2067 B.n331 B.n330 163.367
R2068 B.n335 B.n334 163.367
R2069 B.n339 B.n338 163.367
R2070 B.n343 B.n342 163.367
R2071 B.n347 B.n346 163.367
R2072 B.n351 B.n350 163.367
R2073 B.n355 B.n354 163.367
R2074 B.n359 B.n358 163.367
R2075 B.n363 B.n362 163.367
R2076 B.n367 B.n366 163.367
R2077 B.n371 B.n370 163.367
R2078 B.n375 B.n374 163.367
R2079 B.n379 B.n378 163.367
R2080 B.n383 B.n382 163.367
R2081 B.n387 B.n386 163.367
R2082 B.n391 B.n390 163.367
R2083 B.n393 B.n183 163.367
R2084 B.n811 B.n533 163.367
R2085 B.n811 B.n531 163.367
R2086 B.n815 B.n531 163.367
R2087 B.n815 B.n525 163.367
R2088 B.n823 B.n525 163.367
R2089 B.n823 B.n523 163.367
R2090 B.n827 B.n523 163.367
R2091 B.n827 B.n517 163.367
R2092 B.n835 B.n517 163.367
R2093 B.n835 B.n515 163.367
R2094 B.n839 B.n515 163.367
R2095 B.n839 B.n509 163.367
R2096 B.n847 B.n509 163.367
R2097 B.n847 B.n507 163.367
R2098 B.n851 B.n507 163.367
R2099 B.n851 B.n501 163.367
R2100 B.n859 B.n501 163.367
R2101 B.n859 B.n499 163.367
R2102 B.n863 B.n499 163.367
R2103 B.n863 B.n493 163.367
R2104 B.n871 B.n493 163.367
R2105 B.n871 B.n491 163.367
R2106 B.n875 B.n491 163.367
R2107 B.n875 B.n485 163.367
R2108 B.n883 B.n485 163.367
R2109 B.n883 B.n483 163.367
R2110 B.n887 B.n483 163.367
R2111 B.n887 B.n477 163.367
R2112 B.n895 B.n477 163.367
R2113 B.n895 B.n475 163.367
R2114 B.n899 B.n475 163.367
R2115 B.n899 B.n469 163.367
R2116 B.n907 B.n469 163.367
R2117 B.n907 B.n467 163.367
R2118 B.n911 B.n467 163.367
R2119 B.n911 B.n460 163.367
R2120 B.n919 B.n460 163.367
R2121 B.n919 B.n458 163.367
R2122 B.n923 B.n458 163.367
R2123 B.n923 B.n453 163.367
R2124 B.n931 B.n453 163.367
R2125 B.n931 B.n451 163.367
R2126 B.n935 B.n451 163.367
R2127 B.n935 B.n445 163.367
R2128 B.n943 B.n445 163.367
R2129 B.n943 B.n443 163.367
R2130 B.n947 B.n443 163.367
R2131 B.n947 B.n436 163.367
R2132 B.n955 B.n436 163.367
R2133 B.n955 B.n434 163.367
R2134 B.n959 B.n434 163.367
R2135 B.n959 B.n429 163.367
R2136 B.n967 B.n429 163.367
R2137 B.n967 B.n427 163.367
R2138 B.n971 B.n427 163.367
R2139 B.n971 B.n421 163.367
R2140 B.n979 B.n421 163.367
R2141 B.n979 B.n419 163.367
R2142 B.n983 B.n419 163.367
R2143 B.n983 B.n413 163.367
R2144 B.n991 B.n413 163.367
R2145 B.n991 B.n411 163.367
R2146 B.n995 B.n411 163.367
R2147 B.n995 B.n405 163.367
R2148 B.n1003 B.n405 163.367
R2149 B.n1003 B.n403 163.367
R2150 B.n1008 B.n403 163.367
R2151 B.n1008 B.n397 163.367
R2152 B.n1016 B.n397 163.367
R2153 B.n1017 B.n1016 163.367
R2154 B.n1017 B.n5 163.367
R2155 B.n6 B.n5 163.367
R2156 B.n7 B.n6 163.367
R2157 B.n1023 B.n7 163.367
R2158 B.n1024 B.n1023 163.367
R2159 B.n1024 B.n13 163.367
R2160 B.n14 B.n13 163.367
R2161 B.n15 B.n14 163.367
R2162 B.n1029 B.n15 163.367
R2163 B.n1029 B.n20 163.367
R2164 B.n21 B.n20 163.367
R2165 B.n22 B.n21 163.367
R2166 B.n1034 B.n22 163.367
R2167 B.n1034 B.n27 163.367
R2168 B.n28 B.n27 163.367
R2169 B.n29 B.n28 163.367
R2170 B.n1039 B.n29 163.367
R2171 B.n1039 B.n34 163.367
R2172 B.n35 B.n34 163.367
R2173 B.n36 B.n35 163.367
R2174 B.n1044 B.n36 163.367
R2175 B.n1044 B.n41 163.367
R2176 B.n42 B.n41 163.367
R2177 B.n43 B.n42 163.367
R2178 B.n1049 B.n43 163.367
R2179 B.n1049 B.n48 163.367
R2180 B.n49 B.n48 163.367
R2181 B.n50 B.n49 163.367
R2182 B.n1054 B.n50 163.367
R2183 B.n1054 B.n55 163.367
R2184 B.n56 B.n55 163.367
R2185 B.n57 B.n56 163.367
R2186 B.n1059 B.n57 163.367
R2187 B.n1059 B.n62 163.367
R2188 B.n63 B.n62 163.367
R2189 B.n64 B.n63 163.367
R2190 B.n1064 B.n64 163.367
R2191 B.n1064 B.n69 163.367
R2192 B.n70 B.n69 163.367
R2193 B.n71 B.n70 163.367
R2194 B.n1069 B.n71 163.367
R2195 B.n1069 B.n76 163.367
R2196 B.n77 B.n76 163.367
R2197 B.n78 B.n77 163.367
R2198 B.n1074 B.n78 163.367
R2199 B.n1074 B.n83 163.367
R2200 B.n84 B.n83 163.367
R2201 B.n85 B.n84 163.367
R2202 B.n1079 B.n85 163.367
R2203 B.n1079 B.n90 163.367
R2204 B.n91 B.n90 163.367
R2205 B.n92 B.n91 163.367
R2206 B.n1084 B.n92 163.367
R2207 B.n1084 B.n97 163.367
R2208 B.n98 B.n97 163.367
R2209 B.n99 B.n98 163.367
R2210 B.n1089 B.n99 163.367
R2211 B.n1089 B.n104 163.367
R2212 B.n105 B.n104 163.367
R2213 B.n106 B.n105 163.367
R2214 B.n1094 B.n106 163.367
R2215 B.n1094 B.n111 163.367
R2216 B.n112 B.n111 163.367
R2217 B.n113 B.n112 163.367
R2218 B.n1099 B.n113 163.367
R2219 B.n1099 B.n118 163.367
R2220 B.n119 B.n118 163.367
R2221 B.n120 B.n119 163.367
R2222 B.n1104 B.n120 163.367
R2223 B.n1104 B.n125 163.367
R2224 B.n126 B.n125 163.367
R2225 B.n127 B.n126 163.367
R2226 B.n184 B.n127 163.367
R2227 B.n802 B.n537 163.367
R2228 B.n802 B.n590 163.367
R2229 B.n798 B.n797 163.367
R2230 B.n794 B.n793 163.367
R2231 B.n790 B.n789 163.367
R2232 B.n786 B.n785 163.367
R2233 B.n782 B.n781 163.367
R2234 B.n778 B.n777 163.367
R2235 B.n774 B.n773 163.367
R2236 B.n770 B.n769 163.367
R2237 B.n766 B.n765 163.367
R2238 B.n762 B.n761 163.367
R2239 B.n758 B.n757 163.367
R2240 B.n754 B.n753 163.367
R2241 B.n750 B.n749 163.367
R2242 B.n746 B.n745 163.367
R2243 B.n742 B.n741 163.367
R2244 B.n738 B.n737 163.367
R2245 B.n734 B.n733 163.367
R2246 B.n730 B.n729 163.367
R2247 B.n726 B.n725 163.367
R2248 B.n722 B.n721 163.367
R2249 B.n718 B.n717 163.367
R2250 B.n714 B.n713 163.367
R2251 B.n709 B.n708 163.367
R2252 B.n705 B.n704 163.367
R2253 B.n701 B.n700 163.367
R2254 B.n697 B.n696 163.367
R2255 B.n693 B.n692 163.367
R2256 B.n688 B.n687 163.367
R2257 B.n684 B.n683 163.367
R2258 B.n680 B.n679 163.367
R2259 B.n676 B.n675 163.367
R2260 B.n672 B.n671 163.367
R2261 B.n668 B.n667 163.367
R2262 B.n664 B.n663 163.367
R2263 B.n660 B.n659 163.367
R2264 B.n656 B.n655 163.367
R2265 B.n652 B.n651 163.367
R2266 B.n648 B.n647 163.367
R2267 B.n644 B.n643 163.367
R2268 B.n640 B.n639 163.367
R2269 B.n636 B.n635 163.367
R2270 B.n632 B.n631 163.367
R2271 B.n628 B.n627 163.367
R2272 B.n624 B.n623 163.367
R2273 B.n620 B.n619 163.367
R2274 B.n616 B.n615 163.367
R2275 B.n612 B.n611 163.367
R2276 B.n608 B.n607 163.367
R2277 B.n604 B.n603 163.367
R2278 B.n600 B.n599 163.367
R2279 B.n596 B.n589 163.367
R2280 B.n809 B.n535 163.367
R2281 B.n809 B.n529 163.367
R2282 B.n817 B.n529 163.367
R2283 B.n817 B.n527 163.367
R2284 B.n821 B.n527 163.367
R2285 B.n821 B.n521 163.367
R2286 B.n829 B.n521 163.367
R2287 B.n829 B.n519 163.367
R2288 B.n833 B.n519 163.367
R2289 B.n833 B.n513 163.367
R2290 B.n841 B.n513 163.367
R2291 B.n841 B.n511 163.367
R2292 B.n845 B.n511 163.367
R2293 B.n845 B.n505 163.367
R2294 B.n853 B.n505 163.367
R2295 B.n853 B.n503 163.367
R2296 B.n857 B.n503 163.367
R2297 B.n857 B.n497 163.367
R2298 B.n865 B.n497 163.367
R2299 B.n865 B.n495 163.367
R2300 B.n869 B.n495 163.367
R2301 B.n869 B.n489 163.367
R2302 B.n877 B.n489 163.367
R2303 B.n877 B.n487 163.367
R2304 B.n881 B.n487 163.367
R2305 B.n881 B.n481 163.367
R2306 B.n889 B.n481 163.367
R2307 B.n889 B.n479 163.367
R2308 B.n893 B.n479 163.367
R2309 B.n893 B.n473 163.367
R2310 B.n901 B.n473 163.367
R2311 B.n901 B.n471 163.367
R2312 B.n905 B.n471 163.367
R2313 B.n905 B.n465 163.367
R2314 B.n913 B.n465 163.367
R2315 B.n913 B.n463 163.367
R2316 B.n917 B.n463 163.367
R2317 B.n917 B.n457 163.367
R2318 B.n925 B.n457 163.367
R2319 B.n925 B.n455 163.367
R2320 B.n929 B.n455 163.367
R2321 B.n929 B.n449 163.367
R2322 B.n937 B.n449 163.367
R2323 B.n937 B.n447 163.367
R2324 B.n941 B.n447 163.367
R2325 B.n941 B.n441 163.367
R2326 B.n949 B.n441 163.367
R2327 B.n949 B.n439 163.367
R2328 B.n953 B.n439 163.367
R2329 B.n953 B.n433 163.367
R2330 B.n961 B.n433 163.367
R2331 B.n961 B.n431 163.367
R2332 B.n965 B.n431 163.367
R2333 B.n965 B.n425 163.367
R2334 B.n973 B.n425 163.367
R2335 B.n973 B.n423 163.367
R2336 B.n977 B.n423 163.367
R2337 B.n977 B.n417 163.367
R2338 B.n985 B.n417 163.367
R2339 B.n985 B.n415 163.367
R2340 B.n989 B.n415 163.367
R2341 B.n989 B.n409 163.367
R2342 B.n997 B.n409 163.367
R2343 B.n997 B.n407 163.367
R2344 B.n1001 B.n407 163.367
R2345 B.n1001 B.n401 163.367
R2346 B.n1010 B.n401 163.367
R2347 B.n1010 B.n399 163.367
R2348 B.n1014 B.n399 163.367
R2349 B.n1014 B.n3 163.367
R2350 B.n1260 B.n3 163.367
R2351 B.n1256 B.n2 163.367
R2352 B.n1256 B.n1255 163.367
R2353 B.n1255 B.n9 163.367
R2354 B.n1251 B.n9 163.367
R2355 B.n1251 B.n11 163.367
R2356 B.n1247 B.n11 163.367
R2357 B.n1247 B.n17 163.367
R2358 B.n1243 B.n17 163.367
R2359 B.n1243 B.n19 163.367
R2360 B.n1239 B.n19 163.367
R2361 B.n1239 B.n24 163.367
R2362 B.n1235 B.n24 163.367
R2363 B.n1235 B.n26 163.367
R2364 B.n1231 B.n26 163.367
R2365 B.n1231 B.n31 163.367
R2366 B.n1227 B.n31 163.367
R2367 B.n1227 B.n33 163.367
R2368 B.n1223 B.n33 163.367
R2369 B.n1223 B.n38 163.367
R2370 B.n1219 B.n38 163.367
R2371 B.n1219 B.n40 163.367
R2372 B.n1215 B.n40 163.367
R2373 B.n1215 B.n45 163.367
R2374 B.n1211 B.n45 163.367
R2375 B.n1211 B.n47 163.367
R2376 B.n1207 B.n47 163.367
R2377 B.n1207 B.n52 163.367
R2378 B.n1203 B.n52 163.367
R2379 B.n1203 B.n54 163.367
R2380 B.n1199 B.n54 163.367
R2381 B.n1199 B.n59 163.367
R2382 B.n1195 B.n59 163.367
R2383 B.n1195 B.n61 163.367
R2384 B.n1191 B.n61 163.367
R2385 B.n1191 B.n66 163.367
R2386 B.n1187 B.n66 163.367
R2387 B.n1187 B.n68 163.367
R2388 B.n1183 B.n68 163.367
R2389 B.n1183 B.n73 163.367
R2390 B.n1179 B.n73 163.367
R2391 B.n1179 B.n75 163.367
R2392 B.n1175 B.n75 163.367
R2393 B.n1175 B.n80 163.367
R2394 B.n1171 B.n80 163.367
R2395 B.n1171 B.n82 163.367
R2396 B.n1167 B.n82 163.367
R2397 B.n1167 B.n87 163.367
R2398 B.n1163 B.n87 163.367
R2399 B.n1163 B.n89 163.367
R2400 B.n1159 B.n89 163.367
R2401 B.n1159 B.n94 163.367
R2402 B.n1155 B.n94 163.367
R2403 B.n1155 B.n96 163.367
R2404 B.n1151 B.n96 163.367
R2405 B.n1151 B.n101 163.367
R2406 B.n1147 B.n101 163.367
R2407 B.n1147 B.n103 163.367
R2408 B.n1143 B.n103 163.367
R2409 B.n1143 B.n108 163.367
R2410 B.n1139 B.n108 163.367
R2411 B.n1139 B.n110 163.367
R2412 B.n1135 B.n110 163.367
R2413 B.n1135 B.n115 163.367
R2414 B.n1131 B.n115 163.367
R2415 B.n1131 B.n117 163.367
R2416 B.n1127 B.n117 163.367
R2417 B.n1127 B.n122 163.367
R2418 B.n1123 B.n122 163.367
R2419 B.n1123 B.n124 163.367
R2420 B.n1119 B.n124 163.367
R2421 B.n1119 B.n129 163.367
R2422 B.n189 B.n188 83.7823
R2423 B.n186 B.n185 83.7823
R2424 B.n594 B.n593 83.7823
R2425 B.n592 B.n591 83.7823
R2426 B.n803 B.n534 74.8534
R2427 B.n1113 B.n128 74.8534
R2428 B.n1115 B.n1114 71.676
R2429 B.n191 B.n132 71.676
R2430 B.n195 B.n133 71.676
R2431 B.n199 B.n134 71.676
R2432 B.n203 B.n135 71.676
R2433 B.n207 B.n136 71.676
R2434 B.n211 B.n137 71.676
R2435 B.n215 B.n138 71.676
R2436 B.n219 B.n139 71.676
R2437 B.n223 B.n140 71.676
R2438 B.n227 B.n141 71.676
R2439 B.n231 B.n142 71.676
R2440 B.n235 B.n143 71.676
R2441 B.n239 B.n144 71.676
R2442 B.n243 B.n145 71.676
R2443 B.n247 B.n146 71.676
R2444 B.n251 B.n147 71.676
R2445 B.n255 B.n148 71.676
R2446 B.n259 B.n149 71.676
R2447 B.n263 B.n150 71.676
R2448 B.n267 B.n151 71.676
R2449 B.n271 B.n152 71.676
R2450 B.n275 B.n153 71.676
R2451 B.n279 B.n154 71.676
R2452 B.n283 B.n155 71.676
R2453 B.n287 B.n156 71.676
R2454 B.n291 B.n157 71.676
R2455 B.n295 B.n158 71.676
R2456 B.n299 B.n159 71.676
R2457 B.n303 B.n160 71.676
R2458 B.n307 B.n161 71.676
R2459 B.n311 B.n162 71.676
R2460 B.n315 B.n163 71.676
R2461 B.n319 B.n164 71.676
R2462 B.n323 B.n165 71.676
R2463 B.n327 B.n166 71.676
R2464 B.n331 B.n167 71.676
R2465 B.n335 B.n168 71.676
R2466 B.n339 B.n169 71.676
R2467 B.n343 B.n170 71.676
R2468 B.n347 B.n171 71.676
R2469 B.n351 B.n172 71.676
R2470 B.n355 B.n173 71.676
R2471 B.n359 B.n174 71.676
R2472 B.n363 B.n175 71.676
R2473 B.n367 B.n176 71.676
R2474 B.n371 B.n177 71.676
R2475 B.n375 B.n178 71.676
R2476 B.n379 B.n179 71.676
R2477 B.n383 B.n180 71.676
R2478 B.n387 B.n181 71.676
R2479 B.n391 B.n182 71.676
R2480 B.n1112 B.n183 71.676
R2481 B.n1112 B.n1111 71.676
R2482 B.n393 B.n182 71.676
R2483 B.n390 B.n181 71.676
R2484 B.n386 B.n180 71.676
R2485 B.n382 B.n179 71.676
R2486 B.n378 B.n178 71.676
R2487 B.n374 B.n177 71.676
R2488 B.n370 B.n176 71.676
R2489 B.n366 B.n175 71.676
R2490 B.n362 B.n174 71.676
R2491 B.n358 B.n173 71.676
R2492 B.n354 B.n172 71.676
R2493 B.n350 B.n171 71.676
R2494 B.n346 B.n170 71.676
R2495 B.n342 B.n169 71.676
R2496 B.n338 B.n168 71.676
R2497 B.n334 B.n167 71.676
R2498 B.n330 B.n166 71.676
R2499 B.n326 B.n165 71.676
R2500 B.n322 B.n164 71.676
R2501 B.n318 B.n163 71.676
R2502 B.n314 B.n162 71.676
R2503 B.n310 B.n161 71.676
R2504 B.n306 B.n160 71.676
R2505 B.n302 B.n159 71.676
R2506 B.n298 B.n158 71.676
R2507 B.n294 B.n157 71.676
R2508 B.n290 B.n156 71.676
R2509 B.n286 B.n155 71.676
R2510 B.n282 B.n154 71.676
R2511 B.n278 B.n153 71.676
R2512 B.n274 B.n152 71.676
R2513 B.n270 B.n151 71.676
R2514 B.n266 B.n150 71.676
R2515 B.n262 B.n149 71.676
R2516 B.n258 B.n148 71.676
R2517 B.n254 B.n147 71.676
R2518 B.n250 B.n146 71.676
R2519 B.n246 B.n145 71.676
R2520 B.n242 B.n144 71.676
R2521 B.n238 B.n143 71.676
R2522 B.n234 B.n142 71.676
R2523 B.n230 B.n141 71.676
R2524 B.n226 B.n140 71.676
R2525 B.n222 B.n139 71.676
R2526 B.n218 B.n138 71.676
R2527 B.n214 B.n137 71.676
R2528 B.n210 B.n136 71.676
R2529 B.n206 B.n135 71.676
R2530 B.n202 B.n134 71.676
R2531 B.n198 B.n133 71.676
R2532 B.n194 B.n132 71.676
R2533 B.n1114 B.n131 71.676
R2534 B.n805 B.n804 71.676
R2535 B.n590 B.n538 71.676
R2536 B.n797 B.n539 71.676
R2537 B.n793 B.n540 71.676
R2538 B.n789 B.n541 71.676
R2539 B.n785 B.n542 71.676
R2540 B.n781 B.n543 71.676
R2541 B.n777 B.n544 71.676
R2542 B.n773 B.n545 71.676
R2543 B.n769 B.n546 71.676
R2544 B.n765 B.n547 71.676
R2545 B.n761 B.n548 71.676
R2546 B.n757 B.n549 71.676
R2547 B.n753 B.n550 71.676
R2548 B.n749 B.n551 71.676
R2549 B.n745 B.n552 71.676
R2550 B.n741 B.n553 71.676
R2551 B.n737 B.n554 71.676
R2552 B.n733 B.n555 71.676
R2553 B.n729 B.n556 71.676
R2554 B.n725 B.n557 71.676
R2555 B.n721 B.n558 71.676
R2556 B.n717 B.n559 71.676
R2557 B.n713 B.n560 71.676
R2558 B.n708 B.n561 71.676
R2559 B.n704 B.n562 71.676
R2560 B.n700 B.n563 71.676
R2561 B.n696 B.n564 71.676
R2562 B.n692 B.n565 71.676
R2563 B.n687 B.n566 71.676
R2564 B.n683 B.n567 71.676
R2565 B.n679 B.n568 71.676
R2566 B.n675 B.n569 71.676
R2567 B.n671 B.n570 71.676
R2568 B.n667 B.n571 71.676
R2569 B.n663 B.n572 71.676
R2570 B.n659 B.n573 71.676
R2571 B.n655 B.n574 71.676
R2572 B.n651 B.n575 71.676
R2573 B.n647 B.n576 71.676
R2574 B.n643 B.n577 71.676
R2575 B.n639 B.n578 71.676
R2576 B.n635 B.n579 71.676
R2577 B.n631 B.n580 71.676
R2578 B.n627 B.n581 71.676
R2579 B.n623 B.n582 71.676
R2580 B.n619 B.n583 71.676
R2581 B.n615 B.n584 71.676
R2582 B.n611 B.n585 71.676
R2583 B.n607 B.n586 71.676
R2584 B.n603 B.n587 71.676
R2585 B.n599 B.n588 71.676
R2586 B.n804 B.n537 71.676
R2587 B.n798 B.n538 71.676
R2588 B.n794 B.n539 71.676
R2589 B.n790 B.n540 71.676
R2590 B.n786 B.n541 71.676
R2591 B.n782 B.n542 71.676
R2592 B.n778 B.n543 71.676
R2593 B.n774 B.n544 71.676
R2594 B.n770 B.n545 71.676
R2595 B.n766 B.n546 71.676
R2596 B.n762 B.n547 71.676
R2597 B.n758 B.n548 71.676
R2598 B.n754 B.n549 71.676
R2599 B.n750 B.n550 71.676
R2600 B.n746 B.n551 71.676
R2601 B.n742 B.n552 71.676
R2602 B.n738 B.n553 71.676
R2603 B.n734 B.n554 71.676
R2604 B.n730 B.n555 71.676
R2605 B.n726 B.n556 71.676
R2606 B.n722 B.n557 71.676
R2607 B.n718 B.n558 71.676
R2608 B.n714 B.n559 71.676
R2609 B.n709 B.n560 71.676
R2610 B.n705 B.n561 71.676
R2611 B.n701 B.n562 71.676
R2612 B.n697 B.n563 71.676
R2613 B.n693 B.n564 71.676
R2614 B.n688 B.n565 71.676
R2615 B.n684 B.n566 71.676
R2616 B.n680 B.n567 71.676
R2617 B.n676 B.n568 71.676
R2618 B.n672 B.n569 71.676
R2619 B.n668 B.n570 71.676
R2620 B.n664 B.n571 71.676
R2621 B.n660 B.n572 71.676
R2622 B.n656 B.n573 71.676
R2623 B.n652 B.n574 71.676
R2624 B.n648 B.n575 71.676
R2625 B.n644 B.n576 71.676
R2626 B.n640 B.n577 71.676
R2627 B.n636 B.n578 71.676
R2628 B.n632 B.n579 71.676
R2629 B.n628 B.n580 71.676
R2630 B.n624 B.n581 71.676
R2631 B.n620 B.n582 71.676
R2632 B.n616 B.n583 71.676
R2633 B.n612 B.n584 71.676
R2634 B.n608 B.n585 71.676
R2635 B.n604 B.n586 71.676
R2636 B.n600 B.n587 71.676
R2637 B.n596 B.n588 71.676
R2638 B.n1261 B.n1260 71.676
R2639 B.n1261 B.n2 71.676
R2640 B.n190 B.n189 59.5399
R2641 B.n187 B.n186 59.5399
R2642 B.n690 B.n594 59.5399
R2643 B.n711 B.n592 59.5399
R2644 B.n810 B.n534 38.2712
R2645 B.n810 B.n530 38.2712
R2646 B.n816 B.n530 38.2712
R2647 B.n816 B.n526 38.2712
R2648 B.n822 B.n526 38.2712
R2649 B.n822 B.n522 38.2712
R2650 B.n828 B.n522 38.2712
R2651 B.n828 B.n518 38.2712
R2652 B.n834 B.n518 38.2712
R2653 B.n840 B.n514 38.2712
R2654 B.n840 B.n510 38.2712
R2655 B.n846 B.n510 38.2712
R2656 B.n846 B.n506 38.2712
R2657 B.n852 B.n506 38.2712
R2658 B.n852 B.n502 38.2712
R2659 B.n858 B.n502 38.2712
R2660 B.n858 B.n498 38.2712
R2661 B.n864 B.n498 38.2712
R2662 B.n864 B.n494 38.2712
R2663 B.n870 B.n494 38.2712
R2664 B.n870 B.n490 38.2712
R2665 B.n876 B.n490 38.2712
R2666 B.n876 B.n486 38.2712
R2667 B.n882 B.n486 38.2712
R2668 B.n888 B.n482 38.2712
R2669 B.n888 B.n478 38.2712
R2670 B.n894 B.n478 38.2712
R2671 B.n894 B.n474 38.2712
R2672 B.n900 B.n474 38.2712
R2673 B.n900 B.n470 38.2712
R2674 B.n906 B.n470 38.2712
R2675 B.n906 B.n466 38.2712
R2676 B.n912 B.n466 38.2712
R2677 B.n912 B.n461 38.2712
R2678 B.n918 B.n461 38.2712
R2679 B.n918 B.n462 38.2712
R2680 B.n924 B.n454 38.2712
R2681 B.n930 B.n454 38.2712
R2682 B.n930 B.n450 38.2712
R2683 B.n936 B.n450 38.2712
R2684 B.n936 B.n446 38.2712
R2685 B.n942 B.n446 38.2712
R2686 B.n942 B.n442 38.2712
R2687 B.n948 B.n442 38.2712
R2688 B.n948 B.n437 38.2712
R2689 B.n954 B.n437 38.2712
R2690 B.n954 B.n438 38.2712
R2691 B.n960 B.n430 38.2712
R2692 B.n966 B.n430 38.2712
R2693 B.n966 B.n426 38.2712
R2694 B.n972 B.n426 38.2712
R2695 B.n972 B.n422 38.2712
R2696 B.n978 B.n422 38.2712
R2697 B.n978 B.n418 38.2712
R2698 B.n984 B.n418 38.2712
R2699 B.n984 B.n414 38.2712
R2700 B.n990 B.n414 38.2712
R2701 B.n990 B.n410 38.2712
R2702 B.n996 B.n410 38.2712
R2703 B.n1002 B.n406 38.2712
R2704 B.n1002 B.n402 38.2712
R2705 B.n1009 B.n402 38.2712
R2706 B.n1009 B.n398 38.2712
R2707 B.n1015 B.n398 38.2712
R2708 B.n1015 B.n4 38.2712
R2709 B.n1259 B.n4 38.2712
R2710 B.n1259 B.n1258 38.2712
R2711 B.n1258 B.n1257 38.2712
R2712 B.n1257 B.n8 38.2712
R2713 B.n12 B.n8 38.2712
R2714 B.n1250 B.n12 38.2712
R2715 B.n1250 B.n1249 38.2712
R2716 B.n1249 B.n1248 38.2712
R2717 B.n1248 B.n16 38.2712
R2718 B.n1242 B.n1241 38.2712
R2719 B.n1241 B.n1240 38.2712
R2720 B.n1240 B.n23 38.2712
R2721 B.n1234 B.n23 38.2712
R2722 B.n1234 B.n1233 38.2712
R2723 B.n1233 B.n1232 38.2712
R2724 B.n1232 B.n30 38.2712
R2725 B.n1226 B.n30 38.2712
R2726 B.n1226 B.n1225 38.2712
R2727 B.n1225 B.n1224 38.2712
R2728 B.n1224 B.n37 38.2712
R2729 B.n1218 B.n37 38.2712
R2730 B.n1217 B.n1216 38.2712
R2731 B.n1216 B.n44 38.2712
R2732 B.n1210 B.n44 38.2712
R2733 B.n1210 B.n1209 38.2712
R2734 B.n1209 B.n1208 38.2712
R2735 B.n1208 B.n51 38.2712
R2736 B.n1202 B.n51 38.2712
R2737 B.n1202 B.n1201 38.2712
R2738 B.n1201 B.n1200 38.2712
R2739 B.n1200 B.n58 38.2712
R2740 B.n1194 B.n58 38.2712
R2741 B.n1193 B.n1192 38.2712
R2742 B.n1192 B.n65 38.2712
R2743 B.n1186 B.n65 38.2712
R2744 B.n1186 B.n1185 38.2712
R2745 B.n1185 B.n1184 38.2712
R2746 B.n1184 B.n72 38.2712
R2747 B.n1178 B.n72 38.2712
R2748 B.n1178 B.n1177 38.2712
R2749 B.n1177 B.n1176 38.2712
R2750 B.n1176 B.n79 38.2712
R2751 B.n1170 B.n79 38.2712
R2752 B.n1170 B.n1169 38.2712
R2753 B.n1168 B.n86 38.2712
R2754 B.n1162 B.n86 38.2712
R2755 B.n1162 B.n1161 38.2712
R2756 B.n1161 B.n1160 38.2712
R2757 B.n1160 B.n93 38.2712
R2758 B.n1154 B.n93 38.2712
R2759 B.n1154 B.n1153 38.2712
R2760 B.n1153 B.n1152 38.2712
R2761 B.n1152 B.n100 38.2712
R2762 B.n1146 B.n100 38.2712
R2763 B.n1146 B.n1145 38.2712
R2764 B.n1145 B.n1144 38.2712
R2765 B.n1144 B.n107 38.2712
R2766 B.n1138 B.n107 38.2712
R2767 B.n1138 B.n1137 38.2712
R2768 B.n1136 B.n114 38.2712
R2769 B.n1130 B.n114 38.2712
R2770 B.n1130 B.n1129 38.2712
R2771 B.n1129 B.n1128 38.2712
R2772 B.n1128 B.n121 38.2712
R2773 B.n1122 B.n121 38.2712
R2774 B.n1122 B.n1121 38.2712
R2775 B.n1121 B.n1120 38.2712
R2776 B.n1120 B.n128 38.2712
R2777 B.n807 B.n806 34.8103
R2778 B.n595 B.n532 34.8103
R2779 B.n1110 B.n1109 34.8103
R2780 B.n1117 B.n1116 34.8103
R2781 B.n924 B.t1 33.2059
R2782 B.n1194 B.t3 33.2059
R2783 B.n438 B.t4 32.0803
R2784 B.t6 B.n1217 32.0803
R2785 B.t7 B.n482 21.9498
R2786 B.n1169 B.t2 21.9498
R2787 B.n996 B.t5 20.8242
R2788 B.n1242 B.t0 20.8242
R2789 B.n834 B.t9 19.6986
R2790 B.t13 B.n1136 19.6986
R2791 B.t9 B.n514 18.573
R2792 B.n1137 B.t13 18.573
R2793 B B.n1262 18.0485
R2794 B.t5 B.n406 17.4474
R2795 B.t0 B.n16 17.4474
R2796 B.n882 B.t7 16.3218
R2797 B.t2 B.n1168 16.3218
R2798 B.n808 B.n807 10.6151
R2799 B.n808 B.n528 10.6151
R2800 B.n818 B.n528 10.6151
R2801 B.n819 B.n818 10.6151
R2802 B.n820 B.n819 10.6151
R2803 B.n820 B.n520 10.6151
R2804 B.n830 B.n520 10.6151
R2805 B.n831 B.n830 10.6151
R2806 B.n832 B.n831 10.6151
R2807 B.n832 B.n512 10.6151
R2808 B.n842 B.n512 10.6151
R2809 B.n843 B.n842 10.6151
R2810 B.n844 B.n843 10.6151
R2811 B.n844 B.n504 10.6151
R2812 B.n854 B.n504 10.6151
R2813 B.n855 B.n854 10.6151
R2814 B.n856 B.n855 10.6151
R2815 B.n856 B.n496 10.6151
R2816 B.n866 B.n496 10.6151
R2817 B.n867 B.n866 10.6151
R2818 B.n868 B.n867 10.6151
R2819 B.n868 B.n488 10.6151
R2820 B.n878 B.n488 10.6151
R2821 B.n879 B.n878 10.6151
R2822 B.n880 B.n879 10.6151
R2823 B.n880 B.n480 10.6151
R2824 B.n890 B.n480 10.6151
R2825 B.n891 B.n890 10.6151
R2826 B.n892 B.n891 10.6151
R2827 B.n892 B.n472 10.6151
R2828 B.n902 B.n472 10.6151
R2829 B.n903 B.n902 10.6151
R2830 B.n904 B.n903 10.6151
R2831 B.n904 B.n464 10.6151
R2832 B.n914 B.n464 10.6151
R2833 B.n915 B.n914 10.6151
R2834 B.n916 B.n915 10.6151
R2835 B.n916 B.n456 10.6151
R2836 B.n926 B.n456 10.6151
R2837 B.n927 B.n926 10.6151
R2838 B.n928 B.n927 10.6151
R2839 B.n928 B.n448 10.6151
R2840 B.n938 B.n448 10.6151
R2841 B.n939 B.n938 10.6151
R2842 B.n940 B.n939 10.6151
R2843 B.n940 B.n440 10.6151
R2844 B.n950 B.n440 10.6151
R2845 B.n951 B.n950 10.6151
R2846 B.n952 B.n951 10.6151
R2847 B.n952 B.n432 10.6151
R2848 B.n962 B.n432 10.6151
R2849 B.n963 B.n962 10.6151
R2850 B.n964 B.n963 10.6151
R2851 B.n964 B.n424 10.6151
R2852 B.n974 B.n424 10.6151
R2853 B.n975 B.n974 10.6151
R2854 B.n976 B.n975 10.6151
R2855 B.n976 B.n416 10.6151
R2856 B.n986 B.n416 10.6151
R2857 B.n987 B.n986 10.6151
R2858 B.n988 B.n987 10.6151
R2859 B.n988 B.n408 10.6151
R2860 B.n998 B.n408 10.6151
R2861 B.n999 B.n998 10.6151
R2862 B.n1000 B.n999 10.6151
R2863 B.n1000 B.n400 10.6151
R2864 B.n1011 B.n400 10.6151
R2865 B.n1012 B.n1011 10.6151
R2866 B.n1013 B.n1012 10.6151
R2867 B.n1013 B.n0 10.6151
R2868 B.n806 B.n536 10.6151
R2869 B.n801 B.n536 10.6151
R2870 B.n801 B.n800 10.6151
R2871 B.n800 B.n799 10.6151
R2872 B.n799 B.n796 10.6151
R2873 B.n796 B.n795 10.6151
R2874 B.n795 B.n792 10.6151
R2875 B.n792 B.n791 10.6151
R2876 B.n791 B.n788 10.6151
R2877 B.n788 B.n787 10.6151
R2878 B.n787 B.n784 10.6151
R2879 B.n784 B.n783 10.6151
R2880 B.n783 B.n780 10.6151
R2881 B.n780 B.n779 10.6151
R2882 B.n779 B.n776 10.6151
R2883 B.n776 B.n775 10.6151
R2884 B.n775 B.n772 10.6151
R2885 B.n772 B.n771 10.6151
R2886 B.n771 B.n768 10.6151
R2887 B.n768 B.n767 10.6151
R2888 B.n767 B.n764 10.6151
R2889 B.n764 B.n763 10.6151
R2890 B.n763 B.n760 10.6151
R2891 B.n760 B.n759 10.6151
R2892 B.n759 B.n756 10.6151
R2893 B.n756 B.n755 10.6151
R2894 B.n755 B.n752 10.6151
R2895 B.n752 B.n751 10.6151
R2896 B.n751 B.n748 10.6151
R2897 B.n748 B.n747 10.6151
R2898 B.n747 B.n744 10.6151
R2899 B.n744 B.n743 10.6151
R2900 B.n743 B.n740 10.6151
R2901 B.n740 B.n739 10.6151
R2902 B.n739 B.n736 10.6151
R2903 B.n736 B.n735 10.6151
R2904 B.n735 B.n732 10.6151
R2905 B.n732 B.n731 10.6151
R2906 B.n731 B.n728 10.6151
R2907 B.n728 B.n727 10.6151
R2908 B.n727 B.n724 10.6151
R2909 B.n724 B.n723 10.6151
R2910 B.n723 B.n720 10.6151
R2911 B.n720 B.n719 10.6151
R2912 B.n719 B.n716 10.6151
R2913 B.n716 B.n715 10.6151
R2914 B.n715 B.n712 10.6151
R2915 B.n710 B.n707 10.6151
R2916 B.n707 B.n706 10.6151
R2917 B.n706 B.n703 10.6151
R2918 B.n703 B.n702 10.6151
R2919 B.n702 B.n699 10.6151
R2920 B.n699 B.n698 10.6151
R2921 B.n698 B.n695 10.6151
R2922 B.n695 B.n694 10.6151
R2923 B.n694 B.n691 10.6151
R2924 B.n689 B.n686 10.6151
R2925 B.n686 B.n685 10.6151
R2926 B.n685 B.n682 10.6151
R2927 B.n682 B.n681 10.6151
R2928 B.n681 B.n678 10.6151
R2929 B.n678 B.n677 10.6151
R2930 B.n677 B.n674 10.6151
R2931 B.n674 B.n673 10.6151
R2932 B.n673 B.n670 10.6151
R2933 B.n670 B.n669 10.6151
R2934 B.n669 B.n666 10.6151
R2935 B.n666 B.n665 10.6151
R2936 B.n665 B.n662 10.6151
R2937 B.n662 B.n661 10.6151
R2938 B.n661 B.n658 10.6151
R2939 B.n658 B.n657 10.6151
R2940 B.n657 B.n654 10.6151
R2941 B.n654 B.n653 10.6151
R2942 B.n653 B.n650 10.6151
R2943 B.n650 B.n649 10.6151
R2944 B.n649 B.n646 10.6151
R2945 B.n646 B.n645 10.6151
R2946 B.n645 B.n642 10.6151
R2947 B.n642 B.n641 10.6151
R2948 B.n641 B.n638 10.6151
R2949 B.n638 B.n637 10.6151
R2950 B.n637 B.n634 10.6151
R2951 B.n634 B.n633 10.6151
R2952 B.n633 B.n630 10.6151
R2953 B.n630 B.n629 10.6151
R2954 B.n629 B.n626 10.6151
R2955 B.n626 B.n625 10.6151
R2956 B.n625 B.n622 10.6151
R2957 B.n622 B.n621 10.6151
R2958 B.n621 B.n618 10.6151
R2959 B.n618 B.n617 10.6151
R2960 B.n617 B.n614 10.6151
R2961 B.n614 B.n613 10.6151
R2962 B.n613 B.n610 10.6151
R2963 B.n610 B.n609 10.6151
R2964 B.n609 B.n606 10.6151
R2965 B.n606 B.n605 10.6151
R2966 B.n605 B.n602 10.6151
R2967 B.n602 B.n601 10.6151
R2968 B.n601 B.n598 10.6151
R2969 B.n598 B.n597 10.6151
R2970 B.n597 B.n595 10.6151
R2971 B.n812 B.n532 10.6151
R2972 B.n813 B.n812 10.6151
R2973 B.n814 B.n813 10.6151
R2974 B.n814 B.n524 10.6151
R2975 B.n824 B.n524 10.6151
R2976 B.n825 B.n824 10.6151
R2977 B.n826 B.n825 10.6151
R2978 B.n826 B.n516 10.6151
R2979 B.n836 B.n516 10.6151
R2980 B.n837 B.n836 10.6151
R2981 B.n838 B.n837 10.6151
R2982 B.n838 B.n508 10.6151
R2983 B.n848 B.n508 10.6151
R2984 B.n849 B.n848 10.6151
R2985 B.n850 B.n849 10.6151
R2986 B.n850 B.n500 10.6151
R2987 B.n860 B.n500 10.6151
R2988 B.n861 B.n860 10.6151
R2989 B.n862 B.n861 10.6151
R2990 B.n862 B.n492 10.6151
R2991 B.n872 B.n492 10.6151
R2992 B.n873 B.n872 10.6151
R2993 B.n874 B.n873 10.6151
R2994 B.n874 B.n484 10.6151
R2995 B.n884 B.n484 10.6151
R2996 B.n885 B.n884 10.6151
R2997 B.n886 B.n885 10.6151
R2998 B.n886 B.n476 10.6151
R2999 B.n896 B.n476 10.6151
R3000 B.n897 B.n896 10.6151
R3001 B.n898 B.n897 10.6151
R3002 B.n898 B.n468 10.6151
R3003 B.n908 B.n468 10.6151
R3004 B.n909 B.n908 10.6151
R3005 B.n910 B.n909 10.6151
R3006 B.n910 B.n459 10.6151
R3007 B.n920 B.n459 10.6151
R3008 B.n921 B.n920 10.6151
R3009 B.n922 B.n921 10.6151
R3010 B.n922 B.n452 10.6151
R3011 B.n932 B.n452 10.6151
R3012 B.n933 B.n932 10.6151
R3013 B.n934 B.n933 10.6151
R3014 B.n934 B.n444 10.6151
R3015 B.n944 B.n444 10.6151
R3016 B.n945 B.n944 10.6151
R3017 B.n946 B.n945 10.6151
R3018 B.n946 B.n435 10.6151
R3019 B.n956 B.n435 10.6151
R3020 B.n957 B.n956 10.6151
R3021 B.n958 B.n957 10.6151
R3022 B.n958 B.n428 10.6151
R3023 B.n968 B.n428 10.6151
R3024 B.n969 B.n968 10.6151
R3025 B.n970 B.n969 10.6151
R3026 B.n970 B.n420 10.6151
R3027 B.n980 B.n420 10.6151
R3028 B.n981 B.n980 10.6151
R3029 B.n982 B.n981 10.6151
R3030 B.n982 B.n412 10.6151
R3031 B.n992 B.n412 10.6151
R3032 B.n993 B.n992 10.6151
R3033 B.n994 B.n993 10.6151
R3034 B.n994 B.n404 10.6151
R3035 B.n1004 B.n404 10.6151
R3036 B.n1005 B.n1004 10.6151
R3037 B.n1007 B.n1005 10.6151
R3038 B.n1007 B.n1006 10.6151
R3039 B.n1006 B.n396 10.6151
R3040 B.n1018 B.n396 10.6151
R3041 B.n1019 B.n1018 10.6151
R3042 B.n1020 B.n1019 10.6151
R3043 B.n1021 B.n1020 10.6151
R3044 B.n1022 B.n1021 10.6151
R3045 B.n1025 B.n1022 10.6151
R3046 B.n1026 B.n1025 10.6151
R3047 B.n1027 B.n1026 10.6151
R3048 B.n1028 B.n1027 10.6151
R3049 B.n1030 B.n1028 10.6151
R3050 B.n1031 B.n1030 10.6151
R3051 B.n1032 B.n1031 10.6151
R3052 B.n1033 B.n1032 10.6151
R3053 B.n1035 B.n1033 10.6151
R3054 B.n1036 B.n1035 10.6151
R3055 B.n1037 B.n1036 10.6151
R3056 B.n1038 B.n1037 10.6151
R3057 B.n1040 B.n1038 10.6151
R3058 B.n1041 B.n1040 10.6151
R3059 B.n1042 B.n1041 10.6151
R3060 B.n1043 B.n1042 10.6151
R3061 B.n1045 B.n1043 10.6151
R3062 B.n1046 B.n1045 10.6151
R3063 B.n1047 B.n1046 10.6151
R3064 B.n1048 B.n1047 10.6151
R3065 B.n1050 B.n1048 10.6151
R3066 B.n1051 B.n1050 10.6151
R3067 B.n1052 B.n1051 10.6151
R3068 B.n1053 B.n1052 10.6151
R3069 B.n1055 B.n1053 10.6151
R3070 B.n1056 B.n1055 10.6151
R3071 B.n1057 B.n1056 10.6151
R3072 B.n1058 B.n1057 10.6151
R3073 B.n1060 B.n1058 10.6151
R3074 B.n1061 B.n1060 10.6151
R3075 B.n1062 B.n1061 10.6151
R3076 B.n1063 B.n1062 10.6151
R3077 B.n1065 B.n1063 10.6151
R3078 B.n1066 B.n1065 10.6151
R3079 B.n1067 B.n1066 10.6151
R3080 B.n1068 B.n1067 10.6151
R3081 B.n1070 B.n1068 10.6151
R3082 B.n1071 B.n1070 10.6151
R3083 B.n1072 B.n1071 10.6151
R3084 B.n1073 B.n1072 10.6151
R3085 B.n1075 B.n1073 10.6151
R3086 B.n1076 B.n1075 10.6151
R3087 B.n1077 B.n1076 10.6151
R3088 B.n1078 B.n1077 10.6151
R3089 B.n1080 B.n1078 10.6151
R3090 B.n1081 B.n1080 10.6151
R3091 B.n1082 B.n1081 10.6151
R3092 B.n1083 B.n1082 10.6151
R3093 B.n1085 B.n1083 10.6151
R3094 B.n1086 B.n1085 10.6151
R3095 B.n1087 B.n1086 10.6151
R3096 B.n1088 B.n1087 10.6151
R3097 B.n1090 B.n1088 10.6151
R3098 B.n1091 B.n1090 10.6151
R3099 B.n1092 B.n1091 10.6151
R3100 B.n1093 B.n1092 10.6151
R3101 B.n1095 B.n1093 10.6151
R3102 B.n1096 B.n1095 10.6151
R3103 B.n1097 B.n1096 10.6151
R3104 B.n1098 B.n1097 10.6151
R3105 B.n1100 B.n1098 10.6151
R3106 B.n1101 B.n1100 10.6151
R3107 B.n1102 B.n1101 10.6151
R3108 B.n1103 B.n1102 10.6151
R3109 B.n1105 B.n1103 10.6151
R3110 B.n1106 B.n1105 10.6151
R3111 B.n1107 B.n1106 10.6151
R3112 B.n1108 B.n1107 10.6151
R3113 B.n1109 B.n1108 10.6151
R3114 B.n1254 B.n1 10.6151
R3115 B.n1254 B.n1253 10.6151
R3116 B.n1253 B.n1252 10.6151
R3117 B.n1252 B.n10 10.6151
R3118 B.n1246 B.n10 10.6151
R3119 B.n1246 B.n1245 10.6151
R3120 B.n1245 B.n1244 10.6151
R3121 B.n1244 B.n18 10.6151
R3122 B.n1238 B.n18 10.6151
R3123 B.n1238 B.n1237 10.6151
R3124 B.n1237 B.n1236 10.6151
R3125 B.n1236 B.n25 10.6151
R3126 B.n1230 B.n25 10.6151
R3127 B.n1230 B.n1229 10.6151
R3128 B.n1229 B.n1228 10.6151
R3129 B.n1228 B.n32 10.6151
R3130 B.n1222 B.n32 10.6151
R3131 B.n1222 B.n1221 10.6151
R3132 B.n1221 B.n1220 10.6151
R3133 B.n1220 B.n39 10.6151
R3134 B.n1214 B.n39 10.6151
R3135 B.n1214 B.n1213 10.6151
R3136 B.n1213 B.n1212 10.6151
R3137 B.n1212 B.n46 10.6151
R3138 B.n1206 B.n46 10.6151
R3139 B.n1206 B.n1205 10.6151
R3140 B.n1205 B.n1204 10.6151
R3141 B.n1204 B.n53 10.6151
R3142 B.n1198 B.n53 10.6151
R3143 B.n1198 B.n1197 10.6151
R3144 B.n1197 B.n1196 10.6151
R3145 B.n1196 B.n60 10.6151
R3146 B.n1190 B.n60 10.6151
R3147 B.n1190 B.n1189 10.6151
R3148 B.n1189 B.n1188 10.6151
R3149 B.n1188 B.n67 10.6151
R3150 B.n1182 B.n67 10.6151
R3151 B.n1182 B.n1181 10.6151
R3152 B.n1181 B.n1180 10.6151
R3153 B.n1180 B.n74 10.6151
R3154 B.n1174 B.n74 10.6151
R3155 B.n1174 B.n1173 10.6151
R3156 B.n1173 B.n1172 10.6151
R3157 B.n1172 B.n81 10.6151
R3158 B.n1166 B.n81 10.6151
R3159 B.n1166 B.n1165 10.6151
R3160 B.n1165 B.n1164 10.6151
R3161 B.n1164 B.n88 10.6151
R3162 B.n1158 B.n88 10.6151
R3163 B.n1158 B.n1157 10.6151
R3164 B.n1157 B.n1156 10.6151
R3165 B.n1156 B.n95 10.6151
R3166 B.n1150 B.n95 10.6151
R3167 B.n1150 B.n1149 10.6151
R3168 B.n1149 B.n1148 10.6151
R3169 B.n1148 B.n102 10.6151
R3170 B.n1142 B.n102 10.6151
R3171 B.n1142 B.n1141 10.6151
R3172 B.n1141 B.n1140 10.6151
R3173 B.n1140 B.n109 10.6151
R3174 B.n1134 B.n109 10.6151
R3175 B.n1134 B.n1133 10.6151
R3176 B.n1133 B.n1132 10.6151
R3177 B.n1132 B.n116 10.6151
R3178 B.n1126 B.n116 10.6151
R3179 B.n1126 B.n1125 10.6151
R3180 B.n1125 B.n1124 10.6151
R3181 B.n1124 B.n123 10.6151
R3182 B.n1118 B.n123 10.6151
R3183 B.n1118 B.n1117 10.6151
R3184 B.n1116 B.n130 10.6151
R3185 B.n192 B.n130 10.6151
R3186 B.n193 B.n192 10.6151
R3187 B.n196 B.n193 10.6151
R3188 B.n197 B.n196 10.6151
R3189 B.n200 B.n197 10.6151
R3190 B.n201 B.n200 10.6151
R3191 B.n204 B.n201 10.6151
R3192 B.n205 B.n204 10.6151
R3193 B.n208 B.n205 10.6151
R3194 B.n209 B.n208 10.6151
R3195 B.n212 B.n209 10.6151
R3196 B.n213 B.n212 10.6151
R3197 B.n216 B.n213 10.6151
R3198 B.n217 B.n216 10.6151
R3199 B.n220 B.n217 10.6151
R3200 B.n221 B.n220 10.6151
R3201 B.n224 B.n221 10.6151
R3202 B.n225 B.n224 10.6151
R3203 B.n228 B.n225 10.6151
R3204 B.n229 B.n228 10.6151
R3205 B.n232 B.n229 10.6151
R3206 B.n233 B.n232 10.6151
R3207 B.n236 B.n233 10.6151
R3208 B.n237 B.n236 10.6151
R3209 B.n240 B.n237 10.6151
R3210 B.n241 B.n240 10.6151
R3211 B.n244 B.n241 10.6151
R3212 B.n245 B.n244 10.6151
R3213 B.n248 B.n245 10.6151
R3214 B.n249 B.n248 10.6151
R3215 B.n252 B.n249 10.6151
R3216 B.n253 B.n252 10.6151
R3217 B.n256 B.n253 10.6151
R3218 B.n257 B.n256 10.6151
R3219 B.n260 B.n257 10.6151
R3220 B.n261 B.n260 10.6151
R3221 B.n264 B.n261 10.6151
R3222 B.n265 B.n264 10.6151
R3223 B.n268 B.n265 10.6151
R3224 B.n269 B.n268 10.6151
R3225 B.n272 B.n269 10.6151
R3226 B.n273 B.n272 10.6151
R3227 B.n276 B.n273 10.6151
R3228 B.n277 B.n276 10.6151
R3229 B.n280 B.n277 10.6151
R3230 B.n281 B.n280 10.6151
R3231 B.n285 B.n284 10.6151
R3232 B.n288 B.n285 10.6151
R3233 B.n289 B.n288 10.6151
R3234 B.n292 B.n289 10.6151
R3235 B.n293 B.n292 10.6151
R3236 B.n296 B.n293 10.6151
R3237 B.n297 B.n296 10.6151
R3238 B.n300 B.n297 10.6151
R3239 B.n301 B.n300 10.6151
R3240 B.n305 B.n304 10.6151
R3241 B.n308 B.n305 10.6151
R3242 B.n309 B.n308 10.6151
R3243 B.n312 B.n309 10.6151
R3244 B.n313 B.n312 10.6151
R3245 B.n316 B.n313 10.6151
R3246 B.n317 B.n316 10.6151
R3247 B.n320 B.n317 10.6151
R3248 B.n321 B.n320 10.6151
R3249 B.n324 B.n321 10.6151
R3250 B.n325 B.n324 10.6151
R3251 B.n328 B.n325 10.6151
R3252 B.n329 B.n328 10.6151
R3253 B.n332 B.n329 10.6151
R3254 B.n333 B.n332 10.6151
R3255 B.n336 B.n333 10.6151
R3256 B.n337 B.n336 10.6151
R3257 B.n340 B.n337 10.6151
R3258 B.n341 B.n340 10.6151
R3259 B.n344 B.n341 10.6151
R3260 B.n345 B.n344 10.6151
R3261 B.n348 B.n345 10.6151
R3262 B.n349 B.n348 10.6151
R3263 B.n352 B.n349 10.6151
R3264 B.n353 B.n352 10.6151
R3265 B.n356 B.n353 10.6151
R3266 B.n357 B.n356 10.6151
R3267 B.n360 B.n357 10.6151
R3268 B.n361 B.n360 10.6151
R3269 B.n364 B.n361 10.6151
R3270 B.n365 B.n364 10.6151
R3271 B.n368 B.n365 10.6151
R3272 B.n369 B.n368 10.6151
R3273 B.n372 B.n369 10.6151
R3274 B.n373 B.n372 10.6151
R3275 B.n376 B.n373 10.6151
R3276 B.n377 B.n376 10.6151
R3277 B.n380 B.n377 10.6151
R3278 B.n381 B.n380 10.6151
R3279 B.n384 B.n381 10.6151
R3280 B.n385 B.n384 10.6151
R3281 B.n388 B.n385 10.6151
R3282 B.n389 B.n388 10.6151
R3283 B.n392 B.n389 10.6151
R3284 B.n394 B.n392 10.6151
R3285 B.n395 B.n394 10.6151
R3286 B.n1110 B.n395 10.6151
R3287 B.n712 B.n711 9.36635
R3288 B.n690 B.n689 9.36635
R3289 B.n281 B.n190 9.36635
R3290 B.n304 B.n187 9.36635
R3291 B.n1262 B.n0 8.11757
R3292 B.n1262 B.n1 8.11757
R3293 B.n960 B.t4 6.19134
R3294 B.n1218 B.t6 6.19134
R3295 B.n462 B.t1 5.06573
R3296 B.t3 B.n1193 5.06573
R3297 B.n711 B.n710 1.24928
R3298 B.n691 B.n690 1.24928
R3299 B.n284 B.n190 1.24928
R3300 B.n301 B.n187 1.24928
R3301 VN.n75 VN.n39 161.3
R3302 VN.n74 VN.n73 161.3
R3303 VN.n72 VN.n40 161.3
R3304 VN.n71 VN.n70 161.3
R3305 VN.n69 VN.n41 161.3
R3306 VN.n68 VN.n67 161.3
R3307 VN.n66 VN.n42 161.3
R3308 VN.n65 VN.n64 161.3
R3309 VN.n62 VN.n43 161.3
R3310 VN.n61 VN.n60 161.3
R3311 VN.n59 VN.n44 161.3
R3312 VN.n58 VN.n57 161.3
R3313 VN.n56 VN.n45 161.3
R3314 VN.n55 VN.n54 161.3
R3315 VN.n53 VN.n46 161.3
R3316 VN.n52 VN.n51 161.3
R3317 VN.n50 VN.n47 161.3
R3318 VN.n36 VN.n0 161.3
R3319 VN.n35 VN.n34 161.3
R3320 VN.n33 VN.n1 161.3
R3321 VN.n32 VN.n31 161.3
R3322 VN.n30 VN.n2 161.3
R3323 VN.n29 VN.n28 161.3
R3324 VN.n27 VN.n3 161.3
R3325 VN.n26 VN.n25 161.3
R3326 VN.n23 VN.n4 161.3
R3327 VN.n22 VN.n21 161.3
R3328 VN.n20 VN.n5 161.3
R3329 VN.n19 VN.n18 161.3
R3330 VN.n17 VN.n6 161.3
R3331 VN.n16 VN.n15 161.3
R3332 VN.n14 VN.n7 161.3
R3333 VN.n13 VN.n12 161.3
R3334 VN.n11 VN.n8 161.3
R3335 VN.n9 VN.t7 118.239
R3336 VN.n48 VN.t3 118.239
R3337 VN.n10 VN.t4 86.1927
R3338 VN.n24 VN.t0 86.1927
R3339 VN.n37 VN.t6 86.1927
R3340 VN.n49 VN.t5 86.1927
R3341 VN.n63 VN.t2 86.1927
R3342 VN.n76 VN.t1 86.1927
R3343 VN.n10 VN.n9 67.3496
R3344 VN.n49 VN.n48 67.3496
R3345 VN VN.n77 59.4511
R3346 VN.n38 VN.n37 58.6935
R3347 VN.n77 VN.n76 58.6935
R3348 VN.n31 VN.n30 56.5193
R3349 VN.n70 VN.n69 56.5193
R3350 VN.n17 VN.n16 40.4934
R3351 VN.n18 VN.n17 40.4934
R3352 VN.n56 VN.n55 40.4934
R3353 VN.n57 VN.n56 40.4934
R3354 VN.n12 VN.n11 24.4675
R3355 VN.n12 VN.n7 24.4675
R3356 VN.n16 VN.n7 24.4675
R3357 VN.n18 VN.n5 24.4675
R3358 VN.n22 VN.n5 24.4675
R3359 VN.n23 VN.n22 24.4675
R3360 VN.n25 VN.n3 24.4675
R3361 VN.n29 VN.n3 24.4675
R3362 VN.n30 VN.n29 24.4675
R3363 VN.n31 VN.n1 24.4675
R3364 VN.n35 VN.n1 24.4675
R3365 VN.n36 VN.n35 24.4675
R3366 VN.n55 VN.n46 24.4675
R3367 VN.n51 VN.n46 24.4675
R3368 VN.n51 VN.n50 24.4675
R3369 VN.n69 VN.n68 24.4675
R3370 VN.n68 VN.n42 24.4675
R3371 VN.n64 VN.n42 24.4675
R3372 VN.n62 VN.n61 24.4675
R3373 VN.n61 VN.n44 24.4675
R3374 VN.n57 VN.n44 24.4675
R3375 VN.n75 VN.n74 24.4675
R3376 VN.n74 VN.n40 24.4675
R3377 VN.n70 VN.n40 24.4675
R3378 VN.n37 VN.n36 23.4888
R3379 VN.n76 VN.n75 23.4888
R3380 VN.n25 VN.n24 16.6381
R3381 VN.n64 VN.n63 16.6381
R3382 VN.n11 VN.n10 7.82994
R3383 VN.n24 VN.n23 7.82994
R3384 VN.n50 VN.n49 7.82994
R3385 VN.n63 VN.n62 7.82994
R3386 VN.n48 VN.n47 2.57372
R3387 VN.n9 VN.n8 2.57372
R3388 VN.n77 VN.n39 0.417535
R3389 VN.n38 VN.n0 0.417535
R3390 VN VN.n38 0.394291
R3391 VN.n73 VN.n39 0.189894
R3392 VN.n73 VN.n72 0.189894
R3393 VN.n72 VN.n71 0.189894
R3394 VN.n71 VN.n41 0.189894
R3395 VN.n67 VN.n41 0.189894
R3396 VN.n67 VN.n66 0.189894
R3397 VN.n66 VN.n65 0.189894
R3398 VN.n65 VN.n43 0.189894
R3399 VN.n60 VN.n43 0.189894
R3400 VN.n60 VN.n59 0.189894
R3401 VN.n59 VN.n58 0.189894
R3402 VN.n58 VN.n45 0.189894
R3403 VN.n54 VN.n45 0.189894
R3404 VN.n54 VN.n53 0.189894
R3405 VN.n53 VN.n52 0.189894
R3406 VN.n52 VN.n47 0.189894
R3407 VN.n13 VN.n8 0.189894
R3408 VN.n14 VN.n13 0.189894
R3409 VN.n15 VN.n14 0.189894
R3410 VN.n15 VN.n6 0.189894
R3411 VN.n19 VN.n6 0.189894
R3412 VN.n20 VN.n19 0.189894
R3413 VN.n21 VN.n20 0.189894
R3414 VN.n21 VN.n4 0.189894
R3415 VN.n26 VN.n4 0.189894
R3416 VN.n27 VN.n26 0.189894
R3417 VN.n28 VN.n27 0.189894
R3418 VN.n28 VN.n2 0.189894
R3419 VN.n32 VN.n2 0.189894
R3420 VN.n33 VN.n32 0.189894
R3421 VN.n34 VN.n33 0.189894
R3422 VN.n34 VN.n0 0.189894
R3423 VDD2.n2 VDD2.n1 63.041
R3424 VDD2.n2 VDD2.n0 63.041
R3425 VDD2 VDD2.n5 63.0381
R3426 VDD2.n4 VDD2.n3 61.2342
R3427 VDD2.n4 VDD2.n2 52.7756
R3428 VDD2 VDD2.n4 1.92076
R3429 VDD2.n5 VDD2.t2 1.38803
R3430 VDD2.n5 VDD2.t4 1.38803
R3431 VDD2.n3 VDD2.t6 1.38803
R3432 VDD2.n3 VDD2.t5 1.38803
R3433 VDD2.n1 VDD2.t7 1.38803
R3434 VDD2.n1 VDD2.t1 1.38803
R3435 VDD2.n0 VDD2.t0 1.38803
R3436 VDD2.n0 VDD2.t3 1.38803
C0 VDD1 VN 0.154396f
C1 VTAIL VDD2 9.404691f
C2 VDD1 VDD2 2.5005f
C3 VP VN 9.78361f
C4 VTAIL VDD1 9.340951f
C5 VDD2 VP 0.667736f
C6 VDD2 VN 10.9869f
C7 VTAIL VP 11.7624f
C8 VTAIL VN 11.7482f
C9 VDD1 VP 11.4982f
C10 VDD2 B 6.96879f
C11 VDD1 B 7.5541f
C12 VTAIL B 12.782788f
C13 VN B 21.060152f
C14 VP B 19.715214f
C15 VDD2.t0 B 0.303897f
C16 VDD2.t3 B 0.303897f
C17 VDD2.n0 B 2.75418f
C18 VDD2.t7 B 0.303897f
C19 VDD2.t1 B 0.303897f
C20 VDD2.n1 B 2.75418f
C21 VDD2.n2 B 4.56276f
C22 VDD2.t6 B 0.303897f
C23 VDD2.t5 B 0.303897f
C24 VDD2.n3 B 2.7336f
C25 VDD2.n4 B 3.88963f
C26 VDD2.t2 B 0.303897f
C27 VDD2.t4 B 0.303897f
C28 VDD2.n5 B 2.75413f
C29 VN.n0 B 0.030604f
C30 VN.t6 B 2.53552f
C31 VN.n1 B 0.030324f
C32 VN.n2 B 0.01627f
C33 VN.n3 B 0.030324f
C34 VN.n4 B 0.01627f
C35 VN.t0 B 2.53552f
C36 VN.n5 B 0.030324f
C37 VN.n6 B 0.01627f
C38 VN.n7 B 0.030324f
C39 VN.n8 B 0.215005f
C40 VN.t4 B 2.53552f
C41 VN.t7 B 2.80977f
C42 VN.n9 B 0.894622f
C43 VN.n10 B 0.937325f
C44 VN.n11 B 0.020143f
C45 VN.n12 B 0.030324f
C46 VN.n13 B 0.01627f
C47 VN.n14 B 0.01627f
C48 VN.n15 B 0.01627f
C49 VN.n16 B 0.032337f
C50 VN.n17 B 0.013153f
C51 VN.n18 B 0.032337f
C52 VN.n19 B 0.01627f
C53 VN.n20 B 0.01627f
C54 VN.n21 B 0.01627f
C55 VN.n22 B 0.030324f
C56 VN.n23 B 0.020143f
C57 VN.n24 B 0.88036f
C58 VN.n25 B 0.025533f
C59 VN.n26 B 0.01627f
C60 VN.n27 B 0.01627f
C61 VN.n28 B 0.01627f
C62 VN.n29 B 0.030324f
C63 VN.n30 B 0.026925f
C64 VN.n31 B 0.020578f
C65 VN.n32 B 0.01627f
C66 VN.n33 B 0.01627f
C67 VN.n34 B 0.01627f
C68 VN.n35 B 0.030324f
C69 VN.n36 B 0.029725f
C70 VN.n37 B 0.955904f
C71 VN.n38 B 0.048883f
C72 VN.n39 B 0.030604f
C73 VN.t1 B 2.53552f
C74 VN.n40 B 0.030324f
C75 VN.n41 B 0.01627f
C76 VN.n42 B 0.030324f
C77 VN.n43 B 0.01627f
C78 VN.t2 B 2.53552f
C79 VN.n44 B 0.030324f
C80 VN.n45 B 0.01627f
C81 VN.n46 B 0.030324f
C82 VN.n47 B 0.215005f
C83 VN.t5 B 2.53552f
C84 VN.t3 B 2.80977f
C85 VN.n48 B 0.894622f
C86 VN.n49 B 0.937325f
C87 VN.n50 B 0.020143f
C88 VN.n51 B 0.030324f
C89 VN.n52 B 0.01627f
C90 VN.n53 B 0.01627f
C91 VN.n54 B 0.01627f
C92 VN.n55 B 0.032337f
C93 VN.n56 B 0.013153f
C94 VN.n57 B 0.032337f
C95 VN.n58 B 0.01627f
C96 VN.n59 B 0.01627f
C97 VN.n60 B 0.01627f
C98 VN.n61 B 0.030324f
C99 VN.n62 B 0.020143f
C100 VN.n63 B 0.88036f
C101 VN.n64 B 0.025533f
C102 VN.n65 B 0.01627f
C103 VN.n66 B 0.01627f
C104 VN.n67 B 0.01627f
C105 VN.n68 B 0.030324f
C106 VN.n69 B 0.026925f
C107 VN.n70 B 0.020578f
C108 VN.n71 B 0.01627f
C109 VN.n72 B 0.01627f
C110 VN.n73 B 0.01627f
C111 VN.n74 B 0.030324f
C112 VN.n75 B 0.029725f
C113 VN.n76 B 0.955904f
C114 VN.n77 B 1.19969f
C115 VDD1.t0 B 0.307867f
C116 VDD1.t1 B 0.307867f
C117 VDD1.n0 B 2.79172f
C118 VDD1.t4 B 0.307867f
C119 VDD1.t2 B 0.307867f
C120 VDD1.n1 B 2.79016f
C121 VDD1.t5 B 0.307867f
C122 VDD1.t3 B 0.307867f
C123 VDD1.n2 B 2.79016f
C124 VDD1.n3 B 4.67839f
C125 VDD1.t6 B 0.307867f
C126 VDD1.t7 B 0.307867f
C127 VDD1.n4 B 2.76931f
C128 VDD1.n5 B 3.97503f
C129 VTAIL.t6 B 0.22693f
C130 VTAIL.t3 B 0.22693f
C131 VTAIL.n0 B 1.97936f
C132 VTAIL.n1 B 0.449029f
C133 VTAIL.n2 B 0.02978f
C134 VTAIL.n3 B 0.020124f
C135 VTAIL.n4 B 0.010814f
C136 VTAIL.n5 B 0.02556f
C137 VTAIL.n6 B 0.01145f
C138 VTAIL.n7 B 0.020124f
C139 VTAIL.n8 B 0.010814f
C140 VTAIL.n9 B 0.02556f
C141 VTAIL.n10 B 0.01145f
C142 VTAIL.n11 B 0.020124f
C143 VTAIL.n12 B 0.010814f
C144 VTAIL.n13 B 0.02556f
C145 VTAIL.n14 B 0.01145f
C146 VTAIL.n15 B 0.020124f
C147 VTAIL.n16 B 0.011132f
C148 VTAIL.n17 B 0.02556f
C149 VTAIL.n18 B 0.01145f
C150 VTAIL.n19 B 0.020124f
C151 VTAIL.n20 B 0.010814f
C152 VTAIL.n21 B 0.02556f
C153 VTAIL.n22 B 0.01145f
C154 VTAIL.n23 B 0.020124f
C155 VTAIL.n24 B 0.010814f
C156 VTAIL.n25 B 0.01917f
C157 VTAIL.n26 B 0.018069f
C158 VTAIL.t0 B 0.043415f
C159 VTAIL.n27 B 0.162629f
C160 VTAIL.n28 B 1.21841f
C161 VTAIL.n29 B 0.010814f
C162 VTAIL.n30 B 0.01145f
C163 VTAIL.n31 B 0.02556f
C164 VTAIL.n32 B 0.02556f
C165 VTAIL.n33 B 0.01145f
C166 VTAIL.n34 B 0.010814f
C167 VTAIL.n35 B 0.020124f
C168 VTAIL.n36 B 0.020124f
C169 VTAIL.n37 B 0.010814f
C170 VTAIL.n38 B 0.01145f
C171 VTAIL.n39 B 0.02556f
C172 VTAIL.n40 B 0.02556f
C173 VTAIL.n41 B 0.01145f
C174 VTAIL.n42 B 0.010814f
C175 VTAIL.n43 B 0.020124f
C176 VTAIL.n44 B 0.020124f
C177 VTAIL.n45 B 0.010814f
C178 VTAIL.n46 B 0.010814f
C179 VTAIL.n47 B 0.01145f
C180 VTAIL.n48 B 0.02556f
C181 VTAIL.n49 B 0.02556f
C182 VTAIL.n50 B 0.02556f
C183 VTAIL.n51 B 0.011132f
C184 VTAIL.n52 B 0.010814f
C185 VTAIL.n53 B 0.020124f
C186 VTAIL.n54 B 0.020124f
C187 VTAIL.n55 B 0.010814f
C188 VTAIL.n56 B 0.01145f
C189 VTAIL.n57 B 0.02556f
C190 VTAIL.n58 B 0.02556f
C191 VTAIL.n59 B 0.01145f
C192 VTAIL.n60 B 0.010814f
C193 VTAIL.n61 B 0.020124f
C194 VTAIL.n62 B 0.020124f
C195 VTAIL.n63 B 0.010814f
C196 VTAIL.n64 B 0.01145f
C197 VTAIL.n65 B 0.02556f
C198 VTAIL.n66 B 0.02556f
C199 VTAIL.n67 B 0.01145f
C200 VTAIL.n68 B 0.010814f
C201 VTAIL.n69 B 0.020124f
C202 VTAIL.n70 B 0.020124f
C203 VTAIL.n71 B 0.010814f
C204 VTAIL.n72 B 0.01145f
C205 VTAIL.n73 B 0.02556f
C206 VTAIL.n74 B 0.057974f
C207 VTAIL.n75 B 0.01145f
C208 VTAIL.n76 B 0.010814f
C209 VTAIL.n77 B 0.046241f
C210 VTAIL.n78 B 0.032702f
C211 VTAIL.n79 B 0.288986f
C212 VTAIL.n80 B 0.02978f
C213 VTAIL.n81 B 0.020124f
C214 VTAIL.n82 B 0.010814f
C215 VTAIL.n83 B 0.02556f
C216 VTAIL.n84 B 0.01145f
C217 VTAIL.n85 B 0.020124f
C218 VTAIL.n86 B 0.010814f
C219 VTAIL.n87 B 0.02556f
C220 VTAIL.n88 B 0.01145f
C221 VTAIL.n89 B 0.020124f
C222 VTAIL.n90 B 0.010814f
C223 VTAIL.n91 B 0.02556f
C224 VTAIL.n92 B 0.01145f
C225 VTAIL.n93 B 0.020124f
C226 VTAIL.n94 B 0.011132f
C227 VTAIL.n95 B 0.02556f
C228 VTAIL.n96 B 0.01145f
C229 VTAIL.n97 B 0.020124f
C230 VTAIL.n98 B 0.010814f
C231 VTAIL.n99 B 0.02556f
C232 VTAIL.n100 B 0.01145f
C233 VTAIL.n101 B 0.020124f
C234 VTAIL.n102 B 0.010814f
C235 VTAIL.n103 B 0.01917f
C236 VTAIL.n104 B 0.018069f
C237 VTAIL.t15 B 0.043415f
C238 VTAIL.n105 B 0.162629f
C239 VTAIL.n106 B 1.21841f
C240 VTAIL.n107 B 0.010814f
C241 VTAIL.n108 B 0.01145f
C242 VTAIL.n109 B 0.02556f
C243 VTAIL.n110 B 0.02556f
C244 VTAIL.n111 B 0.01145f
C245 VTAIL.n112 B 0.010814f
C246 VTAIL.n113 B 0.020124f
C247 VTAIL.n114 B 0.020124f
C248 VTAIL.n115 B 0.010814f
C249 VTAIL.n116 B 0.01145f
C250 VTAIL.n117 B 0.02556f
C251 VTAIL.n118 B 0.02556f
C252 VTAIL.n119 B 0.01145f
C253 VTAIL.n120 B 0.010814f
C254 VTAIL.n121 B 0.020124f
C255 VTAIL.n122 B 0.020124f
C256 VTAIL.n123 B 0.010814f
C257 VTAIL.n124 B 0.010814f
C258 VTAIL.n125 B 0.01145f
C259 VTAIL.n126 B 0.02556f
C260 VTAIL.n127 B 0.02556f
C261 VTAIL.n128 B 0.02556f
C262 VTAIL.n129 B 0.011132f
C263 VTAIL.n130 B 0.010814f
C264 VTAIL.n131 B 0.020124f
C265 VTAIL.n132 B 0.020124f
C266 VTAIL.n133 B 0.010814f
C267 VTAIL.n134 B 0.01145f
C268 VTAIL.n135 B 0.02556f
C269 VTAIL.n136 B 0.02556f
C270 VTAIL.n137 B 0.01145f
C271 VTAIL.n138 B 0.010814f
C272 VTAIL.n139 B 0.020124f
C273 VTAIL.n140 B 0.020124f
C274 VTAIL.n141 B 0.010814f
C275 VTAIL.n142 B 0.01145f
C276 VTAIL.n143 B 0.02556f
C277 VTAIL.n144 B 0.02556f
C278 VTAIL.n145 B 0.01145f
C279 VTAIL.n146 B 0.010814f
C280 VTAIL.n147 B 0.020124f
C281 VTAIL.n148 B 0.020124f
C282 VTAIL.n149 B 0.010814f
C283 VTAIL.n150 B 0.01145f
C284 VTAIL.n151 B 0.02556f
C285 VTAIL.n152 B 0.057974f
C286 VTAIL.n153 B 0.01145f
C287 VTAIL.n154 B 0.010814f
C288 VTAIL.n155 B 0.046241f
C289 VTAIL.n156 B 0.032702f
C290 VTAIL.n157 B 0.288986f
C291 VTAIL.t10 B 0.22693f
C292 VTAIL.t11 B 0.22693f
C293 VTAIL.n158 B 1.97936f
C294 VTAIL.n159 B 0.686744f
C295 VTAIL.n160 B 0.02978f
C296 VTAIL.n161 B 0.020124f
C297 VTAIL.n162 B 0.010814f
C298 VTAIL.n163 B 0.02556f
C299 VTAIL.n164 B 0.01145f
C300 VTAIL.n165 B 0.020124f
C301 VTAIL.n166 B 0.010814f
C302 VTAIL.n167 B 0.02556f
C303 VTAIL.n168 B 0.01145f
C304 VTAIL.n169 B 0.020124f
C305 VTAIL.n170 B 0.010814f
C306 VTAIL.n171 B 0.02556f
C307 VTAIL.n172 B 0.01145f
C308 VTAIL.n173 B 0.020124f
C309 VTAIL.n174 B 0.011132f
C310 VTAIL.n175 B 0.02556f
C311 VTAIL.n176 B 0.01145f
C312 VTAIL.n177 B 0.020124f
C313 VTAIL.n178 B 0.010814f
C314 VTAIL.n179 B 0.02556f
C315 VTAIL.n180 B 0.01145f
C316 VTAIL.n181 B 0.020124f
C317 VTAIL.n182 B 0.010814f
C318 VTAIL.n183 B 0.01917f
C319 VTAIL.n184 B 0.018069f
C320 VTAIL.t13 B 0.043415f
C321 VTAIL.n185 B 0.162629f
C322 VTAIL.n186 B 1.21841f
C323 VTAIL.n187 B 0.010814f
C324 VTAIL.n188 B 0.01145f
C325 VTAIL.n189 B 0.02556f
C326 VTAIL.n190 B 0.02556f
C327 VTAIL.n191 B 0.01145f
C328 VTAIL.n192 B 0.010814f
C329 VTAIL.n193 B 0.020124f
C330 VTAIL.n194 B 0.020124f
C331 VTAIL.n195 B 0.010814f
C332 VTAIL.n196 B 0.01145f
C333 VTAIL.n197 B 0.02556f
C334 VTAIL.n198 B 0.02556f
C335 VTAIL.n199 B 0.01145f
C336 VTAIL.n200 B 0.010814f
C337 VTAIL.n201 B 0.020124f
C338 VTAIL.n202 B 0.020124f
C339 VTAIL.n203 B 0.010814f
C340 VTAIL.n204 B 0.010814f
C341 VTAIL.n205 B 0.01145f
C342 VTAIL.n206 B 0.02556f
C343 VTAIL.n207 B 0.02556f
C344 VTAIL.n208 B 0.02556f
C345 VTAIL.n209 B 0.011132f
C346 VTAIL.n210 B 0.010814f
C347 VTAIL.n211 B 0.020124f
C348 VTAIL.n212 B 0.020124f
C349 VTAIL.n213 B 0.010814f
C350 VTAIL.n214 B 0.01145f
C351 VTAIL.n215 B 0.02556f
C352 VTAIL.n216 B 0.02556f
C353 VTAIL.n217 B 0.01145f
C354 VTAIL.n218 B 0.010814f
C355 VTAIL.n219 B 0.020124f
C356 VTAIL.n220 B 0.020124f
C357 VTAIL.n221 B 0.010814f
C358 VTAIL.n222 B 0.01145f
C359 VTAIL.n223 B 0.02556f
C360 VTAIL.n224 B 0.02556f
C361 VTAIL.n225 B 0.01145f
C362 VTAIL.n226 B 0.010814f
C363 VTAIL.n227 B 0.020124f
C364 VTAIL.n228 B 0.020124f
C365 VTAIL.n229 B 0.010814f
C366 VTAIL.n230 B 0.01145f
C367 VTAIL.n231 B 0.02556f
C368 VTAIL.n232 B 0.057974f
C369 VTAIL.n233 B 0.01145f
C370 VTAIL.n234 B 0.010814f
C371 VTAIL.n235 B 0.046241f
C372 VTAIL.n236 B 0.032702f
C373 VTAIL.n237 B 1.57106f
C374 VTAIL.n238 B 0.02978f
C375 VTAIL.n239 B 0.020124f
C376 VTAIL.n240 B 0.010814f
C377 VTAIL.n241 B 0.02556f
C378 VTAIL.n242 B 0.01145f
C379 VTAIL.n243 B 0.020124f
C380 VTAIL.n244 B 0.010814f
C381 VTAIL.n245 B 0.02556f
C382 VTAIL.n246 B 0.01145f
C383 VTAIL.n247 B 0.020124f
C384 VTAIL.n248 B 0.010814f
C385 VTAIL.n249 B 0.02556f
C386 VTAIL.n250 B 0.01145f
C387 VTAIL.n251 B 0.020124f
C388 VTAIL.n252 B 0.011132f
C389 VTAIL.n253 B 0.02556f
C390 VTAIL.n254 B 0.010814f
C391 VTAIL.n255 B 0.01145f
C392 VTAIL.n256 B 0.020124f
C393 VTAIL.n257 B 0.010814f
C394 VTAIL.n258 B 0.02556f
C395 VTAIL.n259 B 0.01145f
C396 VTAIL.n260 B 0.020124f
C397 VTAIL.n261 B 0.010814f
C398 VTAIL.n262 B 0.01917f
C399 VTAIL.n263 B 0.018069f
C400 VTAIL.t7 B 0.043415f
C401 VTAIL.n264 B 0.162629f
C402 VTAIL.n265 B 1.21841f
C403 VTAIL.n266 B 0.010814f
C404 VTAIL.n267 B 0.01145f
C405 VTAIL.n268 B 0.02556f
C406 VTAIL.n269 B 0.02556f
C407 VTAIL.n270 B 0.01145f
C408 VTAIL.n271 B 0.010814f
C409 VTAIL.n272 B 0.020124f
C410 VTAIL.n273 B 0.020124f
C411 VTAIL.n274 B 0.010814f
C412 VTAIL.n275 B 0.01145f
C413 VTAIL.n276 B 0.02556f
C414 VTAIL.n277 B 0.02556f
C415 VTAIL.n278 B 0.01145f
C416 VTAIL.n279 B 0.010814f
C417 VTAIL.n280 B 0.020124f
C418 VTAIL.n281 B 0.020124f
C419 VTAIL.n282 B 0.010814f
C420 VTAIL.n283 B 0.01145f
C421 VTAIL.n284 B 0.02556f
C422 VTAIL.n285 B 0.02556f
C423 VTAIL.n286 B 0.02556f
C424 VTAIL.n287 B 0.011132f
C425 VTAIL.n288 B 0.010814f
C426 VTAIL.n289 B 0.020124f
C427 VTAIL.n290 B 0.020124f
C428 VTAIL.n291 B 0.010814f
C429 VTAIL.n292 B 0.01145f
C430 VTAIL.n293 B 0.02556f
C431 VTAIL.n294 B 0.02556f
C432 VTAIL.n295 B 0.01145f
C433 VTAIL.n296 B 0.010814f
C434 VTAIL.n297 B 0.020124f
C435 VTAIL.n298 B 0.020124f
C436 VTAIL.n299 B 0.010814f
C437 VTAIL.n300 B 0.01145f
C438 VTAIL.n301 B 0.02556f
C439 VTAIL.n302 B 0.02556f
C440 VTAIL.n303 B 0.01145f
C441 VTAIL.n304 B 0.010814f
C442 VTAIL.n305 B 0.020124f
C443 VTAIL.n306 B 0.020124f
C444 VTAIL.n307 B 0.010814f
C445 VTAIL.n308 B 0.01145f
C446 VTAIL.n309 B 0.02556f
C447 VTAIL.n310 B 0.057974f
C448 VTAIL.n311 B 0.01145f
C449 VTAIL.n312 B 0.010814f
C450 VTAIL.n313 B 0.046241f
C451 VTAIL.n314 B 0.032702f
C452 VTAIL.n315 B 1.57106f
C453 VTAIL.t1 B 0.22693f
C454 VTAIL.t4 B 0.22693f
C455 VTAIL.n316 B 1.97936f
C456 VTAIL.n317 B 0.686741f
C457 VTAIL.n318 B 0.02978f
C458 VTAIL.n319 B 0.020124f
C459 VTAIL.n320 B 0.010814f
C460 VTAIL.n321 B 0.02556f
C461 VTAIL.n322 B 0.01145f
C462 VTAIL.n323 B 0.020124f
C463 VTAIL.n324 B 0.010814f
C464 VTAIL.n325 B 0.02556f
C465 VTAIL.n326 B 0.01145f
C466 VTAIL.n327 B 0.020124f
C467 VTAIL.n328 B 0.010814f
C468 VTAIL.n329 B 0.02556f
C469 VTAIL.n330 B 0.01145f
C470 VTAIL.n331 B 0.020124f
C471 VTAIL.n332 B 0.011132f
C472 VTAIL.n333 B 0.02556f
C473 VTAIL.n334 B 0.010814f
C474 VTAIL.n335 B 0.01145f
C475 VTAIL.n336 B 0.020124f
C476 VTAIL.n337 B 0.010814f
C477 VTAIL.n338 B 0.02556f
C478 VTAIL.n339 B 0.01145f
C479 VTAIL.n340 B 0.020124f
C480 VTAIL.n341 B 0.010814f
C481 VTAIL.n342 B 0.01917f
C482 VTAIL.n343 B 0.018069f
C483 VTAIL.t5 B 0.043415f
C484 VTAIL.n344 B 0.162629f
C485 VTAIL.n345 B 1.21841f
C486 VTAIL.n346 B 0.010814f
C487 VTAIL.n347 B 0.01145f
C488 VTAIL.n348 B 0.02556f
C489 VTAIL.n349 B 0.02556f
C490 VTAIL.n350 B 0.01145f
C491 VTAIL.n351 B 0.010814f
C492 VTAIL.n352 B 0.020124f
C493 VTAIL.n353 B 0.020124f
C494 VTAIL.n354 B 0.010814f
C495 VTAIL.n355 B 0.01145f
C496 VTAIL.n356 B 0.02556f
C497 VTAIL.n357 B 0.02556f
C498 VTAIL.n358 B 0.01145f
C499 VTAIL.n359 B 0.010814f
C500 VTAIL.n360 B 0.020124f
C501 VTAIL.n361 B 0.020124f
C502 VTAIL.n362 B 0.010814f
C503 VTAIL.n363 B 0.01145f
C504 VTAIL.n364 B 0.02556f
C505 VTAIL.n365 B 0.02556f
C506 VTAIL.n366 B 0.02556f
C507 VTAIL.n367 B 0.011132f
C508 VTAIL.n368 B 0.010814f
C509 VTAIL.n369 B 0.020124f
C510 VTAIL.n370 B 0.020124f
C511 VTAIL.n371 B 0.010814f
C512 VTAIL.n372 B 0.01145f
C513 VTAIL.n373 B 0.02556f
C514 VTAIL.n374 B 0.02556f
C515 VTAIL.n375 B 0.01145f
C516 VTAIL.n376 B 0.010814f
C517 VTAIL.n377 B 0.020124f
C518 VTAIL.n378 B 0.020124f
C519 VTAIL.n379 B 0.010814f
C520 VTAIL.n380 B 0.01145f
C521 VTAIL.n381 B 0.02556f
C522 VTAIL.n382 B 0.02556f
C523 VTAIL.n383 B 0.01145f
C524 VTAIL.n384 B 0.010814f
C525 VTAIL.n385 B 0.020124f
C526 VTAIL.n386 B 0.020124f
C527 VTAIL.n387 B 0.010814f
C528 VTAIL.n388 B 0.01145f
C529 VTAIL.n389 B 0.02556f
C530 VTAIL.n390 B 0.057974f
C531 VTAIL.n391 B 0.01145f
C532 VTAIL.n392 B 0.010814f
C533 VTAIL.n393 B 0.046241f
C534 VTAIL.n394 B 0.032702f
C535 VTAIL.n395 B 0.288986f
C536 VTAIL.n396 B 0.02978f
C537 VTAIL.n397 B 0.020124f
C538 VTAIL.n398 B 0.010814f
C539 VTAIL.n399 B 0.02556f
C540 VTAIL.n400 B 0.01145f
C541 VTAIL.n401 B 0.020124f
C542 VTAIL.n402 B 0.010814f
C543 VTAIL.n403 B 0.02556f
C544 VTAIL.n404 B 0.01145f
C545 VTAIL.n405 B 0.020124f
C546 VTAIL.n406 B 0.010814f
C547 VTAIL.n407 B 0.02556f
C548 VTAIL.n408 B 0.01145f
C549 VTAIL.n409 B 0.020124f
C550 VTAIL.n410 B 0.011132f
C551 VTAIL.n411 B 0.02556f
C552 VTAIL.n412 B 0.010814f
C553 VTAIL.n413 B 0.01145f
C554 VTAIL.n414 B 0.020124f
C555 VTAIL.n415 B 0.010814f
C556 VTAIL.n416 B 0.02556f
C557 VTAIL.n417 B 0.01145f
C558 VTAIL.n418 B 0.020124f
C559 VTAIL.n419 B 0.010814f
C560 VTAIL.n420 B 0.01917f
C561 VTAIL.n421 B 0.018069f
C562 VTAIL.t12 B 0.043415f
C563 VTAIL.n422 B 0.162629f
C564 VTAIL.n423 B 1.21841f
C565 VTAIL.n424 B 0.010814f
C566 VTAIL.n425 B 0.01145f
C567 VTAIL.n426 B 0.02556f
C568 VTAIL.n427 B 0.02556f
C569 VTAIL.n428 B 0.01145f
C570 VTAIL.n429 B 0.010814f
C571 VTAIL.n430 B 0.020124f
C572 VTAIL.n431 B 0.020124f
C573 VTAIL.n432 B 0.010814f
C574 VTAIL.n433 B 0.01145f
C575 VTAIL.n434 B 0.02556f
C576 VTAIL.n435 B 0.02556f
C577 VTAIL.n436 B 0.01145f
C578 VTAIL.n437 B 0.010814f
C579 VTAIL.n438 B 0.020124f
C580 VTAIL.n439 B 0.020124f
C581 VTAIL.n440 B 0.010814f
C582 VTAIL.n441 B 0.01145f
C583 VTAIL.n442 B 0.02556f
C584 VTAIL.n443 B 0.02556f
C585 VTAIL.n444 B 0.02556f
C586 VTAIL.n445 B 0.011132f
C587 VTAIL.n446 B 0.010814f
C588 VTAIL.n447 B 0.020124f
C589 VTAIL.n448 B 0.020124f
C590 VTAIL.n449 B 0.010814f
C591 VTAIL.n450 B 0.01145f
C592 VTAIL.n451 B 0.02556f
C593 VTAIL.n452 B 0.02556f
C594 VTAIL.n453 B 0.01145f
C595 VTAIL.n454 B 0.010814f
C596 VTAIL.n455 B 0.020124f
C597 VTAIL.n456 B 0.020124f
C598 VTAIL.n457 B 0.010814f
C599 VTAIL.n458 B 0.01145f
C600 VTAIL.n459 B 0.02556f
C601 VTAIL.n460 B 0.02556f
C602 VTAIL.n461 B 0.01145f
C603 VTAIL.n462 B 0.010814f
C604 VTAIL.n463 B 0.020124f
C605 VTAIL.n464 B 0.020124f
C606 VTAIL.n465 B 0.010814f
C607 VTAIL.n466 B 0.01145f
C608 VTAIL.n467 B 0.02556f
C609 VTAIL.n468 B 0.057974f
C610 VTAIL.n469 B 0.01145f
C611 VTAIL.n470 B 0.010814f
C612 VTAIL.n471 B 0.046241f
C613 VTAIL.n472 B 0.032702f
C614 VTAIL.n473 B 0.288986f
C615 VTAIL.t14 B 0.22693f
C616 VTAIL.t8 B 0.22693f
C617 VTAIL.n474 B 1.97936f
C618 VTAIL.n475 B 0.686741f
C619 VTAIL.n476 B 0.02978f
C620 VTAIL.n477 B 0.020124f
C621 VTAIL.n478 B 0.010814f
C622 VTAIL.n479 B 0.02556f
C623 VTAIL.n480 B 0.01145f
C624 VTAIL.n481 B 0.020124f
C625 VTAIL.n482 B 0.010814f
C626 VTAIL.n483 B 0.02556f
C627 VTAIL.n484 B 0.01145f
C628 VTAIL.n485 B 0.020124f
C629 VTAIL.n486 B 0.010814f
C630 VTAIL.n487 B 0.02556f
C631 VTAIL.n488 B 0.01145f
C632 VTAIL.n489 B 0.020124f
C633 VTAIL.n490 B 0.011132f
C634 VTAIL.n491 B 0.02556f
C635 VTAIL.n492 B 0.010814f
C636 VTAIL.n493 B 0.01145f
C637 VTAIL.n494 B 0.020124f
C638 VTAIL.n495 B 0.010814f
C639 VTAIL.n496 B 0.02556f
C640 VTAIL.n497 B 0.01145f
C641 VTAIL.n498 B 0.020124f
C642 VTAIL.n499 B 0.010814f
C643 VTAIL.n500 B 0.01917f
C644 VTAIL.n501 B 0.018069f
C645 VTAIL.t9 B 0.043415f
C646 VTAIL.n502 B 0.162629f
C647 VTAIL.n503 B 1.21841f
C648 VTAIL.n504 B 0.010814f
C649 VTAIL.n505 B 0.01145f
C650 VTAIL.n506 B 0.02556f
C651 VTAIL.n507 B 0.02556f
C652 VTAIL.n508 B 0.01145f
C653 VTAIL.n509 B 0.010814f
C654 VTAIL.n510 B 0.020124f
C655 VTAIL.n511 B 0.020124f
C656 VTAIL.n512 B 0.010814f
C657 VTAIL.n513 B 0.01145f
C658 VTAIL.n514 B 0.02556f
C659 VTAIL.n515 B 0.02556f
C660 VTAIL.n516 B 0.01145f
C661 VTAIL.n517 B 0.010814f
C662 VTAIL.n518 B 0.020124f
C663 VTAIL.n519 B 0.020124f
C664 VTAIL.n520 B 0.010814f
C665 VTAIL.n521 B 0.01145f
C666 VTAIL.n522 B 0.02556f
C667 VTAIL.n523 B 0.02556f
C668 VTAIL.n524 B 0.02556f
C669 VTAIL.n525 B 0.011132f
C670 VTAIL.n526 B 0.010814f
C671 VTAIL.n527 B 0.020124f
C672 VTAIL.n528 B 0.020124f
C673 VTAIL.n529 B 0.010814f
C674 VTAIL.n530 B 0.01145f
C675 VTAIL.n531 B 0.02556f
C676 VTAIL.n532 B 0.02556f
C677 VTAIL.n533 B 0.01145f
C678 VTAIL.n534 B 0.010814f
C679 VTAIL.n535 B 0.020124f
C680 VTAIL.n536 B 0.020124f
C681 VTAIL.n537 B 0.010814f
C682 VTAIL.n538 B 0.01145f
C683 VTAIL.n539 B 0.02556f
C684 VTAIL.n540 B 0.02556f
C685 VTAIL.n541 B 0.01145f
C686 VTAIL.n542 B 0.010814f
C687 VTAIL.n543 B 0.020124f
C688 VTAIL.n544 B 0.020124f
C689 VTAIL.n545 B 0.010814f
C690 VTAIL.n546 B 0.01145f
C691 VTAIL.n547 B 0.02556f
C692 VTAIL.n548 B 0.057974f
C693 VTAIL.n549 B 0.01145f
C694 VTAIL.n550 B 0.010814f
C695 VTAIL.n551 B 0.046241f
C696 VTAIL.n552 B 0.032702f
C697 VTAIL.n553 B 1.57106f
C698 VTAIL.n554 B 0.02978f
C699 VTAIL.n555 B 0.020124f
C700 VTAIL.n556 B 0.010814f
C701 VTAIL.n557 B 0.02556f
C702 VTAIL.n558 B 0.01145f
C703 VTAIL.n559 B 0.020124f
C704 VTAIL.n560 B 0.010814f
C705 VTAIL.n561 B 0.02556f
C706 VTAIL.n562 B 0.01145f
C707 VTAIL.n563 B 0.020124f
C708 VTAIL.n564 B 0.010814f
C709 VTAIL.n565 B 0.02556f
C710 VTAIL.n566 B 0.01145f
C711 VTAIL.n567 B 0.020124f
C712 VTAIL.n568 B 0.011132f
C713 VTAIL.n569 B 0.02556f
C714 VTAIL.n570 B 0.01145f
C715 VTAIL.n571 B 0.020124f
C716 VTAIL.n572 B 0.010814f
C717 VTAIL.n573 B 0.02556f
C718 VTAIL.n574 B 0.01145f
C719 VTAIL.n575 B 0.020124f
C720 VTAIL.n576 B 0.010814f
C721 VTAIL.n577 B 0.01917f
C722 VTAIL.n578 B 0.018069f
C723 VTAIL.t2 B 0.043415f
C724 VTAIL.n579 B 0.162629f
C725 VTAIL.n580 B 1.21841f
C726 VTAIL.n581 B 0.010814f
C727 VTAIL.n582 B 0.01145f
C728 VTAIL.n583 B 0.02556f
C729 VTAIL.n584 B 0.02556f
C730 VTAIL.n585 B 0.01145f
C731 VTAIL.n586 B 0.010814f
C732 VTAIL.n587 B 0.020124f
C733 VTAIL.n588 B 0.020124f
C734 VTAIL.n589 B 0.010814f
C735 VTAIL.n590 B 0.01145f
C736 VTAIL.n591 B 0.02556f
C737 VTAIL.n592 B 0.02556f
C738 VTAIL.n593 B 0.01145f
C739 VTAIL.n594 B 0.010814f
C740 VTAIL.n595 B 0.020124f
C741 VTAIL.n596 B 0.020124f
C742 VTAIL.n597 B 0.010814f
C743 VTAIL.n598 B 0.010814f
C744 VTAIL.n599 B 0.01145f
C745 VTAIL.n600 B 0.02556f
C746 VTAIL.n601 B 0.02556f
C747 VTAIL.n602 B 0.02556f
C748 VTAIL.n603 B 0.011132f
C749 VTAIL.n604 B 0.010814f
C750 VTAIL.n605 B 0.020124f
C751 VTAIL.n606 B 0.020124f
C752 VTAIL.n607 B 0.010814f
C753 VTAIL.n608 B 0.01145f
C754 VTAIL.n609 B 0.02556f
C755 VTAIL.n610 B 0.02556f
C756 VTAIL.n611 B 0.01145f
C757 VTAIL.n612 B 0.010814f
C758 VTAIL.n613 B 0.020124f
C759 VTAIL.n614 B 0.020124f
C760 VTAIL.n615 B 0.010814f
C761 VTAIL.n616 B 0.01145f
C762 VTAIL.n617 B 0.02556f
C763 VTAIL.n618 B 0.02556f
C764 VTAIL.n619 B 0.01145f
C765 VTAIL.n620 B 0.010814f
C766 VTAIL.n621 B 0.020124f
C767 VTAIL.n622 B 0.020124f
C768 VTAIL.n623 B 0.010814f
C769 VTAIL.n624 B 0.01145f
C770 VTAIL.n625 B 0.02556f
C771 VTAIL.n626 B 0.057974f
C772 VTAIL.n627 B 0.01145f
C773 VTAIL.n628 B 0.010814f
C774 VTAIL.n629 B 0.046241f
C775 VTAIL.n630 B 0.032702f
C776 VTAIL.n631 B 1.56729f
C777 VP.n0 B 0.031191f
C778 VP.t4 B 2.58415f
C779 VP.n1 B 0.030905f
C780 VP.n2 B 0.016582f
C781 VP.n3 B 0.030905f
C782 VP.n4 B 0.016582f
C783 VP.t2 B 2.58415f
C784 VP.n5 B 0.030905f
C785 VP.n6 B 0.016582f
C786 VP.n7 B 0.030905f
C787 VP.n8 B 0.016582f
C788 VP.t5 B 2.58415f
C789 VP.n9 B 0.030905f
C790 VP.n10 B 0.016582f
C791 VP.n11 B 0.030905f
C792 VP.n12 B 0.031191f
C793 VP.t3 B 2.58415f
C794 VP.n13 B 0.031191f
C795 VP.t0 B 2.58415f
C796 VP.n14 B 0.030905f
C797 VP.n15 B 0.016582f
C798 VP.n16 B 0.030905f
C799 VP.n17 B 0.016582f
C800 VP.t1 B 2.58415f
C801 VP.n18 B 0.030905f
C802 VP.n19 B 0.016582f
C803 VP.n20 B 0.030905f
C804 VP.n21 B 0.219129f
C805 VP.t6 B 2.58415f
C806 VP.t7 B 2.86366f
C807 VP.n22 B 0.911782f
C808 VP.n23 B 0.955302f
C809 VP.n24 B 0.02053f
C810 VP.n25 B 0.030905f
C811 VP.n26 B 0.016582f
C812 VP.n27 B 0.016582f
C813 VP.n28 B 0.016582f
C814 VP.n29 B 0.032957f
C815 VP.n30 B 0.013405f
C816 VP.n31 B 0.032957f
C817 VP.n32 B 0.016582f
C818 VP.n33 B 0.016582f
C819 VP.n34 B 0.016582f
C820 VP.n35 B 0.030905f
C821 VP.n36 B 0.02053f
C822 VP.n37 B 0.897245f
C823 VP.n38 B 0.026023f
C824 VP.n39 B 0.016582f
C825 VP.n40 B 0.016582f
C826 VP.n41 B 0.016582f
C827 VP.n42 B 0.030905f
C828 VP.n43 B 0.027442f
C829 VP.n44 B 0.020973f
C830 VP.n45 B 0.016582f
C831 VP.n46 B 0.016582f
C832 VP.n47 B 0.016582f
C833 VP.n48 B 0.030905f
C834 VP.n49 B 0.030295f
C835 VP.n50 B 0.974237f
C836 VP.n51 B 1.21889f
C837 VP.n52 B 1.22892f
C838 VP.n53 B 0.974237f
C839 VP.n54 B 0.030295f
C840 VP.n55 B 0.030905f
C841 VP.n56 B 0.016582f
C842 VP.n57 B 0.016582f
C843 VP.n58 B 0.016582f
C844 VP.n59 B 0.020973f
C845 VP.n60 B 0.027442f
C846 VP.n61 B 0.030905f
C847 VP.n62 B 0.016582f
C848 VP.n63 B 0.016582f
C849 VP.n64 B 0.016582f
C850 VP.n65 B 0.026023f
C851 VP.n66 B 0.897245f
C852 VP.n67 B 0.02053f
C853 VP.n68 B 0.030905f
C854 VP.n69 B 0.016582f
C855 VP.n70 B 0.016582f
C856 VP.n71 B 0.016582f
C857 VP.n72 B 0.032957f
C858 VP.n73 B 0.013405f
C859 VP.n74 B 0.032957f
C860 VP.n75 B 0.016582f
C861 VP.n76 B 0.016582f
C862 VP.n77 B 0.016582f
C863 VP.n78 B 0.030905f
C864 VP.n79 B 0.02053f
C865 VP.n80 B 0.897245f
C866 VP.n81 B 0.026023f
C867 VP.n82 B 0.016582f
C868 VP.n83 B 0.016582f
C869 VP.n84 B 0.016582f
C870 VP.n85 B 0.030905f
C871 VP.n86 B 0.027442f
C872 VP.n87 B 0.020973f
C873 VP.n88 B 0.016582f
C874 VP.n89 B 0.016582f
C875 VP.n90 B 0.016582f
C876 VP.n91 B 0.030905f
C877 VP.n92 B 0.030295f
C878 VP.n93 B 0.974237f
C879 VP.n94 B 0.049821f
.ends

