* NGSPICE file created from diff_pair_sample_0184.ext - technology: sky130A

.subckt diff_pair_sample_0184 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VP.t0 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0.3465 ps=2.43 w=2.1 l=0.94
X1 VDD1.t1 VP.t1 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3465 pd=2.43 as=0.819 ps=4.98 w=2.1 l=0.94
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0 ps=0 w=2.1 l=0.94
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0 ps=0 w=2.1 l=0.94
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0 ps=0 w=2.1 l=0.94
X5 VTAIL.t2 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0.3465 ps=2.43 w=2.1 l=0.94
X6 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0.3465 ps=2.43 w=2.1 l=0.94
X7 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3465 pd=2.43 as=0.819 ps=4.98 w=2.1 l=0.94
X8 VDD1.t0 VP.t2 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3465 pd=2.43 as=0.819 ps=4.98 w=2.1 l=0.94
X9 VDD2.t0 VN.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3465 pd=2.43 as=0.819 ps=4.98 w=2.1 l=0.94
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0 ps=0 w=2.1 l=0.94
X11 VTAIL.t3 VP.t3 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.819 pd=4.98 as=0.3465 ps=2.43 w=2.1 l=0.94
R0 VP.n0 VP.t3 114.751
R1 VP.n0 VP.t2 114.663
R2 VP.n2 VP.t0 96.1441
R3 VP.n3 VP.t1 96.1441
R4 VP.n4 VP.n3 80.6037
R5 VP.n2 VP.n1 80.6037
R6 VP.n1 VP.n0 64.935
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.380177
R9 VP VP.n4 0.146778
R10 VDD1 VDD1.n1 121.251
R11 VDD1 VDD1.n0 91.9743
R12 VDD1.n0 VDD1.t3 9.42907
R13 VDD1.n0 VDD1.t0 9.42907
R14 VDD1.n1 VDD1.t2 9.42907
R15 VDD1.n1 VDD1.t1 9.42907
R16 VTAIL.n7 VTAIL.t0 84.6659
R17 VTAIL.n0 VTAIL.t2 84.6659
R18 VTAIL.n1 VTAIL.t5 84.6659
R19 VTAIL.n2 VTAIL.t6 84.6659
R20 VTAIL.n6 VTAIL.t4 84.6659
R21 VTAIL.n5 VTAIL.t3 84.6658
R22 VTAIL.n4 VTAIL.t7 84.6658
R23 VTAIL.n3 VTAIL.t1 84.6658
R24 VTAIL.n7 VTAIL.n6 15.2721
R25 VTAIL.n3 VTAIL.n2 15.2721
R26 VTAIL.n4 VTAIL.n3 1.09533
R27 VTAIL.n6 VTAIL.n5 1.09533
R28 VTAIL.n2 VTAIL.n1 1.09533
R29 VTAIL VTAIL.n0 0.606103
R30 VTAIL VTAIL.n7 0.489724
R31 VTAIL.n5 VTAIL.n4 0.470328
R32 VTAIL.n1 VTAIL.n0 0.470328
R33 B.n341 B.n340 585
R34 B.n342 B.n341 585
R35 B.n127 B.n57 585
R36 B.n126 B.n125 585
R37 B.n124 B.n123 585
R38 B.n122 B.n121 585
R39 B.n120 B.n119 585
R40 B.n118 B.n117 585
R41 B.n116 B.n115 585
R42 B.n114 B.n113 585
R43 B.n112 B.n111 585
R44 B.n110 B.n109 585
R45 B.n108 B.n107 585
R46 B.n106 B.n105 585
R47 B.n104 B.n103 585
R48 B.n102 B.n101 585
R49 B.n100 B.n99 585
R50 B.n98 B.n97 585
R51 B.n96 B.n95 585
R52 B.n94 B.n93 585
R53 B.n92 B.n91 585
R54 B.n90 B.n89 585
R55 B.n88 B.n87 585
R56 B.n85 B.n84 585
R57 B.n83 B.n82 585
R58 B.n81 B.n80 585
R59 B.n79 B.n78 585
R60 B.n77 B.n76 585
R61 B.n75 B.n74 585
R62 B.n73 B.n72 585
R63 B.n71 B.n70 585
R64 B.n69 B.n68 585
R65 B.n67 B.n66 585
R66 B.n65 B.n64 585
R67 B.n40 B.n39 585
R68 B.n345 B.n344 585
R69 B.n339 B.n58 585
R70 B.n58 B.n37 585
R71 B.n338 B.n36 585
R72 B.n349 B.n36 585
R73 B.n337 B.n35 585
R74 B.n350 B.n35 585
R75 B.n336 B.n34 585
R76 B.n351 B.n34 585
R77 B.n335 B.n334 585
R78 B.n334 B.n30 585
R79 B.n333 B.n29 585
R80 B.n357 B.n29 585
R81 B.n332 B.n28 585
R82 B.n358 B.n28 585
R83 B.n331 B.n27 585
R84 B.n359 B.n27 585
R85 B.n330 B.n329 585
R86 B.n329 B.n23 585
R87 B.n328 B.n22 585
R88 B.n365 B.n22 585
R89 B.n327 B.n21 585
R90 B.n366 B.n21 585
R91 B.n326 B.n20 585
R92 B.n367 B.n20 585
R93 B.n325 B.n324 585
R94 B.n324 B.n19 585
R95 B.n323 B.n15 585
R96 B.n373 B.n15 585
R97 B.n322 B.n14 585
R98 B.n374 B.n14 585
R99 B.n321 B.n13 585
R100 B.n375 B.n13 585
R101 B.n320 B.n319 585
R102 B.n319 B.n12 585
R103 B.n318 B.n317 585
R104 B.n318 B.n8 585
R105 B.n316 B.n7 585
R106 B.n382 B.n7 585
R107 B.n315 B.n6 585
R108 B.n383 B.n6 585
R109 B.n314 B.n5 585
R110 B.n384 B.n5 585
R111 B.n313 B.n312 585
R112 B.n312 B.n4 585
R113 B.n311 B.n128 585
R114 B.n311 B.n310 585
R115 B.n300 B.n129 585
R116 B.n303 B.n129 585
R117 B.n302 B.n301 585
R118 B.n304 B.n302 585
R119 B.n299 B.n134 585
R120 B.n134 B.n133 585
R121 B.n298 B.n297 585
R122 B.n297 B.n296 585
R123 B.n136 B.n135 585
R124 B.n289 B.n136 585
R125 B.n288 B.n287 585
R126 B.n290 B.n288 585
R127 B.n286 B.n141 585
R128 B.n141 B.n140 585
R129 B.n285 B.n284 585
R130 B.n284 B.n283 585
R131 B.n143 B.n142 585
R132 B.n144 B.n143 585
R133 B.n276 B.n275 585
R134 B.n277 B.n276 585
R135 B.n274 B.n149 585
R136 B.n149 B.n148 585
R137 B.n273 B.n272 585
R138 B.n272 B.n271 585
R139 B.n151 B.n150 585
R140 B.n152 B.n151 585
R141 B.n264 B.n263 585
R142 B.n265 B.n264 585
R143 B.n262 B.n157 585
R144 B.n157 B.n156 585
R145 B.n261 B.n260 585
R146 B.n260 B.n259 585
R147 B.n159 B.n158 585
R148 B.n160 B.n159 585
R149 B.n255 B.n254 585
R150 B.n163 B.n162 585
R151 B.n251 B.n250 585
R152 B.n252 B.n251 585
R153 B.n249 B.n180 585
R154 B.n248 B.n247 585
R155 B.n246 B.n245 585
R156 B.n244 B.n243 585
R157 B.n242 B.n241 585
R158 B.n240 B.n239 585
R159 B.n238 B.n237 585
R160 B.n236 B.n235 585
R161 B.n234 B.n233 585
R162 B.n232 B.n231 585
R163 B.n230 B.n229 585
R164 B.n228 B.n227 585
R165 B.n226 B.n225 585
R166 B.n224 B.n223 585
R167 B.n222 B.n221 585
R168 B.n220 B.n219 585
R169 B.n218 B.n217 585
R170 B.n216 B.n215 585
R171 B.n214 B.n213 585
R172 B.n211 B.n210 585
R173 B.n209 B.n208 585
R174 B.n207 B.n206 585
R175 B.n205 B.n204 585
R176 B.n203 B.n202 585
R177 B.n201 B.n200 585
R178 B.n199 B.n198 585
R179 B.n197 B.n196 585
R180 B.n195 B.n194 585
R181 B.n193 B.n192 585
R182 B.n191 B.n190 585
R183 B.n189 B.n188 585
R184 B.n187 B.n186 585
R185 B.n256 B.n161 585
R186 B.n161 B.n160 585
R187 B.n258 B.n257 585
R188 B.n259 B.n258 585
R189 B.n155 B.n154 585
R190 B.n156 B.n155 585
R191 B.n267 B.n266 585
R192 B.n266 B.n265 585
R193 B.n268 B.n153 585
R194 B.n153 B.n152 585
R195 B.n270 B.n269 585
R196 B.n271 B.n270 585
R197 B.n147 B.n146 585
R198 B.n148 B.n147 585
R199 B.n279 B.n278 585
R200 B.n278 B.n277 585
R201 B.n280 B.n145 585
R202 B.n145 B.n144 585
R203 B.n282 B.n281 585
R204 B.n283 B.n282 585
R205 B.n139 B.n138 585
R206 B.n140 B.n139 585
R207 B.n292 B.n291 585
R208 B.n291 B.n290 585
R209 B.n293 B.n137 585
R210 B.n289 B.n137 585
R211 B.n295 B.n294 585
R212 B.n296 B.n295 585
R213 B.n132 B.n131 585
R214 B.n133 B.n132 585
R215 B.n306 B.n305 585
R216 B.n305 B.n304 585
R217 B.n307 B.n130 585
R218 B.n303 B.n130 585
R219 B.n309 B.n308 585
R220 B.n310 B.n309 585
R221 B.n3 B.n0 585
R222 B.n4 B.n3 585
R223 B.n381 B.n1 585
R224 B.n382 B.n381 585
R225 B.n380 B.n379 585
R226 B.n380 B.n8 585
R227 B.n378 B.n9 585
R228 B.n12 B.n9 585
R229 B.n377 B.n376 585
R230 B.n376 B.n375 585
R231 B.n11 B.n10 585
R232 B.n374 B.n11 585
R233 B.n372 B.n371 585
R234 B.n373 B.n372 585
R235 B.n370 B.n16 585
R236 B.n19 B.n16 585
R237 B.n369 B.n368 585
R238 B.n368 B.n367 585
R239 B.n18 B.n17 585
R240 B.n366 B.n18 585
R241 B.n364 B.n363 585
R242 B.n365 B.n364 585
R243 B.n362 B.n24 585
R244 B.n24 B.n23 585
R245 B.n361 B.n360 585
R246 B.n360 B.n359 585
R247 B.n26 B.n25 585
R248 B.n358 B.n26 585
R249 B.n356 B.n355 585
R250 B.n357 B.n356 585
R251 B.n354 B.n31 585
R252 B.n31 B.n30 585
R253 B.n353 B.n352 585
R254 B.n352 B.n351 585
R255 B.n33 B.n32 585
R256 B.n350 B.n33 585
R257 B.n348 B.n347 585
R258 B.n349 B.n348 585
R259 B.n346 B.n38 585
R260 B.n38 B.n37 585
R261 B.n385 B.n384 585
R262 B.n383 B.n2 585
R263 B.n344 B.n38 434.841
R264 B.n341 B.n58 434.841
R265 B.n186 B.n159 434.841
R266 B.n254 B.n161 434.841
R267 B.n342 B.n56 256.663
R268 B.n342 B.n55 256.663
R269 B.n342 B.n54 256.663
R270 B.n342 B.n53 256.663
R271 B.n342 B.n52 256.663
R272 B.n342 B.n51 256.663
R273 B.n342 B.n50 256.663
R274 B.n342 B.n49 256.663
R275 B.n342 B.n48 256.663
R276 B.n342 B.n47 256.663
R277 B.n342 B.n46 256.663
R278 B.n342 B.n45 256.663
R279 B.n342 B.n44 256.663
R280 B.n342 B.n43 256.663
R281 B.n342 B.n42 256.663
R282 B.n342 B.n41 256.663
R283 B.n343 B.n342 256.663
R284 B.n253 B.n252 256.663
R285 B.n252 B.n164 256.663
R286 B.n252 B.n165 256.663
R287 B.n252 B.n166 256.663
R288 B.n252 B.n167 256.663
R289 B.n252 B.n168 256.663
R290 B.n252 B.n169 256.663
R291 B.n252 B.n170 256.663
R292 B.n252 B.n171 256.663
R293 B.n252 B.n172 256.663
R294 B.n252 B.n173 256.663
R295 B.n252 B.n174 256.663
R296 B.n252 B.n175 256.663
R297 B.n252 B.n176 256.663
R298 B.n252 B.n177 256.663
R299 B.n252 B.n178 256.663
R300 B.n252 B.n179 256.663
R301 B.n387 B.n386 256.663
R302 B.n62 B.t12 256.341
R303 B.n59 B.t4 256.341
R304 B.n184 B.t8 256.341
R305 B.n181 B.t15 256.341
R306 B.n252 B.n160 165.56
R307 B.n342 B.n37 165.56
R308 B.n64 B.n40 163.367
R309 B.n68 B.n67 163.367
R310 B.n72 B.n71 163.367
R311 B.n76 B.n75 163.367
R312 B.n80 B.n79 163.367
R313 B.n84 B.n83 163.367
R314 B.n89 B.n88 163.367
R315 B.n93 B.n92 163.367
R316 B.n97 B.n96 163.367
R317 B.n101 B.n100 163.367
R318 B.n105 B.n104 163.367
R319 B.n109 B.n108 163.367
R320 B.n113 B.n112 163.367
R321 B.n117 B.n116 163.367
R322 B.n121 B.n120 163.367
R323 B.n125 B.n124 163.367
R324 B.n341 B.n57 163.367
R325 B.n260 B.n159 163.367
R326 B.n260 B.n157 163.367
R327 B.n264 B.n157 163.367
R328 B.n264 B.n151 163.367
R329 B.n272 B.n151 163.367
R330 B.n272 B.n149 163.367
R331 B.n276 B.n149 163.367
R332 B.n276 B.n143 163.367
R333 B.n284 B.n143 163.367
R334 B.n284 B.n141 163.367
R335 B.n288 B.n141 163.367
R336 B.n288 B.n136 163.367
R337 B.n297 B.n136 163.367
R338 B.n297 B.n134 163.367
R339 B.n302 B.n134 163.367
R340 B.n302 B.n129 163.367
R341 B.n311 B.n129 163.367
R342 B.n312 B.n311 163.367
R343 B.n312 B.n5 163.367
R344 B.n6 B.n5 163.367
R345 B.n7 B.n6 163.367
R346 B.n318 B.n7 163.367
R347 B.n319 B.n318 163.367
R348 B.n319 B.n13 163.367
R349 B.n14 B.n13 163.367
R350 B.n15 B.n14 163.367
R351 B.n324 B.n15 163.367
R352 B.n324 B.n20 163.367
R353 B.n21 B.n20 163.367
R354 B.n22 B.n21 163.367
R355 B.n329 B.n22 163.367
R356 B.n329 B.n27 163.367
R357 B.n28 B.n27 163.367
R358 B.n29 B.n28 163.367
R359 B.n334 B.n29 163.367
R360 B.n334 B.n34 163.367
R361 B.n35 B.n34 163.367
R362 B.n36 B.n35 163.367
R363 B.n58 B.n36 163.367
R364 B.n251 B.n163 163.367
R365 B.n251 B.n180 163.367
R366 B.n247 B.n246 163.367
R367 B.n243 B.n242 163.367
R368 B.n239 B.n238 163.367
R369 B.n235 B.n234 163.367
R370 B.n231 B.n230 163.367
R371 B.n227 B.n226 163.367
R372 B.n223 B.n222 163.367
R373 B.n219 B.n218 163.367
R374 B.n215 B.n214 163.367
R375 B.n210 B.n209 163.367
R376 B.n206 B.n205 163.367
R377 B.n202 B.n201 163.367
R378 B.n198 B.n197 163.367
R379 B.n194 B.n193 163.367
R380 B.n190 B.n189 163.367
R381 B.n258 B.n161 163.367
R382 B.n258 B.n155 163.367
R383 B.n266 B.n155 163.367
R384 B.n266 B.n153 163.367
R385 B.n270 B.n153 163.367
R386 B.n270 B.n147 163.367
R387 B.n278 B.n147 163.367
R388 B.n278 B.n145 163.367
R389 B.n282 B.n145 163.367
R390 B.n282 B.n139 163.367
R391 B.n291 B.n139 163.367
R392 B.n291 B.n137 163.367
R393 B.n295 B.n137 163.367
R394 B.n295 B.n132 163.367
R395 B.n305 B.n132 163.367
R396 B.n305 B.n130 163.367
R397 B.n309 B.n130 163.367
R398 B.n309 B.n3 163.367
R399 B.n385 B.n3 163.367
R400 B.n381 B.n2 163.367
R401 B.n381 B.n380 163.367
R402 B.n380 B.n9 163.367
R403 B.n376 B.n9 163.367
R404 B.n376 B.n11 163.367
R405 B.n372 B.n11 163.367
R406 B.n372 B.n16 163.367
R407 B.n368 B.n16 163.367
R408 B.n368 B.n18 163.367
R409 B.n364 B.n18 163.367
R410 B.n364 B.n24 163.367
R411 B.n360 B.n24 163.367
R412 B.n360 B.n26 163.367
R413 B.n356 B.n26 163.367
R414 B.n356 B.n31 163.367
R415 B.n352 B.n31 163.367
R416 B.n352 B.n33 163.367
R417 B.n348 B.n33 163.367
R418 B.n348 B.n38 163.367
R419 B.n59 B.t6 108.828
R420 B.n184 B.t11 108.828
R421 B.n62 B.t13 108.826
R422 B.n181 B.t17 108.826
R423 B.n259 B.n160 101.424
R424 B.n259 B.n156 101.424
R425 B.n265 B.n156 101.424
R426 B.n265 B.n152 101.424
R427 B.n271 B.n152 101.424
R428 B.n277 B.n148 101.424
R429 B.n277 B.n144 101.424
R430 B.n283 B.n144 101.424
R431 B.n283 B.n140 101.424
R432 B.n290 B.n140 101.424
R433 B.n290 B.n289 101.424
R434 B.n296 B.n133 101.424
R435 B.n304 B.n133 101.424
R436 B.n304 B.n303 101.424
R437 B.n310 B.n4 101.424
R438 B.n384 B.n4 101.424
R439 B.n384 B.n383 101.424
R440 B.n383 B.n382 101.424
R441 B.n382 B.n8 101.424
R442 B.n375 B.n12 101.424
R443 B.n375 B.n374 101.424
R444 B.n374 B.n373 101.424
R445 B.n367 B.n19 101.424
R446 B.n367 B.n366 101.424
R447 B.n366 B.n365 101.424
R448 B.n365 B.n23 101.424
R449 B.n359 B.n23 101.424
R450 B.n359 B.n358 101.424
R451 B.n357 B.n30 101.424
R452 B.n351 B.n30 101.424
R453 B.n351 B.n350 101.424
R454 B.n350 B.n349 101.424
R455 B.n349 B.n37 101.424
R456 B.n310 B.t3 98.4412
R457 B.t2 B.n8 98.4412
R458 B.n60 B.t7 84.1969
R459 B.n185 B.t10 84.1969
R460 B.n63 B.t14 84.1967
R461 B.n182 B.t16 84.1967
R462 B.n344 B.n343 71.676
R463 B.n64 B.n41 71.676
R464 B.n68 B.n42 71.676
R465 B.n72 B.n43 71.676
R466 B.n76 B.n44 71.676
R467 B.n80 B.n45 71.676
R468 B.n84 B.n46 71.676
R469 B.n89 B.n47 71.676
R470 B.n93 B.n48 71.676
R471 B.n97 B.n49 71.676
R472 B.n101 B.n50 71.676
R473 B.n105 B.n51 71.676
R474 B.n109 B.n52 71.676
R475 B.n113 B.n53 71.676
R476 B.n117 B.n54 71.676
R477 B.n121 B.n55 71.676
R478 B.n125 B.n56 71.676
R479 B.n57 B.n56 71.676
R480 B.n124 B.n55 71.676
R481 B.n120 B.n54 71.676
R482 B.n116 B.n53 71.676
R483 B.n112 B.n52 71.676
R484 B.n108 B.n51 71.676
R485 B.n104 B.n50 71.676
R486 B.n100 B.n49 71.676
R487 B.n96 B.n48 71.676
R488 B.n92 B.n47 71.676
R489 B.n88 B.n46 71.676
R490 B.n83 B.n45 71.676
R491 B.n79 B.n44 71.676
R492 B.n75 B.n43 71.676
R493 B.n71 B.n42 71.676
R494 B.n67 B.n41 71.676
R495 B.n343 B.n40 71.676
R496 B.n254 B.n253 71.676
R497 B.n180 B.n164 71.676
R498 B.n246 B.n165 71.676
R499 B.n242 B.n166 71.676
R500 B.n238 B.n167 71.676
R501 B.n234 B.n168 71.676
R502 B.n230 B.n169 71.676
R503 B.n226 B.n170 71.676
R504 B.n222 B.n171 71.676
R505 B.n218 B.n172 71.676
R506 B.n214 B.n173 71.676
R507 B.n209 B.n174 71.676
R508 B.n205 B.n175 71.676
R509 B.n201 B.n176 71.676
R510 B.n197 B.n177 71.676
R511 B.n193 B.n178 71.676
R512 B.n189 B.n179 71.676
R513 B.n253 B.n163 71.676
R514 B.n247 B.n164 71.676
R515 B.n243 B.n165 71.676
R516 B.n239 B.n166 71.676
R517 B.n235 B.n167 71.676
R518 B.n231 B.n168 71.676
R519 B.n227 B.n169 71.676
R520 B.n223 B.n170 71.676
R521 B.n219 B.n171 71.676
R522 B.n215 B.n172 71.676
R523 B.n210 B.n173 71.676
R524 B.n206 B.n174 71.676
R525 B.n202 B.n175 71.676
R526 B.n198 B.n176 71.676
R527 B.n194 B.n177 71.676
R528 B.n190 B.n178 71.676
R529 B.n186 B.n179 71.676
R530 B.n386 B.n385 71.676
R531 B.n386 B.n2 71.676
R532 B.n296 B.t1 71.5937
R533 B.n373 B.t0 71.5937
R534 B.t9 B.n148 65.6276
R535 B.n358 B.t5 65.6276
R536 B.n86 B.n63 59.5399
R537 B.n61 B.n60 59.5399
R538 B.n212 B.n185 59.5399
R539 B.n183 B.n182 59.5399
R540 B.n271 B.t9 35.7971
R541 B.t5 B.n357 35.7971
R542 B.n289 B.t1 29.831
R543 B.n19 B.t0 29.831
R544 B.n256 B.n255 28.2542
R545 B.n187 B.n158 28.2542
R546 B.n340 B.n339 28.2542
R547 B.n346 B.n345 28.2542
R548 B.n63 B.n62 24.6308
R549 B.n60 B.n59 24.6308
R550 B.n185 B.n184 24.6308
R551 B.n182 B.n181 24.6308
R552 B B.n387 18.0485
R553 B.n257 B.n256 10.6151
R554 B.n257 B.n154 10.6151
R555 B.n267 B.n154 10.6151
R556 B.n268 B.n267 10.6151
R557 B.n269 B.n268 10.6151
R558 B.n269 B.n146 10.6151
R559 B.n279 B.n146 10.6151
R560 B.n280 B.n279 10.6151
R561 B.n281 B.n280 10.6151
R562 B.n281 B.n138 10.6151
R563 B.n292 B.n138 10.6151
R564 B.n293 B.n292 10.6151
R565 B.n294 B.n293 10.6151
R566 B.n294 B.n131 10.6151
R567 B.n306 B.n131 10.6151
R568 B.n307 B.n306 10.6151
R569 B.n308 B.n307 10.6151
R570 B.n308 B.n0 10.6151
R571 B.n255 B.n162 10.6151
R572 B.n250 B.n162 10.6151
R573 B.n250 B.n249 10.6151
R574 B.n249 B.n248 10.6151
R575 B.n248 B.n245 10.6151
R576 B.n245 B.n244 10.6151
R577 B.n244 B.n241 10.6151
R578 B.n241 B.n240 10.6151
R579 B.n240 B.n237 10.6151
R580 B.n237 B.n236 10.6151
R581 B.n236 B.n233 10.6151
R582 B.n233 B.n232 10.6151
R583 B.n229 B.n228 10.6151
R584 B.n228 B.n225 10.6151
R585 B.n225 B.n224 10.6151
R586 B.n224 B.n221 10.6151
R587 B.n221 B.n220 10.6151
R588 B.n220 B.n217 10.6151
R589 B.n217 B.n216 10.6151
R590 B.n216 B.n213 10.6151
R591 B.n211 B.n208 10.6151
R592 B.n208 B.n207 10.6151
R593 B.n207 B.n204 10.6151
R594 B.n204 B.n203 10.6151
R595 B.n203 B.n200 10.6151
R596 B.n200 B.n199 10.6151
R597 B.n199 B.n196 10.6151
R598 B.n196 B.n195 10.6151
R599 B.n195 B.n192 10.6151
R600 B.n192 B.n191 10.6151
R601 B.n191 B.n188 10.6151
R602 B.n188 B.n187 10.6151
R603 B.n261 B.n158 10.6151
R604 B.n262 B.n261 10.6151
R605 B.n263 B.n262 10.6151
R606 B.n263 B.n150 10.6151
R607 B.n273 B.n150 10.6151
R608 B.n274 B.n273 10.6151
R609 B.n275 B.n274 10.6151
R610 B.n275 B.n142 10.6151
R611 B.n285 B.n142 10.6151
R612 B.n286 B.n285 10.6151
R613 B.n287 B.n286 10.6151
R614 B.n287 B.n135 10.6151
R615 B.n298 B.n135 10.6151
R616 B.n299 B.n298 10.6151
R617 B.n301 B.n299 10.6151
R618 B.n301 B.n300 10.6151
R619 B.n300 B.n128 10.6151
R620 B.n313 B.n128 10.6151
R621 B.n314 B.n313 10.6151
R622 B.n315 B.n314 10.6151
R623 B.n316 B.n315 10.6151
R624 B.n317 B.n316 10.6151
R625 B.n320 B.n317 10.6151
R626 B.n321 B.n320 10.6151
R627 B.n322 B.n321 10.6151
R628 B.n323 B.n322 10.6151
R629 B.n325 B.n323 10.6151
R630 B.n326 B.n325 10.6151
R631 B.n327 B.n326 10.6151
R632 B.n328 B.n327 10.6151
R633 B.n330 B.n328 10.6151
R634 B.n331 B.n330 10.6151
R635 B.n332 B.n331 10.6151
R636 B.n333 B.n332 10.6151
R637 B.n335 B.n333 10.6151
R638 B.n336 B.n335 10.6151
R639 B.n337 B.n336 10.6151
R640 B.n338 B.n337 10.6151
R641 B.n339 B.n338 10.6151
R642 B.n379 B.n1 10.6151
R643 B.n379 B.n378 10.6151
R644 B.n378 B.n377 10.6151
R645 B.n377 B.n10 10.6151
R646 B.n371 B.n10 10.6151
R647 B.n371 B.n370 10.6151
R648 B.n370 B.n369 10.6151
R649 B.n369 B.n17 10.6151
R650 B.n363 B.n17 10.6151
R651 B.n363 B.n362 10.6151
R652 B.n362 B.n361 10.6151
R653 B.n361 B.n25 10.6151
R654 B.n355 B.n25 10.6151
R655 B.n355 B.n354 10.6151
R656 B.n354 B.n353 10.6151
R657 B.n353 B.n32 10.6151
R658 B.n347 B.n32 10.6151
R659 B.n347 B.n346 10.6151
R660 B.n345 B.n39 10.6151
R661 B.n65 B.n39 10.6151
R662 B.n66 B.n65 10.6151
R663 B.n69 B.n66 10.6151
R664 B.n70 B.n69 10.6151
R665 B.n73 B.n70 10.6151
R666 B.n74 B.n73 10.6151
R667 B.n77 B.n74 10.6151
R668 B.n78 B.n77 10.6151
R669 B.n81 B.n78 10.6151
R670 B.n82 B.n81 10.6151
R671 B.n85 B.n82 10.6151
R672 B.n90 B.n87 10.6151
R673 B.n91 B.n90 10.6151
R674 B.n94 B.n91 10.6151
R675 B.n95 B.n94 10.6151
R676 B.n98 B.n95 10.6151
R677 B.n99 B.n98 10.6151
R678 B.n102 B.n99 10.6151
R679 B.n103 B.n102 10.6151
R680 B.n107 B.n106 10.6151
R681 B.n110 B.n107 10.6151
R682 B.n111 B.n110 10.6151
R683 B.n114 B.n111 10.6151
R684 B.n115 B.n114 10.6151
R685 B.n118 B.n115 10.6151
R686 B.n119 B.n118 10.6151
R687 B.n122 B.n119 10.6151
R688 B.n123 B.n122 10.6151
R689 B.n126 B.n123 10.6151
R690 B.n127 B.n126 10.6151
R691 B.n340 B.n127 10.6151
R692 B.n387 B.n0 8.11757
R693 B.n387 B.n1 8.11757
R694 B.n229 B.n183 6.5566
R695 B.n213 B.n212 6.5566
R696 B.n87 B.n86 6.5566
R697 B.n103 B.n61 6.5566
R698 B.n232 B.n183 4.05904
R699 B.n212 B.n211 4.05904
R700 B.n86 B.n85 4.05904
R701 B.n106 B.n61 4.05904
R702 B.n303 B.t3 2.98355
R703 B.n12 B.t2 2.98355
R704 VN.n0 VN.t0 114.751
R705 VN.n1 VN.t3 114.751
R706 VN.n1 VN.t1 114.663
R707 VN.n0 VN.t2 114.663
R708 VN VN.n1 65.2205
R709 VN VN.n0 31.2622
R710 VDD2.n2 VDD2.n0 120.725
R711 VDD2.n2 VDD2.n1 91.9161
R712 VDD2.n1 VDD2.t2 9.42907
R713 VDD2.n1 VDD2.t0 9.42907
R714 VDD2.n0 VDD2.t3 9.42907
R715 VDD2.n0 VDD2.t1 9.42907
R716 VDD2 VDD2.n2 0.0586897
C0 VN VP 3.17405f
C1 VTAIL VDD2 2.44123f
C2 VTAIL VDD1 2.39815f
C3 VDD1 VDD2 0.624597f
C4 VTAIL VP 1.04334f
C5 VTAIL VN 1.02923f
C6 VP VDD2 0.294798f
C7 VP VDD1 1.00768f
C8 VN VDD2 0.866864f
C9 VN VDD1 0.152927f
C10 VDD2 B 2.027741f
C11 VDD1 B 3.82059f
C12 VTAIL B 3.08636f
C13 VN B 6.14986f
C14 VP B 4.593201f
C15 VDD2.t3 B 0.032573f
C16 VDD2.t1 B 0.032573f
C17 VDD2.n0 B 0.379202f
C18 VDD2.t2 B 0.032573f
C19 VDD2.t0 B 0.032573f
C20 VDD2.n1 B 0.220859f
C21 VDD2.n2 B 1.59617f
C22 VN.t0 B 0.206952f
C23 VN.t2 B 0.206822f
C24 VN.n0 B 0.211917f
C25 VN.t3 B 0.206952f
C26 VN.t1 B 0.206822f
C27 VN.n1 B 0.710818f
C28 VTAIL.t2 B 0.206895f
C29 VTAIL.n0 B 0.195161f
C30 VTAIL.t5 B 0.206895f
C31 VTAIL.n1 B 0.220546f
C32 VTAIL.t6 B 0.206895f
C33 VTAIL.n2 B 0.565664f
C34 VTAIL.t1 B 0.206896f
C35 VTAIL.n3 B 0.565663f
C36 VTAIL.t7 B 0.206896f
C37 VTAIL.n4 B 0.220545f
C38 VTAIL.t3 B 0.206896f
C39 VTAIL.n5 B 0.220545f
C40 VTAIL.t4 B 0.206895f
C41 VTAIL.n6 B 0.565664f
C42 VTAIL.t0 B 0.206895f
C43 VTAIL.n7 B 0.53424f
C44 VDD1.t3 B 0.031618f
C45 VDD1.t0 B 0.031618f
C46 VDD1.n0 B 0.214518f
C47 VDD1.t2 B 0.031618f
C48 VDD1.t1 B 0.031618f
C49 VDD1.n1 B 0.379717f
C50 VP.t2 B 0.209636f
C51 VP.t3 B 0.209767f
C52 VP.n0 B 0.709021f
C53 VP.n1 B 1.37222f
C54 VP.t0 B 0.189012f
C55 VP.n2 B 0.127689f
C56 VP.t1 B 0.189012f
C57 VP.n3 B 0.127689f
C58 VP.n4 B 0.039362f
.ends

