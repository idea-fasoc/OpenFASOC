* NGSPICE file created from diff_pair_sample_0234.ext - technology: sky130A

.subckt diff_pair_sample_0234 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.4407 ps=3.04 w=1.13 l=1
X1 VDD1.t4 VP.t1 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.4407 ps=3.04 w=1.13 l=1
X2 VDD2.t5 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.4407 ps=3.04 w=1.13 l=1
X3 VTAIL.t11 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.18645 ps=1.46 w=1.13 l=1
X4 VDD1.t2 VP.t3 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0.18645 ps=1.46 w=1.13 l=1
X5 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0 ps=0 w=1.13 l=1
X6 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0 ps=0 w=1.13 l=1
X7 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.4407 ps=3.04 w=1.13 l=1
X8 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.18645 ps=1.46 w=1.13 l=1
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0 ps=0 w=1.13 l=1
X10 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0.18645 ps=1.46 w=1.13 l=1
X11 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0.18645 ps=1.46 w=1.13 l=1
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0 ps=0 w=1.13 l=1
X13 VTAIL.t4 VN.t5 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.18645 ps=1.46 w=1.13 l=1
X14 VDD1.t1 VP.t4 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4407 pd=3.04 as=0.18645 ps=1.46 w=1.13 l=1
X15 VTAIL.t9 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.18645 pd=1.46 as=0.18645 ps=1.46 w=1.13 l=1
R0 VP.n5 VP.n2 161.3
R1 VP.n13 VP.n0 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n10 VP.n1 161.3
R4 VP.n3 VP.t4 89.1577
R5 VP.n7 VP.n6 80.6037
R6 VP.n15 VP.n14 80.6037
R7 VP.n9 VP.n8 80.6037
R8 VP.n8 VP.t3 66.7575
R9 VP.n14 VP.t1 66.7575
R10 VP.n6 VP.t0 66.7575
R11 VP.n8 VP.n1 48.2005
R12 VP.n14 VP.n13 48.2005
R13 VP.n6 VP.n5 48.2005
R14 VP.n9 VP.n7 34.2552
R15 VP.n4 VP.n3 32.0786
R16 VP.n3 VP.n2 28.4363
R17 VP.n12 VP.t5 27.2335
R18 VP.n4 VP.t2 27.2335
R19 VP.n12 VP.n1 24.4675
R20 VP.n13 VP.n12 24.4675
R21 VP.n5 VP.n4 24.4675
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VTAIL.n11 VTAIL.t5 156.304
R29 VTAIL.n2 VTAIL.t7 156.304
R30 VTAIL.n10 VTAIL.t6 156.304
R31 VTAIL.n7 VTAIL.t0 156.304
R32 VTAIL.n1 VTAIL.n0 130.142
R33 VTAIL.n4 VTAIL.n3 130.142
R34 VTAIL.n9 VTAIL.n8 130.141
R35 VTAIL.n6 VTAIL.n5 130.141
R36 VTAIL.n0 VTAIL.t2 17.5226
R37 VTAIL.n0 VTAIL.t1 17.5226
R38 VTAIL.n3 VTAIL.t8 17.5226
R39 VTAIL.n3 VTAIL.t9 17.5226
R40 VTAIL.n8 VTAIL.t10 17.5226
R41 VTAIL.n8 VTAIL.t11 17.5226
R42 VTAIL.n5 VTAIL.t3 17.5226
R43 VTAIL.n5 VTAIL.t4 17.5226
R44 VTAIL.n6 VTAIL.n4 15.6341
R45 VTAIL.n11 VTAIL.n10 14.4876
R46 VTAIL.n7 VTAIL.n6 1.14705
R47 VTAIL.n10 VTAIL.n9 1.14705
R48 VTAIL.n4 VTAIL.n2 1.14705
R49 VTAIL.n9 VTAIL.n7 1.0436
R50 VTAIL.n2 VTAIL.n1 1.0436
R51 VTAIL VTAIL.n11 0.802224
R52 VTAIL VTAIL.n1 0.345328
R53 VDD1 VDD1.t1 173.9
R54 VDD1.n1 VDD1.t2 173.786
R55 VDD1.n1 VDD1.n0 147.052
R56 VDD1.n3 VDD1.n2 146.821
R57 VDD1.n3 VDD1.n1 29.572
R58 VDD1.n2 VDD1.t3 17.5226
R59 VDD1.n2 VDD1.t5 17.5226
R60 VDD1.n0 VDD1.t0 17.5226
R61 VDD1.n0 VDD1.t4 17.5226
R62 VDD1 VDD1.n3 0.228948
R63 B.n342 B.n341 585
R64 B.n343 B.n342 585
R65 B.n118 B.n60 585
R66 B.n117 B.n116 585
R67 B.n115 B.n114 585
R68 B.n113 B.n112 585
R69 B.n111 B.n110 585
R70 B.n109 B.n108 585
R71 B.n107 B.n106 585
R72 B.n105 B.n104 585
R73 B.n103 B.n102 585
R74 B.n100 B.n99 585
R75 B.n98 B.n97 585
R76 B.n96 B.n95 585
R77 B.n94 B.n93 585
R78 B.n92 B.n91 585
R79 B.n90 B.n89 585
R80 B.n88 B.n87 585
R81 B.n86 B.n85 585
R82 B.n84 B.n83 585
R83 B.n82 B.n81 585
R84 B.n80 B.n79 585
R85 B.n78 B.n77 585
R86 B.n76 B.n75 585
R87 B.n74 B.n73 585
R88 B.n72 B.n71 585
R89 B.n70 B.n69 585
R90 B.n68 B.n67 585
R91 B.n46 B.n45 585
R92 B.n346 B.n345 585
R93 B.n340 B.n61 585
R94 B.n61 B.n43 585
R95 B.n339 B.n42 585
R96 B.n350 B.n42 585
R97 B.n338 B.n41 585
R98 B.n351 B.n41 585
R99 B.n337 B.n40 585
R100 B.n352 B.n40 585
R101 B.n336 B.n335 585
R102 B.n335 B.n36 585
R103 B.n334 B.n35 585
R104 B.t11 B.n35 585
R105 B.n333 B.n34 585
R106 B.n358 B.n34 585
R107 B.n332 B.n33 585
R108 B.n359 B.n33 585
R109 B.n331 B.n330 585
R110 B.n330 B.n29 585
R111 B.n329 B.n28 585
R112 B.n365 B.n28 585
R113 B.n328 B.n27 585
R114 B.n366 B.n27 585
R115 B.n327 B.n26 585
R116 B.n367 B.n26 585
R117 B.n326 B.n325 585
R118 B.n325 B.n25 585
R119 B.n324 B.n21 585
R120 B.n373 B.n21 585
R121 B.n323 B.n20 585
R122 B.n374 B.n20 585
R123 B.n322 B.n19 585
R124 B.n375 B.n19 585
R125 B.n321 B.n320 585
R126 B.n320 B.n18 585
R127 B.n319 B.n14 585
R128 B.n381 B.n14 585
R129 B.n318 B.n13 585
R130 B.n382 B.n13 585
R131 B.n317 B.n12 585
R132 B.n383 B.n12 585
R133 B.n316 B.n315 585
R134 B.n315 B.n314 585
R135 B.n313 B.n312 585
R136 B.n313 B.n8 585
R137 B.n311 B.n7 585
R138 B.n390 B.n7 585
R139 B.n310 B.n6 585
R140 B.n391 B.n6 585
R141 B.n309 B.n5 585
R142 B.n392 B.n5 585
R143 B.n308 B.n307 585
R144 B.n307 B.n4 585
R145 B.n306 B.n119 585
R146 B.n306 B.n305 585
R147 B.n296 B.n120 585
R148 B.n121 B.n120 585
R149 B.n298 B.n297 585
R150 B.n299 B.n298 585
R151 B.n295 B.n126 585
R152 B.n126 B.n125 585
R153 B.n294 B.n293 585
R154 B.n293 B.n292 585
R155 B.n128 B.n127 585
R156 B.n285 B.n128 585
R157 B.n284 B.n283 585
R158 B.n286 B.n284 585
R159 B.n282 B.n133 585
R160 B.n133 B.n132 585
R161 B.n281 B.n280 585
R162 B.n280 B.n279 585
R163 B.n135 B.n134 585
R164 B.n272 B.n135 585
R165 B.n271 B.n270 585
R166 B.n273 B.n271 585
R167 B.n269 B.n140 585
R168 B.n140 B.n139 585
R169 B.n268 B.n267 585
R170 B.n267 B.n266 585
R171 B.n142 B.n141 585
R172 B.n143 B.n142 585
R173 B.n259 B.n258 585
R174 B.n260 B.n259 585
R175 B.n257 B.n148 585
R176 B.n148 B.n147 585
R177 B.n256 B.n255 585
R178 B.n255 B.t7 585
R179 B.n150 B.n149 585
R180 B.n151 B.n150 585
R181 B.n248 B.n247 585
R182 B.n249 B.n248 585
R183 B.n246 B.n156 585
R184 B.n156 B.n155 585
R185 B.n245 B.n244 585
R186 B.n244 B.n243 585
R187 B.n158 B.n157 585
R188 B.n159 B.n158 585
R189 B.n239 B.n238 585
R190 B.n162 B.n161 585
R191 B.n235 B.n234 585
R192 B.n236 B.n235 585
R193 B.n233 B.n176 585
R194 B.n232 B.n231 585
R195 B.n230 B.n229 585
R196 B.n228 B.n227 585
R197 B.n226 B.n225 585
R198 B.n224 B.n223 585
R199 B.n222 B.n221 585
R200 B.n219 B.n218 585
R201 B.n217 B.n216 585
R202 B.n215 B.n214 585
R203 B.n213 B.n212 585
R204 B.n211 B.n210 585
R205 B.n209 B.n208 585
R206 B.n207 B.n206 585
R207 B.n205 B.n204 585
R208 B.n203 B.n202 585
R209 B.n201 B.n200 585
R210 B.n199 B.n198 585
R211 B.n197 B.n196 585
R212 B.n195 B.n194 585
R213 B.n193 B.n192 585
R214 B.n191 B.n190 585
R215 B.n189 B.n188 585
R216 B.n187 B.n186 585
R217 B.n185 B.n184 585
R218 B.n183 B.n182 585
R219 B.n240 B.n160 585
R220 B.n160 B.n159 585
R221 B.n242 B.n241 585
R222 B.n243 B.n242 585
R223 B.n154 B.n153 585
R224 B.n155 B.n154 585
R225 B.n251 B.n250 585
R226 B.n250 B.n249 585
R227 B.n252 B.n152 585
R228 B.n152 B.n151 585
R229 B.n254 B.n253 585
R230 B.t7 B.n254 585
R231 B.n146 B.n145 585
R232 B.n147 B.n146 585
R233 B.n262 B.n261 585
R234 B.n261 B.n260 585
R235 B.n263 B.n144 585
R236 B.n144 B.n143 585
R237 B.n265 B.n264 585
R238 B.n266 B.n265 585
R239 B.n138 B.n137 585
R240 B.n139 B.n138 585
R241 B.n275 B.n274 585
R242 B.n274 B.n273 585
R243 B.n276 B.n136 585
R244 B.n272 B.n136 585
R245 B.n278 B.n277 585
R246 B.n279 B.n278 585
R247 B.n131 B.n130 585
R248 B.n132 B.n131 585
R249 B.n288 B.n287 585
R250 B.n287 B.n286 585
R251 B.n289 B.n129 585
R252 B.n285 B.n129 585
R253 B.n291 B.n290 585
R254 B.n292 B.n291 585
R255 B.n124 B.n123 585
R256 B.n125 B.n124 585
R257 B.n301 B.n300 585
R258 B.n300 B.n299 585
R259 B.n302 B.n122 585
R260 B.n122 B.n121 585
R261 B.n304 B.n303 585
R262 B.n305 B.n304 585
R263 B.n3 B.n0 585
R264 B.n4 B.n3 585
R265 B.n389 B.n1 585
R266 B.n390 B.n389 585
R267 B.n388 B.n387 585
R268 B.n388 B.n8 585
R269 B.n386 B.n9 585
R270 B.n314 B.n9 585
R271 B.n385 B.n384 585
R272 B.n384 B.n383 585
R273 B.n11 B.n10 585
R274 B.n382 B.n11 585
R275 B.n380 B.n379 585
R276 B.n381 B.n380 585
R277 B.n378 B.n15 585
R278 B.n18 B.n15 585
R279 B.n377 B.n376 585
R280 B.n376 B.n375 585
R281 B.n17 B.n16 585
R282 B.n374 B.n17 585
R283 B.n372 B.n371 585
R284 B.n373 B.n372 585
R285 B.n370 B.n22 585
R286 B.n25 B.n22 585
R287 B.n369 B.n368 585
R288 B.n368 B.n367 585
R289 B.n24 B.n23 585
R290 B.n366 B.n24 585
R291 B.n364 B.n363 585
R292 B.n365 B.n364 585
R293 B.n362 B.n30 585
R294 B.n30 B.n29 585
R295 B.n361 B.n360 585
R296 B.n360 B.n359 585
R297 B.n32 B.n31 585
R298 B.n358 B.n32 585
R299 B.n357 B.n356 585
R300 B.t11 B.n357 585
R301 B.n355 B.n37 585
R302 B.n37 B.n36 585
R303 B.n354 B.n353 585
R304 B.n353 B.n352 585
R305 B.n39 B.n38 585
R306 B.n351 B.n39 585
R307 B.n349 B.n348 585
R308 B.n350 B.n349 585
R309 B.n347 B.n44 585
R310 B.n44 B.n43 585
R311 B.n393 B.n392 585
R312 B.n391 B.n2 585
R313 B.n345 B.n44 530.939
R314 B.n342 B.n61 530.939
R315 B.n182 B.n158 530.939
R316 B.n238 B.n160 530.939
R317 B.n343 B.n59 256.663
R318 B.n343 B.n58 256.663
R319 B.n343 B.n57 256.663
R320 B.n343 B.n56 256.663
R321 B.n343 B.n55 256.663
R322 B.n343 B.n54 256.663
R323 B.n343 B.n53 256.663
R324 B.n343 B.n52 256.663
R325 B.n343 B.n51 256.663
R326 B.n343 B.n50 256.663
R327 B.n343 B.n49 256.663
R328 B.n343 B.n48 256.663
R329 B.n343 B.n47 256.663
R330 B.n344 B.n343 256.663
R331 B.n237 B.n236 256.663
R332 B.n236 B.n163 256.663
R333 B.n236 B.n164 256.663
R334 B.n236 B.n165 256.663
R335 B.n236 B.n166 256.663
R336 B.n236 B.n167 256.663
R337 B.n236 B.n168 256.663
R338 B.n236 B.n169 256.663
R339 B.n236 B.n170 256.663
R340 B.n236 B.n171 256.663
R341 B.n236 B.n172 256.663
R342 B.n236 B.n173 256.663
R343 B.n236 B.n174 256.663
R344 B.n236 B.n175 256.663
R345 B.n395 B.n394 256.663
R346 B.n236 B.n159 242.155
R347 B.n343 B.n43 242.155
R348 B.n64 B.t10 230.159
R349 B.n62 B.t17 230.159
R350 B.n179 B.t6 230.159
R351 B.n177 B.t14 230.159
R352 B.n64 B.t12 172.675
R353 B.n177 B.t16 172.675
R354 B.n62 B.t18 172.675
R355 B.n179 B.t9 172.675
R356 B.n67 B.n46 163.367
R357 B.n71 B.n70 163.367
R358 B.n75 B.n74 163.367
R359 B.n79 B.n78 163.367
R360 B.n83 B.n82 163.367
R361 B.n87 B.n86 163.367
R362 B.n91 B.n90 163.367
R363 B.n95 B.n94 163.367
R364 B.n99 B.n98 163.367
R365 B.n104 B.n103 163.367
R366 B.n108 B.n107 163.367
R367 B.n112 B.n111 163.367
R368 B.n116 B.n115 163.367
R369 B.n342 B.n60 163.367
R370 B.n244 B.n158 163.367
R371 B.n244 B.n156 163.367
R372 B.n248 B.n156 163.367
R373 B.n248 B.n150 163.367
R374 B.n255 B.n150 163.367
R375 B.n255 B.n148 163.367
R376 B.n259 B.n148 163.367
R377 B.n259 B.n142 163.367
R378 B.n267 B.n142 163.367
R379 B.n267 B.n140 163.367
R380 B.n271 B.n140 163.367
R381 B.n271 B.n135 163.367
R382 B.n280 B.n135 163.367
R383 B.n280 B.n133 163.367
R384 B.n284 B.n133 163.367
R385 B.n284 B.n128 163.367
R386 B.n293 B.n128 163.367
R387 B.n293 B.n126 163.367
R388 B.n298 B.n126 163.367
R389 B.n298 B.n120 163.367
R390 B.n306 B.n120 163.367
R391 B.n307 B.n306 163.367
R392 B.n307 B.n5 163.367
R393 B.n6 B.n5 163.367
R394 B.n7 B.n6 163.367
R395 B.n313 B.n7 163.367
R396 B.n315 B.n313 163.367
R397 B.n315 B.n12 163.367
R398 B.n13 B.n12 163.367
R399 B.n14 B.n13 163.367
R400 B.n320 B.n14 163.367
R401 B.n320 B.n19 163.367
R402 B.n20 B.n19 163.367
R403 B.n21 B.n20 163.367
R404 B.n325 B.n21 163.367
R405 B.n325 B.n26 163.367
R406 B.n27 B.n26 163.367
R407 B.n28 B.n27 163.367
R408 B.n330 B.n28 163.367
R409 B.n330 B.n33 163.367
R410 B.n34 B.n33 163.367
R411 B.n35 B.n34 163.367
R412 B.n335 B.n35 163.367
R413 B.n335 B.n40 163.367
R414 B.n41 B.n40 163.367
R415 B.n42 B.n41 163.367
R416 B.n61 B.n42 163.367
R417 B.n235 B.n162 163.367
R418 B.n235 B.n176 163.367
R419 B.n231 B.n230 163.367
R420 B.n227 B.n226 163.367
R421 B.n223 B.n222 163.367
R422 B.n218 B.n217 163.367
R423 B.n214 B.n213 163.367
R424 B.n210 B.n209 163.367
R425 B.n206 B.n205 163.367
R426 B.n202 B.n201 163.367
R427 B.n198 B.n197 163.367
R428 B.n194 B.n193 163.367
R429 B.n190 B.n189 163.367
R430 B.n186 B.n185 163.367
R431 B.n242 B.n160 163.367
R432 B.n242 B.n154 163.367
R433 B.n250 B.n154 163.367
R434 B.n250 B.n152 163.367
R435 B.n254 B.n152 163.367
R436 B.n254 B.n146 163.367
R437 B.n261 B.n146 163.367
R438 B.n261 B.n144 163.367
R439 B.n265 B.n144 163.367
R440 B.n265 B.n138 163.367
R441 B.n274 B.n138 163.367
R442 B.n274 B.n136 163.367
R443 B.n278 B.n136 163.367
R444 B.n278 B.n131 163.367
R445 B.n287 B.n131 163.367
R446 B.n287 B.n129 163.367
R447 B.n291 B.n129 163.367
R448 B.n291 B.n124 163.367
R449 B.n300 B.n124 163.367
R450 B.n300 B.n122 163.367
R451 B.n304 B.n122 163.367
R452 B.n304 B.n3 163.367
R453 B.n393 B.n3 163.367
R454 B.n389 B.n2 163.367
R455 B.n389 B.n388 163.367
R456 B.n388 B.n9 163.367
R457 B.n384 B.n9 163.367
R458 B.n384 B.n11 163.367
R459 B.n380 B.n11 163.367
R460 B.n380 B.n15 163.367
R461 B.n376 B.n15 163.367
R462 B.n376 B.n17 163.367
R463 B.n372 B.n17 163.367
R464 B.n372 B.n22 163.367
R465 B.n368 B.n22 163.367
R466 B.n368 B.n24 163.367
R467 B.n364 B.n24 163.367
R468 B.n364 B.n30 163.367
R469 B.n360 B.n30 163.367
R470 B.n360 B.n32 163.367
R471 B.n357 B.n32 163.367
R472 B.n357 B.n37 163.367
R473 B.n353 B.n37 163.367
R474 B.n353 B.n39 163.367
R475 B.n349 B.n39 163.367
R476 B.n349 B.n44 163.367
R477 B.n65 B.t13 146.881
R478 B.n63 B.t19 146.881
R479 B.n180 B.t8 146.881
R480 B.n178 B.t15 146.881
R481 B.n243 B.n159 116.784
R482 B.n243 B.n155 116.784
R483 B.n249 B.n155 116.784
R484 B.n249 B.n151 116.784
R485 B.t7 B.n151 116.784
R486 B.t7 B.n147 116.784
R487 B.n260 B.n147 116.784
R488 B.n260 B.n143 116.784
R489 B.n266 B.n143 116.784
R490 B.n266 B.n139 116.784
R491 B.n273 B.n139 116.784
R492 B.n273 B.n272 116.784
R493 B.n279 B.n132 116.784
R494 B.n286 B.n132 116.784
R495 B.n286 B.n285 116.784
R496 B.n292 B.n125 116.784
R497 B.n299 B.n125 116.784
R498 B.n305 B.n121 116.784
R499 B.n305 B.n4 116.784
R500 B.n392 B.n4 116.784
R501 B.n392 B.n391 116.784
R502 B.n391 B.n390 116.784
R503 B.n390 B.n8 116.784
R504 B.n314 B.n8 116.784
R505 B.n383 B.n382 116.784
R506 B.n382 B.n381 116.784
R507 B.n375 B.n18 116.784
R508 B.n375 B.n374 116.784
R509 B.n374 B.n373 116.784
R510 B.n367 B.n25 116.784
R511 B.n367 B.n366 116.784
R512 B.n366 B.n365 116.784
R513 B.n365 B.n29 116.784
R514 B.n359 B.n29 116.784
R515 B.n359 B.n358 116.784
R516 B.n358 B.t11 116.784
R517 B.t11 B.n36 116.784
R518 B.n352 B.n36 116.784
R519 B.n352 B.n351 116.784
R520 B.n351 B.n350 116.784
R521 B.n350 B.n43 116.784
R522 B.n292 B.t4 113.35
R523 B.n381 B.t1 113.35
R524 B.n299 B.t0 109.915
R525 B.n383 B.t2 109.915
R526 B.n279 B.t3 103.046
R527 B.n373 B.t5 103.046
R528 B.n345 B.n344 71.676
R529 B.n67 B.n47 71.676
R530 B.n71 B.n48 71.676
R531 B.n75 B.n49 71.676
R532 B.n79 B.n50 71.676
R533 B.n83 B.n51 71.676
R534 B.n87 B.n52 71.676
R535 B.n91 B.n53 71.676
R536 B.n95 B.n54 71.676
R537 B.n99 B.n55 71.676
R538 B.n104 B.n56 71.676
R539 B.n108 B.n57 71.676
R540 B.n112 B.n58 71.676
R541 B.n116 B.n59 71.676
R542 B.n60 B.n59 71.676
R543 B.n115 B.n58 71.676
R544 B.n111 B.n57 71.676
R545 B.n107 B.n56 71.676
R546 B.n103 B.n55 71.676
R547 B.n98 B.n54 71.676
R548 B.n94 B.n53 71.676
R549 B.n90 B.n52 71.676
R550 B.n86 B.n51 71.676
R551 B.n82 B.n50 71.676
R552 B.n78 B.n49 71.676
R553 B.n74 B.n48 71.676
R554 B.n70 B.n47 71.676
R555 B.n344 B.n46 71.676
R556 B.n238 B.n237 71.676
R557 B.n176 B.n163 71.676
R558 B.n230 B.n164 71.676
R559 B.n226 B.n165 71.676
R560 B.n222 B.n166 71.676
R561 B.n217 B.n167 71.676
R562 B.n213 B.n168 71.676
R563 B.n209 B.n169 71.676
R564 B.n205 B.n170 71.676
R565 B.n201 B.n171 71.676
R566 B.n197 B.n172 71.676
R567 B.n193 B.n173 71.676
R568 B.n189 B.n174 71.676
R569 B.n185 B.n175 71.676
R570 B.n237 B.n162 71.676
R571 B.n231 B.n163 71.676
R572 B.n227 B.n164 71.676
R573 B.n223 B.n165 71.676
R574 B.n218 B.n166 71.676
R575 B.n214 B.n167 71.676
R576 B.n210 B.n168 71.676
R577 B.n206 B.n169 71.676
R578 B.n202 B.n170 71.676
R579 B.n198 B.n171 71.676
R580 B.n194 B.n172 71.676
R581 B.n190 B.n173 71.676
R582 B.n186 B.n174 71.676
R583 B.n182 B.n175 71.676
R584 B.n394 B.n393 71.676
R585 B.n394 B.n2 71.676
R586 B.n66 B.n65 59.5399
R587 B.n101 B.n63 59.5399
R588 B.n181 B.n180 59.5399
R589 B.n220 B.n178 59.5399
R590 B.n240 B.n239 34.4981
R591 B.n183 B.n157 34.4981
R592 B.n341 B.n340 34.4981
R593 B.n347 B.n346 34.4981
R594 B.n65 B.n64 25.7944
R595 B.n63 B.n62 25.7944
R596 B.n180 B.n179 25.7944
R597 B.n178 B.n177 25.7944
R598 B B.n395 18.0485
R599 B.n272 B.t3 13.7398
R600 B.n25 B.t5 13.7398
R601 B.n241 B.n240 10.6151
R602 B.n241 B.n153 10.6151
R603 B.n251 B.n153 10.6151
R604 B.n252 B.n251 10.6151
R605 B.n253 B.n252 10.6151
R606 B.n253 B.n145 10.6151
R607 B.n262 B.n145 10.6151
R608 B.n263 B.n262 10.6151
R609 B.n264 B.n263 10.6151
R610 B.n264 B.n137 10.6151
R611 B.n275 B.n137 10.6151
R612 B.n276 B.n275 10.6151
R613 B.n277 B.n276 10.6151
R614 B.n277 B.n130 10.6151
R615 B.n288 B.n130 10.6151
R616 B.n289 B.n288 10.6151
R617 B.n290 B.n289 10.6151
R618 B.n290 B.n123 10.6151
R619 B.n301 B.n123 10.6151
R620 B.n302 B.n301 10.6151
R621 B.n303 B.n302 10.6151
R622 B.n303 B.n0 10.6151
R623 B.n239 B.n161 10.6151
R624 B.n234 B.n161 10.6151
R625 B.n234 B.n233 10.6151
R626 B.n233 B.n232 10.6151
R627 B.n232 B.n229 10.6151
R628 B.n229 B.n228 10.6151
R629 B.n228 B.n225 10.6151
R630 B.n225 B.n224 10.6151
R631 B.n224 B.n221 10.6151
R632 B.n219 B.n216 10.6151
R633 B.n216 B.n215 10.6151
R634 B.n215 B.n212 10.6151
R635 B.n212 B.n211 10.6151
R636 B.n211 B.n208 10.6151
R637 B.n208 B.n207 10.6151
R638 B.n207 B.n204 10.6151
R639 B.n204 B.n203 10.6151
R640 B.n200 B.n199 10.6151
R641 B.n199 B.n196 10.6151
R642 B.n196 B.n195 10.6151
R643 B.n195 B.n192 10.6151
R644 B.n192 B.n191 10.6151
R645 B.n191 B.n188 10.6151
R646 B.n188 B.n187 10.6151
R647 B.n187 B.n184 10.6151
R648 B.n184 B.n183 10.6151
R649 B.n245 B.n157 10.6151
R650 B.n246 B.n245 10.6151
R651 B.n247 B.n246 10.6151
R652 B.n247 B.n149 10.6151
R653 B.n256 B.n149 10.6151
R654 B.n257 B.n256 10.6151
R655 B.n258 B.n257 10.6151
R656 B.n258 B.n141 10.6151
R657 B.n268 B.n141 10.6151
R658 B.n269 B.n268 10.6151
R659 B.n270 B.n269 10.6151
R660 B.n270 B.n134 10.6151
R661 B.n281 B.n134 10.6151
R662 B.n282 B.n281 10.6151
R663 B.n283 B.n282 10.6151
R664 B.n283 B.n127 10.6151
R665 B.n294 B.n127 10.6151
R666 B.n295 B.n294 10.6151
R667 B.n297 B.n295 10.6151
R668 B.n297 B.n296 10.6151
R669 B.n296 B.n119 10.6151
R670 B.n308 B.n119 10.6151
R671 B.n309 B.n308 10.6151
R672 B.n310 B.n309 10.6151
R673 B.n311 B.n310 10.6151
R674 B.n312 B.n311 10.6151
R675 B.n316 B.n312 10.6151
R676 B.n317 B.n316 10.6151
R677 B.n318 B.n317 10.6151
R678 B.n319 B.n318 10.6151
R679 B.n321 B.n319 10.6151
R680 B.n322 B.n321 10.6151
R681 B.n323 B.n322 10.6151
R682 B.n324 B.n323 10.6151
R683 B.n326 B.n324 10.6151
R684 B.n327 B.n326 10.6151
R685 B.n328 B.n327 10.6151
R686 B.n329 B.n328 10.6151
R687 B.n331 B.n329 10.6151
R688 B.n332 B.n331 10.6151
R689 B.n333 B.n332 10.6151
R690 B.n334 B.n333 10.6151
R691 B.n336 B.n334 10.6151
R692 B.n337 B.n336 10.6151
R693 B.n338 B.n337 10.6151
R694 B.n339 B.n338 10.6151
R695 B.n340 B.n339 10.6151
R696 B.n387 B.n1 10.6151
R697 B.n387 B.n386 10.6151
R698 B.n386 B.n385 10.6151
R699 B.n385 B.n10 10.6151
R700 B.n379 B.n10 10.6151
R701 B.n379 B.n378 10.6151
R702 B.n378 B.n377 10.6151
R703 B.n377 B.n16 10.6151
R704 B.n371 B.n16 10.6151
R705 B.n371 B.n370 10.6151
R706 B.n370 B.n369 10.6151
R707 B.n369 B.n23 10.6151
R708 B.n363 B.n23 10.6151
R709 B.n363 B.n362 10.6151
R710 B.n362 B.n361 10.6151
R711 B.n361 B.n31 10.6151
R712 B.n356 B.n31 10.6151
R713 B.n356 B.n355 10.6151
R714 B.n355 B.n354 10.6151
R715 B.n354 B.n38 10.6151
R716 B.n348 B.n38 10.6151
R717 B.n348 B.n347 10.6151
R718 B.n346 B.n45 10.6151
R719 B.n68 B.n45 10.6151
R720 B.n69 B.n68 10.6151
R721 B.n72 B.n69 10.6151
R722 B.n73 B.n72 10.6151
R723 B.n76 B.n73 10.6151
R724 B.n77 B.n76 10.6151
R725 B.n80 B.n77 10.6151
R726 B.n81 B.n80 10.6151
R727 B.n85 B.n84 10.6151
R728 B.n88 B.n85 10.6151
R729 B.n89 B.n88 10.6151
R730 B.n92 B.n89 10.6151
R731 B.n93 B.n92 10.6151
R732 B.n96 B.n93 10.6151
R733 B.n97 B.n96 10.6151
R734 B.n100 B.n97 10.6151
R735 B.n105 B.n102 10.6151
R736 B.n106 B.n105 10.6151
R737 B.n109 B.n106 10.6151
R738 B.n110 B.n109 10.6151
R739 B.n113 B.n110 10.6151
R740 B.n114 B.n113 10.6151
R741 B.n117 B.n114 10.6151
R742 B.n118 B.n117 10.6151
R743 B.n341 B.n118 10.6151
R744 B.n395 B.n0 8.11757
R745 B.n395 B.n1 8.11757
R746 B.t0 B.n121 6.87013
R747 B.n314 B.t2 6.87013
R748 B.n220 B.n219 6.5566
R749 B.n203 B.n181 6.5566
R750 B.n84 B.n66 6.5566
R751 B.n101 B.n100 6.5566
R752 B.n221 B.n220 4.05904
R753 B.n200 B.n181 4.05904
R754 B.n81 B.n66 4.05904
R755 B.n102 B.n101 4.05904
R756 B.n285 B.t4 3.43532
R757 B.n18 B.t1 3.43532
R758 VN.n9 VN.n6 161.3
R759 VN.n3 VN.n0 161.3
R760 VN.n7 VN.t1 89.1577
R761 VN.n1 VN.t3 89.1577
R762 VN.n11 VN.n10 80.6037
R763 VN.n5 VN.n4 80.6037
R764 VN.n4 VN.t0 66.7575
R765 VN.n10 VN.t4 66.7575
R766 VN.n4 VN.n3 48.2005
R767 VN.n10 VN.n9 48.2005
R768 VN VN.n11 34.5407
R769 VN.n8 VN.n7 32.0786
R770 VN.n2 VN.n1 32.0786
R771 VN.n7 VN.n6 28.4363
R772 VN.n1 VN.n0 28.4363
R773 VN.n2 VN.t2 27.2335
R774 VN.n8 VN.t5 27.2335
R775 VN.n3 VN.n2 24.4675
R776 VN.n9 VN.n8 24.4675
R777 VN.n11 VN.n6 0.285035
R778 VN.n5 VN.n0 0.285035
R779 VN VN.n5 0.146778
R780 VDD2.n1 VDD2.t2 173.786
R781 VDD2.n2 VDD2.t1 172.982
R782 VDD2.n1 VDD2.n0 147.052
R783 VDD2 VDD2.n3 147.048
R784 VDD2.n2 VDD2.n1 28.4157
R785 VDD2.n3 VDD2.t0 17.5226
R786 VDD2.n3 VDD2.t4 17.5226
R787 VDD2.n0 VDD2.t3 17.5226
R788 VDD2.n0 VDD2.t5 17.5226
R789 VDD2 VDD2.n2 0.918603
C0 VDD2 VP 0.33034f
C1 VP VDD1 0.966559f
C2 VP VTAIL 1.1903f
C3 VDD2 VN 0.794582f
C4 VN VDD1 0.156256f
C5 VN VTAIL 1.17615f
C6 VDD2 VDD1 0.81828f
C7 VDD2 VTAIL 2.77387f
C8 VN VP 3.37123f
C9 VTAIL VDD1 2.7316f
C10 VDD2 B 2.657289f
C11 VDD1 B 2.85567f
C12 VTAIL B 2.254191f
C13 VN B 6.753272f
C14 VP B 5.756616f
C15 VDD2.t2 B 0.110889f
C16 VDD2.t3 B 0.016241f
C17 VDD2.t5 B 0.016241f
C18 VDD2.n0 B 0.083574f
C19 VDD2.n1 B 1.05971f
C20 VDD2.t1 B 0.110009f
C21 VDD2.n2 B 1.01493f
C22 VDD2.t0 B 0.016241f
C23 VDD2.t4 B 0.016241f
C24 VDD2.n3 B 0.083567f
C25 VN.n0 B 0.159327f
C26 VN.t2 B 0.066037f
C27 VN.t3 B 0.138738f
C28 VN.n1 B 0.092363f
C29 VN.n2 B 0.104076f
C30 VN.n3 B 0.033928f
C31 VN.t0 B 0.111351f
C32 VN.n4 B 0.102178f
C33 VN.n5 B 0.027701f
C34 VN.n6 B 0.159327f
C35 VN.t5 B 0.066037f
C36 VN.t1 B 0.138738f
C37 VN.n7 B 0.092363f
C38 VN.n8 B 0.104076f
C39 VN.n9 B 0.033928f
C40 VN.t4 B 0.111351f
C41 VN.n10 B 0.102178f
C42 VN.n11 B 0.872951f
C43 VDD1.t1 B 0.10457f
C44 VDD1.t2 B 0.104423f
C45 VDD1.t0 B 0.015294f
C46 VDD1.t4 B 0.015294f
C47 VDD1.n0 B 0.078701f
C48 VDD1.n1 B 1.05068f
C49 VDD1.t3 B 0.015294f
C50 VDD1.t5 B 0.015294f
C51 VDD1.n2 B 0.078394f
C52 VDD1.n3 B 0.974956f
C53 VTAIL.t2 B 0.021693f
C54 VTAIL.t1 B 0.021693f
C55 VTAIL.n0 B 0.091658f
C56 VTAIL.n1 B 0.252197f
C57 VTAIL.t7 B 0.128172f
C58 VTAIL.n2 B 0.337604f
C59 VTAIL.t8 B 0.021693f
C60 VTAIL.t9 B 0.021693f
C61 VTAIL.n3 B 0.091658f
C62 VTAIL.n4 B 0.819055f
C63 VTAIL.t3 B 0.021693f
C64 VTAIL.t4 B 0.021693f
C65 VTAIL.n5 B 0.091658f
C66 VTAIL.n6 B 0.819056f
C67 VTAIL.t0 B 0.128172f
C68 VTAIL.n7 B 0.337604f
C69 VTAIL.t10 B 0.021693f
C70 VTAIL.t11 B 0.021693f
C71 VTAIL.n8 B 0.091658f
C72 VTAIL.n9 B 0.314955f
C73 VTAIL.t6 B 0.128172f
C74 VTAIL.n10 B 0.751954f
C75 VTAIL.t5 B 0.128172f
C76 VTAIL.n11 B 0.724961f
C77 VP.n0 B 0.039957f
C78 VP.t5 B 0.066854f
C79 VP.n1 B 0.034348f
C80 VP.n2 B 0.1613f
C81 VP.t0 B 0.112729f
C82 VP.t2 B 0.066854f
C83 VP.t4 B 0.140455f
C84 VP.n3 B 0.093506f
C85 VP.n4 B 0.105365f
C86 VP.n5 B 0.034348f
C87 VP.n6 B 0.103443f
C88 VP.n7 B 0.866287f
C89 VP.t3 B 0.112729f
C90 VP.n8 B 0.103443f
C91 VP.n9 B 0.89771f
C92 VP.n10 B 0.039957f
C93 VP.n11 B 0.029944f
C94 VP.n12 B 0.087418f
C95 VP.n13 B 0.034348f
C96 VP.t1 B 0.112729f
C97 VP.n14 B 0.103443f
C98 VP.n15 B 0.028044f
.ends

