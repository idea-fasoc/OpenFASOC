* NGSPICE file created from diff_pair_sample_0999.ext - technology: sky130A

.subckt diff_pair_sample_0999 VTAIL VN VP B VDD2 VDD1
X0 B.t16 B.t14 B.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0 ps=0 w=0.89 l=0.74
X1 VTAIL.t7 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0.14685 ps=1.22 w=0.89 l=0.74
X2 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0 ps=0 w=0.89 l=0.74
X3 VDD2.t0 VN.t1 VTAIL.t6 B.t17 sky130_fd_pr__nfet_01v8 ad=0.14685 pd=1.22 as=0.3471 ps=2.56 w=0.89 l=0.74
X4 VTAIL.t5 VN.t2 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0.14685 ps=1.22 w=0.89 l=0.74
X5 VDD1.t3 VP.t0 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.14685 pd=1.22 as=0.3471 ps=2.56 w=0.89 l=0.74
X6 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0.14685 ps=1.22 w=0.89 l=0.74
X7 VDD2.t1 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.14685 pd=1.22 as=0.3471 ps=2.56 w=0.89 l=0.74
X8 VTAIL.t2 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0.14685 ps=1.22 w=0.89 l=0.74
X9 VDD1.t0 VP.t3 VTAIL.t1 B.t17 sky130_fd_pr__nfet_01v8 ad=0.14685 pd=1.22 as=0.3471 ps=2.56 w=0.89 l=0.74
X10 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0 ps=0 w=0.89 l=0.74
X11 B.t6 B.t3 B.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3471 pd=2.56 as=0 ps=0 w=0.89 l=0.74
R0 B.n288 B.n287 585
R1 B.n289 B.n288 585
R2 B.n106 B.n49 585
R3 B.n105 B.n104 585
R4 B.n103 B.n102 585
R5 B.n101 B.n100 585
R6 B.n99 B.n98 585
R7 B.n97 B.n96 585
R8 B.n95 B.n94 585
R9 B.n93 B.n92 585
R10 B.n91 B.n90 585
R11 B.n89 B.n88 585
R12 B.n87 B.n86 585
R13 B.n85 B.n84 585
R14 B.n83 B.n82 585
R15 B.n81 B.n80 585
R16 B.n79 B.n78 585
R17 B.n77 B.n76 585
R18 B.n75 B.n74 585
R19 B.n72 B.n71 585
R20 B.n70 B.n69 585
R21 B.n68 B.n67 585
R22 B.n66 B.n65 585
R23 B.n64 B.n63 585
R24 B.n62 B.n61 585
R25 B.n60 B.n59 585
R26 B.n58 B.n57 585
R27 B.n56 B.n55 585
R28 B.n286 B.n35 585
R29 B.n290 B.n35 585
R30 B.n285 B.n34 585
R31 B.n291 B.n34 585
R32 B.n284 B.n283 585
R33 B.n283 B.n30 585
R34 B.n282 B.n29 585
R35 B.n297 B.n29 585
R36 B.n281 B.n28 585
R37 B.n298 B.n28 585
R38 B.n280 B.n27 585
R39 B.n299 B.n27 585
R40 B.n279 B.n278 585
R41 B.n278 B.n23 585
R42 B.n277 B.n22 585
R43 B.n305 B.n22 585
R44 B.n276 B.n21 585
R45 B.n306 B.n21 585
R46 B.n275 B.n20 585
R47 B.n307 B.n20 585
R48 B.n274 B.n273 585
R49 B.n273 B.n16 585
R50 B.n272 B.n15 585
R51 B.n313 B.n15 585
R52 B.n271 B.n14 585
R53 B.n314 B.n14 585
R54 B.n270 B.n13 585
R55 B.n315 B.n13 585
R56 B.n269 B.n268 585
R57 B.n268 B.n12 585
R58 B.n267 B.n266 585
R59 B.n267 B.n8 585
R60 B.n265 B.n7 585
R61 B.n322 B.n7 585
R62 B.n264 B.n6 585
R63 B.n323 B.n6 585
R64 B.n263 B.n5 585
R65 B.n324 B.n5 585
R66 B.n262 B.n261 585
R67 B.n261 B.n4 585
R68 B.n260 B.n107 585
R69 B.n260 B.n259 585
R70 B.n249 B.n108 585
R71 B.n252 B.n108 585
R72 B.n251 B.n250 585
R73 B.n253 B.n251 585
R74 B.n248 B.n113 585
R75 B.n113 B.n112 585
R76 B.n247 B.n246 585
R77 B.n246 B.n245 585
R78 B.n115 B.n114 585
R79 B.n116 B.n115 585
R80 B.n238 B.n237 585
R81 B.n239 B.n238 585
R82 B.n236 B.n121 585
R83 B.n121 B.n120 585
R84 B.n235 B.n234 585
R85 B.n234 B.n233 585
R86 B.n123 B.n122 585
R87 B.n124 B.n123 585
R88 B.n226 B.n225 585
R89 B.n227 B.n226 585
R90 B.n224 B.n128 585
R91 B.n132 B.n128 585
R92 B.n223 B.n222 585
R93 B.n222 B.n221 585
R94 B.n130 B.n129 585
R95 B.n131 B.n130 585
R96 B.n214 B.n213 585
R97 B.n215 B.n214 585
R98 B.n212 B.n137 585
R99 B.n137 B.n136 585
R100 B.n206 B.n205 585
R101 B.n204 B.n152 585
R102 B.n203 B.n151 585
R103 B.n208 B.n151 585
R104 B.n202 B.n201 585
R105 B.n200 B.n199 585
R106 B.n198 B.n197 585
R107 B.n196 B.n195 585
R108 B.n194 B.n193 585
R109 B.n192 B.n191 585
R110 B.n190 B.n189 585
R111 B.n188 B.n187 585
R112 B.n186 B.n185 585
R113 B.n184 B.n183 585
R114 B.n182 B.n181 585
R115 B.n180 B.n179 585
R116 B.n178 B.n177 585
R117 B.n176 B.n175 585
R118 B.n174 B.n173 585
R119 B.n171 B.n170 585
R120 B.n169 B.n168 585
R121 B.n167 B.n166 585
R122 B.n165 B.n164 585
R123 B.n163 B.n162 585
R124 B.n161 B.n160 585
R125 B.n159 B.n158 585
R126 B.n139 B.n138 585
R127 B.n211 B.n210 585
R128 B.n135 B.n134 585
R129 B.n136 B.n135 585
R130 B.n217 B.n216 585
R131 B.n216 B.n215 585
R132 B.n218 B.n133 585
R133 B.n133 B.n131 585
R134 B.n220 B.n219 585
R135 B.n221 B.n220 585
R136 B.n127 B.n126 585
R137 B.n132 B.n127 585
R138 B.n229 B.n228 585
R139 B.n228 B.n227 585
R140 B.n230 B.n125 585
R141 B.n125 B.n124 585
R142 B.n232 B.n231 585
R143 B.n233 B.n232 585
R144 B.n119 B.n118 585
R145 B.n120 B.n119 585
R146 B.n241 B.n240 585
R147 B.n240 B.n239 585
R148 B.n242 B.n117 585
R149 B.n117 B.n116 585
R150 B.n244 B.n243 585
R151 B.n245 B.n244 585
R152 B.n111 B.n110 585
R153 B.n112 B.n111 585
R154 B.n255 B.n254 585
R155 B.n254 B.n253 585
R156 B.n256 B.n109 585
R157 B.n252 B.n109 585
R158 B.n258 B.n257 585
R159 B.n259 B.n258 585
R160 B.n3 B.n0 585
R161 B.n4 B.n3 585
R162 B.n321 B.n1 585
R163 B.n322 B.n321 585
R164 B.n320 B.n319 585
R165 B.n320 B.n8 585
R166 B.n318 B.n9 585
R167 B.n12 B.n9 585
R168 B.n317 B.n316 585
R169 B.n316 B.n315 585
R170 B.n11 B.n10 585
R171 B.n314 B.n11 585
R172 B.n312 B.n311 585
R173 B.n313 B.n312 585
R174 B.n310 B.n17 585
R175 B.n17 B.n16 585
R176 B.n309 B.n308 585
R177 B.n308 B.n307 585
R178 B.n19 B.n18 585
R179 B.n306 B.n19 585
R180 B.n304 B.n303 585
R181 B.n305 B.n304 585
R182 B.n302 B.n24 585
R183 B.n24 B.n23 585
R184 B.n301 B.n300 585
R185 B.n300 B.n299 585
R186 B.n26 B.n25 585
R187 B.n298 B.n26 585
R188 B.n296 B.n295 585
R189 B.n297 B.n296 585
R190 B.n294 B.n31 585
R191 B.n31 B.n30 585
R192 B.n293 B.n292 585
R193 B.n292 B.n291 585
R194 B.n33 B.n32 585
R195 B.n290 B.n33 585
R196 B.n325 B.n324 585
R197 B.n323 B.n2 585
R198 B.n55 B.n33 545.355
R199 B.n288 B.n35 545.355
R200 B.n210 B.n137 545.355
R201 B.n206 B.n135 545.355
R202 B.n289 B.n48 256.663
R203 B.n289 B.n47 256.663
R204 B.n289 B.n46 256.663
R205 B.n289 B.n45 256.663
R206 B.n289 B.n44 256.663
R207 B.n289 B.n43 256.663
R208 B.n289 B.n42 256.663
R209 B.n289 B.n41 256.663
R210 B.n289 B.n40 256.663
R211 B.n289 B.n39 256.663
R212 B.n289 B.n38 256.663
R213 B.n289 B.n37 256.663
R214 B.n289 B.n36 256.663
R215 B.n208 B.n207 256.663
R216 B.n208 B.n140 256.663
R217 B.n208 B.n141 256.663
R218 B.n208 B.n142 256.663
R219 B.n208 B.n143 256.663
R220 B.n208 B.n144 256.663
R221 B.n208 B.n145 256.663
R222 B.n208 B.n146 256.663
R223 B.n208 B.n147 256.663
R224 B.n208 B.n148 256.663
R225 B.n208 B.n149 256.663
R226 B.n208 B.n150 256.663
R227 B.n209 B.n208 256.663
R228 B.n327 B.n326 256.663
R229 B.n53 B.t15 255.15
R230 B.n50 B.t5 255.15
R231 B.n156 B.t13 255.15
R232 B.n153 B.t10 255.15
R233 B.n54 B.t16 234.399
R234 B.n51 B.t6 234.399
R235 B.n157 B.t12 234.399
R236 B.n154 B.t9 234.399
R237 B.n50 B.t3 232.215
R238 B.n156 B.t11 232.215
R239 B.n53 B.t14 231.81
R240 B.n153 B.t7 231.81
R241 B.n208 B.n136 226.602
R242 B.n290 B.n289 226.602
R243 B.n59 B.n58 163.367
R244 B.n63 B.n62 163.367
R245 B.n67 B.n66 163.367
R246 B.n71 B.n70 163.367
R247 B.n76 B.n75 163.367
R248 B.n80 B.n79 163.367
R249 B.n84 B.n83 163.367
R250 B.n88 B.n87 163.367
R251 B.n92 B.n91 163.367
R252 B.n96 B.n95 163.367
R253 B.n100 B.n99 163.367
R254 B.n104 B.n103 163.367
R255 B.n288 B.n49 163.367
R256 B.n214 B.n137 163.367
R257 B.n214 B.n130 163.367
R258 B.n222 B.n130 163.367
R259 B.n222 B.n128 163.367
R260 B.n226 B.n128 163.367
R261 B.n226 B.n123 163.367
R262 B.n234 B.n123 163.367
R263 B.n234 B.n121 163.367
R264 B.n238 B.n121 163.367
R265 B.n238 B.n115 163.367
R266 B.n246 B.n115 163.367
R267 B.n246 B.n113 163.367
R268 B.n251 B.n113 163.367
R269 B.n251 B.n108 163.367
R270 B.n260 B.n108 163.367
R271 B.n261 B.n260 163.367
R272 B.n261 B.n5 163.367
R273 B.n6 B.n5 163.367
R274 B.n7 B.n6 163.367
R275 B.n267 B.n7 163.367
R276 B.n268 B.n267 163.367
R277 B.n268 B.n13 163.367
R278 B.n14 B.n13 163.367
R279 B.n15 B.n14 163.367
R280 B.n273 B.n15 163.367
R281 B.n273 B.n20 163.367
R282 B.n21 B.n20 163.367
R283 B.n22 B.n21 163.367
R284 B.n278 B.n22 163.367
R285 B.n278 B.n27 163.367
R286 B.n28 B.n27 163.367
R287 B.n29 B.n28 163.367
R288 B.n283 B.n29 163.367
R289 B.n283 B.n34 163.367
R290 B.n35 B.n34 163.367
R291 B.n152 B.n151 163.367
R292 B.n201 B.n151 163.367
R293 B.n199 B.n198 163.367
R294 B.n195 B.n194 163.367
R295 B.n191 B.n190 163.367
R296 B.n187 B.n186 163.367
R297 B.n183 B.n182 163.367
R298 B.n179 B.n178 163.367
R299 B.n175 B.n174 163.367
R300 B.n170 B.n169 163.367
R301 B.n166 B.n165 163.367
R302 B.n162 B.n161 163.367
R303 B.n158 B.n139 163.367
R304 B.n216 B.n135 163.367
R305 B.n216 B.n133 163.367
R306 B.n220 B.n133 163.367
R307 B.n220 B.n127 163.367
R308 B.n228 B.n127 163.367
R309 B.n228 B.n125 163.367
R310 B.n232 B.n125 163.367
R311 B.n232 B.n119 163.367
R312 B.n240 B.n119 163.367
R313 B.n240 B.n117 163.367
R314 B.n244 B.n117 163.367
R315 B.n244 B.n111 163.367
R316 B.n254 B.n111 163.367
R317 B.n254 B.n109 163.367
R318 B.n258 B.n109 163.367
R319 B.n258 B.n3 163.367
R320 B.n325 B.n3 163.367
R321 B.n321 B.n2 163.367
R322 B.n321 B.n320 163.367
R323 B.n320 B.n9 163.367
R324 B.n316 B.n9 163.367
R325 B.n316 B.n11 163.367
R326 B.n312 B.n11 163.367
R327 B.n312 B.n17 163.367
R328 B.n308 B.n17 163.367
R329 B.n308 B.n19 163.367
R330 B.n304 B.n19 163.367
R331 B.n304 B.n24 163.367
R332 B.n300 B.n24 163.367
R333 B.n300 B.n26 163.367
R334 B.n296 B.n26 163.367
R335 B.n296 B.n31 163.367
R336 B.n292 B.n31 163.367
R337 B.n292 B.n33 163.367
R338 B.n215 B.n136 121.331
R339 B.n215 B.n131 121.331
R340 B.n221 B.n131 121.331
R341 B.n221 B.n132 121.331
R342 B.n227 B.n124 121.331
R343 B.n233 B.n124 121.331
R344 B.n233 B.n120 121.331
R345 B.n239 B.n120 121.331
R346 B.n239 B.n116 121.331
R347 B.n245 B.n116 121.331
R348 B.n253 B.n112 121.331
R349 B.n253 B.n252 121.331
R350 B.n259 B.n4 121.331
R351 B.n324 B.n4 121.331
R352 B.n324 B.n323 121.331
R353 B.n323 B.n322 121.331
R354 B.n322 B.n8 121.331
R355 B.n315 B.n12 121.331
R356 B.n315 B.n314 121.331
R357 B.n313 B.n16 121.331
R358 B.n307 B.n16 121.331
R359 B.n307 B.n306 121.331
R360 B.n306 B.n305 121.331
R361 B.n305 B.n23 121.331
R362 B.n299 B.n23 121.331
R363 B.n298 B.n297 121.331
R364 B.n297 B.n30 121.331
R365 B.n291 B.n30 121.331
R366 B.n291 B.n290 121.331
R367 B.n132 B.t8 99.9194
R368 B.t1 B.n112 99.9194
R369 B.n314 B.t17 99.9194
R370 B.t4 B.n298 99.9194
R371 B.n259 B.t2 82.0767
R372 B.t0 B.n8 82.0767
R373 B.n55 B.n36 71.676
R374 B.n59 B.n37 71.676
R375 B.n63 B.n38 71.676
R376 B.n67 B.n39 71.676
R377 B.n71 B.n40 71.676
R378 B.n76 B.n41 71.676
R379 B.n80 B.n42 71.676
R380 B.n84 B.n43 71.676
R381 B.n88 B.n44 71.676
R382 B.n92 B.n45 71.676
R383 B.n96 B.n46 71.676
R384 B.n100 B.n47 71.676
R385 B.n104 B.n48 71.676
R386 B.n49 B.n48 71.676
R387 B.n103 B.n47 71.676
R388 B.n99 B.n46 71.676
R389 B.n95 B.n45 71.676
R390 B.n91 B.n44 71.676
R391 B.n87 B.n43 71.676
R392 B.n83 B.n42 71.676
R393 B.n79 B.n41 71.676
R394 B.n75 B.n40 71.676
R395 B.n70 B.n39 71.676
R396 B.n66 B.n38 71.676
R397 B.n62 B.n37 71.676
R398 B.n58 B.n36 71.676
R399 B.n207 B.n206 71.676
R400 B.n201 B.n140 71.676
R401 B.n198 B.n141 71.676
R402 B.n194 B.n142 71.676
R403 B.n190 B.n143 71.676
R404 B.n186 B.n144 71.676
R405 B.n182 B.n145 71.676
R406 B.n178 B.n146 71.676
R407 B.n174 B.n147 71.676
R408 B.n169 B.n148 71.676
R409 B.n165 B.n149 71.676
R410 B.n161 B.n150 71.676
R411 B.n209 B.n139 71.676
R412 B.n207 B.n152 71.676
R413 B.n199 B.n140 71.676
R414 B.n195 B.n141 71.676
R415 B.n191 B.n142 71.676
R416 B.n187 B.n143 71.676
R417 B.n183 B.n144 71.676
R418 B.n179 B.n145 71.676
R419 B.n175 B.n146 71.676
R420 B.n170 B.n147 71.676
R421 B.n166 B.n148 71.676
R422 B.n162 B.n149 71.676
R423 B.n158 B.n150 71.676
R424 B.n210 B.n209 71.676
R425 B.n326 B.n325 71.676
R426 B.n326 B.n2 71.676
R427 B.n73 B.n54 59.5399
R428 B.n52 B.n51 59.5399
R429 B.n172 B.n157 59.5399
R430 B.n155 B.n154 59.5399
R431 B.n252 B.t2 39.2544
R432 B.n12 B.t0 39.2544
R433 B.n205 B.n134 35.4346
R434 B.n212 B.n211 35.4346
R435 B.n287 B.n286 35.4346
R436 B.n56 B.n32 35.4346
R437 B.n227 B.t8 21.4117
R438 B.n245 B.t1 21.4117
R439 B.t17 B.n313 21.4117
R440 B.n299 B.t4 21.4117
R441 B.n54 B.n53 20.752
R442 B.n51 B.n50 20.752
R443 B.n157 B.n156 20.752
R444 B.n154 B.n153 20.752
R445 B B.n327 18.0485
R446 B.n217 B.n134 10.6151
R447 B.n218 B.n217 10.6151
R448 B.n219 B.n218 10.6151
R449 B.n219 B.n126 10.6151
R450 B.n229 B.n126 10.6151
R451 B.n230 B.n229 10.6151
R452 B.n231 B.n230 10.6151
R453 B.n231 B.n118 10.6151
R454 B.n241 B.n118 10.6151
R455 B.n242 B.n241 10.6151
R456 B.n243 B.n242 10.6151
R457 B.n243 B.n110 10.6151
R458 B.n255 B.n110 10.6151
R459 B.n256 B.n255 10.6151
R460 B.n257 B.n256 10.6151
R461 B.n257 B.n0 10.6151
R462 B.n205 B.n204 10.6151
R463 B.n204 B.n203 10.6151
R464 B.n203 B.n202 10.6151
R465 B.n202 B.n200 10.6151
R466 B.n200 B.n197 10.6151
R467 B.n197 B.n196 10.6151
R468 B.n196 B.n193 10.6151
R469 B.n193 B.n192 10.6151
R470 B.n189 B.n188 10.6151
R471 B.n188 B.n185 10.6151
R472 B.n185 B.n184 10.6151
R473 B.n184 B.n181 10.6151
R474 B.n181 B.n180 10.6151
R475 B.n180 B.n177 10.6151
R476 B.n177 B.n176 10.6151
R477 B.n176 B.n173 10.6151
R478 B.n171 B.n168 10.6151
R479 B.n168 B.n167 10.6151
R480 B.n167 B.n164 10.6151
R481 B.n164 B.n163 10.6151
R482 B.n163 B.n160 10.6151
R483 B.n160 B.n159 10.6151
R484 B.n159 B.n138 10.6151
R485 B.n211 B.n138 10.6151
R486 B.n213 B.n212 10.6151
R487 B.n213 B.n129 10.6151
R488 B.n223 B.n129 10.6151
R489 B.n224 B.n223 10.6151
R490 B.n225 B.n224 10.6151
R491 B.n225 B.n122 10.6151
R492 B.n235 B.n122 10.6151
R493 B.n236 B.n235 10.6151
R494 B.n237 B.n236 10.6151
R495 B.n237 B.n114 10.6151
R496 B.n247 B.n114 10.6151
R497 B.n248 B.n247 10.6151
R498 B.n250 B.n248 10.6151
R499 B.n250 B.n249 10.6151
R500 B.n249 B.n107 10.6151
R501 B.n262 B.n107 10.6151
R502 B.n263 B.n262 10.6151
R503 B.n264 B.n263 10.6151
R504 B.n265 B.n264 10.6151
R505 B.n266 B.n265 10.6151
R506 B.n269 B.n266 10.6151
R507 B.n270 B.n269 10.6151
R508 B.n271 B.n270 10.6151
R509 B.n272 B.n271 10.6151
R510 B.n274 B.n272 10.6151
R511 B.n275 B.n274 10.6151
R512 B.n276 B.n275 10.6151
R513 B.n277 B.n276 10.6151
R514 B.n279 B.n277 10.6151
R515 B.n280 B.n279 10.6151
R516 B.n281 B.n280 10.6151
R517 B.n282 B.n281 10.6151
R518 B.n284 B.n282 10.6151
R519 B.n285 B.n284 10.6151
R520 B.n286 B.n285 10.6151
R521 B.n319 B.n1 10.6151
R522 B.n319 B.n318 10.6151
R523 B.n318 B.n317 10.6151
R524 B.n317 B.n10 10.6151
R525 B.n311 B.n10 10.6151
R526 B.n311 B.n310 10.6151
R527 B.n310 B.n309 10.6151
R528 B.n309 B.n18 10.6151
R529 B.n303 B.n18 10.6151
R530 B.n303 B.n302 10.6151
R531 B.n302 B.n301 10.6151
R532 B.n301 B.n25 10.6151
R533 B.n295 B.n25 10.6151
R534 B.n295 B.n294 10.6151
R535 B.n294 B.n293 10.6151
R536 B.n293 B.n32 10.6151
R537 B.n57 B.n56 10.6151
R538 B.n60 B.n57 10.6151
R539 B.n61 B.n60 10.6151
R540 B.n64 B.n61 10.6151
R541 B.n65 B.n64 10.6151
R542 B.n68 B.n65 10.6151
R543 B.n69 B.n68 10.6151
R544 B.n72 B.n69 10.6151
R545 B.n77 B.n74 10.6151
R546 B.n78 B.n77 10.6151
R547 B.n81 B.n78 10.6151
R548 B.n82 B.n81 10.6151
R549 B.n85 B.n82 10.6151
R550 B.n86 B.n85 10.6151
R551 B.n89 B.n86 10.6151
R552 B.n90 B.n89 10.6151
R553 B.n94 B.n93 10.6151
R554 B.n97 B.n94 10.6151
R555 B.n98 B.n97 10.6151
R556 B.n101 B.n98 10.6151
R557 B.n102 B.n101 10.6151
R558 B.n105 B.n102 10.6151
R559 B.n106 B.n105 10.6151
R560 B.n287 B.n106 10.6151
R561 B.n327 B.n0 8.11757
R562 B.n327 B.n1 8.11757
R563 B.n189 B.n155 6.4005
R564 B.n173 B.n172 6.4005
R565 B.n74 B.n73 6.4005
R566 B.n90 B.n52 6.4005
R567 B.n192 B.n155 4.21513
R568 B.n172 B.n171 4.21513
R569 B.n73 B.n72 4.21513
R570 B.n93 B.n52 4.21513
R571 VN.n0 VN.t0 103.392
R572 VN.n1 VN.t3 103.392
R573 VN.n0 VN.t1 103.344
R574 VN.n1 VN.t2 103.344
R575 VN VN.n1 77.1867
R576 VN VN.n0 44.7132
R577 VDD2.n2 VDD2.n0 265.248
R578 VDD2.n2 VDD2.n1 238
R579 VDD2.n1 VDD2.t2 22.2477
R580 VDD2.n1 VDD2.t1 22.2477
R581 VDD2.n0 VDD2.t3 22.2477
R582 VDD2.n0 VDD2.t0 22.2477
R583 VDD2 VDD2.n2 0.0586897
R584 VTAIL.n6 VTAIL.t1 243.567
R585 VTAIL.n5 VTAIL.t0 243.567
R586 VTAIL.n4 VTAIL.t4 243.567
R587 VTAIL.n3 VTAIL.t5 243.567
R588 VTAIL.n7 VTAIL.t6 243.566
R589 VTAIL.n0 VTAIL.t7 243.566
R590 VTAIL.n1 VTAIL.t3 243.566
R591 VTAIL.n2 VTAIL.t2 243.566
R592 VTAIL.n7 VTAIL.n6 14.0565
R593 VTAIL.n3 VTAIL.n2 14.0565
R594 VTAIL.n4 VTAIL.n3 0.922914
R595 VTAIL.n6 VTAIL.n5 0.922914
R596 VTAIL.n2 VTAIL.n1 0.922914
R597 VTAIL VTAIL.n0 0.519897
R598 VTAIL.n5 VTAIL.n4 0.470328
R599 VTAIL.n1 VTAIL.n0 0.470328
R600 VTAIL VTAIL.n7 0.403517
R601 VP.n6 VP.n5 161.3
R602 VP.n4 VP.n0 161.3
R603 VP.n3 VP.n2 161.3
R604 VP.n1 VP.t1 103.392
R605 VP.n1 VP.t3 103.344
R606 VP.n3 VP.t2 82.3964
R607 VP.n5 VP.t0 82.3964
R608 VP.n2 VP.n1 76.806
R609 VP.n4 VP.n3 24.1005
R610 VP.n5 VP.n4 24.1005
R611 VP.n2 VP.n0 0.189894
R612 VP.n6 VP.n0 0.189894
R613 VP VP.n6 0.0516364
R614 VDD1 VDD1.n1 265.772
R615 VDD1 VDD1.n0 238.058
R616 VDD1.n0 VDD1.t2 22.2477
R617 VDD1.n0 VDD1.t0 22.2477
R618 VDD1.n1 VDD1.t1 22.2477
R619 VDD1.n1 VDD1.t3 22.2477
C0 VDD1 VDD2 0.576103f
C1 VDD2 VP 0.284075f
C2 VDD1 VN 0.154314f
C3 VP VN 2.8034f
C4 VTAIL VDD2 1.9137f
C5 VTAIL VN 0.728544f
C6 VDD1 VP 0.645296f
C7 VTAIL VDD1 1.87197f
C8 VTAIL VP 0.742651f
C9 VDD2 VN 0.51696f
C10 VDD2 B 1.75364f
C11 VDD1 B 1.91424f
C12 VTAIL B 2.18283f
C13 VN B 5.82108f
C14 VP B 4.041274f
C15 VP.n0 B 0.037543f
C16 VP.t3 B 0.103665f
C17 VP.t1 B 0.103731f
C18 VP.n1 B 0.575886f
C19 VP.n2 B 1.58019f
C20 VP.t2 B 0.085384f
C21 VP.n3 B 0.087489f
C22 VP.n4 B 0.008519f
C23 VP.t0 B 0.085384f
C24 VP.n5 B 0.087489f
C25 VP.n6 B 0.029094f
C26 VN.t0 B 0.101812f
C27 VN.t1 B 0.101747f
C28 VN.n0 B 0.144531f
C29 VN.t3 B 0.101812f
C30 VN.t2 B 0.101747f
C31 VN.n1 B 0.578506f
.ends

