* NGSPICE file created from diff_pair_sample_1257.ext - technology: sky130A

.subckt diff_pair_sample_1257 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=4.407 ps=23.38 w=11.3 l=0.35
X1 VTAIL.t13 VP.t1 VDD1.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X2 VDD1.t7 VP.t2 VTAIL.t12 B.t23 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X3 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=0 ps=0 w=11.3 l=0.35
X4 VDD2.t9 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=1.8645 ps=11.63 w=11.3 l=0.35
X5 VDD1.t6 VP.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=4.407 ps=23.38 w=11.3 l=0.35
X6 VTAIL.t9 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X7 VTAIL.t2 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X8 VDD2.t7 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=4.407 ps=23.38 w=11.3 l=0.35
X9 VTAIL.t4 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X10 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=0 ps=0 w=11.3 l=0.35
X11 VDD2.t5 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=4.407 ps=23.38 w=11.3 l=0.35
X12 VTAIL.t1 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X13 VDD1.t4 VP.t5 VTAIL.t10 B.t22 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=1.8645 ps=11.63 w=11.3 l=0.35
X14 VTAIL.t8 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X15 VTAIL.t5 VN.t6 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X16 VDD2.t2 VN.t7 VTAIL.t17 B.t22 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=1.8645 ps=11.63 w=11.3 l=0.35
X17 VDD2.t1 VN.t8 VTAIL.t18 B.t23 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X18 VDD2.t0 VN.t9 VTAIL.t19 B.t21 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X19 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=0 ps=0 w=11.3 l=0.35
X20 VDD1.t2 VP.t7 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X21 VTAIL.t7 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8645 pd=11.63 as=1.8645 ps=11.63 w=11.3 l=0.35
X22 VDD1.t0 VP.t9 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=1.8645 ps=11.63 w=11.3 l=0.35
X23 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.407 pd=23.38 as=0 ps=0 w=11.3 l=0.35
R0 VP.n21 VP.t3 918.721
R1 VP.n14 VP.t5 918.721
R2 VP.n11 VP.t0 918.721
R3 VP.n5 VP.t9 918.721
R4 VP.n13 VP.t4 891.701
R5 VP.n18 VP.t2 891.701
R6 VP.n20 VP.t6 891.701
R7 VP.n10 VP.t1 891.701
R8 VP.n8 VP.t7 891.701
R9 VP.n4 VP.t8 891.701
R10 VP.n6 VP.n5 161.489
R11 VP.n22 VP.n21 161.3
R12 VP.n7 VP.n6 161.3
R13 VP.n8 VP.n3 161.3
R14 VP.n9 VP.n2 161.3
R15 VP.n12 VP.n11 161.3
R16 VP.n19 VP.n0 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n1 161.3
R19 VP.n15 VP.n14 161.3
R20 VP.n18 VP.n1 47.4702
R21 VP.n19 VP.n18 47.4702
R22 VP.n9 VP.n8 47.4702
R23 VP.n8 VP.n7 47.4702
R24 VP.n15 VP.n12 40.4929
R25 VP.n14 VP.n13 21.1793
R26 VP.n21 VP.n20 21.1793
R27 VP.n11 VP.n10 21.1793
R28 VP.n5 VP.n4 21.1793
R29 VP.n13 VP.n1 0.730803
R30 VP.n20 VP.n19 0.730803
R31 VP.n10 VP.n9 0.730803
R32 VP.n7 VP.n4 0.730803
R33 VP.n6 VP.n3 0.189894
R34 VP.n3 VP.n2 0.189894
R35 VP.n12 VP.n2 0.189894
R36 VP.n16 VP.n15 0.189894
R37 VP.n17 VP.n16 0.189894
R38 VP.n17 VP.n0 0.189894
R39 VP.n22 VP.n0 0.189894
R40 VP VP.n22 0.0516364
R41 VTAIL.n256 VTAIL.n200 289.615
R42 VTAIL.n58 VTAIL.n2 289.615
R43 VTAIL.n194 VTAIL.n138 289.615
R44 VTAIL.n128 VTAIL.n72 289.615
R45 VTAIL.n221 VTAIL.n220 185
R46 VTAIL.n223 VTAIL.n222 185
R47 VTAIL.n216 VTAIL.n215 185
R48 VTAIL.n229 VTAIL.n228 185
R49 VTAIL.n231 VTAIL.n230 185
R50 VTAIL.n212 VTAIL.n211 185
R51 VTAIL.n238 VTAIL.n237 185
R52 VTAIL.n239 VTAIL.n210 185
R53 VTAIL.n241 VTAIL.n240 185
R54 VTAIL.n208 VTAIL.n207 185
R55 VTAIL.n247 VTAIL.n246 185
R56 VTAIL.n249 VTAIL.n248 185
R57 VTAIL.n204 VTAIL.n203 185
R58 VTAIL.n255 VTAIL.n254 185
R59 VTAIL.n257 VTAIL.n256 185
R60 VTAIL.n23 VTAIL.n22 185
R61 VTAIL.n25 VTAIL.n24 185
R62 VTAIL.n18 VTAIL.n17 185
R63 VTAIL.n31 VTAIL.n30 185
R64 VTAIL.n33 VTAIL.n32 185
R65 VTAIL.n14 VTAIL.n13 185
R66 VTAIL.n40 VTAIL.n39 185
R67 VTAIL.n41 VTAIL.n12 185
R68 VTAIL.n43 VTAIL.n42 185
R69 VTAIL.n10 VTAIL.n9 185
R70 VTAIL.n49 VTAIL.n48 185
R71 VTAIL.n51 VTAIL.n50 185
R72 VTAIL.n6 VTAIL.n5 185
R73 VTAIL.n57 VTAIL.n56 185
R74 VTAIL.n59 VTAIL.n58 185
R75 VTAIL.n195 VTAIL.n194 185
R76 VTAIL.n193 VTAIL.n192 185
R77 VTAIL.n142 VTAIL.n141 185
R78 VTAIL.n187 VTAIL.n186 185
R79 VTAIL.n185 VTAIL.n184 185
R80 VTAIL.n146 VTAIL.n145 185
R81 VTAIL.n150 VTAIL.n148 185
R82 VTAIL.n179 VTAIL.n178 185
R83 VTAIL.n177 VTAIL.n176 185
R84 VTAIL.n152 VTAIL.n151 185
R85 VTAIL.n171 VTAIL.n170 185
R86 VTAIL.n169 VTAIL.n168 185
R87 VTAIL.n156 VTAIL.n155 185
R88 VTAIL.n163 VTAIL.n162 185
R89 VTAIL.n161 VTAIL.n160 185
R90 VTAIL.n129 VTAIL.n128 185
R91 VTAIL.n127 VTAIL.n126 185
R92 VTAIL.n76 VTAIL.n75 185
R93 VTAIL.n121 VTAIL.n120 185
R94 VTAIL.n119 VTAIL.n118 185
R95 VTAIL.n80 VTAIL.n79 185
R96 VTAIL.n84 VTAIL.n82 185
R97 VTAIL.n113 VTAIL.n112 185
R98 VTAIL.n111 VTAIL.n110 185
R99 VTAIL.n86 VTAIL.n85 185
R100 VTAIL.n105 VTAIL.n104 185
R101 VTAIL.n103 VTAIL.n102 185
R102 VTAIL.n90 VTAIL.n89 185
R103 VTAIL.n97 VTAIL.n96 185
R104 VTAIL.n95 VTAIL.n94 185
R105 VTAIL.n219 VTAIL.t0 149.524
R106 VTAIL.n21 VTAIL.t11 149.524
R107 VTAIL.n159 VTAIL.t14 149.524
R108 VTAIL.n93 VTAIL.t3 149.524
R109 VTAIL.n222 VTAIL.n221 104.615
R110 VTAIL.n222 VTAIL.n215 104.615
R111 VTAIL.n229 VTAIL.n215 104.615
R112 VTAIL.n230 VTAIL.n229 104.615
R113 VTAIL.n230 VTAIL.n211 104.615
R114 VTAIL.n238 VTAIL.n211 104.615
R115 VTAIL.n239 VTAIL.n238 104.615
R116 VTAIL.n240 VTAIL.n239 104.615
R117 VTAIL.n240 VTAIL.n207 104.615
R118 VTAIL.n247 VTAIL.n207 104.615
R119 VTAIL.n248 VTAIL.n247 104.615
R120 VTAIL.n248 VTAIL.n203 104.615
R121 VTAIL.n255 VTAIL.n203 104.615
R122 VTAIL.n256 VTAIL.n255 104.615
R123 VTAIL.n24 VTAIL.n23 104.615
R124 VTAIL.n24 VTAIL.n17 104.615
R125 VTAIL.n31 VTAIL.n17 104.615
R126 VTAIL.n32 VTAIL.n31 104.615
R127 VTAIL.n32 VTAIL.n13 104.615
R128 VTAIL.n40 VTAIL.n13 104.615
R129 VTAIL.n41 VTAIL.n40 104.615
R130 VTAIL.n42 VTAIL.n41 104.615
R131 VTAIL.n42 VTAIL.n9 104.615
R132 VTAIL.n49 VTAIL.n9 104.615
R133 VTAIL.n50 VTAIL.n49 104.615
R134 VTAIL.n50 VTAIL.n5 104.615
R135 VTAIL.n57 VTAIL.n5 104.615
R136 VTAIL.n58 VTAIL.n57 104.615
R137 VTAIL.n194 VTAIL.n193 104.615
R138 VTAIL.n193 VTAIL.n141 104.615
R139 VTAIL.n186 VTAIL.n141 104.615
R140 VTAIL.n186 VTAIL.n185 104.615
R141 VTAIL.n185 VTAIL.n145 104.615
R142 VTAIL.n150 VTAIL.n145 104.615
R143 VTAIL.n178 VTAIL.n150 104.615
R144 VTAIL.n178 VTAIL.n177 104.615
R145 VTAIL.n177 VTAIL.n151 104.615
R146 VTAIL.n170 VTAIL.n151 104.615
R147 VTAIL.n170 VTAIL.n169 104.615
R148 VTAIL.n169 VTAIL.n155 104.615
R149 VTAIL.n162 VTAIL.n155 104.615
R150 VTAIL.n162 VTAIL.n161 104.615
R151 VTAIL.n128 VTAIL.n127 104.615
R152 VTAIL.n127 VTAIL.n75 104.615
R153 VTAIL.n120 VTAIL.n75 104.615
R154 VTAIL.n120 VTAIL.n119 104.615
R155 VTAIL.n119 VTAIL.n79 104.615
R156 VTAIL.n84 VTAIL.n79 104.615
R157 VTAIL.n112 VTAIL.n84 104.615
R158 VTAIL.n112 VTAIL.n111 104.615
R159 VTAIL.n111 VTAIL.n85 104.615
R160 VTAIL.n104 VTAIL.n85 104.615
R161 VTAIL.n104 VTAIL.n103 104.615
R162 VTAIL.n103 VTAIL.n89 104.615
R163 VTAIL.n96 VTAIL.n89 104.615
R164 VTAIL.n96 VTAIL.n95 104.615
R165 VTAIL.n221 VTAIL.t0 52.3082
R166 VTAIL.n23 VTAIL.t11 52.3082
R167 VTAIL.n161 VTAIL.t14 52.3082
R168 VTAIL.n95 VTAIL.t3 52.3082
R169 VTAIL.n137 VTAIL.n136 43.4717
R170 VTAIL.n135 VTAIL.n134 43.4717
R171 VTAIL.n71 VTAIL.n70 43.4717
R172 VTAIL.n69 VTAIL.n68 43.4717
R173 VTAIL.n263 VTAIL.n262 43.4715
R174 VTAIL.n1 VTAIL.n0 43.4715
R175 VTAIL.n65 VTAIL.n64 43.4715
R176 VTAIL.n67 VTAIL.n66 43.4715
R177 VTAIL.n261 VTAIL.n260 30.246
R178 VTAIL.n63 VTAIL.n62 30.246
R179 VTAIL.n199 VTAIL.n198 30.246
R180 VTAIL.n133 VTAIL.n132 30.246
R181 VTAIL.n69 VTAIL.n67 23.2807
R182 VTAIL.n261 VTAIL.n199 22.6945
R183 VTAIL.n241 VTAIL.n208 13.1884
R184 VTAIL.n43 VTAIL.n10 13.1884
R185 VTAIL.n148 VTAIL.n146 13.1884
R186 VTAIL.n82 VTAIL.n80 13.1884
R187 VTAIL.n242 VTAIL.n210 12.8005
R188 VTAIL.n246 VTAIL.n245 12.8005
R189 VTAIL.n44 VTAIL.n12 12.8005
R190 VTAIL.n48 VTAIL.n47 12.8005
R191 VTAIL.n184 VTAIL.n183 12.8005
R192 VTAIL.n180 VTAIL.n179 12.8005
R193 VTAIL.n118 VTAIL.n117 12.8005
R194 VTAIL.n114 VTAIL.n113 12.8005
R195 VTAIL.n237 VTAIL.n236 12.0247
R196 VTAIL.n249 VTAIL.n206 12.0247
R197 VTAIL.n39 VTAIL.n38 12.0247
R198 VTAIL.n51 VTAIL.n8 12.0247
R199 VTAIL.n187 VTAIL.n144 12.0247
R200 VTAIL.n176 VTAIL.n149 12.0247
R201 VTAIL.n121 VTAIL.n78 12.0247
R202 VTAIL.n110 VTAIL.n83 12.0247
R203 VTAIL.n235 VTAIL.n212 11.249
R204 VTAIL.n250 VTAIL.n204 11.249
R205 VTAIL.n37 VTAIL.n14 11.249
R206 VTAIL.n52 VTAIL.n6 11.249
R207 VTAIL.n188 VTAIL.n142 11.249
R208 VTAIL.n175 VTAIL.n152 11.249
R209 VTAIL.n122 VTAIL.n76 11.249
R210 VTAIL.n109 VTAIL.n86 11.249
R211 VTAIL.n232 VTAIL.n231 10.4732
R212 VTAIL.n254 VTAIL.n253 10.4732
R213 VTAIL.n34 VTAIL.n33 10.4732
R214 VTAIL.n56 VTAIL.n55 10.4732
R215 VTAIL.n192 VTAIL.n191 10.4732
R216 VTAIL.n172 VTAIL.n171 10.4732
R217 VTAIL.n126 VTAIL.n125 10.4732
R218 VTAIL.n106 VTAIL.n105 10.4732
R219 VTAIL.n220 VTAIL.n219 10.2747
R220 VTAIL.n22 VTAIL.n21 10.2747
R221 VTAIL.n160 VTAIL.n159 10.2747
R222 VTAIL.n94 VTAIL.n93 10.2747
R223 VTAIL.n228 VTAIL.n214 9.69747
R224 VTAIL.n257 VTAIL.n202 9.69747
R225 VTAIL.n30 VTAIL.n16 9.69747
R226 VTAIL.n59 VTAIL.n4 9.69747
R227 VTAIL.n195 VTAIL.n140 9.69747
R228 VTAIL.n168 VTAIL.n154 9.69747
R229 VTAIL.n129 VTAIL.n74 9.69747
R230 VTAIL.n102 VTAIL.n88 9.69747
R231 VTAIL.n260 VTAIL.n259 9.45567
R232 VTAIL.n62 VTAIL.n61 9.45567
R233 VTAIL.n198 VTAIL.n197 9.45567
R234 VTAIL.n132 VTAIL.n131 9.45567
R235 VTAIL.n259 VTAIL.n258 9.3005
R236 VTAIL.n202 VTAIL.n201 9.3005
R237 VTAIL.n253 VTAIL.n252 9.3005
R238 VTAIL.n251 VTAIL.n250 9.3005
R239 VTAIL.n206 VTAIL.n205 9.3005
R240 VTAIL.n245 VTAIL.n244 9.3005
R241 VTAIL.n218 VTAIL.n217 9.3005
R242 VTAIL.n225 VTAIL.n224 9.3005
R243 VTAIL.n227 VTAIL.n226 9.3005
R244 VTAIL.n214 VTAIL.n213 9.3005
R245 VTAIL.n233 VTAIL.n232 9.3005
R246 VTAIL.n235 VTAIL.n234 9.3005
R247 VTAIL.n236 VTAIL.n209 9.3005
R248 VTAIL.n243 VTAIL.n242 9.3005
R249 VTAIL.n61 VTAIL.n60 9.3005
R250 VTAIL.n4 VTAIL.n3 9.3005
R251 VTAIL.n55 VTAIL.n54 9.3005
R252 VTAIL.n53 VTAIL.n52 9.3005
R253 VTAIL.n8 VTAIL.n7 9.3005
R254 VTAIL.n47 VTAIL.n46 9.3005
R255 VTAIL.n20 VTAIL.n19 9.3005
R256 VTAIL.n27 VTAIL.n26 9.3005
R257 VTAIL.n29 VTAIL.n28 9.3005
R258 VTAIL.n16 VTAIL.n15 9.3005
R259 VTAIL.n35 VTAIL.n34 9.3005
R260 VTAIL.n37 VTAIL.n36 9.3005
R261 VTAIL.n38 VTAIL.n11 9.3005
R262 VTAIL.n45 VTAIL.n44 9.3005
R263 VTAIL.n158 VTAIL.n157 9.3005
R264 VTAIL.n165 VTAIL.n164 9.3005
R265 VTAIL.n167 VTAIL.n166 9.3005
R266 VTAIL.n154 VTAIL.n153 9.3005
R267 VTAIL.n173 VTAIL.n172 9.3005
R268 VTAIL.n175 VTAIL.n174 9.3005
R269 VTAIL.n149 VTAIL.n147 9.3005
R270 VTAIL.n181 VTAIL.n180 9.3005
R271 VTAIL.n197 VTAIL.n196 9.3005
R272 VTAIL.n140 VTAIL.n139 9.3005
R273 VTAIL.n191 VTAIL.n190 9.3005
R274 VTAIL.n189 VTAIL.n188 9.3005
R275 VTAIL.n144 VTAIL.n143 9.3005
R276 VTAIL.n183 VTAIL.n182 9.3005
R277 VTAIL.n92 VTAIL.n91 9.3005
R278 VTAIL.n99 VTAIL.n98 9.3005
R279 VTAIL.n101 VTAIL.n100 9.3005
R280 VTAIL.n88 VTAIL.n87 9.3005
R281 VTAIL.n107 VTAIL.n106 9.3005
R282 VTAIL.n109 VTAIL.n108 9.3005
R283 VTAIL.n83 VTAIL.n81 9.3005
R284 VTAIL.n115 VTAIL.n114 9.3005
R285 VTAIL.n131 VTAIL.n130 9.3005
R286 VTAIL.n74 VTAIL.n73 9.3005
R287 VTAIL.n125 VTAIL.n124 9.3005
R288 VTAIL.n123 VTAIL.n122 9.3005
R289 VTAIL.n78 VTAIL.n77 9.3005
R290 VTAIL.n117 VTAIL.n116 9.3005
R291 VTAIL.n227 VTAIL.n216 8.92171
R292 VTAIL.n258 VTAIL.n200 8.92171
R293 VTAIL.n29 VTAIL.n18 8.92171
R294 VTAIL.n60 VTAIL.n2 8.92171
R295 VTAIL.n196 VTAIL.n138 8.92171
R296 VTAIL.n167 VTAIL.n156 8.92171
R297 VTAIL.n130 VTAIL.n72 8.92171
R298 VTAIL.n101 VTAIL.n90 8.92171
R299 VTAIL.n224 VTAIL.n223 8.14595
R300 VTAIL.n26 VTAIL.n25 8.14595
R301 VTAIL.n164 VTAIL.n163 8.14595
R302 VTAIL.n98 VTAIL.n97 8.14595
R303 VTAIL.n220 VTAIL.n218 7.3702
R304 VTAIL.n22 VTAIL.n20 7.3702
R305 VTAIL.n160 VTAIL.n158 7.3702
R306 VTAIL.n94 VTAIL.n92 7.3702
R307 VTAIL.n223 VTAIL.n218 5.81868
R308 VTAIL.n25 VTAIL.n20 5.81868
R309 VTAIL.n163 VTAIL.n158 5.81868
R310 VTAIL.n97 VTAIL.n92 5.81868
R311 VTAIL.n224 VTAIL.n216 5.04292
R312 VTAIL.n260 VTAIL.n200 5.04292
R313 VTAIL.n26 VTAIL.n18 5.04292
R314 VTAIL.n62 VTAIL.n2 5.04292
R315 VTAIL.n198 VTAIL.n138 5.04292
R316 VTAIL.n164 VTAIL.n156 5.04292
R317 VTAIL.n132 VTAIL.n72 5.04292
R318 VTAIL.n98 VTAIL.n90 5.04292
R319 VTAIL.n228 VTAIL.n227 4.26717
R320 VTAIL.n258 VTAIL.n257 4.26717
R321 VTAIL.n30 VTAIL.n29 4.26717
R322 VTAIL.n60 VTAIL.n59 4.26717
R323 VTAIL.n196 VTAIL.n195 4.26717
R324 VTAIL.n168 VTAIL.n167 4.26717
R325 VTAIL.n130 VTAIL.n129 4.26717
R326 VTAIL.n102 VTAIL.n101 4.26717
R327 VTAIL.n231 VTAIL.n214 3.49141
R328 VTAIL.n254 VTAIL.n202 3.49141
R329 VTAIL.n33 VTAIL.n16 3.49141
R330 VTAIL.n56 VTAIL.n4 3.49141
R331 VTAIL.n192 VTAIL.n140 3.49141
R332 VTAIL.n171 VTAIL.n154 3.49141
R333 VTAIL.n126 VTAIL.n74 3.49141
R334 VTAIL.n105 VTAIL.n88 3.49141
R335 VTAIL.n219 VTAIL.n217 2.84303
R336 VTAIL.n21 VTAIL.n19 2.84303
R337 VTAIL.n159 VTAIL.n157 2.84303
R338 VTAIL.n93 VTAIL.n91 2.84303
R339 VTAIL.n232 VTAIL.n212 2.71565
R340 VTAIL.n253 VTAIL.n204 2.71565
R341 VTAIL.n34 VTAIL.n14 2.71565
R342 VTAIL.n55 VTAIL.n6 2.71565
R343 VTAIL.n191 VTAIL.n142 2.71565
R344 VTAIL.n172 VTAIL.n152 2.71565
R345 VTAIL.n125 VTAIL.n76 2.71565
R346 VTAIL.n106 VTAIL.n86 2.71565
R347 VTAIL.n237 VTAIL.n235 1.93989
R348 VTAIL.n250 VTAIL.n249 1.93989
R349 VTAIL.n39 VTAIL.n37 1.93989
R350 VTAIL.n52 VTAIL.n51 1.93989
R351 VTAIL.n188 VTAIL.n187 1.93989
R352 VTAIL.n176 VTAIL.n175 1.93989
R353 VTAIL.n122 VTAIL.n121 1.93989
R354 VTAIL.n110 VTAIL.n109 1.93989
R355 VTAIL.n262 VTAIL.t19 1.75271
R356 VTAIL.n262 VTAIL.t2 1.75271
R357 VTAIL.n0 VTAIL.t6 1.75271
R358 VTAIL.n0 VTAIL.t1 1.75271
R359 VTAIL.n64 VTAIL.t12 1.75271
R360 VTAIL.n64 VTAIL.t8 1.75271
R361 VTAIL.n66 VTAIL.t10 1.75271
R362 VTAIL.n66 VTAIL.t9 1.75271
R363 VTAIL.n136 VTAIL.t15 1.75271
R364 VTAIL.n136 VTAIL.t13 1.75271
R365 VTAIL.n134 VTAIL.t16 1.75271
R366 VTAIL.n134 VTAIL.t7 1.75271
R367 VTAIL.n70 VTAIL.t18 1.75271
R368 VTAIL.n70 VTAIL.t4 1.75271
R369 VTAIL.n68 VTAIL.t17 1.75271
R370 VTAIL.n68 VTAIL.t5 1.75271
R371 VTAIL.n236 VTAIL.n210 1.16414
R372 VTAIL.n246 VTAIL.n206 1.16414
R373 VTAIL.n38 VTAIL.n12 1.16414
R374 VTAIL.n48 VTAIL.n8 1.16414
R375 VTAIL.n184 VTAIL.n144 1.16414
R376 VTAIL.n179 VTAIL.n149 1.16414
R377 VTAIL.n118 VTAIL.n78 1.16414
R378 VTAIL.n113 VTAIL.n83 1.16414
R379 VTAIL.n135 VTAIL.n133 0.763431
R380 VTAIL.n63 VTAIL.n1 0.763431
R381 VTAIL.n71 VTAIL.n69 0.586707
R382 VTAIL.n133 VTAIL.n71 0.586707
R383 VTAIL.n137 VTAIL.n135 0.586707
R384 VTAIL.n199 VTAIL.n137 0.586707
R385 VTAIL.n67 VTAIL.n65 0.586707
R386 VTAIL.n65 VTAIL.n63 0.586707
R387 VTAIL.n263 VTAIL.n261 0.586707
R388 VTAIL VTAIL.n1 0.498345
R389 VTAIL.n242 VTAIL.n241 0.388379
R390 VTAIL.n245 VTAIL.n208 0.388379
R391 VTAIL.n44 VTAIL.n43 0.388379
R392 VTAIL.n47 VTAIL.n10 0.388379
R393 VTAIL.n183 VTAIL.n146 0.388379
R394 VTAIL.n180 VTAIL.n148 0.388379
R395 VTAIL.n117 VTAIL.n80 0.388379
R396 VTAIL.n114 VTAIL.n82 0.388379
R397 VTAIL.n225 VTAIL.n217 0.155672
R398 VTAIL.n226 VTAIL.n225 0.155672
R399 VTAIL.n226 VTAIL.n213 0.155672
R400 VTAIL.n233 VTAIL.n213 0.155672
R401 VTAIL.n234 VTAIL.n233 0.155672
R402 VTAIL.n234 VTAIL.n209 0.155672
R403 VTAIL.n243 VTAIL.n209 0.155672
R404 VTAIL.n244 VTAIL.n243 0.155672
R405 VTAIL.n244 VTAIL.n205 0.155672
R406 VTAIL.n251 VTAIL.n205 0.155672
R407 VTAIL.n252 VTAIL.n251 0.155672
R408 VTAIL.n252 VTAIL.n201 0.155672
R409 VTAIL.n259 VTAIL.n201 0.155672
R410 VTAIL.n27 VTAIL.n19 0.155672
R411 VTAIL.n28 VTAIL.n27 0.155672
R412 VTAIL.n28 VTAIL.n15 0.155672
R413 VTAIL.n35 VTAIL.n15 0.155672
R414 VTAIL.n36 VTAIL.n35 0.155672
R415 VTAIL.n36 VTAIL.n11 0.155672
R416 VTAIL.n45 VTAIL.n11 0.155672
R417 VTAIL.n46 VTAIL.n45 0.155672
R418 VTAIL.n46 VTAIL.n7 0.155672
R419 VTAIL.n53 VTAIL.n7 0.155672
R420 VTAIL.n54 VTAIL.n53 0.155672
R421 VTAIL.n54 VTAIL.n3 0.155672
R422 VTAIL.n61 VTAIL.n3 0.155672
R423 VTAIL.n197 VTAIL.n139 0.155672
R424 VTAIL.n190 VTAIL.n139 0.155672
R425 VTAIL.n190 VTAIL.n189 0.155672
R426 VTAIL.n189 VTAIL.n143 0.155672
R427 VTAIL.n182 VTAIL.n143 0.155672
R428 VTAIL.n182 VTAIL.n181 0.155672
R429 VTAIL.n181 VTAIL.n147 0.155672
R430 VTAIL.n174 VTAIL.n147 0.155672
R431 VTAIL.n174 VTAIL.n173 0.155672
R432 VTAIL.n173 VTAIL.n153 0.155672
R433 VTAIL.n166 VTAIL.n153 0.155672
R434 VTAIL.n166 VTAIL.n165 0.155672
R435 VTAIL.n165 VTAIL.n157 0.155672
R436 VTAIL.n131 VTAIL.n73 0.155672
R437 VTAIL.n124 VTAIL.n73 0.155672
R438 VTAIL.n124 VTAIL.n123 0.155672
R439 VTAIL.n123 VTAIL.n77 0.155672
R440 VTAIL.n116 VTAIL.n77 0.155672
R441 VTAIL.n116 VTAIL.n115 0.155672
R442 VTAIL.n115 VTAIL.n81 0.155672
R443 VTAIL.n108 VTAIL.n81 0.155672
R444 VTAIL.n108 VTAIL.n107 0.155672
R445 VTAIL.n107 VTAIL.n87 0.155672
R446 VTAIL.n100 VTAIL.n87 0.155672
R447 VTAIL.n100 VTAIL.n99 0.155672
R448 VTAIL.n99 VTAIL.n91 0.155672
R449 VTAIL VTAIL.n263 0.0888621
R450 VDD1.n56 VDD1.n0 289.615
R451 VDD1.n119 VDD1.n63 289.615
R452 VDD1.n57 VDD1.n56 185
R453 VDD1.n55 VDD1.n54 185
R454 VDD1.n4 VDD1.n3 185
R455 VDD1.n49 VDD1.n48 185
R456 VDD1.n47 VDD1.n46 185
R457 VDD1.n8 VDD1.n7 185
R458 VDD1.n12 VDD1.n10 185
R459 VDD1.n41 VDD1.n40 185
R460 VDD1.n39 VDD1.n38 185
R461 VDD1.n14 VDD1.n13 185
R462 VDD1.n33 VDD1.n32 185
R463 VDD1.n31 VDD1.n30 185
R464 VDD1.n18 VDD1.n17 185
R465 VDD1.n25 VDD1.n24 185
R466 VDD1.n23 VDD1.n22 185
R467 VDD1.n84 VDD1.n83 185
R468 VDD1.n86 VDD1.n85 185
R469 VDD1.n79 VDD1.n78 185
R470 VDD1.n92 VDD1.n91 185
R471 VDD1.n94 VDD1.n93 185
R472 VDD1.n75 VDD1.n74 185
R473 VDD1.n101 VDD1.n100 185
R474 VDD1.n102 VDD1.n73 185
R475 VDD1.n104 VDD1.n103 185
R476 VDD1.n71 VDD1.n70 185
R477 VDD1.n110 VDD1.n109 185
R478 VDD1.n112 VDD1.n111 185
R479 VDD1.n67 VDD1.n66 185
R480 VDD1.n118 VDD1.n117 185
R481 VDD1.n120 VDD1.n119 185
R482 VDD1.n21 VDD1.t0 149.524
R483 VDD1.n82 VDD1.t4 149.524
R484 VDD1.n56 VDD1.n55 104.615
R485 VDD1.n55 VDD1.n3 104.615
R486 VDD1.n48 VDD1.n3 104.615
R487 VDD1.n48 VDD1.n47 104.615
R488 VDD1.n47 VDD1.n7 104.615
R489 VDD1.n12 VDD1.n7 104.615
R490 VDD1.n40 VDD1.n12 104.615
R491 VDD1.n40 VDD1.n39 104.615
R492 VDD1.n39 VDD1.n13 104.615
R493 VDD1.n32 VDD1.n13 104.615
R494 VDD1.n32 VDD1.n31 104.615
R495 VDD1.n31 VDD1.n17 104.615
R496 VDD1.n24 VDD1.n17 104.615
R497 VDD1.n24 VDD1.n23 104.615
R498 VDD1.n85 VDD1.n84 104.615
R499 VDD1.n85 VDD1.n78 104.615
R500 VDD1.n92 VDD1.n78 104.615
R501 VDD1.n93 VDD1.n92 104.615
R502 VDD1.n93 VDD1.n74 104.615
R503 VDD1.n101 VDD1.n74 104.615
R504 VDD1.n102 VDD1.n101 104.615
R505 VDD1.n103 VDD1.n102 104.615
R506 VDD1.n103 VDD1.n70 104.615
R507 VDD1.n110 VDD1.n70 104.615
R508 VDD1.n111 VDD1.n110 104.615
R509 VDD1.n111 VDD1.n66 104.615
R510 VDD1.n118 VDD1.n66 104.615
R511 VDD1.n119 VDD1.n118 104.615
R512 VDD1.n127 VDD1.n126 60.5346
R513 VDD1.n62 VDD1.n61 60.1505
R514 VDD1.n129 VDD1.n128 60.1503
R515 VDD1.n125 VDD1.n124 60.1503
R516 VDD1.n23 VDD1.t0 52.3082
R517 VDD1.n84 VDD1.t4 52.3082
R518 VDD1.n62 VDD1.n60 47.5109
R519 VDD1.n125 VDD1.n123 47.5109
R520 VDD1.n129 VDD1.n127 37.1173
R521 VDD1.n10 VDD1.n8 13.1884
R522 VDD1.n104 VDD1.n71 13.1884
R523 VDD1.n46 VDD1.n45 12.8005
R524 VDD1.n42 VDD1.n41 12.8005
R525 VDD1.n105 VDD1.n73 12.8005
R526 VDD1.n109 VDD1.n108 12.8005
R527 VDD1.n49 VDD1.n6 12.0247
R528 VDD1.n38 VDD1.n11 12.0247
R529 VDD1.n100 VDD1.n99 12.0247
R530 VDD1.n112 VDD1.n69 12.0247
R531 VDD1.n50 VDD1.n4 11.249
R532 VDD1.n37 VDD1.n14 11.249
R533 VDD1.n98 VDD1.n75 11.249
R534 VDD1.n113 VDD1.n67 11.249
R535 VDD1.n54 VDD1.n53 10.4732
R536 VDD1.n34 VDD1.n33 10.4732
R537 VDD1.n95 VDD1.n94 10.4732
R538 VDD1.n117 VDD1.n116 10.4732
R539 VDD1.n22 VDD1.n21 10.2747
R540 VDD1.n83 VDD1.n82 10.2747
R541 VDD1.n57 VDD1.n2 9.69747
R542 VDD1.n30 VDD1.n16 9.69747
R543 VDD1.n91 VDD1.n77 9.69747
R544 VDD1.n120 VDD1.n65 9.69747
R545 VDD1.n60 VDD1.n59 9.45567
R546 VDD1.n123 VDD1.n122 9.45567
R547 VDD1.n20 VDD1.n19 9.3005
R548 VDD1.n27 VDD1.n26 9.3005
R549 VDD1.n29 VDD1.n28 9.3005
R550 VDD1.n16 VDD1.n15 9.3005
R551 VDD1.n35 VDD1.n34 9.3005
R552 VDD1.n37 VDD1.n36 9.3005
R553 VDD1.n11 VDD1.n9 9.3005
R554 VDD1.n43 VDD1.n42 9.3005
R555 VDD1.n59 VDD1.n58 9.3005
R556 VDD1.n2 VDD1.n1 9.3005
R557 VDD1.n53 VDD1.n52 9.3005
R558 VDD1.n51 VDD1.n50 9.3005
R559 VDD1.n6 VDD1.n5 9.3005
R560 VDD1.n45 VDD1.n44 9.3005
R561 VDD1.n122 VDD1.n121 9.3005
R562 VDD1.n65 VDD1.n64 9.3005
R563 VDD1.n116 VDD1.n115 9.3005
R564 VDD1.n114 VDD1.n113 9.3005
R565 VDD1.n69 VDD1.n68 9.3005
R566 VDD1.n108 VDD1.n107 9.3005
R567 VDD1.n81 VDD1.n80 9.3005
R568 VDD1.n88 VDD1.n87 9.3005
R569 VDD1.n90 VDD1.n89 9.3005
R570 VDD1.n77 VDD1.n76 9.3005
R571 VDD1.n96 VDD1.n95 9.3005
R572 VDD1.n98 VDD1.n97 9.3005
R573 VDD1.n99 VDD1.n72 9.3005
R574 VDD1.n106 VDD1.n105 9.3005
R575 VDD1.n58 VDD1.n0 8.92171
R576 VDD1.n29 VDD1.n18 8.92171
R577 VDD1.n90 VDD1.n79 8.92171
R578 VDD1.n121 VDD1.n63 8.92171
R579 VDD1.n26 VDD1.n25 8.14595
R580 VDD1.n87 VDD1.n86 8.14595
R581 VDD1.n22 VDD1.n20 7.3702
R582 VDD1.n83 VDD1.n81 7.3702
R583 VDD1.n25 VDD1.n20 5.81868
R584 VDD1.n86 VDD1.n81 5.81868
R585 VDD1.n60 VDD1.n0 5.04292
R586 VDD1.n26 VDD1.n18 5.04292
R587 VDD1.n87 VDD1.n79 5.04292
R588 VDD1.n123 VDD1.n63 5.04292
R589 VDD1.n58 VDD1.n57 4.26717
R590 VDD1.n30 VDD1.n29 4.26717
R591 VDD1.n91 VDD1.n90 4.26717
R592 VDD1.n121 VDD1.n120 4.26717
R593 VDD1.n54 VDD1.n2 3.49141
R594 VDD1.n33 VDD1.n16 3.49141
R595 VDD1.n94 VDD1.n77 3.49141
R596 VDD1.n117 VDD1.n65 3.49141
R597 VDD1.n21 VDD1.n19 2.84303
R598 VDD1.n82 VDD1.n80 2.84303
R599 VDD1.n53 VDD1.n4 2.71565
R600 VDD1.n34 VDD1.n14 2.71565
R601 VDD1.n95 VDD1.n75 2.71565
R602 VDD1.n116 VDD1.n67 2.71565
R603 VDD1.n50 VDD1.n49 1.93989
R604 VDD1.n38 VDD1.n37 1.93989
R605 VDD1.n100 VDD1.n98 1.93989
R606 VDD1.n113 VDD1.n112 1.93989
R607 VDD1.n128 VDD1.t8 1.75271
R608 VDD1.n128 VDD1.t9 1.75271
R609 VDD1.n61 VDD1.t1 1.75271
R610 VDD1.n61 VDD1.t2 1.75271
R611 VDD1.n126 VDD1.t3 1.75271
R612 VDD1.n126 VDD1.t6 1.75271
R613 VDD1.n124 VDD1.t5 1.75271
R614 VDD1.n124 VDD1.t7 1.75271
R615 VDD1.n46 VDD1.n6 1.16414
R616 VDD1.n41 VDD1.n11 1.16414
R617 VDD1.n99 VDD1.n73 1.16414
R618 VDD1.n109 VDD1.n69 1.16414
R619 VDD1.n45 VDD1.n8 0.388379
R620 VDD1.n42 VDD1.n10 0.388379
R621 VDD1.n105 VDD1.n104 0.388379
R622 VDD1.n108 VDD1.n71 0.388379
R623 VDD1 VDD1.n129 0.381966
R624 VDD1 VDD1.n62 0.205241
R625 VDD1.n59 VDD1.n1 0.155672
R626 VDD1.n52 VDD1.n1 0.155672
R627 VDD1.n52 VDD1.n51 0.155672
R628 VDD1.n51 VDD1.n5 0.155672
R629 VDD1.n44 VDD1.n5 0.155672
R630 VDD1.n44 VDD1.n43 0.155672
R631 VDD1.n43 VDD1.n9 0.155672
R632 VDD1.n36 VDD1.n9 0.155672
R633 VDD1.n36 VDD1.n35 0.155672
R634 VDD1.n35 VDD1.n15 0.155672
R635 VDD1.n28 VDD1.n15 0.155672
R636 VDD1.n28 VDD1.n27 0.155672
R637 VDD1.n27 VDD1.n19 0.155672
R638 VDD1.n88 VDD1.n80 0.155672
R639 VDD1.n89 VDD1.n88 0.155672
R640 VDD1.n89 VDD1.n76 0.155672
R641 VDD1.n96 VDD1.n76 0.155672
R642 VDD1.n97 VDD1.n96 0.155672
R643 VDD1.n97 VDD1.n72 0.155672
R644 VDD1.n106 VDD1.n72 0.155672
R645 VDD1.n107 VDD1.n106 0.155672
R646 VDD1.n107 VDD1.n68 0.155672
R647 VDD1.n114 VDD1.n68 0.155672
R648 VDD1.n115 VDD1.n114 0.155672
R649 VDD1.n115 VDD1.n64 0.155672
R650 VDD1.n122 VDD1.n64 0.155672
R651 VDD1.n127 VDD1.n125 0.0917057
R652 B.n322 B.t7 989.659
R653 B.n328 B.t15 989.659
R654 B.n88 B.t11 989.659
R655 B.n86 B.t18 989.659
R656 B.n618 B.n617 585
R657 B.n619 B.n618 585
R658 B.n264 B.n85 585
R659 B.n263 B.n262 585
R660 B.n261 B.n260 585
R661 B.n259 B.n258 585
R662 B.n257 B.n256 585
R663 B.n255 B.n254 585
R664 B.n253 B.n252 585
R665 B.n251 B.n250 585
R666 B.n249 B.n248 585
R667 B.n247 B.n246 585
R668 B.n245 B.n244 585
R669 B.n243 B.n242 585
R670 B.n241 B.n240 585
R671 B.n239 B.n238 585
R672 B.n237 B.n236 585
R673 B.n235 B.n234 585
R674 B.n233 B.n232 585
R675 B.n231 B.n230 585
R676 B.n229 B.n228 585
R677 B.n227 B.n226 585
R678 B.n225 B.n224 585
R679 B.n223 B.n222 585
R680 B.n221 B.n220 585
R681 B.n219 B.n218 585
R682 B.n217 B.n216 585
R683 B.n215 B.n214 585
R684 B.n213 B.n212 585
R685 B.n211 B.n210 585
R686 B.n209 B.n208 585
R687 B.n207 B.n206 585
R688 B.n205 B.n204 585
R689 B.n203 B.n202 585
R690 B.n201 B.n200 585
R691 B.n199 B.n198 585
R692 B.n197 B.n196 585
R693 B.n195 B.n194 585
R694 B.n193 B.n192 585
R695 B.n191 B.n190 585
R696 B.n189 B.n188 585
R697 B.n186 B.n185 585
R698 B.n184 B.n183 585
R699 B.n182 B.n181 585
R700 B.n180 B.n179 585
R701 B.n178 B.n177 585
R702 B.n176 B.n175 585
R703 B.n174 B.n173 585
R704 B.n172 B.n171 585
R705 B.n170 B.n169 585
R706 B.n168 B.n167 585
R707 B.n166 B.n165 585
R708 B.n164 B.n163 585
R709 B.n162 B.n161 585
R710 B.n160 B.n159 585
R711 B.n158 B.n157 585
R712 B.n156 B.n155 585
R713 B.n154 B.n153 585
R714 B.n152 B.n151 585
R715 B.n150 B.n149 585
R716 B.n148 B.n147 585
R717 B.n146 B.n145 585
R718 B.n144 B.n143 585
R719 B.n142 B.n141 585
R720 B.n140 B.n139 585
R721 B.n138 B.n137 585
R722 B.n136 B.n135 585
R723 B.n134 B.n133 585
R724 B.n132 B.n131 585
R725 B.n130 B.n129 585
R726 B.n128 B.n127 585
R727 B.n126 B.n125 585
R728 B.n124 B.n123 585
R729 B.n122 B.n121 585
R730 B.n120 B.n119 585
R731 B.n118 B.n117 585
R732 B.n116 B.n115 585
R733 B.n114 B.n113 585
R734 B.n112 B.n111 585
R735 B.n110 B.n109 585
R736 B.n108 B.n107 585
R737 B.n106 B.n105 585
R738 B.n104 B.n103 585
R739 B.n102 B.n101 585
R740 B.n100 B.n99 585
R741 B.n98 B.n97 585
R742 B.n96 B.n95 585
R743 B.n94 B.n93 585
R744 B.n92 B.n91 585
R745 B.n39 B.n38 585
R746 B.n616 B.n40 585
R747 B.n620 B.n40 585
R748 B.n615 B.n614 585
R749 B.n614 B.n36 585
R750 B.n613 B.n35 585
R751 B.n626 B.n35 585
R752 B.n612 B.n34 585
R753 B.n627 B.n34 585
R754 B.n611 B.n33 585
R755 B.n628 B.n33 585
R756 B.n610 B.n609 585
R757 B.n609 B.n29 585
R758 B.n608 B.n28 585
R759 B.n634 B.n28 585
R760 B.n607 B.n27 585
R761 B.n635 B.n27 585
R762 B.n606 B.n26 585
R763 B.n636 B.n26 585
R764 B.n605 B.n604 585
R765 B.n604 B.n25 585
R766 B.n603 B.n21 585
R767 B.n642 B.n21 585
R768 B.n602 B.n20 585
R769 B.n643 B.n20 585
R770 B.n601 B.n19 585
R771 B.n644 B.n19 585
R772 B.n600 B.n599 585
R773 B.n599 B.n18 585
R774 B.n598 B.n14 585
R775 B.n650 B.n14 585
R776 B.n597 B.n13 585
R777 B.n651 B.n13 585
R778 B.n596 B.n12 585
R779 B.n652 B.n12 585
R780 B.n595 B.n594 585
R781 B.n594 B.n11 585
R782 B.n593 B.n7 585
R783 B.n658 B.n7 585
R784 B.n592 B.n6 585
R785 B.n659 B.n6 585
R786 B.n591 B.n5 585
R787 B.n660 B.n5 585
R788 B.n590 B.n589 585
R789 B.n589 B.n4 585
R790 B.n588 B.n265 585
R791 B.n588 B.n587 585
R792 B.n577 B.n266 585
R793 B.n580 B.n266 585
R794 B.n579 B.n578 585
R795 B.n581 B.n579 585
R796 B.n576 B.n270 585
R797 B.n273 B.n270 585
R798 B.n575 B.n574 585
R799 B.n574 B.n573 585
R800 B.n272 B.n271 585
R801 B.n566 B.n272 585
R802 B.n565 B.n564 585
R803 B.n567 B.n565 585
R804 B.n563 B.n277 585
R805 B.n280 B.n277 585
R806 B.n562 B.n561 585
R807 B.n561 B.n560 585
R808 B.n279 B.n278 585
R809 B.n553 B.n279 585
R810 B.n552 B.n551 585
R811 B.n554 B.n552 585
R812 B.n550 B.n285 585
R813 B.n285 B.n284 585
R814 B.n549 B.n548 585
R815 B.n548 B.n547 585
R816 B.n287 B.n286 585
R817 B.n288 B.n287 585
R818 B.n540 B.n539 585
R819 B.n541 B.n540 585
R820 B.n538 B.n293 585
R821 B.n293 B.n292 585
R822 B.n537 B.n536 585
R823 B.n536 B.n535 585
R824 B.n295 B.n294 585
R825 B.n296 B.n295 585
R826 B.n528 B.n527 585
R827 B.n529 B.n528 585
R828 B.n299 B.n298 585
R829 B.n351 B.n349 585
R830 B.n352 B.n348 585
R831 B.n352 B.n300 585
R832 B.n355 B.n354 585
R833 B.n356 B.n347 585
R834 B.n358 B.n357 585
R835 B.n360 B.n346 585
R836 B.n363 B.n362 585
R837 B.n364 B.n345 585
R838 B.n366 B.n365 585
R839 B.n368 B.n344 585
R840 B.n371 B.n370 585
R841 B.n372 B.n343 585
R842 B.n374 B.n373 585
R843 B.n376 B.n342 585
R844 B.n379 B.n378 585
R845 B.n380 B.n341 585
R846 B.n382 B.n381 585
R847 B.n384 B.n340 585
R848 B.n387 B.n386 585
R849 B.n388 B.n339 585
R850 B.n390 B.n389 585
R851 B.n392 B.n338 585
R852 B.n395 B.n394 585
R853 B.n396 B.n337 585
R854 B.n398 B.n397 585
R855 B.n400 B.n336 585
R856 B.n403 B.n402 585
R857 B.n404 B.n335 585
R858 B.n406 B.n405 585
R859 B.n408 B.n334 585
R860 B.n411 B.n410 585
R861 B.n412 B.n333 585
R862 B.n414 B.n413 585
R863 B.n416 B.n332 585
R864 B.n419 B.n418 585
R865 B.n420 B.n331 585
R866 B.n422 B.n421 585
R867 B.n424 B.n330 585
R868 B.n427 B.n426 585
R869 B.n429 B.n327 585
R870 B.n431 B.n430 585
R871 B.n433 B.n326 585
R872 B.n436 B.n435 585
R873 B.n437 B.n325 585
R874 B.n439 B.n438 585
R875 B.n441 B.n324 585
R876 B.n444 B.n443 585
R877 B.n445 B.n321 585
R878 B.n448 B.n447 585
R879 B.n450 B.n320 585
R880 B.n453 B.n452 585
R881 B.n454 B.n319 585
R882 B.n456 B.n455 585
R883 B.n458 B.n318 585
R884 B.n461 B.n460 585
R885 B.n462 B.n317 585
R886 B.n464 B.n463 585
R887 B.n466 B.n316 585
R888 B.n469 B.n468 585
R889 B.n470 B.n315 585
R890 B.n472 B.n471 585
R891 B.n474 B.n314 585
R892 B.n477 B.n476 585
R893 B.n478 B.n313 585
R894 B.n480 B.n479 585
R895 B.n482 B.n312 585
R896 B.n485 B.n484 585
R897 B.n486 B.n311 585
R898 B.n488 B.n487 585
R899 B.n490 B.n310 585
R900 B.n493 B.n492 585
R901 B.n494 B.n309 585
R902 B.n496 B.n495 585
R903 B.n498 B.n308 585
R904 B.n501 B.n500 585
R905 B.n502 B.n307 585
R906 B.n504 B.n503 585
R907 B.n506 B.n306 585
R908 B.n509 B.n508 585
R909 B.n510 B.n305 585
R910 B.n512 B.n511 585
R911 B.n514 B.n304 585
R912 B.n517 B.n516 585
R913 B.n518 B.n303 585
R914 B.n520 B.n519 585
R915 B.n522 B.n302 585
R916 B.n525 B.n524 585
R917 B.n526 B.n301 585
R918 B.n531 B.n530 585
R919 B.n530 B.n529 585
R920 B.n532 B.n297 585
R921 B.n297 B.n296 585
R922 B.n534 B.n533 585
R923 B.n535 B.n534 585
R924 B.n291 B.n290 585
R925 B.n292 B.n291 585
R926 B.n543 B.n542 585
R927 B.n542 B.n541 585
R928 B.n544 B.n289 585
R929 B.n289 B.n288 585
R930 B.n546 B.n545 585
R931 B.n547 B.n546 585
R932 B.n283 B.n282 585
R933 B.n284 B.n283 585
R934 B.n556 B.n555 585
R935 B.n555 B.n554 585
R936 B.n557 B.n281 585
R937 B.n553 B.n281 585
R938 B.n559 B.n558 585
R939 B.n560 B.n559 585
R940 B.n276 B.n275 585
R941 B.n280 B.n276 585
R942 B.n569 B.n568 585
R943 B.n568 B.n567 585
R944 B.n570 B.n274 585
R945 B.n566 B.n274 585
R946 B.n572 B.n571 585
R947 B.n573 B.n572 585
R948 B.n269 B.n268 585
R949 B.n273 B.n269 585
R950 B.n583 B.n582 585
R951 B.n582 B.n581 585
R952 B.n584 B.n267 585
R953 B.n580 B.n267 585
R954 B.n586 B.n585 585
R955 B.n587 B.n586 585
R956 B.n2 B.n0 585
R957 B.n4 B.n2 585
R958 B.n3 B.n1 585
R959 B.n659 B.n3 585
R960 B.n657 B.n656 585
R961 B.n658 B.n657 585
R962 B.n655 B.n8 585
R963 B.n11 B.n8 585
R964 B.n654 B.n653 585
R965 B.n653 B.n652 585
R966 B.n10 B.n9 585
R967 B.n651 B.n10 585
R968 B.n649 B.n648 585
R969 B.n650 B.n649 585
R970 B.n647 B.n15 585
R971 B.n18 B.n15 585
R972 B.n646 B.n645 585
R973 B.n645 B.n644 585
R974 B.n17 B.n16 585
R975 B.n643 B.n17 585
R976 B.n641 B.n640 585
R977 B.n642 B.n641 585
R978 B.n639 B.n22 585
R979 B.n25 B.n22 585
R980 B.n638 B.n637 585
R981 B.n637 B.n636 585
R982 B.n24 B.n23 585
R983 B.n635 B.n24 585
R984 B.n633 B.n632 585
R985 B.n634 B.n633 585
R986 B.n631 B.n30 585
R987 B.n30 B.n29 585
R988 B.n630 B.n629 585
R989 B.n629 B.n628 585
R990 B.n32 B.n31 585
R991 B.n627 B.n32 585
R992 B.n625 B.n624 585
R993 B.n626 B.n625 585
R994 B.n623 B.n37 585
R995 B.n37 B.n36 585
R996 B.n622 B.n621 585
R997 B.n621 B.n620 585
R998 B.n662 B.n661 585
R999 B.n661 B.n660 585
R1000 B.n530 B.n299 492.5
R1001 B.n621 B.n39 492.5
R1002 B.n528 B.n301 492.5
R1003 B.n618 B.n40 492.5
R1004 B.n322 B.t10 283.096
R1005 B.n86 B.t19 283.096
R1006 B.n328 B.t17 283.096
R1007 B.n88 B.t13 283.096
R1008 B.n323 B.t9 269.908
R1009 B.n87 B.t20 269.908
R1010 B.n329 B.t16 269.908
R1011 B.n89 B.t14 269.908
R1012 B.n619 B.n84 256.663
R1013 B.n619 B.n83 256.663
R1014 B.n619 B.n82 256.663
R1015 B.n619 B.n81 256.663
R1016 B.n619 B.n80 256.663
R1017 B.n619 B.n79 256.663
R1018 B.n619 B.n78 256.663
R1019 B.n619 B.n77 256.663
R1020 B.n619 B.n76 256.663
R1021 B.n619 B.n75 256.663
R1022 B.n619 B.n74 256.663
R1023 B.n619 B.n73 256.663
R1024 B.n619 B.n72 256.663
R1025 B.n619 B.n71 256.663
R1026 B.n619 B.n70 256.663
R1027 B.n619 B.n69 256.663
R1028 B.n619 B.n68 256.663
R1029 B.n619 B.n67 256.663
R1030 B.n619 B.n66 256.663
R1031 B.n619 B.n65 256.663
R1032 B.n619 B.n64 256.663
R1033 B.n619 B.n63 256.663
R1034 B.n619 B.n62 256.663
R1035 B.n619 B.n61 256.663
R1036 B.n619 B.n60 256.663
R1037 B.n619 B.n59 256.663
R1038 B.n619 B.n58 256.663
R1039 B.n619 B.n57 256.663
R1040 B.n619 B.n56 256.663
R1041 B.n619 B.n55 256.663
R1042 B.n619 B.n54 256.663
R1043 B.n619 B.n53 256.663
R1044 B.n619 B.n52 256.663
R1045 B.n619 B.n51 256.663
R1046 B.n619 B.n50 256.663
R1047 B.n619 B.n49 256.663
R1048 B.n619 B.n48 256.663
R1049 B.n619 B.n47 256.663
R1050 B.n619 B.n46 256.663
R1051 B.n619 B.n45 256.663
R1052 B.n619 B.n44 256.663
R1053 B.n619 B.n43 256.663
R1054 B.n619 B.n42 256.663
R1055 B.n619 B.n41 256.663
R1056 B.n350 B.n300 256.663
R1057 B.n353 B.n300 256.663
R1058 B.n359 B.n300 256.663
R1059 B.n361 B.n300 256.663
R1060 B.n367 B.n300 256.663
R1061 B.n369 B.n300 256.663
R1062 B.n375 B.n300 256.663
R1063 B.n377 B.n300 256.663
R1064 B.n383 B.n300 256.663
R1065 B.n385 B.n300 256.663
R1066 B.n391 B.n300 256.663
R1067 B.n393 B.n300 256.663
R1068 B.n399 B.n300 256.663
R1069 B.n401 B.n300 256.663
R1070 B.n407 B.n300 256.663
R1071 B.n409 B.n300 256.663
R1072 B.n415 B.n300 256.663
R1073 B.n417 B.n300 256.663
R1074 B.n423 B.n300 256.663
R1075 B.n425 B.n300 256.663
R1076 B.n432 B.n300 256.663
R1077 B.n434 B.n300 256.663
R1078 B.n440 B.n300 256.663
R1079 B.n442 B.n300 256.663
R1080 B.n449 B.n300 256.663
R1081 B.n451 B.n300 256.663
R1082 B.n457 B.n300 256.663
R1083 B.n459 B.n300 256.663
R1084 B.n465 B.n300 256.663
R1085 B.n467 B.n300 256.663
R1086 B.n473 B.n300 256.663
R1087 B.n475 B.n300 256.663
R1088 B.n481 B.n300 256.663
R1089 B.n483 B.n300 256.663
R1090 B.n489 B.n300 256.663
R1091 B.n491 B.n300 256.663
R1092 B.n497 B.n300 256.663
R1093 B.n499 B.n300 256.663
R1094 B.n505 B.n300 256.663
R1095 B.n507 B.n300 256.663
R1096 B.n513 B.n300 256.663
R1097 B.n515 B.n300 256.663
R1098 B.n521 B.n300 256.663
R1099 B.n523 B.n300 256.663
R1100 B.n530 B.n297 163.367
R1101 B.n534 B.n297 163.367
R1102 B.n534 B.n291 163.367
R1103 B.n542 B.n291 163.367
R1104 B.n542 B.n289 163.367
R1105 B.n546 B.n289 163.367
R1106 B.n546 B.n283 163.367
R1107 B.n555 B.n283 163.367
R1108 B.n555 B.n281 163.367
R1109 B.n559 B.n281 163.367
R1110 B.n559 B.n276 163.367
R1111 B.n568 B.n276 163.367
R1112 B.n568 B.n274 163.367
R1113 B.n572 B.n274 163.367
R1114 B.n572 B.n269 163.367
R1115 B.n582 B.n269 163.367
R1116 B.n582 B.n267 163.367
R1117 B.n586 B.n267 163.367
R1118 B.n586 B.n2 163.367
R1119 B.n661 B.n2 163.367
R1120 B.n661 B.n3 163.367
R1121 B.n657 B.n3 163.367
R1122 B.n657 B.n8 163.367
R1123 B.n653 B.n8 163.367
R1124 B.n653 B.n10 163.367
R1125 B.n649 B.n10 163.367
R1126 B.n649 B.n15 163.367
R1127 B.n645 B.n15 163.367
R1128 B.n645 B.n17 163.367
R1129 B.n641 B.n17 163.367
R1130 B.n641 B.n22 163.367
R1131 B.n637 B.n22 163.367
R1132 B.n637 B.n24 163.367
R1133 B.n633 B.n24 163.367
R1134 B.n633 B.n30 163.367
R1135 B.n629 B.n30 163.367
R1136 B.n629 B.n32 163.367
R1137 B.n625 B.n32 163.367
R1138 B.n625 B.n37 163.367
R1139 B.n621 B.n37 163.367
R1140 B.n352 B.n351 163.367
R1141 B.n354 B.n352 163.367
R1142 B.n358 B.n347 163.367
R1143 B.n362 B.n360 163.367
R1144 B.n366 B.n345 163.367
R1145 B.n370 B.n368 163.367
R1146 B.n374 B.n343 163.367
R1147 B.n378 B.n376 163.367
R1148 B.n382 B.n341 163.367
R1149 B.n386 B.n384 163.367
R1150 B.n390 B.n339 163.367
R1151 B.n394 B.n392 163.367
R1152 B.n398 B.n337 163.367
R1153 B.n402 B.n400 163.367
R1154 B.n406 B.n335 163.367
R1155 B.n410 B.n408 163.367
R1156 B.n414 B.n333 163.367
R1157 B.n418 B.n416 163.367
R1158 B.n422 B.n331 163.367
R1159 B.n426 B.n424 163.367
R1160 B.n431 B.n327 163.367
R1161 B.n435 B.n433 163.367
R1162 B.n439 B.n325 163.367
R1163 B.n443 B.n441 163.367
R1164 B.n448 B.n321 163.367
R1165 B.n452 B.n450 163.367
R1166 B.n456 B.n319 163.367
R1167 B.n460 B.n458 163.367
R1168 B.n464 B.n317 163.367
R1169 B.n468 B.n466 163.367
R1170 B.n472 B.n315 163.367
R1171 B.n476 B.n474 163.367
R1172 B.n480 B.n313 163.367
R1173 B.n484 B.n482 163.367
R1174 B.n488 B.n311 163.367
R1175 B.n492 B.n490 163.367
R1176 B.n496 B.n309 163.367
R1177 B.n500 B.n498 163.367
R1178 B.n504 B.n307 163.367
R1179 B.n508 B.n506 163.367
R1180 B.n512 B.n305 163.367
R1181 B.n516 B.n514 163.367
R1182 B.n520 B.n303 163.367
R1183 B.n524 B.n522 163.367
R1184 B.n528 B.n295 163.367
R1185 B.n536 B.n295 163.367
R1186 B.n536 B.n293 163.367
R1187 B.n540 B.n293 163.367
R1188 B.n540 B.n287 163.367
R1189 B.n548 B.n287 163.367
R1190 B.n548 B.n285 163.367
R1191 B.n552 B.n285 163.367
R1192 B.n552 B.n279 163.367
R1193 B.n561 B.n279 163.367
R1194 B.n561 B.n277 163.367
R1195 B.n565 B.n277 163.367
R1196 B.n565 B.n272 163.367
R1197 B.n574 B.n272 163.367
R1198 B.n574 B.n270 163.367
R1199 B.n579 B.n270 163.367
R1200 B.n579 B.n266 163.367
R1201 B.n588 B.n266 163.367
R1202 B.n589 B.n588 163.367
R1203 B.n589 B.n5 163.367
R1204 B.n6 B.n5 163.367
R1205 B.n7 B.n6 163.367
R1206 B.n594 B.n7 163.367
R1207 B.n594 B.n12 163.367
R1208 B.n13 B.n12 163.367
R1209 B.n14 B.n13 163.367
R1210 B.n599 B.n14 163.367
R1211 B.n599 B.n19 163.367
R1212 B.n20 B.n19 163.367
R1213 B.n21 B.n20 163.367
R1214 B.n604 B.n21 163.367
R1215 B.n604 B.n26 163.367
R1216 B.n27 B.n26 163.367
R1217 B.n28 B.n27 163.367
R1218 B.n609 B.n28 163.367
R1219 B.n609 B.n33 163.367
R1220 B.n34 B.n33 163.367
R1221 B.n35 B.n34 163.367
R1222 B.n614 B.n35 163.367
R1223 B.n614 B.n40 163.367
R1224 B.n93 B.n92 163.367
R1225 B.n97 B.n96 163.367
R1226 B.n101 B.n100 163.367
R1227 B.n105 B.n104 163.367
R1228 B.n109 B.n108 163.367
R1229 B.n113 B.n112 163.367
R1230 B.n117 B.n116 163.367
R1231 B.n121 B.n120 163.367
R1232 B.n125 B.n124 163.367
R1233 B.n129 B.n128 163.367
R1234 B.n133 B.n132 163.367
R1235 B.n137 B.n136 163.367
R1236 B.n141 B.n140 163.367
R1237 B.n145 B.n144 163.367
R1238 B.n149 B.n148 163.367
R1239 B.n153 B.n152 163.367
R1240 B.n157 B.n156 163.367
R1241 B.n161 B.n160 163.367
R1242 B.n165 B.n164 163.367
R1243 B.n169 B.n168 163.367
R1244 B.n173 B.n172 163.367
R1245 B.n177 B.n176 163.367
R1246 B.n181 B.n180 163.367
R1247 B.n185 B.n184 163.367
R1248 B.n190 B.n189 163.367
R1249 B.n194 B.n193 163.367
R1250 B.n198 B.n197 163.367
R1251 B.n202 B.n201 163.367
R1252 B.n206 B.n205 163.367
R1253 B.n210 B.n209 163.367
R1254 B.n214 B.n213 163.367
R1255 B.n218 B.n217 163.367
R1256 B.n222 B.n221 163.367
R1257 B.n226 B.n225 163.367
R1258 B.n230 B.n229 163.367
R1259 B.n234 B.n233 163.367
R1260 B.n238 B.n237 163.367
R1261 B.n242 B.n241 163.367
R1262 B.n246 B.n245 163.367
R1263 B.n250 B.n249 163.367
R1264 B.n254 B.n253 163.367
R1265 B.n258 B.n257 163.367
R1266 B.n262 B.n261 163.367
R1267 B.n618 B.n85 163.367
R1268 B.n529 B.n300 86.9387
R1269 B.n620 B.n619 86.9387
R1270 B.n350 B.n299 71.676
R1271 B.n354 B.n353 71.676
R1272 B.n359 B.n358 71.676
R1273 B.n362 B.n361 71.676
R1274 B.n367 B.n366 71.676
R1275 B.n370 B.n369 71.676
R1276 B.n375 B.n374 71.676
R1277 B.n378 B.n377 71.676
R1278 B.n383 B.n382 71.676
R1279 B.n386 B.n385 71.676
R1280 B.n391 B.n390 71.676
R1281 B.n394 B.n393 71.676
R1282 B.n399 B.n398 71.676
R1283 B.n402 B.n401 71.676
R1284 B.n407 B.n406 71.676
R1285 B.n410 B.n409 71.676
R1286 B.n415 B.n414 71.676
R1287 B.n418 B.n417 71.676
R1288 B.n423 B.n422 71.676
R1289 B.n426 B.n425 71.676
R1290 B.n432 B.n431 71.676
R1291 B.n435 B.n434 71.676
R1292 B.n440 B.n439 71.676
R1293 B.n443 B.n442 71.676
R1294 B.n449 B.n448 71.676
R1295 B.n452 B.n451 71.676
R1296 B.n457 B.n456 71.676
R1297 B.n460 B.n459 71.676
R1298 B.n465 B.n464 71.676
R1299 B.n468 B.n467 71.676
R1300 B.n473 B.n472 71.676
R1301 B.n476 B.n475 71.676
R1302 B.n481 B.n480 71.676
R1303 B.n484 B.n483 71.676
R1304 B.n489 B.n488 71.676
R1305 B.n492 B.n491 71.676
R1306 B.n497 B.n496 71.676
R1307 B.n500 B.n499 71.676
R1308 B.n505 B.n504 71.676
R1309 B.n508 B.n507 71.676
R1310 B.n513 B.n512 71.676
R1311 B.n516 B.n515 71.676
R1312 B.n521 B.n520 71.676
R1313 B.n524 B.n523 71.676
R1314 B.n41 B.n39 71.676
R1315 B.n93 B.n42 71.676
R1316 B.n97 B.n43 71.676
R1317 B.n101 B.n44 71.676
R1318 B.n105 B.n45 71.676
R1319 B.n109 B.n46 71.676
R1320 B.n113 B.n47 71.676
R1321 B.n117 B.n48 71.676
R1322 B.n121 B.n49 71.676
R1323 B.n125 B.n50 71.676
R1324 B.n129 B.n51 71.676
R1325 B.n133 B.n52 71.676
R1326 B.n137 B.n53 71.676
R1327 B.n141 B.n54 71.676
R1328 B.n145 B.n55 71.676
R1329 B.n149 B.n56 71.676
R1330 B.n153 B.n57 71.676
R1331 B.n157 B.n58 71.676
R1332 B.n161 B.n59 71.676
R1333 B.n165 B.n60 71.676
R1334 B.n169 B.n61 71.676
R1335 B.n173 B.n62 71.676
R1336 B.n177 B.n63 71.676
R1337 B.n181 B.n64 71.676
R1338 B.n185 B.n65 71.676
R1339 B.n190 B.n66 71.676
R1340 B.n194 B.n67 71.676
R1341 B.n198 B.n68 71.676
R1342 B.n202 B.n69 71.676
R1343 B.n206 B.n70 71.676
R1344 B.n210 B.n71 71.676
R1345 B.n214 B.n72 71.676
R1346 B.n218 B.n73 71.676
R1347 B.n222 B.n74 71.676
R1348 B.n226 B.n75 71.676
R1349 B.n230 B.n76 71.676
R1350 B.n234 B.n77 71.676
R1351 B.n238 B.n78 71.676
R1352 B.n242 B.n79 71.676
R1353 B.n246 B.n80 71.676
R1354 B.n250 B.n81 71.676
R1355 B.n254 B.n82 71.676
R1356 B.n258 B.n83 71.676
R1357 B.n262 B.n84 71.676
R1358 B.n85 B.n84 71.676
R1359 B.n261 B.n83 71.676
R1360 B.n257 B.n82 71.676
R1361 B.n253 B.n81 71.676
R1362 B.n249 B.n80 71.676
R1363 B.n245 B.n79 71.676
R1364 B.n241 B.n78 71.676
R1365 B.n237 B.n77 71.676
R1366 B.n233 B.n76 71.676
R1367 B.n229 B.n75 71.676
R1368 B.n225 B.n74 71.676
R1369 B.n221 B.n73 71.676
R1370 B.n217 B.n72 71.676
R1371 B.n213 B.n71 71.676
R1372 B.n209 B.n70 71.676
R1373 B.n205 B.n69 71.676
R1374 B.n201 B.n68 71.676
R1375 B.n197 B.n67 71.676
R1376 B.n193 B.n66 71.676
R1377 B.n189 B.n65 71.676
R1378 B.n184 B.n64 71.676
R1379 B.n180 B.n63 71.676
R1380 B.n176 B.n62 71.676
R1381 B.n172 B.n61 71.676
R1382 B.n168 B.n60 71.676
R1383 B.n164 B.n59 71.676
R1384 B.n160 B.n58 71.676
R1385 B.n156 B.n57 71.676
R1386 B.n152 B.n56 71.676
R1387 B.n148 B.n55 71.676
R1388 B.n144 B.n54 71.676
R1389 B.n140 B.n53 71.676
R1390 B.n136 B.n52 71.676
R1391 B.n132 B.n51 71.676
R1392 B.n128 B.n50 71.676
R1393 B.n124 B.n49 71.676
R1394 B.n120 B.n48 71.676
R1395 B.n116 B.n47 71.676
R1396 B.n112 B.n46 71.676
R1397 B.n108 B.n45 71.676
R1398 B.n104 B.n44 71.676
R1399 B.n100 B.n43 71.676
R1400 B.n96 B.n42 71.676
R1401 B.n92 B.n41 71.676
R1402 B.n351 B.n350 71.676
R1403 B.n353 B.n347 71.676
R1404 B.n360 B.n359 71.676
R1405 B.n361 B.n345 71.676
R1406 B.n368 B.n367 71.676
R1407 B.n369 B.n343 71.676
R1408 B.n376 B.n375 71.676
R1409 B.n377 B.n341 71.676
R1410 B.n384 B.n383 71.676
R1411 B.n385 B.n339 71.676
R1412 B.n392 B.n391 71.676
R1413 B.n393 B.n337 71.676
R1414 B.n400 B.n399 71.676
R1415 B.n401 B.n335 71.676
R1416 B.n408 B.n407 71.676
R1417 B.n409 B.n333 71.676
R1418 B.n416 B.n415 71.676
R1419 B.n417 B.n331 71.676
R1420 B.n424 B.n423 71.676
R1421 B.n425 B.n327 71.676
R1422 B.n433 B.n432 71.676
R1423 B.n434 B.n325 71.676
R1424 B.n441 B.n440 71.676
R1425 B.n442 B.n321 71.676
R1426 B.n450 B.n449 71.676
R1427 B.n451 B.n319 71.676
R1428 B.n458 B.n457 71.676
R1429 B.n459 B.n317 71.676
R1430 B.n466 B.n465 71.676
R1431 B.n467 B.n315 71.676
R1432 B.n474 B.n473 71.676
R1433 B.n475 B.n313 71.676
R1434 B.n482 B.n481 71.676
R1435 B.n483 B.n311 71.676
R1436 B.n490 B.n489 71.676
R1437 B.n491 B.n309 71.676
R1438 B.n498 B.n497 71.676
R1439 B.n499 B.n307 71.676
R1440 B.n506 B.n505 71.676
R1441 B.n507 B.n305 71.676
R1442 B.n514 B.n513 71.676
R1443 B.n515 B.n303 71.676
R1444 B.n522 B.n521 71.676
R1445 B.n523 B.n301 71.676
R1446 B.n446 B.n323 59.5399
R1447 B.n428 B.n329 59.5399
R1448 B.n90 B.n89 59.5399
R1449 B.n187 B.n87 59.5399
R1450 B.n529 B.n296 45.1287
R1451 B.n535 B.n296 45.1287
R1452 B.n535 B.n292 45.1287
R1453 B.n541 B.n292 45.1287
R1454 B.n547 B.n288 45.1287
R1455 B.n547 B.n284 45.1287
R1456 B.n554 B.n284 45.1287
R1457 B.n554 B.n553 45.1287
R1458 B.n560 B.n280 45.1287
R1459 B.n567 B.n566 45.1287
R1460 B.n573 B.n273 45.1287
R1461 B.n581 B.n580 45.1287
R1462 B.n587 B.n4 45.1287
R1463 B.n660 B.n4 45.1287
R1464 B.n660 B.n659 45.1287
R1465 B.n659 B.n658 45.1287
R1466 B.n652 B.n11 45.1287
R1467 B.n651 B.n650 45.1287
R1468 B.n644 B.n18 45.1287
R1469 B.n643 B.n642 45.1287
R1470 B.n636 B.n25 45.1287
R1471 B.n636 B.n635 45.1287
R1472 B.n635 B.n634 45.1287
R1473 B.n634 B.n29 45.1287
R1474 B.n628 B.n627 45.1287
R1475 B.n627 B.n626 45.1287
R1476 B.n626 B.n36 45.1287
R1477 B.n620 B.n36 45.1287
R1478 B.t8 B.n288 36.5013
R1479 B.t12 B.n29 36.5013
R1480 B.n622 B.n38 32.0005
R1481 B.n617 B.n616 32.0005
R1482 B.n527 B.n526 32.0005
R1483 B.n531 B.n298 32.0005
R1484 B.n560 B.t22 27.2102
R1485 B.n567 B.t5 27.2102
R1486 B.n573 B.t23 27.2102
R1487 B.n581 B.t4 27.2102
R1488 B.n587 B.t3 27.2102
R1489 B.n658 B.t6 27.2102
R1490 B.n652 B.t1 27.2102
R1491 B.n650 B.t21 27.2102
R1492 B.n644 B.t2 27.2102
R1493 B.n642 B.t0 27.2102
R1494 B B.n662 18.0485
R1495 B.n553 B.t22 17.9191
R1496 B.n280 B.t5 17.9191
R1497 B.n566 B.t23 17.9191
R1498 B.n273 B.t4 17.9191
R1499 B.n580 B.t3 17.9191
R1500 B.n11 B.t6 17.9191
R1501 B.t1 B.n651 17.9191
R1502 B.n18 B.t21 17.9191
R1503 B.t2 B.n643 17.9191
R1504 B.n25 B.t0 17.9191
R1505 B.n323 B.n322 13.1884
R1506 B.n329 B.n328 13.1884
R1507 B.n89 B.n88 13.1884
R1508 B.n87 B.n86 13.1884
R1509 B.n91 B.n38 10.6151
R1510 B.n94 B.n91 10.6151
R1511 B.n95 B.n94 10.6151
R1512 B.n98 B.n95 10.6151
R1513 B.n99 B.n98 10.6151
R1514 B.n102 B.n99 10.6151
R1515 B.n103 B.n102 10.6151
R1516 B.n106 B.n103 10.6151
R1517 B.n107 B.n106 10.6151
R1518 B.n110 B.n107 10.6151
R1519 B.n111 B.n110 10.6151
R1520 B.n114 B.n111 10.6151
R1521 B.n115 B.n114 10.6151
R1522 B.n118 B.n115 10.6151
R1523 B.n119 B.n118 10.6151
R1524 B.n122 B.n119 10.6151
R1525 B.n123 B.n122 10.6151
R1526 B.n126 B.n123 10.6151
R1527 B.n127 B.n126 10.6151
R1528 B.n130 B.n127 10.6151
R1529 B.n131 B.n130 10.6151
R1530 B.n134 B.n131 10.6151
R1531 B.n135 B.n134 10.6151
R1532 B.n138 B.n135 10.6151
R1533 B.n139 B.n138 10.6151
R1534 B.n142 B.n139 10.6151
R1535 B.n143 B.n142 10.6151
R1536 B.n146 B.n143 10.6151
R1537 B.n147 B.n146 10.6151
R1538 B.n150 B.n147 10.6151
R1539 B.n151 B.n150 10.6151
R1540 B.n154 B.n151 10.6151
R1541 B.n155 B.n154 10.6151
R1542 B.n158 B.n155 10.6151
R1543 B.n159 B.n158 10.6151
R1544 B.n162 B.n159 10.6151
R1545 B.n163 B.n162 10.6151
R1546 B.n166 B.n163 10.6151
R1547 B.n167 B.n166 10.6151
R1548 B.n171 B.n170 10.6151
R1549 B.n174 B.n171 10.6151
R1550 B.n175 B.n174 10.6151
R1551 B.n178 B.n175 10.6151
R1552 B.n179 B.n178 10.6151
R1553 B.n182 B.n179 10.6151
R1554 B.n183 B.n182 10.6151
R1555 B.n186 B.n183 10.6151
R1556 B.n191 B.n188 10.6151
R1557 B.n192 B.n191 10.6151
R1558 B.n195 B.n192 10.6151
R1559 B.n196 B.n195 10.6151
R1560 B.n199 B.n196 10.6151
R1561 B.n200 B.n199 10.6151
R1562 B.n203 B.n200 10.6151
R1563 B.n204 B.n203 10.6151
R1564 B.n207 B.n204 10.6151
R1565 B.n208 B.n207 10.6151
R1566 B.n211 B.n208 10.6151
R1567 B.n212 B.n211 10.6151
R1568 B.n215 B.n212 10.6151
R1569 B.n216 B.n215 10.6151
R1570 B.n219 B.n216 10.6151
R1571 B.n220 B.n219 10.6151
R1572 B.n223 B.n220 10.6151
R1573 B.n224 B.n223 10.6151
R1574 B.n227 B.n224 10.6151
R1575 B.n228 B.n227 10.6151
R1576 B.n231 B.n228 10.6151
R1577 B.n232 B.n231 10.6151
R1578 B.n235 B.n232 10.6151
R1579 B.n236 B.n235 10.6151
R1580 B.n239 B.n236 10.6151
R1581 B.n240 B.n239 10.6151
R1582 B.n243 B.n240 10.6151
R1583 B.n244 B.n243 10.6151
R1584 B.n247 B.n244 10.6151
R1585 B.n248 B.n247 10.6151
R1586 B.n251 B.n248 10.6151
R1587 B.n252 B.n251 10.6151
R1588 B.n255 B.n252 10.6151
R1589 B.n256 B.n255 10.6151
R1590 B.n259 B.n256 10.6151
R1591 B.n260 B.n259 10.6151
R1592 B.n263 B.n260 10.6151
R1593 B.n264 B.n263 10.6151
R1594 B.n617 B.n264 10.6151
R1595 B.n527 B.n294 10.6151
R1596 B.n537 B.n294 10.6151
R1597 B.n538 B.n537 10.6151
R1598 B.n539 B.n538 10.6151
R1599 B.n539 B.n286 10.6151
R1600 B.n549 B.n286 10.6151
R1601 B.n550 B.n549 10.6151
R1602 B.n551 B.n550 10.6151
R1603 B.n551 B.n278 10.6151
R1604 B.n562 B.n278 10.6151
R1605 B.n563 B.n562 10.6151
R1606 B.n564 B.n563 10.6151
R1607 B.n564 B.n271 10.6151
R1608 B.n575 B.n271 10.6151
R1609 B.n576 B.n575 10.6151
R1610 B.n578 B.n576 10.6151
R1611 B.n578 B.n577 10.6151
R1612 B.n577 B.n265 10.6151
R1613 B.n590 B.n265 10.6151
R1614 B.n591 B.n590 10.6151
R1615 B.n592 B.n591 10.6151
R1616 B.n593 B.n592 10.6151
R1617 B.n595 B.n593 10.6151
R1618 B.n596 B.n595 10.6151
R1619 B.n597 B.n596 10.6151
R1620 B.n598 B.n597 10.6151
R1621 B.n600 B.n598 10.6151
R1622 B.n601 B.n600 10.6151
R1623 B.n602 B.n601 10.6151
R1624 B.n603 B.n602 10.6151
R1625 B.n605 B.n603 10.6151
R1626 B.n606 B.n605 10.6151
R1627 B.n607 B.n606 10.6151
R1628 B.n608 B.n607 10.6151
R1629 B.n610 B.n608 10.6151
R1630 B.n611 B.n610 10.6151
R1631 B.n612 B.n611 10.6151
R1632 B.n613 B.n612 10.6151
R1633 B.n615 B.n613 10.6151
R1634 B.n616 B.n615 10.6151
R1635 B.n349 B.n298 10.6151
R1636 B.n349 B.n348 10.6151
R1637 B.n355 B.n348 10.6151
R1638 B.n356 B.n355 10.6151
R1639 B.n357 B.n356 10.6151
R1640 B.n357 B.n346 10.6151
R1641 B.n363 B.n346 10.6151
R1642 B.n364 B.n363 10.6151
R1643 B.n365 B.n364 10.6151
R1644 B.n365 B.n344 10.6151
R1645 B.n371 B.n344 10.6151
R1646 B.n372 B.n371 10.6151
R1647 B.n373 B.n372 10.6151
R1648 B.n373 B.n342 10.6151
R1649 B.n379 B.n342 10.6151
R1650 B.n380 B.n379 10.6151
R1651 B.n381 B.n380 10.6151
R1652 B.n381 B.n340 10.6151
R1653 B.n387 B.n340 10.6151
R1654 B.n388 B.n387 10.6151
R1655 B.n389 B.n388 10.6151
R1656 B.n389 B.n338 10.6151
R1657 B.n395 B.n338 10.6151
R1658 B.n396 B.n395 10.6151
R1659 B.n397 B.n396 10.6151
R1660 B.n397 B.n336 10.6151
R1661 B.n403 B.n336 10.6151
R1662 B.n404 B.n403 10.6151
R1663 B.n405 B.n404 10.6151
R1664 B.n405 B.n334 10.6151
R1665 B.n411 B.n334 10.6151
R1666 B.n412 B.n411 10.6151
R1667 B.n413 B.n412 10.6151
R1668 B.n413 B.n332 10.6151
R1669 B.n419 B.n332 10.6151
R1670 B.n420 B.n419 10.6151
R1671 B.n421 B.n420 10.6151
R1672 B.n421 B.n330 10.6151
R1673 B.n427 B.n330 10.6151
R1674 B.n430 B.n429 10.6151
R1675 B.n430 B.n326 10.6151
R1676 B.n436 B.n326 10.6151
R1677 B.n437 B.n436 10.6151
R1678 B.n438 B.n437 10.6151
R1679 B.n438 B.n324 10.6151
R1680 B.n444 B.n324 10.6151
R1681 B.n445 B.n444 10.6151
R1682 B.n447 B.n320 10.6151
R1683 B.n453 B.n320 10.6151
R1684 B.n454 B.n453 10.6151
R1685 B.n455 B.n454 10.6151
R1686 B.n455 B.n318 10.6151
R1687 B.n461 B.n318 10.6151
R1688 B.n462 B.n461 10.6151
R1689 B.n463 B.n462 10.6151
R1690 B.n463 B.n316 10.6151
R1691 B.n469 B.n316 10.6151
R1692 B.n470 B.n469 10.6151
R1693 B.n471 B.n470 10.6151
R1694 B.n471 B.n314 10.6151
R1695 B.n477 B.n314 10.6151
R1696 B.n478 B.n477 10.6151
R1697 B.n479 B.n478 10.6151
R1698 B.n479 B.n312 10.6151
R1699 B.n485 B.n312 10.6151
R1700 B.n486 B.n485 10.6151
R1701 B.n487 B.n486 10.6151
R1702 B.n487 B.n310 10.6151
R1703 B.n493 B.n310 10.6151
R1704 B.n494 B.n493 10.6151
R1705 B.n495 B.n494 10.6151
R1706 B.n495 B.n308 10.6151
R1707 B.n501 B.n308 10.6151
R1708 B.n502 B.n501 10.6151
R1709 B.n503 B.n502 10.6151
R1710 B.n503 B.n306 10.6151
R1711 B.n509 B.n306 10.6151
R1712 B.n510 B.n509 10.6151
R1713 B.n511 B.n510 10.6151
R1714 B.n511 B.n304 10.6151
R1715 B.n517 B.n304 10.6151
R1716 B.n518 B.n517 10.6151
R1717 B.n519 B.n518 10.6151
R1718 B.n519 B.n302 10.6151
R1719 B.n525 B.n302 10.6151
R1720 B.n526 B.n525 10.6151
R1721 B.n532 B.n531 10.6151
R1722 B.n533 B.n532 10.6151
R1723 B.n533 B.n290 10.6151
R1724 B.n543 B.n290 10.6151
R1725 B.n544 B.n543 10.6151
R1726 B.n545 B.n544 10.6151
R1727 B.n545 B.n282 10.6151
R1728 B.n556 B.n282 10.6151
R1729 B.n557 B.n556 10.6151
R1730 B.n558 B.n557 10.6151
R1731 B.n558 B.n275 10.6151
R1732 B.n569 B.n275 10.6151
R1733 B.n570 B.n569 10.6151
R1734 B.n571 B.n570 10.6151
R1735 B.n571 B.n268 10.6151
R1736 B.n583 B.n268 10.6151
R1737 B.n584 B.n583 10.6151
R1738 B.n585 B.n584 10.6151
R1739 B.n585 B.n0 10.6151
R1740 B.n656 B.n1 10.6151
R1741 B.n656 B.n655 10.6151
R1742 B.n655 B.n654 10.6151
R1743 B.n654 B.n9 10.6151
R1744 B.n648 B.n9 10.6151
R1745 B.n648 B.n647 10.6151
R1746 B.n647 B.n646 10.6151
R1747 B.n646 B.n16 10.6151
R1748 B.n640 B.n16 10.6151
R1749 B.n640 B.n639 10.6151
R1750 B.n639 B.n638 10.6151
R1751 B.n638 B.n23 10.6151
R1752 B.n632 B.n23 10.6151
R1753 B.n632 B.n631 10.6151
R1754 B.n631 B.n630 10.6151
R1755 B.n630 B.n31 10.6151
R1756 B.n624 B.n31 10.6151
R1757 B.n624 B.n623 10.6151
R1758 B.n623 B.n622 10.6151
R1759 B.n541 B.t8 8.62795
R1760 B.n628 B.t12 8.62795
R1761 B.n170 B.n90 6.5566
R1762 B.n187 B.n186 6.5566
R1763 B.n429 B.n428 6.5566
R1764 B.n446 B.n445 6.5566
R1765 B.n167 B.n90 4.05904
R1766 B.n188 B.n187 4.05904
R1767 B.n428 B.n427 4.05904
R1768 B.n447 B.n446 4.05904
R1769 B.n662 B.n0 2.81026
R1770 B.n662 B.n1 2.81026
R1771 VN.n9 VN.t4 918.721
R1772 VN.n3 VN.t0 918.721
R1773 VN.n14 VN.t2 918.721
R1774 VN.n20 VN.t7 918.721
R1775 VN.n2 VN.t5 891.701
R1776 VN.n6 VN.t9 891.701
R1777 VN.n8 VN.t1 891.701
R1778 VN.n13 VN.t3 891.701
R1779 VN.n17 VN.t8 891.701
R1780 VN.n19 VN.t6 891.701
R1781 VN.n15 VN.n14 161.489
R1782 VN.n4 VN.n3 161.489
R1783 VN.n10 VN.n9 161.3
R1784 VN.n21 VN.n20 161.3
R1785 VN.n18 VN.n11 161.3
R1786 VN.n17 VN.n16 161.3
R1787 VN.n15 VN.n12 161.3
R1788 VN.n7 VN.n0 161.3
R1789 VN.n6 VN.n5 161.3
R1790 VN.n4 VN.n1 161.3
R1791 VN.n6 VN.n1 47.4702
R1792 VN.n7 VN.n6 47.4702
R1793 VN.n17 VN.n12 47.4702
R1794 VN.n18 VN.n17 47.4702
R1795 VN VN.n21 40.8736
R1796 VN.n3 VN.n2 21.1793
R1797 VN.n9 VN.n8 21.1793
R1798 VN.n14 VN.n13 21.1793
R1799 VN.n20 VN.n19 21.1793
R1800 VN.n2 VN.n1 0.730803
R1801 VN.n8 VN.n7 0.730803
R1802 VN.n13 VN.n12 0.730803
R1803 VN.n19 VN.n18 0.730803
R1804 VN.n21 VN.n11 0.189894
R1805 VN.n16 VN.n11 0.189894
R1806 VN.n16 VN.n15 0.189894
R1807 VN.n5 VN.n4 0.189894
R1808 VN.n5 VN.n0 0.189894
R1809 VN.n10 VN.n0 0.189894
R1810 VN VN.n10 0.0516364
R1811 VDD2.n121 VDD2.n65 289.615
R1812 VDD2.n56 VDD2.n0 289.615
R1813 VDD2.n122 VDD2.n121 185
R1814 VDD2.n120 VDD2.n119 185
R1815 VDD2.n69 VDD2.n68 185
R1816 VDD2.n114 VDD2.n113 185
R1817 VDD2.n112 VDD2.n111 185
R1818 VDD2.n73 VDD2.n72 185
R1819 VDD2.n77 VDD2.n75 185
R1820 VDD2.n106 VDD2.n105 185
R1821 VDD2.n104 VDD2.n103 185
R1822 VDD2.n79 VDD2.n78 185
R1823 VDD2.n98 VDD2.n97 185
R1824 VDD2.n96 VDD2.n95 185
R1825 VDD2.n83 VDD2.n82 185
R1826 VDD2.n90 VDD2.n89 185
R1827 VDD2.n88 VDD2.n87 185
R1828 VDD2.n21 VDD2.n20 185
R1829 VDD2.n23 VDD2.n22 185
R1830 VDD2.n16 VDD2.n15 185
R1831 VDD2.n29 VDD2.n28 185
R1832 VDD2.n31 VDD2.n30 185
R1833 VDD2.n12 VDD2.n11 185
R1834 VDD2.n38 VDD2.n37 185
R1835 VDD2.n39 VDD2.n10 185
R1836 VDD2.n41 VDD2.n40 185
R1837 VDD2.n8 VDD2.n7 185
R1838 VDD2.n47 VDD2.n46 185
R1839 VDD2.n49 VDD2.n48 185
R1840 VDD2.n4 VDD2.n3 185
R1841 VDD2.n55 VDD2.n54 185
R1842 VDD2.n57 VDD2.n56 185
R1843 VDD2.n86 VDD2.t2 149.524
R1844 VDD2.n19 VDD2.t9 149.524
R1845 VDD2.n121 VDD2.n120 104.615
R1846 VDD2.n120 VDD2.n68 104.615
R1847 VDD2.n113 VDD2.n68 104.615
R1848 VDD2.n113 VDD2.n112 104.615
R1849 VDD2.n112 VDD2.n72 104.615
R1850 VDD2.n77 VDD2.n72 104.615
R1851 VDD2.n105 VDD2.n77 104.615
R1852 VDD2.n105 VDD2.n104 104.615
R1853 VDD2.n104 VDD2.n78 104.615
R1854 VDD2.n97 VDD2.n78 104.615
R1855 VDD2.n97 VDD2.n96 104.615
R1856 VDD2.n96 VDD2.n82 104.615
R1857 VDD2.n89 VDD2.n82 104.615
R1858 VDD2.n89 VDD2.n88 104.615
R1859 VDD2.n22 VDD2.n21 104.615
R1860 VDD2.n22 VDD2.n15 104.615
R1861 VDD2.n29 VDD2.n15 104.615
R1862 VDD2.n30 VDD2.n29 104.615
R1863 VDD2.n30 VDD2.n11 104.615
R1864 VDD2.n38 VDD2.n11 104.615
R1865 VDD2.n39 VDD2.n38 104.615
R1866 VDD2.n40 VDD2.n39 104.615
R1867 VDD2.n40 VDD2.n7 104.615
R1868 VDD2.n47 VDD2.n7 104.615
R1869 VDD2.n48 VDD2.n47 104.615
R1870 VDD2.n48 VDD2.n3 104.615
R1871 VDD2.n55 VDD2.n3 104.615
R1872 VDD2.n56 VDD2.n55 104.615
R1873 VDD2.n64 VDD2.n63 60.5346
R1874 VDD2 VDD2.n129 60.5318
R1875 VDD2.n128 VDD2.n127 60.1505
R1876 VDD2.n62 VDD2.n61 60.1503
R1877 VDD2.n88 VDD2.t2 52.3082
R1878 VDD2.n21 VDD2.t9 52.3082
R1879 VDD2.n62 VDD2.n60 47.5109
R1880 VDD2.n126 VDD2.n125 46.9247
R1881 VDD2.n126 VDD2.n64 36.2412
R1882 VDD2.n75 VDD2.n73 13.1884
R1883 VDD2.n41 VDD2.n8 13.1884
R1884 VDD2.n111 VDD2.n110 12.8005
R1885 VDD2.n107 VDD2.n106 12.8005
R1886 VDD2.n42 VDD2.n10 12.8005
R1887 VDD2.n46 VDD2.n45 12.8005
R1888 VDD2.n114 VDD2.n71 12.0247
R1889 VDD2.n103 VDD2.n76 12.0247
R1890 VDD2.n37 VDD2.n36 12.0247
R1891 VDD2.n49 VDD2.n6 12.0247
R1892 VDD2.n115 VDD2.n69 11.249
R1893 VDD2.n102 VDD2.n79 11.249
R1894 VDD2.n35 VDD2.n12 11.249
R1895 VDD2.n50 VDD2.n4 11.249
R1896 VDD2.n119 VDD2.n118 10.4732
R1897 VDD2.n99 VDD2.n98 10.4732
R1898 VDD2.n32 VDD2.n31 10.4732
R1899 VDD2.n54 VDD2.n53 10.4732
R1900 VDD2.n87 VDD2.n86 10.2747
R1901 VDD2.n20 VDD2.n19 10.2747
R1902 VDD2.n122 VDD2.n67 9.69747
R1903 VDD2.n95 VDD2.n81 9.69747
R1904 VDD2.n28 VDD2.n14 9.69747
R1905 VDD2.n57 VDD2.n2 9.69747
R1906 VDD2.n125 VDD2.n124 9.45567
R1907 VDD2.n60 VDD2.n59 9.45567
R1908 VDD2.n85 VDD2.n84 9.3005
R1909 VDD2.n92 VDD2.n91 9.3005
R1910 VDD2.n94 VDD2.n93 9.3005
R1911 VDD2.n81 VDD2.n80 9.3005
R1912 VDD2.n100 VDD2.n99 9.3005
R1913 VDD2.n102 VDD2.n101 9.3005
R1914 VDD2.n76 VDD2.n74 9.3005
R1915 VDD2.n108 VDD2.n107 9.3005
R1916 VDD2.n124 VDD2.n123 9.3005
R1917 VDD2.n67 VDD2.n66 9.3005
R1918 VDD2.n118 VDD2.n117 9.3005
R1919 VDD2.n116 VDD2.n115 9.3005
R1920 VDD2.n71 VDD2.n70 9.3005
R1921 VDD2.n110 VDD2.n109 9.3005
R1922 VDD2.n59 VDD2.n58 9.3005
R1923 VDD2.n2 VDD2.n1 9.3005
R1924 VDD2.n53 VDD2.n52 9.3005
R1925 VDD2.n51 VDD2.n50 9.3005
R1926 VDD2.n6 VDD2.n5 9.3005
R1927 VDD2.n45 VDD2.n44 9.3005
R1928 VDD2.n18 VDD2.n17 9.3005
R1929 VDD2.n25 VDD2.n24 9.3005
R1930 VDD2.n27 VDD2.n26 9.3005
R1931 VDD2.n14 VDD2.n13 9.3005
R1932 VDD2.n33 VDD2.n32 9.3005
R1933 VDD2.n35 VDD2.n34 9.3005
R1934 VDD2.n36 VDD2.n9 9.3005
R1935 VDD2.n43 VDD2.n42 9.3005
R1936 VDD2.n123 VDD2.n65 8.92171
R1937 VDD2.n94 VDD2.n83 8.92171
R1938 VDD2.n27 VDD2.n16 8.92171
R1939 VDD2.n58 VDD2.n0 8.92171
R1940 VDD2.n91 VDD2.n90 8.14595
R1941 VDD2.n24 VDD2.n23 8.14595
R1942 VDD2.n87 VDD2.n85 7.3702
R1943 VDD2.n20 VDD2.n18 7.3702
R1944 VDD2.n90 VDD2.n85 5.81868
R1945 VDD2.n23 VDD2.n18 5.81868
R1946 VDD2.n125 VDD2.n65 5.04292
R1947 VDD2.n91 VDD2.n83 5.04292
R1948 VDD2.n24 VDD2.n16 5.04292
R1949 VDD2.n60 VDD2.n0 5.04292
R1950 VDD2.n123 VDD2.n122 4.26717
R1951 VDD2.n95 VDD2.n94 4.26717
R1952 VDD2.n28 VDD2.n27 4.26717
R1953 VDD2.n58 VDD2.n57 4.26717
R1954 VDD2.n119 VDD2.n67 3.49141
R1955 VDD2.n98 VDD2.n81 3.49141
R1956 VDD2.n31 VDD2.n14 3.49141
R1957 VDD2.n54 VDD2.n2 3.49141
R1958 VDD2.n86 VDD2.n84 2.84303
R1959 VDD2.n19 VDD2.n17 2.84303
R1960 VDD2.n118 VDD2.n69 2.71565
R1961 VDD2.n99 VDD2.n79 2.71565
R1962 VDD2.n32 VDD2.n12 2.71565
R1963 VDD2.n53 VDD2.n4 2.71565
R1964 VDD2.n115 VDD2.n114 1.93989
R1965 VDD2.n103 VDD2.n102 1.93989
R1966 VDD2.n37 VDD2.n35 1.93989
R1967 VDD2.n50 VDD2.n49 1.93989
R1968 VDD2.n129 VDD2.t6 1.75271
R1969 VDD2.n129 VDD2.t7 1.75271
R1970 VDD2.n127 VDD2.t3 1.75271
R1971 VDD2.n127 VDD2.t1 1.75271
R1972 VDD2.n63 VDD2.t8 1.75271
R1973 VDD2.n63 VDD2.t5 1.75271
R1974 VDD2.n61 VDD2.t4 1.75271
R1975 VDD2.n61 VDD2.t0 1.75271
R1976 VDD2.n111 VDD2.n71 1.16414
R1977 VDD2.n106 VDD2.n76 1.16414
R1978 VDD2.n36 VDD2.n10 1.16414
R1979 VDD2.n46 VDD2.n6 1.16414
R1980 VDD2.n128 VDD2.n126 0.586707
R1981 VDD2.n110 VDD2.n73 0.388379
R1982 VDD2.n107 VDD2.n75 0.388379
R1983 VDD2.n42 VDD2.n41 0.388379
R1984 VDD2.n45 VDD2.n8 0.388379
R1985 VDD2 VDD2.n128 0.205241
R1986 VDD2.n124 VDD2.n66 0.155672
R1987 VDD2.n117 VDD2.n66 0.155672
R1988 VDD2.n117 VDD2.n116 0.155672
R1989 VDD2.n116 VDD2.n70 0.155672
R1990 VDD2.n109 VDD2.n70 0.155672
R1991 VDD2.n109 VDD2.n108 0.155672
R1992 VDD2.n108 VDD2.n74 0.155672
R1993 VDD2.n101 VDD2.n74 0.155672
R1994 VDD2.n101 VDD2.n100 0.155672
R1995 VDD2.n100 VDD2.n80 0.155672
R1996 VDD2.n93 VDD2.n80 0.155672
R1997 VDD2.n93 VDD2.n92 0.155672
R1998 VDD2.n92 VDD2.n84 0.155672
R1999 VDD2.n25 VDD2.n17 0.155672
R2000 VDD2.n26 VDD2.n25 0.155672
R2001 VDD2.n26 VDD2.n13 0.155672
R2002 VDD2.n33 VDD2.n13 0.155672
R2003 VDD2.n34 VDD2.n33 0.155672
R2004 VDD2.n34 VDD2.n9 0.155672
R2005 VDD2.n43 VDD2.n9 0.155672
R2006 VDD2.n44 VDD2.n43 0.155672
R2007 VDD2.n44 VDD2.n5 0.155672
R2008 VDD2.n51 VDD2.n5 0.155672
R2009 VDD2.n52 VDD2.n51 0.155672
R2010 VDD2.n52 VDD2.n1 0.155672
R2011 VDD2.n59 VDD2.n1 0.155672
R2012 VDD2.n64 VDD2.n62 0.0917057
C0 VDD2 VTAIL 18.5186f
C1 VP VTAIL 3.85678f
C2 VDD1 VN 0.147725f
C3 VDD1 VTAIL 18.4878f
C4 VDD2 VP 0.296508f
C5 VN VTAIL 3.84208f
C6 VDD2 VDD1 0.755033f
C7 VDD1 VP 4.31779f
C8 VDD2 VN 4.17384f
C9 VP VN 4.95088f
C10 VDD2 B 4.46696f
C11 VDD1 B 4.336209f
C12 VTAIL B 5.876557f
C13 VN B 7.91159f
C14 VP B 5.766004f
C15 VDD2.n0 B 0.037499f
C16 VDD2.n1 B 0.0286f
C17 VDD2.n2 B 0.015368f
C18 VDD2.n3 B 0.036326f
C19 VDD2.n4 B 0.016272f
C20 VDD2.n5 B 0.0286f
C21 VDD2.n6 B 0.015368f
C22 VDD2.n7 B 0.036326f
C23 VDD2.n8 B 0.015821f
C24 VDD2.n9 B 0.0286f
C25 VDD2.n10 B 0.016272f
C26 VDD2.n11 B 0.036326f
C27 VDD2.n12 B 0.016272f
C28 VDD2.n13 B 0.0286f
C29 VDD2.n14 B 0.015368f
C30 VDD2.n15 B 0.036326f
C31 VDD2.n16 B 0.016272f
C32 VDD2.n17 B 1.35378f
C33 VDD2.n18 B 0.015368f
C34 VDD2.t9 B 0.061244f
C35 VDD2.n19 B 0.198518f
C36 VDD2.n20 B 0.025679f
C37 VDD2.n21 B 0.027244f
C38 VDD2.n22 B 0.036326f
C39 VDD2.n23 B 0.016272f
C40 VDD2.n24 B 0.015368f
C41 VDD2.n25 B 0.0286f
C42 VDD2.n26 B 0.0286f
C43 VDD2.n27 B 0.015368f
C44 VDD2.n28 B 0.016272f
C45 VDD2.n29 B 0.036326f
C46 VDD2.n30 B 0.036326f
C47 VDD2.n31 B 0.016272f
C48 VDD2.n32 B 0.015368f
C49 VDD2.n33 B 0.0286f
C50 VDD2.n34 B 0.0286f
C51 VDD2.n35 B 0.015368f
C52 VDD2.n36 B 0.015368f
C53 VDD2.n37 B 0.016272f
C54 VDD2.n38 B 0.036326f
C55 VDD2.n39 B 0.036326f
C56 VDD2.n40 B 0.036326f
C57 VDD2.n41 B 0.015821f
C58 VDD2.n42 B 0.015368f
C59 VDD2.n43 B 0.0286f
C60 VDD2.n44 B 0.0286f
C61 VDD2.n45 B 0.015368f
C62 VDD2.n46 B 0.016272f
C63 VDD2.n47 B 0.036326f
C64 VDD2.n48 B 0.036326f
C65 VDD2.n49 B 0.016272f
C66 VDD2.n50 B 0.015368f
C67 VDD2.n51 B 0.0286f
C68 VDD2.n52 B 0.0286f
C69 VDD2.n53 B 0.015368f
C70 VDD2.n54 B 0.016272f
C71 VDD2.n55 B 0.036326f
C72 VDD2.n56 B 0.073861f
C73 VDD2.n57 B 0.016272f
C74 VDD2.n58 B 0.015368f
C75 VDD2.n59 B 0.062201f
C76 VDD2.n60 B 0.061813f
C77 VDD2.t4 B 0.255388f
C78 VDD2.t0 B 0.255388f
C79 VDD2.n61 B 2.26465f
C80 VDD2.n62 B 0.413425f
C81 VDD2.t8 B 0.255388f
C82 VDD2.t5 B 0.255388f
C83 VDD2.n63 B 2.26681f
C84 VDD2.n64 B 1.91529f
C85 VDD2.n65 B 0.037499f
C86 VDD2.n66 B 0.0286f
C87 VDD2.n67 B 0.015368f
C88 VDD2.n68 B 0.036326f
C89 VDD2.n69 B 0.016272f
C90 VDD2.n70 B 0.0286f
C91 VDD2.n71 B 0.015368f
C92 VDD2.n72 B 0.036326f
C93 VDD2.n73 B 0.015821f
C94 VDD2.n74 B 0.0286f
C95 VDD2.n75 B 0.015821f
C96 VDD2.n76 B 0.015368f
C97 VDD2.n77 B 0.036326f
C98 VDD2.n78 B 0.036326f
C99 VDD2.n79 B 0.016272f
C100 VDD2.n80 B 0.0286f
C101 VDD2.n81 B 0.015368f
C102 VDD2.n82 B 0.036326f
C103 VDD2.n83 B 0.016272f
C104 VDD2.n84 B 1.35378f
C105 VDD2.n85 B 0.015368f
C106 VDD2.t2 B 0.061244f
C107 VDD2.n86 B 0.198518f
C108 VDD2.n87 B 0.025679f
C109 VDD2.n88 B 0.027244f
C110 VDD2.n89 B 0.036326f
C111 VDD2.n90 B 0.016272f
C112 VDD2.n91 B 0.015368f
C113 VDD2.n92 B 0.0286f
C114 VDD2.n93 B 0.0286f
C115 VDD2.n94 B 0.015368f
C116 VDD2.n95 B 0.016272f
C117 VDD2.n96 B 0.036326f
C118 VDD2.n97 B 0.036326f
C119 VDD2.n98 B 0.016272f
C120 VDD2.n99 B 0.015368f
C121 VDD2.n100 B 0.0286f
C122 VDD2.n101 B 0.0286f
C123 VDD2.n102 B 0.015368f
C124 VDD2.n103 B 0.016272f
C125 VDD2.n104 B 0.036326f
C126 VDD2.n105 B 0.036326f
C127 VDD2.n106 B 0.016272f
C128 VDD2.n107 B 0.015368f
C129 VDD2.n108 B 0.0286f
C130 VDD2.n109 B 0.0286f
C131 VDD2.n110 B 0.015368f
C132 VDD2.n111 B 0.016272f
C133 VDD2.n112 B 0.036326f
C134 VDD2.n113 B 0.036326f
C135 VDD2.n114 B 0.016272f
C136 VDD2.n115 B 0.015368f
C137 VDD2.n116 B 0.0286f
C138 VDD2.n117 B 0.0286f
C139 VDD2.n118 B 0.015368f
C140 VDD2.n119 B 0.016272f
C141 VDD2.n120 B 0.036326f
C142 VDD2.n121 B 0.073861f
C143 VDD2.n122 B 0.016272f
C144 VDD2.n123 B 0.015368f
C145 VDD2.n124 B 0.062201f
C146 VDD2.n125 B 0.060495f
C147 VDD2.n126 B 2.24606f
C148 VDD2.t3 B 0.255388f
C149 VDD2.t1 B 0.255388f
C150 VDD2.n127 B 2.26466f
C151 VDD2.n128 B 0.311068f
C152 VDD2.t6 B 0.255388f
C153 VDD2.t7 B 0.255388f
C154 VDD2.n129 B 2.26678f
C155 VN.n0 B 0.052091f
C156 VN.n1 B 0.011821f
C157 VN.t0 B 0.595426f
C158 VN.t5 B 0.588434f
C159 VN.n2 B 0.236614f
C160 VN.n3 B 0.242649f
C161 VN.n4 B 0.122406f
C162 VN.n5 B 0.052091f
C163 VN.t9 B 0.588434f
C164 VN.n6 B 0.253895f
C165 VN.n7 B 0.011821f
C166 VN.t1 B 0.588434f
C167 VN.n8 B 0.236614f
C168 VN.t4 B 0.595426f
C169 VN.n9 B 0.242567f
C170 VN.n10 B 0.040368f
C171 VN.n11 B 0.052091f
C172 VN.t7 B 0.595426f
C173 VN.n12 B 0.011821f
C174 VN.t8 B 0.588434f
C175 VN.t3 B 0.588434f
C176 VN.n13 B 0.236614f
C177 VN.t2 B 0.595426f
C178 VN.n14 B 0.242649f
C179 VN.n15 B 0.122406f
C180 VN.n16 B 0.052091f
C181 VN.n17 B 0.253895f
C182 VN.n18 B 0.011821f
C183 VN.t6 B 0.588434f
C184 VN.n19 B 0.236614f
C185 VN.n20 B 0.242567f
C186 VN.n21 B 2.05588f
C187 VDD1.n0 B 0.037489f
C188 VDD1.n1 B 0.028593f
C189 VDD1.n2 B 0.015365f
C190 VDD1.n3 B 0.036317f
C191 VDD1.n4 B 0.016268f
C192 VDD1.n5 B 0.028593f
C193 VDD1.n6 B 0.015365f
C194 VDD1.n7 B 0.036317f
C195 VDD1.n8 B 0.015817f
C196 VDD1.n9 B 0.028593f
C197 VDD1.n10 B 0.015817f
C198 VDD1.n11 B 0.015365f
C199 VDD1.n12 B 0.036317f
C200 VDD1.n13 B 0.036317f
C201 VDD1.n14 B 0.016268f
C202 VDD1.n15 B 0.028593f
C203 VDD1.n16 B 0.015365f
C204 VDD1.n17 B 0.036317f
C205 VDD1.n18 B 0.016268f
C206 VDD1.n19 B 1.35345f
C207 VDD1.n20 B 0.015365f
C208 VDD1.t0 B 0.061229f
C209 VDD1.n21 B 0.198469f
C210 VDD1.n22 B 0.025673f
C211 VDD1.n23 B 0.027237f
C212 VDD1.n24 B 0.036317f
C213 VDD1.n25 B 0.016268f
C214 VDD1.n26 B 0.015365f
C215 VDD1.n27 B 0.028593f
C216 VDD1.n28 B 0.028593f
C217 VDD1.n29 B 0.015365f
C218 VDD1.n30 B 0.016268f
C219 VDD1.n31 B 0.036317f
C220 VDD1.n32 B 0.036317f
C221 VDD1.n33 B 0.016268f
C222 VDD1.n34 B 0.015365f
C223 VDD1.n35 B 0.028593f
C224 VDD1.n36 B 0.028593f
C225 VDD1.n37 B 0.015365f
C226 VDD1.n38 B 0.016268f
C227 VDD1.n39 B 0.036317f
C228 VDD1.n40 B 0.036317f
C229 VDD1.n41 B 0.016268f
C230 VDD1.n42 B 0.015365f
C231 VDD1.n43 B 0.028593f
C232 VDD1.n44 B 0.028593f
C233 VDD1.n45 B 0.015365f
C234 VDD1.n46 B 0.016268f
C235 VDD1.n47 B 0.036317f
C236 VDD1.n48 B 0.036317f
C237 VDD1.n49 B 0.016268f
C238 VDD1.n50 B 0.015365f
C239 VDD1.n51 B 0.028593f
C240 VDD1.n52 B 0.028593f
C241 VDD1.n53 B 0.015365f
C242 VDD1.n54 B 0.016268f
C243 VDD1.n55 B 0.036317f
C244 VDD1.n56 B 0.073843f
C245 VDD1.n57 B 0.016268f
C246 VDD1.n58 B 0.015365f
C247 VDD1.n59 B 0.062186f
C248 VDD1.n60 B 0.061798f
C249 VDD1.t1 B 0.255325f
C250 VDD1.t2 B 0.255325f
C251 VDD1.n61 B 2.2641f
C252 VDD1.n62 B 0.416506f
C253 VDD1.n63 B 0.037489f
C254 VDD1.n64 B 0.028593f
C255 VDD1.n65 B 0.015365f
C256 VDD1.n66 B 0.036317f
C257 VDD1.n67 B 0.016268f
C258 VDD1.n68 B 0.028593f
C259 VDD1.n69 B 0.015365f
C260 VDD1.n70 B 0.036317f
C261 VDD1.n71 B 0.015817f
C262 VDD1.n72 B 0.028593f
C263 VDD1.n73 B 0.016268f
C264 VDD1.n74 B 0.036317f
C265 VDD1.n75 B 0.016268f
C266 VDD1.n76 B 0.028593f
C267 VDD1.n77 B 0.015365f
C268 VDD1.n78 B 0.036317f
C269 VDD1.n79 B 0.016268f
C270 VDD1.n80 B 1.35345f
C271 VDD1.n81 B 0.015365f
C272 VDD1.t4 B 0.061229f
C273 VDD1.n82 B 0.198469f
C274 VDD1.n83 B 0.025673f
C275 VDD1.n84 B 0.027237f
C276 VDD1.n85 B 0.036317f
C277 VDD1.n86 B 0.016268f
C278 VDD1.n87 B 0.015365f
C279 VDD1.n88 B 0.028593f
C280 VDD1.n89 B 0.028593f
C281 VDD1.n90 B 0.015365f
C282 VDD1.n91 B 0.016268f
C283 VDD1.n92 B 0.036317f
C284 VDD1.n93 B 0.036317f
C285 VDD1.n94 B 0.016268f
C286 VDD1.n95 B 0.015365f
C287 VDD1.n96 B 0.028593f
C288 VDD1.n97 B 0.028593f
C289 VDD1.n98 B 0.015365f
C290 VDD1.n99 B 0.015365f
C291 VDD1.n100 B 0.016268f
C292 VDD1.n101 B 0.036317f
C293 VDD1.n102 B 0.036317f
C294 VDD1.n103 B 0.036317f
C295 VDD1.n104 B 0.015817f
C296 VDD1.n105 B 0.015365f
C297 VDD1.n106 B 0.028593f
C298 VDD1.n107 B 0.028593f
C299 VDD1.n108 B 0.015365f
C300 VDD1.n109 B 0.016268f
C301 VDD1.n110 B 0.036317f
C302 VDD1.n111 B 0.036317f
C303 VDD1.n112 B 0.016268f
C304 VDD1.n113 B 0.015365f
C305 VDD1.n114 B 0.028593f
C306 VDD1.n115 B 0.028593f
C307 VDD1.n116 B 0.015365f
C308 VDD1.n117 B 0.016268f
C309 VDD1.n118 B 0.036317f
C310 VDD1.n119 B 0.073843f
C311 VDD1.n120 B 0.016268f
C312 VDD1.n121 B 0.015365f
C313 VDD1.n122 B 0.062186f
C314 VDD1.n123 B 0.061798f
C315 VDD1.t5 B 0.255325f
C316 VDD1.t7 B 0.255325f
C317 VDD1.n124 B 2.26409f
C318 VDD1.n125 B 0.413323f
C319 VDD1.t3 B 0.255325f
C320 VDD1.t6 B 0.255325f
C321 VDD1.n126 B 2.26625f
C322 VDD1.n127 B 1.9935f
C323 VDD1.t8 B 0.255325f
C324 VDD1.t9 B 0.255325f
C325 VDD1.n128 B 2.26409f
C326 VDD1.n129 B 2.50439f
C327 VTAIL.t6 B 0.265149f
C328 VTAIL.t1 B 0.265149f
C329 VTAIL.n0 B 2.25849f
C330 VTAIL.n1 B 0.42027f
C331 VTAIL.n2 B 0.038932f
C332 VTAIL.n3 B 0.029693f
C333 VTAIL.n4 B 0.015956f
C334 VTAIL.n5 B 0.037714f
C335 VTAIL.n6 B 0.016895f
C336 VTAIL.n7 B 0.029693f
C337 VTAIL.n8 B 0.015956f
C338 VTAIL.n9 B 0.037714f
C339 VTAIL.n10 B 0.016425f
C340 VTAIL.n11 B 0.029693f
C341 VTAIL.n12 B 0.016895f
C342 VTAIL.n13 B 0.037714f
C343 VTAIL.n14 B 0.016895f
C344 VTAIL.n15 B 0.029693f
C345 VTAIL.n16 B 0.015956f
C346 VTAIL.n17 B 0.037714f
C347 VTAIL.n18 B 0.016895f
C348 VTAIL.n19 B 1.40553f
C349 VTAIL.n20 B 0.015956f
C350 VTAIL.t11 B 0.063585f
C351 VTAIL.n21 B 0.206106f
C352 VTAIL.n22 B 0.026661f
C353 VTAIL.n23 B 0.028285f
C354 VTAIL.n24 B 0.037714f
C355 VTAIL.n25 B 0.016895f
C356 VTAIL.n26 B 0.015956f
C357 VTAIL.n27 B 0.029693f
C358 VTAIL.n28 B 0.029693f
C359 VTAIL.n29 B 0.015956f
C360 VTAIL.n30 B 0.016895f
C361 VTAIL.n31 B 0.037714f
C362 VTAIL.n32 B 0.037714f
C363 VTAIL.n33 B 0.016895f
C364 VTAIL.n34 B 0.015956f
C365 VTAIL.n35 B 0.029693f
C366 VTAIL.n36 B 0.029693f
C367 VTAIL.n37 B 0.015956f
C368 VTAIL.n38 B 0.015956f
C369 VTAIL.n39 B 0.016895f
C370 VTAIL.n40 B 0.037714f
C371 VTAIL.n41 B 0.037714f
C372 VTAIL.n42 B 0.037714f
C373 VTAIL.n43 B 0.016425f
C374 VTAIL.n44 B 0.015956f
C375 VTAIL.n45 B 0.029693f
C376 VTAIL.n46 B 0.029693f
C377 VTAIL.n47 B 0.015956f
C378 VTAIL.n48 B 0.016895f
C379 VTAIL.n49 B 0.037714f
C380 VTAIL.n50 B 0.037714f
C381 VTAIL.n51 B 0.016895f
C382 VTAIL.n52 B 0.015956f
C383 VTAIL.n53 B 0.029693f
C384 VTAIL.n54 B 0.029693f
C385 VTAIL.n55 B 0.015956f
C386 VTAIL.n56 B 0.016895f
C387 VTAIL.n57 B 0.037714f
C388 VTAIL.n58 B 0.076684f
C389 VTAIL.n59 B 0.016895f
C390 VTAIL.n60 B 0.015956f
C391 VTAIL.n61 B 0.064578f
C392 VTAIL.n62 B 0.04227f
C393 VTAIL.n63 B 0.152158f
C394 VTAIL.t12 B 0.265149f
C395 VTAIL.t8 B 0.265149f
C396 VTAIL.n64 B 2.25849f
C397 VTAIL.n65 B 0.411816f
C398 VTAIL.t10 B 0.265149f
C399 VTAIL.t9 B 0.265149f
C400 VTAIL.n66 B 2.25849f
C401 VTAIL.n67 B 1.80329f
C402 VTAIL.t17 B 0.265149f
C403 VTAIL.t5 B 0.265149f
C404 VTAIL.n68 B 2.25851f
C405 VTAIL.n69 B 1.80328f
C406 VTAIL.t18 B 0.265149f
C407 VTAIL.t4 B 0.265149f
C408 VTAIL.n70 B 2.25851f
C409 VTAIL.n71 B 0.411802f
C410 VTAIL.n72 B 0.038932f
C411 VTAIL.n73 B 0.029693f
C412 VTAIL.n74 B 0.015956f
C413 VTAIL.n75 B 0.037714f
C414 VTAIL.n76 B 0.016895f
C415 VTAIL.n77 B 0.029693f
C416 VTAIL.n78 B 0.015956f
C417 VTAIL.n79 B 0.037714f
C418 VTAIL.n80 B 0.016425f
C419 VTAIL.n81 B 0.029693f
C420 VTAIL.n82 B 0.016425f
C421 VTAIL.n83 B 0.015956f
C422 VTAIL.n84 B 0.037714f
C423 VTAIL.n85 B 0.037714f
C424 VTAIL.n86 B 0.016895f
C425 VTAIL.n87 B 0.029693f
C426 VTAIL.n88 B 0.015956f
C427 VTAIL.n89 B 0.037714f
C428 VTAIL.n90 B 0.016895f
C429 VTAIL.n91 B 1.40553f
C430 VTAIL.n92 B 0.015956f
C431 VTAIL.t3 B 0.063585f
C432 VTAIL.n93 B 0.206106f
C433 VTAIL.n94 B 0.026661f
C434 VTAIL.n95 B 0.028285f
C435 VTAIL.n96 B 0.037714f
C436 VTAIL.n97 B 0.016895f
C437 VTAIL.n98 B 0.015956f
C438 VTAIL.n99 B 0.029693f
C439 VTAIL.n100 B 0.029693f
C440 VTAIL.n101 B 0.015956f
C441 VTAIL.n102 B 0.016895f
C442 VTAIL.n103 B 0.037714f
C443 VTAIL.n104 B 0.037714f
C444 VTAIL.n105 B 0.016895f
C445 VTAIL.n106 B 0.015956f
C446 VTAIL.n107 B 0.029693f
C447 VTAIL.n108 B 0.029693f
C448 VTAIL.n109 B 0.015956f
C449 VTAIL.n110 B 0.016895f
C450 VTAIL.n111 B 0.037714f
C451 VTAIL.n112 B 0.037714f
C452 VTAIL.n113 B 0.016895f
C453 VTAIL.n114 B 0.015956f
C454 VTAIL.n115 B 0.029693f
C455 VTAIL.n116 B 0.029693f
C456 VTAIL.n117 B 0.015956f
C457 VTAIL.n118 B 0.016895f
C458 VTAIL.n119 B 0.037714f
C459 VTAIL.n120 B 0.037714f
C460 VTAIL.n121 B 0.016895f
C461 VTAIL.n122 B 0.015956f
C462 VTAIL.n123 B 0.029693f
C463 VTAIL.n124 B 0.029693f
C464 VTAIL.n125 B 0.015956f
C465 VTAIL.n126 B 0.016895f
C466 VTAIL.n127 B 0.037714f
C467 VTAIL.n128 B 0.076684f
C468 VTAIL.n129 B 0.016895f
C469 VTAIL.n130 B 0.015956f
C470 VTAIL.n131 B 0.064578f
C471 VTAIL.n132 B 0.04227f
C472 VTAIL.n133 B 0.152158f
C473 VTAIL.t16 B 0.265149f
C474 VTAIL.t7 B 0.265149f
C475 VTAIL.n134 B 2.25851f
C476 VTAIL.n135 B 0.428711f
C477 VTAIL.t15 B 0.265149f
C478 VTAIL.t13 B 0.265149f
C479 VTAIL.n136 B 2.25851f
C480 VTAIL.n137 B 0.411802f
C481 VTAIL.n138 B 0.038932f
C482 VTAIL.n139 B 0.029693f
C483 VTAIL.n140 B 0.015956f
C484 VTAIL.n141 B 0.037714f
C485 VTAIL.n142 B 0.016895f
C486 VTAIL.n143 B 0.029693f
C487 VTAIL.n144 B 0.015956f
C488 VTAIL.n145 B 0.037714f
C489 VTAIL.n146 B 0.016425f
C490 VTAIL.n147 B 0.029693f
C491 VTAIL.n148 B 0.016425f
C492 VTAIL.n149 B 0.015956f
C493 VTAIL.n150 B 0.037714f
C494 VTAIL.n151 B 0.037714f
C495 VTAIL.n152 B 0.016895f
C496 VTAIL.n153 B 0.029693f
C497 VTAIL.n154 B 0.015956f
C498 VTAIL.n155 B 0.037714f
C499 VTAIL.n156 B 0.016895f
C500 VTAIL.n157 B 1.40553f
C501 VTAIL.n158 B 0.015956f
C502 VTAIL.t14 B 0.063585f
C503 VTAIL.n159 B 0.206106f
C504 VTAIL.n160 B 0.026661f
C505 VTAIL.n161 B 0.028285f
C506 VTAIL.n162 B 0.037714f
C507 VTAIL.n163 B 0.016895f
C508 VTAIL.n164 B 0.015956f
C509 VTAIL.n165 B 0.029693f
C510 VTAIL.n166 B 0.029693f
C511 VTAIL.n167 B 0.015956f
C512 VTAIL.n168 B 0.016895f
C513 VTAIL.n169 B 0.037714f
C514 VTAIL.n170 B 0.037714f
C515 VTAIL.n171 B 0.016895f
C516 VTAIL.n172 B 0.015956f
C517 VTAIL.n173 B 0.029693f
C518 VTAIL.n174 B 0.029693f
C519 VTAIL.n175 B 0.015956f
C520 VTAIL.n176 B 0.016895f
C521 VTAIL.n177 B 0.037714f
C522 VTAIL.n178 B 0.037714f
C523 VTAIL.n179 B 0.016895f
C524 VTAIL.n180 B 0.015956f
C525 VTAIL.n181 B 0.029693f
C526 VTAIL.n182 B 0.029693f
C527 VTAIL.n183 B 0.015956f
C528 VTAIL.n184 B 0.016895f
C529 VTAIL.n185 B 0.037714f
C530 VTAIL.n186 B 0.037714f
C531 VTAIL.n187 B 0.016895f
C532 VTAIL.n188 B 0.015956f
C533 VTAIL.n189 B 0.029693f
C534 VTAIL.n190 B 0.029693f
C535 VTAIL.n191 B 0.015956f
C536 VTAIL.n192 B 0.016895f
C537 VTAIL.n193 B 0.037714f
C538 VTAIL.n194 B 0.076684f
C539 VTAIL.n195 B 0.016895f
C540 VTAIL.n196 B 0.015956f
C541 VTAIL.n197 B 0.064578f
C542 VTAIL.n198 B 0.04227f
C543 VTAIL.n199 B 1.47064f
C544 VTAIL.n200 B 0.038932f
C545 VTAIL.n201 B 0.029693f
C546 VTAIL.n202 B 0.015956f
C547 VTAIL.n203 B 0.037714f
C548 VTAIL.n204 B 0.016895f
C549 VTAIL.n205 B 0.029693f
C550 VTAIL.n206 B 0.015956f
C551 VTAIL.n207 B 0.037714f
C552 VTAIL.n208 B 0.016425f
C553 VTAIL.n209 B 0.029693f
C554 VTAIL.n210 B 0.016895f
C555 VTAIL.n211 B 0.037714f
C556 VTAIL.n212 B 0.016895f
C557 VTAIL.n213 B 0.029693f
C558 VTAIL.n214 B 0.015956f
C559 VTAIL.n215 B 0.037714f
C560 VTAIL.n216 B 0.016895f
C561 VTAIL.n217 B 1.40553f
C562 VTAIL.n218 B 0.015956f
C563 VTAIL.t0 B 0.063585f
C564 VTAIL.n219 B 0.206106f
C565 VTAIL.n220 B 0.026661f
C566 VTAIL.n221 B 0.028285f
C567 VTAIL.n222 B 0.037714f
C568 VTAIL.n223 B 0.016895f
C569 VTAIL.n224 B 0.015956f
C570 VTAIL.n225 B 0.029693f
C571 VTAIL.n226 B 0.029693f
C572 VTAIL.n227 B 0.015956f
C573 VTAIL.n228 B 0.016895f
C574 VTAIL.n229 B 0.037714f
C575 VTAIL.n230 B 0.037714f
C576 VTAIL.n231 B 0.016895f
C577 VTAIL.n232 B 0.015956f
C578 VTAIL.n233 B 0.029693f
C579 VTAIL.n234 B 0.029693f
C580 VTAIL.n235 B 0.015956f
C581 VTAIL.n236 B 0.015956f
C582 VTAIL.n237 B 0.016895f
C583 VTAIL.n238 B 0.037714f
C584 VTAIL.n239 B 0.037714f
C585 VTAIL.n240 B 0.037714f
C586 VTAIL.n241 B 0.016425f
C587 VTAIL.n242 B 0.015956f
C588 VTAIL.n243 B 0.029693f
C589 VTAIL.n244 B 0.029693f
C590 VTAIL.n245 B 0.015956f
C591 VTAIL.n246 B 0.016895f
C592 VTAIL.n247 B 0.037714f
C593 VTAIL.n248 B 0.037714f
C594 VTAIL.n249 B 0.016895f
C595 VTAIL.n250 B 0.015956f
C596 VTAIL.n251 B 0.029693f
C597 VTAIL.n252 B 0.029693f
C598 VTAIL.n253 B 0.015956f
C599 VTAIL.n254 B 0.016895f
C600 VTAIL.n255 B 0.037714f
C601 VTAIL.n256 B 0.076684f
C602 VTAIL.n257 B 0.016895f
C603 VTAIL.n258 B 0.015956f
C604 VTAIL.n259 B 0.064578f
C605 VTAIL.n260 B 0.04227f
C606 VTAIL.n261 B 1.47064f
C607 VTAIL.t19 B 0.265149f
C608 VTAIL.t2 B 0.265149f
C609 VTAIL.n262 B 2.25849f
C610 VTAIL.n263 B 0.364183f
C611 VP.n0 B 0.053192f
C612 VP.n1 B 0.01207f
C613 VP.n2 B 0.053192f
C614 VP.t1 B 0.600871f
C615 VP.t7 B 0.600871f
C616 VP.n3 B 0.053192f
C617 VP.t8 B 0.600871f
C618 VP.n4 B 0.241616f
C619 VP.t9 B 0.608011f
C620 VP.n5 B 0.247778f
C621 VP.n6 B 0.124993f
C622 VP.n7 B 0.01207f
C623 VP.n8 B 0.259261f
C624 VP.n9 B 0.01207f
C625 VP.n10 B 0.241616f
C626 VP.t0 B 0.608011f
C627 VP.n11 B 0.247694f
C628 VP.n12 B 2.06434f
C629 VP.t5 B 0.608011f
C630 VP.t4 B 0.600871f
C631 VP.n13 B 0.241616f
C632 VP.n14 B 0.247694f
C633 VP.n15 B 2.11142f
C634 VP.n16 B 0.053192f
C635 VP.n17 B 0.053192f
C636 VP.t2 B 0.600871f
C637 VP.n18 B 0.259261f
C638 VP.n19 B 0.01207f
C639 VP.t6 B 0.600871f
C640 VP.n20 B 0.241616f
C641 VP.t3 B 0.608011f
C642 VP.n21 B 0.247694f
C643 VP.n22 B 0.041222f
.ends

