* NGSPICE file created from diff_pair_sample_0260.ext - technology: sky130A

.subckt diff_pair_sample_0260 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0493 pd=12.75 as=4.8438 ps=25.62 w=12.42 l=3.29
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=0 ps=0 w=12.42 l=3.29
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=0 ps=0 w=12.42 l=3.29
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=0 ps=0 w=12.42 l=3.29
X4 VTAIL.t7 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=2.0493 ps=12.75 w=12.42 l=3.29
X5 VDD2.t3 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0493 pd=12.75 as=4.8438 ps=25.62 w=12.42 l=3.29
X6 VDD2.t2 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0493 pd=12.75 as=4.8438 ps=25.62 w=12.42 l=3.29
X7 VTAIL.t0 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=2.0493 ps=12.75 w=12.42 l=3.29
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=0 ps=0 w=12.42 l=3.29
X9 VDD1.t1 VP.t2 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0493 pd=12.75 as=4.8438 ps=25.62 w=12.42 l=3.29
X10 VTAIL.t6 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=2.0493 ps=12.75 w=12.42 l=3.29
X11 VTAIL.t1 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8438 pd=25.62 as=2.0493 ps=12.75 w=12.42 l=3.29
R0 VP.n17 VP.n16 161.3
R1 VP.n15 VP.n1 161.3
R2 VP.n14 VP.n13 161.3
R3 VP.n12 VP.n2 161.3
R4 VP.n11 VP.n10 161.3
R5 VP.n9 VP.n3 161.3
R6 VP.n8 VP.n7 161.3
R7 VP.n5 VP.t3 125.968
R8 VP.n5 VP.t0 124.85
R9 VP.n4 VP.t1 90.9798
R10 VP.n0 VP.t2 90.9798
R11 VP.n6 VP.n4 74.9986
R12 VP.n18 VP.n0 74.9986
R13 VP.n6 VP.n5 51.2992
R14 VP.n10 VP.n2 40.577
R15 VP.n14 VP.n2 40.577
R16 VP.n9 VP.n8 24.5923
R17 VP.n10 VP.n9 24.5923
R18 VP.n15 VP.n14 24.5923
R19 VP.n16 VP.n15 24.5923
R20 VP.n8 VP.n4 15.2474
R21 VP.n16 VP.n0 15.2474
R22 VP.n7 VP.n6 0.354861
R23 VP.n18 VP.n17 0.354861
R24 VP VP.n18 0.267071
R25 VP.n7 VP.n3 0.189894
R26 VP.n11 VP.n3 0.189894
R27 VP.n12 VP.n11 0.189894
R28 VP.n13 VP.n12 0.189894
R29 VP.n13 VP.n1 0.189894
R30 VP.n17 VP.n1 0.189894
R31 VTAIL.n5 VTAIL.t6 45.5393
R32 VTAIL.n4 VTAIL.t2 45.5393
R33 VTAIL.n3 VTAIL.t0 45.5393
R34 VTAIL.n7 VTAIL.t3 45.5391
R35 VTAIL.n0 VTAIL.t1 45.5391
R36 VTAIL.n1 VTAIL.t4 45.5391
R37 VTAIL.n2 VTAIL.t7 45.5391
R38 VTAIL.n6 VTAIL.t5 45.5391
R39 VTAIL.n7 VTAIL.n6 26.1945
R40 VTAIL.n3 VTAIL.n2 26.1945
R41 VTAIL.n4 VTAIL.n3 3.12119
R42 VTAIL.n6 VTAIL.n5 3.12119
R43 VTAIL.n2 VTAIL.n1 3.12119
R44 VTAIL VTAIL.n0 1.61903
R45 VTAIL VTAIL.n7 1.50266
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 VDD1 VDD1.n1 104.933
R49 VDD1 VDD1.n0 60.6819
R50 VDD1.n0 VDD1.t0 1.5947
R51 VDD1.n0 VDD1.t3 1.5947
R52 VDD1.n1 VDD1.t2 1.5947
R53 VDD1.n1 VDD1.t1 1.5947
R54 B.n808 B.n807 585
R55 B.n809 B.n808 585
R56 B.n314 B.n123 585
R57 B.n313 B.n312 585
R58 B.n311 B.n310 585
R59 B.n309 B.n308 585
R60 B.n307 B.n306 585
R61 B.n305 B.n304 585
R62 B.n303 B.n302 585
R63 B.n301 B.n300 585
R64 B.n299 B.n298 585
R65 B.n297 B.n296 585
R66 B.n295 B.n294 585
R67 B.n293 B.n292 585
R68 B.n291 B.n290 585
R69 B.n289 B.n288 585
R70 B.n287 B.n286 585
R71 B.n285 B.n284 585
R72 B.n283 B.n282 585
R73 B.n281 B.n280 585
R74 B.n279 B.n278 585
R75 B.n277 B.n276 585
R76 B.n275 B.n274 585
R77 B.n273 B.n272 585
R78 B.n271 B.n270 585
R79 B.n269 B.n268 585
R80 B.n267 B.n266 585
R81 B.n265 B.n264 585
R82 B.n263 B.n262 585
R83 B.n261 B.n260 585
R84 B.n259 B.n258 585
R85 B.n257 B.n256 585
R86 B.n255 B.n254 585
R87 B.n253 B.n252 585
R88 B.n251 B.n250 585
R89 B.n249 B.n248 585
R90 B.n247 B.n246 585
R91 B.n245 B.n244 585
R92 B.n243 B.n242 585
R93 B.n241 B.n240 585
R94 B.n239 B.n238 585
R95 B.n237 B.n236 585
R96 B.n235 B.n234 585
R97 B.n233 B.n232 585
R98 B.n231 B.n230 585
R99 B.n229 B.n228 585
R100 B.n227 B.n226 585
R101 B.n225 B.n224 585
R102 B.n223 B.n222 585
R103 B.n221 B.n220 585
R104 B.n219 B.n218 585
R105 B.n217 B.n216 585
R106 B.n215 B.n214 585
R107 B.n212 B.n211 585
R108 B.n210 B.n209 585
R109 B.n208 B.n207 585
R110 B.n206 B.n205 585
R111 B.n204 B.n203 585
R112 B.n202 B.n201 585
R113 B.n200 B.n199 585
R114 B.n198 B.n197 585
R115 B.n196 B.n195 585
R116 B.n194 B.n193 585
R117 B.n192 B.n191 585
R118 B.n190 B.n189 585
R119 B.n188 B.n187 585
R120 B.n186 B.n185 585
R121 B.n184 B.n183 585
R122 B.n182 B.n181 585
R123 B.n180 B.n179 585
R124 B.n178 B.n177 585
R125 B.n176 B.n175 585
R126 B.n174 B.n173 585
R127 B.n172 B.n171 585
R128 B.n170 B.n169 585
R129 B.n168 B.n167 585
R130 B.n166 B.n165 585
R131 B.n164 B.n163 585
R132 B.n162 B.n161 585
R133 B.n160 B.n159 585
R134 B.n158 B.n157 585
R135 B.n156 B.n155 585
R136 B.n154 B.n153 585
R137 B.n152 B.n151 585
R138 B.n150 B.n149 585
R139 B.n148 B.n147 585
R140 B.n146 B.n145 585
R141 B.n144 B.n143 585
R142 B.n142 B.n141 585
R143 B.n140 B.n139 585
R144 B.n138 B.n137 585
R145 B.n136 B.n135 585
R146 B.n134 B.n133 585
R147 B.n132 B.n131 585
R148 B.n130 B.n129 585
R149 B.n74 B.n73 585
R150 B.n806 B.n75 585
R151 B.n810 B.n75 585
R152 B.n805 B.n804 585
R153 B.n804 B.n71 585
R154 B.n803 B.n70 585
R155 B.n816 B.n70 585
R156 B.n802 B.n69 585
R157 B.n817 B.n69 585
R158 B.n801 B.n68 585
R159 B.n818 B.n68 585
R160 B.n800 B.n799 585
R161 B.n799 B.n64 585
R162 B.n798 B.n63 585
R163 B.n824 B.n63 585
R164 B.n797 B.n62 585
R165 B.n825 B.n62 585
R166 B.n796 B.n61 585
R167 B.n826 B.n61 585
R168 B.n795 B.n794 585
R169 B.n794 B.n57 585
R170 B.n793 B.n56 585
R171 B.n832 B.n56 585
R172 B.n792 B.n55 585
R173 B.n833 B.n55 585
R174 B.n791 B.n54 585
R175 B.n834 B.n54 585
R176 B.n790 B.n789 585
R177 B.n789 B.n50 585
R178 B.n788 B.n49 585
R179 B.n840 B.n49 585
R180 B.n787 B.n48 585
R181 B.n841 B.n48 585
R182 B.n786 B.n47 585
R183 B.n842 B.n47 585
R184 B.n785 B.n784 585
R185 B.n784 B.n43 585
R186 B.n783 B.n42 585
R187 B.n848 B.n42 585
R188 B.n782 B.n41 585
R189 B.n849 B.n41 585
R190 B.n781 B.n40 585
R191 B.n850 B.n40 585
R192 B.n780 B.n779 585
R193 B.n779 B.n36 585
R194 B.n778 B.n35 585
R195 B.n856 B.n35 585
R196 B.n777 B.n34 585
R197 B.n857 B.n34 585
R198 B.n776 B.n33 585
R199 B.n858 B.n33 585
R200 B.n775 B.n774 585
R201 B.n774 B.n29 585
R202 B.n773 B.n28 585
R203 B.n864 B.n28 585
R204 B.n772 B.n27 585
R205 B.n865 B.n27 585
R206 B.n771 B.n26 585
R207 B.n866 B.n26 585
R208 B.n770 B.n769 585
R209 B.n769 B.n22 585
R210 B.n768 B.n21 585
R211 B.n872 B.n21 585
R212 B.n767 B.n20 585
R213 B.n873 B.n20 585
R214 B.n766 B.n19 585
R215 B.n874 B.n19 585
R216 B.n765 B.n764 585
R217 B.n764 B.n18 585
R218 B.n763 B.n14 585
R219 B.n880 B.n14 585
R220 B.n762 B.n13 585
R221 B.n881 B.n13 585
R222 B.n761 B.n12 585
R223 B.n882 B.n12 585
R224 B.n760 B.n759 585
R225 B.n759 B.n8 585
R226 B.n758 B.n7 585
R227 B.n888 B.n7 585
R228 B.n757 B.n6 585
R229 B.n889 B.n6 585
R230 B.n756 B.n5 585
R231 B.n890 B.n5 585
R232 B.n755 B.n754 585
R233 B.n754 B.n4 585
R234 B.n753 B.n315 585
R235 B.n753 B.n752 585
R236 B.n743 B.n316 585
R237 B.n317 B.n316 585
R238 B.n745 B.n744 585
R239 B.n746 B.n745 585
R240 B.n742 B.n322 585
R241 B.n322 B.n321 585
R242 B.n741 B.n740 585
R243 B.n740 B.n739 585
R244 B.n324 B.n323 585
R245 B.n732 B.n324 585
R246 B.n731 B.n730 585
R247 B.n733 B.n731 585
R248 B.n729 B.n329 585
R249 B.n329 B.n328 585
R250 B.n728 B.n727 585
R251 B.n727 B.n726 585
R252 B.n331 B.n330 585
R253 B.n332 B.n331 585
R254 B.n719 B.n718 585
R255 B.n720 B.n719 585
R256 B.n717 B.n337 585
R257 B.n337 B.n336 585
R258 B.n716 B.n715 585
R259 B.n715 B.n714 585
R260 B.n339 B.n338 585
R261 B.n340 B.n339 585
R262 B.n707 B.n706 585
R263 B.n708 B.n707 585
R264 B.n705 B.n345 585
R265 B.n345 B.n344 585
R266 B.n704 B.n703 585
R267 B.n703 B.n702 585
R268 B.n347 B.n346 585
R269 B.n348 B.n347 585
R270 B.n695 B.n694 585
R271 B.n696 B.n695 585
R272 B.n693 B.n353 585
R273 B.n353 B.n352 585
R274 B.n692 B.n691 585
R275 B.n691 B.n690 585
R276 B.n355 B.n354 585
R277 B.n356 B.n355 585
R278 B.n683 B.n682 585
R279 B.n684 B.n683 585
R280 B.n681 B.n361 585
R281 B.n361 B.n360 585
R282 B.n680 B.n679 585
R283 B.n679 B.n678 585
R284 B.n363 B.n362 585
R285 B.n364 B.n363 585
R286 B.n671 B.n670 585
R287 B.n672 B.n671 585
R288 B.n669 B.n369 585
R289 B.n369 B.n368 585
R290 B.n668 B.n667 585
R291 B.n667 B.n666 585
R292 B.n371 B.n370 585
R293 B.n372 B.n371 585
R294 B.n659 B.n658 585
R295 B.n660 B.n659 585
R296 B.n657 B.n377 585
R297 B.n377 B.n376 585
R298 B.n656 B.n655 585
R299 B.n655 B.n654 585
R300 B.n379 B.n378 585
R301 B.n380 B.n379 585
R302 B.n647 B.n646 585
R303 B.n648 B.n647 585
R304 B.n645 B.n385 585
R305 B.n385 B.n384 585
R306 B.n644 B.n643 585
R307 B.n643 B.n642 585
R308 B.n387 B.n386 585
R309 B.n388 B.n387 585
R310 B.n635 B.n634 585
R311 B.n636 B.n635 585
R312 B.n391 B.n390 585
R313 B.n444 B.n443 585
R314 B.n445 B.n441 585
R315 B.n441 B.n392 585
R316 B.n447 B.n446 585
R317 B.n449 B.n440 585
R318 B.n452 B.n451 585
R319 B.n453 B.n439 585
R320 B.n455 B.n454 585
R321 B.n457 B.n438 585
R322 B.n460 B.n459 585
R323 B.n461 B.n437 585
R324 B.n463 B.n462 585
R325 B.n465 B.n436 585
R326 B.n468 B.n467 585
R327 B.n469 B.n435 585
R328 B.n471 B.n470 585
R329 B.n473 B.n434 585
R330 B.n476 B.n475 585
R331 B.n477 B.n433 585
R332 B.n479 B.n478 585
R333 B.n481 B.n432 585
R334 B.n484 B.n483 585
R335 B.n485 B.n431 585
R336 B.n487 B.n486 585
R337 B.n489 B.n430 585
R338 B.n492 B.n491 585
R339 B.n493 B.n429 585
R340 B.n495 B.n494 585
R341 B.n497 B.n428 585
R342 B.n500 B.n499 585
R343 B.n501 B.n427 585
R344 B.n503 B.n502 585
R345 B.n505 B.n426 585
R346 B.n508 B.n507 585
R347 B.n509 B.n425 585
R348 B.n511 B.n510 585
R349 B.n513 B.n424 585
R350 B.n516 B.n515 585
R351 B.n517 B.n423 585
R352 B.n519 B.n518 585
R353 B.n521 B.n422 585
R354 B.n524 B.n523 585
R355 B.n525 B.n419 585
R356 B.n528 B.n527 585
R357 B.n530 B.n418 585
R358 B.n533 B.n532 585
R359 B.n534 B.n417 585
R360 B.n536 B.n535 585
R361 B.n538 B.n416 585
R362 B.n541 B.n540 585
R363 B.n542 B.n415 585
R364 B.n547 B.n546 585
R365 B.n549 B.n414 585
R366 B.n552 B.n551 585
R367 B.n553 B.n413 585
R368 B.n555 B.n554 585
R369 B.n557 B.n412 585
R370 B.n560 B.n559 585
R371 B.n561 B.n411 585
R372 B.n563 B.n562 585
R373 B.n565 B.n410 585
R374 B.n568 B.n567 585
R375 B.n569 B.n409 585
R376 B.n571 B.n570 585
R377 B.n573 B.n408 585
R378 B.n576 B.n575 585
R379 B.n577 B.n407 585
R380 B.n579 B.n578 585
R381 B.n581 B.n406 585
R382 B.n584 B.n583 585
R383 B.n585 B.n405 585
R384 B.n587 B.n586 585
R385 B.n589 B.n404 585
R386 B.n592 B.n591 585
R387 B.n593 B.n403 585
R388 B.n595 B.n594 585
R389 B.n597 B.n402 585
R390 B.n600 B.n599 585
R391 B.n601 B.n401 585
R392 B.n603 B.n602 585
R393 B.n605 B.n400 585
R394 B.n608 B.n607 585
R395 B.n609 B.n399 585
R396 B.n611 B.n610 585
R397 B.n613 B.n398 585
R398 B.n616 B.n615 585
R399 B.n617 B.n397 585
R400 B.n619 B.n618 585
R401 B.n621 B.n396 585
R402 B.n624 B.n623 585
R403 B.n625 B.n395 585
R404 B.n627 B.n626 585
R405 B.n629 B.n394 585
R406 B.n632 B.n631 585
R407 B.n633 B.n393 585
R408 B.n638 B.n637 585
R409 B.n637 B.n636 585
R410 B.n639 B.n389 585
R411 B.n389 B.n388 585
R412 B.n641 B.n640 585
R413 B.n642 B.n641 585
R414 B.n383 B.n382 585
R415 B.n384 B.n383 585
R416 B.n650 B.n649 585
R417 B.n649 B.n648 585
R418 B.n651 B.n381 585
R419 B.n381 B.n380 585
R420 B.n653 B.n652 585
R421 B.n654 B.n653 585
R422 B.n375 B.n374 585
R423 B.n376 B.n375 585
R424 B.n662 B.n661 585
R425 B.n661 B.n660 585
R426 B.n663 B.n373 585
R427 B.n373 B.n372 585
R428 B.n665 B.n664 585
R429 B.n666 B.n665 585
R430 B.n367 B.n366 585
R431 B.n368 B.n367 585
R432 B.n674 B.n673 585
R433 B.n673 B.n672 585
R434 B.n675 B.n365 585
R435 B.n365 B.n364 585
R436 B.n677 B.n676 585
R437 B.n678 B.n677 585
R438 B.n359 B.n358 585
R439 B.n360 B.n359 585
R440 B.n686 B.n685 585
R441 B.n685 B.n684 585
R442 B.n687 B.n357 585
R443 B.n357 B.n356 585
R444 B.n689 B.n688 585
R445 B.n690 B.n689 585
R446 B.n351 B.n350 585
R447 B.n352 B.n351 585
R448 B.n698 B.n697 585
R449 B.n697 B.n696 585
R450 B.n699 B.n349 585
R451 B.n349 B.n348 585
R452 B.n701 B.n700 585
R453 B.n702 B.n701 585
R454 B.n343 B.n342 585
R455 B.n344 B.n343 585
R456 B.n710 B.n709 585
R457 B.n709 B.n708 585
R458 B.n711 B.n341 585
R459 B.n341 B.n340 585
R460 B.n713 B.n712 585
R461 B.n714 B.n713 585
R462 B.n335 B.n334 585
R463 B.n336 B.n335 585
R464 B.n722 B.n721 585
R465 B.n721 B.n720 585
R466 B.n723 B.n333 585
R467 B.n333 B.n332 585
R468 B.n725 B.n724 585
R469 B.n726 B.n725 585
R470 B.n327 B.n326 585
R471 B.n328 B.n327 585
R472 B.n735 B.n734 585
R473 B.n734 B.n733 585
R474 B.n736 B.n325 585
R475 B.n732 B.n325 585
R476 B.n738 B.n737 585
R477 B.n739 B.n738 585
R478 B.n320 B.n319 585
R479 B.n321 B.n320 585
R480 B.n748 B.n747 585
R481 B.n747 B.n746 585
R482 B.n749 B.n318 585
R483 B.n318 B.n317 585
R484 B.n751 B.n750 585
R485 B.n752 B.n751 585
R486 B.n2 B.n0 585
R487 B.n4 B.n2 585
R488 B.n3 B.n1 585
R489 B.n889 B.n3 585
R490 B.n887 B.n886 585
R491 B.n888 B.n887 585
R492 B.n885 B.n9 585
R493 B.n9 B.n8 585
R494 B.n884 B.n883 585
R495 B.n883 B.n882 585
R496 B.n11 B.n10 585
R497 B.n881 B.n11 585
R498 B.n879 B.n878 585
R499 B.n880 B.n879 585
R500 B.n877 B.n15 585
R501 B.n18 B.n15 585
R502 B.n876 B.n875 585
R503 B.n875 B.n874 585
R504 B.n17 B.n16 585
R505 B.n873 B.n17 585
R506 B.n871 B.n870 585
R507 B.n872 B.n871 585
R508 B.n869 B.n23 585
R509 B.n23 B.n22 585
R510 B.n868 B.n867 585
R511 B.n867 B.n866 585
R512 B.n25 B.n24 585
R513 B.n865 B.n25 585
R514 B.n863 B.n862 585
R515 B.n864 B.n863 585
R516 B.n861 B.n30 585
R517 B.n30 B.n29 585
R518 B.n860 B.n859 585
R519 B.n859 B.n858 585
R520 B.n32 B.n31 585
R521 B.n857 B.n32 585
R522 B.n855 B.n854 585
R523 B.n856 B.n855 585
R524 B.n853 B.n37 585
R525 B.n37 B.n36 585
R526 B.n852 B.n851 585
R527 B.n851 B.n850 585
R528 B.n39 B.n38 585
R529 B.n849 B.n39 585
R530 B.n847 B.n846 585
R531 B.n848 B.n847 585
R532 B.n845 B.n44 585
R533 B.n44 B.n43 585
R534 B.n844 B.n843 585
R535 B.n843 B.n842 585
R536 B.n46 B.n45 585
R537 B.n841 B.n46 585
R538 B.n839 B.n838 585
R539 B.n840 B.n839 585
R540 B.n837 B.n51 585
R541 B.n51 B.n50 585
R542 B.n836 B.n835 585
R543 B.n835 B.n834 585
R544 B.n53 B.n52 585
R545 B.n833 B.n53 585
R546 B.n831 B.n830 585
R547 B.n832 B.n831 585
R548 B.n829 B.n58 585
R549 B.n58 B.n57 585
R550 B.n828 B.n827 585
R551 B.n827 B.n826 585
R552 B.n60 B.n59 585
R553 B.n825 B.n60 585
R554 B.n823 B.n822 585
R555 B.n824 B.n823 585
R556 B.n821 B.n65 585
R557 B.n65 B.n64 585
R558 B.n820 B.n819 585
R559 B.n819 B.n818 585
R560 B.n67 B.n66 585
R561 B.n817 B.n67 585
R562 B.n815 B.n814 585
R563 B.n816 B.n815 585
R564 B.n813 B.n72 585
R565 B.n72 B.n71 585
R566 B.n812 B.n811 585
R567 B.n811 B.n810 585
R568 B.n892 B.n891 585
R569 B.n891 B.n890 585
R570 B.n637 B.n391 530.939
R571 B.n811 B.n74 530.939
R572 B.n635 B.n393 530.939
R573 B.n808 B.n75 530.939
R574 B.n543 B.t12 299.875
R575 B.n420 B.t4 299.875
R576 B.n127 B.t8 299.875
R577 B.n124 B.t15 299.875
R578 B.n809 B.n122 256.663
R579 B.n809 B.n121 256.663
R580 B.n809 B.n120 256.663
R581 B.n809 B.n119 256.663
R582 B.n809 B.n118 256.663
R583 B.n809 B.n117 256.663
R584 B.n809 B.n116 256.663
R585 B.n809 B.n115 256.663
R586 B.n809 B.n114 256.663
R587 B.n809 B.n113 256.663
R588 B.n809 B.n112 256.663
R589 B.n809 B.n111 256.663
R590 B.n809 B.n110 256.663
R591 B.n809 B.n109 256.663
R592 B.n809 B.n108 256.663
R593 B.n809 B.n107 256.663
R594 B.n809 B.n106 256.663
R595 B.n809 B.n105 256.663
R596 B.n809 B.n104 256.663
R597 B.n809 B.n103 256.663
R598 B.n809 B.n102 256.663
R599 B.n809 B.n101 256.663
R600 B.n809 B.n100 256.663
R601 B.n809 B.n99 256.663
R602 B.n809 B.n98 256.663
R603 B.n809 B.n97 256.663
R604 B.n809 B.n96 256.663
R605 B.n809 B.n95 256.663
R606 B.n809 B.n94 256.663
R607 B.n809 B.n93 256.663
R608 B.n809 B.n92 256.663
R609 B.n809 B.n91 256.663
R610 B.n809 B.n90 256.663
R611 B.n809 B.n89 256.663
R612 B.n809 B.n88 256.663
R613 B.n809 B.n87 256.663
R614 B.n809 B.n86 256.663
R615 B.n809 B.n85 256.663
R616 B.n809 B.n84 256.663
R617 B.n809 B.n83 256.663
R618 B.n809 B.n82 256.663
R619 B.n809 B.n81 256.663
R620 B.n809 B.n80 256.663
R621 B.n809 B.n79 256.663
R622 B.n809 B.n78 256.663
R623 B.n809 B.n77 256.663
R624 B.n809 B.n76 256.663
R625 B.n442 B.n392 256.663
R626 B.n448 B.n392 256.663
R627 B.n450 B.n392 256.663
R628 B.n456 B.n392 256.663
R629 B.n458 B.n392 256.663
R630 B.n464 B.n392 256.663
R631 B.n466 B.n392 256.663
R632 B.n472 B.n392 256.663
R633 B.n474 B.n392 256.663
R634 B.n480 B.n392 256.663
R635 B.n482 B.n392 256.663
R636 B.n488 B.n392 256.663
R637 B.n490 B.n392 256.663
R638 B.n496 B.n392 256.663
R639 B.n498 B.n392 256.663
R640 B.n504 B.n392 256.663
R641 B.n506 B.n392 256.663
R642 B.n512 B.n392 256.663
R643 B.n514 B.n392 256.663
R644 B.n520 B.n392 256.663
R645 B.n522 B.n392 256.663
R646 B.n529 B.n392 256.663
R647 B.n531 B.n392 256.663
R648 B.n537 B.n392 256.663
R649 B.n539 B.n392 256.663
R650 B.n548 B.n392 256.663
R651 B.n550 B.n392 256.663
R652 B.n556 B.n392 256.663
R653 B.n558 B.n392 256.663
R654 B.n564 B.n392 256.663
R655 B.n566 B.n392 256.663
R656 B.n572 B.n392 256.663
R657 B.n574 B.n392 256.663
R658 B.n580 B.n392 256.663
R659 B.n582 B.n392 256.663
R660 B.n588 B.n392 256.663
R661 B.n590 B.n392 256.663
R662 B.n596 B.n392 256.663
R663 B.n598 B.n392 256.663
R664 B.n604 B.n392 256.663
R665 B.n606 B.n392 256.663
R666 B.n612 B.n392 256.663
R667 B.n614 B.n392 256.663
R668 B.n620 B.n392 256.663
R669 B.n622 B.n392 256.663
R670 B.n628 B.n392 256.663
R671 B.n630 B.n392 256.663
R672 B.n637 B.n389 163.367
R673 B.n641 B.n389 163.367
R674 B.n641 B.n383 163.367
R675 B.n649 B.n383 163.367
R676 B.n649 B.n381 163.367
R677 B.n653 B.n381 163.367
R678 B.n653 B.n375 163.367
R679 B.n661 B.n375 163.367
R680 B.n661 B.n373 163.367
R681 B.n665 B.n373 163.367
R682 B.n665 B.n367 163.367
R683 B.n673 B.n367 163.367
R684 B.n673 B.n365 163.367
R685 B.n677 B.n365 163.367
R686 B.n677 B.n359 163.367
R687 B.n685 B.n359 163.367
R688 B.n685 B.n357 163.367
R689 B.n689 B.n357 163.367
R690 B.n689 B.n351 163.367
R691 B.n697 B.n351 163.367
R692 B.n697 B.n349 163.367
R693 B.n701 B.n349 163.367
R694 B.n701 B.n343 163.367
R695 B.n709 B.n343 163.367
R696 B.n709 B.n341 163.367
R697 B.n713 B.n341 163.367
R698 B.n713 B.n335 163.367
R699 B.n721 B.n335 163.367
R700 B.n721 B.n333 163.367
R701 B.n725 B.n333 163.367
R702 B.n725 B.n327 163.367
R703 B.n734 B.n327 163.367
R704 B.n734 B.n325 163.367
R705 B.n738 B.n325 163.367
R706 B.n738 B.n320 163.367
R707 B.n747 B.n320 163.367
R708 B.n747 B.n318 163.367
R709 B.n751 B.n318 163.367
R710 B.n751 B.n2 163.367
R711 B.n891 B.n2 163.367
R712 B.n891 B.n3 163.367
R713 B.n887 B.n3 163.367
R714 B.n887 B.n9 163.367
R715 B.n883 B.n9 163.367
R716 B.n883 B.n11 163.367
R717 B.n879 B.n11 163.367
R718 B.n879 B.n15 163.367
R719 B.n875 B.n15 163.367
R720 B.n875 B.n17 163.367
R721 B.n871 B.n17 163.367
R722 B.n871 B.n23 163.367
R723 B.n867 B.n23 163.367
R724 B.n867 B.n25 163.367
R725 B.n863 B.n25 163.367
R726 B.n863 B.n30 163.367
R727 B.n859 B.n30 163.367
R728 B.n859 B.n32 163.367
R729 B.n855 B.n32 163.367
R730 B.n855 B.n37 163.367
R731 B.n851 B.n37 163.367
R732 B.n851 B.n39 163.367
R733 B.n847 B.n39 163.367
R734 B.n847 B.n44 163.367
R735 B.n843 B.n44 163.367
R736 B.n843 B.n46 163.367
R737 B.n839 B.n46 163.367
R738 B.n839 B.n51 163.367
R739 B.n835 B.n51 163.367
R740 B.n835 B.n53 163.367
R741 B.n831 B.n53 163.367
R742 B.n831 B.n58 163.367
R743 B.n827 B.n58 163.367
R744 B.n827 B.n60 163.367
R745 B.n823 B.n60 163.367
R746 B.n823 B.n65 163.367
R747 B.n819 B.n65 163.367
R748 B.n819 B.n67 163.367
R749 B.n815 B.n67 163.367
R750 B.n815 B.n72 163.367
R751 B.n811 B.n72 163.367
R752 B.n443 B.n441 163.367
R753 B.n447 B.n441 163.367
R754 B.n451 B.n449 163.367
R755 B.n455 B.n439 163.367
R756 B.n459 B.n457 163.367
R757 B.n463 B.n437 163.367
R758 B.n467 B.n465 163.367
R759 B.n471 B.n435 163.367
R760 B.n475 B.n473 163.367
R761 B.n479 B.n433 163.367
R762 B.n483 B.n481 163.367
R763 B.n487 B.n431 163.367
R764 B.n491 B.n489 163.367
R765 B.n495 B.n429 163.367
R766 B.n499 B.n497 163.367
R767 B.n503 B.n427 163.367
R768 B.n507 B.n505 163.367
R769 B.n511 B.n425 163.367
R770 B.n515 B.n513 163.367
R771 B.n519 B.n423 163.367
R772 B.n523 B.n521 163.367
R773 B.n528 B.n419 163.367
R774 B.n532 B.n530 163.367
R775 B.n536 B.n417 163.367
R776 B.n540 B.n538 163.367
R777 B.n547 B.n415 163.367
R778 B.n551 B.n549 163.367
R779 B.n555 B.n413 163.367
R780 B.n559 B.n557 163.367
R781 B.n563 B.n411 163.367
R782 B.n567 B.n565 163.367
R783 B.n571 B.n409 163.367
R784 B.n575 B.n573 163.367
R785 B.n579 B.n407 163.367
R786 B.n583 B.n581 163.367
R787 B.n587 B.n405 163.367
R788 B.n591 B.n589 163.367
R789 B.n595 B.n403 163.367
R790 B.n599 B.n597 163.367
R791 B.n603 B.n401 163.367
R792 B.n607 B.n605 163.367
R793 B.n611 B.n399 163.367
R794 B.n615 B.n613 163.367
R795 B.n619 B.n397 163.367
R796 B.n623 B.n621 163.367
R797 B.n627 B.n395 163.367
R798 B.n631 B.n629 163.367
R799 B.n635 B.n387 163.367
R800 B.n643 B.n387 163.367
R801 B.n643 B.n385 163.367
R802 B.n647 B.n385 163.367
R803 B.n647 B.n379 163.367
R804 B.n655 B.n379 163.367
R805 B.n655 B.n377 163.367
R806 B.n659 B.n377 163.367
R807 B.n659 B.n371 163.367
R808 B.n667 B.n371 163.367
R809 B.n667 B.n369 163.367
R810 B.n671 B.n369 163.367
R811 B.n671 B.n363 163.367
R812 B.n679 B.n363 163.367
R813 B.n679 B.n361 163.367
R814 B.n683 B.n361 163.367
R815 B.n683 B.n355 163.367
R816 B.n691 B.n355 163.367
R817 B.n691 B.n353 163.367
R818 B.n695 B.n353 163.367
R819 B.n695 B.n347 163.367
R820 B.n703 B.n347 163.367
R821 B.n703 B.n345 163.367
R822 B.n707 B.n345 163.367
R823 B.n707 B.n339 163.367
R824 B.n715 B.n339 163.367
R825 B.n715 B.n337 163.367
R826 B.n719 B.n337 163.367
R827 B.n719 B.n331 163.367
R828 B.n727 B.n331 163.367
R829 B.n727 B.n329 163.367
R830 B.n731 B.n329 163.367
R831 B.n731 B.n324 163.367
R832 B.n740 B.n324 163.367
R833 B.n740 B.n322 163.367
R834 B.n745 B.n322 163.367
R835 B.n745 B.n316 163.367
R836 B.n753 B.n316 163.367
R837 B.n754 B.n753 163.367
R838 B.n754 B.n5 163.367
R839 B.n6 B.n5 163.367
R840 B.n7 B.n6 163.367
R841 B.n759 B.n7 163.367
R842 B.n759 B.n12 163.367
R843 B.n13 B.n12 163.367
R844 B.n14 B.n13 163.367
R845 B.n764 B.n14 163.367
R846 B.n764 B.n19 163.367
R847 B.n20 B.n19 163.367
R848 B.n21 B.n20 163.367
R849 B.n769 B.n21 163.367
R850 B.n769 B.n26 163.367
R851 B.n27 B.n26 163.367
R852 B.n28 B.n27 163.367
R853 B.n774 B.n28 163.367
R854 B.n774 B.n33 163.367
R855 B.n34 B.n33 163.367
R856 B.n35 B.n34 163.367
R857 B.n779 B.n35 163.367
R858 B.n779 B.n40 163.367
R859 B.n41 B.n40 163.367
R860 B.n42 B.n41 163.367
R861 B.n784 B.n42 163.367
R862 B.n784 B.n47 163.367
R863 B.n48 B.n47 163.367
R864 B.n49 B.n48 163.367
R865 B.n789 B.n49 163.367
R866 B.n789 B.n54 163.367
R867 B.n55 B.n54 163.367
R868 B.n56 B.n55 163.367
R869 B.n794 B.n56 163.367
R870 B.n794 B.n61 163.367
R871 B.n62 B.n61 163.367
R872 B.n63 B.n62 163.367
R873 B.n799 B.n63 163.367
R874 B.n799 B.n68 163.367
R875 B.n69 B.n68 163.367
R876 B.n70 B.n69 163.367
R877 B.n804 B.n70 163.367
R878 B.n804 B.n75 163.367
R879 B.n131 B.n130 163.367
R880 B.n135 B.n134 163.367
R881 B.n139 B.n138 163.367
R882 B.n143 B.n142 163.367
R883 B.n147 B.n146 163.367
R884 B.n151 B.n150 163.367
R885 B.n155 B.n154 163.367
R886 B.n159 B.n158 163.367
R887 B.n163 B.n162 163.367
R888 B.n167 B.n166 163.367
R889 B.n171 B.n170 163.367
R890 B.n175 B.n174 163.367
R891 B.n179 B.n178 163.367
R892 B.n183 B.n182 163.367
R893 B.n187 B.n186 163.367
R894 B.n191 B.n190 163.367
R895 B.n195 B.n194 163.367
R896 B.n199 B.n198 163.367
R897 B.n203 B.n202 163.367
R898 B.n207 B.n206 163.367
R899 B.n211 B.n210 163.367
R900 B.n216 B.n215 163.367
R901 B.n220 B.n219 163.367
R902 B.n224 B.n223 163.367
R903 B.n228 B.n227 163.367
R904 B.n232 B.n231 163.367
R905 B.n236 B.n235 163.367
R906 B.n240 B.n239 163.367
R907 B.n244 B.n243 163.367
R908 B.n248 B.n247 163.367
R909 B.n252 B.n251 163.367
R910 B.n256 B.n255 163.367
R911 B.n260 B.n259 163.367
R912 B.n264 B.n263 163.367
R913 B.n268 B.n267 163.367
R914 B.n272 B.n271 163.367
R915 B.n276 B.n275 163.367
R916 B.n280 B.n279 163.367
R917 B.n284 B.n283 163.367
R918 B.n288 B.n287 163.367
R919 B.n292 B.n291 163.367
R920 B.n296 B.n295 163.367
R921 B.n300 B.n299 163.367
R922 B.n304 B.n303 163.367
R923 B.n308 B.n307 163.367
R924 B.n312 B.n311 163.367
R925 B.n808 B.n123 163.367
R926 B.n543 B.t14 141.431
R927 B.n124 B.t16 141.431
R928 B.n420 B.t7 141.416
R929 B.n127 B.t10 141.416
R930 B.n636 B.n392 78.9494
R931 B.n810 B.n809 78.9494
R932 B.n442 B.n391 71.676
R933 B.n448 B.n447 71.676
R934 B.n451 B.n450 71.676
R935 B.n456 B.n455 71.676
R936 B.n459 B.n458 71.676
R937 B.n464 B.n463 71.676
R938 B.n467 B.n466 71.676
R939 B.n472 B.n471 71.676
R940 B.n475 B.n474 71.676
R941 B.n480 B.n479 71.676
R942 B.n483 B.n482 71.676
R943 B.n488 B.n487 71.676
R944 B.n491 B.n490 71.676
R945 B.n496 B.n495 71.676
R946 B.n499 B.n498 71.676
R947 B.n504 B.n503 71.676
R948 B.n507 B.n506 71.676
R949 B.n512 B.n511 71.676
R950 B.n515 B.n514 71.676
R951 B.n520 B.n519 71.676
R952 B.n523 B.n522 71.676
R953 B.n529 B.n528 71.676
R954 B.n532 B.n531 71.676
R955 B.n537 B.n536 71.676
R956 B.n540 B.n539 71.676
R957 B.n548 B.n547 71.676
R958 B.n551 B.n550 71.676
R959 B.n556 B.n555 71.676
R960 B.n559 B.n558 71.676
R961 B.n564 B.n563 71.676
R962 B.n567 B.n566 71.676
R963 B.n572 B.n571 71.676
R964 B.n575 B.n574 71.676
R965 B.n580 B.n579 71.676
R966 B.n583 B.n582 71.676
R967 B.n588 B.n587 71.676
R968 B.n591 B.n590 71.676
R969 B.n596 B.n595 71.676
R970 B.n599 B.n598 71.676
R971 B.n604 B.n603 71.676
R972 B.n607 B.n606 71.676
R973 B.n612 B.n611 71.676
R974 B.n615 B.n614 71.676
R975 B.n620 B.n619 71.676
R976 B.n623 B.n622 71.676
R977 B.n628 B.n627 71.676
R978 B.n631 B.n630 71.676
R979 B.n76 B.n74 71.676
R980 B.n131 B.n77 71.676
R981 B.n135 B.n78 71.676
R982 B.n139 B.n79 71.676
R983 B.n143 B.n80 71.676
R984 B.n147 B.n81 71.676
R985 B.n151 B.n82 71.676
R986 B.n155 B.n83 71.676
R987 B.n159 B.n84 71.676
R988 B.n163 B.n85 71.676
R989 B.n167 B.n86 71.676
R990 B.n171 B.n87 71.676
R991 B.n175 B.n88 71.676
R992 B.n179 B.n89 71.676
R993 B.n183 B.n90 71.676
R994 B.n187 B.n91 71.676
R995 B.n191 B.n92 71.676
R996 B.n195 B.n93 71.676
R997 B.n199 B.n94 71.676
R998 B.n203 B.n95 71.676
R999 B.n207 B.n96 71.676
R1000 B.n211 B.n97 71.676
R1001 B.n216 B.n98 71.676
R1002 B.n220 B.n99 71.676
R1003 B.n224 B.n100 71.676
R1004 B.n228 B.n101 71.676
R1005 B.n232 B.n102 71.676
R1006 B.n236 B.n103 71.676
R1007 B.n240 B.n104 71.676
R1008 B.n244 B.n105 71.676
R1009 B.n248 B.n106 71.676
R1010 B.n252 B.n107 71.676
R1011 B.n256 B.n108 71.676
R1012 B.n260 B.n109 71.676
R1013 B.n264 B.n110 71.676
R1014 B.n268 B.n111 71.676
R1015 B.n272 B.n112 71.676
R1016 B.n276 B.n113 71.676
R1017 B.n280 B.n114 71.676
R1018 B.n284 B.n115 71.676
R1019 B.n288 B.n116 71.676
R1020 B.n292 B.n117 71.676
R1021 B.n296 B.n118 71.676
R1022 B.n300 B.n119 71.676
R1023 B.n304 B.n120 71.676
R1024 B.n308 B.n121 71.676
R1025 B.n312 B.n122 71.676
R1026 B.n123 B.n122 71.676
R1027 B.n311 B.n121 71.676
R1028 B.n307 B.n120 71.676
R1029 B.n303 B.n119 71.676
R1030 B.n299 B.n118 71.676
R1031 B.n295 B.n117 71.676
R1032 B.n291 B.n116 71.676
R1033 B.n287 B.n115 71.676
R1034 B.n283 B.n114 71.676
R1035 B.n279 B.n113 71.676
R1036 B.n275 B.n112 71.676
R1037 B.n271 B.n111 71.676
R1038 B.n267 B.n110 71.676
R1039 B.n263 B.n109 71.676
R1040 B.n259 B.n108 71.676
R1041 B.n255 B.n107 71.676
R1042 B.n251 B.n106 71.676
R1043 B.n247 B.n105 71.676
R1044 B.n243 B.n104 71.676
R1045 B.n239 B.n103 71.676
R1046 B.n235 B.n102 71.676
R1047 B.n231 B.n101 71.676
R1048 B.n227 B.n100 71.676
R1049 B.n223 B.n99 71.676
R1050 B.n219 B.n98 71.676
R1051 B.n215 B.n97 71.676
R1052 B.n210 B.n96 71.676
R1053 B.n206 B.n95 71.676
R1054 B.n202 B.n94 71.676
R1055 B.n198 B.n93 71.676
R1056 B.n194 B.n92 71.676
R1057 B.n190 B.n91 71.676
R1058 B.n186 B.n90 71.676
R1059 B.n182 B.n89 71.676
R1060 B.n178 B.n88 71.676
R1061 B.n174 B.n87 71.676
R1062 B.n170 B.n86 71.676
R1063 B.n166 B.n85 71.676
R1064 B.n162 B.n84 71.676
R1065 B.n158 B.n83 71.676
R1066 B.n154 B.n82 71.676
R1067 B.n150 B.n81 71.676
R1068 B.n146 B.n80 71.676
R1069 B.n142 B.n79 71.676
R1070 B.n138 B.n78 71.676
R1071 B.n134 B.n77 71.676
R1072 B.n130 B.n76 71.676
R1073 B.n443 B.n442 71.676
R1074 B.n449 B.n448 71.676
R1075 B.n450 B.n439 71.676
R1076 B.n457 B.n456 71.676
R1077 B.n458 B.n437 71.676
R1078 B.n465 B.n464 71.676
R1079 B.n466 B.n435 71.676
R1080 B.n473 B.n472 71.676
R1081 B.n474 B.n433 71.676
R1082 B.n481 B.n480 71.676
R1083 B.n482 B.n431 71.676
R1084 B.n489 B.n488 71.676
R1085 B.n490 B.n429 71.676
R1086 B.n497 B.n496 71.676
R1087 B.n498 B.n427 71.676
R1088 B.n505 B.n504 71.676
R1089 B.n506 B.n425 71.676
R1090 B.n513 B.n512 71.676
R1091 B.n514 B.n423 71.676
R1092 B.n521 B.n520 71.676
R1093 B.n522 B.n419 71.676
R1094 B.n530 B.n529 71.676
R1095 B.n531 B.n417 71.676
R1096 B.n538 B.n537 71.676
R1097 B.n539 B.n415 71.676
R1098 B.n549 B.n548 71.676
R1099 B.n550 B.n413 71.676
R1100 B.n557 B.n556 71.676
R1101 B.n558 B.n411 71.676
R1102 B.n565 B.n564 71.676
R1103 B.n566 B.n409 71.676
R1104 B.n573 B.n572 71.676
R1105 B.n574 B.n407 71.676
R1106 B.n581 B.n580 71.676
R1107 B.n582 B.n405 71.676
R1108 B.n589 B.n588 71.676
R1109 B.n590 B.n403 71.676
R1110 B.n597 B.n596 71.676
R1111 B.n598 B.n401 71.676
R1112 B.n605 B.n604 71.676
R1113 B.n606 B.n399 71.676
R1114 B.n613 B.n612 71.676
R1115 B.n614 B.n397 71.676
R1116 B.n621 B.n620 71.676
R1117 B.n622 B.n395 71.676
R1118 B.n629 B.n628 71.676
R1119 B.n630 B.n393 71.676
R1120 B.n544 B.t13 71.2255
R1121 B.n125 B.t17 71.2255
R1122 B.n421 B.t6 71.2098
R1123 B.n128 B.t11 71.2098
R1124 B.n544 B.n543 70.2066
R1125 B.n421 B.n420 70.2066
R1126 B.n128 B.n127 70.2066
R1127 B.n125 B.n124 70.2066
R1128 B.n545 B.n544 59.5399
R1129 B.n526 B.n421 59.5399
R1130 B.n213 B.n128 59.5399
R1131 B.n126 B.n125 59.5399
R1132 B.n636 B.n388 42.2723
R1133 B.n642 B.n388 42.2723
R1134 B.n642 B.n384 42.2723
R1135 B.n648 B.n384 42.2723
R1136 B.n648 B.n380 42.2723
R1137 B.n654 B.n380 42.2723
R1138 B.n654 B.n376 42.2723
R1139 B.n660 B.n376 42.2723
R1140 B.n666 B.n372 42.2723
R1141 B.n666 B.n368 42.2723
R1142 B.n672 B.n368 42.2723
R1143 B.n672 B.n364 42.2723
R1144 B.n678 B.n364 42.2723
R1145 B.n678 B.n360 42.2723
R1146 B.n684 B.n360 42.2723
R1147 B.n684 B.n356 42.2723
R1148 B.n690 B.n356 42.2723
R1149 B.n690 B.n352 42.2723
R1150 B.n696 B.n352 42.2723
R1151 B.n696 B.n348 42.2723
R1152 B.n702 B.n348 42.2723
R1153 B.n708 B.n344 42.2723
R1154 B.n708 B.n340 42.2723
R1155 B.n714 B.n340 42.2723
R1156 B.n714 B.n336 42.2723
R1157 B.n720 B.n336 42.2723
R1158 B.n720 B.n332 42.2723
R1159 B.n726 B.n332 42.2723
R1160 B.n726 B.n328 42.2723
R1161 B.n733 B.n328 42.2723
R1162 B.n733 B.n732 42.2723
R1163 B.n739 B.n321 42.2723
R1164 B.n746 B.n321 42.2723
R1165 B.n746 B.n317 42.2723
R1166 B.n752 B.n317 42.2723
R1167 B.n752 B.n4 42.2723
R1168 B.n890 B.n4 42.2723
R1169 B.n890 B.n889 42.2723
R1170 B.n889 B.n888 42.2723
R1171 B.n888 B.n8 42.2723
R1172 B.n882 B.n8 42.2723
R1173 B.n882 B.n881 42.2723
R1174 B.n881 B.n880 42.2723
R1175 B.n874 B.n18 42.2723
R1176 B.n874 B.n873 42.2723
R1177 B.n873 B.n872 42.2723
R1178 B.n872 B.n22 42.2723
R1179 B.n866 B.n22 42.2723
R1180 B.n866 B.n865 42.2723
R1181 B.n865 B.n864 42.2723
R1182 B.n864 B.n29 42.2723
R1183 B.n858 B.n29 42.2723
R1184 B.n858 B.n857 42.2723
R1185 B.n856 B.n36 42.2723
R1186 B.n850 B.n36 42.2723
R1187 B.n850 B.n849 42.2723
R1188 B.n849 B.n848 42.2723
R1189 B.n848 B.n43 42.2723
R1190 B.n842 B.n43 42.2723
R1191 B.n842 B.n841 42.2723
R1192 B.n841 B.n840 42.2723
R1193 B.n840 B.n50 42.2723
R1194 B.n834 B.n50 42.2723
R1195 B.n834 B.n833 42.2723
R1196 B.n833 B.n832 42.2723
R1197 B.n832 B.n57 42.2723
R1198 B.n826 B.n825 42.2723
R1199 B.n825 B.n824 42.2723
R1200 B.n824 B.n64 42.2723
R1201 B.n818 B.n64 42.2723
R1202 B.n818 B.n817 42.2723
R1203 B.n817 B.n816 42.2723
R1204 B.n816 B.n71 42.2723
R1205 B.n810 B.n71 42.2723
R1206 B.n739 B.t2 39.1641
R1207 B.n880 B.t1 39.1641
R1208 B.n812 B.n73 34.4981
R1209 B.n807 B.n806 34.4981
R1210 B.n634 B.n633 34.4981
R1211 B.n638 B.n390 34.4981
R1212 B.n660 B.t5 24.2446
R1213 B.t0 B.n344 24.2446
R1214 B.n857 B.t3 24.2446
R1215 B.n826 B.t9 24.2446
R1216 B B.n892 18.0485
R1217 B.t5 B.n372 18.0282
R1218 B.n702 B.t0 18.0282
R1219 B.t3 B.n856 18.0282
R1220 B.t9 B.n57 18.0282
R1221 B.n129 B.n73 10.6151
R1222 B.n132 B.n129 10.6151
R1223 B.n133 B.n132 10.6151
R1224 B.n136 B.n133 10.6151
R1225 B.n137 B.n136 10.6151
R1226 B.n140 B.n137 10.6151
R1227 B.n141 B.n140 10.6151
R1228 B.n144 B.n141 10.6151
R1229 B.n145 B.n144 10.6151
R1230 B.n148 B.n145 10.6151
R1231 B.n149 B.n148 10.6151
R1232 B.n152 B.n149 10.6151
R1233 B.n153 B.n152 10.6151
R1234 B.n156 B.n153 10.6151
R1235 B.n157 B.n156 10.6151
R1236 B.n160 B.n157 10.6151
R1237 B.n161 B.n160 10.6151
R1238 B.n164 B.n161 10.6151
R1239 B.n165 B.n164 10.6151
R1240 B.n168 B.n165 10.6151
R1241 B.n169 B.n168 10.6151
R1242 B.n172 B.n169 10.6151
R1243 B.n173 B.n172 10.6151
R1244 B.n176 B.n173 10.6151
R1245 B.n177 B.n176 10.6151
R1246 B.n180 B.n177 10.6151
R1247 B.n181 B.n180 10.6151
R1248 B.n184 B.n181 10.6151
R1249 B.n185 B.n184 10.6151
R1250 B.n188 B.n185 10.6151
R1251 B.n189 B.n188 10.6151
R1252 B.n192 B.n189 10.6151
R1253 B.n193 B.n192 10.6151
R1254 B.n196 B.n193 10.6151
R1255 B.n197 B.n196 10.6151
R1256 B.n200 B.n197 10.6151
R1257 B.n201 B.n200 10.6151
R1258 B.n204 B.n201 10.6151
R1259 B.n205 B.n204 10.6151
R1260 B.n208 B.n205 10.6151
R1261 B.n209 B.n208 10.6151
R1262 B.n212 B.n209 10.6151
R1263 B.n217 B.n214 10.6151
R1264 B.n218 B.n217 10.6151
R1265 B.n221 B.n218 10.6151
R1266 B.n222 B.n221 10.6151
R1267 B.n225 B.n222 10.6151
R1268 B.n226 B.n225 10.6151
R1269 B.n229 B.n226 10.6151
R1270 B.n230 B.n229 10.6151
R1271 B.n234 B.n233 10.6151
R1272 B.n237 B.n234 10.6151
R1273 B.n238 B.n237 10.6151
R1274 B.n241 B.n238 10.6151
R1275 B.n242 B.n241 10.6151
R1276 B.n245 B.n242 10.6151
R1277 B.n246 B.n245 10.6151
R1278 B.n249 B.n246 10.6151
R1279 B.n250 B.n249 10.6151
R1280 B.n253 B.n250 10.6151
R1281 B.n254 B.n253 10.6151
R1282 B.n257 B.n254 10.6151
R1283 B.n258 B.n257 10.6151
R1284 B.n261 B.n258 10.6151
R1285 B.n262 B.n261 10.6151
R1286 B.n265 B.n262 10.6151
R1287 B.n266 B.n265 10.6151
R1288 B.n269 B.n266 10.6151
R1289 B.n270 B.n269 10.6151
R1290 B.n273 B.n270 10.6151
R1291 B.n274 B.n273 10.6151
R1292 B.n277 B.n274 10.6151
R1293 B.n278 B.n277 10.6151
R1294 B.n281 B.n278 10.6151
R1295 B.n282 B.n281 10.6151
R1296 B.n285 B.n282 10.6151
R1297 B.n286 B.n285 10.6151
R1298 B.n289 B.n286 10.6151
R1299 B.n290 B.n289 10.6151
R1300 B.n293 B.n290 10.6151
R1301 B.n294 B.n293 10.6151
R1302 B.n297 B.n294 10.6151
R1303 B.n298 B.n297 10.6151
R1304 B.n301 B.n298 10.6151
R1305 B.n302 B.n301 10.6151
R1306 B.n305 B.n302 10.6151
R1307 B.n306 B.n305 10.6151
R1308 B.n309 B.n306 10.6151
R1309 B.n310 B.n309 10.6151
R1310 B.n313 B.n310 10.6151
R1311 B.n314 B.n313 10.6151
R1312 B.n807 B.n314 10.6151
R1313 B.n634 B.n386 10.6151
R1314 B.n644 B.n386 10.6151
R1315 B.n645 B.n644 10.6151
R1316 B.n646 B.n645 10.6151
R1317 B.n646 B.n378 10.6151
R1318 B.n656 B.n378 10.6151
R1319 B.n657 B.n656 10.6151
R1320 B.n658 B.n657 10.6151
R1321 B.n658 B.n370 10.6151
R1322 B.n668 B.n370 10.6151
R1323 B.n669 B.n668 10.6151
R1324 B.n670 B.n669 10.6151
R1325 B.n670 B.n362 10.6151
R1326 B.n680 B.n362 10.6151
R1327 B.n681 B.n680 10.6151
R1328 B.n682 B.n681 10.6151
R1329 B.n682 B.n354 10.6151
R1330 B.n692 B.n354 10.6151
R1331 B.n693 B.n692 10.6151
R1332 B.n694 B.n693 10.6151
R1333 B.n694 B.n346 10.6151
R1334 B.n704 B.n346 10.6151
R1335 B.n705 B.n704 10.6151
R1336 B.n706 B.n705 10.6151
R1337 B.n706 B.n338 10.6151
R1338 B.n716 B.n338 10.6151
R1339 B.n717 B.n716 10.6151
R1340 B.n718 B.n717 10.6151
R1341 B.n718 B.n330 10.6151
R1342 B.n728 B.n330 10.6151
R1343 B.n729 B.n728 10.6151
R1344 B.n730 B.n729 10.6151
R1345 B.n730 B.n323 10.6151
R1346 B.n741 B.n323 10.6151
R1347 B.n742 B.n741 10.6151
R1348 B.n744 B.n742 10.6151
R1349 B.n744 B.n743 10.6151
R1350 B.n743 B.n315 10.6151
R1351 B.n755 B.n315 10.6151
R1352 B.n756 B.n755 10.6151
R1353 B.n757 B.n756 10.6151
R1354 B.n758 B.n757 10.6151
R1355 B.n760 B.n758 10.6151
R1356 B.n761 B.n760 10.6151
R1357 B.n762 B.n761 10.6151
R1358 B.n763 B.n762 10.6151
R1359 B.n765 B.n763 10.6151
R1360 B.n766 B.n765 10.6151
R1361 B.n767 B.n766 10.6151
R1362 B.n768 B.n767 10.6151
R1363 B.n770 B.n768 10.6151
R1364 B.n771 B.n770 10.6151
R1365 B.n772 B.n771 10.6151
R1366 B.n773 B.n772 10.6151
R1367 B.n775 B.n773 10.6151
R1368 B.n776 B.n775 10.6151
R1369 B.n777 B.n776 10.6151
R1370 B.n778 B.n777 10.6151
R1371 B.n780 B.n778 10.6151
R1372 B.n781 B.n780 10.6151
R1373 B.n782 B.n781 10.6151
R1374 B.n783 B.n782 10.6151
R1375 B.n785 B.n783 10.6151
R1376 B.n786 B.n785 10.6151
R1377 B.n787 B.n786 10.6151
R1378 B.n788 B.n787 10.6151
R1379 B.n790 B.n788 10.6151
R1380 B.n791 B.n790 10.6151
R1381 B.n792 B.n791 10.6151
R1382 B.n793 B.n792 10.6151
R1383 B.n795 B.n793 10.6151
R1384 B.n796 B.n795 10.6151
R1385 B.n797 B.n796 10.6151
R1386 B.n798 B.n797 10.6151
R1387 B.n800 B.n798 10.6151
R1388 B.n801 B.n800 10.6151
R1389 B.n802 B.n801 10.6151
R1390 B.n803 B.n802 10.6151
R1391 B.n805 B.n803 10.6151
R1392 B.n806 B.n805 10.6151
R1393 B.n444 B.n390 10.6151
R1394 B.n445 B.n444 10.6151
R1395 B.n446 B.n445 10.6151
R1396 B.n446 B.n440 10.6151
R1397 B.n452 B.n440 10.6151
R1398 B.n453 B.n452 10.6151
R1399 B.n454 B.n453 10.6151
R1400 B.n454 B.n438 10.6151
R1401 B.n460 B.n438 10.6151
R1402 B.n461 B.n460 10.6151
R1403 B.n462 B.n461 10.6151
R1404 B.n462 B.n436 10.6151
R1405 B.n468 B.n436 10.6151
R1406 B.n469 B.n468 10.6151
R1407 B.n470 B.n469 10.6151
R1408 B.n470 B.n434 10.6151
R1409 B.n476 B.n434 10.6151
R1410 B.n477 B.n476 10.6151
R1411 B.n478 B.n477 10.6151
R1412 B.n478 B.n432 10.6151
R1413 B.n484 B.n432 10.6151
R1414 B.n485 B.n484 10.6151
R1415 B.n486 B.n485 10.6151
R1416 B.n486 B.n430 10.6151
R1417 B.n492 B.n430 10.6151
R1418 B.n493 B.n492 10.6151
R1419 B.n494 B.n493 10.6151
R1420 B.n494 B.n428 10.6151
R1421 B.n500 B.n428 10.6151
R1422 B.n501 B.n500 10.6151
R1423 B.n502 B.n501 10.6151
R1424 B.n502 B.n426 10.6151
R1425 B.n508 B.n426 10.6151
R1426 B.n509 B.n508 10.6151
R1427 B.n510 B.n509 10.6151
R1428 B.n510 B.n424 10.6151
R1429 B.n516 B.n424 10.6151
R1430 B.n517 B.n516 10.6151
R1431 B.n518 B.n517 10.6151
R1432 B.n518 B.n422 10.6151
R1433 B.n524 B.n422 10.6151
R1434 B.n525 B.n524 10.6151
R1435 B.n527 B.n418 10.6151
R1436 B.n533 B.n418 10.6151
R1437 B.n534 B.n533 10.6151
R1438 B.n535 B.n534 10.6151
R1439 B.n535 B.n416 10.6151
R1440 B.n541 B.n416 10.6151
R1441 B.n542 B.n541 10.6151
R1442 B.n546 B.n542 10.6151
R1443 B.n552 B.n414 10.6151
R1444 B.n553 B.n552 10.6151
R1445 B.n554 B.n553 10.6151
R1446 B.n554 B.n412 10.6151
R1447 B.n560 B.n412 10.6151
R1448 B.n561 B.n560 10.6151
R1449 B.n562 B.n561 10.6151
R1450 B.n562 B.n410 10.6151
R1451 B.n568 B.n410 10.6151
R1452 B.n569 B.n568 10.6151
R1453 B.n570 B.n569 10.6151
R1454 B.n570 B.n408 10.6151
R1455 B.n576 B.n408 10.6151
R1456 B.n577 B.n576 10.6151
R1457 B.n578 B.n577 10.6151
R1458 B.n578 B.n406 10.6151
R1459 B.n584 B.n406 10.6151
R1460 B.n585 B.n584 10.6151
R1461 B.n586 B.n585 10.6151
R1462 B.n586 B.n404 10.6151
R1463 B.n592 B.n404 10.6151
R1464 B.n593 B.n592 10.6151
R1465 B.n594 B.n593 10.6151
R1466 B.n594 B.n402 10.6151
R1467 B.n600 B.n402 10.6151
R1468 B.n601 B.n600 10.6151
R1469 B.n602 B.n601 10.6151
R1470 B.n602 B.n400 10.6151
R1471 B.n608 B.n400 10.6151
R1472 B.n609 B.n608 10.6151
R1473 B.n610 B.n609 10.6151
R1474 B.n610 B.n398 10.6151
R1475 B.n616 B.n398 10.6151
R1476 B.n617 B.n616 10.6151
R1477 B.n618 B.n617 10.6151
R1478 B.n618 B.n396 10.6151
R1479 B.n624 B.n396 10.6151
R1480 B.n625 B.n624 10.6151
R1481 B.n626 B.n625 10.6151
R1482 B.n626 B.n394 10.6151
R1483 B.n632 B.n394 10.6151
R1484 B.n633 B.n632 10.6151
R1485 B.n639 B.n638 10.6151
R1486 B.n640 B.n639 10.6151
R1487 B.n640 B.n382 10.6151
R1488 B.n650 B.n382 10.6151
R1489 B.n651 B.n650 10.6151
R1490 B.n652 B.n651 10.6151
R1491 B.n652 B.n374 10.6151
R1492 B.n662 B.n374 10.6151
R1493 B.n663 B.n662 10.6151
R1494 B.n664 B.n663 10.6151
R1495 B.n664 B.n366 10.6151
R1496 B.n674 B.n366 10.6151
R1497 B.n675 B.n674 10.6151
R1498 B.n676 B.n675 10.6151
R1499 B.n676 B.n358 10.6151
R1500 B.n686 B.n358 10.6151
R1501 B.n687 B.n686 10.6151
R1502 B.n688 B.n687 10.6151
R1503 B.n688 B.n350 10.6151
R1504 B.n698 B.n350 10.6151
R1505 B.n699 B.n698 10.6151
R1506 B.n700 B.n699 10.6151
R1507 B.n700 B.n342 10.6151
R1508 B.n710 B.n342 10.6151
R1509 B.n711 B.n710 10.6151
R1510 B.n712 B.n711 10.6151
R1511 B.n712 B.n334 10.6151
R1512 B.n722 B.n334 10.6151
R1513 B.n723 B.n722 10.6151
R1514 B.n724 B.n723 10.6151
R1515 B.n724 B.n326 10.6151
R1516 B.n735 B.n326 10.6151
R1517 B.n736 B.n735 10.6151
R1518 B.n737 B.n736 10.6151
R1519 B.n737 B.n319 10.6151
R1520 B.n748 B.n319 10.6151
R1521 B.n749 B.n748 10.6151
R1522 B.n750 B.n749 10.6151
R1523 B.n750 B.n0 10.6151
R1524 B.n886 B.n1 10.6151
R1525 B.n886 B.n885 10.6151
R1526 B.n885 B.n884 10.6151
R1527 B.n884 B.n10 10.6151
R1528 B.n878 B.n10 10.6151
R1529 B.n878 B.n877 10.6151
R1530 B.n877 B.n876 10.6151
R1531 B.n876 B.n16 10.6151
R1532 B.n870 B.n16 10.6151
R1533 B.n870 B.n869 10.6151
R1534 B.n869 B.n868 10.6151
R1535 B.n868 B.n24 10.6151
R1536 B.n862 B.n24 10.6151
R1537 B.n862 B.n861 10.6151
R1538 B.n861 B.n860 10.6151
R1539 B.n860 B.n31 10.6151
R1540 B.n854 B.n31 10.6151
R1541 B.n854 B.n853 10.6151
R1542 B.n853 B.n852 10.6151
R1543 B.n852 B.n38 10.6151
R1544 B.n846 B.n38 10.6151
R1545 B.n846 B.n845 10.6151
R1546 B.n845 B.n844 10.6151
R1547 B.n844 B.n45 10.6151
R1548 B.n838 B.n45 10.6151
R1549 B.n838 B.n837 10.6151
R1550 B.n837 B.n836 10.6151
R1551 B.n836 B.n52 10.6151
R1552 B.n830 B.n52 10.6151
R1553 B.n830 B.n829 10.6151
R1554 B.n829 B.n828 10.6151
R1555 B.n828 B.n59 10.6151
R1556 B.n822 B.n59 10.6151
R1557 B.n822 B.n821 10.6151
R1558 B.n821 B.n820 10.6151
R1559 B.n820 B.n66 10.6151
R1560 B.n814 B.n66 10.6151
R1561 B.n814 B.n813 10.6151
R1562 B.n813 B.n812 10.6151
R1563 B.n214 B.n213 6.5566
R1564 B.n230 B.n126 6.5566
R1565 B.n527 B.n526 6.5566
R1566 B.n546 B.n545 6.5566
R1567 B.n213 B.n212 4.05904
R1568 B.n233 B.n126 4.05904
R1569 B.n526 B.n525 4.05904
R1570 B.n545 B.n414 4.05904
R1571 B.n732 B.t2 3.10872
R1572 B.n18 B.t1 3.10872
R1573 B.n892 B.n0 2.81026
R1574 B.n892 B.n1 2.81026
R1575 VN.n1 VN.t0 125.968
R1576 VN.n0 VN.t3 125.968
R1577 VN.n0 VN.t1 124.85
R1578 VN.n1 VN.t2 124.85
R1579 VN VN.n1 51.4645
R1580 VN VN.n0 2.49097
R1581 VDD2.n2 VDD2.n0 104.407
R1582 VDD2.n2 VDD2.n1 60.6237
R1583 VDD2.n1 VDD2.t1 1.5947
R1584 VDD2.n1 VDD2.t3 1.5947
R1585 VDD2.n0 VDD2.t0 1.5947
R1586 VDD2.n0 VDD2.t2 1.5947
R1587 VDD2 VDD2.n2 0.0586897
C0 VDD2 VTAIL 5.72287f
C1 VDD2 VN 5.10043f
C2 VN VTAIL 5.0899f
C3 VDD1 VP 5.3881f
C4 VDD2 VDD1 1.18708f
C5 VDD1 VTAIL 5.66404f
C6 VN VDD1 0.149804f
C7 VDD2 VP 0.438392f
C8 VP VTAIL 5.10401f
C9 VN VP 6.76207f
C10 VDD2 B 4.195462f
C11 VDD1 B 8.65426f
C12 VTAIL B 10.712701f
C13 VN B 12.06f
C14 VP B 10.438472f
C15 VDD2.t0 B 0.264957f
C16 VDD2.t2 B 0.264957f
C17 VDD2.n0 B 3.10276f
C18 VDD2.t1 B 0.264957f
C19 VDD2.t3 B 0.264957f
C20 VDD2.n1 B 2.36409f
C21 VDD2.n2 B 3.99605f
C22 VN.t1 B 2.70559f
C23 VN.t3 B 2.71425f
C24 VN.n0 B 1.64248f
C25 VN.t2 B 2.70559f
C26 VN.t0 B 2.71425f
C27 VN.n1 B 3.00295f
C28 VDD1.t0 B 0.269826f
C29 VDD1.t3 B 0.269826f
C30 VDD1.n0 B 2.40803f
C31 VDD1.t2 B 0.269826f
C32 VDD1.t1 B 0.269826f
C33 VDD1.n1 B 3.18792f
C34 VTAIL.t1 B 1.80344f
C35 VTAIL.n0 B 0.341344f
C36 VTAIL.t4 B 1.80344f
C37 VTAIL.n1 B 0.422404f
C38 VTAIL.t7 B 1.80344f
C39 VTAIL.n2 B 1.37071f
C40 VTAIL.t0 B 1.80345f
C41 VTAIL.n3 B 1.3707f
C42 VTAIL.t2 B 1.80345f
C43 VTAIL.n4 B 0.422392f
C44 VTAIL.t6 B 1.80345f
C45 VTAIL.n5 B 0.422392f
C46 VTAIL.t5 B 1.80344f
C47 VTAIL.n6 B 1.37071f
C48 VTAIL.t3 B 1.80344f
C49 VTAIL.n7 B 1.28337f
C50 VP.t2 B 2.4793f
C51 VP.n0 B 0.957024f
C52 VP.n1 B 0.022248f
C53 VP.n2 B 0.017969f
C54 VP.n3 B 0.022248f
C55 VP.t1 B 2.4793f
C56 VP.n4 B 0.957024f
C57 VP.t3 B 2.76714f
C58 VP.t0 B 2.75831f
C59 VP.n5 B 3.0525f
C60 VP.n6 B 1.31175f
C61 VP.n7 B 0.035902f
C62 VP.n8 B 0.033517f
C63 VP.n9 B 0.041256f
C64 VP.n10 B 0.043984f
C65 VP.n11 B 0.022248f
C66 VP.n12 B 0.022248f
C67 VP.n13 B 0.022248f
C68 VP.n14 B 0.043984f
C69 VP.n15 B 0.041256f
C70 VP.n16 B 0.033517f
C71 VP.n17 B 0.035902f
C72 VP.n18 B 0.053252f
.ends

