* NGSPICE file created from diff_pair_sample_0159.ext - technology: sky130A

.subckt diff_pair_sample_0159 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X1 VDD1.t6 VP.t1 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=5.8227 ps=30.64 w=14.93 l=3.12
X2 VDD2.t7 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X3 VDD1.t5 VP.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X4 VDD1.t4 VP.t3 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=5.8227 ps=30.64 w=14.93 l=3.12
X5 VTAIL.t15 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=2.46345 ps=15.26 w=14.93 l=3.12
X6 VTAIL.t5 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X7 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=0 ps=0 w=14.93 l=3.12
X8 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=0 ps=0 w=14.93 l=3.12
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=0 ps=0 w=14.93 l=3.12
X10 VTAIL.t7 VP.t4 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=2.46345 ps=15.26 w=14.93 l=3.12
X11 VTAIL.t6 VP.t5 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X12 VDD2.t4 VN.t3 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=5.8227 ps=30.64 w=14.93 l=3.12
X13 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X14 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=5.8227 ps=30.64 w=14.93 l=3.12
X15 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X16 VTAIL.t12 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.46345 pd=15.26 as=2.46345 ps=15.26 w=14.93 l=3.12
X17 VTAIL.t8 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=2.46345 ps=15.26 w=14.93 l=3.12
X18 VTAIL.t2 VN.t7 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=2.46345 ps=15.26 w=14.93 l=3.12
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.8227 pd=30.64 as=0 ps=0 w=14.93 l=3.12
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n19 VP.t7 148.738
R34 VP.n43 VP.t4 115.326
R35 VP.n55 VP.t2 115.326
R36 VP.n4 VP.t5 115.326
R37 VP.n0 VP.t1 115.326
R38 VP.n11 VP.t3 115.326
R39 VP.n15 VP.t6 115.326
R40 VP.n20 VP.t0 115.326
R41 VP.n43 VP.n42 69.2705
R42 VP.n76 VP.n0 69.2705
R43 VP.n41 VP.n11 69.2705
R44 VP.n49 VP.n48 56.5193
R45 VP.n61 VP.n6 56.5193
R46 VP.n72 VP.n2 56.5193
R47 VP.n37 VP.n13 56.5193
R48 VP.n26 VP.n17 56.5193
R49 VP.n42 VP.n41 55.7114
R50 VP.n20 VP.n19 50.6608
R51 VP.n44 VP.n10 24.4675
R52 VP.n48 VP.n10 24.4675
R53 VP.n50 VP.n49 24.4675
R54 VP.n50 VP.n8 24.4675
R55 VP.n54 VP.n8 24.4675
R56 VP.n57 VP.n56 24.4675
R57 VP.n57 VP.n6 24.4675
R58 VP.n62 VP.n61 24.4675
R59 VP.n63 VP.n62 24.4675
R60 VP.n67 VP.n66 24.4675
R61 VP.n68 VP.n67 24.4675
R62 VP.n68 VP.n2 24.4675
R63 VP.n73 VP.n72 24.4675
R64 VP.n74 VP.n73 24.4675
R65 VP.n38 VP.n37 24.4675
R66 VP.n39 VP.n38 24.4675
R67 VP.n27 VP.n26 24.4675
R68 VP.n28 VP.n27 24.4675
R69 VP.n32 VP.n31 24.4675
R70 VP.n33 VP.n32 24.4675
R71 VP.n33 VP.n13 24.4675
R72 VP.n22 VP.n21 24.4675
R73 VP.n22 VP.n17 24.4675
R74 VP.n56 VP.n55 23.2442
R75 VP.n63 VP.n4 23.2442
R76 VP.n28 VP.n15 23.2442
R77 VP.n21 VP.n20 23.2442
R78 VP.n44 VP.n43 20.7975
R79 VP.n74 VP.n0 20.7975
R80 VP.n39 VP.n11 20.7975
R81 VP.n19 VP.n18 3.87631
R82 VP.n55 VP.n54 1.22385
R83 VP.n66 VP.n4 1.22385
R84 VP.n31 VP.n15 1.22385
R85 VP.n41 VP.n40 0.354971
R86 VP.n45 VP.n42 0.354971
R87 VP.n76 VP.n75 0.354971
R88 VP VP.n76 0.26696
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VTAIL.n658 VTAIL.n582 289.615
R121 VTAIL.n78 VTAIL.n2 289.615
R122 VTAIL.n160 VTAIL.n84 289.615
R123 VTAIL.n244 VTAIL.n168 289.615
R124 VTAIL.n576 VTAIL.n500 289.615
R125 VTAIL.n492 VTAIL.n416 289.615
R126 VTAIL.n410 VTAIL.n334 289.615
R127 VTAIL.n326 VTAIL.n250 289.615
R128 VTAIL.n609 VTAIL.n608 185
R129 VTAIL.n606 VTAIL.n605 185
R130 VTAIL.n615 VTAIL.n614 185
R131 VTAIL.n617 VTAIL.n616 185
R132 VTAIL.n602 VTAIL.n601 185
R133 VTAIL.n623 VTAIL.n622 185
R134 VTAIL.n626 VTAIL.n625 185
R135 VTAIL.n624 VTAIL.n598 185
R136 VTAIL.n631 VTAIL.n597 185
R137 VTAIL.n633 VTAIL.n632 185
R138 VTAIL.n635 VTAIL.n634 185
R139 VTAIL.n594 VTAIL.n593 185
R140 VTAIL.n641 VTAIL.n640 185
R141 VTAIL.n643 VTAIL.n642 185
R142 VTAIL.n590 VTAIL.n589 185
R143 VTAIL.n649 VTAIL.n648 185
R144 VTAIL.n651 VTAIL.n650 185
R145 VTAIL.n586 VTAIL.n585 185
R146 VTAIL.n657 VTAIL.n656 185
R147 VTAIL.n659 VTAIL.n658 185
R148 VTAIL.n29 VTAIL.n28 185
R149 VTAIL.n26 VTAIL.n25 185
R150 VTAIL.n35 VTAIL.n34 185
R151 VTAIL.n37 VTAIL.n36 185
R152 VTAIL.n22 VTAIL.n21 185
R153 VTAIL.n43 VTAIL.n42 185
R154 VTAIL.n46 VTAIL.n45 185
R155 VTAIL.n44 VTAIL.n18 185
R156 VTAIL.n51 VTAIL.n17 185
R157 VTAIL.n53 VTAIL.n52 185
R158 VTAIL.n55 VTAIL.n54 185
R159 VTAIL.n14 VTAIL.n13 185
R160 VTAIL.n61 VTAIL.n60 185
R161 VTAIL.n63 VTAIL.n62 185
R162 VTAIL.n10 VTAIL.n9 185
R163 VTAIL.n69 VTAIL.n68 185
R164 VTAIL.n71 VTAIL.n70 185
R165 VTAIL.n6 VTAIL.n5 185
R166 VTAIL.n77 VTAIL.n76 185
R167 VTAIL.n79 VTAIL.n78 185
R168 VTAIL.n111 VTAIL.n110 185
R169 VTAIL.n108 VTAIL.n107 185
R170 VTAIL.n117 VTAIL.n116 185
R171 VTAIL.n119 VTAIL.n118 185
R172 VTAIL.n104 VTAIL.n103 185
R173 VTAIL.n125 VTAIL.n124 185
R174 VTAIL.n128 VTAIL.n127 185
R175 VTAIL.n126 VTAIL.n100 185
R176 VTAIL.n133 VTAIL.n99 185
R177 VTAIL.n135 VTAIL.n134 185
R178 VTAIL.n137 VTAIL.n136 185
R179 VTAIL.n96 VTAIL.n95 185
R180 VTAIL.n143 VTAIL.n142 185
R181 VTAIL.n145 VTAIL.n144 185
R182 VTAIL.n92 VTAIL.n91 185
R183 VTAIL.n151 VTAIL.n150 185
R184 VTAIL.n153 VTAIL.n152 185
R185 VTAIL.n88 VTAIL.n87 185
R186 VTAIL.n159 VTAIL.n158 185
R187 VTAIL.n161 VTAIL.n160 185
R188 VTAIL.n195 VTAIL.n194 185
R189 VTAIL.n192 VTAIL.n191 185
R190 VTAIL.n201 VTAIL.n200 185
R191 VTAIL.n203 VTAIL.n202 185
R192 VTAIL.n188 VTAIL.n187 185
R193 VTAIL.n209 VTAIL.n208 185
R194 VTAIL.n212 VTAIL.n211 185
R195 VTAIL.n210 VTAIL.n184 185
R196 VTAIL.n217 VTAIL.n183 185
R197 VTAIL.n219 VTAIL.n218 185
R198 VTAIL.n221 VTAIL.n220 185
R199 VTAIL.n180 VTAIL.n179 185
R200 VTAIL.n227 VTAIL.n226 185
R201 VTAIL.n229 VTAIL.n228 185
R202 VTAIL.n176 VTAIL.n175 185
R203 VTAIL.n235 VTAIL.n234 185
R204 VTAIL.n237 VTAIL.n236 185
R205 VTAIL.n172 VTAIL.n171 185
R206 VTAIL.n243 VTAIL.n242 185
R207 VTAIL.n245 VTAIL.n244 185
R208 VTAIL.n577 VTAIL.n576 185
R209 VTAIL.n575 VTAIL.n574 185
R210 VTAIL.n504 VTAIL.n503 185
R211 VTAIL.n569 VTAIL.n568 185
R212 VTAIL.n567 VTAIL.n566 185
R213 VTAIL.n508 VTAIL.n507 185
R214 VTAIL.n561 VTAIL.n560 185
R215 VTAIL.n559 VTAIL.n558 185
R216 VTAIL.n512 VTAIL.n511 185
R217 VTAIL.n553 VTAIL.n552 185
R218 VTAIL.n551 VTAIL.n550 185
R219 VTAIL.n549 VTAIL.n515 185
R220 VTAIL.n519 VTAIL.n516 185
R221 VTAIL.n544 VTAIL.n543 185
R222 VTAIL.n542 VTAIL.n541 185
R223 VTAIL.n521 VTAIL.n520 185
R224 VTAIL.n536 VTAIL.n535 185
R225 VTAIL.n534 VTAIL.n533 185
R226 VTAIL.n525 VTAIL.n524 185
R227 VTAIL.n528 VTAIL.n527 185
R228 VTAIL.n493 VTAIL.n492 185
R229 VTAIL.n491 VTAIL.n490 185
R230 VTAIL.n420 VTAIL.n419 185
R231 VTAIL.n485 VTAIL.n484 185
R232 VTAIL.n483 VTAIL.n482 185
R233 VTAIL.n424 VTAIL.n423 185
R234 VTAIL.n477 VTAIL.n476 185
R235 VTAIL.n475 VTAIL.n474 185
R236 VTAIL.n428 VTAIL.n427 185
R237 VTAIL.n469 VTAIL.n468 185
R238 VTAIL.n467 VTAIL.n466 185
R239 VTAIL.n465 VTAIL.n431 185
R240 VTAIL.n435 VTAIL.n432 185
R241 VTAIL.n460 VTAIL.n459 185
R242 VTAIL.n458 VTAIL.n457 185
R243 VTAIL.n437 VTAIL.n436 185
R244 VTAIL.n452 VTAIL.n451 185
R245 VTAIL.n450 VTAIL.n449 185
R246 VTAIL.n441 VTAIL.n440 185
R247 VTAIL.n444 VTAIL.n443 185
R248 VTAIL.n411 VTAIL.n410 185
R249 VTAIL.n409 VTAIL.n408 185
R250 VTAIL.n338 VTAIL.n337 185
R251 VTAIL.n403 VTAIL.n402 185
R252 VTAIL.n401 VTAIL.n400 185
R253 VTAIL.n342 VTAIL.n341 185
R254 VTAIL.n395 VTAIL.n394 185
R255 VTAIL.n393 VTAIL.n392 185
R256 VTAIL.n346 VTAIL.n345 185
R257 VTAIL.n387 VTAIL.n386 185
R258 VTAIL.n385 VTAIL.n384 185
R259 VTAIL.n383 VTAIL.n349 185
R260 VTAIL.n353 VTAIL.n350 185
R261 VTAIL.n378 VTAIL.n377 185
R262 VTAIL.n376 VTAIL.n375 185
R263 VTAIL.n355 VTAIL.n354 185
R264 VTAIL.n370 VTAIL.n369 185
R265 VTAIL.n368 VTAIL.n367 185
R266 VTAIL.n359 VTAIL.n358 185
R267 VTAIL.n362 VTAIL.n361 185
R268 VTAIL.n327 VTAIL.n326 185
R269 VTAIL.n325 VTAIL.n324 185
R270 VTAIL.n254 VTAIL.n253 185
R271 VTAIL.n319 VTAIL.n318 185
R272 VTAIL.n317 VTAIL.n316 185
R273 VTAIL.n258 VTAIL.n257 185
R274 VTAIL.n311 VTAIL.n310 185
R275 VTAIL.n309 VTAIL.n308 185
R276 VTAIL.n262 VTAIL.n261 185
R277 VTAIL.n303 VTAIL.n302 185
R278 VTAIL.n301 VTAIL.n300 185
R279 VTAIL.n299 VTAIL.n265 185
R280 VTAIL.n269 VTAIL.n266 185
R281 VTAIL.n294 VTAIL.n293 185
R282 VTAIL.n292 VTAIL.n291 185
R283 VTAIL.n271 VTAIL.n270 185
R284 VTAIL.n286 VTAIL.n285 185
R285 VTAIL.n284 VTAIL.n283 185
R286 VTAIL.n275 VTAIL.n274 185
R287 VTAIL.n278 VTAIL.n277 185
R288 VTAIL.t0 VTAIL.n607 149.524
R289 VTAIL.t15 VTAIL.n27 149.524
R290 VTAIL.t11 VTAIL.n109 149.524
R291 VTAIL.t7 VTAIL.n193 149.524
R292 VTAIL.t10 VTAIL.n526 149.524
R293 VTAIL.t8 VTAIL.n442 149.524
R294 VTAIL.t14 VTAIL.n360 149.524
R295 VTAIL.t2 VTAIL.n276 149.524
R296 VTAIL.n608 VTAIL.n605 104.615
R297 VTAIL.n615 VTAIL.n605 104.615
R298 VTAIL.n616 VTAIL.n615 104.615
R299 VTAIL.n616 VTAIL.n601 104.615
R300 VTAIL.n623 VTAIL.n601 104.615
R301 VTAIL.n625 VTAIL.n623 104.615
R302 VTAIL.n625 VTAIL.n624 104.615
R303 VTAIL.n624 VTAIL.n597 104.615
R304 VTAIL.n633 VTAIL.n597 104.615
R305 VTAIL.n634 VTAIL.n633 104.615
R306 VTAIL.n634 VTAIL.n593 104.615
R307 VTAIL.n641 VTAIL.n593 104.615
R308 VTAIL.n642 VTAIL.n641 104.615
R309 VTAIL.n642 VTAIL.n589 104.615
R310 VTAIL.n649 VTAIL.n589 104.615
R311 VTAIL.n650 VTAIL.n649 104.615
R312 VTAIL.n650 VTAIL.n585 104.615
R313 VTAIL.n657 VTAIL.n585 104.615
R314 VTAIL.n658 VTAIL.n657 104.615
R315 VTAIL.n28 VTAIL.n25 104.615
R316 VTAIL.n35 VTAIL.n25 104.615
R317 VTAIL.n36 VTAIL.n35 104.615
R318 VTAIL.n36 VTAIL.n21 104.615
R319 VTAIL.n43 VTAIL.n21 104.615
R320 VTAIL.n45 VTAIL.n43 104.615
R321 VTAIL.n45 VTAIL.n44 104.615
R322 VTAIL.n44 VTAIL.n17 104.615
R323 VTAIL.n53 VTAIL.n17 104.615
R324 VTAIL.n54 VTAIL.n53 104.615
R325 VTAIL.n54 VTAIL.n13 104.615
R326 VTAIL.n61 VTAIL.n13 104.615
R327 VTAIL.n62 VTAIL.n61 104.615
R328 VTAIL.n62 VTAIL.n9 104.615
R329 VTAIL.n69 VTAIL.n9 104.615
R330 VTAIL.n70 VTAIL.n69 104.615
R331 VTAIL.n70 VTAIL.n5 104.615
R332 VTAIL.n77 VTAIL.n5 104.615
R333 VTAIL.n78 VTAIL.n77 104.615
R334 VTAIL.n110 VTAIL.n107 104.615
R335 VTAIL.n117 VTAIL.n107 104.615
R336 VTAIL.n118 VTAIL.n117 104.615
R337 VTAIL.n118 VTAIL.n103 104.615
R338 VTAIL.n125 VTAIL.n103 104.615
R339 VTAIL.n127 VTAIL.n125 104.615
R340 VTAIL.n127 VTAIL.n126 104.615
R341 VTAIL.n126 VTAIL.n99 104.615
R342 VTAIL.n135 VTAIL.n99 104.615
R343 VTAIL.n136 VTAIL.n135 104.615
R344 VTAIL.n136 VTAIL.n95 104.615
R345 VTAIL.n143 VTAIL.n95 104.615
R346 VTAIL.n144 VTAIL.n143 104.615
R347 VTAIL.n144 VTAIL.n91 104.615
R348 VTAIL.n151 VTAIL.n91 104.615
R349 VTAIL.n152 VTAIL.n151 104.615
R350 VTAIL.n152 VTAIL.n87 104.615
R351 VTAIL.n159 VTAIL.n87 104.615
R352 VTAIL.n160 VTAIL.n159 104.615
R353 VTAIL.n194 VTAIL.n191 104.615
R354 VTAIL.n201 VTAIL.n191 104.615
R355 VTAIL.n202 VTAIL.n201 104.615
R356 VTAIL.n202 VTAIL.n187 104.615
R357 VTAIL.n209 VTAIL.n187 104.615
R358 VTAIL.n211 VTAIL.n209 104.615
R359 VTAIL.n211 VTAIL.n210 104.615
R360 VTAIL.n210 VTAIL.n183 104.615
R361 VTAIL.n219 VTAIL.n183 104.615
R362 VTAIL.n220 VTAIL.n219 104.615
R363 VTAIL.n220 VTAIL.n179 104.615
R364 VTAIL.n227 VTAIL.n179 104.615
R365 VTAIL.n228 VTAIL.n227 104.615
R366 VTAIL.n228 VTAIL.n175 104.615
R367 VTAIL.n235 VTAIL.n175 104.615
R368 VTAIL.n236 VTAIL.n235 104.615
R369 VTAIL.n236 VTAIL.n171 104.615
R370 VTAIL.n243 VTAIL.n171 104.615
R371 VTAIL.n244 VTAIL.n243 104.615
R372 VTAIL.n576 VTAIL.n575 104.615
R373 VTAIL.n575 VTAIL.n503 104.615
R374 VTAIL.n568 VTAIL.n503 104.615
R375 VTAIL.n568 VTAIL.n567 104.615
R376 VTAIL.n567 VTAIL.n507 104.615
R377 VTAIL.n560 VTAIL.n507 104.615
R378 VTAIL.n560 VTAIL.n559 104.615
R379 VTAIL.n559 VTAIL.n511 104.615
R380 VTAIL.n552 VTAIL.n511 104.615
R381 VTAIL.n552 VTAIL.n551 104.615
R382 VTAIL.n551 VTAIL.n515 104.615
R383 VTAIL.n519 VTAIL.n515 104.615
R384 VTAIL.n543 VTAIL.n519 104.615
R385 VTAIL.n543 VTAIL.n542 104.615
R386 VTAIL.n542 VTAIL.n520 104.615
R387 VTAIL.n535 VTAIL.n520 104.615
R388 VTAIL.n535 VTAIL.n534 104.615
R389 VTAIL.n534 VTAIL.n524 104.615
R390 VTAIL.n527 VTAIL.n524 104.615
R391 VTAIL.n492 VTAIL.n491 104.615
R392 VTAIL.n491 VTAIL.n419 104.615
R393 VTAIL.n484 VTAIL.n419 104.615
R394 VTAIL.n484 VTAIL.n483 104.615
R395 VTAIL.n483 VTAIL.n423 104.615
R396 VTAIL.n476 VTAIL.n423 104.615
R397 VTAIL.n476 VTAIL.n475 104.615
R398 VTAIL.n475 VTAIL.n427 104.615
R399 VTAIL.n468 VTAIL.n427 104.615
R400 VTAIL.n468 VTAIL.n467 104.615
R401 VTAIL.n467 VTAIL.n431 104.615
R402 VTAIL.n435 VTAIL.n431 104.615
R403 VTAIL.n459 VTAIL.n435 104.615
R404 VTAIL.n459 VTAIL.n458 104.615
R405 VTAIL.n458 VTAIL.n436 104.615
R406 VTAIL.n451 VTAIL.n436 104.615
R407 VTAIL.n451 VTAIL.n450 104.615
R408 VTAIL.n450 VTAIL.n440 104.615
R409 VTAIL.n443 VTAIL.n440 104.615
R410 VTAIL.n410 VTAIL.n409 104.615
R411 VTAIL.n409 VTAIL.n337 104.615
R412 VTAIL.n402 VTAIL.n337 104.615
R413 VTAIL.n402 VTAIL.n401 104.615
R414 VTAIL.n401 VTAIL.n341 104.615
R415 VTAIL.n394 VTAIL.n341 104.615
R416 VTAIL.n394 VTAIL.n393 104.615
R417 VTAIL.n393 VTAIL.n345 104.615
R418 VTAIL.n386 VTAIL.n345 104.615
R419 VTAIL.n386 VTAIL.n385 104.615
R420 VTAIL.n385 VTAIL.n349 104.615
R421 VTAIL.n353 VTAIL.n349 104.615
R422 VTAIL.n377 VTAIL.n353 104.615
R423 VTAIL.n377 VTAIL.n376 104.615
R424 VTAIL.n376 VTAIL.n354 104.615
R425 VTAIL.n369 VTAIL.n354 104.615
R426 VTAIL.n369 VTAIL.n368 104.615
R427 VTAIL.n368 VTAIL.n358 104.615
R428 VTAIL.n361 VTAIL.n358 104.615
R429 VTAIL.n326 VTAIL.n325 104.615
R430 VTAIL.n325 VTAIL.n253 104.615
R431 VTAIL.n318 VTAIL.n253 104.615
R432 VTAIL.n318 VTAIL.n317 104.615
R433 VTAIL.n317 VTAIL.n257 104.615
R434 VTAIL.n310 VTAIL.n257 104.615
R435 VTAIL.n310 VTAIL.n309 104.615
R436 VTAIL.n309 VTAIL.n261 104.615
R437 VTAIL.n302 VTAIL.n261 104.615
R438 VTAIL.n302 VTAIL.n301 104.615
R439 VTAIL.n301 VTAIL.n265 104.615
R440 VTAIL.n269 VTAIL.n265 104.615
R441 VTAIL.n293 VTAIL.n269 104.615
R442 VTAIL.n293 VTAIL.n292 104.615
R443 VTAIL.n292 VTAIL.n270 104.615
R444 VTAIL.n285 VTAIL.n270 104.615
R445 VTAIL.n285 VTAIL.n284 104.615
R446 VTAIL.n284 VTAIL.n274 104.615
R447 VTAIL.n277 VTAIL.n274 104.615
R448 VTAIL.n608 VTAIL.t0 52.3082
R449 VTAIL.n28 VTAIL.t15 52.3082
R450 VTAIL.n110 VTAIL.t11 52.3082
R451 VTAIL.n194 VTAIL.t7 52.3082
R452 VTAIL.n527 VTAIL.t10 52.3082
R453 VTAIL.n443 VTAIL.t8 52.3082
R454 VTAIL.n361 VTAIL.t14 52.3082
R455 VTAIL.n277 VTAIL.t2 52.3082
R456 VTAIL.n499 VTAIL.n498 43.2853
R457 VTAIL.n333 VTAIL.n332 43.2853
R458 VTAIL.n1 VTAIL.n0 43.2851
R459 VTAIL.n167 VTAIL.n166 43.2851
R460 VTAIL.n663 VTAIL.n662 30.8278
R461 VTAIL.n83 VTAIL.n82 30.8278
R462 VTAIL.n165 VTAIL.n164 30.8278
R463 VTAIL.n249 VTAIL.n248 30.8278
R464 VTAIL.n581 VTAIL.n580 30.8278
R465 VTAIL.n497 VTAIL.n496 30.8278
R466 VTAIL.n415 VTAIL.n414 30.8278
R467 VTAIL.n331 VTAIL.n330 30.8278
R468 VTAIL.n663 VTAIL.n581 28.2117
R469 VTAIL.n331 VTAIL.n249 28.2117
R470 VTAIL.n632 VTAIL.n631 13.1884
R471 VTAIL.n52 VTAIL.n51 13.1884
R472 VTAIL.n134 VTAIL.n133 13.1884
R473 VTAIL.n218 VTAIL.n217 13.1884
R474 VTAIL.n550 VTAIL.n549 13.1884
R475 VTAIL.n466 VTAIL.n465 13.1884
R476 VTAIL.n384 VTAIL.n383 13.1884
R477 VTAIL.n300 VTAIL.n299 13.1884
R478 VTAIL.n630 VTAIL.n598 12.8005
R479 VTAIL.n635 VTAIL.n596 12.8005
R480 VTAIL.n50 VTAIL.n18 12.8005
R481 VTAIL.n55 VTAIL.n16 12.8005
R482 VTAIL.n132 VTAIL.n100 12.8005
R483 VTAIL.n137 VTAIL.n98 12.8005
R484 VTAIL.n216 VTAIL.n184 12.8005
R485 VTAIL.n221 VTAIL.n182 12.8005
R486 VTAIL.n553 VTAIL.n514 12.8005
R487 VTAIL.n548 VTAIL.n516 12.8005
R488 VTAIL.n469 VTAIL.n430 12.8005
R489 VTAIL.n464 VTAIL.n432 12.8005
R490 VTAIL.n387 VTAIL.n348 12.8005
R491 VTAIL.n382 VTAIL.n350 12.8005
R492 VTAIL.n303 VTAIL.n264 12.8005
R493 VTAIL.n298 VTAIL.n266 12.8005
R494 VTAIL.n627 VTAIL.n626 12.0247
R495 VTAIL.n636 VTAIL.n594 12.0247
R496 VTAIL.n47 VTAIL.n46 12.0247
R497 VTAIL.n56 VTAIL.n14 12.0247
R498 VTAIL.n129 VTAIL.n128 12.0247
R499 VTAIL.n138 VTAIL.n96 12.0247
R500 VTAIL.n213 VTAIL.n212 12.0247
R501 VTAIL.n222 VTAIL.n180 12.0247
R502 VTAIL.n554 VTAIL.n512 12.0247
R503 VTAIL.n545 VTAIL.n544 12.0247
R504 VTAIL.n470 VTAIL.n428 12.0247
R505 VTAIL.n461 VTAIL.n460 12.0247
R506 VTAIL.n388 VTAIL.n346 12.0247
R507 VTAIL.n379 VTAIL.n378 12.0247
R508 VTAIL.n304 VTAIL.n262 12.0247
R509 VTAIL.n295 VTAIL.n294 12.0247
R510 VTAIL.n622 VTAIL.n600 11.249
R511 VTAIL.n640 VTAIL.n639 11.249
R512 VTAIL.n42 VTAIL.n20 11.249
R513 VTAIL.n60 VTAIL.n59 11.249
R514 VTAIL.n124 VTAIL.n102 11.249
R515 VTAIL.n142 VTAIL.n141 11.249
R516 VTAIL.n208 VTAIL.n186 11.249
R517 VTAIL.n226 VTAIL.n225 11.249
R518 VTAIL.n558 VTAIL.n557 11.249
R519 VTAIL.n541 VTAIL.n518 11.249
R520 VTAIL.n474 VTAIL.n473 11.249
R521 VTAIL.n457 VTAIL.n434 11.249
R522 VTAIL.n392 VTAIL.n391 11.249
R523 VTAIL.n375 VTAIL.n352 11.249
R524 VTAIL.n308 VTAIL.n307 11.249
R525 VTAIL.n291 VTAIL.n268 11.249
R526 VTAIL.n621 VTAIL.n602 10.4732
R527 VTAIL.n643 VTAIL.n592 10.4732
R528 VTAIL.n41 VTAIL.n22 10.4732
R529 VTAIL.n63 VTAIL.n12 10.4732
R530 VTAIL.n123 VTAIL.n104 10.4732
R531 VTAIL.n145 VTAIL.n94 10.4732
R532 VTAIL.n207 VTAIL.n188 10.4732
R533 VTAIL.n229 VTAIL.n178 10.4732
R534 VTAIL.n561 VTAIL.n510 10.4732
R535 VTAIL.n540 VTAIL.n521 10.4732
R536 VTAIL.n477 VTAIL.n426 10.4732
R537 VTAIL.n456 VTAIL.n437 10.4732
R538 VTAIL.n395 VTAIL.n344 10.4732
R539 VTAIL.n374 VTAIL.n355 10.4732
R540 VTAIL.n311 VTAIL.n260 10.4732
R541 VTAIL.n290 VTAIL.n271 10.4732
R542 VTAIL.n609 VTAIL.n607 10.2747
R543 VTAIL.n29 VTAIL.n27 10.2747
R544 VTAIL.n111 VTAIL.n109 10.2747
R545 VTAIL.n195 VTAIL.n193 10.2747
R546 VTAIL.n528 VTAIL.n526 10.2747
R547 VTAIL.n444 VTAIL.n442 10.2747
R548 VTAIL.n362 VTAIL.n360 10.2747
R549 VTAIL.n278 VTAIL.n276 10.2747
R550 VTAIL.n618 VTAIL.n617 9.69747
R551 VTAIL.n644 VTAIL.n590 9.69747
R552 VTAIL.n38 VTAIL.n37 9.69747
R553 VTAIL.n64 VTAIL.n10 9.69747
R554 VTAIL.n120 VTAIL.n119 9.69747
R555 VTAIL.n146 VTAIL.n92 9.69747
R556 VTAIL.n204 VTAIL.n203 9.69747
R557 VTAIL.n230 VTAIL.n176 9.69747
R558 VTAIL.n562 VTAIL.n508 9.69747
R559 VTAIL.n537 VTAIL.n536 9.69747
R560 VTAIL.n478 VTAIL.n424 9.69747
R561 VTAIL.n453 VTAIL.n452 9.69747
R562 VTAIL.n396 VTAIL.n342 9.69747
R563 VTAIL.n371 VTAIL.n370 9.69747
R564 VTAIL.n312 VTAIL.n258 9.69747
R565 VTAIL.n287 VTAIL.n286 9.69747
R566 VTAIL.n662 VTAIL.n661 9.45567
R567 VTAIL.n82 VTAIL.n81 9.45567
R568 VTAIL.n164 VTAIL.n163 9.45567
R569 VTAIL.n248 VTAIL.n247 9.45567
R570 VTAIL.n580 VTAIL.n579 9.45567
R571 VTAIL.n496 VTAIL.n495 9.45567
R572 VTAIL.n414 VTAIL.n413 9.45567
R573 VTAIL.n330 VTAIL.n329 9.45567
R574 VTAIL.n655 VTAIL.n654 9.3005
R575 VTAIL.n584 VTAIL.n583 9.3005
R576 VTAIL.n661 VTAIL.n660 9.3005
R577 VTAIL.n588 VTAIL.n587 9.3005
R578 VTAIL.n647 VTAIL.n646 9.3005
R579 VTAIL.n645 VTAIL.n644 9.3005
R580 VTAIL.n592 VTAIL.n591 9.3005
R581 VTAIL.n639 VTAIL.n638 9.3005
R582 VTAIL.n637 VTAIL.n636 9.3005
R583 VTAIL.n596 VTAIL.n595 9.3005
R584 VTAIL.n611 VTAIL.n610 9.3005
R585 VTAIL.n613 VTAIL.n612 9.3005
R586 VTAIL.n604 VTAIL.n603 9.3005
R587 VTAIL.n619 VTAIL.n618 9.3005
R588 VTAIL.n621 VTAIL.n620 9.3005
R589 VTAIL.n600 VTAIL.n599 9.3005
R590 VTAIL.n628 VTAIL.n627 9.3005
R591 VTAIL.n630 VTAIL.n629 9.3005
R592 VTAIL.n653 VTAIL.n652 9.3005
R593 VTAIL.n75 VTAIL.n74 9.3005
R594 VTAIL.n4 VTAIL.n3 9.3005
R595 VTAIL.n81 VTAIL.n80 9.3005
R596 VTAIL.n8 VTAIL.n7 9.3005
R597 VTAIL.n67 VTAIL.n66 9.3005
R598 VTAIL.n65 VTAIL.n64 9.3005
R599 VTAIL.n12 VTAIL.n11 9.3005
R600 VTAIL.n59 VTAIL.n58 9.3005
R601 VTAIL.n57 VTAIL.n56 9.3005
R602 VTAIL.n16 VTAIL.n15 9.3005
R603 VTAIL.n31 VTAIL.n30 9.3005
R604 VTAIL.n33 VTAIL.n32 9.3005
R605 VTAIL.n24 VTAIL.n23 9.3005
R606 VTAIL.n39 VTAIL.n38 9.3005
R607 VTAIL.n41 VTAIL.n40 9.3005
R608 VTAIL.n20 VTAIL.n19 9.3005
R609 VTAIL.n48 VTAIL.n47 9.3005
R610 VTAIL.n50 VTAIL.n49 9.3005
R611 VTAIL.n73 VTAIL.n72 9.3005
R612 VTAIL.n157 VTAIL.n156 9.3005
R613 VTAIL.n86 VTAIL.n85 9.3005
R614 VTAIL.n163 VTAIL.n162 9.3005
R615 VTAIL.n90 VTAIL.n89 9.3005
R616 VTAIL.n149 VTAIL.n148 9.3005
R617 VTAIL.n147 VTAIL.n146 9.3005
R618 VTAIL.n94 VTAIL.n93 9.3005
R619 VTAIL.n141 VTAIL.n140 9.3005
R620 VTAIL.n139 VTAIL.n138 9.3005
R621 VTAIL.n98 VTAIL.n97 9.3005
R622 VTAIL.n113 VTAIL.n112 9.3005
R623 VTAIL.n115 VTAIL.n114 9.3005
R624 VTAIL.n106 VTAIL.n105 9.3005
R625 VTAIL.n121 VTAIL.n120 9.3005
R626 VTAIL.n123 VTAIL.n122 9.3005
R627 VTAIL.n102 VTAIL.n101 9.3005
R628 VTAIL.n130 VTAIL.n129 9.3005
R629 VTAIL.n132 VTAIL.n131 9.3005
R630 VTAIL.n155 VTAIL.n154 9.3005
R631 VTAIL.n241 VTAIL.n240 9.3005
R632 VTAIL.n170 VTAIL.n169 9.3005
R633 VTAIL.n247 VTAIL.n246 9.3005
R634 VTAIL.n174 VTAIL.n173 9.3005
R635 VTAIL.n233 VTAIL.n232 9.3005
R636 VTAIL.n231 VTAIL.n230 9.3005
R637 VTAIL.n178 VTAIL.n177 9.3005
R638 VTAIL.n225 VTAIL.n224 9.3005
R639 VTAIL.n223 VTAIL.n222 9.3005
R640 VTAIL.n182 VTAIL.n181 9.3005
R641 VTAIL.n197 VTAIL.n196 9.3005
R642 VTAIL.n199 VTAIL.n198 9.3005
R643 VTAIL.n190 VTAIL.n189 9.3005
R644 VTAIL.n205 VTAIL.n204 9.3005
R645 VTAIL.n207 VTAIL.n206 9.3005
R646 VTAIL.n186 VTAIL.n185 9.3005
R647 VTAIL.n214 VTAIL.n213 9.3005
R648 VTAIL.n216 VTAIL.n215 9.3005
R649 VTAIL.n239 VTAIL.n238 9.3005
R650 VTAIL.n502 VTAIL.n501 9.3005
R651 VTAIL.n573 VTAIL.n572 9.3005
R652 VTAIL.n571 VTAIL.n570 9.3005
R653 VTAIL.n506 VTAIL.n505 9.3005
R654 VTAIL.n565 VTAIL.n564 9.3005
R655 VTAIL.n563 VTAIL.n562 9.3005
R656 VTAIL.n510 VTAIL.n509 9.3005
R657 VTAIL.n557 VTAIL.n556 9.3005
R658 VTAIL.n555 VTAIL.n554 9.3005
R659 VTAIL.n514 VTAIL.n513 9.3005
R660 VTAIL.n548 VTAIL.n547 9.3005
R661 VTAIL.n546 VTAIL.n545 9.3005
R662 VTAIL.n518 VTAIL.n517 9.3005
R663 VTAIL.n540 VTAIL.n539 9.3005
R664 VTAIL.n538 VTAIL.n537 9.3005
R665 VTAIL.n523 VTAIL.n522 9.3005
R666 VTAIL.n532 VTAIL.n531 9.3005
R667 VTAIL.n530 VTAIL.n529 9.3005
R668 VTAIL.n579 VTAIL.n578 9.3005
R669 VTAIL.n446 VTAIL.n445 9.3005
R670 VTAIL.n448 VTAIL.n447 9.3005
R671 VTAIL.n439 VTAIL.n438 9.3005
R672 VTAIL.n454 VTAIL.n453 9.3005
R673 VTAIL.n456 VTAIL.n455 9.3005
R674 VTAIL.n434 VTAIL.n433 9.3005
R675 VTAIL.n462 VTAIL.n461 9.3005
R676 VTAIL.n464 VTAIL.n463 9.3005
R677 VTAIL.n418 VTAIL.n417 9.3005
R678 VTAIL.n495 VTAIL.n494 9.3005
R679 VTAIL.n489 VTAIL.n488 9.3005
R680 VTAIL.n487 VTAIL.n486 9.3005
R681 VTAIL.n422 VTAIL.n421 9.3005
R682 VTAIL.n481 VTAIL.n480 9.3005
R683 VTAIL.n479 VTAIL.n478 9.3005
R684 VTAIL.n426 VTAIL.n425 9.3005
R685 VTAIL.n473 VTAIL.n472 9.3005
R686 VTAIL.n471 VTAIL.n470 9.3005
R687 VTAIL.n430 VTAIL.n429 9.3005
R688 VTAIL.n364 VTAIL.n363 9.3005
R689 VTAIL.n366 VTAIL.n365 9.3005
R690 VTAIL.n357 VTAIL.n356 9.3005
R691 VTAIL.n372 VTAIL.n371 9.3005
R692 VTAIL.n374 VTAIL.n373 9.3005
R693 VTAIL.n352 VTAIL.n351 9.3005
R694 VTAIL.n380 VTAIL.n379 9.3005
R695 VTAIL.n382 VTAIL.n381 9.3005
R696 VTAIL.n336 VTAIL.n335 9.3005
R697 VTAIL.n413 VTAIL.n412 9.3005
R698 VTAIL.n407 VTAIL.n406 9.3005
R699 VTAIL.n405 VTAIL.n404 9.3005
R700 VTAIL.n340 VTAIL.n339 9.3005
R701 VTAIL.n399 VTAIL.n398 9.3005
R702 VTAIL.n397 VTAIL.n396 9.3005
R703 VTAIL.n344 VTAIL.n343 9.3005
R704 VTAIL.n391 VTAIL.n390 9.3005
R705 VTAIL.n389 VTAIL.n388 9.3005
R706 VTAIL.n348 VTAIL.n347 9.3005
R707 VTAIL.n280 VTAIL.n279 9.3005
R708 VTAIL.n282 VTAIL.n281 9.3005
R709 VTAIL.n273 VTAIL.n272 9.3005
R710 VTAIL.n288 VTAIL.n287 9.3005
R711 VTAIL.n290 VTAIL.n289 9.3005
R712 VTAIL.n268 VTAIL.n267 9.3005
R713 VTAIL.n296 VTAIL.n295 9.3005
R714 VTAIL.n298 VTAIL.n297 9.3005
R715 VTAIL.n252 VTAIL.n251 9.3005
R716 VTAIL.n329 VTAIL.n328 9.3005
R717 VTAIL.n323 VTAIL.n322 9.3005
R718 VTAIL.n321 VTAIL.n320 9.3005
R719 VTAIL.n256 VTAIL.n255 9.3005
R720 VTAIL.n315 VTAIL.n314 9.3005
R721 VTAIL.n313 VTAIL.n312 9.3005
R722 VTAIL.n260 VTAIL.n259 9.3005
R723 VTAIL.n307 VTAIL.n306 9.3005
R724 VTAIL.n305 VTAIL.n304 9.3005
R725 VTAIL.n264 VTAIL.n263 9.3005
R726 VTAIL.n614 VTAIL.n604 8.92171
R727 VTAIL.n648 VTAIL.n647 8.92171
R728 VTAIL.n662 VTAIL.n582 8.92171
R729 VTAIL.n34 VTAIL.n24 8.92171
R730 VTAIL.n68 VTAIL.n67 8.92171
R731 VTAIL.n82 VTAIL.n2 8.92171
R732 VTAIL.n116 VTAIL.n106 8.92171
R733 VTAIL.n150 VTAIL.n149 8.92171
R734 VTAIL.n164 VTAIL.n84 8.92171
R735 VTAIL.n200 VTAIL.n190 8.92171
R736 VTAIL.n234 VTAIL.n233 8.92171
R737 VTAIL.n248 VTAIL.n168 8.92171
R738 VTAIL.n580 VTAIL.n500 8.92171
R739 VTAIL.n566 VTAIL.n565 8.92171
R740 VTAIL.n533 VTAIL.n523 8.92171
R741 VTAIL.n496 VTAIL.n416 8.92171
R742 VTAIL.n482 VTAIL.n481 8.92171
R743 VTAIL.n449 VTAIL.n439 8.92171
R744 VTAIL.n414 VTAIL.n334 8.92171
R745 VTAIL.n400 VTAIL.n399 8.92171
R746 VTAIL.n367 VTAIL.n357 8.92171
R747 VTAIL.n330 VTAIL.n250 8.92171
R748 VTAIL.n316 VTAIL.n315 8.92171
R749 VTAIL.n283 VTAIL.n273 8.92171
R750 VTAIL.n613 VTAIL.n606 8.14595
R751 VTAIL.n651 VTAIL.n588 8.14595
R752 VTAIL.n660 VTAIL.n659 8.14595
R753 VTAIL.n33 VTAIL.n26 8.14595
R754 VTAIL.n71 VTAIL.n8 8.14595
R755 VTAIL.n80 VTAIL.n79 8.14595
R756 VTAIL.n115 VTAIL.n108 8.14595
R757 VTAIL.n153 VTAIL.n90 8.14595
R758 VTAIL.n162 VTAIL.n161 8.14595
R759 VTAIL.n199 VTAIL.n192 8.14595
R760 VTAIL.n237 VTAIL.n174 8.14595
R761 VTAIL.n246 VTAIL.n245 8.14595
R762 VTAIL.n578 VTAIL.n577 8.14595
R763 VTAIL.n569 VTAIL.n506 8.14595
R764 VTAIL.n532 VTAIL.n525 8.14595
R765 VTAIL.n494 VTAIL.n493 8.14595
R766 VTAIL.n485 VTAIL.n422 8.14595
R767 VTAIL.n448 VTAIL.n441 8.14595
R768 VTAIL.n412 VTAIL.n411 8.14595
R769 VTAIL.n403 VTAIL.n340 8.14595
R770 VTAIL.n366 VTAIL.n359 8.14595
R771 VTAIL.n328 VTAIL.n327 8.14595
R772 VTAIL.n319 VTAIL.n256 8.14595
R773 VTAIL.n282 VTAIL.n275 8.14595
R774 VTAIL.n610 VTAIL.n609 7.3702
R775 VTAIL.n652 VTAIL.n586 7.3702
R776 VTAIL.n656 VTAIL.n584 7.3702
R777 VTAIL.n30 VTAIL.n29 7.3702
R778 VTAIL.n72 VTAIL.n6 7.3702
R779 VTAIL.n76 VTAIL.n4 7.3702
R780 VTAIL.n112 VTAIL.n111 7.3702
R781 VTAIL.n154 VTAIL.n88 7.3702
R782 VTAIL.n158 VTAIL.n86 7.3702
R783 VTAIL.n196 VTAIL.n195 7.3702
R784 VTAIL.n238 VTAIL.n172 7.3702
R785 VTAIL.n242 VTAIL.n170 7.3702
R786 VTAIL.n574 VTAIL.n502 7.3702
R787 VTAIL.n570 VTAIL.n504 7.3702
R788 VTAIL.n529 VTAIL.n528 7.3702
R789 VTAIL.n490 VTAIL.n418 7.3702
R790 VTAIL.n486 VTAIL.n420 7.3702
R791 VTAIL.n445 VTAIL.n444 7.3702
R792 VTAIL.n408 VTAIL.n336 7.3702
R793 VTAIL.n404 VTAIL.n338 7.3702
R794 VTAIL.n363 VTAIL.n362 7.3702
R795 VTAIL.n324 VTAIL.n252 7.3702
R796 VTAIL.n320 VTAIL.n254 7.3702
R797 VTAIL.n279 VTAIL.n278 7.3702
R798 VTAIL.n655 VTAIL.n586 6.59444
R799 VTAIL.n656 VTAIL.n655 6.59444
R800 VTAIL.n75 VTAIL.n6 6.59444
R801 VTAIL.n76 VTAIL.n75 6.59444
R802 VTAIL.n157 VTAIL.n88 6.59444
R803 VTAIL.n158 VTAIL.n157 6.59444
R804 VTAIL.n241 VTAIL.n172 6.59444
R805 VTAIL.n242 VTAIL.n241 6.59444
R806 VTAIL.n574 VTAIL.n573 6.59444
R807 VTAIL.n573 VTAIL.n504 6.59444
R808 VTAIL.n490 VTAIL.n489 6.59444
R809 VTAIL.n489 VTAIL.n420 6.59444
R810 VTAIL.n408 VTAIL.n407 6.59444
R811 VTAIL.n407 VTAIL.n338 6.59444
R812 VTAIL.n324 VTAIL.n323 6.59444
R813 VTAIL.n323 VTAIL.n254 6.59444
R814 VTAIL.n610 VTAIL.n606 5.81868
R815 VTAIL.n652 VTAIL.n651 5.81868
R816 VTAIL.n659 VTAIL.n584 5.81868
R817 VTAIL.n30 VTAIL.n26 5.81868
R818 VTAIL.n72 VTAIL.n71 5.81868
R819 VTAIL.n79 VTAIL.n4 5.81868
R820 VTAIL.n112 VTAIL.n108 5.81868
R821 VTAIL.n154 VTAIL.n153 5.81868
R822 VTAIL.n161 VTAIL.n86 5.81868
R823 VTAIL.n196 VTAIL.n192 5.81868
R824 VTAIL.n238 VTAIL.n237 5.81868
R825 VTAIL.n245 VTAIL.n170 5.81868
R826 VTAIL.n577 VTAIL.n502 5.81868
R827 VTAIL.n570 VTAIL.n569 5.81868
R828 VTAIL.n529 VTAIL.n525 5.81868
R829 VTAIL.n493 VTAIL.n418 5.81868
R830 VTAIL.n486 VTAIL.n485 5.81868
R831 VTAIL.n445 VTAIL.n441 5.81868
R832 VTAIL.n411 VTAIL.n336 5.81868
R833 VTAIL.n404 VTAIL.n403 5.81868
R834 VTAIL.n363 VTAIL.n359 5.81868
R835 VTAIL.n327 VTAIL.n252 5.81868
R836 VTAIL.n320 VTAIL.n319 5.81868
R837 VTAIL.n279 VTAIL.n275 5.81868
R838 VTAIL.n614 VTAIL.n613 5.04292
R839 VTAIL.n648 VTAIL.n588 5.04292
R840 VTAIL.n660 VTAIL.n582 5.04292
R841 VTAIL.n34 VTAIL.n33 5.04292
R842 VTAIL.n68 VTAIL.n8 5.04292
R843 VTAIL.n80 VTAIL.n2 5.04292
R844 VTAIL.n116 VTAIL.n115 5.04292
R845 VTAIL.n150 VTAIL.n90 5.04292
R846 VTAIL.n162 VTAIL.n84 5.04292
R847 VTAIL.n200 VTAIL.n199 5.04292
R848 VTAIL.n234 VTAIL.n174 5.04292
R849 VTAIL.n246 VTAIL.n168 5.04292
R850 VTAIL.n578 VTAIL.n500 5.04292
R851 VTAIL.n566 VTAIL.n506 5.04292
R852 VTAIL.n533 VTAIL.n532 5.04292
R853 VTAIL.n494 VTAIL.n416 5.04292
R854 VTAIL.n482 VTAIL.n422 5.04292
R855 VTAIL.n449 VTAIL.n448 5.04292
R856 VTAIL.n412 VTAIL.n334 5.04292
R857 VTAIL.n400 VTAIL.n340 5.04292
R858 VTAIL.n367 VTAIL.n366 5.04292
R859 VTAIL.n328 VTAIL.n250 5.04292
R860 VTAIL.n316 VTAIL.n256 5.04292
R861 VTAIL.n283 VTAIL.n282 5.04292
R862 VTAIL.n617 VTAIL.n604 4.26717
R863 VTAIL.n647 VTAIL.n590 4.26717
R864 VTAIL.n37 VTAIL.n24 4.26717
R865 VTAIL.n67 VTAIL.n10 4.26717
R866 VTAIL.n119 VTAIL.n106 4.26717
R867 VTAIL.n149 VTAIL.n92 4.26717
R868 VTAIL.n203 VTAIL.n190 4.26717
R869 VTAIL.n233 VTAIL.n176 4.26717
R870 VTAIL.n565 VTAIL.n508 4.26717
R871 VTAIL.n536 VTAIL.n523 4.26717
R872 VTAIL.n481 VTAIL.n424 4.26717
R873 VTAIL.n452 VTAIL.n439 4.26717
R874 VTAIL.n399 VTAIL.n342 4.26717
R875 VTAIL.n370 VTAIL.n357 4.26717
R876 VTAIL.n315 VTAIL.n258 4.26717
R877 VTAIL.n286 VTAIL.n273 4.26717
R878 VTAIL.n618 VTAIL.n602 3.49141
R879 VTAIL.n644 VTAIL.n643 3.49141
R880 VTAIL.n38 VTAIL.n22 3.49141
R881 VTAIL.n64 VTAIL.n63 3.49141
R882 VTAIL.n120 VTAIL.n104 3.49141
R883 VTAIL.n146 VTAIL.n145 3.49141
R884 VTAIL.n204 VTAIL.n188 3.49141
R885 VTAIL.n230 VTAIL.n229 3.49141
R886 VTAIL.n562 VTAIL.n561 3.49141
R887 VTAIL.n537 VTAIL.n521 3.49141
R888 VTAIL.n478 VTAIL.n477 3.49141
R889 VTAIL.n453 VTAIL.n437 3.49141
R890 VTAIL.n396 VTAIL.n395 3.49141
R891 VTAIL.n371 VTAIL.n355 3.49141
R892 VTAIL.n312 VTAIL.n311 3.49141
R893 VTAIL.n287 VTAIL.n271 3.49141
R894 VTAIL.n333 VTAIL.n331 2.97464
R895 VTAIL.n415 VTAIL.n333 2.97464
R896 VTAIL.n499 VTAIL.n497 2.97464
R897 VTAIL.n581 VTAIL.n499 2.97464
R898 VTAIL.n249 VTAIL.n167 2.97464
R899 VTAIL.n167 VTAIL.n165 2.97464
R900 VTAIL.n83 VTAIL.n1 2.97464
R901 VTAIL VTAIL.n663 2.91645
R902 VTAIL.n611 VTAIL.n607 2.84303
R903 VTAIL.n31 VTAIL.n27 2.84303
R904 VTAIL.n113 VTAIL.n109 2.84303
R905 VTAIL.n197 VTAIL.n193 2.84303
R906 VTAIL.n530 VTAIL.n526 2.84303
R907 VTAIL.n446 VTAIL.n442 2.84303
R908 VTAIL.n364 VTAIL.n360 2.84303
R909 VTAIL.n280 VTAIL.n276 2.84303
R910 VTAIL.n622 VTAIL.n621 2.71565
R911 VTAIL.n640 VTAIL.n592 2.71565
R912 VTAIL.n42 VTAIL.n41 2.71565
R913 VTAIL.n60 VTAIL.n12 2.71565
R914 VTAIL.n124 VTAIL.n123 2.71565
R915 VTAIL.n142 VTAIL.n94 2.71565
R916 VTAIL.n208 VTAIL.n207 2.71565
R917 VTAIL.n226 VTAIL.n178 2.71565
R918 VTAIL.n558 VTAIL.n510 2.71565
R919 VTAIL.n541 VTAIL.n540 2.71565
R920 VTAIL.n474 VTAIL.n426 2.71565
R921 VTAIL.n457 VTAIL.n456 2.71565
R922 VTAIL.n392 VTAIL.n344 2.71565
R923 VTAIL.n375 VTAIL.n374 2.71565
R924 VTAIL.n308 VTAIL.n260 2.71565
R925 VTAIL.n291 VTAIL.n290 2.71565
R926 VTAIL.n626 VTAIL.n600 1.93989
R927 VTAIL.n639 VTAIL.n594 1.93989
R928 VTAIL.n46 VTAIL.n20 1.93989
R929 VTAIL.n59 VTAIL.n14 1.93989
R930 VTAIL.n128 VTAIL.n102 1.93989
R931 VTAIL.n141 VTAIL.n96 1.93989
R932 VTAIL.n212 VTAIL.n186 1.93989
R933 VTAIL.n225 VTAIL.n180 1.93989
R934 VTAIL.n557 VTAIL.n512 1.93989
R935 VTAIL.n544 VTAIL.n518 1.93989
R936 VTAIL.n473 VTAIL.n428 1.93989
R937 VTAIL.n460 VTAIL.n434 1.93989
R938 VTAIL.n391 VTAIL.n346 1.93989
R939 VTAIL.n378 VTAIL.n352 1.93989
R940 VTAIL.n307 VTAIL.n262 1.93989
R941 VTAIL.n294 VTAIL.n268 1.93989
R942 VTAIL.n0 VTAIL.t3 1.32669
R943 VTAIL.n0 VTAIL.t5 1.32669
R944 VTAIL.n166 VTAIL.t9 1.32669
R945 VTAIL.n166 VTAIL.t6 1.32669
R946 VTAIL.n498 VTAIL.t13 1.32669
R947 VTAIL.n498 VTAIL.t12 1.32669
R948 VTAIL.n332 VTAIL.t4 1.32669
R949 VTAIL.n332 VTAIL.t1 1.32669
R950 VTAIL.n627 VTAIL.n598 1.16414
R951 VTAIL.n636 VTAIL.n635 1.16414
R952 VTAIL.n47 VTAIL.n18 1.16414
R953 VTAIL.n56 VTAIL.n55 1.16414
R954 VTAIL.n129 VTAIL.n100 1.16414
R955 VTAIL.n138 VTAIL.n137 1.16414
R956 VTAIL.n213 VTAIL.n184 1.16414
R957 VTAIL.n222 VTAIL.n221 1.16414
R958 VTAIL.n554 VTAIL.n553 1.16414
R959 VTAIL.n545 VTAIL.n516 1.16414
R960 VTAIL.n470 VTAIL.n469 1.16414
R961 VTAIL.n461 VTAIL.n432 1.16414
R962 VTAIL.n388 VTAIL.n387 1.16414
R963 VTAIL.n379 VTAIL.n350 1.16414
R964 VTAIL.n304 VTAIL.n303 1.16414
R965 VTAIL.n295 VTAIL.n266 1.16414
R966 VTAIL.n497 VTAIL.n415 0.470328
R967 VTAIL.n165 VTAIL.n83 0.470328
R968 VTAIL.n631 VTAIL.n630 0.388379
R969 VTAIL.n632 VTAIL.n596 0.388379
R970 VTAIL.n51 VTAIL.n50 0.388379
R971 VTAIL.n52 VTAIL.n16 0.388379
R972 VTAIL.n133 VTAIL.n132 0.388379
R973 VTAIL.n134 VTAIL.n98 0.388379
R974 VTAIL.n217 VTAIL.n216 0.388379
R975 VTAIL.n218 VTAIL.n182 0.388379
R976 VTAIL.n550 VTAIL.n514 0.388379
R977 VTAIL.n549 VTAIL.n548 0.388379
R978 VTAIL.n466 VTAIL.n430 0.388379
R979 VTAIL.n465 VTAIL.n464 0.388379
R980 VTAIL.n384 VTAIL.n348 0.388379
R981 VTAIL.n383 VTAIL.n382 0.388379
R982 VTAIL.n300 VTAIL.n264 0.388379
R983 VTAIL.n299 VTAIL.n298 0.388379
R984 VTAIL.n612 VTAIL.n611 0.155672
R985 VTAIL.n612 VTAIL.n603 0.155672
R986 VTAIL.n619 VTAIL.n603 0.155672
R987 VTAIL.n620 VTAIL.n619 0.155672
R988 VTAIL.n620 VTAIL.n599 0.155672
R989 VTAIL.n628 VTAIL.n599 0.155672
R990 VTAIL.n629 VTAIL.n628 0.155672
R991 VTAIL.n629 VTAIL.n595 0.155672
R992 VTAIL.n637 VTAIL.n595 0.155672
R993 VTAIL.n638 VTAIL.n637 0.155672
R994 VTAIL.n638 VTAIL.n591 0.155672
R995 VTAIL.n645 VTAIL.n591 0.155672
R996 VTAIL.n646 VTAIL.n645 0.155672
R997 VTAIL.n646 VTAIL.n587 0.155672
R998 VTAIL.n653 VTAIL.n587 0.155672
R999 VTAIL.n654 VTAIL.n653 0.155672
R1000 VTAIL.n654 VTAIL.n583 0.155672
R1001 VTAIL.n661 VTAIL.n583 0.155672
R1002 VTAIL.n32 VTAIL.n31 0.155672
R1003 VTAIL.n32 VTAIL.n23 0.155672
R1004 VTAIL.n39 VTAIL.n23 0.155672
R1005 VTAIL.n40 VTAIL.n39 0.155672
R1006 VTAIL.n40 VTAIL.n19 0.155672
R1007 VTAIL.n48 VTAIL.n19 0.155672
R1008 VTAIL.n49 VTAIL.n48 0.155672
R1009 VTAIL.n49 VTAIL.n15 0.155672
R1010 VTAIL.n57 VTAIL.n15 0.155672
R1011 VTAIL.n58 VTAIL.n57 0.155672
R1012 VTAIL.n58 VTAIL.n11 0.155672
R1013 VTAIL.n65 VTAIL.n11 0.155672
R1014 VTAIL.n66 VTAIL.n65 0.155672
R1015 VTAIL.n66 VTAIL.n7 0.155672
R1016 VTAIL.n73 VTAIL.n7 0.155672
R1017 VTAIL.n74 VTAIL.n73 0.155672
R1018 VTAIL.n74 VTAIL.n3 0.155672
R1019 VTAIL.n81 VTAIL.n3 0.155672
R1020 VTAIL.n114 VTAIL.n113 0.155672
R1021 VTAIL.n114 VTAIL.n105 0.155672
R1022 VTAIL.n121 VTAIL.n105 0.155672
R1023 VTAIL.n122 VTAIL.n121 0.155672
R1024 VTAIL.n122 VTAIL.n101 0.155672
R1025 VTAIL.n130 VTAIL.n101 0.155672
R1026 VTAIL.n131 VTAIL.n130 0.155672
R1027 VTAIL.n131 VTAIL.n97 0.155672
R1028 VTAIL.n139 VTAIL.n97 0.155672
R1029 VTAIL.n140 VTAIL.n139 0.155672
R1030 VTAIL.n140 VTAIL.n93 0.155672
R1031 VTAIL.n147 VTAIL.n93 0.155672
R1032 VTAIL.n148 VTAIL.n147 0.155672
R1033 VTAIL.n148 VTAIL.n89 0.155672
R1034 VTAIL.n155 VTAIL.n89 0.155672
R1035 VTAIL.n156 VTAIL.n155 0.155672
R1036 VTAIL.n156 VTAIL.n85 0.155672
R1037 VTAIL.n163 VTAIL.n85 0.155672
R1038 VTAIL.n198 VTAIL.n197 0.155672
R1039 VTAIL.n198 VTAIL.n189 0.155672
R1040 VTAIL.n205 VTAIL.n189 0.155672
R1041 VTAIL.n206 VTAIL.n205 0.155672
R1042 VTAIL.n206 VTAIL.n185 0.155672
R1043 VTAIL.n214 VTAIL.n185 0.155672
R1044 VTAIL.n215 VTAIL.n214 0.155672
R1045 VTAIL.n215 VTAIL.n181 0.155672
R1046 VTAIL.n223 VTAIL.n181 0.155672
R1047 VTAIL.n224 VTAIL.n223 0.155672
R1048 VTAIL.n224 VTAIL.n177 0.155672
R1049 VTAIL.n231 VTAIL.n177 0.155672
R1050 VTAIL.n232 VTAIL.n231 0.155672
R1051 VTAIL.n232 VTAIL.n173 0.155672
R1052 VTAIL.n239 VTAIL.n173 0.155672
R1053 VTAIL.n240 VTAIL.n239 0.155672
R1054 VTAIL.n240 VTAIL.n169 0.155672
R1055 VTAIL.n247 VTAIL.n169 0.155672
R1056 VTAIL.n579 VTAIL.n501 0.155672
R1057 VTAIL.n572 VTAIL.n501 0.155672
R1058 VTAIL.n572 VTAIL.n571 0.155672
R1059 VTAIL.n571 VTAIL.n505 0.155672
R1060 VTAIL.n564 VTAIL.n505 0.155672
R1061 VTAIL.n564 VTAIL.n563 0.155672
R1062 VTAIL.n563 VTAIL.n509 0.155672
R1063 VTAIL.n556 VTAIL.n509 0.155672
R1064 VTAIL.n556 VTAIL.n555 0.155672
R1065 VTAIL.n555 VTAIL.n513 0.155672
R1066 VTAIL.n547 VTAIL.n513 0.155672
R1067 VTAIL.n547 VTAIL.n546 0.155672
R1068 VTAIL.n546 VTAIL.n517 0.155672
R1069 VTAIL.n539 VTAIL.n517 0.155672
R1070 VTAIL.n539 VTAIL.n538 0.155672
R1071 VTAIL.n538 VTAIL.n522 0.155672
R1072 VTAIL.n531 VTAIL.n522 0.155672
R1073 VTAIL.n531 VTAIL.n530 0.155672
R1074 VTAIL.n495 VTAIL.n417 0.155672
R1075 VTAIL.n488 VTAIL.n417 0.155672
R1076 VTAIL.n488 VTAIL.n487 0.155672
R1077 VTAIL.n487 VTAIL.n421 0.155672
R1078 VTAIL.n480 VTAIL.n421 0.155672
R1079 VTAIL.n480 VTAIL.n479 0.155672
R1080 VTAIL.n479 VTAIL.n425 0.155672
R1081 VTAIL.n472 VTAIL.n425 0.155672
R1082 VTAIL.n472 VTAIL.n471 0.155672
R1083 VTAIL.n471 VTAIL.n429 0.155672
R1084 VTAIL.n463 VTAIL.n429 0.155672
R1085 VTAIL.n463 VTAIL.n462 0.155672
R1086 VTAIL.n462 VTAIL.n433 0.155672
R1087 VTAIL.n455 VTAIL.n433 0.155672
R1088 VTAIL.n455 VTAIL.n454 0.155672
R1089 VTAIL.n454 VTAIL.n438 0.155672
R1090 VTAIL.n447 VTAIL.n438 0.155672
R1091 VTAIL.n447 VTAIL.n446 0.155672
R1092 VTAIL.n413 VTAIL.n335 0.155672
R1093 VTAIL.n406 VTAIL.n335 0.155672
R1094 VTAIL.n406 VTAIL.n405 0.155672
R1095 VTAIL.n405 VTAIL.n339 0.155672
R1096 VTAIL.n398 VTAIL.n339 0.155672
R1097 VTAIL.n398 VTAIL.n397 0.155672
R1098 VTAIL.n397 VTAIL.n343 0.155672
R1099 VTAIL.n390 VTAIL.n343 0.155672
R1100 VTAIL.n390 VTAIL.n389 0.155672
R1101 VTAIL.n389 VTAIL.n347 0.155672
R1102 VTAIL.n381 VTAIL.n347 0.155672
R1103 VTAIL.n381 VTAIL.n380 0.155672
R1104 VTAIL.n380 VTAIL.n351 0.155672
R1105 VTAIL.n373 VTAIL.n351 0.155672
R1106 VTAIL.n373 VTAIL.n372 0.155672
R1107 VTAIL.n372 VTAIL.n356 0.155672
R1108 VTAIL.n365 VTAIL.n356 0.155672
R1109 VTAIL.n365 VTAIL.n364 0.155672
R1110 VTAIL.n329 VTAIL.n251 0.155672
R1111 VTAIL.n322 VTAIL.n251 0.155672
R1112 VTAIL.n322 VTAIL.n321 0.155672
R1113 VTAIL.n321 VTAIL.n255 0.155672
R1114 VTAIL.n314 VTAIL.n255 0.155672
R1115 VTAIL.n314 VTAIL.n313 0.155672
R1116 VTAIL.n313 VTAIL.n259 0.155672
R1117 VTAIL.n306 VTAIL.n259 0.155672
R1118 VTAIL.n306 VTAIL.n305 0.155672
R1119 VTAIL.n305 VTAIL.n263 0.155672
R1120 VTAIL.n297 VTAIL.n263 0.155672
R1121 VTAIL.n297 VTAIL.n296 0.155672
R1122 VTAIL.n296 VTAIL.n267 0.155672
R1123 VTAIL.n289 VTAIL.n267 0.155672
R1124 VTAIL.n289 VTAIL.n288 0.155672
R1125 VTAIL.n288 VTAIL.n272 0.155672
R1126 VTAIL.n281 VTAIL.n272 0.155672
R1127 VTAIL.n281 VTAIL.n280 0.155672
R1128 VTAIL VTAIL.n1 0.0586897
R1129 VDD1 VDD1.n0 61.5093
R1130 VDD1.n3 VDD1.n2 61.3956
R1131 VDD1.n3 VDD1.n1 61.3956
R1132 VDD1.n5 VDD1.n4 59.9641
R1133 VDD1.n5 VDD1.n3 50.5526
R1134 VDD1 VDD1.n5 1.42938
R1135 VDD1.n4 VDD1.t1 1.32669
R1136 VDD1.n4 VDD1.t4 1.32669
R1137 VDD1.n0 VDD1.t0 1.32669
R1138 VDD1.n0 VDD1.t7 1.32669
R1139 VDD1.n2 VDD1.t2 1.32669
R1140 VDD1.n2 VDD1.t6 1.32669
R1141 VDD1.n1 VDD1.t3 1.32669
R1142 VDD1.n1 VDD1.t5 1.32669
R1143 B.n1032 B.n1031 585
R1144 B.n383 B.n163 585
R1145 B.n382 B.n381 585
R1146 B.n380 B.n379 585
R1147 B.n378 B.n377 585
R1148 B.n376 B.n375 585
R1149 B.n374 B.n373 585
R1150 B.n372 B.n371 585
R1151 B.n370 B.n369 585
R1152 B.n368 B.n367 585
R1153 B.n366 B.n365 585
R1154 B.n364 B.n363 585
R1155 B.n362 B.n361 585
R1156 B.n360 B.n359 585
R1157 B.n358 B.n357 585
R1158 B.n356 B.n355 585
R1159 B.n354 B.n353 585
R1160 B.n352 B.n351 585
R1161 B.n350 B.n349 585
R1162 B.n348 B.n347 585
R1163 B.n346 B.n345 585
R1164 B.n344 B.n343 585
R1165 B.n342 B.n341 585
R1166 B.n340 B.n339 585
R1167 B.n338 B.n337 585
R1168 B.n336 B.n335 585
R1169 B.n334 B.n333 585
R1170 B.n332 B.n331 585
R1171 B.n330 B.n329 585
R1172 B.n328 B.n327 585
R1173 B.n326 B.n325 585
R1174 B.n324 B.n323 585
R1175 B.n322 B.n321 585
R1176 B.n320 B.n319 585
R1177 B.n318 B.n317 585
R1178 B.n316 B.n315 585
R1179 B.n314 B.n313 585
R1180 B.n312 B.n311 585
R1181 B.n310 B.n309 585
R1182 B.n308 B.n307 585
R1183 B.n306 B.n305 585
R1184 B.n304 B.n303 585
R1185 B.n302 B.n301 585
R1186 B.n300 B.n299 585
R1187 B.n298 B.n297 585
R1188 B.n296 B.n295 585
R1189 B.n294 B.n293 585
R1190 B.n292 B.n291 585
R1191 B.n290 B.n289 585
R1192 B.n288 B.n287 585
R1193 B.n286 B.n285 585
R1194 B.n284 B.n283 585
R1195 B.n282 B.n281 585
R1196 B.n280 B.n279 585
R1197 B.n278 B.n277 585
R1198 B.n276 B.n275 585
R1199 B.n274 B.n273 585
R1200 B.n272 B.n271 585
R1201 B.n270 B.n269 585
R1202 B.n268 B.n267 585
R1203 B.n266 B.n265 585
R1204 B.n264 B.n263 585
R1205 B.n262 B.n261 585
R1206 B.n260 B.n259 585
R1207 B.n258 B.n257 585
R1208 B.n256 B.n255 585
R1209 B.n254 B.n253 585
R1210 B.n252 B.n251 585
R1211 B.n250 B.n249 585
R1212 B.n248 B.n247 585
R1213 B.n246 B.n245 585
R1214 B.n244 B.n243 585
R1215 B.n242 B.n241 585
R1216 B.n240 B.n239 585
R1217 B.n238 B.n237 585
R1218 B.n236 B.n235 585
R1219 B.n234 B.n233 585
R1220 B.n232 B.n231 585
R1221 B.n230 B.n229 585
R1222 B.n228 B.n227 585
R1223 B.n226 B.n225 585
R1224 B.n224 B.n223 585
R1225 B.n222 B.n221 585
R1226 B.n220 B.n219 585
R1227 B.n218 B.n217 585
R1228 B.n216 B.n215 585
R1229 B.n214 B.n213 585
R1230 B.n212 B.n211 585
R1231 B.n210 B.n209 585
R1232 B.n208 B.n207 585
R1233 B.n206 B.n205 585
R1234 B.n204 B.n203 585
R1235 B.n202 B.n201 585
R1236 B.n200 B.n199 585
R1237 B.n198 B.n197 585
R1238 B.n196 B.n195 585
R1239 B.n194 B.n193 585
R1240 B.n192 B.n191 585
R1241 B.n190 B.n189 585
R1242 B.n188 B.n187 585
R1243 B.n186 B.n185 585
R1244 B.n184 B.n183 585
R1245 B.n182 B.n181 585
R1246 B.n180 B.n179 585
R1247 B.n178 B.n177 585
R1248 B.n176 B.n175 585
R1249 B.n174 B.n173 585
R1250 B.n172 B.n171 585
R1251 B.n109 B.n108 585
R1252 B.n1037 B.n1036 585
R1253 B.n1030 B.n164 585
R1254 B.n164 B.n106 585
R1255 B.n1029 B.n105 585
R1256 B.n1041 B.n105 585
R1257 B.n1028 B.n104 585
R1258 B.n1042 B.n104 585
R1259 B.n1027 B.n103 585
R1260 B.n1043 B.n103 585
R1261 B.n1026 B.n1025 585
R1262 B.n1025 B.n99 585
R1263 B.n1024 B.n98 585
R1264 B.n1049 B.n98 585
R1265 B.n1023 B.n97 585
R1266 B.n1050 B.n97 585
R1267 B.n1022 B.n96 585
R1268 B.n1051 B.n96 585
R1269 B.n1021 B.n1020 585
R1270 B.n1020 B.n95 585
R1271 B.n1019 B.n91 585
R1272 B.n1057 B.n91 585
R1273 B.n1018 B.n90 585
R1274 B.n1058 B.n90 585
R1275 B.n1017 B.n89 585
R1276 B.n1059 B.n89 585
R1277 B.n1016 B.n1015 585
R1278 B.n1015 B.n85 585
R1279 B.n1014 B.n84 585
R1280 B.n1065 B.n84 585
R1281 B.n1013 B.n83 585
R1282 B.n1066 B.n83 585
R1283 B.n1012 B.n82 585
R1284 B.n1067 B.n82 585
R1285 B.n1011 B.n1010 585
R1286 B.n1010 B.n78 585
R1287 B.n1009 B.n77 585
R1288 B.n1073 B.n77 585
R1289 B.n1008 B.n76 585
R1290 B.n1074 B.n76 585
R1291 B.n1007 B.n75 585
R1292 B.n1075 B.n75 585
R1293 B.n1006 B.n1005 585
R1294 B.n1005 B.n71 585
R1295 B.n1004 B.n70 585
R1296 B.n1081 B.n70 585
R1297 B.n1003 B.n69 585
R1298 B.n1082 B.n69 585
R1299 B.n1002 B.n68 585
R1300 B.n1083 B.n68 585
R1301 B.n1001 B.n1000 585
R1302 B.n1000 B.n64 585
R1303 B.n999 B.n63 585
R1304 B.n1089 B.n63 585
R1305 B.n998 B.n62 585
R1306 B.n1090 B.n62 585
R1307 B.n997 B.n61 585
R1308 B.n1091 B.n61 585
R1309 B.n996 B.n995 585
R1310 B.n995 B.n57 585
R1311 B.n994 B.n56 585
R1312 B.n1097 B.n56 585
R1313 B.n993 B.n55 585
R1314 B.n1098 B.n55 585
R1315 B.n992 B.n54 585
R1316 B.n1099 B.n54 585
R1317 B.n991 B.n990 585
R1318 B.n990 B.n53 585
R1319 B.n989 B.n49 585
R1320 B.n1105 B.n49 585
R1321 B.n988 B.n48 585
R1322 B.n1106 B.n48 585
R1323 B.n987 B.n47 585
R1324 B.n1107 B.n47 585
R1325 B.n986 B.n985 585
R1326 B.n985 B.n43 585
R1327 B.n984 B.n42 585
R1328 B.n1113 B.n42 585
R1329 B.n983 B.n41 585
R1330 B.n1114 B.n41 585
R1331 B.n982 B.n40 585
R1332 B.n1115 B.n40 585
R1333 B.n981 B.n980 585
R1334 B.n980 B.n36 585
R1335 B.n979 B.n35 585
R1336 B.n1121 B.n35 585
R1337 B.n978 B.n34 585
R1338 B.n1122 B.n34 585
R1339 B.n977 B.n33 585
R1340 B.n1123 B.n33 585
R1341 B.n976 B.n975 585
R1342 B.n975 B.n29 585
R1343 B.n974 B.n28 585
R1344 B.n1129 B.n28 585
R1345 B.n973 B.n27 585
R1346 B.n1130 B.n27 585
R1347 B.n972 B.n26 585
R1348 B.n1131 B.n26 585
R1349 B.n971 B.n970 585
R1350 B.n970 B.n22 585
R1351 B.n969 B.n21 585
R1352 B.n1137 B.n21 585
R1353 B.n968 B.n20 585
R1354 B.n1138 B.n20 585
R1355 B.n967 B.n19 585
R1356 B.n1139 B.n19 585
R1357 B.n966 B.n965 585
R1358 B.n965 B.n18 585
R1359 B.n964 B.n14 585
R1360 B.n1145 B.n14 585
R1361 B.n963 B.n13 585
R1362 B.n1146 B.n13 585
R1363 B.n962 B.n12 585
R1364 B.n1147 B.n12 585
R1365 B.n961 B.n960 585
R1366 B.n960 B.n8 585
R1367 B.n959 B.n7 585
R1368 B.n1153 B.n7 585
R1369 B.n958 B.n6 585
R1370 B.n1154 B.n6 585
R1371 B.n957 B.n5 585
R1372 B.n1155 B.n5 585
R1373 B.n956 B.n955 585
R1374 B.n955 B.n4 585
R1375 B.n954 B.n384 585
R1376 B.n954 B.n953 585
R1377 B.n944 B.n385 585
R1378 B.n386 B.n385 585
R1379 B.n946 B.n945 585
R1380 B.n947 B.n946 585
R1381 B.n943 B.n391 585
R1382 B.n391 B.n390 585
R1383 B.n942 B.n941 585
R1384 B.n941 B.n940 585
R1385 B.n393 B.n392 585
R1386 B.n933 B.n393 585
R1387 B.n932 B.n931 585
R1388 B.n934 B.n932 585
R1389 B.n930 B.n398 585
R1390 B.n398 B.n397 585
R1391 B.n929 B.n928 585
R1392 B.n928 B.n927 585
R1393 B.n400 B.n399 585
R1394 B.n401 B.n400 585
R1395 B.n920 B.n919 585
R1396 B.n921 B.n920 585
R1397 B.n918 B.n406 585
R1398 B.n406 B.n405 585
R1399 B.n917 B.n916 585
R1400 B.n916 B.n915 585
R1401 B.n408 B.n407 585
R1402 B.n409 B.n408 585
R1403 B.n908 B.n907 585
R1404 B.n909 B.n908 585
R1405 B.n906 B.n413 585
R1406 B.n417 B.n413 585
R1407 B.n905 B.n904 585
R1408 B.n904 B.n903 585
R1409 B.n415 B.n414 585
R1410 B.n416 B.n415 585
R1411 B.n896 B.n895 585
R1412 B.n897 B.n896 585
R1413 B.n894 B.n422 585
R1414 B.n422 B.n421 585
R1415 B.n893 B.n892 585
R1416 B.n892 B.n891 585
R1417 B.n424 B.n423 585
R1418 B.n425 B.n424 585
R1419 B.n884 B.n883 585
R1420 B.n885 B.n884 585
R1421 B.n882 B.n430 585
R1422 B.n430 B.n429 585
R1423 B.n881 B.n880 585
R1424 B.n880 B.n879 585
R1425 B.n432 B.n431 585
R1426 B.n872 B.n432 585
R1427 B.n871 B.n870 585
R1428 B.n873 B.n871 585
R1429 B.n869 B.n437 585
R1430 B.n437 B.n436 585
R1431 B.n868 B.n867 585
R1432 B.n867 B.n866 585
R1433 B.n439 B.n438 585
R1434 B.n440 B.n439 585
R1435 B.n859 B.n858 585
R1436 B.n860 B.n859 585
R1437 B.n857 B.n445 585
R1438 B.n445 B.n444 585
R1439 B.n856 B.n855 585
R1440 B.n855 B.n854 585
R1441 B.n447 B.n446 585
R1442 B.n448 B.n447 585
R1443 B.n847 B.n846 585
R1444 B.n848 B.n847 585
R1445 B.n845 B.n453 585
R1446 B.n453 B.n452 585
R1447 B.n844 B.n843 585
R1448 B.n843 B.n842 585
R1449 B.n455 B.n454 585
R1450 B.n456 B.n455 585
R1451 B.n835 B.n834 585
R1452 B.n836 B.n835 585
R1453 B.n833 B.n461 585
R1454 B.n461 B.n460 585
R1455 B.n832 B.n831 585
R1456 B.n831 B.n830 585
R1457 B.n463 B.n462 585
R1458 B.n464 B.n463 585
R1459 B.n823 B.n822 585
R1460 B.n824 B.n823 585
R1461 B.n821 B.n469 585
R1462 B.n469 B.n468 585
R1463 B.n820 B.n819 585
R1464 B.n819 B.n818 585
R1465 B.n471 B.n470 585
R1466 B.n472 B.n471 585
R1467 B.n811 B.n810 585
R1468 B.n812 B.n811 585
R1469 B.n809 B.n477 585
R1470 B.n477 B.n476 585
R1471 B.n808 B.n807 585
R1472 B.n807 B.n806 585
R1473 B.n479 B.n478 585
R1474 B.n799 B.n479 585
R1475 B.n798 B.n797 585
R1476 B.n800 B.n798 585
R1477 B.n796 B.n484 585
R1478 B.n484 B.n483 585
R1479 B.n795 B.n794 585
R1480 B.n794 B.n793 585
R1481 B.n486 B.n485 585
R1482 B.n487 B.n486 585
R1483 B.n786 B.n785 585
R1484 B.n787 B.n786 585
R1485 B.n784 B.n492 585
R1486 B.n492 B.n491 585
R1487 B.n783 B.n782 585
R1488 B.n782 B.n781 585
R1489 B.n494 B.n493 585
R1490 B.n495 B.n494 585
R1491 B.n777 B.n776 585
R1492 B.n498 B.n497 585
R1493 B.n773 B.n772 585
R1494 B.n774 B.n773 585
R1495 B.n771 B.n553 585
R1496 B.n770 B.n769 585
R1497 B.n768 B.n767 585
R1498 B.n766 B.n765 585
R1499 B.n764 B.n763 585
R1500 B.n762 B.n761 585
R1501 B.n760 B.n759 585
R1502 B.n758 B.n757 585
R1503 B.n756 B.n755 585
R1504 B.n754 B.n753 585
R1505 B.n752 B.n751 585
R1506 B.n750 B.n749 585
R1507 B.n748 B.n747 585
R1508 B.n746 B.n745 585
R1509 B.n744 B.n743 585
R1510 B.n742 B.n741 585
R1511 B.n740 B.n739 585
R1512 B.n738 B.n737 585
R1513 B.n736 B.n735 585
R1514 B.n734 B.n733 585
R1515 B.n732 B.n731 585
R1516 B.n730 B.n729 585
R1517 B.n728 B.n727 585
R1518 B.n726 B.n725 585
R1519 B.n724 B.n723 585
R1520 B.n722 B.n721 585
R1521 B.n720 B.n719 585
R1522 B.n718 B.n717 585
R1523 B.n716 B.n715 585
R1524 B.n714 B.n713 585
R1525 B.n712 B.n711 585
R1526 B.n710 B.n709 585
R1527 B.n708 B.n707 585
R1528 B.n706 B.n705 585
R1529 B.n704 B.n703 585
R1530 B.n702 B.n701 585
R1531 B.n700 B.n699 585
R1532 B.n698 B.n697 585
R1533 B.n696 B.n695 585
R1534 B.n694 B.n693 585
R1535 B.n692 B.n691 585
R1536 B.n690 B.n689 585
R1537 B.n688 B.n687 585
R1538 B.n686 B.n685 585
R1539 B.n684 B.n683 585
R1540 B.n682 B.n681 585
R1541 B.n680 B.n679 585
R1542 B.n677 B.n676 585
R1543 B.n675 B.n674 585
R1544 B.n673 B.n672 585
R1545 B.n671 B.n670 585
R1546 B.n669 B.n668 585
R1547 B.n667 B.n666 585
R1548 B.n665 B.n664 585
R1549 B.n663 B.n662 585
R1550 B.n661 B.n660 585
R1551 B.n659 B.n658 585
R1552 B.n656 B.n655 585
R1553 B.n654 B.n653 585
R1554 B.n652 B.n651 585
R1555 B.n650 B.n649 585
R1556 B.n648 B.n647 585
R1557 B.n646 B.n645 585
R1558 B.n644 B.n643 585
R1559 B.n642 B.n641 585
R1560 B.n640 B.n639 585
R1561 B.n638 B.n637 585
R1562 B.n636 B.n635 585
R1563 B.n634 B.n633 585
R1564 B.n632 B.n631 585
R1565 B.n630 B.n629 585
R1566 B.n628 B.n627 585
R1567 B.n626 B.n625 585
R1568 B.n624 B.n623 585
R1569 B.n622 B.n621 585
R1570 B.n620 B.n619 585
R1571 B.n618 B.n617 585
R1572 B.n616 B.n615 585
R1573 B.n614 B.n613 585
R1574 B.n612 B.n611 585
R1575 B.n610 B.n609 585
R1576 B.n608 B.n607 585
R1577 B.n606 B.n605 585
R1578 B.n604 B.n603 585
R1579 B.n602 B.n601 585
R1580 B.n600 B.n599 585
R1581 B.n598 B.n597 585
R1582 B.n596 B.n595 585
R1583 B.n594 B.n593 585
R1584 B.n592 B.n591 585
R1585 B.n590 B.n589 585
R1586 B.n588 B.n587 585
R1587 B.n586 B.n585 585
R1588 B.n584 B.n583 585
R1589 B.n582 B.n581 585
R1590 B.n580 B.n579 585
R1591 B.n578 B.n577 585
R1592 B.n576 B.n575 585
R1593 B.n574 B.n573 585
R1594 B.n572 B.n571 585
R1595 B.n570 B.n569 585
R1596 B.n568 B.n567 585
R1597 B.n566 B.n565 585
R1598 B.n564 B.n563 585
R1599 B.n562 B.n561 585
R1600 B.n560 B.n559 585
R1601 B.n558 B.n552 585
R1602 B.n774 B.n552 585
R1603 B.n778 B.n496 585
R1604 B.n496 B.n495 585
R1605 B.n780 B.n779 585
R1606 B.n781 B.n780 585
R1607 B.n490 B.n489 585
R1608 B.n491 B.n490 585
R1609 B.n789 B.n788 585
R1610 B.n788 B.n787 585
R1611 B.n790 B.n488 585
R1612 B.n488 B.n487 585
R1613 B.n792 B.n791 585
R1614 B.n793 B.n792 585
R1615 B.n482 B.n481 585
R1616 B.n483 B.n482 585
R1617 B.n802 B.n801 585
R1618 B.n801 B.n800 585
R1619 B.n803 B.n480 585
R1620 B.n799 B.n480 585
R1621 B.n805 B.n804 585
R1622 B.n806 B.n805 585
R1623 B.n475 B.n474 585
R1624 B.n476 B.n475 585
R1625 B.n814 B.n813 585
R1626 B.n813 B.n812 585
R1627 B.n815 B.n473 585
R1628 B.n473 B.n472 585
R1629 B.n817 B.n816 585
R1630 B.n818 B.n817 585
R1631 B.n467 B.n466 585
R1632 B.n468 B.n467 585
R1633 B.n826 B.n825 585
R1634 B.n825 B.n824 585
R1635 B.n827 B.n465 585
R1636 B.n465 B.n464 585
R1637 B.n829 B.n828 585
R1638 B.n830 B.n829 585
R1639 B.n459 B.n458 585
R1640 B.n460 B.n459 585
R1641 B.n838 B.n837 585
R1642 B.n837 B.n836 585
R1643 B.n839 B.n457 585
R1644 B.n457 B.n456 585
R1645 B.n841 B.n840 585
R1646 B.n842 B.n841 585
R1647 B.n451 B.n450 585
R1648 B.n452 B.n451 585
R1649 B.n850 B.n849 585
R1650 B.n849 B.n848 585
R1651 B.n851 B.n449 585
R1652 B.n449 B.n448 585
R1653 B.n853 B.n852 585
R1654 B.n854 B.n853 585
R1655 B.n443 B.n442 585
R1656 B.n444 B.n443 585
R1657 B.n862 B.n861 585
R1658 B.n861 B.n860 585
R1659 B.n863 B.n441 585
R1660 B.n441 B.n440 585
R1661 B.n865 B.n864 585
R1662 B.n866 B.n865 585
R1663 B.n435 B.n434 585
R1664 B.n436 B.n435 585
R1665 B.n875 B.n874 585
R1666 B.n874 B.n873 585
R1667 B.n876 B.n433 585
R1668 B.n872 B.n433 585
R1669 B.n878 B.n877 585
R1670 B.n879 B.n878 585
R1671 B.n428 B.n427 585
R1672 B.n429 B.n428 585
R1673 B.n887 B.n886 585
R1674 B.n886 B.n885 585
R1675 B.n888 B.n426 585
R1676 B.n426 B.n425 585
R1677 B.n890 B.n889 585
R1678 B.n891 B.n890 585
R1679 B.n420 B.n419 585
R1680 B.n421 B.n420 585
R1681 B.n899 B.n898 585
R1682 B.n898 B.n897 585
R1683 B.n900 B.n418 585
R1684 B.n418 B.n416 585
R1685 B.n902 B.n901 585
R1686 B.n903 B.n902 585
R1687 B.n412 B.n411 585
R1688 B.n417 B.n412 585
R1689 B.n911 B.n910 585
R1690 B.n910 B.n909 585
R1691 B.n912 B.n410 585
R1692 B.n410 B.n409 585
R1693 B.n914 B.n913 585
R1694 B.n915 B.n914 585
R1695 B.n404 B.n403 585
R1696 B.n405 B.n404 585
R1697 B.n923 B.n922 585
R1698 B.n922 B.n921 585
R1699 B.n924 B.n402 585
R1700 B.n402 B.n401 585
R1701 B.n926 B.n925 585
R1702 B.n927 B.n926 585
R1703 B.n396 B.n395 585
R1704 B.n397 B.n396 585
R1705 B.n936 B.n935 585
R1706 B.n935 B.n934 585
R1707 B.n937 B.n394 585
R1708 B.n933 B.n394 585
R1709 B.n939 B.n938 585
R1710 B.n940 B.n939 585
R1711 B.n389 B.n388 585
R1712 B.n390 B.n389 585
R1713 B.n949 B.n948 585
R1714 B.n948 B.n947 585
R1715 B.n950 B.n387 585
R1716 B.n387 B.n386 585
R1717 B.n952 B.n951 585
R1718 B.n953 B.n952 585
R1719 B.n2 B.n0 585
R1720 B.n4 B.n2 585
R1721 B.n3 B.n1 585
R1722 B.n1154 B.n3 585
R1723 B.n1152 B.n1151 585
R1724 B.n1153 B.n1152 585
R1725 B.n1150 B.n9 585
R1726 B.n9 B.n8 585
R1727 B.n1149 B.n1148 585
R1728 B.n1148 B.n1147 585
R1729 B.n11 B.n10 585
R1730 B.n1146 B.n11 585
R1731 B.n1144 B.n1143 585
R1732 B.n1145 B.n1144 585
R1733 B.n1142 B.n15 585
R1734 B.n18 B.n15 585
R1735 B.n1141 B.n1140 585
R1736 B.n1140 B.n1139 585
R1737 B.n17 B.n16 585
R1738 B.n1138 B.n17 585
R1739 B.n1136 B.n1135 585
R1740 B.n1137 B.n1136 585
R1741 B.n1134 B.n23 585
R1742 B.n23 B.n22 585
R1743 B.n1133 B.n1132 585
R1744 B.n1132 B.n1131 585
R1745 B.n25 B.n24 585
R1746 B.n1130 B.n25 585
R1747 B.n1128 B.n1127 585
R1748 B.n1129 B.n1128 585
R1749 B.n1126 B.n30 585
R1750 B.n30 B.n29 585
R1751 B.n1125 B.n1124 585
R1752 B.n1124 B.n1123 585
R1753 B.n32 B.n31 585
R1754 B.n1122 B.n32 585
R1755 B.n1120 B.n1119 585
R1756 B.n1121 B.n1120 585
R1757 B.n1118 B.n37 585
R1758 B.n37 B.n36 585
R1759 B.n1117 B.n1116 585
R1760 B.n1116 B.n1115 585
R1761 B.n39 B.n38 585
R1762 B.n1114 B.n39 585
R1763 B.n1112 B.n1111 585
R1764 B.n1113 B.n1112 585
R1765 B.n1110 B.n44 585
R1766 B.n44 B.n43 585
R1767 B.n1109 B.n1108 585
R1768 B.n1108 B.n1107 585
R1769 B.n46 B.n45 585
R1770 B.n1106 B.n46 585
R1771 B.n1104 B.n1103 585
R1772 B.n1105 B.n1104 585
R1773 B.n1102 B.n50 585
R1774 B.n53 B.n50 585
R1775 B.n1101 B.n1100 585
R1776 B.n1100 B.n1099 585
R1777 B.n52 B.n51 585
R1778 B.n1098 B.n52 585
R1779 B.n1096 B.n1095 585
R1780 B.n1097 B.n1096 585
R1781 B.n1094 B.n58 585
R1782 B.n58 B.n57 585
R1783 B.n1093 B.n1092 585
R1784 B.n1092 B.n1091 585
R1785 B.n60 B.n59 585
R1786 B.n1090 B.n60 585
R1787 B.n1088 B.n1087 585
R1788 B.n1089 B.n1088 585
R1789 B.n1086 B.n65 585
R1790 B.n65 B.n64 585
R1791 B.n1085 B.n1084 585
R1792 B.n1084 B.n1083 585
R1793 B.n67 B.n66 585
R1794 B.n1082 B.n67 585
R1795 B.n1080 B.n1079 585
R1796 B.n1081 B.n1080 585
R1797 B.n1078 B.n72 585
R1798 B.n72 B.n71 585
R1799 B.n1077 B.n1076 585
R1800 B.n1076 B.n1075 585
R1801 B.n74 B.n73 585
R1802 B.n1074 B.n74 585
R1803 B.n1072 B.n1071 585
R1804 B.n1073 B.n1072 585
R1805 B.n1070 B.n79 585
R1806 B.n79 B.n78 585
R1807 B.n1069 B.n1068 585
R1808 B.n1068 B.n1067 585
R1809 B.n81 B.n80 585
R1810 B.n1066 B.n81 585
R1811 B.n1064 B.n1063 585
R1812 B.n1065 B.n1064 585
R1813 B.n1062 B.n86 585
R1814 B.n86 B.n85 585
R1815 B.n1061 B.n1060 585
R1816 B.n1060 B.n1059 585
R1817 B.n88 B.n87 585
R1818 B.n1058 B.n88 585
R1819 B.n1056 B.n1055 585
R1820 B.n1057 B.n1056 585
R1821 B.n1054 B.n92 585
R1822 B.n95 B.n92 585
R1823 B.n1053 B.n1052 585
R1824 B.n1052 B.n1051 585
R1825 B.n94 B.n93 585
R1826 B.n1050 B.n94 585
R1827 B.n1048 B.n1047 585
R1828 B.n1049 B.n1048 585
R1829 B.n1046 B.n100 585
R1830 B.n100 B.n99 585
R1831 B.n1045 B.n1044 585
R1832 B.n1044 B.n1043 585
R1833 B.n102 B.n101 585
R1834 B.n1042 B.n102 585
R1835 B.n1040 B.n1039 585
R1836 B.n1041 B.n1040 585
R1837 B.n1038 B.n107 585
R1838 B.n107 B.n106 585
R1839 B.n1157 B.n1156 585
R1840 B.n1156 B.n1155 585
R1841 B.n776 B.n496 478.086
R1842 B.n1036 B.n107 478.086
R1843 B.n552 B.n494 478.086
R1844 B.n1032 B.n164 478.086
R1845 B.n556 B.t11 399.839
R1846 B.n165 B.t20 399.839
R1847 B.n554 B.t18 399.839
R1848 B.n168 B.t14 399.839
R1849 B.n557 B.t10 332.93
R1850 B.n166 B.t21 332.93
R1851 B.n555 B.t17 332.93
R1852 B.n169 B.t15 332.93
R1853 B.n556 B.t8 324.041
R1854 B.n554 B.t16 324.041
R1855 B.n168 B.t12 324.041
R1856 B.n165 B.t19 324.041
R1857 B.n1034 B.n1033 256.663
R1858 B.n1034 B.n162 256.663
R1859 B.n1034 B.n161 256.663
R1860 B.n1034 B.n160 256.663
R1861 B.n1034 B.n159 256.663
R1862 B.n1034 B.n158 256.663
R1863 B.n1034 B.n157 256.663
R1864 B.n1034 B.n156 256.663
R1865 B.n1034 B.n155 256.663
R1866 B.n1034 B.n154 256.663
R1867 B.n1034 B.n153 256.663
R1868 B.n1034 B.n152 256.663
R1869 B.n1034 B.n151 256.663
R1870 B.n1034 B.n150 256.663
R1871 B.n1034 B.n149 256.663
R1872 B.n1034 B.n148 256.663
R1873 B.n1034 B.n147 256.663
R1874 B.n1034 B.n146 256.663
R1875 B.n1034 B.n145 256.663
R1876 B.n1034 B.n144 256.663
R1877 B.n1034 B.n143 256.663
R1878 B.n1034 B.n142 256.663
R1879 B.n1034 B.n141 256.663
R1880 B.n1034 B.n140 256.663
R1881 B.n1034 B.n139 256.663
R1882 B.n1034 B.n138 256.663
R1883 B.n1034 B.n137 256.663
R1884 B.n1034 B.n136 256.663
R1885 B.n1034 B.n135 256.663
R1886 B.n1034 B.n134 256.663
R1887 B.n1034 B.n133 256.663
R1888 B.n1034 B.n132 256.663
R1889 B.n1034 B.n131 256.663
R1890 B.n1034 B.n130 256.663
R1891 B.n1034 B.n129 256.663
R1892 B.n1034 B.n128 256.663
R1893 B.n1034 B.n127 256.663
R1894 B.n1034 B.n126 256.663
R1895 B.n1034 B.n125 256.663
R1896 B.n1034 B.n124 256.663
R1897 B.n1034 B.n123 256.663
R1898 B.n1034 B.n122 256.663
R1899 B.n1034 B.n121 256.663
R1900 B.n1034 B.n120 256.663
R1901 B.n1034 B.n119 256.663
R1902 B.n1034 B.n118 256.663
R1903 B.n1034 B.n117 256.663
R1904 B.n1034 B.n116 256.663
R1905 B.n1034 B.n115 256.663
R1906 B.n1034 B.n114 256.663
R1907 B.n1034 B.n113 256.663
R1908 B.n1034 B.n112 256.663
R1909 B.n1034 B.n111 256.663
R1910 B.n1034 B.n110 256.663
R1911 B.n1035 B.n1034 256.663
R1912 B.n775 B.n774 256.663
R1913 B.n774 B.n499 256.663
R1914 B.n774 B.n500 256.663
R1915 B.n774 B.n501 256.663
R1916 B.n774 B.n502 256.663
R1917 B.n774 B.n503 256.663
R1918 B.n774 B.n504 256.663
R1919 B.n774 B.n505 256.663
R1920 B.n774 B.n506 256.663
R1921 B.n774 B.n507 256.663
R1922 B.n774 B.n508 256.663
R1923 B.n774 B.n509 256.663
R1924 B.n774 B.n510 256.663
R1925 B.n774 B.n511 256.663
R1926 B.n774 B.n512 256.663
R1927 B.n774 B.n513 256.663
R1928 B.n774 B.n514 256.663
R1929 B.n774 B.n515 256.663
R1930 B.n774 B.n516 256.663
R1931 B.n774 B.n517 256.663
R1932 B.n774 B.n518 256.663
R1933 B.n774 B.n519 256.663
R1934 B.n774 B.n520 256.663
R1935 B.n774 B.n521 256.663
R1936 B.n774 B.n522 256.663
R1937 B.n774 B.n523 256.663
R1938 B.n774 B.n524 256.663
R1939 B.n774 B.n525 256.663
R1940 B.n774 B.n526 256.663
R1941 B.n774 B.n527 256.663
R1942 B.n774 B.n528 256.663
R1943 B.n774 B.n529 256.663
R1944 B.n774 B.n530 256.663
R1945 B.n774 B.n531 256.663
R1946 B.n774 B.n532 256.663
R1947 B.n774 B.n533 256.663
R1948 B.n774 B.n534 256.663
R1949 B.n774 B.n535 256.663
R1950 B.n774 B.n536 256.663
R1951 B.n774 B.n537 256.663
R1952 B.n774 B.n538 256.663
R1953 B.n774 B.n539 256.663
R1954 B.n774 B.n540 256.663
R1955 B.n774 B.n541 256.663
R1956 B.n774 B.n542 256.663
R1957 B.n774 B.n543 256.663
R1958 B.n774 B.n544 256.663
R1959 B.n774 B.n545 256.663
R1960 B.n774 B.n546 256.663
R1961 B.n774 B.n547 256.663
R1962 B.n774 B.n548 256.663
R1963 B.n774 B.n549 256.663
R1964 B.n774 B.n550 256.663
R1965 B.n774 B.n551 256.663
R1966 B.n780 B.n496 163.367
R1967 B.n780 B.n490 163.367
R1968 B.n788 B.n490 163.367
R1969 B.n788 B.n488 163.367
R1970 B.n792 B.n488 163.367
R1971 B.n792 B.n482 163.367
R1972 B.n801 B.n482 163.367
R1973 B.n801 B.n480 163.367
R1974 B.n805 B.n480 163.367
R1975 B.n805 B.n475 163.367
R1976 B.n813 B.n475 163.367
R1977 B.n813 B.n473 163.367
R1978 B.n817 B.n473 163.367
R1979 B.n817 B.n467 163.367
R1980 B.n825 B.n467 163.367
R1981 B.n825 B.n465 163.367
R1982 B.n829 B.n465 163.367
R1983 B.n829 B.n459 163.367
R1984 B.n837 B.n459 163.367
R1985 B.n837 B.n457 163.367
R1986 B.n841 B.n457 163.367
R1987 B.n841 B.n451 163.367
R1988 B.n849 B.n451 163.367
R1989 B.n849 B.n449 163.367
R1990 B.n853 B.n449 163.367
R1991 B.n853 B.n443 163.367
R1992 B.n861 B.n443 163.367
R1993 B.n861 B.n441 163.367
R1994 B.n865 B.n441 163.367
R1995 B.n865 B.n435 163.367
R1996 B.n874 B.n435 163.367
R1997 B.n874 B.n433 163.367
R1998 B.n878 B.n433 163.367
R1999 B.n878 B.n428 163.367
R2000 B.n886 B.n428 163.367
R2001 B.n886 B.n426 163.367
R2002 B.n890 B.n426 163.367
R2003 B.n890 B.n420 163.367
R2004 B.n898 B.n420 163.367
R2005 B.n898 B.n418 163.367
R2006 B.n902 B.n418 163.367
R2007 B.n902 B.n412 163.367
R2008 B.n910 B.n412 163.367
R2009 B.n910 B.n410 163.367
R2010 B.n914 B.n410 163.367
R2011 B.n914 B.n404 163.367
R2012 B.n922 B.n404 163.367
R2013 B.n922 B.n402 163.367
R2014 B.n926 B.n402 163.367
R2015 B.n926 B.n396 163.367
R2016 B.n935 B.n396 163.367
R2017 B.n935 B.n394 163.367
R2018 B.n939 B.n394 163.367
R2019 B.n939 B.n389 163.367
R2020 B.n948 B.n389 163.367
R2021 B.n948 B.n387 163.367
R2022 B.n952 B.n387 163.367
R2023 B.n952 B.n2 163.367
R2024 B.n1156 B.n2 163.367
R2025 B.n1156 B.n3 163.367
R2026 B.n1152 B.n3 163.367
R2027 B.n1152 B.n9 163.367
R2028 B.n1148 B.n9 163.367
R2029 B.n1148 B.n11 163.367
R2030 B.n1144 B.n11 163.367
R2031 B.n1144 B.n15 163.367
R2032 B.n1140 B.n15 163.367
R2033 B.n1140 B.n17 163.367
R2034 B.n1136 B.n17 163.367
R2035 B.n1136 B.n23 163.367
R2036 B.n1132 B.n23 163.367
R2037 B.n1132 B.n25 163.367
R2038 B.n1128 B.n25 163.367
R2039 B.n1128 B.n30 163.367
R2040 B.n1124 B.n30 163.367
R2041 B.n1124 B.n32 163.367
R2042 B.n1120 B.n32 163.367
R2043 B.n1120 B.n37 163.367
R2044 B.n1116 B.n37 163.367
R2045 B.n1116 B.n39 163.367
R2046 B.n1112 B.n39 163.367
R2047 B.n1112 B.n44 163.367
R2048 B.n1108 B.n44 163.367
R2049 B.n1108 B.n46 163.367
R2050 B.n1104 B.n46 163.367
R2051 B.n1104 B.n50 163.367
R2052 B.n1100 B.n50 163.367
R2053 B.n1100 B.n52 163.367
R2054 B.n1096 B.n52 163.367
R2055 B.n1096 B.n58 163.367
R2056 B.n1092 B.n58 163.367
R2057 B.n1092 B.n60 163.367
R2058 B.n1088 B.n60 163.367
R2059 B.n1088 B.n65 163.367
R2060 B.n1084 B.n65 163.367
R2061 B.n1084 B.n67 163.367
R2062 B.n1080 B.n67 163.367
R2063 B.n1080 B.n72 163.367
R2064 B.n1076 B.n72 163.367
R2065 B.n1076 B.n74 163.367
R2066 B.n1072 B.n74 163.367
R2067 B.n1072 B.n79 163.367
R2068 B.n1068 B.n79 163.367
R2069 B.n1068 B.n81 163.367
R2070 B.n1064 B.n81 163.367
R2071 B.n1064 B.n86 163.367
R2072 B.n1060 B.n86 163.367
R2073 B.n1060 B.n88 163.367
R2074 B.n1056 B.n88 163.367
R2075 B.n1056 B.n92 163.367
R2076 B.n1052 B.n92 163.367
R2077 B.n1052 B.n94 163.367
R2078 B.n1048 B.n94 163.367
R2079 B.n1048 B.n100 163.367
R2080 B.n1044 B.n100 163.367
R2081 B.n1044 B.n102 163.367
R2082 B.n1040 B.n102 163.367
R2083 B.n1040 B.n107 163.367
R2084 B.n773 B.n498 163.367
R2085 B.n773 B.n553 163.367
R2086 B.n769 B.n768 163.367
R2087 B.n765 B.n764 163.367
R2088 B.n761 B.n760 163.367
R2089 B.n757 B.n756 163.367
R2090 B.n753 B.n752 163.367
R2091 B.n749 B.n748 163.367
R2092 B.n745 B.n744 163.367
R2093 B.n741 B.n740 163.367
R2094 B.n737 B.n736 163.367
R2095 B.n733 B.n732 163.367
R2096 B.n729 B.n728 163.367
R2097 B.n725 B.n724 163.367
R2098 B.n721 B.n720 163.367
R2099 B.n717 B.n716 163.367
R2100 B.n713 B.n712 163.367
R2101 B.n709 B.n708 163.367
R2102 B.n705 B.n704 163.367
R2103 B.n701 B.n700 163.367
R2104 B.n697 B.n696 163.367
R2105 B.n693 B.n692 163.367
R2106 B.n689 B.n688 163.367
R2107 B.n685 B.n684 163.367
R2108 B.n681 B.n680 163.367
R2109 B.n676 B.n675 163.367
R2110 B.n672 B.n671 163.367
R2111 B.n668 B.n667 163.367
R2112 B.n664 B.n663 163.367
R2113 B.n660 B.n659 163.367
R2114 B.n655 B.n654 163.367
R2115 B.n651 B.n650 163.367
R2116 B.n647 B.n646 163.367
R2117 B.n643 B.n642 163.367
R2118 B.n639 B.n638 163.367
R2119 B.n635 B.n634 163.367
R2120 B.n631 B.n630 163.367
R2121 B.n627 B.n626 163.367
R2122 B.n623 B.n622 163.367
R2123 B.n619 B.n618 163.367
R2124 B.n615 B.n614 163.367
R2125 B.n611 B.n610 163.367
R2126 B.n607 B.n606 163.367
R2127 B.n603 B.n602 163.367
R2128 B.n599 B.n598 163.367
R2129 B.n595 B.n594 163.367
R2130 B.n591 B.n590 163.367
R2131 B.n587 B.n586 163.367
R2132 B.n583 B.n582 163.367
R2133 B.n579 B.n578 163.367
R2134 B.n575 B.n574 163.367
R2135 B.n571 B.n570 163.367
R2136 B.n567 B.n566 163.367
R2137 B.n563 B.n562 163.367
R2138 B.n559 B.n552 163.367
R2139 B.n782 B.n494 163.367
R2140 B.n782 B.n492 163.367
R2141 B.n786 B.n492 163.367
R2142 B.n786 B.n486 163.367
R2143 B.n794 B.n486 163.367
R2144 B.n794 B.n484 163.367
R2145 B.n798 B.n484 163.367
R2146 B.n798 B.n479 163.367
R2147 B.n807 B.n479 163.367
R2148 B.n807 B.n477 163.367
R2149 B.n811 B.n477 163.367
R2150 B.n811 B.n471 163.367
R2151 B.n819 B.n471 163.367
R2152 B.n819 B.n469 163.367
R2153 B.n823 B.n469 163.367
R2154 B.n823 B.n463 163.367
R2155 B.n831 B.n463 163.367
R2156 B.n831 B.n461 163.367
R2157 B.n835 B.n461 163.367
R2158 B.n835 B.n455 163.367
R2159 B.n843 B.n455 163.367
R2160 B.n843 B.n453 163.367
R2161 B.n847 B.n453 163.367
R2162 B.n847 B.n447 163.367
R2163 B.n855 B.n447 163.367
R2164 B.n855 B.n445 163.367
R2165 B.n859 B.n445 163.367
R2166 B.n859 B.n439 163.367
R2167 B.n867 B.n439 163.367
R2168 B.n867 B.n437 163.367
R2169 B.n871 B.n437 163.367
R2170 B.n871 B.n432 163.367
R2171 B.n880 B.n432 163.367
R2172 B.n880 B.n430 163.367
R2173 B.n884 B.n430 163.367
R2174 B.n884 B.n424 163.367
R2175 B.n892 B.n424 163.367
R2176 B.n892 B.n422 163.367
R2177 B.n896 B.n422 163.367
R2178 B.n896 B.n415 163.367
R2179 B.n904 B.n415 163.367
R2180 B.n904 B.n413 163.367
R2181 B.n908 B.n413 163.367
R2182 B.n908 B.n408 163.367
R2183 B.n916 B.n408 163.367
R2184 B.n916 B.n406 163.367
R2185 B.n920 B.n406 163.367
R2186 B.n920 B.n400 163.367
R2187 B.n928 B.n400 163.367
R2188 B.n928 B.n398 163.367
R2189 B.n932 B.n398 163.367
R2190 B.n932 B.n393 163.367
R2191 B.n941 B.n393 163.367
R2192 B.n941 B.n391 163.367
R2193 B.n946 B.n391 163.367
R2194 B.n946 B.n385 163.367
R2195 B.n954 B.n385 163.367
R2196 B.n955 B.n954 163.367
R2197 B.n955 B.n5 163.367
R2198 B.n6 B.n5 163.367
R2199 B.n7 B.n6 163.367
R2200 B.n960 B.n7 163.367
R2201 B.n960 B.n12 163.367
R2202 B.n13 B.n12 163.367
R2203 B.n14 B.n13 163.367
R2204 B.n965 B.n14 163.367
R2205 B.n965 B.n19 163.367
R2206 B.n20 B.n19 163.367
R2207 B.n21 B.n20 163.367
R2208 B.n970 B.n21 163.367
R2209 B.n970 B.n26 163.367
R2210 B.n27 B.n26 163.367
R2211 B.n28 B.n27 163.367
R2212 B.n975 B.n28 163.367
R2213 B.n975 B.n33 163.367
R2214 B.n34 B.n33 163.367
R2215 B.n35 B.n34 163.367
R2216 B.n980 B.n35 163.367
R2217 B.n980 B.n40 163.367
R2218 B.n41 B.n40 163.367
R2219 B.n42 B.n41 163.367
R2220 B.n985 B.n42 163.367
R2221 B.n985 B.n47 163.367
R2222 B.n48 B.n47 163.367
R2223 B.n49 B.n48 163.367
R2224 B.n990 B.n49 163.367
R2225 B.n990 B.n54 163.367
R2226 B.n55 B.n54 163.367
R2227 B.n56 B.n55 163.367
R2228 B.n995 B.n56 163.367
R2229 B.n995 B.n61 163.367
R2230 B.n62 B.n61 163.367
R2231 B.n63 B.n62 163.367
R2232 B.n1000 B.n63 163.367
R2233 B.n1000 B.n68 163.367
R2234 B.n69 B.n68 163.367
R2235 B.n70 B.n69 163.367
R2236 B.n1005 B.n70 163.367
R2237 B.n1005 B.n75 163.367
R2238 B.n76 B.n75 163.367
R2239 B.n77 B.n76 163.367
R2240 B.n1010 B.n77 163.367
R2241 B.n1010 B.n82 163.367
R2242 B.n83 B.n82 163.367
R2243 B.n84 B.n83 163.367
R2244 B.n1015 B.n84 163.367
R2245 B.n1015 B.n89 163.367
R2246 B.n90 B.n89 163.367
R2247 B.n91 B.n90 163.367
R2248 B.n1020 B.n91 163.367
R2249 B.n1020 B.n96 163.367
R2250 B.n97 B.n96 163.367
R2251 B.n98 B.n97 163.367
R2252 B.n1025 B.n98 163.367
R2253 B.n1025 B.n103 163.367
R2254 B.n104 B.n103 163.367
R2255 B.n105 B.n104 163.367
R2256 B.n164 B.n105 163.367
R2257 B.n171 B.n109 163.367
R2258 B.n175 B.n174 163.367
R2259 B.n179 B.n178 163.367
R2260 B.n183 B.n182 163.367
R2261 B.n187 B.n186 163.367
R2262 B.n191 B.n190 163.367
R2263 B.n195 B.n194 163.367
R2264 B.n199 B.n198 163.367
R2265 B.n203 B.n202 163.367
R2266 B.n207 B.n206 163.367
R2267 B.n211 B.n210 163.367
R2268 B.n215 B.n214 163.367
R2269 B.n219 B.n218 163.367
R2270 B.n223 B.n222 163.367
R2271 B.n227 B.n226 163.367
R2272 B.n231 B.n230 163.367
R2273 B.n235 B.n234 163.367
R2274 B.n239 B.n238 163.367
R2275 B.n243 B.n242 163.367
R2276 B.n247 B.n246 163.367
R2277 B.n251 B.n250 163.367
R2278 B.n255 B.n254 163.367
R2279 B.n259 B.n258 163.367
R2280 B.n263 B.n262 163.367
R2281 B.n267 B.n266 163.367
R2282 B.n271 B.n270 163.367
R2283 B.n275 B.n274 163.367
R2284 B.n279 B.n278 163.367
R2285 B.n283 B.n282 163.367
R2286 B.n287 B.n286 163.367
R2287 B.n291 B.n290 163.367
R2288 B.n295 B.n294 163.367
R2289 B.n299 B.n298 163.367
R2290 B.n303 B.n302 163.367
R2291 B.n307 B.n306 163.367
R2292 B.n311 B.n310 163.367
R2293 B.n315 B.n314 163.367
R2294 B.n319 B.n318 163.367
R2295 B.n323 B.n322 163.367
R2296 B.n327 B.n326 163.367
R2297 B.n331 B.n330 163.367
R2298 B.n335 B.n334 163.367
R2299 B.n339 B.n338 163.367
R2300 B.n343 B.n342 163.367
R2301 B.n347 B.n346 163.367
R2302 B.n351 B.n350 163.367
R2303 B.n355 B.n354 163.367
R2304 B.n359 B.n358 163.367
R2305 B.n363 B.n362 163.367
R2306 B.n367 B.n366 163.367
R2307 B.n371 B.n370 163.367
R2308 B.n375 B.n374 163.367
R2309 B.n379 B.n378 163.367
R2310 B.n381 B.n163 163.367
R2311 B.n776 B.n775 71.676
R2312 B.n553 B.n499 71.676
R2313 B.n768 B.n500 71.676
R2314 B.n764 B.n501 71.676
R2315 B.n760 B.n502 71.676
R2316 B.n756 B.n503 71.676
R2317 B.n752 B.n504 71.676
R2318 B.n748 B.n505 71.676
R2319 B.n744 B.n506 71.676
R2320 B.n740 B.n507 71.676
R2321 B.n736 B.n508 71.676
R2322 B.n732 B.n509 71.676
R2323 B.n728 B.n510 71.676
R2324 B.n724 B.n511 71.676
R2325 B.n720 B.n512 71.676
R2326 B.n716 B.n513 71.676
R2327 B.n712 B.n514 71.676
R2328 B.n708 B.n515 71.676
R2329 B.n704 B.n516 71.676
R2330 B.n700 B.n517 71.676
R2331 B.n696 B.n518 71.676
R2332 B.n692 B.n519 71.676
R2333 B.n688 B.n520 71.676
R2334 B.n684 B.n521 71.676
R2335 B.n680 B.n522 71.676
R2336 B.n675 B.n523 71.676
R2337 B.n671 B.n524 71.676
R2338 B.n667 B.n525 71.676
R2339 B.n663 B.n526 71.676
R2340 B.n659 B.n527 71.676
R2341 B.n654 B.n528 71.676
R2342 B.n650 B.n529 71.676
R2343 B.n646 B.n530 71.676
R2344 B.n642 B.n531 71.676
R2345 B.n638 B.n532 71.676
R2346 B.n634 B.n533 71.676
R2347 B.n630 B.n534 71.676
R2348 B.n626 B.n535 71.676
R2349 B.n622 B.n536 71.676
R2350 B.n618 B.n537 71.676
R2351 B.n614 B.n538 71.676
R2352 B.n610 B.n539 71.676
R2353 B.n606 B.n540 71.676
R2354 B.n602 B.n541 71.676
R2355 B.n598 B.n542 71.676
R2356 B.n594 B.n543 71.676
R2357 B.n590 B.n544 71.676
R2358 B.n586 B.n545 71.676
R2359 B.n582 B.n546 71.676
R2360 B.n578 B.n547 71.676
R2361 B.n574 B.n548 71.676
R2362 B.n570 B.n549 71.676
R2363 B.n566 B.n550 71.676
R2364 B.n562 B.n551 71.676
R2365 B.n1036 B.n1035 71.676
R2366 B.n171 B.n110 71.676
R2367 B.n175 B.n111 71.676
R2368 B.n179 B.n112 71.676
R2369 B.n183 B.n113 71.676
R2370 B.n187 B.n114 71.676
R2371 B.n191 B.n115 71.676
R2372 B.n195 B.n116 71.676
R2373 B.n199 B.n117 71.676
R2374 B.n203 B.n118 71.676
R2375 B.n207 B.n119 71.676
R2376 B.n211 B.n120 71.676
R2377 B.n215 B.n121 71.676
R2378 B.n219 B.n122 71.676
R2379 B.n223 B.n123 71.676
R2380 B.n227 B.n124 71.676
R2381 B.n231 B.n125 71.676
R2382 B.n235 B.n126 71.676
R2383 B.n239 B.n127 71.676
R2384 B.n243 B.n128 71.676
R2385 B.n247 B.n129 71.676
R2386 B.n251 B.n130 71.676
R2387 B.n255 B.n131 71.676
R2388 B.n259 B.n132 71.676
R2389 B.n263 B.n133 71.676
R2390 B.n267 B.n134 71.676
R2391 B.n271 B.n135 71.676
R2392 B.n275 B.n136 71.676
R2393 B.n279 B.n137 71.676
R2394 B.n283 B.n138 71.676
R2395 B.n287 B.n139 71.676
R2396 B.n291 B.n140 71.676
R2397 B.n295 B.n141 71.676
R2398 B.n299 B.n142 71.676
R2399 B.n303 B.n143 71.676
R2400 B.n307 B.n144 71.676
R2401 B.n311 B.n145 71.676
R2402 B.n315 B.n146 71.676
R2403 B.n319 B.n147 71.676
R2404 B.n323 B.n148 71.676
R2405 B.n327 B.n149 71.676
R2406 B.n331 B.n150 71.676
R2407 B.n335 B.n151 71.676
R2408 B.n339 B.n152 71.676
R2409 B.n343 B.n153 71.676
R2410 B.n347 B.n154 71.676
R2411 B.n351 B.n155 71.676
R2412 B.n355 B.n156 71.676
R2413 B.n359 B.n157 71.676
R2414 B.n363 B.n158 71.676
R2415 B.n367 B.n159 71.676
R2416 B.n371 B.n160 71.676
R2417 B.n375 B.n161 71.676
R2418 B.n379 B.n162 71.676
R2419 B.n1033 B.n163 71.676
R2420 B.n1033 B.n1032 71.676
R2421 B.n381 B.n162 71.676
R2422 B.n378 B.n161 71.676
R2423 B.n374 B.n160 71.676
R2424 B.n370 B.n159 71.676
R2425 B.n366 B.n158 71.676
R2426 B.n362 B.n157 71.676
R2427 B.n358 B.n156 71.676
R2428 B.n354 B.n155 71.676
R2429 B.n350 B.n154 71.676
R2430 B.n346 B.n153 71.676
R2431 B.n342 B.n152 71.676
R2432 B.n338 B.n151 71.676
R2433 B.n334 B.n150 71.676
R2434 B.n330 B.n149 71.676
R2435 B.n326 B.n148 71.676
R2436 B.n322 B.n147 71.676
R2437 B.n318 B.n146 71.676
R2438 B.n314 B.n145 71.676
R2439 B.n310 B.n144 71.676
R2440 B.n306 B.n143 71.676
R2441 B.n302 B.n142 71.676
R2442 B.n298 B.n141 71.676
R2443 B.n294 B.n140 71.676
R2444 B.n290 B.n139 71.676
R2445 B.n286 B.n138 71.676
R2446 B.n282 B.n137 71.676
R2447 B.n278 B.n136 71.676
R2448 B.n274 B.n135 71.676
R2449 B.n270 B.n134 71.676
R2450 B.n266 B.n133 71.676
R2451 B.n262 B.n132 71.676
R2452 B.n258 B.n131 71.676
R2453 B.n254 B.n130 71.676
R2454 B.n250 B.n129 71.676
R2455 B.n246 B.n128 71.676
R2456 B.n242 B.n127 71.676
R2457 B.n238 B.n126 71.676
R2458 B.n234 B.n125 71.676
R2459 B.n230 B.n124 71.676
R2460 B.n226 B.n123 71.676
R2461 B.n222 B.n122 71.676
R2462 B.n218 B.n121 71.676
R2463 B.n214 B.n120 71.676
R2464 B.n210 B.n119 71.676
R2465 B.n206 B.n118 71.676
R2466 B.n202 B.n117 71.676
R2467 B.n198 B.n116 71.676
R2468 B.n194 B.n115 71.676
R2469 B.n190 B.n114 71.676
R2470 B.n186 B.n113 71.676
R2471 B.n182 B.n112 71.676
R2472 B.n178 B.n111 71.676
R2473 B.n174 B.n110 71.676
R2474 B.n1035 B.n109 71.676
R2475 B.n775 B.n498 71.676
R2476 B.n769 B.n499 71.676
R2477 B.n765 B.n500 71.676
R2478 B.n761 B.n501 71.676
R2479 B.n757 B.n502 71.676
R2480 B.n753 B.n503 71.676
R2481 B.n749 B.n504 71.676
R2482 B.n745 B.n505 71.676
R2483 B.n741 B.n506 71.676
R2484 B.n737 B.n507 71.676
R2485 B.n733 B.n508 71.676
R2486 B.n729 B.n509 71.676
R2487 B.n725 B.n510 71.676
R2488 B.n721 B.n511 71.676
R2489 B.n717 B.n512 71.676
R2490 B.n713 B.n513 71.676
R2491 B.n709 B.n514 71.676
R2492 B.n705 B.n515 71.676
R2493 B.n701 B.n516 71.676
R2494 B.n697 B.n517 71.676
R2495 B.n693 B.n518 71.676
R2496 B.n689 B.n519 71.676
R2497 B.n685 B.n520 71.676
R2498 B.n681 B.n521 71.676
R2499 B.n676 B.n522 71.676
R2500 B.n672 B.n523 71.676
R2501 B.n668 B.n524 71.676
R2502 B.n664 B.n525 71.676
R2503 B.n660 B.n526 71.676
R2504 B.n655 B.n527 71.676
R2505 B.n651 B.n528 71.676
R2506 B.n647 B.n529 71.676
R2507 B.n643 B.n530 71.676
R2508 B.n639 B.n531 71.676
R2509 B.n635 B.n532 71.676
R2510 B.n631 B.n533 71.676
R2511 B.n627 B.n534 71.676
R2512 B.n623 B.n535 71.676
R2513 B.n619 B.n536 71.676
R2514 B.n615 B.n537 71.676
R2515 B.n611 B.n538 71.676
R2516 B.n607 B.n539 71.676
R2517 B.n603 B.n540 71.676
R2518 B.n599 B.n541 71.676
R2519 B.n595 B.n542 71.676
R2520 B.n591 B.n543 71.676
R2521 B.n587 B.n544 71.676
R2522 B.n583 B.n545 71.676
R2523 B.n579 B.n546 71.676
R2524 B.n575 B.n547 71.676
R2525 B.n571 B.n548 71.676
R2526 B.n567 B.n549 71.676
R2527 B.n563 B.n550 71.676
R2528 B.n559 B.n551 71.676
R2529 B.n557 B.n556 66.9096
R2530 B.n555 B.n554 66.9096
R2531 B.n169 B.n168 66.9096
R2532 B.n166 B.n165 66.9096
R2533 B.n774 B.n495 61.5199
R2534 B.n1034 B.n106 61.5199
R2535 B.n657 B.n557 59.5399
R2536 B.n678 B.n555 59.5399
R2537 B.n170 B.n169 59.5399
R2538 B.n167 B.n166 59.5399
R2539 B.n781 B.n495 37.021
R2540 B.n781 B.n491 37.021
R2541 B.n787 B.n491 37.021
R2542 B.n787 B.n487 37.021
R2543 B.n793 B.n487 37.021
R2544 B.n793 B.n483 37.021
R2545 B.n800 B.n483 37.021
R2546 B.n800 B.n799 37.021
R2547 B.n806 B.n476 37.021
R2548 B.n812 B.n476 37.021
R2549 B.n812 B.n472 37.021
R2550 B.n818 B.n472 37.021
R2551 B.n818 B.n468 37.021
R2552 B.n824 B.n468 37.021
R2553 B.n824 B.n464 37.021
R2554 B.n830 B.n464 37.021
R2555 B.n830 B.n460 37.021
R2556 B.n836 B.n460 37.021
R2557 B.n836 B.n456 37.021
R2558 B.n842 B.n456 37.021
R2559 B.n848 B.n452 37.021
R2560 B.n848 B.n448 37.021
R2561 B.n854 B.n448 37.021
R2562 B.n854 B.n444 37.021
R2563 B.n860 B.n444 37.021
R2564 B.n860 B.n440 37.021
R2565 B.n866 B.n440 37.021
R2566 B.n866 B.n436 37.021
R2567 B.n873 B.n436 37.021
R2568 B.n873 B.n872 37.021
R2569 B.n879 B.n429 37.021
R2570 B.n885 B.n429 37.021
R2571 B.n885 B.n425 37.021
R2572 B.n891 B.n425 37.021
R2573 B.n891 B.n421 37.021
R2574 B.n897 B.n421 37.021
R2575 B.n897 B.n416 37.021
R2576 B.n903 B.n416 37.021
R2577 B.n903 B.n417 37.021
R2578 B.n909 B.n409 37.021
R2579 B.n915 B.n409 37.021
R2580 B.n915 B.n405 37.021
R2581 B.n921 B.n405 37.021
R2582 B.n921 B.n401 37.021
R2583 B.n927 B.n401 37.021
R2584 B.n927 B.n397 37.021
R2585 B.n934 B.n397 37.021
R2586 B.n934 B.n933 37.021
R2587 B.n940 B.n390 37.021
R2588 B.n947 B.n390 37.021
R2589 B.n947 B.n386 37.021
R2590 B.n953 B.n386 37.021
R2591 B.n953 B.n4 37.021
R2592 B.n1155 B.n4 37.021
R2593 B.n1155 B.n1154 37.021
R2594 B.n1154 B.n1153 37.021
R2595 B.n1153 B.n8 37.021
R2596 B.n1147 B.n8 37.021
R2597 B.n1147 B.n1146 37.021
R2598 B.n1146 B.n1145 37.021
R2599 B.n1139 B.n18 37.021
R2600 B.n1139 B.n1138 37.021
R2601 B.n1138 B.n1137 37.021
R2602 B.n1137 B.n22 37.021
R2603 B.n1131 B.n22 37.021
R2604 B.n1131 B.n1130 37.021
R2605 B.n1130 B.n1129 37.021
R2606 B.n1129 B.n29 37.021
R2607 B.n1123 B.n29 37.021
R2608 B.n1122 B.n1121 37.021
R2609 B.n1121 B.n36 37.021
R2610 B.n1115 B.n36 37.021
R2611 B.n1115 B.n1114 37.021
R2612 B.n1114 B.n1113 37.021
R2613 B.n1113 B.n43 37.021
R2614 B.n1107 B.n43 37.021
R2615 B.n1107 B.n1106 37.021
R2616 B.n1106 B.n1105 37.021
R2617 B.n1099 B.n53 37.021
R2618 B.n1099 B.n1098 37.021
R2619 B.n1098 B.n1097 37.021
R2620 B.n1097 B.n57 37.021
R2621 B.n1091 B.n57 37.021
R2622 B.n1091 B.n1090 37.021
R2623 B.n1090 B.n1089 37.021
R2624 B.n1089 B.n64 37.021
R2625 B.n1083 B.n64 37.021
R2626 B.n1083 B.n1082 37.021
R2627 B.n1081 B.n71 37.021
R2628 B.n1075 B.n71 37.021
R2629 B.n1075 B.n1074 37.021
R2630 B.n1074 B.n1073 37.021
R2631 B.n1073 B.n78 37.021
R2632 B.n1067 B.n78 37.021
R2633 B.n1067 B.n1066 37.021
R2634 B.n1066 B.n1065 37.021
R2635 B.n1065 B.n85 37.021
R2636 B.n1059 B.n85 37.021
R2637 B.n1059 B.n1058 37.021
R2638 B.n1058 B.n1057 37.021
R2639 B.n1051 B.n95 37.021
R2640 B.n1051 B.n1050 37.021
R2641 B.n1050 B.n1049 37.021
R2642 B.n1049 B.n99 37.021
R2643 B.n1043 B.n99 37.021
R2644 B.n1043 B.n1042 37.021
R2645 B.n1042 B.n1041 37.021
R2646 B.n1041 B.n106 37.021
R2647 B.n879 B.t4 35.9322
R2648 B.n1105 B.t5 35.9322
R2649 B.n842 B.t2 32.6657
R2650 B.t0 B.n1081 32.6657
R2651 B.n1038 B.n1037 31.0639
R2652 B.n1031 B.n1030 31.0639
R2653 B.n558 B.n493 31.0639
R2654 B.n778 B.n777 31.0639
R2655 B.n909 B.t1 30.488
R2656 B.n1123 B.t3 30.488
R2657 B.n940 B.t7 25.0438
R2658 B.n1145 B.t6 25.0438
R2659 B.n799 B.t9 19.5996
R2660 B.n95 B.t13 19.5996
R2661 B B.n1157 18.0485
R2662 B.n806 B.t9 17.4219
R2663 B.n1057 B.t13 17.4219
R2664 B.n933 B.t7 11.9777
R2665 B.n18 B.t6 11.9777
R2666 B.n1037 B.n108 10.6151
R2667 B.n172 B.n108 10.6151
R2668 B.n173 B.n172 10.6151
R2669 B.n176 B.n173 10.6151
R2670 B.n177 B.n176 10.6151
R2671 B.n180 B.n177 10.6151
R2672 B.n181 B.n180 10.6151
R2673 B.n184 B.n181 10.6151
R2674 B.n185 B.n184 10.6151
R2675 B.n188 B.n185 10.6151
R2676 B.n189 B.n188 10.6151
R2677 B.n192 B.n189 10.6151
R2678 B.n193 B.n192 10.6151
R2679 B.n196 B.n193 10.6151
R2680 B.n197 B.n196 10.6151
R2681 B.n200 B.n197 10.6151
R2682 B.n201 B.n200 10.6151
R2683 B.n204 B.n201 10.6151
R2684 B.n205 B.n204 10.6151
R2685 B.n208 B.n205 10.6151
R2686 B.n209 B.n208 10.6151
R2687 B.n212 B.n209 10.6151
R2688 B.n213 B.n212 10.6151
R2689 B.n216 B.n213 10.6151
R2690 B.n217 B.n216 10.6151
R2691 B.n220 B.n217 10.6151
R2692 B.n221 B.n220 10.6151
R2693 B.n224 B.n221 10.6151
R2694 B.n225 B.n224 10.6151
R2695 B.n228 B.n225 10.6151
R2696 B.n229 B.n228 10.6151
R2697 B.n232 B.n229 10.6151
R2698 B.n233 B.n232 10.6151
R2699 B.n236 B.n233 10.6151
R2700 B.n237 B.n236 10.6151
R2701 B.n240 B.n237 10.6151
R2702 B.n241 B.n240 10.6151
R2703 B.n244 B.n241 10.6151
R2704 B.n245 B.n244 10.6151
R2705 B.n248 B.n245 10.6151
R2706 B.n249 B.n248 10.6151
R2707 B.n252 B.n249 10.6151
R2708 B.n253 B.n252 10.6151
R2709 B.n256 B.n253 10.6151
R2710 B.n257 B.n256 10.6151
R2711 B.n260 B.n257 10.6151
R2712 B.n261 B.n260 10.6151
R2713 B.n264 B.n261 10.6151
R2714 B.n265 B.n264 10.6151
R2715 B.n269 B.n268 10.6151
R2716 B.n272 B.n269 10.6151
R2717 B.n273 B.n272 10.6151
R2718 B.n276 B.n273 10.6151
R2719 B.n277 B.n276 10.6151
R2720 B.n280 B.n277 10.6151
R2721 B.n281 B.n280 10.6151
R2722 B.n284 B.n281 10.6151
R2723 B.n285 B.n284 10.6151
R2724 B.n289 B.n288 10.6151
R2725 B.n292 B.n289 10.6151
R2726 B.n293 B.n292 10.6151
R2727 B.n296 B.n293 10.6151
R2728 B.n297 B.n296 10.6151
R2729 B.n300 B.n297 10.6151
R2730 B.n301 B.n300 10.6151
R2731 B.n304 B.n301 10.6151
R2732 B.n305 B.n304 10.6151
R2733 B.n308 B.n305 10.6151
R2734 B.n309 B.n308 10.6151
R2735 B.n312 B.n309 10.6151
R2736 B.n313 B.n312 10.6151
R2737 B.n316 B.n313 10.6151
R2738 B.n317 B.n316 10.6151
R2739 B.n320 B.n317 10.6151
R2740 B.n321 B.n320 10.6151
R2741 B.n324 B.n321 10.6151
R2742 B.n325 B.n324 10.6151
R2743 B.n328 B.n325 10.6151
R2744 B.n329 B.n328 10.6151
R2745 B.n332 B.n329 10.6151
R2746 B.n333 B.n332 10.6151
R2747 B.n336 B.n333 10.6151
R2748 B.n337 B.n336 10.6151
R2749 B.n340 B.n337 10.6151
R2750 B.n341 B.n340 10.6151
R2751 B.n344 B.n341 10.6151
R2752 B.n345 B.n344 10.6151
R2753 B.n348 B.n345 10.6151
R2754 B.n349 B.n348 10.6151
R2755 B.n352 B.n349 10.6151
R2756 B.n353 B.n352 10.6151
R2757 B.n356 B.n353 10.6151
R2758 B.n357 B.n356 10.6151
R2759 B.n360 B.n357 10.6151
R2760 B.n361 B.n360 10.6151
R2761 B.n364 B.n361 10.6151
R2762 B.n365 B.n364 10.6151
R2763 B.n368 B.n365 10.6151
R2764 B.n369 B.n368 10.6151
R2765 B.n372 B.n369 10.6151
R2766 B.n373 B.n372 10.6151
R2767 B.n376 B.n373 10.6151
R2768 B.n377 B.n376 10.6151
R2769 B.n380 B.n377 10.6151
R2770 B.n382 B.n380 10.6151
R2771 B.n383 B.n382 10.6151
R2772 B.n1031 B.n383 10.6151
R2773 B.n783 B.n493 10.6151
R2774 B.n784 B.n783 10.6151
R2775 B.n785 B.n784 10.6151
R2776 B.n785 B.n485 10.6151
R2777 B.n795 B.n485 10.6151
R2778 B.n796 B.n795 10.6151
R2779 B.n797 B.n796 10.6151
R2780 B.n797 B.n478 10.6151
R2781 B.n808 B.n478 10.6151
R2782 B.n809 B.n808 10.6151
R2783 B.n810 B.n809 10.6151
R2784 B.n810 B.n470 10.6151
R2785 B.n820 B.n470 10.6151
R2786 B.n821 B.n820 10.6151
R2787 B.n822 B.n821 10.6151
R2788 B.n822 B.n462 10.6151
R2789 B.n832 B.n462 10.6151
R2790 B.n833 B.n832 10.6151
R2791 B.n834 B.n833 10.6151
R2792 B.n834 B.n454 10.6151
R2793 B.n844 B.n454 10.6151
R2794 B.n845 B.n844 10.6151
R2795 B.n846 B.n845 10.6151
R2796 B.n846 B.n446 10.6151
R2797 B.n856 B.n446 10.6151
R2798 B.n857 B.n856 10.6151
R2799 B.n858 B.n857 10.6151
R2800 B.n858 B.n438 10.6151
R2801 B.n868 B.n438 10.6151
R2802 B.n869 B.n868 10.6151
R2803 B.n870 B.n869 10.6151
R2804 B.n870 B.n431 10.6151
R2805 B.n881 B.n431 10.6151
R2806 B.n882 B.n881 10.6151
R2807 B.n883 B.n882 10.6151
R2808 B.n883 B.n423 10.6151
R2809 B.n893 B.n423 10.6151
R2810 B.n894 B.n893 10.6151
R2811 B.n895 B.n894 10.6151
R2812 B.n895 B.n414 10.6151
R2813 B.n905 B.n414 10.6151
R2814 B.n906 B.n905 10.6151
R2815 B.n907 B.n906 10.6151
R2816 B.n907 B.n407 10.6151
R2817 B.n917 B.n407 10.6151
R2818 B.n918 B.n917 10.6151
R2819 B.n919 B.n918 10.6151
R2820 B.n919 B.n399 10.6151
R2821 B.n929 B.n399 10.6151
R2822 B.n930 B.n929 10.6151
R2823 B.n931 B.n930 10.6151
R2824 B.n931 B.n392 10.6151
R2825 B.n942 B.n392 10.6151
R2826 B.n943 B.n942 10.6151
R2827 B.n945 B.n943 10.6151
R2828 B.n945 B.n944 10.6151
R2829 B.n944 B.n384 10.6151
R2830 B.n956 B.n384 10.6151
R2831 B.n957 B.n956 10.6151
R2832 B.n958 B.n957 10.6151
R2833 B.n959 B.n958 10.6151
R2834 B.n961 B.n959 10.6151
R2835 B.n962 B.n961 10.6151
R2836 B.n963 B.n962 10.6151
R2837 B.n964 B.n963 10.6151
R2838 B.n966 B.n964 10.6151
R2839 B.n967 B.n966 10.6151
R2840 B.n968 B.n967 10.6151
R2841 B.n969 B.n968 10.6151
R2842 B.n971 B.n969 10.6151
R2843 B.n972 B.n971 10.6151
R2844 B.n973 B.n972 10.6151
R2845 B.n974 B.n973 10.6151
R2846 B.n976 B.n974 10.6151
R2847 B.n977 B.n976 10.6151
R2848 B.n978 B.n977 10.6151
R2849 B.n979 B.n978 10.6151
R2850 B.n981 B.n979 10.6151
R2851 B.n982 B.n981 10.6151
R2852 B.n983 B.n982 10.6151
R2853 B.n984 B.n983 10.6151
R2854 B.n986 B.n984 10.6151
R2855 B.n987 B.n986 10.6151
R2856 B.n988 B.n987 10.6151
R2857 B.n989 B.n988 10.6151
R2858 B.n991 B.n989 10.6151
R2859 B.n992 B.n991 10.6151
R2860 B.n993 B.n992 10.6151
R2861 B.n994 B.n993 10.6151
R2862 B.n996 B.n994 10.6151
R2863 B.n997 B.n996 10.6151
R2864 B.n998 B.n997 10.6151
R2865 B.n999 B.n998 10.6151
R2866 B.n1001 B.n999 10.6151
R2867 B.n1002 B.n1001 10.6151
R2868 B.n1003 B.n1002 10.6151
R2869 B.n1004 B.n1003 10.6151
R2870 B.n1006 B.n1004 10.6151
R2871 B.n1007 B.n1006 10.6151
R2872 B.n1008 B.n1007 10.6151
R2873 B.n1009 B.n1008 10.6151
R2874 B.n1011 B.n1009 10.6151
R2875 B.n1012 B.n1011 10.6151
R2876 B.n1013 B.n1012 10.6151
R2877 B.n1014 B.n1013 10.6151
R2878 B.n1016 B.n1014 10.6151
R2879 B.n1017 B.n1016 10.6151
R2880 B.n1018 B.n1017 10.6151
R2881 B.n1019 B.n1018 10.6151
R2882 B.n1021 B.n1019 10.6151
R2883 B.n1022 B.n1021 10.6151
R2884 B.n1023 B.n1022 10.6151
R2885 B.n1024 B.n1023 10.6151
R2886 B.n1026 B.n1024 10.6151
R2887 B.n1027 B.n1026 10.6151
R2888 B.n1028 B.n1027 10.6151
R2889 B.n1029 B.n1028 10.6151
R2890 B.n1030 B.n1029 10.6151
R2891 B.n777 B.n497 10.6151
R2892 B.n772 B.n497 10.6151
R2893 B.n772 B.n771 10.6151
R2894 B.n771 B.n770 10.6151
R2895 B.n770 B.n767 10.6151
R2896 B.n767 B.n766 10.6151
R2897 B.n766 B.n763 10.6151
R2898 B.n763 B.n762 10.6151
R2899 B.n762 B.n759 10.6151
R2900 B.n759 B.n758 10.6151
R2901 B.n758 B.n755 10.6151
R2902 B.n755 B.n754 10.6151
R2903 B.n754 B.n751 10.6151
R2904 B.n751 B.n750 10.6151
R2905 B.n750 B.n747 10.6151
R2906 B.n747 B.n746 10.6151
R2907 B.n746 B.n743 10.6151
R2908 B.n743 B.n742 10.6151
R2909 B.n742 B.n739 10.6151
R2910 B.n739 B.n738 10.6151
R2911 B.n738 B.n735 10.6151
R2912 B.n735 B.n734 10.6151
R2913 B.n734 B.n731 10.6151
R2914 B.n731 B.n730 10.6151
R2915 B.n730 B.n727 10.6151
R2916 B.n727 B.n726 10.6151
R2917 B.n726 B.n723 10.6151
R2918 B.n723 B.n722 10.6151
R2919 B.n722 B.n719 10.6151
R2920 B.n719 B.n718 10.6151
R2921 B.n718 B.n715 10.6151
R2922 B.n715 B.n714 10.6151
R2923 B.n714 B.n711 10.6151
R2924 B.n711 B.n710 10.6151
R2925 B.n710 B.n707 10.6151
R2926 B.n707 B.n706 10.6151
R2927 B.n706 B.n703 10.6151
R2928 B.n703 B.n702 10.6151
R2929 B.n702 B.n699 10.6151
R2930 B.n699 B.n698 10.6151
R2931 B.n698 B.n695 10.6151
R2932 B.n695 B.n694 10.6151
R2933 B.n694 B.n691 10.6151
R2934 B.n691 B.n690 10.6151
R2935 B.n690 B.n687 10.6151
R2936 B.n687 B.n686 10.6151
R2937 B.n686 B.n683 10.6151
R2938 B.n683 B.n682 10.6151
R2939 B.n682 B.n679 10.6151
R2940 B.n677 B.n674 10.6151
R2941 B.n674 B.n673 10.6151
R2942 B.n673 B.n670 10.6151
R2943 B.n670 B.n669 10.6151
R2944 B.n669 B.n666 10.6151
R2945 B.n666 B.n665 10.6151
R2946 B.n665 B.n662 10.6151
R2947 B.n662 B.n661 10.6151
R2948 B.n661 B.n658 10.6151
R2949 B.n656 B.n653 10.6151
R2950 B.n653 B.n652 10.6151
R2951 B.n652 B.n649 10.6151
R2952 B.n649 B.n648 10.6151
R2953 B.n648 B.n645 10.6151
R2954 B.n645 B.n644 10.6151
R2955 B.n644 B.n641 10.6151
R2956 B.n641 B.n640 10.6151
R2957 B.n640 B.n637 10.6151
R2958 B.n637 B.n636 10.6151
R2959 B.n636 B.n633 10.6151
R2960 B.n633 B.n632 10.6151
R2961 B.n632 B.n629 10.6151
R2962 B.n629 B.n628 10.6151
R2963 B.n628 B.n625 10.6151
R2964 B.n625 B.n624 10.6151
R2965 B.n624 B.n621 10.6151
R2966 B.n621 B.n620 10.6151
R2967 B.n620 B.n617 10.6151
R2968 B.n617 B.n616 10.6151
R2969 B.n616 B.n613 10.6151
R2970 B.n613 B.n612 10.6151
R2971 B.n612 B.n609 10.6151
R2972 B.n609 B.n608 10.6151
R2973 B.n608 B.n605 10.6151
R2974 B.n605 B.n604 10.6151
R2975 B.n604 B.n601 10.6151
R2976 B.n601 B.n600 10.6151
R2977 B.n600 B.n597 10.6151
R2978 B.n597 B.n596 10.6151
R2979 B.n596 B.n593 10.6151
R2980 B.n593 B.n592 10.6151
R2981 B.n592 B.n589 10.6151
R2982 B.n589 B.n588 10.6151
R2983 B.n588 B.n585 10.6151
R2984 B.n585 B.n584 10.6151
R2985 B.n584 B.n581 10.6151
R2986 B.n581 B.n580 10.6151
R2987 B.n580 B.n577 10.6151
R2988 B.n577 B.n576 10.6151
R2989 B.n576 B.n573 10.6151
R2990 B.n573 B.n572 10.6151
R2991 B.n572 B.n569 10.6151
R2992 B.n569 B.n568 10.6151
R2993 B.n568 B.n565 10.6151
R2994 B.n565 B.n564 10.6151
R2995 B.n564 B.n561 10.6151
R2996 B.n561 B.n560 10.6151
R2997 B.n560 B.n558 10.6151
R2998 B.n779 B.n778 10.6151
R2999 B.n779 B.n489 10.6151
R3000 B.n789 B.n489 10.6151
R3001 B.n790 B.n789 10.6151
R3002 B.n791 B.n790 10.6151
R3003 B.n791 B.n481 10.6151
R3004 B.n802 B.n481 10.6151
R3005 B.n803 B.n802 10.6151
R3006 B.n804 B.n803 10.6151
R3007 B.n804 B.n474 10.6151
R3008 B.n814 B.n474 10.6151
R3009 B.n815 B.n814 10.6151
R3010 B.n816 B.n815 10.6151
R3011 B.n816 B.n466 10.6151
R3012 B.n826 B.n466 10.6151
R3013 B.n827 B.n826 10.6151
R3014 B.n828 B.n827 10.6151
R3015 B.n828 B.n458 10.6151
R3016 B.n838 B.n458 10.6151
R3017 B.n839 B.n838 10.6151
R3018 B.n840 B.n839 10.6151
R3019 B.n840 B.n450 10.6151
R3020 B.n850 B.n450 10.6151
R3021 B.n851 B.n850 10.6151
R3022 B.n852 B.n851 10.6151
R3023 B.n852 B.n442 10.6151
R3024 B.n862 B.n442 10.6151
R3025 B.n863 B.n862 10.6151
R3026 B.n864 B.n863 10.6151
R3027 B.n864 B.n434 10.6151
R3028 B.n875 B.n434 10.6151
R3029 B.n876 B.n875 10.6151
R3030 B.n877 B.n876 10.6151
R3031 B.n877 B.n427 10.6151
R3032 B.n887 B.n427 10.6151
R3033 B.n888 B.n887 10.6151
R3034 B.n889 B.n888 10.6151
R3035 B.n889 B.n419 10.6151
R3036 B.n899 B.n419 10.6151
R3037 B.n900 B.n899 10.6151
R3038 B.n901 B.n900 10.6151
R3039 B.n901 B.n411 10.6151
R3040 B.n911 B.n411 10.6151
R3041 B.n912 B.n911 10.6151
R3042 B.n913 B.n912 10.6151
R3043 B.n913 B.n403 10.6151
R3044 B.n923 B.n403 10.6151
R3045 B.n924 B.n923 10.6151
R3046 B.n925 B.n924 10.6151
R3047 B.n925 B.n395 10.6151
R3048 B.n936 B.n395 10.6151
R3049 B.n937 B.n936 10.6151
R3050 B.n938 B.n937 10.6151
R3051 B.n938 B.n388 10.6151
R3052 B.n949 B.n388 10.6151
R3053 B.n950 B.n949 10.6151
R3054 B.n951 B.n950 10.6151
R3055 B.n951 B.n0 10.6151
R3056 B.n1151 B.n1 10.6151
R3057 B.n1151 B.n1150 10.6151
R3058 B.n1150 B.n1149 10.6151
R3059 B.n1149 B.n10 10.6151
R3060 B.n1143 B.n10 10.6151
R3061 B.n1143 B.n1142 10.6151
R3062 B.n1142 B.n1141 10.6151
R3063 B.n1141 B.n16 10.6151
R3064 B.n1135 B.n16 10.6151
R3065 B.n1135 B.n1134 10.6151
R3066 B.n1134 B.n1133 10.6151
R3067 B.n1133 B.n24 10.6151
R3068 B.n1127 B.n24 10.6151
R3069 B.n1127 B.n1126 10.6151
R3070 B.n1126 B.n1125 10.6151
R3071 B.n1125 B.n31 10.6151
R3072 B.n1119 B.n31 10.6151
R3073 B.n1119 B.n1118 10.6151
R3074 B.n1118 B.n1117 10.6151
R3075 B.n1117 B.n38 10.6151
R3076 B.n1111 B.n38 10.6151
R3077 B.n1111 B.n1110 10.6151
R3078 B.n1110 B.n1109 10.6151
R3079 B.n1109 B.n45 10.6151
R3080 B.n1103 B.n45 10.6151
R3081 B.n1103 B.n1102 10.6151
R3082 B.n1102 B.n1101 10.6151
R3083 B.n1101 B.n51 10.6151
R3084 B.n1095 B.n51 10.6151
R3085 B.n1095 B.n1094 10.6151
R3086 B.n1094 B.n1093 10.6151
R3087 B.n1093 B.n59 10.6151
R3088 B.n1087 B.n59 10.6151
R3089 B.n1087 B.n1086 10.6151
R3090 B.n1086 B.n1085 10.6151
R3091 B.n1085 B.n66 10.6151
R3092 B.n1079 B.n66 10.6151
R3093 B.n1079 B.n1078 10.6151
R3094 B.n1078 B.n1077 10.6151
R3095 B.n1077 B.n73 10.6151
R3096 B.n1071 B.n73 10.6151
R3097 B.n1071 B.n1070 10.6151
R3098 B.n1070 B.n1069 10.6151
R3099 B.n1069 B.n80 10.6151
R3100 B.n1063 B.n80 10.6151
R3101 B.n1063 B.n1062 10.6151
R3102 B.n1062 B.n1061 10.6151
R3103 B.n1061 B.n87 10.6151
R3104 B.n1055 B.n87 10.6151
R3105 B.n1055 B.n1054 10.6151
R3106 B.n1054 B.n1053 10.6151
R3107 B.n1053 B.n93 10.6151
R3108 B.n1047 B.n93 10.6151
R3109 B.n1047 B.n1046 10.6151
R3110 B.n1046 B.n1045 10.6151
R3111 B.n1045 B.n101 10.6151
R3112 B.n1039 B.n101 10.6151
R3113 B.n1039 B.n1038 10.6151
R3114 B.n265 B.n170 9.36635
R3115 B.n288 B.n167 9.36635
R3116 B.n679 B.n678 9.36635
R3117 B.n657 B.n656 9.36635
R3118 B.n417 B.t1 6.53354
R3119 B.t3 B.n1122 6.53354
R3120 B.t2 B.n452 4.35586
R3121 B.n1082 B.t0 4.35586
R3122 B.n1157 B.n0 2.81026
R3123 B.n1157 B.n1 2.81026
R3124 B.n268 B.n170 1.24928
R3125 B.n285 B.n167 1.24928
R3126 B.n678 B.n677 1.24928
R3127 B.n658 B.n657 1.24928
R3128 B.n872 B.t4 1.08934
R3129 B.n53 B.t5 1.08934
R3130 VN.n60 VN.n59 161.3
R3131 VN.n58 VN.n32 161.3
R3132 VN.n57 VN.n56 161.3
R3133 VN.n55 VN.n33 161.3
R3134 VN.n54 VN.n53 161.3
R3135 VN.n52 VN.n34 161.3
R3136 VN.n51 VN.n50 161.3
R3137 VN.n49 VN.n48 161.3
R3138 VN.n47 VN.n36 161.3
R3139 VN.n46 VN.n45 161.3
R3140 VN.n44 VN.n37 161.3
R3141 VN.n43 VN.n42 161.3
R3142 VN.n41 VN.n38 161.3
R3143 VN.n29 VN.n28 161.3
R3144 VN.n27 VN.n1 161.3
R3145 VN.n26 VN.n25 161.3
R3146 VN.n24 VN.n2 161.3
R3147 VN.n23 VN.n22 161.3
R3148 VN.n21 VN.n3 161.3
R3149 VN.n20 VN.n19 161.3
R3150 VN.n18 VN.n17 161.3
R3151 VN.n16 VN.n5 161.3
R3152 VN.n15 VN.n14 161.3
R3153 VN.n13 VN.n6 161.3
R3154 VN.n12 VN.n11 161.3
R3155 VN.n10 VN.n7 161.3
R3156 VN.n39 VN.t3 148.738
R3157 VN.n8 VN.t1 148.738
R3158 VN.n9 VN.t4 115.326
R3159 VN.n4 VN.t2 115.326
R3160 VN.n0 VN.t5 115.326
R3161 VN.n40 VN.t6 115.326
R3162 VN.n35 VN.t0 115.326
R3163 VN.n31 VN.t7 115.326
R3164 VN.n30 VN.n0 69.2705
R3165 VN.n61 VN.n31 69.2705
R3166 VN.n15 VN.n6 56.5193
R3167 VN.n26 VN.n2 56.5193
R3168 VN.n46 VN.n37 56.5193
R3169 VN.n57 VN.n33 56.5193
R3170 VN VN.n61 55.8768
R3171 VN.n9 VN.n8 50.6608
R3172 VN.n40 VN.n39 50.6608
R3173 VN.n11 VN.n10 24.4675
R3174 VN.n11 VN.n6 24.4675
R3175 VN.n16 VN.n15 24.4675
R3176 VN.n17 VN.n16 24.4675
R3177 VN.n21 VN.n20 24.4675
R3178 VN.n22 VN.n21 24.4675
R3179 VN.n22 VN.n2 24.4675
R3180 VN.n27 VN.n26 24.4675
R3181 VN.n28 VN.n27 24.4675
R3182 VN.n42 VN.n37 24.4675
R3183 VN.n42 VN.n41 24.4675
R3184 VN.n53 VN.n33 24.4675
R3185 VN.n53 VN.n52 24.4675
R3186 VN.n52 VN.n51 24.4675
R3187 VN.n48 VN.n47 24.4675
R3188 VN.n47 VN.n46 24.4675
R3189 VN.n59 VN.n58 24.4675
R3190 VN.n58 VN.n57 24.4675
R3191 VN.n10 VN.n9 23.2442
R3192 VN.n17 VN.n4 23.2442
R3193 VN.n41 VN.n40 23.2442
R3194 VN.n48 VN.n35 23.2442
R3195 VN.n28 VN.n0 20.7975
R3196 VN.n59 VN.n31 20.7975
R3197 VN.n39 VN.n38 3.87633
R3198 VN.n8 VN.n7 3.87633
R3199 VN.n20 VN.n4 1.22385
R3200 VN.n51 VN.n35 1.22385
R3201 VN.n61 VN.n60 0.354971
R3202 VN.n30 VN.n29 0.354971
R3203 VN VN.n30 0.26696
R3204 VN.n60 VN.n32 0.189894
R3205 VN.n56 VN.n32 0.189894
R3206 VN.n56 VN.n55 0.189894
R3207 VN.n55 VN.n54 0.189894
R3208 VN.n54 VN.n34 0.189894
R3209 VN.n50 VN.n34 0.189894
R3210 VN.n50 VN.n49 0.189894
R3211 VN.n49 VN.n36 0.189894
R3212 VN.n45 VN.n36 0.189894
R3213 VN.n45 VN.n44 0.189894
R3214 VN.n44 VN.n43 0.189894
R3215 VN.n43 VN.n38 0.189894
R3216 VN.n12 VN.n7 0.189894
R3217 VN.n13 VN.n12 0.189894
R3218 VN.n14 VN.n13 0.189894
R3219 VN.n14 VN.n5 0.189894
R3220 VN.n18 VN.n5 0.189894
R3221 VN.n19 VN.n18 0.189894
R3222 VN.n19 VN.n3 0.189894
R3223 VN.n23 VN.n3 0.189894
R3224 VN.n24 VN.n23 0.189894
R3225 VN.n25 VN.n24 0.189894
R3226 VN.n25 VN.n1 0.189894
R3227 VN.n29 VN.n1 0.189894
R3228 VDD2.n2 VDD2.n1 61.3956
R3229 VDD2.n2 VDD2.n0 61.3956
R3230 VDD2 VDD2.n5 61.393
R3231 VDD2.n4 VDD2.n3 59.9641
R3232 VDD2.n4 VDD2.n2 49.9696
R3233 VDD2 VDD2.n4 1.54576
R3234 VDD2.n5 VDD2.t1 1.32669
R3235 VDD2.n5 VDD2.t4 1.32669
R3236 VDD2.n3 VDD2.t0 1.32669
R3237 VDD2.n3 VDD2.t7 1.32669
R3238 VDD2.n1 VDD2.t5 1.32669
R3239 VDD2.n1 VDD2.t2 1.32669
R3240 VDD2.n0 VDD2.t6 1.32669
R3241 VDD2.n0 VDD2.t3 1.32669
C0 VDD1 VTAIL 9.13677f
C1 VDD2 VN 11.0618f
C2 VDD1 VDD2 2.04916f
C3 VP VN 8.84095f
C4 VDD1 VP 11.482401f
C5 VDD2 VTAIL 9.19467f
C6 VP VTAIL 11.5151f
C7 VDD2 VP 0.575128f
C8 VDD1 VN 0.152792f
C9 VN VTAIL 11.500999f
C10 VDD2 B 6.152263f
C11 VDD1 B 6.642333f
C12 VTAIL B 12.609422f
C13 VN B 17.738201f
C14 VP B 16.334562f
C15 VDD2.t6 B 0.313674f
C16 VDD2.t3 B 0.313674f
C17 VDD2.n0 B 2.84069f
C18 VDD2.t5 B 0.313674f
C19 VDD2.t2 B 0.313674f
C20 VDD2.n1 B 2.84069f
C21 VDD2.n2 B 4.01548f
C22 VDD2.t0 B 0.313674f
C23 VDD2.t7 B 0.313674f
C24 VDD2.n3 B 2.82637f
C25 VDD2.n4 B 3.57238f
C26 VDD2.t1 B 0.313674f
C27 VDD2.t4 B 0.313674f
C28 VDD2.n5 B 2.84066f
C29 VN.t5 B 2.43872f
C30 VN.n0 B 0.928299f
C31 VN.n1 B 0.019108f
C32 VN.n2 B 0.025232f
C33 VN.n3 B 0.019108f
C34 VN.t2 B 2.43872f
C35 VN.n4 B 0.849049f
C36 VN.n5 B 0.019108f
C37 VN.n6 B 0.027894f
C38 VN.n7 B 0.217948f
C39 VN.t4 B 2.43872f
C40 VN.t1 B 2.66027f
C41 VN.n8 B 0.877333f
C42 VN.n9 B 0.919909f
C43 VN.n10 B 0.034732f
C44 VN.n11 B 0.035612f
C45 VN.n12 B 0.019108f
C46 VN.n13 B 0.019108f
C47 VN.n14 B 0.019108f
C48 VN.n15 B 0.027894f
C49 VN.n16 B 0.035612f
C50 VN.n17 B 0.034732f
C51 VN.n18 B 0.019108f
C52 VN.n19 B 0.019108f
C53 VN.n20 B 0.018909f
C54 VN.n21 B 0.035612f
C55 VN.n22 B 0.035612f
C56 VN.n23 B 0.019108f
C57 VN.n24 B 0.019108f
C58 VN.n25 B 0.019108f
C59 VN.n26 B 0.030556f
C60 VN.n27 B 0.035612f
C61 VN.n28 B 0.032974f
C62 VN.n29 B 0.03084f
C63 VN.n30 B 0.039786f
C64 VN.t7 B 2.43872f
C65 VN.n31 B 0.928299f
C66 VN.n32 B 0.019108f
C67 VN.n33 B 0.025232f
C68 VN.n34 B 0.019108f
C69 VN.t0 B 2.43872f
C70 VN.n35 B 0.849049f
C71 VN.n36 B 0.019108f
C72 VN.n37 B 0.027894f
C73 VN.n38 B 0.217948f
C74 VN.t6 B 2.43872f
C75 VN.t3 B 2.66027f
C76 VN.n39 B 0.877333f
C77 VN.n40 B 0.919909f
C78 VN.n41 B 0.034732f
C79 VN.n42 B 0.035612f
C80 VN.n43 B 0.019108f
C81 VN.n44 B 0.019108f
C82 VN.n45 B 0.019108f
C83 VN.n46 B 0.027894f
C84 VN.n47 B 0.035612f
C85 VN.n48 B 0.034732f
C86 VN.n49 B 0.019108f
C87 VN.n50 B 0.019108f
C88 VN.n51 B 0.018909f
C89 VN.n52 B 0.035612f
C90 VN.n53 B 0.035612f
C91 VN.n54 B 0.019108f
C92 VN.n55 B 0.019108f
C93 VN.n56 B 0.019108f
C94 VN.n57 B 0.030556f
C95 VN.n58 B 0.035612f
C96 VN.n59 B 0.032974f
C97 VN.n60 B 0.03084f
C98 VN.n61 B 1.26697f
C99 VDD1.t0 B 0.3165f
C100 VDD1.t7 B 0.3165f
C101 VDD1.n0 B 2.86765f
C102 VDD1.t3 B 0.3165f
C103 VDD1.t5 B 0.3165f
C104 VDD1.n1 B 2.86629f
C105 VDD1.t2 B 0.3165f
C106 VDD1.t6 B 0.3165f
C107 VDD1.n2 B 2.86629f
C108 VDD1.n3 B 4.10711f
C109 VDD1.t1 B 0.3165f
C110 VDD1.t4 B 0.3165f
C111 VDD1.n4 B 2.85184f
C112 VDD1.n5 B 3.63813f
C113 VTAIL.t3 B 0.228644f
C114 VTAIL.t5 B 0.228644f
C115 VTAIL.n0 B 1.99816f
C116 VTAIL.n1 B 0.389749f
C117 VTAIL.n2 B 0.028417f
C118 VTAIL.n3 B 0.01938f
C119 VTAIL.n4 B 0.010414f
C120 VTAIL.n5 B 0.024614f
C121 VTAIL.n6 B 0.011026f
C122 VTAIL.n7 B 0.01938f
C123 VTAIL.n8 B 0.010414f
C124 VTAIL.n9 B 0.024614f
C125 VTAIL.n10 B 0.011026f
C126 VTAIL.n11 B 0.01938f
C127 VTAIL.n12 B 0.010414f
C128 VTAIL.n13 B 0.024614f
C129 VTAIL.n14 B 0.011026f
C130 VTAIL.n15 B 0.01938f
C131 VTAIL.n16 B 0.010414f
C132 VTAIL.n17 B 0.024614f
C133 VTAIL.n18 B 0.011026f
C134 VTAIL.n19 B 0.01938f
C135 VTAIL.n20 B 0.010414f
C136 VTAIL.n21 B 0.024614f
C137 VTAIL.n22 B 0.011026f
C138 VTAIL.n23 B 0.01938f
C139 VTAIL.n24 B 0.010414f
C140 VTAIL.n25 B 0.024614f
C141 VTAIL.n26 B 0.011026f
C142 VTAIL.n27 B 0.161525f
C143 VTAIL.t15 B 0.041878f
C144 VTAIL.n28 B 0.018461f
C145 VTAIL.n29 B 0.0174f
C146 VTAIL.n30 B 0.010414f
C147 VTAIL.n31 B 1.23023f
C148 VTAIL.n32 B 0.01938f
C149 VTAIL.n33 B 0.010414f
C150 VTAIL.n34 B 0.011026f
C151 VTAIL.n35 B 0.024614f
C152 VTAIL.n36 B 0.024614f
C153 VTAIL.n37 B 0.011026f
C154 VTAIL.n38 B 0.010414f
C155 VTAIL.n39 B 0.01938f
C156 VTAIL.n40 B 0.01938f
C157 VTAIL.n41 B 0.010414f
C158 VTAIL.n42 B 0.011026f
C159 VTAIL.n43 B 0.024614f
C160 VTAIL.n44 B 0.024614f
C161 VTAIL.n45 B 0.024614f
C162 VTAIL.n46 B 0.011026f
C163 VTAIL.n47 B 0.010414f
C164 VTAIL.n48 B 0.01938f
C165 VTAIL.n49 B 0.01938f
C166 VTAIL.n50 B 0.010414f
C167 VTAIL.n51 B 0.01072f
C168 VTAIL.n52 B 0.01072f
C169 VTAIL.n53 B 0.024614f
C170 VTAIL.n54 B 0.024614f
C171 VTAIL.n55 B 0.011026f
C172 VTAIL.n56 B 0.010414f
C173 VTAIL.n57 B 0.01938f
C174 VTAIL.n58 B 0.01938f
C175 VTAIL.n59 B 0.010414f
C176 VTAIL.n60 B 0.011026f
C177 VTAIL.n61 B 0.024614f
C178 VTAIL.n62 B 0.024614f
C179 VTAIL.n63 B 0.011026f
C180 VTAIL.n64 B 0.010414f
C181 VTAIL.n65 B 0.01938f
C182 VTAIL.n66 B 0.01938f
C183 VTAIL.n67 B 0.010414f
C184 VTAIL.n68 B 0.011026f
C185 VTAIL.n69 B 0.024614f
C186 VTAIL.n70 B 0.024614f
C187 VTAIL.n71 B 0.011026f
C188 VTAIL.n72 B 0.010414f
C189 VTAIL.n73 B 0.01938f
C190 VTAIL.n74 B 0.01938f
C191 VTAIL.n75 B 0.010414f
C192 VTAIL.n76 B 0.011026f
C193 VTAIL.n77 B 0.024614f
C194 VTAIL.n78 B 0.055367f
C195 VTAIL.n79 B 0.011026f
C196 VTAIL.n80 B 0.010414f
C197 VTAIL.n81 B 0.042942f
C198 VTAIL.n82 B 0.031136f
C199 VTAIL.n83 B 0.230567f
C200 VTAIL.n84 B 0.028417f
C201 VTAIL.n85 B 0.01938f
C202 VTAIL.n86 B 0.010414f
C203 VTAIL.n87 B 0.024614f
C204 VTAIL.n88 B 0.011026f
C205 VTAIL.n89 B 0.01938f
C206 VTAIL.n90 B 0.010414f
C207 VTAIL.n91 B 0.024614f
C208 VTAIL.n92 B 0.011026f
C209 VTAIL.n93 B 0.01938f
C210 VTAIL.n94 B 0.010414f
C211 VTAIL.n95 B 0.024614f
C212 VTAIL.n96 B 0.011026f
C213 VTAIL.n97 B 0.01938f
C214 VTAIL.n98 B 0.010414f
C215 VTAIL.n99 B 0.024614f
C216 VTAIL.n100 B 0.011026f
C217 VTAIL.n101 B 0.01938f
C218 VTAIL.n102 B 0.010414f
C219 VTAIL.n103 B 0.024614f
C220 VTAIL.n104 B 0.011026f
C221 VTAIL.n105 B 0.01938f
C222 VTAIL.n106 B 0.010414f
C223 VTAIL.n107 B 0.024614f
C224 VTAIL.n108 B 0.011026f
C225 VTAIL.n109 B 0.161525f
C226 VTAIL.t11 B 0.041878f
C227 VTAIL.n110 B 0.018461f
C228 VTAIL.n111 B 0.0174f
C229 VTAIL.n112 B 0.010414f
C230 VTAIL.n113 B 1.23023f
C231 VTAIL.n114 B 0.01938f
C232 VTAIL.n115 B 0.010414f
C233 VTAIL.n116 B 0.011026f
C234 VTAIL.n117 B 0.024614f
C235 VTAIL.n118 B 0.024614f
C236 VTAIL.n119 B 0.011026f
C237 VTAIL.n120 B 0.010414f
C238 VTAIL.n121 B 0.01938f
C239 VTAIL.n122 B 0.01938f
C240 VTAIL.n123 B 0.010414f
C241 VTAIL.n124 B 0.011026f
C242 VTAIL.n125 B 0.024614f
C243 VTAIL.n126 B 0.024614f
C244 VTAIL.n127 B 0.024614f
C245 VTAIL.n128 B 0.011026f
C246 VTAIL.n129 B 0.010414f
C247 VTAIL.n130 B 0.01938f
C248 VTAIL.n131 B 0.01938f
C249 VTAIL.n132 B 0.010414f
C250 VTAIL.n133 B 0.01072f
C251 VTAIL.n134 B 0.01072f
C252 VTAIL.n135 B 0.024614f
C253 VTAIL.n136 B 0.024614f
C254 VTAIL.n137 B 0.011026f
C255 VTAIL.n138 B 0.010414f
C256 VTAIL.n139 B 0.01938f
C257 VTAIL.n140 B 0.01938f
C258 VTAIL.n141 B 0.010414f
C259 VTAIL.n142 B 0.011026f
C260 VTAIL.n143 B 0.024614f
C261 VTAIL.n144 B 0.024614f
C262 VTAIL.n145 B 0.011026f
C263 VTAIL.n146 B 0.010414f
C264 VTAIL.n147 B 0.01938f
C265 VTAIL.n148 B 0.01938f
C266 VTAIL.n149 B 0.010414f
C267 VTAIL.n150 B 0.011026f
C268 VTAIL.n151 B 0.024614f
C269 VTAIL.n152 B 0.024614f
C270 VTAIL.n153 B 0.011026f
C271 VTAIL.n154 B 0.010414f
C272 VTAIL.n155 B 0.01938f
C273 VTAIL.n156 B 0.01938f
C274 VTAIL.n157 B 0.010414f
C275 VTAIL.n158 B 0.011026f
C276 VTAIL.n159 B 0.024614f
C277 VTAIL.n160 B 0.055367f
C278 VTAIL.n161 B 0.011026f
C279 VTAIL.n162 B 0.010414f
C280 VTAIL.n163 B 0.042942f
C281 VTAIL.n164 B 0.031136f
C282 VTAIL.n165 B 0.230567f
C283 VTAIL.t9 B 0.228644f
C284 VTAIL.t6 B 0.228644f
C285 VTAIL.n166 B 1.99816f
C286 VTAIL.n167 B 0.571836f
C287 VTAIL.n168 B 0.028417f
C288 VTAIL.n169 B 0.01938f
C289 VTAIL.n170 B 0.010414f
C290 VTAIL.n171 B 0.024614f
C291 VTAIL.n172 B 0.011026f
C292 VTAIL.n173 B 0.01938f
C293 VTAIL.n174 B 0.010414f
C294 VTAIL.n175 B 0.024614f
C295 VTAIL.n176 B 0.011026f
C296 VTAIL.n177 B 0.01938f
C297 VTAIL.n178 B 0.010414f
C298 VTAIL.n179 B 0.024614f
C299 VTAIL.n180 B 0.011026f
C300 VTAIL.n181 B 0.01938f
C301 VTAIL.n182 B 0.010414f
C302 VTAIL.n183 B 0.024614f
C303 VTAIL.n184 B 0.011026f
C304 VTAIL.n185 B 0.01938f
C305 VTAIL.n186 B 0.010414f
C306 VTAIL.n187 B 0.024614f
C307 VTAIL.n188 B 0.011026f
C308 VTAIL.n189 B 0.01938f
C309 VTAIL.n190 B 0.010414f
C310 VTAIL.n191 B 0.024614f
C311 VTAIL.n192 B 0.011026f
C312 VTAIL.n193 B 0.161525f
C313 VTAIL.t7 B 0.041878f
C314 VTAIL.n194 B 0.018461f
C315 VTAIL.n195 B 0.0174f
C316 VTAIL.n196 B 0.010414f
C317 VTAIL.n197 B 1.23023f
C318 VTAIL.n198 B 0.01938f
C319 VTAIL.n199 B 0.010414f
C320 VTAIL.n200 B 0.011026f
C321 VTAIL.n201 B 0.024614f
C322 VTAIL.n202 B 0.024614f
C323 VTAIL.n203 B 0.011026f
C324 VTAIL.n204 B 0.010414f
C325 VTAIL.n205 B 0.01938f
C326 VTAIL.n206 B 0.01938f
C327 VTAIL.n207 B 0.010414f
C328 VTAIL.n208 B 0.011026f
C329 VTAIL.n209 B 0.024614f
C330 VTAIL.n210 B 0.024614f
C331 VTAIL.n211 B 0.024614f
C332 VTAIL.n212 B 0.011026f
C333 VTAIL.n213 B 0.010414f
C334 VTAIL.n214 B 0.01938f
C335 VTAIL.n215 B 0.01938f
C336 VTAIL.n216 B 0.010414f
C337 VTAIL.n217 B 0.01072f
C338 VTAIL.n218 B 0.01072f
C339 VTAIL.n219 B 0.024614f
C340 VTAIL.n220 B 0.024614f
C341 VTAIL.n221 B 0.011026f
C342 VTAIL.n222 B 0.010414f
C343 VTAIL.n223 B 0.01938f
C344 VTAIL.n224 B 0.01938f
C345 VTAIL.n225 B 0.010414f
C346 VTAIL.n226 B 0.011026f
C347 VTAIL.n227 B 0.024614f
C348 VTAIL.n228 B 0.024614f
C349 VTAIL.n229 B 0.011026f
C350 VTAIL.n230 B 0.010414f
C351 VTAIL.n231 B 0.01938f
C352 VTAIL.n232 B 0.01938f
C353 VTAIL.n233 B 0.010414f
C354 VTAIL.n234 B 0.011026f
C355 VTAIL.n235 B 0.024614f
C356 VTAIL.n236 B 0.024614f
C357 VTAIL.n237 B 0.011026f
C358 VTAIL.n238 B 0.010414f
C359 VTAIL.n239 B 0.01938f
C360 VTAIL.n240 B 0.01938f
C361 VTAIL.n241 B 0.010414f
C362 VTAIL.n242 B 0.011026f
C363 VTAIL.n243 B 0.024614f
C364 VTAIL.n244 B 0.055367f
C365 VTAIL.n245 B 0.011026f
C366 VTAIL.n246 B 0.010414f
C367 VTAIL.n247 B 0.042942f
C368 VTAIL.n248 B 0.031136f
C369 VTAIL.n249 B 1.45392f
C370 VTAIL.n250 B 0.028417f
C371 VTAIL.n251 B 0.01938f
C372 VTAIL.n252 B 0.010414f
C373 VTAIL.n253 B 0.024614f
C374 VTAIL.n254 B 0.011026f
C375 VTAIL.n255 B 0.01938f
C376 VTAIL.n256 B 0.010414f
C377 VTAIL.n257 B 0.024614f
C378 VTAIL.n258 B 0.011026f
C379 VTAIL.n259 B 0.01938f
C380 VTAIL.n260 B 0.010414f
C381 VTAIL.n261 B 0.024614f
C382 VTAIL.n262 B 0.011026f
C383 VTAIL.n263 B 0.01938f
C384 VTAIL.n264 B 0.010414f
C385 VTAIL.n265 B 0.024614f
C386 VTAIL.n266 B 0.011026f
C387 VTAIL.n267 B 0.01938f
C388 VTAIL.n268 B 0.010414f
C389 VTAIL.n269 B 0.024614f
C390 VTAIL.n270 B 0.024614f
C391 VTAIL.n271 B 0.011026f
C392 VTAIL.n272 B 0.01938f
C393 VTAIL.n273 B 0.010414f
C394 VTAIL.n274 B 0.024614f
C395 VTAIL.n275 B 0.011026f
C396 VTAIL.n276 B 0.161525f
C397 VTAIL.t2 B 0.041878f
C398 VTAIL.n277 B 0.018461f
C399 VTAIL.n278 B 0.0174f
C400 VTAIL.n279 B 0.010414f
C401 VTAIL.n280 B 1.23023f
C402 VTAIL.n281 B 0.01938f
C403 VTAIL.n282 B 0.010414f
C404 VTAIL.n283 B 0.011026f
C405 VTAIL.n284 B 0.024614f
C406 VTAIL.n285 B 0.024614f
C407 VTAIL.n286 B 0.011026f
C408 VTAIL.n287 B 0.010414f
C409 VTAIL.n288 B 0.01938f
C410 VTAIL.n289 B 0.01938f
C411 VTAIL.n290 B 0.010414f
C412 VTAIL.n291 B 0.011026f
C413 VTAIL.n292 B 0.024614f
C414 VTAIL.n293 B 0.024614f
C415 VTAIL.n294 B 0.011026f
C416 VTAIL.n295 B 0.010414f
C417 VTAIL.n296 B 0.01938f
C418 VTAIL.n297 B 0.01938f
C419 VTAIL.n298 B 0.010414f
C420 VTAIL.n299 B 0.01072f
C421 VTAIL.n300 B 0.01072f
C422 VTAIL.n301 B 0.024614f
C423 VTAIL.n302 B 0.024614f
C424 VTAIL.n303 B 0.011026f
C425 VTAIL.n304 B 0.010414f
C426 VTAIL.n305 B 0.01938f
C427 VTAIL.n306 B 0.01938f
C428 VTAIL.n307 B 0.010414f
C429 VTAIL.n308 B 0.011026f
C430 VTAIL.n309 B 0.024614f
C431 VTAIL.n310 B 0.024614f
C432 VTAIL.n311 B 0.011026f
C433 VTAIL.n312 B 0.010414f
C434 VTAIL.n313 B 0.01938f
C435 VTAIL.n314 B 0.01938f
C436 VTAIL.n315 B 0.010414f
C437 VTAIL.n316 B 0.011026f
C438 VTAIL.n317 B 0.024614f
C439 VTAIL.n318 B 0.024614f
C440 VTAIL.n319 B 0.011026f
C441 VTAIL.n320 B 0.010414f
C442 VTAIL.n321 B 0.01938f
C443 VTAIL.n322 B 0.01938f
C444 VTAIL.n323 B 0.010414f
C445 VTAIL.n324 B 0.011026f
C446 VTAIL.n325 B 0.024614f
C447 VTAIL.n326 B 0.055367f
C448 VTAIL.n327 B 0.011026f
C449 VTAIL.n328 B 0.010414f
C450 VTAIL.n329 B 0.042942f
C451 VTAIL.n330 B 0.031136f
C452 VTAIL.n331 B 1.45392f
C453 VTAIL.t4 B 0.228644f
C454 VTAIL.t1 B 0.228644f
C455 VTAIL.n332 B 1.99817f
C456 VTAIL.n333 B 0.571826f
C457 VTAIL.n334 B 0.028417f
C458 VTAIL.n335 B 0.01938f
C459 VTAIL.n336 B 0.010414f
C460 VTAIL.n337 B 0.024614f
C461 VTAIL.n338 B 0.011026f
C462 VTAIL.n339 B 0.01938f
C463 VTAIL.n340 B 0.010414f
C464 VTAIL.n341 B 0.024614f
C465 VTAIL.n342 B 0.011026f
C466 VTAIL.n343 B 0.01938f
C467 VTAIL.n344 B 0.010414f
C468 VTAIL.n345 B 0.024614f
C469 VTAIL.n346 B 0.011026f
C470 VTAIL.n347 B 0.01938f
C471 VTAIL.n348 B 0.010414f
C472 VTAIL.n349 B 0.024614f
C473 VTAIL.n350 B 0.011026f
C474 VTAIL.n351 B 0.01938f
C475 VTAIL.n352 B 0.010414f
C476 VTAIL.n353 B 0.024614f
C477 VTAIL.n354 B 0.024614f
C478 VTAIL.n355 B 0.011026f
C479 VTAIL.n356 B 0.01938f
C480 VTAIL.n357 B 0.010414f
C481 VTAIL.n358 B 0.024614f
C482 VTAIL.n359 B 0.011026f
C483 VTAIL.n360 B 0.161525f
C484 VTAIL.t14 B 0.041878f
C485 VTAIL.n361 B 0.018461f
C486 VTAIL.n362 B 0.0174f
C487 VTAIL.n363 B 0.010414f
C488 VTAIL.n364 B 1.23023f
C489 VTAIL.n365 B 0.01938f
C490 VTAIL.n366 B 0.010414f
C491 VTAIL.n367 B 0.011026f
C492 VTAIL.n368 B 0.024614f
C493 VTAIL.n369 B 0.024614f
C494 VTAIL.n370 B 0.011026f
C495 VTAIL.n371 B 0.010414f
C496 VTAIL.n372 B 0.01938f
C497 VTAIL.n373 B 0.01938f
C498 VTAIL.n374 B 0.010414f
C499 VTAIL.n375 B 0.011026f
C500 VTAIL.n376 B 0.024614f
C501 VTAIL.n377 B 0.024614f
C502 VTAIL.n378 B 0.011026f
C503 VTAIL.n379 B 0.010414f
C504 VTAIL.n380 B 0.01938f
C505 VTAIL.n381 B 0.01938f
C506 VTAIL.n382 B 0.010414f
C507 VTAIL.n383 B 0.01072f
C508 VTAIL.n384 B 0.01072f
C509 VTAIL.n385 B 0.024614f
C510 VTAIL.n386 B 0.024614f
C511 VTAIL.n387 B 0.011026f
C512 VTAIL.n388 B 0.010414f
C513 VTAIL.n389 B 0.01938f
C514 VTAIL.n390 B 0.01938f
C515 VTAIL.n391 B 0.010414f
C516 VTAIL.n392 B 0.011026f
C517 VTAIL.n393 B 0.024614f
C518 VTAIL.n394 B 0.024614f
C519 VTAIL.n395 B 0.011026f
C520 VTAIL.n396 B 0.010414f
C521 VTAIL.n397 B 0.01938f
C522 VTAIL.n398 B 0.01938f
C523 VTAIL.n399 B 0.010414f
C524 VTAIL.n400 B 0.011026f
C525 VTAIL.n401 B 0.024614f
C526 VTAIL.n402 B 0.024614f
C527 VTAIL.n403 B 0.011026f
C528 VTAIL.n404 B 0.010414f
C529 VTAIL.n405 B 0.01938f
C530 VTAIL.n406 B 0.01938f
C531 VTAIL.n407 B 0.010414f
C532 VTAIL.n408 B 0.011026f
C533 VTAIL.n409 B 0.024614f
C534 VTAIL.n410 B 0.055367f
C535 VTAIL.n411 B 0.011026f
C536 VTAIL.n412 B 0.010414f
C537 VTAIL.n413 B 0.042942f
C538 VTAIL.n414 B 0.031136f
C539 VTAIL.n415 B 0.230567f
C540 VTAIL.n416 B 0.028417f
C541 VTAIL.n417 B 0.01938f
C542 VTAIL.n418 B 0.010414f
C543 VTAIL.n419 B 0.024614f
C544 VTAIL.n420 B 0.011026f
C545 VTAIL.n421 B 0.01938f
C546 VTAIL.n422 B 0.010414f
C547 VTAIL.n423 B 0.024614f
C548 VTAIL.n424 B 0.011026f
C549 VTAIL.n425 B 0.01938f
C550 VTAIL.n426 B 0.010414f
C551 VTAIL.n427 B 0.024614f
C552 VTAIL.n428 B 0.011026f
C553 VTAIL.n429 B 0.01938f
C554 VTAIL.n430 B 0.010414f
C555 VTAIL.n431 B 0.024614f
C556 VTAIL.n432 B 0.011026f
C557 VTAIL.n433 B 0.01938f
C558 VTAIL.n434 B 0.010414f
C559 VTAIL.n435 B 0.024614f
C560 VTAIL.n436 B 0.024614f
C561 VTAIL.n437 B 0.011026f
C562 VTAIL.n438 B 0.01938f
C563 VTAIL.n439 B 0.010414f
C564 VTAIL.n440 B 0.024614f
C565 VTAIL.n441 B 0.011026f
C566 VTAIL.n442 B 0.161525f
C567 VTAIL.t8 B 0.041878f
C568 VTAIL.n443 B 0.018461f
C569 VTAIL.n444 B 0.0174f
C570 VTAIL.n445 B 0.010414f
C571 VTAIL.n446 B 1.23023f
C572 VTAIL.n447 B 0.01938f
C573 VTAIL.n448 B 0.010414f
C574 VTAIL.n449 B 0.011026f
C575 VTAIL.n450 B 0.024614f
C576 VTAIL.n451 B 0.024614f
C577 VTAIL.n452 B 0.011026f
C578 VTAIL.n453 B 0.010414f
C579 VTAIL.n454 B 0.01938f
C580 VTAIL.n455 B 0.01938f
C581 VTAIL.n456 B 0.010414f
C582 VTAIL.n457 B 0.011026f
C583 VTAIL.n458 B 0.024614f
C584 VTAIL.n459 B 0.024614f
C585 VTAIL.n460 B 0.011026f
C586 VTAIL.n461 B 0.010414f
C587 VTAIL.n462 B 0.01938f
C588 VTAIL.n463 B 0.01938f
C589 VTAIL.n464 B 0.010414f
C590 VTAIL.n465 B 0.01072f
C591 VTAIL.n466 B 0.01072f
C592 VTAIL.n467 B 0.024614f
C593 VTAIL.n468 B 0.024614f
C594 VTAIL.n469 B 0.011026f
C595 VTAIL.n470 B 0.010414f
C596 VTAIL.n471 B 0.01938f
C597 VTAIL.n472 B 0.01938f
C598 VTAIL.n473 B 0.010414f
C599 VTAIL.n474 B 0.011026f
C600 VTAIL.n475 B 0.024614f
C601 VTAIL.n476 B 0.024614f
C602 VTAIL.n477 B 0.011026f
C603 VTAIL.n478 B 0.010414f
C604 VTAIL.n479 B 0.01938f
C605 VTAIL.n480 B 0.01938f
C606 VTAIL.n481 B 0.010414f
C607 VTAIL.n482 B 0.011026f
C608 VTAIL.n483 B 0.024614f
C609 VTAIL.n484 B 0.024614f
C610 VTAIL.n485 B 0.011026f
C611 VTAIL.n486 B 0.010414f
C612 VTAIL.n487 B 0.01938f
C613 VTAIL.n488 B 0.01938f
C614 VTAIL.n489 B 0.010414f
C615 VTAIL.n490 B 0.011026f
C616 VTAIL.n491 B 0.024614f
C617 VTAIL.n492 B 0.055367f
C618 VTAIL.n493 B 0.011026f
C619 VTAIL.n494 B 0.010414f
C620 VTAIL.n495 B 0.042942f
C621 VTAIL.n496 B 0.031136f
C622 VTAIL.n497 B 0.230567f
C623 VTAIL.t13 B 0.228644f
C624 VTAIL.t12 B 0.228644f
C625 VTAIL.n498 B 1.99817f
C626 VTAIL.n499 B 0.571826f
C627 VTAIL.n500 B 0.028417f
C628 VTAIL.n501 B 0.01938f
C629 VTAIL.n502 B 0.010414f
C630 VTAIL.n503 B 0.024614f
C631 VTAIL.n504 B 0.011026f
C632 VTAIL.n505 B 0.01938f
C633 VTAIL.n506 B 0.010414f
C634 VTAIL.n507 B 0.024614f
C635 VTAIL.n508 B 0.011026f
C636 VTAIL.n509 B 0.01938f
C637 VTAIL.n510 B 0.010414f
C638 VTAIL.n511 B 0.024614f
C639 VTAIL.n512 B 0.011026f
C640 VTAIL.n513 B 0.01938f
C641 VTAIL.n514 B 0.010414f
C642 VTAIL.n515 B 0.024614f
C643 VTAIL.n516 B 0.011026f
C644 VTAIL.n517 B 0.01938f
C645 VTAIL.n518 B 0.010414f
C646 VTAIL.n519 B 0.024614f
C647 VTAIL.n520 B 0.024614f
C648 VTAIL.n521 B 0.011026f
C649 VTAIL.n522 B 0.01938f
C650 VTAIL.n523 B 0.010414f
C651 VTAIL.n524 B 0.024614f
C652 VTAIL.n525 B 0.011026f
C653 VTAIL.n526 B 0.161525f
C654 VTAIL.t10 B 0.041878f
C655 VTAIL.n527 B 0.018461f
C656 VTAIL.n528 B 0.0174f
C657 VTAIL.n529 B 0.010414f
C658 VTAIL.n530 B 1.23023f
C659 VTAIL.n531 B 0.01938f
C660 VTAIL.n532 B 0.010414f
C661 VTAIL.n533 B 0.011026f
C662 VTAIL.n534 B 0.024614f
C663 VTAIL.n535 B 0.024614f
C664 VTAIL.n536 B 0.011026f
C665 VTAIL.n537 B 0.010414f
C666 VTAIL.n538 B 0.01938f
C667 VTAIL.n539 B 0.01938f
C668 VTAIL.n540 B 0.010414f
C669 VTAIL.n541 B 0.011026f
C670 VTAIL.n542 B 0.024614f
C671 VTAIL.n543 B 0.024614f
C672 VTAIL.n544 B 0.011026f
C673 VTAIL.n545 B 0.010414f
C674 VTAIL.n546 B 0.01938f
C675 VTAIL.n547 B 0.01938f
C676 VTAIL.n548 B 0.010414f
C677 VTAIL.n549 B 0.01072f
C678 VTAIL.n550 B 0.01072f
C679 VTAIL.n551 B 0.024614f
C680 VTAIL.n552 B 0.024614f
C681 VTAIL.n553 B 0.011026f
C682 VTAIL.n554 B 0.010414f
C683 VTAIL.n555 B 0.01938f
C684 VTAIL.n556 B 0.01938f
C685 VTAIL.n557 B 0.010414f
C686 VTAIL.n558 B 0.011026f
C687 VTAIL.n559 B 0.024614f
C688 VTAIL.n560 B 0.024614f
C689 VTAIL.n561 B 0.011026f
C690 VTAIL.n562 B 0.010414f
C691 VTAIL.n563 B 0.01938f
C692 VTAIL.n564 B 0.01938f
C693 VTAIL.n565 B 0.010414f
C694 VTAIL.n566 B 0.011026f
C695 VTAIL.n567 B 0.024614f
C696 VTAIL.n568 B 0.024614f
C697 VTAIL.n569 B 0.011026f
C698 VTAIL.n570 B 0.010414f
C699 VTAIL.n571 B 0.01938f
C700 VTAIL.n572 B 0.01938f
C701 VTAIL.n573 B 0.010414f
C702 VTAIL.n574 B 0.011026f
C703 VTAIL.n575 B 0.024614f
C704 VTAIL.n576 B 0.055367f
C705 VTAIL.n577 B 0.011026f
C706 VTAIL.n578 B 0.010414f
C707 VTAIL.n579 B 0.042942f
C708 VTAIL.n580 B 0.031136f
C709 VTAIL.n581 B 1.45392f
C710 VTAIL.n582 B 0.028417f
C711 VTAIL.n583 B 0.01938f
C712 VTAIL.n584 B 0.010414f
C713 VTAIL.n585 B 0.024614f
C714 VTAIL.n586 B 0.011026f
C715 VTAIL.n587 B 0.01938f
C716 VTAIL.n588 B 0.010414f
C717 VTAIL.n589 B 0.024614f
C718 VTAIL.n590 B 0.011026f
C719 VTAIL.n591 B 0.01938f
C720 VTAIL.n592 B 0.010414f
C721 VTAIL.n593 B 0.024614f
C722 VTAIL.n594 B 0.011026f
C723 VTAIL.n595 B 0.01938f
C724 VTAIL.n596 B 0.010414f
C725 VTAIL.n597 B 0.024614f
C726 VTAIL.n598 B 0.011026f
C727 VTAIL.n599 B 0.01938f
C728 VTAIL.n600 B 0.010414f
C729 VTAIL.n601 B 0.024614f
C730 VTAIL.n602 B 0.011026f
C731 VTAIL.n603 B 0.01938f
C732 VTAIL.n604 B 0.010414f
C733 VTAIL.n605 B 0.024614f
C734 VTAIL.n606 B 0.011026f
C735 VTAIL.n607 B 0.161525f
C736 VTAIL.t0 B 0.041878f
C737 VTAIL.n608 B 0.018461f
C738 VTAIL.n609 B 0.0174f
C739 VTAIL.n610 B 0.010414f
C740 VTAIL.n611 B 1.23023f
C741 VTAIL.n612 B 0.01938f
C742 VTAIL.n613 B 0.010414f
C743 VTAIL.n614 B 0.011026f
C744 VTAIL.n615 B 0.024614f
C745 VTAIL.n616 B 0.024614f
C746 VTAIL.n617 B 0.011026f
C747 VTAIL.n618 B 0.010414f
C748 VTAIL.n619 B 0.01938f
C749 VTAIL.n620 B 0.01938f
C750 VTAIL.n621 B 0.010414f
C751 VTAIL.n622 B 0.011026f
C752 VTAIL.n623 B 0.024614f
C753 VTAIL.n624 B 0.024614f
C754 VTAIL.n625 B 0.024614f
C755 VTAIL.n626 B 0.011026f
C756 VTAIL.n627 B 0.010414f
C757 VTAIL.n628 B 0.01938f
C758 VTAIL.n629 B 0.01938f
C759 VTAIL.n630 B 0.010414f
C760 VTAIL.n631 B 0.01072f
C761 VTAIL.n632 B 0.01072f
C762 VTAIL.n633 B 0.024614f
C763 VTAIL.n634 B 0.024614f
C764 VTAIL.n635 B 0.011026f
C765 VTAIL.n636 B 0.010414f
C766 VTAIL.n637 B 0.01938f
C767 VTAIL.n638 B 0.01938f
C768 VTAIL.n639 B 0.010414f
C769 VTAIL.n640 B 0.011026f
C770 VTAIL.n641 B 0.024614f
C771 VTAIL.n642 B 0.024614f
C772 VTAIL.n643 B 0.011026f
C773 VTAIL.n644 B 0.010414f
C774 VTAIL.n645 B 0.01938f
C775 VTAIL.n646 B 0.01938f
C776 VTAIL.n647 B 0.010414f
C777 VTAIL.n648 B 0.011026f
C778 VTAIL.n649 B 0.024614f
C779 VTAIL.n650 B 0.024614f
C780 VTAIL.n651 B 0.011026f
C781 VTAIL.n652 B 0.010414f
C782 VTAIL.n653 B 0.01938f
C783 VTAIL.n654 B 0.01938f
C784 VTAIL.n655 B 0.010414f
C785 VTAIL.n656 B 0.011026f
C786 VTAIL.n657 B 0.024614f
C787 VTAIL.n658 B 0.055367f
C788 VTAIL.n659 B 0.011026f
C789 VTAIL.n660 B 0.010414f
C790 VTAIL.n661 B 0.042942f
C791 VTAIL.n662 B 0.031136f
C792 VTAIL.n663 B 1.45028f
C793 VP.t1 B 2.4719f
C794 VP.n0 B 0.940929f
C795 VP.n1 B 0.019368f
C796 VP.n2 B 0.025575f
C797 VP.n3 B 0.019368f
C798 VP.t5 B 2.4719f
C799 VP.n4 B 0.860602f
C800 VP.n5 B 0.019368f
C801 VP.n6 B 0.028274f
C802 VP.n7 B 0.019368f
C803 VP.t2 B 2.4719f
C804 VP.n8 B 0.036097f
C805 VP.n9 B 0.019368f
C806 VP.n10 B 0.036097f
C807 VP.t3 B 2.4719f
C808 VP.n11 B 0.940929f
C809 VP.n12 B 0.019368f
C810 VP.n13 B 0.025575f
C811 VP.n14 B 0.019368f
C812 VP.t6 B 2.4719f
C813 VP.n15 B 0.860602f
C814 VP.n16 B 0.019368f
C815 VP.n17 B 0.028274f
C816 VP.n18 B 0.220914f
C817 VP.t0 B 2.4719f
C818 VP.t7 B 2.69647f
C819 VP.n19 B 0.889271f
C820 VP.n20 B 0.932425f
C821 VP.n21 B 0.035205f
C822 VP.n22 B 0.036097f
C823 VP.n23 B 0.019368f
C824 VP.n24 B 0.019368f
C825 VP.n25 B 0.019368f
C826 VP.n26 B 0.028274f
C827 VP.n27 B 0.036097f
C828 VP.n28 B 0.035205f
C829 VP.n29 B 0.019368f
C830 VP.n30 B 0.019368f
C831 VP.n31 B 0.019166f
C832 VP.n32 B 0.036097f
C833 VP.n33 B 0.036097f
C834 VP.n34 B 0.019368f
C835 VP.n35 B 0.019368f
C836 VP.n36 B 0.019368f
C837 VP.n37 B 0.030972f
C838 VP.n38 B 0.036097f
C839 VP.n39 B 0.033423f
C840 VP.n40 B 0.031259f
C841 VP.n41 B 1.27657f
C842 VP.n42 B 1.28906f
C843 VP.t4 B 2.4719f
C844 VP.n43 B 0.940929f
C845 VP.n44 B 0.033423f
C846 VP.n45 B 0.031259f
C847 VP.n46 B 0.019368f
C848 VP.n47 B 0.019368f
C849 VP.n48 B 0.030972f
C850 VP.n49 B 0.025575f
C851 VP.n50 B 0.036097f
C852 VP.n51 B 0.019368f
C853 VP.n52 B 0.019368f
C854 VP.n53 B 0.019368f
C855 VP.n54 B 0.019166f
C856 VP.n55 B 0.860602f
C857 VP.n56 B 0.035205f
C858 VP.n57 B 0.036097f
C859 VP.n58 B 0.019368f
C860 VP.n59 B 0.019368f
C861 VP.n60 B 0.019368f
C862 VP.n61 B 0.028274f
C863 VP.n62 B 0.036097f
C864 VP.n63 B 0.035205f
C865 VP.n64 B 0.019368f
C866 VP.n65 B 0.019368f
C867 VP.n66 B 0.019166f
C868 VP.n67 B 0.036097f
C869 VP.n68 B 0.036097f
C870 VP.n69 B 0.019368f
C871 VP.n70 B 0.019368f
C872 VP.n71 B 0.019368f
C873 VP.n72 B 0.030972f
C874 VP.n73 B 0.036097f
C875 VP.n74 B 0.033423f
C876 VP.n75 B 0.031259f
C877 VP.n76 B 0.040327f
.ends

