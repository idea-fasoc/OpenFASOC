* NGSPICE file created from diff_pair_sample_1192.ext - technology: sky130A

.subckt diff_pair_sample_1192 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
X1 B.t11 B.t9 B.t10 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=0 ps=0 w=18.94 l=1.74
X2 VDD1.t7 VP.t0 VTAIL.t2 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=7.3866 ps=38.66 w=18.94 l=1.74
X3 B.t8 B.t6 B.t7 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=0 ps=0 w=18.94 l=1.74
X4 VDD2.t6 VN.t1 VTAIL.t10 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=7.3866 ps=38.66 w=18.94 l=1.74
X5 VTAIL.t13 VN.t2 VDD2.t5 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
X6 VDD1.t6 VP.t1 VTAIL.t3 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
X7 VTAIL.t1 VP.t2 VDD1.t5 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=3.1251 ps=19.27 w=18.94 l=1.74
X8 B.t5 B.t3 B.t4 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=0 ps=0 w=18.94 l=1.74
X9 VTAIL.t15 VN.t3 VDD2.t4 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=3.1251 ps=19.27 w=18.94 l=1.74
X10 VTAIL.t6 VP.t3 VDD1.t4 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
X11 VDD1.t3 VP.t4 VTAIL.t0 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
X12 VDD2.t3 VN.t4 VTAIL.t14 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=7.3866 ps=38.66 w=18.94 l=1.74
X13 VTAIL.t5 VP.t5 VDD1.t2 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
X14 B.t2 B.t0 B.t1 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=0 ps=0 w=18.94 l=1.74
X15 VDD1.t1 VP.t6 VTAIL.t7 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=7.3866 ps=38.66 w=18.94 l=1.74
X16 VTAIL.t8 VN.t5 VDD2.t2 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
X17 VTAIL.t11 VN.t6 VDD2.t1 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=3.1251 ps=19.27 w=18.94 l=1.74
X18 VTAIL.t4 VP.t7 VDD1.t0 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=7.3866 pd=38.66 as=3.1251 ps=19.27 w=18.94 l=1.74
X19 VDD2.t0 VN.t7 VTAIL.t12 w_n3040_n4756# sky130_fd_pr__pfet_01v8 ad=3.1251 pd=19.27 as=3.1251 ps=19.27 w=18.94 l=1.74
R0 VN.n5 VN.t6 292.762
R1 VN.n28 VN.t4 292.762
R2 VN.n6 VN.t0 262.33
R3 VN.n14 VN.t2 262.33
R4 VN.n21 VN.t1 262.33
R5 VN.n29 VN.t5 262.33
R6 VN.n37 VN.t7 262.33
R7 VN.n44 VN.t3 262.33
R8 VN.n22 VN.n21 180.531
R9 VN.n45 VN.n44 180.531
R10 VN.n43 VN.n23 161.3
R11 VN.n42 VN.n41 161.3
R12 VN.n40 VN.n24 161.3
R13 VN.n39 VN.n38 161.3
R14 VN.n36 VN.n25 161.3
R15 VN.n35 VN.n34 161.3
R16 VN.n33 VN.n26 161.3
R17 VN.n32 VN.n31 161.3
R18 VN.n30 VN.n27 161.3
R19 VN.n20 VN.n0 161.3
R20 VN.n19 VN.n18 161.3
R21 VN.n17 VN.n1 161.3
R22 VN.n16 VN.n15 161.3
R23 VN.n13 VN.n2 161.3
R24 VN.n12 VN.n11 161.3
R25 VN.n10 VN.n3 161.3
R26 VN.n9 VN.n8 161.3
R27 VN.n7 VN.n4 161.3
R28 VN.n6 VN.n5 66.2123
R29 VN.n29 VN.n28 66.2123
R30 VN VN.n45 52.4191
R31 VN.n19 VN.n1 47.2268
R32 VN.n42 VN.n24 47.2268
R33 VN.n8 VN.n3 40.4106
R34 VN.n12 VN.n3 40.4106
R35 VN.n31 VN.n26 40.4106
R36 VN.n35 VN.n26 40.4106
R37 VN.n15 VN.n1 33.5944
R38 VN.n38 VN.n24 33.5944
R39 VN.n8 VN.n7 24.3439
R40 VN.n13 VN.n12 24.3439
R41 VN.n20 VN.n19 24.3439
R42 VN.n31 VN.n30 24.3439
R43 VN.n36 VN.n35 24.3439
R44 VN.n43 VN.n42 24.3439
R45 VN.n15 VN.n14 22.6399
R46 VN.n38 VN.n37 22.6399
R47 VN.n28 VN.n27 18.4539
R48 VN.n5 VN.n4 18.4539
R49 VN.n21 VN.n20 5.11262
R50 VN.n44 VN.n43 5.11262
R51 VN.n7 VN.n6 1.70454
R52 VN.n14 VN.n13 1.70454
R53 VN.n30 VN.n29 1.70454
R54 VN.n37 VN.n36 1.70454
R55 VN.n45 VN.n23 0.189894
R56 VN.n41 VN.n23 0.189894
R57 VN.n41 VN.n40 0.189894
R58 VN.n40 VN.n39 0.189894
R59 VN.n39 VN.n25 0.189894
R60 VN.n34 VN.n25 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n32 0.189894
R63 VN.n32 VN.n27 0.189894
R64 VN.n9 VN.n4 0.189894
R65 VN.n10 VN.n9 0.189894
R66 VN.n11 VN.n10 0.189894
R67 VN.n11 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n18 VN.n17 0.189894
R71 VN.n18 VN.n0 0.189894
R72 VN.n22 VN.n0 0.189894
R73 VN VN.n22 0.0516364
R74 VTAIL.n850 VTAIL.n750 756.745
R75 VTAIL.n102 VTAIL.n2 756.745
R76 VTAIL.n208 VTAIL.n108 756.745
R77 VTAIL.n316 VTAIL.n216 756.745
R78 VTAIL.n744 VTAIL.n644 756.745
R79 VTAIL.n636 VTAIL.n536 756.745
R80 VTAIL.n530 VTAIL.n430 756.745
R81 VTAIL.n422 VTAIL.n322 756.745
R82 VTAIL.n785 VTAIL.n784 585
R83 VTAIL.n782 VTAIL.n781 585
R84 VTAIL.n791 VTAIL.n790 585
R85 VTAIL.n793 VTAIL.n792 585
R86 VTAIL.n778 VTAIL.n777 585
R87 VTAIL.n799 VTAIL.n798 585
R88 VTAIL.n801 VTAIL.n800 585
R89 VTAIL.n774 VTAIL.n773 585
R90 VTAIL.n807 VTAIL.n806 585
R91 VTAIL.n809 VTAIL.n808 585
R92 VTAIL.n770 VTAIL.n769 585
R93 VTAIL.n815 VTAIL.n814 585
R94 VTAIL.n817 VTAIL.n816 585
R95 VTAIL.n766 VTAIL.n765 585
R96 VTAIL.n823 VTAIL.n822 585
R97 VTAIL.n826 VTAIL.n825 585
R98 VTAIL.n824 VTAIL.n762 585
R99 VTAIL.n831 VTAIL.n761 585
R100 VTAIL.n833 VTAIL.n832 585
R101 VTAIL.n835 VTAIL.n834 585
R102 VTAIL.n758 VTAIL.n757 585
R103 VTAIL.n841 VTAIL.n840 585
R104 VTAIL.n843 VTAIL.n842 585
R105 VTAIL.n754 VTAIL.n753 585
R106 VTAIL.n849 VTAIL.n848 585
R107 VTAIL.n851 VTAIL.n850 585
R108 VTAIL.n37 VTAIL.n36 585
R109 VTAIL.n34 VTAIL.n33 585
R110 VTAIL.n43 VTAIL.n42 585
R111 VTAIL.n45 VTAIL.n44 585
R112 VTAIL.n30 VTAIL.n29 585
R113 VTAIL.n51 VTAIL.n50 585
R114 VTAIL.n53 VTAIL.n52 585
R115 VTAIL.n26 VTAIL.n25 585
R116 VTAIL.n59 VTAIL.n58 585
R117 VTAIL.n61 VTAIL.n60 585
R118 VTAIL.n22 VTAIL.n21 585
R119 VTAIL.n67 VTAIL.n66 585
R120 VTAIL.n69 VTAIL.n68 585
R121 VTAIL.n18 VTAIL.n17 585
R122 VTAIL.n75 VTAIL.n74 585
R123 VTAIL.n78 VTAIL.n77 585
R124 VTAIL.n76 VTAIL.n14 585
R125 VTAIL.n83 VTAIL.n13 585
R126 VTAIL.n85 VTAIL.n84 585
R127 VTAIL.n87 VTAIL.n86 585
R128 VTAIL.n10 VTAIL.n9 585
R129 VTAIL.n93 VTAIL.n92 585
R130 VTAIL.n95 VTAIL.n94 585
R131 VTAIL.n6 VTAIL.n5 585
R132 VTAIL.n101 VTAIL.n100 585
R133 VTAIL.n103 VTAIL.n102 585
R134 VTAIL.n143 VTAIL.n142 585
R135 VTAIL.n140 VTAIL.n139 585
R136 VTAIL.n149 VTAIL.n148 585
R137 VTAIL.n151 VTAIL.n150 585
R138 VTAIL.n136 VTAIL.n135 585
R139 VTAIL.n157 VTAIL.n156 585
R140 VTAIL.n159 VTAIL.n158 585
R141 VTAIL.n132 VTAIL.n131 585
R142 VTAIL.n165 VTAIL.n164 585
R143 VTAIL.n167 VTAIL.n166 585
R144 VTAIL.n128 VTAIL.n127 585
R145 VTAIL.n173 VTAIL.n172 585
R146 VTAIL.n175 VTAIL.n174 585
R147 VTAIL.n124 VTAIL.n123 585
R148 VTAIL.n181 VTAIL.n180 585
R149 VTAIL.n184 VTAIL.n183 585
R150 VTAIL.n182 VTAIL.n120 585
R151 VTAIL.n189 VTAIL.n119 585
R152 VTAIL.n191 VTAIL.n190 585
R153 VTAIL.n193 VTAIL.n192 585
R154 VTAIL.n116 VTAIL.n115 585
R155 VTAIL.n199 VTAIL.n198 585
R156 VTAIL.n201 VTAIL.n200 585
R157 VTAIL.n112 VTAIL.n111 585
R158 VTAIL.n207 VTAIL.n206 585
R159 VTAIL.n209 VTAIL.n208 585
R160 VTAIL.n251 VTAIL.n250 585
R161 VTAIL.n248 VTAIL.n247 585
R162 VTAIL.n257 VTAIL.n256 585
R163 VTAIL.n259 VTAIL.n258 585
R164 VTAIL.n244 VTAIL.n243 585
R165 VTAIL.n265 VTAIL.n264 585
R166 VTAIL.n267 VTAIL.n266 585
R167 VTAIL.n240 VTAIL.n239 585
R168 VTAIL.n273 VTAIL.n272 585
R169 VTAIL.n275 VTAIL.n274 585
R170 VTAIL.n236 VTAIL.n235 585
R171 VTAIL.n281 VTAIL.n280 585
R172 VTAIL.n283 VTAIL.n282 585
R173 VTAIL.n232 VTAIL.n231 585
R174 VTAIL.n289 VTAIL.n288 585
R175 VTAIL.n292 VTAIL.n291 585
R176 VTAIL.n290 VTAIL.n228 585
R177 VTAIL.n297 VTAIL.n227 585
R178 VTAIL.n299 VTAIL.n298 585
R179 VTAIL.n301 VTAIL.n300 585
R180 VTAIL.n224 VTAIL.n223 585
R181 VTAIL.n307 VTAIL.n306 585
R182 VTAIL.n309 VTAIL.n308 585
R183 VTAIL.n220 VTAIL.n219 585
R184 VTAIL.n315 VTAIL.n314 585
R185 VTAIL.n317 VTAIL.n316 585
R186 VTAIL.n745 VTAIL.n744 585
R187 VTAIL.n743 VTAIL.n742 585
R188 VTAIL.n648 VTAIL.n647 585
R189 VTAIL.n737 VTAIL.n736 585
R190 VTAIL.n735 VTAIL.n734 585
R191 VTAIL.n652 VTAIL.n651 585
R192 VTAIL.n729 VTAIL.n728 585
R193 VTAIL.n727 VTAIL.n726 585
R194 VTAIL.n725 VTAIL.n655 585
R195 VTAIL.n659 VTAIL.n656 585
R196 VTAIL.n720 VTAIL.n719 585
R197 VTAIL.n718 VTAIL.n717 585
R198 VTAIL.n661 VTAIL.n660 585
R199 VTAIL.n712 VTAIL.n711 585
R200 VTAIL.n710 VTAIL.n709 585
R201 VTAIL.n665 VTAIL.n664 585
R202 VTAIL.n704 VTAIL.n703 585
R203 VTAIL.n702 VTAIL.n701 585
R204 VTAIL.n669 VTAIL.n668 585
R205 VTAIL.n696 VTAIL.n695 585
R206 VTAIL.n694 VTAIL.n693 585
R207 VTAIL.n673 VTAIL.n672 585
R208 VTAIL.n688 VTAIL.n687 585
R209 VTAIL.n686 VTAIL.n685 585
R210 VTAIL.n677 VTAIL.n676 585
R211 VTAIL.n680 VTAIL.n679 585
R212 VTAIL.n637 VTAIL.n636 585
R213 VTAIL.n635 VTAIL.n634 585
R214 VTAIL.n540 VTAIL.n539 585
R215 VTAIL.n629 VTAIL.n628 585
R216 VTAIL.n627 VTAIL.n626 585
R217 VTAIL.n544 VTAIL.n543 585
R218 VTAIL.n621 VTAIL.n620 585
R219 VTAIL.n619 VTAIL.n618 585
R220 VTAIL.n617 VTAIL.n547 585
R221 VTAIL.n551 VTAIL.n548 585
R222 VTAIL.n612 VTAIL.n611 585
R223 VTAIL.n610 VTAIL.n609 585
R224 VTAIL.n553 VTAIL.n552 585
R225 VTAIL.n604 VTAIL.n603 585
R226 VTAIL.n602 VTAIL.n601 585
R227 VTAIL.n557 VTAIL.n556 585
R228 VTAIL.n596 VTAIL.n595 585
R229 VTAIL.n594 VTAIL.n593 585
R230 VTAIL.n561 VTAIL.n560 585
R231 VTAIL.n588 VTAIL.n587 585
R232 VTAIL.n586 VTAIL.n585 585
R233 VTAIL.n565 VTAIL.n564 585
R234 VTAIL.n580 VTAIL.n579 585
R235 VTAIL.n578 VTAIL.n577 585
R236 VTAIL.n569 VTAIL.n568 585
R237 VTAIL.n572 VTAIL.n571 585
R238 VTAIL.n531 VTAIL.n530 585
R239 VTAIL.n529 VTAIL.n528 585
R240 VTAIL.n434 VTAIL.n433 585
R241 VTAIL.n523 VTAIL.n522 585
R242 VTAIL.n521 VTAIL.n520 585
R243 VTAIL.n438 VTAIL.n437 585
R244 VTAIL.n515 VTAIL.n514 585
R245 VTAIL.n513 VTAIL.n512 585
R246 VTAIL.n511 VTAIL.n441 585
R247 VTAIL.n445 VTAIL.n442 585
R248 VTAIL.n506 VTAIL.n505 585
R249 VTAIL.n504 VTAIL.n503 585
R250 VTAIL.n447 VTAIL.n446 585
R251 VTAIL.n498 VTAIL.n497 585
R252 VTAIL.n496 VTAIL.n495 585
R253 VTAIL.n451 VTAIL.n450 585
R254 VTAIL.n490 VTAIL.n489 585
R255 VTAIL.n488 VTAIL.n487 585
R256 VTAIL.n455 VTAIL.n454 585
R257 VTAIL.n482 VTAIL.n481 585
R258 VTAIL.n480 VTAIL.n479 585
R259 VTAIL.n459 VTAIL.n458 585
R260 VTAIL.n474 VTAIL.n473 585
R261 VTAIL.n472 VTAIL.n471 585
R262 VTAIL.n463 VTAIL.n462 585
R263 VTAIL.n466 VTAIL.n465 585
R264 VTAIL.n423 VTAIL.n422 585
R265 VTAIL.n421 VTAIL.n420 585
R266 VTAIL.n326 VTAIL.n325 585
R267 VTAIL.n415 VTAIL.n414 585
R268 VTAIL.n413 VTAIL.n412 585
R269 VTAIL.n330 VTAIL.n329 585
R270 VTAIL.n407 VTAIL.n406 585
R271 VTAIL.n405 VTAIL.n404 585
R272 VTAIL.n403 VTAIL.n333 585
R273 VTAIL.n337 VTAIL.n334 585
R274 VTAIL.n398 VTAIL.n397 585
R275 VTAIL.n396 VTAIL.n395 585
R276 VTAIL.n339 VTAIL.n338 585
R277 VTAIL.n390 VTAIL.n389 585
R278 VTAIL.n388 VTAIL.n387 585
R279 VTAIL.n343 VTAIL.n342 585
R280 VTAIL.n382 VTAIL.n381 585
R281 VTAIL.n380 VTAIL.n379 585
R282 VTAIL.n347 VTAIL.n346 585
R283 VTAIL.n374 VTAIL.n373 585
R284 VTAIL.n372 VTAIL.n371 585
R285 VTAIL.n351 VTAIL.n350 585
R286 VTAIL.n366 VTAIL.n365 585
R287 VTAIL.n364 VTAIL.n363 585
R288 VTAIL.n355 VTAIL.n354 585
R289 VTAIL.n358 VTAIL.n357 585
R290 VTAIL.t7 VTAIL.n678 327.466
R291 VTAIL.t4 VTAIL.n570 327.466
R292 VTAIL.t14 VTAIL.n464 327.466
R293 VTAIL.t15 VTAIL.n356 327.466
R294 VTAIL.t10 VTAIL.n783 327.466
R295 VTAIL.t11 VTAIL.n35 327.466
R296 VTAIL.t2 VTAIL.n141 327.466
R297 VTAIL.t1 VTAIL.n249 327.466
R298 VTAIL.n784 VTAIL.n781 171.744
R299 VTAIL.n791 VTAIL.n781 171.744
R300 VTAIL.n792 VTAIL.n791 171.744
R301 VTAIL.n792 VTAIL.n777 171.744
R302 VTAIL.n799 VTAIL.n777 171.744
R303 VTAIL.n800 VTAIL.n799 171.744
R304 VTAIL.n800 VTAIL.n773 171.744
R305 VTAIL.n807 VTAIL.n773 171.744
R306 VTAIL.n808 VTAIL.n807 171.744
R307 VTAIL.n808 VTAIL.n769 171.744
R308 VTAIL.n815 VTAIL.n769 171.744
R309 VTAIL.n816 VTAIL.n815 171.744
R310 VTAIL.n816 VTAIL.n765 171.744
R311 VTAIL.n823 VTAIL.n765 171.744
R312 VTAIL.n825 VTAIL.n823 171.744
R313 VTAIL.n825 VTAIL.n824 171.744
R314 VTAIL.n824 VTAIL.n761 171.744
R315 VTAIL.n833 VTAIL.n761 171.744
R316 VTAIL.n834 VTAIL.n833 171.744
R317 VTAIL.n834 VTAIL.n757 171.744
R318 VTAIL.n841 VTAIL.n757 171.744
R319 VTAIL.n842 VTAIL.n841 171.744
R320 VTAIL.n842 VTAIL.n753 171.744
R321 VTAIL.n849 VTAIL.n753 171.744
R322 VTAIL.n850 VTAIL.n849 171.744
R323 VTAIL.n36 VTAIL.n33 171.744
R324 VTAIL.n43 VTAIL.n33 171.744
R325 VTAIL.n44 VTAIL.n43 171.744
R326 VTAIL.n44 VTAIL.n29 171.744
R327 VTAIL.n51 VTAIL.n29 171.744
R328 VTAIL.n52 VTAIL.n51 171.744
R329 VTAIL.n52 VTAIL.n25 171.744
R330 VTAIL.n59 VTAIL.n25 171.744
R331 VTAIL.n60 VTAIL.n59 171.744
R332 VTAIL.n60 VTAIL.n21 171.744
R333 VTAIL.n67 VTAIL.n21 171.744
R334 VTAIL.n68 VTAIL.n67 171.744
R335 VTAIL.n68 VTAIL.n17 171.744
R336 VTAIL.n75 VTAIL.n17 171.744
R337 VTAIL.n77 VTAIL.n75 171.744
R338 VTAIL.n77 VTAIL.n76 171.744
R339 VTAIL.n76 VTAIL.n13 171.744
R340 VTAIL.n85 VTAIL.n13 171.744
R341 VTAIL.n86 VTAIL.n85 171.744
R342 VTAIL.n86 VTAIL.n9 171.744
R343 VTAIL.n93 VTAIL.n9 171.744
R344 VTAIL.n94 VTAIL.n93 171.744
R345 VTAIL.n94 VTAIL.n5 171.744
R346 VTAIL.n101 VTAIL.n5 171.744
R347 VTAIL.n102 VTAIL.n101 171.744
R348 VTAIL.n142 VTAIL.n139 171.744
R349 VTAIL.n149 VTAIL.n139 171.744
R350 VTAIL.n150 VTAIL.n149 171.744
R351 VTAIL.n150 VTAIL.n135 171.744
R352 VTAIL.n157 VTAIL.n135 171.744
R353 VTAIL.n158 VTAIL.n157 171.744
R354 VTAIL.n158 VTAIL.n131 171.744
R355 VTAIL.n165 VTAIL.n131 171.744
R356 VTAIL.n166 VTAIL.n165 171.744
R357 VTAIL.n166 VTAIL.n127 171.744
R358 VTAIL.n173 VTAIL.n127 171.744
R359 VTAIL.n174 VTAIL.n173 171.744
R360 VTAIL.n174 VTAIL.n123 171.744
R361 VTAIL.n181 VTAIL.n123 171.744
R362 VTAIL.n183 VTAIL.n181 171.744
R363 VTAIL.n183 VTAIL.n182 171.744
R364 VTAIL.n182 VTAIL.n119 171.744
R365 VTAIL.n191 VTAIL.n119 171.744
R366 VTAIL.n192 VTAIL.n191 171.744
R367 VTAIL.n192 VTAIL.n115 171.744
R368 VTAIL.n199 VTAIL.n115 171.744
R369 VTAIL.n200 VTAIL.n199 171.744
R370 VTAIL.n200 VTAIL.n111 171.744
R371 VTAIL.n207 VTAIL.n111 171.744
R372 VTAIL.n208 VTAIL.n207 171.744
R373 VTAIL.n250 VTAIL.n247 171.744
R374 VTAIL.n257 VTAIL.n247 171.744
R375 VTAIL.n258 VTAIL.n257 171.744
R376 VTAIL.n258 VTAIL.n243 171.744
R377 VTAIL.n265 VTAIL.n243 171.744
R378 VTAIL.n266 VTAIL.n265 171.744
R379 VTAIL.n266 VTAIL.n239 171.744
R380 VTAIL.n273 VTAIL.n239 171.744
R381 VTAIL.n274 VTAIL.n273 171.744
R382 VTAIL.n274 VTAIL.n235 171.744
R383 VTAIL.n281 VTAIL.n235 171.744
R384 VTAIL.n282 VTAIL.n281 171.744
R385 VTAIL.n282 VTAIL.n231 171.744
R386 VTAIL.n289 VTAIL.n231 171.744
R387 VTAIL.n291 VTAIL.n289 171.744
R388 VTAIL.n291 VTAIL.n290 171.744
R389 VTAIL.n290 VTAIL.n227 171.744
R390 VTAIL.n299 VTAIL.n227 171.744
R391 VTAIL.n300 VTAIL.n299 171.744
R392 VTAIL.n300 VTAIL.n223 171.744
R393 VTAIL.n307 VTAIL.n223 171.744
R394 VTAIL.n308 VTAIL.n307 171.744
R395 VTAIL.n308 VTAIL.n219 171.744
R396 VTAIL.n315 VTAIL.n219 171.744
R397 VTAIL.n316 VTAIL.n315 171.744
R398 VTAIL.n744 VTAIL.n743 171.744
R399 VTAIL.n743 VTAIL.n647 171.744
R400 VTAIL.n736 VTAIL.n647 171.744
R401 VTAIL.n736 VTAIL.n735 171.744
R402 VTAIL.n735 VTAIL.n651 171.744
R403 VTAIL.n728 VTAIL.n651 171.744
R404 VTAIL.n728 VTAIL.n727 171.744
R405 VTAIL.n727 VTAIL.n655 171.744
R406 VTAIL.n659 VTAIL.n655 171.744
R407 VTAIL.n719 VTAIL.n659 171.744
R408 VTAIL.n719 VTAIL.n718 171.744
R409 VTAIL.n718 VTAIL.n660 171.744
R410 VTAIL.n711 VTAIL.n660 171.744
R411 VTAIL.n711 VTAIL.n710 171.744
R412 VTAIL.n710 VTAIL.n664 171.744
R413 VTAIL.n703 VTAIL.n664 171.744
R414 VTAIL.n703 VTAIL.n702 171.744
R415 VTAIL.n702 VTAIL.n668 171.744
R416 VTAIL.n695 VTAIL.n668 171.744
R417 VTAIL.n695 VTAIL.n694 171.744
R418 VTAIL.n694 VTAIL.n672 171.744
R419 VTAIL.n687 VTAIL.n672 171.744
R420 VTAIL.n687 VTAIL.n686 171.744
R421 VTAIL.n686 VTAIL.n676 171.744
R422 VTAIL.n679 VTAIL.n676 171.744
R423 VTAIL.n636 VTAIL.n635 171.744
R424 VTAIL.n635 VTAIL.n539 171.744
R425 VTAIL.n628 VTAIL.n539 171.744
R426 VTAIL.n628 VTAIL.n627 171.744
R427 VTAIL.n627 VTAIL.n543 171.744
R428 VTAIL.n620 VTAIL.n543 171.744
R429 VTAIL.n620 VTAIL.n619 171.744
R430 VTAIL.n619 VTAIL.n547 171.744
R431 VTAIL.n551 VTAIL.n547 171.744
R432 VTAIL.n611 VTAIL.n551 171.744
R433 VTAIL.n611 VTAIL.n610 171.744
R434 VTAIL.n610 VTAIL.n552 171.744
R435 VTAIL.n603 VTAIL.n552 171.744
R436 VTAIL.n603 VTAIL.n602 171.744
R437 VTAIL.n602 VTAIL.n556 171.744
R438 VTAIL.n595 VTAIL.n556 171.744
R439 VTAIL.n595 VTAIL.n594 171.744
R440 VTAIL.n594 VTAIL.n560 171.744
R441 VTAIL.n587 VTAIL.n560 171.744
R442 VTAIL.n587 VTAIL.n586 171.744
R443 VTAIL.n586 VTAIL.n564 171.744
R444 VTAIL.n579 VTAIL.n564 171.744
R445 VTAIL.n579 VTAIL.n578 171.744
R446 VTAIL.n578 VTAIL.n568 171.744
R447 VTAIL.n571 VTAIL.n568 171.744
R448 VTAIL.n530 VTAIL.n529 171.744
R449 VTAIL.n529 VTAIL.n433 171.744
R450 VTAIL.n522 VTAIL.n433 171.744
R451 VTAIL.n522 VTAIL.n521 171.744
R452 VTAIL.n521 VTAIL.n437 171.744
R453 VTAIL.n514 VTAIL.n437 171.744
R454 VTAIL.n514 VTAIL.n513 171.744
R455 VTAIL.n513 VTAIL.n441 171.744
R456 VTAIL.n445 VTAIL.n441 171.744
R457 VTAIL.n505 VTAIL.n445 171.744
R458 VTAIL.n505 VTAIL.n504 171.744
R459 VTAIL.n504 VTAIL.n446 171.744
R460 VTAIL.n497 VTAIL.n446 171.744
R461 VTAIL.n497 VTAIL.n496 171.744
R462 VTAIL.n496 VTAIL.n450 171.744
R463 VTAIL.n489 VTAIL.n450 171.744
R464 VTAIL.n489 VTAIL.n488 171.744
R465 VTAIL.n488 VTAIL.n454 171.744
R466 VTAIL.n481 VTAIL.n454 171.744
R467 VTAIL.n481 VTAIL.n480 171.744
R468 VTAIL.n480 VTAIL.n458 171.744
R469 VTAIL.n473 VTAIL.n458 171.744
R470 VTAIL.n473 VTAIL.n472 171.744
R471 VTAIL.n472 VTAIL.n462 171.744
R472 VTAIL.n465 VTAIL.n462 171.744
R473 VTAIL.n422 VTAIL.n421 171.744
R474 VTAIL.n421 VTAIL.n325 171.744
R475 VTAIL.n414 VTAIL.n325 171.744
R476 VTAIL.n414 VTAIL.n413 171.744
R477 VTAIL.n413 VTAIL.n329 171.744
R478 VTAIL.n406 VTAIL.n329 171.744
R479 VTAIL.n406 VTAIL.n405 171.744
R480 VTAIL.n405 VTAIL.n333 171.744
R481 VTAIL.n337 VTAIL.n333 171.744
R482 VTAIL.n397 VTAIL.n337 171.744
R483 VTAIL.n397 VTAIL.n396 171.744
R484 VTAIL.n396 VTAIL.n338 171.744
R485 VTAIL.n389 VTAIL.n338 171.744
R486 VTAIL.n389 VTAIL.n388 171.744
R487 VTAIL.n388 VTAIL.n342 171.744
R488 VTAIL.n381 VTAIL.n342 171.744
R489 VTAIL.n381 VTAIL.n380 171.744
R490 VTAIL.n380 VTAIL.n346 171.744
R491 VTAIL.n373 VTAIL.n346 171.744
R492 VTAIL.n373 VTAIL.n372 171.744
R493 VTAIL.n372 VTAIL.n350 171.744
R494 VTAIL.n365 VTAIL.n350 171.744
R495 VTAIL.n365 VTAIL.n364 171.744
R496 VTAIL.n364 VTAIL.n354 171.744
R497 VTAIL.n357 VTAIL.n354 171.744
R498 VTAIL.n784 VTAIL.t10 85.8723
R499 VTAIL.n36 VTAIL.t11 85.8723
R500 VTAIL.n142 VTAIL.t2 85.8723
R501 VTAIL.n250 VTAIL.t1 85.8723
R502 VTAIL.n679 VTAIL.t7 85.8723
R503 VTAIL.n571 VTAIL.t4 85.8723
R504 VTAIL.n465 VTAIL.t14 85.8723
R505 VTAIL.n357 VTAIL.t15 85.8723
R506 VTAIL.n1 VTAIL.n0 51.3183
R507 VTAIL.n215 VTAIL.n214 51.3183
R508 VTAIL.n643 VTAIL.n642 51.3182
R509 VTAIL.n429 VTAIL.n428 51.3182
R510 VTAIL.n855 VTAIL.n854 31.7975
R511 VTAIL.n107 VTAIL.n106 31.7975
R512 VTAIL.n213 VTAIL.n212 31.7975
R513 VTAIL.n321 VTAIL.n320 31.7975
R514 VTAIL.n749 VTAIL.n748 31.7975
R515 VTAIL.n641 VTAIL.n640 31.7975
R516 VTAIL.n535 VTAIL.n534 31.7975
R517 VTAIL.n427 VTAIL.n426 31.7975
R518 VTAIL.n855 VTAIL.n749 30.4789
R519 VTAIL.n427 VTAIL.n321 30.4789
R520 VTAIL.n785 VTAIL.n783 16.3895
R521 VTAIL.n37 VTAIL.n35 16.3895
R522 VTAIL.n143 VTAIL.n141 16.3895
R523 VTAIL.n251 VTAIL.n249 16.3895
R524 VTAIL.n680 VTAIL.n678 16.3895
R525 VTAIL.n572 VTAIL.n570 16.3895
R526 VTAIL.n466 VTAIL.n464 16.3895
R527 VTAIL.n358 VTAIL.n356 16.3895
R528 VTAIL.n832 VTAIL.n831 13.1884
R529 VTAIL.n84 VTAIL.n83 13.1884
R530 VTAIL.n190 VTAIL.n189 13.1884
R531 VTAIL.n298 VTAIL.n297 13.1884
R532 VTAIL.n726 VTAIL.n725 13.1884
R533 VTAIL.n618 VTAIL.n617 13.1884
R534 VTAIL.n512 VTAIL.n511 13.1884
R535 VTAIL.n404 VTAIL.n403 13.1884
R536 VTAIL.n786 VTAIL.n782 12.8005
R537 VTAIL.n830 VTAIL.n762 12.8005
R538 VTAIL.n835 VTAIL.n760 12.8005
R539 VTAIL.n38 VTAIL.n34 12.8005
R540 VTAIL.n82 VTAIL.n14 12.8005
R541 VTAIL.n87 VTAIL.n12 12.8005
R542 VTAIL.n144 VTAIL.n140 12.8005
R543 VTAIL.n188 VTAIL.n120 12.8005
R544 VTAIL.n193 VTAIL.n118 12.8005
R545 VTAIL.n252 VTAIL.n248 12.8005
R546 VTAIL.n296 VTAIL.n228 12.8005
R547 VTAIL.n301 VTAIL.n226 12.8005
R548 VTAIL.n729 VTAIL.n654 12.8005
R549 VTAIL.n724 VTAIL.n656 12.8005
R550 VTAIL.n681 VTAIL.n677 12.8005
R551 VTAIL.n621 VTAIL.n546 12.8005
R552 VTAIL.n616 VTAIL.n548 12.8005
R553 VTAIL.n573 VTAIL.n569 12.8005
R554 VTAIL.n515 VTAIL.n440 12.8005
R555 VTAIL.n510 VTAIL.n442 12.8005
R556 VTAIL.n467 VTAIL.n463 12.8005
R557 VTAIL.n407 VTAIL.n332 12.8005
R558 VTAIL.n402 VTAIL.n334 12.8005
R559 VTAIL.n359 VTAIL.n355 12.8005
R560 VTAIL.n790 VTAIL.n789 12.0247
R561 VTAIL.n827 VTAIL.n826 12.0247
R562 VTAIL.n836 VTAIL.n758 12.0247
R563 VTAIL.n42 VTAIL.n41 12.0247
R564 VTAIL.n79 VTAIL.n78 12.0247
R565 VTAIL.n88 VTAIL.n10 12.0247
R566 VTAIL.n148 VTAIL.n147 12.0247
R567 VTAIL.n185 VTAIL.n184 12.0247
R568 VTAIL.n194 VTAIL.n116 12.0247
R569 VTAIL.n256 VTAIL.n255 12.0247
R570 VTAIL.n293 VTAIL.n292 12.0247
R571 VTAIL.n302 VTAIL.n224 12.0247
R572 VTAIL.n730 VTAIL.n652 12.0247
R573 VTAIL.n721 VTAIL.n720 12.0247
R574 VTAIL.n685 VTAIL.n684 12.0247
R575 VTAIL.n622 VTAIL.n544 12.0247
R576 VTAIL.n613 VTAIL.n612 12.0247
R577 VTAIL.n577 VTAIL.n576 12.0247
R578 VTAIL.n516 VTAIL.n438 12.0247
R579 VTAIL.n507 VTAIL.n506 12.0247
R580 VTAIL.n471 VTAIL.n470 12.0247
R581 VTAIL.n408 VTAIL.n330 12.0247
R582 VTAIL.n399 VTAIL.n398 12.0247
R583 VTAIL.n363 VTAIL.n362 12.0247
R584 VTAIL.n793 VTAIL.n780 11.249
R585 VTAIL.n822 VTAIL.n764 11.249
R586 VTAIL.n840 VTAIL.n839 11.249
R587 VTAIL.n45 VTAIL.n32 11.249
R588 VTAIL.n74 VTAIL.n16 11.249
R589 VTAIL.n92 VTAIL.n91 11.249
R590 VTAIL.n151 VTAIL.n138 11.249
R591 VTAIL.n180 VTAIL.n122 11.249
R592 VTAIL.n198 VTAIL.n197 11.249
R593 VTAIL.n259 VTAIL.n246 11.249
R594 VTAIL.n288 VTAIL.n230 11.249
R595 VTAIL.n306 VTAIL.n305 11.249
R596 VTAIL.n734 VTAIL.n733 11.249
R597 VTAIL.n717 VTAIL.n658 11.249
R598 VTAIL.n688 VTAIL.n675 11.249
R599 VTAIL.n626 VTAIL.n625 11.249
R600 VTAIL.n609 VTAIL.n550 11.249
R601 VTAIL.n580 VTAIL.n567 11.249
R602 VTAIL.n520 VTAIL.n519 11.249
R603 VTAIL.n503 VTAIL.n444 11.249
R604 VTAIL.n474 VTAIL.n461 11.249
R605 VTAIL.n412 VTAIL.n411 11.249
R606 VTAIL.n395 VTAIL.n336 11.249
R607 VTAIL.n366 VTAIL.n353 11.249
R608 VTAIL.n794 VTAIL.n778 10.4732
R609 VTAIL.n821 VTAIL.n766 10.4732
R610 VTAIL.n843 VTAIL.n756 10.4732
R611 VTAIL.n46 VTAIL.n30 10.4732
R612 VTAIL.n73 VTAIL.n18 10.4732
R613 VTAIL.n95 VTAIL.n8 10.4732
R614 VTAIL.n152 VTAIL.n136 10.4732
R615 VTAIL.n179 VTAIL.n124 10.4732
R616 VTAIL.n201 VTAIL.n114 10.4732
R617 VTAIL.n260 VTAIL.n244 10.4732
R618 VTAIL.n287 VTAIL.n232 10.4732
R619 VTAIL.n309 VTAIL.n222 10.4732
R620 VTAIL.n737 VTAIL.n650 10.4732
R621 VTAIL.n716 VTAIL.n661 10.4732
R622 VTAIL.n689 VTAIL.n673 10.4732
R623 VTAIL.n629 VTAIL.n542 10.4732
R624 VTAIL.n608 VTAIL.n553 10.4732
R625 VTAIL.n581 VTAIL.n565 10.4732
R626 VTAIL.n523 VTAIL.n436 10.4732
R627 VTAIL.n502 VTAIL.n447 10.4732
R628 VTAIL.n475 VTAIL.n459 10.4732
R629 VTAIL.n415 VTAIL.n328 10.4732
R630 VTAIL.n394 VTAIL.n339 10.4732
R631 VTAIL.n367 VTAIL.n351 10.4732
R632 VTAIL.n798 VTAIL.n797 9.69747
R633 VTAIL.n818 VTAIL.n817 9.69747
R634 VTAIL.n844 VTAIL.n754 9.69747
R635 VTAIL.n50 VTAIL.n49 9.69747
R636 VTAIL.n70 VTAIL.n69 9.69747
R637 VTAIL.n96 VTAIL.n6 9.69747
R638 VTAIL.n156 VTAIL.n155 9.69747
R639 VTAIL.n176 VTAIL.n175 9.69747
R640 VTAIL.n202 VTAIL.n112 9.69747
R641 VTAIL.n264 VTAIL.n263 9.69747
R642 VTAIL.n284 VTAIL.n283 9.69747
R643 VTAIL.n310 VTAIL.n220 9.69747
R644 VTAIL.n738 VTAIL.n648 9.69747
R645 VTAIL.n713 VTAIL.n712 9.69747
R646 VTAIL.n693 VTAIL.n692 9.69747
R647 VTAIL.n630 VTAIL.n540 9.69747
R648 VTAIL.n605 VTAIL.n604 9.69747
R649 VTAIL.n585 VTAIL.n584 9.69747
R650 VTAIL.n524 VTAIL.n434 9.69747
R651 VTAIL.n499 VTAIL.n498 9.69747
R652 VTAIL.n479 VTAIL.n478 9.69747
R653 VTAIL.n416 VTAIL.n326 9.69747
R654 VTAIL.n391 VTAIL.n390 9.69747
R655 VTAIL.n371 VTAIL.n370 9.69747
R656 VTAIL.n854 VTAIL.n853 9.45567
R657 VTAIL.n106 VTAIL.n105 9.45567
R658 VTAIL.n212 VTAIL.n211 9.45567
R659 VTAIL.n320 VTAIL.n319 9.45567
R660 VTAIL.n748 VTAIL.n747 9.45567
R661 VTAIL.n640 VTAIL.n639 9.45567
R662 VTAIL.n534 VTAIL.n533 9.45567
R663 VTAIL.n426 VTAIL.n425 9.45567
R664 VTAIL.n752 VTAIL.n751 9.3005
R665 VTAIL.n847 VTAIL.n846 9.3005
R666 VTAIL.n845 VTAIL.n844 9.3005
R667 VTAIL.n756 VTAIL.n755 9.3005
R668 VTAIL.n839 VTAIL.n838 9.3005
R669 VTAIL.n837 VTAIL.n836 9.3005
R670 VTAIL.n760 VTAIL.n759 9.3005
R671 VTAIL.n805 VTAIL.n804 9.3005
R672 VTAIL.n803 VTAIL.n802 9.3005
R673 VTAIL.n776 VTAIL.n775 9.3005
R674 VTAIL.n797 VTAIL.n796 9.3005
R675 VTAIL.n795 VTAIL.n794 9.3005
R676 VTAIL.n780 VTAIL.n779 9.3005
R677 VTAIL.n789 VTAIL.n788 9.3005
R678 VTAIL.n787 VTAIL.n786 9.3005
R679 VTAIL.n772 VTAIL.n771 9.3005
R680 VTAIL.n811 VTAIL.n810 9.3005
R681 VTAIL.n813 VTAIL.n812 9.3005
R682 VTAIL.n768 VTAIL.n767 9.3005
R683 VTAIL.n819 VTAIL.n818 9.3005
R684 VTAIL.n821 VTAIL.n820 9.3005
R685 VTAIL.n764 VTAIL.n763 9.3005
R686 VTAIL.n828 VTAIL.n827 9.3005
R687 VTAIL.n830 VTAIL.n829 9.3005
R688 VTAIL.n853 VTAIL.n852 9.3005
R689 VTAIL.n4 VTAIL.n3 9.3005
R690 VTAIL.n99 VTAIL.n98 9.3005
R691 VTAIL.n97 VTAIL.n96 9.3005
R692 VTAIL.n8 VTAIL.n7 9.3005
R693 VTAIL.n91 VTAIL.n90 9.3005
R694 VTAIL.n89 VTAIL.n88 9.3005
R695 VTAIL.n12 VTAIL.n11 9.3005
R696 VTAIL.n57 VTAIL.n56 9.3005
R697 VTAIL.n55 VTAIL.n54 9.3005
R698 VTAIL.n28 VTAIL.n27 9.3005
R699 VTAIL.n49 VTAIL.n48 9.3005
R700 VTAIL.n47 VTAIL.n46 9.3005
R701 VTAIL.n32 VTAIL.n31 9.3005
R702 VTAIL.n41 VTAIL.n40 9.3005
R703 VTAIL.n39 VTAIL.n38 9.3005
R704 VTAIL.n24 VTAIL.n23 9.3005
R705 VTAIL.n63 VTAIL.n62 9.3005
R706 VTAIL.n65 VTAIL.n64 9.3005
R707 VTAIL.n20 VTAIL.n19 9.3005
R708 VTAIL.n71 VTAIL.n70 9.3005
R709 VTAIL.n73 VTAIL.n72 9.3005
R710 VTAIL.n16 VTAIL.n15 9.3005
R711 VTAIL.n80 VTAIL.n79 9.3005
R712 VTAIL.n82 VTAIL.n81 9.3005
R713 VTAIL.n105 VTAIL.n104 9.3005
R714 VTAIL.n110 VTAIL.n109 9.3005
R715 VTAIL.n205 VTAIL.n204 9.3005
R716 VTAIL.n203 VTAIL.n202 9.3005
R717 VTAIL.n114 VTAIL.n113 9.3005
R718 VTAIL.n197 VTAIL.n196 9.3005
R719 VTAIL.n195 VTAIL.n194 9.3005
R720 VTAIL.n118 VTAIL.n117 9.3005
R721 VTAIL.n163 VTAIL.n162 9.3005
R722 VTAIL.n161 VTAIL.n160 9.3005
R723 VTAIL.n134 VTAIL.n133 9.3005
R724 VTAIL.n155 VTAIL.n154 9.3005
R725 VTAIL.n153 VTAIL.n152 9.3005
R726 VTAIL.n138 VTAIL.n137 9.3005
R727 VTAIL.n147 VTAIL.n146 9.3005
R728 VTAIL.n145 VTAIL.n144 9.3005
R729 VTAIL.n130 VTAIL.n129 9.3005
R730 VTAIL.n169 VTAIL.n168 9.3005
R731 VTAIL.n171 VTAIL.n170 9.3005
R732 VTAIL.n126 VTAIL.n125 9.3005
R733 VTAIL.n177 VTAIL.n176 9.3005
R734 VTAIL.n179 VTAIL.n178 9.3005
R735 VTAIL.n122 VTAIL.n121 9.3005
R736 VTAIL.n186 VTAIL.n185 9.3005
R737 VTAIL.n188 VTAIL.n187 9.3005
R738 VTAIL.n211 VTAIL.n210 9.3005
R739 VTAIL.n218 VTAIL.n217 9.3005
R740 VTAIL.n313 VTAIL.n312 9.3005
R741 VTAIL.n311 VTAIL.n310 9.3005
R742 VTAIL.n222 VTAIL.n221 9.3005
R743 VTAIL.n305 VTAIL.n304 9.3005
R744 VTAIL.n303 VTAIL.n302 9.3005
R745 VTAIL.n226 VTAIL.n225 9.3005
R746 VTAIL.n271 VTAIL.n270 9.3005
R747 VTAIL.n269 VTAIL.n268 9.3005
R748 VTAIL.n242 VTAIL.n241 9.3005
R749 VTAIL.n263 VTAIL.n262 9.3005
R750 VTAIL.n261 VTAIL.n260 9.3005
R751 VTAIL.n246 VTAIL.n245 9.3005
R752 VTAIL.n255 VTAIL.n254 9.3005
R753 VTAIL.n253 VTAIL.n252 9.3005
R754 VTAIL.n238 VTAIL.n237 9.3005
R755 VTAIL.n277 VTAIL.n276 9.3005
R756 VTAIL.n279 VTAIL.n278 9.3005
R757 VTAIL.n234 VTAIL.n233 9.3005
R758 VTAIL.n285 VTAIL.n284 9.3005
R759 VTAIL.n287 VTAIL.n286 9.3005
R760 VTAIL.n230 VTAIL.n229 9.3005
R761 VTAIL.n294 VTAIL.n293 9.3005
R762 VTAIL.n296 VTAIL.n295 9.3005
R763 VTAIL.n319 VTAIL.n318 9.3005
R764 VTAIL.n706 VTAIL.n705 9.3005
R765 VTAIL.n708 VTAIL.n707 9.3005
R766 VTAIL.n663 VTAIL.n662 9.3005
R767 VTAIL.n714 VTAIL.n713 9.3005
R768 VTAIL.n716 VTAIL.n715 9.3005
R769 VTAIL.n658 VTAIL.n657 9.3005
R770 VTAIL.n722 VTAIL.n721 9.3005
R771 VTAIL.n724 VTAIL.n723 9.3005
R772 VTAIL.n747 VTAIL.n746 9.3005
R773 VTAIL.n646 VTAIL.n645 9.3005
R774 VTAIL.n741 VTAIL.n740 9.3005
R775 VTAIL.n739 VTAIL.n738 9.3005
R776 VTAIL.n650 VTAIL.n649 9.3005
R777 VTAIL.n733 VTAIL.n732 9.3005
R778 VTAIL.n731 VTAIL.n730 9.3005
R779 VTAIL.n654 VTAIL.n653 9.3005
R780 VTAIL.n667 VTAIL.n666 9.3005
R781 VTAIL.n700 VTAIL.n699 9.3005
R782 VTAIL.n698 VTAIL.n697 9.3005
R783 VTAIL.n671 VTAIL.n670 9.3005
R784 VTAIL.n692 VTAIL.n691 9.3005
R785 VTAIL.n690 VTAIL.n689 9.3005
R786 VTAIL.n675 VTAIL.n674 9.3005
R787 VTAIL.n684 VTAIL.n683 9.3005
R788 VTAIL.n682 VTAIL.n681 9.3005
R789 VTAIL.n598 VTAIL.n597 9.3005
R790 VTAIL.n600 VTAIL.n599 9.3005
R791 VTAIL.n555 VTAIL.n554 9.3005
R792 VTAIL.n606 VTAIL.n605 9.3005
R793 VTAIL.n608 VTAIL.n607 9.3005
R794 VTAIL.n550 VTAIL.n549 9.3005
R795 VTAIL.n614 VTAIL.n613 9.3005
R796 VTAIL.n616 VTAIL.n615 9.3005
R797 VTAIL.n639 VTAIL.n638 9.3005
R798 VTAIL.n538 VTAIL.n537 9.3005
R799 VTAIL.n633 VTAIL.n632 9.3005
R800 VTAIL.n631 VTAIL.n630 9.3005
R801 VTAIL.n542 VTAIL.n541 9.3005
R802 VTAIL.n625 VTAIL.n624 9.3005
R803 VTAIL.n623 VTAIL.n622 9.3005
R804 VTAIL.n546 VTAIL.n545 9.3005
R805 VTAIL.n559 VTAIL.n558 9.3005
R806 VTAIL.n592 VTAIL.n591 9.3005
R807 VTAIL.n590 VTAIL.n589 9.3005
R808 VTAIL.n563 VTAIL.n562 9.3005
R809 VTAIL.n584 VTAIL.n583 9.3005
R810 VTAIL.n582 VTAIL.n581 9.3005
R811 VTAIL.n567 VTAIL.n566 9.3005
R812 VTAIL.n576 VTAIL.n575 9.3005
R813 VTAIL.n574 VTAIL.n573 9.3005
R814 VTAIL.n492 VTAIL.n491 9.3005
R815 VTAIL.n494 VTAIL.n493 9.3005
R816 VTAIL.n449 VTAIL.n448 9.3005
R817 VTAIL.n500 VTAIL.n499 9.3005
R818 VTAIL.n502 VTAIL.n501 9.3005
R819 VTAIL.n444 VTAIL.n443 9.3005
R820 VTAIL.n508 VTAIL.n507 9.3005
R821 VTAIL.n510 VTAIL.n509 9.3005
R822 VTAIL.n533 VTAIL.n532 9.3005
R823 VTAIL.n432 VTAIL.n431 9.3005
R824 VTAIL.n527 VTAIL.n526 9.3005
R825 VTAIL.n525 VTAIL.n524 9.3005
R826 VTAIL.n436 VTAIL.n435 9.3005
R827 VTAIL.n519 VTAIL.n518 9.3005
R828 VTAIL.n517 VTAIL.n516 9.3005
R829 VTAIL.n440 VTAIL.n439 9.3005
R830 VTAIL.n453 VTAIL.n452 9.3005
R831 VTAIL.n486 VTAIL.n485 9.3005
R832 VTAIL.n484 VTAIL.n483 9.3005
R833 VTAIL.n457 VTAIL.n456 9.3005
R834 VTAIL.n478 VTAIL.n477 9.3005
R835 VTAIL.n476 VTAIL.n475 9.3005
R836 VTAIL.n461 VTAIL.n460 9.3005
R837 VTAIL.n470 VTAIL.n469 9.3005
R838 VTAIL.n468 VTAIL.n467 9.3005
R839 VTAIL.n384 VTAIL.n383 9.3005
R840 VTAIL.n386 VTAIL.n385 9.3005
R841 VTAIL.n341 VTAIL.n340 9.3005
R842 VTAIL.n392 VTAIL.n391 9.3005
R843 VTAIL.n394 VTAIL.n393 9.3005
R844 VTAIL.n336 VTAIL.n335 9.3005
R845 VTAIL.n400 VTAIL.n399 9.3005
R846 VTAIL.n402 VTAIL.n401 9.3005
R847 VTAIL.n425 VTAIL.n424 9.3005
R848 VTAIL.n324 VTAIL.n323 9.3005
R849 VTAIL.n419 VTAIL.n418 9.3005
R850 VTAIL.n417 VTAIL.n416 9.3005
R851 VTAIL.n328 VTAIL.n327 9.3005
R852 VTAIL.n411 VTAIL.n410 9.3005
R853 VTAIL.n409 VTAIL.n408 9.3005
R854 VTAIL.n332 VTAIL.n331 9.3005
R855 VTAIL.n345 VTAIL.n344 9.3005
R856 VTAIL.n378 VTAIL.n377 9.3005
R857 VTAIL.n376 VTAIL.n375 9.3005
R858 VTAIL.n349 VTAIL.n348 9.3005
R859 VTAIL.n370 VTAIL.n369 9.3005
R860 VTAIL.n368 VTAIL.n367 9.3005
R861 VTAIL.n353 VTAIL.n352 9.3005
R862 VTAIL.n362 VTAIL.n361 9.3005
R863 VTAIL.n360 VTAIL.n359 9.3005
R864 VTAIL.n801 VTAIL.n776 8.92171
R865 VTAIL.n814 VTAIL.n768 8.92171
R866 VTAIL.n848 VTAIL.n847 8.92171
R867 VTAIL.n53 VTAIL.n28 8.92171
R868 VTAIL.n66 VTAIL.n20 8.92171
R869 VTAIL.n100 VTAIL.n99 8.92171
R870 VTAIL.n159 VTAIL.n134 8.92171
R871 VTAIL.n172 VTAIL.n126 8.92171
R872 VTAIL.n206 VTAIL.n205 8.92171
R873 VTAIL.n267 VTAIL.n242 8.92171
R874 VTAIL.n280 VTAIL.n234 8.92171
R875 VTAIL.n314 VTAIL.n313 8.92171
R876 VTAIL.n742 VTAIL.n741 8.92171
R877 VTAIL.n709 VTAIL.n663 8.92171
R878 VTAIL.n696 VTAIL.n671 8.92171
R879 VTAIL.n634 VTAIL.n633 8.92171
R880 VTAIL.n601 VTAIL.n555 8.92171
R881 VTAIL.n588 VTAIL.n563 8.92171
R882 VTAIL.n528 VTAIL.n527 8.92171
R883 VTAIL.n495 VTAIL.n449 8.92171
R884 VTAIL.n482 VTAIL.n457 8.92171
R885 VTAIL.n420 VTAIL.n419 8.92171
R886 VTAIL.n387 VTAIL.n341 8.92171
R887 VTAIL.n374 VTAIL.n349 8.92171
R888 VTAIL.n802 VTAIL.n774 8.14595
R889 VTAIL.n813 VTAIL.n770 8.14595
R890 VTAIL.n851 VTAIL.n752 8.14595
R891 VTAIL.n54 VTAIL.n26 8.14595
R892 VTAIL.n65 VTAIL.n22 8.14595
R893 VTAIL.n103 VTAIL.n4 8.14595
R894 VTAIL.n160 VTAIL.n132 8.14595
R895 VTAIL.n171 VTAIL.n128 8.14595
R896 VTAIL.n209 VTAIL.n110 8.14595
R897 VTAIL.n268 VTAIL.n240 8.14595
R898 VTAIL.n279 VTAIL.n236 8.14595
R899 VTAIL.n317 VTAIL.n218 8.14595
R900 VTAIL.n745 VTAIL.n646 8.14595
R901 VTAIL.n708 VTAIL.n665 8.14595
R902 VTAIL.n697 VTAIL.n669 8.14595
R903 VTAIL.n637 VTAIL.n538 8.14595
R904 VTAIL.n600 VTAIL.n557 8.14595
R905 VTAIL.n589 VTAIL.n561 8.14595
R906 VTAIL.n531 VTAIL.n432 8.14595
R907 VTAIL.n494 VTAIL.n451 8.14595
R908 VTAIL.n483 VTAIL.n455 8.14595
R909 VTAIL.n423 VTAIL.n324 8.14595
R910 VTAIL.n386 VTAIL.n343 8.14595
R911 VTAIL.n375 VTAIL.n347 8.14595
R912 VTAIL.n806 VTAIL.n805 7.3702
R913 VTAIL.n810 VTAIL.n809 7.3702
R914 VTAIL.n852 VTAIL.n750 7.3702
R915 VTAIL.n58 VTAIL.n57 7.3702
R916 VTAIL.n62 VTAIL.n61 7.3702
R917 VTAIL.n104 VTAIL.n2 7.3702
R918 VTAIL.n164 VTAIL.n163 7.3702
R919 VTAIL.n168 VTAIL.n167 7.3702
R920 VTAIL.n210 VTAIL.n108 7.3702
R921 VTAIL.n272 VTAIL.n271 7.3702
R922 VTAIL.n276 VTAIL.n275 7.3702
R923 VTAIL.n318 VTAIL.n216 7.3702
R924 VTAIL.n746 VTAIL.n644 7.3702
R925 VTAIL.n705 VTAIL.n704 7.3702
R926 VTAIL.n701 VTAIL.n700 7.3702
R927 VTAIL.n638 VTAIL.n536 7.3702
R928 VTAIL.n597 VTAIL.n596 7.3702
R929 VTAIL.n593 VTAIL.n592 7.3702
R930 VTAIL.n532 VTAIL.n430 7.3702
R931 VTAIL.n491 VTAIL.n490 7.3702
R932 VTAIL.n487 VTAIL.n486 7.3702
R933 VTAIL.n424 VTAIL.n322 7.3702
R934 VTAIL.n383 VTAIL.n382 7.3702
R935 VTAIL.n379 VTAIL.n378 7.3702
R936 VTAIL.n806 VTAIL.n772 6.59444
R937 VTAIL.n809 VTAIL.n772 6.59444
R938 VTAIL.n854 VTAIL.n750 6.59444
R939 VTAIL.n58 VTAIL.n24 6.59444
R940 VTAIL.n61 VTAIL.n24 6.59444
R941 VTAIL.n106 VTAIL.n2 6.59444
R942 VTAIL.n164 VTAIL.n130 6.59444
R943 VTAIL.n167 VTAIL.n130 6.59444
R944 VTAIL.n212 VTAIL.n108 6.59444
R945 VTAIL.n272 VTAIL.n238 6.59444
R946 VTAIL.n275 VTAIL.n238 6.59444
R947 VTAIL.n320 VTAIL.n216 6.59444
R948 VTAIL.n748 VTAIL.n644 6.59444
R949 VTAIL.n704 VTAIL.n667 6.59444
R950 VTAIL.n701 VTAIL.n667 6.59444
R951 VTAIL.n640 VTAIL.n536 6.59444
R952 VTAIL.n596 VTAIL.n559 6.59444
R953 VTAIL.n593 VTAIL.n559 6.59444
R954 VTAIL.n534 VTAIL.n430 6.59444
R955 VTAIL.n490 VTAIL.n453 6.59444
R956 VTAIL.n487 VTAIL.n453 6.59444
R957 VTAIL.n426 VTAIL.n322 6.59444
R958 VTAIL.n382 VTAIL.n345 6.59444
R959 VTAIL.n379 VTAIL.n345 6.59444
R960 VTAIL.n805 VTAIL.n774 5.81868
R961 VTAIL.n810 VTAIL.n770 5.81868
R962 VTAIL.n852 VTAIL.n851 5.81868
R963 VTAIL.n57 VTAIL.n26 5.81868
R964 VTAIL.n62 VTAIL.n22 5.81868
R965 VTAIL.n104 VTAIL.n103 5.81868
R966 VTAIL.n163 VTAIL.n132 5.81868
R967 VTAIL.n168 VTAIL.n128 5.81868
R968 VTAIL.n210 VTAIL.n209 5.81868
R969 VTAIL.n271 VTAIL.n240 5.81868
R970 VTAIL.n276 VTAIL.n236 5.81868
R971 VTAIL.n318 VTAIL.n317 5.81868
R972 VTAIL.n746 VTAIL.n745 5.81868
R973 VTAIL.n705 VTAIL.n665 5.81868
R974 VTAIL.n700 VTAIL.n669 5.81868
R975 VTAIL.n638 VTAIL.n637 5.81868
R976 VTAIL.n597 VTAIL.n557 5.81868
R977 VTAIL.n592 VTAIL.n561 5.81868
R978 VTAIL.n532 VTAIL.n531 5.81868
R979 VTAIL.n491 VTAIL.n451 5.81868
R980 VTAIL.n486 VTAIL.n455 5.81868
R981 VTAIL.n424 VTAIL.n423 5.81868
R982 VTAIL.n383 VTAIL.n343 5.81868
R983 VTAIL.n378 VTAIL.n347 5.81868
R984 VTAIL.n802 VTAIL.n801 5.04292
R985 VTAIL.n814 VTAIL.n813 5.04292
R986 VTAIL.n848 VTAIL.n752 5.04292
R987 VTAIL.n54 VTAIL.n53 5.04292
R988 VTAIL.n66 VTAIL.n65 5.04292
R989 VTAIL.n100 VTAIL.n4 5.04292
R990 VTAIL.n160 VTAIL.n159 5.04292
R991 VTAIL.n172 VTAIL.n171 5.04292
R992 VTAIL.n206 VTAIL.n110 5.04292
R993 VTAIL.n268 VTAIL.n267 5.04292
R994 VTAIL.n280 VTAIL.n279 5.04292
R995 VTAIL.n314 VTAIL.n218 5.04292
R996 VTAIL.n742 VTAIL.n646 5.04292
R997 VTAIL.n709 VTAIL.n708 5.04292
R998 VTAIL.n697 VTAIL.n696 5.04292
R999 VTAIL.n634 VTAIL.n538 5.04292
R1000 VTAIL.n601 VTAIL.n600 5.04292
R1001 VTAIL.n589 VTAIL.n588 5.04292
R1002 VTAIL.n528 VTAIL.n432 5.04292
R1003 VTAIL.n495 VTAIL.n494 5.04292
R1004 VTAIL.n483 VTAIL.n482 5.04292
R1005 VTAIL.n420 VTAIL.n324 5.04292
R1006 VTAIL.n387 VTAIL.n386 5.04292
R1007 VTAIL.n375 VTAIL.n374 5.04292
R1008 VTAIL.n798 VTAIL.n776 4.26717
R1009 VTAIL.n817 VTAIL.n768 4.26717
R1010 VTAIL.n847 VTAIL.n754 4.26717
R1011 VTAIL.n50 VTAIL.n28 4.26717
R1012 VTAIL.n69 VTAIL.n20 4.26717
R1013 VTAIL.n99 VTAIL.n6 4.26717
R1014 VTAIL.n156 VTAIL.n134 4.26717
R1015 VTAIL.n175 VTAIL.n126 4.26717
R1016 VTAIL.n205 VTAIL.n112 4.26717
R1017 VTAIL.n264 VTAIL.n242 4.26717
R1018 VTAIL.n283 VTAIL.n234 4.26717
R1019 VTAIL.n313 VTAIL.n220 4.26717
R1020 VTAIL.n741 VTAIL.n648 4.26717
R1021 VTAIL.n712 VTAIL.n663 4.26717
R1022 VTAIL.n693 VTAIL.n671 4.26717
R1023 VTAIL.n633 VTAIL.n540 4.26717
R1024 VTAIL.n604 VTAIL.n555 4.26717
R1025 VTAIL.n585 VTAIL.n563 4.26717
R1026 VTAIL.n527 VTAIL.n434 4.26717
R1027 VTAIL.n498 VTAIL.n449 4.26717
R1028 VTAIL.n479 VTAIL.n457 4.26717
R1029 VTAIL.n419 VTAIL.n326 4.26717
R1030 VTAIL.n390 VTAIL.n341 4.26717
R1031 VTAIL.n371 VTAIL.n349 4.26717
R1032 VTAIL.n787 VTAIL.n783 3.70982
R1033 VTAIL.n39 VTAIL.n35 3.70982
R1034 VTAIL.n145 VTAIL.n141 3.70982
R1035 VTAIL.n253 VTAIL.n249 3.70982
R1036 VTAIL.n682 VTAIL.n678 3.70982
R1037 VTAIL.n574 VTAIL.n570 3.70982
R1038 VTAIL.n468 VTAIL.n464 3.70982
R1039 VTAIL.n360 VTAIL.n356 3.70982
R1040 VTAIL.n797 VTAIL.n778 3.49141
R1041 VTAIL.n818 VTAIL.n766 3.49141
R1042 VTAIL.n844 VTAIL.n843 3.49141
R1043 VTAIL.n49 VTAIL.n30 3.49141
R1044 VTAIL.n70 VTAIL.n18 3.49141
R1045 VTAIL.n96 VTAIL.n95 3.49141
R1046 VTAIL.n155 VTAIL.n136 3.49141
R1047 VTAIL.n176 VTAIL.n124 3.49141
R1048 VTAIL.n202 VTAIL.n201 3.49141
R1049 VTAIL.n263 VTAIL.n244 3.49141
R1050 VTAIL.n284 VTAIL.n232 3.49141
R1051 VTAIL.n310 VTAIL.n309 3.49141
R1052 VTAIL.n738 VTAIL.n737 3.49141
R1053 VTAIL.n713 VTAIL.n661 3.49141
R1054 VTAIL.n692 VTAIL.n673 3.49141
R1055 VTAIL.n630 VTAIL.n629 3.49141
R1056 VTAIL.n605 VTAIL.n553 3.49141
R1057 VTAIL.n584 VTAIL.n565 3.49141
R1058 VTAIL.n524 VTAIL.n523 3.49141
R1059 VTAIL.n499 VTAIL.n447 3.49141
R1060 VTAIL.n478 VTAIL.n459 3.49141
R1061 VTAIL.n416 VTAIL.n415 3.49141
R1062 VTAIL.n391 VTAIL.n339 3.49141
R1063 VTAIL.n370 VTAIL.n351 3.49141
R1064 VTAIL.n794 VTAIL.n793 2.71565
R1065 VTAIL.n822 VTAIL.n821 2.71565
R1066 VTAIL.n840 VTAIL.n756 2.71565
R1067 VTAIL.n46 VTAIL.n45 2.71565
R1068 VTAIL.n74 VTAIL.n73 2.71565
R1069 VTAIL.n92 VTAIL.n8 2.71565
R1070 VTAIL.n152 VTAIL.n151 2.71565
R1071 VTAIL.n180 VTAIL.n179 2.71565
R1072 VTAIL.n198 VTAIL.n114 2.71565
R1073 VTAIL.n260 VTAIL.n259 2.71565
R1074 VTAIL.n288 VTAIL.n287 2.71565
R1075 VTAIL.n306 VTAIL.n222 2.71565
R1076 VTAIL.n734 VTAIL.n650 2.71565
R1077 VTAIL.n717 VTAIL.n716 2.71565
R1078 VTAIL.n689 VTAIL.n688 2.71565
R1079 VTAIL.n626 VTAIL.n542 2.71565
R1080 VTAIL.n609 VTAIL.n608 2.71565
R1081 VTAIL.n581 VTAIL.n580 2.71565
R1082 VTAIL.n520 VTAIL.n436 2.71565
R1083 VTAIL.n503 VTAIL.n502 2.71565
R1084 VTAIL.n475 VTAIL.n474 2.71565
R1085 VTAIL.n412 VTAIL.n328 2.71565
R1086 VTAIL.n395 VTAIL.n394 2.71565
R1087 VTAIL.n367 VTAIL.n366 2.71565
R1088 VTAIL.n790 VTAIL.n780 1.93989
R1089 VTAIL.n826 VTAIL.n764 1.93989
R1090 VTAIL.n839 VTAIL.n758 1.93989
R1091 VTAIL.n42 VTAIL.n32 1.93989
R1092 VTAIL.n78 VTAIL.n16 1.93989
R1093 VTAIL.n91 VTAIL.n10 1.93989
R1094 VTAIL.n148 VTAIL.n138 1.93989
R1095 VTAIL.n184 VTAIL.n122 1.93989
R1096 VTAIL.n197 VTAIL.n116 1.93989
R1097 VTAIL.n256 VTAIL.n246 1.93989
R1098 VTAIL.n292 VTAIL.n230 1.93989
R1099 VTAIL.n305 VTAIL.n224 1.93989
R1100 VTAIL.n733 VTAIL.n652 1.93989
R1101 VTAIL.n720 VTAIL.n658 1.93989
R1102 VTAIL.n685 VTAIL.n675 1.93989
R1103 VTAIL.n625 VTAIL.n544 1.93989
R1104 VTAIL.n612 VTAIL.n550 1.93989
R1105 VTAIL.n577 VTAIL.n567 1.93989
R1106 VTAIL.n519 VTAIL.n438 1.93989
R1107 VTAIL.n506 VTAIL.n444 1.93989
R1108 VTAIL.n471 VTAIL.n461 1.93989
R1109 VTAIL.n411 VTAIL.n330 1.93989
R1110 VTAIL.n398 VTAIL.n336 1.93989
R1111 VTAIL.n363 VTAIL.n353 1.93989
R1112 VTAIL.n429 VTAIL.n427 1.78498
R1113 VTAIL.n535 VTAIL.n429 1.78498
R1114 VTAIL.n643 VTAIL.n641 1.78498
R1115 VTAIL.n749 VTAIL.n643 1.78498
R1116 VTAIL.n321 VTAIL.n215 1.78498
R1117 VTAIL.n215 VTAIL.n213 1.78498
R1118 VTAIL.n107 VTAIL.n1 1.78498
R1119 VTAIL VTAIL.n855 1.72679
R1120 VTAIL.n0 VTAIL.t9 1.71671
R1121 VTAIL.n0 VTAIL.t13 1.71671
R1122 VTAIL.n214 VTAIL.t3 1.71671
R1123 VTAIL.n214 VTAIL.t6 1.71671
R1124 VTAIL.n642 VTAIL.t0 1.71671
R1125 VTAIL.n642 VTAIL.t5 1.71671
R1126 VTAIL.n428 VTAIL.t12 1.71671
R1127 VTAIL.n428 VTAIL.t8 1.71671
R1128 VTAIL.n789 VTAIL.n782 1.16414
R1129 VTAIL.n827 VTAIL.n762 1.16414
R1130 VTAIL.n836 VTAIL.n835 1.16414
R1131 VTAIL.n41 VTAIL.n34 1.16414
R1132 VTAIL.n79 VTAIL.n14 1.16414
R1133 VTAIL.n88 VTAIL.n87 1.16414
R1134 VTAIL.n147 VTAIL.n140 1.16414
R1135 VTAIL.n185 VTAIL.n120 1.16414
R1136 VTAIL.n194 VTAIL.n193 1.16414
R1137 VTAIL.n255 VTAIL.n248 1.16414
R1138 VTAIL.n293 VTAIL.n228 1.16414
R1139 VTAIL.n302 VTAIL.n301 1.16414
R1140 VTAIL.n730 VTAIL.n729 1.16414
R1141 VTAIL.n721 VTAIL.n656 1.16414
R1142 VTAIL.n684 VTAIL.n677 1.16414
R1143 VTAIL.n622 VTAIL.n621 1.16414
R1144 VTAIL.n613 VTAIL.n548 1.16414
R1145 VTAIL.n576 VTAIL.n569 1.16414
R1146 VTAIL.n516 VTAIL.n515 1.16414
R1147 VTAIL.n507 VTAIL.n442 1.16414
R1148 VTAIL.n470 VTAIL.n463 1.16414
R1149 VTAIL.n408 VTAIL.n407 1.16414
R1150 VTAIL.n399 VTAIL.n334 1.16414
R1151 VTAIL.n362 VTAIL.n355 1.16414
R1152 VTAIL.n641 VTAIL.n535 0.470328
R1153 VTAIL.n213 VTAIL.n107 0.470328
R1154 VTAIL.n786 VTAIL.n785 0.388379
R1155 VTAIL.n831 VTAIL.n830 0.388379
R1156 VTAIL.n832 VTAIL.n760 0.388379
R1157 VTAIL.n38 VTAIL.n37 0.388379
R1158 VTAIL.n83 VTAIL.n82 0.388379
R1159 VTAIL.n84 VTAIL.n12 0.388379
R1160 VTAIL.n144 VTAIL.n143 0.388379
R1161 VTAIL.n189 VTAIL.n188 0.388379
R1162 VTAIL.n190 VTAIL.n118 0.388379
R1163 VTAIL.n252 VTAIL.n251 0.388379
R1164 VTAIL.n297 VTAIL.n296 0.388379
R1165 VTAIL.n298 VTAIL.n226 0.388379
R1166 VTAIL.n726 VTAIL.n654 0.388379
R1167 VTAIL.n725 VTAIL.n724 0.388379
R1168 VTAIL.n681 VTAIL.n680 0.388379
R1169 VTAIL.n618 VTAIL.n546 0.388379
R1170 VTAIL.n617 VTAIL.n616 0.388379
R1171 VTAIL.n573 VTAIL.n572 0.388379
R1172 VTAIL.n512 VTAIL.n440 0.388379
R1173 VTAIL.n511 VTAIL.n510 0.388379
R1174 VTAIL.n467 VTAIL.n466 0.388379
R1175 VTAIL.n404 VTAIL.n332 0.388379
R1176 VTAIL.n403 VTAIL.n402 0.388379
R1177 VTAIL.n359 VTAIL.n358 0.388379
R1178 VTAIL.n788 VTAIL.n787 0.155672
R1179 VTAIL.n788 VTAIL.n779 0.155672
R1180 VTAIL.n795 VTAIL.n779 0.155672
R1181 VTAIL.n796 VTAIL.n795 0.155672
R1182 VTAIL.n796 VTAIL.n775 0.155672
R1183 VTAIL.n803 VTAIL.n775 0.155672
R1184 VTAIL.n804 VTAIL.n803 0.155672
R1185 VTAIL.n804 VTAIL.n771 0.155672
R1186 VTAIL.n811 VTAIL.n771 0.155672
R1187 VTAIL.n812 VTAIL.n811 0.155672
R1188 VTAIL.n812 VTAIL.n767 0.155672
R1189 VTAIL.n819 VTAIL.n767 0.155672
R1190 VTAIL.n820 VTAIL.n819 0.155672
R1191 VTAIL.n820 VTAIL.n763 0.155672
R1192 VTAIL.n828 VTAIL.n763 0.155672
R1193 VTAIL.n829 VTAIL.n828 0.155672
R1194 VTAIL.n829 VTAIL.n759 0.155672
R1195 VTAIL.n837 VTAIL.n759 0.155672
R1196 VTAIL.n838 VTAIL.n837 0.155672
R1197 VTAIL.n838 VTAIL.n755 0.155672
R1198 VTAIL.n845 VTAIL.n755 0.155672
R1199 VTAIL.n846 VTAIL.n845 0.155672
R1200 VTAIL.n846 VTAIL.n751 0.155672
R1201 VTAIL.n853 VTAIL.n751 0.155672
R1202 VTAIL.n40 VTAIL.n39 0.155672
R1203 VTAIL.n40 VTAIL.n31 0.155672
R1204 VTAIL.n47 VTAIL.n31 0.155672
R1205 VTAIL.n48 VTAIL.n47 0.155672
R1206 VTAIL.n48 VTAIL.n27 0.155672
R1207 VTAIL.n55 VTAIL.n27 0.155672
R1208 VTAIL.n56 VTAIL.n55 0.155672
R1209 VTAIL.n56 VTAIL.n23 0.155672
R1210 VTAIL.n63 VTAIL.n23 0.155672
R1211 VTAIL.n64 VTAIL.n63 0.155672
R1212 VTAIL.n64 VTAIL.n19 0.155672
R1213 VTAIL.n71 VTAIL.n19 0.155672
R1214 VTAIL.n72 VTAIL.n71 0.155672
R1215 VTAIL.n72 VTAIL.n15 0.155672
R1216 VTAIL.n80 VTAIL.n15 0.155672
R1217 VTAIL.n81 VTAIL.n80 0.155672
R1218 VTAIL.n81 VTAIL.n11 0.155672
R1219 VTAIL.n89 VTAIL.n11 0.155672
R1220 VTAIL.n90 VTAIL.n89 0.155672
R1221 VTAIL.n90 VTAIL.n7 0.155672
R1222 VTAIL.n97 VTAIL.n7 0.155672
R1223 VTAIL.n98 VTAIL.n97 0.155672
R1224 VTAIL.n98 VTAIL.n3 0.155672
R1225 VTAIL.n105 VTAIL.n3 0.155672
R1226 VTAIL.n146 VTAIL.n145 0.155672
R1227 VTAIL.n146 VTAIL.n137 0.155672
R1228 VTAIL.n153 VTAIL.n137 0.155672
R1229 VTAIL.n154 VTAIL.n153 0.155672
R1230 VTAIL.n154 VTAIL.n133 0.155672
R1231 VTAIL.n161 VTAIL.n133 0.155672
R1232 VTAIL.n162 VTAIL.n161 0.155672
R1233 VTAIL.n162 VTAIL.n129 0.155672
R1234 VTAIL.n169 VTAIL.n129 0.155672
R1235 VTAIL.n170 VTAIL.n169 0.155672
R1236 VTAIL.n170 VTAIL.n125 0.155672
R1237 VTAIL.n177 VTAIL.n125 0.155672
R1238 VTAIL.n178 VTAIL.n177 0.155672
R1239 VTAIL.n178 VTAIL.n121 0.155672
R1240 VTAIL.n186 VTAIL.n121 0.155672
R1241 VTAIL.n187 VTAIL.n186 0.155672
R1242 VTAIL.n187 VTAIL.n117 0.155672
R1243 VTAIL.n195 VTAIL.n117 0.155672
R1244 VTAIL.n196 VTAIL.n195 0.155672
R1245 VTAIL.n196 VTAIL.n113 0.155672
R1246 VTAIL.n203 VTAIL.n113 0.155672
R1247 VTAIL.n204 VTAIL.n203 0.155672
R1248 VTAIL.n204 VTAIL.n109 0.155672
R1249 VTAIL.n211 VTAIL.n109 0.155672
R1250 VTAIL.n254 VTAIL.n253 0.155672
R1251 VTAIL.n254 VTAIL.n245 0.155672
R1252 VTAIL.n261 VTAIL.n245 0.155672
R1253 VTAIL.n262 VTAIL.n261 0.155672
R1254 VTAIL.n262 VTAIL.n241 0.155672
R1255 VTAIL.n269 VTAIL.n241 0.155672
R1256 VTAIL.n270 VTAIL.n269 0.155672
R1257 VTAIL.n270 VTAIL.n237 0.155672
R1258 VTAIL.n277 VTAIL.n237 0.155672
R1259 VTAIL.n278 VTAIL.n277 0.155672
R1260 VTAIL.n278 VTAIL.n233 0.155672
R1261 VTAIL.n285 VTAIL.n233 0.155672
R1262 VTAIL.n286 VTAIL.n285 0.155672
R1263 VTAIL.n286 VTAIL.n229 0.155672
R1264 VTAIL.n294 VTAIL.n229 0.155672
R1265 VTAIL.n295 VTAIL.n294 0.155672
R1266 VTAIL.n295 VTAIL.n225 0.155672
R1267 VTAIL.n303 VTAIL.n225 0.155672
R1268 VTAIL.n304 VTAIL.n303 0.155672
R1269 VTAIL.n304 VTAIL.n221 0.155672
R1270 VTAIL.n311 VTAIL.n221 0.155672
R1271 VTAIL.n312 VTAIL.n311 0.155672
R1272 VTAIL.n312 VTAIL.n217 0.155672
R1273 VTAIL.n319 VTAIL.n217 0.155672
R1274 VTAIL.n747 VTAIL.n645 0.155672
R1275 VTAIL.n740 VTAIL.n645 0.155672
R1276 VTAIL.n740 VTAIL.n739 0.155672
R1277 VTAIL.n739 VTAIL.n649 0.155672
R1278 VTAIL.n732 VTAIL.n649 0.155672
R1279 VTAIL.n732 VTAIL.n731 0.155672
R1280 VTAIL.n731 VTAIL.n653 0.155672
R1281 VTAIL.n723 VTAIL.n653 0.155672
R1282 VTAIL.n723 VTAIL.n722 0.155672
R1283 VTAIL.n722 VTAIL.n657 0.155672
R1284 VTAIL.n715 VTAIL.n657 0.155672
R1285 VTAIL.n715 VTAIL.n714 0.155672
R1286 VTAIL.n714 VTAIL.n662 0.155672
R1287 VTAIL.n707 VTAIL.n662 0.155672
R1288 VTAIL.n707 VTAIL.n706 0.155672
R1289 VTAIL.n706 VTAIL.n666 0.155672
R1290 VTAIL.n699 VTAIL.n666 0.155672
R1291 VTAIL.n699 VTAIL.n698 0.155672
R1292 VTAIL.n698 VTAIL.n670 0.155672
R1293 VTAIL.n691 VTAIL.n670 0.155672
R1294 VTAIL.n691 VTAIL.n690 0.155672
R1295 VTAIL.n690 VTAIL.n674 0.155672
R1296 VTAIL.n683 VTAIL.n674 0.155672
R1297 VTAIL.n683 VTAIL.n682 0.155672
R1298 VTAIL.n639 VTAIL.n537 0.155672
R1299 VTAIL.n632 VTAIL.n537 0.155672
R1300 VTAIL.n632 VTAIL.n631 0.155672
R1301 VTAIL.n631 VTAIL.n541 0.155672
R1302 VTAIL.n624 VTAIL.n541 0.155672
R1303 VTAIL.n624 VTAIL.n623 0.155672
R1304 VTAIL.n623 VTAIL.n545 0.155672
R1305 VTAIL.n615 VTAIL.n545 0.155672
R1306 VTAIL.n615 VTAIL.n614 0.155672
R1307 VTAIL.n614 VTAIL.n549 0.155672
R1308 VTAIL.n607 VTAIL.n549 0.155672
R1309 VTAIL.n607 VTAIL.n606 0.155672
R1310 VTAIL.n606 VTAIL.n554 0.155672
R1311 VTAIL.n599 VTAIL.n554 0.155672
R1312 VTAIL.n599 VTAIL.n598 0.155672
R1313 VTAIL.n598 VTAIL.n558 0.155672
R1314 VTAIL.n591 VTAIL.n558 0.155672
R1315 VTAIL.n591 VTAIL.n590 0.155672
R1316 VTAIL.n590 VTAIL.n562 0.155672
R1317 VTAIL.n583 VTAIL.n562 0.155672
R1318 VTAIL.n583 VTAIL.n582 0.155672
R1319 VTAIL.n582 VTAIL.n566 0.155672
R1320 VTAIL.n575 VTAIL.n566 0.155672
R1321 VTAIL.n575 VTAIL.n574 0.155672
R1322 VTAIL.n533 VTAIL.n431 0.155672
R1323 VTAIL.n526 VTAIL.n431 0.155672
R1324 VTAIL.n526 VTAIL.n525 0.155672
R1325 VTAIL.n525 VTAIL.n435 0.155672
R1326 VTAIL.n518 VTAIL.n435 0.155672
R1327 VTAIL.n518 VTAIL.n517 0.155672
R1328 VTAIL.n517 VTAIL.n439 0.155672
R1329 VTAIL.n509 VTAIL.n439 0.155672
R1330 VTAIL.n509 VTAIL.n508 0.155672
R1331 VTAIL.n508 VTAIL.n443 0.155672
R1332 VTAIL.n501 VTAIL.n443 0.155672
R1333 VTAIL.n501 VTAIL.n500 0.155672
R1334 VTAIL.n500 VTAIL.n448 0.155672
R1335 VTAIL.n493 VTAIL.n448 0.155672
R1336 VTAIL.n493 VTAIL.n492 0.155672
R1337 VTAIL.n492 VTAIL.n452 0.155672
R1338 VTAIL.n485 VTAIL.n452 0.155672
R1339 VTAIL.n485 VTAIL.n484 0.155672
R1340 VTAIL.n484 VTAIL.n456 0.155672
R1341 VTAIL.n477 VTAIL.n456 0.155672
R1342 VTAIL.n477 VTAIL.n476 0.155672
R1343 VTAIL.n476 VTAIL.n460 0.155672
R1344 VTAIL.n469 VTAIL.n460 0.155672
R1345 VTAIL.n469 VTAIL.n468 0.155672
R1346 VTAIL.n425 VTAIL.n323 0.155672
R1347 VTAIL.n418 VTAIL.n323 0.155672
R1348 VTAIL.n418 VTAIL.n417 0.155672
R1349 VTAIL.n417 VTAIL.n327 0.155672
R1350 VTAIL.n410 VTAIL.n327 0.155672
R1351 VTAIL.n410 VTAIL.n409 0.155672
R1352 VTAIL.n409 VTAIL.n331 0.155672
R1353 VTAIL.n401 VTAIL.n331 0.155672
R1354 VTAIL.n401 VTAIL.n400 0.155672
R1355 VTAIL.n400 VTAIL.n335 0.155672
R1356 VTAIL.n393 VTAIL.n335 0.155672
R1357 VTAIL.n393 VTAIL.n392 0.155672
R1358 VTAIL.n392 VTAIL.n340 0.155672
R1359 VTAIL.n385 VTAIL.n340 0.155672
R1360 VTAIL.n385 VTAIL.n384 0.155672
R1361 VTAIL.n384 VTAIL.n344 0.155672
R1362 VTAIL.n377 VTAIL.n344 0.155672
R1363 VTAIL.n377 VTAIL.n376 0.155672
R1364 VTAIL.n376 VTAIL.n348 0.155672
R1365 VTAIL.n369 VTAIL.n348 0.155672
R1366 VTAIL.n369 VTAIL.n368 0.155672
R1367 VTAIL.n368 VTAIL.n352 0.155672
R1368 VTAIL.n361 VTAIL.n352 0.155672
R1369 VTAIL.n361 VTAIL.n360 0.155672
R1370 VTAIL VTAIL.n1 0.0586897
R1371 VDD2.n2 VDD2.n1 68.8339
R1372 VDD2.n2 VDD2.n0 68.8339
R1373 VDD2 VDD2.n5 68.8309
R1374 VDD2.n4 VDD2.n3 67.997
R1375 VDD2.n4 VDD2.n2 48.0731
R1376 VDD2.n5 VDD2.t2 1.71671
R1377 VDD2.n5 VDD2.t3 1.71671
R1378 VDD2.n3 VDD2.t4 1.71671
R1379 VDD2.n3 VDD2.t0 1.71671
R1380 VDD2.n1 VDD2.t5 1.71671
R1381 VDD2.n1 VDD2.t6 1.71671
R1382 VDD2.n0 VDD2.t1 1.71671
R1383 VDD2.n0 VDD2.t7 1.71671
R1384 VDD2 VDD2.n4 0.950931
R1385 B.n479 B.n478 585
R1386 B.n477 B.n132 585
R1387 B.n476 B.n475 585
R1388 B.n474 B.n133 585
R1389 B.n473 B.n472 585
R1390 B.n471 B.n134 585
R1391 B.n470 B.n469 585
R1392 B.n468 B.n135 585
R1393 B.n467 B.n466 585
R1394 B.n465 B.n136 585
R1395 B.n464 B.n463 585
R1396 B.n462 B.n137 585
R1397 B.n461 B.n460 585
R1398 B.n459 B.n138 585
R1399 B.n458 B.n457 585
R1400 B.n456 B.n139 585
R1401 B.n455 B.n454 585
R1402 B.n453 B.n140 585
R1403 B.n452 B.n451 585
R1404 B.n450 B.n141 585
R1405 B.n449 B.n448 585
R1406 B.n447 B.n142 585
R1407 B.n446 B.n445 585
R1408 B.n444 B.n143 585
R1409 B.n443 B.n442 585
R1410 B.n441 B.n144 585
R1411 B.n440 B.n439 585
R1412 B.n438 B.n145 585
R1413 B.n437 B.n436 585
R1414 B.n435 B.n146 585
R1415 B.n434 B.n433 585
R1416 B.n432 B.n147 585
R1417 B.n431 B.n430 585
R1418 B.n429 B.n148 585
R1419 B.n428 B.n427 585
R1420 B.n426 B.n149 585
R1421 B.n425 B.n424 585
R1422 B.n423 B.n150 585
R1423 B.n422 B.n421 585
R1424 B.n420 B.n151 585
R1425 B.n419 B.n418 585
R1426 B.n417 B.n152 585
R1427 B.n416 B.n415 585
R1428 B.n414 B.n153 585
R1429 B.n413 B.n412 585
R1430 B.n411 B.n154 585
R1431 B.n410 B.n409 585
R1432 B.n408 B.n155 585
R1433 B.n407 B.n406 585
R1434 B.n405 B.n156 585
R1435 B.n404 B.n403 585
R1436 B.n402 B.n157 585
R1437 B.n401 B.n400 585
R1438 B.n399 B.n158 585
R1439 B.n398 B.n397 585
R1440 B.n396 B.n159 585
R1441 B.n395 B.n394 585
R1442 B.n393 B.n160 585
R1443 B.n392 B.n391 585
R1444 B.n390 B.n161 585
R1445 B.n389 B.n388 585
R1446 B.n387 B.n162 585
R1447 B.n386 B.n385 585
R1448 B.n381 B.n163 585
R1449 B.n380 B.n379 585
R1450 B.n378 B.n164 585
R1451 B.n377 B.n376 585
R1452 B.n375 B.n165 585
R1453 B.n374 B.n373 585
R1454 B.n372 B.n166 585
R1455 B.n371 B.n370 585
R1456 B.n369 B.n167 585
R1457 B.n367 B.n366 585
R1458 B.n365 B.n170 585
R1459 B.n364 B.n363 585
R1460 B.n362 B.n171 585
R1461 B.n361 B.n360 585
R1462 B.n359 B.n172 585
R1463 B.n358 B.n357 585
R1464 B.n356 B.n173 585
R1465 B.n355 B.n354 585
R1466 B.n353 B.n174 585
R1467 B.n352 B.n351 585
R1468 B.n350 B.n175 585
R1469 B.n349 B.n348 585
R1470 B.n347 B.n176 585
R1471 B.n346 B.n345 585
R1472 B.n344 B.n177 585
R1473 B.n343 B.n342 585
R1474 B.n341 B.n178 585
R1475 B.n340 B.n339 585
R1476 B.n338 B.n179 585
R1477 B.n337 B.n336 585
R1478 B.n335 B.n180 585
R1479 B.n334 B.n333 585
R1480 B.n332 B.n181 585
R1481 B.n331 B.n330 585
R1482 B.n329 B.n182 585
R1483 B.n328 B.n327 585
R1484 B.n326 B.n183 585
R1485 B.n325 B.n324 585
R1486 B.n323 B.n184 585
R1487 B.n322 B.n321 585
R1488 B.n320 B.n185 585
R1489 B.n319 B.n318 585
R1490 B.n317 B.n186 585
R1491 B.n316 B.n315 585
R1492 B.n314 B.n187 585
R1493 B.n313 B.n312 585
R1494 B.n311 B.n188 585
R1495 B.n310 B.n309 585
R1496 B.n308 B.n189 585
R1497 B.n307 B.n306 585
R1498 B.n305 B.n190 585
R1499 B.n304 B.n303 585
R1500 B.n302 B.n191 585
R1501 B.n301 B.n300 585
R1502 B.n299 B.n192 585
R1503 B.n298 B.n297 585
R1504 B.n296 B.n193 585
R1505 B.n295 B.n294 585
R1506 B.n293 B.n194 585
R1507 B.n292 B.n291 585
R1508 B.n290 B.n195 585
R1509 B.n289 B.n288 585
R1510 B.n287 B.n196 585
R1511 B.n286 B.n285 585
R1512 B.n284 B.n197 585
R1513 B.n283 B.n282 585
R1514 B.n281 B.n198 585
R1515 B.n280 B.n279 585
R1516 B.n278 B.n199 585
R1517 B.n277 B.n276 585
R1518 B.n275 B.n200 585
R1519 B.n480 B.n131 585
R1520 B.n482 B.n481 585
R1521 B.n483 B.n130 585
R1522 B.n485 B.n484 585
R1523 B.n486 B.n129 585
R1524 B.n488 B.n487 585
R1525 B.n489 B.n128 585
R1526 B.n491 B.n490 585
R1527 B.n492 B.n127 585
R1528 B.n494 B.n493 585
R1529 B.n495 B.n126 585
R1530 B.n497 B.n496 585
R1531 B.n498 B.n125 585
R1532 B.n500 B.n499 585
R1533 B.n501 B.n124 585
R1534 B.n503 B.n502 585
R1535 B.n504 B.n123 585
R1536 B.n506 B.n505 585
R1537 B.n507 B.n122 585
R1538 B.n509 B.n508 585
R1539 B.n510 B.n121 585
R1540 B.n512 B.n511 585
R1541 B.n513 B.n120 585
R1542 B.n515 B.n514 585
R1543 B.n516 B.n119 585
R1544 B.n518 B.n517 585
R1545 B.n519 B.n118 585
R1546 B.n521 B.n520 585
R1547 B.n522 B.n117 585
R1548 B.n524 B.n523 585
R1549 B.n525 B.n116 585
R1550 B.n527 B.n526 585
R1551 B.n528 B.n115 585
R1552 B.n530 B.n529 585
R1553 B.n531 B.n114 585
R1554 B.n533 B.n532 585
R1555 B.n534 B.n113 585
R1556 B.n536 B.n535 585
R1557 B.n537 B.n112 585
R1558 B.n539 B.n538 585
R1559 B.n540 B.n111 585
R1560 B.n542 B.n541 585
R1561 B.n543 B.n110 585
R1562 B.n545 B.n544 585
R1563 B.n546 B.n109 585
R1564 B.n548 B.n547 585
R1565 B.n549 B.n108 585
R1566 B.n551 B.n550 585
R1567 B.n552 B.n107 585
R1568 B.n554 B.n553 585
R1569 B.n555 B.n106 585
R1570 B.n557 B.n556 585
R1571 B.n558 B.n105 585
R1572 B.n560 B.n559 585
R1573 B.n561 B.n104 585
R1574 B.n563 B.n562 585
R1575 B.n564 B.n103 585
R1576 B.n566 B.n565 585
R1577 B.n567 B.n102 585
R1578 B.n569 B.n568 585
R1579 B.n570 B.n101 585
R1580 B.n572 B.n571 585
R1581 B.n573 B.n100 585
R1582 B.n575 B.n574 585
R1583 B.n576 B.n99 585
R1584 B.n578 B.n577 585
R1585 B.n579 B.n98 585
R1586 B.n581 B.n580 585
R1587 B.n582 B.n97 585
R1588 B.n584 B.n583 585
R1589 B.n585 B.n96 585
R1590 B.n587 B.n586 585
R1591 B.n588 B.n95 585
R1592 B.n590 B.n589 585
R1593 B.n591 B.n94 585
R1594 B.n593 B.n592 585
R1595 B.n594 B.n93 585
R1596 B.n596 B.n595 585
R1597 B.n798 B.n21 585
R1598 B.n797 B.n796 585
R1599 B.n795 B.n22 585
R1600 B.n794 B.n793 585
R1601 B.n792 B.n23 585
R1602 B.n791 B.n790 585
R1603 B.n789 B.n24 585
R1604 B.n788 B.n787 585
R1605 B.n786 B.n25 585
R1606 B.n785 B.n784 585
R1607 B.n783 B.n26 585
R1608 B.n782 B.n781 585
R1609 B.n780 B.n27 585
R1610 B.n779 B.n778 585
R1611 B.n777 B.n28 585
R1612 B.n776 B.n775 585
R1613 B.n774 B.n29 585
R1614 B.n773 B.n772 585
R1615 B.n771 B.n30 585
R1616 B.n770 B.n769 585
R1617 B.n768 B.n31 585
R1618 B.n767 B.n766 585
R1619 B.n765 B.n32 585
R1620 B.n764 B.n763 585
R1621 B.n762 B.n33 585
R1622 B.n761 B.n760 585
R1623 B.n759 B.n34 585
R1624 B.n758 B.n757 585
R1625 B.n756 B.n35 585
R1626 B.n755 B.n754 585
R1627 B.n753 B.n36 585
R1628 B.n752 B.n751 585
R1629 B.n750 B.n37 585
R1630 B.n749 B.n748 585
R1631 B.n747 B.n38 585
R1632 B.n746 B.n745 585
R1633 B.n744 B.n39 585
R1634 B.n743 B.n742 585
R1635 B.n741 B.n40 585
R1636 B.n740 B.n739 585
R1637 B.n738 B.n41 585
R1638 B.n737 B.n736 585
R1639 B.n735 B.n42 585
R1640 B.n734 B.n733 585
R1641 B.n732 B.n43 585
R1642 B.n731 B.n730 585
R1643 B.n729 B.n44 585
R1644 B.n728 B.n727 585
R1645 B.n726 B.n45 585
R1646 B.n725 B.n724 585
R1647 B.n723 B.n46 585
R1648 B.n722 B.n721 585
R1649 B.n720 B.n47 585
R1650 B.n719 B.n718 585
R1651 B.n717 B.n48 585
R1652 B.n716 B.n715 585
R1653 B.n714 B.n49 585
R1654 B.n713 B.n712 585
R1655 B.n711 B.n50 585
R1656 B.n710 B.n709 585
R1657 B.n708 B.n51 585
R1658 B.n707 B.n706 585
R1659 B.n705 B.n704 585
R1660 B.n703 B.n55 585
R1661 B.n702 B.n701 585
R1662 B.n700 B.n56 585
R1663 B.n699 B.n698 585
R1664 B.n697 B.n57 585
R1665 B.n696 B.n695 585
R1666 B.n694 B.n58 585
R1667 B.n693 B.n692 585
R1668 B.n691 B.n59 585
R1669 B.n689 B.n688 585
R1670 B.n687 B.n62 585
R1671 B.n686 B.n685 585
R1672 B.n684 B.n63 585
R1673 B.n683 B.n682 585
R1674 B.n681 B.n64 585
R1675 B.n680 B.n679 585
R1676 B.n678 B.n65 585
R1677 B.n677 B.n676 585
R1678 B.n675 B.n66 585
R1679 B.n674 B.n673 585
R1680 B.n672 B.n67 585
R1681 B.n671 B.n670 585
R1682 B.n669 B.n68 585
R1683 B.n668 B.n667 585
R1684 B.n666 B.n69 585
R1685 B.n665 B.n664 585
R1686 B.n663 B.n70 585
R1687 B.n662 B.n661 585
R1688 B.n660 B.n71 585
R1689 B.n659 B.n658 585
R1690 B.n657 B.n72 585
R1691 B.n656 B.n655 585
R1692 B.n654 B.n73 585
R1693 B.n653 B.n652 585
R1694 B.n651 B.n74 585
R1695 B.n650 B.n649 585
R1696 B.n648 B.n75 585
R1697 B.n647 B.n646 585
R1698 B.n645 B.n76 585
R1699 B.n644 B.n643 585
R1700 B.n642 B.n77 585
R1701 B.n641 B.n640 585
R1702 B.n639 B.n78 585
R1703 B.n638 B.n637 585
R1704 B.n636 B.n79 585
R1705 B.n635 B.n634 585
R1706 B.n633 B.n80 585
R1707 B.n632 B.n631 585
R1708 B.n630 B.n81 585
R1709 B.n629 B.n628 585
R1710 B.n627 B.n82 585
R1711 B.n626 B.n625 585
R1712 B.n624 B.n83 585
R1713 B.n623 B.n622 585
R1714 B.n621 B.n84 585
R1715 B.n620 B.n619 585
R1716 B.n618 B.n85 585
R1717 B.n617 B.n616 585
R1718 B.n615 B.n86 585
R1719 B.n614 B.n613 585
R1720 B.n612 B.n87 585
R1721 B.n611 B.n610 585
R1722 B.n609 B.n88 585
R1723 B.n608 B.n607 585
R1724 B.n606 B.n89 585
R1725 B.n605 B.n604 585
R1726 B.n603 B.n90 585
R1727 B.n602 B.n601 585
R1728 B.n600 B.n91 585
R1729 B.n599 B.n598 585
R1730 B.n597 B.n92 585
R1731 B.n800 B.n799 585
R1732 B.n801 B.n20 585
R1733 B.n803 B.n802 585
R1734 B.n804 B.n19 585
R1735 B.n806 B.n805 585
R1736 B.n807 B.n18 585
R1737 B.n809 B.n808 585
R1738 B.n810 B.n17 585
R1739 B.n812 B.n811 585
R1740 B.n813 B.n16 585
R1741 B.n815 B.n814 585
R1742 B.n816 B.n15 585
R1743 B.n818 B.n817 585
R1744 B.n819 B.n14 585
R1745 B.n821 B.n820 585
R1746 B.n822 B.n13 585
R1747 B.n824 B.n823 585
R1748 B.n825 B.n12 585
R1749 B.n827 B.n826 585
R1750 B.n828 B.n11 585
R1751 B.n830 B.n829 585
R1752 B.n831 B.n10 585
R1753 B.n833 B.n832 585
R1754 B.n834 B.n9 585
R1755 B.n836 B.n835 585
R1756 B.n837 B.n8 585
R1757 B.n839 B.n838 585
R1758 B.n840 B.n7 585
R1759 B.n842 B.n841 585
R1760 B.n843 B.n6 585
R1761 B.n845 B.n844 585
R1762 B.n846 B.n5 585
R1763 B.n848 B.n847 585
R1764 B.n849 B.n4 585
R1765 B.n851 B.n850 585
R1766 B.n852 B.n3 585
R1767 B.n854 B.n853 585
R1768 B.n855 B.n0 585
R1769 B.n2 B.n1 585
R1770 B.n220 B.n219 585
R1771 B.n221 B.n218 585
R1772 B.n223 B.n222 585
R1773 B.n224 B.n217 585
R1774 B.n226 B.n225 585
R1775 B.n227 B.n216 585
R1776 B.n229 B.n228 585
R1777 B.n230 B.n215 585
R1778 B.n232 B.n231 585
R1779 B.n233 B.n214 585
R1780 B.n235 B.n234 585
R1781 B.n236 B.n213 585
R1782 B.n238 B.n237 585
R1783 B.n239 B.n212 585
R1784 B.n241 B.n240 585
R1785 B.n242 B.n211 585
R1786 B.n244 B.n243 585
R1787 B.n245 B.n210 585
R1788 B.n247 B.n246 585
R1789 B.n248 B.n209 585
R1790 B.n250 B.n249 585
R1791 B.n251 B.n208 585
R1792 B.n253 B.n252 585
R1793 B.n254 B.n207 585
R1794 B.n256 B.n255 585
R1795 B.n257 B.n206 585
R1796 B.n259 B.n258 585
R1797 B.n260 B.n205 585
R1798 B.n262 B.n261 585
R1799 B.n263 B.n204 585
R1800 B.n265 B.n264 585
R1801 B.n266 B.n203 585
R1802 B.n268 B.n267 585
R1803 B.n269 B.n202 585
R1804 B.n271 B.n270 585
R1805 B.n272 B.n201 585
R1806 B.n274 B.n273 585
R1807 B.n382 B.t7 540.87
R1808 B.n60 B.t2 540.87
R1809 B.n168 B.t4 540.87
R1810 B.n52 B.t11 540.87
R1811 B.n383 B.t8 500.726
R1812 B.n61 B.t1 500.726
R1813 B.n169 B.t5 500.724
R1814 B.n53 B.t10 500.724
R1815 B.n275 B.n274 478.086
R1816 B.n478 B.n131 478.086
R1817 B.n597 B.n596 478.086
R1818 B.n800 B.n21 478.086
R1819 B.n168 B.t3 468.565
R1820 B.n382 B.t6 468.565
R1821 B.n60 B.t0 468.565
R1822 B.n52 B.t9 468.565
R1823 B.n857 B.n856 256.663
R1824 B.n856 B.n855 235.042
R1825 B.n856 B.n2 235.042
R1826 B.n276 B.n275 163.367
R1827 B.n276 B.n199 163.367
R1828 B.n280 B.n199 163.367
R1829 B.n281 B.n280 163.367
R1830 B.n282 B.n281 163.367
R1831 B.n282 B.n197 163.367
R1832 B.n286 B.n197 163.367
R1833 B.n287 B.n286 163.367
R1834 B.n288 B.n287 163.367
R1835 B.n288 B.n195 163.367
R1836 B.n292 B.n195 163.367
R1837 B.n293 B.n292 163.367
R1838 B.n294 B.n293 163.367
R1839 B.n294 B.n193 163.367
R1840 B.n298 B.n193 163.367
R1841 B.n299 B.n298 163.367
R1842 B.n300 B.n299 163.367
R1843 B.n300 B.n191 163.367
R1844 B.n304 B.n191 163.367
R1845 B.n305 B.n304 163.367
R1846 B.n306 B.n305 163.367
R1847 B.n306 B.n189 163.367
R1848 B.n310 B.n189 163.367
R1849 B.n311 B.n310 163.367
R1850 B.n312 B.n311 163.367
R1851 B.n312 B.n187 163.367
R1852 B.n316 B.n187 163.367
R1853 B.n317 B.n316 163.367
R1854 B.n318 B.n317 163.367
R1855 B.n318 B.n185 163.367
R1856 B.n322 B.n185 163.367
R1857 B.n323 B.n322 163.367
R1858 B.n324 B.n323 163.367
R1859 B.n324 B.n183 163.367
R1860 B.n328 B.n183 163.367
R1861 B.n329 B.n328 163.367
R1862 B.n330 B.n329 163.367
R1863 B.n330 B.n181 163.367
R1864 B.n334 B.n181 163.367
R1865 B.n335 B.n334 163.367
R1866 B.n336 B.n335 163.367
R1867 B.n336 B.n179 163.367
R1868 B.n340 B.n179 163.367
R1869 B.n341 B.n340 163.367
R1870 B.n342 B.n341 163.367
R1871 B.n342 B.n177 163.367
R1872 B.n346 B.n177 163.367
R1873 B.n347 B.n346 163.367
R1874 B.n348 B.n347 163.367
R1875 B.n348 B.n175 163.367
R1876 B.n352 B.n175 163.367
R1877 B.n353 B.n352 163.367
R1878 B.n354 B.n353 163.367
R1879 B.n354 B.n173 163.367
R1880 B.n358 B.n173 163.367
R1881 B.n359 B.n358 163.367
R1882 B.n360 B.n359 163.367
R1883 B.n360 B.n171 163.367
R1884 B.n364 B.n171 163.367
R1885 B.n365 B.n364 163.367
R1886 B.n366 B.n365 163.367
R1887 B.n366 B.n167 163.367
R1888 B.n371 B.n167 163.367
R1889 B.n372 B.n371 163.367
R1890 B.n373 B.n372 163.367
R1891 B.n373 B.n165 163.367
R1892 B.n377 B.n165 163.367
R1893 B.n378 B.n377 163.367
R1894 B.n379 B.n378 163.367
R1895 B.n379 B.n163 163.367
R1896 B.n386 B.n163 163.367
R1897 B.n387 B.n386 163.367
R1898 B.n388 B.n387 163.367
R1899 B.n388 B.n161 163.367
R1900 B.n392 B.n161 163.367
R1901 B.n393 B.n392 163.367
R1902 B.n394 B.n393 163.367
R1903 B.n394 B.n159 163.367
R1904 B.n398 B.n159 163.367
R1905 B.n399 B.n398 163.367
R1906 B.n400 B.n399 163.367
R1907 B.n400 B.n157 163.367
R1908 B.n404 B.n157 163.367
R1909 B.n405 B.n404 163.367
R1910 B.n406 B.n405 163.367
R1911 B.n406 B.n155 163.367
R1912 B.n410 B.n155 163.367
R1913 B.n411 B.n410 163.367
R1914 B.n412 B.n411 163.367
R1915 B.n412 B.n153 163.367
R1916 B.n416 B.n153 163.367
R1917 B.n417 B.n416 163.367
R1918 B.n418 B.n417 163.367
R1919 B.n418 B.n151 163.367
R1920 B.n422 B.n151 163.367
R1921 B.n423 B.n422 163.367
R1922 B.n424 B.n423 163.367
R1923 B.n424 B.n149 163.367
R1924 B.n428 B.n149 163.367
R1925 B.n429 B.n428 163.367
R1926 B.n430 B.n429 163.367
R1927 B.n430 B.n147 163.367
R1928 B.n434 B.n147 163.367
R1929 B.n435 B.n434 163.367
R1930 B.n436 B.n435 163.367
R1931 B.n436 B.n145 163.367
R1932 B.n440 B.n145 163.367
R1933 B.n441 B.n440 163.367
R1934 B.n442 B.n441 163.367
R1935 B.n442 B.n143 163.367
R1936 B.n446 B.n143 163.367
R1937 B.n447 B.n446 163.367
R1938 B.n448 B.n447 163.367
R1939 B.n448 B.n141 163.367
R1940 B.n452 B.n141 163.367
R1941 B.n453 B.n452 163.367
R1942 B.n454 B.n453 163.367
R1943 B.n454 B.n139 163.367
R1944 B.n458 B.n139 163.367
R1945 B.n459 B.n458 163.367
R1946 B.n460 B.n459 163.367
R1947 B.n460 B.n137 163.367
R1948 B.n464 B.n137 163.367
R1949 B.n465 B.n464 163.367
R1950 B.n466 B.n465 163.367
R1951 B.n466 B.n135 163.367
R1952 B.n470 B.n135 163.367
R1953 B.n471 B.n470 163.367
R1954 B.n472 B.n471 163.367
R1955 B.n472 B.n133 163.367
R1956 B.n476 B.n133 163.367
R1957 B.n477 B.n476 163.367
R1958 B.n478 B.n477 163.367
R1959 B.n596 B.n93 163.367
R1960 B.n592 B.n93 163.367
R1961 B.n592 B.n591 163.367
R1962 B.n591 B.n590 163.367
R1963 B.n590 B.n95 163.367
R1964 B.n586 B.n95 163.367
R1965 B.n586 B.n585 163.367
R1966 B.n585 B.n584 163.367
R1967 B.n584 B.n97 163.367
R1968 B.n580 B.n97 163.367
R1969 B.n580 B.n579 163.367
R1970 B.n579 B.n578 163.367
R1971 B.n578 B.n99 163.367
R1972 B.n574 B.n99 163.367
R1973 B.n574 B.n573 163.367
R1974 B.n573 B.n572 163.367
R1975 B.n572 B.n101 163.367
R1976 B.n568 B.n101 163.367
R1977 B.n568 B.n567 163.367
R1978 B.n567 B.n566 163.367
R1979 B.n566 B.n103 163.367
R1980 B.n562 B.n103 163.367
R1981 B.n562 B.n561 163.367
R1982 B.n561 B.n560 163.367
R1983 B.n560 B.n105 163.367
R1984 B.n556 B.n105 163.367
R1985 B.n556 B.n555 163.367
R1986 B.n555 B.n554 163.367
R1987 B.n554 B.n107 163.367
R1988 B.n550 B.n107 163.367
R1989 B.n550 B.n549 163.367
R1990 B.n549 B.n548 163.367
R1991 B.n548 B.n109 163.367
R1992 B.n544 B.n109 163.367
R1993 B.n544 B.n543 163.367
R1994 B.n543 B.n542 163.367
R1995 B.n542 B.n111 163.367
R1996 B.n538 B.n111 163.367
R1997 B.n538 B.n537 163.367
R1998 B.n537 B.n536 163.367
R1999 B.n536 B.n113 163.367
R2000 B.n532 B.n113 163.367
R2001 B.n532 B.n531 163.367
R2002 B.n531 B.n530 163.367
R2003 B.n530 B.n115 163.367
R2004 B.n526 B.n115 163.367
R2005 B.n526 B.n525 163.367
R2006 B.n525 B.n524 163.367
R2007 B.n524 B.n117 163.367
R2008 B.n520 B.n117 163.367
R2009 B.n520 B.n519 163.367
R2010 B.n519 B.n518 163.367
R2011 B.n518 B.n119 163.367
R2012 B.n514 B.n119 163.367
R2013 B.n514 B.n513 163.367
R2014 B.n513 B.n512 163.367
R2015 B.n512 B.n121 163.367
R2016 B.n508 B.n121 163.367
R2017 B.n508 B.n507 163.367
R2018 B.n507 B.n506 163.367
R2019 B.n506 B.n123 163.367
R2020 B.n502 B.n123 163.367
R2021 B.n502 B.n501 163.367
R2022 B.n501 B.n500 163.367
R2023 B.n500 B.n125 163.367
R2024 B.n496 B.n125 163.367
R2025 B.n496 B.n495 163.367
R2026 B.n495 B.n494 163.367
R2027 B.n494 B.n127 163.367
R2028 B.n490 B.n127 163.367
R2029 B.n490 B.n489 163.367
R2030 B.n489 B.n488 163.367
R2031 B.n488 B.n129 163.367
R2032 B.n484 B.n129 163.367
R2033 B.n484 B.n483 163.367
R2034 B.n483 B.n482 163.367
R2035 B.n482 B.n131 163.367
R2036 B.n796 B.n21 163.367
R2037 B.n796 B.n795 163.367
R2038 B.n795 B.n794 163.367
R2039 B.n794 B.n23 163.367
R2040 B.n790 B.n23 163.367
R2041 B.n790 B.n789 163.367
R2042 B.n789 B.n788 163.367
R2043 B.n788 B.n25 163.367
R2044 B.n784 B.n25 163.367
R2045 B.n784 B.n783 163.367
R2046 B.n783 B.n782 163.367
R2047 B.n782 B.n27 163.367
R2048 B.n778 B.n27 163.367
R2049 B.n778 B.n777 163.367
R2050 B.n777 B.n776 163.367
R2051 B.n776 B.n29 163.367
R2052 B.n772 B.n29 163.367
R2053 B.n772 B.n771 163.367
R2054 B.n771 B.n770 163.367
R2055 B.n770 B.n31 163.367
R2056 B.n766 B.n31 163.367
R2057 B.n766 B.n765 163.367
R2058 B.n765 B.n764 163.367
R2059 B.n764 B.n33 163.367
R2060 B.n760 B.n33 163.367
R2061 B.n760 B.n759 163.367
R2062 B.n759 B.n758 163.367
R2063 B.n758 B.n35 163.367
R2064 B.n754 B.n35 163.367
R2065 B.n754 B.n753 163.367
R2066 B.n753 B.n752 163.367
R2067 B.n752 B.n37 163.367
R2068 B.n748 B.n37 163.367
R2069 B.n748 B.n747 163.367
R2070 B.n747 B.n746 163.367
R2071 B.n746 B.n39 163.367
R2072 B.n742 B.n39 163.367
R2073 B.n742 B.n741 163.367
R2074 B.n741 B.n740 163.367
R2075 B.n740 B.n41 163.367
R2076 B.n736 B.n41 163.367
R2077 B.n736 B.n735 163.367
R2078 B.n735 B.n734 163.367
R2079 B.n734 B.n43 163.367
R2080 B.n730 B.n43 163.367
R2081 B.n730 B.n729 163.367
R2082 B.n729 B.n728 163.367
R2083 B.n728 B.n45 163.367
R2084 B.n724 B.n45 163.367
R2085 B.n724 B.n723 163.367
R2086 B.n723 B.n722 163.367
R2087 B.n722 B.n47 163.367
R2088 B.n718 B.n47 163.367
R2089 B.n718 B.n717 163.367
R2090 B.n717 B.n716 163.367
R2091 B.n716 B.n49 163.367
R2092 B.n712 B.n49 163.367
R2093 B.n712 B.n711 163.367
R2094 B.n711 B.n710 163.367
R2095 B.n710 B.n51 163.367
R2096 B.n706 B.n51 163.367
R2097 B.n706 B.n705 163.367
R2098 B.n705 B.n55 163.367
R2099 B.n701 B.n55 163.367
R2100 B.n701 B.n700 163.367
R2101 B.n700 B.n699 163.367
R2102 B.n699 B.n57 163.367
R2103 B.n695 B.n57 163.367
R2104 B.n695 B.n694 163.367
R2105 B.n694 B.n693 163.367
R2106 B.n693 B.n59 163.367
R2107 B.n688 B.n59 163.367
R2108 B.n688 B.n687 163.367
R2109 B.n687 B.n686 163.367
R2110 B.n686 B.n63 163.367
R2111 B.n682 B.n63 163.367
R2112 B.n682 B.n681 163.367
R2113 B.n681 B.n680 163.367
R2114 B.n680 B.n65 163.367
R2115 B.n676 B.n65 163.367
R2116 B.n676 B.n675 163.367
R2117 B.n675 B.n674 163.367
R2118 B.n674 B.n67 163.367
R2119 B.n670 B.n67 163.367
R2120 B.n670 B.n669 163.367
R2121 B.n669 B.n668 163.367
R2122 B.n668 B.n69 163.367
R2123 B.n664 B.n69 163.367
R2124 B.n664 B.n663 163.367
R2125 B.n663 B.n662 163.367
R2126 B.n662 B.n71 163.367
R2127 B.n658 B.n71 163.367
R2128 B.n658 B.n657 163.367
R2129 B.n657 B.n656 163.367
R2130 B.n656 B.n73 163.367
R2131 B.n652 B.n73 163.367
R2132 B.n652 B.n651 163.367
R2133 B.n651 B.n650 163.367
R2134 B.n650 B.n75 163.367
R2135 B.n646 B.n75 163.367
R2136 B.n646 B.n645 163.367
R2137 B.n645 B.n644 163.367
R2138 B.n644 B.n77 163.367
R2139 B.n640 B.n77 163.367
R2140 B.n640 B.n639 163.367
R2141 B.n639 B.n638 163.367
R2142 B.n638 B.n79 163.367
R2143 B.n634 B.n79 163.367
R2144 B.n634 B.n633 163.367
R2145 B.n633 B.n632 163.367
R2146 B.n632 B.n81 163.367
R2147 B.n628 B.n81 163.367
R2148 B.n628 B.n627 163.367
R2149 B.n627 B.n626 163.367
R2150 B.n626 B.n83 163.367
R2151 B.n622 B.n83 163.367
R2152 B.n622 B.n621 163.367
R2153 B.n621 B.n620 163.367
R2154 B.n620 B.n85 163.367
R2155 B.n616 B.n85 163.367
R2156 B.n616 B.n615 163.367
R2157 B.n615 B.n614 163.367
R2158 B.n614 B.n87 163.367
R2159 B.n610 B.n87 163.367
R2160 B.n610 B.n609 163.367
R2161 B.n609 B.n608 163.367
R2162 B.n608 B.n89 163.367
R2163 B.n604 B.n89 163.367
R2164 B.n604 B.n603 163.367
R2165 B.n603 B.n602 163.367
R2166 B.n602 B.n91 163.367
R2167 B.n598 B.n91 163.367
R2168 B.n598 B.n597 163.367
R2169 B.n801 B.n800 163.367
R2170 B.n802 B.n801 163.367
R2171 B.n802 B.n19 163.367
R2172 B.n806 B.n19 163.367
R2173 B.n807 B.n806 163.367
R2174 B.n808 B.n807 163.367
R2175 B.n808 B.n17 163.367
R2176 B.n812 B.n17 163.367
R2177 B.n813 B.n812 163.367
R2178 B.n814 B.n813 163.367
R2179 B.n814 B.n15 163.367
R2180 B.n818 B.n15 163.367
R2181 B.n819 B.n818 163.367
R2182 B.n820 B.n819 163.367
R2183 B.n820 B.n13 163.367
R2184 B.n824 B.n13 163.367
R2185 B.n825 B.n824 163.367
R2186 B.n826 B.n825 163.367
R2187 B.n826 B.n11 163.367
R2188 B.n830 B.n11 163.367
R2189 B.n831 B.n830 163.367
R2190 B.n832 B.n831 163.367
R2191 B.n832 B.n9 163.367
R2192 B.n836 B.n9 163.367
R2193 B.n837 B.n836 163.367
R2194 B.n838 B.n837 163.367
R2195 B.n838 B.n7 163.367
R2196 B.n842 B.n7 163.367
R2197 B.n843 B.n842 163.367
R2198 B.n844 B.n843 163.367
R2199 B.n844 B.n5 163.367
R2200 B.n848 B.n5 163.367
R2201 B.n849 B.n848 163.367
R2202 B.n850 B.n849 163.367
R2203 B.n850 B.n3 163.367
R2204 B.n854 B.n3 163.367
R2205 B.n855 B.n854 163.367
R2206 B.n220 B.n2 163.367
R2207 B.n221 B.n220 163.367
R2208 B.n222 B.n221 163.367
R2209 B.n222 B.n217 163.367
R2210 B.n226 B.n217 163.367
R2211 B.n227 B.n226 163.367
R2212 B.n228 B.n227 163.367
R2213 B.n228 B.n215 163.367
R2214 B.n232 B.n215 163.367
R2215 B.n233 B.n232 163.367
R2216 B.n234 B.n233 163.367
R2217 B.n234 B.n213 163.367
R2218 B.n238 B.n213 163.367
R2219 B.n239 B.n238 163.367
R2220 B.n240 B.n239 163.367
R2221 B.n240 B.n211 163.367
R2222 B.n244 B.n211 163.367
R2223 B.n245 B.n244 163.367
R2224 B.n246 B.n245 163.367
R2225 B.n246 B.n209 163.367
R2226 B.n250 B.n209 163.367
R2227 B.n251 B.n250 163.367
R2228 B.n252 B.n251 163.367
R2229 B.n252 B.n207 163.367
R2230 B.n256 B.n207 163.367
R2231 B.n257 B.n256 163.367
R2232 B.n258 B.n257 163.367
R2233 B.n258 B.n205 163.367
R2234 B.n262 B.n205 163.367
R2235 B.n263 B.n262 163.367
R2236 B.n264 B.n263 163.367
R2237 B.n264 B.n203 163.367
R2238 B.n268 B.n203 163.367
R2239 B.n269 B.n268 163.367
R2240 B.n270 B.n269 163.367
R2241 B.n270 B.n201 163.367
R2242 B.n274 B.n201 163.367
R2243 B.n368 B.n169 59.5399
R2244 B.n384 B.n383 59.5399
R2245 B.n690 B.n61 59.5399
R2246 B.n54 B.n53 59.5399
R2247 B.n169 B.n168 40.146
R2248 B.n383 B.n382 40.146
R2249 B.n61 B.n60 40.146
R2250 B.n53 B.n52 40.146
R2251 B.n799 B.n798 31.0639
R2252 B.n595 B.n92 31.0639
R2253 B.n480 B.n479 31.0639
R2254 B.n273 B.n200 31.0639
R2255 B B.n857 18.0485
R2256 B.n799 B.n20 10.6151
R2257 B.n803 B.n20 10.6151
R2258 B.n804 B.n803 10.6151
R2259 B.n805 B.n804 10.6151
R2260 B.n805 B.n18 10.6151
R2261 B.n809 B.n18 10.6151
R2262 B.n810 B.n809 10.6151
R2263 B.n811 B.n810 10.6151
R2264 B.n811 B.n16 10.6151
R2265 B.n815 B.n16 10.6151
R2266 B.n816 B.n815 10.6151
R2267 B.n817 B.n816 10.6151
R2268 B.n817 B.n14 10.6151
R2269 B.n821 B.n14 10.6151
R2270 B.n822 B.n821 10.6151
R2271 B.n823 B.n822 10.6151
R2272 B.n823 B.n12 10.6151
R2273 B.n827 B.n12 10.6151
R2274 B.n828 B.n827 10.6151
R2275 B.n829 B.n828 10.6151
R2276 B.n829 B.n10 10.6151
R2277 B.n833 B.n10 10.6151
R2278 B.n834 B.n833 10.6151
R2279 B.n835 B.n834 10.6151
R2280 B.n835 B.n8 10.6151
R2281 B.n839 B.n8 10.6151
R2282 B.n840 B.n839 10.6151
R2283 B.n841 B.n840 10.6151
R2284 B.n841 B.n6 10.6151
R2285 B.n845 B.n6 10.6151
R2286 B.n846 B.n845 10.6151
R2287 B.n847 B.n846 10.6151
R2288 B.n847 B.n4 10.6151
R2289 B.n851 B.n4 10.6151
R2290 B.n852 B.n851 10.6151
R2291 B.n853 B.n852 10.6151
R2292 B.n853 B.n0 10.6151
R2293 B.n798 B.n797 10.6151
R2294 B.n797 B.n22 10.6151
R2295 B.n793 B.n22 10.6151
R2296 B.n793 B.n792 10.6151
R2297 B.n792 B.n791 10.6151
R2298 B.n791 B.n24 10.6151
R2299 B.n787 B.n24 10.6151
R2300 B.n787 B.n786 10.6151
R2301 B.n786 B.n785 10.6151
R2302 B.n785 B.n26 10.6151
R2303 B.n781 B.n26 10.6151
R2304 B.n781 B.n780 10.6151
R2305 B.n780 B.n779 10.6151
R2306 B.n779 B.n28 10.6151
R2307 B.n775 B.n28 10.6151
R2308 B.n775 B.n774 10.6151
R2309 B.n774 B.n773 10.6151
R2310 B.n773 B.n30 10.6151
R2311 B.n769 B.n30 10.6151
R2312 B.n769 B.n768 10.6151
R2313 B.n768 B.n767 10.6151
R2314 B.n767 B.n32 10.6151
R2315 B.n763 B.n32 10.6151
R2316 B.n763 B.n762 10.6151
R2317 B.n762 B.n761 10.6151
R2318 B.n761 B.n34 10.6151
R2319 B.n757 B.n34 10.6151
R2320 B.n757 B.n756 10.6151
R2321 B.n756 B.n755 10.6151
R2322 B.n755 B.n36 10.6151
R2323 B.n751 B.n36 10.6151
R2324 B.n751 B.n750 10.6151
R2325 B.n750 B.n749 10.6151
R2326 B.n749 B.n38 10.6151
R2327 B.n745 B.n38 10.6151
R2328 B.n745 B.n744 10.6151
R2329 B.n744 B.n743 10.6151
R2330 B.n743 B.n40 10.6151
R2331 B.n739 B.n40 10.6151
R2332 B.n739 B.n738 10.6151
R2333 B.n738 B.n737 10.6151
R2334 B.n737 B.n42 10.6151
R2335 B.n733 B.n42 10.6151
R2336 B.n733 B.n732 10.6151
R2337 B.n732 B.n731 10.6151
R2338 B.n731 B.n44 10.6151
R2339 B.n727 B.n44 10.6151
R2340 B.n727 B.n726 10.6151
R2341 B.n726 B.n725 10.6151
R2342 B.n725 B.n46 10.6151
R2343 B.n721 B.n46 10.6151
R2344 B.n721 B.n720 10.6151
R2345 B.n720 B.n719 10.6151
R2346 B.n719 B.n48 10.6151
R2347 B.n715 B.n48 10.6151
R2348 B.n715 B.n714 10.6151
R2349 B.n714 B.n713 10.6151
R2350 B.n713 B.n50 10.6151
R2351 B.n709 B.n50 10.6151
R2352 B.n709 B.n708 10.6151
R2353 B.n708 B.n707 10.6151
R2354 B.n704 B.n703 10.6151
R2355 B.n703 B.n702 10.6151
R2356 B.n702 B.n56 10.6151
R2357 B.n698 B.n56 10.6151
R2358 B.n698 B.n697 10.6151
R2359 B.n697 B.n696 10.6151
R2360 B.n696 B.n58 10.6151
R2361 B.n692 B.n58 10.6151
R2362 B.n692 B.n691 10.6151
R2363 B.n689 B.n62 10.6151
R2364 B.n685 B.n62 10.6151
R2365 B.n685 B.n684 10.6151
R2366 B.n684 B.n683 10.6151
R2367 B.n683 B.n64 10.6151
R2368 B.n679 B.n64 10.6151
R2369 B.n679 B.n678 10.6151
R2370 B.n678 B.n677 10.6151
R2371 B.n677 B.n66 10.6151
R2372 B.n673 B.n66 10.6151
R2373 B.n673 B.n672 10.6151
R2374 B.n672 B.n671 10.6151
R2375 B.n671 B.n68 10.6151
R2376 B.n667 B.n68 10.6151
R2377 B.n667 B.n666 10.6151
R2378 B.n666 B.n665 10.6151
R2379 B.n665 B.n70 10.6151
R2380 B.n661 B.n70 10.6151
R2381 B.n661 B.n660 10.6151
R2382 B.n660 B.n659 10.6151
R2383 B.n659 B.n72 10.6151
R2384 B.n655 B.n72 10.6151
R2385 B.n655 B.n654 10.6151
R2386 B.n654 B.n653 10.6151
R2387 B.n653 B.n74 10.6151
R2388 B.n649 B.n74 10.6151
R2389 B.n649 B.n648 10.6151
R2390 B.n648 B.n647 10.6151
R2391 B.n647 B.n76 10.6151
R2392 B.n643 B.n76 10.6151
R2393 B.n643 B.n642 10.6151
R2394 B.n642 B.n641 10.6151
R2395 B.n641 B.n78 10.6151
R2396 B.n637 B.n78 10.6151
R2397 B.n637 B.n636 10.6151
R2398 B.n636 B.n635 10.6151
R2399 B.n635 B.n80 10.6151
R2400 B.n631 B.n80 10.6151
R2401 B.n631 B.n630 10.6151
R2402 B.n630 B.n629 10.6151
R2403 B.n629 B.n82 10.6151
R2404 B.n625 B.n82 10.6151
R2405 B.n625 B.n624 10.6151
R2406 B.n624 B.n623 10.6151
R2407 B.n623 B.n84 10.6151
R2408 B.n619 B.n84 10.6151
R2409 B.n619 B.n618 10.6151
R2410 B.n618 B.n617 10.6151
R2411 B.n617 B.n86 10.6151
R2412 B.n613 B.n86 10.6151
R2413 B.n613 B.n612 10.6151
R2414 B.n612 B.n611 10.6151
R2415 B.n611 B.n88 10.6151
R2416 B.n607 B.n88 10.6151
R2417 B.n607 B.n606 10.6151
R2418 B.n606 B.n605 10.6151
R2419 B.n605 B.n90 10.6151
R2420 B.n601 B.n90 10.6151
R2421 B.n601 B.n600 10.6151
R2422 B.n600 B.n599 10.6151
R2423 B.n599 B.n92 10.6151
R2424 B.n595 B.n594 10.6151
R2425 B.n594 B.n593 10.6151
R2426 B.n593 B.n94 10.6151
R2427 B.n589 B.n94 10.6151
R2428 B.n589 B.n588 10.6151
R2429 B.n588 B.n587 10.6151
R2430 B.n587 B.n96 10.6151
R2431 B.n583 B.n96 10.6151
R2432 B.n583 B.n582 10.6151
R2433 B.n582 B.n581 10.6151
R2434 B.n581 B.n98 10.6151
R2435 B.n577 B.n98 10.6151
R2436 B.n577 B.n576 10.6151
R2437 B.n576 B.n575 10.6151
R2438 B.n575 B.n100 10.6151
R2439 B.n571 B.n100 10.6151
R2440 B.n571 B.n570 10.6151
R2441 B.n570 B.n569 10.6151
R2442 B.n569 B.n102 10.6151
R2443 B.n565 B.n102 10.6151
R2444 B.n565 B.n564 10.6151
R2445 B.n564 B.n563 10.6151
R2446 B.n563 B.n104 10.6151
R2447 B.n559 B.n104 10.6151
R2448 B.n559 B.n558 10.6151
R2449 B.n558 B.n557 10.6151
R2450 B.n557 B.n106 10.6151
R2451 B.n553 B.n106 10.6151
R2452 B.n553 B.n552 10.6151
R2453 B.n552 B.n551 10.6151
R2454 B.n551 B.n108 10.6151
R2455 B.n547 B.n108 10.6151
R2456 B.n547 B.n546 10.6151
R2457 B.n546 B.n545 10.6151
R2458 B.n545 B.n110 10.6151
R2459 B.n541 B.n110 10.6151
R2460 B.n541 B.n540 10.6151
R2461 B.n540 B.n539 10.6151
R2462 B.n539 B.n112 10.6151
R2463 B.n535 B.n112 10.6151
R2464 B.n535 B.n534 10.6151
R2465 B.n534 B.n533 10.6151
R2466 B.n533 B.n114 10.6151
R2467 B.n529 B.n114 10.6151
R2468 B.n529 B.n528 10.6151
R2469 B.n528 B.n527 10.6151
R2470 B.n527 B.n116 10.6151
R2471 B.n523 B.n116 10.6151
R2472 B.n523 B.n522 10.6151
R2473 B.n522 B.n521 10.6151
R2474 B.n521 B.n118 10.6151
R2475 B.n517 B.n118 10.6151
R2476 B.n517 B.n516 10.6151
R2477 B.n516 B.n515 10.6151
R2478 B.n515 B.n120 10.6151
R2479 B.n511 B.n120 10.6151
R2480 B.n511 B.n510 10.6151
R2481 B.n510 B.n509 10.6151
R2482 B.n509 B.n122 10.6151
R2483 B.n505 B.n122 10.6151
R2484 B.n505 B.n504 10.6151
R2485 B.n504 B.n503 10.6151
R2486 B.n503 B.n124 10.6151
R2487 B.n499 B.n124 10.6151
R2488 B.n499 B.n498 10.6151
R2489 B.n498 B.n497 10.6151
R2490 B.n497 B.n126 10.6151
R2491 B.n493 B.n126 10.6151
R2492 B.n493 B.n492 10.6151
R2493 B.n492 B.n491 10.6151
R2494 B.n491 B.n128 10.6151
R2495 B.n487 B.n128 10.6151
R2496 B.n487 B.n486 10.6151
R2497 B.n486 B.n485 10.6151
R2498 B.n485 B.n130 10.6151
R2499 B.n481 B.n130 10.6151
R2500 B.n481 B.n480 10.6151
R2501 B.n219 B.n1 10.6151
R2502 B.n219 B.n218 10.6151
R2503 B.n223 B.n218 10.6151
R2504 B.n224 B.n223 10.6151
R2505 B.n225 B.n224 10.6151
R2506 B.n225 B.n216 10.6151
R2507 B.n229 B.n216 10.6151
R2508 B.n230 B.n229 10.6151
R2509 B.n231 B.n230 10.6151
R2510 B.n231 B.n214 10.6151
R2511 B.n235 B.n214 10.6151
R2512 B.n236 B.n235 10.6151
R2513 B.n237 B.n236 10.6151
R2514 B.n237 B.n212 10.6151
R2515 B.n241 B.n212 10.6151
R2516 B.n242 B.n241 10.6151
R2517 B.n243 B.n242 10.6151
R2518 B.n243 B.n210 10.6151
R2519 B.n247 B.n210 10.6151
R2520 B.n248 B.n247 10.6151
R2521 B.n249 B.n248 10.6151
R2522 B.n249 B.n208 10.6151
R2523 B.n253 B.n208 10.6151
R2524 B.n254 B.n253 10.6151
R2525 B.n255 B.n254 10.6151
R2526 B.n255 B.n206 10.6151
R2527 B.n259 B.n206 10.6151
R2528 B.n260 B.n259 10.6151
R2529 B.n261 B.n260 10.6151
R2530 B.n261 B.n204 10.6151
R2531 B.n265 B.n204 10.6151
R2532 B.n266 B.n265 10.6151
R2533 B.n267 B.n266 10.6151
R2534 B.n267 B.n202 10.6151
R2535 B.n271 B.n202 10.6151
R2536 B.n272 B.n271 10.6151
R2537 B.n273 B.n272 10.6151
R2538 B.n277 B.n200 10.6151
R2539 B.n278 B.n277 10.6151
R2540 B.n279 B.n278 10.6151
R2541 B.n279 B.n198 10.6151
R2542 B.n283 B.n198 10.6151
R2543 B.n284 B.n283 10.6151
R2544 B.n285 B.n284 10.6151
R2545 B.n285 B.n196 10.6151
R2546 B.n289 B.n196 10.6151
R2547 B.n290 B.n289 10.6151
R2548 B.n291 B.n290 10.6151
R2549 B.n291 B.n194 10.6151
R2550 B.n295 B.n194 10.6151
R2551 B.n296 B.n295 10.6151
R2552 B.n297 B.n296 10.6151
R2553 B.n297 B.n192 10.6151
R2554 B.n301 B.n192 10.6151
R2555 B.n302 B.n301 10.6151
R2556 B.n303 B.n302 10.6151
R2557 B.n303 B.n190 10.6151
R2558 B.n307 B.n190 10.6151
R2559 B.n308 B.n307 10.6151
R2560 B.n309 B.n308 10.6151
R2561 B.n309 B.n188 10.6151
R2562 B.n313 B.n188 10.6151
R2563 B.n314 B.n313 10.6151
R2564 B.n315 B.n314 10.6151
R2565 B.n315 B.n186 10.6151
R2566 B.n319 B.n186 10.6151
R2567 B.n320 B.n319 10.6151
R2568 B.n321 B.n320 10.6151
R2569 B.n321 B.n184 10.6151
R2570 B.n325 B.n184 10.6151
R2571 B.n326 B.n325 10.6151
R2572 B.n327 B.n326 10.6151
R2573 B.n327 B.n182 10.6151
R2574 B.n331 B.n182 10.6151
R2575 B.n332 B.n331 10.6151
R2576 B.n333 B.n332 10.6151
R2577 B.n333 B.n180 10.6151
R2578 B.n337 B.n180 10.6151
R2579 B.n338 B.n337 10.6151
R2580 B.n339 B.n338 10.6151
R2581 B.n339 B.n178 10.6151
R2582 B.n343 B.n178 10.6151
R2583 B.n344 B.n343 10.6151
R2584 B.n345 B.n344 10.6151
R2585 B.n345 B.n176 10.6151
R2586 B.n349 B.n176 10.6151
R2587 B.n350 B.n349 10.6151
R2588 B.n351 B.n350 10.6151
R2589 B.n351 B.n174 10.6151
R2590 B.n355 B.n174 10.6151
R2591 B.n356 B.n355 10.6151
R2592 B.n357 B.n356 10.6151
R2593 B.n357 B.n172 10.6151
R2594 B.n361 B.n172 10.6151
R2595 B.n362 B.n361 10.6151
R2596 B.n363 B.n362 10.6151
R2597 B.n363 B.n170 10.6151
R2598 B.n367 B.n170 10.6151
R2599 B.n370 B.n369 10.6151
R2600 B.n370 B.n166 10.6151
R2601 B.n374 B.n166 10.6151
R2602 B.n375 B.n374 10.6151
R2603 B.n376 B.n375 10.6151
R2604 B.n376 B.n164 10.6151
R2605 B.n380 B.n164 10.6151
R2606 B.n381 B.n380 10.6151
R2607 B.n385 B.n381 10.6151
R2608 B.n389 B.n162 10.6151
R2609 B.n390 B.n389 10.6151
R2610 B.n391 B.n390 10.6151
R2611 B.n391 B.n160 10.6151
R2612 B.n395 B.n160 10.6151
R2613 B.n396 B.n395 10.6151
R2614 B.n397 B.n396 10.6151
R2615 B.n397 B.n158 10.6151
R2616 B.n401 B.n158 10.6151
R2617 B.n402 B.n401 10.6151
R2618 B.n403 B.n402 10.6151
R2619 B.n403 B.n156 10.6151
R2620 B.n407 B.n156 10.6151
R2621 B.n408 B.n407 10.6151
R2622 B.n409 B.n408 10.6151
R2623 B.n409 B.n154 10.6151
R2624 B.n413 B.n154 10.6151
R2625 B.n414 B.n413 10.6151
R2626 B.n415 B.n414 10.6151
R2627 B.n415 B.n152 10.6151
R2628 B.n419 B.n152 10.6151
R2629 B.n420 B.n419 10.6151
R2630 B.n421 B.n420 10.6151
R2631 B.n421 B.n150 10.6151
R2632 B.n425 B.n150 10.6151
R2633 B.n426 B.n425 10.6151
R2634 B.n427 B.n426 10.6151
R2635 B.n427 B.n148 10.6151
R2636 B.n431 B.n148 10.6151
R2637 B.n432 B.n431 10.6151
R2638 B.n433 B.n432 10.6151
R2639 B.n433 B.n146 10.6151
R2640 B.n437 B.n146 10.6151
R2641 B.n438 B.n437 10.6151
R2642 B.n439 B.n438 10.6151
R2643 B.n439 B.n144 10.6151
R2644 B.n443 B.n144 10.6151
R2645 B.n444 B.n443 10.6151
R2646 B.n445 B.n444 10.6151
R2647 B.n445 B.n142 10.6151
R2648 B.n449 B.n142 10.6151
R2649 B.n450 B.n449 10.6151
R2650 B.n451 B.n450 10.6151
R2651 B.n451 B.n140 10.6151
R2652 B.n455 B.n140 10.6151
R2653 B.n456 B.n455 10.6151
R2654 B.n457 B.n456 10.6151
R2655 B.n457 B.n138 10.6151
R2656 B.n461 B.n138 10.6151
R2657 B.n462 B.n461 10.6151
R2658 B.n463 B.n462 10.6151
R2659 B.n463 B.n136 10.6151
R2660 B.n467 B.n136 10.6151
R2661 B.n468 B.n467 10.6151
R2662 B.n469 B.n468 10.6151
R2663 B.n469 B.n134 10.6151
R2664 B.n473 B.n134 10.6151
R2665 B.n474 B.n473 10.6151
R2666 B.n475 B.n474 10.6151
R2667 B.n475 B.n132 10.6151
R2668 B.n479 B.n132 10.6151
R2669 B.n707 B.n54 9.36635
R2670 B.n690 B.n689 9.36635
R2671 B.n368 B.n367 9.36635
R2672 B.n384 B.n162 9.36635
R2673 B.n857 B.n0 8.11757
R2674 B.n857 B.n1 8.11757
R2675 B.n704 B.n54 1.24928
R2676 B.n691 B.n690 1.24928
R2677 B.n369 B.n368 1.24928
R2678 B.n385 B.n384 1.24928
R2679 VP.n12 VP.t7 292.762
R2680 VP.n31 VP.t2 262.33
R2681 VP.n38 VP.t1 262.33
R2682 VP.n46 VP.t3 262.33
R2683 VP.n53 VP.t0 262.33
R2684 VP.n28 VP.t6 262.33
R2685 VP.n21 VP.t5 262.33
R2686 VP.n13 VP.t4 262.33
R2687 VP.n31 VP.n30 180.531
R2688 VP.n54 VP.n53 180.531
R2689 VP.n29 VP.n28 180.531
R2690 VP.n14 VP.n11 161.3
R2691 VP.n16 VP.n15 161.3
R2692 VP.n17 VP.n10 161.3
R2693 VP.n19 VP.n18 161.3
R2694 VP.n20 VP.n9 161.3
R2695 VP.n23 VP.n22 161.3
R2696 VP.n24 VP.n8 161.3
R2697 VP.n26 VP.n25 161.3
R2698 VP.n27 VP.n7 161.3
R2699 VP.n52 VP.n0 161.3
R2700 VP.n51 VP.n50 161.3
R2701 VP.n49 VP.n1 161.3
R2702 VP.n48 VP.n47 161.3
R2703 VP.n45 VP.n2 161.3
R2704 VP.n44 VP.n43 161.3
R2705 VP.n42 VP.n3 161.3
R2706 VP.n41 VP.n40 161.3
R2707 VP.n39 VP.n4 161.3
R2708 VP.n37 VP.n36 161.3
R2709 VP.n35 VP.n5 161.3
R2710 VP.n34 VP.n33 161.3
R2711 VP.n32 VP.n6 161.3
R2712 VP.n13 VP.n12 66.2123
R2713 VP.n30 VP.n29 52.0384
R2714 VP.n33 VP.n5 47.2268
R2715 VP.n51 VP.n1 47.2268
R2716 VP.n26 VP.n8 47.2268
R2717 VP.n40 VP.n3 40.4106
R2718 VP.n44 VP.n3 40.4106
R2719 VP.n19 VP.n10 40.4106
R2720 VP.n15 VP.n10 40.4106
R2721 VP.n37 VP.n5 33.5944
R2722 VP.n47 VP.n1 33.5944
R2723 VP.n22 VP.n8 33.5944
R2724 VP.n33 VP.n32 24.3439
R2725 VP.n40 VP.n39 24.3439
R2726 VP.n45 VP.n44 24.3439
R2727 VP.n52 VP.n51 24.3439
R2728 VP.n27 VP.n26 24.3439
R2729 VP.n20 VP.n19 24.3439
R2730 VP.n15 VP.n14 24.3439
R2731 VP.n38 VP.n37 22.6399
R2732 VP.n47 VP.n46 22.6399
R2733 VP.n22 VP.n21 22.6399
R2734 VP.n12 VP.n11 18.4539
R2735 VP.n32 VP.n31 5.11262
R2736 VP.n53 VP.n52 5.11262
R2737 VP.n28 VP.n27 5.11262
R2738 VP.n39 VP.n38 1.70454
R2739 VP.n46 VP.n45 1.70454
R2740 VP.n21 VP.n20 1.70454
R2741 VP.n14 VP.n13 1.70454
R2742 VP.n16 VP.n11 0.189894
R2743 VP.n17 VP.n16 0.189894
R2744 VP.n18 VP.n17 0.189894
R2745 VP.n18 VP.n9 0.189894
R2746 VP.n23 VP.n9 0.189894
R2747 VP.n24 VP.n23 0.189894
R2748 VP.n25 VP.n24 0.189894
R2749 VP.n25 VP.n7 0.189894
R2750 VP.n29 VP.n7 0.189894
R2751 VP.n30 VP.n6 0.189894
R2752 VP.n34 VP.n6 0.189894
R2753 VP.n35 VP.n34 0.189894
R2754 VP.n36 VP.n35 0.189894
R2755 VP.n36 VP.n4 0.189894
R2756 VP.n41 VP.n4 0.189894
R2757 VP.n42 VP.n41 0.189894
R2758 VP.n43 VP.n42 0.189894
R2759 VP.n43 VP.n2 0.189894
R2760 VP.n48 VP.n2 0.189894
R2761 VP.n49 VP.n48 0.189894
R2762 VP.n50 VP.n49 0.189894
R2763 VP.n50 VP.n0 0.189894
R2764 VP.n54 VP.n0 0.189894
R2765 VP VP.n54 0.0516364
R2766 VDD1 VDD1.n0 68.9475
R2767 VDD1.n3 VDD1.n2 68.8339
R2768 VDD1.n3 VDD1.n1 68.8339
R2769 VDD1.n5 VDD1.n4 67.9968
R2770 VDD1.n5 VDD1.n3 48.6561
R2771 VDD1.n4 VDD1.t2 1.71671
R2772 VDD1.n4 VDD1.t1 1.71671
R2773 VDD1.n0 VDD1.t0 1.71671
R2774 VDD1.n0 VDD1.t3 1.71671
R2775 VDD1.n2 VDD1.t4 1.71671
R2776 VDD1.n2 VDD1.t7 1.71671
R2777 VDD1.n1 VDD1.t5 1.71671
R2778 VDD1.n1 VDD1.t6 1.71671
R2779 VDD1 VDD1.n5 0.834552
C0 B VN 1.10348f
C1 VDD1 w_n3040_n4756# 1.8552f
C2 VP VN 7.89988f
C3 B VP 1.75622f
C4 VN VDD2 12.238f
C5 VTAIL VN 12.069201f
C6 B VDD2 1.6438f
C7 VTAIL B 6.68343f
C8 w_n3040_n4756# VN 6.08603f
C9 VDD1 VN 0.149563f
C10 VP VDD2 0.427547f
C11 VTAIL VP 12.0834f
C12 w_n3040_n4756# B 10.7441f
C13 VDD1 B 1.57483f
C14 VTAIL VDD2 11.2232f
C15 w_n3040_n4756# VP 6.47815f
C16 VDD1 VP 12.5151f
C17 w_n3040_n4756# VDD2 1.93384f
C18 VTAIL w_n3040_n4756# 5.77233f
C19 VDD1 VDD2 1.32805f
C20 VTAIL VDD1 11.1746f
C21 VDD2 VSUBS 1.765094f
C22 VDD1 VSUBS 2.259762f
C23 VTAIL VSUBS 1.484158f
C24 VN VSUBS 6.03106f
C25 VP VSUBS 2.947119f
C26 B VSUBS 4.628628f
C27 w_n3040_n4756# VSUBS 0.176673p
C28 VDD1.t0 VSUBS 0.373638f
C29 VDD1.t3 VSUBS 0.373638f
C30 VDD1.n0 VSUBS 3.13008f
C31 VDD1.t5 VSUBS 0.373638f
C32 VDD1.t6 VSUBS 0.373638f
C33 VDD1.n1 VSUBS 3.12878f
C34 VDD1.t4 VSUBS 0.373638f
C35 VDD1.t7 VSUBS 0.373638f
C36 VDD1.n2 VSUBS 3.12878f
C37 VDD1.n3 VSUBS 3.84286f
C38 VDD1.t2 VSUBS 0.373638f
C39 VDD1.t1 VSUBS 0.373638f
C40 VDD1.n4 VSUBS 3.12002f
C41 VDD1.n5 VSUBS 3.49812f
C42 VP.n0 VSUBS 0.033293f
C43 VP.t0 VSUBS 3.02072f
C44 VP.n1 VSUBS 0.029114f
C45 VP.n2 VSUBS 0.033293f
C46 VP.t3 VSUBS 3.02072f
C47 VP.n3 VSUBS 0.026941f
C48 VP.n4 VSUBS 0.033293f
C49 VP.t1 VSUBS 3.02072f
C50 VP.n5 VSUBS 0.029114f
C51 VP.n6 VSUBS 0.033293f
C52 VP.t2 VSUBS 3.02072f
C53 VP.n7 VSUBS 0.033293f
C54 VP.t6 VSUBS 3.02072f
C55 VP.n8 VSUBS 0.029114f
C56 VP.n9 VSUBS 0.033293f
C57 VP.t5 VSUBS 3.02072f
C58 VP.n10 VSUBS 0.026941f
C59 VP.n11 VSUBS 0.21437f
C60 VP.t4 VSUBS 3.02072f
C61 VP.t7 VSUBS 3.14551f
C62 VP.n12 VSUBS 1.14614f
C63 VP.n13 VSUBS 1.11464f
C64 VP.n14 VSUBS 0.033726f
C65 VP.n15 VSUBS 0.066523f
C66 VP.n16 VSUBS 0.033293f
C67 VP.n17 VSUBS 0.033293f
C68 VP.n18 VSUBS 0.033293f
C69 VP.n19 VSUBS 0.066523f
C70 VP.n20 VSUBS 0.033726f
C71 VP.n21 VSUBS 1.05573f
C72 VP.n22 VSUBS 0.065462f
C73 VP.n23 VSUBS 0.033293f
C74 VP.n24 VSUBS 0.033293f
C75 VP.n25 VSUBS 0.033293f
C76 VP.n26 VSUBS 0.063256f
C77 VP.n27 VSUBS 0.038037f
C78 VP.n28 VSUBS 1.13043f
C79 VP.n29 VSUBS 1.9299f
C80 VP.n30 VSUBS 1.95283f
C81 VP.n31 VSUBS 1.13043f
C82 VP.n32 VSUBS 0.038037f
C83 VP.n33 VSUBS 0.063256f
C84 VP.n34 VSUBS 0.033293f
C85 VP.n35 VSUBS 0.033293f
C86 VP.n36 VSUBS 0.033293f
C87 VP.n37 VSUBS 0.065462f
C88 VP.n38 VSUBS 1.05573f
C89 VP.n39 VSUBS 0.033726f
C90 VP.n40 VSUBS 0.066523f
C91 VP.n41 VSUBS 0.033293f
C92 VP.n42 VSUBS 0.033293f
C93 VP.n43 VSUBS 0.033293f
C94 VP.n44 VSUBS 0.066523f
C95 VP.n45 VSUBS 0.033726f
C96 VP.n46 VSUBS 1.05573f
C97 VP.n47 VSUBS 0.065462f
C98 VP.n48 VSUBS 0.033293f
C99 VP.n49 VSUBS 0.033293f
C100 VP.n50 VSUBS 0.033293f
C101 VP.n51 VSUBS 0.063256f
C102 VP.n52 VSUBS 0.038037f
C103 VP.n53 VSUBS 1.13043f
C104 VP.n54 VSUBS 0.034707f
C105 B.n0 VSUBS 0.005811f
C106 B.n1 VSUBS 0.005811f
C107 B.n2 VSUBS 0.008595f
C108 B.n3 VSUBS 0.006586f
C109 B.n4 VSUBS 0.006586f
C110 B.n5 VSUBS 0.006586f
C111 B.n6 VSUBS 0.006586f
C112 B.n7 VSUBS 0.006586f
C113 B.n8 VSUBS 0.006586f
C114 B.n9 VSUBS 0.006586f
C115 B.n10 VSUBS 0.006586f
C116 B.n11 VSUBS 0.006586f
C117 B.n12 VSUBS 0.006586f
C118 B.n13 VSUBS 0.006586f
C119 B.n14 VSUBS 0.006586f
C120 B.n15 VSUBS 0.006586f
C121 B.n16 VSUBS 0.006586f
C122 B.n17 VSUBS 0.006586f
C123 B.n18 VSUBS 0.006586f
C124 B.n19 VSUBS 0.006586f
C125 B.n20 VSUBS 0.006586f
C126 B.n21 VSUBS 0.015465f
C127 B.n22 VSUBS 0.006586f
C128 B.n23 VSUBS 0.006586f
C129 B.n24 VSUBS 0.006586f
C130 B.n25 VSUBS 0.006586f
C131 B.n26 VSUBS 0.006586f
C132 B.n27 VSUBS 0.006586f
C133 B.n28 VSUBS 0.006586f
C134 B.n29 VSUBS 0.006586f
C135 B.n30 VSUBS 0.006586f
C136 B.n31 VSUBS 0.006586f
C137 B.n32 VSUBS 0.006586f
C138 B.n33 VSUBS 0.006586f
C139 B.n34 VSUBS 0.006586f
C140 B.n35 VSUBS 0.006586f
C141 B.n36 VSUBS 0.006586f
C142 B.n37 VSUBS 0.006586f
C143 B.n38 VSUBS 0.006586f
C144 B.n39 VSUBS 0.006586f
C145 B.n40 VSUBS 0.006586f
C146 B.n41 VSUBS 0.006586f
C147 B.n42 VSUBS 0.006586f
C148 B.n43 VSUBS 0.006586f
C149 B.n44 VSUBS 0.006586f
C150 B.n45 VSUBS 0.006586f
C151 B.n46 VSUBS 0.006586f
C152 B.n47 VSUBS 0.006586f
C153 B.n48 VSUBS 0.006586f
C154 B.n49 VSUBS 0.006586f
C155 B.n50 VSUBS 0.006586f
C156 B.n51 VSUBS 0.006586f
C157 B.t10 VSUBS 0.351898f
C158 B.t11 VSUBS 0.374682f
C159 B.t9 VSUBS 1.32916f
C160 B.n52 VSUBS 0.533376f
C161 B.n53 VSUBS 0.316344f
C162 B.n54 VSUBS 0.01526f
C163 B.n55 VSUBS 0.006586f
C164 B.n56 VSUBS 0.006586f
C165 B.n57 VSUBS 0.006586f
C166 B.n58 VSUBS 0.006586f
C167 B.n59 VSUBS 0.006586f
C168 B.t1 VSUBS 0.351902f
C169 B.t2 VSUBS 0.374685f
C170 B.t0 VSUBS 1.32916f
C171 B.n60 VSUBS 0.533373f
C172 B.n61 VSUBS 0.316341f
C173 B.n62 VSUBS 0.006586f
C174 B.n63 VSUBS 0.006586f
C175 B.n64 VSUBS 0.006586f
C176 B.n65 VSUBS 0.006586f
C177 B.n66 VSUBS 0.006586f
C178 B.n67 VSUBS 0.006586f
C179 B.n68 VSUBS 0.006586f
C180 B.n69 VSUBS 0.006586f
C181 B.n70 VSUBS 0.006586f
C182 B.n71 VSUBS 0.006586f
C183 B.n72 VSUBS 0.006586f
C184 B.n73 VSUBS 0.006586f
C185 B.n74 VSUBS 0.006586f
C186 B.n75 VSUBS 0.006586f
C187 B.n76 VSUBS 0.006586f
C188 B.n77 VSUBS 0.006586f
C189 B.n78 VSUBS 0.006586f
C190 B.n79 VSUBS 0.006586f
C191 B.n80 VSUBS 0.006586f
C192 B.n81 VSUBS 0.006586f
C193 B.n82 VSUBS 0.006586f
C194 B.n83 VSUBS 0.006586f
C195 B.n84 VSUBS 0.006586f
C196 B.n85 VSUBS 0.006586f
C197 B.n86 VSUBS 0.006586f
C198 B.n87 VSUBS 0.006586f
C199 B.n88 VSUBS 0.006586f
C200 B.n89 VSUBS 0.006586f
C201 B.n90 VSUBS 0.006586f
C202 B.n91 VSUBS 0.006586f
C203 B.n92 VSUBS 0.015465f
C204 B.n93 VSUBS 0.006586f
C205 B.n94 VSUBS 0.006586f
C206 B.n95 VSUBS 0.006586f
C207 B.n96 VSUBS 0.006586f
C208 B.n97 VSUBS 0.006586f
C209 B.n98 VSUBS 0.006586f
C210 B.n99 VSUBS 0.006586f
C211 B.n100 VSUBS 0.006586f
C212 B.n101 VSUBS 0.006586f
C213 B.n102 VSUBS 0.006586f
C214 B.n103 VSUBS 0.006586f
C215 B.n104 VSUBS 0.006586f
C216 B.n105 VSUBS 0.006586f
C217 B.n106 VSUBS 0.006586f
C218 B.n107 VSUBS 0.006586f
C219 B.n108 VSUBS 0.006586f
C220 B.n109 VSUBS 0.006586f
C221 B.n110 VSUBS 0.006586f
C222 B.n111 VSUBS 0.006586f
C223 B.n112 VSUBS 0.006586f
C224 B.n113 VSUBS 0.006586f
C225 B.n114 VSUBS 0.006586f
C226 B.n115 VSUBS 0.006586f
C227 B.n116 VSUBS 0.006586f
C228 B.n117 VSUBS 0.006586f
C229 B.n118 VSUBS 0.006586f
C230 B.n119 VSUBS 0.006586f
C231 B.n120 VSUBS 0.006586f
C232 B.n121 VSUBS 0.006586f
C233 B.n122 VSUBS 0.006586f
C234 B.n123 VSUBS 0.006586f
C235 B.n124 VSUBS 0.006586f
C236 B.n125 VSUBS 0.006586f
C237 B.n126 VSUBS 0.006586f
C238 B.n127 VSUBS 0.006586f
C239 B.n128 VSUBS 0.006586f
C240 B.n129 VSUBS 0.006586f
C241 B.n130 VSUBS 0.006586f
C242 B.n131 VSUBS 0.014367f
C243 B.n132 VSUBS 0.006586f
C244 B.n133 VSUBS 0.006586f
C245 B.n134 VSUBS 0.006586f
C246 B.n135 VSUBS 0.006586f
C247 B.n136 VSUBS 0.006586f
C248 B.n137 VSUBS 0.006586f
C249 B.n138 VSUBS 0.006586f
C250 B.n139 VSUBS 0.006586f
C251 B.n140 VSUBS 0.006586f
C252 B.n141 VSUBS 0.006586f
C253 B.n142 VSUBS 0.006586f
C254 B.n143 VSUBS 0.006586f
C255 B.n144 VSUBS 0.006586f
C256 B.n145 VSUBS 0.006586f
C257 B.n146 VSUBS 0.006586f
C258 B.n147 VSUBS 0.006586f
C259 B.n148 VSUBS 0.006586f
C260 B.n149 VSUBS 0.006586f
C261 B.n150 VSUBS 0.006586f
C262 B.n151 VSUBS 0.006586f
C263 B.n152 VSUBS 0.006586f
C264 B.n153 VSUBS 0.006586f
C265 B.n154 VSUBS 0.006586f
C266 B.n155 VSUBS 0.006586f
C267 B.n156 VSUBS 0.006586f
C268 B.n157 VSUBS 0.006586f
C269 B.n158 VSUBS 0.006586f
C270 B.n159 VSUBS 0.006586f
C271 B.n160 VSUBS 0.006586f
C272 B.n161 VSUBS 0.006586f
C273 B.n162 VSUBS 0.006199f
C274 B.n163 VSUBS 0.006586f
C275 B.n164 VSUBS 0.006586f
C276 B.n165 VSUBS 0.006586f
C277 B.n166 VSUBS 0.006586f
C278 B.n167 VSUBS 0.006586f
C279 B.t5 VSUBS 0.351898f
C280 B.t4 VSUBS 0.374682f
C281 B.t3 VSUBS 1.32916f
C282 B.n168 VSUBS 0.533376f
C283 B.n169 VSUBS 0.316344f
C284 B.n170 VSUBS 0.006586f
C285 B.n171 VSUBS 0.006586f
C286 B.n172 VSUBS 0.006586f
C287 B.n173 VSUBS 0.006586f
C288 B.n174 VSUBS 0.006586f
C289 B.n175 VSUBS 0.006586f
C290 B.n176 VSUBS 0.006586f
C291 B.n177 VSUBS 0.006586f
C292 B.n178 VSUBS 0.006586f
C293 B.n179 VSUBS 0.006586f
C294 B.n180 VSUBS 0.006586f
C295 B.n181 VSUBS 0.006586f
C296 B.n182 VSUBS 0.006586f
C297 B.n183 VSUBS 0.006586f
C298 B.n184 VSUBS 0.006586f
C299 B.n185 VSUBS 0.006586f
C300 B.n186 VSUBS 0.006586f
C301 B.n187 VSUBS 0.006586f
C302 B.n188 VSUBS 0.006586f
C303 B.n189 VSUBS 0.006586f
C304 B.n190 VSUBS 0.006586f
C305 B.n191 VSUBS 0.006586f
C306 B.n192 VSUBS 0.006586f
C307 B.n193 VSUBS 0.006586f
C308 B.n194 VSUBS 0.006586f
C309 B.n195 VSUBS 0.006586f
C310 B.n196 VSUBS 0.006586f
C311 B.n197 VSUBS 0.006586f
C312 B.n198 VSUBS 0.006586f
C313 B.n199 VSUBS 0.006586f
C314 B.n200 VSUBS 0.015465f
C315 B.n201 VSUBS 0.006586f
C316 B.n202 VSUBS 0.006586f
C317 B.n203 VSUBS 0.006586f
C318 B.n204 VSUBS 0.006586f
C319 B.n205 VSUBS 0.006586f
C320 B.n206 VSUBS 0.006586f
C321 B.n207 VSUBS 0.006586f
C322 B.n208 VSUBS 0.006586f
C323 B.n209 VSUBS 0.006586f
C324 B.n210 VSUBS 0.006586f
C325 B.n211 VSUBS 0.006586f
C326 B.n212 VSUBS 0.006586f
C327 B.n213 VSUBS 0.006586f
C328 B.n214 VSUBS 0.006586f
C329 B.n215 VSUBS 0.006586f
C330 B.n216 VSUBS 0.006586f
C331 B.n217 VSUBS 0.006586f
C332 B.n218 VSUBS 0.006586f
C333 B.n219 VSUBS 0.006586f
C334 B.n220 VSUBS 0.006586f
C335 B.n221 VSUBS 0.006586f
C336 B.n222 VSUBS 0.006586f
C337 B.n223 VSUBS 0.006586f
C338 B.n224 VSUBS 0.006586f
C339 B.n225 VSUBS 0.006586f
C340 B.n226 VSUBS 0.006586f
C341 B.n227 VSUBS 0.006586f
C342 B.n228 VSUBS 0.006586f
C343 B.n229 VSUBS 0.006586f
C344 B.n230 VSUBS 0.006586f
C345 B.n231 VSUBS 0.006586f
C346 B.n232 VSUBS 0.006586f
C347 B.n233 VSUBS 0.006586f
C348 B.n234 VSUBS 0.006586f
C349 B.n235 VSUBS 0.006586f
C350 B.n236 VSUBS 0.006586f
C351 B.n237 VSUBS 0.006586f
C352 B.n238 VSUBS 0.006586f
C353 B.n239 VSUBS 0.006586f
C354 B.n240 VSUBS 0.006586f
C355 B.n241 VSUBS 0.006586f
C356 B.n242 VSUBS 0.006586f
C357 B.n243 VSUBS 0.006586f
C358 B.n244 VSUBS 0.006586f
C359 B.n245 VSUBS 0.006586f
C360 B.n246 VSUBS 0.006586f
C361 B.n247 VSUBS 0.006586f
C362 B.n248 VSUBS 0.006586f
C363 B.n249 VSUBS 0.006586f
C364 B.n250 VSUBS 0.006586f
C365 B.n251 VSUBS 0.006586f
C366 B.n252 VSUBS 0.006586f
C367 B.n253 VSUBS 0.006586f
C368 B.n254 VSUBS 0.006586f
C369 B.n255 VSUBS 0.006586f
C370 B.n256 VSUBS 0.006586f
C371 B.n257 VSUBS 0.006586f
C372 B.n258 VSUBS 0.006586f
C373 B.n259 VSUBS 0.006586f
C374 B.n260 VSUBS 0.006586f
C375 B.n261 VSUBS 0.006586f
C376 B.n262 VSUBS 0.006586f
C377 B.n263 VSUBS 0.006586f
C378 B.n264 VSUBS 0.006586f
C379 B.n265 VSUBS 0.006586f
C380 B.n266 VSUBS 0.006586f
C381 B.n267 VSUBS 0.006586f
C382 B.n268 VSUBS 0.006586f
C383 B.n269 VSUBS 0.006586f
C384 B.n270 VSUBS 0.006586f
C385 B.n271 VSUBS 0.006586f
C386 B.n272 VSUBS 0.006586f
C387 B.n273 VSUBS 0.014367f
C388 B.n274 VSUBS 0.014367f
C389 B.n275 VSUBS 0.015465f
C390 B.n276 VSUBS 0.006586f
C391 B.n277 VSUBS 0.006586f
C392 B.n278 VSUBS 0.006586f
C393 B.n279 VSUBS 0.006586f
C394 B.n280 VSUBS 0.006586f
C395 B.n281 VSUBS 0.006586f
C396 B.n282 VSUBS 0.006586f
C397 B.n283 VSUBS 0.006586f
C398 B.n284 VSUBS 0.006586f
C399 B.n285 VSUBS 0.006586f
C400 B.n286 VSUBS 0.006586f
C401 B.n287 VSUBS 0.006586f
C402 B.n288 VSUBS 0.006586f
C403 B.n289 VSUBS 0.006586f
C404 B.n290 VSUBS 0.006586f
C405 B.n291 VSUBS 0.006586f
C406 B.n292 VSUBS 0.006586f
C407 B.n293 VSUBS 0.006586f
C408 B.n294 VSUBS 0.006586f
C409 B.n295 VSUBS 0.006586f
C410 B.n296 VSUBS 0.006586f
C411 B.n297 VSUBS 0.006586f
C412 B.n298 VSUBS 0.006586f
C413 B.n299 VSUBS 0.006586f
C414 B.n300 VSUBS 0.006586f
C415 B.n301 VSUBS 0.006586f
C416 B.n302 VSUBS 0.006586f
C417 B.n303 VSUBS 0.006586f
C418 B.n304 VSUBS 0.006586f
C419 B.n305 VSUBS 0.006586f
C420 B.n306 VSUBS 0.006586f
C421 B.n307 VSUBS 0.006586f
C422 B.n308 VSUBS 0.006586f
C423 B.n309 VSUBS 0.006586f
C424 B.n310 VSUBS 0.006586f
C425 B.n311 VSUBS 0.006586f
C426 B.n312 VSUBS 0.006586f
C427 B.n313 VSUBS 0.006586f
C428 B.n314 VSUBS 0.006586f
C429 B.n315 VSUBS 0.006586f
C430 B.n316 VSUBS 0.006586f
C431 B.n317 VSUBS 0.006586f
C432 B.n318 VSUBS 0.006586f
C433 B.n319 VSUBS 0.006586f
C434 B.n320 VSUBS 0.006586f
C435 B.n321 VSUBS 0.006586f
C436 B.n322 VSUBS 0.006586f
C437 B.n323 VSUBS 0.006586f
C438 B.n324 VSUBS 0.006586f
C439 B.n325 VSUBS 0.006586f
C440 B.n326 VSUBS 0.006586f
C441 B.n327 VSUBS 0.006586f
C442 B.n328 VSUBS 0.006586f
C443 B.n329 VSUBS 0.006586f
C444 B.n330 VSUBS 0.006586f
C445 B.n331 VSUBS 0.006586f
C446 B.n332 VSUBS 0.006586f
C447 B.n333 VSUBS 0.006586f
C448 B.n334 VSUBS 0.006586f
C449 B.n335 VSUBS 0.006586f
C450 B.n336 VSUBS 0.006586f
C451 B.n337 VSUBS 0.006586f
C452 B.n338 VSUBS 0.006586f
C453 B.n339 VSUBS 0.006586f
C454 B.n340 VSUBS 0.006586f
C455 B.n341 VSUBS 0.006586f
C456 B.n342 VSUBS 0.006586f
C457 B.n343 VSUBS 0.006586f
C458 B.n344 VSUBS 0.006586f
C459 B.n345 VSUBS 0.006586f
C460 B.n346 VSUBS 0.006586f
C461 B.n347 VSUBS 0.006586f
C462 B.n348 VSUBS 0.006586f
C463 B.n349 VSUBS 0.006586f
C464 B.n350 VSUBS 0.006586f
C465 B.n351 VSUBS 0.006586f
C466 B.n352 VSUBS 0.006586f
C467 B.n353 VSUBS 0.006586f
C468 B.n354 VSUBS 0.006586f
C469 B.n355 VSUBS 0.006586f
C470 B.n356 VSUBS 0.006586f
C471 B.n357 VSUBS 0.006586f
C472 B.n358 VSUBS 0.006586f
C473 B.n359 VSUBS 0.006586f
C474 B.n360 VSUBS 0.006586f
C475 B.n361 VSUBS 0.006586f
C476 B.n362 VSUBS 0.006586f
C477 B.n363 VSUBS 0.006586f
C478 B.n364 VSUBS 0.006586f
C479 B.n365 VSUBS 0.006586f
C480 B.n366 VSUBS 0.006586f
C481 B.n367 VSUBS 0.006199f
C482 B.n368 VSUBS 0.01526f
C483 B.n369 VSUBS 0.003681f
C484 B.n370 VSUBS 0.006586f
C485 B.n371 VSUBS 0.006586f
C486 B.n372 VSUBS 0.006586f
C487 B.n373 VSUBS 0.006586f
C488 B.n374 VSUBS 0.006586f
C489 B.n375 VSUBS 0.006586f
C490 B.n376 VSUBS 0.006586f
C491 B.n377 VSUBS 0.006586f
C492 B.n378 VSUBS 0.006586f
C493 B.n379 VSUBS 0.006586f
C494 B.n380 VSUBS 0.006586f
C495 B.n381 VSUBS 0.006586f
C496 B.t8 VSUBS 0.351902f
C497 B.t7 VSUBS 0.374685f
C498 B.t6 VSUBS 1.32916f
C499 B.n382 VSUBS 0.533373f
C500 B.n383 VSUBS 0.316341f
C501 B.n384 VSUBS 0.01526f
C502 B.n385 VSUBS 0.003681f
C503 B.n386 VSUBS 0.006586f
C504 B.n387 VSUBS 0.006586f
C505 B.n388 VSUBS 0.006586f
C506 B.n389 VSUBS 0.006586f
C507 B.n390 VSUBS 0.006586f
C508 B.n391 VSUBS 0.006586f
C509 B.n392 VSUBS 0.006586f
C510 B.n393 VSUBS 0.006586f
C511 B.n394 VSUBS 0.006586f
C512 B.n395 VSUBS 0.006586f
C513 B.n396 VSUBS 0.006586f
C514 B.n397 VSUBS 0.006586f
C515 B.n398 VSUBS 0.006586f
C516 B.n399 VSUBS 0.006586f
C517 B.n400 VSUBS 0.006586f
C518 B.n401 VSUBS 0.006586f
C519 B.n402 VSUBS 0.006586f
C520 B.n403 VSUBS 0.006586f
C521 B.n404 VSUBS 0.006586f
C522 B.n405 VSUBS 0.006586f
C523 B.n406 VSUBS 0.006586f
C524 B.n407 VSUBS 0.006586f
C525 B.n408 VSUBS 0.006586f
C526 B.n409 VSUBS 0.006586f
C527 B.n410 VSUBS 0.006586f
C528 B.n411 VSUBS 0.006586f
C529 B.n412 VSUBS 0.006586f
C530 B.n413 VSUBS 0.006586f
C531 B.n414 VSUBS 0.006586f
C532 B.n415 VSUBS 0.006586f
C533 B.n416 VSUBS 0.006586f
C534 B.n417 VSUBS 0.006586f
C535 B.n418 VSUBS 0.006586f
C536 B.n419 VSUBS 0.006586f
C537 B.n420 VSUBS 0.006586f
C538 B.n421 VSUBS 0.006586f
C539 B.n422 VSUBS 0.006586f
C540 B.n423 VSUBS 0.006586f
C541 B.n424 VSUBS 0.006586f
C542 B.n425 VSUBS 0.006586f
C543 B.n426 VSUBS 0.006586f
C544 B.n427 VSUBS 0.006586f
C545 B.n428 VSUBS 0.006586f
C546 B.n429 VSUBS 0.006586f
C547 B.n430 VSUBS 0.006586f
C548 B.n431 VSUBS 0.006586f
C549 B.n432 VSUBS 0.006586f
C550 B.n433 VSUBS 0.006586f
C551 B.n434 VSUBS 0.006586f
C552 B.n435 VSUBS 0.006586f
C553 B.n436 VSUBS 0.006586f
C554 B.n437 VSUBS 0.006586f
C555 B.n438 VSUBS 0.006586f
C556 B.n439 VSUBS 0.006586f
C557 B.n440 VSUBS 0.006586f
C558 B.n441 VSUBS 0.006586f
C559 B.n442 VSUBS 0.006586f
C560 B.n443 VSUBS 0.006586f
C561 B.n444 VSUBS 0.006586f
C562 B.n445 VSUBS 0.006586f
C563 B.n446 VSUBS 0.006586f
C564 B.n447 VSUBS 0.006586f
C565 B.n448 VSUBS 0.006586f
C566 B.n449 VSUBS 0.006586f
C567 B.n450 VSUBS 0.006586f
C568 B.n451 VSUBS 0.006586f
C569 B.n452 VSUBS 0.006586f
C570 B.n453 VSUBS 0.006586f
C571 B.n454 VSUBS 0.006586f
C572 B.n455 VSUBS 0.006586f
C573 B.n456 VSUBS 0.006586f
C574 B.n457 VSUBS 0.006586f
C575 B.n458 VSUBS 0.006586f
C576 B.n459 VSUBS 0.006586f
C577 B.n460 VSUBS 0.006586f
C578 B.n461 VSUBS 0.006586f
C579 B.n462 VSUBS 0.006586f
C580 B.n463 VSUBS 0.006586f
C581 B.n464 VSUBS 0.006586f
C582 B.n465 VSUBS 0.006586f
C583 B.n466 VSUBS 0.006586f
C584 B.n467 VSUBS 0.006586f
C585 B.n468 VSUBS 0.006586f
C586 B.n469 VSUBS 0.006586f
C587 B.n470 VSUBS 0.006586f
C588 B.n471 VSUBS 0.006586f
C589 B.n472 VSUBS 0.006586f
C590 B.n473 VSUBS 0.006586f
C591 B.n474 VSUBS 0.006586f
C592 B.n475 VSUBS 0.006586f
C593 B.n476 VSUBS 0.006586f
C594 B.n477 VSUBS 0.006586f
C595 B.n478 VSUBS 0.015465f
C596 B.n479 VSUBS 0.014647f
C597 B.n480 VSUBS 0.015186f
C598 B.n481 VSUBS 0.006586f
C599 B.n482 VSUBS 0.006586f
C600 B.n483 VSUBS 0.006586f
C601 B.n484 VSUBS 0.006586f
C602 B.n485 VSUBS 0.006586f
C603 B.n486 VSUBS 0.006586f
C604 B.n487 VSUBS 0.006586f
C605 B.n488 VSUBS 0.006586f
C606 B.n489 VSUBS 0.006586f
C607 B.n490 VSUBS 0.006586f
C608 B.n491 VSUBS 0.006586f
C609 B.n492 VSUBS 0.006586f
C610 B.n493 VSUBS 0.006586f
C611 B.n494 VSUBS 0.006586f
C612 B.n495 VSUBS 0.006586f
C613 B.n496 VSUBS 0.006586f
C614 B.n497 VSUBS 0.006586f
C615 B.n498 VSUBS 0.006586f
C616 B.n499 VSUBS 0.006586f
C617 B.n500 VSUBS 0.006586f
C618 B.n501 VSUBS 0.006586f
C619 B.n502 VSUBS 0.006586f
C620 B.n503 VSUBS 0.006586f
C621 B.n504 VSUBS 0.006586f
C622 B.n505 VSUBS 0.006586f
C623 B.n506 VSUBS 0.006586f
C624 B.n507 VSUBS 0.006586f
C625 B.n508 VSUBS 0.006586f
C626 B.n509 VSUBS 0.006586f
C627 B.n510 VSUBS 0.006586f
C628 B.n511 VSUBS 0.006586f
C629 B.n512 VSUBS 0.006586f
C630 B.n513 VSUBS 0.006586f
C631 B.n514 VSUBS 0.006586f
C632 B.n515 VSUBS 0.006586f
C633 B.n516 VSUBS 0.006586f
C634 B.n517 VSUBS 0.006586f
C635 B.n518 VSUBS 0.006586f
C636 B.n519 VSUBS 0.006586f
C637 B.n520 VSUBS 0.006586f
C638 B.n521 VSUBS 0.006586f
C639 B.n522 VSUBS 0.006586f
C640 B.n523 VSUBS 0.006586f
C641 B.n524 VSUBS 0.006586f
C642 B.n525 VSUBS 0.006586f
C643 B.n526 VSUBS 0.006586f
C644 B.n527 VSUBS 0.006586f
C645 B.n528 VSUBS 0.006586f
C646 B.n529 VSUBS 0.006586f
C647 B.n530 VSUBS 0.006586f
C648 B.n531 VSUBS 0.006586f
C649 B.n532 VSUBS 0.006586f
C650 B.n533 VSUBS 0.006586f
C651 B.n534 VSUBS 0.006586f
C652 B.n535 VSUBS 0.006586f
C653 B.n536 VSUBS 0.006586f
C654 B.n537 VSUBS 0.006586f
C655 B.n538 VSUBS 0.006586f
C656 B.n539 VSUBS 0.006586f
C657 B.n540 VSUBS 0.006586f
C658 B.n541 VSUBS 0.006586f
C659 B.n542 VSUBS 0.006586f
C660 B.n543 VSUBS 0.006586f
C661 B.n544 VSUBS 0.006586f
C662 B.n545 VSUBS 0.006586f
C663 B.n546 VSUBS 0.006586f
C664 B.n547 VSUBS 0.006586f
C665 B.n548 VSUBS 0.006586f
C666 B.n549 VSUBS 0.006586f
C667 B.n550 VSUBS 0.006586f
C668 B.n551 VSUBS 0.006586f
C669 B.n552 VSUBS 0.006586f
C670 B.n553 VSUBS 0.006586f
C671 B.n554 VSUBS 0.006586f
C672 B.n555 VSUBS 0.006586f
C673 B.n556 VSUBS 0.006586f
C674 B.n557 VSUBS 0.006586f
C675 B.n558 VSUBS 0.006586f
C676 B.n559 VSUBS 0.006586f
C677 B.n560 VSUBS 0.006586f
C678 B.n561 VSUBS 0.006586f
C679 B.n562 VSUBS 0.006586f
C680 B.n563 VSUBS 0.006586f
C681 B.n564 VSUBS 0.006586f
C682 B.n565 VSUBS 0.006586f
C683 B.n566 VSUBS 0.006586f
C684 B.n567 VSUBS 0.006586f
C685 B.n568 VSUBS 0.006586f
C686 B.n569 VSUBS 0.006586f
C687 B.n570 VSUBS 0.006586f
C688 B.n571 VSUBS 0.006586f
C689 B.n572 VSUBS 0.006586f
C690 B.n573 VSUBS 0.006586f
C691 B.n574 VSUBS 0.006586f
C692 B.n575 VSUBS 0.006586f
C693 B.n576 VSUBS 0.006586f
C694 B.n577 VSUBS 0.006586f
C695 B.n578 VSUBS 0.006586f
C696 B.n579 VSUBS 0.006586f
C697 B.n580 VSUBS 0.006586f
C698 B.n581 VSUBS 0.006586f
C699 B.n582 VSUBS 0.006586f
C700 B.n583 VSUBS 0.006586f
C701 B.n584 VSUBS 0.006586f
C702 B.n585 VSUBS 0.006586f
C703 B.n586 VSUBS 0.006586f
C704 B.n587 VSUBS 0.006586f
C705 B.n588 VSUBS 0.006586f
C706 B.n589 VSUBS 0.006586f
C707 B.n590 VSUBS 0.006586f
C708 B.n591 VSUBS 0.006586f
C709 B.n592 VSUBS 0.006586f
C710 B.n593 VSUBS 0.006586f
C711 B.n594 VSUBS 0.006586f
C712 B.n595 VSUBS 0.014367f
C713 B.n596 VSUBS 0.014367f
C714 B.n597 VSUBS 0.015465f
C715 B.n598 VSUBS 0.006586f
C716 B.n599 VSUBS 0.006586f
C717 B.n600 VSUBS 0.006586f
C718 B.n601 VSUBS 0.006586f
C719 B.n602 VSUBS 0.006586f
C720 B.n603 VSUBS 0.006586f
C721 B.n604 VSUBS 0.006586f
C722 B.n605 VSUBS 0.006586f
C723 B.n606 VSUBS 0.006586f
C724 B.n607 VSUBS 0.006586f
C725 B.n608 VSUBS 0.006586f
C726 B.n609 VSUBS 0.006586f
C727 B.n610 VSUBS 0.006586f
C728 B.n611 VSUBS 0.006586f
C729 B.n612 VSUBS 0.006586f
C730 B.n613 VSUBS 0.006586f
C731 B.n614 VSUBS 0.006586f
C732 B.n615 VSUBS 0.006586f
C733 B.n616 VSUBS 0.006586f
C734 B.n617 VSUBS 0.006586f
C735 B.n618 VSUBS 0.006586f
C736 B.n619 VSUBS 0.006586f
C737 B.n620 VSUBS 0.006586f
C738 B.n621 VSUBS 0.006586f
C739 B.n622 VSUBS 0.006586f
C740 B.n623 VSUBS 0.006586f
C741 B.n624 VSUBS 0.006586f
C742 B.n625 VSUBS 0.006586f
C743 B.n626 VSUBS 0.006586f
C744 B.n627 VSUBS 0.006586f
C745 B.n628 VSUBS 0.006586f
C746 B.n629 VSUBS 0.006586f
C747 B.n630 VSUBS 0.006586f
C748 B.n631 VSUBS 0.006586f
C749 B.n632 VSUBS 0.006586f
C750 B.n633 VSUBS 0.006586f
C751 B.n634 VSUBS 0.006586f
C752 B.n635 VSUBS 0.006586f
C753 B.n636 VSUBS 0.006586f
C754 B.n637 VSUBS 0.006586f
C755 B.n638 VSUBS 0.006586f
C756 B.n639 VSUBS 0.006586f
C757 B.n640 VSUBS 0.006586f
C758 B.n641 VSUBS 0.006586f
C759 B.n642 VSUBS 0.006586f
C760 B.n643 VSUBS 0.006586f
C761 B.n644 VSUBS 0.006586f
C762 B.n645 VSUBS 0.006586f
C763 B.n646 VSUBS 0.006586f
C764 B.n647 VSUBS 0.006586f
C765 B.n648 VSUBS 0.006586f
C766 B.n649 VSUBS 0.006586f
C767 B.n650 VSUBS 0.006586f
C768 B.n651 VSUBS 0.006586f
C769 B.n652 VSUBS 0.006586f
C770 B.n653 VSUBS 0.006586f
C771 B.n654 VSUBS 0.006586f
C772 B.n655 VSUBS 0.006586f
C773 B.n656 VSUBS 0.006586f
C774 B.n657 VSUBS 0.006586f
C775 B.n658 VSUBS 0.006586f
C776 B.n659 VSUBS 0.006586f
C777 B.n660 VSUBS 0.006586f
C778 B.n661 VSUBS 0.006586f
C779 B.n662 VSUBS 0.006586f
C780 B.n663 VSUBS 0.006586f
C781 B.n664 VSUBS 0.006586f
C782 B.n665 VSUBS 0.006586f
C783 B.n666 VSUBS 0.006586f
C784 B.n667 VSUBS 0.006586f
C785 B.n668 VSUBS 0.006586f
C786 B.n669 VSUBS 0.006586f
C787 B.n670 VSUBS 0.006586f
C788 B.n671 VSUBS 0.006586f
C789 B.n672 VSUBS 0.006586f
C790 B.n673 VSUBS 0.006586f
C791 B.n674 VSUBS 0.006586f
C792 B.n675 VSUBS 0.006586f
C793 B.n676 VSUBS 0.006586f
C794 B.n677 VSUBS 0.006586f
C795 B.n678 VSUBS 0.006586f
C796 B.n679 VSUBS 0.006586f
C797 B.n680 VSUBS 0.006586f
C798 B.n681 VSUBS 0.006586f
C799 B.n682 VSUBS 0.006586f
C800 B.n683 VSUBS 0.006586f
C801 B.n684 VSUBS 0.006586f
C802 B.n685 VSUBS 0.006586f
C803 B.n686 VSUBS 0.006586f
C804 B.n687 VSUBS 0.006586f
C805 B.n688 VSUBS 0.006586f
C806 B.n689 VSUBS 0.006199f
C807 B.n690 VSUBS 0.01526f
C808 B.n691 VSUBS 0.003681f
C809 B.n692 VSUBS 0.006586f
C810 B.n693 VSUBS 0.006586f
C811 B.n694 VSUBS 0.006586f
C812 B.n695 VSUBS 0.006586f
C813 B.n696 VSUBS 0.006586f
C814 B.n697 VSUBS 0.006586f
C815 B.n698 VSUBS 0.006586f
C816 B.n699 VSUBS 0.006586f
C817 B.n700 VSUBS 0.006586f
C818 B.n701 VSUBS 0.006586f
C819 B.n702 VSUBS 0.006586f
C820 B.n703 VSUBS 0.006586f
C821 B.n704 VSUBS 0.003681f
C822 B.n705 VSUBS 0.006586f
C823 B.n706 VSUBS 0.006586f
C824 B.n707 VSUBS 0.006199f
C825 B.n708 VSUBS 0.006586f
C826 B.n709 VSUBS 0.006586f
C827 B.n710 VSUBS 0.006586f
C828 B.n711 VSUBS 0.006586f
C829 B.n712 VSUBS 0.006586f
C830 B.n713 VSUBS 0.006586f
C831 B.n714 VSUBS 0.006586f
C832 B.n715 VSUBS 0.006586f
C833 B.n716 VSUBS 0.006586f
C834 B.n717 VSUBS 0.006586f
C835 B.n718 VSUBS 0.006586f
C836 B.n719 VSUBS 0.006586f
C837 B.n720 VSUBS 0.006586f
C838 B.n721 VSUBS 0.006586f
C839 B.n722 VSUBS 0.006586f
C840 B.n723 VSUBS 0.006586f
C841 B.n724 VSUBS 0.006586f
C842 B.n725 VSUBS 0.006586f
C843 B.n726 VSUBS 0.006586f
C844 B.n727 VSUBS 0.006586f
C845 B.n728 VSUBS 0.006586f
C846 B.n729 VSUBS 0.006586f
C847 B.n730 VSUBS 0.006586f
C848 B.n731 VSUBS 0.006586f
C849 B.n732 VSUBS 0.006586f
C850 B.n733 VSUBS 0.006586f
C851 B.n734 VSUBS 0.006586f
C852 B.n735 VSUBS 0.006586f
C853 B.n736 VSUBS 0.006586f
C854 B.n737 VSUBS 0.006586f
C855 B.n738 VSUBS 0.006586f
C856 B.n739 VSUBS 0.006586f
C857 B.n740 VSUBS 0.006586f
C858 B.n741 VSUBS 0.006586f
C859 B.n742 VSUBS 0.006586f
C860 B.n743 VSUBS 0.006586f
C861 B.n744 VSUBS 0.006586f
C862 B.n745 VSUBS 0.006586f
C863 B.n746 VSUBS 0.006586f
C864 B.n747 VSUBS 0.006586f
C865 B.n748 VSUBS 0.006586f
C866 B.n749 VSUBS 0.006586f
C867 B.n750 VSUBS 0.006586f
C868 B.n751 VSUBS 0.006586f
C869 B.n752 VSUBS 0.006586f
C870 B.n753 VSUBS 0.006586f
C871 B.n754 VSUBS 0.006586f
C872 B.n755 VSUBS 0.006586f
C873 B.n756 VSUBS 0.006586f
C874 B.n757 VSUBS 0.006586f
C875 B.n758 VSUBS 0.006586f
C876 B.n759 VSUBS 0.006586f
C877 B.n760 VSUBS 0.006586f
C878 B.n761 VSUBS 0.006586f
C879 B.n762 VSUBS 0.006586f
C880 B.n763 VSUBS 0.006586f
C881 B.n764 VSUBS 0.006586f
C882 B.n765 VSUBS 0.006586f
C883 B.n766 VSUBS 0.006586f
C884 B.n767 VSUBS 0.006586f
C885 B.n768 VSUBS 0.006586f
C886 B.n769 VSUBS 0.006586f
C887 B.n770 VSUBS 0.006586f
C888 B.n771 VSUBS 0.006586f
C889 B.n772 VSUBS 0.006586f
C890 B.n773 VSUBS 0.006586f
C891 B.n774 VSUBS 0.006586f
C892 B.n775 VSUBS 0.006586f
C893 B.n776 VSUBS 0.006586f
C894 B.n777 VSUBS 0.006586f
C895 B.n778 VSUBS 0.006586f
C896 B.n779 VSUBS 0.006586f
C897 B.n780 VSUBS 0.006586f
C898 B.n781 VSUBS 0.006586f
C899 B.n782 VSUBS 0.006586f
C900 B.n783 VSUBS 0.006586f
C901 B.n784 VSUBS 0.006586f
C902 B.n785 VSUBS 0.006586f
C903 B.n786 VSUBS 0.006586f
C904 B.n787 VSUBS 0.006586f
C905 B.n788 VSUBS 0.006586f
C906 B.n789 VSUBS 0.006586f
C907 B.n790 VSUBS 0.006586f
C908 B.n791 VSUBS 0.006586f
C909 B.n792 VSUBS 0.006586f
C910 B.n793 VSUBS 0.006586f
C911 B.n794 VSUBS 0.006586f
C912 B.n795 VSUBS 0.006586f
C913 B.n796 VSUBS 0.006586f
C914 B.n797 VSUBS 0.006586f
C915 B.n798 VSUBS 0.015465f
C916 B.n799 VSUBS 0.014367f
C917 B.n800 VSUBS 0.014367f
C918 B.n801 VSUBS 0.006586f
C919 B.n802 VSUBS 0.006586f
C920 B.n803 VSUBS 0.006586f
C921 B.n804 VSUBS 0.006586f
C922 B.n805 VSUBS 0.006586f
C923 B.n806 VSUBS 0.006586f
C924 B.n807 VSUBS 0.006586f
C925 B.n808 VSUBS 0.006586f
C926 B.n809 VSUBS 0.006586f
C927 B.n810 VSUBS 0.006586f
C928 B.n811 VSUBS 0.006586f
C929 B.n812 VSUBS 0.006586f
C930 B.n813 VSUBS 0.006586f
C931 B.n814 VSUBS 0.006586f
C932 B.n815 VSUBS 0.006586f
C933 B.n816 VSUBS 0.006586f
C934 B.n817 VSUBS 0.006586f
C935 B.n818 VSUBS 0.006586f
C936 B.n819 VSUBS 0.006586f
C937 B.n820 VSUBS 0.006586f
C938 B.n821 VSUBS 0.006586f
C939 B.n822 VSUBS 0.006586f
C940 B.n823 VSUBS 0.006586f
C941 B.n824 VSUBS 0.006586f
C942 B.n825 VSUBS 0.006586f
C943 B.n826 VSUBS 0.006586f
C944 B.n827 VSUBS 0.006586f
C945 B.n828 VSUBS 0.006586f
C946 B.n829 VSUBS 0.006586f
C947 B.n830 VSUBS 0.006586f
C948 B.n831 VSUBS 0.006586f
C949 B.n832 VSUBS 0.006586f
C950 B.n833 VSUBS 0.006586f
C951 B.n834 VSUBS 0.006586f
C952 B.n835 VSUBS 0.006586f
C953 B.n836 VSUBS 0.006586f
C954 B.n837 VSUBS 0.006586f
C955 B.n838 VSUBS 0.006586f
C956 B.n839 VSUBS 0.006586f
C957 B.n840 VSUBS 0.006586f
C958 B.n841 VSUBS 0.006586f
C959 B.n842 VSUBS 0.006586f
C960 B.n843 VSUBS 0.006586f
C961 B.n844 VSUBS 0.006586f
C962 B.n845 VSUBS 0.006586f
C963 B.n846 VSUBS 0.006586f
C964 B.n847 VSUBS 0.006586f
C965 B.n848 VSUBS 0.006586f
C966 B.n849 VSUBS 0.006586f
C967 B.n850 VSUBS 0.006586f
C968 B.n851 VSUBS 0.006586f
C969 B.n852 VSUBS 0.006586f
C970 B.n853 VSUBS 0.006586f
C971 B.n854 VSUBS 0.006586f
C972 B.n855 VSUBS 0.008595f
C973 B.n856 VSUBS 0.009156f
C974 B.n857 VSUBS 0.018207f
C975 VDD2.t1 VSUBS 0.370349f
C976 VDD2.t7 VSUBS 0.370349f
C977 VDD2.n0 VSUBS 3.10124f
C978 VDD2.t5 VSUBS 0.370349f
C979 VDD2.t6 VSUBS 0.370349f
C980 VDD2.n1 VSUBS 3.10124f
C981 VDD2.n2 VSUBS 3.75732f
C982 VDD2.t4 VSUBS 0.370349f
C983 VDD2.t0 VSUBS 0.370349f
C984 VDD2.n3 VSUBS 3.09257f
C985 VDD2.n4 VSUBS 3.43692f
C986 VDD2.t2 VSUBS 0.370349f
C987 VDD2.t3 VSUBS 0.370349f
C988 VDD2.n5 VSUBS 3.1012f
C989 VTAIL.t9 VSUBS 0.346162f
C990 VTAIL.t13 VSUBS 0.346162f
C991 VTAIL.n0 VSUBS 2.74185f
C992 VTAIL.n1 VSUBS 0.716672f
C993 VTAIL.n2 VSUBS 0.025512f
C994 VTAIL.n3 VSUBS 0.023128f
C995 VTAIL.n4 VSUBS 0.012428f
C996 VTAIL.n5 VSUBS 0.029376f
C997 VTAIL.n6 VSUBS 0.013159f
C998 VTAIL.n7 VSUBS 0.023128f
C999 VTAIL.n8 VSUBS 0.012428f
C1000 VTAIL.n9 VSUBS 0.029376f
C1001 VTAIL.n10 VSUBS 0.013159f
C1002 VTAIL.n11 VSUBS 0.023128f
C1003 VTAIL.n12 VSUBS 0.012428f
C1004 VTAIL.n13 VSUBS 0.029376f
C1005 VTAIL.n14 VSUBS 0.013159f
C1006 VTAIL.n15 VSUBS 0.023128f
C1007 VTAIL.n16 VSUBS 0.012428f
C1008 VTAIL.n17 VSUBS 0.029376f
C1009 VTAIL.n18 VSUBS 0.013159f
C1010 VTAIL.n19 VSUBS 0.023128f
C1011 VTAIL.n20 VSUBS 0.012428f
C1012 VTAIL.n21 VSUBS 0.029376f
C1013 VTAIL.n22 VSUBS 0.013159f
C1014 VTAIL.n23 VSUBS 0.023128f
C1015 VTAIL.n24 VSUBS 0.012428f
C1016 VTAIL.n25 VSUBS 0.029376f
C1017 VTAIL.n26 VSUBS 0.013159f
C1018 VTAIL.n27 VSUBS 0.023128f
C1019 VTAIL.n28 VSUBS 0.012428f
C1020 VTAIL.n29 VSUBS 0.029376f
C1021 VTAIL.n30 VSUBS 0.013159f
C1022 VTAIL.n31 VSUBS 0.023128f
C1023 VTAIL.n32 VSUBS 0.012428f
C1024 VTAIL.n33 VSUBS 0.029376f
C1025 VTAIL.n34 VSUBS 0.013159f
C1026 VTAIL.n35 VSUBS 0.189913f
C1027 VTAIL.t11 VSUBS 0.063114f
C1028 VTAIL.n36 VSUBS 0.022032f
C1029 VTAIL.n37 VSUBS 0.018687f
C1030 VTAIL.n38 VSUBS 0.012428f
C1031 VTAIL.n39 VSUBS 1.89048f
C1032 VTAIL.n40 VSUBS 0.023128f
C1033 VTAIL.n41 VSUBS 0.012428f
C1034 VTAIL.n42 VSUBS 0.013159f
C1035 VTAIL.n43 VSUBS 0.029376f
C1036 VTAIL.n44 VSUBS 0.029376f
C1037 VTAIL.n45 VSUBS 0.013159f
C1038 VTAIL.n46 VSUBS 0.012428f
C1039 VTAIL.n47 VSUBS 0.023128f
C1040 VTAIL.n48 VSUBS 0.023128f
C1041 VTAIL.n49 VSUBS 0.012428f
C1042 VTAIL.n50 VSUBS 0.013159f
C1043 VTAIL.n51 VSUBS 0.029376f
C1044 VTAIL.n52 VSUBS 0.029376f
C1045 VTAIL.n53 VSUBS 0.013159f
C1046 VTAIL.n54 VSUBS 0.012428f
C1047 VTAIL.n55 VSUBS 0.023128f
C1048 VTAIL.n56 VSUBS 0.023128f
C1049 VTAIL.n57 VSUBS 0.012428f
C1050 VTAIL.n58 VSUBS 0.013159f
C1051 VTAIL.n59 VSUBS 0.029376f
C1052 VTAIL.n60 VSUBS 0.029376f
C1053 VTAIL.n61 VSUBS 0.013159f
C1054 VTAIL.n62 VSUBS 0.012428f
C1055 VTAIL.n63 VSUBS 0.023128f
C1056 VTAIL.n64 VSUBS 0.023128f
C1057 VTAIL.n65 VSUBS 0.012428f
C1058 VTAIL.n66 VSUBS 0.013159f
C1059 VTAIL.n67 VSUBS 0.029376f
C1060 VTAIL.n68 VSUBS 0.029376f
C1061 VTAIL.n69 VSUBS 0.013159f
C1062 VTAIL.n70 VSUBS 0.012428f
C1063 VTAIL.n71 VSUBS 0.023128f
C1064 VTAIL.n72 VSUBS 0.023128f
C1065 VTAIL.n73 VSUBS 0.012428f
C1066 VTAIL.n74 VSUBS 0.013159f
C1067 VTAIL.n75 VSUBS 0.029376f
C1068 VTAIL.n76 VSUBS 0.029376f
C1069 VTAIL.n77 VSUBS 0.029376f
C1070 VTAIL.n78 VSUBS 0.013159f
C1071 VTAIL.n79 VSUBS 0.012428f
C1072 VTAIL.n80 VSUBS 0.023128f
C1073 VTAIL.n81 VSUBS 0.023128f
C1074 VTAIL.n82 VSUBS 0.012428f
C1075 VTAIL.n83 VSUBS 0.012794f
C1076 VTAIL.n84 VSUBS 0.012794f
C1077 VTAIL.n85 VSUBS 0.029376f
C1078 VTAIL.n86 VSUBS 0.029376f
C1079 VTAIL.n87 VSUBS 0.013159f
C1080 VTAIL.n88 VSUBS 0.012428f
C1081 VTAIL.n89 VSUBS 0.023128f
C1082 VTAIL.n90 VSUBS 0.023128f
C1083 VTAIL.n91 VSUBS 0.012428f
C1084 VTAIL.n92 VSUBS 0.013159f
C1085 VTAIL.n93 VSUBS 0.029376f
C1086 VTAIL.n94 VSUBS 0.029376f
C1087 VTAIL.n95 VSUBS 0.013159f
C1088 VTAIL.n96 VSUBS 0.012428f
C1089 VTAIL.n97 VSUBS 0.023128f
C1090 VTAIL.n98 VSUBS 0.023128f
C1091 VTAIL.n99 VSUBS 0.012428f
C1092 VTAIL.n100 VSUBS 0.013159f
C1093 VTAIL.n101 VSUBS 0.029376f
C1094 VTAIL.n102 VSUBS 0.071454f
C1095 VTAIL.n103 VSUBS 0.013159f
C1096 VTAIL.n104 VSUBS 0.012428f
C1097 VTAIL.n105 VSUBS 0.052828f
C1098 VTAIL.n106 VSUBS 0.035929f
C1099 VTAIL.n107 VSUBS 0.187399f
C1100 VTAIL.n108 VSUBS 0.025512f
C1101 VTAIL.n109 VSUBS 0.023128f
C1102 VTAIL.n110 VSUBS 0.012428f
C1103 VTAIL.n111 VSUBS 0.029376f
C1104 VTAIL.n112 VSUBS 0.013159f
C1105 VTAIL.n113 VSUBS 0.023128f
C1106 VTAIL.n114 VSUBS 0.012428f
C1107 VTAIL.n115 VSUBS 0.029376f
C1108 VTAIL.n116 VSUBS 0.013159f
C1109 VTAIL.n117 VSUBS 0.023128f
C1110 VTAIL.n118 VSUBS 0.012428f
C1111 VTAIL.n119 VSUBS 0.029376f
C1112 VTAIL.n120 VSUBS 0.013159f
C1113 VTAIL.n121 VSUBS 0.023128f
C1114 VTAIL.n122 VSUBS 0.012428f
C1115 VTAIL.n123 VSUBS 0.029376f
C1116 VTAIL.n124 VSUBS 0.013159f
C1117 VTAIL.n125 VSUBS 0.023128f
C1118 VTAIL.n126 VSUBS 0.012428f
C1119 VTAIL.n127 VSUBS 0.029376f
C1120 VTAIL.n128 VSUBS 0.013159f
C1121 VTAIL.n129 VSUBS 0.023128f
C1122 VTAIL.n130 VSUBS 0.012428f
C1123 VTAIL.n131 VSUBS 0.029376f
C1124 VTAIL.n132 VSUBS 0.013159f
C1125 VTAIL.n133 VSUBS 0.023128f
C1126 VTAIL.n134 VSUBS 0.012428f
C1127 VTAIL.n135 VSUBS 0.029376f
C1128 VTAIL.n136 VSUBS 0.013159f
C1129 VTAIL.n137 VSUBS 0.023128f
C1130 VTAIL.n138 VSUBS 0.012428f
C1131 VTAIL.n139 VSUBS 0.029376f
C1132 VTAIL.n140 VSUBS 0.013159f
C1133 VTAIL.n141 VSUBS 0.189913f
C1134 VTAIL.t2 VSUBS 0.063114f
C1135 VTAIL.n142 VSUBS 0.022032f
C1136 VTAIL.n143 VSUBS 0.018687f
C1137 VTAIL.n144 VSUBS 0.012428f
C1138 VTAIL.n145 VSUBS 1.89048f
C1139 VTAIL.n146 VSUBS 0.023128f
C1140 VTAIL.n147 VSUBS 0.012428f
C1141 VTAIL.n148 VSUBS 0.013159f
C1142 VTAIL.n149 VSUBS 0.029376f
C1143 VTAIL.n150 VSUBS 0.029376f
C1144 VTAIL.n151 VSUBS 0.013159f
C1145 VTAIL.n152 VSUBS 0.012428f
C1146 VTAIL.n153 VSUBS 0.023128f
C1147 VTAIL.n154 VSUBS 0.023128f
C1148 VTAIL.n155 VSUBS 0.012428f
C1149 VTAIL.n156 VSUBS 0.013159f
C1150 VTAIL.n157 VSUBS 0.029376f
C1151 VTAIL.n158 VSUBS 0.029376f
C1152 VTAIL.n159 VSUBS 0.013159f
C1153 VTAIL.n160 VSUBS 0.012428f
C1154 VTAIL.n161 VSUBS 0.023128f
C1155 VTAIL.n162 VSUBS 0.023128f
C1156 VTAIL.n163 VSUBS 0.012428f
C1157 VTAIL.n164 VSUBS 0.013159f
C1158 VTAIL.n165 VSUBS 0.029376f
C1159 VTAIL.n166 VSUBS 0.029376f
C1160 VTAIL.n167 VSUBS 0.013159f
C1161 VTAIL.n168 VSUBS 0.012428f
C1162 VTAIL.n169 VSUBS 0.023128f
C1163 VTAIL.n170 VSUBS 0.023128f
C1164 VTAIL.n171 VSUBS 0.012428f
C1165 VTAIL.n172 VSUBS 0.013159f
C1166 VTAIL.n173 VSUBS 0.029376f
C1167 VTAIL.n174 VSUBS 0.029376f
C1168 VTAIL.n175 VSUBS 0.013159f
C1169 VTAIL.n176 VSUBS 0.012428f
C1170 VTAIL.n177 VSUBS 0.023128f
C1171 VTAIL.n178 VSUBS 0.023128f
C1172 VTAIL.n179 VSUBS 0.012428f
C1173 VTAIL.n180 VSUBS 0.013159f
C1174 VTAIL.n181 VSUBS 0.029376f
C1175 VTAIL.n182 VSUBS 0.029376f
C1176 VTAIL.n183 VSUBS 0.029376f
C1177 VTAIL.n184 VSUBS 0.013159f
C1178 VTAIL.n185 VSUBS 0.012428f
C1179 VTAIL.n186 VSUBS 0.023128f
C1180 VTAIL.n187 VSUBS 0.023128f
C1181 VTAIL.n188 VSUBS 0.012428f
C1182 VTAIL.n189 VSUBS 0.012794f
C1183 VTAIL.n190 VSUBS 0.012794f
C1184 VTAIL.n191 VSUBS 0.029376f
C1185 VTAIL.n192 VSUBS 0.029376f
C1186 VTAIL.n193 VSUBS 0.013159f
C1187 VTAIL.n194 VSUBS 0.012428f
C1188 VTAIL.n195 VSUBS 0.023128f
C1189 VTAIL.n196 VSUBS 0.023128f
C1190 VTAIL.n197 VSUBS 0.012428f
C1191 VTAIL.n198 VSUBS 0.013159f
C1192 VTAIL.n199 VSUBS 0.029376f
C1193 VTAIL.n200 VSUBS 0.029376f
C1194 VTAIL.n201 VSUBS 0.013159f
C1195 VTAIL.n202 VSUBS 0.012428f
C1196 VTAIL.n203 VSUBS 0.023128f
C1197 VTAIL.n204 VSUBS 0.023128f
C1198 VTAIL.n205 VSUBS 0.012428f
C1199 VTAIL.n206 VSUBS 0.013159f
C1200 VTAIL.n207 VSUBS 0.029376f
C1201 VTAIL.n208 VSUBS 0.071454f
C1202 VTAIL.n209 VSUBS 0.013159f
C1203 VTAIL.n210 VSUBS 0.012428f
C1204 VTAIL.n211 VSUBS 0.052828f
C1205 VTAIL.n212 VSUBS 0.035929f
C1206 VTAIL.n213 VSUBS 0.187399f
C1207 VTAIL.t3 VSUBS 0.346162f
C1208 VTAIL.t6 VSUBS 0.346162f
C1209 VTAIL.n214 VSUBS 2.74185f
C1210 VTAIL.n215 VSUBS 0.845324f
C1211 VTAIL.n216 VSUBS 0.025512f
C1212 VTAIL.n217 VSUBS 0.023128f
C1213 VTAIL.n218 VSUBS 0.012428f
C1214 VTAIL.n219 VSUBS 0.029376f
C1215 VTAIL.n220 VSUBS 0.013159f
C1216 VTAIL.n221 VSUBS 0.023128f
C1217 VTAIL.n222 VSUBS 0.012428f
C1218 VTAIL.n223 VSUBS 0.029376f
C1219 VTAIL.n224 VSUBS 0.013159f
C1220 VTAIL.n225 VSUBS 0.023128f
C1221 VTAIL.n226 VSUBS 0.012428f
C1222 VTAIL.n227 VSUBS 0.029376f
C1223 VTAIL.n228 VSUBS 0.013159f
C1224 VTAIL.n229 VSUBS 0.023128f
C1225 VTAIL.n230 VSUBS 0.012428f
C1226 VTAIL.n231 VSUBS 0.029376f
C1227 VTAIL.n232 VSUBS 0.013159f
C1228 VTAIL.n233 VSUBS 0.023128f
C1229 VTAIL.n234 VSUBS 0.012428f
C1230 VTAIL.n235 VSUBS 0.029376f
C1231 VTAIL.n236 VSUBS 0.013159f
C1232 VTAIL.n237 VSUBS 0.023128f
C1233 VTAIL.n238 VSUBS 0.012428f
C1234 VTAIL.n239 VSUBS 0.029376f
C1235 VTAIL.n240 VSUBS 0.013159f
C1236 VTAIL.n241 VSUBS 0.023128f
C1237 VTAIL.n242 VSUBS 0.012428f
C1238 VTAIL.n243 VSUBS 0.029376f
C1239 VTAIL.n244 VSUBS 0.013159f
C1240 VTAIL.n245 VSUBS 0.023128f
C1241 VTAIL.n246 VSUBS 0.012428f
C1242 VTAIL.n247 VSUBS 0.029376f
C1243 VTAIL.n248 VSUBS 0.013159f
C1244 VTAIL.n249 VSUBS 0.189913f
C1245 VTAIL.t1 VSUBS 0.063114f
C1246 VTAIL.n250 VSUBS 0.022032f
C1247 VTAIL.n251 VSUBS 0.018687f
C1248 VTAIL.n252 VSUBS 0.012428f
C1249 VTAIL.n253 VSUBS 1.89048f
C1250 VTAIL.n254 VSUBS 0.023128f
C1251 VTAIL.n255 VSUBS 0.012428f
C1252 VTAIL.n256 VSUBS 0.013159f
C1253 VTAIL.n257 VSUBS 0.029376f
C1254 VTAIL.n258 VSUBS 0.029376f
C1255 VTAIL.n259 VSUBS 0.013159f
C1256 VTAIL.n260 VSUBS 0.012428f
C1257 VTAIL.n261 VSUBS 0.023128f
C1258 VTAIL.n262 VSUBS 0.023128f
C1259 VTAIL.n263 VSUBS 0.012428f
C1260 VTAIL.n264 VSUBS 0.013159f
C1261 VTAIL.n265 VSUBS 0.029376f
C1262 VTAIL.n266 VSUBS 0.029376f
C1263 VTAIL.n267 VSUBS 0.013159f
C1264 VTAIL.n268 VSUBS 0.012428f
C1265 VTAIL.n269 VSUBS 0.023128f
C1266 VTAIL.n270 VSUBS 0.023128f
C1267 VTAIL.n271 VSUBS 0.012428f
C1268 VTAIL.n272 VSUBS 0.013159f
C1269 VTAIL.n273 VSUBS 0.029376f
C1270 VTAIL.n274 VSUBS 0.029376f
C1271 VTAIL.n275 VSUBS 0.013159f
C1272 VTAIL.n276 VSUBS 0.012428f
C1273 VTAIL.n277 VSUBS 0.023128f
C1274 VTAIL.n278 VSUBS 0.023128f
C1275 VTAIL.n279 VSUBS 0.012428f
C1276 VTAIL.n280 VSUBS 0.013159f
C1277 VTAIL.n281 VSUBS 0.029376f
C1278 VTAIL.n282 VSUBS 0.029376f
C1279 VTAIL.n283 VSUBS 0.013159f
C1280 VTAIL.n284 VSUBS 0.012428f
C1281 VTAIL.n285 VSUBS 0.023128f
C1282 VTAIL.n286 VSUBS 0.023128f
C1283 VTAIL.n287 VSUBS 0.012428f
C1284 VTAIL.n288 VSUBS 0.013159f
C1285 VTAIL.n289 VSUBS 0.029376f
C1286 VTAIL.n290 VSUBS 0.029376f
C1287 VTAIL.n291 VSUBS 0.029376f
C1288 VTAIL.n292 VSUBS 0.013159f
C1289 VTAIL.n293 VSUBS 0.012428f
C1290 VTAIL.n294 VSUBS 0.023128f
C1291 VTAIL.n295 VSUBS 0.023128f
C1292 VTAIL.n296 VSUBS 0.012428f
C1293 VTAIL.n297 VSUBS 0.012794f
C1294 VTAIL.n298 VSUBS 0.012794f
C1295 VTAIL.n299 VSUBS 0.029376f
C1296 VTAIL.n300 VSUBS 0.029376f
C1297 VTAIL.n301 VSUBS 0.013159f
C1298 VTAIL.n302 VSUBS 0.012428f
C1299 VTAIL.n303 VSUBS 0.023128f
C1300 VTAIL.n304 VSUBS 0.023128f
C1301 VTAIL.n305 VSUBS 0.012428f
C1302 VTAIL.n306 VSUBS 0.013159f
C1303 VTAIL.n307 VSUBS 0.029376f
C1304 VTAIL.n308 VSUBS 0.029376f
C1305 VTAIL.n309 VSUBS 0.013159f
C1306 VTAIL.n310 VSUBS 0.012428f
C1307 VTAIL.n311 VSUBS 0.023128f
C1308 VTAIL.n312 VSUBS 0.023128f
C1309 VTAIL.n313 VSUBS 0.012428f
C1310 VTAIL.n314 VSUBS 0.013159f
C1311 VTAIL.n315 VSUBS 0.029376f
C1312 VTAIL.n316 VSUBS 0.071454f
C1313 VTAIL.n317 VSUBS 0.013159f
C1314 VTAIL.n318 VSUBS 0.012428f
C1315 VTAIL.n319 VSUBS 0.052828f
C1316 VTAIL.n320 VSUBS 0.035929f
C1317 VTAIL.n321 VSUBS 1.81636f
C1318 VTAIL.n322 VSUBS 0.025512f
C1319 VTAIL.n323 VSUBS 0.023128f
C1320 VTAIL.n324 VSUBS 0.012428f
C1321 VTAIL.n325 VSUBS 0.029376f
C1322 VTAIL.n326 VSUBS 0.013159f
C1323 VTAIL.n327 VSUBS 0.023128f
C1324 VTAIL.n328 VSUBS 0.012428f
C1325 VTAIL.n329 VSUBS 0.029376f
C1326 VTAIL.n330 VSUBS 0.013159f
C1327 VTAIL.n331 VSUBS 0.023128f
C1328 VTAIL.n332 VSUBS 0.012428f
C1329 VTAIL.n333 VSUBS 0.029376f
C1330 VTAIL.n334 VSUBS 0.013159f
C1331 VTAIL.n335 VSUBS 0.023128f
C1332 VTAIL.n336 VSUBS 0.012428f
C1333 VTAIL.n337 VSUBS 0.029376f
C1334 VTAIL.n338 VSUBS 0.029376f
C1335 VTAIL.n339 VSUBS 0.013159f
C1336 VTAIL.n340 VSUBS 0.023128f
C1337 VTAIL.n341 VSUBS 0.012428f
C1338 VTAIL.n342 VSUBS 0.029376f
C1339 VTAIL.n343 VSUBS 0.013159f
C1340 VTAIL.n344 VSUBS 0.023128f
C1341 VTAIL.n345 VSUBS 0.012428f
C1342 VTAIL.n346 VSUBS 0.029376f
C1343 VTAIL.n347 VSUBS 0.013159f
C1344 VTAIL.n348 VSUBS 0.023128f
C1345 VTAIL.n349 VSUBS 0.012428f
C1346 VTAIL.n350 VSUBS 0.029376f
C1347 VTAIL.n351 VSUBS 0.013159f
C1348 VTAIL.n352 VSUBS 0.023128f
C1349 VTAIL.n353 VSUBS 0.012428f
C1350 VTAIL.n354 VSUBS 0.029376f
C1351 VTAIL.n355 VSUBS 0.013159f
C1352 VTAIL.n356 VSUBS 0.189913f
C1353 VTAIL.t15 VSUBS 0.063114f
C1354 VTAIL.n357 VSUBS 0.022032f
C1355 VTAIL.n358 VSUBS 0.018687f
C1356 VTAIL.n359 VSUBS 0.012428f
C1357 VTAIL.n360 VSUBS 1.89048f
C1358 VTAIL.n361 VSUBS 0.023128f
C1359 VTAIL.n362 VSUBS 0.012428f
C1360 VTAIL.n363 VSUBS 0.013159f
C1361 VTAIL.n364 VSUBS 0.029376f
C1362 VTAIL.n365 VSUBS 0.029376f
C1363 VTAIL.n366 VSUBS 0.013159f
C1364 VTAIL.n367 VSUBS 0.012428f
C1365 VTAIL.n368 VSUBS 0.023128f
C1366 VTAIL.n369 VSUBS 0.023128f
C1367 VTAIL.n370 VSUBS 0.012428f
C1368 VTAIL.n371 VSUBS 0.013159f
C1369 VTAIL.n372 VSUBS 0.029376f
C1370 VTAIL.n373 VSUBS 0.029376f
C1371 VTAIL.n374 VSUBS 0.013159f
C1372 VTAIL.n375 VSUBS 0.012428f
C1373 VTAIL.n376 VSUBS 0.023128f
C1374 VTAIL.n377 VSUBS 0.023128f
C1375 VTAIL.n378 VSUBS 0.012428f
C1376 VTAIL.n379 VSUBS 0.013159f
C1377 VTAIL.n380 VSUBS 0.029376f
C1378 VTAIL.n381 VSUBS 0.029376f
C1379 VTAIL.n382 VSUBS 0.013159f
C1380 VTAIL.n383 VSUBS 0.012428f
C1381 VTAIL.n384 VSUBS 0.023128f
C1382 VTAIL.n385 VSUBS 0.023128f
C1383 VTAIL.n386 VSUBS 0.012428f
C1384 VTAIL.n387 VSUBS 0.013159f
C1385 VTAIL.n388 VSUBS 0.029376f
C1386 VTAIL.n389 VSUBS 0.029376f
C1387 VTAIL.n390 VSUBS 0.013159f
C1388 VTAIL.n391 VSUBS 0.012428f
C1389 VTAIL.n392 VSUBS 0.023128f
C1390 VTAIL.n393 VSUBS 0.023128f
C1391 VTAIL.n394 VSUBS 0.012428f
C1392 VTAIL.n395 VSUBS 0.013159f
C1393 VTAIL.n396 VSUBS 0.029376f
C1394 VTAIL.n397 VSUBS 0.029376f
C1395 VTAIL.n398 VSUBS 0.013159f
C1396 VTAIL.n399 VSUBS 0.012428f
C1397 VTAIL.n400 VSUBS 0.023128f
C1398 VTAIL.n401 VSUBS 0.023128f
C1399 VTAIL.n402 VSUBS 0.012428f
C1400 VTAIL.n403 VSUBS 0.012794f
C1401 VTAIL.n404 VSUBS 0.012794f
C1402 VTAIL.n405 VSUBS 0.029376f
C1403 VTAIL.n406 VSUBS 0.029376f
C1404 VTAIL.n407 VSUBS 0.013159f
C1405 VTAIL.n408 VSUBS 0.012428f
C1406 VTAIL.n409 VSUBS 0.023128f
C1407 VTAIL.n410 VSUBS 0.023128f
C1408 VTAIL.n411 VSUBS 0.012428f
C1409 VTAIL.n412 VSUBS 0.013159f
C1410 VTAIL.n413 VSUBS 0.029376f
C1411 VTAIL.n414 VSUBS 0.029376f
C1412 VTAIL.n415 VSUBS 0.013159f
C1413 VTAIL.n416 VSUBS 0.012428f
C1414 VTAIL.n417 VSUBS 0.023128f
C1415 VTAIL.n418 VSUBS 0.023128f
C1416 VTAIL.n419 VSUBS 0.012428f
C1417 VTAIL.n420 VSUBS 0.013159f
C1418 VTAIL.n421 VSUBS 0.029376f
C1419 VTAIL.n422 VSUBS 0.071454f
C1420 VTAIL.n423 VSUBS 0.013159f
C1421 VTAIL.n424 VSUBS 0.012428f
C1422 VTAIL.n425 VSUBS 0.052828f
C1423 VTAIL.n426 VSUBS 0.035929f
C1424 VTAIL.n427 VSUBS 1.81636f
C1425 VTAIL.t12 VSUBS 0.346162f
C1426 VTAIL.t8 VSUBS 0.346162f
C1427 VTAIL.n428 VSUBS 2.74186f
C1428 VTAIL.n429 VSUBS 0.845314f
C1429 VTAIL.n430 VSUBS 0.025512f
C1430 VTAIL.n431 VSUBS 0.023128f
C1431 VTAIL.n432 VSUBS 0.012428f
C1432 VTAIL.n433 VSUBS 0.029376f
C1433 VTAIL.n434 VSUBS 0.013159f
C1434 VTAIL.n435 VSUBS 0.023128f
C1435 VTAIL.n436 VSUBS 0.012428f
C1436 VTAIL.n437 VSUBS 0.029376f
C1437 VTAIL.n438 VSUBS 0.013159f
C1438 VTAIL.n439 VSUBS 0.023128f
C1439 VTAIL.n440 VSUBS 0.012428f
C1440 VTAIL.n441 VSUBS 0.029376f
C1441 VTAIL.n442 VSUBS 0.013159f
C1442 VTAIL.n443 VSUBS 0.023128f
C1443 VTAIL.n444 VSUBS 0.012428f
C1444 VTAIL.n445 VSUBS 0.029376f
C1445 VTAIL.n446 VSUBS 0.029376f
C1446 VTAIL.n447 VSUBS 0.013159f
C1447 VTAIL.n448 VSUBS 0.023128f
C1448 VTAIL.n449 VSUBS 0.012428f
C1449 VTAIL.n450 VSUBS 0.029376f
C1450 VTAIL.n451 VSUBS 0.013159f
C1451 VTAIL.n452 VSUBS 0.023128f
C1452 VTAIL.n453 VSUBS 0.012428f
C1453 VTAIL.n454 VSUBS 0.029376f
C1454 VTAIL.n455 VSUBS 0.013159f
C1455 VTAIL.n456 VSUBS 0.023128f
C1456 VTAIL.n457 VSUBS 0.012428f
C1457 VTAIL.n458 VSUBS 0.029376f
C1458 VTAIL.n459 VSUBS 0.013159f
C1459 VTAIL.n460 VSUBS 0.023128f
C1460 VTAIL.n461 VSUBS 0.012428f
C1461 VTAIL.n462 VSUBS 0.029376f
C1462 VTAIL.n463 VSUBS 0.013159f
C1463 VTAIL.n464 VSUBS 0.189913f
C1464 VTAIL.t14 VSUBS 0.063114f
C1465 VTAIL.n465 VSUBS 0.022032f
C1466 VTAIL.n466 VSUBS 0.018687f
C1467 VTAIL.n467 VSUBS 0.012428f
C1468 VTAIL.n468 VSUBS 1.89048f
C1469 VTAIL.n469 VSUBS 0.023128f
C1470 VTAIL.n470 VSUBS 0.012428f
C1471 VTAIL.n471 VSUBS 0.013159f
C1472 VTAIL.n472 VSUBS 0.029376f
C1473 VTAIL.n473 VSUBS 0.029376f
C1474 VTAIL.n474 VSUBS 0.013159f
C1475 VTAIL.n475 VSUBS 0.012428f
C1476 VTAIL.n476 VSUBS 0.023128f
C1477 VTAIL.n477 VSUBS 0.023128f
C1478 VTAIL.n478 VSUBS 0.012428f
C1479 VTAIL.n479 VSUBS 0.013159f
C1480 VTAIL.n480 VSUBS 0.029376f
C1481 VTAIL.n481 VSUBS 0.029376f
C1482 VTAIL.n482 VSUBS 0.013159f
C1483 VTAIL.n483 VSUBS 0.012428f
C1484 VTAIL.n484 VSUBS 0.023128f
C1485 VTAIL.n485 VSUBS 0.023128f
C1486 VTAIL.n486 VSUBS 0.012428f
C1487 VTAIL.n487 VSUBS 0.013159f
C1488 VTAIL.n488 VSUBS 0.029376f
C1489 VTAIL.n489 VSUBS 0.029376f
C1490 VTAIL.n490 VSUBS 0.013159f
C1491 VTAIL.n491 VSUBS 0.012428f
C1492 VTAIL.n492 VSUBS 0.023128f
C1493 VTAIL.n493 VSUBS 0.023128f
C1494 VTAIL.n494 VSUBS 0.012428f
C1495 VTAIL.n495 VSUBS 0.013159f
C1496 VTAIL.n496 VSUBS 0.029376f
C1497 VTAIL.n497 VSUBS 0.029376f
C1498 VTAIL.n498 VSUBS 0.013159f
C1499 VTAIL.n499 VSUBS 0.012428f
C1500 VTAIL.n500 VSUBS 0.023128f
C1501 VTAIL.n501 VSUBS 0.023128f
C1502 VTAIL.n502 VSUBS 0.012428f
C1503 VTAIL.n503 VSUBS 0.013159f
C1504 VTAIL.n504 VSUBS 0.029376f
C1505 VTAIL.n505 VSUBS 0.029376f
C1506 VTAIL.n506 VSUBS 0.013159f
C1507 VTAIL.n507 VSUBS 0.012428f
C1508 VTAIL.n508 VSUBS 0.023128f
C1509 VTAIL.n509 VSUBS 0.023128f
C1510 VTAIL.n510 VSUBS 0.012428f
C1511 VTAIL.n511 VSUBS 0.012794f
C1512 VTAIL.n512 VSUBS 0.012794f
C1513 VTAIL.n513 VSUBS 0.029376f
C1514 VTAIL.n514 VSUBS 0.029376f
C1515 VTAIL.n515 VSUBS 0.013159f
C1516 VTAIL.n516 VSUBS 0.012428f
C1517 VTAIL.n517 VSUBS 0.023128f
C1518 VTAIL.n518 VSUBS 0.023128f
C1519 VTAIL.n519 VSUBS 0.012428f
C1520 VTAIL.n520 VSUBS 0.013159f
C1521 VTAIL.n521 VSUBS 0.029376f
C1522 VTAIL.n522 VSUBS 0.029376f
C1523 VTAIL.n523 VSUBS 0.013159f
C1524 VTAIL.n524 VSUBS 0.012428f
C1525 VTAIL.n525 VSUBS 0.023128f
C1526 VTAIL.n526 VSUBS 0.023128f
C1527 VTAIL.n527 VSUBS 0.012428f
C1528 VTAIL.n528 VSUBS 0.013159f
C1529 VTAIL.n529 VSUBS 0.029376f
C1530 VTAIL.n530 VSUBS 0.071454f
C1531 VTAIL.n531 VSUBS 0.013159f
C1532 VTAIL.n532 VSUBS 0.012428f
C1533 VTAIL.n533 VSUBS 0.052828f
C1534 VTAIL.n534 VSUBS 0.035929f
C1535 VTAIL.n535 VSUBS 0.187399f
C1536 VTAIL.n536 VSUBS 0.025512f
C1537 VTAIL.n537 VSUBS 0.023128f
C1538 VTAIL.n538 VSUBS 0.012428f
C1539 VTAIL.n539 VSUBS 0.029376f
C1540 VTAIL.n540 VSUBS 0.013159f
C1541 VTAIL.n541 VSUBS 0.023128f
C1542 VTAIL.n542 VSUBS 0.012428f
C1543 VTAIL.n543 VSUBS 0.029376f
C1544 VTAIL.n544 VSUBS 0.013159f
C1545 VTAIL.n545 VSUBS 0.023128f
C1546 VTAIL.n546 VSUBS 0.012428f
C1547 VTAIL.n547 VSUBS 0.029376f
C1548 VTAIL.n548 VSUBS 0.013159f
C1549 VTAIL.n549 VSUBS 0.023128f
C1550 VTAIL.n550 VSUBS 0.012428f
C1551 VTAIL.n551 VSUBS 0.029376f
C1552 VTAIL.n552 VSUBS 0.029376f
C1553 VTAIL.n553 VSUBS 0.013159f
C1554 VTAIL.n554 VSUBS 0.023128f
C1555 VTAIL.n555 VSUBS 0.012428f
C1556 VTAIL.n556 VSUBS 0.029376f
C1557 VTAIL.n557 VSUBS 0.013159f
C1558 VTAIL.n558 VSUBS 0.023128f
C1559 VTAIL.n559 VSUBS 0.012428f
C1560 VTAIL.n560 VSUBS 0.029376f
C1561 VTAIL.n561 VSUBS 0.013159f
C1562 VTAIL.n562 VSUBS 0.023128f
C1563 VTAIL.n563 VSUBS 0.012428f
C1564 VTAIL.n564 VSUBS 0.029376f
C1565 VTAIL.n565 VSUBS 0.013159f
C1566 VTAIL.n566 VSUBS 0.023128f
C1567 VTAIL.n567 VSUBS 0.012428f
C1568 VTAIL.n568 VSUBS 0.029376f
C1569 VTAIL.n569 VSUBS 0.013159f
C1570 VTAIL.n570 VSUBS 0.189913f
C1571 VTAIL.t4 VSUBS 0.063114f
C1572 VTAIL.n571 VSUBS 0.022032f
C1573 VTAIL.n572 VSUBS 0.018687f
C1574 VTAIL.n573 VSUBS 0.012428f
C1575 VTAIL.n574 VSUBS 1.89048f
C1576 VTAIL.n575 VSUBS 0.023128f
C1577 VTAIL.n576 VSUBS 0.012428f
C1578 VTAIL.n577 VSUBS 0.013159f
C1579 VTAIL.n578 VSUBS 0.029376f
C1580 VTAIL.n579 VSUBS 0.029376f
C1581 VTAIL.n580 VSUBS 0.013159f
C1582 VTAIL.n581 VSUBS 0.012428f
C1583 VTAIL.n582 VSUBS 0.023128f
C1584 VTAIL.n583 VSUBS 0.023128f
C1585 VTAIL.n584 VSUBS 0.012428f
C1586 VTAIL.n585 VSUBS 0.013159f
C1587 VTAIL.n586 VSUBS 0.029376f
C1588 VTAIL.n587 VSUBS 0.029376f
C1589 VTAIL.n588 VSUBS 0.013159f
C1590 VTAIL.n589 VSUBS 0.012428f
C1591 VTAIL.n590 VSUBS 0.023128f
C1592 VTAIL.n591 VSUBS 0.023128f
C1593 VTAIL.n592 VSUBS 0.012428f
C1594 VTAIL.n593 VSUBS 0.013159f
C1595 VTAIL.n594 VSUBS 0.029376f
C1596 VTAIL.n595 VSUBS 0.029376f
C1597 VTAIL.n596 VSUBS 0.013159f
C1598 VTAIL.n597 VSUBS 0.012428f
C1599 VTAIL.n598 VSUBS 0.023128f
C1600 VTAIL.n599 VSUBS 0.023128f
C1601 VTAIL.n600 VSUBS 0.012428f
C1602 VTAIL.n601 VSUBS 0.013159f
C1603 VTAIL.n602 VSUBS 0.029376f
C1604 VTAIL.n603 VSUBS 0.029376f
C1605 VTAIL.n604 VSUBS 0.013159f
C1606 VTAIL.n605 VSUBS 0.012428f
C1607 VTAIL.n606 VSUBS 0.023128f
C1608 VTAIL.n607 VSUBS 0.023128f
C1609 VTAIL.n608 VSUBS 0.012428f
C1610 VTAIL.n609 VSUBS 0.013159f
C1611 VTAIL.n610 VSUBS 0.029376f
C1612 VTAIL.n611 VSUBS 0.029376f
C1613 VTAIL.n612 VSUBS 0.013159f
C1614 VTAIL.n613 VSUBS 0.012428f
C1615 VTAIL.n614 VSUBS 0.023128f
C1616 VTAIL.n615 VSUBS 0.023128f
C1617 VTAIL.n616 VSUBS 0.012428f
C1618 VTAIL.n617 VSUBS 0.012794f
C1619 VTAIL.n618 VSUBS 0.012794f
C1620 VTAIL.n619 VSUBS 0.029376f
C1621 VTAIL.n620 VSUBS 0.029376f
C1622 VTAIL.n621 VSUBS 0.013159f
C1623 VTAIL.n622 VSUBS 0.012428f
C1624 VTAIL.n623 VSUBS 0.023128f
C1625 VTAIL.n624 VSUBS 0.023128f
C1626 VTAIL.n625 VSUBS 0.012428f
C1627 VTAIL.n626 VSUBS 0.013159f
C1628 VTAIL.n627 VSUBS 0.029376f
C1629 VTAIL.n628 VSUBS 0.029376f
C1630 VTAIL.n629 VSUBS 0.013159f
C1631 VTAIL.n630 VSUBS 0.012428f
C1632 VTAIL.n631 VSUBS 0.023128f
C1633 VTAIL.n632 VSUBS 0.023128f
C1634 VTAIL.n633 VSUBS 0.012428f
C1635 VTAIL.n634 VSUBS 0.013159f
C1636 VTAIL.n635 VSUBS 0.029376f
C1637 VTAIL.n636 VSUBS 0.071454f
C1638 VTAIL.n637 VSUBS 0.013159f
C1639 VTAIL.n638 VSUBS 0.012428f
C1640 VTAIL.n639 VSUBS 0.052828f
C1641 VTAIL.n640 VSUBS 0.035929f
C1642 VTAIL.n641 VSUBS 0.187399f
C1643 VTAIL.t0 VSUBS 0.346162f
C1644 VTAIL.t5 VSUBS 0.346162f
C1645 VTAIL.n642 VSUBS 2.74186f
C1646 VTAIL.n643 VSUBS 0.845314f
C1647 VTAIL.n644 VSUBS 0.025512f
C1648 VTAIL.n645 VSUBS 0.023128f
C1649 VTAIL.n646 VSUBS 0.012428f
C1650 VTAIL.n647 VSUBS 0.029376f
C1651 VTAIL.n648 VSUBS 0.013159f
C1652 VTAIL.n649 VSUBS 0.023128f
C1653 VTAIL.n650 VSUBS 0.012428f
C1654 VTAIL.n651 VSUBS 0.029376f
C1655 VTAIL.n652 VSUBS 0.013159f
C1656 VTAIL.n653 VSUBS 0.023128f
C1657 VTAIL.n654 VSUBS 0.012428f
C1658 VTAIL.n655 VSUBS 0.029376f
C1659 VTAIL.n656 VSUBS 0.013159f
C1660 VTAIL.n657 VSUBS 0.023128f
C1661 VTAIL.n658 VSUBS 0.012428f
C1662 VTAIL.n659 VSUBS 0.029376f
C1663 VTAIL.n660 VSUBS 0.029376f
C1664 VTAIL.n661 VSUBS 0.013159f
C1665 VTAIL.n662 VSUBS 0.023128f
C1666 VTAIL.n663 VSUBS 0.012428f
C1667 VTAIL.n664 VSUBS 0.029376f
C1668 VTAIL.n665 VSUBS 0.013159f
C1669 VTAIL.n666 VSUBS 0.023128f
C1670 VTAIL.n667 VSUBS 0.012428f
C1671 VTAIL.n668 VSUBS 0.029376f
C1672 VTAIL.n669 VSUBS 0.013159f
C1673 VTAIL.n670 VSUBS 0.023128f
C1674 VTAIL.n671 VSUBS 0.012428f
C1675 VTAIL.n672 VSUBS 0.029376f
C1676 VTAIL.n673 VSUBS 0.013159f
C1677 VTAIL.n674 VSUBS 0.023128f
C1678 VTAIL.n675 VSUBS 0.012428f
C1679 VTAIL.n676 VSUBS 0.029376f
C1680 VTAIL.n677 VSUBS 0.013159f
C1681 VTAIL.n678 VSUBS 0.189913f
C1682 VTAIL.t7 VSUBS 0.063114f
C1683 VTAIL.n679 VSUBS 0.022032f
C1684 VTAIL.n680 VSUBS 0.018687f
C1685 VTAIL.n681 VSUBS 0.012428f
C1686 VTAIL.n682 VSUBS 1.89048f
C1687 VTAIL.n683 VSUBS 0.023128f
C1688 VTAIL.n684 VSUBS 0.012428f
C1689 VTAIL.n685 VSUBS 0.013159f
C1690 VTAIL.n686 VSUBS 0.029376f
C1691 VTAIL.n687 VSUBS 0.029376f
C1692 VTAIL.n688 VSUBS 0.013159f
C1693 VTAIL.n689 VSUBS 0.012428f
C1694 VTAIL.n690 VSUBS 0.023128f
C1695 VTAIL.n691 VSUBS 0.023128f
C1696 VTAIL.n692 VSUBS 0.012428f
C1697 VTAIL.n693 VSUBS 0.013159f
C1698 VTAIL.n694 VSUBS 0.029376f
C1699 VTAIL.n695 VSUBS 0.029376f
C1700 VTAIL.n696 VSUBS 0.013159f
C1701 VTAIL.n697 VSUBS 0.012428f
C1702 VTAIL.n698 VSUBS 0.023128f
C1703 VTAIL.n699 VSUBS 0.023128f
C1704 VTAIL.n700 VSUBS 0.012428f
C1705 VTAIL.n701 VSUBS 0.013159f
C1706 VTAIL.n702 VSUBS 0.029376f
C1707 VTAIL.n703 VSUBS 0.029376f
C1708 VTAIL.n704 VSUBS 0.013159f
C1709 VTAIL.n705 VSUBS 0.012428f
C1710 VTAIL.n706 VSUBS 0.023128f
C1711 VTAIL.n707 VSUBS 0.023128f
C1712 VTAIL.n708 VSUBS 0.012428f
C1713 VTAIL.n709 VSUBS 0.013159f
C1714 VTAIL.n710 VSUBS 0.029376f
C1715 VTAIL.n711 VSUBS 0.029376f
C1716 VTAIL.n712 VSUBS 0.013159f
C1717 VTAIL.n713 VSUBS 0.012428f
C1718 VTAIL.n714 VSUBS 0.023128f
C1719 VTAIL.n715 VSUBS 0.023128f
C1720 VTAIL.n716 VSUBS 0.012428f
C1721 VTAIL.n717 VSUBS 0.013159f
C1722 VTAIL.n718 VSUBS 0.029376f
C1723 VTAIL.n719 VSUBS 0.029376f
C1724 VTAIL.n720 VSUBS 0.013159f
C1725 VTAIL.n721 VSUBS 0.012428f
C1726 VTAIL.n722 VSUBS 0.023128f
C1727 VTAIL.n723 VSUBS 0.023128f
C1728 VTAIL.n724 VSUBS 0.012428f
C1729 VTAIL.n725 VSUBS 0.012794f
C1730 VTAIL.n726 VSUBS 0.012794f
C1731 VTAIL.n727 VSUBS 0.029376f
C1732 VTAIL.n728 VSUBS 0.029376f
C1733 VTAIL.n729 VSUBS 0.013159f
C1734 VTAIL.n730 VSUBS 0.012428f
C1735 VTAIL.n731 VSUBS 0.023128f
C1736 VTAIL.n732 VSUBS 0.023128f
C1737 VTAIL.n733 VSUBS 0.012428f
C1738 VTAIL.n734 VSUBS 0.013159f
C1739 VTAIL.n735 VSUBS 0.029376f
C1740 VTAIL.n736 VSUBS 0.029376f
C1741 VTAIL.n737 VSUBS 0.013159f
C1742 VTAIL.n738 VSUBS 0.012428f
C1743 VTAIL.n739 VSUBS 0.023128f
C1744 VTAIL.n740 VSUBS 0.023128f
C1745 VTAIL.n741 VSUBS 0.012428f
C1746 VTAIL.n742 VSUBS 0.013159f
C1747 VTAIL.n743 VSUBS 0.029376f
C1748 VTAIL.n744 VSUBS 0.071454f
C1749 VTAIL.n745 VSUBS 0.013159f
C1750 VTAIL.n746 VSUBS 0.012428f
C1751 VTAIL.n747 VSUBS 0.052828f
C1752 VTAIL.n748 VSUBS 0.035929f
C1753 VTAIL.n749 VSUBS 1.81636f
C1754 VTAIL.n750 VSUBS 0.025512f
C1755 VTAIL.n751 VSUBS 0.023128f
C1756 VTAIL.n752 VSUBS 0.012428f
C1757 VTAIL.n753 VSUBS 0.029376f
C1758 VTAIL.n754 VSUBS 0.013159f
C1759 VTAIL.n755 VSUBS 0.023128f
C1760 VTAIL.n756 VSUBS 0.012428f
C1761 VTAIL.n757 VSUBS 0.029376f
C1762 VTAIL.n758 VSUBS 0.013159f
C1763 VTAIL.n759 VSUBS 0.023128f
C1764 VTAIL.n760 VSUBS 0.012428f
C1765 VTAIL.n761 VSUBS 0.029376f
C1766 VTAIL.n762 VSUBS 0.013159f
C1767 VTAIL.n763 VSUBS 0.023128f
C1768 VTAIL.n764 VSUBS 0.012428f
C1769 VTAIL.n765 VSUBS 0.029376f
C1770 VTAIL.n766 VSUBS 0.013159f
C1771 VTAIL.n767 VSUBS 0.023128f
C1772 VTAIL.n768 VSUBS 0.012428f
C1773 VTAIL.n769 VSUBS 0.029376f
C1774 VTAIL.n770 VSUBS 0.013159f
C1775 VTAIL.n771 VSUBS 0.023128f
C1776 VTAIL.n772 VSUBS 0.012428f
C1777 VTAIL.n773 VSUBS 0.029376f
C1778 VTAIL.n774 VSUBS 0.013159f
C1779 VTAIL.n775 VSUBS 0.023128f
C1780 VTAIL.n776 VSUBS 0.012428f
C1781 VTAIL.n777 VSUBS 0.029376f
C1782 VTAIL.n778 VSUBS 0.013159f
C1783 VTAIL.n779 VSUBS 0.023128f
C1784 VTAIL.n780 VSUBS 0.012428f
C1785 VTAIL.n781 VSUBS 0.029376f
C1786 VTAIL.n782 VSUBS 0.013159f
C1787 VTAIL.n783 VSUBS 0.189913f
C1788 VTAIL.t10 VSUBS 0.063114f
C1789 VTAIL.n784 VSUBS 0.022032f
C1790 VTAIL.n785 VSUBS 0.018687f
C1791 VTAIL.n786 VSUBS 0.012428f
C1792 VTAIL.n787 VSUBS 1.89048f
C1793 VTAIL.n788 VSUBS 0.023128f
C1794 VTAIL.n789 VSUBS 0.012428f
C1795 VTAIL.n790 VSUBS 0.013159f
C1796 VTAIL.n791 VSUBS 0.029376f
C1797 VTAIL.n792 VSUBS 0.029376f
C1798 VTAIL.n793 VSUBS 0.013159f
C1799 VTAIL.n794 VSUBS 0.012428f
C1800 VTAIL.n795 VSUBS 0.023128f
C1801 VTAIL.n796 VSUBS 0.023128f
C1802 VTAIL.n797 VSUBS 0.012428f
C1803 VTAIL.n798 VSUBS 0.013159f
C1804 VTAIL.n799 VSUBS 0.029376f
C1805 VTAIL.n800 VSUBS 0.029376f
C1806 VTAIL.n801 VSUBS 0.013159f
C1807 VTAIL.n802 VSUBS 0.012428f
C1808 VTAIL.n803 VSUBS 0.023128f
C1809 VTAIL.n804 VSUBS 0.023128f
C1810 VTAIL.n805 VSUBS 0.012428f
C1811 VTAIL.n806 VSUBS 0.013159f
C1812 VTAIL.n807 VSUBS 0.029376f
C1813 VTAIL.n808 VSUBS 0.029376f
C1814 VTAIL.n809 VSUBS 0.013159f
C1815 VTAIL.n810 VSUBS 0.012428f
C1816 VTAIL.n811 VSUBS 0.023128f
C1817 VTAIL.n812 VSUBS 0.023128f
C1818 VTAIL.n813 VSUBS 0.012428f
C1819 VTAIL.n814 VSUBS 0.013159f
C1820 VTAIL.n815 VSUBS 0.029376f
C1821 VTAIL.n816 VSUBS 0.029376f
C1822 VTAIL.n817 VSUBS 0.013159f
C1823 VTAIL.n818 VSUBS 0.012428f
C1824 VTAIL.n819 VSUBS 0.023128f
C1825 VTAIL.n820 VSUBS 0.023128f
C1826 VTAIL.n821 VSUBS 0.012428f
C1827 VTAIL.n822 VSUBS 0.013159f
C1828 VTAIL.n823 VSUBS 0.029376f
C1829 VTAIL.n824 VSUBS 0.029376f
C1830 VTAIL.n825 VSUBS 0.029376f
C1831 VTAIL.n826 VSUBS 0.013159f
C1832 VTAIL.n827 VSUBS 0.012428f
C1833 VTAIL.n828 VSUBS 0.023128f
C1834 VTAIL.n829 VSUBS 0.023128f
C1835 VTAIL.n830 VSUBS 0.012428f
C1836 VTAIL.n831 VSUBS 0.012794f
C1837 VTAIL.n832 VSUBS 0.012794f
C1838 VTAIL.n833 VSUBS 0.029376f
C1839 VTAIL.n834 VSUBS 0.029376f
C1840 VTAIL.n835 VSUBS 0.013159f
C1841 VTAIL.n836 VSUBS 0.012428f
C1842 VTAIL.n837 VSUBS 0.023128f
C1843 VTAIL.n838 VSUBS 0.023128f
C1844 VTAIL.n839 VSUBS 0.012428f
C1845 VTAIL.n840 VSUBS 0.013159f
C1846 VTAIL.n841 VSUBS 0.029376f
C1847 VTAIL.n842 VSUBS 0.029376f
C1848 VTAIL.n843 VSUBS 0.013159f
C1849 VTAIL.n844 VSUBS 0.012428f
C1850 VTAIL.n845 VSUBS 0.023128f
C1851 VTAIL.n846 VSUBS 0.023128f
C1852 VTAIL.n847 VSUBS 0.012428f
C1853 VTAIL.n848 VSUBS 0.013159f
C1854 VTAIL.n849 VSUBS 0.029376f
C1855 VTAIL.n850 VSUBS 0.071454f
C1856 VTAIL.n851 VSUBS 0.013159f
C1857 VTAIL.n852 VSUBS 0.012428f
C1858 VTAIL.n853 VSUBS 0.052828f
C1859 VTAIL.n854 VSUBS 0.035929f
C1860 VTAIL.n855 VSUBS 1.81202f
C1861 VN.n0 VSUBS 0.032656f
C1862 VN.t1 VSUBS 2.96295f
C1863 VN.n1 VSUBS 0.028557f
C1864 VN.n2 VSUBS 0.032656f
C1865 VN.t2 VSUBS 2.96295f
C1866 VN.n3 VSUBS 0.026426f
C1867 VN.n4 VSUBS 0.21027f
C1868 VN.t0 VSUBS 2.96295f
C1869 VN.t6 VSUBS 3.08535f
C1870 VN.n5 VSUBS 1.12422f
C1871 VN.n6 VSUBS 1.09332f
C1872 VN.n7 VSUBS 0.033081f
C1873 VN.n8 VSUBS 0.065251f
C1874 VN.n9 VSUBS 0.032656f
C1875 VN.n10 VSUBS 0.032656f
C1876 VN.n11 VSUBS 0.032656f
C1877 VN.n12 VSUBS 0.065251f
C1878 VN.n13 VSUBS 0.033081f
C1879 VN.n14 VSUBS 1.03554f
C1880 VN.n15 VSUBS 0.06421f
C1881 VN.n16 VSUBS 0.032656f
C1882 VN.n17 VSUBS 0.032656f
C1883 VN.n18 VSUBS 0.032656f
C1884 VN.n19 VSUBS 0.062046f
C1885 VN.n20 VSUBS 0.037309f
C1886 VN.n21 VSUBS 1.10881f
C1887 VN.n22 VSUBS 0.034043f
C1888 VN.n23 VSUBS 0.032656f
C1889 VN.t3 VSUBS 2.96295f
C1890 VN.n24 VSUBS 0.028557f
C1891 VN.n25 VSUBS 0.032656f
C1892 VN.t7 VSUBS 2.96295f
C1893 VN.n26 VSUBS 0.026426f
C1894 VN.n27 VSUBS 0.21027f
C1895 VN.t5 VSUBS 2.96295f
C1896 VN.t4 VSUBS 3.08535f
C1897 VN.n28 VSUBS 1.12422f
C1898 VN.n29 VSUBS 1.09332f
C1899 VN.n30 VSUBS 0.033081f
C1900 VN.n31 VSUBS 0.065251f
C1901 VN.n32 VSUBS 0.032656f
C1902 VN.n33 VSUBS 0.032656f
C1903 VN.n34 VSUBS 0.032656f
C1904 VN.n35 VSUBS 0.065251f
C1905 VN.n36 VSUBS 0.033081f
C1906 VN.n37 VSUBS 1.03554f
C1907 VN.n38 VSUBS 0.06421f
C1908 VN.n39 VSUBS 0.032656f
C1909 VN.n40 VSUBS 0.032656f
C1910 VN.n41 VSUBS 0.032656f
C1911 VN.n42 VSUBS 0.062046f
C1912 VN.n43 VSUBS 0.037309f
C1913 VN.n44 VSUBS 1.10881f
C1914 VN.n45 VSUBS 1.91417f
.ends

