* NGSPICE file created from diff_pair_sample_0457.ext - technology: sky130A

.subckt diff_pair_sample_0457 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=3.2
X1 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=3.2
X2 VTAIL.t7 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=3.2
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=3.2
X4 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=3.2
X5 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=3.2
X6 VDD1.t1 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=3.2
X7 VTAIL.t1 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=3.2
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=3.2
X9 VDD1.t2 VP.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=3.2
X10 VTAIL.t4 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=3.2
X11 VDD2.t0 VN.t3 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=3.2
R0 B.n1018 B.n1017 585
R1 B.n1019 B.n1018 585
R2 B.n421 B.n143 585
R3 B.n420 B.n419 585
R4 B.n418 B.n417 585
R5 B.n416 B.n415 585
R6 B.n414 B.n413 585
R7 B.n412 B.n411 585
R8 B.n410 B.n409 585
R9 B.n408 B.n407 585
R10 B.n406 B.n405 585
R11 B.n404 B.n403 585
R12 B.n402 B.n401 585
R13 B.n400 B.n399 585
R14 B.n398 B.n397 585
R15 B.n396 B.n395 585
R16 B.n394 B.n393 585
R17 B.n392 B.n391 585
R18 B.n390 B.n389 585
R19 B.n388 B.n387 585
R20 B.n386 B.n385 585
R21 B.n384 B.n383 585
R22 B.n382 B.n381 585
R23 B.n380 B.n379 585
R24 B.n378 B.n377 585
R25 B.n376 B.n375 585
R26 B.n374 B.n373 585
R27 B.n372 B.n371 585
R28 B.n370 B.n369 585
R29 B.n368 B.n367 585
R30 B.n366 B.n365 585
R31 B.n364 B.n363 585
R32 B.n362 B.n361 585
R33 B.n360 B.n359 585
R34 B.n358 B.n357 585
R35 B.n356 B.n355 585
R36 B.n354 B.n353 585
R37 B.n352 B.n351 585
R38 B.n350 B.n349 585
R39 B.n348 B.n347 585
R40 B.n346 B.n345 585
R41 B.n344 B.n343 585
R42 B.n342 B.n341 585
R43 B.n340 B.n339 585
R44 B.n338 B.n337 585
R45 B.n336 B.n335 585
R46 B.n334 B.n333 585
R47 B.n332 B.n331 585
R48 B.n330 B.n329 585
R49 B.n328 B.n327 585
R50 B.n326 B.n325 585
R51 B.n324 B.n323 585
R52 B.n322 B.n321 585
R53 B.n320 B.n319 585
R54 B.n318 B.n317 585
R55 B.n316 B.n315 585
R56 B.n314 B.n313 585
R57 B.n312 B.n311 585
R58 B.n310 B.n309 585
R59 B.n308 B.n307 585
R60 B.n306 B.n305 585
R61 B.n304 B.n303 585
R62 B.n302 B.n301 585
R63 B.n300 B.n299 585
R64 B.n298 B.n297 585
R65 B.n296 B.n295 585
R66 B.n294 B.n293 585
R67 B.n292 B.n291 585
R68 B.n290 B.n289 585
R69 B.n288 B.n287 585
R70 B.n286 B.n285 585
R71 B.n284 B.n283 585
R72 B.n282 B.n281 585
R73 B.n280 B.n279 585
R74 B.n278 B.n277 585
R75 B.n275 B.n274 585
R76 B.n273 B.n272 585
R77 B.n271 B.n270 585
R78 B.n269 B.n268 585
R79 B.n267 B.n266 585
R80 B.n265 B.n264 585
R81 B.n263 B.n262 585
R82 B.n261 B.n260 585
R83 B.n259 B.n258 585
R84 B.n257 B.n256 585
R85 B.n255 B.n254 585
R86 B.n253 B.n252 585
R87 B.n251 B.n250 585
R88 B.n249 B.n248 585
R89 B.n247 B.n246 585
R90 B.n245 B.n244 585
R91 B.n243 B.n242 585
R92 B.n241 B.n240 585
R93 B.n239 B.n238 585
R94 B.n237 B.n236 585
R95 B.n235 B.n234 585
R96 B.n233 B.n232 585
R97 B.n231 B.n230 585
R98 B.n229 B.n228 585
R99 B.n227 B.n226 585
R100 B.n225 B.n224 585
R101 B.n223 B.n222 585
R102 B.n221 B.n220 585
R103 B.n219 B.n218 585
R104 B.n217 B.n216 585
R105 B.n215 B.n214 585
R106 B.n213 B.n212 585
R107 B.n211 B.n210 585
R108 B.n209 B.n208 585
R109 B.n207 B.n206 585
R110 B.n205 B.n204 585
R111 B.n203 B.n202 585
R112 B.n201 B.n200 585
R113 B.n199 B.n198 585
R114 B.n197 B.n196 585
R115 B.n195 B.n194 585
R116 B.n193 B.n192 585
R117 B.n191 B.n190 585
R118 B.n189 B.n188 585
R119 B.n187 B.n186 585
R120 B.n185 B.n184 585
R121 B.n183 B.n182 585
R122 B.n181 B.n180 585
R123 B.n179 B.n178 585
R124 B.n177 B.n176 585
R125 B.n175 B.n174 585
R126 B.n173 B.n172 585
R127 B.n171 B.n170 585
R128 B.n169 B.n168 585
R129 B.n167 B.n166 585
R130 B.n165 B.n164 585
R131 B.n163 B.n162 585
R132 B.n161 B.n160 585
R133 B.n159 B.n158 585
R134 B.n157 B.n156 585
R135 B.n155 B.n154 585
R136 B.n153 B.n152 585
R137 B.n151 B.n150 585
R138 B.n74 B.n73 585
R139 B.n1022 B.n1021 585
R140 B.n1016 B.n144 585
R141 B.n144 B.n71 585
R142 B.n1015 B.n70 585
R143 B.n1026 B.n70 585
R144 B.n1014 B.n69 585
R145 B.n1027 B.n69 585
R146 B.n1013 B.n68 585
R147 B.n1028 B.n68 585
R148 B.n1012 B.n1011 585
R149 B.n1011 B.n64 585
R150 B.n1010 B.n63 585
R151 B.n1034 B.n63 585
R152 B.n1009 B.n62 585
R153 B.n1035 B.n62 585
R154 B.n1008 B.n61 585
R155 B.n1036 B.n61 585
R156 B.n1007 B.n1006 585
R157 B.n1006 B.n60 585
R158 B.n1005 B.n56 585
R159 B.n1042 B.n56 585
R160 B.n1004 B.n55 585
R161 B.n1043 B.n55 585
R162 B.n1003 B.n54 585
R163 B.n1044 B.n54 585
R164 B.n1002 B.n1001 585
R165 B.n1001 B.n50 585
R166 B.n1000 B.n49 585
R167 B.n1050 B.n49 585
R168 B.n999 B.n48 585
R169 B.n1051 B.n48 585
R170 B.n998 B.n47 585
R171 B.n1052 B.n47 585
R172 B.n997 B.n996 585
R173 B.n996 B.n43 585
R174 B.n995 B.n42 585
R175 B.n1058 B.n42 585
R176 B.n994 B.n41 585
R177 B.n1059 B.n41 585
R178 B.n993 B.n40 585
R179 B.n1060 B.n40 585
R180 B.n992 B.n991 585
R181 B.n991 B.n36 585
R182 B.n990 B.n35 585
R183 B.n1066 B.n35 585
R184 B.n989 B.n34 585
R185 B.n1067 B.n34 585
R186 B.n988 B.n33 585
R187 B.n1068 B.n33 585
R188 B.n987 B.n986 585
R189 B.n986 B.n29 585
R190 B.n985 B.n28 585
R191 B.n1074 B.n28 585
R192 B.n984 B.n27 585
R193 B.n1075 B.n27 585
R194 B.n983 B.n26 585
R195 B.n1076 B.n26 585
R196 B.n982 B.n981 585
R197 B.n981 B.n22 585
R198 B.n980 B.n21 585
R199 B.n1082 B.n21 585
R200 B.n979 B.n20 585
R201 B.n1083 B.n20 585
R202 B.n978 B.n19 585
R203 B.n1084 B.n19 585
R204 B.n977 B.n976 585
R205 B.n976 B.n18 585
R206 B.n975 B.n14 585
R207 B.n1090 B.n14 585
R208 B.n974 B.n13 585
R209 B.n1091 B.n13 585
R210 B.n973 B.n12 585
R211 B.n1092 B.n12 585
R212 B.n972 B.n971 585
R213 B.n971 B.n8 585
R214 B.n970 B.n7 585
R215 B.n1098 B.n7 585
R216 B.n969 B.n6 585
R217 B.n1099 B.n6 585
R218 B.n968 B.n5 585
R219 B.n1100 B.n5 585
R220 B.n967 B.n966 585
R221 B.n966 B.n4 585
R222 B.n965 B.n422 585
R223 B.n965 B.n964 585
R224 B.n955 B.n423 585
R225 B.n424 B.n423 585
R226 B.n957 B.n956 585
R227 B.n958 B.n957 585
R228 B.n954 B.n429 585
R229 B.n429 B.n428 585
R230 B.n953 B.n952 585
R231 B.n952 B.n951 585
R232 B.n431 B.n430 585
R233 B.n944 B.n431 585
R234 B.n943 B.n942 585
R235 B.n945 B.n943 585
R236 B.n941 B.n436 585
R237 B.n436 B.n435 585
R238 B.n940 B.n939 585
R239 B.n939 B.n938 585
R240 B.n438 B.n437 585
R241 B.n439 B.n438 585
R242 B.n931 B.n930 585
R243 B.n932 B.n931 585
R244 B.n929 B.n444 585
R245 B.n444 B.n443 585
R246 B.n928 B.n927 585
R247 B.n927 B.n926 585
R248 B.n446 B.n445 585
R249 B.n447 B.n446 585
R250 B.n919 B.n918 585
R251 B.n920 B.n919 585
R252 B.n917 B.n452 585
R253 B.n452 B.n451 585
R254 B.n916 B.n915 585
R255 B.n915 B.n914 585
R256 B.n454 B.n453 585
R257 B.n455 B.n454 585
R258 B.n907 B.n906 585
R259 B.n908 B.n907 585
R260 B.n905 B.n460 585
R261 B.n460 B.n459 585
R262 B.n904 B.n903 585
R263 B.n903 B.n902 585
R264 B.n462 B.n461 585
R265 B.n463 B.n462 585
R266 B.n895 B.n894 585
R267 B.n896 B.n895 585
R268 B.n893 B.n468 585
R269 B.n468 B.n467 585
R270 B.n892 B.n891 585
R271 B.n891 B.n890 585
R272 B.n470 B.n469 585
R273 B.n471 B.n470 585
R274 B.n883 B.n882 585
R275 B.n884 B.n883 585
R276 B.n881 B.n476 585
R277 B.n476 B.n475 585
R278 B.n880 B.n879 585
R279 B.n879 B.n878 585
R280 B.n478 B.n477 585
R281 B.n871 B.n478 585
R282 B.n870 B.n869 585
R283 B.n872 B.n870 585
R284 B.n868 B.n483 585
R285 B.n483 B.n482 585
R286 B.n867 B.n866 585
R287 B.n866 B.n865 585
R288 B.n485 B.n484 585
R289 B.n486 B.n485 585
R290 B.n858 B.n857 585
R291 B.n859 B.n858 585
R292 B.n856 B.n491 585
R293 B.n491 B.n490 585
R294 B.n855 B.n854 585
R295 B.n854 B.n853 585
R296 B.n493 B.n492 585
R297 B.n494 B.n493 585
R298 B.n849 B.n848 585
R299 B.n497 B.n496 585
R300 B.n845 B.n844 585
R301 B.n846 B.n845 585
R302 B.n843 B.n566 585
R303 B.n842 B.n841 585
R304 B.n840 B.n839 585
R305 B.n838 B.n837 585
R306 B.n836 B.n835 585
R307 B.n834 B.n833 585
R308 B.n832 B.n831 585
R309 B.n830 B.n829 585
R310 B.n828 B.n827 585
R311 B.n826 B.n825 585
R312 B.n824 B.n823 585
R313 B.n822 B.n821 585
R314 B.n820 B.n819 585
R315 B.n818 B.n817 585
R316 B.n816 B.n815 585
R317 B.n814 B.n813 585
R318 B.n812 B.n811 585
R319 B.n810 B.n809 585
R320 B.n808 B.n807 585
R321 B.n806 B.n805 585
R322 B.n804 B.n803 585
R323 B.n802 B.n801 585
R324 B.n800 B.n799 585
R325 B.n798 B.n797 585
R326 B.n796 B.n795 585
R327 B.n794 B.n793 585
R328 B.n792 B.n791 585
R329 B.n790 B.n789 585
R330 B.n788 B.n787 585
R331 B.n786 B.n785 585
R332 B.n784 B.n783 585
R333 B.n782 B.n781 585
R334 B.n780 B.n779 585
R335 B.n778 B.n777 585
R336 B.n776 B.n775 585
R337 B.n774 B.n773 585
R338 B.n772 B.n771 585
R339 B.n770 B.n769 585
R340 B.n768 B.n767 585
R341 B.n766 B.n765 585
R342 B.n764 B.n763 585
R343 B.n762 B.n761 585
R344 B.n760 B.n759 585
R345 B.n758 B.n757 585
R346 B.n756 B.n755 585
R347 B.n754 B.n753 585
R348 B.n752 B.n751 585
R349 B.n750 B.n749 585
R350 B.n748 B.n747 585
R351 B.n746 B.n745 585
R352 B.n744 B.n743 585
R353 B.n742 B.n741 585
R354 B.n740 B.n739 585
R355 B.n738 B.n737 585
R356 B.n736 B.n735 585
R357 B.n734 B.n733 585
R358 B.n732 B.n731 585
R359 B.n730 B.n729 585
R360 B.n728 B.n727 585
R361 B.n726 B.n725 585
R362 B.n724 B.n723 585
R363 B.n722 B.n721 585
R364 B.n720 B.n719 585
R365 B.n718 B.n717 585
R366 B.n716 B.n715 585
R367 B.n714 B.n713 585
R368 B.n712 B.n711 585
R369 B.n710 B.n709 585
R370 B.n708 B.n707 585
R371 B.n706 B.n705 585
R372 B.n704 B.n703 585
R373 B.n701 B.n700 585
R374 B.n699 B.n698 585
R375 B.n697 B.n696 585
R376 B.n695 B.n694 585
R377 B.n693 B.n692 585
R378 B.n691 B.n690 585
R379 B.n689 B.n688 585
R380 B.n687 B.n686 585
R381 B.n685 B.n684 585
R382 B.n683 B.n682 585
R383 B.n681 B.n680 585
R384 B.n679 B.n678 585
R385 B.n677 B.n676 585
R386 B.n675 B.n674 585
R387 B.n673 B.n672 585
R388 B.n671 B.n670 585
R389 B.n669 B.n668 585
R390 B.n667 B.n666 585
R391 B.n665 B.n664 585
R392 B.n663 B.n662 585
R393 B.n661 B.n660 585
R394 B.n659 B.n658 585
R395 B.n657 B.n656 585
R396 B.n655 B.n654 585
R397 B.n653 B.n652 585
R398 B.n651 B.n650 585
R399 B.n649 B.n648 585
R400 B.n647 B.n646 585
R401 B.n645 B.n644 585
R402 B.n643 B.n642 585
R403 B.n641 B.n640 585
R404 B.n639 B.n638 585
R405 B.n637 B.n636 585
R406 B.n635 B.n634 585
R407 B.n633 B.n632 585
R408 B.n631 B.n630 585
R409 B.n629 B.n628 585
R410 B.n627 B.n626 585
R411 B.n625 B.n624 585
R412 B.n623 B.n622 585
R413 B.n621 B.n620 585
R414 B.n619 B.n618 585
R415 B.n617 B.n616 585
R416 B.n615 B.n614 585
R417 B.n613 B.n612 585
R418 B.n611 B.n610 585
R419 B.n609 B.n608 585
R420 B.n607 B.n606 585
R421 B.n605 B.n604 585
R422 B.n603 B.n602 585
R423 B.n601 B.n600 585
R424 B.n599 B.n598 585
R425 B.n597 B.n596 585
R426 B.n595 B.n594 585
R427 B.n593 B.n592 585
R428 B.n591 B.n590 585
R429 B.n589 B.n588 585
R430 B.n587 B.n586 585
R431 B.n585 B.n584 585
R432 B.n583 B.n582 585
R433 B.n581 B.n580 585
R434 B.n579 B.n578 585
R435 B.n577 B.n576 585
R436 B.n575 B.n574 585
R437 B.n573 B.n572 585
R438 B.n850 B.n495 585
R439 B.n495 B.n494 585
R440 B.n852 B.n851 585
R441 B.n853 B.n852 585
R442 B.n489 B.n488 585
R443 B.n490 B.n489 585
R444 B.n861 B.n860 585
R445 B.n860 B.n859 585
R446 B.n862 B.n487 585
R447 B.n487 B.n486 585
R448 B.n864 B.n863 585
R449 B.n865 B.n864 585
R450 B.n481 B.n480 585
R451 B.n482 B.n481 585
R452 B.n874 B.n873 585
R453 B.n873 B.n872 585
R454 B.n875 B.n479 585
R455 B.n871 B.n479 585
R456 B.n877 B.n876 585
R457 B.n878 B.n877 585
R458 B.n474 B.n473 585
R459 B.n475 B.n474 585
R460 B.n886 B.n885 585
R461 B.n885 B.n884 585
R462 B.n887 B.n472 585
R463 B.n472 B.n471 585
R464 B.n889 B.n888 585
R465 B.n890 B.n889 585
R466 B.n466 B.n465 585
R467 B.n467 B.n466 585
R468 B.n898 B.n897 585
R469 B.n897 B.n896 585
R470 B.n899 B.n464 585
R471 B.n464 B.n463 585
R472 B.n901 B.n900 585
R473 B.n902 B.n901 585
R474 B.n458 B.n457 585
R475 B.n459 B.n458 585
R476 B.n910 B.n909 585
R477 B.n909 B.n908 585
R478 B.n911 B.n456 585
R479 B.n456 B.n455 585
R480 B.n913 B.n912 585
R481 B.n914 B.n913 585
R482 B.n450 B.n449 585
R483 B.n451 B.n450 585
R484 B.n922 B.n921 585
R485 B.n921 B.n920 585
R486 B.n923 B.n448 585
R487 B.n448 B.n447 585
R488 B.n925 B.n924 585
R489 B.n926 B.n925 585
R490 B.n442 B.n441 585
R491 B.n443 B.n442 585
R492 B.n934 B.n933 585
R493 B.n933 B.n932 585
R494 B.n935 B.n440 585
R495 B.n440 B.n439 585
R496 B.n937 B.n936 585
R497 B.n938 B.n937 585
R498 B.n434 B.n433 585
R499 B.n435 B.n434 585
R500 B.n947 B.n946 585
R501 B.n946 B.n945 585
R502 B.n948 B.n432 585
R503 B.n944 B.n432 585
R504 B.n950 B.n949 585
R505 B.n951 B.n950 585
R506 B.n427 B.n426 585
R507 B.n428 B.n427 585
R508 B.n960 B.n959 585
R509 B.n959 B.n958 585
R510 B.n961 B.n425 585
R511 B.n425 B.n424 585
R512 B.n963 B.n962 585
R513 B.n964 B.n963 585
R514 B.n2 B.n0 585
R515 B.n4 B.n2 585
R516 B.n3 B.n1 585
R517 B.n1099 B.n3 585
R518 B.n1097 B.n1096 585
R519 B.n1098 B.n1097 585
R520 B.n1095 B.n9 585
R521 B.n9 B.n8 585
R522 B.n1094 B.n1093 585
R523 B.n1093 B.n1092 585
R524 B.n11 B.n10 585
R525 B.n1091 B.n11 585
R526 B.n1089 B.n1088 585
R527 B.n1090 B.n1089 585
R528 B.n1087 B.n15 585
R529 B.n18 B.n15 585
R530 B.n1086 B.n1085 585
R531 B.n1085 B.n1084 585
R532 B.n17 B.n16 585
R533 B.n1083 B.n17 585
R534 B.n1081 B.n1080 585
R535 B.n1082 B.n1081 585
R536 B.n1079 B.n23 585
R537 B.n23 B.n22 585
R538 B.n1078 B.n1077 585
R539 B.n1077 B.n1076 585
R540 B.n25 B.n24 585
R541 B.n1075 B.n25 585
R542 B.n1073 B.n1072 585
R543 B.n1074 B.n1073 585
R544 B.n1071 B.n30 585
R545 B.n30 B.n29 585
R546 B.n1070 B.n1069 585
R547 B.n1069 B.n1068 585
R548 B.n32 B.n31 585
R549 B.n1067 B.n32 585
R550 B.n1065 B.n1064 585
R551 B.n1066 B.n1065 585
R552 B.n1063 B.n37 585
R553 B.n37 B.n36 585
R554 B.n1062 B.n1061 585
R555 B.n1061 B.n1060 585
R556 B.n39 B.n38 585
R557 B.n1059 B.n39 585
R558 B.n1057 B.n1056 585
R559 B.n1058 B.n1057 585
R560 B.n1055 B.n44 585
R561 B.n44 B.n43 585
R562 B.n1054 B.n1053 585
R563 B.n1053 B.n1052 585
R564 B.n46 B.n45 585
R565 B.n1051 B.n46 585
R566 B.n1049 B.n1048 585
R567 B.n1050 B.n1049 585
R568 B.n1047 B.n51 585
R569 B.n51 B.n50 585
R570 B.n1046 B.n1045 585
R571 B.n1045 B.n1044 585
R572 B.n53 B.n52 585
R573 B.n1043 B.n53 585
R574 B.n1041 B.n1040 585
R575 B.n1042 B.n1041 585
R576 B.n1039 B.n57 585
R577 B.n60 B.n57 585
R578 B.n1038 B.n1037 585
R579 B.n1037 B.n1036 585
R580 B.n59 B.n58 585
R581 B.n1035 B.n59 585
R582 B.n1033 B.n1032 585
R583 B.n1034 B.n1033 585
R584 B.n1031 B.n65 585
R585 B.n65 B.n64 585
R586 B.n1030 B.n1029 585
R587 B.n1029 B.n1028 585
R588 B.n67 B.n66 585
R589 B.n1027 B.n67 585
R590 B.n1025 B.n1024 585
R591 B.n1026 B.n1025 585
R592 B.n1023 B.n72 585
R593 B.n72 B.n71 585
R594 B.n1102 B.n1101 585
R595 B.n1101 B.n1100 585
R596 B.n848 B.n495 564.573
R597 B.n1021 B.n72 564.573
R598 B.n572 B.n493 564.573
R599 B.n1018 B.n144 564.573
R600 B.n570 B.t8 358.675
R601 B.n567 B.t12 358.675
R602 B.n148 B.t15 358.675
R603 B.n145 B.t4 358.675
R604 B.n1019 B.n142 256.663
R605 B.n1019 B.n141 256.663
R606 B.n1019 B.n140 256.663
R607 B.n1019 B.n139 256.663
R608 B.n1019 B.n138 256.663
R609 B.n1019 B.n137 256.663
R610 B.n1019 B.n136 256.663
R611 B.n1019 B.n135 256.663
R612 B.n1019 B.n134 256.663
R613 B.n1019 B.n133 256.663
R614 B.n1019 B.n132 256.663
R615 B.n1019 B.n131 256.663
R616 B.n1019 B.n130 256.663
R617 B.n1019 B.n129 256.663
R618 B.n1019 B.n128 256.663
R619 B.n1019 B.n127 256.663
R620 B.n1019 B.n126 256.663
R621 B.n1019 B.n125 256.663
R622 B.n1019 B.n124 256.663
R623 B.n1019 B.n123 256.663
R624 B.n1019 B.n122 256.663
R625 B.n1019 B.n121 256.663
R626 B.n1019 B.n120 256.663
R627 B.n1019 B.n119 256.663
R628 B.n1019 B.n118 256.663
R629 B.n1019 B.n117 256.663
R630 B.n1019 B.n116 256.663
R631 B.n1019 B.n115 256.663
R632 B.n1019 B.n114 256.663
R633 B.n1019 B.n113 256.663
R634 B.n1019 B.n112 256.663
R635 B.n1019 B.n111 256.663
R636 B.n1019 B.n110 256.663
R637 B.n1019 B.n109 256.663
R638 B.n1019 B.n108 256.663
R639 B.n1019 B.n107 256.663
R640 B.n1019 B.n106 256.663
R641 B.n1019 B.n105 256.663
R642 B.n1019 B.n104 256.663
R643 B.n1019 B.n103 256.663
R644 B.n1019 B.n102 256.663
R645 B.n1019 B.n101 256.663
R646 B.n1019 B.n100 256.663
R647 B.n1019 B.n99 256.663
R648 B.n1019 B.n98 256.663
R649 B.n1019 B.n97 256.663
R650 B.n1019 B.n96 256.663
R651 B.n1019 B.n95 256.663
R652 B.n1019 B.n94 256.663
R653 B.n1019 B.n93 256.663
R654 B.n1019 B.n92 256.663
R655 B.n1019 B.n91 256.663
R656 B.n1019 B.n90 256.663
R657 B.n1019 B.n89 256.663
R658 B.n1019 B.n88 256.663
R659 B.n1019 B.n87 256.663
R660 B.n1019 B.n86 256.663
R661 B.n1019 B.n85 256.663
R662 B.n1019 B.n84 256.663
R663 B.n1019 B.n83 256.663
R664 B.n1019 B.n82 256.663
R665 B.n1019 B.n81 256.663
R666 B.n1019 B.n80 256.663
R667 B.n1019 B.n79 256.663
R668 B.n1019 B.n78 256.663
R669 B.n1019 B.n77 256.663
R670 B.n1019 B.n76 256.663
R671 B.n1019 B.n75 256.663
R672 B.n1020 B.n1019 256.663
R673 B.n847 B.n846 256.663
R674 B.n846 B.n498 256.663
R675 B.n846 B.n499 256.663
R676 B.n846 B.n500 256.663
R677 B.n846 B.n501 256.663
R678 B.n846 B.n502 256.663
R679 B.n846 B.n503 256.663
R680 B.n846 B.n504 256.663
R681 B.n846 B.n505 256.663
R682 B.n846 B.n506 256.663
R683 B.n846 B.n507 256.663
R684 B.n846 B.n508 256.663
R685 B.n846 B.n509 256.663
R686 B.n846 B.n510 256.663
R687 B.n846 B.n511 256.663
R688 B.n846 B.n512 256.663
R689 B.n846 B.n513 256.663
R690 B.n846 B.n514 256.663
R691 B.n846 B.n515 256.663
R692 B.n846 B.n516 256.663
R693 B.n846 B.n517 256.663
R694 B.n846 B.n518 256.663
R695 B.n846 B.n519 256.663
R696 B.n846 B.n520 256.663
R697 B.n846 B.n521 256.663
R698 B.n846 B.n522 256.663
R699 B.n846 B.n523 256.663
R700 B.n846 B.n524 256.663
R701 B.n846 B.n525 256.663
R702 B.n846 B.n526 256.663
R703 B.n846 B.n527 256.663
R704 B.n846 B.n528 256.663
R705 B.n846 B.n529 256.663
R706 B.n846 B.n530 256.663
R707 B.n846 B.n531 256.663
R708 B.n846 B.n532 256.663
R709 B.n846 B.n533 256.663
R710 B.n846 B.n534 256.663
R711 B.n846 B.n535 256.663
R712 B.n846 B.n536 256.663
R713 B.n846 B.n537 256.663
R714 B.n846 B.n538 256.663
R715 B.n846 B.n539 256.663
R716 B.n846 B.n540 256.663
R717 B.n846 B.n541 256.663
R718 B.n846 B.n542 256.663
R719 B.n846 B.n543 256.663
R720 B.n846 B.n544 256.663
R721 B.n846 B.n545 256.663
R722 B.n846 B.n546 256.663
R723 B.n846 B.n547 256.663
R724 B.n846 B.n548 256.663
R725 B.n846 B.n549 256.663
R726 B.n846 B.n550 256.663
R727 B.n846 B.n551 256.663
R728 B.n846 B.n552 256.663
R729 B.n846 B.n553 256.663
R730 B.n846 B.n554 256.663
R731 B.n846 B.n555 256.663
R732 B.n846 B.n556 256.663
R733 B.n846 B.n557 256.663
R734 B.n846 B.n558 256.663
R735 B.n846 B.n559 256.663
R736 B.n846 B.n560 256.663
R737 B.n846 B.n561 256.663
R738 B.n846 B.n562 256.663
R739 B.n846 B.n563 256.663
R740 B.n846 B.n564 256.663
R741 B.n846 B.n565 256.663
R742 B.n852 B.n495 163.367
R743 B.n852 B.n489 163.367
R744 B.n860 B.n489 163.367
R745 B.n860 B.n487 163.367
R746 B.n864 B.n487 163.367
R747 B.n864 B.n481 163.367
R748 B.n873 B.n481 163.367
R749 B.n873 B.n479 163.367
R750 B.n877 B.n479 163.367
R751 B.n877 B.n474 163.367
R752 B.n885 B.n474 163.367
R753 B.n885 B.n472 163.367
R754 B.n889 B.n472 163.367
R755 B.n889 B.n466 163.367
R756 B.n897 B.n466 163.367
R757 B.n897 B.n464 163.367
R758 B.n901 B.n464 163.367
R759 B.n901 B.n458 163.367
R760 B.n909 B.n458 163.367
R761 B.n909 B.n456 163.367
R762 B.n913 B.n456 163.367
R763 B.n913 B.n450 163.367
R764 B.n921 B.n450 163.367
R765 B.n921 B.n448 163.367
R766 B.n925 B.n448 163.367
R767 B.n925 B.n442 163.367
R768 B.n933 B.n442 163.367
R769 B.n933 B.n440 163.367
R770 B.n937 B.n440 163.367
R771 B.n937 B.n434 163.367
R772 B.n946 B.n434 163.367
R773 B.n946 B.n432 163.367
R774 B.n950 B.n432 163.367
R775 B.n950 B.n427 163.367
R776 B.n959 B.n427 163.367
R777 B.n959 B.n425 163.367
R778 B.n963 B.n425 163.367
R779 B.n963 B.n2 163.367
R780 B.n1101 B.n2 163.367
R781 B.n1101 B.n3 163.367
R782 B.n1097 B.n3 163.367
R783 B.n1097 B.n9 163.367
R784 B.n1093 B.n9 163.367
R785 B.n1093 B.n11 163.367
R786 B.n1089 B.n11 163.367
R787 B.n1089 B.n15 163.367
R788 B.n1085 B.n15 163.367
R789 B.n1085 B.n17 163.367
R790 B.n1081 B.n17 163.367
R791 B.n1081 B.n23 163.367
R792 B.n1077 B.n23 163.367
R793 B.n1077 B.n25 163.367
R794 B.n1073 B.n25 163.367
R795 B.n1073 B.n30 163.367
R796 B.n1069 B.n30 163.367
R797 B.n1069 B.n32 163.367
R798 B.n1065 B.n32 163.367
R799 B.n1065 B.n37 163.367
R800 B.n1061 B.n37 163.367
R801 B.n1061 B.n39 163.367
R802 B.n1057 B.n39 163.367
R803 B.n1057 B.n44 163.367
R804 B.n1053 B.n44 163.367
R805 B.n1053 B.n46 163.367
R806 B.n1049 B.n46 163.367
R807 B.n1049 B.n51 163.367
R808 B.n1045 B.n51 163.367
R809 B.n1045 B.n53 163.367
R810 B.n1041 B.n53 163.367
R811 B.n1041 B.n57 163.367
R812 B.n1037 B.n57 163.367
R813 B.n1037 B.n59 163.367
R814 B.n1033 B.n59 163.367
R815 B.n1033 B.n65 163.367
R816 B.n1029 B.n65 163.367
R817 B.n1029 B.n67 163.367
R818 B.n1025 B.n67 163.367
R819 B.n1025 B.n72 163.367
R820 B.n845 B.n497 163.367
R821 B.n845 B.n566 163.367
R822 B.n841 B.n840 163.367
R823 B.n837 B.n836 163.367
R824 B.n833 B.n832 163.367
R825 B.n829 B.n828 163.367
R826 B.n825 B.n824 163.367
R827 B.n821 B.n820 163.367
R828 B.n817 B.n816 163.367
R829 B.n813 B.n812 163.367
R830 B.n809 B.n808 163.367
R831 B.n805 B.n804 163.367
R832 B.n801 B.n800 163.367
R833 B.n797 B.n796 163.367
R834 B.n793 B.n792 163.367
R835 B.n789 B.n788 163.367
R836 B.n785 B.n784 163.367
R837 B.n781 B.n780 163.367
R838 B.n777 B.n776 163.367
R839 B.n773 B.n772 163.367
R840 B.n769 B.n768 163.367
R841 B.n765 B.n764 163.367
R842 B.n761 B.n760 163.367
R843 B.n757 B.n756 163.367
R844 B.n753 B.n752 163.367
R845 B.n749 B.n748 163.367
R846 B.n745 B.n744 163.367
R847 B.n741 B.n740 163.367
R848 B.n737 B.n736 163.367
R849 B.n733 B.n732 163.367
R850 B.n729 B.n728 163.367
R851 B.n725 B.n724 163.367
R852 B.n721 B.n720 163.367
R853 B.n717 B.n716 163.367
R854 B.n713 B.n712 163.367
R855 B.n709 B.n708 163.367
R856 B.n705 B.n704 163.367
R857 B.n700 B.n699 163.367
R858 B.n696 B.n695 163.367
R859 B.n692 B.n691 163.367
R860 B.n688 B.n687 163.367
R861 B.n684 B.n683 163.367
R862 B.n680 B.n679 163.367
R863 B.n676 B.n675 163.367
R864 B.n672 B.n671 163.367
R865 B.n668 B.n667 163.367
R866 B.n664 B.n663 163.367
R867 B.n660 B.n659 163.367
R868 B.n656 B.n655 163.367
R869 B.n652 B.n651 163.367
R870 B.n648 B.n647 163.367
R871 B.n644 B.n643 163.367
R872 B.n640 B.n639 163.367
R873 B.n636 B.n635 163.367
R874 B.n632 B.n631 163.367
R875 B.n628 B.n627 163.367
R876 B.n624 B.n623 163.367
R877 B.n620 B.n619 163.367
R878 B.n616 B.n615 163.367
R879 B.n612 B.n611 163.367
R880 B.n608 B.n607 163.367
R881 B.n604 B.n603 163.367
R882 B.n600 B.n599 163.367
R883 B.n596 B.n595 163.367
R884 B.n592 B.n591 163.367
R885 B.n588 B.n587 163.367
R886 B.n584 B.n583 163.367
R887 B.n580 B.n579 163.367
R888 B.n576 B.n575 163.367
R889 B.n854 B.n493 163.367
R890 B.n854 B.n491 163.367
R891 B.n858 B.n491 163.367
R892 B.n858 B.n485 163.367
R893 B.n866 B.n485 163.367
R894 B.n866 B.n483 163.367
R895 B.n870 B.n483 163.367
R896 B.n870 B.n478 163.367
R897 B.n879 B.n478 163.367
R898 B.n879 B.n476 163.367
R899 B.n883 B.n476 163.367
R900 B.n883 B.n470 163.367
R901 B.n891 B.n470 163.367
R902 B.n891 B.n468 163.367
R903 B.n895 B.n468 163.367
R904 B.n895 B.n462 163.367
R905 B.n903 B.n462 163.367
R906 B.n903 B.n460 163.367
R907 B.n907 B.n460 163.367
R908 B.n907 B.n454 163.367
R909 B.n915 B.n454 163.367
R910 B.n915 B.n452 163.367
R911 B.n919 B.n452 163.367
R912 B.n919 B.n446 163.367
R913 B.n927 B.n446 163.367
R914 B.n927 B.n444 163.367
R915 B.n931 B.n444 163.367
R916 B.n931 B.n438 163.367
R917 B.n939 B.n438 163.367
R918 B.n939 B.n436 163.367
R919 B.n943 B.n436 163.367
R920 B.n943 B.n431 163.367
R921 B.n952 B.n431 163.367
R922 B.n952 B.n429 163.367
R923 B.n957 B.n429 163.367
R924 B.n957 B.n423 163.367
R925 B.n965 B.n423 163.367
R926 B.n966 B.n965 163.367
R927 B.n966 B.n5 163.367
R928 B.n6 B.n5 163.367
R929 B.n7 B.n6 163.367
R930 B.n971 B.n7 163.367
R931 B.n971 B.n12 163.367
R932 B.n13 B.n12 163.367
R933 B.n14 B.n13 163.367
R934 B.n976 B.n14 163.367
R935 B.n976 B.n19 163.367
R936 B.n20 B.n19 163.367
R937 B.n21 B.n20 163.367
R938 B.n981 B.n21 163.367
R939 B.n981 B.n26 163.367
R940 B.n27 B.n26 163.367
R941 B.n28 B.n27 163.367
R942 B.n986 B.n28 163.367
R943 B.n986 B.n33 163.367
R944 B.n34 B.n33 163.367
R945 B.n35 B.n34 163.367
R946 B.n991 B.n35 163.367
R947 B.n991 B.n40 163.367
R948 B.n41 B.n40 163.367
R949 B.n42 B.n41 163.367
R950 B.n996 B.n42 163.367
R951 B.n996 B.n47 163.367
R952 B.n48 B.n47 163.367
R953 B.n49 B.n48 163.367
R954 B.n1001 B.n49 163.367
R955 B.n1001 B.n54 163.367
R956 B.n55 B.n54 163.367
R957 B.n56 B.n55 163.367
R958 B.n1006 B.n56 163.367
R959 B.n1006 B.n61 163.367
R960 B.n62 B.n61 163.367
R961 B.n63 B.n62 163.367
R962 B.n1011 B.n63 163.367
R963 B.n1011 B.n68 163.367
R964 B.n69 B.n68 163.367
R965 B.n70 B.n69 163.367
R966 B.n144 B.n70 163.367
R967 B.n150 B.n74 163.367
R968 B.n154 B.n153 163.367
R969 B.n158 B.n157 163.367
R970 B.n162 B.n161 163.367
R971 B.n166 B.n165 163.367
R972 B.n170 B.n169 163.367
R973 B.n174 B.n173 163.367
R974 B.n178 B.n177 163.367
R975 B.n182 B.n181 163.367
R976 B.n186 B.n185 163.367
R977 B.n190 B.n189 163.367
R978 B.n194 B.n193 163.367
R979 B.n198 B.n197 163.367
R980 B.n202 B.n201 163.367
R981 B.n206 B.n205 163.367
R982 B.n210 B.n209 163.367
R983 B.n214 B.n213 163.367
R984 B.n218 B.n217 163.367
R985 B.n222 B.n221 163.367
R986 B.n226 B.n225 163.367
R987 B.n230 B.n229 163.367
R988 B.n234 B.n233 163.367
R989 B.n238 B.n237 163.367
R990 B.n242 B.n241 163.367
R991 B.n246 B.n245 163.367
R992 B.n250 B.n249 163.367
R993 B.n254 B.n253 163.367
R994 B.n258 B.n257 163.367
R995 B.n262 B.n261 163.367
R996 B.n266 B.n265 163.367
R997 B.n270 B.n269 163.367
R998 B.n274 B.n273 163.367
R999 B.n279 B.n278 163.367
R1000 B.n283 B.n282 163.367
R1001 B.n287 B.n286 163.367
R1002 B.n291 B.n290 163.367
R1003 B.n295 B.n294 163.367
R1004 B.n299 B.n298 163.367
R1005 B.n303 B.n302 163.367
R1006 B.n307 B.n306 163.367
R1007 B.n311 B.n310 163.367
R1008 B.n315 B.n314 163.367
R1009 B.n319 B.n318 163.367
R1010 B.n323 B.n322 163.367
R1011 B.n327 B.n326 163.367
R1012 B.n331 B.n330 163.367
R1013 B.n335 B.n334 163.367
R1014 B.n339 B.n338 163.367
R1015 B.n343 B.n342 163.367
R1016 B.n347 B.n346 163.367
R1017 B.n351 B.n350 163.367
R1018 B.n355 B.n354 163.367
R1019 B.n359 B.n358 163.367
R1020 B.n363 B.n362 163.367
R1021 B.n367 B.n366 163.367
R1022 B.n371 B.n370 163.367
R1023 B.n375 B.n374 163.367
R1024 B.n379 B.n378 163.367
R1025 B.n383 B.n382 163.367
R1026 B.n387 B.n386 163.367
R1027 B.n391 B.n390 163.367
R1028 B.n395 B.n394 163.367
R1029 B.n399 B.n398 163.367
R1030 B.n403 B.n402 163.367
R1031 B.n407 B.n406 163.367
R1032 B.n411 B.n410 163.367
R1033 B.n415 B.n414 163.367
R1034 B.n419 B.n418 163.367
R1035 B.n1018 B.n143 163.367
R1036 B.n570 B.t11 139.097
R1037 B.n145 B.t6 139.097
R1038 B.n567 B.t14 139.071
R1039 B.n148 B.t16 139.071
R1040 B.n848 B.n847 71.676
R1041 B.n566 B.n498 71.676
R1042 B.n840 B.n499 71.676
R1043 B.n836 B.n500 71.676
R1044 B.n832 B.n501 71.676
R1045 B.n828 B.n502 71.676
R1046 B.n824 B.n503 71.676
R1047 B.n820 B.n504 71.676
R1048 B.n816 B.n505 71.676
R1049 B.n812 B.n506 71.676
R1050 B.n808 B.n507 71.676
R1051 B.n804 B.n508 71.676
R1052 B.n800 B.n509 71.676
R1053 B.n796 B.n510 71.676
R1054 B.n792 B.n511 71.676
R1055 B.n788 B.n512 71.676
R1056 B.n784 B.n513 71.676
R1057 B.n780 B.n514 71.676
R1058 B.n776 B.n515 71.676
R1059 B.n772 B.n516 71.676
R1060 B.n768 B.n517 71.676
R1061 B.n764 B.n518 71.676
R1062 B.n760 B.n519 71.676
R1063 B.n756 B.n520 71.676
R1064 B.n752 B.n521 71.676
R1065 B.n748 B.n522 71.676
R1066 B.n744 B.n523 71.676
R1067 B.n740 B.n524 71.676
R1068 B.n736 B.n525 71.676
R1069 B.n732 B.n526 71.676
R1070 B.n728 B.n527 71.676
R1071 B.n724 B.n528 71.676
R1072 B.n720 B.n529 71.676
R1073 B.n716 B.n530 71.676
R1074 B.n712 B.n531 71.676
R1075 B.n708 B.n532 71.676
R1076 B.n704 B.n533 71.676
R1077 B.n699 B.n534 71.676
R1078 B.n695 B.n535 71.676
R1079 B.n691 B.n536 71.676
R1080 B.n687 B.n537 71.676
R1081 B.n683 B.n538 71.676
R1082 B.n679 B.n539 71.676
R1083 B.n675 B.n540 71.676
R1084 B.n671 B.n541 71.676
R1085 B.n667 B.n542 71.676
R1086 B.n663 B.n543 71.676
R1087 B.n659 B.n544 71.676
R1088 B.n655 B.n545 71.676
R1089 B.n651 B.n546 71.676
R1090 B.n647 B.n547 71.676
R1091 B.n643 B.n548 71.676
R1092 B.n639 B.n549 71.676
R1093 B.n635 B.n550 71.676
R1094 B.n631 B.n551 71.676
R1095 B.n627 B.n552 71.676
R1096 B.n623 B.n553 71.676
R1097 B.n619 B.n554 71.676
R1098 B.n615 B.n555 71.676
R1099 B.n611 B.n556 71.676
R1100 B.n607 B.n557 71.676
R1101 B.n603 B.n558 71.676
R1102 B.n599 B.n559 71.676
R1103 B.n595 B.n560 71.676
R1104 B.n591 B.n561 71.676
R1105 B.n587 B.n562 71.676
R1106 B.n583 B.n563 71.676
R1107 B.n579 B.n564 71.676
R1108 B.n575 B.n565 71.676
R1109 B.n1021 B.n1020 71.676
R1110 B.n150 B.n75 71.676
R1111 B.n154 B.n76 71.676
R1112 B.n158 B.n77 71.676
R1113 B.n162 B.n78 71.676
R1114 B.n166 B.n79 71.676
R1115 B.n170 B.n80 71.676
R1116 B.n174 B.n81 71.676
R1117 B.n178 B.n82 71.676
R1118 B.n182 B.n83 71.676
R1119 B.n186 B.n84 71.676
R1120 B.n190 B.n85 71.676
R1121 B.n194 B.n86 71.676
R1122 B.n198 B.n87 71.676
R1123 B.n202 B.n88 71.676
R1124 B.n206 B.n89 71.676
R1125 B.n210 B.n90 71.676
R1126 B.n214 B.n91 71.676
R1127 B.n218 B.n92 71.676
R1128 B.n222 B.n93 71.676
R1129 B.n226 B.n94 71.676
R1130 B.n230 B.n95 71.676
R1131 B.n234 B.n96 71.676
R1132 B.n238 B.n97 71.676
R1133 B.n242 B.n98 71.676
R1134 B.n246 B.n99 71.676
R1135 B.n250 B.n100 71.676
R1136 B.n254 B.n101 71.676
R1137 B.n258 B.n102 71.676
R1138 B.n262 B.n103 71.676
R1139 B.n266 B.n104 71.676
R1140 B.n270 B.n105 71.676
R1141 B.n274 B.n106 71.676
R1142 B.n279 B.n107 71.676
R1143 B.n283 B.n108 71.676
R1144 B.n287 B.n109 71.676
R1145 B.n291 B.n110 71.676
R1146 B.n295 B.n111 71.676
R1147 B.n299 B.n112 71.676
R1148 B.n303 B.n113 71.676
R1149 B.n307 B.n114 71.676
R1150 B.n311 B.n115 71.676
R1151 B.n315 B.n116 71.676
R1152 B.n319 B.n117 71.676
R1153 B.n323 B.n118 71.676
R1154 B.n327 B.n119 71.676
R1155 B.n331 B.n120 71.676
R1156 B.n335 B.n121 71.676
R1157 B.n339 B.n122 71.676
R1158 B.n343 B.n123 71.676
R1159 B.n347 B.n124 71.676
R1160 B.n351 B.n125 71.676
R1161 B.n355 B.n126 71.676
R1162 B.n359 B.n127 71.676
R1163 B.n363 B.n128 71.676
R1164 B.n367 B.n129 71.676
R1165 B.n371 B.n130 71.676
R1166 B.n375 B.n131 71.676
R1167 B.n379 B.n132 71.676
R1168 B.n383 B.n133 71.676
R1169 B.n387 B.n134 71.676
R1170 B.n391 B.n135 71.676
R1171 B.n395 B.n136 71.676
R1172 B.n399 B.n137 71.676
R1173 B.n403 B.n138 71.676
R1174 B.n407 B.n139 71.676
R1175 B.n411 B.n140 71.676
R1176 B.n415 B.n141 71.676
R1177 B.n419 B.n142 71.676
R1178 B.n143 B.n142 71.676
R1179 B.n418 B.n141 71.676
R1180 B.n414 B.n140 71.676
R1181 B.n410 B.n139 71.676
R1182 B.n406 B.n138 71.676
R1183 B.n402 B.n137 71.676
R1184 B.n398 B.n136 71.676
R1185 B.n394 B.n135 71.676
R1186 B.n390 B.n134 71.676
R1187 B.n386 B.n133 71.676
R1188 B.n382 B.n132 71.676
R1189 B.n378 B.n131 71.676
R1190 B.n374 B.n130 71.676
R1191 B.n370 B.n129 71.676
R1192 B.n366 B.n128 71.676
R1193 B.n362 B.n127 71.676
R1194 B.n358 B.n126 71.676
R1195 B.n354 B.n125 71.676
R1196 B.n350 B.n124 71.676
R1197 B.n346 B.n123 71.676
R1198 B.n342 B.n122 71.676
R1199 B.n338 B.n121 71.676
R1200 B.n334 B.n120 71.676
R1201 B.n330 B.n119 71.676
R1202 B.n326 B.n118 71.676
R1203 B.n322 B.n117 71.676
R1204 B.n318 B.n116 71.676
R1205 B.n314 B.n115 71.676
R1206 B.n310 B.n114 71.676
R1207 B.n306 B.n113 71.676
R1208 B.n302 B.n112 71.676
R1209 B.n298 B.n111 71.676
R1210 B.n294 B.n110 71.676
R1211 B.n290 B.n109 71.676
R1212 B.n286 B.n108 71.676
R1213 B.n282 B.n107 71.676
R1214 B.n278 B.n106 71.676
R1215 B.n273 B.n105 71.676
R1216 B.n269 B.n104 71.676
R1217 B.n265 B.n103 71.676
R1218 B.n261 B.n102 71.676
R1219 B.n257 B.n101 71.676
R1220 B.n253 B.n100 71.676
R1221 B.n249 B.n99 71.676
R1222 B.n245 B.n98 71.676
R1223 B.n241 B.n97 71.676
R1224 B.n237 B.n96 71.676
R1225 B.n233 B.n95 71.676
R1226 B.n229 B.n94 71.676
R1227 B.n225 B.n93 71.676
R1228 B.n221 B.n92 71.676
R1229 B.n217 B.n91 71.676
R1230 B.n213 B.n90 71.676
R1231 B.n209 B.n89 71.676
R1232 B.n205 B.n88 71.676
R1233 B.n201 B.n87 71.676
R1234 B.n197 B.n86 71.676
R1235 B.n193 B.n85 71.676
R1236 B.n189 B.n84 71.676
R1237 B.n185 B.n83 71.676
R1238 B.n181 B.n82 71.676
R1239 B.n177 B.n81 71.676
R1240 B.n173 B.n80 71.676
R1241 B.n169 B.n79 71.676
R1242 B.n165 B.n78 71.676
R1243 B.n161 B.n77 71.676
R1244 B.n157 B.n76 71.676
R1245 B.n153 B.n75 71.676
R1246 B.n1020 B.n74 71.676
R1247 B.n847 B.n497 71.676
R1248 B.n841 B.n498 71.676
R1249 B.n837 B.n499 71.676
R1250 B.n833 B.n500 71.676
R1251 B.n829 B.n501 71.676
R1252 B.n825 B.n502 71.676
R1253 B.n821 B.n503 71.676
R1254 B.n817 B.n504 71.676
R1255 B.n813 B.n505 71.676
R1256 B.n809 B.n506 71.676
R1257 B.n805 B.n507 71.676
R1258 B.n801 B.n508 71.676
R1259 B.n797 B.n509 71.676
R1260 B.n793 B.n510 71.676
R1261 B.n789 B.n511 71.676
R1262 B.n785 B.n512 71.676
R1263 B.n781 B.n513 71.676
R1264 B.n777 B.n514 71.676
R1265 B.n773 B.n515 71.676
R1266 B.n769 B.n516 71.676
R1267 B.n765 B.n517 71.676
R1268 B.n761 B.n518 71.676
R1269 B.n757 B.n519 71.676
R1270 B.n753 B.n520 71.676
R1271 B.n749 B.n521 71.676
R1272 B.n745 B.n522 71.676
R1273 B.n741 B.n523 71.676
R1274 B.n737 B.n524 71.676
R1275 B.n733 B.n525 71.676
R1276 B.n729 B.n526 71.676
R1277 B.n725 B.n527 71.676
R1278 B.n721 B.n528 71.676
R1279 B.n717 B.n529 71.676
R1280 B.n713 B.n530 71.676
R1281 B.n709 B.n531 71.676
R1282 B.n705 B.n532 71.676
R1283 B.n700 B.n533 71.676
R1284 B.n696 B.n534 71.676
R1285 B.n692 B.n535 71.676
R1286 B.n688 B.n536 71.676
R1287 B.n684 B.n537 71.676
R1288 B.n680 B.n538 71.676
R1289 B.n676 B.n539 71.676
R1290 B.n672 B.n540 71.676
R1291 B.n668 B.n541 71.676
R1292 B.n664 B.n542 71.676
R1293 B.n660 B.n543 71.676
R1294 B.n656 B.n544 71.676
R1295 B.n652 B.n545 71.676
R1296 B.n648 B.n546 71.676
R1297 B.n644 B.n547 71.676
R1298 B.n640 B.n548 71.676
R1299 B.n636 B.n549 71.676
R1300 B.n632 B.n550 71.676
R1301 B.n628 B.n551 71.676
R1302 B.n624 B.n552 71.676
R1303 B.n620 B.n553 71.676
R1304 B.n616 B.n554 71.676
R1305 B.n612 B.n555 71.676
R1306 B.n608 B.n556 71.676
R1307 B.n604 B.n557 71.676
R1308 B.n600 B.n558 71.676
R1309 B.n596 B.n559 71.676
R1310 B.n592 B.n560 71.676
R1311 B.n588 B.n561 71.676
R1312 B.n584 B.n562 71.676
R1313 B.n580 B.n563 71.676
R1314 B.n576 B.n564 71.676
R1315 B.n572 B.n565 71.676
R1316 B.n571 B.t10 70.6373
R1317 B.n146 B.t7 70.6373
R1318 B.n568 B.t13 70.6105
R1319 B.n149 B.t17 70.6105
R1320 B.n571 B.n570 68.4611
R1321 B.n568 B.n567 68.4611
R1322 B.n149 B.n148 68.4611
R1323 B.n146 B.n145 68.4611
R1324 B.n846 B.n494 61.6092
R1325 B.n1019 B.n71 61.6092
R1326 B.n702 B.n571 59.5399
R1327 B.n569 B.n568 59.5399
R1328 B.n276 B.n149 59.5399
R1329 B.n147 B.n146 59.5399
R1330 B.n1023 B.n1022 36.6834
R1331 B.n1017 B.n1016 36.6834
R1332 B.n573 B.n492 36.6834
R1333 B.n850 B.n849 36.6834
R1334 B.n853 B.n494 29.7125
R1335 B.n853 B.n490 29.7125
R1336 B.n859 B.n490 29.7125
R1337 B.n859 B.n486 29.7125
R1338 B.n865 B.n486 29.7125
R1339 B.n865 B.n482 29.7125
R1340 B.n872 B.n482 29.7125
R1341 B.n872 B.n871 29.7125
R1342 B.n878 B.n475 29.7125
R1343 B.n884 B.n475 29.7125
R1344 B.n884 B.n471 29.7125
R1345 B.n890 B.n471 29.7125
R1346 B.n890 B.n467 29.7125
R1347 B.n896 B.n467 29.7125
R1348 B.n896 B.n463 29.7125
R1349 B.n902 B.n463 29.7125
R1350 B.n902 B.n459 29.7125
R1351 B.n908 B.n459 29.7125
R1352 B.n908 B.n455 29.7125
R1353 B.n914 B.n455 29.7125
R1354 B.n920 B.n451 29.7125
R1355 B.n920 B.n447 29.7125
R1356 B.n926 B.n447 29.7125
R1357 B.n926 B.n443 29.7125
R1358 B.n932 B.n443 29.7125
R1359 B.n932 B.n439 29.7125
R1360 B.n938 B.n439 29.7125
R1361 B.n938 B.n435 29.7125
R1362 B.n945 B.n435 29.7125
R1363 B.n945 B.n944 29.7125
R1364 B.n951 B.n428 29.7125
R1365 B.n958 B.n428 29.7125
R1366 B.n958 B.n424 29.7125
R1367 B.n964 B.n424 29.7125
R1368 B.n964 B.n4 29.7125
R1369 B.n1100 B.n4 29.7125
R1370 B.n1100 B.n1099 29.7125
R1371 B.n1099 B.n1098 29.7125
R1372 B.n1098 B.n8 29.7125
R1373 B.n1092 B.n8 29.7125
R1374 B.n1092 B.n1091 29.7125
R1375 B.n1091 B.n1090 29.7125
R1376 B.n1084 B.n18 29.7125
R1377 B.n1084 B.n1083 29.7125
R1378 B.n1083 B.n1082 29.7125
R1379 B.n1082 B.n22 29.7125
R1380 B.n1076 B.n22 29.7125
R1381 B.n1076 B.n1075 29.7125
R1382 B.n1075 B.n1074 29.7125
R1383 B.n1074 B.n29 29.7125
R1384 B.n1068 B.n29 29.7125
R1385 B.n1068 B.n1067 29.7125
R1386 B.n1066 B.n36 29.7125
R1387 B.n1060 B.n36 29.7125
R1388 B.n1060 B.n1059 29.7125
R1389 B.n1059 B.n1058 29.7125
R1390 B.n1058 B.n43 29.7125
R1391 B.n1052 B.n43 29.7125
R1392 B.n1052 B.n1051 29.7125
R1393 B.n1051 B.n1050 29.7125
R1394 B.n1050 B.n50 29.7125
R1395 B.n1044 B.n50 29.7125
R1396 B.n1044 B.n1043 29.7125
R1397 B.n1043 B.n1042 29.7125
R1398 B.n1036 B.n60 29.7125
R1399 B.n1036 B.n1035 29.7125
R1400 B.n1035 B.n1034 29.7125
R1401 B.n1034 B.n64 29.7125
R1402 B.n1028 B.n64 29.7125
R1403 B.n1028 B.n1027 29.7125
R1404 B.n1027 B.n1026 29.7125
R1405 B.n1026 B.n71 29.7125
R1406 B.n914 B.t0 24.4692
R1407 B.t1 B.n1066 24.4692
R1408 B.n951 B.t2 23.5953
R1409 B.n1090 B.t3 23.5953
R1410 B.n878 B.t9 22.7215
R1411 B.n1042 B.t5 22.7215
R1412 B B.n1102 18.0485
R1413 B.n1022 B.n73 10.6151
R1414 B.n151 B.n73 10.6151
R1415 B.n152 B.n151 10.6151
R1416 B.n155 B.n152 10.6151
R1417 B.n156 B.n155 10.6151
R1418 B.n159 B.n156 10.6151
R1419 B.n160 B.n159 10.6151
R1420 B.n163 B.n160 10.6151
R1421 B.n164 B.n163 10.6151
R1422 B.n167 B.n164 10.6151
R1423 B.n168 B.n167 10.6151
R1424 B.n171 B.n168 10.6151
R1425 B.n172 B.n171 10.6151
R1426 B.n175 B.n172 10.6151
R1427 B.n176 B.n175 10.6151
R1428 B.n179 B.n176 10.6151
R1429 B.n180 B.n179 10.6151
R1430 B.n183 B.n180 10.6151
R1431 B.n184 B.n183 10.6151
R1432 B.n187 B.n184 10.6151
R1433 B.n188 B.n187 10.6151
R1434 B.n191 B.n188 10.6151
R1435 B.n192 B.n191 10.6151
R1436 B.n195 B.n192 10.6151
R1437 B.n196 B.n195 10.6151
R1438 B.n199 B.n196 10.6151
R1439 B.n200 B.n199 10.6151
R1440 B.n203 B.n200 10.6151
R1441 B.n204 B.n203 10.6151
R1442 B.n207 B.n204 10.6151
R1443 B.n208 B.n207 10.6151
R1444 B.n211 B.n208 10.6151
R1445 B.n212 B.n211 10.6151
R1446 B.n215 B.n212 10.6151
R1447 B.n216 B.n215 10.6151
R1448 B.n219 B.n216 10.6151
R1449 B.n220 B.n219 10.6151
R1450 B.n223 B.n220 10.6151
R1451 B.n224 B.n223 10.6151
R1452 B.n227 B.n224 10.6151
R1453 B.n228 B.n227 10.6151
R1454 B.n231 B.n228 10.6151
R1455 B.n232 B.n231 10.6151
R1456 B.n235 B.n232 10.6151
R1457 B.n236 B.n235 10.6151
R1458 B.n239 B.n236 10.6151
R1459 B.n240 B.n239 10.6151
R1460 B.n243 B.n240 10.6151
R1461 B.n244 B.n243 10.6151
R1462 B.n247 B.n244 10.6151
R1463 B.n248 B.n247 10.6151
R1464 B.n251 B.n248 10.6151
R1465 B.n252 B.n251 10.6151
R1466 B.n255 B.n252 10.6151
R1467 B.n256 B.n255 10.6151
R1468 B.n259 B.n256 10.6151
R1469 B.n260 B.n259 10.6151
R1470 B.n263 B.n260 10.6151
R1471 B.n264 B.n263 10.6151
R1472 B.n267 B.n264 10.6151
R1473 B.n268 B.n267 10.6151
R1474 B.n271 B.n268 10.6151
R1475 B.n272 B.n271 10.6151
R1476 B.n275 B.n272 10.6151
R1477 B.n280 B.n277 10.6151
R1478 B.n281 B.n280 10.6151
R1479 B.n284 B.n281 10.6151
R1480 B.n285 B.n284 10.6151
R1481 B.n288 B.n285 10.6151
R1482 B.n289 B.n288 10.6151
R1483 B.n292 B.n289 10.6151
R1484 B.n293 B.n292 10.6151
R1485 B.n297 B.n296 10.6151
R1486 B.n300 B.n297 10.6151
R1487 B.n301 B.n300 10.6151
R1488 B.n304 B.n301 10.6151
R1489 B.n305 B.n304 10.6151
R1490 B.n308 B.n305 10.6151
R1491 B.n309 B.n308 10.6151
R1492 B.n312 B.n309 10.6151
R1493 B.n313 B.n312 10.6151
R1494 B.n316 B.n313 10.6151
R1495 B.n317 B.n316 10.6151
R1496 B.n320 B.n317 10.6151
R1497 B.n321 B.n320 10.6151
R1498 B.n324 B.n321 10.6151
R1499 B.n325 B.n324 10.6151
R1500 B.n328 B.n325 10.6151
R1501 B.n329 B.n328 10.6151
R1502 B.n332 B.n329 10.6151
R1503 B.n333 B.n332 10.6151
R1504 B.n336 B.n333 10.6151
R1505 B.n337 B.n336 10.6151
R1506 B.n340 B.n337 10.6151
R1507 B.n341 B.n340 10.6151
R1508 B.n344 B.n341 10.6151
R1509 B.n345 B.n344 10.6151
R1510 B.n348 B.n345 10.6151
R1511 B.n349 B.n348 10.6151
R1512 B.n352 B.n349 10.6151
R1513 B.n353 B.n352 10.6151
R1514 B.n356 B.n353 10.6151
R1515 B.n357 B.n356 10.6151
R1516 B.n360 B.n357 10.6151
R1517 B.n361 B.n360 10.6151
R1518 B.n364 B.n361 10.6151
R1519 B.n365 B.n364 10.6151
R1520 B.n368 B.n365 10.6151
R1521 B.n369 B.n368 10.6151
R1522 B.n372 B.n369 10.6151
R1523 B.n373 B.n372 10.6151
R1524 B.n376 B.n373 10.6151
R1525 B.n377 B.n376 10.6151
R1526 B.n380 B.n377 10.6151
R1527 B.n381 B.n380 10.6151
R1528 B.n384 B.n381 10.6151
R1529 B.n385 B.n384 10.6151
R1530 B.n388 B.n385 10.6151
R1531 B.n389 B.n388 10.6151
R1532 B.n392 B.n389 10.6151
R1533 B.n393 B.n392 10.6151
R1534 B.n396 B.n393 10.6151
R1535 B.n397 B.n396 10.6151
R1536 B.n400 B.n397 10.6151
R1537 B.n401 B.n400 10.6151
R1538 B.n404 B.n401 10.6151
R1539 B.n405 B.n404 10.6151
R1540 B.n408 B.n405 10.6151
R1541 B.n409 B.n408 10.6151
R1542 B.n412 B.n409 10.6151
R1543 B.n413 B.n412 10.6151
R1544 B.n416 B.n413 10.6151
R1545 B.n417 B.n416 10.6151
R1546 B.n420 B.n417 10.6151
R1547 B.n421 B.n420 10.6151
R1548 B.n1017 B.n421 10.6151
R1549 B.n855 B.n492 10.6151
R1550 B.n856 B.n855 10.6151
R1551 B.n857 B.n856 10.6151
R1552 B.n857 B.n484 10.6151
R1553 B.n867 B.n484 10.6151
R1554 B.n868 B.n867 10.6151
R1555 B.n869 B.n868 10.6151
R1556 B.n869 B.n477 10.6151
R1557 B.n880 B.n477 10.6151
R1558 B.n881 B.n880 10.6151
R1559 B.n882 B.n881 10.6151
R1560 B.n882 B.n469 10.6151
R1561 B.n892 B.n469 10.6151
R1562 B.n893 B.n892 10.6151
R1563 B.n894 B.n893 10.6151
R1564 B.n894 B.n461 10.6151
R1565 B.n904 B.n461 10.6151
R1566 B.n905 B.n904 10.6151
R1567 B.n906 B.n905 10.6151
R1568 B.n906 B.n453 10.6151
R1569 B.n916 B.n453 10.6151
R1570 B.n917 B.n916 10.6151
R1571 B.n918 B.n917 10.6151
R1572 B.n918 B.n445 10.6151
R1573 B.n928 B.n445 10.6151
R1574 B.n929 B.n928 10.6151
R1575 B.n930 B.n929 10.6151
R1576 B.n930 B.n437 10.6151
R1577 B.n940 B.n437 10.6151
R1578 B.n941 B.n940 10.6151
R1579 B.n942 B.n941 10.6151
R1580 B.n942 B.n430 10.6151
R1581 B.n953 B.n430 10.6151
R1582 B.n954 B.n953 10.6151
R1583 B.n956 B.n954 10.6151
R1584 B.n956 B.n955 10.6151
R1585 B.n955 B.n422 10.6151
R1586 B.n967 B.n422 10.6151
R1587 B.n968 B.n967 10.6151
R1588 B.n969 B.n968 10.6151
R1589 B.n970 B.n969 10.6151
R1590 B.n972 B.n970 10.6151
R1591 B.n973 B.n972 10.6151
R1592 B.n974 B.n973 10.6151
R1593 B.n975 B.n974 10.6151
R1594 B.n977 B.n975 10.6151
R1595 B.n978 B.n977 10.6151
R1596 B.n979 B.n978 10.6151
R1597 B.n980 B.n979 10.6151
R1598 B.n982 B.n980 10.6151
R1599 B.n983 B.n982 10.6151
R1600 B.n984 B.n983 10.6151
R1601 B.n985 B.n984 10.6151
R1602 B.n987 B.n985 10.6151
R1603 B.n988 B.n987 10.6151
R1604 B.n989 B.n988 10.6151
R1605 B.n990 B.n989 10.6151
R1606 B.n992 B.n990 10.6151
R1607 B.n993 B.n992 10.6151
R1608 B.n994 B.n993 10.6151
R1609 B.n995 B.n994 10.6151
R1610 B.n997 B.n995 10.6151
R1611 B.n998 B.n997 10.6151
R1612 B.n999 B.n998 10.6151
R1613 B.n1000 B.n999 10.6151
R1614 B.n1002 B.n1000 10.6151
R1615 B.n1003 B.n1002 10.6151
R1616 B.n1004 B.n1003 10.6151
R1617 B.n1005 B.n1004 10.6151
R1618 B.n1007 B.n1005 10.6151
R1619 B.n1008 B.n1007 10.6151
R1620 B.n1009 B.n1008 10.6151
R1621 B.n1010 B.n1009 10.6151
R1622 B.n1012 B.n1010 10.6151
R1623 B.n1013 B.n1012 10.6151
R1624 B.n1014 B.n1013 10.6151
R1625 B.n1015 B.n1014 10.6151
R1626 B.n1016 B.n1015 10.6151
R1627 B.n849 B.n496 10.6151
R1628 B.n844 B.n496 10.6151
R1629 B.n844 B.n843 10.6151
R1630 B.n843 B.n842 10.6151
R1631 B.n842 B.n839 10.6151
R1632 B.n839 B.n838 10.6151
R1633 B.n838 B.n835 10.6151
R1634 B.n835 B.n834 10.6151
R1635 B.n834 B.n831 10.6151
R1636 B.n831 B.n830 10.6151
R1637 B.n830 B.n827 10.6151
R1638 B.n827 B.n826 10.6151
R1639 B.n826 B.n823 10.6151
R1640 B.n823 B.n822 10.6151
R1641 B.n822 B.n819 10.6151
R1642 B.n819 B.n818 10.6151
R1643 B.n818 B.n815 10.6151
R1644 B.n815 B.n814 10.6151
R1645 B.n814 B.n811 10.6151
R1646 B.n811 B.n810 10.6151
R1647 B.n810 B.n807 10.6151
R1648 B.n807 B.n806 10.6151
R1649 B.n806 B.n803 10.6151
R1650 B.n803 B.n802 10.6151
R1651 B.n802 B.n799 10.6151
R1652 B.n799 B.n798 10.6151
R1653 B.n798 B.n795 10.6151
R1654 B.n795 B.n794 10.6151
R1655 B.n794 B.n791 10.6151
R1656 B.n791 B.n790 10.6151
R1657 B.n790 B.n787 10.6151
R1658 B.n787 B.n786 10.6151
R1659 B.n786 B.n783 10.6151
R1660 B.n783 B.n782 10.6151
R1661 B.n782 B.n779 10.6151
R1662 B.n779 B.n778 10.6151
R1663 B.n778 B.n775 10.6151
R1664 B.n775 B.n774 10.6151
R1665 B.n774 B.n771 10.6151
R1666 B.n771 B.n770 10.6151
R1667 B.n770 B.n767 10.6151
R1668 B.n767 B.n766 10.6151
R1669 B.n766 B.n763 10.6151
R1670 B.n763 B.n762 10.6151
R1671 B.n762 B.n759 10.6151
R1672 B.n759 B.n758 10.6151
R1673 B.n758 B.n755 10.6151
R1674 B.n755 B.n754 10.6151
R1675 B.n754 B.n751 10.6151
R1676 B.n751 B.n750 10.6151
R1677 B.n750 B.n747 10.6151
R1678 B.n747 B.n746 10.6151
R1679 B.n746 B.n743 10.6151
R1680 B.n743 B.n742 10.6151
R1681 B.n742 B.n739 10.6151
R1682 B.n739 B.n738 10.6151
R1683 B.n738 B.n735 10.6151
R1684 B.n735 B.n734 10.6151
R1685 B.n734 B.n731 10.6151
R1686 B.n731 B.n730 10.6151
R1687 B.n730 B.n727 10.6151
R1688 B.n727 B.n726 10.6151
R1689 B.n726 B.n723 10.6151
R1690 B.n723 B.n722 10.6151
R1691 B.n719 B.n718 10.6151
R1692 B.n718 B.n715 10.6151
R1693 B.n715 B.n714 10.6151
R1694 B.n714 B.n711 10.6151
R1695 B.n711 B.n710 10.6151
R1696 B.n710 B.n707 10.6151
R1697 B.n707 B.n706 10.6151
R1698 B.n706 B.n703 10.6151
R1699 B.n701 B.n698 10.6151
R1700 B.n698 B.n697 10.6151
R1701 B.n697 B.n694 10.6151
R1702 B.n694 B.n693 10.6151
R1703 B.n693 B.n690 10.6151
R1704 B.n690 B.n689 10.6151
R1705 B.n689 B.n686 10.6151
R1706 B.n686 B.n685 10.6151
R1707 B.n685 B.n682 10.6151
R1708 B.n682 B.n681 10.6151
R1709 B.n681 B.n678 10.6151
R1710 B.n678 B.n677 10.6151
R1711 B.n677 B.n674 10.6151
R1712 B.n674 B.n673 10.6151
R1713 B.n673 B.n670 10.6151
R1714 B.n670 B.n669 10.6151
R1715 B.n669 B.n666 10.6151
R1716 B.n666 B.n665 10.6151
R1717 B.n665 B.n662 10.6151
R1718 B.n662 B.n661 10.6151
R1719 B.n661 B.n658 10.6151
R1720 B.n658 B.n657 10.6151
R1721 B.n657 B.n654 10.6151
R1722 B.n654 B.n653 10.6151
R1723 B.n653 B.n650 10.6151
R1724 B.n650 B.n649 10.6151
R1725 B.n649 B.n646 10.6151
R1726 B.n646 B.n645 10.6151
R1727 B.n645 B.n642 10.6151
R1728 B.n642 B.n641 10.6151
R1729 B.n641 B.n638 10.6151
R1730 B.n638 B.n637 10.6151
R1731 B.n637 B.n634 10.6151
R1732 B.n634 B.n633 10.6151
R1733 B.n633 B.n630 10.6151
R1734 B.n630 B.n629 10.6151
R1735 B.n629 B.n626 10.6151
R1736 B.n626 B.n625 10.6151
R1737 B.n625 B.n622 10.6151
R1738 B.n622 B.n621 10.6151
R1739 B.n621 B.n618 10.6151
R1740 B.n618 B.n617 10.6151
R1741 B.n617 B.n614 10.6151
R1742 B.n614 B.n613 10.6151
R1743 B.n613 B.n610 10.6151
R1744 B.n610 B.n609 10.6151
R1745 B.n609 B.n606 10.6151
R1746 B.n606 B.n605 10.6151
R1747 B.n605 B.n602 10.6151
R1748 B.n602 B.n601 10.6151
R1749 B.n601 B.n598 10.6151
R1750 B.n598 B.n597 10.6151
R1751 B.n597 B.n594 10.6151
R1752 B.n594 B.n593 10.6151
R1753 B.n593 B.n590 10.6151
R1754 B.n590 B.n589 10.6151
R1755 B.n589 B.n586 10.6151
R1756 B.n586 B.n585 10.6151
R1757 B.n585 B.n582 10.6151
R1758 B.n582 B.n581 10.6151
R1759 B.n581 B.n578 10.6151
R1760 B.n578 B.n577 10.6151
R1761 B.n577 B.n574 10.6151
R1762 B.n574 B.n573 10.6151
R1763 B.n851 B.n850 10.6151
R1764 B.n851 B.n488 10.6151
R1765 B.n861 B.n488 10.6151
R1766 B.n862 B.n861 10.6151
R1767 B.n863 B.n862 10.6151
R1768 B.n863 B.n480 10.6151
R1769 B.n874 B.n480 10.6151
R1770 B.n875 B.n874 10.6151
R1771 B.n876 B.n875 10.6151
R1772 B.n876 B.n473 10.6151
R1773 B.n886 B.n473 10.6151
R1774 B.n887 B.n886 10.6151
R1775 B.n888 B.n887 10.6151
R1776 B.n888 B.n465 10.6151
R1777 B.n898 B.n465 10.6151
R1778 B.n899 B.n898 10.6151
R1779 B.n900 B.n899 10.6151
R1780 B.n900 B.n457 10.6151
R1781 B.n910 B.n457 10.6151
R1782 B.n911 B.n910 10.6151
R1783 B.n912 B.n911 10.6151
R1784 B.n912 B.n449 10.6151
R1785 B.n922 B.n449 10.6151
R1786 B.n923 B.n922 10.6151
R1787 B.n924 B.n923 10.6151
R1788 B.n924 B.n441 10.6151
R1789 B.n934 B.n441 10.6151
R1790 B.n935 B.n934 10.6151
R1791 B.n936 B.n935 10.6151
R1792 B.n936 B.n433 10.6151
R1793 B.n947 B.n433 10.6151
R1794 B.n948 B.n947 10.6151
R1795 B.n949 B.n948 10.6151
R1796 B.n949 B.n426 10.6151
R1797 B.n960 B.n426 10.6151
R1798 B.n961 B.n960 10.6151
R1799 B.n962 B.n961 10.6151
R1800 B.n962 B.n0 10.6151
R1801 B.n1096 B.n1 10.6151
R1802 B.n1096 B.n1095 10.6151
R1803 B.n1095 B.n1094 10.6151
R1804 B.n1094 B.n10 10.6151
R1805 B.n1088 B.n10 10.6151
R1806 B.n1088 B.n1087 10.6151
R1807 B.n1087 B.n1086 10.6151
R1808 B.n1086 B.n16 10.6151
R1809 B.n1080 B.n16 10.6151
R1810 B.n1080 B.n1079 10.6151
R1811 B.n1079 B.n1078 10.6151
R1812 B.n1078 B.n24 10.6151
R1813 B.n1072 B.n24 10.6151
R1814 B.n1072 B.n1071 10.6151
R1815 B.n1071 B.n1070 10.6151
R1816 B.n1070 B.n31 10.6151
R1817 B.n1064 B.n31 10.6151
R1818 B.n1064 B.n1063 10.6151
R1819 B.n1063 B.n1062 10.6151
R1820 B.n1062 B.n38 10.6151
R1821 B.n1056 B.n38 10.6151
R1822 B.n1056 B.n1055 10.6151
R1823 B.n1055 B.n1054 10.6151
R1824 B.n1054 B.n45 10.6151
R1825 B.n1048 B.n45 10.6151
R1826 B.n1048 B.n1047 10.6151
R1827 B.n1047 B.n1046 10.6151
R1828 B.n1046 B.n52 10.6151
R1829 B.n1040 B.n52 10.6151
R1830 B.n1040 B.n1039 10.6151
R1831 B.n1039 B.n1038 10.6151
R1832 B.n1038 B.n58 10.6151
R1833 B.n1032 B.n58 10.6151
R1834 B.n1032 B.n1031 10.6151
R1835 B.n1031 B.n1030 10.6151
R1836 B.n1030 B.n66 10.6151
R1837 B.n1024 B.n66 10.6151
R1838 B.n1024 B.n1023 10.6151
R1839 B.n871 B.t9 6.99156
R1840 B.n60 B.t5 6.99156
R1841 B.n277 B.n276 6.5566
R1842 B.n293 B.n147 6.5566
R1843 B.n719 B.n569 6.5566
R1844 B.n703 B.n702 6.5566
R1845 B.n944 B.t2 6.11768
R1846 B.n18 B.t3 6.11768
R1847 B.t0 B.n451 5.2438
R1848 B.n1067 B.t1 5.2438
R1849 B.n276 B.n275 4.05904
R1850 B.n296 B.n147 4.05904
R1851 B.n722 B.n569 4.05904
R1852 B.n702 B.n701 4.05904
R1853 B.n1102 B.n0 2.81026
R1854 B.n1102 B.n1 2.81026
R1855 VP.n5 VP.t3 184.6
R1856 VP.n5 VP.t1 183.504
R1857 VP.n17 VP.n16 161.3
R1858 VP.n15 VP.n1 161.3
R1859 VP.n14 VP.n13 161.3
R1860 VP.n12 VP.n2 161.3
R1861 VP.n11 VP.n10 161.3
R1862 VP.n9 VP.n3 161.3
R1863 VP.n8 VP.n7 161.3
R1864 VP.n4 VP.t0 149.873
R1865 VP.n0 VP.t2 149.873
R1866 VP.n6 VP.n4 77.2119
R1867 VP.n18 VP.n0 77.2119
R1868 VP.n6 VP.n5 56.7471
R1869 VP.n10 VP.n2 40.577
R1870 VP.n14 VP.n2 40.577
R1871 VP.n9 VP.n8 24.5923
R1872 VP.n10 VP.n9 24.5923
R1873 VP.n15 VP.n14 24.5923
R1874 VP.n16 VP.n15 24.5923
R1875 VP.n8 VP.n4 13.0342
R1876 VP.n16 VP.n0 13.0342
R1877 VP.n7 VP.n6 0.354861
R1878 VP.n18 VP.n17 0.354861
R1879 VP VP.n18 0.267071
R1880 VP.n7 VP.n3 0.189894
R1881 VP.n11 VP.n3 0.189894
R1882 VP.n12 VP.n11 0.189894
R1883 VP.n13 VP.n12 0.189894
R1884 VP.n13 VP.n1 0.189894
R1885 VP.n17 VP.n1 0.189894
R1886 VDD1 VDD1.n1 114.996
R1887 VDD1 VDD1.n0 64.5295
R1888 VDD1.n0 VDD1.t0 0.995475
R1889 VDD1.n0 VDD1.t1 0.995475
R1890 VDD1.n1 VDD1.t3 0.995475
R1891 VDD1.n1 VDD1.t2 0.995475
R1892 VTAIL.n5 VTAIL.t4 48.7877
R1893 VTAIL.n4 VTAIL.t2 48.7877
R1894 VTAIL.n3 VTAIL.t1 48.7877
R1895 VTAIL.n7 VTAIL.t0 48.7875
R1896 VTAIL.n0 VTAIL.t3 48.7875
R1897 VTAIL.n1 VTAIL.t5 48.7875
R1898 VTAIL.n2 VTAIL.t7 48.7875
R1899 VTAIL.n6 VTAIL.t6 48.7875
R1900 VTAIL.n7 VTAIL.n6 32.5652
R1901 VTAIL.n3 VTAIL.n2 32.5652
R1902 VTAIL.n4 VTAIL.n3 3.0436
R1903 VTAIL.n6 VTAIL.n5 3.0436
R1904 VTAIL.n2 VTAIL.n1 3.0436
R1905 VTAIL VTAIL.n0 1.58024
R1906 VTAIL VTAIL.n7 1.46386
R1907 VTAIL.n5 VTAIL.n4 0.470328
R1908 VTAIL.n1 VTAIL.n0 0.470328
R1909 VN.n1 VN.t2 184.6
R1910 VN.n0 VN.t0 184.6
R1911 VN.n0 VN.t3 183.504
R1912 VN.n1 VN.t1 183.504
R1913 VN VN.n1 56.9124
R1914 VN VN.n0 2.61312
R1915 VDD2.n2 VDD2.n0 114.471
R1916 VDD2.n2 VDD2.n1 64.4713
R1917 VDD2.n1 VDD2.t2 0.995475
R1918 VDD2.n1 VDD2.t1 0.995475
R1919 VDD2.n0 VDD2.t3 0.995475
R1920 VDD2.n0 VDD2.t0 0.995475
R1921 VDD2 VDD2.n2 0.0586897
C0 VN VTAIL 7.57529f
C1 VDD2 VTAIL 7.3437f
C2 VDD1 VP 8.225241f
C3 VP VTAIL 7.5894f
C4 VDD2 VN 7.94318f
C5 VDD1 VTAIL 7.28547f
C6 VP VN 8.085381f
C7 VDD2 VP 0.432663f
C8 VDD1 VN 0.149721f
C9 VDD2 VDD1 1.17282f
C10 VDD2 B 4.712392f
C11 VDD1 B 9.864051f
C12 VTAIL B 15.195141f
C13 VN B 12.49422f
C14 VP B 10.757277f
C15 VDD2.t3 B 0.414625f
C16 VDD2.t0 B 0.414625f
C17 VDD2.n0 B 4.76587f
C18 VDD2.t2 B 0.414625f
C19 VDD2.t1 B 0.414625f
C20 VDD2.n1 B 3.80176f
C21 VDD2.n2 B 4.709661f
C22 VN.t3 B 3.9011f
C23 VN.t0 B 3.90921f
C24 VN.n0 B 2.44143f
C25 VN.t1 B 3.9011f
C26 VN.t2 B 3.90921f
C27 VN.n1 B 3.91204f
C28 VTAIL.t3 B 2.76651f
C29 VTAIL.n0 B 0.296496f
C30 VTAIL.t5 B 2.76651f
C31 VTAIL.n1 B 0.368599f
C32 VTAIL.t7 B 2.76651f
C33 VTAIL.n2 B 1.54838f
C34 VTAIL.t1 B 2.76651f
C35 VTAIL.n3 B 1.54838f
C36 VTAIL.t2 B 2.76651f
C37 VTAIL.n4 B 0.368599f
C38 VTAIL.t4 B 2.76651f
C39 VTAIL.n5 B 0.368599f
C40 VTAIL.t6 B 2.76651f
C41 VTAIL.n6 B 1.54838f
C42 VTAIL.t0 B 2.76651f
C43 VTAIL.n7 B 1.47054f
C44 VDD1.t0 B 0.420116f
C45 VDD1.t1 B 0.420116f
C46 VDD1.n0 B 3.85256f
C47 VDD1.t3 B 0.420116f
C48 VDD1.t2 B 0.420116f
C49 VDD1.n1 B 4.85763f
C50 VP.t2 B 3.69563f
C51 VP.n0 B 1.35003f
C52 VP.n1 B 0.021061f
C53 VP.n2 B 0.01701f
C54 VP.n3 B 0.021061f
C55 VP.t0 B 3.69563f
C56 VP.n4 B 1.35003f
C57 VP.t3 B 3.96381f
C58 VP.t1 B 3.95558f
C59 VP.n5 B 3.95845f
C60 VP.n6 B 1.42798f
C61 VP.n7 B 0.033987f
C62 VP.n8 B 0.029994f
C63 VP.n9 B 0.039056f
C64 VP.n10 B 0.041638f
C65 VP.n11 B 0.021061f
C66 VP.n12 B 0.021061f
C67 VP.n13 B 0.021061f
C68 VP.n14 B 0.041638f
C69 VP.n15 B 0.039056f
C70 VP.n16 B 0.029994f
C71 VP.n17 B 0.033987f
C72 VP.n18 B 0.0514f
.ends

