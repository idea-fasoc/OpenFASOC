* NGSPICE file created from diff_pair_sample_1144.ext - technology: sky130A

.subckt diff_pair_sample_1144 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=0 ps=0 w=19.56 l=0.26
X1 B.t8 B.t6 B.t7 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=0 ps=0 w=19.56 l=0.26
X2 VDD2.t1 VN.t0 VTAIL.t2 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=7.6284 ps=39.9 w=19.56 l=0.26
X3 B.t5 B.t3 B.t4 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=0 ps=0 w=19.56 l=0.26
X4 VDD1.t1 VP.t0 VTAIL.t0 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=7.6284 ps=39.9 w=19.56 l=0.26
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=7.6284 ps=39.9 w=19.56 l=0.26
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=7.6284 ps=39.9 w=19.56 l=0.26
X7 B.t2 B.t0 B.t1 w_n1206_n4884# sky130_fd_pr__pfet_01v8 ad=7.6284 pd=39.9 as=0 ps=0 w=19.56 l=0.26
R0 B.n130 B.t3 2035.51
R1 B.n292 B.t0 2035.51
R2 B.n46 B.t9 2035.51
R3 B.n40 B.t6 2035.51
R4 B.n392 B.n391 585
R5 B.n390 B.n93 585
R6 B.n389 B.n388 585
R7 B.n387 B.n94 585
R8 B.n386 B.n385 585
R9 B.n384 B.n95 585
R10 B.n383 B.n382 585
R11 B.n381 B.n96 585
R12 B.n380 B.n379 585
R13 B.n378 B.n97 585
R14 B.n377 B.n376 585
R15 B.n375 B.n98 585
R16 B.n374 B.n373 585
R17 B.n372 B.n99 585
R18 B.n371 B.n370 585
R19 B.n369 B.n100 585
R20 B.n368 B.n367 585
R21 B.n366 B.n101 585
R22 B.n365 B.n364 585
R23 B.n363 B.n102 585
R24 B.n362 B.n361 585
R25 B.n360 B.n103 585
R26 B.n359 B.n358 585
R27 B.n357 B.n104 585
R28 B.n356 B.n355 585
R29 B.n354 B.n105 585
R30 B.n353 B.n352 585
R31 B.n351 B.n106 585
R32 B.n350 B.n349 585
R33 B.n348 B.n107 585
R34 B.n347 B.n346 585
R35 B.n345 B.n108 585
R36 B.n344 B.n343 585
R37 B.n342 B.n109 585
R38 B.n341 B.n340 585
R39 B.n339 B.n110 585
R40 B.n338 B.n337 585
R41 B.n336 B.n111 585
R42 B.n335 B.n334 585
R43 B.n333 B.n112 585
R44 B.n332 B.n331 585
R45 B.n330 B.n113 585
R46 B.n329 B.n328 585
R47 B.n327 B.n114 585
R48 B.n326 B.n325 585
R49 B.n324 B.n115 585
R50 B.n323 B.n322 585
R51 B.n321 B.n116 585
R52 B.n320 B.n319 585
R53 B.n318 B.n117 585
R54 B.n317 B.n316 585
R55 B.n315 B.n118 585
R56 B.n314 B.n313 585
R57 B.n312 B.n119 585
R58 B.n311 B.n310 585
R59 B.n309 B.n120 585
R60 B.n308 B.n307 585
R61 B.n306 B.n121 585
R62 B.n305 B.n304 585
R63 B.n303 B.n122 585
R64 B.n302 B.n301 585
R65 B.n300 B.n123 585
R66 B.n299 B.n298 585
R67 B.n297 B.n124 585
R68 B.n296 B.n295 585
R69 B.n291 B.n125 585
R70 B.n290 B.n289 585
R71 B.n288 B.n126 585
R72 B.n287 B.n286 585
R73 B.n285 B.n127 585
R74 B.n284 B.n283 585
R75 B.n282 B.n128 585
R76 B.n281 B.n280 585
R77 B.n278 B.n129 585
R78 B.n277 B.n276 585
R79 B.n275 B.n132 585
R80 B.n274 B.n273 585
R81 B.n272 B.n133 585
R82 B.n271 B.n270 585
R83 B.n269 B.n134 585
R84 B.n268 B.n267 585
R85 B.n266 B.n135 585
R86 B.n265 B.n264 585
R87 B.n263 B.n136 585
R88 B.n262 B.n261 585
R89 B.n260 B.n137 585
R90 B.n259 B.n258 585
R91 B.n257 B.n138 585
R92 B.n256 B.n255 585
R93 B.n254 B.n139 585
R94 B.n253 B.n252 585
R95 B.n251 B.n140 585
R96 B.n250 B.n249 585
R97 B.n248 B.n141 585
R98 B.n247 B.n246 585
R99 B.n245 B.n142 585
R100 B.n244 B.n243 585
R101 B.n242 B.n143 585
R102 B.n241 B.n240 585
R103 B.n239 B.n144 585
R104 B.n238 B.n237 585
R105 B.n236 B.n145 585
R106 B.n235 B.n234 585
R107 B.n233 B.n146 585
R108 B.n232 B.n231 585
R109 B.n230 B.n147 585
R110 B.n229 B.n228 585
R111 B.n227 B.n148 585
R112 B.n226 B.n225 585
R113 B.n224 B.n149 585
R114 B.n223 B.n222 585
R115 B.n221 B.n150 585
R116 B.n220 B.n219 585
R117 B.n218 B.n151 585
R118 B.n217 B.n216 585
R119 B.n215 B.n152 585
R120 B.n214 B.n213 585
R121 B.n212 B.n153 585
R122 B.n211 B.n210 585
R123 B.n209 B.n154 585
R124 B.n208 B.n207 585
R125 B.n206 B.n155 585
R126 B.n205 B.n204 585
R127 B.n203 B.n156 585
R128 B.n202 B.n201 585
R129 B.n200 B.n157 585
R130 B.n199 B.n198 585
R131 B.n197 B.n158 585
R132 B.n196 B.n195 585
R133 B.n194 B.n159 585
R134 B.n193 B.n192 585
R135 B.n191 B.n160 585
R136 B.n190 B.n189 585
R137 B.n188 B.n161 585
R138 B.n187 B.n186 585
R139 B.n185 B.n162 585
R140 B.n184 B.n183 585
R141 B.n393 B.n92 585
R142 B.n395 B.n394 585
R143 B.n396 B.n91 585
R144 B.n398 B.n397 585
R145 B.n399 B.n90 585
R146 B.n401 B.n400 585
R147 B.n402 B.n89 585
R148 B.n404 B.n403 585
R149 B.n405 B.n88 585
R150 B.n407 B.n406 585
R151 B.n408 B.n87 585
R152 B.n410 B.n409 585
R153 B.n411 B.n86 585
R154 B.n413 B.n412 585
R155 B.n414 B.n85 585
R156 B.n416 B.n415 585
R157 B.n417 B.n84 585
R158 B.n419 B.n418 585
R159 B.n420 B.n83 585
R160 B.n422 B.n421 585
R161 B.n423 B.n82 585
R162 B.n425 B.n424 585
R163 B.n426 B.n81 585
R164 B.n428 B.n427 585
R165 B.n635 B.n634 585
R166 B.n633 B.n8 585
R167 B.n632 B.n631 585
R168 B.n630 B.n9 585
R169 B.n629 B.n628 585
R170 B.n627 B.n10 585
R171 B.n626 B.n625 585
R172 B.n624 B.n11 585
R173 B.n623 B.n622 585
R174 B.n621 B.n12 585
R175 B.n620 B.n619 585
R176 B.n618 B.n13 585
R177 B.n617 B.n616 585
R178 B.n615 B.n14 585
R179 B.n614 B.n613 585
R180 B.n612 B.n15 585
R181 B.n611 B.n610 585
R182 B.n609 B.n16 585
R183 B.n608 B.n607 585
R184 B.n606 B.n17 585
R185 B.n605 B.n604 585
R186 B.n603 B.n18 585
R187 B.n602 B.n601 585
R188 B.n600 B.n19 585
R189 B.n599 B.n598 585
R190 B.n597 B.n20 585
R191 B.n596 B.n595 585
R192 B.n594 B.n21 585
R193 B.n593 B.n592 585
R194 B.n591 B.n22 585
R195 B.n590 B.n589 585
R196 B.n588 B.n23 585
R197 B.n587 B.n586 585
R198 B.n585 B.n24 585
R199 B.n584 B.n583 585
R200 B.n582 B.n25 585
R201 B.n581 B.n580 585
R202 B.n579 B.n26 585
R203 B.n578 B.n577 585
R204 B.n576 B.n27 585
R205 B.n575 B.n574 585
R206 B.n573 B.n28 585
R207 B.n572 B.n571 585
R208 B.n570 B.n29 585
R209 B.n569 B.n568 585
R210 B.n567 B.n30 585
R211 B.n566 B.n565 585
R212 B.n564 B.n31 585
R213 B.n563 B.n562 585
R214 B.n561 B.n32 585
R215 B.n560 B.n559 585
R216 B.n558 B.n33 585
R217 B.n557 B.n556 585
R218 B.n555 B.n34 585
R219 B.n554 B.n553 585
R220 B.n552 B.n35 585
R221 B.n551 B.n550 585
R222 B.n549 B.n36 585
R223 B.n548 B.n547 585
R224 B.n546 B.n37 585
R225 B.n545 B.n544 585
R226 B.n543 B.n38 585
R227 B.n542 B.n541 585
R228 B.n540 B.n39 585
R229 B.n538 B.n537 585
R230 B.n536 B.n42 585
R231 B.n535 B.n534 585
R232 B.n533 B.n43 585
R233 B.n532 B.n531 585
R234 B.n530 B.n44 585
R235 B.n529 B.n528 585
R236 B.n527 B.n45 585
R237 B.n526 B.n525 585
R238 B.n524 B.n523 585
R239 B.n522 B.n49 585
R240 B.n521 B.n520 585
R241 B.n519 B.n50 585
R242 B.n518 B.n517 585
R243 B.n516 B.n51 585
R244 B.n515 B.n514 585
R245 B.n513 B.n52 585
R246 B.n512 B.n511 585
R247 B.n510 B.n53 585
R248 B.n509 B.n508 585
R249 B.n507 B.n54 585
R250 B.n506 B.n505 585
R251 B.n504 B.n55 585
R252 B.n503 B.n502 585
R253 B.n501 B.n56 585
R254 B.n500 B.n499 585
R255 B.n498 B.n57 585
R256 B.n497 B.n496 585
R257 B.n495 B.n58 585
R258 B.n494 B.n493 585
R259 B.n492 B.n59 585
R260 B.n491 B.n490 585
R261 B.n489 B.n60 585
R262 B.n488 B.n487 585
R263 B.n486 B.n61 585
R264 B.n485 B.n484 585
R265 B.n483 B.n62 585
R266 B.n482 B.n481 585
R267 B.n480 B.n63 585
R268 B.n479 B.n478 585
R269 B.n477 B.n64 585
R270 B.n476 B.n475 585
R271 B.n474 B.n65 585
R272 B.n473 B.n472 585
R273 B.n471 B.n66 585
R274 B.n470 B.n469 585
R275 B.n468 B.n67 585
R276 B.n467 B.n466 585
R277 B.n465 B.n68 585
R278 B.n464 B.n463 585
R279 B.n462 B.n69 585
R280 B.n461 B.n460 585
R281 B.n459 B.n70 585
R282 B.n458 B.n457 585
R283 B.n456 B.n71 585
R284 B.n455 B.n454 585
R285 B.n453 B.n72 585
R286 B.n452 B.n451 585
R287 B.n450 B.n73 585
R288 B.n449 B.n448 585
R289 B.n447 B.n74 585
R290 B.n446 B.n445 585
R291 B.n444 B.n75 585
R292 B.n443 B.n442 585
R293 B.n441 B.n76 585
R294 B.n440 B.n439 585
R295 B.n438 B.n77 585
R296 B.n437 B.n436 585
R297 B.n435 B.n78 585
R298 B.n434 B.n433 585
R299 B.n432 B.n79 585
R300 B.n431 B.n430 585
R301 B.n429 B.n80 585
R302 B.n636 B.n7 585
R303 B.n638 B.n637 585
R304 B.n639 B.n6 585
R305 B.n641 B.n640 585
R306 B.n642 B.n5 585
R307 B.n644 B.n643 585
R308 B.n645 B.n4 585
R309 B.n647 B.n646 585
R310 B.n648 B.n3 585
R311 B.n650 B.n649 585
R312 B.n651 B.n0 585
R313 B.n2 B.n1 585
R314 B.n169 B.n168 585
R315 B.n170 B.n167 585
R316 B.n172 B.n171 585
R317 B.n173 B.n166 585
R318 B.n175 B.n174 585
R319 B.n176 B.n165 585
R320 B.n178 B.n177 585
R321 B.n179 B.n164 585
R322 B.n181 B.n180 585
R323 B.n182 B.n163 585
R324 B.n184 B.n163 545.355
R325 B.n393 B.n392 545.355
R326 B.n429 B.n428 545.355
R327 B.n634 B.n7 545.355
R328 B.n292 B.t1 523.253
R329 B.n46 B.t11 523.253
R330 B.n130 B.t4 523.253
R331 B.n40 B.t8 523.253
R332 B.n293 B.t2 511.81
R333 B.n47 B.t10 511.81
R334 B.n131 B.t5 511.81
R335 B.n41 B.t7 511.81
R336 B.n653 B.n652 256.663
R337 B.n652 B.n651 235.042
R338 B.n652 B.n2 235.042
R339 B.n185 B.n184 163.367
R340 B.n186 B.n185 163.367
R341 B.n186 B.n161 163.367
R342 B.n190 B.n161 163.367
R343 B.n191 B.n190 163.367
R344 B.n192 B.n191 163.367
R345 B.n192 B.n159 163.367
R346 B.n196 B.n159 163.367
R347 B.n197 B.n196 163.367
R348 B.n198 B.n197 163.367
R349 B.n198 B.n157 163.367
R350 B.n202 B.n157 163.367
R351 B.n203 B.n202 163.367
R352 B.n204 B.n203 163.367
R353 B.n204 B.n155 163.367
R354 B.n208 B.n155 163.367
R355 B.n209 B.n208 163.367
R356 B.n210 B.n209 163.367
R357 B.n210 B.n153 163.367
R358 B.n214 B.n153 163.367
R359 B.n215 B.n214 163.367
R360 B.n216 B.n215 163.367
R361 B.n216 B.n151 163.367
R362 B.n220 B.n151 163.367
R363 B.n221 B.n220 163.367
R364 B.n222 B.n221 163.367
R365 B.n222 B.n149 163.367
R366 B.n226 B.n149 163.367
R367 B.n227 B.n226 163.367
R368 B.n228 B.n227 163.367
R369 B.n228 B.n147 163.367
R370 B.n232 B.n147 163.367
R371 B.n233 B.n232 163.367
R372 B.n234 B.n233 163.367
R373 B.n234 B.n145 163.367
R374 B.n238 B.n145 163.367
R375 B.n239 B.n238 163.367
R376 B.n240 B.n239 163.367
R377 B.n240 B.n143 163.367
R378 B.n244 B.n143 163.367
R379 B.n245 B.n244 163.367
R380 B.n246 B.n245 163.367
R381 B.n246 B.n141 163.367
R382 B.n250 B.n141 163.367
R383 B.n251 B.n250 163.367
R384 B.n252 B.n251 163.367
R385 B.n252 B.n139 163.367
R386 B.n256 B.n139 163.367
R387 B.n257 B.n256 163.367
R388 B.n258 B.n257 163.367
R389 B.n258 B.n137 163.367
R390 B.n262 B.n137 163.367
R391 B.n263 B.n262 163.367
R392 B.n264 B.n263 163.367
R393 B.n264 B.n135 163.367
R394 B.n268 B.n135 163.367
R395 B.n269 B.n268 163.367
R396 B.n270 B.n269 163.367
R397 B.n270 B.n133 163.367
R398 B.n274 B.n133 163.367
R399 B.n275 B.n274 163.367
R400 B.n276 B.n275 163.367
R401 B.n276 B.n129 163.367
R402 B.n281 B.n129 163.367
R403 B.n282 B.n281 163.367
R404 B.n283 B.n282 163.367
R405 B.n283 B.n127 163.367
R406 B.n287 B.n127 163.367
R407 B.n288 B.n287 163.367
R408 B.n289 B.n288 163.367
R409 B.n289 B.n125 163.367
R410 B.n296 B.n125 163.367
R411 B.n297 B.n296 163.367
R412 B.n298 B.n297 163.367
R413 B.n298 B.n123 163.367
R414 B.n302 B.n123 163.367
R415 B.n303 B.n302 163.367
R416 B.n304 B.n303 163.367
R417 B.n304 B.n121 163.367
R418 B.n308 B.n121 163.367
R419 B.n309 B.n308 163.367
R420 B.n310 B.n309 163.367
R421 B.n310 B.n119 163.367
R422 B.n314 B.n119 163.367
R423 B.n315 B.n314 163.367
R424 B.n316 B.n315 163.367
R425 B.n316 B.n117 163.367
R426 B.n320 B.n117 163.367
R427 B.n321 B.n320 163.367
R428 B.n322 B.n321 163.367
R429 B.n322 B.n115 163.367
R430 B.n326 B.n115 163.367
R431 B.n327 B.n326 163.367
R432 B.n328 B.n327 163.367
R433 B.n328 B.n113 163.367
R434 B.n332 B.n113 163.367
R435 B.n333 B.n332 163.367
R436 B.n334 B.n333 163.367
R437 B.n334 B.n111 163.367
R438 B.n338 B.n111 163.367
R439 B.n339 B.n338 163.367
R440 B.n340 B.n339 163.367
R441 B.n340 B.n109 163.367
R442 B.n344 B.n109 163.367
R443 B.n345 B.n344 163.367
R444 B.n346 B.n345 163.367
R445 B.n346 B.n107 163.367
R446 B.n350 B.n107 163.367
R447 B.n351 B.n350 163.367
R448 B.n352 B.n351 163.367
R449 B.n352 B.n105 163.367
R450 B.n356 B.n105 163.367
R451 B.n357 B.n356 163.367
R452 B.n358 B.n357 163.367
R453 B.n358 B.n103 163.367
R454 B.n362 B.n103 163.367
R455 B.n363 B.n362 163.367
R456 B.n364 B.n363 163.367
R457 B.n364 B.n101 163.367
R458 B.n368 B.n101 163.367
R459 B.n369 B.n368 163.367
R460 B.n370 B.n369 163.367
R461 B.n370 B.n99 163.367
R462 B.n374 B.n99 163.367
R463 B.n375 B.n374 163.367
R464 B.n376 B.n375 163.367
R465 B.n376 B.n97 163.367
R466 B.n380 B.n97 163.367
R467 B.n381 B.n380 163.367
R468 B.n382 B.n381 163.367
R469 B.n382 B.n95 163.367
R470 B.n386 B.n95 163.367
R471 B.n387 B.n386 163.367
R472 B.n388 B.n387 163.367
R473 B.n388 B.n93 163.367
R474 B.n392 B.n93 163.367
R475 B.n428 B.n81 163.367
R476 B.n424 B.n81 163.367
R477 B.n424 B.n423 163.367
R478 B.n423 B.n422 163.367
R479 B.n422 B.n83 163.367
R480 B.n418 B.n83 163.367
R481 B.n418 B.n417 163.367
R482 B.n417 B.n416 163.367
R483 B.n416 B.n85 163.367
R484 B.n412 B.n85 163.367
R485 B.n412 B.n411 163.367
R486 B.n411 B.n410 163.367
R487 B.n410 B.n87 163.367
R488 B.n406 B.n87 163.367
R489 B.n406 B.n405 163.367
R490 B.n405 B.n404 163.367
R491 B.n404 B.n89 163.367
R492 B.n400 B.n89 163.367
R493 B.n400 B.n399 163.367
R494 B.n399 B.n398 163.367
R495 B.n398 B.n91 163.367
R496 B.n394 B.n91 163.367
R497 B.n394 B.n393 163.367
R498 B.n634 B.n633 163.367
R499 B.n633 B.n632 163.367
R500 B.n632 B.n9 163.367
R501 B.n628 B.n9 163.367
R502 B.n628 B.n627 163.367
R503 B.n627 B.n626 163.367
R504 B.n626 B.n11 163.367
R505 B.n622 B.n11 163.367
R506 B.n622 B.n621 163.367
R507 B.n621 B.n620 163.367
R508 B.n620 B.n13 163.367
R509 B.n616 B.n13 163.367
R510 B.n616 B.n615 163.367
R511 B.n615 B.n614 163.367
R512 B.n614 B.n15 163.367
R513 B.n610 B.n15 163.367
R514 B.n610 B.n609 163.367
R515 B.n609 B.n608 163.367
R516 B.n608 B.n17 163.367
R517 B.n604 B.n17 163.367
R518 B.n604 B.n603 163.367
R519 B.n603 B.n602 163.367
R520 B.n602 B.n19 163.367
R521 B.n598 B.n19 163.367
R522 B.n598 B.n597 163.367
R523 B.n597 B.n596 163.367
R524 B.n596 B.n21 163.367
R525 B.n592 B.n21 163.367
R526 B.n592 B.n591 163.367
R527 B.n591 B.n590 163.367
R528 B.n590 B.n23 163.367
R529 B.n586 B.n23 163.367
R530 B.n586 B.n585 163.367
R531 B.n585 B.n584 163.367
R532 B.n584 B.n25 163.367
R533 B.n580 B.n25 163.367
R534 B.n580 B.n579 163.367
R535 B.n579 B.n578 163.367
R536 B.n578 B.n27 163.367
R537 B.n574 B.n27 163.367
R538 B.n574 B.n573 163.367
R539 B.n573 B.n572 163.367
R540 B.n572 B.n29 163.367
R541 B.n568 B.n29 163.367
R542 B.n568 B.n567 163.367
R543 B.n567 B.n566 163.367
R544 B.n566 B.n31 163.367
R545 B.n562 B.n31 163.367
R546 B.n562 B.n561 163.367
R547 B.n561 B.n560 163.367
R548 B.n560 B.n33 163.367
R549 B.n556 B.n33 163.367
R550 B.n556 B.n555 163.367
R551 B.n555 B.n554 163.367
R552 B.n554 B.n35 163.367
R553 B.n550 B.n35 163.367
R554 B.n550 B.n549 163.367
R555 B.n549 B.n548 163.367
R556 B.n548 B.n37 163.367
R557 B.n544 B.n37 163.367
R558 B.n544 B.n543 163.367
R559 B.n543 B.n542 163.367
R560 B.n542 B.n39 163.367
R561 B.n537 B.n39 163.367
R562 B.n537 B.n536 163.367
R563 B.n536 B.n535 163.367
R564 B.n535 B.n43 163.367
R565 B.n531 B.n43 163.367
R566 B.n531 B.n530 163.367
R567 B.n530 B.n529 163.367
R568 B.n529 B.n45 163.367
R569 B.n525 B.n45 163.367
R570 B.n525 B.n524 163.367
R571 B.n524 B.n49 163.367
R572 B.n520 B.n49 163.367
R573 B.n520 B.n519 163.367
R574 B.n519 B.n518 163.367
R575 B.n518 B.n51 163.367
R576 B.n514 B.n51 163.367
R577 B.n514 B.n513 163.367
R578 B.n513 B.n512 163.367
R579 B.n512 B.n53 163.367
R580 B.n508 B.n53 163.367
R581 B.n508 B.n507 163.367
R582 B.n507 B.n506 163.367
R583 B.n506 B.n55 163.367
R584 B.n502 B.n55 163.367
R585 B.n502 B.n501 163.367
R586 B.n501 B.n500 163.367
R587 B.n500 B.n57 163.367
R588 B.n496 B.n57 163.367
R589 B.n496 B.n495 163.367
R590 B.n495 B.n494 163.367
R591 B.n494 B.n59 163.367
R592 B.n490 B.n59 163.367
R593 B.n490 B.n489 163.367
R594 B.n489 B.n488 163.367
R595 B.n488 B.n61 163.367
R596 B.n484 B.n61 163.367
R597 B.n484 B.n483 163.367
R598 B.n483 B.n482 163.367
R599 B.n482 B.n63 163.367
R600 B.n478 B.n63 163.367
R601 B.n478 B.n477 163.367
R602 B.n477 B.n476 163.367
R603 B.n476 B.n65 163.367
R604 B.n472 B.n65 163.367
R605 B.n472 B.n471 163.367
R606 B.n471 B.n470 163.367
R607 B.n470 B.n67 163.367
R608 B.n466 B.n67 163.367
R609 B.n466 B.n465 163.367
R610 B.n465 B.n464 163.367
R611 B.n464 B.n69 163.367
R612 B.n460 B.n69 163.367
R613 B.n460 B.n459 163.367
R614 B.n459 B.n458 163.367
R615 B.n458 B.n71 163.367
R616 B.n454 B.n71 163.367
R617 B.n454 B.n453 163.367
R618 B.n453 B.n452 163.367
R619 B.n452 B.n73 163.367
R620 B.n448 B.n73 163.367
R621 B.n448 B.n447 163.367
R622 B.n447 B.n446 163.367
R623 B.n446 B.n75 163.367
R624 B.n442 B.n75 163.367
R625 B.n442 B.n441 163.367
R626 B.n441 B.n440 163.367
R627 B.n440 B.n77 163.367
R628 B.n436 B.n77 163.367
R629 B.n436 B.n435 163.367
R630 B.n435 B.n434 163.367
R631 B.n434 B.n79 163.367
R632 B.n430 B.n79 163.367
R633 B.n430 B.n429 163.367
R634 B.n638 B.n7 163.367
R635 B.n639 B.n638 163.367
R636 B.n640 B.n639 163.367
R637 B.n640 B.n5 163.367
R638 B.n644 B.n5 163.367
R639 B.n645 B.n644 163.367
R640 B.n646 B.n645 163.367
R641 B.n646 B.n3 163.367
R642 B.n650 B.n3 163.367
R643 B.n651 B.n650 163.367
R644 B.n168 B.n2 163.367
R645 B.n168 B.n167 163.367
R646 B.n172 B.n167 163.367
R647 B.n173 B.n172 163.367
R648 B.n174 B.n173 163.367
R649 B.n174 B.n165 163.367
R650 B.n178 B.n165 163.367
R651 B.n179 B.n178 163.367
R652 B.n180 B.n179 163.367
R653 B.n180 B.n163 163.367
R654 B.n279 B.n131 59.5399
R655 B.n294 B.n293 59.5399
R656 B.n48 B.n47 59.5399
R657 B.n539 B.n41 59.5399
R658 B.n636 B.n635 35.4346
R659 B.n427 B.n80 35.4346
R660 B.n183 B.n182 35.4346
R661 B.n391 B.n92 35.4346
R662 B B.n653 18.0485
R663 B.n131 B.n130 11.4429
R664 B.n293 B.n292 11.4429
R665 B.n47 B.n46 11.4429
R666 B.n41 B.n40 11.4429
R667 B.n637 B.n636 10.6151
R668 B.n637 B.n6 10.6151
R669 B.n641 B.n6 10.6151
R670 B.n642 B.n641 10.6151
R671 B.n643 B.n642 10.6151
R672 B.n643 B.n4 10.6151
R673 B.n647 B.n4 10.6151
R674 B.n648 B.n647 10.6151
R675 B.n649 B.n648 10.6151
R676 B.n649 B.n0 10.6151
R677 B.n635 B.n8 10.6151
R678 B.n631 B.n8 10.6151
R679 B.n631 B.n630 10.6151
R680 B.n630 B.n629 10.6151
R681 B.n629 B.n10 10.6151
R682 B.n625 B.n10 10.6151
R683 B.n625 B.n624 10.6151
R684 B.n624 B.n623 10.6151
R685 B.n623 B.n12 10.6151
R686 B.n619 B.n12 10.6151
R687 B.n619 B.n618 10.6151
R688 B.n618 B.n617 10.6151
R689 B.n617 B.n14 10.6151
R690 B.n613 B.n14 10.6151
R691 B.n613 B.n612 10.6151
R692 B.n612 B.n611 10.6151
R693 B.n611 B.n16 10.6151
R694 B.n607 B.n16 10.6151
R695 B.n607 B.n606 10.6151
R696 B.n606 B.n605 10.6151
R697 B.n605 B.n18 10.6151
R698 B.n601 B.n18 10.6151
R699 B.n601 B.n600 10.6151
R700 B.n600 B.n599 10.6151
R701 B.n599 B.n20 10.6151
R702 B.n595 B.n20 10.6151
R703 B.n595 B.n594 10.6151
R704 B.n594 B.n593 10.6151
R705 B.n593 B.n22 10.6151
R706 B.n589 B.n22 10.6151
R707 B.n589 B.n588 10.6151
R708 B.n588 B.n587 10.6151
R709 B.n587 B.n24 10.6151
R710 B.n583 B.n24 10.6151
R711 B.n583 B.n582 10.6151
R712 B.n582 B.n581 10.6151
R713 B.n581 B.n26 10.6151
R714 B.n577 B.n26 10.6151
R715 B.n577 B.n576 10.6151
R716 B.n576 B.n575 10.6151
R717 B.n575 B.n28 10.6151
R718 B.n571 B.n28 10.6151
R719 B.n571 B.n570 10.6151
R720 B.n570 B.n569 10.6151
R721 B.n569 B.n30 10.6151
R722 B.n565 B.n30 10.6151
R723 B.n565 B.n564 10.6151
R724 B.n564 B.n563 10.6151
R725 B.n563 B.n32 10.6151
R726 B.n559 B.n32 10.6151
R727 B.n559 B.n558 10.6151
R728 B.n558 B.n557 10.6151
R729 B.n557 B.n34 10.6151
R730 B.n553 B.n34 10.6151
R731 B.n553 B.n552 10.6151
R732 B.n552 B.n551 10.6151
R733 B.n551 B.n36 10.6151
R734 B.n547 B.n36 10.6151
R735 B.n547 B.n546 10.6151
R736 B.n546 B.n545 10.6151
R737 B.n545 B.n38 10.6151
R738 B.n541 B.n38 10.6151
R739 B.n541 B.n540 10.6151
R740 B.n538 B.n42 10.6151
R741 B.n534 B.n42 10.6151
R742 B.n534 B.n533 10.6151
R743 B.n533 B.n532 10.6151
R744 B.n532 B.n44 10.6151
R745 B.n528 B.n44 10.6151
R746 B.n528 B.n527 10.6151
R747 B.n527 B.n526 10.6151
R748 B.n523 B.n522 10.6151
R749 B.n522 B.n521 10.6151
R750 B.n521 B.n50 10.6151
R751 B.n517 B.n50 10.6151
R752 B.n517 B.n516 10.6151
R753 B.n516 B.n515 10.6151
R754 B.n515 B.n52 10.6151
R755 B.n511 B.n52 10.6151
R756 B.n511 B.n510 10.6151
R757 B.n510 B.n509 10.6151
R758 B.n509 B.n54 10.6151
R759 B.n505 B.n54 10.6151
R760 B.n505 B.n504 10.6151
R761 B.n504 B.n503 10.6151
R762 B.n503 B.n56 10.6151
R763 B.n499 B.n56 10.6151
R764 B.n499 B.n498 10.6151
R765 B.n498 B.n497 10.6151
R766 B.n497 B.n58 10.6151
R767 B.n493 B.n58 10.6151
R768 B.n493 B.n492 10.6151
R769 B.n492 B.n491 10.6151
R770 B.n491 B.n60 10.6151
R771 B.n487 B.n60 10.6151
R772 B.n487 B.n486 10.6151
R773 B.n486 B.n485 10.6151
R774 B.n485 B.n62 10.6151
R775 B.n481 B.n62 10.6151
R776 B.n481 B.n480 10.6151
R777 B.n480 B.n479 10.6151
R778 B.n479 B.n64 10.6151
R779 B.n475 B.n64 10.6151
R780 B.n475 B.n474 10.6151
R781 B.n474 B.n473 10.6151
R782 B.n473 B.n66 10.6151
R783 B.n469 B.n66 10.6151
R784 B.n469 B.n468 10.6151
R785 B.n468 B.n467 10.6151
R786 B.n467 B.n68 10.6151
R787 B.n463 B.n68 10.6151
R788 B.n463 B.n462 10.6151
R789 B.n462 B.n461 10.6151
R790 B.n461 B.n70 10.6151
R791 B.n457 B.n70 10.6151
R792 B.n457 B.n456 10.6151
R793 B.n456 B.n455 10.6151
R794 B.n455 B.n72 10.6151
R795 B.n451 B.n72 10.6151
R796 B.n451 B.n450 10.6151
R797 B.n450 B.n449 10.6151
R798 B.n449 B.n74 10.6151
R799 B.n445 B.n74 10.6151
R800 B.n445 B.n444 10.6151
R801 B.n444 B.n443 10.6151
R802 B.n443 B.n76 10.6151
R803 B.n439 B.n76 10.6151
R804 B.n439 B.n438 10.6151
R805 B.n438 B.n437 10.6151
R806 B.n437 B.n78 10.6151
R807 B.n433 B.n78 10.6151
R808 B.n433 B.n432 10.6151
R809 B.n432 B.n431 10.6151
R810 B.n431 B.n80 10.6151
R811 B.n427 B.n426 10.6151
R812 B.n426 B.n425 10.6151
R813 B.n425 B.n82 10.6151
R814 B.n421 B.n82 10.6151
R815 B.n421 B.n420 10.6151
R816 B.n420 B.n419 10.6151
R817 B.n419 B.n84 10.6151
R818 B.n415 B.n84 10.6151
R819 B.n415 B.n414 10.6151
R820 B.n414 B.n413 10.6151
R821 B.n413 B.n86 10.6151
R822 B.n409 B.n86 10.6151
R823 B.n409 B.n408 10.6151
R824 B.n408 B.n407 10.6151
R825 B.n407 B.n88 10.6151
R826 B.n403 B.n88 10.6151
R827 B.n403 B.n402 10.6151
R828 B.n402 B.n401 10.6151
R829 B.n401 B.n90 10.6151
R830 B.n397 B.n90 10.6151
R831 B.n397 B.n396 10.6151
R832 B.n396 B.n395 10.6151
R833 B.n395 B.n92 10.6151
R834 B.n169 B.n1 10.6151
R835 B.n170 B.n169 10.6151
R836 B.n171 B.n170 10.6151
R837 B.n171 B.n166 10.6151
R838 B.n175 B.n166 10.6151
R839 B.n176 B.n175 10.6151
R840 B.n177 B.n176 10.6151
R841 B.n177 B.n164 10.6151
R842 B.n181 B.n164 10.6151
R843 B.n182 B.n181 10.6151
R844 B.n183 B.n162 10.6151
R845 B.n187 B.n162 10.6151
R846 B.n188 B.n187 10.6151
R847 B.n189 B.n188 10.6151
R848 B.n189 B.n160 10.6151
R849 B.n193 B.n160 10.6151
R850 B.n194 B.n193 10.6151
R851 B.n195 B.n194 10.6151
R852 B.n195 B.n158 10.6151
R853 B.n199 B.n158 10.6151
R854 B.n200 B.n199 10.6151
R855 B.n201 B.n200 10.6151
R856 B.n201 B.n156 10.6151
R857 B.n205 B.n156 10.6151
R858 B.n206 B.n205 10.6151
R859 B.n207 B.n206 10.6151
R860 B.n207 B.n154 10.6151
R861 B.n211 B.n154 10.6151
R862 B.n212 B.n211 10.6151
R863 B.n213 B.n212 10.6151
R864 B.n213 B.n152 10.6151
R865 B.n217 B.n152 10.6151
R866 B.n218 B.n217 10.6151
R867 B.n219 B.n218 10.6151
R868 B.n219 B.n150 10.6151
R869 B.n223 B.n150 10.6151
R870 B.n224 B.n223 10.6151
R871 B.n225 B.n224 10.6151
R872 B.n225 B.n148 10.6151
R873 B.n229 B.n148 10.6151
R874 B.n230 B.n229 10.6151
R875 B.n231 B.n230 10.6151
R876 B.n231 B.n146 10.6151
R877 B.n235 B.n146 10.6151
R878 B.n236 B.n235 10.6151
R879 B.n237 B.n236 10.6151
R880 B.n237 B.n144 10.6151
R881 B.n241 B.n144 10.6151
R882 B.n242 B.n241 10.6151
R883 B.n243 B.n242 10.6151
R884 B.n243 B.n142 10.6151
R885 B.n247 B.n142 10.6151
R886 B.n248 B.n247 10.6151
R887 B.n249 B.n248 10.6151
R888 B.n249 B.n140 10.6151
R889 B.n253 B.n140 10.6151
R890 B.n254 B.n253 10.6151
R891 B.n255 B.n254 10.6151
R892 B.n255 B.n138 10.6151
R893 B.n259 B.n138 10.6151
R894 B.n260 B.n259 10.6151
R895 B.n261 B.n260 10.6151
R896 B.n261 B.n136 10.6151
R897 B.n265 B.n136 10.6151
R898 B.n266 B.n265 10.6151
R899 B.n267 B.n266 10.6151
R900 B.n267 B.n134 10.6151
R901 B.n271 B.n134 10.6151
R902 B.n272 B.n271 10.6151
R903 B.n273 B.n272 10.6151
R904 B.n273 B.n132 10.6151
R905 B.n277 B.n132 10.6151
R906 B.n278 B.n277 10.6151
R907 B.n280 B.n128 10.6151
R908 B.n284 B.n128 10.6151
R909 B.n285 B.n284 10.6151
R910 B.n286 B.n285 10.6151
R911 B.n286 B.n126 10.6151
R912 B.n290 B.n126 10.6151
R913 B.n291 B.n290 10.6151
R914 B.n295 B.n291 10.6151
R915 B.n299 B.n124 10.6151
R916 B.n300 B.n299 10.6151
R917 B.n301 B.n300 10.6151
R918 B.n301 B.n122 10.6151
R919 B.n305 B.n122 10.6151
R920 B.n306 B.n305 10.6151
R921 B.n307 B.n306 10.6151
R922 B.n307 B.n120 10.6151
R923 B.n311 B.n120 10.6151
R924 B.n312 B.n311 10.6151
R925 B.n313 B.n312 10.6151
R926 B.n313 B.n118 10.6151
R927 B.n317 B.n118 10.6151
R928 B.n318 B.n317 10.6151
R929 B.n319 B.n318 10.6151
R930 B.n319 B.n116 10.6151
R931 B.n323 B.n116 10.6151
R932 B.n324 B.n323 10.6151
R933 B.n325 B.n324 10.6151
R934 B.n325 B.n114 10.6151
R935 B.n329 B.n114 10.6151
R936 B.n330 B.n329 10.6151
R937 B.n331 B.n330 10.6151
R938 B.n331 B.n112 10.6151
R939 B.n335 B.n112 10.6151
R940 B.n336 B.n335 10.6151
R941 B.n337 B.n336 10.6151
R942 B.n337 B.n110 10.6151
R943 B.n341 B.n110 10.6151
R944 B.n342 B.n341 10.6151
R945 B.n343 B.n342 10.6151
R946 B.n343 B.n108 10.6151
R947 B.n347 B.n108 10.6151
R948 B.n348 B.n347 10.6151
R949 B.n349 B.n348 10.6151
R950 B.n349 B.n106 10.6151
R951 B.n353 B.n106 10.6151
R952 B.n354 B.n353 10.6151
R953 B.n355 B.n354 10.6151
R954 B.n355 B.n104 10.6151
R955 B.n359 B.n104 10.6151
R956 B.n360 B.n359 10.6151
R957 B.n361 B.n360 10.6151
R958 B.n361 B.n102 10.6151
R959 B.n365 B.n102 10.6151
R960 B.n366 B.n365 10.6151
R961 B.n367 B.n366 10.6151
R962 B.n367 B.n100 10.6151
R963 B.n371 B.n100 10.6151
R964 B.n372 B.n371 10.6151
R965 B.n373 B.n372 10.6151
R966 B.n373 B.n98 10.6151
R967 B.n377 B.n98 10.6151
R968 B.n378 B.n377 10.6151
R969 B.n379 B.n378 10.6151
R970 B.n379 B.n96 10.6151
R971 B.n383 B.n96 10.6151
R972 B.n384 B.n383 10.6151
R973 B.n385 B.n384 10.6151
R974 B.n385 B.n94 10.6151
R975 B.n389 B.n94 10.6151
R976 B.n390 B.n389 10.6151
R977 B.n391 B.n390 10.6151
R978 B.n653 B.n0 8.11757
R979 B.n653 B.n1 8.11757
R980 B.n539 B.n538 7.18099
R981 B.n526 B.n48 7.18099
R982 B.n280 B.n279 7.18099
R983 B.n295 B.n294 7.18099
R984 B.n540 B.n539 3.43465
R985 B.n523 B.n48 3.43465
R986 B.n279 B.n278 3.43465
R987 B.n294 B.n124 3.43465
R988 VN VN.t1 2163.54
R989 VN VN.t0 2119.01
R990 VTAIL.n353 VTAIL.n352 585
R991 VTAIL.n350 VTAIL.n349 585
R992 VTAIL.n359 VTAIL.n358 585
R993 VTAIL.n361 VTAIL.n360 585
R994 VTAIL.n346 VTAIL.n345 585
R995 VTAIL.n367 VTAIL.n366 585
R996 VTAIL.n370 VTAIL.n369 585
R997 VTAIL.n368 VTAIL.n342 585
R998 VTAIL.n375 VTAIL.n341 585
R999 VTAIL.n377 VTAIL.n376 585
R1000 VTAIL.n379 VTAIL.n378 585
R1001 VTAIL.n338 VTAIL.n337 585
R1002 VTAIL.n385 VTAIL.n384 585
R1003 VTAIL.n387 VTAIL.n386 585
R1004 VTAIL.n334 VTAIL.n333 585
R1005 VTAIL.n393 VTAIL.n392 585
R1006 VTAIL.n395 VTAIL.n394 585
R1007 VTAIL.n330 VTAIL.n329 585
R1008 VTAIL.n401 VTAIL.n400 585
R1009 VTAIL.n403 VTAIL.n402 585
R1010 VTAIL.n326 VTAIL.n325 585
R1011 VTAIL.n409 VTAIL.n408 585
R1012 VTAIL.n411 VTAIL.n410 585
R1013 VTAIL.n322 VTAIL.n321 585
R1014 VTAIL.n417 VTAIL.n416 585
R1015 VTAIL.n419 VTAIL.n418 585
R1016 VTAIL.n35 VTAIL.n34 585
R1017 VTAIL.n32 VTAIL.n31 585
R1018 VTAIL.n41 VTAIL.n40 585
R1019 VTAIL.n43 VTAIL.n42 585
R1020 VTAIL.n28 VTAIL.n27 585
R1021 VTAIL.n49 VTAIL.n48 585
R1022 VTAIL.n52 VTAIL.n51 585
R1023 VTAIL.n50 VTAIL.n24 585
R1024 VTAIL.n57 VTAIL.n23 585
R1025 VTAIL.n59 VTAIL.n58 585
R1026 VTAIL.n61 VTAIL.n60 585
R1027 VTAIL.n20 VTAIL.n19 585
R1028 VTAIL.n67 VTAIL.n66 585
R1029 VTAIL.n69 VTAIL.n68 585
R1030 VTAIL.n16 VTAIL.n15 585
R1031 VTAIL.n75 VTAIL.n74 585
R1032 VTAIL.n77 VTAIL.n76 585
R1033 VTAIL.n12 VTAIL.n11 585
R1034 VTAIL.n83 VTAIL.n82 585
R1035 VTAIL.n85 VTAIL.n84 585
R1036 VTAIL.n8 VTAIL.n7 585
R1037 VTAIL.n91 VTAIL.n90 585
R1038 VTAIL.n93 VTAIL.n92 585
R1039 VTAIL.n4 VTAIL.n3 585
R1040 VTAIL.n99 VTAIL.n98 585
R1041 VTAIL.n101 VTAIL.n100 585
R1042 VTAIL.n313 VTAIL.n312 585
R1043 VTAIL.n311 VTAIL.n310 585
R1044 VTAIL.n216 VTAIL.n215 585
R1045 VTAIL.n305 VTAIL.n304 585
R1046 VTAIL.n303 VTAIL.n302 585
R1047 VTAIL.n220 VTAIL.n219 585
R1048 VTAIL.n297 VTAIL.n296 585
R1049 VTAIL.n295 VTAIL.n294 585
R1050 VTAIL.n224 VTAIL.n223 585
R1051 VTAIL.n289 VTAIL.n288 585
R1052 VTAIL.n287 VTAIL.n286 585
R1053 VTAIL.n228 VTAIL.n227 585
R1054 VTAIL.n281 VTAIL.n280 585
R1055 VTAIL.n279 VTAIL.n278 585
R1056 VTAIL.n232 VTAIL.n231 585
R1057 VTAIL.n273 VTAIL.n272 585
R1058 VTAIL.n271 VTAIL.n270 585
R1059 VTAIL.n269 VTAIL.n235 585
R1060 VTAIL.n239 VTAIL.n236 585
R1061 VTAIL.n264 VTAIL.n263 585
R1062 VTAIL.n262 VTAIL.n261 585
R1063 VTAIL.n241 VTAIL.n240 585
R1064 VTAIL.n256 VTAIL.n255 585
R1065 VTAIL.n254 VTAIL.n253 585
R1066 VTAIL.n245 VTAIL.n244 585
R1067 VTAIL.n248 VTAIL.n247 585
R1068 VTAIL.n207 VTAIL.n206 585
R1069 VTAIL.n205 VTAIL.n204 585
R1070 VTAIL.n110 VTAIL.n109 585
R1071 VTAIL.n199 VTAIL.n198 585
R1072 VTAIL.n197 VTAIL.n196 585
R1073 VTAIL.n114 VTAIL.n113 585
R1074 VTAIL.n191 VTAIL.n190 585
R1075 VTAIL.n189 VTAIL.n188 585
R1076 VTAIL.n118 VTAIL.n117 585
R1077 VTAIL.n183 VTAIL.n182 585
R1078 VTAIL.n181 VTAIL.n180 585
R1079 VTAIL.n122 VTAIL.n121 585
R1080 VTAIL.n175 VTAIL.n174 585
R1081 VTAIL.n173 VTAIL.n172 585
R1082 VTAIL.n126 VTAIL.n125 585
R1083 VTAIL.n167 VTAIL.n166 585
R1084 VTAIL.n165 VTAIL.n164 585
R1085 VTAIL.n163 VTAIL.n129 585
R1086 VTAIL.n133 VTAIL.n130 585
R1087 VTAIL.n158 VTAIL.n157 585
R1088 VTAIL.n156 VTAIL.n155 585
R1089 VTAIL.n135 VTAIL.n134 585
R1090 VTAIL.n150 VTAIL.n149 585
R1091 VTAIL.n148 VTAIL.n147 585
R1092 VTAIL.n139 VTAIL.n138 585
R1093 VTAIL.n142 VTAIL.n141 585
R1094 VTAIL.n418 VTAIL.n318 498.474
R1095 VTAIL.n100 VTAIL.n0 498.474
R1096 VTAIL.n312 VTAIL.n212 498.474
R1097 VTAIL.n206 VTAIL.n106 498.474
R1098 VTAIL.t2 VTAIL.n351 329.036
R1099 VTAIL.t1 VTAIL.n33 329.036
R1100 VTAIL.t0 VTAIL.n246 329.036
R1101 VTAIL.t3 VTAIL.n140 329.036
R1102 VTAIL.n352 VTAIL.n349 171.744
R1103 VTAIL.n359 VTAIL.n349 171.744
R1104 VTAIL.n360 VTAIL.n359 171.744
R1105 VTAIL.n360 VTAIL.n345 171.744
R1106 VTAIL.n367 VTAIL.n345 171.744
R1107 VTAIL.n369 VTAIL.n367 171.744
R1108 VTAIL.n369 VTAIL.n368 171.744
R1109 VTAIL.n368 VTAIL.n341 171.744
R1110 VTAIL.n377 VTAIL.n341 171.744
R1111 VTAIL.n378 VTAIL.n377 171.744
R1112 VTAIL.n378 VTAIL.n337 171.744
R1113 VTAIL.n385 VTAIL.n337 171.744
R1114 VTAIL.n386 VTAIL.n385 171.744
R1115 VTAIL.n386 VTAIL.n333 171.744
R1116 VTAIL.n393 VTAIL.n333 171.744
R1117 VTAIL.n394 VTAIL.n393 171.744
R1118 VTAIL.n394 VTAIL.n329 171.744
R1119 VTAIL.n401 VTAIL.n329 171.744
R1120 VTAIL.n402 VTAIL.n401 171.744
R1121 VTAIL.n402 VTAIL.n325 171.744
R1122 VTAIL.n409 VTAIL.n325 171.744
R1123 VTAIL.n410 VTAIL.n409 171.744
R1124 VTAIL.n410 VTAIL.n321 171.744
R1125 VTAIL.n417 VTAIL.n321 171.744
R1126 VTAIL.n418 VTAIL.n417 171.744
R1127 VTAIL.n34 VTAIL.n31 171.744
R1128 VTAIL.n41 VTAIL.n31 171.744
R1129 VTAIL.n42 VTAIL.n41 171.744
R1130 VTAIL.n42 VTAIL.n27 171.744
R1131 VTAIL.n49 VTAIL.n27 171.744
R1132 VTAIL.n51 VTAIL.n49 171.744
R1133 VTAIL.n51 VTAIL.n50 171.744
R1134 VTAIL.n50 VTAIL.n23 171.744
R1135 VTAIL.n59 VTAIL.n23 171.744
R1136 VTAIL.n60 VTAIL.n59 171.744
R1137 VTAIL.n60 VTAIL.n19 171.744
R1138 VTAIL.n67 VTAIL.n19 171.744
R1139 VTAIL.n68 VTAIL.n67 171.744
R1140 VTAIL.n68 VTAIL.n15 171.744
R1141 VTAIL.n75 VTAIL.n15 171.744
R1142 VTAIL.n76 VTAIL.n75 171.744
R1143 VTAIL.n76 VTAIL.n11 171.744
R1144 VTAIL.n83 VTAIL.n11 171.744
R1145 VTAIL.n84 VTAIL.n83 171.744
R1146 VTAIL.n84 VTAIL.n7 171.744
R1147 VTAIL.n91 VTAIL.n7 171.744
R1148 VTAIL.n92 VTAIL.n91 171.744
R1149 VTAIL.n92 VTAIL.n3 171.744
R1150 VTAIL.n99 VTAIL.n3 171.744
R1151 VTAIL.n100 VTAIL.n99 171.744
R1152 VTAIL.n312 VTAIL.n311 171.744
R1153 VTAIL.n311 VTAIL.n215 171.744
R1154 VTAIL.n304 VTAIL.n215 171.744
R1155 VTAIL.n304 VTAIL.n303 171.744
R1156 VTAIL.n303 VTAIL.n219 171.744
R1157 VTAIL.n296 VTAIL.n219 171.744
R1158 VTAIL.n296 VTAIL.n295 171.744
R1159 VTAIL.n295 VTAIL.n223 171.744
R1160 VTAIL.n288 VTAIL.n223 171.744
R1161 VTAIL.n288 VTAIL.n287 171.744
R1162 VTAIL.n287 VTAIL.n227 171.744
R1163 VTAIL.n280 VTAIL.n227 171.744
R1164 VTAIL.n280 VTAIL.n279 171.744
R1165 VTAIL.n279 VTAIL.n231 171.744
R1166 VTAIL.n272 VTAIL.n231 171.744
R1167 VTAIL.n272 VTAIL.n271 171.744
R1168 VTAIL.n271 VTAIL.n235 171.744
R1169 VTAIL.n239 VTAIL.n235 171.744
R1170 VTAIL.n263 VTAIL.n239 171.744
R1171 VTAIL.n263 VTAIL.n262 171.744
R1172 VTAIL.n262 VTAIL.n240 171.744
R1173 VTAIL.n255 VTAIL.n240 171.744
R1174 VTAIL.n255 VTAIL.n254 171.744
R1175 VTAIL.n254 VTAIL.n244 171.744
R1176 VTAIL.n247 VTAIL.n244 171.744
R1177 VTAIL.n206 VTAIL.n205 171.744
R1178 VTAIL.n205 VTAIL.n109 171.744
R1179 VTAIL.n198 VTAIL.n109 171.744
R1180 VTAIL.n198 VTAIL.n197 171.744
R1181 VTAIL.n197 VTAIL.n113 171.744
R1182 VTAIL.n190 VTAIL.n113 171.744
R1183 VTAIL.n190 VTAIL.n189 171.744
R1184 VTAIL.n189 VTAIL.n117 171.744
R1185 VTAIL.n182 VTAIL.n117 171.744
R1186 VTAIL.n182 VTAIL.n181 171.744
R1187 VTAIL.n181 VTAIL.n121 171.744
R1188 VTAIL.n174 VTAIL.n121 171.744
R1189 VTAIL.n174 VTAIL.n173 171.744
R1190 VTAIL.n173 VTAIL.n125 171.744
R1191 VTAIL.n166 VTAIL.n125 171.744
R1192 VTAIL.n166 VTAIL.n165 171.744
R1193 VTAIL.n165 VTAIL.n129 171.744
R1194 VTAIL.n133 VTAIL.n129 171.744
R1195 VTAIL.n157 VTAIL.n133 171.744
R1196 VTAIL.n157 VTAIL.n156 171.744
R1197 VTAIL.n156 VTAIL.n134 171.744
R1198 VTAIL.n149 VTAIL.n134 171.744
R1199 VTAIL.n149 VTAIL.n148 171.744
R1200 VTAIL.n148 VTAIL.n138 171.744
R1201 VTAIL.n141 VTAIL.n138 171.744
R1202 VTAIL.n352 VTAIL.t2 85.8723
R1203 VTAIL.n34 VTAIL.t1 85.8723
R1204 VTAIL.n247 VTAIL.t0 85.8723
R1205 VTAIL.n141 VTAIL.t3 85.8723
R1206 VTAIL.n423 VTAIL.n422 36.8399
R1207 VTAIL.n105 VTAIL.n104 36.8399
R1208 VTAIL.n317 VTAIL.n316 36.8399
R1209 VTAIL.n211 VTAIL.n210 36.8399
R1210 VTAIL.n211 VTAIL.n105 30.2634
R1211 VTAIL.n423 VTAIL.n317 29.7548
R1212 VTAIL.n376 VTAIL.n375 13.1884
R1213 VTAIL.n58 VTAIL.n57 13.1884
R1214 VTAIL.n270 VTAIL.n269 13.1884
R1215 VTAIL.n164 VTAIL.n163 13.1884
R1216 VTAIL.n374 VTAIL.n342 12.8005
R1217 VTAIL.n379 VTAIL.n340 12.8005
R1218 VTAIL.n420 VTAIL.n419 12.8005
R1219 VTAIL.n56 VTAIL.n24 12.8005
R1220 VTAIL.n61 VTAIL.n22 12.8005
R1221 VTAIL.n102 VTAIL.n101 12.8005
R1222 VTAIL.n314 VTAIL.n313 12.8005
R1223 VTAIL.n273 VTAIL.n234 12.8005
R1224 VTAIL.n268 VTAIL.n236 12.8005
R1225 VTAIL.n208 VTAIL.n207 12.8005
R1226 VTAIL.n167 VTAIL.n128 12.8005
R1227 VTAIL.n162 VTAIL.n130 12.8005
R1228 VTAIL.n371 VTAIL.n370 12.0247
R1229 VTAIL.n380 VTAIL.n338 12.0247
R1230 VTAIL.n416 VTAIL.n320 12.0247
R1231 VTAIL.n53 VTAIL.n52 12.0247
R1232 VTAIL.n62 VTAIL.n20 12.0247
R1233 VTAIL.n98 VTAIL.n2 12.0247
R1234 VTAIL.n310 VTAIL.n214 12.0247
R1235 VTAIL.n274 VTAIL.n232 12.0247
R1236 VTAIL.n265 VTAIL.n264 12.0247
R1237 VTAIL.n204 VTAIL.n108 12.0247
R1238 VTAIL.n168 VTAIL.n126 12.0247
R1239 VTAIL.n159 VTAIL.n158 12.0247
R1240 VTAIL.n366 VTAIL.n344 11.249
R1241 VTAIL.n384 VTAIL.n383 11.249
R1242 VTAIL.n415 VTAIL.n322 11.249
R1243 VTAIL.n48 VTAIL.n26 11.249
R1244 VTAIL.n66 VTAIL.n65 11.249
R1245 VTAIL.n97 VTAIL.n4 11.249
R1246 VTAIL.n309 VTAIL.n216 11.249
R1247 VTAIL.n278 VTAIL.n277 11.249
R1248 VTAIL.n261 VTAIL.n238 11.249
R1249 VTAIL.n203 VTAIL.n110 11.249
R1250 VTAIL.n172 VTAIL.n171 11.249
R1251 VTAIL.n155 VTAIL.n132 11.249
R1252 VTAIL.n353 VTAIL.n351 10.7239
R1253 VTAIL.n35 VTAIL.n33 10.7239
R1254 VTAIL.n248 VTAIL.n246 10.7239
R1255 VTAIL.n142 VTAIL.n140 10.7239
R1256 VTAIL.n365 VTAIL.n346 10.4732
R1257 VTAIL.n387 VTAIL.n336 10.4732
R1258 VTAIL.n412 VTAIL.n411 10.4732
R1259 VTAIL.n47 VTAIL.n28 10.4732
R1260 VTAIL.n69 VTAIL.n18 10.4732
R1261 VTAIL.n94 VTAIL.n93 10.4732
R1262 VTAIL.n306 VTAIL.n305 10.4732
R1263 VTAIL.n281 VTAIL.n230 10.4732
R1264 VTAIL.n260 VTAIL.n241 10.4732
R1265 VTAIL.n200 VTAIL.n199 10.4732
R1266 VTAIL.n175 VTAIL.n124 10.4732
R1267 VTAIL.n154 VTAIL.n135 10.4732
R1268 VTAIL.n362 VTAIL.n361 9.69747
R1269 VTAIL.n388 VTAIL.n334 9.69747
R1270 VTAIL.n408 VTAIL.n324 9.69747
R1271 VTAIL.n44 VTAIL.n43 9.69747
R1272 VTAIL.n70 VTAIL.n16 9.69747
R1273 VTAIL.n90 VTAIL.n6 9.69747
R1274 VTAIL.n302 VTAIL.n218 9.69747
R1275 VTAIL.n282 VTAIL.n228 9.69747
R1276 VTAIL.n257 VTAIL.n256 9.69747
R1277 VTAIL.n196 VTAIL.n112 9.69747
R1278 VTAIL.n176 VTAIL.n122 9.69747
R1279 VTAIL.n151 VTAIL.n150 9.69747
R1280 VTAIL.n422 VTAIL.n421 9.45567
R1281 VTAIL.n104 VTAIL.n103 9.45567
R1282 VTAIL.n316 VTAIL.n315 9.45567
R1283 VTAIL.n210 VTAIL.n209 9.45567
R1284 VTAIL.n397 VTAIL.n396 9.3005
R1285 VTAIL.n332 VTAIL.n331 9.3005
R1286 VTAIL.n391 VTAIL.n390 9.3005
R1287 VTAIL.n389 VTAIL.n388 9.3005
R1288 VTAIL.n336 VTAIL.n335 9.3005
R1289 VTAIL.n383 VTAIL.n382 9.3005
R1290 VTAIL.n381 VTAIL.n380 9.3005
R1291 VTAIL.n340 VTAIL.n339 9.3005
R1292 VTAIL.n355 VTAIL.n354 9.3005
R1293 VTAIL.n357 VTAIL.n356 9.3005
R1294 VTAIL.n348 VTAIL.n347 9.3005
R1295 VTAIL.n363 VTAIL.n362 9.3005
R1296 VTAIL.n365 VTAIL.n364 9.3005
R1297 VTAIL.n344 VTAIL.n343 9.3005
R1298 VTAIL.n372 VTAIL.n371 9.3005
R1299 VTAIL.n374 VTAIL.n373 9.3005
R1300 VTAIL.n399 VTAIL.n398 9.3005
R1301 VTAIL.n328 VTAIL.n327 9.3005
R1302 VTAIL.n405 VTAIL.n404 9.3005
R1303 VTAIL.n407 VTAIL.n406 9.3005
R1304 VTAIL.n324 VTAIL.n323 9.3005
R1305 VTAIL.n413 VTAIL.n412 9.3005
R1306 VTAIL.n415 VTAIL.n414 9.3005
R1307 VTAIL.n320 VTAIL.n319 9.3005
R1308 VTAIL.n421 VTAIL.n420 9.3005
R1309 VTAIL.n79 VTAIL.n78 9.3005
R1310 VTAIL.n14 VTAIL.n13 9.3005
R1311 VTAIL.n73 VTAIL.n72 9.3005
R1312 VTAIL.n71 VTAIL.n70 9.3005
R1313 VTAIL.n18 VTAIL.n17 9.3005
R1314 VTAIL.n65 VTAIL.n64 9.3005
R1315 VTAIL.n63 VTAIL.n62 9.3005
R1316 VTAIL.n22 VTAIL.n21 9.3005
R1317 VTAIL.n37 VTAIL.n36 9.3005
R1318 VTAIL.n39 VTAIL.n38 9.3005
R1319 VTAIL.n30 VTAIL.n29 9.3005
R1320 VTAIL.n45 VTAIL.n44 9.3005
R1321 VTAIL.n47 VTAIL.n46 9.3005
R1322 VTAIL.n26 VTAIL.n25 9.3005
R1323 VTAIL.n54 VTAIL.n53 9.3005
R1324 VTAIL.n56 VTAIL.n55 9.3005
R1325 VTAIL.n81 VTAIL.n80 9.3005
R1326 VTAIL.n10 VTAIL.n9 9.3005
R1327 VTAIL.n87 VTAIL.n86 9.3005
R1328 VTAIL.n89 VTAIL.n88 9.3005
R1329 VTAIL.n6 VTAIL.n5 9.3005
R1330 VTAIL.n95 VTAIL.n94 9.3005
R1331 VTAIL.n97 VTAIL.n96 9.3005
R1332 VTAIL.n2 VTAIL.n1 9.3005
R1333 VTAIL.n103 VTAIL.n102 9.3005
R1334 VTAIL.n250 VTAIL.n249 9.3005
R1335 VTAIL.n252 VTAIL.n251 9.3005
R1336 VTAIL.n243 VTAIL.n242 9.3005
R1337 VTAIL.n258 VTAIL.n257 9.3005
R1338 VTAIL.n260 VTAIL.n259 9.3005
R1339 VTAIL.n238 VTAIL.n237 9.3005
R1340 VTAIL.n266 VTAIL.n265 9.3005
R1341 VTAIL.n268 VTAIL.n267 9.3005
R1342 VTAIL.n222 VTAIL.n221 9.3005
R1343 VTAIL.n299 VTAIL.n298 9.3005
R1344 VTAIL.n301 VTAIL.n300 9.3005
R1345 VTAIL.n218 VTAIL.n217 9.3005
R1346 VTAIL.n307 VTAIL.n306 9.3005
R1347 VTAIL.n309 VTAIL.n308 9.3005
R1348 VTAIL.n214 VTAIL.n213 9.3005
R1349 VTAIL.n315 VTAIL.n314 9.3005
R1350 VTAIL.n293 VTAIL.n292 9.3005
R1351 VTAIL.n291 VTAIL.n290 9.3005
R1352 VTAIL.n226 VTAIL.n225 9.3005
R1353 VTAIL.n285 VTAIL.n284 9.3005
R1354 VTAIL.n283 VTAIL.n282 9.3005
R1355 VTAIL.n230 VTAIL.n229 9.3005
R1356 VTAIL.n277 VTAIL.n276 9.3005
R1357 VTAIL.n275 VTAIL.n274 9.3005
R1358 VTAIL.n234 VTAIL.n233 9.3005
R1359 VTAIL.n144 VTAIL.n143 9.3005
R1360 VTAIL.n146 VTAIL.n145 9.3005
R1361 VTAIL.n137 VTAIL.n136 9.3005
R1362 VTAIL.n152 VTAIL.n151 9.3005
R1363 VTAIL.n154 VTAIL.n153 9.3005
R1364 VTAIL.n132 VTAIL.n131 9.3005
R1365 VTAIL.n160 VTAIL.n159 9.3005
R1366 VTAIL.n162 VTAIL.n161 9.3005
R1367 VTAIL.n116 VTAIL.n115 9.3005
R1368 VTAIL.n193 VTAIL.n192 9.3005
R1369 VTAIL.n195 VTAIL.n194 9.3005
R1370 VTAIL.n112 VTAIL.n111 9.3005
R1371 VTAIL.n201 VTAIL.n200 9.3005
R1372 VTAIL.n203 VTAIL.n202 9.3005
R1373 VTAIL.n108 VTAIL.n107 9.3005
R1374 VTAIL.n209 VTAIL.n208 9.3005
R1375 VTAIL.n187 VTAIL.n186 9.3005
R1376 VTAIL.n185 VTAIL.n184 9.3005
R1377 VTAIL.n120 VTAIL.n119 9.3005
R1378 VTAIL.n179 VTAIL.n178 9.3005
R1379 VTAIL.n177 VTAIL.n176 9.3005
R1380 VTAIL.n124 VTAIL.n123 9.3005
R1381 VTAIL.n171 VTAIL.n170 9.3005
R1382 VTAIL.n169 VTAIL.n168 9.3005
R1383 VTAIL.n128 VTAIL.n127 9.3005
R1384 VTAIL.n358 VTAIL.n348 8.92171
R1385 VTAIL.n392 VTAIL.n391 8.92171
R1386 VTAIL.n407 VTAIL.n326 8.92171
R1387 VTAIL.n40 VTAIL.n30 8.92171
R1388 VTAIL.n74 VTAIL.n73 8.92171
R1389 VTAIL.n89 VTAIL.n8 8.92171
R1390 VTAIL.n301 VTAIL.n220 8.92171
R1391 VTAIL.n286 VTAIL.n285 8.92171
R1392 VTAIL.n253 VTAIL.n243 8.92171
R1393 VTAIL.n195 VTAIL.n114 8.92171
R1394 VTAIL.n180 VTAIL.n179 8.92171
R1395 VTAIL.n147 VTAIL.n137 8.92171
R1396 VTAIL.n357 VTAIL.n350 8.14595
R1397 VTAIL.n395 VTAIL.n332 8.14595
R1398 VTAIL.n404 VTAIL.n403 8.14595
R1399 VTAIL.n39 VTAIL.n32 8.14595
R1400 VTAIL.n77 VTAIL.n14 8.14595
R1401 VTAIL.n86 VTAIL.n85 8.14595
R1402 VTAIL.n298 VTAIL.n297 8.14595
R1403 VTAIL.n289 VTAIL.n226 8.14595
R1404 VTAIL.n252 VTAIL.n245 8.14595
R1405 VTAIL.n192 VTAIL.n191 8.14595
R1406 VTAIL.n183 VTAIL.n120 8.14595
R1407 VTAIL.n146 VTAIL.n139 8.14595
R1408 VTAIL.n422 VTAIL.n318 7.75445
R1409 VTAIL.n104 VTAIL.n0 7.75445
R1410 VTAIL.n316 VTAIL.n212 7.75445
R1411 VTAIL.n210 VTAIL.n106 7.75445
R1412 VTAIL.n354 VTAIL.n353 7.3702
R1413 VTAIL.n396 VTAIL.n330 7.3702
R1414 VTAIL.n400 VTAIL.n328 7.3702
R1415 VTAIL.n36 VTAIL.n35 7.3702
R1416 VTAIL.n78 VTAIL.n12 7.3702
R1417 VTAIL.n82 VTAIL.n10 7.3702
R1418 VTAIL.n294 VTAIL.n222 7.3702
R1419 VTAIL.n290 VTAIL.n224 7.3702
R1420 VTAIL.n249 VTAIL.n248 7.3702
R1421 VTAIL.n188 VTAIL.n116 7.3702
R1422 VTAIL.n184 VTAIL.n118 7.3702
R1423 VTAIL.n143 VTAIL.n142 7.3702
R1424 VTAIL.n399 VTAIL.n330 6.59444
R1425 VTAIL.n400 VTAIL.n399 6.59444
R1426 VTAIL.n81 VTAIL.n12 6.59444
R1427 VTAIL.n82 VTAIL.n81 6.59444
R1428 VTAIL.n294 VTAIL.n293 6.59444
R1429 VTAIL.n293 VTAIL.n224 6.59444
R1430 VTAIL.n188 VTAIL.n187 6.59444
R1431 VTAIL.n187 VTAIL.n118 6.59444
R1432 VTAIL.n420 VTAIL.n318 6.08283
R1433 VTAIL.n102 VTAIL.n0 6.08283
R1434 VTAIL.n314 VTAIL.n212 6.08283
R1435 VTAIL.n208 VTAIL.n106 6.08283
R1436 VTAIL.n354 VTAIL.n350 5.81868
R1437 VTAIL.n396 VTAIL.n395 5.81868
R1438 VTAIL.n403 VTAIL.n328 5.81868
R1439 VTAIL.n36 VTAIL.n32 5.81868
R1440 VTAIL.n78 VTAIL.n77 5.81868
R1441 VTAIL.n85 VTAIL.n10 5.81868
R1442 VTAIL.n297 VTAIL.n222 5.81868
R1443 VTAIL.n290 VTAIL.n289 5.81868
R1444 VTAIL.n249 VTAIL.n245 5.81868
R1445 VTAIL.n191 VTAIL.n116 5.81868
R1446 VTAIL.n184 VTAIL.n183 5.81868
R1447 VTAIL.n143 VTAIL.n139 5.81868
R1448 VTAIL.n358 VTAIL.n357 5.04292
R1449 VTAIL.n392 VTAIL.n332 5.04292
R1450 VTAIL.n404 VTAIL.n326 5.04292
R1451 VTAIL.n40 VTAIL.n39 5.04292
R1452 VTAIL.n74 VTAIL.n14 5.04292
R1453 VTAIL.n86 VTAIL.n8 5.04292
R1454 VTAIL.n298 VTAIL.n220 5.04292
R1455 VTAIL.n286 VTAIL.n226 5.04292
R1456 VTAIL.n253 VTAIL.n252 5.04292
R1457 VTAIL.n192 VTAIL.n114 5.04292
R1458 VTAIL.n180 VTAIL.n120 5.04292
R1459 VTAIL.n147 VTAIL.n146 5.04292
R1460 VTAIL.n361 VTAIL.n348 4.26717
R1461 VTAIL.n391 VTAIL.n334 4.26717
R1462 VTAIL.n408 VTAIL.n407 4.26717
R1463 VTAIL.n43 VTAIL.n30 4.26717
R1464 VTAIL.n73 VTAIL.n16 4.26717
R1465 VTAIL.n90 VTAIL.n89 4.26717
R1466 VTAIL.n302 VTAIL.n301 4.26717
R1467 VTAIL.n285 VTAIL.n228 4.26717
R1468 VTAIL.n256 VTAIL.n243 4.26717
R1469 VTAIL.n196 VTAIL.n195 4.26717
R1470 VTAIL.n179 VTAIL.n122 4.26717
R1471 VTAIL.n150 VTAIL.n137 4.26717
R1472 VTAIL.n362 VTAIL.n346 3.49141
R1473 VTAIL.n388 VTAIL.n387 3.49141
R1474 VTAIL.n411 VTAIL.n324 3.49141
R1475 VTAIL.n44 VTAIL.n28 3.49141
R1476 VTAIL.n70 VTAIL.n69 3.49141
R1477 VTAIL.n93 VTAIL.n6 3.49141
R1478 VTAIL.n305 VTAIL.n218 3.49141
R1479 VTAIL.n282 VTAIL.n281 3.49141
R1480 VTAIL.n257 VTAIL.n241 3.49141
R1481 VTAIL.n199 VTAIL.n112 3.49141
R1482 VTAIL.n176 VTAIL.n175 3.49141
R1483 VTAIL.n151 VTAIL.n135 3.49141
R1484 VTAIL.n366 VTAIL.n365 2.71565
R1485 VTAIL.n384 VTAIL.n336 2.71565
R1486 VTAIL.n412 VTAIL.n322 2.71565
R1487 VTAIL.n48 VTAIL.n47 2.71565
R1488 VTAIL.n66 VTAIL.n18 2.71565
R1489 VTAIL.n94 VTAIL.n4 2.71565
R1490 VTAIL.n306 VTAIL.n216 2.71565
R1491 VTAIL.n278 VTAIL.n230 2.71565
R1492 VTAIL.n261 VTAIL.n260 2.71565
R1493 VTAIL.n200 VTAIL.n110 2.71565
R1494 VTAIL.n172 VTAIL.n124 2.71565
R1495 VTAIL.n155 VTAIL.n154 2.71565
R1496 VTAIL.n250 VTAIL.n246 2.41282
R1497 VTAIL.n144 VTAIL.n140 2.41282
R1498 VTAIL.n355 VTAIL.n351 2.41282
R1499 VTAIL.n37 VTAIL.n33 2.41282
R1500 VTAIL.n370 VTAIL.n344 1.93989
R1501 VTAIL.n383 VTAIL.n338 1.93989
R1502 VTAIL.n416 VTAIL.n415 1.93989
R1503 VTAIL.n52 VTAIL.n26 1.93989
R1504 VTAIL.n65 VTAIL.n20 1.93989
R1505 VTAIL.n98 VTAIL.n97 1.93989
R1506 VTAIL.n310 VTAIL.n309 1.93989
R1507 VTAIL.n277 VTAIL.n232 1.93989
R1508 VTAIL.n264 VTAIL.n238 1.93989
R1509 VTAIL.n204 VTAIL.n203 1.93989
R1510 VTAIL.n171 VTAIL.n126 1.93989
R1511 VTAIL.n158 VTAIL.n132 1.93989
R1512 VTAIL.n371 VTAIL.n342 1.16414
R1513 VTAIL.n380 VTAIL.n379 1.16414
R1514 VTAIL.n419 VTAIL.n320 1.16414
R1515 VTAIL.n53 VTAIL.n24 1.16414
R1516 VTAIL.n62 VTAIL.n61 1.16414
R1517 VTAIL.n101 VTAIL.n2 1.16414
R1518 VTAIL.n313 VTAIL.n214 1.16414
R1519 VTAIL.n274 VTAIL.n273 1.16414
R1520 VTAIL.n265 VTAIL.n236 1.16414
R1521 VTAIL.n207 VTAIL.n108 1.16414
R1522 VTAIL.n168 VTAIL.n167 1.16414
R1523 VTAIL.n159 VTAIL.n130 1.16414
R1524 VTAIL.n317 VTAIL.n211 0.724638
R1525 VTAIL VTAIL.n105 0.655672
R1526 VTAIL.n375 VTAIL.n374 0.388379
R1527 VTAIL.n376 VTAIL.n340 0.388379
R1528 VTAIL.n57 VTAIL.n56 0.388379
R1529 VTAIL.n58 VTAIL.n22 0.388379
R1530 VTAIL.n270 VTAIL.n234 0.388379
R1531 VTAIL.n269 VTAIL.n268 0.388379
R1532 VTAIL.n164 VTAIL.n128 0.388379
R1533 VTAIL.n163 VTAIL.n162 0.388379
R1534 VTAIL.n356 VTAIL.n355 0.155672
R1535 VTAIL.n356 VTAIL.n347 0.155672
R1536 VTAIL.n363 VTAIL.n347 0.155672
R1537 VTAIL.n364 VTAIL.n363 0.155672
R1538 VTAIL.n364 VTAIL.n343 0.155672
R1539 VTAIL.n372 VTAIL.n343 0.155672
R1540 VTAIL.n373 VTAIL.n372 0.155672
R1541 VTAIL.n373 VTAIL.n339 0.155672
R1542 VTAIL.n381 VTAIL.n339 0.155672
R1543 VTAIL.n382 VTAIL.n381 0.155672
R1544 VTAIL.n382 VTAIL.n335 0.155672
R1545 VTAIL.n389 VTAIL.n335 0.155672
R1546 VTAIL.n390 VTAIL.n389 0.155672
R1547 VTAIL.n390 VTAIL.n331 0.155672
R1548 VTAIL.n397 VTAIL.n331 0.155672
R1549 VTAIL.n398 VTAIL.n397 0.155672
R1550 VTAIL.n398 VTAIL.n327 0.155672
R1551 VTAIL.n405 VTAIL.n327 0.155672
R1552 VTAIL.n406 VTAIL.n405 0.155672
R1553 VTAIL.n406 VTAIL.n323 0.155672
R1554 VTAIL.n413 VTAIL.n323 0.155672
R1555 VTAIL.n414 VTAIL.n413 0.155672
R1556 VTAIL.n414 VTAIL.n319 0.155672
R1557 VTAIL.n421 VTAIL.n319 0.155672
R1558 VTAIL.n38 VTAIL.n37 0.155672
R1559 VTAIL.n38 VTAIL.n29 0.155672
R1560 VTAIL.n45 VTAIL.n29 0.155672
R1561 VTAIL.n46 VTAIL.n45 0.155672
R1562 VTAIL.n46 VTAIL.n25 0.155672
R1563 VTAIL.n54 VTAIL.n25 0.155672
R1564 VTAIL.n55 VTAIL.n54 0.155672
R1565 VTAIL.n55 VTAIL.n21 0.155672
R1566 VTAIL.n63 VTAIL.n21 0.155672
R1567 VTAIL.n64 VTAIL.n63 0.155672
R1568 VTAIL.n64 VTAIL.n17 0.155672
R1569 VTAIL.n71 VTAIL.n17 0.155672
R1570 VTAIL.n72 VTAIL.n71 0.155672
R1571 VTAIL.n72 VTAIL.n13 0.155672
R1572 VTAIL.n79 VTAIL.n13 0.155672
R1573 VTAIL.n80 VTAIL.n79 0.155672
R1574 VTAIL.n80 VTAIL.n9 0.155672
R1575 VTAIL.n87 VTAIL.n9 0.155672
R1576 VTAIL.n88 VTAIL.n87 0.155672
R1577 VTAIL.n88 VTAIL.n5 0.155672
R1578 VTAIL.n95 VTAIL.n5 0.155672
R1579 VTAIL.n96 VTAIL.n95 0.155672
R1580 VTAIL.n96 VTAIL.n1 0.155672
R1581 VTAIL.n103 VTAIL.n1 0.155672
R1582 VTAIL.n315 VTAIL.n213 0.155672
R1583 VTAIL.n308 VTAIL.n213 0.155672
R1584 VTAIL.n308 VTAIL.n307 0.155672
R1585 VTAIL.n307 VTAIL.n217 0.155672
R1586 VTAIL.n300 VTAIL.n217 0.155672
R1587 VTAIL.n300 VTAIL.n299 0.155672
R1588 VTAIL.n299 VTAIL.n221 0.155672
R1589 VTAIL.n292 VTAIL.n221 0.155672
R1590 VTAIL.n292 VTAIL.n291 0.155672
R1591 VTAIL.n291 VTAIL.n225 0.155672
R1592 VTAIL.n284 VTAIL.n225 0.155672
R1593 VTAIL.n284 VTAIL.n283 0.155672
R1594 VTAIL.n283 VTAIL.n229 0.155672
R1595 VTAIL.n276 VTAIL.n229 0.155672
R1596 VTAIL.n276 VTAIL.n275 0.155672
R1597 VTAIL.n275 VTAIL.n233 0.155672
R1598 VTAIL.n267 VTAIL.n233 0.155672
R1599 VTAIL.n267 VTAIL.n266 0.155672
R1600 VTAIL.n266 VTAIL.n237 0.155672
R1601 VTAIL.n259 VTAIL.n237 0.155672
R1602 VTAIL.n259 VTAIL.n258 0.155672
R1603 VTAIL.n258 VTAIL.n242 0.155672
R1604 VTAIL.n251 VTAIL.n242 0.155672
R1605 VTAIL.n251 VTAIL.n250 0.155672
R1606 VTAIL.n209 VTAIL.n107 0.155672
R1607 VTAIL.n202 VTAIL.n107 0.155672
R1608 VTAIL.n202 VTAIL.n201 0.155672
R1609 VTAIL.n201 VTAIL.n111 0.155672
R1610 VTAIL.n194 VTAIL.n111 0.155672
R1611 VTAIL.n194 VTAIL.n193 0.155672
R1612 VTAIL.n193 VTAIL.n115 0.155672
R1613 VTAIL.n186 VTAIL.n115 0.155672
R1614 VTAIL.n186 VTAIL.n185 0.155672
R1615 VTAIL.n185 VTAIL.n119 0.155672
R1616 VTAIL.n178 VTAIL.n119 0.155672
R1617 VTAIL.n178 VTAIL.n177 0.155672
R1618 VTAIL.n177 VTAIL.n123 0.155672
R1619 VTAIL.n170 VTAIL.n123 0.155672
R1620 VTAIL.n170 VTAIL.n169 0.155672
R1621 VTAIL.n169 VTAIL.n127 0.155672
R1622 VTAIL.n161 VTAIL.n127 0.155672
R1623 VTAIL.n161 VTAIL.n160 0.155672
R1624 VTAIL.n160 VTAIL.n131 0.155672
R1625 VTAIL.n153 VTAIL.n131 0.155672
R1626 VTAIL.n153 VTAIL.n152 0.155672
R1627 VTAIL.n152 VTAIL.n136 0.155672
R1628 VTAIL.n145 VTAIL.n136 0.155672
R1629 VTAIL.n145 VTAIL.n144 0.155672
R1630 VTAIL VTAIL.n423 0.0694655
R1631 VDD2.n206 VDD2.n205 585
R1632 VDD2.n204 VDD2.n203 585
R1633 VDD2.n109 VDD2.n108 585
R1634 VDD2.n198 VDD2.n197 585
R1635 VDD2.n196 VDD2.n195 585
R1636 VDD2.n113 VDD2.n112 585
R1637 VDD2.n190 VDD2.n189 585
R1638 VDD2.n188 VDD2.n187 585
R1639 VDD2.n117 VDD2.n116 585
R1640 VDD2.n182 VDD2.n181 585
R1641 VDD2.n180 VDD2.n179 585
R1642 VDD2.n121 VDD2.n120 585
R1643 VDD2.n174 VDD2.n173 585
R1644 VDD2.n172 VDD2.n171 585
R1645 VDD2.n125 VDD2.n124 585
R1646 VDD2.n166 VDD2.n165 585
R1647 VDD2.n164 VDD2.n163 585
R1648 VDD2.n162 VDD2.n128 585
R1649 VDD2.n132 VDD2.n129 585
R1650 VDD2.n157 VDD2.n156 585
R1651 VDD2.n155 VDD2.n154 585
R1652 VDD2.n134 VDD2.n133 585
R1653 VDD2.n149 VDD2.n148 585
R1654 VDD2.n147 VDD2.n146 585
R1655 VDD2.n138 VDD2.n137 585
R1656 VDD2.n141 VDD2.n140 585
R1657 VDD2.n35 VDD2.n34 585
R1658 VDD2.n32 VDD2.n31 585
R1659 VDD2.n41 VDD2.n40 585
R1660 VDD2.n43 VDD2.n42 585
R1661 VDD2.n28 VDD2.n27 585
R1662 VDD2.n49 VDD2.n48 585
R1663 VDD2.n52 VDD2.n51 585
R1664 VDD2.n50 VDD2.n24 585
R1665 VDD2.n57 VDD2.n23 585
R1666 VDD2.n59 VDD2.n58 585
R1667 VDD2.n61 VDD2.n60 585
R1668 VDD2.n20 VDD2.n19 585
R1669 VDD2.n67 VDD2.n66 585
R1670 VDD2.n69 VDD2.n68 585
R1671 VDD2.n16 VDD2.n15 585
R1672 VDD2.n75 VDD2.n74 585
R1673 VDD2.n77 VDD2.n76 585
R1674 VDD2.n12 VDD2.n11 585
R1675 VDD2.n83 VDD2.n82 585
R1676 VDD2.n85 VDD2.n84 585
R1677 VDD2.n8 VDD2.n7 585
R1678 VDD2.n91 VDD2.n90 585
R1679 VDD2.n93 VDD2.n92 585
R1680 VDD2.n4 VDD2.n3 585
R1681 VDD2.n99 VDD2.n98 585
R1682 VDD2.n101 VDD2.n100 585
R1683 VDD2.n205 VDD2.n105 498.474
R1684 VDD2.n100 VDD2.n0 498.474
R1685 VDD2.t0 VDD2.n139 329.036
R1686 VDD2.t1 VDD2.n33 329.036
R1687 VDD2.n205 VDD2.n204 171.744
R1688 VDD2.n204 VDD2.n108 171.744
R1689 VDD2.n197 VDD2.n108 171.744
R1690 VDD2.n197 VDD2.n196 171.744
R1691 VDD2.n196 VDD2.n112 171.744
R1692 VDD2.n189 VDD2.n112 171.744
R1693 VDD2.n189 VDD2.n188 171.744
R1694 VDD2.n188 VDD2.n116 171.744
R1695 VDD2.n181 VDD2.n116 171.744
R1696 VDD2.n181 VDD2.n180 171.744
R1697 VDD2.n180 VDD2.n120 171.744
R1698 VDD2.n173 VDD2.n120 171.744
R1699 VDD2.n173 VDD2.n172 171.744
R1700 VDD2.n172 VDD2.n124 171.744
R1701 VDD2.n165 VDD2.n124 171.744
R1702 VDD2.n165 VDD2.n164 171.744
R1703 VDD2.n164 VDD2.n128 171.744
R1704 VDD2.n132 VDD2.n128 171.744
R1705 VDD2.n156 VDD2.n132 171.744
R1706 VDD2.n156 VDD2.n155 171.744
R1707 VDD2.n155 VDD2.n133 171.744
R1708 VDD2.n148 VDD2.n133 171.744
R1709 VDD2.n148 VDD2.n147 171.744
R1710 VDD2.n147 VDD2.n137 171.744
R1711 VDD2.n140 VDD2.n137 171.744
R1712 VDD2.n34 VDD2.n31 171.744
R1713 VDD2.n41 VDD2.n31 171.744
R1714 VDD2.n42 VDD2.n41 171.744
R1715 VDD2.n42 VDD2.n27 171.744
R1716 VDD2.n49 VDD2.n27 171.744
R1717 VDD2.n51 VDD2.n49 171.744
R1718 VDD2.n51 VDD2.n50 171.744
R1719 VDD2.n50 VDD2.n23 171.744
R1720 VDD2.n59 VDD2.n23 171.744
R1721 VDD2.n60 VDD2.n59 171.744
R1722 VDD2.n60 VDD2.n19 171.744
R1723 VDD2.n67 VDD2.n19 171.744
R1724 VDD2.n68 VDD2.n67 171.744
R1725 VDD2.n68 VDD2.n15 171.744
R1726 VDD2.n75 VDD2.n15 171.744
R1727 VDD2.n76 VDD2.n75 171.744
R1728 VDD2.n76 VDD2.n11 171.744
R1729 VDD2.n83 VDD2.n11 171.744
R1730 VDD2.n84 VDD2.n83 171.744
R1731 VDD2.n84 VDD2.n7 171.744
R1732 VDD2.n91 VDD2.n7 171.744
R1733 VDD2.n92 VDD2.n91 171.744
R1734 VDD2.n92 VDD2.n3 171.744
R1735 VDD2.n99 VDD2.n3 171.744
R1736 VDD2.n100 VDD2.n99 171.744
R1737 VDD2.n210 VDD2.n104 95.0747
R1738 VDD2.n140 VDD2.t0 85.8723
R1739 VDD2.n34 VDD2.t1 85.8723
R1740 VDD2.n210 VDD2.n209 53.5187
R1741 VDD2.n163 VDD2.n162 13.1884
R1742 VDD2.n58 VDD2.n57 13.1884
R1743 VDD2.n207 VDD2.n206 12.8005
R1744 VDD2.n166 VDD2.n127 12.8005
R1745 VDD2.n161 VDD2.n129 12.8005
R1746 VDD2.n56 VDD2.n24 12.8005
R1747 VDD2.n61 VDD2.n22 12.8005
R1748 VDD2.n102 VDD2.n101 12.8005
R1749 VDD2.n203 VDD2.n107 12.0247
R1750 VDD2.n167 VDD2.n125 12.0247
R1751 VDD2.n158 VDD2.n157 12.0247
R1752 VDD2.n53 VDD2.n52 12.0247
R1753 VDD2.n62 VDD2.n20 12.0247
R1754 VDD2.n98 VDD2.n2 12.0247
R1755 VDD2.n202 VDD2.n109 11.249
R1756 VDD2.n171 VDD2.n170 11.249
R1757 VDD2.n154 VDD2.n131 11.249
R1758 VDD2.n48 VDD2.n26 11.249
R1759 VDD2.n66 VDD2.n65 11.249
R1760 VDD2.n97 VDD2.n4 11.249
R1761 VDD2.n141 VDD2.n139 10.7239
R1762 VDD2.n35 VDD2.n33 10.7239
R1763 VDD2.n199 VDD2.n198 10.4732
R1764 VDD2.n174 VDD2.n123 10.4732
R1765 VDD2.n153 VDD2.n134 10.4732
R1766 VDD2.n47 VDD2.n28 10.4732
R1767 VDD2.n69 VDD2.n18 10.4732
R1768 VDD2.n94 VDD2.n93 10.4732
R1769 VDD2.n195 VDD2.n111 9.69747
R1770 VDD2.n175 VDD2.n121 9.69747
R1771 VDD2.n150 VDD2.n149 9.69747
R1772 VDD2.n44 VDD2.n43 9.69747
R1773 VDD2.n70 VDD2.n16 9.69747
R1774 VDD2.n90 VDD2.n6 9.69747
R1775 VDD2.n209 VDD2.n208 9.45567
R1776 VDD2.n104 VDD2.n103 9.45567
R1777 VDD2.n143 VDD2.n142 9.3005
R1778 VDD2.n145 VDD2.n144 9.3005
R1779 VDD2.n136 VDD2.n135 9.3005
R1780 VDD2.n151 VDD2.n150 9.3005
R1781 VDD2.n153 VDD2.n152 9.3005
R1782 VDD2.n131 VDD2.n130 9.3005
R1783 VDD2.n159 VDD2.n158 9.3005
R1784 VDD2.n161 VDD2.n160 9.3005
R1785 VDD2.n115 VDD2.n114 9.3005
R1786 VDD2.n192 VDD2.n191 9.3005
R1787 VDD2.n194 VDD2.n193 9.3005
R1788 VDD2.n111 VDD2.n110 9.3005
R1789 VDD2.n200 VDD2.n199 9.3005
R1790 VDD2.n202 VDD2.n201 9.3005
R1791 VDD2.n107 VDD2.n106 9.3005
R1792 VDD2.n208 VDD2.n207 9.3005
R1793 VDD2.n186 VDD2.n185 9.3005
R1794 VDD2.n184 VDD2.n183 9.3005
R1795 VDD2.n119 VDD2.n118 9.3005
R1796 VDD2.n178 VDD2.n177 9.3005
R1797 VDD2.n176 VDD2.n175 9.3005
R1798 VDD2.n123 VDD2.n122 9.3005
R1799 VDD2.n170 VDD2.n169 9.3005
R1800 VDD2.n168 VDD2.n167 9.3005
R1801 VDD2.n127 VDD2.n126 9.3005
R1802 VDD2.n79 VDD2.n78 9.3005
R1803 VDD2.n14 VDD2.n13 9.3005
R1804 VDD2.n73 VDD2.n72 9.3005
R1805 VDD2.n71 VDD2.n70 9.3005
R1806 VDD2.n18 VDD2.n17 9.3005
R1807 VDD2.n65 VDD2.n64 9.3005
R1808 VDD2.n63 VDD2.n62 9.3005
R1809 VDD2.n22 VDD2.n21 9.3005
R1810 VDD2.n37 VDD2.n36 9.3005
R1811 VDD2.n39 VDD2.n38 9.3005
R1812 VDD2.n30 VDD2.n29 9.3005
R1813 VDD2.n45 VDD2.n44 9.3005
R1814 VDD2.n47 VDD2.n46 9.3005
R1815 VDD2.n26 VDD2.n25 9.3005
R1816 VDD2.n54 VDD2.n53 9.3005
R1817 VDD2.n56 VDD2.n55 9.3005
R1818 VDD2.n81 VDD2.n80 9.3005
R1819 VDD2.n10 VDD2.n9 9.3005
R1820 VDD2.n87 VDD2.n86 9.3005
R1821 VDD2.n89 VDD2.n88 9.3005
R1822 VDD2.n6 VDD2.n5 9.3005
R1823 VDD2.n95 VDD2.n94 9.3005
R1824 VDD2.n97 VDD2.n96 9.3005
R1825 VDD2.n2 VDD2.n1 9.3005
R1826 VDD2.n103 VDD2.n102 9.3005
R1827 VDD2.n194 VDD2.n113 8.92171
R1828 VDD2.n179 VDD2.n178 8.92171
R1829 VDD2.n146 VDD2.n136 8.92171
R1830 VDD2.n40 VDD2.n30 8.92171
R1831 VDD2.n74 VDD2.n73 8.92171
R1832 VDD2.n89 VDD2.n8 8.92171
R1833 VDD2.n191 VDD2.n190 8.14595
R1834 VDD2.n182 VDD2.n119 8.14595
R1835 VDD2.n145 VDD2.n138 8.14595
R1836 VDD2.n39 VDD2.n32 8.14595
R1837 VDD2.n77 VDD2.n14 8.14595
R1838 VDD2.n86 VDD2.n85 8.14595
R1839 VDD2.n209 VDD2.n105 7.75445
R1840 VDD2.n104 VDD2.n0 7.75445
R1841 VDD2.n187 VDD2.n115 7.3702
R1842 VDD2.n183 VDD2.n117 7.3702
R1843 VDD2.n142 VDD2.n141 7.3702
R1844 VDD2.n36 VDD2.n35 7.3702
R1845 VDD2.n78 VDD2.n12 7.3702
R1846 VDD2.n82 VDD2.n10 7.3702
R1847 VDD2.n187 VDD2.n186 6.59444
R1848 VDD2.n186 VDD2.n117 6.59444
R1849 VDD2.n81 VDD2.n12 6.59444
R1850 VDD2.n82 VDD2.n81 6.59444
R1851 VDD2.n207 VDD2.n105 6.08283
R1852 VDD2.n102 VDD2.n0 6.08283
R1853 VDD2.n190 VDD2.n115 5.81868
R1854 VDD2.n183 VDD2.n182 5.81868
R1855 VDD2.n142 VDD2.n138 5.81868
R1856 VDD2.n36 VDD2.n32 5.81868
R1857 VDD2.n78 VDD2.n77 5.81868
R1858 VDD2.n85 VDD2.n10 5.81868
R1859 VDD2.n191 VDD2.n113 5.04292
R1860 VDD2.n179 VDD2.n119 5.04292
R1861 VDD2.n146 VDD2.n145 5.04292
R1862 VDD2.n40 VDD2.n39 5.04292
R1863 VDD2.n74 VDD2.n14 5.04292
R1864 VDD2.n86 VDD2.n8 5.04292
R1865 VDD2.n195 VDD2.n194 4.26717
R1866 VDD2.n178 VDD2.n121 4.26717
R1867 VDD2.n149 VDD2.n136 4.26717
R1868 VDD2.n43 VDD2.n30 4.26717
R1869 VDD2.n73 VDD2.n16 4.26717
R1870 VDD2.n90 VDD2.n89 4.26717
R1871 VDD2.n198 VDD2.n111 3.49141
R1872 VDD2.n175 VDD2.n174 3.49141
R1873 VDD2.n150 VDD2.n134 3.49141
R1874 VDD2.n44 VDD2.n28 3.49141
R1875 VDD2.n70 VDD2.n69 3.49141
R1876 VDD2.n93 VDD2.n6 3.49141
R1877 VDD2.n199 VDD2.n109 2.71565
R1878 VDD2.n171 VDD2.n123 2.71565
R1879 VDD2.n154 VDD2.n153 2.71565
R1880 VDD2.n48 VDD2.n47 2.71565
R1881 VDD2.n66 VDD2.n18 2.71565
R1882 VDD2.n94 VDD2.n4 2.71565
R1883 VDD2.n143 VDD2.n139 2.41282
R1884 VDD2.n37 VDD2.n33 2.41282
R1885 VDD2.n203 VDD2.n202 1.93989
R1886 VDD2.n170 VDD2.n125 1.93989
R1887 VDD2.n157 VDD2.n131 1.93989
R1888 VDD2.n52 VDD2.n26 1.93989
R1889 VDD2.n65 VDD2.n20 1.93989
R1890 VDD2.n98 VDD2.n97 1.93989
R1891 VDD2.n206 VDD2.n107 1.16414
R1892 VDD2.n167 VDD2.n166 1.16414
R1893 VDD2.n158 VDD2.n129 1.16414
R1894 VDD2.n53 VDD2.n24 1.16414
R1895 VDD2.n62 VDD2.n61 1.16414
R1896 VDD2.n101 VDD2.n2 1.16414
R1897 VDD2.n163 VDD2.n127 0.388379
R1898 VDD2.n162 VDD2.n161 0.388379
R1899 VDD2.n57 VDD2.n56 0.388379
R1900 VDD2.n58 VDD2.n22 0.388379
R1901 VDD2 VDD2.n210 0.185845
R1902 VDD2.n208 VDD2.n106 0.155672
R1903 VDD2.n201 VDD2.n106 0.155672
R1904 VDD2.n201 VDD2.n200 0.155672
R1905 VDD2.n200 VDD2.n110 0.155672
R1906 VDD2.n193 VDD2.n110 0.155672
R1907 VDD2.n193 VDD2.n192 0.155672
R1908 VDD2.n192 VDD2.n114 0.155672
R1909 VDD2.n185 VDD2.n114 0.155672
R1910 VDD2.n185 VDD2.n184 0.155672
R1911 VDD2.n184 VDD2.n118 0.155672
R1912 VDD2.n177 VDD2.n118 0.155672
R1913 VDD2.n177 VDD2.n176 0.155672
R1914 VDD2.n176 VDD2.n122 0.155672
R1915 VDD2.n169 VDD2.n122 0.155672
R1916 VDD2.n169 VDD2.n168 0.155672
R1917 VDD2.n168 VDD2.n126 0.155672
R1918 VDD2.n160 VDD2.n126 0.155672
R1919 VDD2.n160 VDD2.n159 0.155672
R1920 VDD2.n159 VDD2.n130 0.155672
R1921 VDD2.n152 VDD2.n130 0.155672
R1922 VDD2.n152 VDD2.n151 0.155672
R1923 VDD2.n151 VDD2.n135 0.155672
R1924 VDD2.n144 VDD2.n135 0.155672
R1925 VDD2.n144 VDD2.n143 0.155672
R1926 VDD2.n38 VDD2.n37 0.155672
R1927 VDD2.n38 VDD2.n29 0.155672
R1928 VDD2.n45 VDD2.n29 0.155672
R1929 VDD2.n46 VDD2.n45 0.155672
R1930 VDD2.n46 VDD2.n25 0.155672
R1931 VDD2.n54 VDD2.n25 0.155672
R1932 VDD2.n55 VDD2.n54 0.155672
R1933 VDD2.n55 VDD2.n21 0.155672
R1934 VDD2.n63 VDD2.n21 0.155672
R1935 VDD2.n64 VDD2.n63 0.155672
R1936 VDD2.n64 VDD2.n17 0.155672
R1937 VDD2.n71 VDD2.n17 0.155672
R1938 VDD2.n72 VDD2.n71 0.155672
R1939 VDD2.n72 VDD2.n13 0.155672
R1940 VDD2.n79 VDD2.n13 0.155672
R1941 VDD2.n80 VDD2.n79 0.155672
R1942 VDD2.n80 VDD2.n9 0.155672
R1943 VDD2.n87 VDD2.n9 0.155672
R1944 VDD2.n88 VDD2.n87 0.155672
R1945 VDD2.n88 VDD2.n5 0.155672
R1946 VDD2.n95 VDD2.n5 0.155672
R1947 VDD2.n96 VDD2.n95 0.155672
R1948 VDD2.n96 VDD2.n1 0.155672
R1949 VDD2.n103 VDD2.n1 0.155672
R1950 VP.n0 VP.t0 2163.15
R1951 VP.n0 VP.t1 2118.96
R1952 VP VP.n0 0.0516364
R1953 VDD1.n101 VDD1.n100 585
R1954 VDD1.n99 VDD1.n98 585
R1955 VDD1.n4 VDD1.n3 585
R1956 VDD1.n93 VDD1.n92 585
R1957 VDD1.n91 VDD1.n90 585
R1958 VDD1.n8 VDD1.n7 585
R1959 VDD1.n85 VDD1.n84 585
R1960 VDD1.n83 VDD1.n82 585
R1961 VDD1.n12 VDD1.n11 585
R1962 VDD1.n77 VDD1.n76 585
R1963 VDD1.n75 VDD1.n74 585
R1964 VDD1.n16 VDD1.n15 585
R1965 VDD1.n69 VDD1.n68 585
R1966 VDD1.n67 VDD1.n66 585
R1967 VDD1.n20 VDD1.n19 585
R1968 VDD1.n61 VDD1.n60 585
R1969 VDD1.n59 VDD1.n58 585
R1970 VDD1.n57 VDD1.n23 585
R1971 VDD1.n27 VDD1.n24 585
R1972 VDD1.n52 VDD1.n51 585
R1973 VDD1.n50 VDD1.n49 585
R1974 VDD1.n29 VDD1.n28 585
R1975 VDD1.n44 VDD1.n43 585
R1976 VDD1.n42 VDD1.n41 585
R1977 VDD1.n33 VDD1.n32 585
R1978 VDD1.n36 VDD1.n35 585
R1979 VDD1.n140 VDD1.n139 585
R1980 VDD1.n137 VDD1.n136 585
R1981 VDD1.n146 VDD1.n145 585
R1982 VDD1.n148 VDD1.n147 585
R1983 VDD1.n133 VDD1.n132 585
R1984 VDD1.n154 VDD1.n153 585
R1985 VDD1.n157 VDD1.n156 585
R1986 VDD1.n155 VDD1.n129 585
R1987 VDD1.n162 VDD1.n128 585
R1988 VDD1.n164 VDD1.n163 585
R1989 VDD1.n166 VDD1.n165 585
R1990 VDD1.n125 VDD1.n124 585
R1991 VDD1.n172 VDD1.n171 585
R1992 VDD1.n174 VDD1.n173 585
R1993 VDD1.n121 VDD1.n120 585
R1994 VDD1.n180 VDD1.n179 585
R1995 VDD1.n182 VDD1.n181 585
R1996 VDD1.n117 VDD1.n116 585
R1997 VDD1.n188 VDD1.n187 585
R1998 VDD1.n190 VDD1.n189 585
R1999 VDD1.n113 VDD1.n112 585
R2000 VDD1.n196 VDD1.n195 585
R2001 VDD1.n198 VDD1.n197 585
R2002 VDD1.n109 VDD1.n108 585
R2003 VDD1.n204 VDD1.n203 585
R2004 VDD1.n206 VDD1.n205 585
R2005 VDD1.n100 VDD1.n0 498.474
R2006 VDD1.n205 VDD1.n105 498.474
R2007 VDD1.t1 VDD1.n34 329.036
R2008 VDD1.t0 VDD1.n138 329.036
R2009 VDD1.n100 VDD1.n99 171.744
R2010 VDD1.n99 VDD1.n3 171.744
R2011 VDD1.n92 VDD1.n3 171.744
R2012 VDD1.n92 VDD1.n91 171.744
R2013 VDD1.n91 VDD1.n7 171.744
R2014 VDD1.n84 VDD1.n7 171.744
R2015 VDD1.n84 VDD1.n83 171.744
R2016 VDD1.n83 VDD1.n11 171.744
R2017 VDD1.n76 VDD1.n11 171.744
R2018 VDD1.n76 VDD1.n75 171.744
R2019 VDD1.n75 VDD1.n15 171.744
R2020 VDD1.n68 VDD1.n15 171.744
R2021 VDD1.n68 VDD1.n67 171.744
R2022 VDD1.n67 VDD1.n19 171.744
R2023 VDD1.n60 VDD1.n19 171.744
R2024 VDD1.n60 VDD1.n59 171.744
R2025 VDD1.n59 VDD1.n23 171.744
R2026 VDD1.n27 VDD1.n23 171.744
R2027 VDD1.n51 VDD1.n27 171.744
R2028 VDD1.n51 VDD1.n50 171.744
R2029 VDD1.n50 VDD1.n28 171.744
R2030 VDD1.n43 VDD1.n28 171.744
R2031 VDD1.n43 VDD1.n42 171.744
R2032 VDD1.n42 VDD1.n32 171.744
R2033 VDD1.n35 VDD1.n32 171.744
R2034 VDD1.n139 VDD1.n136 171.744
R2035 VDD1.n146 VDD1.n136 171.744
R2036 VDD1.n147 VDD1.n146 171.744
R2037 VDD1.n147 VDD1.n132 171.744
R2038 VDD1.n154 VDD1.n132 171.744
R2039 VDD1.n156 VDD1.n154 171.744
R2040 VDD1.n156 VDD1.n155 171.744
R2041 VDD1.n155 VDD1.n128 171.744
R2042 VDD1.n164 VDD1.n128 171.744
R2043 VDD1.n165 VDD1.n164 171.744
R2044 VDD1.n165 VDD1.n124 171.744
R2045 VDD1.n172 VDD1.n124 171.744
R2046 VDD1.n173 VDD1.n172 171.744
R2047 VDD1.n173 VDD1.n120 171.744
R2048 VDD1.n180 VDD1.n120 171.744
R2049 VDD1.n181 VDD1.n180 171.744
R2050 VDD1.n181 VDD1.n116 171.744
R2051 VDD1.n188 VDD1.n116 171.744
R2052 VDD1.n189 VDD1.n188 171.744
R2053 VDD1.n189 VDD1.n112 171.744
R2054 VDD1.n196 VDD1.n112 171.744
R2055 VDD1.n197 VDD1.n196 171.744
R2056 VDD1.n197 VDD1.n108 171.744
R2057 VDD1.n204 VDD1.n108 171.744
R2058 VDD1.n205 VDD1.n204 171.744
R2059 VDD1 VDD1.n209 95.7267
R2060 VDD1.n35 VDD1.t1 85.8723
R2061 VDD1.n139 VDD1.t0 85.8723
R2062 VDD1 VDD1.n104 53.704
R2063 VDD1.n58 VDD1.n57 13.1884
R2064 VDD1.n163 VDD1.n162 13.1884
R2065 VDD1.n102 VDD1.n101 12.8005
R2066 VDD1.n61 VDD1.n22 12.8005
R2067 VDD1.n56 VDD1.n24 12.8005
R2068 VDD1.n161 VDD1.n129 12.8005
R2069 VDD1.n166 VDD1.n127 12.8005
R2070 VDD1.n207 VDD1.n206 12.8005
R2071 VDD1.n98 VDD1.n2 12.0247
R2072 VDD1.n62 VDD1.n20 12.0247
R2073 VDD1.n53 VDD1.n52 12.0247
R2074 VDD1.n158 VDD1.n157 12.0247
R2075 VDD1.n167 VDD1.n125 12.0247
R2076 VDD1.n203 VDD1.n107 12.0247
R2077 VDD1.n97 VDD1.n4 11.249
R2078 VDD1.n66 VDD1.n65 11.249
R2079 VDD1.n49 VDD1.n26 11.249
R2080 VDD1.n153 VDD1.n131 11.249
R2081 VDD1.n171 VDD1.n170 11.249
R2082 VDD1.n202 VDD1.n109 11.249
R2083 VDD1.n36 VDD1.n34 10.7239
R2084 VDD1.n140 VDD1.n138 10.7239
R2085 VDD1.n94 VDD1.n93 10.4732
R2086 VDD1.n69 VDD1.n18 10.4732
R2087 VDD1.n48 VDD1.n29 10.4732
R2088 VDD1.n152 VDD1.n133 10.4732
R2089 VDD1.n174 VDD1.n123 10.4732
R2090 VDD1.n199 VDD1.n198 10.4732
R2091 VDD1.n90 VDD1.n6 9.69747
R2092 VDD1.n70 VDD1.n16 9.69747
R2093 VDD1.n45 VDD1.n44 9.69747
R2094 VDD1.n149 VDD1.n148 9.69747
R2095 VDD1.n175 VDD1.n121 9.69747
R2096 VDD1.n195 VDD1.n111 9.69747
R2097 VDD1.n104 VDD1.n103 9.45567
R2098 VDD1.n209 VDD1.n208 9.45567
R2099 VDD1.n38 VDD1.n37 9.3005
R2100 VDD1.n40 VDD1.n39 9.3005
R2101 VDD1.n31 VDD1.n30 9.3005
R2102 VDD1.n46 VDD1.n45 9.3005
R2103 VDD1.n48 VDD1.n47 9.3005
R2104 VDD1.n26 VDD1.n25 9.3005
R2105 VDD1.n54 VDD1.n53 9.3005
R2106 VDD1.n56 VDD1.n55 9.3005
R2107 VDD1.n10 VDD1.n9 9.3005
R2108 VDD1.n87 VDD1.n86 9.3005
R2109 VDD1.n89 VDD1.n88 9.3005
R2110 VDD1.n6 VDD1.n5 9.3005
R2111 VDD1.n95 VDD1.n94 9.3005
R2112 VDD1.n97 VDD1.n96 9.3005
R2113 VDD1.n2 VDD1.n1 9.3005
R2114 VDD1.n103 VDD1.n102 9.3005
R2115 VDD1.n81 VDD1.n80 9.3005
R2116 VDD1.n79 VDD1.n78 9.3005
R2117 VDD1.n14 VDD1.n13 9.3005
R2118 VDD1.n73 VDD1.n72 9.3005
R2119 VDD1.n71 VDD1.n70 9.3005
R2120 VDD1.n18 VDD1.n17 9.3005
R2121 VDD1.n65 VDD1.n64 9.3005
R2122 VDD1.n63 VDD1.n62 9.3005
R2123 VDD1.n22 VDD1.n21 9.3005
R2124 VDD1.n184 VDD1.n183 9.3005
R2125 VDD1.n119 VDD1.n118 9.3005
R2126 VDD1.n178 VDD1.n177 9.3005
R2127 VDD1.n176 VDD1.n175 9.3005
R2128 VDD1.n123 VDD1.n122 9.3005
R2129 VDD1.n170 VDD1.n169 9.3005
R2130 VDD1.n168 VDD1.n167 9.3005
R2131 VDD1.n127 VDD1.n126 9.3005
R2132 VDD1.n142 VDD1.n141 9.3005
R2133 VDD1.n144 VDD1.n143 9.3005
R2134 VDD1.n135 VDD1.n134 9.3005
R2135 VDD1.n150 VDD1.n149 9.3005
R2136 VDD1.n152 VDD1.n151 9.3005
R2137 VDD1.n131 VDD1.n130 9.3005
R2138 VDD1.n159 VDD1.n158 9.3005
R2139 VDD1.n161 VDD1.n160 9.3005
R2140 VDD1.n186 VDD1.n185 9.3005
R2141 VDD1.n115 VDD1.n114 9.3005
R2142 VDD1.n192 VDD1.n191 9.3005
R2143 VDD1.n194 VDD1.n193 9.3005
R2144 VDD1.n111 VDD1.n110 9.3005
R2145 VDD1.n200 VDD1.n199 9.3005
R2146 VDD1.n202 VDD1.n201 9.3005
R2147 VDD1.n107 VDD1.n106 9.3005
R2148 VDD1.n208 VDD1.n207 9.3005
R2149 VDD1.n89 VDD1.n8 8.92171
R2150 VDD1.n74 VDD1.n73 8.92171
R2151 VDD1.n41 VDD1.n31 8.92171
R2152 VDD1.n145 VDD1.n135 8.92171
R2153 VDD1.n179 VDD1.n178 8.92171
R2154 VDD1.n194 VDD1.n113 8.92171
R2155 VDD1.n86 VDD1.n85 8.14595
R2156 VDD1.n77 VDD1.n14 8.14595
R2157 VDD1.n40 VDD1.n33 8.14595
R2158 VDD1.n144 VDD1.n137 8.14595
R2159 VDD1.n182 VDD1.n119 8.14595
R2160 VDD1.n191 VDD1.n190 8.14595
R2161 VDD1.n104 VDD1.n0 7.75445
R2162 VDD1.n209 VDD1.n105 7.75445
R2163 VDD1.n82 VDD1.n10 7.3702
R2164 VDD1.n78 VDD1.n12 7.3702
R2165 VDD1.n37 VDD1.n36 7.3702
R2166 VDD1.n141 VDD1.n140 7.3702
R2167 VDD1.n183 VDD1.n117 7.3702
R2168 VDD1.n187 VDD1.n115 7.3702
R2169 VDD1.n82 VDD1.n81 6.59444
R2170 VDD1.n81 VDD1.n12 6.59444
R2171 VDD1.n186 VDD1.n117 6.59444
R2172 VDD1.n187 VDD1.n186 6.59444
R2173 VDD1.n102 VDD1.n0 6.08283
R2174 VDD1.n207 VDD1.n105 6.08283
R2175 VDD1.n85 VDD1.n10 5.81868
R2176 VDD1.n78 VDD1.n77 5.81868
R2177 VDD1.n37 VDD1.n33 5.81868
R2178 VDD1.n141 VDD1.n137 5.81868
R2179 VDD1.n183 VDD1.n182 5.81868
R2180 VDD1.n190 VDD1.n115 5.81868
R2181 VDD1.n86 VDD1.n8 5.04292
R2182 VDD1.n74 VDD1.n14 5.04292
R2183 VDD1.n41 VDD1.n40 5.04292
R2184 VDD1.n145 VDD1.n144 5.04292
R2185 VDD1.n179 VDD1.n119 5.04292
R2186 VDD1.n191 VDD1.n113 5.04292
R2187 VDD1.n90 VDD1.n89 4.26717
R2188 VDD1.n73 VDD1.n16 4.26717
R2189 VDD1.n44 VDD1.n31 4.26717
R2190 VDD1.n148 VDD1.n135 4.26717
R2191 VDD1.n178 VDD1.n121 4.26717
R2192 VDD1.n195 VDD1.n194 4.26717
R2193 VDD1.n93 VDD1.n6 3.49141
R2194 VDD1.n70 VDD1.n69 3.49141
R2195 VDD1.n45 VDD1.n29 3.49141
R2196 VDD1.n149 VDD1.n133 3.49141
R2197 VDD1.n175 VDD1.n174 3.49141
R2198 VDD1.n198 VDD1.n111 3.49141
R2199 VDD1.n94 VDD1.n4 2.71565
R2200 VDD1.n66 VDD1.n18 2.71565
R2201 VDD1.n49 VDD1.n48 2.71565
R2202 VDD1.n153 VDD1.n152 2.71565
R2203 VDD1.n171 VDD1.n123 2.71565
R2204 VDD1.n199 VDD1.n109 2.71565
R2205 VDD1.n38 VDD1.n34 2.41282
R2206 VDD1.n142 VDD1.n138 2.41282
R2207 VDD1.n98 VDD1.n97 1.93989
R2208 VDD1.n65 VDD1.n20 1.93989
R2209 VDD1.n52 VDD1.n26 1.93989
R2210 VDD1.n157 VDD1.n131 1.93989
R2211 VDD1.n170 VDD1.n125 1.93989
R2212 VDD1.n203 VDD1.n202 1.93989
R2213 VDD1.n101 VDD1.n2 1.16414
R2214 VDD1.n62 VDD1.n61 1.16414
R2215 VDD1.n53 VDD1.n24 1.16414
R2216 VDD1.n158 VDD1.n129 1.16414
R2217 VDD1.n167 VDD1.n166 1.16414
R2218 VDD1.n206 VDD1.n107 1.16414
R2219 VDD1.n58 VDD1.n22 0.388379
R2220 VDD1.n57 VDD1.n56 0.388379
R2221 VDD1.n162 VDD1.n161 0.388379
R2222 VDD1.n163 VDD1.n127 0.388379
R2223 VDD1.n103 VDD1.n1 0.155672
R2224 VDD1.n96 VDD1.n1 0.155672
R2225 VDD1.n96 VDD1.n95 0.155672
R2226 VDD1.n95 VDD1.n5 0.155672
R2227 VDD1.n88 VDD1.n5 0.155672
R2228 VDD1.n88 VDD1.n87 0.155672
R2229 VDD1.n87 VDD1.n9 0.155672
R2230 VDD1.n80 VDD1.n9 0.155672
R2231 VDD1.n80 VDD1.n79 0.155672
R2232 VDD1.n79 VDD1.n13 0.155672
R2233 VDD1.n72 VDD1.n13 0.155672
R2234 VDD1.n72 VDD1.n71 0.155672
R2235 VDD1.n71 VDD1.n17 0.155672
R2236 VDD1.n64 VDD1.n17 0.155672
R2237 VDD1.n64 VDD1.n63 0.155672
R2238 VDD1.n63 VDD1.n21 0.155672
R2239 VDD1.n55 VDD1.n21 0.155672
R2240 VDD1.n55 VDD1.n54 0.155672
R2241 VDD1.n54 VDD1.n25 0.155672
R2242 VDD1.n47 VDD1.n25 0.155672
R2243 VDD1.n47 VDD1.n46 0.155672
R2244 VDD1.n46 VDD1.n30 0.155672
R2245 VDD1.n39 VDD1.n30 0.155672
R2246 VDD1.n39 VDD1.n38 0.155672
R2247 VDD1.n143 VDD1.n142 0.155672
R2248 VDD1.n143 VDD1.n134 0.155672
R2249 VDD1.n150 VDD1.n134 0.155672
R2250 VDD1.n151 VDD1.n150 0.155672
R2251 VDD1.n151 VDD1.n130 0.155672
R2252 VDD1.n159 VDD1.n130 0.155672
R2253 VDD1.n160 VDD1.n159 0.155672
R2254 VDD1.n160 VDD1.n126 0.155672
R2255 VDD1.n168 VDD1.n126 0.155672
R2256 VDD1.n169 VDD1.n168 0.155672
R2257 VDD1.n169 VDD1.n122 0.155672
R2258 VDD1.n176 VDD1.n122 0.155672
R2259 VDD1.n177 VDD1.n176 0.155672
R2260 VDD1.n177 VDD1.n118 0.155672
R2261 VDD1.n184 VDD1.n118 0.155672
R2262 VDD1.n185 VDD1.n184 0.155672
R2263 VDD1.n185 VDD1.n114 0.155672
R2264 VDD1.n192 VDD1.n114 0.155672
R2265 VDD1.n193 VDD1.n192 0.155672
R2266 VDD1.n193 VDD1.n110 0.155672
R2267 VDD1.n200 VDD1.n110 0.155672
R2268 VDD1.n201 VDD1.n200 0.155672
R2269 VDD1.n201 VDD1.n106 0.155672
R2270 VDD1.n208 VDD1.n106 0.155672
C0 VP w_n1206_n4884# 1.78978f
C1 VP VN 5.76475f
C2 VP VDD1 2.18068f
C3 VP VDD2 0.238484f
C4 B w_n1206_n4884# 8.432321f
C5 VP VTAIL 1.15704f
C6 B VN 0.741617f
C7 B VDD1 1.85966f
C8 B VDD2 1.87134f
C9 VN w_n1206_n4884# 1.6412f
C10 B VTAIL 3.68923f
C11 VDD1 w_n1206_n4884# 2.09612f
C12 VN VDD1 0.148711f
C13 VDD2 w_n1206_n4884# 2.09644f
C14 VTAIL w_n1206_n4884# 4.34893f
C15 VN VDD2 2.09921f
C16 VDD1 VDD2 0.426016f
C17 VN VTAIL 1.14184f
C18 VTAIL VDD1 11.090199f
C19 B VP 0.976494f
C20 VTAIL VDD2 11.1135f
C21 VDD2 VSUBS 0.988413f
C22 VDD1 VSUBS 4.99871f
C23 VTAIL VSUBS 0.216309f
C24 VN VSUBS 7.79426f
C25 VP VSUBS 1.269279f
C26 B VSUBS 2.814605f
C27 w_n1206_n4884# VSUBS 71.9403f
C28 VDD1.n0 VSUBS 0.031292f
C29 VDD1.n1 VSUBS 0.027865f
C30 VDD1.n2 VSUBS 0.014974f
C31 VDD1.n3 VSUBS 0.035392f
C32 VDD1.n4 VSUBS 0.015854f
C33 VDD1.n5 VSUBS 0.027865f
C34 VDD1.n6 VSUBS 0.014974f
C35 VDD1.n7 VSUBS 0.035392f
C36 VDD1.n8 VSUBS 0.015854f
C37 VDD1.n9 VSUBS 0.027865f
C38 VDD1.n10 VSUBS 0.014974f
C39 VDD1.n11 VSUBS 0.035392f
C40 VDD1.n12 VSUBS 0.015854f
C41 VDD1.n13 VSUBS 0.027865f
C42 VDD1.n14 VSUBS 0.014974f
C43 VDD1.n15 VSUBS 0.035392f
C44 VDD1.n16 VSUBS 0.015854f
C45 VDD1.n17 VSUBS 0.027865f
C46 VDD1.n18 VSUBS 0.014974f
C47 VDD1.n19 VSUBS 0.035392f
C48 VDD1.n20 VSUBS 0.015854f
C49 VDD1.n21 VSUBS 0.027865f
C50 VDD1.n22 VSUBS 0.014974f
C51 VDD1.n23 VSUBS 0.035392f
C52 VDD1.n24 VSUBS 0.015854f
C53 VDD1.n25 VSUBS 0.027865f
C54 VDD1.n26 VSUBS 0.014974f
C55 VDD1.n27 VSUBS 0.035392f
C56 VDD1.n28 VSUBS 0.035392f
C57 VDD1.n29 VSUBS 0.015854f
C58 VDD1.n30 VSUBS 0.027865f
C59 VDD1.n31 VSUBS 0.014974f
C60 VDD1.n32 VSUBS 0.035392f
C61 VDD1.n33 VSUBS 0.015854f
C62 VDD1.n34 VSUBS 0.314705f
C63 VDD1.t1 VSUBS 0.076977f
C64 VDD1.n35 VSUBS 0.026544f
C65 VDD1.n36 VSUBS 0.026624f
C66 VDD1.n37 VSUBS 0.014974f
C67 VDD1.n38 VSUBS 2.29213f
C68 VDD1.n39 VSUBS 0.027865f
C69 VDD1.n40 VSUBS 0.014974f
C70 VDD1.n41 VSUBS 0.015854f
C71 VDD1.n42 VSUBS 0.035392f
C72 VDD1.n43 VSUBS 0.035392f
C73 VDD1.n44 VSUBS 0.015854f
C74 VDD1.n45 VSUBS 0.014974f
C75 VDD1.n46 VSUBS 0.027865f
C76 VDD1.n47 VSUBS 0.027865f
C77 VDD1.n48 VSUBS 0.014974f
C78 VDD1.n49 VSUBS 0.015854f
C79 VDD1.n50 VSUBS 0.035392f
C80 VDD1.n51 VSUBS 0.035392f
C81 VDD1.n52 VSUBS 0.015854f
C82 VDD1.n53 VSUBS 0.014974f
C83 VDD1.n54 VSUBS 0.027865f
C84 VDD1.n55 VSUBS 0.027865f
C85 VDD1.n56 VSUBS 0.014974f
C86 VDD1.n57 VSUBS 0.015414f
C87 VDD1.n58 VSUBS 0.015414f
C88 VDD1.n59 VSUBS 0.035392f
C89 VDD1.n60 VSUBS 0.035392f
C90 VDD1.n61 VSUBS 0.015854f
C91 VDD1.n62 VSUBS 0.014974f
C92 VDD1.n63 VSUBS 0.027865f
C93 VDD1.n64 VSUBS 0.027865f
C94 VDD1.n65 VSUBS 0.014974f
C95 VDD1.n66 VSUBS 0.015854f
C96 VDD1.n67 VSUBS 0.035392f
C97 VDD1.n68 VSUBS 0.035392f
C98 VDD1.n69 VSUBS 0.015854f
C99 VDD1.n70 VSUBS 0.014974f
C100 VDD1.n71 VSUBS 0.027865f
C101 VDD1.n72 VSUBS 0.027865f
C102 VDD1.n73 VSUBS 0.014974f
C103 VDD1.n74 VSUBS 0.015854f
C104 VDD1.n75 VSUBS 0.035392f
C105 VDD1.n76 VSUBS 0.035392f
C106 VDD1.n77 VSUBS 0.015854f
C107 VDD1.n78 VSUBS 0.014974f
C108 VDD1.n79 VSUBS 0.027865f
C109 VDD1.n80 VSUBS 0.027865f
C110 VDD1.n81 VSUBS 0.014974f
C111 VDD1.n82 VSUBS 0.015854f
C112 VDD1.n83 VSUBS 0.035392f
C113 VDD1.n84 VSUBS 0.035392f
C114 VDD1.n85 VSUBS 0.015854f
C115 VDD1.n86 VSUBS 0.014974f
C116 VDD1.n87 VSUBS 0.027865f
C117 VDD1.n88 VSUBS 0.027865f
C118 VDD1.n89 VSUBS 0.014974f
C119 VDD1.n90 VSUBS 0.015854f
C120 VDD1.n91 VSUBS 0.035392f
C121 VDD1.n92 VSUBS 0.035392f
C122 VDD1.n93 VSUBS 0.015854f
C123 VDD1.n94 VSUBS 0.014974f
C124 VDD1.n95 VSUBS 0.027865f
C125 VDD1.n96 VSUBS 0.027865f
C126 VDD1.n97 VSUBS 0.014974f
C127 VDD1.n98 VSUBS 0.015854f
C128 VDD1.n99 VSUBS 0.035392f
C129 VDD1.n100 VSUBS 0.090237f
C130 VDD1.n101 VSUBS 0.015854f
C131 VDD1.n102 VSUBS 0.029404f
C132 VDD1.n103 VSUBS 0.073545f
C133 VDD1.n104 VSUBS 0.089802f
C134 VDD1.n105 VSUBS 0.031292f
C135 VDD1.n106 VSUBS 0.027865f
C136 VDD1.n107 VSUBS 0.014974f
C137 VDD1.n108 VSUBS 0.035392f
C138 VDD1.n109 VSUBS 0.015854f
C139 VDD1.n110 VSUBS 0.027865f
C140 VDD1.n111 VSUBS 0.014974f
C141 VDD1.n112 VSUBS 0.035392f
C142 VDD1.n113 VSUBS 0.015854f
C143 VDD1.n114 VSUBS 0.027865f
C144 VDD1.n115 VSUBS 0.014974f
C145 VDD1.n116 VSUBS 0.035392f
C146 VDD1.n117 VSUBS 0.015854f
C147 VDD1.n118 VSUBS 0.027865f
C148 VDD1.n119 VSUBS 0.014974f
C149 VDD1.n120 VSUBS 0.035392f
C150 VDD1.n121 VSUBS 0.015854f
C151 VDD1.n122 VSUBS 0.027865f
C152 VDD1.n123 VSUBS 0.014974f
C153 VDD1.n124 VSUBS 0.035392f
C154 VDD1.n125 VSUBS 0.015854f
C155 VDD1.n126 VSUBS 0.027865f
C156 VDD1.n127 VSUBS 0.014974f
C157 VDD1.n128 VSUBS 0.035392f
C158 VDD1.n129 VSUBS 0.015854f
C159 VDD1.n130 VSUBS 0.027865f
C160 VDD1.n131 VSUBS 0.014974f
C161 VDD1.n132 VSUBS 0.035392f
C162 VDD1.n133 VSUBS 0.015854f
C163 VDD1.n134 VSUBS 0.027865f
C164 VDD1.n135 VSUBS 0.014974f
C165 VDD1.n136 VSUBS 0.035392f
C166 VDD1.n137 VSUBS 0.015854f
C167 VDD1.n138 VSUBS 0.314705f
C168 VDD1.t0 VSUBS 0.076977f
C169 VDD1.n139 VSUBS 0.026544f
C170 VDD1.n140 VSUBS 0.026624f
C171 VDD1.n141 VSUBS 0.014974f
C172 VDD1.n142 VSUBS 2.29213f
C173 VDD1.n143 VSUBS 0.027865f
C174 VDD1.n144 VSUBS 0.014974f
C175 VDD1.n145 VSUBS 0.015854f
C176 VDD1.n146 VSUBS 0.035392f
C177 VDD1.n147 VSUBS 0.035392f
C178 VDD1.n148 VSUBS 0.015854f
C179 VDD1.n149 VSUBS 0.014974f
C180 VDD1.n150 VSUBS 0.027865f
C181 VDD1.n151 VSUBS 0.027865f
C182 VDD1.n152 VSUBS 0.014974f
C183 VDD1.n153 VSUBS 0.015854f
C184 VDD1.n154 VSUBS 0.035392f
C185 VDD1.n155 VSUBS 0.035392f
C186 VDD1.n156 VSUBS 0.035392f
C187 VDD1.n157 VSUBS 0.015854f
C188 VDD1.n158 VSUBS 0.014974f
C189 VDD1.n159 VSUBS 0.027865f
C190 VDD1.n160 VSUBS 0.027865f
C191 VDD1.n161 VSUBS 0.014974f
C192 VDD1.n162 VSUBS 0.015414f
C193 VDD1.n163 VSUBS 0.015414f
C194 VDD1.n164 VSUBS 0.035392f
C195 VDD1.n165 VSUBS 0.035392f
C196 VDD1.n166 VSUBS 0.015854f
C197 VDD1.n167 VSUBS 0.014974f
C198 VDD1.n168 VSUBS 0.027865f
C199 VDD1.n169 VSUBS 0.027865f
C200 VDD1.n170 VSUBS 0.014974f
C201 VDD1.n171 VSUBS 0.015854f
C202 VDD1.n172 VSUBS 0.035392f
C203 VDD1.n173 VSUBS 0.035392f
C204 VDD1.n174 VSUBS 0.015854f
C205 VDD1.n175 VSUBS 0.014974f
C206 VDD1.n176 VSUBS 0.027865f
C207 VDD1.n177 VSUBS 0.027865f
C208 VDD1.n178 VSUBS 0.014974f
C209 VDD1.n179 VSUBS 0.015854f
C210 VDD1.n180 VSUBS 0.035392f
C211 VDD1.n181 VSUBS 0.035392f
C212 VDD1.n182 VSUBS 0.015854f
C213 VDD1.n183 VSUBS 0.014974f
C214 VDD1.n184 VSUBS 0.027865f
C215 VDD1.n185 VSUBS 0.027865f
C216 VDD1.n186 VSUBS 0.014974f
C217 VDD1.n187 VSUBS 0.015854f
C218 VDD1.n188 VSUBS 0.035392f
C219 VDD1.n189 VSUBS 0.035392f
C220 VDD1.n190 VSUBS 0.015854f
C221 VDD1.n191 VSUBS 0.014974f
C222 VDD1.n192 VSUBS 0.027865f
C223 VDD1.n193 VSUBS 0.027865f
C224 VDD1.n194 VSUBS 0.014974f
C225 VDD1.n195 VSUBS 0.015854f
C226 VDD1.n196 VSUBS 0.035392f
C227 VDD1.n197 VSUBS 0.035392f
C228 VDD1.n198 VSUBS 0.015854f
C229 VDD1.n199 VSUBS 0.014974f
C230 VDD1.n200 VSUBS 0.027865f
C231 VDD1.n201 VSUBS 0.027865f
C232 VDD1.n202 VSUBS 0.014974f
C233 VDD1.n203 VSUBS 0.015854f
C234 VDD1.n204 VSUBS 0.035392f
C235 VDD1.n205 VSUBS 0.090237f
C236 VDD1.n206 VSUBS 0.015854f
C237 VDD1.n207 VSUBS 0.029404f
C238 VDD1.n208 VSUBS 0.073545f
C239 VDD1.n209 VSUBS 0.97527f
C240 VP.t0 VSUBS 0.973604f
C241 VP.t1 VSUBS 0.911015f
C242 VP.n0 VSUBS 6.10798f
C243 VDD2.n0 VSUBS 0.031298f
C244 VDD2.n1 VSUBS 0.02787f
C245 VDD2.n2 VSUBS 0.014976f
C246 VDD2.n3 VSUBS 0.035399f
C247 VDD2.n4 VSUBS 0.015857f
C248 VDD2.n5 VSUBS 0.02787f
C249 VDD2.n6 VSUBS 0.014976f
C250 VDD2.n7 VSUBS 0.035399f
C251 VDD2.n8 VSUBS 0.015857f
C252 VDD2.n9 VSUBS 0.02787f
C253 VDD2.n10 VSUBS 0.014976f
C254 VDD2.n11 VSUBS 0.035399f
C255 VDD2.n12 VSUBS 0.015857f
C256 VDD2.n13 VSUBS 0.02787f
C257 VDD2.n14 VSUBS 0.014976f
C258 VDD2.n15 VSUBS 0.035399f
C259 VDD2.n16 VSUBS 0.015857f
C260 VDD2.n17 VSUBS 0.02787f
C261 VDD2.n18 VSUBS 0.014976f
C262 VDD2.n19 VSUBS 0.035399f
C263 VDD2.n20 VSUBS 0.015857f
C264 VDD2.n21 VSUBS 0.02787f
C265 VDD2.n22 VSUBS 0.014976f
C266 VDD2.n23 VSUBS 0.035399f
C267 VDD2.n24 VSUBS 0.015857f
C268 VDD2.n25 VSUBS 0.02787f
C269 VDD2.n26 VSUBS 0.014976f
C270 VDD2.n27 VSUBS 0.035399f
C271 VDD2.n28 VSUBS 0.015857f
C272 VDD2.n29 VSUBS 0.02787f
C273 VDD2.n30 VSUBS 0.014976f
C274 VDD2.n31 VSUBS 0.035399f
C275 VDD2.n32 VSUBS 0.015857f
C276 VDD2.n33 VSUBS 0.314765f
C277 VDD2.t1 VSUBS 0.076992f
C278 VDD2.n34 VSUBS 0.026549f
C279 VDD2.n35 VSUBS 0.026629f
C280 VDD2.n36 VSUBS 0.014976f
C281 VDD2.n37 VSUBS 2.29257f
C282 VDD2.n38 VSUBS 0.02787f
C283 VDD2.n39 VSUBS 0.014976f
C284 VDD2.n40 VSUBS 0.015857f
C285 VDD2.n41 VSUBS 0.035399f
C286 VDD2.n42 VSUBS 0.035399f
C287 VDD2.n43 VSUBS 0.015857f
C288 VDD2.n44 VSUBS 0.014976f
C289 VDD2.n45 VSUBS 0.02787f
C290 VDD2.n46 VSUBS 0.02787f
C291 VDD2.n47 VSUBS 0.014976f
C292 VDD2.n48 VSUBS 0.015857f
C293 VDD2.n49 VSUBS 0.035399f
C294 VDD2.n50 VSUBS 0.035399f
C295 VDD2.n51 VSUBS 0.035399f
C296 VDD2.n52 VSUBS 0.015857f
C297 VDD2.n53 VSUBS 0.014976f
C298 VDD2.n54 VSUBS 0.02787f
C299 VDD2.n55 VSUBS 0.02787f
C300 VDD2.n56 VSUBS 0.014976f
C301 VDD2.n57 VSUBS 0.015417f
C302 VDD2.n58 VSUBS 0.015417f
C303 VDD2.n59 VSUBS 0.035399f
C304 VDD2.n60 VSUBS 0.035399f
C305 VDD2.n61 VSUBS 0.015857f
C306 VDD2.n62 VSUBS 0.014976f
C307 VDD2.n63 VSUBS 0.02787f
C308 VDD2.n64 VSUBS 0.02787f
C309 VDD2.n65 VSUBS 0.014976f
C310 VDD2.n66 VSUBS 0.015857f
C311 VDD2.n67 VSUBS 0.035399f
C312 VDD2.n68 VSUBS 0.035399f
C313 VDD2.n69 VSUBS 0.015857f
C314 VDD2.n70 VSUBS 0.014976f
C315 VDD2.n71 VSUBS 0.02787f
C316 VDD2.n72 VSUBS 0.02787f
C317 VDD2.n73 VSUBS 0.014976f
C318 VDD2.n74 VSUBS 0.015857f
C319 VDD2.n75 VSUBS 0.035399f
C320 VDD2.n76 VSUBS 0.035399f
C321 VDD2.n77 VSUBS 0.015857f
C322 VDD2.n78 VSUBS 0.014976f
C323 VDD2.n79 VSUBS 0.02787f
C324 VDD2.n80 VSUBS 0.02787f
C325 VDD2.n81 VSUBS 0.014976f
C326 VDD2.n82 VSUBS 0.015857f
C327 VDD2.n83 VSUBS 0.035399f
C328 VDD2.n84 VSUBS 0.035399f
C329 VDD2.n85 VSUBS 0.015857f
C330 VDD2.n86 VSUBS 0.014976f
C331 VDD2.n87 VSUBS 0.02787f
C332 VDD2.n88 VSUBS 0.02787f
C333 VDD2.n89 VSUBS 0.014976f
C334 VDD2.n90 VSUBS 0.015857f
C335 VDD2.n91 VSUBS 0.035399f
C336 VDD2.n92 VSUBS 0.035399f
C337 VDD2.n93 VSUBS 0.015857f
C338 VDD2.n94 VSUBS 0.014976f
C339 VDD2.n95 VSUBS 0.02787f
C340 VDD2.n96 VSUBS 0.02787f
C341 VDD2.n97 VSUBS 0.014976f
C342 VDD2.n98 VSUBS 0.015857f
C343 VDD2.n99 VSUBS 0.035399f
C344 VDD2.n100 VSUBS 0.090254f
C345 VDD2.n101 VSUBS 0.015857f
C346 VDD2.n102 VSUBS 0.02941f
C347 VDD2.n103 VSUBS 0.073559f
C348 VDD2.n104 VSUBS 0.939767f
C349 VDD2.n105 VSUBS 0.031298f
C350 VDD2.n106 VSUBS 0.02787f
C351 VDD2.n107 VSUBS 0.014976f
C352 VDD2.n108 VSUBS 0.035399f
C353 VDD2.n109 VSUBS 0.015857f
C354 VDD2.n110 VSUBS 0.02787f
C355 VDD2.n111 VSUBS 0.014976f
C356 VDD2.n112 VSUBS 0.035399f
C357 VDD2.n113 VSUBS 0.015857f
C358 VDD2.n114 VSUBS 0.02787f
C359 VDD2.n115 VSUBS 0.014976f
C360 VDD2.n116 VSUBS 0.035399f
C361 VDD2.n117 VSUBS 0.015857f
C362 VDD2.n118 VSUBS 0.02787f
C363 VDD2.n119 VSUBS 0.014976f
C364 VDD2.n120 VSUBS 0.035399f
C365 VDD2.n121 VSUBS 0.015857f
C366 VDD2.n122 VSUBS 0.02787f
C367 VDD2.n123 VSUBS 0.014976f
C368 VDD2.n124 VSUBS 0.035399f
C369 VDD2.n125 VSUBS 0.015857f
C370 VDD2.n126 VSUBS 0.02787f
C371 VDD2.n127 VSUBS 0.014976f
C372 VDD2.n128 VSUBS 0.035399f
C373 VDD2.n129 VSUBS 0.015857f
C374 VDD2.n130 VSUBS 0.02787f
C375 VDD2.n131 VSUBS 0.014976f
C376 VDD2.n132 VSUBS 0.035399f
C377 VDD2.n133 VSUBS 0.035399f
C378 VDD2.n134 VSUBS 0.015857f
C379 VDD2.n135 VSUBS 0.02787f
C380 VDD2.n136 VSUBS 0.014976f
C381 VDD2.n137 VSUBS 0.035399f
C382 VDD2.n138 VSUBS 0.015857f
C383 VDD2.n139 VSUBS 0.314765f
C384 VDD2.t0 VSUBS 0.076992f
C385 VDD2.n140 VSUBS 0.026549f
C386 VDD2.n141 VSUBS 0.026629f
C387 VDD2.n142 VSUBS 0.014976f
C388 VDD2.n143 VSUBS 2.29257f
C389 VDD2.n144 VSUBS 0.02787f
C390 VDD2.n145 VSUBS 0.014976f
C391 VDD2.n146 VSUBS 0.015857f
C392 VDD2.n147 VSUBS 0.035399f
C393 VDD2.n148 VSUBS 0.035399f
C394 VDD2.n149 VSUBS 0.015857f
C395 VDD2.n150 VSUBS 0.014976f
C396 VDD2.n151 VSUBS 0.02787f
C397 VDD2.n152 VSUBS 0.02787f
C398 VDD2.n153 VSUBS 0.014976f
C399 VDD2.n154 VSUBS 0.015857f
C400 VDD2.n155 VSUBS 0.035399f
C401 VDD2.n156 VSUBS 0.035399f
C402 VDD2.n157 VSUBS 0.015857f
C403 VDD2.n158 VSUBS 0.014976f
C404 VDD2.n159 VSUBS 0.02787f
C405 VDD2.n160 VSUBS 0.02787f
C406 VDD2.n161 VSUBS 0.014976f
C407 VDD2.n162 VSUBS 0.015417f
C408 VDD2.n163 VSUBS 0.015417f
C409 VDD2.n164 VSUBS 0.035399f
C410 VDD2.n165 VSUBS 0.035399f
C411 VDD2.n166 VSUBS 0.015857f
C412 VDD2.n167 VSUBS 0.014976f
C413 VDD2.n168 VSUBS 0.02787f
C414 VDD2.n169 VSUBS 0.02787f
C415 VDD2.n170 VSUBS 0.014976f
C416 VDD2.n171 VSUBS 0.015857f
C417 VDD2.n172 VSUBS 0.035399f
C418 VDD2.n173 VSUBS 0.035399f
C419 VDD2.n174 VSUBS 0.015857f
C420 VDD2.n175 VSUBS 0.014976f
C421 VDD2.n176 VSUBS 0.02787f
C422 VDD2.n177 VSUBS 0.02787f
C423 VDD2.n178 VSUBS 0.014976f
C424 VDD2.n179 VSUBS 0.015857f
C425 VDD2.n180 VSUBS 0.035399f
C426 VDD2.n181 VSUBS 0.035399f
C427 VDD2.n182 VSUBS 0.015857f
C428 VDD2.n183 VSUBS 0.014976f
C429 VDD2.n184 VSUBS 0.02787f
C430 VDD2.n185 VSUBS 0.02787f
C431 VDD2.n186 VSUBS 0.014976f
C432 VDD2.n187 VSUBS 0.015857f
C433 VDD2.n188 VSUBS 0.035399f
C434 VDD2.n189 VSUBS 0.035399f
C435 VDD2.n190 VSUBS 0.015857f
C436 VDD2.n191 VSUBS 0.014976f
C437 VDD2.n192 VSUBS 0.02787f
C438 VDD2.n193 VSUBS 0.02787f
C439 VDD2.n194 VSUBS 0.014976f
C440 VDD2.n195 VSUBS 0.015857f
C441 VDD2.n196 VSUBS 0.035399f
C442 VDD2.n197 VSUBS 0.035399f
C443 VDD2.n198 VSUBS 0.015857f
C444 VDD2.n199 VSUBS 0.014976f
C445 VDD2.n200 VSUBS 0.02787f
C446 VDD2.n201 VSUBS 0.02787f
C447 VDD2.n202 VSUBS 0.014976f
C448 VDD2.n203 VSUBS 0.015857f
C449 VDD2.n204 VSUBS 0.035399f
C450 VDD2.n205 VSUBS 0.090254f
C451 VDD2.n206 VSUBS 0.015857f
C452 VDD2.n207 VSUBS 0.02941f
C453 VDD2.n208 VSUBS 0.073559f
C454 VDD2.n209 VSUBS 0.089558f
C455 VDD2.n210 VSUBS 3.81523f
C456 VTAIL.n0 VSUBS 0.032216f
C457 VTAIL.n1 VSUBS 0.028688f
C458 VTAIL.n2 VSUBS 0.015415f
C459 VTAIL.n3 VSUBS 0.036437f
C460 VTAIL.n4 VSUBS 0.016322f
C461 VTAIL.n5 VSUBS 0.028688f
C462 VTAIL.n6 VSUBS 0.015415f
C463 VTAIL.n7 VSUBS 0.036437f
C464 VTAIL.n8 VSUBS 0.016322f
C465 VTAIL.n9 VSUBS 0.028688f
C466 VTAIL.n10 VSUBS 0.015415f
C467 VTAIL.n11 VSUBS 0.036437f
C468 VTAIL.n12 VSUBS 0.016322f
C469 VTAIL.n13 VSUBS 0.028688f
C470 VTAIL.n14 VSUBS 0.015415f
C471 VTAIL.n15 VSUBS 0.036437f
C472 VTAIL.n16 VSUBS 0.016322f
C473 VTAIL.n17 VSUBS 0.028688f
C474 VTAIL.n18 VSUBS 0.015415f
C475 VTAIL.n19 VSUBS 0.036437f
C476 VTAIL.n20 VSUBS 0.016322f
C477 VTAIL.n21 VSUBS 0.028688f
C478 VTAIL.n22 VSUBS 0.015415f
C479 VTAIL.n23 VSUBS 0.036437f
C480 VTAIL.n24 VSUBS 0.016322f
C481 VTAIL.n25 VSUBS 0.028688f
C482 VTAIL.n26 VSUBS 0.015415f
C483 VTAIL.n27 VSUBS 0.036437f
C484 VTAIL.n28 VSUBS 0.016322f
C485 VTAIL.n29 VSUBS 0.028688f
C486 VTAIL.n30 VSUBS 0.015415f
C487 VTAIL.n31 VSUBS 0.036437f
C488 VTAIL.n32 VSUBS 0.016322f
C489 VTAIL.n33 VSUBS 0.323995f
C490 VTAIL.t1 VSUBS 0.07925f
C491 VTAIL.n34 VSUBS 0.027327f
C492 VTAIL.n35 VSUBS 0.02741f
C493 VTAIL.n36 VSUBS 0.015415f
C494 VTAIL.n37 VSUBS 2.3598f
C495 VTAIL.n38 VSUBS 0.028688f
C496 VTAIL.n39 VSUBS 0.015415f
C497 VTAIL.n40 VSUBS 0.016322f
C498 VTAIL.n41 VSUBS 0.036437f
C499 VTAIL.n42 VSUBS 0.036437f
C500 VTAIL.n43 VSUBS 0.016322f
C501 VTAIL.n44 VSUBS 0.015415f
C502 VTAIL.n45 VSUBS 0.028688f
C503 VTAIL.n46 VSUBS 0.028688f
C504 VTAIL.n47 VSUBS 0.015415f
C505 VTAIL.n48 VSUBS 0.016322f
C506 VTAIL.n49 VSUBS 0.036437f
C507 VTAIL.n50 VSUBS 0.036437f
C508 VTAIL.n51 VSUBS 0.036437f
C509 VTAIL.n52 VSUBS 0.016322f
C510 VTAIL.n53 VSUBS 0.015415f
C511 VTAIL.n54 VSUBS 0.028688f
C512 VTAIL.n55 VSUBS 0.028688f
C513 VTAIL.n56 VSUBS 0.015415f
C514 VTAIL.n57 VSUBS 0.015869f
C515 VTAIL.n58 VSUBS 0.015869f
C516 VTAIL.n59 VSUBS 0.036437f
C517 VTAIL.n60 VSUBS 0.036437f
C518 VTAIL.n61 VSUBS 0.016322f
C519 VTAIL.n62 VSUBS 0.015415f
C520 VTAIL.n63 VSUBS 0.028688f
C521 VTAIL.n64 VSUBS 0.028688f
C522 VTAIL.n65 VSUBS 0.015415f
C523 VTAIL.n66 VSUBS 0.016322f
C524 VTAIL.n67 VSUBS 0.036437f
C525 VTAIL.n68 VSUBS 0.036437f
C526 VTAIL.n69 VSUBS 0.016322f
C527 VTAIL.n70 VSUBS 0.015415f
C528 VTAIL.n71 VSUBS 0.028688f
C529 VTAIL.n72 VSUBS 0.028688f
C530 VTAIL.n73 VSUBS 0.015415f
C531 VTAIL.n74 VSUBS 0.016322f
C532 VTAIL.n75 VSUBS 0.036437f
C533 VTAIL.n76 VSUBS 0.036437f
C534 VTAIL.n77 VSUBS 0.016322f
C535 VTAIL.n78 VSUBS 0.015415f
C536 VTAIL.n79 VSUBS 0.028688f
C537 VTAIL.n80 VSUBS 0.028688f
C538 VTAIL.n81 VSUBS 0.015415f
C539 VTAIL.n82 VSUBS 0.016322f
C540 VTAIL.n83 VSUBS 0.036437f
C541 VTAIL.n84 VSUBS 0.036437f
C542 VTAIL.n85 VSUBS 0.016322f
C543 VTAIL.n86 VSUBS 0.015415f
C544 VTAIL.n87 VSUBS 0.028688f
C545 VTAIL.n88 VSUBS 0.028688f
C546 VTAIL.n89 VSUBS 0.015415f
C547 VTAIL.n90 VSUBS 0.016322f
C548 VTAIL.n91 VSUBS 0.036437f
C549 VTAIL.n92 VSUBS 0.036437f
C550 VTAIL.n93 VSUBS 0.016322f
C551 VTAIL.n94 VSUBS 0.015415f
C552 VTAIL.n95 VSUBS 0.028688f
C553 VTAIL.n96 VSUBS 0.028688f
C554 VTAIL.n97 VSUBS 0.015415f
C555 VTAIL.n98 VSUBS 0.016322f
C556 VTAIL.n99 VSUBS 0.036437f
C557 VTAIL.n100 VSUBS 0.0929f
C558 VTAIL.n101 VSUBS 0.016322f
C559 VTAIL.n102 VSUBS 0.030272f
C560 VTAIL.n103 VSUBS 0.075716f
C561 VTAIL.n104 VSUBS 0.07244f
C562 VTAIL.n105 VSUBS 2.1344f
C563 VTAIL.n106 VSUBS 0.032216f
C564 VTAIL.n107 VSUBS 0.028688f
C565 VTAIL.n108 VSUBS 0.015415f
C566 VTAIL.n109 VSUBS 0.036437f
C567 VTAIL.n110 VSUBS 0.016322f
C568 VTAIL.n111 VSUBS 0.028688f
C569 VTAIL.n112 VSUBS 0.015415f
C570 VTAIL.n113 VSUBS 0.036437f
C571 VTAIL.n114 VSUBS 0.016322f
C572 VTAIL.n115 VSUBS 0.028688f
C573 VTAIL.n116 VSUBS 0.015415f
C574 VTAIL.n117 VSUBS 0.036437f
C575 VTAIL.n118 VSUBS 0.016322f
C576 VTAIL.n119 VSUBS 0.028688f
C577 VTAIL.n120 VSUBS 0.015415f
C578 VTAIL.n121 VSUBS 0.036437f
C579 VTAIL.n122 VSUBS 0.016322f
C580 VTAIL.n123 VSUBS 0.028688f
C581 VTAIL.n124 VSUBS 0.015415f
C582 VTAIL.n125 VSUBS 0.036437f
C583 VTAIL.n126 VSUBS 0.016322f
C584 VTAIL.n127 VSUBS 0.028688f
C585 VTAIL.n128 VSUBS 0.015415f
C586 VTAIL.n129 VSUBS 0.036437f
C587 VTAIL.n130 VSUBS 0.016322f
C588 VTAIL.n131 VSUBS 0.028688f
C589 VTAIL.n132 VSUBS 0.015415f
C590 VTAIL.n133 VSUBS 0.036437f
C591 VTAIL.n134 VSUBS 0.036437f
C592 VTAIL.n135 VSUBS 0.016322f
C593 VTAIL.n136 VSUBS 0.028688f
C594 VTAIL.n137 VSUBS 0.015415f
C595 VTAIL.n138 VSUBS 0.036437f
C596 VTAIL.n139 VSUBS 0.016322f
C597 VTAIL.n140 VSUBS 0.323995f
C598 VTAIL.t3 VSUBS 0.07925f
C599 VTAIL.n141 VSUBS 0.027327f
C600 VTAIL.n142 VSUBS 0.02741f
C601 VTAIL.n143 VSUBS 0.015415f
C602 VTAIL.n144 VSUBS 2.3598f
C603 VTAIL.n145 VSUBS 0.028688f
C604 VTAIL.n146 VSUBS 0.015415f
C605 VTAIL.n147 VSUBS 0.016322f
C606 VTAIL.n148 VSUBS 0.036437f
C607 VTAIL.n149 VSUBS 0.036437f
C608 VTAIL.n150 VSUBS 0.016322f
C609 VTAIL.n151 VSUBS 0.015415f
C610 VTAIL.n152 VSUBS 0.028688f
C611 VTAIL.n153 VSUBS 0.028688f
C612 VTAIL.n154 VSUBS 0.015415f
C613 VTAIL.n155 VSUBS 0.016322f
C614 VTAIL.n156 VSUBS 0.036437f
C615 VTAIL.n157 VSUBS 0.036437f
C616 VTAIL.n158 VSUBS 0.016322f
C617 VTAIL.n159 VSUBS 0.015415f
C618 VTAIL.n160 VSUBS 0.028688f
C619 VTAIL.n161 VSUBS 0.028688f
C620 VTAIL.n162 VSUBS 0.015415f
C621 VTAIL.n163 VSUBS 0.015869f
C622 VTAIL.n164 VSUBS 0.015869f
C623 VTAIL.n165 VSUBS 0.036437f
C624 VTAIL.n166 VSUBS 0.036437f
C625 VTAIL.n167 VSUBS 0.016322f
C626 VTAIL.n168 VSUBS 0.015415f
C627 VTAIL.n169 VSUBS 0.028688f
C628 VTAIL.n170 VSUBS 0.028688f
C629 VTAIL.n171 VSUBS 0.015415f
C630 VTAIL.n172 VSUBS 0.016322f
C631 VTAIL.n173 VSUBS 0.036437f
C632 VTAIL.n174 VSUBS 0.036437f
C633 VTAIL.n175 VSUBS 0.016322f
C634 VTAIL.n176 VSUBS 0.015415f
C635 VTAIL.n177 VSUBS 0.028688f
C636 VTAIL.n178 VSUBS 0.028688f
C637 VTAIL.n179 VSUBS 0.015415f
C638 VTAIL.n180 VSUBS 0.016322f
C639 VTAIL.n181 VSUBS 0.036437f
C640 VTAIL.n182 VSUBS 0.036437f
C641 VTAIL.n183 VSUBS 0.016322f
C642 VTAIL.n184 VSUBS 0.015415f
C643 VTAIL.n185 VSUBS 0.028688f
C644 VTAIL.n186 VSUBS 0.028688f
C645 VTAIL.n187 VSUBS 0.015415f
C646 VTAIL.n188 VSUBS 0.016322f
C647 VTAIL.n189 VSUBS 0.036437f
C648 VTAIL.n190 VSUBS 0.036437f
C649 VTAIL.n191 VSUBS 0.016322f
C650 VTAIL.n192 VSUBS 0.015415f
C651 VTAIL.n193 VSUBS 0.028688f
C652 VTAIL.n194 VSUBS 0.028688f
C653 VTAIL.n195 VSUBS 0.015415f
C654 VTAIL.n196 VSUBS 0.016322f
C655 VTAIL.n197 VSUBS 0.036437f
C656 VTAIL.n198 VSUBS 0.036437f
C657 VTAIL.n199 VSUBS 0.016322f
C658 VTAIL.n200 VSUBS 0.015415f
C659 VTAIL.n201 VSUBS 0.028688f
C660 VTAIL.n202 VSUBS 0.028688f
C661 VTAIL.n203 VSUBS 0.015415f
C662 VTAIL.n204 VSUBS 0.016322f
C663 VTAIL.n205 VSUBS 0.036437f
C664 VTAIL.n206 VSUBS 0.0929f
C665 VTAIL.n207 VSUBS 0.016322f
C666 VTAIL.n208 VSUBS 0.030272f
C667 VTAIL.n209 VSUBS 0.075716f
C668 VTAIL.n210 VSUBS 0.07244f
C669 VTAIL.n211 VSUBS 2.14077f
C670 VTAIL.n212 VSUBS 0.032216f
C671 VTAIL.n213 VSUBS 0.028688f
C672 VTAIL.n214 VSUBS 0.015415f
C673 VTAIL.n215 VSUBS 0.036437f
C674 VTAIL.n216 VSUBS 0.016322f
C675 VTAIL.n217 VSUBS 0.028688f
C676 VTAIL.n218 VSUBS 0.015415f
C677 VTAIL.n219 VSUBS 0.036437f
C678 VTAIL.n220 VSUBS 0.016322f
C679 VTAIL.n221 VSUBS 0.028688f
C680 VTAIL.n222 VSUBS 0.015415f
C681 VTAIL.n223 VSUBS 0.036437f
C682 VTAIL.n224 VSUBS 0.016322f
C683 VTAIL.n225 VSUBS 0.028688f
C684 VTAIL.n226 VSUBS 0.015415f
C685 VTAIL.n227 VSUBS 0.036437f
C686 VTAIL.n228 VSUBS 0.016322f
C687 VTAIL.n229 VSUBS 0.028688f
C688 VTAIL.n230 VSUBS 0.015415f
C689 VTAIL.n231 VSUBS 0.036437f
C690 VTAIL.n232 VSUBS 0.016322f
C691 VTAIL.n233 VSUBS 0.028688f
C692 VTAIL.n234 VSUBS 0.015415f
C693 VTAIL.n235 VSUBS 0.036437f
C694 VTAIL.n236 VSUBS 0.016322f
C695 VTAIL.n237 VSUBS 0.028688f
C696 VTAIL.n238 VSUBS 0.015415f
C697 VTAIL.n239 VSUBS 0.036437f
C698 VTAIL.n240 VSUBS 0.036437f
C699 VTAIL.n241 VSUBS 0.016322f
C700 VTAIL.n242 VSUBS 0.028688f
C701 VTAIL.n243 VSUBS 0.015415f
C702 VTAIL.n244 VSUBS 0.036437f
C703 VTAIL.n245 VSUBS 0.016322f
C704 VTAIL.n246 VSUBS 0.323995f
C705 VTAIL.t0 VSUBS 0.07925f
C706 VTAIL.n247 VSUBS 0.027327f
C707 VTAIL.n248 VSUBS 0.02741f
C708 VTAIL.n249 VSUBS 0.015415f
C709 VTAIL.n250 VSUBS 2.3598f
C710 VTAIL.n251 VSUBS 0.028688f
C711 VTAIL.n252 VSUBS 0.015415f
C712 VTAIL.n253 VSUBS 0.016322f
C713 VTAIL.n254 VSUBS 0.036437f
C714 VTAIL.n255 VSUBS 0.036437f
C715 VTAIL.n256 VSUBS 0.016322f
C716 VTAIL.n257 VSUBS 0.015415f
C717 VTAIL.n258 VSUBS 0.028688f
C718 VTAIL.n259 VSUBS 0.028688f
C719 VTAIL.n260 VSUBS 0.015415f
C720 VTAIL.n261 VSUBS 0.016322f
C721 VTAIL.n262 VSUBS 0.036437f
C722 VTAIL.n263 VSUBS 0.036437f
C723 VTAIL.n264 VSUBS 0.016322f
C724 VTAIL.n265 VSUBS 0.015415f
C725 VTAIL.n266 VSUBS 0.028688f
C726 VTAIL.n267 VSUBS 0.028688f
C727 VTAIL.n268 VSUBS 0.015415f
C728 VTAIL.n269 VSUBS 0.015869f
C729 VTAIL.n270 VSUBS 0.015869f
C730 VTAIL.n271 VSUBS 0.036437f
C731 VTAIL.n272 VSUBS 0.036437f
C732 VTAIL.n273 VSUBS 0.016322f
C733 VTAIL.n274 VSUBS 0.015415f
C734 VTAIL.n275 VSUBS 0.028688f
C735 VTAIL.n276 VSUBS 0.028688f
C736 VTAIL.n277 VSUBS 0.015415f
C737 VTAIL.n278 VSUBS 0.016322f
C738 VTAIL.n279 VSUBS 0.036437f
C739 VTAIL.n280 VSUBS 0.036437f
C740 VTAIL.n281 VSUBS 0.016322f
C741 VTAIL.n282 VSUBS 0.015415f
C742 VTAIL.n283 VSUBS 0.028688f
C743 VTAIL.n284 VSUBS 0.028688f
C744 VTAIL.n285 VSUBS 0.015415f
C745 VTAIL.n286 VSUBS 0.016322f
C746 VTAIL.n287 VSUBS 0.036437f
C747 VTAIL.n288 VSUBS 0.036437f
C748 VTAIL.n289 VSUBS 0.016322f
C749 VTAIL.n290 VSUBS 0.015415f
C750 VTAIL.n291 VSUBS 0.028688f
C751 VTAIL.n292 VSUBS 0.028688f
C752 VTAIL.n293 VSUBS 0.015415f
C753 VTAIL.n294 VSUBS 0.016322f
C754 VTAIL.n295 VSUBS 0.036437f
C755 VTAIL.n296 VSUBS 0.036437f
C756 VTAIL.n297 VSUBS 0.016322f
C757 VTAIL.n298 VSUBS 0.015415f
C758 VTAIL.n299 VSUBS 0.028688f
C759 VTAIL.n300 VSUBS 0.028688f
C760 VTAIL.n301 VSUBS 0.015415f
C761 VTAIL.n302 VSUBS 0.016322f
C762 VTAIL.n303 VSUBS 0.036437f
C763 VTAIL.n304 VSUBS 0.036437f
C764 VTAIL.n305 VSUBS 0.016322f
C765 VTAIL.n306 VSUBS 0.015415f
C766 VTAIL.n307 VSUBS 0.028688f
C767 VTAIL.n308 VSUBS 0.028688f
C768 VTAIL.n309 VSUBS 0.015415f
C769 VTAIL.n310 VSUBS 0.016322f
C770 VTAIL.n311 VSUBS 0.036437f
C771 VTAIL.n312 VSUBS 0.0929f
C772 VTAIL.n313 VSUBS 0.016322f
C773 VTAIL.n314 VSUBS 0.030272f
C774 VTAIL.n315 VSUBS 0.075716f
C775 VTAIL.n316 VSUBS 0.07244f
C776 VTAIL.n317 VSUBS 2.09376f
C777 VTAIL.n318 VSUBS 0.032216f
C778 VTAIL.n319 VSUBS 0.028688f
C779 VTAIL.n320 VSUBS 0.015415f
C780 VTAIL.n321 VSUBS 0.036437f
C781 VTAIL.n322 VSUBS 0.016322f
C782 VTAIL.n323 VSUBS 0.028688f
C783 VTAIL.n324 VSUBS 0.015415f
C784 VTAIL.n325 VSUBS 0.036437f
C785 VTAIL.n326 VSUBS 0.016322f
C786 VTAIL.n327 VSUBS 0.028688f
C787 VTAIL.n328 VSUBS 0.015415f
C788 VTAIL.n329 VSUBS 0.036437f
C789 VTAIL.n330 VSUBS 0.016322f
C790 VTAIL.n331 VSUBS 0.028688f
C791 VTAIL.n332 VSUBS 0.015415f
C792 VTAIL.n333 VSUBS 0.036437f
C793 VTAIL.n334 VSUBS 0.016322f
C794 VTAIL.n335 VSUBS 0.028688f
C795 VTAIL.n336 VSUBS 0.015415f
C796 VTAIL.n337 VSUBS 0.036437f
C797 VTAIL.n338 VSUBS 0.016322f
C798 VTAIL.n339 VSUBS 0.028688f
C799 VTAIL.n340 VSUBS 0.015415f
C800 VTAIL.n341 VSUBS 0.036437f
C801 VTAIL.n342 VSUBS 0.016322f
C802 VTAIL.n343 VSUBS 0.028688f
C803 VTAIL.n344 VSUBS 0.015415f
C804 VTAIL.n345 VSUBS 0.036437f
C805 VTAIL.n346 VSUBS 0.016322f
C806 VTAIL.n347 VSUBS 0.028688f
C807 VTAIL.n348 VSUBS 0.015415f
C808 VTAIL.n349 VSUBS 0.036437f
C809 VTAIL.n350 VSUBS 0.016322f
C810 VTAIL.n351 VSUBS 0.323995f
C811 VTAIL.t2 VSUBS 0.07925f
C812 VTAIL.n352 VSUBS 0.027327f
C813 VTAIL.n353 VSUBS 0.02741f
C814 VTAIL.n354 VSUBS 0.015415f
C815 VTAIL.n355 VSUBS 2.3598f
C816 VTAIL.n356 VSUBS 0.028688f
C817 VTAIL.n357 VSUBS 0.015415f
C818 VTAIL.n358 VSUBS 0.016322f
C819 VTAIL.n359 VSUBS 0.036437f
C820 VTAIL.n360 VSUBS 0.036437f
C821 VTAIL.n361 VSUBS 0.016322f
C822 VTAIL.n362 VSUBS 0.015415f
C823 VTAIL.n363 VSUBS 0.028688f
C824 VTAIL.n364 VSUBS 0.028688f
C825 VTAIL.n365 VSUBS 0.015415f
C826 VTAIL.n366 VSUBS 0.016322f
C827 VTAIL.n367 VSUBS 0.036437f
C828 VTAIL.n368 VSUBS 0.036437f
C829 VTAIL.n369 VSUBS 0.036437f
C830 VTAIL.n370 VSUBS 0.016322f
C831 VTAIL.n371 VSUBS 0.015415f
C832 VTAIL.n372 VSUBS 0.028688f
C833 VTAIL.n373 VSUBS 0.028688f
C834 VTAIL.n374 VSUBS 0.015415f
C835 VTAIL.n375 VSUBS 0.015869f
C836 VTAIL.n376 VSUBS 0.015869f
C837 VTAIL.n377 VSUBS 0.036437f
C838 VTAIL.n378 VSUBS 0.036437f
C839 VTAIL.n379 VSUBS 0.016322f
C840 VTAIL.n380 VSUBS 0.015415f
C841 VTAIL.n381 VSUBS 0.028688f
C842 VTAIL.n382 VSUBS 0.028688f
C843 VTAIL.n383 VSUBS 0.015415f
C844 VTAIL.n384 VSUBS 0.016322f
C845 VTAIL.n385 VSUBS 0.036437f
C846 VTAIL.n386 VSUBS 0.036437f
C847 VTAIL.n387 VSUBS 0.016322f
C848 VTAIL.n388 VSUBS 0.015415f
C849 VTAIL.n389 VSUBS 0.028688f
C850 VTAIL.n390 VSUBS 0.028688f
C851 VTAIL.n391 VSUBS 0.015415f
C852 VTAIL.n392 VSUBS 0.016322f
C853 VTAIL.n393 VSUBS 0.036437f
C854 VTAIL.n394 VSUBS 0.036437f
C855 VTAIL.n395 VSUBS 0.016322f
C856 VTAIL.n396 VSUBS 0.015415f
C857 VTAIL.n397 VSUBS 0.028688f
C858 VTAIL.n398 VSUBS 0.028688f
C859 VTAIL.n399 VSUBS 0.015415f
C860 VTAIL.n400 VSUBS 0.016322f
C861 VTAIL.n401 VSUBS 0.036437f
C862 VTAIL.n402 VSUBS 0.036437f
C863 VTAIL.n403 VSUBS 0.016322f
C864 VTAIL.n404 VSUBS 0.015415f
C865 VTAIL.n405 VSUBS 0.028688f
C866 VTAIL.n406 VSUBS 0.028688f
C867 VTAIL.n407 VSUBS 0.015415f
C868 VTAIL.n408 VSUBS 0.016322f
C869 VTAIL.n409 VSUBS 0.036437f
C870 VTAIL.n410 VSUBS 0.036437f
C871 VTAIL.n411 VSUBS 0.016322f
C872 VTAIL.n412 VSUBS 0.015415f
C873 VTAIL.n413 VSUBS 0.028688f
C874 VTAIL.n414 VSUBS 0.028688f
C875 VTAIL.n415 VSUBS 0.015415f
C876 VTAIL.n416 VSUBS 0.016322f
C877 VTAIL.n417 VSUBS 0.036437f
C878 VTAIL.n418 VSUBS 0.0929f
C879 VTAIL.n419 VSUBS 0.016322f
C880 VTAIL.n420 VSUBS 0.030272f
C881 VTAIL.n421 VSUBS 0.075716f
C882 VTAIL.n422 VSUBS 0.07244f
C883 VTAIL.n423 VSUBS 2.03319f
C884 VN.t0 VSUBS 0.890011f
C885 VN.t1 VSUBS 0.952475f
C886 B.n0 VSUBS 0.006459f
C887 B.n1 VSUBS 0.006459f
C888 B.n2 VSUBS 0.009552f
C889 B.n3 VSUBS 0.00732f
C890 B.n4 VSUBS 0.00732f
C891 B.n5 VSUBS 0.00732f
C892 B.n6 VSUBS 0.00732f
C893 B.n7 VSUBS 0.017783f
C894 B.n8 VSUBS 0.00732f
C895 B.n9 VSUBS 0.00732f
C896 B.n10 VSUBS 0.00732f
C897 B.n11 VSUBS 0.00732f
C898 B.n12 VSUBS 0.00732f
C899 B.n13 VSUBS 0.00732f
C900 B.n14 VSUBS 0.00732f
C901 B.n15 VSUBS 0.00732f
C902 B.n16 VSUBS 0.00732f
C903 B.n17 VSUBS 0.00732f
C904 B.n18 VSUBS 0.00732f
C905 B.n19 VSUBS 0.00732f
C906 B.n20 VSUBS 0.00732f
C907 B.n21 VSUBS 0.00732f
C908 B.n22 VSUBS 0.00732f
C909 B.n23 VSUBS 0.00732f
C910 B.n24 VSUBS 0.00732f
C911 B.n25 VSUBS 0.00732f
C912 B.n26 VSUBS 0.00732f
C913 B.n27 VSUBS 0.00732f
C914 B.n28 VSUBS 0.00732f
C915 B.n29 VSUBS 0.00732f
C916 B.n30 VSUBS 0.00732f
C917 B.n31 VSUBS 0.00732f
C918 B.n32 VSUBS 0.00732f
C919 B.n33 VSUBS 0.00732f
C920 B.n34 VSUBS 0.00732f
C921 B.n35 VSUBS 0.00732f
C922 B.n36 VSUBS 0.00732f
C923 B.n37 VSUBS 0.00732f
C924 B.n38 VSUBS 0.00732f
C925 B.n39 VSUBS 0.00732f
C926 B.t7 VSUBS 0.406849f
C927 B.t8 VSUBS 0.414337f
C928 B.t6 VSUBS 0.204946f
C929 B.n40 VSUBS 0.407858f
C930 B.n41 VSUBS 0.352855f
C931 B.n42 VSUBS 0.00732f
C932 B.n43 VSUBS 0.00732f
C933 B.n44 VSUBS 0.00732f
C934 B.n45 VSUBS 0.00732f
C935 B.t10 VSUBS 0.406853f
C936 B.t11 VSUBS 0.41434f
C937 B.t9 VSUBS 0.204946f
C938 B.n46 VSUBS 0.407854f
C939 B.n47 VSUBS 0.352851f
C940 B.n48 VSUBS 0.01696f
C941 B.n49 VSUBS 0.00732f
C942 B.n50 VSUBS 0.00732f
C943 B.n51 VSUBS 0.00732f
C944 B.n52 VSUBS 0.00732f
C945 B.n53 VSUBS 0.00732f
C946 B.n54 VSUBS 0.00732f
C947 B.n55 VSUBS 0.00732f
C948 B.n56 VSUBS 0.00732f
C949 B.n57 VSUBS 0.00732f
C950 B.n58 VSUBS 0.00732f
C951 B.n59 VSUBS 0.00732f
C952 B.n60 VSUBS 0.00732f
C953 B.n61 VSUBS 0.00732f
C954 B.n62 VSUBS 0.00732f
C955 B.n63 VSUBS 0.00732f
C956 B.n64 VSUBS 0.00732f
C957 B.n65 VSUBS 0.00732f
C958 B.n66 VSUBS 0.00732f
C959 B.n67 VSUBS 0.00732f
C960 B.n68 VSUBS 0.00732f
C961 B.n69 VSUBS 0.00732f
C962 B.n70 VSUBS 0.00732f
C963 B.n71 VSUBS 0.00732f
C964 B.n72 VSUBS 0.00732f
C965 B.n73 VSUBS 0.00732f
C966 B.n74 VSUBS 0.00732f
C967 B.n75 VSUBS 0.00732f
C968 B.n76 VSUBS 0.00732f
C969 B.n77 VSUBS 0.00732f
C970 B.n78 VSUBS 0.00732f
C971 B.n79 VSUBS 0.00732f
C972 B.n80 VSUBS 0.018386f
C973 B.n81 VSUBS 0.00732f
C974 B.n82 VSUBS 0.00732f
C975 B.n83 VSUBS 0.00732f
C976 B.n84 VSUBS 0.00732f
C977 B.n85 VSUBS 0.00732f
C978 B.n86 VSUBS 0.00732f
C979 B.n87 VSUBS 0.00732f
C980 B.n88 VSUBS 0.00732f
C981 B.n89 VSUBS 0.00732f
C982 B.n90 VSUBS 0.00732f
C983 B.n91 VSUBS 0.00732f
C984 B.n92 VSUBS 0.01858f
C985 B.n93 VSUBS 0.00732f
C986 B.n94 VSUBS 0.00732f
C987 B.n95 VSUBS 0.00732f
C988 B.n96 VSUBS 0.00732f
C989 B.n97 VSUBS 0.00732f
C990 B.n98 VSUBS 0.00732f
C991 B.n99 VSUBS 0.00732f
C992 B.n100 VSUBS 0.00732f
C993 B.n101 VSUBS 0.00732f
C994 B.n102 VSUBS 0.00732f
C995 B.n103 VSUBS 0.00732f
C996 B.n104 VSUBS 0.00732f
C997 B.n105 VSUBS 0.00732f
C998 B.n106 VSUBS 0.00732f
C999 B.n107 VSUBS 0.00732f
C1000 B.n108 VSUBS 0.00732f
C1001 B.n109 VSUBS 0.00732f
C1002 B.n110 VSUBS 0.00732f
C1003 B.n111 VSUBS 0.00732f
C1004 B.n112 VSUBS 0.00732f
C1005 B.n113 VSUBS 0.00732f
C1006 B.n114 VSUBS 0.00732f
C1007 B.n115 VSUBS 0.00732f
C1008 B.n116 VSUBS 0.00732f
C1009 B.n117 VSUBS 0.00732f
C1010 B.n118 VSUBS 0.00732f
C1011 B.n119 VSUBS 0.00732f
C1012 B.n120 VSUBS 0.00732f
C1013 B.n121 VSUBS 0.00732f
C1014 B.n122 VSUBS 0.00732f
C1015 B.n123 VSUBS 0.00732f
C1016 B.n124 VSUBS 0.004844f
C1017 B.n125 VSUBS 0.00732f
C1018 B.n126 VSUBS 0.00732f
C1019 B.n127 VSUBS 0.00732f
C1020 B.n128 VSUBS 0.00732f
C1021 B.n129 VSUBS 0.00732f
C1022 B.t5 VSUBS 0.406849f
C1023 B.t4 VSUBS 0.414337f
C1024 B.t3 VSUBS 0.204946f
C1025 B.n130 VSUBS 0.407858f
C1026 B.n131 VSUBS 0.352855f
C1027 B.n132 VSUBS 0.00732f
C1028 B.n133 VSUBS 0.00732f
C1029 B.n134 VSUBS 0.00732f
C1030 B.n135 VSUBS 0.00732f
C1031 B.n136 VSUBS 0.00732f
C1032 B.n137 VSUBS 0.00732f
C1033 B.n138 VSUBS 0.00732f
C1034 B.n139 VSUBS 0.00732f
C1035 B.n140 VSUBS 0.00732f
C1036 B.n141 VSUBS 0.00732f
C1037 B.n142 VSUBS 0.00732f
C1038 B.n143 VSUBS 0.00732f
C1039 B.n144 VSUBS 0.00732f
C1040 B.n145 VSUBS 0.00732f
C1041 B.n146 VSUBS 0.00732f
C1042 B.n147 VSUBS 0.00732f
C1043 B.n148 VSUBS 0.00732f
C1044 B.n149 VSUBS 0.00732f
C1045 B.n150 VSUBS 0.00732f
C1046 B.n151 VSUBS 0.00732f
C1047 B.n152 VSUBS 0.00732f
C1048 B.n153 VSUBS 0.00732f
C1049 B.n154 VSUBS 0.00732f
C1050 B.n155 VSUBS 0.00732f
C1051 B.n156 VSUBS 0.00732f
C1052 B.n157 VSUBS 0.00732f
C1053 B.n158 VSUBS 0.00732f
C1054 B.n159 VSUBS 0.00732f
C1055 B.n160 VSUBS 0.00732f
C1056 B.n161 VSUBS 0.00732f
C1057 B.n162 VSUBS 0.00732f
C1058 B.n163 VSUBS 0.017783f
C1059 B.n164 VSUBS 0.00732f
C1060 B.n165 VSUBS 0.00732f
C1061 B.n166 VSUBS 0.00732f
C1062 B.n167 VSUBS 0.00732f
C1063 B.n168 VSUBS 0.00732f
C1064 B.n169 VSUBS 0.00732f
C1065 B.n170 VSUBS 0.00732f
C1066 B.n171 VSUBS 0.00732f
C1067 B.n172 VSUBS 0.00732f
C1068 B.n173 VSUBS 0.00732f
C1069 B.n174 VSUBS 0.00732f
C1070 B.n175 VSUBS 0.00732f
C1071 B.n176 VSUBS 0.00732f
C1072 B.n177 VSUBS 0.00732f
C1073 B.n178 VSUBS 0.00732f
C1074 B.n179 VSUBS 0.00732f
C1075 B.n180 VSUBS 0.00732f
C1076 B.n181 VSUBS 0.00732f
C1077 B.n182 VSUBS 0.017783f
C1078 B.n183 VSUBS 0.018386f
C1079 B.n184 VSUBS 0.018386f
C1080 B.n185 VSUBS 0.00732f
C1081 B.n186 VSUBS 0.00732f
C1082 B.n187 VSUBS 0.00732f
C1083 B.n188 VSUBS 0.00732f
C1084 B.n189 VSUBS 0.00732f
C1085 B.n190 VSUBS 0.00732f
C1086 B.n191 VSUBS 0.00732f
C1087 B.n192 VSUBS 0.00732f
C1088 B.n193 VSUBS 0.00732f
C1089 B.n194 VSUBS 0.00732f
C1090 B.n195 VSUBS 0.00732f
C1091 B.n196 VSUBS 0.00732f
C1092 B.n197 VSUBS 0.00732f
C1093 B.n198 VSUBS 0.00732f
C1094 B.n199 VSUBS 0.00732f
C1095 B.n200 VSUBS 0.00732f
C1096 B.n201 VSUBS 0.00732f
C1097 B.n202 VSUBS 0.00732f
C1098 B.n203 VSUBS 0.00732f
C1099 B.n204 VSUBS 0.00732f
C1100 B.n205 VSUBS 0.00732f
C1101 B.n206 VSUBS 0.00732f
C1102 B.n207 VSUBS 0.00732f
C1103 B.n208 VSUBS 0.00732f
C1104 B.n209 VSUBS 0.00732f
C1105 B.n210 VSUBS 0.00732f
C1106 B.n211 VSUBS 0.00732f
C1107 B.n212 VSUBS 0.00732f
C1108 B.n213 VSUBS 0.00732f
C1109 B.n214 VSUBS 0.00732f
C1110 B.n215 VSUBS 0.00732f
C1111 B.n216 VSUBS 0.00732f
C1112 B.n217 VSUBS 0.00732f
C1113 B.n218 VSUBS 0.00732f
C1114 B.n219 VSUBS 0.00732f
C1115 B.n220 VSUBS 0.00732f
C1116 B.n221 VSUBS 0.00732f
C1117 B.n222 VSUBS 0.00732f
C1118 B.n223 VSUBS 0.00732f
C1119 B.n224 VSUBS 0.00732f
C1120 B.n225 VSUBS 0.00732f
C1121 B.n226 VSUBS 0.00732f
C1122 B.n227 VSUBS 0.00732f
C1123 B.n228 VSUBS 0.00732f
C1124 B.n229 VSUBS 0.00732f
C1125 B.n230 VSUBS 0.00732f
C1126 B.n231 VSUBS 0.00732f
C1127 B.n232 VSUBS 0.00732f
C1128 B.n233 VSUBS 0.00732f
C1129 B.n234 VSUBS 0.00732f
C1130 B.n235 VSUBS 0.00732f
C1131 B.n236 VSUBS 0.00732f
C1132 B.n237 VSUBS 0.00732f
C1133 B.n238 VSUBS 0.00732f
C1134 B.n239 VSUBS 0.00732f
C1135 B.n240 VSUBS 0.00732f
C1136 B.n241 VSUBS 0.00732f
C1137 B.n242 VSUBS 0.00732f
C1138 B.n243 VSUBS 0.00732f
C1139 B.n244 VSUBS 0.00732f
C1140 B.n245 VSUBS 0.00732f
C1141 B.n246 VSUBS 0.00732f
C1142 B.n247 VSUBS 0.00732f
C1143 B.n248 VSUBS 0.00732f
C1144 B.n249 VSUBS 0.00732f
C1145 B.n250 VSUBS 0.00732f
C1146 B.n251 VSUBS 0.00732f
C1147 B.n252 VSUBS 0.00732f
C1148 B.n253 VSUBS 0.00732f
C1149 B.n254 VSUBS 0.00732f
C1150 B.n255 VSUBS 0.00732f
C1151 B.n256 VSUBS 0.00732f
C1152 B.n257 VSUBS 0.00732f
C1153 B.n258 VSUBS 0.00732f
C1154 B.n259 VSUBS 0.00732f
C1155 B.n260 VSUBS 0.00732f
C1156 B.n261 VSUBS 0.00732f
C1157 B.n262 VSUBS 0.00732f
C1158 B.n263 VSUBS 0.00732f
C1159 B.n264 VSUBS 0.00732f
C1160 B.n265 VSUBS 0.00732f
C1161 B.n266 VSUBS 0.00732f
C1162 B.n267 VSUBS 0.00732f
C1163 B.n268 VSUBS 0.00732f
C1164 B.n269 VSUBS 0.00732f
C1165 B.n270 VSUBS 0.00732f
C1166 B.n271 VSUBS 0.00732f
C1167 B.n272 VSUBS 0.00732f
C1168 B.n273 VSUBS 0.00732f
C1169 B.n274 VSUBS 0.00732f
C1170 B.n275 VSUBS 0.00732f
C1171 B.n276 VSUBS 0.00732f
C1172 B.n277 VSUBS 0.00732f
C1173 B.n278 VSUBS 0.004844f
C1174 B.n279 VSUBS 0.01696f
C1175 B.n280 VSUBS 0.006136f
C1176 B.n281 VSUBS 0.00732f
C1177 B.n282 VSUBS 0.00732f
C1178 B.n283 VSUBS 0.00732f
C1179 B.n284 VSUBS 0.00732f
C1180 B.n285 VSUBS 0.00732f
C1181 B.n286 VSUBS 0.00732f
C1182 B.n287 VSUBS 0.00732f
C1183 B.n288 VSUBS 0.00732f
C1184 B.n289 VSUBS 0.00732f
C1185 B.n290 VSUBS 0.00732f
C1186 B.n291 VSUBS 0.00732f
C1187 B.t2 VSUBS 0.406853f
C1188 B.t1 VSUBS 0.41434f
C1189 B.t0 VSUBS 0.204946f
C1190 B.n292 VSUBS 0.407854f
C1191 B.n293 VSUBS 0.352851f
C1192 B.n294 VSUBS 0.01696f
C1193 B.n295 VSUBS 0.006136f
C1194 B.n296 VSUBS 0.00732f
C1195 B.n297 VSUBS 0.00732f
C1196 B.n298 VSUBS 0.00732f
C1197 B.n299 VSUBS 0.00732f
C1198 B.n300 VSUBS 0.00732f
C1199 B.n301 VSUBS 0.00732f
C1200 B.n302 VSUBS 0.00732f
C1201 B.n303 VSUBS 0.00732f
C1202 B.n304 VSUBS 0.00732f
C1203 B.n305 VSUBS 0.00732f
C1204 B.n306 VSUBS 0.00732f
C1205 B.n307 VSUBS 0.00732f
C1206 B.n308 VSUBS 0.00732f
C1207 B.n309 VSUBS 0.00732f
C1208 B.n310 VSUBS 0.00732f
C1209 B.n311 VSUBS 0.00732f
C1210 B.n312 VSUBS 0.00732f
C1211 B.n313 VSUBS 0.00732f
C1212 B.n314 VSUBS 0.00732f
C1213 B.n315 VSUBS 0.00732f
C1214 B.n316 VSUBS 0.00732f
C1215 B.n317 VSUBS 0.00732f
C1216 B.n318 VSUBS 0.00732f
C1217 B.n319 VSUBS 0.00732f
C1218 B.n320 VSUBS 0.00732f
C1219 B.n321 VSUBS 0.00732f
C1220 B.n322 VSUBS 0.00732f
C1221 B.n323 VSUBS 0.00732f
C1222 B.n324 VSUBS 0.00732f
C1223 B.n325 VSUBS 0.00732f
C1224 B.n326 VSUBS 0.00732f
C1225 B.n327 VSUBS 0.00732f
C1226 B.n328 VSUBS 0.00732f
C1227 B.n329 VSUBS 0.00732f
C1228 B.n330 VSUBS 0.00732f
C1229 B.n331 VSUBS 0.00732f
C1230 B.n332 VSUBS 0.00732f
C1231 B.n333 VSUBS 0.00732f
C1232 B.n334 VSUBS 0.00732f
C1233 B.n335 VSUBS 0.00732f
C1234 B.n336 VSUBS 0.00732f
C1235 B.n337 VSUBS 0.00732f
C1236 B.n338 VSUBS 0.00732f
C1237 B.n339 VSUBS 0.00732f
C1238 B.n340 VSUBS 0.00732f
C1239 B.n341 VSUBS 0.00732f
C1240 B.n342 VSUBS 0.00732f
C1241 B.n343 VSUBS 0.00732f
C1242 B.n344 VSUBS 0.00732f
C1243 B.n345 VSUBS 0.00732f
C1244 B.n346 VSUBS 0.00732f
C1245 B.n347 VSUBS 0.00732f
C1246 B.n348 VSUBS 0.00732f
C1247 B.n349 VSUBS 0.00732f
C1248 B.n350 VSUBS 0.00732f
C1249 B.n351 VSUBS 0.00732f
C1250 B.n352 VSUBS 0.00732f
C1251 B.n353 VSUBS 0.00732f
C1252 B.n354 VSUBS 0.00732f
C1253 B.n355 VSUBS 0.00732f
C1254 B.n356 VSUBS 0.00732f
C1255 B.n357 VSUBS 0.00732f
C1256 B.n358 VSUBS 0.00732f
C1257 B.n359 VSUBS 0.00732f
C1258 B.n360 VSUBS 0.00732f
C1259 B.n361 VSUBS 0.00732f
C1260 B.n362 VSUBS 0.00732f
C1261 B.n363 VSUBS 0.00732f
C1262 B.n364 VSUBS 0.00732f
C1263 B.n365 VSUBS 0.00732f
C1264 B.n366 VSUBS 0.00732f
C1265 B.n367 VSUBS 0.00732f
C1266 B.n368 VSUBS 0.00732f
C1267 B.n369 VSUBS 0.00732f
C1268 B.n370 VSUBS 0.00732f
C1269 B.n371 VSUBS 0.00732f
C1270 B.n372 VSUBS 0.00732f
C1271 B.n373 VSUBS 0.00732f
C1272 B.n374 VSUBS 0.00732f
C1273 B.n375 VSUBS 0.00732f
C1274 B.n376 VSUBS 0.00732f
C1275 B.n377 VSUBS 0.00732f
C1276 B.n378 VSUBS 0.00732f
C1277 B.n379 VSUBS 0.00732f
C1278 B.n380 VSUBS 0.00732f
C1279 B.n381 VSUBS 0.00732f
C1280 B.n382 VSUBS 0.00732f
C1281 B.n383 VSUBS 0.00732f
C1282 B.n384 VSUBS 0.00732f
C1283 B.n385 VSUBS 0.00732f
C1284 B.n386 VSUBS 0.00732f
C1285 B.n387 VSUBS 0.00732f
C1286 B.n388 VSUBS 0.00732f
C1287 B.n389 VSUBS 0.00732f
C1288 B.n390 VSUBS 0.00732f
C1289 B.n391 VSUBS 0.017589f
C1290 B.n392 VSUBS 0.018386f
C1291 B.n393 VSUBS 0.017783f
C1292 B.n394 VSUBS 0.00732f
C1293 B.n395 VSUBS 0.00732f
C1294 B.n396 VSUBS 0.00732f
C1295 B.n397 VSUBS 0.00732f
C1296 B.n398 VSUBS 0.00732f
C1297 B.n399 VSUBS 0.00732f
C1298 B.n400 VSUBS 0.00732f
C1299 B.n401 VSUBS 0.00732f
C1300 B.n402 VSUBS 0.00732f
C1301 B.n403 VSUBS 0.00732f
C1302 B.n404 VSUBS 0.00732f
C1303 B.n405 VSUBS 0.00732f
C1304 B.n406 VSUBS 0.00732f
C1305 B.n407 VSUBS 0.00732f
C1306 B.n408 VSUBS 0.00732f
C1307 B.n409 VSUBS 0.00732f
C1308 B.n410 VSUBS 0.00732f
C1309 B.n411 VSUBS 0.00732f
C1310 B.n412 VSUBS 0.00732f
C1311 B.n413 VSUBS 0.00732f
C1312 B.n414 VSUBS 0.00732f
C1313 B.n415 VSUBS 0.00732f
C1314 B.n416 VSUBS 0.00732f
C1315 B.n417 VSUBS 0.00732f
C1316 B.n418 VSUBS 0.00732f
C1317 B.n419 VSUBS 0.00732f
C1318 B.n420 VSUBS 0.00732f
C1319 B.n421 VSUBS 0.00732f
C1320 B.n422 VSUBS 0.00732f
C1321 B.n423 VSUBS 0.00732f
C1322 B.n424 VSUBS 0.00732f
C1323 B.n425 VSUBS 0.00732f
C1324 B.n426 VSUBS 0.00732f
C1325 B.n427 VSUBS 0.017783f
C1326 B.n428 VSUBS 0.017783f
C1327 B.n429 VSUBS 0.018386f
C1328 B.n430 VSUBS 0.00732f
C1329 B.n431 VSUBS 0.00732f
C1330 B.n432 VSUBS 0.00732f
C1331 B.n433 VSUBS 0.00732f
C1332 B.n434 VSUBS 0.00732f
C1333 B.n435 VSUBS 0.00732f
C1334 B.n436 VSUBS 0.00732f
C1335 B.n437 VSUBS 0.00732f
C1336 B.n438 VSUBS 0.00732f
C1337 B.n439 VSUBS 0.00732f
C1338 B.n440 VSUBS 0.00732f
C1339 B.n441 VSUBS 0.00732f
C1340 B.n442 VSUBS 0.00732f
C1341 B.n443 VSUBS 0.00732f
C1342 B.n444 VSUBS 0.00732f
C1343 B.n445 VSUBS 0.00732f
C1344 B.n446 VSUBS 0.00732f
C1345 B.n447 VSUBS 0.00732f
C1346 B.n448 VSUBS 0.00732f
C1347 B.n449 VSUBS 0.00732f
C1348 B.n450 VSUBS 0.00732f
C1349 B.n451 VSUBS 0.00732f
C1350 B.n452 VSUBS 0.00732f
C1351 B.n453 VSUBS 0.00732f
C1352 B.n454 VSUBS 0.00732f
C1353 B.n455 VSUBS 0.00732f
C1354 B.n456 VSUBS 0.00732f
C1355 B.n457 VSUBS 0.00732f
C1356 B.n458 VSUBS 0.00732f
C1357 B.n459 VSUBS 0.00732f
C1358 B.n460 VSUBS 0.00732f
C1359 B.n461 VSUBS 0.00732f
C1360 B.n462 VSUBS 0.00732f
C1361 B.n463 VSUBS 0.00732f
C1362 B.n464 VSUBS 0.00732f
C1363 B.n465 VSUBS 0.00732f
C1364 B.n466 VSUBS 0.00732f
C1365 B.n467 VSUBS 0.00732f
C1366 B.n468 VSUBS 0.00732f
C1367 B.n469 VSUBS 0.00732f
C1368 B.n470 VSUBS 0.00732f
C1369 B.n471 VSUBS 0.00732f
C1370 B.n472 VSUBS 0.00732f
C1371 B.n473 VSUBS 0.00732f
C1372 B.n474 VSUBS 0.00732f
C1373 B.n475 VSUBS 0.00732f
C1374 B.n476 VSUBS 0.00732f
C1375 B.n477 VSUBS 0.00732f
C1376 B.n478 VSUBS 0.00732f
C1377 B.n479 VSUBS 0.00732f
C1378 B.n480 VSUBS 0.00732f
C1379 B.n481 VSUBS 0.00732f
C1380 B.n482 VSUBS 0.00732f
C1381 B.n483 VSUBS 0.00732f
C1382 B.n484 VSUBS 0.00732f
C1383 B.n485 VSUBS 0.00732f
C1384 B.n486 VSUBS 0.00732f
C1385 B.n487 VSUBS 0.00732f
C1386 B.n488 VSUBS 0.00732f
C1387 B.n489 VSUBS 0.00732f
C1388 B.n490 VSUBS 0.00732f
C1389 B.n491 VSUBS 0.00732f
C1390 B.n492 VSUBS 0.00732f
C1391 B.n493 VSUBS 0.00732f
C1392 B.n494 VSUBS 0.00732f
C1393 B.n495 VSUBS 0.00732f
C1394 B.n496 VSUBS 0.00732f
C1395 B.n497 VSUBS 0.00732f
C1396 B.n498 VSUBS 0.00732f
C1397 B.n499 VSUBS 0.00732f
C1398 B.n500 VSUBS 0.00732f
C1399 B.n501 VSUBS 0.00732f
C1400 B.n502 VSUBS 0.00732f
C1401 B.n503 VSUBS 0.00732f
C1402 B.n504 VSUBS 0.00732f
C1403 B.n505 VSUBS 0.00732f
C1404 B.n506 VSUBS 0.00732f
C1405 B.n507 VSUBS 0.00732f
C1406 B.n508 VSUBS 0.00732f
C1407 B.n509 VSUBS 0.00732f
C1408 B.n510 VSUBS 0.00732f
C1409 B.n511 VSUBS 0.00732f
C1410 B.n512 VSUBS 0.00732f
C1411 B.n513 VSUBS 0.00732f
C1412 B.n514 VSUBS 0.00732f
C1413 B.n515 VSUBS 0.00732f
C1414 B.n516 VSUBS 0.00732f
C1415 B.n517 VSUBS 0.00732f
C1416 B.n518 VSUBS 0.00732f
C1417 B.n519 VSUBS 0.00732f
C1418 B.n520 VSUBS 0.00732f
C1419 B.n521 VSUBS 0.00732f
C1420 B.n522 VSUBS 0.00732f
C1421 B.n523 VSUBS 0.004844f
C1422 B.n524 VSUBS 0.00732f
C1423 B.n525 VSUBS 0.00732f
C1424 B.n526 VSUBS 0.006136f
C1425 B.n527 VSUBS 0.00732f
C1426 B.n528 VSUBS 0.00732f
C1427 B.n529 VSUBS 0.00732f
C1428 B.n530 VSUBS 0.00732f
C1429 B.n531 VSUBS 0.00732f
C1430 B.n532 VSUBS 0.00732f
C1431 B.n533 VSUBS 0.00732f
C1432 B.n534 VSUBS 0.00732f
C1433 B.n535 VSUBS 0.00732f
C1434 B.n536 VSUBS 0.00732f
C1435 B.n537 VSUBS 0.00732f
C1436 B.n538 VSUBS 0.006136f
C1437 B.n539 VSUBS 0.01696f
C1438 B.n540 VSUBS 0.004844f
C1439 B.n541 VSUBS 0.00732f
C1440 B.n542 VSUBS 0.00732f
C1441 B.n543 VSUBS 0.00732f
C1442 B.n544 VSUBS 0.00732f
C1443 B.n545 VSUBS 0.00732f
C1444 B.n546 VSUBS 0.00732f
C1445 B.n547 VSUBS 0.00732f
C1446 B.n548 VSUBS 0.00732f
C1447 B.n549 VSUBS 0.00732f
C1448 B.n550 VSUBS 0.00732f
C1449 B.n551 VSUBS 0.00732f
C1450 B.n552 VSUBS 0.00732f
C1451 B.n553 VSUBS 0.00732f
C1452 B.n554 VSUBS 0.00732f
C1453 B.n555 VSUBS 0.00732f
C1454 B.n556 VSUBS 0.00732f
C1455 B.n557 VSUBS 0.00732f
C1456 B.n558 VSUBS 0.00732f
C1457 B.n559 VSUBS 0.00732f
C1458 B.n560 VSUBS 0.00732f
C1459 B.n561 VSUBS 0.00732f
C1460 B.n562 VSUBS 0.00732f
C1461 B.n563 VSUBS 0.00732f
C1462 B.n564 VSUBS 0.00732f
C1463 B.n565 VSUBS 0.00732f
C1464 B.n566 VSUBS 0.00732f
C1465 B.n567 VSUBS 0.00732f
C1466 B.n568 VSUBS 0.00732f
C1467 B.n569 VSUBS 0.00732f
C1468 B.n570 VSUBS 0.00732f
C1469 B.n571 VSUBS 0.00732f
C1470 B.n572 VSUBS 0.00732f
C1471 B.n573 VSUBS 0.00732f
C1472 B.n574 VSUBS 0.00732f
C1473 B.n575 VSUBS 0.00732f
C1474 B.n576 VSUBS 0.00732f
C1475 B.n577 VSUBS 0.00732f
C1476 B.n578 VSUBS 0.00732f
C1477 B.n579 VSUBS 0.00732f
C1478 B.n580 VSUBS 0.00732f
C1479 B.n581 VSUBS 0.00732f
C1480 B.n582 VSUBS 0.00732f
C1481 B.n583 VSUBS 0.00732f
C1482 B.n584 VSUBS 0.00732f
C1483 B.n585 VSUBS 0.00732f
C1484 B.n586 VSUBS 0.00732f
C1485 B.n587 VSUBS 0.00732f
C1486 B.n588 VSUBS 0.00732f
C1487 B.n589 VSUBS 0.00732f
C1488 B.n590 VSUBS 0.00732f
C1489 B.n591 VSUBS 0.00732f
C1490 B.n592 VSUBS 0.00732f
C1491 B.n593 VSUBS 0.00732f
C1492 B.n594 VSUBS 0.00732f
C1493 B.n595 VSUBS 0.00732f
C1494 B.n596 VSUBS 0.00732f
C1495 B.n597 VSUBS 0.00732f
C1496 B.n598 VSUBS 0.00732f
C1497 B.n599 VSUBS 0.00732f
C1498 B.n600 VSUBS 0.00732f
C1499 B.n601 VSUBS 0.00732f
C1500 B.n602 VSUBS 0.00732f
C1501 B.n603 VSUBS 0.00732f
C1502 B.n604 VSUBS 0.00732f
C1503 B.n605 VSUBS 0.00732f
C1504 B.n606 VSUBS 0.00732f
C1505 B.n607 VSUBS 0.00732f
C1506 B.n608 VSUBS 0.00732f
C1507 B.n609 VSUBS 0.00732f
C1508 B.n610 VSUBS 0.00732f
C1509 B.n611 VSUBS 0.00732f
C1510 B.n612 VSUBS 0.00732f
C1511 B.n613 VSUBS 0.00732f
C1512 B.n614 VSUBS 0.00732f
C1513 B.n615 VSUBS 0.00732f
C1514 B.n616 VSUBS 0.00732f
C1515 B.n617 VSUBS 0.00732f
C1516 B.n618 VSUBS 0.00732f
C1517 B.n619 VSUBS 0.00732f
C1518 B.n620 VSUBS 0.00732f
C1519 B.n621 VSUBS 0.00732f
C1520 B.n622 VSUBS 0.00732f
C1521 B.n623 VSUBS 0.00732f
C1522 B.n624 VSUBS 0.00732f
C1523 B.n625 VSUBS 0.00732f
C1524 B.n626 VSUBS 0.00732f
C1525 B.n627 VSUBS 0.00732f
C1526 B.n628 VSUBS 0.00732f
C1527 B.n629 VSUBS 0.00732f
C1528 B.n630 VSUBS 0.00732f
C1529 B.n631 VSUBS 0.00732f
C1530 B.n632 VSUBS 0.00732f
C1531 B.n633 VSUBS 0.00732f
C1532 B.n634 VSUBS 0.018386f
C1533 B.n635 VSUBS 0.018386f
C1534 B.n636 VSUBS 0.017783f
C1535 B.n637 VSUBS 0.00732f
C1536 B.n638 VSUBS 0.00732f
C1537 B.n639 VSUBS 0.00732f
C1538 B.n640 VSUBS 0.00732f
C1539 B.n641 VSUBS 0.00732f
C1540 B.n642 VSUBS 0.00732f
C1541 B.n643 VSUBS 0.00732f
C1542 B.n644 VSUBS 0.00732f
C1543 B.n645 VSUBS 0.00732f
C1544 B.n646 VSUBS 0.00732f
C1545 B.n647 VSUBS 0.00732f
C1546 B.n648 VSUBS 0.00732f
C1547 B.n649 VSUBS 0.00732f
C1548 B.n650 VSUBS 0.00732f
C1549 B.n651 VSUBS 0.009552f
C1550 B.n652 VSUBS 0.010176f
C1551 B.n653 VSUBS 0.020235f
.ends

