* NGSPICE file created from diff_pair_sample_0385.ext - technology: sky130A

.subckt diff_pair_sample_0385 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t14 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=3
X1 B.t11 B.t9 B.t10 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=3
X2 B.t8 B.t6 B.t7 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=3
X3 VTAIL.t15 VN.t1 VDD2.t6 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=3
X4 B.t5 B.t3 B.t4 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=3
X5 VDD2.t5 VN.t2 VTAIL.t13 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
X6 B.t2 B.t0 B.t1 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=3
X7 VDD2.t4 VN.t3 VTAIL.t11 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=3
X8 VTAIL.t12 VN.t4 VDD2.t3 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
X9 VDD1.t7 VP.t0 VTAIL.t6 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=3
X10 VDD1.t6 VP.t1 VTAIL.t4 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
X11 VTAIL.t5 VP.t2 VDD1.t5 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=3
X12 VTAIL.t9 VN.t5 VDD2.t2 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
X13 VDD2.t1 VN.t6 VTAIL.t10 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
X14 VDD1.t4 VP.t3 VTAIL.t2 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
X15 VDD1.t3 VP.t4 VTAIL.t7 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=3
X16 VTAIL.t3 VP.t5 VDD1.t2 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
X17 VTAIL.t8 VN.t7 VDD2.t0 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=3
X18 VTAIL.t1 VP.t6 VDD1.t1 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=3
X19 VTAIL.t0 VP.t7 VDD1.t0 w_n4300_n2640# sky130_fd_pr__pfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=3
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n50 VN.n49 161.3
R7 VN.n48 VN.n35 161.3
R8 VN.n47 VN.n46 161.3
R9 VN.n45 VN.n36 161.3
R10 VN.n44 VN.n43 161.3
R11 VN.n42 VN.n37 161.3
R12 VN.n41 VN.n40 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n4 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n14 VN.n5 161.3
R23 VN.n13 VN.n12 161.3
R24 VN.n11 VN.n6 161.3
R25 VN.n10 VN.n9 161.3
R26 VN.n38 VN.t3 98.9905
R27 VN.n7 VN.t1 98.9905
R28 VN.n8 VN.t6 67.1592
R29 VN.n20 VN.t5 67.1592
R30 VN.n0 VN.t0 67.1592
R31 VN.n39 VN.t4 67.1592
R32 VN.n51 VN.t2 67.1592
R33 VN.n31 VN.t7 67.1592
R34 VN.n8 VN.n7 66.0722
R35 VN.n39 VN.n38 66.0722
R36 VN.n30 VN.n0 65.8996
R37 VN.n61 VN.n31 65.8996
R38 VN.n26 VN.n2 56.5617
R39 VN.n57 VN.n33 56.5617
R40 VN VN.n61 50.3618
R41 VN.n14 VN.n13 40.577
R42 VN.n15 VN.n14 40.577
R43 VN.n45 VN.n44 40.577
R44 VN.n46 VN.n45 40.577
R45 VN.n9 VN.n6 24.5923
R46 VN.n13 VN.n6 24.5923
R47 VN.n15 VN.n4 24.5923
R48 VN.n19 VN.n4 24.5923
R49 VN.n22 VN.n21 24.5923
R50 VN.n22 VN.n2 24.5923
R51 VN.n27 VN.n26 24.5923
R52 VN.n28 VN.n27 24.5923
R53 VN.n44 VN.n37 24.5923
R54 VN.n40 VN.n37 24.5923
R55 VN.n53 VN.n33 24.5923
R56 VN.n53 VN.n52 24.5923
R57 VN.n50 VN.n35 24.5923
R58 VN.n46 VN.n35 24.5923
R59 VN.n59 VN.n58 24.5923
R60 VN.n58 VN.n57 24.5923
R61 VN.n28 VN.n0 24.3464
R62 VN.n59 VN.n31 24.3464
R63 VN.n21 VN.n20 16.477
R64 VN.n52 VN.n51 16.477
R65 VN.n9 VN.n8 8.11581
R66 VN.n20 VN.n19 8.11581
R67 VN.n40 VN.n39 8.11581
R68 VN.n51 VN.n50 8.11581
R69 VN.n41 VN.n38 5.23312
R70 VN.n10 VN.n7 5.23312
R71 VN.n61 VN.n60 0.354861
R72 VN.n30 VN.n29 0.354861
R73 VN VN.n30 0.267071
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n49 VN.n34 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n47 0.189894
R82 VN.n47 VN.n36 0.189894
R83 VN.n43 VN.n36 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n41 0.189894
R86 VN.n11 VN.n10 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n12 VN.n5 0.189894
R89 VN.n16 VN.n5 0.189894
R90 VN.n17 VN.n16 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n18 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VTAIL.n11 VTAIL.t5 72.3729
R99 VTAIL.n10 VTAIL.t11 72.3729
R100 VTAIL.n7 VTAIL.t8 72.3729
R101 VTAIL.n14 VTAIL.t7 72.3728
R102 VTAIL.n15 VTAIL.t14 72.3728
R103 VTAIL.n2 VTAIL.t15 72.3728
R104 VTAIL.n3 VTAIL.t6 72.3728
R105 VTAIL.n6 VTAIL.t1 72.3728
R106 VTAIL.n13 VTAIL.n12 68.4849
R107 VTAIL.n9 VTAIL.n8 68.4849
R108 VTAIL.n1 VTAIL.n0 68.4846
R109 VTAIL.n5 VTAIL.n4 68.4846
R110 VTAIL.n15 VTAIL.n14 22.4445
R111 VTAIL.n7 VTAIL.n6 22.4445
R112 VTAIL.n0 VTAIL.t10 3.88866
R113 VTAIL.n0 VTAIL.t9 3.88866
R114 VTAIL.n4 VTAIL.t2 3.88866
R115 VTAIL.n4 VTAIL.t0 3.88866
R116 VTAIL.n12 VTAIL.t4 3.88866
R117 VTAIL.n12 VTAIL.t3 3.88866
R118 VTAIL.n8 VTAIL.t13 3.88866
R119 VTAIL.n8 VTAIL.t12 3.88866
R120 VTAIL.n9 VTAIL.n7 2.87119
R121 VTAIL.n10 VTAIL.n9 2.87119
R122 VTAIL.n13 VTAIL.n11 2.87119
R123 VTAIL.n14 VTAIL.n13 2.87119
R124 VTAIL.n6 VTAIL.n5 2.87119
R125 VTAIL.n5 VTAIL.n3 2.87119
R126 VTAIL.n2 VTAIL.n1 2.87119
R127 VTAIL VTAIL.n15 2.813
R128 VTAIL.n11 VTAIL.n10 0.470328
R129 VTAIL.n3 VTAIL.n2 0.470328
R130 VTAIL VTAIL.n1 0.0586897
R131 VDD2.n2 VDD2.n1 86.5434
R132 VDD2.n2 VDD2.n0 86.5434
R133 VDD2 VDD2.n5 86.5406
R134 VDD2.n4 VDD2.n3 85.1636
R135 VDD2.n4 VDD2.n2 43.8403
R136 VDD2.n5 VDD2.t3 3.88866
R137 VDD2.n5 VDD2.t4 3.88866
R138 VDD2.n3 VDD2.t0 3.88866
R139 VDD2.n3 VDD2.t5 3.88866
R140 VDD2.n1 VDD2.t2 3.88866
R141 VDD2.n1 VDD2.t7 3.88866
R142 VDD2.n0 VDD2.t6 3.88866
R143 VDD2.n0 VDD2.t1 3.88866
R144 VDD2 VDD2.n4 1.49403
R145 B.n561 B.n70 585
R146 B.n563 B.n562 585
R147 B.n564 B.n69 585
R148 B.n566 B.n565 585
R149 B.n567 B.n68 585
R150 B.n569 B.n568 585
R151 B.n570 B.n67 585
R152 B.n572 B.n571 585
R153 B.n573 B.n66 585
R154 B.n575 B.n574 585
R155 B.n576 B.n65 585
R156 B.n578 B.n577 585
R157 B.n579 B.n64 585
R158 B.n581 B.n580 585
R159 B.n582 B.n63 585
R160 B.n584 B.n583 585
R161 B.n585 B.n62 585
R162 B.n587 B.n586 585
R163 B.n588 B.n61 585
R164 B.n590 B.n589 585
R165 B.n591 B.n60 585
R166 B.n593 B.n592 585
R167 B.n594 B.n59 585
R168 B.n596 B.n595 585
R169 B.n597 B.n58 585
R170 B.n599 B.n598 585
R171 B.n600 B.n57 585
R172 B.n602 B.n601 585
R173 B.n603 B.n56 585
R174 B.n605 B.n604 585
R175 B.n606 B.n53 585
R176 B.n609 B.n608 585
R177 B.n610 B.n52 585
R178 B.n612 B.n611 585
R179 B.n613 B.n51 585
R180 B.n615 B.n614 585
R181 B.n616 B.n50 585
R182 B.n618 B.n617 585
R183 B.n619 B.n49 585
R184 B.n621 B.n620 585
R185 B.n623 B.n622 585
R186 B.n624 B.n45 585
R187 B.n626 B.n625 585
R188 B.n627 B.n44 585
R189 B.n629 B.n628 585
R190 B.n630 B.n43 585
R191 B.n632 B.n631 585
R192 B.n633 B.n42 585
R193 B.n635 B.n634 585
R194 B.n636 B.n41 585
R195 B.n638 B.n637 585
R196 B.n639 B.n40 585
R197 B.n641 B.n640 585
R198 B.n642 B.n39 585
R199 B.n644 B.n643 585
R200 B.n645 B.n38 585
R201 B.n647 B.n646 585
R202 B.n648 B.n37 585
R203 B.n650 B.n649 585
R204 B.n651 B.n36 585
R205 B.n653 B.n652 585
R206 B.n654 B.n35 585
R207 B.n656 B.n655 585
R208 B.n657 B.n34 585
R209 B.n659 B.n658 585
R210 B.n660 B.n33 585
R211 B.n662 B.n661 585
R212 B.n663 B.n32 585
R213 B.n665 B.n664 585
R214 B.n666 B.n31 585
R215 B.n668 B.n667 585
R216 B.n560 B.n559 585
R217 B.n558 B.n71 585
R218 B.n557 B.n556 585
R219 B.n555 B.n72 585
R220 B.n554 B.n553 585
R221 B.n552 B.n73 585
R222 B.n551 B.n550 585
R223 B.n549 B.n74 585
R224 B.n548 B.n547 585
R225 B.n546 B.n75 585
R226 B.n545 B.n544 585
R227 B.n543 B.n76 585
R228 B.n542 B.n541 585
R229 B.n540 B.n77 585
R230 B.n539 B.n538 585
R231 B.n537 B.n78 585
R232 B.n536 B.n535 585
R233 B.n534 B.n79 585
R234 B.n533 B.n532 585
R235 B.n531 B.n80 585
R236 B.n530 B.n529 585
R237 B.n528 B.n81 585
R238 B.n527 B.n526 585
R239 B.n525 B.n82 585
R240 B.n524 B.n523 585
R241 B.n522 B.n83 585
R242 B.n521 B.n520 585
R243 B.n519 B.n84 585
R244 B.n518 B.n517 585
R245 B.n516 B.n85 585
R246 B.n515 B.n514 585
R247 B.n513 B.n86 585
R248 B.n512 B.n511 585
R249 B.n510 B.n87 585
R250 B.n509 B.n508 585
R251 B.n507 B.n88 585
R252 B.n506 B.n505 585
R253 B.n504 B.n89 585
R254 B.n503 B.n502 585
R255 B.n501 B.n90 585
R256 B.n500 B.n499 585
R257 B.n498 B.n91 585
R258 B.n497 B.n496 585
R259 B.n495 B.n92 585
R260 B.n494 B.n493 585
R261 B.n492 B.n93 585
R262 B.n491 B.n490 585
R263 B.n489 B.n94 585
R264 B.n488 B.n487 585
R265 B.n486 B.n95 585
R266 B.n485 B.n484 585
R267 B.n483 B.n96 585
R268 B.n482 B.n481 585
R269 B.n480 B.n97 585
R270 B.n479 B.n478 585
R271 B.n477 B.n98 585
R272 B.n476 B.n475 585
R273 B.n474 B.n99 585
R274 B.n473 B.n472 585
R275 B.n471 B.n100 585
R276 B.n470 B.n469 585
R277 B.n468 B.n101 585
R278 B.n467 B.n466 585
R279 B.n465 B.n102 585
R280 B.n464 B.n463 585
R281 B.n462 B.n103 585
R282 B.n461 B.n460 585
R283 B.n459 B.n104 585
R284 B.n458 B.n457 585
R285 B.n456 B.n105 585
R286 B.n455 B.n454 585
R287 B.n453 B.n106 585
R288 B.n452 B.n451 585
R289 B.n450 B.n107 585
R290 B.n449 B.n448 585
R291 B.n447 B.n108 585
R292 B.n446 B.n445 585
R293 B.n444 B.n109 585
R294 B.n443 B.n442 585
R295 B.n441 B.n110 585
R296 B.n440 B.n439 585
R297 B.n438 B.n111 585
R298 B.n437 B.n436 585
R299 B.n435 B.n112 585
R300 B.n434 B.n433 585
R301 B.n432 B.n113 585
R302 B.n431 B.n430 585
R303 B.n429 B.n114 585
R304 B.n428 B.n427 585
R305 B.n426 B.n115 585
R306 B.n425 B.n424 585
R307 B.n423 B.n116 585
R308 B.n422 B.n421 585
R309 B.n420 B.n117 585
R310 B.n419 B.n418 585
R311 B.n417 B.n118 585
R312 B.n416 B.n415 585
R313 B.n414 B.n119 585
R314 B.n413 B.n412 585
R315 B.n411 B.n120 585
R316 B.n410 B.n409 585
R317 B.n408 B.n121 585
R318 B.n407 B.n406 585
R319 B.n405 B.n122 585
R320 B.n404 B.n403 585
R321 B.n402 B.n123 585
R322 B.n401 B.n400 585
R323 B.n399 B.n124 585
R324 B.n398 B.n397 585
R325 B.n396 B.n125 585
R326 B.n395 B.n394 585
R327 B.n393 B.n126 585
R328 B.n392 B.n391 585
R329 B.n390 B.n127 585
R330 B.n389 B.n388 585
R331 B.n281 B.n280 585
R332 B.n282 B.n167 585
R333 B.n284 B.n283 585
R334 B.n285 B.n166 585
R335 B.n287 B.n286 585
R336 B.n288 B.n165 585
R337 B.n290 B.n289 585
R338 B.n291 B.n164 585
R339 B.n293 B.n292 585
R340 B.n294 B.n163 585
R341 B.n296 B.n295 585
R342 B.n297 B.n162 585
R343 B.n299 B.n298 585
R344 B.n300 B.n161 585
R345 B.n302 B.n301 585
R346 B.n303 B.n160 585
R347 B.n305 B.n304 585
R348 B.n306 B.n159 585
R349 B.n308 B.n307 585
R350 B.n309 B.n158 585
R351 B.n311 B.n310 585
R352 B.n312 B.n157 585
R353 B.n314 B.n313 585
R354 B.n315 B.n156 585
R355 B.n317 B.n316 585
R356 B.n318 B.n155 585
R357 B.n320 B.n319 585
R358 B.n321 B.n154 585
R359 B.n323 B.n322 585
R360 B.n324 B.n153 585
R361 B.n326 B.n325 585
R362 B.n328 B.n327 585
R363 B.n329 B.n149 585
R364 B.n331 B.n330 585
R365 B.n332 B.n148 585
R366 B.n334 B.n333 585
R367 B.n335 B.n147 585
R368 B.n337 B.n336 585
R369 B.n338 B.n146 585
R370 B.n340 B.n339 585
R371 B.n342 B.n143 585
R372 B.n344 B.n343 585
R373 B.n345 B.n142 585
R374 B.n347 B.n346 585
R375 B.n348 B.n141 585
R376 B.n350 B.n349 585
R377 B.n351 B.n140 585
R378 B.n353 B.n352 585
R379 B.n354 B.n139 585
R380 B.n356 B.n355 585
R381 B.n357 B.n138 585
R382 B.n359 B.n358 585
R383 B.n360 B.n137 585
R384 B.n362 B.n361 585
R385 B.n363 B.n136 585
R386 B.n365 B.n364 585
R387 B.n366 B.n135 585
R388 B.n368 B.n367 585
R389 B.n369 B.n134 585
R390 B.n371 B.n370 585
R391 B.n372 B.n133 585
R392 B.n374 B.n373 585
R393 B.n375 B.n132 585
R394 B.n377 B.n376 585
R395 B.n378 B.n131 585
R396 B.n380 B.n379 585
R397 B.n381 B.n130 585
R398 B.n383 B.n382 585
R399 B.n384 B.n129 585
R400 B.n386 B.n385 585
R401 B.n387 B.n128 585
R402 B.n279 B.n168 585
R403 B.n278 B.n277 585
R404 B.n276 B.n169 585
R405 B.n275 B.n274 585
R406 B.n273 B.n170 585
R407 B.n272 B.n271 585
R408 B.n270 B.n171 585
R409 B.n269 B.n268 585
R410 B.n267 B.n172 585
R411 B.n266 B.n265 585
R412 B.n264 B.n173 585
R413 B.n263 B.n262 585
R414 B.n261 B.n174 585
R415 B.n260 B.n259 585
R416 B.n258 B.n175 585
R417 B.n257 B.n256 585
R418 B.n255 B.n176 585
R419 B.n254 B.n253 585
R420 B.n252 B.n177 585
R421 B.n251 B.n250 585
R422 B.n249 B.n178 585
R423 B.n248 B.n247 585
R424 B.n246 B.n179 585
R425 B.n245 B.n244 585
R426 B.n243 B.n180 585
R427 B.n242 B.n241 585
R428 B.n240 B.n181 585
R429 B.n239 B.n238 585
R430 B.n237 B.n182 585
R431 B.n236 B.n235 585
R432 B.n234 B.n183 585
R433 B.n233 B.n232 585
R434 B.n231 B.n184 585
R435 B.n230 B.n229 585
R436 B.n228 B.n185 585
R437 B.n227 B.n226 585
R438 B.n225 B.n186 585
R439 B.n224 B.n223 585
R440 B.n222 B.n187 585
R441 B.n221 B.n220 585
R442 B.n219 B.n188 585
R443 B.n218 B.n217 585
R444 B.n216 B.n189 585
R445 B.n215 B.n214 585
R446 B.n213 B.n190 585
R447 B.n212 B.n211 585
R448 B.n210 B.n191 585
R449 B.n209 B.n208 585
R450 B.n207 B.n192 585
R451 B.n206 B.n205 585
R452 B.n204 B.n193 585
R453 B.n203 B.n202 585
R454 B.n201 B.n194 585
R455 B.n200 B.n199 585
R456 B.n198 B.n195 585
R457 B.n197 B.n196 585
R458 B.n2 B.n0 585
R459 B.n753 B.n1 585
R460 B.n752 B.n751 585
R461 B.n750 B.n3 585
R462 B.n749 B.n748 585
R463 B.n747 B.n4 585
R464 B.n746 B.n745 585
R465 B.n744 B.n5 585
R466 B.n743 B.n742 585
R467 B.n741 B.n6 585
R468 B.n740 B.n739 585
R469 B.n738 B.n7 585
R470 B.n737 B.n736 585
R471 B.n735 B.n8 585
R472 B.n734 B.n733 585
R473 B.n732 B.n9 585
R474 B.n731 B.n730 585
R475 B.n729 B.n10 585
R476 B.n728 B.n727 585
R477 B.n726 B.n11 585
R478 B.n725 B.n724 585
R479 B.n723 B.n12 585
R480 B.n722 B.n721 585
R481 B.n720 B.n13 585
R482 B.n719 B.n718 585
R483 B.n717 B.n14 585
R484 B.n716 B.n715 585
R485 B.n714 B.n15 585
R486 B.n713 B.n712 585
R487 B.n711 B.n16 585
R488 B.n710 B.n709 585
R489 B.n708 B.n17 585
R490 B.n707 B.n706 585
R491 B.n705 B.n18 585
R492 B.n704 B.n703 585
R493 B.n702 B.n19 585
R494 B.n701 B.n700 585
R495 B.n699 B.n20 585
R496 B.n698 B.n697 585
R497 B.n696 B.n21 585
R498 B.n695 B.n694 585
R499 B.n693 B.n22 585
R500 B.n692 B.n691 585
R501 B.n690 B.n23 585
R502 B.n689 B.n688 585
R503 B.n687 B.n24 585
R504 B.n686 B.n685 585
R505 B.n684 B.n25 585
R506 B.n683 B.n682 585
R507 B.n681 B.n26 585
R508 B.n680 B.n679 585
R509 B.n678 B.n27 585
R510 B.n677 B.n676 585
R511 B.n675 B.n28 585
R512 B.n674 B.n673 585
R513 B.n672 B.n29 585
R514 B.n671 B.n670 585
R515 B.n669 B.n30 585
R516 B.n755 B.n754 585
R517 B.n280 B.n279 545.355
R518 B.n669 B.n668 545.355
R519 B.n388 B.n387 545.355
R520 B.n561 B.n560 545.355
R521 B.n144 B.t0 275.738
R522 B.n150 B.t3 275.738
R523 B.n46 B.t9 275.738
R524 B.n54 B.t6 275.738
R525 B.n144 B.t2 176.911
R526 B.n54 B.t7 176.911
R527 B.n150 B.t5 176.901
R528 B.n46 B.t10 176.901
R529 B.n279 B.n278 163.367
R530 B.n278 B.n169 163.367
R531 B.n274 B.n169 163.367
R532 B.n274 B.n273 163.367
R533 B.n273 B.n272 163.367
R534 B.n272 B.n171 163.367
R535 B.n268 B.n171 163.367
R536 B.n268 B.n267 163.367
R537 B.n267 B.n266 163.367
R538 B.n266 B.n173 163.367
R539 B.n262 B.n173 163.367
R540 B.n262 B.n261 163.367
R541 B.n261 B.n260 163.367
R542 B.n260 B.n175 163.367
R543 B.n256 B.n175 163.367
R544 B.n256 B.n255 163.367
R545 B.n255 B.n254 163.367
R546 B.n254 B.n177 163.367
R547 B.n250 B.n177 163.367
R548 B.n250 B.n249 163.367
R549 B.n249 B.n248 163.367
R550 B.n248 B.n179 163.367
R551 B.n244 B.n179 163.367
R552 B.n244 B.n243 163.367
R553 B.n243 B.n242 163.367
R554 B.n242 B.n181 163.367
R555 B.n238 B.n181 163.367
R556 B.n238 B.n237 163.367
R557 B.n237 B.n236 163.367
R558 B.n236 B.n183 163.367
R559 B.n232 B.n183 163.367
R560 B.n232 B.n231 163.367
R561 B.n231 B.n230 163.367
R562 B.n230 B.n185 163.367
R563 B.n226 B.n185 163.367
R564 B.n226 B.n225 163.367
R565 B.n225 B.n224 163.367
R566 B.n224 B.n187 163.367
R567 B.n220 B.n187 163.367
R568 B.n220 B.n219 163.367
R569 B.n219 B.n218 163.367
R570 B.n218 B.n189 163.367
R571 B.n214 B.n189 163.367
R572 B.n214 B.n213 163.367
R573 B.n213 B.n212 163.367
R574 B.n212 B.n191 163.367
R575 B.n208 B.n191 163.367
R576 B.n208 B.n207 163.367
R577 B.n207 B.n206 163.367
R578 B.n206 B.n193 163.367
R579 B.n202 B.n193 163.367
R580 B.n202 B.n201 163.367
R581 B.n201 B.n200 163.367
R582 B.n200 B.n195 163.367
R583 B.n196 B.n195 163.367
R584 B.n196 B.n2 163.367
R585 B.n754 B.n2 163.367
R586 B.n754 B.n753 163.367
R587 B.n753 B.n752 163.367
R588 B.n752 B.n3 163.367
R589 B.n748 B.n3 163.367
R590 B.n748 B.n747 163.367
R591 B.n747 B.n746 163.367
R592 B.n746 B.n5 163.367
R593 B.n742 B.n5 163.367
R594 B.n742 B.n741 163.367
R595 B.n741 B.n740 163.367
R596 B.n740 B.n7 163.367
R597 B.n736 B.n7 163.367
R598 B.n736 B.n735 163.367
R599 B.n735 B.n734 163.367
R600 B.n734 B.n9 163.367
R601 B.n730 B.n9 163.367
R602 B.n730 B.n729 163.367
R603 B.n729 B.n728 163.367
R604 B.n728 B.n11 163.367
R605 B.n724 B.n11 163.367
R606 B.n724 B.n723 163.367
R607 B.n723 B.n722 163.367
R608 B.n722 B.n13 163.367
R609 B.n718 B.n13 163.367
R610 B.n718 B.n717 163.367
R611 B.n717 B.n716 163.367
R612 B.n716 B.n15 163.367
R613 B.n712 B.n15 163.367
R614 B.n712 B.n711 163.367
R615 B.n711 B.n710 163.367
R616 B.n710 B.n17 163.367
R617 B.n706 B.n17 163.367
R618 B.n706 B.n705 163.367
R619 B.n705 B.n704 163.367
R620 B.n704 B.n19 163.367
R621 B.n700 B.n19 163.367
R622 B.n700 B.n699 163.367
R623 B.n699 B.n698 163.367
R624 B.n698 B.n21 163.367
R625 B.n694 B.n21 163.367
R626 B.n694 B.n693 163.367
R627 B.n693 B.n692 163.367
R628 B.n692 B.n23 163.367
R629 B.n688 B.n23 163.367
R630 B.n688 B.n687 163.367
R631 B.n687 B.n686 163.367
R632 B.n686 B.n25 163.367
R633 B.n682 B.n25 163.367
R634 B.n682 B.n681 163.367
R635 B.n681 B.n680 163.367
R636 B.n680 B.n27 163.367
R637 B.n676 B.n27 163.367
R638 B.n676 B.n675 163.367
R639 B.n675 B.n674 163.367
R640 B.n674 B.n29 163.367
R641 B.n670 B.n29 163.367
R642 B.n670 B.n669 163.367
R643 B.n280 B.n167 163.367
R644 B.n284 B.n167 163.367
R645 B.n285 B.n284 163.367
R646 B.n286 B.n285 163.367
R647 B.n286 B.n165 163.367
R648 B.n290 B.n165 163.367
R649 B.n291 B.n290 163.367
R650 B.n292 B.n291 163.367
R651 B.n292 B.n163 163.367
R652 B.n296 B.n163 163.367
R653 B.n297 B.n296 163.367
R654 B.n298 B.n297 163.367
R655 B.n298 B.n161 163.367
R656 B.n302 B.n161 163.367
R657 B.n303 B.n302 163.367
R658 B.n304 B.n303 163.367
R659 B.n304 B.n159 163.367
R660 B.n308 B.n159 163.367
R661 B.n309 B.n308 163.367
R662 B.n310 B.n309 163.367
R663 B.n310 B.n157 163.367
R664 B.n314 B.n157 163.367
R665 B.n315 B.n314 163.367
R666 B.n316 B.n315 163.367
R667 B.n316 B.n155 163.367
R668 B.n320 B.n155 163.367
R669 B.n321 B.n320 163.367
R670 B.n322 B.n321 163.367
R671 B.n322 B.n153 163.367
R672 B.n326 B.n153 163.367
R673 B.n327 B.n326 163.367
R674 B.n327 B.n149 163.367
R675 B.n331 B.n149 163.367
R676 B.n332 B.n331 163.367
R677 B.n333 B.n332 163.367
R678 B.n333 B.n147 163.367
R679 B.n337 B.n147 163.367
R680 B.n338 B.n337 163.367
R681 B.n339 B.n338 163.367
R682 B.n339 B.n143 163.367
R683 B.n344 B.n143 163.367
R684 B.n345 B.n344 163.367
R685 B.n346 B.n345 163.367
R686 B.n346 B.n141 163.367
R687 B.n350 B.n141 163.367
R688 B.n351 B.n350 163.367
R689 B.n352 B.n351 163.367
R690 B.n352 B.n139 163.367
R691 B.n356 B.n139 163.367
R692 B.n357 B.n356 163.367
R693 B.n358 B.n357 163.367
R694 B.n358 B.n137 163.367
R695 B.n362 B.n137 163.367
R696 B.n363 B.n362 163.367
R697 B.n364 B.n363 163.367
R698 B.n364 B.n135 163.367
R699 B.n368 B.n135 163.367
R700 B.n369 B.n368 163.367
R701 B.n370 B.n369 163.367
R702 B.n370 B.n133 163.367
R703 B.n374 B.n133 163.367
R704 B.n375 B.n374 163.367
R705 B.n376 B.n375 163.367
R706 B.n376 B.n131 163.367
R707 B.n380 B.n131 163.367
R708 B.n381 B.n380 163.367
R709 B.n382 B.n381 163.367
R710 B.n382 B.n129 163.367
R711 B.n386 B.n129 163.367
R712 B.n387 B.n386 163.367
R713 B.n388 B.n127 163.367
R714 B.n392 B.n127 163.367
R715 B.n393 B.n392 163.367
R716 B.n394 B.n393 163.367
R717 B.n394 B.n125 163.367
R718 B.n398 B.n125 163.367
R719 B.n399 B.n398 163.367
R720 B.n400 B.n399 163.367
R721 B.n400 B.n123 163.367
R722 B.n404 B.n123 163.367
R723 B.n405 B.n404 163.367
R724 B.n406 B.n405 163.367
R725 B.n406 B.n121 163.367
R726 B.n410 B.n121 163.367
R727 B.n411 B.n410 163.367
R728 B.n412 B.n411 163.367
R729 B.n412 B.n119 163.367
R730 B.n416 B.n119 163.367
R731 B.n417 B.n416 163.367
R732 B.n418 B.n417 163.367
R733 B.n418 B.n117 163.367
R734 B.n422 B.n117 163.367
R735 B.n423 B.n422 163.367
R736 B.n424 B.n423 163.367
R737 B.n424 B.n115 163.367
R738 B.n428 B.n115 163.367
R739 B.n429 B.n428 163.367
R740 B.n430 B.n429 163.367
R741 B.n430 B.n113 163.367
R742 B.n434 B.n113 163.367
R743 B.n435 B.n434 163.367
R744 B.n436 B.n435 163.367
R745 B.n436 B.n111 163.367
R746 B.n440 B.n111 163.367
R747 B.n441 B.n440 163.367
R748 B.n442 B.n441 163.367
R749 B.n442 B.n109 163.367
R750 B.n446 B.n109 163.367
R751 B.n447 B.n446 163.367
R752 B.n448 B.n447 163.367
R753 B.n448 B.n107 163.367
R754 B.n452 B.n107 163.367
R755 B.n453 B.n452 163.367
R756 B.n454 B.n453 163.367
R757 B.n454 B.n105 163.367
R758 B.n458 B.n105 163.367
R759 B.n459 B.n458 163.367
R760 B.n460 B.n459 163.367
R761 B.n460 B.n103 163.367
R762 B.n464 B.n103 163.367
R763 B.n465 B.n464 163.367
R764 B.n466 B.n465 163.367
R765 B.n466 B.n101 163.367
R766 B.n470 B.n101 163.367
R767 B.n471 B.n470 163.367
R768 B.n472 B.n471 163.367
R769 B.n472 B.n99 163.367
R770 B.n476 B.n99 163.367
R771 B.n477 B.n476 163.367
R772 B.n478 B.n477 163.367
R773 B.n478 B.n97 163.367
R774 B.n482 B.n97 163.367
R775 B.n483 B.n482 163.367
R776 B.n484 B.n483 163.367
R777 B.n484 B.n95 163.367
R778 B.n488 B.n95 163.367
R779 B.n489 B.n488 163.367
R780 B.n490 B.n489 163.367
R781 B.n490 B.n93 163.367
R782 B.n494 B.n93 163.367
R783 B.n495 B.n494 163.367
R784 B.n496 B.n495 163.367
R785 B.n496 B.n91 163.367
R786 B.n500 B.n91 163.367
R787 B.n501 B.n500 163.367
R788 B.n502 B.n501 163.367
R789 B.n502 B.n89 163.367
R790 B.n506 B.n89 163.367
R791 B.n507 B.n506 163.367
R792 B.n508 B.n507 163.367
R793 B.n508 B.n87 163.367
R794 B.n512 B.n87 163.367
R795 B.n513 B.n512 163.367
R796 B.n514 B.n513 163.367
R797 B.n514 B.n85 163.367
R798 B.n518 B.n85 163.367
R799 B.n519 B.n518 163.367
R800 B.n520 B.n519 163.367
R801 B.n520 B.n83 163.367
R802 B.n524 B.n83 163.367
R803 B.n525 B.n524 163.367
R804 B.n526 B.n525 163.367
R805 B.n526 B.n81 163.367
R806 B.n530 B.n81 163.367
R807 B.n531 B.n530 163.367
R808 B.n532 B.n531 163.367
R809 B.n532 B.n79 163.367
R810 B.n536 B.n79 163.367
R811 B.n537 B.n536 163.367
R812 B.n538 B.n537 163.367
R813 B.n538 B.n77 163.367
R814 B.n542 B.n77 163.367
R815 B.n543 B.n542 163.367
R816 B.n544 B.n543 163.367
R817 B.n544 B.n75 163.367
R818 B.n548 B.n75 163.367
R819 B.n549 B.n548 163.367
R820 B.n550 B.n549 163.367
R821 B.n550 B.n73 163.367
R822 B.n554 B.n73 163.367
R823 B.n555 B.n554 163.367
R824 B.n556 B.n555 163.367
R825 B.n556 B.n71 163.367
R826 B.n560 B.n71 163.367
R827 B.n668 B.n31 163.367
R828 B.n664 B.n31 163.367
R829 B.n664 B.n663 163.367
R830 B.n663 B.n662 163.367
R831 B.n662 B.n33 163.367
R832 B.n658 B.n33 163.367
R833 B.n658 B.n657 163.367
R834 B.n657 B.n656 163.367
R835 B.n656 B.n35 163.367
R836 B.n652 B.n35 163.367
R837 B.n652 B.n651 163.367
R838 B.n651 B.n650 163.367
R839 B.n650 B.n37 163.367
R840 B.n646 B.n37 163.367
R841 B.n646 B.n645 163.367
R842 B.n645 B.n644 163.367
R843 B.n644 B.n39 163.367
R844 B.n640 B.n39 163.367
R845 B.n640 B.n639 163.367
R846 B.n639 B.n638 163.367
R847 B.n638 B.n41 163.367
R848 B.n634 B.n41 163.367
R849 B.n634 B.n633 163.367
R850 B.n633 B.n632 163.367
R851 B.n632 B.n43 163.367
R852 B.n628 B.n43 163.367
R853 B.n628 B.n627 163.367
R854 B.n627 B.n626 163.367
R855 B.n626 B.n45 163.367
R856 B.n622 B.n45 163.367
R857 B.n622 B.n621 163.367
R858 B.n621 B.n49 163.367
R859 B.n617 B.n49 163.367
R860 B.n617 B.n616 163.367
R861 B.n616 B.n615 163.367
R862 B.n615 B.n51 163.367
R863 B.n611 B.n51 163.367
R864 B.n611 B.n610 163.367
R865 B.n610 B.n609 163.367
R866 B.n609 B.n53 163.367
R867 B.n604 B.n53 163.367
R868 B.n604 B.n603 163.367
R869 B.n603 B.n602 163.367
R870 B.n602 B.n57 163.367
R871 B.n598 B.n57 163.367
R872 B.n598 B.n597 163.367
R873 B.n597 B.n596 163.367
R874 B.n596 B.n59 163.367
R875 B.n592 B.n59 163.367
R876 B.n592 B.n591 163.367
R877 B.n591 B.n590 163.367
R878 B.n590 B.n61 163.367
R879 B.n586 B.n61 163.367
R880 B.n586 B.n585 163.367
R881 B.n585 B.n584 163.367
R882 B.n584 B.n63 163.367
R883 B.n580 B.n63 163.367
R884 B.n580 B.n579 163.367
R885 B.n579 B.n578 163.367
R886 B.n578 B.n65 163.367
R887 B.n574 B.n65 163.367
R888 B.n574 B.n573 163.367
R889 B.n573 B.n572 163.367
R890 B.n572 B.n67 163.367
R891 B.n568 B.n67 163.367
R892 B.n568 B.n567 163.367
R893 B.n567 B.n566 163.367
R894 B.n566 B.n69 163.367
R895 B.n562 B.n69 163.367
R896 B.n562 B.n561 163.367
R897 B.n145 B.t1 112.329
R898 B.n55 B.t8 112.329
R899 B.n151 B.t4 112.32
R900 B.n47 B.t11 112.32
R901 B.n145 B.n144 64.5823
R902 B.n151 B.n150 64.5823
R903 B.n47 B.n46 64.5823
R904 B.n55 B.n54 64.5823
R905 B.n341 B.n145 59.5399
R906 B.n152 B.n151 59.5399
R907 B.n48 B.n47 59.5399
R908 B.n607 B.n55 59.5399
R909 B.n667 B.n30 35.4346
R910 B.n389 B.n128 35.4346
R911 B.n281 B.n168 35.4346
R912 B.n559 B.n70 35.4346
R913 B B.n755 18.0485
R914 B.n667 B.n666 10.6151
R915 B.n666 B.n665 10.6151
R916 B.n665 B.n32 10.6151
R917 B.n661 B.n32 10.6151
R918 B.n661 B.n660 10.6151
R919 B.n660 B.n659 10.6151
R920 B.n659 B.n34 10.6151
R921 B.n655 B.n34 10.6151
R922 B.n655 B.n654 10.6151
R923 B.n654 B.n653 10.6151
R924 B.n653 B.n36 10.6151
R925 B.n649 B.n36 10.6151
R926 B.n649 B.n648 10.6151
R927 B.n648 B.n647 10.6151
R928 B.n647 B.n38 10.6151
R929 B.n643 B.n38 10.6151
R930 B.n643 B.n642 10.6151
R931 B.n642 B.n641 10.6151
R932 B.n641 B.n40 10.6151
R933 B.n637 B.n40 10.6151
R934 B.n637 B.n636 10.6151
R935 B.n636 B.n635 10.6151
R936 B.n635 B.n42 10.6151
R937 B.n631 B.n42 10.6151
R938 B.n631 B.n630 10.6151
R939 B.n630 B.n629 10.6151
R940 B.n629 B.n44 10.6151
R941 B.n625 B.n44 10.6151
R942 B.n625 B.n624 10.6151
R943 B.n624 B.n623 10.6151
R944 B.n620 B.n619 10.6151
R945 B.n619 B.n618 10.6151
R946 B.n618 B.n50 10.6151
R947 B.n614 B.n50 10.6151
R948 B.n614 B.n613 10.6151
R949 B.n613 B.n612 10.6151
R950 B.n612 B.n52 10.6151
R951 B.n608 B.n52 10.6151
R952 B.n606 B.n605 10.6151
R953 B.n605 B.n56 10.6151
R954 B.n601 B.n56 10.6151
R955 B.n601 B.n600 10.6151
R956 B.n600 B.n599 10.6151
R957 B.n599 B.n58 10.6151
R958 B.n595 B.n58 10.6151
R959 B.n595 B.n594 10.6151
R960 B.n594 B.n593 10.6151
R961 B.n593 B.n60 10.6151
R962 B.n589 B.n60 10.6151
R963 B.n589 B.n588 10.6151
R964 B.n588 B.n587 10.6151
R965 B.n587 B.n62 10.6151
R966 B.n583 B.n62 10.6151
R967 B.n583 B.n582 10.6151
R968 B.n582 B.n581 10.6151
R969 B.n581 B.n64 10.6151
R970 B.n577 B.n64 10.6151
R971 B.n577 B.n576 10.6151
R972 B.n576 B.n575 10.6151
R973 B.n575 B.n66 10.6151
R974 B.n571 B.n66 10.6151
R975 B.n571 B.n570 10.6151
R976 B.n570 B.n569 10.6151
R977 B.n569 B.n68 10.6151
R978 B.n565 B.n68 10.6151
R979 B.n565 B.n564 10.6151
R980 B.n564 B.n563 10.6151
R981 B.n563 B.n70 10.6151
R982 B.n390 B.n389 10.6151
R983 B.n391 B.n390 10.6151
R984 B.n391 B.n126 10.6151
R985 B.n395 B.n126 10.6151
R986 B.n396 B.n395 10.6151
R987 B.n397 B.n396 10.6151
R988 B.n397 B.n124 10.6151
R989 B.n401 B.n124 10.6151
R990 B.n402 B.n401 10.6151
R991 B.n403 B.n402 10.6151
R992 B.n403 B.n122 10.6151
R993 B.n407 B.n122 10.6151
R994 B.n408 B.n407 10.6151
R995 B.n409 B.n408 10.6151
R996 B.n409 B.n120 10.6151
R997 B.n413 B.n120 10.6151
R998 B.n414 B.n413 10.6151
R999 B.n415 B.n414 10.6151
R1000 B.n415 B.n118 10.6151
R1001 B.n419 B.n118 10.6151
R1002 B.n420 B.n419 10.6151
R1003 B.n421 B.n420 10.6151
R1004 B.n421 B.n116 10.6151
R1005 B.n425 B.n116 10.6151
R1006 B.n426 B.n425 10.6151
R1007 B.n427 B.n426 10.6151
R1008 B.n427 B.n114 10.6151
R1009 B.n431 B.n114 10.6151
R1010 B.n432 B.n431 10.6151
R1011 B.n433 B.n432 10.6151
R1012 B.n433 B.n112 10.6151
R1013 B.n437 B.n112 10.6151
R1014 B.n438 B.n437 10.6151
R1015 B.n439 B.n438 10.6151
R1016 B.n439 B.n110 10.6151
R1017 B.n443 B.n110 10.6151
R1018 B.n444 B.n443 10.6151
R1019 B.n445 B.n444 10.6151
R1020 B.n445 B.n108 10.6151
R1021 B.n449 B.n108 10.6151
R1022 B.n450 B.n449 10.6151
R1023 B.n451 B.n450 10.6151
R1024 B.n451 B.n106 10.6151
R1025 B.n455 B.n106 10.6151
R1026 B.n456 B.n455 10.6151
R1027 B.n457 B.n456 10.6151
R1028 B.n457 B.n104 10.6151
R1029 B.n461 B.n104 10.6151
R1030 B.n462 B.n461 10.6151
R1031 B.n463 B.n462 10.6151
R1032 B.n463 B.n102 10.6151
R1033 B.n467 B.n102 10.6151
R1034 B.n468 B.n467 10.6151
R1035 B.n469 B.n468 10.6151
R1036 B.n469 B.n100 10.6151
R1037 B.n473 B.n100 10.6151
R1038 B.n474 B.n473 10.6151
R1039 B.n475 B.n474 10.6151
R1040 B.n475 B.n98 10.6151
R1041 B.n479 B.n98 10.6151
R1042 B.n480 B.n479 10.6151
R1043 B.n481 B.n480 10.6151
R1044 B.n481 B.n96 10.6151
R1045 B.n485 B.n96 10.6151
R1046 B.n486 B.n485 10.6151
R1047 B.n487 B.n486 10.6151
R1048 B.n487 B.n94 10.6151
R1049 B.n491 B.n94 10.6151
R1050 B.n492 B.n491 10.6151
R1051 B.n493 B.n492 10.6151
R1052 B.n493 B.n92 10.6151
R1053 B.n497 B.n92 10.6151
R1054 B.n498 B.n497 10.6151
R1055 B.n499 B.n498 10.6151
R1056 B.n499 B.n90 10.6151
R1057 B.n503 B.n90 10.6151
R1058 B.n504 B.n503 10.6151
R1059 B.n505 B.n504 10.6151
R1060 B.n505 B.n88 10.6151
R1061 B.n509 B.n88 10.6151
R1062 B.n510 B.n509 10.6151
R1063 B.n511 B.n510 10.6151
R1064 B.n511 B.n86 10.6151
R1065 B.n515 B.n86 10.6151
R1066 B.n516 B.n515 10.6151
R1067 B.n517 B.n516 10.6151
R1068 B.n517 B.n84 10.6151
R1069 B.n521 B.n84 10.6151
R1070 B.n522 B.n521 10.6151
R1071 B.n523 B.n522 10.6151
R1072 B.n523 B.n82 10.6151
R1073 B.n527 B.n82 10.6151
R1074 B.n528 B.n527 10.6151
R1075 B.n529 B.n528 10.6151
R1076 B.n529 B.n80 10.6151
R1077 B.n533 B.n80 10.6151
R1078 B.n534 B.n533 10.6151
R1079 B.n535 B.n534 10.6151
R1080 B.n535 B.n78 10.6151
R1081 B.n539 B.n78 10.6151
R1082 B.n540 B.n539 10.6151
R1083 B.n541 B.n540 10.6151
R1084 B.n541 B.n76 10.6151
R1085 B.n545 B.n76 10.6151
R1086 B.n546 B.n545 10.6151
R1087 B.n547 B.n546 10.6151
R1088 B.n547 B.n74 10.6151
R1089 B.n551 B.n74 10.6151
R1090 B.n552 B.n551 10.6151
R1091 B.n553 B.n552 10.6151
R1092 B.n553 B.n72 10.6151
R1093 B.n557 B.n72 10.6151
R1094 B.n558 B.n557 10.6151
R1095 B.n559 B.n558 10.6151
R1096 B.n282 B.n281 10.6151
R1097 B.n283 B.n282 10.6151
R1098 B.n283 B.n166 10.6151
R1099 B.n287 B.n166 10.6151
R1100 B.n288 B.n287 10.6151
R1101 B.n289 B.n288 10.6151
R1102 B.n289 B.n164 10.6151
R1103 B.n293 B.n164 10.6151
R1104 B.n294 B.n293 10.6151
R1105 B.n295 B.n294 10.6151
R1106 B.n295 B.n162 10.6151
R1107 B.n299 B.n162 10.6151
R1108 B.n300 B.n299 10.6151
R1109 B.n301 B.n300 10.6151
R1110 B.n301 B.n160 10.6151
R1111 B.n305 B.n160 10.6151
R1112 B.n306 B.n305 10.6151
R1113 B.n307 B.n306 10.6151
R1114 B.n307 B.n158 10.6151
R1115 B.n311 B.n158 10.6151
R1116 B.n312 B.n311 10.6151
R1117 B.n313 B.n312 10.6151
R1118 B.n313 B.n156 10.6151
R1119 B.n317 B.n156 10.6151
R1120 B.n318 B.n317 10.6151
R1121 B.n319 B.n318 10.6151
R1122 B.n319 B.n154 10.6151
R1123 B.n323 B.n154 10.6151
R1124 B.n324 B.n323 10.6151
R1125 B.n325 B.n324 10.6151
R1126 B.n329 B.n328 10.6151
R1127 B.n330 B.n329 10.6151
R1128 B.n330 B.n148 10.6151
R1129 B.n334 B.n148 10.6151
R1130 B.n335 B.n334 10.6151
R1131 B.n336 B.n335 10.6151
R1132 B.n336 B.n146 10.6151
R1133 B.n340 B.n146 10.6151
R1134 B.n343 B.n342 10.6151
R1135 B.n343 B.n142 10.6151
R1136 B.n347 B.n142 10.6151
R1137 B.n348 B.n347 10.6151
R1138 B.n349 B.n348 10.6151
R1139 B.n349 B.n140 10.6151
R1140 B.n353 B.n140 10.6151
R1141 B.n354 B.n353 10.6151
R1142 B.n355 B.n354 10.6151
R1143 B.n355 B.n138 10.6151
R1144 B.n359 B.n138 10.6151
R1145 B.n360 B.n359 10.6151
R1146 B.n361 B.n360 10.6151
R1147 B.n361 B.n136 10.6151
R1148 B.n365 B.n136 10.6151
R1149 B.n366 B.n365 10.6151
R1150 B.n367 B.n366 10.6151
R1151 B.n367 B.n134 10.6151
R1152 B.n371 B.n134 10.6151
R1153 B.n372 B.n371 10.6151
R1154 B.n373 B.n372 10.6151
R1155 B.n373 B.n132 10.6151
R1156 B.n377 B.n132 10.6151
R1157 B.n378 B.n377 10.6151
R1158 B.n379 B.n378 10.6151
R1159 B.n379 B.n130 10.6151
R1160 B.n383 B.n130 10.6151
R1161 B.n384 B.n383 10.6151
R1162 B.n385 B.n384 10.6151
R1163 B.n385 B.n128 10.6151
R1164 B.n277 B.n168 10.6151
R1165 B.n277 B.n276 10.6151
R1166 B.n276 B.n275 10.6151
R1167 B.n275 B.n170 10.6151
R1168 B.n271 B.n170 10.6151
R1169 B.n271 B.n270 10.6151
R1170 B.n270 B.n269 10.6151
R1171 B.n269 B.n172 10.6151
R1172 B.n265 B.n172 10.6151
R1173 B.n265 B.n264 10.6151
R1174 B.n264 B.n263 10.6151
R1175 B.n263 B.n174 10.6151
R1176 B.n259 B.n174 10.6151
R1177 B.n259 B.n258 10.6151
R1178 B.n258 B.n257 10.6151
R1179 B.n257 B.n176 10.6151
R1180 B.n253 B.n176 10.6151
R1181 B.n253 B.n252 10.6151
R1182 B.n252 B.n251 10.6151
R1183 B.n251 B.n178 10.6151
R1184 B.n247 B.n178 10.6151
R1185 B.n247 B.n246 10.6151
R1186 B.n246 B.n245 10.6151
R1187 B.n245 B.n180 10.6151
R1188 B.n241 B.n180 10.6151
R1189 B.n241 B.n240 10.6151
R1190 B.n240 B.n239 10.6151
R1191 B.n239 B.n182 10.6151
R1192 B.n235 B.n182 10.6151
R1193 B.n235 B.n234 10.6151
R1194 B.n234 B.n233 10.6151
R1195 B.n233 B.n184 10.6151
R1196 B.n229 B.n184 10.6151
R1197 B.n229 B.n228 10.6151
R1198 B.n228 B.n227 10.6151
R1199 B.n227 B.n186 10.6151
R1200 B.n223 B.n186 10.6151
R1201 B.n223 B.n222 10.6151
R1202 B.n222 B.n221 10.6151
R1203 B.n221 B.n188 10.6151
R1204 B.n217 B.n188 10.6151
R1205 B.n217 B.n216 10.6151
R1206 B.n216 B.n215 10.6151
R1207 B.n215 B.n190 10.6151
R1208 B.n211 B.n190 10.6151
R1209 B.n211 B.n210 10.6151
R1210 B.n210 B.n209 10.6151
R1211 B.n209 B.n192 10.6151
R1212 B.n205 B.n192 10.6151
R1213 B.n205 B.n204 10.6151
R1214 B.n204 B.n203 10.6151
R1215 B.n203 B.n194 10.6151
R1216 B.n199 B.n194 10.6151
R1217 B.n199 B.n198 10.6151
R1218 B.n198 B.n197 10.6151
R1219 B.n197 B.n0 10.6151
R1220 B.n751 B.n1 10.6151
R1221 B.n751 B.n750 10.6151
R1222 B.n750 B.n749 10.6151
R1223 B.n749 B.n4 10.6151
R1224 B.n745 B.n4 10.6151
R1225 B.n745 B.n744 10.6151
R1226 B.n744 B.n743 10.6151
R1227 B.n743 B.n6 10.6151
R1228 B.n739 B.n6 10.6151
R1229 B.n739 B.n738 10.6151
R1230 B.n738 B.n737 10.6151
R1231 B.n737 B.n8 10.6151
R1232 B.n733 B.n8 10.6151
R1233 B.n733 B.n732 10.6151
R1234 B.n732 B.n731 10.6151
R1235 B.n731 B.n10 10.6151
R1236 B.n727 B.n10 10.6151
R1237 B.n727 B.n726 10.6151
R1238 B.n726 B.n725 10.6151
R1239 B.n725 B.n12 10.6151
R1240 B.n721 B.n12 10.6151
R1241 B.n721 B.n720 10.6151
R1242 B.n720 B.n719 10.6151
R1243 B.n719 B.n14 10.6151
R1244 B.n715 B.n14 10.6151
R1245 B.n715 B.n714 10.6151
R1246 B.n714 B.n713 10.6151
R1247 B.n713 B.n16 10.6151
R1248 B.n709 B.n16 10.6151
R1249 B.n709 B.n708 10.6151
R1250 B.n708 B.n707 10.6151
R1251 B.n707 B.n18 10.6151
R1252 B.n703 B.n18 10.6151
R1253 B.n703 B.n702 10.6151
R1254 B.n702 B.n701 10.6151
R1255 B.n701 B.n20 10.6151
R1256 B.n697 B.n20 10.6151
R1257 B.n697 B.n696 10.6151
R1258 B.n696 B.n695 10.6151
R1259 B.n695 B.n22 10.6151
R1260 B.n691 B.n22 10.6151
R1261 B.n691 B.n690 10.6151
R1262 B.n690 B.n689 10.6151
R1263 B.n689 B.n24 10.6151
R1264 B.n685 B.n24 10.6151
R1265 B.n685 B.n684 10.6151
R1266 B.n684 B.n683 10.6151
R1267 B.n683 B.n26 10.6151
R1268 B.n679 B.n26 10.6151
R1269 B.n679 B.n678 10.6151
R1270 B.n678 B.n677 10.6151
R1271 B.n677 B.n28 10.6151
R1272 B.n673 B.n28 10.6151
R1273 B.n673 B.n672 10.6151
R1274 B.n672 B.n671 10.6151
R1275 B.n671 B.n30 10.6151
R1276 B.n620 B.n48 6.5566
R1277 B.n608 B.n607 6.5566
R1278 B.n328 B.n152 6.5566
R1279 B.n341 B.n340 6.5566
R1280 B.n623 B.n48 4.05904
R1281 B.n607 B.n606 4.05904
R1282 B.n325 B.n152 4.05904
R1283 B.n342 B.n341 4.05904
R1284 B.n755 B.n0 2.81026
R1285 B.n755 B.n1 2.81026
R1286 VP.n21 VP.n20 161.3
R1287 VP.n22 VP.n17 161.3
R1288 VP.n24 VP.n23 161.3
R1289 VP.n25 VP.n16 161.3
R1290 VP.n27 VP.n26 161.3
R1291 VP.n28 VP.n15 161.3
R1292 VP.n30 VP.n29 161.3
R1293 VP.n32 VP.n14 161.3
R1294 VP.n34 VP.n33 161.3
R1295 VP.n35 VP.n13 161.3
R1296 VP.n37 VP.n36 161.3
R1297 VP.n38 VP.n12 161.3
R1298 VP.n40 VP.n39 161.3
R1299 VP.n73 VP.n72 161.3
R1300 VP.n71 VP.n1 161.3
R1301 VP.n70 VP.n69 161.3
R1302 VP.n68 VP.n2 161.3
R1303 VP.n67 VP.n66 161.3
R1304 VP.n65 VP.n3 161.3
R1305 VP.n63 VP.n62 161.3
R1306 VP.n61 VP.n4 161.3
R1307 VP.n60 VP.n59 161.3
R1308 VP.n58 VP.n5 161.3
R1309 VP.n57 VP.n56 161.3
R1310 VP.n55 VP.n6 161.3
R1311 VP.n54 VP.n53 161.3
R1312 VP.n51 VP.n7 161.3
R1313 VP.n50 VP.n49 161.3
R1314 VP.n48 VP.n8 161.3
R1315 VP.n47 VP.n46 161.3
R1316 VP.n45 VP.n9 161.3
R1317 VP.n44 VP.n43 161.3
R1318 VP.n18 VP.t2 98.9902
R1319 VP.n10 VP.t6 67.1592
R1320 VP.n52 VP.t3 67.1592
R1321 VP.n64 VP.t7 67.1592
R1322 VP.n0 VP.t0 67.1592
R1323 VP.n11 VP.t4 67.1592
R1324 VP.n31 VP.t5 67.1592
R1325 VP.n19 VP.t1 67.1592
R1326 VP.n19 VP.n18 66.0722
R1327 VP.n42 VP.n10 65.8996
R1328 VP.n74 VP.n0 65.8996
R1329 VP.n41 VP.n11 65.8996
R1330 VP.n46 VP.n8 56.5617
R1331 VP.n70 VP.n2 56.5617
R1332 VP.n37 VP.n13 56.5617
R1333 VP.n42 VP.n41 50.1965
R1334 VP.n58 VP.n57 40.577
R1335 VP.n59 VP.n58 40.577
R1336 VP.n26 VP.n25 40.577
R1337 VP.n25 VP.n24 40.577
R1338 VP.n45 VP.n44 24.5923
R1339 VP.n46 VP.n45 24.5923
R1340 VP.n50 VP.n8 24.5923
R1341 VP.n51 VP.n50 24.5923
R1342 VP.n53 VP.n6 24.5923
R1343 VP.n57 VP.n6 24.5923
R1344 VP.n59 VP.n4 24.5923
R1345 VP.n63 VP.n4 24.5923
R1346 VP.n66 VP.n65 24.5923
R1347 VP.n66 VP.n2 24.5923
R1348 VP.n71 VP.n70 24.5923
R1349 VP.n72 VP.n71 24.5923
R1350 VP.n38 VP.n37 24.5923
R1351 VP.n39 VP.n38 24.5923
R1352 VP.n26 VP.n15 24.5923
R1353 VP.n30 VP.n15 24.5923
R1354 VP.n33 VP.n32 24.5923
R1355 VP.n33 VP.n13 24.5923
R1356 VP.n20 VP.n17 24.5923
R1357 VP.n24 VP.n17 24.5923
R1358 VP.n44 VP.n10 24.3464
R1359 VP.n72 VP.n0 24.3464
R1360 VP.n39 VP.n11 24.3464
R1361 VP.n52 VP.n51 16.477
R1362 VP.n65 VP.n64 16.477
R1363 VP.n32 VP.n31 16.477
R1364 VP.n53 VP.n52 8.11581
R1365 VP.n64 VP.n63 8.11581
R1366 VP.n31 VP.n30 8.11581
R1367 VP.n20 VP.n19 8.11581
R1368 VP.n21 VP.n18 5.23308
R1369 VP.n41 VP.n40 0.354861
R1370 VP.n43 VP.n42 0.354861
R1371 VP.n74 VP.n73 0.354861
R1372 VP VP.n74 0.267071
R1373 VP.n22 VP.n21 0.189894
R1374 VP.n23 VP.n22 0.189894
R1375 VP.n23 VP.n16 0.189894
R1376 VP.n27 VP.n16 0.189894
R1377 VP.n28 VP.n27 0.189894
R1378 VP.n29 VP.n28 0.189894
R1379 VP.n29 VP.n14 0.189894
R1380 VP.n34 VP.n14 0.189894
R1381 VP.n35 VP.n34 0.189894
R1382 VP.n36 VP.n35 0.189894
R1383 VP.n36 VP.n12 0.189894
R1384 VP.n40 VP.n12 0.189894
R1385 VP.n43 VP.n9 0.189894
R1386 VP.n47 VP.n9 0.189894
R1387 VP.n48 VP.n47 0.189894
R1388 VP.n49 VP.n48 0.189894
R1389 VP.n49 VP.n7 0.189894
R1390 VP.n54 VP.n7 0.189894
R1391 VP.n55 VP.n54 0.189894
R1392 VP.n56 VP.n55 0.189894
R1393 VP.n56 VP.n5 0.189894
R1394 VP.n60 VP.n5 0.189894
R1395 VP.n61 VP.n60 0.189894
R1396 VP.n62 VP.n61 0.189894
R1397 VP.n62 VP.n3 0.189894
R1398 VP.n67 VP.n3 0.189894
R1399 VP.n68 VP.n67 0.189894
R1400 VP.n69 VP.n68 0.189894
R1401 VP.n69 VP.n1 0.189894
R1402 VP.n73 VP.n1 0.189894
R1403 VDD1 VDD1.n0 86.6572
R1404 VDD1.n3 VDD1.n2 86.5434
R1405 VDD1.n3 VDD1.n1 86.5434
R1406 VDD1.n5 VDD1.n4 85.1635
R1407 VDD1.n5 VDD1.n3 44.4233
R1408 VDD1.n4 VDD1.t2 3.88866
R1409 VDD1.n4 VDD1.t3 3.88866
R1410 VDD1.n0 VDD1.t5 3.88866
R1411 VDD1.n0 VDD1.t6 3.88866
R1412 VDD1.n2 VDD1.t0 3.88866
R1413 VDD1.n2 VDD1.t7 3.88866
R1414 VDD1.n1 VDD1.t1 3.88866
R1415 VDD1.n1 VDD1.t4 3.88866
R1416 VDD1 VDD1.n5 1.37766
C0 B VDD2 1.78136f
C1 VDD1 B 1.67275f
C2 VDD1 VDD2 1.98659f
C3 w_n4300_n2640# VN 8.78036f
C4 VN VP 7.4706f
C5 w_n4300_n2640# VP 9.339769f
C6 VTAIL VN 7.05774f
C7 w_n4300_n2640# VTAIL 3.42919f
C8 VTAIL VP 7.07185f
C9 VN B 1.27967f
C10 w_n4300_n2640# B 9.70764f
C11 B VP 2.21956f
C12 VN VDD2 6.35126f
C13 VDD1 VN 0.152903f
C14 w_n4300_n2640# VDD2 2.12035f
C15 w_n4300_n2640# VDD1 1.98886f
C16 VP VDD2 0.562687f
C17 VDD1 VP 6.75945f
C18 VTAIL B 3.93817f
C19 VTAIL VDD2 7.11567f
C20 VDD1 VTAIL 7.05857f
C21 VDD2 VSUBS 1.907411f
C22 VDD1 VSUBS 2.489123f
C23 VTAIL VSUBS 1.255376f
C24 VN VSUBS 7.22556f
C25 VP VSUBS 3.885092f
C26 B VSUBS 5.14383f
C27 w_n4300_n2640# VSUBS 0.140713p
C28 VDD1.t5 VSUBS 0.163544f
C29 VDD1.t6 VSUBS 0.163544f
C30 VDD1.n0 VSUBS 1.21277f
C31 VDD1.t1 VSUBS 0.163544f
C32 VDD1.t4 VSUBS 0.163544f
C33 VDD1.n1 VSUBS 1.21163f
C34 VDD1.t0 VSUBS 0.163544f
C35 VDD1.t7 VSUBS 0.163544f
C36 VDD1.n2 VSUBS 1.21163f
C37 VDD1.n3 VSUBS 3.73353f
C38 VDD1.t2 VSUBS 0.163544f
C39 VDD1.t3 VSUBS 0.163544f
C40 VDD1.n4 VSUBS 1.19936f
C41 VDD1.n5 VSUBS 3.02926f
C42 VP.t0 VSUBS 2.27459f
C43 VP.n0 VSUBS 0.963238f
C44 VP.n1 VSUBS 0.033706f
C45 VP.n2 VSUBS 0.056457f
C46 VP.n3 VSUBS 0.033706f
C47 VP.t7 VSUBS 2.27459f
C48 VP.n4 VSUBS 0.062505f
C49 VP.n5 VSUBS 0.033706f
C50 VP.n6 VSUBS 0.062505f
C51 VP.n7 VSUBS 0.033706f
C52 VP.t3 VSUBS 2.27459f
C53 VP.n8 VSUBS 0.056457f
C54 VP.n9 VSUBS 0.033706f
C55 VP.t6 VSUBS 2.27459f
C56 VP.n10 VSUBS 0.963238f
C57 VP.t4 VSUBS 2.27459f
C58 VP.n11 VSUBS 0.963238f
C59 VP.n12 VSUBS 0.033706f
C60 VP.n13 VSUBS 0.056457f
C61 VP.n14 VSUBS 0.033706f
C62 VP.t5 VSUBS 2.27459f
C63 VP.n15 VSUBS 0.062505f
C64 VP.n16 VSUBS 0.033706f
C65 VP.n17 VSUBS 0.062505f
C66 VP.t2 VSUBS 2.61274f
C67 VP.n18 VSUBS 0.89123f
C68 VP.t1 VSUBS 2.27459f
C69 VP.n19 VSUBS 0.92223f
C70 VP.n20 VSUBS 0.04183f
C71 VP.n21 VSUBS 0.361433f
C72 VP.n22 VSUBS 0.033706f
C73 VP.n23 VSUBS 0.033706f
C74 VP.n24 VSUBS 0.066637f
C75 VP.n25 VSUBS 0.027223f
C76 VP.n26 VSUBS 0.066637f
C77 VP.n27 VSUBS 0.033706f
C78 VP.n28 VSUBS 0.033706f
C79 VP.n29 VSUBS 0.033706f
C80 VP.n30 VSUBS 0.04183f
C81 VP.n31 VSUBS 0.82054f
C82 VP.n32 VSUBS 0.052322f
C83 VP.n33 VSUBS 0.062505f
C84 VP.n34 VSUBS 0.033706f
C85 VP.n35 VSUBS 0.033706f
C86 VP.n36 VSUBS 0.033706f
C87 VP.n37 VSUBS 0.041536f
C88 VP.n38 VSUBS 0.062505f
C89 VP.n39 VSUBS 0.062196f
C90 VP.n40 VSUBS 0.054392f
C91 VP.n41 VSUBS 1.91087f
C92 VP.n42 VSUBS 1.93508f
C93 VP.n43 VSUBS 0.054392f
C94 VP.n44 VSUBS 0.062196f
C95 VP.n45 VSUBS 0.062505f
C96 VP.n46 VSUBS 0.041536f
C97 VP.n47 VSUBS 0.033706f
C98 VP.n48 VSUBS 0.033706f
C99 VP.n49 VSUBS 0.033706f
C100 VP.n50 VSUBS 0.062505f
C101 VP.n51 VSUBS 0.052322f
C102 VP.n52 VSUBS 0.82054f
C103 VP.n53 VSUBS 0.04183f
C104 VP.n54 VSUBS 0.033706f
C105 VP.n55 VSUBS 0.033706f
C106 VP.n56 VSUBS 0.033706f
C107 VP.n57 VSUBS 0.066637f
C108 VP.n58 VSUBS 0.027223f
C109 VP.n59 VSUBS 0.066637f
C110 VP.n60 VSUBS 0.033706f
C111 VP.n61 VSUBS 0.033706f
C112 VP.n62 VSUBS 0.033706f
C113 VP.n63 VSUBS 0.04183f
C114 VP.n64 VSUBS 0.82054f
C115 VP.n65 VSUBS 0.052322f
C116 VP.n66 VSUBS 0.062505f
C117 VP.n67 VSUBS 0.033706f
C118 VP.n68 VSUBS 0.033706f
C119 VP.n69 VSUBS 0.033706f
C120 VP.n70 VSUBS 0.041536f
C121 VP.n71 VSUBS 0.062505f
C122 VP.n72 VSUBS 0.062196f
C123 VP.n73 VSUBS 0.054392f
C124 VP.n74 VSUBS 0.063029f
C125 B.n0 VSUBS 0.005287f
C126 B.n1 VSUBS 0.005287f
C127 B.n2 VSUBS 0.00836f
C128 B.n3 VSUBS 0.00836f
C129 B.n4 VSUBS 0.00836f
C130 B.n5 VSUBS 0.00836f
C131 B.n6 VSUBS 0.00836f
C132 B.n7 VSUBS 0.00836f
C133 B.n8 VSUBS 0.00836f
C134 B.n9 VSUBS 0.00836f
C135 B.n10 VSUBS 0.00836f
C136 B.n11 VSUBS 0.00836f
C137 B.n12 VSUBS 0.00836f
C138 B.n13 VSUBS 0.00836f
C139 B.n14 VSUBS 0.00836f
C140 B.n15 VSUBS 0.00836f
C141 B.n16 VSUBS 0.00836f
C142 B.n17 VSUBS 0.00836f
C143 B.n18 VSUBS 0.00836f
C144 B.n19 VSUBS 0.00836f
C145 B.n20 VSUBS 0.00836f
C146 B.n21 VSUBS 0.00836f
C147 B.n22 VSUBS 0.00836f
C148 B.n23 VSUBS 0.00836f
C149 B.n24 VSUBS 0.00836f
C150 B.n25 VSUBS 0.00836f
C151 B.n26 VSUBS 0.00836f
C152 B.n27 VSUBS 0.00836f
C153 B.n28 VSUBS 0.00836f
C154 B.n29 VSUBS 0.00836f
C155 B.n30 VSUBS 0.02031f
C156 B.n31 VSUBS 0.00836f
C157 B.n32 VSUBS 0.00836f
C158 B.n33 VSUBS 0.00836f
C159 B.n34 VSUBS 0.00836f
C160 B.n35 VSUBS 0.00836f
C161 B.n36 VSUBS 0.00836f
C162 B.n37 VSUBS 0.00836f
C163 B.n38 VSUBS 0.00836f
C164 B.n39 VSUBS 0.00836f
C165 B.n40 VSUBS 0.00836f
C166 B.n41 VSUBS 0.00836f
C167 B.n42 VSUBS 0.00836f
C168 B.n43 VSUBS 0.00836f
C169 B.n44 VSUBS 0.00836f
C170 B.n45 VSUBS 0.00836f
C171 B.t11 VSUBS 0.310278f
C172 B.t10 VSUBS 0.337804f
C173 B.t9 VSUBS 1.40453f
C174 B.n46 VSUBS 0.186944f
C175 B.n47 VSUBS 0.087325f
C176 B.n48 VSUBS 0.01937f
C177 B.n49 VSUBS 0.00836f
C178 B.n50 VSUBS 0.00836f
C179 B.n51 VSUBS 0.00836f
C180 B.n52 VSUBS 0.00836f
C181 B.n53 VSUBS 0.00836f
C182 B.t8 VSUBS 0.310275f
C183 B.t7 VSUBS 0.337801f
C184 B.t6 VSUBS 1.40453f
C185 B.n54 VSUBS 0.186948f
C186 B.n55 VSUBS 0.087327f
C187 B.n56 VSUBS 0.00836f
C188 B.n57 VSUBS 0.00836f
C189 B.n58 VSUBS 0.00836f
C190 B.n59 VSUBS 0.00836f
C191 B.n60 VSUBS 0.00836f
C192 B.n61 VSUBS 0.00836f
C193 B.n62 VSUBS 0.00836f
C194 B.n63 VSUBS 0.00836f
C195 B.n64 VSUBS 0.00836f
C196 B.n65 VSUBS 0.00836f
C197 B.n66 VSUBS 0.00836f
C198 B.n67 VSUBS 0.00836f
C199 B.n68 VSUBS 0.00836f
C200 B.n69 VSUBS 0.00836f
C201 B.n70 VSUBS 0.020088f
C202 B.n71 VSUBS 0.00836f
C203 B.n72 VSUBS 0.00836f
C204 B.n73 VSUBS 0.00836f
C205 B.n74 VSUBS 0.00836f
C206 B.n75 VSUBS 0.00836f
C207 B.n76 VSUBS 0.00836f
C208 B.n77 VSUBS 0.00836f
C209 B.n78 VSUBS 0.00836f
C210 B.n79 VSUBS 0.00836f
C211 B.n80 VSUBS 0.00836f
C212 B.n81 VSUBS 0.00836f
C213 B.n82 VSUBS 0.00836f
C214 B.n83 VSUBS 0.00836f
C215 B.n84 VSUBS 0.00836f
C216 B.n85 VSUBS 0.00836f
C217 B.n86 VSUBS 0.00836f
C218 B.n87 VSUBS 0.00836f
C219 B.n88 VSUBS 0.00836f
C220 B.n89 VSUBS 0.00836f
C221 B.n90 VSUBS 0.00836f
C222 B.n91 VSUBS 0.00836f
C223 B.n92 VSUBS 0.00836f
C224 B.n93 VSUBS 0.00836f
C225 B.n94 VSUBS 0.00836f
C226 B.n95 VSUBS 0.00836f
C227 B.n96 VSUBS 0.00836f
C228 B.n97 VSUBS 0.00836f
C229 B.n98 VSUBS 0.00836f
C230 B.n99 VSUBS 0.00836f
C231 B.n100 VSUBS 0.00836f
C232 B.n101 VSUBS 0.00836f
C233 B.n102 VSUBS 0.00836f
C234 B.n103 VSUBS 0.00836f
C235 B.n104 VSUBS 0.00836f
C236 B.n105 VSUBS 0.00836f
C237 B.n106 VSUBS 0.00836f
C238 B.n107 VSUBS 0.00836f
C239 B.n108 VSUBS 0.00836f
C240 B.n109 VSUBS 0.00836f
C241 B.n110 VSUBS 0.00836f
C242 B.n111 VSUBS 0.00836f
C243 B.n112 VSUBS 0.00836f
C244 B.n113 VSUBS 0.00836f
C245 B.n114 VSUBS 0.00836f
C246 B.n115 VSUBS 0.00836f
C247 B.n116 VSUBS 0.00836f
C248 B.n117 VSUBS 0.00836f
C249 B.n118 VSUBS 0.00836f
C250 B.n119 VSUBS 0.00836f
C251 B.n120 VSUBS 0.00836f
C252 B.n121 VSUBS 0.00836f
C253 B.n122 VSUBS 0.00836f
C254 B.n123 VSUBS 0.00836f
C255 B.n124 VSUBS 0.00836f
C256 B.n125 VSUBS 0.00836f
C257 B.n126 VSUBS 0.00836f
C258 B.n127 VSUBS 0.00836f
C259 B.n128 VSUBS 0.020999f
C260 B.n129 VSUBS 0.00836f
C261 B.n130 VSUBS 0.00836f
C262 B.n131 VSUBS 0.00836f
C263 B.n132 VSUBS 0.00836f
C264 B.n133 VSUBS 0.00836f
C265 B.n134 VSUBS 0.00836f
C266 B.n135 VSUBS 0.00836f
C267 B.n136 VSUBS 0.00836f
C268 B.n137 VSUBS 0.00836f
C269 B.n138 VSUBS 0.00836f
C270 B.n139 VSUBS 0.00836f
C271 B.n140 VSUBS 0.00836f
C272 B.n141 VSUBS 0.00836f
C273 B.n142 VSUBS 0.00836f
C274 B.n143 VSUBS 0.00836f
C275 B.t1 VSUBS 0.310275f
C276 B.t2 VSUBS 0.337801f
C277 B.t0 VSUBS 1.40453f
C278 B.n144 VSUBS 0.186948f
C279 B.n145 VSUBS 0.087327f
C280 B.n146 VSUBS 0.00836f
C281 B.n147 VSUBS 0.00836f
C282 B.n148 VSUBS 0.00836f
C283 B.n149 VSUBS 0.00836f
C284 B.t4 VSUBS 0.310278f
C285 B.t5 VSUBS 0.337804f
C286 B.t3 VSUBS 1.40453f
C287 B.n150 VSUBS 0.186944f
C288 B.n151 VSUBS 0.087325f
C289 B.n152 VSUBS 0.01937f
C290 B.n153 VSUBS 0.00836f
C291 B.n154 VSUBS 0.00836f
C292 B.n155 VSUBS 0.00836f
C293 B.n156 VSUBS 0.00836f
C294 B.n157 VSUBS 0.00836f
C295 B.n158 VSUBS 0.00836f
C296 B.n159 VSUBS 0.00836f
C297 B.n160 VSUBS 0.00836f
C298 B.n161 VSUBS 0.00836f
C299 B.n162 VSUBS 0.00836f
C300 B.n163 VSUBS 0.00836f
C301 B.n164 VSUBS 0.00836f
C302 B.n165 VSUBS 0.00836f
C303 B.n166 VSUBS 0.00836f
C304 B.n167 VSUBS 0.00836f
C305 B.n168 VSUBS 0.02031f
C306 B.n169 VSUBS 0.00836f
C307 B.n170 VSUBS 0.00836f
C308 B.n171 VSUBS 0.00836f
C309 B.n172 VSUBS 0.00836f
C310 B.n173 VSUBS 0.00836f
C311 B.n174 VSUBS 0.00836f
C312 B.n175 VSUBS 0.00836f
C313 B.n176 VSUBS 0.00836f
C314 B.n177 VSUBS 0.00836f
C315 B.n178 VSUBS 0.00836f
C316 B.n179 VSUBS 0.00836f
C317 B.n180 VSUBS 0.00836f
C318 B.n181 VSUBS 0.00836f
C319 B.n182 VSUBS 0.00836f
C320 B.n183 VSUBS 0.00836f
C321 B.n184 VSUBS 0.00836f
C322 B.n185 VSUBS 0.00836f
C323 B.n186 VSUBS 0.00836f
C324 B.n187 VSUBS 0.00836f
C325 B.n188 VSUBS 0.00836f
C326 B.n189 VSUBS 0.00836f
C327 B.n190 VSUBS 0.00836f
C328 B.n191 VSUBS 0.00836f
C329 B.n192 VSUBS 0.00836f
C330 B.n193 VSUBS 0.00836f
C331 B.n194 VSUBS 0.00836f
C332 B.n195 VSUBS 0.00836f
C333 B.n196 VSUBS 0.00836f
C334 B.n197 VSUBS 0.00836f
C335 B.n198 VSUBS 0.00836f
C336 B.n199 VSUBS 0.00836f
C337 B.n200 VSUBS 0.00836f
C338 B.n201 VSUBS 0.00836f
C339 B.n202 VSUBS 0.00836f
C340 B.n203 VSUBS 0.00836f
C341 B.n204 VSUBS 0.00836f
C342 B.n205 VSUBS 0.00836f
C343 B.n206 VSUBS 0.00836f
C344 B.n207 VSUBS 0.00836f
C345 B.n208 VSUBS 0.00836f
C346 B.n209 VSUBS 0.00836f
C347 B.n210 VSUBS 0.00836f
C348 B.n211 VSUBS 0.00836f
C349 B.n212 VSUBS 0.00836f
C350 B.n213 VSUBS 0.00836f
C351 B.n214 VSUBS 0.00836f
C352 B.n215 VSUBS 0.00836f
C353 B.n216 VSUBS 0.00836f
C354 B.n217 VSUBS 0.00836f
C355 B.n218 VSUBS 0.00836f
C356 B.n219 VSUBS 0.00836f
C357 B.n220 VSUBS 0.00836f
C358 B.n221 VSUBS 0.00836f
C359 B.n222 VSUBS 0.00836f
C360 B.n223 VSUBS 0.00836f
C361 B.n224 VSUBS 0.00836f
C362 B.n225 VSUBS 0.00836f
C363 B.n226 VSUBS 0.00836f
C364 B.n227 VSUBS 0.00836f
C365 B.n228 VSUBS 0.00836f
C366 B.n229 VSUBS 0.00836f
C367 B.n230 VSUBS 0.00836f
C368 B.n231 VSUBS 0.00836f
C369 B.n232 VSUBS 0.00836f
C370 B.n233 VSUBS 0.00836f
C371 B.n234 VSUBS 0.00836f
C372 B.n235 VSUBS 0.00836f
C373 B.n236 VSUBS 0.00836f
C374 B.n237 VSUBS 0.00836f
C375 B.n238 VSUBS 0.00836f
C376 B.n239 VSUBS 0.00836f
C377 B.n240 VSUBS 0.00836f
C378 B.n241 VSUBS 0.00836f
C379 B.n242 VSUBS 0.00836f
C380 B.n243 VSUBS 0.00836f
C381 B.n244 VSUBS 0.00836f
C382 B.n245 VSUBS 0.00836f
C383 B.n246 VSUBS 0.00836f
C384 B.n247 VSUBS 0.00836f
C385 B.n248 VSUBS 0.00836f
C386 B.n249 VSUBS 0.00836f
C387 B.n250 VSUBS 0.00836f
C388 B.n251 VSUBS 0.00836f
C389 B.n252 VSUBS 0.00836f
C390 B.n253 VSUBS 0.00836f
C391 B.n254 VSUBS 0.00836f
C392 B.n255 VSUBS 0.00836f
C393 B.n256 VSUBS 0.00836f
C394 B.n257 VSUBS 0.00836f
C395 B.n258 VSUBS 0.00836f
C396 B.n259 VSUBS 0.00836f
C397 B.n260 VSUBS 0.00836f
C398 B.n261 VSUBS 0.00836f
C399 B.n262 VSUBS 0.00836f
C400 B.n263 VSUBS 0.00836f
C401 B.n264 VSUBS 0.00836f
C402 B.n265 VSUBS 0.00836f
C403 B.n266 VSUBS 0.00836f
C404 B.n267 VSUBS 0.00836f
C405 B.n268 VSUBS 0.00836f
C406 B.n269 VSUBS 0.00836f
C407 B.n270 VSUBS 0.00836f
C408 B.n271 VSUBS 0.00836f
C409 B.n272 VSUBS 0.00836f
C410 B.n273 VSUBS 0.00836f
C411 B.n274 VSUBS 0.00836f
C412 B.n275 VSUBS 0.00836f
C413 B.n276 VSUBS 0.00836f
C414 B.n277 VSUBS 0.00836f
C415 B.n278 VSUBS 0.00836f
C416 B.n279 VSUBS 0.02031f
C417 B.n280 VSUBS 0.020999f
C418 B.n281 VSUBS 0.020999f
C419 B.n282 VSUBS 0.00836f
C420 B.n283 VSUBS 0.00836f
C421 B.n284 VSUBS 0.00836f
C422 B.n285 VSUBS 0.00836f
C423 B.n286 VSUBS 0.00836f
C424 B.n287 VSUBS 0.00836f
C425 B.n288 VSUBS 0.00836f
C426 B.n289 VSUBS 0.00836f
C427 B.n290 VSUBS 0.00836f
C428 B.n291 VSUBS 0.00836f
C429 B.n292 VSUBS 0.00836f
C430 B.n293 VSUBS 0.00836f
C431 B.n294 VSUBS 0.00836f
C432 B.n295 VSUBS 0.00836f
C433 B.n296 VSUBS 0.00836f
C434 B.n297 VSUBS 0.00836f
C435 B.n298 VSUBS 0.00836f
C436 B.n299 VSUBS 0.00836f
C437 B.n300 VSUBS 0.00836f
C438 B.n301 VSUBS 0.00836f
C439 B.n302 VSUBS 0.00836f
C440 B.n303 VSUBS 0.00836f
C441 B.n304 VSUBS 0.00836f
C442 B.n305 VSUBS 0.00836f
C443 B.n306 VSUBS 0.00836f
C444 B.n307 VSUBS 0.00836f
C445 B.n308 VSUBS 0.00836f
C446 B.n309 VSUBS 0.00836f
C447 B.n310 VSUBS 0.00836f
C448 B.n311 VSUBS 0.00836f
C449 B.n312 VSUBS 0.00836f
C450 B.n313 VSUBS 0.00836f
C451 B.n314 VSUBS 0.00836f
C452 B.n315 VSUBS 0.00836f
C453 B.n316 VSUBS 0.00836f
C454 B.n317 VSUBS 0.00836f
C455 B.n318 VSUBS 0.00836f
C456 B.n319 VSUBS 0.00836f
C457 B.n320 VSUBS 0.00836f
C458 B.n321 VSUBS 0.00836f
C459 B.n322 VSUBS 0.00836f
C460 B.n323 VSUBS 0.00836f
C461 B.n324 VSUBS 0.00836f
C462 B.n325 VSUBS 0.005778f
C463 B.n326 VSUBS 0.00836f
C464 B.n327 VSUBS 0.00836f
C465 B.n328 VSUBS 0.006762f
C466 B.n329 VSUBS 0.00836f
C467 B.n330 VSUBS 0.00836f
C468 B.n331 VSUBS 0.00836f
C469 B.n332 VSUBS 0.00836f
C470 B.n333 VSUBS 0.00836f
C471 B.n334 VSUBS 0.00836f
C472 B.n335 VSUBS 0.00836f
C473 B.n336 VSUBS 0.00836f
C474 B.n337 VSUBS 0.00836f
C475 B.n338 VSUBS 0.00836f
C476 B.n339 VSUBS 0.00836f
C477 B.n340 VSUBS 0.006762f
C478 B.n341 VSUBS 0.01937f
C479 B.n342 VSUBS 0.005778f
C480 B.n343 VSUBS 0.00836f
C481 B.n344 VSUBS 0.00836f
C482 B.n345 VSUBS 0.00836f
C483 B.n346 VSUBS 0.00836f
C484 B.n347 VSUBS 0.00836f
C485 B.n348 VSUBS 0.00836f
C486 B.n349 VSUBS 0.00836f
C487 B.n350 VSUBS 0.00836f
C488 B.n351 VSUBS 0.00836f
C489 B.n352 VSUBS 0.00836f
C490 B.n353 VSUBS 0.00836f
C491 B.n354 VSUBS 0.00836f
C492 B.n355 VSUBS 0.00836f
C493 B.n356 VSUBS 0.00836f
C494 B.n357 VSUBS 0.00836f
C495 B.n358 VSUBS 0.00836f
C496 B.n359 VSUBS 0.00836f
C497 B.n360 VSUBS 0.00836f
C498 B.n361 VSUBS 0.00836f
C499 B.n362 VSUBS 0.00836f
C500 B.n363 VSUBS 0.00836f
C501 B.n364 VSUBS 0.00836f
C502 B.n365 VSUBS 0.00836f
C503 B.n366 VSUBS 0.00836f
C504 B.n367 VSUBS 0.00836f
C505 B.n368 VSUBS 0.00836f
C506 B.n369 VSUBS 0.00836f
C507 B.n370 VSUBS 0.00836f
C508 B.n371 VSUBS 0.00836f
C509 B.n372 VSUBS 0.00836f
C510 B.n373 VSUBS 0.00836f
C511 B.n374 VSUBS 0.00836f
C512 B.n375 VSUBS 0.00836f
C513 B.n376 VSUBS 0.00836f
C514 B.n377 VSUBS 0.00836f
C515 B.n378 VSUBS 0.00836f
C516 B.n379 VSUBS 0.00836f
C517 B.n380 VSUBS 0.00836f
C518 B.n381 VSUBS 0.00836f
C519 B.n382 VSUBS 0.00836f
C520 B.n383 VSUBS 0.00836f
C521 B.n384 VSUBS 0.00836f
C522 B.n385 VSUBS 0.00836f
C523 B.n386 VSUBS 0.00836f
C524 B.n387 VSUBS 0.020999f
C525 B.n388 VSUBS 0.02031f
C526 B.n389 VSUBS 0.02031f
C527 B.n390 VSUBS 0.00836f
C528 B.n391 VSUBS 0.00836f
C529 B.n392 VSUBS 0.00836f
C530 B.n393 VSUBS 0.00836f
C531 B.n394 VSUBS 0.00836f
C532 B.n395 VSUBS 0.00836f
C533 B.n396 VSUBS 0.00836f
C534 B.n397 VSUBS 0.00836f
C535 B.n398 VSUBS 0.00836f
C536 B.n399 VSUBS 0.00836f
C537 B.n400 VSUBS 0.00836f
C538 B.n401 VSUBS 0.00836f
C539 B.n402 VSUBS 0.00836f
C540 B.n403 VSUBS 0.00836f
C541 B.n404 VSUBS 0.00836f
C542 B.n405 VSUBS 0.00836f
C543 B.n406 VSUBS 0.00836f
C544 B.n407 VSUBS 0.00836f
C545 B.n408 VSUBS 0.00836f
C546 B.n409 VSUBS 0.00836f
C547 B.n410 VSUBS 0.00836f
C548 B.n411 VSUBS 0.00836f
C549 B.n412 VSUBS 0.00836f
C550 B.n413 VSUBS 0.00836f
C551 B.n414 VSUBS 0.00836f
C552 B.n415 VSUBS 0.00836f
C553 B.n416 VSUBS 0.00836f
C554 B.n417 VSUBS 0.00836f
C555 B.n418 VSUBS 0.00836f
C556 B.n419 VSUBS 0.00836f
C557 B.n420 VSUBS 0.00836f
C558 B.n421 VSUBS 0.00836f
C559 B.n422 VSUBS 0.00836f
C560 B.n423 VSUBS 0.00836f
C561 B.n424 VSUBS 0.00836f
C562 B.n425 VSUBS 0.00836f
C563 B.n426 VSUBS 0.00836f
C564 B.n427 VSUBS 0.00836f
C565 B.n428 VSUBS 0.00836f
C566 B.n429 VSUBS 0.00836f
C567 B.n430 VSUBS 0.00836f
C568 B.n431 VSUBS 0.00836f
C569 B.n432 VSUBS 0.00836f
C570 B.n433 VSUBS 0.00836f
C571 B.n434 VSUBS 0.00836f
C572 B.n435 VSUBS 0.00836f
C573 B.n436 VSUBS 0.00836f
C574 B.n437 VSUBS 0.00836f
C575 B.n438 VSUBS 0.00836f
C576 B.n439 VSUBS 0.00836f
C577 B.n440 VSUBS 0.00836f
C578 B.n441 VSUBS 0.00836f
C579 B.n442 VSUBS 0.00836f
C580 B.n443 VSUBS 0.00836f
C581 B.n444 VSUBS 0.00836f
C582 B.n445 VSUBS 0.00836f
C583 B.n446 VSUBS 0.00836f
C584 B.n447 VSUBS 0.00836f
C585 B.n448 VSUBS 0.00836f
C586 B.n449 VSUBS 0.00836f
C587 B.n450 VSUBS 0.00836f
C588 B.n451 VSUBS 0.00836f
C589 B.n452 VSUBS 0.00836f
C590 B.n453 VSUBS 0.00836f
C591 B.n454 VSUBS 0.00836f
C592 B.n455 VSUBS 0.00836f
C593 B.n456 VSUBS 0.00836f
C594 B.n457 VSUBS 0.00836f
C595 B.n458 VSUBS 0.00836f
C596 B.n459 VSUBS 0.00836f
C597 B.n460 VSUBS 0.00836f
C598 B.n461 VSUBS 0.00836f
C599 B.n462 VSUBS 0.00836f
C600 B.n463 VSUBS 0.00836f
C601 B.n464 VSUBS 0.00836f
C602 B.n465 VSUBS 0.00836f
C603 B.n466 VSUBS 0.00836f
C604 B.n467 VSUBS 0.00836f
C605 B.n468 VSUBS 0.00836f
C606 B.n469 VSUBS 0.00836f
C607 B.n470 VSUBS 0.00836f
C608 B.n471 VSUBS 0.00836f
C609 B.n472 VSUBS 0.00836f
C610 B.n473 VSUBS 0.00836f
C611 B.n474 VSUBS 0.00836f
C612 B.n475 VSUBS 0.00836f
C613 B.n476 VSUBS 0.00836f
C614 B.n477 VSUBS 0.00836f
C615 B.n478 VSUBS 0.00836f
C616 B.n479 VSUBS 0.00836f
C617 B.n480 VSUBS 0.00836f
C618 B.n481 VSUBS 0.00836f
C619 B.n482 VSUBS 0.00836f
C620 B.n483 VSUBS 0.00836f
C621 B.n484 VSUBS 0.00836f
C622 B.n485 VSUBS 0.00836f
C623 B.n486 VSUBS 0.00836f
C624 B.n487 VSUBS 0.00836f
C625 B.n488 VSUBS 0.00836f
C626 B.n489 VSUBS 0.00836f
C627 B.n490 VSUBS 0.00836f
C628 B.n491 VSUBS 0.00836f
C629 B.n492 VSUBS 0.00836f
C630 B.n493 VSUBS 0.00836f
C631 B.n494 VSUBS 0.00836f
C632 B.n495 VSUBS 0.00836f
C633 B.n496 VSUBS 0.00836f
C634 B.n497 VSUBS 0.00836f
C635 B.n498 VSUBS 0.00836f
C636 B.n499 VSUBS 0.00836f
C637 B.n500 VSUBS 0.00836f
C638 B.n501 VSUBS 0.00836f
C639 B.n502 VSUBS 0.00836f
C640 B.n503 VSUBS 0.00836f
C641 B.n504 VSUBS 0.00836f
C642 B.n505 VSUBS 0.00836f
C643 B.n506 VSUBS 0.00836f
C644 B.n507 VSUBS 0.00836f
C645 B.n508 VSUBS 0.00836f
C646 B.n509 VSUBS 0.00836f
C647 B.n510 VSUBS 0.00836f
C648 B.n511 VSUBS 0.00836f
C649 B.n512 VSUBS 0.00836f
C650 B.n513 VSUBS 0.00836f
C651 B.n514 VSUBS 0.00836f
C652 B.n515 VSUBS 0.00836f
C653 B.n516 VSUBS 0.00836f
C654 B.n517 VSUBS 0.00836f
C655 B.n518 VSUBS 0.00836f
C656 B.n519 VSUBS 0.00836f
C657 B.n520 VSUBS 0.00836f
C658 B.n521 VSUBS 0.00836f
C659 B.n522 VSUBS 0.00836f
C660 B.n523 VSUBS 0.00836f
C661 B.n524 VSUBS 0.00836f
C662 B.n525 VSUBS 0.00836f
C663 B.n526 VSUBS 0.00836f
C664 B.n527 VSUBS 0.00836f
C665 B.n528 VSUBS 0.00836f
C666 B.n529 VSUBS 0.00836f
C667 B.n530 VSUBS 0.00836f
C668 B.n531 VSUBS 0.00836f
C669 B.n532 VSUBS 0.00836f
C670 B.n533 VSUBS 0.00836f
C671 B.n534 VSUBS 0.00836f
C672 B.n535 VSUBS 0.00836f
C673 B.n536 VSUBS 0.00836f
C674 B.n537 VSUBS 0.00836f
C675 B.n538 VSUBS 0.00836f
C676 B.n539 VSUBS 0.00836f
C677 B.n540 VSUBS 0.00836f
C678 B.n541 VSUBS 0.00836f
C679 B.n542 VSUBS 0.00836f
C680 B.n543 VSUBS 0.00836f
C681 B.n544 VSUBS 0.00836f
C682 B.n545 VSUBS 0.00836f
C683 B.n546 VSUBS 0.00836f
C684 B.n547 VSUBS 0.00836f
C685 B.n548 VSUBS 0.00836f
C686 B.n549 VSUBS 0.00836f
C687 B.n550 VSUBS 0.00836f
C688 B.n551 VSUBS 0.00836f
C689 B.n552 VSUBS 0.00836f
C690 B.n553 VSUBS 0.00836f
C691 B.n554 VSUBS 0.00836f
C692 B.n555 VSUBS 0.00836f
C693 B.n556 VSUBS 0.00836f
C694 B.n557 VSUBS 0.00836f
C695 B.n558 VSUBS 0.00836f
C696 B.n559 VSUBS 0.021221f
C697 B.n560 VSUBS 0.02031f
C698 B.n561 VSUBS 0.020999f
C699 B.n562 VSUBS 0.00836f
C700 B.n563 VSUBS 0.00836f
C701 B.n564 VSUBS 0.00836f
C702 B.n565 VSUBS 0.00836f
C703 B.n566 VSUBS 0.00836f
C704 B.n567 VSUBS 0.00836f
C705 B.n568 VSUBS 0.00836f
C706 B.n569 VSUBS 0.00836f
C707 B.n570 VSUBS 0.00836f
C708 B.n571 VSUBS 0.00836f
C709 B.n572 VSUBS 0.00836f
C710 B.n573 VSUBS 0.00836f
C711 B.n574 VSUBS 0.00836f
C712 B.n575 VSUBS 0.00836f
C713 B.n576 VSUBS 0.00836f
C714 B.n577 VSUBS 0.00836f
C715 B.n578 VSUBS 0.00836f
C716 B.n579 VSUBS 0.00836f
C717 B.n580 VSUBS 0.00836f
C718 B.n581 VSUBS 0.00836f
C719 B.n582 VSUBS 0.00836f
C720 B.n583 VSUBS 0.00836f
C721 B.n584 VSUBS 0.00836f
C722 B.n585 VSUBS 0.00836f
C723 B.n586 VSUBS 0.00836f
C724 B.n587 VSUBS 0.00836f
C725 B.n588 VSUBS 0.00836f
C726 B.n589 VSUBS 0.00836f
C727 B.n590 VSUBS 0.00836f
C728 B.n591 VSUBS 0.00836f
C729 B.n592 VSUBS 0.00836f
C730 B.n593 VSUBS 0.00836f
C731 B.n594 VSUBS 0.00836f
C732 B.n595 VSUBS 0.00836f
C733 B.n596 VSUBS 0.00836f
C734 B.n597 VSUBS 0.00836f
C735 B.n598 VSUBS 0.00836f
C736 B.n599 VSUBS 0.00836f
C737 B.n600 VSUBS 0.00836f
C738 B.n601 VSUBS 0.00836f
C739 B.n602 VSUBS 0.00836f
C740 B.n603 VSUBS 0.00836f
C741 B.n604 VSUBS 0.00836f
C742 B.n605 VSUBS 0.00836f
C743 B.n606 VSUBS 0.005778f
C744 B.n607 VSUBS 0.01937f
C745 B.n608 VSUBS 0.006762f
C746 B.n609 VSUBS 0.00836f
C747 B.n610 VSUBS 0.00836f
C748 B.n611 VSUBS 0.00836f
C749 B.n612 VSUBS 0.00836f
C750 B.n613 VSUBS 0.00836f
C751 B.n614 VSUBS 0.00836f
C752 B.n615 VSUBS 0.00836f
C753 B.n616 VSUBS 0.00836f
C754 B.n617 VSUBS 0.00836f
C755 B.n618 VSUBS 0.00836f
C756 B.n619 VSUBS 0.00836f
C757 B.n620 VSUBS 0.006762f
C758 B.n621 VSUBS 0.00836f
C759 B.n622 VSUBS 0.00836f
C760 B.n623 VSUBS 0.005778f
C761 B.n624 VSUBS 0.00836f
C762 B.n625 VSUBS 0.00836f
C763 B.n626 VSUBS 0.00836f
C764 B.n627 VSUBS 0.00836f
C765 B.n628 VSUBS 0.00836f
C766 B.n629 VSUBS 0.00836f
C767 B.n630 VSUBS 0.00836f
C768 B.n631 VSUBS 0.00836f
C769 B.n632 VSUBS 0.00836f
C770 B.n633 VSUBS 0.00836f
C771 B.n634 VSUBS 0.00836f
C772 B.n635 VSUBS 0.00836f
C773 B.n636 VSUBS 0.00836f
C774 B.n637 VSUBS 0.00836f
C775 B.n638 VSUBS 0.00836f
C776 B.n639 VSUBS 0.00836f
C777 B.n640 VSUBS 0.00836f
C778 B.n641 VSUBS 0.00836f
C779 B.n642 VSUBS 0.00836f
C780 B.n643 VSUBS 0.00836f
C781 B.n644 VSUBS 0.00836f
C782 B.n645 VSUBS 0.00836f
C783 B.n646 VSUBS 0.00836f
C784 B.n647 VSUBS 0.00836f
C785 B.n648 VSUBS 0.00836f
C786 B.n649 VSUBS 0.00836f
C787 B.n650 VSUBS 0.00836f
C788 B.n651 VSUBS 0.00836f
C789 B.n652 VSUBS 0.00836f
C790 B.n653 VSUBS 0.00836f
C791 B.n654 VSUBS 0.00836f
C792 B.n655 VSUBS 0.00836f
C793 B.n656 VSUBS 0.00836f
C794 B.n657 VSUBS 0.00836f
C795 B.n658 VSUBS 0.00836f
C796 B.n659 VSUBS 0.00836f
C797 B.n660 VSUBS 0.00836f
C798 B.n661 VSUBS 0.00836f
C799 B.n662 VSUBS 0.00836f
C800 B.n663 VSUBS 0.00836f
C801 B.n664 VSUBS 0.00836f
C802 B.n665 VSUBS 0.00836f
C803 B.n666 VSUBS 0.00836f
C804 B.n667 VSUBS 0.020999f
C805 B.n668 VSUBS 0.020999f
C806 B.n669 VSUBS 0.02031f
C807 B.n670 VSUBS 0.00836f
C808 B.n671 VSUBS 0.00836f
C809 B.n672 VSUBS 0.00836f
C810 B.n673 VSUBS 0.00836f
C811 B.n674 VSUBS 0.00836f
C812 B.n675 VSUBS 0.00836f
C813 B.n676 VSUBS 0.00836f
C814 B.n677 VSUBS 0.00836f
C815 B.n678 VSUBS 0.00836f
C816 B.n679 VSUBS 0.00836f
C817 B.n680 VSUBS 0.00836f
C818 B.n681 VSUBS 0.00836f
C819 B.n682 VSUBS 0.00836f
C820 B.n683 VSUBS 0.00836f
C821 B.n684 VSUBS 0.00836f
C822 B.n685 VSUBS 0.00836f
C823 B.n686 VSUBS 0.00836f
C824 B.n687 VSUBS 0.00836f
C825 B.n688 VSUBS 0.00836f
C826 B.n689 VSUBS 0.00836f
C827 B.n690 VSUBS 0.00836f
C828 B.n691 VSUBS 0.00836f
C829 B.n692 VSUBS 0.00836f
C830 B.n693 VSUBS 0.00836f
C831 B.n694 VSUBS 0.00836f
C832 B.n695 VSUBS 0.00836f
C833 B.n696 VSUBS 0.00836f
C834 B.n697 VSUBS 0.00836f
C835 B.n698 VSUBS 0.00836f
C836 B.n699 VSUBS 0.00836f
C837 B.n700 VSUBS 0.00836f
C838 B.n701 VSUBS 0.00836f
C839 B.n702 VSUBS 0.00836f
C840 B.n703 VSUBS 0.00836f
C841 B.n704 VSUBS 0.00836f
C842 B.n705 VSUBS 0.00836f
C843 B.n706 VSUBS 0.00836f
C844 B.n707 VSUBS 0.00836f
C845 B.n708 VSUBS 0.00836f
C846 B.n709 VSUBS 0.00836f
C847 B.n710 VSUBS 0.00836f
C848 B.n711 VSUBS 0.00836f
C849 B.n712 VSUBS 0.00836f
C850 B.n713 VSUBS 0.00836f
C851 B.n714 VSUBS 0.00836f
C852 B.n715 VSUBS 0.00836f
C853 B.n716 VSUBS 0.00836f
C854 B.n717 VSUBS 0.00836f
C855 B.n718 VSUBS 0.00836f
C856 B.n719 VSUBS 0.00836f
C857 B.n720 VSUBS 0.00836f
C858 B.n721 VSUBS 0.00836f
C859 B.n722 VSUBS 0.00836f
C860 B.n723 VSUBS 0.00836f
C861 B.n724 VSUBS 0.00836f
C862 B.n725 VSUBS 0.00836f
C863 B.n726 VSUBS 0.00836f
C864 B.n727 VSUBS 0.00836f
C865 B.n728 VSUBS 0.00836f
C866 B.n729 VSUBS 0.00836f
C867 B.n730 VSUBS 0.00836f
C868 B.n731 VSUBS 0.00836f
C869 B.n732 VSUBS 0.00836f
C870 B.n733 VSUBS 0.00836f
C871 B.n734 VSUBS 0.00836f
C872 B.n735 VSUBS 0.00836f
C873 B.n736 VSUBS 0.00836f
C874 B.n737 VSUBS 0.00836f
C875 B.n738 VSUBS 0.00836f
C876 B.n739 VSUBS 0.00836f
C877 B.n740 VSUBS 0.00836f
C878 B.n741 VSUBS 0.00836f
C879 B.n742 VSUBS 0.00836f
C880 B.n743 VSUBS 0.00836f
C881 B.n744 VSUBS 0.00836f
C882 B.n745 VSUBS 0.00836f
C883 B.n746 VSUBS 0.00836f
C884 B.n747 VSUBS 0.00836f
C885 B.n748 VSUBS 0.00836f
C886 B.n749 VSUBS 0.00836f
C887 B.n750 VSUBS 0.00836f
C888 B.n751 VSUBS 0.00836f
C889 B.n752 VSUBS 0.00836f
C890 B.n753 VSUBS 0.00836f
C891 B.n754 VSUBS 0.00836f
C892 B.n755 VSUBS 0.01893f
C893 VDD2.t6 VSUBS 0.184761f
C894 VDD2.t1 VSUBS 0.184761f
C895 VDD2.n0 VSUBS 1.36882f
C896 VDD2.t2 VSUBS 0.184761f
C897 VDD2.t7 VSUBS 0.184761f
C898 VDD2.n1 VSUBS 1.36882f
C899 VDD2.n2 VSUBS 4.15976f
C900 VDD2.t0 VSUBS 0.184761f
C901 VDD2.t5 VSUBS 0.184761f
C902 VDD2.n3 VSUBS 1.35497f
C903 VDD2.n4 VSUBS 3.38758f
C904 VDD2.t3 VSUBS 0.184761f
C905 VDD2.t4 VSUBS 0.184761f
C906 VDD2.n5 VSUBS 1.36878f
C907 VTAIL.t10 VSUBS 0.180889f
C908 VTAIL.t9 VSUBS 0.180889f
C909 VTAIL.n0 VSUBS 1.21476f
C910 VTAIL.n1 VSUBS 0.797293f
C911 VTAIL.t15 VSUBS 1.62604f
C912 VTAIL.n2 VSUBS 0.915663f
C913 VTAIL.t6 VSUBS 1.62604f
C914 VTAIL.n3 VSUBS 0.915663f
C915 VTAIL.t2 VSUBS 0.180889f
C916 VTAIL.t0 VSUBS 0.180889f
C917 VTAIL.n4 VSUBS 1.21476f
C918 VTAIL.n5 VSUBS 1.04544f
C919 VTAIL.t1 VSUBS 1.62604f
C920 VTAIL.n6 VSUBS 2.13528f
C921 VTAIL.t8 VSUBS 1.62605f
C922 VTAIL.n7 VSUBS 2.13527f
C923 VTAIL.t13 VSUBS 0.180889f
C924 VTAIL.t12 VSUBS 0.180889f
C925 VTAIL.n8 VSUBS 1.21476f
C926 VTAIL.n9 VSUBS 1.04543f
C927 VTAIL.t11 VSUBS 1.62605f
C928 VTAIL.n10 VSUBS 0.915652f
C929 VTAIL.t5 VSUBS 1.62605f
C930 VTAIL.n11 VSUBS 0.915652f
C931 VTAIL.t4 VSUBS 0.180889f
C932 VTAIL.t3 VSUBS 0.180889f
C933 VTAIL.n12 VSUBS 1.21476f
C934 VTAIL.n13 VSUBS 1.04543f
C935 VTAIL.t7 VSUBS 1.62604f
C936 VTAIL.n14 VSUBS 2.13528f
C937 VTAIL.t14 VSUBS 1.62604f
C938 VTAIL.n15 VSUBS 2.13015f
C939 VN.t0 VSUBS 2.0573f
C940 VN.n0 VSUBS 0.871222f
C941 VN.n1 VSUBS 0.030486f
C942 VN.n2 VSUBS 0.051064f
C943 VN.n3 VSUBS 0.030486f
C944 VN.t5 VSUBS 2.0573f
C945 VN.n4 VSUBS 0.056534f
C946 VN.n5 VSUBS 0.030486f
C947 VN.n6 VSUBS 0.056534f
C948 VN.t1 VSUBS 2.36315f
C949 VN.n7 VSUBS 0.806092f
C950 VN.t6 VSUBS 2.0573f
C951 VN.n8 VSUBS 0.834132f
C952 VN.n9 VSUBS 0.037834f
C953 VN.n10 VSUBS 0.326906f
C954 VN.n11 VSUBS 0.030486f
C955 VN.n12 VSUBS 0.030486f
C956 VN.n13 VSUBS 0.060272f
C957 VN.n14 VSUBS 0.024622f
C958 VN.n15 VSUBS 0.060272f
C959 VN.n16 VSUBS 0.030486f
C960 VN.n17 VSUBS 0.030486f
C961 VN.n18 VSUBS 0.030486f
C962 VN.n19 VSUBS 0.037834f
C963 VN.n20 VSUBS 0.742156f
C964 VN.n21 VSUBS 0.047324f
C965 VN.n22 VSUBS 0.056534f
C966 VN.n23 VSUBS 0.030486f
C967 VN.n24 VSUBS 0.030486f
C968 VN.n25 VSUBS 0.030486f
C969 VN.n26 VSUBS 0.037569f
C970 VN.n27 VSUBS 0.056534f
C971 VN.n28 VSUBS 0.056255f
C972 VN.n29 VSUBS 0.049196f
C973 VN.n30 VSUBS 0.057008f
C974 VN.t7 VSUBS 2.0573f
C975 VN.n31 VSUBS 0.871222f
C976 VN.n32 VSUBS 0.030486f
C977 VN.n33 VSUBS 0.051064f
C978 VN.n34 VSUBS 0.030486f
C979 VN.t2 VSUBS 2.0573f
C980 VN.n35 VSUBS 0.056534f
C981 VN.n36 VSUBS 0.030486f
C982 VN.n37 VSUBS 0.056534f
C983 VN.t3 VSUBS 2.36315f
C984 VN.n38 VSUBS 0.806092f
C985 VN.t4 VSUBS 2.0573f
C986 VN.n39 VSUBS 0.834132f
C987 VN.n40 VSUBS 0.037834f
C988 VN.n41 VSUBS 0.326906f
C989 VN.n42 VSUBS 0.030486f
C990 VN.n43 VSUBS 0.030486f
C991 VN.n44 VSUBS 0.060272f
C992 VN.n45 VSUBS 0.024622f
C993 VN.n46 VSUBS 0.060272f
C994 VN.n47 VSUBS 0.030486f
C995 VN.n48 VSUBS 0.030486f
C996 VN.n49 VSUBS 0.030486f
C997 VN.n50 VSUBS 0.037834f
C998 VN.n51 VSUBS 0.742156f
C999 VN.n52 VSUBS 0.047324f
C1000 VN.n53 VSUBS 0.056534f
C1001 VN.n54 VSUBS 0.030486f
C1002 VN.n55 VSUBS 0.030486f
C1003 VN.n56 VSUBS 0.030486f
C1004 VN.n57 VSUBS 0.037569f
C1005 VN.n58 VSUBS 0.056534f
C1006 VN.n59 VSUBS 0.056255f
C1007 VN.n60 VSUBS 0.049196f
C1008 VN.n61 VSUBS 1.74077f
.ends

