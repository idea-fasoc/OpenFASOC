* NGSPICE file created from diff_pair_sample_1628.ext - technology: sky130A

.subckt diff_pair_sample_1628 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X1 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=0 ps=0 w=8.56 l=1.03
X2 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=1.4124 ps=8.89 w=8.56 l=1.03
X3 VTAIL.t14 VP.t1 VDD1.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X4 VDD1.t2 VP.t2 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=3.3384 ps=17.9 w=8.56 l=1.03
X5 VDD1.t0 VP.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X6 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=0 ps=0 w=8.56 l=1.03
X7 VDD1.t4 VP.t4 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=3.3384 ps=17.9 w=8.56 l=1.03
X8 VDD2.t6 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X9 VTAIL.t10 VP.t5 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=1.4124 ps=8.89 w=8.56 l=1.03
X10 VDD2.t5 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=3.3384 ps=17.9 w=8.56 l=1.03
X11 VTAIL.t5 VN.t3 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=1.4124 ps=8.89 w=8.56 l=1.03
X12 VDD1.t1 VP.t6 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X13 VTAIL.t7 VN.t4 VDD2.t3 B.t21 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X14 VDD2.t2 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=3.3384 ps=17.9 w=8.56 l=1.03
X15 VDD2.t1 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X16 VTAIL.t0 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4124 pd=8.89 as=1.4124 ps=8.89 w=8.56 l=1.03
X17 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=0 ps=0 w=8.56 l=1.03
X18 VTAIL.t8 VP.t7 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=1.4124 ps=8.89 w=8.56 l=1.03
X19 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=3.3384 pd=17.9 as=0 ps=0 w=8.56 l=1.03
R0 VP.n9 VP.t7 255.736
R1 VP.n21 VP.t5 238.894
R2 VP.n33 VP.t2 238.894
R3 VP.n18 VP.t4 238.894
R4 VP.n3 VP.t6 200.287
R5 VP.n1 VP.t0 200.287
R6 VP.n6 VP.t1 200.287
R7 VP.n8 VP.t3 200.287
R8 VP.n34 VP.n33 161.3
R9 VP.n11 VP.n10 161.3
R10 VP.n12 VP.n7 161.3
R11 VP.n14 VP.n13 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n5 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n32 VP.n0 161.3
R16 VP.n31 VP.n30 161.3
R17 VP.n29 VP.n28 161.3
R18 VP.n27 VP.n2 161.3
R19 VP.n26 VP.n25 161.3
R20 VP.n24 VP.n23 161.3
R21 VP.n22 VP.n4 161.3
R22 VP.n21 VP.n20 161.3
R23 VP.n23 VP.n22 54.0429
R24 VP.n32 VP.n31 54.0429
R25 VP.n17 VP.n16 54.0429
R26 VP.n9 VP.n8 45.8978
R27 VP.n10 VP.n9 43.6106
R28 VP.n20 VP.n19 41.0081
R29 VP.n27 VP.n26 40.4106
R30 VP.n28 VP.n27 40.4106
R31 VP.n13 VP.n12 40.4106
R32 VP.n12 VP.n11 40.4106
R33 VP.n23 VP.n3 15.5803
R34 VP.n31 VP.n1 15.5803
R35 VP.n16 VP.n6 15.5803
R36 VP.n26 VP.n3 8.76414
R37 VP.n28 VP.n1 8.76414
R38 VP.n13 VP.n6 8.76414
R39 VP.n11 VP.n8 8.76414
R40 VP.n22 VP.n21 3.65202
R41 VP.n33 VP.n32 3.65202
R42 VP.n18 VP.n17 3.65202
R43 VP.n10 VP.n7 0.189894
R44 VP.n14 VP.n7 0.189894
R45 VP.n15 VP.n14 0.189894
R46 VP.n15 VP.n5 0.189894
R47 VP.n19 VP.n5 0.189894
R48 VP.n20 VP.n4 0.189894
R49 VP.n24 VP.n4 0.189894
R50 VP.n25 VP.n24 0.189894
R51 VP.n25 VP.n2 0.189894
R52 VP.n29 VP.n2 0.189894
R53 VP.n30 VP.n29 0.189894
R54 VP.n30 VP.n0 0.189894
R55 VP.n34 VP.n0 0.189894
R56 VP VP.n34 0.0516364
R57 VDD1 VDD1.n0 64.8613
R58 VDD1.n3 VDD1.n2 64.7476
R59 VDD1.n3 VDD1.n1 64.7476
R60 VDD1.n5 VDD1.n4 64.2168
R61 VDD1.n5 VDD1.n3 36.9535
R62 VDD1.n4 VDD1.t7 2.31358
R63 VDD1.n4 VDD1.t4 2.31358
R64 VDD1.n0 VDD1.t6 2.31358
R65 VDD1.n0 VDD1.t0 2.31358
R66 VDD1.n2 VDD1.t5 2.31358
R67 VDD1.n2 VDD1.t2 2.31358
R68 VDD1.n1 VDD1.t3 2.31358
R69 VDD1.n1 VDD1.t1 2.31358
R70 VDD1 VDD1.n5 0.528517
R71 VTAIL.n370 VTAIL.n330 289.615
R72 VTAIL.n42 VTAIL.n2 289.615
R73 VTAIL.n88 VTAIL.n48 289.615
R74 VTAIL.n136 VTAIL.n96 289.615
R75 VTAIL.n324 VTAIL.n284 289.615
R76 VTAIL.n276 VTAIL.n236 289.615
R77 VTAIL.n230 VTAIL.n190 289.615
R78 VTAIL.n182 VTAIL.n142 289.615
R79 VTAIL.n345 VTAIL.n344 185
R80 VTAIL.n342 VTAIL.n341 185
R81 VTAIL.n351 VTAIL.n350 185
R82 VTAIL.n353 VTAIL.n352 185
R83 VTAIL.n338 VTAIL.n337 185
R84 VTAIL.n359 VTAIL.n358 185
R85 VTAIL.n362 VTAIL.n361 185
R86 VTAIL.n360 VTAIL.n334 185
R87 VTAIL.n367 VTAIL.n333 185
R88 VTAIL.n369 VTAIL.n368 185
R89 VTAIL.n371 VTAIL.n370 185
R90 VTAIL.n17 VTAIL.n16 185
R91 VTAIL.n14 VTAIL.n13 185
R92 VTAIL.n23 VTAIL.n22 185
R93 VTAIL.n25 VTAIL.n24 185
R94 VTAIL.n10 VTAIL.n9 185
R95 VTAIL.n31 VTAIL.n30 185
R96 VTAIL.n34 VTAIL.n33 185
R97 VTAIL.n32 VTAIL.n6 185
R98 VTAIL.n39 VTAIL.n5 185
R99 VTAIL.n41 VTAIL.n40 185
R100 VTAIL.n43 VTAIL.n42 185
R101 VTAIL.n63 VTAIL.n62 185
R102 VTAIL.n60 VTAIL.n59 185
R103 VTAIL.n69 VTAIL.n68 185
R104 VTAIL.n71 VTAIL.n70 185
R105 VTAIL.n56 VTAIL.n55 185
R106 VTAIL.n77 VTAIL.n76 185
R107 VTAIL.n80 VTAIL.n79 185
R108 VTAIL.n78 VTAIL.n52 185
R109 VTAIL.n85 VTAIL.n51 185
R110 VTAIL.n87 VTAIL.n86 185
R111 VTAIL.n89 VTAIL.n88 185
R112 VTAIL.n111 VTAIL.n110 185
R113 VTAIL.n108 VTAIL.n107 185
R114 VTAIL.n117 VTAIL.n116 185
R115 VTAIL.n119 VTAIL.n118 185
R116 VTAIL.n104 VTAIL.n103 185
R117 VTAIL.n125 VTAIL.n124 185
R118 VTAIL.n128 VTAIL.n127 185
R119 VTAIL.n126 VTAIL.n100 185
R120 VTAIL.n133 VTAIL.n99 185
R121 VTAIL.n135 VTAIL.n134 185
R122 VTAIL.n137 VTAIL.n136 185
R123 VTAIL.n325 VTAIL.n324 185
R124 VTAIL.n323 VTAIL.n322 185
R125 VTAIL.n321 VTAIL.n287 185
R126 VTAIL.n291 VTAIL.n288 185
R127 VTAIL.n316 VTAIL.n315 185
R128 VTAIL.n314 VTAIL.n313 185
R129 VTAIL.n293 VTAIL.n292 185
R130 VTAIL.n308 VTAIL.n307 185
R131 VTAIL.n306 VTAIL.n305 185
R132 VTAIL.n297 VTAIL.n296 185
R133 VTAIL.n300 VTAIL.n299 185
R134 VTAIL.n277 VTAIL.n276 185
R135 VTAIL.n275 VTAIL.n274 185
R136 VTAIL.n273 VTAIL.n239 185
R137 VTAIL.n243 VTAIL.n240 185
R138 VTAIL.n268 VTAIL.n267 185
R139 VTAIL.n266 VTAIL.n265 185
R140 VTAIL.n245 VTAIL.n244 185
R141 VTAIL.n260 VTAIL.n259 185
R142 VTAIL.n258 VTAIL.n257 185
R143 VTAIL.n249 VTAIL.n248 185
R144 VTAIL.n252 VTAIL.n251 185
R145 VTAIL.n231 VTAIL.n230 185
R146 VTAIL.n229 VTAIL.n228 185
R147 VTAIL.n227 VTAIL.n193 185
R148 VTAIL.n197 VTAIL.n194 185
R149 VTAIL.n222 VTAIL.n221 185
R150 VTAIL.n220 VTAIL.n219 185
R151 VTAIL.n199 VTAIL.n198 185
R152 VTAIL.n214 VTAIL.n213 185
R153 VTAIL.n212 VTAIL.n211 185
R154 VTAIL.n203 VTAIL.n202 185
R155 VTAIL.n206 VTAIL.n205 185
R156 VTAIL.n183 VTAIL.n182 185
R157 VTAIL.n181 VTAIL.n180 185
R158 VTAIL.n179 VTAIL.n145 185
R159 VTAIL.n149 VTAIL.n146 185
R160 VTAIL.n174 VTAIL.n173 185
R161 VTAIL.n172 VTAIL.n171 185
R162 VTAIL.n151 VTAIL.n150 185
R163 VTAIL.n166 VTAIL.n165 185
R164 VTAIL.n164 VTAIL.n163 185
R165 VTAIL.n155 VTAIL.n154 185
R166 VTAIL.n158 VTAIL.n157 185
R167 VTAIL.t3 VTAIL.n343 149.524
R168 VTAIL.t5 VTAIL.n15 149.524
R169 VTAIL.t13 VTAIL.n61 149.524
R170 VTAIL.t10 VTAIL.n109 149.524
R171 VTAIL.t11 VTAIL.n298 149.524
R172 VTAIL.t8 VTAIL.n250 149.524
R173 VTAIL.t6 VTAIL.n204 149.524
R174 VTAIL.t2 VTAIL.n156 149.524
R175 VTAIL.n344 VTAIL.n341 104.615
R176 VTAIL.n351 VTAIL.n341 104.615
R177 VTAIL.n352 VTAIL.n351 104.615
R178 VTAIL.n352 VTAIL.n337 104.615
R179 VTAIL.n359 VTAIL.n337 104.615
R180 VTAIL.n361 VTAIL.n359 104.615
R181 VTAIL.n361 VTAIL.n360 104.615
R182 VTAIL.n360 VTAIL.n333 104.615
R183 VTAIL.n369 VTAIL.n333 104.615
R184 VTAIL.n370 VTAIL.n369 104.615
R185 VTAIL.n16 VTAIL.n13 104.615
R186 VTAIL.n23 VTAIL.n13 104.615
R187 VTAIL.n24 VTAIL.n23 104.615
R188 VTAIL.n24 VTAIL.n9 104.615
R189 VTAIL.n31 VTAIL.n9 104.615
R190 VTAIL.n33 VTAIL.n31 104.615
R191 VTAIL.n33 VTAIL.n32 104.615
R192 VTAIL.n32 VTAIL.n5 104.615
R193 VTAIL.n41 VTAIL.n5 104.615
R194 VTAIL.n42 VTAIL.n41 104.615
R195 VTAIL.n62 VTAIL.n59 104.615
R196 VTAIL.n69 VTAIL.n59 104.615
R197 VTAIL.n70 VTAIL.n69 104.615
R198 VTAIL.n70 VTAIL.n55 104.615
R199 VTAIL.n77 VTAIL.n55 104.615
R200 VTAIL.n79 VTAIL.n77 104.615
R201 VTAIL.n79 VTAIL.n78 104.615
R202 VTAIL.n78 VTAIL.n51 104.615
R203 VTAIL.n87 VTAIL.n51 104.615
R204 VTAIL.n88 VTAIL.n87 104.615
R205 VTAIL.n110 VTAIL.n107 104.615
R206 VTAIL.n117 VTAIL.n107 104.615
R207 VTAIL.n118 VTAIL.n117 104.615
R208 VTAIL.n118 VTAIL.n103 104.615
R209 VTAIL.n125 VTAIL.n103 104.615
R210 VTAIL.n127 VTAIL.n125 104.615
R211 VTAIL.n127 VTAIL.n126 104.615
R212 VTAIL.n126 VTAIL.n99 104.615
R213 VTAIL.n135 VTAIL.n99 104.615
R214 VTAIL.n136 VTAIL.n135 104.615
R215 VTAIL.n324 VTAIL.n323 104.615
R216 VTAIL.n323 VTAIL.n287 104.615
R217 VTAIL.n291 VTAIL.n287 104.615
R218 VTAIL.n315 VTAIL.n291 104.615
R219 VTAIL.n315 VTAIL.n314 104.615
R220 VTAIL.n314 VTAIL.n292 104.615
R221 VTAIL.n307 VTAIL.n292 104.615
R222 VTAIL.n307 VTAIL.n306 104.615
R223 VTAIL.n306 VTAIL.n296 104.615
R224 VTAIL.n299 VTAIL.n296 104.615
R225 VTAIL.n276 VTAIL.n275 104.615
R226 VTAIL.n275 VTAIL.n239 104.615
R227 VTAIL.n243 VTAIL.n239 104.615
R228 VTAIL.n267 VTAIL.n243 104.615
R229 VTAIL.n267 VTAIL.n266 104.615
R230 VTAIL.n266 VTAIL.n244 104.615
R231 VTAIL.n259 VTAIL.n244 104.615
R232 VTAIL.n259 VTAIL.n258 104.615
R233 VTAIL.n258 VTAIL.n248 104.615
R234 VTAIL.n251 VTAIL.n248 104.615
R235 VTAIL.n230 VTAIL.n229 104.615
R236 VTAIL.n229 VTAIL.n193 104.615
R237 VTAIL.n197 VTAIL.n193 104.615
R238 VTAIL.n221 VTAIL.n197 104.615
R239 VTAIL.n221 VTAIL.n220 104.615
R240 VTAIL.n220 VTAIL.n198 104.615
R241 VTAIL.n213 VTAIL.n198 104.615
R242 VTAIL.n213 VTAIL.n212 104.615
R243 VTAIL.n212 VTAIL.n202 104.615
R244 VTAIL.n205 VTAIL.n202 104.615
R245 VTAIL.n182 VTAIL.n181 104.615
R246 VTAIL.n181 VTAIL.n145 104.615
R247 VTAIL.n149 VTAIL.n145 104.615
R248 VTAIL.n173 VTAIL.n149 104.615
R249 VTAIL.n173 VTAIL.n172 104.615
R250 VTAIL.n172 VTAIL.n150 104.615
R251 VTAIL.n165 VTAIL.n150 104.615
R252 VTAIL.n165 VTAIL.n164 104.615
R253 VTAIL.n164 VTAIL.n154 104.615
R254 VTAIL.n157 VTAIL.n154 104.615
R255 VTAIL.n344 VTAIL.t3 52.3082
R256 VTAIL.n16 VTAIL.t5 52.3082
R257 VTAIL.n62 VTAIL.t13 52.3082
R258 VTAIL.n110 VTAIL.t10 52.3082
R259 VTAIL.n299 VTAIL.t11 52.3082
R260 VTAIL.n251 VTAIL.t8 52.3082
R261 VTAIL.n205 VTAIL.t6 52.3082
R262 VTAIL.n157 VTAIL.t2 52.3082
R263 VTAIL.n283 VTAIL.n282 47.5381
R264 VTAIL.n189 VTAIL.n188 47.5381
R265 VTAIL.n1 VTAIL.n0 47.538
R266 VTAIL.n95 VTAIL.n94 47.538
R267 VTAIL.n375 VTAIL.n374 32.9611
R268 VTAIL.n47 VTAIL.n46 32.9611
R269 VTAIL.n93 VTAIL.n92 32.9611
R270 VTAIL.n141 VTAIL.n140 32.9611
R271 VTAIL.n329 VTAIL.n328 32.9611
R272 VTAIL.n281 VTAIL.n280 32.9611
R273 VTAIL.n235 VTAIL.n234 32.9611
R274 VTAIL.n187 VTAIL.n186 32.9611
R275 VTAIL.n375 VTAIL.n329 20.9186
R276 VTAIL.n187 VTAIL.n141 20.9186
R277 VTAIL.n368 VTAIL.n367 13.1884
R278 VTAIL.n40 VTAIL.n39 13.1884
R279 VTAIL.n86 VTAIL.n85 13.1884
R280 VTAIL.n134 VTAIL.n133 13.1884
R281 VTAIL.n322 VTAIL.n321 13.1884
R282 VTAIL.n274 VTAIL.n273 13.1884
R283 VTAIL.n228 VTAIL.n227 13.1884
R284 VTAIL.n180 VTAIL.n179 13.1884
R285 VTAIL.n366 VTAIL.n334 12.8005
R286 VTAIL.n371 VTAIL.n332 12.8005
R287 VTAIL.n38 VTAIL.n6 12.8005
R288 VTAIL.n43 VTAIL.n4 12.8005
R289 VTAIL.n84 VTAIL.n52 12.8005
R290 VTAIL.n89 VTAIL.n50 12.8005
R291 VTAIL.n132 VTAIL.n100 12.8005
R292 VTAIL.n137 VTAIL.n98 12.8005
R293 VTAIL.n325 VTAIL.n286 12.8005
R294 VTAIL.n320 VTAIL.n288 12.8005
R295 VTAIL.n277 VTAIL.n238 12.8005
R296 VTAIL.n272 VTAIL.n240 12.8005
R297 VTAIL.n231 VTAIL.n192 12.8005
R298 VTAIL.n226 VTAIL.n194 12.8005
R299 VTAIL.n183 VTAIL.n144 12.8005
R300 VTAIL.n178 VTAIL.n146 12.8005
R301 VTAIL.n363 VTAIL.n362 12.0247
R302 VTAIL.n372 VTAIL.n330 12.0247
R303 VTAIL.n35 VTAIL.n34 12.0247
R304 VTAIL.n44 VTAIL.n2 12.0247
R305 VTAIL.n81 VTAIL.n80 12.0247
R306 VTAIL.n90 VTAIL.n48 12.0247
R307 VTAIL.n129 VTAIL.n128 12.0247
R308 VTAIL.n138 VTAIL.n96 12.0247
R309 VTAIL.n326 VTAIL.n284 12.0247
R310 VTAIL.n317 VTAIL.n316 12.0247
R311 VTAIL.n278 VTAIL.n236 12.0247
R312 VTAIL.n269 VTAIL.n268 12.0247
R313 VTAIL.n232 VTAIL.n190 12.0247
R314 VTAIL.n223 VTAIL.n222 12.0247
R315 VTAIL.n184 VTAIL.n142 12.0247
R316 VTAIL.n175 VTAIL.n174 12.0247
R317 VTAIL.n358 VTAIL.n336 11.249
R318 VTAIL.n30 VTAIL.n8 11.249
R319 VTAIL.n76 VTAIL.n54 11.249
R320 VTAIL.n124 VTAIL.n102 11.249
R321 VTAIL.n313 VTAIL.n290 11.249
R322 VTAIL.n265 VTAIL.n242 11.249
R323 VTAIL.n219 VTAIL.n196 11.249
R324 VTAIL.n171 VTAIL.n148 11.249
R325 VTAIL.n357 VTAIL.n338 10.4732
R326 VTAIL.n29 VTAIL.n10 10.4732
R327 VTAIL.n75 VTAIL.n56 10.4732
R328 VTAIL.n123 VTAIL.n104 10.4732
R329 VTAIL.n312 VTAIL.n293 10.4732
R330 VTAIL.n264 VTAIL.n245 10.4732
R331 VTAIL.n218 VTAIL.n199 10.4732
R332 VTAIL.n170 VTAIL.n151 10.4732
R333 VTAIL.n345 VTAIL.n343 10.2747
R334 VTAIL.n17 VTAIL.n15 10.2747
R335 VTAIL.n63 VTAIL.n61 10.2747
R336 VTAIL.n111 VTAIL.n109 10.2747
R337 VTAIL.n300 VTAIL.n298 10.2747
R338 VTAIL.n252 VTAIL.n250 10.2747
R339 VTAIL.n206 VTAIL.n204 10.2747
R340 VTAIL.n158 VTAIL.n156 10.2747
R341 VTAIL.n354 VTAIL.n353 9.69747
R342 VTAIL.n26 VTAIL.n25 9.69747
R343 VTAIL.n72 VTAIL.n71 9.69747
R344 VTAIL.n120 VTAIL.n119 9.69747
R345 VTAIL.n309 VTAIL.n308 9.69747
R346 VTAIL.n261 VTAIL.n260 9.69747
R347 VTAIL.n215 VTAIL.n214 9.69747
R348 VTAIL.n167 VTAIL.n166 9.69747
R349 VTAIL.n374 VTAIL.n373 9.45567
R350 VTAIL.n46 VTAIL.n45 9.45567
R351 VTAIL.n92 VTAIL.n91 9.45567
R352 VTAIL.n140 VTAIL.n139 9.45567
R353 VTAIL.n328 VTAIL.n327 9.45567
R354 VTAIL.n280 VTAIL.n279 9.45567
R355 VTAIL.n234 VTAIL.n233 9.45567
R356 VTAIL.n186 VTAIL.n185 9.45567
R357 VTAIL.n373 VTAIL.n372 9.3005
R358 VTAIL.n332 VTAIL.n331 9.3005
R359 VTAIL.n347 VTAIL.n346 9.3005
R360 VTAIL.n349 VTAIL.n348 9.3005
R361 VTAIL.n340 VTAIL.n339 9.3005
R362 VTAIL.n355 VTAIL.n354 9.3005
R363 VTAIL.n357 VTAIL.n356 9.3005
R364 VTAIL.n336 VTAIL.n335 9.3005
R365 VTAIL.n364 VTAIL.n363 9.3005
R366 VTAIL.n366 VTAIL.n365 9.3005
R367 VTAIL.n45 VTAIL.n44 9.3005
R368 VTAIL.n4 VTAIL.n3 9.3005
R369 VTAIL.n19 VTAIL.n18 9.3005
R370 VTAIL.n21 VTAIL.n20 9.3005
R371 VTAIL.n12 VTAIL.n11 9.3005
R372 VTAIL.n27 VTAIL.n26 9.3005
R373 VTAIL.n29 VTAIL.n28 9.3005
R374 VTAIL.n8 VTAIL.n7 9.3005
R375 VTAIL.n36 VTAIL.n35 9.3005
R376 VTAIL.n38 VTAIL.n37 9.3005
R377 VTAIL.n91 VTAIL.n90 9.3005
R378 VTAIL.n50 VTAIL.n49 9.3005
R379 VTAIL.n65 VTAIL.n64 9.3005
R380 VTAIL.n67 VTAIL.n66 9.3005
R381 VTAIL.n58 VTAIL.n57 9.3005
R382 VTAIL.n73 VTAIL.n72 9.3005
R383 VTAIL.n75 VTAIL.n74 9.3005
R384 VTAIL.n54 VTAIL.n53 9.3005
R385 VTAIL.n82 VTAIL.n81 9.3005
R386 VTAIL.n84 VTAIL.n83 9.3005
R387 VTAIL.n139 VTAIL.n138 9.3005
R388 VTAIL.n98 VTAIL.n97 9.3005
R389 VTAIL.n113 VTAIL.n112 9.3005
R390 VTAIL.n115 VTAIL.n114 9.3005
R391 VTAIL.n106 VTAIL.n105 9.3005
R392 VTAIL.n121 VTAIL.n120 9.3005
R393 VTAIL.n123 VTAIL.n122 9.3005
R394 VTAIL.n102 VTAIL.n101 9.3005
R395 VTAIL.n130 VTAIL.n129 9.3005
R396 VTAIL.n132 VTAIL.n131 9.3005
R397 VTAIL.n302 VTAIL.n301 9.3005
R398 VTAIL.n304 VTAIL.n303 9.3005
R399 VTAIL.n295 VTAIL.n294 9.3005
R400 VTAIL.n310 VTAIL.n309 9.3005
R401 VTAIL.n312 VTAIL.n311 9.3005
R402 VTAIL.n290 VTAIL.n289 9.3005
R403 VTAIL.n318 VTAIL.n317 9.3005
R404 VTAIL.n320 VTAIL.n319 9.3005
R405 VTAIL.n327 VTAIL.n326 9.3005
R406 VTAIL.n286 VTAIL.n285 9.3005
R407 VTAIL.n254 VTAIL.n253 9.3005
R408 VTAIL.n256 VTAIL.n255 9.3005
R409 VTAIL.n247 VTAIL.n246 9.3005
R410 VTAIL.n262 VTAIL.n261 9.3005
R411 VTAIL.n264 VTAIL.n263 9.3005
R412 VTAIL.n242 VTAIL.n241 9.3005
R413 VTAIL.n270 VTAIL.n269 9.3005
R414 VTAIL.n272 VTAIL.n271 9.3005
R415 VTAIL.n279 VTAIL.n278 9.3005
R416 VTAIL.n238 VTAIL.n237 9.3005
R417 VTAIL.n208 VTAIL.n207 9.3005
R418 VTAIL.n210 VTAIL.n209 9.3005
R419 VTAIL.n201 VTAIL.n200 9.3005
R420 VTAIL.n216 VTAIL.n215 9.3005
R421 VTAIL.n218 VTAIL.n217 9.3005
R422 VTAIL.n196 VTAIL.n195 9.3005
R423 VTAIL.n224 VTAIL.n223 9.3005
R424 VTAIL.n226 VTAIL.n225 9.3005
R425 VTAIL.n233 VTAIL.n232 9.3005
R426 VTAIL.n192 VTAIL.n191 9.3005
R427 VTAIL.n160 VTAIL.n159 9.3005
R428 VTAIL.n162 VTAIL.n161 9.3005
R429 VTAIL.n153 VTAIL.n152 9.3005
R430 VTAIL.n168 VTAIL.n167 9.3005
R431 VTAIL.n170 VTAIL.n169 9.3005
R432 VTAIL.n148 VTAIL.n147 9.3005
R433 VTAIL.n176 VTAIL.n175 9.3005
R434 VTAIL.n178 VTAIL.n177 9.3005
R435 VTAIL.n185 VTAIL.n184 9.3005
R436 VTAIL.n144 VTAIL.n143 9.3005
R437 VTAIL.n350 VTAIL.n340 8.92171
R438 VTAIL.n22 VTAIL.n12 8.92171
R439 VTAIL.n68 VTAIL.n58 8.92171
R440 VTAIL.n116 VTAIL.n106 8.92171
R441 VTAIL.n305 VTAIL.n295 8.92171
R442 VTAIL.n257 VTAIL.n247 8.92171
R443 VTAIL.n211 VTAIL.n201 8.92171
R444 VTAIL.n163 VTAIL.n153 8.92171
R445 VTAIL.n349 VTAIL.n342 8.14595
R446 VTAIL.n21 VTAIL.n14 8.14595
R447 VTAIL.n67 VTAIL.n60 8.14595
R448 VTAIL.n115 VTAIL.n108 8.14595
R449 VTAIL.n304 VTAIL.n297 8.14595
R450 VTAIL.n256 VTAIL.n249 8.14595
R451 VTAIL.n210 VTAIL.n203 8.14595
R452 VTAIL.n162 VTAIL.n155 8.14595
R453 VTAIL.n346 VTAIL.n345 7.3702
R454 VTAIL.n18 VTAIL.n17 7.3702
R455 VTAIL.n64 VTAIL.n63 7.3702
R456 VTAIL.n112 VTAIL.n111 7.3702
R457 VTAIL.n301 VTAIL.n300 7.3702
R458 VTAIL.n253 VTAIL.n252 7.3702
R459 VTAIL.n207 VTAIL.n206 7.3702
R460 VTAIL.n159 VTAIL.n158 7.3702
R461 VTAIL.n346 VTAIL.n342 5.81868
R462 VTAIL.n18 VTAIL.n14 5.81868
R463 VTAIL.n64 VTAIL.n60 5.81868
R464 VTAIL.n112 VTAIL.n108 5.81868
R465 VTAIL.n301 VTAIL.n297 5.81868
R466 VTAIL.n253 VTAIL.n249 5.81868
R467 VTAIL.n207 VTAIL.n203 5.81868
R468 VTAIL.n159 VTAIL.n155 5.81868
R469 VTAIL.n350 VTAIL.n349 5.04292
R470 VTAIL.n22 VTAIL.n21 5.04292
R471 VTAIL.n68 VTAIL.n67 5.04292
R472 VTAIL.n116 VTAIL.n115 5.04292
R473 VTAIL.n305 VTAIL.n304 5.04292
R474 VTAIL.n257 VTAIL.n256 5.04292
R475 VTAIL.n211 VTAIL.n210 5.04292
R476 VTAIL.n163 VTAIL.n162 5.04292
R477 VTAIL.n353 VTAIL.n340 4.26717
R478 VTAIL.n25 VTAIL.n12 4.26717
R479 VTAIL.n71 VTAIL.n58 4.26717
R480 VTAIL.n119 VTAIL.n106 4.26717
R481 VTAIL.n308 VTAIL.n295 4.26717
R482 VTAIL.n260 VTAIL.n247 4.26717
R483 VTAIL.n214 VTAIL.n201 4.26717
R484 VTAIL.n166 VTAIL.n153 4.26717
R485 VTAIL.n354 VTAIL.n338 3.49141
R486 VTAIL.n26 VTAIL.n10 3.49141
R487 VTAIL.n72 VTAIL.n56 3.49141
R488 VTAIL.n120 VTAIL.n104 3.49141
R489 VTAIL.n309 VTAIL.n293 3.49141
R490 VTAIL.n261 VTAIL.n245 3.49141
R491 VTAIL.n215 VTAIL.n199 3.49141
R492 VTAIL.n167 VTAIL.n151 3.49141
R493 VTAIL.n347 VTAIL.n343 2.84303
R494 VTAIL.n19 VTAIL.n15 2.84303
R495 VTAIL.n65 VTAIL.n61 2.84303
R496 VTAIL.n113 VTAIL.n109 2.84303
R497 VTAIL.n302 VTAIL.n298 2.84303
R498 VTAIL.n254 VTAIL.n250 2.84303
R499 VTAIL.n208 VTAIL.n204 2.84303
R500 VTAIL.n160 VTAIL.n156 2.84303
R501 VTAIL.n358 VTAIL.n357 2.71565
R502 VTAIL.n30 VTAIL.n29 2.71565
R503 VTAIL.n76 VTAIL.n75 2.71565
R504 VTAIL.n124 VTAIL.n123 2.71565
R505 VTAIL.n313 VTAIL.n312 2.71565
R506 VTAIL.n265 VTAIL.n264 2.71565
R507 VTAIL.n219 VTAIL.n218 2.71565
R508 VTAIL.n171 VTAIL.n170 2.71565
R509 VTAIL.n0 VTAIL.t1 2.31358
R510 VTAIL.n0 VTAIL.t7 2.31358
R511 VTAIL.n94 VTAIL.t9 2.31358
R512 VTAIL.n94 VTAIL.t15 2.31358
R513 VTAIL.n282 VTAIL.t12 2.31358
R514 VTAIL.n282 VTAIL.t14 2.31358
R515 VTAIL.n188 VTAIL.t4 2.31358
R516 VTAIL.n188 VTAIL.t0 2.31358
R517 VTAIL.n362 VTAIL.n336 1.93989
R518 VTAIL.n374 VTAIL.n330 1.93989
R519 VTAIL.n34 VTAIL.n8 1.93989
R520 VTAIL.n46 VTAIL.n2 1.93989
R521 VTAIL.n80 VTAIL.n54 1.93989
R522 VTAIL.n92 VTAIL.n48 1.93989
R523 VTAIL.n128 VTAIL.n102 1.93989
R524 VTAIL.n140 VTAIL.n96 1.93989
R525 VTAIL.n328 VTAIL.n284 1.93989
R526 VTAIL.n316 VTAIL.n290 1.93989
R527 VTAIL.n280 VTAIL.n236 1.93989
R528 VTAIL.n268 VTAIL.n242 1.93989
R529 VTAIL.n234 VTAIL.n190 1.93989
R530 VTAIL.n222 VTAIL.n196 1.93989
R531 VTAIL.n186 VTAIL.n142 1.93989
R532 VTAIL.n174 VTAIL.n148 1.93989
R533 VTAIL.n189 VTAIL.n187 1.17291
R534 VTAIL.n235 VTAIL.n189 1.17291
R535 VTAIL.n283 VTAIL.n281 1.17291
R536 VTAIL.n329 VTAIL.n283 1.17291
R537 VTAIL.n141 VTAIL.n95 1.17291
R538 VTAIL.n95 VTAIL.n93 1.17291
R539 VTAIL.n47 VTAIL.n1 1.17291
R540 VTAIL.n363 VTAIL.n334 1.16414
R541 VTAIL.n372 VTAIL.n371 1.16414
R542 VTAIL.n35 VTAIL.n6 1.16414
R543 VTAIL.n44 VTAIL.n43 1.16414
R544 VTAIL.n81 VTAIL.n52 1.16414
R545 VTAIL.n90 VTAIL.n89 1.16414
R546 VTAIL.n129 VTAIL.n100 1.16414
R547 VTAIL.n138 VTAIL.n137 1.16414
R548 VTAIL.n326 VTAIL.n325 1.16414
R549 VTAIL.n317 VTAIL.n288 1.16414
R550 VTAIL.n278 VTAIL.n277 1.16414
R551 VTAIL.n269 VTAIL.n240 1.16414
R552 VTAIL.n232 VTAIL.n231 1.16414
R553 VTAIL.n223 VTAIL.n194 1.16414
R554 VTAIL.n184 VTAIL.n183 1.16414
R555 VTAIL.n175 VTAIL.n146 1.16414
R556 VTAIL VTAIL.n375 1.11472
R557 VTAIL.n281 VTAIL.n235 0.470328
R558 VTAIL.n93 VTAIL.n47 0.470328
R559 VTAIL.n367 VTAIL.n366 0.388379
R560 VTAIL.n368 VTAIL.n332 0.388379
R561 VTAIL.n39 VTAIL.n38 0.388379
R562 VTAIL.n40 VTAIL.n4 0.388379
R563 VTAIL.n85 VTAIL.n84 0.388379
R564 VTAIL.n86 VTAIL.n50 0.388379
R565 VTAIL.n133 VTAIL.n132 0.388379
R566 VTAIL.n134 VTAIL.n98 0.388379
R567 VTAIL.n322 VTAIL.n286 0.388379
R568 VTAIL.n321 VTAIL.n320 0.388379
R569 VTAIL.n274 VTAIL.n238 0.388379
R570 VTAIL.n273 VTAIL.n272 0.388379
R571 VTAIL.n228 VTAIL.n192 0.388379
R572 VTAIL.n227 VTAIL.n226 0.388379
R573 VTAIL.n180 VTAIL.n144 0.388379
R574 VTAIL.n179 VTAIL.n178 0.388379
R575 VTAIL.n348 VTAIL.n347 0.155672
R576 VTAIL.n348 VTAIL.n339 0.155672
R577 VTAIL.n355 VTAIL.n339 0.155672
R578 VTAIL.n356 VTAIL.n355 0.155672
R579 VTAIL.n356 VTAIL.n335 0.155672
R580 VTAIL.n364 VTAIL.n335 0.155672
R581 VTAIL.n365 VTAIL.n364 0.155672
R582 VTAIL.n365 VTAIL.n331 0.155672
R583 VTAIL.n373 VTAIL.n331 0.155672
R584 VTAIL.n20 VTAIL.n19 0.155672
R585 VTAIL.n20 VTAIL.n11 0.155672
R586 VTAIL.n27 VTAIL.n11 0.155672
R587 VTAIL.n28 VTAIL.n27 0.155672
R588 VTAIL.n28 VTAIL.n7 0.155672
R589 VTAIL.n36 VTAIL.n7 0.155672
R590 VTAIL.n37 VTAIL.n36 0.155672
R591 VTAIL.n37 VTAIL.n3 0.155672
R592 VTAIL.n45 VTAIL.n3 0.155672
R593 VTAIL.n66 VTAIL.n65 0.155672
R594 VTAIL.n66 VTAIL.n57 0.155672
R595 VTAIL.n73 VTAIL.n57 0.155672
R596 VTAIL.n74 VTAIL.n73 0.155672
R597 VTAIL.n74 VTAIL.n53 0.155672
R598 VTAIL.n82 VTAIL.n53 0.155672
R599 VTAIL.n83 VTAIL.n82 0.155672
R600 VTAIL.n83 VTAIL.n49 0.155672
R601 VTAIL.n91 VTAIL.n49 0.155672
R602 VTAIL.n114 VTAIL.n113 0.155672
R603 VTAIL.n114 VTAIL.n105 0.155672
R604 VTAIL.n121 VTAIL.n105 0.155672
R605 VTAIL.n122 VTAIL.n121 0.155672
R606 VTAIL.n122 VTAIL.n101 0.155672
R607 VTAIL.n130 VTAIL.n101 0.155672
R608 VTAIL.n131 VTAIL.n130 0.155672
R609 VTAIL.n131 VTAIL.n97 0.155672
R610 VTAIL.n139 VTAIL.n97 0.155672
R611 VTAIL.n327 VTAIL.n285 0.155672
R612 VTAIL.n319 VTAIL.n285 0.155672
R613 VTAIL.n319 VTAIL.n318 0.155672
R614 VTAIL.n318 VTAIL.n289 0.155672
R615 VTAIL.n311 VTAIL.n289 0.155672
R616 VTAIL.n311 VTAIL.n310 0.155672
R617 VTAIL.n310 VTAIL.n294 0.155672
R618 VTAIL.n303 VTAIL.n294 0.155672
R619 VTAIL.n303 VTAIL.n302 0.155672
R620 VTAIL.n279 VTAIL.n237 0.155672
R621 VTAIL.n271 VTAIL.n237 0.155672
R622 VTAIL.n271 VTAIL.n270 0.155672
R623 VTAIL.n270 VTAIL.n241 0.155672
R624 VTAIL.n263 VTAIL.n241 0.155672
R625 VTAIL.n263 VTAIL.n262 0.155672
R626 VTAIL.n262 VTAIL.n246 0.155672
R627 VTAIL.n255 VTAIL.n246 0.155672
R628 VTAIL.n255 VTAIL.n254 0.155672
R629 VTAIL.n233 VTAIL.n191 0.155672
R630 VTAIL.n225 VTAIL.n191 0.155672
R631 VTAIL.n225 VTAIL.n224 0.155672
R632 VTAIL.n224 VTAIL.n195 0.155672
R633 VTAIL.n217 VTAIL.n195 0.155672
R634 VTAIL.n217 VTAIL.n216 0.155672
R635 VTAIL.n216 VTAIL.n200 0.155672
R636 VTAIL.n209 VTAIL.n200 0.155672
R637 VTAIL.n209 VTAIL.n208 0.155672
R638 VTAIL.n185 VTAIL.n143 0.155672
R639 VTAIL.n177 VTAIL.n143 0.155672
R640 VTAIL.n177 VTAIL.n176 0.155672
R641 VTAIL.n176 VTAIL.n147 0.155672
R642 VTAIL.n169 VTAIL.n147 0.155672
R643 VTAIL.n169 VTAIL.n168 0.155672
R644 VTAIL.n168 VTAIL.n152 0.155672
R645 VTAIL.n161 VTAIL.n152 0.155672
R646 VTAIL.n161 VTAIL.n160 0.155672
R647 VTAIL VTAIL.n1 0.0586897
R648 B.n602 B.n601 585
R649 B.n603 B.n602 585
R650 B.n238 B.n91 585
R651 B.n237 B.n236 585
R652 B.n235 B.n234 585
R653 B.n233 B.n232 585
R654 B.n231 B.n230 585
R655 B.n229 B.n228 585
R656 B.n227 B.n226 585
R657 B.n225 B.n224 585
R658 B.n223 B.n222 585
R659 B.n221 B.n220 585
R660 B.n219 B.n218 585
R661 B.n217 B.n216 585
R662 B.n215 B.n214 585
R663 B.n213 B.n212 585
R664 B.n211 B.n210 585
R665 B.n209 B.n208 585
R666 B.n207 B.n206 585
R667 B.n205 B.n204 585
R668 B.n203 B.n202 585
R669 B.n201 B.n200 585
R670 B.n199 B.n198 585
R671 B.n197 B.n196 585
R672 B.n195 B.n194 585
R673 B.n193 B.n192 585
R674 B.n191 B.n190 585
R675 B.n189 B.n188 585
R676 B.n187 B.n186 585
R677 B.n185 B.n184 585
R678 B.n183 B.n182 585
R679 B.n181 B.n180 585
R680 B.n179 B.n178 585
R681 B.n176 B.n175 585
R682 B.n174 B.n173 585
R683 B.n172 B.n171 585
R684 B.n170 B.n169 585
R685 B.n168 B.n167 585
R686 B.n166 B.n165 585
R687 B.n164 B.n163 585
R688 B.n162 B.n161 585
R689 B.n160 B.n159 585
R690 B.n158 B.n157 585
R691 B.n156 B.n155 585
R692 B.n154 B.n153 585
R693 B.n152 B.n151 585
R694 B.n150 B.n149 585
R695 B.n148 B.n147 585
R696 B.n146 B.n145 585
R697 B.n144 B.n143 585
R698 B.n142 B.n141 585
R699 B.n140 B.n139 585
R700 B.n138 B.n137 585
R701 B.n136 B.n135 585
R702 B.n134 B.n133 585
R703 B.n132 B.n131 585
R704 B.n130 B.n129 585
R705 B.n128 B.n127 585
R706 B.n126 B.n125 585
R707 B.n124 B.n123 585
R708 B.n122 B.n121 585
R709 B.n120 B.n119 585
R710 B.n118 B.n117 585
R711 B.n116 B.n115 585
R712 B.n114 B.n113 585
R713 B.n112 B.n111 585
R714 B.n110 B.n109 585
R715 B.n108 B.n107 585
R716 B.n106 B.n105 585
R717 B.n104 B.n103 585
R718 B.n102 B.n101 585
R719 B.n100 B.n99 585
R720 B.n98 B.n97 585
R721 B.n53 B.n52 585
R722 B.n600 B.n54 585
R723 B.n604 B.n54 585
R724 B.n599 B.n598 585
R725 B.n598 B.n50 585
R726 B.n597 B.n49 585
R727 B.n610 B.n49 585
R728 B.n596 B.n48 585
R729 B.n611 B.n48 585
R730 B.n595 B.n47 585
R731 B.n612 B.n47 585
R732 B.n594 B.n593 585
R733 B.n593 B.n46 585
R734 B.n592 B.n42 585
R735 B.n618 B.n42 585
R736 B.n591 B.n41 585
R737 B.n619 B.n41 585
R738 B.n590 B.n40 585
R739 B.n620 B.n40 585
R740 B.n589 B.n588 585
R741 B.n588 B.n36 585
R742 B.n587 B.n35 585
R743 B.n626 B.n35 585
R744 B.n586 B.n34 585
R745 B.n627 B.n34 585
R746 B.n585 B.n33 585
R747 B.n628 B.n33 585
R748 B.n584 B.n583 585
R749 B.n583 B.n29 585
R750 B.n582 B.n28 585
R751 B.n634 B.n28 585
R752 B.n581 B.n27 585
R753 B.n635 B.n27 585
R754 B.n580 B.n26 585
R755 B.n636 B.n26 585
R756 B.n579 B.n578 585
R757 B.n578 B.n22 585
R758 B.n577 B.n21 585
R759 B.n642 B.n21 585
R760 B.n576 B.n20 585
R761 B.n643 B.n20 585
R762 B.n575 B.n19 585
R763 B.n644 B.n19 585
R764 B.n574 B.n573 585
R765 B.n573 B.n15 585
R766 B.n572 B.n14 585
R767 B.n650 B.n14 585
R768 B.n571 B.n13 585
R769 B.n651 B.n13 585
R770 B.n570 B.n12 585
R771 B.n652 B.n12 585
R772 B.n569 B.n568 585
R773 B.n568 B.n8 585
R774 B.n567 B.n7 585
R775 B.n658 B.n7 585
R776 B.n566 B.n6 585
R777 B.n659 B.n6 585
R778 B.n565 B.n5 585
R779 B.n660 B.n5 585
R780 B.n564 B.n563 585
R781 B.n563 B.n4 585
R782 B.n562 B.n239 585
R783 B.n562 B.n561 585
R784 B.n552 B.n240 585
R785 B.n241 B.n240 585
R786 B.n554 B.n553 585
R787 B.n555 B.n554 585
R788 B.n551 B.n246 585
R789 B.n246 B.n245 585
R790 B.n550 B.n549 585
R791 B.n549 B.n548 585
R792 B.n248 B.n247 585
R793 B.n249 B.n248 585
R794 B.n541 B.n540 585
R795 B.n542 B.n541 585
R796 B.n539 B.n254 585
R797 B.n254 B.n253 585
R798 B.n538 B.n537 585
R799 B.n537 B.n536 585
R800 B.n256 B.n255 585
R801 B.n257 B.n256 585
R802 B.n529 B.n528 585
R803 B.n530 B.n529 585
R804 B.n527 B.n262 585
R805 B.n262 B.n261 585
R806 B.n526 B.n525 585
R807 B.n525 B.n524 585
R808 B.n264 B.n263 585
R809 B.n265 B.n264 585
R810 B.n517 B.n516 585
R811 B.n518 B.n517 585
R812 B.n515 B.n270 585
R813 B.n270 B.n269 585
R814 B.n514 B.n513 585
R815 B.n513 B.n512 585
R816 B.n272 B.n271 585
R817 B.n273 B.n272 585
R818 B.n505 B.n504 585
R819 B.n506 B.n505 585
R820 B.n503 B.n278 585
R821 B.n278 B.n277 585
R822 B.n502 B.n501 585
R823 B.n501 B.n500 585
R824 B.n280 B.n279 585
R825 B.n493 B.n280 585
R826 B.n492 B.n491 585
R827 B.n494 B.n492 585
R828 B.n490 B.n285 585
R829 B.n285 B.n284 585
R830 B.n489 B.n488 585
R831 B.n488 B.n487 585
R832 B.n287 B.n286 585
R833 B.n288 B.n287 585
R834 B.n480 B.n479 585
R835 B.n481 B.n480 585
R836 B.n291 B.n290 585
R837 B.n335 B.n333 585
R838 B.n336 B.n332 585
R839 B.n336 B.n292 585
R840 B.n339 B.n338 585
R841 B.n340 B.n331 585
R842 B.n342 B.n341 585
R843 B.n344 B.n330 585
R844 B.n347 B.n346 585
R845 B.n348 B.n329 585
R846 B.n350 B.n349 585
R847 B.n352 B.n328 585
R848 B.n355 B.n354 585
R849 B.n356 B.n327 585
R850 B.n358 B.n357 585
R851 B.n360 B.n326 585
R852 B.n363 B.n362 585
R853 B.n364 B.n325 585
R854 B.n366 B.n365 585
R855 B.n368 B.n324 585
R856 B.n371 B.n370 585
R857 B.n372 B.n323 585
R858 B.n374 B.n373 585
R859 B.n376 B.n322 585
R860 B.n379 B.n378 585
R861 B.n380 B.n321 585
R862 B.n382 B.n381 585
R863 B.n384 B.n320 585
R864 B.n387 B.n386 585
R865 B.n388 B.n319 585
R866 B.n390 B.n389 585
R867 B.n392 B.n318 585
R868 B.n395 B.n394 585
R869 B.n397 B.n315 585
R870 B.n399 B.n398 585
R871 B.n401 B.n314 585
R872 B.n404 B.n403 585
R873 B.n405 B.n313 585
R874 B.n407 B.n406 585
R875 B.n409 B.n312 585
R876 B.n412 B.n411 585
R877 B.n413 B.n309 585
R878 B.n416 B.n415 585
R879 B.n418 B.n308 585
R880 B.n421 B.n420 585
R881 B.n422 B.n307 585
R882 B.n424 B.n423 585
R883 B.n426 B.n306 585
R884 B.n429 B.n428 585
R885 B.n430 B.n305 585
R886 B.n432 B.n431 585
R887 B.n434 B.n304 585
R888 B.n437 B.n436 585
R889 B.n438 B.n303 585
R890 B.n440 B.n439 585
R891 B.n442 B.n302 585
R892 B.n445 B.n444 585
R893 B.n446 B.n301 585
R894 B.n448 B.n447 585
R895 B.n450 B.n300 585
R896 B.n453 B.n452 585
R897 B.n454 B.n299 585
R898 B.n456 B.n455 585
R899 B.n458 B.n298 585
R900 B.n461 B.n460 585
R901 B.n462 B.n297 585
R902 B.n464 B.n463 585
R903 B.n466 B.n296 585
R904 B.n469 B.n468 585
R905 B.n470 B.n295 585
R906 B.n472 B.n471 585
R907 B.n474 B.n294 585
R908 B.n477 B.n476 585
R909 B.n478 B.n293 585
R910 B.n483 B.n482 585
R911 B.n482 B.n481 585
R912 B.n484 B.n289 585
R913 B.n289 B.n288 585
R914 B.n486 B.n485 585
R915 B.n487 B.n486 585
R916 B.n283 B.n282 585
R917 B.n284 B.n283 585
R918 B.n496 B.n495 585
R919 B.n495 B.n494 585
R920 B.n497 B.n281 585
R921 B.n493 B.n281 585
R922 B.n499 B.n498 585
R923 B.n500 B.n499 585
R924 B.n276 B.n275 585
R925 B.n277 B.n276 585
R926 B.n508 B.n507 585
R927 B.n507 B.n506 585
R928 B.n509 B.n274 585
R929 B.n274 B.n273 585
R930 B.n511 B.n510 585
R931 B.n512 B.n511 585
R932 B.n268 B.n267 585
R933 B.n269 B.n268 585
R934 B.n520 B.n519 585
R935 B.n519 B.n518 585
R936 B.n521 B.n266 585
R937 B.n266 B.n265 585
R938 B.n523 B.n522 585
R939 B.n524 B.n523 585
R940 B.n260 B.n259 585
R941 B.n261 B.n260 585
R942 B.n532 B.n531 585
R943 B.n531 B.n530 585
R944 B.n533 B.n258 585
R945 B.n258 B.n257 585
R946 B.n535 B.n534 585
R947 B.n536 B.n535 585
R948 B.n252 B.n251 585
R949 B.n253 B.n252 585
R950 B.n544 B.n543 585
R951 B.n543 B.n542 585
R952 B.n545 B.n250 585
R953 B.n250 B.n249 585
R954 B.n547 B.n546 585
R955 B.n548 B.n547 585
R956 B.n244 B.n243 585
R957 B.n245 B.n244 585
R958 B.n557 B.n556 585
R959 B.n556 B.n555 585
R960 B.n558 B.n242 585
R961 B.n242 B.n241 585
R962 B.n560 B.n559 585
R963 B.n561 B.n560 585
R964 B.n2 B.n0 585
R965 B.n4 B.n2 585
R966 B.n3 B.n1 585
R967 B.n659 B.n3 585
R968 B.n657 B.n656 585
R969 B.n658 B.n657 585
R970 B.n655 B.n9 585
R971 B.n9 B.n8 585
R972 B.n654 B.n653 585
R973 B.n653 B.n652 585
R974 B.n11 B.n10 585
R975 B.n651 B.n11 585
R976 B.n649 B.n648 585
R977 B.n650 B.n649 585
R978 B.n647 B.n16 585
R979 B.n16 B.n15 585
R980 B.n646 B.n645 585
R981 B.n645 B.n644 585
R982 B.n18 B.n17 585
R983 B.n643 B.n18 585
R984 B.n641 B.n640 585
R985 B.n642 B.n641 585
R986 B.n639 B.n23 585
R987 B.n23 B.n22 585
R988 B.n638 B.n637 585
R989 B.n637 B.n636 585
R990 B.n25 B.n24 585
R991 B.n635 B.n25 585
R992 B.n633 B.n632 585
R993 B.n634 B.n633 585
R994 B.n631 B.n30 585
R995 B.n30 B.n29 585
R996 B.n630 B.n629 585
R997 B.n629 B.n628 585
R998 B.n32 B.n31 585
R999 B.n627 B.n32 585
R1000 B.n625 B.n624 585
R1001 B.n626 B.n625 585
R1002 B.n623 B.n37 585
R1003 B.n37 B.n36 585
R1004 B.n622 B.n621 585
R1005 B.n621 B.n620 585
R1006 B.n39 B.n38 585
R1007 B.n619 B.n39 585
R1008 B.n617 B.n616 585
R1009 B.n618 B.n617 585
R1010 B.n615 B.n43 585
R1011 B.n46 B.n43 585
R1012 B.n614 B.n613 585
R1013 B.n613 B.n612 585
R1014 B.n45 B.n44 585
R1015 B.n611 B.n45 585
R1016 B.n609 B.n608 585
R1017 B.n610 B.n609 585
R1018 B.n607 B.n51 585
R1019 B.n51 B.n50 585
R1020 B.n606 B.n605 585
R1021 B.n605 B.n604 585
R1022 B.n662 B.n661 585
R1023 B.n661 B.n660 585
R1024 B.n482 B.n291 482.89
R1025 B.n605 B.n53 482.89
R1026 B.n480 B.n293 482.89
R1027 B.n602 B.n54 482.89
R1028 B.n310 B.t7 403.413
R1029 B.n316 B.t11 403.413
R1030 B.n94 B.t18 403.413
R1031 B.n92 B.t14 403.413
R1032 B.n603 B.n90 256.663
R1033 B.n603 B.n89 256.663
R1034 B.n603 B.n88 256.663
R1035 B.n603 B.n87 256.663
R1036 B.n603 B.n86 256.663
R1037 B.n603 B.n85 256.663
R1038 B.n603 B.n84 256.663
R1039 B.n603 B.n83 256.663
R1040 B.n603 B.n82 256.663
R1041 B.n603 B.n81 256.663
R1042 B.n603 B.n80 256.663
R1043 B.n603 B.n79 256.663
R1044 B.n603 B.n78 256.663
R1045 B.n603 B.n77 256.663
R1046 B.n603 B.n76 256.663
R1047 B.n603 B.n75 256.663
R1048 B.n603 B.n74 256.663
R1049 B.n603 B.n73 256.663
R1050 B.n603 B.n72 256.663
R1051 B.n603 B.n71 256.663
R1052 B.n603 B.n70 256.663
R1053 B.n603 B.n69 256.663
R1054 B.n603 B.n68 256.663
R1055 B.n603 B.n67 256.663
R1056 B.n603 B.n66 256.663
R1057 B.n603 B.n65 256.663
R1058 B.n603 B.n64 256.663
R1059 B.n603 B.n63 256.663
R1060 B.n603 B.n62 256.663
R1061 B.n603 B.n61 256.663
R1062 B.n603 B.n60 256.663
R1063 B.n603 B.n59 256.663
R1064 B.n603 B.n58 256.663
R1065 B.n603 B.n57 256.663
R1066 B.n603 B.n56 256.663
R1067 B.n603 B.n55 256.663
R1068 B.n334 B.n292 256.663
R1069 B.n337 B.n292 256.663
R1070 B.n343 B.n292 256.663
R1071 B.n345 B.n292 256.663
R1072 B.n351 B.n292 256.663
R1073 B.n353 B.n292 256.663
R1074 B.n359 B.n292 256.663
R1075 B.n361 B.n292 256.663
R1076 B.n367 B.n292 256.663
R1077 B.n369 B.n292 256.663
R1078 B.n375 B.n292 256.663
R1079 B.n377 B.n292 256.663
R1080 B.n383 B.n292 256.663
R1081 B.n385 B.n292 256.663
R1082 B.n391 B.n292 256.663
R1083 B.n393 B.n292 256.663
R1084 B.n400 B.n292 256.663
R1085 B.n402 B.n292 256.663
R1086 B.n408 B.n292 256.663
R1087 B.n410 B.n292 256.663
R1088 B.n417 B.n292 256.663
R1089 B.n419 B.n292 256.663
R1090 B.n425 B.n292 256.663
R1091 B.n427 B.n292 256.663
R1092 B.n433 B.n292 256.663
R1093 B.n435 B.n292 256.663
R1094 B.n441 B.n292 256.663
R1095 B.n443 B.n292 256.663
R1096 B.n449 B.n292 256.663
R1097 B.n451 B.n292 256.663
R1098 B.n457 B.n292 256.663
R1099 B.n459 B.n292 256.663
R1100 B.n465 B.n292 256.663
R1101 B.n467 B.n292 256.663
R1102 B.n473 B.n292 256.663
R1103 B.n475 B.n292 256.663
R1104 B.n310 B.t10 249.048
R1105 B.n92 B.t16 249.048
R1106 B.n316 B.t13 249.048
R1107 B.n94 B.t19 249.048
R1108 B.n311 B.t9 222.673
R1109 B.n93 B.t17 222.673
R1110 B.n317 B.t12 222.673
R1111 B.n95 B.t20 222.673
R1112 B.n482 B.n289 163.367
R1113 B.n486 B.n289 163.367
R1114 B.n486 B.n283 163.367
R1115 B.n495 B.n283 163.367
R1116 B.n495 B.n281 163.367
R1117 B.n499 B.n281 163.367
R1118 B.n499 B.n276 163.367
R1119 B.n507 B.n276 163.367
R1120 B.n507 B.n274 163.367
R1121 B.n511 B.n274 163.367
R1122 B.n511 B.n268 163.367
R1123 B.n519 B.n268 163.367
R1124 B.n519 B.n266 163.367
R1125 B.n523 B.n266 163.367
R1126 B.n523 B.n260 163.367
R1127 B.n531 B.n260 163.367
R1128 B.n531 B.n258 163.367
R1129 B.n535 B.n258 163.367
R1130 B.n535 B.n252 163.367
R1131 B.n543 B.n252 163.367
R1132 B.n543 B.n250 163.367
R1133 B.n547 B.n250 163.367
R1134 B.n547 B.n244 163.367
R1135 B.n556 B.n244 163.367
R1136 B.n556 B.n242 163.367
R1137 B.n560 B.n242 163.367
R1138 B.n560 B.n2 163.367
R1139 B.n661 B.n2 163.367
R1140 B.n661 B.n3 163.367
R1141 B.n657 B.n3 163.367
R1142 B.n657 B.n9 163.367
R1143 B.n653 B.n9 163.367
R1144 B.n653 B.n11 163.367
R1145 B.n649 B.n11 163.367
R1146 B.n649 B.n16 163.367
R1147 B.n645 B.n16 163.367
R1148 B.n645 B.n18 163.367
R1149 B.n641 B.n18 163.367
R1150 B.n641 B.n23 163.367
R1151 B.n637 B.n23 163.367
R1152 B.n637 B.n25 163.367
R1153 B.n633 B.n25 163.367
R1154 B.n633 B.n30 163.367
R1155 B.n629 B.n30 163.367
R1156 B.n629 B.n32 163.367
R1157 B.n625 B.n32 163.367
R1158 B.n625 B.n37 163.367
R1159 B.n621 B.n37 163.367
R1160 B.n621 B.n39 163.367
R1161 B.n617 B.n39 163.367
R1162 B.n617 B.n43 163.367
R1163 B.n613 B.n43 163.367
R1164 B.n613 B.n45 163.367
R1165 B.n609 B.n45 163.367
R1166 B.n609 B.n51 163.367
R1167 B.n605 B.n51 163.367
R1168 B.n336 B.n335 163.367
R1169 B.n338 B.n336 163.367
R1170 B.n342 B.n331 163.367
R1171 B.n346 B.n344 163.367
R1172 B.n350 B.n329 163.367
R1173 B.n354 B.n352 163.367
R1174 B.n358 B.n327 163.367
R1175 B.n362 B.n360 163.367
R1176 B.n366 B.n325 163.367
R1177 B.n370 B.n368 163.367
R1178 B.n374 B.n323 163.367
R1179 B.n378 B.n376 163.367
R1180 B.n382 B.n321 163.367
R1181 B.n386 B.n384 163.367
R1182 B.n390 B.n319 163.367
R1183 B.n394 B.n392 163.367
R1184 B.n399 B.n315 163.367
R1185 B.n403 B.n401 163.367
R1186 B.n407 B.n313 163.367
R1187 B.n411 B.n409 163.367
R1188 B.n416 B.n309 163.367
R1189 B.n420 B.n418 163.367
R1190 B.n424 B.n307 163.367
R1191 B.n428 B.n426 163.367
R1192 B.n432 B.n305 163.367
R1193 B.n436 B.n434 163.367
R1194 B.n440 B.n303 163.367
R1195 B.n444 B.n442 163.367
R1196 B.n448 B.n301 163.367
R1197 B.n452 B.n450 163.367
R1198 B.n456 B.n299 163.367
R1199 B.n460 B.n458 163.367
R1200 B.n464 B.n297 163.367
R1201 B.n468 B.n466 163.367
R1202 B.n472 B.n295 163.367
R1203 B.n476 B.n474 163.367
R1204 B.n480 B.n287 163.367
R1205 B.n488 B.n287 163.367
R1206 B.n488 B.n285 163.367
R1207 B.n492 B.n285 163.367
R1208 B.n492 B.n280 163.367
R1209 B.n501 B.n280 163.367
R1210 B.n501 B.n278 163.367
R1211 B.n505 B.n278 163.367
R1212 B.n505 B.n272 163.367
R1213 B.n513 B.n272 163.367
R1214 B.n513 B.n270 163.367
R1215 B.n517 B.n270 163.367
R1216 B.n517 B.n264 163.367
R1217 B.n525 B.n264 163.367
R1218 B.n525 B.n262 163.367
R1219 B.n529 B.n262 163.367
R1220 B.n529 B.n256 163.367
R1221 B.n537 B.n256 163.367
R1222 B.n537 B.n254 163.367
R1223 B.n541 B.n254 163.367
R1224 B.n541 B.n248 163.367
R1225 B.n549 B.n248 163.367
R1226 B.n549 B.n246 163.367
R1227 B.n554 B.n246 163.367
R1228 B.n554 B.n240 163.367
R1229 B.n562 B.n240 163.367
R1230 B.n563 B.n562 163.367
R1231 B.n563 B.n5 163.367
R1232 B.n6 B.n5 163.367
R1233 B.n7 B.n6 163.367
R1234 B.n568 B.n7 163.367
R1235 B.n568 B.n12 163.367
R1236 B.n13 B.n12 163.367
R1237 B.n14 B.n13 163.367
R1238 B.n573 B.n14 163.367
R1239 B.n573 B.n19 163.367
R1240 B.n20 B.n19 163.367
R1241 B.n21 B.n20 163.367
R1242 B.n578 B.n21 163.367
R1243 B.n578 B.n26 163.367
R1244 B.n27 B.n26 163.367
R1245 B.n28 B.n27 163.367
R1246 B.n583 B.n28 163.367
R1247 B.n583 B.n33 163.367
R1248 B.n34 B.n33 163.367
R1249 B.n35 B.n34 163.367
R1250 B.n588 B.n35 163.367
R1251 B.n588 B.n40 163.367
R1252 B.n41 B.n40 163.367
R1253 B.n42 B.n41 163.367
R1254 B.n593 B.n42 163.367
R1255 B.n593 B.n47 163.367
R1256 B.n48 B.n47 163.367
R1257 B.n49 B.n48 163.367
R1258 B.n598 B.n49 163.367
R1259 B.n598 B.n54 163.367
R1260 B.n99 B.n98 163.367
R1261 B.n103 B.n102 163.367
R1262 B.n107 B.n106 163.367
R1263 B.n111 B.n110 163.367
R1264 B.n115 B.n114 163.367
R1265 B.n119 B.n118 163.367
R1266 B.n123 B.n122 163.367
R1267 B.n127 B.n126 163.367
R1268 B.n131 B.n130 163.367
R1269 B.n135 B.n134 163.367
R1270 B.n139 B.n138 163.367
R1271 B.n143 B.n142 163.367
R1272 B.n147 B.n146 163.367
R1273 B.n151 B.n150 163.367
R1274 B.n155 B.n154 163.367
R1275 B.n159 B.n158 163.367
R1276 B.n163 B.n162 163.367
R1277 B.n167 B.n166 163.367
R1278 B.n171 B.n170 163.367
R1279 B.n175 B.n174 163.367
R1280 B.n180 B.n179 163.367
R1281 B.n184 B.n183 163.367
R1282 B.n188 B.n187 163.367
R1283 B.n192 B.n191 163.367
R1284 B.n196 B.n195 163.367
R1285 B.n200 B.n199 163.367
R1286 B.n204 B.n203 163.367
R1287 B.n208 B.n207 163.367
R1288 B.n212 B.n211 163.367
R1289 B.n216 B.n215 163.367
R1290 B.n220 B.n219 163.367
R1291 B.n224 B.n223 163.367
R1292 B.n228 B.n227 163.367
R1293 B.n232 B.n231 163.367
R1294 B.n236 B.n235 163.367
R1295 B.n602 B.n91 163.367
R1296 B.n481 B.n292 104.156
R1297 B.n604 B.n603 104.156
R1298 B.n334 B.n291 71.676
R1299 B.n338 B.n337 71.676
R1300 B.n343 B.n342 71.676
R1301 B.n346 B.n345 71.676
R1302 B.n351 B.n350 71.676
R1303 B.n354 B.n353 71.676
R1304 B.n359 B.n358 71.676
R1305 B.n362 B.n361 71.676
R1306 B.n367 B.n366 71.676
R1307 B.n370 B.n369 71.676
R1308 B.n375 B.n374 71.676
R1309 B.n378 B.n377 71.676
R1310 B.n383 B.n382 71.676
R1311 B.n386 B.n385 71.676
R1312 B.n391 B.n390 71.676
R1313 B.n394 B.n393 71.676
R1314 B.n400 B.n399 71.676
R1315 B.n403 B.n402 71.676
R1316 B.n408 B.n407 71.676
R1317 B.n411 B.n410 71.676
R1318 B.n417 B.n416 71.676
R1319 B.n420 B.n419 71.676
R1320 B.n425 B.n424 71.676
R1321 B.n428 B.n427 71.676
R1322 B.n433 B.n432 71.676
R1323 B.n436 B.n435 71.676
R1324 B.n441 B.n440 71.676
R1325 B.n444 B.n443 71.676
R1326 B.n449 B.n448 71.676
R1327 B.n452 B.n451 71.676
R1328 B.n457 B.n456 71.676
R1329 B.n460 B.n459 71.676
R1330 B.n465 B.n464 71.676
R1331 B.n468 B.n467 71.676
R1332 B.n473 B.n472 71.676
R1333 B.n476 B.n475 71.676
R1334 B.n55 B.n53 71.676
R1335 B.n99 B.n56 71.676
R1336 B.n103 B.n57 71.676
R1337 B.n107 B.n58 71.676
R1338 B.n111 B.n59 71.676
R1339 B.n115 B.n60 71.676
R1340 B.n119 B.n61 71.676
R1341 B.n123 B.n62 71.676
R1342 B.n127 B.n63 71.676
R1343 B.n131 B.n64 71.676
R1344 B.n135 B.n65 71.676
R1345 B.n139 B.n66 71.676
R1346 B.n143 B.n67 71.676
R1347 B.n147 B.n68 71.676
R1348 B.n151 B.n69 71.676
R1349 B.n155 B.n70 71.676
R1350 B.n159 B.n71 71.676
R1351 B.n163 B.n72 71.676
R1352 B.n167 B.n73 71.676
R1353 B.n171 B.n74 71.676
R1354 B.n175 B.n75 71.676
R1355 B.n180 B.n76 71.676
R1356 B.n184 B.n77 71.676
R1357 B.n188 B.n78 71.676
R1358 B.n192 B.n79 71.676
R1359 B.n196 B.n80 71.676
R1360 B.n200 B.n81 71.676
R1361 B.n204 B.n82 71.676
R1362 B.n208 B.n83 71.676
R1363 B.n212 B.n84 71.676
R1364 B.n216 B.n85 71.676
R1365 B.n220 B.n86 71.676
R1366 B.n224 B.n87 71.676
R1367 B.n228 B.n88 71.676
R1368 B.n232 B.n89 71.676
R1369 B.n236 B.n90 71.676
R1370 B.n91 B.n90 71.676
R1371 B.n235 B.n89 71.676
R1372 B.n231 B.n88 71.676
R1373 B.n227 B.n87 71.676
R1374 B.n223 B.n86 71.676
R1375 B.n219 B.n85 71.676
R1376 B.n215 B.n84 71.676
R1377 B.n211 B.n83 71.676
R1378 B.n207 B.n82 71.676
R1379 B.n203 B.n81 71.676
R1380 B.n199 B.n80 71.676
R1381 B.n195 B.n79 71.676
R1382 B.n191 B.n78 71.676
R1383 B.n187 B.n77 71.676
R1384 B.n183 B.n76 71.676
R1385 B.n179 B.n75 71.676
R1386 B.n174 B.n74 71.676
R1387 B.n170 B.n73 71.676
R1388 B.n166 B.n72 71.676
R1389 B.n162 B.n71 71.676
R1390 B.n158 B.n70 71.676
R1391 B.n154 B.n69 71.676
R1392 B.n150 B.n68 71.676
R1393 B.n146 B.n67 71.676
R1394 B.n142 B.n66 71.676
R1395 B.n138 B.n65 71.676
R1396 B.n134 B.n64 71.676
R1397 B.n130 B.n63 71.676
R1398 B.n126 B.n62 71.676
R1399 B.n122 B.n61 71.676
R1400 B.n118 B.n60 71.676
R1401 B.n114 B.n59 71.676
R1402 B.n110 B.n58 71.676
R1403 B.n106 B.n57 71.676
R1404 B.n102 B.n56 71.676
R1405 B.n98 B.n55 71.676
R1406 B.n335 B.n334 71.676
R1407 B.n337 B.n331 71.676
R1408 B.n344 B.n343 71.676
R1409 B.n345 B.n329 71.676
R1410 B.n352 B.n351 71.676
R1411 B.n353 B.n327 71.676
R1412 B.n360 B.n359 71.676
R1413 B.n361 B.n325 71.676
R1414 B.n368 B.n367 71.676
R1415 B.n369 B.n323 71.676
R1416 B.n376 B.n375 71.676
R1417 B.n377 B.n321 71.676
R1418 B.n384 B.n383 71.676
R1419 B.n385 B.n319 71.676
R1420 B.n392 B.n391 71.676
R1421 B.n393 B.n315 71.676
R1422 B.n401 B.n400 71.676
R1423 B.n402 B.n313 71.676
R1424 B.n409 B.n408 71.676
R1425 B.n410 B.n309 71.676
R1426 B.n418 B.n417 71.676
R1427 B.n419 B.n307 71.676
R1428 B.n426 B.n425 71.676
R1429 B.n427 B.n305 71.676
R1430 B.n434 B.n433 71.676
R1431 B.n435 B.n303 71.676
R1432 B.n442 B.n441 71.676
R1433 B.n443 B.n301 71.676
R1434 B.n450 B.n449 71.676
R1435 B.n451 B.n299 71.676
R1436 B.n458 B.n457 71.676
R1437 B.n459 B.n297 71.676
R1438 B.n466 B.n465 71.676
R1439 B.n467 B.n295 71.676
R1440 B.n474 B.n473 71.676
R1441 B.n475 B.n293 71.676
R1442 B.n414 B.n311 59.5399
R1443 B.n396 B.n317 59.5399
R1444 B.n96 B.n95 59.5399
R1445 B.n177 B.n93 59.5399
R1446 B.n481 B.n288 54.0663
R1447 B.n487 B.n288 54.0663
R1448 B.n487 B.n284 54.0663
R1449 B.n494 B.n284 54.0663
R1450 B.n494 B.n493 54.0663
R1451 B.n500 B.n277 54.0663
R1452 B.n506 B.n277 54.0663
R1453 B.n506 B.n273 54.0663
R1454 B.n512 B.n273 54.0663
R1455 B.n512 B.n269 54.0663
R1456 B.n518 B.n269 54.0663
R1457 B.n524 B.n265 54.0663
R1458 B.n524 B.n261 54.0663
R1459 B.n530 B.n261 54.0663
R1460 B.n536 B.n257 54.0663
R1461 B.n536 B.n253 54.0663
R1462 B.n542 B.n253 54.0663
R1463 B.n548 B.n249 54.0663
R1464 B.n548 B.n245 54.0663
R1465 B.n555 B.n245 54.0663
R1466 B.n561 B.n241 54.0663
R1467 B.n561 B.n4 54.0663
R1468 B.n660 B.n4 54.0663
R1469 B.n660 B.n659 54.0663
R1470 B.n659 B.n658 54.0663
R1471 B.n658 B.n8 54.0663
R1472 B.n652 B.n651 54.0663
R1473 B.n651 B.n650 54.0663
R1474 B.n650 B.n15 54.0663
R1475 B.n644 B.n643 54.0663
R1476 B.n643 B.n642 54.0663
R1477 B.n642 B.n22 54.0663
R1478 B.n636 B.n635 54.0663
R1479 B.n635 B.n634 54.0663
R1480 B.n634 B.n29 54.0663
R1481 B.n628 B.n627 54.0663
R1482 B.n627 B.n626 54.0663
R1483 B.n626 B.n36 54.0663
R1484 B.n620 B.n36 54.0663
R1485 B.n620 B.n619 54.0663
R1486 B.n619 B.n618 54.0663
R1487 B.n612 B.n46 54.0663
R1488 B.n612 B.n611 54.0663
R1489 B.n611 B.n610 54.0663
R1490 B.n610 B.n50 54.0663
R1491 B.n604 B.n50 54.0663
R1492 B.n500 B.t8 43.7302
R1493 B.n618 B.t15 43.7302
R1494 B.t2 B.n265 32.599
R1495 B.t4 B.n257 32.599
R1496 B.t0 B.n249 32.599
R1497 B.t6 B.n241 32.599
R1498 B.t5 B.n8 32.599
R1499 B.t1 B.n15 32.599
R1500 B.t21 B.n22 32.599
R1501 B.t3 B.n29 32.599
R1502 B.n606 B.n52 31.3761
R1503 B.n601 B.n600 31.3761
R1504 B.n479 B.n478 31.3761
R1505 B.n483 B.n290 31.3761
R1506 B.n311 B.n310 26.3763
R1507 B.n317 B.n316 26.3763
R1508 B.n95 B.n94 26.3763
R1509 B.n93 B.n92 26.3763
R1510 B.n518 B.t2 21.4678
R1511 B.n530 B.t4 21.4678
R1512 B.n542 B.t0 21.4678
R1513 B.n555 B.t6 21.4678
R1514 B.n652 B.t5 21.4678
R1515 B.n644 B.t1 21.4678
R1516 B.n636 B.t21 21.4678
R1517 B.n628 B.t3 21.4678
R1518 B B.n662 18.0485
R1519 B.n97 B.n52 10.6151
R1520 B.n100 B.n97 10.6151
R1521 B.n101 B.n100 10.6151
R1522 B.n104 B.n101 10.6151
R1523 B.n105 B.n104 10.6151
R1524 B.n108 B.n105 10.6151
R1525 B.n109 B.n108 10.6151
R1526 B.n112 B.n109 10.6151
R1527 B.n113 B.n112 10.6151
R1528 B.n116 B.n113 10.6151
R1529 B.n117 B.n116 10.6151
R1530 B.n120 B.n117 10.6151
R1531 B.n121 B.n120 10.6151
R1532 B.n124 B.n121 10.6151
R1533 B.n125 B.n124 10.6151
R1534 B.n128 B.n125 10.6151
R1535 B.n129 B.n128 10.6151
R1536 B.n132 B.n129 10.6151
R1537 B.n133 B.n132 10.6151
R1538 B.n136 B.n133 10.6151
R1539 B.n137 B.n136 10.6151
R1540 B.n140 B.n137 10.6151
R1541 B.n141 B.n140 10.6151
R1542 B.n144 B.n141 10.6151
R1543 B.n145 B.n144 10.6151
R1544 B.n148 B.n145 10.6151
R1545 B.n149 B.n148 10.6151
R1546 B.n152 B.n149 10.6151
R1547 B.n153 B.n152 10.6151
R1548 B.n156 B.n153 10.6151
R1549 B.n157 B.n156 10.6151
R1550 B.n161 B.n160 10.6151
R1551 B.n164 B.n161 10.6151
R1552 B.n165 B.n164 10.6151
R1553 B.n168 B.n165 10.6151
R1554 B.n169 B.n168 10.6151
R1555 B.n172 B.n169 10.6151
R1556 B.n173 B.n172 10.6151
R1557 B.n176 B.n173 10.6151
R1558 B.n181 B.n178 10.6151
R1559 B.n182 B.n181 10.6151
R1560 B.n185 B.n182 10.6151
R1561 B.n186 B.n185 10.6151
R1562 B.n189 B.n186 10.6151
R1563 B.n190 B.n189 10.6151
R1564 B.n193 B.n190 10.6151
R1565 B.n194 B.n193 10.6151
R1566 B.n197 B.n194 10.6151
R1567 B.n198 B.n197 10.6151
R1568 B.n201 B.n198 10.6151
R1569 B.n202 B.n201 10.6151
R1570 B.n205 B.n202 10.6151
R1571 B.n206 B.n205 10.6151
R1572 B.n209 B.n206 10.6151
R1573 B.n210 B.n209 10.6151
R1574 B.n213 B.n210 10.6151
R1575 B.n214 B.n213 10.6151
R1576 B.n217 B.n214 10.6151
R1577 B.n218 B.n217 10.6151
R1578 B.n221 B.n218 10.6151
R1579 B.n222 B.n221 10.6151
R1580 B.n225 B.n222 10.6151
R1581 B.n226 B.n225 10.6151
R1582 B.n229 B.n226 10.6151
R1583 B.n230 B.n229 10.6151
R1584 B.n233 B.n230 10.6151
R1585 B.n234 B.n233 10.6151
R1586 B.n237 B.n234 10.6151
R1587 B.n238 B.n237 10.6151
R1588 B.n601 B.n238 10.6151
R1589 B.n479 B.n286 10.6151
R1590 B.n489 B.n286 10.6151
R1591 B.n490 B.n489 10.6151
R1592 B.n491 B.n490 10.6151
R1593 B.n491 B.n279 10.6151
R1594 B.n502 B.n279 10.6151
R1595 B.n503 B.n502 10.6151
R1596 B.n504 B.n503 10.6151
R1597 B.n504 B.n271 10.6151
R1598 B.n514 B.n271 10.6151
R1599 B.n515 B.n514 10.6151
R1600 B.n516 B.n515 10.6151
R1601 B.n516 B.n263 10.6151
R1602 B.n526 B.n263 10.6151
R1603 B.n527 B.n526 10.6151
R1604 B.n528 B.n527 10.6151
R1605 B.n528 B.n255 10.6151
R1606 B.n538 B.n255 10.6151
R1607 B.n539 B.n538 10.6151
R1608 B.n540 B.n539 10.6151
R1609 B.n540 B.n247 10.6151
R1610 B.n550 B.n247 10.6151
R1611 B.n551 B.n550 10.6151
R1612 B.n553 B.n551 10.6151
R1613 B.n553 B.n552 10.6151
R1614 B.n552 B.n239 10.6151
R1615 B.n564 B.n239 10.6151
R1616 B.n565 B.n564 10.6151
R1617 B.n566 B.n565 10.6151
R1618 B.n567 B.n566 10.6151
R1619 B.n569 B.n567 10.6151
R1620 B.n570 B.n569 10.6151
R1621 B.n571 B.n570 10.6151
R1622 B.n572 B.n571 10.6151
R1623 B.n574 B.n572 10.6151
R1624 B.n575 B.n574 10.6151
R1625 B.n576 B.n575 10.6151
R1626 B.n577 B.n576 10.6151
R1627 B.n579 B.n577 10.6151
R1628 B.n580 B.n579 10.6151
R1629 B.n581 B.n580 10.6151
R1630 B.n582 B.n581 10.6151
R1631 B.n584 B.n582 10.6151
R1632 B.n585 B.n584 10.6151
R1633 B.n586 B.n585 10.6151
R1634 B.n587 B.n586 10.6151
R1635 B.n589 B.n587 10.6151
R1636 B.n590 B.n589 10.6151
R1637 B.n591 B.n590 10.6151
R1638 B.n592 B.n591 10.6151
R1639 B.n594 B.n592 10.6151
R1640 B.n595 B.n594 10.6151
R1641 B.n596 B.n595 10.6151
R1642 B.n597 B.n596 10.6151
R1643 B.n599 B.n597 10.6151
R1644 B.n600 B.n599 10.6151
R1645 B.n333 B.n290 10.6151
R1646 B.n333 B.n332 10.6151
R1647 B.n339 B.n332 10.6151
R1648 B.n340 B.n339 10.6151
R1649 B.n341 B.n340 10.6151
R1650 B.n341 B.n330 10.6151
R1651 B.n347 B.n330 10.6151
R1652 B.n348 B.n347 10.6151
R1653 B.n349 B.n348 10.6151
R1654 B.n349 B.n328 10.6151
R1655 B.n355 B.n328 10.6151
R1656 B.n356 B.n355 10.6151
R1657 B.n357 B.n356 10.6151
R1658 B.n357 B.n326 10.6151
R1659 B.n363 B.n326 10.6151
R1660 B.n364 B.n363 10.6151
R1661 B.n365 B.n364 10.6151
R1662 B.n365 B.n324 10.6151
R1663 B.n371 B.n324 10.6151
R1664 B.n372 B.n371 10.6151
R1665 B.n373 B.n372 10.6151
R1666 B.n373 B.n322 10.6151
R1667 B.n379 B.n322 10.6151
R1668 B.n380 B.n379 10.6151
R1669 B.n381 B.n380 10.6151
R1670 B.n381 B.n320 10.6151
R1671 B.n387 B.n320 10.6151
R1672 B.n388 B.n387 10.6151
R1673 B.n389 B.n388 10.6151
R1674 B.n389 B.n318 10.6151
R1675 B.n395 B.n318 10.6151
R1676 B.n398 B.n397 10.6151
R1677 B.n398 B.n314 10.6151
R1678 B.n404 B.n314 10.6151
R1679 B.n405 B.n404 10.6151
R1680 B.n406 B.n405 10.6151
R1681 B.n406 B.n312 10.6151
R1682 B.n412 B.n312 10.6151
R1683 B.n413 B.n412 10.6151
R1684 B.n415 B.n308 10.6151
R1685 B.n421 B.n308 10.6151
R1686 B.n422 B.n421 10.6151
R1687 B.n423 B.n422 10.6151
R1688 B.n423 B.n306 10.6151
R1689 B.n429 B.n306 10.6151
R1690 B.n430 B.n429 10.6151
R1691 B.n431 B.n430 10.6151
R1692 B.n431 B.n304 10.6151
R1693 B.n437 B.n304 10.6151
R1694 B.n438 B.n437 10.6151
R1695 B.n439 B.n438 10.6151
R1696 B.n439 B.n302 10.6151
R1697 B.n445 B.n302 10.6151
R1698 B.n446 B.n445 10.6151
R1699 B.n447 B.n446 10.6151
R1700 B.n447 B.n300 10.6151
R1701 B.n453 B.n300 10.6151
R1702 B.n454 B.n453 10.6151
R1703 B.n455 B.n454 10.6151
R1704 B.n455 B.n298 10.6151
R1705 B.n461 B.n298 10.6151
R1706 B.n462 B.n461 10.6151
R1707 B.n463 B.n462 10.6151
R1708 B.n463 B.n296 10.6151
R1709 B.n469 B.n296 10.6151
R1710 B.n470 B.n469 10.6151
R1711 B.n471 B.n470 10.6151
R1712 B.n471 B.n294 10.6151
R1713 B.n477 B.n294 10.6151
R1714 B.n478 B.n477 10.6151
R1715 B.n484 B.n483 10.6151
R1716 B.n485 B.n484 10.6151
R1717 B.n485 B.n282 10.6151
R1718 B.n496 B.n282 10.6151
R1719 B.n497 B.n496 10.6151
R1720 B.n498 B.n497 10.6151
R1721 B.n498 B.n275 10.6151
R1722 B.n508 B.n275 10.6151
R1723 B.n509 B.n508 10.6151
R1724 B.n510 B.n509 10.6151
R1725 B.n510 B.n267 10.6151
R1726 B.n520 B.n267 10.6151
R1727 B.n521 B.n520 10.6151
R1728 B.n522 B.n521 10.6151
R1729 B.n522 B.n259 10.6151
R1730 B.n532 B.n259 10.6151
R1731 B.n533 B.n532 10.6151
R1732 B.n534 B.n533 10.6151
R1733 B.n534 B.n251 10.6151
R1734 B.n544 B.n251 10.6151
R1735 B.n545 B.n544 10.6151
R1736 B.n546 B.n545 10.6151
R1737 B.n546 B.n243 10.6151
R1738 B.n557 B.n243 10.6151
R1739 B.n558 B.n557 10.6151
R1740 B.n559 B.n558 10.6151
R1741 B.n559 B.n0 10.6151
R1742 B.n656 B.n1 10.6151
R1743 B.n656 B.n655 10.6151
R1744 B.n655 B.n654 10.6151
R1745 B.n654 B.n10 10.6151
R1746 B.n648 B.n10 10.6151
R1747 B.n648 B.n647 10.6151
R1748 B.n647 B.n646 10.6151
R1749 B.n646 B.n17 10.6151
R1750 B.n640 B.n17 10.6151
R1751 B.n640 B.n639 10.6151
R1752 B.n639 B.n638 10.6151
R1753 B.n638 B.n24 10.6151
R1754 B.n632 B.n24 10.6151
R1755 B.n632 B.n631 10.6151
R1756 B.n631 B.n630 10.6151
R1757 B.n630 B.n31 10.6151
R1758 B.n624 B.n31 10.6151
R1759 B.n624 B.n623 10.6151
R1760 B.n623 B.n622 10.6151
R1761 B.n622 B.n38 10.6151
R1762 B.n616 B.n38 10.6151
R1763 B.n616 B.n615 10.6151
R1764 B.n615 B.n614 10.6151
R1765 B.n614 B.n44 10.6151
R1766 B.n608 B.n44 10.6151
R1767 B.n608 B.n607 10.6151
R1768 B.n607 B.n606 10.6151
R1769 B.n493 B.t8 10.3366
R1770 B.n46 B.t15 10.3366
R1771 B.n160 B.n96 6.5566
R1772 B.n177 B.n176 6.5566
R1773 B.n397 B.n396 6.5566
R1774 B.n414 B.n413 6.5566
R1775 B.n157 B.n96 4.05904
R1776 B.n178 B.n177 4.05904
R1777 B.n396 B.n395 4.05904
R1778 B.n415 B.n414 4.05904
R1779 B.n662 B.n0 2.81026
R1780 B.n662 B.n1 2.81026
R1781 VN.n4 VN.t3 255.736
R1782 VN.n19 VN.t5 255.736
R1783 VN.n13 VN.t2 238.894
R1784 VN.n28 VN.t0 238.894
R1785 VN.n3 VN.t1 200.287
R1786 VN.n1 VN.t4 200.287
R1787 VN.n18 VN.t7 200.287
R1788 VN.n16 VN.t6 200.287
R1789 VN.n14 VN.n13 161.3
R1790 VN.n29 VN.n28 161.3
R1791 VN.n27 VN.n15 161.3
R1792 VN.n26 VN.n25 161.3
R1793 VN.n24 VN.n23 161.3
R1794 VN.n22 VN.n17 161.3
R1795 VN.n21 VN.n20 161.3
R1796 VN.n12 VN.n0 161.3
R1797 VN.n11 VN.n10 161.3
R1798 VN.n9 VN.n8 161.3
R1799 VN.n7 VN.n2 161.3
R1800 VN.n6 VN.n5 161.3
R1801 VN.n12 VN.n11 54.0429
R1802 VN.n27 VN.n26 54.0429
R1803 VN.n4 VN.n3 45.8978
R1804 VN.n19 VN.n18 45.8978
R1805 VN.n20 VN.n19 43.6106
R1806 VN.n5 VN.n4 43.6106
R1807 VN VN.n29 41.3888
R1808 VN.n7 VN.n6 40.4106
R1809 VN.n8 VN.n7 40.4106
R1810 VN.n22 VN.n21 40.4106
R1811 VN.n23 VN.n22 40.4106
R1812 VN.n11 VN.n1 15.5803
R1813 VN.n26 VN.n16 15.5803
R1814 VN.n6 VN.n3 8.76414
R1815 VN.n8 VN.n1 8.76414
R1816 VN.n21 VN.n18 8.76414
R1817 VN.n23 VN.n16 8.76414
R1818 VN.n13 VN.n12 3.65202
R1819 VN.n28 VN.n27 3.65202
R1820 VN.n29 VN.n15 0.189894
R1821 VN.n25 VN.n15 0.189894
R1822 VN.n25 VN.n24 0.189894
R1823 VN.n24 VN.n17 0.189894
R1824 VN.n20 VN.n17 0.189894
R1825 VN.n5 VN.n2 0.189894
R1826 VN.n9 VN.n2 0.189894
R1827 VN.n10 VN.n9 0.189894
R1828 VN.n10 VN.n0 0.189894
R1829 VN.n14 VN.n0 0.189894
R1830 VN VN.n14 0.0516364
R1831 VDD2.n2 VDD2.n1 64.7476
R1832 VDD2.n2 VDD2.n0 64.7476
R1833 VDD2 VDD2.n5 64.7448
R1834 VDD2.n4 VDD2.n3 64.2169
R1835 VDD2.n4 VDD2.n2 36.3705
R1836 VDD2.n5 VDD2.t0 2.31358
R1837 VDD2.n5 VDD2.t2 2.31358
R1838 VDD2.n3 VDD2.t7 2.31358
R1839 VDD2.n3 VDD2.t1 2.31358
R1840 VDD2.n1 VDD2.t3 2.31358
R1841 VDD2.n1 VDD2.t5 2.31358
R1842 VDD2.n0 VDD2.t4 2.31358
R1843 VDD2.n0 VDD2.t6 2.31358
R1844 VDD2 VDD2.n4 0.644897
C0 VDD1 VN 0.148504f
C1 VTAIL VN 4.84202f
C2 VN VDD2 4.81485f
C3 VN VP 5.1051f
C4 VDD1 VTAIL 7.454589f
C5 VDD1 VDD2 0.990541f
C6 VDD1 VP 5.01796f
C7 VTAIL VDD2 7.49848f
C8 VTAIL VP 4.85613f
C9 VDD2 VP 0.352221f
C10 VDD2 B 3.535875f
C11 VDD1 B 3.807036f
C12 VTAIL B 7.277006f
C13 VN B 9.32815f
C14 VP B 7.688151f
C15 VDD2.t4 B 0.173834f
C16 VDD2.t6 B 0.173834f
C17 VDD2.n0 B 1.51633f
C18 VDD2.t3 B 0.173834f
C19 VDD2.t5 B 0.173834f
C20 VDD2.n1 B 1.51633f
C21 VDD2.n2 B 2.20518f
C22 VDD2.t7 B 0.173834f
C23 VDD2.t1 B 0.173834f
C24 VDD2.n3 B 1.51339f
C25 VDD2.n4 B 2.19043f
C26 VDD2.t0 B 0.173834f
C27 VDD2.t2 B 0.173834f
C28 VDD2.n5 B 1.5163f
C29 VN.n0 B 0.037931f
C30 VN.t4 B 0.900729f
C31 VN.n1 B 0.347488f
C32 VN.n2 B 0.037931f
C33 VN.t1 B 0.900729f
C34 VN.n3 B 0.383537f
C35 VN.t3 B 0.987885f
C36 VN.n4 B 0.402476f
C37 VN.n5 B 0.165159f
C38 VN.n6 B 0.053339f
C39 VN.n7 B 0.030694f
C40 VN.n8 B 0.053339f
C41 VN.n9 B 0.037931f
C42 VN.n10 B 0.037931f
C43 VN.n11 B 0.054178f
C44 VN.n12 B 0.012264f
C45 VN.t2 B 0.960948f
C46 VN.n13 B 0.39819f
C47 VN.n14 B 0.029395f
C48 VN.n15 B 0.037931f
C49 VN.t6 B 0.900729f
C50 VN.n16 B 0.347488f
C51 VN.n17 B 0.037931f
C52 VN.t7 B 0.900729f
C53 VN.n18 B 0.383537f
C54 VN.t5 B 0.987885f
C55 VN.n19 B 0.402476f
C56 VN.n20 B 0.165159f
C57 VN.n21 B 0.053339f
C58 VN.n22 B 0.030694f
C59 VN.n23 B 0.053339f
C60 VN.n24 B 0.037931f
C61 VN.n25 B 0.037931f
C62 VN.n26 B 0.054178f
C63 VN.n27 B 0.012264f
C64 VN.t0 B 0.960948f
C65 VN.n28 B 0.39819f
C66 VN.n29 B 1.52902f
C67 VTAIL.t1 B 0.137024f
C68 VTAIL.t7 B 0.137024f
C69 VTAIL.n0 B 1.13729f
C70 VTAIL.n1 B 0.270849f
C71 VTAIL.n2 B 0.026286f
C72 VTAIL.n3 B 0.020257f
C73 VTAIL.n4 B 0.010885f
C74 VTAIL.n5 B 0.025728f
C75 VTAIL.n6 B 0.011525f
C76 VTAIL.n7 B 0.020257f
C77 VTAIL.n8 B 0.010885f
C78 VTAIL.n9 B 0.025728f
C79 VTAIL.n10 B 0.011525f
C80 VTAIL.n11 B 0.020257f
C81 VTAIL.n12 B 0.010885f
C82 VTAIL.n13 B 0.025728f
C83 VTAIL.n14 B 0.011525f
C84 VTAIL.n15 B 0.119306f
C85 VTAIL.t5 B 0.043084f
C86 VTAIL.n16 B 0.019296f
C87 VTAIL.n17 B 0.018188f
C88 VTAIL.n18 B 0.010885f
C89 VTAIL.n19 B 0.711958f
C90 VTAIL.n20 B 0.020257f
C91 VTAIL.n21 B 0.010885f
C92 VTAIL.n22 B 0.011525f
C93 VTAIL.n23 B 0.025728f
C94 VTAIL.n24 B 0.025728f
C95 VTAIL.n25 B 0.011525f
C96 VTAIL.n26 B 0.010885f
C97 VTAIL.n27 B 0.020257f
C98 VTAIL.n28 B 0.020257f
C99 VTAIL.n29 B 0.010885f
C100 VTAIL.n30 B 0.011525f
C101 VTAIL.n31 B 0.025728f
C102 VTAIL.n32 B 0.025728f
C103 VTAIL.n33 B 0.025728f
C104 VTAIL.n34 B 0.011525f
C105 VTAIL.n35 B 0.010885f
C106 VTAIL.n36 B 0.020257f
C107 VTAIL.n37 B 0.020257f
C108 VTAIL.n38 B 0.010885f
C109 VTAIL.n39 B 0.011205f
C110 VTAIL.n40 B 0.011205f
C111 VTAIL.n41 B 0.025728f
C112 VTAIL.n42 B 0.051831f
C113 VTAIL.n43 B 0.011525f
C114 VTAIL.n44 B 0.010885f
C115 VTAIL.n45 B 0.047929f
C116 VTAIL.n46 B 0.028637f
C117 VTAIL.n47 B 0.125117f
C118 VTAIL.n48 B 0.026286f
C119 VTAIL.n49 B 0.020257f
C120 VTAIL.n50 B 0.010885f
C121 VTAIL.n51 B 0.025728f
C122 VTAIL.n52 B 0.011525f
C123 VTAIL.n53 B 0.020257f
C124 VTAIL.n54 B 0.010885f
C125 VTAIL.n55 B 0.025728f
C126 VTAIL.n56 B 0.011525f
C127 VTAIL.n57 B 0.020257f
C128 VTAIL.n58 B 0.010885f
C129 VTAIL.n59 B 0.025728f
C130 VTAIL.n60 B 0.011525f
C131 VTAIL.n61 B 0.119306f
C132 VTAIL.t13 B 0.043084f
C133 VTAIL.n62 B 0.019296f
C134 VTAIL.n63 B 0.018188f
C135 VTAIL.n64 B 0.010885f
C136 VTAIL.n65 B 0.711958f
C137 VTAIL.n66 B 0.020257f
C138 VTAIL.n67 B 0.010885f
C139 VTAIL.n68 B 0.011525f
C140 VTAIL.n69 B 0.025728f
C141 VTAIL.n70 B 0.025728f
C142 VTAIL.n71 B 0.011525f
C143 VTAIL.n72 B 0.010885f
C144 VTAIL.n73 B 0.020257f
C145 VTAIL.n74 B 0.020257f
C146 VTAIL.n75 B 0.010885f
C147 VTAIL.n76 B 0.011525f
C148 VTAIL.n77 B 0.025728f
C149 VTAIL.n78 B 0.025728f
C150 VTAIL.n79 B 0.025728f
C151 VTAIL.n80 B 0.011525f
C152 VTAIL.n81 B 0.010885f
C153 VTAIL.n82 B 0.020257f
C154 VTAIL.n83 B 0.020257f
C155 VTAIL.n84 B 0.010885f
C156 VTAIL.n85 B 0.011205f
C157 VTAIL.n86 B 0.011205f
C158 VTAIL.n87 B 0.025728f
C159 VTAIL.n88 B 0.051831f
C160 VTAIL.n89 B 0.011525f
C161 VTAIL.n90 B 0.010885f
C162 VTAIL.n91 B 0.047929f
C163 VTAIL.n92 B 0.028637f
C164 VTAIL.n93 B 0.125117f
C165 VTAIL.t9 B 0.137024f
C166 VTAIL.t15 B 0.137024f
C167 VTAIL.n94 B 1.13729f
C168 VTAIL.n95 B 0.343576f
C169 VTAIL.n96 B 0.026286f
C170 VTAIL.n97 B 0.020257f
C171 VTAIL.n98 B 0.010885f
C172 VTAIL.n99 B 0.025728f
C173 VTAIL.n100 B 0.011525f
C174 VTAIL.n101 B 0.020257f
C175 VTAIL.n102 B 0.010885f
C176 VTAIL.n103 B 0.025728f
C177 VTAIL.n104 B 0.011525f
C178 VTAIL.n105 B 0.020257f
C179 VTAIL.n106 B 0.010885f
C180 VTAIL.n107 B 0.025728f
C181 VTAIL.n108 B 0.011525f
C182 VTAIL.n109 B 0.119306f
C183 VTAIL.t10 B 0.043084f
C184 VTAIL.n110 B 0.019296f
C185 VTAIL.n111 B 0.018188f
C186 VTAIL.n112 B 0.010885f
C187 VTAIL.n113 B 0.711958f
C188 VTAIL.n114 B 0.020257f
C189 VTAIL.n115 B 0.010885f
C190 VTAIL.n116 B 0.011525f
C191 VTAIL.n117 B 0.025728f
C192 VTAIL.n118 B 0.025728f
C193 VTAIL.n119 B 0.011525f
C194 VTAIL.n120 B 0.010885f
C195 VTAIL.n121 B 0.020257f
C196 VTAIL.n122 B 0.020257f
C197 VTAIL.n123 B 0.010885f
C198 VTAIL.n124 B 0.011525f
C199 VTAIL.n125 B 0.025728f
C200 VTAIL.n126 B 0.025728f
C201 VTAIL.n127 B 0.025728f
C202 VTAIL.n128 B 0.011525f
C203 VTAIL.n129 B 0.010885f
C204 VTAIL.n130 B 0.020257f
C205 VTAIL.n131 B 0.020257f
C206 VTAIL.n132 B 0.010885f
C207 VTAIL.n133 B 0.011205f
C208 VTAIL.n134 B 0.011205f
C209 VTAIL.n135 B 0.025728f
C210 VTAIL.n136 B 0.051831f
C211 VTAIL.n137 B 0.011525f
C212 VTAIL.n138 B 0.010885f
C213 VTAIL.n139 B 0.047929f
C214 VTAIL.n140 B 0.028637f
C215 VTAIL.n141 B 0.927798f
C216 VTAIL.n142 B 0.026286f
C217 VTAIL.n143 B 0.020257f
C218 VTAIL.n144 B 0.010885f
C219 VTAIL.n145 B 0.025728f
C220 VTAIL.n146 B 0.011525f
C221 VTAIL.n147 B 0.020257f
C222 VTAIL.n148 B 0.010885f
C223 VTAIL.n149 B 0.025728f
C224 VTAIL.n150 B 0.025728f
C225 VTAIL.n151 B 0.011525f
C226 VTAIL.n152 B 0.020257f
C227 VTAIL.n153 B 0.010885f
C228 VTAIL.n154 B 0.025728f
C229 VTAIL.n155 B 0.011525f
C230 VTAIL.n156 B 0.119306f
C231 VTAIL.t2 B 0.043084f
C232 VTAIL.n157 B 0.019296f
C233 VTAIL.n158 B 0.018188f
C234 VTAIL.n159 B 0.010885f
C235 VTAIL.n160 B 0.711958f
C236 VTAIL.n161 B 0.020257f
C237 VTAIL.n162 B 0.010885f
C238 VTAIL.n163 B 0.011525f
C239 VTAIL.n164 B 0.025728f
C240 VTAIL.n165 B 0.025728f
C241 VTAIL.n166 B 0.011525f
C242 VTAIL.n167 B 0.010885f
C243 VTAIL.n168 B 0.020257f
C244 VTAIL.n169 B 0.020257f
C245 VTAIL.n170 B 0.010885f
C246 VTAIL.n171 B 0.011525f
C247 VTAIL.n172 B 0.025728f
C248 VTAIL.n173 B 0.025728f
C249 VTAIL.n174 B 0.011525f
C250 VTAIL.n175 B 0.010885f
C251 VTAIL.n176 B 0.020257f
C252 VTAIL.n177 B 0.020257f
C253 VTAIL.n178 B 0.010885f
C254 VTAIL.n179 B 0.011205f
C255 VTAIL.n180 B 0.011205f
C256 VTAIL.n181 B 0.025728f
C257 VTAIL.n182 B 0.051831f
C258 VTAIL.n183 B 0.011525f
C259 VTAIL.n184 B 0.010885f
C260 VTAIL.n185 B 0.047929f
C261 VTAIL.n186 B 0.028637f
C262 VTAIL.n187 B 0.927798f
C263 VTAIL.t4 B 0.137024f
C264 VTAIL.t0 B 0.137024f
C265 VTAIL.n188 B 1.13729f
C266 VTAIL.n189 B 0.343569f
C267 VTAIL.n190 B 0.026286f
C268 VTAIL.n191 B 0.020257f
C269 VTAIL.n192 B 0.010885f
C270 VTAIL.n193 B 0.025728f
C271 VTAIL.n194 B 0.011525f
C272 VTAIL.n195 B 0.020257f
C273 VTAIL.n196 B 0.010885f
C274 VTAIL.n197 B 0.025728f
C275 VTAIL.n198 B 0.025728f
C276 VTAIL.n199 B 0.011525f
C277 VTAIL.n200 B 0.020257f
C278 VTAIL.n201 B 0.010885f
C279 VTAIL.n202 B 0.025728f
C280 VTAIL.n203 B 0.011525f
C281 VTAIL.n204 B 0.119306f
C282 VTAIL.t6 B 0.043084f
C283 VTAIL.n205 B 0.019296f
C284 VTAIL.n206 B 0.018188f
C285 VTAIL.n207 B 0.010885f
C286 VTAIL.n208 B 0.711958f
C287 VTAIL.n209 B 0.020257f
C288 VTAIL.n210 B 0.010885f
C289 VTAIL.n211 B 0.011525f
C290 VTAIL.n212 B 0.025728f
C291 VTAIL.n213 B 0.025728f
C292 VTAIL.n214 B 0.011525f
C293 VTAIL.n215 B 0.010885f
C294 VTAIL.n216 B 0.020257f
C295 VTAIL.n217 B 0.020257f
C296 VTAIL.n218 B 0.010885f
C297 VTAIL.n219 B 0.011525f
C298 VTAIL.n220 B 0.025728f
C299 VTAIL.n221 B 0.025728f
C300 VTAIL.n222 B 0.011525f
C301 VTAIL.n223 B 0.010885f
C302 VTAIL.n224 B 0.020257f
C303 VTAIL.n225 B 0.020257f
C304 VTAIL.n226 B 0.010885f
C305 VTAIL.n227 B 0.011205f
C306 VTAIL.n228 B 0.011205f
C307 VTAIL.n229 B 0.025728f
C308 VTAIL.n230 B 0.051831f
C309 VTAIL.n231 B 0.011525f
C310 VTAIL.n232 B 0.010885f
C311 VTAIL.n233 B 0.047929f
C312 VTAIL.n234 B 0.028637f
C313 VTAIL.n235 B 0.125117f
C314 VTAIL.n236 B 0.026286f
C315 VTAIL.n237 B 0.020257f
C316 VTAIL.n238 B 0.010885f
C317 VTAIL.n239 B 0.025728f
C318 VTAIL.n240 B 0.011525f
C319 VTAIL.n241 B 0.020257f
C320 VTAIL.n242 B 0.010885f
C321 VTAIL.n243 B 0.025728f
C322 VTAIL.n244 B 0.025728f
C323 VTAIL.n245 B 0.011525f
C324 VTAIL.n246 B 0.020257f
C325 VTAIL.n247 B 0.010885f
C326 VTAIL.n248 B 0.025728f
C327 VTAIL.n249 B 0.011525f
C328 VTAIL.n250 B 0.119306f
C329 VTAIL.t8 B 0.043084f
C330 VTAIL.n251 B 0.019296f
C331 VTAIL.n252 B 0.018188f
C332 VTAIL.n253 B 0.010885f
C333 VTAIL.n254 B 0.711958f
C334 VTAIL.n255 B 0.020257f
C335 VTAIL.n256 B 0.010885f
C336 VTAIL.n257 B 0.011525f
C337 VTAIL.n258 B 0.025728f
C338 VTAIL.n259 B 0.025728f
C339 VTAIL.n260 B 0.011525f
C340 VTAIL.n261 B 0.010885f
C341 VTAIL.n262 B 0.020257f
C342 VTAIL.n263 B 0.020257f
C343 VTAIL.n264 B 0.010885f
C344 VTAIL.n265 B 0.011525f
C345 VTAIL.n266 B 0.025728f
C346 VTAIL.n267 B 0.025728f
C347 VTAIL.n268 B 0.011525f
C348 VTAIL.n269 B 0.010885f
C349 VTAIL.n270 B 0.020257f
C350 VTAIL.n271 B 0.020257f
C351 VTAIL.n272 B 0.010885f
C352 VTAIL.n273 B 0.011205f
C353 VTAIL.n274 B 0.011205f
C354 VTAIL.n275 B 0.025728f
C355 VTAIL.n276 B 0.051831f
C356 VTAIL.n277 B 0.011525f
C357 VTAIL.n278 B 0.010885f
C358 VTAIL.n279 B 0.047929f
C359 VTAIL.n280 B 0.028637f
C360 VTAIL.n281 B 0.125117f
C361 VTAIL.t12 B 0.137024f
C362 VTAIL.t14 B 0.137024f
C363 VTAIL.n282 B 1.13729f
C364 VTAIL.n283 B 0.343569f
C365 VTAIL.n284 B 0.026286f
C366 VTAIL.n285 B 0.020257f
C367 VTAIL.n286 B 0.010885f
C368 VTAIL.n287 B 0.025728f
C369 VTAIL.n288 B 0.011525f
C370 VTAIL.n289 B 0.020257f
C371 VTAIL.n290 B 0.010885f
C372 VTAIL.n291 B 0.025728f
C373 VTAIL.n292 B 0.025728f
C374 VTAIL.n293 B 0.011525f
C375 VTAIL.n294 B 0.020257f
C376 VTAIL.n295 B 0.010885f
C377 VTAIL.n296 B 0.025728f
C378 VTAIL.n297 B 0.011525f
C379 VTAIL.n298 B 0.119306f
C380 VTAIL.t11 B 0.043084f
C381 VTAIL.n299 B 0.019296f
C382 VTAIL.n300 B 0.018188f
C383 VTAIL.n301 B 0.010885f
C384 VTAIL.n302 B 0.711958f
C385 VTAIL.n303 B 0.020257f
C386 VTAIL.n304 B 0.010885f
C387 VTAIL.n305 B 0.011525f
C388 VTAIL.n306 B 0.025728f
C389 VTAIL.n307 B 0.025728f
C390 VTAIL.n308 B 0.011525f
C391 VTAIL.n309 B 0.010885f
C392 VTAIL.n310 B 0.020257f
C393 VTAIL.n311 B 0.020257f
C394 VTAIL.n312 B 0.010885f
C395 VTAIL.n313 B 0.011525f
C396 VTAIL.n314 B 0.025728f
C397 VTAIL.n315 B 0.025728f
C398 VTAIL.n316 B 0.011525f
C399 VTAIL.n317 B 0.010885f
C400 VTAIL.n318 B 0.020257f
C401 VTAIL.n319 B 0.020257f
C402 VTAIL.n320 B 0.010885f
C403 VTAIL.n321 B 0.011205f
C404 VTAIL.n322 B 0.011205f
C405 VTAIL.n323 B 0.025728f
C406 VTAIL.n324 B 0.051831f
C407 VTAIL.n325 B 0.011525f
C408 VTAIL.n326 B 0.010885f
C409 VTAIL.n327 B 0.047929f
C410 VTAIL.n328 B 0.028637f
C411 VTAIL.n329 B 0.927798f
C412 VTAIL.n330 B 0.026286f
C413 VTAIL.n331 B 0.020257f
C414 VTAIL.n332 B 0.010885f
C415 VTAIL.n333 B 0.025728f
C416 VTAIL.n334 B 0.011525f
C417 VTAIL.n335 B 0.020257f
C418 VTAIL.n336 B 0.010885f
C419 VTAIL.n337 B 0.025728f
C420 VTAIL.n338 B 0.011525f
C421 VTAIL.n339 B 0.020257f
C422 VTAIL.n340 B 0.010885f
C423 VTAIL.n341 B 0.025728f
C424 VTAIL.n342 B 0.011525f
C425 VTAIL.n343 B 0.119306f
C426 VTAIL.t3 B 0.043084f
C427 VTAIL.n344 B 0.019296f
C428 VTAIL.n345 B 0.018188f
C429 VTAIL.n346 B 0.010885f
C430 VTAIL.n347 B 0.711958f
C431 VTAIL.n348 B 0.020257f
C432 VTAIL.n349 B 0.010885f
C433 VTAIL.n350 B 0.011525f
C434 VTAIL.n351 B 0.025728f
C435 VTAIL.n352 B 0.025728f
C436 VTAIL.n353 B 0.011525f
C437 VTAIL.n354 B 0.010885f
C438 VTAIL.n355 B 0.020257f
C439 VTAIL.n356 B 0.020257f
C440 VTAIL.n357 B 0.010885f
C441 VTAIL.n358 B 0.011525f
C442 VTAIL.n359 B 0.025728f
C443 VTAIL.n360 B 0.025728f
C444 VTAIL.n361 B 0.025728f
C445 VTAIL.n362 B 0.011525f
C446 VTAIL.n363 B 0.010885f
C447 VTAIL.n364 B 0.020257f
C448 VTAIL.n365 B 0.020257f
C449 VTAIL.n366 B 0.010885f
C450 VTAIL.n367 B 0.011205f
C451 VTAIL.n368 B 0.011205f
C452 VTAIL.n369 B 0.025728f
C453 VTAIL.n370 B 0.051831f
C454 VTAIL.n371 B 0.011525f
C455 VTAIL.n372 B 0.010885f
C456 VTAIL.n373 B 0.047929f
C457 VTAIL.n374 B 0.028637f
C458 VTAIL.n375 B 0.924f
C459 VDD1.t6 B 0.175307f
C460 VDD1.t0 B 0.175307f
C461 VDD1.n0 B 1.5299f
C462 VDD1.t3 B 0.175307f
C463 VDD1.t1 B 0.175307f
C464 VDD1.n1 B 1.52918f
C465 VDD1.t5 B 0.175307f
C466 VDD1.t2 B 0.175307f
C467 VDD1.n2 B 1.52918f
C468 VDD1.n3 B 2.27907f
C469 VDD1.t7 B 0.175307f
C470 VDD1.t4 B 0.175307f
C471 VDD1.n4 B 1.52622f
C472 VDD1.n5 B 2.23981f
C473 VP.n0 B 0.038846f
C474 VP.t0 B 0.922458f
C475 VP.n1 B 0.35587f
C476 VP.n2 B 0.038846f
C477 VP.t6 B 0.922458f
C478 VP.n3 B 0.35587f
C479 VP.n4 B 0.038846f
C480 VP.n5 B 0.038846f
C481 VP.t4 B 0.984129f
C482 VP.t1 B 0.922458f
C483 VP.n6 B 0.35587f
C484 VP.n7 B 0.038846f
C485 VP.t3 B 0.922458f
C486 VP.n8 B 0.392789f
C487 VP.t7 B 1.01172f
C488 VP.n9 B 0.412185f
C489 VP.n10 B 0.169144f
C490 VP.n11 B 0.054626f
C491 VP.n12 B 0.031435f
C492 VP.n13 B 0.054626f
C493 VP.n14 B 0.038846f
C494 VP.n15 B 0.038846f
C495 VP.n16 B 0.055485f
C496 VP.n17 B 0.01256f
C497 VP.n18 B 0.407795f
C498 VP.n19 B 1.54037f
C499 VP.n20 B 1.57432f
C500 VP.t5 B 0.984129f
C501 VP.n21 B 0.407795f
C502 VP.n22 B 0.01256f
C503 VP.n23 B 0.055485f
C504 VP.n24 B 0.038846f
C505 VP.n25 B 0.038846f
C506 VP.n26 B 0.054626f
C507 VP.n27 B 0.031435f
C508 VP.n28 B 0.054626f
C509 VP.n29 B 0.038846f
C510 VP.n30 B 0.038846f
C511 VP.n31 B 0.055485f
C512 VP.n32 B 0.01256f
C513 VP.t2 B 0.984129f
C514 VP.n33 B 0.407795f
C515 VP.n34 B 0.030104f
.ends

