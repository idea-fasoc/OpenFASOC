* NGSPICE file created from diff_pair_sample_0022.ext - technology: sky130A

.subckt diff_pair_sample_0022 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=0 ps=0 w=10.52 l=3.69
X1 VDD1.t5 VP.t0 VTAIL.t11 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=4.1028 ps=21.82 w=10.52 l=3.69
X2 VTAIL.t6 VP.t1 VDD1.t4 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=1.7358 ps=10.85 w=10.52 l=3.69
X3 VTAIL.t9 VP.t2 VDD1.t3 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=1.7358 ps=10.85 w=10.52 l=3.69
X4 VDD2.t5 VN.t0 VTAIL.t2 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=1.7358 ps=10.85 w=10.52 l=3.69
X5 VDD1.t2 VP.t3 VTAIL.t7 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=4.1028 ps=21.82 w=10.52 l=3.69
X6 VDD2.t4 VN.t1 VTAIL.t0 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=4.1028 ps=21.82 w=10.52 l=3.69
X7 VTAIL.t5 VN.t2 VDD2.t3 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=1.7358 ps=10.85 w=10.52 l=3.69
X8 VDD2.t2 VN.t3 VTAIL.t1 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=4.1028 ps=21.82 w=10.52 l=3.69
X9 B.t8 B.t6 B.t7 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=0 ps=0 w=10.52 l=3.69
X10 VDD2.t1 VN.t4 VTAIL.t4 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=1.7358 ps=10.85 w=10.52 l=3.69
X11 B.t5 B.t3 B.t4 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=0 ps=0 w=10.52 l=3.69
X12 B.t2 B.t0 B.t1 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=0 ps=0 w=10.52 l=3.69
X13 VDD1.t1 VP.t4 VTAIL.t10 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=1.7358 ps=10.85 w=10.52 l=3.69
X14 VTAIL.t3 VN.t5 VDD2.t0 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=1.7358 pd=10.85 as=1.7358 ps=10.85 w=10.52 l=3.69
X15 VDD1.t0 VP.t5 VTAIL.t8 w_n4186_n3072# sky130_fd_pr__pfet_01v8 ad=4.1028 pd=21.82 as=1.7358 ps=10.85 w=10.52 l=3.69
R0 B.n413 B.n132 585
R1 B.n412 B.n411 585
R2 B.n410 B.n133 585
R3 B.n409 B.n408 585
R4 B.n407 B.n134 585
R5 B.n406 B.n405 585
R6 B.n404 B.n135 585
R7 B.n403 B.n402 585
R8 B.n401 B.n136 585
R9 B.n400 B.n399 585
R10 B.n398 B.n137 585
R11 B.n397 B.n396 585
R12 B.n395 B.n138 585
R13 B.n394 B.n393 585
R14 B.n392 B.n139 585
R15 B.n391 B.n390 585
R16 B.n389 B.n140 585
R17 B.n388 B.n387 585
R18 B.n386 B.n141 585
R19 B.n385 B.n384 585
R20 B.n383 B.n142 585
R21 B.n382 B.n381 585
R22 B.n380 B.n143 585
R23 B.n379 B.n378 585
R24 B.n377 B.n144 585
R25 B.n376 B.n375 585
R26 B.n374 B.n145 585
R27 B.n373 B.n372 585
R28 B.n371 B.n146 585
R29 B.n370 B.n369 585
R30 B.n368 B.n147 585
R31 B.n367 B.n366 585
R32 B.n365 B.n148 585
R33 B.n364 B.n363 585
R34 B.n362 B.n149 585
R35 B.n361 B.n360 585
R36 B.n359 B.n150 585
R37 B.n358 B.n357 585
R38 B.n353 B.n151 585
R39 B.n352 B.n351 585
R40 B.n350 B.n152 585
R41 B.n349 B.n348 585
R42 B.n347 B.n153 585
R43 B.n346 B.n345 585
R44 B.n344 B.n154 585
R45 B.n343 B.n342 585
R46 B.n341 B.n155 585
R47 B.n339 B.n338 585
R48 B.n337 B.n158 585
R49 B.n336 B.n335 585
R50 B.n334 B.n159 585
R51 B.n333 B.n332 585
R52 B.n331 B.n160 585
R53 B.n330 B.n329 585
R54 B.n328 B.n161 585
R55 B.n327 B.n326 585
R56 B.n325 B.n162 585
R57 B.n324 B.n323 585
R58 B.n322 B.n163 585
R59 B.n321 B.n320 585
R60 B.n319 B.n164 585
R61 B.n318 B.n317 585
R62 B.n316 B.n165 585
R63 B.n315 B.n314 585
R64 B.n313 B.n166 585
R65 B.n312 B.n311 585
R66 B.n310 B.n167 585
R67 B.n309 B.n308 585
R68 B.n307 B.n168 585
R69 B.n306 B.n305 585
R70 B.n304 B.n169 585
R71 B.n303 B.n302 585
R72 B.n301 B.n170 585
R73 B.n300 B.n299 585
R74 B.n298 B.n171 585
R75 B.n297 B.n296 585
R76 B.n295 B.n172 585
R77 B.n294 B.n293 585
R78 B.n292 B.n173 585
R79 B.n291 B.n290 585
R80 B.n289 B.n174 585
R81 B.n288 B.n287 585
R82 B.n286 B.n175 585
R83 B.n285 B.n284 585
R84 B.n415 B.n414 585
R85 B.n416 B.n131 585
R86 B.n418 B.n417 585
R87 B.n419 B.n130 585
R88 B.n421 B.n420 585
R89 B.n422 B.n129 585
R90 B.n424 B.n423 585
R91 B.n425 B.n128 585
R92 B.n427 B.n426 585
R93 B.n428 B.n127 585
R94 B.n430 B.n429 585
R95 B.n431 B.n126 585
R96 B.n433 B.n432 585
R97 B.n434 B.n125 585
R98 B.n436 B.n435 585
R99 B.n437 B.n124 585
R100 B.n439 B.n438 585
R101 B.n440 B.n123 585
R102 B.n442 B.n441 585
R103 B.n443 B.n122 585
R104 B.n445 B.n444 585
R105 B.n446 B.n121 585
R106 B.n448 B.n447 585
R107 B.n449 B.n120 585
R108 B.n451 B.n450 585
R109 B.n452 B.n119 585
R110 B.n454 B.n453 585
R111 B.n455 B.n118 585
R112 B.n457 B.n456 585
R113 B.n458 B.n117 585
R114 B.n460 B.n459 585
R115 B.n461 B.n116 585
R116 B.n463 B.n462 585
R117 B.n464 B.n115 585
R118 B.n466 B.n465 585
R119 B.n467 B.n114 585
R120 B.n469 B.n468 585
R121 B.n470 B.n113 585
R122 B.n472 B.n471 585
R123 B.n473 B.n112 585
R124 B.n475 B.n474 585
R125 B.n476 B.n111 585
R126 B.n478 B.n477 585
R127 B.n479 B.n110 585
R128 B.n481 B.n480 585
R129 B.n482 B.n109 585
R130 B.n484 B.n483 585
R131 B.n485 B.n108 585
R132 B.n487 B.n486 585
R133 B.n488 B.n107 585
R134 B.n490 B.n489 585
R135 B.n491 B.n106 585
R136 B.n493 B.n492 585
R137 B.n494 B.n105 585
R138 B.n496 B.n495 585
R139 B.n497 B.n104 585
R140 B.n499 B.n498 585
R141 B.n500 B.n103 585
R142 B.n502 B.n501 585
R143 B.n503 B.n102 585
R144 B.n505 B.n504 585
R145 B.n506 B.n101 585
R146 B.n508 B.n507 585
R147 B.n509 B.n100 585
R148 B.n511 B.n510 585
R149 B.n512 B.n99 585
R150 B.n514 B.n513 585
R151 B.n515 B.n98 585
R152 B.n517 B.n516 585
R153 B.n518 B.n97 585
R154 B.n520 B.n519 585
R155 B.n521 B.n96 585
R156 B.n523 B.n522 585
R157 B.n524 B.n95 585
R158 B.n526 B.n525 585
R159 B.n527 B.n94 585
R160 B.n529 B.n528 585
R161 B.n530 B.n93 585
R162 B.n532 B.n531 585
R163 B.n533 B.n92 585
R164 B.n535 B.n534 585
R165 B.n536 B.n91 585
R166 B.n538 B.n537 585
R167 B.n539 B.n90 585
R168 B.n541 B.n540 585
R169 B.n542 B.n89 585
R170 B.n544 B.n543 585
R171 B.n545 B.n88 585
R172 B.n547 B.n546 585
R173 B.n548 B.n87 585
R174 B.n550 B.n549 585
R175 B.n551 B.n86 585
R176 B.n553 B.n552 585
R177 B.n554 B.n85 585
R178 B.n556 B.n555 585
R179 B.n557 B.n84 585
R180 B.n559 B.n558 585
R181 B.n560 B.n83 585
R182 B.n562 B.n561 585
R183 B.n563 B.n82 585
R184 B.n565 B.n564 585
R185 B.n566 B.n81 585
R186 B.n568 B.n567 585
R187 B.n569 B.n80 585
R188 B.n571 B.n570 585
R189 B.n572 B.n79 585
R190 B.n574 B.n573 585
R191 B.n575 B.n78 585
R192 B.n577 B.n576 585
R193 B.n578 B.n77 585
R194 B.n580 B.n579 585
R195 B.n581 B.n76 585
R196 B.n709 B.n708 585
R197 B.n707 B.n30 585
R198 B.n706 B.n705 585
R199 B.n704 B.n31 585
R200 B.n703 B.n702 585
R201 B.n701 B.n32 585
R202 B.n700 B.n699 585
R203 B.n698 B.n33 585
R204 B.n697 B.n696 585
R205 B.n695 B.n34 585
R206 B.n694 B.n693 585
R207 B.n692 B.n35 585
R208 B.n691 B.n690 585
R209 B.n689 B.n36 585
R210 B.n688 B.n687 585
R211 B.n686 B.n37 585
R212 B.n685 B.n684 585
R213 B.n683 B.n38 585
R214 B.n682 B.n681 585
R215 B.n680 B.n39 585
R216 B.n679 B.n678 585
R217 B.n677 B.n40 585
R218 B.n676 B.n675 585
R219 B.n674 B.n41 585
R220 B.n673 B.n672 585
R221 B.n671 B.n42 585
R222 B.n670 B.n669 585
R223 B.n668 B.n43 585
R224 B.n667 B.n666 585
R225 B.n665 B.n44 585
R226 B.n664 B.n663 585
R227 B.n662 B.n45 585
R228 B.n661 B.n660 585
R229 B.n659 B.n46 585
R230 B.n658 B.n657 585
R231 B.n656 B.n47 585
R232 B.n655 B.n654 585
R233 B.n653 B.n652 585
R234 B.n651 B.n51 585
R235 B.n650 B.n649 585
R236 B.n648 B.n52 585
R237 B.n647 B.n646 585
R238 B.n645 B.n53 585
R239 B.n644 B.n643 585
R240 B.n642 B.n54 585
R241 B.n641 B.n640 585
R242 B.n639 B.n55 585
R243 B.n637 B.n636 585
R244 B.n635 B.n58 585
R245 B.n634 B.n633 585
R246 B.n632 B.n59 585
R247 B.n631 B.n630 585
R248 B.n629 B.n60 585
R249 B.n628 B.n627 585
R250 B.n626 B.n61 585
R251 B.n625 B.n624 585
R252 B.n623 B.n62 585
R253 B.n622 B.n621 585
R254 B.n620 B.n63 585
R255 B.n619 B.n618 585
R256 B.n617 B.n64 585
R257 B.n616 B.n615 585
R258 B.n614 B.n65 585
R259 B.n613 B.n612 585
R260 B.n611 B.n66 585
R261 B.n610 B.n609 585
R262 B.n608 B.n67 585
R263 B.n607 B.n606 585
R264 B.n605 B.n68 585
R265 B.n604 B.n603 585
R266 B.n602 B.n69 585
R267 B.n601 B.n600 585
R268 B.n599 B.n70 585
R269 B.n598 B.n597 585
R270 B.n596 B.n71 585
R271 B.n595 B.n594 585
R272 B.n593 B.n72 585
R273 B.n592 B.n591 585
R274 B.n590 B.n73 585
R275 B.n589 B.n588 585
R276 B.n587 B.n74 585
R277 B.n586 B.n585 585
R278 B.n584 B.n75 585
R279 B.n583 B.n582 585
R280 B.n710 B.n29 585
R281 B.n712 B.n711 585
R282 B.n713 B.n28 585
R283 B.n715 B.n714 585
R284 B.n716 B.n27 585
R285 B.n718 B.n717 585
R286 B.n719 B.n26 585
R287 B.n721 B.n720 585
R288 B.n722 B.n25 585
R289 B.n724 B.n723 585
R290 B.n725 B.n24 585
R291 B.n727 B.n726 585
R292 B.n728 B.n23 585
R293 B.n730 B.n729 585
R294 B.n731 B.n22 585
R295 B.n733 B.n732 585
R296 B.n734 B.n21 585
R297 B.n736 B.n735 585
R298 B.n737 B.n20 585
R299 B.n739 B.n738 585
R300 B.n740 B.n19 585
R301 B.n742 B.n741 585
R302 B.n743 B.n18 585
R303 B.n745 B.n744 585
R304 B.n746 B.n17 585
R305 B.n748 B.n747 585
R306 B.n749 B.n16 585
R307 B.n751 B.n750 585
R308 B.n752 B.n15 585
R309 B.n754 B.n753 585
R310 B.n755 B.n14 585
R311 B.n757 B.n756 585
R312 B.n758 B.n13 585
R313 B.n760 B.n759 585
R314 B.n761 B.n12 585
R315 B.n763 B.n762 585
R316 B.n764 B.n11 585
R317 B.n766 B.n765 585
R318 B.n767 B.n10 585
R319 B.n769 B.n768 585
R320 B.n770 B.n9 585
R321 B.n772 B.n771 585
R322 B.n773 B.n8 585
R323 B.n775 B.n774 585
R324 B.n776 B.n7 585
R325 B.n778 B.n777 585
R326 B.n779 B.n6 585
R327 B.n781 B.n780 585
R328 B.n782 B.n5 585
R329 B.n784 B.n783 585
R330 B.n785 B.n4 585
R331 B.n787 B.n786 585
R332 B.n788 B.n3 585
R333 B.n790 B.n789 585
R334 B.n791 B.n0 585
R335 B.n2 B.n1 585
R336 B.n204 B.n203 585
R337 B.n205 B.n202 585
R338 B.n207 B.n206 585
R339 B.n208 B.n201 585
R340 B.n210 B.n209 585
R341 B.n211 B.n200 585
R342 B.n213 B.n212 585
R343 B.n214 B.n199 585
R344 B.n216 B.n215 585
R345 B.n217 B.n198 585
R346 B.n219 B.n218 585
R347 B.n220 B.n197 585
R348 B.n222 B.n221 585
R349 B.n223 B.n196 585
R350 B.n225 B.n224 585
R351 B.n226 B.n195 585
R352 B.n228 B.n227 585
R353 B.n229 B.n194 585
R354 B.n231 B.n230 585
R355 B.n232 B.n193 585
R356 B.n234 B.n233 585
R357 B.n235 B.n192 585
R358 B.n237 B.n236 585
R359 B.n238 B.n191 585
R360 B.n240 B.n239 585
R361 B.n241 B.n190 585
R362 B.n243 B.n242 585
R363 B.n244 B.n189 585
R364 B.n246 B.n245 585
R365 B.n247 B.n188 585
R366 B.n249 B.n248 585
R367 B.n250 B.n187 585
R368 B.n252 B.n251 585
R369 B.n253 B.n186 585
R370 B.n255 B.n254 585
R371 B.n256 B.n185 585
R372 B.n258 B.n257 585
R373 B.n259 B.n184 585
R374 B.n261 B.n260 585
R375 B.n262 B.n183 585
R376 B.n264 B.n263 585
R377 B.n265 B.n182 585
R378 B.n267 B.n266 585
R379 B.n268 B.n181 585
R380 B.n270 B.n269 585
R381 B.n271 B.n180 585
R382 B.n273 B.n272 585
R383 B.n274 B.n179 585
R384 B.n276 B.n275 585
R385 B.n277 B.n178 585
R386 B.n279 B.n278 585
R387 B.n280 B.n177 585
R388 B.n282 B.n281 585
R389 B.n283 B.n176 585
R390 B.n284 B.n283 492.5
R391 B.n414 B.n413 492.5
R392 B.n582 B.n581 492.5
R393 B.n708 B.n29 492.5
R394 B.n156 B.t9 277.964
R395 B.n354 B.t6 277.964
R396 B.n56 B.t3 277.964
R397 B.n48 B.t0 277.964
R398 B.n793 B.n792 256.663
R399 B.n792 B.n791 235.042
R400 B.n792 B.n2 235.042
R401 B.n354 B.t7 191.675
R402 B.n56 B.t5 191.675
R403 B.n156 B.t10 191.663
R404 B.n48 B.t2 191.663
R405 B.n284 B.n175 163.367
R406 B.n288 B.n175 163.367
R407 B.n289 B.n288 163.367
R408 B.n290 B.n289 163.367
R409 B.n290 B.n173 163.367
R410 B.n294 B.n173 163.367
R411 B.n295 B.n294 163.367
R412 B.n296 B.n295 163.367
R413 B.n296 B.n171 163.367
R414 B.n300 B.n171 163.367
R415 B.n301 B.n300 163.367
R416 B.n302 B.n301 163.367
R417 B.n302 B.n169 163.367
R418 B.n306 B.n169 163.367
R419 B.n307 B.n306 163.367
R420 B.n308 B.n307 163.367
R421 B.n308 B.n167 163.367
R422 B.n312 B.n167 163.367
R423 B.n313 B.n312 163.367
R424 B.n314 B.n313 163.367
R425 B.n314 B.n165 163.367
R426 B.n318 B.n165 163.367
R427 B.n319 B.n318 163.367
R428 B.n320 B.n319 163.367
R429 B.n320 B.n163 163.367
R430 B.n324 B.n163 163.367
R431 B.n325 B.n324 163.367
R432 B.n326 B.n325 163.367
R433 B.n326 B.n161 163.367
R434 B.n330 B.n161 163.367
R435 B.n331 B.n330 163.367
R436 B.n332 B.n331 163.367
R437 B.n332 B.n159 163.367
R438 B.n336 B.n159 163.367
R439 B.n337 B.n336 163.367
R440 B.n338 B.n337 163.367
R441 B.n338 B.n155 163.367
R442 B.n343 B.n155 163.367
R443 B.n344 B.n343 163.367
R444 B.n345 B.n344 163.367
R445 B.n345 B.n153 163.367
R446 B.n349 B.n153 163.367
R447 B.n350 B.n349 163.367
R448 B.n351 B.n350 163.367
R449 B.n351 B.n151 163.367
R450 B.n358 B.n151 163.367
R451 B.n359 B.n358 163.367
R452 B.n360 B.n359 163.367
R453 B.n360 B.n149 163.367
R454 B.n364 B.n149 163.367
R455 B.n365 B.n364 163.367
R456 B.n366 B.n365 163.367
R457 B.n366 B.n147 163.367
R458 B.n370 B.n147 163.367
R459 B.n371 B.n370 163.367
R460 B.n372 B.n371 163.367
R461 B.n372 B.n145 163.367
R462 B.n376 B.n145 163.367
R463 B.n377 B.n376 163.367
R464 B.n378 B.n377 163.367
R465 B.n378 B.n143 163.367
R466 B.n382 B.n143 163.367
R467 B.n383 B.n382 163.367
R468 B.n384 B.n383 163.367
R469 B.n384 B.n141 163.367
R470 B.n388 B.n141 163.367
R471 B.n389 B.n388 163.367
R472 B.n390 B.n389 163.367
R473 B.n390 B.n139 163.367
R474 B.n394 B.n139 163.367
R475 B.n395 B.n394 163.367
R476 B.n396 B.n395 163.367
R477 B.n396 B.n137 163.367
R478 B.n400 B.n137 163.367
R479 B.n401 B.n400 163.367
R480 B.n402 B.n401 163.367
R481 B.n402 B.n135 163.367
R482 B.n406 B.n135 163.367
R483 B.n407 B.n406 163.367
R484 B.n408 B.n407 163.367
R485 B.n408 B.n133 163.367
R486 B.n412 B.n133 163.367
R487 B.n413 B.n412 163.367
R488 B.n581 B.n580 163.367
R489 B.n580 B.n77 163.367
R490 B.n576 B.n77 163.367
R491 B.n576 B.n575 163.367
R492 B.n575 B.n574 163.367
R493 B.n574 B.n79 163.367
R494 B.n570 B.n79 163.367
R495 B.n570 B.n569 163.367
R496 B.n569 B.n568 163.367
R497 B.n568 B.n81 163.367
R498 B.n564 B.n81 163.367
R499 B.n564 B.n563 163.367
R500 B.n563 B.n562 163.367
R501 B.n562 B.n83 163.367
R502 B.n558 B.n83 163.367
R503 B.n558 B.n557 163.367
R504 B.n557 B.n556 163.367
R505 B.n556 B.n85 163.367
R506 B.n552 B.n85 163.367
R507 B.n552 B.n551 163.367
R508 B.n551 B.n550 163.367
R509 B.n550 B.n87 163.367
R510 B.n546 B.n87 163.367
R511 B.n546 B.n545 163.367
R512 B.n545 B.n544 163.367
R513 B.n544 B.n89 163.367
R514 B.n540 B.n89 163.367
R515 B.n540 B.n539 163.367
R516 B.n539 B.n538 163.367
R517 B.n538 B.n91 163.367
R518 B.n534 B.n91 163.367
R519 B.n534 B.n533 163.367
R520 B.n533 B.n532 163.367
R521 B.n532 B.n93 163.367
R522 B.n528 B.n93 163.367
R523 B.n528 B.n527 163.367
R524 B.n527 B.n526 163.367
R525 B.n526 B.n95 163.367
R526 B.n522 B.n95 163.367
R527 B.n522 B.n521 163.367
R528 B.n521 B.n520 163.367
R529 B.n520 B.n97 163.367
R530 B.n516 B.n97 163.367
R531 B.n516 B.n515 163.367
R532 B.n515 B.n514 163.367
R533 B.n514 B.n99 163.367
R534 B.n510 B.n99 163.367
R535 B.n510 B.n509 163.367
R536 B.n509 B.n508 163.367
R537 B.n508 B.n101 163.367
R538 B.n504 B.n101 163.367
R539 B.n504 B.n503 163.367
R540 B.n503 B.n502 163.367
R541 B.n502 B.n103 163.367
R542 B.n498 B.n103 163.367
R543 B.n498 B.n497 163.367
R544 B.n497 B.n496 163.367
R545 B.n496 B.n105 163.367
R546 B.n492 B.n105 163.367
R547 B.n492 B.n491 163.367
R548 B.n491 B.n490 163.367
R549 B.n490 B.n107 163.367
R550 B.n486 B.n107 163.367
R551 B.n486 B.n485 163.367
R552 B.n485 B.n484 163.367
R553 B.n484 B.n109 163.367
R554 B.n480 B.n109 163.367
R555 B.n480 B.n479 163.367
R556 B.n479 B.n478 163.367
R557 B.n478 B.n111 163.367
R558 B.n474 B.n111 163.367
R559 B.n474 B.n473 163.367
R560 B.n473 B.n472 163.367
R561 B.n472 B.n113 163.367
R562 B.n468 B.n113 163.367
R563 B.n468 B.n467 163.367
R564 B.n467 B.n466 163.367
R565 B.n466 B.n115 163.367
R566 B.n462 B.n115 163.367
R567 B.n462 B.n461 163.367
R568 B.n461 B.n460 163.367
R569 B.n460 B.n117 163.367
R570 B.n456 B.n117 163.367
R571 B.n456 B.n455 163.367
R572 B.n455 B.n454 163.367
R573 B.n454 B.n119 163.367
R574 B.n450 B.n119 163.367
R575 B.n450 B.n449 163.367
R576 B.n449 B.n448 163.367
R577 B.n448 B.n121 163.367
R578 B.n444 B.n121 163.367
R579 B.n444 B.n443 163.367
R580 B.n443 B.n442 163.367
R581 B.n442 B.n123 163.367
R582 B.n438 B.n123 163.367
R583 B.n438 B.n437 163.367
R584 B.n437 B.n436 163.367
R585 B.n436 B.n125 163.367
R586 B.n432 B.n125 163.367
R587 B.n432 B.n431 163.367
R588 B.n431 B.n430 163.367
R589 B.n430 B.n127 163.367
R590 B.n426 B.n127 163.367
R591 B.n426 B.n425 163.367
R592 B.n425 B.n424 163.367
R593 B.n424 B.n129 163.367
R594 B.n420 B.n129 163.367
R595 B.n420 B.n419 163.367
R596 B.n419 B.n418 163.367
R597 B.n418 B.n131 163.367
R598 B.n414 B.n131 163.367
R599 B.n708 B.n707 163.367
R600 B.n707 B.n706 163.367
R601 B.n706 B.n31 163.367
R602 B.n702 B.n31 163.367
R603 B.n702 B.n701 163.367
R604 B.n701 B.n700 163.367
R605 B.n700 B.n33 163.367
R606 B.n696 B.n33 163.367
R607 B.n696 B.n695 163.367
R608 B.n695 B.n694 163.367
R609 B.n694 B.n35 163.367
R610 B.n690 B.n35 163.367
R611 B.n690 B.n689 163.367
R612 B.n689 B.n688 163.367
R613 B.n688 B.n37 163.367
R614 B.n684 B.n37 163.367
R615 B.n684 B.n683 163.367
R616 B.n683 B.n682 163.367
R617 B.n682 B.n39 163.367
R618 B.n678 B.n39 163.367
R619 B.n678 B.n677 163.367
R620 B.n677 B.n676 163.367
R621 B.n676 B.n41 163.367
R622 B.n672 B.n41 163.367
R623 B.n672 B.n671 163.367
R624 B.n671 B.n670 163.367
R625 B.n670 B.n43 163.367
R626 B.n666 B.n43 163.367
R627 B.n666 B.n665 163.367
R628 B.n665 B.n664 163.367
R629 B.n664 B.n45 163.367
R630 B.n660 B.n45 163.367
R631 B.n660 B.n659 163.367
R632 B.n659 B.n658 163.367
R633 B.n658 B.n47 163.367
R634 B.n654 B.n47 163.367
R635 B.n654 B.n653 163.367
R636 B.n653 B.n51 163.367
R637 B.n649 B.n51 163.367
R638 B.n649 B.n648 163.367
R639 B.n648 B.n647 163.367
R640 B.n647 B.n53 163.367
R641 B.n643 B.n53 163.367
R642 B.n643 B.n642 163.367
R643 B.n642 B.n641 163.367
R644 B.n641 B.n55 163.367
R645 B.n636 B.n55 163.367
R646 B.n636 B.n635 163.367
R647 B.n635 B.n634 163.367
R648 B.n634 B.n59 163.367
R649 B.n630 B.n59 163.367
R650 B.n630 B.n629 163.367
R651 B.n629 B.n628 163.367
R652 B.n628 B.n61 163.367
R653 B.n624 B.n61 163.367
R654 B.n624 B.n623 163.367
R655 B.n623 B.n622 163.367
R656 B.n622 B.n63 163.367
R657 B.n618 B.n63 163.367
R658 B.n618 B.n617 163.367
R659 B.n617 B.n616 163.367
R660 B.n616 B.n65 163.367
R661 B.n612 B.n65 163.367
R662 B.n612 B.n611 163.367
R663 B.n611 B.n610 163.367
R664 B.n610 B.n67 163.367
R665 B.n606 B.n67 163.367
R666 B.n606 B.n605 163.367
R667 B.n605 B.n604 163.367
R668 B.n604 B.n69 163.367
R669 B.n600 B.n69 163.367
R670 B.n600 B.n599 163.367
R671 B.n599 B.n598 163.367
R672 B.n598 B.n71 163.367
R673 B.n594 B.n71 163.367
R674 B.n594 B.n593 163.367
R675 B.n593 B.n592 163.367
R676 B.n592 B.n73 163.367
R677 B.n588 B.n73 163.367
R678 B.n588 B.n587 163.367
R679 B.n587 B.n586 163.367
R680 B.n586 B.n75 163.367
R681 B.n582 B.n75 163.367
R682 B.n712 B.n29 163.367
R683 B.n713 B.n712 163.367
R684 B.n714 B.n713 163.367
R685 B.n714 B.n27 163.367
R686 B.n718 B.n27 163.367
R687 B.n719 B.n718 163.367
R688 B.n720 B.n719 163.367
R689 B.n720 B.n25 163.367
R690 B.n724 B.n25 163.367
R691 B.n725 B.n724 163.367
R692 B.n726 B.n725 163.367
R693 B.n726 B.n23 163.367
R694 B.n730 B.n23 163.367
R695 B.n731 B.n730 163.367
R696 B.n732 B.n731 163.367
R697 B.n732 B.n21 163.367
R698 B.n736 B.n21 163.367
R699 B.n737 B.n736 163.367
R700 B.n738 B.n737 163.367
R701 B.n738 B.n19 163.367
R702 B.n742 B.n19 163.367
R703 B.n743 B.n742 163.367
R704 B.n744 B.n743 163.367
R705 B.n744 B.n17 163.367
R706 B.n748 B.n17 163.367
R707 B.n749 B.n748 163.367
R708 B.n750 B.n749 163.367
R709 B.n750 B.n15 163.367
R710 B.n754 B.n15 163.367
R711 B.n755 B.n754 163.367
R712 B.n756 B.n755 163.367
R713 B.n756 B.n13 163.367
R714 B.n760 B.n13 163.367
R715 B.n761 B.n760 163.367
R716 B.n762 B.n761 163.367
R717 B.n762 B.n11 163.367
R718 B.n766 B.n11 163.367
R719 B.n767 B.n766 163.367
R720 B.n768 B.n767 163.367
R721 B.n768 B.n9 163.367
R722 B.n772 B.n9 163.367
R723 B.n773 B.n772 163.367
R724 B.n774 B.n773 163.367
R725 B.n774 B.n7 163.367
R726 B.n778 B.n7 163.367
R727 B.n779 B.n778 163.367
R728 B.n780 B.n779 163.367
R729 B.n780 B.n5 163.367
R730 B.n784 B.n5 163.367
R731 B.n785 B.n784 163.367
R732 B.n786 B.n785 163.367
R733 B.n786 B.n3 163.367
R734 B.n790 B.n3 163.367
R735 B.n791 B.n790 163.367
R736 B.n204 B.n2 163.367
R737 B.n205 B.n204 163.367
R738 B.n206 B.n205 163.367
R739 B.n206 B.n201 163.367
R740 B.n210 B.n201 163.367
R741 B.n211 B.n210 163.367
R742 B.n212 B.n211 163.367
R743 B.n212 B.n199 163.367
R744 B.n216 B.n199 163.367
R745 B.n217 B.n216 163.367
R746 B.n218 B.n217 163.367
R747 B.n218 B.n197 163.367
R748 B.n222 B.n197 163.367
R749 B.n223 B.n222 163.367
R750 B.n224 B.n223 163.367
R751 B.n224 B.n195 163.367
R752 B.n228 B.n195 163.367
R753 B.n229 B.n228 163.367
R754 B.n230 B.n229 163.367
R755 B.n230 B.n193 163.367
R756 B.n234 B.n193 163.367
R757 B.n235 B.n234 163.367
R758 B.n236 B.n235 163.367
R759 B.n236 B.n191 163.367
R760 B.n240 B.n191 163.367
R761 B.n241 B.n240 163.367
R762 B.n242 B.n241 163.367
R763 B.n242 B.n189 163.367
R764 B.n246 B.n189 163.367
R765 B.n247 B.n246 163.367
R766 B.n248 B.n247 163.367
R767 B.n248 B.n187 163.367
R768 B.n252 B.n187 163.367
R769 B.n253 B.n252 163.367
R770 B.n254 B.n253 163.367
R771 B.n254 B.n185 163.367
R772 B.n258 B.n185 163.367
R773 B.n259 B.n258 163.367
R774 B.n260 B.n259 163.367
R775 B.n260 B.n183 163.367
R776 B.n264 B.n183 163.367
R777 B.n265 B.n264 163.367
R778 B.n266 B.n265 163.367
R779 B.n266 B.n181 163.367
R780 B.n270 B.n181 163.367
R781 B.n271 B.n270 163.367
R782 B.n272 B.n271 163.367
R783 B.n272 B.n179 163.367
R784 B.n276 B.n179 163.367
R785 B.n277 B.n276 163.367
R786 B.n278 B.n277 163.367
R787 B.n278 B.n177 163.367
R788 B.n282 B.n177 163.367
R789 B.n283 B.n282 163.367
R790 B.n355 B.t8 113.713
R791 B.n57 B.t4 113.713
R792 B.n157 B.t11 113.701
R793 B.n49 B.t1 113.701
R794 B.n157 B.n156 77.9641
R795 B.n355 B.n354 77.9641
R796 B.n57 B.n56 77.9641
R797 B.n49 B.n48 77.9641
R798 B.n340 B.n157 59.5399
R799 B.n356 B.n355 59.5399
R800 B.n638 B.n57 59.5399
R801 B.n50 B.n49 59.5399
R802 B.n710 B.n709 32.0005
R803 B.n583 B.n76 32.0005
R804 B.n415 B.n132 32.0005
R805 B.n285 B.n176 32.0005
R806 B B.n793 18.0485
R807 B.n711 B.n710 10.6151
R808 B.n711 B.n28 10.6151
R809 B.n715 B.n28 10.6151
R810 B.n716 B.n715 10.6151
R811 B.n717 B.n716 10.6151
R812 B.n717 B.n26 10.6151
R813 B.n721 B.n26 10.6151
R814 B.n722 B.n721 10.6151
R815 B.n723 B.n722 10.6151
R816 B.n723 B.n24 10.6151
R817 B.n727 B.n24 10.6151
R818 B.n728 B.n727 10.6151
R819 B.n729 B.n728 10.6151
R820 B.n729 B.n22 10.6151
R821 B.n733 B.n22 10.6151
R822 B.n734 B.n733 10.6151
R823 B.n735 B.n734 10.6151
R824 B.n735 B.n20 10.6151
R825 B.n739 B.n20 10.6151
R826 B.n740 B.n739 10.6151
R827 B.n741 B.n740 10.6151
R828 B.n741 B.n18 10.6151
R829 B.n745 B.n18 10.6151
R830 B.n746 B.n745 10.6151
R831 B.n747 B.n746 10.6151
R832 B.n747 B.n16 10.6151
R833 B.n751 B.n16 10.6151
R834 B.n752 B.n751 10.6151
R835 B.n753 B.n752 10.6151
R836 B.n753 B.n14 10.6151
R837 B.n757 B.n14 10.6151
R838 B.n758 B.n757 10.6151
R839 B.n759 B.n758 10.6151
R840 B.n759 B.n12 10.6151
R841 B.n763 B.n12 10.6151
R842 B.n764 B.n763 10.6151
R843 B.n765 B.n764 10.6151
R844 B.n765 B.n10 10.6151
R845 B.n769 B.n10 10.6151
R846 B.n770 B.n769 10.6151
R847 B.n771 B.n770 10.6151
R848 B.n771 B.n8 10.6151
R849 B.n775 B.n8 10.6151
R850 B.n776 B.n775 10.6151
R851 B.n777 B.n776 10.6151
R852 B.n777 B.n6 10.6151
R853 B.n781 B.n6 10.6151
R854 B.n782 B.n781 10.6151
R855 B.n783 B.n782 10.6151
R856 B.n783 B.n4 10.6151
R857 B.n787 B.n4 10.6151
R858 B.n788 B.n787 10.6151
R859 B.n789 B.n788 10.6151
R860 B.n789 B.n0 10.6151
R861 B.n709 B.n30 10.6151
R862 B.n705 B.n30 10.6151
R863 B.n705 B.n704 10.6151
R864 B.n704 B.n703 10.6151
R865 B.n703 B.n32 10.6151
R866 B.n699 B.n32 10.6151
R867 B.n699 B.n698 10.6151
R868 B.n698 B.n697 10.6151
R869 B.n697 B.n34 10.6151
R870 B.n693 B.n34 10.6151
R871 B.n693 B.n692 10.6151
R872 B.n692 B.n691 10.6151
R873 B.n691 B.n36 10.6151
R874 B.n687 B.n36 10.6151
R875 B.n687 B.n686 10.6151
R876 B.n686 B.n685 10.6151
R877 B.n685 B.n38 10.6151
R878 B.n681 B.n38 10.6151
R879 B.n681 B.n680 10.6151
R880 B.n680 B.n679 10.6151
R881 B.n679 B.n40 10.6151
R882 B.n675 B.n40 10.6151
R883 B.n675 B.n674 10.6151
R884 B.n674 B.n673 10.6151
R885 B.n673 B.n42 10.6151
R886 B.n669 B.n42 10.6151
R887 B.n669 B.n668 10.6151
R888 B.n668 B.n667 10.6151
R889 B.n667 B.n44 10.6151
R890 B.n663 B.n44 10.6151
R891 B.n663 B.n662 10.6151
R892 B.n662 B.n661 10.6151
R893 B.n661 B.n46 10.6151
R894 B.n657 B.n46 10.6151
R895 B.n657 B.n656 10.6151
R896 B.n656 B.n655 10.6151
R897 B.n652 B.n651 10.6151
R898 B.n651 B.n650 10.6151
R899 B.n650 B.n52 10.6151
R900 B.n646 B.n52 10.6151
R901 B.n646 B.n645 10.6151
R902 B.n645 B.n644 10.6151
R903 B.n644 B.n54 10.6151
R904 B.n640 B.n54 10.6151
R905 B.n640 B.n639 10.6151
R906 B.n637 B.n58 10.6151
R907 B.n633 B.n58 10.6151
R908 B.n633 B.n632 10.6151
R909 B.n632 B.n631 10.6151
R910 B.n631 B.n60 10.6151
R911 B.n627 B.n60 10.6151
R912 B.n627 B.n626 10.6151
R913 B.n626 B.n625 10.6151
R914 B.n625 B.n62 10.6151
R915 B.n621 B.n62 10.6151
R916 B.n621 B.n620 10.6151
R917 B.n620 B.n619 10.6151
R918 B.n619 B.n64 10.6151
R919 B.n615 B.n64 10.6151
R920 B.n615 B.n614 10.6151
R921 B.n614 B.n613 10.6151
R922 B.n613 B.n66 10.6151
R923 B.n609 B.n66 10.6151
R924 B.n609 B.n608 10.6151
R925 B.n608 B.n607 10.6151
R926 B.n607 B.n68 10.6151
R927 B.n603 B.n68 10.6151
R928 B.n603 B.n602 10.6151
R929 B.n602 B.n601 10.6151
R930 B.n601 B.n70 10.6151
R931 B.n597 B.n70 10.6151
R932 B.n597 B.n596 10.6151
R933 B.n596 B.n595 10.6151
R934 B.n595 B.n72 10.6151
R935 B.n591 B.n72 10.6151
R936 B.n591 B.n590 10.6151
R937 B.n590 B.n589 10.6151
R938 B.n589 B.n74 10.6151
R939 B.n585 B.n74 10.6151
R940 B.n585 B.n584 10.6151
R941 B.n584 B.n583 10.6151
R942 B.n579 B.n76 10.6151
R943 B.n579 B.n578 10.6151
R944 B.n578 B.n577 10.6151
R945 B.n577 B.n78 10.6151
R946 B.n573 B.n78 10.6151
R947 B.n573 B.n572 10.6151
R948 B.n572 B.n571 10.6151
R949 B.n571 B.n80 10.6151
R950 B.n567 B.n80 10.6151
R951 B.n567 B.n566 10.6151
R952 B.n566 B.n565 10.6151
R953 B.n565 B.n82 10.6151
R954 B.n561 B.n82 10.6151
R955 B.n561 B.n560 10.6151
R956 B.n560 B.n559 10.6151
R957 B.n559 B.n84 10.6151
R958 B.n555 B.n84 10.6151
R959 B.n555 B.n554 10.6151
R960 B.n554 B.n553 10.6151
R961 B.n553 B.n86 10.6151
R962 B.n549 B.n86 10.6151
R963 B.n549 B.n548 10.6151
R964 B.n548 B.n547 10.6151
R965 B.n547 B.n88 10.6151
R966 B.n543 B.n88 10.6151
R967 B.n543 B.n542 10.6151
R968 B.n542 B.n541 10.6151
R969 B.n541 B.n90 10.6151
R970 B.n537 B.n90 10.6151
R971 B.n537 B.n536 10.6151
R972 B.n536 B.n535 10.6151
R973 B.n535 B.n92 10.6151
R974 B.n531 B.n92 10.6151
R975 B.n531 B.n530 10.6151
R976 B.n530 B.n529 10.6151
R977 B.n529 B.n94 10.6151
R978 B.n525 B.n94 10.6151
R979 B.n525 B.n524 10.6151
R980 B.n524 B.n523 10.6151
R981 B.n523 B.n96 10.6151
R982 B.n519 B.n96 10.6151
R983 B.n519 B.n518 10.6151
R984 B.n518 B.n517 10.6151
R985 B.n517 B.n98 10.6151
R986 B.n513 B.n98 10.6151
R987 B.n513 B.n512 10.6151
R988 B.n512 B.n511 10.6151
R989 B.n511 B.n100 10.6151
R990 B.n507 B.n100 10.6151
R991 B.n507 B.n506 10.6151
R992 B.n506 B.n505 10.6151
R993 B.n505 B.n102 10.6151
R994 B.n501 B.n102 10.6151
R995 B.n501 B.n500 10.6151
R996 B.n500 B.n499 10.6151
R997 B.n499 B.n104 10.6151
R998 B.n495 B.n104 10.6151
R999 B.n495 B.n494 10.6151
R1000 B.n494 B.n493 10.6151
R1001 B.n493 B.n106 10.6151
R1002 B.n489 B.n106 10.6151
R1003 B.n489 B.n488 10.6151
R1004 B.n488 B.n487 10.6151
R1005 B.n487 B.n108 10.6151
R1006 B.n483 B.n108 10.6151
R1007 B.n483 B.n482 10.6151
R1008 B.n482 B.n481 10.6151
R1009 B.n481 B.n110 10.6151
R1010 B.n477 B.n110 10.6151
R1011 B.n477 B.n476 10.6151
R1012 B.n476 B.n475 10.6151
R1013 B.n475 B.n112 10.6151
R1014 B.n471 B.n112 10.6151
R1015 B.n471 B.n470 10.6151
R1016 B.n470 B.n469 10.6151
R1017 B.n469 B.n114 10.6151
R1018 B.n465 B.n114 10.6151
R1019 B.n465 B.n464 10.6151
R1020 B.n464 B.n463 10.6151
R1021 B.n463 B.n116 10.6151
R1022 B.n459 B.n116 10.6151
R1023 B.n459 B.n458 10.6151
R1024 B.n458 B.n457 10.6151
R1025 B.n457 B.n118 10.6151
R1026 B.n453 B.n118 10.6151
R1027 B.n453 B.n452 10.6151
R1028 B.n452 B.n451 10.6151
R1029 B.n451 B.n120 10.6151
R1030 B.n447 B.n120 10.6151
R1031 B.n447 B.n446 10.6151
R1032 B.n446 B.n445 10.6151
R1033 B.n445 B.n122 10.6151
R1034 B.n441 B.n122 10.6151
R1035 B.n441 B.n440 10.6151
R1036 B.n440 B.n439 10.6151
R1037 B.n439 B.n124 10.6151
R1038 B.n435 B.n124 10.6151
R1039 B.n435 B.n434 10.6151
R1040 B.n434 B.n433 10.6151
R1041 B.n433 B.n126 10.6151
R1042 B.n429 B.n126 10.6151
R1043 B.n429 B.n428 10.6151
R1044 B.n428 B.n427 10.6151
R1045 B.n427 B.n128 10.6151
R1046 B.n423 B.n128 10.6151
R1047 B.n423 B.n422 10.6151
R1048 B.n422 B.n421 10.6151
R1049 B.n421 B.n130 10.6151
R1050 B.n417 B.n130 10.6151
R1051 B.n417 B.n416 10.6151
R1052 B.n416 B.n415 10.6151
R1053 B.n203 B.n1 10.6151
R1054 B.n203 B.n202 10.6151
R1055 B.n207 B.n202 10.6151
R1056 B.n208 B.n207 10.6151
R1057 B.n209 B.n208 10.6151
R1058 B.n209 B.n200 10.6151
R1059 B.n213 B.n200 10.6151
R1060 B.n214 B.n213 10.6151
R1061 B.n215 B.n214 10.6151
R1062 B.n215 B.n198 10.6151
R1063 B.n219 B.n198 10.6151
R1064 B.n220 B.n219 10.6151
R1065 B.n221 B.n220 10.6151
R1066 B.n221 B.n196 10.6151
R1067 B.n225 B.n196 10.6151
R1068 B.n226 B.n225 10.6151
R1069 B.n227 B.n226 10.6151
R1070 B.n227 B.n194 10.6151
R1071 B.n231 B.n194 10.6151
R1072 B.n232 B.n231 10.6151
R1073 B.n233 B.n232 10.6151
R1074 B.n233 B.n192 10.6151
R1075 B.n237 B.n192 10.6151
R1076 B.n238 B.n237 10.6151
R1077 B.n239 B.n238 10.6151
R1078 B.n239 B.n190 10.6151
R1079 B.n243 B.n190 10.6151
R1080 B.n244 B.n243 10.6151
R1081 B.n245 B.n244 10.6151
R1082 B.n245 B.n188 10.6151
R1083 B.n249 B.n188 10.6151
R1084 B.n250 B.n249 10.6151
R1085 B.n251 B.n250 10.6151
R1086 B.n251 B.n186 10.6151
R1087 B.n255 B.n186 10.6151
R1088 B.n256 B.n255 10.6151
R1089 B.n257 B.n256 10.6151
R1090 B.n257 B.n184 10.6151
R1091 B.n261 B.n184 10.6151
R1092 B.n262 B.n261 10.6151
R1093 B.n263 B.n262 10.6151
R1094 B.n263 B.n182 10.6151
R1095 B.n267 B.n182 10.6151
R1096 B.n268 B.n267 10.6151
R1097 B.n269 B.n268 10.6151
R1098 B.n269 B.n180 10.6151
R1099 B.n273 B.n180 10.6151
R1100 B.n274 B.n273 10.6151
R1101 B.n275 B.n274 10.6151
R1102 B.n275 B.n178 10.6151
R1103 B.n279 B.n178 10.6151
R1104 B.n280 B.n279 10.6151
R1105 B.n281 B.n280 10.6151
R1106 B.n281 B.n176 10.6151
R1107 B.n286 B.n285 10.6151
R1108 B.n287 B.n286 10.6151
R1109 B.n287 B.n174 10.6151
R1110 B.n291 B.n174 10.6151
R1111 B.n292 B.n291 10.6151
R1112 B.n293 B.n292 10.6151
R1113 B.n293 B.n172 10.6151
R1114 B.n297 B.n172 10.6151
R1115 B.n298 B.n297 10.6151
R1116 B.n299 B.n298 10.6151
R1117 B.n299 B.n170 10.6151
R1118 B.n303 B.n170 10.6151
R1119 B.n304 B.n303 10.6151
R1120 B.n305 B.n304 10.6151
R1121 B.n305 B.n168 10.6151
R1122 B.n309 B.n168 10.6151
R1123 B.n310 B.n309 10.6151
R1124 B.n311 B.n310 10.6151
R1125 B.n311 B.n166 10.6151
R1126 B.n315 B.n166 10.6151
R1127 B.n316 B.n315 10.6151
R1128 B.n317 B.n316 10.6151
R1129 B.n317 B.n164 10.6151
R1130 B.n321 B.n164 10.6151
R1131 B.n322 B.n321 10.6151
R1132 B.n323 B.n322 10.6151
R1133 B.n323 B.n162 10.6151
R1134 B.n327 B.n162 10.6151
R1135 B.n328 B.n327 10.6151
R1136 B.n329 B.n328 10.6151
R1137 B.n329 B.n160 10.6151
R1138 B.n333 B.n160 10.6151
R1139 B.n334 B.n333 10.6151
R1140 B.n335 B.n334 10.6151
R1141 B.n335 B.n158 10.6151
R1142 B.n339 B.n158 10.6151
R1143 B.n342 B.n341 10.6151
R1144 B.n342 B.n154 10.6151
R1145 B.n346 B.n154 10.6151
R1146 B.n347 B.n346 10.6151
R1147 B.n348 B.n347 10.6151
R1148 B.n348 B.n152 10.6151
R1149 B.n352 B.n152 10.6151
R1150 B.n353 B.n352 10.6151
R1151 B.n357 B.n353 10.6151
R1152 B.n361 B.n150 10.6151
R1153 B.n362 B.n361 10.6151
R1154 B.n363 B.n362 10.6151
R1155 B.n363 B.n148 10.6151
R1156 B.n367 B.n148 10.6151
R1157 B.n368 B.n367 10.6151
R1158 B.n369 B.n368 10.6151
R1159 B.n369 B.n146 10.6151
R1160 B.n373 B.n146 10.6151
R1161 B.n374 B.n373 10.6151
R1162 B.n375 B.n374 10.6151
R1163 B.n375 B.n144 10.6151
R1164 B.n379 B.n144 10.6151
R1165 B.n380 B.n379 10.6151
R1166 B.n381 B.n380 10.6151
R1167 B.n381 B.n142 10.6151
R1168 B.n385 B.n142 10.6151
R1169 B.n386 B.n385 10.6151
R1170 B.n387 B.n386 10.6151
R1171 B.n387 B.n140 10.6151
R1172 B.n391 B.n140 10.6151
R1173 B.n392 B.n391 10.6151
R1174 B.n393 B.n392 10.6151
R1175 B.n393 B.n138 10.6151
R1176 B.n397 B.n138 10.6151
R1177 B.n398 B.n397 10.6151
R1178 B.n399 B.n398 10.6151
R1179 B.n399 B.n136 10.6151
R1180 B.n403 B.n136 10.6151
R1181 B.n404 B.n403 10.6151
R1182 B.n405 B.n404 10.6151
R1183 B.n405 B.n134 10.6151
R1184 B.n409 B.n134 10.6151
R1185 B.n410 B.n409 10.6151
R1186 B.n411 B.n410 10.6151
R1187 B.n411 B.n132 10.6151
R1188 B.n655 B.n50 9.36635
R1189 B.n638 B.n637 9.36635
R1190 B.n340 B.n339 9.36635
R1191 B.n356 B.n150 9.36635
R1192 B.n793 B.n0 8.11757
R1193 B.n793 B.n1 8.11757
R1194 B.n652 B.n50 1.24928
R1195 B.n639 B.n638 1.24928
R1196 B.n341 B.n340 1.24928
R1197 B.n357 B.n356 1.24928
R1198 VP.n16 VP.n13 161.3
R1199 VP.n18 VP.n17 161.3
R1200 VP.n19 VP.n12 161.3
R1201 VP.n21 VP.n20 161.3
R1202 VP.n22 VP.n11 161.3
R1203 VP.n24 VP.n23 161.3
R1204 VP.n25 VP.n10 161.3
R1205 VP.n27 VP.n26 161.3
R1206 VP.n56 VP.n55 161.3
R1207 VP.n54 VP.n1 161.3
R1208 VP.n53 VP.n52 161.3
R1209 VP.n51 VP.n2 161.3
R1210 VP.n50 VP.n49 161.3
R1211 VP.n48 VP.n3 161.3
R1212 VP.n47 VP.n46 161.3
R1213 VP.n45 VP.n4 161.3
R1214 VP.n44 VP.n43 161.3
R1215 VP.n42 VP.n5 161.3
R1216 VP.n41 VP.n40 161.3
R1217 VP.n39 VP.n6 161.3
R1218 VP.n38 VP.n37 161.3
R1219 VP.n36 VP.n7 161.3
R1220 VP.n35 VP.n34 161.3
R1221 VP.n33 VP.n8 161.3
R1222 VP.n32 VP.n31 161.3
R1223 VP.n15 VP.t5 101.177
R1224 VP.n30 VP.n29 89.2619
R1225 VP.n57 VP.n0 89.2619
R1226 VP.n28 VP.n9 89.2619
R1227 VP.n43 VP.t1 68.7084
R1228 VP.n30 VP.t4 68.7084
R1229 VP.n0 VP.t0 68.7084
R1230 VP.n14 VP.t2 68.7084
R1231 VP.n9 VP.t3 68.7084
R1232 VP.n29 VP.n28 51.8253
R1233 VP.n15 VP.n14 50.5885
R1234 VP.n37 VP.n36 41.5458
R1235 VP.n49 VP.n2 41.5458
R1236 VP.n20 VP.n11 41.5458
R1237 VP.n37 VP.n6 39.6083
R1238 VP.n49 VP.n48 39.6083
R1239 VP.n20 VP.n19 39.6083
R1240 VP.n31 VP.n8 24.5923
R1241 VP.n35 VP.n8 24.5923
R1242 VP.n36 VP.n35 24.5923
R1243 VP.n41 VP.n6 24.5923
R1244 VP.n42 VP.n41 24.5923
R1245 VP.n43 VP.n42 24.5923
R1246 VP.n43 VP.n4 24.5923
R1247 VP.n47 VP.n4 24.5923
R1248 VP.n48 VP.n47 24.5923
R1249 VP.n53 VP.n2 24.5923
R1250 VP.n54 VP.n53 24.5923
R1251 VP.n55 VP.n54 24.5923
R1252 VP.n24 VP.n11 24.5923
R1253 VP.n25 VP.n24 24.5923
R1254 VP.n26 VP.n25 24.5923
R1255 VP.n14 VP.n13 24.5923
R1256 VP.n18 VP.n13 24.5923
R1257 VP.n19 VP.n18 24.5923
R1258 VP.n16 VP.n15 2.49421
R1259 VP.n31 VP.n30 0.984173
R1260 VP.n55 VP.n0 0.984173
R1261 VP.n26 VP.n9 0.984173
R1262 VP.n28 VP.n27 0.354861
R1263 VP.n32 VP.n29 0.354861
R1264 VP.n57 VP.n56 0.354861
R1265 VP VP.n57 0.267071
R1266 VP.n17 VP.n16 0.189894
R1267 VP.n17 VP.n12 0.189894
R1268 VP.n21 VP.n12 0.189894
R1269 VP.n22 VP.n21 0.189894
R1270 VP.n23 VP.n22 0.189894
R1271 VP.n23 VP.n10 0.189894
R1272 VP.n27 VP.n10 0.189894
R1273 VP.n33 VP.n32 0.189894
R1274 VP.n34 VP.n33 0.189894
R1275 VP.n34 VP.n7 0.189894
R1276 VP.n38 VP.n7 0.189894
R1277 VP.n39 VP.n38 0.189894
R1278 VP.n40 VP.n39 0.189894
R1279 VP.n40 VP.n5 0.189894
R1280 VP.n44 VP.n5 0.189894
R1281 VP.n45 VP.n44 0.189894
R1282 VP.n46 VP.n45 0.189894
R1283 VP.n46 VP.n3 0.189894
R1284 VP.n50 VP.n3 0.189894
R1285 VP.n51 VP.n50 0.189894
R1286 VP.n52 VP.n51 0.189894
R1287 VP.n52 VP.n1 0.189894
R1288 VP.n56 VP.n1 0.189894
R1289 VTAIL.n7 VTAIL.t1 66.7585
R1290 VTAIL.n10 VTAIL.t7 66.7583
R1291 VTAIL.n11 VTAIL.t0 66.7583
R1292 VTAIL.n2 VTAIL.t11 66.7583
R1293 VTAIL.n9 VTAIL.n8 63.6687
R1294 VTAIL.n6 VTAIL.n5 63.6687
R1295 VTAIL.n1 VTAIL.n0 63.6684
R1296 VTAIL.n4 VTAIL.n3 63.6684
R1297 VTAIL.n6 VTAIL.n4 28.3669
R1298 VTAIL.n11 VTAIL.n10 24.9014
R1299 VTAIL.n7 VTAIL.n6 3.46602
R1300 VTAIL.n10 VTAIL.n9 3.46602
R1301 VTAIL.n4 VTAIL.n2 3.46602
R1302 VTAIL.n0 VTAIL.t4 3.09033
R1303 VTAIL.n0 VTAIL.t5 3.09033
R1304 VTAIL.n3 VTAIL.t10 3.09033
R1305 VTAIL.n3 VTAIL.t6 3.09033
R1306 VTAIL.n8 VTAIL.t8 3.09033
R1307 VTAIL.n8 VTAIL.t9 3.09033
R1308 VTAIL.n5 VTAIL.t2 3.09033
R1309 VTAIL.n5 VTAIL.t3 3.09033
R1310 VTAIL VTAIL.n11 2.54145
R1311 VTAIL.n9 VTAIL.n7 2.20309
R1312 VTAIL.n2 VTAIL.n1 2.20309
R1313 VTAIL VTAIL.n1 0.925069
R1314 VDD1 VDD1.t0 86.0946
R1315 VDD1.n1 VDD1.t1 85.9809
R1316 VDD1.n1 VDD1.n0 81.1583
R1317 VDD1.n3 VDD1.n2 80.3473
R1318 VDD1.n3 VDD1.n1 46.363
R1319 VDD1.n2 VDD1.t3 3.09033
R1320 VDD1.n2 VDD1.t2 3.09033
R1321 VDD1.n0 VDD1.t4 3.09033
R1322 VDD1.n0 VDD1.t5 3.09033
R1323 VDD1 VDD1.n3 0.80869
R1324 VN.n38 VN.n37 161.3
R1325 VN.n36 VN.n21 161.3
R1326 VN.n35 VN.n34 161.3
R1327 VN.n33 VN.n22 161.3
R1328 VN.n32 VN.n31 161.3
R1329 VN.n30 VN.n23 161.3
R1330 VN.n29 VN.n28 161.3
R1331 VN.n27 VN.n24 161.3
R1332 VN.n18 VN.n17 161.3
R1333 VN.n16 VN.n1 161.3
R1334 VN.n15 VN.n14 161.3
R1335 VN.n13 VN.n2 161.3
R1336 VN.n12 VN.n11 161.3
R1337 VN.n10 VN.n3 161.3
R1338 VN.n9 VN.n8 161.3
R1339 VN.n7 VN.n4 161.3
R1340 VN.n26 VN.t3 101.177
R1341 VN.n6 VN.t4 101.177
R1342 VN.n19 VN.n0 89.2619
R1343 VN.n39 VN.n20 89.2619
R1344 VN.n5 VN.t2 68.7084
R1345 VN.n0 VN.t1 68.7084
R1346 VN.n25 VN.t5 68.7084
R1347 VN.n20 VN.t0 68.7084
R1348 VN VN.n39 51.9906
R1349 VN.n6 VN.n5 50.5885
R1350 VN.n26 VN.n25 50.5885
R1351 VN.n11 VN.n2 41.5458
R1352 VN.n31 VN.n22 41.5458
R1353 VN.n11 VN.n10 39.6083
R1354 VN.n31 VN.n30 39.6083
R1355 VN.n5 VN.n4 24.5923
R1356 VN.n9 VN.n4 24.5923
R1357 VN.n10 VN.n9 24.5923
R1358 VN.n15 VN.n2 24.5923
R1359 VN.n16 VN.n15 24.5923
R1360 VN.n17 VN.n16 24.5923
R1361 VN.n30 VN.n29 24.5923
R1362 VN.n29 VN.n24 24.5923
R1363 VN.n25 VN.n24 24.5923
R1364 VN.n37 VN.n36 24.5923
R1365 VN.n36 VN.n35 24.5923
R1366 VN.n35 VN.n22 24.5923
R1367 VN.n7 VN.n6 2.49422
R1368 VN.n27 VN.n26 2.49422
R1369 VN.n17 VN.n0 0.984173
R1370 VN.n37 VN.n20 0.984173
R1371 VN.n39 VN.n38 0.354861
R1372 VN.n19 VN.n18 0.354861
R1373 VN VN.n19 0.267071
R1374 VN.n38 VN.n21 0.189894
R1375 VN.n34 VN.n21 0.189894
R1376 VN.n34 VN.n33 0.189894
R1377 VN.n33 VN.n32 0.189894
R1378 VN.n32 VN.n23 0.189894
R1379 VN.n28 VN.n23 0.189894
R1380 VN.n28 VN.n27 0.189894
R1381 VN.n8 VN.n7 0.189894
R1382 VN.n8 VN.n3 0.189894
R1383 VN.n12 VN.n3 0.189894
R1384 VN.n13 VN.n12 0.189894
R1385 VN.n14 VN.n13 0.189894
R1386 VN.n14 VN.n1 0.189894
R1387 VN.n18 VN.n1 0.189894
R1388 VDD2.n1 VDD2.t1 85.9809
R1389 VDD2.n2 VDD2.t5 83.4373
R1390 VDD2.n1 VDD2.n0 81.1583
R1391 VDD2 VDD2.n3 81.1555
R1392 VDD2.n2 VDD2.n1 44.0472
R1393 VDD2.n3 VDD2.t0 3.09033
R1394 VDD2.n3 VDD2.t2 3.09033
R1395 VDD2.n0 VDD2.t3 3.09033
R1396 VDD2.n0 VDD2.t4 3.09033
R1397 VDD2 VDD2.n2 2.65783
C0 VDD2 VN 6.29444f
C1 VDD2 VTAIL 7.69298f
C2 w_n4186_n3072# VDD2 2.57042f
C3 VDD2 VP 0.550582f
C4 VDD2 VDD1 1.83089f
C5 VN B 1.38452f
C6 VTAIL B 3.74742f
C7 w_n4186_n3072# B 10.7666f
C8 B VP 2.29866f
C9 VDD1 B 2.25693f
C10 VTAIL VN 6.78667f
C11 w_n4186_n3072# VN 8.169499f
C12 w_n4186_n3072# VTAIL 2.86403f
C13 VDD2 B 2.35716f
C14 VN VP 7.70971f
C15 VDD1 VN 0.152378f
C16 VTAIL VP 6.80112f
C17 VDD1 VTAIL 7.63371f
C18 w_n4186_n3072# VP 8.71373f
C19 w_n4186_n3072# VDD1 2.45049f
C20 VDD1 VP 6.69002f
C21 VDD2 VSUBS 2.157594f
C22 VDD1 VSUBS 2.72551f
C23 VTAIL VSUBS 1.349888f
C24 VN VSUBS 6.87923f
C25 VP VSUBS 3.723007f
C26 B VSUBS 5.589375f
C27 w_n4186_n3072# VSUBS 0.158683p
C28 VDD2.t1 VSUBS 2.46093f
C29 VDD2.t3 VSUBS 0.242223f
C30 VDD2.t4 VSUBS 0.242223f
C31 VDD2.n0 VSUBS 1.86871f
C32 VDD2.n1 VSUBS 4.3894f
C33 VDD2.t5 VSUBS 2.43564f
C34 VDD2.n2 VSUBS 3.75915f
C35 VDD2.t0 VSUBS 0.242223f
C36 VDD2.t2 VSUBS 0.242223f
C37 VDD2.n3 VSUBS 1.86866f
C38 VN.t1 VSUBS 2.79474f
C39 VN.n0 VSUBS 1.07997f
C40 VN.n1 VSUBS 0.02653f
C41 VN.n2 VSUBS 0.052171f
C42 VN.n3 VSUBS 0.02653f
C43 VN.n4 VSUBS 0.049198f
C44 VN.t2 VSUBS 2.79474f
C45 VN.n5 VSUBS 1.09411f
C46 VN.t4 VSUBS 3.17763f
C47 VN.n6 VSUBS 1.03808f
C48 VN.n7 VSUBS 0.338001f
C49 VN.n8 VSUBS 0.02653f
C50 VN.n9 VSUBS 0.049198f
C51 VN.n10 VSUBS 0.052697f
C52 VN.n11 VSUBS 0.021461f
C53 VN.n12 VSUBS 0.02653f
C54 VN.n13 VSUBS 0.02653f
C55 VN.n14 VSUBS 0.02653f
C56 VN.n15 VSUBS 0.049198f
C57 VN.n16 VSUBS 0.049198f
C58 VN.n17 VSUBS 0.025882f
C59 VN.n18 VSUBS 0.042813f
C60 VN.n19 VSUBS 0.08114f
C61 VN.t0 VSUBS 2.79474f
C62 VN.n20 VSUBS 1.07997f
C63 VN.n21 VSUBS 0.02653f
C64 VN.n22 VSUBS 0.052171f
C65 VN.n23 VSUBS 0.02653f
C66 VN.n24 VSUBS 0.049198f
C67 VN.t3 VSUBS 3.17763f
C68 VN.t5 VSUBS 2.79474f
C69 VN.n25 VSUBS 1.09411f
C70 VN.n26 VSUBS 1.03808f
C71 VN.n27 VSUBS 0.338001f
C72 VN.n28 VSUBS 0.02653f
C73 VN.n29 VSUBS 0.049198f
C74 VN.n30 VSUBS 0.052697f
C75 VN.n31 VSUBS 0.021461f
C76 VN.n32 VSUBS 0.02653f
C77 VN.n33 VSUBS 0.02653f
C78 VN.n34 VSUBS 0.02653f
C79 VN.n35 VSUBS 0.049198f
C80 VN.n36 VSUBS 0.049198f
C81 VN.n37 VSUBS 0.025882f
C82 VN.n38 VSUBS 0.042813f
C83 VN.n39 VSUBS 1.61457f
C84 VDD1.t0 VSUBS 2.46136f
C85 VDD1.t1 VSUBS 2.45995f
C86 VDD1.t4 VSUBS 0.242127f
C87 VDD1.t5 VSUBS 0.242127f
C88 VDD1.n0 VSUBS 1.86797f
C89 VDD1.n1 VSUBS 4.56444f
C90 VDD1.t3 VSUBS 0.242127f
C91 VDD1.t2 VSUBS 0.242127f
C92 VDD1.n2 VSUBS 1.85864f
C93 VDD1.n3 VSUBS 3.75582f
C94 VTAIL.t4 VSUBS 0.255418f
C95 VTAIL.t5 VSUBS 0.255418f
C96 VTAIL.n0 VSUBS 1.81868f
C97 VTAIL.n1 VSUBS 0.957668f
C98 VTAIL.t11 VSUBS 2.41068f
C99 VTAIL.n2 VSUBS 1.31382f
C100 VTAIL.t10 VSUBS 0.255418f
C101 VTAIL.t6 VSUBS 0.255418f
C102 VTAIL.n3 VSUBS 1.81868f
C103 VTAIL.n4 VSUBS 2.99253f
C104 VTAIL.t2 VSUBS 0.255418f
C105 VTAIL.t3 VSUBS 0.255418f
C106 VTAIL.n5 VSUBS 1.81869f
C107 VTAIL.n6 VSUBS 2.99252f
C108 VTAIL.t1 VSUBS 2.41069f
C109 VTAIL.n7 VSUBS 1.31381f
C110 VTAIL.t8 VSUBS 0.255418f
C111 VTAIL.t9 VSUBS 0.255418f
C112 VTAIL.n8 VSUBS 1.81869f
C113 VTAIL.n9 VSUBS 1.20922f
C114 VTAIL.t7 VSUBS 2.41068f
C115 VTAIL.n10 VSUBS 2.75404f
C116 VTAIL.t0 VSUBS 2.41068f
C117 VTAIL.n11 VSUBS 2.6625f
C118 VP.t0 VSUBS 3.10713f
C119 VP.n0 VSUBS 1.20069f
C120 VP.n1 VSUBS 0.029496f
C121 VP.n2 VSUBS 0.058003f
C122 VP.n3 VSUBS 0.029496f
C123 VP.n4 VSUBS 0.054697f
C124 VP.n5 VSUBS 0.029496f
C125 VP.t1 VSUBS 3.10713f
C126 VP.n6 VSUBS 0.058587f
C127 VP.n7 VSUBS 0.029496f
C128 VP.n8 VSUBS 0.054697f
C129 VP.t3 VSUBS 3.10713f
C130 VP.n9 VSUBS 1.20069f
C131 VP.n10 VSUBS 0.029496f
C132 VP.n11 VSUBS 0.058003f
C133 VP.n12 VSUBS 0.029496f
C134 VP.n13 VSUBS 0.054697f
C135 VP.t5 VSUBS 3.5328f
C136 VP.t2 VSUBS 3.10713f
C137 VP.n14 VSUBS 1.2164f
C138 VP.n15 VSUBS 1.15411f
C139 VP.n16 VSUBS 0.375782f
C140 VP.n17 VSUBS 0.029496f
C141 VP.n18 VSUBS 0.054697f
C142 VP.n19 VSUBS 0.058587f
C143 VP.n20 VSUBS 0.02386f
C144 VP.n21 VSUBS 0.029496f
C145 VP.n22 VSUBS 0.029496f
C146 VP.n23 VSUBS 0.029496f
C147 VP.n24 VSUBS 0.054697f
C148 VP.n25 VSUBS 0.054697f
C149 VP.n26 VSUBS 0.028775f
C150 VP.n27 VSUBS 0.047598f
C151 VP.n28 VSUBS 1.78312f
C152 VP.n29 VSUBS 1.80364f
C153 VP.t4 VSUBS 3.10713f
C154 VP.n30 VSUBS 1.20069f
C155 VP.n31 VSUBS 0.028775f
C156 VP.n32 VSUBS 0.047598f
C157 VP.n33 VSUBS 0.029496f
C158 VP.n34 VSUBS 0.029496f
C159 VP.n35 VSUBS 0.054697f
C160 VP.n36 VSUBS 0.058003f
C161 VP.n37 VSUBS 0.02386f
C162 VP.n38 VSUBS 0.029496f
C163 VP.n39 VSUBS 0.029496f
C164 VP.n40 VSUBS 0.029496f
C165 VP.n41 VSUBS 0.054697f
C166 VP.n42 VSUBS 0.054697f
C167 VP.n43 VSUBS 1.1243f
C168 VP.n44 VSUBS 0.029496f
C169 VP.n45 VSUBS 0.029496f
C170 VP.n46 VSUBS 0.029496f
C171 VP.n47 VSUBS 0.054697f
C172 VP.n48 VSUBS 0.058587f
C173 VP.n49 VSUBS 0.02386f
C174 VP.n50 VSUBS 0.029496f
C175 VP.n51 VSUBS 0.029496f
C176 VP.n52 VSUBS 0.029496f
C177 VP.n53 VSUBS 0.054697f
C178 VP.n54 VSUBS 0.054697f
C179 VP.n55 VSUBS 0.028775f
C180 VP.n56 VSUBS 0.047598f
C181 VP.n57 VSUBS 0.090209f
C182 B.n0 VSUBS 0.007848f
C183 B.n1 VSUBS 0.007848f
C184 B.n2 VSUBS 0.011606f
C185 B.n3 VSUBS 0.008894f
C186 B.n4 VSUBS 0.008894f
C187 B.n5 VSUBS 0.008894f
C188 B.n6 VSUBS 0.008894f
C189 B.n7 VSUBS 0.008894f
C190 B.n8 VSUBS 0.008894f
C191 B.n9 VSUBS 0.008894f
C192 B.n10 VSUBS 0.008894f
C193 B.n11 VSUBS 0.008894f
C194 B.n12 VSUBS 0.008894f
C195 B.n13 VSUBS 0.008894f
C196 B.n14 VSUBS 0.008894f
C197 B.n15 VSUBS 0.008894f
C198 B.n16 VSUBS 0.008894f
C199 B.n17 VSUBS 0.008894f
C200 B.n18 VSUBS 0.008894f
C201 B.n19 VSUBS 0.008894f
C202 B.n20 VSUBS 0.008894f
C203 B.n21 VSUBS 0.008894f
C204 B.n22 VSUBS 0.008894f
C205 B.n23 VSUBS 0.008894f
C206 B.n24 VSUBS 0.008894f
C207 B.n25 VSUBS 0.008894f
C208 B.n26 VSUBS 0.008894f
C209 B.n27 VSUBS 0.008894f
C210 B.n28 VSUBS 0.008894f
C211 B.n29 VSUBS 0.020156f
C212 B.n30 VSUBS 0.008894f
C213 B.n31 VSUBS 0.008894f
C214 B.n32 VSUBS 0.008894f
C215 B.n33 VSUBS 0.008894f
C216 B.n34 VSUBS 0.008894f
C217 B.n35 VSUBS 0.008894f
C218 B.n36 VSUBS 0.008894f
C219 B.n37 VSUBS 0.008894f
C220 B.n38 VSUBS 0.008894f
C221 B.n39 VSUBS 0.008894f
C222 B.n40 VSUBS 0.008894f
C223 B.n41 VSUBS 0.008894f
C224 B.n42 VSUBS 0.008894f
C225 B.n43 VSUBS 0.008894f
C226 B.n44 VSUBS 0.008894f
C227 B.n45 VSUBS 0.008894f
C228 B.n46 VSUBS 0.008894f
C229 B.n47 VSUBS 0.008894f
C230 B.t1 VSUBS 0.429014f
C231 B.t2 VSUBS 0.463245f
C232 B.t0 VSUBS 2.31209f
C233 B.n48 VSUBS 0.263858f
C234 B.n49 VSUBS 0.096838f
C235 B.n50 VSUBS 0.020607f
C236 B.n51 VSUBS 0.008894f
C237 B.n52 VSUBS 0.008894f
C238 B.n53 VSUBS 0.008894f
C239 B.n54 VSUBS 0.008894f
C240 B.n55 VSUBS 0.008894f
C241 B.t4 VSUBS 0.429008f
C242 B.t5 VSUBS 0.46324f
C243 B.t3 VSUBS 2.31209f
C244 B.n56 VSUBS 0.263863f
C245 B.n57 VSUBS 0.096844f
C246 B.n58 VSUBS 0.008894f
C247 B.n59 VSUBS 0.008894f
C248 B.n60 VSUBS 0.008894f
C249 B.n61 VSUBS 0.008894f
C250 B.n62 VSUBS 0.008894f
C251 B.n63 VSUBS 0.008894f
C252 B.n64 VSUBS 0.008894f
C253 B.n65 VSUBS 0.008894f
C254 B.n66 VSUBS 0.008894f
C255 B.n67 VSUBS 0.008894f
C256 B.n68 VSUBS 0.008894f
C257 B.n69 VSUBS 0.008894f
C258 B.n70 VSUBS 0.008894f
C259 B.n71 VSUBS 0.008894f
C260 B.n72 VSUBS 0.008894f
C261 B.n73 VSUBS 0.008894f
C262 B.n74 VSUBS 0.008894f
C263 B.n75 VSUBS 0.008894f
C264 B.n76 VSUBS 0.020156f
C265 B.n77 VSUBS 0.008894f
C266 B.n78 VSUBS 0.008894f
C267 B.n79 VSUBS 0.008894f
C268 B.n80 VSUBS 0.008894f
C269 B.n81 VSUBS 0.008894f
C270 B.n82 VSUBS 0.008894f
C271 B.n83 VSUBS 0.008894f
C272 B.n84 VSUBS 0.008894f
C273 B.n85 VSUBS 0.008894f
C274 B.n86 VSUBS 0.008894f
C275 B.n87 VSUBS 0.008894f
C276 B.n88 VSUBS 0.008894f
C277 B.n89 VSUBS 0.008894f
C278 B.n90 VSUBS 0.008894f
C279 B.n91 VSUBS 0.008894f
C280 B.n92 VSUBS 0.008894f
C281 B.n93 VSUBS 0.008894f
C282 B.n94 VSUBS 0.008894f
C283 B.n95 VSUBS 0.008894f
C284 B.n96 VSUBS 0.008894f
C285 B.n97 VSUBS 0.008894f
C286 B.n98 VSUBS 0.008894f
C287 B.n99 VSUBS 0.008894f
C288 B.n100 VSUBS 0.008894f
C289 B.n101 VSUBS 0.008894f
C290 B.n102 VSUBS 0.008894f
C291 B.n103 VSUBS 0.008894f
C292 B.n104 VSUBS 0.008894f
C293 B.n105 VSUBS 0.008894f
C294 B.n106 VSUBS 0.008894f
C295 B.n107 VSUBS 0.008894f
C296 B.n108 VSUBS 0.008894f
C297 B.n109 VSUBS 0.008894f
C298 B.n110 VSUBS 0.008894f
C299 B.n111 VSUBS 0.008894f
C300 B.n112 VSUBS 0.008894f
C301 B.n113 VSUBS 0.008894f
C302 B.n114 VSUBS 0.008894f
C303 B.n115 VSUBS 0.008894f
C304 B.n116 VSUBS 0.008894f
C305 B.n117 VSUBS 0.008894f
C306 B.n118 VSUBS 0.008894f
C307 B.n119 VSUBS 0.008894f
C308 B.n120 VSUBS 0.008894f
C309 B.n121 VSUBS 0.008894f
C310 B.n122 VSUBS 0.008894f
C311 B.n123 VSUBS 0.008894f
C312 B.n124 VSUBS 0.008894f
C313 B.n125 VSUBS 0.008894f
C314 B.n126 VSUBS 0.008894f
C315 B.n127 VSUBS 0.008894f
C316 B.n128 VSUBS 0.008894f
C317 B.n129 VSUBS 0.008894f
C318 B.n130 VSUBS 0.008894f
C319 B.n131 VSUBS 0.008894f
C320 B.n132 VSUBS 0.019842f
C321 B.n133 VSUBS 0.008894f
C322 B.n134 VSUBS 0.008894f
C323 B.n135 VSUBS 0.008894f
C324 B.n136 VSUBS 0.008894f
C325 B.n137 VSUBS 0.008894f
C326 B.n138 VSUBS 0.008894f
C327 B.n139 VSUBS 0.008894f
C328 B.n140 VSUBS 0.008894f
C329 B.n141 VSUBS 0.008894f
C330 B.n142 VSUBS 0.008894f
C331 B.n143 VSUBS 0.008894f
C332 B.n144 VSUBS 0.008894f
C333 B.n145 VSUBS 0.008894f
C334 B.n146 VSUBS 0.008894f
C335 B.n147 VSUBS 0.008894f
C336 B.n148 VSUBS 0.008894f
C337 B.n149 VSUBS 0.008894f
C338 B.n150 VSUBS 0.008371f
C339 B.n151 VSUBS 0.008894f
C340 B.n152 VSUBS 0.008894f
C341 B.n153 VSUBS 0.008894f
C342 B.n154 VSUBS 0.008894f
C343 B.n155 VSUBS 0.008894f
C344 B.t11 VSUBS 0.429014f
C345 B.t10 VSUBS 0.463245f
C346 B.t9 VSUBS 2.31209f
C347 B.n156 VSUBS 0.263858f
C348 B.n157 VSUBS 0.096838f
C349 B.n158 VSUBS 0.008894f
C350 B.n159 VSUBS 0.008894f
C351 B.n160 VSUBS 0.008894f
C352 B.n161 VSUBS 0.008894f
C353 B.n162 VSUBS 0.008894f
C354 B.n163 VSUBS 0.008894f
C355 B.n164 VSUBS 0.008894f
C356 B.n165 VSUBS 0.008894f
C357 B.n166 VSUBS 0.008894f
C358 B.n167 VSUBS 0.008894f
C359 B.n168 VSUBS 0.008894f
C360 B.n169 VSUBS 0.008894f
C361 B.n170 VSUBS 0.008894f
C362 B.n171 VSUBS 0.008894f
C363 B.n172 VSUBS 0.008894f
C364 B.n173 VSUBS 0.008894f
C365 B.n174 VSUBS 0.008894f
C366 B.n175 VSUBS 0.008894f
C367 B.n176 VSUBS 0.020156f
C368 B.n177 VSUBS 0.008894f
C369 B.n178 VSUBS 0.008894f
C370 B.n179 VSUBS 0.008894f
C371 B.n180 VSUBS 0.008894f
C372 B.n181 VSUBS 0.008894f
C373 B.n182 VSUBS 0.008894f
C374 B.n183 VSUBS 0.008894f
C375 B.n184 VSUBS 0.008894f
C376 B.n185 VSUBS 0.008894f
C377 B.n186 VSUBS 0.008894f
C378 B.n187 VSUBS 0.008894f
C379 B.n188 VSUBS 0.008894f
C380 B.n189 VSUBS 0.008894f
C381 B.n190 VSUBS 0.008894f
C382 B.n191 VSUBS 0.008894f
C383 B.n192 VSUBS 0.008894f
C384 B.n193 VSUBS 0.008894f
C385 B.n194 VSUBS 0.008894f
C386 B.n195 VSUBS 0.008894f
C387 B.n196 VSUBS 0.008894f
C388 B.n197 VSUBS 0.008894f
C389 B.n198 VSUBS 0.008894f
C390 B.n199 VSUBS 0.008894f
C391 B.n200 VSUBS 0.008894f
C392 B.n201 VSUBS 0.008894f
C393 B.n202 VSUBS 0.008894f
C394 B.n203 VSUBS 0.008894f
C395 B.n204 VSUBS 0.008894f
C396 B.n205 VSUBS 0.008894f
C397 B.n206 VSUBS 0.008894f
C398 B.n207 VSUBS 0.008894f
C399 B.n208 VSUBS 0.008894f
C400 B.n209 VSUBS 0.008894f
C401 B.n210 VSUBS 0.008894f
C402 B.n211 VSUBS 0.008894f
C403 B.n212 VSUBS 0.008894f
C404 B.n213 VSUBS 0.008894f
C405 B.n214 VSUBS 0.008894f
C406 B.n215 VSUBS 0.008894f
C407 B.n216 VSUBS 0.008894f
C408 B.n217 VSUBS 0.008894f
C409 B.n218 VSUBS 0.008894f
C410 B.n219 VSUBS 0.008894f
C411 B.n220 VSUBS 0.008894f
C412 B.n221 VSUBS 0.008894f
C413 B.n222 VSUBS 0.008894f
C414 B.n223 VSUBS 0.008894f
C415 B.n224 VSUBS 0.008894f
C416 B.n225 VSUBS 0.008894f
C417 B.n226 VSUBS 0.008894f
C418 B.n227 VSUBS 0.008894f
C419 B.n228 VSUBS 0.008894f
C420 B.n229 VSUBS 0.008894f
C421 B.n230 VSUBS 0.008894f
C422 B.n231 VSUBS 0.008894f
C423 B.n232 VSUBS 0.008894f
C424 B.n233 VSUBS 0.008894f
C425 B.n234 VSUBS 0.008894f
C426 B.n235 VSUBS 0.008894f
C427 B.n236 VSUBS 0.008894f
C428 B.n237 VSUBS 0.008894f
C429 B.n238 VSUBS 0.008894f
C430 B.n239 VSUBS 0.008894f
C431 B.n240 VSUBS 0.008894f
C432 B.n241 VSUBS 0.008894f
C433 B.n242 VSUBS 0.008894f
C434 B.n243 VSUBS 0.008894f
C435 B.n244 VSUBS 0.008894f
C436 B.n245 VSUBS 0.008894f
C437 B.n246 VSUBS 0.008894f
C438 B.n247 VSUBS 0.008894f
C439 B.n248 VSUBS 0.008894f
C440 B.n249 VSUBS 0.008894f
C441 B.n250 VSUBS 0.008894f
C442 B.n251 VSUBS 0.008894f
C443 B.n252 VSUBS 0.008894f
C444 B.n253 VSUBS 0.008894f
C445 B.n254 VSUBS 0.008894f
C446 B.n255 VSUBS 0.008894f
C447 B.n256 VSUBS 0.008894f
C448 B.n257 VSUBS 0.008894f
C449 B.n258 VSUBS 0.008894f
C450 B.n259 VSUBS 0.008894f
C451 B.n260 VSUBS 0.008894f
C452 B.n261 VSUBS 0.008894f
C453 B.n262 VSUBS 0.008894f
C454 B.n263 VSUBS 0.008894f
C455 B.n264 VSUBS 0.008894f
C456 B.n265 VSUBS 0.008894f
C457 B.n266 VSUBS 0.008894f
C458 B.n267 VSUBS 0.008894f
C459 B.n268 VSUBS 0.008894f
C460 B.n269 VSUBS 0.008894f
C461 B.n270 VSUBS 0.008894f
C462 B.n271 VSUBS 0.008894f
C463 B.n272 VSUBS 0.008894f
C464 B.n273 VSUBS 0.008894f
C465 B.n274 VSUBS 0.008894f
C466 B.n275 VSUBS 0.008894f
C467 B.n276 VSUBS 0.008894f
C468 B.n277 VSUBS 0.008894f
C469 B.n278 VSUBS 0.008894f
C470 B.n279 VSUBS 0.008894f
C471 B.n280 VSUBS 0.008894f
C472 B.n281 VSUBS 0.008894f
C473 B.n282 VSUBS 0.008894f
C474 B.n283 VSUBS 0.020156f
C475 B.n284 VSUBS 0.020914f
C476 B.n285 VSUBS 0.020914f
C477 B.n286 VSUBS 0.008894f
C478 B.n287 VSUBS 0.008894f
C479 B.n288 VSUBS 0.008894f
C480 B.n289 VSUBS 0.008894f
C481 B.n290 VSUBS 0.008894f
C482 B.n291 VSUBS 0.008894f
C483 B.n292 VSUBS 0.008894f
C484 B.n293 VSUBS 0.008894f
C485 B.n294 VSUBS 0.008894f
C486 B.n295 VSUBS 0.008894f
C487 B.n296 VSUBS 0.008894f
C488 B.n297 VSUBS 0.008894f
C489 B.n298 VSUBS 0.008894f
C490 B.n299 VSUBS 0.008894f
C491 B.n300 VSUBS 0.008894f
C492 B.n301 VSUBS 0.008894f
C493 B.n302 VSUBS 0.008894f
C494 B.n303 VSUBS 0.008894f
C495 B.n304 VSUBS 0.008894f
C496 B.n305 VSUBS 0.008894f
C497 B.n306 VSUBS 0.008894f
C498 B.n307 VSUBS 0.008894f
C499 B.n308 VSUBS 0.008894f
C500 B.n309 VSUBS 0.008894f
C501 B.n310 VSUBS 0.008894f
C502 B.n311 VSUBS 0.008894f
C503 B.n312 VSUBS 0.008894f
C504 B.n313 VSUBS 0.008894f
C505 B.n314 VSUBS 0.008894f
C506 B.n315 VSUBS 0.008894f
C507 B.n316 VSUBS 0.008894f
C508 B.n317 VSUBS 0.008894f
C509 B.n318 VSUBS 0.008894f
C510 B.n319 VSUBS 0.008894f
C511 B.n320 VSUBS 0.008894f
C512 B.n321 VSUBS 0.008894f
C513 B.n322 VSUBS 0.008894f
C514 B.n323 VSUBS 0.008894f
C515 B.n324 VSUBS 0.008894f
C516 B.n325 VSUBS 0.008894f
C517 B.n326 VSUBS 0.008894f
C518 B.n327 VSUBS 0.008894f
C519 B.n328 VSUBS 0.008894f
C520 B.n329 VSUBS 0.008894f
C521 B.n330 VSUBS 0.008894f
C522 B.n331 VSUBS 0.008894f
C523 B.n332 VSUBS 0.008894f
C524 B.n333 VSUBS 0.008894f
C525 B.n334 VSUBS 0.008894f
C526 B.n335 VSUBS 0.008894f
C527 B.n336 VSUBS 0.008894f
C528 B.n337 VSUBS 0.008894f
C529 B.n338 VSUBS 0.008894f
C530 B.n339 VSUBS 0.008371f
C531 B.n340 VSUBS 0.020607f
C532 B.n341 VSUBS 0.00497f
C533 B.n342 VSUBS 0.008894f
C534 B.n343 VSUBS 0.008894f
C535 B.n344 VSUBS 0.008894f
C536 B.n345 VSUBS 0.008894f
C537 B.n346 VSUBS 0.008894f
C538 B.n347 VSUBS 0.008894f
C539 B.n348 VSUBS 0.008894f
C540 B.n349 VSUBS 0.008894f
C541 B.n350 VSUBS 0.008894f
C542 B.n351 VSUBS 0.008894f
C543 B.n352 VSUBS 0.008894f
C544 B.n353 VSUBS 0.008894f
C545 B.t8 VSUBS 0.429008f
C546 B.t7 VSUBS 0.46324f
C547 B.t6 VSUBS 2.31209f
C548 B.n354 VSUBS 0.263863f
C549 B.n355 VSUBS 0.096844f
C550 B.n356 VSUBS 0.020607f
C551 B.n357 VSUBS 0.00497f
C552 B.n358 VSUBS 0.008894f
C553 B.n359 VSUBS 0.008894f
C554 B.n360 VSUBS 0.008894f
C555 B.n361 VSUBS 0.008894f
C556 B.n362 VSUBS 0.008894f
C557 B.n363 VSUBS 0.008894f
C558 B.n364 VSUBS 0.008894f
C559 B.n365 VSUBS 0.008894f
C560 B.n366 VSUBS 0.008894f
C561 B.n367 VSUBS 0.008894f
C562 B.n368 VSUBS 0.008894f
C563 B.n369 VSUBS 0.008894f
C564 B.n370 VSUBS 0.008894f
C565 B.n371 VSUBS 0.008894f
C566 B.n372 VSUBS 0.008894f
C567 B.n373 VSUBS 0.008894f
C568 B.n374 VSUBS 0.008894f
C569 B.n375 VSUBS 0.008894f
C570 B.n376 VSUBS 0.008894f
C571 B.n377 VSUBS 0.008894f
C572 B.n378 VSUBS 0.008894f
C573 B.n379 VSUBS 0.008894f
C574 B.n380 VSUBS 0.008894f
C575 B.n381 VSUBS 0.008894f
C576 B.n382 VSUBS 0.008894f
C577 B.n383 VSUBS 0.008894f
C578 B.n384 VSUBS 0.008894f
C579 B.n385 VSUBS 0.008894f
C580 B.n386 VSUBS 0.008894f
C581 B.n387 VSUBS 0.008894f
C582 B.n388 VSUBS 0.008894f
C583 B.n389 VSUBS 0.008894f
C584 B.n390 VSUBS 0.008894f
C585 B.n391 VSUBS 0.008894f
C586 B.n392 VSUBS 0.008894f
C587 B.n393 VSUBS 0.008894f
C588 B.n394 VSUBS 0.008894f
C589 B.n395 VSUBS 0.008894f
C590 B.n396 VSUBS 0.008894f
C591 B.n397 VSUBS 0.008894f
C592 B.n398 VSUBS 0.008894f
C593 B.n399 VSUBS 0.008894f
C594 B.n400 VSUBS 0.008894f
C595 B.n401 VSUBS 0.008894f
C596 B.n402 VSUBS 0.008894f
C597 B.n403 VSUBS 0.008894f
C598 B.n404 VSUBS 0.008894f
C599 B.n405 VSUBS 0.008894f
C600 B.n406 VSUBS 0.008894f
C601 B.n407 VSUBS 0.008894f
C602 B.n408 VSUBS 0.008894f
C603 B.n409 VSUBS 0.008894f
C604 B.n410 VSUBS 0.008894f
C605 B.n411 VSUBS 0.008894f
C606 B.n412 VSUBS 0.008894f
C607 B.n413 VSUBS 0.020914f
C608 B.n414 VSUBS 0.020156f
C609 B.n415 VSUBS 0.021228f
C610 B.n416 VSUBS 0.008894f
C611 B.n417 VSUBS 0.008894f
C612 B.n418 VSUBS 0.008894f
C613 B.n419 VSUBS 0.008894f
C614 B.n420 VSUBS 0.008894f
C615 B.n421 VSUBS 0.008894f
C616 B.n422 VSUBS 0.008894f
C617 B.n423 VSUBS 0.008894f
C618 B.n424 VSUBS 0.008894f
C619 B.n425 VSUBS 0.008894f
C620 B.n426 VSUBS 0.008894f
C621 B.n427 VSUBS 0.008894f
C622 B.n428 VSUBS 0.008894f
C623 B.n429 VSUBS 0.008894f
C624 B.n430 VSUBS 0.008894f
C625 B.n431 VSUBS 0.008894f
C626 B.n432 VSUBS 0.008894f
C627 B.n433 VSUBS 0.008894f
C628 B.n434 VSUBS 0.008894f
C629 B.n435 VSUBS 0.008894f
C630 B.n436 VSUBS 0.008894f
C631 B.n437 VSUBS 0.008894f
C632 B.n438 VSUBS 0.008894f
C633 B.n439 VSUBS 0.008894f
C634 B.n440 VSUBS 0.008894f
C635 B.n441 VSUBS 0.008894f
C636 B.n442 VSUBS 0.008894f
C637 B.n443 VSUBS 0.008894f
C638 B.n444 VSUBS 0.008894f
C639 B.n445 VSUBS 0.008894f
C640 B.n446 VSUBS 0.008894f
C641 B.n447 VSUBS 0.008894f
C642 B.n448 VSUBS 0.008894f
C643 B.n449 VSUBS 0.008894f
C644 B.n450 VSUBS 0.008894f
C645 B.n451 VSUBS 0.008894f
C646 B.n452 VSUBS 0.008894f
C647 B.n453 VSUBS 0.008894f
C648 B.n454 VSUBS 0.008894f
C649 B.n455 VSUBS 0.008894f
C650 B.n456 VSUBS 0.008894f
C651 B.n457 VSUBS 0.008894f
C652 B.n458 VSUBS 0.008894f
C653 B.n459 VSUBS 0.008894f
C654 B.n460 VSUBS 0.008894f
C655 B.n461 VSUBS 0.008894f
C656 B.n462 VSUBS 0.008894f
C657 B.n463 VSUBS 0.008894f
C658 B.n464 VSUBS 0.008894f
C659 B.n465 VSUBS 0.008894f
C660 B.n466 VSUBS 0.008894f
C661 B.n467 VSUBS 0.008894f
C662 B.n468 VSUBS 0.008894f
C663 B.n469 VSUBS 0.008894f
C664 B.n470 VSUBS 0.008894f
C665 B.n471 VSUBS 0.008894f
C666 B.n472 VSUBS 0.008894f
C667 B.n473 VSUBS 0.008894f
C668 B.n474 VSUBS 0.008894f
C669 B.n475 VSUBS 0.008894f
C670 B.n476 VSUBS 0.008894f
C671 B.n477 VSUBS 0.008894f
C672 B.n478 VSUBS 0.008894f
C673 B.n479 VSUBS 0.008894f
C674 B.n480 VSUBS 0.008894f
C675 B.n481 VSUBS 0.008894f
C676 B.n482 VSUBS 0.008894f
C677 B.n483 VSUBS 0.008894f
C678 B.n484 VSUBS 0.008894f
C679 B.n485 VSUBS 0.008894f
C680 B.n486 VSUBS 0.008894f
C681 B.n487 VSUBS 0.008894f
C682 B.n488 VSUBS 0.008894f
C683 B.n489 VSUBS 0.008894f
C684 B.n490 VSUBS 0.008894f
C685 B.n491 VSUBS 0.008894f
C686 B.n492 VSUBS 0.008894f
C687 B.n493 VSUBS 0.008894f
C688 B.n494 VSUBS 0.008894f
C689 B.n495 VSUBS 0.008894f
C690 B.n496 VSUBS 0.008894f
C691 B.n497 VSUBS 0.008894f
C692 B.n498 VSUBS 0.008894f
C693 B.n499 VSUBS 0.008894f
C694 B.n500 VSUBS 0.008894f
C695 B.n501 VSUBS 0.008894f
C696 B.n502 VSUBS 0.008894f
C697 B.n503 VSUBS 0.008894f
C698 B.n504 VSUBS 0.008894f
C699 B.n505 VSUBS 0.008894f
C700 B.n506 VSUBS 0.008894f
C701 B.n507 VSUBS 0.008894f
C702 B.n508 VSUBS 0.008894f
C703 B.n509 VSUBS 0.008894f
C704 B.n510 VSUBS 0.008894f
C705 B.n511 VSUBS 0.008894f
C706 B.n512 VSUBS 0.008894f
C707 B.n513 VSUBS 0.008894f
C708 B.n514 VSUBS 0.008894f
C709 B.n515 VSUBS 0.008894f
C710 B.n516 VSUBS 0.008894f
C711 B.n517 VSUBS 0.008894f
C712 B.n518 VSUBS 0.008894f
C713 B.n519 VSUBS 0.008894f
C714 B.n520 VSUBS 0.008894f
C715 B.n521 VSUBS 0.008894f
C716 B.n522 VSUBS 0.008894f
C717 B.n523 VSUBS 0.008894f
C718 B.n524 VSUBS 0.008894f
C719 B.n525 VSUBS 0.008894f
C720 B.n526 VSUBS 0.008894f
C721 B.n527 VSUBS 0.008894f
C722 B.n528 VSUBS 0.008894f
C723 B.n529 VSUBS 0.008894f
C724 B.n530 VSUBS 0.008894f
C725 B.n531 VSUBS 0.008894f
C726 B.n532 VSUBS 0.008894f
C727 B.n533 VSUBS 0.008894f
C728 B.n534 VSUBS 0.008894f
C729 B.n535 VSUBS 0.008894f
C730 B.n536 VSUBS 0.008894f
C731 B.n537 VSUBS 0.008894f
C732 B.n538 VSUBS 0.008894f
C733 B.n539 VSUBS 0.008894f
C734 B.n540 VSUBS 0.008894f
C735 B.n541 VSUBS 0.008894f
C736 B.n542 VSUBS 0.008894f
C737 B.n543 VSUBS 0.008894f
C738 B.n544 VSUBS 0.008894f
C739 B.n545 VSUBS 0.008894f
C740 B.n546 VSUBS 0.008894f
C741 B.n547 VSUBS 0.008894f
C742 B.n548 VSUBS 0.008894f
C743 B.n549 VSUBS 0.008894f
C744 B.n550 VSUBS 0.008894f
C745 B.n551 VSUBS 0.008894f
C746 B.n552 VSUBS 0.008894f
C747 B.n553 VSUBS 0.008894f
C748 B.n554 VSUBS 0.008894f
C749 B.n555 VSUBS 0.008894f
C750 B.n556 VSUBS 0.008894f
C751 B.n557 VSUBS 0.008894f
C752 B.n558 VSUBS 0.008894f
C753 B.n559 VSUBS 0.008894f
C754 B.n560 VSUBS 0.008894f
C755 B.n561 VSUBS 0.008894f
C756 B.n562 VSUBS 0.008894f
C757 B.n563 VSUBS 0.008894f
C758 B.n564 VSUBS 0.008894f
C759 B.n565 VSUBS 0.008894f
C760 B.n566 VSUBS 0.008894f
C761 B.n567 VSUBS 0.008894f
C762 B.n568 VSUBS 0.008894f
C763 B.n569 VSUBS 0.008894f
C764 B.n570 VSUBS 0.008894f
C765 B.n571 VSUBS 0.008894f
C766 B.n572 VSUBS 0.008894f
C767 B.n573 VSUBS 0.008894f
C768 B.n574 VSUBS 0.008894f
C769 B.n575 VSUBS 0.008894f
C770 B.n576 VSUBS 0.008894f
C771 B.n577 VSUBS 0.008894f
C772 B.n578 VSUBS 0.008894f
C773 B.n579 VSUBS 0.008894f
C774 B.n580 VSUBS 0.008894f
C775 B.n581 VSUBS 0.020156f
C776 B.n582 VSUBS 0.020914f
C777 B.n583 VSUBS 0.020914f
C778 B.n584 VSUBS 0.008894f
C779 B.n585 VSUBS 0.008894f
C780 B.n586 VSUBS 0.008894f
C781 B.n587 VSUBS 0.008894f
C782 B.n588 VSUBS 0.008894f
C783 B.n589 VSUBS 0.008894f
C784 B.n590 VSUBS 0.008894f
C785 B.n591 VSUBS 0.008894f
C786 B.n592 VSUBS 0.008894f
C787 B.n593 VSUBS 0.008894f
C788 B.n594 VSUBS 0.008894f
C789 B.n595 VSUBS 0.008894f
C790 B.n596 VSUBS 0.008894f
C791 B.n597 VSUBS 0.008894f
C792 B.n598 VSUBS 0.008894f
C793 B.n599 VSUBS 0.008894f
C794 B.n600 VSUBS 0.008894f
C795 B.n601 VSUBS 0.008894f
C796 B.n602 VSUBS 0.008894f
C797 B.n603 VSUBS 0.008894f
C798 B.n604 VSUBS 0.008894f
C799 B.n605 VSUBS 0.008894f
C800 B.n606 VSUBS 0.008894f
C801 B.n607 VSUBS 0.008894f
C802 B.n608 VSUBS 0.008894f
C803 B.n609 VSUBS 0.008894f
C804 B.n610 VSUBS 0.008894f
C805 B.n611 VSUBS 0.008894f
C806 B.n612 VSUBS 0.008894f
C807 B.n613 VSUBS 0.008894f
C808 B.n614 VSUBS 0.008894f
C809 B.n615 VSUBS 0.008894f
C810 B.n616 VSUBS 0.008894f
C811 B.n617 VSUBS 0.008894f
C812 B.n618 VSUBS 0.008894f
C813 B.n619 VSUBS 0.008894f
C814 B.n620 VSUBS 0.008894f
C815 B.n621 VSUBS 0.008894f
C816 B.n622 VSUBS 0.008894f
C817 B.n623 VSUBS 0.008894f
C818 B.n624 VSUBS 0.008894f
C819 B.n625 VSUBS 0.008894f
C820 B.n626 VSUBS 0.008894f
C821 B.n627 VSUBS 0.008894f
C822 B.n628 VSUBS 0.008894f
C823 B.n629 VSUBS 0.008894f
C824 B.n630 VSUBS 0.008894f
C825 B.n631 VSUBS 0.008894f
C826 B.n632 VSUBS 0.008894f
C827 B.n633 VSUBS 0.008894f
C828 B.n634 VSUBS 0.008894f
C829 B.n635 VSUBS 0.008894f
C830 B.n636 VSUBS 0.008894f
C831 B.n637 VSUBS 0.008371f
C832 B.n638 VSUBS 0.020607f
C833 B.n639 VSUBS 0.00497f
C834 B.n640 VSUBS 0.008894f
C835 B.n641 VSUBS 0.008894f
C836 B.n642 VSUBS 0.008894f
C837 B.n643 VSUBS 0.008894f
C838 B.n644 VSUBS 0.008894f
C839 B.n645 VSUBS 0.008894f
C840 B.n646 VSUBS 0.008894f
C841 B.n647 VSUBS 0.008894f
C842 B.n648 VSUBS 0.008894f
C843 B.n649 VSUBS 0.008894f
C844 B.n650 VSUBS 0.008894f
C845 B.n651 VSUBS 0.008894f
C846 B.n652 VSUBS 0.00497f
C847 B.n653 VSUBS 0.008894f
C848 B.n654 VSUBS 0.008894f
C849 B.n655 VSUBS 0.008371f
C850 B.n656 VSUBS 0.008894f
C851 B.n657 VSUBS 0.008894f
C852 B.n658 VSUBS 0.008894f
C853 B.n659 VSUBS 0.008894f
C854 B.n660 VSUBS 0.008894f
C855 B.n661 VSUBS 0.008894f
C856 B.n662 VSUBS 0.008894f
C857 B.n663 VSUBS 0.008894f
C858 B.n664 VSUBS 0.008894f
C859 B.n665 VSUBS 0.008894f
C860 B.n666 VSUBS 0.008894f
C861 B.n667 VSUBS 0.008894f
C862 B.n668 VSUBS 0.008894f
C863 B.n669 VSUBS 0.008894f
C864 B.n670 VSUBS 0.008894f
C865 B.n671 VSUBS 0.008894f
C866 B.n672 VSUBS 0.008894f
C867 B.n673 VSUBS 0.008894f
C868 B.n674 VSUBS 0.008894f
C869 B.n675 VSUBS 0.008894f
C870 B.n676 VSUBS 0.008894f
C871 B.n677 VSUBS 0.008894f
C872 B.n678 VSUBS 0.008894f
C873 B.n679 VSUBS 0.008894f
C874 B.n680 VSUBS 0.008894f
C875 B.n681 VSUBS 0.008894f
C876 B.n682 VSUBS 0.008894f
C877 B.n683 VSUBS 0.008894f
C878 B.n684 VSUBS 0.008894f
C879 B.n685 VSUBS 0.008894f
C880 B.n686 VSUBS 0.008894f
C881 B.n687 VSUBS 0.008894f
C882 B.n688 VSUBS 0.008894f
C883 B.n689 VSUBS 0.008894f
C884 B.n690 VSUBS 0.008894f
C885 B.n691 VSUBS 0.008894f
C886 B.n692 VSUBS 0.008894f
C887 B.n693 VSUBS 0.008894f
C888 B.n694 VSUBS 0.008894f
C889 B.n695 VSUBS 0.008894f
C890 B.n696 VSUBS 0.008894f
C891 B.n697 VSUBS 0.008894f
C892 B.n698 VSUBS 0.008894f
C893 B.n699 VSUBS 0.008894f
C894 B.n700 VSUBS 0.008894f
C895 B.n701 VSUBS 0.008894f
C896 B.n702 VSUBS 0.008894f
C897 B.n703 VSUBS 0.008894f
C898 B.n704 VSUBS 0.008894f
C899 B.n705 VSUBS 0.008894f
C900 B.n706 VSUBS 0.008894f
C901 B.n707 VSUBS 0.008894f
C902 B.n708 VSUBS 0.020914f
C903 B.n709 VSUBS 0.020914f
C904 B.n710 VSUBS 0.020156f
C905 B.n711 VSUBS 0.008894f
C906 B.n712 VSUBS 0.008894f
C907 B.n713 VSUBS 0.008894f
C908 B.n714 VSUBS 0.008894f
C909 B.n715 VSUBS 0.008894f
C910 B.n716 VSUBS 0.008894f
C911 B.n717 VSUBS 0.008894f
C912 B.n718 VSUBS 0.008894f
C913 B.n719 VSUBS 0.008894f
C914 B.n720 VSUBS 0.008894f
C915 B.n721 VSUBS 0.008894f
C916 B.n722 VSUBS 0.008894f
C917 B.n723 VSUBS 0.008894f
C918 B.n724 VSUBS 0.008894f
C919 B.n725 VSUBS 0.008894f
C920 B.n726 VSUBS 0.008894f
C921 B.n727 VSUBS 0.008894f
C922 B.n728 VSUBS 0.008894f
C923 B.n729 VSUBS 0.008894f
C924 B.n730 VSUBS 0.008894f
C925 B.n731 VSUBS 0.008894f
C926 B.n732 VSUBS 0.008894f
C927 B.n733 VSUBS 0.008894f
C928 B.n734 VSUBS 0.008894f
C929 B.n735 VSUBS 0.008894f
C930 B.n736 VSUBS 0.008894f
C931 B.n737 VSUBS 0.008894f
C932 B.n738 VSUBS 0.008894f
C933 B.n739 VSUBS 0.008894f
C934 B.n740 VSUBS 0.008894f
C935 B.n741 VSUBS 0.008894f
C936 B.n742 VSUBS 0.008894f
C937 B.n743 VSUBS 0.008894f
C938 B.n744 VSUBS 0.008894f
C939 B.n745 VSUBS 0.008894f
C940 B.n746 VSUBS 0.008894f
C941 B.n747 VSUBS 0.008894f
C942 B.n748 VSUBS 0.008894f
C943 B.n749 VSUBS 0.008894f
C944 B.n750 VSUBS 0.008894f
C945 B.n751 VSUBS 0.008894f
C946 B.n752 VSUBS 0.008894f
C947 B.n753 VSUBS 0.008894f
C948 B.n754 VSUBS 0.008894f
C949 B.n755 VSUBS 0.008894f
C950 B.n756 VSUBS 0.008894f
C951 B.n757 VSUBS 0.008894f
C952 B.n758 VSUBS 0.008894f
C953 B.n759 VSUBS 0.008894f
C954 B.n760 VSUBS 0.008894f
C955 B.n761 VSUBS 0.008894f
C956 B.n762 VSUBS 0.008894f
C957 B.n763 VSUBS 0.008894f
C958 B.n764 VSUBS 0.008894f
C959 B.n765 VSUBS 0.008894f
C960 B.n766 VSUBS 0.008894f
C961 B.n767 VSUBS 0.008894f
C962 B.n768 VSUBS 0.008894f
C963 B.n769 VSUBS 0.008894f
C964 B.n770 VSUBS 0.008894f
C965 B.n771 VSUBS 0.008894f
C966 B.n772 VSUBS 0.008894f
C967 B.n773 VSUBS 0.008894f
C968 B.n774 VSUBS 0.008894f
C969 B.n775 VSUBS 0.008894f
C970 B.n776 VSUBS 0.008894f
C971 B.n777 VSUBS 0.008894f
C972 B.n778 VSUBS 0.008894f
C973 B.n779 VSUBS 0.008894f
C974 B.n780 VSUBS 0.008894f
C975 B.n781 VSUBS 0.008894f
C976 B.n782 VSUBS 0.008894f
C977 B.n783 VSUBS 0.008894f
C978 B.n784 VSUBS 0.008894f
C979 B.n785 VSUBS 0.008894f
C980 B.n786 VSUBS 0.008894f
C981 B.n787 VSUBS 0.008894f
C982 B.n788 VSUBS 0.008894f
C983 B.n789 VSUBS 0.008894f
C984 B.n790 VSUBS 0.008894f
C985 B.n791 VSUBS 0.011606f
C986 B.n792 VSUBS 0.012364f
C987 B.n793 VSUBS 0.024586f
.ends

