* NGSPICE file created from diff_pair_sample_0090.ext - technology: sky130A

.subckt diff_pair_sample_0090 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=0.47
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=0.47
X2 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=0.47
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=0.47
X4 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=0.47
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=0.47
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=0.47
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=0.47
R0 B.n323 B.n322 585
R1 B.n324 B.n323 585
R2 B.n133 B.n48 585
R3 B.n132 B.n131 585
R4 B.n130 B.n129 585
R5 B.n128 B.n127 585
R6 B.n126 B.n125 585
R7 B.n124 B.n123 585
R8 B.n122 B.n121 585
R9 B.n120 B.n119 585
R10 B.n118 B.n117 585
R11 B.n116 B.n115 585
R12 B.n114 B.n113 585
R13 B.n112 B.n111 585
R14 B.n110 B.n109 585
R15 B.n108 B.n107 585
R16 B.n106 B.n105 585
R17 B.n103 B.n102 585
R18 B.n101 B.n100 585
R19 B.n99 B.n98 585
R20 B.n97 B.n96 585
R21 B.n95 B.n94 585
R22 B.n93 B.n92 585
R23 B.n91 B.n90 585
R24 B.n89 B.n88 585
R25 B.n87 B.n86 585
R26 B.n85 B.n84 585
R27 B.n83 B.n82 585
R28 B.n81 B.n80 585
R29 B.n79 B.n78 585
R30 B.n77 B.n76 585
R31 B.n75 B.n74 585
R32 B.n73 B.n72 585
R33 B.n71 B.n70 585
R34 B.n69 B.n68 585
R35 B.n67 B.n66 585
R36 B.n65 B.n64 585
R37 B.n63 B.n62 585
R38 B.n61 B.n60 585
R39 B.n59 B.n58 585
R40 B.n57 B.n56 585
R41 B.n55 B.n54 585
R42 B.n321 B.n27 585
R43 B.n325 B.n27 585
R44 B.n320 B.n26 585
R45 B.n326 B.n26 585
R46 B.n319 B.n318 585
R47 B.n318 B.n22 585
R48 B.n317 B.n21 585
R49 B.n332 B.n21 585
R50 B.n316 B.n20 585
R51 B.n333 B.n20 585
R52 B.n315 B.n19 585
R53 B.n334 B.n19 585
R54 B.n314 B.n313 585
R55 B.n313 B.n15 585
R56 B.n312 B.n14 585
R57 B.n340 B.n14 585
R58 B.n311 B.n13 585
R59 B.n341 B.n13 585
R60 B.n310 B.n12 585
R61 B.n342 B.n12 585
R62 B.n309 B.n308 585
R63 B.n308 B.n11 585
R64 B.n307 B.n7 585
R65 B.n348 B.n7 585
R66 B.n306 B.n6 585
R67 B.n349 B.n6 585
R68 B.n305 B.n5 585
R69 B.n350 B.n5 585
R70 B.n304 B.n303 585
R71 B.n303 B.n4 585
R72 B.n302 B.n134 585
R73 B.n302 B.n301 585
R74 B.n291 B.n135 585
R75 B.n294 B.n135 585
R76 B.n293 B.n292 585
R77 B.n295 B.n293 585
R78 B.n290 B.n140 585
R79 B.n140 B.n139 585
R80 B.n289 B.n288 585
R81 B.n288 B.n287 585
R82 B.n142 B.n141 585
R83 B.n143 B.n142 585
R84 B.n280 B.n279 585
R85 B.n281 B.n280 585
R86 B.n278 B.n147 585
R87 B.n151 B.n147 585
R88 B.n277 B.n276 585
R89 B.n276 B.n275 585
R90 B.n149 B.n148 585
R91 B.n150 B.n149 585
R92 B.n268 B.n267 585
R93 B.n269 B.n268 585
R94 B.n266 B.n156 585
R95 B.n156 B.n155 585
R96 B.n260 B.n259 585
R97 B.n258 B.n178 585
R98 B.n257 B.n177 585
R99 B.n262 B.n177 585
R100 B.n256 B.n255 585
R101 B.n254 B.n253 585
R102 B.n252 B.n251 585
R103 B.n250 B.n249 585
R104 B.n248 B.n247 585
R105 B.n246 B.n245 585
R106 B.n244 B.n243 585
R107 B.n242 B.n241 585
R108 B.n240 B.n239 585
R109 B.n238 B.n237 585
R110 B.n236 B.n235 585
R111 B.n234 B.n233 585
R112 B.n232 B.n231 585
R113 B.n229 B.n228 585
R114 B.n227 B.n226 585
R115 B.n225 B.n224 585
R116 B.n223 B.n222 585
R117 B.n221 B.n220 585
R118 B.n219 B.n218 585
R119 B.n217 B.n216 585
R120 B.n215 B.n214 585
R121 B.n213 B.n212 585
R122 B.n211 B.n210 585
R123 B.n209 B.n208 585
R124 B.n207 B.n206 585
R125 B.n205 B.n204 585
R126 B.n203 B.n202 585
R127 B.n201 B.n200 585
R128 B.n199 B.n198 585
R129 B.n197 B.n196 585
R130 B.n195 B.n194 585
R131 B.n193 B.n192 585
R132 B.n191 B.n190 585
R133 B.n189 B.n188 585
R134 B.n187 B.n186 585
R135 B.n185 B.n184 585
R136 B.n158 B.n157 585
R137 B.n265 B.n264 585
R138 B.n154 B.n153 585
R139 B.n155 B.n154 585
R140 B.n271 B.n270 585
R141 B.n270 B.n269 585
R142 B.n272 B.n152 585
R143 B.n152 B.n150 585
R144 B.n274 B.n273 585
R145 B.n275 B.n274 585
R146 B.n146 B.n145 585
R147 B.n151 B.n146 585
R148 B.n283 B.n282 585
R149 B.n282 B.n281 585
R150 B.n284 B.n144 585
R151 B.n144 B.n143 585
R152 B.n286 B.n285 585
R153 B.n287 B.n286 585
R154 B.n138 B.n137 585
R155 B.n139 B.n138 585
R156 B.n297 B.n296 585
R157 B.n296 B.n295 585
R158 B.n298 B.n136 585
R159 B.n294 B.n136 585
R160 B.n300 B.n299 585
R161 B.n301 B.n300 585
R162 B.n2 B.n0 585
R163 B.n4 B.n2 585
R164 B.n3 B.n1 585
R165 B.n349 B.n3 585
R166 B.n347 B.n346 585
R167 B.n348 B.n347 585
R168 B.n345 B.n8 585
R169 B.n11 B.n8 585
R170 B.n344 B.n343 585
R171 B.n343 B.n342 585
R172 B.n10 B.n9 585
R173 B.n341 B.n10 585
R174 B.n339 B.n338 585
R175 B.n340 B.n339 585
R176 B.n337 B.n16 585
R177 B.n16 B.n15 585
R178 B.n336 B.n335 585
R179 B.n335 B.n334 585
R180 B.n18 B.n17 585
R181 B.n333 B.n18 585
R182 B.n331 B.n330 585
R183 B.n332 B.n331 585
R184 B.n329 B.n23 585
R185 B.n23 B.n22 585
R186 B.n328 B.n327 585
R187 B.n327 B.n326 585
R188 B.n25 B.n24 585
R189 B.n325 B.n25 585
R190 B.n352 B.n351 585
R191 B.n351 B.n350 585
R192 B.n260 B.n154 473.281
R193 B.n54 B.n25 473.281
R194 B.n264 B.n156 473.281
R195 B.n323 B.n27 473.281
R196 B.n181 B.t6 370.236
R197 B.n179 B.t13 370.236
R198 B.n51 B.t10 370.236
R199 B.n49 B.t2 370.236
R200 B.n324 B.n47 256.663
R201 B.n324 B.n46 256.663
R202 B.n324 B.n45 256.663
R203 B.n324 B.n44 256.663
R204 B.n324 B.n43 256.663
R205 B.n324 B.n42 256.663
R206 B.n324 B.n41 256.663
R207 B.n324 B.n40 256.663
R208 B.n324 B.n39 256.663
R209 B.n324 B.n38 256.663
R210 B.n324 B.n37 256.663
R211 B.n324 B.n36 256.663
R212 B.n324 B.n35 256.663
R213 B.n324 B.n34 256.663
R214 B.n324 B.n33 256.663
R215 B.n324 B.n32 256.663
R216 B.n324 B.n31 256.663
R217 B.n324 B.n30 256.663
R218 B.n324 B.n29 256.663
R219 B.n324 B.n28 256.663
R220 B.n262 B.n261 256.663
R221 B.n262 B.n159 256.663
R222 B.n262 B.n160 256.663
R223 B.n262 B.n161 256.663
R224 B.n262 B.n162 256.663
R225 B.n262 B.n163 256.663
R226 B.n262 B.n164 256.663
R227 B.n262 B.n165 256.663
R228 B.n262 B.n166 256.663
R229 B.n262 B.n167 256.663
R230 B.n262 B.n168 256.663
R231 B.n262 B.n169 256.663
R232 B.n262 B.n170 256.663
R233 B.n262 B.n171 256.663
R234 B.n262 B.n172 256.663
R235 B.n262 B.n173 256.663
R236 B.n262 B.n174 256.663
R237 B.n262 B.n175 256.663
R238 B.n262 B.n176 256.663
R239 B.n263 B.n262 256.663
R240 B.n270 B.n154 163.367
R241 B.n270 B.n152 163.367
R242 B.n274 B.n152 163.367
R243 B.n274 B.n146 163.367
R244 B.n282 B.n146 163.367
R245 B.n282 B.n144 163.367
R246 B.n286 B.n144 163.367
R247 B.n286 B.n138 163.367
R248 B.n296 B.n138 163.367
R249 B.n296 B.n136 163.367
R250 B.n300 B.n136 163.367
R251 B.n300 B.n2 163.367
R252 B.n351 B.n2 163.367
R253 B.n351 B.n3 163.367
R254 B.n347 B.n3 163.367
R255 B.n347 B.n8 163.367
R256 B.n343 B.n8 163.367
R257 B.n343 B.n10 163.367
R258 B.n339 B.n10 163.367
R259 B.n339 B.n16 163.367
R260 B.n335 B.n16 163.367
R261 B.n335 B.n18 163.367
R262 B.n331 B.n18 163.367
R263 B.n331 B.n23 163.367
R264 B.n327 B.n23 163.367
R265 B.n327 B.n25 163.367
R266 B.n178 B.n177 163.367
R267 B.n255 B.n177 163.367
R268 B.n253 B.n252 163.367
R269 B.n249 B.n248 163.367
R270 B.n245 B.n244 163.367
R271 B.n241 B.n240 163.367
R272 B.n237 B.n236 163.367
R273 B.n233 B.n232 163.367
R274 B.n228 B.n227 163.367
R275 B.n224 B.n223 163.367
R276 B.n220 B.n219 163.367
R277 B.n216 B.n215 163.367
R278 B.n212 B.n211 163.367
R279 B.n208 B.n207 163.367
R280 B.n204 B.n203 163.367
R281 B.n200 B.n199 163.367
R282 B.n196 B.n195 163.367
R283 B.n192 B.n191 163.367
R284 B.n188 B.n187 163.367
R285 B.n184 B.n158 163.367
R286 B.n268 B.n156 163.367
R287 B.n268 B.n149 163.367
R288 B.n276 B.n149 163.367
R289 B.n276 B.n147 163.367
R290 B.n280 B.n147 163.367
R291 B.n280 B.n142 163.367
R292 B.n288 B.n142 163.367
R293 B.n288 B.n140 163.367
R294 B.n293 B.n140 163.367
R295 B.n293 B.n135 163.367
R296 B.n302 B.n135 163.367
R297 B.n303 B.n302 163.367
R298 B.n303 B.n5 163.367
R299 B.n6 B.n5 163.367
R300 B.n7 B.n6 163.367
R301 B.n308 B.n7 163.367
R302 B.n308 B.n12 163.367
R303 B.n13 B.n12 163.367
R304 B.n14 B.n13 163.367
R305 B.n313 B.n14 163.367
R306 B.n313 B.n19 163.367
R307 B.n20 B.n19 163.367
R308 B.n21 B.n20 163.367
R309 B.n318 B.n21 163.367
R310 B.n318 B.n26 163.367
R311 B.n27 B.n26 163.367
R312 B.n58 B.n57 163.367
R313 B.n62 B.n61 163.367
R314 B.n66 B.n65 163.367
R315 B.n70 B.n69 163.367
R316 B.n74 B.n73 163.367
R317 B.n78 B.n77 163.367
R318 B.n82 B.n81 163.367
R319 B.n86 B.n85 163.367
R320 B.n90 B.n89 163.367
R321 B.n94 B.n93 163.367
R322 B.n98 B.n97 163.367
R323 B.n102 B.n101 163.367
R324 B.n107 B.n106 163.367
R325 B.n111 B.n110 163.367
R326 B.n115 B.n114 163.367
R327 B.n119 B.n118 163.367
R328 B.n123 B.n122 163.367
R329 B.n127 B.n126 163.367
R330 B.n131 B.n130 163.367
R331 B.n323 B.n48 163.367
R332 B.n181 B.t9 147.306
R333 B.n49 B.t4 147.306
R334 B.n179 B.t15 147.306
R335 B.n51 B.t11 147.306
R336 B.n262 B.n155 144.071
R337 B.n325 B.n324 144.071
R338 B.n182 B.t8 131.792
R339 B.n50 B.t5 131.792
R340 B.n180 B.t14 131.792
R341 B.n52 B.t12 131.792
R342 B.n269 B.n155 88.2601
R343 B.n269 B.n150 88.2601
R344 B.n275 B.n150 88.2601
R345 B.n275 B.n151 88.2601
R346 B.n281 B.n143 88.2601
R347 B.n287 B.n143 88.2601
R348 B.n287 B.n139 88.2601
R349 B.n295 B.n139 88.2601
R350 B.n295 B.n294 88.2601
R351 B.n301 B.n4 88.2601
R352 B.n350 B.n4 88.2601
R353 B.n350 B.n349 88.2601
R354 B.n349 B.n348 88.2601
R355 B.n342 B.n11 88.2601
R356 B.n342 B.n341 88.2601
R357 B.n341 B.n340 88.2601
R358 B.n340 B.n15 88.2601
R359 B.n334 B.n15 88.2601
R360 B.n333 B.n332 88.2601
R361 B.n332 B.n22 88.2601
R362 B.n326 B.n22 88.2601
R363 B.n326 B.n325 88.2601
R364 B.n261 B.n260 71.676
R365 B.n255 B.n159 71.676
R366 B.n252 B.n160 71.676
R367 B.n248 B.n161 71.676
R368 B.n244 B.n162 71.676
R369 B.n240 B.n163 71.676
R370 B.n236 B.n164 71.676
R371 B.n232 B.n165 71.676
R372 B.n227 B.n166 71.676
R373 B.n223 B.n167 71.676
R374 B.n219 B.n168 71.676
R375 B.n215 B.n169 71.676
R376 B.n211 B.n170 71.676
R377 B.n207 B.n171 71.676
R378 B.n203 B.n172 71.676
R379 B.n199 B.n173 71.676
R380 B.n195 B.n174 71.676
R381 B.n191 B.n175 71.676
R382 B.n187 B.n176 71.676
R383 B.n263 B.n158 71.676
R384 B.n54 B.n28 71.676
R385 B.n58 B.n29 71.676
R386 B.n62 B.n30 71.676
R387 B.n66 B.n31 71.676
R388 B.n70 B.n32 71.676
R389 B.n74 B.n33 71.676
R390 B.n78 B.n34 71.676
R391 B.n82 B.n35 71.676
R392 B.n86 B.n36 71.676
R393 B.n90 B.n37 71.676
R394 B.n94 B.n38 71.676
R395 B.n98 B.n39 71.676
R396 B.n102 B.n40 71.676
R397 B.n107 B.n41 71.676
R398 B.n111 B.n42 71.676
R399 B.n115 B.n43 71.676
R400 B.n119 B.n44 71.676
R401 B.n123 B.n45 71.676
R402 B.n127 B.n46 71.676
R403 B.n131 B.n47 71.676
R404 B.n48 B.n47 71.676
R405 B.n130 B.n46 71.676
R406 B.n126 B.n45 71.676
R407 B.n122 B.n44 71.676
R408 B.n118 B.n43 71.676
R409 B.n114 B.n42 71.676
R410 B.n110 B.n41 71.676
R411 B.n106 B.n40 71.676
R412 B.n101 B.n39 71.676
R413 B.n97 B.n38 71.676
R414 B.n93 B.n37 71.676
R415 B.n89 B.n36 71.676
R416 B.n85 B.n35 71.676
R417 B.n81 B.n34 71.676
R418 B.n77 B.n33 71.676
R419 B.n73 B.n32 71.676
R420 B.n69 B.n31 71.676
R421 B.n65 B.n30 71.676
R422 B.n61 B.n29 71.676
R423 B.n57 B.n28 71.676
R424 B.n261 B.n178 71.676
R425 B.n253 B.n159 71.676
R426 B.n249 B.n160 71.676
R427 B.n245 B.n161 71.676
R428 B.n241 B.n162 71.676
R429 B.n237 B.n163 71.676
R430 B.n233 B.n164 71.676
R431 B.n228 B.n165 71.676
R432 B.n224 B.n166 71.676
R433 B.n220 B.n167 71.676
R434 B.n216 B.n168 71.676
R435 B.n212 B.n169 71.676
R436 B.n208 B.n170 71.676
R437 B.n204 B.n171 71.676
R438 B.n200 B.n172 71.676
R439 B.n196 B.n173 71.676
R440 B.n192 B.n174 71.676
R441 B.n188 B.n175 71.676
R442 B.n184 B.n176 71.676
R443 B.n264 B.n263 71.676
R444 B.n301 B.t1 68.7911
R445 B.n348 B.t0 68.7911
R446 B.n183 B.n182 59.5399
R447 B.n230 B.n180 59.5399
R448 B.n53 B.n52 59.5399
R449 B.n104 B.n50 59.5399
R450 B.n151 B.t7 58.4076
R451 B.t3 B.n333 58.4076
R452 B.n55 B.n24 30.7517
R453 B.n266 B.n265 30.7517
R454 B.n259 B.n153 30.7517
R455 B.n322 B.n321 30.7517
R456 B.n281 B.t7 29.853
R457 B.n334 B.t3 29.853
R458 B.n294 B.t1 19.4695
R459 B.n11 B.t0 19.4695
R460 B B.n352 18.0485
R461 B.n182 B.n181 15.5157
R462 B.n180 B.n179 15.5157
R463 B.n52 B.n51 15.5157
R464 B.n50 B.n49 15.5157
R465 B.n56 B.n55 10.6151
R466 B.n59 B.n56 10.6151
R467 B.n60 B.n59 10.6151
R468 B.n63 B.n60 10.6151
R469 B.n64 B.n63 10.6151
R470 B.n67 B.n64 10.6151
R471 B.n68 B.n67 10.6151
R472 B.n71 B.n68 10.6151
R473 B.n72 B.n71 10.6151
R474 B.n75 B.n72 10.6151
R475 B.n76 B.n75 10.6151
R476 B.n79 B.n76 10.6151
R477 B.n80 B.n79 10.6151
R478 B.n83 B.n80 10.6151
R479 B.n84 B.n83 10.6151
R480 B.n88 B.n87 10.6151
R481 B.n91 B.n88 10.6151
R482 B.n92 B.n91 10.6151
R483 B.n95 B.n92 10.6151
R484 B.n96 B.n95 10.6151
R485 B.n99 B.n96 10.6151
R486 B.n100 B.n99 10.6151
R487 B.n103 B.n100 10.6151
R488 B.n108 B.n105 10.6151
R489 B.n109 B.n108 10.6151
R490 B.n112 B.n109 10.6151
R491 B.n113 B.n112 10.6151
R492 B.n116 B.n113 10.6151
R493 B.n117 B.n116 10.6151
R494 B.n120 B.n117 10.6151
R495 B.n121 B.n120 10.6151
R496 B.n124 B.n121 10.6151
R497 B.n125 B.n124 10.6151
R498 B.n128 B.n125 10.6151
R499 B.n129 B.n128 10.6151
R500 B.n132 B.n129 10.6151
R501 B.n133 B.n132 10.6151
R502 B.n322 B.n133 10.6151
R503 B.n267 B.n266 10.6151
R504 B.n267 B.n148 10.6151
R505 B.n277 B.n148 10.6151
R506 B.n278 B.n277 10.6151
R507 B.n279 B.n278 10.6151
R508 B.n279 B.n141 10.6151
R509 B.n289 B.n141 10.6151
R510 B.n290 B.n289 10.6151
R511 B.n292 B.n290 10.6151
R512 B.n292 B.n291 10.6151
R513 B.n291 B.n134 10.6151
R514 B.n304 B.n134 10.6151
R515 B.n305 B.n304 10.6151
R516 B.n306 B.n305 10.6151
R517 B.n307 B.n306 10.6151
R518 B.n309 B.n307 10.6151
R519 B.n310 B.n309 10.6151
R520 B.n311 B.n310 10.6151
R521 B.n312 B.n311 10.6151
R522 B.n314 B.n312 10.6151
R523 B.n315 B.n314 10.6151
R524 B.n316 B.n315 10.6151
R525 B.n317 B.n316 10.6151
R526 B.n319 B.n317 10.6151
R527 B.n320 B.n319 10.6151
R528 B.n321 B.n320 10.6151
R529 B.n259 B.n258 10.6151
R530 B.n258 B.n257 10.6151
R531 B.n257 B.n256 10.6151
R532 B.n256 B.n254 10.6151
R533 B.n254 B.n251 10.6151
R534 B.n251 B.n250 10.6151
R535 B.n250 B.n247 10.6151
R536 B.n247 B.n246 10.6151
R537 B.n246 B.n243 10.6151
R538 B.n243 B.n242 10.6151
R539 B.n242 B.n239 10.6151
R540 B.n239 B.n238 10.6151
R541 B.n238 B.n235 10.6151
R542 B.n235 B.n234 10.6151
R543 B.n234 B.n231 10.6151
R544 B.n229 B.n226 10.6151
R545 B.n226 B.n225 10.6151
R546 B.n225 B.n222 10.6151
R547 B.n222 B.n221 10.6151
R548 B.n221 B.n218 10.6151
R549 B.n218 B.n217 10.6151
R550 B.n217 B.n214 10.6151
R551 B.n214 B.n213 10.6151
R552 B.n210 B.n209 10.6151
R553 B.n209 B.n206 10.6151
R554 B.n206 B.n205 10.6151
R555 B.n205 B.n202 10.6151
R556 B.n202 B.n201 10.6151
R557 B.n201 B.n198 10.6151
R558 B.n198 B.n197 10.6151
R559 B.n197 B.n194 10.6151
R560 B.n194 B.n193 10.6151
R561 B.n193 B.n190 10.6151
R562 B.n190 B.n189 10.6151
R563 B.n189 B.n186 10.6151
R564 B.n186 B.n185 10.6151
R565 B.n185 B.n157 10.6151
R566 B.n265 B.n157 10.6151
R567 B.n271 B.n153 10.6151
R568 B.n272 B.n271 10.6151
R569 B.n273 B.n272 10.6151
R570 B.n273 B.n145 10.6151
R571 B.n283 B.n145 10.6151
R572 B.n284 B.n283 10.6151
R573 B.n285 B.n284 10.6151
R574 B.n285 B.n137 10.6151
R575 B.n297 B.n137 10.6151
R576 B.n298 B.n297 10.6151
R577 B.n299 B.n298 10.6151
R578 B.n299 B.n0 10.6151
R579 B.n346 B.n1 10.6151
R580 B.n346 B.n345 10.6151
R581 B.n345 B.n344 10.6151
R582 B.n344 B.n9 10.6151
R583 B.n338 B.n9 10.6151
R584 B.n338 B.n337 10.6151
R585 B.n337 B.n336 10.6151
R586 B.n336 B.n17 10.6151
R587 B.n330 B.n17 10.6151
R588 B.n330 B.n329 10.6151
R589 B.n329 B.n328 10.6151
R590 B.n328 B.n24 10.6151
R591 B.n87 B.n53 7.18099
R592 B.n104 B.n103 7.18099
R593 B.n230 B.n229 7.18099
R594 B.n213 B.n183 7.18099
R595 B.n84 B.n53 3.43465
R596 B.n105 B.n104 3.43465
R597 B.n231 B.n230 3.43465
R598 B.n210 B.n183 3.43465
R599 B.n352 B.n0 2.81026
R600 B.n352 B.n1 2.81026
R601 VN VN.t0 440.663
R602 VN VN.t1 407.993
R603 VTAIL.n58 VTAIL.n48 289.615
R604 VTAIL.n10 VTAIL.n0 289.615
R605 VTAIL.n42 VTAIL.n32 289.615
R606 VTAIL.n26 VTAIL.n16 289.615
R607 VTAIL.n52 VTAIL.n51 185
R608 VTAIL.n57 VTAIL.n56 185
R609 VTAIL.n59 VTAIL.n58 185
R610 VTAIL.n4 VTAIL.n3 185
R611 VTAIL.n9 VTAIL.n8 185
R612 VTAIL.n11 VTAIL.n10 185
R613 VTAIL.n43 VTAIL.n42 185
R614 VTAIL.n41 VTAIL.n40 185
R615 VTAIL.n36 VTAIL.n35 185
R616 VTAIL.n27 VTAIL.n26 185
R617 VTAIL.n25 VTAIL.n24 185
R618 VTAIL.n20 VTAIL.n19 185
R619 VTAIL.n53 VTAIL.t3 148.606
R620 VTAIL.n5 VTAIL.t0 148.606
R621 VTAIL.n37 VTAIL.t1 148.606
R622 VTAIL.n21 VTAIL.t2 148.606
R623 VTAIL.n57 VTAIL.n51 104.615
R624 VTAIL.n58 VTAIL.n57 104.615
R625 VTAIL.n9 VTAIL.n3 104.615
R626 VTAIL.n10 VTAIL.n9 104.615
R627 VTAIL.n42 VTAIL.n41 104.615
R628 VTAIL.n41 VTAIL.n35 104.615
R629 VTAIL.n26 VTAIL.n25 104.615
R630 VTAIL.n25 VTAIL.n19 104.615
R631 VTAIL.t3 VTAIL.n51 52.3082
R632 VTAIL.t0 VTAIL.n3 52.3082
R633 VTAIL.t1 VTAIL.n35 52.3082
R634 VTAIL.t2 VTAIL.n19 52.3082
R635 VTAIL.n63 VTAIL.n62 33.349
R636 VTAIL.n15 VTAIL.n14 33.349
R637 VTAIL.n47 VTAIL.n46 33.349
R638 VTAIL.n31 VTAIL.n30 33.349
R639 VTAIL.n31 VTAIL.n15 16.5048
R640 VTAIL.n63 VTAIL.n47 15.8152
R641 VTAIL.n53 VTAIL.n52 15.5966
R642 VTAIL.n5 VTAIL.n4 15.5966
R643 VTAIL.n37 VTAIL.n36 15.5966
R644 VTAIL.n21 VTAIL.n20 15.5966
R645 VTAIL.n56 VTAIL.n55 12.8005
R646 VTAIL.n8 VTAIL.n7 12.8005
R647 VTAIL.n40 VTAIL.n39 12.8005
R648 VTAIL.n24 VTAIL.n23 12.8005
R649 VTAIL.n59 VTAIL.n50 12.0247
R650 VTAIL.n11 VTAIL.n2 12.0247
R651 VTAIL.n43 VTAIL.n34 12.0247
R652 VTAIL.n27 VTAIL.n18 12.0247
R653 VTAIL.n60 VTAIL.n48 11.249
R654 VTAIL.n12 VTAIL.n0 11.249
R655 VTAIL.n44 VTAIL.n32 11.249
R656 VTAIL.n28 VTAIL.n16 11.249
R657 VTAIL.n62 VTAIL.n61 9.45567
R658 VTAIL.n14 VTAIL.n13 9.45567
R659 VTAIL.n46 VTAIL.n45 9.45567
R660 VTAIL.n30 VTAIL.n29 9.45567
R661 VTAIL.n61 VTAIL.n60 9.3005
R662 VTAIL.n50 VTAIL.n49 9.3005
R663 VTAIL.n55 VTAIL.n54 9.3005
R664 VTAIL.n13 VTAIL.n12 9.3005
R665 VTAIL.n2 VTAIL.n1 9.3005
R666 VTAIL.n7 VTAIL.n6 9.3005
R667 VTAIL.n45 VTAIL.n44 9.3005
R668 VTAIL.n34 VTAIL.n33 9.3005
R669 VTAIL.n39 VTAIL.n38 9.3005
R670 VTAIL.n29 VTAIL.n28 9.3005
R671 VTAIL.n18 VTAIL.n17 9.3005
R672 VTAIL.n23 VTAIL.n22 9.3005
R673 VTAIL.n54 VTAIL.n53 4.46457
R674 VTAIL.n6 VTAIL.n5 4.46457
R675 VTAIL.n38 VTAIL.n37 4.46457
R676 VTAIL.n22 VTAIL.n21 4.46457
R677 VTAIL.n62 VTAIL.n48 2.71565
R678 VTAIL.n14 VTAIL.n0 2.71565
R679 VTAIL.n46 VTAIL.n32 2.71565
R680 VTAIL.n30 VTAIL.n16 2.71565
R681 VTAIL.n60 VTAIL.n59 1.93989
R682 VTAIL.n12 VTAIL.n11 1.93989
R683 VTAIL.n44 VTAIL.n43 1.93989
R684 VTAIL.n28 VTAIL.n27 1.93989
R685 VTAIL.n56 VTAIL.n50 1.16414
R686 VTAIL.n8 VTAIL.n2 1.16414
R687 VTAIL.n40 VTAIL.n34 1.16414
R688 VTAIL.n24 VTAIL.n18 1.16414
R689 VTAIL.n47 VTAIL.n31 0.815155
R690 VTAIL VTAIL.n15 0.700931
R691 VTAIL.n55 VTAIL.n52 0.388379
R692 VTAIL.n7 VTAIL.n4 0.388379
R693 VTAIL.n39 VTAIL.n36 0.388379
R694 VTAIL.n23 VTAIL.n20 0.388379
R695 VTAIL.n54 VTAIL.n49 0.155672
R696 VTAIL.n61 VTAIL.n49 0.155672
R697 VTAIL.n6 VTAIL.n1 0.155672
R698 VTAIL.n13 VTAIL.n1 0.155672
R699 VTAIL.n45 VTAIL.n33 0.155672
R700 VTAIL.n38 VTAIL.n33 0.155672
R701 VTAIL.n29 VTAIL.n17 0.155672
R702 VTAIL.n22 VTAIL.n17 0.155672
R703 VTAIL VTAIL.n63 0.114724
R704 VDD2.n25 VDD2.n15 289.615
R705 VDD2.n10 VDD2.n0 289.615
R706 VDD2.n26 VDD2.n25 185
R707 VDD2.n24 VDD2.n23 185
R708 VDD2.n19 VDD2.n18 185
R709 VDD2.n4 VDD2.n3 185
R710 VDD2.n9 VDD2.n8 185
R711 VDD2.n11 VDD2.n10 185
R712 VDD2.n20 VDD2.t1 148.606
R713 VDD2.n5 VDD2.t0 148.606
R714 VDD2.n25 VDD2.n24 104.615
R715 VDD2.n24 VDD2.n18 104.615
R716 VDD2.n9 VDD2.n3 104.615
R717 VDD2.n10 VDD2.n9 104.615
R718 VDD2.n30 VDD2.n14 77.8252
R719 VDD2.t1 VDD2.n18 52.3082
R720 VDD2.t0 VDD2.n3 52.3082
R721 VDD2.n30 VDD2.n29 50.0278
R722 VDD2.n20 VDD2.n19 15.5966
R723 VDD2.n5 VDD2.n4 15.5966
R724 VDD2.n23 VDD2.n22 12.8005
R725 VDD2.n8 VDD2.n7 12.8005
R726 VDD2.n26 VDD2.n17 12.0247
R727 VDD2.n11 VDD2.n2 12.0247
R728 VDD2.n27 VDD2.n15 11.249
R729 VDD2.n12 VDD2.n0 11.249
R730 VDD2.n29 VDD2.n28 9.45567
R731 VDD2.n14 VDD2.n13 9.45567
R732 VDD2.n28 VDD2.n27 9.3005
R733 VDD2.n17 VDD2.n16 9.3005
R734 VDD2.n22 VDD2.n21 9.3005
R735 VDD2.n13 VDD2.n12 9.3005
R736 VDD2.n2 VDD2.n1 9.3005
R737 VDD2.n7 VDD2.n6 9.3005
R738 VDD2.n21 VDD2.n20 4.46457
R739 VDD2.n6 VDD2.n5 4.46457
R740 VDD2.n29 VDD2.n15 2.71565
R741 VDD2.n14 VDD2.n0 2.71565
R742 VDD2.n27 VDD2.n26 1.93989
R743 VDD2.n12 VDD2.n11 1.93989
R744 VDD2.n23 VDD2.n17 1.16414
R745 VDD2.n8 VDD2.n2 1.16414
R746 VDD2.n22 VDD2.n19 0.388379
R747 VDD2.n7 VDD2.n4 0.388379
R748 VDD2 VDD2.n30 0.231103
R749 VDD2.n28 VDD2.n16 0.155672
R750 VDD2.n21 VDD2.n16 0.155672
R751 VDD2.n6 VDD2.n1 0.155672
R752 VDD2.n13 VDD2.n1 0.155672
R753 VP.n0 VP.t0 440.281
R754 VP.n0 VP.t1 407.94
R755 VP VP.n0 0.0516364
R756 VDD1.n10 VDD1.n0 289.615
R757 VDD1.n25 VDD1.n15 289.615
R758 VDD1.n11 VDD1.n10 185
R759 VDD1.n9 VDD1.n8 185
R760 VDD1.n4 VDD1.n3 185
R761 VDD1.n19 VDD1.n18 185
R762 VDD1.n24 VDD1.n23 185
R763 VDD1.n26 VDD1.n25 185
R764 VDD1.n5 VDD1.t1 148.606
R765 VDD1.n20 VDD1.t0 148.606
R766 VDD1.n10 VDD1.n9 104.615
R767 VDD1.n9 VDD1.n3 104.615
R768 VDD1.n24 VDD1.n18 104.615
R769 VDD1.n25 VDD1.n24 104.615
R770 VDD1 VDD1.n29 78.5224
R771 VDD1.t1 VDD1.n3 52.3082
R772 VDD1.t0 VDD1.n18 52.3082
R773 VDD1 VDD1.n14 50.2584
R774 VDD1.n5 VDD1.n4 15.5966
R775 VDD1.n20 VDD1.n19 15.5966
R776 VDD1.n8 VDD1.n7 12.8005
R777 VDD1.n23 VDD1.n22 12.8005
R778 VDD1.n11 VDD1.n2 12.0247
R779 VDD1.n26 VDD1.n17 12.0247
R780 VDD1.n12 VDD1.n0 11.249
R781 VDD1.n27 VDD1.n15 11.249
R782 VDD1.n14 VDD1.n13 9.45567
R783 VDD1.n29 VDD1.n28 9.45567
R784 VDD1.n13 VDD1.n12 9.3005
R785 VDD1.n2 VDD1.n1 9.3005
R786 VDD1.n7 VDD1.n6 9.3005
R787 VDD1.n28 VDD1.n27 9.3005
R788 VDD1.n17 VDD1.n16 9.3005
R789 VDD1.n22 VDD1.n21 9.3005
R790 VDD1.n6 VDD1.n5 4.46457
R791 VDD1.n21 VDD1.n20 4.46457
R792 VDD1.n14 VDD1.n0 2.71565
R793 VDD1.n29 VDD1.n15 2.71565
R794 VDD1.n12 VDD1.n11 1.93989
R795 VDD1.n27 VDD1.n26 1.93989
R796 VDD1.n8 VDD1.n2 1.16414
R797 VDD1.n23 VDD1.n17 1.16414
R798 VDD1.n7 VDD1.n4 0.388379
R799 VDD1.n22 VDD1.n19 0.388379
R800 VDD1.n13 VDD1.n1 0.155672
R801 VDD1.n6 VDD1.n1 0.155672
R802 VDD1.n21 VDD1.n16 0.155672
R803 VDD1.n28 VDD1.n16 0.155672
C0 VP VN 2.82856f
C1 VDD2 VDD1 0.438221f
C2 VDD1 VTAIL 2.49069f
C3 VDD1 VN 0.153721f
C4 VDD1 VP 0.719044f
C5 VDD2 VTAIL 2.52762f
C6 VDD2 VN 0.624919f
C7 VTAIL VN 0.541999f
C8 VDD2 VP 0.249655f
C9 VTAIL VP 0.55626f
C10 VDD2 B 2.061049f
C11 VDD1 B 3.3676f
C12 VTAIL B 2.607353f
C13 VN B 5.419611f
C14 VP B 3.057911f
C15 VDD1.n0 B 0.022702f
C16 VDD1.n1 B 0.016966f
C17 VDD1.n2 B 0.009117f
C18 VDD1.n3 B 0.016161f
C19 VDD1.n4 B 0.012565f
C20 VDD1.t1 B 0.036239f
C21 VDD1.n5 B 0.062469f
C22 VDD1.n6 B 0.181432f
C23 VDD1.n7 B 0.009117f
C24 VDD1.n8 B 0.009653f
C25 VDD1.n9 B 0.021548f
C26 VDD1.n10 B 0.044624f
C27 VDD1.n11 B 0.009653f
C28 VDD1.n12 B 0.009117f
C29 VDD1.n13 B 0.040606f
C30 VDD1.n14 B 0.036718f
C31 VDD1.n15 B 0.022702f
C32 VDD1.n16 B 0.016966f
C33 VDD1.n17 B 0.009117f
C34 VDD1.n18 B 0.016161f
C35 VDD1.n19 B 0.012565f
C36 VDD1.t0 B 0.036239f
C37 VDD1.n20 B 0.062469f
C38 VDD1.n21 B 0.181432f
C39 VDD1.n22 B 0.009117f
C40 VDD1.n23 B 0.009653f
C41 VDD1.n24 B 0.021548f
C42 VDD1.n25 B 0.044624f
C43 VDD1.n26 B 0.009653f
C44 VDD1.n27 B 0.009117f
C45 VDD1.n28 B 0.040606f
C46 VDD1.n29 B 0.24426f
C47 VP.t0 B 0.315218f
C48 VP.t1 B 0.231123f
C49 VP.n0 B 2.24486f
C50 VDD2.n0 B 0.023286f
C51 VDD2.n1 B 0.017402f
C52 VDD2.n2 B 0.009351f
C53 VDD2.n3 B 0.016577f
C54 VDD2.n4 B 0.012888f
C55 VDD2.t0 B 0.03717f
C56 VDD2.n5 B 0.064075f
C57 VDD2.n6 B 0.186096f
C58 VDD2.n7 B 0.009351f
C59 VDD2.n8 B 0.009901f
C60 VDD2.n9 B 0.022102f
C61 VDD2.n10 B 0.045771f
C62 VDD2.n11 B 0.009901f
C63 VDD2.n12 B 0.009351f
C64 VDD2.n13 B 0.04165f
C65 VDD2.n14 B 0.232572f
C66 VDD2.n15 B 0.023286f
C67 VDD2.n16 B 0.017402f
C68 VDD2.n17 B 0.009351f
C69 VDD2.n18 B 0.016577f
C70 VDD2.n19 B 0.012888f
C71 VDD2.t1 B 0.03717f
C72 VDD2.n20 B 0.064075f
C73 VDD2.n21 B 0.186096f
C74 VDD2.n22 B 0.009351f
C75 VDD2.n23 B 0.009901f
C76 VDD2.n24 B 0.022102f
C77 VDD2.n25 B 0.045771f
C78 VDD2.n26 B 0.009901f
C79 VDD2.n27 B 0.009351f
C80 VDD2.n28 B 0.04165f
C81 VDD2.n29 B 0.037445f
C82 VDD2.n30 B 1.16749f
C83 VTAIL.n0 B 0.027702f
C84 VTAIL.n1 B 0.020702f
C85 VTAIL.n2 B 0.011124f
C86 VTAIL.n3 B 0.01972f
C87 VTAIL.n4 B 0.015332f
C88 VTAIL.t0 B 0.04422f
C89 VTAIL.n5 B 0.076227f
C90 VTAIL.n6 B 0.221389f
C91 VTAIL.n7 B 0.011124f
C92 VTAIL.n8 B 0.011779f
C93 VTAIL.n9 B 0.026294f
C94 VTAIL.n10 B 0.054452f
C95 VTAIL.n11 B 0.011779f
C96 VTAIL.n12 B 0.011124f
C97 VTAIL.n13 B 0.049548f
C98 VTAIL.n14 B 0.030265f
C99 VTAIL.n15 B 0.6226f
C100 VTAIL.n16 B 0.027702f
C101 VTAIL.n17 B 0.020702f
C102 VTAIL.n18 B 0.011124f
C103 VTAIL.n19 B 0.01972f
C104 VTAIL.n20 B 0.015332f
C105 VTAIL.t2 B 0.04422f
C106 VTAIL.n21 B 0.076227f
C107 VTAIL.n22 B 0.221389f
C108 VTAIL.n23 B 0.011124f
C109 VTAIL.n24 B 0.011779f
C110 VTAIL.n25 B 0.026294f
C111 VTAIL.n26 B 0.054452f
C112 VTAIL.n27 B 0.011779f
C113 VTAIL.n28 B 0.011124f
C114 VTAIL.n29 B 0.049548f
C115 VTAIL.n30 B 0.030265f
C116 VTAIL.n31 B 0.63022f
C117 VTAIL.n32 B 0.027702f
C118 VTAIL.n33 B 0.020702f
C119 VTAIL.n34 B 0.011124f
C120 VTAIL.n35 B 0.01972f
C121 VTAIL.n36 B 0.015332f
C122 VTAIL.t1 B 0.04422f
C123 VTAIL.n37 B 0.076227f
C124 VTAIL.n38 B 0.221389f
C125 VTAIL.n39 B 0.011124f
C126 VTAIL.n40 B 0.011779f
C127 VTAIL.n41 B 0.026294f
C128 VTAIL.n42 B 0.054452f
C129 VTAIL.n43 B 0.011779f
C130 VTAIL.n44 B 0.011124f
C131 VTAIL.n45 B 0.049548f
C132 VTAIL.n46 B 0.030265f
C133 VTAIL.n47 B 0.584216f
C134 VTAIL.n48 B 0.027702f
C135 VTAIL.n49 B 0.020702f
C136 VTAIL.n50 B 0.011124f
C137 VTAIL.n51 B 0.01972f
C138 VTAIL.n52 B 0.015332f
C139 VTAIL.t3 B 0.04422f
C140 VTAIL.n53 B 0.076227f
C141 VTAIL.n54 B 0.221389f
C142 VTAIL.n55 B 0.011124f
C143 VTAIL.n56 B 0.011779f
C144 VTAIL.n57 B 0.026294f
C145 VTAIL.n58 B 0.054452f
C146 VTAIL.n59 B 0.011779f
C147 VTAIL.n60 B 0.011124f
C148 VTAIL.n61 B 0.049548f
C149 VTAIL.n62 B 0.030265f
C150 VTAIL.n63 B 0.537492f
C151 VN.t1 B 0.226294f
C152 VN.t0 B 0.311586f
.ends

