* NGSPICE file created from diff_pair_sample_1672.ext - technology: sky130A

.subckt diff_pair_sample_1672 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0.54615 ps=3.64 w=3.31 l=1.01
X1 VDD2.t7 VN.t0 VTAIL.t6 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
X2 VTAIL.t2 VN.t1 VDD2.t6 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
X3 VTAIL.t3 VN.t2 VDD2.t5 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0.54615 ps=3.64 w=3.31 l=1.01
X4 VDD1.t7 VP.t1 VTAIL.t14 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=1.2909 ps=7.4 w=3.31 l=1.01
X5 B.t11 B.t9 B.t10 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0 ps=0 w=3.31 l=1.01
X6 VDD2.t4 VN.t3 VTAIL.t7 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=1.2909 ps=7.4 w=3.31 l=1.01
X7 VDD2.t3 VN.t4 VTAIL.t1 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
X8 B.t8 B.t6 B.t7 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0 ps=0 w=3.31 l=1.01
X9 VDD2.t2 VN.t5 VTAIL.t4 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=1.2909 ps=7.4 w=3.31 l=1.01
X10 VDD1.t5 VP.t2 VTAIL.t13 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
X11 B.t5 B.t3 B.t4 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0 ps=0 w=3.31 l=1.01
X12 VTAIL.t0 VN.t6 VDD2.t1 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0.54615 ps=3.64 w=3.31 l=1.01
X13 VDD1.t2 VP.t3 VTAIL.t12 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=1.2909 ps=7.4 w=3.31 l=1.01
X14 VDD1.t0 VP.t4 VTAIL.t11 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
X15 VTAIL.t10 VP.t5 VDD1.t6 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
X16 VTAIL.t9 VP.t6 VDD1.t3 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0.54615 ps=3.64 w=3.31 l=1.01
X17 VTAIL.t8 VP.t7 VDD1.t4 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
X18 B.t2 B.t0 B.t1 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=1.2909 pd=7.4 as=0 ps=0 w=3.31 l=1.01
X19 VTAIL.t5 VN.t7 VDD2.t0 w_n2310_n1630# sky130_fd_pr__pfet_01v8 ad=0.54615 pd=3.64 as=0.54615 ps=3.64 w=3.31 l=1.01
R0 VP.n34 VP.n33 161.3
R1 VP.n11 VP.n10 161.3
R2 VP.n12 VP.n7 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n16 VP.n15 161.3
R5 VP.n17 VP.n5 161.3
R6 VP.n19 VP.n18 161.3
R7 VP.n32 VP.n0 161.3
R8 VP.n31 VP.n30 161.3
R9 VP.n29 VP.n28 161.3
R10 VP.n27 VP.n2 161.3
R11 VP.n26 VP.n25 161.3
R12 VP.n24 VP.n23 161.3
R13 VP.n22 VP.n4 161.3
R14 VP.n21 VP.n20 161.3
R15 VP.n9 VP.t0 133.733
R16 VP.n21 VP.t6 118.115
R17 VP.n33 VP.t3 118.115
R18 VP.n18 VP.t1 118.115
R19 VP.n3 VP.t4 78.9817
R20 VP.n1 VP.t5 78.9817
R21 VP.n6 VP.t7 78.9817
R22 VP.n8 VP.t2 78.9817
R23 VP.n23 VP.n22 56.0336
R24 VP.n32 VP.n31 56.0336
R25 VP.n17 VP.n16 56.0336
R26 VP.n9 VP.n8 46.6347
R27 VP.n10 VP.n9 43.8151
R28 VP.n27 VP.n26 40.4934
R29 VP.n28 VP.n27 40.4934
R30 VP.n13 VP.n12 40.4934
R31 VP.n12 VP.n11 40.4934
R32 VP.n20 VP.n19 36.9096
R33 VP.n23 VP.n3 16.1487
R34 VP.n31 VP.n1 16.1487
R35 VP.n16 VP.n6 16.1487
R36 VP.n26 VP.n3 8.31928
R37 VP.n28 VP.n1 8.31928
R38 VP.n13 VP.n6 8.31928
R39 VP.n11 VP.n8 8.31928
R40 VP.n22 VP.n21 0.730803
R41 VP.n33 VP.n32 0.730803
R42 VP.n18 VP.n17 0.730803
R43 VP.n10 VP.n7 0.189894
R44 VP.n14 VP.n7 0.189894
R45 VP.n15 VP.n14 0.189894
R46 VP.n15 VP.n5 0.189894
R47 VP.n19 VP.n5 0.189894
R48 VP.n20 VP.n4 0.189894
R49 VP.n24 VP.n4 0.189894
R50 VP.n25 VP.n24 0.189894
R51 VP.n25 VP.n2 0.189894
R52 VP.n29 VP.n2 0.189894
R53 VP.n30 VP.n29 0.189894
R54 VP.n30 VP.n0 0.189894
R55 VP.n34 VP.n0 0.189894
R56 VP VP.n34 0.0516364
R57 VDD1 VDD1.n0 132.172
R58 VDD1.n3 VDD1.n2 132.058
R59 VDD1.n3 VDD1.n1 132.058
R60 VDD1.n5 VDD1.n4 131.536
R61 VDD1.n5 VDD1.n3 32.35
R62 VDD1.n4 VDD1.t4 9.82074
R63 VDD1.n4 VDD1.t7 9.82074
R64 VDD1.n0 VDD1.t1 9.82074
R65 VDD1.n0 VDD1.t5 9.82074
R66 VDD1.n2 VDD1.t6 9.82074
R67 VDD1.n2 VDD1.t2 9.82074
R68 VDD1.n1 VDD1.t3 9.82074
R69 VDD1.n1 VDD1.t0 9.82074
R70 VDD1 VDD1.n5 0.519897
R71 VTAIL.n130 VTAIL.n120 756.745
R72 VTAIL.n12 VTAIL.n2 756.745
R73 VTAIL.n28 VTAIL.n18 756.745
R74 VTAIL.n46 VTAIL.n36 756.745
R75 VTAIL.n114 VTAIL.n104 756.745
R76 VTAIL.n96 VTAIL.n86 756.745
R77 VTAIL.n80 VTAIL.n70 756.745
R78 VTAIL.n62 VTAIL.n52 756.745
R79 VTAIL.n124 VTAIL.n123 585
R80 VTAIL.n129 VTAIL.n128 585
R81 VTAIL.n131 VTAIL.n130 585
R82 VTAIL.n6 VTAIL.n5 585
R83 VTAIL.n11 VTAIL.n10 585
R84 VTAIL.n13 VTAIL.n12 585
R85 VTAIL.n22 VTAIL.n21 585
R86 VTAIL.n27 VTAIL.n26 585
R87 VTAIL.n29 VTAIL.n28 585
R88 VTAIL.n40 VTAIL.n39 585
R89 VTAIL.n45 VTAIL.n44 585
R90 VTAIL.n47 VTAIL.n46 585
R91 VTAIL.n115 VTAIL.n114 585
R92 VTAIL.n113 VTAIL.n112 585
R93 VTAIL.n108 VTAIL.n107 585
R94 VTAIL.n97 VTAIL.n96 585
R95 VTAIL.n95 VTAIL.n94 585
R96 VTAIL.n90 VTAIL.n89 585
R97 VTAIL.n81 VTAIL.n80 585
R98 VTAIL.n79 VTAIL.n78 585
R99 VTAIL.n74 VTAIL.n73 585
R100 VTAIL.n63 VTAIL.n62 585
R101 VTAIL.n61 VTAIL.n60 585
R102 VTAIL.n56 VTAIL.n55 585
R103 VTAIL.n125 VTAIL.t7 336.901
R104 VTAIL.n7 VTAIL.t3 336.901
R105 VTAIL.n23 VTAIL.t12 336.901
R106 VTAIL.n41 VTAIL.t9 336.901
R107 VTAIL.n109 VTAIL.t14 336.901
R108 VTAIL.n91 VTAIL.t15 336.901
R109 VTAIL.n75 VTAIL.t4 336.901
R110 VTAIL.n57 VTAIL.t0 336.901
R111 VTAIL.n129 VTAIL.n123 171.744
R112 VTAIL.n130 VTAIL.n129 171.744
R113 VTAIL.n11 VTAIL.n5 171.744
R114 VTAIL.n12 VTAIL.n11 171.744
R115 VTAIL.n27 VTAIL.n21 171.744
R116 VTAIL.n28 VTAIL.n27 171.744
R117 VTAIL.n45 VTAIL.n39 171.744
R118 VTAIL.n46 VTAIL.n45 171.744
R119 VTAIL.n114 VTAIL.n113 171.744
R120 VTAIL.n113 VTAIL.n107 171.744
R121 VTAIL.n96 VTAIL.n95 171.744
R122 VTAIL.n95 VTAIL.n89 171.744
R123 VTAIL.n80 VTAIL.n79 171.744
R124 VTAIL.n79 VTAIL.n73 171.744
R125 VTAIL.n62 VTAIL.n61 171.744
R126 VTAIL.n61 VTAIL.n55 171.744
R127 VTAIL.n103 VTAIL.n102 114.856
R128 VTAIL.n69 VTAIL.n68 114.856
R129 VTAIL.n1 VTAIL.n0 114.856
R130 VTAIL.n35 VTAIL.n34 114.856
R131 VTAIL.t7 VTAIL.n123 85.8723
R132 VTAIL.t3 VTAIL.n5 85.8723
R133 VTAIL.t12 VTAIL.n21 85.8723
R134 VTAIL.t9 VTAIL.n39 85.8723
R135 VTAIL.t14 VTAIL.n107 85.8723
R136 VTAIL.t15 VTAIL.n89 85.8723
R137 VTAIL.t4 VTAIL.n73 85.8723
R138 VTAIL.t0 VTAIL.n55 85.8723
R139 VTAIL.n135 VTAIL.n134 35.8702
R140 VTAIL.n17 VTAIL.n16 35.8702
R141 VTAIL.n33 VTAIL.n32 35.8702
R142 VTAIL.n51 VTAIL.n50 35.8702
R143 VTAIL.n119 VTAIL.n118 35.8702
R144 VTAIL.n101 VTAIL.n100 35.8702
R145 VTAIL.n85 VTAIL.n84 35.8702
R146 VTAIL.n67 VTAIL.n66 35.8702
R147 VTAIL.n135 VTAIL.n119 16.3755
R148 VTAIL.n67 VTAIL.n51 16.3755
R149 VTAIL.n125 VTAIL.n124 16.193
R150 VTAIL.n7 VTAIL.n6 16.193
R151 VTAIL.n23 VTAIL.n22 16.193
R152 VTAIL.n41 VTAIL.n40 16.193
R153 VTAIL.n109 VTAIL.n108 16.193
R154 VTAIL.n91 VTAIL.n90 16.193
R155 VTAIL.n75 VTAIL.n74 16.193
R156 VTAIL.n57 VTAIL.n56 16.193
R157 VTAIL.n128 VTAIL.n127 12.8005
R158 VTAIL.n10 VTAIL.n9 12.8005
R159 VTAIL.n26 VTAIL.n25 12.8005
R160 VTAIL.n44 VTAIL.n43 12.8005
R161 VTAIL.n112 VTAIL.n111 12.8005
R162 VTAIL.n94 VTAIL.n93 12.8005
R163 VTAIL.n78 VTAIL.n77 12.8005
R164 VTAIL.n60 VTAIL.n59 12.8005
R165 VTAIL.n131 VTAIL.n122 12.0247
R166 VTAIL.n13 VTAIL.n4 12.0247
R167 VTAIL.n29 VTAIL.n20 12.0247
R168 VTAIL.n47 VTAIL.n38 12.0247
R169 VTAIL.n115 VTAIL.n106 12.0247
R170 VTAIL.n97 VTAIL.n88 12.0247
R171 VTAIL.n81 VTAIL.n72 12.0247
R172 VTAIL.n63 VTAIL.n54 12.0247
R173 VTAIL.n132 VTAIL.n120 11.249
R174 VTAIL.n14 VTAIL.n2 11.249
R175 VTAIL.n30 VTAIL.n18 11.249
R176 VTAIL.n48 VTAIL.n36 11.249
R177 VTAIL.n116 VTAIL.n104 11.249
R178 VTAIL.n98 VTAIL.n86 11.249
R179 VTAIL.n82 VTAIL.n70 11.249
R180 VTAIL.n64 VTAIL.n52 11.249
R181 VTAIL.n0 VTAIL.t1 9.82074
R182 VTAIL.n0 VTAIL.t2 9.82074
R183 VTAIL.n34 VTAIL.t11 9.82074
R184 VTAIL.n34 VTAIL.t10 9.82074
R185 VTAIL.n102 VTAIL.t13 9.82074
R186 VTAIL.n102 VTAIL.t8 9.82074
R187 VTAIL.n68 VTAIL.t6 9.82074
R188 VTAIL.n68 VTAIL.t5 9.82074
R189 VTAIL.n134 VTAIL.n133 9.45567
R190 VTAIL.n16 VTAIL.n15 9.45567
R191 VTAIL.n32 VTAIL.n31 9.45567
R192 VTAIL.n50 VTAIL.n49 9.45567
R193 VTAIL.n118 VTAIL.n117 9.45567
R194 VTAIL.n100 VTAIL.n99 9.45567
R195 VTAIL.n84 VTAIL.n83 9.45567
R196 VTAIL.n66 VTAIL.n65 9.45567
R197 VTAIL.n133 VTAIL.n132 9.3005
R198 VTAIL.n122 VTAIL.n121 9.3005
R199 VTAIL.n127 VTAIL.n126 9.3005
R200 VTAIL.n15 VTAIL.n14 9.3005
R201 VTAIL.n4 VTAIL.n3 9.3005
R202 VTAIL.n9 VTAIL.n8 9.3005
R203 VTAIL.n31 VTAIL.n30 9.3005
R204 VTAIL.n20 VTAIL.n19 9.3005
R205 VTAIL.n25 VTAIL.n24 9.3005
R206 VTAIL.n49 VTAIL.n48 9.3005
R207 VTAIL.n38 VTAIL.n37 9.3005
R208 VTAIL.n43 VTAIL.n42 9.3005
R209 VTAIL.n117 VTAIL.n116 9.3005
R210 VTAIL.n106 VTAIL.n105 9.3005
R211 VTAIL.n111 VTAIL.n110 9.3005
R212 VTAIL.n99 VTAIL.n98 9.3005
R213 VTAIL.n88 VTAIL.n87 9.3005
R214 VTAIL.n93 VTAIL.n92 9.3005
R215 VTAIL.n83 VTAIL.n82 9.3005
R216 VTAIL.n72 VTAIL.n71 9.3005
R217 VTAIL.n77 VTAIL.n76 9.3005
R218 VTAIL.n65 VTAIL.n64 9.3005
R219 VTAIL.n54 VTAIL.n53 9.3005
R220 VTAIL.n59 VTAIL.n58 9.3005
R221 VTAIL.n110 VTAIL.n109 3.91276
R222 VTAIL.n92 VTAIL.n91 3.91276
R223 VTAIL.n76 VTAIL.n75 3.91276
R224 VTAIL.n58 VTAIL.n57 3.91276
R225 VTAIL.n126 VTAIL.n125 3.91276
R226 VTAIL.n8 VTAIL.n7 3.91276
R227 VTAIL.n24 VTAIL.n23 3.91276
R228 VTAIL.n42 VTAIL.n41 3.91276
R229 VTAIL.n134 VTAIL.n120 2.71565
R230 VTAIL.n16 VTAIL.n2 2.71565
R231 VTAIL.n32 VTAIL.n18 2.71565
R232 VTAIL.n50 VTAIL.n36 2.71565
R233 VTAIL.n118 VTAIL.n104 2.71565
R234 VTAIL.n100 VTAIL.n86 2.71565
R235 VTAIL.n84 VTAIL.n70 2.71565
R236 VTAIL.n66 VTAIL.n52 2.71565
R237 VTAIL.n132 VTAIL.n131 1.93989
R238 VTAIL.n14 VTAIL.n13 1.93989
R239 VTAIL.n30 VTAIL.n29 1.93989
R240 VTAIL.n48 VTAIL.n47 1.93989
R241 VTAIL.n116 VTAIL.n115 1.93989
R242 VTAIL.n98 VTAIL.n97 1.93989
R243 VTAIL.n82 VTAIL.n81 1.93989
R244 VTAIL.n64 VTAIL.n63 1.93989
R245 VTAIL.n128 VTAIL.n122 1.16414
R246 VTAIL.n10 VTAIL.n4 1.16414
R247 VTAIL.n26 VTAIL.n20 1.16414
R248 VTAIL.n44 VTAIL.n38 1.16414
R249 VTAIL.n112 VTAIL.n106 1.16414
R250 VTAIL.n94 VTAIL.n88 1.16414
R251 VTAIL.n78 VTAIL.n72 1.16414
R252 VTAIL.n60 VTAIL.n54 1.16414
R253 VTAIL.n69 VTAIL.n67 1.15567
R254 VTAIL.n85 VTAIL.n69 1.15567
R255 VTAIL.n103 VTAIL.n101 1.15567
R256 VTAIL.n119 VTAIL.n103 1.15567
R257 VTAIL.n51 VTAIL.n35 1.15567
R258 VTAIL.n35 VTAIL.n33 1.15567
R259 VTAIL.n17 VTAIL.n1 1.15567
R260 VTAIL VTAIL.n135 1.09748
R261 VTAIL.n101 VTAIL.n85 0.470328
R262 VTAIL.n33 VTAIL.n17 0.470328
R263 VTAIL.n127 VTAIL.n124 0.388379
R264 VTAIL.n9 VTAIL.n6 0.388379
R265 VTAIL.n25 VTAIL.n22 0.388379
R266 VTAIL.n43 VTAIL.n40 0.388379
R267 VTAIL.n111 VTAIL.n108 0.388379
R268 VTAIL.n93 VTAIL.n90 0.388379
R269 VTAIL.n77 VTAIL.n74 0.388379
R270 VTAIL.n59 VTAIL.n56 0.388379
R271 VTAIL.n126 VTAIL.n121 0.155672
R272 VTAIL.n133 VTAIL.n121 0.155672
R273 VTAIL.n8 VTAIL.n3 0.155672
R274 VTAIL.n15 VTAIL.n3 0.155672
R275 VTAIL.n24 VTAIL.n19 0.155672
R276 VTAIL.n31 VTAIL.n19 0.155672
R277 VTAIL.n42 VTAIL.n37 0.155672
R278 VTAIL.n49 VTAIL.n37 0.155672
R279 VTAIL.n117 VTAIL.n105 0.155672
R280 VTAIL.n110 VTAIL.n105 0.155672
R281 VTAIL.n99 VTAIL.n87 0.155672
R282 VTAIL.n92 VTAIL.n87 0.155672
R283 VTAIL.n83 VTAIL.n71 0.155672
R284 VTAIL.n76 VTAIL.n71 0.155672
R285 VTAIL.n65 VTAIL.n53 0.155672
R286 VTAIL.n58 VTAIL.n53 0.155672
R287 VTAIL VTAIL.n1 0.0586897
R288 VN.n14 VN.n13 161.3
R289 VN.n29 VN.n28 161.3
R290 VN.n27 VN.n15 161.3
R291 VN.n26 VN.n25 161.3
R292 VN.n24 VN.n23 161.3
R293 VN.n22 VN.n17 161.3
R294 VN.n21 VN.n20 161.3
R295 VN.n12 VN.n0 161.3
R296 VN.n11 VN.n10 161.3
R297 VN.n9 VN.n8 161.3
R298 VN.n7 VN.n2 161.3
R299 VN.n6 VN.n5 161.3
R300 VN.n4 VN.t2 133.733
R301 VN.n19 VN.t5 133.733
R302 VN.n13 VN.t3 118.115
R303 VN.n28 VN.t6 118.115
R304 VN.n3 VN.t4 78.9817
R305 VN.n1 VN.t1 78.9817
R306 VN.n18 VN.t7 78.9817
R307 VN.n16 VN.t0 78.9817
R308 VN.n12 VN.n11 56.0336
R309 VN.n27 VN.n26 56.0336
R310 VN.n4 VN.n3 46.6347
R311 VN.n19 VN.n18 46.6347
R312 VN.n20 VN.n19 43.8151
R313 VN.n5 VN.n4 43.8151
R314 VN.n7 VN.n6 40.4934
R315 VN.n8 VN.n7 40.4934
R316 VN.n22 VN.n21 40.4934
R317 VN.n23 VN.n22 40.4934
R318 VN VN.n29 37.2903
R319 VN.n11 VN.n1 16.1487
R320 VN.n26 VN.n16 16.1487
R321 VN.n6 VN.n3 8.31928
R322 VN.n8 VN.n1 8.31928
R323 VN.n21 VN.n18 8.31928
R324 VN.n23 VN.n16 8.31928
R325 VN.n13 VN.n12 0.730803
R326 VN.n28 VN.n27 0.730803
R327 VN.n29 VN.n15 0.189894
R328 VN.n25 VN.n15 0.189894
R329 VN.n25 VN.n24 0.189894
R330 VN.n24 VN.n17 0.189894
R331 VN.n20 VN.n17 0.189894
R332 VN.n5 VN.n2 0.189894
R333 VN.n9 VN.n2 0.189894
R334 VN.n10 VN.n9 0.189894
R335 VN.n10 VN.n0 0.189894
R336 VN.n14 VN.n0 0.189894
R337 VN VN.n14 0.0516364
R338 VDD2.n2 VDD2.n1 132.058
R339 VDD2.n2 VDD2.n0 132.058
R340 VDD2 VDD2.n5 132.054
R341 VDD2.n4 VDD2.n3 131.536
R342 VDD2.n4 VDD2.n2 31.767
R343 VDD2.n5 VDD2.t0 9.82074
R344 VDD2.n5 VDD2.t2 9.82074
R345 VDD2.n3 VDD2.t1 9.82074
R346 VDD2.n3 VDD2.t7 9.82074
R347 VDD2.n1 VDD2.t6 9.82074
R348 VDD2.n1 VDD2.t4 9.82074
R349 VDD2.n0 VDD2.t5 9.82074
R350 VDD2.n0 VDD2.t3 9.82074
R351 VDD2 VDD2.n4 0.636276
R352 B.n300 B.n41 585
R353 B.n302 B.n301 585
R354 B.n303 B.n40 585
R355 B.n305 B.n304 585
R356 B.n306 B.n39 585
R357 B.n308 B.n307 585
R358 B.n309 B.n38 585
R359 B.n311 B.n310 585
R360 B.n312 B.n37 585
R361 B.n314 B.n313 585
R362 B.n315 B.n36 585
R363 B.n317 B.n316 585
R364 B.n318 B.n35 585
R365 B.n320 B.n319 585
R366 B.n321 B.n34 585
R367 B.n323 B.n322 585
R368 B.n325 B.n31 585
R369 B.n327 B.n326 585
R370 B.n328 B.n30 585
R371 B.n330 B.n329 585
R372 B.n331 B.n29 585
R373 B.n333 B.n332 585
R374 B.n334 B.n28 585
R375 B.n336 B.n335 585
R376 B.n337 B.n27 585
R377 B.n339 B.n338 585
R378 B.n341 B.n340 585
R379 B.n342 B.n23 585
R380 B.n344 B.n343 585
R381 B.n345 B.n22 585
R382 B.n347 B.n346 585
R383 B.n348 B.n21 585
R384 B.n350 B.n349 585
R385 B.n351 B.n20 585
R386 B.n353 B.n352 585
R387 B.n354 B.n19 585
R388 B.n356 B.n355 585
R389 B.n357 B.n18 585
R390 B.n359 B.n358 585
R391 B.n360 B.n17 585
R392 B.n362 B.n361 585
R393 B.n363 B.n16 585
R394 B.n299 B.n298 585
R395 B.n297 B.n42 585
R396 B.n296 B.n295 585
R397 B.n294 B.n43 585
R398 B.n293 B.n292 585
R399 B.n291 B.n44 585
R400 B.n290 B.n289 585
R401 B.n288 B.n45 585
R402 B.n287 B.n286 585
R403 B.n285 B.n46 585
R404 B.n284 B.n283 585
R405 B.n282 B.n47 585
R406 B.n281 B.n280 585
R407 B.n279 B.n48 585
R408 B.n278 B.n277 585
R409 B.n276 B.n49 585
R410 B.n275 B.n274 585
R411 B.n273 B.n50 585
R412 B.n272 B.n271 585
R413 B.n270 B.n51 585
R414 B.n269 B.n268 585
R415 B.n267 B.n52 585
R416 B.n266 B.n265 585
R417 B.n264 B.n53 585
R418 B.n263 B.n262 585
R419 B.n261 B.n54 585
R420 B.n260 B.n259 585
R421 B.n258 B.n55 585
R422 B.n257 B.n256 585
R423 B.n255 B.n56 585
R424 B.n254 B.n253 585
R425 B.n252 B.n57 585
R426 B.n251 B.n250 585
R427 B.n249 B.n58 585
R428 B.n248 B.n247 585
R429 B.n246 B.n59 585
R430 B.n245 B.n244 585
R431 B.n243 B.n60 585
R432 B.n242 B.n241 585
R433 B.n240 B.n61 585
R434 B.n239 B.n238 585
R435 B.n237 B.n62 585
R436 B.n236 B.n235 585
R437 B.n234 B.n63 585
R438 B.n233 B.n232 585
R439 B.n231 B.n64 585
R440 B.n230 B.n229 585
R441 B.n228 B.n65 585
R442 B.n227 B.n226 585
R443 B.n225 B.n66 585
R444 B.n224 B.n223 585
R445 B.n222 B.n67 585
R446 B.n221 B.n220 585
R447 B.n219 B.n68 585
R448 B.n218 B.n217 585
R449 B.n216 B.n69 585
R450 B.n215 B.n214 585
R451 B.n150 B.n95 585
R452 B.n152 B.n151 585
R453 B.n153 B.n94 585
R454 B.n155 B.n154 585
R455 B.n156 B.n93 585
R456 B.n158 B.n157 585
R457 B.n159 B.n92 585
R458 B.n161 B.n160 585
R459 B.n162 B.n91 585
R460 B.n164 B.n163 585
R461 B.n165 B.n90 585
R462 B.n167 B.n166 585
R463 B.n168 B.n89 585
R464 B.n170 B.n169 585
R465 B.n171 B.n88 585
R466 B.n173 B.n172 585
R467 B.n175 B.n85 585
R468 B.n177 B.n176 585
R469 B.n178 B.n84 585
R470 B.n180 B.n179 585
R471 B.n181 B.n83 585
R472 B.n183 B.n182 585
R473 B.n184 B.n82 585
R474 B.n186 B.n185 585
R475 B.n187 B.n81 585
R476 B.n189 B.n188 585
R477 B.n191 B.n190 585
R478 B.n192 B.n77 585
R479 B.n194 B.n193 585
R480 B.n195 B.n76 585
R481 B.n197 B.n196 585
R482 B.n198 B.n75 585
R483 B.n200 B.n199 585
R484 B.n201 B.n74 585
R485 B.n203 B.n202 585
R486 B.n204 B.n73 585
R487 B.n206 B.n205 585
R488 B.n207 B.n72 585
R489 B.n209 B.n208 585
R490 B.n210 B.n71 585
R491 B.n212 B.n211 585
R492 B.n213 B.n70 585
R493 B.n149 B.n148 585
R494 B.n147 B.n96 585
R495 B.n146 B.n145 585
R496 B.n144 B.n97 585
R497 B.n143 B.n142 585
R498 B.n141 B.n98 585
R499 B.n140 B.n139 585
R500 B.n138 B.n99 585
R501 B.n137 B.n136 585
R502 B.n135 B.n100 585
R503 B.n134 B.n133 585
R504 B.n132 B.n101 585
R505 B.n131 B.n130 585
R506 B.n129 B.n102 585
R507 B.n128 B.n127 585
R508 B.n126 B.n103 585
R509 B.n125 B.n124 585
R510 B.n123 B.n104 585
R511 B.n122 B.n121 585
R512 B.n120 B.n105 585
R513 B.n119 B.n118 585
R514 B.n117 B.n106 585
R515 B.n116 B.n115 585
R516 B.n114 B.n107 585
R517 B.n113 B.n112 585
R518 B.n111 B.n108 585
R519 B.n110 B.n109 585
R520 B.n2 B.n0 585
R521 B.n405 B.n1 585
R522 B.n404 B.n403 585
R523 B.n402 B.n3 585
R524 B.n401 B.n400 585
R525 B.n399 B.n4 585
R526 B.n398 B.n397 585
R527 B.n396 B.n5 585
R528 B.n395 B.n394 585
R529 B.n393 B.n6 585
R530 B.n392 B.n391 585
R531 B.n390 B.n7 585
R532 B.n389 B.n388 585
R533 B.n387 B.n8 585
R534 B.n386 B.n385 585
R535 B.n384 B.n9 585
R536 B.n383 B.n382 585
R537 B.n381 B.n10 585
R538 B.n380 B.n379 585
R539 B.n378 B.n11 585
R540 B.n377 B.n376 585
R541 B.n375 B.n12 585
R542 B.n374 B.n373 585
R543 B.n372 B.n13 585
R544 B.n371 B.n370 585
R545 B.n369 B.n14 585
R546 B.n368 B.n367 585
R547 B.n366 B.n15 585
R548 B.n365 B.n364 585
R549 B.n407 B.n406 585
R550 B.n148 B.n95 444.452
R551 B.n364 B.n363 444.452
R552 B.n214 B.n213 444.452
R553 B.n298 B.n41 444.452
R554 B.n78 B.t3 281.976
R555 B.n86 B.t0 281.976
R556 B.n24 B.t6 281.976
R557 B.n32 B.t9 281.976
R558 B.n78 B.t5 253.683
R559 B.n32 B.t10 253.683
R560 B.n86 B.t2 253.681
R561 B.n24 B.t7 253.681
R562 B.n79 B.t4 227.695
R563 B.n33 B.t11 227.695
R564 B.n87 B.t1 227.695
R565 B.n25 B.t8 227.695
R566 B.n148 B.n147 163.367
R567 B.n147 B.n146 163.367
R568 B.n146 B.n97 163.367
R569 B.n142 B.n97 163.367
R570 B.n142 B.n141 163.367
R571 B.n141 B.n140 163.367
R572 B.n140 B.n99 163.367
R573 B.n136 B.n99 163.367
R574 B.n136 B.n135 163.367
R575 B.n135 B.n134 163.367
R576 B.n134 B.n101 163.367
R577 B.n130 B.n101 163.367
R578 B.n130 B.n129 163.367
R579 B.n129 B.n128 163.367
R580 B.n128 B.n103 163.367
R581 B.n124 B.n103 163.367
R582 B.n124 B.n123 163.367
R583 B.n123 B.n122 163.367
R584 B.n122 B.n105 163.367
R585 B.n118 B.n105 163.367
R586 B.n118 B.n117 163.367
R587 B.n117 B.n116 163.367
R588 B.n116 B.n107 163.367
R589 B.n112 B.n107 163.367
R590 B.n112 B.n111 163.367
R591 B.n111 B.n110 163.367
R592 B.n110 B.n2 163.367
R593 B.n406 B.n2 163.367
R594 B.n406 B.n405 163.367
R595 B.n405 B.n404 163.367
R596 B.n404 B.n3 163.367
R597 B.n400 B.n3 163.367
R598 B.n400 B.n399 163.367
R599 B.n399 B.n398 163.367
R600 B.n398 B.n5 163.367
R601 B.n394 B.n5 163.367
R602 B.n394 B.n393 163.367
R603 B.n393 B.n392 163.367
R604 B.n392 B.n7 163.367
R605 B.n388 B.n7 163.367
R606 B.n388 B.n387 163.367
R607 B.n387 B.n386 163.367
R608 B.n386 B.n9 163.367
R609 B.n382 B.n9 163.367
R610 B.n382 B.n381 163.367
R611 B.n381 B.n380 163.367
R612 B.n380 B.n11 163.367
R613 B.n376 B.n11 163.367
R614 B.n376 B.n375 163.367
R615 B.n375 B.n374 163.367
R616 B.n374 B.n13 163.367
R617 B.n370 B.n13 163.367
R618 B.n370 B.n369 163.367
R619 B.n369 B.n368 163.367
R620 B.n368 B.n15 163.367
R621 B.n364 B.n15 163.367
R622 B.n152 B.n95 163.367
R623 B.n153 B.n152 163.367
R624 B.n154 B.n153 163.367
R625 B.n154 B.n93 163.367
R626 B.n158 B.n93 163.367
R627 B.n159 B.n158 163.367
R628 B.n160 B.n159 163.367
R629 B.n160 B.n91 163.367
R630 B.n164 B.n91 163.367
R631 B.n165 B.n164 163.367
R632 B.n166 B.n165 163.367
R633 B.n166 B.n89 163.367
R634 B.n170 B.n89 163.367
R635 B.n171 B.n170 163.367
R636 B.n172 B.n171 163.367
R637 B.n172 B.n85 163.367
R638 B.n177 B.n85 163.367
R639 B.n178 B.n177 163.367
R640 B.n179 B.n178 163.367
R641 B.n179 B.n83 163.367
R642 B.n183 B.n83 163.367
R643 B.n184 B.n183 163.367
R644 B.n185 B.n184 163.367
R645 B.n185 B.n81 163.367
R646 B.n189 B.n81 163.367
R647 B.n190 B.n189 163.367
R648 B.n190 B.n77 163.367
R649 B.n194 B.n77 163.367
R650 B.n195 B.n194 163.367
R651 B.n196 B.n195 163.367
R652 B.n196 B.n75 163.367
R653 B.n200 B.n75 163.367
R654 B.n201 B.n200 163.367
R655 B.n202 B.n201 163.367
R656 B.n202 B.n73 163.367
R657 B.n206 B.n73 163.367
R658 B.n207 B.n206 163.367
R659 B.n208 B.n207 163.367
R660 B.n208 B.n71 163.367
R661 B.n212 B.n71 163.367
R662 B.n213 B.n212 163.367
R663 B.n214 B.n69 163.367
R664 B.n218 B.n69 163.367
R665 B.n219 B.n218 163.367
R666 B.n220 B.n219 163.367
R667 B.n220 B.n67 163.367
R668 B.n224 B.n67 163.367
R669 B.n225 B.n224 163.367
R670 B.n226 B.n225 163.367
R671 B.n226 B.n65 163.367
R672 B.n230 B.n65 163.367
R673 B.n231 B.n230 163.367
R674 B.n232 B.n231 163.367
R675 B.n232 B.n63 163.367
R676 B.n236 B.n63 163.367
R677 B.n237 B.n236 163.367
R678 B.n238 B.n237 163.367
R679 B.n238 B.n61 163.367
R680 B.n242 B.n61 163.367
R681 B.n243 B.n242 163.367
R682 B.n244 B.n243 163.367
R683 B.n244 B.n59 163.367
R684 B.n248 B.n59 163.367
R685 B.n249 B.n248 163.367
R686 B.n250 B.n249 163.367
R687 B.n250 B.n57 163.367
R688 B.n254 B.n57 163.367
R689 B.n255 B.n254 163.367
R690 B.n256 B.n255 163.367
R691 B.n256 B.n55 163.367
R692 B.n260 B.n55 163.367
R693 B.n261 B.n260 163.367
R694 B.n262 B.n261 163.367
R695 B.n262 B.n53 163.367
R696 B.n266 B.n53 163.367
R697 B.n267 B.n266 163.367
R698 B.n268 B.n267 163.367
R699 B.n268 B.n51 163.367
R700 B.n272 B.n51 163.367
R701 B.n273 B.n272 163.367
R702 B.n274 B.n273 163.367
R703 B.n274 B.n49 163.367
R704 B.n278 B.n49 163.367
R705 B.n279 B.n278 163.367
R706 B.n280 B.n279 163.367
R707 B.n280 B.n47 163.367
R708 B.n284 B.n47 163.367
R709 B.n285 B.n284 163.367
R710 B.n286 B.n285 163.367
R711 B.n286 B.n45 163.367
R712 B.n290 B.n45 163.367
R713 B.n291 B.n290 163.367
R714 B.n292 B.n291 163.367
R715 B.n292 B.n43 163.367
R716 B.n296 B.n43 163.367
R717 B.n297 B.n296 163.367
R718 B.n298 B.n297 163.367
R719 B.n363 B.n362 163.367
R720 B.n362 B.n17 163.367
R721 B.n358 B.n17 163.367
R722 B.n358 B.n357 163.367
R723 B.n357 B.n356 163.367
R724 B.n356 B.n19 163.367
R725 B.n352 B.n19 163.367
R726 B.n352 B.n351 163.367
R727 B.n351 B.n350 163.367
R728 B.n350 B.n21 163.367
R729 B.n346 B.n21 163.367
R730 B.n346 B.n345 163.367
R731 B.n345 B.n344 163.367
R732 B.n344 B.n23 163.367
R733 B.n340 B.n23 163.367
R734 B.n340 B.n339 163.367
R735 B.n339 B.n27 163.367
R736 B.n335 B.n27 163.367
R737 B.n335 B.n334 163.367
R738 B.n334 B.n333 163.367
R739 B.n333 B.n29 163.367
R740 B.n329 B.n29 163.367
R741 B.n329 B.n328 163.367
R742 B.n328 B.n327 163.367
R743 B.n327 B.n31 163.367
R744 B.n322 B.n31 163.367
R745 B.n322 B.n321 163.367
R746 B.n321 B.n320 163.367
R747 B.n320 B.n35 163.367
R748 B.n316 B.n35 163.367
R749 B.n316 B.n315 163.367
R750 B.n315 B.n314 163.367
R751 B.n314 B.n37 163.367
R752 B.n310 B.n37 163.367
R753 B.n310 B.n309 163.367
R754 B.n309 B.n308 163.367
R755 B.n308 B.n39 163.367
R756 B.n304 B.n39 163.367
R757 B.n304 B.n303 163.367
R758 B.n303 B.n302 163.367
R759 B.n302 B.n41 163.367
R760 B.n80 B.n79 59.5399
R761 B.n174 B.n87 59.5399
R762 B.n26 B.n25 59.5399
R763 B.n324 B.n33 59.5399
R764 B.n365 B.n16 28.8785
R765 B.n215 B.n70 28.8785
R766 B.n150 B.n149 28.8785
R767 B.n300 B.n299 28.8785
R768 B.n79 B.n78 25.9884
R769 B.n87 B.n86 25.9884
R770 B.n25 B.n24 25.9884
R771 B.n33 B.n32 25.9884
R772 B B.n407 18.0485
R773 B.n361 B.n16 10.6151
R774 B.n361 B.n360 10.6151
R775 B.n360 B.n359 10.6151
R776 B.n359 B.n18 10.6151
R777 B.n355 B.n18 10.6151
R778 B.n355 B.n354 10.6151
R779 B.n354 B.n353 10.6151
R780 B.n353 B.n20 10.6151
R781 B.n349 B.n20 10.6151
R782 B.n349 B.n348 10.6151
R783 B.n348 B.n347 10.6151
R784 B.n347 B.n22 10.6151
R785 B.n343 B.n22 10.6151
R786 B.n343 B.n342 10.6151
R787 B.n342 B.n341 10.6151
R788 B.n338 B.n337 10.6151
R789 B.n337 B.n336 10.6151
R790 B.n336 B.n28 10.6151
R791 B.n332 B.n28 10.6151
R792 B.n332 B.n331 10.6151
R793 B.n331 B.n330 10.6151
R794 B.n330 B.n30 10.6151
R795 B.n326 B.n30 10.6151
R796 B.n326 B.n325 10.6151
R797 B.n323 B.n34 10.6151
R798 B.n319 B.n34 10.6151
R799 B.n319 B.n318 10.6151
R800 B.n318 B.n317 10.6151
R801 B.n317 B.n36 10.6151
R802 B.n313 B.n36 10.6151
R803 B.n313 B.n312 10.6151
R804 B.n312 B.n311 10.6151
R805 B.n311 B.n38 10.6151
R806 B.n307 B.n38 10.6151
R807 B.n307 B.n306 10.6151
R808 B.n306 B.n305 10.6151
R809 B.n305 B.n40 10.6151
R810 B.n301 B.n40 10.6151
R811 B.n301 B.n300 10.6151
R812 B.n216 B.n215 10.6151
R813 B.n217 B.n216 10.6151
R814 B.n217 B.n68 10.6151
R815 B.n221 B.n68 10.6151
R816 B.n222 B.n221 10.6151
R817 B.n223 B.n222 10.6151
R818 B.n223 B.n66 10.6151
R819 B.n227 B.n66 10.6151
R820 B.n228 B.n227 10.6151
R821 B.n229 B.n228 10.6151
R822 B.n229 B.n64 10.6151
R823 B.n233 B.n64 10.6151
R824 B.n234 B.n233 10.6151
R825 B.n235 B.n234 10.6151
R826 B.n235 B.n62 10.6151
R827 B.n239 B.n62 10.6151
R828 B.n240 B.n239 10.6151
R829 B.n241 B.n240 10.6151
R830 B.n241 B.n60 10.6151
R831 B.n245 B.n60 10.6151
R832 B.n246 B.n245 10.6151
R833 B.n247 B.n246 10.6151
R834 B.n247 B.n58 10.6151
R835 B.n251 B.n58 10.6151
R836 B.n252 B.n251 10.6151
R837 B.n253 B.n252 10.6151
R838 B.n253 B.n56 10.6151
R839 B.n257 B.n56 10.6151
R840 B.n258 B.n257 10.6151
R841 B.n259 B.n258 10.6151
R842 B.n259 B.n54 10.6151
R843 B.n263 B.n54 10.6151
R844 B.n264 B.n263 10.6151
R845 B.n265 B.n264 10.6151
R846 B.n265 B.n52 10.6151
R847 B.n269 B.n52 10.6151
R848 B.n270 B.n269 10.6151
R849 B.n271 B.n270 10.6151
R850 B.n271 B.n50 10.6151
R851 B.n275 B.n50 10.6151
R852 B.n276 B.n275 10.6151
R853 B.n277 B.n276 10.6151
R854 B.n277 B.n48 10.6151
R855 B.n281 B.n48 10.6151
R856 B.n282 B.n281 10.6151
R857 B.n283 B.n282 10.6151
R858 B.n283 B.n46 10.6151
R859 B.n287 B.n46 10.6151
R860 B.n288 B.n287 10.6151
R861 B.n289 B.n288 10.6151
R862 B.n289 B.n44 10.6151
R863 B.n293 B.n44 10.6151
R864 B.n294 B.n293 10.6151
R865 B.n295 B.n294 10.6151
R866 B.n295 B.n42 10.6151
R867 B.n299 B.n42 10.6151
R868 B.n151 B.n150 10.6151
R869 B.n151 B.n94 10.6151
R870 B.n155 B.n94 10.6151
R871 B.n156 B.n155 10.6151
R872 B.n157 B.n156 10.6151
R873 B.n157 B.n92 10.6151
R874 B.n161 B.n92 10.6151
R875 B.n162 B.n161 10.6151
R876 B.n163 B.n162 10.6151
R877 B.n163 B.n90 10.6151
R878 B.n167 B.n90 10.6151
R879 B.n168 B.n167 10.6151
R880 B.n169 B.n168 10.6151
R881 B.n169 B.n88 10.6151
R882 B.n173 B.n88 10.6151
R883 B.n176 B.n175 10.6151
R884 B.n176 B.n84 10.6151
R885 B.n180 B.n84 10.6151
R886 B.n181 B.n180 10.6151
R887 B.n182 B.n181 10.6151
R888 B.n182 B.n82 10.6151
R889 B.n186 B.n82 10.6151
R890 B.n187 B.n186 10.6151
R891 B.n188 B.n187 10.6151
R892 B.n192 B.n191 10.6151
R893 B.n193 B.n192 10.6151
R894 B.n193 B.n76 10.6151
R895 B.n197 B.n76 10.6151
R896 B.n198 B.n197 10.6151
R897 B.n199 B.n198 10.6151
R898 B.n199 B.n74 10.6151
R899 B.n203 B.n74 10.6151
R900 B.n204 B.n203 10.6151
R901 B.n205 B.n204 10.6151
R902 B.n205 B.n72 10.6151
R903 B.n209 B.n72 10.6151
R904 B.n210 B.n209 10.6151
R905 B.n211 B.n210 10.6151
R906 B.n211 B.n70 10.6151
R907 B.n149 B.n96 10.6151
R908 B.n145 B.n96 10.6151
R909 B.n145 B.n144 10.6151
R910 B.n144 B.n143 10.6151
R911 B.n143 B.n98 10.6151
R912 B.n139 B.n98 10.6151
R913 B.n139 B.n138 10.6151
R914 B.n138 B.n137 10.6151
R915 B.n137 B.n100 10.6151
R916 B.n133 B.n100 10.6151
R917 B.n133 B.n132 10.6151
R918 B.n132 B.n131 10.6151
R919 B.n131 B.n102 10.6151
R920 B.n127 B.n102 10.6151
R921 B.n127 B.n126 10.6151
R922 B.n126 B.n125 10.6151
R923 B.n125 B.n104 10.6151
R924 B.n121 B.n104 10.6151
R925 B.n121 B.n120 10.6151
R926 B.n120 B.n119 10.6151
R927 B.n119 B.n106 10.6151
R928 B.n115 B.n106 10.6151
R929 B.n115 B.n114 10.6151
R930 B.n114 B.n113 10.6151
R931 B.n113 B.n108 10.6151
R932 B.n109 B.n108 10.6151
R933 B.n109 B.n0 10.6151
R934 B.n403 B.n1 10.6151
R935 B.n403 B.n402 10.6151
R936 B.n402 B.n401 10.6151
R937 B.n401 B.n4 10.6151
R938 B.n397 B.n4 10.6151
R939 B.n397 B.n396 10.6151
R940 B.n396 B.n395 10.6151
R941 B.n395 B.n6 10.6151
R942 B.n391 B.n6 10.6151
R943 B.n391 B.n390 10.6151
R944 B.n390 B.n389 10.6151
R945 B.n389 B.n8 10.6151
R946 B.n385 B.n8 10.6151
R947 B.n385 B.n384 10.6151
R948 B.n384 B.n383 10.6151
R949 B.n383 B.n10 10.6151
R950 B.n379 B.n10 10.6151
R951 B.n379 B.n378 10.6151
R952 B.n378 B.n377 10.6151
R953 B.n377 B.n12 10.6151
R954 B.n373 B.n12 10.6151
R955 B.n373 B.n372 10.6151
R956 B.n372 B.n371 10.6151
R957 B.n371 B.n14 10.6151
R958 B.n367 B.n14 10.6151
R959 B.n367 B.n366 10.6151
R960 B.n366 B.n365 10.6151
R961 B.n341 B.n26 9.36635
R962 B.n324 B.n323 9.36635
R963 B.n174 B.n173 9.36635
R964 B.n191 B.n80 9.36635
R965 B.n407 B.n0 2.81026
R966 B.n407 B.n1 2.81026
R967 B.n338 B.n26 1.24928
R968 B.n325 B.n324 1.24928
R969 B.n175 B.n174 1.24928
R970 B.n188 B.n80 1.24928
C0 VDD2 B 0.976247f
C1 B VN 0.754656f
C2 VTAIL VDD2 4.4288f
C3 VTAIL VN 2.42762f
C4 VDD2 w_n2310_n1630# 1.23007f
C5 VN w_n2310_n1630# 4.07826f
C6 VP VDD1 2.29302f
C7 B VDD1 0.929892f
C8 B VP 1.24069f
C9 VTAIL VDD1 4.38504f
C10 VTAIL VP 2.44173f
C11 VDD2 VN 2.09203f
C12 VDD1 w_n2310_n1630# 1.18276f
C13 VP w_n2310_n1630# 4.37162f
C14 VTAIL B 1.58799f
C15 B w_n2310_n1630# 5.2475f
C16 VTAIL w_n2310_n1630# 2.0146f
C17 VDD2 VDD1 0.980981f
C18 VDD1 VN 0.153604f
C19 VDD2 VP 0.355736f
C20 VP VN 4.11235f
C21 VDD2 VSUBS 1.01688f
C22 VDD1 VSUBS 1.3856f
C23 VTAIL VSUBS 0.444132f
C24 VN VSUBS 4.44179f
C25 VP VSUBS 1.507008f
C26 B VSUBS 2.373058f
C27 w_n2310_n1630# VSUBS 47.5952f
C28 B.n0 VSUBS 0.004795f
C29 B.n1 VSUBS 0.004795f
C30 B.n2 VSUBS 0.007583f
C31 B.n3 VSUBS 0.007583f
C32 B.n4 VSUBS 0.007583f
C33 B.n5 VSUBS 0.007583f
C34 B.n6 VSUBS 0.007583f
C35 B.n7 VSUBS 0.007583f
C36 B.n8 VSUBS 0.007583f
C37 B.n9 VSUBS 0.007583f
C38 B.n10 VSUBS 0.007583f
C39 B.n11 VSUBS 0.007583f
C40 B.n12 VSUBS 0.007583f
C41 B.n13 VSUBS 0.007583f
C42 B.n14 VSUBS 0.007583f
C43 B.n15 VSUBS 0.007583f
C44 B.n16 VSUBS 0.01685f
C45 B.n17 VSUBS 0.007583f
C46 B.n18 VSUBS 0.007583f
C47 B.n19 VSUBS 0.007583f
C48 B.n20 VSUBS 0.007583f
C49 B.n21 VSUBS 0.007583f
C50 B.n22 VSUBS 0.007583f
C51 B.n23 VSUBS 0.007583f
C52 B.t8 VSUBS 0.05307f
C53 B.t7 VSUBS 0.062294f
C54 B.t6 VSUBS 0.168352f
C55 B.n24 VSUBS 0.112274f
C56 B.n25 VSUBS 0.100853f
C57 B.n26 VSUBS 0.017569f
C58 B.n27 VSUBS 0.007583f
C59 B.n28 VSUBS 0.007583f
C60 B.n29 VSUBS 0.007583f
C61 B.n30 VSUBS 0.007583f
C62 B.n31 VSUBS 0.007583f
C63 B.t11 VSUBS 0.053071f
C64 B.t10 VSUBS 0.062294f
C65 B.t9 VSUBS 0.168352f
C66 B.n32 VSUBS 0.112274f
C67 B.n33 VSUBS 0.100853f
C68 B.n34 VSUBS 0.007583f
C69 B.n35 VSUBS 0.007583f
C70 B.n36 VSUBS 0.007583f
C71 B.n37 VSUBS 0.007583f
C72 B.n38 VSUBS 0.007583f
C73 B.n39 VSUBS 0.007583f
C74 B.n40 VSUBS 0.007583f
C75 B.n41 VSUBS 0.01685f
C76 B.n42 VSUBS 0.007583f
C77 B.n43 VSUBS 0.007583f
C78 B.n44 VSUBS 0.007583f
C79 B.n45 VSUBS 0.007583f
C80 B.n46 VSUBS 0.007583f
C81 B.n47 VSUBS 0.007583f
C82 B.n48 VSUBS 0.007583f
C83 B.n49 VSUBS 0.007583f
C84 B.n50 VSUBS 0.007583f
C85 B.n51 VSUBS 0.007583f
C86 B.n52 VSUBS 0.007583f
C87 B.n53 VSUBS 0.007583f
C88 B.n54 VSUBS 0.007583f
C89 B.n55 VSUBS 0.007583f
C90 B.n56 VSUBS 0.007583f
C91 B.n57 VSUBS 0.007583f
C92 B.n58 VSUBS 0.007583f
C93 B.n59 VSUBS 0.007583f
C94 B.n60 VSUBS 0.007583f
C95 B.n61 VSUBS 0.007583f
C96 B.n62 VSUBS 0.007583f
C97 B.n63 VSUBS 0.007583f
C98 B.n64 VSUBS 0.007583f
C99 B.n65 VSUBS 0.007583f
C100 B.n66 VSUBS 0.007583f
C101 B.n67 VSUBS 0.007583f
C102 B.n68 VSUBS 0.007583f
C103 B.n69 VSUBS 0.007583f
C104 B.n70 VSUBS 0.01685f
C105 B.n71 VSUBS 0.007583f
C106 B.n72 VSUBS 0.007583f
C107 B.n73 VSUBS 0.007583f
C108 B.n74 VSUBS 0.007583f
C109 B.n75 VSUBS 0.007583f
C110 B.n76 VSUBS 0.007583f
C111 B.n77 VSUBS 0.007583f
C112 B.t4 VSUBS 0.053071f
C113 B.t5 VSUBS 0.062294f
C114 B.t3 VSUBS 0.168352f
C115 B.n78 VSUBS 0.112274f
C116 B.n79 VSUBS 0.100853f
C117 B.n80 VSUBS 0.017569f
C118 B.n81 VSUBS 0.007583f
C119 B.n82 VSUBS 0.007583f
C120 B.n83 VSUBS 0.007583f
C121 B.n84 VSUBS 0.007583f
C122 B.n85 VSUBS 0.007583f
C123 B.t1 VSUBS 0.05307f
C124 B.t2 VSUBS 0.062294f
C125 B.t0 VSUBS 0.168352f
C126 B.n86 VSUBS 0.112274f
C127 B.n87 VSUBS 0.100853f
C128 B.n88 VSUBS 0.007583f
C129 B.n89 VSUBS 0.007583f
C130 B.n90 VSUBS 0.007583f
C131 B.n91 VSUBS 0.007583f
C132 B.n92 VSUBS 0.007583f
C133 B.n93 VSUBS 0.007583f
C134 B.n94 VSUBS 0.007583f
C135 B.n95 VSUBS 0.01685f
C136 B.n96 VSUBS 0.007583f
C137 B.n97 VSUBS 0.007583f
C138 B.n98 VSUBS 0.007583f
C139 B.n99 VSUBS 0.007583f
C140 B.n100 VSUBS 0.007583f
C141 B.n101 VSUBS 0.007583f
C142 B.n102 VSUBS 0.007583f
C143 B.n103 VSUBS 0.007583f
C144 B.n104 VSUBS 0.007583f
C145 B.n105 VSUBS 0.007583f
C146 B.n106 VSUBS 0.007583f
C147 B.n107 VSUBS 0.007583f
C148 B.n108 VSUBS 0.007583f
C149 B.n109 VSUBS 0.007583f
C150 B.n110 VSUBS 0.007583f
C151 B.n111 VSUBS 0.007583f
C152 B.n112 VSUBS 0.007583f
C153 B.n113 VSUBS 0.007583f
C154 B.n114 VSUBS 0.007583f
C155 B.n115 VSUBS 0.007583f
C156 B.n116 VSUBS 0.007583f
C157 B.n117 VSUBS 0.007583f
C158 B.n118 VSUBS 0.007583f
C159 B.n119 VSUBS 0.007583f
C160 B.n120 VSUBS 0.007583f
C161 B.n121 VSUBS 0.007583f
C162 B.n122 VSUBS 0.007583f
C163 B.n123 VSUBS 0.007583f
C164 B.n124 VSUBS 0.007583f
C165 B.n125 VSUBS 0.007583f
C166 B.n126 VSUBS 0.007583f
C167 B.n127 VSUBS 0.007583f
C168 B.n128 VSUBS 0.007583f
C169 B.n129 VSUBS 0.007583f
C170 B.n130 VSUBS 0.007583f
C171 B.n131 VSUBS 0.007583f
C172 B.n132 VSUBS 0.007583f
C173 B.n133 VSUBS 0.007583f
C174 B.n134 VSUBS 0.007583f
C175 B.n135 VSUBS 0.007583f
C176 B.n136 VSUBS 0.007583f
C177 B.n137 VSUBS 0.007583f
C178 B.n138 VSUBS 0.007583f
C179 B.n139 VSUBS 0.007583f
C180 B.n140 VSUBS 0.007583f
C181 B.n141 VSUBS 0.007583f
C182 B.n142 VSUBS 0.007583f
C183 B.n143 VSUBS 0.007583f
C184 B.n144 VSUBS 0.007583f
C185 B.n145 VSUBS 0.007583f
C186 B.n146 VSUBS 0.007583f
C187 B.n147 VSUBS 0.007583f
C188 B.n148 VSUBS 0.015936f
C189 B.n149 VSUBS 0.015936f
C190 B.n150 VSUBS 0.01685f
C191 B.n151 VSUBS 0.007583f
C192 B.n152 VSUBS 0.007583f
C193 B.n153 VSUBS 0.007583f
C194 B.n154 VSUBS 0.007583f
C195 B.n155 VSUBS 0.007583f
C196 B.n156 VSUBS 0.007583f
C197 B.n157 VSUBS 0.007583f
C198 B.n158 VSUBS 0.007583f
C199 B.n159 VSUBS 0.007583f
C200 B.n160 VSUBS 0.007583f
C201 B.n161 VSUBS 0.007583f
C202 B.n162 VSUBS 0.007583f
C203 B.n163 VSUBS 0.007583f
C204 B.n164 VSUBS 0.007583f
C205 B.n165 VSUBS 0.007583f
C206 B.n166 VSUBS 0.007583f
C207 B.n167 VSUBS 0.007583f
C208 B.n168 VSUBS 0.007583f
C209 B.n169 VSUBS 0.007583f
C210 B.n170 VSUBS 0.007583f
C211 B.n171 VSUBS 0.007583f
C212 B.n172 VSUBS 0.007583f
C213 B.n173 VSUBS 0.007137f
C214 B.n174 VSUBS 0.017569f
C215 B.n175 VSUBS 0.004238f
C216 B.n176 VSUBS 0.007583f
C217 B.n177 VSUBS 0.007583f
C218 B.n178 VSUBS 0.007583f
C219 B.n179 VSUBS 0.007583f
C220 B.n180 VSUBS 0.007583f
C221 B.n181 VSUBS 0.007583f
C222 B.n182 VSUBS 0.007583f
C223 B.n183 VSUBS 0.007583f
C224 B.n184 VSUBS 0.007583f
C225 B.n185 VSUBS 0.007583f
C226 B.n186 VSUBS 0.007583f
C227 B.n187 VSUBS 0.007583f
C228 B.n188 VSUBS 0.004238f
C229 B.n189 VSUBS 0.007583f
C230 B.n190 VSUBS 0.007583f
C231 B.n191 VSUBS 0.007137f
C232 B.n192 VSUBS 0.007583f
C233 B.n193 VSUBS 0.007583f
C234 B.n194 VSUBS 0.007583f
C235 B.n195 VSUBS 0.007583f
C236 B.n196 VSUBS 0.007583f
C237 B.n197 VSUBS 0.007583f
C238 B.n198 VSUBS 0.007583f
C239 B.n199 VSUBS 0.007583f
C240 B.n200 VSUBS 0.007583f
C241 B.n201 VSUBS 0.007583f
C242 B.n202 VSUBS 0.007583f
C243 B.n203 VSUBS 0.007583f
C244 B.n204 VSUBS 0.007583f
C245 B.n205 VSUBS 0.007583f
C246 B.n206 VSUBS 0.007583f
C247 B.n207 VSUBS 0.007583f
C248 B.n208 VSUBS 0.007583f
C249 B.n209 VSUBS 0.007583f
C250 B.n210 VSUBS 0.007583f
C251 B.n211 VSUBS 0.007583f
C252 B.n212 VSUBS 0.007583f
C253 B.n213 VSUBS 0.01685f
C254 B.n214 VSUBS 0.015936f
C255 B.n215 VSUBS 0.015936f
C256 B.n216 VSUBS 0.007583f
C257 B.n217 VSUBS 0.007583f
C258 B.n218 VSUBS 0.007583f
C259 B.n219 VSUBS 0.007583f
C260 B.n220 VSUBS 0.007583f
C261 B.n221 VSUBS 0.007583f
C262 B.n222 VSUBS 0.007583f
C263 B.n223 VSUBS 0.007583f
C264 B.n224 VSUBS 0.007583f
C265 B.n225 VSUBS 0.007583f
C266 B.n226 VSUBS 0.007583f
C267 B.n227 VSUBS 0.007583f
C268 B.n228 VSUBS 0.007583f
C269 B.n229 VSUBS 0.007583f
C270 B.n230 VSUBS 0.007583f
C271 B.n231 VSUBS 0.007583f
C272 B.n232 VSUBS 0.007583f
C273 B.n233 VSUBS 0.007583f
C274 B.n234 VSUBS 0.007583f
C275 B.n235 VSUBS 0.007583f
C276 B.n236 VSUBS 0.007583f
C277 B.n237 VSUBS 0.007583f
C278 B.n238 VSUBS 0.007583f
C279 B.n239 VSUBS 0.007583f
C280 B.n240 VSUBS 0.007583f
C281 B.n241 VSUBS 0.007583f
C282 B.n242 VSUBS 0.007583f
C283 B.n243 VSUBS 0.007583f
C284 B.n244 VSUBS 0.007583f
C285 B.n245 VSUBS 0.007583f
C286 B.n246 VSUBS 0.007583f
C287 B.n247 VSUBS 0.007583f
C288 B.n248 VSUBS 0.007583f
C289 B.n249 VSUBS 0.007583f
C290 B.n250 VSUBS 0.007583f
C291 B.n251 VSUBS 0.007583f
C292 B.n252 VSUBS 0.007583f
C293 B.n253 VSUBS 0.007583f
C294 B.n254 VSUBS 0.007583f
C295 B.n255 VSUBS 0.007583f
C296 B.n256 VSUBS 0.007583f
C297 B.n257 VSUBS 0.007583f
C298 B.n258 VSUBS 0.007583f
C299 B.n259 VSUBS 0.007583f
C300 B.n260 VSUBS 0.007583f
C301 B.n261 VSUBS 0.007583f
C302 B.n262 VSUBS 0.007583f
C303 B.n263 VSUBS 0.007583f
C304 B.n264 VSUBS 0.007583f
C305 B.n265 VSUBS 0.007583f
C306 B.n266 VSUBS 0.007583f
C307 B.n267 VSUBS 0.007583f
C308 B.n268 VSUBS 0.007583f
C309 B.n269 VSUBS 0.007583f
C310 B.n270 VSUBS 0.007583f
C311 B.n271 VSUBS 0.007583f
C312 B.n272 VSUBS 0.007583f
C313 B.n273 VSUBS 0.007583f
C314 B.n274 VSUBS 0.007583f
C315 B.n275 VSUBS 0.007583f
C316 B.n276 VSUBS 0.007583f
C317 B.n277 VSUBS 0.007583f
C318 B.n278 VSUBS 0.007583f
C319 B.n279 VSUBS 0.007583f
C320 B.n280 VSUBS 0.007583f
C321 B.n281 VSUBS 0.007583f
C322 B.n282 VSUBS 0.007583f
C323 B.n283 VSUBS 0.007583f
C324 B.n284 VSUBS 0.007583f
C325 B.n285 VSUBS 0.007583f
C326 B.n286 VSUBS 0.007583f
C327 B.n287 VSUBS 0.007583f
C328 B.n288 VSUBS 0.007583f
C329 B.n289 VSUBS 0.007583f
C330 B.n290 VSUBS 0.007583f
C331 B.n291 VSUBS 0.007583f
C332 B.n292 VSUBS 0.007583f
C333 B.n293 VSUBS 0.007583f
C334 B.n294 VSUBS 0.007583f
C335 B.n295 VSUBS 0.007583f
C336 B.n296 VSUBS 0.007583f
C337 B.n297 VSUBS 0.007583f
C338 B.n298 VSUBS 0.015936f
C339 B.n299 VSUBS 0.016949f
C340 B.n300 VSUBS 0.015837f
C341 B.n301 VSUBS 0.007583f
C342 B.n302 VSUBS 0.007583f
C343 B.n303 VSUBS 0.007583f
C344 B.n304 VSUBS 0.007583f
C345 B.n305 VSUBS 0.007583f
C346 B.n306 VSUBS 0.007583f
C347 B.n307 VSUBS 0.007583f
C348 B.n308 VSUBS 0.007583f
C349 B.n309 VSUBS 0.007583f
C350 B.n310 VSUBS 0.007583f
C351 B.n311 VSUBS 0.007583f
C352 B.n312 VSUBS 0.007583f
C353 B.n313 VSUBS 0.007583f
C354 B.n314 VSUBS 0.007583f
C355 B.n315 VSUBS 0.007583f
C356 B.n316 VSUBS 0.007583f
C357 B.n317 VSUBS 0.007583f
C358 B.n318 VSUBS 0.007583f
C359 B.n319 VSUBS 0.007583f
C360 B.n320 VSUBS 0.007583f
C361 B.n321 VSUBS 0.007583f
C362 B.n322 VSUBS 0.007583f
C363 B.n323 VSUBS 0.007137f
C364 B.n324 VSUBS 0.017569f
C365 B.n325 VSUBS 0.004238f
C366 B.n326 VSUBS 0.007583f
C367 B.n327 VSUBS 0.007583f
C368 B.n328 VSUBS 0.007583f
C369 B.n329 VSUBS 0.007583f
C370 B.n330 VSUBS 0.007583f
C371 B.n331 VSUBS 0.007583f
C372 B.n332 VSUBS 0.007583f
C373 B.n333 VSUBS 0.007583f
C374 B.n334 VSUBS 0.007583f
C375 B.n335 VSUBS 0.007583f
C376 B.n336 VSUBS 0.007583f
C377 B.n337 VSUBS 0.007583f
C378 B.n338 VSUBS 0.004238f
C379 B.n339 VSUBS 0.007583f
C380 B.n340 VSUBS 0.007583f
C381 B.n341 VSUBS 0.007137f
C382 B.n342 VSUBS 0.007583f
C383 B.n343 VSUBS 0.007583f
C384 B.n344 VSUBS 0.007583f
C385 B.n345 VSUBS 0.007583f
C386 B.n346 VSUBS 0.007583f
C387 B.n347 VSUBS 0.007583f
C388 B.n348 VSUBS 0.007583f
C389 B.n349 VSUBS 0.007583f
C390 B.n350 VSUBS 0.007583f
C391 B.n351 VSUBS 0.007583f
C392 B.n352 VSUBS 0.007583f
C393 B.n353 VSUBS 0.007583f
C394 B.n354 VSUBS 0.007583f
C395 B.n355 VSUBS 0.007583f
C396 B.n356 VSUBS 0.007583f
C397 B.n357 VSUBS 0.007583f
C398 B.n358 VSUBS 0.007583f
C399 B.n359 VSUBS 0.007583f
C400 B.n360 VSUBS 0.007583f
C401 B.n361 VSUBS 0.007583f
C402 B.n362 VSUBS 0.007583f
C403 B.n363 VSUBS 0.01685f
C404 B.n364 VSUBS 0.015936f
C405 B.n365 VSUBS 0.015936f
C406 B.n366 VSUBS 0.007583f
C407 B.n367 VSUBS 0.007583f
C408 B.n368 VSUBS 0.007583f
C409 B.n369 VSUBS 0.007583f
C410 B.n370 VSUBS 0.007583f
C411 B.n371 VSUBS 0.007583f
C412 B.n372 VSUBS 0.007583f
C413 B.n373 VSUBS 0.007583f
C414 B.n374 VSUBS 0.007583f
C415 B.n375 VSUBS 0.007583f
C416 B.n376 VSUBS 0.007583f
C417 B.n377 VSUBS 0.007583f
C418 B.n378 VSUBS 0.007583f
C419 B.n379 VSUBS 0.007583f
C420 B.n380 VSUBS 0.007583f
C421 B.n381 VSUBS 0.007583f
C422 B.n382 VSUBS 0.007583f
C423 B.n383 VSUBS 0.007583f
C424 B.n384 VSUBS 0.007583f
C425 B.n385 VSUBS 0.007583f
C426 B.n386 VSUBS 0.007583f
C427 B.n387 VSUBS 0.007583f
C428 B.n388 VSUBS 0.007583f
C429 B.n389 VSUBS 0.007583f
C430 B.n390 VSUBS 0.007583f
C431 B.n391 VSUBS 0.007583f
C432 B.n392 VSUBS 0.007583f
C433 B.n393 VSUBS 0.007583f
C434 B.n394 VSUBS 0.007583f
C435 B.n395 VSUBS 0.007583f
C436 B.n396 VSUBS 0.007583f
C437 B.n397 VSUBS 0.007583f
C438 B.n398 VSUBS 0.007583f
C439 B.n399 VSUBS 0.007583f
C440 B.n400 VSUBS 0.007583f
C441 B.n401 VSUBS 0.007583f
C442 B.n402 VSUBS 0.007583f
C443 B.n403 VSUBS 0.007583f
C444 B.n404 VSUBS 0.007583f
C445 B.n405 VSUBS 0.007583f
C446 B.n406 VSUBS 0.007583f
C447 B.n407 VSUBS 0.017171f
C448 VDD2.t5 VSUBS 0.066031f
C449 VDD2.t3 VSUBS 0.066031f
C450 VDD2.n0 VSUBS 0.361504f
C451 VDD2.t6 VSUBS 0.066031f
C452 VDD2.t4 VSUBS 0.066031f
C453 VDD2.n1 VSUBS 0.361504f
C454 VDD2.n2 VSUBS 2.10601f
C455 VDD2.t1 VSUBS 0.066031f
C456 VDD2.t7 VSUBS 0.066031f
C457 VDD2.n3 VSUBS 0.359605f
C458 VDD2.n4 VSUBS 1.85024f
C459 VDD2.t0 VSUBS 0.066031f
C460 VDD2.t2 VSUBS 0.066031f
C461 VDD2.n5 VSUBS 0.361489f
C462 VN.n0 VSUBS 0.060509f
C463 VN.t1 VSUBS 0.509812f
C464 VN.n1 VSUBS 0.244644f
C465 VN.n2 VSUBS 0.060509f
C466 VN.t4 VSUBS 0.509812f
C467 VN.n3 VSUBS 0.299915f
C468 VN.t2 VSUBS 0.643184f
C469 VN.n4 VSUBS 0.331146f
C470 VN.n5 VSUBS 0.260514f
C471 VN.n6 VSUBS 0.083514f
C472 VN.n7 VSUBS 0.048916f
C473 VN.n8 VSUBS 0.083514f
C474 VN.n9 VSUBS 0.060509f
C475 VN.n10 VSUBS 0.060509f
C476 VN.n11 VSUBS 0.084428f
C477 VN.n12 VSUBS 0.018561f
C478 VN.t3 VSUBS 0.603439f
C479 VN.n13 VSUBS 0.32188f
C480 VN.n14 VSUBS 0.046892f
C481 VN.n15 VSUBS 0.060509f
C482 VN.t0 VSUBS 0.509812f
C483 VN.n16 VSUBS 0.244644f
C484 VN.n17 VSUBS 0.060509f
C485 VN.t7 VSUBS 0.509812f
C486 VN.n18 VSUBS 0.299915f
C487 VN.t5 VSUBS 0.643184f
C488 VN.n19 VSUBS 0.331146f
C489 VN.n20 VSUBS 0.260514f
C490 VN.n21 VSUBS 0.083514f
C491 VN.n22 VSUBS 0.048916f
C492 VN.n23 VSUBS 0.083514f
C493 VN.n24 VSUBS 0.060509f
C494 VN.n25 VSUBS 0.060509f
C495 VN.n26 VSUBS 0.084428f
C496 VN.n27 VSUBS 0.018561f
C497 VN.t6 VSUBS 0.603439f
C498 VN.n28 VSUBS 0.32188f
C499 VN.n29 VSUBS 2.03276f
C500 VTAIL.t1 VSUBS 0.072542f
C501 VTAIL.t2 VSUBS 0.072542f
C502 VTAIL.n0 VSUBS 0.342714f
C503 VTAIL.n1 VSUBS 0.488839f
C504 VTAIL.n2 VSUBS 0.03071f
C505 VTAIL.n3 VSUBS 0.027734f
C506 VTAIL.n4 VSUBS 0.014903f
C507 VTAIL.n5 VSUBS 0.026419f
C508 VTAIL.n6 VSUBS 0.021747f
C509 VTAIL.t3 VSUBS 0.079879f
C510 VTAIL.n7 VSUBS 0.103045f
C511 VTAIL.n8 VSUBS 0.291255f
C512 VTAIL.n9 VSUBS 0.014903f
C513 VTAIL.n10 VSUBS 0.015779f
C514 VTAIL.n11 VSUBS 0.035225f
C515 VTAIL.n12 VSUBS 0.086082f
C516 VTAIL.n13 VSUBS 0.015779f
C517 VTAIL.n14 VSUBS 0.014903f
C518 VTAIL.n15 VSUBS 0.071304f
C519 VTAIL.n16 VSUBS 0.043537f
C520 VTAIL.n17 VSUBS 0.172977f
C521 VTAIL.n18 VSUBS 0.03071f
C522 VTAIL.n19 VSUBS 0.027734f
C523 VTAIL.n20 VSUBS 0.014903f
C524 VTAIL.n21 VSUBS 0.026419f
C525 VTAIL.n22 VSUBS 0.021747f
C526 VTAIL.t12 VSUBS 0.079879f
C527 VTAIL.n23 VSUBS 0.103045f
C528 VTAIL.n24 VSUBS 0.291255f
C529 VTAIL.n25 VSUBS 0.014903f
C530 VTAIL.n26 VSUBS 0.015779f
C531 VTAIL.n27 VSUBS 0.035225f
C532 VTAIL.n28 VSUBS 0.086082f
C533 VTAIL.n29 VSUBS 0.015779f
C534 VTAIL.n30 VSUBS 0.014903f
C535 VTAIL.n31 VSUBS 0.071304f
C536 VTAIL.n32 VSUBS 0.043537f
C537 VTAIL.n33 VSUBS 0.172977f
C538 VTAIL.t11 VSUBS 0.072542f
C539 VTAIL.t10 VSUBS 0.072542f
C540 VTAIL.n34 VSUBS 0.342714f
C541 VTAIL.n35 VSUBS 0.58687f
C542 VTAIL.n36 VSUBS 0.03071f
C543 VTAIL.n37 VSUBS 0.027734f
C544 VTAIL.n38 VSUBS 0.014903f
C545 VTAIL.n39 VSUBS 0.026419f
C546 VTAIL.n40 VSUBS 0.021747f
C547 VTAIL.t9 VSUBS 0.079879f
C548 VTAIL.n41 VSUBS 0.103045f
C549 VTAIL.n42 VSUBS 0.291255f
C550 VTAIL.n43 VSUBS 0.014903f
C551 VTAIL.n44 VSUBS 0.015779f
C552 VTAIL.n45 VSUBS 0.035225f
C553 VTAIL.n46 VSUBS 0.086082f
C554 VTAIL.n47 VSUBS 0.015779f
C555 VTAIL.n48 VSUBS 0.014903f
C556 VTAIL.n49 VSUBS 0.071304f
C557 VTAIL.n50 VSUBS 0.043537f
C558 VTAIL.n51 VSUBS 0.865948f
C559 VTAIL.n52 VSUBS 0.03071f
C560 VTAIL.n53 VSUBS 0.027734f
C561 VTAIL.n54 VSUBS 0.014903f
C562 VTAIL.n55 VSUBS 0.026419f
C563 VTAIL.n56 VSUBS 0.021747f
C564 VTAIL.t0 VSUBS 0.079879f
C565 VTAIL.n57 VSUBS 0.103045f
C566 VTAIL.n58 VSUBS 0.291255f
C567 VTAIL.n59 VSUBS 0.014903f
C568 VTAIL.n60 VSUBS 0.015779f
C569 VTAIL.n61 VSUBS 0.035225f
C570 VTAIL.n62 VSUBS 0.086082f
C571 VTAIL.n63 VSUBS 0.015779f
C572 VTAIL.n64 VSUBS 0.014903f
C573 VTAIL.n65 VSUBS 0.071304f
C574 VTAIL.n66 VSUBS 0.043537f
C575 VTAIL.n67 VSUBS 0.865948f
C576 VTAIL.t6 VSUBS 0.072542f
C577 VTAIL.t5 VSUBS 0.072542f
C578 VTAIL.n68 VSUBS 0.342716f
C579 VTAIL.n69 VSUBS 0.586868f
C580 VTAIL.n70 VSUBS 0.03071f
C581 VTAIL.n71 VSUBS 0.027734f
C582 VTAIL.n72 VSUBS 0.014903f
C583 VTAIL.n73 VSUBS 0.026419f
C584 VTAIL.n74 VSUBS 0.021747f
C585 VTAIL.t4 VSUBS 0.079879f
C586 VTAIL.n75 VSUBS 0.103045f
C587 VTAIL.n76 VSUBS 0.291255f
C588 VTAIL.n77 VSUBS 0.014903f
C589 VTAIL.n78 VSUBS 0.015779f
C590 VTAIL.n79 VSUBS 0.035225f
C591 VTAIL.n80 VSUBS 0.086082f
C592 VTAIL.n81 VSUBS 0.015779f
C593 VTAIL.n82 VSUBS 0.014903f
C594 VTAIL.n83 VSUBS 0.071304f
C595 VTAIL.n84 VSUBS 0.043537f
C596 VTAIL.n85 VSUBS 0.172977f
C597 VTAIL.n86 VSUBS 0.03071f
C598 VTAIL.n87 VSUBS 0.027734f
C599 VTAIL.n88 VSUBS 0.014903f
C600 VTAIL.n89 VSUBS 0.026419f
C601 VTAIL.n90 VSUBS 0.021747f
C602 VTAIL.t15 VSUBS 0.079879f
C603 VTAIL.n91 VSUBS 0.103045f
C604 VTAIL.n92 VSUBS 0.291255f
C605 VTAIL.n93 VSUBS 0.014903f
C606 VTAIL.n94 VSUBS 0.015779f
C607 VTAIL.n95 VSUBS 0.035225f
C608 VTAIL.n96 VSUBS 0.086082f
C609 VTAIL.n97 VSUBS 0.015779f
C610 VTAIL.n98 VSUBS 0.014903f
C611 VTAIL.n99 VSUBS 0.071304f
C612 VTAIL.n100 VSUBS 0.043537f
C613 VTAIL.n101 VSUBS 0.172977f
C614 VTAIL.t13 VSUBS 0.072542f
C615 VTAIL.t8 VSUBS 0.072542f
C616 VTAIL.n102 VSUBS 0.342716f
C617 VTAIL.n103 VSUBS 0.586868f
C618 VTAIL.n104 VSUBS 0.03071f
C619 VTAIL.n105 VSUBS 0.027734f
C620 VTAIL.n106 VSUBS 0.014903f
C621 VTAIL.n107 VSUBS 0.026419f
C622 VTAIL.n108 VSUBS 0.021747f
C623 VTAIL.t14 VSUBS 0.079879f
C624 VTAIL.n109 VSUBS 0.103045f
C625 VTAIL.n110 VSUBS 0.291255f
C626 VTAIL.n111 VSUBS 0.014903f
C627 VTAIL.n112 VSUBS 0.015779f
C628 VTAIL.n113 VSUBS 0.035225f
C629 VTAIL.n114 VSUBS 0.086082f
C630 VTAIL.n115 VSUBS 0.015779f
C631 VTAIL.n116 VSUBS 0.014903f
C632 VTAIL.n117 VSUBS 0.071304f
C633 VTAIL.n118 VSUBS 0.043537f
C634 VTAIL.n119 VSUBS 0.865948f
C635 VTAIL.n120 VSUBS 0.03071f
C636 VTAIL.n121 VSUBS 0.027734f
C637 VTAIL.n122 VSUBS 0.014903f
C638 VTAIL.n123 VSUBS 0.026419f
C639 VTAIL.n124 VSUBS 0.021747f
C640 VTAIL.t7 VSUBS 0.079879f
C641 VTAIL.n125 VSUBS 0.103045f
C642 VTAIL.n126 VSUBS 0.291255f
C643 VTAIL.n127 VSUBS 0.014903f
C644 VTAIL.n128 VSUBS 0.015779f
C645 VTAIL.n129 VSUBS 0.035225f
C646 VTAIL.n130 VSUBS 0.086082f
C647 VTAIL.n131 VSUBS 0.015779f
C648 VTAIL.n132 VSUBS 0.014903f
C649 VTAIL.n133 VSUBS 0.071304f
C650 VTAIL.n134 VSUBS 0.043537f
C651 VTAIL.n135 VSUBS 0.860748f
C652 VDD1.t1 VSUBS 0.067101f
C653 VDD1.t5 VSUBS 0.067101f
C654 VDD1.n0 VSUBS 0.367817f
C655 VDD1.t3 VSUBS 0.067101f
C656 VDD1.t0 VSUBS 0.067101f
C657 VDD1.n1 VSUBS 0.367358f
C658 VDD1.t6 VSUBS 0.067101f
C659 VDD1.t2 VSUBS 0.067101f
C660 VDD1.n2 VSUBS 0.367358f
C661 VDD1.n3 VSUBS 2.19486f
C662 VDD1.t4 VSUBS 0.067101f
C663 VDD1.t7 VSUBS 0.067101f
C664 VDD1.n4 VSUBS 0.365426f
C665 VDD1.n5 VSUBS 1.91059f
C666 VP.n0 VSUBS 0.063315f
C667 VP.t5 VSUBS 0.533456f
C668 VP.n1 VSUBS 0.25599f
C669 VP.n2 VSUBS 0.063315f
C670 VP.t4 VSUBS 0.533456f
C671 VP.n3 VSUBS 0.25599f
C672 VP.n4 VSUBS 0.063315f
C673 VP.n5 VSUBS 0.063315f
C674 VP.t1 VSUBS 0.631425f
C675 VP.t7 VSUBS 0.533456f
C676 VP.n6 VSUBS 0.25599f
C677 VP.n7 VSUBS 0.063315f
C678 VP.t2 VSUBS 0.533456f
C679 VP.n8 VSUBS 0.313825f
C680 VP.t0 VSUBS 0.673013f
C681 VP.n9 VSUBS 0.346504f
C682 VP.n10 VSUBS 0.272596f
C683 VP.n11 VSUBS 0.087387f
C684 VP.n12 VSUBS 0.051184f
C685 VP.n13 VSUBS 0.087387f
C686 VP.n14 VSUBS 0.063315f
C687 VP.n15 VSUBS 0.063315f
C688 VP.n16 VSUBS 0.088344f
C689 VP.n17 VSUBS 0.019422f
C690 VP.n18 VSUBS 0.336808f
C691 VP.n19 VSUBS 2.08511f
C692 VP.n20 VSUBS 2.14677f
C693 VP.t6 VSUBS 0.631425f
C694 VP.n21 VSUBS 0.336808f
C695 VP.n22 VSUBS 0.019422f
C696 VP.n23 VSUBS 0.088344f
C697 VP.n24 VSUBS 0.063315f
C698 VP.n25 VSUBS 0.063315f
C699 VP.n26 VSUBS 0.087387f
C700 VP.n27 VSUBS 0.051184f
C701 VP.n28 VSUBS 0.087387f
C702 VP.n29 VSUBS 0.063315f
C703 VP.n30 VSUBS 0.063315f
C704 VP.n31 VSUBS 0.088344f
C705 VP.n32 VSUBS 0.019422f
C706 VP.t3 VSUBS 0.631425f
C707 VP.n33 VSUBS 0.336808f
C708 VP.n34 VSUBS 0.049067f
.ends

