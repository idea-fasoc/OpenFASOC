* NGSPICE file created from diff_pair_sample_1075.ext - technology: sky130A

.subckt diff_pair_sample_1075 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=0.50325 ps=3.38 w=3.05 l=2.34
X1 VDD2.t4 VN.t1 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=1.1895 ps=6.88 w=3.05 l=2.34
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0 ps=0 w=3.05 l=2.34
X3 VDD2.t5 VN.t2 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0.50325 ps=3.38 w=3.05 l=2.34
X4 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=1.1895 ps=6.88 w=3.05 l=2.34
X5 VTAIL.t4 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=0.50325 ps=3.38 w=3.05 l=2.34
X6 VDD1.t3 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0.50325 ps=3.38 w=3.05 l=2.34
X7 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0 ps=0 w=3.05 l=2.34
X8 VTAIL.t8 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=0.50325 ps=3.38 w=3.05 l=2.34
X9 VDD2.t3 VN.t4 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=1.1895 ps=6.88 w=3.05 l=2.34
X10 VTAIL.t1 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=0.50325 ps=3.38 w=3.05 l=2.34
X11 VDD2.t1 VN.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0.50325 ps=3.38 w=3.05 l=2.34
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0 ps=0 w=3.05 l=2.34
X13 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.50325 pd=3.38 as=1.1895 ps=6.88 w=3.05 l=2.34
X14 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0.50325 ps=3.38 w=3.05 l=2.34
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1895 pd=6.88 as=0 ps=0 w=3.05 l=2.34
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n13 VN.n12 102.438
R11 VN.n27 VN.n26 102.438
R12 VN.n3 VN.t2 64.5298
R13 VN.n17 VN.t4 64.5298
R14 VN.n6 VN.n1 56.5193
R15 VN.n20 VN.n15 56.5193
R16 VN.n18 VN.n17 47.8803
R17 VN.n4 VN.n3 47.8803
R18 VN VN.n27 41.0853
R19 VN.n4 VN.t3 31.4129
R20 VN.n12 VN.t1 31.4129
R21 VN.n18 VN.t0 31.4129
R22 VN.n26 VN.t5 31.4129
R23 VN.n5 VN.n4 24.4675
R24 VN.n6 VN.n5 24.4675
R25 VN.n10 VN.n1 24.4675
R26 VN.n11 VN.n10 24.4675
R27 VN.n20 VN.n19 24.4675
R28 VN.n19 VN.n18 24.4675
R29 VN.n25 VN.n24 24.4675
R30 VN.n24 VN.n15 24.4675
R31 VN.n12 VN.n11 8.31928
R32 VN.n26 VN.n25 8.31928
R33 VN.n17 VN.n16 6.95571
R34 VN.n3 VN.n2 6.95571
R35 VN.n27 VN.n14 0.278367
R36 VN.n13 VN.n0 0.278367
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153454
R46 VDD2.n1 VDD2.t5 88.9055
R47 VDD2.n2 VDD2.t1 87.2346
R48 VDD2.n1 VDD2.n0 81.2628
R49 VDD2 VDD2.n3 81.2601
R50 VDD2.n2 VDD2.n1 33.8252
R51 VDD2.n3 VDD2.t2 6.4923
R52 VDD2.n3 VDD2.t3 6.4923
R53 VDD2.n0 VDD2.t0 6.4923
R54 VDD2.n0 VDD2.t4 6.4923
R55 VDD2 VDD2.n2 1.78498
R56 VTAIL.n10 VTAIL.t2 70.5558
R57 VTAIL.n7 VTAIL.t7 70.5558
R58 VTAIL.n11 VTAIL.t10 70.5557
R59 VTAIL.n2 VTAIL.t3 70.5557
R60 VTAIL.n9 VTAIL.n8 64.064
R61 VTAIL.n6 VTAIL.n5 64.064
R62 VTAIL.n1 VTAIL.n0 64.0639
R63 VTAIL.n4 VTAIL.n3 64.0639
R64 VTAIL.n6 VTAIL.n4 19.5996
R65 VTAIL.n11 VTAIL.n10 17.2979
R66 VTAIL.n0 VTAIL.t9 6.4923
R67 VTAIL.n0 VTAIL.t8 6.4923
R68 VTAIL.n3 VTAIL.t0 6.4923
R69 VTAIL.n3 VTAIL.t4 6.4923
R70 VTAIL.n8 VTAIL.t5 6.4923
R71 VTAIL.n8 VTAIL.t1 6.4923
R72 VTAIL.n5 VTAIL.t6 6.4923
R73 VTAIL.n5 VTAIL.t11 6.4923
R74 VTAIL.n7 VTAIL.n6 2.30222
R75 VTAIL.n10 VTAIL.n9 2.30222
R76 VTAIL.n4 VTAIL.n2 2.30222
R77 VTAIL VTAIL.n11 1.6686
R78 VTAIL.n9 VTAIL.n7 1.62119
R79 VTAIL.n2 VTAIL.n1 1.62119
R80 VTAIL VTAIL.n1 0.634121
R81 B.n525 B.n524 585
R82 B.n174 B.n94 585
R83 B.n173 B.n172 585
R84 B.n171 B.n170 585
R85 B.n169 B.n168 585
R86 B.n167 B.n166 585
R87 B.n165 B.n164 585
R88 B.n163 B.n162 585
R89 B.n161 B.n160 585
R90 B.n159 B.n158 585
R91 B.n157 B.n156 585
R92 B.n155 B.n154 585
R93 B.n153 B.n152 585
R94 B.n151 B.n150 585
R95 B.n149 B.n148 585
R96 B.n146 B.n145 585
R97 B.n144 B.n143 585
R98 B.n142 B.n141 585
R99 B.n140 B.n139 585
R100 B.n138 B.n137 585
R101 B.n136 B.n135 585
R102 B.n134 B.n133 585
R103 B.n132 B.n131 585
R104 B.n130 B.n129 585
R105 B.n128 B.n127 585
R106 B.n125 B.n124 585
R107 B.n123 B.n122 585
R108 B.n121 B.n120 585
R109 B.n119 B.n118 585
R110 B.n117 B.n116 585
R111 B.n115 B.n114 585
R112 B.n113 B.n112 585
R113 B.n111 B.n110 585
R114 B.n109 B.n108 585
R115 B.n107 B.n106 585
R116 B.n105 B.n104 585
R117 B.n103 B.n102 585
R118 B.n101 B.n100 585
R119 B.n75 B.n74 585
R120 B.n530 B.n529 585
R121 B.n523 B.n95 585
R122 B.n95 B.n72 585
R123 B.n522 B.n71 585
R124 B.n534 B.n71 585
R125 B.n521 B.n70 585
R126 B.n535 B.n70 585
R127 B.n520 B.n69 585
R128 B.n536 B.n69 585
R129 B.n519 B.n518 585
R130 B.n518 B.n65 585
R131 B.n517 B.n64 585
R132 B.n542 B.n64 585
R133 B.n516 B.n63 585
R134 B.n543 B.n63 585
R135 B.n515 B.n62 585
R136 B.n544 B.n62 585
R137 B.n514 B.n513 585
R138 B.n513 B.n58 585
R139 B.n512 B.n57 585
R140 B.n550 B.n57 585
R141 B.n511 B.n56 585
R142 B.n551 B.n56 585
R143 B.n510 B.n55 585
R144 B.n552 B.n55 585
R145 B.n509 B.n508 585
R146 B.n508 B.n51 585
R147 B.n507 B.n50 585
R148 B.n558 B.n50 585
R149 B.n506 B.n49 585
R150 B.n559 B.n49 585
R151 B.n505 B.n48 585
R152 B.n560 B.n48 585
R153 B.n504 B.n503 585
R154 B.n503 B.n44 585
R155 B.n502 B.n43 585
R156 B.n566 B.n43 585
R157 B.n501 B.n42 585
R158 B.n567 B.n42 585
R159 B.n500 B.n41 585
R160 B.n568 B.n41 585
R161 B.n499 B.n498 585
R162 B.n498 B.n37 585
R163 B.n497 B.n36 585
R164 B.n574 B.n36 585
R165 B.n496 B.n35 585
R166 B.n575 B.n35 585
R167 B.n495 B.n34 585
R168 B.n576 B.n34 585
R169 B.n494 B.n493 585
R170 B.n493 B.n30 585
R171 B.n492 B.n29 585
R172 B.n582 B.n29 585
R173 B.n491 B.n28 585
R174 B.n583 B.n28 585
R175 B.n490 B.n27 585
R176 B.n584 B.n27 585
R177 B.n489 B.n488 585
R178 B.n488 B.n23 585
R179 B.n487 B.n22 585
R180 B.n590 B.n22 585
R181 B.n486 B.n21 585
R182 B.n591 B.n21 585
R183 B.n485 B.n20 585
R184 B.n592 B.n20 585
R185 B.n484 B.n483 585
R186 B.n483 B.n16 585
R187 B.n482 B.n15 585
R188 B.n598 B.n15 585
R189 B.n481 B.n14 585
R190 B.n599 B.n14 585
R191 B.n480 B.n13 585
R192 B.n600 B.n13 585
R193 B.n479 B.n478 585
R194 B.n478 B.n12 585
R195 B.n477 B.n476 585
R196 B.n477 B.n8 585
R197 B.n475 B.n7 585
R198 B.n607 B.n7 585
R199 B.n474 B.n6 585
R200 B.n608 B.n6 585
R201 B.n473 B.n5 585
R202 B.n609 B.n5 585
R203 B.n472 B.n471 585
R204 B.n471 B.n4 585
R205 B.n470 B.n175 585
R206 B.n470 B.n469 585
R207 B.n460 B.n176 585
R208 B.n177 B.n176 585
R209 B.n462 B.n461 585
R210 B.n463 B.n462 585
R211 B.n459 B.n182 585
R212 B.n182 B.n181 585
R213 B.n458 B.n457 585
R214 B.n457 B.n456 585
R215 B.n184 B.n183 585
R216 B.n185 B.n184 585
R217 B.n449 B.n448 585
R218 B.n450 B.n449 585
R219 B.n447 B.n190 585
R220 B.n190 B.n189 585
R221 B.n446 B.n445 585
R222 B.n445 B.n444 585
R223 B.n192 B.n191 585
R224 B.n193 B.n192 585
R225 B.n437 B.n436 585
R226 B.n438 B.n437 585
R227 B.n435 B.n197 585
R228 B.n201 B.n197 585
R229 B.n434 B.n433 585
R230 B.n433 B.n432 585
R231 B.n199 B.n198 585
R232 B.n200 B.n199 585
R233 B.n425 B.n424 585
R234 B.n426 B.n425 585
R235 B.n423 B.n206 585
R236 B.n206 B.n205 585
R237 B.n422 B.n421 585
R238 B.n421 B.n420 585
R239 B.n208 B.n207 585
R240 B.n209 B.n208 585
R241 B.n413 B.n412 585
R242 B.n414 B.n413 585
R243 B.n411 B.n213 585
R244 B.n217 B.n213 585
R245 B.n410 B.n409 585
R246 B.n409 B.n408 585
R247 B.n215 B.n214 585
R248 B.n216 B.n215 585
R249 B.n401 B.n400 585
R250 B.n402 B.n401 585
R251 B.n399 B.n222 585
R252 B.n222 B.n221 585
R253 B.n398 B.n397 585
R254 B.n397 B.n396 585
R255 B.n224 B.n223 585
R256 B.n225 B.n224 585
R257 B.n389 B.n388 585
R258 B.n390 B.n389 585
R259 B.n387 B.n230 585
R260 B.n230 B.n229 585
R261 B.n386 B.n385 585
R262 B.n385 B.n384 585
R263 B.n232 B.n231 585
R264 B.n233 B.n232 585
R265 B.n377 B.n376 585
R266 B.n378 B.n377 585
R267 B.n375 B.n238 585
R268 B.n238 B.n237 585
R269 B.n374 B.n373 585
R270 B.n373 B.n372 585
R271 B.n240 B.n239 585
R272 B.n241 B.n240 585
R273 B.n365 B.n364 585
R274 B.n366 B.n365 585
R275 B.n363 B.n246 585
R276 B.n246 B.n245 585
R277 B.n362 B.n361 585
R278 B.n361 B.n360 585
R279 B.n248 B.n247 585
R280 B.n249 B.n248 585
R281 B.n356 B.n355 585
R282 B.n252 B.n251 585
R283 B.n352 B.n351 585
R284 B.n353 B.n352 585
R285 B.n350 B.n272 585
R286 B.n349 B.n348 585
R287 B.n347 B.n346 585
R288 B.n345 B.n344 585
R289 B.n343 B.n342 585
R290 B.n341 B.n340 585
R291 B.n339 B.n338 585
R292 B.n337 B.n336 585
R293 B.n335 B.n334 585
R294 B.n333 B.n332 585
R295 B.n331 B.n330 585
R296 B.n329 B.n328 585
R297 B.n327 B.n326 585
R298 B.n325 B.n324 585
R299 B.n323 B.n322 585
R300 B.n321 B.n320 585
R301 B.n319 B.n318 585
R302 B.n317 B.n316 585
R303 B.n315 B.n314 585
R304 B.n313 B.n312 585
R305 B.n311 B.n310 585
R306 B.n309 B.n308 585
R307 B.n307 B.n306 585
R308 B.n305 B.n304 585
R309 B.n303 B.n302 585
R310 B.n301 B.n300 585
R311 B.n299 B.n298 585
R312 B.n297 B.n296 585
R313 B.n295 B.n294 585
R314 B.n293 B.n292 585
R315 B.n291 B.n290 585
R316 B.n289 B.n288 585
R317 B.n287 B.n286 585
R318 B.n285 B.n284 585
R319 B.n283 B.n282 585
R320 B.n281 B.n280 585
R321 B.n279 B.n271 585
R322 B.n353 B.n271 585
R323 B.n357 B.n250 585
R324 B.n250 B.n249 585
R325 B.n359 B.n358 585
R326 B.n360 B.n359 585
R327 B.n244 B.n243 585
R328 B.n245 B.n244 585
R329 B.n368 B.n367 585
R330 B.n367 B.n366 585
R331 B.n369 B.n242 585
R332 B.n242 B.n241 585
R333 B.n371 B.n370 585
R334 B.n372 B.n371 585
R335 B.n236 B.n235 585
R336 B.n237 B.n236 585
R337 B.n380 B.n379 585
R338 B.n379 B.n378 585
R339 B.n381 B.n234 585
R340 B.n234 B.n233 585
R341 B.n383 B.n382 585
R342 B.n384 B.n383 585
R343 B.n228 B.n227 585
R344 B.n229 B.n228 585
R345 B.n392 B.n391 585
R346 B.n391 B.n390 585
R347 B.n393 B.n226 585
R348 B.n226 B.n225 585
R349 B.n395 B.n394 585
R350 B.n396 B.n395 585
R351 B.n220 B.n219 585
R352 B.n221 B.n220 585
R353 B.n404 B.n403 585
R354 B.n403 B.n402 585
R355 B.n405 B.n218 585
R356 B.n218 B.n216 585
R357 B.n407 B.n406 585
R358 B.n408 B.n407 585
R359 B.n212 B.n211 585
R360 B.n217 B.n212 585
R361 B.n416 B.n415 585
R362 B.n415 B.n414 585
R363 B.n417 B.n210 585
R364 B.n210 B.n209 585
R365 B.n419 B.n418 585
R366 B.n420 B.n419 585
R367 B.n204 B.n203 585
R368 B.n205 B.n204 585
R369 B.n428 B.n427 585
R370 B.n427 B.n426 585
R371 B.n429 B.n202 585
R372 B.n202 B.n200 585
R373 B.n431 B.n430 585
R374 B.n432 B.n431 585
R375 B.n196 B.n195 585
R376 B.n201 B.n196 585
R377 B.n440 B.n439 585
R378 B.n439 B.n438 585
R379 B.n441 B.n194 585
R380 B.n194 B.n193 585
R381 B.n443 B.n442 585
R382 B.n444 B.n443 585
R383 B.n188 B.n187 585
R384 B.n189 B.n188 585
R385 B.n452 B.n451 585
R386 B.n451 B.n450 585
R387 B.n453 B.n186 585
R388 B.n186 B.n185 585
R389 B.n455 B.n454 585
R390 B.n456 B.n455 585
R391 B.n180 B.n179 585
R392 B.n181 B.n180 585
R393 B.n465 B.n464 585
R394 B.n464 B.n463 585
R395 B.n466 B.n178 585
R396 B.n178 B.n177 585
R397 B.n468 B.n467 585
R398 B.n469 B.n468 585
R399 B.n3 B.n0 585
R400 B.n4 B.n3 585
R401 B.n606 B.n1 585
R402 B.n607 B.n606 585
R403 B.n605 B.n604 585
R404 B.n605 B.n8 585
R405 B.n603 B.n9 585
R406 B.n12 B.n9 585
R407 B.n602 B.n601 585
R408 B.n601 B.n600 585
R409 B.n11 B.n10 585
R410 B.n599 B.n11 585
R411 B.n597 B.n596 585
R412 B.n598 B.n597 585
R413 B.n595 B.n17 585
R414 B.n17 B.n16 585
R415 B.n594 B.n593 585
R416 B.n593 B.n592 585
R417 B.n19 B.n18 585
R418 B.n591 B.n19 585
R419 B.n589 B.n588 585
R420 B.n590 B.n589 585
R421 B.n587 B.n24 585
R422 B.n24 B.n23 585
R423 B.n586 B.n585 585
R424 B.n585 B.n584 585
R425 B.n26 B.n25 585
R426 B.n583 B.n26 585
R427 B.n581 B.n580 585
R428 B.n582 B.n581 585
R429 B.n579 B.n31 585
R430 B.n31 B.n30 585
R431 B.n578 B.n577 585
R432 B.n577 B.n576 585
R433 B.n33 B.n32 585
R434 B.n575 B.n33 585
R435 B.n573 B.n572 585
R436 B.n574 B.n573 585
R437 B.n571 B.n38 585
R438 B.n38 B.n37 585
R439 B.n570 B.n569 585
R440 B.n569 B.n568 585
R441 B.n40 B.n39 585
R442 B.n567 B.n40 585
R443 B.n565 B.n564 585
R444 B.n566 B.n565 585
R445 B.n563 B.n45 585
R446 B.n45 B.n44 585
R447 B.n562 B.n561 585
R448 B.n561 B.n560 585
R449 B.n47 B.n46 585
R450 B.n559 B.n47 585
R451 B.n557 B.n556 585
R452 B.n558 B.n557 585
R453 B.n555 B.n52 585
R454 B.n52 B.n51 585
R455 B.n554 B.n553 585
R456 B.n553 B.n552 585
R457 B.n54 B.n53 585
R458 B.n551 B.n54 585
R459 B.n549 B.n548 585
R460 B.n550 B.n549 585
R461 B.n547 B.n59 585
R462 B.n59 B.n58 585
R463 B.n546 B.n545 585
R464 B.n545 B.n544 585
R465 B.n61 B.n60 585
R466 B.n543 B.n61 585
R467 B.n541 B.n540 585
R468 B.n542 B.n541 585
R469 B.n539 B.n66 585
R470 B.n66 B.n65 585
R471 B.n538 B.n537 585
R472 B.n537 B.n536 585
R473 B.n68 B.n67 585
R474 B.n535 B.n68 585
R475 B.n533 B.n532 585
R476 B.n534 B.n533 585
R477 B.n531 B.n73 585
R478 B.n73 B.n72 585
R479 B.n610 B.n609 585
R480 B.n608 B.n2 585
R481 B.n529 B.n73 516.524
R482 B.n525 B.n95 516.524
R483 B.n271 B.n248 516.524
R484 B.n355 B.n250 516.524
R485 B.n527 B.n526 256.663
R486 B.n527 B.n93 256.663
R487 B.n527 B.n92 256.663
R488 B.n527 B.n91 256.663
R489 B.n527 B.n90 256.663
R490 B.n527 B.n89 256.663
R491 B.n527 B.n88 256.663
R492 B.n527 B.n87 256.663
R493 B.n527 B.n86 256.663
R494 B.n527 B.n85 256.663
R495 B.n527 B.n84 256.663
R496 B.n527 B.n83 256.663
R497 B.n527 B.n82 256.663
R498 B.n527 B.n81 256.663
R499 B.n527 B.n80 256.663
R500 B.n527 B.n79 256.663
R501 B.n527 B.n78 256.663
R502 B.n527 B.n77 256.663
R503 B.n527 B.n76 256.663
R504 B.n528 B.n527 256.663
R505 B.n354 B.n353 256.663
R506 B.n353 B.n253 256.663
R507 B.n353 B.n254 256.663
R508 B.n353 B.n255 256.663
R509 B.n353 B.n256 256.663
R510 B.n353 B.n257 256.663
R511 B.n353 B.n258 256.663
R512 B.n353 B.n259 256.663
R513 B.n353 B.n260 256.663
R514 B.n353 B.n261 256.663
R515 B.n353 B.n262 256.663
R516 B.n353 B.n263 256.663
R517 B.n353 B.n264 256.663
R518 B.n353 B.n265 256.663
R519 B.n353 B.n266 256.663
R520 B.n353 B.n267 256.663
R521 B.n353 B.n268 256.663
R522 B.n353 B.n269 256.663
R523 B.n353 B.n270 256.663
R524 B.n612 B.n611 256.663
R525 B.n98 B.t17 239.03
R526 B.n96 B.t6 239.03
R527 B.n276 B.t14 239.03
R528 B.n273 B.t10 239.03
R529 B.n353 B.n249 165.166
R530 B.n527 B.n72 165.166
R531 B.n100 B.n75 163.367
R532 B.n104 B.n103 163.367
R533 B.n108 B.n107 163.367
R534 B.n112 B.n111 163.367
R535 B.n116 B.n115 163.367
R536 B.n120 B.n119 163.367
R537 B.n124 B.n123 163.367
R538 B.n129 B.n128 163.367
R539 B.n133 B.n132 163.367
R540 B.n137 B.n136 163.367
R541 B.n141 B.n140 163.367
R542 B.n145 B.n144 163.367
R543 B.n150 B.n149 163.367
R544 B.n154 B.n153 163.367
R545 B.n158 B.n157 163.367
R546 B.n162 B.n161 163.367
R547 B.n166 B.n165 163.367
R548 B.n170 B.n169 163.367
R549 B.n172 B.n94 163.367
R550 B.n361 B.n248 163.367
R551 B.n361 B.n246 163.367
R552 B.n365 B.n246 163.367
R553 B.n365 B.n240 163.367
R554 B.n373 B.n240 163.367
R555 B.n373 B.n238 163.367
R556 B.n377 B.n238 163.367
R557 B.n377 B.n232 163.367
R558 B.n385 B.n232 163.367
R559 B.n385 B.n230 163.367
R560 B.n389 B.n230 163.367
R561 B.n389 B.n224 163.367
R562 B.n397 B.n224 163.367
R563 B.n397 B.n222 163.367
R564 B.n401 B.n222 163.367
R565 B.n401 B.n215 163.367
R566 B.n409 B.n215 163.367
R567 B.n409 B.n213 163.367
R568 B.n413 B.n213 163.367
R569 B.n413 B.n208 163.367
R570 B.n421 B.n208 163.367
R571 B.n421 B.n206 163.367
R572 B.n425 B.n206 163.367
R573 B.n425 B.n199 163.367
R574 B.n433 B.n199 163.367
R575 B.n433 B.n197 163.367
R576 B.n437 B.n197 163.367
R577 B.n437 B.n192 163.367
R578 B.n445 B.n192 163.367
R579 B.n445 B.n190 163.367
R580 B.n449 B.n190 163.367
R581 B.n449 B.n184 163.367
R582 B.n457 B.n184 163.367
R583 B.n457 B.n182 163.367
R584 B.n462 B.n182 163.367
R585 B.n462 B.n176 163.367
R586 B.n470 B.n176 163.367
R587 B.n471 B.n470 163.367
R588 B.n471 B.n5 163.367
R589 B.n6 B.n5 163.367
R590 B.n7 B.n6 163.367
R591 B.n477 B.n7 163.367
R592 B.n478 B.n477 163.367
R593 B.n478 B.n13 163.367
R594 B.n14 B.n13 163.367
R595 B.n15 B.n14 163.367
R596 B.n483 B.n15 163.367
R597 B.n483 B.n20 163.367
R598 B.n21 B.n20 163.367
R599 B.n22 B.n21 163.367
R600 B.n488 B.n22 163.367
R601 B.n488 B.n27 163.367
R602 B.n28 B.n27 163.367
R603 B.n29 B.n28 163.367
R604 B.n493 B.n29 163.367
R605 B.n493 B.n34 163.367
R606 B.n35 B.n34 163.367
R607 B.n36 B.n35 163.367
R608 B.n498 B.n36 163.367
R609 B.n498 B.n41 163.367
R610 B.n42 B.n41 163.367
R611 B.n43 B.n42 163.367
R612 B.n503 B.n43 163.367
R613 B.n503 B.n48 163.367
R614 B.n49 B.n48 163.367
R615 B.n50 B.n49 163.367
R616 B.n508 B.n50 163.367
R617 B.n508 B.n55 163.367
R618 B.n56 B.n55 163.367
R619 B.n57 B.n56 163.367
R620 B.n513 B.n57 163.367
R621 B.n513 B.n62 163.367
R622 B.n63 B.n62 163.367
R623 B.n64 B.n63 163.367
R624 B.n518 B.n64 163.367
R625 B.n518 B.n69 163.367
R626 B.n70 B.n69 163.367
R627 B.n71 B.n70 163.367
R628 B.n95 B.n71 163.367
R629 B.n352 B.n252 163.367
R630 B.n352 B.n272 163.367
R631 B.n348 B.n347 163.367
R632 B.n344 B.n343 163.367
R633 B.n340 B.n339 163.367
R634 B.n336 B.n335 163.367
R635 B.n332 B.n331 163.367
R636 B.n328 B.n327 163.367
R637 B.n324 B.n323 163.367
R638 B.n320 B.n319 163.367
R639 B.n316 B.n315 163.367
R640 B.n312 B.n311 163.367
R641 B.n308 B.n307 163.367
R642 B.n304 B.n303 163.367
R643 B.n300 B.n299 163.367
R644 B.n296 B.n295 163.367
R645 B.n292 B.n291 163.367
R646 B.n288 B.n287 163.367
R647 B.n284 B.n283 163.367
R648 B.n280 B.n271 163.367
R649 B.n359 B.n250 163.367
R650 B.n359 B.n244 163.367
R651 B.n367 B.n244 163.367
R652 B.n367 B.n242 163.367
R653 B.n371 B.n242 163.367
R654 B.n371 B.n236 163.367
R655 B.n379 B.n236 163.367
R656 B.n379 B.n234 163.367
R657 B.n383 B.n234 163.367
R658 B.n383 B.n228 163.367
R659 B.n391 B.n228 163.367
R660 B.n391 B.n226 163.367
R661 B.n395 B.n226 163.367
R662 B.n395 B.n220 163.367
R663 B.n403 B.n220 163.367
R664 B.n403 B.n218 163.367
R665 B.n407 B.n218 163.367
R666 B.n407 B.n212 163.367
R667 B.n415 B.n212 163.367
R668 B.n415 B.n210 163.367
R669 B.n419 B.n210 163.367
R670 B.n419 B.n204 163.367
R671 B.n427 B.n204 163.367
R672 B.n427 B.n202 163.367
R673 B.n431 B.n202 163.367
R674 B.n431 B.n196 163.367
R675 B.n439 B.n196 163.367
R676 B.n439 B.n194 163.367
R677 B.n443 B.n194 163.367
R678 B.n443 B.n188 163.367
R679 B.n451 B.n188 163.367
R680 B.n451 B.n186 163.367
R681 B.n455 B.n186 163.367
R682 B.n455 B.n180 163.367
R683 B.n464 B.n180 163.367
R684 B.n464 B.n178 163.367
R685 B.n468 B.n178 163.367
R686 B.n468 B.n3 163.367
R687 B.n610 B.n3 163.367
R688 B.n606 B.n2 163.367
R689 B.n606 B.n605 163.367
R690 B.n605 B.n9 163.367
R691 B.n601 B.n9 163.367
R692 B.n601 B.n11 163.367
R693 B.n597 B.n11 163.367
R694 B.n597 B.n17 163.367
R695 B.n593 B.n17 163.367
R696 B.n593 B.n19 163.367
R697 B.n589 B.n19 163.367
R698 B.n589 B.n24 163.367
R699 B.n585 B.n24 163.367
R700 B.n585 B.n26 163.367
R701 B.n581 B.n26 163.367
R702 B.n581 B.n31 163.367
R703 B.n577 B.n31 163.367
R704 B.n577 B.n33 163.367
R705 B.n573 B.n33 163.367
R706 B.n573 B.n38 163.367
R707 B.n569 B.n38 163.367
R708 B.n569 B.n40 163.367
R709 B.n565 B.n40 163.367
R710 B.n565 B.n45 163.367
R711 B.n561 B.n45 163.367
R712 B.n561 B.n47 163.367
R713 B.n557 B.n47 163.367
R714 B.n557 B.n52 163.367
R715 B.n553 B.n52 163.367
R716 B.n553 B.n54 163.367
R717 B.n549 B.n54 163.367
R718 B.n549 B.n59 163.367
R719 B.n545 B.n59 163.367
R720 B.n545 B.n61 163.367
R721 B.n541 B.n61 163.367
R722 B.n541 B.n66 163.367
R723 B.n537 B.n66 163.367
R724 B.n537 B.n68 163.367
R725 B.n533 B.n68 163.367
R726 B.n533 B.n73 163.367
R727 B.n96 B.t8 133.258
R728 B.n276 B.t16 133.258
R729 B.n98 B.t18 133.256
R730 B.n273 B.t13 133.256
R731 B.n360 B.n249 89.8504
R732 B.n360 B.n245 89.8504
R733 B.n366 B.n245 89.8504
R734 B.n366 B.n241 89.8504
R735 B.n372 B.n241 89.8504
R736 B.n372 B.n237 89.8504
R737 B.n378 B.n237 89.8504
R738 B.n384 B.n233 89.8504
R739 B.n384 B.n229 89.8504
R740 B.n390 B.n229 89.8504
R741 B.n390 B.n225 89.8504
R742 B.n396 B.n225 89.8504
R743 B.n396 B.n221 89.8504
R744 B.n402 B.n221 89.8504
R745 B.n402 B.n216 89.8504
R746 B.n408 B.n216 89.8504
R747 B.n408 B.n217 89.8504
R748 B.n414 B.n209 89.8504
R749 B.n420 B.n209 89.8504
R750 B.n420 B.n205 89.8504
R751 B.n426 B.n205 89.8504
R752 B.n426 B.n200 89.8504
R753 B.n432 B.n200 89.8504
R754 B.n432 B.n201 89.8504
R755 B.n438 B.n193 89.8504
R756 B.n444 B.n193 89.8504
R757 B.n444 B.n189 89.8504
R758 B.n450 B.n189 89.8504
R759 B.n450 B.n185 89.8504
R760 B.n456 B.n185 89.8504
R761 B.n463 B.n181 89.8504
R762 B.n463 B.n177 89.8504
R763 B.n469 B.n177 89.8504
R764 B.n469 B.n4 89.8504
R765 B.n609 B.n4 89.8504
R766 B.n609 B.n608 89.8504
R767 B.n608 B.n607 89.8504
R768 B.n607 B.n8 89.8504
R769 B.n12 B.n8 89.8504
R770 B.n600 B.n12 89.8504
R771 B.n600 B.n599 89.8504
R772 B.n598 B.n16 89.8504
R773 B.n592 B.n16 89.8504
R774 B.n592 B.n591 89.8504
R775 B.n591 B.n590 89.8504
R776 B.n590 B.n23 89.8504
R777 B.n584 B.n23 89.8504
R778 B.n583 B.n582 89.8504
R779 B.n582 B.n30 89.8504
R780 B.n576 B.n30 89.8504
R781 B.n576 B.n575 89.8504
R782 B.n575 B.n574 89.8504
R783 B.n574 B.n37 89.8504
R784 B.n568 B.n37 89.8504
R785 B.n567 B.n566 89.8504
R786 B.n566 B.n44 89.8504
R787 B.n560 B.n44 89.8504
R788 B.n560 B.n559 89.8504
R789 B.n559 B.n558 89.8504
R790 B.n558 B.n51 89.8504
R791 B.n552 B.n51 89.8504
R792 B.n552 B.n551 89.8504
R793 B.n551 B.n550 89.8504
R794 B.n550 B.n58 89.8504
R795 B.n544 B.n543 89.8504
R796 B.n543 B.n542 89.8504
R797 B.n542 B.n65 89.8504
R798 B.n536 B.n65 89.8504
R799 B.n536 B.n535 89.8504
R800 B.n535 B.n534 89.8504
R801 B.n534 B.n72 89.8504
R802 B.n456 B.t3 87.2077
R803 B.t5 B.n598 87.2077
R804 B.n97 B.t9 81.4763
R805 B.n277 B.t15 81.4763
R806 B.n99 B.t19 81.4745
R807 B.n274 B.t12 81.4745
R808 B.n438 B.t4 79.2798
R809 B.n584 B.t1 79.2798
R810 B.n529 B.n528 71.676
R811 B.n100 B.n76 71.676
R812 B.n104 B.n77 71.676
R813 B.n108 B.n78 71.676
R814 B.n112 B.n79 71.676
R815 B.n116 B.n80 71.676
R816 B.n120 B.n81 71.676
R817 B.n124 B.n82 71.676
R818 B.n129 B.n83 71.676
R819 B.n133 B.n84 71.676
R820 B.n137 B.n85 71.676
R821 B.n141 B.n86 71.676
R822 B.n145 B.n87 71.676
R823 B.n150 B.n88 71.676
R824 B.n154 B.n89 71.676
R825 B.n158 B.n90 71.676
R826 B.n162 B.n91 71.676
R827 B.n166 B.n92 71.676
R828 B.n170 B.n93 71.676
R829 B.n526 B.n94 71.676
R830 B.n526 B.n525 71.676
R831 B.n172 B.n93 71.676
R832 B.n169 B.n92 71.676
R833 B.n165 B.n91 71.676
R834 B.n161 B.n90 71.676
R835 B.n157 B.n89 71.676
R836 B.n153 B.n88 71.676
R837 B.n149 B.n87 71.676
R838 B.n144 B.n86 71.676
R839 B.n140 B.n85 71.676
R840 B.n136 B.n84 71.676
R841 B.n132 B.n83 71.676
R842 B.n128 B.n82 71.676
R843 B.n123 B.n81 71.676
R844 B.n119 B.n80 71.676
R845 B.n115 B.n79 71.676
R846 B.n111 B.n78 71.676
R847 B.n107 B.n77 71.676
R848 B.n103 B.n76 71.676
R849 B.n528 B.n75 71.676
R850 B.n355 B.n354 71.676
R851 B.n272 B.n253 71.676
R852 B.n347 B.n254 71.676
R853 B.n343 B.n255 71.676
R854 B.n339 B.n256 71.676
R855 B.n335 B.n257 71.676
R856 B.n331 B.n258 71.676
R857 B.n327 B.n259 71.676
R858 B.n323 B.n260 71.676
R859 B.n319 B.n261 71.676
R860 B.n315 B.n262 71.676
R861 B.n311 B.n263 71.676
R862 B.n307 B.n264 71.676
R863 B.n303 B.n265 71.676
R864 B.n299 B.n266 71.676
R865 B.n295 B.n267 71.676
R866 B.n291 B.n268 71.676
R867 B.n287 B.n269 71.676
R868 B.n283 B.n270 71.676
R869 B.n354 B.n252 71.676
R870 B.n348 B.n253 71.676
R871 B.n344 B.n254 71.676
R872 B.n340 B.n255 71.676
R873 B.n336 B.n256 71.676
R874 B.n332 B.n257 71.676
R875 B.n328 B.n258 71.676
R876 B.n324 B.n259 71.676
R877 B.n320 B.n260 71.676
R878 B.n316 B.n261 71.676
R879 B.n312 B.n262 71.676
R880 B.n308 B.n263 71.676
R881 B.n304 B.n264 71.676
R882 B.n300 B.n265 71.676
R883 B.n296 B.n266 71.676
R884 B.n292 B.n267 71.676
R885 B.n288 B.n268 71.676
R886 B.n284 B.n269 71.676
R887 B.n280 B.n270 71.676
R888 B.n611 B.n610 71.676
R889 B.n611 B.n2 71.676
R890 B.t11 B.n233 71.3518
R891 B.t7 B.n58 71.3518
R892 B.n414 B.t0 66.0666
R893 B.n568 B.t2 66.0666
R894 B.n126 B.n99 59.5399
R895 B.n147 B.n97 59.5399
R896 B.n278 B.n277 59.5399
R897 B.n275 B.n274 59.5399
R898 B.n99 B.n98 51.7823
R899 B.n97 B.n96 51.7823
R900 B.n277 B.n276 51.7823
R901 B.n274 B.n273 51.7823
R902 B.n357 B.n356 33.5615
R903 B.n279 B.n247 33.5615
R904 B.n524 B.n523 33.5615
R905 B.n531 B.n530 33.5615
R906 B.n217 B.t0 23.7843
R907 B.t2 B.n567 23.7843
R908 B.n378 B.t11 18.499
R909 B.n544 B.t7 18.499
R910 B B.n612 18.0485
R911 B.n358 B.n357 10.6151
R912 B.n358 B.n243 10.6151
R913 B.n368 B.n243 10.6151
R914 B.n369 B.n368 10.6151
R915 B.n370 B.n369 10.6151
R916 B.n370 B.n235 10.6151
R917 B.n380 B.n235 10.6151
R918 B.n381 B.n380 10.6151
R919 B.n382 B.n381 10.6151
R920 B.n382 B.n227 10.6151
R921 B.n392 B.n227 10.6151
R922 B.n393 B.n392 10.6151
R923 B.n394 B.n393 10.6151
R924 B.n394 B.n219 10.6151
R925 B.n404 B.n219 10.6151
R926 B.n405 B.n404 10.6151
R927 B.n406 B.n405 10.6151
R928 B.n406 B.n211 10.6151
R929 B.n416 B.n211 10.6151
R930 B.n417 B.n416 10.6151
R931 B.n418 B.n417 10.6151
R932 B.n418 B.n203 10.6151
R933 B.n428 B.n203 10.6151
R934 B.n429 B.n428 10.6151
R935 B.n430 B.n429 10.6151
R936 B.n430 B.n195 10.6151
R937 B.n440 B.n195 10.6151
R938 B.n441 B.n440 10.6151
R939 B.n442 B.n441 10.6151
R940 B.n442 B.n187 10.6151
R941 B.n452 B.n187 10.6151
R942 B.n453 B.n452 10.6151
R943 B.n454 B.n453 10.6151
R944 B.n454 B.n179 10.6151
R945 B.n465 B.n179 10.6151
R946 B.n466 B.n465 10.6151
R947 B.n467 B.n466 10.6151
R948 B.n467 B.n0 10.6151
R949 B.n356 B.n251 10.6151
R950 B.n351 B.n251 10.6151
R951 B.n351 B.n350 10.6151
R952 B.n350 B.n349 10.6151
R953 B.n349 B.n346 10.6151
R954 B.n346 B.n345 10.6151
R955 B.n345 B.n342 10.6151
R956 B.n342 B.n341 10.6151
R957 B.n341 B.n338 10.6151
R958 B.n338 B.n337 10.6151
R959 B.n337 B.n334 10.6151
R960 B.n334 B.n333 10.6151
R961 B.n333 B.n330 10.6151
R962 B.n330 B.n329 10.6151
R963 B.n326 B.n325 10.6151
R964 B.n325 B.n322 10.6151
R965 B.n322 B.n321 10.6151
R966 B.n321 B.n318 10.6151
R967 B.n318 B.n317 10.6151
R968 B.n317 B.n314 10.6151
R969 B.n314 B.n313 10.6151
R970 B.n313 B.n310 10.6151
R971 B.n310 B.n309 10.6151
R972 B.n306 B.n305 10.6151
R973 B.n305 B.n302 10.6151
R974 B.n302 B.n301 10.6151
R975 B.n301 B.n298 10.6151
R976 B.n298 B.n297 10.6151
R977 B.n297 B.n294 10.6151
R978 B.n294 B.n293 10.6151
R979 B.n293 B.n290 10.6151
R980 B.n290 B.n289 10.6151
R981 B.n289 B.n286 10.6151
R982 B.n286 B.n285 10.6151
R983 B.n285 B.n282 10.6151
R984 B.n282 B.n281 10.6151
R985 B.n281 B.n279 10.6151
R986 B.n362 B.n247 10.6151
R987 B.n363 B.n362 10.6151
R988 B.n364 B.n363 10.6151
R989 B.n364 B.n239 10.6151
R990 B.n374 B.n239 10.6151
R991 B.n375 B.n374 10.6151
R992 B.n376 B.n375 10.6151
R993 B.n376 B.n231 10.6151
R994 B.n386 B.n231 10.6151
R995 B.n387 B.n386 10.6151
R996 B.n388 B.n387 10.6151
R997 B.n388 B.n223 10.6151
R998 B.n398 B.n223 10.6151
R999 B.n399 B.n398 10.6151
R1000 B.n400 B.n399 10.6151
R1001 B.n400 B.n214 10.6151
R1002 B.n410 B.n214 10.6151
R1003 B.n411 B.n410 10.6151
R1004 B.n412 B.n411 10.6151
R1005 B.n412 B.n207 10.6151
R1006 B.n422 B.n207 10.6151
R1007 B.n423 B.n422 10.6151
R1008 B.n424 B.n423 10.6151
R1009 B.n424 B.n198 10.6151
R1010 B.n434 B.n198 10.6151
R1011 B.n435 B.n434 10.6151
R1012 B.n436 B.n435 10.6151
R1013 B.n436 B.n191 10.6151
R1014 B.n446 B.n191 10.6151
R1015 B.n447 B.n446 10.6151
R1016 B.n448 B.n447 10.6151
R1017 B.n448 B.n183 10.6151
R1018 B.n458 B.n183 10.6151
R1019 B.n459 B.n458 10.6151
R1020 B.n461 B.n459 10.6151
R1021 B.n461 B.n460 10.6151
R1022 B.n460 B.n175 10.6151
R1023 B.n472 B.n175 10.6151
R1024 B.n473 B.n472 10.6151
R1025 B.n474 B.n473 10.6151
R1026 B.n475 B.n474 10.6151
R1027 B.n476 B.n475 10.6151
R1028 B.n479 B.n476 10.6151
R1029 B.n480 B.n479 10.6151
R1030 B.n481 B.n480 10.6151
R1031 B.n482 B.n481 10.6151
R1032 B.n484 B.n482 10.6151
R1033 B.n485 B.n484 10.6151
R1034 B.n486 B.n485 10.6151
R1035 B.n487 B.n486 10.6151
R1036 B.n489 B.n487 10.6151
R1037 B.n490 B.n489 10.6151
R1038 B.n491 B.n490 10.6151
R1039 B.n492 B.n491 10.6151
R1040 B.n494 B.n492 10.6151
R1041 B.n495 B.n494 10.6151
R1042 B.n496 B.n495 10.6151
R1043 B.n497 B.n496 10.6151
R1044 B.n499 B.n497 10.6151
R1045 B.n500 B.n499 10.6151
R1046 B.n501 B.n500 10.6151
R1047 B.n502 B.n501 10.6151
R1048 B.n504 B.n502 10.6151
R1049 B.n505 B.n504 10.6151
R1050 B.n506 B.n505 10.6151
R1051 B.n507 B.n506 10.6151
R1052 B.n509 B.n507 10.6151
R1053 B.n510 B.n509 10.6151
R1054 B.n511 B.n510 10.6151
R1055 B.n512 B.n511 10.6151
R1056 B.n514 B.n512 10.6151
R1057 B.n515 B.n514 10.6151
R1058 B.n516 B.n515 10.6151
R1059 B.n517 B.n516 10.6151
R1060 B.n519 B.n517 10.6151
R1061 B.n520 B.n519 10.6151
R1062 B.n521 B.n520 10.6151
R1063 B.n522 B.n521 10.6151
R1064 B.n523 B.n522 10.6151
R1065 B.n604 B.n1 10.6151
R1066 B.n604 B.n603 10.6151
R1067 B.n603 B.n602 10.6151
R1068 B.n602 B.n10 10.6151
R1069 B.n596 B.n10 10.6151
R1070 B.n596 B.n595 10.6151
R1071 B.n595 B.n594 10.6151
R1072 B.n594 B.n18 10.6151
R1073 B.n588 B.n18 10.6151
R1074 B.n588 B.n587 10.6151
R1075 B.n587 B.n586 10.6151
R1076 B.n586 B.n25 10.6151
R1077 B.n580 B.n25 10.6151
R1078 B.n580 B.n579 10.6151
R1079 B.n579 B.n578 10.6151
R1080 B.n578 B.n32 10.6151
R1081 B.n572 B.n32 10.6151
R1082 B.n572 B.n571 10.6151
R1083 B.n571 B.n570 10.6151
R1084 B.n570 B.n39 10.6151
R1085 B.n564 B.n39 10.6151
R1086 B.n564 B.n563 10.6151
R1087 B.n563 B.n562 10.6151
R1088 B.n562 B.n46 10.6151
R1089 B.n556 B.n46 10.6151
R1090 B.n556 B.n555 10.6151
R1091 B.n555 B.n554 10.6151
R1092 B.n554 B.n53 10.6151
R1093 B.n548 B.n53 10.6151
R1094 B.n548 B.n547 10.6151
R1095 B.n547 B.n546 10.6151
R1096 B.n546 B.n60 10.6151
R1097 B.n540 B.n60 10.6151
R1098 B.n540 B.n539 10.6151
R1099 B.n539 B.n538 10.6151
R1100 B.n538 B.n67 10.6151
R1101 B.n532 B.n67 10.6151
R1102 B.n532 B.n531 10.6151
R1103 B.n530 B.n74 10.6151
R1104 B.n101 B.n74 10.6151
R1105 B.n102 B.n101 10.6151
R1106 B.n105 B.n102 10.6151
R1107 B.n106 B.n105 10.6151
R1108 B.n109 B.n106 10.6151
R1109 B.n110 B.n109 10.6151
R1110 B.n113 B.n110 10.6151
R1111 B.n114 B.n113 10.6151
R1112 B.n117 B.n114 10.6151
R1113 B.n118 B.n117 10.6151
R1114 B.n121 B.n118 10.6151
R1115 B.n122 B.n121 10.6151
R1116 B.n125 B.n122 10.6151
R1117 B.n130 B.n127 10.6151
R1118 B.n131 B.n130 10.6151
R1119 B.n134 B.n131 10.6151
R1120 B.n135 B.n134 10.6151
R1121 B.n138 B.n135 10.6151
R1122 B.n139 B.n138 10.6151
R1123 B.n142 B.n139 10.6151
R1124 B.n143 B.n142 10.6151
R1125 B.n146 B.n143 10.6151
R1126 B.n151 B.n148 10.6151
R1127 B.n152 B.n151 10.6151
R1128 B.n155 B.n152 10.6151
R1129 B.n156 B.n155 10.6151
R1130 B.n159 B.n156 10.6151
R1131 B.n160 B.n159 10.6151
R1132 B.n163 B.n160 10.6151
R1133 B.n164 B.n163 10.6151
R1134 B.n167 B.n164 10.6151
R1135 B.n168 B.n167 10.6151
R1136 B.n171 B.n168 10.6151
R1137 B.n173 B.n171 10.6151
R1138 B.n174 B.n173 10.6151
R1139 B.n524 B.n174 10.6151
R1140 B.n201 B.t4 10.5711
R1141 B.t1 B.n583 10.5711
R1142 B.n329 B.n275 9.36635
R1143 B.n306 B.n278 9.36635
R1144 B.n126 B.n125 9.36635
R1145 B.n148 B.n147 9.36635
R1146 B.n612 B.n0 8.11757
R1147 B.n612 B.n1 8.11757
R1148 B.t3 B.n181 2.64314
R1149 B.n599 B.t5 2.64314
R1150 B.n326 B.n275 1.24928
R1151 B.n309 B.n278 1.24928
R1152 B.n127 B.n126 1.24928
R1153 B.n147 B.n146 1.24928
R1154 VP.n11 VP.n8 161.3
R1155 VP.n13 VP.n12 161.3
R1156 VP.n14 VP.n7 161.3
R1157 VP.n16 VP.n15 161.3
R1158 VP.n17 VP.n6 161.3
R1159 VP.n37 VP.n0 161.3
R1160 VP.n36 VP.n35 161.3
R1161 VP.n34 VP.n1 161.3
R1162 VP.n33 VP.n32 161.3
R1163 VP.n31 VP.n2 161.3
R1164 VP.n30 VP.n29 161.3
R1165 VP.n28 VP.n3 161.3
R1166 VP.n27 VP.n26 161.3
R1167 VP.n25 VP.n4 161.3
R1168 VP.n24 VP.n23 161.3
R1169 VP.n22 VP.n5 161.3
R1170 VP.n21 VP.n20 102.438
R1171 VP.n39 VP.n38 102.438
R1172 VP.n19 VP.n18 102.438
R1173 VP.n9 VP.t2 64.5298
R1174 VP.n26 VP.n25 56.5193
R1175 VP.n32 VP.n1 56.5193
R1176 VP.n12 VP.n7 56.5193
R1177 VP.n10 VP.n9 47.8803
R1178 VP.n21 VP.n19 40.8064
R1179 VP.n30 VP.t1 31.4129
R1180 VP.n20 VP.t5 31.4129
R1181 VP.n38 VP.t4 31.4129
R1182 VP.n10 VP.t3 31.4129
R1183 VP.n18 VP.t0 31.4129
R1184 VP.n24 VP.n5 24.4675
R1185 VP.n25 VP.n24 24.4675
R1186 VP.n26 VP.n3 24.4675
R1187 VP.n30 VP.n3 24.4675
R1188 VP.n31 VP.n30 24.4675
R1189 VP.n32 VP.n31 24.4675
R1190 VP.n36 VP.n1 24.4675
R1191 VP.n37 VP.n36 24.4675
R1192 VP.n16 VP.n7 24.4675
R1193 VP.n17 VP.n16 24.4675
R1194 VP.n11 VP.n10 24.4675
R1195 VP.n12 VP.n11 24.4675
R1196 VP.n20 VP.n5 8.31928
R1197 VP.n38 VP.n37 8.31928
R1198 VP.n18 VP.n17 8.31928
R1199 VP.n9 VP.n8 6.95571
R1200 VP.n19 VP.n6 0.278367
R1201 VP.n22 VP.n21 0.278367
R1202 VP.n39 VP.n0 0.278367
R1203 VP.n13 VP.n8 0.189894
R1204 VP.n14 VP.n13 0.189894
R1205 VP.n15 VP.n14 0.189894
R1206 VP.n15 VP.n6 0.189894
R1207 VP.n23 VP.n22 0.189894
R1208 VP.n23 VP.n4 0.189894
R1209 VP.n27 VP.n4 0.189894
R1210 VP.n28 VP.n27 0.189894
R1211 VP.n29 VP.n28 0.189894
R1212 VP.n29 VP.n2 0.189894
R1213 VP.n33 VP.n2 0.189894
R1214 VP.n34 VP.n33 0.189894
R1215 VP.n35 VP.n34 0.189894
R1216 VP.n35 VP.n0 0.189894
R1217 VP VP.n39 0.153454
R1218 VDD1 VDD1.t3 89.0191
R1219 VDD1.n1 VDD1.t0 88.9055
R1220 VDD1.n1 VDD1.n0 81.2628
R1221 VDD1.n3 VDD1.n2 80.7428
R1222 VDD1.n3 VDD1.n1 35.5591
R1223 VDD1.n2 VDD1.t2 6.4923
R1224 VDD1.n2 VDD1.t5 6.4923
R1225 VDD1.n0 VDD1.t4 6.4923
R1226 VDD1.n0 VDD1.t1 6.4923
R1227 VDD1 VDD1.n3 0.517741
C0 VDD1 VDD2 1.30508f
C1 VDD2 VN 1.95691f
C2 VP VDD2 0.441367f
C3 VTAIL VDD2 4.3711f
C4 VDD1 VN 0.155545f
C5 VP VDD1 2.24035f
C6 VP VN 5.02707f
C7 VTAIL VDD1 4.32001f
C8 VTAIL VN 2.6294f
C9 VTAIL VP 2.64356f
C10 VDD2 B 4.028777f
C11 VDD1 B 4.48963f
C12 VTAIL B 3.755956f
C13 VN B 11.056931f
C14 VP B 9.92531f
C15 VDD1.t3 B 0.514412f
C16 VDD1.t0 B 0.513812f
C17 VDD1.t4 B 0.054601f
C18 VDD1.t1 B 0.054601f
C19 VDD1.n0 B 0.39726f
C20 VDD1.n1 B 2.11887f
C21 VDD1.t2 B 0.054601f
C22 VDD1.t5 B 0.054601f
C23 VDD1.n2 B 0.394711f
C24 VDD1.n3 B 1.82346f
C25 VP.n0 B 0.041951f
C26 VP.t4 B 0.566879f
C27 VP.n1 B 0.038918f
C28 VP.n2 B 0.03182f
C29 VP.t1 B 0.566879f
C30 VP.n3 B 0.059304f
C31 VP.n4 B 0.03182f
C32 VP.n5 B 0.03998f
C33 VP.n6 B 0.041951f
C34 VP.t0 B 0.566879f
C35 VP.n7 B 0.038918f
C36 VP.n8 B 0.299022f
C37 VP.t3 B 0.566879f
C38 VP.t2 B 0.784226f
C39 VP.n9 B 0.31219f
C40 VP.n10 B 0.344913f
C41 VP.n11 B 0.059304f
C42 VP.n12 B 0.053991f
C43 VP.n13 B 0.03182f
C44 VP.n14 B 0.03182f
C45 VP.n15 B 0.03182f
C46 VP.n16 B 0.059304f
C47 VP.n17 B 0.03998f
C48 VP.n18 B 0.334079f
C49 VP.n19 B 1.28889f
C50 VP.t5 B 0.566879f
C51 VP.n20 B 0.334079f
C52 VP.n21 B 1.31692f
C53 VP.n22 B 0.041951f
C54 VP.n23 B 0.03182f
C55 VP.n24 B 0.059304f
C56 VP.n25 B 0.038918f
C57 VP.n26 B 0.053991f
C58 VP.n27 B 0.03182f
C59 VP.n28 B 0.03182f
C60 VP.n29 B 0.03182f
C61 VP.n30 B 0.271449f
C62 VP.n31 B 0.059304f
C63 VP.n32 B 0.053991f
C64 VP.n33 B 0.03182f
C65 VP.n34 B 0.03182f
C66 VP.n35 B 0.03182f
C67 VP.n36 B 0.059304f
C68 VP.n37 B 0.03998f
C69 VP.n38 B 0.334079f
C70 VP.n39 B 0.050348f
C71 VTAIL.t9 B 0.074206f
C72 VTAIL.t8 B 0.074206f
C73 VTAIL.n0 B 0.473398f
C74 VTAIL.n1 B 0.492818f
C75 VTAIL.t3 B 0.620427f
C76 VTAIL.n2 B 0.713656f
C77 VTAIL.t0 B 0.074206f
C78 VTAIL.t4 B 0.074206f
C79 VTAIL.n3 B 0.473398f
C80 VTAIL.n4 B 1.63328f
C81 VTAIL.t6 B 0.074206f
C82 VTAIL.t11 B 0.074206f
C83 VTAIL.n5 B 0.473402f
C84 VTAIL.n6 B 1.63328f
C85 VTAIL.t7 B 0.62043f
C86 VTAIL.n7 B 0.713653f
C87 VTAIL.t5 B 0.074206f
C88 VTAIL.t1 B 0.074206f
C89 VTAIL.n8 B 0.473402f
C90 VTAIL.n9 B 0.658302f
C91 VTAIL.t2 B 0.62043f
C92 VTAIL.n10 B 1.46028f
C93 VTAIL.t10 B 0.620427f
C94 VTAIL.n11 B 1.39743f
C95 VDD2.t5 B 0.352347f
C96 VDD2.t0 B 0.037443f
C97 VDD2.t4 B 0.037443f
C98 VDD2.n0 B 0.272422f
C99 VDD2.n1 B 1.38549f
C100 VDD2.t1 B 0.347834f
C101 VDD2.n2 B 1.23375f
C102 VDD2.t2 B 0.037443f
C103 VDD2.t3 B 0.037443f
C104 VDD2.n3 B 0.272408f
C105 VN.n0 B 0.032386f
C106 VN.t1 B 0.437623f
C107 VN.n1 B 0.030044f
C108 VN.n2 B 0.230841f
C109 VN.t3 B 0.437623f
C110 VN.t2 B 0.605412f
C111 VN.n3 B 0.241007f
C112 VN.n4 B 0.266269f
C113 VN.n5 B 0.045782f
C114 VN.n6 B 0.04168f
C115 VN.n7 B 0.024565f
C116 VN.n8 B 0.024565f
C117 VN.n9 B 0.024565f
C118 VN.n10 B 0.045782f
C119 VN.n11 B 0.030864f
C120 VN.n12 B 0.257905f
C121 VN.n13 B 0.038868f
C122 VN.n14 B 0.032386f
C123 VN.t5 B 0.437623f
C124 VN.n15 B 0.030044f
C125 VN.n16 B 0.230841f
C126 VN.t0 B 0.437623f
C127 VN.t4 B 0.605412f
C128 VN.n17 B 0.241007f
C129 VN.n18 B 0.266269f
C130 VN.n19 B 0.045782f
C131 VN.n20 B 0.04168f
C132 VN.n21 B 0.024565f
C133 VN.n22 B 0.024565f
C134 VN.n23 B 0.024565f
C135 VN.n24 B 0.045782f
C136 VN.n25 B 0.030864f
C137 VN.n26 B 0.257905f
C138 VN.n27 B 1.00868f
.ends

