* NGSPICE file created from diff_pair_sample_1040.ext - technology: sky130A

.subckt diff_pair_sample_1040 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
X1 VDD1.t7 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
X2 VTAIL.t13 VN.t1 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
X3 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=0 ps=0 w=18.92 l=0.34
X4 VTAIL.t15 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
X5 VDD2.t4 VN.t3 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
X6 VDD2.t3 VN.t4 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=7.3788 ps=38.62 w=18.92 l=0.34
X7 VDD2.t2 VN.t5 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=7.3788 ps=38.62 w=18.92 l=0.34
X8 VTAIL.t0 VP.t1 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=3.1218 ps=19.25 w=18.92 l=0.34
X9 VTAIL.t10 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=3.1218 ps=19.25 w=18.92 l=0.34
X10 VDD1.t5 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=7.3788 ps=38.62 w=18.92 l=0.34
X11 VTAIL.t14 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=3.1218 ps=19.25 w=18.92 l=0.34
X12 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=0 ps=0 w=18.92 l=0.34
X13 VTAIL.t4 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
X14 VTAIL.t6 VP.t4 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
X15 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=7.3788 ps=38.62 w=18.92 l=0.34
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=0 ps=0 w=18.92 l=0.34
X17 VTAIL.t7 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=3.1218 ps=19.25 w=18.92 l=0.34
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.3788 pd=38.62 as=0 ps=0 w=18.92 l=0.34
X19 VDD1.t0 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1218 pd=19.25 as=3.1218 ps=19.25 w=18.92 l=0.34
R0 VN.n1 VN.t6 1486.58
R1 VN.n7 VN.t5 1486.58
R2 VN.n4 VN.t4 1470.47
R3 VN.n10 VN.t7 1470.47
R4 VN.n2 VN.t3 1458.05
R5 VN.n3 VN.t2 1458.05
R6 VN.n8 VN.t1 1458.05
R7 VN.n9 VN.t0 1458.05
R8 VN.n5 VN.n4 161.3
R9 VN.n11 VN.n10 161.3
R10 VN.n9 VN.n6 161.3
R11 VN.n3 VN.n0 161.3
R12 VN.n7 VN.n6 72.8343
R13 VN.n1 VN.n0 72.8343
R14 VN.n3 VN.n2 48.2005
R15 VN.n9 VN.n8 48.2005
R16 VN VN.n11 46.0024
R17 VN.n4 VN.n3 35.7853
R18 VN.n10 VN.n9 35.7853
R19 VN.n8 VN.n7 16.0984
R20 VN.n2 VN.n1 16.0984
R21 VN.n11 VN.n6 0.189894
R22 VN.n5 VN.n0 0.189894
R23 VN VN.n5 0.0516364
R24 VTAIL.n850 VTAIL.n750 289.615
R25 VTAIL.n102 VTAIL.n2 289.615
R26 VTAIL.n208 VTAIL.n108 289.615
R27 VTAIL.n316 VTAIL.n216 289.615
R28 VTAIL.n744 VTAIL.n644 289.615
R29 VTAIL.n636 VTAIL.n536 289.615
R30 VTAIL.n530 VTAIL.n430 289.615
R31 VTAIL.n422 VTAIL.n322 289.615
R32 VTAIL.n785 VTAIL.n784 185
R33 VTAIL.n782 VTAIL.n781 185
R34 VTAIL.n791 VTAIL.n790 185
R35 VTAIL.n793 VTAIL.n792 185
R36 VTAIL.n778 VTAIL.n777 185
R37 VTAIL.n799 VTAIL.n798 185
R38 VTAIL.n801 VTAIL.n800 185
R39 VTAIL.n774 VTAIL.n773 185
R40 VTAIL.n807 VTAIL.n806 185
R41 VTAIL.n809 VTAIL.n808 185
R42 VTAIL.n770 VTAIL.n769 185
R43 VTAIL.n815 VTAIL.n814 185
R44 VTAIL.n817 VTAIL.n816 185
R45 VTAIL.n766 VTAIL.n765 185
R46 VTAIL.n823 VTAIL.n822 185
R47 VTAIL.n826 VTAIL.n825 185
R48 VTAIL.n824 VTAIL.n762 185
R49 VTAIL.n831 VTAIL.n761 185
R50 VTAIL.n833 VTAIL.n832 185
R51 VTAIL.n835 VTAIL.n834 185
R52 VTAIL.n758 VTAIL.n757 185
R53 VTAIL.n841 VTAIL.n840 185
R54 VTAIL.n843 VTAIL.n842 185
R55 VTAIL.n754 VTAIL.n753 185
R56 VTAIL.n849 VTAIL.n848 185
R57 VTAIL.n851 VTAIL.n850 185
R58 VTAIL.n37 VTAIL.n36 185
R59 VTAIL.n34 VTAIL.n33 185
R60 VTAIL.n43 VTAIL.n42 185
R61 VTAIL.n45 VTAIL.n44 185
R62 VTAIL.n30 VTAIL.n29 185
R63 VTAIL.n51 VTAIL.n50 185
R64 VTAIL.n53 VTAIL.n52 185
R65 VTAIL.n26 VTAIL.n25 185
R66 VTAIL.n59 VTAIL.n58 185
R67 VTAIL.n61 VTAIL.n60 185
R68 VTAIL.n22 VTAIL.n21 185
R69 VTAIL.n67 VTAIL.n66 185
R70 VTAIL.n69 VTAIL.n68 185
R71 VTAIL.n18 VTAIL.n17 185
R72 VTAIL.n75 VTAIL.n74 185
R73 VTAIL.n78 VTAIL.n77 185
R74 VTAIL.n76 VTAIL.n14 185
R75 VTAIL.n83 VTAIL.n13 185
R76 VTAIL.n85 VTAIL.n84 185
R77 VTAIL.n87 VTAIL.n86 185
R78 VTAIL.n10 VTAIL.n9 185
R79 VTAIL.n93 VTAIL.n92 185
R80 VTAIL.n95 VTAIL.n94 185
R81 VTAIL.n6 VTAIL.n5 185
R82 VTAIL.n101 VTAIL.n100 185
R83 VTAIL.n103 VTAIL.n102 185
R84 VTAIL.n143 VTAIL.n142 185
R85 VTAIL.n140 VTAIL.n139 185
R86 VTAIL.n149 VTAIL.n148 185
R87 VTAIL.n151 VTAIL.n150 185
R88 VTAIL.n136 VTAIL.n135 185
R89 VTAIL.n157 VTAIL.n156 185
R90 VTAIL.n159 VTAIL.n158 185
R91 VTAIL.n132 VTAIL.n131 185
R92 VTAIL.n165 VTAIL.n164 185
R93 VTAIL.n167 VTAIL.n166 185
R94 VTAIL.n128 VTAIL.n127 185
R95 VTAIL.n173 VTAIL.n172 185
R96 VTAIL.n175 VTAIL.n174 185
R97 VTAIL.n124 VTAIL.n123 185
R98 VTAIL.n181 VTAIL.n180 185
R99 VTAIL.n184 VTAIL.n183 185
R100 VTAIL.n182 VTAIL.n120 185
R101 VTAIL.n189 VTAIL.n119 185
R102 VTAIL.n191 VTAIL.n190 185
R103 VTAIL.n193 VTAIL.n192 185
R104 VTAIL.n116 VTAIL.n115 185
R105 VTAIL.n199 VTAIL.n198 185
R106 VTAIL.n201 VTAIL.n200 185
R107 VTAIL.n112 VTAIL.n111 185
R108 VTAIL.n207 VTAIL.n206 185
R109 VTAIL.n209 VTAIL.n208 185
R110 VTAIL.n251 VTAIL.n250 185
R111 VTAIL.n248 VTAIL.n247 185
R112 VTAIL.n257 VTAIL.n256 185
R113 VTAIL.n259 VTAIL.n258 185
R114 VTAIL.n244 VTAIL.n243 185
R115 VTAIL.n265 VTAIL.n264 185
R116 VTAIL.n267 VTAIL.n266 185
R117 VTAIL.n240 VTAIL.n239 185
R118 VTAIL.n273 VTAIL.n272 185
R119 VTAIL.n275 VTAIL.n274 185
R120 VTAIL.n236 VTAIL.n235 185
R121 VTAIL.n281 VTAIL.n280 185
R122 VTAIL.n283 VTAIL.n282 185
R123 VTAIL.n232 VTAIL.n231 185
R124 VTAIL.n289 VTAIL.n288 185
R125 VTAIL.n292 VTAIL.n291 185
R126 VTAIL.n290 VTAIL.n228 185
R127 VTAIL.n297 VTAIL.n227 185
R128 VTAIL.n299 VTAIL.n298 185
R129 VTAIL.n301 VTAIL.n300 185
R130 VTAIL.n224 VTAIL.n223 185
R131 VTAIL.n307 VTAIL.n306 185
R132 VTAIL.n309 VTAIL.n308 185
R133 VTAIL.n220 VTAIL.n219 185
R134 VTAIL.n315 VTAIL.n314 185
R135 VTAIL.n317 VTAIL.n316 185
R136 VTAIL.n745 VTAIL.n744 185
R137 VTAIL.n743 VTAIL.n742 185
R138 VTAIL.n648 VTAIL.n647 185
R139 VTAIL.n737 VTAIL.n736 185
R140 VTAIL.n735 VTAIL.n734 185
R141 VTAIL.n652 VTAIL.n651 185
R142 VTAIL.n729 VTAIL.n728 185
R143 VTAIL.n727 VTAIL.n726 185
R144 VTAIL.n725 VTAIL.n655 185
R145 VTAIL.n659 VTAIL.n656 185
R146 VTAIL.n720 VTAIL.n719 185
R147 VTAIL.n718 VTAIL.n717 185
R148 VTAIL.n661 VTAIL.n660 185
R149 VTAIL.n712 VTAIL.n711 185
R150 VTAIL.n710 VTAIL.n709 185
R151 VTAIL.n665 VTAIL.n664 185
R152 VTAIL.n704 VTAIL.n703 185
R153 VTAIL.n702 VTAIL.n701 185
R154 VTAIL.n669 VTAIL.n668 185
R155 VTAIL.n696 VTAIL.n695 185
R156 VTAIL.n694 VTAIL.n693 185
R157 VTAIL.n673 VTAIL.n672 185
R158 VTAIL.n688 VTAIL.n687 185
R159 VTAIL.n686 VTAIL.n685 185
R160 VTAIL.n677 VTAIL.n676 185
R161 VTAIL.n680 VTAIL.n679 185
R162 VTAIL.n637 VTAIL.n636 185
R163 VTAIL.n635 VTAIL.n634 185
R164 VTAIL.n540 VTAIL.n539 185
R165 VTAIL.n629 VTAIL.n628 185
R166 VTAIL.n627 VTAIL.n626 185
R167 VTAIL.n544 VTAIL.n543 185
R168 VTAIL.n621 VTAIL.n620 185
R169 VTAIL.n619 VTAIL.n618 185
R170 VTAIL.n617 VTAIL.n547 185
R171 VTAIL.n551 VTAIL.n548 185
R172 VTAIL.n612 VTAIL.n611 185
R173 VTAIL.n610 VTAIL.n609 185
R174 VTAIL.n553 VTAIL.n552 185
R175 VTAIL.n604 VTAIL.n603 185
R176 VTAIL.n602 VTAIL.n601 185
R177 VTAIL.n557 VTAIL.n556 185
R178 VTAIL.n596 VTAIL.n595 185
R179 VTAIL.n594 VTAIL.n593 185
R180 VTAIL.n561 VTAIL.n560 185
R181 VTAIL.n588 VTAIL.n587 185
R182 VTAIL.n586 VTAIL.n585 185
R183 VTAIL.n565 VTAIL.n564 185
R184 VTAIL.n580 VTAIL.n579 185
R185 VTAIL.n578 VTAIL.n577 185
R186 VTAIL.n569 VTAIL.n568 185
R187 VTAIL.n572 VTAIL.n571 185
R188 VTAIL.n531 VTAIL.n530 185
R189 VTAIL.n529 VTAIL.n528 185
R190 VTAIL.n434 VTAIL.n433 185
R191 VTAIL.n523 VTAIL.n522 185
R192 VTAIL.n521 VTAIL.n520 185
R193 VTAIL.n438 VTAIL.n437 185
R194 VTAIL.n515 VTAIL.n514 185
R195 VTAIL.n513 VTAIL.n512 185
R196 VTAIL.n511 VTAIL.n441 185
R197 VTAIL.n445 VTAIL.n442 185
R198 VTAIL.n506 VTAIL.n505 185
R199 VTAIL.n504 VTAIL.n503 185
R200 VTAIL.n447 VTAIL.n446 185
R201 VTAIL.n498 VTAIL.n497 185
R202 VTAIL.n496 VTAIL.n495 185
R203 VTAIL.n451 VTAIL.n450 185
R204 VTAIL.n490 VTAIL.n489 185
R205 VTAIL.n488 VTAIL.n487 185
R206 VTAIL.n455 VTAIL.n454 185
R207 VTAIL.n482 VTAIL.n481 185
R208 VTAIL.n480 VTAIL.n479 185
R209 VTAIL.n459 VTAIL.n458 185
R210 VTAIL.n474 VTAIL.n473 185
R211 VTAIL.n472 VTAIL.n471 185
R212 VTAIL.n463 VTAIL.n462 185
R213 VTAIL.n466 VTAIL.n465 185
R214 VTAIL.n423 VTAIL.n422 185
R215 VTAIL.n421 VTAIL.n420 185
R216 VTAIL.n326 VTAIL.n325 185
R217 VTAIL.n415 VTAIL.n414 185
R218 VTAIL.n413 VTAIL.n412 185
R219 VTAIL.n330 VTAIL.n329 185
R220 VTAIL.n407 VTAIL.n406 185
R221 VTAIL.n405 VTAIL.n404 185
R222 VTAIL.n403 VTAIL.n333 185
R223 VTAIL.n337 VTAIL.n334 185
R224 VTAIL.n398 VTAIL.n397 185
R225 VTAIL.n396 VTAIL.n395 185
R226 VTAIL.n339 VTAIL.n338 185
R227 VTAIL.n390 VTAIL.n389 185
R228 VTAIL.n388 VTAIL.n387 185
R229 VTAIL.n343 VTAIL.n342 185
R230 VTAIL.n382 VTAIL.n381 185
R231 VTAIL.n380 VTAIL.n379 185
R232 VTAIL.n347 VTAIL.n346 185
R233 VTAIL.n374 VTAIL.n373 185
R234 VTAIL.n372 VTAIL.n371 185
R235 VTAIL.n351 VTAIL.n350 185
R236 VTAIL.n366 VTAIL.n365 185
R237 VTAIL.n364 VTAIL.n363 185
R238 VTAIL.n355 VTAIL.n354 185
R239 VTAIL.n358 VTAIL.n357 185
R240 VTAIL.t2 VTAIL.n678 147.659
R241 VTAIL.t0 VTAIL.n570 147.659
R242 VTAIL.t8 VTAIL.n464 147.659
R243 VTAIL.t14 VTAIL.n356 147.659
R244 VTAIL.t9 VTAIL.n783 147.659
R245 VTAIL.t10 VTAIL.n35 147.659
R246 VTAIL.t3 VTAIL.n141 147.659
R247 VTAIL.t7 VTAIL.n249 147.659
R248 VTAIL.n784 VTAIL.n781 104.615
R249 VTAIL.n791 VTAIL.n781 104.615
R250 VTAIL.n792 VTAIL.n791 104.615
R251 VTAIL.n792 VTAIL.n777 104.615
R252 VTAIL.n799 VTAIL.n777 104.615
R253 VTAIL.n800 VTAIL.n799 104.615
R254 VTAIL.n800 VTAIL.n773 104.615
R255 VTAIL.n807 VTAIL.n773 104.615
R256 VTAIL.n808 VTAIL.n807 104.615
R257 VTAIL.n808 VTAIL.n769 104.615
R258 VTAIL.n815 VTAIL.n769 104.615
R259 VTAIL.n816 VTAIL.n815 104.615
R260 VTAIL.n816 VTAIL.n765 104.615
R261 VTAIL.n823 VTAIL.n765 104.615
R262 VTAIL.n825 VTAIL.n823 104.615
R263 VTAIL.n825 VTAIL.n824 104.615
R264 VTAIL.n824 VTAIL.n761 104.615
R265 VTAIL.n833 VTAIL.n761 104.615
R266 VTAIL.n834 VTAIL.n833 104.615
R267 VTAIL.n834 VTAIL.n757 104.615
R268 VTAIL.n841 VTAIL.n757 104.615
R269 VTAIL.n842 VTAIL.n841 104.615
R270 VTAIL.n842 VTAIL.n753 104.615
R271 VTAIL.n849 VTAIL.n753 104.615
R272 VTAIL.n850 VTAIL.n849 104.615
R273 VTAIL.n36 VTAIL.n33 104.615
R274 VTAIL.n43 VTAIL.n33 104.615
R275 VTAIL.n44 VTAIL.n43 104.615
R276 VTAIL.n44 VTAIL.n29 104.615
R277 VTAIL.n51 VTAIL.n29 104.615
R278 VTAIL.n52 VTAIL.n51 104.615
R279 VTAIL.n52 VTAIL.n25 104.615
R280 VTAIL.n59 VTAIL.n25 104.615
R281 VTAIL.n60 VTAIL.n59 104.615
R282 VTAIL.n60 VTAIL.n21 104.615
R283 VTAIL.n67 VTAIL.n21 104.615
R284 VTAIL.n68 VTAIL.n67 104.615
R285 VTAIL.n68 VTAIL.n17 104.615
R286 VTAIL.n75 VTAIL.n17 104.615
R287 VTAIL.n77 VTAIL.n75 104.615
R288 VTAIL.n77 VTAIL.n76 104.615
R289 VTAIL.n76 VTAIL.n13 104.615
R290 VTAIL.n85 VTAIL.n13 104.615
R291 VTAIL.n86 VTAIL.n85 104.615
R292 VTAIL.n86 VTAIL.n9 104.615
R293 VTAIL.n93 VTAIL.n9 104.615
R294 VTAIL.n94 VTAIL.n93 104.615
R295 VTAIL.n94 VTAIL.n5 104.615
R296 VTAIL.n101 VTAIL.n5 104.615
R297 VTAIL.n102 VTAIL.n101 104.615
R298 VTAIL.n142 VTAIL.n139 104.615
R299 VTAIL.n149 VTAIL.n139 104.615
R300 VTAIL.n150 VTAIL.n149 104.615
R301 VTAIL.n150 VTAIL.n135 104.615
R302 VTAIL.n157 VTAIL.n135 104.615
R303 VTAIL.n158 VTAIL.n157 104.615
R304 VTAIL.n158 VTAIL.n131 104.615
R305 VTAIL.n165 VTAIL.n131 104.615
R306 VTAIL.n166 VTAIL.n165 104.615
R307 VTAIL.n166 VTAIL.n127 104.615
R308 VTAIL.n173 VTAIL.n127 104.615
R309 VTAIL.n174 VTAIL.n173 104.615
R310 VTAIL.n174 VTAIL.n123 104.615
R311 VTAIL.n181 VTAIL.n123 104.615
R312 VTAIL.n183 VTAIL.n181 104.615
R313 VTAIL.n183 VTAIL.n182 104.615
R314 VTAIL.n182 VTAIL.n119 104.615
R315 VTAIL.n191 VTAIL.n119 104.615
R316 VTAIL.n192 VTAIL.n191 104.615
R317 VTAIL.n192 VTAIL.n115 104.615
R318 VTAIL.n199 VTAIL.n115 104.615
R319 VTAIL.n200 VTAIL.n199 104.615
R320 VTAIL.n200 VTAIL.n111 104.615
R321 VTAIL.n207 VTAIL.n111 104.615
R322 VTAIL.n208 VTAIL.n207 104.615
R323 VTAIL.n250 VTAIL.n247 104.615
R324 VTAIL.n257 VTAIL.n247 104.615
R325 VTAIL.n258 VTAIL.n257 104.615
R326 VTAIL.n258 VTAIL.n243 104.615
R327 VTAIL.n265 VTAIL.n243 104.615
R328 VTAIL.n266 VTAIL.n265 104.615
R329 VTAIL.n266 VTAIL.n239 104.615
R330 VTAIL.n273 VTAIL.n239 104.615
R331 VTAIL.n274 VTAIL.n273 104.615
R332 VTAIL.n274 VTAIL.n235 104.615
R333 VTAIL.n281 VTAIL.n235 104.615
R334 VTAIL.n282 VTAIL.n281 104.615
R335 VTAIL.n282 VTAIL.n231 104.615
R336 VTAIL.n289 VTAIL.n231 104.615
R337 VTAIL.n291 VTAIL.n289 104.615
R338 VTAIL.n291 VTAIL.n290 104.615
R339 VTAIL.n290 VTAIL.n227 104.615
R340 VTAIL.n299 VTAIL.n227 104.615
R341 VTAIL.n300 VTAIL.n299 104.615
R342 VTAIL.n300 VTAIL.n223 104.615
R343 VTAIL.n307 VTAIL.n223 104.615
R344 VTAIL.n308 VTAIL.n307 104.615
R345 VTAIL.n308 VTAIL.n219 104.615
R346 VTAIL.n315 VTAIL.n219 104.615
R347 VTAIL.n316 VTAIL.n315 104.615
R348 VTAIL.n744 VTAIL.n743 104.615
R349 VTAIL.n743 VTAIL.n647 104.615
R350 VTAIL.n736 VTAIL.n647 104.615
R351 VTAIL.n736 VTAIL.n735 104.615
R352 VTAIL.n735 VTAIL.n651 104.615
R353 VTAIL.n728 VTAIL.n651 104.615
R354 VTAIL.n728 VTAIL.n727 104.615
R355 VTAIL.n727 VTAIL.n655 104.615
R356 VTAIL.n659 VTAIL.n655 104.615
R357 VTAIL.n719 VTAIL.n659 104.615
R358 VTAIL.n719 VTAIL.n718 104.615
R359 VTAIL.n718 VTAIL.n660 104.615
R360 VTAIL.n711 VTAIL.n660 104.615
R361 VTAIL.n711 VTAIL.n710 104.615
R362 VTAIL.n710 VTAIL.n664 104.615
R363 VTAIL.n703 VTAIL.n664 104.615
R364 VTAIL.n703 VTAIL.n702 104.615
R365 VTAIL.n702 VTAIL.n668 104.615
R366 VTAIL.n695 VTAIL.n668 104.615
R367 VTAIL.n695 VTAIL.n694 104.615
R368 VTAIL.n694 VTAIL.n672 104.615
R369 VTAIL.n687 VTAIL.n672 104.615
R370 VTAIL.n687 VTAIL.n686 104.615
R371 VTAIL.n686 VTAIL.n676 104.615
R372 VTAIL.n679 VTAIL.n676 104.615
R373 VTAIL.n636 VTAIL.n635 104.615
R374 VTAIL.n635 VTAIL.n539 104.615
R375 VTAIL.n628 VTAIL.n539 104.615
R376 VTAIL.n628 VTAIL.n627 104.615
R377 VTAIL.n627 VTAIL.n543 104.615
R378 VTAIL.n620 VTAIL.n543 104.615
R379 VTAIL.n620 VTAIL.n619 104.615
R380 VTAIL.n619 VTAIL.n547 104.615
R381 VTAIL.n551 VTAIL.n547 104.615
R382 VTAIL.n611 VTAIL.n551 104.615
R383 VTAIL.n611 VTAIL.n610 104.615
R384 VTAIL.n610 VTAIL.n552 104.615
R385 VTAIL.n603 VTAIL.n552 104.615
R386 VTAIL.n603 VTAIL.n602 104.615
R387 VTAIL.n602 VTAIL.n556 104.615
R388 VTAIL.n595 VTAIL.n556 104.615
R389 VTAIL.n595 VTAIL.n594 104.615
R390 VTAIL.n594 VTAIL.n560 104.615
R391 VTAIL.n587 VTAIL.n560 104.615
R392 VTAIL.n587 VTAIL.n586 104.615
R393 VTAIL.n586 VTAIL.n564 104.615
R394 VTAIL.n579 VTAIL.n564 104.615
R395 VTAIL.n579 VTAIL.n578 104.615
R396 VTAIL.n578 VTAIL.n568 104.615
R397 VTAIL.n571 VTAIL.n568 104.615
R398 VTAIL.n530 VTAIL.n529 104.615
R399 VTAIL.n529 VTAIL.n433 104.615
R400 VTAIL.n522 VTAIL.n433 104.615
R401 VTAIL.n522 VTAIL.n521 104.615
R402 VTAIL.n521 VTAIL.n437 104.615
R403 VTAIL.n514 VTAIL.n437 104.615
R404 VTAIL.n514 VTAIL.n513 104.615
R405 VTAIL.n513 VTAIL.n441 104.615
R406 VTAIL.n445 VTAIL.n441 104.615
R407 VTAIL.n505 VTAIL.n445 104.615
R408 VTAIL.n505 VTAIL.n504 104.615
R409 VTAIL.n504 VTAIL.n446 104.615
R410 VTAIL.n497 VTAIL.n446 104.615
R411 VTAIL.n497 VTAIL.n496 104.615
R412 VTAIL.n496 VTAIL.n450 104.615
R413 VTAIL.n489 VTAIL.n450 104.615
R414 VTAIL.n489 VTAIL.n488 104.615
R415 VTAIL.n488 VTAIL.n454 104.615
R416 VTAIL.n481 VTAIL.n454 104.615
R417 VTAIL.n481 VTAIL.n480 104.615
R418 VTAIL.n480 VTAIL.n458 104.615
R419 VTAIL.n473 VTAIL.n458 104.615
R420 VTAIL.n473 VTAIL.n472 104.615
R421 VTAIL.n472 VTAIL.n462 104.615
R422 VTAIL.n465 VTAIL.n462 104.615
R423 VTAIL.n422 VTAIL.n421 104.615
R424 VTAIL.n421 VTAIL.n325 104.615
R425 VTAIL.n414 VTAIL.n325 104.615
R426 VTAIL.n414 VTAIL.n413 104.615
R427 VTAIL.n413 VTAIL.n329 104.615
R428 VTAIL.n406 VTAIL.n329 104.615
R429 VTAIL.n406 VTAIL.n405 104.615
R430 VTAIL.n405 VTAIL.n333 104.615
R431 VTAIL.n337 VTAIL.n333 104.615
R432 VTAIL.n397 VTAIL.n337 104.615
R433 VTAIL.n397 VTAIL.n396 104.615
R434 VTAIL.n396 VTAIL.n338 104.615
R435 VTAIL.n389 VTAIL.n338 104.615
R436 VTAIL.n389 VTAIL.n388 104.615
R437 VTAIL.n388 VTAIL.n342 104.615
R438 VTAIL.n381 VTAIL.n342 104.615
R439 VTAIL.n381 VTAIL.n380 104.615
R440 VTAIL.n380 VTAIL.n346 104.615
R441 VTAIL.n373 VTAIL.n346 104.615
R442 VTAIL.n373 VTAIL.n372 104.615
R443 VTAIL.n372 VTAIL.n350 104.615
R444 VTAIL.n365 VTAIL.n350 104.615
R445 VTAIL.n365 VTAIL.n364 104.615
R446 VTAIL.n364 VTAIL.n354 104.615
R447 VTAIL.n357 VTAIL.n354 104.615
R448 VTAIL.n784 VTAIL.t9 52.3082
R449 VTAIL.n36 VTAIL.t10 52.3082
R450 VTAIL.n142 VTAIL.t3 52.3082
R451 VTAIL.n250 VTAIL.t7 52.3082
R452 VTAIL.n679 VTAIL.t2 52.3082
R453 VTAIL.n571 VTAIL.t0 52.3082
R454 VTAIL.n465 VTAIL.t8 52.3082
R455 VTAIL.n357 VTAIL.t14 52.3082
R456 VTAIL.n1 VTAIL.n0 43.1674
R457 VTAIL.n215 VTAIL.n214 43.1674
R458 VTAIL.n643 VTAIL.n642 43.1674
R459 VTAIL.n429 VTAIL.n428 43.1674
R460 VTAIL.n855 VTAIL.n854 31.4096
R461 VTAIL.n107 VTAIL.n106 31.4096
R462 VTAIL.n213 VTAIL.n212 31.4096
R463 VTAIL.n321 VTAIL.n320 31.4096
R464 VTAIL.n749 VTAIL.n748 31.4096
R465 VTAIL.n641 VTAIL.n640 31.4096
R466 VTAIL.n535 VTAIL.n534 31.4096
R467 VTAIL.n427 VTAIL.n426 31.4096
R468 VTAIL.n855 VTAIL.n749 29.2548
R469 VTAIL.n427 VTAIL.n321 29.2548
R470 VTAIL.n785 VTAIL.n783 15.6677
R471 VTAIL.n37 VTAIL.n35 15.6677
R472 VTAIL.n143 VTAIL.n141 15.6677
R473 VTAIL.n251 VTAIL.n249 15.6677
R474 VTAIL.n680 VTAIL.n678 15.6677
R475 VTAIL.n572 VTAIL.n570 15.6677
R476 VTAIL.n466 VTAIL.n464 15.6677
R477 VTAIL.n358 VTAIL.n356 15.6677
R478 VTAIL.n832 VTAIL.n831 13.1884
R479 VTAIL.n84 VTAIL.n83 13.1884
R480 VTAIL.n190 VTAIL.n189 13.1884
R481 VTAIL.n298 VTAIL.n297 13.1884
R482 VTAIL.n726 VTAIL.n725 13.1884
R483 VTAIL.n618 VTAIL.n617 13.1884
R484 VTAIL.n512 VTAIL.n511 13.1884
R485 VTAIL.n404 VTAIL.n403 13.1884
R486 VTAIL.n786 VTAIL.n782 12.8005
R487 VTAIL.n830 VTAIL.n762 12.8005
R488 VTAIL.n835 VTAIL.n760 12.8005
R489 VTAIL.n38 VTAIL.n34 12.8005
R490 VTAIL.n82 VTAIL.n14 12.8005
R491 VTAIL.n87 VTAIL.n12 12.8005
R492 VTAIL.n144 VTAIL.n140 12.8005
R493 VTAIL.n188 VTAIL.n120 12.8005
R494 VTAIL.n193 VTAIL.n118 12.8005
R495 VTAIL.n252 VTAIL.n248 12.8005
R496 VTAIL.n296 VTAIL.n228 12.8005
R497 VTAIL.n301 VTAIL.n226 12.8005
R498 VTAIL.n729 VTAIL.n654 12.8005
R499 VTAIL.n724 VTAIL.n656 12.8005
R500 VTAIL.n681 VTAIL.n677 12.8005
R501 VTAIL.n621 VTAIL.n546 12.8005
R502 VTAIL.n616 VTAIL.n548 12.8005
R503 VTAIL.n573 VTAIL.n569 12.8005
R504 VTAIL.n515 VTAIL.n440 12.8005
R505 VTAIL.n510 VTAIL.n442 12.8005
R506 VTAIL.n467 VTAIL.n463 12.8005
R507 VTAIL.n407 VTAIL.n332 12.8005
R508 VTAIL.n402 VTAIL.n334 12.8005
R509 VTAIL.n359 VTAIL.n355 12.8005
R510 VTAIL.n790 VTAIL.n789 12.0247
R511 VTAIL.n827 VTAIL.n826 12.0247
R512 VTAIL.n836 VTAIL.n758 12.0247
R513 VTAIL.n42 VTAIL.n41 12.0247
R514 VTAIL.n79 VTAIL.n78 12.0247
R515 VTAIL.n88 VTAIL.n10 12.0247
R516 VTAIL.n148 VTAIL.n147 12.0247
R517 VTAIL.n185 VTAIL.n184 12.0247
R518 VTAIL.n194 VTAIL.n116 12.0247
R519 VTAIL.n256 VTAIL.n255 12.0247
R520 VTAIL.n293 VTAIL.n292 12.0247
R521 VTAIL.n302 VTAIL.n224 12.0247
R522 VTAIL.n730 VTAIL.n652 12.0247
R523 VTAIL.n721 VTAIL.n720 12.0247
R524 VTAIL.n685 VTAIL.n684 12.0247
R525 VTAIL.n622 VTAIL.n544 12.0247
R526 VTAIL.n613 VTAIL.n612 12.0247
R527 VTAIL.n577 VTAIL.n576 12.0247
R528 VTAIL.n516 VTAIL.n438 12.0247
R529 VTAIL.n507 VTAIL.n506 12.0247
R530 VTAIL.n471 VTAIL.n470 12.0247
R531 VTAIL.n408 VTAIL.n330 12.0247
R532 VTAIL.n399 VTAIL.n398 12.0247
R533 VTAIL.n363 VTAIL.n362 12.0247
R534 VTAIL.n793 VTAIL.n780 11.249
R535 VTAIL.n822 VTAIL.n764 11.249
R536 VTAIL.n840 VTAIL.n839 11.249
R537 VTAIL.n45 VTAIL.n32 11.249
R538 VTAIL.n74 VTAIL.n16 11.249
R539 VTAIL.n92 VTAIL.n91 11.249
R540 VTAIL.n151 VTAIL.n138 11.249
R541 VTAIL.n180 VTAIL.n122 11.249
R542 VTAIL.n198 VTAIL.n197 11.249
R543 VTAIL.n259 VTAIL.n246 11.249
R544 VTAIL.n288 VTAIL.n230 11.249
R545 VTAIL.n306 VTAIL.n305 11.249
R546 VTAIL.n734 VTAIL.n733 11.249
R547 VTAIL.n717 VTAIL.n658 11.249
R548 VTAIL.n688 VTAIL.n675 11.249
R549 VTAIL.n626 VTAIL.n625 11.249
R550 VTAIL.n609 VTAIL.n550 11.249
R551 VTAIL.n580 VTAIL.n567 11.249
R552 VTAIL.n520 VTAIL.n519 11.249
R553 VTAIL.n503 VTAIL.n444 11.249
R554 VTAIL.n474 VTAIL.n461 11.249
R555 VTAIL.n412 VTAIL.n411 11.249
R556 VTAIL.n395 VTAIL.n336 11.249
R557 VTAIL.n366 VTAIL.n353 11.249
R558 VTAIL.n794 VTAIL.n778 10.4732
R559 VTAIL.n821 VTAIL.n766 10.4732
R560 VTAIL.n843 VTAIL.n756 10.4732
R561 VTAIL.n46 VTAIL.n30 10.4732
R562 VTAIL.n73 VTAIL.n18 10.4732
R563 VTAIL.n95 VTAIL.n8 10.4732
R564 VTAIL.n152 VTAIL.n136 10.4732
R565 VTAIL.n179 VTAIL.n124 10.4732
R566 VTAIL.n201 VTAIL.n114 10.4732
R567 VTAIL.n260 VTAIL.n244 10.4732
R568 VTAIL.n287 VTAIL.n232 10.4732
R569 VTAIL.n309 VTAIL.n222 10.4732
R570 VTAIL.n737 VTAIL.n650 10.4732
R571 VTAIL.n716 VTAIL.n661 10.4732
R572 VTAIL.n689 VTAIL.n673 10.4732
R573 VTAIL.n629 VTAIL.n542 10.4732
R574 VTAIL.n608 VTAIL.n553 10.4732
R575 VTAIL.n581 VTAIL.n565 10.4732
R576 VTAIL.n523 VTAIL.n436 10.4732
R577 VTAIL.n502 VTAIL.n447 10.4732
R578 VTAIL.n475 VTAIL.n459 10.4732
R579 VTAIL.n415 VTAIL.n328 10.4732
R580 VTAIL.n394 VTAIL.n339 10.4732
R581 VTAIL.n367 VTAIL.n351 10.4732
R582 VTAIL.n798 VTAIL.n797 9.69747
R583 VTAIL.n818 VTAIL.n817 9.69747
R584 VTAIL.n844 VTAIL.n754 9.69747
R585 VTAIL.n50 VTAIL.n49 9.69747
R586 VTAIL.n70 VTAIL.n69 9.69747
R587 VTAIL.n96 VTAIL.n6 9.69747
R588 VTAIL.n156 VTAIL.n155 9.69747
R589 VTAIL.n176 VTAIL.n175 9.69747
R590 VTAIL.n202 VTAIL.n112 9.69747
R591 VTAIL.n264 VTAIL.n263 9.69747
R592 VTAIL.n284 VTAIL.n283 9.69747
R593 VTAIL.n310 VTAIL.n220 9.69747
R594 VTAIL.n738 VTAIL.n648 9.69747
R595 VTAIL.n713 VTAIL.n712 9.69747
R596 VTAIL.n693 VTAIL.n692 9.69747
R597 VTAIL.n630 VTAIL.n540 9.69747
R598 VTAIL.n605 VTAIL.n604 9.69747
R599 VTAIL.n585 VTAIL.n584 9.69747
R600 VTAIL.n524 VTAIL.n434 9.69747
R601 VTAIL.n499 VTAIL.n498 9.69747
R602 VTAIL.n479 VTAIL.n478 9.69747
R603 VTAIL.n416 VTAIL.n326 9.69747
R604 VTAIL.n391 VTAIL.n390 9.69747
R605 VTAIL.n371 VTAIL.n370 9.69747
R606 VTAIL.n854 VTAIL.n853 9.45567
R607 VTAIL.n106 VTAIL.n105 9.45567
R608 VTAIL.n212 VTAIL.n211 9.45567
R609 VTAIL.n320 VTAIL.n319 9.45567
R610 VTAIL.n748 VTAIL.n747 9.45567
R611 VTAIL.n640 VTAIL.n639 9.45567
R612 VTAIL.n534 VTAIL.n533 9.45567
R613 VTAIL.n426 VTAIL.n425 9.45567
R614 VTAIL.n752 VTAIL.n751 9.3005
R615 VTAIL.n847 VTAIL.n846 9.3005
R616 VTAIL.n845 VTAIL.n844 9.3005
R617 VTAIL.n756 VTAIL.n755 9.3005
R618 VTAIL.n839 VTAIL.n838 9.3005
R619 VTAIL.n837 VTAIL.n836 9.3005
R620 VTAIL.n760 VTAIL.n759 9.3005
R621 VTAIL.n805 VTAIL.n804 9.3005
R622 VTAIL.n803 VTAIL.n802 9.3005
R623 VTAIL.n776 VTAIL.n775 9.3005
R624 VTAIL.n797 VTAIL.n796 9.3005
R625 VTAIL.n795 VTAIL.n794 9.3005
R626 VTAIL.n780 VTAIL.n779 9.3005
R627 VTAIL.n789 VTAIL.n788 9.3005
R628 VTAIL.n787 VTAIL.n786 9.3005
R629 VTAIL.n772 VTAIL.n771 9.3005
R630 VTAIL.n811 VTAIL.n810 9.3005
R631 VTAIL.n813 VTAIL.n812 9.3005
R632 VTAIL.n768 VTAIL.n767 9.3005
R633 VTAIL.n819 VTAIL.n818 9.3005
R634 VTAIL.n821 VTAIL.n820 9.3005
R635 VTAIL.n764 VTAIL.n763 9.3005
R636 VTAIL.n828 VTAIL.n827 9.3005
R637 VTAIL.n830 VTAIL.n829 9.3005
R638 VTAIL.n853 VTAIL.n852 9.3005
R639 VTAIL.n4 VTAIL.n3 9.3005
R640 VTAIL.n99 VTAIL.n98 9.3005
R641 VTAIL.n97 VTAIL.n96 9.3005
R642 VTAIL.n8 VTAIL.n7 9.3005
R643 VTAIL.n91 VTAIL.n90 9.3005
R644 VTAIL.n89 VTAIL.n88 9.3005
R645 VTAIL.n12 VTAIL.n11 9.3005
R646 VTAIL.n57 VTAIL.n56 9.3005
R647 VTAIL.n55 VTAIL.n54 9.3005
R648 VTAIL.n28 VTAIL.n27 9.3005
R649 VTAIL.n49 VTAIL.n48 9.3005
R650 VTAIL.n47 VTAIL.n46 9.3005
R651 VTAIL.n32 VTAIL.n31 9.3005
R652 VTAIL.n41 VTAIL.n40 9.3005
R653 VTAIL.n39 VTAIL.n38 9.3005
R654 VTAIL.n24 VTAIL.n23 9.3005
R655 VTAIL.n63 VTAIL.n62 9.3005
R656 VTAIL.n65 VTAIL.n64 9.3005
R657 VTAIL.n20 VTAIL.n19 9.3005
R658 VTAIL.n71 VTAIL.n70 9.3005
R659 VTAIL.n73 VTAIL.n72 9.3005
R660 VTAIL.n16 VTAIL.n15 9.3005
R661 VTAIL.n80 VTAIL.n79 9.3005
R662 VTAIL.n82 VTAIL.n81 9.3005
R663 VTAIL.n105 VTAIL.n104 9.3005
R664 VTAIL.n110 VTAIL.n109 9.3005
R665 VTAIL.n205 VTAIL.n204 9.3005
R666 VTAIL.n203 VTAIL.n202 9.3005
R667 VTAIL.n114 VTAIL.n113 9.3005
R668 VTAIL.n197 VTAIL.n196 9.3005
R669 VTAIL.n195 VTAIL.n194 9.3005
R670 VTAIL.n118 VTAIL.n117 9.3005
R671 VTAIL.n163 VTAIL.n162 9.3005
R672 VTAIL.n161 VTAIL.n160 9.3005
R673 VTAIL.n134 VTAIL.n133 9.3005
R674 VTAIL.n155 VTAIL.n154 9.3005
R675 VTAIL.n153 VTAIL.n152 9.3005
R676 VTAIL.n138 VTAIL.n137 9.3005
R677 VTAIL.n147 VTAIL.n146 9.3005
R678 VTAIL.n145 VTAIL.n144 9.3005
R679 VTAIL.n130 VTAIL.n129 9.3005
R680 VTAIL.n169 VTAIL.n168 9.3005
R681 VTAIL.n171 VTAIL.n170 9.3005
R682 VTAIL.n126 VTAIL.n125 9.3005
R683 VTAIL.n177 VTAIL.n176 9.3005
R684 VTAIL.n179 VTAIL.n178 9.3005
R685 VTAIL.n122 VTAIL.n121 9.3005
R686 VTAIL.n186 VTAIL.n185 9.3005
R687 VTAIL.n188 VTAIL.n187 9.3005
R688 VTAIL.n211 VTAIL.n210 9.3005
R689 VTAIL.n218 VTAIL.n217 9.3005
R690 VTAIL.n313 VTAIL.n312 9.3005
R691 VTAIL.n311 VTAIL.n310 9.3005
R692 VTAIL.n222 VTAIL.n221 9.3005
R693 VTAIL.n305 VTAIL.n304 9.3005
R694 VTAIL.n303 VTAIL.n302 9.3005
R695 VTAIL.n226 VTAIL.n225 9.3005
R696 VTAIL.n271 VTAIL.n270 9.3005
R697 VTAIL.n269 VTAIL.n268 9.3005
R698 VTAIL.n242 VTAIL.n241 9.3005
R699 VTAIL.n263 VTAIL.n262 9.3005
R700 VTAIL.n261 VTAIL.n260 9.3005
R701 VTAIL.n246 VTAIL.n245 9.3005
R702 VTAIL.n255 VTAIL.n254 9.3005
R703 VTAIL.n253 VTAIL.n252 9.3005
R704 VTAIL.n238 VTAIL.n237 9.3005
R705 VTAIL.n277 VTAIL.n276 9.3005
R706 VTAIL.n279 VTAIL.n278 9.3005
R707 VTAIL.n234 VTAIL.n233 9.3005
R708 VTAIL.n285 VTAIL.n284 9.3005
R709 VTAIL.n287 VTAIL.n286 9.3005
R710 VTAIL.n230 VTAIL.n229 9.3005
R711 VTAIL.n294 VTAIL.n293 9.3005
R712 VTAIL.n296 VTAIL.n295 9.3005
R713 VTAIL.n319 VTAIL.n318 9.3005
R714 VTAIL.n706 VTAIL.n705 9.3005
R715 VTAIL.n708 VTAIL.n707 9.3005
R716 VTAIL.n663 VTAIL.n662 9.3005
R717 VTAIL.n714 VTAIL.n713 9.3005
R718 VTAIL.n716 VTAIL.n715 9.3005
R719 VTAIL.n658 VTAIL.n657 9.3005
R720 VTAIL.n722 VTAIL.n721 9.3005
R721 VTAIL.n724 VTAIL.n723 9.3005
R722 VTAIL.n747 VTAIL.n746 9.3005
R723 VTAIL.n646 VTAIL.n645 9.3005
R724 VTAIL.n741 VTAIL.n740 9.3005
R725 VTAIL.n739 VTAIL.n738 9.3005
R726 VTAIL.n650 VTAIL.n649 9.3005
R727 VTAIL.n733 VTAIL.n732 9.3005
R728 VTAIL.n731 VTAIL.n730 9.3005
R729 VTAIL.n654 VTAIL.n653 9.3005
R730 VTAIL.n667 VTAIL.n666 9.3005
R731 VTAIL.n700 VTAIL.n699 9.3005
R732 VTAIL.n698 VTAIL.n697 9.3005
R733 VTAIL.n671 VTAIL.n670 9.3005
R734 VTAIL.n692 VTAIL.n691 9.3005
R735 VTAIL.n690 VTAIL.n689 9.3005
R736 VTAIL.n675 VTAIL.n674 9.3005
R737 VTAIL.n684 VTAIL.n683 9.3005
R738 VTAIL.n682 VTAIL.n681 9.3005
R739 VTAIL.n598 VTAIL.n597 9.3005
R740 VTAIL.n600 VTAIL.n599 9.3005
R741 VTAIL.n555 VTAIL.n554 9.3005
R742 VTAIL.n606 VTAIL.n605 9.3005
R743 VTAIL.n608 VTAIL.n607 9.3005
R744 VTAIL.n550 VTAIL.n549 9.3005
R745 VTAIL.n614 VTAIL.n613 9.3005
R746 VTAIL.n616 VTAIL.n615 9.3005
R747 VTAIL.n639 VTAIL.n638 9.3005
R748 VTAIL.n538 VTAIL.n537 9.3005
R749 VTAIL.n633 VTAIL.n632 9.3005
R750 VTAIL.n631 VTAIL.n630 9.3005
R751 VTAIL.n542 VTAIL.n541 9.3005
R752 VTAIL.n625 VTAIL.n624 9.3005
R753 VTAIL.n623 VTAIL.n622 9.3005
R754 VTAIL.n546 VTAIL.n545 9.3005
R755 VTAIL.n559 VTAIL.n558 9.3005
R756 VTAIL.n592 VTAIL.n591 9.3005
R757 VTAIL.n590 VTAIL.n589 9.3005
R758 VTAIL.n563 VTAIL.n562 9.3005
R759 VTAIL.n584 VTAIL.n583 9.3005
R760 VTAIL.n582 VTAIL.n581 9.3005
R761 VTAIL.n567 VTAIL.n566 9.3005
R762 VTAIL.n576 VTAIL.n575 9.3005
R763 VTAIL.n574 VTAIL.n573 9.3005
R764 VTAIL.n492 VTAIL.n491 9.3005
R765 VTAIL.n494 VTAIL.n493 9.3005
R766 VTAIL.n449 VTAIL.n448 9.3005
R767 VTAIL.n500 VTAIL.n499 9.3005
R768 VTAIL.n502 VTAIL.n501 9.3005
R769 VTAIL.n444 VTAIL.n443 9.3005
R770 VTAIL.n508 VTAIL.n507 9.3005
R771 VTAIL.n510 VTAIL.n509 9.3005
R772 VTAIL.n533 VTAIL.n532 9.3005
R773 VTAIL.n432 VTAIL.n431 9.3005
R774 VTAIL.n527 VTAIL.n526 9.3005
R775 VTAIL.n525 VTAIL.n524 9.3005
R776 VTAIL.n436 VTAIL.n435 9.3005
R777 VTAIL.n519 VTAIL.n518 9.3005
R778 VTAIL.n517 VTAIL.n516 9.3005
R779 VTAIL.n440 VTAIL.n439 9.3005
R780 VTAIL.n453 VTAIL.n452 9.3005
R781 VTAIL.n486 VTAIL.n485 9.3005
R782 VTAIL.n484 VTAIL.n483 9.3005
R783 VTAIL.n457 VTAIL.n456 9.3005
R784 VTAIL.n478 VTAIL.n477 9.3005
R785 VTAIL.n476 VTAIL.n475 9.3005
R786 VTAIL.n461 VTAIL.n460 9.3005
R787 VTAIL.n470 VTAIL.n469 9.3005
R788 VTAIL.n468 VTAIL.n467 9.3005
R789 VTAIL.n384 VTAIL.n383 9.3005
R790 VTAIL.n386 VTAIL.n385 9.3005
R791 VTAIL.n341 VTAIL.n340 9.3005
R792 VTAIL.n392 VTAIL.n391 9.3005
R793 VTAIL.n394 VTAIL.n393 9.3005
R794 VTAIL.n336 VTAIL.n335 9.3005
R795 VTAIL.n400 VTAIL.n399 9.3005
R796 VTAIL.n402 VTAIL.n401 9.3005
R797 VTAIL.n425 VTAIL.n424 9.3005
R798 VTAIL.n324 VTAIL.n323 9.3005
R799 VTAIL.n419 VTAIL.n418 9.3005
R800 VTAIL.n417 VTAIL.n416 9.3005
R801 VTAIL.n328 VTAIL.n327 9.3005
R802 VTAIL.n411 VTAIL.n410 9.3005
R803 VTAIL.n409 VTAIL.n408 9.3005
R804 VTAIL.n332 VTAIL.n331 9.3005
R805 VTAIL.n345 VTAIL.n344 9.3005
R806 VTAIL.n378 VTAIL.n377 9.3005
R807 VTAIL.n376 VTAIL.n375 9.3005
R808 VTAIL.n349 VTAIL.n348 9.3005
R809 VTAIL.n370 VTAIL.n369 9.3005
R810 VTAIL.n368 VTAIL.n367 9.3005
R811 VTAIL.n353 VTAIL.n352 9.3005
R812 VTAIL.n362 VTAIL.n361 9.3005
R813 VTAIL.n360 VTAIL.n359 9.3005
R814 VTAIL.n801 VTAIL.n776 8.92171
R815 VTAIL.n814 VTAIL.n768 8.92171
R816 VTAIL.n848 VTAIL.n847 8.92171
R817 VTAIL.n53 VTAIL.n28 8.92171
R818 VTAIL.n66 VTAIL.n20 8.92171
R819 VTAIL.n100 VTAIL.n99 8.92171
R820 VTAIL.n159 VTAIL.n134 8.92171
R821 VTAIL.n172 VTAIL.n126 8.92171
R822 VTAIL.n206 VTAIL.n205 8.92171
R823 VTAIL.n267 VTAIL.n242 8.92171
R824 VTAIL.n280 VTAIL.n234 8.92171
R825 VTAIL.n314 VTAIL.n313 8.92171
R826 VTAIL.n742 VTAIL.n741 8.92171
R827 VTAIL.n709 VTAIL.n663 8.92171
R828 VTAIL.n696 VTAIL.n671 8.92171
R829 VTAIL.n634 VTAIL.n633 8.92171
R830 VTAIL.n601 VTAIL.n555 8.92171
R831 VTAIL.n588 VTAIL.n563 8.92171
R832 VTAIL.n528 VTAIL.n527 8.92171
R833 VTAIL.n495 VTAIL.n449 8.92171
R834 VTAIL.n482 VTAIL.n457 8.92171
R835 VTAIL.n420 VTAIL.n419 8.92171
R836 VTAIL.n387 VTAIL.n341 8.92171
R837 VTAIL.n374 VTAIL.n349 8.92171
R838 VTAIL.n802 VTAIL.n774 8.14595
R839 VTAIL.n813 VTAIL.n770 8.14595
R840 VTAIL.n851 VTAIL.n752 8.14595
R841 VTAIL.n54 VTAIL.n26 8.14595
R842 VTAIL.n65 VTAIL.n22 8.14595
R843 VTAIL.n103 VTAIL.n4 8.14595
R844 VTAIL.n160 VTAIL.n132 8.14595
R845 VTAIL.n171 VTAIL.n128 8.14595
R846 VTAIL.n209 VTAIL.n110 8.14595
R847 VTAIL.n268 VTAIL.n240 8.14595
R848 VTAIL.n279 VTAIL.n236 8.14595
R849 VTAIL.n317 VTAIL.n218 8.14595
R850 VTAIL.n745 VTAIL.n646 8.14595
R851 VTAIL.n708 VTAIL.n665 8.14595
R852 VTAIL.n697 VTAIL.n669 8.14595
R853 VTAIL.n637 VTAIL.n538 8.14595
R854 VTAIL.n600 VTAIL.n557 8.14595
R855 VTAIL.n589 VTAIL.n561 8.14595
R856 VTAIL.n531 VTAIL.n432 8.14595
R857 VTAIL.n494 VTAIL.n451 8.14595
R858 VTAIL.n483 VTAIL.n455 8.14595
R859 VTAIL.n423 VTAIL.n324 8.14595
R860 VTAIL.n386 VTAIL.n343 8.14595
R861 VTAIL.n375 VTAIL.n347 8.14595
R862 VTAIL.n806 VTAIL.n805 7.3702
R863 VTAIL.n810 VTAIL.n809 7.3702
R864 VTAIL.n852 VTAIL.n750 7.3702
R865 VTAIL.n58 VTAIL.n57 7.3702
R866 VTAIL.n62 VTAIL.n61 7.3702
R867 VTAIL.n104 VTAIL.n2 7.3702
R868 VTAIL.n164 VTAIL.n163 7.3702
R869 VTAIL.n168 VTAIL.n167 7.3702
R870 VTAIL.n210 VTAIL.n108 7.3702
R871 VTAIL.n272 VTAIL.n271 7.3702
R872 VTAIL.n276 VTAIL.n275 7.3702
R873 VTAIL.n318 VTAIL.n216 7.3702
R874 VTAIL.n746 VTAIL.n644 7.3702
R875 VTAIL.n705 VTAIL.n704 7.3702
R876 VTAIL.n701 VTAIL.n700 7.3702
R877 VTAIL.n638 VTAIL.n536 7.3702
R878 VTAIL.n597 VTAIL.n596 7.3702
R879 VTAIL.n593 VTAIL.n592 7.3702
R880 VTAIL.n532 VTAIL.n430 7.3702
R881 VTAIL.n491 VTAIL.n490 7.3702
R882 VTAIL.n487 VTAIL.n486 7.3702
R883 VTAIL.n424 VTAIL.n322 7.3702
R884 VTAIL.n383 VTAIL.n382 7.3702
R885 VTAIL.n379 VTAIL.n378 7.3702
R886 VTAIL.n806 VTAIL.n772 6.59444
R887 VTAIL.n809 VTAIL.n772 6.59444
R888 VTAIL.n854 VTAIL.n750 6.59444
R889 VTAIL.n58 VTAIL.n24 6.59444
R890 VTAIL.n61 VTAIL.n24 6.59444
R891 VTAIL.n106 VTAIL.n2 6.59444
R892 VTAIL.n164 VTAIL.n130 6.59444
R893 VTAIL.n167 VTAIL.n130 6.59444
R894 VTAIL.n212 VTAIL.n108 6.59444
R895 VTAIL.n272 VTAIL.n238 6.59444
R896 VTAIL.n275 VTAIL.n238 6.59444
R897 VTAIL.n320 VTAIL.n216 6.59444
R898 VTAIL.n748 VTAIL.n644 6.59444
R899 VTAIL.n704 VTAIL.n667 6.59444
R900 VTAIL.n701 VTAIL.n667 6.59444
R901 VTAIL.n640 VTAIL.n536 6.59444
R902 VTAIL.n596 VTAIL.n559 6.59444
R903 VTAIL.n593 VTAIL.n559 6.59444
R904 VTAIL.n534 VTAIL.n430 6.59444
R905 VTAIL.n490 VTAIL.n453 6.59444
R906 VTAIL.n487 VTAIL.n453 6.59444
R907 VTAIL.n426 VTAIL.n322 6.59444
R908 VTAIL.n382 VTAIL.n345 6.59444
R909 VTAIL.n379 VTAIL.n345 6.59444
R910 VTAIL.n805 VTAIL.n774 5.81868
R911 VTAIL.n810 VTAIL.n770 5.81868
R912 VTAIL.n852 VTAIL.n851 5.81868
R913 VTAIL.n57 VTAIL.n26 5.81868
R914 VTAIL.n62 VTAIL.n22 5.81868
R915 VTAIL.n104 VTAIL.n103 5.81868
R916 VTAIL.n163 VTAIL.n132 5.81868
R917 VTAIL.n168 VTAIL.n128 5.81868
R918 VTAIL.n210 VTAIL.n209 5.81868
R919 VTAIL.n271 VTAIL.n240 5.81868
R920 VTAIL.n276 VTAIL.n236 5.81868
R921 VTAIL.n318 VTAIL.n317 5.81868
R922 VTAIL.n746 VTAIL.n745 5.81868
R923 VTAIL.n705 VTAIL.n665 5.81868
R924 VTAIL.n700 VTAIL.n669 5.81868
R925 VTAIL.n638 VTAIL.n637 5.81868
R926 VTAIL.n597 VTAIL.n557 5.81868
R927 VTAIL.n592 VTAIL.n561 5.81868
R928 VTAIL.n532 VTAIL.n531 5.81868
R929 VTAIL.n491 VTAIL.n451 5.81868
R930 VTAIL.n486 VTAIL.n455 5.81868
R931 VTAIL.n424 VTAIL.n423 5.81868
R932 VTAIL.n383 VTAIL.n343 5.81868
R933 VTAIL.n378 VTAIL.n347 5.81868
R934 VTAIL.n802 VTAIL.n801 5.04292
R935 VTAIL.n814 VTAIL.n813 5.04292
R936 VTAIL.n848 VTAIL.n752 5.04292
R937 VTAIL.n54 VTAIL.n53 5.04292
R938 VTAIL.n66 VTAIL.n65 5.04292
R939 VTAIL.n100 VTAIL.n4 5.04292
R940 VTAIL.n160 VTAIL.n159 5.04292
R941 VTAIL.n172 VTAIL.n171 5.04292
R942 VTAIL.n206 VTAIL.n110 5.04292
R943 VTAIL.n268 VTAIL.n267 5.04292
R944 VTAIL.n280 VTAIL.n279 5.04292
R945 VTAIL.n314 VTAIL.n218 5.04292
R946 VTAIL.n742 VTAIL.n646 5.04292
R947 VTAIL.n709 VTAIL.n708 5.04292
R948 VTAIL.n697 VTAIL.n696 5.04292
R949 VTAIL.n634 VTAIL.n538 5.04292
R950 VTAIL.n601 VTAIL.n600 5.04292
R951 VTAIL.n589 VTAIL.n588 5.04292
R952 VTAIL.n528 VTAIL.n432 5.04292
R953 VTAIL.n495 VTAIL.n494 5.04292
R954 VTAIL.n483 VTAIL.n482 5.04292
R955 VTAIL.n420 VTAIL.n324 5.04292
R956 VTAIL.n387 VTAIL.n386 5.04292
R957 VTAIL.n375 VTAIL.n374 5.04292
R958 VTAIL.n682 VTAIL.n678 4.38563
R959 VTAIL.n574 VTAIL.n570 4.38563
R960 VTAIL.n468 VTAIL.n464 4.38563
R961 VTAIL.n360 VTAIL.n356 4.38563
R962 VTAIL.n787 VTAIL.n783 4.38563
R963 VTAIL.n39 VTAIL.n35 4.38563
R964 VTAIL.n145 VTAIL.n141 4.38563
R965 VTAIL.n253 VTAIL.n249 4.38563
R966 VTAIL.n798 VTAIL.n776 4.26717
R967 VTAIL.n817 VTAIL.n768 4.26717
R968 VTAIL.n847 VTAIL.n754 4.26717
R969 VTAIL.n50 VTAIL.n28 4.26717
R970 VTAIL.n69 VTAIL.n20 4.26717
R971 VTAIL.n99 VTAIL.n6 4.26717
R972 VTAIL.n156 VTAIL.n134 4.26717
R973 VTAIL.n175 VTAIL.n126 4.26717
R974 VTAIL.n205 VTAIL.n112 4.26717
R975 VTAIL.n264 VTAIL.n242 4.26717
R976 VTAIL.n283 VTAIL.n234 4.26717
R977 VTAIL.n313 VTAIL.n220 4.26717
R978 VTAIL.n741 VTAIL.n648 4.26717
R979 VTAIL.n712 VTAIL.n663 4.26717
R980 VTAIL.n693 VTAIL.n671 4.26717
R981 VTAIL.n633 VTAIL.n540 4.26717
R982 VTAIL.n604 VTAIL.n555 4.26717
R983 VTAIL.n585 VTAIL.n563 4.26717
R984 VTAIL.n527 VTAIL.n434 4.26717
R985 VTAIL.n498 VTAIL.n449 4.26717
R986 VTAIL.n479 VTAIL.n457 4.26717
R987 VTAIL.n419 VTAIL.n326 4.26717
R988 VTAIL.n390 VTAIL.n341 4.26717
R989 VTAIL.n371 VTAIL.n349 4.26717
R990 VTAIL.n797 VTAIL.n778 3.49141
R991 VTAIL.n818 VTAIL.n766 3.49141
R992 VTAIL.n844 VTAIL.n843 3.49141
R993 VTAIL.n49 VTAIL.n30 3.49141
R994 VTAIL.n70 VTAIL.n18 3.49141
R995 VTAIL.n96 VTAIL.n95 3.49141
R996 VTAIL.n155 VTAIL.n136 3.49141
R997 VTAIL.n176 VTAIL.n124 3.49141
R998 VTAIL.n202 VTAIL.n201 3.49141
R999 VTAIL.n263 VTAIL.n244 3.49141
R1000 VTAIL.n284 VTAIL.n232 3.49141
R1001 VTAIL.n310 VTAIL.n309 3.49141
R1002 VTAIL.n738 VTAIL.n737 3.49141
R1003 VTAIL.n713 VTAIL.n661 3.49141
R1004 VTAIL.n692 VTAIL.n673 3.49141
R1005 VTAIL.n630 VTAIL.n629 3.49141
R1006 VTAIL.n605 VTAIL.n553 3.49141
R1007 VTAIL.n584 VTAIL.n565 3.49141
R1008 VTAIL.n524 VTAIL.n523 3.49141
R1009 VTAIL.n499 VTAIL.n447 3.49141
R1010 VTAIL.n478 VTAIL.n459 3.49141
R1011 VTAIL.n416 VTAIL.n415 3.49141
R1012 VTAIL.n391 VTAIL.n339 3.49141
R1013 VTAIL.n370 VTAIL.n351 3.49141
R1014 VTAIL.n794 VTAIL.n793 2.71565
R1015 VTAIL.n822 VTAIL.n821 2.71565
R1016 VTAIL.n840 VTAIL.n756 2.71565
R1017 VTAIL.n46 VTAIL.n45 2.71565
R1018 VTAIL.n74 VTAIL.n73 2.71565
R1019 VTAIL.n92 VTAIL.n8 2.71565
R1020 VTAIL.n152 VTAIL.n151 2.71565
R1021 VTAIL.n180 VTAIL.n179 2.71565
R1022 VTAIL.n198 VTAIL.n114 2.71565
R1023 VTAIL.n260 VTAIL.n259 2.71565
R1024 VTAIL.n288 VTAIL.n287 2.71565
R1025 VTAIL.n306 VTAIL.n222 2.71565
R1026 VTAIL.n734 VTAIL.n650 2.71565
R1027 VTAIL.n717 VTAIL.n716 2.71565
R1028 VTAIL.n689 VTAIL.n688 2.71565
R1029 VTAIL.n626 VTAIL.n542 2.71565
R1030 VTAIL.n609 VTAIL.n608 2.71565
R1031 VTAIL.n581 VTAIL.n580 2.71565
R1032 VTAIL.n520 VTAIL.n436 2.71565
R1033 VTAIL.n503 VTAIL.n502 2.71565
R1034 VTAIL.n475 VTAIL.n474 2.71565
R1035 VTAIL.n412 VTAIL.n328 2.71565
R1036 VTAIL.n395 VTAIL.n394 2.71565
R1037 VTAIL.n367 VTAIL.n366 2.71565
R1038 VTAIL.n790 VTAIL.n780 1.93989
R1039 VTAIL.n826 VTAIL.n764 1.93989
R1040 VTAIL.n839 VTAIL.n758 1.93989
R1041 VTAIL.n42 VTAIL.n32 1.93989
R1042 VTAIL.n78 VTAIL.n16 1.93989
R1043 VTAIL.n91 VTAIL.n10 1.93989
R1044 VTAIL.n148 VTAIL.n138 1.93989
R1045 VTAIL.n184 VTAIL.n122 1.93989
R1046 VTAIL.n197 VTAIL.n116 1.93989
R1047 VTAIL.n256 VTAIL.n246 1.93989
R1048 VTAIL.n292 VTAIL.n230 1.93989
R1049 VTAIL.n305 VTAIL.n224 1.93989
R1050 VTAIL.n733 VTAIL.n652 1.93989
R1051 VTAIL.n720 VTAIL.n658 1.93989
R1052 VTAIL.n685 VTAIL.n675 1.93989
R1053 VTAIL.n625 VTAIL.n544 1.93989
R1054 VTAIL.n612 VTAIL.n550 1.93989
R1055 VTAIL.n577 VTAIL.n567 1.93989
R1056 VTAIL.n519 VTAIL.n438 1.93989
R1057 VTAIL.n506 VTAIL.n444 1.93989
R1058 VTAIL.n471 VTAIL.n461 1.93989
R1059 VTAIL.n411 VTAIL.n330 1.93989
R1060 VTAIL.n398 VTAIL.n336 1.93989
R1061 VTAIL.n363 VTAIL.n353 1.93989
R1062 VTAIL.n789 VTAIL.n782 1.16414
R1063 VTAIL.n827 VTAIL.n762 1.16414
R1064 VTAIL.n836 VTAIL.n835 1.16414
R1065 VTAIL.n41 VTAIL.n34 1.16414
R1066 VTAIL.n79 VTAIL.n14 1.16414
R1067 VTAIL.n88 VTAIL.n87 1.16414
R1068 VTAIL.n147 VTAIL.n140 1.16414
R1069 VTAIL.n185 VTAIL.n120 1.16414
R1070 VTAIL.n194 VTAIL.n193 1.16414
R1071 VTAIL.n255 VTAIL.n248 1.16414
R1072 VTAIL.n293 VTAIL.n228 1.16414
R1073 VTAIL.n302 VTAIL.n301 1.16414
R1074 VTAIL.n730 VTAIL.n729 1.16414
R1075 VTAIL.n721 VTAIL.n656 1.16414
R1076 VTAIL.n684 VTAIL.n677 1.16414
R1077 VTAIL.n622 VTAIL.n621 1.16414
R1078 VTAIL.n613 VTAIL.n548 1.16414
R1079 VTAIL.n576 VTAIL.n569 1.16414
R1080 VTAIL.n516 VTAIL.n515 1.16414
R1081 VTAIL.n507 VTAIL.n442 1.16414
R1082 VTAIL.n470 VTAIL.n463 1.16414
R1083 VTAIL.n408 VTAIL.n407 1.16414
R1084 VTAIL.n399 VTAIL.n334 1.16414
R1085 VTAIL.n362 VTAIL.n355 1.16414
R1086 VTAIL.n0 VTAIL.t11 1.04701
R1087 VTAIL.n0 VTAIL.t15 1.04701
R1088 VTAIL.n214 VTAIL.t5 1.04701
R1089 VTAIL.n214 VTAIL.t4 1.04701
R1090 VTAIL.n642 VTAIL.t1 1.04701
R1091 VTAIL.n642 VTAIL.t6 1.04701
R1092 VTAIL.n428 VTAIL.t12 1.04701
R1093 VTAIL.n428 VTAIL.t13 1.04701
R1094 VTAIL.n429 VTAIL.n427 0.578086
R1095 VTAIL.n535 VTAIL.n429 0.578086
R1096 VTAIL.n643 VTAIL.n641 0.578086
R1097 VTAIL.n749 VTAIL.n643 0.578086
R1098 VTAIL.n321 VTAIL.n215 0.578086
R1099 VTAIL.n215 VTAIL.n213 0.578086
R1100 VTAIL.n107 VTAIL.n1 0.578086
R1101 VTAIL VTAIL.n855 0.519897
R1102 VTAIL.n641 VTAIL.n535 0.470328
R1103 VTAIL.n213 VTAIL.n107 0.470328
R1104 VTAIL.n786 VTAIL.n785 0.388379
R1105 VTAIL.n831 VTAIL.n830 0.388379
R1106 VTAIL.n832 VTAIL.n760 0.388379
R1107 VTAIL.n38 VTAIL.n37 0.388379
R1108 VTAIL.n83 VTAIL.n82 0.388379
R1109 VTAIL.n84 VTAIL.n12 0.388379
R1110 VTAIL.n144 VTAIL.n143 0.388379
R1111 VTAIL.n189 VTAIL.n188 0.388379
R1112 VTAIL.n190 VTAIL.n118 0.388379
R1113 VTAIL.n252 VTAIL.n251 0.388379
R1114 VTAIL.n297 VTAIL.n296 0.388379
R1115 VTAIL.n298 VTAIL.n226 0.388379
R1116 VTAIL.n726 VTAIL.n654 0.388379
R1117 VTAIL.n725 VTAIL.n724 0.388379
R1118 VTAIL.n681 VTAIL.n680 0.388379
R1119 VTAIL.n618 VTAIL.n546 0.388379
R1120 VTAIL.n617 VTAIL.n616 0.388379
R1121 VTAIL.n573 VTAIL.n572 0.388379
R1122 VTAIL.n512 VTAIL.n440 0.388379
R1123 VTAIL.n511 VTAIL.n510 0.388379
R1124 VTAIL.n467 VTAIL.n466 0.388379
R1125 VTAIL.n404 VTAIL.n332 0.388379
R1126 VTAIL.n403 VTAIL.n402 0.388379
R1127 VTAIL.n359 VTAIL.n358 0.388379
R1128 VTAIL.n788 VTAIL.n787 0.155672
R1129 VTAIL.n788 VTAIL.n779 0.155672
R1130 VTAIL.n795 VTAIL.n779 0.155672
R1131 VTAIL.n796 VTAIL.n795 0.155672
R1132 VTAIL.n796 VTAIL.n775 0.155672
R1133 VTAIL.n803 VTAIL.n775 0.155672
R1134 VTAIL.n804 VTAIL.n803 0.155672
R1135 VTAIL.n804 VTAIL.n771 0.155672
R1136 VTAIL.n811 VTAIL.n771 0.155672
R1137 VTAIL.n812 VTAIL.n811 0.155672
R1138 VTAIL.n812 VTAIL.n767 0.155672
R1139 VTAIL.n819 VTAIL.n767 0.155672
R1140 VTAIL.n820 VTAIL.n819 0.155672
R1141 VTAIL.n820 VTAIL.n763 0.155672
R1142 VTAIL.n828 VTAIL.n763 0.155672
R1143 VTAIL.n829 VTAIL.n828 0.155672
R1144 VTAIL.n829 VTAIL.n759 0.155672
R1145 VTAIL.n837 VTAIL.n759 0.155672
R1146 VTAIL.n838 VTAIL.n837 0.155672
R1147 VTAIL.n838 VTAIL.n755 0.155672
R1148 VTAIL.n845 VTAIL.n755 0.155672
R1149 VTAIL.n846 VTAIL.n845 0.155672
R1150 VTAIL.n846 VTAIL.n751 0.155672
R1151 VTAIL.n853 VTAIL.n751 0.155672
R1152 VTAIL.n40 VTAIL.n39 0.155672
R1153 VTAIL.n40 VTAIL.n31 0.155672
R1154 VTAIL.n47 VTAIL.n31 0.155672
R1155 VTAIL.n48 VTAIL.n47 0.155672
R1156 VTAIL.n48 VTAIL.n27 0.155672
R1157 VTAIL.n55 VTAIL.n27 0.155672
R1158 VTAIL.n56 VTAIL.n55 0.155672
R1159 VTAIL.n56 VTAIL.n23 0.155672
R1160 VTAIL.n63 VTAIL.n23 0.155672
R1161 VTAIL.n64 VTAIL.n63 0.155672
R1162 VTAIL.n64 VTAIL.n19 0.155672
R1163 VTAIL.n71 VTAIL.n19 0.155672
R1164 VTAIL.n72 VTAIL.n71 0.155672
R1165 VTAIL.n72 VTAIL.n15 0.155672
R1166 VTAIL.n80 VTAIL.n15 0.155672
R1167 VTAIL.n81 VTAIL.n80 0.155672
R1168 VTAIL.n81 VTAIL.n11 0.155672
R1169 VTAIL.n89 VTAIL.n11 0.155672
R1170 VTAIL.n90 VTAIL.n89 0.155672
R1171 VTAIL.n90 VTAIL.n7 0.155672
R1172 VTAIL.n97 VTAIL.n7 0.155672
R1173 VTAIL.n98 VTAIL.n97 0.155672
R1174 VTAIL.n98 VTAIL.n3 0.155672
R1175 VTAIL.n105 VTAIL.n3 0.155672
R1176 VTAIL.n146 VTAIL.n145 0.155672
R1177 VTAIL.n146 VTAIL.n137 0.155672
R1178 VTAIL.n153 VTAIL.n137 0.155672
R1179 VTAIL.n154 VTAIL.n153 0.155672
R1180 VTAIL.n154 VTAIL.n133 0.155672
R1181 VTAIL.n161 VTAIL.n133 0.155672
R1182 VTAIL.n162 VTAIL.n161 0.155672
R1183 VTAIL.n162 VTAIL.n129 0.155672
R1184 VTAIL.n169 VTAIL.n129 0.155672
R1185 VTAIL.n170 VTAIL.n169 0.155672
R1186 VTAIL.n170 VTAIL.n125 0.155672
R1187 VTAIL.n177 VTAIL.n125 0.155672
R1188 VTAIL.n178 VTAIL.n177 0.155672
R1189 VTAIL.n178 VTAIL.n121 0.155672
R1190 VTAIL.n186 VTAIL.n121 0.155672
R1191 VTAIL.n187 VTAIL.n186 0.155672
R1192 VTAIL.n187 VTAIL.n117 0.155672
R1193 VTAIL.n195 VTAIL.n117 0.155672
R1194 VTAIL.n196 VTAIL.n195 0.155672
R1195 VTAIL.n196 VTAIL.n113 0.155672
R1196 VTAIL.n203 VTAIL.n113 0.155672
R1197 VTAIL.n204 VTAIL.n203 0.155672
R1198 VTAIL.n204 VTAIL.n109 0.155672
R1199 VTAIL.n211 VTAIL.n109 0.155672
R1200 VTAIL.n254 VTAIL.n253 0.155672
R1201 VTAIL.n254 VTAIL.n245 0.155672
R1202 VTAIL.n261 VTAIL.n245 0.155672
R1203 VTAIL.n262 VTAIL.n261 0.155672
R1204 VTAIL.n262 VTAIL.n241 0.155672
R1205 VTAIL.n269 VTAIL.n241 0.155672
R1206 VTAIL.n270 VTAIL.n269 0.155672
R1207 VTAIL.n270 VTAIL.n237 0.155672
R1208 VTAIL.n277 VTAIL.n237 0.155672
R1209 VTAIL.n278 VTAIL.n277 0.155672
R1210 VTAIL.n278 VTAIL.n233 0.155672
R1211 VTAIL.n285 VTAIL.n233 0.155672
R1212 VTAIL.n286 VTAIL.n285 0.155672
R1213 VTAIL.n286 VTAIL.n229 0.155672
R1214 VTAIL.n294 VTAIL.n229 0.155672
R1215 VTAIL.n295 VTAIL.n294 0.155672
R1216 VTAIL.n295 VTAIL.n225 0.155672
R1217 VTAIL.n303 VTAIL.n225 0.155672
R1218 VTAIL.n304 VTAIL.n303 0.155672
R1219 VTAIL.n304 VTAIL.n221 0.155672
R1220 VTAIL.n311 VTAIL.n221 0.155672
R1221 VTAIL.n312 VTAIL.n311 0.155672
R1222 VTAIL.n312 VTAIL.n217 0.155672
R1223 VTAIL.n319 VTAIL.n217 0.155672
R1224 VTAIL.n747 VTAIL.n645 0.155672
R1225 VTAIL.n740 VTAIL.n645 0.155672
R1226 VTAIL.n740 VTAIL.n739 0.155672
R1227 VTAIL.n739 VTAIL.n649 0.155672
R1228 VTAIL.n732 VTAIL.n649 0.155672
R1229 VTAIL.n732 VTAIL.n731 0.155672
R1230 VTAIL.n731 VTAIL.n653 0.155672
R1231 VTAIL.n723 VTAIL.n653 0.155672
R1232 VTAIL.n723 VTAIL.n722 0.155672
R1233 VTAIL.n722 VTAIL.n657 0.155672
R1234 VTAIL.n715 VTAIL.n657 0.155672
R1235 VTAIL.n715 VTAIL.n714 0.155672
R1236 VTAIL.n714 VTAIL.n662 0.155672
R1237 VTAIL.n707 VTAIL.n662 0.155672
R1238 VTAIL.n707 VTAIL.n706 0.155672
R1239 VTAIL.n706 VTAIL.n666 0.155672
R1240 VTAIL.n699 VTAIL.n666 0.155672
R1241 VTAIL.n699 VTAIL.n698 0.155672
R1242 VTAIL.n698 VTAIL.n670 0.155672
R1243 VTAIL.n691 VTAIL.n670 0.155672
R1244 VTAIL.n691 VTAIL.n690 0.155672
R1245 VTAIL.n690 VTAIL.n674 0.155672
R1246 VTAIL.n683 VTAIL.n674 0.155672
R1247 VTAIL.n683 VTAIL.n682 0.155672
R1248 VTAIL.n639 VTAIL.n537 0.155672
R1249 VTAIL.n632 VTAIL.n537 0.155672
R1250 VTAIL.n632 VTAIL.n631 0.155672
R1251 VTAIL.n631 VTAIL.n541 0.155672
R1252 VTAIL.n624 VTAIL.n541 0.155672
R1253 VTAIL.n624 VTAIL.n623 0.155672
R1254 VTAIL.n623 VTAIL.n545 0.155672
R1255 VTAIL.n615 VTAIL.n545 0.155672
R1256 VTAIL.n615 VTAIL.n614 0.155672
R1257 VTAIL.n614 VTAIL.n549 0.155672
R1258 VTAIL.n607 VTAIL.n549 0.155672
R1259 VTAIL.n607 VTAIL.n606 0.155672
R1260 VTAIL.n606 VTAIL.n554 0.155672
R1261 VTAIL.n599 VTAIL.n554 0.155672
R1262 VTAIL.n599 VTAIL.n598 0.155672
R1263 VTAIL.n598 VTAIL.n558 0.155672
R1264 VTAIL.n591 VTAIL.n558 0.155672
R1265 VTAIL.n591 VTAIL.n590 0.155672
R1266 VTAIL.n590 VTAIL.n562 0.155672
R1267 VTAIL.n583 VTAIL.n562 0.155672
R1268 VTAIL.n583 VTAIL.n582 0.155672
R1269 VTAIL.n582 VTAIL.n566 0.155672
R1270 VTAIL.n575 VTAIL.n566 0.155672
R1271 VTAIL.n575 VTAIL.n574 0.155672
R1272 VTAIL.n533 VTAIL.n431 0.155672
R1273 VTAIL.n526 VTAIL.n431 0.155672
R1274 VTAIL.n526 VTAIL.n525 0.155672
R1275 VTAIL.n525 VTAIL.n435 0.155672
R1276 VTAIL.n518 VTAIL.n435 0.155672
R1277 VTAIL.n518 VTAIL.n517 0.155672
R1278 VTAIL.n517 VTAIL.n439 0.155672
R1279 VTAIL.n509 VTAIL.n439 0.155672
R1280 VTAIL.n509 VTAIL.n508 0.155672
R1281 VTAIL.n508 VTAIL.n443 0.155672
R1282 VTAIL.n501 VTAIL.n443 0.155672
R1283 VTAIL.n501 VTAIL.n500 0.155672
R1284 VTAIL.n500 VTAIL.n448 0.155672
R1285 VTAIL.n493 VTAIL.n448 0.155672
R1286 VTAIL.n493 VTAIL.n492 0.155672
R1287 VTAIL.n492 VTAIL.n452 0.155672
R1288 VTAIL.n485 VTAIL.n452 0.155672
R1289 VTAIL.n485 VTAIL.n484 0.155672
R1290 VTAIL.n484 VTAIL.n456 0.155672
R1291 VTAIL.n477 VTAIL.n456 0.155672
R1292 VTAIL.n477 VTAIL.n476 0.155672
R1293 VTAIL.n476 VTAIL.n460 0.155672
R1294 VTAIL.n469 VTAIL.n460 0.155672
R1295 VTAIL.n469 VTAIL.n468 0.155672
R1296 VTAIL.n425 VTAIL.n323 0.155672
R1297 VTAIL.n418 VTAIL.n323 0.155672
R1298 VTAIL.n418 VTAIL.n417 0.155672
R1299 VTAIL.n417 VTAIL.n327 0.155672
R1300 VTAIL.n410 VTAIL.n327 0.155672
R1301 VTAIL.n410 VTAIL.n409 0.155672
R1302 VTAIL.n409 VTAIL.n331 0.155672
R1303 VTAIL.n401 VTAIL.n331 0.155672
R1304 VTAIL.n401 VTAIL.n400 0.155672
R1305 VTAIL.n400 VTAIL.n335 0.155672
R1306 VTAIL.n393 VTAIL.n335 0.155672
R1307 VTAIL.n393 VTAIL.n392 0.155672
R1308 VTAIL.n392 VTAIL.n340 0.155672
R1309 VTAIL.n385 VTAIL.n340 0.155672
R1310 VTAIL.n385 VTAIL.n384 0.155672
R1311 VTAIL.n384 VTAIL.n344 0.155672
R1312 VTAIL.n377 VTAIL.n344 0.155672
R1313 VTAIL.n377 VTAIL.n376 0.155672
R1314 VTAIL.n376 VTAIL.n348 0.155672
R1315 VTAIL.n369 VTAIL.n348 0.155672
R1316 VTAIL.n369 VTAIL.n368 0.155672
R1317 VTAIL.n368 VTAIL.n352 0.155672
R1318 VTAIL.n361 VTAIL.n352 0.155672
R1319 VTAIL.n361 VTAIL.n360 0.155672
R1320 VTAIL VTAIL.n1 0.0586897
R1321 VDD2.n2 VDD2.n1 60.0797
R1322 VDD2.n2 VDD2.n0 60.0797
R1323 VDD2 VDD2.n5 60.0767
R1324 VDD2.n4 VDD2.n3 59.8462
R1325 VDD2.n4 VDD2.n2 42.6248
R1326 VDD2.n5 VDD2.t6 1.04701
R1327 VDD2.n5 VDD2.t2 1.04701
R1328 VDD2.n3 VDD2.t0 1.04701
R1329 VDD2.n3 VDD2.t7 1.04701
R1330 VDD2.n1 VDD2.t5 1.04701
R1331 VDD2.n1 VDD2.t3 1.04701
R1332 VDD2.n0 VDD2.t1 1.04701
R1333 VDD2.n0 VDD2.t4 1.04701
R1334 VDD2 VDD2.n4 0.347483
R1335 B.n183 B.t16 1553.17
R1336 B.n176 B.t8 1553.17
R1337 B.n68 B.t12 1553.17
R1338 B.n76 B.t19 1553.17
R1339 B.n563 B.n562 585
R1340 B.n564 B.n109 585
R1341 B.n566 B.n565 585
R1342 B.n568 B.n108 585
R1343 B.n571 B.n570 585
R1344 B.n572 B.n107 585
R1345 B.n574 B.n573 585
R1346 B.n576 B.n106 585
R1347 B.n579 B.n578 585
R1348 B.n580 B.n105 585
R1349 B.n582 B.n581 585
R1350 B.n584 B.n104 585
R1351 B.n587 B.n586 585
R1352 B.n588 B.n103 585
R1353 B.n590 B.n589 585
R1354 B.n592 B.n102 585
R1355 B.n595 B.n594 585
R1356 B.n596 B.n101 585
R1357 B.n598 B.n597 585
R1358 B.n600 B.n100 585
R1359 B.n603 B.n602 585
R1360 B.n604 B.n99 585
R1361 B.n606 B.n605 585
R1362 B.n608 B.n98 585
R1363 B.n611 B.n610 585
R1364 B.n612 B.n97 585
R1365 B.n614 B.n613 585
R1366 B.n616 B.n96 585
R1367 B.n619 B.n618 585
R1368 B.n620 B.n95 585
R1369 B.n622 B.n621 585
R1370 B.n624 B.n94 585
R1371 B.n627 B.n626 585
R1372 B.n628 B.n93 585
R1373 B.n630 B.n629 585
R1374 B.n632 B.n92 585
R1375 B.n635 B.n634 585
R1376 B.n636 B.n91 585
R1377 B.n638 B.n637 585
R1378 B.n640 B.n90 585
R1379 B.n643 B.n642 585
R1380 B.n644 B.n89 585
R1381 B.n646 B.n645 585
R1382 B.n648 B.n88 585
R1383 B.n651 B.n650 585
R1384 B.n652 B.n87 585
R1385 B.n654 B.n653 585
R1386 B.n656 B.n86 585
R1387 B.n659 B.n658 585
R1388 B.n660 B.n85 585
R1389 B.n662 B.n661 585
R1390 B.n664 B.n84 585
R1391 B.n667 B.n666 585
R1392 B.n668 B.n83 585
R1393 B.n670 B.n669 585
R1394 B.n672 B.n82 585
R1395 B.n675 B.n674 585
R1396 B.n676 B.n81 585
R1397 B.n678 B.n677 585
R1398 B.n680 B.n80 585
R1399 B.n682 B.n681 585
R1400 B.n684 B.n683 585
R1401 B.n687 B.n686 585
R1402 B.n688 B.n75 585
R1403 B.n690 B.n689 585
R1404 B.n692 B.n74 585
R1405 B.n695 B.n694 585
R1406 B.n696 B.n73 585
R1407 B.n698 B.n697 585
R1408 B.n700 B.n72 585
R1409 B.n702 B.n701 585
R1410 B.n704 B.n703 585
R1411 B.n707 B.n706 585
R1412 B.n708 B.n67 585
R1413 B.n710 B.n709 585
R1414 B.n712 B.n66 585
R1415 B.n715 B.n714 585
R1416 B.n716 B.n65 585
R1417 B.n718 B.n717 585
R1418 B.n720 B.n64 585
R1419 B.n723 B.n722 585
R1420 B.n724 B.n63 585
R1421 B.n726 B.n725 585
R1422 B.n728 B.n62 585
R1423 B.n731 B.n730 585
R1424 B.n732 B.n61 585
R1425 B.n734 B.n733 585
R1426 B.n736 B.n60 585
R1427 B.n739 B.n738 585
R1428 B.n740 B.n59 585
R1429 B.n742 B.n741 585
R1430 B.n744 B.n58 585
R1431 B.n747 B.n746 585
R1432 B.n748 B.n57 585
R1433 B.n750 B.n749 585
R1434 B.n752 B.n56 585
R1435 B.n755 B.n754 585
R1436 B.n756 B.n55 585
R1437 B.n758 B.n757 585
R1438 B.n760 B.n54 585
R1439 B.n763 B.n762 585
R1440 B.n764 B.n53 585
R1441 B.n766 B.n765 585
R1442 B.n768 B.n52 585
R1443 B.n771 B.n770 585
R1444 B.n772 B.n51 585
R1445 B.n774 B.n773 585
R1446 B.n776 B.n50 585
R1447 B.n779 B.n778 585
R1448 B.n780 B.n49 585
R1449 B.n782 B.n781 585
R1450 B.n784 B.n48 585
R1451 B.n787 B.n786 585
R1452 B.n788 B.n47 585
R1453 B.n790 B.n789 585
R1454 B.n792 B.n46 585
R1455 B.n795 B.n794 585
R1456 B.n796 B.n45 585
R1457 B.n798 B.n797 585
R1458 B.n800 B.n44 585
R1459 B.n803 B.n802 585
R1460 B.n804 B.n43 585
R1461 B.n806 B.n805 585
R1462 B.n808 B.n42 585
R1463 B.n811 B.n810 585
R1464 B.n812 B.n41 585
R1465 B.n814 B.n813 585
R1466 B.n816 B.n40 585
R1467 B.n819 B.n818 585
R1468 B.n820 B.n39 585
R1469 B.n822 B.n821 585
R1470 B.n824 B.n38 585
R1471 B.n827 B.n826 585
R1472 B.n828 B.n37 585
R1473 B.n560 B.n35 585
R1474 B.n831 B.n35 585
R1475 B.n559 B.n34 585
R1476 B.n832 B.n34 585
R1477 B.n558 B.n33 585
R1478 B.n833 B.n33 585
R1479 B.n557 B.n556 585
R1480 B.n556 B.n29 585
R1481 B.n555 B.n28 585
R1482 B.n839 B.n28 585
R1483 B.n554 B.n27 585
R1484 B.n840 B.n27 585
R1485 B.n553 B.n26 585
R1486 B.n841 B.n26 585
R1487 B.n552 B.n551 585
R1488 B.n551 B.n22 585
R1489 B.n550 B.n21 585
R1490 B.n847 B.n21 585
R1491 B.n549 B.n20 585
R1492 B.n848 B.n20 585
R1493 B.n548 B.n19 585
R1494 B.n849 B.n19 585
R1495 B.n547 B.n546 585
R1496 B.n546 B.n18 585
R1497 B.n545 B.n14 585
R1498 B.n855 B.n14 585
R1499 B.n544 B.n13 585
R1500 B.n856 B.n13 585
R1501 B.n543 B.n12 585
R1502 B.n857 B.n12 585
R1503 B.n542 B.n541 585
R1504 B.n541 B.n11 585
R1505 B.n540 B.n7 585
R1506 B.n863 B.n7 585
R1507 B.n539 B.n6 585
R1508 B.n864 B.n6 585
R1509 B.n538 B.n5 585
R1510 B.n865 B.n5 585
R1511 B.n537 B.n536 585
R1512 B.n536 B.n4 585
R1513 B.n535 B.n110 585
R1514 B.n535 B.n534 585
R1515 B.n524 B.n111 585
R1516 B.n527 B.n111 585
R1517 B.n526 B.n525 585
R1518 B.n528 B.n526 585
R1519 B.n523 B.n115 585
R1520 B.n118 B.n115 585
R1521 B.n522 B.n521 585
R1522 B.n521 B.n520 585
R1523 B.n117 B.n116 585
R1524 B.n513 B.n117 585
R1525 B.n512 B.n511 585
R1526 B.n514 B.n512 585
R1527 B.n510 B.n122 585
R1528 B.n126 B.n122 585
R1529 B.n509 B.n508 585
R1530 B.n508 B.n507 585
R1531 B.n124 B.n123 585
R1532 B.n125 B.n124 585
R1533 B.n500 B.n499 585
R1534 B.n501 B.n500 585
R1535 B.n498 B.n131 585
R1536 B.n131 B.n130 585
R1537 B.n497 B.n496 585
R1538 B.n496 B.n495 585
R1539 B.n133 B.n132 585
R1540 B.n134 B.n133 585
R1541 B.n488 B.n487 585
R1542 B.n489 B.n488 585
R1543 B.n486 B.n139 585
R1544 B.n139 B.n138 585
R1545 B.n485 B.n484 585
R1546 B.n484 B.n483 585
R1547 B.n480 B.n143 585
R1548 B.n479 B.n478 585
R1549 B.n476 B.n144 585
R1550 B.n476 B.n142 585
R1551 B.n475 B.n474 585
R1552 B.n473 B.n472 585
R1553 B.n471 B.n146 585
R1554 B.n469 B.n468 585
R1555 B.n467 B.n147 585
R1556 B.n466 B.n465 585
R1557 B.n463 B.n148 585
R1558 B.n461 B.n460 585
R1559 B.n459 B.n149 585
R1560 B.n458 B.n457 585
R1561 B.n455 B.n150 585
R1562 B.n453 B.n452 585
R1563 B.n451 B.n151 585
R1564 B.n450 B.n449 585
R1565 B.n447 B.n152 585
R1566 B.n445 B.n444 585
R1567 B.n443 B.n153 585
R1568 B.n442 B.n441 585
R1569 B.n439 B.n154 585
R1570 B.n437 B.n436 585
R1571 B.n435 B.n155 585
R1572 B.n434 B.n433 585
R1573 B.n431 B.n156 585
R1574 B.n429 B.n428 585
R1575 B.n427 B.n157 585
R1576 B.n426 B.n425 585
R1577 B.n423 B.n158 585
R1578 B.n421 B.n420 585
R1579 B.n419 B.n159 585
R1580 B.n418 B.n417 585
R1581 B.n415 B.n160 585
R1582 B.n413 B.n412 585
R1583 B.n411 B.n161 585
R1584 B.n410 B.n409 585
R1585 B.n407 B.n162 585
R1586 B.n405 B.n404 585
R1587 B.n403 B.n163 585
R1588 B.n402 B.n401 585
R1589 B.n399 B.n164 585
R1590 B.n397 B.n396 585
R1591 B.n395 B.n165 585
R1592 B.n394 B.n393 585
R1593 B.n391 B.n166 585
R1594 B.n389 B.n388 585
R1595 B.n387 B.n167 585
R1596 B.n386 B.n385 585
R1597 B.n383 B.n168 585
R1598 B.n381 B.n380 585
R1599 B.n379 B.n169 585
R1600 B.n378 B.n377 585
R1601 B.n375 B.n170 585
R1602 B.n373 B.n372 585
R1603 B.n371 B.n171 585
R1604 B.n370 B.n369 585
R1605 B.n367 B.n172 585
R1606 B.n365 B.n364 585
R1607 B.n363 B.n173 585
R1608 B.n362 B.n361 585
R1609 B.n359 B.n174 585
R1610 B.n357 B.n356 585
R1611 B.n355 B.n175 585
R1612 B.n354 B.n353 585
R1613 B.n351 B.n179 585
R1614 B.n349 B.n348 585
R1615 B.n347 B.n180 585
R1616 B.n346 B.n345 585
R1617 B.n343 B.n181 585
R1618 B.n341 B.n340 585
R1619 B.n339 B.n182 585
R1620 B.n337 B.n336 585
R1621 B.n334 B.n185 585
R1622 B.n332 B.n331 585
R1623 B.n330 B.n186 585
R1624 B.n329 B.n328 585
R1625 B.n326 B.n187 585
R1626 B.n324 B.n323 585
R1627 B.n322 B.n188 585
R1628 B.n321 B.n320 585
R1629 B.n318 B.n189 585
R1630 B.n316 B.n315 585
R1631 B.n314 B.n190 585
R1632 B.n313 B.n312 585
R1633 B.n310 B.n191 585
R1634 B.n308 B.n307 585
R1635 B.n306 B.n192 585
R1636 B.n305 B.n304 585
R1637 B.n302 B.n193 585
R1638 B.n300 B.n299 585
R1639 B.n298 B.n194 585
R1640 B.n297 B.n296 585
R1641 B.n294 B.n195 585
R1642 B.n292 B.n291 585
R1643 B.n290 B.n196 585
R1644 B.n289 B.n288 585
R1645 B.n286 B.n197 585
R1646 B.n284 B.n283 585
R1647 B.n282 B.n198 585
R1648 B.n281 B.n280 585
R1649 B.n278 B.n199 585
R1650 B.n276 B.n275 585
R1651 B.n274 B.n200 585
R1652 B.n273 B.n272 585
R1653 B.n270 B.n201 585
R1654 B.n268 B.n267 585
R1655 B.n266 B.n202 585
R1656 B.n265 B.n264 585
R1657 B.n262 B.n203 585
R1658 B.n260 B.n259 585
R1659 B.n258 B.n204 585
R1660 B.n257 B.n256 585
R1661 B.n254 B.n205 585
R1662 B.n252 B.n251 585
R1663 B.n250 B.n206 585
R1664 B.n249 B.n248 585
R1665 B.n246 B.n207 585
R1666 B.n244 B.n243 585
R1667 B.n242 B.n208 585
R1668 B.n241 B.n240 585
R1669 B.n238 B.n209 585
R1670 B.n236 B.n235 585
R1671 B.n234 B.n210 585
R1672 B.n233 B.n232 585
R1673 B.n230 B.n211 585
R1674 B.n228 B.n227 585
R1675 B.n226 B.n212 585
R1676 B.n225 B.n224 585
R1677 B.n222 B.n213 585
R1678 B.n220 B.n219 585
R1679 B.n218 B.n214 585
R1680 B.n217 B.n216 585
R1681 B.n141 B.n140 585
R1682 B.n142 B.n141 585
R1683 B.n482 B.n481 585
R1684 B.n483 B.n482 585
R1685 B.n137 B.n136 585
R1686 B.n138 B.n137 585
R1687 B.n491 B.n490 585
R1688 B.n490 B.n489 585
R1689 B.n492 B.n135 585
R1690 B.n135 B.n134 585
R1691 B.n494 B.n493 585
R1692 B.n495 B.n494 585
R1693 B.n129 B.n128 585
R1694 B.n130 B.n129 585
R1695 B.n503 B.n502 585
R1696 B.n502 B.n501 585
R1697 B.n504 B.n127 585
R1698 B.n127 B.n125 585
R1699 B.n506 B.n505 585
R1700 B.n507 B.n506 585
R1701 B.n121 B.n120 585
R1702 B.n126 B.n121 585
R1703 B.n516 B.n515 585
R1704 B.n515 B.n514 585
R1705 B.n517 B.n119 585
R1706 B.n513 B.n119 585
R1707 B.n519 B.n518 585
R1708 B.n520 B.n519 585
R1709 B.n114 B.n113 585
R1710 B.n118 B.n114 585
R1711 B.n530 B.n529 585
R1712 B.n529 B.n528 585
R1713 B.n531 B.n112 585
R1714 B.n527 B.n112 585
R1715 B.n533 B.n532 585
R1716 B.n534 B.n533 585
R1717 B.n2 B.n0 585
R1718 B.n4 B.n2 585
R1719 B.n3 B.n1 585
R1720 B.n864 B.n3 585
R1721 B.n862 B.n861 585
R1722 B.n863 B.n862 585
R1723 B.n860 B.n8 585
R1724 B.n11 B.n8 585
R1725 B.n859 B.n858 585
R1726 B.n858 B.n857 585
R1727 B.n10 B.n9 585
R1728 B.n856 B.n10 585
R1729 B.n854 B.n853 585
R1730 B.n855 B.n854 585
R1731 B.n852 B.n15 585
R1732 B.n18 B.n15 585
R1733 B.n851 B.n850 585
R1734 B.n850 B.n849 585
R1735 B.n17 B.n16 585
R1736 B.n848 B.n17 585
R1737 B.n846 B.n845 585
R1738 B.n847 B.n846 585
R1739 B.n844 B.n23 585
R1740 B.n23 B.n22 585
R1741 B.n843 B.n842 585
R1742 B.n842 B.n841 585
R1743 B.n25 B.n24 585
R1744 B.n840 B.n25 585
R1745 B.n838 B.n837 585
R1746 B.n839 B.n838 585
R1747 B.n836 B.n30 585
R1748 B.n30 B.n29 585
R1749 B.n835 B.n834 585
R1750 B.n834 B.n833 585
R1751 B.n32 B.n31 585
R1752 B.n832 B.n32 585
R1753 B.n830 B.n829 585
R1754 B.n831 B.n830 585
R1755 B.n867 B.n866 585
R1756 B.n866 B.n865 585
R1757 B.n482 B.n143 454.062
R1758 B.n830 B.n37 454.062
R1759 B.n484 B.n141 454.062
R1760 B.n562 B.n35 454.062
R1761 B.n183 B.t18 414.454
R1762 B.n76 B.t20 414.454
R1763 B.n176 B.t11 414.454
R1764 B.n68 B.t14 414.454
R1765 B.n184 B.t17 401.459
R1766 B.n77 B.t21 401.459
R1767 B.n177 B.t10 401.459
R1768 B.n69 B.t15 401.459
R1769 B.n561 B.n36 256.663
R1770 B.n567 B.n36 256.663
R1771 B.n569 B.n36 256.663
R1772 B.n575 B.n36 256.663
R1773 B.n577 B.n36 256.663
R1774 B.n583 B.n36 256.663
R1775 B.n585 B.n36 256.663
R1776 B.n591 B.n36 256.663
R1777 B.n593 B.n36 256.663
R1778 B.n599 B.n36 256.663
R1779 B.n601 B.n36 256.663
R1780 B.n607 B.n36 256.663
R1781 B.n609 B.n36 256.663
R1782 B.n615 B.n36 256.663
R1783 B.n617 B.n36 256.663
R1784 B.n623 B.n36 256.663
R1785 B.n625 B.n36 256.663
R1786 B.n631 B.n36 256.663
R1787 B.n633 B.n36 256.663
R1788 B.n639 B.n36 256.663
R1789 B.n641 B.n36 256.663
R1790 B.n647 B.n36 256.663
R1791 B.n649 B.n36 256.663
R1792 B.n655 B.n36 256.663
R1793 B.n657 B.n36 256.663
R1794 B.n663 B.n36 256.663
R1795 B.n665 B.n36 256.663
R1796 B.n671 B.n36 256.663
R1797 B.n673 B.n36 256.663
R1798 B.n679 B.n36 256.663
R1799 B.n79 B.n36 256.663
R1800 B.n685 B.n36 256.663
R1801 B.n691 B.n36 256.663
R1802 B.n693 B.n36 256.663
R1803 B.n699 B.n36 256.663
R1804 B.n71 B.n36 256.663
R1805 B.n705 B.n36 256.663
R1806 B.n711 B.n36 256.663
R1807 B.n713 B.n36 256.663
R1808 B.n719 B.n36 256.663
R1809 B.n721 B.n36 256.663
R1810 B.n727 B.n36 256.663
R1811 B.n729 B.n36 256.663
R1812 B.n735 B.n36 256.663
R1813 B.n737 B.n36 256.663
R1814 B.n743 B.n36 256.663
R1815 B.n745 B.n36 256.663
R1816 B.n751 B.n36 256.663
R1817 B.n753 B.n36 256.663
R1818 B.n759 B.n36 256.663
R1819 B.n761 B.n36 256.663
R1820 B.n767 B.n36 256.663
R1821 B.n769 B.n36 256.663
R1822 B.n775 B.n36 256.663
R1823 B.n777 B.n36 256.663
R1824 B.n783 B.n36 256.663
R1825 B.n785 B.n36 256.663
R1826 B.n791 B.n36 256.663
R1827 B.n793 B.n36 256.663
R1828 B.n799 B.n36 256.663
R1829 B.n801 B.n36 256.663
R1830 B.n807 B.n36 256.663
R1831 B.n809 B.n36 256.663
R1832 B.n815 B.n36 256.663
R1833 B.n817 B.n36 256.663
R1834 B.n823 B.n36 256.663
R1835 B.n825 B.n36 256.663
R1836 B.n477 B.n142 256.663
R1837 B.n145 B.n142 256.663
R1838 B.n470 B.n142 256.663
R1839 B.n464 B.n142 256.663
R1840 B.n462 B.n142 256.663
R1841 B.n456 B.n142 256.663
R1842 B.n454 B.n142 256.663
R1843 B.n448 B.n142 256.663
R1844 B.n446 B.n142 256.663
R1845 B.n440 B.n142 256.663
R1846 B.n438 B.n142 256.663
R1847 B.n432 B.n142 256.663
R1848 B.n430 B.n142 256.663
R1849 B.n424 B.n142 256.663
R1850 B.n422 B.n142 256.663
R1851 B.n416 B.n142 256.663
R1852 B.n414 B.n142 256.663
R1853 B.n408 B.n142 256.663
R1854 B.n406 B.n142 256.663
R1855 B.n400 B.n142 256.663
R1856 B.n398 B.n142 256.663
R1857 B.n392 B.n142 256.663
R1858 B.n390 B.n142 256.663
R1859 B.n384 B.n142 256.663
R1860 B.n382 B.n142 256.663
R1861 B.n376 B.n142 256.663
R1862 B.n374 B.n142 256.663
R1863 B.n368 B.n142 256.663
R1864 B.n366 B.n142 256.663
R1865 B.n360 B.n142 256.663
R1866 B.n358 B.n142 256.663
R1867 B.n352 B.n142 256.663
R1868 B.n350 B.n142 256.663
R1869 B.n344 B.n142 256.663
R1870 B.n342 B.n142 256.663
R1871 B.n335 B.n142 256.663
R1872 B.n333 B.n142 256.663
R1873 B.n327 B.n142 256.663
R1874 B.n325 B.n142 256.663
R1875 B.n319 B.n142 256.663
R1876 B.n317 B.n142 256.663
R1877 B.n311 B.n142 256.663
R1878 B.n309 B.n142 256.663
R1879 B.n303 B.n142 256.663
R1880 B.n301 B.n142 256.663
R1881 B.n295 B.n142 256.663
R1882 B.n293 B.n142 256.663
R1883 B.n287 B.n142 256.663
R1884 B.n285 B.n142 256.663
R1885 B.n279 B.n142 256.663
R1886 B.n277 B.n142 256.663
R1887 B.n271 B.n142 256.663
R1888 B.n269 B.n142 256.663
R1889 B.n263 B.n142 256.663
R1890 B.n261 B.n142 256.663
R1891 B.n255 B.n142 256.663
R1892 B.n253 B.n142 256.663
R1893 B.n247 B.n142 256.663
R1894 B.n245 B.n142 256.663
R1895 B.n239 B.n142 256.663
R1896 B.n237 B.n142 256.663
R1897 B.n231 B.n142 256.663
R1898 B.n229 B.n142 256.663
R1899 B.n223 B.n142 256.663
R1900 B.n221 B.n142 256.663
R1901 B.n215 B.n142 256.663
R1902 B.n482 B.n137 163.367
R1903 B.n490 B.n137 163.367
R1904 B.n490 B.n135 163.367
R1905 B.n494 B.n135 163.367
R1906 B.n494 B.n129 163.367
R1907 B.n502 B.n129 163.367
R1908 B.n502 B.n127 163.367
R1909 B.n506 B.n127 163.367
R1910 B.n506 B.n121 163.367
R1911 B.n515 B.n121 163.367
R1912 B.n515 B.n119 163.367
R1913 B.n519 B.n119 163.367
R1914 B.n519 B.n114 163.367
R1915 B.n529 B.n114 163.367
R1916 B.n529 B.n112 163.367
R1917 B.n533 B.n112 163.367
R1918 B.n533 B.n2 163.367
R1919 B.n866 B.n2 163.367
R1920 B.n866 B.n3 163.367
R1921 B.n862 B.n3 163.367
R1922 B.n862 B.n8 163.367
R1923 B.n858 B.n8 163.367
R1924 B.n858 B.n10 163.367
R1925 B.n854 B.n10 163.367
R1926 B.n854 B.n15 163.367
R1927 B.n850 B.n15 163.367
R1928 B.n850 B.n17 163.367
R1929 B.n846 B.n17 163.367
R1930 B.n846 B.n23 163.367
R1931 B.n842 B.n23 163.367
R1932 B.n842 B.n25 163.367
R1933 B.n838 B.n25 163.367
R1934 B.n838 B.n30 163.367
R1935 B.n834 B.n30 163.367
R1936 B.n834 B.n32 163.367
R1937 B.n830 B.n32 163.367
R1938 B.n478 B.n476 163.367
R1939 B.n476 B.n475 163.367
R1940 B.n472 B.n471 163.367
R1941 B.n469 B.n147 163.367
R1942 B.n465 B.n463 163.367
R1943 B.n461 B.n149 163.367
R1944 B.n457 B.n455 163.367
R1945 B.n453 B.n151 163.367
R1946 B.n449 B.n447 163.367
R1947 B.n445 B.n153 163.367
R1948 B.n441 B.n439 163.367
R1949 B.n437 B.n155 163.367
R1950 B.n433 B.n431 163.367
R1951 B.n429 B.n157 163.367
R1952 B.n425 B.n423 163.367
R1953 B.n421 B.n159 163.367
R1954 B.n417 B.n415 163.367
R1955 B.n413 B.n161 163.367
R1956 B.n409 B.n407 163.367
R1957 B.n405 B.n163 163.367
R1958 B.n401 B.n399 163.367
R1959 B.n397 B.n165 163.367
R1960 B.n393 B.n391 163.367
R1961 B.n389 B.n167 163.367
R1962 B.n385 B.n383 163.367
R1963 B.n381 B.n169 163.367
R1964 B.n377 B.n375 163.367
R1965 B.n373 B.n171 163.367
R1966 B.n369 B.n367 163.367
R1967 B.n365 B.n173 163.367
R1968 B.n361 B.n359 163.367
R1969 B.n357 B.n175 163.367
R1970 B.n353 B.n351 163.367
R1971 B.n349 B.n180 163.367
R1972 B.n345 B.n343 163.367
R1973 B.n341 B.n182 163.367
R1974 B.n336 B.n334 163.367
R1975 B.n332 B.n186 163.367
R1976 B.n328 B.n326 163.367
R1977 B.n324 B.n188 163.367
R1978 B.n320 B.n318 163.367
R1979 B.n316 B.n190 163.367
R1980 B.n312 B.n310 163.367
R1981 B.n308 B.n192 163.367
R1982 B.n304 B.n302 163.367
R1983 B.n300 B.n194 163.367
R1984 B.n296 B.n294 163.367
R1985 B.n292 B.n196 163.367
R1986 B.n288 B.n286 163.367
R1987 B.n284 B.n198 163.367
R1988 B.n280 B.n278 163.367
R1989 B.n276 B.n200 163.367
R1990 B.n272 B.n270 163.367
R1991 B.n268 B.n202 163.367
R1992 B.n264 B.n262 163.367
R1993 B.n260 B.n204 163.367
R1994 B.n256 B.n254 163.367
R1995 B.n252 B.n206 163.367
R1996 B.n248 B.n246 163.367
R1997 B.n244 B.n208 163.367
R1998 B.n240 B.n238 163.367
R1999 B.n236 B.n210 163.367
R2000 B.n232 B.n230 163.367
R2001 B.n228 B.n212 163.367
R2002 B.n224 B.n222 163.367
R2003 B.n220 B.n214 163.367
R2004 B.n216 B.n141 163.367
R2005 B.n484 B.n139 163.367
R2006 B.n488 B.n139 163.367
R2007 B.n488 B.n133 163.367
R2008 B.n496 B.n133 163.367
R2009 B.n496 B.n131 163.367
R2010 B.n500 B.n131 163.367
R2011 B.n500 B.n124 163.367
R2012 B.n508 B.n124 163.367
R2013 B.n508 B.n122 163.367
R2014 B.n512 B.n122 163.367
R2015 B.n512 B.n117 163.367
R2016 B.n521 B.n117 163.367
R2017 B.n521 B.n115 163.367
R2018 B.n526 B.n115 163.367
R2019 B.n526 B.n111 163.367
R2020 B.n535 B.n111 163.367
R2021 B.n536 B.n535 163.367
R2022 B.n536 B.n5 163.367
R2023 B.n6 B.n5 163.367
R2024 B.n7 B.n6 163.367
R2025 B.n541 B.n7 163.367
R2026 B.n541 B.n12 163.367
R2027 B.n13 B.n12 163.367
R2028 B.n14 B.n13 163.367
R2029 B.n546 B.n14 163.367
R2030 B.n546 B.n19 163.367
R2031 B.n20 B.n19 163.367
R2032 B.n21 B.n20 163.367
R2033 B.n551 B.n21 163.367
R2034 B.n551 B.n26 163.367
R2035 B.n27 B.n26 163.367
R2036 B.n28 B.n27 163.367
R2037 B.n556 B.n28 163.367
R2038 B.n556 B.n33 163.367
R2039 B.n34 B.n33 163.367
R2040 B.n35 B.n34 163.367
R2041 B.n826 B.n824 163.367
R2042 B.n822 B.n39 163.367
R2043 B.n818 B.n816 163.367
R2044 B.n814 B.n41 163.367
R2045 B.n810 B.n808 163.367
R2046 B.n806 B.n43 163.367
R2047 B.n802 B.n800 163.367
R2048 B.n798 B.n45 163.367
R2049 B.n794 B.n792 163.367
R2050 B.n790 B.n47 163.367
R2051 B.n786 B.n784 163.367
R2052 B.n782 B.n49 163.367
R2053 B.n778 B.n776 163.367
R2054 B.n774 B.n51 163.367
R2055 B.n770 B.n768 163.367
R2056 B.n766 B.n53 163.367
R2057 B.n762 B.n760 163.367
R2058 B.n758 B.n55 163.367
R2059 B.n754 B.n752 163.367
R2060 B.n750 B.n57 163.367
R2061 B.n746 B.n744 163.367
R2062 B.n742 B.n59 163.367
R2063 B.n738 B.n736 163.367
R2064 B.n734 B.n61 163.367
R2065 B.n730 B.n728 163.367
R2066 B.n726 B.n63 163.367
R2067 B.n722 B.n720 163.367
R2068 B.n718 B.n65 163.367
R2069 B.n714 B.n712 163.367
R2070 B.n710 B.n67 163.367
R2071 B.n706 B.n704 163.367
R2072 B.n701 B.n700 163.367
R2073 B.n698 B.n73 163.367
R2074 B.n694 B.n692 163.367
R2075 B.n690 B.n75 163.367
R2076 B.n686 B.n684 163.367
R2077 B.n681 B.n680 163.367
R2078 B.n678 B.n81 163.367
R2079 B.n674 B.n672 163.367
R2080 B.n670 B.n83 163.367
R2081 B.n666 B.n664 163.367
R2082 B.n662 B.n85 163.367
R2083 B.n658 B.n656 163.367
R2084 B.n654 B.n87 163.367
R2085 B.n650 B.n648 163.367
R2086 B.n646 B.n89 163.367
R2087 B.n642 B.n640 163.367
R2088 B.n638 B.n91 163.367
R2089 B.n634 B.n632 163.367
R2090 B.n630 B.n93 163.367
R2091 B.n626 B.n624 163.367
R2092 B.n622 B.n95 163.367
R2093 B.n618 B.n616 163.367
R2094 B.n614 B.n97 163.367
R2095 B.n610 B.n608 163.367
R2096 B.n606 B.n99 163.367
R2097 B.n602 B.n600 163.367
R2098 B.n598 B.n101 163.367
R2099 B.n594 B.n592 163.367
R2100 B.n590 B.n103 163.367
R2101 B.n586 B.n584 163.367
R2102 B.n582 B.n105 163.367
R2103 B.n578 B.n576 163.367
R2104 B.n574 B.n107 163.367
R2105 B.n570 B.n568 163.367
R2106 B.n566 B.n109 163.367
R2107 B.n477 B.n143 71.676
R2108 B.n475 B.n145 71.676
R2109 B.n471 B.n470 71.676
R2110 B.n464 B.n147 71.676
R2111 B.n463 B.n462 71.676
R2112 B.n456 B.n149 71.676
R2113 B.n455 B.n454 71.676
R2114 B.n448 B.n151 71.676
R2115 B.n447 B.n446 71.676
R2116 B.n440 B.n153 71.676
R2117 B.n439 B.n438 71.676
R2118 B.n432 B.n155 71.676
R2119 B.n431 B.n430 71.676
R2120 B.n424 B.n157 71.676
R2121 B.n423 B.n422 71.676
R2122 B.n416 B.n159 71.676
R2123 B.n415 B.n414 71.676
R2124 B.n408 B.n161 71.676
R2125 B.n407 B.n406 71.676
R2126 B.n400 B.n163 71.676
R2127 B.n399 B.n398 71.676
R2128 B.n392 B.n165 71.676
R2129 B.n391 B.n390 71.676
R2130 B.n384 B.n167 71.676
R2131 B.n383 B.n382 71.676
R2132 B.n376 B.n169 71.676
R2133 B.n375 B.n374 71.676
R2134 B.n368 B.n171 71.676
R2135 B.n367 B.n366 71.676
R2136 B.n360 B.n173 71.676
R2137 B.n359 B.n358 71.676
R2138 B.n352 B.n175 71.676
R2139 B.n351 B.n350 71.676
R2140 B.n344 B.n180 71.676
R2141 B.n343 B.n342 71.676
R2142 B.n335 B.n182 71.676
R2143 B.n334 B.n333 71.676
R2144 B.n327 B.n186 71.676
R2145 B.n326 B.n325 71.676
R2146 B.n319 B.n188 71.676
R2147 B.n318 B.n317 71.676
R2148 B.n311 B.n190 71.676
R2149 B.n310 B.n309 71.676
R2150 B.n303 B.n192 71.676
R2151 B.n302 B.n301 71.676
R2152 B.n295 B.n194 71.676
R2153 B.n294 B.n293 71.676
R2154 B.n287 B.n196 71.676
R2155 B.n286 B.n285 71.676
R2156 B.n279 B.n198 71.676
R2157 B.n278 B.n277 71.676
R2158 B.n271 B.n200 71.676
R2159 B.n270 B.n269 71.676
R2160 B.n263 B.n202 71.676
R2161 B.n262 B.n261 71.676
R2162 B.n255 B.n204 71.676
R2163 B.n254 B.n253 71.676
R2164 B.n247 B.n206 71.676
R2165 B.n246 B.n245 71.676
R2166 B.n239 B.n208 71.676
R2167 B.n238 B.n237 71.676
R2168 B.n231 B.n210 71.676
R2169 B.n230 B.n229 71.676
R2170 B.n223 B.n212 71.676
R2171 B.n222 B.n221 71.676
R2172 B.n215 B.n214 71.676
R2173 B.n825 B.n37 71.676
R2174 B.n824 B.n823 71.676
R2175 B.n817 B.n39 71.676
R2176 B.n816 B.n815 71.676
R2177 B.n809 B.n41 71.676
R2178 B.n808 B.n807 71.676
R2179 B.n801 B.n43 71.676
R2180 B.n800 B.n799 71.676
R2181 B.n793 B.n45 71.676
R2182 B.n792 B.n791 71.676
R2183 B.n785 B.n47 71.676
R2184 B.n784 B.n783 71.676
R2185 B.n777 B.n49 71.676
R2186 B.n776 B.n775 71.676
R2187 B.n769 B.n51 71.676
R2188 B.n768 B.n767 71.676
R2189 B.n761 B.n53 71.676
R2190 B.n760 B.n759 71.676
R2191 B.n753 B.n55 71.676
R2192 B.n752 B.n751 71.676
R2193 B.n745 B.n57 71.676
R2194 B.n744 B.n743 71.676
R2195 B.n737 B.n59 71.676
R2196 B.n736 B.n735 71.676
R2197 B.n729 B.n61 71.676
R2198 B.n728 B.n727 71.676
R2199 B.n721 B.n63 71.676
R2200 B.n720 B.n719 71.676
R2201 B.n713 B.n65 71.676
R2202 B.n712 B.n711 71.676
R2203 B.n705 B.n67 71.676
R2204 B.n704 B.n71 71.676
R2205 B.n700 B.n699 71.676
R2206 B.n693 B.n73 71.676
R2207 B.n692 B.n691 71.676
R2208 B.n685 B.n75 71.676
R2209 B.n684 B.n79 71.676
R2210 B.n680 B.n679 71.676
R2211 B.n673 B.n81 71.676
R2212 B.n672 B.n671 71.676
R2213 B.n665 B.n83 71.676
R2214 B.n664 B.n663 71.676
R2215 B.n657 B.n85 71.676
R2216 B.n656 B.n655 71.676
R2217 B.n649 B.n87 71.676
R2218 B.n648 B.n647 71.676
R2219 B.n641 B.n89 71.676
R2220 B.n640 B.n639 71.676
R2221 B.n633 B.n91 71.676
R2222 B.n632 B.n631 71.676
R2223 B.n625 B.n93 71.676
R2224 B.n624 B.n623 71.676
R2225 B.n617 B.n95 71.676
R2226 B.n616 B.n615 71.676
R2227 B.n609 B.n97 71.676
R2228 B.n608 B.n607 71.676
R2229 B.n601 B.n99 71.676
R2230 B.n600 B.n599 71.676
R2231 B.n593 B.n101 71.676
R2232 B.n592 B.n591 71.676
R2233 B.n585 B.n103 71.676
R2234 B.n584 B.n583 71.676
R2235 B.n577 B.n105 71.676
R2236 B.n576 B.n575 71.676
R2237 B.n569 B.n107 71.676
R2238 B.n568 B.n567 71.676
R2239 B.n561 B.n109 71.676
R2240 B.n562 B.n561 71.676
R2241 B.n567 B.n566 71.676
R2242 B.n570 B.n569 71.676
R2243 B.n575 B.n574 71.676
R2244 B.n578 B.n577 71.676
R2245 B.n583 B.n582 71.676
R2246 B.n586 B.n585 71.676
R2247 B.n591 B.n590 71.676
R2248 B.n594 B.n593 71.676
R2249 B.n599 B.n598 71.676
R2250 B.n602 B.n601 71.676
R2251 B.n607 B.n606 71.676
R2252 B.n610 B.n609 71.676
R2253 B.n615 B.n614 71.676
R2254 B.n618 B.n617 71.676
R2255 B.n623 B.n622 71.676
R2256 B.n626 B.n625 71.676
R2257 B.n631 B.n630 71.676
R2258 B.n634 B.n633 71.676
R2259 B.n639 B.n638 71.676
R2260 B.n642 B.n641 71.676
R2261 B.n647 B.n646 71.676
R2262 B.n650 B.n649 71.676
R2263 B.n655 B.n654 71.676
R2264 B.n658 B.n657 71.676
R2265 B.n663 B.n662 71.676
R2266 B.n666 B.n665 71.676
R2267 B.n671 B.n670 71.676
R2268 B.n674 B.n673 71.676
R2269 B.n679 B.n678 71.676
R2270 B.n681 B.n79 71.676
R2271 B.n686 B.n685 71.676
R2272 B.n691 B.n690 71.676
R2273 B.n694 B.n693 71.676
R2274 B.n699 B.n698 71.676
R2275 B.n701 B.n71 71.676
R2276 B.n706 B.n705 71.676
R2277 B.n711 B.n710 71.676
R2278 B.n714 B.n713 71.676
R2279 B.n719 B.n718 71.676
R2280 B.n722 B.n721 71.676
R2281 B.n727 B.n726 71.676
R2282 B.n730 B.n729 71.676
R2283 B.n735 B.n734 71.676
R2284 B.n738 B.n737 71.676
R2285 B.n743 B.n742 71.676
R2286 B.n746 B.n745 71.676
R2287 B.n751 B.n750 71.676
R2288 B.n754 B.n753 71.676
R2289 B.n759 B.n758 71.676
R2290 B.n762 B.n761 71.676
R2291 B.n767 B.n766 71.676
R2292 B.n770 B.n769 71.676
R2293 B.n775 B.n774 71.676
R2294 B.n778 B.n777 71.676
R2295 B.n783 B.n782 71.676
R2296 B.n786 B.n785 71.676
R2297 B.n791 B.n790 71.676
R2298 B.n794 B.n793 71.676
R2299 B.n799 B.n798 71.676
R2300 B.n802 B.n801 71.676
R2301 B.n807 B.n806 71.676
R2302 B.n810 B.n809 71.676
R2303 B.n815 B.n814 71.676
R2304 B.n818 B.n817 71.676
R2305 B.n823 B.n822 71.676
R2306 B.n826 B.n825 71.676
R2307 B.n478 B.n477 71.676
R2308 B.n472 B.n145 71.676
R2309 B.n470 B.n469 71.676
R2310 B.n465 B.n464 71.676
R2311 B.n462 B.n461 71.676
R2312 B.n457 B.n456 71.676
R2313 B.n454 B.n453 71.676
R2314 B.n449 B.n448 71.676
R2315 B.n446 B.n445 71.676
R2316 B.n441 B.n440 71.676
R2317 B.n438 B.n437 71.676
R2318 B.n433 B.n432 71.676
R2319 B.n430 B.n429 71.676
R2320 B.n425 B.n424 71.676
R2321 B.n422 B.n421 71.676
R2322 B.n417 B.n416 71.676
R2323 B.n414 B.n413 71.676
R2324 B.n409 B.n408 71.676
R2325 B.n406 B.n405 71.676
R2326 B.n401 B.n400 71.676
R2327 B.n398 B.n397 71.676
R2328 B.n393 B.n392 71.676
R2329 B.n390 B.n389 71.676
R2330 B.n385 B.n384 71.676
R2331 B.n382 B.n381 71.676
R2332 B.n377 B.n376 71.676
R2333 B.n374 B.n373 71.676
R2334 B.n369 B.n368 71.676
R2335 B.n366 B.n365 71.676
R2336 B.n361 B.n360 71.676
R2337 B.n358 B.n357 71.676
R2338 B.n353 B.n352 71.676
R2339 B.n350 B.n349 71.676
R2340 B.n345 B.n344 71.676
R2341 B.n342 B.n341 71.676
R2342 B.n336 B.n335 71.676
R2343 B.n333 B.n332 71.676
R2344 B.n328 B.n327 71.676
R2345 B.n325 B.n324 71.676
R2346 B.n320 B.n319 71.676
R2347 B.n317 B.n316 71.676
R2348 B.n312 B.n311 71.676
R2349 B.n309 B.n308 71.676
R2350 B.n304 B.n303 71.676
R2351 B.n301 B.n300 71.676
R2352 B.n296 B.n295 71.676
R2353 B.n293 B.n292 71.676
R2354 B.n288 B.n287 71.676
R2355 B.n285 B.n284 71.676
R2356 B.n280 B.n279 71.676
R2357 B.n277 B.n276 71.676
R2358 B.n272 B.n271 71.676
R2359 B.n269 B.n268 71.676
R2360 B.n264 B.n263 71.676
R2361 B.n261 B.n260 71.676
R2362 B.n256 B.n255 71.676
R2363 B.n253 B.n252 71.676
R2364 B.n248 B.n247 71.676
R2365 B.n245 B.n244 71.676
R2366 B.n240 B.n239 71.676
R2367 B.n237 B.n236 71.676
R2368 B.n232 B.n231 71.676
R2369 B.n229 B.n228 71.676
R2370 B.n224 B.n223 71.676
R2371 B.n221 B.n220 71.676
R2372 B.n216 B.n215 71.676
R2373 B.n338 B.n184 59.5399
R2374 B.n178 B.n177 59.5399
R2375 B.n70 B.n69 59.5399
R2376 B.n78 B.n77 59.5399
R2377 B.n483 B.n142 55.0119
R2378 B.n831 B.n36 55.0119
R2379 B.n483 B.n138 30.916
R2380 B.n489 B.n138 30.916
R2381 B.n489 B.n134 30.916
R2382 B.n495 B.n134 30.916
R2383 B.n501 B.n130 30.916
R2384 B.n501 B.n125 30.916
R2385 B.n507 B.n125 30.916
R2386 B.n507 B.n126 30.916
R2387 B.n514 B.n513 30.916
R2388 B.n520 B.n118 30.916
R2389 B.n528 B.n527 30.916
R2390 B.n534 B.n4 30.916
R2391 B.n865 B.n4 30.916
R2392 B.n865 B.n864 30.916
R2393 B.n864 B.n863 30.916
R2394 B.n857 B.n11 30.916
R2395 B.n856 B.n855 30.916
R2396 B.n849 B.n18 30.916
R2397 B.n848 B.n847 30.916
R2398 B.n847 B.n22 30.916
R2399 B.n841 B.n22 30.916
R2400 B.n841 B.n840 30.916
R2401 B.n839 B.n29 30.916
R2402 B.n833 B.n29 30.916
R2403 B.n833 B.n832 30.916
R2404 B.n832 B.n831 30.916
R2405 B.n563 B.n560 29.5029
R2406 B.n829 B.n828 29.5029
R2407 B.n485 B.n140 29.5029
R2408 B.n481 B.n480 29.5029
R2409 B.t9 B.n130 20.9139
R2410 B.n840 B.t13 20.9139
R2411 B.n534 B.t3 18.1861
R2412 B.n863 B.t0 18.1861
R2413 B B.n867 18.0485
R2414 B.n528 B.t4 17.2768
R2415 B.n857 B.t1 17.2768
R2416 B.n520 B.t5 16.3675
R2417 B.n855 B.t6 16.3675
R2418 B.n126 B.t7 15.4582
R2419 B.n514 B.t7 15.4582
R2420 B.n849 B.t2 15.4582
R2421 B.t2 B.n848 15.4582
R2422 B.n513 B.t5 14.549
R2423 B.n18 B.t6 14.549
R2424 B.n118 B.t4 13.6397
R2425 B.t1 B.n856 13.6397
R2426 B.n184 B.n183 12.9944
R2427 B.n177 B.n176 12.9944
R2428 B.n69 B.n68 12.9944
R2429 B.n77 B.n76 12.9944
R2430 B.n527 B.t3 12.7304
R2431 B.n11 B.t0 12.7304
R2432 B.n828 B.n827 10.6151
R2433 B.n827 B.n38 10.6151
R2434 B.n821 B.n38 10.6151
R2435 B.n821 B.n820 10.6151
R2436 B.n820 B.n819 10.6151
R2437 B.n819 B.n40 10.6151
R2438 B.n813 B.n40 10.6151
R2439 B.n813 B.n812 10.6151
R2440 B.n812 B.n811 10.6151
R2441 B.n811 B.n42 10.6151
R2442 B.n805 B.n42 10.6151
R2443 B.n805 B.n804 10.6151
R2444 B.n804 B.n803 10.6151
R2445 B.n803 B.n44 10.6151
R2446 B.n797 B.n44 10.6151
R2447 B.n797 B.n796 10.6151
R2448 B.n796 B.n795 10.6151
R2449 B.n795 B.n46 10.6151
R2450 B.n789 B.n46 10.6151
R2451 B.n789 B.n788 10.6151
R2452 B.n788 B.n787 10.6151
R2453 B.n787 B.n48 10.6151
R2454 B.n781 B.n48 10.6151
R2455 B.n781 B.n780 10.6151
R2456 B.n780 B.n779 10.6151
R2457 B.n779 B.n50 10.6151
R2458 B.n773 B.n50 10.6151
R2459 B.n773 B.n772 10.6151
R2460 B.n772 B.n771 10.6151
R2461 B.n771 B.n52 10.6151
R2462 B.n765 B.n52 10.6151
R2463 B.n765 B.n764 10.6151
R2464 B.n764 B.n763 10.6151
R2465 B.n763 B.n54 10.6151
R2466 B.n757 B.n54 10.6151
R2467 B.n757 B.n756 10.6151
R2468 B.n756 B.n755 10.6151
R2469 B.n755 B.n56 10.6151
R2470 B.n749 B.n56 10.6151
R2471 B.n749 B.n748 10.6151
R2472 B.n748 B.n747 10.6151
R2473 B.n747 B.n58 10.6151
R2474 B.n741 B.n58 10.6151
R2475 B.n741 B.n740 10.6151
R2476 B.n740 B.n739 10.6151
R2477 B.n739 B.n60 10.6151
R2478 B.n733 B.n60 10.6151
R2479 B.n733 B.n732 10.6151
R2480 B.n732 B.n731 10.6151
R2481 B.n731 B.n62 10.6151
R2482 B.n725 B.n62 10.6151
R2483 B.n725 B.n724 10.6151
R2484 B.n724 B.n723 10.6151
R2485 B.n723 B.n64 10.6151
R2486 B.n717 B.n64 10.6151
R2487 B.n717 B.n716 10.6151
R2488 B.n716 B.n715 10.6151
R2489 B.n715 B.n66 10.6151
R2490 B.n709 B.n66 10.6151
R2491 B.n709 B.n708 10.6151
R2492 B.n708 B.n707 10.6151
R2493 B.n703 B.n702 10.6151
R2494 B.n702 B.n72 10.6151
R2495 B.n697 B.n72 10.6151
R2496 B.n697 B.n696 10.6151
R2497 B.n696 B.n695 10.6151
R2498 B.n695 B.n74 10.6151
R2499 B.n689 B.n74 10.6151
R2500 B.n689 B.n688 10.6151
R2501 B.n688 B.n687 10.6151
R2502 B.n683 B.n682 10.6151
R2503 B.n682 B.n80 10.6151
R2504 B.n677 B.n80 10.6151
R2505 B.n677 B.n676 10.6151
R2506 B.n676 B.n675 10.6151
R2507 B.n675 B.n82 10.6151
R2508 B.n669 B.n82 10.6151
R2509 B.n669 B.n668 10.6151
R2510 B.n668 B.n667 10.6151
R2511 B.n667 B.n84 10.6151
R2512 B.n661 B.n84 10.6151
R2513 B.n661 B.n660 10.6151
R2514 B.n660 B.n659 10.6151
R2515 B.n659 B.n86 10.6151
R2516 B.n653 B.n86 10.6151
R2517 B.n653 B.n652 10.6151
R2518 B.n652 B.n651 10.6151
R2519 B.n651 B.n88 10.6151
R2520 B.n645 B.n88 10.6151
R2521 B.n645 B.n644 10.6151
R2522 B.n644 B.n643 10.6151
R2523 B.n643 B.n90 10.6151
R2524 B.n637 B.n90 10.6151
R2525 B.n637 B.n636 10.6151
R2526 B.n636 B.n635 10.6151
R2527 B.n635 B.n92 10.6151
R2528 B.n629 B.n92 10.6151
R2529 B.n629 B.n628 10.6151
R2530 B.n628 B.n627 10.6151
R2531 B.n627 B.n94 10.6151
R2532 B.n621 B.n94 10.6151
R2533 B.n621 B.n620 10.6151
R2534 B.n620 B.n619 10.6151
R2535 B.n619 B.n96 10.6151
R2536 B.n613 B.n96 10.6151
R2537 B.n613 B.n612 10.6151
R2538 B.n612 B.n611 10.6151
R2539 B.n611 B.n98 10.6151
R2540 B.n605 B.n98 10.6151
R2541 B.n605 B.n604 10.6151
R2542 B.n604 B.n603 10.6151
R2543 B.n603 B.n100 10.6151
R2544 B.n597 B.n100 10.6151
R2545 B.n597 B.n596 10.6151
R2546 B.n596 B.n595 10.6151
R2547 B.n595 B.n102 10.6151
R2548 B.n589 B.n102 10.6151
R2549 B.n589 B.n588 10.6151
R2550 B.n588 B.n587 10.6151
R2551 B.n587 B.n104 10.6151
R2552 B.n581 B.n104 10.6151
R2553 B.n581 B.n580 10.6151
R2554 B.n580 B.n579 10.6151
R2555 B.n579 B.n106 10.6151
R2556 B.n573 B.n106 10.6151
R2557 B.n573 B.n572 10.6151
R2558 B.n572 B.n571 10.6151
R2559 B.n571 B.n108 10.6151
R2560 B.n565 B.n108 10.6151
R2561 B.n565 B.n564 10.6151
R2562 B.n564 B.n563 10.6151
R2563 B.n486 B.n485 10.6151
R2564 B.n487 B.n486 10.6151
R2565 B.n487 B.n132 10.6151
R2566 B.n497 B.n132 10.6151
R2567 B.n498 B.n497 10.6151
R2568 B.n499 B.n498 10.6151
R2569 B.n499 B.n123 10.6151
R2570 B.n509 B.n123 10.6151
R2571 B.n510 B.n509 10.6151
R2572 B.n511 B.n510 10.6151
R2573 B.n511 B.n116 10.6151
R2574 B.n522 B.n116 10.6151
R2575 B.n523 B.n522 10.6151
R2576 B.n525 B.n523 10.6151
R2577 B.n525 B.n524 10.6151
R2578 B.n524 B.n110 10.6151
R2579 B.n537 B.n110 10.6151
R2580 B.n538 B.n537 10.6151
R2581 B.n539 B.n538 10.6151
R2582 B.n540 B.n539 10.6151
R2583 B.n542 B.n540 10.6151
R2584 B.n543 B.n542 10.6151
R2585 B.n544 B.n543 10.6151
R2586 B.n545 B.n544 10.6151
R2587 B.n547 B.n545 10.6151
R2588 B.n548 B.n547 10.6151
R2589 B.n549 B.n548 10.6151
R2590 B.n550 B.n549 10.6151
R2591 B.n552 B.n550 10.6151
R2592 B.n553 B.n552 10.6151
R2593 B.n554 B.n553 10.6151
R2594 B.n555 B.n554 10.6151
R2595 B.n557 B.n555 10.6151
R2596 B.n558 B.n557 10.6151
R2597 B.n559 B.n558 10.6151
R2598 B.n560 B.n559 10.6151
R2599 B.n480 B.n479 10.6151
R2600 B.n479 B.n144 10.6151
R2601 B.n474 B.n144 10.6151
R2602 B.n474 B.n473 10.6151
R2603 B.n473 B.n146 10.6151
R2604 B.n468 B.n146 10.6151
R2605 B.n468 B.n467 10.6151
R2606 B.n467 B.n466 10.6151
R2607 B.n466 B.n148 10.6151
R2608 B.n460 B.n148 10.6151
R2609 B.n460 B.n459 10.6151
R2610 B.n459 B.n458 10.6151
R2611 B.n458 B.n150 10.6151
R2612 B.n452 B.n150 10.6151
R2613 B.n452 B.n451 10.6151
R2614 B.n451 B.n450 10.6151
R2615 B.n450 B.n152 10.6151
R2616 B.n444 B.n152 10.6151
R2617 B.n444 B.n443 10.6151
R2618 B.n443 B.n442 10.6151
R2619 B.n442 B.n154 10.6151
R2620 B.n436 B.n154 10.6151
R2621 B.n436 B.n435 10.6151
R2622 B.n435 B.n434 10.6151
R2623 B.n434 B.n156 10.6151
R2624 B.n428 B.n156 10.6151
R2625 B.n428 B.n427 10.6151
R2626 B.n427 B.n426 10.6151
R2627 B.n426 B.n158 10.6151
R2628 B.n420 B.n158 10.6151
R2629 B.n420 B.n419 10.6151
R2630 B.n419 B.n418 10.6151
R2631 B.n418 B.n160 10.6151
R2632 B.n412 B.n160 10.6151
R2633 B.n412 B.n411 10.6151
R2634 B.n411 B.n410 10.6151
R2635 B.n410 B.n162 10.6151
R2636 B.n404 B.n162 10.6151
R2637 B.n404 B.n403 10.6151
R2638 B.n403 B.n402 10.6151
R2639 B.n402 B.n164 10.6151
R2640 B.n396 B.n164 10.6151
R2641 B.n396 B.n395 10.6151
R2642 B.n395 B.n394 10.6151
R2643 B.n394 B.n166 10.6151
R2644 B.n388 B.n166 10.6151
R2645 B.n388 B.n387 10.6151
R2646 B.n387 B.n386 10.6151
R2647 B.n386 B.n168 10.6151
R2648 B.n380 B.n168 10.6151
R2649 B.n380 B.n379 10.6151
R2650 B.n379 B.n378 10.6151
R2651 B.n378 B.n170 10.6151
R2652 B.n372 B.n170 10.6151
R2653 B.n372 B.n371 10.6151
R2654 B.n371 B.n370 10.6151
R2655 B.n370 B.n172 10.6151
R2656 B.n364 B.n172 10.6151
R2657 B.n364 B.n363 10.6151
R2658 B.n363 B.n362 10.6151
R2659 B.n362 B.n174 10.6151
R2660 B.n356 B.n355 10.6151
R2661 B.n355 B.n354 10.6151
R2662 B.n354 B.n179 10.6151
R2663 B.n348 B.n179 10.6151
R2664 B.n348 B.n347 10.6151
R2665 B.n347 B.n346 10.6151
R2666 B.n346 B.n181 10.6151
R2667 B.n340 B.n181 10.6151
R2668 B.n340 B.n339 10.6151
R2669 B.n337 B.n185 10.6151
R2670 B.n331 B.n185 10.6151
R2671 B.n331 B.n330 10.6151
R2672 B.n330 B.n329 10.6151
R2673 B.n329 B.n187 10.6151
R2674 B.n323 B.n187 10.6151
R2675 B.n323 B.n322 10.6151
R2676 B.n322 B.n321 10.6151
R2677 B.n321 B.n189 10.6151
R2678 B.n315 B.n189 10.6151
R2679 B.n315 B.n314 10.6151
R2680 B.n314 B.n313 10.6151
R2681 B.n313 B.n191 10.6151
R2682 B.n307 B.n191 10.6151
R2683 B.n307 B.n306 10.6151
R2684 B.n306 B.n305 10.6151
R2685 B.n305 B.n193 10.6151
R2686 B.n299 B.n193 10.6151
R2687 B.n299 B.n298 10.6151
R2688 B.n298 B.n297 10.6151
R2689 B.n297 B.n195 10.6151
R2690 B.n291 B.n195 10.6151
R2691 B.n291 B.n290 10.6151
R2692 B.n290 B.n289 10.6151
R2693 B.n289 B.n197 10.6151
R2694 B.n283 B.n197 10.6151
R2695 B.n283 B.n282 10.6151
R2696 B.n282 B.n281 10.6151
R2697 B.n281 B.n199 10.6151
R2698 B.n275 B.n199 10.6151
R2699 B.n275 B.n274 10.6151
R2700 B.n274 B.n273 10.6151
R2701 B.n273 B.n201 10.6151
R2702 B.n267 B.n201 10.6151
R2703 B.n267 B.n266 10.6151
R2704 B.n266 B.n265 10.6151
R2705 B.n265 B.n203 10.6151
R2706 B.n259 B.n203 10.6151
R2707 B.n259 B.n258 10.6151
R2708 B.n258 B.n257 10.6151
R2709 B.n257 B.n205 10.6151
R2710 B.n251 B.n205 10.6151
R2711 B.n251 B.n250 10.6151
R2712 B.n250 B.n249 10.6151
R2713 B.n249 B.n207 10.6151
R2714 B.n243 B.n207 10.6151
R2715 B.n243 B.n242 10.6151
R2716 B.n242 B.n241 10.6151
R2717 B.n241 B.n209 10.6151
R2718 B.n235 B.n209 10.6151
R2719 B.n235 B.n234 10.6151
R2720 B.n234 B.n233 10.6151
R2721 B.n233 B.n211 10.6151
R2722 B.n227 B.n211 10.6151
R2723 B.n227 B.n226 10.6151
R2724 B.n226 B.n225 10.6151
R2725 B.n225 B.n213 10.6151
R2726 B.n219 B.n213 10.6151
R2727 B.n219 B.n218 10.6151
R2728 B.n218 B.n217 10.6151
R2729 B.n217 B.n140 10.6151
R2730 B.n481 B.n136 10.6151
R2731 B.n491 B.n136 10.6151
R2732 B.n492 B.n491 10.6151
R2733 B.n493 B.n492 10.6151
R2734 B.n493 B.n128 10.6151
R2735 B.n503 B.n128 10.6151
R2736 B.n504 B.n503 10.6151
R2737 B.n505 B.n504 10.6151
R2738 B.n505 B.n120 10.6151
R2739 B.n516 B.n120 10.6151
R2740 B.n517 B.n516 10.6151
R2741 B.n518 B.n517 10.6151
R2742 B.n518 B.n113 10.6151
R2743 B.n530 B.n113 10.6151
R2744 B.n531 B.n530 10.6151
R2745 B.n532 B.n531 10.6151
R2746 B.n532 B.n0 10.6151
R2747 B.n861 B.n1 10.6151
R2748 B.n861 B.n860 10.6151
R2749 B.n860 B.n859 10.6151
R2750 B.n859 B.n9 10.6151
R2751 B.n853 B.n9 10.6151
R2752 B.n853 B.n852 10.6151
R2753 B.n852 B.n851 10.6151
R2754 B.n851 B.n16 10.6151
R2755 B.n845 B.n16 10.6151
R2756 B.n845 B.n844 10.6151
R2757 B.n844 B.n843 10.6151
R2758 B.n843 B.n24 10.6151
R2759 B.n837 B.n24 10.6151
R2760 B.n837 B.n836 10.6151
R2761 B.n836 B.n835 10.6151
R2762 B.n835 B.n31 10.6151
R2763 B.n829 B.n31 10.6151
R2764 B.n495 B.t9 10.0026
R2765 B.t13 B.n839 10.0026
R2766 B.n707 B.n70 9.36635
R2767 B.n683 B.n78 9.36635
R2768 B.n178 B.n174 9.36635
R2769 B.n338 B.n337 9.36635
R2770 B.n867 B.n0 2.81026
R2771 B.n867 B.n1 2.81026
R2772 B.n703 B.n70 1.24928
R2773 B.n687 B.n78 1.24928
R2774 B.n356 B.n178 1.24928
R2775 B.n339 B.n338 1.24928
R2776 VP.n3 VP.t1 1486.58
R2777 VP.n12 VP.t5 1470.47
R2778 VP.n1 VP.t6 1470.47
R2779 VP.n6 VP.t2 1470.47
R2780 VP.n10 VP.t7 1458.05
R2781 VP.n11 VP.t3 1458.05
R2782 VP.n5 VP.t4 1458.05
R2783 VP.n4 VP.t0 1458.05
R2784 VP.n13 VP.n12 161.3
R2785 VP.n5 VP.n2 161.3
R2786 VP.n7 VP.n6 161.3
R2787 VP.n11 VP.n0 161.3
R2788 VP.n10 VP.n9 161.3
R2789 VP.n8 VP.n1 161.3
R2790 VP.n3 VP.n2 72.8343
R2791 VP.n11 VP.n10 48.2005
R2792 VP.n5 VP.n4 48.2005
R2793 VP.n8 VP.n7 45.6217
R2794 VP.n10 VP.n1 35.7853
R2795 VP.n12 VP.n11 35.7853
R2796 VP.n6 VP.n5 35.7853
R2797 VP.n4 VP.n3 16.0984
R2798 VP.n7 VP.n2 0.189894
R2799 VP.n9 VP.n8 0.189894
R2800 VP.n9 VP.n0 0.189894
R2801 VP.n13 VP.n0 0.189894
R2802 VP VP.n13 0.0516364
R2803 VDD1 VDD1.n0 60.1932
R2804 VDD1.n3 VDD1.n2 60.0797
R2805 VDD1.n3 VDD1.n1 60.0797
R2806 VDD1.n5 VDD1.n4 59.846
R2807 VDD1.n5 VDD1.n3 43.2078
R2808 VDD1.n4 VDD1.t3 1.04701
R2809 VDD1.n4 VDD1.t5 1.04701
R2810 VDD1.n0 VDD1.t6 1.04701
R2811 VDD1.n0 VDD1.t7 1.04701
R2812 VDD1.n2 VDD1.t4 1.04701
R2813 VDD1.n2 VDD1.t2 1.04701
R2814 VDD1.n1 VDD1.t1 1.04701
R2815 VDD1.n1 VDD1.t0 1.04701
R2816 VDD1 VDD1.n5 0.231103
C0 VDD2 VN 5.50508f
C1 VDD1 VP 5.63637f
C2 VP VTAIL 4.82677f
C3 VDD1 VTAIL 23.403101f
C4 VDD2 VP 0.278563f
C5 VP VN 6.18262f
C6 VDD1 VDD2 0.649374f
C7 VDD2 VTAIL 23.4424f
C8 VDD1 VN 0.147023f
C9 VN VTAIL 4.81267f
C10 VDD2 B 3.716774f
C11 VDD1 B 3.907419f
C12 VTAIL B 12.298511f
C13 VN B 8.36322f
C14 VP B 5.691056f
C15 VDD1.t6 B 0.489207f
C16 VDD1.t7 B 0.489207f
C17 VDD1.n0 B 4.46557f
C18 VDD1.t1 B 0.489207f
C19 VDD1.t0 B 0.489207f
C20 VDD1.n1 B 4.46481f
C21 VDD1.t4 B 0.489207f
C22 VDD1.t2 B 0.489207f
C23 VDD1.n2 B 4.46481f
C24 VDD1.n3 B 3.20953f
C25 VDD1.t3 B 0.489207f
C26 VDD1.t5 B 0.489207f
C27 VDD1.n4 B 4.46333f
C28 VDD1.n5 B 3.57417f
C29 VP.n0 B 0.054591f
C30 VP.t6 B 0.998561f
C31 VP.n1 B 0.380222f
C32 VP.n2 B 0.175162f
C33 VP.t4 B 0.995428f
C34 VP.t0 B 0.995428f
C35 VP.t1 B 1.00268f
C36 VP.n3 B 0.376492f
C37 VP.n4 B 0.38874f
C38 VP.n5 B 0.38874f
C39 VP.t2 B 0.998561f
C40 VP.n6 B 0.380222f
C41 VP.n7 B 2.57709f
C42 VP.n8 B 2.61999f
C43 VP.n9 B 0.054591f
C44 VP.t7 B 0.995428f
C45 VP.n10 B 0.38874f
C46 VP.t3 B 0.995428f
C47 VP.n11 B 0.38874f
C48 VP.t5 B 0.998561f
C49 VP.n12 B 0.380222f
C50 VP.n13 B 0.042306f
C51 VDD2.t1 B 0.48956f
C52 VDD2.t4 B 0.48956f
C53 VDD2.n0 B 4.46803f
C54 VDD2.t5 B 0.48956f
C55 VDD2.t3 B 0.48956f
C56 VDD2.n1 B 4.46803f
C57 VDD2.n2 B 3.14217f
C58 VDD2.t0 B 0.48956f
C59 VDD2.t7 B 0.48956f
C60 VDD2.n3 B 4.46657f
C61 VDD2.n4 B 3.53775f
C62 VDD2.t6 B 0.48956f
C63 VDD2.t2 B 0.48956f
C64 VDD2.n5 B 4.46799f
C65 VTAIL.t11 B 0.340702f
C66 VTAIL.t15 B 0.340702f
C67 VTAIL.n0 B 3.03617f
C68 VTAIL.n1 B 0.279349f
C69 VTAIL.n2 B 0.03203f
C70 VTAIL.n3 B 0.022788f
C71 VTAIL.n4 B 0.012245f
C72 VTAIL.n5 B 0.028943f
C73 VTAIL.n6 B 0.012965f
C74 VTAIL.n7 B 0.022788f
C75 VTAIL.n8 B 0.012245f
C76 VTAIL.n9 B 0.028943f
C77 VTAIL.n10 B 0.012965f
C78 VTAIL.n11 B 0.022788f
C79 VTAIL.n12 B 0.012245f
C80 VTAIL.n13 B 0.028943f
C81 VTAIL.n14 B 0.012965f
C82 VTAIL.n15 B 0.022788f
C83 VTAIL.n16 B 0.012245f
C84 VTAIL.n17 B 0.028943f
C85 VTAIL.n18 B 0.012965f
C86 VTAIL.n19 B 0.022788f
C87 VTAIL.n20 B 0.012245f
C88 VTAIL.n21 B 0.028943f
C89 VTAIL.n22 B 0.012965f
C90 VTAIL.n23 B 0.022788f
C91 VTAIL.n24 B 0.012245f
C92 VTAIL.n25 B 0.028943f
C93 VTAIL.n26 B 0.012965f
C94 VTAIL.n27 B 0.022788f
C95 VTAIL.n28 B 0.012245f
C96 VTAIL.n29 B 0.028943f
C97 VTAIL.n30 B 0.012965f
C98 VTAIL.n31 B 0.022788f
C99 VTAIL.n32 B 0.012245f
C100 VTAIL.n33 B 0.028943f
C101 VTAIL.n34 B 0.012965f
C102 VTAIL.n35 B 0.171022f
C103 VTAIL.t10 B 0.04803f
C104 VTAIL.n36 B 0.021707f
C105 VTAIL.n37 B 0.017098f
C106 VTAIL.n38 B 0.012245f
C107 VTAIL.n39 B 1.89199f
C108 VTAIL.n40 B 0.022788f
C109 VTAIL.n41 B 0.012245f
C110 VTAIL.n42 B 0.012965f
C111 VTAIL.n43 B 0.028943f
C112 VTAIL.n44 B 0.028943f
C113 VTAIL.n45 B 0.012965f
C114 VTAIL.n46 B 0.012245f
C115 VTAIL.n47 B 0.022788f
C116 VTAIL.n48 B 0.022788f
C117 VTAIL.n49 B 0.012245f
C118 VTAIL.n50 B 0.012965f
C119 VTAIL.n51 B 0.028943f
C120 VTAIL.n52 B 0.028943f
C121 VTAIL.n53 B 0.012965f
C122 VTAIL.n54 B 0.012245f
C123 VTAIL.n55 B 0.022788f
C124 VTAIL.n56 B 0.022788f
C125 VTAIL.n57 B 0.012245f
C126 VTAIL.n58 B 0.012965f
C127 VTAIL.n59 B 0.028943f
C128 VTAIL.n60 B 0.028943f
C129 VTAIL.n61 B 0.012965f
C130 VTAIL.n62 B 0.012245f
C131 VTAIL.n63 B 0.022788f
C132 VTAIL.n64 B 0.022788f
C133 VTAIL.n65 B 0.012245f
C134 VTAIL.n66 B 0.012965f
C135 VTAIL.n67 B 0.028943f
C136 VTAIL.n68 B 0.028943f
C137 VTAIL.n69 B 0.012965f
C138 VTAIL.n70 B 0.012245f
C139 VTAIL.n71 B 0.022788f
C140 VTAIL.n72 B 0.022788f
C141 VTAIL.n73 B 0.012245f
C142 VTAIL.n74 B 0.012965f
C143 VTAIL.n75 B 0.028943f
C144 VTAIL.n76 B 0.028943f
C145 VTAIL.n77 B 0.028943f
C146 VTAIL.n78 B 0.012965f
C147 VTAIL.n79 B 0.012245f
C148 VTAIL.n80 B 0.022788f
C149 VTAIL.n81 B 0.022788f
C150 VTAIL.n82 B 0.012245f
C151 VTAIL.n83 B 0.012605f
C152 VTAIL.n84 B 0.012605f
C153 VTAIL.n85 B 0.028943f
C154 VTAIL.n86 B 0.028943f
C155 VTAIL.n87 B 0.012965f
C156 VTAIL.n88 B 0.012245f
C157 VTAIL.n89 B 0.022788f
C158 VTAIL.n90 B 0.022788f
C159 VTAIL.n91 B 0.012245f
C160 VTAIL.n92 B 0.012965f
C161 VTAIL.n93 B 0.028943f
C162 VTAIL.n94 B 0.028943f
C163 VTAIL.n95 B 0.012965f
C164 VTAIL.n96 B 0.012245f
C165 VTAIL.n97 B 0.022788f
C166 VTAIL.n98 B 0.022788f
C167 VTAIL.n99 B 0.012245f
C168 VTAIL.n100 B 0.012965f
C169 VTAIL.n101 B 0.028943f
C170 VTAIL.n102 B 0.062657f
C171 VTAIL.n103 B 0.012965f
C172 VTAIL.n104 B 0.012245f
C173 VTAIL.n105 B 0.051427f
C174 VTAIL.n106 B 0.03502f
C175 VTAIL.n107 B 0.095668f
C176 VTAIL.n108 B 0.03203f
C177 VTAIL.n109 B 0.022788f
C178 VTAIL.n110 B 0.012245f
C179 VTAIL.n111 B 0.028943f
C180 VTAIL.n112 B 0.012965f
C181 VTAIL.n113 B 0.022788f
C182 VTAIL.n114 B 0.012245f
C183 VTAIL.n115 B 0.028943f
C184 VTAIL.n116 B 0.012965f
C185 VTAIL.n117 B 0.022788f
C186 VTAIL.n118 B 0.012245f
C187 VTAIL.n119 B 0.028943f
C188 VTAIL.n120 B 0.012965f
C189 VTAIL.n121 B 0.022788f
C190 VTAIL.n122 B 0.012245f
C191 VTAIL.n123 B 0.028943f
C192 VTAIL.n124 B 0.012965f
C193 VTAIL.n125 B 0.022788f
C194 VTAIL.n126 B 0.012245f
C195 VTAIL.n127 B 0.028943f
C196 VTAIL.n128 B 0.012965f
C197 VTAIL.n129 B 0.022788f
C198 VTAIL.n130 B 0.012245f
C199 VTAIL.n131 B 0.028943f
C200 VTAIL.n132 B 0.012965f
C201 VTAIL.n133 B 0.022788f
C202 VTAIL.n134 B 0.012245f
C203 VTAIL.n135 B 0.028943f
C204 VTAIL.n136 B 0.012965f
C205 VTAIL.n137 B 0.022788f
C206 VTAIL.n138 B 0.012245f
C207 VTAIL.n139 B 0.028943f
C208 VTAIL.n140 B 0.012965f
C209 VTAIL.n141 B 0.171022f
C210 VTAIL.t3 B 0.04803f
C211 VTAIL.n142 B 0.021707f
C212 VTAIL.n143 B 0.017098f
C213 VTAIL.n144 B 0.012245f
C214 VTAIL.n145 B 1.89199f
C215 VTAIL.n146 B 0.022788f
C216 VTAIL.n147 B 0.012245f
C217 VTAIL.n148 B 0.012965f
C218 VTAIL.n149 B 0.028943f
C219 VTAIL.n150 B 0.028943f
C220 VTAIL.n151 B 0.012965f
C221 VTAIL.n152 B 0.012245f
C222 VTAIL.n153 B 0.022788f
C223 VTAIL.n154 B 0.022788f
C224 VTAIL.n155 B 0.012245f
C225 VTAIL.n156 B 0.012965f
C226 VTAIL.n157 B 0.028943f
C227 VTAIL.n158 B 0.028943f
C228 VTAIL.n159 B 0.012965f
C229 VTAIL.n160 B 0.012245f
C230 VTAIL.n161 B 0.022788f
C231 VTAIL.n162 B 0.022788f
C232 VTAIL.n163 B 0.012245f
C233 VTAIL.n164 B 0.012965f
C234 VTAIL.n165 B 0.028943f
C235 VTAIL.n166 B 0.028943f
C236 VTAIL.n167 B 0.012965f
C237 VTAIL.n168 B 0.012245f
C238 VTAIL.n169 B 0.022788f
C239 VTAIL.n170 B 0.022788f
C240 VTAIL.n171 B 0.012245f
C241 VTAIL.n172 B 0.012965f
C242 VTAIL.n173 B 0.028943f
C243 VTAIL.n174 B 0.028943f
C244 VTAIL.n175 B 0.012965f
C245 VTAIL.n176 B 0.012245f
C246 VTAIL.n177 B 0.022788f
C247 VTAIL.n178 B 0.022788f
C248 VTAIL.n179 B 0.012245f
C249 VTAIL.n180 B 0.012965f
C250 VTAIL.n181 B 0.028943f
C251 VTAIL.n182 B 0.028943f
C252 VTAIL.n183 B 0.028943f
C253 VTAIL.n184 B 0.012965f
C254 VTAIL.n185 B 0.012245f
C255 VTAIL.n186 B 0.022788f
C256 VTAIL.n187 B 0.022788f
C257 VTAIL.n188 B 0.012245f
C258 VTAIL.n189 B 0.012605f
C259 VTAIL.n190 B 0.012605f
C260 VTAIL.n191 B 0.028943f
C261 VTAIL.n192 B 0.028943f
C262 VTAIL.n193 B 0.012965f
C263 VTAIL.n194 B 0.012245f
C264 VTAIL.n195 B 0.022788f
C265 VTAIL.n196 B 0.022788f
C266 VTAIL.n197 B 0.012245f
C267 VTAIL.n198 B 0.012965f
C268 VTAIL.n199 B 0.028943f
C269 VTAIL.n200 B 0.028943f
C270 VTAIL.n201 B 0.012965f
C271 VTAIL.n202 B 0.012245f
C272 VTAIL.n203 B 0.022788f
C273 VTAIL.n204 B 0.022788f
C274 VTAIL.n205 B 0.012245f
C275 VTAIL.n206 B 0.012965f
C276 VTAIL.n207 B 0.028943f
C277 VTAIL.n208 B 0.062657f
C278 VTAIL.n209 B 0.012965f
C279 VTAIL.n210 B 0.012245f
C280 VTAIL.n211 B 0.051427f
C281 VTAIL.n212 B 0.03502f
C282 VTAIL.n213 B 0.095668f
C283 VTAIL.t5 B 0.340702f
C284 VTAIL.t4 B 0.340702f
C285 VTAIL.n214 B 3.03617f
C286 VTAIL.n215 B 0.317486f
C287 VTAIL.n216 B 0.03203f
C288 VTAIL.n217 B 0.022788f
C289 VTAIL.n218 B 0.012245f
C290 VTAIL.n219 B 0.028943f
C291 VTAIL.n220 B 0.012965f
C292 VTAIL.n221 B 0.022788f
C293 VTAIL.n222 B 0.012245f
C294 VTAIL.n223 B 0.028943f
C295 VTAIL.n224 B 0.012965f
C296 VTAIL.n225 B 0.022788f
C297 VTAIL.n226 B 0.012245f
C298 VTAIL.n227 B 0.028943f
C299 VTAIL.n228 B 0.012965f
C300 VTAIL.n229 B 0.022788f
C301 VTAIL.n230 B 0.012245f
C302 VTAIL.n231 B 0.028943f
C303 VTAIL.n232 B 0.012965f
C304 VTAIL.n233 B 0.022788f
C305 VTAIL.n234 B 0.012245f
C306 VTAIL.n235 B 0.028943f
C307 VTAIL.n236 B 0.012965f
C308 VTAIL.n237 B 0.022788f
C309 VTAIL.n238 B 0.012245f
C310 VTAIL.n239 B 0.028943f
C311 VTAIL.n240 B 0.012965f
C312 VTAIL.n241 B 0.022788f
C313 VTAIL.n242 B 0.012245f
C314 VTAIL.n243 B 0.028943f
C315 VTAIL.n244 B 0.012965f
C316 VTAIL.n245 B 0.022788f
C317 VTAIL.n246 B 0.012245f
C318 VTAIL.n247 B 0.028943f
C319 VTAIL.n248 B 0.012965f
C320 VTAIL.n249 B 0.171022f
C321 VTAIL.t7 B 0.04803f
C322 VTAIL.n250 B 0.021707f
C323 VTAIL.n251 B 0.017098f
C324 VTAIL.n252 B 0.012245f
C325 VTAIL.n253 B 1.89199f
C326 VTAIL.n254 B 0.022788f
C327 VTAIL.n255 B 0.012245f
C328 VTAIL.n256 B 0.012965f
C329 VTAIL.n257 B 0.028943f
C330 VTAIL.n258 B 0.028943f
C331 VTAIL.n259 B 0.012965f
C332 VTAIL.n260 B 0.012245f
C333 VTAIL.n261 B 0.022788f
C334 VTAIL.n262 B 0.022788f
C335 VTAIL.n263 B 0.012245f
C336 VTAIL.n264 B 0.012965f
C337 VTAIL.n265 B 0.028943f
C338 VTAIL.n266 B 0.028943f
C339 VTAIL.n267 B 0.012965f
C340 VTAIL.n268 B 0.012245f
C341 VTAIL.n269 B 0.022788f
C342 VTAIL.n270 B 0.022788f
C343 VTAIL.n271 B 0.012245f
C344 VTAIL.n272 B 0.012965f
C345 VTAIL.n273 B 0.028943f
C346 VTAIL.n274 B 0.028943f
C347 VTAIL.n275 B 0.012965f
C348 VTAIL.n276 B 0.012245f
C349 VTAIL.n277 B 0.022788f
C350 VTAIL.n278 B 0.022788f
C351 VTAIL.n279 B 0.012245f
C352 VTAIL.n280 B 0.012965f
C353 VTAIL.n281 B 0.028943f
C354 VTAIL.n282 B 0.028943f
C355 VTAIL.n283 B 0.012965f
C356 VTAIL.n284 B 0.012245f
C357 VTAIL.n285 B 0.022788f
C358 VTAIL.n286 B 0.022788f
C359 VTAIL.n287 B 0.012245f
C360 VTAIL.n288 B 0.012965f
C361 VTAIL.n289 B 0.028943f
C362 VTAIL.n290 B 0.028943f
C363 VTAIL.n291 B 0.028943f
C364 VTAIL.n292 B 0.012965f
C365 VTAIL.n293 B 0.012245f
C366 VTAIL.n294 B 0.022788f
C367 VTAIL.n295 B 0.022788f
C368 VTAIL.n296 B 0.012245f
C369 VTAIL.n297 B 0.012605f
C370 VTAIL.n298 B 0.012605f
C371 VTAIL.n299 B 0.028943f
C372 VTAIL.n300 B 0.028943f
C373 VTAIL.n301 B 0.012965f
C374 VTAIL.n302 B 0.012245f
C375 VTAIL.n303 B 0.022788f
C376 VTAIL.n304 B 0.022788f
C377 VTAIL.n305 B 0.012245f
C378 VTAIL.n306 B 0.012965f
C379 VTAIL.n307 B 0.028943f
C380 VTAIL.n308 B 0.028943f
C381 VTAIL.n309 B 0.012965f
C382 VTAIL.n310 B 0.012245f
C383 VTAIL.n311 B 0.022788f
C384 VTAIL.n312 B 0.022788f
C385 VTAIL.n313 B 0.012245f
C386 VTAIL.n314 B 0.012965f
C387 VTAIL.n315 B 0.028943f
C388 VTAIL.n316 B 0.062657f
C389 VTAIL.n317 B 0.012965f
C390 VTAIL.n318 B 0.012245f
C391 VTAIL.n319 B 0.051427f
C392 VTAIL.n320 B 0.03502f
C393 VTAIL.n321 B 1.61074f
C394 VTAIL.n322 B 0.03203f
C395 VTAIL.n323 B 0.022788f
C396 VTAIL.n324 B 0.012245f
C397 VTAIL.n325 B 0.028943f
C398 VTAIL.n326 B 0.012965f
C399 VTAIL.n327 B 0.022788f
C400 VTAIL.n328 B 0.012245f
C401 VTAIL.n329 B 0.028943f
C402 VTAIL.n330 B 0.012965f
C403 VTAIL.n331 B 0.022788f
C404 VTAIL.n332 B 0.012245f
C405 VTAIL.n333 B 0.028943f
C406 VTAIL.n334 B 0.012965f
C407 VTAIL.n335 B 0.022788f
C408 VTAIL.n336 B 0.012245f
C409 VTAIL.n337 B 0.028943f
C410 VTAIL.n338 B 0.028943f
C411 VTAIL.n339 B 0.012965f
C412 VTAIL.n340 B 0.022788f
C413 VTAIL.n341 B 0.012245f
C414 VTAIL.n342 B 0.028943f
C415 VTAIL.n343 B 0.012965f
C416 VTAIL.n344 B 0.022788f
C417 VTAIL.n345 B 0.012245f
C418 VTAIL.n346 B 0.028943f
C419 VTAIL.n347 B 0.012965f
C420 VTAIL.n348 B 0.022788f
C421 VTAIL.n349 B 0.012245f
C422 VTAIL.n350 B 0.028943f
C423 VTAIL.n351 B 0.012965f
C424 VTAIL.n352 B 0.022788f
C425 VTAIL.n353 B 0.012245f
C426 VTAIL.n354 B 0.028943f
C427 VTAIL.n355 B 0.012965f
C428 VTAIL.n356 B 0.171022f
C429 VTAIL.t14 B 0.04803f
C430 VTAIL.n357 B 0.021707f
C431 VTAIL.n358 B 0.017098f
C432 VTAIL.n359 B 0.012245f
C433 VTAIL.n360 B 1.89199f
C434 VTAIL.n361 B 0.022788f
C435 VTAIL.n362 B 0.012245f
C436 VTAIL.n363 B 0.012965f
C437 VTAIL.n364 B 0.028943f
C438 VTAIL.n365 B 0.028943f
C439 VTAIL.n366 B 0.012965f
C440 VTAIL.n367 B 0.012245f
C441 VTAIL.n368 B 0.022788f
C442 VTAIL.n369 B 0.022788f
C443 VTAIL.n370 B 0.012245f
C444 VTAIL.n371 B 0.012965f
C445 VTAIL.n372 B 0.028943f
C446 VTAIL.n373 B 0.028943f
C447 VTAIL.n374 B 0.012965f
C448 VTAIL.n375 B 0.012245f
C449 VTAIL.n376 B 0.022788f
C450 VTAIL.n377 B 0.022788f
C451 VTAIL.n378 B 0.012245f
C452 VTAIL.n379 B 0.012965f
C453 VTAIL.n380 B 0.028943f
C454 VTAIL.n381 B 0.028943f
C455 VTAIL.n382 B 0.012965f
C456 VTAIL.n383 B 0.012245f
C457 VTAIL.n384 B 0.022788f
C458 VTAIL.n385 B 0.022788f
C459 VTAIL.n386 B 0.012245f
C460 VTAIL.n387 B 0.012965f
C461 VTAIL.n388 B 0.028943f
C462 VTAIL.n389 B 0.028943f
C463 VTAIL.n390 B 0.012965f
C464 VTAIL.n391 B 0.012245f
C465 VTAIL.n392 B 0.022788f
C466 VTAIL.n393 B 0.022788f
C467 VTAIL.n394 B 0.012245f
C468 VTAIL.n395 B 0.012965f
C469 VTAIL.n396 B 0.028943f
C470 VTAIL.n397 B 0.028943f
C471 VTAIL.n398 B 0.012965f
C472 VTAIL.n399 B 0.012245f
C473 VTAIL.n400 B 0.022788f
C474 VTAIL.n401 B 0.022788f
C475 VTAIL.n402 B 0.012245f
C476 VTAIL.n403 B 0.012605f
C477 VTAIL.n404 B 0.012605f
C478 VTAIL.n405 B 0.028943f
C479 VTAIL.n406 B 0.028943f
C480 VTAIL.n407 B 0.012965f
C481 VTAIL.n408 B 0.012245f
C482 VTAIL.n409 B 0.022788f
C483 VTAIL.n410 B 0.022788f
C484 VTAIL.n411 B 0.012245f
C485 VTAIL.n412 B 0.012965f
C486 VTAIL.n413 B 0.028943f
C487 VTAIL.n414 B 0.028943f
C488 VTAIL.n415 B 0.012965f
C489 VTAIL.n416 B 0.012245f
C490 VTAIL.n417 B 0.022788f
C491 VTAIL.n418 B 0.022788f
C492 VTAIL.n419 B 0.012245f
C493 VTAIL.n420 B 0.012965f
C494 VTAIL.n421 B 0.028943f
C495 VTAIL.n422 B 0.062657f
C496 VTAIL.n423 B 0.012965f
C497 VTAIL.n424 B 0.012245f
C498 VTAIL.n425 B 0.051427f
C499 VTAIL.n426 B 0.03502f
C500 VTAIL.n427 B 1.61074f
C501 VTAIL.t12 B 0.340702f
C502 VTAIL.t13 B 0.340702f
C503 VTAIL.n428 B 3.03617f
C504 VTAIL.n429 B 0.317484f
C505 VTAIL.n430 B 0.03203f
C506 VTAIL.n431 B 0.022788f
C507 VTAIL.n432 B 0.012245f
C508 VTAIL.n433 B 0.028943f
C509 VTAIL.n434 B 0.012965f
C510 VTAIL.n435 B 0.022788f
C511 VTAIL.n436 B 0.012245f
C512 VTAIL.n437 B 0.028943f
C513 VTAIL.n438 B 0.012965f
C514 VTAIL.n439 B 0.022788f
C515 VTAIL.n440 B 0.012245f
C516 VTAIL.n441 B 0.028943f
C517 VTAIL.n442 B 0.012965f
C518 VTAIL.n443 B 0.022788f
C519 VTAIL.n444 B 0.012245f
C520 VTAIL.n445 B 0.028943f
C521 VTAIL.n446 B 0.028943f
C522 VTAIL.n447 B 0.012965f
C523 VTAIL.n448 B 0.022788f
C524 VTAIL.n449 B 0.012245f
C525 VTAIL.n450 B 0.028943f
C526 VTAIL.n451 B 0.012965f
C527 VTAIL.n452 B 0.022788f
C528 VTAIL.n453 B 0.012245f
C529 VTAIL.n454 B 0.028943f
C530 VTAIL.n455 B 0.012965f
C531 VTAIL.n456 B 0.022788f
C532 VTAIL.n457 B 0.012245f
C533 VTAIL.n458 B 0.028943f
C534 VTAIL.n459 B 0.012965f
C535 VTAIL.n460 B 0.022788f
C536 VTAIL.n461 B 0.012245f
C537 VTAIL.n462 B 0.028943f
C538 VTAIL.n463 B 0.012965f
C539 VTAIL.n464 B 0.171022f
C540 VTAIL.t8 B 0.04803f
C541 VTAIL.n465 B 0.021707f
C542 VTAIL.n466 B 0.017098f
C543 VTAIL.n467 B 0.012245f
C544 VTAIL.n468 B 1.89199f
C545 VTAIL.n469 B 0.022788f
C546 VTAIL.n470 B 0.012245f
C547 VTAIL.n471 B 0.012965f
C548 VTAIL.n472 B 0.028943f
C549 VTAIL.n473 B 0.028943f
C550 VTAIL.n474 B 0.012965f
C551 VTAIL.n475 B 0.012245f
C552 VTAIL.n476 B 0.022788f
C553 VTAIL.n477 B 0.022788f
C554 VTAIL.n478 B 0.012245f
C555 VTAIL.n479 B 0.012965f
C556 VTAIL.n480 B 0.028943f
C557 VTAIL.n481 B 0.028943f
C558 VTAIL.n482 B 0.012965f
C559 VTAIL.n483 B 0.012245f
C560 VTAIL.n484 B 0.022788f
C561 VTAIL.n485 B 0.022788f
C562 VTAIL.n486 B 0.012245f
C563 VTAIL.n487 B 0.012965f
C564 VTAIL.n488 B 0.028943f
C565 VTAIL.n489 B 0.028943f
C566 VTAIL.n490 B 0.012965f
C567 VTAIL.n491 B 0.012245f
C568 VTAIL.n492 B 0.022788f
C569 VTAIL.n493 B 0.022788f
C570 VTAIL.n494 B 0.012245f
C571 VTAIL.n495 B 0.012965f
C572 VTAIL.n496 B 0.028943f
C573 VTAIL.n497 B 0.028943f
C574 VTAIL.n498 B 0.012965f
C575 VTAIL.n499 B 0.012245f
C576 VTAIL.n500 B 0.022788f
C577 VTAIL.n501 B 0.022788f
C578 VTAIL.n502 B 0.012245f
C579 VTAIL.n503 B 0.012965f
C580 VTAIL.n504 B 0.028943f
C581 VTAIL.n505 B 0.028943f
C582 VTAIL.n506 B 0.012965f
C583 VTAIL.n507 B 0.012245f
C584 VTAIL.n508 B 0.022788f
C585 VTAIL.n509 B 0.022788f
C586 VTAIL.n510 B 0.012245f
C587 VTAIL.n511 B 0.012605f
C588 VTAIL.n512 B 0.012605f
C589 VTAIL.n513 B 0.028943f
C590 VTAIL.n514 B 0.028943f
C591 VTAIL.n515 B 0.012965f
C592 VTAIL.n516 B 0.012245f
C593 VTAIL.n517 B 0.022788f
C594 VTAIL.n518 B 0.022788f
C595 VTAIL.n519 B 0.012245f
C596 VTAIL.n520 B 0.012965f
C597 VTAIL.n521 B 0.028943f
C598 VTAIL.n522 B 0.028943f
C599 VTAIL.n523 B 0.012965f
C600 VTAIL.n524 B 0.012245f
C601 VTAIL.n525 B 0.022788f
C602 VTAIL.n526 B 0.022788f
C603 VTAIL.n527 B 0.012245f
C604 VTAIL.n528 B 0.012965f
C605 VTAIL.n529 B 0.028943f
C606 VTAIL.n530 B 0.062657f
C607 VTAIL.n531 B 0.012965f
C608 VTAIL.n532 B 0.012245f
C609 VTAIL.n533 B 0.051427f
C610 VTAIL.n534 B 0.03502f
C611 VTAIL.n535 B 0.095668f
C612 VTAIL.n536 B 0.03203f
C613 VTAIL.n537 B 0.022788f
C614 VTAIL.n538 B 0.012245f
C615 VTAIL.n539 B 0.028943f
C616 VTAIL.n540 B 0.012965f
C617 VTAIL.n541 B 0.022788f
C618 VTAIL.n542 B 0.012245f
C619 VTAIL.n543 B 0.028943f
C620 VTAIL.n544 B 0.012965f
C621 VTAIL.n545 B 0.022788f
C622 VTAIL.n546 B 0.012245f
C623 VTAIL.n547 B 0.028943f
C624 VTAIL.n548 B 0.012965f
C625 VTAIL.n549 B 0.022788f
C626 VTAIL.n550 B 0.012245f
C627 VTAIL.n551 B 0.028943f
C628 VTAIL.n552 B 0.028943f
C629 VTAIL.n553 B 0.012965f
C630 VTAIL.n554 B 0.022788f
C631 VTAIL.n555 B 0.012245f
C632 VTAIL.n556 B 0.028943f
C633 VTAIL.n557 B 0.012965f
C634 VTAIL.n558 B 0.022788f
C635 VTAIL.n559 B 0.012245f
C636 VTAIL.n560 B 0.028943f
C637 VTAIL.n561 B 0.012965f
C638 VTAIL.n562 B 0.022788f
C639 VTAIL.n563 B 0.012245f
C640 VTAIL.n564 B 0.028943f
C641 VTAIL.n565 B 0.012965f
C642 VTAIL.n566 B 0.022788f
C643 VTAIL.n567 B 0.012245f
C644 VTAIL.n568 B 0.028943f
C645 VTAIL.n569 B 0.012965f
C646 VTAIL.n570 B 0.171022f
C647 VTAIL.t0 B 0.04803f
C648 VTAIL.n571 B 0.021707f
C649 VTAIL.n572 B 0.017098f
C650 VTAIL.n573 B 0.012245f
C651 VTAIL.n574 B 1.89199f
C652 VTAIL.n575 B 0.022788f
C653 VTAIL.n576 B 0.012245f
C654 VTAIL.n577 B 0.012965f
C655 VTAIL.n578 B 0.028943f
C656 VTAIL.n579 B 0.028943f
C657 VTAIL.n580 B 0.012965f
C658 VTAIL.n581 B 0.012245f
C659 VTAIL.n582 B 0.022788f
C660 VTAIL.n583 B 0.022788f
C661 VTAIL.n584 B 0.012245f
C662 VTAIL.n585 B 0.012965f
C663 VTAIL.n586 B 0.028943f
C664 VTAIL.n587 B 0.028943f
C665 VTAIL.n588 B 0.012965f
C666 VTAIL.n589 B 0.012245f
C667 VTAIL.n590 B 0.022788f
C668 VTAIL.n591 B 0.022788f
C669 VTAIL.n592 B 0.012245f
C670 VTAIL.n593 B 0.012965f
C671 VTAIL.n594 B 0.028943f
C672 VTAIL.n595 B 0.028943f
C673 VTAIL.n596 B 0.012965f
C674 VTAIL.n597 B 0.012245f
C675 VTAIL.n598 B 0.022788f
C676 VTAIL.n599 B 0.022788f
C677 VTAIL.n600 B 0.012245f
C678 VTAIL.n601 B 0.012965f
C679 VTAIL.n602 B 0.028943f
C680 VTAIL.n603 B 0.028943f
C681 VTAIL.n604 B 0.012965f
C682 VTAIL.n605 B 0.012245f
C683 VTAIL.n606 B 0.022788f
C684 VTAIL.n607 B 0.022788f
C685 VTAIL.n608 B 0.012245f
C686 VTAIL.n609 B 0.012965f
C687 VTAIL.n610 B 0.028943f
C688 VTAIL.n611 B 0.028943f
C689 VTAIL.n612 B 0.012965f
C690 VTAIL.n613 B 0.012245f
C691 VTAIL.n614 B 0.022788f
C692 VTAIL.n615 B 0.022788f
C693 VTAIL.n616 B 0.012245f
C694 VTAIL.n617 B 0.012605f
C695 VTAIL.n618 B 0.012605f
C696 VTAIL.n619 B 0.028943f
C697 VTAIL.n620 B 0.028943f
C698 VTAIL.n621 B 0.012965f
C699 VTAIL.n622 B 0.012245f
C700 VTAIL.n623 B 0.022788f
C701 VTAIL.n624 B 0.022788f
C702 VTAIL.n625 B 0.012245f
C703 VTAIL.n626 B 0.012965f
C704 VTAIL.n627 B 0.028943f
C705 VTAIL.n628 B 0.028943f
C706 VTAIL.n629 B 0.012965f
C707 VTAIL.n630 B 0.012245f
C708 VTAIL.n631 B 0.022788f
C709 VTAIL.n632 B 0.022788f
C710 VTAIL.n633 B 0.012245f
C711 VTAIL.n634 B 0.012965f
C712 VTAIL.n635 B 0.028943f
C713 VTAIL.n636 B 0.062657f
C714 VTAIL.n637 B 0.012965f
C715 VTAIL.n638 B 0.012245f
C716 VTAIL.n639 B 0.051427f
C717 VTAIL.n640 B 0.03502f
C718 VTAIL.n641 B 0.095668f
C719 VTAIL.t1 B 0.340702f
C720 VTAIL.t6 B 0.340702f
C721 VTAIL.n642 B 3.03617f
C722 VTAIL.n643 B 0.317484f
C723 VTAIL.n644 B 0.03203f
C724 VTAIL.n645 B 0.022788f
C725 VTAIL.n646 B 0.012245f
C726 VTAIL.n647 B 0.028943f
C727 VTAIL.n648 B 0.012965f
C728 VTAIL.n649 B 0.022788f
C729 VTAIL.n650 B 0.012245f
C730 VTAIL.n651 B 0.028943f
C731 VTAIL.n652 B 0.012965f
C732 VTAIL.n653 B 0.022788f
C733 VTAIL.n654 B 0.012245f
C734 VTAIL.n655 B 0.028943f
C735 VTAIL.n656 B 0.012965f
C736 VTAIL.n657 B 0.022788f
C737 VTAIL.n658 B 0.012245f
C738 VTAIL.n659 B 0.028943f
C739 VTAIL.n660 B 0.028943f
C740 VTAIL.n661 B 0.012965f
C741 VTAIL.n662 B 0.022788f
C742 VTAIL.n663 B 0.012245f
C743 VTAIL.n664 B 0.028943f
C744 VTAIL.n665 B 0.012965f
C745 VTAIL.n666 B 0.022788f
C746 VTAIL.n667 B 0.012245f
C747 VTAIL.n668 B 0.028943f
C748 VTAIL.n669 B 0.012965f
C749 VTAIL.n670 B 0.022788f
C750 VTAIL.n671 B 0.012245f
C751 VTAIL.n672 B 0.028943f
C752 VTAIL.n673 B 0.012965f
C753 VTAIL.n674 B 0.022788f
C754 VTAIL.n675 B 0.012245f
C755 VTAIL.n676 B 0.028943f
C756 VTAIL.n677 B 0.012965f
C757 VTAIL.n678 B 0.171022f
C758 VTAIL.t2 B 0.04803f
C759 VTAIL.n679 B 0.021707f
C760 VTAIL.n680 B 0.017098f
C761 VTAIL.n681 B 0.012245f
C762 VTAIL.n682 B 1.89199f
C763 VTAIL.n683 B 0.022788f
C764 VTAIL.n684 B 0.012245f
C765 VTAIL.n685 B 0.012965f
C766 VTAIL.n686 B 0.028943f
C767 VTAIL.n687 B 0.028943f
C768 VTAIL.n688 B 0.012965f
C769 VTAIL.n689 B 0.012245f
C770 VTAIL.n690 B 0.022788f
C771 VTAIL.n691 B 0.022788f
C772 VTAIL.n692 B 0.012245f
C773 VTAIL.n693 B 0.012965f
C774 VTAIL.n694 B 0.028943f
C775 VTAIL.n695 B 0.028943f
C776 VTAIL.n696 B 0.012965f
C777 VTAIL.n697 B 0.012245f
C778 VTAIL.n698 B 0.022788f
C779 VTAIL.n699 B 0.022788f
C780 VTAIL.n700 B 0.012245f
C781 VTAIL.n701 B 0.012965f
C782 VTAIL.n702 B 0.028943f
C783 VTAIL.n703 B 0.028943f
C784 VTAIL.n704 B 0.012965f
C785 VTAIL.n705 B 0.012245f
C786 VTAIL.n706 B 0.022788f
C787 VTAIL.n707 B 0.022788f
C788 VTAIL.n708 B 0.012245f
C789 VTAIL.n709 B 0.012965f
C790 VTAIL.n710 B 0.028943f
C791 VTAIL.n711 B 0.028943f
C792 VTAIL.n712 B 0.012965f
C793 VTAIL.n713 B 0.012245f
C794 VTAIL.n714 B 0.022788f
C795 VTAIL.n715 B 0.022788f
C796 VTAIL.n716 B 0.012245f
C797 VTAIL.n717 B 0.012965f
C798 VTAIL.n718 B 0.028943f
C799 VTAIL.n719 B 0.028943f
C800 VTAIL.n720 B 0.012965f
C801 VTAIL.n721 B 0.012245f
C802 VTAIL.n722 B 0.022788f
C803 VTAIL.n723 B 0.022788f
C804 VTAIL.n724 B 0.012245f
C805 VTAIL.n725 B 0.012605f
C806 VTAIL.n726 B 0.012605f
C807 VTAIL.n727 B 0.028943f
C808 VTAIL.n728 B 0.028943f
C809 VTAIL.n729 B 0.012965f
C810 VTAIL.n730 B 0.012245f
C811 VTAIL.n731 B 0.022788f
C812 VTAIL.n732 B 0.022788f
C813 VTAIL.n733 B 0.012245f
C814 VTAIL.n734 B 0.012965f
C815 VTAIL.n735 B 0.028943f
C816 VTAIL.n736 B 0.028943f
C817 VTAIL.n737 B 0.012965f
C818 VTAIL.n738 B 0.012245f
C819 VTAIL.n739 B 0.022788f
C820 VTAIL.n740 B 0.022788f
C821 VTAIL.n741 B 0.012245f
C822 VTAIL.n742 B 0.012965f
C823 VTAIL.n743 B 0.028943f
C824 VTAIL.n744 B 0.062657f
C825 VTAIL.n745 B 0.012965f
C826 VTAIL.n746 B 0.012245f
C827 VTAIL.n747 B 0.051427f
C828 VTAIL.n748 B 0.03502f
C829 VTAIL.n749 B 1.61074f
C830 VTAIL.n750 B 0.03203f
C831 VTAIL.n751 B 0.022788f
C832 VTAIL.n752 B 0.012245f
C833 VTAIL.n753 B 0.028943f
C834 VTAIL.n754 B 0.012965f
C835 VTAIL.n755 B 0.022788f
C836 VTAIL.n756 B 0.012245f
C837 VTAIL.n757 B 0.028943f
C838 VTAIL.n758 B 0.012965f
C839 VTAIL.n759 B 0.022788f
C840 VTAIL.n760 B 0.012245f
C841 VTAIL.n761 B 0.028943f
C842 VTAIL.n762 B 0.012965f
C843 VTAIL.n763 B 0.022788f
C844 VTAIL.n764 B 0.012245f
C845 VTAIL.n765 B 0.028943f
C846 VTAIL.n766 B 0.012965f
C847 VTAIL.n767 B 0.022788f
C848 VTAIL.n768 B 0.012245f
C849 VTAIL.n769 B 0.028943f
C850 VTAIL.n770 B 0.012965f
C851 VTAIL.n771 B 0.022788f
C852 VTAIL.n772 B 0.012245f
C853 VTAIL.n773 B 0.028943f
C854 VTAIL.n774 B 0.012965f
C855 VTAIL.n775 B 0.022788f
C856 VTAIL.n776 B 0.012245f
C857 VTAIL.n777 B 0.028943f
C858 VTAIL.n778 B 0.012965f
C859 VTAIL.n779 B 0.022788f
C860 VTAIL.n780 B 0.012245f
C861 VTAIL.n781 B 0.028943f
C862 VTAIL.n782 B 0.012965f
C863 VTAIL.n783 B 0.171022f
C864 VTAIL.t9 B 0.04803f
C865 VTAIL.n784 B 0.021707f
C866 VTAIL.n785 B 0.017098f
C867 VTAIL.n786 B 0.012245f
C868 VTAIL.n787 B 1.89199f
C869 VTAIL.n788 B 0.022788f
C870 VTAIL.n789 B 0.012245f
C871 VTAIL.n790 B 0.012965f
C872 VTAIL.n791 B 0.028943f
C873 VTAIL.n792 B 0.028943f
C874 VTAIL.n793 B 0.012965f
C875 VTAIL.n794 B 0.012245f
C876 VTAIL.n795 B 0.022788f
C877 VTAIL.n796 B 0.022788f
C878 VTAIL.n797 B 0.012245f
C879 VTAIL.n798 B 0.012965f
C880 VTAIL.n799 B 0.028943f
C881 VTAIL.n800 B 0.028943f
C882 VTAIL.n801 B 0.012965f
C883 VTAIL.n802 B 0.012245f
C884 VTAIL.n803 B 0.022788f
C885 VTAIL.n804 B 0.022788f
C886 VTAIL.n805 B 0.012245f
C887 VTAIL.n806 B 0.012965f
C888 VTAIL.n807 B 0.028943f
C889 VTAIL.n808 B 0.028943f
C890 VTAIL.n809 B 0.012965f
C891 VTAIL.n810 B 0.012245f
C892 VTAIL.n811 B 0.022788f
C893 VTAIL.n812 B 0.022788f
C894 VTAIL.n813 B 0.012245f
C895 VTAIL.n814 B 0.012965f
C896 VTAIL.n815 B 0.028943f
C897 VTAIL.n816 B 0.028943f
C898 VTAIL.n817 B 0.012965f
C899 VTAIL.n818 B 0.012245f
C900 VTAIL.n819 B 0.022788f
C901 VTAIL.n820 B 0.022788f
C902 VTAIL.n821 B 0.012245f
C903 VTAIL.n822 B 0.012965f
C904 VTAIL.n823 B 0.028943f
C905 VTAIL.n824 B 0.028943f
C906 VTAIL.n825 B 0.028943f
C907 VTAIL.n826 B 0.012965f
C908 VTAIL.n827 B 0.012245f
C909 VTAIL.n828 B 0.022788f
C910 VTAIL.n829 B 0.022788f
C911 VTAIL.n830 B 0.012245f
C912 VTAIL.n831 B 0.012605f
C913 VTAIL.n832 B 0.012605f
C914 VTAIL.n833 B 0.028943f
C915 VTAIL.n834 B 0.028943f
C916 VTAIL.n835 B 0.012965f
C917 VTAIL.n836 B 0.012245f
C918 VTAIL.n837 B 0.022788f
C919 VTAIL.n838 B 0.022788f
C920 VTAIL.n839 B 0.012245f
C921 VTAIL.n840 B 0.012965f
C922 VTAIL.n841 B 0.028943f
C923 VTAIL.n842 B 0.028943f
C924 VTAIL.n843 B 0.012965f
C925 VTAIL.n844 B 0.012245f
C926 VTAIL.n845 B 0.022788f
C927 VTAIL.n846 B 0.022788f
C928 VTAIL.n847 B 0.012245f
C929 VTAIL.n848 B 0.012965f
C930 VTAIL.n849 B 0.028943f
C931 VTAIL.n850 B 0.062657f
C932 VTAIL.n851 B 0.012965f
C933 VTAIL.n852 B 0.012245f
C934 VTAIL.n853 B 0.051427f
C935 VTAIL.n854 B 0.03502f
C936 VTAIL.n855 B 1.60647f
C937 VN.n0 B 0.173306f
C938 VN.t6 B 0.992057f
C939 VN.n1 B 0.372502f
C940 VN.t3 B 0.984879f
C941 VN.n2 B 0.38462f
C942 VN.t2 B 0.984879f
C943 VN.n3 B 0.38462f
C944 VN.t4 B 0.987978f
C945 VN.n4 B 0.376193f
C946 VN.n5 B 0.041858f
C947 VN.n6 B 0.173306f
C948 VN.t7 B 0.987978f
C949 VN.t1 B 0.984879f
C950 VN.t5 B 0.992057f
C951 VN.n7 B 0.372502f
C952 VN.n8 B 0.38462f
C953 VN.t0 B 0.984879f
C954 VN.n9 B 0.38462f
C955 VN.n10 B 0.376193f
C956 VN.n11 B 2.58507f
.ends

