* NGSPICE file created from diff_pair_sample_1327.ext - technology: sky130A

.subckt diff_pair_sample_1327 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=0 ps=0 w=12.46 l=3.65
X1 VTAIL.t15 VP.t0 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X2 VDD2.t7 VN.t0 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=4.8594 ps=25.7 w=12.46 l=3.65
X3 VTAIL.t2 VN.t1 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=2.0559 ps=12.79 w=12.46 l=3.65
X4 VDD2.t5 VN.t2 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X5 VTAIL.t14 VP.t1 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=0 ps=0 w=12.46 l=3.65
X7 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=0 ps=0 w=12.46 l=3.65
X8 VTAIL.t7 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=2.0559 ps=12.79 w=12.46 l=3.65
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=0 ps=0 w=12.46 l=3.65
X10 VDD1.t2 VP.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X11 VTAIL.t5 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X12 VDD2.t2 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X13 VDD1.t7 VP.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=4.8594 ps=25.7 w=12.46 l=3.65
X14 VDD1.t3 VP.t4 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X15 VTAIL.t4 VN.t6 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=2.0559 ps=12.79 w=12.46 l=3.65
X16 VTAIL.t10 VP.t5 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=2.0559 ps=12.79 w=12.46 l=3.65
X17 VDD2.t0 VN.t7 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=4.8594 ps=25.7 w=12.46 l=3.65
X18 VDD1.t4 VP.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0559 pd=12.79 as=4.8594 ps=25.7 w=12.46 l=3.65
X19 VTAIL.t8 VP.t7 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=4.8594 pd=25.7 as=2.0559 ps=12.79 w=12.46 l=3.65
R0 B.n831 B.n830 585
R1 B.n831 B.n121 585
R2 B.n834 B.n833 585
R3 B.n835 B.n173 585
R4 B.n837 B.n836 585
R5 B.n839 B.n172 585
R6 B.n842 B.n841 585
R7 B.n843 B.n171 585
R8 B.n845 B.n844 585
R9 B.n847 B.n170 585
R10 B.n850 B.n849 585
R11 B.n851 B.n169 585
R12 B.n853 B.n852 585
R13 B.n855 B.n168 585
R14 B.n858 B.n857 585
R15 B.n859 B.n167 585
R16 B.n861 B.n860 585
R17 B.n863 B.n166 585
R18 B.n866 B.n865 585
R19 B.n867 B.n165 585
R20 B.n869 B.n868 585
R21 B.n871 B.n164 585
R22 B.n874 B.n873 585
R23 B.n875 B.n163 585
R24 B.n877 B.n876 585
R25 B.n879 B.n162 585
R26 B.n882 B.n881 585
R27 B.n883 B.n161 585
R28 B.n885 B.n884 585
R29 B.n887 B.n160 585
R30 B.n890 B.n889 585
R31 B.n891 B.n159 585
R32 B.n893 B.n892 585
R33 B.n895 B.n158 585
R34 B.n898 B.n897 585
R35 B.n899 B.n157 585
R36 B.n901 B.n900 585
R37 B.n903 B.n156 585
R38 B.n906 B.n905 585
R39 B.n907 B.n155 585
R40 B.n909 B.n908 585
R41 B.n911 B.n154 585
R42 B.n914 B.n913 585
R43 B.n915 B.n151 585
R44 B.n918 B.n917 585
R45 B.n920 B.n150 585
R46 B.n923 B.n922 585
R47 B.n924 B.n149 585
R48 B.n926 B.n925 585
R49 B.n928 B.n148 585
R50 B.n931 B.n930 585
R51 B.n932 B.n144 585
R52 B.n934 B.n933 585
R53 B.n936 B.n143 585
R54 B.n939 B.n938 585
R55 B.n940 B.n142 585
R56 B.n942 B.n941 585
R57 B.n944 B.n141 585
R58 B.n947 B.n946 585
R59 B.n948 B.n140 585
R60 B.n950 B.n949 585
R61 B.n952 B.n139 585
R62 B.n955 B.n954 585
R63 B.n956 B.n138 585
R64 B.n958 B.n957 585
R65 B.n960 B.n137 585
R66 B.n963 B.n962 585
R67 B.n964 B.n136 585
R68 B.n966 B.n965 585
R69 B.n968 B.n135 585
R70 B.n971 B.n970 585
R71 B.n972 B.n134 585
R72 B.n974 B.n973 585
R73 B.n976 B.n133 585
R74 B.n979 B.n978 585
R75 B.n980 B.n132 585
R76 B.n982 B.n981 585
R77 B.n984 B.n131 585
R78 B.n987 B.n986 585
R79 B.n988 B.n130 585
R80 B.n990 B.n989 585
R81 B.n992 B.n129 585
R82 B.n995 B.n994 585
R83 B.n996 B.n128 585
R84 B.n998 B.n997 585
R85 B.n1000 B.n127 585
R86 B.n1003 B.n1002 585
R87 B.n1004 B.n126 585
R88 B.n1006 B.n1005 585
R89 B.n1008 B.n125 585
R90 B.n1011 B.n1010 585
R91 B.n1012 B.n124 585
R92 B.n1014 B.n1013 585
R93 B.n1016 B.n123 585
R94 B.n1019 B.n1018 585
R95 B.n1020 B.n122 585
R96 B.n829 B.n120 585
R97 B.n1023 B.n120 585
R98 B.n828 B.n119 585
R99 B.n1024 B.n119 585
R100 B.n827 B.n118 585
R101 B.n1025 B.n118 585
R102 B.n826 B.n825 585
R103 B.n825 B.n114 585
R104 B.n824 B.n113 585
R105 B.n1031 B.n113 585
R106 B.n823 B.n112 585
R107 B.n1032 B.n112 585
R108 B.n822 B.n111 585
R109 B.n1033 B.n111 585
R110 B.n821 B.n820 585
R111 B.n820 B.n107 585
R112 B.n819 B.n106 585
R113 B.n1039 B.n106 585
R114 B.n818 B.n105 585
R115 B.n1040 B.n105 585
R116 B.n817 B.n104 585
R117 B.n1041 B.n104 585
R118 B.n816 B.n815 585
R119 B.n815 B.n100 585
R120 B.n814 B.n99 585
R121 B.n1047 B.n99 585
R122 B.n813 B.n98 585
R123 B.n1048 B.n98 585
R124 B.n812 B.n97 585
R125 B.n1049 B.n97 585
R126 B.n811 B.n810 585
R127 B.n810 B.n93 585
R128 B.n809 B.n92 585
R129 B.n1055 B.n92 585
R130 B.n808 B.n91 585
R131 B.n1056 B.n91 585
R132 B.n807 B.n90 585
R133 B.n1057 B.n90 585
R134 B.n806 B.n805 585
R135 B.n805 B.n86 585
R136 B.n804 B.n85 585
R137 B.n1063 B.n85 585
R138 B.n803 B.n84 585
R139 B.n1064 B.n84 585
R140 B.n802 B.n83 585
R141 B.n1065 B.n83 585
R142 B.n801 B.n800 585
R143 B.n800 B.n82 585
R144 B.n799 B.n78 585
R145 B.n1071 B.n78 585
R146 B.n798 B.n77 585
R147 B.n1072 B.n77 585
R148 B.n797 B.n76 585
R149 B.n1073 B.n76 585
R150 B.n796 B.n795 585
R151 B.n795 B.n72 585
R152 B.n794 B.n71 585
R153 B.n1079 B.n71 585
R154 B.n793 B.n70 585
R155 B.n1080 B.n70 585
R156 B.n792 B.n69 585
R157 B.n1081 B.n69 585
R158 B.n791 B.n790 585
R159 B.n790 B.n65 585
R160 B.n789 B.n64 585
R161 B.n1087 B.n64 585
R162 B.n788 B.n63 585
R163 B.n1088 B.n63 585
R164 B.n787 B.n62 585
R165 B.n1089 B.n62 585
R166 B.n786 B.n785 585
R167 B.n785 B.n61 585
R168 B.n784 B.n57 585
R169 B.n1095 B.n57 585
R170 B.n783 B.n56 585
R171 B.n1096 B.n56 585
R172 B.n782 B.n55 585
R173 B.n1097 B.n55 585
R174 B.n781 B.n780 585
R175 B.n780 B.n51 585
R176 B.n779 B.n50 585
R177 B.n1103 B.n50 585
R178 B.n778 B.n49 585
R179 B.n1104 B.n49 585
R180 B.n777 B.n48 585
R181 B.n1105 B.n48 585
R182 B.n776 B.n775 585
R183 B.n775 B.n44 585
R184 B.n774 B.n43 585
R185 B.n1111 B.n43 585
R186 B.n773 B.n42 585
R187 B.n1112 B.n42 585
R188 B.n772 B.n41 585
R189 B.n1113 B.n41 585
R190 B.n771 B.n770 585
R191 B.n770 B.n40 585
R192 B.n769 B.n36 585
R193 B.n1119 B.n36 585
R194 B.n768 B.n35 585
R195 B.n1120 B.n35 585
R196 B.n767 B.n34 585
R197 B.n1121 B.n34 585
R198 B.n766 B.n765 585
R199 B.n765 B.n30 585
R200 B.n764 B.n29 585
R201 B.n1127 B.n29 585
R202 B.n763 B.n28 585
R203 B.n1128 B.n28 585
R204 B.n762 B.n27 585
R205 B.n1129 B.n27 585
R206 B.n761 B.n760 585
R207 B.n760 B.n23 585
R208 B.n759 B.n22 585
R209 B.n1135 B.n22 585
R210 B.n758 B.n21 585
R211 B.n1136 B.n21 585
R212 B.n757 B.n20 585
R213 B.n1137 B.n20 585
R214 B.n756 B.n755 585
R215 B.n755 B.n19 585
R216 B.n754 B.n15 585
R217 B.n1143 B.n15 585
R218 B.n753 B.n14 585
R219 B.n1144 B.n14 585
R220 B.n752 B.n13 585
R221 B.n1145 B.n13 585
R222 B.n751 B.n750 585
R223 B.n750 B.n12 585
R224 B.n749 B.n748 585
R225 B.n749 B.n8 585
R226 B.n747 B.n7 585
R227 B.n1152 B.n7 585
R228 B.n746 B.n6 585
R229 B.n1153 B.n6 585
R230 B.n745 B.n5 585
R231 B.n1154 B.n5 585
R232 B.n744 B.n743 585
R233 B.n743 B.n4 585
R234 B.n742 B.n174 585
R235 B.n742 B.n741 585
R236 B.n732 B.n175 585
R237 B.n176 B.n175 585
R238 B.n734 B.n733 585
R239 B.n735 B.n734 585
R240 B.n731 B.n181 585
R241 B.n181 B.n180 585
R242 B.n730 B.n729 585
R243 B.n729 B.n728 585
R244 B.n183 B.n182 585
R245 B.n721 B.n183 585
R246 B.n720 B.n719 585
R247 B.n722 B.n720 585
R248 B.n718 B.n188 585
R249 B.n188 B.n187 585
R250 B.n717 B.n716 585
R251 B.n716 B.n715 585
R252 B.n190 B.n189 585
R253 B.n191 B.n190 585
R254 B.n708 B.n707 585
R255 B.n709 B.n708 585
R256 B.n706 B.n196 585
R257 B.n196 B.n195 585
R258 B.n705 B.n704 585
R259 B.n704 B.n703 585
R260 B.n198 B.n197 585
R261 B.n199 B.n198 585
R262 B.n696 B.n695 585
R263 B.n697 B.n696 585
R264 B.n694 B.n204 585
R265 B.n204 B.n203 585
R266 B.n693 B.n692 585
R267 B.n692 B.n691 585
R268 B.n206 B.n205 585
R269 B.n684 B.n206 585
R270 B.n683 B.n682 585
R271 B.n685 B.n683 585
R272 B.n681 B.n211 585
R273 B.n211 B.n210 585
R274 B.n680 B.n679 585
R275 B.n679 B.n678 585
R276 B.n213 B.n212 585
R277 B.n214 B.n213 585
R278 B.n671 B.n670 585
R279 B.n672 B.n671 585
R280 B.n669 B.n219 585
R281 B.n219 B.n218 585
R282 B.n668 B.n667 585
R283 B.n667 B.n666 585
R284 B.n221 B.n220 585
R285 B.n222 B.n221 585
R286 B.n659 B.n658 585
R287 B.n660 B.n659 585
R288 B.n657 B.n227 585
R289 B.n227 B.n226 585
R290 B.n656 B.n655 585
R291 B.n655 B.n654 585
R292 B.n229 B.n228 585
R293 B.n647 B.n229 585
R294 B.n646 B.n645 585
R295 B.n648 B.n646 585
R296 B.n644 B.n234 585
R297 B.n234 B.n233 585
R298 B.n643 B.n642 585
R299 B.n642 B.n641 585
R300 B.n236 B.n235 585
R301 B.n237 B.n236 585
R302 B.n634 B.n633 585
R303 B.n635 B.n634 585
R304 B.n632 B.n242 585
R305 B.n242 B.n241 585
R306 B.n631 B.n630 585
R307 B.n630 B.n629 585
R308 B.n244 B.n243 585
R309 B.n245 B.n244 585
R310 B.n622 B.n621 585
R311 B.n623 B.n622 585
R312 B.n620 B.n250 585
R313 B.n250 B.n249 585
R314 B.n619 B.n618 585
R315 B.n618 B.n617 585
R316 B.n252 B.n251 585
R317 B.n610 B.n252 585
R318 B.n609 B.n608 585
R319 B.n611 B.n609 585
R320 B.n607 B.n257 585
R321 B.n257 B.n256 585
R322 B.n606 B.n605 585
R323 B.n605 B.n604 585
R324 B.n259 B.n258 585
R325 B.n260 B.n259 585
R326 B.n597 B.n596 585
R327 B.n598 B.n597 585
R328 B.n595 B.n265 585
R329 B.n265 B.n264 585
R330 B.n594 B.n593 585
R331 B.n593 B.n592 585
R332 B.n267 B.n266 585
R333 B.n268 B.n267 585
R334 B.n585 B.n584 585
R335 B.n586 B.n585 585
R336 B.n583 B.n273 585
R337 B.n273 B.n272 585
R338 B.n582 B.n581 585
R339 B.n581 B.n580 585
R340 B.n275 B.n274 585
R341 B.n276 B.n275 585
R342 B.n573 B.n572 585
R343 B.n574 B.n573 585
R344 B.n571 B.n280 585
R345 B.n284 B.n280 585
R346 B.n570 B.n569 585
R347 B.n569 B.n568 585
R348 B.n282 B.n281 585
R349 B.n283 B.n282 585
R350 B.n561 B.n560 585
R351 B.n562 B.n561 585
R352 B.n559 B.n289 585
R353 B.n289 B.n288 585
R354 B.n558 B.n557 585
R355 B.n557 B.n556 585
R356 B.n291 B.n290 585
R357 B.n292 B.n291 585
R358 B.n549 B.n548 585
R359 B.n550 B.n549 585
R360 B.n547 B.n297 585
R361 B.n297 B.n296 585
R362 B.n546 B.n545 585
R363 B.n545 B.n544 585
R364 B.n541 B.n301 585
R365 B.n540 B.n539 585
R366 B.n537 B.n302 585
R367 B.n537 B.n300 585
R368 B.n536 B.n535 585
R369 B.n534 B.n533 585
R370 B.n532 B.n304 585
R371 B.n530 B.n529 585
R372 B.n528 B.n305 585
R373 B.n527 B.n526 585
R374 B.n524 B.n306 585
R375 B.n522 B.n521 585
R376 B.n520 B.n307 585
R377 B.n519 B.n518 585
R378 B.n516 B.n308 585
R379 B.n514 B.n513 585
R380 B.n512 B.n309 585
R381 B.n511 B.n510 585
R382 B.n508 B.n310 585
R383 B.n506 B.n505 585
R384 B.n504 B.n311 585
R385 B.n503 B.n502 585
R386 B.n500 B.n312 585
R387 B.n498 B.n497 585
R388 B.n496 B.n313 585
R389 B.n495 B.n494 585
R390 B.n492 B.n314 585
R391 B.n490 B.n489 585
R392 B.n488 B.n315 585
R393 B.n487 B.n486 585
R394 B.n484 B.n316 585
R395 B.n482 B.n481 585
R396 B.n480 B.n317 585
R397 B.n479 B.n478 585
R398 B.n476 B.n318 585
R399 B.n474 B.n473 585
R400 B.n472 B.n319 585
R401 B.n471 B.n470 585
R402 B.n468 B.n320 585
R403 B.n466 B.n465 585
R404 B.n464 B.n321 585
R405 B.n463 B.n462 585
R406 B.n460 B.n322 585
R407 B.n458 B.n457 585
R408 B.n455 B.n323 585
R409 B.n454 B.n453 585
R410 B.n451 B.n326 585
R411 B.n449 B.n448 585
R412 B.n447 B.n327 585
R413 B.n446 B.n445 585
R414 B.n443 B.n328 585
R415 B.n441 B.n440 585
R416 B.n439 B.n329 585
R417 B.n437 B.n436 585
R418 B.n434 B.n332 585
R419 B.n432 B.n431 585
R420 B.n430 B.n333 585
R421 B.n429 B.n428 585
R422 B.n426 B.n334 585
R423 B.n424 B.n423 585
R424 B.n422 B.n335 585
R425 B.n421 B.n420 585
R426 B.n418 B.n336 585
R427 B.n416 B.n415 585
R428 B.n414 B.n337 585
R429 B.n413 B.n412 585
R430 B.n410 B.n338 585
R431 B.n408 B.n407 585
R432 B.n406 B.n339 585
R433 B.n405 B.n404 585
R434 B.n402 B.n340 585
R435 B.n400 B.n399 585
R436 B.n398 B.n341 585
R437 B.n397 B.n396 585
R438 B.n394 B.n342 585
R439 B.n392 B.n391 585
R440 B.n390 B.n343 585
R441 B.n389 B.n388 585
R442 B.n386 B.n344 585
R443 B.n384 B.n383 585
R444 B.n382 B.n345 585
R445 B.n381 B.n380 585
R446 B.n378 B.n346 585
R447 B.n376 B.n375 585
R448 B.n374 B.n347 585
R449 B.n373 B.n372 585
R450 B.n370 B.n348 585
R451 B.n368 B.n367 585
R452 B.n366 B.n349 585
R453 B.n365 B.n364 585
R454 B.n362 B.n350 585
R455 B.n360 B.n359 585
R456 B.n358 B.n351 585
R457 B.n357 B.n356 585
R458 B.n354 B.n352 585
R459 B.n299 B.n298 585
R460 B.n543 B.n542 585
R461 B.n544 B.n543 585
R462 B.n295 B.n294 585
R463 B.n296 B.n295 585
R464 B.n552 B.n551 585
R465 B.n551 B.n550 585
R466 B.n553 B.n293 585
R467 B.n293 B.n292 585
R468 B.n555 B.n554 585
R469 B.n556 B.n555 585
R470 B.n287 B.n286 585
R471 B.n288 B.n287 585
R472 B.n564 B.n563 585
R473 B.n563 B.n562 585
R474 B.n565 B.n285 585
R475 B.n285 B.n283 585
R476 B.n567 B.n566 585
R477 B.n568 B.n567 585
R478 B.n279 B.n278 585
R479 B.n284 B.n279 585
R480 B.n576 B.n575 585
R481 B.n575 B.n574 585
R482 B.n577 B.n277 585
R483 B.n277 B.n276 585
R484 B.n579 B.n578 585
R485 B.n580 B.n579 585
R486 B.n271 B.n270 585
R487 B.n272 B.n271 585
R488 B.n588 B.n587 585
R489 B.n587 B.n586 585
R490 B.n589 B.n269 585
R491 B.n269 B.n268 585
R492 B.n591 B.n590 585
R493 B.n592 B.n591 585
R494 B.n263 B.n262 585
R495 B.n264 B.n263 585
R496 B.n600 B.n599 585
R497 B.n599 B.n598 585
R498 B.n601 B.n261 585
R499 B.n261 B.n260 585
R500 B.n603 B.n602 585
R501 B.n604 B.n603 585
R502 B.n255 B.n254 585
R503 B.n256 B.n255 585
R504 B.n613 B.n612 585
R505 B.n612 B.n611 585
R506 B.n614 B.n253 585
R507 B.n610 B.n253 585
R508 B.n616 B.n615 585
R509 B.n617 B.n616 585
R510 B.n248 B.n247 585
R511 B.n249 B.n248 585
R512 B.n625 B.n624 585
R513 B.n624 B.n623 585
R514 B.n626 B.n246 585
R515 B.n246 B.n245 585
R516 B.n628 B.n627 585
R517 B.n629 B.n628 585
R518 B.n240 B.n239 585
R519 B.n241 B.n240 585
R520 B.n637 B.n636 585
R521 B.n636 B.n635 585
R522 B.n638 B.n238 585
R523 B.n238 B.n237 585
R524 B.n640 B.n639 585
R525 B.n641 B.n640 585
R526 B.n232 B.n231 585
R527 B.n233 B.n232 585
R528 B.n650 B.n649 585
R529 B.n649 B.n648 585
R530 B.n651 B.n230 585
R531 B.n647 B.n230 585
R532 B.n653 B.n652 585
R533 B.n654 B.n653 585
R534 B.n225 B.n224 585
R535 B.n226 B.n225 585
R536 B.n662 B.n661 585
R537 B.n661 B.n660 585
R538 B.n663 B.n223 585
R539 B.n223 B.n222 585
R540 B.n665 B.n664 585
R541 B.n666 B.n665 585
R542 B.n217 B.n216 585
R543 B.n218 B.n217 585
R544 B.n674 B.n673 585
R545 B.n673 B.n672 585
R546 B.n675 B.n215 585
R547 B.n215 B.n214 585
R548 B.n677 B.n676 585
R549 B.n678 B.n677 585
R550 B.n209 B.n208 585
R551 B.n210 B.n209 585
R552 B.n687 B.n686 585
R553 B.n686 B.n685 585
R554 B.n688 B.n207 585
R555 B.n684 B.n207 585
R556 B.n690 B.n689 585
R557 B.n691 B.n690 585
R558 B.n202 B.n201 585
R559 B.n203 B.n202 585
R560 B.n699 B.n698 585
R561 B.n698 B.n697 585
R562 B.n700 B.n200 585
R563 B.n200 B.n199 585
R564 B.n702 B.n701 585
R565 B.n703 B.n702 585
R566 B.n194 B.n193 585
R567 B.n195 B.n194 585
R568 B.n711 B.n710 585
R569 B.n710 B.n709 585
R570 B.n712 B.n192 585
R571 B.n192 B.n191 585
R572 B.n714 B.n713 585
R573 B.n715 B.n714 585
R574 B.n186 B.n185 585
R575 B.n187 B.n186 585
R576 B.n724 B.n723 585
R577 B.n723 B.n722 585
R578 B.n725 B.n184 585
R579 B.n721 B.n184 585
R580 B.n727 B.n726 585
R581 B.n728 B.n727 585
R582 B.n179 B.n178 585
R583 B.n180 B.n179 585
R584 B.n737 B.n736 585
R585 B.n736 B.n735 585
R586 B.n738 B.n177 585
R587 B.n177 B.n176 585
R588 B.n740 B.n739 585
R589 B.n741 B.n740 585
R590 B.n3 B.n0 585
R591 B.n4 B.n3 585
R592 B.n1151 B.n1 585
R593 B.n1152 B.n1151 585
R594 B.n1150 B.n1149 585
R595 B.n1150 B.n8 585
R596 B.n1148 B.n9 585
R597 B.n12 B.n9 585
R598 B.n1147 B.n1146 585
R599 B.n1146 B.n1145 585
R600 B.n11 B.n10 585
R601 B.n1144 B.n11 585
R602 B.n1142 B.n1141 585
R603 B.n1143 B.n1142 585
R604 B.n1140 B.n16 585
R605 B.n19 B.n16 585
R606 B.n1139 B.n1138 585
R607 B.n1138 B.n1137 585
R608 B.n18 B.n17 585
R609 B.n1136 B.n18 585
R610 B.n1134 B.n1133 585
R611 B.n1135 B.n1134 585
R612 B.n1132 B.n24 585
R613 B.n24 B.n23 585
R614 B.n1131 B.n1130 585
R615 B.n1130 B.n1129 585
R616 B.n26 B.n25 585
R617 B.n1128 B.n26 585
R618 B.n1126 B.n1125 585
R619 B.n1127 B.n1126 585
R620 B.n1124 B.n31 585
R621 B.n31 B.n30 585
R622 B.n1123 B.n1122 585
R623 B.n1122 B.n1121 585
R624 B.n33 B.n32 585
R625 B.n1120 B.n33 585
R626 B.n1118 B.n1117 585
R627 B.n1119 B.n1118 585
R628 B.n1116 B.n37 585
R629 B.n40 B.n37 585
R630 B.n1115 B.n1114 585
R631 B.n1114 B.n1113 585
R632 B.n39 B.n38 585
R633 B.n1112 B.n39 585
R634 B.n1110 B.n1109 585
R635 B.n1111 B.n1110 585
R636 B.n1108 B.n45 585
R637 B.n45 B.n44 585
R638 B.n1107 B.n1106 585
R639 B.n1106 B.n1105 585
R640 B.n47 B.n46 585
R641 B.n1104 B.n47 585
R642 B.n1102 B.n1101 585
R643 B.n1103 B.n1102 585
R644 B.n1100 B.n52 585
R645 B.n52 B.n51 585
R646 B.n1099 B.n1098 585
R647 B.n1098 B.n1097 585
R648 B.n54 B.n53 585
R649 B.n1096 B.n54 585
R650 B.n1094 B.n1093 585
R651 B.n1095 B.n1094 585
R652 B.n1092 B.n58 585
R653 B.n61 B.n58 585
R654 B.n1091 B.n1090 585
R655 B.n1090 B.n1089 585
R656 B.n60 B.n59 585
R657 B.n1088 B.n60 585
R658 B.n1086 B.n1085 585
R659 B.n1087 B.n1086 585
R660 B.n1084 B.n66 585
R661 B.n66 B.n65 585
R662 B.n1083 B.n1082 585
R663 B.n1082 B.n1081 585
R664 B.n68 B.n67 585
R665 B.n1080 B.n68 585
R666 B.n1078 B.n1077 585
R667 B.n1079 B.n1078 585
R668 B.n1076 B.n73 585
R669 B.n73 B.n72 585
R670 B.n1075 B.n1074 585
R671 B.n1074 B.n1073 585
R672 B.n75 B.n74 585
R673 B.n1072 B.n75 585
R674 B.n1070 B.n1069 585
R675 B.n1071 B.n1070 585
R676 B.n1068 B.n79 585
R677 B.n82 B.n79 585
R678 B.n1067 B.n1066 585
R679 B.n1066 B.n1065 585
R680 B.n81 B.n80 585
R681 B.n1064 B.n81 585
R682 B.n1062 B.n1061 585
R683 B.n1063 B.n1062 585
R684 B.n1060 B.n87 585
R685 B.n87 B.n86 585
R686 B.n1059 B.n1058 585
R687 B.n1058 B.n1057 585
R688 B.n89 B.n88 585
R689 B.n1056 B.n89 585
R690 B.n1054 B.n1053 585
R691 B.n1055 B.n1054 585
R692 B.n1052 B.n94 585
R693 B.n94 B.n93 585
R694 B.n1051 B.n1050 585
R695 B.n1050 B.n1049 585
R696 B.n96 B.n95 585
R697 B.n1048 B.n96 585
R698 B.n1046 B.n1045 585
R699 B.n1047 B.n1046 585
R700 B.n1044 B.n101 585
R701 B.n101 B.n100 585
R702 B.n1043 B.n1042 585
R703 B.n1042 B.n1041 585
R704 B.n103 B.n102 585
R705 B.n1040 B.n103 585
R706 B.n1038 B.n1037 585
R707 B.n1039 B.n1038 585
R708 B.n1036 B.n108 585
R709 B.n108 B.n107 585
R710 B.n1035 B.n1034 585
R711 B.n1034 B.n1033 585
R712 B.n110 B.n109 585
R713 B.n1032 B.n110 585
R714 B.n1030 B.n1029 585
R715 B.n1031 B.n1030 585
R716 B.n1028 B.n115 585
R717 B.n115 B.n114 585
R718 B.n1027 B.n1026 585
R719 B.n1026 B.n1025 585
R720 B.n117 B.n116 585
R721 B.n1024 B.n117 585
R722 B.n1022 B.n1021 585
R723 B.n1023 B.n1022 585
R724 B.n1155 B.n1154 585
R725 B.n1153 B.n2 585
R726 B.n1022 B.n122 564.573
R727 B.n831 B.n120 564.573
R728 B.n545 B.n299 564.573
R729 B.n543 B.n301 564.573
R730 B.n145 B.t19 291.493
R731 B.n152 B.t12 291.493
R732 B.n330 B.t8 291.493
R733 B.n324 B.t16 291.493
R734 B.n832 B.n121 256.663
R735 B.n838 B.n121 256.663
R736 B.n840 B.n121 256.663
R737 B.n846 B.n121 256.663
R738 B.n848 B.n121 256.663
R739 B.n854 B.n121 256.663
R740 B.n856 B.n121 256.663
R741 B.n862 B.n121 256.663
R742 B.n864 B.n121 256.663
R743 B.n870 B.n121 256.663
R744 B.n872 B.n121 256.663
R745 B.n878 B.n121 256.663
R746 B.n880 B.n121 256.663
R747 B.n886 B.n121 256.663
R748 B.n888 B.n121 256.663
R749 B.n894 B.n121 256.663
R750 B.n896 B.n121 256.663
R751 B.n902 B.n121 256.663
R752 B.n904 B.n121 256.663
R753 B.n910 B.n121 256.663
R754 B.n912 B.n121 256.663
R755 B.n919 B.n121 256.663
R756 B.n921 B.n121 256.663
R757 B.n927 B.n121 256.663
R758 B.n929 B.n121 256.663
R759 B.n935 B.n121 256.663
R760 B.n937 B.n121 256.663
R761 B.n943 B.n121 256.663
R762 B.n945 B.n121 256.663
R763 B.n951 B.n121 256.663
R764 B.n953 B.n121 256.663
R765 B.n959 B.n121 256.663
R766 B.n961 B.n121 256.663
R767 B.n967 B.n121 256.663
R768 B.n969 B.n121 256.663
R769 B.n975 B.n121 256.663
R770 B.n977 B.n121 256.663
R771 B.n983 B.n121 256.663
R772 B.n985 B.n121 256.663
R773 B.n991 B.n121 256.663
R774 B.n993 B.n121 256.663
R775 B.n999 B.n121 256.663
R776 B.n1001 B.n121 256.663
R777 B.n1007 B.n121 256.663
R778 B.n1009 B.n121 256.663
R779 B.n1015 B.n121 256.663
R780 B.n1017 B.n121 256.663
R781 B.n538 B.n300 256.663
R782 B.n303 B.n300 256.663
R783 B.n531 B.n300 256.663
R784 B.n525 B.n300 256.663
R785 B.n523 B.n300 256.663
R786 B.n517 B.n300 256.663
R787 B.n515 B.n300 256.663
R788 B.n509 B.n300 256.663
R789 B.n507 B.n300 256.663
R790 B.n501 B.n300 256.663
R791 B.n499 B.n300 256.663
R792 B.n493 B.n300 256.663
R793 B.n491 B.n300 256.663
R794 B.n485 B.n300 256.663
R795 B.n483 B.n300 256.663
R796 B.n477 B.n300 256.663
R797 B.n475 B.n300 256.663
R798 B.n469 B.n300 256.663
R799 B.n467 B.n300 256.663
R800 B.n461 B.n300 256.663
R801 B.n459 B.n300 256.663
R802 B.n452 B.n300 256.663
R803 B.n450 B.n300 256.663
R804 B.n444 B.n300 256.663
R805 B.n442 B.n300 256.663
R806 B.n435 B.n300 256.663
R807 B.n433 B.n300 256.663
R808 B.n427 B.n300 256.663
R809 B.n425 B.n300 256.663
R810 B.n419 B.n300 256.663
R811 B.n417 B.n300 256.663
R812 B.n411 B.n300 256.663
R813 B.n409 B.n300 256.663
R814 B.n403 B.n300 256.663
R815 B.n401 B.n300 256.663
R816 B.n395 B.n300 256.663
R817 B.n393 B.n300 256.663
R818 B.n387 B.n300 256.663
R819 B.n385 B.n300 256.663
R820 B.n379 B.n300 256.663
R821 B.n377 B.n300 256.663
R822 B.n371 B.n300 256.663
R823 B.n369 B.n300 256.663
R824 B.n363 B.n300 256.663
R825 B.n361 B.n300 256.663
R826 B.n355 B.n300 256.663
R827 B.n353 B.n300 256.663
R828 B.n1157 B.n1156 256.663
R829 B.n1018 B.n1016 163.367
R830 B.n1014 B.n124 163.367
R831 B.n1010 B.n1008 163.367
R832 B.n1006 B.n126 163.367
R833 B.n1002 B.n1000 163.367
R834 B.n998 B.n128 163.367
R835 B.n994 B.n992 163.367
R836 B.n990 B.n130 163.367
R837 B.n986 B.n984 163.367
R838 B.n982 B.n132 163.367
R839 B.n978 B.n976 163.367
R840 B.n974 B.n134 163.367
R841 B.n970 B.n968 163.367
R842 B.n966 B.n136 163.367
R843 B.n962 B.n960 163.367
R844 B.n958 B.n138 163.367
R845 B.n954 B.n952 163.367
R846 B.n950 B.n140 163.367
R847 B.n946 B.n944 163.367
R848 B.n942 B.n142 163.367
R849 B.n938 B.n936 163.367
R850 B.n934 B.n144 163.367
R851 B.n930 B.n928 163.367
R852 B.n926 B.n149 163.367
R853 B.n922 B.n920 163.367
R854 B.n918 B.n151 163.367
R855 B.n913 B.n911 163.367
R856 B.n909 B.n155 163.367
R857 B.n905 B.n903 163.367
R858 B.n901 B.n157 163.367
R859 B.n897 B.n895 163.367
R860 B.n893 B.n159 163.367
R861 B.n889 B.n887 163.367
R862 B.n885 B.n161 163.367
R863 B.n881 B.n879 163.367
R864 B.n877 B.n163 163.367
R865 B.n873 B.n871 163.367
R866 B.n869 B.n165 163.367
R867 B.n865 B.n863 163.367
R868 B.n861 B.n167 163.367
R869 B.n857 B.n855 163.367
R870 B.n853 B.n169 163.367
R871 B.n849 B.n847 163.367
R872 B.n845 B.n171 163.367
R873 B.n841 B.n839 163.367
R874 B.n837 B.n173 163.367
R875 B.n833 B.n831 163.367
R876 B.n545 B.n297 163.367
R877 B.n549 B.n297 163.367
R878 B.n549 B.n291 163.367
R879 B.n557 B.n291 163.367
R880 B.n557 B.n289 163.367
R881 B.n561 B.n289 163.367
R882 B.n561 B.n282 163.367
R883 B.n569 B.n282 163.367
R884 B.n569 B.n280 163.367
R885 B.n573 B.n280 163.367
R886 B.n573 B.n275 163.367
R887 B.n581 B.n275 163.367
R888 B.n581 B.n273 163.367
R889 B.n585 B.n273 163.367
R890 B.n585 B.n267 163.367
R891 B.n593 B.n267 163.367
R892 B.n593 B.n265 163.367
R893 B.n597 B.n265 163.367
R894 B.n597 B.n259 163.367
R895 B.n605 B.n259 163.367
R896 B.n605 B.n257 163.367
R897 B.n609 B.n257 163.367
R898 B.n609 B.n252 163.367
R899 B.n618 B.n252 163.367
R900 B.n618 B.n250 163.367
R901 B.n622 B.n250 163.367
R902 B.n622 B.n244 163.367
R903 B.n630 B.n244 163.367
R904 B.n630 B.n242 163.367
R905 B.n634 B.n242 163.367
R906 B.n634 B.n236 163.367
R907 B.n642 B.n236 163.367
R908 B.n642 B.n234 163.367
R909 B.n646 B.n234 163.367
R910 B.n646 B.n229 163.367
R911 B.n655 B.n229 163.367
R912 B.n655 B.n227 163.367
R913 B.n659 B.n227 163.367
R914 B.n659 B.n221 163.367
R915 B.n667 B.n221 163.367
R916 B.n667 B.n219 163.367
R917 B.n671 B.n219 163.367
R918 B.n671 B.n213 163.367
R919 B.n679 B.n213 163.367
R920 B.n679 B.n211 163.367
R921 B.n683 B.n211 163.367
R922 B.n683 B.n206 163.367
R923 B.n692 B.n206 163.367
R924 B.n692 B.n204 163.367
R925 B.n696 B.n204 163.367
R926 B.n696 B.n198 163.367
R927 B.n704 B.n198 163.367
R928 B.n704 B.n196 163.367
R929 B.n708 B.n196 163.367
R930 B.n708 B.n190 163.367
R931 B.n716 B.n190 163.367
R932 B.n716 B.n188 163.367
R933 B.n720 B.n188 163.367
R934 B.n720 B.n183 163.367
R935 B.n729 B.n183 163.367
R936 B.n729 B.n181 163.367
R937 B.n734 B.n181 163.367
R938 B.n734 B.n175 163.367
R939 B.n742 B.n175 163.367
R940 B.n743 B.n742 163.367
R941 B.n743 B.n5 163.367
R942 B.n6 B.n5 163.367
R943 B.n7 B.n6 163.367
R944 B.n749 B.n7 163.367
R945 B.n750 B.n749 163.367
R946 B.n750 B.n13 163.367
R947 B.n14 B.n13 163.367
R948 B.n15 B.n14 163.367
R949 B.n755 B.n15 163.367
R950 B.n755 B.n20 163.367
R951 B.n21 B.n20 163.367
R952 B.n22 B.n21 163.367
R953 B.n760 B.n22 163.367
R954 B.n760 B.n27 163.367
R955 B.n28 B.n27 163.367
R956 B.n29 B.n28 163.367
R957 B.n765 B.n29 163.367
R958 B.n765 B.n34 163.367
R959 B.n35 B.n34 163.367
R960 B.n36 B.n35 163.367
R961 B.n770 B.n36 163.367
R962 B.n770 B.n41 163.367
R963 B.n42 B.n41 163.367
R964 B.n43 B.n42 163.367
R965 B.n775 B.n43 163.367
R966 B.n775 B.n48 163.367
R967 B.n49 B.n48 163.367
R968 B.n50 B.n49 163.367
R969 B.n780 B.n50 163.367
R970 B.n780 B.n55 163.367
R971 B.n56 B.n55 163.367
R972 B.n57 B.n56 163.367
R973 B.n785 B.n57 163.367
R974 B.n785 B.n62 163.367
R975 B.n63 B.n62 163.367
R976 B.n64 B.n63 163.367
R977 B.n790 B.n64 163.367
R978 B.n790 B.n69 163.367
R979 B.n70 B.n69 163.367
R980 B.n71 B.n70 163.367
R981 B.n795 B.n71 163.367
R982 B.n795 B.n76 163.367
R983 B.n77 B.n76 163.367
R984 B.n78 B.n77 163.367
R985 B.n800 B.n78 163.367
R986 B.n800 B.n83 163.367
R987 B.n84 B.n83 163.367
R988 B.n85 B.n84 163.367
R989 B.n805 B.n85 163.367
R990 B.n805 B.n90 163.367
R991 B.n91 B.n90 163.367
R992 B.n92 B.n91 163.367
R993 B.n810 B.n92 163.367
R994 B.n810 B.n97 163.367
R995 B.n98 B.n97 163.367
R996 B.n99 B.n98 163.367
R997 B.n815 B.n99 163.367
R998 B.n815 B.n104 163.367
R999 B.n105 B.n104 163.367
R1000 B.n106 B.n105 163.367
R1001 B.n820 B.n106 163.367
R1002 B.n820 B.n111 163.367
R1003 B.n112 B.n111 163.367
R1004 B.n113 B.n112 163.367
R1005 B.n825 B.n113 163.367
R1006 B.n825 B.n118 163.367
R1007 B.n119 B.n118 163.367
R1008 B.n120 B.n119 163.367
R1009 B.n539 B.n537 163.367
R1010 B.n537 B.n536 163.367
R1011 B.n533 B.n532 163.367
R1012 B.n530 B.n305 163.367
R1013 B.n526 B.n524 163.367
R1014 B.n522 B.n307 163.367
R1015 B.n518 B.n516 163.367
R1016 B.n514 B.n309 163.367
R1017 B.n510 B.n508 163.367
R1018 B.n506 B.n311 163.367
R1019 B.n502 B.n500 163.367
R1020 B.n498 B.n313 163.367
R1021 B.n494 B.n492 163.367
R1022 B.n490 B.n315 163.367
R1023 B.n486 B.n484 163.367
R1024 B.n482 B.n317 163.367
R1025 B.n478 B.n476 163.367
R1026 B.n474 B.n319 163.367
R1027 B.n470 B.n468 163.367
R1028 B.n466 B.n321 163.367
R1029 B.n462 B.n460 163.367
R1030 B.n458 B.n323 163.367
R1031 B.n453 B.n451 163.367
R1032 B.n449 B.n327 163.367
R1033 B.n445 B.n443 163.367
R1034 B.n441 B.n329 163.367
R1035 B.n436 B.n434 163.367
R1036 B.n432 B.n333 163.367
R1037 B.n428 B.n426 163.367
R1038 B.n424 B.n335 163.367
R1039 B.n420 B.n418 163.367
R1040 B.n416 B.n337 163.367
R1041 B.n412 B.n410 163.367
R1042 B.n408 B.n339 163.367
R1043 B.n404 B.n402 163.367
R1044 B.n400 B.n341 163.367
R1045 B.n396 B.n394 163.367
R1046 B.n392 B.n343 163.367
R1047 B.n388 B.n386 163.367
R1048 B.n384 B.n345 163.367
R1049 B.n380 B.n378 163.367
R1050 B.n376 B.n347 163.367
R1051 B.n372 B.n370 163.367
R1052 B.n368 B.n349 163.367
R1053 B.n364 B.n362 163.367
R1054 B.n360 B.n351 163.367
R1055 B.n356 B.n354 163.367
R1056 B.n543 B.n295 163.367
R1057 B.n551 B.n295 163.367
R1058 B.n551 B.n293 163.367
R1059 B.n555 B.n293 163.367
R1060 B.n555 B.n287 163.367
R1061 B.n563 B.n287 163.367
R1062 B.n563 B.n285 163.367
R1063 B.n567 B.n285 163.367
R1064 B.n567 B.n279 163.367
R1065 B.n575 B.n279 163.367
R1066 B.n575 B.n277 163.367
R1067 B.n579 B.n277 163.367
R1068 B.n579 B.n271 163.367
R1069 B.n587 B.n271 163.367
R1070 B.n587 B.n269 163.367
R1071 B.n591 B.n269 163.367
R1072 B.n591 B.n263 163.367
R1073 B.n599 B.n263 163.367
R1074 B.n599 B.n261 163.367
R1075 B.n603 B.n261 163.367
R1076 B.n603 B.n255 163.367
R1077 B.n612 B.n255 163.367
R1078 B.n612 B.n253 163.367
R1079 B.n616 B.n253 163.367
R1080 B.n616 B.n248 163.367
R1081 B.n624 B.n248 163.367
R1082 B.n624 B.n246 163.367
R1083 B.n628 B.n246 163.367
R1084 B.n628 B.n240 163.367
R1085 B.n636 B.n240 163.367
R1086 B.n636 B.n238 163.367
R1087 B.n640 B.n238 163.367
R1088 B.n640 B.n232 163.367
R1089 B.n649 B.n232 163.367
R1090 B.n649 B.n230 163.367
R1091 B.n653 B.n230 163.367
R1092 B.n653 B.n225 163.367
R1093 B.n661 B.n225 163.367
R1094 B.n661 B.n223 163.367
R1095 B.n665 B.n223 163.367
R1096 B.n665 B.n217 163.367
R1097 B.n673 B.n217 163.367
R1098 B.n673 B.n215 163.367
R1099 B.n677 B.n215 163.367
R1100 B.n677 B.n209 163.367
R1101 B.n686 B.n209 163.367
R1102 B.n686 B.n207 163.367
R1103 B.n690 B.n207 163.367
R1104 B.n690 B.n202 163.367
R1105 B.n698 B.n202 163.367
R1106 B.n698 B.n200 163.367
R1107 B.n702 B.n200 163.367
R1108 B.n702 B.n194 163.367
R1109 B.n710 B.n194 163.367
R1110 B.n710 B.n192 163.367
R1111 B.n714 B.n192 163.367
R1112 B.n714 B.n186 163.367
R1113 B.n723 B.n186 163.367
R1114 B.n723 B.n184 163.367
R1115 B.n727 B.n184 163.367
R1116 B.n727 B.n179 163.367
R1117 B.n736 B.n179 163.367
R1118 B.n736 B.n177 163.367
R1119 B.n740 B.n177 163.367
R1120 B.n740 B.n3 163.367
R1121 B.n1155 B.n3 163.367
R1122 B.n1151 B.n2 163.367
R1123 B.n1151 B.n1150 163.367
R1124 B.n1150 B.n9 163.367
R1125 B.n1146 B.n9 163.367
R1126 B.n1146 B.n11 163.367
R1127 B.n1142 B.n11 163.367
R1128 B.n1142 B.n16 163.367
R1129 B.n1138 B.n16 163.367
R1130 B.n1138 B.n18 163.367
R1131 B.n1134 B.n18 163.367
R1132 B.n1134 B.n24 163.367
R1133 B.n1130 B.n24 163.367
R1134 B.n1130 B.n26 163.367
R1135 B.n1126 B.n26 163.367
R1136 B.n1126 B.n31 163.367
R1137 B.n1122 B.n31 163.367
R1138 B.n1122 B.n33 163.367
R1139 B.n1118 B.n33 163.367
R1140 B.n1118 B.n37 163.367
R1141 B.n1114 B.n37 163.367
R1142 B.n1114 B.n39 163.367
R1143 B.n1110 B.n39 163.367
R1144 B.n1110 B.n45 163.367
R1145 B.n1106 B.n45 163.367
R1146 B.n1106 B.n47 163.367
R1147 B.n1102 B.n47 163.367
R1148 B.n1102 B.n52 163.367
R1149 B.n1098 B.n52 163.367
R1150 B.n1098 B.n54 163.367
R1151 B.n1094 B.n54 163.367
R1152 B.n1094 B.n58 163.367
R1153 B.n1090 B.n58 163.367
R1154 B.n1090 B.n60 163.367
R1155 B.n1086 B.n60 163.367
R1156 B.n1086 B.n66 163.367
R1157 B.n1082 B.n66 163.367
R1158 B.n1082 B.n68 163.367
R1159 B.n1078 B.n68 163.367
R1160 B.n1078 B.n73 163.367
R1161 B.n1074 B.n73 163.367
R1162 B.n1074 B.n75 163.367
R1163 B.n1070 B.n75 163.367
R1164 B.n1070 B.n79 163.367
R1165 B.n1066 B.n79 163.367
R1166 B.n1066 B.n81 163.367
R1167 B.n1062 B.n81 163.367
R1168 B.n1062 B.n87 163.367
R1169 B.n1058 B.n87 163.367
R1170 B.n1058 B.n89 163.367
R1171 B.n1054 B.n89 163.367
R1172 B.n1054 B.n94 163.367
R1173 B.n1050 B.n94 163.367
R1174 B.n1050 B.n96 163.367
R1175 B.n1046 B.n96 163.367
R1176 B.n1046 B.n101 163.367
R1177 B.n1042 B.n101 163.367
R1178 B.n1042 B.n103 163.367
R1179 B.n1038 B.n103 163.367
R1180 B.n1038 B.n108 163.367
R1181 B.n1034 B.n108 163.367
R1182 B.n1034 B.n110 163.367
R1183 B.n1030 B.n110 163.367
R1184 B.n1030 B.n115 163.367
R1185 B.n1026 B.n115 163.367
R1186 B.n1026 B.n117 163.367
R1187 B.n1022 B.n117 163.367
R1188 B.n152 B.t14 149.185
R1189 B.n330 B.t11 149.185
R1190 B.n145 B.t20 149.168
R1191 B.n324 B.t18 149.168
R1192 B.n544 B.n300 82.4927
R1193 B.n1023 B.n121 82.4927
R1194 B.n146 B.n145 77.1884
R1195 B.n153 B.n152 77.1884
R1196 B.n331 B.n330 77.1884
R1197 B.n325 B.n324 77.1884
R1198 B.n153 B.t15 71.9961
R1199 B.n331 B.t10 71.9961
R1200 B.n146 B.t21 71.9804
R1201 B.n325 B.t17 71.9804
R1202 B.n1017 B.n122 71.676
R1203 B.n1016 B.n1015 71.676
R1204 B.n1009 B.n124 71.676
R1205 B.n1008 B.n1007 71.676
R1206 B.n1001 B.n126 71.676
R1207 B.n1000 B.n999 71.676
R1208 B.n993 B.n128 71.676
R1209 B.n992 B.n991 71.676
R1210 B.n985 B.n130 71.676
R1211 B.n984 B.n983 71.676
R1212 B.n977 B.n132 71.676
R1213 B.n976 B.n975 71.676
R1214 B.n969 B.n134 71.676
R1215 B.n968 B.n967 71.676
R1216 B.n961 B.n136 71.676
R1217 B.n960 B.n959 71.676
R1218 B.n953 B.n138 71.676
R1219 B.n952 B.n951 71.676
R1220 B.n945 B.n140 71.676
R1221 B.n944 B.n943 71.676
R1222 B.n937 B.n142 71.676
R1223 B.n936 B.n935 71.676
R1224 B.n929 B.n144 71.676
R1225 B.n928 B.n927 71.676
R1226 B.n921 B.n149 71.676
R1227 B.n920 B.n919 71.676
R1228 B.n912 B.n151 71.676
R1229 B.n911 B.n910 71.676
R1230 B.n904 B.n155 71.676
R1231 B.n903 B.n902 71.676
R1232 B.n896 B.n157 71.676
R1233 B.n895 B.n894 71.676
R1234 B.n888 B.n159 71.676
R1235 B.n887 B.n886 71.676
R1236 B.n880 B.n161 71.676
R1237 B.n879 B.n878 71.676
R1238 B.n872 B.n163 71.676
R1239 B.n871 B.n870 71.676
R1240 B.n864 B.n165 71.676
R1241 B.n863 B.n862 71.676
R1242 B.n856 B.n167 71.676
R1243 B.n855 B.n854 71.676
R1244 B.n848 B.n169 71.676
R1245 B.n847 B.n846 71.676
R1246 B.n840 B.n171 71.676
R1247 B.n839 B.n838 71.676
R1248 B.n832 B.n173 71.676
R1249 B.n833 B.n832 71.676
R1250 B.n838 B.n837 71.676
R1251 B.n841 B.n840 71.676
R1252 B.n846 B.n845 71.676
R1253 B.n849 B.n848 71.676
R1254 B.n854 B.n853 71.676
R1255 B.n857 B.n856 71.676
R1256 B.n862 B.n861 71.676
R1257 B.n865 B.n864 71.676
R1258 B.n870 B.n869 71.676
R1259 B.n873 B.n872 71.676
R1260 B.n878 B.n877 71.676
R1261 B.n881 B.n880 71.676
R1262 B.n886 B.n885 71.676
R1263 B.n889 B.n888 71.676
R1264 B.n894 B.n893 71.676
R1265 B.n897 B.n896 71.676
R1266 B.n902 B.n901 71.676
R1267 B.n905 B.n904 71.676
R1268 B.n910 B.n909 71.676
R1269 B.n913 B.n912 71.676
R1270 B.n919 B.n918 71.676
R1271 B.n922 B.n921 71.676
R1272 B.n927 B.n926 71.676
R1273 B.n930 B.n929 71.676
R1274 B.n935 B.n934 71.676
R1275 B.n938 B.n937 71.676
R1276 B.n943 B.n942 71.676
R1277 B.n946 B.n945 71.676
R1278 B.n951 B.n950 71.676
R1279 B.n954 B.n953 71.676
R1280 B.n959 B.n958 71.676
R1281 B.n962 B.n961 71.676
R1282 B.n967 B.n966 71.676
R1283 B.n970 B.n969 71.676
R1284 B.n975 B.n974 71.676
R1285 B.n978 B.n977 71.676
R1286 B.n983 B.n982 71.676
R1287 B.n986 B.n985 71.676
R1288 B.n991 B.n990 71.676
R1289 B.n994 B.n993 71.676
R1290 B.n999 B.n998 71.676
R1291 B.n1002 B.n1001 71.676
R1292 B.n1007 B.n1006 71.676
R1293 B.n1010 B.n1009 71.676
R1294 B.n1015 B.n1014 71.676
R1295 B.n1018 B.n1017 71.676
R1296 B.n538 B.n301 71.676
R1297 B.n536 B.n303 71.676
R1298 B.n532 B.n531 71.676
R1299 B.n525 B.n305 71.676
R1300 B.n524 B.n523 71.676
R1301 B.n517 B.n307 71.676
R1302 B.n516 B.n515 71.676
R1303 B.n509 B.n309 71.676
R1304 B.n508 B.n507 71.676
R1305 B.n501 B.n311 71.676
R1306 B.n500 B.n499 71.676
R1307 B.n493 B.n313 71.676
R1308 B.n492 B.n491 71.676
R1309 B.n485 B.n315 71.676
R1310 B.n484 B.n483 71.676
R1311 B.n477 B.n317 71.676
R1312 B.n476 B.n475 71.676
R1313 B.n469 B.n319 71.676
R1314 B.n468 B.n467 71.676
R1315 B.n461 B.n321 71.676
R1316 B.n460 B.n459 71.676
R1317 B.n452 B.n323 71.676
R1318 B.n451 B.n450 71.676
R1319 B.n444 B.n327 71.676
R1320 B.n443 B.n442 71.676
R1321 B.n435 B.n329 71.676
R1322 B.n434 B.n433 71.676
R1323 B.n427 B.n333 71.676
R1324 B.n426 B.n425 71.676
R1325 B.n419 B.n335 71.676
R1326 B.n418 B.n417 71.676
R1327 B.n411 B.n337 71.676
R1328 B.n410 B.n409 71.676
R1329 B.n403 B.n339 71.676
R1330 B.n402 B.n401 71.676
R1331 B.n395 B.n341 71.676
R1332 B.n394 B.n393 71.676
R1333 B.n387 B.n343 71.676
R1334 B.n386 B.n385 71.676
R1335 B.n379 B.n345 71.676
R1336 B.n378 B.n377 71.676
R1337 B.n371 B.n347 71.676
R1338 B.n370 B.n369 71.676
R1339 B.n363 B.n349 71.676
R1340 B.n362 B.n361 71.676
R1341 B.n355 B.n351 71.676
R1342 B.n354 B.n353 71.676
R1343 B.n539 B.n538 71.676
R1344 B.n533 B.n303 71.676
R1345 B.n531 B.n530 71.676
R1346 B.n526 B.n525 71.676
R1347 B.n523 B.n522 71.676
R1348 B.n518 B.n517 71.676
R1349 B.n515 B.n514 71.676
R1350 B.n510 B.n509 71.676
R1351 B.n507 B.n506 71.676
R1352 B.n502 B.n501 71.676
R1353 B.n499 B.n498 71.676
R1354 B.n494 B.n493 71.676
R1355 B.n491 B.n490 71.676
R1356 B.n486 B.n485 71.676
R1357 B.n483 B.n482 71.676
R1358 B.n478 B.n477 71.676
R1359 B.n475 B.n474 71.676
R1360 B.n470 B.n469 71.676
R1361 B.n467 B.n466 71.676
R1362 B.n462 B.n461 71.676
R1363 B.n459 B.n458 71.676
R1364 B.n453 B.n452 71.676
R1365 B.n450 B.n449 71.676
R1366 B.n445 B.n444 71.676
R1367 B.n442 B.n441 71.676
R1368 B.n436 B.n435 71.676
R1369 B.n433 B.n432 71.676
R1370 B.n428 B.n427 71.676
R1371 B.n425 B.n424 71.676
R1372 B.n420 B.n419 71.676
R1373 B.n417 B.n416 71.676
R1374 B.n412 B.n411 71.676
R1375 B.n409 B.n408 71.676
R1376 B.n404 B.n403 71.676
R1377 B.n401 B.n400 71.676
R1378 B.n396 B.n395 71.676
R1379 B.n393 B.n392 71.676
R1380 B.n388 B.n387 71.676
R1381 B.n385 B.n384 71.676
R1382 B.n380 B.n379 71.676
R1383 B.n377 B.n376 71.676
R1384 B.n372 B.n371 71.676
R1385 B.n369 B.n368 71.676
R1386 B.n364 B.n363 71.676
R1387 B.n361 B.n360 71.676
R1388 B.n356 B.n355 71.676
R1389 B.n353 B.n299 71.676
R1390 B.n1156 B.n1155 71.676
R1391 B.n1156 B.n2 71.676
R1392 B.n147 B.n146 59.5399
R1393 B.n916 B.n153 59.5399
R1394 B.n438 B.n331 59.5399
R1395 B.n456 B.n325 59.5399
R1396 B.n544 B.n296 42.177
R1397 B.n550 B.n296 42.177
R1398 B.n550 B.n292 42.177
R1399 B.n556 B.n292 42.177
R1400 B.n556 B.n288 42.177
R1401 B.n562 B.n288 42.177
R1402 B.n562 B.n283 42.177
R1403 B.n568 B.n283 42.177
R1404 B.n568 B.n284 42.177
R1405 B.n574 B.n276 42.177
R1406 B.n580 B.n276 42.177
R1407 B.n580 B.n272 42.177
R1408 B.n586 B.n272 42.177
R1409 B.n586 B.n268 42.177
R1410 B.n592 B.n268 42.177
R1411 B.n592 B.n264 42.177
R1412 B.n598 B.n264 42.177
R1413 B.n598 B.n260 42.177
R1414 B.n604 B.n260 42.177
R1415 B.n604 B.n256 42.177
R1416 B.n611 B.n256 42.177
R1417 B.n611 B.n610 42.177
R1418 B.n617 B.n249 42.177
R1419 B.n623 B.n249 42.177
R1420 B.n623 B.n245 42.177
R1421 B.n629 B.n245 42.177
R1422 B.n629 B.n241 42.177
R1423 B.n635 B.n241 42.177
R1424 B.n635 B.n237 42.177
R1425 B.n641 B.n237 42.177
R1426 B.n641 B.n233 42.177
R1427 B.n648 B.n233 42.177
R1428 B.n648 B.n647 42.177
R1429 B.n654 B.n226 42.177
R1430 B.n660 B.n226 42.177
R1431 B.n660 B.n222 42.177
R1432 B.n666 B.n222 42.177
R1433 B.n666 B.n218 42.177
R1434 B.n672 B.n218 42.177
R1435 B.n672 B.n214 42.177
R1436 B.n678 B.n214 42.177
R1437 B.n678 B.n210 42.177
R1438 B.n685 B.n210 42.177
R1439 B.n685 B.n684 42.177
R1440 B.n691 B.n203 42.177
R1441 B.n697 B.n203 42.177
R1442 B.n697 B.n199 42.177
R1443 B.n703 B.n199 42.177
R1444 B.n703 B.n195 42.177
R1445 B.n709 B.n195 42.177
R1446 B.n709 B.n191 42.177
R1447 B.n715 B.n191 42.177
R1448 B.n715 B.n187 42.177
R1449 B.n722 B.n187 42.177
R1450 B.n722 B.n721 42.177
R1451 B.n728 B.n180 42.177
R1452 B.n735 B.n180 42.177
R1453 B.n735 B.n176 42.177
R1454 B.n741 B.n176 42.177
R1455 B.n741 B.n4 42.177
R1456 B.n1154 B.n4 42.177
R1457 B.n1154 B.n1153 42.177
R1458 B.n1153 B.n1152 42.177
R1459 B.n1152 B.n8 42.177
R1460 B.n12 B.n8 42.177
R1461 B.n1145 B.n12 42.177
R1462 B.n1145 B.n1144 42.177
R1463 B.n1144 B.n1143 42.177
R1464 B.n1137 B.n19 42.177
R1465 B.n1137 B.n1136 42.177
R1466 B.n1136 B.n1135 42.177
R1467 B.n1135 B.n23 42.177
R1468 B.n1129 B.n23 42.177
R1469 B.n1129 B.n1128 42.177
R1470 B.n1128 B.n1127 42.177
R1471 B.n1127 B.n30 42.177
R1472 B.n1121 B.n30 42.177
R1473 B.n1121 B.n1120 42.177
R1474 B.n1120 B.n1119 42.177
R1475 B.n1113 B.n40 42.177
R1476 B.n1113 B.n1112 42.177
R1477 B.n1112 B.n1111 42.177
R1478 B.n1111 B.n44 42.177
R1479 B.n1105 B.n44 42.177
R1480 B.n1105 B.n1104 42.177
R1481 B.n1104 B.n1103 42.177
R1482 B.n1103 B.n51 42.177
R1483 B.n1097 B.n51 42.177
R1484 B.n1097 B.n1096 42.177
R1485 B.n1096 B.n1095 42.177
R1486 B.n1089 B.n61 42.177
R1487 B.n1089 B.n1088 42.177
R1488 B.n1088 B.n1087 42.177
R1489 B.n1087 B.n65 42.177
R1490 B.n1081 B.n65 42.177
R1491 B.n1081 B.n1080 42.177
R1492 B.n1080 B.n1079 42.177
R1493 B.n1079 B.n72 42.177
R1494 B.n1073 B.n72 42.177
R1495 B.n1073 B.n1072 42.177
R1496 B.n1072 B.n1071 42.177
R1497 B.n1065 B.n82 42.177
R1498 B.n1065 B.n1064 42.177
R1499 B.n1064 B.n1063 42.177
R1500 B.n1063 B.n86 42.177
R1501 B.n1057 B.n86 42.177
R1502 B.n1057 B.n1056 42.177
R1503 B.n1056 B.n1055 42.177
R1504 B.n1055 B.n93 42.177
R1505 B.n1049 B.n93 42.177
R1506 B.n1049 B.n1048 42.177
R1507 B.n1048 B.n1047 42.177
R1508 B.n1047 B.n100 42.177
R1509 B.n1041 B.n100 42.177
R1510 B.n1040 B.n1039 42.177
R1511 B.n1039 B.n107 42.177
R1512 B.n1033 B.n107 42.177
R1513 B.n1033 B.n1032 42.177
R1514 B.n1032 B.n1031 42.177
R1515 B.n1031 B.n114 42.177
R1516 B.n1025 B.n114 42.177
R1517 B.n1025 B.n1024 42.177
R1518 B.n1024 B.n1023 42.177
R1519 B.n574 B.t9 41.5567
R1520 B.n1041 B.t13 41.5567
R1521 B.n728 B.t2 40.3163
R1522 B.n1143 B.t7 40.3163
R1523 B.n610 B.t4 39.0758
R1524 B.n82 B.t5 39.0758
R1525 B.n542 B.n541 36.6834
R1526 B.n546 B.n298 36.6834
R1527 B.n1021 B.n1020 36.6834
R1528 B.n830 B.n829 36.6834
R1529 B.n691 B.t6 27.9114
R1530 B.n1119 B.t0 27.9114
R1531 B.n647 B.t1 26.6709
R1532 B.n61 B.t3 26.6709
R1533 B B.n1157 18.0485
R1534 B.n654 B.t1 15.5066
R1535 B.n1095 B.t3 15.5066
R1536 B.n684 B.t6 14.2661
R1537 B.n40 B.t0 14.2661
R1538 B.n542 B.n294 10.6151
R1539 B.n552 B.n294 10.6151
R1540 B.n553 B.n552 10.6151
R1541 B.n554 B.n553 10.6151
R1542 B.n554 B.n286 10.6151
R1543 B.n564 B.n286 10.6151
R1544 B.n565 B.n564 10.6151
R1545 B.n566 B.n565 10.6151
R1546 B.n566 B.n278 10.6151
R1547 B.n576 B.n278 10.6151
R1548 B.n577 B.n576 10.6151
R1549 B.n578 B.n577 10.6151
R1550 B.n578 B.n270 10.6151
R1551 B.n588 B.n270 10.6151
R1552 B.n589 B.n588 10.6151
R1553 B.n590 B.n589 10.6151
R1554 B.n590 B.n262 10.6151
R1555 B.n600 B.n262 10.6151
R1556 B.n601 B.n600 10.6151
R1557 B.n602 B.n601 10.6151
R1558 B.n602 B.n254 10.6151
R1559 B.n613 B.n254 10.6151
R1560 B.n614 B.n613 10.6151
R1561 B.n615 B.n614 10.6151
R1562 B.n615 B.n247 10.6151
R1563 B.n625 B.n247 10.6151
R1564 B.n626 B.n625 10.6151
R1565 B.n627 B.n626 10.6151
R1566 B.n627 B.n239 10.6151
R1567 B.n637 B.n239 10.6151
R1568 B.n638 B.n637 10.6151
R1569 B.n639 B.n638 10.6151
R1570 B.n639 B.n231 10.6151
R1571 B.n650 B.n231 10.6151
R1572 B.n651 B.n650 10.6151
R1573 B.n652 B.n651 10.6151
R1574 B.n652 B.n224 10.6151
R1575 B.n662 B.n224 10.6151
R1576 B.n663 B.n662 10.6151
R1577 B.n664 B.n663 10.6151
R1578 B.n664 B.n216 10.6151
R1579 B.n674 B.n216 10.6151
R1580 B.n675 B.n674 10.6151
R1581 B.n676 B.n675 10.6151
R1582 B.n676 B.n208 10.6151
R1583 B.n687 B.n208 10.6151
R1584 B.n688 B.n687 10.6151
R1585 B.n689 B.n688 10.6151
R1586 B.n689 B.n201 10.6151
R1587 B.n699 B.n201 10.6151
R1588 B.n700 B.n699 10.6151
R1589 B.n701 B.n700 10.6151
R1590 B.n701 B.n193 10.6151
R1591 B.n711 B.n193 10.6151
R1592 B.n712 B.n711 10.6151
R1593 B.n713 B.n712 10.6151
R1594 B.n713 B.n185 10.6151
R1595 B.n724 B.n185 10.6151
R1596 B.n725 B.n724 10.6151
R1597 B.n726 B.n725 10.6151
R1598 B.n726 B.n178 10.6151
R1599 B.n737 B.n178 10.6151
R1600 B.n738 B.n737 10.6151
R1601 B.n739 B.n738 10.6151
R1602 B.n739 B.n0 10.6151
R1603 B.n541 B.n540 10.6151
R1604 B.n540 B.n302 10.6151
R1605 B.n535 B.n302 10.6151
R1606 B.n535 B.n534 10.6151
R1607 B.n534 B.n304 10.6151
R1608 B.n529 B.n304 10.6151
R1609 B.n529 B.n528 10.6151
R1610 B.n528 B.n527 10.6151
R1611 B.n527 B.n306 10.6151
R1612 B.n521 B.n306 10.6151
R1613 B.n521 B.n520 10.6151
R1614 B.n520 B.n519 10.6151
R1615 B.n519 B.n308 10.6151
R1616 B.n513 B.n308 10.6151
R1617 B.n513 B.n512 10.6151
R1618 B.n512 B.n511 10.6151
R1619 B.n511 B.n310 10.6151
R1620 B.n505 B.n310 10.6151
R1621 B.n505 B.n504 10.6151
R1622 B.n504 B.n503 10.6151
R1623 B.n503 B.n312 10.6151
R1624 B.n497 B.n312 10.6151
R1625 B.n497 B.n496 10.6151
R1626 B.n496 B.n495 10.6151
R1627 B.n495 B.n314 10.6151
R1628 B.n489 B.n314 10.6151
R1629 B.n489 B.n488 10.6151
R1630 B.n488 B.n487 10.6151
R1631 B.n487 B.n316 10.6151
R1632 B.n481 B.n316 10.6151
R1633 B.n481 B.n480 10.6151
R1634 B.n480 B.n479 10.6151
R1635 B.n479 B.n318 10.6151
R1636 B.n473 B.n318 10.6151
R1637 B.n473 B.n472 10.6151
R1638 B.n472 B.n471 10.6151
R1639 B.n471 B.n320 10.6151
R1640 B.n465 B.n320 10.6151
R1641 B.n465 B.n464 10.6151
R1642 B.n464 B.n463 10.6151
R1643 B.n463 B.n322 10.6151
R1644 B.n457 B.n322 10.6151
R1645 B.n455 B.n454 10.6151
R1646 B.n454 B.n326 10.6151
R1647 B.n448 B.n326 10.6151
R1648 B.n448 B.n447 10.6151
R1649 B.n447 B.n446 10.6151
R1650 B.n446 B.n328 10.6151
R1651 B.n440 B.n328 10.6151
R1652 B.n440 B.n439 10.6151
R1653 B.n437 B.n332 10.6151
R1654 B.n431 B.n332 10.6151
R1655 B.n431 B.n430 10.6151
R1656 B.n430 B.n429 10.6151
R1657 B.n429 B.n334 10.6151
R1658 B.n423 B.n334 10.6151
R1659 B.n423 B.n422 10.6151
R1660 B.n422 B.n421 10.6151
R1661 B.n421 B.n336 10.6151
R1662 B.n415 B.n336 10.6151
R1663 B.n415 B.n414 10.6151
R1664 B.n414 B.n413 10.6151
R1665 B.n413 B.n338 10.6151
R1666 B.n407 B.n338 10.6151
R1667 B.n407 B.n406 10.6151
R1668 B.n406 B.n405 10.6151
R1669 B.n405 B.n340 10.6151
R1670 B.n399 B.n340 10.6151
R1671 B.n399 B.n398 10.6151
R1672 B.n398 B.n397 10.6151
R1673 B.n397 B.n342 10.6151
R1674 B.n391 B.n342 10.6151
R1675 B.n391 B.n390 10.6151
R1676 B.n390 B.n389 10.6151
R1677 B.n389 B.n344 10.6151
R1678 B.n383 B.n344 10.6151
R1679 B.n383 B.n382 10.6151
R1680 B.n382 B.n381 10.6151
R1681 B.n381 B.n346 10.6151
R1682 B.n375 B.n346 10.6151
R1683 B.n375 B.n374 10.6151
R1684 B.n374 B.n373 10.6151
R1685 B.n373 B.n348 10.6151
R1686 B.n367 B.n348 10.6151
R1687 B.n367 B.n366 10.6151
R1688 B.n366 B.n365 10.6151
R1689 B.n365 B.n350 10.6151
R1690 B.n359 B.n350 10.6151
R1691 B.n359 B.n358 10.6151
R1692 B.n358 B.n357 10.6151
R1693 B.n357 B.n352 10.6151
R1694 B.n352 B.n298 10.6151
R1695 B.n547 B.n546 10.6151
R1696 B.n548 B.n547 10.6151
R1697 B.n548 B.n290 10.6151
R1698 B.n558 B.n290 10.6151
R1699 B.n559 B.n558 10.6151
R1700 B.n560 B.n559 10.6151
R1701 B.n560 B.n281 10.6151
R1702 B.n570 B.n281 10.6151
R1703 B.n571 B.n570 10.6151
R1704 B.n572 B.n571 10.6151
R1705 B.n572 B.n274 10.6151
R1706 B.n582 B.n274 10.6151
R1707 B.n583 B.n582 10.6151
R1708 B.n584 B.n583 10.6151
R1709 B.n584 B.n266 10.6151
R1710 B.n594 B.n266 10.6151
R1711 B.n595 B.n594 10.6151
R1712 B.n596 B.n595 10.6151
R1713 B.n596 B.n258 10.6151
R1714 B.n606 B.n258 10.6151
R1715 B.n607 B.n606 10.6151
R1716 B.n608 B.n607 10.6151
R1717 B.n608 B.n251 10.6151
R1718 B.n619 B.n251 10.6151
R1719 B.n620 B.n619 10.6151
R1720 B.n621 B.n620 10.6151
R1721 B.n621 B.n243 10.6151
R1722 B.n631 B.n243 10.6151
R1723 B.n632 B.n631 10.6151
R1724 B.n633 B.n632 10.6151
R1725 B.n633 B.n235 10.6151
R1726 B.n643 B.n235 10.6151
R1727 B.n644 B.n643 10.6151
R1728 B.n645 B.n644 10.6151
R1729 B.n645 B.n228 10.6151
R1730 B.n656 B.n228 10.6151
R1731 B.n657 B.n656 10.6151
R1732 B.n658 B.n657 10.6151
R1733 B.n658 B.n220 10.6151
R1734 B.n668 B.n220 10.6151
R1735 B.n669 B.n668 10.6151
R1736 B.n670 B.n669 10.6151
R1737 B.n670 B.n212 10.6151
R1738 B.n680 B.n212 10.6151
R1739 B.n681 B.n680 10.6151
R1740 B.n682 B.n681 10.6151
R1741 B.n682 B.n205 10.6151
R1742 B.n693 B.n205 10.6151
R1743 B.n694 B.n693 10.6151
R1744 B.n695 B.n694 10.6151
R1745 B.n695 B.n197 10.6151
R1746 B.n705 B.n197 10.6151
R1747 B.n706 B.n705 10.6151
R1748 B.n707 B.n706 10.6151
R1749 B.n707 B.n189 10.6151
R1750 B.n717 B.n189 10.6151
R1751 B.n718 B.n717 10.6151
R1752 B.n719 B.n718 10.6151
R1753 B.n719 B.n182 10.6151
R1754 B.n730 B.n182 10.6151
R1755 B.n731 B.n730 10.6151
R1756 B.n733 B.n731 10.6151
R1757 B.n733 B.n732 10.6151
R1758 B.n732 B.n174 10.6151
R1759 B.n744 B.n174 10.6151
R1760 B.n745 B.n744 10.6151
R1761 B.n746 B.n745 10.6151
R1762 B.n747 B.n746 10.6151
R1763 B.n748 B.n747 10.6151
R1764 B.n751 B.n748 10.6151
R1765 B.n752 B.n751 10.6151
R1766 B.n753 B.n752 10.6151
R1767 B.n754 B.n753 10.6151
R1768 B.n756 B.n754 10.6151
R1769 B.n757 B.n756 10.6151
R1770 B.n758 B.n757 10.6151
R1771 B.n759 B.n758 10.6151
R1772 B.n761 B.n759 10.6151
R1773 B.n762 B.n761 10.6151
R1774 B.n763 B.n762 10.6151
R1775 B.n764 B.n763 10.6151
R1776 B.n766 B.n764 10.6151
R1777 B.n767 B.n766 10.6151
R1778 B.n768 B.n767 10.6151
R1779 B.n769 B.n768 10.6151
R1780 B.n771 B.n769 10.6151
R1781 B.n772 B.n771 10.6151
R1782 B.n773 B.n772 10.6151
R1783 B.n774 B.n773 10.6151
R1784 B.n776 B.n774 10.6151
R1785 B.n777 B.n776 10.6151
R1786 B.n778 B.n777 10.6151
R1787 B.n779 B.n778 10.6151
R1788 B.n781 B.n779 10.6151
R1789 B.n782 B.n781 10.6151
R1790 B.n783 B.n782 10.6151
R1791 B.n784 B.n783 10.6151
R1792 B.n786 B.n784 10.6151
R1793 B.n787 B.n786 10.6151
R1794 B.n788 B.n787 10.6151
R1795 B.n789 B.n788 10.6151
R1796 B.n791 B.n789 10.6151
R1797 B.n792 B.n791 10.6151
R1798 B.n793 B.n792 10.6151
R1799 B.n794 B.n793 10.6151
R1800 B.n796 B.n794 10.6151
R1801 B.n797 B.n796 10.6151
R1802 B.n798 B.n797 10.6151
R1803 B.n799 B.n798 10.6151
R1804 B.n801 B.n799 10.6151
R1805 B.n802 B.n801 10.6151
R1806 B.n803 B.n802 10.6151
R1807 B.n804 B.n803 10.6151
R1808 B.n806 B.n804 10.6151
R1809 B.n807 B.n806 10.6151
R1810 B.n808 B.n807 10.6151
R1811 B.n809 B.n808 10.6151
R1812 B.n811 B.n809 10.6151
R1813 B.n812 B.n811 10.6151
R1814 B.n813 B.n812 10.6151
R1815 B.n814 B.n813 10.6151
R1816 B.n816 B.n814 10.6151
R1817 B.n817 B.n816 10.6151
R1818 B.n818 B.n817 10.6151
R1819 B.n819 B.n818 10.6151
R1820 B.n821 B.n819 10.6151
R1821 B.n822 B.n821 10.6151
R1822 B.n823 B.n822 10.6151
R1823 B.n824 B.n823 10.6151
R1824 B.n826 B.n824 10.6151
R1825 B.n827 B.n826 10.6151
R1826 B.n828 B.n827 10.6151
R1827 B.n829 B.n828 10.6151
R1828 B.n1149 B.n1 10.6151
R1829 B.n1149 B.n1148 10.6151
R1830 B.n1148 B.n1147 10.6151
R1831 B.n1147 B.n10 10.6151
R1832 B.n1141 B.n10 10.6151
R1833 B.n1141 B.n1140 10.6151
R1834 B.n1140 B.n1139 10.6151
R1835 B.n1139 B.n17 10.6151
R1836 B.n1133 B.n17 10.6151
R1837 B.n1133 B.n1132 10.6151
R1838 B.n1132 B.n1131 10.6151
R1839 B.n1131 B.n25 10.6151
R1840 B.n1125 B.n25 10.6151
R1841 B.n1125 B.n1124 10.6151
R1842 B.n1124 B.n1123 10.6151
R1843 B.n1123 B.n32 10.6151
R1844 B.n1117 B.n32 10.6151
R1845 B.n1117 B.n1116 10.6151
R1846 B.n1116 B.n1115 10.6151
R1847 B.n1115 B.n38 10.6151
R1848 B.n1109 B.n38 10.6151
R1849 B.n1109 B.n1108 10.6151
R1850 B.n1108 B.n1107 10.6151
R1851 B.n1107 B.n46 10.6151
R1852 B.n1101 B.n46 10.6151
R1853 B.n1101 B.n1100 10.6151
R1854 B.n1100 B.n1099 10.6151
R1855 B.n1099 B.n53 10.6151
R1856 B.n1093 B.n53 10.6151
R1857 B.n1093 B.n1092 10.6151
R1858 B.n1092 B.n1091 10.6151
R1859 B.n1091 B.n59 10.6151
R1860 B.n1085 B.n59 10.6151
R1861 B.n1085 B.n1084 10.6151
R1862 B.n1084 B.n1083 10.6151
R1863 B.n1083 B.n67 10.6151
R1864 B.n1077 B.n67 10.6151
R1865 B.n1077 B.n1076 10.6151
R1866 B.n1076 B.n1075 10.6151
R1867 B.n1075 B.n74 10.6151
R1868 B.n1069 B.n74 10.6151
R1869 B.n1069 B.n1068 10.6151
R1870 B.n1068 B.n1067 10.6151
R1871 B.n1067 B.n80 10.6151
R1872 B.n1061 B.n80 10.6151
R1873 B.n1061 B.n1060 10.6151
R1874 B.n1060 B.n1059 10.6151
R1875 B.n1059 B.n88 10.6151
R1876 B.n1053 B.n88 10.6151
R1877 B.n1053 B.n1052 10.6151
R1878 B.n1052 B.n1051 10.6151
R1879 B.n1051 B.n95 10.6151
R1880 B.n1045 B.n95 10.6151
R1881 B.n1045 B.n1044 10.6151
R1882 B.n1044 B.n1043 10.6151
R1883 B.n1043 B.n102 10.6151
R1884 B.n1037 B.n102 10.6151
R1885 B.n1037 B.n1036 10.6151
R1886 B.n1036 B.n1035 10.6151
R1887 B.n1035 B.n109 10.6151
R1888 B.n1029 B.n109 10.6151
R1889 B.n1029 B.n1028 10.6151
R1890 B.n1028 B.n1027 10.6151
R1891 B.n1027 B.n116 10.6151
R1892 B.n1021 B.n116 10.6151
R1893 B.n1020 B.n1019 10.6151
R1894 B.n1019 B.n123 10.6151
R1895 B.n1013 B.n123 10.6151
R1896 B.n1013 B.n1012 10.6151
R1897 B.n1012 B.n1011 10.6151
R1898 B.n1011 B.n125 10.6151
R1899 B.n1005 B.n125 10.6151
R1900 B.n1005 B.n1004 10.6151
R1901 B.n1004 B.n1003 10.6151
R1902 B.n1003 B.n127 10.6151
R1903 B.n997 B.n127 10.6151
R1904 B.n997 B.n996 10.6151
R1905 B.n996 B.n995 10.6151
R1906 B.n995 B.n129 10.6151
R1907 B.n989 B.n129 10.6151
R1908 B.n989 B.n988 10.6151
R1909 B.n988 B.n987 10.6151
R1910 B.n987 B.n131 10.6151
R1911 B.n981 B.n131 10.6151
R1912 B.n981 B.n980 10.6151
R1913 B.n980 B.n979 10.6151
R1914 B.n979 B.n133 10.6151
R1915 B.n973 B.n133 10.6151
R1916 B.n973 B.n972 10.6151
R1917 B.n972 B.n971 10.6151
R1918 B.n971 B.n135 10.6151
R1919 B.n965 B.n135 10.6151
R1920 B.n965 B.n964 10.6151
R1921 B.n964 B.n963 10.6151
R1922 B.n963 B.n137 10.6151
R1923 B.n957 B.n137 10.6151
R1924 B.n957 B.n956 10.6151
R1925 B.n956 B.n955 10.6151
R1926 B.n955 B.n139 10.6151
R1927 B.n949 B.n139 10.6151
R1928 B.n949 B.n948 10.6151
R1929 B.n948 B.n947 10.6151
R1930 B.n947 B.n141 10.6151
R1931 B.n941 B.n141 10.6151
R1932 B.n941 B.n940 10.6151
R1933 B.n940 B.n939 10.6151
R1934 B.n939 B.n143 10.6151
R1935 B.n933 B.n932 10.6151
R1936 B.n932 B.n931 10.6151
R1937 B.n931 B.n148 10.6151
R1938 B.n925 B.n148 10.6151
R1939 B.n925 B.n924 10.6151
R1940 B.n924 B.n923 10.6151
R1941 B.n923 B.n150 10.6151
R1942 B.n917 B.n150 10.6151
R1943 B.n915 B.n914 10.6151
R1944 B.n914 B.n154 10.6151
R1945 B.n908 B.n154 10.6151
R1946 B.n908 B.n907 10.6151
R1947 B.n907 B.n906 10.6151
R1948 B.n906 B.n156 10.6151
R1949 B.n900 B.n156 10.6151
R1950 B.n900 B.n899 10.6151
R1951 B.n899 B.n898 10.6151
R1952 B.n898 B.n158 10.6151
R1953 B.n892 B.n158 10.6151
R1954 B.n892 B.n891 10.6151
R1955 B.n891 B.n890 10.6151
R1956 B.n890 B.n160 10.6151
R1957 B.n884 B.n160 10.6151
R1958 B.n884 B.n883 10.6151
R1959 B.n883 B.n882 10.6151
R1960 B.n882 B.n162 10.6151
R1961 B.n876 B.n162 10.6151
R1962 B.n876 B.n875 10.6151
R1963 B.n875 B.n874 10.6151
R1964 B.n874 B.n164 10.6151
R1965 B.n868 B.n164 10.6151
R1966 B.n868 B.n867 10.6151
R1967 B.n867 B.n866 10.6151
R1968 B.n866 B.n166 10.6151
R1969 B.n860 B.n166 10.6151
R1970 B.n860 B.n859 10.6151
R1971 B.n859 B.n858 10.6151
R1972 B.n858 B.n168 10.6151
R1973 B.n852 B.n168 10.6151
R1974 B.n852 B.n851 10.6151
R1975 B.n851 B.n850 10.6151
R1976 B.n850 B.n170 10.6151
R1977 B.n844 B.n170 10.6151
R1978 B.n844 B.n843 10.6151
R1979 B.n843 B.n842 10.6151
R1980 B.n842 B.n172 10.6151
R1981 B.n836 B.n172 10.6151
R1982 B.n836 B.n835 10.6151
R1983 B.n835 B.n834 10.6151
R1984 B.n834 B.n830 10.6151
R1985 B.n1157 B.n0 8.11757
R1986 B.n1157 B.n1 8.11757
R1987 B.n456 B.n455 6.5566
R1988 B.n439 B.n438 6.5566
R1989 B.n933 B.n147 6.5566
R1990 B.n917 B.n916 6.5566
R1991 B.n457 B.n456 4.05904
R1992 B.n438 B.n437 4.05904
R1993 B.n147 B.n143 4.05904
R1994 B.n916 B.n915 4.05904
R1995 B.n617 B.t4 3.10171
R1996 B.n1071 B.t5 3.10171
R1997 B.n721 B.t2 1.86123
R1998 B.n19 B.t7 1.86123
R1999 B.n284 B.t9 0.620742
R2000 B.t13 B.n1040 0.620742
R2001 VP.n24 VP.n21 161.3
R2002 VP.n26 VP.n25 161.3
R2003 VP.n27 VP.n20 161.3
R2004 VP.n29 VP.n28 161.3
R2005 VP.n30 VP.n19 161.3
R2006 VP.n32 VP.n31 161.3
R2007 VP.n33 VP.n18 161.3
R2008 VP.n36 VP.n35 161.3
R2009 VP.n37 VP.n17 161.3
R2010 VP.n39 VP.n38 161.3
R2011 VP.n40 VP.n16 161.3
R2012 VP.n42 VP.n41 161.3
R2013 VP.n43 VP.n15 161.3
R2014 VP.n45 VP.n44 161.3
R2015 VP.n46 VP.n14 161.3
R2016 VP.n48 VP.n47 161.3
R2017 VP.n89 VP.n88 161.3
R2018 VP.n87 VP.n1 161.3
R2019 VP.n86 VP.n85 161.3
R2020 VP.n84 VP.n2 161.3
R2021 VP.n83 VP.n82 161.3
R2022 VP.n81 VP.n3 161.3
R2023 VP.n80 VP.n79 161.3
R2024 VP.n78 VP.n4 161.3
R2025 VP.n77 VP.n76 161.3
R2026 VP.n74 VP.n5 161.3
R2027 VP.n73 VP.n72 161.3
R2028 VP.n71 VP.n6 161.3
R2029 VP.n70 VP.n69 161.3
R2030 VP.n68 VP.n7 161.3
R2031 VP.n67 VP.n66 161.3
R2032 VP.n65 VP.n8 161.3
R2033 VP.n64 VP.n63 161.3
R2034 VP.n61 VP.n9 161.3
R2035 VP.n60 VP.n59 161.3
R2036 VP.n58 VP.n10 161.3
R2037 VP.n57 VP.n56 161.3
R2038 VP.n55 VP.n11 161.3
R2039 VP.n54 VP.n53 161.3
R2040 VP.n52 VP.n12 161.3
R2041 VP.n23 VP.t5 115.698
R2042 VP.n50 VP.t7 82.2706
R2043 VP.n62 VP.t4 82.2706
R2044 VP.n75 VP.t1 82.2706
R2045 VP.n0 VP.t3 82.2706
R2046 VP.n13 VP.t6 82.2706
R2047 VP.n34 VP.t0 82.2706
R2048 VP.n22 VP.t2 82.2706
R2049 VP.n51 VP.n50 79.1799
R2050 VP.n90 VP.n0 79.1799
R2051 VP.n49 VP.n13 79.1799
R2052 VP.n23 VP.n22 62.7141
R2053 VP.n56 VP.n10 56.4773
R2054 VP.n41 VP.n15 56.4773
R2055 VP.n69 VP.n6 56.4773
R2056 VP.n82 VP.n2 56.4773
R2057 VP.n28 VP.n19 56.4773
R2058 VP.n51 VP.n49 56.2946
R2059 VP.n54 VP.n12 24.3439
R2060 VP.n55 VP.n54 24.3439
R2061 VP.n56 VP.n55 24.3439
R2062 VP.n60 VP.n10 24.3439
R2063 VP.n61 VP.n60 24.3439
R2064 VP.n63 VP.n61 24.3439
R2065 VP.n67 VP.n8 24.3439
R2066 VP.n68 VP.n67 24.3439
R2067 VP.n69 VP.n68 24.3439
R2068 VP.n73 VP.n6 24.3439
R2069 VP.n74 VP.n73 24.3439
R2070 VP.n76 VP.n74 24.3439
R2071 VP.n80 VP.n4 24.3439
R2072 VP.n81 VP.n80 24.3439
R2073 VP.n82 VP.n81 24.3439
R2074 VP.n86 VP.n2 24.3439
R2075 VP.n87 VP.n86 24.3439
R2076 VP.n88 VP.n87 24.3439
R2077 VP.n45 VP.n15 24.3439
R2078 VP.n46 VP.n45 24.3439
R2079 VP.n47 VP.n46 24.3439
R2080 VP.n32 VP.n19 24.3439
R2081 VP.n33 VP.n32 24.3439
R2082 VP.n35 VP.n33 24.3439
R2083 VP.n39 VP.n17 24.3439
R2084 VP.n40 VP.n39 24.3439
R2085 VP.n41 VP.n40 24.3439
R2086 VP.n26 VP.n21 24.3439
R2087 VP.n27 VP.n26 24.3439
R2088 VP.n28 VP.n27 24.3439
R2089 VP.n63 VP.n62 12.6591
R2090 VP.n75 VP.n4 12.6591
R2091 VP.n34 VP.n17 12.6591
R2092 VP.n62 VP.n8 11.6853
R2093 VP.n76 VP.n75 11.6853
R2094 VP.n35 VP.n34 11.6853
R2095 VP.n22 VP.n21 11.6853
R2096 VP.n50 VP.n12 10.7116
R2097 VP.n88 VP.n0 10.7116
R2098 VP.n47 VP.n13 10.7116
R2099 VP.n24 VP.n23 3.1448
R2100 VP.n49 VP.n48 0.355081
R2101 VP.n52 VP.n51 0.355081
R2102 VP.n90 VP.n89 0.355081
R2103 VP VP.n90 0.26685
R2104 VP.n25 VP.n24 0.189894
R2105 VP.n25 VP.n20 0.189894
R2106 VP.n29 VP.n20 0.189894
R2107 VP.n30 VP.n29 0.189894
R2108 VP.n31 VP.n30 0.189894
R2109 VP.n31 VP.n18 0.189894
R2110 VP.n36 VP.n18 0.189894
R2111 VP.n37 VP.n36 0.189894
R2112 VP.n38 VP.n37 0.189894
R2113 VP.n38 VP.n16 0.189894
R2114 VP.n42 VP.n16 0.189894
R2115 VP.n43 VP.n42 0.189894
R2116 VP.n44 VP.n43 0.189894
R2117 VP.n44 VP.n14 0.189894
R2118 VP.n48 VP.n14 0.189894
R2119 VP.n53 VP.n52 0.189894
R2120 VP.n53 VP.n11 0.189894
R2121 VP.n57 VP.n11 0.189894
R2122 VP.n58 VP.n57 0.189894
R2123 VP.n59 VP.n58 0.189894
R2124 VP.n59 VP.n9 0.189894
R2125 VP.n64 VP.n9 0.189894
R2126 VP.n65 VP.n64 0.189894
R2127 VP.n66 VP.n65 0.189894
R2128 VP.n66 VP.n7 0.189894
R2129 VP.n70 VP.n7 0.189894
R2130 VP.n71 VP.n70 0.189894
R2131 VP.n72 VP.n71 0.189894
R2132 VP.n72 VP.n5 0.189894
R2133 VP.n77 VP.n5 0.189894
R2134 VP.n78 VP.n77 0.189894
R2135 VP.n79 VP.n78 0.189894
R2136 VP.n79 VP.n3 0.189894
R2137 VP.n83 VP.n3 0.189894
R2138 VP.n84 VP.n83 0.189894
R2139 VP.n85 VP.n84 0.189894
R2140 VP.n85 VP.n1 0.189894
R2141 VP.n89 VP.n1 0.189894
R2142 VDD1 VDD1.n0 63.1734
R2143 VDD1.n3 VDD1.n2 63.0596
R2144 VDD1.n3 VDD1.n1 63.0596
R2145 VDD1.n5 VDD1.n4 61.3995
R2146 VDD1.n5 VDD1.n3 50.4793
R2147 VDD1 VDD1.n5 1.65783
R2148 VDD1.n4 VDD1.t0 1.58959
R2149 VDD1.n4 VDD1.t4 1.58959
R2150 VDD1.n0 VDD1.t5 1.58959
R2151 VDD1.n0 VDD1.t2 1.58959
R2152 VDD1.n2 VDD1.t1 1.58959
R2153 VDD1.n2 VDD1.t7 1.58959
R2154 VDD1.n1 VDD1.t6 1.58959
R2155 VDD1.n1 VDD1.t3 1.58959
R2156 VTAIL.n11 VTAIL.t10 46.3099
R2157 VTAIL.n10 VTAIL.t0 46.3099
R2158 VTAIL.n7 VTAIL.t2 46.3099
R2159 VTAIL.n15 VTAIL.t3 46.3098
R2160 VTAIL.n2 VTAIL.t7 46.3098
R2161 VTAIL.n3 VTAIL.t12 46.3098
R2162 VTAIL.n6 VTAIL.t8 46.3098
R2163 VTAIL.n14 VTAIL.t9 46.3098
R2164 VTAIL.n13 VTAIL.n12 44.7209
R2165 VTAIL.n9 VTAIL.n8 44.7209
R2166 VTAIL.n1 VTAIL.n0 44.7206
R2167 VTAIL.n5 VTAIL.n4 44.7206
R2168 VTAIL.n15 VTAIL.n14 26.5393
R2169 VTAIL.n7 VTAIL.n6 26.5393
R2170 VTAIL.n9 VTAIL.n7 3.43153
R2171 VTAIL.n10 VTAIL.n9 3.43153
R2172 VTAIL.n13 VTAIL.n11 3.43153
R2173 VTAIL.n14 VTAIL.n13 3.43153
R2174 VTAIL.n6 VTAIL.n5 3.43153
R2175 VTAIL.n5 VTAIL.n3 3.43153
R2176 VTAIL.n2 VTAIL.n1 3.43153
R2177 VTAIL VTAIL.n15 3.37334
R2178 VTAIL.n0 VTAIL.t6 1.58959
R2179 VTAIL.n0 VTAIL.t5 1.58959
R2180 VTAIL.n4 VTAIL.t11 1.58959
R2181 VTAIL.n4 VTAIL.t14 1.58959
R2182 VTAIL.n12 VTAIL.t13 1.58959
R2183 VTAIL.n12 VTAIL.t15 1.58959
R2184 VTAIL.n8 VTAIL.t1 1.58959
R2185 VTAIL.n8 VTAIL.t4 1.58959
R2186 VTAIL.n11 VTAIL.n10 0.470328
R2187 VTAIL.n3 VTAIL.n2 0.470328
R2188 VTAIL VTAIL.n1 0.0586897
R2189 VN.n72 VN.n71 161.3
R2190 VN.n70 VN.n38 161.3
R2191 VN.n69 VN.n68 161.3
R2192 VN.n67 VN.n39 161.3
R2193 VN.n66 VN.n65 161.3
R2194 VN.n64 VN.n40 161.3
R2195 VN.n63 VN.n62 161.3
R2196 VN.n61 VN.n41 161.3
R2197 VN.n60 VN.n59 161.3
R2198 VN.n58 VN.n42 161.3
R2199 VN.n57 VN.n56 161.3
R2200 VN.n55 VN.n44 161.3
R2201 VN.n54 VN.n53 161.3
R2202 VN.n52 VN.n45 161.3
R2203 VN.n51 VN.n50 161.3
R2204 VN.n49 VN.n46 161.3
R2205 VN.n35 VN.n34 161.3
R2206 VN.n33 VN.n1 161.3
R2207 VN.n32 VN.n31 161.3
R2208 VN.n30 VN.n2 161.3
R2209 VN.n29 VN.n28 161.3
R2210 VN.n27 VN.n3 161.3
R2211 VN.n26 VN.n25 161.3
R2212 VN.n24 VN.n4 161.3
R2213 VN.n23 VN.n22 161.3
R2214 VN.n20 VN.n5 161.3
R2215 VN.n19 VN.n18 161.3
R2216 VN.n17 VN.n6 161.3
R2217 VN.n16 VN.n15 161.3
R2218 VN.n14 VN.n7 161.3
R2219 VN.n13 VN.n12 161.3
R2220 VN.n11 VN.n8 161.3
R2221 VN.n48 VN.t7 115.698
R2222 VN.n10 VN.t3 115.698
R2223 VN.n9 VN.t2 82.2706
R2224 VN.n21 VN.t4 82.2706
R2225 VN.n0 VN.t0 82.2706
R2226 VN.n47 VN.t6 82.2706
R2227 VN.n43 VN.t5 82.2706
R2228 VN.n37 VN.t1 82.2706
R2229 VN.n36 VN.n0 79.1799
R2230 VN.n73 VN.n37 79.1799
R2231 VN.n10 VN.n9 62.7141
R2232 VN.n48 VN.n47 62.7141
R2233 VN.n15 VN.n6 56.4773
R2234 VN.n28 VN.n2 56.4773
R2235 VN.n53 VN.n44 56.4773
R2236 VN.n65 VN.n39 56.4773
R2237 VN VN.n73 56.46
R2238 VN.n13 VN.n8 24.3439
R2239 VN.n14 VN.n13 24.3439
R2240 VN.n15 VN.n14 24.3439
R2241 VN.n19 VN.n6 24.3439
R2242 VN.n20 VN.n19 24.3439
R2243 VN.n22 VN.n20 24.3439
R2244 VN.n26 VN.n4 24.3439
R2245 VN.n27 VN.n26 24.3439
R2246 VN.n28 VN.n27 24.3439
R2247 VN.n32 VN.n2 24.3439
R2248 VN.n33 VN.n32 24.3439
R2249 VN.n34 VN.n33 24.3439
R2250 VN.n53 VN.n52 24.3439
R2251 VN.n52 VN.n51 24.3439
R2252 VN.n51 VN.n46 24.3439
R2253 VN.n65 VN.n64 24.3439
R2254 VN.n64 VN.n63 24.3439
R2255 VN.n63 VN.n41 24.3439
R2256 VN.n59 VN.n58 24.3439
R2257 VN.n58 VN.n57 24.3439
R2258 VN.n57 VN.n44 24.3439
R2259 VN.n71 VN.n70 24.3439
R2260 VN.n70 VN.n69 24.3439
R2261 VN.n69 VN.n39 24.3439
R2262 VN.n21 VN.n4 12.6591
R2263 VN.n43 VN.n41 12.6591
R2264 VN.n9 VN.n8 11.6853
R2265 VN.n22 VN.n21 11.6853
R2266 VN.n47 VN.n46 11.6853
R2267 VN.n59 VN.n43 11.6853
R2268 VN.n34 VN.n0 10.7116
R2269 VN.n71 VN.n37 10.7116
R2270 VN.n49 VN.n48 3.14482
R2271 VN.n11 VN.n10 3.14482
R2272 VN.n73 VN.n72 0.355081
R2273 VN.n36 VN.n35 0.355081
R2274 VN VN.n36 0.26685
R2275 VN.n72 VN.n38 0.189894
R2276 VN.n68 VN.n38 0.189894
R2277 VN.n68 VN.n67 0.189894
R2278 VN.n67 VN.n66 0.189894
R2279 VN.n66 VN.n40 0.189894
R2280 VN.n62 VN.n40 0.189894
R2281 VN.n62 VN.n61 0.189894
R2282 VN.n61 VN.n60 0.189894
R2283 VN.n60 VN.n42 0.189894
R2284 VN.n56 VN.n42 0.189894
R2285 VN.n56 VN.n55 0.189894
R2286 VN.n55 VN.n54 0.189894
R2287 VN.n54 VN.n45 0.189894
R2288 VN.n50 VN.n45 0.189894
R2289 VN.n50 VN.n49 0.189894
R2290 VN.n12 VN.n11 0.189894
R2291 VN.n12 VN.n7 0.189894
R2292 VN.n16 VN.n7 0.189894
R2293 VN.n17 VN.n16 0.189894
R2294 VN.n18 VN.n17 0.189894
R2295 VN.n18 VN.n5 0.189894
R2296 VN.n23 VN.n5 0.189894
R2297 VN.n24 VN.n23 0.189894
R2298 VN.n25 VN.n24 0.189894
R2299 VN.n25 VN.n3 0.189894
R2300 VN.n29 VN.n3 0.189894
R2301 VN.n30 VN.n29 0.189894
R2302 VN.n31 VN.n30 0.189894
R2303 VN.n31 VN.n1 0.189894
R2304 VN.n35 VN.n1 0.189894
R2305 VDD2.n2 VDD2.n1 63.0596
R2306 VDD2.n2 VDD2.n0 63.0596
R2307 VDD2 VDD2.n5 63.0568
R2308 VDD2.n4 VDD2.n3 61.3997
R2309 VDD2.n4 VDD2.n2 49.8963
R2310 VDD2 VDD2.n4 1.77421
R2311 VDD2.n5 VDD2.t1 1.58959
R2312 VDD2.n5 VDD2.t0 1.58959
R2313 VDD2.n3 VDD2.t6 1.58959
R2314 VDD2.n3 VDD2.t2 1.58959
R2315 VDD2.n1 VDD2.t3 1.58959
R2316 VDD2.n1 VDD2.t7 1.58959
R2317 VDD2.n0 VDD2.t4 1.58959
R2318 VDD2.n0 VDD2.t5 1.58959
C0 VTAIL VP 10.276599f
C1 VDD1 VDD2 2.32301f
C2 VN VDD1 0.153436f
C3 VTAIL VDD1 8.64439f
C4 VP VDD1 10.0107f
C5 VN VDD2 9.53488f
C6 VTAIL VDD2 8.70585f
C7 VP VDD2 0.631212f
C8 VN VTAIL 10.262501f
C9 VN VP 9.03754f
C10 VDD2 B 6.492256f
C11 VDD1 B 7.04331f
C12 VTAIL B 11.473742f
C13 VN B 19.58943f
C14 VP B 18.246763f
C15 VDD2.t4 B 0.266047f
C16 VDD2.t5 B 0.266047f
C17 VDD2.n0 B 2.39313f
C18 VDD2.t3 B 0.266047f
C19 VDD2.t7 B 0.266047f
C20 VDD2.n1 B 2.39313f
C21 VDD2.n2 B 4.23455f
C22 VDD2.t6 B 0.266047f
C23 VDD2.t2 B 0.266047f
C24 VDD2.n3 B 2.37525f
C25 VDD2.n4 B 3.6227f
C26 VDD2.t1 B 0.266047f
C27 VDD2.t0 B 0.266047f
C28 VDD2.n5 B 2.39308f
C29 VN.t0 B 2.18798f
C30 VN.n0 B 0.837757f
C31 VN.n1 B 0.017639f
C32 VN.n2 B 0.026851f
C33 VN.n3 B 0.017639f
C34 VN.n4 B 0.025209f
C35 VN.n5 B 0.017639f
C36 VN.n6 B 0.025861f
C37 VN.n7 B 0.017639f
C38 VN.n8 B 0.024556f
C39 VN.t2 B 2.18798f
C40 VN.n9 B 0.827434f
C41 VN.t3 B 2.44873f
C42 VN.n10 B 0.784433f
C43 VN.n11 B 0.221007f
C44 VN.n12 B 0.017639f
C45 VN.n13 B 0.033039f
C46 VN.n14 B 0.033039f
C47 VN.n15 B 0.025861f
C48 VN.n16 B 0.017639f
C49 VN.n17 B 0.017639f
C50 VN.n18 B 0.017639f
C51 VN.n19 B 0.033039f
C52 VN.n20 B 0.033039f
C53 VN.t4 B 2.18798f
C54 VN.n21 B 0.765686f
C55 VN.n22 B 0.024556f
C56 VN.n23 B 0.017639f
C57 VN.n24 B 0.017639f
C58 VN.n25 B 0.017639f
C59 VN.n26 B 0.033039f
C60 VN.n27 B 0.033039f
C61 VN.n28 B 0.024871f
C62 VN.n29 B 0.017639f
C63 VN.n30 B 0.017639f
C64 VN.n31 B 0.017639f
C65 VN.n32 B 0.033039f
C66 VN.n33 B 0.033039f
C67 VN.n34 B 0.023904f
C68 VN.n35 B 0.028473f
C69 VN.n36 B 0.04817f
C70 VN.t1 B 2.18798f
C71 VN.n37 B 0.837757f
C72 VN.n38 B 0.017639f
C73 VN.n39 B 0.026851f
C74 VN.n40 B 0.017639f
C75 VN.n41 B 0.025209f
C76 VN.n42 B 0.017639f
C77 VN.t5 B 2.18798f
C78 VN.n43 B 0.765686f
C79 VN.n44 B 0.025861f
C80 VN.n45 B 0.017639f
C81 VN.n46 B 0.024556f
C82 VN.t7 B 2.44873f
C83 VN.t6 B 2.18798f
C84 VN.n47 B 0.827434f
C85 VN.n48 B 0.784433f
C86 VN.n49 B 0.221007f
C87 VN.n50 B 0.017639f
C88 VN.n51 B 0.033039f
C89 VN.n52 B 0.033039f
C90 VN.n53 B 0.025861f
C91 VN.n54 B 0.017639f
C92 VN.n55 B 0.017639f
C93 VN.n56 B 0.017639f
C94 VN.n57 B 0.033039f
C95 VN.n58 B 0.033039f
C96 VN.n59 B 0.024556f
C97 VN.n60 B 0.017639f
C98 VN.n61 B 0.017639f
C99 VN.n62 B 0.017639f
C100 VN.n63 B 0.033039f
C101 VN.n64 B 0.033039f
C102 VN.n65 B 0.024871f
C103 VN.n66 B 0.017639f
C104 VN.n67 B 0.017639f
C105 VN.n68 B 0.017639f
C106 VN.n69 B 0.033039f
C107 VN.n70 B 0.033039f
C108 VN.n71 B 0.023904f
C109 VN.n72 B 0.028473f
C110 VN.n73 B 1.19854f
C111 VTAIL.t6 B 0.201494f
C112 VTAIL.t5 B 0.201494f
C113 VTAIL.n0 B 1.73682f
C114 VTAIL.n1 B 0.434764f
C115 VTAIL.t7 B 2.2148f
C116 VTAIL.n2 B 0.533452f
C117 VTAIL.t12 B 2.2148f
C118 VTAIL.n3 B 0.533452f
C119 VTAIL.t11 B 0.201494f
C120 VTAIL.t14 B 0.201494f
C121 VTAIL.n4 B 1.73682f
C122 VTAIL.n5 B 0.657167f
C123 VTAIL.t8 B 2.2148f
C124 VTAIL.n6 B 1.71497f
C125 VTAIL.t2 B 2.21481f
C126 VTAIL.n7 B 1.71496f
C127 VTAIL.t1 B 0.201494f
C128 VTAIL.t4 B 0.201494f
C129 VTAIL.n8 B 1.73682f
C130 VTAIL.n9 B 0.657162f
C131 VTAIL.t0 B 2.21481f
C132 VTAIL.n10 B 0.533438f
C133 VTAIL.t10 B 2.21481f
C134 VTAIL.n11 B 0.533438f
C135 VTAIL.t13 B 0.201494f
C136 VTAIL.t15 B 0.201494f
C137 VTAIL.n12 B 1.73682f
C138 VTAIL.n13 B 0.657162f
C139 VTAIL.t9 B 2.2148f
C140 VTAIL.n14 B 1.71497f
C141 VTAIL.t3 B 2.2148f
C142 VTAIL.n15 B 1.71114f
C143 VDD1.t5 B 0.269925f
C144 VDD1.t2 B 0.269925f
C145 VDD1.n0 B 2.42949f
C146 VDD1.t6 B 0.269925f
C147 VDD1.t3 B 0.269925f
C148 VDD1.n1 B 2.42801f
C149 VDD1.t1 B 0.269925f
C150 VDD1.t7 B 0.269925f
C151 VDD1.n2 B 2.42801f
C152 VDD1.n3 B 4.35275f
C153 VDD1.t0 B 0.269925f
C154 VDD1.t4 B 0.269925f
C155 VDD1.n4 B 2.40985f
C156 VDD1.n5 B 3.70999f
C157 VP.t3 B 2.22788f
C158 VP.n0 B 0.853036f
C159 VP.n1 B 0.01796f
C160 VP.n2 B 0.027341f
C161 VP.n3 B 0.01796f
C162 VP.n4 B 0.025669f
C163 VP.n5 B 0.01796f
C164 VP.n6 B 0.026333f
C165 VP.n7 B 0.01796f
C166 VP.n8 B 0.025004f
C167 VP.n9 B 0.01796f
C168 VP.n10 B 0.025325f
C169 VP.n11 B 0.01796f
C170 VP.n12 B 0.02434f
C171 VP.t6 B 2.22788f
C172 VP.n13 B 0.853036f
C173 VP.n14 B 0.01796f
C174 VP.n15 B 0.027341f
C175 VP.n16 B 0.01796f
C176 VP.n17 B 0.025669f
C177 VP.n18 B 0.01796f
C178 VP.n19 B 0.026333f
C179 VP.n20 B 0.01796f
C180 VP.n21 B 0.025004f
C181 VP.t5 B 2.49339f
C182 VP.t2 B 2.22788f
C183 VP.n22 B 0.842524f
C184 VP.n23 B 0.798741f
C185 VP.n24 B 0.225038f
C186 VP.n25 B 0.01796f
C187 VP.n26 B 0.033641f
C188 VP.n27 B 0.033641f
C189 VP.n28 B 0.026333f
C190 VP.n29 B 0.01796f
C191 VP.n30 B 0.01796f
C192 VP.n31 B 0.01796f
C193 VP.n32 B 0.033641f
C194 VP.n33 B 0.033641f
C195 VP.t0 B 2.22788f
C196 VP.n34 B 0.77965f
C197 VP.n35 B 0.025004f
C198 VP.n36 B 0.01796f
C199 VP.n37 B 0.01796f
C200 VP.n38 B 0.01796f
C201 VP.n39 B 0.033641f
C202 VP.n40 B 0.033641f
C203 VP.n41 B 0.025325f
C204 VP.n42 B 0.01796f
C205 VP.n43 B 0.01796f
C206 VP.n44 B 0.01796f
C207 VP.n45 B 0.033641f
C208 VP.n46 B 0.033641f
C209 VP.n47 B 0.02434f
C210 VP.n48 B 0.028992f
C211 VP.n49 B 1.21334f
C212 VP.t7 B 2.22788f
C213 VP.n50 B 0.853036f
C214 VP.n51 B 1.22477f
C215 VP.n52 B 0.028992f
C216 VP.n53 B 0.01796f
C217 VP.n54 B 0.033641f
C218 VP.n55 B 0.033641f
C219 VP.n56 B 0.027341f
C220 VP.n57 B 0.01796f
C221 VP.n58 B 0.01796f
C222 VP.n59 B 0.01796f
C223 VP.n60 B 0.033641f
C224 VP.n61 B 0.033641f
C225 VP.t4 B 2.22788f
C226 VP.n62 B 0.77965f
C227 VP.n63 B 0.025669f
C228 VP.n64 B 0.01796f
C229 VP.n65 B 0.01796f
C230 VP.n66 B 0.01796f
C231 VP.n67 B 0.033641f
C232 VP.n68 B 0.033641f
C233 VP.n69 B 0.026333f
C234 VP.n70 B 0.01796f
C235 VP.n71 B 0.01796f
C236 VP.n72 B 0.01796f
C237 VP.n73 B 0.033641f
C238 VP.n74 B 0.033641f
C239 VP.t1 B 2.22788f
C240 VP.n75 B 0.77965f
C241 VP.n76 B 0.025004f
C242 VP.n77 B 0.01796f
C243 VP.n78 B 0.01796f
C244 VP.n79 B 0.01796f
C245 VP.n80 B 0.033641f
C246 VP.n81 B 0.033641f
C247 VP.n82 B 0.025325f
C248 VP.n83 B 0.01796f
C249 VP.n84 B 0.01796f
C250 VP.n85 B 0.01796f
C251 VP.n86 B 0.033641f
C252 VP.n87 B 0.033641f
C253 VP.n88 B 0.02434f
C254 VP.n89 B 0.028992f
C255 VP.n90 B 0.049048f
.ends

