* NGSPICE file created from diff_pair_sample_1059.ext - technology: sky130A

.subckt diff_pair_sample_1059 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0.4836 ps=3.26 w=1.24 l=2.91
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0 ps=0 w=1.24 l=2.91
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0 ps=0 w=1.24 l=2.91
X3 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0.4836 ps=3.26 w=1.24 l=2.91
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0.4836 ps=3.26 w=1.24 l=2.91
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0 ps=0 w=1.24 l=2.91
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0 ps=0 w=1.24 l=2.91
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4836 pd=3.26 as=0.4836 ps=3.26 w=1.24 l=2.91
R0 VP.n0 VP.t1 88.7351
R1 VP.n0 VP.t0 51.4077
R2 VP VP.n0 0.431812
R3 VTAIL.n3 VTAIL.t0 155.132
R4 VTAIL.n0 VTAIL.t2 155.132
R5 VTAIL.n2 VTAIL.t3 155.132
R6 VTAIL.n1 VTAIL.t1 155.132
R7 VTAIL.n1 VTAIL.n0 19.0221
R8 VTAIL.n3 VTAIL.n2 16.2289
R9 VTAIL.n2 VTAIL.n1 1.86688
R10 VTAIL VTAIL.n0 1.22679
R11 VTAIL VTAIL.n3 0.640586
R12 VDD1 VDD1.t1 203.349
R13 VDD1 VDD1.t0 172.567
R14 B.n372 B.n371 585
R15 B.n373 B.n372 585
R16 B.n125 B.n67 585
R17 B.n124 B.n123 585
R18 B.n122 B.n121 585
R19 B.n120 B.n119 585
R20 B.n118 B.n117 585
R21 B.n116 B.n115 585
R22 B.n114 B.n113 585
R23 B.n112 B.n111 585
R24 B.n110 B.n109 585
R25 B.n107 B.n106 585
R26 B.n105 B.n104 585
R27 B.n103 B.n102 585
R28 B.n101 B.n100 585
R29 B.n99 B.n98 585
R30 B.n97 B.n96 585
R31 B.n95 B.n94 585
R32 B.n93 B.n92 585
R33 B.n91 B.n90 585
R34 B.n89 B.n88 585
R35 B.n87 B.n86 585
R36 B.n85 B.n84 585
R37 B.n83 B.n82 585
R38 B.n81 B.n80 585
R39 B.n79 B.n78 585
R40 B.n77 B.n76 585
R41 B.n75 B.n74 585
R42 B.n53 B.n52 585
R43 B.n376 B.n375 585
R44 B.n370 B.n68 585
R45 B.n68 B.n50 585
R46 B.n369 B.n49 585
R47 B.n380 B.n49 585
R48 B.n368 B.n48 585
R49 B.n381 B.n48 585
R50 B.n367 B.n47 585
R51 B.n382 B.n47 585
R52 B.n366 B.n365 585
R53 B.n365 B.n43 585
R54 B.n364 B.n42 585
R55 B.n388 B.n42 585
R56 B.n363 B.n41 585
R57 B.n389 B.n41 585
R58 B.n362 B.n40 585
R59 B.n390 B.n40 585
R60 B.n361 B.n360 585
R61 B.n360 B.n36 585
R62 B.n359 B.n35 585
R63 B.n396 B.n35 585
R64 B.n358 B.n34 585
R65 B.n397 B.n34 585
R66 B.n357 B.n33 585
R67 B.n398 B.n33 585
R68 B.n356 B.n355 585
R69 B.n355 B.n29 585
R70 B.n354 B.n28 585
R71 B.n404 B.n28 585
R72 B.n353 B.n27 585
R73 B.n405 B.n27 585
R74 B.n352 B.n26 585
R75 B.n406 B.n26 585
R76 B.n351 B.n350 585
R77 B.n350 B.n22 585
R78 B.n349 B.n21 585
R79 B.n412 B.n21 585
R80 B.n348 B.n20 585
R81 B.n413 B.n20 585
R82 B.n347 B.n19 585
R83 B.n414 B.n19 585
R84 B.n346 B.n345 585
R85 B.n345 B.n18 585
R86 B.n344 B.n14 585
R87 B.n420 B.n14 585
R88 B.n343 B.n13 585
R89 B.n421 B.n13 585
R90 B.n342 B.n12 585
R91 B.n422 B.n12 585
R92 B.n341 B.n340 585
R93 B.n340 B.n8 585
R94 B.n339 B.n7 585
R95 B.n428 B.n7 585
R96 B.n338 B.n6 585
R97 B.n429 B.n6 585
R98 B.n337 B.n5 585
R99 B.n430 B.n5 585
R100 B.n336 B.n335 585
R101 B.n335 B.n4 585
R102 B.n334 B.n126 585
R103 B.n334 B.n333 585
R104 B.n324 B.n127 585
R105 B.n128 B.n127 585
R106 B.n326 B.n325 585
R107 B.n327 B.n326 585
R108 B.n323 B.n133 585
R109 B.n133 B.n132 585
R110 B.n322 B.n321 585
R111 B.n321 B.n320 585
R112 B.n135 B.n134 585
R113 B.n313 B.n135 585
R114 B.n312 B.n311 585
R115 B.n314 B.n312 585
R116 B.n310 B.n140 585
R117 B.n140 B.n139 585
R118 B.n309 B.n308 585
R119 B.n308 B.n307 585
R120 B.n142 B.n141 585
R121 B.n143 B.n142 585
R122 B.n300 B.n299 585
R123 B.n301 B.n300 585
R124 B.n298 B.n148 585
R125 B.n148 B.n147 585
R126 B.n297 B.n296 585
R127 B.n296 B.n295 585
R128 B.n150 B.n149 585
R129 B.n151 B.n150 585
R130 B.n288 B.n287 585
R131 B.n289 B.n288 585
R132 B.n286 B.n156 585
R133 B.n156 B.n155 585
R134 B.n285 B.n284 585
R135 B.n284 B.n283 585
R136 B.n158 B.n157 585
R137 B.n159 B.n158 585
R138 B.n276 B.n275 585
R139 B.n277 B.n276 585
R140 B.n274 B.n164 585
R141 B.n164 B.n163 585
R142 B.n273 B.n272 585
R143 B.n272 B.n271 585
R144 B.n166 B.n165 585
R145 B.n167 B.n166 585
R146 B.n264 B.n263 585
R147 B.n265 B.n264 585
R148 B.n262 B.n172 585
R149 B.n172 B.n171 585
R150 B.n261 B.n260 585
R151 B.n260 B.n259 585
R152 B.n174 B.n173 585
R153 B.n175 B.n174 585
R154 B.n255 B.n254 585
R155 B.n178 B.n177 585
R156 B.n251 B.n250 585
R157 B.n252 B.n251 585
R158 B.n249 B.n192 585
R159 B.n248 B.n247 585
R160 B.n246 B.n245 585
R161 B.n244 B.n243 585
R162 B.n242 B.n241 585
R163 B.n240 B.n239 585
R164 B.n238 B.n237 585
R165 B.n235 B.n234 585
R166 B.n233 B.n232 585
R167 B.n231 B.n230 585
R168 B.n229 B.n228 585
R169 B.n227 B.n226 585
R170 B.n225 B.n224 585
R171 B.n223 B.n222 585
R172 B.n221 B.n220 585
R173 B.n219 B.n218 585
R174 B.n217 B.n216 585
R175 B.n215 B.n214 585
R176 B.n213 B.n212 585
R177 B.n211 B.n210 585
R178 B.n209 B.n208 585
R179 B.n207 B.n206 585
R180 B.n205 B.n204 585
R181 B.n203 B.n202 585
R182 B.n201 B.n200 585
R183 B.n199 B.n198 585
R184 B.n256 B.n176 585
R185 B.n176 B.n175 585
R186 B.n258 B.n257 585
R187 B.n259 B.n258 585
R188 B.n170 B.n169 585
R189 B.n171 B.n170 585
R190 B.n267 B.n266 585
R191 B.n266 B.n265 585
R192 B.n268 B.n168 585
R193 B.n168 B.n167 585
R194 B.n270 B.n269 585
R195 B.n271 B.n270 585
R196 B.n162 B.n161 585
R197 B.n163 B.n162 585
R198 B.n279 B.n278 585
R199 B.n278 B.n277 585
R200 B.n280 B.n160 585
R201 B.n160 B.n159 585
R202 B.n282 B.n281 585
R203 B.n283 B.n282 585
R204 B.n154 B.n153 585
R205 B.n155 B.n154 585
R206 B.n291 B.n290 585
R207 B.n290 B.n289 585
R208 B.n292 B.n152 585
R209 B.n152 B.n151 585
R210 B.n294 B.n293 585
R211 B.n295 B.n294 585
R212 B.n146 B.n145 585
R213 B.n147 B.n146 585
R214 B.n303 B.n302 585
R215 B.n302 B.n301 585
R216 B.n304 B.n144 585
R217 B.n144 B.n143 585
R218 B.n306 B.n305 585
R219 B.n307 B.n306 585
R220 B.n138 B.n137 585
R221 B.n139 B.n138 585
R222 B.n316 B.n315 585
R223 B.n315 B.n314 585
R224 B.n317 B.n136 585
R225 B.n313 B.n136 585
R226 B.n319 B.n318 585
R227 B.n320 B.n319 585
R228 B.n131 B.n130 585
R229 B.n132 B.n131 585
R230 B.n329 B.n328 585
R231 B.n328 B.n327 585
R232 B.n330 B.n129 585
R233 B.n129 B.n128 585
R234 B.n332 B.n331 585
R235 B.n333 B.n332 585
R236 B.n2 B.n0 585
R237 B.n4 B.n2 585
R238 B.n3 B.n1 585
R239 B.n429 B.n3 585
R240 B.n427 B.n426 585
R241 B.n428 B.n427 585
R242 B.n425 B.n9 585
R243 B.n9 B.n8 585
R244 B.n424 B.n423 585
R245 B.n423 B.n422 585
R246 B.n11 B.n10 585
R247 B.n421 B.n11 585
R248 B.n419 B.n418 585
R249 B.n420 B.n419 585
R250 B.n417 B.n15 585
R251 B.n18 B.n15 585
R252 B.n416 B.n415 585
R253 B.n415 B.n414 585
R254 B.n17 B.n16 585
R255 B.n413 B.n17 585
R256 B.n411 B.n410 585
R257 B.n412 B.n411 585
R258 B.n409 B.n23 585
R259 B.n23 B.n22 585
R260 B.n408 B.n407 585
R261 B.n407 B.n406 585
R262 B.n25 B.n24 585
R263 B.n405 B.n25 585
R264 B.n403 B.n402 585
R265 B.n404 B.n403 585
R266 B.n401 B.n30 585
R267 B.n30 B.n29 585
R268 B.n400 B.n399 585
R269 B.n399 B.n398 585
R270 B.n32 B.n31 585
R271 B.n397 B.n32 585
R272 B.n395 B.n394 585
R273 B.n396 B.n395 585
R274 B.n393 B.n37 585
R275 B.n37 B.n36 585
R276 B.n392 B.n391 585
R277 B.n391 B.n390 585
R278 B.n39 B.n38 585
R279 B.n389 B.n39 585
R280 B.n387 B.n386 585
R281 B.n388 B.n387 585
R282 B.n385 B.n44 585
R283 B.n44 B.n43 585
R284 B.n384 B.n383 585
R285 B.n383 B.n382 585
R286 B.n46 B.n45 585
R287 B.n381 B.n46 585
R288 B.n379 B.n378 585
R289 B.n380 B.n379 585
R290 B.n377 B.n51 585
R291 B.n51 B.n50 585
R292 B.n432 B.n431 585
R293 B.n431 B.n430 585
R294 B.n254 B.n176 569.379
R295 B.n375 B.n51 569.379
R296 B.n198 B.n174 569.379
R297 B.n372 B.n68 569.379
R298 B.n373 B.n66 256.663
R299 B.n373 B.n65 256.663
R300 B.n373 B.n64 256.663
R301 B.n373 B.n63 256.663
R302 B.n373 B.n62 256.663
R303 B.n373 B.n61 256.663
R304 B.n373 B.n60 256.663
R305 B.n373 B.n59 256.663
R306 B.n373 B.n58 256.663
R307 B.n373 B.n57 256.663
R308 B.n373 B.n56 256.663
R309 B.n373 B.n55 256.663
R310 B.n373 B.n54 256.663
R311 B.n374 B.n373 256.663
R312 B.n253 B.n252 256.663
R313 B.n252 B.n179 256.663
R314 B.n252 B.n180 256.663
R315 B.n252 B.n181 256.663
R316 B.n252 B.n182 256.663
R317 B.n252 B.n183 256.663
R318 B.n252 B.n184 256.663
R319 B.n252 B.n185 256.663
R320 B.n252 B.n186 256.663
R321 B.n252 B.n187 256.663
R322 B.n252 B.n188 256.663
R323 B.n252 B.n189 256.663
R324 B.n252 B.n190 256.663
R325 B.n252 B.n191 256.663
R326 B.n252 B.n175 227.936
R327 B.n373 B.n50 227.936
R328 B.n195 B.t12 211.851
R329 B.n193 B.t15 211.851
R330 B.n71 B.t7 211.851
R331 B.n69 B.t4 211.851
R332 B.n195 B.t9 209.149
R333 B.n193 B.t13 209.149
R334 B.n71 B.t6 209.149
R335 B.n69 B.t2 209.149
R336 B.n258 B.n176 163.367
R337 B.n258 B.n170 163.367
R338 B.n266 B.n170 163.367
R339 B.n266 B.n168 163.367
R340 B.n270 B.n168 163.367
R341 B.n270 B.n162 163.367
R342 B.n278 B.n162 163.367
R343 B.n278 B.n160 163.367
R344 B.n282 B.n160 163.367
R345 B.n282 B.n154 163.367
R346 B.n290 B.n154 163.367
R347 B.n290 B.n152 163.367
R348 B.n294 B.n152 163.367
R349 B.n294 B.n146 163.367
R350 B.n302 B.n146 163.367
R351 B.n302 B.n144 163.367
R352 B.n306 B.n144 163.367
R353 B.n306 B.n138 163.367
R354 B.n315 B.n138 163.367
R355 B.n315 B.n136 163.367
R356 B.n319 B.n136 163.367
R357 B.n319 B.n131 163.367
R358 B.n328 B.n131 163.367
R359 B.n328 B.n129 163.367
R360 B.n332 B.n129 163.367
R361 B.n332 B.n2 163.367
R362 B.n431 B.n2 163.367
R363 B.n431 B.n3 163.367
R364 B.n427 B.n3 163.367
R365 B.n427 B.n9 163.367
R366 B.n423 B.n9 163.367
R367 B.n423 B.n11 163.367
R368 B.n419 B.n11 163.367
R369 B.n419 B.n15 163.367
R370 B.n415 B.n15 163.367
R371 B.n415 B.n17 163.367
R372 B.n411 B.n17 163.367
R373 B.n411 B.n23 163.367
R374 B.n407 B.n23 163.367
R375 B.n407 B.n25 163.367
R376 B.n403 B.n25 163.367
R377 B.n403 B.n30 163.367
R378 B.n399 B.n30 163.367
R379 B.n399 B.n32 163.367
R380 B.n395 B.n32 163.367
R381 B.n395 B.n37 163.367
R382 B.n391 B.n37 163.367
R383 B.n391 B.n39 163.367
R384 B.n387 B.n39 163.367
R385 B.n387 B.n44 163.367
R386 B.n383 B.n44 163.367
R387 B.n383 B.n46 163.367
R388 B.n379 B.n46 163.367
R389 B.n379 B.n51 163.367
R390 B.n251 B.n178 163.367
R391 B.n251 B.n192 163.367
R392 B.n247 B.n246 163.367
R393 B.n243 B.n242 163.367
R394 B.n239 B.n238 163.367
R395 B.n234 B.n233 163.367
R396 B.n230 B.n229 163.367
R397 B.n226 B.n225 163.367
R398 B.n222 B.n221 163.367
R399 B.n218 B.n217 163.367
R400 B.n214 B.n213 163.367
R401 B.n210 B.n209 163.367
R402 B.n206 B.n205 163.367
R403 B.n202 B.n201 163.367
R404 B.n260 B.n174 163.367
R405 B.n260 B.n172 163.367
R406 B.n264 B.n172 163.367
R407 B.n264 B.n166 163.367
R408 B.n272 B.n166 163.367
R409 B.n272 B.n164 163.367
R410 B.n276 B.n164 163.367
R411 B.n276 B.n158 163.367
R412 B.n284 B.n158 163.367
R413 B.n284 B.n156 163.367
R414 B.n288 B.n156 163.367
R415 B.n288 B.n150 163.367
R416 B.n296 B.n150 163.367
R417 B.n296 B.n148 163.367
R418 B.n300 B.n148 163.367
R419 B.n300 B.n142 163.367
R420 B.n308 B.n142 163.367
R421 B.n308 B.n140 163.367
R422 B.n312 B.n140 163.367
R423 B.n312 B.n135 163.367
R424 B.n321 B.n135 163.367
R425 B.n321 B.n133 163.367
R426 B.n326 B.n133 163.367
R427 B.n326 B.n127 163.367
R428 B.n334 B.n127 163.367
R429 B.n335 B.n334 163.367
R430 B.n335 B.n5 163.367
R431 B.n6 B.n5 163.367
R432 B.n7 B.n6 163.367
R433 B.n340 B.n7 163.367
R434 B.n340 B.n12 163.367
R435 B.n13 B.n12 163.367
R436 B.n14 B.n13 163.367
R437 B.n345 B.n14 163.367
R438 B.n345 B.n19 163.367
R439 B.n20 B.n19 163.367
R440 B.n21 B.n20 163.367
R441 B.n350 B.n21 163.367
R442 B.n350 B.n26 163.367
R443 B.n27 B.n26 163.367
R444 B.n28 B.n27 163.367
R445 B.n355 B.n28 163.367
R446 B.n355 B.n33 163.367
R447 B.n34 B.n33 163.367
R448 B.n35 B.n34 163.367
R449 B.n360 B.n35 163.367
R450 B.n360 B.n40 163.367
R451 B.n41 B.n40 163.367
R452 B.n42 B.n41 163.367
R453 B.n365 B.n42 163.367
R454 B.n365 B.n47 163.367
R455 B.n48 B.n47 163.367
R456 B.n49 B.n48 163.367
R457 B.n68 B.n49 163.367
R458 B.n74 B.n53 163.367
R459 B.n78 B.n77 163.367
R460 B.n82 B.n81 163.367
R461 B.n86 B.n85 163.367
R462 B.n90 B.n89 163.367
R463 B.n94 B.n93 163.367
R464 B.n98 B.n97 163.367
R465 B.n102 B.n101 163.367
R466 B.n106 B.n105 163.367
R467 B.n111 B.n110 163.367
R468 B.n115 B.n114 163.367
R469 B.n119 B.n118 163.367
R470 B.n123 B.n122 163.367
R471 B.n372 B.n67 163.367
R472 B.n196 B.t11 149.014
R473 B.n194 B.t14 149.014
R474 B.n72 B.t8 149.014
R475 B.n70 B.t5 149.014
R476 B.n259 B.n175 114.812
R477 B.n259 B.n171 114.812
R478 B.n265 B.n171 114.812
R479 B.n265 B.n167 114.812
R480 B.n271 B.n167 114.812
R481 B.n271 B.n163 114.812
R482 B.n277 B.n163 114.812
R483 B.n283 B.n159 114.812
R484 B.n283 B.n155 114.812
R485 B.n289 B.n155 114.812
R486 B.n289 B.n151 114.812
R487 B.n295 B.n151 114.812
R488 B.n295 B.n147 114.812
R489 B.n301 B.n147 114.812
R490 B.n301 B.n143 114.812
R491 B.n307 B.n143 114.812
R492 B.n307 B.n139 114.812
R493 B.n314 B.n139 114.812
R494 B.n314 B.n313 114.812
R495 B.n320 B.n132 114.812
R496 B.n327 B.n132 114.812
R497 B.n327 B.n128 114.812
R498 B.n333 B.n128 114.812
R499 B.n333 B.n4 114.812
R500 B.n430 B.n4 114.812
R501 B.n430 B.n429 114.812
R502 B.n429 B.n428 114.812
R503 B.n428 B.n8 114.812
R504 B.n422 B.n8 114.812
R505 B.n422 B.n421 114.812
R506 B.n421 B.n420 114.812
R507 B.n414 B.n18 114.812
R508 B.n414 B.n413 114.812
R509 B.n413 B.n412 114.812
R510 B.n412 B.n22 114.812
R511 B.n406 B.n22 114.812
R512 B.n406 B.n405 114.812
R513 B.n405 B.n404 114.812
R514 B.n404 B.n29 114.812
R515 B.n398 B.n29 114.812
R516 B.n398 B.n397 114.812
R517 B.n397 B.n396 114.812
R518 B.n396 B.n36 114.812
R519 B.n390 B.n389 114.812
R520 B.n389 B.n388 114.812
R521 B.n388 B.n43 114.812
R522 B.n382 B.n43 114.812
R523 B.n382 B.n381 114.812
R524 B.n381 B.n380 114.812
R525 B.n380 B.n50 114.812
R526 B.n277 B.t10 102.993
R527 B.n390 B.t3 102.993
R528 B.n313 B.t1 72.6022
R529 B.n18 B.t0 72.6022
R530 B.n254 B.n253 71.676
R531 B.n192 B.n179 71.676
R532 B.n246 B.n180 71.676
R533 B.n242 B.n181 71.676
R534 B.n238 B.n182 71.676
R535 B.n233 B.n183 71.676
R536 B.n229 B.n184 71.676
R537 B.n225 B.n185 71.676
R538 B.n221 B.n186 71.676
R539 B.n217 B.n187 71.676
R540 B.n213 B.n188 71.676
R541 B.n209 B.n189 71.676
R542 B.n205 B.n190 71.676
R543 B.n201 B.n191 71.676
R544 B.n375 B.n374 71.676
R545 B.n74 B.n54 71.676
R546 B.n78 B.n55 71.676
R547 B.n82 B.n56 71.676
R548 B.n86 B.n57 71.676
R549 B.n90 B.n58 71.676
R550 B.n94 B.n59 71.676
R551 B.n98 B.n60 71.676
R552 B.n102 B.n61 71.676
R553 B.n106 B.n62 71.676
R554 B.n111 B.n63 71.676
R555 B.n115 B.n64 71.676
R556 B.n119 B.n65 71.676
R557 B.n123 B.n66 71.676
R558 B.n67 B.n66 71.676
R559 B.n122 B.n65 71.676
R560 B.n118 B.n64 71.676
R561 B.n114 B.n63 71.676
R562 B.n110 B.n62 71.676
R563 B.n105 B.n61 71.676
R564 B.n101 B.n60 71.676
R565 B.n97 B.n59 71.676
R566 B.n93 B.n58 71.676
R567 B.n89 B.n57 71.676
R568 B.n85 B.n56 71.676
R569 B.n81 B.n55 71.676
R570 B.n77 B.n54 71.676
R571 B.n374 B.n53 71.676
R572 B.n253 B.n178 71.676
R573 B.n247 B.n179 71.676
R574 B.n243 B.n180 71.676
R575 B.n239 B.n181 71.676
R576 B.n234 B.n182 71.676
R577 B.n230 B.n183 71.676
R578 B.n226 B.n184 71.676
R579 B.n222 B.n185 71.676
R580 B.n218 B.n186 71.676
R581 B.n214 B.n187 71.676
R582 B.n210 B.n188 71.676
R583 B.n206 B.n189 71.676
R584 B.n202 B.n190 71.676
R585 B.n198 B.n191 71.676
R586 B.n196 B.n195 62.8369
R587 B.n194 B.n193 62.8369
R588 B.n72 B.n71 62.8369
R589 B.n70 B.n69 62.8369
R590 B.n197 B.n196 59.5399
R591 B.n236 B.n194 59.5399
R592 B.n73 B.n72 59.5399
R593 B.n108 B.n70 59.5399
R594 B.n320 B.t1 42.2108
R595 B.n420 B.t0 42.2108
R596 B.n377 B.n376 36.9956
R597 B.n371 B.n370 36.9956
R598 B.n199 B.n173 36.9956
R599 B.n256 B.n255 36.9956
R600 B B.n432 18.0485
R601 B.t10 B.n159 11.8194
R602 B.t3 B.n36 11.8194
R603 B.n376 B.n52 10.6151
R604 B.n75 B.n52 10.6151
R605 B.n76 B.n75 10.6151
R606 B.n79 B.n76 10.6151
R607 B.n80 B.n79 10.6151
R608 B.n83 B.n80 10.6151
R609 B.n84 B.n83 10.6151
R610 B.n87 B.n84 10.6151
R611 B.n88 B.n87 10.6151
R612 B.n92 B.n91 10.6151
R613 B.n95 B.n92 10.6151
R614 B.n96 B.n95 10.6151
R615 B.n99 B.n96 10.6151
R616 B.n100 B.n99 10.6151
R617 B.n103 B.n100 10.6151
R618 B.n104 B.n103 10.6151
R619 B.n107 B.n104 10.6151
R620 B.n112 B.n109 10.6151
R621 B.n113 B.n112 10.6151
R622 B.n116 B.n113 10.6151
R623 B.n117 B.n116 10.6151
R624 B.n120 B.n117 10.6151
R625 B.n121 B.n120 10.6151
R626 B.n124 B.n121 10.6151
R627 B.n125 B.n124 10.6151
R628 B.n371 B.n125 10.6151
R629 B.n261 B.n173 10.6151
R630 B.n262 B.n261 10.6151
R631 B.n263 B.n262 10.6151
R632 B.n263 B.n165 10.6151
R633 B.n273 B.n165 10.6151
R634 B.n274 B.n273 10.6151
R635 B.n275 B.n274 10.6151
R636 B.n275 B.n157 10.6151
R637 B.n285 B.n157 10.6151
R638 B.n286 B.n285 10.6151
R639 B.n287 B.n286 10.6151
R640 B.n287 B.n149 10.6151
R641 B.n297 B.n149 10.6151
R642 B.n298 B.n297 10.6151
R643 B.n299 B.n298 10.6151
R644 B.n299 B.n141 10.6151
R645 B.n309 B.n141 10.6151
R646 B.n310 B.n309 10.6151
R647 B.n311 B.n310 10.6151
R648 B.n311 B.n134 10.6151
R649 B.n322 B.n134 10.6151
R650 B.n323 B.n322 10.6151
R651 B.n325 B.n323 10.6151
R652 B.n325 B.n324 10.6151
R653 B.n324 B.n126 10.6151
R654 B.n336 B.n126 10.6151
R655 B.n337 B.n336 10.6151
R656 B.n338 B.n337 10.6151
R657 B.n339 B.n338 10.6151
R658 B.n341 B.n339 10.6151
R659 B.n342 B.n341 10.6151
R660 B.n343 B.n342 10.6151
R661 B.n344 B.n343 10.6151
R662 B.n346 B.n344 10.6151
R663 B.n347 B.n346 10.6151
R664 B.n348 B.n347 10.6151
R665 B.n349 B.n348 10.6151
R666 B.n351 B.n349 10.6151
R667 B.n352 B.n351 10.6151
R668 B.n353 B.n352 10.6151
R669 B.n354 B.n353 10.6151
R670 B.n356 B.n354 10.6151
R671 B.n357 B.n356 10.6151
R672 B.n358 B.n357 10.6151
R673 B.n359 B.n358 10.6151
R674 B.n361 B.n359 10.6151
R675 B.n362 B.n361 10.6151
R676 B.n363 B.n362 10.6151
R677 B.n364 B.n363 10.6151
R678 B.n366 B.n364 10.6151
R679 B.n367 B.n366 10.6151
R680 B.n368 B.n367 10.6151
R681 B.n369 B.n368 10.6151
R682 B.n370 B.n369 10.6151
R683 B.n255 B.n177 10.6151
R684 B.n250 B.n177 10.6151
R685 B.n250 B.n249 10.6151
R686 B.n249 B.n248 10.6151
R687 B.n248 B.n245 10.6151
R688 B.n245 B.n244 10.6151
R689 B.n244 B.n241 10.6151
R690 B.n241 B.n240 10.6151
R691 B.n240 B.n237 10.6151
R692 B.n235 B.n232 10.6151
R693 B.n232 B.n231 10.6151
R694 B.n231 B.n228 10.6151
R695 B.n228 B.n227 10.6151
R696 B.n227 B.n224 10.6151
R697 B.n224 B.n223 10.6151
R698 B.n223 B.n220 10.6151
R699 B.n220 B.n219 10.6151
R700 B.n216 B.n215 10.6151
R701 B.n215 B.n212 10.6151
R702 B.n212 B.n211 10.6151
R703 B.n211 B.n208 10.6151
R704 B.n208 B.n207 10.6151
R705 B.n207 B.n204 10.6151
R706 B.n204 B.n203 10.6151
R707 B.n203 B.n200 10.6151
R708 B.n200 B.n199 10.6151
R709 B.n257 B.n256 10.6151
R710 B.n257 B.n169 10.6151
R711 B.n267 B.n169 10.6151
R712 B.n268 B.n267 10.6151
R713 B.n269 B.n268 10.6151
R714 B.n269 B.n161 10.6151
R715 B.n279 B.n161 10.6151
R716 B.n280 B.n279 10.6151
R717 B.n281 B.n280 10.6151
R718 B.n281 B.n153 10.6151
R719 B.n291 B.n153 10.6151
R720 B.n292 B.n291 10.6151
R721 B.n293 B.n292 10.6151
R722 B.n293 B.n145 10.6151
R723 B.n303 B.n145 10.6151
R724 B.n304 B.n303 10.6151
R725 B.n305 B.n304 10.6151
R726 B.n305 B.n137 10.6151
R727 B.n316 B.n137 10.6151
R728 B.n317 B.n316 10.6151
R729 B.n318 B.n317 10.6151
R730 B.n318 B.n130 10.6151
R731 B.n329 B.n130 10.6151
R732 B.n330 B.n329 10.6151
R733 B.n331 B.n330 10.6151
R734 B.n331 B.n0 10.6151
R735 B.n426 B.n1 10.6151
R736 B.n426 B.n425 10.6151
R737 B.n425 B.n424 10.6151
R738 B.n424 B.n10 10.6151
R739 B.n418 B.n10 10.6151
R740 B.n418 B.n417 10.6151
R741 B.n417 B.n416 10.6151
R742 B.n416 B.n16 10.6151
R743 B.n410 B.n16 10.6151
R744 B.n410 B.n409 10.6151
R745 B.n409 B.n408 10.6151
R746 B.n408 B.n24 10.6151
R747 B.n402 B.n24 10.6151
R748 B.n402 B.n401 10.6151
R749 B.n401 B.n400 10.6151
R750 B.n400 B.n31 10.6151
R751 B.n394 B.n31 10.6151
R752 B.n394 B.n393 10.6151
R753 B.n393 B.n392 10.6151
R754 B.n392 B.n38 10.6151
R755 B.n386 B.n38 10.6151
R756 B.n386 B.n385 10.6151
R757 B.n385 B.n384 10.6151
R758 B.n384 B.n45 10.6151
R759 B.n378 B.n45 10.6151
R760 B.n378 B.n377 10.6151
R761 B.n91 B.n73 6.5566
R762 B.n108 B.n107 6.5566
R763 B.n236 B.n235 6.5566
R764 B.n219 B.n197 6.5566
R765 B.n88 B.n73 4.05904
R766 B.n109 B.n108 4.05904
R767 B.n237 B.n236 4.05904
R768 B.n216 B.n197 4.05904
R769 B.n432 B.n0 2.81026
R770 B.n432 B.n1 2.81026
R771 VN VN.t0 88.7367
R772 VN VN.t1 51.839
R773 VDD2.n0 VDD2.t0 202.125
R774 VDD2.n0 VDD2.t1 171.811
R775 VDD2 VDD2.n0 0.756965
C0 VN VDD2 0.524266f
C1 VDD1 VP 0.720548f
C2 VDD1 VTAIL 2.32559f
C3 VDD1 VN 0.156008f
C4 VP VTAIL 0.958055f
C5 VDD1 VDD2 0.711054f
C6 VN VP 3.6137f
C7 VN VTAIL 0.943932f
C8 VP VDD2 0.354115f
C9 VDD2 VTAIL 2.38082f
C10 VDD2 B 2.578298f
C11 VDD1 B 4.59558f
C12 VTAIL B 2.701302f
C13 VN B 7.915061f
C14 VP B 5.806601f
C15 VDD2.t0 B 0.249803f
C16 VDD2.t1 B 0.124346f
C17 VDD2.n0 B 1.8929f
C18 VN.t1 B 0.508324f
C19 VN.t0 B 1.03926f
C20 VDD1.t0 B 0.116611f
C21 VDD1.t1 B 0.245453f
C22 VTAIL.t2 B 0.134037f
C23 VTAIL.n0 B 1.09856f
C24 VTAIL.t1 B 0.134037f
C25 VTAIL.n1 B 1.1473f
C26 VTAIL.t3 B 0.134037f
C27 VTAIL.n2 B 0.934626f
C28 VTAIL.t0 B 0.134037f
C29 VTAIL.n3 B 0.841252f
C30 VP.t0 B 0.512511f
C31 VP.t1 B 1.04788f
C32 VP.n0 B 1.95106f
.ends

