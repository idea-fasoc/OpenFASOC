* NGSPICE file created from diff_pair_sample_0538.ext - technology: sky130A

.subckt diff_pair_sample_0538 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=1.52
X1 B.t11 B.t9 B.t10 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=1.52
X2 B.t8 B.t6 B.t7 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=1.52
X3 VTAIL.t1 VP.t0 VDD1.t3 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=1.52
X4 B.t5 B.t3 B.t4 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=1.52
X5 VTAIL.t6 VN.t1 VDD2.t0 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=1.52
X6 VDD2.t3 VN.t2 VTAIL.t5 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=1.52
X7 VDD1.t2 VP.t1 VTAIL.t2 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=1.52
X8 VDD1.t1 VP.t2 VTAIL.t3 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=1.52
X9 B.t2 B.t0 B.t1 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=1.52
X10 VDD2.t1 VN.t3 VTAIL.t4 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=1.52
X11 VTAIL.t0 VP.t3 VDD1.t0 w_n2080_n1940# sky130_fd_pr__pfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=1.52
R0 VN.n0 VN.t1 113.791
R1 VN.n1 VN.t2 113.791
R2 VN.n0 VN.t3 113.472
R3 VN.n1 VN.t0 113.472
R4 VN VN.n1 50.8393
R5 VN VN.n0 12.9719
R6 VDD2.n2 VDD2.n0 131.965
R7 VDD2.n2 VDD2.n1 99.277
R8 VDD2.n1 VDD2.t2 6.68877
R9 VDD2.n1 VDD2.t3 6.68877
R10 VDD2.n0 VDD2.t0 6.68877
R11 VDD2.n0 VDD2.t1 6.68877
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t1 89.2866
R14 VTAIL.n4 VTAIL.t5 89.2866
R15 VTAIL.n3 VTAIL.t7 89.2866
R16 VTAIL.n7 VTAIL.t4 89.2865
R17 VTAIL.n0 VTAIL.t6 89.2865
R18 VTAIL.n1 VTAIL.t2 89.2865
R19 VTAIL.n2 VTAIL.t0 89.2865
R20 VTAIL.n6 VTAIL.t3 89.2865
R21 VTAIL.n7 VTAIL.n6 18.1514
R22 VTAIL.n3 VTAIL.n2 18.1514
R23 VTAIL.n4 VTAIL.n3 1.59533
R24 VTAIL.n6 VTAIL.n5 1.59533
R25 VTAIL.n2 VTAIL.n1 1.59533
R26 VTAIL VTAIL.n0 0.856103
R27 VTAIL VTAIL.n7 0.739724
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n223 B.n222 585
R31 B.n221 B.n70 585
R32 B.n220 B.n219 585
R33 B.n218 B.n71 585
R34 B.n217 B.n216 585
R35 B.n215 B.n72 585
R36 B.n214 B.n213 585
R37 B.n212 B.n73 585
R38 B.n211 B.n210 585
R39 B.n209 B.n74 585
R40 B.n208 B.n207 585
R41 B.n206 B.n75 585
R42 B.n205 B.n204 585
R43 B.n203 B.n76 585
R44 B.n202 B.n201 585
R45 B.n200 B.n77 585
R46 B.n199 B.n198 585
R47 B.n197 B.n78 585
R48 B.n196 B.n195 585
R49 B.n194 B.n79 585
R50 B.n193 B.n192 585
R51 B.n190 B.n80 585
R52 B.n189 B.n188 585
R53 B.n187 B.n83 585
R54 B.n186 B.n185 585
R55 B.n184 B.n84 585
R56 B.n183 B.n182 585
R57 B.n181 B.n85 585
R58 B.n180 B.n179 585
R59 B.n178 B.n86 585
R60 B.n176 B.n175 585
R61 B.n174 B.n89 585
R62 B.n173 B.n172 585
R63 B.n171 B.n90 585
R64 B.n170 B.n169 585
R65 B.n168 B.n91 585
R66 B.n167 B.n166 585
R67 B.n165 B.n92 585
R68 B.n164 B.n163 585
R69 B.n162 B.n93 585
R70 B.n161 B.n160 585
R71 B.n159 B.n94 585
R72 B.n158 B.n157 585
R73 B.n156 B.n95 585
R74 B.n155 B.n154 585
R75 B.n153 B.n96 585
R76 B.n152 B.n151 585
R77 B.n150 B.n97 585
R78 B.n149 B.n148 585
R79 B.n147 B.n98 585
R80 B.n146 B.n145 585
R81 B.n224 B.n69 585
R82 B.n226 B.n225 585
R83 B.n227 B.n68 585
R84 B.n229 B.n228 585
R85 B.n230 B.n67 585
R86 B.n232 B.n231 585
R87 B.n233 B.n66 585
R88 B.n235 B.n234 585
R89 B.n236 B.n65 585
R90 B.n238 B.n237 585
R91 B.n239 B.n64 585
R92 B.n241 B.n240 585
R93 B.n242 B.n63 585
R94 B.n244 B.n243 585
R95 B.n245 B.n62 585
R96 B.n247 B.n246 585
R97 B.n248 B.n61 585
R98 B.n250 B.n249 585
R99 B.n251 B.n60 585
R100 B.n253 B.n252 585
R101 B.n254 B.n59 585
R102 B.n256 B.n255 585
R103 B.n257 B.n58 585
R104 B.n259 B.n258 585
R105 B.n260 B.n57 585
R106 B.n262 B.n261 585
R107 B.n263 B.n56 585
R108 B.n265 B.n264 585
R109 B.n266 B.n55 585
R110 B.n268 B.n267 585
R111 B.n269 B.n54 585
R112 B.n271 B.n270 585
R113 B.n272 B.n53 585
R114 B.n274 B.n273 585
R115 B.n275 B.n52 585
R116 B.n277 B.n276 585
R117 B.n278 B.n51 585
R118 B.n280 B.n279 585
R119 B.n281 B.n50 585
R120 B.n283 B.n282 585
R121 B.n284 B.n49 585
R122 B.n286 B.n285 585
R123 B.n287 B.n48 585
R124 B.n289 B.n288 585
R125 B.n290 B.n47 585
R126 B.n292 B.n291 585
R127 B.n293 B.n46 585
R128 B.n295 B.n294 585
R129 B.n296 B.n45 585
R130 B.n298 B.n297 585
R131 B.n375 B.n14 585
R132 B.n374 B.n373 585
R133 B.n372 B.n15 585
R134 B.n371 B.n370 585
R135 B.n369 B.n16 585
R136 B.n368 B.n367 585
R137 B.n366 B.n17 585
R138 B.n365 B.n364 585
R139 B.n363 B.n18 585
R140 B.n362 B.n361 585
R141 B.n360 B.n19 585
R142 B.n359 B.n358 585
R143 B.n357 B.n20 585
R144 B.n356 B.n355 585
R145 B.n354 B.n21 585
R146 B.n353 B.n352 585
R147 B.n351 B.n22 585
R148 B.n350 B.n349 585
R149 B.n348 B.n23 585
R150 B.n347 B.n346 585
R151 B.n345 B.n24 585
R152 B.n344 B.n343 585
R153 B.n342 B.n25 585
R154 B.n341 B.n340 585
R155 B.n339 B.n29 585
R156 B.n338 B.n337 585
R157 B.n336 B.n30 585
R158 B.n335 B.n334 585
R159 B.n333 B.n31 585
R160 B.n332 B.n331 585
R161 B.n329 B.n32 585
R162 B.n328 B.n327 585
R163 B.n326 B.n35 585
R164 B.n325 B.n324 585
R165 B.n323 B.n36 585
R166 B.n322 B.n321 585
R167 B.n320 B.n37 585
R168 B.n319 B.n318 585
R169 B.n317 B.n38 585
R170 B.n316 B.n315 585
R171 B.n314 B.n39 585
R172 B.n313 B.n312 585
R173 B.n311 B.n40 585
R174 B.n310 B.n309 585
R175 B.n308 B.n41 585
R176 B.n307 B.n306 585
R177 B.n305 B.n42 585
R178 B.n304 B.n303 585
R179 B.n302 B.n43 585
R180 B.n301 B.n300 585
R181 B.n299 B.n44 585
R182 B.n377 B.n376 585
R183 B.n378 B.n13 585
R184 B.n380 B.n379 585
R185 B.n381 B.n12 585
R186 B.n383 B.n382 585
R187 B.n384 B.n11 585
R188 B.n386 B.n385 585
R189 B.n387 B.n10 585
R190 B.n389 B.n388 585
R191 B.n390 B.n9 585
R192 B.n392 B.n391 585
R193 B.n393 B.n8 585
R194 B.n395 B.n394 585
R195 B.n396 B.n7 585
R196 B.n398 B.n397 585
R197 B.n399 B.n6 585
R198 B.n401 B.n400 585
R199 B.n402 B.n5 585
R200 B.n404 B.n403 585
R201 B.n405 B.n4 585
R202 B.n407 B.n406 585
R203 B.n408 B.n3 585
R204 B.n410 B.n409 585
R205 B.n411 B.n0 585
R206 B.n2 B.n1 585
R207 B.n111 B.n110 585
R208 B.n113 B.n112 585
R209 B.n114 B.n109 585
R210 B.n116 B.n115 585
R211 B.n117 B.n108 585
R212 B.n119 B.n118 585
R213 B.n120 B.n107 585
R214 B.n122 B.n121 585
R215 B.n123 B.n106 585
R216 B.n125 B.n124 585
R217 B.n126 B.n105 585
R218 B.n128 B.n127 585
R219 B.n129 B.n104 585
R220 B.n131 B.n130 585
R221 B.n132 B.n103 585
R222 B.n134 B.n133 585
R223 B.n135 B.n102 585
R224 B.n137 B.n136 585
R225 B.n138 B.n101 585
R226 B.n140 B.n139 585
R227 B.n141 B.n100 585
R228 B.n143 B.n142 585
R229 B.n144 B.n99 585
R230 B.n145 B.n144 473.281
R231 B.n224 B.n223 473.281
R232 B.n297 B.n44 473.281
R233 B.n376 B.n375 473.281
R234 B.n87 B.t0 282.57
R235 B.n81 B.t9 282.57
R236 B.n33 B.t6 282.57
R237 B.n26 B.t3 282.57
R238 B.n413 B.n412 256.663
R239 B.n412 B.n411 235.042
R240 B.n412 B.n2 235.042
R241 B.n145 B.n98 163.367
R242 B.n149 B.n98 163.367
R243 B.n150 B.n149 163.367
R244 B.n151 B.n150 163.367
R245 B.n151 B.n96 163.367
R246 B.n155 B.n96 163.367
R247 B.n156 B.n155 163.367
R248 B.n157 B.n156 163.367
R249 B.n157 B.n94 163.367
R250 B.n161 B.n94 163.367
R251 B.n162 B.n161 163.367
R252 B.n163 B.n162 163.367
R253 B.n163 B.n92 163.367
R254 B.n167 B.n92 163.367
R255 B.n168 B.n167 163.367
R256 B.n169 B.n168 163.367
R257 B.n169 B.n90 163.367
R258 B.n173 B.n90 163.367
R259 B.n174 B.n173 163.367
R260 B.n175 B.n174 163.367
R261 B.n175 B.n86 163.367
R262 B.n180 B.n86 163.367
R263 B.n181 B.n180 163.367
R264 B.n182 B.n181 163.367
R265 B.n182 B.n84 163.367
R266 B.n186 B.n84 163.367
R267 B.n187 B.n186 163.367
R268 B.n188 B.n187 163.367
R269 B.n188 B.n80 163.367
R270 B.n193 B.n80 163.367
R271 B.n194 B.n193 163.367
R272 B.n195 B.n194 163.367
R273 B.n195 B.n78 163.367
R274 B.n199 B.n78 163.367
R275 B.n200 B.n199 163.367
R276 B.n201 B.n200 163.367
R277 B.n201 B.n76 163.367
R278 B.n205 B.n76 163.367
R279 B.n206 B.n205 163.367
R280 B.n207 B.n206 163.367
R281 B.n207 B.n74 163.367
R282 B.n211 B.n74 163.367
R283 B.n212 B.n211 163.367
R284 B.n213 B.n212 163.367
R285 B.n213 B.n72 163.367
R286 B.n217 B.n72 163.367
R287 B.n218 B.n217 163.367
R288 B.n219 B.n218 163.367
R289 B.n219 B.n70 163.367
R290 B.n223 B.n70 163.367
R291 B.n297 B.n296 163.367
R292 B.n296 B.n295 163.367
R293 B.n295 B.n46 163.367
R294 B.n291 B.n46 163.367
R295 B.n291 B.n290 163.367
R296 B.n290 B.n289 163.367
R297 B.n289 B.n48 163.367
R298 B.n285 B.n48 163.367
R299 B.n285 B.n284 163.367
R300 B.n284 B.n283 163.367
R301 B.n283 B.n50 163.367
R302 B.n279 B.n50 163.367
R303 B.n279 B.n278 163.367
R304 B.n278 B.n277 163.367
R305 B.n277 B.n52 163.367
R306 B.n273 B.n52 163.367
R307 B.n273 B.n272 163.367
R308 B.n272 B.n271 163.367
R309 B.n271 B.n54 163.367
R310 B.n267 B.n54 163.367
R311 B.n267 B.n266 163.367
R312 B.n266 B.n265 163.367
R313 B.n265 B.n56 163.367
R314 B.n261 B.n56 163.367
R315 B.n261 B.n260 163.367
R316 B.n260 B.n259 163.367
R317 B.n259 B.n58 163.367
R318 B.n255 B.n58 163.367
R319 B.n255 B.n254 163.367
R320 B.n254 B.n253 163.367
R321 B.n253 B.n60 163.367
R322 B.n249 B.n60 163.367
R323 B.n249 B.n248 163.367
R324 B.n248 B.n247 163.367
R325 B.n247 B.n62 163.367
R326 B.n243 B.n62 163.367
R327 B.n243 B.n242 163.367
R328 B.n242 B.n241 163.367
R329 B.n241 B.n64 163.367
R330 B.n237 B.n64 163.367
R331 B.n237 B.n236 163.367
R332 B.n236 B.n235 163.367
R333 B.n235 B.n66 163.367
R334 B.n231 B.n66 163.367
R335 B.n231 B.n230 163.367
R336 B.n230 B.n229 163.367
R337 B.n229 B.n68 163.367
R338 B.n225 B.n68 163.367
R339 B.n225 B.n224 163.367
R340 B.n375 B.n374 163.367
R341 B.n374 B.n15 163.367
R342 B.n370 B.n15 163.367
R343 B.n370 B.n369 163.367
R344 B.n369 B.n368 163.367
R345 B.n368 B.n17 163.367
R346 B.n364 B.n17 163.367
R347 B.n364 B.n363 163.367
R348 B.n363 B.n362 163.367
R349 B.n362 B.n19 163.367
R350 B.n358 B.n19 163.367
R351 B.n358 B.n357 163.367
R352 B.n357 B.n356 163.367
R353 B.n356 B.n21 163.367
R354 B.n352 B.n21 163.367
R355 B.n352 B.n351 163.367
R356 B.n351 B.n350 163.367
R357 B.n350 B.n23 163.367
R358 B.n346 B.n23 163.367
R359 B.n346 B.n345 163.367
R360 B.n345 B.n344 163.367
R361 B.n344 B.n25 163.367
R362 B.n340 B.n25 163.367
R363 B.n340 B.n339 163.367
R364 B.n339 B.n338 163.367
R365 B.n338 B.n30 163.367
R366 B.n334 B.n30 163.367
R367 B.n334 B.n333 163.367
R368 B.n333 B.n332 163.367
R369 B.n332 B.n32 163.367
R370 B.n327 B.n32 163.367
R371 B.n327 B.n326 163.367
R372 B.n326 B.n325 163.367
R373 B.n325 B.n36 163.367
R374 B.n321 B.n36 163.367
R375 B.n321 B.n320 163.367
R376 B.n320 B.n319 163.367
R377 B.n319 B.n38 163.367
R378 B.n315 B.n38 163.367
R379 B.n315 B.n314 163.367
R380 B.n314 B.n313 163.367
R381 B.n313 B.n40 163.367
R382 B.n309 B.n40 163.367
R383 B.n309 B.n308 163.367
R384 B.n308 B.n307 163.367
R385 B.n307 B.n42 163.367
R386 B.n303 B.n42 163.367
R387 B.n303 B.n302 163.367
R388 B.n302 B.n301 163.367
R389 B.n301 B.n44 163.367
R390 B.n376 B.n13 163.367
R391 B.n380 B.n13 163.367
R392 B.n381 B.n380 163.367
R393 B.n382 B.n381 163.367
R394 B.n382 B.n11 163.367
R395 B.n386 B.n11 163.367
R396 B.n387 B.n386 163.367
R397 B.n388 B.n387 163.367
R398 B.n388 B.n9 163.367
R399 B.n392 B.n9 163.367
R400 B.n393 B.n392 163.367
R401 B.n394 B.n393 163.367
R402 B.n394 B.n7 163.367
R403 B.n398 B.n7 163.367
R404 B.n399 B.n398 163.367
R405 B.n400 B.n399 163.367
R406 B.n400 B.n5 163.367
R407 B.n404 B.n5 163.367
R408 B.n405 B.n404 163.367
R409 B.n406 B.n405 163.367
R410 B.n406 B.n3 163.367
R411 B.n410 B.n3 163.367
R412 B.n411 B.n410 163.367
R413 B.n110 B.n2 163.367
R414 B.n113 B.n110 163.367
R415 B.n114 B.n113 163.367
R416 B.n115 B.n114 163.367
R417 B.n115 B.n108 163.367
R418 B.n119 B.n108 163.367
R419 B.n120 B.n119 163.367
R420 B.n121 B.n120 163.367
R421 B.n121 B.n106 163.367
R422 B.n125 B.n106 163.367
R423 B.n126 B.n125 163.367
R424 B.n127 B.n126 163.367
R425 B.n127 B.n104 163.367
R426 B.n131 B.n104 163.367
R427 B.n132 B.n131 163.367
R428 B.n133 B.n132 163.367
R429 B.n133 B.n102 163.367
R430 B.n137 B.n102 163.367
R431 B.n138 B.n137 163.367
R432 B.n139 B.n138 163.367
R433 B.n139 B.n100 163.367
R434 B.n143 B.n100 163.367
R435 B.n144 B.n143 163.367
R436 B.n81 B.t10 152.524
R437 B.n33 B.t8 152.524
R438 B.n87 B.t1 152.52
R439 B.n26 B.t5 152.52
R440 B.n82 B.t11 116.647
R441 B.n34 B.t7 116.647
R442 B.n88 B.t2 116.641
R443 B.n27 B.t4 116.641
R444 B.n177 B.n88 59.5399
R445 B.n191 B.n82 59.5399
R446 B.n330 B.n34 59.5399
R447 B.n28 B.n27 59.5399
R448 B.n88 B.n87 35.8793
R449 B.n82 B.n81 35.8793
R450 B.n34 B.n33 35.8793
R451 B.n27 B.n26 35.8793
R452 B.n377 B.n14 30.7517
R453 B.n299 B.n298 30.7517
R454 B.n222 B.n69 30.7517
R455 B.n146 B.n99 30.7517
R456 B B.n413 18.0485
R457 B.n378 B.n377 10.6151
R458 B.n379 B.n378 10.6151
R459 B.n379 B.n12 10.6151
R460 B.n383 B.n12 10.6151
R461 B.n384 B.n383 10.6151
R462 B.n385 B.n384 10.6151
R463 B.n385 B.n10 10.6151
R464 B.n389 B.n10 10.6151
R465 B.n390 B.n389 10.6151
R466 B.n391 B.n390 10.6151
R467 B.n391 B.n8 10.6151
R468 B.n395 B.n8 10.6151
R469 B.n396 B.n395 10.6151
R470 B.n397 B.n396 10.6151
R471 B.n397 B.n6 10.6151
R472 B.n401 B.n6 10.6151
R473 B.n402 B.n401 10.6151
R474 B.n403 B.n402 10.6151
R475 B.n403 B.n4 10.6151
R476 B.n407 B.n4 10.6151
R477 B.n408 B.n407 10.6151
R478 B.n409 B.n408 10.6151
R479 B.n409 B.n0 10.6151
R480 B.n373 B.n14 10.6151
R481 B.n373 B.n372 10.6151
R482 B.n372 B.n371 10.6151
R483 B.n371 B.n16 10.6151
R484 B.n367 B.n16 10.6151
R485 B.n367 B.n366 10.6151
R486 B.n366 B.n365 10.6151
R487 B.n365 B.n18 10.6151
R488 B.n361 B.n18 10.6151
R489 B.n361 B.n360 10.6151
R490 B.n360 B.n359 10.6151
R491 B.n359 B.n20 10.6151
R492 B.n355 B.n20 10.6151
R493 B.n355 B.n354 10.6151
R494 B.n354 B.n353 10.6151
R495 B.n353 B.n22 10.6151
R496 B.n349 B.n22 10.6151
R497 B.n349 B.n348 10.6151
R498 B.n348 B.n347 10.6151
R499 B.n347 B.n24 10.6151
R500 B.n343 B.n342 10.6151
R501 B.n342 B.n341 10.6151
R502 B.n341 B.n29 10.6151
R503 B.n337 B.n29 10.6151
R504 B.n337 B.n336 10.6151
R505 B.n336 B.n335 10.6151
R506 B.n335 B.n31 10.6151
R507 B.n331 B.n31 10.6151
R508 B.n329 B.n328 10.6151
R509 B.n328 B.n35 10.6151
R510 B.n324 B.n35 10.6151
R511 B.n324 B.n323 10.6151
R512 B.n323 B.n322 10.6151
R513 B.n322 B.n37 10.6151
R514 B.n318 B.n37 10.6151
R515 B.n318 B.n317 10.6151
R516 B.n317 B.n316 10.6151
R517 B.n316 B.n39 10.6151
R518 B.n312 B.n39 10.6151
R519 B.n312 B.n311 10.6151
R520 B.n311 B.n310 10.6151
R521 B.n310 B.n41 10.6151
R522 B.n306 B.n41 10.6151
R523 B.n306 B.n305 10.6151
R524 B.n305 B.n304 10.6151
R525 B.n304 B.n43 10.6151
R526 B.n300 B.n43 10.6151
R527 B.n300 B.n299 10.6151
R528 B.n298 B.n45 10.6151
R529 B.n294 B.n45 10.6151
R530 B.n294 B.n293 10.6151
R531 B.n293 B.n292 10.6151
R532 B.n292 B.n47 10.6151
R533 B.n288 B.n47 10.6151
R534 B.n288 B.n287 10.6151
R535 B.n287 B.n286 10.6151
R536 B.n286 B.n49 10.6151
R537 B.n282 B.n49 10.6151
R538 B.n282 B.n281 10.6151
R539 B.n281 B.n280 10.6151
R540 B.n280 B.n51 10.6151
R541 B.n276 B.n51 10.6151
R542 B.n276 B.n275 10.6151
R543 B.n275 B.n274 10.6151
R544 B.n274 B.n53 10.6151
R545 B.n270 B.n53 10.6151
R546 B.n270 B.n269 10.6151
R547 B.n269 B.n268 10.6151
R548 B.n268 B.n55 10.6151
R549 B.n264 B.n55 10.6151
R550 B.n264 B.n263 10.6151
R551 B.n263 B.n262 10.6151
R552 B.n262 B.n57 10.6151
R553 B.n258 B.n57 10.6151
R554 B.n258 B.n257 10.6151
R555 B.n257 B.n256 10.6151
R556 B.n256 B.n59 10.6151
R557 B.n252 B.n59 10.6151
R558 B.n252 B.n251 10.6151
R559 B.n251 B.n250 10.6151
R560 B.n250 B.n61 10.6151
R561 B.n246 B.n61 10.6151
R562 B.n246 B.n245 10.6151
R563 B.n245 B.n244 10.6151
R564 B.n244 B.n63 10.6151
R565 B.n240 B.n63 10.6151
R566 B.n240 B.n239 10.6151
R567 B.n239 B.n238 10.6151
R568 B.n238 B.n65 10.6151
R569 B.n234 B.n65 10.6151
R570 B.n234 B.n233 10.6151
R571 B.n233 B.n232 10.6151
R572 B.n232 B.n67 10.6151
R573 B.n228 B.n67 10.6151
R574 B.n228 B.n227 10.6151
R575 B.n227 B.n226 10.6151
R576 B.n226 B.n69 10.6151
R577 B.n111 B.n1 10.6151
R578 B.n112 B.n111 10.6151
R579 B.n112 B.n109 10.6151
R580 B.n116 B.n109 10.6151
R581 B.n117 B.n116 10.6151
R582 B.n118 B.n117 10.6151
R583 B.n118 B.n107 10.6151
R584 B.n122 B.n107 10.6151
R585 B.n123 B.n122 10.6151
R586 B.n124 B.n123 10.6151
R587 B.n124 B.n105 10.6151
R588 B.n128 B.n105 10.6151
R589 B.n129 B.n128 10.6151
R590 B.n130 B.n129 10.6151
R591 B.n130 B.n103 10.6151
R592 B.n134 B.n103 10.6151
R593 B.n135 B.n134 10.6151
R594 B.n136 B.n135 10.6151
R595 B.n136 B.n101 10.6151
R596 B.n140 B.n101 10.6151
R597 B.n141 B.n140 10.6151
R598 B.n142 B.n141 10.6151
R599 B.n142 B.n99 10.6151
R600 B.n147 B.n146 10.6151
R601 B.n148 B.n147 10.6151
R602 B.n148 B.n97 10.6151
R603 B.n152 B.n97 10.6151
R604 B.n153 B.n152 10.6151
R605 B.n154 B.n153 10.6151
R606 B.n154 B.n95 10.6151
R607 B.n158 B.n95 10.6151
R608 B.n159 B.n158 10.6151
R609 B.n160 B.n159 10.6151
R610 B.n160 B.n93 10.6151
R611 B.n164 B.n93 10.6151
R612 B.n165 B.n164 10.6151
R613 B.n166 B.n165 10.6151
R614 B.n166 B.n91 10.6151
R615 B.n170 B.n91 10.6151
R616 B.n171 B.n170 10.6151
R617 B.n172 B.n171 10.6151
R618 B.n172 B.n89 10.6151
R619 B.n176 B.n89 10.6151
R620 B.n179 B.n178 10.6151
R621 B.n179 B.n85 10.6151
R622 B.n183 B.n85 10.6151
R623 B.n184 B.n183 10.6151
R624 B.n185 B.n184 10.6151
R625 B.n185 B.n83 10.6151
R626 B.n189 B.n83 10.6151
R627 B.n190 B.n189 10.6151
R628 B.n192 B.n79 10.6151
R629 B.n196 B.n79 10.6151
R630 B.n197 B.n196 10.6151
R631 B.n198 B.n197 10.6151
R632 B.n198 B.n77 10.6151
R633 B.n202 B.n77 10.6151
R634 B.n203 B.n202 10.6151
R635 B.n204 B.n203 10.6151
R636 B.n204 B.n75 10.6151
R637 B.n208 B.n75 10.6151
R638 B.n209 B.n208 10.6151
R639 B.n210 B.n209 10.6151
R640 B.n210 B.n73 10.6151
R641 B.n214 B.n73 10.6151
R642 B.n215 B.n214 10.6151
R643 B.n216 B.n215 10.6151
R644 B.n216 B.n71 10.6151
R645 B.n220 B.n71 10.6151
R646 B.n221 B.n220 10.6151
R647 B.n222 B.n221 10.6151
R648 B.n413 B.n0 8.11757
R649 B.n413 B.n1 8.11757
R650 B.n343 B.n28 6.5566
R651 B.n331 B.n330 6.5566
R652 B.n178 B.n177 6.5566
R653 B.n191 B.n190 6.5566
R654 B.n28 B.n24 4.05904
R655 B.n330 B.n329 4.05904
R656 B.n177 B.n176 4.05904
R657 B.n192 B.n191 4.05904
R658 VP.n4 VP.n3 177.286
R659 VP.n12 VP.n11 177.286
R660 VP.n10 VP.n0 161.3
R661 VP.n9 VP.n8 161.3
R662 VP.n7 VP.n1 161.3
R663 VP.n6 VP.n5 161.3
R664 VP.n2 VP.t0 113.791
R665 VP.n2 VP.t2 113.472
R666 VP.n4 VP.t3 77.0571
R667 VP.n11 VP.t1 77.0571
R668 VP.n9 VP.n1 56.5617
R669 VP.n3 VP.n2 50.4587
R670 VP.n5 VP.n1 24.5923
R671 VP.n10 VP.n9 24.5923
R672 VP.n5 VP.n4 8.60764
R673 VP.n11 VP.n10 8.60764
R674 VP.n6 VP.n3 0.189894
R675 VP.n7 VP.n6 0.189894
R676 VP.n8 VP.n7 0.189894
R677 VP.n8 VP.n0 0.189894
R678 VP.n12 VP.n0 0.189894
R679 VP VP.n12 0.0516364
R680 VDD1 VDD1.n1 132.49
R681 VDD1 VDD1.n0 99.3352
R682 VDD1.n0 VDD1.t3 6.68877
R683 VDD1.n0 VDD1.t1 6.68877
R684 VDD1.n1 VDD1.t0 6.68877
R685 VDD1.n1 VDD1.t2 6.68877
C0 w_n2080_n1940# VDD2 1.08117f
C1 VTAIL VN 2.01454f
C2 VN B 0.827581f
C3 w_n2080_n1940# VP 3.44774f
C4 VDD2 VTAIL 3.43147f
C5 VDD2 B 0.913795f
C6 VTAIL VP 2.02864f
C7 B VP 1.26166f
C8 w_n2080_n1940# VTAIL 2.30656f
C9 w_n2080_n1940# B 5.9206f
C10 VDD1 VN 0.152293f
C11 VTAIL B 2.21811f
C12 VDD2 VDD1 0.764639f
C13 VDD1 VP 2.05793f
C14 w_n2080_n1940# VDD1 1.04947f
C15 VDD1 VTAIL 3.38451f
C16 VDD2 VN 1.88088f
C17 VDD1 B 0.879206f
C18 VN VP 4.0877f
C19 w_n2080_n1940# VN 3.18317f
C20 VDD2 VP 0.330187f
C21 VDD2 VSUBS 0.55118f
C22 VDD1 VSUBS 4.146778f
C23 VTAIL VSUBS 0.555296f
C24 VN VSUBS 4.41713f
C25 VP VSUBS 1.337291f
C26 B VSUBS 2.608517f
C27 w_n2080_n1940# VSUBS 50.5939f
C28 VDD1.t3 VSUBS 0.105835f
C29 VDD1.t1 VSUBS 0.105835f
C30 VDD1.n0 VSUBS 0.658304f
C31 VDD1.t0 VSUBS 0.105835f
C32 VDD1.t2 VSUBS 0.105835f
C33 VDD1.n1 VSUBS 1.01365f
C34 VP.n0 VSUBS 0.055921f
C35 VP.t1 VSUBS 1.0783f
C36 VP.n1 VSUBS 0.08129f
C37 VP.t0 VSUBS 1.29246f
C38 VP.t2 VSUBS 1.29056f
C39 VP.n2 VSUBS 2.62477f
C40 VP.n3 VSUBS 2.52944f
C41 VP.t3 VSUBS 1.0783f
C42 VP.n4 VSUBS 0.549612f
C43 VP.n5 VSUBS 0.070424f
C44 VP.n6 VSUBS 0.055921f
C45 VP.n7 VSUBS 0.055921f
C46 VP.n8 VSUBS 0.055921f
C47 VP.n9 VSUBS 0.08129f
C48 VP.n10 VSUBS 0.070424f
C49 VP.n11 VSUBS 0.549612f
C50 VP.n12 VSUBS 0.054487f
C51 B.n0 VSUBS 0.008121f
C52 B.n1 VSUBS 0.008121f
C53 B.n2 VSUBS 0.012011f
C54 B.n3 VSUBS 0.009204f
C55 B.n4 VSUBS 0.009204f
C56 B.n5 VSUBS 0.009204f
C57 B.n6 VSUBS 0.009204f
C58 B.n7 VSUBS 0.009204f
C59 B.n8 VSUBS 0.009204f
C60 B.n9 VSUBS 0.009204f
C61 B.n10 VSUBS 0.009204f
C62 B.n11 VSUBS 0.009204f
C63 B.n12 VSUBS 0.009204f
C64 B.n13 VSUBS 0.009204f
C65 B.n14 VSUBS 0.021286f
C66 B.n15 VSUBS 0.009204f
C67 B.n16 VSUBS 0.009204f
C68 B.n17 VSUBS 0.009204f
C69 B.n18 VSUBS 0.009204f
C70 B.n19 VSUBS 0.009204f
C71 B.n20 VSUBS 0.009204f
C72 B.n21 VSUBS 0.009204f
C73 B.n22 VSUBS 0.009204f
C74 B.n23 VSUBS 0.009204f
C75 B.n24 VSUBS 0.006362f
C76 B.n25 VSUBS 0.009204f
C77 B.t4 VSUBS 0.177278f
C78 B.t5 VSUBS 0.194422f
C79 B.t3 VSUBS 0.451229f
C80 B.n26 VSUBS 0.119595f
C81 B.n27 VSUBS 0.086006f
C82 B.n28 VSUBS 0.021325f
C83 B.n29 VSUBS 0.009204f
C84 B.n30 VSUBS 0.009204f
C85 B.n31 VSUBS 0.009204f
C86 B.n32 VSUBS 0.009204f
C87 B.t7 VSUBS 0.177278f
C88 B.t8 VSUBS 0.194422f
C89 B.t6 VSUBS 0.451229f
C90 B.n33 VSUBS 0.119595f
C91 B.n34 VSUBS 0.086006f
C92 B.n35 VSUBS 0.009204f
C93 B.n36 VSUBS 0.009204f
C94 B.n37 VSUBS 0.009204f
C95 B.n38 VSUBS 0.009204f
C96 B.n39 VSUBS 0.009204f
C97 B.n40 VSUBS 0.009204f
C98 B.n41 VSUBS 0.009204f
C99 B.n42 VSUBS 0.009204f
C100 B.n43 VSUBS 0.009204f
C101 B.n44 VSUBS 0.021286f
C102 B.n45 VSUBS 0.009204f
C103 B.n46 VSUBS 0.009204f
C104 B.n47 VSUBS 0.009204f
C105 B.n48 VSUBS 0.009204f
C106 B.n49 VSUBS 0.009204f
C107 B.n50 VSUBS 0.009204f
C108 B.n51 VSUBS 0.009204f
C109 B.n52 VSUBS 0.009204f
C110 B.n53 VSUBS 0.009204f
C111 B.n54 VSUBS 0.009204f
C112 B.n55 VSUBS 0.009204f
C113 B.n56 VSUBS 0.009204f
C114 B.n57 VSUBS 0.009204f
C115 B.n58 VSUBS 0.009204f
C116 B.n59 VSUBS 0.009204f
C117 B.n60 VSUBS 0.009204f
C118 B.n61 VSUBS 0.009204f
C119 B.n62 VSUBS 0.009204f
C120 B.n63 VSUBS 0.009204f
C121 B.n64 VSUBS 0.009204f
C122 B.n65 VSUBS 0.009204f
C123 B.n66 VSUBS 0.009204f
C124 B.n67 VSUBS 0.009204f
C125 B.n68 VSUBS 0.009204f
C126 B.n69 VSUBS 0.021286f
C127 B.n70 VSUBS 0.009204f
C128 B.n71 VSUBS 0.009204f
C129 B.n72 VSUBS 0.009204f
C130 B.n73 VSUBS 0.009204f
C131 B.n74 VSUBS 0.009204f
C132 B.n75 VSUBS 0.009204f
C133 B.n76 VSUBS 0.009204f
C134 B.n77 VSUBS 0.009204f
C135 B.n78 VSUBS 0.009204f
C136 B.n79 VSUBS 0.009204f
C137 B.n80 VSUBS 0.009204f
C138 B.t11 VSUBS 0.177278f
C139 B.t10 VSUBS 0.194422f
C140 B.t9 VSUBS 0.451229f
C141 B.n81 VSUBS 0.119595f
C142 B.n82 VSUBS 0.086006f
C143 B.n83 VSUBS 0.009204f
C144 B.n84 VSUBS 0.009204f
C145 B.n85 VSUBS 0.009204f
C146 B.n86 VSUBS 0.009204f
C147 B.t2 VSUBS 0.177278f
C148 B.t1 VSUBS 0.194422f
C149 B.t0 VSUBS 0.451229f
C150 B.n87 VSUBS 0.119595f
C151 B.n88 VSUBS 0.086006f
C152 B.n89 VSUBS 0.009204f
C153 B.n90 VSUBS 0.009204f
C154 B.n91 VSUBS 0.009204f
C155 B.n92 VSUBS 0.009204f
C156 B.n93 VSUBS 0.009204f
C157 B.n94 VSUBS 0.009204f
C158 B.n95 VSUBS 0.009204f
C159 B.n96 VSUBS 0.009204f
C160 B.n97 VSUBS 0.009204f
C161 B.n98 VSUBS 0.009204f
C162 B.n99 VSUBS 0.020132f
C163 B.n100 VSUBS 0.009204f
C164 B.n101 VSUBS 0.009204f
C165 B.n102 VSUBS 0.009204f
C166 B.n103 VSUBS 0.009204f
C167 B.n104 VSUBS 0.009204f
C168 B.n105 VSUBS 0.009204f
C169 B.n106 VSUBS 0.009204f
C170 B.n107 VSUBS 0.009204f
C171 B.n108 VSUBS 0.009204f
C172 B.n109 VSUBS 0.009204f
C173 B.n110 VSUBS 0.009204f
C174 B.n111 VSUBS 0.009204f
C175 B.n112 VSUBS 0.009204f
C176 B.n113 VSUBS 0.009204f
C177 B.n114 VSUBS 0.009204f
C178 B.n115 VSUBS 0.009204f
C179 B.n116 VSUBS 0.009204f
C180 B.n117 VSUBS 0.009204f
C181 B.n118 VSUBS 0.009204f
C182 B.n119 VSUBS 0.009204f
C183 B.n120 VSUBS 0.009204f
C184 B.n121 VSUBS 0.009204f
C185 B.n122 VSUBS 0.009204f
C186 B.n123 VSUBS 0.009204f
C187 B.n124 VSUBS 0.009204f
C188 B.n125 VSUBS 0.009204f
C189 B.n126 VSUBS 0.009204f
C190 B.n127 VSUBS 0.009204f
C191 B.n128 VSUBS 0.009204f
C192 B.n129 VSUBS 0.009204f
C193 B.n130 VSUBS 0.009204f
C194 B.n131 VSUBS 0.009204f
C195 B.n132 VSUBS 0.009204f
C196 B.n133 VSUBS 0.009204f
C197 B.n134 VSUBS 0.009204f
C198 B.n135 VSUBS 0.009204f
C199 B.n136 VSUBS 0.009204f
C200 B.n137 VSUBS 0.009204f
C201 B.n138 VSUBS 0.009204f
C202 B.n139 VSUBS 0.009204f
C203 B.n140 VSUBS 0.009204f
C204 B.n141 VSUBS 0.009204f
C205 B.n142 VSUBS 0.009204f
C206 B.n143 VSUBS 0.009204f
C207 B.n144 VSUBS 0.020132f
C208 B.n145 VSUBS 0.021286f
C209 B.n146 VSUBS 0.021286f
C210 B.n147 VSUBS 0.009204f
C211 B.n148 VSUBS 0.009204f
C212 B.n149 VSUBS 0.009204f
C213 B.n150 VSUBS 0.009204f
C214 B.n151 VSUBS 0.009204f
C215 B.n152 VSUBS 0.009204f
C216 B.n153 VSUBS 0.009204f
C217 B.n154 VSUBS 0.009204f
C218 B.n155 VSUBS 0.009204f
C219 B.n156 VSUBS 0.009204f
C220 B.n157 VSUBS 0.009204f
C221 B.n158 VSUBS 0.009204f
C222 B.n159 VSUBS 0.009204f
C223 B.n160 VSUBS 0.009204f
C224 B.n161 VSUBS 0.009204f
C225 B.n162 VSUBS 0.009204f
C226 B.n163 VSUBS 0.009204f
C227 B.n164 VSUBS 0.009204f
C228 B.n165 VSUBS 0.009204f
C229 B.n166 VSUBS 0.009204f
C230 B.n167 VSUBS 0.009204f
C231 B.n168 VSUBS 0.009204f
C232 B.n169 VSUBS 0.009204f
C233 B.n170 VSUBS 0.009204f
C234 B.n171 VSUBS 0.009204f
C235 B.n172 VSUBS 0.009204f
C236 B.n173 VSUBS 0.009204f
C237 B.n174 VSUBS 0.009204f
C238 B.n175 VSUBS 0.009204f
C239 B.n176 VSUBS 0.006362f
C240 B.n177 VSUBS 0.021325f
C241 B.n178 VSUBS 0.007444f
C242 B.n179 VSUBS 0.009204f
C243 B.n180 VSUBS 0.009204f
C244 B.n181 VSUBS 0.009204f
C245 B.n182 VSUBS 0.009204f
C246 B.n183 VSUBS 0.009204f
C247 B.n184 VSUBS 0.009204f
C248 B.n185 VSUBS 0.009204f
C249 B.n186 VSUBS 0.009204f
C250 B.n187 VSUBS 0.009204f
C251 B.n188 VSUBS 0.009204f
C252 B.n189 VSUBS 0.009204f
C253 B.n190 VSUBS 0.007444f
C254 B.n191 VSUBS 0.021325f
C255 B.n192 VSUBS 0.006362f
C256 B.n193 VSUBS 0.009204f
C257 B.n194 VSUBS 0.009204f
C258 B.n195 VSUBS 0.009204f
C259 B.n196 VSUBS 0.009204f
C260 B.n197 VSUBS 0.009204f
C261 B.n198 VSUBS 0.009204f
C262 B.n199 VSUBS 0.009204f
C263 B.n200 VSUBS 0.009204f
C264 B.n201 VSUBS 0.009204f
C265 B.n202 VSUBS 0.009204f
C266 B.n203 VSUBS 0.009204f
C267 B.n204 VSUBS 0.009204f
C268 B.n205 VSUBS 0.009204f
C269 B.n206 VSUBS 0.009204f
C270 B.n207 VSUBS 0.009204f
C271 B.n208 VSUBS 0.009204f
C272 B.n209 VSUBS 0.009204f
C273 B.n210 VSUBS 0.009204f
C274 B.n211 VSUBS 0.009204f
C275 B.n212 VSUBS 0.009204f
C276 B.n213 VSUBS 0.009204f
C277 B.n214 VSUBS 0.009204f
C278 B.n215 VSUBS 0.009204f
C279 B.n216 VSUBS 0.009204f
C280 B.n217 VSUBS 0.009204f
C281 B.n218 VSUBS 0.009204f
C282 B.n219 VSUBS 0.009204f
C283 B.n220 VSUBS 0.009204f
C284 B.n221 VSUBS 0.009204f
C285 B.n222 VSUBS 0.020132f
C286 B.n223 VSUBS 0.021286f
C287 B.n224 VSUBS 0.020132f
C288 B.n225 VSUBS 0.009204f
C289 B.n226 VSUBS 0.009204f
C290 B.n227 VSUBS 0.009204f
C291 B.n228 VSUBS 0.009204f
C292 B.n229 VSUBS 0.009204f
C293 B.n230 VSUBS 0.009204f
C294 B.n231 VSUBS 0.009204f
C295 B.n232 VSUBS 0.009204f
C296 B.n233 VSUBS 0.009204f
C297 B.n234 VSUBS 0.009204f
C298 B.n235 VSUBS 0.009204f
C299 B.n236 VSUBS 0.009204f
C300 B.n237 VSUBS 0.009204f
C301 B.n238 VSUBS 0.009204f
C302 B.n239 VSUBS 0.009204f
C303 B.n240 VSUBS 0.009204f
C304 B.n241 VSUBS 0.009204f
C305 B.n242 VSUBS 0.009204f
C306 B.n243 VSUBS 0.009204f
C307 B.n244 VSUBS 0.009204f
C308 B.n245 VSUBS 0.009204f
C309 B.n246 VSUBS 0.009204f
C310 B.n247 VSUBS 0.009204f
C311 B.n248 VSUBS 0.009204f
C312 B.n249 VSUBS 0.009204f
C313 B.n250 VSUBS 0.009204f
C314 B.n251 VSUBS 0.009204f
C315 B.n252 VSUBS 0.009204f
C316 B.n253 VSUBS 0.009204f
C317 B.n254 VSUBS 0.009204f
C318 B.n255 VSUBS 0.009204f
C319 B.n256 VSUBS 0.009204f
C320 B.n257 VSUBS 0.009204f
C321 B.n258 VSUBS 0.009204f
C322 B.n259 VSUBS 0.009204f
C323 B.n260 VSUBS 0.009204f
C324 B.n261 VSUBS 0.009204f
C325 B.n262 VSUBS 0.009204f
C326 B.n263 VSUBS 0.009204f
C327 B.n264 VSUBS 0.009204f
C328 B.n265 VSUBS 0.009204f
C329 B.n266 VSUBS 0.009204f
C330 B.n267 VSUBS 0.009204f
C331 B.n268 VSUBS 0.009204f
C332 B.n269 VSUBS 0.009204f
C333 B.n270 VSUBS 0.009204f
C334 B.n271 VSUBS 0.009204f
C335 B.n272 VSUBS 0.009204f
C336 B.n273 VSUBS 0.009204f
C337 B.n274 VSUBS 0.009204f
C338 B.n275 VSUBS 0.009204f
C339 B.n276 VSUBS 0.009204f
C340 B.n277 VSUBS 0.009204f
C341 B.n278 VSUBS 0.009204f
C342 B.n279 VSUBS 0.009204f
C343 B.n280 VSUBS 0.009204f
C344 B.n281 VSUBS 0.009204f
C345 B.n282 VSUBS 0.009204f
C346 B.n283 VSUBS 0.009204f
C347 B.n284 VSUBS 0.009204f
C348 B.n285 VSUBS 0.009204f
C349 B.n286 VSUBS 0.009204f
C350 B.n287 VSUBS 0.009204f
C351 B.n288 VSUBS 0.009204f
C352 B.n289 VSUBS 0.009204f
C353 B.n290 VSUBS 0.009204f
C354 B.n291 VSUBS 0.009204f
C355 B.n292 VSUBS 0.009204f
C356 B.n293 VSUBS 0.009204f
C357 B.n294 VSUBS 0.009204f
C358 B.n295 VSUBS 0.009204f
C359 B.n296 VSUBS 0.009204f
C360 B.n297 VSUBS 0.020132f
C361 B.n298 VSUBS 0.020132f
C362 B.n299 VSUBS 0.021286f
C363 B.n300 VSUBS 0.009204f
C364 B.n301 VSUBS 0.009204f
C365 B.n302 VSUBS 0.009204f
C366 B.n303 VSUBS 0.009204f
C367 B.n304 VSUBS 0.009204f
C368 B.n305 VSUBS 0.009204f
C369 B.n306 VSUBS 0.009204f
C370 B.n307 VSUBS 0.009204f
C371 B.n308 VSUBS 0.009204f
C372 B.n309 VSUBS 0.009204f
C373 B.n310 VSUBS 0.009204f
C374 B.n311 VSUBS 0.009204f
C375 B.n312 VSUBS 0.009204f
C376 B.n313 VSUBS 0.009204f
C377 B.n314 VSUBS 0.009204f
C378 B.n315 VSUBS 0.009204f
C379 B.n316 VSUBS 0.009204f
C380 B.n317 VSUBS 0.009204f
C381 B.n318 VSUBS 0.009204f
C382 B.n319 VSUBS 0.009204f
C383 B.n320 VSUBS 0.009204f
C384 B.n321 VSUBS 0.009204f
C385 B.n322 VSUBS 0.009204f
C386 B.n323 VSUBS 0.009204f
C387 B.n324 VSUBS 0.009204f
C388 B.n325 VSUBS 0.009204f
C389 B.n326 VSUBS 0.009204f
C390 B.n327 VSUBS 0.009204f
C391 B.n328 VSUBS 0.009204f
C392 B.n329 VSUBS 0.006362f
C393 B.n330 VSUBS 0.021325f
C394 B.n331 VSUBS 0.007444f
C395 B.n332 VSUBS 0.009204f
C396 B.n333 VSUBS 0.009204f
C397 B.n334 VSUBS 0.009204f
C398 B.n335 VSUBS 0.009204f
C399 B.n336 VSUBS 0.009204f
C400 B.n337 VSUBS 0.009204f
C401 B.n338 VSUBS 0.009204f
C402 B.n339 VSUBS 0.009204f
C403 B.n340 VSUBS 0.009204f
C404 B.n341 VSUBS 0.009204f
C405 B.n342 VSUBS 0.009204f
C406 B.n343 VSUBS 0.007444f
C407 B.n344 VSUBS 0.009204f
C408 B.n345 VSUBS 0.009204f
C409 B.n346 VSUBS 0.009204f
C410 B.n347 VSUBS 0.009204f
C411 B.n348 VSUBS 0.009204f
C412 B.n349 VSUBS 0.009204f
C413 B.n350 VSUBS 0.009204f
C414 B.n351 VSUBS 0.009204f
C415 B.n352 VSUBS 0.009204f
C416 B.n353 VSUBS 0.009204f
C417 B.n354 VSUBS 0.009204f
C418 B.n355 VSUBS 0.009204f
C419 B.n356 VSUBS 0.009204f
C420 B.n357 VSUBS 0.009204f
C421 B.n358 VSUBS 0.009204f
C422 B.n359 VSUBS 0.009204f
C423 B.n360 VSUBS 0.009204f
C424 B.n361 VSUBS 0.009204f
C425 B.n362 VSUBS 0.009204f
C426 B.n363 VSUBS 0.009204f
C427 B.n364 VSUBS 0.009204f
C428 B.n365 VSUBS 0.009204f
C429 B.n366 VSUBS 0.009204f
C430 B.n367 VSUBS 0.009204f
C431 B.n368 VSUBS 0.009204f
C432 B.n369 VSUBS 0.009204f
C433 B.n370 VSUBS 0.009204f
C434 B.n371 VSUBS 0.009204f
C435 B.n372 VSUBS 0.009204f
C436 B.n373 VSUBS 0.009204f
C437 B.n374 VSUBS 0.009204f
C438 B.n375 VSUBS 0.021286f
C439 B.n376 VSUBS 0.020132f
C440 B.n377 VSUBS 0.020132f
C441 B.n378 VSUBS 0.009204f
C442 B.n379 VSUBS 0.009204f
C443 B.n380 VSUBS 0.009204f
C444 B.n381 VSUBS 0.009204f
C445 B.n382 VSUBS 0.009204f
C446 B.n383 VSUBS 0.009204f
C447 B.n384 VSUBS 0.009204f
C448 B.n385 VSUBS 0.009204f
C449 B.n386 VSUBS 0.009204f
C450 B.n387 VSUBS 0.009204f
C451 B.n388 VSUBS 0.009204f
C452 B.n389 VSUBS 0.009204f
C453 B.n390 VSUBS 0.009204f
C454 B.n391 VSUBS 0.009204f
C455 B.n392 VSUBS 0.009204f
C456 B.n393 VSUBS 0.009204f
C457 B.n394 VSUBS 0.009204f
C458 B.n395 VSUBS 0.009204f
C459 B.n396 VSUBS 0.009204f
C460 B.n397 VSUBS 0.009204f
C461 B.n398 VSUBS 0.009204f
C462 B.n399 VSUBS 0.009204f
C463 B.n400 VSUBS 0.009204f
C464 B.n401 VSUBS 0.009204f
C465 B.n402 VSUBS 0.009204f
C466 B.n403 VSUBS 0.009204f
C467 B.n404 VSUBS 0.009204f
C468 B.n405 VSUBS 0.009204f
C469 B.n406 VSUBS 0.009204f
C470 B.n407 VSUBS 0.009204f
C471 B.n408 VSUBS 0.009204f
C472 B.n409 VSUBS 0.009204f
C473 B.n410 VSUBS 0.009204f
C474 B.n411 VSUBS 0.012011f
C475 B.n412 VSUBS 0.012795f
C476 B.n413 VSUBS 0.025443f
C477 VTAIL.t6 VSUBS 0.797003f
C478 VTAIL.n0 VSUBS 0.632362f
C479 VTAIL.t2 VSUBS 0.797003f
C480 VTAIL.n1 VSUBS 0.697246f
C481 VTAIL.t0 VSUBS 0.797003f
C482 VTAIL.n2 VSUBS 1.53375f
C483 VTAIL.t7 VSUBS 0.797008f
C484 VTAIL.n3 VSUBS 1.53374f
C485 VTAIL.t5 VSUBS 0.797008f
C486 VTAIL.n4 VSUBS 0.697241f
C487 VTAIL.t1 VSUBS 0.797008f
C488 VTAIL.n5 VSUBS 0.697241f
C489 VTAIL.t3 VSUBS 0.797003f
C490 VTAIL.n6 VSUBS 1.53375f
C491 VTAIL.t4 VSUBS 0.797003f
C492 VTAIL.n7 VSUBS 1.45865f
C493 VDD2.t0 VSUBS 0.066659f
C494 VDD2.t1 VSUBS 0.066659f
C495 VDD2.n0 VSUBS 0.626999f
C496 VDD2.t2 VSUBS 0.066659f
C497 VDD2.t3 VSUBS 0.066659f
C498 VDD2.n1 VSUBS 0.414411f
C499 VDD2.n2 VSUBS 1.99902f
C500 VN.t1 VSUBS 1.02922f
C501 VN.t3 VSUBS 1.02771f
C502 VN.n0 VSUBS 0.783263f
C503 VN.t2 VSUBS 1.02922f
C504 VN.t0 VSUBS 1.02771f
C505 VN.n1 VSUBS 2.11551f
.ends

