* NGSPICE file created from diff_pair_sample_1360.ext - technology: sky130A

.subckt diff_pair_sample_1360 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t3 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0.7854 ps=5.09 w=4.76 l=2.57
X1 VTAIL.t1 VN.t0 VDD2.t3 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0.7854 ps=5.09 w=4.76 l=2.57
X2 VDD1.t1 VP.t1 VTAIL.t6 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=0.7854 pd=5.09 as=1.8564 ps=10.3 w=4.76 l=2.57
X3 B.t11 B.t9 B.t10 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0 ps=0 w=4.76 l=2.57
X4 VTAIL.t5 VP.t2 VDD1.t0 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0.7854 ps=5.09 w=4.76 l=2.57
X5 VDD2.t2 VN.t1 VTAIL.t3 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=0.7854 pd=5.09 as=1.8564 ps=10.3 w=4.76 l=2.57
X6 VDD2.t1 VN.t2 VTAIL.t0 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=0.7854 pd=5.09 as=1.8564 ps=10.3 w=4.76 l=2.57
X7 B.t8 B.t6 B.t7 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0 ps=0 w=4.76 l=2.57
X8 VTAIL.t2 VN.t3 VDD2.t0 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0.7854 ps=5.09 w=4.76 l=2.57
X9 B.t5 B.t3 B.t4 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0 ps=0 w=4.76 l=2.57
X10 B.t2 B.t0 B.t1 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=1.8564 pd=10.3 as=0 ps=0 w=4.76 l=2.57
X11 VDD1.t2 VP.t3 VTAIL.t4 w_n2710_n1920# sky130_fd_pr__pfet_01v8 ad=0.7854 pd=5.09 as=1.8564 ps=10.3 w=4.76 l=2.57
R0 VP.n14 VP.n0 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n11 VP.n1 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n8 VP.n2 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n5 VP.n3 101.072
R7 VP.n16 VP.n15 101.072
R8 VP.n4 VP.t2 80.6876
R9 VP.n4 VP.t3 79.9167
R10 VP.n9 VP.n1 56.5617
R11 VP.n5 VP.n4 45.1091
R12 VP.n3 VP.t0 44.6371
R13 VP.n15 VP.t1 44.6371
R14 VP.n8 VP.n7 24.5923
R15 VP.n9 VP.n8 24.5923
R16 VP.n13 VP.n1 24.5923
R17 VP.n14 VP.n13 24.5923
R18 VP.n7 VP.n3 9.83723
R19 VP.n15 VP.n14 9.83723
R20 VP.n6 VP.n5 0.278335
R21 VP.n16 VP.n0 0.278335
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153485
R28 VDD1 VDD1.n1 143.802
R29 VDD1 VDD1.n0 108.016
R30 VDD1.n0 VDD1.t0 6.82928
R31 VDD1.n0 VDD1.t2 6.82928
R32 VDD1.n1 VDD1.t3 6.82928
R33 VDD1.n1 VDD1.t1 6.82928
R34 VTAIL.n186 VTAIL.n168 756.745
R35 VTAIL.n18 VTAIL.n0 756.745
R36 VTAIL.n42 VTAIL.n24 756.745
R37 VTAIL.n66 VTAIL.n48 756.745
R38 VTAIL.n162 VTAIL.n144 756.745
R39 VTAIL.n138 VTAIL.n120 756.745
R40 VTAIL.n114 VTAIL.n96 756.745
R41 VTAIL.n90 VTAIL.n72 756.745
R42 VTAIL.n177 VTAIL.n176 585
R43 VTAIL.n179 VTAIL.n178 585
R44 VTAIL.n172 VTAIL.n171 585
R45 VTAIL.n185 VTAIL.n184 585
R46 VTAIL.n187 VTAIL.n186 585
R47 VTAIL.n9 VTAIL.n8 585
R48 VTAIL.n11 VTAIL.n10 585
R49 VTAIL.n4 VTAIL.n3 585
R50 VTAIL.n17 VTAIL.n16 585
R51 VTAIL.n19 VTAIL.n18 585
R52 VTAIL.n33 VTAIL.n32 585
R53 VTAIL.n35 VTAIL.n34 585
R54 VTAIL.n28 VTAIL.n27 585
R55 VTAIL.n41 VTAIL.n40 585
R56 VTAIL.n43 VTAIL.n42 585
R57 VTAIL.n57 VTAIL.n56 585
R58 VTAIL.n59 VTAIL.n58 585
R59 VTAIL.n52 VTAIL.n51 585
R60 VTAIL.n65 VTAIL.n64 585
R61 VTAIL.n67 VTAIL.n66 585
R62 VTAIL.n163 VTAIL.n162 585
R63 VTAIL.n161 VTAIL.n160 585
R64 VTAIL.n148 VTAIL.n147 585
R65 VTAIL.n155 VTAIL.n154 585
R66 VTAIL.n153 VTAIL.n152 585
R67 VTAIL.n139 VTAIL.n138 585
R68 VTAIL.n137 VTAIL.n136 585
R69 VTAIL.n124 VTAIL.n123 585
R70 VTAIL.n131 VTAIL.n130 585
R71 VTAIL.n129 VTAIL.n128 585
R72 VTAIL.n115 VTAIL.n114 585
R73 VTAIL.n113 VTAIL.n112 585
R74 VTAIL.n100 VTAIL.n99 585
R75 VTAIL.n107 VTAIL.n106 585
R76 VTAIL.n105 VTAIL.n104 585
R77 VTAIL.n91 VTAIL.n90 585
R78 VTAIL.n89 VTAIL.n88 585
R79 VTAIL.n76 VTAIL.n75 585
R80 VTAIL.n83 VTAIL.n82 585
R81 VTAIL.n81 VTAIL.n80 585
R82 VTAIL.n175 VTAIL.t0 328.587
R83 VTAIL.n7 VTAIL.t2 328.587
R84 VTAIL.n31 VTAIL.t6 328.587
R85 VTAIL.n55 VTAIL.t7 328.587
R86 VTAIL.n151 VTAIL.t4 328.587
R87 VTAIL.n127 VTAIL.t5 328.587
R88 VTAIL.n103 VTAIL.t3 328.587
R89 VTAIL.n79 VTAIL.t1 328.587
R90 VTAIL.n178 VTAIL.n177 171.744
R91 VTAIL.n178 VTAIL.n171 171.744
R92 VTAIL.n185 VTAIL.n171 171.744
R93 VTAIL.n186 VTAIL.n185 171.744
R94 VTAIL.n10 VTAIL.n9 171.744
R95 VTAIL.n10 VTAIL.n3 171.744
R96 VTAIL.n17 VTAIL.n3 171.744
R97 VTAIL.n18 VTAIL.n17 171.744
R98 VTAIL.n34 VTAIL.n33 171.744
R99 VTAIL.n34 VTAIL.n27 171.744
R100 VTAIL.n41 VTAIL.n27 171.744
R101 VTAIL.n42 VTAIL.n41 171.744
R102 VTAIL.n58 VTAIL.n57 171.744
R103 VTAIL.n58 VTAIL.n51 171.744
R104 VTAIL.n65 VTAIL.n51 171.744
R105 VTAIL.n66 VTAIL.n65 171.744
R106 VTAIL.n162 VTAIL.n161 171.744
R107 VTAIL.n161 VTAIL.n147 171.744
R108 VTAIL.n154 VTAIL.n147 171.744
R109 VTAIL.n154 VTAIL.n153 171.744
R110 VTAIL.n138 VTAIL.n137 171.744
R111 VTAIL.n137 VTAIL.n123 171.744
R112 VTAIL.n130 VTAIL.n123 171.744
R113 VTAIL.n130 VTAIL.n129 171.744
R114 VTAIL.n114 VTAIL.n113 171.744
R115 VTAIL.n113 VTAIL.n99 171.744
R116 VTAIL.n106 VTAIL.n99 171.744
R117 VTAIL.n106 VTAIL.n105 171.744
R118 VTAIL.n90 VTAIL.n89 171.744
R119 VTAIL.n89 VTAIL.n75 171.744
R120 VTAIL.n82 VTAIL.n75 171.744
R121 VTAIL.n82 VTAIL.n81 171.744
R122 VTAIL.n177 VTAIL.t0 85.8723
R123 VTAIL.n9 VTAIL.t2 85.8723
R124 VTAIL.n33 VTAIL.t6 85.8723
R125 VTAIL.n57 VTAIL.t7 85.8723
R126 VTAIL.n153 VTAIL.t4 85.8723
R127 VTAIL.n129 VTAIL.t5 85.8723
R128 VTAIL.n105 VTAIL.t3 85.8723
R129 VTAIL.n81 VTAIL.t1 85.8723
R130 VTAIL.n191 VTAIL.n190 36.0641
R131 VTAIL.n23 VTAIL.n22 36.0641
R132 VTAIL.n47 VTAIL.n46 36.0641
R133 VTAIL.n71 VTAIL.n70 36.0641
R134 VTAIL.n167 VTAIL.n166 36.0641
R135 VTAIL.n143 VTAIL.n142 36.0641
R136 VTAIL.n119 VTAIL.n118 36.0641
R137 VTAIL.n95 VTAIL.n94 36.0641
R138 VTAIL.n191 VTAIL.n167 18.9703
R139 VTAIL.n95 VTAIL.n71 18.9703
R140 VTAIL.n176 VTAIL.n175 16.3651
R141 VTAIL.n8 VTAIL.n7 16.3651
R142 VTAIL.n32 VTAIL.n31 16.3651
R143 VTAIL.n56 VTAIL.n55 16.3651
R144 VTAIL.n152 VTAIL.n151 16.3651
R145 VTAIL.n128 VTAIL.n127 16.3651
R146 VTAIL.n104 VTAIL.n103 16.3651
R147 VTAIL.n80 VTAIL.n79 16.3651
R148 VTAIL.n179 VTAIL.n174 12.8005
R149 VTAIL.n11 VTAIL.n6 12.8005
R150 VTAIL.n35 VTAIL.n30 12.8005
R151 VTAIL.n59 VTAIL.n54 12.8005
R152 VTAIL.n155 VTAIL.n150 12.8005
R153 VTAIL.n131 VTAIL.n126 12.8005
R154 VTAIL.n107 VTAIL.n102 12.8005
R155 VTAIL.n83 VTAIL.n78 12.8005
R156 VTAIL.n180 VTAIL.n172 12.0247
R157 VTAIL.n12 VTAIL.n4 12.0247
R158 VTAIL.n36 VTAIL.n28 12.0247
R159 VTAIL.n60 VTAIL.n52 12.0247
R160 VTAIL.n156 VTAIL.n148 12.0247
R161 VTAIL.n132 VTAIL.n124 12.0247
R162 VTAIL.n108 VTAIL.n100 12.0247
R163 VTAIL.n84 VTAIL.n76 12.0247
R164 VTAIL.n184 VTAIL.n183 11.249
R165 VTAIL.n16 VTAIL.n15 11.249
R166 VTAIL.n40 VTAIL.n39 11.249
R167 VTAIL.n64 VTAIL.n63 11.249
R168 VTAIL.n160 VTAIL.n159 11.249
R169 VTAIL.n136 VTAIL.n135 11.249
R170 VTAIL.n112 VTAIL.n111 11.249
R171 VTAIL.n88 VTAIL.n87 11.249
R172 VTAIL.n187 VTAIL.n170 10.4732
R173 VTAIL.n19 VTAIL.n2 10.4732
R174 VTAIL.n43 VTAIL.n26 10.4732
R175 VTAIL.n67 VTAIL.n50 10.4732
R176 VTAIL.n163 VTAIL.n146 10.4732
R177 VTAIL.n139 VTAIL.n122 10.4732
R178 VTAIL.n115 VTAIL.n98 10.4732
R179 VTAIL.n91 VTAIL.n74 10.4732
R180 VTAIL.n188 VTAIL.n168 9.69747
R181 VTAIL.n20 VTAIL.n0 9.69747
R182 VTAIL.n44 VTAIL.n24 9.69747
R183 VTAIL.n68 VTAIL.n48 9.69747
R184 VTAIL.n164 VTAIL.n144 9.69747
R185 VTAIL.n140 VTAIL.n120 9.69747
R186 VTAIL.n116 VTAIL.n96 9.69747
R187 VTAIL.n92 VTAIL.n72 9.69747
R188 VTAIL.n190 VTAIL.n189 9.45567
R189 VTAIL.n22 VTAIL.n21 9.45567
R190 VTAIL.n46 VTAIL.n45 9.45567
R191 VTAIL.n70 VTAIL.n69 9.45567
R192 VTAIL.n166 VTAIL.n165 9.45567
R193 VTAIL.n142 VTAIL.n141 9.45567
R194 VTAIL.n118 VTAIL.n117 9.45567
R195 VTAIL.n94 VTAIL.n93 9.45567
R196 VTAIL.n189 VTAIL.n188 9.3005
R197 VTAIL.n170 VTAIL.n169 9.3005
R198 VTAIL.n183 VTAIL.n182 9.3005
R199 VTAIL.n181 VTAIL.n180 9.3005
R200 VTAIL.n174 VTAIL.n173 9.3005
R201 VTAIL.n21 VTAIL.n20 9.3005
R202 VTAIL.n2 VTAIL.n1 9.3005
R203 VTAIL.n15 VTAIL.n14 9.3005
R204 VTAIL.n13 VTAIL.n12 9.3005
R205 VTAIL.n6 VTAIL.n5 9.3005
R206 VTAIL.n45 VTAIL.n44 9.3005
R207 VTAIL.n26 VTAIL.n25 9.3005
R208 VTAIL.n39 VTAIL.n38 9.3005
R209 VTAIL.n37 VTAIL.n36 9.3005
R210 VTAIL.n30 VTAIL.n29 9.3005
R211 VTAIL.n69 VTAIL.n68 9.3005
R212 VTAIL.n50 VTAIL.n49 9.3005
R213 VTAIL.n63 VTAIL.n62 9.3005
R214 VTAIL.n61 VTAIL.n60 9.3005
R215 VTAIL.n54 VTAIL.n53 9.3005
R216 VTAIL.n165 VTAIL.n164 9.3005
R217 VTAIL.n146 VTAIL.n145 9.3005
R218 VTAIL.n159 VTAIL.n158 9.3005
R219 VTAIL.n157 VTAIL.n156 9.3005
R220 VTAIL.n150 VTAIL.n149 9.3005
R221 VTAIL.n141 VTAIL.n140 9.3005
R222 VTAIL.n122 VTAIL.n121 9.3005
R223 VTAIL.n135 VTAIL.n134 9.3005
R224 VTAIL.n133 VTAIL.n132 9.3005
R225 VTAIL.n126 VTAIL.n125 9.3005
R226 VTAIL.n117 VTAIL.n116 9.3005
R227 VTAIL.n98 VTAIL.n97 9.3005
R228 VTAIL.n111 VTAIL.n110 9.3005
R229 VTAIL.n109 VTAIL.n108 9.3005
R230 VTAIL.n102 VTAIL.n101 9.3005
R231 VTAIL.n93 VTAIL.n92 9.3005
R232 VTAIL.n74 VTAIL.n73 9.3005
R233 VTAIL.n87 VTAIL.n86 9.3005
R234 VTAIL.n85 VTAIL.n84 9.3005
R235 VTAIL.n78 VTAIL.n77 9.3005
R236 VTAIL.n190 VTAIL.n168 4.26717
R237 VTAIL.n22 VTAIL.n0 4.26717
R238 VTAIL.n46 VTAIL.n24 4.26717
R239 VTAIL.n70 VTAIL.n48 4.26717
R240 VTAIL.n166 VTAIL.n144 4.26717
R241 VTAIL.n142 VTAIL.n120 4.26717
R242 VTAIL.n118 VTAIL.n96 4.26717
R243 VTAIL.n94 VTAIL.n72 4.26717
R244 VTAIL.n175 VTAIL.n173 3.73474
R245 VTAIL.n7 VTAIL.n5 3.73474
R246 VTAIL.n31 VTAIL.n29 3.73474
R247 VTAIL.n55 VTAIL.n53 3.73474
R248 VTAIL.n151 VTAIL.n149 3.73474
R249 VTAIL.n127 VTAIL.n125 3.73474
R250 VTAIL.n103 VTAIL.n101 3.73474
R251 VTAIL.n79 VTAIL.n77 3.73474
R252 VTAIL.n188 VTAIL.n187 3.49141
R253 VTAIL.n20 VTAIL.n19 3.49141
R254 VTAIL.n44 VTAIL.n43 3.49141
R255 VTAIL.n68 VTAIL.n67 3.49141
R256 VTAIL.n164 VTAIL.n163 3.49141
R257 VTAIL.n140 VTAIL.n139 3.49141
R258 VTAIL.n116 VTAIL.n115 3.49141
R259 VTAIL.n92 VTAIL.n91 3.49141
R260 VTAIL.n184 VTAIL.n170 2.71565
R261 VTAIL.n16 VTAIL.n2 2.71565
R262 VTAIL.n40 VTAIL.n26 2.71565
R263 VTAIL.n64 VTAIL.n50 2.71565
R264 VTAIL.n160 VTAIL.n146 2.71565
R265 VTAIL.n136 VTAIL.n122 2.71565
R266 VTAIL.n112 VTAIL.n98 2.71565
R267 VTAIL.n88 VTAIL.n74 2.71565
R268 VTAIL.n119 VTAIL.n95 2.5005
R269 VTAIL.n167 VTAIL.n143 2.5005
R270 VTAIL.n71 VTAIL.n47 2.5005
R271 VTAIL.n183 VTAIL.n172 1.93989
R272 VTAIL.n15 VTAIL.n4 1.93989
R273 VTAIL.n39 VTAIL.n28 1.93989
R274 VTAIL.n63 VTAIL.n52 1.93989
R275 VTAIL.n159 VTAIL.n148 1.93989
R276 VTAIL.n135 VTAIL.n124 1.93989
R277 VTAIL.n111 VTAIL.n100 1.93989
R278 VTAIL.n87 VTAIL.n76 1.93989
R279 VTAIL VTAIL.n23 1.30869
R280 VTAIL VTAIL.n191 1.19231
R281 VTAIL.n180 VTAIL.n179 1.16414
R282 VTAIL.n12 VTAIL.n11 1.16414
R283 VTAIL.n36 VTAIL.n35 1.16414
R284 VTAIL.n60 VTAIL.n59 1.16414
R285 VTAIL.n156 VTAIL.n155 1.16414
R286 VTAIL.n132 VTAIL.n131 1.16414
R287 VTAIL.n108 VTAIL.n107 1.16414
R288 VTAIL.n84 VTAIL.n83 1.16414
R289 VTAIL.n143 VTAIL.n119 0.470328
R290 VTAIL.n47 VTAIL.n23 0.470328
R291 VTAIL.n176 VTAIL.n174 0.388379
R292 VTAIL.n8 VTAIL.n6 0.388379
R293 VTAIL.n32 VTAIL.n30 0.388379
R294 VTAIL.n56 VTAIL.n54 0.388379
R295 VTAIL.n152 VTAIL.n150 0.388379
R296 VTAIL.n128 VTAIL.n126 0.388379
R297 VTAIL.n104 VTAIL.n102 0.388379
R298 VTAIL.n80 VTAIL.n78 0.388379
R299 VTAIL.n181 VTAIL.n173 0.155672
R300 VTAIL.n182 VTAIL.n181 0.155672
R301 VTAIL.n182 VTAIL.n169 0.155672
R302 VTAIL.n189 VTAIL.n169 0.155672
R303 VTAIL.n13 VTAIL.n5 0.155672
R304 VTAIL.n14 VTAIL.n13 0.155672
R305 VTAIL.n14 VTAIL.n1 0.155672
R306 VTAIL.n21 VTAIL.n1 0.155672
R307 VTAIL.n37 VTAIL.n29 0.155672
R308 VTAIL.n38 VTAIL.n37 0.155672
R309 VTAIL.n38 VTAIL.n25 0.155672
R310 VTAIL.n45 VTAIL.n25 0.155672
R311 VTAIL.n61 VTAIL.n53 0.155672
R312 VTAIL.n62 VTAIL.n61 0.155672
R313 VTAIL.n62 VTAIL.n49 0.155672
R314 VTAIL.n69 VTAIL.n49 0.155672
R315 VTAIL.n165 VTAIL.n145 0.155672
R316 VTAIL.n158 VTAIL.n145 0.155672
R317 VTAIL.n158 VTAIL.n157 0.155672
R318 VTAIL.n157 VTAIL.n149 0.155672
R319 VTAIL.n141 VTAIL.n121 0.155672
R320 VTAIL.n134 VTAIL.n121 0.155672
R321 VTAIL.n134 VTAIL.n133 0.155672
R322 VTAIL.n133 VTAIL.n125 0.155672
R323 VTAIL.n117 VTAIL.n97 0.155672
R324 VTAIL.n110 VTAIL.n97 0.155672
R325 VTAIL.n110 VTAIL.n109 0.155672
R326 VTAIL.n109 VTAIL.n101 0.155672
R327 VTAIL.n93 VTAIL.n73 0.155672
R328 VTAIL.n86 VTAIL.n73 0.155672
R329 VTAIL.n86 VTAIL.n85 0.155672
R330 VTAIL.n85 VTAIL.n77 0.155672
R331 VN.n0 VN.t3 80.6876
R332 VN.n1 VN.t1 80.6876
R333 VN.n0 VN.t2 79.9167
R334 VN.n1 VN.t0 79.9167
R335 VN VN.n1 45.3879
R336 VN VN.n0 4.37656
R337 VDD2.n2 VDD2.n0 143.276
R338 VDD2.n2 VDD2.n1 107.959
R339 VDD2.n1 VDD2.t3 6.82928
R340 VDD2.n1 VDD2.t2 6.82928
R341 VDD2.n0 VDD2.t0 6.82928
R342 VDD2.n0 VDD2.t1 6.82928
R343 VDD2 VDD2.n2 0.0586897
R344 B.n252 B.n251 585
R345 B.n250 B.n83 585
R346 B.n249 B.n248 585
R347 B.n247 B.n84 585
R348 B.n246 B.n245 585
R349 B.n244 B.n85 585
R350 B.n243 B.n242 585
R351 B.n241 B.n86 585
R352 B.n240 B.n239 585
R353 B.n238 B.n87 585
R354 B.n237 B.n236 585
R355 B.n235 B.n88 585
R356 B.n234 B.n233 585
R357 B.n232 B.n89 585
R358 B.n231 B.n230 585
R359 B.n229 B.n90 585
R360 B.n228 B.n227 585
R361 B.n226 B.n91 585
R362 B.n225 B.n224 585
R363 B.n223 B.n92 585
R364 B.n221 B.n220 585
R365 B.n219 B.n95 585
R366 B.n218 B.n217 585
R367 B.n216 B.n96 585
R368 B.n215 B.n214 585
R369 B.n213 B.n97 585
R370 B.n212 B.n211 585
R371 B.n210 B.n98 585
R372 B.n209 B.n208 585
R373 B.n207 B.n99 585
R374 B.n206 B.n205 585
R375 B.n201 B.n100 585
R376 B.n200 B.n199 585
R377 B.n198 B.n101 585
R378 B.n197 B.n196 585
R379 B.n195 B.n102 585
R380 B.n194 B.n193 585
R381 B.n192 B.n103 585
R382 B.n191 B.n190 585
R383 B.n189 B.n104 585
R384 B.n188 B.n187 585
R385 B.n186 B.n105 585
R386 B.n185 B.n184 585
R387 B.n183 B.n106 585
R388 B.n182 B.n181 585
R389 B.n180 B.n107 585
R390 B.n179 B.n178 585
R391 B.n177 B.n108 585
R392 B.n176 B.n175 585
R393 B.n174 B.n109 585
R394 B.n253 B.n82 585
R395 B.n255 B.n254 585
R396 B.n256 B.n81 585
R397 B.n258 B.n257 585
R398 B.n259 B.n80 585
R399 B.n261 B.n260 585
R400 B.n262 B.n79 585
R401 B.n264 B.n263 585
R402 B.n265 B.n78 585
R403 B.n267 B.n266 585
R404 B.n268 B.n77 585
R405 B.n270 B.n269 585
R406 B.n271 B.n76 585
R407 B.n273 B.n272 585
R408 B.n274 B.n75 585
R409 B.n276 B.n275 585
R410 B.n277 B.n74 585
R411 B.n279 B.n278 585
R412 B.n280 B.n73 585
R413 B.n282 B.n281 585
R414 B.n283 B.n72 585
R415 B.n285 B.n284 585
R416 B.n286 B.n71 585
R417 B.n288 B.n287 585
R418 B.n289 B.n70 585
R419 B.n291 B.n290 585
R420 B.n292 B.n69 585
R421 B.n294 B.n293 585
R422 B.n295 B.n68 585
R423 B.n297 B.n296 585
R424 B.n298 B.n67 585
R425 B.n300 B.n299 585
R426 B.n301 B.n66 585
R427 B.n303 B.n302 585
R428 B.n304 B.n65 585
R429 B.n306 B.n305 585
R430 B.n307 B.n64 585
R431 B.n309 B.n308 585
R432 B.n310 B.n63 585
R433 B.n312 B.n311 585
R434 B.n313 B.n62 585
R435 B.n315 B.n314 585
R436 B.n316 B.n61 585
R437 B.n318 B.n317 585
R438 B.n319 B.n60 585
R439 B.n321 B.n320 585
R440 B.n322 B.n59 585
R441 B.n324 B.n323 585
R442 B.n325 B.n58 585
R443 B.n327 B.n326 585
R444 B.n328 B.n57 585
R445 B.n330 B.n329 585
R446 B.n331 B.n56 585
R447 B.n333 B.n332 585
R448 B.n334 B.n55 585
R449 B.n336 B.n335 585
R450 B.n337 B.n54 585
R451 B.n339 B.n338 585
R452 B.n340 B.n53 585
R453 B.n342 B.n341 585
R454 B.n343 B.n52 585
R455 B.n345 B.n344 585
R456 B.n346 B.n51 585
R457 B.n348 B.n347 585
R458 B.n349 B.n50 585
R459 B.n351 B.n350 585
R460 B.n352 B.n49 585
R461 B.n354 B.n353 585
R462 B.n430 B.n429 585
R463 B.n428 B.n19 585
R464 B.n427 B.n426 585
R465 B.n425 B.n20 585
R466 B.n424 B.n423 585
R467 B.n422 B.n21 585
R468 B.n421 B.n420 585
R469 B.n419 B.n22 585
R470 B.n418 B.n417 585
R471 B.n416 B.n23 585
R472 B.n415 B.n414 585
R473 B.n413 B.n24 585
R474 B.n412 B.n411 585
R475 B.n410 B.n25 585
R476 B.n409 B.n408 585
R477 B.n407 B.n26 585
R478 B.n406 B.n405 585
R479 B.n404 B.n27 585
R480 B.n403 B.n402 585
R481 B.n401 B.n28 585
R482 B.n400 B.n399 585
R483 B.n398 B.n29 585
R484 B.n397 B.n396 585
R485 B.n395 B.n33 585
R486 B.n394 B.n393 585
R487 B.n392 B.n34 585
R488 B.n391 B.n390 585
R489 B.n389 B.n35 585
R490 B.n388 B.n387 585
R491 B.n386 B.n36 585
R492 B.n384 B.n383 585
R493 B.n382 B.n39 585
R494 B.n381 B.n380 585
R495 B.n379 B.n40 585
R496 B.n378 B.n377 585
R497 B.n376 B.n41 585
R498 B.n375 B.n374 585
R499 B.n373 B.n42 585
R500 B.n372 B.n371 585
R501 B.n370 B.n43 585
R502 B.n369 B.n368 585
R503 B.n367 B.n44 585
R504 B.n366 B.n365 585
R505 B.n364 B.n45 585
R506 B.n363 B.n362 585
R507 B.n361 B.n46 585
R508 B.n360 B.n359 585
R509 B.n358 B.n47 585
R510 B.n357 B.n356 585
R511 B.n355 B.n48 585
R512 B.n431 B.n18 585
R513 B.n433 B.n432 585
R514 B.n434 B.n17 585
R515 B.n436 B.n435 585
R516 B.n437 B.n16 585
R517 B.n439 B.n438 585
R518 B.n440 B.n15 585
R519 B.n442 B.n441 585
R520 B.n443 B.n14 585
R521 B.n445 B.n444 585
R522 B.n446 B.n13 585
R523 B.n448 B.n447 585
R524 B.n449 B.n12 585
R525 B.n451 B.n450 585
R526 B.n452 B.n11 585
R527 B.n454 B.n453 585
R528 B.n455 B.n10 585
R529 B.n457 B.n456 585
R530 B.n458 B.n9 585
R531 B.n460 B.n459 585
R532 B.n461 B.n8 585
R533 B.n463 B.n462 585
R534 B.n464 B.n7 585
R535 B.n466 B.n465 585
R536 B.n467 B.n6 585
R537 B.n469 B.n468 585
R538 B.n470 B.n5 585
R539 B.n472 B.n471 585
R540 B.n473 B.n4 585
R541 B.n475 B.n474 585
R542 B.n476 B.n3 585
R543 B.n478 B.n477 585
R544 B.n479 B.n0 585
R545 B.n2 B.n1 585
R546 B.n126 B.n125 585
R547 B.n128 B.n127 585
R548 B.n129 B.n124 585
R549 B.n131 B.n130 585
R550 B.n132 B.n123 585
R551 B.n134 B.n133 585
R552 B.n135 B.n122 585
R553 B.n137 B.n136 585
R554 B.n138 B.n121 585
R555 B.n140 B.n139 585
R556 B.n141 B.n120 585
R557 B.n143 B.n142 585
R558 B.n144 B.n119 585
R559 B.n146 B.n145 585
R560 B.n147 B.n118 585
R561 B.n149 B.n148 585
R562 B.n150 B.n117 585
R563 B.n152 B.n151 585
R564 B.n153 B.n116 585
R565 B.n155 B.n154 585
R566 B.n156 B.n115 585
R567 B.n158 B.n157 585
R568 B.n159 B.n114 585
R569 B.n161 B.n160 585
R570 B.n162 B.n113 585
R571 B.n164 B.n163 585
R572 B.n165 B.n112 585
R573 B.n167 B.n166 585
R574 B.n168 B.n111 585
R575 B.n170 B.n169 585
R576 B.n171 B.n110 585
R577 B.n173 B.n172 585
R578 B.n174 B.n173 550.159
R579 B.n251 B.n82 550.159
R580 B.n353 B.n48 550.159
R581 B.n431 B.n430 550.159
R582 B.n93 B.t10 303.69
R583 B.n37 B.t5 303.69
R584 B.n202 B.t1 303.69
R585 B.n30 B.t8 303.69
R586 B.n481 B.n480 256.663
R587 B.n202 B.t0 252.637
R588 B.n93 B.t9 252.637
R589 B.n37 B.t3 252.637
R590 B.n30 B.t6 252.637
R591 B.n94 B.t11 247.447
R592 B.n38 B.t4 247.447
R593 B.n203 B.t2 247.447
R594 B.n31 B.t7 247.447
R595 B.n480 B.n479 235.042
R596 B.n480 B.n2 235.042
R597 B.n175 B.n174 163.367
R598 B.n175 B.n108 163.367
R599 B.n179 B.n108 163.367
R600 B.n180 B.n179 163.367
R601 B.n181 B.n180 163.367
R602 B.n181 B.n106 163.367
R603 B.n185 B.n106 163.367
R604 B.n186 B.n185 163.367
R605 B.n187 B.n186 163.367
R606 B.n187 B.n104 163.367
R607 B.n191 B.n104 163.367
R608 B.n192 B.n191 163.367
R609 B.n193 B.n192 163.367
R610 B.n193 B.n102 163.367
R611 B.n197 B.n102 163.367
R612 B.n198 B.n197 163.367
R613 B.n199 B.n198 163.367
R614 B.n199 B.n100 163.367
R615 B.n206 B.n100 163.367
R616 B.n207 B.n206 163.367
R617 B.n208 B.n207 163.367
R618 B.n208 B.n98 163.367
R619 B.n212 B.n98 163.367
R620 B.n213 B.n212 163.367
R621 B.n214 B.n213 163.367
R622 B.n214 B.n96 163.367
R623 B.n218 B.n96 163.367
R624 B.n219 B.n218 163.367
R625 B.n220 B.n219 163.367
R626 B.n220 B.n92 163.367
R627 B.n225 B.n92 163.367
R628 B.n226 B.n225 163.367
R629 B.n227 B.n226 163.367
R630 B.n227 B.n90 163.367
R631 B.n231 B.n90 163.367
R632 B.n232 B.n231 163.367
R633 B.n233 B.n232 163.367
R634 B.n233 B.n88 163.367
R635 B.n237 B.n88 163.367
R636 B.n238 B.n237 163.367
R637 B.n239 B.n238 163.367
R638 B.n239 B.n86 163.367
R639 B.n243 B.n86 163.367
R640 B.n244 B.n243 163.367
R641 B.n245 B.n244 163.367
R642 B.n245 B.n84 163.367
R643 B.n249 B.n84 163.367
R644 B.n250 B.n249 163.367
R645 B.n251 B.n250 163.367
R646 B.n353 B.n352 163.367
R647 B.n352 B.n351 163.367
R648 B.n351 B.n50 163.367
R649 B.n347 B.n50 163.367
R650 B.n347 B.n346 163.367
R651 B.n346 B.n345 163.367
R652 B.n345 B.n52 163.367
R653 B.n341 B.n52 163.367
R654 B.n341 B.n340 163.367
R655 B.n340 B.n339 163.367
R656 B.n339 B.n54 163.367
R657 B.n335 B.n54 163.367
R658 B.n335 B.n334 163.367
R659 B.n334 B.n333 163.367
R660 B.n333 B.n56 163.367
R661 B.n329 B.n56 163.367
R662 B.n329 B.n328 163.367
R663 B.n328 B.n327 163.367
R664 B.n327 B.n58 163.367
R665 B.n323 B.n58 163.367
R666 B.n323 B.n322 163.367
R667 B.n322 B.n321 163.367
R668 B.n321 B.n60 163.367
R669 B.n317 B.n60 163.367
R670 B.n317 B.n316 163.367
R671 B.n316 B.n315 163.367
R672 B.n315 B.n62 163.367
R673 B.n311 B.n62 163.367
R674 B.n311 B.n310 163.367
R675 B.n310 B.n309 163.367
R676 B.n309 B.n64 163.367
R677 B.n305 B.n64 163.367
R678 B.n305 B.n304 163.367
R679 B.n304 B.n303 163.367
R680 B.n303 B.n66 163.367
R681 B.n299 B.n66 163.367
R682 B.n299 B.n298 163.367
R683 B.n298 B.n297 163.367
R684 B.n297 B.n68 163.367
R685 B.n293 B.n68 163.367
R686 B.n293 B.n292 163.367
R687 B.n292 B.n291 163.367
R688 B.n291 B.n70 163.367
R689 B.n287 B.n70 163.367
R690 B.n287 B.n286 163.367
R691 B.n286 B.n285 163.367
R692 B.n285 B.n72 163.367
R693 B.n281 B.n72 163.367
R694 B.n281 B.n280 163.367
R695 B.n280 B.n279 163.367
R696 B.n279 B.n74 163.367
R697 B.n275 B.n74 163.367
R698 B.n275 B.n274 163.367
R699 B.n274 B.n273 163.367
R700 B.n273 B.n76 163.367
R701 B.n269 B.n76 163.367
R702 B.n269 B.n268 163.367
R703 B.n268 B.n267 163.367
R704 B.n267 B.n78 163.367
R705 B.n263 B.n78 163.367
R706 B.n263 B.n262 163.367
R707 B.n262 B.n261 163.367
R708 B.n261 B.n80 163.367
R709 B.n257 B.n80 163.367
R710 B.n257 B.n256 163.367
R711 B.n256 B.n255 163.367
R712 B.n255 B.n82 163.367
R713 B.n430 B.n19 163.367
R714 B.n426 B.n19 163.367
R715 B.n426 B.n425 163.367
R716 B.n425 B.n424 163.367
R717 B.n424 B.n21 163.367
R718 B.n420 B.n21 163.367
R719 B.n420 B.n419 163.367
R720 B.n419 B.n418 163.367
R721 B.n418 B.n23 163.367
R722 B.n414 B.n23 163.367
R723 B.n414 B.n413 163.367
R724 B.n413 B.n412 163.367
R725 B.n412 B.n25 163.367
R726 B.n408 B.n25 163.367
R727 B.n408 B.n407 163.367
R728 B.n407 B.n406 163.367
R729 B.n406 B.n27 163.367
R730 B.n402 B.n27 163.367
R731 B.n402 B.n401 163.367
R732 B.n401 B.n400 163.367
R733 B.n400 B.n29 163.367
R734 B.n396 B.n29 163.367
R735 B.n396 B.n395 163.367
R736 B.n395 B.n394 163.367
R737 B.n394 B.n34 163.367
R738 B.n390 B.n34 163.367
R739 B.n390 B.n389 163.367
R740 B.n389 B.n388 163.367
R741 B.n388 B.n36 163.367
R742 B.n383 B.n36 163.367
R743 B.n383 B.n382 163.367
R744 B.n382 B.n381 163.367
R745 B.n381 B.n40 163.367
R746 B.n377 B.n40 163.367
R747 B.n377 B.n376 163.367
R748 B.n376 B.n375 163.367
R749 B.n375 B.n42 163.367
R750 B.n371 B.n42 163.367
R751 B.n371 B.n370 163.367
R752 B.n370 B.n369 163.367
R753 B.n369 B.n44 163.367
R754 B.n365 B.n44 163.367
R755 B.n365 B.n364 163.367
R756 B.n364 B.n363 163.367
R757 B.n363 B.n46 163.367
R758 B.n359 B.n46 163.367
R759 B.n359 B.n358 163.367
R760 B.n358 B.n357 163.367
R761 B.n357 B.n48 163.367
R762 B.n432 B.n431 163.367
R763 B.n432 B.n17 163.367
R764 B.n436 B.n17 163.367
R765 B.n437 B.n436 163.367
R766 B.n438 B.n437 163.367
R767 B.n438 B.n15 163.367
R768 B.n442 B.n15 163.367
R769 B.n443 B.n442 163.367
R770 B.n444 B.n443 163.367
R771 B.n444 B.n13 163.367
R772 B.n448 B.n13 163.367
R773 B.n449 B.n448 163.367
R774 B.n450 B.n449 163.367
R775 B.n450 B.n11 163.367
R776 B.n454 B.n11 163.367
R777 B.n455 B.n454 163.367
R778 B.n456 B.n455 163.367
R779 B.n456 B.n9 163.367
R780 B.n460 B.n9 163.367
R781 B.n461 B.n460 163.367
R782 B.n462 B.n461 163.367
R783 B.n462 B.n7 163.367
R784 B.n466 B.n7 163.367
R785 B.n467 B.n466 163.367
R786 B.n468 B.n467 163.367
R787 B.n468 B.n5 163.367
R788 B.n472 B.n5 163.367
R789 B.n473 B.n472 163.367
R790 B.n474 B.n473 163.367
R791 B.n474 B.n3 163.367
R792 B.n478 B.n3 163.367
R793 B.n479 B.n478 163.367
R794 B.n126 B.n2 163.367
R795 B.n127 B.n126 163.367
R796 B.n127 B.n124 163.367
R797 B.n131 B.n124 163.367
R798 B.n132 B.n131 163.367
R799 B.n133 B.n132 163.367
R800 B.n133 B.n122 163.367
R801 B.n137 B.n122 163.367
R802 B.n138 B.n137 163.367
R803 B.n139 B.n138 163.367
R804 B.n139 B.n120 163.367
R805 B.n143 B.n120 163.367
R806 B.n144 B.n143 163.367
R807 B.n145 B.n144 163.367
R808 B.n145 B.n118 163.367
R809 B.n149 B.n118 163.367
R810 B.n150 B.n149 163.367
R811 B.n151 B.n150 163.367
R812 B.n151 B.n116 163.367
R813 B.n155 B.n116 163.367
R814 B.n156 B.n155 163.367
R815 B.n157 B.n156 163.367
R816 B.n157 B.n114 163.367
R817 B.n161 B.n114 163.367
R818 B.n162 B.n161 163.367
R819 B.n163 B.n162 163.367
R820 B.n163 B.n112 163.367
R821 B.n167 B.n112 163.367
R822 B.n168 B.n167 163.367
R823 B.n169 B.n168 163.367
R824 B.n169 B.n110 163.367
R825 B.n173 B.n110 163.367
R826 B.n204 B.n203 59.5399
R827 B.n222 B.n94 59.5399
R828 B.n385 B.n38 59.5399
R829 B.n32 B.n31 59.5399
R830 B.n203 B.n202 56.2429
R831 B.n94 B.n93 56.2429
R832 B.n38 B.n37 56.2429
R833 B.n31 B.n30 56.2429
R834 B.n253 B.n252 35.7468
R835 B.n429 B.n18 35.7468
R836 B.n355 B.n354 35.7468
R837 B.n172 B.n109 35.7468
R838 B B.n481 18.0485
R839 B.n433 B.n18 10.6151
R840 B.n434 B.n433 10.6151
R841 B.n435 B.n434 10.6151
R842 B.n435 B.n16 10.6151
R843 B.n439 B.n16 10.6151
R844 B.n440 B.n439 10.6151
R845 B.n441 B.n440 10.6151
R846 B.n441 B.n14 10.6151
R847 B.n445 B.n14 10.6151
R848 B.n446 B.n445 10.6151
R849 B.n447 B.n446 10.6151
R850 B.n447 B.n12 10.6151
R851 B.n451 B.n12 10.6151
R852 B.n452 B.n451 10.6151
R853 B.n453 B.n452 10.6151
R854 B.n453 B.n10 10.6151
R855 B.n457 B.n10 10.6151
R856 B.n458 B.n457 10.6151
R857 B.n459 B.n458 10.6151
R858 B.n459 B.n8 10.6151
R859 B.n463 B.n8 10.6151
R860 B.n464 B.n463 10.6151
R861 B.n465 B.n464 10.6151
R862 B.n465 B.n6 10.6151
R863 B.n469 B.n6 10.6151
R864 B.n470 B.n469 10.6151
R865 B.n471 B.n470 10.6151
R866 B.n471 B.n4 10.6151
R867 B.n475 B.n4 10.6151
R868 B.n476 B.n475 10.6151
R869 B.n477 B.n476 10.6151
R870 B.n477 B.n0 10.6151
R871 B.n429 B.n428 10.6151
R872 B.n428 B.n427 10.6151
R873 B.n427 B.n20 10.6151
R874 B.n423 B.n20 10.6151
R875 B.n423 B.n422 10.6151
R876 B.n422 B.n421 10.6151
R877 B.n421 B.n22 10.6151
R878 B.n417 B.n22 10.6151
R879 B.n417 B.n416 10.6151
R880 B.n416 B.n415 10.6151
R881 B.n415 B.n24 10.6151
R882 B.n411 B.n24 10.6151
R883 B.n411 B.n410 10.6151
R884 B.n410 B.n409 10.6151
R885 B.n409 B.n26 10.6151
R886 B.n405 B.n26 10.6151
R887 B.n405 B.n404 10.6151
R888 B.n404 B.n403 10.6151
R889 B.n403 B.n28 10.6151
R890 B.n399 B.n398 10.6151
R891 B.n398 B.n397 10.6151
R892 B.n397 B.n33 10.6151
R893 B.n393 B.n33 10.6151
R894 B.n393 B.n392 10.6151
R895 B.n392 B.n391 10.6151
R896 B.n391 B.n35 10.6151
R897 B.n387 B.n35 10.6151
R898 B.n387 B.n386 10.6151
R899 B.n384 B.n39 10.6151
R900 B.n380 B.n39 10.6151
R901 B.n380 B.n379 10.6151
R902 B.n379 B.n378 10.6151
R903 B.n378 B.n41 10.6151
R904 B.n374 B.n41 10.6151
R905 B.n374 B.n373 10.6151
R906 B.n373 B.n372 10.6151
R907 B.n372 B.n43 10.6151
R908 B.n368 B.n43 10.6151
R909 B.n368 B.n367 10.6151
R910 B.n367 B.n366 10.6151
R911 B.n366 B.n45 10.6151
R912 B.n362 B.n45 10.6151
R913 B.n362 B.n361 10.6151
R914 B.n361 B.n360 10.6151
R915 B.n360 B.n47 10.6151
R916 B.n356 B.n47 10.6151
R917 B.n356 B.n355 10.6151
R918 B.n354 B.n49 10.6151
R919 B.n350 B.n49 10.6151
R920 B.n350 B.n349 10.6151
R921 B.n349 B.n348 10.6151
R922 B.n348 B.n51 10.6151
R923 B.n344 B.n51 10.6151
R924 B.n344 B.n343 10.6151
R925 B.n343 B.n342 10.6151
R926 B.n342 B.n53 10.6151
R927 B.n338 B.n53 10.6151
R928 B.n338 B.n337 10.6151
R929 B.n337 B.n336 10.6151
R930 B.n336 B.n55 10.6151
R931 B.n332 B.n55 10.6151
R932 B.n332 B.n331 10.6151
R933 B.n331 B.n330 10.6151
R934 B.n330 B.n57 10.6151
R935 B.n326 B.n57 10.6151
R936 B.n326 B.n325 10.6151
R937 B.n325 B.n324 10.6151
R938 B.n324 B.n59 10.6151
R939 B.n320 B.n59 10.6151
R940 B.n320 B.n319 10.6151
R941 B.n319 B.n318 10.6151
R942 B.n318 B.n61 10.6151
R943 B.n314 B.n61 10.6151
R944 B.n314 B.n313 10.6151
R945 B.n313 B.n312 10.6151
R946 B.n312 B.n63 10.6151
R947 B.n308 B.n63 10.6151
R948 B.n308 B.n307 10.6151
R949 B.n307 B.n306 10.6151
R950 B.n306 B.n65 10.6151
R951 B.n302 B.n65 10.6151
R952 B.n302 B.n301 10.6151
R953 B.n301 B.n300 10.6151
R954 B.n300 B.n67 10.6151
R955 B.n296 B.n67 10.6151
R956 B.n296 B.n295 10.6151
R957 B.n295 B.n294 10.6151
R958 B.n294 B.n69 10.6151
R959 B.n290 B.n69 10.6151
R960 B.n290 B.n289 10.6151
R961 B.n289 B.n288 10.6151
R962 B.n288 B.n71 10.6151
R963 B.n284 B.n71 10.6151
R964 B.n284 B.n283 10.6151
R965 B.n283 B.n282 10.6151
R966 B.n282 B.n73 10.6151
R967 B.n278 B.n73 10.6151
R968 B.n278 B.n277 10.6151
R969 B.n277 B.n276 10.6151
R970 B.n276 B.n75 10.6151
R971 B.n272 B.n75 10.6151
R972 B.n272 B.n271 10.6151
R973 B.n271 B.n270 10.6151
R974 B.n270 B.n77 10.6151
R975 B.n266 B.n77 10.6151
R976 B.n266 B.n265 10.6151
R977 B.n265 B.n264 10.6151
R978 B.n264 B.n79 10.6151
R979 B.n260 B.n79 10.6151
R980 B.n260 B.n259 10.6151
R981 B.n259 B.n258 10.6151
R982 B.n258 B.n81 10.6151
R983 B.n254 B.n81 10.6151
R984 B.n254 B.n253 10.6151
R985 B.n125 B.n1 10.6151
R986 B.n128 B.n125 10.6151
R987 B.n129 B.n128 10.6151
R988 B.n130 B.n129 10.6151
R989 B.n130 B.n123 10.6151
R990 B.n134 B.n123 10.6151
R991 B.n135 B.n134 10.6151
R992 B.n136 B.n135 10.6151
R993 B.n136 B.n121 10.6151
R994 B.n140 B.n121 10.6151
R995 B.n141 B.n140 10.6151
R996 B.n142 B.n141 10.6151
R997 B.n142 B.n119 10.6151
R998 B.n146 B.n119 10.6151
R999 B.n147 B.n146 10.6151
R1000 B.n148 B.n147 10.6151
R1001 B.n148 B.n117 10.6151
R1002 B.n152 B.n117 10.6151
R1003 B.n153 B.n152 10.6151
R1004 B.n154 B.n153 10.6151
R1005 B.n154 B.n115 10.6151
R1006 B.n158 B.n115 10.6151
R1007 B.n159 B.n158 10.6151
R1008 B.n160 B.n159 10.6151
R1009 B.n160 B.n113 10.6151
R1010 B.n164 B.n113 10.6151
R1011 B.n165 B.n164 10.6151
R1012 B.n166 B.n165 10.6151
R1013 B.n166 B.n111 10.6151
R1014 B.n170 B.n111 10.6151
R1015 B.n171 B.n170 10.6151
R1016 B.n172 B.n171 10.6151
R1017 B.n176 B.n109 10.6151
R1018 B.n177 B.n176 10.6151
R1019 B.n178 B.n177 10.6151
R1020 B.n178 B.n107 10.6151
R1021 B.n182 B.n107 10.6151
R1022 B.n183 B.n182 10.6151
R1023 B.n184 B.n183 10.6151
R1024 B.n184 B.n105 10.6151
R1025 B.n188 B.n105 10.6151
R1026 B.n189 B.n188 10.6151
R1027 B.n190 B.n189 10.6151
R1028 B.n190 B.n103 10.6151
R1029 B.n194 B.n103 10.6151
R1030 B.n195 B.n194 10.6151
R1031 B.n196 B.n195 10.6151
R1032 B.n196 B.n101 10.6151
R1033 B.n200 B.n101 10.6151
R1034 B.n201 B.n200 10.6151
R1035 B.n205 B.n201 10.6151
R1036 B.n209 B.n99 10.6151
R1037 B.n210 B.n209 10.6151
R1038 B.n211 B.n210 10.6151
R1039 B.n211 B.n97 10.6151
R1040 B.n215 B.n97 10.6151
R1041 B.n216 B.n215 10.6151
R1042 B.n217 B.n216 10.6151
R1043 B.n217 B.n95 10.6151
R1044 B.n221 B.n95 10.6151
R1045 B.n224 B.n223 10.6151
R1046 B.n224 B.n91 10.6151
R1047 B.n228 B.n91 10.6151
R1048 B.n229 B.n228 10.6151
R1049 B.n230 B.n229 10.6151
R1050 B.n230 B.n89 10.6151
R1051 B.n234 B.n89 10.6151
R1052 B.n235 B.n234 10.6151
R1053 B.n236 B.n235 10.6151
R1054 B.n236 B.n87 10.6151
R1055 B.n240 B.n87 10.6151
R1056 B.n241 B.n240 10.6151
R1057 B.n242 B.n241 10.6151
R1058 B.n242 B.n85 10.6151
R1059 B.n246 B.n85 10.6151
R1060 B.n247 B.n246 10.6151
R1061 B.n248 B.n247 10.6151
R1062 B.n248 B.n83 10.6151
R1063 B.n252 B.n83 10.6151
R1064 B.n32 B.n28 9.36635
R1065 B.n385 B.n384 9.36635
R1066 B.n205 B.n204 9.36635
R1067 B.n223 B.n222 9.36635
R1068 B.n481 B.n0 8.11757
R1069 B.n481 B.n1 8.11757
R1070 B.n399 B.n32 1.24928
R1071 B.n386 B.n385 1.24928
R1072 B.n204 B.n99 1.24928
R1073 B.n222 B.n221 1.24928
C0 VP VDD2 0.397113f
C1 VP B 1.6086f
C2 VP VTAIL 2.44276f
C3 VN w_n2710_n1920# 4.44082f
C4 VDD2 VN 2.0713f
C5 B VN 1.03083f
C6 VN VTAIL 2.42865f
C7 VDD1 w_n2710_n1920# 1.25529f
C8 VP VN 4.8239f
C9 VDD1 VDD2 1.0153f
C10 B VDD1 1.06038f
C11 VDD1 VTAIL 3.67297f
C12 VP VDD1 2.31393f
C13 VDD2 w_n2710_n1920# 1.31043f
C14 B w_n2710_n1920# 7.19242f
C15 VTAIL w_n2710_n1920# 2.33374f
C16 VDD1 VN 0.15331f
C17 B VDD2 1.11213f
C18 VDD2 VTAIL 3.72698f
C19 B VTAIL 2.53657f
C20 VP w_n2710_n1920# 4.78903f
C21 VDD2 VSUBS 0.772283f
C22 VDD1 VSUBS 4.796306f
C23 VTAIL VSUBS 0.647217f
C24 VN VSUBS 5.30658f
C25 VP VSUBS 1.853972f
C26 B VSUBS 3.450163f
C27 w_n2710_n1920# VSUBS 65.2676f
C28 B.n0 VSUBS 0.007804f
C29 B.n1 VSUBS 0.007804f
C30 B.n2 VSUBS 0.011542f
C31 B.n3 VSUBS 0.008845f
C32 B.n4 VSUBS 0.008845f
C33 B.n5 VSUBS 0.008845f
C34 B.n6 VSUBS 0.008845f
C35 B.n7 VSUBS 0.008845f
C36 B.n8 VSUBS 0.008845f
C37 B.n9 VSUBS 0.008845f
C38 B.n10 VSUBS 0.008845f
C39 B.n11 VSUBS 0.008845f
C40 B.n12 VSUBS 0.008845f
C41 B.n13 VSUBS 0.008845f
C42 B.n14 VSUBS 0.008845f
C43 B.n15 VSUBS 0.008845f
C44 B.n16 VSUBS 0.008845f
C45 B.n17 VSUBS 0.008845f
C46 B.n18 VSUBS 0.021458f
C47 B.n19 VSUBS 0.008845f
C48 B.n20 VSUBS 0.008845f
C49 B.n21 VSUBS 0.008845f
C50 B.n22 VSUBS 0.008845f
C51 B.n23 VSUBS 0.008845f
C52 B.n24 VSUBS 0.008845f
C53 B.n25 VSUBS 0.008845f
C54 B.n26 VSUBS 0.008845f
C55 B.n27 VSUBS 0.008845f
C56 B.n28 VSUBS 0.008325f
C57 B.n29 VSUBS 0.008845f
C58 B.t7 VSUBS 0.087738f
C59 B.t8 VSUBS 0.116182f
C60 B.t6 VSUBS 0.738238f
C61 B.n30 VSUBS 0.200364f
C62 B.n31 VSUBS 0.166201f
C63 B.n32 VSUBS 0.020493f
C64 B.n33 VSUBS 0.008845f
C65 B.n34 VSUBS 0.008845f
C66 B.n35 VSUBS 0.008845f
C67 B.n36 VSUBS 0.008845f
C68 B.t4 VSUBS 0.08774f
C69 B.t5 VSUBS 0.116183f
C70 B.t3 VSUBS 0.738238f
C71 B.n37 VSUBS 0.200363f
C72 B.n38 VSUBS 0.166199f
C73 B.n39 VSUBS 0.008845f
C74 B.n40 VSUBS 0.008845f
C75 B.n41 VSUBS 0.008845f
C76 B.n42 VSUBS 0.008845f
C77 B.n43 VSUBS 0.008845f
C78 B.n44 VSUBS 0.008845f
C79 B.n45 VSUBS 0.008845f
C80 B.n46 VSUBS 0.008845f
C81 B.n47 VSUBS 0.008845f
C82 B.n48 VSUBS 0.022506f
C83 B.n49 VSUBS 0.008845f
C84 B.n50 VSUBS 0.008845f
C85 B.n51 VSUBS 0.008845f
C86 B.n52 VSUBS 0.008845f
C87 B.n53 VSUBS 0.008845f
C88 B.n54 VSUBS 0.008845f
C89 B.n55 VSUBS 0.008845f
C90 B.n56 VSUBS 0.008845f
C91 B.n57 VSUBS 0.008845f
C92 B.n58 VSUBS 0.008845f
C93 B.n59 VSUBS 0.008845f
C94 B.n60 VSUBS 0.008845f
C95 B.n61 VSUBS 0.008845f
C96 B.n62 VSUBS 0.008845f
C97 B.n63 VSUBS 0.008845f
C98 B.n64 VSUBS 0.008845f
C99 B.n65 VSUBS 0.008845f
C100 B.n66 VSUBS 0.008845f
C101 B.n67 VSUBS 0.008845f
C102 B.n68 VSUBS 0.008845f
C103 B.n69 VSUBS 0.008845f
C104 B.n70 VSUBS 0.008845f
C105 B.n71 VSUBS 0.008845f
C106 B.n72 VSUBS 0.008845f
C107 B.n73 VSUBS 0.008845f
C108 B.n74 VSUBS 0.008845f
C109 B.n75 VSUBS 0.008845f
C110 B.n76 VSUBS 0.008845f
C111 B.n77 VSUBS 0.008845f
C112 B.n78 VSUBS 0.008845f
C113 B.n79 VSUBS 0.008845f
C114 B.n80 VSUBS 0.008845f
C115 B.n81 VSUBS 0.008845f
C116 B.n82 VSUBS 0.021458f
C117 B.n83 VSUBS 0.008845f
C118 B.n84 VSUBS 0.008845f
C119 B.n85 VSUBS 0.008845f
C120 B.n86 VSUBS 0.008845f
C121 B.n87 VSUBS 0.008845f
C122 B.n88 VSUBS 0.008845f
C123 B.n89 VSUBS 0.008845f
C124 B.n90 VSUBS 0.008845f
C125 B.n91 VSUBS 0.008845f
C126 B.n92 VSUBS 0.008845f
C127 B.t11 VSUBS 0.08774f
C128 B.t10 VSUBS 0.116183f
C129 B.t9 VSUBS 0.738238f
C130 B.n93 VSUBS 0.200363f
C131 B.n94 VSUBS 0.166199f
C132 B.n95 VSUBS 0.008845f
C133 B.n96 VSUBS 0.008845f
C134 B.n97 VSUBS 0.008845f
C135 B.n98 VSUBS 0.008845f
C136 B.n99 VSUBS 0.004943f
C137 B.n100 VSUBS 0.008845f
C138 B.n101 VSUBS 0.008845f
C139 B.n102 VSUBS 0.008845f
C140 B.n103 VSUBS 0.008845f
C141 B.n104 VSUBS 0.008845f
C142 B.n105 VSUBS 0.008845f
C143 B.n106 VSUBS 0.008845f
C144 B.n107 VSUBS 0.008845f
C145 B.n108 VSUBS 0.008845f
C146 B.n109 VSUBS 0.022506f
C147 B.n110 VSUBS 0.008845f
C148 B.n111 VSUBS 0.008845f
C149 B.n112 VSUBS 0.008845f
C150 B.n113 VSUBS 0.008845f
C151 B.n114 VSUBS 0.008845f
C152 B.n115 VSUBS 0.008845f
C153 B.n116 VSUBS 0.008845f
C154 B.n117 VSUBS 0.008845f
C155 B.n118 VSUBS 0.008845f
C156 B.n119 VSUBS 0.008845f
C157 B.n120 VSUBS 0.008845f
C158 B.n121 VSUBS 0.008845f
C159 B.n122 VSUBS 0.008845f
C160 B.n123 VSUBS 0.008845f
C161 B.n124 VSUBS 0.008845f
C162 B.n125 VSUBS 0.008845f
C163 B.n126 VSUBS 0.008845f
C164 B.n127 VSUBS 0.008845f
C165 B.n128 VSUBS 0.008845f
C166 B.n129 VSUBS 0.008845f
C167 B.n130 VSUBS 0.008845f
C168 B.n131 VSUBS 0.008845f
C169 B.n132 VSUBS 0.008845f
C170 B.n133 VSUBS 0.008845f
C171 B.n134 VSUBS 0.008845f
C172 B.n135 VSUBS 0.008845f
C173 B.n136 VSUBS 0.008845f
C174 B.n137 VSUBS 0.008845f
C175 B.n138 VSUBS 0.008845f
C176 B.n139 VSUBS 0.008845f
C177 B.n140 VSUBS 0.008845f
C178 B.n141 VSUBS 0.008845f
C179 B.n142 VSUBS 0.008845f
C180 B.n143 VSUBS 0.008845f
C181 B.n144 VSUBS 0.008845f
C182 B.n145 VSUBS 0.008845f
C183 B.n146 VSUBS 0.008845f
C184 B.n147 VSUBS 0.008845f
C185 B.n148 VSUBS 0.008845f
C186 B.n149 VSUBS 0.008845f
C187 B.n150 VSUBS 0.008845f
C188 B.n151 VSUBS 0.008845f
C189 B.n152 VSUBS 0.008845f
C190 B.n153 VSUBS 0.008845f
C191 B.n154 VSUBS 0.008845f
C192 B.n155 VSUBS 0.008845f
C193 B.n156 VSUBS 0.008845f
C194 B.n157 VSUBS 0.008845f
C195 B.n158 VSUBS 0.008845f
C196 B.n159 VSUBS 0.008845f
C197 B.n160 VSUBS 0.008845f
C198 B.n161 VSUBS 0.008845f
C199 B.n162 VSUBS 0.008845f
C200 B.n163 VSUBS 0.008845f
C201 B.n164 VSUBS 0.008845f
C202 B.n165 VSUBS 0.008845f
C203 B.n166 VSUBS 0.008845f
C204 B.n167 VSUBS 0.008845f
C205 B.n168 VSUBS 0.008845f
C206 B.n169 VSUBS 0.008845f
C207 B.n170 VSUBS 0.008845f
C208 B.n171 VSUBS 0.008845f
C209 B.n172 VSUBS 0.021458f
C210 B.n173 VSUBS 0.021458f
C211 B.n174 VSUBS 0.022506f
C212 B.n175 VSUBS 0.008845f
C213 B.n176 VSUBS 0.008845f
C214 B.n177 VSUBS 0.008845f
C215 B.n178 VSUBS 0.008845f
C216 B.n179 VSUBS 0.008845f
C217 B.n180 VSUBS 0.008845f
C218 B.n181 VSUBS 0.008845f
C219 B.n182 VSUBS 0.008845f
C220 B.n183 VSUBS 0.008845f
C221 B.n184 VSUBS 0.008845f
C222 B.n185 VSUBS 0.008845f
C223 B.n186 VSUBS 0.008845f
C224 B.n187 VSUBS 0.008845f
C225 B.n188 VSUBS 0.008845f
C226 B.n189 VSUBS 0.008845f
C227 B.n190 VSUBS 0.008845f
C228 B.n191 VSUBS 0.008845f
C229 B.n192 VSUBS 0.008845f
C230 B.n193 VSUBS 0.008845f
C231 B.n194 VSUBS 0.008845f
C232 B.n195 VSUBS 0.008845f
C233 B.n196 VSUBS 0.008845f
C234 B.n197 VSUBS 0.008845f
C235 B.n198 VSUBS 0.008845f
C236 B.n199 VSUBS 0.008845f
C237 B.n200 VSUBS 0.008845f
C238 B.n201 VSUBS 0.008845f
C239 B.t2 VSUBS 0.087738f
C240 B.t1 VSUBS 0.116182f
C241 B.t0 VSUBS 0.738238f
C242 B.n202 VSUBS 0.200364f
C243 B.n203 VSUBS 0.166201f
C244 B.n204 VSUBS 0.020493f
C245 B.n205 VSUBS 0.008325f
C246 B.n206 VSUBS 0.008845f
C247 B.n207 VSUBS 0.008845f
C248 B.n208 VSUBS 0.008845f
C249 B.n209 VSUBS 0.008845f
C250 B.n210 VSUBS 0.008845f
C251 B.n211 VSUBS 0.008845f
C252 B.n212 VSUBS 0.008845f
C253 B.n213 VSUBS 0.008845f
C254 B.n214 VSUBS 0.008845f
C255 B.n215 VSUBS 0.008845f
C256 B.n216 VSUBS 0.008845f
C257 B.n217 VSUBS 0.008845f
C258 B.n218 VSUBS 0.008845f
C259 B.n219 VSUBS 0.008845f
C260 B.n220 VSUBS 0.008845f
C261 B.n221 VSUBS 0.004943f
C262 B.n222 VSUBS 0.020493f
C263 B.n223 VSUBS 0.008325f
C264 B.n224 VSUBS 0.008845f
C265 B.n225 VSUBS 0.008845f
C266 B.n226 VSUBS 0.008845f
C267 B.n227 VSUBS 0.008845f
C268 B.n228 VSUBS 0.008845f
C269 B.n229 VSUBS 0.008845f
C270 B.n230 VSUBS 0.008845f
C271 B.n231 VSUBS 0.008845f
C272 B.n232 VSUBS 0.008845f
C273 B.n233 VSUBS 0.008845f
C274 B.n234 VSUBS 0.008845f
C275 B.n235 VSUBS 0.008845f
C276 B.n236 VSUBS 0.008845f
C277 B.n237 VSUBS 0.008845f
C278 B.n238 VSUBS 0.008845f
C279 B.n239 VSUBS 0.008845f
C280 B.n240 VSUBS 0.008845f
C281 B.n241 VSUBS 0.008845f
C282 B.n242 VSUBS 0.008845f
C283 B.n243 VSUBS 0.008845f
C284 B.n244 VSUBS 0.008845f
C285 B.n245 VSUBS 0.008845f
C286 B.n246 VSUBS 0.008845f
C287 B.n247 VSUBS 0.008845f
C288 B.n248 VSUBS 0.008845f
C289 B.n249 VSUBS 0.008845f
C290 B.n250 VSUBS 0.008845f
C291 B.n251 VSUBS 0.022506f
C292 B.n252 VSUBS 0.021551f
C293 B.n253 VSUBS 0.022413f
C294 B.n254 VSUBS 0.008845f
C295 B.n255 VSUBS 0.008845f
C296 B.n256 VSUBS 0.008845f
C297 B.n257 VSUBS 0.008845f
C298 B.n258 VSUBS 0.008845f
C299 B.n259 VSUBS 0.008845f
C300 B.n260 VSUBS 0.008845f
C301 B.n261 VSUBS 0.008845f
C302 B.n262 VSUBS 0.008845f
C303 B.n263 VSUBS 0.008845f
C304 B.n264 VSUBS 0.008845f
C305 B.n265 VSUBS 0.008845f
C306 B.n266 VSUBS 0.008845f
C307 B.n267 VSUBS 0.008845f
C308 B.n268 VSUBS 0.008845f
C309 B.n269 VSUBS 0.008845f
C310 B.n270 VSUBS 0.008845f
C311 B.n271 VSUBS 0.008845f
C312 B.n272 VSUBS 0.008845f
C313 B.n273 VSUBS 0.008845f
C314 B.n274 VSUBS 0.008845f
C315 B.n275 VSUBS 0.008845f
C316 B.n276 VSUBS 0.008845f
C317 B.n277 VSUBS 0.008845f
C318 B.n278 VSUBS 0.008845f
C319 B.n279 VSUBS 0.008845f
C320 B.n280 VSUBS 0.008845f
C321 B.n281 VSUBS 0.008845f
C322 B.n282 VSUBS 0.008845f
C323 B.n283 VSUBS 0.008845f
C324 B.n284 VSUBS 0.008845f
C325 B.n285 VSUBS 0.008845f
C326 B.n286 VSUBS 0.008845f
C327 B.n287 VSUBS 0.008845f
C328 B.n288 VSUBS 0.008845f
C329 B.n289 VSUBS 0.008845f
C330 B.n290 VSUBS 0.008845f
C331 B.n291 VSUBS 0.008845f
C332 B.n292 VSUBS 0.008845f
C333 B.n293 VSUBS 0.008845f
C334 B.n294 VSUBS 0.008845f
C335 B.n295 VSUBS 0.008845f
C336 B.n296 VSUBS 0.008845f
C337 B.n297 VSUBS 0.008845f
C338 B.n298 VSUBS 0.008845f
C339 B.n299 VSUBS 0.008845f
C340 B.n300 VSUBS 0.008845f
C341 B.n301 VSUBS 0.008845f
C342 B.n302 VSUBS 0.008845f
C343 B.n303 VSUBS 0.008845f
C344 B.n304 VSUBS 0.008845f
C345 B.n305 VSUBS 0.008845f
C346 B.n306 VSUBS 0.008845f
C347 B.n307 VSUBS 0.008845f
C348 B.n308 VSUBS 0.008845f
C349 B.n309 VSUBS 0.008845f
C350 B.n310 VSUBS 0.008845f
C351 B.n311 VSUBS 0.008845f
C352 B.n312 VSUBS 0.008845f
C353 B.n313 VSUBS 0.008845f
C354 B.n314 VSUBS 0.008845f
C355 B.n315 VSUBS 0.008845f
C356 B.n316 VSUBS 0.008845f
C357 B.n317 VSUBS 0.008845f
C358 B.n318 VSUBS 0.008845f
C359 B.n319 VSUBS 0.008845f
C360 B.n320 VSUBS 0.008845f
C361 B.n321 VSUBS 0.008845f
C362 B.n322 VSUBS 0.008845f
C363 B.n323 VSUBS 0.008845f
C364 B.n324 VSUBS 0.008845f
C365 B.n325 VSUBS 0.008845f
C366 B.n326 VSUBS 0.008845f
C367 B.n327 VSUBS 0.008845f
C368 B.n328 VSUBS 0.008845f
C369 B.n329 VSUBS 0.008845f
C370 B.n330 VSUBS 0.008845f
C371 B.n331 VSUBS 0.008845f
C372 B.n332 VSUBS 0.008845f
C373 B.n333 VSUBS 0.008845f
C374 B.n334 VSUBS 0.008845f
C375 B.n335 VSUBS 0.008845f
C376 B.n336 VSUBS 0.008845f
C377 B.n337 VSUBS 0.008845f
C378 B.n338 VSUBS 0.008845f
C379 B.n339 VSUBS 0.008845f
C380 B.n340 VSUBS 0.008845f
C381 B.n341 VSUBS 0.008845f
C382 B.n342 VSUBS 0.008845f
C383 B.n343 VSUBS 0.008845f
C384 B.n344 VSUBS 0.008845f
C385 B.n345 VSUBS 0.008845f
C386 B.n346 VSUBS 0.008845f
C387 B.n347 VSUBS 0.008845f
C388 B.n348 VSUBS 0.008845f
C389 B.n349 VSUBS 0.008845f
C390 B.n350 VSUBS 0.008845f
C391 B.n351 VSUBS 0.008845f
C392 B.n352 VSUBS 0.008845f
C393 B.n353 VSUBS 0.021458f
C394 B.n354 VSUBS 0.021458f
C395 B.n355 VSUBS 0.022506f
C396 B.n356 VSUBS 0.008845f
C397 B.n357 VSUBS 0.008845f
C398 B.n358 VSUBS 0.008845f
C399 B.n359 VSUBS 0.008845f
C400 B.n360 VSUBS 0.008845f
C401 B.n361 VSUBS 0.008845f
C402 B.n362 VSUBS 0.008845f
C403 B.n363 VSUBS 0.008845f
C404 B.n364 VSUBS 0.008845f
C405 B.n365 VSUBS 0.008845f
C406 B.n366 VSUBS 0.008845f
C407 B.n367 VSUBS 0.008845f
C408 B.n368 VSUBS 0.008845f
C409 B.n369 VSUBS 0.008845f
C410 B.n370 VSUBS 0.008845f
C411 B.n371 VSUBS 0.008845f
C412 B.n372 VSUBS 0.008845f
C413 B.n373 VSUBS 0.008845f
C414 B.n374 VSUBS 0.008845f
C415 B.n375 VSUBS 0.008845f
C416 B.n376 VSUBS 0.008845f
C417 B.n377 VSUBS 0.008845f
C418 B.n378 VSUBS 0.008845f
C419 B.n379 VSUBS 0.008845f
C420 B.n380 VSUBS 0.008845f
C421 B.n381 VSUBS 0.008845f
C422 B.n382 VSUBS 0.008845f
C423 B.n383 VSUBS 0.008845f
C424 B.n384 VSUBS 0.008325f
C425 B.n385 VSUBS 0.020493f
C426 B.n386 VSUBS 0.004943f
C427 B.n387 VSUBS 0.008845f
C428 B.n388 VSUBS 0.008845f
C429 B.n389 VSUBS 0.008845f
C430 B.n390 VSUBS 0.008845f
C431 B.n391 VSUBS 0.008845f
C432 B.n392 VSUBS 0.008845f
C433 B.n393 VSUBS 0.008845f
C434 B.n394 VSUBS 0.008845f
C435 B.n395 VSUBS 0.008845f
C436 B.n396 VSUBS 0.008845f
C437 B.n397 VSUBS 0.008845f
C438 B.n398 VSUBS 0.008845f
C439 B.n399 VSUBS 0.004943f
C440 B.n400 VSUBS 0.008845f
C441 B.n401 VSUBS 0.008845f
C442 B.n402 VSUBS 0.008845f
C443 B.n403 VSUBS 0.008845f
C444 B.n404 VSUBS 0.008845f
C445 B.n405 VSUBS 0.008845f
C446 B.n406 VSUBS 0.008845f
C447 B.n407 VSUBS 0.008845f
C448 B.n408 VSUBS 0.008845f
C449 B.n409 VSUBS 0.008845f
C450 B.n410 VSUBS 0.008845f
C451 B.n411 VSUBS 0.008845f
C452 B.n412 VSUBS 0.008845f
C453 B.n413 VSUBS 0.008845f
C454 B.n414 VSUBS 0.008845f
C455 B.n415 VSUBS 0.008845f
C456 B.n416 VSUBS 0.008845f
C457 B.n417 VSUBS 0.008845f
C458 B.n418 VSUBS 0.008845f
C459 B.n419 VSUBS 0.008845f
C460 B.n420 VSUBS 0.008845f
C461 B.n421 VSUBS 0.008845f
C462 B.n422 VSUBS 0.008845f
C463 B.n423 VSUBS 0.008845f
C464 B.n424 VSUBS 0.008845f
C465 B.n425 VSUBS 0.008845f
C466 B.n426 VSUBS 0.008845f
C467 B.n427 VSUBS 0.008845f
C468 B.n428 VSUBS 0.008845f
C469 B.n429 VSUBS 0.022506f
C470 B.n430 VSUBS 0.022506f
C471 B.n431 VSUBS 0.021458f
C472 B.n432 VSUBS 0.008845f
C473 B.n433 VSUBS 0.008845f
C474 B.n434 VSUBS 0.008845f
C475 B.n435 VSUBS 0.008845f
C476 B.n436 VSUBS 0.008845f
C477 B.n437 VSUBS 0.008845f
C478 B.n438 VSUBS 0.008845f
C479 B.n439 VSUBS 0.008845f
C480 B.n440 VSUBS 0.008845f
C481 B.n441 VSUBS 0.008845f
C482 B.n442 VSUBS 0.008845f
C483 B.n443 VSUBS 0.008845f
C484 B.n444 VSUBS 0.008845f
C485 B.n445 VSUBS 0.008845f
C486 B.n446 VSUBS 0.008845f
C487 B.n447 VSUBS 0.008845f
C488 B.n448 VSUBS 0.008845f
C489 B.n449 VSUBS 0.008845f
C490 B.n450 VSUBS 0.008845f
C491 B.n451 VSUBS 0.008845f
C492 B.n452 VSUBS 0.008845f
C493 B.n453 VSUBS 0.008845f
C494 B.n454 VSUBS 0.008845f
C495 B.n455 VSUBS 0.008845f
C496 B.n456 VSUBS 0.008845f
C497 B.n457 VSUBS 0.008845f
C498 B.n458 VSUBS 0.008845f
C499 B.n459 VSUBS 0.008845f
C500 B.n460 VSUBS 0.008845f
C501 B.n461 VSUBS 0.008845f
C502 B.n462 VSUBS 0.008845f
C503 B.n463 VSUBS 0.008845f
C504 B.n464 VSUBS 0.008845f
C505 B.n465 VSUBS 0.008845f
C506 B.n466 VSUBS 0.008845f
C507 B.n467 VSUBS 0.008845f
C508 B.n468 VSUBS 0.008845f
C509 B.n469 VSUBS 0.008845f
C510 B.n470 VSUBS 0.008845f
C511 B.n471 VSUBS 0.008845f
C512 B.n472 VSUBS 0.008845f
C513 B.n473 VSUBS 0.008845f
C514 B.n474 VSUBS 0.008845f
C515 B.n475 VSUBS 0.008845f
C516 B.n476 VSUBS 0.008845f
C517 B.n477 VSUBS 0.008845f
C518 B.n478 VSUBS 0.008845f
C519 B.n479 VSUBS 0.011542f
C520 B.n480 VSUBS 0.012295f
C521 B.n481 VSUBS 0.02445f
C522 VDD2.t0 VSUBS 0.104839f
C523 VDD2.t1 VSUBS 0.104839f
C524 VDD2.n0 VSUBS 1.00307f
C525 VDD2.t3 VSUBS 0.104839f
C526 VDD2.t2 VSUBS 0.104839f
C527 VDD2.n1 VSUBS 0.650516f
C528 VDD2.n2 VSUBS 3.49654f
C529 VN.t3 VSUBS 1.77163f
C530 VN.t2 VSUBS 1.76397f
C531 VN.n0 VSUBS 1.09927f
C532 VN.t1 VSUBS 1.77163f
C533 VN.t0 VSUBS 1.76397f
C534 VN.n1 VSUBS 3.08335f
C535 VTAIL.n0 VSUBS 0.033127f
C536 VTAIL.n1 VSUBS 0.02892f
C537 VTAIL.n2 VSUBS 0.01554f
C538 VTAIL.n3 VSUBS 0.036732f
C539 VTAIL.n4 VSUBS 0.016454f
C540 VTAIL.n5 VSUBS 0.49709f
C541 VTAIL.n6 VSUBS 0.01554f
C542 VTAIL.t2 VSUBS 0.080673f
C543 VTAIL.n7 VSUBS 0.118949f
C544 VTAIL.n8 VSUBS 0.02327f
C545 VTAIL.n9 VSUBS 0.027549f
C546 VTAIL.n10 VSUBS 0.036732f
C547 VTAIL.n11 VSUBS 0.016454f
C548 VTAIL.n12 VSUBS 0.01554f
C549 VTAIL.n13 VSUBS 0.02892f
C550 VTAIL.n14 VSUBS 0.02892f
C551 VTAIL.n15 VSUBS 0.01554f
C552 VTAIL.n16 VSUBS 0.016454f
C553 VTAIL.n17 VSUBS 0.036732f
C554 VTAIL.n18 VSUBS 0.093523f
C555 VTAIL.n19 VSUBS 0.016454f
C556 VTAIL.n20 VSUBS 0.01554f
C557 VTAIL.n21 VSUBS 0.074749f
C558 VTAIL.n22 VSUBS 0.047467f
C559 VTAIL.n23 VSUBS 0.194859f
C560 VTAIL.n24 VSUBS 0.033127f
C561 VTAIL.n25 VSUBS 0.02892f
C562 VTAIL.n26 VSUBS 0.01554f
C563 VTAIL.n27 VSUBS 0.036732f
C564 VTAIL.n28 VSUBS 0.016454f
C565 VTAIL.n29 VSUBS 0.49709f
C566 VTAIL.n30 VSUBS 0.01554f
C567 VTAIL.t6 VSUBS 0.080673f
C568 VTAIL.n31 VSUBS 0.118949f
C569 VTAIL.n32 VSUBS 0.02327f
C570 VTAIL.n33 VSUBS 0.027549f
C571 VTAIL.n34 VSUBS 0.036732f
C572 VTAIL.n35 VSUBS 0.016454f
C573 VTAIL.n36 VSUBS 0.01554f
C574 VTAIL.n37 VSUBS 0.02892f
C575 VTAIL.n38 VSUBS 0.02892f
C576 VTAIL.n39 VSUBS 0.01554f
C577 VTAIL.n40 VSUBS 0.016454f
C578 VTAIL.n41 VSUBS 0.036732f
C579 VTAIL.n42 VSUBS 0.093523f
C580 VTAIL.n43 VSUBS 0.016454f
C581 VTAIL.n44 VSUBS 0.01554f
C582 VTAIL.n45 VSUBS 0.074749f
C583 VTAIL.n46 VSUBS 0.047467f
C584 VTAIL.n47 VSUBS 0.30592f
C585 VTAIL.n48 VSUBS 0.033127f
C586 VTAIL.n49 VSUBS 0.02892f
C587 VTAIL.n50 VSUBS 0.01554f
C588 VTAIL.n51 VSUBS 0.036732f
C589 VTAIL.n52 VSUBS 0.016454f
C590 VTAIL.n53 VSUBS 0.49709f
C591 VTAIL.n54 VSUBS 0.01554f
C592 VTAIL.t7 VSUBS 0.080673f
C593 VTAIL.n55 VSUBS 0.118949f
C594 VTAIL.n56 VSUBS 0.02327f
C595 VTAIL.n57 VSUBS 0.027549f
C596 VTAIL.n58 VSUBS 0.036732f
C597 VTAIL.n59 VSUBS 0.016454f
C598 VTAIL.n60 VSUBS 0.01554f
C599 VTAIL.n61 VSUBS 0.02892f
C600 VTAIL.n62 VSUBS 0.02892f
C601 VTAIL.n63 VSUBS 0.01554f
C602 VTAIL.n64 VSUBS 0.016454f
C603 VTAIL.n65 VSUBS 0.036732f
C604 VTAIL.n66 VSUBS 0.093523f
C605 VTAIL.n67 VSUBS 0.016454f
C606 VTAIL.n68 VSUBS 0.01554f
C607 VTAIL.n69 VSUBS 0.074749f
C608 VTAIL.n70 VSUBS 0.047467f
C609 VTAIL.n71 VSUBS 1.27034f
C610 VTAIL.n72 VSUBS 0.033127f
C611 VTAIL.n73 VSUBS 0.02892f
C612 VTAIL.n74 VSUBS 0.01554f
C613 VTAIL.n75 VSUBS 0.036732f
C614 VTAIL.n76 VSUBS 0.016454f
C615 VTAIL.n77 VSUBS 0.49709f
C616 VTAIL.n78 VSUBS 0.01554f
C617 VTAIL.t1 VSUBS 0.080673f
C618 VTAIL.n79 VSUBS 0.118949f
C619 VTAIL.n80 VSUBS 0.02327f
C620 VTAIL.n81 VSUBS 0.027549f
C621 VTAIL.n82 VSUBS 0.036732f
C622 VTAIL.n83 VSUBS 0.016454f
C623 VTAIL.n84 VSUBS 0.01554f
C624 VTAIL.n85 VSUBS 0.02892f
C625 VTAIL.n86 VSUBS 0.02892f
C626 VTAIL.n87 VSUBS 0.01554f
C627 VTAIL.n88 VSUBS 0.016454f
C628 VTAIL.n89 VSUBS 0.036732f
C629 VTAIL.n90 VSUBS 0.093523f
C630 VTAIL.n91 VSUBS 0.016454f
C631 VTAIL.n92 VSUBS 0.01554f
C632 VTAIL.n93 VSUBS 0.074749f
C633 VTAIL.n94 VSUBS 0.047467f
C634 VTAIL.n95 VSUBS 1.27034f
C635 VTAIL.n96 VSUBS 0.033127f
C636 VTAIL.n97 VSUBS 0.02892f
C637 VTAIL.n98 VSUBS 0.01554f
C638 VTAIL.n99 VSUBS 0.036732f
C639 VTAIL.n100 VSUBS 0.016454f
C640 VTAIL.n101 VSUBS 0.49709f
C641 VTAIL.n102 VSUBS 0.01554f
C642 VTAIL.t3 VSUBS 0.080673f
C643 VTAIL.n103 VSUBS 0.118949f
C644 VTAIL.n104 VSUBS 0.02327f
C645 VTAIL.n105 VSUBS 0.027549f
C646 VTAIL.n106 VSUBS 0.036732f
C647 VTAIL.n107 VSUBS 0.016454f
C648 VTAIL.n108 VSUBS 0.01554f
C649 VTAIL.n109 VSUBS 0.02892f
C650 VTAIL.n110 VSUBS 0.02892f
C651 VTAIL.n111 VSUBS 0.01554f
C652 VTAIL.n112 VSUBS 0.016454f
C653 VTAIL.n113 VSUBS 0.036732f
C654 VTAIL.n114 VSUBS 0.093523f
C655 VTAIL.n115 VSUBS 0.016454f
C656 VTAIL.n116 VSUBS 0.01554f
C657 VTAIL.n117 VSUBS 0.074749f
C658 VTAIL.n118 VSUBS 0.047467f
C659 VTAIL.n119 VSUBS 0.30592f
C660 VTAIL.n120 VSUBS 0.033127f
C661 VTAIL.n121 VSUBS 0.02892f
C662 VTAIL.n122 VSUBS 0.01554f
C663 VTAIL.n123 VSUBS 0.036732f
C664 VTAIL.n124 VSUBS 0.016454f
C665 VTAIL.n125 VSUBS 0.49709f
C666 VTAIL.n126 VSUBS 0.01554f
C667 VTAIL.t5 VSUBS 0.080673f
C668 VTAIL.n127 VSUBS 0.118949f
C669 VTAIL.n128 VSUBS 0.02327f
C670 VTAIL.n129 VSUBS 0.027549f
C671 VTAIL.n130 VSUBS 0.036732f
C672 VTAIL.n131 VSUBS 0.016454f
C673 VTAIL.n132 VSUBS 0.01554f
C674 VTAIL.n133 VSUBS 0.02892f
C675 VTAIL.n134 VSUBS 0.02892f
C676 VTAIL.n135 VSUBS 0.01554f
C677 VTAIL.n136 VSUBS 0.016454f
C678 VTAIL.n137 VSUBS 0.036732f
C679 VTAIL.n138 VSUBS 0.093523f
C680 VTAIL.n139 VSUBS 0.016454f
C681 VTAIL.n140 VSUBS 0.01554f
C682 VTAIL.n141 VSUBS 0.074749f
C683 VTAIL.n142 VSUBS 0.047467f
C684 VTAIL.n143 VSUBS 0.30592f
C685 VTAIL.n144 VSUBS 0.033127f
C686 VTAIL.n145 VSUBS 0.02892f
C687 VTAIL.n146 VSUBS 0.01554f
C688 VTAIL.n147 VSUBS 0.036732f
C689 VTAIL.n148 VSUBS 0.016454f
C690 VTAIL.n149 VSUBS 0.49709f
C691 VTAIL.n150 VSUBS 0.01554f
C692 VTAIL.t4 VSUBS 0.080673f
C693 VTAIL.n151 VSUBS 0.118949f
C694 VTAIL.n152 VSUBS 0.02327f
C695 VTAIL.n153 VSUBS 0.027549f
C696 VTAIL.n154 VSUBS 0.036732f
C697 VTAIL.n155 VSUBS 0.016454f
C698 VTAIL.n156 VSUBS 0.01554f
C699 VTAIL.n157 VSUBS 0.02892f
C700 VTAIL.n158 VSUBS 0.02892f
C701 VTAIL.n159 VSUBS 0.01554f
C702 VTAIL.n160 VSUBS 0.016454f
C703 VTAIL.n161 VSUBS 0.036732f
C704 VTAIL.n162 VSUBS 0.093523f
C705 VTAIL.n163 VSUBS 0.016454f
C706 VTAIL.n164 VSUBS 0.01554f
C707 VTAIL.n165 VSUBS 0.074749f
C708 VTAIL.n166 VSUBS 0.047467f
C709 VTAIL.n167 VSUBS 1.27034f
C710 VTAIL.n168 VSUBS 0.033127f
C711 VTAIL.n169 VSUBS 0.02892f
C712 VTAIL.n170 VSUBS 0.01554f
C713 VTAIL.n171 VSUBS 0.036732f
C714 VTAIL.n172 VSUBS 0.016454f
C715 VTAIL.n173 VSUBS 0.49709f
C716 VTAIL.n174 VSUBS 0.01554f
C717 VTAIL.t0 VSUBS 0.080673f
C718 VTAIL.n175 VSUBS 0.118949f
C719 VTAIL.n176 VSUBS 0.02327f
C720 VTAIL.n177 VSUBS 0.027549f
C721 VTAIL.n178 VSUBS 0.036732f
C722 VTAIL.n179 VSUBS 0.016454f
C723 VTAIL.n180 VSUBS 0.01554f
C724 VTAIL.n181 VSUBS 0.02892f
C725 VTAIL.n182 VSUBS 0.02892f
C726 VTAIL.n183 VSUBS 0.01554f
C727 VTAIL.n184 VSUBS 0.016454f
C728 VTAIL.n185 VSUBS 0.036732f
C729 VTAIL.n186 VSUBS 0.093523f
C730 VTAIL.n187 VSUBS 0.016454f
C731 VTAIL.n188 VSUBS 0.01554f
C732 VTAIL.n189 VSUBS 0.074749f
C733 VTAIL.n190 VSUBS 0.047467f
C734 VTAIL.n191 VSUBS 1.14843f
C735 VDD1.t0 VSUBS 0.106563f
C736 VDD1.t2 VSUBS 0.106563f
C737 VDD1.n0 VSUBS 0.661572f
C738 VDD1.t3 VSUBS 0.106563f
C739 VDD1.t1 VSUBS 0.106563f
C740 VDD1.n1 VSUBS 1.03781f
C741 VP.n0 VSUBS 0.060839f
C742 VP.t1 VSUBS 1.47133f
C743 VP.n1 VSUBS 0.067084f
C744 VP.n2 VSUBS 0.046149f
C745 VP.t0 VSUBS 1.47133f
C746 VP.n3 VSUBS 0.721122f
C747 VP.t3 VSUBS 1.84958f
C748 VP.t2 VSUBS 1.85761f
C749 VP.n4 VSUBS 3.20839f
C750 VP.n5 VSUBS 2.13401f
C751 VP.n6 VSUBS 0.060839f
C752 VP.n7 VSUBS 0.06023f
C753 VP.n8 VSUBS 0.085579f
C754 VP.n9 VSUBS 0.067084f
C755 VP.n10 VSUBS 0.046149f
C756 VP.n11 VSUBS 0.046149f
C757 VP.n12 VSUBS 0.046149f
C758 VP.n13 VSUBS 0.085579f
C759 VP.n14 VSUBS 0.06023f
C760 VP.n15 VSUBS 0.721122f
C761 VP.n16 VSUBS 0.074851f
.ends

