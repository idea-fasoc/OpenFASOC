* NGSPICE file created from diff_pair_sample_1456.ext - technology: sky130A

.subckt diff_pair_sample_1456 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t17 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=6.2088 ps=32.62 w=15.92 l=0.31
X1 VTAIL.t1 VN.t0 VDD2.t9 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X2 B.t11 B.t9 B.t10 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=0 ps=0 w=15.92 l=0.31
X3 VDD2.t8 VN.t1 VTAIL.t6 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=2.6268 ps=16.25 w=15.92 l=0.31
X4 B.t8 B.t6 B.t7 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=0 ps=0 w=15.92 l=0.31
X5 VDD2.t7 VN.t2 VTAIL.t4 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=2.6268 ps=16.25 w=15.92 l=0.31
X6 VTAIL.t16 VP.t1 VDD1.t8 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X7 VDD1.t7 VP.t2 VTAIL.t19 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=2.6268 ps=16.25 w=15.92 l=0.31
X8 VTAIL.t18 VP.t3 VDD1.t6 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X9 VDD1.t5 VP.t4 VTAIL.t14 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X10 VDD1.t4 VP.t5 VTAIL.t15 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=2.6268 ps=16.25 w=15.92 l=0.31
X11 VDD2.t6 VN.t3 VTAIL.t8 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=6.2088 ps=32.62 w=15.92 l=0.31
X12 VTAIL.t9 VN.t4 VDD2.t5 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X13 VTAIL.t13 VP.t6 VDD1.t3 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X14 B.t5 B.t3 B.t4 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=0 ps=0 w=15.92 l=0.31
X15 B.t2 B.t0 B.t1 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=6.2088 pd=32.62 as=0 ps=0 w=15.92 l=0.31
X16 VDD1.t2 VP.t7 VTAIL.t11 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=6.2088 ps=32.62 w=15.92 l=0.31
X17 VDD1.t1 VP.t8 VTAIL.t10 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X18 VDD2.t4 VN.t5 VTAIL.t3 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X19 VTAIL.t0 VN.t6 VDD2.t3 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X20 VDD2.t2 VN.t7 VTAIL.t5 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=6.2088 ps=32.62 w=15.92 l=0.31
X21 VTAIL.t2 VN.t8 VDD2.t1 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X22 VDD2.t0 VN.t9 VTAIL.t7 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
X23 VTAIL.t12 VP.t9 VDD1.t0 w_n1738_n4152# sky130_fd_pr__pfet_01v8 ad=2.6268 pd=16.25 as=2.6268 ps=16.25 w=15.92 l=0.31
R0 VP.n21 VP.t7 1381.17
R1 VP.n14 VP.t2 1381.17
R2 VP.n5 VP.t5 1381.17
R3 VP.n11 VP.t0 1381.17
R4 VP.n18 VP.t4 1340.27
R5 VP.n20 VP.t3 1340.27
R6 VP.n13 VP.t6 1340.27
R7 VP.n8 VP.t8 1340.27
R8 VP.n4 VP.t9 1340.27
R9 VP.n10 VP.t1 1340.27
R10 VP.n6 VP.n5 161.489
R11 VP.n22 VP.n21 161.3
R12 VP.n6 VP.n3 161.3
R13 VP.n8 VP.n7 161.3
R14 VP.n9 VP.n2 161.3
R15 VP.n12 VP.n11 161.3
R16 VP.n19 VP.n0 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n1 161.3
R19 VP.n15 VP.n14 161.3
R20 VP.n18 VP.n1 73.0308
R21 VP.n19 VP.n18 73.0308
R22 VP.n8 VP.n3 73.0308
R23 VP.n9 VP.n8 73.0308
R24 VP.n14 VP.n13 52.5823
R25 VP.n21 VP.n20 52.5823
R26 VP.n5 VP.n4 52.5823
R27 VP.n11 VP.n10 52.5823
R28 VP.n15 VP.n12 43.705
R29 VP.n13 VP.n1 20.449
R30 VP.n20 VP.n19 20.449
R31 VP.n4 VP.n3 20.449
R32 VP.n10 VP.n9 20.449
R33 VP.n7 VP.n6 0.189894
R34 VP.n7 VP.n2 0.189894
R35 VP.n12 VP.n2 0.189894
R36 VP.n16 VP.n15 0.189894
R37 VP.n17 VP.n16 0.189894
R38 VP.n17 VP.n0 0.189894
R39 VP.n22 VP.n0 0.189894
R40 VP VP.n22 0.0516364
R41 VTAIL.n11 VTAIL.t8 59.2655
R42 VTAIL.n16 VTAIL.t17 59.2654
R43 VTAIL.n17 VTAIL.t5 59.2654
R44 VTAIL.n2 VTAIL.t11 59.2654
R45 VTAIL.n15 VTAIL.n14 57.2238
R46 VTAIL.n13 VTAIL.n12 57.2238
R47 VTAIL.n10 VTAIL.n9 57.2238
R48 VTAIL.n8 VTAIL.n7 57.2238
R49 VTAIL.n19 VTAIL.n18 57.2235
R50 VTAIL.n1 VTAIL.n0 57.2235
R51 VTAIL.n4 VTAIL.n3 57.2235
R52 VTAIL.n6 VTAIL.n5 57.2235
R53 VTAIL.n8 VTAIL.n6 27.1945
R54 VTAIL.n17 VTAIL.n16 26.6427
R55 VTAIL.n18 VTAIL.t7 2.04227
R56 VTAIL.n18 VTAIL.t0 2.04227
R57 VTAIL.n0 VTAIL.t4 2.04227
R58 VTAIL.n0 VTAIL.t2 2.04227
R59 VTAIL.n3 VTAIL.t14 2.04227
R60 VTAIL.n3 VTAIL.t18 2.04227
R61 VTAIL.n5 VTAIL.t19 2.04227
R62 VTAIL.n5 VTAIL.t13 2.04227
R63 VTAIL.n14 VTAIL.t10 2.04227
R64 VTAIL.n14 VTAIL.t16 2.04227
R65 VTAIL.n12 VTAIL.t15 2.04227
R66 VTAIL.n12 VTAIL.t12 2.04227
R67 VTAIL.n9 VTAIL.t3 2.04227
R68 VTAIL.n9 VTAIL.t1 2.04227
R69 VTAIL.n7 VTAIL.t6 2.04227
R70 VTAIL.n7 VTAIL.t9 2.04227
R71 VTAIL.n13 VTAIL.n11 0.74619
R72 VTAIL.n2 VTAIL.n1 0.74619
R73 VTAIL.n10 VTAIL.n8 0.552224
R74 VTAIL.n11 VTAIL.n10 0.552224
R75 VTAIL.n15 VTAIL.n13 0.552224
R76 VTAIL.n16 VTAIL.n15 0.552224
R77 VTAIL.n6 VTAIL.n4 0.552224
R78 VTAIL.n4 VTAIL.n2 0.552224
R79 VTAIL.n19 VTAIL.n17 0.552224
R80 VTAIL VTAIL.n1 0.472483
R81 VTAIL VTAIL.n19 0.0802414
R82 VDD1.n1 VDD1.t4 76.496
R83 VDD1.n3 VDD1.t7 76.4959
R84 VDD1.n5 VDD1.n4 74.2607
R85 VDD1.n1 VDD1.n0 73.9026
R86 VDD1.n7 VDD1.n6 73.9024
R87 VDD1.n3 VDD1.n2 73.9023
R88 VDD1.n7 VDD1.n5 40.919
R89 VDD1.n6 VDD1.t8 2.04227
R90 VDD1.n6 VDD1.t9 2.04227
R91 VDD1.n0 VDD1.t0 2.04227
R92 VDD1.n0 VDD1.t1 2.04227
R93 VDD1.n4 VDD1.t6 2.04227
R94 VDD1.n4 VDD1.t2 2.04227
R95 VDD1.n2 VDD1.t3 2.04227
R96 VDD1.n2 VDD1.t5 2.04227
R97 VDD1 VDD1.n7 0.356103
R98 VDD1 VDD1.n1 0.196621
R99 VDD1.n5 VDD1.n3 0.083085
R100 VN.n9 VN.t7 1381.17
R101 VN.n3 VN.t2 1381.17
R102 VN.n20 VN.t1 1381.17
R103 VN.n14 VN.t3 1381.17
R104 VN.n6 VN.t9 1340.27
R105 VN.n8 VN.t6 1340.27
R106 VN.n2 VN.t8 1340.27
R107 VN.n17 VN.t5 1340.27
R108 VN.n19 VN.t4 1340.27
R109 VN.n13 VN.t0 1340.27
R110 VN.n15 VN.n14 161.489
R111 VN.n4 VN.n3 161.489
R112 VN.n10 VN.n9 161.3
R113 VN.n21 VN.n20 161.3
R114 VN.n18 VN.n11 161.3
R115 VN.n17 VN.n16 161.3
R116 VN.n15 VN.n12 161.3
R117 VN.n7 VN.n0 161.3
R118 VN.n6 VN.n5 161.3
R119 VN.n4 VN.n1 161.3
R120 VN.n6 VN.n1 73.0308
R121 VN.n7 VN.n6 73.0308
R122 VN.n18 VN.n17 73.0308
R123 VN.n17 VN.n12 73.0308
R124 VN.n3 VN.n2 52.5823
R125 VN.n9 VN.n8 52.5823
R126 VN.n20 VN.n19 52.5823
R127 VN.n14 VN.n13 52.5823
R128 VN VN.n21 44.0857
R129 VN.n2 VN.n1 20.449
R130 VN.n8 VN.n7 20.449
R131 VN.n19 VN.n18 20.449
R132 VN.n13 VN.n12 20.449
R133 VN.n21 VN.n11 0.189894
R134 VN.n16 VN.n11 0.189894
R135 VN.n16 VN.n15 0.189894
R136 VN.n5 VN.n4 0.189894
R137 VN.n5 VN.n0 0.189894
R138 VN.n10 VN.n0 0.189894
R139 VN VN.n10 0.0516364
R140 VDD2.n1 VDD2.t7 76.4959
R141 VDD2.n4 VDD2.t8 75.9443
R142 VDD2.n3 VDD2.n2 74.2607
R143 VDD2 VDD2.n7 74.258
R144 VDD2.n6 VDD2.n5 73.9026
R145 VDD2.n1 VDD2.n0 73.9023
R146 VDD2.n4 VDD2.n3 40.0601
R147 VDD2.n7 VDD2.t9 2.04227
R148 VDD2.n7 VDD2.t6 2.04227
R149 VDD2.n5 VDD2.t5 2.04227
R150 VDD2.n5 VDD2.t4 2.04227
R151 VDD2.n2 VDD2.t3 2.04227
R152 VDD2.n2 VDD2.t2 2.04227
R153 VDD2.n0 VDD2.t1 2.04227
R154 VDD2.n0 VDD2.t0 2.04227
R155 VDD2.n6 VDD2.n4 0.552224
R156 VDD2 VDD2.n6 0.196621
R157 VDD2.n3 VDD2.n1 0.083085
R158 B.n126 B.t9 1452.62
R159 B.n284 B.t0 1452.62
R160 B.n46 B.t6 1452.62
R161 B.n38 B.t3 1452.62
R162 B.n367 B.n94 585
R163 B.n366 B.n365 585
R164 B.n364 B.n95 585
R165 B.n363 B.n362 585
R166 B.n361 B.n96 585
R167 B.n360 B.n359 585
R168 B.n358 B.n97 585
R169 B.n357 B.n356 585
R170 B.n355 B.n98 585
R171 B.n354 B.n353 585
R172 B.n352 B.n99 585
R173 B.n351 B.n350 585
R174 B.n349 B.n100 585
R175 B.n348 B.n347 585
R176 B.n346 B.n101 585
R177 B.n345 B.n344 585
R178 B.n343 B.n102 585
R179 B.n342 B.n341 585
R180 B.n340 B.n103 585
R181 B.n339 B.n338 585
R182 B.n337 B.n104 585
R183 B.n336 B.n335 585
R184 B.n334 B.n105 585
R185 B.n333 B.n332 585
R186 B.n331 B.n106 585
R187 B.n330 B.n329 585
R188 B.n328 B.n107 585
R189 B.n327 B.n326 585
R190 B.n325 B.n108 585
R191 B.n324 B.n323 585
R192 B.n322 B.n109 585
R193 B.n321 B.n320 585
R194 B.n319 B.n110 585
R195 B.n318 B.n317 585
R196 B.n316 B.n111 585
R197 B.n315 B.n314 585
R198 B.n313 B.n112 585
R199 B.n312 B.n311 585
R200 B.n310 B.n113 585
R201 B.n309 B.n308 585
R202 B.n307 B.n114 585
R203 B.n306 B.n305 585
R204 B.n304 B.n115 585
R205 B.n303 B.n302 585
R206 B.n301 B.n116 585
R207 B.n300 B.n299 585
R208 B.n298 B.n117 585
R209 B.n297 B.n296 585
R210 B.n295 B.n118 585
R211 B.n294 B.n293 585
R212 B.n292 B.n119 585
R213 B.n291 B.n290 585
R214 B.n289 B.n120 585
R215 B.n288 B.n287 585
R216 B.n283 B.n121 585
R217 B.n282 B.n281 585
R218 B.n280 B.n122 585
R219 B.n279 B.n278 585
R220 B.n277 B.n123 585
R221 B.n276 B.n275 585
R222 B.n274 B.n124 585
R223 B.n273 B.n272 585
R224 B.n271 B.n125 585
R225 B.n269 B.n268 585
R226 B.n267 B.n128 585
R227 B.n266 B.n265 585
R228 B.n264 B.n129 585
R229 B.n263 B.n262 585
R230 B.n261 B.n130 585
R231 B.n260 B.n259 585
R232 B.n258 B.n131 585
R233 B.n257 B.n256 585
R234 B.n255 B.n132 585
R235 B.n254 B.n253 585
R236 B.n252 B.n133 585
R237 B.n251 B.n250 585
R238 B.n249 B.n134 585
R239 B.n248 B.n247 585
R240 B.n246 B.n135 585
R241 B.n245 B.n244 585
R242 B.n243 B.n136 585
R243 B.n242 B.n241 585
R244 B.n240 B.n137 585
R245 B.n239 B.n238 585
R246 B.n237 B.n138 585
R247 B.n236 B.n235 585
R248 B.n234 B.n139 585
R249 B.n233 B.n232 585
R250 B.n231 B.n140 585
R251 B.n230 B.n229 585
R252 B.n228 B.n141 585
R253 B.n227 B.n226 585
R254 B.n225 B.n142 585
R255 B.n224 B.n223 585
R256 B.n222 B.n143 585
R257 B.n221 B.n220 585
R258 B.n219 B.n144 585
R259 B.n218 B.n217 585
R260 B.n216 B.n145 585
R261 B.n215 B.n214 585
R262 B.n213 B.n146 585
R263 B.n212 B.n211 585
R264 B.n210 B.n147 585
R265 B.n209 B.n208 585
R266 B.n207 B.n148 585
R267 B.n206 B.n205 585
R268 B.n204 B.n149 585
R269 B.n203 B.n202 585
R270 B.n201 B.n150 585
R271 B.n200 B.n199 585
R272 B.n198 B.n151 585
R273 B.n197 B.n196 585
R274 B.n195 B.n152 585
R275 B.n194 B.n193 585
R276 B.n192 B.n153 585
R277 B.n191 B.n190 585
R278 B.n369 B.n368 585
R279 B.n370 B.n93 585
R280 B.n372 B.n371 585
R281 B.n373 B.n92 585
R282 B.n375 B.n374 585
R283 B.n376 B.n91 585
R284 B.n378 B.n377 585
R285 B.n379 B.n90 585
R286 B.n381 B.n380 585
R287 B.n382 B.n89 585
R288 B.n384 B.n383 585
R289 B.n385 B.n88 585
R290 B.n387 B.n386 585
R291 B.n388 B.n87 585
R292 B.n390 B.n389 585
R293 B.n391 B.n86 585
R294 B.n393 B.n392 585
R295 B.n394 B.n85 585
R296 B.n396 B.n395 585
R297 B.n397 B.n84 585
R298 B.n399 B.n398 585
R299 B.n400 B.n83 585
R300 B.n402 B.n401 585
R301 B.n403 B.n82 585
R302 B.n405 B.n404 585
R303 B.n406 B.n81 585
R304 B.n408 B.n407 585
R305 B.n409 B.n80 585
R306 B.n411 B.n410 585
R307 B.n412 B.n79 585
R308 B.n414 B.n413 585
R309 B.n415 B.n78 585
R310 B.n417 B.n416 585
R311 B.n418 B.n77 585
R312 B.n420 B.n419 585
R313 B.n421 B.n76 585
R314 B.n423 B.n422 585
R315 B.n424 B.n75 585
R316 B.n426 B.n425 585
R317 B.n427 B.n74 585
R318 B.n603 B.n602 585
R319 B.n601 B.n12 585
R320 B.n600 B.n599 585
R321 B.n598 B.n13 585
R322 B.n597 B.n596 585
R323 B.n595 B.n14 585
R324 B.n594 B.n593 585
R325 B.n592 B.n15 585
R326 B.n591 B.n590 585
R327 B.n589 B.n16 585
R328 B.n588 B.n587 585
R329 B.n586 B.n17 585
R330 B.n585 B.n584 585
R331 B.n583 B.n18 585
R332 B.n582 B.n581 585
R333 B.n580 B.n19 585
R334 B.n579 B.n578 585
R335 B.n577 B.n20 585
R336 B.n576 B.n575 585
R337 B.n574 B.n21 585
R338 B.n573 B.n572 585
R339 B.n571 B.n22 585
R340 B.n570 B.n569 585
R341 B.n568 B.n23 585
R342 B.n567 B.n566 585
R343 B.n565 B.n24 585
R344 B.n564 B.n563 585
R345 B.n562 B.n25 585
R346 B.n561 B.n560 585
R347 B.n559 B.n26 585
R348 B.n558 B.n557 585
R349 B.n556 B.n27 585
R350 B.n555 B.n554 585
R351 B.n553 B.n28 585
R352 B.n552 B.n551 585
R353 B.n550 B.n29 585
R354 B.n549 B.n548 585
R355 B.n547 B.n30 585
R356 B.n546 B.n545 585
R357 B.n544 B.n31 585
R358 B.n543 B.n542 585
R359 B.n541 B.n32 585
R360 B.n540 B.n539 585
R361 B.n538 B.n33 585
R362 B.n537 B.n536 585
R363 B.n535 B.n34 585
R364 B.n534 B.n533 585
R365 B.n532 B.n35 585
R366 B.n531 B.n530 585
R367 B.n529 B.n36 585
R368 B.n528 B.n527 585
R369 B.n526 B.n37 585
R370 B.n525 B.n524 585
R371 B.n523 B.n522 585
R372 B.n521 B.n41 585
R373 B.n520 B.n519 585
R374 B.n518 B.n42 585
R375 B.n517 B.n516 585
R376 B.n515 B.n43 585
R377 B.n514 B.n513 585
R378 B.n512 B.n44 585
R379 B.n511 B.n510 585
R380 B.n509 B.n45 585
R381 B.n507 B.n506 585
R382 B.n505 B.n48 585
R383 B.n504 B.n503 585
R384 B.n502 B.n49 585
R385 B.n501 B.n500 585
R386 B.n499 B.n50 585
R387 B.n498 B.n497 585
R388 B.n496 B.n51 585
R389 B.n495 B.n494 585
R390 B.n493 B.n52 585
R391 B.n492 B.n491 585
R392 B.n490 B.n53 585
R393 B.n489 B.n488 585
R394 B.n487 B.n54 585
R395 B.n486 B.n485 585
R396 B.n484 B.n55 585
R397 B.n483 B.n482 585
R398 B.n481 B.n56 585
R399 B.n480 B.n479 585
R400 B.n478 B.n57 585
R401 B.n477 B.n476 585
R402 B.n475 B.n58 585
R403 B.n474 B.n473 585
R404 B.n472 B.n59 585
R405 B.n471 B.n470 585
R406 B.n469 B.n60 585
R407 B.n468 B.n467 585
R408 B.n466 B.n61 585
R409 B.n465 B.n464 585
R410 B.n463 B.n62 585
R411 B.n462 B.n461 585
R412 B.n460 B.n63 585
R413 B.n459 B.n458 585
R414 B.n457 B.n64 585
R415 B.n456 B.n455 585
R416 B.n454 B.n65 585
R417 B.n453 B.n452 585
R418 B.n451 B.n66 585
R419 B.n450 B.n449 585
R420 B.n448 B.n67 585
R421 B.n447 B.n446 585
R422 B.n445 B.n68 585
R423 B.n444 B.n443 585
R424 B.n442 B.n69 585
R425 B.n441 B.n440 585
R426 B.n439 B.n70 585
R427 B.n438 B.n437 585
R428 B.n436 B.n71 585
R429 B.n435 B.n434 585
R430 B.n433 B.n72 585
R431 B.n432 B.n431 585
R432 B.n430 B.n73 585
R433 B.n429 B.n428 585
R434 B.n604 B.n11 585
R435 B.n606 B.n605 585
R436 B.n607 B.n10 585
R437 B.n609 B.n608 585
R438 B.n610 B.n9 585
R439 B.n612 B.n611 585
R440 B.n613 B.n8 585
R441 B.n615 B.n614 585
R442 B.n616 B.n7 585
R443 B.n618 B.n617 585
R444 B.n619 B.n6 585
R445 B.n621 B.n620 585
R446 B.n622 B.n5 585
R447 B.n624 B.n623 585
R448 B.n625 B.n4 585
R449 B.n627 B.n626 585
R450 B.n628 B.n3 585
R451 B.n630 B.n629 585
R452 B.n631 B.n0 585
R453 B.n2 B.n1 585
R454 B.n164 B.n163 585
R455 B.n165 B.n162 585
R456 B.n167 B.n166 585
R457 B.n168 B.n161 585
R458 B.n170 B.n169 585
R459 B.n171 B.n160 585
R460 B.n173 B.n172 585
R461 B.n174 B.n159 585
R462 B.n176 B.n175 585
R463 B.n177 B.n158 585
R464 B.n179 B.n178 585
R465 B.n180 B.n157 585
R466 B.n182 B.n181 585
R467 B.n183 B.n156 585
R468 B.n185 B.n184 585
R469 B.n186 B.n155 585
R470 B.n188 B.n187 585
R471 B.n189 B.n154 585
R472 B.n190 B.n189 473.281
R473 B.n368 B.n367 473.281
R474 B.n428 B.n427 473.281
R475 B.n602 B.n11 473.281
R476 B.n633 B.n632 256.663
R477 B.n632 B.n631 235.042
R478 B.n632 B.n2 235.042
R479 B.n190 B.n153 163.367
R480 B.n194 B.n153 163.367
R481 B.n195 B.n194 163.367
R482 B.n196 B.n195 163.367
R483 B.n196 B.n151 163.367
R484 B.n200 B.n151 163.367
R485 B.n201 B.n200 163.367
R486 B.n202 B.n201 163.367
R487 B.n202 B.n149 163.367
R488 B.n206 B.n149 163.367
R489 B.n207 B.n206 163.367
R490 B.n208 B.n207 163.367
R491 B.n208 B.n147 163.367
R492 B.n212 B.n147 163.367
R493 B.n213 B.n212 163.367
R494 B.n214 B.n213 163.367
R495 B.n214 B.n145 163.367
R496 B.n218 B.n145 163.367
R497 B.n219 B.n218 163.367
R498 B.n220 B.n219 163.367
R499 B.n220 B.n143 163.367
R500 B.n224 B.n143 163.367
R501 B.n225 B.n224 163.367
R502 B.n226 B.n225 163.367
R503 B.n226 B.n141 163.367
R504 B.n230 B.n141 163.367
R505 B.n231 B.n230 163.367
R506 B.n232 B.n231 163.367
R507 B.n232 B.n139 163.367
R508 B.n236 B.n139 163.367
R509 B.n237 B.n236 163.367
R510 B.n238 B.n237 163.367
R511 B.n238 B.n137 163.367
R512 B.n242 B.n137 163.367
R513 B.n243 B.n242 163.367
R514 B.n244 B.n243 163.367
R515 B.n244 B.n135 163.367
R516 B.n248 B.n135 163.367
R517 B.n249 B.n248 163.367
R518 B.n250 B.n249 163.367
R519 B.n250 B.n133 163.367
R520 B.n254 B.n133 163.367
R521 B.n255 B.n254 163.367
R522 B.n256 B.n255 163.367
R523 B.n256 B.n131 163.367
R524 B.n260 B.n131 163.367
R525 B.n261 B.n260 163.367
R526 B.n262 B.n261 163.367
R527 B.n262 B.n129 163.367
R528 B.n266 B.n129 163.367
R529 B.n267 B.n266 163.367
R530 B.n268 B.n267 163.367
R531 B.n268 B.n125 163.367
R532 B.n273 B.n125 163.367
R533 B.n274 B.n273 163.367
R534 B.n275 B.n274 163.367
R535 B.n275 B.n123 163.367
R536 B.n279 B.n123 163.367
R537 B.n280 B.n279 163.367
R538 B.n281 B.n280 163.367
R539 B.n281 B.n121 163.367
R540 B.n288 B.n121 163.367
R541 B.n289 B.n288 163.367
R542 B.n290 B.n289 163.367
R543 B.n290 B.n119 163.367
R544 B.n294 B.n119 163.367
R545 B.n295 B.n294 163.367
R546 B.n296 B.n295 163.367
R547 B.n296 B.n117 163.367
R548 B.n300 B.n117 163.367
R549 B.n301 B.n300 163.367
R550 B.n302 B.n301 163.367
R551 B.n302 B.n115 163.367
R552 B.n306 B.n115 163.367
R553 B.n307 B.n306 163.367
R554 B.n308 B.n307 163.367
R555 B.n308 B.n113 163.367
R556 B.n312 B.n113 163.367
R557 B.n313 B.n312 163.367
R558 B.n314 B.n313 163.367
R559 B.n314 B.n111 163.367
R560 B.n318 B.n111 163.367
R561 B.n319 B.n318 163.367
R562 B.n320 B.n319 163.367
R563 B.n320 B.n109 163.367
R564 B.n324 B.n109 163.367
R565 B.n325 B.n324 163.367
R566 B.n326 B.n325 163.367
R567 B.n326 B.n107 163.367
R568 B.n330 B.n107 163.367
R569 B.n331 B.n330 163.367
R570 B.n332 B.n331 163.367
R571 B.n332 B.n105 163.367
R572 B.n336 B.n105 163.367
R573 B.n337 B.n336 163.367
R574 B.n338 B.n337 163.367
R575 B.n338 B.n103 163.367
R576 B.n342 B.n103 163.367
R577 B.n343 B.n342 163.367
R578 B.n344 B.n343 163.367
R579 B.n344 B.n101 163.367
R580 B.n348 B.n101 163.367
R581 B.n349 B.n348 163.367
R582 B.n350 B.n349 163.367
R583 B.n350 B.n99 163.367
R584 B.n354 B.n99 163.367
R585 B.n355 B.n354 163.367
R586 B.n356 B.n355 163.367
R587 B.n356 B.n97 163.367
R588 B.n360 B.n97 163.367
R589 B.n361 B.n360 163.367
R590 B.n362 B.n361 163.367
R591 B.n362 B.n95 163.367
R592 B.n366 B.n95 163.367
R593 B.n367 B.n366 163.367
R594 B.n427 B.n426 163.367
R595 B.n426 B.n75 163.367
R596 B.n422 B.n75 163.367
R597 B.n422 B.n421 163.367
R598 B.n421 B.n420 163.367
R599 B.n420 B.n77 163.367
R600 B.n416 B.n77 163.367
R601 B.n416 B.n415 163.367
R602 B.n415 B.n414 163.367
R603 B.n414 B.n79 163.367
R604 B.n410 B.n79 163.367
R605 B.n410 B.n409 163.367
R606 B.n409 B.n408 163.367
R607 B.n408 B.n81 163.367
R608 B.n404 B.n81 163.367
R609 B.n404 B.n403 163.367
R610 B.n403 B.n402 163.367
R611 B.n402 B.n83 163.367
R612 B.n398 B.n83 163.367
R613 B.n398 B.n397 163.367
R614 B.n397 B.n396 163.367
R615 B.n396 B.n85 163.367
R616 B.n392 B.n85 163.367
R617 B.n392 B.n391 163.367
R618 B.n391 B.n390 163.367
R619 B.n390 B.n87 163.367
R620 B.n386 B.n87 163.367
R621 B.n386 B.n385 163.367
R622 B.n385 B.n384 163.367
R623 B.n384 B.n89 163.367
R624 B.n380 B.n89 163.367
R625 B.n380 B.n379 163.367
R626 B.n379 B.n378 163.367
R627 B.n378 B.n91 163.367
R628 B.n374 B.n91 163.367
R629 B.n374 B.n373 163.367
R630 B.n373 B.n372 163.367
R631 B.n372 B.n93 163.367
R632 B.n368 B.n93 163.367
R633 B.n602 B.n601 163.367
R634 B.n601 B.n600 163.367
R635 B.n600 B.n13 163.367
R636 B.n596 B.n13 163.367
R637 B.n596 B.n595 163.367
R638 B.n595 B.n594 163.367
R639 B.n594 B.n15 163.367
R640 B.n590 B.n15 163.367
R641 B.n590 B.n589 163.367
R642 B.n589 B.n588 163.367
R643 B.n588 B.n17 163.367
R644 B.n584 B.n17 163.367
R645 B.n584 B.n583 163.367
R646 B.n583 B.n582 163.367
R647 B.n582 B.n19 163.367
R648 B.n578 B.n19 163.367
R649 B.n578 B.n577 163.367
R650 B.n577 B.n576 163.367
R651 B.n576 B.n21 163.367
R652 B.n572 B.n21 163.367
R653 B.n572 B.n571 163.367
R654 B.n571 B.n570 163.367
R655 B.n570 B.n23 163.367
R656 B.n566 B.n23 163.367
R657 B.n566 B.n565 163.367
R658 B.n565 B.n564 163.367
R659 B.n564 B.n25 163.367
R660 B.n560 B.n25 163.367
R661 B.n560 B.n559 163.367
R662 B.n559 B.n558 163.367
R663 B.n558 B.n27 163.367
R664 B.n554 B.n27 163.367
R665 B.n554 B.n553 163.367
R666 B.n553 B.n552 163.367
R667 B.n552 B.n29 163.367
R668 B.n548 B.n29 163.367
R669 B.n548 B.n547 163.367
R670 B.n547 B.n546 163.367
R671 B.n546 B.n31 163.367
R672 B.n542 B.n31 163.367
R673 B.n542 B.n541 163.367
R674 B.n541 B.n540 163.367
R675 B.n540 B.n33 163.367
R676 B.n536 B.n33 163.367
R677 B.n536 B.n535 163.367
R678 B.n535 B.n534 163.367
R679 B.n534 B.n35 163.367
R680 B.n530 B.n35 163.367
R681 B.n530 B.n529 163.367
R682 B.n529 B.n528 163.367
R683 B.n528 B.n37 163.367
R684 B.n524 B.n37 163.367
R685 B.n524 B.n523 163.367
R686 B.n523 B.n41 163.367
R687 B.n519 B.n41 163.367
R688 B.n519 B.n518 163.367
R689 B.n518 B.n517 163.367
R690 B.n517 B.n43 163.367
R691 B.n513 B.n43 163.367
R692 B.n513 B.n512 163.367
R693 B.n512 B.n511 163.367
R694 B.n511 B.n45 163.367
R695 B.n506 B.n45 163.367
R696 B.n506 B.n505 163.367
R697 B.n505 B.n504 163.367
R698 B.n504 B.n49 163.367
R699 B.n500 B.n49 163.367
R700 B.n500 B.n499 163.367
R701 B.n499 B.n498 163.367
R702 B.n498 B.n51 163.367
R703 B.n494 B.n51 163.367
R704 B.n494 B.n493 163.367
R705 B.n493 B.n492 163.367
R706 B.n492 B.n53 163.367
R707 B.n488 B.n53 163.367
R708 B.n488 B.n487 163.367
R709 B.n487 B.n486 163.367
R710 B.n486 B.n55 163.367
R711 B.n482 B.n55 163.367
R712 B.n482 B.n481 163.367
R713 B.n481 B.n480 163.367
R714 B.n480 B.n57 163.367
R715 B.n476 B.n57 163.367
R716 B.n476 B.n475 163.367
R717 B.n475 B.n474 163.367
R718 B.n474 B.n59 163.367
R719 B.n470 B.n59 163.367
R720 B.n470 B.n469 163.367
R721 B.n469 B.n468 163.367
R722 B.n468 B.n61 163.367
R723 B.n464 B.n61 163.367
R724 B.n464 B.n463 163.367
R725 B.n463 B.n462 163.367
R726 B.n462 B.n63 163.367
R727 B.n458 B.n63 163.367
R728 B.n458 B.n457 163.367
R729 B.n457 B.n456 163.367
R730 B.n456 B.n65 163.367
R731 B.n452 B.n65 163.367
R732 B.n452 B.n451 163.367
R733 B.n451 B.n450 163.367
R734 B.n450 B.n67 163.367
R735 B.n446 B.n67 163.367
R736 B.n446 B.n445 163.367
R737 B.n445 B.n444 163.367
R738 B.n444 B.n69 163.367
R739 B.n440 B.n69 163.367
R740 B.n440 B.n439 163.367
R741 B.n439 B.n438 163.367
R742 B.n438 B.n71 163.367
R743 B.n434 B.n71 163.367
R744 B.n434 B.n433 163.367
R745 B.n433 B.n432 163.367
R746 B.n432 B.n73 163.367
R747 B.n428 B.n73 163.367
R748 B.n606 B.n11 163.367
R749 B.n607 B.n606 163.367
R750 B.n608 B.n607 163.367
R751 B.n608 B.n9 163.367
R752 B.n612 B.n9 163.367
R753 B.n613 B.n612 163.367
R754 B.n614 B.n613 163.367
R755 B.n614 B.n7 163.367
R756 B.n618 B.n7 163.367
R757 B.n619 B.n618 163.367
R758 B.n620 B.n619 163.367
R759 B.n620 B.n5 163.367
R760 B.n624 B.n5 163.367
R761 B.n625 B.n624 163.367
R762 B.n626 B.n625 163.367
R763 B.n626 B.n3 163.367
R764 B.n630 B.n3 163.367
R765 B.n631 B.n630 163.367
R766 B.n164 B.n2 163.367
R767 B.n165 B.n164 163.367
R768 B.n166 B.n165 163.367
R769 B.n166 B.n161 163.367
R770 B.n170 B.n161 163.367
R771 B.n171 B.n170 163.367
R772 B.n172 B.n171 163.367
R773 B.n172 B.n159 163.367
R774 B.n176 B.n159 163.367
R775 B.n177 B.n176 163.367
R776 B.n178 B.n177 163.367
R777 B.n178 B.n157 163.367
R778 B.n182 B.n157 163.367
R779 B.n183 B.n182 163.367
R780 B.n184 B.n183 163.367
R781 B.n184 B.n155 163.367
R782 B.n188 B.n155 163.367
R783 B.n189 B.n188 163.367
R784 B.n284 B.t1 124.279
R785 B.n46 B.t8 124.279
R786 B.n126 B.t10 124.26
R787 B.n38 B.t5 124.26
R788 B.n285 B.t2 111.868
R789 B.n47 B.t7 111.868
R790 B.n127 B.t11 111.847
R791 B.n39 B.t4 111.847
R792 B.n270 B.n127 59.5399
R793 B.n286 B.n285 59.5399
R794 B.n508 B.n47 59.5399
R795 B.n40 B.n39 59.5399
R796 B.n604 B.n603 30.7517
R797 B.n429 B.n74 30.7517
R798 B.n369 B.n94 30.7517
R799 B.n191 B.n154 30.7517
R800 B B.n633 18.0485
R801 B.n127 B.n126 12.4126
R802 B.n285 B.n284 12.4126
R803 B.n47 B.n46 12.4126
R804 B.n39 B.n38 12.4126
R805 B.n605 B.n604 10.6151
R806 B.n605 B.n10 10.6151
R807 B.n609 B.n10 10.6151
R808 B.n610 B.n609 10.6151
R809 B.n611 B.n610 10.6151
R810 B.n611 B.n8 10.6151
R811 B.n615 B.n8 10.6151
R812 B.n616 B.n615 10.6151
R813 B.n617 B.n616 10.6151
R814 B.n617 B.n6 10.6151
R815 B.n621 B.n6 10.6151
R816 B.n622 B.n621 10.6151
R817 B.n623 B.n622 10.6151
R818 B.n623 B.n4 10.6151
R819 B.n627 B.n4 10.6151
R820 B.n628 B.n627 10.6151
R821 B.n629 B.n628 10.6151
R822 B.n629 B.n0 10.6151
R823 B.n603 B.n12 10.6151
R824 B.n599 B.n12 10.6151
R825 B.n599 B.n598 10.6151
R826 B.n598 B.n597 10.6151
R827 B.n597 B.n14 10.6151
R828 B.n593 B.n14 10.6151
R829 B.n593 B.n592 10.6151
R830 B.n592 B.n591 10.6151
R831 B.n591 B.n16 10.6151
R832 B.n587 B.n16 10.6151
R833 B.n587 B.n586 10.6151
R834 B.n586 B.n585 10.6151
R835 B.n585 B.n18 10.6151
R836 B.n581 B.n18 10.6151
R837 B.n581 B.n580 10.6151
R838 B.n580 B.n579 10.6151
R839 B.n579 B.n20 10.6151
R840 B.n575 B.n20 10.6151
R841 B.n575 B.n574 10.6151
R842 B.n574 B.n573 10.6151
R843 B.n573 B.n22 10.6151
R844 B.n569 B.n22 10.6151
R845 B.n569 B.n568 10.6151
R846 B.n568 B.n567 10.6151
R847 B.n567 B.n24 10.6151
R848 B.n563 B.n24 10.6151
R849 B.n563 B.n562 10.6151
R850 B.n562 B.n561 10.6151
R851 B.n561 B.n26 10.6151
R852 B.n557 B.n26 10.6151
R853 B.n557 B.n556 10.6151
R854 B.n556 B.n555 10.6151
R855 B.n555 B.n28 10.6151
R856 B.n551 B.n28 10.6151
R857 B.n551 B.n550 10.6151
R858 B.n550 B.n549 10.6151
R859 B.n549 B.n30 10.6151
R860 B.n545 B.n30 10.6151
R861 B.n545 B.n544 10.6151
R862 B.n544 B.n543 10.6151
R863 B.n543 B.n32 10.6151
R864 B.n539 B.n32 10.6151
R865 B.n539 B.n538 10.6151
R866 B.n538 B.n537 10.6151
R867 B.n537 B.n34 10.6151
R868 B.n533 B.n34 10.6151
R869 B.n533 B.n532 10.6151
R870 B.n532 B.n531 10.6151
R871 B.n531 B.n36 10.6151
R872 B.n527 B.n36 10.6151
R873 B.n527 B.n526 10.6151
R874 B.n526 B.n525 10.6151
R875 B.n522 B.n521 10.6151
R876 B.n521 B.n520 10.6151
R877 B.n520 B.n42 10.6151
R878 B.n516 B.n42 10.6151
R879 B.n516 B.n515 10.6151
R880 B.n515 B.n514 10.6151
R881 B.n514 B.n44 10.6151
R882 B.n510 B.n44 10.6151
R883 B.n510 B.n509 10.6151
R884 B.n507 B.n48 10.6151
R885 B.n503 B.n48 10.6151
R886 B.n503 B.n502 10.6151
R887 B.n502 B.n501 10.6151
R888 B.n501 B.n50 10.6151
R889 B.n497 B.n50 10.6151
R890 B.n497 B.n496 10.6151
R891 B.n496 B.n495 10.6151
R892 B.n495 B.n52 10.6151
R893 B.n491 B.n52 10.6151
R894 B.n491 B.n490 10.6151
R895 B.n490 B.n489 10.6151
R896 B.n489 B.n54 10.6151
R897 B.n485 B.n54 10.6151
R898 B.n485 B.n484 10.6151
R899 B.n484 B.n483 10.6151
R900 B.n483 B.n56 10.6151
R901 B.n479 B.n56 10.6151
R902 B.n479 B.n478 10.6151
R903 B.n478 B.n477 10.6151
R904 B.n477 B.n58 10.6151
R905 B.n473 B.n58 10.6151
R906 B.n473 B.n472 10.6151
R907 B.n472 B.n471 10.6151
R908 B.n471 B.n60 10.6151
R909 B.n467 B.n60 10.6151
R910 B.n467 B.n466 10.6151
R911 B.n466 B.n465 10.6151
R912 B.n465 B.n62 10.6151
R913 B.n461 B.n62 10.6151
R914 B.n461 B.n460 10.6151
R915 B.n460 B.n459 10.6151
R916 B.n459 B.n64 10.6151
R917 B.n455 B.n64 10.6151
R918 B.n455 B.n454 10.6151
R919 B.n454 B.n453 10.6151
R920 B.n453 B.n66 10.6151
R921 B.n449 B.n66 10.6151
R922 B.n449 B.n448 10.6151
R923 B.n448 B.n447 10.6151
R924 B.n447 B.n68 10.6151
R925 B.n443 B.n68 10.6151
R926 B.n443 B.n442 10.6151
R927 B.n442 B.n441 10.6151
R928 B.n441 B.n70 10.6151
R929 B.n437 B.n70 10.6151
R930 B.n437 B.n436 10.6151
R931 B.n436 B.n435 10.6151
R932 B.n435 B.n72 10.6151
R933 B.n431 B.n72 10.6151
R934 B.n431 B.n430 10.6151
R935 B.n430 B.n429 10.6151
R936 B.n425 B.n74 10.6151
R937 B.n425 B.n424 10.6151
R938 B.n424 B.n423 10.6151
R939 B.n423 B.n76 10.6151
R940 B.n419 B.n76 10.6151
R941 B.n419 B.n418 10.6151
R942 B.n418 B.n417 10.6151
R943 B.n417 B.n78 10.6151
R944 B.n413 B.n78 10.6151
R945 B.n413 B.n412 10.6151
R946 B.n412 B.n411 10.6151
R947 B.n411 B.n80 10.6151
R948 B.n407 B.n80 10.6151
R949 B.n407 B.n406 10.6151
R950 B.n406 B.n405 10.6151
R951 B.n405 B.n82 10.6151
R952 B.n401 B.n82 10.6151
R953 B.n401 B.n400 10.6151
R954 B.n400 B.n399 10.6151
R955 B.n399 B.n84 10.6151
R956 B.n395 B.n84 10.6151
R957 B.n395 B.n394 10.6151
R958 B.n394 B.n393 10.6151
R959 B.n393 B.n86 10.6151
R960 B.n389 B.n86 10.6151
R961 B.n389 B.n388 10.6151
R962 B.n388 B.n387 10.6151
R963 B.n387 B.n88 10.6151
R964 B.n383 B.n88 10.6151
R965 B.n383 B.n382 10.6151
R966 B.n382 B.n381 10.6151
R967 B.n381 B.n90 10.6151
R968 B.n377 B.n90 10.6151
R969 B.n377 B.n376 10.6151
R970 B.n376 B.n375 10.6151
R971 B.n375 B.n92 10.6151
R972 B.n371 B.n92 10.6151
R973 B.n371 B.n370 10.6151
R974 B.n370 B.n369 10.6151
R975 B.n163 B.n1 10.6151
R976 B.n163 B.n162 10.6151
R977 B.n167 B.n162 10.6151
R978 B.n168 B.n167 10.6151
R979 B.n169 B.n168 10.6151
R980 B.n169 B.n160 10.6151
R981 B.n173 B.n160 10.6151
R982 B.n174 B.n173 10.6151
R983 B.n175 B.n174 10.6151
R984 B.n175 B.n158 10.6151
R985 B.n179 B.n158 10.6151
R986 B.n180 B.n179 10.6151
R987 B.n181 B.n180 10.6151
R988 B.n181 B.n156 10.6151
R989 B.n185 B.n156 10.6151
R990 B.n186 B.n185 10.6151
R991 B.n187 B.n186 10.6151
R992 B.n187 B.n154 10.6151
R993 B.n192 B.n191 10.6151
R994 B.n193 B.n192 10.6151
R995 B.n193 B.n152 10.6151
R996 B.n197 B.n152 10.6151
R997 B.n198 B.n197 10.6151
R998 B.n199 B.n198 10.6151
R999 B.n199 B.n150 10.6151
R1000 B.n203 B.n150 10.6151
R1001 B.n204 B.n203 10.6151
R1002 B.n205 B.n204 10.6151
R1003 B.n205 B.n148 10.6151
R1004 B.n209 B.n148 10.6151
R1005 B.n210 B.n209 10.6151
R1006 B.n211 B.n210 10.6151
R1007 B.n211 B.n146 10.6151
R1008 B.n215 B.n146 10.6151
R1009 B.n216 B.n215 10.6151
R1010 B.n217 B.n216 10.6151
R1011 B.n217 B.n144 10.6151
R1012 B.n221 B.n144 10.6151
R1013 B.n222 B.n221 10.6151
R1014 B.n223 B.n222 10.6151
R1015 B.n223 B.n142 10.6151
R1016 B.n227 B.n142 10.6151
R1017 B.n228 B.n227 10.6151
R1018 B.n229 B.n228 10.6151
R1019 B.n229 B.n140 10.6151
R1020 B.n233 B.n140 10.6151
R1021 B.n234 B.n233 10.6151
R1022 B.n235 B.n234 10.6151
R1023 B.n235 B.n138 10.6151
R1024 B.n239 B.n138 10.6151
R1025 B.n240 B.n239 10.6151
R1026 B.n241 B.n240 10.6151
R1027 B.n241 B.n136 10.6151
R1028 B.n245 B.n136 10.6151
R1029 B.n246 B.n245 10.6151
R1030 B.n247 B.n246 10.6151
R1031 B.n247 B.n134 10.6151
R1032 B.n251 B.n134 10.6151
R1033 B.n252 B.n251 10.6151
R1034 B.n253 B.n252 10.6151
R1035 B.n253 B.n132 10.6151
R1036 B.n257 B.n132 10.6151
R1037 B.n258 B.n257 10.6151
R1038 B.n259 B.n258 10.6151
R1039 B.n259 B.n130 10.6151
R1040 B.n263 B.n130 10.6151
R1041 B.n264 B.n263 10.6151
R1042 B.n265 B.n264 10.6151
R1043 B.n265 B.n128 10.6151
R1044 B.n269 B.n128 10.6151
R1045 B.n272 B.n271 10.6151
R1046 B.n272 B.n124 10.6151
R1047 B.n276 B.n124 10.6151
R1048 B.n277 B.n276 10.6151
R1049 B.n278 B.n277 10.6151
R1050 B.n278 B.n122 10.6151
R1051 B.n282 B.n122 10.6151
R1052 B.n283 B.n282 10.6151
R1053 B.n287 B.n283 10.6151
R1054 B.n291 B.n120 10.6151
R1055 B.n292 B.n291 10.6151
R1056 B.n293 B.n292 10.6151
R1057 B.n293 B.n118 10.6151
R1058 B.n297 B.n118 10.6151
R1059 B.n298 B.n297 10.6151
R1060 B.n299 B.n298 10.6151
R1061 B.n299 B.n116 10.6151
R1062 B.n303 B.n116 10.6151
R1063 B.n304 B.n303 10.6151
R1064 B.n305 B.n304 10.6151
R1065 B.n305 B.n114 10.6151
R1066 B.n309 B.n114 10.6151
R1067 B.n310 B.n309 10.6151
R1068 B.n311 B.n310 10.6151
R1069 B.n311 B.n112 10.6151
R1070 B.n315 B.n112 10.6151
R1071 B.n316 B.n315 10.6151
R1072 B.n317 B.n316 10.6151
R1073 B.n317 B.n110 10.6151
R1074 B.n321 B.n110 10.6151
R1075 B.n322 B.n321 10.6151
R1076 B.n323 B.n322 10.6151
R1077 B.n323 B.n108 10.6151
R1078 B.n327 B.n108 10.6151
R1079 B.n328 B.n327 10.6151
R1080 B.n329 B.n328 10.6151
R1081 B.n329 B.n106 10.6151
R1082 B.n333 B.n106 10.6151
R1083 B.n334 B.n333 10.6151
R1084 B.n335 B.n334 10.6151
R1085 B.n335 B.n104 10.6151
R1086 B.n339 B.n104 10.6151
R1087 B.n340 B.n339 10.6151
R1088 B.n341 B.n340 10.6151
R1089 B.n341 B.n102 10.6151
R1090 B.n345 B.n102 10.6151
R1091 B.n346 B.n345 10.6151
R1092 B.n347 B.n346 10.6151
R1093 B.n347 B.n100 10.6151
R1094 B.n351 B.n100 10.6151
R1095 B.n352 B.n351 10.6151
R1096 B.n353 B.n352 10.6151
R1097 B.n353 B.n98 10.6151
R1098 B.n357 B.n98 10.6151
R1099 B.n358 B.n357 10.6151
R1100 B.n359 B.n358 10.6151
R1101 B.n359 B.n96 10.6151
R1102 B.n363 B.n96 10.6151
R1103 B.n364 B.n363 10.6151
R1104 B.n365 B.n364 10.6151
R1105 B.n365 B.n94 10.6151
R1106 B.n525 B.n40 9.36635
R1107 B.n508 B.n507 9.36635
R1108 B.n270 B.n269 9.36635
R1109 B.n286 B.n120 9.36635
R1110 B.n633 B.n0 8.11757
R1111 B.n633 B.n1 8.11757
R1112 B.n522 B.n40 1.24928
R1113 B.n509 B.n508 1.24928
R1114 B.n271 B.n270 1.24928
R1115 B.n287 B.n286 1.24928
C0 VDD1 VN 0.147686f
C1 w_n1738_n4152# VP 3.3155f
C2 VTAIL B 3.0909f
C3 B VDD2 1.83439f
C4 VTAIL w_n1738_n4152# 3.68416f
C5 B VDD1 1.80502f
C6 w_n1738_n4152# VDD2 2.18033f
C7 w_n1738_n4152# VDD1 2.15571f
C8 VTAIL VP 4.73622f
C9 B VN 0.740957f
C10 VDD2 VP 0.292309f
C11 w_n1738_n4152# VN 3.09629f
C12 VDD1 VP 5.4099f
C13 VTAIL VDD2 26.6618f
C14 VTAIL VDD1 26.634699f
C15 B w_n1738_n4152# 7.81058f
C16 VN VP 5.75072f
C17 VDD1 VDD2 0.732832f
C18 VTAIL VN 4.72125f
C19 B VP 1.09694f
C20 VDD2 VN 5.27205f
C21 VDD2 VSUBS 1.595016f
C22 VDD1 VSUBS 1.150298f
C23 VTAIL VSUBS 0.649368f
C24 VN VSUBS 5.00641f
C25 VP VSUBS 1.480785f
C26 B VSUBS 2.850952f
C27 w_n1738_n4152# VSUBS 88.4086f
C28 B.n0 VSUBS 0.006519f
C29 B.n1 VSUBS 0.006519f
C30 B.n2 VSUBS 0.009642f
C31 B.n3 VSUBS 0.007389f
C32 B.n4 VSUBS 0.007389f
C33 B.n5 VSUBS 0.007389f
C34 B.n6 VSUBS 0.007389f
C35 B.n7 VSUBS 0.007389f
C36 B.n8 VSUBS 0.007389f
C37 B.n9 VSUBS 0.007389f
C38 B.n10 VSUBS 0.007389f
C39 B.n11 VSUBS 0.016206f
C40 B.n12 VSUBS 0.007389f
C41 B.n13 VSUBS 0.007389f
C42 B.n14 VSUBS 0.007389f
C43 B.n15 VSUBS 0.007389f
C44 B.n16 VSUBS 0.007389f
C45 B.n17 VSUBS 0.007389f
C46 B.n18 VSUBS 0.007389f
C47 B.n19 VSUBS 0.007389f
C48 B.n20 VSUBS 0.007389f
C49 B.n21 VSUBS 0.007389f
C50 B.n22 VSUBS 0.007389f
C51 B.n23 VSUBS 0.007389f
C52 B.n24 VSUBS 0.007389f
C53 B.n25 VSUBS 0.007389f
C54 B.n26 VSUBS 0.007389f
C55 B.n27 VSUBS 0.007389f
C56 B.n28 VSUBS 0.007389f
C57 B.n29 VSUBS 0.007389f
C58 B.n30 VSUBS 0.007389f
C59 B.n31 VSUBS 0.007389f
C60 B.n32 VSUBS 0.007389f
C61 B.n33 VSUBS 0.007389f
C62 B.n34 VSUBS 0.007389f
C63 B.n35 VSUBS 0.007389f
C64 B.n36 VSUBS 0.007389f
C65 B.n37 VSUBS 0.007389f
C66 B.t4 VSUBS 0.562149f
C67 B.t5 VSUBS 0.567688f
C68 B.t3 VSUBS 0.202937f
C69 B.n38 VSUBS 0.119927f
C70 B.n39 VSUBS 0.06599f
C71 B.n40 VSUBS 0.017119f
C72 B.n41 VSUBS 0.007389f
C73 B.n42 VSUBS 0.007389f
C74 B.n43 VSUBS 0.007389f
C75 B.n44 VSUBS 0.007389f
C76 B.n45 VSUBS 0.007389f
C77 B.t7 VSUBS 0.562132f
C78 B.t8 VSUBS 0.567672f
C79 B.t6 VSUBS 0.202937f
C80 B.n46 VSUBS 0.119943f
C81 B.n47 VSUBS 0.066007f
C82 B.n48 VSUBS 0.007389f
C83 B.n49 VSUBS 0.007389f
C84 B.n50 VSUBS 0.007389f
C85 B.n51 VSUBS 0.007389f
C86 B.n52 VSUBS 0.007389f
C87 B.n53 VSUBS 0.007389f
C88 B.n54 VSUBS 0.007389f
C89 B.n55 VSUBS 0.007389f
C90 B.n56 VSUBS 0.007389f
C91 B.n57 VSUBS 0.007389f
C92 B.n58 VSUBS 0.007389f
C93 B.n59 VSUBS 0.007389f
C94 B.n60 VSUBS 0.007389f
C95 B.n61 VSUBS 0.007389f
C96 B.n62 VSUBS 0.007389f
C97 B.n63 VSUBS 0.007389f
C98 B.n64 VSUBS 0.007389f
C99 B.n65 VSUBS 0.007389f
C100 B.n66 VSUBS 0.007389f
C101 B.n67 VSUBS 0.007389f
C102 B.n68 VSUBS 0.007389f
C103 B.n69 VSUBS 0.007389f
C104 B.n70 VSUBS 0.007389f
C105 B.n71 VSUBS 0.007389f
C106 B.n72 VSUBS 0.007389f
C107 B.n73 VSUBS 0.007389f
C108 B.n74 VSUBS 0.016206f
C109 B.n75 VSUBS 0.007389f
C110 B.n76 VSUBS 0.007389f
C111 B.n77 VSUBS 0.007389f
C112 B.n78 VSUBS 0.007389f
C113 B.n79 VSUBS 0.007389f
C114 B.n80 VSUBS 0.007389f
C115 B.n81 VSUBS 0.007389f
C116 B.n82 VSUBS 0.007389f
C117 B.n83 VSUBS 0.007389f
C118 B.n84 VSUBS 0.007389f
C119 B.n85 VSUBS 0.007389f
C120 B.n86 VSUBS 0.007389f
C121 B.n87 VSUBS 0.007389f
C122 B.n88 VSUBS 0.007389f
C123 B.n89 VSUBS 0.007389f
C124 B.n90 VSUBS 0.007389f
C125 B.n91 VSUBS 0.007389f
C126 B.n92 VSUBS 0.007389f
C127 B.n93 VSUBS 0.007389f
C128 B.n94 VSUBS 0.016116f
C129 B.n95 VSUBS 0.007389f
C130 B.n96 VSUBS 0.007389f
C131 B.n97 VSUBS 0.007389f
C132 B.n98 VSUBS 0.007389f
C133 B.n99 VSUBS 0.007389f
C134 B.n100 VSUBS 0.007389f
C135 B.n101 VSUBS 0.007389f
C136 B.n102 VSUBS 0.007389f
C137 B.n103 VSUBS 0.007389f
C138 B.n104 VSUBS 0.007389f
C139 B.n105 VSUBS 0.007389f
C140 B.n106 VSUBS 0.007389f
C141 B.n107 VSUBS 0.007389f
C142 B.n108 VSUBS 0.007389f
C143 B.n109 VSUBS 0.007389f
C144 B.n110 VSUBS 0.007389f
C145 B.n111 VSUBS 0.007389f
C146 B.n112 VSUBS 0.007389f
C147 B.n113 VSUBS 0.007389f
C148 B.n114 VSUBS 0.007389f
C149 B.n115 VSUBS 0.007389f
C150 B.n116 VSUBS 0.007389f
C151 B.n117 VSUBS 0.007389f
C152 B.n118 VSUBS 0.007389f
C153 B.n119 VSUBS 0.007389f
C154 B.n120 VSUBS 0.006954f
C155 B.n121 VSUBS 0.007389f
C156 B.n122 VSUBS 0.007389f
C157 B.n123 VSUBS 0.007389f
C158 B.n124 VSUBS 0.007389f
C159 B.n125 VSUBS 0.007389f
C160 B.t11 VSUBS 0.562149f
C161 B.t10 VSUBS 0.567688f
C162 B.t9 VSUBS 0.202937f
C163 B.n126 VSUBS 0.119927f
C164 B.n127 VSUBS 0.06599f
C165 B.n128 VSUBS 0.007389f
C166 B.n129 VSUBS 0.007389f
C167 B.n130 VSUBS 0.007389f
C168 B.n131 VSUBS 0.007389f
C169 B.n132 VSUBS 0.007389f
C170 B.n133 VSUBS 0.007389f
C171 B.n134 VSUBS 0.007389f
C172 B.n135 VSUBS 0.007389f
C173 B.n136 VSUBS 0.007389f
C174 B.n137 VSUBS 0.007389f
C175 B.n138 VSUBS 0.007389f
C176 B.n139 VSUBS 0.007389f
C177 B.n140 VSUBS 0.007389f
C178 B.n141 VSUBS 0.007389f
C179 B.n142 VSUBS 0.007389f
C180 B.n143 VSUBS 0.007389f
C181 B.n144 VSUBS 0.007389f
C182 B.n145 VSUBS 0.007389f
C183 B.n146 VSUBS 0.007389f
C184 B.n147 VSUBS 0.007389f
C185 B.n148 VSUBS 0.007389f
C186 B.n149 VSUBS 0.007389f
C187 B.n150 VSUBS 0.007389f
C188 B.n151 VSUBS 0.007389f
C189 B.n152 VSUBS 0.007389f
C190 B.n153 VSUBS 0.007389f
C191 B.n154 VSUBS 0.016206f
C192 B.n155 VSUBS 0.007389f
C193 B.n156 VSUBS 0.007389f
C194 B.n157 VSUBS 0.007389f
C195 B.n158 VSUBS 0.007389f
C196 B.n159 VSUBS 0.007389f
C197 B.n160 VSUBS 0.007389f
C198 B.n161 VSUBS 0.007389f
C199 B.n162 VSUBS 0.007389f
C200 B.n163 VSUBS 0.007389f
C201 B.n164 VSUBS 0.007389f
C202 B.n165 VSUBS 0.007389f
C203 B.n166 VSUBS 0.007389f
C204 B.n167 VSUBS 0.007389f
C205 B.n168 VSUBS 0.007389f
C206 B.n169 VSUBS 0.007389f
C207 B.n170 VSUBS 0.007389f
C208 B.n171 VSUBS 0.007389f
C209 B.n172 VSUBS 0.007389f
C210 B.n173 VSUBS 0.007389f
C211 B.n174 VSUBS 0.007389f
C212 B.n175 VSUBS 0.007389f
C213 B.n176 VSUBS 0.007389f
C214 B.n177 VSUBS 0.007389f
C215 B.n178 VSUBS 0.007389f
C216 B.n179 VSUBS 0.007389f
C217 B.n180 VSUBS 0.007389f
C218 B.n181 VSUBS 0.007389f
C219 B.n182 VSUBS 0.007389f
C220 B.n183 VSUBS 0.007389f
C221 B.n184 VSUBS 0.007389f
C222 B.n185 VSUBS 0.007389f
C223 B.n186 VSUBS 0.007389f
C224 B.n187 VSUBS 0.007389f
C225 B.n188 VSUBS 0.007389f
C226 B.n189 VSUBS 0.016206f
C227 B.n190 VSUBS 0.017043f
C228 B.n191 VSUBS 0.017043f
C229 B.n192 VSUBS 0.007389f
C230 B.n193 VSUBS 0.007389f
C231 B.n194 VSUBS 0.007389f
C232 B.n195 VSUBS 0.007389f
C233 B.n196 VSUBS 0.007389f
C234 B.n197 VSUBS 0.007389f
C235 B.n198 VSUBS 0.007389f
C236 B.n199 VSUBS 0.007389f
C237 B.n200 VSUBS 0.007389f
C238 B.n201 VSUBS 0.007389f
C239 B.n202 VSUBS 0.007389f
C240 B.n203 VSUBS 0.007389f
C241 B.n204 VSUBS 0.007389f
C242 B.n205 VSUBS 0.007389f
C243 B.n206 VSUBS 0.007389f
C244 B.n207 VSUBS 0.007389f
C245 B.n208 VSUBS 0.007389f
C246 B.n209 VSUBS 0.007389f
C247 B.n210 VSUBS 0.007389f
C248 B.n211 VSUBS 0.007389f
C249 B.n212 VSUBS 0.007389f
C250 B.n213 VSUBS 0.007389f
C251 B.n214 VSUBS 0.007389f
C252 B.n215 VSUBS 0.007389f
C253 B.n216 VSUBS 0.007389f
C254 B.n217 VSUBS 0.007389f
C255 B.n218 VSUBS 0.007389f
C256 B.n219 VSUBS 0.007389f
C257 B.n220 VSUBS 0.007389f
C258 B.n221 VSUBS 0.007389f
C259 B.n222 VSUBS 0.007389f
C260 B.n223 VSUBS 0.007389f
C261 B.n224 VSUBS 0.007389f
C262 B.n225 VSUBS 0.007389f
C263 B.n226 VSUBS 0.007389f
C264 B.n227 VSUBS 0.007389f
C265 B.n228 VSUBS 0.007389f
C266 B.n229 VSUBS 0.007389f
C267 B.n230 VSUBS 0.007389f
C268 B.n231 VSUBS 0.007389f
C269 B.n232 VSUBS 0.007389f
C270 B.n233 VSUBS 0.007389f
C271 B.n234 VSUBS 0.007389f
C272 B.n235 VSUBS 0.007389f
C273 B.n236 VSUBS 0.007389f
C274 B.n237 VSUBS 0.007389f
C275 B.n238 VSUBS 0.007389f
C276 B.n239 VSUBS 0.007389f
C277 B.n240 VSUBS 0.007389f
C278 B.n241 VSUBS 0.007389f
C279 B.n242 VSUBS 0.007389f
C280 B.n243 VSUBS 0.007389f
C281 B.n244 VSUBS 0.007389f
C282 B.n245 VSUBS 0.007389f
C283 B.n246 VSUBS 0.007389f
C284 B.n247 VSUBS 0.007389f
C285 B.n248 VSUBS 0.007389f
C286 B.n249 VSUBS 0.007389f
C287 B.n250 VSUBS 0.007389f
C288 B.n251 VSUBS 0.007389f
C289 B.n252 VSUBS 0.007389f
C290 B.n253 VSUBS 0.007389f
C291 B.n254 VSUBS 0.007389f
C292 B.n255 VSUBS 0.007389f
C293 B.n256 VSUBS 0.007389f
C294 B.n257 VSUBS 0.007389f
C295 B.n258 VSUBS 0.007389f
C296 B.n259 VSUBS 0.007389f
C297 B.n260 VSUBS 0.007389f
C298 B.n261 VSUBS 0.007389f
C299 B.n262 VSUBS 0.007389f
C300 B.n263 VSUBS 0.007389f
C301 B.n264 VSUBS 0.007389f
C302 B.n265 VSUBS 0.007389f
C303 B.n266 VSUBS 0.007389f
C304 B.n267 VSUBS 0.007389f
C305 B.n268 VSUBS 0.007389f
C306 B.n269 VSUBS 0.006954f
C307 B.n270 VSUBS 0.017119f
C308 B.n271 VSUBS 0.004129f
C309 B.n272 VSUBS 0.007389f
C310 B.n273 VSUBS 0.007389f
C311 B.n274 VSUBS 0.007389f
C312 B.n275 VSUBS 0.007389f
C313 B.n276 VSUBS 0.007389f
C314 B.n277 VSUBS 0.007389f
C315 B.n278 VSUBS 0.007389f
C316 B.n279 VSUBS 0.007389f
C317 B.n280 VSUBS 0.007389f
C318 B.n281 VSUBS 0.007389f
C319 B.n282 VSUBS 0.007389f
C320 B.n283 VSUBS 0.007389f
C321 B.t2 VSUBS 0.562132f
C322 B.t1 VSUBS 0.567672f
C323 B.t0 VSUBS 0.202937f
C324 B.n284 VSUBS 0.119943f
C325 B.n285 VSUBS 0.066007f
C326 B.n286 VSUBS 0.017119f
C327 B.n287 VSUBS 0.004129f
C328 B.n288 VSUBS 0.007389f
C329 B.n289 VSUBS 0.007389f
C330 B.n290 VSUBS 0.007389f
C331 B.n291 VSUBS 0.007389f
C332 B.n292 VSUBS 0.007389f
C333 B.n293 VSUBS 0.007389f
C334 B.n294 VSUBS 0.007389f
C335 B.n295 VSUBS 0.007389f
C336 B.n296 VSUBS 0.007389f
C337 B.n297 VSUBS 0.007389f
C338 B.n298 VSUBS 0.007389f
C339 B.n299 VSUBS 0.007389f
C340 B.n300 VSUBS 0.007389f
C341 B.n301 VSUBS 0.007389f
C342 B.n302 VSUBS 0.007389f
C343 B.n303 VSUBS 0.007389f
C344 B.n304 VSUBS 0.007389f
C345 B.n305 VSUBS 0.007389f
C346 B.n306 VSUBS 0.007389f
C347 B.n307 VSUBS 0.007389f
C348 B.n308 VSUBS 0.007389f
C349 B.n309 VSUBS 0.007389f
C350 B.n310 VSUBS 0.007389f
C351 B.n311 VSUBS 0.007389f
C352 B.n312 VSUBS 0.007389f
C353 B.n313 VSUBS 0.007389f
C354 B.n314 VSUBS 0.007389f
C355 B.n315 VSUBS 0.007389f
C356 B.n316 VSUBS 0.007389f
C357 B.n317 VSUBS 0.007389f
C358 B.n318 VSUBS 0.007389f
C359 B.n319 VSUBS 0.007389f
C360 B.n320 VSUBS 0.007389f
C361 B.n321 VSUBS 0.007389f
C362 B.n322 VSUBS 0.007389f
C363 B.n323 VSUBS 0.007389f
C364 B.n324 VSUBS 0.007389f
C365 B.n325 VSUBS 0.007389f
C366 B.n326 VSUBS 0.007389f
C367 B.n327 VSUBS 0.007389f
C368 B.n328 VSUBS 0.007389f
C369 B.n329 VSUBS 0.007389f
C370 B.n330 VSUBS 0.007389f
C371 B.n331 VSUBS 0.007389f
C372 B.n332 VSUBS 0.007389f
C373 B.n333 VSUBS 0.007389f
C374 B.n334 VSUBS 0.007389f
C375 B.n335 VSUBS 0.007389f
C376 B.n336 VSUBS 0.007389f
C377 B.n337 VSUBS 0.007389f
C378 B.n338 VSUBS 0.007389f
C379 B.n339 VSUBS 0.007389f
C380 B.n340 VSUBS 0.007389f
C381 B.n341 VSUBS 0.007389f
C382 B.n342 VSUBS 0.007389f
C383 B.n343 VSUBS 0.007389f
C384 B.n344 VSUBS 0.007389f
C385 B.n345 VSUBS 0.007389f
C386 B.n346 VSUBS 0.007389f
C387 B.n347 VSUBS 0.007389f
C388 B.n348 VSUBS 0.007389f
C389 B.n349 VSUBS 0.007389f
C390 B.n350 VSUBS 0.007389f
C391 B.n351 VSUBS 0.007389f
C392 B.n352 VSUBS 0.007389f
C393 B.n353 VSUBS 0.007389f
C394 B.n354 VSUBS 0.007389f
C395 B.n355 VSUBS 0.007389f
C396 B.n356 VSUBS 0.007389f
C397 B.n357 VSUBS 0.007389f
C398 B.n358 VSUBS 0.007389f
C399 B.n359 VSUBS 0.007389f
C400 B.n360 VSUBS 0.007389f
C401 B.n361 VSUBS 0.007389f
C402 B.n362 VSUBS 0.007389f
C403 B.n363 VSUBS 0.007389f
C404 B.n364 VSUBS 0.007389f
C405 B.n365 VSUBS 0.007389f
C406 B.n366 VSUBS 0.007389f
C407 B.n367 VSUBS 0.017043f
C408 B.n368 VSUBS 0.016206f
C409 B.n369 VSUBS 0.017133f
C410 B.n370 VSUBS 0.007389f
C411 B.n371 VSUBS 0.007389f
C412 B.n372 VSUBS 0.007389f
C413 B.n373 VSUBS 0.007389f
C414 B.n374 VSUBS 0.007389f
C415 B.n375 VSUBS 0.007389f
C416 B.n376 VSUBS 0.007389f
C417 B.n377 VSUBS 0.007389f
C418 B.n378 VSUBS 0.007389f
C419 B.n379 VSUBS 0.007389f
C420 B.n380 VSUBS 0.007389f
C421 B.n381 VSUBS 0.007389f
C422 B.n382 VSUBS 0.007389f
C423 B.n383 VSUBS 0.007389f
C424 B.n384 VSUBS 0.007389f
C425 B.n385 VSUBS 0.007389f
C426 B.n386 VSUBS 0.007389f
C427 B.n387 VSUBS 0.007389f
C428 B.n388 VSUBS 0.007389f
C429 B.n389 VSUBS 0.007389f
C430 B.n390 VSUBS 0.007389f
C431 B.n391 VSUBS 0.007389f
C432 B.n392 VSUBS 0.007389f
C433 B.n393 VSUBS 0.007389f
C434 B.n394 VSUBS 0.007389f
C435 B.n395 VSUBS 0.007389f
C436 B.n396 VSUBS 0.007389f
C437 B.n397 VSUBS 0.007389f
C438 B.n398 VSUBS 0.007389f
C439 B.n399 VSUBS 0.007389f
C440 B.n400 VSUBS 0.007389f
C441 B.n401 VSUBS 0.007389f
C442 B.n402 VSUBS 0.007389f
C443 B.n403 VSUBS 0.007389f
C444 B.n404 VSUBS 0.007389f
C445 B.n405 VSUBS 0.007389f
C446 B.n406 VSUBS 0.007389f
C447 B.n407 VSUBS 0.007389f
C448 B.n408 VSUBS 0.007389f
C449 B.n409 VSUBS 0.007389f
C450 B.n410 VSUBS 0.007389f
C451 B.n411 VSUBS 0.007389f
C452 B.n412 VSUBS 0.007389f
C453 B.n413 VSUBS 0.007389f
C454 B.n414 VSUBS 0.007389f
C455 B.n415 VSUBS 0.007389f
C456 B.n416 VSUBS 0.007389f
C457 B.n417 VSUBS 0.007389f
C458 B.n418 VSUBS 0.007389f
C459 B.n419 VSUBS 0.007389f
C460 B.n420 VSUBS 0.007389f
C461 B.n421 VSUBS 0.007389f
C462 B.n422 VSUBS 0.007389f
C463 B.n423 VSUBS 0.007389f
C464 B.n424 VSUBS 0.007389f
C465 B.n425 VSUBS 0.007389f
C466 B.n426 VSUBS 0.007389f
C467 B.n427 VSUBS 0.016206f
C468 B.n428 VSUBS 0.017043f
C469 B.n429 VSUBS 0.017043f
C470 B.n430 VSUBS 0.007389f
C471 B.n431 VSUBS 0.007389f
C472 B.n432 VSUBS 0.007389f
C473 B.n433 VSUBS 0.007389f
C474 B.n434 VSUBS 0.007389f
C475 B.n435 VSUBS 0.007389f
C476 B.n436 VSUBS 0.007389f
C477 B.n437 VSUBS 0.007389f
C478 B.n438 VSUBS 0.007389f
C479 B.n439 VSUBS 0.007389f
C480 B.n440 VSUBS 0.007389f
C481 B.n441 VSUBS 0.007389f
C482 B.n442 VSUBS 0.007389f
C483 B.n443 VSUBS 0.007389f
C484 B.n444 VSUBS 0.007389f
C485 B.n445 VSUBS 0.007389f
C486 B.n446 VSUBS 0.007389f
C487 B.n447 VSUBS 0.007389f
C488 B.n448 VSUBS 0.007389f
C489 B.n449 VSUBS 0.007389f
C490 B.n450 VSUBS 0.007389f
C491 B.n451 VSUBS 0.007389f
C492 B.n452 VSUBS 0.007389f
C493 B.n453 VSUBS 0.007389f
C494 B.n454 VSUBS 0.007389f
C495 B.n455 VSUBS 0.007389f
C496 B.n456 VSUBS 0.007389f
C497 B.n457 VSUBS 0.007389f
C498 B.n458 VSUBS 0.007389f
C499 B.n459 VSUBS 0.007389f
C500 B.n460 VSUBS 0.007389f
C501 B.n461 VSUBS 0.007389f
C502 B.n462 VSUBS 0.007389f
C503 B.n463 VSUBS 0.007389f
C504 B.n464 VSUBS 0.007389f
C505 B.n465 VSUBS 0.007389f
C506 B.n466 VSUBS 0.007389f
C507 B.n467 VSUBS 0.007389f
C508 B.n468 VSUBS 0.007389f
C509 B.n469 VSUBS 0.007389f
C510 B.n470 VSUBS 0.007389f
C511 B.n471 VSUBS 0.007389f
C512 B.n472 VSUBS 0.007389f
C513 B.n473 VSUBS 0.007389f
C514 B.n474 VSUBS 0.007389f
C515 B.n475 VSUBS 0.007389f
C516 B.n476 VSUBS 0.007389f
C517 B.n477 VSUBS 0.007389f
C518 B.n478 VSUBS 0.007389f
C519 B.n479 VSUBS 0.007389f
C520 B.n480 VSUBS 0.007389f
C521 B.n481 VSUBS 0.007389f
C522 B.n482 VSUBS 0.007389f
C523 B.n483 VSUBS 0.007389f
C524 B.n484 VSUBS 0.007389f
C525 B.n485 VSUBS 0.007389f
C526 B.n486 VSUBS 0.007389f
C527 B.n487 VSUBS 0.007389f
C528 B.n488 VSUBS 0.007389f
C529 B.n489 VSUBS 0.007389f
C530 B.n490 VSUBS 0.007389f
C531 B.n491 VSUBS 0.007389f
C532 B.n492 VSUBS 0.007389f
C533 B.n493 VSUBS 0.007389f
C534 B.n494 VSUBS 0.007389f
C535 B.n495 VSUBS 0.007389f
C536 B.n496 VSUBS 0.007389f
C537 B.n497 VSUBS 0.007389f
C538 B.n498 VSUBS 0.007389f
C539 B.n499 VSUBS 0.007389f
C540 B.n500 VSUBS 0.007389f
C541 B.n501 VSUBS 0.007389f
C542 B.n502 VSUBS 0.007389f
C543 B.n503 VSUBS 0.007389f
C544 B.n504 VSUBS 0.007389f
C545 B.n505 VSUBS 0.007389f
C546 B.n506 VSUBS 0.007389f
C547 B.n507 VSUBS 0.006954f
C548 B.n508 VSUBS 0.017119f
C549 B.n509 VSUBS 0.004129f
C550 B.n510 VSUBS 0.007389f
C551 B.n511 VSUBS 0.007389f
C552 B.n512 VSUBS 0.007389f
C553 B.n513 VSUBS 0.007389f
C554 B.n514 VSUBS 0.007389f
C555 B.n515 VSUBS 0.007389f
C556 B.n516 VSUBS 0.007389f
C557 B.n517 VSUBS 0.007389f
C558 B.n518 VSUBS 0.007389f
C559 B.n519 VSUBS 0.007389f
C560 B.n520 VSUBS 0.007389f
C561 B.n521 VSUBS 0.007389f
C562 B.n522 VSUBS 0.004129f
C563 B.n523 VSUBS 0.007389f
C564 B.n524 VSUBS 0.007389f
C565 B.n525 VSUBS 0.006954f
C566 B.n526 VSUBS 0.007389f
C567 B.n527 VSUBS 0.007389f
C568 B.n528 VSUBS 0.007389f
C569 B.n529 VSUBS 0.007389f
C570 B.n530 VSUBS 0.007389f
C571 B.n531 VSUBS 0.007389f
C572 B.n532 VSUBS 0.007389f
C573 B.n533 VSUBS 0.007389f
C574 B.n534 VSUBS 0.007389f
C575 B.n535 VSUBS 0.007389f
C576 B.n536 VSUBS 0.007389f
C577 B.n537 VSUBS 0.007389f
C578 B.n538 VSUBS 0.007389f
C579 B.n539 VSUBS 0.007389f
C580 B.n540 VSUBS 0.007389f
C581 B.n541 VSUBS 0.007389f
C582 B.n542 VSUBS 0.007389f
C583 B.n543 VSUBS 0.007389f
C584 B.n544 VSUBS 0.007389f
C585 B.n545 VSUBS 0.007389f
C586 B.n546 VSUBS 0.007389f
C587 B.n547 VSUBS 0.007389f
C588 B.n548 VSUBS 0.007389f
C589 B.n549 VSUBS 0.007389f
C590 B.n550 VSUBS 0.007389f
C591 B.n551 VSUBS 0.007389f
C592 B.n552 VSUBS 0.007389f
C593 B.n553 VSUBS 0.007389f
C594 B.n554 VSUBS 0.007389f
C595 B.n555 VSUBS 0.007389f
C596 B.n556 VSUBS 0.007389f
C597 B.n557 VSUBS 0.007389f
C598 B.n558 VSUBS 0.007389f
C599 B.n559 VSUBS 0.007389f
C600 B.n560 VSUBS 0.007389f
C601 B.n561 VSUBS 0.007389f
C602 B.n562 VSUBS 0.007389f
C603 B.n563 VSUBS 0.007389f
C604 B.n564 VSUBS 0.007389f
C605 B.n565 VSUBS 0.007389f
C606 B.n566 VSUBS 0.007389f
C607 B.n567 VSUBS 0.007389f
C608 B.n568 VSUBS 0.007389f
C609 B.n569 VSUBS 0.007389f
C610 B.n570 VSUBS 0.007389f
C611 B.n571 VSUBS 0.007389f
C612 B.n572 VSUBS 0.007389f
C613 B.n573 VSUBS 0.007389f
C614 B.n574 VSUBS 0.007389f
C615 B.n575 VSUBS 0.007389f
C616 B.n576 VSUBS 0.007389f
C617 B.n577 VSUBS 0.007389f
C618 B.n578 VSUBS 0.007389f
C619 B.n579 VSUBS 0.007389f
C620 B.n580 VSUBS 0.007389f
C621 B.n581 VSUBS 0.007389f
C622 B.n582 VSUBS 0.007389f
C623 B.n583 VSUBS 0.007389f
C624 B.n584 VSUBS 0.007389f
C625 B.n585 VSUBS 0.007389f
C626 B.n586 VSUBS 0.007389f
C627 B.n587 VSUBS 0.007389f
C628 B.n588 VSUBS 0.007389f
C629 B.n589 VSUBS 0.007389f
C630 B.n590 VSUBS 0.007389f
C631 B.n591 VSUBS 0.007389f
C632 B.n592 VSUBS 0.007389f
C633 B.n593 VSUBS 0.007389f
C634 B.n594 VSUBS 0.007389f
C635 B.n595 VSUBS 0.007389f
C636 B.n596 VSUBS 0.007389f
C637 B.n597 VSUBS 0.007389f
C638 B.n598 VSUBS 0.007389f
C639 B.n599 VSUBS 0.007389f
C640 B.n600 VSUBS 0.007389f
C641 B.n601 VSUBS 0.007389f
C642 B.n602 VSUBS 0.017043f
C643 B.n603 VSUBS 0.017043f
C644 B.n604 VSUBS 0.016206f
C645 B.n605 VSUBS 0.007389f
C646 B.n606 VSUBS 0.007389f
C647 B.n607 VSUBS 0.007389f
C648 B.n608 VSUBS 0.007389f
C649 B.n609 VSUBS 0.007389f
C650 B.n610 VSUBS 0.007389f
C651 B.n611 VSUBS 0.007389f
C652 B.n612 VSUBS 0.007389f
C653 B.n613 VSUBS 0.007389f
C654 B.n614 VSUBS 0.007389f
C655 B.n615 VSUBS 0.007389f
C656 B.n616 VSUBS 0.007389f
C657 B.n617 VSUBS 0.007389f
C658 B.n618 VSUBS 0.007389f
C659 B.n619 VSUBS 0.007389f
C660 B.n620 VSUBS 0.007389f
C661 B.n621 VSUBS 0.007389f
C662 B.n622 VSUBS 0.007389f
C663 B.n623 VSUBS 0.007389f
C664 B.n624 VSUBS 0.007389f
C665 B.n625 VSUBS 0.007389f
C666 B.n626 VSUBS 0.007389f
C667 B.n627 VSUBS 0.007389f
C668 B.n628 VSUBS 0.007389f
C669 B.n629 VSUBS 0.007389f
C670 B.n630 VSUBS 0.007389f
C671 B.n631 VSUBS 0.009642f
C672 B.n632 VSUBS 0.010271f
C673 B.n633 VSUBS 0.020425f
C674 VDD2.t7 VSUBS 4.28354f
C675 VDD2.t1 VSUBS 0.400327f
C676 VDD2.t0 VSUBS 0.400327f
C677 VDD2.n0 VSUBS 3.2933f
C678 VDD2.n1 VSUBS 1.4386f
C679 VDD2.t3 VSUBS 0.400327f
C680 VDD2.t2 VSUBS 0.400327f
C681 VDD2.n2 VSUBS 3.2967f
C682 VDD2.n3 VSUBS 2.79369f
C683 VDD2.t8 VSUBS 4.27798f
C684 VDD2.n4 VSUBS 3.5942f
C685 VDD2.t5 VSUBS 0.400327f
C686 VDD2.t4 VSUBS 0.400327f
C687 VDD2.n5 VSUBS 3.2933f
C688 VDD2.n6 VSUBS 0.673516f
C689 VDD2.t9 VSUBS 0.400327f
C690 VDD2.t6 VSUBS 0.400327f
C691 VDD2.n7 VSUBS 3.29665f
C692 VN.n0 VSUBS 0.064004f
C693 VN.t6 VSUBS 0.891155f
C694 VN.t9 VSUBS 0.891155f
C695 VN.n1 VSUBS 0.026757f
C696 VN.t2 VSUBS 0.901306f
C697 VN.t8 VSUBS 0.891155f
C698 VN.n2 VSUBS 0.339271f
C699 VN.n3 VSUBS 0.359521f
C700 VN.n4 VSUBS 0.142517f
C701 VN.n5 VSUBS 0.064004f
C702 VN.n6 VSUBS 0.360503f
C703 VN.n7 VSUBS 0.026757f
C704 VN.n8 VSUBS 0.339271f
C705 VN.t7 VSUBS 0.901306f
C706 VN.n9 VSUBS 0.359428f
C707 VN.n10 VSUBS 0.049601f
C708 VN.n11 VSUBS 0.064004f
C709 VN.t1 VSUBS 0.901306f
C710 VN.t4 VSUBS 0.891155f
C711 VN.t5 VSUBS 0.891155f
C712 VN.n12 VSUBS 0.026757f
C713 VN.t0 VSUBS 0.891155f
C714 VN.n13 VSUBS 0.339271f
C715 VN.t3 VSUBS 0.901306f
C716 VN.n14 VSUBS 0.359521f
C717 VN.n15 VSUBS 0.142517f
C718 VN.n16 VSUBS 0.064004f
C719 VN.n17 VSUBS 0.360503f
C720 VN.n18 VSUBS 0.026757f
C721 VN.n19 VSUBS 0.339271f
C722 VN.n20 VSUBS 0.359428f
C723 VN.n21 VSUBS 2.86258f
C724 VDD1.t4 VSUBS 4.26889f
C725 VDD1.t0 VSUBS 0.398956f
C726 VDD1.t1 VSUBS 0.398956f
C727 VDD1.n0 VSUBS 3.28202f
C728 VDD1.n1 VSUBS 1.43635f
C729 VDD1.t7 VSUBS 4.26887f
C730 VDD1.t3 VSUBS 0.398956f
C731 VDD1.t5 VSUBS 0.398956f
C732 VDD1.n2 VSUBS 3.28202f
C733 VDD1.n3 VSUBS 1.43368f
C734 VDD1.t6 VSUBS 0.398956f
C735 VDD1.t2 VSUBS 0.398956f
C736 VDD1.n4 VSUBS 3.28541f
C737 VDD1.n5 VSUBS 2.87124f
C738 VDD1.t8 VSUBS 0.398956f
C739 VDD1.t9 VSUBS 0.398956f
C740 VDD1.n6 VSUBS 3.28201f
C741 VDD1.n7 VSUBS 3.5415f
C742 VTAIL.t4 VSUBS 0.422559f
C743 VTAIL.t2 VSUBS 0.422559f
C744 VTAIL.n0 VSUBS 3.29444f
C745 VTAIL.n1 VSUBS 0.897879f
C746 VTAIL.t11 VSUBS 4.30822f
C747 VTAIL.n2 VSUBS 1.04517f
C748 VTAIL.t14 VSUBS 0.422559f
C749 VTAIL.t18 VSUBS 0.422559f
C750 VTAIL.n3 VSUBS 3.29444f
C751 VTAIL.n4 VSUBS 0.885516f
C752 VTAIL.t19 VSUBS 0.422559f
C753 VTAIL.t13 VSUBS 0.422559f
C754 VTAIL.n5 VSUBS 3.29444f
C755 VTAIL.n6 VSUBS 2.88685f
C756 VTAIL.t6 VSUBS 0.422559f
C757 VTAIL.t9 VSUBS 0.422559f
C758 VTAIL.n7 VSUBS 3.29444f
C759 VTAIL.n8 VSUBS 2.88684f
C760 VTAIL.t3 VSUBS 0.422559f
C761 VTAIL.t1 VSUBS 0.422559f
C762 VTAIL.n9 VSUBS 3.29444f
C763 VTAIL.n10 VSUBS 0.88551f
C764 VTAIL.t8 VSUBS 4.30825f
C765 VTAIL.n11 VSUBS 1.04513f
C766 VTAIL.t15 VSUBS 0.422559f
C767 VTAIL.t12 VSUBS 0.422559f
C768 VTAIL.n12 VSUBS 3.29444f
C769 VTAIL.n13 VSUBS 0.906503f
C770 VTAIL.t10 VSUBS 0.422559f
C771 VTAIL.t16 VSUBS 0.422559f
C772 VTAIL.n14 VSUBS 3.29444f
C773 VTAIL.n15 VSUBS 0.88551f
C774 VTAIL.t17 VSUBS 4.30821f
C775 VTAIL.n16 VSUBS 2.96579f
C776 VTAIL.t5 VSUBS 4.30822f
C777 VTAIL.n17 VSUBS 2.96579f
C778 VTAIL.t7 VSUBS 0.422559f
C779 VTAIL.t0 VSUBS 0.422559f
C780 VTAIL.n18 VSUBS 3.29444f
C781 VTAIL.n19 VSUBS 0.834434f
C782 VP.n0 VSUBS 0.065331f
C783 VP.t3 VSUBS 0.90963f
C784 VP.t4 VSUBS 0.90963f
C785 VP.n1 VSUBS 0.027312f
C786 VP.n2 VSUBS 0.065331f
C787 VP.t1 VSUBS 0.90963f
C788 VP.t8 VSUBS 0.90963f
C789 VP.n3 VSUBS 0.027312f
C790 VP.t5 VSUBS 0.919992f
C791 VP.t9 VSUBS 0.90963f
C792 VP.n4 VSUBS 0.346305f
C793 VP.n5 VSUBS 0.366974f
C794 VP.n6 VSUBS 0.145471f
C795 VP.n7 VSUBS 0.065331f
C796 VP.n8 VSUBS 0.367977f
C797 VP.n9 VSUBS 0.027312f
C798 VP.n10 VSUBS 0.346305f
C799 VP.t0 VSUBS 0.919992f
C800 VP.n11 VSUBS 0.36688f
C801 VP.n12 VSUBS 2.87914f
C802 VP.t2 VSUBS 0.919992f
C803 VP.t6 VSUBS 0.90963f
C804 VP.n13 VSUBS 0.346305f
C805 VP.n14 VSUBS 0.36688f
C806 VP.n15 VSUBS 2.93272f
C807 VP.n16 VSUBS 0.065331f
C808 VP.n17 VSUBS 0.065331f
C809 VP.n18 VSUBS 0.367977f
C810 VP.n19 VSUBS 0.027312f
C811 VP.n20 VSUBS 0.346305f
C812 VP.t7 VSUBS 0.919992f
C813 VP.n21 VSUBS 0.36688f
C814 VP.n22 VSUBS 0.050629f
.ends

