* NGSPICE file created from diff_pair_sample_0690.ext - technology: sky130A

.subckt diff_pair_sample_0690 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.4719 ps=3.2 w=1.21 l=2.52
X1 VTAIL.t3 VP.t1 VDD1.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X2 VDD2.t9 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.4719 ps=3.2 w=1.21 l=2.52
X3 VDD1.t7 VP.t2 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0.19965 ps=1.54 w=1.21 l=2.52
X4 VDD2.t8 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0.19965 ps=1.54 w=1.21 l=2.52
X5 VTAIL.t0 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X6 VTAIL.t10 VP.t3 VDD1.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X7 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0 ps=0 w=1.21 l=2.52
X8 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0 ps=0 w=1.21 l=2.52
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0 ps=0 w=1.21 l=2.52
X10 VTAIL.t4 VP.t4 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X11 VDD1.t4 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X12 VTAIL.t16 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0 ps=0 w=1.21 l=2.52
X14 VDD2.t5 VN.t4 VTAIL.t19 B.t3 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X15 VTAIL.t17 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X16 VTAIL.t11 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X17 VDD2.t3 VN.t6 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.4719 ps=3.2 w=1.21 l=2.52
X18 VTAIL.t14 VN.t7 VDD2.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X19 VDD2.t1 VN.t8 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0.19965 ps=1.54 w=1.21 l=2.52
X20 VDD1.t2 VP.t7 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4719 pd=3.2 as=0.19965 ps=1.54 w=1.21 l=2.52
X21 VDD1.t1 VP.t8 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.4719 ps=3.2 w=1.21 l=2.52
X22 VDD2.t0 VN.t9 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
X23 VDD1.t0 VP.t9 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.19965 pd=1.54 as=0.19965 ps=1.54 w=1.21 l=2.52
R0 VP.n25 VP.n24 161.3
R1 VP.n26 VP.n21 161.3
R2 VP.n28 VP.n27 161.3
R3 VP.n29 VP.n20 161.3
R4 VP.n31 VP.n30 161.3
R5 VP.n32 VP.n19 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n18 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n17 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n13 161.3
R17 VP.n88 VP.n0 161.3
R18 VP.n87 VP.n86 161.3
R19 VP.n85 VP.n1 161.3
R20 VP.n84 VP.n83 161.3
R21 VP.n82 VP.n2 161.3
R22 VP.n81 VP.n80 161.3
R23 VP.n79 VP.n78 161.3
R24 VP.n77 VP.n4 161.3
R25 VP.n76 VP.n75 161.3
R26 VP.n74 VP.n5 161.3
R27 VP.n73 VP.n72 161.3
R28 VP.n71 VP.n6 161.3
R29 VP.n70 VP.n69 161.3
R30 VP.n68 VP.n7 161.3
R31 VP.n67 VP.n66 161.3
R32 VP.n65 VP.n8 161.3
R33 VP.n64 VP.n63 161.3
R34 VP.n62 VP.n61 161.3
R35 VP.n60 VP.n10 161.3
R36 VP.n59 VP.n58 161.3
R37 VP.n57 VP.n11 161.3
R38 VP.n56 VP.n55 161.3
R39 VP.n54 VP.n12 161.3
R40 VP.n53 VP.n52 100.969
R41 VP.n90 VP.n89 100.969
R42 VP.n51 VP.n50 100.969
R43 VP.n59 VP.n11 56.5193
R44 VP.n83 VP.n1 56.5193
R45 VP.n44 VP.n14 56.5193
R46 VP.n23 VP.n22 55.3127
R47 VP.n66 VP.n7 47.7779
R48 VP.n76 VP.n5 47.7779
R49 VP.n37 VP.n18 47.7779
R50 VP.n27 VP.n20 47.7779
R51 VP.n23 VP.t7 45.1187
R52 VP.n52 VP.n51 44.5034
R53 VP.n66 VP.n65 33.2089
R54 VP.n77 VP.n76 33.2089
R55 VP.n38 VP.n37 33.2089
R56 VP.n27 VP.n26 33.2089
R57 VP.n55 VP.n54 24.4675
R58 VP.n55 VP.n11 24.4675
R59 VP.n60 VP.n59 24.4675
R60 VP.n61 VP.n60 24.4675
R61 VP.n65 VP.n64 24.4675
R62 VP.n70 VP.n7 24.4675
R63 VP.n71 VP.n70 24.4675
R64 VP.n72 VP.n71 24.4675
R65 VP.n72 VP.n5 24.4675
R66 VP.n78 VP.n77 24.4675
R67 VP.n82 VP.n81 24.4675
R68 VP.n83 VP.n82 24.4675
R69 VP.n87 VP.n1 24.4675
R70 VP.n88 VP.n87 24.4675
R71 VP.n48 VP.n14 24.4675
R72 VP.n49 VP.n48 24.4675
R73 VP.n39 VP.n38 24.4675
R74 VP.n43 VP.n42 24.4675
R75 VP.n44 VP.n43 24.4675
R76 VP.n31 VP.n20 24.4675
R77 VP.n32 VP.n31 24.4675
R78 VP.n33 VP.n32 24.4675
R79 VP.n33 VP.n18 24.4675
R80 VP.n26 VP.n25 24.4675
R81 VP.n64 VP.n9 17.1274
R82 VP.n78 VP.n3 17.1274
R83 VP.n39 VP.n16 17.1274
R84 VP.n25 VP.n22 17.1274
R85 VP.n71 VP.t9 11.5723
R86 VP.n53 VP.t2 11.5723
R87 VP.n9 VP.t4 11.5723
R88 VP.n3 VP.t3 11.5723
R89 VP.n89 VP.t8 11.5723
R90 VP.n32 VP.t5 11.5723
R91 VP.n50 VP.t0 11.5723
R92 VP.n16 VP.t1 11.5723
R93 VP.n22 VP.t6 11.5723
R94 VP.n54 VP.n53 9.7873
R95 VP.n89 VP.n88 9.7873
R96 VP.n50 VP.n49 9.7873
R97 VP.n61 VP.n9 7.3406
R98 VP.n81 VP.n3 7.3406
R99 VP.n42 VP.n16 7.3406
R100 VP.n24 VP.n23 6.86339
R101 VP.n51 VP.n13 0.278367
R102 VP.n52 VP.n12 0.278367
R103 VP.n90 VP.n0 0.278367
R104 VP.n24 VP.n21 0.189894
R105 VP.n28 VP.n21 0.189894
R106 VP.n29 VP.n28 0.189894
R107 VP.n30 VP.n29 0.189894
R108 VP.n30 VP.n19 0.189894
R109 VP.n34 VP.n19 0.189894
R110 VP.n35 VP.n34 0.189894
R111 VP.n36 VP.n35 0.189894
R112 VP.n36 VP.n17 0.189894
R113 VP.n40 VP.n17 0.189894
R114 VP.n41 VP.n40 0.189894
R115 VP.n41 VP.n15 0.189894
R116 VP.n45 VP.n15 0.189894
R117 VP.n46 VP.n45 0.189894
R118 VP.n47 VP.n46 0.189894
R119 VP.n47 VP.n13 0.189894
R120 VP.n56 VP.n12 0.189894
R121 VP.n57 VP.n56 0.189894
R122 VP.n58 VP.n57 0.189894
R123 VP.n58 VP.n10 0.189894
R124 VP.n62 VP.n10 0.189894
R125 VP.n63 VP.n62 0.189894
R126 VP.n63 VP.n8 0.189894
R127 VP.n67 VP.n8 0.189894
R128 VP.n68 VP.n67 0.189894
R129 VP.n69 VP.n68 0.189894
R130 VP.n69 VP.n6 0.189894
R131 VP.n73 VP.n6 0.189894
R132 VP.n74 VP.n73 0.189894
R133 VP.n75 VP.n74 0.189894
R134 VP.n75 VP.n4 0.189894
R135 VP.n79 VP.n4 0.189894
R136 VP.n80 VP.n79 0.189894
R137 VP.n80 VP.n2 0.189894
R138 VP.n84 VP.n2 0.189894
R139 VP.n85 VP.n84 0.189894
R140 VP.n86 VP.n85 0.189894
R141 VP.n86 VP.n0 0.189894
R142 VP VP.n90 0.153454
R143 VTAIL.n17 VTAIL.t2 154.55
R144 VTAIL.n2 VTAIL.t8 154.55
R145 VTAIL.n16 VTAIL.t5 154.55
R146 VTAIL.n11 VTAIL.t15 154.55
R147 VTAIL.n19 VTAIL.n18 128.393
R148 VTAIL.n1 VTAIL.n0 128.393
R149 VTAIL.n4 VTAIL.n3 128.393
R150 VTAIL.n6 VTAIL.n5 128.393
R151 VTAIL.n15 VTAIL.n14 128.392
R152 VTAIL.n13 VTAIL.n12 128.392
R153 VTAIL.n10 VTAIL.n9 128.392
R154 VTAIL.n8 VTAIL.n7 128.392
R155 VTAIL.n8 VTAIL.n6 18.3238
R156 VTAIL.n18 VTAIL.t18 16.3641
R157 VTAIL.n18 VTAIL.t14 16.3641
R158 VTAIL.n0 VTAIL.t13 16.3641
R159 VTAIL.n0 VTAIL.t0 16.3641
R160 VTAIL.n3 VTAIL.t9 16.3641
R161 VTAIL.n3 VTAIL.t10 16.3641
R162 VTAIL.n5 VTAIL.t7 16.3641
R163 VTAIL.n5 VTAIL.t4 16.3641
R164 VTAIL.n14 VTAIL.t6 16.3641
R165 VTAIL.n14 VTAIL.t3 16.3641
R166 VTAIL.n12 VTAIL.t12 16.3641
R167 VTAIL.n12 VTAIL.t11 16.3641
R168 VTAIL.n9 VTAIL.t19 16.3641
R169 VTAIL.n9 VTAIL.t17 16.3641
R170 VTAIL.n7 VTAIL.t1 16.3641
R171 VTAIL.n7 VTAIL.t16 16.3641
R172 VTAIL.n17 VTAIL.n16 15.8669
R173 VTAIL.n10 VTAIL.n8 2.4574
R174 VTAIL.n11 VTAIL.n10 2.4574
R175 VTAIL.n15 VTAIL.n13 2.4574
R176 VTAIL.n16 VTAIL.n15 2.4574
R177 VTAIL.n6 VTAIL.n4 2.4574
R178 VTAIL.n4 VTAIL.n2 2.4574
R179 VTAIL.n19 VTAIL.n17 2.4574
R180 VTAIL VTAIL.n1 1.90136
R181 VTAIL.n13 VTAIL.n11 1.69878
R182 VTAIL.n2 VTAIL.n1 1.69878
R183 VTAIL VTAIL.n19 0.556535
R184 VDD1.n1 VDD1.t2 173.686
R185 VDD1.n3 VDD1.t7 173.686
R186 VDD1.n5 VDD1.n4 146.858
R187 VDD1.n3 VDD1.n2 145.071
R188 VDD1.n7 VDD1.n6 145.071
R189 VDD1.n1 VDD1.n0 145.071
R190 VDD1.n7 VDD1.n5 38.2401
R191 VDD1.n6 VDD1.t8 16.3641
R192 VDD1.n6 VDD1.t9 16.3641
R193 VDD1.n0 VDD1.t3 16.3641
R194 VDD1.n0 VDD1.t4 16.3641
R195 VDD1.n4 VDD1.t6 16.3641
R196 VDD1.n4 VDD1.t1 16.3641
R197 VDD1.n2 VDD1.t5 16.3641
R198 VDD1.n2 VDD1.t0 16.3641
R199 VDD1 VDD1.n7 1.78498
R200 VDD1 VDD1.n1 0.672914
R201 VDD1.n5 VDD1.n3 0.559378
R202 B.n569 B.n568 585
R203 B.n569 B.n107 585
R204 B.n572 B.n571 585
R205 B.n573 B.n126 585
R206 B.n575 B.n574 585
R207 B.n577 B.n125 585
R208 B.n580 B.n579 585
R209 B.n581 B.n124 585
R210 B.n583 B.n582 585
R211 B.n585 B.n123 585
R212 B.n588 B.n587 585
R213 B.n590 B.n120 585
R214 B.n592 B.n591 585
R215 B.n594 B.n119 585
R216 B.n597 B.n596 585
R217 B.n598 B.n118 585
R218 B.n600 B.n599 585
R219 B.n602 B.n117 585
R220 B.n604 B.n603 585
R221 B.n606 B.n605 585
R222 B.n609 B.n608 585
R223 B.n610 B.n112 585
R224 B.n612 B.n611 585
R225 B.n614 B.n111 585
R226 B.n617 B.n616 585
R227 B.n618 B.n110 585
R228 B.n620 B.n619 585
R229 B.n622 B.n109 585
R230 B.n625 B.n624 585
R231 B.n626 B.n108 585
R232 B.n567 B.n106 585
R233 B.n629 B.n106 585
R234 B.n566 B.n105 585
R235 B.n630 B.n105 585
R236 B.n565 B.n104 585
R237 B.n631 B.n104 585
R238 B.n564 B.n563 585
R239 B.n563 B.n100 585
R240 B.n562 B.n99 585
R241 B.n637 B.n99 585
R242 B.n561 B.n98 585
R243 B.n638 B.n98 585
R244 B.n560 B.n97 585
R245 B.n639 B.n97 585
R246 B.n559 B.n558 585
R247 B.n558 B.n96 585
R248 B.n557 B.n92 585
R249 B.n645 B.n92 585
R250 B.n556 B.n91 585
R251 B.n646 B.n91 585
R252 B.n555 B.n90 585
R253 B.n647 B.n90 585
R254 B.n554 B.n553 585
R255 B.n553 B.n86 585
R256 B.n552 B.n85 585
R257 B.n653 B.n85 585
R258 B.n551 B.n84 585
R259 B.n654 B.n84 585
R260 B.n550 B.n83 585
R261 B.n655 B.n83 585
R262 B.n549 B.n548 585
R263 B.n548 B.n79 585
R264 B.n547 B.n78 585
R265 B.n661 B.n78 585
R266 B.n546 B.n77 585
R267 B.n662 B.n77 585
R268 B.n545 B.n76 585
R269 B.n663 B.n76 585
R270 B.n544 B.n543 585
R271 B.n543 B.n75 585
R272 B.n542 B.n71 585
R273 B.n669 B.n71 585
R274 B.n541 B.n70 585
R275 B.n670 B.n70 585
R276 B.n540 B.n69 585
R277 B.n671 B.n69 585
R278 B.n539 B.n538 585
R279 B.n538 B.n65 585
R280 B.n537 B.n64 585
R281 B.n677 B.n64 585
R282 B.n536 B.n63 585
R283 B.n678 B.n63 585
R284 B.n535 B.n62 585
R285 B.n679 B.n62 585
R286 B.n534 B.n533 585
R287 B.n533 B.n61 585
R288 B.n532 B.n57 585
R289 B.n685 B.n57 585
R290 B.n531 B.n56 585
R291 B.n686 B.n56 585
R292 B.n530 B.n55 585
R293 B.n687 B.n55 585
R294 B.n529 B.n528 585
R295 B.n528 B.n51 585
R296 B.n527 B.n50 585
R297 B.n693 B.n50 585
R298 B.n526 B.n49 585
R299 B.n694 B.n49 585
R300 B.n525 B.n48 585
R301 B.n695 B.n48 585
R302 B.n524 B.n523 585
R303 B.n523 B.n47 585
R304 B.n522 B.n43 585
R305 B.n701 B.n43 585
R306 B.n521 B.n42 585
R307 B.n702 B.n42 585
R308 B.n520 B.n41 585
R309 B.n703 B.n41 585
R310 B.n519 B.n518 585
R311 B.n518 B.n37 585
R312 B.n517 B.n36 585
R313 B.n709 B.n36 585
R314 B.n516 B.n35 585
R315 B.n710 B.n35 585
R316 B.n515 B.n34 585
R317 B.n711 B.n34 585
R318 B.n514 B.n513 585
R319 B.n513 B.n30 585
R320 B.n512 B.n29 585
R321 B.n717 B.n29 585
R322 B.n511 B.n28 585
R323 B.n718 B.n28 585
R324 B.n510 B.n27 585
R325 B.n719 B.n27 585
R326 B.n509 B.n508 585
R327 B.n508 B.n23 585
R328 B.n507 B.n22 585
R329 B.n725 B.n22 585
R330 B.n506 B.n21 585
R331 B.n726 B.n21 585
R332 B.n505 B.n20 585
R333 B.n727 B.n20 585
R334 B.n504 B.n503 585
R335 B.n503 B.n16 585
R336 B.n502 B.n15 585
R337 B.n733 B.n15 585
R338 B.n501 B.n14 585
R339 B.n734 B.n14 585
R340 B.n500 B.n13 585
R341 B.n735 B.n13 585
R342 B.n499 B.n498 585
R343 B.n498 B.n12 585
R344 B.n497 B.n496 585
R345 B.n497 B.n8 585
R346 B.n495 B.n7 585
R347 B.n742 B.n7 585
R348 B.n494 B.n6 585
R349 B.n743 B.n6 585
R350 B.n493 B.n5 585
R351 B.n744 B.n5 585
R352 B.n492 B.n491 585
R353 B.n491 B.n4 585
R354 B.n490 B.n127 585
R355 B.n490 B.n489 585
R356 B.n480 B.n128 585
R357 B.n129 B.n128 585
R358 B.n482 B.n481 585
R359 B.n483 B.n482 585
R360 B.n479 B.n134 585
R361 B.n134 B.n133 585
R362 B.n478 B.n477 585
R363 B.n477 B.n476 585
R364 B.n136 B.n135 585
R365 B.n137 B.n136 585
R366 B.n469 B.n468 585
R367 B.n470 B.n469 585
R368 B.n467 B.n142 585
R369 B.n142 B.n141 585
R370 B.n466 B.n465 585
R371 B.n465 B.n464 585
R372 B.n144 B.n143 585
R373 B.n145 B.n144 585
R374 B.n457 B.n456 585
R375 B.n458 B.n457 585
R376 B.n455 B.n150 585
R377 B.n150 B.n149 585
R378 B.n454 B.n453 585
R379 B.n453 B.n452 585
R380 B.n152 B.n151 585
R381 B.n153 B.n152 585
R382 B.n445 B.n444 585
R383 B.n446 B.n445 585
R384 B.n443 B.n158 585
R385 B.n158 B.n157 585
R386 B.n442 B.n441 585
R387 B.n441 B.n440 585
R388 B.n160 B.n159 585
R389 B.n161 B.n160 585
R390 B.n433 B.n432 585
R391 B.n434 B.n433 585
R392 B.n431 B.n166 585
R393 B.n166 B.n165 585
R394 B.n430 B.n429 585
R395 B.n429 B.n428 585
R396 B.n168 B.n167 585
R397 B.n421 B.n168 585
R398 B.n420 B.n419 585
R399 B.n422 B.n420 585
R400 B.n418 B.n173 585
R401 B.n173 B.n172 585
R402 B.n417 B.n416 585
R403 B.n416 B.n415 585
R404 B.n175 B.n174 585
R405 B.n176 B.n175 585
R406 B.n408 B.n407 585
R407 B.n409 B.n408 585
R408 B.n406 B.n181 585
R409 B.n181 B.n180 585
R410 B.n405 B.n404 585
R411 B.n404 B.n403 585
R412 B.n183 B.n182 585
R413 B.n396 B.n183 585
R414 B.n395 B.n394 585
R415 B.n397 B.n395 585
R416 B.n393 B.n188 585
R417 B.n188 B.n187 585
R418 B.n392 B.n391 585
R419 B.n391 B.n390 585
R420 B.n190 B.n189 585
R421 B.n191 B.n190 585
R422 B.n383 B.n382 585
R423 B.n384 B.n383 585
R424 B.n381 B.n196 585
R425 B.n196 B.n195 585
R426 B.n380 B.n379 585
R427 B.n379 B.n378 585
R428 B.n198 B.n197 585
R429 B.n371 B.n198 585
R430 B.n370 B.n369 585
R431 B.n372 B.n370 585
R432 B.n368 B.n203 585
R433 B.n203 B.n202 585
R434 B.n367 B.n366 585
R435 B.n366 B.n365 585
R436 B.n205 B.n204 585
R437 B.n206 B.n205 585
R438 B.n358 B.n357 585
R439 B.n359 B.n358 585
R440 B.n356 B.n211 585
R441 B.n211 B.n210 585
R442 B.n355 B.n354 585
R443 B.n354 B.n353 585
R444 B.n213 B.n212 585
R445 B.n214 B.n213 585
R446 B.n346 B.n345 585
R447 B.n347 B.n346 585
R448 B.n344 B.n219 585
R449 B.n219 B.n218 585
R450 B.n343 B.n342 585
R451 B.n342 B.n341 585
R452 B.n221 B.n220 585
R453 B.n334 B.n221 585
R454 B.n333 B.n332 585
R455 B.n335 B.n333 585
R456 B.n331 B.n226 585
R457 B.n226 B.n225 585
R458 B.n330 B.n329 585
R459 B.n329 B.n328 585
R460 B.n228 B.n227 585
R461 B.n229 B.n228 585
R462 B.n321 B.n320 585
R463 B.n322 B.n321 585
R464 B.n319 B.n234 585
R465 B.n234 B.n233 585
R466 B.n318 B.n317 585
R467 B.n317 B.n316 585
R468 B.n313 B.n238 585
R469 B.n312 B.n311 585
R470 B.n309 B.n239 585
R471 B.n309 B.n237 585
R472 B.n308 B.n307 585
R473 B.n306 B.n305 585
R474 B.n304 B.n241 585
R475 B.n302 B.n301 585
R476 B.n300 B.n242 585
R477 B.n299 B.n298 585
R478 B.n296 B.n243 585
R479 B.n294 B.n293 585
R480 B.n292 B.n244 585
R481 B.n291 B.n290 585
R482 B.n288 B.n248 585
R483 B.n286 B.n285 585
R484 B.n284 B.n249 585
R485 B.n283 B.n282 585
R486 B.n280 B.n250 585
R487 B.n278 B.n277 585
R488 B.n275 B.n251 585
R489 B.n274 B.n273 585
R490 B.n271 B.n254 585
R491 B.n269 B.n268 585
R492 B.n267 B.n255 585
R493 B.n266 B.n265 585
R494 B.n263 B.n256 585
R495 B.n261 B.n260 585
R496 B.n259 B.n258 585
R497 B.n236 B.n235 585
R498 B.n315 B.n314 585
R499 B.n316 B.n315 585
R500 B.n232 B.n231 585
R501 B.n233 B.n232 585
R502 B.n324 B.n323 585
R503 B.n323 B.n322 585
R504 B.n325 B.n230 585
R505 B.n230 B.n229 585
R506 B.n327 B.n326 585
R507 B.n328 B.n327 585
R508 B.n224 B.n223 585
R509 B.n225 B.n224 585
R510 B.n337 B.n336 585
R511 B.n336 B.n335 585
R512 B.n338 B.n222 585
R513 B.n334 B.n222 585
R514 B.n340 B.n339 585
R515 B.n341 B.n340 585
R516 B.n217 B.n216 585
R517 B.n218 B.n217 585
R518 B.n349 B.n348 585
R519 B.n348 B.n347 585
R520 B.n350 B.n215 585
R521 B.n215 B.n214 585
R522 B.n352 B.n351 585
R523 B.n353 B.n352 585
R524 B.n209 B.n208 585
R525 B.n210 B.n209 585
R526 B.n361 B.n360 585
R527 B.n360 B.n359 585
R528 B.n362 B.n207 585
R529 B.n207 B.n206 585
R530 B.n364 B.n363 585
R531 B.n365 B.n364 585
R532 B.n201 B.n200 585
R533 B.n202 B.n201 585
R534 B.n374 B.n373 585
R535 B.n373 B.n372 585
R536 B.n375 B.n199 585
R537 B.n371 B.n199 585
R538 B.n377 B.n376 585
R539 B.n378 B.n377 585
R540 B.n194 B.n193 585
R541 B.n195 B.n194 585
R542 B.n386 B.n385 585
R543 B.n385 B.n384 585
R544 B.n387 B.n192 585
R545 B.n192 B.n191 585
R546 B.n389 B.n388 585
R547 B.n390 B.n389 585
R548 B.n186 B.n185 585
R549 B.n187 B.n186 585
R550 B.n399 B.n398 585
R551 B.n398 B.n397 585
R552 B.n400 B.n184 585
R553 B.n396 B.n184 585
R554 B.n402 B.n401 585
R555 B.n403 B.n402 585
R556 B.n179 B.n178 585
R557 B.n180 B.n179 585
R558 B.n411 B.n410 585
R559 B.n410 B.n409 585
R560 B.n412 B.n177 585
R561 B.n177 B.n176 585
R562 B.n414 B.n413 585
R563 B.n415 B.n414 585
R564 B.n171 B.n170 585
R565 B.n172 B.n171 585
R566 B.n424 B.n423 585
R567 B.n423 B.n422 585
R568 B.n425 B.n169 585
R569 B.n421 B.n169 585
R570 B.n427 B.n426 585
R571 B.n428 B.n427 585
R572 B.n164 B.n163 585
R573 B.n165 B.n164 585
R574 B.n436 B.n435 585
R575 B.n435 B.n434 585
R576 B.n437 B.n162 585
R577 B.n162 B.n161 585
R578 B.n439 B.n438 585
R579 B.n440 B.n439 585
R580 B.n156 B.n155 585
R581 B.n157 B.n156 585
R582 B.n448 B.n447 585
R583 B.n447 B.n446 585
R584 B.n449 B.n154 585
R585 B.n154 B.n153 585
R586 B.n451 B.n450 585
R587 B.n452 B.n451 585
R588 B.n148 B.n147 585
R589 B.n149 B.n148 585
R590 B.n460 B.n459 585
R591 B.n459 B.n458 585
R592 B.n461 B.n146 585
R593 B.n146 B.n145 585
R594 B.n463 B.n462 585
R595 B.n464 B.n463 585
R596 B.n140 B.n139 585
R597 B.n141 B.n140 585
R598 B.n472 B.n471 585
R599 B.n471 B.n470 585
R600 B.n473 B.n138 585
R601 B.n138 B.n137 585
R602 B.n475 B.n474 585
R603 B.n476 B.n475 585
R604 B.n132 B.n131 585
R605 B.n133 B.n132 585
R606 B.n485 B.n484 585
R607 B.n484 B.n483 585
R608 B.n486 B.n130 585
R609 B.n130 B.n129 585
R610 B.n488 B.n487 585
R611 B.n489 B.n488 585
R612 B.n3 B.n0 585
R613 B.n4 B.n3 585
R614 B.n741 B.n1 585
R615 B.n742 B.n741 585
R616 B.n740 B.n739 585
R617 B.n740 B.n8 585
R618 B.n738 B.n9 585
R619 B.n12 B.n9 585
R620 B.n737 B.n736 585
R621 B.n736 B.n735 585
R622 B.n11 B.n10 585
R623 B.n734 B.n11 585
R624 B.n732 B.n731 585
R625 B.n733 B.n732 585
R626 B.n730 B.n17 585
R627 B.n17 B.n16 585
R628 B.n729 B.n728 585
R629 B.n728 B.n727 585
R630 B.n19 B.n18 585
R631 B.n726 B.n19 585
R632 B.n724 B.n723 585
R633 B.n725 B.n724 585
R634 B.n722 B.n24 585
R635 B.n24 B.n23 585
R636 B.n721 B.n720 585
R637 B.n720 B.n719 585
R638 B.n26 B.n25 585
R639 B.n718 B.n26 585
R640 B.n716 B.n715 585
R641 B.n717 B.n716 585
R642 B.n714 B.n31 585
R643 B.n31 B.n30 585
R644 B.n713 B.n712 585
R645 B.n712 B.n711 585
R646 B.n33 B.n32 585
R647 B.n710 B.n33 585
R648 B.n708 B.n707 585
R649 B.n709 B.n708 585
R650 B.n706 B.n38 585
R651 B.n38 B.n37 585
R652 B.n705 B.n704 585
R653 B.n704 B.n703 585
R654 B.n40 B.n39 585
R655 B.n702 B.n40 585
R656 B.n700 B.n699 585
R657 B.n701 B.n700 585
R658 B.n698 B.n44 585
R659 B.n47 B.n44 585
R660 B.n697 B.n696 585
R661 B.n696 B.n695 585
R662 B.n46 B.n45 585
R663 B.n694 B.n46 585
R664 B.n692 B.n691 585
R665 B.n693 B.n692 585
R666 B.n690 B.n52 585
R667 B.n52 B.n51 585
R668 B.n689 B.n688 585
R669 B.n688 B.n687 585
R670 B.n54 B.n53 585
R671 B.n686 B.n54 585
R672 B.n684 B.n683 585
R673 B.n685 B.n684 585
R674 B.n682 B.n58 585
R675 B.n61 B.n58 585
R676 B.n681 B.n680 585
R677 B.n680 B.n679 585
R678 B.n60 B.n59 585
R679 B.n678 B.n60 585
R680 B.n676 B.n675 585
R681 B.n677 B.n676 585
R682 B.n674 B.n66 585
R683 B.n66 B.n65 585
R684 B.n673 B.n672 585
R685 B.n672 B.n671 585
R686 B.n68 B.n67 585
R687 B.n670 B.n68 585
R688 B.n668 B.n667 585
R689 B.n669 B.n668 585
R690 B.n666 B.n72 585
R691 B.n75 B.n72 585
R692 B.n665 B.n664 585
R693 B.n664 B.n663 585
R694 B.n74 B.n73 585
R695 B.n662 B.n74 585
R696 B.n660 B.n659 585
R697 B.n661 B.n660 585
R698 B.n658 B.n80 585
R699 B.n80 B.n79 585
R700 B.n657 B.n656 585
R701 B.n656 B.n655 585
R702 B.n82 B.n81 585
R703 B.n654 B.n82 585
R704 B.n652 B.n651 585
R705 B.n653 B.n652 585
R706 B.n650 B.n87 585
R707 B.n87 B.n86 585
R708 B.n649 B.n648 585
R709 B.n648 B.n647 585
R710 B.n89 B.n88 585
R711 B.n646 B.n89 585
R712 B.n644 B.n643 585
R713 B.n645 B.n644 585
R714 B.n642 B.n93 585
R715 B.n96 B.n93 585
R716 B.n641 B.n640 585
R717 B.n640 B.n639 585
R718 B.n95 B.n94 585
R719 B.n638 B.n95 585
R720 B.n636 B.n635 585
R721 B.n637 B.n636 585
R722 B.n634 B.n101 585
R723 B.n101 B.n100 585
R724 B.n633 B.n632 585
R725 B.n632 B.n631 585
R726 B.n103 B.n102 585
R727 B.n630 B.n103 585
R728 B.n628 B.n627 585
R729 B.n629 B.n628 585
R730 B.n745 B.n744 585
R731 B.n743 B.n2 585
R732 B.n628 B.n108 511.721
R733 B.n569 B.n106 511.721
R734 B.n317 B.n236 511.721
R735 B.n315 B.n238 511.721
R736 B.n570 B.n107 256.663
R737 B.n576 B.n107 256.663
R738 B.n578 B.n107 256.663
R739 B.n584 B.n107 256.663
R740 B.n586 B.n107 256.663
R741 B.n593 B.n107 256.663
R742 B.n595 B.n107 256.663
R743 B.n601 B.n107 256.663
R744 B.n116 B.n107 256.663
R745 B.n607 B.n107 256.663
R746 B.n613 B.n107 256.663
R747 B.n615 B.n107 256.663
R748 B.n621 B.n107 256.663
R749 B.n623 B.n107 256.663
R750 B.n310 B.n237 256.663
R751 B.n240 B.n237 256.663
R752 B.n303 B.n237 256.663
R753 B.n297 B.n237 256.663
R754 B.n295 B.n237 256.663
R755 B.n289 B.n237 256.663
R756 B.n287 B.n237 256.663
R757 B.n281 B.n237 256.663
R758 B.n279 B.n237 256.663
R759 B.n272 B.n237 256.663
R760 B.n270 B.n237 256.663
R761 B.n264 B.n237 256.663
R762 B.n262 B.n237 256.663
R763 B.n257 B.n237 256.663
R764 B.n747 B.n746 256.663
R765 B.n113 B.t18 208.704
R766 B.n121 B.t14 208.704
R767 B.n252 B.t21 208.704
R768 B.n245 B.t10 208.704
R769 B.n113 B.t19 203.706
R770 B.n245 B.t13 203.706
R771 B.n121 B.t16 203.706
R772 B.n252 B.t23 203.706
R773 B.n316 B.n237 198.458
R774 B.n629 B.n107 198.458
R775 B.n624 B.n622 163.367
R776 B.n620 B.n110 163.367
R777 B.n616 B.n614 163.367
R778 B.n612 B.n112 163.367
R779 B.n608 B.n606 163.367
R780 B.n603 B.n602 163.367
R781 B.n600 B.n118 163.367
R782 B.n596 B.n594 163.367
R783 B.n592 B.n120 163.367
R784 B.n587 B.n585 163.367
R785 B.n583 B.n124 163.367
R786 B.n579 B.n577 163.367
R787 B.n575 B.n126 163.367
R788 B.n571 B.n569 163.367
R789 B.n317 B.n234 163.367
R790 B.n321 B.n234 163.367
R791 B.n321 B.n228 163.367
R792 B.n329 B.n228 163.367
R793 B.n329 B.n226 163.367
R794 B.n333 B.n226 163.367
R795 B.n333 B.n221 163.367
R796 B.n342 B.n221 163.367
R797 B.n342 B.n219 163.367
R798 B.n346 B.n219 163.367
R799 B.n346 B.n213 163.367
R800 B.n354 B.n213 163.367
R801 B.n354 B.n211 163.367
R802 B.n358 B.n211 163.367
R803 B.n358 B.n205 163.367
R804 B.n366 B.n205 163.367
R805 B.n366 B.n203 163.367
R806 B.n370 B.n203 163.367
R807 B.n370 B.n198 163.367
R808 B.n379 B.n198 163.367
R809 B.n379 B.n196 163.367
R810 B.n383 B.n196 163.367
R811 B.n383 B.n190 163.367
R812 B.n391 B.n190 163.367
R813 B.n391 B.n188 163.367
R814 B.n395 B.n188 163.367
R815 B.n395 B.n183 163.367
R816 B.n404 B.n183 163.367
R817 B.n404 B.n181 163.367
R818 B.n408 B.n181 163.367
R819 B.n408 B.n175 163.367
R820 B.n416 B.n175 163.367
R821 B.n416 B.n173 163.367
R822 B.n420 B.n173 163.367
R823 B.n420 B.n168 163.367
R824 B.n429 B.n168 163.367
R825 B.n429 B.n166 163.367
R826 B.n433 B.n166 163.367
R827 B.n433 B.n160 163.367
R828 B.n441 B.n160 163.367
R829 B.n441 B.n158 163.367
R830 B.n445 B.n158 163.367
R831 B.n445 B.n152 163.367
R832 B.n453 B.n152 163.367
R833 B.n453 B.n150 163.367
R834 B.n457 B.n150 163.367
R835 B.n457 B.n144 163.367
R836 B.n465 B.n144 163.367
R837 B.n465 B.n142 163.367
R838 B.n469 B.n142 163.367
R839 B.n469 B.n136 163.367
R840 B.n477 B.n136 163.367
R841 B.n477 B.n134 163.367
R842 B.n482 B.n134 163.367
R843 B.n482 B.n128 163.367
R844 B.n490 B.n128 163.367
R845 B.n491 B.n490 163.367
R846 B.n491 B.n5 163.367
R847 B.n6 B.n5 163.367
R848 B.n7 B.n6 163.367
R849 B.n497 B.n7 163.367
R850 B.n498 B.n497 163.367
R851 B.n498 B.n13 163.367
R852 B.n14 B.n13 163.367
R853 B.n15 B.n14 163.367
R854 B.n503 B.n15 163.367
R855 B.n503 B.n20 163.367
R856 B.n21 B.n20 163.367
R857 B.n22 B.n21 163.367
R858 B.n508 B.n22 163.367
R859 B.n508 B.n27 163.367
R860 B.n28 B.n27 163.367
R861 B.n29 B.n28 163.367
R862 B.n513 B.n29 163.367
R863 B.n513 B.n34 163.367
R864 B.n35 B.n34 163.367
R865 B.n36 B.n35 163.367
R866 B.n518 B.n36 163.367
R867 B.n518 B.n41 163.367
R868 B.n42 B.n41 163.367
R869 B.n43 B.n42 163.367
R870 B.n523 B.n43 163.367
R871 B.n523 B.n48 163.367
R872 B.n49 B.n48 163.367
R873 B.n50 B.n49 163.367
R874 B.n528 B.n50 163.367
R875 B.n528 B.n55 163.367
R876 B.n56 B.n55 163.367
R877 B.n57 B.n56 163.367
R878 B.n533 B.n57 163.367
R879 B.n533 B.n62 163.367
R880 B.n63 B.n62 163.367
R881 B.n64 B.n63 163.367
R882 B.n538 B.n64 163.367
R883 B.n538 B.n69 163.367
R884 B.n70 B.n69 163.367
R885 B.n71 B.n70 163.367
R886 B.n543 B.n71 163.367
R887 B.n543 B.n76 163.367
R888 B.n77 B.n76 163.367
R889 B.n78 B.n77 163.367
R890 B.n548 B.n78 163.367
R891 B.n548 B.n83 163.367
R892 B.n84 B.n83 163.367
R893 B.n85 B.n84 163.367
R894 B.n553 B.n85 163.367
R895 B.n553 B.n90 163.367
R896 B.n91 B.n90 163.367
R897 B.n92 B.n91 163.367
R898 B.n558 B.n92 163.367
R899 B.n558 B.n97 163.367
R900 B.n98 B.n97 163.367
R901 B.n99 B.n98 163.367
R902 B.n563 B.n99 163.367
R903 B.n563 B.n104 163.367
R904 B.n105 B.n104 163.367
R905 B.n106 B.n105 163.367
R906 B.n311 B.n309 163.367
R907 B.n309 B.n308 163.367
R908 B.n305 B.n304 163.367
R909 B.n302 B.n242 163.367
R910 B.n298 B.n296 163.367
R911 B.n294 B.n244 163.367
R912 B.n290 B.n288 163.367
R913 B.n286 B.n249 163.367
R914 B.n282 B.n280 163.367
R915 B.n278 B.n251 163.367
R916 B.n273 B.n271 163.367
R917 B.n269 B.n255 163.367
R918 B.n265 B.n263 163.367
R919 B.n261 B.n258 163.367
R920 B.n315 B.n232 163.367
R921 B.n323 B.n232 163.367
R922 B.n323 B.n230 163.367
R923 B.n327 B.n230 163.367
R924 B.n327 B.n224 163.367
R925 B.n336 B.n224 163.367
R926 B.n336 B.n222 163.367
R927 B.n340 B.n222 163.367
R928 B.n340 B.n217 163.367
R929 B.n348 B.n217 163.367
R930 B.n348 B.n215 163.367
R931 B.n352 B.n215 163.367
R932 B.n352 B.n209 163.367
R933 B.n360 B.n209 163.367
R934 B.n360 B.n207 163.367
R935 B.n364 B.n207 163.367
R936 B.n364 B.n201 163.367
R937 B.n373 B.n201 163.367
R938 B.n373 B.n199 163.367
R939 B.n377 B.n199 163.367
R940 B.n377 B.n194 163.367
R941 B.n385 B.n194 163.367
R942 B.n385 B.n192 163.367
R943 B.n389 B.n192 163.367
R944 B.n389 B.n186 163.367
R945 B.n398 B.n186 163.367
R946 B.n398 B.n184 163.367
R947 B.n402 B.n184 163.367
R948 B.n402 B.n179 163.367
R949 B.n410 B.n179 163.367
R950 B.n410 B.n177 163.367
R951 B.n414 B.n177 163.367
R952 B.n414 B.n171 163.367
R953 B.n423 B.n171 163.367
R954 B.n423 B.n169 163.367
R955 B.n427 B.n169 163.367
R956 B.n427 B.n164 163.367
R957 B.n435 B.n164 163.367
R958 B.n435 B.n162 163.367
R959 B.n439 B.n162 163.367
R960 B.n439 B.n156 163.367
R961 B.n447 B.n156 163.367
R962 B.n447 B.n154 163.367
R963 B.n451 B.n154 163.367
R964 B.n451 B.n148 163.367
R965 B.n459 B.n148 163.367
R966 B.n459 B.n146 163.367
R967 B.n463 B.n146 163.367
R968 B.n463 B.n140 163.367
R969 B.n471 B.n140 163.367
R970 B.n471 B.n138 163.367
R971 B.n475 B.n138 163.367
R972 B.n475 B.n132 163.367
R973 B.n484 B.n132 163.367
R974 B.n484 B.n130 163.367
R975 B.n488 B.n130 163.367
R976 B.n488 B.n3 163.367
R977 B.n745 B.n3 163.367
R978 B.n741 B.n2 163.367
R979 B.n741 B.n740 163.367
R980 B.n740 B.n9 163.367
R981 B.n736 B.n9 163.367
R982 B.n736 B.n11 163.367
R983 B.n732 B.n11 163.367
R984 B.n732 B.n17 163.367
R985 B.n728 B.n17 163.367
R986 B.n728 B.n19 163.367
R987 B.n724 B.n19 163.367
R988 B.n724 B.n24 163.367
R989 B.n720 B.n24 163.367
R990 B.n720 B.n26 163.367
R991 B.n716 B.n26 163.367
R992 B.n716 B.n31 163.367
R993 B.n712 B.n31 163.367
R994 B.n712 B.n33 163.367
R995 B.n708 B.n33 163.367
R996 B.n708 B.n38 163.367
R997 B.n704 B.n38 163.367
R998 B.n704 B.n40 163.367
R999 B.n700 B.n40 163.367
R1000 B.n700 B.n44 163.367
R1001 B.n696 B.n44 163.367
R1002 B.n696 B.n46 163.367
R1003 B.n692 B.n46 163.367
R1004 B.n692 B.n52 163.367
R1005 B.n688 B.n52 163.367
R1006 B.n688 B.n54 163.367
R1007 B.n684 B.n54 163.367
R1008 B.n684 B.n58 163.367
R1009 B.n680 B.n58 163.367
R1010 B.n680 B.n60 163.367
R1011 B.n676 B.n60 163.367
R1012 B.n676 B.n66 163.367
R1013 B.n672 B.n66 163.367
R1014 B.n672 B.n68 163.367
R1015 B.n668 B.n68 163.367
R1016 B.n668 B.n72 163.367
R1017 B.n664 B.n72 163.367
R1018 B.n664 B.n74 163.367
R1019 B.n660 B.n74 163.367
R1020 B.n660 B.n80 163.367
R1021 B.n656 B.n80 163.367
R1022 B.n656 B.n82 163.367
R1023 B.n652 B.n82 163.367
R1024 B.n652 B.n87 163.367
R1025 B.n648 B.n87 163.367
R1026 B.n648 B.n89 163.367
R1027 B.n644 B.n89 163.367
R1028 B.n644 B.n93 163.367
R1029 B.n640 B.n93 163.367
R1030 B.n640 B.n95 163.367
R1031 B.n636 B.n95 163.367
R1032 B.n636 B.n101 163.367
R1033 B.n632 B.n101 163.367
R1034 B.n632 B.n103 163.367
R1035 B.n628 B.n103 163.367
R1036 B.n114 B.t20 148.433
R1037 B.n122 B.t17 148.433
R1038 B.n253 B.t22 148.433
R1039 B.n246 B.t12 148.433
R1040 B.n316 B.n233 115.344
R1041 B.n322 B.n233 115.344
R1042 B.n322 B.n229 115.344
R1043 B.n328 B.n229 115.344
R1044 B.n328 B.n225 115.344
R1045 B.n335 B.n225 115.344
R1046 B.n335 B.n334 115.344
R1047 B.n341 B.n218 115.344
R1048 B.n347 B.n218 115.344
R1049 B.n347 B.n214 115.344
R1050 B.n353 B.n214 115.344
R1051 B.n353 B.n210 115.344
R1052 B.n359 B.n210 115.344
R1053 B.n359 B.n206 115.344
R1054 B.n365 B.n206 115.344
R1055 B.n365 B.n202 115.344
R1056 B.n372 B.n202 115.344
R1057 B.n372 B.n371 115.344
R1058 B.n378 B.n195 115.344
R1059 B.n384 B.n195 115.344
R1060 B.n384 B.n191 115.344
R1061 B.n390 B.n191 115.344
R1062 B.n390 B.n187 115.344
R1063 B.n397 B.n187 115.344
R1064 B.n397 B.n396 115.344
R1065 B.n403 B.n180 115.344
R1066 B.n409 B.n180 115.344
R1067 B.n409 B.n176 115.344
R1068 B.n415 B.n176 115.344
R1069 B.n415 B.n172 115.344
R1070 B.n422 B.n172 115.344
R1071 B.n422 B.n421 115.344
R1072 B.n428 B.n165 115.344
R1073 B.n434 B.n165 115.344
R1074 B.n434 B.n161 115.344
R1075 B.n440 B.n161 115.344
R1076 B.n440 B.n157 115.344
R1077 B.n446 B.n157 115.344
R1078 B.n446 B.n153 115.344
R1079 B.n452 B.n153 115.344
R1080 B.n458 B.n149 115.344
R1081 B.n458 B.n145 115.344
R1082 B.n464 B.n145 115.344
R1083 B.n464 B.n141 115.344
R1084 B.n470 B.n141 115.344
R1085 B.n470 B.n137 115.344
R1086 B.n476 B.n137 115.344
R1087 B.n483 B.n133 115.344
R1088 B.n483 B.n129 115.344
R1089 B.n489 B.n129 115.344
R1090 B.n489 B.n4 115.344
R1091 B.n744 B.n4 115.344
R1092 B.n744 B.n743 115.344
R1093 B.n743 B.n742 115.344
R1094 B.n742 B.n8 115.344
R1095 B.n12 B.n8 115.344
R1096 B.n735 B.n12 115.344
R1097 B.n735 B.n734 115.344
R1098 B.n733 B.n16 115.344
R1099 B.n727 B.n16 115.344
R1100 B.n727 B.n726 115.344
R1101 B.n726 B.n725 115.344
R1102 B.n725 B.n23 115.344
R1103 B.n719 B.n23 115.344
R1104 B.n719 B.n718 115.344
R1105 B.n717 B.n30 115.344
R1106 B.n711 B.n30 115.344
R1107 B.n711 B.n710 115.344
R1108 B.n710 B.n709 115.344
R1109 B.n709 B.n37 115.344
R1110 B.n703 B.n37 115.344
R1111 B.n703 B.n702 115.344
R1112 B.n702 B.n701 115.344
R1113 B.n695 B.n47 115.344
R1114 B.n695 B.n694 115.344
R1115 B.n694 B.n693 115.344
R1116 B.n693 B.n51 115.344
R1117 B.n687 B.n51 115.344
R1118 B.n687 B.n686 115.344
R1119 B.n686 B.n685 115.344
R1120 B.n679 B.n61 115.344
R1121 B.n679 B.n678 115.344
R1122 B.n678 B.n677 115.344
R1123 B.n677 B.n65 115.344
R1124 B.n671 B.n65 115.344
R1125 B.n671 B.n670 115.344
R1126 B.n670 B.n669 115.344
R1127 B.n663 B.n75 115.344
R1128 B.n663 B.n662 115.344
R1129 B.n662 B.n661 115.344
R1130 B.n661 B.n79 115.344
R1131 B.n655 B.n79 115.344
R1132 B.n655 B.n654 115.344
R1133 B.n654 B.n653 115.344
R1134 B.n653 B.n86 115.344
R1135 B.n647 B.n86 115.344
R1136 B.n647 B.n646 115.344
R1137 B.n646 B.n645 115.344
R1138 B.n639 B.n96 115.344
R1139 B.n639 B.n638 115.344
R1140 B.n638 B.n637 115.344
R1141 B.n637 B.n100 115.344
R1142 B.n631 B.n100 115.344
R1143 B.n631 B.n630 115.344
R1144 B.n630 B.n629 115.344
R1145 B.n421 B.t3 108.558
R1146 B.n47 B.t6 108.558
R1147 B.n378 B.t1 94.9889
R1148 B.n669 B.t2 94.9889
R1149 B.n476 B.t4 81.4192
R1150 B.t5 B.n733 81.4192
R1151 B.t8 B.n149 78.0267
R1152 B.n718 B.t0 78.0267
R1153 B.n623 B.n108 71.676
R1154 B.n622 B.n621 71.676
R1155 B.n615 B.n110 71.676
R1156 B.n614 B.n613 71.676
R1157 B.n607 B.n112 71.676
R1158 B.n606 B.n116 71.676
R1159 B.n602 B.n601 71.676
R1160 B.n595 B.n118 71.676
R1161 B.n594 B.n593 71.676
R1162 B.n586 B.n120 71.676
R1163 B.n585 B.n584 71.676
R1164 B.n578 B.n124 71.676
R1165 B.n577 B.n576 71.676
R1166 B.n570 B.n126 71.676
R1167 B.n571 B.n570 71.676
R1168 B.n576 B.n575 71.676
R1169 B.n579 B.n578 71.676
R1170 B.n584 B.n583 71.676
R1171 B.n587 B.n586 71.676
R1172 B.n593 B.n592 71.676
R1173 B.n596 B.n595 71.676
R1174 B.n601 B.n600 71.676
R1175 B.n603 B.n116 71.676
R1176 B.n608 B.n607 71.676
R1177 B.n613 B.n612 71.676
R1178 B.n616 B.n615 71.676
R1179 B.n621 B.n620 71.676
R1180 B.n624 B.n623 71.676
R1181 B.n310 B.n238 71.676
R1182 B.n308 B.n240 71.676
R1183 B.n304 B.n303 71.676
R1184 B.n297 B.n242 71.676
R1185 B.n296 B.n295 71.676
R1186 B.n289 B.n244 71.676
R1187 B.n288 B.n287 71.676
R1188 B.n281 B.n249 71.676
R1189 B.n280 B.n279 71.676
R1190 B.n272 B.n251 71.676
R1191 B.n271 B.n270 71.676
R1192 B.n264 B.n255 71.676
R1193 B.n263 B.n262 71.676
R1194 B.n258 B.n257 71.676
R1195 B.n311 B.n310 71.676
R1196 B.n305 B.n240 71.676
R1197 B.n303 B.n302 71.676
R1198 B.n298 B.n297 71.676
R1199 B.n295 B.n294 71.676
R1200 B.n290 B.n289 71.676
R1201 B.n287 B.n286 71.676
R1202 B.n282 B.n281 71.676
R1203 B.n279 B.n278 71.676
R1204 B.n273 B.n272 71.676
R1205 B.n270 B.n269 71.676
R1206 B.n265 B.n264 71.676
R1207 B.n262 B.n261 71.676
R1208 B.n257 B.n236 71.676
R1209 B.n746 B.n745 71.676
R1210 B.n746 B.n2 71.676
R1211 B.n334 B.t11 67.8494
R1212 B.n96 B.t15 67.8494
R1213 B.n396 B.t7 64.4569
R1214 B.n61 B.t9 64.4569
R1215 B.n115 B.n114 59.5399
R1216 B.n589 B.n122 59.5399
R1217 B.n276 B.n253 59.5399
R1218 B.n247 B.n246 59.5399
R1219 B.n114 B.n113 55.2732
R1220 B.n122 B.n121 55.2732
R1221 B.n253 B.n252 55.2732
R1222 B.n246 B.n245 55.2732
R1223 B.n403 B.t7 50.8872
R1224 B.n685 B.t9 50.8872
R1225 B.n341 B.t11 47.4947
R1226 B.n645 B.t15 47.4947
R1227 B.n452 B.t8 37.3174
R1228 B.t0 B.n717 37.3174
R1229 B.t4 B.n133 33.9249
R1230 B.n734 B.t5 33.9249
R1231 B.n314 B.n313 33.2493
R1232 B.n318 B.n235 33.2493
R1233 B.n568 B.n567 33.2493
R1234 B.n627 B.n626 33.2493
R1235 B.n371 B.t1 20.3552
R1236 B.n75 B.t2 20.3552
R1237 B B.n747 18.0485
R1238 B.n314 B.n231 10.6151
R1239 B.n324 B.n231 10.6151
R1240 B.n325 B.n324 10.6151
R1241 B.n326 B.n325 10.6151
R1242 B.n326 B.n223 10.6151
R1243 B.n337 B.n223 10.6151
R1244 B.n338 B.n337 10.6151
R1245 B.n339 B.n338 10.6151
R1246 B.n339 B.n216 10.6151
R1247 B.n349 B.n216 10.6151
R1248 B.n350 B.n349 10.6151
R1249 B.n351 B.n350 10.6151
R1250 B.n351 B.n208 10.6151
R1251 B.n361 B.n208 10.6151
R1252 B.n362 B.n361 10.6151
R1253 B.n363 B.n362 10.6151
R1254 B.n363 B.n200 10.6151
R1255 B.n374 B.n200 10.6151
R1256 B.n375 B.n374 10.6151
R1257 B.n376 B.n375 10.6151
R1258 B.n376 B.n193 10.6151
R1259 B.n386 B.n193 10.6151
R1260 B.n387 B.n386 10.6151
R1261 B.n388 B.n387 10.6151
R1262 B.n388 B.n185 10.6151
R1263 B.n399 B.n185 10.6151
R1264 B.n400 B.n399 10.6151
R1265 B.n401 B.n400 10.6151
R1266 B.n401 B.n178 10.6151
R1267 B.n411 B.n178 10.6151
R1268 B.n412 B.n411 10.6151
R1269 B.n413 B.n412 10.6151
R1270 B.n413 B.n170 10.6151
R1271 B.n424 B.n170 10.6151
R1272 B.n425 B.n424 10.6151
R1273 B.n426 B.n425 10.6151
R1274 B.n426 B.n163 10.6151
R1275 B.n436 B.n163 10.6151
R1276 B.n437 B.n436 10.6151
R1277 B.n438 B.n437 10.6151
R1278 B.n438 B.n155 10.6151
R1279 B.n448 B.n155 10.6151
R1280 B.n449 B.n448 10.6151
R1281 B.n450 B.n449 10.6151
R1282 B.n450 B.n147 10.6151
R1283 B.n460 B.n147 10.6151
R1284 B.n461 B.n460 10.6151
R1285 B.n462 B.n461 10.6151
R1286 B.n462 B.n139 10.6151
R1287 B.n472 B.n139 10.6151
R1288 B.n473 B.n472 10.6151
R1289 B.n474 B.n473 10.6151
R1290 B.n474 B.n131 10.6151
R1291 B.n485 B.n131 10.6151
R1292 B.n486 B.n485 10.6151
R1293 B.n487 B.n486 10.6151
R1294 B.n487 B.n0 10.6151
R1295 B.n313 B.n312 10.6151
R1296 B.n312 B.n239 10.6151
R1297 B.n307 B.n239 10.6151
R1298 B.n307 B.n306 10.6151
R1299 B.n306 B.n241 10.6151
R1300 B.n301 B.n241 10.6151
R1301 B.n301 B.n300 10.6151
R1302 B.n300 B.n299 10.6151
R1303 B.n299 B.n243 10.6151
R1304 B.n293 B.n292 10.6151
R1305 B.n292 B.n291 10.6151
R1306 B.n291 B.n248 10.6151
R1307 B.n285 B.n248 10.6151
R1308 B.n285 B.n284 10.6151
R1309 B.n284 B.n283 10.6151
R1310 B.n283 B.n250 10.6151
R1311 B.n277 B.n250 10.6151
R1312 B.n275 B.n274 10.6151
R1313 B.n274 B.n254 10.6151
R1314 B.n268 B.n254 10.6151
R1315 B.n268 B.n267 10.6151
R1316 B.n267 B.n266 10.6151
R1317 B.n266 B.n256 10.6151
R1318 B.n260 B.n256 10.6151
R1319 B.n260 B.n259 10.6151
R1320 B.n259 B.n235 10.6151
R1321 B.n319 B.n318 10.6151
R1322 B.n320 B.n319 10.6151
R1323 B.n320 B.n227 10.6151
R1324 B.n330 B.n227 10.6151
R1325 B.n331 B.n330 10.6151
R1326 B.n332 B.n331 10.6151
R1327 B.n332 B.n220 10.6151
R1328 B.n343 B.n220 10.6151
R1329 B.n344 B.n343 10.6151
R1330 B.n345 B.n344 10.6151
R1331 B.n345 B.n212 10.6151
R1332 B.n355 B.n212 10.6151
R1333 B.n356 B.n355 10.6151
R1334 B.n357 B.n356 10.6151
R1335 B.n357 B.n204 10.6151
R1336 B.n367 B.n204 10.6151
R1337 B.n368 B.n367 10.6151
R1338 B.n369 B.n368 10.6151
R1339 B.n369 B.n197 10.6151
R1340 B.n380 B.n197 10.6151
R1341 B.n381 B.n380 10.6151
R1342 B.n382 B.n381 10.6151
R1343 B.n382 B.n189 10.6151
R1344 B.n392 B.n189 10.6151
R1345 B.n393 B.n392 10.6151
R1346 B.n394 B.n393 10.6151
R1347 B.n394 B.n182 10.6151
R1348 B.n405 B.n182 10.6151
R1349 B.n406 B.n405 10.6151
R1350 B.n407 B.n406 10.6151
R1351 B.n407 B.n174 10.6151
R1352 B.n417 B.n174 10.6151
R1353 B.n418 B.n417 10.6151
R1354 B.n419 B.n418 10.6151
R1355 B.n419 B.n167 10.6151
R1356 B.n430 B.n167 10.6151
R1357 B.n431 B.n430 10.6151
R1358 B.n432 B.n431 10.6151
R1359 B.n432 B.n159 10.6151
R1360 B.n442 B.n159 10.6151
R1361 B.n443 B.n442 10.6151
R1362 B.n444 B.n443 10.6151
R1363 B.n444 B.n151 10.6151
R1364 B.n454 B.n151 10.6151
R1365 B.n455 B.n454 10.6151
R1366 B.n456 B.n455 10.6151
R1367 B.n456 B.n143 10.6151
R1368 B.n466 B.n143 10.6151
R1369 B.n467 B.n466 10.6151
R1370 B.n468 B.n467 10.6151
R1371 B.n468 B.n135 10.6151
R1372 B.n478 B.n135 10.6151
R1373 B.n479 B.n478 10.6151
R1374 B.n481 B.n479 10.6151
R1375 B.n481 B.n480 10.6151
R1376 B.n480 B.n127 10.6151
R1377 B.n492 B.n127 10.6151
R1378 B.n493 B.n492 10.6151
R1379 B.n494 B.n493 10.6151
R1380 B.n495 B.n494 10.6151
R1381 B.n496 B.n495 10.6151
R1382 B.n499 B.n496 10.6151
R1383 B.n500 B.n499 10.6151
R1384 B.n501 B.n500 10.6151
R1385 B.n502 B.n501 10.6151
R1386 B.n504 B.n502 10.6151
R1387 B.n505 B.n504 10.6151
R1388 B.n506 B.n505 10.6151
R1389 B.n507 B.n506 10.6151
R1390 B.n509 B.n507 10.6151
R1391 B.n510 B.n509 10.6151
R1392 B.n511 B.n510 10.6151
R1393 B.n512 B.n511 10.6151
R1394 B.n514 B.n512 10.6151
R1395 B.n515 B.n514 10.6151
R1396 B.n516 B.n515 10.6151
R1397 B.n517 B.n516 10.6151
R1398 B.n519 B.n517 10.6151
R1399 B.n520 B.n519 10.6151
R1400 B.n521 B.n520 10.6151
R1401 B.n522 B.n521 10.6151
R1402 B.n524 B.n522 10.6151
R1403 B.n525 B.n524 10.6151
R1404 B.n526 B.n525 10.6151
R1405 B.n527 B.n526 10.6151
R1406 B.n529 B.n527 10.6151
R1407 B.n530 B.n529 10.6151
R1408 B.n531 B.n530 10.6151
R1409 B.n532 B.n531 10.6151
R1410 B.n534 B.n532 10.6151
R1411 B.n535 B.n534 10.6151
R1412 B.n536 B.n535 10.6151
R1413 B.n537 B.n536 10.6151
R1414 B.n539 B.n537 10.6151
R1415 B.n540 B.n539 10.6151
R1416 B.n541 B.n540 10.6151
R1417 B.n542 B.n541 10.6151
R1418 B.n544 B.n542 10.6151
R1419 B.n545 B.n544 10.6151
R1420 B.n546 B.n545 10.6151
R1421 B.n547 B.n546 10.6151
R1422 B.n549 B.n547 10.6151
R1423 B.n550 B.n549 10.6151
R1424 B.n551 B.n550 10.6151
R1425 B.n552 B.n551 10.6151
R1426 B.n554 B.n552 10.6151
R1427 B.n555 B.n554 10.6151
R1428 B.n556 B.n555 10.6151
R1429 B.n557 B.n556 10.6151
R1430 B.n559 B.n557 10.6151
R1431 B.n560 B.n559 10.6151
R1432 B.n561 B.n560 10.6151
R1433 B.n562 B.n561 10.6151
R1434 B.n564 B.n562 10.6151
R1435 B.n565 B.n564 10.6151
R1436 B.n566 B.n565 10.6151
R1437 B.n567 B.n566 10.6151
R1438 B.n739 B.n1 10.6151
R1439 B.n739 B.n738 10.6151
R1440 B.n738 B.n737 10.6151
R1441 B.n737 B.n10 10.6151
R1442 B.n731 B.n10 10.6151
R1443 B.n731 B.n730 10.6151
R1444 B.n730 B.n729 10.6151
R1445 B.n729 B.n18 10.6151
R1446 B.n723 B.n18 10.6151
R1447 B.n723 B.n722 10.6151
R1448 B.n722 B.n721 10.6151
R1449 B.n721 B.n25 10.6151
R1450 B.n715 B.n25 10.6151
R1451 B.n715 B.n714 10.6151
R1452 B.n714 B.n713 10.6151
R1453 B.n713 B.n32 10.6151
R1454 B.n707 B.n32 10.6151
R1455 B.n707 B.n706 10.6151
R1456 B.n706 B.n705 10.6151
R1457 B.n705 B.n39 10.6151
R1458 B.n699 B.n39 10.6151
R1459 B.n699 B.n698 10.6151
R1460 B.n698 B.n697 10.6151
R1461 B.n697 B.n45 10.6151
R1462 B.n691 B.n45 10.6151
R1463 B.n691 B.n690 10.6151
R1464 B.n690 B.n689 10.6151
R1465 B.n689 B.n53 10.6151
R1466 B.n683 B.n53 10.6151
R1467 B.n683 B.n682 10.6151
R1468 B.n682 B.n681 10.6151
R1469 B.n681 B.n59 10.6151
R1470 B.n675 B.n59 10.6151
R1471 B.n675 B.n674 10.6151
R1472 B.n674 B.n673 10.6151
R1473 B.n673 B.n67 10.6151
R1474 B.n667 B.n67 10.6151
R1475 B.n667 B.n666 10.6151
R1476 B.n666 B.n665 10.6151
R1477 B.n665 B.n73 10.6151
R1478 B.n659 B.n73 10.6151
R1479 B.n659 B.n658 10.6151
R1480 B.n658 B.n657 10.6151
R1481 B.n657 B.n81 10.6151
R1482 B.n651 B.n81 10.6151
R1483 B.n651 B.n650 10.6151
R1484 B.n650 B.n649 10.6151
R1485 B.n649 B.n88 10.6151
R1486 B.n643 B.n88 10.6151
R1487 B.n643 B.n642 10.6151
R1488 B.n642 B.n641 10.6151
R1489 B.n641 B.n94 10.6151
R1490 B.n635 B.n94 10.6151
R1491 B.n635 B.n634 10.6151
R1492 B.n634 B.n633 10.6151
R1493 B.n633 B.n102 10.6151
R1494 B.n627 B.n102 10.6151
R1495 B.n626 B.n625 10.6151
R1496 B.n625 B.n109 10.6151
R1497 B.n619 B.n109 10.6151
R1498 B.n619 B.n618 10.6151
R1499 B.n618 B.n617 10.6151
R1500 B.n617 B.n111 10.6151
R1501 B.n611 B.n111 10.6151
R1502 B.n611 B.n610 10.6151
R1503 B.n610 B.n609 10.6151
R1504 B.n605 B.n604 10.6151
R1505 B.n604 B.n117 10.6151
R1506 B.n599 B.n117 10.6151
R1507 B.n599 B.n598 10.6151
R1508 B.n598 B.n597 10.6151
R1509 B.n597 B.n119 10.6151
R1510 B.n591 B.n119 10.6151
R1511 B.n591 B.n590 10.6151
R1512 B.n588 B.n123 10.6151
R1513 B.n582 B.n123 10.6151
R1514 B.n582 B.n581 10.6151
R1515 B.n581 B.n580 10.6151
R1516 B.n580 B.n125 10.6151
R1517 B.n574 B.n125 10.6151
R1518 B.n574 B.n573 10.6151
R1519 B.n573 B.n572 10.6151
R1520 B.n572 B.n568 10.6151
R1521 B.n747 B.n0 8.11757
R1522 B.n747 B.n1 8.11757
R1523 B.n428 B.t3 6.78539
R1524 B.n701 B.t6 6.78539
R1525 B.n293 B.n247 6.5566
R1526 B.n277 B.n276 6.5566
R1527 B.n605 B.n115 6.5566
R1528 B.n590 B.n589 6.5566
R1529 B.n247 B.n243 4.05904
R1530 B.n276 B.n275 4.05904
R1531 B.n609 B.n115 4.05904
R1532 B.n589 B.n588 4.05904
R1533 VN.n75 VN.n39 161.3
R1534 VN.n74 VN.n73 161.3
R1535 VN.n72 VN.n40 161.3
R1536 VN.n71 VN.n70 161.3
R1537 VN.n69 VN.n41 161.3
R1538 VN.n68 VN.n67 161.3
R1539 VN.n66 VN.n65 161.3
R1540 VN.n64 VN.n43 161.3
R1541 VN.n63 VN.n62 161.3
R1542 VN.n61 VN.n44 161.3
R1543 VN.n60 VN.n59 161.3
R1544 VN.n58 VN.n45 161.3
R1545 VN.n57 VN.n56 161.3
R1546 VN.n55 VN.n46 161.3
R1547 VN.n54 VN.n53 161.3
R1548 VN.n52 VN.n47 161.3
R1549 VN.n51 VN.n50 161.3
R1550 VN.n36 VN.n0 161.3
R1551 VN.n35 VN.n34 161.3
R1552 VN.n33 VN.n1 161.3
R1553 VN.n32 VN.n31 161.3
R1554 VN.n30 VN.n2 161.3
R1555 VN.n29 VN.n28 161.3
R1556 VN.n27 VN.n26 161.3
R1557 VN.n25 VN.n4 161.3
R1558 VN.n24 VN.n23 161.3
R1559 VN.n22 VN.n5 161.3
R1560 VN.n21 VN.n20 161.3
R1561 VN.n19 VN.n6 161.3
R1562 VN.n18 VN.n17 161.3
R1563 VN.n16 VN.n7 161.3
R1564 VN.n15 VN.n14 161.3
R1565 VN.n13 VN.n8 161.3
R1566 VN.n12 VN.n11 161.3
R1567 VN.n38 VN.n37 100.969
R1568 VN.n77 VN.n76 100.969
R1569 VN.n31 VN.n1 56.5193
R1570 VN.n70 VN.n40 56.5193
R1571 VN.n10 VN.n9 55.3127
R1572 VN.n49 VN.n48 55.3127
R1573 VN.n14 VN.n7 47.7779
R1574 VN.n24 VN.n5 47.7779
R1575 VN.n53 VN.n46 47.7779
R1576 VN.n63 VN.n44 47.7779
R1577 VN.n10 VN.t8 45.1187
R1578 VN.n49 VN.t6 45.1187
R1579 VN VN.n77 44.7822
R1580 VN.n14 VN.n13 33.2089
R1581 VN.n25 VN.n24 33.2089
R1582 VN.n53 VN.n52 33.2089
R1583 VN.n64 VN.n63 33.2089
R1584 VN.n13 VN.n12 24.4675
R1585 VN.n18 VN.n7 24.4675
R1586 VN.n19 VN.n18 24.4675
R1587 VN.n20 VN.n19 24.4675
R1588 VN.n20 VN.n5 24.4675
R1589 VN.n26 VN.n25 24.4675
R1590 VN.n30 VN.n29 24.4675
R1591 VN.n31 VN.n30 24.4675
R1592 VN.n35 VN.n1 24.4675
R1593 VN.n36 VN.n35 24.4675
R1594 VN.n52 VN.n51 24.4675
R1595 VN.n59 VN.n44 24.4675
R1596 VN.n59 VN.n58 24.4675
R1597 VN.n58 VN.n57 24.4675
R1598 VN.n57 VN.n46 24.4675
R1599 VN.n70 VN.n69 24.4675
R1600 VN.n69 VN.n68 24.4675
R1601 VN.n65 VN.n64 24.4675
R1602 VN.n75 VN.n74 24.4675
R1603 VN.n74 VN.n40 24.4675
R1604 VN.n12 VN.n9 17.1274
R1605 VN.n26 VN.n3 17.1274
R1606 VN.n51 VN.n48 17.1274
R1607 VN.n65 VN.n42 17.1274
R1608 VN.n19 VN.t9 11.5723
R1609 VN.n9 VN.t2 11.5723
R1610 VN.n3 VN.t7 11.5723
R1611 VN.n37 VN.t0 11.5723
R1612 VN.n58 VN.t4 11.5723
R1613 VN.n48 VN.t5 11.5723
R1614 VN.n42 VN.t3 11.5723
R1615 VN.n76 VN.t1 11.5723
R1616 VN.n37 VN.n36 9.7873
R1617 VN.n76 VN.n75 9.7873
R1618 VN.n29 VN.n3 7.3406
R1619 VN.n68 VN.n42 7.3406
R1620 VN.n50 VN.n49 6.86339
R1621 VN.n11 VN.n10 6.86339
R1622 VN.n77 VN.n39 0.278367
R1623 VN.n38 VN.n0 0.278367
R1624 VN.n73 VN.n39 0.189894
R1625 VN.n73 VN.n72 0.189894
R1626 VN.n72 VN.n71 0.189894
R1627 VN.n71 VN.n41 0.189894
R1628 VN.n67 VN.n41 0.189894
R1629 VN.n67 VN.n66 0.189894
R1630 VN.n66 VN.n43 0.189894
R1631 VN.n62 VN.n43 0.189894
R1632 VN.n62 VN.n61 0.189894
R1633 VN.n61 VN.n60 0.189894
R1634 VN.n60 VN.n45 0.189894
R1635 VN.n56 VN.n45 0.189894
R1636 VN.n56 VN.n55 0.189894
R1637 VN.n55 VN.n54 0.189894
R1638 VN.n54 VN.n47 0.189894
R1639 VN.n50 VN.n47 0.189894
R1640 VN.n11 VN.n8 0.189894
R1641 VN.n15 VN.n8 0.189894
R1642 VN.n16 VN.n15 0.189894
R1643 VN.n17 VN.n16 0.189894
R1644 VN.n17 VN.n6 0.189894
R1645 VN.n21 VN.n6 0.189894
R1646 VN.n22 VN.n21 0.189894
R1647 VN.n23 VN.n22 0.189894
R1648 VN.n23 VN.n4 0.189894
R1649 VN.n27 VN.n4 0.189894
R1650 VN.n28 VN.n27 0.189894
R1651 VN.n28 VN.n2 0.189894
R1652 VN.n32 VN.n2 0.189894
R1653 VN.n33 VN.n32 0.189894
R1654 VN.n34 VN.n33 0.189894
R1655 VN.n34 VN.n0 0.189894
R1656 VN VN.n38 0.153454
R1657 VDD2.n1 VDD2.t1 173.686
R1658 VDD2.n4 VDD2.t8 171.23
R1659 VDD2.n3 VDD2.n2 146.858
R1660 VDD2 VDD2.n7 146.856
R1661 VDD2.n1 VDD2.n0 145.071
R1662 VDD2.n6 VDD2.n5 145.071
R1663 VDD2.n4 VDD2.n3 36.4287
R1664 VDD2.n7 VDD2.t4 16.3641
R1665 VDD2.n7 VDD2.t3 16.3641
R1666 VDD2.n5 VDD2.t6 16.3641
R1667 VDD2.n5 VDD2.t5 16.3641
R1668 VDD2.n2 VDD2.t2 16.3641
R1669 VDD2.n2 VDD2.t9 16.3641
R1670 VDD2.n0 VDD2.t7 16.3641
R1671 VDD2.n0 VDD2.t0 16.3641
R1672 VDD2.n6 VDD2.n4 2.4574
R1673 VDD2 VDD2.n6 0.672914
R1674 VDD2.n3 VDD2.n1 0.559378
C0 VDD2 VP 0.582007f
C1 VN VDD1 0.160806f
C2 VN VTAIL 3.0226f
C3 VDD1 VTAIL 5.32167f
C4 VP VN 6.2915f
C5 VP VDD1 1.95485f
C6 VDD2 VN 1.53793f
C7 VDD2 VDD1 2.12098f
C8 VP VTAIL 3.03673f
C9 VDD2 VTAIL 5.37458f
C10 VDD2 B 5.210944f
C11 VDD1 B 5.159465f
C12 VTAIL B 3.314782f
C13 VN B 16.74843f
C14 VP B 15.264479f
C15 VDD2.t1 B 0.168635f
C16 VDD2.t7 B 0.024501f
C17 VDD2.t0 B 0.024501f
C18 VDD2.n0 B 0.122341f
C19 VDD2.n1 B 0.835739f
C20 VDD2.t2 B 0.024501f
C21 VDD2.t9 B 0.024501f
C22 VDD2.n2 B 0.128878f
C23 VDD2.n3 B 2.24721f
C24 VDD2.t8 B 0.162757f
C25 VDD2.n4 B 2.22004f
C26 VDD2.t6 B 0.024501f
C27 VDD2.t5 B 0.024501f
C28 VDD2.n5 B 0.122341f
C29 VDD2.n6 B 0.434361f
C30 VDD2.t4 B 0.024501f
C31 VDD2.t3 B 0.024501f
C32 VDD2.n7 B 0.128861f
C33 VN.n0 B 0.036877f
C34 VN.t0 B 0.173173f
C35 VN.n1 B 0.038887f
C36 VN.n2 B 0.027971f
C37 VN.t7 B 0.173173f
C38 VN.n3 B 0.10541f
C39 VN.n4 B 0.027971f
C40 VN.n5 B 0.052633f
C41 VN.n6 B 0.027971f
C42 VN.t9 B 0.173173f
C43 VN.n7 B 0.052633f
C44 VN.n8 B 0.027971f
C45 VN.t2 B 0.173173f
C46 VN.n9 B 0.190087f
C47 VN.t8 B 0.377628f
C48 VN.n10 B 0.179457f
C49 VN.n11 B 0.268122f
C50 VN.n12 B 0.04441f
C51 VN.n13 B 0.056466f
C52 VN.n14 B 0.024701f
C53 VN.n15 B 0.027971f
C54 VN.n16 B 0.027971f
C55 VN.n17 B 0.027971f
C56 VN.n18 B 0.052131f
C57 VN.n19 B 0.131804f
C58 VN.n20 B 0.052131f
C59 VN.n21 B 0.027971f
C60 VN.n22 B 0.027971f
C61 VN.n23 B 0.027971f
C62 VN.n24 B 0.024701f
C63 VN.n25 B 0.056466f
C64 VN.n26 B 0.04441f
C65 VN.n27 B 0.027971f
C66 VN.n28 B 0.027971f
C67 VN.n29 B 0.034115f
C68 VN.n30 B 0.052131f
C69 VN.n31 B 0.042784f
C70 VN.n32 B 0.027971f
C71 VN.n33 B 0.027971f
C72 VN.n34 B 0.027971f
C73 VN.n35 B 0.052131f
C74 VN.n36 B 0.036688f
C75 VN.n37 B 0.195889f
C76 VN.n38 B 0.044952f
C77 VN.n39 B 0.036877f
C78 VN.t1 B 0.173173f
C79 VN.n40 B 0.038887f
C80 VN.n41 B 0.027971f
C81 VN.t3 B 0.173173f
C82 VN.n42 B 0.10541f
C83 VN.n43 B 0.027971f
C84 VN.n44 B 0.052633f
C85 VN.n45 B 0.027971f
C86 VN.t4 B 0.173173f
C87 VN.n46 B 0.052633f
C88 VN.n47 B 0.027971f
C89 VN.t5 B 0.173173f
C90 VN.n48 B 0.190087f
C91 VN.t6 B 0.377628f
C92 VN.n49 B 0.179457f
C93 VN.n50 B 0.268122f
C94 VN.n51 B 0.04441f
C95 VN.n52 B 0.056466f
C96 VN.n53 B 0.024701f
C97 VN.n54 B 0.027971f
C98 VN.n55 B 0.027971f
C99 VN.n56 B 0.027971f
C100 VN.n57 B 0.052131f
C101 VN.n58 B 0.131804f
C102 VN.n59 B 0.052131f
C103 VN.n60 B 0.027971f
C104 VN.n61 B 0.027971f
C105 VN.n62 B 0.027971f
C106 VN.n63 B 0.024701f
C107 VN.n64 B 0.056466f
C108 VN.n65 B 0.04441f
C109 VN.n66 B 0.027971f
C110 VN.n67 B 0.027971f
C111 VN.n68 B 0.034115f
C112 VN.n69 B 0.052131f
C113 VN.n70 B 0.042784f
C114 VN.n71 B 0.027971f
C115 VN.n72 B 0.027971f
C116 VN.n73 B 0.027971f
C117 VN.n74 B 0.052131f
C118 VN.n75 B 0.036688f
C119 VN.n76 B 0.195889f
C120 VN.n77 B 1.31942f
C121 VDD1.t2 B 0.164313f
C122 VDD1.t3 B 0.023873f
C123 VDD1.t4 B 0.023873f
C124 VDD1.n0 B 0.119206f
C125 VDD1.n1 B 0.822418f
C126 VDD1.t7 B 0.164313f
C127 VDD1.t5 B 0.023873f
C128 VDD1.t0 B 0.023873f
C129 VDD1.n2 B 0.119206f
C130 VDD1.n3 B 0.81432f
C131 VDD1.t6 B 0.023873f
C132 VDD1.t1 B 0.023873f
C133 VDD1.n4 B 0.125575f
C134 VDD1.n5 B 2.3023f
C135 VDD1.t8 B 0.023873f
C136 VDD1.t9 B 0.023873f
C137 VDD1.n6 B 0.119206f
C138 VDD1.n7 B 2.26051f
C139 VTAIL.t13 B 0.038667f
C140 VTAIL.t0 B 0.038667f
C141 VTAIL.n0 B 0.157998f
C142 VTAIL.n1 B 0.726838f
C143 VTAIL.t8 B 0.223221f
C144 VTAIL.n2 B 0.839524f
C145 VTAIL.t9 B 0.038667f
C146 VTAIL.t10 B 0.038667f
C147 VTAIL.n3 B 0.157998f
C148 VTAIL.n4 B 0.898142f
C149 VTAIL.t7 B 0.038667f
C150 VTAIL.t4 B 0.038667f
C151 VTAIL.n5 B 0.157998f
C152 VTAIL.n6 B 1.90352f
C153 VTAIL.t1 B 0.038667f
C154 VTAIL.t16 B 0.038667f
C155 VTAIL.n7 B 0.157997f
C156 VTAIL.n8 B 1.90352f
C157 VTAIL.t19 B 0.038667f
C158 VTAIL.t17 B 0.038667f
C159 VTAIL.n9 B 0.157997f
C160 VTAIL.n10 B 0.898143f
C161 VTAIL.t15 B 0.223221f
C162 VTAIL.n11 B 0.839524f
C163 VTAIL.t12 B 0.038667f
C164 VTAIL.t11 B 0.038667f
C165 VTAIL.n12 B 0.157997f
C166 VTAIL.n13 B 0.799292f
C167 VTAIL.t6 B 0.038667f
C168 VTAIL.t3 B 0.038667f
C169 VTAIL.n14 B 0.157997f
C170 VTAIL.n15 B 0.898143f
C171 VTAIL.t5 B 0.223221f
C172 VTAIL.n16 B 1.62361f
C173 VTAIL.t2 B 0.223221f
C174 VTAIL.n17 B 1.62361f
C175 VTAIL.t18 B 0.038667f
C176 VTAIL.t14 B 0.038667f
C177 VTAIL.n18 B 0.157998f
C178 VTAIL.n19 B 0.650453f
C179 VP.n0 B 0.037033f
C180 VP.t8 B 0.173909f
C181 VP.n1 B 0.039052f
C182 VP.n2 B 0.02809f
C183 VP.t3 B 0.173909f
C184 VP.n3 B 0.105858f
C185 VP.n4 B 0.02809f
C186 VP.n5 B 0.052856f
C187 VP.n6 B 0.02809f
C188 VP.t9 B 0.173909f
C189 VP.n7 B 0.052856f
C190 VP.n8 B 0.02809f
C191 VP.t4 B 0.173909f
C192 VP.n9 B 0.105858f
C193 VP.n10 B 0.02809f
C194 VP.n11 B 0.039052f
C195 VP.n12 B 0.037033f
C196 VP.t2 B 0.173909f
C197 VP.n13 B 0.037033f
C198 VP.t0 B 0.173909f
C199 VP.n14 B 0.039052f
C200 VP.n15 B 0.02809f
C201 VP.t1 B 0.173909f
C202 VP.n16 B 0.105858f
C203 VP.n17 B 0.02809f
C204 VP.n18 B 0.052856f
C205 VP.n19 B 0.02809f
C206 VP.t5 B 0.173909f
C207 VP.n20 B 0.052856f
C208 VP.n21 B 0.02809f
C209 VP.t6 B 0.173909f
C210 VP.n22 B 0.190894f
C211 VP.t7 B 0.379231f
C212 VP.n23 B 0.180219f
C213 VP.n24 B 0.269261f
C214 VP.n25 B 0.044598f
C215 VP.n26 B 0.056706f
C216 VP.n27 B 0.024806f
C217 VP.n28 B 0.02809f
C218 VP.n29 B 0.02809f
C219 VP.n30 B 0.02809f
C220 VP.n31 B 0.052352f
C221 VP.n32 B 0.132363f
C222 VP.n33 B 0.052352f
C223 VP.n34 B 0.02809f
C224 VP.n35 B 0.02809f
C225 VP.n36 B 0.02809f
C226 VP.n37 B 0.024806f
C227 VP.n38 B 0.056706f
C228 VP.n39 B 0.044598f
C229 VP.n40 B 0.02809f
C230 VP.n41 B 0.02809f
C231 VP.n42 B 0.034259f
C232 VP.n43 B 0.052352f
C233 VP.n44 B 0.042965f
C234 VP.n45 B 0.02809f
C235 VP.n46 B 0.02809f
C236 VP.n47 B 0.02809f
C237 VP.n48 B 0.052352f
C238 VP.n49 B 0.036844f
C239 VP.n50 B 0.196721f
C240 VP.n51 B 1.30963f
C241 VP.n52 B 1.33232f
C242 VP.n53 B 0.196721f
C243 VP.n54 B 0.036844f
C244 VP.n55 B 0.052352f
C245 VP.n56 B 0.02809f
C246 VP.n57 B 0.02809f
C247 VP.n58 B 0.02809f
C248 VP.n59 B 0.042965f
C249 VP.n60 B 0.052352f
C250 VP.n61 B 0.034259f
C251 VP.n62 B 0.02809f
C252 VP.n63 B 0.02809f
C253 VP.n64 B 0.044598f
C254 VP.n65 B 0.056706f
C255 VP.n66 B 0.024806f
C256 VP.n67 B 0.02809f
C257 VP.n68 B 0.02809f
C258 VP.n69 B 0.02809f
C259 VP.n70 B 0.052352f
C260 VP.n71 B 0.132363f
C261 VP.n72 B 0.052352f
C262 VP.n73 B 0.02809f
C263 VP.n74 B 0.02809f
C264 VP.n75 B 0.02809f
C265 VP.n76 B 0.024806f
C266 VP.n77 B 0.056706f
C267 VP.n78 B 0.044598f
C268 VP.n79 B 0.02809f
C269 VP.n80 B 0.02809f
C270 VP.n81 B 0.034259f
C271 VP.n82 B 0.052352f
C272 VP.n83 B 0.042965f
C273 VP.n84 B 0.02809f
C274 VP.n85 B 0.02809f
C275 VP.n86 B 0.02809f
C276 VP.n87 B 0.052352f
C277 VP.n88 B 0.036844f
C278 VP.n89 B 0.196721f
C279 VP.n90 B 0.045143f
.ends

