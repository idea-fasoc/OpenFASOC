* NGSPICE file created from diff_pair_sample_0130.ext - technology: sky130A

.subckt diff_pair_sample_0130 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=1.27
X1 VTAIL.t19 VN.t1 VDD2.t8 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X2 VDD2.t7 VN.t2 VTAIL.t15 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=1.27
X3 VDD1.t9 VP.t0 VTAIL.t7 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X4 VTAIL.t16 VN.t3 VDD2.t6 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X5 VTAIL.t8 VP.t1 VDD1.t8 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X6 VDD2.t5 VN.t4 VTAIL.t11 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X7 VDD2.t4 VN.t5 VTAIL.t12 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=1.27
X8 VDD1.t7 VP.t2 VTAIL.t2 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=1.27
X9 VDD1.t6 VP.t3 VTAIL.t9 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=1.27
X10 VDD1.t5 VP.t4 VTAIL.t5 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=1.27
X11 B.t11 B.t9 B.t10 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=1.27
X12 VTAIL.t1 VP.t5 VDD1.t4 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X13 VTAIL.t10 VN.t6 VDD2.t3 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X14 B.t8 B.t6 B.t7 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=1.27
X15 VTAIL.t6 VP.t6 VDD1.t3 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X16 VTAIL.t17 VN.t7 VDD2.t2 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X17 B.t5 B.t3 B.t4 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=1.27
X18 VTAIL.t3 VP.t7 VDD1.t2 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X19 VDD1.t1 VP.t8 VTAIL.t4 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=1.27
X20 VDD2.t1 VN.t8 VTAIL.t14 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=1.27
X21 VDD2.t0 VN.t9 VTAIL.t13 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X22 VDD1.t0 VP.t9 VTAIL.t0 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=1.27
X23 B.t2 B.t0 B.t1 w_n2890_n2544# sky130_fd_pr__pfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=1.27
R0 VN.n6 VN.t0 176.614
R1 VN.n32 VN.t2 176.614
R2 VN.n24 VN.n23 175.833
R3 VN.n49 VN.n48 175.833
R4 VN.n47 VN.n25 161.3
R5 VN.n46 VN.n45 161.3
R6 VN.n44 VN.n26 161.3
R7 VN.n43 VN.n42 161.3
R8 VN.n41 VN.n27 161.3
R9 VN.n40 VN.n39 161.3
R10 VN.n38 VN.n29 161.3
R11 VN.n37 VN.n36 161.3
R12 VN.n35 VN.n30 161.3
R13 VN.n34 VN.n33 161.3
R14 VN.n22 VN.n0 161.3
R15 VN.n21 VN.n20 161.3
R16 VN.n19 VN.n1 161.3
R17 VN.n18 VN.n17 161.3
R18 VN.n15 VN.n2 161.3
R19 VN.n14 VN.n13 161.3
R20 VN.n12 VN.n3 161.3
R21 VN.n11 VN.n10 161.3
R22 VN.n9 VN.n4 161.3
R23 VN.n8 VN.n7 161.3
R24 VN.n3 VN.t9 149.345
R25 VN.n5 VN.t6 149.345
R26 VN.n16 VN.t1 149.345
R27 VN.n23 VN.t5 149.345
R28 VN.n29 VN.t4 149.345
R29 VN.n31 VN.t7 149.345
R30 VN.n28 VN.t3 149.345
R31 VN.n48 VN.t8 149.345
R32 VN.n6 VN.n5 60.024
R33 VN.n32 VN.n31 60.024
R34 VN.n10 VN.n9 56.4357
R35 VN.n15 VN.n14 56.4357
R36 VN.n36 VN.n35 56.4357
R37 VN.n41 VN.n40 56.4357
R38 VN.n21 VN.n1 50.0905
R39 VN.n46 VN.n26 50.0905
R40 VN VN.n49 43.01
R41 VN.n22 VN.n21 30.5668
R42 VN.n47 VN.n46 30.5668
R43 VN.n33 VN.n32 27.7309
R44 VN.n7 VN.n6 27.7309
R45 VN.n9 VN.n8 24.2216
R46 VN.n10 VN.n3 24.2216
R47 VN.n14 VN.n3 24.2216
R48 VN.n17 VN.n15 24.2216
R49 VN.n35 VN.n34 24.2216
R50 VN.n40 VN.n29 24.2216
R51 VN.n36 VN.n29 24.2216
R52 VN.n42 VN.n41 24.2216
R53 VN.n16 VN.n1 19.3774
R54 VN.n28 VN.n26 19.3774
R55 VN.n23 VN.n22 9.68894
R56 VN.n48 VN.n47 9.68894
R57 VN.n8 VN.n5 4.84472
R58 VN.n17 VN.n16 4.84472
R59 VN.n34 VN.n31 4.84472
R60 VN.n42 VN.n28 4.84472
R61 VN.n49 VN.n25 0.189894
R62 VN.n45 VN.n25 0.189894
R63 VN.n45 VN.n44 0.189894
R64 VN.n44 VN.n43 0.189894
R65 VN.n43 VN.n27 0.189894
R66 VN.n39 VN.n27 0.189894
R67 VN.n39 VN.n38 0.189894
R68 VN.n38 VN.n37 0.189894
R69 VN.n37 VN.n30 0.189894
R70 VN.n33 VN.n30 0.189894
R71 VN.n7 VN.n4 0.189894
R72 VN.n11 VN.n4 0.189894
R73 VN.n12 VN.n11 0.189894
R74 VN.n13 VN.n12 0.189894
R75 VN.n13 VN.n2 0.189894
R76 VN.n18 VN.n2 0.189894
R77 VN.n19 VN.n18 0.189894
R78 VN.n20 VN.n19 0.189894
R79 VN.n20 VN.n0 0.189894
R80 VN.n24 VN.n0 0.189894
R81 VN VN.n24 0.0516364
R82 VTAIL.n176 VTAIL.n140 756.745
R83 VTAIL.n38 VTAIL.n2 756.745
R84 VTAIL.n134 VTAIL.n98 756.745
R85 VTAIL.n88 VTAIL.n52 756.745
R86 VTAIL.n152 VTAIL.n151 585
R87 VTAIL.n157 VTAIL.n156 585
R88 VTAIL.n159 VTAIL.n158 585
R89 VTAIL.n148 VTAIL.n147 585
R90 VTAIL.n165 VTAIL.n164 585
R91 VTAIL.n167 VTAIL.n166 585
R92 VTAIL.n144 VTAIL.n143 585
R93 VTAIL.n174 VTAIL.n173 585
R94 VTAIL.n175 VTAIL.n142 585
R95 VTAIL.n177 VTAIL.n176 585
R96 VTAIL.n14 VTAIL.n13 585
R97 VTAIL.n19 VTAIL.n18 585
R98 VTAIL.n21 VTAIL.n20 585
R99 VTAIL.n10 VTAIL.n9 585
R100 VTAIL.n27 VTAIL.n26 585
R101 VTAIL.n29 VTAIL.n28 585
R102 VTAIL.n6 VTAIL.n5 585
R103 VTAIL.n36 VTAIL.n35 585
R104 VTAIL.n37 VTAIL.n4 585
R105 VTAIL.n39 VTAIL.n38 585
R106 VTAIL.n135 VTAIL.n134 585
R107 VTAIL.n133 VTAIL.n100 585
R108 VTAIL.n132 VTAIL.n131 585
R109 VTAIL.n103 VTAIL.n101 585
R110 VTAIL.n126 VTAIL.n125 585
R111 VTAIL.n124 VTAIL.n123 585
R112 VTAIL.n107 VTAIL.n106 585
R113 VTAIL.n118 VTAIL.n117 585
R114 VTAIL.n116 VTAIL.n115 585
R115 VTAIL.n111 VTAIL.n110 585
R116 VTAIL.n89 VTAIL.n88 585
R117 VTAIL.n87 VTAIL.n54 585
R118 VTAIL.n86 VTAIL.n85 585
R119 VTAIL.n57 VTAIL.n55 585
R120 VTAIL.n80 VTAIL.n79 585
R121 VTAIL.n78 VTAIL.n77 585
R122 VTAIL.n61 VTAIL.n60 585
R123 VTAIL.n72 VTAIL.n71 585
R124 VTAIL.n70 VTAIL.n69 585
R125 VTAIL.n65 VTAIL.n64 585
R126 VTAIL.n153 VTAIL.t12 329.043
R127 VTAIL.n15 VTAIL.t2 329.043
R128 VTAIL.n112 VTAIL.t9 329.043
R129 VTAIL.n66 VTAIL.t15 329.043
R130 VTAIL.n157 VTAIL.n151 171.744
R131 VTAIL.n158 VTAIL.n157 171.744
R132 VTAIL.n158 VTAIL.n147 171.744
R133 VTAIL.n165 VTAIL.n147 171.744
R134 VTAIL.n166 VTAIL.n165 171.744
R135 VTAIL.n166 VTAIL.n143 171.744
R136 VTAIL.n174 VTAIL.n143 171.744
R137 VTAIL.n175 VTAIL.n174 171.744
R138 VTAIL.n176 VTAIL.n175 171.744
R139 VTAIL.n19 VTAIL.n13 171.744
R140 VTAIL.n20 VTAIL.n19 171.744
R141 VTAIL.n20 VTAIL.n9 171.744
R142 VTAIL.n27 VTAIL.n9 171.744
R143 VTAIL.n28 VTAIL.n27 171.744
R144 VTAIL.n28 VTAIL.n5 171.744
R145 VTAIL.n36 VTAIL.n5 171.744
R146 VTAIL.n37 VTAIL.n36 171.744
R147 VTAIL.n38 VTAIL.n37 171.744
R148 VTAIL.n134 VTAIL.n133 171.744
R149 VTAIL.n133 VTAIL.n132 171.744
R150 VTAIL.n132 VTAIL.n101 171.744
R151 VTAIL.n125 VTAIL.n101 171.744
R152 VTAIL.n125 VTAIL.n124 171.744
R153 VTAIL.n124 VTAIL.n106 171.744
R154 VTAIL.n117 VTAIL.n106 171.744
R155 VTAIL.n117 VTAIL.n116 171.744
R156 VTAIL.n116 VTAIL.n110 171.744
R157 VTAIL.n88 VTAIL.n87 171.744
R158 VTAIL.n87 VTAIL.n86 171.744
R159 VTAIL.n86 VTAIL.n55 171.744
R160 VTAIL.n79 VTAIL.n55 171.744
R161 VTAIL.n79 VTAIL.n78 171.744
R162 VTAIL.n78 VTAIL.n60 171.744
R163 VTAIL.n71 VTAIL.n60 171.744
R164 VTAIL.n71 VTAIL.n70 171.744
R165 VTAIL.n70 VTAIL.n64 171.744
R166 VTAIL.t12 VTAIL.n151 85.8723
R167 VTAIL.t2 VTAIL.n13 85.8723
R168 VTAIL.t9 VTAIL.n110 85.8723
R169 VTAIL.t15 VTAIL.n64 85.8723
R170 VTAIL.n97 VTAIL.n96 67.038
R171 VTAIL.n95 VTAIL.n94 67.038
R172 VTAIL.n51 VTAIL.n50 67.038
R173 VTAIL.n49 VTAIL.n48 67.038
R174 VTAIL.n183 VTAIL.n182 67.0378
R175 VTAIL.n1 VTAIL.n0 67.0378
R176 VTAIL.n45 VTAIL.n44 67.0378
R177 VTAIL.n47 VTAIL.n46 67.0378
R178 VTAIL.n181 VTAIL.n180 33.5429
R179 VTAIL.n43 VTAIL.n42 33.5429
R180 VTAIL.n139 VTAIL.n138 33.5429
R181 VTAIL.n93 VTAIL.n92 33.5429
R182 VTAIL.n49 VTAIL.n47 21.9186
R183 VTAIL.n181 VTAIL.n139 20.5393
R184 VTAIL.n177 VTAIL.n142 13.1884
R185 VTAIL.n39 VTAIL.n4 13.1884
R186 VTAIL.n135 VTAIL.n100 13.1884
R187 VTAIL.n89 VTAIL.n54 13.1884
R188 VTAIL.n173 VTAIL.n172 12.8005
R189 VTAIL.n178 VTAIL.n140 12.8005
R190 VTAIL.n35 VTAIL.n34 12.8005
R191 VTAIL.n40 VTAIL.n2 12.8005
R192 VTAIL.n136 VTAIL.n98 12.8005
R193 VTAIL.n131 VTAIL.n102 12.8005
R194 VTAIL.n90 VTAIL.n52 12.8005
R195 VTAIL.n85 VTAIL.n56 12.8005
R196 VTAIL.n171 VTAIL.n144 12.0247
R197 VTAIL.n33 VTAIL.n6 12.0247
R198 VTAIL.n130 VTAIL.n103 12.0247
R199 VTAIL.n84 VTAIL.n57 12.0247
R200 VTAIL.n168 VTAIL.n167 11.249
R201 VTAIL.n30 VTAIL.n29 11.249
R202 VTAIL.n127 VTAIL.n126 11.249
R203 VTAIL.n81 VTAIL.n80 11.249
R204 VTAIL.n153 VTAIL.n152 10.7238
R205 VTAIL.n15 VTAIL.n14 10.7238
R206 VTAIL.n112 VTAIL.n111 10.7238
R207 VTAIL.n66 VTAIL.n65 10.7238
R208 VTAIL.n164 VTAIL.n146 10.4732
R209 VTAIL.n26 VTAIL.n8 10.4732
R210 VTAIL.n123 VTAIL.n105 10.4732
R211 VTAIL.n77 VTAIL.n59 10.4732
R212 VTAIL.n163 VTAIL.n148 9.69747
R213 VTAIL.n25 VTAIL.n10 9.69747
R214 VTAIL.n122 VTAIL.n107 9.69747
R215 VTAIL.n76 VTAIL.n61 9.69747
R216 VTAIL.n180 VTAIL.n179 9.45567
R217 VTAIL.n42 VTAIL.n41 9.45567
R218 VTAIL.n138 VTAIL.n137 9.45567
R219 VTAIL.n92 VTAIL.n91 9.45567
R220 VTAIL.n179 VTAIL.n178 9.3005
R221 VTAIL.n155 VTAIL.n154 9.3005
R222 VTAIL.n150 VTAIL.n149 9.3005
R223 VTAIL.n161 VTAIL.n160 9.3005
R224 VTAIL.n163 VTAIL.n162 9.3005
R225 VTAIL.n146 VTAIL.n145 9.3005
R226 VTAIL.n169 VTAIL.n168 9.3005
R227 VTAIL.n171 VTAIL.n170 9.3005
R228 VTAIL.n172 VTAIL.n141 9.3005
R229 VTAIL.n41 VTAIL.n40 9.3005
R230 VTAIL.n17 VTAIL.n16 9.3005
R231 VTAIL.n12 VTAIL.n11 9.3005
R232 VTAIL.n23 VTAIL.n22 9.3005
R233 VTAIL.n25 VTAIL.n24 9.3005
R234 VTAIL.n8 VTAIL.n7 9.3005
R235 VTAIL.n31 VTAIL.n30 9.3005
R236 VTAIL.n33 VTAIL.n32 9.3005
R237 VTAIL.n34 VTAIL.n3 9.3005
R238 VTAIL.n114 VTAIL.n113 9.3005
R239 VTAIL.n109 VTAIL.n108 9.3005
R240 VTAIL.n120 VTAIL.n119 9.3005
R241 VTAIL.n122 VTAIL.n121 9.3005
R242 VTAIL.n105 VTAIL.n104 9.3005
R243 VTAIL.n128 VTAIL.n127 9.3005
R244 VTAIL.n130 VTAIL.n129 9.3005
R245 VTAIL.n102 VTAIL.n99 9.3005
R246 VTAIL.n137 VTAIL.n136 9.3005
R247 VTAIL.n68 VTAIL.n67 9.3005
R248 VTAIL.n63 VTAIL.n62 9.3005
R249 VTAIL.n74 VTAIL.n73 9.3005
R250 VTAIL.n76 VTAIL.n75 9.3005
R251 VTAIL.n59 VTAIL.n58 9.3005
R252 VTAIL.n82 VTAIL.n81 9.3005
R253 VTAIL.n84 VTAIL.n83 9.3005
R254 VTAIL.n56 VTAIL.n53 9.3005
R255 VTAIL.n91 VTAIL.n90 9.3005
R256 VTAIL.n160 VTAIL.n159 8.92171
R257 VTAIL.n22 VTAIL.n21 8.92171
R258 VTAIL.n119 VTAIL.n118 8.92171
R259 VTAIL.n73 VTAIL.n72 8.92171
R260 VTAIL.n156 VTAIL.n150 8.14595
R261 VTAIL.n18 VTAIL.n12 8.14595
R262 VTAIL.n115 VTAIL.n109 8.14595
R263 VTAIL.n69 VTAIL.n63 8.14595
R264 VTAIL.n155 VTAIL.n152 7.3702
R265 VTAIL.n17 VTAIL.n14 7.3702
R266 VTAIL.n114 VTAIL.n111 7.3702
R267 VTAIL.n68 VTAIL.n65 7.3702
R268 VTAIL.n156 VTAIL.n155 5.81868
R269 VTAIL.n18 VTAIL.n17 5.81868
R270 VTAIL.n115 VTAIL.n114 5.81868
R271 VTAIL.n69 VTAIL.n68 5.81868
R272 VTAIL.n159 VTAIL.n150 5.04292
R273 VTAIL.n21 VTAIL.n12 5.04292
R274 VTAIL.n118 VTAIL.n109 5.04292
R275 VTAIL.n72 VTAIL.n63 5.04292
R276 VTAIL.n160 VTAIL.n148 4.26717
R277 VTAIL.n22 VTAIL.n10 4.26717
R278 VTAIL.n119 VTAIL.n107 4.26717
R279 VTAIL.n73 VTAIL.n61 4.26717
R280 VTAIL.n182 VTAIL.t13 4.13074
R281 VTAIL.n182 VTAIL.t19 4.13074
R282 VTAIL.n0 VTAIL.t18 4.13074
R283 VTAIL.n0 VTAIL.t10 4.13074
R284 VTAIL.n44 VTAIL.t0 4.13074
R285 VTAIL.n44 VTAIL.t1 4.13074
R286 VTAIL.n46 VTAIL.t5 4.13074
R287 VTAIL.n46 VTAIL.t8 4.13074
R288 VTAIL.n96 VTAIL.t7 4.13074
R289 VTAIL.n96 VTAIL.t3 4.13074
R290 VTAIL.n94 VTAIL.t4 4.13074
R291 VTAIL.n94 VTAIL.t6 4.13074
R292 VTAIL.n50 VTAIL.t11 4.13074
R293 VTAIL.n50 VTAIL.t17 4.13074
R294 VTAIL.n48 VTAIL.t14 4.13074
R295 VTAIL.n48 VTAIL.t16 4.13074
R296 VTAIL.n164 VTAIL.n163 3.49141
R297 VTAIL.n26 VTAIL.n25 3.49141
R298 VTAIL.n123 VTAIL.n122 3.49141
R299 VTAIL.n77 VTAIL.n76 3.49141
R300 VTAIL.n167 VTAIL.n146 2.71565
R301 VTAIL.n29 VTAIL.n8 2.71565
R302 VTAIL.n126 VTAIL.n105 2.71565
R303 VTAIL.n80 VTAIL.n59 2.71565
R304 VTAIL.n154 VTAIL.n153 2.4129
R305 VTAIL.n16 VTAIL.n15 2.4129
R306 VTAIL.n113 VTAIL.n112 2.4129
R307 VTAIL.n67 VTAIL.n66 2.4129
R308 VTAIL.n168 VTAIL.n144 1.93989
R309 VTAIL.n30 VTAIL.n6 1.93989
R310 VTAIL.n127 VTAIL.n103 1.93989
R311 VTAIL.n81 VTAIL.n57 1.93989
R312 VTAIL.n51 VTAIL.n49 1.37981
R313 VTAIL.n93 VTAIL.n51 1.37981
R314 VTAIL.n97 VTAIL.n95 1.37981
R315 VTAIL.n139 VTAIL.n97 1.37981
R316 VTAIL.n47 VTAIL.n45 1.37981
R317 VTAIL.n45 VTAIL.n43 1.37981
R318 VTAIL.n183 VTAIL.n181 1.37981
R319 VTAIL.n173 VTAIL.n171 1.16414
R320 VTAIL.n180 VTAIL.n140 1.16414
R321 VTAIL.n35 VTAIL.n33 1.16414
R322 VTAIL.n42 VTAIL.n2 1.16414
R323 VTAIL.n138 VTAIL.n98 1.16414
R324 VTAIL.n131 VTAIL.n130 1.16414
R325 VTAIL.n92 VTAIL.n52 1.16414
R326 VTAIL.n85 VTAIL.n84 1.16414
R327 VTAIL.n95 VTAIL.n93 1.15998
R328 VTAIL.n43 VTAIL.n1 1.15998
R329 VTAIL VTAIL.n1 1.09317
R330 VTAIL.n172 VTAIL.n142 0.388379
R331 VTAIL.n178 VTAIL.n177 0.388379
R332 VTAIL.n34 VTAIL.n4 0.388379
R333 VTAIL.n40 VTAIL.n39 0.388379
R334 VTAIL.n136 VTAIL.n135 0.388379
R335 VTAIL.n102 VTAIL.n100 0.388379
R336 VTAIL.n90 VTAIL.n89 0.388379
R337 VTAIL.n56 VTAIL.n54 0.388379
R338 VTAIL VTAIL.n183 0.287138
R339 VTAIL.n154 VTAIL.n149 0.155672
R340 VTAIL.n161 VTAIL.n149 0.155672
R341 VTAIL.n162 VTAIL.n161 0.155672
R342 VTAIL.n162 VTAIL.n145 0.155672
R343 VTAIL.n169 VTAIL.n145 0.155672
R344 VTAIL.n170 VTAIL.n169 0.155672
R345 VTAIL.n170 VTAIL.n141 0.155672
R346 VTAIL.n179 VTAIL.n141 0.155672
R347 VTAIL.n16 VTAIL.n11 0.155672
R348 VTAIL.n23 VTAIL.n11 0.155672
R349 VTAIL.n24 VTAIL.n23 0.155672
R350 VTAIL.n24 VTAIL.n7 0.155672
R351 VTAIL.n31 VTAIL.n7 0.155672
R352 VTAIL.n32 VTAIL.n31 0.155672
R353 VTAIL.n32 VTAIL.n3 0.155672
R354 VTAIL.n41 VTAIL.n3 0.155672
R355 VTAIL.n137 VTAIL.n99 0.155672
R356 VTAIL.n129 VTAIL.n99 0.155672
R357 VTAIL.n129 VTAIL.n128 0.155672
R358 VTAIL.n128 VTAIL.n104 0.155672
R359 VTAIL.n121 VTAIL.n104 0.155672
R360 VTAIL.n121 VTAIL.n120 0.155672
R361 VTAIL.n120 VTAIL.n108 0.155672
R362 VTAIL.n113 VTAIL.n108 0.155672
R363 VTAIL.n91 VTAIL.n53 0.155672
R364 VTAIL.n83 VTAIL.n53 0.155672
R365 VTAIL.n83 VTAIL.n82 0.155672
R366 VTAIL.n82 VTAIL.n58 0.155672
R367 VTAIL.n75 VTAIL.n58 0.155672
R368 VTAIL.n75 VTAIL.n74 0.155672
R369 VTAIL.n74 VTAIL.n62 0.155672
R370 VTAIL.n67 VTAIL.n62 0.155672
R371 VDD2.n81 VDD2.n45 756.745
R372 VDD2.n36 VDD2.n0 756.745
R373 VDD2.n82 VDD2.n81 585
R374 VDD2.n80 VDD2.n47 585
R375 VDD2.n79 VDD2.n78 585
R376 VDD2.n50 VDD2.n48 585
R377 VDD2.n73 VDD2.n72 585
R378 VDD2.n71 VDD2.n70 585
R379 VDD2.n54 VDD2.n53 585
R380 VDD2.n65 VDD2.n64 585
R381 VDD2.n63 VDD2.n62 585
R382 VDD2.n58 VDD2.n57 585
R383 VDD2.n12 VDD2.n11 585
R384 VDD2.n17 VDD2.n16 585
R385 VDD2.n19 VDD2.n18 585
R386 VDD2.n8 VDD2.n7 585
R387 VDD2.n25 VDD2.n24 585
R388 VDD2.n27 VDD2.n26 585
R389 VDD2.n4 VDD2.n3 585
R390 VDD2.n34 VDD2.n33 585
R391 VDD2.n35 VDD2.n2 585
R392 VDD2.n37 VDD2.n36 585
R393 VDD2.n59 VDD2.t1 329.043
R394 VDD2.n13 VDD2.t9 329.043
R395 VDD2.n81 VDD2.n80 171.744
R396 VDD2.n80 VDD2.n79 171.744
R397 VDD2.n79 VDD2.n48 171.744
R398 VDD2.n72 VDD2.n48 171.744
R399 VDD2.n72 VDD2.n71 171.744
R400 VDD2.n71 VDD2.n53 171.744
R401 VDD2.n64 VDD2.n53 171.744
R402 VDD2.n64 VDD2.n63 171.744
R403 VDD2.n63 VDD2.n57 171.744
R404 VDD2.n17 VDD2.n11 171.744
R405 VDD2.n18 VDD2.n17 171.744
R406 VDD2.n18 VDD2.n7 171.744
R407 VDD2.n25 VDD2.n7 171.744
R408 VDD2.n26 VDD2.n25 171.744
R409 VDD2.n26 VDD2.n3 171.744
R410 VDD2.n34 VDD2.n3 171.744
R411 VDD2.n35 VDD2.n34 171.744
R412 VDD2.n36 VDD2.n35 171.744
R413 VDD2.t1 VDD2.n57 85.8723
R414 VDD2.t9 VDD2.n11 85.8723
R415 VDD2.n44 VDD2.n43 84.6958
R416 VDD2 VDD2.n89 84.6929
R417 VDD2.n88 VDD2.n87 83.7168
R418 VDD2.n42 VDD2.n41 83.7166
R419 VDD2.n42 VDD2.n40 51.601
R420 VDD2.n86 VDD2.n85 50.2217
R421 VDD2.n86 VDD2.n44 37.0601
R422 VDD2.n82 VDD2.n47 13.1884
R423 VDD2.n37 VDD2.n2 13.1884
R424 VDD2.n83 VDD2.n45 12.8005
R425 VDD2.n78 VDD2.n49 12.8005
R426 VDD2.n33 VDD2.n32 12.8005
R427 VDD2.n38 VDD2.n0 12.8005
R428 VDD2.n77 VDD2.n50 12.0247
R429 VDD2.n31 VDD2.n4 12.0247
R430 VDD2.n74 VDD2.n73 11.249
R431 VDD2.n28 VDD2.n27 11.249
R432 VDD2.n59 VDD2.n58 10.7238
R433 VDD2.n13 VDD2.n12 10.7238
R434 VDD2.n70 VDD2.n52 10.4732
R435 VDD2.n24 VDD2.n6 10.4732
R436 VDD2.n69 VDD2.n54 9.69747
R437 VDD2.n23 VDD2.n8 9.69747
R438 VDD2.n85 VDD2.n84 9.45567
R439 VDD2.n40 VDD2.n39 9.45567
R440 VDD2.n61 VDD2.n60 9.3005
R441 VDD2.n56 VDD2.n55 9.3005
R442 VDD2.n67 VDD2.n66 9.3005
R443 VDD2.n69 VDD2.n68 9.3005
R444 VDD2.n52 VDD2.n51 9.3005
R445 VDD2.n75 VDD2.n74 9.3005
R446 VDD2.n77 VDD2.n76 9.3005
R447 VDD2.n49 VDD2.n46 9.3005
R448 VDD2.n84 VDD2.n83 9.3005
R449 VDD2.n39 VDD2.n38 9.3005
R450 VDD2.n15 VDD2.n14 9.3005
R451 VDD2.n10 VDD2.n9 9.3005
R452 VDD2.n21 VDD2.n20 9.3005
R453 VDD2.n23 VDD2.n22 9.3005
R454 VDD2.n6 VDD2.n5 9.3005
R455 VDD2.n29 VDD2.n28 9.3005
R456 VDD2.n31 VDD2.n30 9.3005
R457 VDD2.n32 VDD2.n1 9.3005
R458 VDD2.n66 VDD2.n65 8.92171
R459 VDD2.n20 VDD2.n19 8.92171
R460 VDD2.n62 VDD2.n56 8.14595
R461 VDD2.n16 VDD2.n10 8.14595
R462 VDD2.n61 VDD2.n58 7.3702
R463 VDD2.n15 VDD2.n12 7.3702
R464 VDD2.n62 VDD2.n61 5.81868
R465 VDD2.n16 VDD2.n15 5.81868
R466 VDD2.n65 VDD2.n56 5.04292
R467 VDD2.n19 VDD2.n10 5.04292
R468 VDD2.n66 VDD2.n54 4.26717
R469 VDD2.n20 VDD2.n8 4.26717
R470 VDD2.n89 VDD2.t2 4.13074
R471 VDD2.n89 VDD2.t7 4.13074
R472 VDD2.n87 VDD2.t6 4.13074
R473 VDD2.n87 VDD2.t5 4.13074
R474 VDD2.n43 VDD2.t8 4.13074
R475 VDD2.n43 VDD2.t4 4.13074
R476 VDD2.n41 VDD2.t3 4.13074
R477 VDD2.n41 VDD2.t0 4.13074
R478 VDD2.n70 VDD2.n69 3.49141
R479 VDD2.n24 VDD2.n23 3.49141
R480 VDD2.n73 VDD2.n52 2.71565
R481 VDD2.n27 VDD2.n6 2.71565
R482 VDD2.n60 VDD2.n59 2.4129
R483 VDD2.n14 VDD2.n13 2.4129
R484 VDD2.n74 VDD2.n50 1.93989
R485 VDD2.n28 VDD2.n4 1.93989
R486 VDD2.n88 VDD2.n86 1.37981
R487 VDD2.n85 VDD2.n45 1.16414
R488 VDD2.n78 VDD2.n77 1.16414
R489 VDD2.n33 VDD2.n31 1.16414
R490 VDD2.n40 VDD2.n0 1.16414
R491 VDD2 VDD2.n88 0.403517
R492 VDD2.n83 VDD2.n82 0.388379
R493 VDD2.n49 VDD2.n47 0.388379
R494 VDD2.n32 VDD2.n2 0.388379
R495 VDD2.n38 VDD2.n37 0.388379
R496 VDD2.n44 VDD2.n42 0.289982
R497 VDD2.n84 VDD2.n46 0.155672
R498 VDD2.n76 VDD2.n46 0.155672
R499 VDD2.n76 VDD2.n75 0.155672
R500 VDD2.n75 VDD2.n51 0.155672
R501 VDD2.n68 VDD2.n51 0.155672
R502 VDD2.n68 VDD2.n67 0.155672
R503 VDD2.n67 VDD2.n55 0.155672
R504 VDD2.n60 VDD2.n55 0.155672
R505 VDD2.n14 VDD2.n9 0.155672
R506 VDD2.n21 VDD2.n9 0.155672
R507 VDD2.n22 VDD2.n21 0.155672
R508 VDD2.n22 VDD2.n5 0.155672
R509 VDD2.n29 VDD2.n5 0.155672
R510 VDD2.n30 VDD2.n29 0.155672
R511 VDD2.n30 VDD2.n1 0.155672
R512 VDD2.n39 VDD2.n1 0.155672
R513 VP.n14 VP.t8 176.614
R514 VP.n33 VP.n7 175.833
R515 VP.n56 VP.n55 175.833
R516 VP.n32 VP.n31 175.833
R517 VP.n16 VP.n15 161.3
R518 VP.n17 VP.n12 161.3
R519 VP.n19 VP.n18 161.3
R520 VP.n20 VP.n11 161.3
R521 VP.n22 VP.n21 161.3
R522 VP.n23 VP.n10 161.3
R523 VP.n26 VP.n25 161.3
R524 VP.n27 VP.n9 161.3
R525 VP.n29 VP.n28 161.3
R526 VP.n30 VP.n8 161.3
R527 VP.n54 VP.n0 161.3
R528 VP.n53 VP.n52 161.3
R529 VP.n51 VP.n1 161.3
R530 VP.n50 VP.n49 161.3
R531 VP.n47 VP.n2 161.3
R532 VP.n46 VP.n45 161.3
R533 VP.n44 VP.n3 161.3
R534 VP.n43 VP.n42 161.3
R535 VP.n41 VP.n4 161.3
R536 VP.n40 VP.n39 161.3
R537 VP.n38 VP.n37 161.3
R538 VP.n36 VP.n6 161.3
R539 VP.n35 VP.n34 161.3
R540 VP.n3 VP.t9 149.345
R541 VP.n7 VP.t4 149.345
R542 VP.n5 VP.t1 149.345
R543 VP.n48 VP.t5 149.345
R544 VP.n55 VP.t2 149.345
R545 VP.n11 VP.t0 149.345
R546 VP.n31 VP.t3 149.345
R547 VP.n24 VP.t7 149.345
R548 VP.n13 VP.t6 149.345
R549 VP.n14 VP.n13 60.024
R550 VP.n42 VP.n41 56.4357
R551 VP.n47 VP.n46 56.4357
R552 VP.n23 VP.n22 56.4357
R553 VP.n18 VP.n17 56.4357
R554 VP.n37 VP.n36 50.0905
R555 VP.n53 VP.n1 50.0905
R556 VP.n29 VP.n9 50.0905
R557 VP.n33 VP.n32 42.6293
R558 VP.n36 VP.n35 30.5668
R559 VP.n54 VP.n53 30.5668
R560 VP.n30 VP.n29 30.5668
R561 VP.n15 VP.n14 27.7309
R562 VP.n41 VP.n40 24.2216
R563 VP.n42 VP.n3 24.2216
R564 VP.n46 VP.n3 24.2216
R565 VP.n49 VP.n47 24.2216
R566 VP.n25 VP.n23 24.2216
R567 VP.n18 VP.n11 24.2216
R568 VP.n22 VP.n11 24.2216
R569 VP.n17 VP.n16 24.2216
R570 VP.n37 VP.n5 19.3774
R571 VP.n48 VP.n1 19.3774
R572 VP.n24 VP.n9 19.3774
R573 VP.n35 VP.n7 9.68894
R574 VP.n55 VP.n54 9.68894
R575 VP.n31 VP.n30 9.68894
R576 VP.n40 VP.n5 4.84472
R577 VP.n49 VP.n48 4.84472
R578 VP.n25 VP.n24 4.84472
R579 VP.n16 VP.n13 4.84472
R580 VP.n15 VP.n12 0.189894
R581 VP.n19 VP.n12 0.189894
R582 VP.n20 VP.n19 0.189894
R583 VP.n21 VP.n20 0.189894
R584 VP.n21 VP.n10 0.189894
R585 VP.n26 VP.n10 0.189894
R586 VP.n27 VP.n26 0.189894
R587 VP.n28 VP.n27 0.189894
R588 VP.n28 VP.n8 0.189894
R589 VP.n32 VP.n8 0.189894
R590 VP.n34 VP.n33 0.189894
R591 VP.n34 VP.n6 0.189894
R592 VP.n38 VP.n6 0.189894
R593 VP.n39 VP.n38 0.189894
R594 VP.n39 VP.n4 0.189894
R595 VP.n43 VP.n4 0.189894
R596 VP.n44 VP.n43 0.189894
R597 VP.n45 VP.n44 0.189894
R598 VP.n45 VP.n2 0.189894
R599 VP.n50 VP.n2 0.189894
R600 VP.n51 VP.n50 0.189894
R601 VP.n52 VP.n51 0.189894
R602 VP.n52 VP.n0 0.189894
R603 VP.n56 VP.n0 0.189894
R604 VP VP.n56 0.0516364
R605 VDD1.n36 VDD1.n0 756.745
R606 VDD1.n79 VDD1.n43 756.745
R607 VDD1.n37 VDD1.n36 585
R608 VDD1.n35 VDD1.n2 585
R609 VDD1.n34 VDD1.n33 585
R610 VDD1.n5 VDD1.n3 585
R611 VDD1.n28 VDD1.n27 585
R612 VDD1.n26 VDD1.n25 585
R613 VDD1.n9 VDD1.n8 585
R614 VDD1.n20 VDD1.n19 585
R615 VDD1.n18 VDD1.n17 585
R616 VDD1.n13 VDD1.n12 585
R617 VDD1.n55 VDD1.n54 585
R618 VDD1.n60 VDD1.n59 585
R619 VDD1.n62 VDD1.n61 585
R620 VDD1.n51 VDD1.n50 585
R621 VDD1.n68 VDD1.n67 585
R622 VDD1.n70 VDD1.n69 585
R623 VDD1.n47 VDD1.n46 585
R624 VDD1.n77 VDD1.n76 585
R625 VDD1.n78 VDD1.n45 585
R626 VDD1.n80 VDD1.n79 585
R627 VDD1.n14 VDD1.t1 329.043
R628 VDD1.n56 VDD1.t5 329.043
R629 VDD1.n36 VDD1.n35 171.744
R630 VDD1.n35 VDD1.n34 171.744
R631 VDD1.n34 VDD1.n3 171.744
R632 VDD1.n27 VDD1.n3 171.744
R633 VDD1.n27 VDD1.n26 171.744
R634 VDD1.n26 VDD1.n8 171.744
R635 VDD1.n19 VDD1.n8 171.744
R636 VDD1.n19 VDD1.n18 171.744
R637 VDD1.n18 VDD1.n12 171.744
R638 VDD1.n60 VDD1.n54 171.744
R639 VDD1.n61 VDD1.n60 171.744
R640 VDD1.n61 VDD1.n50 171.744
R641 VDD1.n68 VDD1.n50 171.744
R642 VDD1.n69 VDD1.n68 171.744
R643 VDD1.n69 VDD1.n46 171.744
R644 VDD1.n77 VDD1.n46 171.744
R645 VDD1.n78 VDD1.n77 171.744
R646 VDD1.n79 VDD1.n78 171.744
R647 VDD1.t1 VDD1.n12 85.8723
R648 VDD1.t5 VDD1.n54 85.8723
R649 VDD1.n87 VDD1.n86 84.6958
R650 VDD1.n42 VDD1.n41 83.7168
R651 VDD1.n89 VDD1.n88 83.7166
R652 VDD1.n85 VDD1.n84 83.7166
R653 VDD1.n42 VDD1.n40 51.601
R654 VDD1.n85 VDD1.n83 51.601
R655 VDD1.n89 VDD1.n87 38.3328
R656 VDD1.n37 VDD1.n2 13.1884
R657 VDD1.n80 VDD1.n45 13.1884
R658 VDD1.n38 VDD1.n0 12.8005
R659 VDD1.n33 VDD1.n4 12.8005
R660 VDD1.n76 VDD1.n75 12.8005
R661 VDD1.n81 VDD1.n43 12.8005
R662 VDD1.n32 VDD1.n5 12.0247
R663 VDD1.n74 VDD1.n47 12.0247
R664 VDD1.n29 VDD1.n28 11.249
R665 VDD1.n71 VDD1.n70 11.249
R666 VDD1.n14 VDD1.n13 10.7238
R667 VDD1.n56 VDD1.n55 10.7238
R668 VDD1.n25 VDD1.n7 10.4732
R669 VDD1.n67 VDD1.n49 10.4732
R670 VDD1.n24 VDD1.n9 9.69747
R671 VDD1.n66 VDD1.n51 9.69747
R672 VDD1.n40 VDD1.n39 9.45567
R673 VDD1.n83 VDD1.n82 9.45567
R674 VDD1.n16 VDD1.n15 9.3005
R675 VDD1.n11 VDD1.n10 9.3005
R676 VDD1.n22 VDD1.n21 9.3005
R677 VDD1.n24 VDD1.n23 9.3005
R678 VDD1.n7 VDD1.n6 9.3005
R679 VDD1.n30 VDD1.n29 9.3005
R680 VDD1.n32 VDD1.n31 9.3005
R681 VDD1.n4 VDD1.n1 9.3005
R682 VDD1.n39 VDD1.n38 9.3005
R683 VDD1.n82 VDD1.n81 9.3005
R684 VDD1.n58 VDD1.n57 9.3005
R685 VDD1.n53 VDD1.n52 9.3005
R686 VDD1.n64 VDD1.n63 9.3005
R687 VDD1.n66 VDD1.n65 9.3005
R688 VDD1.n49 VDD1.n48 9.3005
R689 VDD1.n72 VDD1.n71 9.3005
R690 VDD1.n74 VDD1.n73 9.3005
R691 VDD1.n75 VDD1.n44 9.3005
R692 VDD1.n21 VDD1.n20 8.92171
R693 VDD1.n63 VDD1.n62 8.92171
R694 VDD1.n17 VDD1.n11 8.14595
R695 VDD1.n59 VDD1.n53 8.14595
R696 VDD1.n16 VDD1.n13 7.3702
R697 VDD1.n58 VDD1.n55 7.3702
R698 VDD1.n17 VDD1.n16 5.81868
R699 VDD1.n59 VDD1.n58 5.81868
R700 VDD1.n20 VDD1.n11 5.04292
R701 VDD1.n62 VDD1.n53 5.04292
R702 VDD1.n21 VDD1.n9 4.26717
R703 VDD1.n63 VDD1.n51 4.26717
R704 VDD1.n88 VDD1.t2 4.13074
R705 VDD1.n88 VDD1.t6 4.13074
R706 VDD1.n41 VDD1.t3 4.13074
R707 VDD1.n41 VDD1.t9 4.13074
R708 VDD1.n86 VDD1.t4 4.13074
R709 VDD1.n86 VDD1.t7 4.13074
R710 VDD1.n84 VDD1.t8 4.13074
R711 VDD1.n84 VDD1.t0 4.13074
R712 VDD1.n25 VDD1.n24 3.49141
R713 VDD1.n67 VDD1.n66 3.49141
R714 VDD1.n28 VDD1.n7 2.71565
R715 VDD1.n70 VDD1.n49 2.71565
R716 VDD1.n15 VDD1.n14 2.4129
R717 VDD1.n57 VDD1.n56 2.4129
R718 VDD1.n29 VDD1.n5 1.93989
R719 VDD1.n71 VDD1.n47 1.93989
R720 VDD1.n40 VDD1.n0 1.16414
R721 VDD1.n33 VDD1.n32 1.16414
R722 VDD1.n76 VDD1.n74 1.16414
R723 VDD1.n83 VDD1.n43 1.16414
R724 VDD1 VDD1.n89 0.976793
R725 VDD1 VDD1.n42 0.403517
R726 VDD1.n38 VDD1.n37 0.388379
R727 VDD1.n4 VDD1.n2 0.388379
R728 VDD1.n75 VDD1.n45 0.388379
R729 VDD1.n81 VDD1.n80 0.388379
R730 VDD1.n87 VDD1.n85 0.289982
R731 VDD1.n39 VDD1.n1 0.155672
R732 VDD1.n31 VDD1.n1 0.155672
R733 VDD1.n31 VDD1.n30 0.155672
R734 VDD1.n30 VDD1.n6 0.155672
R735 VDD1.n23 VDD1.n6 0.155672
R736 VDD1.n23 VDD1.n22 0.155672
R737 VDD1.n22 VDD1.n10 0.155672
R738 VDD1.n15 VDD1.n10 0.155672
R739 VDD1.n57 VDD1.n52 0.155672
R740 VDD1.n64 VDD1.n52 0.155672
R741 VDD1.n65 VDD1.n64 0.155672
R742 VDD1.n65 VDD1.n48 0.155672
R743 VDD1.n72 VDD1.n48 0.155672
R744 VDD1.n73 VDD1.n72 0.155672
R745 VDD1.n73 VDD1.n44 0.155672
R746 VDD1.n82 VDD1.n44 0.155672
R747 B.n309 B.n308 585
R748 B.n307 B.n96 585
R749 B.n306 B.n305 585
R750 B.n304 B.n97 585
R751 B.n303 B.n302 585
R752 B.n301 B.n98 585
R753 B.n300 B.n299 585
R754 B.n298 B.n99 585
R755 B.n297 B.n296 585
R756 B.n295 B.n100 585
R757 B.n294 B.n293 585
R758 B.n292 B.n101 585
R759 B.n291 B.n290 585
R760 B.n289 B.n102 585
R761 B.n288 B.n287 585
R762 B.n286 B.n103 585
R763 B.n285 B.n284 585
R764 B.n283 B.n104 585
R765 B.n282 B.n281 585
R766 B.n280 B.n105 585
R767 B.n279 B.n278 585
R768 B.n277 B.n106 585
R769 B.n276 B.n275 585
R770 B.n274 B.n107 585
R771 B.n273 B.n272 585
R772 B.n271 B.n108 585
R773 B.n270 B.n269 585
R774 B.n268 B.n109 585
R775 B.n267 B.n266 585
R776 B.n265 B.n110 585
R777 B.n264 B.n263 585
R778 B.n259 B.n111 585
R779 B.n258 B.n257 585
R780 B.n256 B.n112 585
R781 B.n255 B.n254 585
R782 B.n253 B.n113 585
R783 B.n252 B.n251 585
R784 B.n250 B.n114 585
R785 B.n249 B.n248 585
R786 B.n246 B.n115 585
R787 B.n245 B.n244 585
R788 B.n243 B.n118 585
R789 B.n242 B.n241 585
R790 B.n240 B.n119 585
R791 B.n239 B.n238 585
R792 B.n237 B.n120 585
R793 B.n236 B.n235 585
R794 B.n234 B.n121 585
R795 B.n233 B.n232 585
R796 B.n231 B.n122 585
R797 B.n230 B.n229 585
R798 B.n228 B.n123 585
R799 B.n227 B.n226 585
R800 B.n225 B.n124 585
R801 B.n224 B.n223 585
R802 B.n222 B.n125 585
R803 B.n221 B.n220 585
R804 B.n219 B.n126 585
R805 B.n218 B.n217 585
R806 B.n216 B.n127 585
R807 B.n215 B.n214 585
R808 B.n213 B.n128 585
R809 B.n212 B.n211 585
R810 B.n210 B.n129 585
R811 B.n209 B.n208 585
R812 B.n207 B.n130 585
R813 B.n206 B.n205 585
R814 B.n204 B.n131 585
R815 B.n203 B.n202 585
R816 B.n310 B.n95 585
R817 B.n312 B.n311 585
R818 B.n313 B.n94 585
R819 B.n315 B.n314 585
R820 B.n316 B.n93 585
R821 B.n318 B.n317 585
R822 B.n319 B.n92 585
R823 B.n321 B.n320 585
R824 B.n322 B.n91 585
R825 B.n324 B.n323 585
R826 B.n325 B.n90 585
R827 B.n327 B.n326 585
R828 B.n328 B.n89 585
R829 B.n330 B.n329 585
R830 B.n331 B.n88 585
R831 B.n333 B.n332 585
R832 B.n334 B.n87 585
R833 B.n336 B.n335 585
R834 B.n337 B.n86 585
R835 B.n339 B.n338 585
R836 B.n340 B.n85 585
R837 B.n342 B.n341 585
R838 B.n343 B.n84 585
R839 B.n345 B.n344 585
R840 B.n346 B.n83 585
R841 B.n348 B.n347 585
R842 B.n349 B.n82 585
R843 B.n351 B.n350 585
R844 B.n352 B.n81 585
R845 B.n354 B.n353 585
R846 B.n355 B.n80 585
R847 B.n357 B.n356 585
R848 B.n358 B.n79 585
R849 B.n360 B.n359 585
R850 B.n361 B.n78 585
R851 B.n363 B.n362 585
R852 B.n364 B.n77 585
R853 B.n366 B.n365 585
R854 B.n367 B.n76 585
R855 B.n369 B.n368 585
R856 B.n370 B.n75 585
R857 B.n372 B.n371 585
R858 B.n373 B.n74 585
R859 B.n375 B.n374 585
R860 B.n376 B.n73 585
R861 B.n378 B.n377 585
R862 B.n379 B.n72 585
R863 B.n381 B.n380 585
R864 B.n382 B.n71 585
R865 B.n384 B.n383 585
R866 B.n385 B.n70 585
R867 B.n387 B.n386 585
R868 B.n388 B.n69 585
R869 B.n390 B.n389 585
R870 B.n391 B.n68 585
R871 B.n393 B.n392 585
R872 B.n394 B.n67 585
R873 B.n396 B.n395 585
R874 B.n397 B.n66 585
R875 B.n399 B.n398 585
R876 B.n400 B.n65 585
R877 B.n402 B.n401 585
R878 B.n403 B.n64 585
R879 B.n405 B.n404 585
R880 B.n406 B.n63 585
R881 B.n408 B.n407 585
R882 B.n409 B.n62 585
R883 B.n411 B.n410 585
R884 B.n412 B.n61 585
R885 B.n414 B.n413 585
R886 B.n415 B.n60 585
R887 B.n417 B.n416 585
R888 B.n418 B.n59 585
R889 B.n420 B.n419 585
R890 B.n525 B.n20 585
R891 B.n524 B.n523 585
R892 B.n522 B.n21 585
R893 B.n521 B.n520 585
R894 B.n519 B.n22 585
R895 B.n518 B.n517 585
R896 B.n516 B.n23 585
R897 B.n515 B.n514 585
R898 B.n513 B.n24 585
R899 B.n512 B.n511 585
R900 B.n510 B.n25 585
R901 B.n509 B.n508 585
R902 B.n507 B.n26 585
R903 B.n506 B.n505 585
R904 B.n504 B.n27 585
R905 B.n503 B.n502 585
R906 B.n501 B.n28 585
R907 B.n500 B.n499 585
R908 B.n498 B.n29 585
R909 B.n497 B.n496 585
R910 B.n495 B.n30 585
R911 B.n494 B.n493 585
R912 B.n492 B.n31 585
R913 B.n491 B.n490 585
R914 B.n489 B.n32 585
R915 B.n488 B.n487 585
R916 B.n486 B.n33 585
R917 B.n485 B.n484 585
R918 B.n483 B.n34 585
R919 B.n482 B.n481 585
R920 B.n479 B.n35 585
R921 B.n478 B.n477 585
R922 B.n476 B.n38 585
R923 B.n475 B.n474 585
R924 B.n473 B.n39 585
R925 B.n472 B.n471 585
R926 B.n470 B.n40 585
R927 B.n469 B.n468 585
R928 B.n467 B.n41 585
R929 B.n465 B.n464 585
R930 B.n463 B.n44 585
R931 B.n462 B.n461 585
R932 B.n460 B.n45 585
R933 B.n459 B.n458 585
R934 B.n457 B.n46 585
R935 B.n456 B.n455 585
R936 B.n454 B.n47 585
R937 B.n453 B.n452 585
R938 B.n451 B.n48 585
R939 B.n450 B.n449 585
R940 B.n448 B.n49 585
R941 B.n447 B.n446 585
R942 B.n445 B.n50 585
R943 B.n444 B.n443 585
R944 B.n442 B.n51 585
R945 B.n441 B.n440 585
R946 B.n439 B.n52 585
R947 B.n438 B.n437 585
R948 B.n436 B.n53 585
R949 B.n435 B.n434 585
R950 B.n433 B.n54 585
R951 B.n432 B.n431 585
R952 B.n430 B.n55 585
R953 B.n429 B.n428 585
R954 B.n427 B.n56 585
R955 B.n426 B.n425 585
R956 B.n424 B.n57 585
R957 B.n423 B.n422 585
R958 B.n421 B.n58 585
R959 B.n527 B.n526 585
R960 B.n528 B.n19 585
R961 B.n530 B.n529 585
R962 B.n531 B.n18 585
R963 B.n533 B.n532 585
R964 B.n534 B.n17 585
R965 B.n536 B.n535 585
R966 B.n537 B.n16 585
R967 B.n539 B.n538 585
R968 B.n540 B.n15 585
R969 B.n542 B.n541 585
R970 B.n543 B.n14 585
R971 B.n545 B.n544 585
R972 B.n546 B.n13 585
R973 B.n548 B.n547 585
R974 B.n549 B.n12 585
R975 B.n551 B.n550 585
R976 B.n552 B.n11 585
R977 B.n554 B.n553 585
R978 B.n555 B.n10 585
R979 B.n557 B.n556 585
R980 B.n558 B.n9 585
R981 B.n560 B.n559 585
R982 B.n561 B.n8 585
R983 B.n563 B.n562 585
R984 B.n564 B.n7 585
R985 B.n566 B.n565 585
R986 B.n567 B.n6 585
R987 B.n569 B.n568 585
R988 B.n570 B.n5 585
R989 B.n572 B.n571 585
R990 B.n573 B.n4 585
R991 B.n575 B.n574 585
R992 B.n576 B.n3 585
R993 B.n578 B.n577 585
R994 B.n579 B.n0 585
R995 B.n2 B.n1 585
R996 B.n150 B.n149 585
R997 B.n152 B.n151 585
R998 B.n153 B.n148 585
R999 B.n155 B.n154 585
R1000 B.n156 B.n147 585
R1001 B.n158 B.n157 585
R1002 B.n159 B.n146 585
R1003 B.n161 B.n160 585
R1004 B.n162 B.n145 585
R1005 B.n164 B.n163 585
R1006 B.n165 B.n144 585
R1007 B.n167 B.n166 585
R1008 B.n168 B.n143 585
R1009 B.n170 B.n169 585
R1010 B.n171 B.n142 585
R1011 B.n173 B.n172 585
R1012 B.n174 B.n141 585
R1013 B.n176 B.n175 585
R1014 B.n177 B.n140 585
R1015 B.n179 B.n178 585
R1016 B.n180 B.n139 585
R1017 B.n182 B.n181 585
R1018 B.n183 B.n138 585
R1019 B.n185 B.n184 585
R1020 B.n186 B.n137 585
R1021 B.n188 B.n187 585
R1022 B.n189 B.n136 585
R1023 B.n191 B.n190 585
R1024 B.n192 B.n135 585
R1025 B.n194 B.n193 585
R1026 B.n195 B.n134 585
R1027 B.n197 B.n196 585
R1028 B.n198 B.n133 585
R1029 B.n200 B.n199 585
R1030 B.n201 B.n132 585
R1031 B.n202 B.n201 439.647
R1032 B.n308 B.n95 439.647
R1033 B.n421 B.n420 439.647
R1034 B.n526 B.n525 439.647
R1035 B.n260 B.t3 354.452
R1036 B.n42 B.t6 354.452
R1037 B.n116 B.t9 353.938
R1038 B.n36 B.t0 353.938
R1039 B.n260 B.t4 332.394
R1040 B.n42 B.t8 332.394
R1041 B.n116 B.t10 332.394
R1042 B.n36 B.t2 332.394
R1043 B.n261 B.t5 301.363
R1044 B.n43 B.t7 301.363
R1045 B.n117 B.t11 301.363
R1046 B.n37 B.t1 301.363
R1047 B.n581 B.n580 256.663
R1048 B.n580 B.n579 235.042
R1049 B.n580 B.n2 235.042
R1050 B.n202 B.n131 163.367
R1051 B.n206 B.n131 163.367
R1052 B.n207 B.n206 163.367
R1053 B.n208 B.n207 163.367
R1054 B.n208 B.n129 163.367
R1055 B.n212 B.n129 163.367
R1056 B.n213 B.n212 163.367
R1057 B.n214 B.n213 163.367
R1058 B.n214 B.n127 163.367
R1059 B.n218 B.n127 163.367
R1060 B.n219 B.n218 163.367
R1061 B.n220 B.n219 163.367
R1062 B.n220 B.n125 163.367
R1063 B.n224 B.n125 163.367
R1064 B.n225 B.n224 163.367
R1065 B.n226 B.n225 163.367
R1066 B.n226 B.n123 163.367
R1067 B.n230 B.n123 163.367
R1068 B.n231 B.n230 163.367
R1069 B.n232 B.n231 163.367
R1070 B.n232 B.n121 163.367
R1071 B.n236 B.n121 163.367
R1072 B.n237 B.n236 163.367
R1073 B.n238 B.n237 163.367
R1074 B.n238 B.n119 163.367
R1075 B.n242 B.n119 163.367
R1076 B.n243 B.n242 163.367
R1077 B.n244 B.n243 163.367
R1078 B.n244 B.n115 163.367
R1079 B.n249 B.n115 163.367
R1080 B.n250 B.n249 163.367
R1081 B.n251 B.n250 163.367
R1082 B.n251 B.n113 163.367
R1083 B.n255 B.n113 163.367
R1084 B.n256 B.n255 163.367
R1085 B.n257 B.n256 163.367
R1086 B.n257 B.n111 163.367
R1087 B.n264 B.n111 163.367
R1088 B.n265 B.n264 163.367
R1089 B.n266 B.n265 163.367
R1090 B.n266 B.n109 163.367
R1091 B.n270 B.n109 163.367
R1092 B.n271 B.n270 163.367
R1093 B.n272 B.n271 163.367
R1094 B.n272 B.n107 163.367
R1095 B.n276 B.n107 163.367
R1096 B.n277 B.n276 163.367
R1097 B.n278 B.n277 163.367
R1098 B.n278 B.n105 163.367
R1099 B.n282 B.n105 163.367
R1100 B.n283 B.n282 163.367
R1101 B.n284 B.n283 163.367
R1102 B.n284 B.n103 163.367
R1103 B.n288 B.n103 163.367
R1104 B.n289 B.n288 163.367
R1105 B.n290 B.n289 163.367
R1106 B.n290 B.n101 163.367
R1107 B.n294 B.n101 163.367
R1108 B.n295 B.n294 163.367
R1109 B.n296 B.n295 163.367
R1110 B.n296 B.n99 163.367
R1111 B.n300 B.n99 163.367
R1112 B.n301 B.n300 163.367
R1113 B.n302 B.n301 163.367
R1114 B.n302 B.n97 163.367
R1115 B.n306 B.n97 163.367
R1116 B.n307 B.n306 163.367
R1117 B.n308 B.n307 163.367
R1118 B.n420 B.n59 163.367
R1119 B.n416 B.n59 163.367
R1120 B.n416 B.n415 163.367
R1121 B.n415 B.n414 163.367
R1122 B.n414 B.n61 163.367
R1123 B.n410 B.n61 163.367
R1124 B.n410 B.n409 163.367
R1125 B.n409 B.n408 163.367
R1126 B.n408 B.n63 163.367
R1127 B.n404 B.n63 163.367
R1128 B.n404 B.n403 163.367
R1129 B.n403 B.n402 163.367
R1130 B.n402 B.n65 163.367
R1131 B.n398 B.n65 163.367
R1132 B.n398 B.n397 163.367
R1133 B.n397 B.n396 163.367
R1134 B.n396 B.n67 163.367
R1135 B.n392 B.n67 163.367
R1136 B.n392 B.n391 163.367
R1137 B.n391 B.n390 163.367
R1138 B.n390 B.n69 163.367
R1139 B.n386 B.n69 163.367
R1140 B.n386 B.n385 163.367
R1141 B.n385 B.n384 163.367
R1142 B.n384 B.n71 163.367
R1143 B.n380 B.n71 163.367
R1144 B.n380 B.n379 163.367
R1145 B.n379 B.n378 163.367
R1146 B.n378 B.n73 163.367
R1147 B.n374 B.n73 163.367
R1148 B.n374 B.n373 163.367
R1149 B.n373 B.n372 163.367
R1150 B.n372 B.n75 163.367
R1151 B.n368 B.n75 163.367
R1152 B.n368 B.n367 163.367
R1153 B.n367 B.n366 163.367
R1154 B.n366 B.n77 163.367
R1155 B.n362 B.n77 163.367
R1156 B.n362 B.n361 163.367
R1157 B.n361 B.n360 163.367
R1158 B.n360 B.n79 163.367
R1159 B.n356 B.n79 163.367
R1160 B.n356 B.n355 163.367
R1161 B.n355 B.n354 163.367
R1162 B.n354 B.n81 163.367
R1163 B.n350 B.n81 163.367
R1164 B.n350 B.n349 163.367
R1165 B.n349 B.n348 163.367
R1166 B.n348 B.n83 163.367
R1167 B.n344 B.n83 163.367
R1168 B.n344 B.n343 163.367
R1169 B.n343 B.n342 163.367
R1170 B.n342 B.n85 163.367
R1171 B.n338 B.n85 163.367
R1172 B.n338 B.n337 163.367
R1173 B.n337 B.n336 163.367
R1174 B.n336 B.n87 163.367
R1175 B.n332 B.n87 163.367
R1176 B.n332 B.n331 163.367
R1177 B.n331 B.n330 163.367
R1178 B.n330 B.n89 163.367
R1179 B.n326 B.n89 163.367
R1180 B.n326 B.n325 163.367
R1181 B.n325 B.n324 163.367
R1182 B.n324 B.n91 163.367
R1183 B.n320 B.n91 163.367
R1184 B.n320 B.n319 163.367
R1185 B.n319 B.n318 163.367
R1186 B.n318 B.n93 163.367
R1187 B.n314 B.n93 163.367
R1188 B.n314 B.n313 163.367
R1189 B.n313 B.n312 163.367
R1190 B.n312 B.n95 163.367
R1191 B.n525 B.n524 163.367
R1192 B.n524 B.n21 163.367
R1193 B.n520 B.n21 163.367
R1194 B.n520 B.n519 163.367
R1195 B.n519 B.n518 163.367
R1196 B.n518 B.n23 163.367
R1197 B.n514 B.n23 163.367
R1198 B.n514 B.n513 163.367
R1199 B.n513 B.n512 163.367
R1200 B.n512 B.n25 163.367
R1201 B.n508 B.n25 163.367
R1202 B.n508 B.n507 163.367
R1203 B.n507 B.n506 163.367
R1204 B.n506 B.n27 163.367
R1205 B.n502 B.n27 163.367
R1206 B.n502 B.n501 163.367
R1207 B.n501 B.n500 163.367
R1208 B.n500 B.n29 163.367
R1209 B.n496 B.n29 163.367
R1210 B.n496 B.n495 163.367
R1211 B.n495 B.n494 163.367
R1212 B.n494 B.n31 163.367
R1213 B.n490 B.n31 163.367
R1214 B.n490 B.n489 163.367
R1215 B.n489 B.n488 163.367
R1216 B.n488 B.n33 163.367
R1217 B.n484 B.n33 163.367
R1218 B.n484 B.n483 163.367
R1219 B.n483 B.n482 163.367
R1220 B.n482 B.n35 163.367
R1221 B.n477 B.n35 163.367
R1222 B.n477 B.n476 163.367
R1223 B.n476 B.n475 163.367
R1224 B.n475 B.n39 163.367
R1225 B.n471 B.n39 163.367
R1226 B.n471 B.n470 163.367
R1227 B.n470 B.n469 163.367
R1228 B.n469 B.n41 163.367
R1229 B.n464 B.n41 163.367
R1230 B.n464 B.n463 163.367
R1231 B.n463 B.n462 163.367
R1232 B.n462 B.n45 163.367
R1233 B.n458 B.n45 163.367
R1234 B.n458 B.n457 163.367
R1235 B.n457 B.n456 163.367
R1236 B.n456 B.n47 163.367
R1237 B.n452 B.n47 163.367
R1238 B.n452 B.n451 163.367
R1239 B.n451 B.n450 163.367
R1240 B.n450 B.n49 163.367
R1241 B.n446 B.n49 163.367
R1242 B.n446 B.n445 163.367
R1243 B.n445 B.n444 163.367
R1244 B.n444 B.n51 163.367
R1245 B.n440 B.n51 163.367
R1246 B.n440 B.n439 163.367
R1247 B.n439 B.n438 163.367
R1248 B.n438 B.n53 163.367
R1249 B.n434 B.n53 163.367
R1250 B.n434 B.n433 163.367
R1251 B.n433 B.n432 163.367
R1252 B.n432 B.n55 163.367
R1253 B.n428 B.n55 163.367
R1254 B.n428 B.n427 163.367
R1255 B.n427 B.n426 163.367
R1256 B.n426 B.n57 163.367
R1257 B.n422 B.n57 163.367
R1258 B.n422 B.n421 163.367
R1259 B.n526 B.n19 163.367
R1260 B.n530 B.n19 163.367
R1261 B.n531 B.n530 163.367
R1262 B.n532 B.n531 163.367
R1263 B.n532 B.n17 163.367
R1264 B.n536 B.n17 163.367
R1265 B.n537 B.n536 163.367
R1266 B.n538 B.n537 163.367
R1267 B.n538 B.n15 163.367
R1268 B.n542 B.n15 163.367
R1269 B.n543 B.n542 163.367
R1270 B.n544 B.n543 163.367
R1271 B.n544 B.n13 163.367
R1272 B.n548 B.n13 163.367
R1273 B.n549 B.n548 163.367
R1274 B.n550 B.n549 163.367
R1275 B.n550 B.n11 163.367
R1276 B.n554 B.n11 163.367
R1277 B.n555 B.n554 163.367
R1278 B.n556 B.n555 163.367
R1279 B.n556 B.n9 163.367
R1280 B.n560 B.n9 163.367
R1281 B.n561 B.n560 163.367
R1282 B.n562 B.n561 163.367
R1283 B.n562 B.n7 163.367
R1284 B.n566 B.n7 163.367
R1285 B.n567 B.n566 163.367
R1286 B.n568 B.n567 163.367
R1287 B.n568 B.n5 163.367
R1288 B.n572 B.n5 163.367
R1289 B.n573 B.n572 163.367
R1290 B.n574 B.n573 163.367
R1291 B.n574 B.n3 163.367
R1292 B.n578 B.n3 163.367
R1293 B.n579 B.n578 163.367
R1294 B.n149 B.n2 163.367
R1295 B.n152 B.n149 163.367
R1296 B.n153 B.n152 163.367
R1297 B.n154 B.n153 163.367
R1298 B.n154 B.n147 163.367
R1299 B.n158 B.n147 163.367
R1300 B.n159 B.n158 163.367
R1301 B.n160 B.n159 163.367
R1302 B.n160 B.n145 163.367
R1303 B.n164 B.n145 163.367
R1304 B.n165 B.n164 163.367
R1305 B.n166 B.n165 163.367
R1306 B.n166 B.n143 163.367
R1307 B.n170 B.n143 163.367
R1308 B.n171 B.n170 163.367
R1309 B.n172 B.n171 163.367
R1310 B.n172 B.n141 163.367
R1311 B.n176 B.n141 163.367
R1312 B.n177 B.n176 163.367
R1313 B.n178 B.n177 163.367
R1314 B.n178 B.n139 163.367
R1315 B.n182 B.n139 163.367
R1316 B.n183 B.n182 163.367
R1317 B.n184 B.n183 163.367
R1318 B.n184 B.n137 163.367
R1319 B.n188 B.n137 163.367
R1320 B.n189 B.n188 163.367
R1321 B.n190 B.n189 163.367
R1322 B.n190 B.n135 163.367
R1323 B.n194 B.n135 163.367
R1324 B.n195 B.n194 163.367
R1325 B.n196 B.n195 163.367
R1326 B.n196 B.n133 163.367
R1327 B.n200 B.n133 163.367
R1328 B.n201 B.n200 163.367
R1329 B.n247 B.n117 59.5399
R1330 B.n262 B.n261 59.5399
R1331 B.n466 B.n43 59.5399
R1332 B.n480 B.n37 59.5399
R1333 B.n117 B.n116 31.0308
R1334 B.n261 B.n260 31.0308
R1335 B.n43 B.n42 31.0308
R1336 B.n37 B.n36 31.0308
R1337 B.n310 B.n309 28.5664
R1338 B.n527 B.n20 28.5664
R1339 B.n419 B.n58 28.5664
R1340 B.n203 B.n132 28.5664
R1341 B B.n581 18.0485
R1342 B.n528 B.n527 10.6151
R1343 B.n529 B.n528 10.6151
R1344 B.n529 B.n18 10.6151
R1345 B.n533 B.n18 10.6151
R1346 B.n534 B.n533 10.6151
R1347 B.n535 B.n534 10.6151
R1348 B.n535 B.n16 10.6151
R1349 B.n539 B.n16 10.6151
R1350 B.n540 B.n539 10.6151
R1351 B.n541 B.n540 10.6151
R1352 B.n541 B.n14 10.6151
R1353 B.n545 B.n14 10.6151
R1354 B.n546 B.n545 10.6151
R1355 B.n547 B.n546 10.6151
R1356 B.n547 B.n12 10.6151
R1357 B.n551 B.n12 10.6151
R1358 B.n552 B.n551 10.6151
R1359 B.n553 B.n552 10.6151
R1360 B.n553 B.n10 10.6151
R1361 B.n557 B.n10 10.6151
R1362 B.n558 B.n557 10.6151
R1363 B.n559 B.n558 10.6151
R1364 B.n559 B.n8 10.6151
R1365 B.n563 B.n8 10.6151
R1366 B.n564 B.n563 10.6151
R1367 B.n565 B.n564 10.6151
R1368 B.n565 B.n6 10.6151
R1369 B.n569 B.n6 10.6151
R1370 B.n570 B.n569 10.6151
R1371 B.n571 B.n570 10.6151
R1372 B.n571 B.n4 10.6151
R1373 B.n575 B.n4 10.6151
R1374 B.n576 B.n575 10.6151
R1375 B.n577 B.n576 10.6151
R1376 B.n577 B.n0 10.6151
R1377 B.n523 B.n20 10.6151
R1378 B.n523 B.n522 10.6151
R1379 B.n522 B.n521 10.6151
R1380 B.n521 B.n22 10.6151
R1381 B.n517 B.n22 10.6151
R1382 B.n517 B.n516 10.6151
R1383 B.n516 B.n515 10.6151
R1384 B.n515 B.n24 10.6151
R1385 B.n511 B.n24 10.6151
R1386 B.n511 B.n510 10.6151
R1387 B.n510 B.n509 10.6151
R1388 B.n509 B.n26 10.6151
R1389 B.n505 B.n26 10.6151
R1390 B.n505 B.n504 10.6151
R1391 B.n504 B.n503 10.6151
R1392 B.n503 B.n28 10.6151
R1393 B.n499 B.n28 10.6151
R1394 B.n499 B.n498 10.6151
R1395 B.n498 B.n497 10.6151
R1396 B.n497 B.n30 10.6151
R1397 B.n493 B.n30 10.6151
R1398 B.n493 B.n492 10.6151
R1399 B.n492 B.n491 10.6151
R1400 B.n491 B.n32 10.6151
R1401 B.n487 B.n32 10.6151
R1402 B.n487 B.n486 10.6151
R1403 B.n486 B.n485 10.6151
R1404 B.n485 B.n34 10.6151
R1405 B.n481 B.n34 10.6151
R1406 B.n479 B.n478 10.6151
R1407 B.n478 B.n38 10.6151
R1408 B.n474 B.n38 10.6151
R1409 B.n474 B.n473 10.6151
R1410 B.n473 B.n472 10.6151
R1411 B.n472 B.n40 10.6151
R1412 B.n468 B.n40 10.6151
R1413 B.n468 B.n467 10.6151
R1414 B.n465 B.n44 10.6151
R1415 B.n461 B.n44 10.6151
R1416 B.n461 B.n460 10.6151
R1417 B.n460 B.n459 10.6151
R1418 B.n459 B.n46 10.6151
R1419 B.n455 B.n46 10.6151
R1420 B.n455 B.n454 10.6151
R1421 B.n454 B.n453 10.6151
R1422 B.n453 B.n48 10.6151
R1423 B.n449 B.n48 10.6151
R1424 B.n449 B.n448 10.6151
R1425 B.n448 B.n447 10.6151
R1426 B.n447 B.n50 10.6151
R1427 B.n443 B.n50 10.6151
R1428 B.n443 B.n442 10.6151
R1429 B.n442 B.n441 10.6151
R1430 B.n441 B.n52 10.6151
R1431 B.n437 B.n52 10.6151
R1432 B.n437 B.n436 10.6151
R1433 B.n436 B.n435 10.6151
R1434 B.n435 B.n54 10.6151
R1435 B.n431 B.n54 10.6151
R1436 B.n431 B.n430 10.6151
R1437 B.n430 B.n429 10.6151
R1438 B.n429 B.n56 10.6151
R1439 B.n425 B.n56 10.6151
R1440 B.n425 B.n424 10.6151
R1441 B.n424 B.n423 10.6151
R1442 B.n423 B.n58 10.6151
R1443 B.n419 B.n418 10.6151
R1444 B.n418 B.n417 10.6151
R1445 B.n417 B.n60 10.6151
R1446 B.n413 B.n60 10.6151
R1447 B.n413 B.n412 10.6151
R1448 B.n412 B.n411 10.6151
R1449 B.n411 B.n62 10.6151
R1450 B.n407 B.n62 10.6151
R1451 B.n407 B.n406 10.6151
R1452 B.n406 B.n405 10.6151
R1453 B.n405 B.n64 10.6151
R1454 B.n401 B.n64 10.6151
R1455 B.n401 B.n400 10.6151
R1456 B.n400 B.n399 10.6151
R1457 B.n399 B.n66 10.6151
R1458 B.n395 B.n66 10.6151
R1459 B.n395 B.n394 10.6151
R1460 B.n394 B.n393 10.6151
R1461 B.n393 B.n68 10.6151
R1462 B.n389 B.n68 10.6151
R1463 B.n389 B.n388 10.6151
R1464 B.n388 B.n387 10.6151
R1465 B.n387 B.n70 10.6151
R1466 B.n383 B.n70 10.6151
R1467 B.n383 B.n382 10.6151
R1468 B.n382 B.n381 10.6151
R1469 B.n381 B.n72 10.6151
R1470 B.n377 B.n72 10.6151
R1471 B.n377 B.n376 10.6151
R1472 B.n376 B.n375 10.6151
R1473 B.n375 B.n74 10.6151
R1474 B.n371 B.n74 10.6151
R1475 B.n371 B.n370 10.6151
R1476 B.n370 B.n369 10.6151
R1477 B.n369 B.n76 10.6151
R1478 B.n365 B.n76 10.6151
R1479 B.n365 B.n364 10.6151
R1480 B.n364 B.n363 10.6151
R1481 B.n363 B.n78 10.6151
R1482 B.n359 B.n78 10.6151
R1483 B.n359 B.n358 10.6151
R1484 B.n358 B.n357 10.6151
R1485 B.n357 B.n80 10.6151
R1486 B.n353 B.n80 10.6151
R1487 B.n353 B.n352 10.6151
R1488 B.n352 B.n351 10.6151
R1489 B.n351 B.n82 10.6151
R1490 B.n347 B.n82 10.6151
R1491 B.n347 B.n346 10.6151
R1492 B.n346 B.n345 10.6151
R1493 B.n345 B.n84 10.6151
R1494 B.n341 B.n84 10.6151
R1495 B.n341 B.n340 10.6151
R1496 B.n340 B.n339 10.6151
R1497 B.n339 B.n86 10.6151
R1498 B.n335 B.n86 10.6151
R1499 B.n335 B.n334 10.6151
R1500 B.n334 B.n333 10.6151
R1501 B.n333 B.n88 10.6151
R1502 B.n329 B.n88 10.6151
R1503 B.n329 B.n328 10.6151
R1504 B.n328 B.n327 10.6151
R1505 B.n327 B.n90 10.6151
R1506 B.n323 B.n90 10.6151
R1507 B.n323 B.n322 10.6151
R1508 B.n322 B.n321 10.6151
R1509 B.n321 B.n92 10.6151
R1510 B.n317 B.n92 10.6151
R1511 B.n317 B.n316 10.6151
R1512 B.n316 B.n315 10.6151
R1513 B.n315 B.n94 10.6151
R1514 B.n311 B.n94 10.6151
R1515 B.n311 B.n310 10.6151
R1516 B.n150 B.n1 10.6151
R1517 B.n151 B.n150 10.6151
R1518 B.n151 B.n148 10.6151
R1519 B.n155 B.n148 10.6151
R1520 B.n156 B.n155 10.6151
R1521 B.n157 B.n156 10.6151
R1522 B.n157 B.n146 10.6151
R1523 B.n161 B.n146 10.6151
R1524 B.n162 B.n161 10.6151
R1525 B.n163 B.n162 10.6151
R1526 B.n163 B.n144 10.6151
R1527 B.n167 B.n144 10.6151
R1528 B.n168 B.n167 10.6151
R1529 B.n169 B.n168 10.6151
R1530 B.n169 B.n142 10.6151
R1531 B.n173 B.n142 10.6151
R1532 B.n174 B.n173 10.6151
R1533 B.n175 B.n174 10.6151
R1534 B.n175 B.n140 10.6151
R1535 B.n179 B.n140 10.6151
R1536 B.n180 B.n179 10.6151
R1537 B.n181 B.n180 10.6151
R1538 B.n181 B.n138 10.6151
R1539 B.n185 B.n138 10.6151
R1540 B.n186 B.n185 10.6151
R1541 B.n187 B.n186 10.6151
R1542 B.n187 B.n136 10.6151
R1543 B.n191 B.n136 10.6151
R1544 B.n192 B.n191 10.6151
R1545 B.n193 B.n192 10.6151
R1546 B.n193 B.n134 10.6151
R1547 B.n197 B.n134 10.6151
R1548 B.n198 B.n197 10.6151
R1549 B.n199 B.n198 10.6151
R1550 B.n199 B.n132 10.6151
R1551 B.n204 B.n203 10.6151
R1552 B.n205 B.n204 10.6151
R1553 B.n205 B.n130 10.6151
R1554 B.n209 B.n130 10.6151
R1555 B.n210 B.n209 10.6151
R1556 B.n211 B.n210 10.6151
R1557 B.n211 B.n128 10.6151
R1558 B.n215 B.n128 10.6151
R1559 B.n216 B.n215 10.6151
R1560 B.n217 B.n216 10.6151
R1561 B.n217 B.n126 10.6151
R1562 B.n221 B.n126 10.6151
R1563 B.n222 B.n221 10.6151
R1564 B.n223 B.n222 10.6151
R1565 B.n223 B.n124 10.6151
R1566 B.n227 B.n124 10.6151
R1567 B.n228 B.n227 10.6151
R1568 B.n229 B.n228 10.6151
R1569 B.n229 B.n122 10.6151
R1570 B.n233 B.n122 10.6151
R1571 B.n234 B.n233 10.6151
R1572 B.n235 B.n234 10.6151
R1573 B.n235 B.n120 10.6151
R1574 B.n239 B.n120 10.6151
R1575 B.n240 B.n239 10.6151
R1576 B.n241 B.n240 10.6151
R1577 B.n241 B.n118 10.6151
R1578 B.n245 B.n118 10.6151
R1579 B.n246 B.n245 10.6151
R1580 B.n248 B.n114 10.6151
R1581 B.n252 B.n114 10.6151
R1582 B.n253 B.n252 10.6151
R1583 B.n254 B.n253 10.6151
R1584 B.n254 B.n112 10.6151
R1585 B.n258 B.n112 10.6151
R1586 B.n259 B.n258 10.6151
R1587 B.n263 B.n259 10.6151
R1588 B.n267 B.n110 10.6151
R1589 B.n268 B.n267 10.6151
R1590 B.n269 B.n268 10.6151
R1591 B.n269 B.n108 10.6151
R1592 B.n273 B.n108 10.6151
R1593 B.n274 B.n273 10.6151
R1594 B.n275 B.n274 10.6151
R1595 B.n275 B.n106 10.6151
R1596 B.n279 B.n106 10.6151
R1597 B.n280 B.n279 10.6151
R1598 B.n281 B.n280 10.6151
R1599 B.n281 B.n104 10.6151
R1600 B.n285 B.n104 10.6151
R1601 B.n286 B.n285 10.6151
R1602 B.n287 B.n286 10.6151
R1603 B.n287 B.n102 10.6151
R1604 B.n291 B.n102 10.6151
R1605 B.n292 B.n291 10.6151
R1606 B.n293 B.n292 10.6151
R1607 B.n293 B.n100 10.6151
R1608 B.n297 B.n100 10.6151
R1609 B.n298 B.n297 10.6151
R1610 B.n299 B.n298 10.6151
R1611 B.n299 B.n98 10.6151
R1612 B.n303 B.n98 10.6151
R1613 B.n304 B.n303 10.6151
R1614 B.n305 B.n304 10.6151
R1615 B.n305 B.n96 10.6151
R1616 B.n309 B.n96 10.6151
R1617 B.n581 B.n0 8.11757
R1618 B.n581 B.n1 8.11757
R1619 B.n480 B.n479 6.7127
R1620 B.n467 B.n466 6.7127
R1621 B.n248 B.n247 6.7127
R1622 B.n263 B.n262 6.7127
R1623 B.n481 B.n480 3.90294
R1624 B.n466 B.n465 3.90294
R1625 B.n247 B.n246 3.90294
R1626 B.n262 B.n110 3.90294
C0 VN w_n2890_n2544# 5.73596f
C1 VN VTAIL 6.14566f
C2 w_n2890_n2544# VDD1 1.9813f
C3 VDD1 VTAIL 8.57761f
C4 w_n2890_n2544# B 7.1638f
C5 VTAIL B 2.27829f
C6 VN VDD1 0.150348f
C7 VN B 0.894428f
C8 VP w_n2890_n2544# 6.10812f
C9 VP VTAIL 6.16f
C10 VDD1 B 1.63508f
C11 VN VP 5.67861f
C12 VP VDD1 6.15186f
C13 VP B 1.5129f
C14 VDD2 w_n2890_n2544# 2.05577f
C15 VDD2 VTAIL 8.619121f
C16 VN VDD2 5.89167f
C17 VDD2 VDD1 1.32416f
C18 VDD2 B 1.70122f
C19 VDD2 VP 0.41361f
C20 w_n2890_n2544# VTAIL 2.43899f
C21 VDD2 VSUBS 1.445874f
C22 VDD1 VSUBS 1.251509f
C23 VTAIL VSUBS 0.833277f
C24 VN VSUBS 5.41377f
C25 VP VSUBS 2.380649f
C26 B VSUBS 3.367971f
C27 w_n2890_n2544# VSUBS 91.2431f
C28 B.n0 VSUBS 0.006742f
C29 B.n1 VSUBS 0.006742f
C30 B.n2 VSUBS 0.009971f
C31 B.n3 VSUBS 0.007641f
C32 B.n4 VSUBS 0.007641f
C33 B.n5 VSUBS 0.007641f
C34 B.n6 VSUBS 0.007641f
C35 B.n7 VSUBS 0.007641f
C36 B.n8 VSUBS 0.007641f
C37 B.n9 VSUBS 0.007641f
C38 B.n10 VSUBS 0.007641f
C39 B.n11 VSUBS 0.007641f
C40 B.n12 VSUBS 0.007641f
C41 B.n13 VSUBS 0.007641f
C42 B.n14 VSUBS 0.007641f
C43 B.n15 VSUBS 0.007641f
C44 B.n16 VSUBS 0.007641f
C45 B.n17 VSUBS 0.007641f
C46 B.n18 VSUBS 0.007641f
C47 B.n19 VSUBS 0.007641f
C48 B.n20 VSUBS 0.016946f
C49 B.n21 VSUBS 0.007641f
C50 B.n22 VSUBS 0.007641f
C51 B.n23 VSUBS 0.007641f
C52 B.n24 VSUBS 0.007641f
C53 B.n25 VSUBS 0.007641f
C54 B.n26 VSUBS 0.007641f
C55 B.n27 VSUBS 0.007641f
C56 B.n28 VSUBS 0.007641f
C57 B.n29 VSUBS 0.007641f
C58 B.n30 VSUBS 0.007641f
C59 B.n31 VSUBS 0.007641f
C60 B.n32 VSUBS 0.007641f
C61 B.n33 VSUBS 0.007641f
C62 B.n34 VSUBS 0.007641f
C63 B.n35 VSUBS 0.007641f
C64 B.t1 VSUBS 0.135326f
C65 B.t2 VSUBS 0.153072f
C66 B.t0 VSUBS 0.484968f
C67 B.n36 VSUBS 0.255651f
C68 B.n37 VSUBS 0.200989f
C69 B.n38 VSUBS 0.007641f
C70 B.n39 VSUBS 0.007641f
C71 B.n40 VSUBS 0.007641f
C72 B.n41 VSUBS 0.007641f
C73 B.t7 VSUBS 0.135329f
C74 B.t8 VSUBS 0.153074f
C75 B.t6 VSUBS 0.485058f
C76 B.n42 VSUBS 0.255559f
C77 B.n43 VSUBS 0.200986f
C78 B.n44 VSUBS 0.007641f
C79 B.n45 VSUBS 0.007641f
C80 B.n46 VSUBS 0.007641f
C81 B.n47 VSUBS 0.007641f
C82 B.n48 VSUBS 0.007641f
C83 B.n49 VSUBS 0.007641f
C84 B.n50 VSUBS 0.007641f
C85 B.n51 VSUBS 0.007641f
C86 B.n52 VSUBS 0.007641f
C87 B.n53 VSUBS 0.007641f
C88 B.n54 VSUBS 0.007641f
C89 B.n55 VSUBS 0.007641f
C90 B.n56 VSUBS 0.007641f
C91 B.n57 VSUBS 0.007641f
C92 B.n58 VSUBS 0.016946f
C93 B.n59 VSUBS 0.007641f
C94 B.n60 VSUBS 0.007641f
C95 B.n61 VSUBS 0.007641f
C96 B.n62 VSUBS 0.007641f
C97 B.n63 VSUBS 0.007641f
C98 B.n64 VSUBS 0.007641f
C99 B.n65 VSUBS 0.007641f
C100 B.n66 VSUBS 0.007641f
C101 B.n67 VSUBS 0.007641f
C102 B.n68 VSUBS 0.007641f
C103 B.n69 VSUBS 0.007641f
C104 B.n70 VSUBS 0.007641f
C105 B.n71 VSUBS 0.007641f
C106 B.n72 VSUBS 0.007641f
C107 B.n73 VSUBS 0.007641f
C108 B.n74 VSUBS 0.007641f
C109 B.n75 VSUBS 0.007641f
C110 B.n76 VSUBS 0.007641f
C111 B.n77 VSUBS 0.007641f
C112 B.n78 VSUBS 0.007641f
C113 B.n79 VSUBS 0.007641f
C114 B.n80 VSUBS 0.007641f
C115 B.n81 VSUBS 0.007641f
C116 B.n82 VSUBS 0.007641f
C117 B.n83 VSUBS 0.007641f
C118 B.n84 VSUBS 0.007641f
C119 B.n85 VSUBS 0.007641f
C120 B.n86 VSUBS 0.007641f
C121 B.n87 VSUBS 0.007641f
C122 B.n88 VSUBS 0.007641f
C123 B.n89 VSUBS 0.007641f
C124 B.n90 VSUBS 0.007641f
C125 B.n91 VSUBS 0.007641f
C126 B.n92 VSUBS 0.007641f
C127 B.n93 VSUBS 0.007641f
C128 B.n94 VSUBS 0.007641f
C129 B.n95 VSUBS 0.015864f
C130 B.n96 VSUBS 0.007641f
C131 B.n97 VSUBS 0.007641f
C132 B.n98 VSUBS 0.007641f
C133 B.n99 VSUBS 0.007641f
C134 B.n100 VSUBS 0.007641f
C135 B.n101 VSUBS 0.007641f
C136 B.n102 VSUBS 0.007641f
C137 B.n103 VSUBS 0.007641f
C138 B.n104 VSUBS 0.007641f
C139 B.n105 VSUBS 0.007641f
C140 B.n106 VSUBS 0.007641f
C141 B.n107 VSUBS 0.007641f
C142 B.n108 VSUBS 0.007641f
C143 B.n109 VSUBS 0.007641f
C144 B.n110 VSUBS 0.005225f
C145 B.n111 VSUBS 0.007641f
C146 B.n112 VSUBS 0.007641f
C147 B.n113 VSUBS 0.007641f
C148 B.n114 VSUBS 0.007641f
C149 B.n115 VSUBS 0.007641f
C150 B.t11 VSUBS 0.135326f
C151 B.t10 VSUBS 0.153072f
C152 B.t9 VSUBS 0.484968f
C153 B.n116 VSUBS 0.255651f
C154 B.n117 VSUBS 0.200989f
C155 B.n118 VSUBS 0.007641f
C156 B.n119 VSUBS 0.007641f
C157 B.n120 VSUBS 0.007641f
C158 B.n121 VSUBS 0.007641f
C159 B.n122 VSUBS 0.007641f
C160 B.n123 VSUBS 0.007641f
C161 B.n124 VSUBS 0.007641f
C162 B.n125 VSUBS 0.007641f
C163 B.n126 VSUBS 0.007641f
C164 B.n127 VSUBS 0.007641f
C165 B.n128 VSUBS 0.007641f
C166 B.n129 VSUBS 0.007641f
C167 B.n130 VSUBS 0.007641f
C168 B.n131 VSUBS 0.007641f
C169 B.n132 VSUBS 0.015864f
C170 B.n133 VSUBS 0.007641f
C171 B.n134 VSUBS 0.007641f
C172 B.n135 VSUBS 0.007641f
C173 B.n136 VSUBS 0.007641f
C174 B.n137 VSUBS 0.007641f
C175 B.n138 VSUBS 0.007641f
C176 B.n139 VSUBS 0.007641f
C177 B.n140 VSUBS 0.007641f
C178 B.n141 VSUBS 0.007641f
C179 B.n142 VSUBS 0.007641f
C180 B.n143 VSUBS 0.007641f
C181 B.n144 VSUBS 0.007641f
C182 B.n145 VSUBS 0.007641f
C183 B.n146 VSUBS 0.007641f
C184 B.n147 VSUBS 0.007641f
C185 B.n148 VSUBS 0.007641f
C186 B.n149 VSUBS 0.007641f
C187 B.n150 VSUBS 0.007641f
C188 B.n151 VSUBS 0.007641f
C189 B.n152 VSUBS 0.007641f
C190 B.n153 VSUBS 0.007641f
C191 B.n154 VSUBS 0.007641f
C192 B.n155 VSUBS 0.007641f
C193 B.n156 VSUBS 0.007641f
C194 B.n157 VSUBS 0.007641f
C195 B.n158 VSUBS 0.007641f
C196 B.n159 VSUBS 0.007641f
C197 B.n160 VSUBS 0.007641f
C198 B.n161 VSUBS 0.007641f
C199 B.n162 VSUBS 0.007641f
C200 B.n163 VSUBS 0.007641f
C201 B.n164 VSUBS 0.007641f
C202 B.n165 VSUBS 0.007641f
C203 B.n166 VSUBS 0.007641f
C204 B.n167 VSUBS 0.007641f
C205 B.n168 VSUBS 0.007641f
C206 B.n169 VSUBS 0.007641f
C207 B.n170 VSUBS 0.007641f
C208 B.n171 VSUBS 0.007641f
C209 B.n172 VSUBS 0.007641f
C210 B.n173 VSUBS 0.007641f
C211 B.n174 VSUBS 0.007641f
C212 B.n175 VSUBS 0.007641f
C213 B.n176 VSUBS 0.007641f
C214 B.n177 VSUBS 0.007641f
C215 B.n178 VSUBS 0.007641f
C216 B.n179 VSUBS 0.007641f
C217 B.n180 VSUBS 0.007641f
C218 B.n181 VSUBS 0.007641f
C219 B.n182 VSUBS 0.007641f
C220 B.n183 VSUBS 0.007641f
C221 B.n184 VSUBS 0.007641f
C222 B.n185 VSUBS 0.007641f
C223 B.n186 VSUBS 0.007641f
C224 B.n187 VSUBS 0.007641f
C225 B.n188 VSUBS 0.007641f
C226 B.n189 VSUBS 0.007641f
C227 B.n190 VSUBS 0.007641f
C228 B.n191 VSUBS 0.007641f
C229 B.n192 VSUBS 0.007641f
C230 B.n193 VSUBS 0.007641f
C231 B.n194 VSUBS 0.007641f
C232 B.n195 VSUBS 0.007641f
C233 B.n196 VSUBS 0.007641f
C234 B.n197 VSUBS 0.007641f
C235 B.n198 VSUBS 0.007641f
C236 B.n199 VSUBS 0.007641f
C237 B.n200 VSUBS 0.007641f
C238 B.n201 VSUBS 0.015864f
C239 B.n202 VSUBS 0.016946f
C240 B.n203 VSUBS 0.016946f
C241 B.n204 VSUBS 0.007641f
C242 B.n205 VSUBS 0.007641f
C243 B.n206 VSUBS 0.007641f
C244 B.n207 VSUBS 0.007641f
C245 B.n208 VSUBS 0.007641f
C246 B.n209 VSUBS 0.007641f
C247 B.n210 VSUBS 0.007641f
C248 B.n211 VSUBS 0.007641f
C249 B.n212 VSUBS 0.007641f
C250 B.n213 VSUBS 0.007641f
C251 B.n214 VSUBS 0.007641f
C252 B.n215 VSUBS 0.007641f
C253 B.n216 VSUBS 0.007641f
C254 B.n217 VSUBS 0.007641f
C255 B.n218 VSUBS 0.007641f
C256 B.n219 VSUBS 0.007641f
C257 B.n220 VSUBS 0.007641f
C258 B.n221 VSUBS 0.007641f
C259 B.n222 VSUBS 0.007641f
C260 B.n223 VSUBS 0.007641f
C261 B.n224 VSUBS 0.007641f
C262 B.n225 VSUBS 0.007641f
C263 B.n226 VSUBS 0.007641f
C264 B.n227 VSUBS 0.007641f
C265 B.n228 VSUBS 0.007641f
C266 B.n229 VSUBS 0.007641f
C267 B.n230 VSUBS 0.007641f
C268 B.n231 VSUBS 0.007641f
C269 B.n232 VSUBS 0.007641f
C270 B.n233 VSUBS 0.007641f
C271 B.n234 VSUBS 0.007641f
C272 B.n235 VSUBS 0.007641f
C273 B.n236 VSUBS 0.007641f
C274 B.n237 VSUBS 0.007641f
C275 B.n238 VSUBS 0.007641f
C276 B.n239 VSUBS 0.007641f
C277 B.n240 VSUBS 0.007641f
C278 B.n241 VSUBS 0.007641f
C279 B.n242 VSUBS 0.007641f
C280 B.n243 VSUBS 0.007641f
C281 B.n244 VSUBS 0.007641f
C282 B.n245 VSUBS 0.007641f
C283 B.n246 VSUBS 0.005225f
C284 B.n247 VSUBS 0.017703f
C285 B.n248 VSUBS 0.006236f
C286 B.n249 VSUBS 0.007641f
C287 B.n250 VSUBS 0.007641f
C288 B.n251 VSUBS 0.007641f
C289 B.n252 VSUBS 0.007641f
C290 B.n253 VSUBS 0.007641f
C291 B.n254 VSUBS 0.007641f
C292 B.n255 VSUBS 0.007641f
C293 B.n256 VSUBS 0.007641f
C294 B.n257 VSUBS 0.007641f
C295 B.n258 VSUBS 0.007641f
C296 B.n259 VSUBS 0.007641f
C297 B.t5 VSUBS 0.135329f
C298 B.t4 VSUBS 0.153074f
C299 B.t3 VSUBS 0.485058f
C300 B.n260 VSUBS 0.255559f
C301 B.n261 VSUBS 0.200986f
C302 B.n262 VSUBS 0.017703f
C303 B.n263 VSUBS 0.006236f
C304 B.n264 VSUBS 0.007641f
C305 B.n265 VSUBS 0.007641f
C306 B.n266 VSUBS 0.007641f
C307 B.n267 VSUBS 0.007641f
C308 B.n268 VSUBS 0.007641f
C309 B.n269 VSUBS 0.007641f
C310 B.n270 VSUBS 0.007641f
C311 B.n271 VSUBS 0.007641f
C312 B.n272 VSUBS 0.007641f
C313 B.n273 VSUBS 0.007641f
C314 B.n274 VSUBS 0.007641f
C315 B.n275 VSUBS 0.007641f
C316 B.n276 VSUBS 0.007641f
C317 B.n277 VSUBS 0.007641f
C318 B.n278 VSUBS 0.007641f
C319 B.n279 VSUBS 0.007641f
C320 B.n280 VSUBS 0.007641f
C321 B.n281 VSUBS 0.007641f
C322 B.n282 VSUBS 0.007641f
C323 B.n283 VSUBS 0.007641f
C324 B.n284 VSUBS 0.007641f
C325 B.n285 VSUBS 0.007641f
C326 B.n286 VSUBS 0.007641f
C327 B.n287 VSUBS 0.007641f
C328 B.n288 VSUBS 0.007641f
C329 B.n289 VSUBS 0.007641f
C330 B.n290 VSUBS 0.007641f
C331 B.n291 VSUBS 0.007641f
C332 B.n292 VSUBS 0.007641f
C333 B.n293 VSUBS 0.007641f
C334 B.n294 VSUBS 0.007641f
C335 B.n295 VSUBS 0.007641f
C336 B.n296 VSUBS 0.007641f
C337 B.n297 VSUBS 0.007641f
C338 B.n298 VSUBS 0.007641f
C339 B.n299 VSUBS 0.007641f
C340 B.n300 VSUBS 0.007641f
C341 B.n301 VSUBS 0.007641f
C342 B.n302 VSUBS 0.007641f
C343 B.n303 VSUBS 0.007641f
C344 B.n304 VSUBS 0.007641f
C345 B.n305 VSUBS 0.007641f
C346 B.n306 VSUBS 0.007641f
C347 B.n307 VSUBS 0.007641f
C348 B.n308 VSUBS 0.016946f
C349 B.n309 VSUBS 0.015914f
C350 B.n310 VSUBS 0.016896f
C351 B.n311 VSUBS 0.007641f
C352 B.n312 VSUBS 0.007641f
C353 B.n313 VSUBS 0.007641f
C354 B.n314 VSUBS 0.007641f
C355 B.n315 VSUBS 0.007641f
C356 B.n316 VSUBS 0.007641f
C357 B.n317 VSUBS 0.007641f
C358 B.n318 VSUBS 0.007641f
C359 B.n319 VSUBS 0.007641f
C360 B.n320 VSUBS 0.007641f
C361 B.n321 VSUBS 0.007641f
C362 B.n322 VSUBS 0.007641f
C363 B.n323 VSUBS 0.007641f
C364 B.n324 VSUBS 0.007641f
C365 B.n325 VSUBS 0.007641f
C366 B.n326 VSUBS 0.007641f
C367 B.n327 VSUBS 0.007641f
C368 B.n328 VSUBS 0.007641f
C369 B.n329 VSUBS 0.007641f
C370 B.n330 VSUBS 0.007641f
C371 B.n331 VSUBS 0.007641f
C372 B.n332 VSUBS 0.007641f
C373 B.n333 VSUBS 0.007641f
C374 B.n334 VSUBS 0.007641f
C375 B.n335 VSUBS 0.007641f
C376 B.n336 VSUBS 0.007641f
C377 B.n337 VSUBS 0.007641f
C378 B.n338 VSUBS 0.007641f
C379 B.n339 VSUBS 0.007641f
C380 B.n340 VSUBS 0.007641f
C381 B.n341 VSUBS 0.007641f
C382 B.n342 VSUBS 0.007641f
C383 B.n343 VSUBS 0.007641f
C384 B.n344 VSUBS 0.007641f
C385 B.n345 VSUBS 0.007641f
C386 B.n346 VSUBS 0.007641f
C387 B.n347 VSUBS 0.007641f
C388 B.n348 VSUBS 0.007641f
C389 B.n349 VSUBS 0.007641f
C390 B.n350 VSUBS 0.007641f
C391 B.n351 VSUBS 0.007641f
C392 B.n352 VSUBS 0.007641f
C393 B.n353 VSUBS 0.007641f
C394 B.n354 VSUBS 0.007641f
C395 B.n355 VSUBS 0.007641f
C396 B.n356 VSUBS 0.007641f
C397 B.n357 VSUBS 0.007641f
C398 B.n358 VSUBS 0.007641f
C399 B.n359 VSUBS 0.007641f
C400 B.n360 VSUBS 0.007641f
C401 B.n361 VSUBS 0.007641f
C402 B.n362 VSUBS 0.007641f
C403 B.n363 VSUBS 0.007641f
C404 B.n364 VSUBS 0.007641f
C405 B.n365 VSUBS 0.007641f
C406 B.n366 VSUBS 0.007641f
C407 B.n367 VSUBS 0.007641f
C408 B.n368 VSUBS 0.007641f
C409 B.n369 VSUBS 0.007641f
C410 B.n370 VSUBS 0.007641f
C411 B.n371 VSUBS 0.007641f
C412 B.n372 VSUBS 0.007641f
C413 B.n373 VSUBS 0.007641f
C414 B.n374 VSUBS 0.007641f
C415 B.n375 VSUBS 0.007641f
C416 B.n376 VSUBS 0.007641f
C417 B.n377 VSUBS 0.007641f
C418 B.n378 VSUBS 0.007641f
C419 B.n379 VSUBS 0.007641f
C420 B.n380 VSUBS 0.007641f
C421 B.n381 VSUBS 0.007641f
C422 B.n382 VSUBS 0.007641f
C423 B.n383 VSUBS 0.007641f
C424 B.n384 VSUBS 0.007641f
C425 B.n385 VSUBS 0.007641f
C426 B.n386 VSUBS 0.007641f
C427 B.n387 VSUBS 0.007641f
C428 B.n388 VSUBS 0.007641f
C429 B.n389 VSUBS 0.007641f
C430 B.n390 VSUBS 0.007641f
C431 B.n391 VSUBS 0.007641f
C432 B.n392 VSUBS 0.007641f
C433 B.n393 VSUBS 0.007641f
C434 B.n394 VSUBS 0.007641f
C435 B.n395 VSUBS 0.007641f
C436 B.n396 VSUBS 0.007641f
C437 B.n397 VSUBS 0.007641f
C438 B.n398 VSUBS 0.007641f
C439 B.n399 VSUBS 0.007641f
C440 B.n400 VSUBS 0.007641f
C441 B.n401 VSUBS 0.007641f
C442 B.n402 VSUBS 0.007641f
C443 B.n403 VSUBS 0.007641f
C444 B.n404 VSUBS 0.007641f
C445 B.n405 VSUBS 0.007641f
C446 B.n406 VSUBS 0.007641f
C447 B.n407 VSUBS 0.007641f
C448 B.n408 VSUBS 0.007641f
C449 B.n409 VSUBS 0.007641f
C450 B.n410 VSUBS 0.007641f
C451 B.n411 VSUBS 0.007641f
C452 B.n412 VSUBS 0.007641f
C453 B.n413 VSUBS 0.007641f
C454 B.n414 VSUBS 0.007641f
C455 B.n415 VSUBS 0.007641f
C456 B.n416 VSUBS 0.007641f
C457 B.n417 VSUBS 0.007641f
C458 B.n418 VSUBS 0.007641f
C459 B.n419 VSUBS 0.015864f
C460 B.n420 VSUBS 0.015864f
C461 B.n421 VSUBS 0.016946f
C462 B.n422 VSUBS 0.007641f
C463 B.n423 VSUBS 0.007641f
C464 B.n424 VSUBS 0.007641f
C465 B.n425 VSUBS 0.007641f
C466 B.n426 VSUBS 0.007641f
C467 B.n427 VSUBS 0.007641f
C468 B.n428 VSUBS 0.007641f
C469 B.n429 VSUBS 0.007641f
C470 B.n430 VSUBS 0.007641f
C471 B.n431 VSUBS 0.007641f
C472 B.n432 VSUBS 0.007641f
C473 B.n433 VSUBS 0.007641f
C474 B.n434 VSUBS 0.007641f
C475 B.n435 VSUBS 0.007641f
C476 B.n436 VSUBS 0.007641f
C477 B.n437 VSUBS 0.007641f
C478 B.n438 VSUBS 0.007641f
C479 B.n439 VSUBS 0.007641f
C480 B.n440 VSUBS 0.007641f
C481 B.n441 VSUBS 0.007641f
C482 B.n442 VSUBS 0.007641f
C483 B.n443 VSUBS 0.007641f
C484 B.n444 VSUBS 0.007641f
C485 B.n445 VSUBS 0.007641f
C486 B.n446 VSUBS 0.007641f
C487 B.n447 VSUBS 0.007641f
C488 B.n448 VSUBS 0.007641f
C489 B.n449 VSUBS 0.007641f
C490 B.n450 VSUBS 0.007641f
C491 B.n451 VSUBS 0.007641f
C492 B.n452 VSUBS 0.007641f
C493 B.n453 VSUBS 0.007641f
C494 B.n454 VSUBS 0.007641f
C495 B.n455 VSUBS 0.007641f
C496 B.n456 VSUBS 0.007641f
C497 B.n457 VSUBS 0.007641f
C498 B.n458 VSUBS 0.007641f
C499 B.n459 VSUBS 0.007641f
C500 B.n460 VSUBS 0.007641f
C501 B.n461 VSUBS 0.007641f
C502 B.n462 VSUBS 0.007641f
C503 B.n463 VSUBS 0.007641f
C504 B.n464 VSUBS 0.007641f
C505 B.n465 VSUBS 0.005225f
C506 B.n466 VSUBS 0.017703f
C507 B.n467 VSUBS 0.006236f
C508 B.n468 VSUBS 0.007641f
C509 B.n469 VSUBS 0.007641f
C510 B.n470 VSUBS 0.007641f
C511 B.n471 VSUBS 0.007641f
C512 B.n472 VSUBS 0.007641f
C513 B.n473 VSUBS 0.007641f
C514 B.n474 VSUBS 0.007641f
C515 B.n475 VSUBS 0.007641f
C516 B.n476 VSUBS 0.007641f
C517 B.n477 VSUBS 0.007641f
C518 B.n478 VSUBS 0.007641f
C519 B.n479 VSUBS 0.006236f
C520 B.n480 VSUBS 0.017703f
C521 B.n481 VSUBS 0.005225f
C522 B.n482 VSUBS 0.007641f
C523 B.n483 VSUBS 0.007641f
C524 B.n484 VSUBS 0.007641f
C525 B.n485 VSUBS 0.007641f
C526 B.n486 VSUBS 0.007641f
C527 B.n487 VSUBS 0.007641f
C528 B.n488 VSUBS 0.007641f
C529 B.n489 VSUBS 0.007641f
C530 B.n490 VSUBS 0.007641f
C531 B.n491 VSUBS 0.007641f
C532 B.n492 VSUBS 0.007641f
C533 B.n493 VSUBS 0.007641f
C534 B.n494 VSUBS 0.007641f
C535 B.n495 VSUBS 0.007641f
C536 B.n496 VSUBS 0.007641f
C537 B.n497 VSUBS 0.007641f
C538 B.n498 VSUBS 0.007641f
C539 B.n499 VSUBS 0.007641f
C540 B.n500 VSUBS 0.007641f
C541 B.n501 VSUBS 0.007641f
C542 B.n502 VSUBS 0.007641f
C543 B.n503 VSUBS 0.007641f
C544 B.n504 VSUBS 0.007641f
C545 B.n505 VSUBS 0.007641f
C546 B.n506 VSUBS 0.007641f
C547 B.n507 VSUBS 0.007641f
C548 B.n508 VSUBS 0.007641f
C549 B.n509 VSUBS 0.007641f
C550 B.n510 VSUBS 0.007641f
C551 B.n511 VSUBS 0.007641f
C552 B.n512 VSUBS 0.007641f
C553 B.n513 VSUBS 0.007641f
C554 B.n514 VSUBS 0.007641f
C555 B.n515 VSUBS 0.007641f
C556 B.n516 VSUBS 0.007641f
C557 B.n517 VSUBS 0.007641f
C558 B.n518 VSUBS 0.007641f
C559 B.n519 VSUBS 0.007641f
C560 B.n520 VSUBS 0.007641f
C561 B.n521 VSUBS 0.007641f
C562 B.n522 VSUBS 0.007641f
C563 B.n523 VSUBS 0.007641f
C564 B.n524 VSUBS 0.007641f
C565 B.n525 VSUBS 0.016946f
C566 B.n526 VSUBS 0.015864f
C567 B.n527 VSUBS 0.015864f
C568 B.n528 VSUBS 0.007641f
C569 B.n529 VSUBS 0.007641f
C570 B.n530 VSUBS 0.007641f
C571 B.n531 VSUBS 0.007641f
C572 B.n532 VSUBS 0.007641f
C573 B.n533 VSUBS 0.007641f
C574 B.n534 VSUBS 0.007641f
C575 B.n535 VSUBS 0.007641f
C576 B.n536 VSUBS 0.007641f
C577 B.n537 VSUBS 0.007641f
C578 B.n538 VSUBS 0.007641f
C579 B.n539 VSUBS 0.007641f
C580 B.n540 VSUBS 0.007641f
C581 B.n541 VSUBS 0.007641f
C582 B.n542 VSUBS 0.007641f
C583 B.n543 VSUBS 0.007641f
C584 B.n544 VSUBS 0.007641f
C585 B.n545 VSUBS 0.007641f
C586 B.n546 VSUBS 0.007641f
C587 B.n547 VSUBS 0.007641f
C588 B.n548 VSUBS 0.007641f
C589 B.n549 VSUBS 0.007641f
C590 B.n550 VSUBS 0.007641f
C591 B.n551 VSUBS 0.007641f
C592 B.n552 VSUBS 0.007641f
C593 B.n553 VSUBS 0.007641f
C594 B.n554 VSUBS 0.007641f
C595 B.n555 VSUBS 0.007641f
C596 B.n556 VSUBS 0.007641f
C597 B.n557 VSUBS 0.007641f
C598 B.n558 VSUBS 0.007641f
C599 B.n559 VSUBS 0.007641f
C600 B.n560 VSUBS 0.007641f
C601 B.n561 VSUBS 0.007641f
C602 B.n562 VSUBS 0.007641f
C603 B.n563 VSUBS 0.007641f
C604 B.n564 VSUBS 0.007641f
C605 B.n565 VSUBS 0.007641f
C606 B.n566 VSUBS 0.007641f
C607 B.n567 VSUBS 0.007641f
C608 B.n568 VSUBS 0.007641f
C609 B.n569 VSUBS 0.007641f
C610 B.n570 VSUBS 0.007641f
C611 B.n571 VSUBS 0.007641f
C612 B.n572 VSUBS 0.007641f
C613 B.n573 VSUBS 0.007641f
C614 B.n574 VSUBS 0.007641f
C615 B.n575 VSUBS 0.007641f
C616 B.n576 VSUBS 0.007641f
C617 B.n577 VSUBS 0.007641f
C618 B.n578 VSUBS 0.007641f
C619 B.n579 VSUBS 0.009971f
C620 B.n580 VSUBS 0.010621f
C621 B.n581 VSUBS 0.021122f
C622 VDD1.n0 VSUBS 0.023757f
C623 VDD1.n1 VSUBS 0.023233f
C624 VDD1.n2 VSUBS 0.012852f
C625 VDD1.n3 VSUBS 0.029509f
C626 VDD1.n4 VSUBS 0.012485f
C627 VDD1.n5 VSUBS 0.013219f
C628 VDD1.n6 VSUBS 0.023233f
C629 VDD1.n7 VSUBS 0.012485f
C630 VDD1.n8 VSUBS 0.029509f
C631 VDD1.n9 VSUBS 0.013219f
C632 VDD1.n10 VSUBS 0.023233f
C633 VDD1.n11 VSUBS 0.012485f
C634 VDD1.n12 VSUBS 0.022132f
C635 VDD1.n13 VSUBS 0.022198f
C636 VDD1.t1 VSUBS 0.063354f
C637 VDD1.n14 VSUBS 0.139664f
C638 VDD1.n15 VSUBS 0.720932f
C639 VDD1.n16 VSUBS 0.012485f
C640 VDD1.n17 VSUBS 0.013219f
C641 VDD1.n18 VSUBS 0.029509f
C642 VDD1.n19 VSUBS 0.029509f
C643 VDD1.n20 VSUBS 0.013219f
C644 VDD1.n21 VSUBS 0.012485f
C645 VDD1.n22 VSUBS 0.023233f
C646 VDD1.n23 VSUBS 0.023233f
C647 VDD1.n24 VSUBS 0.012485f
C648 VDD1.n25 VSUBS 0.013219f
C649 VDD1.n26 VSUBS 0.029509f
C650 VDD1.n27 VSUBS 0.029509f
C651 VDD1.n28 VSUBS 0.013219f
C652 VDD1.n29 VSUBS 0.012485f
C653 VDD1.n30 VSUBS 0.023233f
C654 VDD1.n31 VSUBS 0.023233f
C655 VDD1.n32 VSUBS 0.012485f
C656 VDD1.n33 VSUBS 0.013219f
C657 VDD1.n34 VSUBS 0.029509f
C658 VDD1.n35 VSUBS 0.029509f
C659 VDD1.n36 VSUBS 0.065404f
C660 VDD1.n37 VSUBS 0.012852f
C661 VDD1.n38 VSUBS 0.012485f
C662 VDD1.n39 VSUBS 0.055925f
C663 VDD1.n40 VSUBS 0.052706f
C664 VDD1.t3 VSUBS 0.144491f
C665 VDD1.t9 VSUBS 0.144491f
C666 VDD1.n41 VSUBS 1.04111f
C667 VDD1.n42 VSUBS 0.671566f
C668 VDD1.n43 VSUBS 0.023757f
C669 VDD1.n44 VSUBS 0.023233f
C670 VDD1.n45 VSUBS 0.012852f
C671 VDD1.n46 VSUBS 0.029509f
C672 VDD1.n47 VSUBS 0.013219f
C673 VDD1.n48 VSUBS 0.023233f
C674 VDD1.n49 VSUBS 0.012485f
C675 VDD1.n50 VSUBS 0.029509f
C676 VDD1.n51 VSUBS 0.013219f
C677 VDD1.n52 VSUBS 0.023233f
C678 VDD1.n53 VSUBS 0.012485f
C679 VDD1.n54 VSUBS 0.022132f
C680 VDD1.n55 VSUBS 0.022198f
C681 VDD1.t5 VSUBS 0.063354f
C682 VDD1.n56 VSUBS 0.139664f
C683 VDD1.n57 VSUBS 0.720932f
C684 VDD1.n58 VSUBS 0.012485f
C685 VDD1.n59 VSUBS 0.013219f
C686 VDD1.n60 VSUBS 0.029509f
C687 VDD1.n61 VSUBS 0.029509f
C688 VDD1.n62 VSUBS 0.013219f
C689 VDD1.n63 VSUBS 0.012485f
C690 VDD1.n64 VSUBS 0.023233f
C691 VDD1.n65 VSUBS 0.023233f
C692 VDD1.n66 VSUBS 0.012485f
C693 VDD1.n67 VSUBS 0.013219f
C694 VDD1.n68 VSUBS 0.029509f
C695 VDD1.n69 VSUBS 0.029509f
C696 VDD1.n70 VSUBS 0.013219f
C697 VDD1.n71 VSUBS 0.012485f
C698 VDD1.n72 VSUBS 0.023233f
C699 VDD1.n73 VSUBS 0.023233f
C700 VDD1.n74 VSUBS 0.012485f
C701 VDD1.n75 VSUBS 0.012485f
C702 VDD1.n76 VSUBS 0.013219f
C703 VDD1.n77 VSUBS 0.029509f
C704 VDD1.n78 VSUBS 0.029509f
C705 VDD1.n79 VSUBS 0.065404f
C706 VDD1.n80 VSUBS 0.012852f
C707 VDD1.n81 VSUBS 0.012485f
C708 VDD1.n82 VSUBS 0.055925f
C709 VDD1.n83 VSUBS 0.052706f
C710 VDD1.t8 VSUBS 0.144491f
C711 VDD1.t0 VSUBS 0.144491f
C712 VDD1.n84 VSUBS 1.04111f
C713 VDD1.n85 VSUBS 0.664933f
C714 VDD1.t4 VSUBS 0.144491f
C715 VDD1.t7 VSUBS 0.144491f
C716 VDD1.n86 VSUBS 1.04781f
C717 VDD1.n87 VSUBS 2.10233f
C718 VDD1.t2 VSUBS 0.144491f
C719 VDD1.t6 VSUBS 0.144491f
C720 VDD1.n88 VSUBS 1.04111f
C721 VDD1.n89 VSUBS 2.34009f
C722 VP.n0 VSUBS 0.045989f
C723 VP.t2 VSUBS 1.23251f
C724 VP.n1 VSUBS 0.076693f
C725 VP.n2 VSUBS 0.045989f
C726 VP.t9 VSUBS 1.23251f
C727 VP.n3 VSUBS 0.51596f
C728 VP.n4 VSUBS 0.045989f
C729 VP.t1 VSUBS 1.23251f
C730 VP.n5 VSUBS 0.472135f
C731 VP.n6 VSUBS 0.045989f
C732 VP.t4 VSUBS 1.23251f
C733 VP.n7 VSUBS 0.549198f
C734 VP.n8 VSUBS 0.045989f
C735 VP.t3 VSUBS 1.23251f
C736 VP.n9 VSUBS 0.076693f
C737 VP.n10 VSUBS 0.045989f
C738 VP.t0 VSUBS 1.23251f
C739 VP.n11 VSUBS 0.51596f
C740 VP.n12 VSUBS 0.045989f
C741 VP.t6 VSUBS 1.23251f
C742 VP.n13 VSUBS 0.534288f
C743 VP.t8 VSUBS 1.32737f
C744 VP.n14 VSUBS 0.582212f
C745 VP.n15 VSUBS 0.239482f
C746 VP.n16 VSUBS 0.052374f
C747 VP.n17 VSUBS 0.061212f
C748 VP.n18 VSUBS 0.07421f
C749 VP.n19 VSUBS 0.045989f
C750 VP.n20 VSUBS 0.045989f
C751 VP.n21 VSUBS 0.045989f
C752 VP.n22 VSUBS 0.07421f
C753 VP.n23 VSUBS 0.061212f
C754 VP.t7 VSUBS 1.23251f
C755 VP.n24 VSUBS 0.472135f
C756 VP.n25 VSUBS 0.052374f
C757 VP.n26 VSUBS 0.045989f
C758 VP.n27 VSUBS 0.045989f
C759 VP.n28 VSUBS 0.045989f
C760 VP.n29 VSUBS 0.043616f
C761 VP.n30 VSUBS 0.067487f
C762 VP.n31 VSUBS 0.549198f
C763 VP.n32 VSUBS 1.95262f
C764 VP.n33 VSUBS 1.9914f
C765 VP.n34 VSUBS 0.045989f
C766 VP.n35 VSUBS 0.067487f
C767 VP.n36 VSUBS 0.043616f
C768 VP.n37 VSUBS 0.076693f
C769 VP.n38 VSUBS 0.045989f
C770 VP.n39 VSUBS 0.045989f
C771 VP.n40 VSUBS 0.052374f
C772 VP.n41 VSUBS 0.061212f
C773 VP.n42 VSUBS 0.07421f
C774 VP.n43 VSUBS 0.045989f
C775 VP.n44 VSUBS 0.045989f
C776 VP.n45 VSUBS 0.045989f
C777 VP.n46 VSUBS 0.07421f
C778 VP.n47 VSUBS 0.061212f
C779 VP.t5 VSUBS 1.23251f
C780 VP.n48 VSUBS 0.472135f
C781 VP.n49 VSUBS 0.052374f
C782 VP.n50 VSUBS 0.045989f
C783 VP.n51 VSUBS 0.045989f
C784 VP.n52 VSUBS 0.045989f
C785 VP.n53 VSUBS 0.043616f
C786 VP.n54 VSUBS 0.067487f
C787 VP.n55 VSUBS 0.549198f
C788 VP.n56 VSUBS 0.042583f
C789 VDD2.n0 VSUBS 0.026802f
C790 VDD2.n1 VSUBS 0.026211f
C791 VDD2.n2 VSUBS 0.014499f
C792 VDD2.n3 VSUBS 0.033291f
C793 VDD2.n4 VSUBS 0.014913f
C794 VDD2.n5 VSUBS 0.026211f
C795 VDD2.n6 VSUBS 0.014085f
C796 VDD2.n7 VSUBS 0.033291f
C797 VDD2.n8 VSUBS 0.014913f
C798 VDD2.n9 VSUBS 0.026211f
C799 VDD2.n10 VSUBS 0.014085f
C800 VDD2.n11 VSUBS 0.024968f
C801 VDD2.n12 VSUBS 0.025043f
C802 VDD2.t9 VSUBS 0.071473f
C803 VDD2.n13 VSUBS 0.157564f
C804 VDD2.n14 VSUBS 0.813329f
C805 VDD2.n15 VSUBS 0.014085f
C806 VDD2.n16 VSUBS 0.014913f
C807 VDD2.n17 VSUBS 0.033291f
C808 VDD2.n18 VSUBS 0.033291f
C809 VDD2.n19 VSUBS 0.014913f
C810 VDD2.n20 VSUBS 0.014085f
C811 VDD2.n21 VSUBS 0.026211f
C812 VDD2.n22 VSUBS 0.026211f
C813 VDD2.n23 VSUBS 0.014085f
C814 VDD2.n24 VSUBS 0.014913f
C815 VDD2.n25 VSUBS 0.033291f
C816 VDD2.n26 VSUBS 0.033291f
C817 VDD2.n27 VSUBS 0.014913f
C818 VDD2.n28 VSUBS 0.014085f
C819 VDD2.n29 VSUBS 0.026211f
C820 VDD2.n30 VSUBS 0.026211f
C821 VDD2.n31 VSUBS 0.014085f
C822 VDD2.n32 VSUBS 0.014085f
C823 VDD2.n33 VSUBS 0.014913f
C824 VDD2.n34 VSUBS 0.033291f
C825 VDD2.n35 VSUBS 0.033291f
C826 VDD2.n36 VSUBS 0.073787f
C827 VDD2.n37 VSUBS 0.014499f
C828 VDD2.n38 VSUBS 0.014085f
C829 VDD2.n39 VSUBS 0.063092f
C830 VDD2.n40 VSUBS 0.059461f
C831 VDD2.t3 VSUBS 0.163009f
C832 VDD2.t0 VSUBS 0.163009f
C833 VDD2.n41 VSUBS 1.17454f
C834 VDD2.n42 VSUBS 0.750152f
C835 VDD2.t8 VSUBS 0.163009f
C836 VDD2.t4 VSUBS 0.163009f
C837 VDD2.n43 VSUBS 1.1821f
C838 VDD2.n44 VSUBS 2.27896f
C839 VDD2.n45 VSUBS 0.026802f
C840 VDD2.n46 VSUBS 0.026211f
C841 VDD2.n47 VSUBS 0.014499f
C842 VDD2.n48 VSUBS 0.033291f
C843 VDD2.n49 VSUBS 0.014085f
C844 VDD2.n50 VSUBS 0.014913f
C845 VDD2.n51 VSUBS 0.026211f
C846 VDD2.n52 VSUBS 0.014085f
C847 VDD2.n53 VSUBS 0.033291f
C848 VDD2.n54 VSUBS 0.014913f
C849 VDD2.n55 VSUBS 0.026211f
C850 VDD2.n56 VSUBS 0.014085f
C851 VDD2.n57 VSUBS 0.024968f
C852 VDD2.n58 VSUBS 0.025043f
C853 VDD2.t1 VSUBS 0.071473f
C854 VDD2.n59 VSUBS 0.157564f
C855 VDD2.n60 VSUBS 0.813329f
C856 VDD2.n61 VSUBS 0.014085f
C857 VDD2.n62 VSUBS 0.014913f
C858 VDD2.n63 VSUBS 0.033291f
C859 VDD2.n64 VSUBS 0.033291f
C860 VDD2.n65 VSUBS 0.014913f
C861 VDD2.n66 VSUBS 0.014085f
C862 VDD2.n67 VSUBS 0.026211f
C863 VDD2.n68 VSUBS 0.026211f
C864 VDD2.n69 VSUBS 0.014085f
C865 VDD2.n70 VSUBS 0.014913f
C866 VDD2.n71 VSUBS 0.033291f
C867 VDD2.n72 VSUBS 0.033291f
C868 VDD2.n73 VSUBS 0.014913f
C869 VDD2.n74 VSUBS 0.014085f
C870 VDD2.n75 VSUBS 0.026211f
C871 VDD2.n76 VSUBS 0.026211f
C872 VDD2.n77 VSUBS 0.014085f
C873 VDD2.n78 VSUBS 0.014913f
C874 VDD2.n79 VSUBS 0.033291f
C875 VDD2.n80 VSUBS 0.033291f
C876 VDD2.n81 VSUBS 0.073787f
C877 VDD2.n82 VSUBS 0.014499f
C878 VDD2.n83 VSUBS 0.014085f
C879 VDD2.n84 VSUBS 0.063092f
C880 VDD2.n85 VSUBS 0.054959f
C881 VDD2.n86 VSUBS 2.15169f
C882 VDD2.t6 VSUBS 0.163009f
C883 VDD2.t5 VSUBS 0.163009f
C884 VDD2.n87 VSUBS 1.17455f
C885 VDD2.n88 VSUBS 0.593738f
C886 VDD2.t2 VSUBS 0.163009f
C887 VDD2.t7 VSUBS 0.163009f
C888 VDD2.n89 VSUBS 1.18207f
C889 VTAIL.t18 VSUBS 0.185548f
C890 VTAIL.t10 VSUBS 0.185548f
C891 VTAIL.n0 VSUBS 1.21284f
C892 VTAIL.n1 VSUBS 0.804559f
C893 VTAIL.n2 VSUBS 0.030508f
C894 VTAIL.n3 VSUBS 0.029835f
C895 VTAIL.n4 VSUBS 0.016504f
C896 VTAIL.n5 VSUBS 0.037894f
C897 VTAIL.n6 VSUBS 0.016975f
C898 VTAIL.n7 VSUBS 0.029835f
C899 VTAIL.n8 VSUBS 0.016032f
C900 VTAIL.n9 VSUBS 0.037894f
C901 VTAIL.n10 VSUBS 0.016975f
C902 VTAIL.n11 VSUBS 0.029835f
C903 VTAIL.n12 VSUBS 0.016032f
C904 VTAIL.n13 VSUBS 0.028421f
C905 VTAIL.n14 VSUBS 0.028506f
C906 VTAIL.t2 VSUBS 0.081356f
C907 VTAIL.n15 VSUBS 0.17935f
C908 VTAIL.n16 VSUBS 0.925787f
C909 VTAIL.n17 VSUBS 0.016032f
C910 VTAIL.n18 VSUBS 0.016975f
C911 VTAIL.n19 VSUBS 0.037894f
C912 VTAIL.n20 VSUBS 0.037894f
C913 VTAIL.n21 VSUBS 0.016975f
C914 VTAIL.n22 VSUBS 0.016032f
C915 VTAIL.n23 VSUBS 0.029835f
C916 VTAIL.n24 VSUBS 0.029835f
C917 VTAIL.n25 VSUBS 0.016032f
C918 VTAIL.n26 VSUBS 0.016975f
C919 VTAIL.n27 VSUBS 0.037894f
C920 VTAIL.n28 VSUBS 0.037894f
C921 VTAIL.n29 VSUBS 0.016975f
C922 VTAIL.n30 VSUBS 0.016032f
C923 VTAIL.n31 VSUBS 0.029835f
C924 VTAIL.n32 VSUBS 0.029835f
C925 VTAIL.n33 VSUBS 0.016032f
C926 VTAIL.n34 VSUBS 0.016032f
C927 VTAIL.n35 VSUBS 0.016975f
C928 VTAIL.n36 VSUBS 0.037894f
C929 VTAIL.n37 VSUBS 0.037894f
C930 VTAIL.n38 VSUBS 0.083989f
C931 VTAIL.n39 VSUBS 0.016504f
C932 VTAIL.n40 VSUBS 0.016032f
C933 VTAIL.n41 VSUBS 0.071816f
C934 VTAIL.n42 VSUBS 0.041979f
C935 VTAIL.n43 VSUBS 0.271162f
C936 VTAIL.t0 VSUBS 0.185548f
C937 VTAIL.t1 VSUBS 0.185548f
C938 VTAIL.n44 VSUBS 1.21284f
C939 VTAIL.n45 VSUBS 0.853249f
C940 VTAIL.t5 VSUBS 0.185548f
C941 VTAIL.t8 VSUBS 0.185548f
C942 VTAIL.n46 VSUBS 1.21284f
C943 VTAIL.n47 VSUBS 2.04418f
C944 VTAIL.t14 VSUBS 0.185548f
C945 VTAIL.t16 VSUBS 0.185548f
C946 VTAIL.n48 VSUBS 1.21285f
C947 VTAIL.n49 VSUBS 2.04418f
C948 VTAIL.t11 VSUBS 0.185548f
C949 VTAIL.t17 VSUBS 0.185548f
C950 VTAIL.n50 VSUBS 1.21285f
C951 VTAIL.n51 VSUBS 0.85324f
C952 VTAIL.n52 VSUBS 0.030508f
C953 VTAIL.n53 VSUBS 0.029835f
C954 VTAIL.n54 VSUBS 0.016504f
C955 VTAIL.n55 VSUBS 0.037894f
C956 VTAIL.n56 VSUBS 0.016032f
C957 VTAIL.n57 VSUBS 0.016975f
C958 VTAIL.n58 VSUBS 0.029835f
C959 VTAIL.n59 VSUBS 0.016032f
C960 VTAIL.n60 VSUBS 0.037894f
C961 VTAIL.n61 VSUBS 0.016975f
C962 VTAIL.n62 VSUBS 0.029835f
C963 VTAIL.n63 VSUBS 0.016032f
C964 VTAIL.n64 VSUBS 0.028421f
C965 VTAIL.n65 VSUBS 0.028506f
C966 VTAIL.t15 VSUBS 0.081356f
C967 VTAIL.n66 VSUBS 0.17935f
C968 VTAIL.n67 VSUBS 0.925787f
C969 VTAIL.n68 VSUBS 0.016032f
C970 VTAIL.n69 VSUBS 0.016975f
C971 VTAIL.n70 VSUBS 0.037894f
C972 VTAIL.n71 VSUBS 0.037894f
C973 VTAIL.n72 VSUBS 0.016975f
C974 VTAIL.n73 VSUBS 0.016032f
C975 VTAIL.n74 VSUBS 0.029835f
C976 VTAIL.n75 VSUBS 0.029835f
C977 VTAIL.n76 VSUBS 0.016032f
C978 VTAIL.n77 VSUBS 0.016975f
C979 VTAIL.n78 VSUBS 0.037894f
C980 VTAIL.n79 VSUBS 0.037894f
C981 VTAIL.n80 VSUBS 0.016975f
C982 VTAIL.n81 VSUBS 0.016032f
C983 VTAIL.n82 VSUBS 0.029835f
C984 VTAIL.n83 VSUBS 0.029835f
C985 VTAIL.n84 VSUBS 0.016032f
C986 VTAIL.n85 VSUBS 0.016975f
C987 VTAIL.n86 VSUBS 0.037894f
C988 VTAIL.n87 VSUBS 0.037894f
C989 VTAIL.n88 VSUBS 0.083989f
C990 VTAIL.n89 VSUBS 0.016504f
C991 VTAIL.n90 VSUBS 0.016032f
C992 VTAIL.n91 VSUBS 0.071816f
C993 VTAIL.n92 VSUBS 0.041979f
C994 VTAIL.n93 VSUBS 0.271162f
C995 VTAIL.t4 VSUBS 0.185548f
C996 VTAIL.t6 VSUBS 0.185548f
C997 VTAIL.n94 VSUBS 1.21285f
C998 VTAIL.n95 VSUBS 0.832107f
C999 VTAIL.t7 VSUBS 0.185548f
C1000 VTAIL.t3 VSUBS 0.185548f
C1001 VTAIL.n96 VSUBS 1.21285f
C1002 VTAIL.n97 VSUBS 0.85324f
C1003 VTAIL.n98 VSUBS 0.030508f
C1004 VTAIL.n99 VSUBS 0.029835f
C1005 VTAIL.n100 VSUBS 0.016504f
C1006 VTAIL.n101 VSUBS 0.037894f
C1007 VTAIL.n102 VSUBS 0.016032f
C1008 VTAIL.n103 VSUBS 0.016975f
C1009 VTAIL.n104 VSUBS 0.029835f
C1010 VTAIL.n105 VSUBS 0.016032f
C1011 VTAIL.n106 VSUBS 0.037894f
C1012 VTAIL.n107 VSUBS 0.016975f
C1013 VTAIL.n108 VSUBS 0.029835f
C1014 VTAIL.n109 VSUBS 0.016032f
C1015 VTAIL.n110 VSUBS 0.028421f
C1016 VTAIL.n111 VSUBS 0.028506f
C1017 VTAIL.t9 VSUBS 0.081356f
C1018 VTAIL.n112 VSUBS 0.17935f
C1019 VTAIL.n113 VSUBS 0.925787f
C1020 VTAIL.n114 VSUBS 0.016032f
C1021 VTAIL.n115 VSUBS 0.016975f
C1022 VTAIL.n116 VSUBS 0.037894f
C1023 VTAIL.n117 VSUBS 0.037894f
C1024 VTAIL.n118 VSUBS 0.016975f
C1025 VTAIL.n119 VSUBS 0.016032f
C1026 VTAIL.n120 VSUBS 0.029835f
C1027 VTAIL.n121 VSUBS 0.029835f
C1028 VTAIL.n122 VSUBS 0.016032f
C1029 VTAIL.n123 VSUBS 0.016975f
C1030 VTAIL.n124 VSUBS 0.037894f
C1031 VTAIL.n125 VSUBS 0.037894f
C1032 VTAIL.n126 VSUBS 0.016975f
C1033 VTAIL.n127 VSUBS 0.016032f
C1034 VTAIL.n128 VSUBS 0.029835f
C1035 VTAIL.n129 VSUBS 0.029835f
C1036 VTAIL.n130 VSUBS 0.016032f
C1037 VTAIL.n131 VSUBS 0.016975f
C1038 VTAIL.n132 VSUBS 0.037894f
C1039 VTAIL.n133 VSUBS 0.037894f
C1040 VTAIL.n134 VSUBS 0.083989f
C1041 VTAIL.n135 VSUBS 0.016504f
C1042 VTAIL.n136 VSUBS 0.016032f
C1043 VTAIL.n137 VSUBS 0.071816f
C1044 VTAIL.n138 VSUBS 0.041979f
C1045 VTAIL.n139 VSUBS 1.35063f
C1046 VTAIL.n140 VSUBS 0.030508f
C1047 VTAIL.n141 VSUBS 0.029835f
C1048 VTAIL.n142 VSUBS 0.016504f
C1049 VTAIL.n143 VSUBS 0.037894f
C1050 VTAIL.n144 VSUBS 0.016975f
C1051 VTAIL.n145 VSUBS 0.029835f
C1052 VTAIL.n146 VSUBS 0.016032f
C1053 VTAIL.n147 VSUBS 0.037894f
C1054 VTAIL.n148 VSUBS 0.016975f
C1055 VTAIL.n149 VSUBS 0.029835f
C1056 VTAIL.n150 VSUBS 0.016032f
C1057 VTAIL.n151 VSUBS 0.028421f
C1058 VTAIL.n152 VSUBS 0.028506f
C1059 VTAIL.t12 VSUBS 0.081356f
C1060 VTAIL.n153 VSUBS 0.17935f
C1061 VTAIL.n154 VSUBS 0.925787f
C1062 VTAIL.n155 VSUBS 0.016032f
C1063 VTAIL.n156 VSUBS 0.016975f
C1064 VTAIL.n157 VSUBS 0.037894f
C1065 VTAIL.n158 VSUBS 0.037894f
C1066 VTAIL.n159 VSUBS 0.016975f
C1067 VTAIL.n160 VSUBS 0.016032f
C1068 VTAIL.n161 VSUBS 0.029835f
C1069 VTAIL.n162 VSUBS 0.029835f
C1070 VTAIL.n163 VSUBS 0.016032f
C1071 VTAIL.n164 VSUBS 0.016975f
C1072 VTAIL.n165 VSUBS 0.037894f
C1073 VTAIL.n166 VSUBS 0.037894f
C1074 VTAIL.n167 VSUBS 0.016975f
C1075 VTAIL.n168 VSUBS 0.016032f
C1076 VTAIL.n169 VSUBS 0.029835f
C1077 VTAIL.n170 VSUBS 0.029835f
C1078 VTAIL.n171 VSUBS 0.016032f
C1079 VTAIL.n172 VSUBS 0.016032f
C1080 VTAIL.n173 VSUBS 0.016975f
C1081 VTAIL.n174 VSUBS 0.037894f
C1082 VTAIL.n175 VSUBS 0.037894f
C1083 VTAIL.n176 VSUBS 0.083989f
C1084 VTAIL.n177 VSUBS 0.016504f
C1085 VTAIL.n178 VSUBS 0.016032f
C1086 VTAIL.n179 VSUBS 0.071816f
C1087 VTAIL.n180 VSUBS 0.041979f
C1088 VTAIL.n181 VSUBS 1.35063f
C1089 VTAIL.t13 VSUBS 0.185548f
C1090 VTAIL.t19 VSUBS 0.185548f
C1091 VTAIL.n182 VSUBS 1.21284f
C1092 VTAIL.n183 VSUBS 0.748204f
C1093 VN.n0 VSUBS 0.04435f
C1094 VN.t5 VSUBS 1.1886f
C1095 VN.n1 VSUBS 0.07396f
C1096 VN.n2 VSUBS 0.04435f
C1097 VN.t9 VSUBS 1.1886f
C1098 VN.n3 VSUBS 0.497574f
C1099 VN.n4 VSUBS 0.04435f
C1100 VN.t6 VSUBS 1.1886f
C1101 VN.n5 VSUBS 0.515249f
C1102 VN.t0 VSUBS 1.28007f
C1103 VN.n6 VSUBS 0.561465f
C1104 VN.n7 VSUBS 0.230949f
C1105 VN.n8 VSUBS 0.050508f
C1106 VN.n9 VSUBS 0.059031f
C1107 VN.n10 VSUBS 0.071565f
C1108 VN.n11 VSUBS 0.04435f
C1109 VN.n12 VSUBS 0.04435f
C1110 VN.n13 VSUBS 0.04435f
C1111 VN.n14 VSUBS 0.071565f
C1112 VN.n15 VSUBS 0.059031f
C1113 VN.t1 VSUBS 1.1886f
C1114 VN.n16 VSUBS 0.455311f
C1115 VN.n17 VSUBS 0.050508f
C1116 VN.n18 VSUBS 0.04435f
C1117 VN.n19 VSUBS 0.04435f
C1118 VN.n20 VSUBS 0.04435f
C1119 VN.n21 VSUBS 0.042062f
C1120 VN.n22 VSUBS 0.065082f
C1121 VN.n23 VSUBS 0.529628f
C1122 VN.n24 VSUBS 0.041065f
C1123 VN.n25 VSUBS 0.04435f
C1124 VN.t8 VSUBS 1.1886f
C1125 VN.n26 VSUBS 0.07396f
C1126 VN.n27 VSUBS 0.04435f
C1127 VN.t3 VSUBS 1.1886f
C1128 VN.n28 VSUBS 0.455311f
C1129 VN.t4 VSUBS 1.1886f
C1130 VN.n29 VSUBS 0.497574f
C1131 VN.n30 VSUBS 0.04435f
C1132 VN.t7 VSUBS 1.1886f
C1133 VN.n31 VSUBS 0.515249f
C1134 VN.t2 VSUBS 1.28007f
C1135 VN.n32 VSUBS 0.561465f
C1136 VN.n33 VSUBS 0.230949f
C1137 VN.n34 VSUBS 0.050508f
C1138 VN.n35 VSUBS 0.059031f
C1139 VN.n36 VSUBS 0.071565f
C1140 VN.n37 VSUBS 0.04435f
C1141 VN.n38 VSUBS 0.04435f
C1142 VN.n39 VSUBS 0.04435f
C1143 VN.n40 VSUBS 0.071565f
C1144 VN.n41 VSUBS 0.059031f
C1145 VN.n42 VSUBS 0.050508f
C1146 VN.n43 VSUBS 0.04435f
C1147 VN.n44 VSUBS 0.04435f
C1148 VN.n45 VSUBS 0.04435f
C1149 VN.n46 VSUBS 0.042062f
C1150 VN.n47 VSUBS 0.065082f
C1151 VN.n48 VSUBS 0.529628f
C1152 VN.n49 VSUBS 1.91213f
.ends

