* NGSPICE file created from diff_pair_sample_1258.ext - technology: sky130A

.subckt diff_pair_sample_1258 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.6435 ps=4.08 w=1.65 l=0.53
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0 ps=0 w=1.65 l=0.53
X2 VDD1.t4 VP.t1 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.6435 ps=4.08 w=1.65 l=0.53
X3 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0 ps=0 w=1.65 l=0.53
X4 VDD1.t3 VP.t2 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0.27225 ps=1.98 w=1.65 l=0.53
X5 VTAIL.t10 VN.t0 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.27225 ps=1.98 w=1.65 l=0.53
X6 VDD1.t2 VP.t3 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0.27225 ps=1.98 w=1.65 l=0.53
X7 VTAIL.t3 VN.t1 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.27225 ps=1.98 w=1.65 l=0.53
X8 VDD2.t3 VN.t2 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0.27225 ps=1.98 w=1.65 l=0.53
X9 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0.27225 ps=1.98 w=1.65 l=0.53
X10 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0 ps=0 w=1.65 l=0.53
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6435 pd=4.08 as=0 ps=0 w=1.65 l=0.53
X12 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.6435 ps=4.08 w=1.65 l=0.53
X13 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.6435 ps=4.08 w=1.65 l=0.53
X14 VTAIL.t7 VP.t4 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.27225 ps=1.98 w=1.65 l=0.53
X15 VTAIL.t9 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.27225 pd=1.98 as=0.27225 ps=1.98 w=1.65 l=0.53
R0 VP.n1 VP.t3 176.423
R1 VP.n9 VP.n8 161.3
R2 VP.n4 VP.n3 161.3
R3 VP.n6 VP.n5 161.3
R4 VP.n6 VP.t2 149.602
R5 VP.n7 VP.t5 149.602
R6 VP.n8 VP.t1 149.602
R7 VP.n3 VP.t0 149.602
R8 VP.n2 VP.t4 149.602
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 32.7126
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VTAIL.n11 VTAIL.t2 111.492
R20 VTAIL.n2 VTAIL.t5 111.492
R21 VTAIL.n10 VTAIL.t8 111.492
R22 VTAIL.n7 VTAIL.t1 111.492
R23 VTAIL.n1 VTAIL.n0 99.4915
R24 VTAIL.n4 VTAIL.n3 99.4915
R25 VTAIL.n9 VTAIL.n8 99.4915
R26 VTAIL.n6 VTAIL.n5 99.4915
R27 VTAIL.n6 VTAIL.n4 15.2721
R28 VTAIL.n11 VTAIL.n10 14.5307
R29 VTAIL.n0 VTAIL.t0 12.0005
R30 VTAIL.n0 VTAIL.t3 12.0005
R31 VTAIL.n3 VTAIL.t4 12.0005
R32 VTAIL.n3 VTAIL.t9 12.0005
R33 VTAIL.n8 VTAIL.t6 12.0005
R34 VTAIL.n8 VTAIL.t7 12.0005
R35 VTAIL.n5 VTAIL.t11 12.0005
R36 VTAIL.n5 VTAIL.t10 12.0005
R37 VTAIL.n9 VTAIL.n7 0.841017
R38 VTAIL.n2 VTAIL.n1 0.841017
R39 VTAIL.n7 VTAIL.n6 0.741879
R40 VTAIL.n10 VTAIL.n9 0.741879
R41 VTAIL.n4 VTAIL.n2 0.741879
R42 VTAIL VTAIL.n11 0.498345
R43 VTAIL VTAIL.n1 0.244034
R44 VDD1 VDD1.t2 128.785
R45 VDD1.n1 VDD1.t3 128.671
R46 VDD1.n1 VDD1.n0 116.3
R47 VDD1.n3 VDD1.n2 116.171
R48 VDD1.n3 VDD1.n1 28.5009
R49 VDD1.n2 VDD1.t1 12.0005
R50 VDD1.n2 VDD1.t5 12.0005
R51 VDD1.n0 VDD1.t0 12.0005
R52 VDD1.n0 VDD1.t4 12.0005
R53 VDD1 VDD1.n3 0.127655
R54 B.n255 B.n254 585
R55 B.n257 B.n57 585
R56 B.n260 B.n259 585
R57 B.n261 B.n56 585
R58 B.n263 B.n262 585
R59 B.n265 B.n55 585
R60 B.n268 B.n267 585
R61 B.n269 B.n54 585
R62 B.n271 B.n270 585
R63 B.n273 B.n53 585
R64 B.n276 B.n275 585
R65 B.n278 B.n50 585
R66 B.n280 B.n279 585
R67 B.n282 B.n49 585
R68 B.n285 B.n284 585
R69 B.n286 B.n48 585
R70 B.n288 B.n287 585
R71 B.n290 B.n47 585
R72 B.n293 B.n292 585
R73 B.n294 B.n43 585
R74 B.n296 B.n295 585
R75 B.n298 B.n42 585
R76 B.n301 B.n300 585
R77 B.n302 B.n41 585
R78 B.n304 B.n303 585
R79 B.n306 B.n40 585
R80 B.n309 B.n308 585
R81 B.n310 B.n39 585
R82 B.n312 B.n311 585
R83 B.n314 B.n38 585
R84 B.n317 B.n316 585
R85 B.n318 B.n37 585
R86 B.n253 B.n35 585
R87 B.n321 B.n35 585
R88 B.n252 B.n34 585
R89 B.n322 B.n34 585
R90 B.n251 B.n33 585
R91 B.n323 B.n33 585
R92 B.n250 B.n249 585
R93 B.n249 B.n29 585
R94 B.n248 B.n28 585
R95 B.n329 B.n28 585
R96 B.n247 B.n27 585
R97 B.n330 B.n27 585
R98 B.n246 B.n26 585
R99 B.n331 B.n26 585
R100 B.n245 B.n244 585
R101 B.n244 B.n22 585
R102 B.n243 B.n21 585
R103 B.n337 B.n21 585
R104 B.n242 B.n20 585
R105 B.n338 B.n20 585
R106 B.n241 B.n19 585
R107 B.n339 B.n19 585
R108 B.n240 B.n239 585
R109 B.n239 B.n15 585
R110 B.n238 B.n14 585
R111 B.n345 B.n14 585
R112 B.n237 B.n13 585
R113 B.n346 B.n13 585
R114 B.n236 B.n12 585
R115 B.n347 B.n12 585
R116 B.n235 B.n234 585
R117 B.n234 B.n11 585
R118 B.n233 B.n7 585
R119 B.n353 B.n7 585
R120 B.n232 B.n6 585
R121 B.n354 B.n6 585
R122 B.n231 B.n5 585
R123 B.n355 B.n5 585
R124 B.n230 B.n229 585
R125 B.n229 B.n4 585
R126 B.n228 B.n58 585
R127 B.n228 B.n227 585
R128 B.n217 B.n59 585
R129 B.n220 B.n59 585
R130 B.n219 B.n218 585
R131 B.n221 B.n219 585
R132 B.n216 B.n64 585
R133 B.n64 B.n63 585
R134 B.n215 B.n214 585
R135 B.n214 B.n213 585
R136 B.n66 B.n65 585
R137 B.n67 B.n66 585
R138 B.n206 B.n205 585
R139 B.n207 B.n206 585
R140 B.n204 B.n72 585
R141 B.n72 B.n71 585
R142 B.n203 B.n202 585
R143 B.n202 B.n201 585
R144 B.n74 B.n73 585
R145 B.n75 B.n74 585
R146 B.n194 B.n193 585
R147 B.n195 B.n194 585
R148 B.n192 B.n80 585
R149 B.n80 B.n79 585
R150 B.n191 B.n190 585
R151 B.n190 B.n189 585
R152 B.n82 B.n81 585
R153 B.n83 B.n82 585
R154 B.n182 B.n181 585
R155 B.n183 B.n182 585
R156 B.n180 B.n88 585
R157 B.n88 B.n87 585
R158 B.n179 B.n178 585
R159 B.n178 B.n177 585
R160 B.n174 B.n92 585
R161 B.n173 B.n172 585
R162 B.n170 B.n93 585
R163 B.n170 B.n91 585
R164 B.n169 B.n168 585
R165 B.n167 B.n166 585
R166 B.n165 B.n95 585
R167 B.n163 B.n162 585
R168 B.n161 B.n96 585
R169 B.n160 B.n159 585
R170 B.n157 B.n97 585
R171 B.n155 B.n154 585
R172 B.n152 B.n98 585
R173 B.n151 B.n150 585
R174 B.n148 B.n101 585
R175 B.n146 B.n145 585
R176 B.n144 B.n102 585
R177 B.n143 B.n142 585
R178 B.n140 B.n103 585
R179 B.n138 B.n137 585
R180 B.n136 B.n104 585
R181 B.n135 B.n134 585
R182 B.n132 B.n131 585
R183 B.n130 B.n129 585
R184 B.n128 B.n109 585
R185 B.n126 B.n125 585
R186 B.n124 B.n110 585
R187 B.n123 B.n122 585
R188 B.n120 B.n111 585
R189 B.n118 B.n117 585
R190 B.n116 B.n112 585
R191 B.n115 B.n114 585
R192 B.n90 B.n89 585
R193 B.n91 B.n90 585
R194 B.n176 B.n175 585
R195 B.n177 B.n176 585
R196 B.n86 B.n85 585
R197 B.n87 B.n86 585
R198 B.n185 B.n184 585
R199 B.n184 B.n183 585
R200 B.n186 B.n84 585
R201 B.n84 B.n83 585
R202 B.n188 B.n187 585
R203 B.n189 B.n188 585
R204 B.n78 B.n77 585
R205 B.n79 B.n78 585
R206 B.n197 B.n196 585
R207 B.n196 B.n195 585
R208 B.n198 B.n76 585
R209 B.n76 B.n75 585
R210 B.n200 B.n199 585
R211 B.n201 B.n200 585
R212 B.n70 B.n69 585
R213 B.n71 B.n70 585
R214 B.n209 B.n208 585
R215 B.n208 B.n207 585
R216 B.n210 B.n68 585
R217 B.n68 B.n67 585
R218 B.n212 B.n211 585
R219 B.n213 B.n212 585
R220 B.n62 B.n61 585
R221 B.n63 B.n62 585
R222 B.n223 B.n222 585
R223 B.n222 B.n221 585
R224 B.n224 B.n60 585
R225 B.n220 B.n60 585
R226 B.n226 B.n225 585
R227 B.n227 B.n226 585
R228 B.n2 B.n0 585
R229 B.n4 B.n2 585
R230 B.n3 B.n1 585
R231 B.n354 B.n3 585
R232 B.n352 B.n351 585
R233 B.n353 B.n352 585
R234 B.n350 B.n8 585
R235 B.n11 B.n8 585
R236 B.n349 B.n348 585
R237 B.n348 B.n347 585
R238 B.n10 B.n9 585
R239 B.n346 B.n10 585
R240 B.n344 B.n343 585
R241 B.n345 B.n344 585
R242 B.n342 B.n16 585
R243 B.n16 B.n15 585
R244 B.n341 B.n340 585
R245 B.n340 B.n339 585
R246 B.n18 B.n17 585
R247 B.n338 B.n18 585
R248 B.n336 B.n335 585
R249 B.n337 B.n336 585
R250 B.n334 B.n23 585
R251 B.n23 B.n22 585
R252 B.n333 B.n332 585
R253 B.n332 B.n331 585
R254 B.n25 B.n24 585
R255 B.n330 B.n25 585
R256 B.n328 B.n327 585
R257 B.n329 B.n328 585
R258 B.n326 B.n30 585
R259 B.n30 B.n29 585
R260 B.n325 B.n324 585
R261 B.n324 B.n323 585
R262 B.n32 B.n31 585
R263 B.n322 B.n32 585
R264 B.n320 B.n319 585
R265 B.n321 B.n320 585
R266 B.n357 B.n356 585
R267 B.n356 B.n355 585
R268 B.n176 B.n92 530.939
R269 B.n320 B.n37 530.939
R270 B.n178 B.n90 530.939
R271 B.n255 B.n35 530.939
R272 B.n105 B.t10 280.755
R273 B.n99 B.t6 280.755
R274 B.n44 B.t13 280.755
R275 B.n51 B.t17 280.755
R276 B.n256 B.n36 256.663
R277 B.n258 B.n36 256.663
R278 B.n264 B.n36 256.663
R279 B.n266 B.n36 256.663
R280 B.n272 B.n36 256.663
R281 B.n274 B.n36 256.663
R282 B.n281 B.n36 256.663
R283 B.n283 B.n36 256.663
R284 B.n289 B.n36 256.663
R285 B.n291 B.n36 256.663
R286 B.n297 B.n36 256.663
R287 B.n299 B.n36 256.663
R288 B.n305 B.n36 256.663
R289 B.n307 B.n36 256.663
R290 B.n313 B.n36 256.663
R291 B.n315 B.n36 256.663
R292 B.n171 B.n91 256.663
R293 B.n94 B.n91 256.663
R294 B.n164 B.n91 256.663
R295 B.n158 B.n91 256.663
R296 B.n156 B.n91 256.663
R297 B.n149 B.n91 256.663
R298 B.n147 B.n91 256.663
R299 B.n141 B.n91 256.663
R300 B.n139 B.n91 256.663
R301 B.n133 B.n91 256.663
R302 B.n108 B.n91 256.663
R303 B.n127 B.n91 256.663
R304 B.n121 B.n91 256.663
R305 B.n119 B.n91 256.663
R306 B.n113 B.n91 256.663
R307 B.n177 B.n91 220.794
R308 B.n321 B.n36 220.794
R309 B.n176 B.n86 163.367
R310 B.n184 B.n86 163.367
R311 B.n184 B.n84 163.367
R312 B.n188 B.n84 163.367
R313 B.n188 B.n78 163.367
R314 B.n196 B.n78 163.367
R315 B.n196 B.n76 163.367
R316 B.n200 B.n76 163.367
R317 B.n200 B.n70 163.367
R318 B.n208 B.n70 163.367
R319 B.n208 B.n68 163.367
R320 B.n212 B.n68 163.367
R321 B.n212 B.n62 163.367
R322 B.n222 B.n62 163.367
R323 B.n222 B.n60 163.367
R324 B.n226 B.n60 163.367
R325 B.n226 B.n2 163.367
R326 B.n356 B.n2 163.367
R327 B.n356 B.n3 163.367
R328 B.n352 B.n3 163.367
R329 B.n352 B.n8 163.367
R330 B.n348 B.n8 163.367
R331 B.n348 B.n10 163.367
R332 B.n344 B.n10 163.367
R333 B.n344 B.n16 163.367
R334 B.n340 B.n16 163.367
R335 B.n340 B.n18 163.367
R336 B.n336 B.n18 163.367
R337 B.n336 B.n23 163.367
R338 B.n332 B.n23 163.367
R339 B.n332 B.n25 163.367
R340 B.n328 B.n25 163.367
R341 B.n328 B.n30 163.367
R342 B.n324 B.n30 163.367
R343 B.n324 B.n32 163.367
R344 B.n320 B.n32 163.367
R345 B.n172 B.n170 163.367
R346 B.n170 B.n169 163.367
R347 B.n166 B.n165 163.367
R348 B.n163 B.n96 163.367
R349 B.n159 B.n157 163.367
R350 B.n155 B.n98 163.367
R351 B.n150 B.n148 163.367
R352 B.n146 B.n102 163.367
R353 B.n142 B.n140 163.367
R354 B.n138 B.n104 163.367
R355 B.n134 B.n132 163.367
R356 B.n129 B.n128 163.367
R357 B.n126 B.n110 163.367
R358 B.n122 B.n120 163.367
R359 B.n118 B.n112 163.367
R360 B.n114 B.n90 163.367
R361 B.n178 B.n88 163.367
R362 B.n182 B.n88 163.367
R363 B.n182 B.n82 163.367
R364 B.n190 B.n82 163.367
R365 B.n190 B.n80 163.367
R366 B.n194 B.n80 163.367
R367 B.n194 B.n74 163.367
R368 B.n202 B.n74 163.367
R369 B.n202 B.n72 163.367
R370 B.n206 B.n72 163.367
R371 B.n206 B.n66 163.367
R372 B.n214 B.n66 163.367
R373 B.n214 B.n64 163.367
R374 B.n219 B.n64 163.367
R375 B.n219 B.n59 163.367
R376 B.n228 B.n59 163.367
R377 B.n229 B.n228 163.367
R378 B.n229 B.n5 163.367
R379 B.n6 B.n5 163.367
R380 B.n7 B.n6 163.367
R381 B.n234 B.n7 163.367
R382 B.n234 B.n12 163.367
R383 B.n13 B.n12 163.367
R384 B.n14 B.n13 163.367
R385 B.n239 B.n14 163.367
R386 B.n239 B.n19 163.367
R387 B.n20 B.n19 163.367
R388 B.n21 B.n20 163.367
R389 B.n244 B.n21 163.367
R390 B.n244 B.n26 163.367
R391 B.n27 B.n26 163.367
R392 B.n28 B.n27 163.367
R393 B.n249 B.n28 163.367
R394 B.n249 B.n33 163.367
R395 B.n34 B.n33 163.367
R396 B.n35 B.n34 163.367
R397 B.n316 B.n314 163.367
R398 B.n312 B.n39 163.367
R399 B.n308 B.n306 163.367
R400 B.n304 B.n41 163.367
R401 B.n300 B.n298 163.367
R402 B.n296 B.n43 163.367
R403 B.n292 B.n290 163.367
R404 B.n288 B.n48 163.367
R405 B.n284 B.n282 163.367
R406 B.n280 B.n50 163.367
R407 B.n275 B.n273 163.367
R408 B.n271 B.n54 163.367
R409 B.n267 B.n265 163.367
R410 B.n263 B.n56 163.367
R411 B.n259 B.n257 163.367
R412 B.n105 B.t12 125.728
R413 B.n51 B.t18 125.728
R414 B.n99 B.t9 125.727
R415 B.n44 B.t15 125.727
R416 B.n106 B.t11 109.049
R417 B.n52 B.t19 109.049
R418 B.n100 B.t8 109.049
R419 B.n45 B.t16 109.049
R420 B.n177 B.n87 108.014
R421 B.n183 B.n87 108.014
R422 B.n183 B.n83 108.014
R423 B.n189 B.n83 108.014
R424 B.n195 B.n79 108.014
R425 B.n195 B.n75 108.014
R426 B.n201 B.n75 108.014
R427 B.n201 B.n71 108.014
R428 B.n207 B.n71 108.014
R429 B.n213 B.n67 108.014
R430 B.n221 B.n63 108.014
R431 B.n221 B.n220 108.014
R432 B.n227 B.n4 108.014
R433 B.n355 B.n4 108.014
R434 B.n355 B.n354 108.014
R435 B.n354 B.n353 108.014
R436 B.n347 B.n11 108.014
R437 B.n347 B.n346 108.014
R438 B.n345 B.n15 108.014
R439 B.n339 B.n338 108.014
R440 B.n338 B.n337 108.014
R441 B.n337 B.n22 108.014
R442 B.n331 B.n22 108.014
R443 B.n331 B.n330 108.014
R444 B.n329 B.n29 108.014
R445 B.n323 B.n29 108.014
R446 B.n323 B.n322 108.014
R447 B.n322 B.n321 108.014
R448 B.t5 B.n67 100.073
R449 B.t2 B.n15 100.073
R450 B.n227 B.t1 93.7189
R451 B.n353 B.t0 93.7189
R452 B.n171 B.n92 71.676
R453 B.n169 B.n94 71.676
R454 B.n165 B.n164 71.676
R455 B.n158 B.n96 71.676
R456 B.n157 B.n156 71.676
R457 B.n149 B.n98 71.676
R458 B.n148 B.n147 71.676
R459 B.n141 B.n102 71.676
R460 B.n140 B.n139 71.676
R461 B.n133 B.n104 71.676
R462 B.n132 B.n108 71.676
R463 B.n128 B.n127 71.676
R464 B.n121 B.n110 71.676
R465 B.n120 B.n119 71.676
R466 B.n113 B.n112 71.676
R467 B.n315 B.n37 71.676
R468 B.n314 B.n313 71.676
R469 B.n307 B.n39 71.676
R470 B.n306 B.n305 71.676
R471 B.n299 B.n41 71.676
R472 B.n298 B.n297 71.676
R473 B.n291 B.n43 71.676
R474 B.n290 B.n289 71.676
R475 B.n283 B.n48 71.676
R476 B.n282 B.n281 71.676
R477 B.n274 B.n50 71.676
R478 B.n273 B.n272 71.676
R479 B.n266 B.n54 71.676
R480 B.n265 B.n264 71.676
R481 B.n258 B.n56 71.676
R482 B.n257 B.n256 71.676
R483 B.n256 B.n255 71.676
R484 B.n259 B.n258 71.676
R485 B.n264 B.n263 71.676
R486 B.n267 B.n266 71.676
R487 B.n272 B.n271 71.676
R488 B.n275 B.n274 71.676
R489 B.n281 B.n280 71.676
R490 B.n284 B.n283 71.676
R491 B.n289 B.n288 71.676
R492 B.n292 B.n291 71.676
R493 B.n297 B.n296 71.676
R494 B.n300 B.n299 71.676
R495 B.n305 B.n304 71.676
R496 B.n308 B.n307 71.676
R497 B.n313 B.n312 71.676
R498 B.n316 B.n315 71.676
R499 B.n172 B.n171 71.676
R500 B.n166 B.n94 71.676
R501 B.n164 B.n163 71.676
R502 B.n159 B.n158 71.676
R503 B.n156 B.n155 71.676
R504 B.n150 B.n149 71.676
R505 B.n147 B.n146 71.676
R506 B.n142 B.n141 71.676
R507 B.n139 B.n138 71.676
R508 B.n134 B.n133 71.676
R509 B.n129 B.n108 71.676
R510 B.n127 B.n126 71.676
R511 B.n122 B.n121 71.676
R512 B.n119 B.n118 71.676
R513 B.n114 B.n113 71.676
R514 B.t7 B.n79 71.4806
R515 B.n330 B.t14 71.4806
R516 B.n213 B.t4 65.1269
R517 B.t3 B.n345 65.1269
R518 B.n107 B.n106 59.5399
R519 B.n153 B.n100 59.5399
R520 B.n46 B.n45 59.5399
R521 B.n277 B.n52 59.5399
R522 B.t4 B.n63 42.8886
R523 B.n346 B.t3 42.8886
R524 B.n189 B.t7 36.5348
R525 B.t14 B.n329 36.5348
R526 B.n319 B.n318 34.4981
R527 B.n254 B.n253 34.4981
R528 B.n179 B.n89 34.4981
R529 B.n175 B.n174 34.4981
R530 B B.n357 18.0485
R531 B.n106 B.n105 16.6793
R532 B.n100 B.n99 16.6793
R533 B.n45 B.n44 16.6793
R534 B.n52 B.n51 16.6793
R535 B.n220 B.t1 14.2965
R536 B.n11 B.t0 14.2965
R537 B.n318 B.n317 10.6151
R538 B.n317 B.n38 10.6151
R539 B.n311 B.n38 10.6151
R540 B.n311 B.n310 10.6151
R541 B.n310 B.n309 10.6151
R542 B.n309 B.n40 10.6151
R543 B.n303 B.n40 10.6151
R544 B.n303 B.n302 10.6151
R545 B.n302 B.n301 10.6151
R546 B.n301 B.n42 10.6151
R547 B.n295 B.n294 10.6151
R548 B.n294 B.n293 10.6151
R549 B.n293 B.n47 10.6151
R550 B.n287 B.n47 10.6151
R551 B.n287 B.n286 10.6151
R552 B.n286 B.n285 10.6151
R553 B.n285 B.n49 10.6151
R554 B.n279 B.n49 10.6151
R555 B.n279 B.n278 10.6151
R556 B.n276 B.n53 10.6151
R557 B.n270 B.n53 10.6151
R558 B.n270 B.n269 10.6151
R559 B.n269 B.n268 10.6151
R560 B.n268 B.n55 10.6151
R561 B.n262 B.n55 10.6151
R562 B.n262 B.n261 10.6151
R563 B.n261 B.n260 10.6151
R564 B.n260 B.n57 10.6151
R565 B.n254 B.n57 10.6151
R566 B.n180 B.n179 10.6151
R567 B.n181 B.n180 10.6151
R568 B.n181 B.n81 10.6151
R569 B.n191 B.n81 10.6151
R570 B.n192 B.n191 10.6151
R571 B.n193 B.n192 10.6151
R572 B.n193 B.n73 10.6151
R573 B.n203 B.n73 10.6151
R574 B.n204 B.n203 10.6151
R575 B.n205 B.n204 10.6151
R576 B.n205 B.n65 10.6151
R577 B.n215 B.n65 10.6151
R578 B.n216 B.n215 10.6151
R579 B.n218 B.n216 10.6151
R580 B.n218 B.n217 10.6151
R581 B.n217 B.n58 10.6151
R582 B.n230 B.n58 10.6151
R583 B.n231 B.n230 10.6151
R584 B.n232 B.n231 10.6151
R585 B.n233 B.n232 10.6151
R586 B.n235 B.n233 10.6151
R587 B.n236 B.n235 10.6151
R588 B.n237 B.n236 10.6151
R589 B.n238 B.n237 10.6151
R590 B.n240 B.n238 10.6151
R591 B.n241 B.n240 10.6151
R592 B.n242 B.n241 10.6151
R593 B.n243 B.n242 10.6151
R594 B.n245 B.n243 10.6151
R595 B.n246 B.n245 10.6151
R596 B.n247 B.n246 10.6151
R597 B.n248 B.n247 10.6151
R598 B.n250 B.n248 10.6151
R599 B.n251 B.n250 10.6151
R600 B.n252 B.n251 10.6151
R601 B.n253 B.n252 10.6151
R602 B.n174 B.n173 10.6151
R603 B.n173 B.n93 10.6151
R604 B.n168 B.n93 10.6151
R605 B.n168 B.n167 10.6151
R606 B.n167 B.n95 10.6151
R607 B.n162 B.n95 10.6151
R608 B.n162 B.n161 10.6151
R609 B.n161 B.n160 10.6151
R610 B.n160 B.n97 10.6151
R611 B.n154 B.n97 10.6151
R612 B.n152 B.n151 10.6151
R613 B.n151 B.n101 10.6151
R614 B.n145 B.n101 10.6151
R615 B.n145 B.n144 10.6151
R616 B.n144 B.n143 10.6151
R617 B.n143 B.n103 10.6151
R618 B.n137 B.n103 10.6151
R619 B.n137 B.n136 10.6151
R620 B.n136 B.n135 10.6151
R621 B.n131 B.n130 10.6151
R622 B.n130 B.n109 10.6151
R623 B.n125 B.n109 10.6151
R624 B.n125 B.n124 10.6151
R625 B.n124 B.n123 10.6151
R626 B.n123 B.n111 10.6151
R627 B.n117 B.n111 10.6151
R628 B.n117 B.n116 10.6151
R629 B.n116 B.n115 10.6151
R630 B.n115 B.n89 10.6151
R631 B.n175 B.n85 10.6151
R632 B.n185 B.n85 10.6151
R633 B.n186 B.n185 10.6151
R634 B.n187 B.n186 10.6151
R635 B.n187 B.n77 10.6151
R636 B.n197 B.n77 10.6151
R637 B.n198 B.n197 10.6151
R638 B.n199 B.n198 10.6151
R639 B.n199 B.n69 10.6151
R640 B.n209 B.n69 10.6151
R641 B.n210 B.n209 10.6151
R642 B.n211 B.n210 10.6151
R643 B.n211 B.n61 10.6151
R644 B.n223 B.n61 10.6151
R645 B.n224 B.n223 10.6151
R646 B.n225 B.n224 10.6151
R647 B.n225 B.n0 10.6151
R648 B.n351 B.n1 10.6151
R649 B.n351 B.n350 10.6151
R650 B.n350 B.n349 10.6151
R651 B.n349 B.n9 10.6151
R652 B.n343 B.n9 10.6151
R653 B.n343 B.n342 10.6151
R654 B.n342 B.n341 10.6151
R655 B.n341 B.n17 10.6151
R656 B.n335 B.n17 10.6151
R657 B.n335 B.n334 10.6151
R658 B.n334 B.n333 10.6151
R659 B.n333 B.n24 10.6151
R660 B.n327 B.n24 10.6151
R661 B.n327 B.n326 10.6151
R662 B.n326 B.n325 10.6151
R663 B.n325 B.n31 10.6151
R664 B.n319 B.n31 10.6151
R665 B.n46 B.n42 9.36635
R666 B.n277 B.n276 9.36635
R667 B.n154 B.n153 9.36635
R668 B.n131 B.n107 9.36635
R669 B.n207 B.t5 7.94274
R670 B.n339 B.t2 7.94274
R671 B.n357 B.n0 2.81026
R672 B.n357 B.n1 2.81026
R673 B.n295 B.n46 1.24928
R674 B.n278 B.n277 1.24928
R675 B.n153 B.n152 1.24928
R676 B.n135 B.n107 1.24928
R677 VN.n0 VN.t3 176.423
R678 VN.n4 VN.t4 176.423
R679 VN.n3 VN.n2 161.3
R680 VN.n7 VN.n6 161.3
R681 VN.n1 VN.t1 149.602
R682 VN.n2 VN.t5 149.602
R683 VN.n5 VN.t0 149.602
R684 VN.n6 VN.t2 149.602
R685 VN.n2 VN.n1 48.2005
R686 VN.n6 VN.n5 48.2005
R687 VN.n7 VN.n4 45.1367
R688 VN.n3 VN.n0 45.1367
R689 VN VN.n7 33.0933
R690 VN.n5 VN.n4 13.3799
R691 VN.n1 VN.n0 13.3799
R692 VN VN.n3 0.0516364
R693 VDD2.n1 VDD2.t2 128.671
R694 VDD2.n2 VDD2.t3 128.171
R695 VDD2.n1 VDD2.n0 116.3
R696 VDD2 VDD2.n3 116.297
R697 VDD2.n2 VDD2.n1 27.5472
R698 VDD2.n3 VDD2.t5 12.0005
R699 VDD2.n3 VDD2.t1 12.0005
R700 VDD2.n0 VDD2.t4 12.0005
R701 VDD2.n0 VDD2.t0 12.0005
R702 VDD2 VDD2.n2 0.614724
C0 VDD2 VDD1 0.647384f
C1 VTAIL VP 0.970176f
C2 VDD1 VTAIL 3.02808f
C3 VDD2 VN 0.795877f
C4 VDD1 VP 0.928598f
C5 VTAIL VN 0.955993f
C6 VDD2 VTAIL 3.06666f
C7 VN VP 3.0082f
C8 VDD1 VN 0.154872f
C9 VDD2 VP 0.289398f
C10 VDD2 B 2.40908f
C11 VDD1 B 2.575455f
C12 VTAIL B 2.26642f
C13 VN B 5.397115f
C14 VP B 4.39247f
C15 VDD2.t2 B 0.197303f
C16 VDD2.t4 B 0.025257f
C17 VDD2.t0 B 0.025257f
C18 VDD2.n0 B 0.145562f
C19 VDD2.n1 B 1.03122f
C20 VDD2.t3 B 0.196518f
C21 VDD2.n2 B 1.03048f
C22 VDD2.t5 B 0.025257f
C23 VDD2.t1 B 0.025257f
C24 VDD2.n3 B 0.145553f
C25 VN.t3 B 0.102142f
C26 VN.n0 B 0.061642f
C27 VN.t1 B 0.091195f
C28 VN.n1 B 0.079395f
C29 VN.t5 B 0.091195f
C30 VN.n2 B 0.071917f
C31 VN.n3 B 0.128795f
C32 VN.t4 B 0.102142f
C33 VN.n4 B 0.061642f
C34 VN.t0 B 0.091195f
C35 VN.n5 B 0.079395f
C36 VN.t2 B 0.091195f
C37 VN.n6 B 0.071917f
C38 VN.n7 B 0.983267f
C39 VDD1.t2 B 0.186827f
C40 VDD1.t3 B 0.186631f
C41 VDD1.t0 B 0.02389f
C42 VDD1.t4 B 0.02389f
C43 VDD1.n0 B 0.137688f
C44 VDD1.n1 B 1.02568f
C45 VDD1.t1 B 0.02389f
C46 VDD1.t5 B 0.02389f
C47 VDD1.n2 B 0.137467f
C48 VDD1.n3 B 0.990462f
C49 VTAIL.t0 B 0.031772f
C50 VTAIL.t3 B 0.031772f
C51 VTAIL.n0 B 0.153167f
C52 VTAIL.n1 B 0.263145f
C53 VTAIL.t5 B 0.217425f
C54 VTAIL.n2 B 0.324627f
C55 VTAIL.t4 B 0.031772f
C56 VTAIL.t9 B 0.031772f
C57 VTAIL.n3 B 0.153167f
C58 VTAIL.n4 B 0.795342f
C59 VTAIL.t11 B 0.031772f
C60 VTAIL.t10 B 0.031772f
C61 VTAIL.n5 B 0.153168f
C62 VTAIL.n6 B 0.795341f
C63 VTAIL.t1 B 0.217426f
C64 VTAIL.n7 B 0.324626f
C65 VTAIL.t6 B 0.031772f
C66 VTAIL.t7 B 0.031772f
C67 VTAIL.n8 B 0.153168f
C68 VTAIL.n9 B 0.302234f
C69 VTAIL.t8 B 0.217426f
C70 VTAIL.n10 B 0.759523f
C71 VTAIL.t2 B 0.217425f
C72 VTAIL.n11 B 0.740403f
C73 VP.n0 B 0.044553f
C74 VP.t3 B 0.103743f
C75 VP.n1 B 0.062609f
C76 VP.t0 B 0.092625f
C77 VP.t4 B 0.092625f
C78 VP.n2 B 0.08064f
C79 VP.n3 B 0.073045f
C80 VP.n4 B 0.976324f
C81 VP.n5 B 0.919412f
C82 VP.t2 B 0.092625f
C83 VP.n6 B 0.073045f
C84 VP.t5 B 0.092625f
C85 VP.n7 B 0.08064f
C86 VP.t1 B 0.092625f
C87 VP.n8 B 0.073045f
C88 VP.n9 B 0.037127f
.ends

