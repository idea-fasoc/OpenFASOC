* NGSPICE file created from diff_pair_sample_0277.ext - technology: sky130A

.subckt diff_pair_sample_0277 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=2.6091 ps=14.16 w=6.69 l=2.01
X1 VTAIL.t0 VN.t0 VDD2.t5 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=1.10385 ps=7.02 w=6.69 l=2.01
X2 VDD2.t4 VN.t1 VTAIL.t1 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=1.10385 ps=7.02 w=6.69 l=2.01
X3 B.t11 B.t9 B.t10 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=0 ps=0 w=6.69 l=2.01
X4 B.t8 B.t6 B.t7 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=0 ps=0 w=6.69 l=2.01
X5 VDD2.t3 VN.t2 VTAIL.t2 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=1.10385 ps=7.02 w=6.69 l=2.01
X6 VTAIL.t10 VP.t1 VDD1.t4 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=1.10385 ps=7.02 w=6.69 l=2.01
X7 VDD1.t3 VP.t2 VTAIL.t9 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=1.10385 ps=7.02 w=6.69 l=2.01
X8 VTAIL.t3 VN.t3 VDD2.t2 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=1.10385 ps=7.02 w=6.69 l=2.01
X9 VDD2.t1 VN.t4 VTAIL.t5 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=2.6091 ps=14.16 w=6.69 l=2.01
X10 VDD1.t2 VP.t3 VTAIL.t7 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=1.10385 ps=7.02 w=6.69 l=2.01
X11 B.t5 B.t3 B.t4 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=0 ps=0 w=6.69 l=2.01
X12 B.t2 B.t0 B.t1 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=2.6091 pd=14.16 as=0 ps=0 w=6.69 l=2.01
X13 VTAIL.t6 VP.t4 VDD1.t1 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=1.10385 ps=7.02 w=6.69 l=2.01
X14 VDD2.t0 VN.t5 VTAIL.t4 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=2.6091 ps=14.16 w=6.69 l=2.01
X15 VDD1.t0 VP.t5 VTAIL.t11 w_n2842_n2306# sky130_fd_pr__pfet_01v8 ad=1.10385 pd=7.02 as=2.6091 ps=14.16 w=6.69 l=2.01
R0 VP.n10 VP.n9 161.3
R1 VP.n11 VP.n6 161.3
R2 VP.n13 VP.n12 161.3
R3 VP.n14 VP.n5 161.3
R4 VP.n31 VP.n0 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n28 VP.n1 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n25 VP.n2 161.3
R9 VP.n24 VP.n23 161.3
R10 VP.n22 VP.n3 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n19 VP.n4 161.3
R13 VP.n7 VP.t3 113.751
R14 VP.n18 VP.n17 94.1189
R15 VP.n33 VP.n32 94.1189
R16 VP.n16 VP.n15 94.1189
R17 VP.n25 VP.t4 80.2139
R18 VP.n18 VP.t2 80.2139
R19 VP.n32 VP.t5 80.2139
R20 VP.n8 VP.t1 80.2139
R21 VP.n15 VP.t0 80.2139
R22 VP.n20 VP.n3 56.5193
R23 VP.n30 VP.n1 56.5193
R24 VP.n13 VP.n6 56.5193
R25 VP.n8 VP.n7 45.7559
R26 VP.n17 VP.n16 42.3178
R27 VP.n20 VP.n19 24.4675
R28 VP.n24 VP.n3 24.4675
R29 VP.n25 VP.n24 24.4675
R30 VP.n26 VP.n25 24.4675
R31 VP.n26 VP.n1 24.4675
R32 VP.n31 VP.n30 24.4675
R33 VP.n14 VP.n13 24.4675
R34 VP.n9 VP.n8 24.4675
R35 VP.n9 VP.n6 24.4675
R36 VP.n19 VP.n18 16.6381
R37 VP.n32 VP.n31 16.6381
R38 VP.n15 VP.n14 16.6381
R39 VP.n10 VP.n7 9.28439
R40 VP.n16 VP.n5 0.278367
R41 VP.n17 VP.n4 0.278367
R42 VP.n33 VP.n0 0.278367
R43 VP.n11 VP.n10 0.189894
R44 VP.n12 VP.n11 0.189894
R45 VP.n12 VP.n5 0.189894
R46 VP.n21 VP.n4 0.189894
R47 VP.n22 VP.n21 0.189894
R48 VP.n23 VP.n22 0.189894
R49 VP.n23 VP.n2 0.189894
R50 VP.n27 VP.n2 0.189894
R51 VP.n28 VP.n27 0.189894
R52 VP.n29 VP.n28 0.189894
R53 VP.n29 VP.n0 0.189894
R54 VP VP.n33 0.153454
R55 VTAIL.n146 VTAIL.n116 756.745
R56 VTAIL.n32 VTAIL.n2 756.745
R57 VTAIL.n110 VTAIL.n80 756.745
R58 VTAIL.n72 VTAIL.n42 756.745
R59 VTAIL.n129 VTAIL.n128 585
R60 VTAIL.n131 VTAIL.n130 585
R61 VTAIL.n124 VTAIL.n123 585
R62 VTAIL.n137 VTAIL.n136 585
R63 VTAIL.n139 VTAIL.n138 585
R64 VTAIL.n120 VTAIL.n119 585
R65 VTAIL.n145 VTAIL.n144 585
R66 VTAIL.n147 VTAIL.n146 585
R67 VTAIL.n15 VTAIL.n14 585
R68 VTAIL.n17 VTAIL.n16 585
R69 VTAIL.n10 VTAIL.n9 585
R70 VTAIL.n23 VTAIL.n22 585
R71 VTAIL.n25 VTAIL.n24 585
R72 VTAIL.n6 VTAIL.n5 585
R73 VTAIL.n31 VTAIL.n30 585
R74 VTAIL.n33 VTAIL.n32 585
R75 VTAIL.n111 VTAIL.n110 585
R76 VTAIL.n109 VTAIL.n108 585
R77 VTAIL.n84 VTAIL.n83 585
R78 VTAIL.n103 VTAIL.n102 585
R79 VTAIL.n101 VTAIL.n100 585
R80 VTAIL.n88 VTAIL.n87 585
R81 VTAIL.n95 VTAIL.n94 585
R82 VTAIL.n93 VTAIL.n92 585
R83 VTAIL.n73 VTAIL.n72 585
R84 VTAIL.n71 VTAIL.n70 585
R85 VTAIL.n46 VTAIL.n45 585
R86 VTAIL.n65 VTAIL.n64 585
R87 VTAIL.n63 VTAIL.n62 585
R88 VTAIL.n50 VTAIL.n49 585
R89 VTAIL.n57 VTAIL.n56 585
R90 VTAIL.n55 VTAIL.n54 585
R91 VTAIL.n127 VTAIL.t4 327.514
R92 VTAIL.n13 VTAIL.t11 327.514
R93 VTAIL.n91 VTAIL.t8 327.514
R94 VTAIL.n53 VTAIL.t5 327.514
R95 VTAIL.n130 VTAIL.n129 171.744
R96 VTAIL.n130 VTAIL.n123 171.744
R97 VTAIL.n137 VTAIL.n123 171.744
R98 VTAIL.n138 VTAIL.n137 171.744
R99 VTAIL.n138 VTAIL.n119 171.744
R100 VTAIL.n145 VTAIL.n119 171.744
R101 VTAIL.n146 VTAIL.n145 171.744
R102 VTAIL.n16 VTAIL.n15 171.744
R103 VTAIL.n16 VTAIL.n9 171.744
R104 VTAIL.n23 VTAIL.n9 171.744
R105 VTAIL.n24 VTAIL.n23 171.744
R106 VTAIL.n24 VTAIL.n5 171.744
R107 VTAIL.n31 VTAIL.n5 171.744
R108 VTAIL.n32 VTAIL.n31 171.744
R109 VTAIL.n110 VTAIL.n109 171.744
R110 VTAIL.n109 VTAIL.n83 171.744
R111 VTAIL.n102 VTAIL.n83 171.744
R112 VTAIL.n102 VTAIL.n101 171.744
R113 VTAIL.n101 VTAIL.n87 171.744
R114 VTAIL.n94 VTAIL.n87 171.744
R115 VTAIL.n94 VTAIL.n93 171.744
R116 VTAIL.n72 VTAIL.n71 171.744
R117 VTAIL.n71 VTAIL.n45 171.744
R118 VTAIL.n64 VTAIL.n45 171.744
R119 VTAIL.n64 VTAIL.n63 171.744
R120 VTAIL.n63 VTAIL.n49 171.744
R121 VTAIL.n56 VTAIL.n49 171.744
R122 VTAIL.n56 VTAIL.n55 171.744
R123 VTAIL.n129 VTAIL.t4 85.8723
R124 VTAIL.n15 VTAIL.t11 85.8723
R125 VTAIL.n93 VTAIL.t8 85.8723
R126 VTAIL.n55 VTAIL.t5 85.8723
R127 VTAIL.n79 VTAIL.n78 71.1384
R128 VTAIL.n41 VTAIL.n40 71.1384
R129 VTAIL.n1 VTAIL.n0 71.1382
R130 VTAIL.n39 VTAIL.n38 71.1382
R131 VTAIL.n151 VTAIL.n150 31.6035
R132 VTAIL.n37 VTAIL.n36 31.6035
R133 VTAIL.n115 VTAIL.n114 31.6035
R134 VTAIL.n77 VTAIL.n76 31.6035
R135 VTAIL.n41 VTAIL.n39 22.1686
R136 VTAIL.n151 VTAIL.n115 20.1514
R137 VTAIL.n128 VTAIL.n127 16.3884
R138 VTAIL.n14 VTAIL.n13 16.3884
R139 VTAIL.n92 VTAIL.n91 16.3884
R140 VTAIL.n54 VTAIL.n53 16.3884
R141 VTAIL.n131 VTAIL.n126 12.8005
R142 VTAIL.n17 VTAIL.n12 12.8005
R143 VTAIL.n95 VTAIL.n90 12.8005
R144 VTAIL.n57 VTAIL.n52 12.8005
R145 VTAIL.n132 VTAIL.n124 12.0247
R146 VTAIL.n18 VTAIL.n10 12.0247
R147 VTAIL.n96 VTAIL.n88 12.0247
R148 VTAIL.n58 VTAIL.n50 12.0247
R149 VTAIL.n136 VTAIL.n135 11.249
R150 VTAIL.n22 VTAIL.n21 11.249
R151 VTAIL.n100 VTAIL.n99 11.249
R152 VTAIL.n62 VTAIL.n61 11.249
R153 VTAIL.n139 VTAIL.n122 10.4732
R154 VTAIL.n25 VTAIL.n8 10.4732
R155 VTAIL.n103 VTAIL.n86 10.4732
R156 VTAIL.n65 VTAIL.n48 10.4732
R157 VTAIL.n140 VTAIL.n120 9.69747
R158 VTAIL.n26 VTAIL.n6 9.69747
R159 VTAIL.n104 VTAIL.n84 9.69747
R160 VTAIL.n66 VTAIL.n46 9.69747
R161 VTAIL.n150 VTAIL.n149 9.45567
R162 VTAIL.n36 VTAIL.n35 9.45567
R163 VTAIL.n114 VTAIL.n113 9.45567
R164 VTAIL.n76 VTAIL.n75 9.45567
R165 VTAIL.n118 VTAIL.n117 9.3005
R166 VTAIL.n143 VTAIL.n142 9.3005
R167 VTAIL.n141 VTAIL.n140 9.3005
R168 VTAIL.n122 VTAIL.n121 9.3005
R169 VTAIL.n135 VTAIL.n134 9.3005
R170 VTAIL.n133 VTAIL.n132 9.3005
R171 VTAIL.n126 VTAIL.n125 9.3005
R172 VTAIL.n149 VTAIL.n148 9.3005
R173 VTAIL.n4 VTAIL.n3 9.3005
R174 VTAIL.n29 VTAIL.n28 9.3005
R175 VTAIL.n27 VTAIL.n26 9.3005
R176 VTAIL.n8 VTAIL.n7 9.3005
R177 VTAIL.n21 VTAIL.n20 9.3005
R178 VTAIL.n19 VTAIL.n18 9.3005
R179 VTAIL.n12 VTAIL.n11 9.3005
R180 VTAIL.n35 VTAIL.n34 9.3005
R181 VTAIL.n113 VTAIL.n112 9.3005
R182 VTAIL.n82 VTAIL.n81 9.3005
R183 VTAIL.n107 VTAIL.n106 9.3005
R184 VTAIL.n105 VTAIL.n104 9.3005
R185 VTAIL.n86 VTAIL.n85 9.3005
R186 VTAIL.n99 VTAIL.n98 9.3005
R187 VTAIL.n97 VTAIL.n96 9.3005
R188 VTAIL.n90 VTAIL.n89 9.3005
R189 VTAIL.n75 VTAIL.n74 9.3005
R190 VTAIL.n44 VTAIL.n43 9.3005
R191 VTAIL.n69 VTAIL.n68 9.3005
R192 VTAIL.n67 VTAIL.n66 9.3005
R193 VTAIL.n48 VTAIL.n47 9.3005
R194 VTAIL.n61 VTAIL.n60 9.3005
R195 VTAIL.n59 VTAIL.n58 9.3005
R196 VTAIL.n52 VTAIL.n51 9.3005
R197 VTAIL.n144 VTAIL.n143 8.92171
R198 VTAIL.n30 VTAIL.n29 8.92171
R199 VTAIL.n108 VTAIL.n107 8.92171
R200 VTAIL.n70 VTAIL.n69 8.92171
R201 VTAIL.n147 VTAIL.n118 8.14595
R202 VTAIL.n33 VTAIL.n4 8.14595
R203 VTAIL.n111 VTAIL.n82 8.14595
R204 VTAIL.n73 VTAIL.n44 8.14595
R205 VTAIL.n148 VTAIL.n116 7.3702
R206 VTAIL.n34 VTAIL.n2 7.3702
R207 VTAIL.n112 VTAIL.n80 7.3702
R208 VTAIL.n74 VTAIL.n42 7.3702
R209 VTAIL.n150 VTAIL.n116 6.59444
R210 VTAIL.n36 VTAIL.n2 6.59444
R211 VTAIL.n114 VTAIL.n80 6.59444
R212 VTAIL.n76 VTAIL.n42 6.59444
R213 VTAIL.n148 VTAIL.n147 5.81868
R214 VTAIL.n34 VTAIL.n33 5.81868
R215 VTAIL.n112 VTAIL.n111 5.81868
R216 VTAIL.n74 VTAIL.n73 5.81868
R217 VTAIL.n144 VTAIL.n118 5.04292
R218 VTAIL.n30 VTAIL.n4 5.04292
R219 VTAIL.n108 VTAIL.n82 5.04292
R220 VTAIL.n70 VTAIL.n44 5.04292
R221 VTAIL.n0 VTAIL.t2 4.85924
R222 VTAIL.n0 VTAIL.t0 4.85924
R223 VTAIL.n38 VTAIL.t9 4.85924
R224 VTAIL.n38 VTAIL.t6 4.85924
R225 VTAIL.n78 VTAIL.t7 4.85924
R226 VTAIL.n78 VTAIL.t10 4.85924
R227 VTAIL.n40 VTAIL.t1 4.85924
R228 VTAIL.n40 VTAIL.t3 4.85924
R229 VTAIL.n143 VTAIL.n120 4.26717
R230 VTAIL.n29 VTAIL.n6 4.26717
R231 VTAIL.n107 VTAIL.n84 4.26717
R232 VTAIL.n69 VTAIL.n46 4.26717
R233 VTAIL.n127 VTAIL.n125 3.71088
R234 VTAIL.n13 VTAIL.n11 3.71088
R235 VTAIL.n91 VTAIL.n89 3.71088
R236 VTAIL.n53 VTAIL.n51 3.71088
R237 VTAIL.n140 VTAIL.n139 3.49141
R238 VTAIL.n26 VTAIL.n25 3.49141
R239 VTAIL.n104 VTAIL.n103 3.49141
R240 VTAIL.n66 VTAIL.n65 3.49141
R241 VTAIL.n136 VTAIL.n122 2.71565
R242 VTAIL.n22 VTAIL.n8 2.71565
R243 VTAIL.n100 VTAIL.n86 2.71565
R244 VTAIL.n62 VTAIL.n48 2.71565
R245 VTAIL.n77 VTAIL.n41 2.01774
R246 VTAIL.n115 VTAIL.n79 2.01774
R247 VTAIL.n39 VTAIL.n37 2.01774
R248 VTAIL.n135 VTAIL.n124 1.93989
R249 VTAIL.n21 VTAIL.n10 1.93989
R250 VTAIL.n99 VTAIL.n88 1.93989
R251 VTAIL.n61 VTAIL.n50 1.93989
R252 VTAIL.n79 VTAIL.n77 1.47895
R253 VTAIL.n37 VTAIL.n1 1.47895
R254 VTAIL VTAIL.n151 1.45524
R255 VTAIL.n132 VTAIL.n131 1.16414
R256 VTAIL.n18 VTAIL.n17 1.16414
R257 VTAIL.n96 VTAIL.n95 1.16414
R258 VTAIL.n58 VTAIL.n57 1.16414
R259 VTAIL VTAIL.n1 0.563
R260 VTAIL.n128 VTAIL.n126 0.388379
R261 VTAIL.n14 VTAIL.n12 0.388379
R262 VTAIL.n92 VTAIL.n90 0.388379
R263 VTAIL.n54 VTAIL.n52 0.388379
R264 VTAIL.n133 VTAIL.n125 0.155672
R265 VTAIL.n134 VTAIL.n133 0.155672
R266 VTAIL.n134 VTAIL.n121 0.155672
R267 VTAIL.n141 VTAIL.n121 0.155672
R268 VTAIL.n142 VTAIL.n141 0.155672
R269 VTAIL.n142 VTAIL.n117 0.155672
R270 VTAIL.n149 VTAIL.n117 0.155672
R271 VTAIL.n19 VTAIL.n11 0.155672
R272 VTAIL.n20 VTAIL.n19 0.155672
R273 VTAIL.n20 VTAIL.n7 0.155672
R274 VTAIL.n27 VTAIL.n7 0.155672
R275 VTAIL.n28 VTAIL.n27 0.155672
R276 VTAIL.n28 VTAIL.n3 0.155672
R277 VTAIL.n35 VTAIL.n3 0.155672
R278 VTAIL.n113 VTAIL.n81 0.155672
R279 VTAIL.n106 VTAIL.n81 0.155672
R280 VTAIL.n106 VTAIL.n105 0.155672
R281 VTAIL.n105 VTAIL.n85 0.155672
R282 VTAIL.n98 VTAIL.n85 0.155672
R283 VTAIL.n98 VTAIL.n97 0.155672
R284 VTAIL.n97 VTAIL.n89 0.155672
R285 VTAIL.n75 VTAIL.n43 0.155672
R286 VTAIL.n68 VTAIL.n43 0.155672
R287 VTAIL.n68 VTAIL.n67 0.155672
R288 VTAIL.n67 VTAIL.n47 0.155672
R289 VTAIL.n60 VTAIL.n47 0.155672
R290 VTAIL.n60 VTAIL.n59 0.155672
R291 VTAIL.n59 VTAIL.n51 0.155672
R292 VDD1.n30 VDD1.n0 756.745
R293 VDD1.n65 VDD1.n35 756.745
R294 VDD1.n31 VDD1.n30 585
R295 VDD1.n29 VDD1.n28 585
R296 VDD1.n4 VDD1.n3 585
R297 VDD1.n23 VDD1.n22 585
R298 VDD1.n21 VDD1.n20 585
R299 VDD1.n8 VDD1.n7 585
R300 VDD1.n15 VDD1.n14 585
R301 VDD1.n13 VDD1.n12 585
R302 VDD1.n48 VDD1.n47 585
R303 VDD1.n50 VDD1.n49 585
R304 VDD1.n43 VDD1.n42 585
R305 VDD1.n56 VDD1.n55 585
R306 VDD1.n58 VDD1.n57 585
R307 VDD1.n39 VDD1.n38 585
R308 VDD1.n64 VDD1.n63 585
R309 VDD1.n66 VDD1.n65 585
R310 VDD1.n11 VDD1.t2 327.514
R311 VDD1.n46 VDD1.t3 327.514
R312 VDD1.n30 VDD1.n29 171.744
R313 VDD1.n29 VDD1.n3 171.744
R314 VDD1.n22 VDD1.n3 171.744
R315 VDD1.n22 VDD1.n21 171.744
R316 VDD1.n21 VDD1.n7 171.744
R317 VDD1.n14 VDD1.n7 171.744
R318 VDD1.n14 VDD1.n13 171.744
R319 VDD1.n49 VDD1.n48 171.744
R320 VDD1.n49 VDD1.n42 171.744
R321 VDD1.n56 VDD1.n42 171.744
R322 VDD1.n57 VDD1.n56 171.744
R323 VDD1.n57 VDD1.n38 171.744
R324 VDD1.n64 VDD1.n38 171.744
R325 VDD1.n65 VDD1.n64 171.744
R326 VDD1.n71 VDD1.n70 88.2659
R327 VDD1.n73 VDD1.n72 87.817
R328 VDD1.n13 VDD1.t2 85.8723
R329 VDD1.n48 VDD1.t3 85.8723
R330 VDD1 VDD1.n34 49.8534
R331 VDD1.n71 VDD1.n69 49.7399
R332 VDD1.n73 VDD1.n71 37.6302
R333 VDD1.n47 VDD1.n46 16.3884
R334 VDD1.n12 VDD1.n11 16.3884
R335 VDD1.n15 VDD1.n10 12.8005
R336 VDD1.n50 VDD1.n45 12.8005
R337 VDD1.n16 VDD1.n8 12.0247
R338 VDD1.n51 VDD1.n43 12.0247
R339 VDD1.n20 VDD1.n19 11.249
R340 VDD1.n55 VDD1.n54 11.249
R341 VDD1.n23 VDD1.n6 10.4732
R342 VDD1.n58 VDD1.n41 10.4732
R343 VDD1.n24 VDD1.n4 9.69747
R344 VDD1.n59 VDD1.n39 9.69747
R345 VDD1.n34 VDD1.n33 9.45567
R346 VDD1.n69 VDD1.n68 9.45567
R347 VDD1.n33 VDD1.n32 9.3005
R348 VDD1.n2 VDD1.n1 9.3005
R349 VDD1.n27 VDD1.n26 9.3005
R350 VDD1.n25 VDD1.n24 9.3005
R351 VDD1.n6 VDD1.n5 9.3005
R352 VDD1.n19 VDD1.n18 9.3005
R353 VDD1.n17 VDD1.n16 9.3005
R354 VDD1.n10 VDD1.n9 9.3005
R355 VDD1.n37 VDD1.n36 9.3005
R356 VDD1.n62 VDD1.n61 9.3005
R357 VDD1.n60 VDD1.n59 9.3005
R358 VDD1.n41 VDD1.n40 9.3005
R359 VDD1.n54 VDD1.n53 9.3005
R360 VDD1.n52 VDD1.n51 9.3005
R361 VDD1.n45 VDD1.n44 9.3005
R362 VDD1.n68 VDD1.n67 9.3005
R363 VDD1.n28 VDD1.n27 8.92171
R364 VDD1.n63 VDD1.n62 8.92171
R365 VDD1.n31 VDD1.n2 8.14595
R366 VDD1.n66 VDD1.n37 8.14595
R367 VDD1.n32 VDD1.n0 7.3702
R368 VDD1.n67 VDD1.n35 7.3702
R369 VDD1.n34 VDD1.n0 6.59444
R370 VDD1.n69 VDD1.n35 6.59444
R371 VDD1.n32 VDD1.n31 5.81868
R372 VDD1.n67 VDD1.n66 5.81868
R373 VDD1.n28 VDD1.n2 5.04292
R374 VDD1.n63 VDD1.n37 5.04292
R375 VDD1.n72 VDD1.t4 4.85924
R376 VDD1.n72 VDD1.t5 4.85924
R377 VDD1.n70 VDD1.t1 4.85924
R378 VDD1.n70 VDD1.t0 4.85924
R379 VDD1.n27 VDD1.n4 4.26717
R380 VDD1.n62 VDD1.n39 4.26717
R381 VDD1.n11 VDD1.n9 3.71088
R382 VDD1.n46 VDD1.n44 3.71088
R383 VDD1.n24 VDD1.n23 3.49141
R384 VDD1.n59 VDD1.n58 3.49141
R385 VDD1.n20 VDD1.n6 2.71565
R386 VDD1.n55 VDD1.n41 2.71565
R387 VDD1.n19 VDD1.n8 1.93989
R388 VDD1.n54 VDD1.n43 1.93989
R389 VDD1.n16 VDD1.n15 1.16414
R390 VDD1.n51 VDD1.n50 1.16414
R391 VDD1 VDD1.n73 0.446621
R392 VDD1.n12 VDD1.n10 0.388379
R393 VDD1.n47 VDD1.n45 0.388379
R394 VDD1.n33 VDD1.n1 0.155672
R395 VDD1.n26 VDD1.n1 0.155672
R396 VDD1.n26 VDD1.n25 0.155672
R397 VDD1.n25 VDD1.n5 0.155672
R398 VDD1.n18 VDD1.n5 0.155672
R399 VDD1.n18 VDD1.n17 0.155672
R400 VDD1.n17 VDD1.n9 0.155672
R401 VDD1.n52 VDD1.n44 0.155672
R402 VDD1.n53 VDD1.n52 0.155672
R403 VDD1.n53 VDD1.n40 0.155672
R404 VDD1.n60 VDD1.n40 0.155672
R405 VDD1.n61 VDD1.n60 0.155672
R406 VDD1.n61 VDD1.n36 0.155672
R407 VDD1.n68 VDD1.n36 0.155672
R408 VN.n21 VN.n12 161.3
R409 VN.n20 VN.n19 161.3
R410 VN.n18 VN.n13 161.3
R411 VN.n17 VN.n16 161.3
R412 VN.n9 VN.n0 161.3
R413 VN.n8 VN.n7 161.3
R414 VN.n6 VN.n1 161.3
R415 VN.n5 VN.n4 161.3
R416 VN.n2 VN.t2 113.751
R417 VN.n14 VN.t4 113.751
R418 VN.n11 VN.n10 94.1189
R419 VN.n23 VN.n22 94.1189
R420 VN.n3 VN.t0 80.2139
R421 VN.n10 VN.t5 80.2139
R422 VN.n15 VN.t3 80.2139
R423 VN.n22 VN.t1 80.2139
R424 VN.n8 VN.n1 56.5193
R425 VN.n20 VN.n13 56.5193
R426 VN.n15 VN.n14 45.7559
R427 VN.n3 VN.n2 45.7559
R428 VN VN.n23 42.5966
R429 VN.n4 VN.n3 24.4675
R430 VN.n4 VN.n1 24.4675
R431 VN.n9 VN.n8 24.4675
R432 VN.n16 VN.n13 24.4675
R433 VN.n16 VN.n15 24.4675
R434 VN.n21 VN.n20 24.4675
R435 VN.n10 VN.n9 16.6381
R436 VN.n22 VN.n21 16.6381
R437 VN.n17 VN.n14 9.28439
R438 VN.n5 VN.n2 9.28439
R439 VN.n23 VN.n12 0.278367
R440 VN.n11 VN.n0 0.278367
R441 VN.n19 VN.n12 0.189894
R442 VN.n19 VN.n18 0.189894
R443 VN.n18 VN.n17 0.189894
R444 VN.n6 VN.n5 0.189894
R445 VN.n7 VN.n6 0.189894
R446 VN.n7 VN.n0 0.189894
R447 VN VN.n11 0.153454
R448 VDD2.n67 VDD2.n37 756.745
R449 VDD2.n30 VDD2.n0 756.745
R450 VDD2.n68 VDD2.n67 585
R451 VDD2.n66 VDD2.n65 585
R452 VDD2.n41 VDD2.n40 585
R453 VDD2.n60 VDD2.n59 585
R454 VDD2.n58 VDD2.n57 585
R455 VDD2.n45 VDD2.n44 585
R456 VDD2.n52 VDD2.n51 585
R457 VDD2.n50 VDD2.n49 585
R458 VDD2.n13 VDD2.n12 585
R459 VDD2.n15 VDD2.n14 585
R460 VDD2.n8 VDD2.n7 585
R461 VDD2.n21 VDD2.n20 585
R462 VDD2.n23 VDD2.n22 585
R463 VDD2.n4 VDD2.n3 585
R464 VDD2.n29 VDD2.n28 585
R465 VDD2.n31 VDD2.n30 585
R466 VDD2.n48 VDD2.t4 327.514
R467 VDD2.n11 VDD2.t3 327.514
R468 VDD2.n67 VDD2.n66 171.744
R469 VDD2.n66 VDD2.n40 171.744
R470 VDD2.n59 VDD2.n40 171.744
R471 VDD2.n59 VDD2.n58 171.744
R472 VDD2.n58 VDD2.n44 171.744
R473 VDD2.n51 VDD2.n44 171.744
R474 VDD2.n51 VDD2.n50 171.744
R475 VDD2.n14 VDD2.n13 171.744
R476 VDD2.n14 VDD2.n7 171.744
R477 VDD2.n21 VDD2.n7 171.744
R478 VDD2.n22 VDD2.n21 171.744
R479 VDD2.n22 VDD2.n3 171.744
R480 VDD2.n29 VDD2.n3 171.744
R481 VDD2.n30 VDD2.n29 171.744
R482 VDD2.n36 VDD2.n35 88.2659
R483 VDD2 VDD2.n73 88.2631
R484 VDD2.n50 VDD2.t4 85.8723
R485 VDD2.n13 VDD2.t3 85.8723
R486 VDD2.n36 VDD2.n34 49.7399
R487 VDD2.n72 VDD2.n71 48.2823
R488 VDD2.n72 VDD2.n36 36.0386
R489 VDD2.n12 VDD2.n11 16.3884
R490 VDD2.n49 VDD2.n48 16.3884
R491 VDD2.n52 VDD2.n47 12.8005
R492 VDD2.n15 VDD2.n10 12.8005
R493 VDD2.n53 VDD2.n45 12.0247
R494 VDD2.n16 VDD2.n8 12.0247
R495 VDD2.n57 VDD2.n56 11.249
R496 VDD2.n20 VDD2.n19 11.249
R497 VDD2.n60 VDD2.n43 10.4732
R498 VDD2.n23 VDD2.n6 10.4732
R499 VDD2.n61 VDD2.n41 9.69747
R500 VDD2.n24 VDD2.n4 9.69747
R501 VDD2.n71 VDD2.n70 9.45567
R502 VDD2.n34 VDD2.n33 9.45567
R503 VDD2.n70 VDD2.n69 9.3005
R504 VDD2.n39 VDD2.n38 9.3005
R505 VDD2.n64 VDD2.n63 9.3005
R506 VDD2.n62 VDD2.n61 9.3005
R507 VDD2.n43 VDD2.n42 9.3005
R508 VDD2.n56 VDD2.n55 9.3005
R509 VDD2.n54 VDD2.n53 9.3005
R510 VDD2.n47 VDD2.n46 9.3005
R511 VDD2.n2 VDD2.n1 9.3005
R512 VDD2.n27 VDD2.n26 9.3005
R513 VDD2.n25 VDD2.n24 9.3005
R514 VDD2.n6 VDD2.n5 9.3005
R515 VDD2.n19 VDD2.n18 9.3005
R516 VDD2.n17 VDD2.n16 9.3005
R517 VDD2.n10 VDD2.n9 9.3005
R518 VDD2.n33 VDD2.n32 9.3005
R519 VDD2.n65 VDD2.n64 8.92171
R520 VDD2.n28 VDD2.n27 8.92171
R521 VDD2.n68 VDD2.n39 8.14595
R522 VDD2.n31 VDD2.n2 8.14595
R523 VDD2.n69 VDD2.n37 7.3702
R524 VDD2.n32 VDD2.n0 7.3702
R525 VDD2.n71 VDD2.n37 6.59444
R526 VDD2.n34 VDD2.n0 6.59444
R527 VDD2.n69 VDD2.n68 5.81868
R528 VDD2.n32 VDD2.n31 5.81868
R529 VDD2.n65 VDD2.n39 5.04292
R530 VDD2.n28 VDD2.n2 5.04292
R531 VDD2.n73 VDD2.t2 4.85924
R532 VDD2.n73 VDD2.t1 4.85924
R533 VDD2.n35 VDD2.t5 4.85924
R534 VDD2.n35 VDD2.t0 4.85924
R535 VDD2.n64 VDD2.n41 4.26717
R536 VDD2.n27 VDD2.n4 4.26717
R537 VDD2.n48 VDD2.n46 3.71088
R538 VDD2.n11 VDD2.n9 3.71088
R539 VDD2.n61 VDD2.n60 3.49141
R540 VDD2.n24 VDD2.n23 3.49141
R541 VDD2.n57 VDD2.n43 2.71565
R542 VDD2.n20 VDD2.n6 2.71565
R543 VDD2.n56 VDD2.n45 1.93989
R544 VDD2.n19 VDD2.n8 1.93989
R545 VDD2 VDD2.n72 1.57162
R546 VDD2.n53 VDD2.n52 1.16414
R547 VDD2.n16 VDD2.n15 1.16414
R548 VDD2.n49 VDD2.n47 0.388379
R549 VDD2.n12 VDD2.n10 0.388379
R550 VDD2.n70 VDD2.n38 0.155672
R551 VDD2.n63 VDD2.n38 0.155672
R552 VDD2.n63 VDD2.n62 0.155672
R553 VDD2.n62 VDD2.n42 0.155672
R554 VDD2.n55 VDD2.n42 0.155672
R555 VDD2.n55 VDD2.n54 0.155672
R556 VDD2.n54 VDD2.n46 0.155672
R557 VDD2.n17 VDD2.n9 0.155672
R558 VDD2.n18 VDD2.n17 0.155672
R559 VDD2.n18 VDD2.n5 0.155672
R560 VDD2.n25 VDD2.n5 0.155672
R561 VDD2.n26 VDD2.n25 0.155672
R562 VDD2.n26 VDD2.n1 0.155672
R563 VDD2.n33 VDD2.n1 0.155672
R564 B.n289 B.n288 585
R565 B.n287 B.n92 585
R566 B.n286 B.n285 585
R567 B.n284 B.n93 585
R568 B.n283 B.n282 585
R569 B.n281 B.n94 585
R570 B.n280 B.n279 585
R571 B.n278 B.n95 585
R572 B.n277 B.n276 585
R573 B.n275 B.n96 585
R574 B.n274 B.n273 585
R575 B.n272 B.n97 585
R576 B.n271 B.n270 585
R577 B.n269 B.n98 585
R578 B.n268 B.n267 585
R579 B.n266 B.n99 585
R580 B.n265 B.n264 585
R581 B.n263 B.n100 585
R582 B.n262 B.n261 585
R583 B.n260 B.n101 585
R584 B.n259 B.n258 585
R585 B.n257 B.n102 585
R586 B.n256 B.n255 585
R587 B.n254 B.n103 585
R588 B.n253 B.n252 585
R589 B.n251 B.n104 585
R590 B.n249 B.n248 585
R591 B.n247 B.n107 585
R592 B.n246 B.n245 585
R593 B.n244 B.n108 585
R594 B.n243 B.n242 585
R595 B.n241 B.n109 585
R596 B.n240 B.n239 585
R597 B.n238 B.n110 585
R598 B.n237 B.n236 585
R599 B.n235 B.n111 585
R600 B.n234 B.n233 585
R601 B.n229 B.n112 585
R602 B.n228 B.n227 585
R603 B.n226 B.n113 585
R604 B.n225 B.n224 585
R605 B.n223 B.n114 585
R606 B.n222 B.n221 585
R607 B.n220 B.n115 585
R608 B.n219 B.n218 585
R609 B.n217 B.n116 585
R610 B.n216 B.n215 585
R611 B.n214 B.n117 585
R612 B.n213 B.n212 585
R613 B.n211 B.n118 585
R614 B.n210 B.n209 585
R615 B.n208 B.n119 585
R616 B.n207 B.n206 585
R617 B.n205 B.n120 585
R618 B.n204 B.n203 585
R619 B.n202 B.n121 585
R620 B.n201 B.n200 585
R621 B.n199 B.n122 585
R622 B.n198 B.n197 585
R623 B.n196 B.n123 585
R624 B.n195 B.n194 585
R625 B.n193 B.n124 585
R626 B.n290 B.n91 585
R627 B.n292 B.n291 585
R628 B.n293 B.n90 585
R629 B.n295 B.n294 585
R630 B.n296 B.n89 585
R631 B.n298 B.n297 585
R632 B.n299 B.n88 585
R633 B.n301 B.n300 585
R634 B.n302 B.n87 585
R635 B.n304 B.n303 585
R636 B.n305 B.n86 585
R637 B.n307 B.n306 585
R638 B.n308 B.n85 585
R639 B.n310 B.n309 585
R640 B.n311 B.n84 585
R641 B.n313 B.n312 585
R642 B.n314 B.n83 585
R643 B.n316 B.n315 585
R644 B.n317 B.n82 585
R645 B.n319 B.n318 585
R646 B.n320 B.n81 585
R647 B.n322 B.n321 585
R648 B.n323 B.n80 585
R649 B.n325 B.n324 585
R650 B.n326 B.n79 585
R651 B.n328 B.n327 585
R652 B.n329 B.n78 585
R653 B.n331 B.n330 585
R654 B.n332 B.n77 585
R655 B.n334 B.n333 585
R656 B.n335 B.n76 585
R657 B.n337 B.n336 585
R658 B.n338 B.n75 585
R659 B.n340 B.n339 585
R660 B.n341 B.n74 585
R661 B.n343 B.n342 585
R662 B.n344 B.n73 585
R663 B.n346 B.n345 585
R664 B.n347 B.n72 585
R665 B.n349 B.n348 585
R666 B.n350 B.n71 585
R667 B.n352 B.n351 585
R668 B.n353 B.n70 585
R669 B.n355 B.n354 585
R670 B.n356 B.n69 585
R671 B.n358 B.n357 585
R672 B.n359 B.n68 585
R673 B.n361 B.n360 585
R674 B.n362 B.n67 585
R675 B.n364 B.n363 585
R676 B.n365 B.n66 585
R677 B.n367 B.n366 585
R678 B.n368 B.n65 585
R679 B.n370 B.n369 585
R680 B.n371 B.n64 585
R681 B.n373 B.n372 585
R682 B.n374 B.n63 585
R683 B.n376 B.n375 585
R684 B.n377 B.n62 585
R685 B.n379 B.n378 585
R686 B.n380 B.n61 585
R687 B.n382 B.n381 585
R688 B.n383 B.n60 585
R689 B.n385 B.n384 585
R690 B.n386 B.n59 585
R691 B.n388 B.n387 585
R692 B.n389 B.n58 585
R693 B.n391 B.n390 585
R694 B.n392 B.n57 585
R695 B.n394 B.n393 585
R696 B.n395 B.n56 585
R697 B.n397 B.n396 585
R698 B.n491 B.n490 585
R699 B.n489 B.n20 585
R700 B.n488 B.n487 585
R701 B.n486 B.n21 585
R702 B.n485 B.n484 585
R703 B.n483 B.n22 585
R704 B.n482 B.n481 585
R705 B.n480 B.n23 585
R706 B.n479 B.n478 585
R707 B.n477 B.n24 585
R708 B.n476 B.n475 585
R709 B.n474 B.n25 585
R710 B.n473 B.n472 585
R711 B.n471 B.n26 585
R712 B.n470 B.n469 585
R713 B.n468 B.n27 585
R714 B.n467 B.n466 585
R715 B.n465 B.n28 585
R716 B.n464 B.n463 585
R717 B.n462 B.n29 585
R718 B.n461 B.n460 585
R719 B.n459 B.n30 585
R720 B.n458 B.n457 585
R721 B.n456 B.n31 585
R722 B.n455 B.n454 585
R723 B.n453 B.n32 585
R724 B.n452 B.n451 585
R725 B.n450 B.n33 585
R726 B.n449 B.n448 585
R727 B.n447 B.n37 585
R728 B.n446 B.n445 585
R729 B.n444 B.n38 585
R730 B.n443 B.n442 585
R731 B.n441 B.n39 585
R732 B.n440 B.n439 585
R733 B.n438 B.n40 585
R734 B.n436 B.n435 585
R735 B.n434 B.n43 585
R736 B.n433 B.n432 585
R737 B.n431 B.n44 585
R738 B.n430 B.n429 585
R739 B.n428 B.n45 585
R740 B.n427 B.n426 585
R741 B.n425 B.n46 585
R742 B.n424 B.n423 585
R743 B.n422 B.n47 585
R744 B.n421 B.n420 585
R745 B.n419 B.n48 585
R746 B.n418 B.n417 585
R747 B.n416 B.n49 585
R748 B.n415 B.n414 585
R749 B.n413 B.n50 585
R750 B.n412 B.n411 585
R751 B.n410 B.n51 585
R752 B.n409 B.n408 585
R753 B.n407 B.n52 585
R754 B.n406 B.n405 585
R755 B.n404 B.n53 585
R756 B.n403 B.n402 585
R757 B.n401 B.n54 585
R758 B.n400 B.n399 585
R759 B.n398 B.n55 585
R760 B.n492 B.n19 585
R761 B.n494 B.n493 585
R762 B.n495 B.n18 585
R763 B.n497 B.n496 585
R764 B.n498 B.n17 585
R765 B.n500 B.n499 585
R766 B.n501 B.n16 585
R767 B.n503 B.n502 585
R768 B.n504 B.n15 585
R769 B.n506 B.n505 585
R770 B.n507 B.n14 585
R771 B.n509 B.n508 585
R772 B.n510 B.n13 585
R773 B.n512 B.n511 585
R774 B.n513 B.n12 585
R775 B.n515 B.n514 585
R776 B.n516 B.n11 585
R777 B.n518 B.n517 585
R778 B.n519 B.n10 585
R779 B.n521 B.n520 585
R780 B.n522 B.n9 585
R781 B.n524 B.n523 585
R782 B.n525 B.n8 585
R783 B.n527 B.n526 585
R784 B.n528 B.n7 585
R785 B.n530 B.n529 585
R786 B.n531 B.n6 585
R787 B.n533 B.n532 585
R788 B.n534 B.n5 585
R789 B.n536 B.n535 585
R790 B.n537 B.n4 585
R791 B.n539 B.n538 585
R792 B.n540 B.n3 585
R793 B.n542 B.n541 585
R794 B.n543 B.n0 585
R795 B.n2 B.n1 585
R796 B.n142 B.n141 585
R797 B.n144 B.n143 585
R798 B.n145 B.n140 585
R799 B.n147 B.n146 585
R800 B.n148 B.n139 585
R801 B.n150 B.n149 585
R802 B.n151 B.n138 585
R803 B.n153 B.n152 585
R804 B.n154 B.n137 585
R805 B.n156 B.n155 585
R806 B.n157 B.n136 585
R807 B.n159 B.n158 585
R808 B.n160 B.n135 585
R809 B.n162 B.n161 585
R810 B.n163 B.n134 585
R811 B.n165 B.n164 585
R812 B.n166 B.n133 585
R813 B.n168 B.n167 585
R814 B.n169 B.n132 585
R815 B.n171 B.n170 585
R816 B.n172 B.n131 585
R817 B.n174 B.n173 585
R818 B.n175 B.n130 585
R819 B.n177 B.n176 585
R820 B.n178 B.n129 585
R821 B.n180 B.n179 585
R822 B.n181 B.n128 585
R823 B.n183 B.n182 585
R824 B.n184 B.n127 585
R825 B.n186 B.n185 585
R826 B.n187 B.n126 585
R827 B.n189 B.n188 585
R828 B.n190 B.n125 585
R829 B.n192 B.n191 585
R830 B.n191 B.n124 487.695
R831 B.n290 B.n289 487.695
R832 B.n398 B.n397 487.695
R833 B.n490 B.n19 487.695
R834 B.n105 B.t4 325.762
R835 B.n41 B.t11 325.762
R836 B.n230 B.t7 325.762
R837 B.n34 B.t2 325.762
R838 B.n230 B.t6 287.154
R839 B.n105 B.t3 287.154
R840 B.n41 B.t9 287.154
R841 B.n34 B.t0 287.154
R842 B.n106 B.t5 280.38
R843 B.n42 B.t10 280.38
R844 B.n231 B.t8 280.38
R845 B.n35 B.t1 280.38
R846 B.n545 B.n544 256.663
R847 B.n544 B.n543 235.042
R848 B.n544 B.n2 235.042
R849 B.n195 B.n124 163.367
R850 B.n196 B.n195 163.367
R851 B.n197 B.n196 163.367
R852 B.n197 B.n122 163.367
R853 B.n201 B.n122 163.367
R854 B.n202 B.n201 163.367
R855 B.n203 B.n202 163.367
R856 B.n203 B.n120 163.367
R857 B.n207 B.n120 163.367
R858 B.n208 B.n207 163.367
R859 B.n209 B.n208 163.367
R860 B.n209 B.n118 163.367
R861 B.n213 B.n118 163.367
R862 B.n214 B.n213 163.367
R863 B.n215 B.n214 163.367
R864 B.n215 B.n116 163.367
R865 B.n219 B.n116 163.367
R866 B.n220 B.n219 163.367
R867 B.n221 B.n220 163.367
R868 B.n221 B.n114 163.367
R869 B.n225 B.n114 163.367
R870 B.n226 B.n225 163.367
R871 B.n227 B.n226 163.367
R872 B.n227 B.n112 163.367
R873 B.n234 B.n112 163.367
R874 B.n235 B.n234 163.367
R875 B.n236 B.n235 163.367
R876 B.n236 B.n110 163.367
R877 B.n240 B.n110 163.367
R878 B.n241 B.n240 163.367
R879 B.n242 B.n241 163.367
R880 B.n242 B.n108 163.367
R881 B.n246 B.n108 163.367
R882 B.n247 B.n246 163.367
R883 B.n248 B.n247 163.367
R884 B.n248 B.n104 163.367
R885 B.n253 B.n104 163.367
R886 B.n254 B.n253 163.367
R887 B.n255 B.n254 163.367
R888 B.n255 B.n102 163.367
R889 B.n259 B.n102 163.367
R890 B.n260 B.n259 163.367
R891 B.n261 B.n260 163.367
R892 B.n261 B.n100 163.367
R893 B.n265 B.n100 163.367
R894 B.n266 B.n265 163.367
R895 B.n267 B.n266 163.367
R896 B.n267 B.n98 163.367
R897 B.n271 B.n98 163.367
R898 B.n272 B.n271 163.367
R899 B.n273 B.n272 163.367
R900 B.n273 B.n96 163.367
R901 B.n277 B.n96 163.367
R902 B.n278 B.n277 163.367
R903 B.n279 B.n278 163.367
R904 B.n279 B.n94 163.367
R905 B.n283 B.n94 163.367
R906 B.n284 B.n283 163.367
R907 B.n285 B.n284 163.367
R908 B.n285 B.n92 163.367
R909 B.n289 B.n92 163.367
R910 B.n397 B.n56 163.367
R911 B.n393 B.n56 163.367
R912 B.n393 B.n392 163.367
R913 B.n392 B.n391 163.367
R914 B.n391 B.n58 163.367
R915 B.n387 B.n58 163.367
R916 B.n387 B.n386 163.367
R917 B.n386 B.n385 163.367
R918 B.n385 B.n60 163.367
R919 B.n381 B.n60 163.367
R920 B.n381 B.n380 163.367
R921 B.n380 B.n379 163.367
R922 B.n379 B.n62 163.367
R923 B.n375 B.n62 163.367
R924 B.n375 B.n374 163.367
R925 B.n374 B.n373 163.367
R926 B.n373 B.n64 163.367
R927 B.n369 B.n64 163.367
R928 B.n369 B.n368 163.367
R929 B.n368 B.n367 163.367
R930 B.n367 B.n66 163.367
R931 B.n363 B.n66 163.367
R932 B.n363 B.n362 163.367
R933 B.n362 B.n361 163.367
R934 B.n361 B.n68 163.367
R935 B.n357 B.n68 163.367
R936 B.n357 B.n356 163.367
R937 B.n356 B.n355 163.367
R938 B.n355 B.n70 163.367
R939 B.n351 B.n70 163.367
R940 B.n351 B.n350 163.367
R941 B.n350 B.n349 163.367
R942 B.n349 B.n72 163.367
R943 B.n345 B.n72 163.367
R944 B.n345 B.n344 163.367
R945 B.n344 B.n343 163.367
R946 B.n343 B.n74 163.367
R947 B.n339 B.n74 163.367
R948 B.n339 B.n338 163.367
R949 B.n338 B.n337 163.367
R950 B.n337 B.n76 163.367
R951 B.n333 B.n76 163.367
R952 B.n333 B.n332 163.367
R953 B.n332 B.n331 163.367
R954 B.n331 B.n78 163.367
R955 B.n327 B.n78 163.367
R956 B.n327 B.n326 163.367
R957 B.n326 B.n325 163.367
R958 B.n325 B.n80 163.367
R959 B.n321 B.n80 163.367
R960 B.n321 B.n320 163.367
R961 B.n320 B.n319 163.367
R962 B.n319 B.n82 163.367
R963 B.n315 B.n82 163.367
R964 B.n315 B.n314 163.367
R965 B.n314 B.n313 163.367
R966 B.n313 B.n84 163.367
R967 B.n309 B.n84 163.367
R968 B.n309 B.n308 163.367
R969 B.n308 B.n307 163.367
R970 B.n307 B.n86 163.367
R971 B.n303 B.n86 163.367
R972 B.n303 B.n302 163.367
R973 B.n302 B.n301 163.367
R974 B.n301 B.n88 163.367
R975 B.n297 B.n88 163.367
R976 B.n297 B.n296 163.367
R977 B.n296 B.n295 163.367
R978 B.n295 B.n90 163.367
R979 B.n291 B.n90 163.367
R980 B.n291 B.n290 163.367
R981 B.n490 B.n489 163.367
R982 B.n489 B.n488 163.367
R983 B.n488 B.n21 163.367
R984 B.n484 B.n21 163.367
R985 B.n484 B.n483 163.367
R986 B.n483 B.n482 163.367
R987 B.n482 B.n23 163.367
R988 B.n478 B.n23 163.367
R989 B.n478 B.n477 163.367
R990 B.n477 B.n476 163.367
R991 B.n476 B.n25 163.367
R992 B.n472 B.n25 163.367
R993 B.n472 B.n471 163.367
R994 B.n471 B.n470 163.367
R995 B.n470 B.n27 163.367
R996 B.n466 B.n27 163.367
R997 B.n466 B.n465 163.367
R998 B.n465 B.n464 163.367
R999 B.n464 B.n29 163.367
R1000 B.n460 B.n29 163.367
R1001 B.n460 B.n459 163.367
R1002 B.n459 B.n458 163.367
R1003 B.n458 B.n31 163.367
R1004 B.n454 B.n31 163.367
R1005 B.n454 B.n453 163.367
R1006 B.n453 B.n452 163.367
R1007 B.n452 B.n33 163.367
R1008 B.n448 B.n33 163.367
R1009 B.n448 B.n447 163.367
R1010 B.n447 B.n446 163.367
R1011 B.n446 B.n38 163.367
R1012 B.n442 B.n38 163.367
R1013 B.n442 B.n441 163.367
R1014 B.n441 B.n440 163.367
R1015 B.n440 B.n40 163.367
R1016 B.n435 B.n40 163.367
R1017 B.n435 B.n434 163.367
R1018 B.n434 B.n433 163.367
R1019 B.n433 B.n44 163.367
R1020 B.n429 B.n44 163.367
R1021 B.n429 B.n428 163.367
R1022 B.n428 B.n427 163.367
R1023 B.n427 B.n46 163.367
R1024 B.n423 B.n46 163.367
R1025 B.n423 B.n422 163.367
R1026 B.n422 B.n421 163.367
R1027 B.n421 B.n48 163.367
R1028 B.n417 B.n48 163.367
R1029 B.n417 B.n416 163.367
R1030 B.n416 B.n415 163.367
R1031 B.n415 B.n50 163.367
R1032 B.n411 B.n50 163.367
R1033 B.n411 B.n410 163.367
R1034 B.n410 B.n409 163.367
R1035 B.n409 B.n52 163.367
R1036 B.n405 B.n52 163.367
R1037 B.n405 B.n404 163.367
R1038 B.n404 B.n403 163.367
R1039 B.n403 B.n54 163.367
R1040 B.n399 B.n54 163.367
R1041 B.n399 B.n398 163.367
R1042 B.n494 B.n19 163.367
R1043 B.n495 B.n494 163.367
R1044 B.n496 B.n495 163.367
R1045 B.n496 B.n17 163.367
R1046 B.n500 B.n17 163.367
R1047 B.n501 B.n500 163.367
R1048 B.n502 B.n501 163.367
R1049 B.n502 B.n15 163.367
R1050 B.n506 B.n15 163.367
R1051 B.n507 B.n506 163.367
R1052 B.n508 B.n507 163.367
R1053 B.n508 B.n13 163.367
R1054 B.n512 B.n13 163.367
R1055 B.n513 B.n512 163.367
R1056 B.n514 B.n513 163.367
R1057 B.n514 B.n11 163.367
R1058 B.n518 B.n11 163.367
R1059 B.n519 B.n518 163.367
R1060 B.n520 B.n519 163.367
R1061 B.n520 B.n9 163.367
R1062 B.n524 B.n9 163.367
R1063 B.n525 B.n524 163.367
R1064 B.n526 B.n525 163.367
R1065 B.n526 B.n7 163.367
R1066 B.n530 B.n7 163.367
R1067 B.n531 B.n530 163.367
R1068 B.n532 B.n531 163.367
R1069 B.n532 B.n5 163.367
R1070 B.n536 B.n5 163.367
R1071 B.n537 B.n536 163.367
R1072 B.n538 B.n537 163.367
R1073 B.n538 B.n3 163.367
R1074 B.n542 B.n3 163.367
R1075 B.n543 B.n542 163.367
R1076 B.n142 B.n2 163.367
R1077 B.n143 B.n142 163.367
R1078 B.n143 B.n140 163.367
R1079 B.n147 B.n140 163.367
R1080 B.n148 B.n147 163.367
R1081 B.n149 B.n148 163.367
R1082 B.n149 B.n138 163.367
R1083 B.n153 B.n138 163.367
R1084 B.n154 B.n153 163.367
R1085 B.n155 B.n154 163.367
R1086 B.n155 B.n136 163.367
R1087 B.n159 B.n136 163.367
R1088 B.n160 B.n159 163.367
R1089 B.n161 B.n160 163.367
R1090 B.n161 B.n134 163.367
R1091 B.n165 B.n134 163.367
R1092 B.n166 B.n165 163.367
R1093 B.n167 B.n166 163.367
R1094 B.n167 B.n132 163.367
R1095 B.n171 B.n132 163.367
R1096 B.n172 B.n171 163.367
R1097 B.n173 B.n172 163.367
R1098 B.n173 B.n130 163.367
R1099 B.n177 B.n130 163.367
R1100 B.n178 B.n177 163.367
R1101 B.n179 B.n178 163.367
R1102 B.n179 B.n128 163.367
R1103 B.n183 B.n128 163.367
R1104 B.n184 B.n183 163.367
R1105 B.n185 B.n184 163.367
R1106 B.n185 B.n126 163.367
R1107 B.n189 B.n126 163.367
R1108 B.n190 B.n189 163.367
R1109 B.n191 B.n190 163.367
R1110 B.n232 B.n231 59.5399
R1111 B.n250 B.n106 59.5399
R1112 B.n437 B.n42 59.5399
R1113 B.n36 B.n35 59.5399
R1114 B.n231 B.n230 45.3823
R1115 B.n106 B.n105 45.3823
R1116 B.n42 B.n41 45.3823
R1117 B.n35 B.n34 45.3823
R1118 B.n492 B.n491 31.6883
R1119 B.n396 B.n55 31.6883
R1120 B.n288 B.n91 31.6883
R1121 B.n193 B.n192 31.6883
R1122 B B.n545 18.0485
R1123 B.n493 B.n492 10.6151
R1124 B.n493 B.n18 10.6151
R1125 B.n497 B.n18 10.6151
R1126 B.n498 B.n497 10.6151
R1127 B.n499 B.n498 10.6151
R1128 B.n499 B.n16 10.6151
R1129 B.n503 B.n16 10.6151
R1130 B.n504 B.n503 10.6151
R1131 B.n505 B.n504 10.6151
R1132 B.n505 B.n14 10.6151
R1133 B.n509 B.n14 10.6151
R1134 B.n510 B.n509 10.6151
R1135 B.n511 B.n510 10.6151
R1136 B.n511 B.n12 10.6151
R1137 B.n515 B.n12 10.6151
R1138 B.n516 B.n515 10.6151
R1139 B.n517 B.n516 10.6151
R1140 B.n517 B.n10 10.6151
R1141 B.n521 B.n10 10.6151
R1142 B.n522 B.n521 10.6151
R1143 B.n523 B.n522 10.6151
R1144 B.n523 B.n8 10.6151
R1145 B.n527 B.n8 10.6151
R1146 B.n528 B.n527 10.6151
R1147 B.n529 B.n528 10.6151
R1148 B.n529 B.n6 10.6151
R1149 B.n533 B.n6 10.6151
R1150 B.n534 B.n533 10.6151
R1151 B.n535 B.n534 10.6151
R1152 B.n535 B.n4 10.6151
R1153 B.n539 B.n4 10.6151
R1154 B.n540 B.n539 10.6151
R1155 B.n541 B.n540 10.6151
R1156 B.n541 B.n0 10.6151
R1157 B.n491 B.n20 10.6151
R1158 B.n487 B.n20 10.6151
R1159 B.n487 B.n486 10.6151
R1160 B.n486 B.n485 10.6151
R1161 B.n485 B.n22 10.6151
R1162 B.n481 B.n22 10.6151
R1163 B.n481 B.n480 10.6151
R1164 B.n480 B.n479 10.6151
R1165 B.n479 B.n24 10.6151
R1166 B.n475 B.n24 10.6151
R1167 B.n475 B.n474 10.6151
R1168 B.n474 B.n473 10.6151
R1169 B.n473 B.n26 10.6151
R1170 B.n469 B.n26 10.6151
R1171 B.n469 B.n468 10.6151
R1172 B.n468 B.n467 10.6151
R1173 B.n467 B.n28 10.6151
R1174 B.n463 B.n28 10.6151
R1175 B.n463 B.n462 10.6151
R1176 B.n462 B.n461 10.6151
R1177 B.n461 B.n30 10.6151
R1178 B.n457 B.n30 10.6151
R1179 B.n457 B.n456 10.6151
R1180 B.n456 B.n455 10.6151
R1181 B.n455 B.n32 10.6151
R1182 B.n451 B.n450 10.6151
R1183 B.n450 B.n449 10.6151
R1184 B.n449 B.n37 10.6151
R1185 B.n445 B.n37 10.6151
R1186 B.n445 B.n444 10.6151
R1187 B.n444 B.n443 10.6151
R1188 B.n443 B.n39 10.6151
R1189 B.n439 B.n39 10.6151
R1190 B.n439 B.n438 10.6151
R1191 B.n436 B.n43 10.6151
R1192 B.n432 B.n43 10.6151
R1193 B.n432 B.n431 10.6151
R1194 B.n431 B.n430 10.6151
R1195 B.n430 B.n45 10.6151
R1196 B.n426 B.n45 10.6151
R1197 B.n426 B.n425 10.6151
R1198 B.n425 B.n424 10.6151
R1199 B.n424 B.n47 10.6151
R1200 B.n420 B.n47 10.6151
R1201 B.n420 B.n419 10.6151
R1202 B.n419 B.n418 10.6151
R1203 B.n418 B.n49 10.6151
R1204 B.n414 B.n49 10.6151
R1205 B.n414 B.n413 10.6151
R1206 B.n413 B.n412 10.6151
R1207 B.n412 B.n51 10.6151
R1208 B.n408 B.n51 10.6151
R1209 B.n408 B.n407 10.6151
R1210 B.n407 B.n406 10.6151
R1211 B.n406 B.n53 10.6151
R1212 B.n402 B.n53 10.6151
R1213 B.n402 B.n401 10.6151
R1214 B.n401 B.n400 10.6151
R1215 B.n400 B.n55 10.6151
R1216 B.n396 B.n395 10.6151
R1217 B.n395 B.n394 10.6151
R1218 B.n394 B.n57 10.6151
R1219 B.n390 B.n57 10.6151
R1220 B.n390 B.n389 10.6151
R1221 B.n389 B.n388 10.6151
R1222 B.n388 B.n59 10.6151
R1223 B.n384 B.n59 10.6151
R1224 B.n384 B.n383 10.6151
R1225 B.n383 B.n382 10.6151
R1226 B.n382 B.n61 10.6151
R1227 B.n378 B.n61 10.6151
R1228 B.n378 B.n377 10.6151
R1229 B.n377 B.n376 10.6151
R1230 B.n376 B.n63 10.6151
R1231 B.n372 B.n63 10.6151
R1232 B.n372 B.n371 10.6151
R1233 B.n371 B.n370 10.6151
R1234 B.n370 B.n65 10.6151
R1235 B.n366 B.n65 10.6151
R1236 B.n366 B.n365 10.6151
R1237 B.n365 B.n364 10.6151
R1238 B.n364 B.n67 10.6151
R1239 B.n360 B.n67 10.6151
R1240 B.n360 B.n359 10.6151
R1241 B.n359 B.n358 10.6151
R1242 B.n358 B.n69 10.6151
R1243 B.n354 B.n69 10.6151
R1244 B.n354 B.n353 10.6151
R1245 B.n353 B.n352 10.6151
R1246 B.n352 B.n71 10.6151
R1247 B.n348 B.n71 10.6151
R1248 B.n348 B.n347 10.6151
R1249 B.n347 B.n346 10.6151
R1250 B.n346 B.n73 10.6151
R1251 B.n342 B.n73 10.6151
R1252 B.n342 B.n341 10.6151
R1253 B.n341 B.n340 10.6151
R1254 B.n340 B.n75 10.6151
R1255 B.n336 B.n75 10.6151
R1256 B.n336 B.n335 10.6151
R1257 B.n335 B.n334 10.6151
R1258 B.n334 B.n77 10.6151
R1259 B.n330 B.n77 10.6151
R1260 B.n330 B.n329 10.6151
R1261 B.n329 B.n328 10.6151
R1262 B.n328 B.n79 10.6151
R1263 B.n324 B.n79 10.6151
R1264 B.n324 B.n323 10.6151
R1265 B.n323 B.n322 10.6151
R1266 B.n322 B.n81 10.6151
R1267 B.n318 B.n81 10.6151
R1268 B.n318 B.n317 10.6151
R1269 B.n317 B.n316 10.6151
R1270 B.n316 B.n83 10.6151
R1271 B.n312 B.n83 10.6151
R1272 B.n312 B.n311 10.6151
R1273 B.n311 B.n310 10.6151
R1274 B.n310 B.n85 10.6151
R1275 B.n306 B.n85 10.6151
R1276 B.n306 B.n305 10.6151
R1277 B.n305 B.n304 10.6151
R1278 B.n304 B.n87 10.6151
R1279 B.n300 B.n87 10.6151
R1280 B.n300 B.n299 10.6151
R1281 B.n299 B.n298 10.6151
R1282 B.n298 B.n89 10.6151
R1283 B.n294 B.n89 10.6151
R1284 B.n294 B.n293 10.6151
R1285 B.n293 B.n292 10.6151
R1286 B.n292 B.n91 10.6151
R1287 B.n141 B.n1 10.6151
R1288 B.n144 B.n141 10.6151
R1289 B.n145 B.n144 10.6151
R1290 B.n146 B.n145 10.6151
R1291 B.n146 B.n139 10.6151
R1292 B.n150 B.n139 10.6151
R1293 B.n151 B.n150 10.6151
R1294 B.n152 B.n151 10.6151
R1295 B.n152 B.n137 10.6151
R1296 B.n156 B.n137 10.6151
R1297 B.n157 B.n156 10.6151
R1298 B.n158 B.n157 10.6151
R1299 B.n158 B.n135 10.6151
R1300 B.n162 B.n135 10.6151
R1301 B.n163 B.n162 10.6151
R1302 B.n164 B.n163 10.6151
R1303 B.n164 B.n133 10.6151
R1304 B.n168 B.n133 10.6151
R1305 B.n169 B.n168 10.6151
R1306 B.n170 B.n169 10.6151
R1307 B.n170 B.n131 10.6151
R1308 B.n174 B.n131 10.6151
R1309 B.n175 B.n174 10.6151
R1310 B.n176 B.n175 10.6151
R1311 B.n176 B.n129 10.6151
R1312 B.n180 B.n129 10.6151
R1313 B.n181 B.n180 10.6151
R1314 B.n182 B.n181 10.6151
R1315 B.n182 B.n127 10.6151
R1316 B.n186 B.n127 10.6151
R1317 B.n187 B.n186 10.6151
R1318 B.n188 B.n187 10.6151
R1319 B.n188 B.n125 10.6151
R1320 B.n192 B.n125 10.6151
R1321 B.n194 B.n193 10.6151
R1322 B.n194 B.n123 10.6151
R1323 B.n198 B.n123 10.6151
R1324 B.n199 B.n198 10.6151
R1325 B.n200 B.n199 10.6151
R1326 B.n200 B.n121 10.6151
R1327 B.n204 B.n121 10.6151
R1328 B.n205 B.n204 10.6151
R1329 B.n206 B.n205 10.6151
R1330 B.n206 B.n119 10.6151
R1331 B.n210 B.n119 10.6151
R1332 B.n211 B.n210 10.6151
R1333 B.n212 B.n211 10.6151
R1334 B.n212 B.n117 10.6151
R1335 B.n216 B.n117 10.6151
R1336 B.n217 B.n216 10.6151
R1337 B.n218 B.n217 10.6151
R1338 B.n218 B.n115 10.6151
R1339 B.n222 B.n115 10.6151
R1340 B.n223 B.n222 10.6151
R1341 B.n224 B.n223 10.6151
R1342 B.n224 B.n113 10.6151
R1343 B.n228 B.n113 10.6151
R1344 B.n229 B.n228 10.6151
R1345 B.n233 B.n229 10.6151
R1346 B.n237 B.n111 10.6151
R1347 B.n238 B.n237 10.6151
R1348 B.n239 B.n238 10.6151
R1349 B.n239 B.n109 10.6151
R1350 B.n243 B.n109 10.6151
R1351 B.n244 B.n243 10.6151
R1352 B.n245 B.n244 10.6151
R1353 B.n245 B.n107 10.6151
R1354 B.n249 B.n107 10.6151
R1355 B.n252 B.n251 10.6151
R1356 B.n252 B.n103 10.6151
R1357 B.n256 B.n103 10.6151
R1358 B.n257 B.n256 10.6151
R1359 B.n258 B.n257 10.6151
R1360 B.n258 B.n101 10.6151
R1361 B.n262 B.n101 10.6151
R1362 B.n263 B.n262 10.6151
R1363 B.n264 B.n263 10.6151
R1364 B.n264 B.n99 10.6151
R1365 B.n268 B.n99 10.6151
R1366 B.n269 B.n268 10.6151
R1367 B.n270 B.n269 10.6151
R1368 B.n270 B.n97 10.6151
R1369 B.n274 B.n97 10.6151
R1370 B.n275 B.n274 10.6151
R1371 B.n276 B.n275 10.6151
R1372 B.n276 B.n95 10.6151
R1373 B.n280 B.n95 10.6151
R1374 B.n281 B.n280 10.6151
R1375 B.n282 B.n281 10.6151
R1376 B.n282 B.n93 10.6151
R1377 B.n286 B.n93 10.6151
R1378 B.n287 B.n286 10.6151
R1379 B.n288 B.n287 10.6151
R1380 B.n36 B.n32 9.36635
R1381 B.n437 B.n436 9.36635
R1382 B.n233 B.n232 9.36635
R1383 B.n251 B.n250 9.36635
R1384 B.n545 B.n0 8.11757
R1385 B.n545 B.n1 8.11757
R1386 B.n451 B.n36 1.24928
R1387 B.n438 B.n437 1.24928
R1388 B.n232 B.n111 1.24928
R1389 B.n250 B.n249 1.24928
C0 w_n2842_n2306# VDD2 1.84232f
C1 VP w_n2842_n2306# 5.51535f
C2 w_n2842_n2306# VDD1 1.77605f
C3 VDD2 B 1.58334f
C4 VP B 1.58651f
C5 VTAIL VDD2 5.64163f
C6 VP VTAIL 4.08427f
C7 VDD1 B 1.5234f
C8 VTAIL VDD1 5.59395f
C9 VN w_n2842_n2306# 5.14956f
C10 VP VDD2 0.407906f
C11 VN B 0.978763f
C12 VDD2 VDD1 1.1859f
C13 VN VTAIL 4.07003f
C14 VP VDD1 3.96777f
C15 VN VDD2 3.71215f
C16 VN VP 5.37369f
C17 w_n2842_n2306# B 7.37598f
C18 VN VDD1 0.150006f
C19 VTAIL w_n2842_n2306# 2.17569f
C20 VTAIL B 2.29971f
C21 VDD2 VSUBS 1.340137f
C22 VDD1 VSUBS 1.377849f
C23 VTAIL VSUBS 0.641323f
C24 VN VSUBS 4.99858f
C25 VP VSUBS 2.159117f
C26 B VSUBS 3.60392f
C27 w_n2842_n2306# VSUBS 81.6109f
C28 B.n0 VSUBS 0.006756f
C29 B.n1 VSUBS 0.006756f
C30 B.n2 VSUBS 0.009991f
C31 B.n3 VSUBS 0.007657f
C32 B.n4 VSUBS 0.007657f
C33 B.n5 VSUBS 0.007657f
C34 B.n6 VSUBS 0.007657f
C35 B.n7 VSUBS 0.007657f
C36 B.n8 VSUBS 0.007657f
C37 B.n9 VSUBS 0.007657f
C38 B.n10 VSUBS 0.007657f
C39 B.n11 VSUBS 0.007657f
C40 B.n12 VSUBS 0.007657f
C41 B.n13 VSUBS 0.007657f
C42 B.n14 VSUBS 0.007657f
C43 B.n15 VSUBS 0.007657f
C44 B.n16 VSUBS 0.007657f
C45 B.n17 VSUBS 0.007657f
C46 B.n18 VSUBS 0.007657f
C47 B.n19 VSUBS 0.016849f
C48 B.n20 VSUBS 0.007657f
C49 B.n21 VSUBS 0.007657f
C50 B.n22 VSUBS 0.007657f
C51 B.n23 VSUBS 0.007657f
C52 B.n24 VSUBS 0.007657f
C53 B.n25 VSUBS 0.007657f
C54 B.n26 VSUBS 0.007657f
C55 B.n27 VSUBS 0.007657f
C56 B.n28 VSUBS 0.007657f
C57 B.n29 VSUBS 0.007657f
C58 B.n30 VSUBS 0.007657f
C59 B.n31 VSUBS 0.007657f
C60 B.n32 VSUBS 0.007206f
C61 B.n33 VSUBS 0.007657f
C62 B.t1 VSUBS 0.111394f
C63 B.t2 VSUBS 0.135257f
C64 B.t0 VSUBS 0.682098f
C65 B.n34 VSUBS 0.231088f
C66 B.n35 VSUBS 0.182214f
C67 B.n36 VSUBS 0.017739f
C68 B.n37 VSUBS 0.007657f
C69 B.n38 VSUBS 0.007657f
C70 B.n39 VSUBS 0.007657f
C71 B.n40 VSUBS 0.007657f
C72 B.t10 VSUBS 0.111396f
C73 B.t11 VSUBS 0.135258f
C74 B.t9 VSUBS 0.682098f
C75 B.n41 VSUBS 0.231086f
C76 B.n42 VSUBS 0.182211f
C77 B.n43 VSUBS 0.007657f
C78 B.n44 VSUBS 0.007657f
C79 B.n45 VSUBS 0.007657f
C80 B.n46 VSUBS 0.007657f
C81 B.n47 VSUBS 0.007657f
C82 B.n48 VSUBS 0.007657f
C83 B.n49 VSUBS 0.007657f
C84 B.n50 VSUBS 0.007657f
C85 B.n51 VSUBS 0.007657f
C86 B.n52 VSUBS 0.007657f
C87 B.n53 VSUBS 0.007657f
C88 B.n54 VSUBS 0.007657f
C89 B.n55 VSUBS 0.018281f
C90 B.n56 VSUBS 0.007657f
C91 B.n57 VSUBS 0.007657f
C92 B.n58 VSUBS 0.007657f
C93 B.n59 VSUBS 0.007657f
C94 B.n60 VSUBS 0.007657f
C95 B.n61 VSUBS 0.007657f
C96 B.n62 VSUBS 0.007657f
C97 B.n63 VSUBS 0.007657f
C98 B.n64 VSUBS 0.007657f
C99 B.n65 VSUBS 0.007657f
C100 B.n66 VSUBS 0.007657f
C101 B.n67 VSUBS 0.007657f
C102 B.n68 VSUBS 0.007657f
C103 B.n69 VSUBS 0.007657f
C104 B.n70 VSUBS 0.007657f
C105 B.n71 VSUBS 0.007657f
C106 B.n72 VSUBS 0.007657f
C107 B.n73 VSUBS 0.007657f
C108 B.n74 VSUBS 0.007657f
C109 B.n75 VSUBS 0.007657f
C110 B.n76 VSUBS 0.007657f
C111 B.n77 VSUBS 0.007657f
C112 B.n78 VSUBS 0.007657f
C113 B.n79 VSUBS 0.007657f
C114 B.n80 VSUBS 0.007657f
C115 B.n81 VSUBS 0.007657f
C116 B.n82 VSUBS 0.007657f
C117 B.n83 VSUBS 0.007657f
C118 B.n84 VSUBS 0.007657f
C119 B.n85 VSUBS 0.007657f
C120 B.n86 VSUBS 0.007657f
C121 B.n87 VSUBS 0.007657f
C122 B.n88 VSUBS 0.007657f
C123 B.n89 VSUBS 0.007657f
C124 B.n90 VSUBS 0.007657f
C125 B.n91 VSUBS 0.017781f
C126 B.n92 VSUBS 0.007657f
C127 B.n93 VSUBS 0.007657f
C128 B.n94 VSUBS 0.007657f
C129 B.n95 VSUBS 0.007657f
C130 B.n96 VSUBS 0.007657f
C131 B.n97 VSUBS 0.007657f
C132 B.n98 VSUBS 0.007657f
C133 B.n99 VSUBS 0.007657f
C134 B.n100 VSUBS 0.007657f
C135 B.n101 VSUBS 0.007657f
C136 B.n102 VSUBS 0.007657f
C137 B.n103 VSUBS 0.007657f
C138 B.n104 VSUBS 0.007657f
C139 B.t5 VSUBS 0.111396f
C140 B.t4 VSUBS 0.135258f
C141 B.t3 VSUBS 0.682098f
C142 B.n105 VSUBS 0.231086f
C143 B.n106 VSUBS 0.182211f
C144 B.n107 VSUBS 0.007657f
C145 B.n108 VSUBS 0.007657f
C146 B.n109 VSUBS 0.007657f
C147 B.n110 VSUBS 0.007657f
C148 B.n111 VSUBS 0.004279f
C149 B.n112 VSUBS 0.007657f
C150 B.n113 VSUBS 0.007657f
C151 B.n114 VSUBS 0.007657f
C152 B.n115 VSUBS 0.007657f
C153 B.n116 VSUBS 0.007657f
C154 B.n117 VSUBS 0.007657f
C155 B.n118 VSUBS 0.007657f
C156 B.n119 VSUBS 0.007657f
C157 B.n120 VSUBS 0.007657f
C158 B.n121 VSUBS 0.007657f
C159 B.n122 VSUBS 0.007657f
C160 B.n123 VSUBS 0.007657f
C161 B.n124 VSUBS 0.018281f
C162 B.n125 VSUBS 0.007657f
C163 B.n126 VSUBS 0.007657f
C164 B.n127 VSUBS 0.007657f
C165 B.n128 VSUBS 0.007657f
C166 B.n129 VSUBS 0.007657f
C167 B.n130 VSUBS 0.007657f
C168 B.n131 VSUBS 0.007657f
C169 B.n132 VSUBS 0.007657f
C170 B.n133 VSUBS 0.007657f
C171 B.n134 VSUBS 0.007657f
C172 B.n135 VSUBS 0.007657f
C173 B.n136 VSUBS 0.007657f
C174 B.n137 VSUBS 0.007657f
C175 B.n138 VSUBS 0.007657f
C176 B.n139 VSUBS 0.007657f
C177 B.n140 VSUBS 0.007657f
C178 B.n141 VSUBS 0.007657f
C179 B.n142 VSUBS 0.007657f
C180 B.n143 VSUBS 0.007657f
C181 B.n144 VSUBS 0.007657f
C182 B.n145 VSUBS 0.007657f
C183 B.n146 VSUBS 0.007657f
C184 B.n147 VSUBS 0.007657f
C185 B.n148 VSUBS 0.007657f
C186 B.n149 VSUBS 0.007657f
C187 B.n150 VSUBS 0.007657f
C188 B.n151 VSUBS 0.007657f
C189 B.n152 VSUBS 0.007657f
C190 B.n153 VSUBS 0.007657f
C191 B.n154 VSUBS 0.007657f
C192 B.n155 VSUBS 0.007657f
C193 B.n156 VSUBS 0.007657f
C194 B.n157 VSUBS 0.007657f
C195 B.n158 VSUBS 0.007657f
C196 B.n159 VSUBS 0.007657f
C197 B.n160 VSUBS 0.007657f
C198 B.n161 VSUBS 0.007657f
C199 B.n162 VSUBS 0.007657f
C200 B.n163 VSUBS 0.007657f
C201 B.n164 VSUBS 0.007657f
C202 B.n165 VSUBS 0.007657f
C203 B.n166 VSUBS 0.007657f
C204 B.n167 VSUBS 0.007657f
C205 B.n168 VSUBS 0.007657f
C206 B.n169 VSUBS 0.007657f
C207 B.n170 VSUBS 0.007657f
C208 B.n171 VSUBS 0.007657f
C209 B.n172 VSUBS 0.007657f
C210 B.n173 VSUBS 0.007657f
C211 B.n174 VSUBS 0.007657f
C212 B.n175 VSUBS 0.007657f
C213 B.n176 VSUBS 0.007657f
C214 B.n177 VSUBS 0.007657f
C215 B.n178 VSUBS 0.007657f
C216 B.n179 VSUBS 0.007657f
C217 B.n180 VSUBS 0.007657f
C218 B.n181 VSUBS 0.007657f
C219 B.n182 VSUBS 0.007657f
C220 B.n183 VSUBS 0.007657f
C221 B.n184 VSUBS 0.007657f
C222 B.n185 VSUBS 0.007657f
C223 B.n186 VSUBS 0.007657f
C224 B.n187 VSUBS 0.007657f
C225 B.n188 VSUBS 0.007657f
C226 B.n189 VSUBS 0.007657f
C227 B.n190 VSUBS 0.007657f
C228 B.n191 VSUBS 0.016849f
C229 B.n192 VSUBS 0.016849f
C230 B.n193 VSUBS 0.018281f
C231 B.n194 VSUBS 0.007657f
C232 B.n195 VSUBS 0.007657f
C233 B.n196 VSUBS 0.007657f
C234 B.n197 VSUBS 0.007657f
C235 B.n198 VSUBS 0.007657f
C236 B.n199 VSUBS 0.007657f
C237 B.n200 VSUBS 0.007657f
C238 B.n201 VSUBS 0.007657f
C239 B.n202 VSUBS 0.007657f
C240 B.n203 VSUBS 0.007657f
C241 B.n204 VSUBS 0.007657f
C242 B.n205 VSUBS 0.007657f
C243 B.n206 VSUBS 0.007657f
C244 B.n207 VSUBS 0.007657f
C245 B.n208 VSUBS 0.007657f
C246 B.n209 VSUBS 0.007657f
C247 B.n210 VSUBS 0.007657f
C248 B.n211 VSUBS 0.007657f
C249 B.n212 VSUBS 0.007657f
C250 B.n213 VSUBS 0.007657f
C251 B.n214 VSUBS 0.007657f
C252 B.n215 VSUBS 0.007657f
C253 B.n216 VSUBS 0.007657f
C254 B.n217 VSUBS 0.007657f
C255 B.n218 VSUBS 0.007657f
C256 B.n219 VSUBS 0.007657f
C257 B.n220 VSUBS 0.007657f
C258 B.n221 VSUBS 0.007657f
C259 B.n222 VSUBS 0.007657f
C260 B.n223 VSUBS 0.007657f
C261 B.n224 VSUBS 0.007657f
C262 B.n225 VSUBS 0.007657f
C263 B.n226 VSUBS 0.007657f
C264 B.n227 VSUBS 0.007657f
C265 B.n228 VSUBS 0.007657f
C266 B.n229 VSUBS 0.007657f
C267 B.t8 VSUBS 0.111394f
C268 B.t7 VSUBS 0.135257f
C269 B.t6 VSUBS 0.682098f
C270 B.n230 VSUBS 0.231088f
C271 B.n231 VSUBS 0.182214f
C272 B.n232 VSUBS 0.017739f
C273 B.n233 VSUBS 0.007206f
C274 B.n234 VSUBS 0.007657f
C275 B.n235 VSUBS 0.007657f
C276 B.n236 VSUBS 0.007657f
C277 B.n237 VSUBS 0.007657f
C278 B.n238 VSUBS 0.007657f
C279 B.n239 VSUBS 0.007657f
C280 B.n240 VSUBS 0.007657f
C281 B.n241 VSUBS 0.007657f
C282 B.n242 VSUBS 0.007657f
C283 B.n243 VSUBS 0.007657f
C284 B.n244 VSUBS 0.007657f
C285 B.n245 VSUBS 0.007657f
C286 B.n246 VSUBS 0.007657f
C287 B.n247 VSUBS 0.007657f
C288 B.n248 VSUBS 0.007657f
C289 B.n249 VSUBS 0.004279f
C290 B.n250 VSUBS 0.017739f
C291 B.n251 VSUBS 0.007206f
C292 B.n252 VSUBS 0.007657f
C293 B.n253 VSUBS 0.007657f
C294 B.n254 VSUBS 0.007657f
C295 B.n255 VSUBS 0.007657f
C296 B.n256 VSUBS 0.007657f
C297 B.n257 VSUBS 0.007657f
C298 B.n258 VSUBS 0.007657f
C299 B.n259 VSUBS 0.007657f
C300 B.n260 VSUBS 0.007657f
C301 B.n261 VSUBS 0.007657f
C302 B.n262 VSUBS 0.007657f
C303 B.n263 VSUBS 0.007657f
C304 B.n264 VSUBS 0.007657f
C305 B.n265 VSUBS 0.007657f
C306 B.n266 VSUBS 0.007657f
C307 B.n267 VSUBS 0.007657f
C308 B.n268 VSUBS 0.007657f
C309 B.n269 VSUBS 0.007657f
C310 B.n270 VSUBS 0.007657f
C311 B.n271 VSUBS 0.007657f
C312 B.n272 VSUBS 0.007657f
C313 B.n273 VSUBS 0.007657f
C314 B.n274 VSUBS 0.007657f
C315 B.n275 VSUBS 0.007657f
C316 B.n276 VSUBS 0.007657f
C317 B.n277 VSUBS 0.007657f
C318 B.n278 VSUBS 0.007657f
C319 B.n279 VSUBS 0.007657f
C320 B.n280 VSUBS 0.007657f
C321 B.n281 VSUBS 0.007657f
C322 B.n282 VSUBS 0.007657f
C323 B.n283 VSUBS 0.007657f
C324 B.n284 VSUBS 0.007657f
C325 B.n285 VSUBS 0.007657f
C326 B.n286 VSUBS 0.007657f
C327 B.n287 VSUBS 0.007657f
C328 B.n288 VSUBS 0.017349f
C329 B.n289 VSUBS 0.018281f
C330 B.n290 VSUBS 0.016849f
C331 B.n291 VSUBS 0.007657f
C332 B.n292 VSUBS 0.007657f
C333 B.n293 VSUBS 0.007657f
C334 B.n294 VSUBS 0.007657f
C335 B.n295 VSUBS 0.007657f
C336 B.n296 VSUBS 0.007657f
C337 B.n297 VSUBS 0.007657f
C338 B.n298 VSUBS 0.007657f
C339 B.n299 VSUBS 0.007657f
C340 B.n300 VSUBS 0.007657f
C341 B.n301 VSUBS 0.007657f
C342 B.n302 VSUBS 0.007657f
C343 B.n303 VSUBS 0.007657f
C344 B.n304 VSUBS 0.007657f
C345 B.n305 VSUBS 0.007657f
C346 B.n306 VSUBS 0.007657f
C347 B.n307 VSUBS 0.007657f
C348 B.n308 VSUBS 0.007657f
C349 B.n309 VSUBS 0.007657f
C350 B.n310 VSUBS 0.007657f
C351 B.n311 VSUBS 0.007657f
C352 B.n312 VSUBS 0.007657f
C353 B.n313 VSUBS 0.007657f
C354 B.n314 VSUBS 0.007657f
C355 B.n315 VSUBS 0.007657f
C356 B.n316 VSUBS 0.007657f
C357 B.n317 VSUBS 0.007657f
C358 B.n318 VSUBS 0.007657f
C359 B.n319 VSUBS 0.007657f
C360 B.n320 VSUBS 0.007657f
C361 B.n321 VSUBS 0.007657f
C362 B.n322 VSUBS 0.007657f
C363 B.n323 VSUBS 0.007657f
C364 B.n324 VSUBS 0.007657f
C365 B.n325 VSUBS 0.007657f
C366 B.n326 VSUBS 0.007657f
C367 B.n327 VSUBS 0.007657f
C368 B.n328 VSUBS 0.007657f
C369 B.n329 VSUBS 0.007657f
C370 B.n330 VSUBS 0.007657f
C371 B.n331 VSUBS 0.007657f
C372 B.n332 VSUBS 0.007657f
C373 B.n333 VSUBS 0.007657f
C374 B.n334 VSUBS 0.007657f
C375 B.n335 VSUBS 0.007657f
C376 B.n336 VSUBS 0.007657f
C377 B.n337 VSUBS 0.007657f
C378 B.n338 VSUBS 0.007657f
C379 B.n339 VSUBS 0.007657f
C380 B.n340 VSUBS 0.007657f
C381 B.n341 VSUBS 0.007657f
C382 B.n342 VSUBS 0.007657f
C383 B.n343 VSUBS 0.007657f
C384 B.n344 VSUBS 0.007657f
C385 B.n345 VSUBS 0.007657f
C386 B.n346 VSUBS 0.007657f
C387 B.n347 VSUBS 0.007657f
C388 B.n348 VSUBS 0.007657f
C389 B.n349 VSUBS 0.007657f
C390 B.n350 VSUBS 0.007657f
C391 B.n351 VSUBS 0.007657f
C392 B.n352 VSUBS 0.007657f
C393 B.n353 VSUBS 0.007657f
C394 B.n354 VSUBS 0.007657f
C395 B.n355 VSUBS 0.007657f
C396 B.n356 VSUBS 0.007657f
C397 B.n357 VSUBS 0.007657f
C398 B.n358 VSUBS 0.007657f
C399 B.n359 VSUBS 0.007657f
C400 B.n360 VSUBS 0.007657f
C401 B.n361 VSUBS 0.007657f
C402 B.n362 VSUBS 0.007657f
C403 B.n363 VSUBS 0.007657f
C404 B.n364 VSUBS 0.007657f
C405 B.n365 VSUBS 0.007657f
C406 B.n366 VSUBS 0.007657f
C407 B.n367 VSUBS 0.007657f
C408 B.n368 VSUBS 0.007657f
C409 B.n369 VSUBS 0.007657f
C410 B.n370 VSUBS 0.007657f
C411 B.n371 VSUBS 0.007657f
C412 B.n372 VSUBS 0.007657f
C413 B.n373 VSUBS 0.007657f
C414 B.n374 VSUBS 0.007657f
C415 B.n375 VSUBS 0.007657f
C416 B.n376 VSUBS 0.007657f
C417 B.n377 VSUBS 0.007657f
C418 B.n378 VSUBS 0.007657f
C419 B.n379 VSUBS 0.007657f
C420 B.n380 VSUBS 0.007657f
C421 B.n381 VSUBS 0.007657f
C422 B.n382 VSUBS 0.007657f
C423 B.n383 VSUBS 0.007657f
C424 B.n384 VSUBS 0.007657f
C425 B.n385 VSUBS 0.007657f
C426 B.n386 VSUBS 0.007657f
C427 B.n387 VSUBS 0.007657f
C428 B.n388 VSUBS 0.007657f
C429 B.n389 VSUBS 0.007657f
C430 B.n390 VSUBS 0.007657f
C431 B.n391 VSUBS 0.007657f
C432 B.n392 VSUBS 0.007657f
C433 B.n393 VSUBS 0.007657f
C434 B.n394 VSUBS 0.007657f
C435 B.n395 VSUBS 0.007657f
C436 B.n396 VSUBS 0.016849f
C437 B.n397 VSUBS 0.016849f
C438 B.n398 VSUBS 0.018281f
C439 B.n399 VSUBS 0.007657f
C440 B.n400 VSUBS 0.007657f
C441 B.n401 VSUBS 0.007657f
C442 B.n402 VSUBS 0.007657f
C443 B.n403 VSUBS 0.007657f
C444 B.n404 VSUBS 0.007657f
C445 B.n405 VSUBS 0.007657f
C446 B.n406 VSUBS 0.007657f
C447 B.n407 VSUBS 0.007657f
C448 B.n408 VSUBS 0.007657f
C449 B.n409 VSUBS 0.007657f
C450 B.n410 VSUBS 0.007657f
C451 B.n411 VSUBS 0.007657f
C452 B.n412 VSUBS 0.007657f
C453 B.n413 VSUBS 0.007657f
C454 B.n414 VSUBS 0.007657f
C455 B.n415 VSUBS 0.007657f
C456 B.n416 VSUBS 0.007657f
C457 B.n417 VSUBS 0.007657f
C458 B.n418 VSUBS 0.007657f
C459 B.n419 VSUBS 0.007657f
C460 B.n420 VSUBS 0.007657f
C461 B.n421 VSUBS 0.007657f
C462 B.n422 VSUBS 0.007657f
C463 B.n423 VSUBS 0.007657f
C464 B.n424 VSUBS 0.007657f
C465 B.n425 VSUBS 0.007657f
C466 B.n426 VSUBS 0.007657f
C467 B.n427 VSUBS 0.007657f
C468 B.n428 VSUBS 0.007657f
C469 B.n429 VSUBS 0.007657f
C470 B.n430 VSUBS 0.007657f
C471 B.n431 VSUBS 0.007657f
C472 B.n432 VSUBS 0.007657f
C473 B.n433 VSUBS 0.007657f
C474 B.n434 VSUBS 0.007657f
C475 B.n435 VSUBS 0.007657f
C476 B.n436 VSUBS 0.007206f
C477 B.n437 VSUBS 0.017739f
C478 B.n438 VSUBS 0.004279f
C479 B.n439 VSUBS 0.007657f
C480 B.n440 VSUBS 0.007657f
C481 B.n441 VSUBS 0.007657f
C482 B.n442 VSUBS 0.007657f
C483 B.n443 VSUBS 0.007657f
C484 B.n444 VSUBS 0.007657f
C485 B.n445 VSUBS 0.007657f
C486 B.n446 VSUBS 0.007657f
C487 B.n447 VSUBS 0.007657f
C488 B.n448 VSUBS 0.007657f
C489 B.n449 VSUBS 0.007657f
C490 B.n450 VSUBS 0.007657f
C491 B.n451 VSUBS 0.004279f
C492 B.n452 VSUBS 0.007657f
C493 B.n453 VSUBS 0.007657f
C494 B.n454 VSUBS 0.007657f
C495 B.n455 VSUBS 0.007657f
C496 B.n456 VSUBS 0.007657f
C497 B.n457 VSUBS 0.007657f
C498 B.n458 VSUBS 0.007657f
C499 B.n459 VSUBS 0.007657f
C500 B.n460 VSUBS 0.007657f
C501 B.n461 VSUBS 0.007657f
C502 B.n462 VSUBS 0.007657f
C503 B.n463 VSUBS 0.007657f
C504 B.n464 VSUBS 0.007657f
C505 B.n465 VSUBS 0.007657f
C506 B.n466 VSUBS 0.007657f
C507 B.n467 VSUBS 0.007657f
C508 B.n468 VSUBS 0.007657f
C509 B.n469 VSUBS 0.007657f
C510 B.n470 VSUBS 0.007657f
C511 B.n471 VSUBS 0.007657f
C512 B.n472 VSUBS 0.007657f
C513 B.n473 VSUBS 0.007657f
C514 B.n474 VSUBS 0.007657f
C515 B.n475 VSUBS 0.007657f
C516 B.n476 VSUBS 0.007657f
C517 B.n477 VSUBS 0.007657f
C518 B.n478 VSUBS 0.007657f
C519 B.n479 VSUBS 0.007657f
C520 B.n480 VSUBS 0.007657f
C521 B.n481 VSUBS 0.007657f
C522 B.n482 VSUBS 0.007657f
C523 B.n483 VSUBS 0.007657f
C524 B.n484 VSUBS 0.007657f
C525 B.n485 VSUBS 0.007657f
C526 B.n486 VSUBS 0.007657f
C527 B.n487 VSUBS 0.007657f
C528 B.n488 VSUBS 0.007657f
C529 B.n489 VSUBS 0.007657f
C530 B.n490 VSUBS 0.018281f
C531 B.n491 VSUBS 0.018281f
C532 B.n492 VSUBS 0.016849f
C533 B.n493 VSUBS 0.007657f
C534 B.n494 VSUBS 0.007657f
C535 B.n495 VSUBS 0.007657f
C536 B.n496 VSUBS 0.007657f
C537 B.n497 VSUBS 0.007657f
C538 B.n498 VSUBS 0.007657f
C539 B.n499 VSUBS 0.007657f
C540 B.n500 VSUBS 0.007657f
C541 B.n501 VSUBS 0.007657f
C542 B.n502 VSUBS 0.007657f
C543 B.n503 VSUBS 0.007657f
C544 B.n504 VSUBS 0.007657f
C545 B.n505 VSUBS 0.007657f
C546 B.n506 VSUBS 0.007657f
C547 B.n507 VSUBS 0.007657f
C548 B.n508 VSUBS 0.007657f
C549 B.n509 VSUBS 0.007657f
C550 B.n510 VSUBS 0.007657f
C551 B.n511 VSUBS 0.007657f
C552 B.n512 VSUBS 0.007657f
C553 B.n513 VSUBS 0.007657f
C554 B.n514 VSUBS 0.007657f
C555 B.n515 VSUBS 0.007657f
C556 B.n516 VSUBS 0.007657f
C557 B.n517 VSUBS 0.007657f
C558 B.n518 VSUBS 0.007657f
C559 B.n519 VSUBS 0.007657f
C560 B.n520 VSUBS 0.007657f
C561 B.n521 VSUBS 0.007657f
C562 B.n522 VSUBS 0.007657f
C563 B.n523 VSUBS 0.007657f
C564 B.n524 VSUBS 0.007657f
C565 B.n525 VSUBS 0.007657f
C566 B.n526 VSUBS 0.007657f
C567 B.n527 VSUBS 0.007657f
C568 B.n528 VSUBS 0.007657f
C569 B.n529 VSUBS 0.007657f
C570 B.n530 VSUBS 0.007657f
C571 B.n531 VSUBS 0.007657f
C572 B.n532 VSUBS 0.007657f
C573 B.n533 VSUBS 0.007657f
C574 B.n534 VSUBS 0.007657f
C575 B.n535 VSUBS 0.007657f
C576 B.n536 VSUBS 0.007657f
C577 B.n537 VSUBS 0.007657f
C578 B.n538 VSUBS 0.007657f
C579 B.n539 VSUBS 0.007657f
C580 B.n540 VSUBS 0.007657f
C581 B.n541 VSUBS 0.007657f
C582 B.n542 VSUBS 0.007657f
C583 B.n543 VSUBS 0.009991f
C584 B.n544 VSUBS 0.010643f
C585 B.n545 VSUBS 0.021165f
C586 VDD2.n0 VSUBS 0.023839f
C587 VDD2.n1 VSUBS 0.021695f
C588 VDD2.n2 VSUBS 0.011658f
C589 VDD2.n3 VSUBS 0.027555f
C590 VDD2.n4 VSUBS 0.012344f
C591 VDD2.n5 VSUBS 0.021695f
C592 VDD2.n6 VSUBS 0.011658f
C593 VDD2.n7 VSUBS 0.027555f
C594 VDD2.n8 VSUBS 0.012344f
C595 VDD2.n9 VSUBS 0.566085f
C596 VDD2.n10 VSUBS 0.011658f
C597 VDD2.t3 VSUBS 0.05892f
C598 VDD2.n11 VSUBS 0.100119f
C599 VDD2.n12 VSUBS 0.017526f
C600 VDD2.n13 VSUBS 0.020666f
C601 VDD2.n14 VSUBS 0.027555f
C602 VDD2.n15 VSUBS 0.012344f
C603 VDD2.n16 VSUBS 0.011658f
C604 VDD2.n17 VSUBS 0.021695f
C605 VDD2.n18 VSUBS 0.021695f
C606 VDD2.n19 VSUBS 0.011658f
C607 VDD2.n20 VSUBS 0.012344f
C608 VDD2.n21 VSUBS 0.027555f
C609 VDD2.n22 VSUBS 0.027555f
C610 VDD2.n23 VSUBS 0.012344f
C611 VDD2.n24 VSUBS 0.011658f
C612 VDD2.n25 VSUBS 0.021695f
C613 VDD2.n26 VSUBS 0.021695f
C614 VDD2.n27 VSUBS 0.011658f
C615 VDD2.n28 VSUBS 0.012344f
C616 VDD2.n29 VSUBS 0.027555f
C617 VDD2.n30 VSUBS 0.066712f
C618 VDD2.n31 VSUBS 0.012344f
C619 VDD2.n32 VSUBS 0.011658f
C620 VDD2.n33 VSUBS 0.049258f
C621 VDD2.n34 VSUBS 0.052714f
C622 VDD2.t5 VSUBS 0.114694f
C623 VDD2.t0 VSUBS 0.114694f
C624 VDD2.n35 VSUBS 0.784298f
C625 VDD2.n36 VSUBS 2.00984f
C626 VDD2.n37 VSUBS 0.023839f
C627 VDD2.n38 VSUBS 0.021695f
C628 VDD2.n39 VSUBS 0.011658f
C629 VDD2.n40 VSUBS 0.027555f
C630 VDD2.n41 VSUBS 0.012344f
C631 VDD2.n42 VSUBS 0.021695f
C632 VDD2.n43 VSUBS 0.011658f
C633 VDD2.n44 VSUBS 0.027555f
C634 VDD2.n45 VSUBS 0.012344f
C635 VDD2.n46 VSUBS 0.566085f
C636 VDD2.n47 VSUBS 0.011658f
C637 VDD2.t4 VSUBS 0.05892f
C638 VDD2.n48 VSUBS 0.100119f
C639 VDD2.n49 VSUBS 0.017526f
C640 VDD2.n50 VSUBS 0.020666f
C641 VDD2.n51 VSUBS 0.027555f
C642 VDD2.n52 VSUBS 0.012344f
C643 VDD2.n53 VSUBS 0.011658f
C644 VDD2.n54 VSUBS 0.021695f
C645 VDD2.n55 VSUBS 0.021695f
C646 VDD2.n56 VSUBS 0.011658f
C647 VDD2.n57 VSUBS 0.012344f
C648 VDD2.n58 VSUBS 0.027555f
C649 VDD2.n59 VSUBS 0.027555f
C650 VDD2.n60 VSUBS 0.012344f
C651 VDD2.n61 VSUBS 0.011658f
C652 VDD2.n62 VSUBS 0.021695f
C653 VDD2.n63 VSUBS 0.021695f
C654 VDD2.n64 VSUBS 0.011658f
C655 VDD2.n65 VSUBS 0.012344f
C656 VDD2.n66 VSUBS 0.027555f
C657 VDD2.n67 VSUBS 0.066712f
C658 VDD2.n68 VSUBS 0.012344f
C659 VDD2.n69 VSUBS 0.011658f
C660 VDD2.n70 VSUBS 0.049258f
C661 VDD2.n71 VSUBS 0.048509f
C662 VDD2.n72 VSUBS 1.72078f
C663 VDD2.t2 VSUBS 0.114694f
C664 VDD2.t1 VSUBS 0.114694f
C665 VDD2.n73 VSUBS 0.784274f
C666 VN.n0 VSUBS 0.054065f
C667 VN.t5 VSUBS 1.46836f
C668 VN.n1 VSUBS 0.050722f
C669 VN.t2 VSUBS 1.6932f
C670 VN.n2 VSUBS 0.639934f
C671 VN.t0 VSUBS 1.46836f
C672 VN.n3 VSUBS 0.672757f
C673 VN.n4 VSUBS 0.076428f
C674 VN.n5 VSUBS 0.341788f
C675 VN.n6 VSUBS 0.041008f
C676 VN.n7 VSUBS 0.041008f
C677 VN.n8 VSUBS 0.069006f
C678 VN.n9 VSUBS 0.064354f
C679 VN.n10 VSUBS 0.671656f
C680 VN.n11 VSUBS 0.053352f
C681 VN.n12 VSUBS 0.054065f
C682 VN.t1 VSUBS 1.46836f
C683 VN.n13 VSUBS 0.050722f
C684 VN.t4 VSUBS 1.6932f
C685 VN.n14 VSUBS 0.639934f
C686 VN.t3 VSUBS 1.46836f
C687 VN.n15 VSUBS 0.672757f
C688 VN.n16 VSUBS 0.076428f
C689 VN.n17 VSUBS 0.341788f
C690 VN.n18 VSUBS 0.041008f
C691 VN.n19 VSUBS 0.041008f
C692 VN.n20 VSUBS 0.069006f
C693 VN.n21 VSUBS 0.064354f
C694 VN.n22 VSUBS 0.671656f
C695 VN.n23 VSUBS 1.77379f
C696 VDD1.n0 VSUBS 0.024398f
C697 VDD1.n1 VSUBS 0.022204f
C698 VDD1.n2 VSUBS 0.011931f
C699 VDD1.n3 VSUBS 0.028201f
C700 VDD1.n4 VSUBS 0.012633f
C701 VDD1.n5 VSUBS 0.022204f
C702 VDD1.n6 VSUBS 0.011931f
C703 VDD1.n7 VSUBS 0.028201f
C704 VDD1.n8 VSUBS 0.012633f
C705 VDD1.n9 VSUBS 0.579354f
C706 VDD1.n10 VSUBS 0.011931f
C707 VDD1.t2 VSUBS 0.060301f
C708 VDD1.n11 VSUBS 0.102466f
C709 VDD1.n12 VSUBS 0.017937f
C710 VDD1.n13 VSUBS 0.021151f
C711 VDD1.n14 VSUBS 0.028201f
C712 VDD1.n15 VSUBS 0.012633f
C713 VDD1.n16 VSUBS 0.011931f
C714 VDD1.n17 VSUBS 0.022204f
C715 VDD1.n18 VSUBS 0.022204f
C716 VDD1.n19 VSUBS 0.011931f
C717 VDD1.n20 VSUBS 0.012633f
C718 VDD1.n21 VSUBS 0.028201f
C719 VDD1.n22 VSUBS 0.028201f
C720 VDD1.n23 VSUBS 0.012633f
C721 VDD1.n24 VSUBS 0.011931f
C722 VDD1.n25 VSUBS 0.022204f
C723 VDD1.n26 VSUBS 0.022204f
C724 VDD1.n27 VSUBS 0.011931f
C725 VDD1.n28 VSUBS 0.012633f
C726 VDD1.n29 VSUBS 0.028201f
C727 VDD1.n30 VSUBS 0.068276f
C728 VDD1.n31 VSUBS 0.012633f
C729 VDD1.n32 VSUBS 0.011931f
C730 VDD1.n33 VSUBS 0.050412f
C731 VDD1.n34 VSUBS 0.054519f
C732 VDD1.n35 VSUBS 0.024398f
C733 VDD1.n36 VSUBS 0.022204f
C734 VDD1.n37 VSUBS 0.011931f
C735 VDD1.n38 VSUBS 0.028201f
C736 VDD1.n39 VSUBS 0.012633f
C737 VDD1.n40 VSUBS 0.022204f
C738 VDD1.n41 VSUBS 0.011931f
C739 VDD1.n42 VSUBS 0.028201f
C740 VDD1.n43 VSUBS 0.012633f
C741 VDD1.n44 VSUBS 0.579354f
C742 VDD1.n45 VSUBS 0.011931f
C743 VDD1.t3 VSUBS 0.060301f
C744 VDD1.n46 VSUBS 0.102466f
C745 VDD1.n47 VSUBS 0.017937f
C746 VDD1.n48 VSUBS 0.021151f
C747 VDD1.n49 VSUBS 0.028201f
C748 VDD1.n50 VSUBS 0.012633f
C749 VDD1.n51 VSUBS 0.011931f
C750 VDD1.n52 VSUBS 0.022204f
C751 VDD1.n53 VSUBS 0.022204f
C752 VDD1.n54 VSUBS 0.011931f
C753 VDD1.n55 VSUBS 0.012633f
C754 VDD1.n56 VSUBS 0.028201f
C755 VDD1.n57 VSUBS 0.028201f
C756 VDD1.n58 VSUBS 0.012633f
C757 VDD1.n59 VSUBS 0.011931f
C758 VDD1.n60 VSUBS 0.022204f
C759 VDD1.n61 VSUBS 0.022204f
C760 VDD1.n62 VSUBS 0.011931f
C761 VDD1.n63 VSUBS 0.012633f
C762 VDD1.n64 VSUBS 0.028201f
C763 VDD1.n65 VSUBS 0.068276f
C764 VDD1.n66 VSUBS 0.012633f
C765 VDD1.n67 VSUBS 0.011931f
C766 VDD1.n68 VSUBS 0.050412f
C767 VDD1.n69 VSUBS 0.05395f
C768 VDD1.t1 VSUBS 0.117382f
C769 VDD1.t0 VSUBS 0.117382f
C770 VDD1.n70 VSUBS 0.802682f
C771 VDD1.n71 VSUBS 2.15001f
C772 VDD1.t4 VSUBS 0.117382f
C773 VDD1.t5 VSUBS 0.117382f
C774 VDD1.n72 VSUBS 0.799833f
C775 VDD1.n73 VSUBS 2.15418f
C776 VTAIL.t2 VSUBS 0.168333f
C777 VTAIL.t0 VSUBS 0.168333f
C778 VTAIL.n0 VSUBS 1.02283f
C779 VTAIL.n1 VSUBS 0.826035f
C780 VTAIL.n2 VSUBS 0.034989f
C781 VTAIL.n3 VSUBS 0.031841f
C782 VTAIL.n4 VSUBS 0.01711f
C783 VTAIL.n5 VSUBS 0.040442f
C784 VTAIL.n6 VSUBS 0.018117f
C785 VTAIL.n7 VSUBS 0.031841f
C786 VTAIL.n8 VSUBS 0.01711f
C787 VTAIL.n9 VSUBS 0.040442f
C788 VTAIL.n10 VSUBS 0.018117f
C789 VTAIL.n11 VSUBS 0.830829f
C790 VTAIL.n12 VSUBS 0.01711f
C791 VTAIL.t11 VSUBS 0.086475f
C792 VTAIL.n13 VSUBS 0.146942f
C793 VTAIL.n14 VSUBS 0.025723f
C794 VTAIL.n15 VSUBS 0.030332f
C795 VTAIL.n16 VSUBS 0.040442f
C796 VTAIL.n17 VSUBS 0.018117f
C797 VTAIL.n18 VSUBS 0.01711f
C798 VTAIL.n19 VSUBS 0.031841f
C799 VTAIL.n20 VSUBS 0.031841f
C800 VTAIL.n21 VSUBS 0.01711f
C801 VTAIL.n22 VSUBS 0.018117f
C802 VTAIL.n23 VSUBS 0.040442f
C803 VTAIL.n24 VSUBS 0.040442f
C804 VTAIL.n25 VSUBS 0.018117f
C805 VTAIL.n26 VSUBS 0.01711f
C806 VTAIL.n27 VSUBS 0.031841f
C807 VTAIL.n28 VSUBS 0.031841f
C808 VTAIL.n29 VSUBS 0.01711f
C809 VTAIL.n30 VSUBS 0.018117f
C810 VTAIL.n31 VSUBS 0.040442f
C811 VTAIL.n32 VSUBS 0.097912f
C812 VTAIL.n33 VSUBS 0.018117f
C813 VTAIL.n34 VSUBS 0.01711f
C814 VTAIL.n35 VSUBS 0.072295f
C815 VTAIL.n36 VSUBS 0.049199f
C816 VTAIL.n37 VSUBS 0.385115f
C817 VTAIL.t9 VSUBS 0.168333f
C818 VTAIL.t6 VSUBS 0.168333f
C819 VTAIL.n38 VSUBS 1.02283f
C820 VTAIL.n39 VSUBS 2.26178f
C821 VTAIL.t1 VSUBS 0.168333f
C822 VTAIL.t3 VSUBS 0.168333f
C823 VTAIL.n40 VSUBS 1.02283f
C824 VTAIL.n41 VSUBS 2.26178f
C825 VTAIL.n42 VSUBS 0.034989f
C826 VTAIL.n43 VSUBS 0.031841f
C827 VTAIL.n44 VSUBS 0.01711f
C828 VTAIL.n45 VSUBS 0.040442f
C829 VTAIL.n46 VSUBS 0.018117f
C830 VTAIL.n47 VSUBS 0.031841f
C831 VTAIL.n48 VSUBS 0.01711f
C832 VTAIL.n49 VSUBS 0.040442f
C833 VTAIL.n50 VSUBS 0.018117f
C834 VTAIL.n51 VSUBS 0.830829f
C835 VTAIL.n52 VSUBS 0.01711f
C836 VTAIL.t5 VSUBS 0.086475f
C837 VTAIL.n53 VSUBS 0.146942f
C838 VTAIL.n54 VSUBS 0.025723f
C839 VTAIL.n55 VSUBS 0.030332f
C840 VTAIL.n56 VSUBS 0.040442f
C841 VTAIL.n57 VSUBS 0.018117f
C842 VTAIL.n58 VSUBS 0.01711f
C843 VTAIL.n59 VSUBS 0.031841f
C844 VTAIL.n60 VSUBS 0.031841f
C845 VTAIL.n61 VSUBS 0.01711f
C846 VTAIL.n62 VSUBS 0.018117f
C847 VTAIL.n63 VSUBS 0.040442f
C848 VTAIL.n64 VSUBS 0.040442f
C849 VTAIL.n65 VSUBS 0.018117f
C850 VTAIL.n66 VSUBS 0.01711f
C851 VTAIL.n67 VSUBS 0.031841f
C852 VTAIL.n68 VSUBS 0.031841f
C853 VTAIL.n69 VSUBS 0.01711f
C854 VTAIL.n70 VSUBS 0.018117f
C855 VTAIL.n71 VSUBS 0.040442f
C856 VTAIL.n72 VSUBS 0.097912f
C857 VTAIL.n73 VSUBS 0.018117f
C858 VTAIL.n74 VSUBS 0.01711f
C859 VTAIL.n75 VSUBS 0.072295f
C860 VTAIL.n76 VSUBS 0.049199f
C861 VTAIL.n77 VSUBS 0.385115f
C862 VTAIL.t7 VSUBS 0.168333f
C863 VTAIL.t10 VSUBS 0.168333f
C864 VTAIL.n78 VSUBS 1.02283f
C865 VTAIL.n79 VSUBS 0.975284f
C866 VTAIL.n80 VSUBS 0.034989f
C867 VTAIL.n81 VSUBS 0.031841f
C868 VTAIL.n82 VSUBS 0.01711f
C869 VTAIL.n83 VSUBS 0.040442f
C870 VTAIL.n84 VSUBS 0.018117f
C871 VTAIL.n85 VSUBS 0.031841f
C872 VTAIL.n86 VSUBS 0.01711f
C873 VTAIL.n87 VSUBS 0.040442f
C874 VTAIL.n88 VSUBS 0.018117f
C875 VTAIL.n89 VSUBS 0.830829f
C876 VTAIL.n90 VSUBS 0.01711f
C877 VTAIL.t8 VSUBS 0.086475f
C878 VTAIL.n91 VSUBS 0.146942f
C879 VTAIL.n92 VSUBS 0.025723f
C880 VTAIL.n93 VSUBS 0.030332f
C881 VTAIL.n94 VSUBS 0.040442f
C882 VTAIL.n95 VSUBS 0.018117f
C883 VTAIL.n96 VSUBS 0.01711f
C884 VTAIL.n97 VSUBS 0.031841f
C885 VTAIL.n98 VSUBS 0.031841f
C886 VTAIL.n99 VSUBS 0.01711f
C887 VTAIL.n100 VSUBS 0.018117f
C888 VTAIL.n101 VSUBS 0.040442f
C889 VTAIL.n102 VSUBS 0.040442f
C890 VTAIL.n103 VSUBS 0.018117f
C891 VTAIL.n104 VSUBS 0.01711f
C892 VTAIL.n105 VSUBS 0.031841f
C893 VTAIL.n106 VSUBS 0.031841f
C894 VTAIL.n107 VSUBS 0.01711f
C895 VTAIL.n108 VSUBS 0.018117f
C896 VTAIL.n109 VSUBS 0.040442f
C897 VTAIL.n110 VSUBS 0.097912f
C898 VTAIL.n111 VSUBS 0.018117f
C899 VTAIL.n112 VSUBS 0.01711f
C900 VTAIL.n113 VSUBS 0.072295f
C901 VTAIL.n114 VSUBS 0.049199f
C902 VTAIL.n115 VSUBS 1.46464f
C903 VTAIL.n116 VSUBS 0.034989f
C904 VTAIL.n117 VSUBS 0.031841f
C905 VTAIL.n118 VSUBS 0.01711f
C906 VTAIL.n119 VSUBS 0.040442f
C907 VTAIL.n120 VSUBS 0.018117f
C908 VTAIL.n121 VSUBS 0.031841f
C909 VTAIL.n122 VSUBS 0.01711f
C910 VTAIL.n123 VSUBS 0.040442f
C911 VTAIL.n124 VSUBS 0.018117f
C912 VTAIL.n125 VSUBS 0.830829f
C913 VTAIL.n126 VSUBS 0.01711f
C914 VTAIL.t4 VSUBS 0.086475f
C915 VTAIL.n127 VSUBS 0.146942f
C916 VTAIL.n128 VSUBS 0.025723f
C917 VTAIL.n129 VSUBS 0.030332f
C918 VTAIL.n130 VSUBS 0.040442f
C919 VTAIL.n131 VSUBS 0.018117f
C920 VTAIL.n132 VSUBS 0.01711f
C921 VTAIL.n133 VSUBS 0.031841f
C922 VTAIL.n134 VSUBS 0.031841f
C923 VTAIL.n135 VSUBS 0.01711f
C924 VTAIL.n136 VSUBS 0.018117f
C925 VTAIL.n137 VSUBS 0.040442f
C926 VTAIL.n138 VSUBS 0.040442f
C927 VTAIL.n139 VSUBS 0.018117f
C928 VTAIL.n140 VSUBS 0.01711f
C929 VTAIL.n141 VSUBS 0.031841f
C930 VTAIL.n142 VSUBS 0.031841f
C931 VTAIL.n143 VSUBS 0.01711f
C932 VTAIL.n144 VSUBS 0.018117f
C933 VTAIL.n145 VSUBS 0.040442f
C934 VTAIL.n146 VSUBS 0.097912f
C935 VTAIL.n147 VSUBS 0.018117f
C936 VTAIL.n148 VSUBS 0.01711f
C937 VTAIL.n149 VSUBS 0.072295f
C938 VTAIL.n150 VSUBS 0.049199f
C939 VTAIL.n151 VSUBS 1.40693f
C940 VP.n0 VSUBS 0.05631f
C941 VP.t5 VSUBS 1.52935f
C942 VP.n1 VSUBS 0.052829f
C943 VP.n2 VSUBS 0.042711f
C944 VP.t4 VSUBS 1.52935f
C945 VP.n3 VSUBS 0.052829f
C946 VP.n4 VSUBS 0.05631f
C947 VP.t2 VSUBS 1.52935f
C948 VP.n5 VSUBS 0.05631f
C949 VP.t0 VSUBS 1.52935f
C950 VP.n6 VSUBS 0.052829f
C951 VP.t3 VSUBS 1.76352f
C952 VP.n7 VSUBS 0.666512f
C953 VP.t1 VSUBS 1.52935f
C954 VP.n8 VSUBS 0.700698f
C955 VP.n9 VSUBS 0.079603f
C956 VP.n10 VSUBS 0.355983f
C957 VP.n11 VSUBS 0.042711f
C958 VP.n12 VSUBS 0.042711f
C959 VP.n13 VSUBS 0.071872f
C960 VP.n14 VSUBS 0.067026f
C961 VP.n15 VSUBS 0.699551f
C962 VP.n16 VSUBS 1.82384f
C963 VP.n17 VSUBS 1.86012f
C964 VP.n18 VSUBS 0.699551f
C965 VP.n19 VSUBS 0.067026f
C966 VP.n20 VSUBS 0.071872f
C967 VP.n21 VSUBS 0.042711f
C968 VP.n22 VSUBS 0.042711f
C969 VP.n23 VSUBS 0.042711f
C970 VP.n24 VSUBS 0.079603f
C971 VP.n25 VSUBS 0.616117f
C972 VP.n26 VSUBS 0.079603f
C973 VP.n27 VSUBS 0.042711f
C974 VP.n28 VSUBS 0.042711f
C975 VP.n29 VSUBS 0.042711f
C976 VP.n30 VSUBS 0.071872f
C977 VP.n31 VSUBS 0.067026f
C978 VP.n32 VSUBS 0.699551f
C979 VP.n33 VSUBS 0.055568f
.ends

