* NGSPICE file created from diff_pair_sample_1160.ext - technology: sky130A

.subckt diff_pair_sample_1160 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=3.69
X1 VDD1.t9 VP.t0 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=3.69
X2 VDD2.t9 VN.t0 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=3.69
X3 VTAIL.t8 VN.t1 VDD2.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X4 VDD1.t8 VP.t1 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=3.69
X5 VTAIL.t18 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X6 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=3.69
X7 VDD2.t7 VN.t2 VTAIL.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X8 VDD1.t6 VP.t3 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X9 VTAIL.t11 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X10 VTAIL.t12 VP.t5 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X11 VTAIL.t0 VN.t3 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X12 VDD1.t3 VP.t6 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=3.69
X13 VDD2.t5 VN.t4 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=3.69
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=3.69
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=3.69
X16 VDD2.t4 VN.t5 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X17 VTAIL.t2 VN.t6 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X18 VDD2.t2 VN.t7 VTAIL.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=3.69
X19 VDD2.t1 VN.t8 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=3.69
X20 VDD1.t2 VP.t7 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=3.69
X21 VTAIL.t1 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X22 VTAIL.t19 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
X23 VDD1.t0 VP.t9 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=3.69
R0 B.n888 B.n887 585
R1 B.n889 B.n888 585
R2 B.n266 B.n168 585
R3 B.n265 B.n264 585
R4 B.n263 B.n262 585
R5 B.n261 B.n260 585
R6 B.n259 B.n258 585
R7 B.n257 B.n256 585
R8 B.n255 B.n254 585
R9 B.n253 B.n252 585
R10 B.n251 B.n250 585
R11 B.n249 B.n248 585
R12 B.n247 B.n246 585
R13 B.n245 B.n244 585
R14 B.n243 B.n242 585
R15 B.n241 B.n240 585
R16 B.n239 B.n238 585
R17 B.n237 B.n236 585
R18 B.n235 B.n234 585
R19 B.n233 B.n232 585
R20 B.n231 B.n230 585
R21 B.n228 B.n227 585
R22 B.n226 B.n225 585
R23 B.n224 B.n223 585
R24 B.n222 B.n221 585
R25 B.n220 B.n219 585
R26 B.n218 B.n217 585
R27 B.n216 B.n215 585
R28 B.n214 B.n213 585
R29 B.n212 B.n211 585
R30 B.n210 B.n209 585
R31 B.n208 B.n207 585
R32 B.n206 B.n205 585
R33 B.n204 B.n203 585
R34 B.n202 B.n201 585
R35 B.n200 B.n199 585
R36 B.n198 B.n197 585
R37 B.n196 B.n195 585
R38 B.n194 B.n193 585
R39 B.n192 B.n191 585
R40 B.n190 B.n189 585
R41 B.n188 B.n187 585
R42 B.n186 B.n185 585
R43 B.n184 B.n183 585
R44 B.n182 B.n181 585
R45 B.n180 B.n179 585
R46 B.n178 B.n177 585
R47 B.n176 B.n175 585
R48 B.n144 B.n143 585
R49 B.n892 B.n891 585
R50 B.n886 B.n169 585
R51 B.n169 B.n141 585
R52 B.n885 B.n140 585
R53 B.n896 B.n140 585
R54 B.n884 B.n139 585
R55 B.n897 B.n139 585
R56 B.n883 B.n138 585
R57 B.n898 B.n138 585
R58 B.n882 B.n881 585
R59 B.n881 B.n134 585
R60 B.n880 B.n133 585
R61 B.n904 B.n133 585
R62 B.n879 B.n132 585
R63 B.n905 B.n132 585
R64 B.n878 B.n131 585
R65 B.n906 B.n131 585
R66 B.n877 B.n876 585
R67 B.n876 B.n127 585
R68 B.n875 B.n126 585
R69 B.n912 B.n126 585
R70 B.n874 B.n125 585
R71 B.n913 B.n125 585
R72 B.n873 B.n124 585
R73 B.n914 B.n124 585
R74 B.n872 B.n871 585
R75 B.n871 B.n120 585
R76 B.n870 B.n119 585
R77 B.n920 B.n119 585
R78 B.n869 B.n118 585
R79 B.n921 B.n118 585
R80 B.n868 B.n117 585
R81 B.n922 B.n117 585
R82 B.n867 B.n866 585
R83 B.n866 B.n113 585
R84 B.n865 B.n112 585
R85 B.n928 B.n112 585
R86 B.n864 B.n111 585
R87 B.n929 B.n111 585
R88 B.n863 B.n110 585
R89 B.n930 B.n110 585
R90 B.n862 B.n861 585
R91 B.n861 B.n106 585
R92 B.n860 B.n105 585
R93 B.n936 B.n105 585
R94 B.n859 B.n104 585
R95 B.n937 B.n104 585
R96 B.n858 B.n103 585
R97 B.n938 B.n103 585
R98 B.n857 B.n856 585
R99 B.n856 B.n102 585
R100 B.n855 B.n98 585
R101 B.n944 B.n98 585
R102 B.n854 B.n97 585
R103 B.n945 B.n97 585
R104 B.n853 B.n96 585
R105 B.n946 B.n96 585
R106 B.n852 B.n851 585
R107 B.n851 B.n92 585
R108 B.n850 B.n91 585
R109 B.n952 B.n91 585
R110 B.n849 B.n90 585
R111 B.n953 B.n90 585
R112 B.n848 B.n89 585
R113 B.n954 B.n89 585
R114 B.n847 B.n846 585
R115 B.n846 B.n85 585
R116 B.n845 B.n84 585
R117 B.n960 B.n84 585
R118 B.n844 B.n83 585
R119 B.n961 B.n83 585
R120 B.n843 B.n82 585
R121 B.n962 B.n82 585
R122 B.n842 B.n841 585
R123 B.n841 B.n81 585
R124 B.n840 B.n77 585
R125 B.n968 B.n77 585
R126 B.n839 B.n76 585
R127 B.n969 B.n76 585
R128 B.n838 B.n75 585
R129 B.n970 B.n75 585
R130 B.n837 B.n836 585
R131 B.n836 B.n71 585
R132 B.n835 B.n70 585
R133 B.n976 B.n70 585
R134 B.n834 B.n69 585
R135 B.n977 B.n69 585
R136 B.n833 B.n68 585
R137 B.n978 B.n68 585
R138 B.n832 B.n831 585
R139 B.n831 B.n64 585
R140 B.n830 B.n63 585
R141 B.n984 B.n63 585
R142 B.n829 B.n62 585
R143 B.n985 B.n62 585
R144 B.n828 B.n61 585
R145 B.n986 B.n61 585
R146 B.n827 B.n826 585
R147 B.n826 B.n57 585
R148 B.n825 B.n56 585
R149 B.n992 B.n56 585
R150 B.n824 B.n55 585
R151 B.n993 B.n55 585
R152 B.n823 B.n54 585
R153 B.n994 B.n54 585
R154 B.n822 B.n821 585
R155 B.n821 B.n50 585
R156 B.n820 B.n49 585
R157 B.n1000 B.n49 585
R158 B.n819 B.n48 585
R159 B.n1001 B.n48 585
R160 B.n818 B.n47 585
R161 B.n1002 B.n47 585
R162 B.n817 B.n816 585
R163 B.n816 B.n43 585
R164 B.n815 B.n42 585
R165 B.n1008 B.n42 585
R166 B.n814 B.n41 585
R167 B.n1009 B.n41 585
R168 B.n813 B.n40 585
R169 B.n1010 B.n40 585
R170 B.n812 B.n811 585
R171 B.n811 B.n36 585
R172 B.n810 B.n35 585
R173 B.n1016 B.n35 585
R174 B.n809 B.n34 585
R175 B.n1017 B.n34 585
R176 B.n808 B.n33 585
R177 B.n1018 B.n33 585
R178 B.n807 B.n806 585
R179 B.n806 B.n29 585
R180 B.n805 B.n28 585
R181 B.n1024 B.n28 585
R182 B.n804 B.n27 585
R183 B.n1025 B.n27 585
R184 B.n803 B.n26 585
R185 B.n1026 B.n26 585
R186 B.n802 B.n801 585
R187 B.n801 B.n22 585
R188 B.n800 B.n21 585
R189 B.n1032 B.n21 585
R190 B.n799 B.n20 585
R191 B.n1033 B.n20 585
R192 B.n798 B.n19 585
R193 B.n1034 B.n19 585
R194 B.n797 B.n796 585
R195 B.n796 B.n15 585
R196 B.n795 B.n14 585
R197 B.n1040 B.n14 585
R198 B.n794 B.n13 585
R199 B.n1041 B.n13 585
R200 B.n793 B.n12 585
R201 B.n1042 B.n12 585
R202 B.n792 B.n791 585
R203 B.n791 B.n8 585
R204 B.n790 B.n7 585
R205 B.n1048 B.n7 585
R206 B.n789 B.n6 585
R207 B.n1049 B.n6 585
R208 B.n788 B.n5 585
R209 B.n1050 B.n5 585
R210 B.n787 B.n786 585
R211 B.n786 B.n4 585
R212 B.n785 B.n267 585
R213 B.n785 B.n784 585
R214 B.n775 B.n268 585
R215 B.n269 B.n268 585
R216 B.n777 B.n776 585
R217 B.n778 B.n777 585
R218 B.n774 B.n274 585
R219 B.n274 B.n273 585
R220 B.n773 B.n772 585
R221 B.n772 B.n771 585
R222 B.n276 B.n275 585
R223 B.n277 B.n276 585
R224 B.n764 B.n763 585
R225 B.n765 B.n764 585
R226 B.n762 B.n282 585
R227 B.n282 B.n281 585
R228 B.n761 B.n760 585
R229 B.n760 B.n759 585
R230 B.n284 B.n283 585
R231 B.n285 B.n284 585
R232 B.n752 B.n751 585
R233 B.n753 B.n752 585
R234 B.n750 B.n290 585
R235 B.n290 B.n289 585
R236 B.n749 B.n748 585
R237 B.n748 B.n747 585
R238 B.n292 B.n291 585
R239 B.n293 B.n292 585
R240 B.n740 B.n739 585
R241 B.n741 B.n740 585
R242 B.n738 B.n298 585
R243 B.n298 B.n297 585
R244 B.n737 B.n736 585
R245 B.n736 B.n735 585
R246 B.n300 B.n299 585
R247 B.n301 B.n300 585
R248 B.n728 B.n727 585
R249 B.n729 B.n728 585
R250 B.n726 B.n306 585
R251 B.n306 B.n305 585
R252 B.n725 B.n724 585
R253 B.n724 B.n723 585
R254 B.n308 B.n307 585
R255 B.n309 B.n308 585
R256 B.n716 B.n715 585
R257 B.n717 B.n716 585
R258 B.n714 B.n314 585
R259 B.n314 B.n313 585
R260 B.n713 B.n712 585
R261 B.n712 B.n711 585
R262 B.n316 B.n315 585
R263 B.n317 B.n316 585
R264 B.n704 B.n703 585
R265 B.n705 B.n704 585
R266 B.n702 B.n322 585
R267 B.n322 B.n321 585
R268 B.n701 B.n700 585
R269 B.n700 B.n699 585
R270 B.n324 B.n323 585
R271 B.n325 B.n324 585
R272 B.n692 B.n691 585
R273 B.n693 B.n692 585
R274 B.n690 B.n330 585
R275 B.n330 B.n329 585
R276 B.n689 B.n688 585
R277 B.n688 B.n687 585
R278 B.n332 B.n331 585
R279 B.n333 B.n332 585
R280 B.n680 B.n679 585
R281 B.n681 B.n680 585
R282 B.n678 B.n338 585
R283 B.n338 B.n337 585
R284 B.n677 B.n676 585
R285 B.n676 B.n675 585
R286 B.n340 B.n339 585
R287 B.n341 B.n340 585
R288 B.n668 B.n667 585
R289 B.n669 B.n668 585
R290 B.n666 B.n346 585
R291 B.n346 B.n345 585
R292 B.n665 B.n664 585
R293 B.n664 B.n663 585
R294 B.n348 B.n347 585
R295 B.n656 B.n348 585
R296 B.n655 B.n654 585
R297 B.n657 B.n655 585
R298 B.n653 B.n353 585
R299 B.n353 B.n352 585
R300 B.n652 B.n651 585
R301 B.n651 B.n650 585
R302 B.n355 B.n354 585
R303 B.n356 B.n355 585
R304 B.n643 B.n642 585
R305 B.n644 B.n643 585
R306 B.n641 B.n361 585
R307 B.n361 B.n360 585
R308 B.n640 B.n639 585
R309 B.n639 B.n638 585
R310 B.n363 B.n362 585
R311 B.n364 B.n363 585
R312 B.n631 B.n630 585
R313 B.n632 B.n631 585
R314 B.n629 B.n369 585
R315 B.n369 B.n368 585
R316 B.n628 B.n627 585
R317 B.n627 B.n626 585
R318 B.n371 B.n370 585
R319 B.n619 B.n371 585
R320 B.n618 B.n617 585
R321 B.n620 B.n618 585
R322 B.n616 B.n376 585
R323 B.n376 B.n375 585
R324 B.n615 B.n614 585
R325 B.n614 B.n613 585
R326 B.n378 B.n377 585
R327 B.n379 B.n378 585
R328 B.n606 B.n605 585
R329 B.n607 B.n606 585
R330 B.n604 B.n384 585
R331 B.n384 B.n383 585
R332 B.n603 B.n602 585
R333 B.n602 B.n601 585
R334 B.n386 B.n385 585
R335 B.n387 B.n386 585
R336 B.n594 B.n593 585
R337 B.n595 B.n594 585
R338 B.n592 B.n392 585
R339 B.n392 B.n391 585
R340 B.n591 B.n590 585
R341 B.n590 B.n589 585
R342 B.n394 B.n393 585
R343 B.n395 B.n394 585
R344 B.n582 B.n581 585
R345 B.n583 B.n582 585
R346 B.n580 B.n400 585
R347 B.n400 B.n399 585
R348 B.n579 B.n578 585
R349 B.n578 B.n577 585
R350 B.n402 B.n401 585
R351 B.n403 B.n402 585
R352 B.n570 B.n569 585
R353 B.n571 B.n570 585
R354 B.n568 B.n408 585
R355 B.n408 B.n407 585
R356 B.n567 B.n566 585
R357 B.n566 B.n565 585
R358 B.n410 B.n409 585
R359 B.n411 B.n410 585
R360 B.n558 B.n557 585
R361 B.n559 B.n558 585
R362 B.n556 B.n416 585
R363 B.n416 B.n415 585
R364 B.n555 B.n554 585
R365 B.n554 B.n553 585
R366 B.n418 B.n417 585
R367 B.n419 B.n418 585
R368 B.n549 B.n548 585
R369 B.n422 B.n421 585
R370 B.n545 B.n544 585
R371 B.n546 B.n545 585
R372 B.n543 B.n446 585
R373 B.n542 B.n541 585
R374 B.n540 B.n539 585
R375 B.n538 B.n537 585
R376 B.n536 B.n535 585
R377 B.n534 B.n533 585
R378 B.n532 B.n531 585
R379 B.n530 B.n529 585
R380 B.n528 B.n527 585
R381 B.n526 B.n525 585
R382 B.n524 B.n523 585
R383 B.n522 B.n521 585
R384 B.n520 B.n519 585
R385 B.n518 B.n517 585
R386 B.n516 B.n515 585
R387 B.n514 B.n513 585
R388 B.n512 B.n511 585
R389 B.n509 B.n508 585
R390 B.n507 B.n506 585
R391 B.n505 B.n504 585
R392 B.n503 B.n502 585
R393 B.n501 B.n500 585
R394 B.n499 B.n498 585
R395 B.n497 B.n496 585
R396 B.n495 B.n494 585
R397 B.n493 B.n492 585
R398 B.n491 B.n490 585
R399 B.n489 B.n488 585
R400 B.n487 B.n486 585
R401 B.n485 B.n484 585
R402 B.n483 B.n482 585
R403 B.n481 B.n480 585
R404 B.n479 B.n478 585
R405 B.n477 B.n476 585
R406 B.n475 B.n474 585
R407 B.n473 B.n472 585
R408 B.n471 B.n470 585
R409 B.n469 B.n468 585
R410 B.n467 B.n466 585
R411 B.n465 B.n464 585
R412 B.n463 B.n462 585
R413 B.n461 B.n460 585
R414 B.n459 B.n458 585
R415 B.n457 B.n456 585
R416 B.n455 B.n454 585
R417 B.n453 B.n452 585
R418 B.n550 B.n420 585
R419 B.n420 B.n419 585
R420 B.n552 B.n551 585
R421 B.n553 B.n552 585
R422 B.n414 B.n413 585
R423 B.n415 B.n414 585
R424 B.n561 B.n560 585
R425 B.n560 B.n559 585
R426 B.n562 B.n412 585
R427 B.n412 B.n411 585
R428 B.n564 B.n563 585
R429 B.n565 B.n564 585
R430 B.n406 B.n405 585
R431 B.n407 B.n406 585
R432 B.n573 B.n572 585
R433 B.n572 B.n571 585
R434 B.n574 B.n404 585
R435 B.n404 B.n403 585
R436 B.n576 B.n575 585
R437 B.n577 B.n576 585
R438 B.n398 B.n397 585
R439 B.n399 B.n398 585
R440 B.n585 B.n584 585
R441 B.n584 B.n583 585
R442 B.n586 B.n396 585
R443 B.n396 B.n395 585
R444 B.n588 B.n587 585
R445 B.n589 B.n588 585
R446 B.n390 B.n389 585
R447 B.n391 B.n390 585
R448 B.n597 B.n596 585
R449 B.n596 B.n595 585
R450 B.n598 B.n388 585
R451 B.n388 B.n387 585
R452 B.n600 B.n599 585
R453 B.n601 B.n600 585
R454 B.n382 B.n381 585
R455 B.n383 B.n382 585
R456 B.n609 B.n608 585
R457 B.n608 B.n607 585
R458 B.n610 B.n380 585
R459 B.n380 B.n379 585
R460 B.n612 B.n611 585
R461 B.n613 B.n612 585
R462 B.n374 B.n373 585
R463 B.n375 B.n374 585
R464 B.n622 B.n621 585
R465 B.n621 B.n620 585
R466 B.n623 B.n372 585
R467 B.n619 B.n372 585
R468 B.n625 B.n624 585
R469 B.n626 B.n625 585
R470 B.n367 B.n366 585
R471 B.n368 B.n367 585
R472 B.n634 B.n633 585
R473 B.n633 B.n632 585
R474 B.n635 B.n365 585
R475 B.n365 B.n364 585
R476 B.n637 B.n636 585
R477 B.n638 B.n637 585
R478 B.n359 B.n358 585
R479 B.n360 B.n359 585
R480 B.n646 B.n645 585
R481 B.n645 B.n644 585
R482 B.n647 B.n357 585
R483 B.n357 B.n356 585
R484 B.n649 B.n648 585
R485 B.n650 B.n649 585
R486 B.n351 B.n350 585
R487 B.n352 B.n351 585
R488 B.n659 B.n658 585
R489 B.n658 B.n657 585
R490 B.n660 B.n349 585
R491 B.n656 B.n349 585
R492 B.n662 B.n661 585
R493 B.n663 B.n662 585
R494 B.n344 B.n343 585
R495 B.n345 B.n344 585
R496 B.n671 B.n670 585
R497 B.n670 B.n669 585
R498 B.n672 B.n342 585
R499 B.n342 B.n341 585
R500 B.n674 B.n673 585
R501 B.n675 B.n674 585
R502 B.n336 B.n335 585
R503 B.n337 B.n336 585
R504 B.n683 B.n682 585
R505 B.n682 B.n681 585
R506 B.n684 B.n334 585
R507 B.n334 B.n333 585
R508 B.n686 B.n685 585
R509 B.n687 B.n686 585
R510 B.n328 B.n327 585
R511 B.n329 B.n328 585
R512 B.n695 B.n694 585
R513 B.n694 B.n693 585
R514 B.n696 B.n326 585
R515 B.n326 B.n325 585
R516 B.n698 B.n697 585
R517 B.n699 B.n698 585
R518 B.n320 B.n319 585
R519 B.n321 B.n320 585
R520 B.n707 B.n706 585
R521 B.n706 B.n705 585
R522 B.n708 B.n318 585
R523 B.n318 B.n317 585
R524 B.n710 B.n709 585
R525 B.n711 B.n710 585
R526 B.n312 B.n311 585
R527 B.n313 B.n312 585
R528 B.n719 B.n718 585
R529 B.n718 B.n717 585
R530 B.n720 B.n310 585
R531 B.n310 B.n309 585
R532 B.n722 B.n721 585
R533 B.n723 B.n722 585
R534 B.n304 B.n303 585
R535 B.n305 B.n304 585
R536 B.n731 B.n730 585
R537 B.n730 B.n729 585
R538 B.n732 B.n302 585
R539 B.n302 B.n301 585
R540 B.n734 B.n733 585
R541 B.n735 B.n734 585
R542 B.n296 B.n295 585
R543 B.n297 B.n296 585
R544 B.n743 B.n742 585
R545 B.n742 B.n741 585
R546 B.n744 B.n294 585
R547 B.n294 B.n293 585
R548 B.n746 B.n745 585
R549 B.n747 B.n746 585
R550 B.n288 B.n287 585
R551 B.n289 B.n288 585
R552 B.n755 B.n754 585
R553 B.n754 B.n753 585
R554 B.n756 B.n286 585
R555 B.n286 B.n285 585
R556 B.n758 B.n757 585
R557 B.n759 B.n758 585
R558 B.n280 B.n279 585
R559 B.n281 B.n280 585
R560 B.n767 B.n766 585
R561 B.n766 B.n765 585
R562 B.n768 B.n278 585
R563 B.n278 B.n277 585
R564 B.n770 B.n769 585
R565 B.n771 B.n770 585
R566 B.n272 B.n271 585
R567 B.n273 B.n272 585
R568 B.n780 B.n779 585
R569 B.n779 B.n778 585
R570 B.n781 B.n270 585
R571 B.n270 B.n269 585
R572 B.n783 B.n782 585
R573 B.n784 B.n783 585
R574 B.n2 B.n0 585
R575 B.n4 B.n2 585
R576 B.n3 B.n1 585
R577 B.n1049 B.n3 585
R578 B.n1047 B.n1046 585
R579 B.n1048 B.n1047 585
R580 B.n1045 B.n9 585
R581 B.n9 B.n8 585
R582 B.n1044 B.n1043 585
R583 B.n1043 B.n1042 585
R584 B.n11 B.n10 585
R585 B.n1041 B.n11 585
R586 B.n1039 B.n1038 585
R587 B.n1040 B.n1039 585
R588 B.n1037 B.n16 585
R589 B.n16 B.n15 585
R590 B.n1036 B.n1035 585
R591 B.n1035 B.n1034 585
R592 B.n18 B.n17 585
R593 B.n1033 B.n18 585
R594 B.n1031 B.n1030 585
R595 B.n1032 B.n1031 585
R596 B.n1029 B.n23 585
R597 B.n23 B.n22 585
R598 B.n1028 B.n1027 585
R599 B.n1027 B.n1026 585
R600 B.n25 B.n24 585
R601 B.n1025 B.n25 585
R602 B.n1023 B.n1022 585
R603 B.n1024 B.n1023 585
R604 B.n1021 B.n30 585
R605 B.n30 B.n29 585
R606 B.n1020 B.n1019 585
R607 B.n1019 B.n1018 585
R608 B.n32 B.n31 585
R609 B.n1017 B.n32 585
R610 B.n1015 B.n1014 585
R611 B.n1016 B.n1015 585
R612 B.n1013 B.n37 585
R613 B.n37 B.n36 585
R614 B.n1012 B.n1011 585
R615 B.n1011 B.n1010 585
R616 B.n39 B.n38 585
R617 B.n1009 B.n39 585
R618 B.n1007 B.n1006 585
R619 B.n1008 B.n1007 585
R620 B.n1005 B.n44 585
R621 B.n44 B.n43 585
R622 B.n1004 B.n1003 585
R623 B.n1003 B.n1002 585
R624 B.n46 B.n45 585
R625 B.n1001 B.n46 585
R626 B.n999 B.n998 585
R627 B.n1000 B.n999 585
R628 B.n997 B.n51 585
R629 B.n51 B.n50 585
R630 B.n996 B.n995 585
R631 B.n995 B.n994 585
R632 B.n53 B.n52 585
R633 B.n993 B.n53 585
R634 B.n991 B.n990 585
R635 B.n992 B.n991 585
R636 B.n989 B.n58 585
R637 B.n58 B.n57 585
R638 B.n988 B.n987 585
R639 B.n987 B.n986 585
R640 B.n60 B.n59 585
R641 B.n985 B.n60 585
R642 B.n983 B.n982 585
R643 B.n984 B.n983 585
R644 B.n981 B.n65 585
R645 B.n65 B.n64 585
R646 B.n980 B.n979 585
R647 B.n979 B.n978 585
R648 B.n67 B.n66 585
R649 B.n977 B.n67 585
R650 B.n975 B.n974 585
R651 B.n976 B.n975 585
R652 B.n973 B.n72 585
R653 B.n72 B.n71 585
R654 B.n972 B.n971 585
R655 B.n971 B.n970 585
R656 B.n74 B.n73 585
R657 B.n969 B.n74 585
R658 B.n967 B.n966 585
R659 B.n968 B.n967 585
R660 B.n965 B.n78 585
R661 B.n81 B.n78 585
R662 B.n964 B.n963 585
R663 B.n963 B.n962 585
R664 B.n80 B.n79 585
R665 B.n961 B.n80 585
R666 B.n959 B.n958 585
R667 B.n960 B.n959 585
R668 B.n957 B.n86 585
R669 B.n86 B.n85 585
R670 B.n956 B.n955 585
R671 B.n955 B.n954 585
R672 B.n88 B.n87 585
R673 B.n953 B.n88 585
R674 B.n951 B.n950 585
R675 B.n952 B.n951 585
R676 B.n949 B.n93 585
R677 B.n93 B.n92 585
R678 B.n948 B.n947 585
R679 B.n947 B.n946 585
R680 B.n95 B.n94 585
R681 B.n945 B.n95 585
R682 B.n943 B.n942 585
R683 B.n944 B.n943 585
R684 B.n941 B.n99 585
R685 B.n102 B.n99 585
R686 B.n940 B.n939 585
R687 B.n939 B.n938 585
R688 B.n101 B.n100 585
R689 B.n937 B.n101 585
R690 B.n935 B.n934 585
R691 B.n936 B.n935 585
R692 B.n933 B.n107 585
R693 B.n107 B.n106 585
R694 B.n932 B.n931 585
R695 B.n931 B.n930 585
R696 B.n109 B.n108 585
R697 B.n929 B.n109 585
R698 B.n927 B.n926 585
R699 B.n928 B.n927 585
R700 B.n925 B.n114 585
R701 B.n114 B.n113 585
R702 B.n924 B.n923 585
R703 B.n923 B.n922 585
R704 B.n116 B.n115 585
R705 B.n921 B.n116 585
R706 B.n919 B.n918 585
R707 B.n920 B.n919 585
R708 B.n917 B.n121 585
R709 B.n121 B.n120 585
R710 B.n916 B.n915 585
R711 B.n915 B.n914 585
R712 B.n123 B.n122 585
R713 B.n913 B.n123 585
R714 B.n911 B.n910 585
R715 B.n912 B.n911 585
R716 B.n909 B.n128 585
R717 B.n128 B.n127 585
R718 B.n908 B.n907 585
R719 B.n907 B.n906 585
R720 B.n130 B.n129 585
R721 B.n905 B.n130 585
R722 B.n903 B.n902 585
R723 B.n904 B.n903 585
R724 B.n901 B.n135 585
R725 B.n135 B.n134 585
R726 B.n900 B.n899 585
R727 B.n899 B.n898 585
R728 B.n137 B.n136 585
R729 B.n897 B.n137 585
R730 B.n895 B.n894 585
R731 B.n896 B.n895 585
R732 B.n893 B.n142 585
R733 B.n142 B.n141 585
R734 B.n1052 B.n1051 585
R735 B.n1051 B.n1050 585
R736 B.n548 B.n420 535.745
R737 B.n891 B.n142 535.745
R738 B.n452 B.n418 535.745
R739 B.n888 B.n169 535.745
R740 B.n889 B.n167 256.663
R741 B.n889 B.n166 256.663
R742 B.n889 B.n165 256.663
R743 B.n889 B.n164 256.663
R744 B.n889 B.n163 256.663
R745 B.n889 B.n162 256.663
R746 B.n889 B.n161 256.663
R747 B.n889 B.n160 256.663
R748 B.n889 B.n159 256.663
R749 B.n889 B.n158 256.663
R750 B.n889 B.n157 256.663
R751 B.n889 B.n156 256.663
R752 B.n889 B.n155 256.663
R753 B.n889 B.n154 256.663
R754 B.n889 B.n153 256.663
R755 B.n889 B.n152 256.663
R756 B.n889 B.n151 256.663
R757 B.n889 B.n150 256.663
R758 B.n889 B.n149 256.663
R759 B.n889 B.n148 256.663
R760 B.n889 B.n147 256.663
R761 B.n889 B.n146 256.663
R762 B.n889 B.n145 256.663
R763 B.n890 B.n889 256.663
R764 B.n547 B.n546 256.663
R765 B.n546 B.n423 256.663
R766 B.n546 B.n424 256.663
R767 B.n546 B.n425 256.663
R768 B.n546 B.n426 256.663
R769 B.n546 B.n427 256.663
R770 B.n546 B.n428 256.663
R771 B.n546 B.n429 256.663
R772 B.n546 B.n430 256.663
R773 B.n546 B.n431 256.663
R774 B.n546 B.n432 256.663
R775 B.n546 B.n433 256.663
R776 B.n546 B.n434 256.663
R777 B.n546 B.n435 256.663
R778 B.n546 B.n436 256.663
R779 B.n546 B.n437 256.663
R780 B.n546 B.n438 256.663
R781 B.n546 B.n439 256.663
R782 B.n546 B.n440 256.663
R783 B.n546 B.n441 256.663
R784 B.n546 B.n442 256.663
R785 B.n546 B.n443 256.663
R786 B.n546 B.n444 256.663
R787 B.n546 B.n445 256.663
R788 B.n449 B.t10 239.365
R789 B.n447 B.t21 239.365
R790 B.n172 B.t18 239.365
R791 B.n170 B.t14 239.365
R792 B.n449 B.t13 233.189
R793 B.n170 B.t16 233.189
R794 B.n447 B.t23 233.189
R795 B.n172 B.t19 233.189
R796 B.n552 B.n420 163.367
R797 B.n552 B.n414 163.367
R798 B.n560 B.n414 163.367
R799 B.n560 B.n412 163.367
R800 B.n564 B.n412 163.367
R801 B.n564 B.n406 163.367
R802 B.n572 B.n406 163.367
R803 B.n572 B.n404 163.367
R804 B.n576 B.n404 163.367
R805 B.n576 B.n398 163.367
R806 B.n584 B.n398 163.367
R807 B.n584 B.n396 163.367
R808 B.n588 B.n396 163.367
R809 B.n588 B.n390 163.367
R810 B.n596 B.n390 163.367
R811 B.n596 B.n388 163.367
R812 B.n600 B.n388 163.367
R813 B.n600 B.n382 163.367
R814 B.n608 B.n382 163.367
R815 B.n608 B.n380 163.367
R816 B.n612 B.n380 163.367
R817 B.n612 B.n374 163.367
R818 B.n621 B.n374 163.367
R819 B.n621 B.n372 163.367
R820 B.n625 B.n372 163.367
R821 B.n625 B.n367 163.367
R822 B.n633 B.n367 163.367
R823 B.n633 B.n365 163.367
R824 B.n637 B.n365 163.367
R825 B.n637 B.n359 163.367
R826 B.n645 B.n359 163.367
R827 B.n645 B.n357 163.367
R828 B.n649 B.n357 163.367
R829 B.n649 B.n351 163.367
R830 B.n658 B.n351 163.367
R831 B.n658 B.n349 163.367
R832 B.n662 B.n349 163.367
R833 B.n662 B.n344 163.367
R834 B.n670 B.n344 163.367
R835 B.n670 B.n342 163.367
R836 B.n674 B.n342 163.367
R837 B.n674 B.n336 163.367
R838 B.n682 B.n336 163.367
R839 B.n682 B.n334 163.367
R840 B.n686 B.n334 163.367
R841 B.n686 B.n328 163.367
R842 B.n694 B.n328 163.367
R843 B.n694 B.n326 163.367
R844 B.n698 B.n326 163.367
R845 B.n698 B.n320 163.367
R846 B.n706 B.n320 163.367
R847 B.n706 B.n318 163.367
R848 B.n710 B.n318 163.367
R849 B.n710 B.n312 163.367
R850 B.n718 B.n312 163.367
R851 B.n718 B.n310 163.367
R852 B.n722 B.n310 163.367
R853 B.n722 B.n304 163.367
R854 B.n730 B.n304 163.367
R855 B.n730 B.n302 163.367
R856 B.n734 B.n302 163.367
R857 B.n734 B.n296 163.367
R858 B.n742 B.n296 163.367
R859 B.n742 B.n294 163.367
R860 B.n746 B.n294 163.367
R861 B.n746 B.n288 163.367
R862 B.n754 B.n288 163.367
R863 B.n754 B.n286 163.367
R864 B.n758 B.n286 163.367
R865 B.n758 B.n280 163.367
R866 B.n766 B.n280 163.367
R867 B.n766 B.n278 163.367
R868 B.n770 B.n278 163.367
R869 B.n770 B.n272 163.367
R870 B.n779 B.n272 163.367
R871 B.n779 B.n270 163.367
R872 B.n783 B.n270 163.367
R873 B.n783 B.n2 163.367
R874 B.n1051 B.n2 163.367
R875 B.n1051 B.n3 163.367
R876 B.n1047 B.n3 163.367
R877 B.n1047 B.n9 163.367
R878 B.n1043 B.n9 163.367
R879 B.n1043 B.n11 163.367
R880 B.n1039 B.n11 163.367
R881 B.n1039 B.n16 163.367
R882 B.n1035 B.n16 163.367
R883 B.n1035 B.n18 163.367
R884 B.n1031 B.n18 163.367
R885 B.n1031 B.n23 163.367
R886 B.n1027 B.n23 163.367
R887 B.n1027 B.n25 163.367
R888 B.n1023 B.n25 163.367
R889 B.n1023 B.n30 163.367
R890 B.n1019 B.n30 163.367
R891 B.n1019 B.n32 163.367
R892 B.n1015 B.n32 163.367
R893 B.n1015 B.n37 163.367
R894 B.n1011 B.n37 163.367
R895 B.n1011 B.n39 163.367
R896 B.n1007 B.n39 163.367
R897 B.n1007 B.n44 163.367
R898 B.n1003 B.n44 163.367
R899 B.n1003 B.n46 163.367
R900 B.n999 B.n46 163.367
R901 B.n999 B.n51 163.367
R902 B.n995 B.n51 163.367
R903 B.n995 B.n53 163.367
R904 B.n991 B.n53 163.367
R905 B.n991 B.n58 163.367
R906 B.n987 B.n58 163.367
R907 B.n987 B.n60 163.367
R908 B.n983 B.n60 163.367
R909 B.n983 B.n65 163.367
R910 B.n979 B.n65 163.367
R911 B.n979 B.n67 163.367
R912 B.n975 B.n67 163.367
R913 B.n975 B.n72 163.367
R914 B.n971 B.n72 163.367
R915 B.n971 B.n74 163.367
R916 B.n967 B.n74 163.367
R917 B.n967 B.n78 163.367
R918 B.n963 B.n78 163.367
R919 B.n963 B.n80 163.367
R920 B.n959 B.n80 163.367
R921 B.n959 B.n86 163.367
R922 B.n955 B.n86 163.367
R923 B.n955 B.n88 163.367
R924 B.n951 B.n88 163.367
R925 B.n951 B.n93 163.367
R926 B.n947 B.n93 163.367
R927 B.n947 B.n95 163.367
R928 B.n943 B.n95 163.367
R929 B.n943 B.n99 163.367
R930 B.n939 B.n99 163.367
R931 B.n939 B.n101 163.367
R932 B.n935 B.n101 163.367
R933 B.n935 B.n107 163.367
R934 B.n931 B.n107 163.367
R935 B.n931 B.n109 163.367
R936 B.n927 B.n109 163.367
R937 B.n927 B.n114 163.367
R938 B.n923 B.n114 163.367
R939 B.n923 B.n116 163.367
R940 B.n919 B.n116 163.367
R941 B.n919 B.n121 163.367
R942 B.n915 B.n121 163.367
R943 B.n915 B.n123 163.367
R944 B.n911 B.n123 163.367
R945 B.n911 B.n128 163.367
R946 B.n907 B.n128 163.367
R947 B.n907 B.n130 163.367
R948 B.n903 B.n130 163.367
R949 B.n903 B.n135 163.367
R950 B.n899 B.n135 163.367
R951 B.n899 B.n137 163.367
R952 B.n895 B.n137 163.367
R953 B.n895 B.n142 163.367
R954 B.n545 B.n422 163.367
R955 B.n545 B.n446 163.367
R956 B.n541 B.n540 163.367
R957 B.n537 B.n536 163.367
R958 B.n533 B.n532 163.367
R959 B.n529 B.n528 163.367
R960 B.n525 B.n524 163.367
R961 B.n521 B.n520 163.367
R962 B.n517 B.n516 163.367
R963 B.n513 B.n512 163.367
R964 B.n508 B.n507 163.367
R965 B.n504 B.n503 163.367
R966 B.n500 B.n499 163.367
R967 B.n496 B.n495 163.367
R968 B.n492 B.n491 163.367
R969 B.n488 B.n487 163.367
R970 B.n484 B.n483 163.367
R971 B.n480 B.n479 163.367
R972 B.n476 B.n475 163.367
R973 B.n472 B.n471 163.367
R974 B.n468 B.n467 163.367
R975 B.n464 B.n463 163.367
R976 B.n460 B.n459 163.367
R977 B.n456 B.n455 163.367
R978 B.n554 B.n418 163.367
R979 B.n554 B.n416 163.367
R980 B.n558 B.n416 163.367
R981 B.n558 B.n410 163.367
R982 B.n566 B.n410 163.367
R983 B.n566 B.n408 163.367
R984 B.n570 B.n408 163.367
R985 B.n570 B.n402 163.367
R986 B.n578 B.n402 163.367
R987 B.n578 B.n400 163.367
R988 B.n582 B.n400 163.367
R989 B.n582 B.n394 163.367
R990 B.n590 B.n394 163.367
R991 B.n590 B.n392 163.367
R992 B.n594 B.n392 163.367
R993 B.n594 B.n386 163.367
R994 B.n602 B.n386 163.367
R995 B.n602 B.n384 163.367
R996 B.n606 B.n384 163.367
R997 B.n606 B.n378 163.367
R998 B.n614 B.n378 163.367
R999 B.n614 B.n376 163.367
R1000 B.n618 B.n376 163.367
R1001 B.n618 B.n371 163.367
R1002 B.n627 B.n371 163.367
R1003 B.n627 B.n369 163.367
R1004 B.n631 B.n369 163.367
R1005 B.n631 B.n363 163.367
R1006 B.n639 B.n363 163.367
R1007 B.n639 B.n361 163.367
R1008 B.n643 B.n361 163.367
R1009 B.n643 B.n355 163.367
R1010 B.n651 B.n355 163.367
R1011 B.n651 B.n353 163.367
R1012 B.n655 B.n353 163.367
R1013 B.n655 B.n348 163.367
R1014 B.n664 B.n348 163.367
R1015 B.n664 B.n346 163.367
R1016 B.n668 B.n346 163.367
R1017 B.n668 B.n340 163.367
R1018 B.n676 B.n340 163.367
R1019 B.n676 B.n338 163.367
R1020 B.n680 B.n338 163.367
R1021 B.n680 B.n332 163.367
R1022 B.n688 B.n332 163.367
R1023 B.n688 B.n330 163.367
R1024 B.n692 B.n330 163.367
R1025 B.n692 B.n324 163.367
R1026 B.n700 B.n324 163.367
R1027 B.n700 B.n322 163.367
R1028 B.n704 B.n322 163.367
R1029 B.n704 B.n316 163.367
R1030 B.n712 B.n316 163.367
R1031 B.n712 B.n314 163.367
R1032 B.n716 B.n314 163.367
R1033 B.n716 B.n308 163.367
R1034 B.n724 B.n308 163.367
R1035 B.n724 B.n306 163.367
R1036 B.n728 B.n306 163.367
R1037 B.n728 B.n300 163.367
R1038 B.n736 B.n300 163.367
R1039 B.n736 B.n298 163.367
R1040 B.n740 B.n298 163.367
R1041 B.n740 B.n292 163.367
R1042 B.n748 B.n292 163.367
R1043 B.n748 B.n290 163.367
R1044 B.n752 B.n290 163.367
R1045 B.n752 B.n284 163.367
R1046 B.n760 B.n284 163.367
R1047 B.n760 B.n282 163.367
R1048 B.n764 B.n282 163.367
R1049 B.n764 B.n276 163.367
R1050 B.n772 B.n276 163.367
R1051 B.n772 B.n274 163.367
R1052 B.n777 B.n274 163.367
R1053 B.n777 B.n268 163.367
R1054 B.n785 B.n268 163.367
R1055 B.n786 B.n785 163.367
R1056 B.n786 B.n5 163.367
R1057 B.n6 B.n5 163.367
R1058 B.n7 B.n6 163.367
R1059 B.n791 B.n7 163.367
R1060 B.n791 B.n12 163.367
R1061 B.n13 B.n12 163.367
R1062 B.n14 B.n13 163.367
R1063 B.n796 B.n14 163.367
R1064 B.n796 B.n19 163.367
R1065 B.n20 B.n19 163.367
R1066 B.n21 B.n20 163.367
R1067 B.n801 B.n21 163.367
R1068 B.n801 B.n26 163.367
R1069 B.n27 B.n26 163.367
R1070 B.n28 B.n27 163.367
R1071 B.n806 B.n28 163.367
R1072 B.n806 B.n33 163.367
R1073 B.n34 B.n33 163.367
R1074 B.n35 B.n34 163.367
R1075 B.n811 B.n35 163.367
R1076 B.n811 B.n40 163.367
R1077 B.n41 B.n40 163.367
R1078 B.n42 B.n41 163.367
R1079 B.n816 B.n42 163.367
R1080 B.n816 B.n47 163.367
R1081 B.n48 B.n47 163.367
R1082 B.n49 B.n48 163.367
R1083 B.n821 B.n49 163.367
R1084 B.n821 B.n54 163.367
R1085 B.n55 B.n54 163.367
R1086 B.n56 B.n55 163.367
R1087 B.n826 B.n56 163.367
R1088 B.n826 B.n61 163.367
R1089 B.n62 B.n61 163.367
R1090 B.n63 B.n62 163.367
R1091 B.n831 B.n63 163.367
R1092 B.n831 B.n68 163.367
R1093 B.n69 B.n68 163.367
R1094 B.n70 B.n69 163.367
R1095 B.n836 B.n70 163.367
R1096 B.n836 B.n75 163.367
R1097 B.n76 B.n75 163.367
R1098 B.n77 B.n76 163.367
R1099 B.n841 B.n77 163.367
R1100 B.n841 B.n82 163.367
R1101 B.n83 B.n82 163.367
R1102 B.n84 B.n83 163.367
R1103 B.n846 B.n84 163.367
R1104 B.n846 B.n89 163.367
R1105 B.n90 B.n89 163.367
R1106 B.n91 B.n90 163.367
R1107 B.n851 B.n91 163.367
R1108 B.n851 B.n96 163.367
R1109 B.n97 B.n96 163.367
R1110 B.n98 B.n97 163.367
R1111 B.n856 B.n98 163.367
R1112 B.n856 B.n103 163.367
R1113 B.n104 B.n103 163.367
R1114 B.n105 B.n104 163.367
R1115 B.n861 B.n105 163.367
R1116 B.n861 B.n110 163.367
R1117 B.n111 B.n110 163.367
R1118 B.n112 B.n111 163.367
R1119 B.n866 B.n112 163.367
R1120 B.n866 B.n117 163.367
R1121 B.n118 B.n117 163.367
R1122 B.n119 B.n118 163.367
R1123 B.n871 B.n119 163.367
R1124 B.n871 B.n124 163.367
R1125 B.n125 B.n124 163.367
R1126 B.n126 B.n125 163.367
R1127 B.n876 B.n126 163.367
R1128 B.n876 B.n131 163.367
R1129 B.n132 B.n131 163.367
R1130 B.n133 B.n132 163.367
R1131 B.n881 B.n133 163.367
R1132 B.n881 B.n138 163.367
R1133 B.n139 B.n138 163.367
R1134 B.n140 B.n139 163.367
R1135 B.n169 B.n140 163.367
R1136 B.n175 B.n144 163.367
R1137 B.n179 B.n178 163.367
R1138 B.n183 B.n182 163.367
R1139 B.n187 B.n186 163.367
R1140 B.n191 B.n190 163.367
R1141 B.n195 B.n194 163.367
R1142 B.n199 B.n198 163.367
R1143 B.n203 B.n202 163.367
R1144 B.n207 B.n206 163.367
R1145 B.n211 B.n210 163.367
R1146 B.n215 B.n214 163.367
R1147 B.n219 B.n218 163.367
R1148 B.n223 B.n222 163.367
R1149 B.n227 B.n226 163.367
R1150 B.n232 B.n231 163.367
R1151 B.n236 B.n235 163.367
R1152 B.n240 B.n239 163.367
R1153 B.n244 B.n243 163.367
R1154 B.n248 B.n247 163.367
R1155 B.n252 B.n251 163.367
R1156 B.n256 B.n255 163.367
R1157 B.n260 B.n259 163.367
R1158 B.n264 B.n263 163.367
R1159 B.n888 B.n168 163.367
R1160 B.n450 B.t12 155.225
R1161 B.n171 B.t17 155.225
R1162 B.n448 B.t22 155.225
R1163 B.n173 B.t20 155.225
R1164 B.n546 B.n419 141.326
R1165 B.n889 B.n141 141.326
R1166 B.n450 B.n449 77.9641
R1167 B.n448 B.n447 77.9641
R1168 B.n173 B.n172 77.9641
R1169 B.n171 B.n170 77.9641
R1170 B.n553 B.n419 75.6707
R1171 B.n553 B.n415 75.6707
R1172 B.n559 B.n415 75.6707
R1173 B.n559 B.n411 75.6707
R1174 B.n565 B.n411 75.6707
R1175 B.n565 B.n407 75.6707
R1176 B.n571 B.n407 75.6707
R1177 B.n571 B.n403 75.6707
R1178 B.n577 B.n403 75.6707
R1179 B.n583 B.n399 75.6707
R1180 B.n583 B.n395 75.6707
R1181 B.n589 B.n395 75.6707
R1182 B.n589 B.n391 75.6707
R1183 B.n595 B.n391 75.6707
R1184 B.n595 B.n387 75.6707
R1185 B.n601 B.n387 75.6707
R1186 B.n601 B.n383 75.6707
R1187 B.n607 B.n383 75.6707
R1188 B.n607 B.n379 75.6707
R1189 B.n613 B.n379 75.6707
R1190 B.n613 B.n375 75.6707
R1191 B.n620 B.n375 75.6707
R1192 B.n620 B.n619 75.6707
R1193 B.n626 B.n368 75.6707
R1194 B.n632 B.n368 75.6707
R1195 B.n632 B.n364 75.6707
R1196 B.n638 B.n364 75.6707
R1197 B.n638 B.n360 75.6707
R1198 B.n644 B.n360 75.6707
R1199 B.n644 B.n356 75.6707
R1200 B.n650 B.n356 75.6707
R1201 B.n650 B.n352 75.6707
R1202 B.n657 B.n352 75.6707
R1203 B.n657 B.n656 75.6707
R1204 B.n663 B.n345 75.6707
R1205 B.n669 B.n345 75.6707
R1206 B.n669 B.n341 75.6707
R1207 B.n675 B.n341 75.6707
R1208 B.n675 B.n337 75.6707
R1209 B.n681 B.n337 75.6707
R1210 B.n681 B.n333 75.6707
R1211 B.n687 B.n333 75.6707
R1212 B.n687 B.n329 75.6707
R1213 B.n693 B.n329 75.6707
R1214 B.n699 B.n325 75.6707
R1215 B.n699 B.n321 75.6707
R1216 B.n705 B.n321 75.6707
R1217 B.n705 B.n317 75.6707
R1218 B.n711 B.n317 75.6707
R1219 B.n711 B.n313 75.6707
R1220 B.n717 B.n313 75.6707
R1221 B.n717 B.n309 75.6707
R1222 B.n723 B.n309 75.6707
R1223 B.n723 B.n305 75.6707
R1224 B.n729 B.n305 75.6707
R1225 B.n735 B.n301 75.6707
R1226 B.n735 B.n297 75.6707
R1227 B.n741 B.n297 75.6707
R1228 B.n741 B.n293 75.6707
R1229 B.n747 B.n293 75.6707
R1230 B.n747 B.n289 75.6707
R1231 B.n753 B.n289 75.6707
R1232 B.n753 B.n285 75.6707
R1233 B.n759 B.n285 75.6707
R1234 B.n759 B.n281 75.6707
R1235 B.n765 B.n281 75.6707
R1236 B.n771 B.n277 75.6707
R1237 B.n771 B.n273 75.6707
R1238 B.n778 B.n273 75.6707
R1239 B.n778 B.n269 75.6707
R1240 B.n784 B.n269 75.6707
R1241 B.n784 B.n4 75.6707
R1242 B.n1050 B.n4 75.6707
R1243 B.n1050 B.n1049 75.6707
R1244 B.n1049 B.n1048 75.6707
R1245 B.n1048 B.n8 75.6707
R1246 B.n1042 B.n8 75.6707
R1247 B.n1042 B.n1041 75.6707
R1248 B.n1041 B.n1040 75.6707
R1249 B.n1040 B.n15 75.6707
R1250 B.n1034 B.n1033 75.6707
R1251 B.n1033 B.n1032 75.6707
R1252 B.n1032 B.n22 75.6707
R1253 B.n1026 B.n22 75.6707
R1254 B.n1026 B.n1025 75.6707
R1255 B.n1025 B.n1024 75.6707
R1256 B.n1024 B.n29 75.6707
R1257 B.n1018 B.n29 75.6707
R1258 B.n1018 B.n1017 75.6707
R1259 B.n1017 B.n1016 75.6707
R1260 B.n1016 B.n36 75.6707
R1261 B.n1010 B.n1009 75.6707
R1262 B.n1009 B.n1008 75.6707
R1263 B.n1008 B.n43 75.6707
R1264 B.n1002 B.n43 75.6707
R1265 B.n1002 B.n1001 75.6707
R1266 B.n1001 B.n1000 75.6707
R1267 B.n1000 B.n50 75.6707
R1268 B.n994 B.n50 75.6707
R1269 B.n994 B.n993 75.6707
R1270 B.n993 B.n992 75.6707
R1271 B.n992 B.n57 75.6707
R1272 B.n986 B.n985 75.6707
R1273 B.n985 B.n984 75.6707
R1274 B.n984 B.n64 75.6707
R1275 B.n978 B.n64 75.6707
R1276 B.n978 B.n977 75.6707
R1277 B.n977 B.n976 75.6707
R1278 B.n976 B.n71 75.6707
R1279 B.n970 B.n71 75.6707
R1280 B.n970 B.n969 75.6707
R1281 B.n969 B.n968 75.6707
R1282 B.n962 B.n81 75.6707
R1283 B.n962 B.n961 75.6707
R1284 B.n961 B.n960 75.6707
R1285 B.n960 B.n85 75.6707
R1286 B.n954 B.n85 75.6707
R1287 B.n954 B.n953 75.6707
R1288 B.n953 B.n952 75.6707
R1289 B.n952 B.n92 75.6707
R1290 B.n946 B.n92 75.6707
R1291 B.n946 B.n945 75.6707
R1292 B.n945 B.n944 75.6707
R1293 B.n938 B.n102 75.6707
R1294 B.n938 B.n937 75.6707
R1295 B.n937 B.n936 75.6707
R1296 B.n936 B.n106 75.6707
R1297 B.n930 B.n106 75.6707
R1298 B.n930 B.n929 75.6707
R1299 B.n929 B.n928 75.6707
R1300 B.n928 B.n113 75.6707
R1301 B.n922 B.n113 75.6707
R1302 B.n922 B.n921 75.6707
R1303 B.n921 B.n920 75.6707
R1304 B.n920 B.n120 75.6707
R1305 B.n914 B.n120 75.6707
R1306 B.n914 B.n913 75.6707
R1307 B.n912 B.n127 75.6707
R1308 B.n906 B.n127 75.6707
R1309 B.n906 B.n905 75.6707
R1310 B.n905 B.n904 75.6707
R1311 B.n904 B.n134 75.6707
R1312 B.n898 B.n134 75.6707
R1313 B.n898 B.n897 75.6707
R1314 B.n897 B.n896 75.6707
R1315 B.n896 B.n141 75.6707
R1316 B.n663 B.t0 74.5579
R1317 B.n968 B.t1 74.5579
R1318 B.n548 B.n547 71.676
R1319 B.n446 B.n423 71.676
R1320 B.n540 B.n424 71.676
R1321 B.n536 B.n425 71.676
R1322 B.n532 B.n426 71.676
R1323 B.n528 B.n427 71.676
R1324 B.n524 B.n428 71.676
R1325 B.n520 B.n429 71.676
R1326 B.n516 B.n430 71.676
R1327 B.n512 B.n431 71.676
R1328 B.n507 B.n432 71.676
R1329 B.n503 B.n433 71.676
R1330 B.n499 B.n434 71.676
R1331 B.n495 B.n435 71.676
R1332 B.n491 B.n436 71.676
R1333 B.n487 B.n437 71.676
R1334 B.n483 B.n438 71.676
R1335 B.n479 B.n439 71.676
R1336 B.n475 B.n440 71.676
R1337 B.n471 B.n441 71.676
R1338 B.n467 B.n442 71.676
R1339 B.n463 B.n443 71.676
R1340 B.n459 B.n444 71.676
R1341 B.n455 B.n445 71.676
R1342 B.n891 B.n890 71.676
R1343 B.n175 B.n145 71.676
R1344 B.n179 B.n146 71.676
R1345 B.n183 B.n147 71.676
R1346 B.n187 B.n148 71.676
R1347 B.n191 B.n149 71.676
R1348 B.n195 B.n150 71.676
R1349 B.n199 B.n151 71.676
R1350 B.n203 B.n152 71.676
R1351 B.n207 B.n153 71.676
R1352 B.n211 B.n154 71.676
R1353 B.n215 B.n155 71.676
R1354 B.n219 B.n156 71.676
R1355 B.n223 B.n157 71.676
R1356 B.n227 B.n158 71.676
R1357 B.n232 B.n159 71.676
R1358 B.n236 B.n160 71.676
R1359 B.n240 B.n161 71.676
R1360 B.n244 B.n162 71.676
R1361 B.n248 B.n163 71.676
R1362 B.n252 B.n164 71.676
R1363 B.n256 B.n165 71.676
R1364 B.n260 B.n166 71.676
R1365 B.n264 B.n167 71.676
R1366 B.n168 B.n167 71.676
R1367 B.n263 B.n166 71.676
R1368 B.n259 B.n165 71.676
R1369 B.n255 B.n164 71.676
R1370 B.n251 B.n163 71.676
R1371 B.n247 B.n162 71.676
R1372 B.n243 B.n161 71.676
R1373 B.n239 B.n160 71.676
R1374 B.n235 B.n159 71.676
R1375 B.n231 B.n158 71.676
R1376 B.n226 B.n157 71.676
R1377 B.n222 B.n156 71.676
R1378 B.n218 B.n155 71.676
R1379 B.n214 B.n154 71.676
R1380 B.n210 B.n153 71.676
R1381 B.n206 B.n152 71.676
R1382 B.n202 B.n151 71.676
R1383 B.n198 B.n150 71.676
R1384 B.n194 B.n149 71.676
R1385 B.n190 B.n148 71.676
R1386 B.n186 B.n147 71.676
R1387 B.n182 B.n146 71.676
R1388 B.n178 B.n145 71.676
R1389 B.n890 B.n144 71.676
R1390 B.n547 B.n422 71.676
R1391 B.n541 B.n423 71.676
R1392 B.n537 B.n424 71.676
R1393 B.n533 B.n425 71.676
R1394 B.n529 B.n426 71.676
R1395 B.n525 B.n427 71.676
R1396 B.n521 B.n428 71.676
R1397 B.n517 B.n429 71.676
R1398 B.n513 B.n430 71.676
R1399 B.n508 B.n431 71.676
R1400 B.n504 B.n432 71.676
R1401 B.n500 B.n433 71.676
R1402 B.n496 B.n434 71.676
R1403 B.n492 B.n435 71.676
R1404 B.n488 B.n436 71.676
R1405 B.n484 B.n437 71.676
R1406 B.n480 B.n438 71.676
R1407 B.n476 B.n439 71.676
R1408 B.n472 B.n440 71.676
R1409 B.n468 B.n441 71.676
R1410 B.n464 B.n442 71.676
R1411 B.n460 B.n443 71.676
R1412 B.n456 B.n444 71.676
R1413 B.n452 B.n445 71.676
R1414 B.t11 B.n399 63.4299
R1415 B.n693 B.t8 63.4299
R1416 B.n986 B.t7 63.4299
R1417 B.n913 B.t15 63.4299
R1418 B.n626 B.t6 61.2043
R1419 B.n944 B.t5 61.2043
R1420 B.n451 B.n450 59.5399
R1421 B.n510 B.n448 59.5399
R1422 B.n174 B.n173 59.5399
R1423 B.n229 B.n171 59.5399
R1424 B.n729 B.t2 50.0764
R1425 B.n1010 B.t3 50.0764
R1426 B.t9 B.n277 38.9484
R1427 B.t4 B.n15 38.9484
R1428 B.n765 B.t9 36.7228
R1429 B.n1034 B.t4 36.7228
R1430 B.n893 B.n892 34.8103
R1431 B.n887 B.n886 34.8103
R1432 B.n453 B.n417 34.8103
R1433 B.n550 B.n549 34.8103
R1434 B.t2 B.n301 25.5948
R1435 B.t3 B.n36 25.5948
R1436 B B.n1052 18.0485
R1437 B.n619 B.t6 14.4669
R1438 B.n102 B.t5 14.4669
R1439 B.n577 B.t11 12.2413
R1440 B.t8 B.n325 12.2413
R1441 B.t7 B.n57 12.2413
R1442 B.t15 B.n912 12.2413
R1443 B.n892 B.n143 10.6151
R1444 B.n176 B.n143 10.6151
R1445 B.n177 B.n176 10.6151
R1446 B.n180 B.n177 10.6151
R1447 B.n181 B.n180 10.6151
R1448 B.n184 B.n181 10.6151
R1449 B.n185 B.n184 10.6151
R1450 B.n188 B.n185 10.6151
R1451 B.n189 B.n188 10.6151
R1452 B.n192 B.n189 10.6151
R1453 B.n193 B.n192 10.6151
R1454 B.n196 B.n193 10.6151
R1455 B.n197 B.n196 10.6151
R1456 B.n200 B.n197 10.6151
R1457 B.n201 B.n200 10.6151
R1458 B.n204 B.n201 10.6151
R1459 B.n205 B.n204 10.6151
R1460 B.n208 B.n205 10.6151
R1461 B.n209 B.n208 10.6151
R1462 B.n213 B.n212 10.6151
R1463 B.n216 B.n213 10.6151
R1464 B.n217 B.n216 10.6151
R1465 B.n220 B.n217 10.6151
R1466 B.n221 B.n220 10.6151
R1467 B.n224 B.n221 10.6151
R1468 B.n225 B.n224 10.6151
R1469 B.n228 B.n225 10.6151
R1470 B.n233 B.n230 10.6151
R1471 B.n234 B.n233 10.6151
R1472 B.n237 B.n234 10.6151
R1473 B.n238 B.n237 10.6151
R1474 B.n241 B.n238 10.6151
R1475 B.n242 B.n241 10.6151
R1476 B.n245 B.n242 10.6151
R1477 B.n246 B.n245 10.6151
R1478 B.n249 B.n246 10.6151
R1479 B.n250 B.n249 10.6151
R1480 B.n253 B.n250 10.6151
R1481 B.n254 B.n253 10.6151
R1482 B.n257 B.n254 10.6151
R1483 B.n258 B.n257 10.6151
R1484 B.n261 B.n258 10.6151
R1485 B.n262 B.n261 10.6151
R1486 B.n265 B.n262 10.6151
R1487 B.n266 B.n265 10.6151
R1488 B.n887 B.n266 10.6151
R1489 B.n555 B.n417 10.6151
R1490 B.n556 B.n555 10.6151
R1491 B.n557 B.n556 10.6151
R1492 B.n557 B.n409 10.6151
R1493 B.n567 B.n409 10.6151
R1494 B.n568 B.n567 10.6151
R1495 B.n569 B.n568 10.6151
R1496 B.n569 B.n401 10.6151
R1497 B.n579 B.n401 10.6151
R1498 B.n580 B.n579 10.6151
R1499 B.n581 B.n580 10.6151
R1500 B.n581 B.n393 10.6151
R1501 B.n591 B.n393 10.6151
R1502 B.n592 B.n591 10.6151
R1503 B.n593 B.n592 10.6151
R1504 B.n593 B.n385 10.6151
R1505 B.n603 B.n385 10.6151
R1506 B.n604 B.n603 10.6151
R1507 B.n605 B.n604 10.6151
R1508 B.n605 B.n377 10.6151
R1509 B.n615 B.n377 10.6151
R1510 B.n616 B.n615 10.6151
R1511 B.n617 B.n616 10.6151
R1512 B.n617 B.n370 10.6151
R1513 B.n628 B.n370 10.6151
R1514 B.n629 B.n628 10.6151
R1515 B.n630 B.n629 10.6151
R1516 B.n630 B.n362 10.6151
R1517 B.n640 B.n362 10.6151
R1518 B.n641 B.n640 10.6151
R1519 B.n642 B.n641 10.6151
R1520 B.n642 B.n354 10.6151
R1521 B.n652 B.n354 10.6151
R1522 B.n653 B.n652 10.6151
R1523 B.n654 B.n653 10.6151
R1524 B.n654 B.n347 10.6151
R1525 B.n665 B.n347 10.6151
R1526 B.n666 B.n665 10.6151
R1527 B.n667 B.n666 10.6151
R1528 B.n667 B.n339 10.6151
R1529 B.n677 B.n339 10.6151
R1530 B.n678 B.n677 10.6151
R1531 B.n679 B.n678 10.6151
R1532 B.n679 B.n331 10.6151
R1533 B.n689 B.n331 10.6151
R1534 B.n690 B.n689 10.6151
R1535 B.n691 B.n690 10.6151
R1536 B.n691 B.n323 10.6151
R1537 B.n701 B.n323 10.6151
R1538 B.n702 B.n701 10.6151
R1539 B.n703 B.n702 10.6151
R1540 B.n703 B.n315 10.6151
R1541 B.n713 B.n315 10.6151
R1542 B.n714 B.n713 10.6151
R1543 B.n715 B.n714 10.6151
R1544 B.n715 B.n307 10.6151
R1545 B.n725 B.n307 10.6151
R1546 B.n726 B.n725 10.6151
R1547 B.n727 B.n726 10.6151
R1548 B.n727 B.n299 10.6151
R1549 B.n737 B.n299 10.6151
R1550 B.n738 B.n737 10.6151
R1551 B.n739 B.n738 10.6151
R1552 B.n739 B.n291 10.6151
R1553 B.n749 B.n291 10.6151
R1554 B.n750 B.n749 10.6151
R1555 B.n751 B.n750 10.6151
R1556 B.n751 B.n283 10.6151
R1557 B.n761 B.n283 10.6151
R1558 B.n762 B.n761 10.6151
R1559 B.n763 B.n762 10.6151
R1560 B.n763 B.n275 10.6151
R1561 B.n773 B.n275 10.6151
R1562 B.n774 B.n773 10.6151
R1563 B.n776 B.n774 10.6151
R1564 B.n776 B.n775 10.6151
R1565 B.n775 B.n267 10.6151
R1566 B.n787 B.n267 10.6151
R1567 B.n788 B.n787 10.6151
R1568 B.n789 B.n788 10.6151
R1569 B.n790 B.n789 10.6151
R1570 B.n792 B.n790 10.6151
R1571 B.n793 B.n792 10.6151
R1572 B.n794 B.n793 10.6151
R1573 B.n795 B.n794 10.6151
R1574 B.n797 B.n795 10.6151
R1575 B.n798 B.n797 10.6151
R1576 B.n799 B.n798 10.6151
R1577 B.n800 B.n799 10.6151
R1578 B.n802 B.n800 10.6151
R1579 B.n803 B.n802 10.6151
R1580 B.n804 B.n803 10.6151
R1581 B.n805 B.n804 10.6151
R1582 B.n807 B.n805 10.6151
R1583 B.n808 B.n807 10.6151
R1584 B.n809 B.n808 10.6151
R1585 B.n810 B.n809 10.6151
R1586 B.n812 B.n810 10.6151
R1587 B.n813 B.n812 10.6151
R1588 B.n814 B.n813 10.6151
R1589 B.n815 B.n814 10.6151
R1590 B.n817 B.n815 10.6151
R1591 B.n818 B.n817 10.6151
R1592 B.n819 B.n818 10.6151
R1593 B.n820 B.n819 10.6151
R1594 B.n822 B.n820 10.6151
R1595 B.n823 B.n822 10.6151
R1596 B.n824 B.n823 10.6151
R1597 B.n825 B.n824 10.6151
R1598 B.n827 B.n825 10.6151
R1599 B.n828 B.n827 10.6151
R1600 B.n829 B.n828 10.6151
R1601 B.n830 B.n829 10.6151
R1602 B.n832 B.n830 10.6151
R1603 B.n833 B.n832 10.6151
R1604 B.n834 B.n833 10.6151
R1605 B.n835 B.n834 10.6151
R1606 B.n837 B.n835 10.6151
R1607 B.n838 B.n837 10.6151
R1608 B.n839 B.n838 10.6151
R1609 B.n840 B.n839 10.6151
R1610 B.n842 B.n840 10.6151
R1611 B.n843 B.n842 10.6151
R1612 B.n844 B.n843 10.6151
R1613 B.n845 B.n844 10.6151
R1614 B.n847 B.n845 10.6151
R1615 B.n848 B.n847 10.6151
R1616 B.n849 B.n848 10.6151
R1617 B.n850 B.n849 10.6151
R1618 B.n852 B.n850 10.6151
R1619 B.n853 B.n852 10.6151
R1620 B.n854 B.n853 10.6151
R1621 B.n855 B.n854 10.6151
R1622 B.n857 B.n855 10.6151
R1623 B.n858 B.n857 10.6151
R1624 B.n859 B.n858 10.6151
R1625 B.n860 B.n859 10.6151
R1626 B.n862 B.n860 10.6151
R1627 B.n863 B.n862 10.6151
R1628 B.n864 B.n863 10.6151
R1629 B.n865 B.n864 10.6151
R1630 B.n867 B.n865 10.6151
R1631 B.n868 B.n867 10.6151
R1632 B.n869 B.n868 10.6151
R1633 B.n870 B.n869 10.6151
R1634 B.n872 B.n870 10.6151
R1635 B.n873 B.n872 10.6151
R1636 B.n874 B.n873 10.6151
R1637 B.n875 B.n874 10.6151
R1638 B.n877 B.n875 10.6151
R1639 B.n878 B.n877 10.6151
R1640 B.n879 B.n878 10.6151
R1641 B.n880 B.n879 10.6151
R1642 B.n882 B.n880 10.6151
R1643 B.n883 B.n882 10.6151
R1644 B.n884 B.n883 10.6151
R1645 B.n885 B.n884 10.6151
R1646 B.n886 B.n885 10.6151
R1647 B.n549 B.n421 10.6151
R1648 B.n544 B.n421 10.6151
R1649 B.n544 B.n543 10.6151
R1650 B.n543 B.n542 10.6151
R1651 B.n542 B.n539 10.6151
R1652 B.n539 B.n538 10.6151
R1653 B.n538 B.n535 10.6151
R1654 B.n535 B.n534 10.6151
R1655 B.n534 B.n531 10.6151
R1656 B.n531 B.n530 10.6151
R1657 B.n530 B.n527 10.6151
R1658 B.n527 B.n526 10.6151
R1659 B.n526 B.n523 10.6151
R1660 B.n523 B.n522 10.6151
R1661 B.n522 B.n519 10.6151
R1662 B.n519 B.n518 10.6151
R1663 B.n518 B.n515 10.6151
R1664 B.n515 B.n514 10.6151
R1665 B.n514 B.n511 10.6151
R1666 B.n509 B.n506 10.6151
R1667 B.n506 B.n505 10.6151
R1668 B.n505 B.n502 10.6151
R1669 B.n502 B.n501 10.6151
R1670 B.n501 B.n498 10.6151
R1671 B.n498 B.n497 10.6151
R1672 B.n497 B.n494 10.6151
R1673 B.n494 B.n493 10.6151
R1674 B.n490 B.n489 10.6151
R1675 B.n489 B.n486 10.6151
R1676 B.n486 B.n485 10.6151
R1677 B.n485 B.n482 10.6151
R1678 B.n482 B.n481 10.6151
R1679 B.n481 B.n478 10.6151
R1680 B.n478 B.n477 10.6151
R1681 B.n477 B.n474 10.6151
R1682 B.n474 B.n473 10.6151
R1683 B.n473 B.n470 10.6151
R1684 B.n470 B.n469 10.6151
R1685 B.n469 B.n466 10.6151
R1686 B.n466 B.n465 10.6151
R1687 B.n465 B.n462 10.6151
R1688 B.n462 B.n461 10.6151
R1689 B.n461 B.n458 10.6151
R1690 B.n458 B.n457 10.6151
R1691 B.n457 B.n454 10.6151
R1692 B.n454 B.n453 10.6151
R1693 B.n551 B.n550 10.6151
R1694 B.n551 B.n413 10.6151
R1695 B.n561 B.n413 10.6151
R1696 B.n562 B.n561 10.6151
R1697 B.n563 B.n562 10.6151
R1698 B.n563 B.n405 10.6151
R1699 B.n573 B.n405 10.6151
R1700 B.n574 B.n573 10.6151
R1701 B.n575 B.n574 10.6151
R1702 B.n575 B.n397 10.6151
R1703 B.n585 B.n397 10.6151
R1704 B.n586 B.n585 10.6151
R1705 B.n587 B.n586 10.6151
R1706 B.n587 B.n389 10.6151
R1707 B.n597 B.n389 10.6151
R1708 B.n598 B.n597 10.6151
R1709 B.n599 B.n598 10.6151
R1710 B.n599 B.n381 10.6151
R1711 B.n609 B.n381 10.6151
R1712 B.n610 B.n609 10.6151
R1713 B.n611 B.n610 10.6151
R1714 B.n611 B.n373 10.6151
R1715 B.n622 B.n373 10.6151
R1716 B.n623 B.n622 10.6151
R1717 B.n624 B.n623 10.6151
R1718 B.n624 B.n366 10.6151
R1719 B.n634 B.n366 10.6151
R1720 B.n635 B.n634 10.6151
R1721 B.n636 B.n635 10.6151
R1722 B.n636 B.n358 10.6151
R1723 B.n646 B.n358 10.6151
R1724 B.n647 B.n646 10.6151
R1725 B.n648 B.n647 10.6151
R1726 B.n648 B.n350 10.6151
R1727 B.n659 B.n350 10.6151
R1728 B.n660 B.n659 10.6151
R1729 B.n661 B.n660 10.6151
R1730 B.n661 B.n343 10.6151
R1731 B.n671 B.n343 10.6151
R1732 B.n672 B.n671 10.6151
R1733 B.n673 B.n672 10.6151
R1734 B.n673 B.n335 10.6151
R1735 B.n683 B.n335 10.6151
R1736 B.n684 B.n683 10.6151
R1737 B.n685 B.n684 10.6151
R1738 B.n685 B.n327 10.6151
R1739 B.n695 B.n327 10.6151
R1740 B.n696 B.n695 10.6151
R1741 B.n697 B.n696 10.6151
R1742 B.n697 B.n319 10.6151
R1743 B.n707 B.n319 10.6151
R1744 B.n708 B.n707 10.6151
R1745 B.n709 B.n708 10.6151
R1746 B.n709 B.n311 10.6151
R1747 B.n719 B.n311 10.6151
R1748 B.n720 B.n719 10.6151
R1749 B.n721 B.n720 10.6151
R1750 B.n721 B.n303 10.6151
R1751 B.n731 B.n303 10.6151
R1752 B.n732 B.n731 10.6151
R1753 B.n733 B.n732 10.6151
R1754 B.n733 B.n295 10.6151
R1755 B.n743 B.n295 10.6151
R1756 B.n744 B.n743 10.6151
R1757 B.n745 B.n744 10.6151
R1758 B.n745 B.n287 10.6151
R1759 B.n755 B.n287 10.6151
R1760 B.n756 B.n755 10.6151
R1761 B.n757 B.n756 10.6151
R1762 B.n757 B.n279 10.6151
R1763 B.n767 B.n279 10.6151
R1764 B.n768 B.n767 10.6151
R1765 B.n769 B.n768 10.6151
R1766 B.n769 B.n271 10.6151
R1767 B.n780 B.n271 10.6151
R1768 B.n781 B.n780 10.6151
R1769 B.n782 B.n781 10.6151
R1770 B.n782 B.n0 10.6151
R1771 B.n1046 B.n1 10.6151
R1772 B.n1046 B.n1045 10.6151
R1773 B.n1045 B.n1044 10.6151
R1774 B.n1044 B.n10 10.6151
R1775 B.n1038 B.n10 10.6151
R1776 B.n1038 B.n1037 10.6151
R1777 B.n1037 B.n1036 10.6151
R1778 B.n1036 B.n17 10.6151
R1779 B.n1030 B.n17 10.6151
R1780 B.n1030 B.n1029 10.6151
R1781 B.n1029 B.n1028 10.6151
R1782 B.n1028 B.n24 10.6151
R1783 B.n1022 B.n24 10.6151
R1784 B.n1022 B.n1021 10.6151
R1785 B.n1021 B.n1020 10.6151
R1786 B.n1020 B.n31 10.6151
R1787 B.n1014 B.n31 10.6151
R1788 B.n1014 B.n1013 10.6151
R1789 B.n1013 B.n1012 10.6151
R1790 B.n1012 B.n38 10.6151
R1791 B.n1006 B.n38 10.6151
R1792 B.n1006 B.n1005 10.6151
R1793 B.n1005 B.n1004 10.6151
R1794 B.n1004 B.n45 10.6151
R1795 B.n998 B.n45 10.6151
R1796 B.n998 B.n997 10.6151
R1797 B.n997 B.n996 10.6151
R1798 B.n996 B.n52 10.6151
R1799 B.n990 B.n52 10.6151
R1800 B.n990 B.n989 10.6151
R1801 B.n989 B.n988 10.6151
R1802 B.n988 B.n59 10.6151
R1803 B.n982 B.n59 10.6151
R1804 B.n982 B.n981 10.6151
R1805 B.n981 B.n980 10.6151
R1806 B.n980 B.n66 10.6151
R1807 B.n974 B.n66 10.6151
R1808 B.n974 B.n973 10.6151
R1809 B.n973 B.n972 10.6151
R1810 B.n972 B.n73 10.6151
R1811 B.n966 B.n73 10.6151
R1812 B.n966 B.n965 10.6151
R1813 B.n965 B.n964 10.6151
R1814 B.n964 B.n79 10.6151
R1815 B.n958 B.n79 10.6151
R1816 B.n958 B.n957 10.6151
R1817 B.n957 B.n956 10.6151
R1818 B.n956 B.n87 10.6151
R1819 B.n950 B.n87 10.6151
R1820 B.n950 B.n949 10.6151
R1821 B.n949 B.n948 10.6151
R1822 B.n948 B.n94 10.6151
R1823 B.n942 B.n94 10.6151
R1824 B.n942 B.n941 10.6151
R1825 B.n941 B.n940 10.6151
R1826 B.n940 B.n100 10.6151
R1827 B.n934 B.n100 10.6151
R1828 B.n934 B.n933 10.6151
R1829 B.n933 B.n932 10.6151
R1830 B.n932 B.n108 10.6151
R1831 B.n926 B.n108 10.6151
R1832 B.n926 B.n925 10.6151
R1833 B.n925 B.n924 10.6151
R1834 B.n924 B.n115 10.6151
R1835 B.n918 B.n115 10.6151
R1836 B.n918 B.n917 10.6151
R1837 B.n917 B.n916 10.6151
R1838 B.n916 B.n122 10.6151
R1839 B.n910 B.n122 10.6151
R1840 B.n910 B.n909 10.6151
R1841 B.n909 B.n908 10.6151
R1842 B.n908 B.n129 10.6151
R1843 B.n902 B.n129 10.6151
R1844 B.n902 B.n901 10.6151
R1845 B.n901 B.n900 10.6151
R1846 B.n900 B.n136 10.6151
R1847 B.n894 B.n136 10.6151
R1848 B.n894 B.n893 10.6151
R1849 B.n212 B.n174 6.5566
R1850 B.n229 B.n228 6.5566
R1851 B.n510 B.n509 6.5566
R1852 B.n493 B.n451 6.5566
R1853 B.n209 B.n174 4.05904
R1854 B.n230 B.n229 4.05904
R1855 B.n511 B.n510 4.05904
R1856 B.n490 B.n451 4.05904
R1857 B.n1052 B.n0 2.81026
R1858 B.n1052 B.n1 2.81026
R1859 B.n656 B.t0 1.1133
R1860 B.n81 B.t1 1.1133
R1861 VP.n33 VP.n32 161.3
R1862 VP.n34 VP.n29 161.3
R1863 VP.n36 VP.n35 161.3
R1864 VP.n37 VP.n28 161.3
R1865 VP.n39 VP.n38 161.3
R1866 VP.n40 VP.n27 161.3
R1867 VP.n42 VP.n41 161.3
R1868 VP.n43 VP.n26 161.3
R1869 VP.n45 VP.n44 161.3
R1870 VP.n46 VP.n25 161.3
R1871 VP.n48 VP.n47 161.3
R1872 VP.n49 VP.n24 161.3
R1873 VP.n51 VP.n50 161.3
R1874 VP.n52 VP.n23 161.3
R1875 VP.n54 VP.n53 161.3
R1876 VP.n55 VP.n22 161.3
R1877 VP.n58 VP.n57 161.3
R1878 VP.n59 VP.n21 161.3
R1879 VP.n61 VP.n60 161.3
R1880 VP.n62 VP.n20 161.3
R1881 VP.n64 VP.n63 161.3
R1882 VP.n65 VP.n19 161.3
R1883 VP.n67 VP.n66 161.3
R1884 VP.n68 VP.n18 161.3
R1885 VP.n70 VP.n69 161.3
R1886 VP.n125 VP.n124 161.3
R1887 VP.n123 VP.n1 161.3
R1888 VP.n122 VP.n121 161.3
R1889 VP.n120 VP.n2 161.3
R1890 VP.n119 VP.n118 161.3
R1891 VP.n117 VP.n3 161.3
R1892 VP.n116 VP.n115 161.3
R1893 VP.n114 VP.n4 161.3
R1894 VP.n113 VP.n112 161.3
R1895 VP.n110 VP.n5 161.3
R1896 VP.n109 VP.n108 161.3
R1897 VP.n107 VP.n6 161.3
R1898 VP.n106 VP.n105 161.3
R1899 VP.n104 VP.n7 161.3
R1900 VP.n103 VP.n102 161.3
R1901 VP.n101 VP.n8 161.3
R1902 VP.n100 VP.n99 161.3
R1903 VP.n98 VP.n9 161.3
R1904 VP.n97 VP.n96 161.3
R1905 VP.n95 VP.n10 161.3
R1906 VP.n94 VP.n93 161.3
R1907 VP.n92 VP.n11 161.3
R1908 VP.n91 VP.n90 161.3
R1909 VP.n89 VP.n12 161.3
R1910 VP.n88 VP.n87 161.3
R1911 VP.n85 VP.n13 161.3
R1912 VP.n84 VP.n83 161.3
R1913 VP.n82 VP.n14 161.3
R1914 VP.n81 VP.n80 161.3
R1915 VP.n79 VP.n15 161.3
R1916 VP.n78 VP.n77 161.3
R1917 VP.n76 VP.n16 161.3
R1918 VP.n75 VP.n74 161.3
R1919 VP.n73 VP.n72 88.1101
R1920 VP.n126 VP.n0 88.1101
R1921 VP.n71 VP.n17 88.1101
R1922 VP.n31 VP.n30 74.0089
R1923 VP.n30 VP.t0 61.7127
R1924 VP.n72 VP.n71 53.4539
R1925 VP.n80 VP.n79 43.4072
R1926 VP.n118 VP.n2 43.4072
R1927 VP.n63 VP.n19 43.4072
R1928 VP.n93 VP.n92 41.4647
R1929 VP.n105 VP.n6 41.4647
R1930 VP.n50 VP.n23 41.4647
R1931 VP.n38 VP.n37 41.4647
R1932 VP.n93 VP.n10 39.5221
R1933 VP.n105 VP.n104 39.5221
R1934 VP.n50 VP.n49 39.5221
R1935 VP.n38 VP.n27 39.5221
R1936 VP.n80 VP.n14 37.5796
R1937 VP.n118 VP.n117 37.5796
R1938 VP.n63 VP.n62 37.5796
R1939 VP.n99 VP.t9 30.1092
R1940 VP.n73 VP.t7 30.1092
R1941 VP.n86 VP.t8 30.1092
R1942 VP.n111 VP.t4 30.1092
R1943 VP.n0 VP.t1 30.1092
R1944 VP.n44 VP.t3 30.1092
R1945 VP.n17 VP.t6 30.1092
R1946 VP.n56 VP.t5 30.1092
R1947 VP.n31 VP.t2 30.1092
R1948 VP.n74 VP.n16 24.4675
R1949 VP.n78 VP.n16 24.4675
R1950 VP.n79 VP.n78 24.4675
R1951 VP.n84 VP.n14 24.4675
R1952 VP.n85 VP.n84 24.4675
R1953 VP.n87 VP.n12 24.4675
R1954 VP.n91 VP.n12 24.4675
R1955 VP.n92 VP.n91 24.4675
R1956 VP.n97 VP.n10 24.4675
R1957 VP.n98 VP.n97 24.4675
R1958 VP.n99 VP.n98 24.4675
R1959 VP.n99 VP.n8 24.4675
R1960 VP.n103 VP.n8 24.4675
R1961 VP.n104 VP.n103 24.4675
R1962 VP.n109 VP.n6 24.4675
R1963 VP.n110 VP.n109 24.4675
R1964 VP.n112 VP.n110 24.4675
R1965 VP.n116 VP.n4 24.4675
R1966 VP.n117 VP.n116 24.4675
R1967 VP.n122 VP.n2 24.4675
R1968 VP.n123 VP.n122 24.4675
R1969 VP.n124 VP.n123 24.4675
R1970 VP.n67 VP.n19 24.4675
R1971 VP.n68 VP.n67 24.4675
R1972 VP.n69 VP.n68 24.4675
R1973 VP.n54 VP.n23 24.4675
R1974 VP.n55 VP.n54 24.4675
R1975 VP.n57 VP.n55 24.4675
R1976 VP.n61 VP.n21 24.4675
R1977 VP.n62 VP.n61 24.4675
R1978 VP.n42 VP.n27 24.4675
R1979 VP.n43 VP.n42 24.4675
R1980 VP.n44 VP.n43 24.4675
R1981 VP.n44 VP.n25 24.4675
R1982 VP.n48 VP.n25 24.4675
R1983 VP.n49 VP.n48 24.4675
R1984 VP.n32 VP.n29 24.4675
R1985 VP.n36 VP.n29 24.4675
R1986 VP.n37 VP.n36 24.4675
R1987 VP.n86 VP.n85 23.4888
R1988 VP.n111 VP.n4 23.4888
R1989 VP.n56 VP.n21 23.4888
R1990 VP.n33 VP.n30 3.40896
R1991 VP.n74 VP.n73 1.95786
R1992 VP.n124 VP.n0 1.95786
R1993 VP.n69 VP.n17 1.95786
R1994 VP.n87 VP.n86 0.97918
R1995 VP.n112 VP.n111 0.97918
R1996 VP.n57 VP.n56 0.97918
R1997 VP.n32 VP.n31 0.97918
R1998 VP.n71 VP.n70 0.354971
R1999 VP.n75 VP.n72 0.354971
R2000 VP.n126 VP.n125 0.354971
R2001 VP VP.n126 0.26696
R2002 VP.n34 VP.n33 0.189894
R2003 VP.n35 VP.n34 0.189894
R2004 VP.n35 VP.n28 0.189894
R2005 VP.n39 VP.n28 0.189894
R2006 VP.n40 VP.n39 0.189894
R2007 VP.n41 VP.n40 0.189894
R2008 VP.n41 VP.n26 0.189894
R2009 VP.n45 VP.n26 0.189894
R2010 VP.n46 VP.n45 0.189894
R2011 VP.n47 VP.n46 0.189894
R2012 VP.n47 VP.n24 0.189894
R2013 VP.n51 VP.n24 0.189894
R2014 VP.n52 VP.n51 0.189894
R2015 VP.n53 VP.n52 0.189894
R2016 VP.n53 VP.n22 0.189894
R2017 VP.n58 VP.n22 0.189894
R2018 VP.n59 VP.n58 0.189894
R2019 VP.n60 VP.n59 0.189894
R2020 VP.n60 VP.n20 0.189894
R2021 VP.n64 VP.n20 0.189894
R2022 VP.n65 VP.n64 0.189894
R2023 VP.n66 VP.n65 0.189894
R2024 VP.n66 VP.n18 0.189894
R2025 VP.n70 VP.n18 0.189894
R2026 VP.n76 VP.n75 0.189894
R2027 VP.n77 VP.n76 0.189894
R2028 VP.n77 VP.n15 0.189894
R2029 VP.n81 VP.n15 0.189894
R2030 VP.n82 VP.n81 0.189894
R2031 VP.n83 VP.n82 0.189894
R2032 VP.n83 VP.n13 0.189894
R2033 VP.n88 VP.n13 0.189894
R2034 VP.n89 VP.n88 0.189894
R2035 VP.n90 VP.n89 0.189894
R2036 VP.n90 VP.n11 0.189894
R2037 VP.n94 VP.n11 0.189894
R2038 VP.n95 VP.n94 0.189894
R2039 VP.n96 VP.n95 0.189894
R2040 VP.n96 VP.n9 0.189894
R2041 VP.n100 VP.n9 0.189894
R2042 VP.n101 VP.n100 0.189894
R2043 VP.n102 VP.n101 0.189894
R2044 VP.n102 VP.n7 0.189894
R2045 VP.n106 VP.n7 0.189894
R2046 VP.n107 VP.n106 0.189894
R2047 VP.n108 VP.n107 0.189894
R2048 VP.n108 VP.n5 0.189894
R2049 VP.n113 VP.n5 0.189894
R2050 VP.n114 VP.n113 0.189894
R2051 VP.n115 VP.n114 0.189894
R2052 VP.n115 VP.n3 0.189894
R2053 VP.n119 VP.n3 0.189894
R2054 VP.n120 VP.n119 0.189894
R2055 VP.n121 VP.n120 0.189894
R2056 VP.n121 VP.n1 0.189894
R2057 VP.n125 VP.n1 0.189894
R2058 VTAIL.n104 VTAIL.n86 289.615
R2059 VTAIL.n20 VTAIL.n2 289.615
R2060 VTAIL.n80 VTAIL.n62 289.615
R2061 VTAIL.n52 VTAIL.n34 289.615
R2062 VTAIL.n95 VTAIL.n94 185
R2063 VTAIL.n97 VTAIL.n96 185
R2064 VTAIL.n90 VTAIL.n89 185
R2065 VTAIL.n103 VTAIL.n102 185
R2066 VTAIL.n105 VTAIL.n104 185
R2067 VTAIL.n11 VTAIL.n10 185
R2068 VTAIL.n13 VTAIL.n12 185
R2069 VTAIL.n6 VTAIL.n5 185
R2070 VTAIL.n19 VTAIL.n18 185
R2071 VTAIL.n21 VTAIL.n20 185
R2072 VTAIL.n81 VTAIL.n80 185
R2073 VTAIL.n79 VTAIL.n78 185
R2074 VTAIL.n66 VTAIL.n65 185
R2075 VTAIL.n73 VTAIL.n72 185
R2076 VTAIL.n71 VTAIL.n70 185
R2077 VTAIL.n53 VTAIL.n52 185
R2078 VTAIL.n51 VTAIL.n50 185
R2079 VTAIL.n38 VTAIL.n37 185
R2080 VTAIL.n45 VTAIL.n44 185
R2081 VTAIL.n43 VTAIL.n42 185
R2082 VTAIL.n93 VTAIL.t9 147.714
R2083 VTAIL.n9 VTAIL.t15 147.714
R2084 VTAIL.n69 VTAIL.t13 147.714
R2085 VTAIL.n41 VTAIL.t7 147.714
R2086 VTAIL.n96 VTAIL.n95 104.615
R2087 VTAIL.n96 VTAIL.n89 104.615
R2088 VTAIL.n103 VTAIL.n89 104.615
R2089 VTAIL.n104 VTAIL.n103 104.615
R2090 VTAIL.n12 VTAIL.n11 104.615
R2091 VTAIL.n12 VTAIL.n5 104.615
R2092 VTAIL.n19 VTAIL.n5 104.615
R2093 VTAIL.n20 VTAIL.n19 104.615
R2094 VTAIL.n80 VTAIL.n79 104.615
R2095 VTAIL.n79 VTAIL.n65 104.615
R2096 VTAIL.n72 VTAIL.n65 104.615
R2097 VTAIL.n72 VTAIL.n71 104.615
R2098 VTAIL.n52 VTAIL.n51 104.615
R2099 VTAIL.n51 VTAIL.n37 104.615
R2100 VTAIL.n44 VTAIL.n37 104.615
R2101 VTAIL.n44 VTAIL.n43 104.615
R2102 VTAIL.n61 VTAIL.n60 54.9327
R2103 VTAIL.n59 VTAIL.n58 54.9327
R2104 VTAIL.n33 VTAIL.n32 54.9327
R2105 VTAIL.n31 VTAIL.n30 54.9327
R2106 VTAIL.n111 VTAIL.n110 54.9326
R2107 VTAIL.n1 VTAIL.n0 54.9326
R2108 VTAIL.n27 VTAIL.n26 54.9326
R2109 VTAIL.n29 VTAIL.n28 54.9326
R2110 VTAIL.n95 VTAIL.t9 52.3082
R2111 VTAIL.n11 VTAIL.t15 52.3082
R2112 VTAIL.n71 VTAIL.t13 52.3082
R2113 VTAIL.n43 VTAIL.t7 52.3082
R2114 VTAIL.n109 VTAIL.n108 33.155
R2115 VTAIL.n25 VTAIL.n24 33.155
R2116 VTAIL.n85 VTAIL.n84 33.155
R2117 VTAIL.n57 VTAIL.n56 33.155
R2118 VTAIL.n31 VTAIL.n29 23.2721
R2119 VTAIL.n109 VTAIL.n85 19.8065
R2120 VTAIL.n94 VTAIL.n93 15.6631
R2121 VTAIL.n10 VTAIL.n9 15.6631
R2122 VTAIL.n70 VTAIL.n69 15.6631
R2123 VTAIL.n42 VTAIL.n41 15.6631
R2124 VTAIL.n97 VTAIL.n92 12.8005
R2125 VTAIL.n13 VTAIL.n8 12.8005
R2126 VTAIL.n73 VTAIL.n68 12.8005
R2127 VTAIL.n45 VTAIL.n40 12.8005
R2128 VTAIL.n98 VTAIL.n90 12.0247
R2129 VTAIL.n14 VTAIL.n6 12.0247
R2130 VTAIL.n74 VTAIL.n66 12.0247
R2131 VTAIL.n46 VTAIL.n38 12.0247
R2132 VTAIL.n102 VTAIL.n101 11.249
R2133 VTAIL.n18 VTAIL.n17 11.249
R2134 VTAIL.n78 VTAIL.n77 11.249
R2135 VTAIL.n50 VTAIL.n49 11.249
R2136 VTAIL.n105 VTAIL.n88 10.4732
R2137 VTAIL.n21 VTAIL.n4 10.4732
R2138 VTAIL.n81 VTAIL.n64 10.4732
R2139 VTAIL.n53 VTAIL.n36 10.4732
R2140 VTAIL.n106 VTAIL.n86 9.69747
R2141 VTAIL.n22 VTAIL.n2 9.69747
R2142 VTAIL.n82 VTAIL.n62 9.69747
R2143 VTAIL.n54 VTAIL.n34 9.69747
R2144 VTAIL.n108 VTAIL.n107 9.45567
R2145 VTAIL.n24 VTAIL.n23 9.45567
R2146 VTAIL.n84 VTAIL.n83 9.45567
R2147 VTAIL.n56 VTAIL.n55 9.45567
R2148 VTAIL.n107 VTAIL.n106 9.3005
R2149 VTAIL.n88 VTAIL.n87 9.3005
R2150 VTAIL.n101 VTAIL.n100 9.3005
R2151 VTAIL.n99 VTAIL.n98 9.3005
R2152 VTAIL.n92 VTAIL.n91 9.3005
R2153 VTAIL.n23 VTAIL.n22 9.3005
R2154 VTAIL.n4 VTAIL.n3 9.3005
R2155 VTAIL.n17 VTAIL.n16 9.3005
R2156 VTAIL.n15 VTAIL.n14 9.3005
R2157 VTAIL.n8 VTAIL.n7 9.3005
R2158 VTAIL.n83 VTAIL.n82 9.3005
R2159 VTAIL.n64 VTAIL.n63 9.3005
R2160 VTAIL.n77 VTAIL.n76 9.3005
R2161 VTAIL.n75 VTAIL.n74 9.3005
R2162 VTAIL.n68 VTAIL.n67 9.3005
R2163 VTAIL.n55 VTAIL.n54 9.3005
R2164 VTAIL.n36 VTAIL.n35 9.3005
R2165 VTAIL.n49 VTAIL.n48 9.3005
R2166 VTAIL.n47 VTAIL.n46 9.3005
R2167 VTAIL.n40 VTAIL.n39 9.3005
R2168 VTAIL.n93 VTAIL.n91 4.39059
R2169 VTAIL.n9 VTAIL.n7 4.39059
R2170 VTAIL.n69 VTAIL.n67 4.39059
R2171 VTAIL.n41 VTAIL.n39 4.39059
R2172 VTAIL.n110 VTAIL.t4 4.29551
R2173 VTAIL.n110 VTAIL.t8 4.29551
R2174 VTAIL.n0 VTAIL.t3 4.29551
R2175 VTAIL.n0 VTAIL.t2 4.29551
R2176 VTAIL.n26 VTAIL.t10 4.29551
R2177 VTAIL.n26 VTAIL.t11 4.29551
R2178 VTAIL.n28 VTAIL.t16 4.29551
R2179 VTAIL.n28 VTAIL.t19 4.29551
R2180 VTAIL.n60 VTAIL.t14 4.29551
R2181 VTAIL.n60 VTAIL.t12 4.29551
R2182 VTAIL.n58 VTAIL.t17 4.29551
R2183 VTAIL.n58 VTAIL.t18 4.29551
R2184 VTAIL.n32 VTAIL.t6 4.29551
R2185 VTAIL.n32 VTAIL.t1 4.29551
R2186 VTAIL.n30 VTAIL.t5 4.29551
R2187 VTAIL.n30 VTAIL.t0 4.29551
R2188 VTAIL.n108 VTAIL.n86 4.26717
R2189 VTAIL.n24 VTAIL.n2 4.26717
R2190 VTAIL.n84 VTAIL.n62 4.26717
R2191 VTAIL.n56 VTAIL.n34 4.26717
R2192 VTAIL.n106 VTAIL.n105 3.49141
R2193 VTAIL.n22 VTAIL.n21 3.49141
R2194 VTAIL.n82 VTAIL.n81 3.49141
R2195 VTAIL.n54 VTAIL.n53 3.49141
R2196 VTAIL.n33 VTAIL.n31 3.46602
R2197 VTAIL.n57 VTAIL.n33 3.46602
R2198 VTAIL.n61 VTAIL.n59 3.46602
R2199 VTAIL.n85 VTAIL.n61 3.46602
R2200 VTAIL.n29 VTAIL.n27 3.46602
R2201 VTAIL.n27 VTAIL.n25 3.46602
R2202 VTAIL.n111 VTAIL.n109 3.46602
R2203 VTAIL.n102 VTAIL.n88 2.71565
R2204 VTAIL.n18 VTAIL.n4 2.71565
R2205 VTAIL.n78 VTAIL.n64 2.71565
R2206 VTAIL.n50 VTAIL.n36 2.71565
R2207 VTAIL VTAIL.n1 2.65783
R2208 VTAIL.n59 VTAIL.n57 2.20309
R2209 VTAIL.n25 VTAIL.n1 2.20309
R2210 VTAIL.n101 VTAIL.n90 1.93989
R2211 VTAIL.n17 VTAIL.n6 1.93989
R2212 VTAIL.n77 VTAIL.n66 1.93989
R2213 VTAIL.n49 VTAIL.n38 1.93989
R2214 VTAIL.n98 VTAIL.n97 1.16414
R2215 VTAIL.n14 VTAIL.n13 1.16414
R2216 VTAIL.n74 VTAIL.n73 1.16414
R2217 VTAIL.n46 VTAIL.n45 1.16414
R2218 VTAIL VTAIL.n111 0.80869
R2219 VTAIL.n94 VTAIL.n92 0.388379
R2220 VTAIL.n10 VTAIL.n8 0.388379
R2221 VTAIL.n70 VTAIL.n68 0.388379
R2222 VTAIL.n42 VTAIL.n40 0.388379
R2223 VTAIL.n99 VTAIL.n91 0.155672
R2224 VTAIL.n100 VTAIL.n99 0.155672
R2225 VTAIL.n100 VTAIL.n87 0.155672
R2226 VTAIL.n107 VTAIL.n87 0.155672
R2227 VTAIL.n15 VTAIL.n7 0.155672
R2228 VTAIL.n16 VTAIL.n15 0.155672
R2229 VTAIL.n16 VTAIL.n3 0.155672
R2230 VTAIL.n23 VTAIL.n3 0.155672
R2231 VTAIL.n83 VTAIL.n63 0.155672
R2232 VTAIL.n76 VTAIL.n63 0.155672
R2233 VTAIL.n76 VTAIL.n75 0.155672
R2234 VTAIL.n75 VTAIL.n67 0.155672
R2235 VTAIL.n55 VTAIL.n35 0.155672
R2236 VTAIL.n48 VTAIL.n35 0.155672
R2237 VTAIL.n48 VTAIL.n47 0.155672
R2238 VTAIL.n47 VTAIL.n39 0.155672
R2239 VDD1.n18 VDD1.n0 289.615
R2240 VDD1.n43 VDD1.n25 289.615
R2241 VDD1.n19 VDD1.n18 185
R2242 VDD1.n17 VDD1.n16 185
R2243 VDD1.n4 VDD1.n3 185
R2244 VDD1.n11 VDD1.n10 185
R2245 VDD1.n9 VDD1.n8 185
R2246 VDD1.n34 VDD1.n33 185
R2247 VDD1.n36 VDD1.n35 185
R2248 VDD1.n29 VDD1.n28 185
R2249 VDD1.n42 VDD1.n41 185
R2250 VDD1.n44 VDD1.n43 185
R2251 VDD1.n7 VDD1.t9 147.714
R2252 VDD1.n32 VDD1.t2 147.714
R2253 VDD1.n18 VDD1.n17 104.615
R2254 VDD1.n17 VDD1.n3 104.615
R2255 VDD1.n10 VDD1.n3 104.615
R2256 VDD1.n10 VDD1.n9 104.615
R2257 VDD1.n35 VDD1.n34 104.615
R2258 VDD1.n35 VDD1.n28 104.615
R2259 VDD1.n42 VDD1.n28 104.615
R2260 VDD1.n43 VDD1.n42 104.615
R2261 VDD1.n51 VDD1.n50 74.1551
R2262 VDD1.n24 VDD1.n23 71.6115
R2263 VDD1.n53 VDD1.n52 71.6113
R2264 VDD1.n49 VDD1.n48 71.6113
R2265 VDD1.n24 VDD1.n22 53.2994
R2266 VDD1.n49 VDD1.n47 53.2994
R2267 VDD1.n9 VDD1.t9 52.3082
R2268 VDD1.n34 VDD1.t2 52.3082
R2269 VDD1.n53 VDD1.n51 46.4664
R2270 VDD1.n8 VDD1.n7 15.6631
R2271 VDD1.n33 VDD1.n32 15.6631
R2272 VDD1.n11 VDD1.n6 12.8005
R2273 VDD1.n36 VDD1.n31 12.8005
R2274 VDD1.n12 VDD1.n4 12.0247
R2275 VDD1.n37 VDD1.n29 12.0247
R2276 VDD1.n16 VDD1.n15 11.249
R2277 VDD1.n41 VDD1.n40 11.249
R2278 VDD1.n19 VDD1.n2 10.4732
R2279 VDD1.n44 VDD1.n27 10.4732
R2280 VDD1.n20 VDD1.n0 9.69747
R2281 VDD1.n45 VDD1.n25 9.69747
R2282 VDD1.n22 VDD1.n21 9.45567
R2283 VDD1.n47 VDD1.n46 9.45567
R2284 VDD1.n21 VDD1.n20 9.3005
R2285 VDD1.n2 VDD1.n1 9.3005
R2286 VDD1.n15 VDD1.n14 9.3005
R2287 VDD1.n13 VDD1.n12 9.3005
R2288 VDD1.n6 VDD1.n5 9.3005
R2289 VDD1.n46 VDD1.n45 9.3005
R2290 VDD1.n27 VDD1.n26 9.3005
R2291 VDD1.n40 VDD1.n39 9.3005
R2292 VDD1.n38 VDD1.n37 9.3005
R2293 VDD1.n31 VDD1.n30 9.3005
R2294 VDD1.n7 VDD1.n5 4.39059
R2295 VDD1.n32 VDD1.n30 4.39059
R2296 VDD1.n52 VDD1.t4 4.29551
R2297 VDD1.n52 VDD1.t3 4.29551
R2298 VDD1.n23 VDD1.t7 4.29551
R2299 VDD1.n23 VDD1.t6 4.29551
R2300 VDD1.n50 VDD1.t5 4.29551
R2301 VDD1.n50 VDD1.t8 4.29551
R2302 VDD1.n48 VDD1.t1 4.29551
R2303 VDD1.n48 VDD1.t0 4.29551
R2304 VDD1.n22 VDD1.n0 4.26717
R2305 VDD1.n47 VDD1.n25 4.26717
R2306 VDD1.n20 VDD1.n19 3.49141
R2307 VDD1.n45 VDD1.n44 3.49141
R2308 VDD1.n16 VDD1.n2 2.71565
R2309 VDD1.n41 VDD1.n27 2.71565
R2310 VDD1 VDD1.n53 2.54145
R2311 VDD1.n15 VDD1.n4 1.93989
R2312 VDD1.n40 VDD1.n29 1.93989
R2313 VDD1.n12 VDD1.n11 1.16414
R2314 VDD1.n37 VDD1.n36 1.16414
R2315 VDD1 VDD1.n24 0.925069
R2316 VDD1.n51 VDD1.n49 0.811533
R2317 VDD1.n8 VDD1.n6 0.388379
R2318 VDD1.n33 VDD1.n31 0.388379
R2319 VDD1.n21 VDD1.n1 0.155672
R2320 VDD1.n14 VDD1.n1 0.155672
R2321 VDD1.n14 VDD1.n13 0.155672
R2322 VDD1.n13 VDD1.n5 0.155672
R2323 VDD1.n38 VDD1.n30 0.155672
R2324 VDD1.n39 VDD1.n38 0.155672
R2325 VDD1.n39 VDD1.n26 0.155672
R2326 VDD1.n46 VDD1.n26 0.155672
R2327 VN.n108 VN.n107 161.3
R2328 VN.n106 VN.n56 161.3
R2329 VN.n105 VN.n104 161.3
R2330 VN.n103 VN.n57 161.3
R2331 VN.n102 VN.n101 161.3
R2332 VN.n100 VN.n58 161.3
R2333 VN.n99 VN.n98 161.3
R2334 VN.n97 VN.n59 161.3
R2335 VN.n96 VN.n95 161.3
R2336 VN.n94 VN.n60 161.3
R2337 VN.n93 VN.n92 161.3
R2338 VN.n91 VN.n62 161.3
R2339 VN.n90 VN.n89 161.3
R2340 VN.n88 VN.n63 161.3
R2341 VN.n87 VN.n86 161.3
R2342 VN.n85 VN.n64 161.3
R2343 VN.n84 VN.n83 161.3
R2344 VN.n82 VN.n65 161.3
R2345 VN.n81 VN.n80 161.3
R2346 VN.n79 VN.n66 161.3
R2347 VN.n78 VN.n77 161.3
R2348 VN.n76 VN.n67 161.3
R2349 VN.n75 VN.n74 161.3
R2350 VN.n73 VN.n68 161.3
R2351 VN.n72 VN.n71 161.3
R2352 VN.n53 VN.n52 161.3
R2353 VN.n51 VN.n1 161.3
R2354 VN.n50 VN.n49 161.3
R2355 VN.n48 VN.n2 161.3
R2356 VN.n47 VN.n46 161.3
R2357 VN.n45 VN.n3 161.3
R2358 VN.n44 VN.n43 161.3
R2359 VN.n42 VN.n4 161.3
R2360 VN.n41 VN.n40 161.3
R2361 VN.n38 VN.n5 161.3
R2362 VN.n37 VN.n36 161.3
R2363 VN.n35 VN.n6 161.3
R2364 VN.n34 VN.n33 161.3
R2365 VN.n32 VN.n7 161.3
R2366 VN.n31 VN.n30 161.3
R2367 VN.n29 VN.n8 161.3
R2368 VN.n28 VN.n27 161.3
R2369 VN.n26 VN.n9 161.3
R2370 VN.n25 VN.n24 161.3
R2371 VN.n23 VN.n10 161.3
R2372 VN.n22 VN.n21 161.3
R2373 VN.n20 VN.n11 161.3
R2374 VN.n19 VN.n18 161.3
R2375 VN.n17 VN.n12 161.3
R2376 VN.n16 VN.n15 161.3
R2377 VN.n54 VN.n0 88.1101
R2378 VN.n109 VN.n55 88.1101
R2379 VN.n14 VN.n13 74.0089
R2380 VN.n70 VN.n69 74.0089
R2381 VN.n69 VN.t7 61.7129
R2382 VN.n13 VN.t8 61.7129
R2383 VN VN.n109 53.6192
R2384 VN.n46 VN.n2 43.4072
R2385 VN.n101 VN.n57 43.4072
R2386 VN.n21 VN.n20 41.4647
R2387 VN.n33 VN.n6 41.4647
R2388 VN.n77 VN.n76 41.4647
R2389 VN.n89 VN.n62 41.4647
R2390 VN.n21 VN.n10 39.5221
R2391 VN.n33 VN.n32 39.5221
R2392 VN.n77 VN.n66 39.5221
R2393 VN.n89 VN.n88 39.5221
R2394 VN.n46 VN.n45 37.5796
R2395 VN.n101 VN.n100 37.5796
R2396 VN.n27 VN.t5 30.1092
R2397 VN.n14 VN.t6 30.1092
R2398 VN.n39 VN.t1 30.1092
R2399 VN.n0 VN.t0 30.1092
R2400 VN.n83 VN.t2 30.1092
R2401 VN.n70 VN.t9 30.1092
R2402 VN.n61 VN.t3 30.1092
R2403 VN.n55 VN.t4 30.1092
R2404 VN.n15 VN.n12 24.4675
R2405 VN.n19 VN.n12 24.4675
R2406 VN.n20 VN.n19 24.4675
R2407 VN.n25 VN.n10 24.4675
R2408 VN.n26 VN.n25 24.4675
R2409 VN.n27 VN.n26 24.4675
R2410 VN.n27 VN.n8 24.4675
R2411 VN.n31 VN.n8 24.4675
R2412 VN.n32 VN.n31 24.4675
R2413 VN.n37 VN.n6 24.4675
R2414 VN.n38 VN.n37 24.4675
R2415 VN.n40 VN.n38 24.4675
R2416 VN.n44 VN.n4 24.4675
R2417 VN.n45 VN.n44 24.4675
R2418 VN.n50 VN.n2 24.4675
R2419 VN.n51 VN.n50 24.4675
R2420 VN.n52 VN.n51 24.4675
R2421 VN.n76 VN.n75 24.4675
R2422 VN.n75 VN.n68 24.4675
R2423 VN.n71 VN.n68 24.4675
R2424 VN.n88 VN.n87 24.4675
R2425 VN.n87 VN.n64 24.4675
R2426 VN.n83 VN.n64 24.4675
R2427 VN.n83 VN.n82 24.4675
R2428 VN.n82 VN.n81 24.4675
R2429 VN.n81 VN.n66 24.4675
R2430 VN.n100 VN.n99 24.4675
R2431 VN.n99 VN.n59 24.4675
R2432 VN.n95 VN.n94 24.4675
R2433 VN.n94 VN.n93 24.4675
R2434 VN.n93 VN.n62 24.4675
R2435 VN.n107 VN.n106 24.4675
R2436 VN.n106 VN.n105 24.4675
R2437 VN.n105 VN.n57 24.4675
R2438 VN.n39 VN.n4 23.4888
R2439 VN.n61 VN.n59 23.4888
R2440 VN.n72 VN.n69 3.40897
R2441 VN.n16 VN.n13 3.40897
R2442 VN.n52 VN.n0 1.95786
R2443 VN.n107 VN.n55 1.95786
R2444 VN.n15 VN.n14 0.97918
R2445 VN.n40 VN.n39 0.97918
R2446 VN.n71 VN.n70 0.97918
R2447 VN.n95 VN.n61 0.97918
R2448 VN.n109 VN.n108 0.354971
R2449 VN.n54 VN.n53 0.354971
R2450 VN VN.n54 0.26696
R2451 VN.n108 VN.n56 0.189894
R2452 VN.n104 VN.n56 0.189894
R2453 VN.n104 VN.n103 0.189894
R2454 VN.n103 VN.n102 0.189894
R2455 VN.n102 VN.n58 0.189894
R2456 VN.n98 VN.n58 0.189894
R2457 VN.n98 VN.n97 0.189894
R2458 VN.n97 VN.n96 0.189894
R2459 VN.n96 VN.n60 0.189894
R2460 VN.n92 VN.n60 0.189894
R2461 VN.n92 VN.n91 0.189894
R2462 VN.n91 VN.n90 0.189894
R2463 VN.n90 VN.n63 0.189894
R2464 VN.n86 VN.n63 0.189894
R2465 VN.n86 VN.n85 0.189894
R2466 VN.n85 VN.n84 0.189894
R2467 VN.n84 VN.n65 0.189894
R2468 VN.n80 VN.n65 0.189894
R2469 VN.n80 VN.n79 0.189894
R2470 VN.n79 VN.n78 0.189894
R2471 VN.n78 VN.n67 0.189894
R2472 VN.n74 VN.n67 0.189894
R2473 VN.n74 VN.n73 0.189894
R2474 VN.n73 VN.n72 0.189894
R2475 VN.n17 VN.n16 0.189894
R2476 VN.n18 VN.n17 0.189894
R2477 VN.n18 VN.n11 0.189894
R2478 VN.n22 VN.n11 0.189894
R2479 VN.n23 VN.n22 0.189894
R2480 VN.n24 VN.n23 0.189894
R2481 VN.n24 VN.n9 0.189894
R2482 VN.n28 VN.n9 0.189894
R2483 VN.n29 VN.n28 0.189894
R2484 VN.n30 VN.n29 0.189894
R2485 VN.n30 VN.n7 0.189894
R2486 VN.n34 VN.n7 0.189894
R2487 VN.n35 VN.n34 0.189894
R2488 VN.n36 VN.n35 0.189894
R2489 VN.n36 VN.n5 0.189894
R2490 VN.n41 VN.n5 0.189894
R2491 VN.n42 VN.n41 0.189894
R2492 VN.n43 VN.n42 0.189894
R2493 VN.n43 VN.n3 0.189894
R2494 VN.n47 VN.n3 0.189894
R2495 VN.n48 VN.n47 0.189894
R2496 VN.n49 VN.n48 0.189894
R2497 VN.n49 VN.n1 0.189894
R2498 VN.n53 VN.n1 0.189894
R2499 VDD2.n45 VDD2.n27 289.615
R2500 VDD2.n18 VDD2.n0 289.615
R2501 VDD2.n46 VDD2.n45 185
R2502 VDD2.n44 VDD2.n43 185
R2503 VDD2.n31 VDD2.n30 185
R2504 VDD2.n38 VDD2.n37 185
R2505 VDD2.n36 VDD2.n35 185
R2506 VDD2.n9 VDD2.n8 185
R2507 VDD2.n11 VDD2.n10 185
R2508 VDD2.n4 VDD2.n3 185
R2509 VDD2.n17 VDD2.n16 185
R2510 VDD2.n19 VDD2.n18 185
R2511 VDD2.n34 VDD2.t5 147.714
R2512 VDD2.n7 VDD2.t1 147.714
R2513 VDD2.n45 VDD2.n44 104.615
R2514 VDD2.n44 VDD2.n30 104.615
R2515 VDD2.n37 VDD2.n30 104.615
R2516 VDD2.n37 VDD2.n36 104.615
R2517 VDD2.n10 VDD2.n9 104.615
R2518 VDD2.n10 VDD2.n3 104.615
R2519 VDD2.n17 VDD2.n3 104.615
R2520 VDD2.n18 VDD2.n17 104.615
R2521 VDD2.n26 VDD2.n25 74.1551
R2522 VDD2 VDD2.n53 74.1523
R2523 VDD2.n52 VDD2.n51 71.6115
R2524 VDD2.n24 VDD2.n23 71.6113
R2525 VDD2.n24 VDD2.n22 53.2994
R2526 VDD2.n36 VDD2.t5 52.3082
R2527 VDD2.n9 VDD2.t1 52.3082
R2528 VDD2.n50 VDD2.n49 49.8338
R2529 VDD2.n50 VDD2.n26 44.1506
R2530 VDD2.n35 VDD2.n34 15.6631
R2531 VDD2.n8 VDD2.n7 15.6631
R2532 VDD2.n38 VDD2.n33 12.8005
R2533 VDD2.n11 VDD2.n6 12.8005
R2534 VDD2.n39 VDD2.n31 12.0247
R2535 VDD2.n12 VDD2.n4 12.0247
R2536 VDD2.n43 VDD2.n42 11.249
R2537 VDD2.n16 VDD2.n15 11.249
R2538 VDD2.n46 VDD2.n29 10.4732
R2539 VDD2.n19 VDD2.n2 10.4732
R2540 VDD2.n47 VDD2.n27 9.69747
R2541 VDD2.n20 VDD2.n0 9.69747
R2542 VDD2.n49 VDD2.n48 9.45567
R2543 VDD2.n22 VDD2.n21 9.45567
R2544 VDD2.n48 VDD2.n47 9.3005
R2545 VDD2.n29 VDD2.n28 9.3005
R2546 VDD2.n42 VDD2.n41 9.3005
R2547 VDD2.n40 VDD2.n39 9.3005
R2548 VDD2.n33 VDD2.n32 9.3005
R2549 VDD2.n21 VDD2.n20 9.3005
R2550 VDD2.n2 VDD2.n1 9.3005
R2551 VDD2.n15 VDD2.n14 9.3005
R2552 VDD2.n13 VDD2.n12 9.3005
R2553 VDD2.n6 VDD2.n5 9.3005
R2554 VDD2.n34 VDD2.n32 4.39059
R2555 VDD2.n7 VDD2.n5 4.39059
R2556 VDD2.n53 VDD2.t0 4.29551
R2557 VDD2.n53 VDD2.t2 4.29551
R2558 VDD2.n51 VDD2.t6 4.29551
R2559 VDD2.n51 VDD2.t7 4.29551
R2560 VDD2.n25 VDD2.t8 4.29551
R2561 VDD2.n25 VDD2.t9 4.29551
R2562 VDD2.n23 VDD2.t3 4.29551
R2563 VDD2.n23 VDD2.t4 4.29551
R2564 VDD2.n49 VDD2.n27 4.26717
R2565 VDD2.n22 VDD2.n0 4.26717
R2566 VDD2.n47 VDD2.n46 3.49141
R2567 VDD2.n20 VDD2.n19 3.49141
R2568 VDD2.n52 VDD2.n50 3.46602
R2569 VDD2.n43 VDD2.n29 2.71565
R2570 VDD2.n16 VDD2.n2 2.71565
R2571 VDD2.n42 VDD2.n31 1.93989
R2572 VDD2.n15 VDD2.n4 1.93989
R2573 VDD2.n39 VDD2.n38 1.16414
R2574 VDD2.n12 VDD2.n11 1.16414
R2575 VDD2 VDD2.n52 0.925069
R2576 VDD2.n26 VDD2.n24 0.811533
R2577 VDD2.n35 VDD2.n33 0.388379
R2578 VDD2.n8 VDD2.n6 0.388379
R2579 VDD2.n48 VDD2.n28 0.155672
R2580 VDD2.n41 VDD2.n28 0.155672
R2581 VDD2.n41 VDD2.n40 0.155672
R2582 VDD2.n40 VDD2.n32 0.155672
R2583 VDD2.n13 VDD2.n5 0.155672
R2584 VDD2.n14 VDD2.n13 0.155672
R2585 VDD2.n14 VDD2.n1 0.155672
R2586 VDD2.n21 VDD2.n1 0.155672
C0 VP VTAIL 6.4817f
C1 VDD1 VDD2 2.88147f
C2 VN VDD1 0.159493f
C3 VN VDD2 4.70036f
C4 VTAIL VDD1 8.033319f
C5 VTAIL VDD2 8.093659f
C6 VN VTAIL 6.46744f
C7 VP VDD1 5.26351f
C8 VP VDD2 0.726435f
C9 VP VN 8.645519f
C10 VDD2 B 7.26434f
C11 VDD1 B 7.162355f
C12 VTAIL B 5.410303f
C13 VN B 22.613949f
C14 VP B 21.102837f
C15 VDD2.n0 B 0.03853f
C16 VDD2.n1 B 0.027812f
C17 VDD2.n2 B 0.014945f
C18 VDD2.n3 B 0.035325f
C19 VDD2.n4 B 0.015824f
C20 VDD2.n5 B 0.483113f
C21 VDD2.n6 B 0.014945f
C22 VDD2.t1 B 0.057967f
C23 VDD2.n7 B 0.110293f
C24 VDD2.n8 B 0.020847f
C25 VDD2.n9 B 0.026493f
C26 VDD2.n10 B 0.035325f
C27 VDD2.n11 B 0.015824f
C28 VDD2.n12 B 0.014945f
C29 VDD2.n13 B 0.027812f
C30 VDD2.n14 B 0.027812f
C31 VDD2.n15 B 0.014945f
C32 VDD2.n16 B 0.015824f
C33 VDD2.n17 B 0.035325f
C34 VDD2.n18 B 0.075476f
C35 VDD2.n19 B 0.015824f
C36 VDD2.n20 B 0.014945f
C37 VDD2.n21 B 0.066186f
C38 VDD2.n22 B 0.085122f
C39 VDD2.t3 B 0.101318f
C40 VDD2.t4 B 0.101318f
C41 VDD2.n23 B 0.815208f
C42 VDD2.n24 B 0.945132f
C43 VDD2.t8 B 0.101318f
C44 VDD2.t9 B 0.101318f
C45 VDD2.n25 B 0.841609f
C46 VDD2.n26 B 3.35325f
C47 VDD2.n27 B 0.03853f
C48 VDD2.n28 B 0.027812f
C49 VDD2.n29 B 0.014945f
C50 VDD2.n30 B 0.035325f
C51 VDD2.n31 B 0.015824f
C52 VDD2.n32 B 0.483113f
C53 VDD2.n33 B 0.014945f
C54 VDD2.t5 B 0.057967f
C55 VDD2.n34 B 0.110293f
C56 VDD2.n35 B 0.020847f
C57 VDD2.n36 B 0.026493f
C58 VDD2.n37 B 0.035325f
C59 VDD2.n38 B 0.015824f
C60 VDD2.n39 B 0.014945f
C61 VDD2.n40 B 0.027812f
C62 VDD2.n41 B 0.027812f
C63 VDD2.n42 B 0.014945f
C64 VDD2.n43 B 0.015824f
C65 VDD2.n44 B 0.035325f
C66 VDD2.n45 B 0.075476f
C67 VDD2.n46 B 0.015824f
C68 VDD2.n47 B 0.014945f
C69 VDD2.n48 B 0.066186f
C70 VDD2.n49 B 0.061376f
C71 VDD2.n50 B 3.05194f
C72 VDD2.t6 B 0.101318f
C73 VDD2.t7 B 0.101318f
C74 VDD2.n51 B 0.815212f
C75 VDD2.n52 B 0.613043f
C76 VDD2.t0 B 0.101318f
C77 VDD2.t2 B 0.101318f
C78 VDD2.n53 B 0.841563f
C79 VN.t0 B 0.932457f
C80 VN.n0 B 0.430408f
C81 VN.n1 B 0.021084f
C82 VN.n2 B 0.041156f
C83 VN.n3 B 0.021084f
C84 VN.n4 B 0.03852f
C85 VN.n5 B 0.021084f
C86 VN.n6 B 0.04168f
C87 VN.n7 B 0.021084f
C88 VN.n8 B 0.039296f
C89 VN.n9 B 0.021084f
C90 VN.t5 B 0.932457f
C91 VN.n10 B 0.042102f
C92 VN.n11 B 0.021084f
C93 VN.n12 B 0.039296f
C94 VN.t8 B 1.19591f
C95 VN.n13 B 0.418355f
C96 VN.t6 B 0.932457f
C97 VN.n14 B 0.421249f
C98 VN.n15 B 0.020671f
C99 VN.n16 B 0.267876f
C100 VN.n17 B 0.021084f
C101 VN.n18 B 0.021084f
C102 VN.n19 B 0.039296f
C103 VN.n20 B 0.04168f
C104 VN.n21 B 0.017072f
C105 VN.n22 B 0.021084f
C106 VN.n23 B 0.021084f
C107 VN.n24 B 0.021084f
C108 VN.n25 B 0.039296f
C109 VN.n26 B 0.039296f
C110 VN.n27 B 0.374341f
C111 VN.n28 B 0.021084f
C112 VN.n29 B 0.021084f
C113 VN.n30 B 0.021084f
C114 VN.n31 B 0.039296f
C115 VN.n32 B 0.042102f
C116 VN.n33 B 0.017072f
C117 VN.n34 B 0.021084f
C118 VN.n35 B 0.021084f
C119 VN.n36 B 0.021084f
C120 VN.n37 B 0.039296f
C121 VN.n38 B 0.039296f
C122 VN.t1 B 0.932457f
C123 VN.n39 B 0.354446f
C124 VN.n40 B 0.020671f
C125 VN.n41 B 0.021084f
C126 VN.n42 B 0.021084f
C127 VN.n43 B 0.021084f
C128 VN.n44 B 0.039296f
C129 VN.n45 B 0.042408f
C130 VN.n46 B 0.01729f
C131 VN.n47 B 0.021084f
C132 VN.n48 B 0.021084f
C133 VN.n49 B 0.021084f
C134 VN.n50 B 0.039296f
C135 VN.n51 B 0.039296f
C136 VN.n52 B 0.021447f
C137 VN.n53 B 0.034029f
C138 VN.n54 B 0.064024f
C139 VN.t4 B 0.932457f
C140 VN.n55 B 0.430408f
C141 VN.n56 B 0.021084f
C142 VN.n57 B 0.041156f
C143 VN.n58 B 0.021084f
C144 VN.n59 B 0.03852f
C145 VN.n60 B 0.021084f
C146 VN.t3 B 0.932457f
C147 VN.n61 B 0.354446f
C148 VN.n62 B 0.04168f
C149 VN.n63 B 0.021084f
C150 VN.n64 B 0.039296f
C151 VN.n65 B 0.021084f
C152 VN.t2 B 0.932457f
C153 VN.n66 B 0.042102f
C154 VN.n67 B 0.021084f
C155 VN.n68 B 0.039296f
C156 VN.t7 B 1.19591f
C157 VN.n69 B 0.418355f
C158 VN.t9 B 0.932457f
C159 VN.n70 B 0.421249f
C160 VN.n71 B 0.020671f
C161 VN.n72 B 0.267876f
C162 VN.n73 B 0.021084f
C163 VN.n74 B 0.021084f
C164 VN.n75 B 0.039296f
C165 VN.n76 B 0.04168f
C166 VN.n77 B 0.017072f
C167 VN.n78 B 0.021084f
C168 VN.n79 B 0.021084f
C169 VN.n80 B 0.021084f
C170 VN.n81 B 0.039296f
C171 VN.n82 B 0.039296f
C172 VN.n83 B 0.374341f
C173 VN.n84 B 0.021084f
C174 VN.n85 B 0.021084f
C175 VN.n86 B 0.021084f
C176 VN.n87 B 0.039296f
C177 VN.n88 B 0.042102f
C178 VN.n89 B 0.017072f
C179 VN.n90 B 0.021084f
C180 VN.n91 B 0.021084f
C181 VN.n92 B 0.021084f
C182 VN.n93 B 0.039296f
C183 VN.n94 B 0.039296f
C184 VN.n95 B 0.020671f
C185 VN.n96 B 0.021084f
C186 VN.n97 B 0.021084f
C187 VN.n98 B 0.021084f
C188 VN.n99 B 0.039296f
C189 VN.n100 B 0.042408f
C190 VN.n101 B 0.01729f
C191 VN.n102 B 0.021084f
C192 VN.n103 B 0.021084f
C193 VN.n104 B 0.021084f
C194 VN.n105 B 0.039296f
C195 VN.n106 B 0.039296f
C196 VN.n107 B 0.021447f
C197 VN.n108 B 0.034029f
C198 VN.n109 B 1.33903f
C199 VDD1.n0 B 0.039498f
C200 VDD1.n1 B 0.028511f
C201 VDD1.n2 B 0.015321f
C202 VDD1.n3 B 0.036213f
C203 VDD1.n4 B 0.016222f
C204 VDD1.n5 B 0.495258f
C205 VDD1.n6 B 0.015321f
C206 VDD1.t9 B 0.059424f
C207 VDD1.n7 B 0.113065f
C208 VDD1.n8 B 0.021371f
C209 VDD1.n9 B 0.027159f
C210 VDD1.n10 B 0.036213f
C211 VDD1.n11 B 0.016222f
C212 VDD1.n12 B 0.015321f
C213 VDD1.n13 B 0.028511f
C214 VDD1.n14 B 0.028511f
C215 VDD1.n15 B 0.015321f
C216 VDD1.n16 B 0.016222f
C217 VDD1.n17 B 0.036213f
C218 VDD1.n18 B 0.077374f
C219 VDD1.n19 B 0.016222f
C220 VDD1.n20 B 0.015321f
C221 VDD1.n21 B 0.06785f
C222 VDD1.n22 B 0.087262f
C223 VDD1.t7 B 0.103866f
C224 VDD1.t6 B 0.103866f
C225 VDD1.n23 B 0.835706f
C226 VDD1.n24 B 0.978504f
C227 VDD1.n25 B 0.039498f
C228 VDD1.n26 B 0.028511f
C229 VDD1.n27 B 0.015321f
C230 VDD1.n28 B 0.036213f
C231 VDD1.n29 B 0.016222f
C232 VDD1.n30 B 0.495258f
C233 VDD1.n31 B 0.015321f
C234 VDD1.t2 B 0.059424f
C235 VDD1.n32 B 0.113065f
C236 VDD1.n33 B 0.021371f
C237 VDD1.n34 B 0.027159f
C238 VDD1.n35 B 0.036213f
C239 VDD1.n36 B 0.016222f
C240 VDD1.n37 B 0.015321f
C241 VDD1.n38 B 0.028511f
C242 VDD1.n39 B 0.028511f
C243 VDD1.n40 B 0.015321f
C244 VDD1.n41 B 0.016222f
C245 VDD1.n42 B 0.036213f
C246 VDD1.n43 B 0.077374f
C247 VDD1.n44 B 0.016222f
C248 VDD1.n45 B 0.015321f
C249 VDD1.n46 B 0.06785f
C250 VDD1.n47 B 0.087262f
C251 VDD1.t1 B 0.103866f
C252 VDD1.t0 B 0.103866f
C253 VDD1.n48 B 0.835702f
C254 VDD1.n49 B 0.968892f
C255 VDD1.t5 B 0.103866f
C256 VDD1.t8 B 0.103866f
C257 VDD1.n50 B 0.862767f
C258 VDD1.n51 B 3.60636f
C259 VDD1.t4 B 0.103866f
C260 VDD1.t3 B 0.103866f
C261 VDD1.n52 B 0.835702f
C262 VDD1.n53 B 3.47921f
C263 VTAIL.t3 B 0.116774f
C264 VTAIL.t2 B 0.116774f
C265 VTAIL.n0 B 0.864559f
C266 VTAIL.n1 B 0.786522f
C267 VTAIL.n2 B 0.044407f
C268 VTAIL.n3 B 0.032055f
C269 VTAIL.n4 B 0.017225f
C270 VTAIL.n5 B 0.040713f
C271 VTAIL.n6 B 0.018238f
C272 VTAIL.n7 B 0.556808f
C273 VTAIL.n8 B 0.017225f
C274 VTAIL.t15 B 0.06681f
C275 VTAIL.n9 B 0.127117f
C276 VTAIL.n10 B 0.024027f
C277 VTAIL.n11 B 0.030535f
C278 VTAIL.n12 B 0.040713f
C279 VTAIL.n13 B 0.018238f
C280 VTAIL.n14 B 0.017225f
C281 VTAIL.n15 B 0.032055f
C282 VTAIL.n16 B 0.032055f
C283 VTAIL.n17 B 0.017225f
C284 VTAIL.n18 B 0.018238f
C285 VTAIL.n19 B 0.040713f
C286 VTAIL.n20 B 0.086989f
C287 VTAIL.n21 B 0.018238f
C288 VTAIL.n22 B 0.017225f
C289 VTAIL.n23 B 0.076282f
C290 VTAIL.n24 B 0.048623f
C291 VTAIL.n25 B 0.614055f
C292 VTAIL.t10 B 0.116774f
C293 VTAIL.t11 B 0.116774f
C294 VTAIL.n26 B 0.864559f
C295 VTAIL.n27 B 1.00044f
C296 VTAIL.t16 B 0.116774f
C297 VTAIL.t19 B 0.116774f
C298 VTAIL.n28 B 0.864559f
C299 VTAIL.n29 B 2.20429f
C300 VTAIL.t5 B 0.116774f
C301 VTAIL.t0 B 0.116774f
C302 VTAIL.n30 B 0.864565f
C303 VTAIL.n31 B 2.20428f
C304 VTAIL.t6 B 0.116774f
C305 VTAIL.t1 B 0.116774f
C306 VTAIL.n32 B 0.864565f
C307 VTAIL.n33 B 1.00044f
C308 VTAIL.n34 B 0.044407f
C309 VTAIL.n35 B 0.032055f
C310 VTAIL.n36 B 0.017225f
C311 VTAIL.n37 B 0.040713f
C312 VTAIL.n38 B 0.018238f
C313 VTAIL.n39 B 0.556807f
C314 VTAIL.n40 B 0.017225f
C315 VTAIL.t7 B 0.06681f
C316 VTAIL.n41 B 0.127117f
C317 VTAIL.n42 B 0.024027f
C318 VTAIL.n43 B 0.030535f
C319 VTAIL.n44 B 0.040713f
C320 VTAIL.n45 B 0.018238f
C321 VTAIL.n46 B 0.017225f
C322 VTAIL.n47 B 0.032055f
C323 VTAIL.n48 B 0.032055f
C324 VTAIL.n49 B 0.017225f
C325 VTAIL.n50 B 0.018238f
C326 VTAIL.n51 B 0.040713f
C327 VTAIL.n52 B 0.086989f
C328 VTAIL.n53 B 0.018238f
C329 VTAIL.n54 B 0.017225f
C330 VTAIL.n55 B 0.076282f
C331 VTAIL.n56 B 0.048623f
C332 VTAIL.n57 B 0.614055f
C333 VTAIL.t17 B 0.116774f
C334 VTAIL.t18 B 0.116774f
C335 VTAIL.n58 B 0.864565f
C336 VTAIL.n59 B 0.869992f
C337 VTAIL.t14 B 0.116774f
C338 VTAIL.t12 B 0.116774f
C339 VTAIL.n60 B 0.864565f
C340 VTAIL.n61 B 1.00044f
C341 VTAIL.n62 B 0.044407f
C342 VTAIL.n63 B 0.032055f
C343 VTAIL.n64 B 0.017225f
C344 VTAIL.n65 B 0.040713f
C345 VTAIL.n66 B 0.018238f
C346 VTAIL.n67 B 0.556807f
C347 VTAIL.n68 B 0.017225f
C348 VTAIL.t13 B 0.06681f
C349 VTAIL.n69 B 0.127117f
C350 VTAIL.n70 B 0.024027f
C351 VTAIL.n71 B 0.030535f
C352 VTAIL.n72 B 0.040713f
C353 VTAIL.n73 B 0.018238f
C354 VTAIL.n74 B 0.017225f
C355 VTAIL.n75 B 0.032055f
C356 VTAIL.n76 B 0.032055f
C357 VTAIL.n77 B 0.017225f
C358 VTAIL.n78 B 0.018238f
C359 VTAIL.n79 B 0.040713f
C360 VTAIL.n80 B 0.086989f
C361 VTAIL.n81 B 0.018238f
C362 VTAIL.n82 B 0.017225f
C363 VTAIL.n83 B 0.076282f
C364 VTAIL.n84 B 0.048623f
C365 VTAIL.n85 B 1.5904f
C366 VTAIL.n86 B 0.044407f
C367 VTAIL.n87 B 0.032055f
C368 VTAIL.n88 B 0.017225f
C369 VTAIL.n89 B 0.040713f
C370 VTAIL.n90 B 0.018238f
C371 VTAIL.n91 B 0.556808f
C372 VTAIL.n92 B 0.017225f
C373 VTAIL.t9 B 0.06681f
C374 VTAIL.n93 B 0.127117f
C375 VTAIL.n94 B 0.024027f
C376 VTAIL.n95 B 0.030535f
C377 VTAIL.n96 B 0.040713f
C378 VTAIL.n97 B 0.018238f
C379 VTAIL.n98 B 0.017225f
C380 VTAIL.n99 B 0.032055f
C381 VTAIL.n100 B 0.032055f
C382 VTAIL.n101 B 0.017225f
C383 VTAIL.n102 B 0.018238f
C384 VTAIL.n103 B 0.040713f
C385 VTAIL.n104 B 0.086989f
C386 VTAIL.n105 B 0.018238f
C387 VTAIL.n106 B 0.017225f
C388 VTAIL.n107 B 0.076282f
C389 VTAIL.n108 B 0.048623f
C390 VTAIL.n109 B 1.5904f
C391 VTAIL.t4 B 0.116774f
C392 VTAIL.t8 B 0.116774f
C393 VTAIL.n110 B 0.864559f
C394 VTAIL.n111 B 0.725974f
C395 VP.t1 B 0.962154f
C396 VP.n0 B 0.444116f
C397 VP.n1 B 0.021756f
C398 VP.n2 B 0.042467f
C399 VP.n3 B 0.021756f
C400 VP.n4 B 0.039746f
C401 VP.n5 B 0.021756f
C402 VP.n6 B 0.043007f
C403 VP.n7 B 0.021756f
C404 VP.n8 B 0.040547f
C405 VP.n9 B 0.021756f
C406 VP.t9 B 0.962154f
C407 VP.n10 B 0.043443f
C408 VP.n11 B 0.021756f
C409 VP.n12 B 0.040547f
C410 VP.n13 B 0.021756f
C411 VP.t8 B 0.962154f
C412 VP.n14 B 0.043759f
C413 VP.n15 B 0.021756f
C414 VP.n16 B 0.040547f
C415 VP.t6 B 0.962154f
C416 VP.n17 B 0.444116f
C417 VP.n18 B 0.021756f
C418 VP.n19 B 0.042467f
C419 VP.n20 B 0.021756f
C420 VP.n21 B 0.039746f
C421 VP.n22 B 0.021756f
C422 VP.n23 B 0.043007f
C423 VP.n24 B 0.021756f
C424 VP.n25 B 0.040547f
C425 VP.n26 B 0.021756f
C426 VP.t3 B 0.962154f
C427 VP.n27 B 0.043443f
C428 VP.n28 B 0.021756f
C429 VP.n29 B 0.040547f
C430 VP.t0 B 1.23399f
C431 VP.n30 B 0.431679f
C432 VP.t2 B 0.962154f
C433 VP.n31 B 0.434665f
C434 VP.n32 B 0.021329f
C435 VP.n33 B 0.276408f
C436 VP.n34 B 0.021756f
C437 VP.n35 B 0.021756f
C438 VP.n36 B 0.040547f
C439 VP.n37 B 0.043007f
C440 VP.n38 B 0.017615f
C441 VP.n39 B 0.021756f
C442 VP.n40 B 0.021756f
C443 VP.n41 B 0.021756f
C444 VP.n42 B 0.040547f
C445 VP.n43 B 0.040547f
C446 VP.n44 B 0.386263f
C447 VP.n45 B 0.021756f
C448 VP.n46 B 0.021756f
C449 VP.n47 B 0.021756f
C450 VP.n48 B 0.040547f
C451 VP.n49 B 0.043443f
C452 VP.n50 B 0.017615f
C453 VP.n51 B 0.021756f
C454 VP.n52 B 0.021756f
C455 VP.n53 B 0.021756f
C456 VP.n54 B 0.040547f
C457 VP.n55 B 0.040547f
C458 VP.t5 B 0.962154f
C459 VP.n56 B 0.365734f
C460 VP.n57 B 0.021329f
C461 VP.n58 B 0.021756f
C462 VP.n59 B 0.021756f
C463 VP.n60 B 0.021756f
C464 VP.n61 B 0.040547f
C465 VP.n62 B 0.043759f
C466 VP.n63 B 0.01784f
C467 VP.n64 B 0.021756f
C468 VP.n65 B 0.021756f
C469 VP.n66 B 0.021756f
C470 VP.n67 B 0.040547f
C471 VP.n68 B 0.040547f
C472 VP.n69 B 0.02213f
C473 VP.n70 B 0.035113f
C474 VP.n71 B 1.37297f
C475 VP.n72 B 1.3876f
C476 VP.t7 B 0.962154f
C477 VP.n73 B 0.444116f
C478 VP.n74 B 0.02213f
C479 VP.n75 B 0.035113f
C480 VP.n76 B 0.021756f
C481 VP.n77 B 0.021756f
C482 VP.n78 B 0.040547f
C483 VP.n79 B 0.042467f
C484 VP.n80 B 0.01784f
C485 VP.n81 B 0.021756f
C486 VP.n82 B 0.021756f
C487 VP.n83 B 0.021756f
C488 VP.n84 B 0.040547f
C489 VP.n85 B 0.039746f
C490 VP.n86 B 0.365734f
C491 VP.n87 B 0.021329f
C492 VP.n88 B 0.021756f
C493 VP.n89 B 0.021756f
C494 VP.n90 B 0.021756f
C495 VP.n91 B 0.040547f
C496 VP.n92 B 0.043007f
C497 VP.n93 B 0.017615f
C498 VP.n94 B 0.021756f
C499 VP.n95 B 0.021756f
C500 VP.n96 B 0.021756f
C501 VP.n97 B 0.040547f
C502 VP.n98 B 0.040547f
C503 VP.n99 B 0.386263f
C504 VP.n100 B 0.021756f
C505 VP.n101 B 0.021756f
C506 VP.n102 B 0.021756f
C507 VP.n103 B 0.040547f
C508 VP.n104 B 0.043443f
C509 VP.n105 B 0.017615f
C510 VP.n106 B 0.021756f
C511 VP.n107 B 0.021756f
C512 VP.n108 B 0.021756f
C513 VP.n109 B 0.040547f
C514 VP.n110 B 0.040547f
C515 VP.t4 B 0.962154f
C516 VP.n111 B 0.365734f
C517 VP.n112 B 0.021329f
C518 VP.n113 B 0.021756f
C519 VP.n114 B 0.021756f
C520 VP.n115 B 0.021756f
C521 VP.n116 B 0.040547f
C522 VP.n117 B 0.043759f
C523 VP.n118 B 0.01784f
C524 VP.n119 B 0.021756f
C525 VP.n120 B 0.021756f
C526 VP.n121 B 0.021756f
C527 VP.n122 B 0.040547f
C528 VP.n123 B 0.040547f
C529 VP.n124 B 0.02213f
C530 VP.n125 B 0.035113f
C531 VP.n126 B 0.066063f
.ends

