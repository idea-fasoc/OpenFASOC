* NGSPICE file created from diff_pair_sample_1438.ext - technology: sky130A

.subckt diff_pair_sample_1438 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=0 ps=0 w=6.36 l=2.48
X1 VTAIL.t15 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=1.0494 ps=6.69 w=6.36 l=2.48
X2 VTAIL.t5 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
X3 VTAIL.t14 VN.t1 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
X4 VTAIL.t13 VN.t2 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
X5 VTAIL.t12 VN.t3 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=1.0494 ps=6.69 w=6.36 l=2.48
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=0 ps=0 w=6.36 l=2.48
X7 VTAIL.t2 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=1.0494 ps=6.69 w=6.36 l=2.48
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=0 ps=0 w=6.36 l=2.48
X9 VDD1.t5 VP.t2 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=2.4804 ps=13.5 w=6.36 l=2.48
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=0 ps=0 w=6.36 l=2.48
X11 VDD2.t4 VN.t4 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
X12 VDD1.t4 VP.t3 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
X13 VDD2.t5 VN.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=2.4804 ps=13.5 w=6.36 l=2.48
X14 VDD2.t6 VN.t6 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
X15 VTAIL.t0 VP.t4 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
X16 VTAIL.t6 VP.t5 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4804 pd=13.5 as=1.0494 ps=6.69 w=6.36 l=2.48
X17 VDD1.t1 VP.t6 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=2.4804 ps=13.5 w=6.36 l=2.48
X18 VDD2.t3 VN.t7 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=2.4804 ps=13.5 w=6.36 l=2.48
X19 VDD1.t0 VP.t7 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0494 pd=6.69 as=1.0494 ps=6.69 w=6.36 l=2.48
R0 B.n708 B.n707 585
R1 B.n244 B.n121 585
R2 B.n243 B.n242 585
R3 B.n241 B.n240 585
R4 B.n239 B.n238 585
R5 B.n237 B.n236 585
R6 B.n235 B.n234 585
R7 B.n233 B.n232 585
R8 B.n231 B.n230 585
R9 B.n229 B.n228 585
R10 B.n227 B.n226 585
R11 B.n225 B.n224 585
R12 B.n223 B.n222 585
R13 B.n221 B.n220 585
R14 B.n219 B.n218 585
R15 B.n217 B.n216 585
R16 B.n215 B.n214 585
R17 B.n213 B.n212 585
R18 B.n211 B.n210 585
R19 B.n209 B.n208 585
R20 B.n207 B.n206 585
R21 B.n205 B.n204 585
R22 B.n203 B.n202 585
R23 B.n201 B.n200 585
R24 B.n199 B.n198 585
R25 B.n196 B.n195 585
R26 B.n194 B.n193 585
R27 B.n192 B.n191 585
R28 B.n190 B.n189 585
R29 B.n188 B.n187 585
R30 B.n186 B.n185 585
R31 B.n184 B.n183 585
R32 B.n182 B.n181 585
R33 B.n180 B.n179 585
R34 B.n178 B.n177 585
R35 B.n175 B.n174 585
R36 B.n173 B.n172 585
R37 B.n171 B.n170 585
R38 B.n169 B.n168 585
R39 B.n167 B.n166 585
R40 B.n165 B.n164 585
R41 B.n163 B.n162 585
R42 B.n161 B.n160 585
R43 B.n159 B.n158 585
R44 B.n157 B.n156 585
R45 B.n155 B.n154 585
R46 B.n153 B.n152 585
R47 B.n151 B.n150 585
R48 B.n149 B.n148 585
R49 B.n147 B.n146 585
R50 B.n145 B.n144 585
R51 B.n143 B.n142 585
R52 B.n141 B.n140 585
R53 B.n139 B.n138 585
R54 B.n137 B.n136 585
R55 B.n135 B.n134 585
R56 B.n133 B.n132 585
R57 B.n131 B.n130 585
R58 B.n129 B.n128 585
R59 B.n127 B.n126 585
R60 B.n706 B.n91 585
R61 B.n711 B.n91 585
R62 B.n705 B.n90 585
R63 B.n712 B.n90 585
R64 B.n704 B.n703 585
R65 B.n703 B.n86 585
R66 B.n702 B.n85 585
R67 B.n718 B.n85 585
R68 B.n701 B.n84 585
R69 B.n719 B.n84 585
R70 B.n700 B.n83 585
R71 B.n720 B.n83 585
R72 B.n699 B.n698 585
R73 B.n698 B.n79 585
R74 B.n697 B.n78 585
R75 B.n726 B.n78 585
R76 B.n696 B.n77 585
R77 B.n727 B.n77 585
R78 B.n695 B.n76 585
R79 B.n728 B.n76 585
R80 B.n694 B.n693 585
R81 B.n693 B.n72 585
R82 B.n692 B.n71 585
R83 B.n734 B.n71 585
R84 B.n691 B.n70 585
R85 B.n735 B.n70 585
R86 B.n690 B.n69 585
R87 B.n736 B.n69 585
R88 B.n689 B.n688 585
R89 B.n688 B.n65 585
R90 B.n687 B.n64 585
R91 B.n742 B.n64 585
R92 B.n686 B.n63 585
R93 B.n743 B.n63 585
R94 B.n685 B.n62 585
R95 B.n744 B.n62 585
R96 B.n684 B.n683 585
R97 B.n683 B.n61 585
R98 B.n682 B.n57 585
R99 B.n750 B.n57 585
R100 B.n681 B.n56 585
R101 B.n751 B.n56 585
R102 B.n680 B.n55 585
R103 B.n752 B.n55 585
R104 B.n679 B.n678 585
R105 B.n678 B.n51 585
R106 B.n677 B.n50 585
R107 B.n758 B.n50 585
R108 B.n676 B.n49 585
R109 B.n759 B.n49 585
R110 B.n675 B.n48 585
R111 B.n760 B.n48 585
R112 B.n674 B.n673 585
R113 B.n673 B.n44 585
R114 B.n672 B.n43 585
R115 B.n766 B.n43 585
R116 B.n671 B.n42 585
R117 B.n767 B.n42 585
R118 B.n670 B.n41 585
R119 B.n768 B.n41 585
R120 B.n669 B.n668 585
R121 B.n668 B.n37 585
R122 B.n667 B.n36 585
R123 B.n774 B.n36 585
R124 B.n666 B.n35 585
R125 B.n775 B.n35 585
R126 B.n665 B.n34 585
R127 B.n776 B.n34 585
R128 B.n664 B.n663 585
R129 B.n663 B.n30 585
R130 B.n662 B.n29 585
R131 B.n782 B.n29 585
R132 B.n661 B.n28 585
R133 B.n783 B.n28 585
R134 B.n660 B.n27 585
R135 B.n784 B.n27 585
R136 B.n659 B.n658 585
R137 B.n658 B.n23 585
R138 B.n657 B.n22 585
R139 B.n790 B.n22 585
R140 B.n656 B.n21 585
R141 B.n791 B.n21 585
R142 B.n655 B.n20 585
R143 B.n792 B.n20 585
R144 B.n654 B.n653 585
R145 B.n653 B.n16 585
R146 B.n652 B.n15 585
R147 B.n798 B.n15 585
R148 B.n651 B.n14 585
R149 B.n799 B.n14 585
R150 B.n650 B.n13 585
R151 B.n800 B.n13 585
R152 B.n649 B.n648 585
R153 B.n648 B.n12 585
R154 B.n647 B.n646 585
R155 B.n647 B.n8 585
R156 B.n645 B.n7 585
R157 B.n807 B.n7 585
R158 B.n644 B.n6 585
R159 B.n808 B.n6 585
R160 B.n643 B.n5 585
R161 B.n809 B.n5 585
R162 B.n642 B.n641 585
R163 B.n641 B.n4 585
R164 B.n640 B.n245 585
R165 B.n640 B.n639 585
R166 B.n630 B.n246 585
R167 B.n247 B.n246 585
R168 B.n632 B.n631 585
R169 B.n633 B.n632 585
R170 B.n629 B.n252 585
R171 B.n252 B.n251 585
R172 B.n628 B.n627 585
R173 B.n627 B.n626 585
R174 B.n254 B.n253 585
R175 B.n255 B.n254 585
R176 B.n619 B.n618 585
R177 B.n620 B.n619 585
R178 B.n617 B.n260 585
R179 B.n260 B.n259 585
R180 B.n616 B.n615 585
R181 B.n615 B.n614 585
R182 B.n262 B.n261 585
R183 B.n263 B.n262 585
R184 B.n607 B.n606 585
R185 B.n608 B.n607 585
R186 B.n605 B.n268 585
R187 B.n268 B.n267 585
R188 B.n604 B.n603 585
R189 B.n603 B.n602 585
R190 B.n270 B.n269 585
R191 B.n271 B.n270 585
R192 B.n595 B.n594 585
R193 B.n596 B.n595 585
R194 B.n593 B.n276 585
R195 B.n276 B.n275 585
R196 B.n592 B.n591 585
R197 B.n591 B.n590 585
R198 B.n278 B.n277 585
R199 B.n279 B.n278 585
R200 B.n583 B.n582 585
R201 B.n584 B.n583 585
R202 B.n581 B.n284 585
R203 B.n284 B.n283 585
R204 B.n580 B.n579 585
R205 B.n579 B.n578 585
R206 B.n286 B.n285 585
R207 B.n287 B.n286 585
R208 B.n571 B.n570 585
R209 B.n572 B.n571 585
R210 B.n569 B.n292 585
R211 B.n292 B.n291 585
R212 B.n568 B.n567 585
R213 B.n567 B.n566 585
R214 B.n294 B.n293 585
R215 B.n295 B.n294 585
R216 B.n559 B.n558 585
R217 B.n560 B.n559 585
R218 B.n557 B.n300 585
R219 B.n300 B.n299 585
R220 B.n556 B.n555 585
R221 B.n555 B.n554 585
R222 B.n302 B.n301 585
R223 B.n547 B.n302 585
R224 B.n546 B.n545 585
R225 B.n548 B.n546 585
R226 B.n544 B.n307 585
R227 B.n307 B.n306 585
R228 B.n543 B.n542 585
R229 B.n542 B.n541 585
R230 B.n309 B.n308 585
R231 B.n310 B.n309 585
R232 B.n534 B.n533 585
R233 B.n535 B.n534 585
R234 B.n532 B.n315 585
R235 B.n315 B.n314 585
R236 B.n531 B.n530 585
R237 B.n530 B.n529 585
R238 B.n317 B.n316 585
R239 B.n318 B.n317 585
R240 B.n522 B.n521 585
R241 B.n523 B.n522 585
R242 B.n520 B.n323 585
R243 B.n323 B.n322 585
R244 B.n519 B.n518 585
R245 B.n518 B.n517 585
R246 B.n325 B.n324 585
R247 B.n326 B.n325 585
R248 B.n510 B.n509 585
R249 B.n511 B.n510 585
R250 B.n508 B.n331 585
R251 B.n331 B.n330 585
R252 B.n507 B.n506 585
R253 B.n506 B.n505 585
R254 B.n333 B.n332 585
R255 B.n334 B.n333 585
R256 B.n498 B.n497 585
R257 B.n499 B.n498 585
R258 B.n496 B.n339 585
R259 B.n339 B.n338 585
R260 B.n491 B.n490 585
R261 B.n489 B.n371 585
R262 B.n488 B.n370 585
R263 B.n493 B.n370 585
R264 B.n487 B.n486 585
R265 B.n485 B.n484 585
R266 B.n483 B.n482 585
R267 B.n481 B.n480 585
R268 B.n479 B.n478 585
R269 B.n477 B.n476 585
R270 B.n475 B.n474 585
R271 B.n473 B.n472 585
R272 B.n471 B.n470 585
R273 B.n469 B.n468 585
R274 B.n467 B.n466 585
R275 B.n465 B.n464 585
R276 B.n463 B.n462 585
R277 B.n461 B.n460 585
R278 B.n459 B.n458 585
R279 B.n457 B.n456 585
R280 B.n455 B.n454 585
R281 B.n453 B.n452 585
R282 B.n451 B.n450 585
R283 B.n449 B.n448 585
R284 B.n447 B.n446 585
R285 B.n445 B.n444 585
R286 B.n443 B.n442 585
R287 B.n441 B.n440 585
R288 B.n439 B.n438 585
R289 B.n437 B.n436 585
R290 B.n435 B.n434 585
R291 B.n433 B.n432 585
R292 B.n431 B.n430 585
R293 B.n429 B.n428 585
R294 B.n427 B.n426 585
R295 B.n425 B.n424 585
R296 B.n423 B.n422 585
R297 B.n421 B.n420 585
R298 B.n419 B.n418 585
R299 B.n417 B.n416 585
R300 B.n415 B.n414 585
R301 B.n413 B.n412 585
R302 B.n411 B.n410 585
R303 B.n409 B.n408 585
R304 B.n407 B.n406 585
R305 B.n405 B.n404 585
R306 B.n403 B.n402 585
R307 B.n401 B.n400 585
R308 B.n399 B.n398 585
R309 B.n397 B.n396 585
R310 B.n395 B.n394 585
R311 B.n393 B.n392 585
R312 B.n391 B.n390 585
R313 B.n389 B.n388 585
R314 B.n387 B.n386 585
R315 B.n385 B.n384 585
R316 B.n383 B.n382 585
R317 B.n381 B.n380 585
R318 B.n379 B.n378 585
R319 B.n341 B.n340 585
R320 B.n495 B.n494 585
R321 B.n494 B.n493 585
R322 B.n337 B.n336 585
R323 B.n338 B.n337 585
R324 B.n501 B.n500 585
R325 B.n500 B.n499 585
R326 B.n502 B.n335 585
R327 B.n335 B.n334 585
R328 B.n504 B.n503 585
R329 B.n505 B.n504 585
R330 B.n329 B.n328 585
R331 B.n330 B.n329 585
R332 B.n513 B.n512 585
R333 B.n512 B.n511 585
R334 B.n514 B.n327 585
R335 B.n327 B.n326 585
R336 B.n516 B.n515 585
R337 B.n517 B.n516 585
R338 B.n321 B.n320 585
R339 B.n322 B.n321 585
R340 B.n525 B.n524 585
R341 B.n524 B.n523 585
R342 B.n526 B.n319 585
R343 B.n319 B.n318 585
R344 B.n528 B.n527 585
R345 B.n529 B.n528 585
R346 B.n313 B.n312 585
R347 B.n314 B.n313 585
R348 B.n537 B.n536 585
R349 B.n536 B.n535 585
R350 B.n538 B.n311 585
R351 B.n311 B.n310 585
R352 B.n540 B.n539 585
R353 B.n541 B.n540 585
R354 B.n305 B.n304 585
R355 B.n306 B.n305 585
R356 B.n550 B.n549 585
R357 B.n549 B.n548 585
R358 B.n551 B.n303 585
R359 B.n547 B.n303 585
R360 B.n553 B.n552 585
R361 B.n554 B.n553 585
R362 B.n298 B.n297 585
R363 B.n299 B.n298 585
R364 B.n562 B.n561 585
R365 B.n561 B.n560 585
R366 B.n563 B.n296 585
R367 B.n296 B.n295 585
R368 B.n565 B.n564 585
R369 B.n566 B.n565 585
R370 B.n290 B.n289 585
R371 B.n291 B.n290 585
R372 B.n574 B.n573 585
R373 B.n573 B.n572 585
R374 B.n575 B.n288 585
R375 B.n288 B.n287 585
R376 B.n577 B.n576 585
R377 B.n578 B.n577 585
R378 B.n282 B.n281 585
R379 B.n283 B.n282 585
R380 B.n586 B.n585 585
R381 B.n585 B.n584 585
R382 B.n587 B.n280 585
R383 B.n280 B.n279 585
R384 B.n589 B.n588 585
R385 B.n590 B.n589 585
R386 B.n274 B.n273 585
R387 B.n275 B.n274 585
R388 B.n598 B.n597 585
R389 B.n597 B.n596 585
R390 B.n599 B.n272 585
R391 B.n272 B.n271 585
R392 B.n601 B.n600 585
R393 B.n602 B.n601 585
R394 B.n266 B.n265 585
R395 B.n267 B.n266 585
R396 B.n610 B.n609 585
R397 B.n609 B.n608 585
R398 B.n611 B.n264 585
R399 B.n264 B.n263 585
R400 B.n613 B.n612 585
R401 B.n614 B.n613 585
R402 B.n258 B.n257 585
R403 B.n259 B.n258 585
R404 B.n622 B.n621 585
R405 B.n621 B.n620 585
R406 B.n623 B.n256 585
R407 B.n256 B.n255 585
R408 B.n625 B.n624 585
R409 B.n626 B.n625 585
R410 B.n250 B.n249 585
R411 B.n251 B.n250 585
R412 B.n635 B.n634 585
R413 B.n634 B.n633 585
R414 B.n636 B.n248 585
R415 B.n248 B.n247 585
R416 B.n638 B.n637 585
R417 B.n639 B.n638 585
R418 B.n3 B.n0 585
R419 B.n4 B.n3 585
R420 B.n806 B.n1 585
R421 B.n807 B.n806 585
R422 B.n805 B.n804 585
R423 B.n805 B.n8 585
R424 B.n803 B.n9 585
R425 B.n12 B.n9 585
R426 B.n802 B.n801 585
R427 B.n801 B.n800 585
R428 B.n11 B.n10 585
R429 B.n799 B.n11 585
R430 B.n797 B.n796 585
R431 B.n798 B.n797 585
R432 B.n795 B.n17 585
R433 B.n17 B.n16 585
R434 B.n794 B.n793 585
R435 B.n793 B.n792 585
R436 B.n19 B.n18 585
R437 B.n791 B.n19 585
R438 B.n789 B.n788 585
R439 B.n790 B.n789 585
R440 B.n787 B.n24 585
R441 B.n24 B.n23 585
R442 B.n786 B.n785 585
R443 B.n785 B.n784 585
R444 B.n26 B.n25 585
R445 B.n783 B.n26 585
R446 B.n781 B.n780 585
R447 B.n782 B.n781 585
R448 B.n779 B.n31 585
R449 B.n31 B.n30 585
R450 B.n778 B.n777 585
R451 B.n777 B.n776 585
R452 B.n33 B.n32 585
R453 B.n775 B.n33 585
R454 B.n773 B.n772 585
R455 B.n774 B.n773 585
R456 B.n771 B.n38 585
R457 B.n38 B.n37 585
R458 B.n770 B.n769 585
R459 B.n769 B.n768 585
R460 B.n40 B.n39 585
R461 B.n767 B.n40 585
R462 B.n765 B.n764 585
R463 B.n766 B.n765 585
R464 B.n763 B.n45 585
R465 B.n45 B.n44 585
R466 B.n762 B.n761 585
R467 B.n761 B.n760 585
R468 B.n47 B.n46 585
R469 B.n759 B.n47 585
R470 B.n757 B.n756 585
R471 B.n758 B.n757 585
R472 B.n755 B.n52 585
R473 B.n52 B.n51 585
R474 B.n754 B.n753 585
R475 B.n753 B.n752 585
R476 B.n54 B.n53 585
R477 B.n751 B.n54 585
R478 B.n749 B.n748 585
R479 B.n750 B.n749 585
R480 B.n747 B.n58 585
R481 B.n61 B.n58 585
R482 B.n746 B.n745 585
R483 B.n745 B.n744 585
R484 B.n60 B.n59 585
R485 B.n743 B.n60 585
R486 B.n741 B.n740 585
R487 B.n742 B.n741 585
R488 B.n739 B.n66 585
R489 B.n66 B.n65 585
R490 B.n738 B.n737 585
R491 B.n737 B.n736 585
R492 B.n68 B.n67 585
R493 B.n735 B.n68 585
R494 B.n733 B.n732 585
R495 B.n734 B.n733 585
R496 B.n731 B.n73 585
R497 B.n73 B.n72 585
R498 B.n730 B.n729 585
R499 B.n729 B.n728 585
R500 B.n75 B.n74 585
R501 B.n727 B.n75 585
R502 B.n725 B.n724 585
R503 B.n726 B.n725 585
R504 B.n723 B.n80 585
R505 B.n80 B.n79 585
R506 B.n722 B.n721 585
R507 B.n721 B.n720 585
R508 B.n82 B.n81 585
R509 B.n719 B.n82 585
R510 B.n717 B.n716 585
R511 B.n718 B.n717 585
R512 B.n715 B.n87 585
R513 B.n87 B.n86 585
R514 B.n714 B.n713 585
R515 B.n713 B.n712 585
R516 B.n89 B.n88 585
R517 B.n711 B.n89 585
R518 B.n810 B.n809 585
R519 B.n808 B.n2 585
R520 B.n126 B.n89 458.866
R521 B.n708 B.n91 458.866
R522 B.n494 B.n339 458.866
R523 B.n491 B.n337 458.866
R524 B.n124 B.t16 269.663
R525 B.n122 B.t8 269.663
R526 B.n375 B.t12 269.663
R527 B.n372 B.t19 269.663
R528 B.n710 B.n709 256.663
R529 B.n710 B.n120 256.663
R530 B.n710 B.n119 256.663
R531 B.n710 B.n118 256.663
R532 B.n710 B.n117 256.663
R533 B.n710 B.n116 256.663
R534 B.n710 B.n115 256.663
R535 B.n710 B.n114 256.663
R536 B.n710 B.n113 256.663
R537 B.n710 B.n112 256.663
R538 B.n710 B.n111 256.663
R539 B.n710 B.n110 256.663
R540 B.n710 B.n109 256.663
R541 B.n710 B.n108 256.663
R542 B.n710 B.n107 256.663
R543 B.n710 B.n106 256.663
R544 B.n710 B.n105 256.663
R545 B.n710 B.n104 256.663
R546 B.n710 B.n103 256.663
R547 B.n710 B.n102 256.663
R548 B.n710 B.n101 256.663
R549 B.n710 B.n100 256.663
R550 B.n710 B.n99 256.663
R551 B.n710 B.n98 256.663
R552 B.n710 B.n97 256.663
R553 B.n710 B.n96 256.663
R554 B.n710 B.n95 256.663
R555 B.n710 B.n94 256.663
R556 B.n710 B.n93 256.663
R557 B.n710 B.n92 256.663
R558 B.n493 B.n492 256.663
R559 B.n493 B.n342 256.663
R560 B.n493 B.n343 256.663
R561 B.n493 B.n344 256.663
R562 B.n493 B.n345 256.663
R563 B.n493 B.n346 256.663
R564 B.n493 B.n347 256.663
R565 B.n493 B.n348 256.663
R566 B.n493 B.n349 256.663
R567 B.n493 B.n350 256.663
R568 B.n493 B.n351 256.663
R569 B.n493 B.n352 256.663
R570 B.n493 B.n353 256.663
R571 B.n493 B.n354 256.663
R572 B.n493 B.n355 256.663
R573 B.n493 B.n356 256.663
R574 B.n493 B.n357 256.663
R575 B.n493 B.n358 256.663
R576 B.n493 B.n359 256.663
R577 B.n493 B.n360 256.663
R578 B.n493 B.n361 256.663
R579 B.n493 B.n362 256.663
R580 B.n493 B.n363 256.663
R581 B.n493 B.n364 256.663
R582 B.n493 B.n365 256.663
R583 B.n493 B.n366 256.663
R584 B.n493 B.n367 256.663
R585 B.n493 B.n368 256.663
R586 B.n493 B.n369 256.663
R587 B.n812 B.n811 256.663
R588 B.n130 B.n129 163.367
R589 B.n134 B.n133 163.367
R590 B.n138 B.n137 163.367
R591 B.n142 B.n141 163.367
R592 B.n146 B.n145 163.367
R593 B.n150 B.n149 163.367
R594 B.n154 B.n153 163.367
R595 B.n158 B.n157 163.367
R596 B.n162 B.n161 163.367
R597 B.n166 B.n165 163.367
R598 B.n170 B.n169 163.367
R599 B.n174 B.n173 163.367
R600 B.n179 B.n178 163.367
R601 B.n183 B.n182 163.367
R602 B.n187 B.n186 163.367
R603 B.n191 B.n190 163.367
R604 B.n195 B.n194 163.367
R605 B.n200 B.n199 163.367
R606 B.n204 B.n203 163.367
R607 B.n208 B.n207 163.367
R608 B.n212 B.n211 163.367
R609 B.n216 B.n215 163.367
R610 B.n220 B.n219 163.367
R611 B.n224 B.n223 163.367
R612 B.n228 B.n227 163.367
R613 B.n232 B.n231 163.367
R614 B.n236 B.n235 163.367
R615 B.n240 B.n239 163.367
R616 B.n242 B.n121 163.367
R617 B.n498 B.n339 163.367
R618 B.n498 B.n333 163.367
R619 B.n506 B.n333 163.367
R620 B.n506 B.n331 163.367
R621 B.n510 B.n331 163.367
R622 B.n510 B.n325 163.367
R623 B.n518 B.n325 163.367
R624 B.n518 B.n323 163.367
R625 B.n522 B.n323 163.367
R626 B.n522 B.n317 163.367
R627 B.n530 B.n317 163.367
R628 B.n530 B.n315 163.367
R629 B.n534 B.n315 163.367
R630 B.n534 B.n309 163.367
R631 B.n542 B.n309 163.367
R632 B.n542 B.n307 163.367
R633 B.n546 B.n307 163.367
R634 B.n546 B.n302 163.367
R635 B.n555 B.n302 163.367
R636 B.n555 B.n300 163.367
R637 B.n559 B.n300 163.367
R638 B.n559 B.n294 163.367
R639 B.n567 B.n294 163.367
R640 B.n567 B.n292 163.367
R641 B.n571 B.n292 163.367
R642 B.n571 B.n286 163.367
R643 B.n579 B.n286 163.367
R644 B.n579 B.n284 163.367
R645 B.n583 B.n284 163.367
R646 B.n583 B.n278 163.367
R647 B.n591 B.n278 163.367
R648 B.n591 B.n276 163.367
R649 B.n595 B.n276 163.367
R650 B.n595 B.n270 163.367
R651 B.n603 B.n270 163.367
R652 B.n603 B.n268 163.367
R653 B.n607 B.n268 163.367
R654 B.n607 B.n262 163.367
R655 B.n615 B.n262 163.367
R656 B.n615 B.n260 163.367
R657 B.n619 B.n260 163.367
R658 B.n619 B.n254 163.367
R659 B.n627 B.n254 163.367
R660 B.n627 B.n252 163.367
R661 B.n632 B.n252 163.367
R662 B.n632 B.n246 163.367
R663 B.n640 B.n246 163.367
R664 B.n641 B.n640 163.367
R665 B.n641 B.n5 163.367
R666 B.n6 B.n5 163.367
R667 B.n7 B.n6 163.367
R668 B.n647 B.n7 163.367
R669 B.n648 B.n647 163.367
R670 B.n648 B.n13 163.367
R671 B.n14 B.n13 163.367
R672 B.n15 B.n14 163.367
R673 B.n653 B.n15 163.367
R674 B.n653 B.n20 163.367
R675 B.n21 B.n20 163.367
R676 B.n22 B.n21 163.367
R677 B.n658 B.n22 163.367
R678 B.n658 B.n27 163.367
R679 B.n28 B.n27 163.367
R680 B.n29 B.n28 163.367
R681 B.n663 B.n29 163.367
R682 B.n663 B.n34 163.367
R683 B.n35 B.n34 163.367
R684 B.n36 B.n35 163.367
R685 B.n668 B.n36 163.367
R686 B.n668 B.n41 163.367
R687 B.n42 B.n41 163.367
R688 B.n43 B.n42 163.367
R689 B.n673 B.n43 163.367
R690 B.n673 B.n48 163.367
R691 B.n49 B.n48 163.367
R692 B.n50 B.n49 163.367
R693 B.n678 B.n50 163.367
R694 B.n678 B.n55 163.367
R695 B.n56 B.n55 163.367
R696 B.n57 B.n56 163.367
R697 B.n683 B.n57 163.367
R698 B.n683 B.n62 163.367
R699 B.n63 B.n62 163.367
R700 B.n64 B.n63 163.367
R701 B.n688 B.n64 163.367
R702 B.n688 B.n69 163.367
R703 B.n70 B.n69 163.367
R704 B.n71 B.n70 163.367
R705 B.n693 B.n71 163.367
R706 B.n693 B.n76 163.367
R707 B.n77 B.n76 163.367
R708 B.n78 B.n77 163.367
R709 B.n698 B.n78 163.367
R710 B.n698 B.n83 163.367
R711 B.n84 B.n83 163.367
R712 B.n85 B.n84 163.367
R713 B.n703 B.n85 163.367
R714 B.n703 B.n90 163.367
R715 B.n91 B.n90 163.367
R716 B.n371 B.n370 163.367
R717 B.n486 B.n370 163.367
R718 B.n484 B.n483 163.367
R719 B.n480 B.n479 163.367
R720 B.n476 B.n475 163.367
R721 B.n472 B.n471 163.367
R722 B.n468 B.n467 163.367
R723 B.n464 B.n463 163.367
R724 B.n460 B.n459 163.367
R725 B.n456 B.n455 163.367
R726 B.n452 B.n451 163.367
R727 B.n448 B.n447 163.367
R728 B.n444 B.n443 163.367
R729 B.n440 B.n439 163.367
R730 B.n436 B.n435 163.367
R731 B.n432 B.n431 163.367
R732 B.n428 B.n427 163.367
R733 B.n424 B.n423 163.367
R734 B.n420 B.n419 163.367
R735 B.n416 B.n415 163.367
R736 B.n412 B.n411 163.367
R737 B.n408 B.n407 163.367
R738 B.n404 B.n403 163.367
R739 B.n400 B.n399 163.367
R740 B.n396 B.n395 163.367
R741 B.n392 B.n391 163.367
R742 B.n388 B.n387 163.367
R743 B.n384 B.n383 163.367
R744 B.n380 B.n379 163.367
R745 B.n494 B.n341 163.367
R746 B.n500 B.n337 163.367
R747 B.n500 B.n335 163.367
R748 B.n504 B.n335 163.367
R749 B.n504 B.n329 163.367
R750 B.n512 B.n329 163.367
R751 B.n512 B.n327 163.367
R752 B.n516 B.n327 163.367
R753 B.n516 B.n321 163.367
R754 B.n524 B.n321 163.367
R755 B.n524 B.n319 163.367
R756 B.n528 B.n319 163.367
R757 B.n528 B.n313 163.367
R758 B.n536 B.n313 163.367
R759 B.n536 B.n311 163.367
R760 B.n540 B.n311 163.367
R761 B.n540 B.n305 163.367
R762 B.n549 B.n305 163.367
R763 B.n549 B.n303 163.367
R764 B.n553 B.n303 163.367
R765 B.n553 B.n298 163.367
R766 B.n561 B.n298 163.367
R767 B.n561 B.n296 163.367
R768 B.n565 B.n296 163.367
R769 B.n565 B.n290 163.367
R770 B.n573 B.n290 163.367
R771 B.n573 B.n288 163.367
R772 B.n577 B.n288 163.367
R773 B.n577 B.n282 163.367
R774 B.n585 B.n282 163.367
R775 B.n585 B.n280 163.367
R776 B.n589 B.n280 163.367
R777 B.n589 B.n274 163.367
R778 B.n597 B.n274 163.367
R779 B.n597 B.n272 163.367
R780 B.n601 B.n272 163.367
R781 B.n601 B.n266 163.367
R782 B.n609 B.n266 163.367
R783 B.n609 B.n264 163.367
R784 B.n613 B.n264 163.367
R785 B.n613 B.n258 163.367
R786 B.n621 B.n258 163.367
R787 B.n621 B.n256 163.367
R788 B.n625 B.n256 163.367
R789 B.n625 B.n250 163.367
R790 B.n634 B.n250 163.367
R791 B.n634 B.n248 163.367
R792 B.n638 B.n248 163.367
R793 B.n638 B.n3 163.367
R794 B.n810 B.n3 163.367
R795 B.n806 B.n2 163.367
R796 B.n806 B.n805 163.367
R797 B.n805 B.n9 163.367
R798 B.n801 B.n9 163.367
R799 B.n801 B.n11 163.367
R800 B.n797 B.n11 163.367
R801 B.n797 B.n17 163.367
R802 B.n793 B.n17 163.367
R803 B.n793 B.n19 163.367
R804 B.n789 B.n19 163.367
R805 B.n789 B.n24 163.367
R806 B.n785 B.n24 163.367
R807 B.n785 B.n26 163.367
R808 B.n781 B.n26 163.367
R809 B.n781 B.n31 163.367
R810 B.n777 B.n31 163.367
R811 B.n777 B.n33 163.367
R812 B.n773 B.n33 163.367
R813 B.n773 B.n38 163.367
R814 B.n769 B.n38 163.367
R815 B.n769 B.n40 163.367
R816 B.n765 B.n40 163.367
R817 B.n765 B.n45 163.367
R818 B.n761 B.n45 163.367
R819 B.n761 B.n47 163.367
R820 B.n757 B.n47 163.367
R821 B.n757 B.n52 163.367
R822 B.n753 B.n52 163.367
R823 B.n753 B.n54 163.367
R824 B.n749 B.n54 163.367
R825 B.n749 B.n58 163.367
R826 B.n745 B.n58 163.367
R827 B.n745 B.n60 163.367
R828 B.n741 B.n60 163.367
R829 B.n741 B.n66 163.367
R830 B.n737 B.n66 163.367
R831 B.n737 B.n68 163.367
R832 B.n733 B.n68 163.367
R833 B.n733 B.n73 163.367
R834 B.n729 B.n73 163.367
R835 B.n729 B.n75 163.367
R836 B.n725 B.n75 163.367
R837 B.n725 B.n80 163.367
R838 B.n721 B.n80 163.367
R839 B.n721 B.n82 163.367
R840 B.n717 B.n82 163.367
R841 B.n717 B.n87 163.367
R842 B.n713 B.n87 163.367
R843 B.n713 B.n89 163.367
R844 B.n122 B.t10 128.407
R845 B.n375 B.t15 128.407
R846 B.n124 B.t17 128.401
R847 B.n372 B.t21 128.401
R848 B.n493 B.n338 112.505
R849 B.n711 B.n710 112.505
R850 B.n123 B.t11 73.9109
R851 B.n376 B.t14 73.9109
R852 B.n125 B.t18 73.9041
R853 B.n373 B.t20 73.9041
R854 B.n126 B.n92 71.676
R855 B.n130 B.n93 71.676
R856 B.n134 B.n94 71.676
R857 B.n138 B.n95 71.676
R858 B.n142 B.n96 71.676
R859 B.n146 B.n97 71.676
R860 B.n150 B.n98 71.676
R861 B.n154 B.n99 71.676
R862 B.n158 B.n100 71.676
R863 B.n162 B.n101 71.676
R864 B.n166 B.n102 71.676
R865 B.n170 B.n103 71.676
R866 B.n174 B.n104 71.676
R867 B.n179 B.n105 71.676
R868 B.n183 B.n106 71.676
R869 B.n187 B.n107 71.676
R870 B.n191 B.n108 71.676
R871 B.n195 B.n109 71.676
R872 B.n200 B.n110 71.676
R873 B.n204 B.n111 71.676
R874 B.n208 B.n112 71.676
R875 B.n212 B.n113 71.676
R876 B.n216 B.n114 71.676
R877 B.n220 B.n115 71.676
R878 B.n224 B.n116 71.676
R879 B.n228 B.n117 71.676
R880 B.n232 B.n118 71.676
R881 B.n236 B.n119 71.676
R882 B.n240 B.n120 71.676
R883 B.n709 B.n121 71.676
R884 B.n709 B.n708 71.676
R885 B.n242 B.n120 71.676
R886 B.n239 B.n119 71.676
R887 B.n235 B.n118 71.676
R888 B.n231 B.n117 71.676
R889 B.n227 B.n116 71.676
R890 B.n223 B.n115 71.676
R891 B.n219 B.n114 71.676
R892 B.n215 B.n113 71.676
R893 B.n211 B.n112 71.676
R894 B.n207 B.n111 71.676
R895 B.n203 B.n110 71.676
R896 B.n199 B.n109 71.676
R897 B.n194 B.n108 71.676
R898 B.n190 B.n107 71.676
R899 B.n186 B.n106 71.676
R900 B.n182 B.n105 71.676
R901 B.n178 B.n104 71.676
R902 B.n173 B.n103 71.676
R903 B.n169 B.n102 71.676
R904 B.n165 B.n101 71.676
R905 B.n161 B.n100 71.676
R906 B.n157 B.n99 71.676
R907 B.n153 B.n98 71.676
R908 B.n149 B.n97 71.676
R909 B.n145 B.n96 71.676
R910 B.n141 B.n95 71.676
R911 B.n137 B.n94 71.676
R912 B.n133 B.n93 71.676
R913 B.n129 B.n92 71.676
R914 B.n492 B.n491 71.676
R915 B.n486 B.n342 71.676
R916 B.n483 B.n343 71.676
R917 B.n479 B.n344 71.676
R918 B.n475 B.n345 71.676
R919 B.n471 B.n346 71.676
R920 B.n467 B.n347 71.676
R921 B.n463 B.n348 71.676
R922 B.n459 B.n349 71.676
R923 B.n455 B.n350 71.676
R924 B.n451 B.n351 71.676
R925 B.n447 B.n352 71.676
R926 B.n443 B.n353 71.676
R927 B.n439 B.n354 71.676
R928 B.n435 B.n355 71.676
R929 B.n431 B.n356 71.676
R930 B.n427 B.n357 71.676
R931 B.n423 B.n358 71.676
R932 B.n419 B.n359 71.676
R933 B.n415 B.n360 71.676
R934 B.n411 B.n361 71.676
R935 B.n407 B.n362 71.676
R936 B.n403 B.n363 71.676
R937 B.n399 B.n364 71.676
R938 B.n395 B.n365 71.676
R939 B.n391 B.n366 71.676
R940 B.n387 B.n367 71.676
R941 B.n383 B.n368 71.676
R942 B.n379 B.n369 71.676
R943 B.n492 B.n371 71.676
R944 B.n484 B.n342 71.676
R945 B.n480 B.n343 71.676
R946 B.n476 B.n344 71.676
R947 B.n472 B.n345 71.676
R948 B.n468 B.n346 71.676
R949 B.n464 B.n347 71.676
R950 B.n460 B.n348 71.676
R951 B.n456 B.n349 71.676
R952 B.n452 B.n350 71.676
R953 B.n448 B.n351 71.676
R954 B.n444 B.n352 71.676
R955 B.n440 B.n353 71.676
R956 B.n436 B.n354 71.676
R957 B.n432 B.n355 71.676
R958 B.n428 B.n356 71.676
R959 B.n424 B.n357 71.676
R960 B.n420 B.n358 71.676
R961 B.n416 B.n359 71.676
R962 B.n412 B.n360 71.676
R963 B.n408 B.n361 71.676
R964 B.n404 B.n362 71.676
R965 B.n400 B.n363 71.676
R966 B.n396 B.n364 71.676
R967 B.n392 B.n365 71.676
R968 B.n388 B.n366 71.676
R969 B.n384 B.n367 71.676
R970 B.n380 B.n368 71.676
R971 B.n369 B.n341 71.676
R972 B.n811 B.n810 71.676
R973 B.n811 B.n2 71.676
R974 B.n499 B.n338 64.2893
R975 B.n499 B.n334 64.2893
R976 B.n505 B.n334 64.2893
R977 B.n505 B.n330 64.2893
R978 B.n511 B.n330 64.2893
R979 B.n511 B.n326 64.2893
R980 B.n517 B.n326 64.2893
R981 B.n523 B.n322 64.2893
R982 B.n523 B.n318 64.2893
R983 B.n529 B.n318 64.2893
R984 B.n529 B.n314 64.2893
R985 B.n535 B.n314 64.2893
R986 B.n535 B.n310 64.2893
R987 B.n541 B.n310 64.2893
R988 B.n541 B.n306 64.2893
R989 B.n548 B.n306 64.2893
R990 B.n548 B.n547 64.2893
R991 B.n554 B.n299 64.2893
R992 B.n560 B.n299 64.2893
R993 B.n560 B.n295 64.2893
R994 B.n566 B.n295 64.2893
R995 B.n566 B.n291 64.2893
R996 B.n572 B.n291 64.2893
R997 B.n572 B.n287 64.2893
R998 B.n578 B.n287 64.2893
R999 B.n584 B.n283 64.2893
R1000 B.n584 B.n279 64.2893
R1001 B.n590 B.n279 64.2893
R1002 B.n590 B.n275 64.2893
R1003 B.n596 B.n275 64.2893
R1004 B.n596 B.n271 64.2893
R1005 B.n602 B.n271 64.2893
R1006 B.n608 B.n267 64.2893
R1007 B.n608 B.n263 64.2893
R1008 B.n614 B.n263 64.2893
R1009 B.n614 B.n259 64.2893
R1010 B.n620 B.n259 64.2893
R1011 B.n620 B.n255 64.2893
R1012 B.n626 B.n255 64.2893
R1013 B.n633 B.n251 64.2893
R1014 B.n633 B.n247 64.2893
R1015 B.n639 B.n247 64.2893
R1016 B.n639 B.n4 64.2893
R1017 B.n809 B.n4 64.2893
R1018 B.n809 B.n808 64.2893
R1019 B.n808 B.n807 64.2893
R1020 B.n807 B.n8 64.2893
R1021 B.n12 B.n8 64.2893
R1022 B.n800 B.n12 64.2893
R1023 B.n800 B.n799 64.2893
R1024 B.n798 B.n16 64.2893
R1025 B.n792 B.n16 64.2893
R1026 B.n792 B.n791 64.2893
R1027 B.n791 B.n790 64.2893
R1028 B.n790 B.n23 64.2893
R1029 B.n784 B.n23 64.2893
R1030 B.n784 B.n783 64.2893
R1031 B.n782 B.n30 64.2893
R1032 B.n776 B.n30 64.2893
R1033 B.n776 B.n775 64.2893
R1034 B.n775 B.n774 64.2893
R1035 B.n774 B.n37 64.2893
R1036 B.n768 B.n37 64.2893
R1037 B.n768 B.n767 64.2893
R1038 B.n766 B.n44 64.2893
R1039 B.n760 B.n44 64.2893
R1040 B.n760 B.n759 64.2893
R1041 B.n759 B.n758 64.2893
R1042 B.n758 B.n51 64.2893
R1043 B.n752 B.n51 64.2893
R1044 B.n752 B.n751 64.2893
R1045 B.n751 B.n750 64.2893
R1046 B.n744 B.n61 64.2893
R1047 B.n744 B.n743 64.2893
R1048 B.n743 B.n742 64.2893
R1049 B.n742 B.n65 64.2893
R1050 B.n736 B.n65 64.2893
R1051 B.n736 B.n735 64.2893
R1052 B.n735 B.n734 64.2893
R1053 B.n734 B.n72 64.2893
R1054 B.n728 B.n72 64.2893
R1055 B.n728 B.n727 64.2893
R1056 B.n726 B.n79 64.2893
R1057 B.n720 B.n79 64.2893
R1058 B.n720 B.n719 64.2893
R1059 B.n719 B.n718 64.2893
R1060 B.n718 B.n86 64.2893
R1061 B.n712 B.n86 64.2893
R1062 B.n712 B.n711 64.2893
R1063 B.n547 B.t5 62.3984
R1064 B.n61 B.t7 62.3984
R1065 B.n176 B.n125 59.5399
R1066 B.n197 B.n123 59.5399
R1067 B.n377 B.n376 59.5399
R1068 B.n374 B.n373 59.5399
R1069 B.n125 B.n124 54.4975
R1070 B.n123 B.n122 54.4975
R1071 B.n376 B.n375 54.4975
R1072 B.n373 B.n372 54.4975
R1073 B.t4 B.n283 49.1625
R1074 B.n626 B.t0 49.1625
R1075 B.t6 B.n798 49.1625
R1076 B.n767 B.t2 49.1625
R1077 B.n517 B.t13 32.1449
R1078 B.t13 B.n322 32.1449
R1079 B.n602 B.t3 32.1449
R1080 B.t3 B.n267 32.1449
R1081 B.n783 B.t1 32.1449
R1082 B.t1 B.n782 32.1449
R1083 B.n727 B.t9 32.1449
R1084 B.t9 B.n726 32.1449
R1085 B.n490 B.n336 29.8151
R1086 B.n496 B.n495 29.8151
R1087 B.n707 B.n706 29.8151
R1088 B.n127 B.n88 29.8151
R1089 B B.n812 18.0485
R1090 B.n578 B.t4 15.1273
R1091 B.t0 B.n251 15.1273
R1092 B.n799 B.t6 15.1273
R1093 B.t2 B.n766 15.1273
R1094 B.n501 B.n336 10.6151
R1095 B.n502 B.n501 10.6151
R1096 B.n503 B.n502 10.6151
R1097 B.n503 B.n328 10.6151
R1098 B.n513 B.n328 10.6151
R1099 B.n514 B.n513 10.6151
R1100 B.n515 B.n514 10.6151
R1101 B.n515 B.n320 10.6151
R1102 B.n525 B.n320 10.6151
R1103 B.n526 B.n525 10.6151
R1104 B.n527 B.n526 10.6151
R1105 B.n527 B.n312 10.6151
R1106 B.n537 B.n312 10.6151
R1107 B.n538 B.n537 10.6151
R1108 B.n539 B.n538 10.6151
R1109 B.n539 B.n304 10.6151
R1110 B.n550 B.n304 10.6151
R1111 B.n551 B.n550 10.6151
R1112 B.n552 B.n551 10.6151
R1113 B.n552 B.n297 10.6151
R1114 B.n562 B.n297 10.6151
R1115 B.n563 B.n562 10.6151
R1116 B.n564 B.n563 10.6151
R1117 B.n564 B.n289 10.6151
R1118 B.n574 B.n289 10.6151
R1119 B.n575 B.n574 10.6151
R1120 B.n576 B.n575 10.6151
R1121 B.n576 B.n281 10.6151
R1122 B.n586 B.n281 10.6151
R1123 B.n587 B.n586 10.6151
R1124 B.n588 B.n587 10.6151
R1125 B.n588 B.n273 10.6151
R1126 B.n598 B.n273 10.6151
R1127 B.n599 B.n598 10.6151
R1128 B.n600 B.n599 10.6151
R1129 B.n600 B.n265 10.6151
R1130 B.n610 B.n265 10.6151
R1131 B.n611 B.n610 10.6151
R1132 B.n612 B.n611 10.6151
R1133 B.n612 B.n257 10.6151
R1134 B.n622 B.n257 10.6151
R1135 B.n623 B.n622 10.6151
R1136 B.n624 B.n623 10.6151
R1137 B.n624 B.n249 10.6151
R1138 B.n635 B.n249 10.6151
R1139 B.n636 B.n635 10.6151
R1140 B.n637 B.n636 10.6151
R1141 B.n637 B.n0 10.6151
R1142 B.n490 B.n489 10.6151
R1143 B.n489 B.n488 10.6151
R1144 B.n488 B.n487 10.6151
R1145 B.n487 B.n485 10.6151
R1146 B.n485 B.n482 10.6151
R1147 B.n482 B.n481 10.6151
R1148 B.n481 B.n478 10.6151
R1149 B.n478 B.n477 10.6151
R1150 B.n477 B.n474 10.6151
R1151 B.n474 B.n473 10.6151
R1152 B.n473 B.n470 10.6151
R1153 B.n470 B.n469 10.6151
R1154 B.n469 B.n466 10.6151
R1155 B.n466 B.n465 10.6151
R1156 B.n465 B.n462 10.6151
R1157 B.n462 B.n461 10.6151
R1158 B.n461 B.n458 10.6151
R1159 B.n458 B.n457 10.6151
R1160 B.n457 B.n454 10.6151
R1161 B.n454 B.n453 10.6151
R1162 B.n453 B.n450 10.6151
R1163 B.n450 B.n449 10.6151
R1164 B.n449 B.n446 10.6151
R1165 B.n446 B.n445 10.6151
R1166 B.n442 B.n441 10.6151
R1167 B.n441 B.n438 10.6151
R1168 B.n438 B.n437 10.6151
R1169 B.n437 B.n434 10.6151
R1170 B.n434 B.n433 10.6151
R1171 B.n433 B.n430 10.6151
R1172 B.n430 B.n429 10.6151
R1173 B.n429 B.n426 10.6151
R1174 B.n426 B.n425 10.6151
R1175 B.n422 B.n421 10.6151
R1176 B.n421 B.n418 10.6151
R1177 B.n418 B.n417 10.6151
R1178 B.n417 B.n414 10.6151
R1179 B.n414 B.n413 10.6151
R1180 B.n413 B.n410 10.6151
R1181 B.n410 B.n409 10.6151
R1182 B.n409 B.n406 10.6151
R1183 B.n406 B.n405 10.6151
R1184 B.n405 B.n402 10.6151
R1185 B.n402 B.n401 10.6151
R1186 B.n401 B.n398 10.6151
R1187 B.n398 B.n397 10.6151
R1188 B.n397 B.n394 10.6151
R1189 B.n394 B.n393 10.6151
R1190 B.n393 B.n390 10.6151
R1191 B.n390 B.n389 10.6151
R1192 B.n389 B.n386 10.6151
R1193 B.n386 B.n385 10.6151
R1194 B.n385 B.n382 10.6151
R1195 B.n382 B.n381 10.6151
R1196 B.n381 B.n378 10.6151
R1197 B.n378 B.n340 10.6151
R1198 B.n495 B.n340 10.6151
R1199 B.n497 B.n496 10.6151
R1200 B.n497 B.n332 10.6151
R1201 B.n507 B.n332 10.6151
R1202 B.n508 B.n507 10.6151
R1203 B.n509 B.n508 10.6151
R1204 B.n509 B.n324 10.6151
R1205 B.n519 B.n324 10.6151
R1206 B.n520 B.n519 10.6151
R1207 B.n521 B.n520 10.6151
R1208 B.n521 B.n316 10.6151
R1209 B.n531 B.n316 10.6151
R1210 B.n532 B.n531 10.6151
R1211 B.n533 B.n532 10.6151
R1212 B.n533 B.n308 10.6151
R1213 B.n543 B.n308 10.6151
R1214 B.n544 B.n543 10.6151
R1215 B.n545 B.n544 10.6151
R1216 B.n545 B.n301 10.6151
R1217 B.n556 B.n301 10.6151
R1218 B.n557 B.n556 10.6151
R1219 B.n558 B.n557 10.6151
R1220 B.n558 B.n293 10.6151
R1221 B.n568 B.n293 10.6151
R1222 B.n569 B.n568 10.6151
R1223 B.n570 B.n569 10.6151
R1224 B.n570 B.n285 10.6151
R1225 B.n580 B.n285 10.6151
R1226 B.n581 B.n580 10.6151
R1227 B.n582 B.n581 10.6151
R1228 B.n582 B.n277 10.6151
R1229 B.n592 B.n277 10.6151
R1230 B.n593 B.n592 10.6151
R1231 B.n594 B.n593 10.6151
R1232 B.n594 B.n269 10.6151
R1233 B.n604 B.n269 10.6151
R1234 B.n605 B.n604 10.6151
R1235 B.n606 B.n605 10.6151
R1236 B.n606 B.n261 10.6151
R1237 B.n616 B.n261 10.6151
R1238 B.n617 B.n616 10.6151
R1239 B.n618 B.n617 10.6151
R1240 B.n618 B.n253 10.6151
R1241 B.n628 B.n253 10.6151
R1242 B.n629 B.n628 10.6151
R1243 B.n631 B.n629 10.6151
R1244 B.n631 B.n630 10.6151
R1245 B.n630 B.n245 10.6151
R1246 B.n642 B.n245 10.6151
R1247 B.n643 B.n642 10.6151
R1248 B.n644 B.n643 10.6151
R1249 B.n645 B.n644 10.6151
R1250 B.n646 B.n645 10.6151
R1251 B.n649 B.n646 10.6151
R1252 B.n650 B.n649 10.6151
R1253 B.n651 B.n650 10.6151
R1254 B.n652 B.n651 10.6151
R1255 B.n654 B.n652 10.6151
R1256 B.n655 B.n654 10.6151
R1257 B.n656 B.n655 10.6151
R1258 B.n657 B.n656 10.6151
R1259 B.n659 B.n657 10.6151
R1260 B.n660 B.n659 10.6151
R1261 B.n661 B.n660 10.6151
R1262 B.n662 B.n661 10.6151
R1263 B.n664 B.n662 10.6151
R1264 B.n665 B.n664 10.6151
R1265 B.n666 B.n665 10.6151
R1266 B.n667 B.n666 10.6151
R1267 B.n669 B.n667 10.6151
R1268 B.n670 B.n669 10.6151
R1269 B.n671 B.n670 10.6151
R1270 B.n672 B.n671 10.6151
R1271 B.n674 B.n672 10.6151
R1272 B.n675 B.n674 10.6151
R1273 B.n676 B.n675 10.6151
R1274 B.n677 B.n676 10.6151
R1275 B.n679 B.n677 10.6151
R1276 B.n680 B.n679 10.6151
R1277 B.n681 B.n680 10.6151
R1278 B.n682 B.n681 10.6151
R1279 B.n684 B.n682 10.6151
R1280 B.n685 B.n684 10.6151
R1281 B.n686 B.n685 10.6151
R1282 B.n687 B.n686 10.6151
R1283 B.n689 B.n687 10.6151
R1284 B.n690 B.n689 10.6151
R1285 B.n691 B.n690 10.6151
R1286 B.n692 B.n691 10.6151
R1287 B.n694 B.n692 10.6151
R1288 B.n695 B.n694 10.6151
R1289 B.n696 B.n695 10.6151
R1290 B.n697 B.n696 10.6151
R1291 B.n699 B.n697 10.6151
R1292 B.n700 B.n699 10.6151
R1293 B.n701 B.n700 10.6151
R1294 B.n702 B.n701 10.6151
R1295 B.n704 B.n702 10.6151
R1296 B.n705 B.n704 10.6151
R1297 B.n706 B.n705 10.6151
R1298 B.n804 B.n1 10.6151
R1299 B.n804 B.n803 10.6151
R1300 B.n803 B.n802 10.6151
R1301 B.n802 B.n10 10.6151
R1302 B.n796 B.n10 10.6151
R1303 B.n796 B.n795 10.6151
R1304 B.n795 B.n794 10.6151
R1305 B.n794 B.n18 10.6151
R1306 B.n788 B.n18 10.6151
R1307 B.n788 B.n787 10.6151
R1308 B.n787 B.n786 10.6151
R1309 B.n786 B.n25 10.6151
R1310 B.n780 B.n25 10.6151
R1311 B.n780 B.n779 10.6151
R1312 B.n779 B.n778 10.6151
R1313 B.n778 B.n32 10.6151
R1314 B.n772 B.n32 10.6151
R1315 B.n772 B.n771 10.6151
R1316 B.n771 B.n770 10.6151
R1317 B.n770 B.n39 10.6151
R1318 B.n764 B.n39 10.6151
R1319 B.n764 B.n763 10.6151
R1320 B.n763 B.n762 10.6151
R1321 B.n762 B.n46 10.6151
R1322 B.n756 B.n46 10.6151
R1323 B.n756 B.n755 10.6151
R1324 B.n755 B.n754 10.6151
R1325 B.n754 B.n53 10.6151
R1326 B.n748 B.n53 10.6151
R1327 B.n748 B.n747 10.6151
R1328 B.n747 B.n746 10.6151
R1329 B.n746 B.n59 10.6151
R1330 B.n740 B.n59 10.6151
R1331 B.n740 B.n739 10.6151
R1332 B.n739 B.n738 10.6151
R1333 B.n738 B.n67 10.6151
R1334 B.n732 B.n67 10.6151
R1335 B.n732 B.n731 10.6151
R1336 B.n731 B.n730 10.6151
R1337 B.n730 B.n74 10.6151
R1338 B.n724 B.n74 10.6151
R1339 B.n724 B.n723 10.6151
R1340 B.n723 B.n722 10.6151
R1341 B.n722 B.n81 10.6151
R1342 B.n716 B.n81 10.6151
R1343 B.n716 B.n715 10.6151
R1344 B.n715 B.n714 10.6151
R1345 B.n714 B.n88 10.6151
R1346 B.n128 B.n127 10.6151
R1347 B.n131 B.n128 10.6151
R1348 B.n132 B.n131 10.6151
R1349 B.n135 B.n132 10.6151
R1350 B.n136 B.n135 10.6151
R1351 B.n139 B.n136 10.6151
R1352 B.n140 B.n139 10.6151
R1353 B.n143 B.n140 10.6151
R1354 B.n144 B.n143 10.6151
R1355 B.n147 B.n144 10.6151
R1356 B.n148 B.n147 10.6151
R1357 B.n151 B.n148 10.6151
R1358 B.n152 B.n151 10.6151
R1359 B.n155 B.n152 10.6151
R1360 B.n156 B.n155 10.6151
R1361 B.n159 B.n156 10.6151
R1362 B.n160 B.n159 10.6151
R1363 B.n163 B.n160 10.6151
R1364 B.n164 B.n163 10.6151
R1365 B.n167 B.n164 10.6151
R1366 B.n168 B.n167 10.6151
R1367 B.n171 B.n168 10.6151
R1368 B.n172 B.n171 10.6151
R1369 B.n175 B.n172 10.6151
R1370 B.n180 B.n177 10.6151
R1371 B.n181 B.n180 10.6151
R1372 B.n184 B.n181 10.6151
R1373 B.n185 B.n184 10.6151
R1374 B.n188 B.n185 10.6151
R1375 B.n189 B.n188 10.6151
R1376 B.n192 B.n189 10.6151
R1377 B.n193 B.n192 10.6151
R1378 B.n196 B.n193 10.6151
R1379 B.n201 B.n198 10.6151
R1380 B.n202 B.n201 10.6151
R1381 B.n205 B.n202 10.6151
R1382 B.n206 B.n205 10.6151
R1383 B.n209 B.n206 10.6151
R1384 B.n210 B.n209 10.6151
R1385 B.n213 B.n210 10.6151
R1386 B.n214 B.n213 10.6151
R1387 B.n217 B.n214 10.6151
R1388 B.n218 B.n217 10.6151
R1389 B.n221 B.n218 10.6151
R1390 B.n222 B.n221 10.6151
R1391 B.n225 B.n222 10.6151
R1392 B.n226 B.n225 10.6151
R1393 B.n229 B.n226 10.6151
R1394 B.n230 B.n229 10.6151
R1395 B.n233 B.n230 10.6151
R1396 B.n234 B.n233 10.6151
R1397 B.n237 B.n234 10.6151
R1398 B.n238 B.n237 10.6151
R1399 B.n241 B.n238 10.6151
R1400 B.n243 B.n241 10.6151
R1401 B.n244 B.n243 10.6151
R1402 B.n707 B.n244 10.6151
R1403 B.n445 B.n374 9.36635
R1404 B.n422 B.n377 9.36635
R1405 B.n176 B.n175 9.36635
R1406 B.n198 B.n197 9.36635
R1407 B.n812 B.n0 8.11757
R1408 B.n812 B.n1 8.11757
R1409 B.n554 B.t5 1.89135
R1410 B.n750 B.t7 1.89135
R1411 B.n442 B.n374 1.24928
R1412 B.n425 B.n377 1.24928
R1413 B.n177 B.n176 1.24928
R1414 B.n197 B.n196 1.24928
R1415 VN.n51 VN.n27 161.3
R1416 VN.n50 VN.n49 161.3
R1417 VN.n48 VN.n28 161.3
R1418 VN.n47 VN.n46 161.3
R1419 VN.n45 VN.n29 161.3
R1420 VN.n44 VN.n43 161.3
R1421 VN.n42 VN.n41 161.3
R1422 VN.n40 VN.n31 161.3
R1423 VN.n39 VN.n38 161.3
R1424 VN.n37 VN.n32 161.3
R1425 VN.n36 VN.n35 161.3
R1426 VN.n24 VN.n0 161.3
R1427 VN.n23 VN.n22 161.3
R1428 VN.n21 VN.n1 161.3
R1429 VN.n20 VN.n19 161.3
R1430 VN.n18 VN.n2 161.3
R1431 VN.n17 VN.n16 161.3
R1432 VN.n15 VN.n14 161.3
R1433 VN.n13 VN.n4 161.3
R1434 VN.n12 VN.n11 161.3
R1435 VN.n10 VN.n5 161.3
R1436 VN.n9 VN.n8 161.3
R1437 VN.n26 VN.n25 100.334
R1438 VN.n53 VN.n52 100.334
R1439 VN.n6 VN.t0 95.6414
R1440 VN.n33 VN.t5 95.6414
R1441 VN.n7 VN.t4 61.8053
R1442 VN.n3 VN.t1 61.8053
R1443 VN.n25 VN.t7 61.8053
R1444 VN.n34 VN.t2 61.8053
R1445 VN.n30 VN.t6 61.8053
R1446 VN.n52 VN.t3 61.8053
R1447 VN.n19 VN.n1 56.5617
R1448 VN.n46 VN.n28 56.5617
R1449 VN.n7 VN.n6 52.7959
R1450 VN.n34 VN.n33 52.7959
R1451 VN VN.n53 46.3391
R1452 VN.n12 VN.n5 40.577
R1453 VN.n13 VN.n12 40.577
R1454 VN.n39 VN.n32 40.577
R1455 VN.n40 VN.n39 40.577
R1456 VN.n8 VN.n5 24.5923
R1457 VN.n14 VN.n13 24.5923
R1458 VN.n18 VN.n17 24.5923
R1459 VN.n19 VN.n18 24.5923
R1460 VN.n23 VN.n1 24.5923
R1461 VN.n24 VN.n23 24.5923
R1462 VN.n35 VN.n32 24.5923
R1463 VN.n46 VN.n45 24.5923
R1464 VN.n45 VN.n44 24.5923
R1465 VN.n41 VN.n40 24.5923
R1466 VN.n51 VN.n50 24.5923
R1467 VN.n50 VN.n28 24.5923
R1468 VN.n8 VN.n7 19.9199
R1469 VN.n14 VN.n3 19.9199
R1470 VN.n35 VN.n34 19.9199
R1471 VN.n41 VN.n30 19.9199
R1472 VN.n25 VN.n24 10.575
R1473 VN.n52 VN.n51 10.575
R1474 VN.n36 VN.n33 6.79754
R1475 VN.n9 VN.n6 6.79754
R1476 VN.n17 VN.n3 4.67295
R1477 VN.n44 VN.n30 4.67295
R1478 VN.n53 VN.n27 0.278335
R1479 VN.n26 VN.n0 0.278335
R1480 VN.n49 VN.n27 0.189894
R1481 VN.n49 VN.n48 0.189894
R1482 VN.n48 VN.n47 0.189894
R1483 VN.n47 VN.n29 0.189894
R1484 VN.n43 VN.n29 0.189894
R1485 VN.n43 VN.n42 0.189894
R1486 VN.n42 VN.n31 0.189894
R1487 VN.n38 VN.n31 0.189894
R1488 VN.n38 VN.n37 0.189894
R1489 VN.n37 VN.n36 0.189894
R1490 VN.n10 VN.n9 0.189894
R1491 VN.n11 VN.n10 0.189894
R1492 VN.n11 VN.n4 0.189894
R1493 VN.n15 VN.n4 0.189894
R1494 VN.n16 VN.n15 0.189894
R1495 VN.n16 VN.n2 0.189894
R1496 VN.n20 VN.n2 0.189894
R1497 VN.n21 VN.n20 0.189894
R1498 VN.n22 VN.n21 0.189894
R1499 VN.n22 VN.n0 0.189894
R1500 VN VN.n26 0.153485
R1501 VDD2.n2 VDD2.n1 67.7517
R1502 VDD2.n2 VDD2.n0 67.7517
R1503 VDD2 VDD2.n5 67.7489
R1504 VDD2.n4 VDD2.n3 66.5961
R1505 VDD2.n4 VDD2.n2 40.0989
R1506 VDD2.n5 VDD2.t2 3.11371
R1507 VDD2.n5 VDD2.t5 3.11371
R1508 VDD2.n3 VDD2.t1 3.11371
R1509 VDD2.n3 VDD2.t6 3.11371
R1510 VDD2.n1 VDD2.t0 3.11371
R1511 VDD2.n1 VDD2.t3 3.11371
R1512 VDD2.n0 VDD2.t7 3.11371
R1513 VDD2.n0 VDD2.t4 3.11371
R1514 VDD2 VDD2.n4 1.2699
R1515 VTAIL.n11 VTAIL.t2 53.0304
R1516 VTAIL.n10 VTAIL.t10 53.0304
R1517 VTAIL.n7 VTAIL.t12 53.0304
R1518 VTAIL.n15 VTAIL.t8 53.0303
R1519 VTAIL.n2 VTAIL.t15 53.0303
R1520 VTAIL.n3 VTAIL.t1 53.0303
R1521 VTAIL.n6 VTAIL.t6 53.0303
R1522 VTAIL.n14 VTAIL.t4 53.0303
R1523 VTAIL.n13 VTAIL.n12 49.9173
R1524 VTAIL.n9 VTAIL.n8 49.9173
R1525 VTAIL.n1 VTAIL.n0 49.917
R1526 VTAIL.n5 VTAIL.n4 49.917
R1527 VTAIL.n15 VTAIL.n14 20.2721
R1528 VTAIL.n7 VTAIL.n6 20.2721
R1529 VTAIL.n0 VTAIL.t11 3.11371
R1530 VTAIL.n0 VTAIL.t14 3.11371
R1531 VTAIL.n4 VTAIL.t3 3.11371
R1532 VTAIL.n4 VTAIL.t0 3.11371
R1533 VTAIL.n12 VTAIL.t7 3.11371
R1534 VTAIL.n12 VTAIL.t5 3.11371
R1535 VTAIL.n8 VTAIL.t9 3.11371
R1536 VTAIL.n8 VTAIL.t13 3.11371
R1537 VTAIL.n9 VTAIL.n7 2.42291
R1538 VTAIL.n10 VTAIL.n9 2.42291
R1539 VTAIL.n13 VTAIL.n11 2.42291
R1540 VTAIL.n14 VTAIL.n13 2.42291
R1541 VTAIL.n6 VTAIL.n5 2.42291
R1542 VTAIL.n5 VTAIL.n3 2.42291
R1543 VTAIL.n2 VTAIL.n1 2.42291
R1544 VTAIL VTAIL.n15 2.36472
R1545 VTAIL.n11 VTAIL.n10 0.470328
R1546 VTAIL.n3 VTAIL.n2 0.470328
R1547 VTAIL VTAIL.n1 0.0586897
R1548 VP.n19 VP.n18 161.3
R1549 VP.n20 VP.n15 161.3
R1550 VP.n22 VP.n21 161.3
R1551 VP.n23 VP.n14 161.3
R1552 VP.n25 VP.n24 161.3
R1553 VP.n27 VP.n26 161.3
R1554 VP.n28 VP.n12 161.3
R1555 VP.n30 VP.n29 161.3
R1556 VP.n31 VP.n11 161.3
R1557 VP.n33 VP.n32 161.3
R1558 VP.n34 VP.n10 161.3
R1559 VP.n64 VP.n0 161.3
R1560 VP.n63 VP.n62 161.3
R1561 VP.n61 VP.n1 161.3
R1562 VP.n60 VP.n59 161.3
R1563 VP.n58 VP.n2 161.3
R1564 VP.n57 VP.n56 161.3
R1565 VP.n55 VP.n54 161.3
R1566 VP.n53 VP.n4 161.3
R1567 VP.n52 VP.n51 161.3
R1568 VP.n50 VP.n5 161.3
R1569 VP.n49 VP.n48 161.3
R1570 VP.n46 VP.n6 161.3
R1571 VP.n45 VP.n44 161.3
R1572 VP.n43 VP.n7 161.3
R1573 VP.n42 VP.n41 161.3
R1574 VP.n40 VP.n8 161.3
R1575 VP.n39 VP.n38 161.3
R1576 VP.n37 VP.n9 100.334
R1577 VP.n66 VP.n65 100.334
R1578 VP.n36 VP.n35 100.334
R1579 VP.n16 VP.t1 95.6414
R1580 VP.n9 VP.t5 61.8053
R1581 VP.n47 VP.t7 61.8053
R1582 VP.n3 VP.t4 61.8053
R1583 VP.n65 VP.t6 61.8053
R1584 VP.n35 VP.t2 61.8053
R1585 VP.n13 VP.t0 61.8053
R1586 VP.n17 VP.t3 61.8053
R1587 VP.n41 VP.n7 56.5617
R1588 VP.n59 VP.n1 56.5617
R1589 VP.n29 VP.n11 56.5617
R1590 VP.n17 VP.n16 52.7959
R1591 VP.n37 VP.n36 46.0603
R1592 VP.n52 VP.n5 40.577
R1593 VP.n53 VP.n52 40.577
R1594 VP.n23 VP.n22 40.577
R1595 VP.n22 VP.n15 40.577
R1596 VP.n40 VP.n39 24.5923
R1597 VP.n41 VP.n40 24.5923
R1598 VP.n45 VP.n7 24.5923
R1599 VP.n46 VP.n45 24.5923
R1600 VP.n48 VP.n5 24.5923
R1601 VP.n54 VP.n53 24.5923
R1602 VP.n58 VP.n57 24.5923
R1603 VP.n59 VP.n58 24.5923
R1604 VP.n63 VP.n1 24.5923
R1605 VP.n64 VP.n63 24.5923
R1606 VP.n33 VP.n11 24.5923
R1607 VP.n34 VP.n33 24.5923
R1608 VP.n24 VP.n23 24.5923
R1609 VP.n28 VP.n27 24.5923
R1610 VP.n29 VP.n28 24.5923
R1611 VP.n18 VP.n15 24.5923
R1612 VP.n48 VP.n47 19.9199
R1613 VP.n54 VP.n3 19.9199
R1614 VP.n24 VP.n13 19.9199
R1615 VP.n18 VP.n17 19.9199
R1616 VP.n39 VP.n9 10.575
R1617 VP.n65 VP.n64 10.575
R1618 VP.n35 VP.n34 10.575
R1619 VP.n19 VP.n16 6.79754
R1620 VP.n47 VP.n46 4.67295
R1621 VP.n57 VP.n3 4.67295
R1622 VP.n27 VP.n13 4.67295
R1623 VP.n36 VP.n10 0.278335
R1624 VP.n38 VP.n37 0.278335
R1625 VP.n66 VP.n0 0.278335
R1626 VP.n20 VP.n19 0.189894
R1627 VP.n21 VP.n20 0.189894
R1628 VP.n21 VP.n14 0.189894
R1629 VP.n25 VP.n14 0.189894
R1630 VP.n26 VP.n25 0.189894
R1631 VP.n26 VP.n12 0.189894
R1632 VP.n30 VP.n12 0.189894
R1633 VP.n31 VP.n30 0.189894
R1634 VP.n32 VP.n31 0.189894
R1635 VP.n32 VP.n10 0.189894
R1636 VP.n38 VP.n8 0.189894
R1637 VP.n42 VP.n8 0.189894
R1638 VP.n43 VP.n42 0.189894
R1639 VP.n44 VP.n43 0.189894
R1640 VP.n44 VP.n6 0.189894
R1641 VP.n49 VP.n6 0.189894
R1642 VP.n50 VP.n49 0.189894
R1643 VP.n51 VP.n50 0.189894
R1644 VP.n51 VP.n4 0.189894
R1645 VP.n55 VP.n4 0.189894
R1646 VP.n56 VP.n55 0.189894
R1647 VP.n56 VP.n2 0.189894
R1648 VP.n60 VP.n2 0.189894
R1649 VP.n61 VP.n60 0.189894
R1650 VP.n62 VP.n61 0.189894
R1651 VP.n62 VP.n0 0.189894
R1652 VP VP.n66 0.153485
R1653 VDD1 VDD1.n0 67.8654
R1654 VDD1.n3 VDD1.n2 67.7517
R1655 VDD1.n3 VDD1.n1 67.7517
R1656 VDD1.n5 VDD1.n4 66.5959
R1657 VDD1.n5 VDD1.n3 40.6819
R1658 VDD1.n4 VDD1.t7 3.11371
R1659 VDD1.n4 VDD1.t5 3.11371
R1660 VDD1.n0 VDD1.t6 3.11371
R1661 VDD1.n0 VDD1.t4 3.11371
R1662 VDD1.n2 VDD1.t3 3.11371
R1663 VDD1.n2 VDD1.t1 3.11371
R1664 VDD1.n1 VDD1.t2 3.11371
R1665 VDD1.n1 VDD1.t0 3.11371
R1666 VDD1 VDD1.n5 1.15352
C0 VP VDD2 0.507336f
C1 VN VDD2 4.77167f
C2 VTAIL VDD1 6.11368f
C3 VP VN 6.46601f
C4 VDD2 VDD1 1.71564f
C5 VP VDD1 5.12573f
C6 VN VDD1 0.151945f
C7 VTAIL VDD2 6.16729f
C8 VP VTAIL 5.56129f
C9 VN VTAIL 5.54718f
C10 VDD2 B 4.795033f
C11 VDD1 B 5.217693f
C12 VTAIL B 6.669565f
C13 VN B 14.430301f
C14 VP B 13.049212f
C15 VDD1.t6 B 0.123859f
C16 VDD1.t4 B 0.123859f
C17 VDD1.n0 B 1.04956f
C18 VDD1.t2 B 0.123859f
C19 VDD1.t0 B 0.123859f
C20 VDD1.n1 B 1.04858f
C21 VDD1.t3 B 0.123859f
C22 VDD1.t1 B 0.123859f
C23 VDD1.n2 B 1.04858f
C24 VDD1.n3 B 2.86942f
C25 VDD1.t7 B 0.123859f
C26 VDD1.t5 B 0.123859f
C27 VDD1.n4 B 1.04012f
C28 VDD1.n5 B 2.46574f
C29 VP.n0 B 0.034072f
C30 VP.t6 B 1.08254f
C31 VP.n1 B 0.033279f
C32 VP.n2 B 0.025845f
C33 VP.t4 B 1.08254f
C34 VP.n3 B 0.404464f
C35 VP.n4 B 0.025845f
C36 VP.n5 B 0.051096f
C37 VP.n6 B 0.025845f
C38 VP.t7 B 1.08254f
C39 VP.n7 B 0.04186f
C40 VP.n8 B 0.025845f
C41 VP.t5 B 1.08254f
C42 VP.n9 B 0.487202f
C43 VP.n10 B 0.034072f
C44 VP.t2 B 1.08254f
C45 VP.n11 B 0.033279f
C46 VP.n12 B 0.025845f
C47 VP.t0 B 1.08254f
C48 VP.n13 B 0.404464f
C49 VP.n14 B 0.025845f
C50 VP.n15 B 0.051096f
C51 VP.t1 B 1.28026f
C52 VP.n16 B 0.45829f
C53 VP.t3 B 1.08254f
C54 VP.n17 B 0.484659f
C55 VP.n18 B 0.043431f
C56 VP.n19 B 0.246673f
C57 VP.n20 B 0.025845f
C58 VP.n21 B 0.025845f
C59 VP.n22 B 0.020874f
C60 VP.n23 B 0.051096f
C61 VP.n24 B 0.043431f
C62 VP.n25 B 0.025845f
C63 VP.n26 B 0.025845f
C64 VP.n27 B 0.028762f
C65 VP.n28 B 0.047927f
C66 VP.n29 B 0.04186f
C67 VP.n30 B 0.025845f
C68 VP.n31 B 0.025845f
C69 VP.n32 B 0.025845f
C70 VP.n33 B 0.047927f
C71 VP.n34 B 0.03444f
C72 VP.n35 B 0.487202f
C73 VP.n36 B 1.26993f
C74 VP.n37 B 1.29016f
C75 VP.n38 B 0.034072f
C76 VP.n39 B 0.03444f
C77 VP.n40 B 0.047927f
C78 VP.n41 B 0.033279f
C79 VP.n42 B 0.025845f
C80 VP.n43 B 0.025845f
C81 VP.n44 B 0.025845f
C82 VP.n45 B 0.047927f
C83 VP.n46 B 0.028762f
C84 VP.n47 B 0.404464f
C85 VP.n48 B 0.043431f
C86 VP.n49 B 0.025845f
C87 VP.n50 B 0.025845f
C88 VP.n51 B 0.025845f
C89 VP.n52 B 0.020874f
C90 VP.n53 B 0.051096f
C91 VP.n54 B 0.043431f
C92 VP.n55 B 0.025845f
C93 VP.n56 B 0.025845f
C94 VP.n57 B 0.028762f
C95 VP.n58 B 0.047927f
C96 VP.n59 B 0.04186f
C97 VP.n60 B 0.025845f
C98 VP.n61 B 0.025845f
C99 VP.n62 B 0.025845f
C100 VP.n63 B 0.047927f
C101 VP.n64 B 0.03444f
C102 VP.n65 B 0.487202f
C103 VP.n66 B 0.040726f
C104 VTAIL.t11 B 0.114724f
C105 VTAIL.t14 B 0.114724f
C106 VTAIL.n0 B 0.902622f
C107 VTAIL.n1 B 0.398503f
C108 VTAIL.t15 B 1.15088f
C109 VTAIL.n2 B 0.493405f
C110 VTAIL.t1 B 1.15088f
C111 VTAIL.n3 B 0.493405f
C112 VTAIL.t3 B 0.114724f
C113 VTAIL.t0 B 0.114724f
C114 VTAIL.n4 B 0.902622f
C115 VTAIL.n5 B 0.572398f
C116 VTAIL.t6 B 1.15088f
C117 VTAIL.n6 B 1.35037f
C118 VTAIL.t12 B 1.15089f
C119 VTAIL.n7 B 1.35036f
C120 VTAIL.t9 B 0.114724f
C121 VTAIL.t13 B 0.114724f
C122 VTAIL.n8 B 0.902627f
C123 VTAIL.n9 B 0.572393f
C124 VTAIL.t10 B 1.15089f
C125 VTAIL.n10 B 0.493398f
C126 VTAIL.t2 B 1.15089f
C127 VTAIL.n11 B 0.493398f
C128 VTAIL.t7 B 0.114724f
C129 VTAIL.t5 B 0.114724f
C130 VTAIL.n12 B 0.902627f
C131 VTAIL.n13 B 0.572393f
C132 VTAIL.t4 B 1.15088f
C133 VTAIL.n14 B 1.35037f
C134 VTAIL.t8 B 1.15088f
C135 VTAIL.n15 B 1.34609f
C136 VDD2.t7 B 0.122643f
C137 VDD2.t4 B 0.122643f
C138 VDD2.n0 B 1.03829f
C139 VDD2.t0 B 0.122643f
C140 VDD2.t3 B 0.122643f
C141 VDD2.n1 B 1.03829f
C142 VDD2.n2 B 2.7902f
C143 VDD2.t1 B 0.122643f
C144 VDD2.t6 B 0.122643f
C145 VDD2.n3 B 1.02993f
C146 VDD2.n4 B 2.41163f
C147 VDD2.t2 B 0.122643f
C148 VDD2.t5 B 0.122643f
C149 VDD2.n5 B 1.03826f
C150 VN.n0 B 0.033209f
C151 VN.t7 B 1.05513f
C152 VN.n1 B 0.032437f
C153 VN.n2 B 0.025191f
C154 VN.t1 B 1.05513f
C155 VN.n3 B 0.394225f
C156 VN.n4 B 0.025191f
C157 VN.n5 B 0.049802f
C158 VN.t0 B 1.24785f
C159 VN.n6 B 0.446688f
C160 VN.t4 B 1.05513f
C161 VN.n7 B 0.47239f
C162 VN.n8 B 0.042332f
C163 VN.n9 B 0.240429f
C164 VN.n10 B 0.025191f
C165 VN.n11 B 0.025191f
C166 VN.n12 B 0.020346f
C167 VN.n13 B 0.049802f
C168 VN.n14 B 0.042332f
C169 VN.n15 B 0.025191f
C170 VN.n16 B 0.025191f
C171 VN.n17 B 0.028034f
C172 VN.n18 B 0.046714f
C173 VN.n19 B 0.0408f
C174 VN.n20 B 0.025191f
C175 VN.n21 B 0.025191f
C176 VN.n22 B 0.025191f
C177 VN.n23 B 0.046714f
C178 VN.n24 B 0.033569f
C179 VN.n25 B 0.474869f
C180 VN.n26 B 0.039695f
C181 VN.n27 B 0.033209f
C182 VN.t3 B 1.05513f
C183 VN.n28 B 0.032437f
C184 VN.n29 B 0.025191f
C185 VN.t6 B 1.05513f
C186 VN.n30 B 0.394225f
C187 VN.n31 B 0.025191f
C188 VN.n32 B 0.049802f
C189 VN.t5 B 1.24785f
C190 VN.n33 B 0.446688f
C191 VN.t2 B 1.05513f
C192 VN.n34 B 0.47239f
C193 VN.n35 B 0.042332f
C194 VN.n36 B 0.240429f
C195 VN.n37 B 0.025191f
C196 VN.n38 B 0.025191f
C197 VN.n39 B 0.020346f
C198 VN.n40 B 0.049802f
C199 VN.n41 B 0.042332f
C200 VN.n42 B 0.025191f
C201 VN.n43 B 0.025191f
C202 VN.n44 B 0.028034f
C203 VN.n45 B 0.046714f
C204 VN.n46 B 0.0408f
C205 VN.n47 B 0.025191f
C206 VN.n48 B 0.025191f
C207 VN.n49 B 0.025191f
C208 VN.n50 B 0.046714f
C209 VN.n51 B 0.033569f
C210 VN.n52 B 0.474869f
C211 VN.n53 B 1.2515f
.ends

