* NGSPICE file created from diff_pair_sample_0498.ext - technology: sky130A

.subckt diff_pair_sample_0498 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=6.0801 ps=31.96 w=15.59 l=3.4
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=0 ps=0 w=15.59 l=3.4
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=6.0801 ps=31.96 w=15.59 l=3.4
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=0 ps=0 w=15.59 l=3.4
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=6.0801 ps=31.96 w=15.59 l=3.4
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=0 ps=0 w=15.59 l=3.4
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=0 ps=0 w=15.59 l=3.4
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.0801 pd=31.96 as=6.0801 ps=31.96 w=15.59 l=3.4
R0 VP.n0 VP.t1 198.792
R1 VP.n0 VP.t0 149.293
R2 VP VP.n0 0.52637
R3 VTAIL.n338 VTAIL.n258 289.615
R4 VTAIL.n80 VTAIL.n0 289.615
R5 VTAIL.n252 VTAIL.n172 289.615
R6 VTAIL.n166 VTAIL.n86 289.615
R7 VTAIL.n287 VTAIL.n286 185
R8 VTAIL.n289 VTAIL.n288 185
R9 VTAIL.n282 VTAIL.n281 185
R10 VTAIL.n295 VTAIL.n294 185
R11 VTAIL.n297 VTAIL.n296 185
R12 VTAIL.n278 VTAIL.n277 185
R13 VTAIL.n303 VTAIL.n302 185
R14 VTAIL.n305 VTAIL.n304 185
R15 VTAIL.n274 VTAIL.n273 185
R16 VTAIL.n311 VTAIL.n310 185
R17 VTAIL.n313 VTAIL.n312 185
R18 VTAIL.n270 VTAIL.n269 185
R19 VTAIL.n319 VTAIL.n318 185
R20 VTAIL.n321 VTAIL.n320 185
R21 VTAIL.n266 VTAIL.n265 185
R22 VTAIL.n328 VTAIL.n327 185
R23 VTAIL.n329 VTAIL.n264 185
R24 VTAIL.n331 VTAIL.n330 185
R25 VTAIL.n262 VTAIL.n261 185
R26 VTAIL.n337 VTAIL.n336 185
R27 VTAIL.n339 VTAIL.n338 185
R28 VTAIL.n29 VTAIL.n28 185
R29 VTAIL.n31 VTAIL.n30 185
R30 VTAIL.n24 VTAIL.n23 185
R31 VTAIL.n37 VTAIL.n36 185
R32 VTAIL.n39 VTAIL.n38 185
R33 VTAIL.n20 VTAIL.n19 185
R34 VTAIL.n45 VTAIL.n44 185
R35 VTAIL.n47 VTAIL.n46 185
R36 VTAIL.n16 VTAIL.n15 185
R37 VTAIL.n53 VTAIL.n52 185
R38 VTAIL.n55 VTAIL.n54 185
R39 VTAIL.n12 VTAIL.n11 185
R40 VTAIL.n61 VTAIL.n60 185
R41 VTAIL.n63 VTAIL.n62 185
R42 VTAIL.n8 VTAIL.n7 185
R43 VTAIL.n70 VTAIL.n69 185
R44 VTAIL.n71 VTAIL.n6 185
R45 VTAIL.n73 VTAIL.n72 185
R46 VTAIL.n4 VTAIL.n3 185
R47 VTAIL.n79 VTAIL.n78 185
R48 VTAIL.n81 VTAIL.n80 185
R49 VTAIL.n253 VTAIL.n252 185
R50 VTAIL.n251 VTAIL.n250 185
R51 VTAIL.n176 VTAIL.n175 185
R52 VTAIL.n180 VTAIL.n178 185
R53 VTAIL.n245 VTAIL.n244 185
R54 VTAIL.n243 VTAIL.n242 185
R55 VTAIL.n182 VTAIL.n181 185
R56 VTAIL.n237 VTAIL.n236 185
R57 VTAIL.n235 VTAIL.n234 185
R58 VTAIL.n186 VTAIL.n185 185
R59 VTAIL.n229 VTAIL.n228 185
R60 VTAIL.n227 VTAIL.n226 185
R61 VTAIL.n190 VTAIL.n189 185
R62 VTAIL.n221 VTAIL.n220 185
R63 VTAIL.n219 VTAIL.n218 185
R64 VTAIL.n194 VTAIL.n193 185
R65 VTAIL.n213 VTAIL.n212 185
R66 VTAIL.n211 VTAIL.n210 185
R67 VTAIL.n198 VTAIL.n197 185
R68 VTAIL.n205 VTAIL.n204 185
R69 VTAIL.n203 VTAIL.n202 185
R70 VTAIL.n167 VTAIL.n166 185
R71 VTAIL.n165 VTAIL.n164 185
R72 VTAIL.n90 VTAIL.n89 185
R73 VTAIL.n94 VTAIL.n92 185
R74 VTAIL.n159 VTAIL.n158 185
R75 VTAIL.n157 VTAIL.n156 185
R76 VTAIL.n96 VTAIL.n95 185
R77 VTAIL.n151 VTAIL.n150 185
R78 VTAIL.n149 VTAIL.n148 185
R79 VTAIL.n100 VTAIL.n99 185
R80 VTAIL.n143 VTAIL.n142 185
R81 VTAIL.n141 VTAIL.n140 185
R82 VTAIL.n104 VTAIL.n103 185
R83 VTAIL.n135 VTAIL.n134 185
R84 VTAIL.n133 VTAIL.n132 185
R85 VTAIL.n108 VTAIL.n107 185
R86 VTAIL.n127 VTAIL.n126 185
R87 VTAIL.n125 VTAIL.n124 185
R88 VTAIL.n112 VTAIL.n111 185
R89 VTAIL.n119 VTAIL.n118 185
R90 VTAIL.n117 VTAIL.n116 185
R91 VTAIL.n285 VTAIL.t0 147.659
R92 VTAIL.n27 VTAIL.t3 147.659
R93 VTAIL.n201 VTAIL.t2 147.659
R94 VTAIL.n115 VTAIL.t1 147.659
R95 VTAIL.n288 VTAIL.n287 104.615
R96 VTAIL.n288 VTAIL.n281 104.615
R97 VTAIL.n295 VTAIL.n281 104.615
R98 VTAIL.n296 VTAIL.n295 104.615
R99 VTAIL.n296 VTAIL.n277 104.615
R100 VTAIL.n303 VTAIL.n277 104.615
R101 VTAIL.n304 VTAIL.n303 104.615
R102 VTAIL.n304 VTAIL.n273 104.615
R103 VTAIL.n311 VTAIL.n273 104.615
R104 VTAIL.n312 VTAIL.n311 104.615
R105 VTAIL.n312 VTAIL.n269 104.615
R106 VTAIL.n319 VTAIL.n269 104.615
R107 VTAIL.n320 VTAIL.n319 104.615
R108 VTAIL.n320 VTAIL.n265 104.615
R109 VTAIL.n328 VTAIL.n265 104.615
R110 VTAIL.n329 VTAIL.n328 104.615
R111 VTAIL.n330 VTAIL.n329 104.615
R112 VTAIL.n330 VTAIL.n261 104.615
R113 VTAIL.n337 VTAIL.n261 104.615
R114 VTAIL.n338 VTAIL.n337 104.615
R115 VTAIL.n30 VTAIL.n29 104.615
R116 VTAIL.n30 VTAIL.n23 104.615
R117 VTAIL.n37 VTAIL.n23 104.615
R118 VTAIL.n38 VTAIL.n37 104.615
R119 VTAIL.n38 VTAIL.n19 104.615
R120 VTAIL.n45 VTAIL.n19 104.615
R121 VTAIL.n46 VTAIL.n45 104.615
R122 VTAIL.n46 VTAIL.n15 104.615
R123 VTAIL.n53 VTAIL.n15 104.615
R124 VTAIL.n54 VTAIL.n53 104.615
R125 VTAIL.n54 VTAIL.n11 104.615
R126 VTAIL.n61 VTAIL.n11 104.615
R127 VTAIL.n62 VTAIL.n61 104.615
R128 VTAIL.n62 VTAIL.n7 104.615
R129 VTAIL.n70 VTAIL.n7 104.615
R130 VTAIL.n71 VTAIL.n70 104.615
R131 VTAIL.n72 VTAIL.n71 104.615
R132 VTAIL.n72 VTAIL.n3 104.615
R133 VTAIL.n79 VTAIL.n3 104.615
R134 VTAIL.n80 VTAIL.n79 104.615
R135 VTAIL.n252 VTAIL.n251 104.615
R136 VTAIL.n251 VTAIL.n175 104.615
R137 VTAIL.n180 VTAIL.n175 104.615
R138 VTAIL.n244 VTAIL.n180 104.615
R139 VTAIL.n244 VTAIL.n243 104.615
R140 VTAIL.n243 VTAIL.n181 104.615
R141 VTAIL.n236 VTAIL.n181 104.615
R142 VTAIL.n236 VTAIL.n235 104.615
R143 VTAIL.n235 VTAIL.n185 104.615
R144 VTAIL.n228 VTAIL.n185 104.615
R145 VTAIL.n228 VTAIL.n227 104.615
R146 VTAIL.n227 VTAIL.n189 104.615
R147 VTAIL.n220 VTAIL.n189 104.615
R148 VTAIL.n220 VTAIL.n219 104.615
R149 VTAIL.n219 VTAIL.n193 104.615
R150 VTAIL.n212 VTAIL.n193 104.615
R151 VTAIL.n212 VTAIL.n211 104.615
R152 VTAIL.n211 VTAIL.n197 104.615
R153 VTAIL.n204 VTAIL.n197 104.615
R154 VTAIL.n204 VTAIL.n203 104.615
R155 VTAIL.n166 VTAIL.n165 104.615
R156 VTAIL.n165 VTAIL.n89 104.615
R157 VTAIL.n94 VTAIL.n89 104.615
R158 VTAIL.n158 VTAIL.n94 104.615
R159 VTAIL.n158 VTAIL.n157 104.615
R160 VTAIL.n157 VTAIL.n95 104.615
R161 VTAIL.n150 VTAIL.n95 104.615
R162 VTAIL.n150 VTAIL.n149 104.615
R163 VTAIL.n149 VTAIL.n99 104.615
R164 VTAIL.n142 VTAIL.n99 104.615
R165 VTAIL.n142 VTAIL.n141 104.615
R166 VTAIL.n141 VTAIL.n103 104.615
R167 VTAIL.n134 VTAIL.n103 104.615
R168 VTAIL.n134 VTAIL.n133 104.615
R169 VTAIL.n133 VTAIL.n107 104.615
R170 VTAIL.n126 VTAIL.n107 104.615
R171 VTAIL.n126 VTAIL.n125 104.615
R172 VTAIL.n125 VTAIL.n111 104.615
R173 VTAIL.n118 VTAIL.n111 104.615
R174 VTAIL.n118 VTAIL.n117 104.615
R175 VTAIL.n287 VTAIL.t0 52.3082
R176 VTAIL.n29 VTAIL.t3 52.3082
R177 VTAIL.n203 VTAIL.t2 52.3082
R178 VTAIL.n117 VTAIL.t1 52.3082
R179 VTAIL.n343 VTAIL.n342 36.646
R180 VTAIL.n85 VTAIL.n84 36.646
R181 VTAIL.n257 VTAIL.n256 36.646
R182 VTAIL.n171 VTAIL.n170 36.646
R183 VTAIL.n171 VTAIL.n85 32.2376
R184 VTAIL.n343 VTAIL.n257 29.0221
R185 VTAIL.n286 VTAIL.n285 15.6677
R186 VTAIL.n28 VTAIL.n27 15.6677
R187 VTAIL.n202 VTAIL.n201 15.6677
R188 VTAIL.n116 VTAIL.n115 15.6677
R189 VTAIL.n331 VTAIL.n262 13.1884
R190 VTAIL.n73 VTAIL.n4 13.1884
R191 VTAIL.n178 VTAIL.n176 13.1884
R192 VTAIL.n92 VTAIL.n90 13.1884
R193 VTAIL.n289 VTAIL.n284 12.8005
R194 VTAIL.n332 VTAIL.n264 12.8005
R195 VTAIL.n336 VTAIL.n335 12.8005
R196 VTAIL.n31 VTAIL.n26 12.8005
R197 VTAIL.n74 VTAIL.n6 12.8005
R198 VTAIL.n78 VTAIL.n77 12.8005
R199 VTAIL.n250 VTAIL.n249 12.8005
R200 VTAIL.n246 VTAIL.n245 12.8005
R201 VTAIL.n205 VTAIL.n200 12.8005
R202 VTAIL.n164 VTAIL.n163 12.8005
R203 VTAIL.n160 VTAIL.n159 12.8005
R204 VTAIL.n119 VTAIL.n114 12.8005
R205 VTAIL.n290 VTAIL.n282 12.0247
R206 VTAIL.n327 VTAIL.n326 12.0247
R207 VTAIL.n339 VTAIL.n260 12.0247
R208 VTAIL.n32 VTAIL.n24 12.0247
R209 VTAIL.n69 VTAIL.n68 12.0247
R210 VTAIL.n81 VTAIL.n2 12.0247
R211 VTAIL.n253 VTAIL.n174 12.0247
R212 VTAIL.n242 VTAIL.n179 12.0247
R213 VTAIL.n206 VTAIL.n198 12.0247
R214 VTAIL.n167 VTAIL.n88 12.0247
R215 VTAIL.n156 VTAIL.n93 12.0247
R216 VTAIL.n120 VTAIL.n112 12.0247
R217 VTAIL.n294 VTAIL.n293 11.249
R218 VTAIL.n325 VTAIL.n266 11.249
R219 VTAIL.n340 VTAIL.n258 11.249
R220 VTAIL.n36 VTAIL.n35 11.249
R221 VTAIL.n67 VTAIL.n8 11.249
R222 VTAIL.n82 VTAIL.n0 11.249
R223 VTAIL.n254 VTAIL.n172 11.249
R224 VTAIL.n241 VTAIL.n182 11.249
R225 VTAIL.n210 VTAIL.n209 11.249
R226 VTAIL.n168 VTAIL.n86 11.249
R227 VTAIL.n155 VTAIL.n96 11.249
R228 VTAIL.n124 VTAIL.n123 11.249
R229 VTAIL.n297 VTAIL.n280 10.4732
R230 VTAIL.n322 VTAIL.n321 10.4732
R231 VTAIL.n39 VTAIL.n22 10.4732
R232 VTAIL.n64 VTAIL.n63 10.4732
R233 VTAIL.n238 VTAIL.n237 10.4732
R234 VTAIL.n213 VTAIL.n196 10.4732
R235 VTAIL.n152 VTAIL.n151 10.4732
R236 VTAIL.n127 VTAIL.n110 10.4732
R237 VTAIL.n298 VTAIL.n278 9.69747
R238 VTAIL.n318 VTAIL.n268 9.69747
R239 VTAIL.n40 VTAIL.n20 9.69747
R240 VTAIL.n60 VTAIL.n10 9.69747
R241 VTAIL.n234 VTAIL.n184 9.69747
R242 VTAIL.n214 VTAIL.n194 9.69747
R243 VTAIL.n148 VTAIL.n98 9.69747
R244 VTAIL.n128 VTAIL.n108 9.69747
R245 VTAIL.n342 VTAIL.n341 9.45567
R246 VTAIL.n84 VTAIL.n83 9.45567
R247 VTAIL.n256 VTAIL.n255 9.45567
R248 VTAIL.n170 VTAIL.n169 9.45567
R249 VTAIL.n341 VTAIL.n340 9.3005
R250 VTAIL.n260 VTAIL.n259 9.3005
R251 VTAIL.n335 VTAIL.n334 9.3005
R252 VTAIL.n307 VTAIL.n306 9.3005
R253 VTAIL.n276 VTAIL.n275 9.3005
R254 VTAIL.n301 VTAIL.n300 9.3005
R255 VTAIL.n299 VTAIL.n298 9.3005
R256 VTAIL.n280 VTAIL.n279 9.3005
R257 VTAIL.n293 VTAIL.n292 9.3005
R258 VTAIL.n291 VTAIL.n290 9.3005
R259 VTAIL.n284 VTAIL.n283 9.3005
R260 VTAIL.n309 VTAIL.n308 9.3005
R261 VTAIL.n272 VTAIL.n271 9.3005
R262 VTAIL.n315 VTAIL.n314 9.3005
R263 VTAIL.n317 VTAIL.n316 9.3005
R264 VTAIL.n268 VTAIL.n267 9.3005
R265 VTAIL.n323 VTAIL.n322 9.3005
R266 VTAIL.n325 VTAIL.n324 9.3005
R267 VTAIL.n326 VTAIL.n263 9.3005
R268 VTAIL.n333 VTAIL.n332 9.3005
R269 VTAIL.n83 VTAIL.n82 9.3005
R270 VTAIL.n2 VTAIL.n1 9.3005
R271 VTAIL.n77 VTAIL.n76 9.3005
R272 VTAIL.n49 VTAIL.n48 9.3005
R273 VTAIL.n18 VTAIL.n17 9.3005
R274 VTAIL.n43 VTAIL.n42 9.3005
R275 VTAIL.n41 VTAIL.n40 9.3005
R276 VTAIL.n22 VTAIL.n21 9.3005
R277 VTAIL.n35 VTAIL.n34 9.3005
R278 VTAIL.n33 VTAIL.n32 9.3005
R279 VTAIL.n26 VTAIL.n25 9.3005
R280 VTAIL.n51 VTAIL.n50 9.3005
R281 VTAIL.n14 VTAIL.n13 9.3005
R282 VTAIL.n57 VTAIL.n56 9.3005
R283 VTAIL.n59 VTAIL.n58 9.3005
R284 VTAIL.n10 VTAIL.n9 9.3005
R285 VTAIL.n65 VTAIL.n64 9.3005
R286 VTAIL.n67 VTAIL.n66 9.3005
R287 VTAIL.n68 VTAIL.n5 9.3005
R288 VTAIL.n75 VTAIL.n74 9.3005
R289 VTAIL.n188 VTAIL.n187 9.3005
R290 VTAIL.n231 VTAIL.n230 9.3005
R291 VTAIL.n233 VTAIL.n232 9.3005
R292 VTAIL.n184 VTAIL.n183 9.3005
R293 VTAIL.n239 VTAIL.n238 9.3005
R294 VTAIL.n241 VTAIL.n240 9.3005
R295 VTAIL.n179 VTAIL.n177 9.3005
R296 VTAIL.n247 VTAIL.n246 9.3005
R297 VTAIL.n255 VTAIL.n254 9.3005
R298 VTAIL.n174 VTAIL.n173 9.3005
R299 VTAIL.n249 VTAIL.n248 9.3005
R300 VTAIL.n225 VTAIL.n224 9.3005
R301 VTAIL.n223 VTAIL.n222 9.3005
R302 VTAIL.n192 VTAIL.n191 9.3005
R303 VTAIL.n217 VTAIL.n216 9.3005
R304 VTAIL.n215 VTAIL.n214 9.3005
R305 VTAIL.n196 VTAIL.n195 9.3005
R306 VTAIL.n209 VTAIL.n208 9.3005
R307 VTAIL.n207 VTAIL.n206 9.3005
R308 VTAIL.n200 VTAIL.n199 9.3005
R309 VTAIL.n102 VTAIL.n101 9.3005
R310 VTAIL.n145 VTAIL.n144 9.3005
R311 VTAIL.n147 VTAIL.n146 9.3005
R312 VTAIL.n98 VTAIL.n97 9.3005
R313 VTAIL.n153 VTAIL.n152 9.3005
R314 VTAIL.n155 VTAIL.n154 9.3005
R315 VTAIL.n93 VTAIL.n91 9.3005
R316 VTAIL.n161 VTAIL.n160 9.3005
R317 VTAIL.n169 VTAIL.n168 9.3005
R318 VTAIL.n88 VTAIL.n87 9.3005
R319 VTAIL.n163 VTAIL.n162 9.3005
R320 VTAIL.n139 VTAIL.n138 9.3005
R321 VTAIL.n137 VTAIL.n136 9.3005
R322 VTAIL.n106 VTAIL.n105 9.3005
R323 VTAIL.n131 VTAIL.n130 9.3005
R324 VTAIL.n129 VTAIL.n128 9.3005
R325 VTAIL.n110 VTAIL.n109 9.3005
R326 VTAIL.n123 VTAIL.n122 9.3005
R327 VTAIL.n121 VTAIL.n120 9.3005
R328 VTAIL.n114 VTAIL.n113 9.3005
R329 VTAIL.n302 VTAIL.n301 8.92171
R330 VTAIL.n317 VTAIL.n270 8.92171
R331 VTAIL.n44 VTAIL.n43 8.92171
R332 VTAIL.n59 VTAIL.n12 8.92171
R333 VTAIL.n233 VTAIL.n186 8.92171
R334 VTAIL.n218 VTAIL.n217 8.92171
R335 VTAIL.n147 VTAIL.n100 8.92171
R336 VTAIL.n132 VTAIL.n131 8.92171
R337 VTAIL.n305 VTAIL.n276 8.14595
R338 VTAIL.n314 VTAIL.n313 8.14595
R339 VTAIL.n47 VTAIL.n18 8.14595
R340 VTAIL.n56 VTAIL.n55 8.14595
R341 VTAIL.n230 VTAIL.n229 8.14595
R342 VTAIL.n221 VTAIL.n192 8.14595
R343 VTAIL.n144 VTAIL.n143 8.14595
R344 VTAIL.n135 VTAIL.n106 8.14595
R345 VTAIL.n306 VTAIL.n274 7.3702
R346 VTAIL.n310 VTAIL.n272 7.3702
R347 VTAIL.n48 VTAIL.n16 7.3702
R348 VTAIL.n52 VTAIL.n14 7.3702
R349 VTAIL.n226 VTAIL.n188 7.3702
R350 VTAIL.n222 VTAIL.n190 7.3702
R351 VTAIL.n140 VTAIL.n102 7.3702
R352 VTAIL.n136 VTAIL.n104 7.3702
R353 VTAIL.n309 VTAIL.n274 6.59444
R354 VTAIL.n310 VTAIL.n309 6.59444
R355 VTAIL.n51 VTAIL.n16 6.59444
R356 VTAIL.n52 VTAIL.n51 6.59444
R357 VTAIL.n226 VTAIL.n225 6.59444
R358 VTAIL.n225 VTAIL.n190 6.59444
R359 VTAIL.n140 VTAIL.n139 6.59444
R360 VTAIL.n139 VTAIL.n104 6.59444
R361 VTAIL.n306 VTAIL.n305 5.81868
R362 VTAIL.n313 VTAIL.n272 5.81868
R363 VTAIL.n48 VTAIL.n47 5.81868
R364 VTAIL.n55 VTAIL.n14 5.81868
R365 VTAIL.n229 VTAIL.n188 5.81868
R366 VTAIL.n222 VTAIL.n221 5.81868
R367 VTAIL.n143 VTAIL.n102 5.81868
R368 VTAIL.n136 VTAIL.n135 5.81868
R369 VTAIL.n302 VTAIL.n276 5.04292
R370 VTAIL.n314 VTAIL.n270 5.04292
R371 VTAIL.n44 VTAIL.n18 5.04292
R372 VTAIL.n56 VTAIL.n12 5.04292
R373 VTAIL.n230 VTAIL.n186 5.04292
R374 VTAIL.n218 VTAIL.n192 5.04292
R375 VTAIL.n144 VTAIL.n100 5.04292
R376 VTAIL.n132 VTAIL.n106 5.04292
R377 VTAIL.n285 VTAIL.n283 4.38563
R378 VTAIL.n27 VTAIL.n25 4.38563
R379 VTAIL.n201 VTAIL.n199 4.38563
R380 VTAIL.n115 VTAIL.n113 4.38563
R381 VTAIL.n301 VTAIL.n278 4.26717
R382 VTAIL.n318 VTAIL.n317 4.26717
R383 VTAIL.n43 VTAIL.n20 4.26717
R384 VTAIL.n60 VTAIL.n59 4.26717
R385 VTAIL.n234 VTAIL.n233 4.26717
R386 VTAIL.n217 VTAIL.n194 4.26717
R387 VTAIL.n148 VTAIL.n147 4.26717
R388 VTAIL.n131 VTAIL.n108 4.26717
R389 VTAIL.n298 VTAIL.n297 3.49141
R390 VTAIL.n321 VTAIL.n268 3.49141
R391 VTAIL.n40 VTAIL.n39 3.49141
R392 VTAIL.n63 VTAIL.n10 3.49141
R393 VTAIL.n237 VTAIL.n184 3.49141
R394 VTAIL.n214 VTAIL.n213 3.49141
R395 VTAIL.n151 VTAIL.n98 3.49141
R396 VTAIL.n128 VTAIL.n127 3.49141
R397 VTAIL.n294 VTAIL.n280 2.71565
R398 VTAIL.n322 VTAIL.n266 2.71565
R399 VTAIL.n342 VTAIL.n258 2.71565
R400 VTAIL.n36 VTAIL.n22 2.71565
R401 VTAIL.n64 VTAIL.n8 2.71565
R402 VTAIL.n84 VTAIL.n0 2.71565
R403 VTAIL.n256 VTAIL.n172 2.71565
R404 VTAIL.n238 VTAIL.n182 2.71565
R405 VTAIL.n210 VTAIL.n196 2.71565
R406 VTAIL.n170 VTAIL.n86 2.71565
R407 VTAIL.n152 VTAIL.n96 2.71565
R408 VTAIL.n124 VTAIL.n110 2.71565
R409 VTAIL.n257 VTAIL.n171 2.07809
R410 VTAIL.n293 VTAIL.n282 1.93989
R411 VTAIL.n327 VTAIL.n325 1.93989
R412 VTAIL.n340 VTAIL.n339 1.93989
R413 VTAIL.n35 VTAIL.n24 1.93989
R414 VTAIL.n69 VTAIL.n67 1.93989
R415 VTAIL.n82 VTAIL.n81 1.93989
R416 VTAIL.n254 VTAIL.n253 1.93989
R417 VTAIL.n242 VTAIL.n241 1.93989
R418 VTAIL.n209 VTAIL.n198 1.93989
R419 VTAIL.n168 VTAIL.n167 1.93989
R420 VTAIL.n156 VTAIL.n155 1.93989
R421 VTAIL.n123 VTAIL.n112 1.93989
R422 VTAIL VTAIL.n85 1.3324
R423 VTAIL.n290 VTAIL.n289 1.16414
R424 VTAIL.n326 VTAIL.n264 1.16414
R425 VTAIL.n336 VTAIL.n260 1.16414
R426 VTAIL.n32 VTAIL.n31 1.16414
R427 VTAIL.n68 VTAIL.n6 1.16414
R428 VTAIL.n78 VTAIL.n2 1.16414
R429 VTAIL.n250 VTAIL.n174 1.16414
R430 VTAIL.n245 VTAIL.n179 1.16414
R431 VTAIL.n206 VTAIL.n205 1.16414
R432 VTAIL.n164 VTAIL.n88 1.16414
R433 VTAIL.n159 VTAIL.n93 1.16414
R434 VTAIL.n120 VTAIL.n119 1.16414
R435 VTAIL VTAIL.n343 0.74619
R436 VTAIL.n286 VTAIL.n284 0.388379
R437 VTAIL.n332 VTAIL.n331 0.388379
R438 VTAIL.n335 VTAIL.n262 0.388379
R439 VTAIL.n28 VTAIL.n26 0.388379
R440 VTAIL.n74 VTAIL.n73 0.388379
R441 VTAIL.n77 VTAIL.n4 0.388379
R442 VTAIL.n249 VTAIL.n176 0.388379
R443 VTAIL.n246 VTAIL.n178 0.388379
R444 VTAIL.n202 VTAIL.n200 0.388379
R445 VTAIL.n163 VTAIL.n90 0.388379
R446 VTAIL.n160 VTAIL.n92 0.388379
R447 VTAIL.n116 VTAIL.n114 0.388379
R448 VTAIL.n291 VTAIL.n283 0.155672
R449 VTAIL.n292 VTAIL.n291 0.155672
R450 VTAIL.n292 VTAIL.n279 0.155672
R451 VTAIL.n299 VTAIL.n279 0.155672
R452 VTAIL.n300 VTAIL.n299 0.155672
R453 VTAIL.n300 VTAIL.n275 0.155672
R454 VTAIL.n307 VTAIL.n275 0.155672
R455 VTAIL.n308 VTAIL.n307 0.155672
R456 VTAIL.n308 VTAIL.n271 0.155672
R457 VTAIL.n315 VTAIL.n271 0.155672
R458 VTAIL.n316 VTAIL.n315 0.155672
R459 VTAIL.n316 VTAIL.n267 0.155672
R460 VTAIL.n323 VTAIL.n267 0.155672
R461 VTAIL.n324 VTAIL.n323 0.155672
R462 VTAIL.n324 VTAIL.n263 0.155672
R463 VTAIL.n333 VTAIL.n263 0.155672
R464 VTAIL.n334 VTAIL.n333 0.155672
R465 VTAIL.n334 VTAIL.n259 0.155672
R466 VTAIL.n341 VTAIL.n259 0.155672
R467 VTAIL.n33 VTAIL.n25 0.155672
R468 VTAIL.n34 VTAIL.n33 0.155672
R469 VTAIL.n34 VTAIL.n21 0.155672
R470 VTAIL.n41 VTAIL.n21 0.155672
R471 VTAIL.n42 VTAIL.n41 0.155672
R472 VTAIL.n42 VTAIL.n17 0.155672
R473 VTAIL.n49 VTAIL.n17 0.155672
R474 VTAIL.n50 VTAIL.n49 0.155672
R475 VTAIL.n50 VTAIL.n13 0.155672
R476 VTAIL.n57 VTAIL.n13 0.155672
R477 VTAIL.n58 VTAIL.n57 0.155672
R478 VTAIL.n58 VTAIL.n9 0.155672
R479 VTAIL.n65 VTAIL.n9 0.155672
R480 VTAIL.n66 VTAIL.n65 0.155672
R481 VTAIL.n66 VTAIL.n5 0.155672
R482 VTAIL.n75 VTAIL.n5 0.155672
R483 VTAIL.n76 VTAIL.n75 0.155672
R484 VTAIL.n76 VTAIL.n1 0.155672
R485 VTAIL.n83 VTAIL.n1 0.155672
R486 VTAIL.n255 VTAIL.n173 0.155672
R487 VTAIL.n248 VTAIL.n173 0.155672
R488 VTAIL.n248 VTAIL.n247 0.155672
R489 VTAIL.n247 VTAIL.n177 0.155672
R490 VTAIL.n240 VTAIL.n177 0.155672
R491 VTAIL.n240 VTAIL.n239 0.155672
R492 VTAIL.n239 VTAIL.n183 0.155672
R493 VTAIL.n232 VTAIL.n183 0.155672
R494 VTAIL.n232 VTAIL.n231 0.155672
R495 VTAIL.n231 VTAIL.n187 0.155672
R496 VTAIL.n224 VTAIL.n187 0.155672
R497 VTAIL.n224 VTAIL.n223 0.155672
R498 VTAIL.n223 VTAIL.n191 0.155672
R499 VTAIL.n216 VTAIL.n191 0.155672
R500 VTAIL.n216 VTAIL.n215 0.155672
R501 VTAIL.n215 VTAIL.n195 0.155672
R502 VTAIL.n208 VTAIL.n195 0.155672
R503 VTAIL.n208 VTAIL.n207 0.155672
R504 VTAIL.n207 VTAIL.n199 0.155672
R505 VTAIL.n169 VTAIL.n87 0.155672
R506 VTAIL.n162 VTAIL.n87 0.155672
R507 VTAIL.n162 VTAIL.n161 0.155672
R508 VTAIL.n161 VTAIL.n91 0.155672
R509 VTAIL.n154 VTAIL.n91 0.155672
R510 VTAIL.n154 VTAIL.n153 0.155672
R511 VTAIL.n153 VTAIL.n97 0.155672
R512 VTAIL.n146 VTAIL.n97 0.155672
R513 VTAIL.n146 VTAIL.n145 0.155672
R514 VTAIL.n145 VTAIL.n101 0.155672
R515 VTAIL.n138 VTAIL.n101 0.155672
R516 VTAIL.n138 VTAIL.n137 0.155672
R517 VTAIL.n137 VTAIL.n105 0.155672
R518 VTAIL.n130 VTAIL.n105 0.155672
R519 VTAIL.n130 VTAIL.n129 0.155672
R520 VTAIL.n129 VTAIL.n109 0.155672
R521 VTAIL.n122 VTAIL.n109 0.155672
R522 VTAIL.n122 VTAIL.n121 0.155672
R523 VTAIL.n121 VTAIL.n113 0.155672
R524 VDD1.n80 VDD1.n0 289.615
R525 VDD1.n165 VDD1.n85 289.615
R526 VDD1.n81 VDD1.n80 185
R527 VDD1.n79 VDD1.n78 185
R528 VDD1.n4 VDD1.n3 185
R529 VDD1.n8 VDD1.n6 185
R530 VDD1.n73 VDD1.n72 185
R531 VDD1.n71 VDD1.n70 185
R532 VDD1.n10 VDD1.n9 185
R533 VDD1.n65 VDD1.n64 185
R534 VDD1.n63 VDD1.n62 185
R535 VDD1.n14 VDD1.n13 185
R536 VDD1.n57 VDD1.n56 185
R537 VDD1.n55 VDD1.n54 185
R538 VDD1.n18 VDD1.n17 185
R539 VDD1.n49 VDD1.n48 185
R540 VDD1.n47 VDD1.n46 185
R541 VDD1.n22 VDD1.n21 185
R542 VDD1.n41 VDD1.n40 185
R543 VDD1.n39 VDD1.n38 185
R544 VDD1.n26 VDD1.n25 185
R545 VDD1.n33 VDD1.n32 185
R546 VDD1.n31 VDD1.n30 185
R547 VDD1.n114 VDD1.n113 185
R548 VDD1.n116 VDD1.n115 185
R549 VDD1.n109 VDD1.n108 185
R550 VDD1.n122 VDD1.n121 185
R551 VDD1.n124 VDD1.n123 185
R552 VDD1.n105 VDD1.n104 185
R553 VDD1.n130 VDD1.n129 185
R554 VDD1.n132 VDD1.n131 185
R555 VDD1.n101 VDD1.n100 185
R556 VDD1.n138 VDD1.n137 185
R557 VDD1.n140 VDD1.n139 185
R558 VDD1.n97 VDD1.n96 185
R559 VDD1.n146 VDD1.n145 185
R560 VDD1.n148 VDD1.n147 185
R561 VDD1.n93 VDD1.n92 185
R562 VDD1.n155 VDD1.n154 185
R563 VDD1.n156 VDD1.n91 185
R564 VDD1.n158 VDD1.n157 185
R565 VDD1.n89 VDD1.n88 185
R566 VDD1.n164 VDD1.n163 185
R567 VDD1.n166 VDD1.n165 185
R568 VDD1.n29 VDD1.t0 147.659
R569 VDD1.n112 VDD1.t1 147.659
R570 VDD1.n80 VDD1.n79 104.615
R571 VDD1.n79 VDD1.n3 104.615
R572 VDD1.n8 VDD1.n3 104.615
R573 VDD1.n72 VDD1.n8 104.615
R574 VDD1.n72 VDD1.n71 104.615
R575 VDD1.n71 VDD1.n9 104.615
R576 VDD1.n64 VDD1.n9 104.615
R577 VDD1.n64 VDD1.n63 104.615
R578 VDD1.n63 VDD1.n13 104.615
R579 VDD1.n56 VDD1.n13 104.615
R580 VDD1.n56 VDD1.n55 104.615
R581 VDD1.n55 VDD1.n17 104.615
R582 VDD1.n48 VDD1.n17 104.615
R583 VDD1.n48 VDD1.n47 104.615
R584 VDD1.n47 VDD1.n21 104.615
R585 VDD1.n40 VDD1.n21 104.615
R586 VDD1.n40 VDD1.n39 104.615
R587 VDD1.n39 VDD1.n25 104.615
R588 VDD1.n32 VDD1.n25 104.615
R589 VDD1.n32 VDD1.n31 104.615
R590 VDD1.n115 VDD1.n114 104.615
R591 VDD1.n115 VDD1.n108 104.615
R592 VDD1.n122 VDD1.n108 104.615
R593 VDD1.n123 VDD1.n122 104.615
R594 VDD1.n123 VDD1.n104 104.615
R595 VDD1.n130 VDD1.n104 104.615
R596 VDD1.n131 VDD1.n130 104.615
R597 VDD1.n131 VDD1.n100 104.615
R598 VDD1.n138 VDD1.n100 104.615
R599 VDD1.n139 VDD1.n138 104.615
R600 VDD1.n139 VDD1.n96 104.615
R601 VDD1.n146 VDD1.n96 104.615
R602 VDD1.n147 VDD1.n146 104.615
R603 VDD1.n147 VDD1.n92 104.615
R604 VDD1.n155 VDD1.n92 104.615
R605 VDD1.n156 VDD1.n155 104.615
R606 VDD1.n157 VDD1.n156 104.615
R607 VDD1.n157 VDD1.n88 104.615
R608 VDD1.n164 VDD1.n88 104.615
R609 VDD1.n165 VDD1.n164 104.615
R610 VDD1 VDD1.n169 98.1836
R611 VDD1 VDD1.n84 54.1868
R612 VDD1.n31 VDD1.t0 52.3082
R613 VDD1.n114 VDD1.t1 52.3082
R614 VDD1.n30 VDD1.n29 15.6677
R615 VDD1.n113 VDD1.n112 15.6677
R616 VDD1.n6 VDD1.n4 13.1884
R617 VDD1.n158 VDD1.n89 13.1884
R618 VDD1.n78 VDD1.n77 12.8005
R619 VDD1.n74 VDD1.n73 12.8005
R620 VDD1.n33 VDD1.n28 12.8005
R621 VDD1.n116 VDD1.n111 12.8005
R622 VDD1.n159 VDD1.n91 12.8005
R623 VDD1.n163 VDD1.n162 12.8005
R624 VDD1.n81 VDD1.n2 12.0247
R625 VDD1.n70 VDD1.n7 12.0247
R626 VDD1.n34 VDD1.n26 12.0247
R627 VDD1.n117 VDD1.n109 12.0247
R628 VDD1.n154 VDD1.n153 12.0247
R629 VDD1.n166 VDD1.n87 12.0247
R630 VDD1.n82 VDD1.n0 11.249
R631 VDD1.n69 VDD1.n10 11.249
R632 VDD1.n38 VDD1.n37 11.249
R633 VDD1.n121 VDD1.n120 11.249
R634 VDD1.n152 VDD1.n93 11.249
R635 VDD1.n167 VDD1.n85 11.249
R636 VDD1.n66 VDD1.n65 10.4732
R637 VDD1.n41 VDD1.n24 10.4732
R638 VDD1.n124 VDD1.n107 10.4732
R639 VDD1.n149 VDD1.n148 10.4732
R640 VDD1.n62 VDD1.n12 9.69747
R641 VDD1.n42 VDD1.n22 9.69747
R642 VDD1.n125 VDD1.n105 9.69747
R643 VDD1.n145 VDD1.n95 9.69747
R644 VDD1.n84 VDD1.n83 9.45567
R645 VDD1.n169 VDD1.n168 9.45567
R646 VDD1.n16 VDD1.n15 9.3005
R647 VDD1.n59 VDD1.n58 9.3005
R648 VDD1.n61 VDD1.n60 9.3005
R649 VDD1.n12 VDD1.n11 9.3005
R650 VDD1.n67 VDD1.n66 9.3005
R651 VDD1.n69 VDD1.n68 9.3005
R652 VDD1.n7 VDD1.n5 9.3005
R653 VDD1.n75 VDD1.n74 9.3005
R654 VDD1.n83 VDD1.n82 9.3005
R655 VDD1.n2 VDD1.n1 9.3005
R656 VDD1.n77 VDD1.n76 9.3005
R657 VDD1.n53 VDD1.n52 9.3005
R658 VDD1.n51 VDD1.n50 9.3005
R659 VDD1.n20 VDD1.n19 9.3005
R660 VDD1.n45 VDD1.n44 9.3005
R661 VDD1.n43 VDD1.n42 9.3005
R662 VDD1.n24 VDD1.n23 9.3005
R663 VDD1.n37 VDD1.n36 9.3005
R664 VDD1.n35 VDD1.n34 9.3005
R665 VDD1.n28 VDD1.n27 9.3005
R666 VDD1.n168 VDD1.n167 9.3005
R667 VDD1.n87 VDD1.n86 9.3005
R668 VDD1.n162 VDD1.n161 9.3005
R669 VDD1.n134 VDD1.n133 9.3005
R670 VDD1.n103 VDD1.n102 9.3005
R671 VDD1.n128 VDD1.n127 9.3005
R672 VDD1.n126 VDD1.n125 9.3005
R673 VDD1.n107 VDD1.n106 9.3005
R674 VDD1.n120 VDD1.n119 9.3005
R675 VDD1.n118 VDD1.n117 9.3005
R676 VDD1.n111 VDD1.n110 9.3005
R677 VDD1.n136 VDD1.n135 9.3005
R678 VDD1.n99 VDD1.n98 9.3005
R679 VDD1.n142 VDD1.n141 9.3005
R680 VDD1.n144 VDD1.n143 9.3005
R681 VDD1.n95 VDD1.n94 9.3005
R682 VDD1.n150 VDD1.n149 9.3005
R683 VDD1.n152 VDD1.n151 9.3005
R684 VDD1.n153 VDD1.n90 9.3005
R685 VDD1.n160 VDD1.n159 9.3005
R686 VDD1.n61 VDD1.n14 8.92171
R687 VDD1.n46 VDD1.n45 8.92171
R688 VDD1.n129 VDD1.n128 8.92171
R689 VDD1.n144 VDD1.n97 8.92171
R690 VDD1.n58 VDD1.n57 8.14595
R691 VDD1.n49 VDD1.n20 8.14595
R692 VDD1.n132 VDD1.n103 8.14595
R693 VDD1.n141 VDD1.n140 8.14595
R694 VDD1.n54 VDD1.n16 7.3702
R695 VDD1.n50 VDD1.n18 7.3702
R696 VDD1.n133 VDD1.n101 7.3702
R697 VDD1.n137 VDD1.n99 7.3702
R698 VDD1.n54 VDD1.n53 6.59444
R699 VDD1.n53 VDD1.n18 6.59444
R700 VDD1.n136 VDD1.n101 6.59444
R701 VDD1.n137 VDD1.n136 6.59444
R702 VDD1.n57 VDD1.n16 5.81868
R703 VDD1.n50 VDD1.n49 5.81868
R704 VDD1.n133 VDD1.n132 5.81868
R705 VDD1.n140 VDD1.n99 5.81868
R706 VDD1.n58 VDD1.n14 5.04292
R707 VDD1.n46 VDD1.n20 5.04292
R708 VDD1.n129 VDD1.n103 5.04292
R709 VDD1.n141 VDD1.n97 5.04292
R710 VDD1.n29 VDD1.n27 4.38563
R711 VDD1.n112 VDD1.n110 4.38563
R712 VDD1.n62 VDD1.n61 4.26717
R713 VDD1.n45 VDD1.n22 4.26717
R714 VDD1.n128 VDD1.n105 4.26717
R715 VDD1.n145 VDD1.n144 4.26717
R716 VDD1.n65 VDD1.n12 3.49141
R717 VDD1.n42 VDD1.n41 3.49141
R718 VDD1.n125 VDD1.n124 3.49141
R719 VDD1.n148 VDD1.n95 3.49141
R720 VDD1.n84 VDD1.n0 2.71565
R721 VDD1.n66 VDD1.n10 2.71565
R722 VDD1.n38 VDD1.n24 2.71565
R723 VDD1.n121 VDD1.n107 2.71565
R724 VDD1.n149 VDD1.n93 2.71565
R725 VDD1.n169 VDD1.n85 2.71565
R726 VDD1.n82 VDD1.n81 1.93989
R727 VDD1.n70 VDD1.n69 1.93989
R728 VDD1.n37 VDD1.n26 1.93989
R729 VDD1.n120 VDD1.n109 1.93989
R730 VDD1.n154 VDD1.n152 1.93989
R731 VDD1.n167 VDD1.n166 1.93989
R732 VDD1.n78 VDD1.n2 1.16414
R733 VDD1.n73 VDD1.n7 1.16414
R734 VDD1.n34 VDD1.n33 1.16414
R735 VDD1.n117 VDD1.n116 1.16414
R736 VDD1.n153 VDD1.n91 1.16414
R737 VDD1.n163 VDD1.n87 1.16414
R738 VDD1.n77 VDD1.n4 0.388379
R739 VDD1.n74 VDD1.n6 0.388379
R740 VDD1.n30 VDD1.n28 0.388379
R741 VDD1.n113 VDD1.n111 0.388379
R742 VDD1.n159 VDD1.n158 0.388379
R743 VDD1.n162 VDD1.n89 0.388379
R744 VDD1.n83 VDD1.n1 0.155672
R745 VDD1.n76 VDD1.n1 0.155672
R746 VDD1.n76 VDD1.n75 0.155672
R747 VDD1.n75 VDD1.n5 0.155672
R748 VDD1.n68 VDD1.n5 0.155672
R749 VDD1.n68 VDD1.n67 0.155672
R750 VDD1.n67 VDD1.n11 0.155672
R751 VDD1.n60 VDD1.n11 0.155672
R752 VDD1.n60 VDD1.n59 0.155672
R753 VDD1.n59 VDD1.n15 0.155672
R754 VDD1.n52 VDD1.n15 0.155672
R755 VDD1.n52 VDD1.n51 0.155672
R756 VDD1.n51 VDD1.n19 0.155672
R757 VDD1.n44 VDD1.n19 0.155672
R758 VDD1.n44 VDD1.n43 0.155672
R759 VDD1.n43 VDD1.n23 0.155672
R760 VDD1.n36 VDD1.n23 0.155672
R761 VDD1.n36 VDD1.n35 0.155672
R762 VDD1.n35 VDD1.n27 0.155672
R763 VDD1.n118 VDD1.n110 0.155672
R764 VDD1.n119 VDD1.n118 0.155672
R765 VDD1.n119 VDD1.n106 0.155672
R766 VDD1.n126 VDD1.n106 0.155672
R767 VDD1.n127 VDD1.n126 0.155672
R768 VDD1.n127 VDD1.n102 0.155672
R769 VDD1.n134 VDD1.n102 0.155672
R770 VDD1.n135 VDD1.n134 0.155672
R771 VDD1.n135 VDD1.n98 0.155672
R772 VDD1.n142 VDD1.n98 0.155672
R773 VDD1.n143 VDD1.n142 0.155672
R774 VDD1.n143 VDD1.n94 0.155672
R775 VDD1.n150 VDD1.n94 0.155672
R776 VDD1.n151 VDD1.n150 0.155672
R777 VDD1.n151 VDD1.n90 0.155672
R778 VDD1.n160 VDD1.n90 0.155672
R779 VDD1.n161 VDD1.n160 0.155672
R780 VDD1.n161 VDD1.n86 0.155672
R781 VDD1.n168 VDD1.n86 0.155672
R782 B.n597 B.n596 585
R783 B.n599 B.n119 585
R784 B.n602 B.n601 585
R785 B.n603 B.n118 585
R786 B.n605 B.n604 585
R787 B.n607 B.n117 585
R788 B.n610 B.n609 585
R789 B.n611 B.n116 585
R790 B.n613 B.n612 585
R791 B.n615 B.n115 585
R792 B.n618 B.n617 585
R793 B.n619 B.n114 585
R794 B.n621 B.n620 585
R795 B.n623 B.n113 585
R796 B.n626 B.n625 585
R797 B.n627 B.n112 585
R798 B.n629 B.n628 585
R799 B.n631 B.n111 585
R800 B.n634 B.n633 585
R801 B.n635 B.n110 585
R802 B.n637 B.n636 585
R803 B.n639 B.n109 585
R804 B.n642 B.n641 585
R805 B.n643 B.n108 585
R806 B.n645 B.n644 585
R807 B.n647 B.n107 585
R808 B.n650 B.n649 585
R809 B.n651 B.n106 585
R810 B.n653 B.n652 585
R811 B.n655 B.n105 585
R812 B.n658 B.n657 585
R813 B.n659 B.n104 585
R814 B.n661 B.n660 585
R815 B.n663 B.n103 585
R816 B.n666 B.n665 585
R817 B.n667 B.n102 585
R818 B.n669 B.n668 585
R819 B.n671 B.n101 585
R820 B.n674 B.n673 585
R821 B.n675 B.n100 585
R822 B.n677 B.n676 585
R823 B.n679 B.n99 585
R824 B.n682 B.n681 585
R825 B.n683 B.n98 585
R826 B.n685 B.n684 585
R827 B.n687 B.n97 585
R828 B.n690 B.n689 585
R829 B.n691 B.n96 585
R830 B.n693 B.n692 585
R831 B.n695 B.n95 585
R832 B.n697 B.n696 585
R833 B.n699 B.n698 585
R834 B.n702 B.n701 585
R835 B.n703 B.n90 585
R836 B.n705 B.n704 585
R837 B.n707 B.n89 585
R838 B.n710 B.n709 585
R839 B.n711 B.n88 585
R840 B.n713 B.n712 585
R841 B.n715 B.n87 585
R842 B.n718 B.n717 585
R843 B.n719 B.n84 585
R844 B.n722 B.n721 585
R845 B.n724 B.n83 585
R846 B.n727 B.n726 585
R847 B.n728 B.n82 585
R848 B.n730 B.n729 585
R849 B.n732 B.n81 585
R850 B.n735 B.n734 585
R851 B.n736 B.n80 585
R852 B.n738 B.n737 585
R853 B.n740 B.n79 585
R854 B.n743 B.n742 585
R855 B.n744 B.n78 585
R856 B.n746 B.n745 585
R857 B.n748 B.n77 585
R858 B.n751 B.n750 585
R859 B.n752 B.n76 585
R860 B.n754 B.n753 585
R861 B.n756 B.n75 585
R862 B.n759 B.n758 585
R863 B.n760 B.n74 585
R864 B.n762 B.n761 585
R865 B.n764 B.n73 585
R866 B.n767 B.n766 585
R867 B.n768 B.n72 585
R868 B.n770 B.n769 585
R869 B.n772 B.n71 585
R870 B.n775 B.n774 585
R871 B.n776 B.n70 585
R872 B.n778 B.n777 585
R873 B.n780 B.n69 585
R874 B.n783 B.n782 585
R875 B.n784 B.n68 585
R876 B.n786 B.n785 585
R877 B.n788 B.n67 585
R878 B.n791 B.n790 585
R879 B.n792 B.n66 585
R880 B.n794 B.n793 585
R881 B.n796 B.n65 585
R882 B.n799 B.n798 585
R883 B.n800 B.n64 585
R884 B.n802 B.n801 585
R885 B.n804 B.n63 585
R886 B.n807 B.n806 585
R887 B.n808 B.n62 585
R888 B.n810 B.n809 585
R889 B.n812 B.n61 585
R890 B.n815 B.n814 585
R891 B.n816 B.n60 585
R892 B.n818 B.n817 585
R893 B.n820 B.n59 585
R894 B.n823 B.n822 585
R895 B.n824 B.n58 585
R896 B.n595 B.n56 585
R897 B.n827 B.n56 585
R898 B.n594 B.n55 585
R899 B.n828 B.n55 585
R900 B.n593 B.n54 585
R901 B.n829 B.n54 585
R902 B.n592 B.n591 585
R903 B.n591 B.n50 585
R904 B.n590 B.n49 585
R905 B.n835 B.n49 585
R906 B.n589 B.n48 585
R907 B.n836 B.n48 585
R908 B.n588 B.n47 585
R909 B.n837 B.n47 585
R910 B.n587 B.n586 585
R911 B.n586 B.n43 585
R912 B.n585 B.n42 585
R913 B.n843 B.n42 585
R914 B.n584 B.n41 585
R915 B.n844 B.n41 585
R916 B.n583 B.n40 585
R917 B.n845 B.n40 585
R918 B.n582 B.n581 585
R919 B.n581 B.n36 585
R920 B.n580 B.n35 585
R921 B.n851 B.n35 585
R922 B.n579 B.n34 585
R923 B.n852 B.n34 585
R924 B.n578 B.n33 585
R925 B.n853 B.n33 585
R926 B.n577 B.n576 585
R927 B.n576 B.n29 585
R928 B.n575 B.n28 585
R929 B.n859 B.n28 585
R930 B.n574 B.n27 585
R931 B.n860 B.n27 585
R932 B.n573 B.n26 585
R933 B.n861 B.n26 585
R934 B.n572 B.n571 585
R935 B.n571 B.n22 585
R936 B.n570 B.n21 585
R937 B.n867 B.n21 585
R938 B.n569 B.n20 585
R939 B.n868 B.n20 585
R940 B.n568 B.n19 585
R941 B.n869 B.n19 585
R942 B.n567 B.n566 585
R943 B.n566 B.n15 585
R944 B.n565 B.n14 585
R945 B.n875 B.n14 585
R946 B.n564 B.n13 585
R947 B.n876 B.n13 585
R948 B.n563 B.n12 585
R949 B.n877 B.n12 585
R950 B.n562 B.n561 585
R951 B.n561 B.n8 585
R952 B.n560 B.n7 585
R953 B.n883 B.n7 585
R954 B.n559 B.n6 585
R955 B.n884 B.n6 585
R956 B.n558 B.n5 585
R957 B.n885 B.n5 585
R958 B.n557 B.n556 585
R959 B.n556 B.n4 585
R960 B.n555 B.n120 585
R961 B.n555 B.n554 585
R962 B.n545 B.n121 585
R963 B.n122 B.n121 585
R964 B.n547 B.n546 585
R965 B.n548 B.n547 585
R966 B.n544 B.n127 585
R967 B.n127 B.n126 585
R968 B.n543 B.n542 585
R969 B.n542 B.n541 585
R970 B.n129 B.n128 585
R971 B.n130 B.n129 585
R972 B.n534 B.n533 585
R973 B.n535 B.n534 585
R974 B.n532 B.n135 585
R975 B.n135 B.n134 585
R976 B.n531 B.n530 585
R977 B.n530 B.n529 585
R978 B.n137 B.n136 585
R979 B.n138 B.n137 585
R980 B.n522 B.n521 585
R981 B.n523 B.n522 585
R982 B.n520 B.n143 585
R983 B.n143 B.n142 585
R984 B.n519 B.n518 585
R985 B.n518 B.n517 585
R986 B.n145 B.n144 585
R987 B.n146 B.n145 585
R988 B.n510 B.n509 585
R989 B.n511 B.n510 585
R990 B.n508 B.n151 585
R991 B.n151 B.n150 585
R992 B.n507 B.n506 585
R993 B.n506 B.n505 585
R994 B.n153 B.n152 585
R995 B.n154 B.n153 585
R996 B.n498 B.n497 585
R997 B.n499 B.n498 585
R998 B.n496 B.n159 585
R999 B.n159 B.n158 585
R1000 B.n495 B.n494 585
R1001 B.n494 B.n493 585
R1002 B.n161 B.n160 585
R1003 B.n162 B.n161 585
R1004 B.n486 B.n485 585
R1005 B.n487 B.n486 585
R1006 B.n484 B.n167 585
R1007 B.n167 B.n166 585
R1008 B.n483 B.n482 585
R1009 B.n482 B.n481 585
R1010 B.n169 B.n168 585
R1011 B.n170 B.n169 585
R1012 B.n474 B.n473 585
R1013 B.n475 B.n474 585
R1014 B.n472 B.n175 585
R1015 B.n175 B.n174 585
R1016 B.n471 B.n470 585
R1017 B.n470 B.n469 585
R1018 B.n466 B.n179 585
R1019 B.n465 B.n464 585
R1020 B.n462 B.n180 585
R1021 B.n462 B.n178 585
R1022 B.n461 B.n460 585
R1023 B.n459 B.n458 585
R1024 B.n457 B.n182 585
R1025 B.n455 B.n454 585
R1026 B.n453 B.n183 585
R1027 B.n452 B.n451 585
R1028 B.n449 B.n184 585
R1029 B.n447 B.n446 585
R1030 B.n445 B.n185 585
R1031 B.n444 B.n443 585
R1032 B.n441 B.n186 585
R1033 B.n439 B.n438 585
R1034 B.n437 B.n187 585
R1035 B.n436 B.n435 585
R1036 B.n433 B.n188 585
R1037 B.n431 B.n430 585
R1038 B.n429 B.n189 585
R1039 B.n428 B.n427 585
R1040 B.n425 B.n190 585
R1041 B.n423 B.n422 585
R1042 B.n421 B.n191 585
R1043 B.n420 B.n419 585
R1044 B.n417 B.n192 585
R1045 B.n415 B.n414 585
R1046 B.n413 B.n193 585
R1047 B.n412 B.n411 585
R1048 B.n409 B.n194 585
R1049 B.n407 B.n406 585
R1050 B.n405 B.n195 585
R1051 B.n404 B.n403 585
R1052 B.n401 B.n196 585
R1053 B.n399 B.n398 585
R1054 B.n397 B.n197 585
R1055 B.n396 B.n395 585
R1056 B.n393 B.n198 585
R1057 B.n391 B.n390 585
R1058 B.n389 B.n199 585
R1059 B.n388 B.n387 585
R1060 B.n385 B.n200 585
R1061 B.n383 B.n382 585
R1062 B.n381 B.n201 585
R1063 B.n380 B.n379 585
R1064 B.n377 B.n202 585
R1065 B.n375 B.n374 585
R1066 B.n373 B.n203 585
R1067 B.n372 B.n371 585
R1068 B.n369 B.n204 585
R1069 B.n367 B.n366 585
R1070 B.n365 B.n205 585
R1071 B.n363 B.n362 585
R1072 B.n360 B.n208 585
R1073 B.n358 B.n357 585
R1074 B.n356 B.n209 585
R1075 B.n355 B.n354 585
R1076 B.n352 B.n210 585
R1077 B.n350 B.n349 585
R1078 B.n348 B.n211 585
R1079 B.n347 B.n346 585
R1080 B.n344 B.n212 585
R1081 B.n342 B.n341 585
R1082 B.n340 B.n213 585
R1083 B.n339 B.n338 585
R1084 B.n336 B.n217 585
R1085 B.n334 B.n333 585
R1086 B.n332 B.n218 585
R1087 B.n331 B.n330 585
R1088 B.n328 B.n219 585
R1089 B.n326 B.n325 585
R1090 B.n324 B.n220 585
R1091 B.n323 B.n322 585
R1092 B.n320 B.n221 585
R1093 B.n318 B.n317 585
R1094 B.n316 B.n222 585
R1095 B.n315 B.n314 585
R1096 B.n312 B.n223 585
R1097 B.n310 B.n309 585
R1098 B.n308 B.n224 585
R1099 B.n307 B.n306 585
R1100 B.n304 B.n225 585
R1101 B.n302 B.n301 585
R1102 B.n300 B.n226 585
R1103 B.n299 B.n298 585
R1104 B.n296 B.n227 585
R1105 B.n294 B.n293 585
R1106 B.n292 B.n228 585
R1107 B.n291 B.n290 585
R1108 B.n288 B.n229 585
R1109 B.n286 B.n285 585
R1110 B.n284 B.n230 585
R1111 B.n283 B.n282 585
R1112 B.n280 B.n231 585
R1113 B.n278 B.n277 585
R1114 B.n276 B.n232 585
R1115 B.n275 B.n274 585
R1116 B.n272 B.n233 585
R1117 B.n270 B.n269 585
R1118 B.n268 B.n234 585
R1119 B.n267 B.n266 585
R1120 B.n264 B.n235 585
R1121 B.n262 B.n261 585
R1122 B.n260 B.n236 585
R1123 B.n259 B.n258 585
R1124 B.n256 B.n237 585
R1125 B.n254 B.n253 585
R1126 B.n252 B.n238 585
R1127 B.n251 B.n250 585
R1128 B.n248 B.n239 585
R1129 B.n246 B.n245 585
R1130 B.n244 B.n240 585
R1131 B.n243 B.n242 585
R1132 B.n177 B.n176 585
R1133 B.n178 B.n177 585
R1134 B.n468 B.n467 585
R1135 B.n469 B.n468 585
R1136 B.n173 B.n172 585
R1137 B.n174 B.n173 585
R1138 B.n477 B.n476 585
R1139 B.n476 B.n475 585
R1140 B.n478 B.n171 585
R1141 B.n171 B.n170 585
R1142 B.n480 B.n479 585
R1143 B.n481 B.n480 585
R1144 B.n165 B.n164 585
R1145 B.n166 B.n165 585
R1146 B.n489 B.n488 585
R1147 B.n488 B.n487 585
R1148 B.n490 B.n163 585
R1149 B.n163 B.n162 585
R1150 B.n492 B.n491 585
R1151 B.n493 B.n492 585
R1152 B.n157 B.n156 585
R1153 B.n158 B.n157 585
R1154 B.n501 B.n500 585
R1155 B.n500 B.n499 585
R1156 B.n502 B.n155 585
R1157 B.n155 B.n154 585
R1158 B.n504 B.n503 585
R1159 B.n505 B.n504 585
R1160 B.n149 B.n148 585
R1161 B.n150 B.n149 585
R1162 B.n513 B.n512 585
R1163 B.n512 B.n511 585
R1164 B.n514 B.n147 585
R1165 B.n147 B.n146 585
R1166 B.n516 B.n515 585
R1167 B.n517 B.n516 585
R1168 B.n141 B.n140 585
R1169 B.n142 B.n141 585
R1170 B.n525 B.n524 585
R1171 B.n524 B.n523 585
R1172 B.n526 B.n139 585
R1173 B.n139 B.n138 585
R1174 B.n528 B.n527 585
R1175 B.n529 B.n528 585
R1176 B.n133 B.n132 585
R1177 B.n134 B.n133 585
R1178 B.n537 B.n536 585
R1179 B.n536 B.n535 585
R1180 B.n538 B.n131 585
R1181 B.n131 B.n130 585
R1182 B.n540 B.n539 585
R1183 B.n541 B.n540 585
R1184 B.n125 B.n124 585
R1185 B.n126 B.n125 585
R1186 B.n550 B.n549 585
R1187 B.n549 B.n548 585
R1188 B.n551 B.n123 585
R1189 B.n123 B.n122 585
R1190 B.n553 B.n552 585
R1191 B.n554 B.n553 585
R1192 B.n2 B.n0 585
R1193 B.n4 B.n2 585
R1194 B.n3 B.n1 585
R1195 B.n884 B.n3 585
R1196 B.n882 B.n881 585
R1197 B.n883 B.n882 585
R1198 B.n880 B.n9 585
R1199 B.n9 B.n8 585
R1200 B.n879 B.n878 585
R1201 B.n878 B.n877 585
R1202 B.n11 B.n10 585
R1203 B.n876 B.n11 585
R1204 B.n874 B.n873 585
R1205 B.n875 B.n874 585
R1206 B.n872 B.n16 585
R1207 B.n16 B.n15 585
R1208 B.n871 B.n870 585
R1209 B.n870 B.n869 585
R1210 B.n18 B.n17 585
R1211 B.n868 B.n18 585
R1212 B.n866 B.n865 585
R1213 B.n867 B.n866 585
R1214 B.n864 B.n23 585
R1215 B.n23 B.n22 585
R1216 B.n863 B.n862 585
R1217 B.n862 B.n861 585
R1218 B.n25 B.n24 585
R1219 B.n860 B.n25 585
R1220 B.n858 B.n857 585
R1221 B.n859 B.n858 585
R1222 B.n856 B.n30 585
R1223 B.n30 B.n29 585
R1224 B.n855 B.n854 585
R1225 B.n854 B.n853 585
R1226 B.n32 B.n31 585
R1227 B.n852 B.n32 585
R1228 B.n850 B.n849 585
R1229 B.n851 B.n850 585
R1230 B.n848 B.n37 585
R1231 B.n37 B.n36 585
R1232 B.n847 B.n846 585
R1233 B.n846 B.n845 585
R1234 B.n39 B.n38 585
R1235 B.n844 B.n39 585
R1236 B.n842 B.n841 585
R1237 B.n843 B.n842 585
R1238 B.n840 B.n44 585
R1239 B.n44 B.n43 585
R1240 B.n839 B.n838 585
R1241 B.n838 B.n837 585
R1242 B.n46 B.n45 585
R1243 B.n836 B.n46 585
R1244 B.n834 B.n833 585
R1245 B.n835 B.n834 585
R1246 B.n832 B.n51 585
R1247 B.n51 B.n50 585
R1248 B.n831 B.n830 585
R1249 B.n830 B.n829 585
R1250 B.n53 B.n52 585
R1251 B.n828 B.n53 585
R1252 B.n826 B.n825 585
R1253 B.n827 B.n826 585
R1254 B.n887 B.n886 585
R1255 B.n886 B.n885 585
R1256 B.n468 B.n179 502.111
R1257 B.n826 B.n58 502.111
R1258 B.n470 B.n177 502.111
R1259 B.n597 B.n56 502.111
R1260 B.n214 B.t5 416.594
R1261 B.n91 B.t8 416.594
R1262 B.n206 B.t12 416.594
R1263 B.n85 B.t14 416.594
R1264 B.n215 B.t4 344.255
R1265 B.n92 B.t9 344.255
R1266 B.n207 B.t11 344.255
R1267 B.n86 B.t15 344.255
R1268 B.n214 B.t2 319.507
R1269 B.n206 B.t10 319.507
R1270 B.n85 B.t13 319.507
R1271 B.n91 B.t6 319.507
R1272 B.n598 B.n57 256.663
R1273 B.n600 B.n57 256.663
R1274 B.n606 B.n57 256.663
R1275 B.n608 B.n57 256.663
R1276 B.n614 B.n57 256.663
R1277 B.n616 B.n57 256.663
R1278 B.n622 B.n57 256.663
R1279 B.n624 B.n57 256.663
R1280 B.n630 B.n57 256.663
R1281 B.n632 B.n57 256.663
R1282 B.n638 B.n57 256.663
R1283 B.n640 B.n57 256.663
R1284 B.n646 B.n57 256.663
R1285 B.n648 B.n57 256.663
R1286 B.n654 B.n57 256.663
R1287 B.n656 B.n57 256.663
R1288 B.n662 B.n57 256.663
R1289 B.n664 B.n57 256.663
R1290 B.n670 B.n57 256.663
R1291 B.n672 B.n57 256.663
R1292 B.n678 B.n57 256.663
R1293 B.n680 B.n57 256.663
R1294 B.n686 B.n57 256.663
R1295 B.n688 B.n57 256.663
R1296 B.n694 B.n57 256.663
R1297 B.n94 B.n57 256.663
R1298 B.n700 B.n57 256.663
R1299 B.n706 B.n57 256.663
R1300 B.n708 B.n57 256.663
R1301 B.n714 B.n57 256.663
R1302 B.n716 B.n57 256.663
R1303 B.n723 B.n57 256.663
R1304 B.n725 B.n57 256.663
R1305 B.n731 B.n57 256.663
R1306 B.n733 B.n57 256.663
R1307 B.n739 B.n57 256.663
R1308 B.n741 B.n57 256.663
R1309 B.n747 B.n57 256.663
R1310 B.n749 B.n57 256.663
R1311 B.n755 B.n57 256.663
R1312 B.n757 B.n57 256.663
R1313 B.n763 B.n57 256.663
R1314 B.n765 B.n57 256.663
R1315 B.n771 B.n57 256.663
R1316 B.n773 B.n57 256.663
R1317 B.n779 B.n57 256.663
R1318 B.n781 B.n57 256.663
R1319 B.n787 B.n57 256.663
R1320 B.n789 B.n57 256.663
R1321 B.n795 B.n57 256.663
R1322 B.n797 B.n57 256.663
R1323 B.n803 B.n57 256.663
R1324 B.n805 B.n57 256.663
R1325 B.n811 B.n57 256.663
R1326 B.n813 B.n57 256.663
R1327 B.n819 B.n57 256.663
R1328 B.n821 B.n57 256.663
R1329 B.n463 B.n178 256.663
R1330 B.n181 B.n178 256.663
R1331 B.n456 B.n178 256.663
R1332 B.n450 B.n178 256.663
R1333 B.n448 B.n178 256.663
R1334 B.n442 B.n178 256.663
R1335 B.n440 B.n178 256.663
R1336 B.n434 B.n178 256.663
R1337 B.n432 B.n178 256.663
R1338 B.n426 B.n178 256.663
R1339 B.n424 B.n178 256.663
R1340 B.n418 B.n178 256.663
R1341 B.n416 B.n178 256.663
R1342 B.n410 B.n178 256.663
R1343 B.n408 B.n178 256.663
R1344 B.n402 B.n178 256.663
R1345 B.n400 B.n178 256.663
R1346 B.n394 B.n178 256.663
R1347 B.n392 B.n178 256.663
R1348 B.n386 B.n178 256.663
R1349 B.n384 B.n178 256.663
R1350 B.n378 B.n178 256.663
R1351 B.n376 B.n178 256.663
R1352 B.n370 B.n178 256.663
R1353 B.n368 B.n178 256.663
R1354 B.n361 B.n178 256.663
R1355 B.n359 B.n178 256.663
R1356 B.n353 B.n178 256.663
R1357 B.n351 B.n178 256.663
R1358 B.n345 B.n178 256.663
R1359 B.n343 B.n178 256.663
R1360 B.n337 B.n178 256.663
R1361 B.n335 B.n178 256.663
R1362 B.n329 B.n178 256.663
R1363 B.n327 B.n178 256.663
R1364 B.n321 B.n178 256.663
R1365 B.n319 B.n178 256.663
R1366 B.n313 B.n178 256.663
R1367 B.n311 B.n178 256.663
R1368 B.n305 B.n178 256.663
R1369 B.n303 B.n178 256.663
R1370 B.n297 B.n178 256.663
R1371 B.n295 B.n178 256.663
R1372 B.n289 B.n178 256.663
R1373 B.n287 B.n178 256.663
R1374 B.n281 B.n178 256.663
R1375 B.n279 B.n178 256.663
R1376 B.n273 B.n178 256.663
R1377 B.n271 B.n178 256.663
R1378 B.n265 B.n178 256.663
R1379 B.n263 B.n178 256.663
R1380 B.n257 B.n178 256.663
R1381 B.n255 B.n178 256.663
R1382 B.n249 B.n178 256.663
R1383 B.n247 B.n178 256.663
R1384 B.n241 B.n178 256.663
R1385 B.n468 B.n173 163.367
R1386 B.n476 B.n173 163.367
R1387 B.n476 B.n171 163.367
R1388 B.n480 B.n171 163.367
R1389 B.n480 B.n165 163.367
R1390 B.n488 B.n165 163.367
R1391 B.n488 B.n163 163.367
R1392 B.n492 B.n163 163.367
R1393 B.n492 B.n157 163.367
R1394 B.n500 B.n157 163.367
R1395 B.n500 B.n155 163.367
R1396 B.n504 B.n155 163.367
R1397 B.n504 B.n149 163.367
R1398 B.n512 B.n149 163.367
R1399 B.n512 B.n147 163.367
R1400 B.n516 B.n147 163.367
R1401 B.n516 B.n141 163.367
R1402 B.n524 B.n141 163.367
R1403 B.n524 B.n139 163.367
R1404 B.n528 B.n139 163.367
R1405 B.n528 B.n133 163.367
R1406 B.n536 B.n133 163.367
R1407 B.n536 B.n131 163.367
R1408 B.n540 B.n131 163.367
R1409 B.n540 B.n125 163.367
R1410 B.n549 B.n125 163.367
R1411 B.n549 B.n123 163.367
R1412 B.n553 B.n123 163.367
R1413 B.n553 B.n2 163.367
R1414 B.n886 B.n2 163.367
R1415 B.n886 B.n3 163.367
R1416 B.n882 B.n3 163.367
R1417 B.n882 B.n9 163.367
R1418 B.n878 B.n9 163.367
R1419 B.n878 B.n11 163.367
R1420 B.n874 B.n11 163.367
R1421 B.n874 B.n16 163.367
R1422 B.n870 B.n16 163.367
R1423 B.n870 B.n18 163.367
R1424 B.n866 B.n18 163.367
R1425 B.n866 B.n23 163.367
R1426 B.n862 B.n23 163.367
R1427 B.n862 B.n25 163.367
R1428 B.n858 B.n25 163.367
R1429 B.n858 B.n30 163.367
R1430 B.n854 B.n30 163.367
R1431 B.n854 B.n32 163.367
R1432 B.n850 B.n32 163.367
R1433 B.n850 B.n37 163.367
R1434 B.n846 B.n37 163.367
R1435 B.n846 B.n39 163.367
R1436 B.n842 B.n39 163.367
R1437 B.n842 B.n44 163.367
R1438 B.n838 B.n44 163.367
R1439 B.n838 B.n46 163.367
R1440 B.n834 B.n46 163.367
R1441 B.n834 B.n51 163.367
R1442 B.n830 B.n51 163.367
R1443 B.n830 B.n53 163.367
R1444 B.n826 B.n53 163.367
R1445 B.n464 B.n462 163.367
R1446 B.n462 B.n461 163.367
R1447 B.n458 B.n457 163.367
R1448 B.n455 B.n183 163.367
R1449 B.n451 B.n449 163.367
R1450 B.n447 B.n185 163.367
R1451 B.n443 B.n441 163.367
R1452 B.n439 B.n187 163.367
R1453 B.n435 B.n433 163.367
R1454 B.n431 B.n189 163.367
R1455 B.n427 B.n425 163.367
R1456 B.n423 B.n191 163.367
R1457 B.n419 B.n417 163.367
R1458 B.n415 B.n193 163.367
R1459 B.n411 B.n409 163.367
R1460 B.n407 B.n195 163.367
R1461 B.n403 B.n401 163.367
R1462 B.n399 B.n197 163.367
R1463 B.n395 B.n393 163.367
R1464 B.n391 B.n199 163.367
R1465 B.n387 B.n385 163.367
R1466 B.n383 B.n201 163.367
R1467 B.n379 B.n377 163.367
R1468 B.n375 B.n203 163.367
R1469 B.n371 B.n369 163.367
R1470 B.n367 B.n205 163.367
R1471 B.n362 B.n360 163.367
R1472 B.n358 B.n209 163.367
R1473 B.n354 B.n352 163.367
R1474 B.n350 B.n211 163.367
R1475 B.n346 B.n344 163.367
R1476 B.n342 B.n213 163.367
R1477 B.n338 B.n336 163.367
R1478 B.n334 B.n218 163.367
R1479 B.n330 B.n328 163.367
R1480 B.n326 B.n220 163.367
R1481 B.n322 B.n320 163.367
R1482 B.n318 B.n222 163.367
R1483 B.n314 B.n312 163.367
R1484 B.n310 B.n224 163.367
R1485 B.n306 B.n304 163.367
R1486 B.n302 B.n226 163.367
R1487 B.n298 B.n296 163.367
R1488 B.n294 B.n228 163.367
R1489 B.n290 B.n288 163.367
R1490 B.n286 B.n230 163.367
R1491 B.n282 B.n280 163.367
R1492 B.n278 B.n232 163.367
R1493 B.n274 B.n272 163.367
R1494 B.n270 B.n234 163.367
R1495 B.n266 B.n264 163.367
R1496 B.n262 B.n236 163.367
R1497 B.n258 B.n256 163.367
R1498 B.n254 B.n238 163.367
R1499 B.n250 B.n248 163.367
R1500 B.n246 B.n240 163.367
R1501 B.n242 B.n177 163.367
R1502 B.n470 B.n175 163.367
R1503 B.n474 B.n175 163.367
R1504 B.n474 B.n169 163.367
R1505 B.n482 B.n169 163.367
R1506 B.n482 B.n167 163.367
R1507 B.n486 B.n167 163.367
R1508 B.n486 B.n161 163.367
R1509 B.n494 B.n161 163.367
R1510 B.n494 B.n159 163.367
R1511 B.n498 B.n159 163.367
R1512 B.n498 B.n153 163.367
R1513 B.n506 B.n153 163.367
R1514 B.n506 B.n151 163.367
R1515 B.n510 B.n151 163.367
R1516 B.n510 B.n145 163.367
R1517 B.n518 B.n145 163.367
R1518 B.n518 B.n143 163.367
R1519 B.n522 B.n143 163.367
R1520 B.n522 B.n137 163.367
R1521 B.n530 B.n137 163.367
R1522 B.n530 B.n135 163.367
R1523 B.n534 B.n135 163.367
R1524 B.n534 B.n129 163.367
R1525 B.n542 B.n129 163.367
R1526 B.n542 B.n127 163.367
R1527 B.n547 B.n127 163.367
R1528 B.n547 B.n121 163.367
R1529 B.n555 B.n121 163.367
R1530 B.n556 B.n555 163.367
R1531 B.n556 B.n5 163.367
R1532 B.n6 B.n5 163.367
R1533 B.n7 B.n6 163.367
R1534 B.n561 B.n7 163.367
R1535 B.n561 B.n12 163.367
R1536 B.n13 B.n12 163.367
R1537 B.n14 B.n13 163.367
R1538 B.n566 B.n14 163.367
R1539 B.n566 B.n19 163.367
R1540 B.n20 B.n19 163.367
R1541 B.n21 B.n20 163.367
R1542 B.n571 B.n21 163.367
R1543 B.n571 B.n26 163.367
R1544 B.n27 B.n26 163.367
R1545 B.n28 B.n27 163.367
R1546 B.n576 B.n28 163.367
R1547 B.n576 B.n33 163.367
R1548 B.n34 B.n33 163.367
R1549 B.n35 B.n34 163.367
R1550 B.n581 B.n35 163.367
R1551 B.n581 B.n40 163.367
R1552 B.n41 B.n40 163.367
R1553 B.n42 B.n41 163.367
R1554 B.n586 B.n42 163.367
R1555 B.n586 B.n47 163.367
R1556 B.n48 B.n47 163.367
R1557 B.n49 B.n48 163.367
R1558 B.n591 B.n49 163.367
R1559 B.n591 B.n54 163.367
R1560 B.n55 B.n54 163.367
R1561 B.n56 B.n55 163.367
R1562 B.n822 B.n820 163.367
R1563 B.n818 B.n60 163.367
R1564 B.n814 B.n812 163.367
R1565 B.n810 B.n62 163.367
R1566 B.n806 B.n804 163.367
R1567 B.n802 B.n64 163.367
R1568 B.n798 B.n796 163.367
R1569 B.n794 B.n66 163.367
R1570 B.n790 B.n788 163.367
R1571 B.n786 B.n68 163.367
R1572 B.n782 B.n780 163.367
R1573 B.n778 B.n70 163.367
R1574 B.n774 B.n772 163.367
R1575 B.n770 B.n72 163.367
R1576 B.n766 B.n764 163.367
R1577 B.n762 B.n74 163.367
R1578 B.n758 B.n756 163.367
R1579 B.n754 B.n76 163.367
R1580 B.n750 B.n748 163.367
R1581 B.n746 B.n78 163.367
R1582 B.n742 B.n740 163.367
R1583 B.n738 B.n80 163.367
R1584 B.n734 B.n732 163.367
R1585 B.n730 B.n82 163.367
R1586 B.n726 B.n724 163.367
R1587 B.n722 B.n84 163.367
R1588 B.n717 B.n715 163.367
R1589 B.n713 B.n88 163.367
R1590 B.n709 B.n707 163.367
R1591 B.n705 B.n90 163.367
R1592 B.n701 B.n699 163.367
R1593 B.n696 B.n695 163.367
R1594 B.n693 B.n96 163.367
R1595 B.n689 B.n687 163.367
R1596 B.n685 B.n98 163.367
R1597 B.n681 B.n679 163.367
R1598 B.n677 B.n100 163.367
R1599 B.n673 B.n671 163.367
R1600 B.n669 B.n102 163.367
R1601 B.n665 B.n663 163.367
R1602 B.n661 B.n104 163.367
R1603 B.n657 B.n655 163.367
R1604 B.n653 B.n106 163.367
R1605 B.n649 B.n647 163.367
R1606 B.n645 B.n108 163.367
R1607 B.n641 B.n639 163.367
R1608 B.n637 B.n110 163.367
R1609 B.n633 B.n631 163.367
R1610 B.n629 B.n112 163.367
R1611 B.n625 B.n623 163.367
R1612 B.n621 B.n114 163.367
R1613 B.n617 B.n615 163.367
R1614 B.n613 B.n116 163.367
R1615 B.n609 B.n607 163.367
R1616 B.n605 B.n118 163.367
R1617 B.n601 B.n599 163.367
R1618 B.n215 B.n214 72.3399
R1619 B.n207 B.n206 72.3399
R1620 B.n86 B.n85 72.3399
R1621 B.n92 B.n91 72.3399
R1622 B.n463 B.n179 71.676
R1623 B.n461 B.n181 71.676
R1624 B.n457 B.n456 71.676
R1625 B.n450 B.n183 71.676
R1626 B.n449 B.n448 71.676
R1627 B.n442 B.n185 71.676
R1628 B.n441 B.n440 71.676
R1629 B.n434 B.n187 71.676
R1630 B.n433 B.n432 71.676
R1631 B.n426 B.n189 71.676
R1632 B.n425 B.n424 71.676
R1633 B.n418 B.n191 71.676
R1634 B.n417 B.n416 71.676
R1635 B.n410 B.n193 71.676
R1636 B.n409 B.n408 71.676
R1637 B.n402 B.n195 71.676
R1638 B.n401 B.n400 71.676
R1639 B.n394 B.n197 71.676
R1640 B.n393 B.n392 71.676
R1641 B.n386 B.n199 71.676
R1642 B.n385 B.n384 71.676
R1643 B.n378 B.n201 71.676
R1644 B.n377 B.n376 71.676
R1645 B.n370 B.n203 71.676
R1646 B.n369 B.n368 71.676
R1647 B.n361 B.n205 71.676
R1648 B.n360 B.n359 71.676
R1649 B.n353 B.n209 71.676
R1650 B.n352 B.n351 71.676
R1651 B.n345 B.n211 71.676
R1652 B.n344 B.n343 71.676
R1653 B.n337 B.n213 71.676
R1654 B.n336 B.n335 71.676
R1655 B.n329 B.n218 71.676
R1656 B.n328 B.n327 71.676
R1657 B.n321 B.n220 71.676
R1658 B.n320 B.n319 71.676
R1659 B.n313 B.n222 71.676
R1660 B.n312 B.n311 71.676
R1661 B.n305 B.n224 71.676
R1662 B.n304 B.n303 71.676
R1663 B.n297 B.n226 71.676
R1664 B.n296 B.n295 71.676
R1665 B.n289 B.n228 71.676
R1666 B.n288 B.n287 71.676
R1667 B.n281 B.n230 71.676
R1668 B.n280 B.n279 71.676
R1669 B.n273 B.n232 71.676
R1670 B.n272 B.n271 71.676
R1671 B.n265 B.n234 71.676
R1672 B.n264 B.n263 71.676
R1673 B.n257 B.n236 71.676
R1674 B.n256 B.n255 71.676
R1675 B.n249 B.n238 71.676
R1676 B.n248 B.n247 71.676
R1677 B.n241 B.n240 71.676
R1678 B.n821 B.n58 71.676
R1679 B.n820 B.n819 71.676
R1680 B.n813 B.n60 71.676
R1681 B.n812 B.n811 71.676
R1682 B.n805 B.n62 71.676
R1683 B.n804 B.n803 71.676
R1684 B.n797 B.n64 71.676
R1685 B.n796 B.n795 71.676
R1686 B.n789 B.n66 71.676
R1687 B.n788 B.n787 71.676
R1688 B.n781 B.n68 71.676
R1689 B.n780 B.n779 71.676
R1690 B.n773 B.n70 71.676
R1691 B.n772 B.n771 71.676
R1692 B.n765 B.n72 71.676
R1693 B.n764 B.n763 71.676
R1694 B.n757 B.n74 71.676
R1695 B.n756 B.n755 71.676
R1696 B.n749 B.n76 71.676
R1697 B.n748 B.n747 71.676
R1698 B.n741 B.n78 71.676
R1699 B.n740 B.n739 71.676
R1700 B.n733 B.n80 71.676
R1701 B.n732 B.n731 71.676
R1702 B.n725 B.n82 71.676
R1703 B.n724 B.n723 71.676
R1704 B.n716 B.n84 71.676
R1705 B.n715 B.n714 71.676
R1706 B.n708 B.n88 71.676
R1707 B.n707 B.n706 71.676
R1708 B.n700 B.n90 71.676
R1709 B.n699 B.n94 71.676
R1710 B.n695 B.n694 71.676
R1711 B.n688 B.n96 71.676
R1712 B.n687 B.n686 71.676
R1713 B.n680 B.n98 71.676
R1714 B.n679 B.n678 71.676
R1715 B.n672 B.n100 71.676
R1716 B.n671 B.n670 71.676
R1717 B.n664 B.n102 71.676
R1718 B.n663 B.n662 71.676
R1719 B.n656 B.n104 71.676
R1720 B.n655 B.n654 71.676
R1721 B.n648 B.n106 71.676
R1722 B.n647 B.n646 71.676
R1723 B.n640 B.n108 71.676
R1724 B.n639 B.n638 71.676
R1725 B.n632 B.n110 71.676
R1726 B.n631 B.n630 71.676
R1727 B.n624 B.n112 71.676
R1728 B.n623 B.n622 71.676
R1729 B.n616 B.n114 71.676
R1730 B.n615 B.n614 71.676
R1731 B.n608 B.n116 71.676
R1732 B.n607 B.n606 71.676
R1733 B.n600 B.n118 71.676
R1734 B.n599 B.n598 71.676
R1735 B.n598 B.n597 71.676
R1736 B.n601 B.n600 71.676
R1737 B.n606 B.n605 71.676
R1738 B.n609 B.n608 71.676
R1739 B.n614 B.n613 71.676
R1740 B.n617 B.n616 71.676
R1741 B.n622 B.n621 71.676
R1742 B.n625 B.n624 71.676
R1743 B.n630 B.n629 71.676
R1744 B.n633 B.n632 71.676
R1745 B.n638 B.n637 71.676
R1746 B.n641 B.n640 71.676
R1747 B.n646 B.n645 71.676
R1748 B.n649 B.n648 71.676
R1749 B.n654 B.n653 71.676
R1750 B.n657 B.n656 71.676
R1751 B.n662 B.n661 71.676
R1752 B.n665 B.n664 71.676
R1753 B.n670 B.n669 71.676
R1754 B.n673 B.n672 71.676
R1755 B.n678 B.n677 71.676
R1756 B.n681 B.n680 71.676
R1757 B.n686 B.n685 71.676
R1758 B.n689 B.n688 71.676
R1759 B.n694 B.n693 71.676
R1760 B.n696 B.n94 71.676
R1761 B.n701 B.n700 71.676
R1762 B.n706 B.n705 71.676
R1763 B.n709 B.n708 71.676
R1764 B.n714 B.n713 71.676
R1765 B.n717 B.n716 71.676
R1766 B.n723 B.n722 71.676
R1767 B.n726 B.n725 71.676
R1768 B.n731 B.n730 71.676
R1769 B.n734 B.n733 71.676
R1770 B.n739 B.n738 71.676
R1771 B.n742 B.n741 71.676
R1772 B.n747 B.n746 71.676
R1773 B.n750 B.n749 71.676
R1774 B.n755 B.n754 71.676
R1775 B.n758 B.n757 71.676
R1776 B.n763 B.n762 71.676
R1777 B.n766 B.n765 71.676
R1778 B.n771 B.n770 71.676
R1779 B.n774 B.n773 71.676
R1780 B.n779 B.n778 71.676
R1781 B.n782 B.n781 71.676
R1782 B.n787 B.n786 71.676
R1783 B.n790 B.n789 71.676
R1784 B.n795 B.n794 71.676
R1785 B.n798 B.n797 71.676
R1786 B.n803 B.n802 71.676
R1787 B.n806 B.n805 71.676
R1788 B.n811 B.n810 71.676
R1789 B.n814 B.n813 71.676
R1790 B.n819 B.n818 71.676
R1791 B.n822 B.n821 71.676
R1792 B.n464 B.n463 71.676
R1793 B.n458 B.n181 71.676
R1794 B.n456 B.n455 71.676
R1795 B.n451 B.n450 71.676
R1796 B.n448 B.n447 71.676
R1797 B.n443 B.n442 71.676
R1798 B.n440 B.n439 71.676
R1799 B.n435 B.n434 71.676
R1800 B.n432 B.n431 71.676
R1801 B.n427 B.n426 71.676
R1802 B.n424 B.n423 71.676
R1803 B.n419 B.n418 71.676
R1804 B.n416 B.n415 71.676
R1805 B.n411 B.n410 71.676
R1806 B.n408 B.n407 71.676
R1807 B.n403 B.n402 71.676
R1808 B.n400 B.n399 71.676
R1809 B.n395 B.n394 71.676
R1810 B.n392 B.n391 71.676
R1811 B.n387 B.n386 71.676
R1812 B.n384 B.n383 71.676
R1813 B.n379 B.n378 71.676
R1814 B.n376 B.n375 71.676
R1815 B.n371 B.n370 71.676
R1816 B.n368 B.n367 71.676
R1817 B.n362 B.n361 71.676
R1818 B.n359 B.n358 71.676
R1819 B.n354 B.n353 71.676
R1820 B.n351 B.n350 71.676
R1821 B.n346 B.n345 71.676
R1822 B.n343 B.n342 71.676
R1823 B.n338 B.n337 71.676
R1824 B.n335 B.n334 71.676
R1825 B.n330 B.n329 71.676
R1826 B.n327 B.n326 71.676
R1827 B.n322 B.n321 71.676
R1828 B.n319 B.n318 71.676
R1829 B.n314 B.n313 71.676
R1830 B.n311 B.n310 71.676
R1831 B.n306 B.n305 71.676
R1832 B.n303 B.n302 71.676
R1833 B.n298 B.n297 71.676
R1834 B.n295 B.n294 71.676
R1835 B.n290 B.n289 71.676
R1836 B.n287 B.n286 71.676
R1837 B.n282 B.n281 71.676
R1838 B.n279 B.n278 71.676
R1839 B.n274 B.n273 71.676
R1840 B.n271 B.n270 71.676
R1841 B.n266 B.n265 71.676
R1842 B.n263 B.n262 71.676
R1843 B.n258 B.n257 71.676
R1844 B.n255 B.n254 71.676
R1845 B.n250 B.n249 71.676
R1846 B.n247 B.n246 71.676
R1847 B.n242 B.n241 71.676
R1848 B.n469 B.n178 66.9547
R1849 B.n827 B.n57 66.9547
R1850 B.n216 B.n215 59.5399
R1851 B.n364 B.n207 59.5399
R1852 B.n720 B.n86 59.5399
R1853 B.n93 B.n92 59.5399
R1854 B.n469 B.n174 35.85
R1855 B.n475 B.n174 35.85
R1856 B.n475 B.n170 35.85
R1857 B.n481 B.n170 35.85
R1858 B.n481 B.n166 35.85
R1859 B.n487 B.n166 35.85
R1860 B.n487 B.n162 35.85
R1861 B.n493 B.n162 35.85
R1862 B.n499 B.n158 35.85
R1863 B.n499 B.n154 35.85
R1864 B.n505 B.n154 35.85
R1865 B.n505 B.n150 35.85
R1866 B.n511 B.n150 35.85
R1867 B.n511 B.n146 35.85
R1868 B.n517 B.n146 35.85
R1869 B.n517 B.n142 35.85
R1870 B.n523 B.n142 35.85
R1871 B.n523 B.n138 35.85
R1872 B.n529 B.n138 35.85
R1873 B.n529 B.n134 35.85
R1874 B.n535 B.n134 35.85
R1875 B.n541 B.n130 35.85
R1876 B.n541 B.n126 35.85
R1877 B.n548 B.n126 35.85
R1878 B.n548 B.n122 35.85
R1879 B.n554 B.n122 35.85
R1880 B.n554 B.n4 35.85
R1881 B.n885 B.n4 35.85
R1882 B.n885 B.n884 35.85
R1883 B.n884 B.n883 35.85
R1884 B.n883 B.n8 35.85
R1885 B.n877 B.n8 35.85
R1886 B.n877 B.n876 35.85
R1887 B.n876 B.n875 35.85
R1888 B.n875 B.n15 35.85
R1889 B.n869 B.n868 35.85
R1890 B.n868 B.n867 35.85
R1891 B.n867 B.n22 35.85
R1892 B.n861 B.n22 35.85
R1893 B.n861 B.n860 35.85
R1894 B.n860 B.n859 35.85
R1895 B.n859 B.n29 35.85
R1896 B.n853 B.n29 35.85
R1897 B.n853 B.n852 35.85
R1898 B.n852 B.n851 35.85
R1899 B.n851 B.n36 35.85
R1900 B.n845 B.n36 35.85
R1901 B.n845 B.n844 35.85
R1902 B.n843 B.n43 35.85
R1903 B.n837 B.n43 35.85
R1904 B.n837 B.n836 35.85
R1905 B.n836 B.n835 35.85
R1906 B.n835 B.n50 35.85
R1907 B.n829 B.n50 35.85
R1908 B.n829 B.n828 35.85
R1909 B.n828 B.n827 35.85
R1910 B.n535 B.t1 32.6868
R1911 B.n869 B.t0 32.6868
R1912 B.n825 B.n824 32.6249
R1913 B.n596 B.n595 32.6249
R1914 B.n471 B.n176 32.6249
R1915 B.n467 B.n466 32.6249
R1916 B.n493 B.t3 26.3604
R1917 B.t7 B.n843 26.3604
R1918 B B.n887 18.0485
R1919 B.n824 B.n823 10.6151
R1920 B.n823 B.n59 10.6151
R1921 B.n817 B.n59 10.6151
R1922 B.n817 B.n816 10.6151
R1923 B.n816 B.n815 10.6151
R1924 B.n815 B.n61 10.6151
R1925 B.n809 B.n61 10.6151
R1926 B.n809 B.n808 10.6151
R1927 B.n808 B.n807 10.6151
R1928 B.n807 B.n63 10.6151
R1929 B.n801 B.n63 10.6151
R1930 B.n801 B.n800 10.6151
R1931 B.n800 B.n799 10.6151
R1932 B.n799 B.n65 10.6151
R1933 B.n793 B.n65 10.6151
R1934 B.n793 B.n792 10.6151
R1935 B.n792 B.n791 10.6151
R1936 B.n791 B.n67 10.6151
R1937 B.n785 B.n67 10.6151
R1938 B.n785 B.n784 10.6151
R1939 B.n784 B.n783 10.6151
R1940 B.n783 B.n69 10.6151
R1941 B.n777 B.n69 10.6151
R1942 B.n777 B.n776 10.6151
R1943 B.n776 B.n775 10.6151
R1944 B.n775 B.n71 10.6151
R1945 B.n769 B.n71 10.6151
R1946 B.n769 B.n768 10.6151
R1947 B.n768 B.n767 10.6151
R1948 B.n767 B.n73 10.6151
R1949 B.n761 B.n73 10.6151
R1950 B.n761 B.n760 10.6151
R1951 B.n760 B.n759 10.6151
R1952 B.n759 B.n75 10.6151
R1953 B.n753 B.n75 10.6151
R1954 B.n753 B.n752 10.6151
R1955 B.n752 B.n751 10.6151
R1956 B.n751 B.n77 10.6151
R1957 B.n745 B.n77 10.6151
R1958 B.n745 B.n744 10.6151
R1959 B.n744 B.n743 10.6151
R1960 B.n743 B.n79 10.6151
R1961 B.n737 B.n79 10.6151
R1962 B.n737 B.n736 10.6151
R1963 B.n736 B.n735 10.6151
R1964 B.n735 B.n81 10.6151
R1965 B.n729 B.n81 10.6151
R1966 B.n729 B.n728 10.6151
R1967 B.n728 B.n727 10.6151
R1968 B.n727 B.n83 10.6151
R1969 B.n721 B.n83 10.6151
R1970 B.n719 B.n718 10.6151
R1971 B.n718 B.n87 10.6151
R1972 B.n712 B.n87 10.6151
R1973 B.n712 B.n711 10.6151
R1974 B.n711 B.n710 10.6151
R1975 B.n710 B.n89 10.6151
R1976 B.n704 B.n89 10.6151
R1977 B.n704 B.n703 10.6151
R1978 B.n703 B.n702 10.6151
R1979 B.n698 B.n697 10.6151
R1980 B.n697 B.n95 10.6151
R1981 B.n692 B.n95 10.6151
R1982 B.n692 B.n691 10.6151
R1983 B.n691 B.n690 10.6151
R1984 B.n690 B.n97 10.6151
R1985 B.n684 B.n97 10.6151
R1986 B.n684 B.n683 10.6151
R1987 B.n683 B.n682 10.6151
R1988 B.n682 B.n99 10.6151
R1989 B.n676 B.n99 10.6151
R1990 B.n676 B.n675 10.6151
R1991 B.n675 B.n674 10.6151
R1992 B.n674 B.n101 10.6151
R1993 B.n668 B.n101 10.6151
R1994 B.n668 B.n667 10.6151
R1995 B.n667 B.n666 10.6151
R1996 B.n666 B.n103 10.6151
R1997 B.n660 B.n103 10.6151
R1998 B.n660 B.n659 10.6151
R1999 B.n659 B.n658 10.6151
R2000 B.n658 B.n105 10.6151
R2001 B.n652 B.n105 10.6151
R2002 B.n652 B.n651 10.6151
R2003 B.n651 B.n650 10.6151
R2004 B.n650 B.n107 10.6151
R2005 B.n644 B.n107 10.6151
R2006 B.n644 B.n643 10.6151
R2007 B.n643 B.n642 10.6151
R2008 B.n642 B.n109 10.6151
R2009 B.n636 B.n109 10.6151
R2010 B.n636 B.n635 10.6151
R2011 B.n635 B.n634 10.6151
R2012 B.n634 B.n111 10.6151
R2013 B.n628 B.n111 10.6151
R2014 B.n628 B.n627 10.6151
R2015 B.n627 B.n626 10.6151
R2016 B.n626 B.n113 10.6151
R2017 B.n620 B.n113 10.6151
R2018 B.n620 B.n619 10.6151
R2019 B.n619 B.n618 10.6151
R2020 B.n618 B.n115 10.6151
R2021 B.n612 B.n115 10.6151
R2022 B.n612 B.n611 10.6151
R2023 B.n611 B.n610 10.6151
R2024 B.n610 B.n117 10.6151
R2025 B.n604 B.n117 10.6151
R2026 B.n604 B.n603 10.6151
R2027 B.n603 B.n602 10.6151
R2028 B.n602 B.n119 10.6151
R2029 B.n596 B.n119 10.6151
R2030 B.n472 B.n471 10.6151
R2031 B.n473 B.n472 10.6151
R2032 B.n473 B.n168 10.6151
R2033 B.n483 B.n168 10.6151
R2034 B.n484 B.n483 10.6151
R2035 B.n485 B.n484 10.6151
R2036 B.n485 B.n160 10.6151
R2037 B.n495 B.n160 10.6151
R2038 B.n496 B.n495 10.6151
R2039 B.n497 B.n496 10.6151
R2040 B.n497 B.n152 10.6151
R2041 B.n507 B.n152 10.6151
R2042 B.n508 B.n507 10.6151
R2043 B.n509 B.n508 10.6151
R2044 B.n509 B.n144 10.6151
R2045 B.n519 B.n144 10.6151
R2046 B.n520 B.n519 10.6151
R2047 B.n521 B.n520 10.6151
R2048 B.n521 B.n136 10.6151
R2049 B.n531 B.n136 10.6151
R2050 B.n532 B.n531 10.6151
R2051 B.n533 B.n532 10.6151
R2052 B.n533 B.n128 10.6151
R2053 B.n543 B.n128 10.6151
R2054 B.n544 B.n543 10.6151
R2055 B.n546 B.n544 10.6151
R2056 B.n546 B.n545 10.6151
R2057 B.n545 B.n120 10.6151
R2058 B.n557 B.n120 10.6151
R2059 B.n558 B.n557 10.6151
R2060 B.n559 B.n558 10.6151
R2061 B.n560 B.n559 10.6151
R2062 B.n562 B.n560 10.6151
R2063 B.n563 B.n562 10.6151
R2064 B.n564 B.n563 10.6151
R2065 B.n565 B.n564 10.6151
R2066 B.n567 B.n565 10.6151
R2067 B.n568 B.n567 10.6151
R2068 B.n569 B.n568 10.6151
R2069 B.n570 B.n569 10.6151
R2070 B.n572 B.n570 10.6151
R2071 B.n573 B.n572 10.6151
R2072 B.n574 B.n573 10.6151
R2073 B.n575 B.n574 10.6151
R2074 B.n577 B.n575 10.6151
R2075 B.n578 B.n577 10.6151
R2076 B.n579 B.n578 10.6151
R2077 B.n580 B.n579 10.6151
R2078 B.n582 B.n580 10.6151
R2079 B.n583 B.n582 10.6151
R2080 B.n584 B.n583 10.6151
R2081 B.n585 B.n584 10.6151
R2082 B.n587 B.n585 10.6151
R2083 B.n588 B.n587 10.6151
R2084 B.n589 B.n588 10.6151
R2085 B.n590 B.n589 10.6151
R2086 B.n592 B.n590 10.6151
R2087 B.n593 B.n592 10.6151
R2088 B.n594 B.n593 10.6151
R2089 B.n595 B.n594 10.6151
R2090 B.n466 B.n465 10.6151
R2091 B.n465 B.n180 10.6151
R2092 B.n460 B.n180 10.6151
R2093 B.n460 B.n459 10.6151
R2094 B.n459 B.n182 10.6151
R2095 B.n454 B.n182 10.6151
R2096 B.n454 B.n453 10.6151
R2097 B.n453 B.n452 10.6151
R2098 B.n452 B.n184 10.6151
R2099 B.n446 B.n184 10.6151
R2100 B.n446 B.n445 10.6151
R2101 B.n445 B.n444 10.6151
R2102 B.n444 B.n186 10.6151
R2103 B.n438 B.n186 10.6151
R2104 B.n438 B.n437 10.6151
R2105 B.n437 B.n436 10.6151
R2106 B.n436 B.n188 10.6151
R2107 B.n430 B.n188 10.6151
R2108 B.n430 B.n429 10.6151
R2109 B.n429 B.n428 10.6151
R2110 B.n428 B.n190 10.6151
R2111 B.n422 B.n190 10.6151
R2112 B.n422 B.n421 10.6151
R2113 B.n421 B.n420 10.6151
R2114 B.n420 B.n192 10.6151
R2115 B.n414 B.n192 10.6151
R2116 B.n414 B.n413 10.6151
R2117 B.n413 B.n412 10.6151
R2118 B.n412 B.n194 10.6151
R2119 B.n406 B.n194 10.6151
R2120 B.n406 B.n405 10.6151
R2121 B.n405 B.n404 10.6151
R2122 B.n404 B.n196 10.6151
R2123 B.n398 B.n196 10.6151
R2124 B.n398 B.n397 10.6151
R2125 B.n397 B.n396 10.6151
R2126 B.n396 B.n198 10.6151
R2127 B.n390 B.n198 10.6151
R2128 B.n390 B.n389 10.6151
R2129 B.n389 B.n388 10.6151
R2130 B.n388 B.n200 10.6151
R2131 B.n382 B.n200 10.6151
R2132 B.n382 B.n381 10.6151
R2133 B.n381 B.n380 10.6151
R2134 B.n380 B.n202 10.6151
R2135 B.n374 B.n202 10.6151
R2136 B.n374 B.n373 10.6151
R2137 B.n373 B.n372 10.6151
R2138 B.n372 B.n204 10.6151
R2139 B.n366 B.n204 10.6151
R2140 B.n366 B.n365 10.6151
R2141 B.n363 B.n208 10.6151
R2142 B.n357 B.n208 10.6151
R2143 B.n357 B.n356 10.6151
R2144 B.n356 B.n355 10.6151
R2145 B.n355 B.n210 10.6151
R2146 B.n349 B.n210 10.6151
R2147 B.n349 B.n348 10.6151
R2148 B.n348 B.n347 10.6151
R2149 B.n347 B.n212 10.6151
R2150 B.n341 B.n340 10.6151
R2151 B.n340 B.n339 10.6151
R2152 B.n339 B.n217 10.6151
R2153 B.n333 B.n217 10.6151
R2154 B.n333 B.n332 10.6151
R2155 B.n332 B.n331 10.6151
R2156 B.n331 B.n219 10.6151
R2157 B.n325 B.n219 10.6151
R2158 B.n325 B.n324 10.6151
R2159 B.n324 B.n323 10.6151
R2160 B.n323 B.n221 10.6151
R2161 B.n317 B.n221 10.6151
R2162 B.n317 B.n316 10.6151
R2163 B.n316 B.n315 10.6151
R2164 B.n315 B.n223 10.6151
R2165 B.n309 B.n223 10.6151
R2166 B.n309 B.n308 10.6151
R2167 B.n308 B.n307 10.6151
R2168 B.n307 B.n225 10.6151
R2169 B.n301 B.n225 10.6151
R2170 B.n301 B.n300 10.6151
R2171 B.n300 B.n299 10.6151
R2172 B.n299 B.n227 10.6151
R2173 B.n293 B.n227 10.6151
R2174 B.n293 B.n292 10.6151
R2175 B.n292 B.n291 10.6151
R2176 B.n291 B.n229 10.6151
R2177 B.n285 B.n229 10.6151
R2178 B.n285 B.n284 10.6151
R2179 B.n284 B.n283 10.6151
R2180 B.n283 B.n231 10.6151
R2181 B.n277 B.n231 10.6151
R2182 B.n277 B.n276 10.6151
R2183 B.n276 B.n275 10.6151
R2184 B.n275 B.n233 10.6151
R2185 B.n269 B.n233 10.6151
R2186 B.n269 B.n268 10.6151
R2187 B.n268 B.n267 10.6151
R2188 B.n267 B.n235 10.6151
R2189 B.n261 B.n235 10.6151
R2190 B.n261 B.n260 10.6151
R2191 B.n260 B.n259 10.6151
R2192 B.n259 B.n237 10.6151
R2193 B.n253 B.n237 10.6151
R2194 B.n253 B.n252 10.6151
R2195 B.n252 B.n251 10.6151
R2196 B.n251 B.n239 10.6151
R2197 B.n245 B.n239 10.6151
R2198 B.n245 B.n244 10.6151
R2199 B.n244 B.n243 10.6151
R2200 B.n243 B.n176 10.6151
R2201 B.n467 B.n172 10.6151
R2202 B.n477 B.n172 10.6151
R2203 B.n478 B.n477 10.6151
R2204 B.n479 B.n478 10.6151
R2205 B.n479 B.n164 10.6151
R2206 B.n489 B.n164 10.6151
R2207 B.n490 B.n489 10.6151
R2208 B.n491 B.n490 10.6151
R2209 B.n491 B.n156 10.6151
R2210 B.n501 B.n156 10.6151
R2211 B.n502 B.n501 10.6151
R2212 B.n503 B.n502 10.6151
R2213 B.n503 B.n148 10.6151
R2214 B.n513 B.n148 10.6151
R2215 B.n514 B.n513 10.6151
R2216 B.n515 B.n514 10.6151
R2217 B.n515 B.n140 10.6151
R2218 B.n525 B.n140 10.6151
R2219 B.n526 B.n525 10.6151
R2220 B.n527 B.n526 10.6151
R2221 B.n527 B.n132 10.6151
R2222 B.n537 B.n132 10.6151
R2223 B.n538 B.n537 10.6151
R2224 B.n539 B.n538 10.6151
R2225 B.n539 B.n124 10.6151
R2226 B.n550 B.n124 10.6151
R2227 B.n551 B.n550 10.6151
R2228 B.n552 B.n551 10.6151
R2229 B.n552 B.n0 10.6151
R2230 B.n881 B.n1 10.6151
R2231 B.n881 B.n880 10.6151
R2232 B.n880 B.n879 10.6151
R2233 B.n879 B.n10 10.6151
R2234 B.n873 B.n10 10.6151
R2235 B.n873 B.n872 10.6151
R2236 B.n872 B.n871 10.6151
R2237 B.n871 B.n17 10.6151
R2238 B.n865 B.n17 10.6151
R2239 B.n865 B.n864 10.6151
R2240 B.n864 B.n863 10.6151
R2241 B.n863 B.n24 10.6151
R2242 B.n857 B.n24 10.6151
R2243 B.n857 B.n856 10.6151
R2244 B.n856 B.n855 10.6151
R2245 B.n855 B.n31 10.6151
R2246 B.n849 B.n31 10.6151
R2247 B.n849 B.n848 10.6151
R2248 B.n848 B.n847 10.6151
R2249 B.n847 B.n38 10.6151
R2250 B.n841 B.n38 10.6151
R2251 B.n841 B.n840 10.6151
R2252 B.n840 B.n839 10.6151
R2253 B.n839 B.n45 10.6151
R2254 B.n833 B.n45 10.6151
R2255 B.n833 B.n832 10.6151
R2256 B.n832 B.n831 10.6151
R2257 B.n831 B.n52 10.6151
R2258 B.n825 B.n52 10.6151
R2259 B.t3 B.n158 9.49008
R2260 B.n844 B.t7 9.49008
R2261 B.n721 B.n720 9.36635
R2262 B.n698 B.n93 9.36635
R2263 B.n365 B.n364 9.36635
R2264 B.n341 B.n216 9.36635
R2265 B.t1 B.n130 3.16369
R2266 B.t0 B.n15 3.16369
R2267 B.n887 B.n0 2.81026
R2268 B.n887 B.n1 2.81026
R2269 B.n720 B.n719 1.24928
R2270 B.n702 B.n93 1.24928
R2271 B.n364 B.n363 1.24928
R2272 B.n216 B.n212 1.24928
R2273 VN VN.t1 198.698
R2274 VN VN.t0 149.82
R2275 VDD2.n165 VDD2.n85 289.615
R2276 VDD2.n80 VDD2.n0 289.615
R2277 VDD2.n166 VDD2.n165 185
R2278 VDD2.n164 VDD2.n163 185
R2279 VDD2.n89 VDD2.n88 185
R2280 VDD2.n93 VDD2.n91 185
R2281 VDD2.n158 VDD2.n157 185
R2282 VDD2.n156 VDD2.n155 185
R2283 VDD2.n95 VDD2.n94 185
R2284 VDD2.n150 VDD2.n149 185
R2285 VDD2.n148 VDD2.n147 185
R2286 VDD2.n99 VDD2.n98 185
R2287 VDD2.n142 VDD2.n141 185
R2288 VDD2.n140 VDD2.n139 185
R2289 VDD2.n103 VDD2.n102 185
R2290 VDD2.n134 VDD2.n133 185
R2291 VDD2.n132 VDD2.n131 185
R2292 VDD2.n107 VDD2.n106 185
R2293 VDD2.n126 VDD2.n125 185
R2294 VDD2.n124 VDD2.n123 185
R2295 VDD2.n111 VDD2.n110 185
R2296 VDD2.n118 VDD2.n117 185
R2297 VDD2.n116 VDD2.n115 185
R2298 VDD2.n29 VDD2.n28 185
R2299 VDD2.n31 VDD2.n30 185
R2300 VDD2.n24 VDD2.n23 185
R2301 VDD2.n37 VDD2.n36 185
R2302 VDD2.n39 VDD2.n38 185
R2303 VDD2.n20 VDD2.n19 185
R2304 VDD2.n45 VDD2.n44 185
R2305 VDD2.n47 VDD2.n46 185
R2306 VDD2.n16 VDD2.n15 185
R2307 VDD2.n53 VDD2.n52 185
R2308 VDD2.n55 VDD2.n54 185
R2309 VDD2.n12 VDD2.n11 185
R2310 VDD2.n61 VDD2.n60 185
R2311 VDD2.n63 VDD2.n62 185
R2312 VDD2.n8 VDD2.n7 185
R2313 VDD2.n70 VDD2.n69 185
R2314 VDD2.n71 VDD2.n6 185
R2315 VDD2.n73 VDD2.n72 185
R2316 VDD2.n4 VDD2.n3 185
R2317 VDD2.n79 VDD2.n78 185
R2318 VDD2.n81 VDD2.n80 185
R2319 VDD2.n114 VDD2.t0 147.659
R2320 VDD2.n27 VDD2.t1 147.659
R2321 VDD2.n165 VDD2.n164 104.615
R2322 VDD2.n164 VDD2.n88 104.615
R2323 VDD2.n93 VDD2.n88 104.615
R2324 VDD2.n157 VDD2.n93 104.615
R2325 VDD2.n157 VDD2.n156 104.615
R2326 VDD2.n156 VDD2.n94 104.615
R2327 VDD2.n149 VDD2.n94 104.615
R2328 VDD2.n149 VDD2.n148 104.615
R2329 VDD2.n148 VDD2.n98 104.615
R2330 VDD2.n141 VDD2.n98 104.615
R2331 VDD2.n141 VDD2.n140 104.615
R2332 VDD2.n140 VDD2.n102 104.615
R2333 VDD2.n133 VDD2.n102 104.615
R2334 VDD2.n133 VDD2.n132 104.615
R2335 VDD2.n132 VDD2.n106 104.615
R2336 VDD2.n125 VDD2.n106 104.615
R2337 VDD2.n125 VDD2.n124 104.615
R2338 VDD2.n124 VDD2.n110 104.615
R2339 VDD2.n117 VDD2.n110 104.615
R2340 VDD2.n117 VDD2.n116 104.615
R2341 VDD2.n30 VDD2.n29 104.615
R2342 VDD2.n30 VDD2.n23 104.615
R2343 VDD2.n37 VDD2.n23 104.615
R2344 VDD2.n38 VDD2.n37 104.615
R2345 VDD2.n38 VDD2.n19 104.615
R2346 VDD2.n45 VDD2.n19 104.615
R2347 VDD2.n46 VDD2.n45 104.615
R2348 VDD2.n46 VDD2.n15 104.615
R2349 VDD2.n53 VDD2.n15 104.615
R2350 VDD2.n54 VDD2.n53 104.615
R2351 VDD2.n54 VDD2.n11 104.615
R2352 VDD2.n61 VDD2.n11 104.615
R2353 VDD2.n62 VDD2.n61 104.615
R2354 VDD2.n62 VDD2.n7 104.615
R2355 VDD2.n70 VDD2.n7 104.615
R2356 VDD2.n71 VDD2.n70 104.615
R2357 VDD2.n72 VDD2.n71 104.615
R2358 VDD2.n72 VDD2.n3 104.615
R2359 VDD2.n79 VDD2.n3 104.615
R2360 VDD2.n80 VDD2.n79 104.615
R2361 VDD2.n170 VDD2.n84 96.8549
R2362 VDD2.n170 VDD2.n169 53.3247
R2363 VDD2.n116 VDD2.t0 52.3082
R2364 VDD2.n29 VDD2.t1 52.3082
R2365 VDD2.n115 VDD2.n114 15.6677
R2366 VDD2.n28 VDD2.n27 15.6677
R2367 VDD2.n91 VDD2.n89 13.1884
R2368 VDD2.n73 VDD2.n4 13.1884
R2369 VDD2.n163 VDD2.n162 12.8005
R2370 VDD2.n159 VDD2.n158 12.8005
R2371 VDD2.n118 VDD2.n113 12.8005
R2372 VDD2.n31 VDD2.n26 12.8005
R2373 VDD2.n74 VDD2.n6 12.8005
R2374 VDD2.n78 VDD2.n77 12.8005
R2375 VDD2.n166 VDD2.n87 12.0247
R2376 VDD2.n155 VDD2.n92 12.0247
R2377 VDD2.n119 VDD2.n111 12.0247
R2378 VDD2.n32 VDD2.n24 12.0247
R2379 VDD2.n69 VDD2.n68 12.0247
R2380 VDD2.n81 VDD2.n2 12.0247
R2381 VDD2.n167 VDD2.n85 11.249
R2382 VDD2.n154 VDD2.n95 11.249
R2383 VDD2.n123 VDD2.n122 11.249
R2384 VDD2.n36 VDD2.n35 11.249
R2385 VDD2.n67 VDD2.n8 11.249
R2386 VDD2.n82 VDD2.n0 11.249
R2387 VDD2.n151 VDD2.n150 10.4732
R2388 VDD2.n126 VDD2.n109 10.4732
R2389 VDD2.n39 VDD2.n22 10.4732
R2390 VDD2.n64 VDD2.n63 10.4732
R2391 VDD2.n147 VDD2.n97 9.69747
R2392 VDD2.n127 VDD2.n107 9.69747
R2393 VDD2.n40 VDD2.n20 9.69747
R2394 VDD2.n60 VDD2.n10 9.69747
R2395 VDD2.n169 VDD2.n168 9.45567
R2396 VDD2.n84 VDD2.n83 9.45567
R2397 VDD2.n101 VDD2.n100 9.3005
R2398 VDD2.n144 VDD2.n143 9.3005
R2399 VDD2.n146 VDD2.n145 9.3005
R2400 VDD2.n97 VDD2.n96 9.3005
R2401 VDD2.n152 VDD2.n151 9.3005
R2402 VDD2.n154 VDD2.n153 9.3005
R2403 VDD2.n92 VDD2.n90 9.3005
R2404 VDD2.n160 VDD2.n159 9.3005
R2405 VDD2.n168 VDD2.n167 9.3005
R2406 VDD2.n87 VDD2.n86 9.3005
R2407 VDD2.n162 VDD2.n161 9.3005
R2408 VDD2.n138 VDD2.n137 9.3005
R2409 VDD2.n136 VDD2.n135 9.3005
R2410 VDD2.n105 VDD2.n104 9.3005
R2411 VDD2.n130 VDD2.n129 9.3005
R2412 VDD2.n128 VDD2.n127 9.3005
R2413 VDD2.n109 VDD2.n108 9.3005
R2414 VDD2.n122 VDD2.n121 9.3005
R2415 VDD2.n120 VDD2.n119 9.3005
R2416 VDD2.n113 VDD2.n112 9.3005
R2417 VDD2.n83 VDD2.n82 9.3005
R2418 VDD2.n2 VDD2.n1 9.3005
R2419 VDD2.n77 VDD2.n76 9.3005
R2420 VDD2.n49 VDD2.n48 9.3005
R2421 VDD2.n18 VDD2.n17 9.3005
R2422 VDD2.n43 VDD2.n42 9.3005
R2423 VDD2.n41 VDD2.n40 9.3005
R2424 VDD2.n22 VDD2.n21 9.3005
R2425 VDD2.n35 VDD2.n34 9.3005
R2426 VDD2.n33 VDD2.n32 9.3005
R2427 VDD2.n26 VDD2.n25 9.3005
R2428 VDD2.n51 VDD2.n50 9.3005
R2429 VDD2.n14 VDD2.n13 9.3005
R2430 VDD2.n57 VDD2.n56 9.3005
R2431 VDD2.n59 VDD2.n58 9.3005
R2432 VDD2.n10 VDD2.n9 9.3005
R2433 VDD2.n65 VDD2.n64 9.3005
R2434 VDD2.n67 VDD2.n66 9.3005
R2435 VDD2.n68 VDD2.n5 9.3005
R2436 VDD2.n75 VDD2.n74 9.3005
R2437 VDD2.n146 VDD2.n99 8.92171
R2438 VDD2.n131 VDD2.n130 8.92171
R2439 VDD2.n44 VDD2.n43 8.92171
R2440 VDD2.n59 VDD2.n12 8.92171
R2441 VDD2.n143 VDD2.n142 8.14595
R2442 VDD2.n134 VDD2.n105 8.14595
R2443 VDD2.n47 VDD2.n18 8.14595
R2444 VDD2.n56 VDD2.n55 8.14595
R2445 VDD2.n139 VDD2.n101 7.3702
R2446 VDD2.n135 VDD2.n103 7.3702
R2447 VDD2.n48 VDD2.n16 7.3702
R2448 VDD2.n52 VDD2.n14 7.3702
R2449 VDD2.n139 VDD2.n138 6.59444
R2450 VDD2.n138 VDD2.n103 6.59444
R2451 VDD2.n51 VDD2.n16 6.59444
R2452 VDD2.n52 VDD2.n51 6.59444
R2453 VDD2.n142 VDD2.n101 5.81868
R2454 VDD2.n135 VDD2.n134 5.81868
R2455 VDD2.n48 VDD2.n47 5.81868
R2456 VDD2.n55 VDD2.n14 5.81868
R2457 VDD2.n143 VDD2.n99 5.04292
R2458 VDD2.n131 VDD2.n105 5.04292
R2459 VDD2.n44 VDD2.n18 5.04292
R2460 VDD2.n56 VDD2.n12 5.04292
R2461 VDD2.n114 VDD2.n112 4.38563
R2462 VDD2.n27 VDD2.n25 4.38563
R2463 VDD2.n147 VDD2.n146 4.26717
R2464 VDD2.n130 VDD2.n107 4.26717
R2465 VDD2.n43 VDD2.n20 4.26717
R2466 VDD2.n60 VDD2.n59 4.26717
R2467 VDD2.n150 VDD2.n97 3.49141
R2468 VDD2.n127 VDD2.n126 3.49141
R2469 VDD2.n40 VDD2.n39 3.49141
R2470 VDD2.n63 VDD2.n10 3.49141
R2471 VDD2.n169 VDD2.n85 2.71565
R2472 VDD2.n151 VDD2.n95 2.71565
R2473 VDD2.n123 VDD2.n109 2.71565
R2474 VDD2.n36 VDD2.n22 2.71565
R2475 VDD2.n64 VDD2.n8 2.71565
R2476 VDD2.n84 VDD2.n0 2.71565
R2477 VDD2.n167 VDD2.n166 1.93989
R2478 VDD2.n155 VDD2.n154 1.93989
R2479 VDD2.n122 VDD2.n111 1.93989
R2480 VDD2.n35 VDD2.n24 1.93989
R2481 VDD2.n69 VDD2.n67 1.93989
R2482 VDD2.n82 VDD2.n81 1.93989
R2483 VDD2.n163 VDD2.n87 1.16414
R2484 VDD2.n158 VDD2.n92 1.16414
R2485 VDD2.n119 VDD2.n118 1.16414
R2486 VDD2.n32 VDD2.n31 1.16414
R2487 VDD2.n68 VDD2.n6 1.16414
R2488 VDD2.n78 VDD2.n2 1.16414
R2489 VDD2 VDD2.n170 0.862569
R2490 VDD2.n162 VDD2.n89 0.388379
R2491 VDD2.n159 VDD2.n91 0.388379
R2492 VDD2.n115 VDD2.n113 0.388379
R2493 VDD2.n28 VDD2.n26 0.388379
R2494 VDD2.n74 VDD2.n73 0.388379
R2495 VDD2.n77 VDD2.n4 0.388379
R2496 VDD2.n168 VDD2.n86 0.155672
R2497 VDD2.n161 VDD2.n86 0.155672
R2498 VDD2.n161 VDD2.n160 0.155672
R2499 VDD2.n160 VDD2.n90 0.155672
R2500 VDD2.n153 VDD2.n90 0.155672
R2501 VDD2.n153 VDD2.n152 0.155672
R2502 VDD2.n152 VDD2.n96 0.155672
R2503 VDD2.n145 VDD2.n96 0.155672
R2504 VDD2.n145 VDD2.n144 0.155672
R2505 VDD2.n144 VDD2.n100 0.155672
R2506 VDD2.n137 VDD2.n100 0.155672
R2507 VDD2.n137 VDD2.n136 0.155672
R2508 VDD2.n136 VDD2.n104 0.155672
R2509 VDD2.n129 VDD2.n104 0.155672
R2510 VDD2.n129 VDD2.n128 0.155672
R2511 VDD2.n128 VDD2.n108 0.155672
R2512 VDD2.n121 VDD2.n108 0.155672
R2513 VDD2.n121 VDD2.n120 0.155672
R2514 VDD2.n120 VDD2.n112 0.155672
R2515 VDD2.n33 VDD2.n25 0.155672
R2516 VDD2.n34 VDD2.n33 0.155672
R2517 VDD2.n34 VDD2.n21 0.155672
R2518 VDD2.n41 VDD2.n21 0.155672
R2519 VDD2.n42 VDD2.n41 0.155672
R2520 VDD2.n42 VDD2.n17 0.155672
R2521 VDD2.n49 VDD2.n17 0.155672
R2522 VDD2.n50 VDD2.n49 0.155672
R2523 VDD2.n50 VDD2.n13 0.155672
R2524 VDD2.n57 VDD2.n13 0.155672
R2525 VDD2.n58 VDD2.n57 0.155672
R2526 VDD2.n58 VDD2.n9 0.155672
R2527 VDD2.n65 VDD2.n9 0.155672
R2528 VDD2.n66 VDD2.n65 0.155672
R2529 VDD2.n66 VDD2.n5 0.155672
R2530 VDD2.n75 VDD2.n5 0.155672
R2531 VDD2.n76 VDD2.n75 0.155672
R2532 VDD2.n76 VDD2.n1 0.155672
R2533 VDD2.n83 VDD2.n1 0.155672
C0 VDD1 VDD2 0.772565f
C1 VP VDD1 3.88633f
C2 VN VDD1 0.148489f
C3 VP VDD2 0.366907f
C4 VN VDD2 3.67061f
C5 VTAIL VDD1 6.12527f
C6 VP VN 6.49627f
C7 VTAIL VDD2 6.18132f
C8 VP VTAIL 3.23484f
C9 VN VTAIL 3.22056f
C10 VDD2 B 5.352203f
C11 VDD1 B 8.54216f
C12 VTAIL B 9.218194f
C13 VN B 12.32251f
C14 VP B 7.632671f
C15 VDD2.n0 B 0.029399f
C16 VDD2.n1 B 0.020235f
C17 VDD2.n2 B 0.010874f
C18 VDD2.n3 B 0.025701f
C19 VDD2.n4 B 0.011193f
C20 VDD2.n5 B 0.020235f
C21 VDD2.n6 B 0.011513f
C22 VDD2.n7 B 0.025701f
C23 VDD2.n8 B 0.011513f
C24 VDD2.n9 B 0.020235f
C25 VDD2.n10 B 0.010874f
C26 VDD2.n11 B 0.025701f
C27 VDD2.n12 B 0.011513f
C28 VDD2.n13 B 0.020235f
C29 VDD2.n14 B 0.010874f
C30 VDD2.n15 B 0.025701f
C31 VDD2.n16 B 0.011513f
C32 VDD2.n17 B 0.020235f
C33 VDD2.n18 B 0.010874f
C34 VDD2.n19 B 0.025701f
C35 VDD2.n20 B 0.011513f
C36 VDD2.n21 B 0.020235f
C37 VDD2.n22 B 0.010874f
C38 VDD2.n23 B 0.025701f
C39 VDD2.n24 B 0.011513f
C40 VDD2.n25 B 1.37127f
C41 VDD2.n26 B 0.010874f
C42 VDD2.t1 B 0.04242f
C43 VDD2.n27 B 0.134974f
C44 VDD2.n28 B 0.015183f
C45 VDD2.n29 B 0.019276f
C46 VDD2.n30 B 0.025701f
C47 VDD2.n31 B 0.011513f
C48 VDD2.n32 B 0.010874f
C49 VDD2.n33 B 0.020235f
C50 VDD2.n34 B 0.020235f
C51 VDD2.n35 B 0.010874f
C52 VDD2.n36 B 0.011513f
C53 VDD2.n37 B 0.025701f
C54 VDD2.n38 B 0.025701f
C55 VDD2.n39 B 0.011513f
C56 VDD2.n40 B 0.010874f
C57 VDD2.n41 B 0.020235f
C58 VDD2.n42 B 0.020235f
C59 VDD2.n43 B 0.010874f
C60 VDD2.n44 B 0.011513f
C61 VDD2.n45 B 0.025701f
C62 VDD2.n46 B 0.025701f
C63 VDD2.n47 B 0.011513f
C64 VDD2.n48 B 0.010874f
C65 VDD2.n49 B 0.020235f
C66 VDD2.n50 B 0.020235f
C67 VDD2.n51 B 0.010874f
C68 VDD2.n52 B 0.011513f
C69 VDD2.n53 B 0.025701f
C70 VDD2.n54 B 0.025701f
C71 VDD2.n55 B 0.011513f
C72 VDD2.n56 B 0.010874f
C73 VDD2.n57 B 0.020235f
C74 VDD2.n58 B 0.020235f
C75 VDD2.n59 B 0.010874f
C76 VDD2.n60 B 0.011513f
C77 VDD2.n61 B 0.025701f
C78 VDD2.n62 B 0.025701f
C79 VDD2.n63 B 0.011513f
C80 VDD2.n64 B 0.010874f
C81 VDD2.n65 B 0.020235f
C82 VDD2.n66 B 0.020235f
C83 VDD2.n67 B 0.010874f
C84 VDD2.n68 B 0.010874f
C85 VDD2.n69 B 0.011513f
C86 VDD2.n70 B 0.025701f
C87 VDD2.n71 B 0.025701f
C88 VDD2.n72 B 0.025701f
C89 VDD2.n73 B 0.011193f
C90 VDD2.n74 B 0.010874f
C91 VDD2.n75 B 0.020235f
C92 VDD2.n76 B 0.020235f
C93 VDD2.n77 B 0.010874f
C94 VDD2.n78 B 0.011513f
C95 VDD2.n79 B 0.025701f
C96 VDD2.n80 B 0.057329f
C97 VDD2.n81 B 0.011513f
C98 VDD2.n82 B 0.010874f
C99 VDD2.n83 B 0.053131f
C100 VDD2.n84 B 0.717063f
C101 VDD2.n85 B 0.029399f
C102 VDD2.n86 B 0.020235f
C103 VDD2.n87 B 0.010874f
C104 VDD2.n88 B 0.025701f
C105 VDD2.n89 B 0.011193f
C106 VDD2.n90 B 0.020235f
C107 VDD2.n91 B 0.011193f
C108 VDD2.n92 B 0.010874f
C109 VDD2.n93 B 0.025701f
C110 VDD2.n94 B 0.025701f
C111 VDD2.n95 B 0.011513f
C112 VDD2.n96 B 0.020235f
C113 VDD2.n97 B 0.010874f
C114 VDD2.n98 B 0.025701f
C115 VDD2.n99 B 0.011513f
C116 VDD2.n100 B 0.020235f
C117 VDD2.n101 B 0.010874f
C118 VDD2.n102 B 0.025701f
C119 VDD2.n103 B 0.011513f
C120 VDD2.n104 B 0.020235f
C121 VDD2.n105 B 0.010874f
C122 VDD2.n106 B 0.025701f
C123 VDD2.n107 B 0.011513f
C124 VDD2.n108 B 0.020235f
C125 VDD2.n109 B 0.010874f
C126 VDD2.n110 B 0.025701f
C127 VDD2.n111 B 0.011513f
C128 VDD2.n112 B 1.37127f
C129 VDD2.n113 B 0.010874f
C130 VDD2.t0 B 0.04242f
C131 VDD2.n114 B 0.134974f
C132 VDD2.n115 B 0.015183f
C133 VDD2.n116 B 0.019276f
C134 VDD2.n117 B 0.025701f
C135 VDD2.n118 B 0.011513f
C136 VDD2.n119 B 0.010874f
C137 VDD2.n120 B 0.020235f
C138 VDD2.n121 B 0.020235f
C139 VDD2.n122 B 0.010874f
C140 VDD2.n123 B 0.011513f
C141 VDD2.n124 B 0.025701f
C142 VDD2.n125 B 0.025701f
C143 VDD2.n126 B 0.011513f
C144 VDD2.n127 B 0.010874f
C145 VDD2.n128 B 0.020235f
C146 VDD2.n129 B 0.020235f
C147 VDD2.n130 B 0.010874f
C148 VDD2.n131 B 0.011513f
C149 VDD2.n132 B 0.025701f
C150 VDD2.n133 B 0.025701f
C151 VDD2.n134 B 0.011513f
C152 VDD2.n135 B 0.010874f
C153 VDD2.n136 B 0.020235f
C154 VDD2.n137 B 0.020235f
C155 VDD2.n138 B 0.010874f
C156 VDD2.n139 B 0.011513f
C157 VDD2.n140 B 0.025701f
C158 VDD2.n141 B 0.025701f
C159 VDD2.n142 B 0.011513f
C160 VDD2.n143 B 0.010874f
C161 VDD2.n144 B 0.020235f
C162 VDD2.n145 B 0.020235f
C163 VDD2.n146 B 0.010874f
C164 VDD2.n147 B 0.011513f
C165 VDD2.n148 B 0.025701f
C166 VDD2.n149 B 0.025701f
C167 VDD2.n150 B 0.011513f
C168 VDD2.n151 B 0.010874f
C169 VDD2.n152 B 0.020235f
C170 VDD2.n153 B 0.020235f
C171 VDD2.n154 B 0.010874f
C172 VDD2.n155 B 0.011513f
C173 VDD2.n156 B 0.025701f
C174 VDD2.n157 B 0.025701f
C175 VDD2.n158 B 0.011513f
C176 VDD2.n159 B 0.010874f
C177 VDD2.n160 B 0.020235f
C178 VDD2.n161 B 0.020235f
C179 VDD2.n162 B 0.010874f
C180 VDD2.n163 B 0.011513f
C181 VDD2.n164 B 0.025701f
C182 VDD2.n165 B 0.057329f
C183 VDD2.n166 B 0.011513f
C184 VDD2.n167 B 0.010874f
C185 VDD2.n168 B 0.053131f
C186 VDD2.n169 B 0.046365f
C187 VDD2.n170 B 2.92968f
C188 VN.t0 B 4.04916f
C189 VN.t1 B 4.69897f
C190 VDD1.n0 B 0.029473f
C191 VDD1.n1 B 0.020287f
C192 VDD1.n2 B 0.010901f
C193 VDD1.n3 B 0.025767f
C194 VDD1.n4 B 0.011222f
C195 VDD1.n5 B 0.020287f
C196 VDD1.n6 B 0.011222f
C197 VDD1.n7 B 0.010901f
C198 VDD1.n8 B 0.025767f
C199 VDD1.n9 B 0.025767f
C200 VDD1.n10 B 0.011542f
C201 VDD1.n11 B 0.020287f
C202 VDD1.n12 B 0.010901f
C203 VDD1.n13 B 0.025767f
C204 VDD1.n14 B 0.011542f
C205 VDD1.n15 B 0.020287f
C206 VDD1.n16 B 0.010901f
C207 VDD1.n17 B 0.025767f
C208 VDD1.n18 B 0.011542f
C209 VDD1.n19 B 0.020287f
C210 VDD1.n20 B 0.010901f
C211 VDD1.n21 B 0.025767f
C212 VDD1.n22 B 0.011542f
C213 VDD1.n23 B 0.020287f
C214 VDD1.n24 B 0.010901f
C215 VDD1.n25 B 0.025767f
C216 VDD1.n26 B 0.011542f
C217 VDD1.n27 B 1.37474f
C218 VDD1.n28 B 0.010901f
C219 VDD1.t0 B 0.042527f
C220 VDD1.n29 B 0.135315f
C221 VDD1.n30 B 0.015221f
C222 VDD1.n31 B 0.019325f
C223 VDD1.n32 B 0.025767f
C224 VDD1.n33 B 0.011542f
C225 VDD1.n34 B 0.010901f
C226 VDD1.n35 B 0.020287f
C227 VDD1.n36 B 0.020287f
C228 VDD1.n37 B 0.010901f
C229 VDD1.n38 B 0.011542f
C230 VDD1.n39 B 0.025767f
C231 VDD1.n40 B 0.025767f
C232 VDD1.n41 B 0.011542f
C233 VDD1.n42 B 0.010901f
C234 VDD1.n43 B 0.020287f
C235 VDD1.n44 B 0.020287f
C236 VDD1.n45 B 0.010901f
C237 VDD1.n46 B 0.011542f
C238 VDD1.n47 B 0.025767f
C239 VDD1.n48 B 0.025767f
C240 VDD1.n49 B 0.011542f
C241 VDD1.n50 B 0.010901f
C242 VDD1.n51 B 0.020287f
C243 VDD1.n52 B 0.020287f
C244 VDD1.n53 B 0.010901f
C245 VDD1.n54 B 0.011542f
C246 VDD1.n55 B 0.025767f
C247 VDD1.n56 B 0.025767f
C248 VDD1.n57 B 0.011542f
C249 VDD1.n58 B 0.010901f
C250 VDD1.n59 B 0.020287f
C251 VDD1.n60 B 0.020287f
C252 VDD1.n61 B 0.010901f
C253 VDD1.n62 B 0.011542f
C254 VDD1.n63 B 0.025767f
C255 VDD1.n64 B 0.025767f
C256 VDD1.n65 B 0.011542f
C257 VDD1.n66 B 0.010901f
C258 VDD1.n67 B 0.020287f
C259 VDD1.n68 B 0.020287f
C260 VDD1.n69 B 0.010901f
C261 VDD1.n70 B 0.011542f
C262 VDD1.n71 B 0.025767f
C263 VDD1.n72 B 0.025767f
C264 VDD1.n73 B 0.011542f
C265 VDD1.n74 B 0.010901f
C266 VDD1.n75 B 0.020287f
C267 VDD1.n76 B 0.020287f
C268 VDD1.n77 B 0.010901f
C269 VDD1.n78 B 0.011542f
C270 VDD1.n79 B 0.025767f
C271 VDD1.n80 B 0.057475f
C272 VDD1.n81 B 0.011542f
C273 VDD1.n82 B 0.010901f
C274 VDD1.n83 B 0.053266f
C275 VDD1.n84 B 0.048059f
C276 VDD1.n85 B 0.029473f
C277 VDD1.n86 B 0.020287f
C278 VDD1.n87 B 0.010901f
C279 VDD1.n88 B 0.025767f
C280 VDD1.n89 B 0.011222f
C281 VDD1.n90 B 0.020287f
C282 VDD1.n91 B 0.011542f
C283 VDD1.n92 B 0.025767f
C284 VDD1.n93 B 0.011542f
C285 VDD1.n94 B 0.020287f
C286 VDD1.n95 B 0.010901f
C287 VDD1.n96 B 0.025767f
C288 VDD1.n97 B 0.011542f
C289 VDD1.n98 B 0.020287f
C290 VDD1.n99 B 0.010901f
C291 VDD1.n100 B 0.025767f
C292 VDD1.n101 B 0.011542f
C293 VDD1.n102 B 0.020287f
C294 VDD1.n103 B 0.010901f
C295 VDD1.n104 B 0.025767f
C296 VDD1.n105 B 0.011542f
C297 VDD1.n106 B 0.020287f
C298 VDD1.n107 B 0.010901f
C299 VDD1.n108 B 0.025767f
C300 VDD1.n109 B 0.011542f
C301 VDD1.n110 B 1.37474f
C302 VDD1.n111 B 0.010901f
C303 VDD1.t1 B 0.042527f
C304 VDD1.n112 B 0.135315f
C305 VDD1.n113 B 0.015221f
C306 VDD1.n114 B 0.019325f
C307 VDD1.n115 B 0.025767f
C308 VDD1.n116 B 0.011542f
C309 VDD1.n117 B 0.010901f
C310 VDD1.n118 B 0.020287f
C311 VDD1.n119 B 0.020287f
C312 VDD1.n120 B 0.010901f
C313 VDD1.n121 B 0.011542f
C314 VDD1.n122 B 0.025767f
C315 VDD1.n123 B 0.025767f
C316 VDD1.n124 B 0.011542f
C317 VDD1.n125 B 0.010901f
C318 VDD1.n126 B 0.020287f
C319 VDD1.n127 B 0.020287f
C320 VDD1.n128 B 0.010901f
C321 VDD1.n129 B 0.011542f
C322 VDD1.n130 B 0.025767f
C323 VDD1.n131 B 0.025767f
C324 VDD1.n132 B 0.011542f
C325 VDD1.n133 B 0.010901f
C326 VDD1.n134 B 0.020287f
C327 VDD1.n135 B 0.020287f
C328 VDD1.n136 B 0.010901f
C329 VDD1.n137 B 0.011542f
C330 VDD1.n138 B 0.025767f
C331 VDD1.n139 B 0.025767f
C332 VDD1.n140 B 0.011542f
C333 VDD1.n141 B 0.010901f
C334 VDD1.n142 B 0.020287f
C335 VDD1.n143 B 0.020287f
C336 VDD1.n144 B 0.010901f
C337 VDD1.n145 B 0.011542f
C338 VDD1.n146 B 0.025767f
C339 VDD1.n147 B 0.025767f
C340 VDD1.n148 B 0.011542f
C341 VDD1.n149 B 0.010901f
C342 VDD1.n150 B 0.020287f
C343 VDD1.n151 B 0.020287f
C344 VDD1.n152 B 0.010901f
C345 VDD1.n153 B 0.010901f
C346 VDD1.n154 B 0.011542f
C347 VDD1.n155 B 0.025767f
C348 VDD1.n156 B 0.025767f
C349 VDD1.n157 B 0.025767f
C350 VDD1.n158 B 0.011222f
C351 VDD1.n159 B 0.010901f
C352 VDD1.n160 B 0.020287f
C353 VDD1.n161 B 0.020287f
C354 VDD1.n162 B 0.010901f
C355 VDD1.n163 B 0.011542f
C356 VDD1.n164 B 0.025767f
C357 VDD1.n165 B 0.057475f
C358 VDD1.n166 B 0.011542f
C359 VDD1.n167 B 0.010901f
C360 VDD1.n168 B 0.053266f
C361 VDD1.n169 B 0.765461f
C362 VTAIL.n0 B 0.029385f
C363 VTAIL.n1 B 0.020226f
C364 VTAIL.n2 B 0.010869f
C365 VTAIL.n3 B 0.02569f
C366 VTAIL.n4 B 0.011189f
C367 VTAIL.n5 B 0.020226f
C368 VTAIL.n6 B 0.011508f
C369 VTAIL.n7 B 0.02569f
C370 VTAIL.n8 B 0.011508f
C371 VTAIL.n9 B 0.020226f
C372 VTAIL.n10 B 0.010869f
C373 VTAIL.n11 B 0.02569f
C374 VTAIL.n12 B 0.011508f
C375 VTAIL.n13 B 0.020226f
C376 VTAIL.n14 B 0.010869f
C377 VTAIL.n15 B 0.02569f
C378 VTAIL.n16 B 0.011508f
C379 VTAIL.n17 B 0.020226f
C380 VTAIL.n18 B 0.010869f
C381 VTAIL.n19 B 0.02569f
C382 VTAIL.n20 B 0.011508f
C383 VTAIL.n21 B 0.020226f
C384 VTAIL.n22 B 0.010869f
C385 VTAIL.n23 B 0.02569f
C386 VTAIL.n24 B 0.011508f
C387 VTAIL.n25 B 1.37065f
C388 VTAIL.n26 B 0.010869f
C389 VTAIL.t3 B 0.0424f
C390 VTAIL.n27 B 0.134913f
C391 VTAIL.n28 B 0.015176f
C392 VTAIL.n29 B 0.019267f
C393 VTAIL.n30 B 0.02569f
C394 VTAIL.n31 B 0.011508f
C395 VTAIL.n32 B 0.010869f
C396 VTAIL.n33 B 0.020226f
C397 VTAIL.n34 B 0.020226f
C398 VTAIL.n35 B 0.010869f
C399 VTAIL.n36 B 0.011508f
C400 VTAIL.n37 B 0.02569f
C401 VTAIL.n38 B 0.02569f
C402 VTAIL.n39 B 0.011508f
C403 VTAIL.n40 B 0.010869f
C404 VTAIL.n41 B 0.020226f
C405 VTAIL.n42 B 0.020226f
C406 VTAIL.n43 B 0.010869f
C407 VTAIL.n44 B 0.011508f
C408 VTAIL.n45 B 0.02569f
C409 VTAIL.n46 B 0.02569f
C410 VTAIL.n47 B 0.011508f
C411 VTAIL.n48 B 0.010869f
C412 VTAIL.n49 B 0.020226f
C413 VTAIL.n50 B 0.020226f
C414 VTAIL.n51 B 0.010869f
C415 VTAIL.n52 B 0.011508f
C416 VTAIL.n53 B 0.02569f
C417 VTAIL.n54 B 0.02569f
C418 VTAIL.n55 B 0.011508f
C419 VTAIL.n56 B 0.010869f
C420 VTAIL.n57 B 0.020226f
C421 VTAIL.n58 B 0.020226f
C422 VTAIL.n59 B 0.010869f
C423 VTAIL.n60 B 0.011508f
C424 VTAIL.n61 B 0.02569f
C425 VTAIL.n62 B 0.02569f
C426 VTAIL.n63 B 0.011508f
C427 VTAIL.n64 B 0.010869f
C428 VTAIL.n65 B 0.020226f
C429 VTAIL.n66 B 0.020226f
C430 VTAIL.n67 B 0.010869f
C431 VTAIL.n68 B 0.010869f
C432 VTAIL.n69 B 0.011508f
C433 VTAIL.n70 B 0.02569f
C434 VTAIL.n71 B 0.02569f
C435 VTAIL.n72 B 0.02569f
C436 VTAIL.n73 B 0.011189f
C437 VTAIL.n74 B 0.010869f
C438 VTAIL.n75 B 0.020226f
C439 VTAIL.n76 B 0.020226f
C440 VTAIL.n77 B 0.010869f
C441 VTAIL.n78 B 0.011508f
C442 VTAIL.n79 B 0.02569f
C443 VTAIL.n80 B 0.057303f
C444 VTAIL.n81 B 0.011508f
C445 VTAIL.n82 B 0.010869f
C446 VTAIL.n83 B 0.053107f
C447 VTAIL.n84 B 0.032422f
C448 VTAIL.n85 B 1.67748f
C449 VTAIL.n86 B 0.029385f
C450 VTAIL.n87 B 0.020226f
C451 VTAIL.n88 B 0.010869f
C452 VTAIL.n89 B 0.02569f
C453 VTAIL.n90 B 0.011189f
C454 VTAIL.n91 B 0.020226f
C455 VTAIL.n92 B 0.011189f
C456 VTAIL.n93 B 0.010869f
C457 VTAIL.n94 B 0.02569f
C458 VTAIL.n95 B 0.02569f
C459 VTAIL.n96 B 0.011508f
C460 VTAIL.n97 B 0.020226f
C461 VTAIL.n98 B 0.010869f
C462 VTAIL.n99 B 0.02569f
C463 VTAIL.n100 B 0.011508f
C464 VTAIL.n101 B 0.020226f
C465 VTAIL.n102 B 0.010869f
C466 VTAIL.n103 B 0.02569f
C467 VTAIL.n104 B 0.011508f
C468 VTAIL.n105 B 0.020226f
C469 VTAIL.n106 B 0.010869f
C470 VTAIL.n107 B 0.02569f
C471 VTAIL.n108 B 0.011508f
C472 VTAIL.n109 B 0.020226f
C473 VTAIL.n110 B 0.010869f
C474 VTAIL.n111 B 0.02569f
C475 VTAIL.n112 B 0.011508f
C476 VTAIL.n113 B 1.37065f
C477 VTAIL.n114 B 0.010869f
C478 VTAIL.t1 B 0.0424f
C479 VTAIL.n115 B 0.134913f
C480 VTAIL.n116 B 0.015176f
C481 VTAIL.n117 B 0.019267f
C482 VTAIL.n118 B 0.02569f
C483 VTAIL.n119 B 0.011508f
C484 VTAIL.n120 B 0.010869f
C485 VTAIL.n121 B 0.020226f
C486 VTAIL.n122 B 0.020226f
C487 VTAIL.n123 B 0.010869f
C488 VTAIL.n124 B 0.011508f
C489 VTAIL.n125 B 0.02569f
C490 VTAIL.n126 B 0.02569f
C491 VTAIL.n127 B 0.011508f
C492 VTAIL.n128 B 0.010869f
C493 VTAIL.n129 B 0.020226f
C494 VTAIL.n130 B 0.020226f
C495 VTAIL.n131 B 0.010869f
C496 VTAIL.n132 B 0.011508f
C497 VTAIL.n133 B 0.02569f
C498 VTAIL.n134 B 0.02569f
C499 VTAIL.n135 B 0.011508f
C500 VTAIL.n136 B 0.010869f
C501 VTAIL.n137 B 0.020226f
C502 VTAIL.n138 B 0.020226f
C503 VTAIL.n139 B 0.010869f
C504 VTAIL.n140 B 0.011508f
C505 VTAIL.n141 B 0.02569f
C506 VTAIL.n142 B 0.02569f
C507 VTAIL.n143 B 0.011508f
C508 VTAIL.n144 B 0.010869f
C509 VTAIL.n145 B 0.020226f
C510 VTAIL.n146 B 0.020226f
C511 VTAIL.n147 B 0.010869f
C512 VTAIL.n148 B 0.011508f
C513 VTAIL.n149 B 0.02569f
C514 VTAIL.n150 B 0.02569f
C515 VTAIL.n151 B 0.011508f
C516 VTAIL.n152 B 0.010869f
C517 VTAIL.n153 B 0.020226f
C518 VTAIL.n154 B 0.020226f
C519 VTAIL.n155 B 0.010869f
C520 VTAIL.n156 B 0.011508f
C521 VTAIL.n157 B 0.02569f
C522 VTAIL.n158 B 0.02569f
C523 VTAIL.n159 B 0.011508f
C524 VTAIL.n160 B 0.010869f
C525 VTAIL.n161 B 0.020226f
C526 VTAIL.n162 B 0.020226f
C527 VTAIL.n163 B 0.010869f
C528 VTAIL.n164 B 0.011508f
C529 VTAIL.n165 B 0.02569f
C530 VTAIL.n166 B 0.057303f
C531 VTAIL.n167 B 0.011508f
C532 VTAIL.n168 B 0.010869f
C533 VTAIL.n169 B 0.053107f
C534 VTAIL.n170 B 0.032422f
C535 VTAIL.n171 B 1.72608f
C536 VTAIL.n172 B 0.029385f
C537 VTAIL.n173 B 0.020226f
C538 VTAIL.n174 B 0.010869f
C539 VTAIL.n175 B 0.02569f
C540 VTAIL.n176 B 0.011189f
C541 VTAIL.n177 B 0.020226f
C542 VTAIL.n178 B 0.011189f
C543 VTAIL.n179 B 0.010869f
C544 VTAIL.n180 B 0.02569f
C545 VTAIL.n181 B 0.02569f
C546 VTAIL.n182 B 0.011508f
C547 VTAIL.n183 B 0.020226f
C548 VTAIL.n184 B 0.010869f
C549 VTAIL.n185 B 0.02569f
C550 VTAIL.n186 B 0.011508f
C551 VTAIL.n187 B 0.020226f
C552 VTAIL.n188 B 0.010869f
C553 VTAIL.n189 B 0.02569f
C554 VTAIL.n190 B 0.011508f
C555 VTAIL.n191 B 0.020226f
C556 VTAIL.n192 B 0.010869f
C557 VTAIL.n193 B 0.02569f
C558 VTAIL.n194 B 0.011508f
C559 VTAIL.n195 B 0.020226f
C560 VTAIL.n196 B 0.010869f
C561 VTAIL.n197 B 0.02569f
C562 VTAIL.n198 B 0.011508f
C563 VTAIL.n199 B 1.37065f
C564 VTAIL.n200 B 0.010869f
C565 VTAIL.t2 B 0.0424f
C566 VTAIL.n201 B 0.134913f
C567 VTAIL.n202 B 0.015176f
C568 VTAIL.n203 B 0.019267f
C569 VTAIL.n204 B 0.02569f
C570 VTAIL.n205 B 0.011508f
C571 VTAIL.n206 B 0.010869f
C572 VTAIL.n207 B 0.020226f
C573 VTAIL.n208 B 0.020226f
C574 VTAIL.n209 B 0.010869f
C575 VTAIL.n210 B 0.011508f
C576 VTAIL.n211 B 0.02569f
C577 VTAIL.n212 B 0.02569f
C578 VTAIL.n213 B 0.011508f
C579 VTAIL.n214 B 0.010869f
C580 VTAIL.n215 B 0.020226f
C581 VTAIL.n216 B 0.020226f
C582 VTAIL.n217 B 0.010869f
C583 VTAIL.n218 B 0.011508f
C584 VTAIL.n219 B 0.02569f
C585 VTAIL.n220 B 0.02569f
C586 VTAIL.n221 B 0.011508f
C587 VTAIL.n222 B 0.010869f
C588 VTAIL.n223 B 0.020226f
C589 VTAIL.n224 B 0.020226f
C590 VTAIL.n225 B 0.010869f
C591 VTAIL.n226 B 0.011508f
C592 VTAIL.n227 B 0.02569f
C593 VTAIL.n228 B 0.02569f
C594 VTAIL.n229 B 0.011508f
C595 VTAIL.n230 B 0.010869f
C596 VTAIL.n231 B 0.020226f
C597 VTAIL.n232 B 0.020226f
C598 VTAIL.n233 B 0.010869f
C599 VTAIL.n234 B 0.011508f
C600 VTAIL.n235 B 0.02569f
C601 VTAIL.n236 B 0.02569f
C602 VTAIL.n237 B 0.011508f
C603 VTAIL.n238 B 0.010869f
C604 VTAIL.n239 B 0.020226f
C605 VTAIL.n240 B 0.020226f
C606 VTAIL.n241 B 0.010869f
C607 VTAIL.n242 B 0.011508f
C608 VTAIL.n243 B 0.02569f
C609 VTAIL.n244 B 0.02569f
C610 VTAIL.n245 B 0.011508f
C611 VTAIL.n246 B 0.010869f
C612 VTAIL.n247 B 0.020226f
C613 VTAIL.n248 B 0.020226f
C614 VTAIL.n249 B 0.010869f
C615 VTAIL.n250 B 0.011508f
C616 VTAIL.n251 B 0.02569f
C617 VTAIL.n252 B 0.057303f
C618 VTAIL.n253 B 0.011508f
C619 VTAIL.n254 B 0.010869f
C620 VTAIL.n255 B 0.053107f
C621 VTAIL.n256 B 0.032422f
C622 VTAIL.n257 B 1.51651f
C623 VTAIL.n258 B 0.029385f
C624 VTAIL.n259 B 0.020226f
C625 VTAIL.n260 B 0.010869f
C626 VTAIL.n261 B 0.02569f
C627 VTAIL.n262 B 0.011189f
C628 VTAIL.n263 B 0.020226f
C629 VTAIL.n264 B 0.011508f
C630 VTAIL.n265 B 0.02569f
C631 VTAIL.n266 B 0.011508f
C632 VTAIL.n267 B 0.020226f
C633 VTAIL.n268 B 0.010869f
C634 VTAIL.n269 B 0.02569f
C635 VTAIL.n270 B 0.011508f
C636 VTAIL.n271 B 0.020226f
C637 VTAIL.n272 B 0.010869f
C638 VTAIL.n273 B 0.02569f
C639 VTAIL.n274 B 0.011508f
C640 VTAIL.n275 B 0.020226f
C641 VTAIL.n276 B 0.010869f
C642 VTAIL.n277 B 0.02569f
C643 VTAIL.n278 B 0.011508f
C644 VTAIL.n279 B 0.020226f
C645 VTAIL.n280 B 0.010869f
C646 VTAIL.n281 B 0.02569f
C647 VTAIL.n282 B 0.011508f
C648 VTAIL.n283 B 1.37065f
C649 VTAIL.n284 B 0.010869f
C650 VTAIL.t0 B 0.0424f
C651 VTAIL.n285 B 0.134913f
C652 VTAIL.n286 B 0.015176f
C653 VTAIL.n287 B 0.019267f
C654 VTAIL.n288 B 0.02569f
C655 VTAIL.n289 B 0.011508f
C656 VTAIL.n290 B 0.010869f
C657 VTAIL.n291 B 0.020226f
C658 VTAIL.n292 B 0.020226f
C659 VTAIL.n293 B 0.010869f
C660 VTAIL.n294 B 0.011508f
C661 VTAIL.n295 B 0.02569f
C662 VTAIL.n296 B 0.02569f
C663 VTAIL.n297 B 0.011508f
C664 VTAIL.n298 B 0.010869f
C665 VTAIL.n299 B 0.020226f
C666 VTAIL.n300 B 0.020226f
C667 VTAIL.n301 B 0.010869f
C668 VTAIL.n302 B 0.011508f
C669 VTAIL.n303 B 0.02569f
C670 VTAIL.n304 B 0.02569f
C671 VTAIL.n305 B 0.011508f
C672 VTAIL.n306 B 0.010869f
C673 VTAIL.n307 B 0.020226f
C674 VTAIL.n308 B 0.020226f
C675 VTAIL.n309 B 0.010869f
C676 VTAIL.n310 B 0.011508f
C677 VTAIL.n311 B 0.02569f
C678 VTAIL.n312 B 0.02569f
C679 VTAIL.n313 B 0.011508f
C680 VTAIL.n314 B 0.010869f
C681 VTAIL.n315 B 0.020226f
C682 VTAIL.n316 B 0.020226f
C683 VTAIL.n317 B 0.010869f
C684 VTAIL.n318 B 0.011508f
C685 VTAIL.n319 B 0.02569f
C686 VTAIL.n320 B 0.02569f
C687 VTAIL.n321 B 0.011508f
C688 VTAIL.n322 B 0.010869f
C689 VTAIL.n323 B 0.020226f
C690 VTAIL.n324 B 0.020226f
C691 VTAIL.n325 B 0.010869f
C692 VTAIL.n326 B 0.010869f
C693 VTAIL.n327 B 0.011508f
C694 VTAIL.n328 B 0.02569f
C695 VTAIL.n329 B 0.02569f
C696 VTAIL.n330 B 0.02569f
C697 VTAIL.n331 B 0.011189f
C698 VTAIL.n332 B 0.010869f
C699 VTAIL.n333 B 0.020226f
C700 VTAIL.n334 B 0.020226f
C701 VTAIL.n335 B 0.010869f
C702 VTAIL.n336 B 0.011508f
C703 VTAIL.n337 B 0.02569f
C704 VTAIL.n338 B 0.057303f
C705 VTAIL.n339 B 0.011508f
C706 VTAIL.n340 B 0.010869f
C707 VTAIL.n341 B 0.053107f
C708 VTAIL.n342 B 0.032422f
C709 VTAIL.n343 B 1.42971f
C710 VP.t1 B 4.78198f
C711 VP.t0 B 4.11599f
C712 VP.n0 B 4.60925f
.ends

