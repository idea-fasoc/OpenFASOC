* NGSPICE file created from diff_pair_sample_1711.ext - technology: sky130A

.subckt diff_pair_sample_1711 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=3.46
X1 VDD1.t4 VP.t1 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=3.46
X2 VDD2.t5 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=3.46
X3 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=3.46
X4 VTAIL.t11 VN.t2 VDD2.t3 B.t19 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=0.82335 ps=5.32 w=4.99 l=3.46
X5 VTAIL.t8 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=0.82335 ps=5.32 w=4.99 l=3.46
X6 VDD1.t2 VP.t3 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=3.46
X7 B.t18 B.t16 B.t17 B.t10 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=3.46
X8 B.t15 B.t13 B.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=3.46
X9 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=3.46
X10 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=3.46
X11 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=3.46
X12 VDD1.t1 VP.t4 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=3.46
X13 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=0.82335 ps=5.32 w=4.99 l=3.46
X14 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=3.46
X15 VTAIL.t5 VP.t5 VDD1.t0 B.t19 sky130_fd_pr__nfet_01v8 ad=0.82335 pd=5.32 as=0.82335 ps=5.32 w=4.99 l=3.46
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n50 VP.n49 161.3
R8 VP.n48 VP.n1 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n2 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n42 VP.n3 161.3
R13 VP.n41 VP.n40 161.3
R14 VP.n39 VP.n4 161.3
R15 VP.n38 VP.n37 161.3
R16 VP.n36 VP.n5 161.3
R17 VP.n35 VP.n34 161.3
R18 VP.n33 VP.n6 161.3
R19 VP.n32 VP.n31 161.3
R20 VP.n30 VP.n7 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n27 VP.n8 75.8765
R23 VP.n51 VP.n0 75.8765
R24 VP.n26 VP.n9 75.8765
R25 VP.n14 VP.t1 68.783
R26 VP.n35 VP.n6 50.6917
R27 VP.n43 VP.n2 50.6917
R28 VP.n18 VP.n11 50.6917
R29 VP.n14 VP.n13 50.1886
R30 VP.n27 VP.n26 46.8819
R31 VP.n4 VP.t2 34.7574
R32 VP.n8 VP.t4 34.7574
R33 VP.n0 VP.t3 34.7574
R34 VP.n13 VP.t5 34.7574
R35 VP.n9 VP.t0 34.7574
R36 VP.n31 VP.n6 30.2951
R37 VP.n47 VP.n2 30.2951
R38 VP.n22 VP.n11 30.2951
R39 VP.n30 VP.n29 24.4675
R40 VP.n31 VP.n30 24.4675
R41 VP.n36 VP.n35 24.4675
R42 VP.n37 VP.n36 24.4675
R43 VP.n37 VP.n4 24.4675
R44 VP.n41 VP.n4 24.4675
R45 VP.n42 VP.n41 24.4675
R46 VP.n43 VP.n42 24.4675
R47 VP.n48 VP.n47 24.4675
R48 VP.n49 VP.n48 24.4675
R49 VP.n23 VP.n22 24.4675
R50 VP.n24 VP.n23 24.4675
R51 VP.n16 VP.n13 24.4675
R52 VP.n17 VP.n16 24.4675
R53 VP.n18 VP.n17 24.4675
R54 VP.n29 VP.n8 14.1914
R55 VP.n49 VP.n0 14.1914
R56 VP.n24 VP.n9 14.1914
R57 VP.n15 VP.n14 3.01035
R58 VP.n26 VP.n25 0.354971
R59 VP.n28 VP.n27 0.354971
R60 VP.n51 VP.n50 0.354971
R61 VP VP.n51 0.26696
R62 VP.n15 VP.n12 0.189894
R63 VP.n19 VP.n12 0.189894
R64 VP.n20 VP.n19 0.189894
R65 VP.n21 VP.n20 0.189894
R66 VP.n21 VP.n10 0.189894
R67 VP.n25 VP.n10 0.189894
R68 VP.n28 VP.n7 0.189894
R69 VP.n32 VP.n7 0.189894
R70 VP.n33 VP.n32 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n34 VP.n5 0.189894
R73 VP.n38 VP.n5 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n40 VP.n3 0.189894
R77 VP.n44 VP.n3 0.189894
R78 VP.n45 VP.n44 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n46 VP.n1 0.189894
R81 VP.n50 VP.n1 0.189894
R82 VTAIL.n7 VTAIL.t4 58.2137
R83 VTAIL.n11 VTAIL.t3 58.2137
R84 VTAIL.n2 VTAIL.t9 58.2137
R85 VTAIL.n10 VTAIL.t6 58.2137
R86 VTAIL.n9 VTAIL.n8 54.2459
R87 VTAIL.n6 VTAIL.n5 54.2459
R88 VTAIL.n1 VTAIL.n0 54.2456
R89 VTAIL.n4 VTAIL.n3 54.2456
R90 VTAIL.n6 VTAIL.n4 23.2031
R91 VTAIL.n11 VTAIL.n10 19.9358
R92 VTAIL.n0 VTAIL.t1 3.96844
R93 VTAIL.n0 VTAIL.t11 3.96844
R94 VTAIL.n3 VTAIL.t10 3.96844
R95 VTAIL.n3 VTAIL.t8 3.96844
R96 VTAIL.n8 VTAIL.t7 3.96844
R97 VTAIL.n8 VTAIL.t5 3.96844
R98 VTAIL.n5 VTAIL.t2 3.96844
R99 VTAIL.n5 VTAIL.t0 3.96844
R100 VTAIL.n7 VTAIL.n6 3.26774
R101 VTAIL.n10 VTAIL.n9 3.26774
R102 VTAIL.n4 VTAIL.n2 3.26774
R103 VTAIL VTAIL.n11 2.39274
R104 VTAIL.n9 VTAIL.n7 2.10395
R105 VTAIL.n2 VTAIL.n1 2.10395
R106 VTAIL VTAIL.n1 0.8755
R107 VDD1 VDD1.t4 77.4011
R108 VDD1.n1 VDD1.t1 77.2875
R109 VDD1.n1 VDD1.n0 71.6859
R110 VDD1.n3 VDD1.n2 70.9245
R111 VDD1.n3 VDD1.n1 40.8522
R112 VDD1.n2 VDD1.t0 3.96844
R113 VDD1.n2 VDD1.t5 3.96844
R114 VDD1.n0 VDD1.t3 3.96844
R115 VDD1.n0 VDD1.t2 3.96844
R116 VDD1 VDD1.n3 0.759121
R117 B.n691 B.n690 585
R118 B.n228 B.n123 585
R119 B.n227 B.n226 585
R120 B.n225 B.n224 585
R121 B.n223 B.n222 585
R122 B.n221 B.n220 585
R123 B.n219 B.n218 585
R124 B.n217 B.n216 585
R125 B.n215 B.n214 585
R126 B.n213 B.n212 585
R127 B.n211 B.n210 585
R128 B.n209 B.n208 585
R129 B.n207 B.n206 585
R130 B.n205 B.n204 585
R131 B.n203 B.n202 585
R132 B.n201 B.n200 585
R133 B.n199 B.n198 585
R134 B.n197 B.n196 585
R135 B.n195 B.n194 585
R136 B.n193 B.n192 585
R137 B.n191 B.n190 585
R138 B.n188 B.n187 585
R139 B.n186 B.n185 585
R140 B.n184 B.n183 585
R141 B.n182 B.n181 585
R142 B.n180 B.n179 585
R143 B.n178 B.n177 585
R144 B.n176 B.n175 585
R145 B.n174 B.n173 585
R146 B.n172 B.n171 585
R147 B.n170 B.n169 585
R148 B.n167 B.n166 585
R149 B.n165 B.n164 585
R150 B.n163 B.n162 585
R151 B.n161 B.n160 585
R152 B.n159 B.n158 585
R153 B.n157 B.n156 585
R154 B.n155 B.n154 585
R155 B.n153 B.n152 585
R156 B.n151 B.n150 585
R157 B.n149 B.n148 585
R158 B.n147 B.n146 585
R159 B.n145 B.n144 585
R160 B.n143 B.n142 585
R161 B.n141 B.n140 585
R162 B.n139 B.n138 585
R163 B.n137 B.n136 585
R164 B.n135 B.n134 585
R165 B.n133 B.n132 585
R166 B.n131 B.n130 585
R167 B.n129 B.n128 585
R168 B.n96 B.n95 585
R169 B.n689 B.n97 585
R170 B.n694 B.n97 585
R171 B.n688 B.n687 585
R172 B.n687 B.n93 585
R173 B.n686 B.n92 585
R174 B.n700 B.n92 585
R175 B.n685 B.n91 585
R176 B.n701 B.n91 585
R177 B.n684 B.n90 585
R178 B.n702 B.n90 585
R179 B.n683 B.n682 585
R180 B.n682 B.n86 585
R181 B.n681 B.n85 585
R182 B.n708 B.n85 585
R183 B.n680 B.n84 585
R184 B.n709 B.n84 585
R185 B.n679 B.n83 585
R186 B.n710 B.n83 585
R187 B.n678 B.n677 585
R188 B.n677 B.n79 585
R189 B.n676 B.n78 585
R190 B.n716 B.n78 585
R191 B.n675 B.n77 585
R192 B.n717 B.n77 585
R193 B.n674 B.n76 585
R194 B.n718 B.n76 585
R195 B.n673 B.n672 585
R196 B.n672 B.n72 585
R197 B.n671 B.n71 585
R198 B.n724 B.n71 585
R199 B.n670 B.n70 585
R200 B.n725 B.n70 585
R201 B.n669 B.n69 585
R202 B.n726 B.n69 585
R203 B.n668 B.n667 585
R204 B.n667 B.n65 585
R205 B.n666 B.n64 585
R206 B.n732 B.n64 585
R207 B.n665 B.n63 585
R208 B.n733 B.n63 585
R209 B.n664 B.n62 585
R210 B.n734 B.n62 585
R211 B.n663 B.n662 585
R212 B.n662 B.n58 585
R213 B.n661 B.n57 585
R214 B.n740 B.n57 585
R215 B.n660 B.n56 585
R216 B.n741 B.n56 585
R217 B.n659 B.n55 585
R218 B.n742 B.n55 585
R219 B.n658 B.n657 585
R220 B.n657 B.n51 585
R221 B.n656 B.n50 585
R222 B.n748 B.n50 585
R223 B.n655 B.n49 585
R224 B.n749 B.n49 585
R225 B.n654 B.n48 585
R226 B.n750 B.n48 585
R227 B.n653 B.n652 585
R228 B.n652 B.n44 585
R229 B.n651 B.n43 585
R230 B.n756 B.n43 585
R231 B.n650 B.n42 585
R232 B.n757 B.n42 585
R233 B.n649 B.n41 585
R234 B.n758 B.n41 585
R235 B.n648 B.n647 585
R236 B.n647 B.n37 585
R237 B.n646 B.n36 585
R238 B.n764 B.n36 585
R239 B.n645 B.n35 585
R240 B.n765 B.n35 585
R241 B.n644 B.n34 585
R242 B.n766 B.n34 585
R243 B.n643 B.n642 585
R244 B.n642 B.n30 585
R245 B.n641 B.n29 585
R246 B.n772 B.n29 585
R247 B.n640 B.n28 585
R248 B.n773 B.n28 585
R249 B.n639 B.n27 585
R250 B.n774 B.n27 585
R251 B.n638 B.n637 585
R252 B.n637 B.n23 585
R253 B.n636 B.n22 585
R254 B.n780 B.n22 585
R255 B.n635 B.n21 585
R256 B.n781 B.n21 585
R257 B.n634 B.n20 585
R258 B.n782 B.n20 585
R259 B.n633 B.n632 585
R260 B.n632 B.n19 585
R261 B.n631 B.n15 585
R262 B.n788 B.n15 585
R263 B.n630 B.n14 585
R264 B.n789 B.n14 585
R265 B.n629 B.n13 585
R266 B.n790 B.n13 585
R267 B.n628 B.n627 585
R268 B.n627 B.n12 585
R269 B.n626 B.n625 585
R270 B.n626 B.n8 585
R271 B.n624 B.n7 585
R272 B.n797 B.n7 585
R273 B.n623 B.n6 585
R274 B.n798 B.n6 585
R275 B.n622 B.n5 585
R276 B.n799 B.n5 585
R277 B.n621 B.n620 585
R278 B.n620 B.n4 585
R279 B.n619 B.n229 585
R280 B.n619 B.n618 585
R281 B.n609 B.n230 585
R282 B.n231 B.n230 585
R283 B.n611 B.n610 585
R284 B.n612 B.n611 585
R285 B.n608 B.n236 585
R286 B.n236 B.n235 585
R287 B.n607 B.n606 585
R288 B.n606 B.n605 585
R289 B.n238 B.n237 585
R290 B.n598 B.n238 585
R291 B.n597 B.n596 585
R292 B.n599 B.n597 585
R293 B.n595 B.n243 585
R294 B.n243 B.n242 585
R295 B.n594 B.n593 585
R296 B.n593 B.n592 585
R297 B.n245 B.n244 585
R298 B.n246 B.n245 585
R299 B.n585 B.n584 585
R300 B.n586 B.n585 585
R301 B.n583 B.n251 585
R302 B.n251 B.n250 585
R303 B.n582 B.n581 585
R304 B.n581 B.n580 585
R305 B.n253 B.n252 585
R306 B.n254 B.n253 585
R307 B.n573 B.n572 585
R308 B.n574 B.n573 585
R309 B.n571 B.n259 585
R310 B.n259 B.n258 585
R311 B.n570 B.n569 585
R312 B.n569 B.n568 585
R313 B.n261 B.n260 585
R314 B.n262 B.n261 585
R315 B.n561 B.n560 585
R316 B.n562 B.n561 585
R317 B.n559 B.n267 585
R318 B.n267 B.n266 585
R319 B.n558 B.n557 585
R320 B.n557 B.n556 585
R321 B.n269 B.n268 585
R322 B.n270 B.n269 585
R323 B.n549 B.n548 585
R324 B.n550 B.n549 585
R325 B.n547 B.n275 585
R326 B.n275 B.n274 585
R327 B.n546 B.n545 585
R328 B.n545 B.n544 585
R329 B.n277 B.n276 585
R330 B.n278 B.n277 585
R331 B.n537 B.n536 585
R332 B.n538 B.n537 585
R333 B.n535 B.n282 585
R334 B.n286 B.n282 585
R335 B.n534 B.n533 585
R336 B.n533 B.n532 585
R337 B.n284 B.n283 585
R338 B.n285 B.n284 585
R339 B.n525 B.n524 585
R340 B.n526 B.n525 585
R341 B.n523 B.n291 585
R342 B.n291 B.n290 585
R343 B.n522 B.n521 585
R344 B.n521 B.n520 585
R345 B.n293 B.n292 585
R346 B.n294 B.n293 585
R347 B.n513 B.n512 585
R348 B.n514 B.n513 585
R349 B.n511 B.n299 585
R350 B.n299 B.n298 585
R351 B.n510 B.n509 585
R352 B.n509 B.n508 585
R353 B.n301 B.n300 585
R354 B.n302 B.n301 585
R355 B.n501 B.n500 585
R356 B.n502 B.n501 585
R357 B.n499 B.n307 585
R358 B.n307 B.n306 585
R359 B.n498 B.n497 585
R360 B.n497 B.n496 585
R361 B.n309 B.n308 585
R362 B.n310 B.n309 585
R363 B.n489 B.n488 585
R364 B.n490 B.n489 585
R365 B.n487 B.n315 585
R366 B.n315 B.n314 585
R367 B.n486 B.n485 585
R368 B.n485 B.n484 585
R369 B.n317 B.n316 585
R370 B.n318 B.n317 585
R371 B.n477 B.n476 585
R372 B.n478 B.n477 585
R373 B.n475 B.n323 585
R374 B.n323 B.n322 585
R375 B.n474 B.n473 585
R376 B.n473 B.n472 585
R377 B.n325 B.n324 585
R378 B.n326 B.n325 585
R379 B.n465 B.n464 585
R380 B.n466 B.n465 585
R381 B.n329 B.n328 585
R382 B.n364 B.n363 585
R383 B.n365 B.n361 585
R384 B.n361 B.n330 585
R385 B.n367 B.n366 585
R386 B.n369 B.n360 585
R387 B.n372 B.n371 585
R388 B.n373 B.n359 585
R389 B.n375 B.n374 585
R390 B.n377 B.n358 585
R391 B.n380 B.n379 585
R392 B.n381 B.n357 585
R393 B.n383 B.n382 585
R394 B.n385 B.n356 585
R395 B.n388 B.n387 585
R396 B.n389 B.n355 585
R397 B.n391 B.n390 585
R398 B.n393 B.n354 585
R399 B.n396 B.n395 585
R400 B.n397 B.n353 585
R401 B.n399 B.n398 585
R402 B.n401 B.n352 585
R403 B.n404 B.n403 585
R404 B.n405 B.n348 585
R405 B.n407 B.n406 585
R406 B.n409 B.n347 585
R407 B.n412 B.n411 585
R408 B.n413 B.n346 585
R409 B.n415 B.n414 585
R410 B.n417 B.n345 585
R411 B.n420 B.n419 585
R412 B.n421 B.n342 585
R413 B.n424 B.n423 585
R414 B.n426 B.n341 585
R415 B.n429 B.n428 585
R416 B.n430 B.n340 585
R417 B.n432 B.n431 585
R418 B.n434 B.n339 585
R419 B.n437 B.n436 585
R420 B.n438 B.n338 585
R421 B.n440 B.n439 585
R422 B.n442 B.n337 585
R423 B.n445 B.n444 585
R424 B.n446 B.n336 585
R425 B.n448 B.n447 585
R426 B.n450 B.n335 585
R427 B.n453 B.n452 585
R428 B.n454 B.n334 585
R429 B.n456 B.n455 585
R430 B.n458 B.n333 585
R431 B.n459 B.n332 585
R432 B.n462 B.n461 585
R433 B.n463 B.n331 585
R434 B.n331 B.n330 585
R435 B.n468 B.n467 585
R436 B.n467 B.n466 585
R437 B.n469 B.n327 585
R438 B.n327 B.n326 585
R439 B.n471 B.n470 585
R440 B.n472 B.n471 585
R441 B.n321 B.n320 585
R442 B.n322 B.n321 585
R443 B.n480 B.n479 585
R444 B.n479 B.n478 585
R445 B.n481 B.n319 585
R446 B.n319 B.n318 585
R447 B.n483 B.n482 585
R448 B.n484 B.n483 585
R449 B.n313 B.n312 585
R450 B.n314 B.n313 585
R451 B.n492 B.n491 585
R452 B.n491 B.n490 585
R453 B.n493 B.n311 585
R454 B.n311 B.n310 585
R455 B.n495 B.n494 585
R456 B.n496 B.n495 585
R457 B.n305 B.n304 585
R458 B.n306 B.n305 585
R459 B.n504 B.n503 585
R460 B.n503 B.n502 585
R461 B.n505 B.n303 585
R462 B.n303 B.n302 585
R463 B.n507 B.n506 585
R464 B.n508 B.n507 585
R465 B.n297 B.n296 585
R466 B.n298 B.n297 585
R467 B.n516 B.n515 585
R468 B.n515 B.n514 585
R469 B.n517 B.n295 585
R470 B.n295 B.n294 585
R471 B.n519 B.n518 585
R472 B.n520 B.n519 585
R473 B.n289 B.n288 585
R474 B.n290 B.n289 585
R475 B.n528 B.n527 585
R476 B.n527 B.n526 585
R477 B.n529 B.n287 585
R478 B.n287 B.n285 585
R479 B.n531 B.n530 585
R480 B.n532 B.n531 585
R481 B.n281 B.n280 585
R482 B.n286 B.n281 585
R483 B.n540 B.n539 585
R484 B.n539 B.n538 585
R485 B.n541 B.n279 585
R486 B.n279 B.n278 585
R487 B.n543 B.n542 585
R488 B.n544 B.n543 585
R489 B.n273 B.n272 585
R490 B.n274 B.n273 585
R491 B.n552 B.n551 585
R492 B.n551 B.n550 585
R493 B.n553 B.n271 585
R494 B.n271 B.n270 585
R495 B.n555 B.n554 585
R496 B.n556 B.n555 585
R497 B.n265 B.n264 585
R498 B.n266 B.n265 585
R499 B.n564 B.n563 585
R500 B.n563 B.n562 585
R501 B.n565 B.n263 585
R502 B.n263 B.n262 585
R503 B.n567 B.n566 585
R504 B.n568 B.n567 585
R505 B.n257 B.n256 585
R506 B.n258 B.n257 585
R507 B.n576 B.n575 585
R508 B.n575 B.n574 585
R509 B.n577 B.n255 585
R510 B.n255 B.n254 585
R511 B.n579 B.n578 585
R512 B.n580 B.n579 585
R513 B.n249 B.n248 585
R514 B.n250 B.n249 585
R515 B.n588 B.n587 585
R516 B.n587 B.n586 585
R517 B.n589 B.n247 585
R518 B.n247 B.n246 585
R519 B.n591 B.n590 585
R520 B.n592 B.n591 585
R521 B.n241 B.n240 585
R522 B.n242 B.n241 585
R523 B.n601 B.n600 585
R524 B.n600 B.n599 585
R525 B.n602 B.n239 585
R526 B.n598 B.n239 585
R527 B.n604 B.n603 585
R528 B.n605 B.n604 585
R529 B.n234 B.n233 585
R530 B.n235 B.n234 585
R531 B.n614 B.n613 585
R532 B.n613 B.n612 585
R533 B.n615 B.n232 585
R534 B.n232 B.n231 585
R535 B.n617 B.n616 585
R536 B.n618 B.n617 585
R537 B.n3 B.n0 585
R538 B.n4 B.n3 585
R539 B.n796 B.n1 585
R540 B.n797 B.n796 585
R541 B.n795 B.n794 585
R542 B.n795 B.n8 585
R543 B.n793 B.n9 585
R544 B.n12 B.n9 585
R545 B.n792 B.n791 585
R546 B.n791 B.n790 585
R547 B.n11 B.n10 585
R548 B.n789 B.n11 585
R549 B.n787 B.n786 585
R550 B.n788 B.n787 585
R551 B.n785 B.n16 585
R552 B.n19 B.n16 585
R553 B.n784 B.n783 585
R554 B.n783 B.n782 585
R555 B.n18 B.n17 585
R556 B.n781 B.n18 585
R557 B.n779 B.n778 585
R558 B.n780 B.n779 585
R559 B.n777 B.n24 585
R560 B.n24 B.n23 585
R561 B.n776 B.n775 585
R562 B.n775 B.n774 585
R563 B.n26 B.n25 585
R564 B.n773 B.n26 585
R565 B.n771 B.n770 585
R566 B.n772 B.n771 585
R567 B.n769 B.n31 585
R568 B.n31 B.n30 585
R569 B.n768 B.n767 585
R570 B.n767 B.n766 585
R571 B.n33 B.n32 585
R572 B.n765 B.n33 585
R573 B.n763 B.n762 585
R574 B.n764 B.n763 585
R575 B.n761 B.n38 585
R576 B.n38 B.n37 585
R577 B.n760 B.n759 585
R578 B.n759 B.n758 585
R579 B.n40 B.n39 585
R580 B.n757 B.n40 585
R581 B.n755 B.n754 585
R582 B.n756 B.n755 585
R583 B.n753 B.n45 585
R584 B.n45 B.n44 585
R585 B.n752 B.n751 585
R586 B.n751 B.n750 585
R587 B.n47 B.n46 585
R588 B.n749 B.n47 585
R589 B.n747 B.n746 585
R590 B.n748 B.n747 585
R591 B.n745 B.n52 585
R592 B.n52 B.n51 585
R593 B.n744 B.n743 585
R594 B.n743 B.n742 585
R595 B.n54 B.n53 585
R596 B.n741 B.n54 585
R597 B.n739 B.n738 585
R598 B.n740 B.n739 585
R599 B.n737 B.n59 585
R600 B.n59 B.n58 585
R601 B.n736 B.n735 585
R602 B.n735 B.n734 585
R603 B.n61 B.n60 585
R604 B.n733 B.n61 585
R605 B.n731 B.n730 585
R606 B.n732 B.n731 585
R607 B.n729 B.n66 585
R608 B.n66 B.n65 585
R609 B.n728 B.n727 585
R610 B.n727 B.n726 585
R611 B.n68 B.n67 585
R612 B.n725 B.n68 585
R613 B.n723 B.n722 585
R614 B.n724 B.n723 585
R615 B.n721 B.n73 585
R616 B.n73 B.n72 585
R617 B.n720 B.n719 585
R618 B.n719 B.n718 585
R619 B.n75 B.n74 585
R620 B.n717 B.n75 585
R621 B.n715 B.n714 585
R622 B.n716 B.n715 585
R623 B.n713 B.n80 585
R624 B.n80 B.n79 585
R625 B.n712 B.n711 585
R626 B.n711 B.n710 585
R627 B.n82 B.n81 585
R628 B.n709 B.n82 585
R629 B.n707 B.n706 585
R630 B.n708 B.n707 585
R631 B.n705 B.n87 585
R632 B.n87 B.n86 585
R633 B.n704 B.n703 585
R634 B.n703 B.n702 585
R635 B.n89 B.n88 585
R636 B.n701 B.n89 585
R637 B.n699 B.n698 585
R638 B.n700 B.n699 585
R639 B.n697 B.n94 585
R640 B.n94 B.n93 585
R641 B.n696 B.n695 585
R642 B.n695 B.n694 585
R643 B.n800 B.n799 585
R644 B.n798 B.n2 585
R645 B.n695 B.n96 497.305
R646 B.n691 B.n97 497.305
R647 B.n465 B.n331 497.305
R648 B.n467 B.n329 497.305
R649 B.n693 B.n692 256.663
R650 B.n693 B.n122 256.663
R651 B.n693 B.n121 256.663
R652 B.n693 B.n120 256.663
R653 B.n693 B.n119 256.663
R654 B.n693 B.n118 256.663
R655 B.n693 B.n117 256.663
R656 B.n693 B.n116 256.663
R657 B.n693 B.n115 256.663
R658 B.n693 B.n114 256.663
R659 B.n693 B.n113 256.663
R660 B.n693 B.n112 256.663
R661 B.n693 B.n111 256.663
R662 B.n693 B.n110 256.663
R663 B.n693 B.n109 256.663
R664 B.n693 B.n108 256.663
R665 B.n693 B.n107 256.663
R666 B.n693 B.n106 256.663
R667 B.n693 B.n105 256.663
R668 B.n693 B.n104 256.663
R669 B.n693 B.n103 256.663
R670 B.n693 B.n102 256.663
R671 B.n693 B.n101 256.663
R672 B.n693 B.n100 256.663
R673 B.n693 B.n99 256.663
R674 B.n693 B.n98 256.663
R675 B.n362 B.n330 256.663
R676 B.n368 B.n330 256.663
R677 B.n370 B.n330 256.663
R678 B.n376 B.n330 256.663
R679 B.n378 B.n330 256.663
R680 B.n384 B.n330 256.663
R681 B.n386 B.n330 256.663
R682 B.n392 B.n330 256.663
R683 B.n394 B.n330 256.663
R684 B.n400 B.n330 256.663
R685 B.n402 B.n330 256.663
R686 B.n408 B.n330 256.663
R687 B.n410 B.n330 256.663
R688 B.n416 B.n330 256.663
R689 B.n418 B.n330 256.663
R690 B.n425 B.n330 256.663
R691 B.n427 B.n330 256.663
R692 B.n433 B.n330 256.663
R693 B.n435 B.n330 256.663
R694 B.n441 B.n330 256.663
R695 B.n443 B.n330 256.663
R696 B.n449 B.n330 256.663
R697 B.n451 B.n330 256.663
R698 B.n457 B.n330 256.663
R699 B.n460 B.n330 256.663
R700 B.n802 B.n801 256.663
R701 B.n126 B.t13 243.815
R702 B.n124 B.t5 243.815
R703 B.n343 B.t16 243.815
R704 B.n349 B.t9 243.815
R705 B.n130 B.n129 163.367
R706 B.n134 B.n133 163.367
R707 B.n138 B.n137 163.367
R708 B.n142 B.n141 163.367
R709 B.n146 B.n145 163.367
R710 B.n150 B.n149 163.367
R711 B.n154 B.n153 163.367
R712 B.n158 B.n157 163.367
R713 B.n162 B.n161 163.367
R714 B.n166 B.n165 163.367
R715 B.n171 B.n170 163.367
R716 B.n175 B.n174 163.367
R717 B.n179 B.n178 163.367
R718 B.n183 B.n182 163.367
R719 B.n187 B.n186 163.367
R720 B.n192 B.n191 163.367
R721 B.n196 B.n195 163.367
R722 B.n200 B.n199 163.367
R723 B.n204 B.n203 163.367
R724 B.n208 B.n207 163.367
R725 B.n212 B.n211 163.367
R726 B.n216 B.n215 163.367
R727 B.n220 B.n219 163.367
R728 B.n224 B.n223 163.367
R729 B.n226 B.n123 163.367
R730 B.n465 B.n325 163.367
R731 B.n473 B.n325 163.367
R732 B.n473 B.n323 163.367
R733 B.n477 B.n323 163.367
R734 B.n477 B.n317 163.367
R735 B.n485 B.n317 163.367
R736 B.n485 B.n315 163.367
R737 B.n489 B.n315 163.367
R738 B.n489 B.n309 163.367
R739 B.n497 B.n309 163.367
R740 B.n497 B.n307 163.367
R741 B.n501 B.n307 163.367
R742 B.n501 B.n301 163.367
R743 B.n509 B.n301 163.367
R744 B.n509 B.n299 163.367
R745 B.n513 B.n299 163.367
R746 B.n513 B.n293 163.367
R747 B.n521 B.n293 163.367
R748 B.n521 B.n291 163.367
R749 B.n525 B.n291 163.367
R750 B.n525 B.n284 163.367
R751 B.n533 B.n284 163.367
R752 B.n533 B.n282 163.367
R753 B.n537 B.n282 163.367
R754 B.n537 B.n277 163.367
R755 B.n545 B.n277 163.367
R756 B.n545 B.n275 163.367
R757 B.n549 B.n275 163.367
R758 B.n549 B.n269 163.367
R759 B.n557 B.n269 163.367
R760 B.n557 B.n267 163.367
R761 B.n561 B.n267 163.367
R762 B.n561 B.n261 163.367
R763 B.n569 B.n261 163.367
R764 B.n569 B.n259 163.367
R765 B.n573 B.n259 163.367
R766 B.n573 B.n253 163.367
R767 B.n581 B.n253 163.367
R768 B.n581 B.n251 163.367
R769 B.n585 B.n251 163.367
R770 B.n585 B.n245 163.367
R771 B.n593 B.n245 163.367
R772 B.n593 B.n243 163.367
R773 B.n597 B.n243 163.367
R774 B.n597 B.n238 163.367
R775 B.n606 B.n238 163.367
R776 B.n606 B.n236 163.367
R777 B.n611 B.n236 163.367
R778 B.n611 B.n230 163.367
R779 B.n619 B.n230 163.367
R780 B.n620 B.n619 163.367
R781 B.n620 B.n5 163.367
R782 B.n6 B.n5 163.367
R783 B.n7 B.n6 163.367
R784 B.n626 B.n7 163.367
R785 B.n627 B.n626 163.367
R786 B.n627 B.n13 163.367
R787 B.n14 B.n13 163.367
R788 B.n15 B.n14 163.367
R789 B.n632 B.n15 163.367
R790 B.n632 B.n20 163.367
R791 B.n21 B.n20 163.367
R792 B.n22 B.n21 163.367
R793 B.n637 B.n22 163.367
R794 B.n637 B.n27 163.367
R795 B.n28 B.n27 163.367
R796 B.n29 B.n28 163.367
R797 B.n642 B.n29 163.367
R798 B.n642 B.n34 163.367
R799 B.n35 B.n34 163.367
R800 B.n36 B.n35 163.367
R801 B.n647 B.n36 163.367
R802 B.n647 B.n41 163.367
R803 B.n42 B.n41 163.367
R804 B.n43 B.n42 163.367
R805 B.n652 B.n43 163.367
R806 B.n652 B.n48 163.367
R807 B.n49 B.n48 163.367
R808 B.n50 B.n49 163.367
R809 B.n657 B.n50 163.367
R810 B.n657 B.n55 163.367
R811 B.n56 B.n55 163.367
R812 B.n57 B.n56 163.367
R813 B.n662 B.n57 163.367
R814 B.n662 B.n62 163.367
R815 B.n63 B.n62 163.367
R816 B.n64 B.n63 163.367
R817 B.n667 B.n64 163.367
R818 B.n667 B.n69 163.367
R819 B.n70 B.n69 163.367
R820 B.n71 B.n70 163.367
R821 B.n672 B.n71 163.367
R822 B.n672 B.n76 163.367
R823 B.n77 B.n76 163.367
R824 B.n78 B.n77 163.367
R825 B.n677 B.n78 163.367
R826 B.n677 B.n83 163.367
R827 B.n84 B.n83 163.367
R828 B.n85 B.n84 163.367
R829 B.n682 B.n85 163.367
R830 B.n682 B.n90 163.367
R831 B.n91 B.n90 163.367
R832 B.n92 B.n91 163.367
R833 B.n687 B.n92 163.367
R834 B.n687 B.n97 163.367
R835 B.n363 B.n361 163.367
R836 B.n367 B.n361 163.367
R837 B.n371 B.n369 163.367
R838 B.n375 B.n359 163.367
R839 B.n379 B.n377 163.367
R840 B.n383 B.n357 163.367
R841 B.n387 B.n385 163.367
R842 B.n391 B.n355 163.367
R843 B.n395 B.n393 163.367
R844 B.n399 B.n353 163.367
R845 B.n403 B.n401 163.367
R846 B.n407 B.n348 163.367
R847 B.n411 B.n409 163.367
R848 B.n415 B.n346 163.367
R849 B.n419 B.n417 163.367
R850 B.n424 B.n342 163.367
R851 B.n428 B.n426 163.367
R852 B.n432 B.n340 163.367
R853 B.n436 B.n434 163.367
R854 B.n440 B.n338 163.367
R855 B.n444 B.n442 163.367
R856 B.n448 B.n336 163.367
R857 B.n452 B.n450 163.367
R858 B.n456 B.n334 163.367
R859 B.n459 B.n458 163.367
R860 B.n461 B.n331 163.367
R861 B.n467 B.n327 163.367
R862 B.n471 B.n327 163.367
R863 B.n471 B.n321 163.367
R864 B.n479 B.n321 163.367
R865 B.n479 B.n319 163.367
R866 B.n483 B.n319 163.367
R867 B.n483 B.n313 163.367
R868 B.n491 B.n313 163.367
R869 B.n491 B.n311 163.367
R870 B.n495 B.n311 163.367
R871 B.n495 B.n305 163.367
R872 B.n503 B.n305 163.367
R873 B.n503 B.n303 163.367
R874 B.n507 B.n303 163.367
R875 B.n507 B.n297 163.367
R876 B.n515 B.n297 163.367
R877 B.n515 B.n295 163.367
R878 B.n519 B.n295 163.367
R879 B.n519 B.n289 163.367
R880 B.n527 B.n289 163.367
R881 B.n527 B.n287 163.367
R882 B.n531 B.n287 163.367
R883 B.n531 B.n281 163.367
R884 B.n539 B.n281 163.367
R885 B.n539 B.n279 163.367
R886 B.n543 B.n279 163.367
R887 B.n543 B.n273 163.367
R888 B.n551 B.n273 163.367
R889 B.n551 B.n271 163.367
R890 B.n555 B.n271 163.367
R891 B.n555 B.n265 163.367
R892 B.n563 B.n265 163.367
R893 B.n563 B.n263 163.367
R894 B.n567 B.n263 163.367
R895 B.n567 B.n257 163.367
R896 B.n575 B.n257 163.367
R897 B.n575 B.n255 163.367
R898 B.n579 B.n255 163.367
R899 B.n579 B.n249 163.367
R900 B.n587 B.n249 163.367
R901 B.n587 B.n247 163.367
R902 B.n591 B.n247 163.367
R903 B.n591 B.n241 163.367
R904 B.n600 B.n241 163.367
R905 B.n600 B.n239 163.367
R906 B.n604 B.n239 163.367
R907 B.n604 B.n234 163.367
R908 B.n613 B.n234 163.367
R909 B.n613 B.n232 163.367
R910 B.n617 B.n232 163.367
R911 B.n617 B.n3 163.367
R912 B.n800 B.n3 163.367
R913 B.n796 B.n2 163.367
R914 B.n796 B.n795 163.367
R915 B.n795 B.n9 163.367
R916 B.n791 B.n9 163.367
R917 B.n791 B.n11 163.367
R918 B.n787 B.n11 163.367
R919 B.n787 B.n16 163.367
R920 B.n783 B.n16 163.367
R921 B.n783 B.n18 163.367
R922 B.n779 B.n18 163.367
R923 B.n779 B.n24 163.367
R924 B.n775 B.n24 163.367
R925 B.n775 B.n26 163.367
R926 B.n771 B.n26 163.367
R927 B.n771 B.n31 163.367
R928 B.n767 B.n31 163.367
R929 B.n767 B.n33 163.367
R930 B.n763 B.n33 163.367
R931 B.n763 B.n38 163.367
R932 B.n759 B.n38 163.367
R933 B.n759 B.n40 163.367
R934 B.n755 B.n40 163.367
R935 B.n755 B.n45 163.367
R936 B.n751 B.n45 163.367
R937 B.n751 B.n47 163.367
R938 B.n747 B.n47 163.367
R939 B.n747 B.n52 163.367
R940 B.n743 B.n52 163.367
R941 B.n743 B.n54 163.367
R942 B.n739 B.n54 163.367
R943 B.n739 B.n59 163.367
R944 B.n735 B.n59 163.367
R945 B.n735 B.n61 163.367
R946 B.n731 B.n61 163.367
R947 B.n731 B.n66 163.367
R948 B.n727 B.n66 163.367
R949 B.n727 B.n68 163.367
R950 B.n723 B.n68 163.367
R951 B.n723 B.n73 163.367
R952 B.n719 B.n73 163.367
R953 B.n719 B.n75 163.367
R954 B.n715 B.n75 163.367
R955 B.n715 B.n80 163.367
R956 B.n711 B.n80 163.367
R957 B.n711 B.n82 163.367
R958 B.n707 B.n82 163.367
R959 B.n707 B.n87 163.367
R960 B.n703 B.n87 163.367
R961 B.n703 B.n89 163.367
R962 B.n699 B.n89 163.367
R963 B.n699 B.n94 163.367
R964 B.n695 B.n94 163.367
R965 B.n124 B.t7 148.16
R966 B.n343 B.t18 148.16
R967 B.n126 B.t14 148.155
R968 B.n349 B.t12 148.155
R969 B.n466 B.n330 146.81
R970 B.n694 B.n693 146.81
R971 B.n125 B.t8 74.6564
R972 B.n344 B.t17 74.6564
R973 B.n127 B.t15 74.6516
R974 B.n350 B.t11 74.6516
R975 B.n127 B.n126 73.5035
R976 B.n125 B.n124 73.5035
R977 B.n344 B.n343 73.5035
R978 B.n350 B.n349 73.5035
R979 B.n466 B.n326 72.8695
R980 B.n472 B.n326 72.8695
R981 B.n472 B.n322 72.8695
R982 B.n478 B.n322 72.8695
R983 B.n478 B.n318 72.8695
R984 B.n484 B.n318 72.8695
R985 B.n484 B.n314 72.8695
R986 B.n490 B.n314 72.8695
R987 B.n496 B.n310 72.8695
R988 B.n496 B.n306 72.8695
R989 B.n502 B.n306 72.8695
R990 B.n502 B.n302 72.8695
R991 B.n508 B.n302 72.8695
R992 B.n508 B.n298 72.8695
R993 B.n514 B.n298 72.8695
R994 B.n514 B.n294 72.8695
R995 B.n520 B.n294 72.8695
R996 B.n520 B.n290 72.8695
R997 B.n526 B.n290 72.8695
R998 B.n526 B.n285 72.8695
R999 B.n532 B.n285 72.8695
R1000 B.n532 B.n286 72.8695
R1001 B.n538 B.n278 72.8695
R1002 B.n544 B.n278 72.8695
R1003 B.n544 B.n274 72.8695
R1004 B.n550 B.n274 72.8695
R1005 B.n550 B.n270 72.8695
R1006 B.n556 B.n270 72.8695
R1007 B.n556 B.n266 72.8695
R1008 B.n562 B.n266 72.8695
R1009 B.n562 B.n262 72.8695
R1010 B.n568 B.n262 72.8695
R1011 B.n574 B.n258 72.8695
R1012 B.n574 B.n254 72.8695
R1013 B.n580 B.n254 72.8695
R1014 B.n580 B.n250 72.8695
R1015 B.n586 B.n250 72.8695
R1016 B.n586 B.n246 72.8695
R1017 B.n592 B.n246 72.8695
R1018 B.n592 B.n242 72.8695
R1019 B.n599 B.n242 72.8695
R1020 B.n599 B.n598 72.8695
R1021 B.n605 B.n235 72.8695
R1022 B.n612 B.n235 72.8695
R1023 B.n612 B.n231 72.8695
R1024 B.n618 B.n231 72.8695
R1025 B.n618 B.n4 72.8695
R1026 B.n799 B.n4 72.8695
R1027 B.n799 B.n798 72.8695
R1028 B.n798 B.n797 72.8695
R1029 B.n797 B.n8 72.8695
R1030 B.n12 B.n8 72.8695
R1031 B.n790 B.n12 72.8695
R1032 B.n790 B.n789 72.8695
R1033 B.n789 B.n788 72.8695
R1034 B.n782 B.n19 72.8695
R1035 B.n782 B.n781 72.8695
R1036 B.n781 B.n780 72.8695
R1037 B.n780 B.n23 72.8695
R1038 B.n774 B.n23 72.8695
R1039 B.n774 B.n773 72.8695
R1040 B.n773 B.n772 72.8695
R1041 B.n772 B.n30 72.8695
R1042 B.n766 B.n30 72.8695
R1043 B.n766 B.n765 72.8695
R1044 B.n764 B.n37 72.8695
R1045 B.n758 B.n37 72.8695
R1046 B.n758 B.n757 72.8695
R1047 B.n757 B.n756 72.8695
R1048 B.n756 B.n44 72.8695
R1049 B.n750 B.n44 72.8695
R1050 B.n750 B.n749 72.8695
R1051 B.n749 B.n748 72.8695
R1052 B.n748 B.n51 72.8695
R1053 B.n742 B.n51 72.8695
R1054 B.n741 B.n740 72.8695
R1055 B.n740 B.n58 72.8695
R1056 B.n734 B.n58 72.8695
R1057 B.n734 B.n733 72.8695
R1058 B.n733 B.n732 72.8695
R1059 B.n732 B.n65 72.8695
R1060 B.n726 B.n65 72.8695
R1061 B.n726 B.n725 72.8695
R1062 B.n725 B.n724 72.8695
R1063 B.n724 B.n72 72.8695
R1064 B.n718 B.n72 72.8695
R1065 B.n718 B.n717 72.8695
R1066 B.n717 B.n716 72.8695
R1067 B.n716 B.n79 72.8695
R1068 B.n710 B.n709 72.8695
R1069 B.n709 B.n708 72.8695
R1070 B.n708 B.n86 72.8695
R1071 B.n702 B.n86 72.8695
R1072 B.n702 B.n701 72.8695
R1073 B.n701 B.n700 72.8695
R1074 B.n700 B.n93 72.8695
R1075 B.n694 B.n93 72.8695
R1076 B.n98 B.n96 71.676
R1077 B.n130 B.n99 71.676
R1078 B.n134 B.n100 71.676
R1079 B.n138 B.n101 71.676
R1080 B.n142 B.n102 71.676
R1081 B.n146 B.n103 71.676
R1082 B.n150 B.n104 71.676
R1083 B.n154 B.n105 71.676
R1084 B.n158 B.n106 71.676
R1085 B.n162 B.n107 71.676
R1086 B.n166 B.n108 71.676
R1087 B.n171 B.n109 71.676
R1088 B.n175 B.n110 71.676
R1089 B.n179 B.n111 71.676
R1090 B.n183 B.n112 71.676
R1091 B.n187 B.n113 71.676
R1092 B.n192 B.n114 71.676
R1093 B.n196 B.n115 71.676
R1094 B.n200 B.n116 71.676
R1095 B.n204 B.n117 71.676
R1096 B.n208 B.n118 71.676
R1097 B.n212 B.n119 71.676
R1098 B.n216 B.n120 71.676
R1099 B.n220 B.n121 71.676
R1100 B.n224 B.n122 71.676
R1101 B.n692 B.n123 71.676
R1102 B.n692 B.n691 71.676
R1103 B.n226 B.n122 71.676
R1104 B.n223 B.n121 71.676
R1105 B.n219 B.n120 71.676
R1106 B.n215 B.n119 71.676
R1107 B.n211 B.n118 71.676
R1108 B.n207 B.n117 71.676
R1109 B.n203 B.n116 71.676
R1110 B.n199 B.n115 71.676
R1111 B.n195 B.n114 71.676
R1112 B.n191 B.n113 71.676
R1113 B.n186 B.n112 71.676
R1114 B.n182 B.n111 71.676
R1115 B.n178 B.n110 71.676
R1116 B.n174 B.n109 71.676
R1117 B.n170 B.n108 71.676
R1118 B.n165 B.n107 71.676
R1119 B.n161 B.n106 71.676
R1120 B.n157 B.n105 71.676
R1121 B.n153 B.n104 71.676
R1122 B.n149 B.n103 71.676
R1123 B.n145 B.n102 71.676
R1124 B.n141 B.n101 71.676
R1125 B.n137 B.n100 71.676
R1126 B.n133 B.n99 71.676
R1127 B.n129 B.n98 71.676
R1128 B.n362 B.n329 71.676
R1129 B.n368 B.n367 71.676
R1130 B.n371 B.n370 71.676
R1131 B.n376 B.n375 71.676
R1132 B.n379 B.n378 71.676
R1133 B.n384 B.n383 71.676
R1134 B.n387 B.n386 71.676
R1135 B.n392 B.n391 71.676
R1136 B.n395 B.n394 71.676
R1137 B.n400 B.n399 71.676
R1138 B.n403 B.n402 71.676
R1139 B.n408 B.n407 71.676
R1140 B.n411 B.n410 71.676
R1141 B.n416 B.n415 71.676
R1142 B.n419 B.n418 71.676
R1143 B.n425 B.n424 71.676
R1144 B.n428 B.n427 71.676
R1145 B.n433 B.n432 71.676
R1146 B.n436 B.n435 71.676
R1147 B.n441 B.n440 71.676
R1148 B.n444 B.n443 71.676
R1149 B.n449 B.n448 71.676
R1150 B.n452 B.n451 71.676
R1151 B.n457 B.n456 71.676
R1152 B.n460 B.n459 71.676
R1153 B.n363 B.n362 71.676
R1154 B.n369 B.n368 71.676
R1155 B.n370 B.n359 71.676
R1156 B.n377 B.n376 71.676
R1157 B.n378 B.n357 71.676
R1158 B.n385 B.n384 71.676
R1159 B.n386 B.n355 71.676
R1160 B.n393 B.n392 71.676
R1161 B.n394 B.n353 71.676
R1162 B.n401 B.n400 71.676
R1163 B.n402 B.n348 71.676
R1164 B.n409 B.n408 71.676
R1165 B.n410 B.n346 71.676
R1166 B.n417 B.n416 71.676
R1167 B.n418 B.n342 71.676
R1168 B.n426 B.n425 71.676
R1169 B.n427 B.n340 71.676
R1170 B.n434 B.n433 71.676
R1171 B.n435 B.n338 71.676
R1172 B.n442 B.n441 71.676
R1173 B.n443 B.n336 71.676
R1174 B.n450 B.n449 71.676
R1175 B.n451 B.n334 71.676
R1176 B.n458 B.n457 71.676
R1177 B.n461 B.n460 71.676
R1178 B.n801 B.n800 71.676
R1179 B.n801 B.n2 71.676
R1180 B.n538 B.t2 70.7263
R1181 B.n742 B.t3 70.7263
R1182 B.t0 B.n258 60.0102
R1183 B.n765 B.t19 60.0102
R1184 B.n168 B.n127 59.5399
R1185 B.n189 B.n125 59.5399
R1186 B.n422 B.n344 59.5399
R1187 B.n351 B.n350 59.5399
R1188 B.n490 B.t10 49.2942
R1189 B.n605 B.t4 49.2942
R1190 B.n788 B.t1 49.2942
R1191 B.n710 B.t6 49.2942
R1192 B.n468 B.n328 32.3127
R1193 B.n464 B.n463 32.3127
R1194 B.n690 B.n689 32.3127
R1195 B.n696 B.n95 32.3127
R1196 B.t10 B.n310 23.5758
R1197 B.n598 B.t4 23.5758
R1198 B.n19 B.t1 23.5758
R1199 B.t6 B.n79 23.5758
R1200 B B.n802 18.0485
R1201 B.n568 B.t0 12.8597
R1202 B.t19 B.n764 12.8597
R1203 B.n469 B.n468 10.6151
R1204 B.n470 B.n469 10.6151
R1205 B.n470 B.n320 10.6151
R1206 B.n480 B.n320 10.6151
R1207 B.n481 B.n480 10.6151
R1208 B.n482 B.n481 10.6151
R1209 B.n482 B.n312 10.6151
R1210 B.n492 B.n312 10.6151
R1211 B.n493 B.n492 10.6151
R1212 B.n494 B.n493 10.6151
R1213 B.n494 B.n304 10.6151
R1214 B.n504 B.n304 10.6151
R1215 B.n505 B.n504 10.6151
R1216 B.n506 B.n505 10.6151
R1217 B.n506 B.n296 10.6151
R1218 B.n516 B.n296 10.6151
R1219 B.n517 B.n516 10.6151
R1220 B.n518 B.n517 10.6151
R1221 B.n518 B.n288 10.6151
R1222 B.n528 B.n288 10.6151
R1223 B.n529 B.n528 10.6151
R1224 B.n530 B.n529 10.6151
R1225 B.n530 B.n280 10.6151
R1226 B.n540 B.n280 10.6151
R1227 B.n541 B.n540 10.6151
R1228 B.n542 B.n541 10.6151
R1229 B.n542 B.n272 10.6151
R1230 B.n552 B.n272 10.6151
R1231 B.n553 B.n552 10.6151
R1232 B.n554 B.n553 10.6151
R1233 B.n554 B.n264 10.6151
R1234 B.n564 B.n264 10.6151
R1235 B.n565 B.n564 10.6151
R1236 B.n566 B.n565 10.6151
R1237 B.n566 B.n256 10.6151
R1238 B.n576 B.n256 10.6151
R1239 B.n577 B.n576 10.6151
R1240 B.n578 B.n577 10.6151
R1241 B.n578 B.n248 10.6151
R1242 B.n588 B.n248 10.6151
R1243 B.n589 B.n588 10.6151
R1244 B.n590 B.n589 10.6151
R1245 B.n590 B.n240 10.6151
R1246 B.n601 B.n240 10.6151
R1247 B.n602 B.n601 10.6151
R1248 B.n603 B.n602 10.6151
R1249 B.n603 B.n233 10.6151
R1250 B.n614 B.n233 10.6151
R1251 B.n615 B.n614 10.6151
R1252 B.n616 B.n615 10.6151
R1253 B.n616 B.n0 10.6151
R1254 B.n364 B.n328 10.6151
R1255 B.n365 B.n364 10.6151
R1256 B.n366 B.n365 10.6151
R1257 B.n366 B.n360 10.6151
R1258 B.n372 B.n360 10.6151
R1259 B.n373 B.n372 10.6151
R1260 B.n374 B.n373 10.6151
R1261 B.n374 B.n358 10.6151
R1262 B.n380 B.n358 10.6151
R1263 B.n381 B.n380 10.6151
R1264 B.n382 B.n381 10.6151
R1265 B.n382 B.n356 10.6151
R1266 B.n388 B.n356 10.6151
R1267 B.n389 B.n388 10.6151
R1268 B.n390 B.n389 10.6151
R1269 B.n390 B.n354 10.6151
R1270 B.n396 B.n354 10.6151
R1271 B.n397 B.n396 10.6151
R1272 B.n398 B.n397 10.6151
R1273 B.n398 B.n352 10.6151
R1274 B.n405 B.n404 10.6151
R1275 B.n406 B.n405 10.6151
R1276 B.n406 B.n347 10.6151
R1277 B.n412 B.n347 10.6151
R1278 B.n413 B.n412 10.6151
R1279 B.n414 B.n413 10.6151
R1280 B.n414 B.n345 10.6151
R1281 B.n420 B.n345 10.6151
R1282 B.n421 B.n420 10.6151
R1283 B.n423 B.n341 10.6151
R1284 B.n429 B.n341 10.6151
R1285 B.n430 B.n429 10.6151
R1286 B.n431 B.n430 10.6151
R1287 B.n431 B.n339 10.6151
R1288 B.n437 B.n339 10.6151
R1289 B.n438 B.n437 10.6151
R1290 B.n439 B.n438 10.6151
R1291 B.n439 B.n337 10.6151
R1292 B.n445 B.n337 10.6151
R1293 B.n446 B.n445 10.6151
R1294 B.n447 B.n446 10.6151
R1295 B.n447 B.n335 10.6151
R1296 B.n453 B.n335 10.6151
R1297 B.n454 B.n453 10.6151
R1298 B.n455 B.n454 10.6151
R1299 B.n455 B.n333 10.6151
R1300 B.n333 B.n332 10.6151
R1301 B.n462 B.n332 10.6151
R1302 B.n463 B.n462 10.6151
R1303 B.n464 B.n324 10.6151
R1304 B.n474 B.n324 10.6151
R1305 B.n475 B.n474 10.6151
R1306 B.n476 B.n475 10.6151
R1307 B.n476 B.n316 10.6151
R1308 B.n486 B.n316 10.6151
R1309 B.n487 B.n486 10.6151
R1310 B.n488 B.n487 10.6151
R1311 B.n488 B.n308 10.6151
R1312 B.n498 B.n308 10.6151
R1313 B.n499 B.n498 10.6151
R1314 B.n500 B.n499 10.6151
R1315 B.n500 B.n300 10.6151
R1316 B.n510 B.n300 10.6151
R1317 B.n511 B.n510 10.6151
R1318 B.n512 B.n511 10.6151
R1319 B.n512 B.n292 10.6151
R1320 B.n522 B.n292 10.6151
R1321 B.n523 B.n522 10.6151
R1322 B.n524 B.n523 10.6151
R1323 B.n524 B.n283 10.6151
R1324 B.n534 B.n283 10.6151
R1325 B.n535 B.n534 10.6151
R1326 B.n536 B.n535 10.6151
R1327 B.n536 B.n276 10.6151
R1328 B.n546 B.n276 10.6151
R1329 B.n547 B.n546 10.6151
R1330 B.n548 B.n547 10.6151
R1331 B.n548 B.n268 10.6151
R1332 B.n558 B.n268 10.6151
R1333 B.n559 B.n558 10.6151
R1334 B.n560 B.n559 10.6151
R1335 B.n560 B.n260 10.6151
R1336 B.n570 B.n260 10.6151
R1337 B.n571 B.n570 10.6151
R1338 B.n572 B.n571 10.6151
R1339 B.n572 B.n252 10.6151
R1340 B.n582 B.n252 10.6151
R1341 B.n583 B.n582 10.6151
R1342 B.n584 B.n583 10.6151
R1343 B.n584 B.n244 10.6151
R1344 B.n594 B.n244 10.6151
R1345 B.n595 B.n594 10.6151
R1346 B.n596 B.n595 10.6151
R1347 B.n596 B.n237 10.6151
R1348 B.n607 B.n237 10.6151
R1349 B.n608 B.n607 10.6151
R1350 B.n610 B.n608 10.6151
R1351 B.n610 B.n609 10.6151
R1352 B.n609 B.n229 10.6151
R1353 B.n621 B.n229 10.6151
R1354 B.n622 B.n621 10.6151
R1355 B.n623 B.n622 10.6151
R1356 B.n624 B.n623 10.6151
R1357 B.n625 B.n624 10.6151
R1358 B.n628 B.n625 10.6151
R1359 B.n629 B.n628 10.6151
R1360 B.n630 B.n629 10.6151
R1361 B.n631 B.n630 10.6151
R1362 B.n633 B.n631 10.6151
R1363 B.n634 B.n633 10.6151
R1364 B.n635 B.n634 10.6151
R1365 B.n636 B.n635 10.6151
R1366 B.n638 B.n636 10.6151
R1367 B.n639 B.n638 10.6151
R1368 B.n640 B.n639 10.6151
R1369 B.n641 B.n640 10.6151
R1370 B.n643 B.n641 10.6151
R1371 B.n644 B.n643 10.6151
R1372 B.n645 B.n644 10.6151
R1373 B.n646 B.n645 10.6151
R1374 B.n648 B.n646 10.6151
R1375 B.n649 B.n648 10.6151
R1376 B.n650 B.n649 10.6151
R1377 B.n651 B.n650 10.6151
R1378 B.n653 B.n651 10.6151
R1379 B.n654 B.n653 10.6151
R1380 B.n655 B.n654 10.6151
R1381 B.n656 B.n655 10.6151
R1382 B.n658 B.n656 10.6151
R1383 B.n659 B.n658 10.6151
R1384 B.n660 B.n659 10.6151
R1385 B.n661 B.n660 10.6151
R1386 B.n663 B.n661 10.6151
R1387 B.n664 B.n663 10.6151
R1388 B.n665 B.n664 10.6151
R1389 B.n666 B.n665 10.6151
R1390 B.n668 B.n666 10.6151
R1391 B.n669 B.n668 10.6151
R1392 B.n670 B.n669 10.6151
R1393 B.n671 B.n670 10.6151
R1394 B.n673 B.n671 10.6151
R1395 B.n674 B.n673 10.6151
R1396 B.n675 B.n674 10.6151
R1397 B.n676 B.n675 10.6151
R1398 B.n678 B.n676 10.6151
R1399 B.n679 B.n678 10.6151
R1400 B.n680 B.n679 10.6151
R1401 B.n681 B.n680 10.6151
R1402 B.n683 B.n681 10.6151
R1403 B.n684 B.n683 10.6151
R1404 B.n685 B.n684 10.6151
R1405 B.n686 B.n685 10.6151
R1406 B.n688 B.n686 10.6151
R1407 B.n689 B.n688 10.6151
R1408 B.n794 B.n1 10.6151
R1409 B.n794 B.n793 10.6151
R1410 B.n793 B.n792 10.6151
R1411 B.n792 B.n10 10.6151
R1412 B.n786 B.n10 10.6151
R1413 B.n786 B.n785 10.6151
R1414 B.n785 B.n784 10.6151
R1415 B.n784 B.n17 10.6151
R1416 B.n778 B.n17 10.6151
R1417 B.n778 B.n777 10.6151
R1418 B.n777 B.n776 10.6151
R1419 B.n776 B.n25 10.6151
R1420 B.n770 B.n25 10.6151
R1421 B.n770 B.n769 10.6151
R1422 B.n769 B.n768 10.6151
R1423 B.n768 B.n32 10.6151
R1424 B.n762 B.n32 10.6151
R1425 B.n762 B.n761 10.6151
R1426 B.n761 B.n760 10.6151
R1427 B.n760 B.n39 10.6151
R1428 B.n754 B.n39 10.6151
R1429 B.n754 B.n753 10.6151
R1430 B.n753 B.n752 10.6151
R1431 B.n752 B.n46 10.6151
R1432 B.n746 B.n46 10.6151
R1433 B.n746 B.n745 10.6151
R1434 B.n745 B.n744 10.6151
R1435 B.n744 B.n53 10.6151
R1436 B.n738 B.n53 10.6151
R1437 B.n738 B.n737 10.6151
R1438 B.n737 B.n736 10.6151
R1439 B.n736 B.n60 10.6151
R1440 B.n730 B.n60 10.6151
R1441 B.n730 B.n729 10.6151
R1442 B.n729 B.n728 10.6151
R1443 B.n728 B.n67 10.6151
R1444 B.n722 B.n67 10.6151
R1445 B.n722 B.n721 10.6151
R1446 B.n721 B.n720 10.6151
R1447 B.n720 B.n74 10.6151
R1448 B.n714 B.n74 10.6151
R1449 B.n714 B.n713 10.6151
R1450 B.n713 B.n712 10.6151
R1451 B.n712 B.n81 10.6151
R1452 B.n706 B.n81 10.6151
R1453 B.n706 B.n705 10.6151
R1454 B.n705 B.n704 10.6151
R1455 B.n704 B.n88 10.6151
R1456 B.n698 B.n88 10.6151
R1457 B.n698 B.n697 10.6151
R1458 B.n697 B.n696 10.6151
R1459 B.n128 B.n95 10.6151
R1460 B.n131 B.n128 10.6151
R1461 B.n132 B.n131 10.6151
R1462 B.n135 B.n132 10.6151
R1463 B.n136 B.n135 10.6151
R1464 B.n139 B.n136 10.6151
R1465 B.n140 B.n139 10.6151
R1466 B.n143 B.n140 10.6151
R1467 B.n144 B.n143 10.6151
R1468 B.n147 B.n144 10.6151
R1469 B.n148 B.n147 10.6151
R1470 B.n151 B.n148 10.6151
R1471 B.n152 B.n151 10.6151
R1472 B.n155 B.n152 10.6151
R1473 B.n156 B.n155 10.6151
R1474 B.n159 B.n156 10.6151
R1475 B.n160 B.n159 10.6151
R1476 B.n163 B.n160 10.6151
R1477 B.n164 B.n163 10.6151
R1478 B.n167 B.n164 10.6151
R1479 B.n172 B.n169 10.6151
R1480 B.n173 B.n172 10.6151
R1481 B.n176 B.n173 10.6151
R1482 B.n177 B.n176 10.6151
R1483 B.n180 B.n177 10.6151
R1484 B.n181 B.n180 10.6151
R1485 B.n184 B.n181 10.6151
R1486 B.n185 B.n184 10.6151
R1487 B.n188 B.n185 10.6151
R1488 B.n193 B.n190 10.6151
R1489 B.n194 B.n193 10.6151
R1490 B.n197 B.n194 10.6151
R1491 B.n198 B.n197 10.6151
R1492 B.n201 B.n198 10.6151
R1493 B.n202 B.n201 10.6151
R1494 B.n205 B.n202 10.6151
R1495 B.n206 B.n205 10.6151
R1496 B.n209 B.n206 10.6151
R1497 B.n210 B.n209 10.6151
R1498 B.n213 B.n210 10.6151
R1499 B.n214 B.n213 10.6151
R1500 B.n217 B.n214 10.6151
R1501 B.n218 B.n217 10.6151
R1502 B.n221 B.n218 10.6151
R1503 B.n222 B.n221 10.6151
R1504 B.n225 B.n222 10.6151
R1505 B.n227 B.n225 10.6151
R1506 B.n228 B.n227 10.6151
R1507 B.n690 B.n228 10.6151
R1508 B.n352 B.n351 9.36635
R1509 B.n423 B.n422 9.36635
R1510 B.n168 B.n167 9.36635
R1511 B.n190 B.n189 9.36635
R1512 B.n802 B.n0 8.11757
R1513 B.n802 B.n1 8.11757
R1514 B.n286 B.t2 2.14371
R1515 B.t3 B.n741 2.14371
R1516 B.n404 B.n351 1.24928
R1517 B.n422 B.n421 1.24928
R1518 B.n169 B.n168 1.24928
R1519 B.n189 B.n188 1.24928
R1520 VN.n34 VN.n33 161.3
R1521 VN.n32 VN.n19 161.3
R1522 VN.n31 VN.n30 161.3
R1523 VN.n29 VN.n20 161.3
R1524 VN.n28 VN.n27 161.3
R1525 VN.n26 VN.n21 161.3
R1526 VN.n25 VN.n24 161.3
R1527 VN.n16 VN.n15 161.3
R1528 VN.n14 VN.n1 161.3
R1529 VN.n13 VN.n12 161.3
R1530 VN.n11 VN.n2 161.3
R1531 VN.n10 VN.n9 161.3
R1532 VN.n8 VN.n3 161.3
R1533 VN.n7 VN.n6 161.3
R1534 VN.n17 VN.n0 75.8765
R1535 VN.n35 VN.n18 75.8765
R1536 VN.n23 VN.t3 68.7832
R1537 VN.n5 VN.t4 68.7832
R1538 VN.n9 VN.n2 50.6917
R1539 VN.n27 VN.n20 50.6917
R1540 VN.n23 VN.n22 50.1886
R1541 VN.n5 VN.n4 50.1886
R1542 VN VN.n35 47.0473
R1543 VN.n4 VN.t2 34.7574
R1544 VN.n0 VN.t1 34.7574
R1545 VN.n22 VN.t5 34.7574
R1546 VN.n18 VN.t0 34.7574
R1547 VN.n13 VN.n2 30.2951
R1548 VN.n31 VN.n20 30.2951
R1549 VN.n7 VN.n4 24.4675
R1550 VN.n8 VN.n7 24.4675
R1551 VN.n9 VN.n8 24.4675
R1552 VN.n14 VN.n13 24.4675
R1553 VN.n15 VN.n14 24.4675
R1554 VN.n27 VN.n26 24.4675
R1555 VN.n26 VN.n25 24.4675
R1556 VN.n25 VN.n22 24.4675
R1557 VN.n33 VN.n32 24.4675
R1558 VN.n32 VN.n31 24.4675
R1559 VN.n15 VN.n0 14.1914
R1560 VN.n33 VN.n18 14.1914
R1561 VN.n24 VN.n23 3.01037
R1562 VN.n6 VN.n5 3.01037
R1563 VN.n35 VN.n34 0.354971
R1564 VN.n17 VN.n16 0.354971
R1565 VN VN.n17 0.26696
R1566 VN.n34 VN.n19 0.189894
R1567 VN.n30 VN.n19 0.189894
R1568 VN.n30 VN.n29 0.189894
R1569 VN.n29 VN.n28 0.189894
R1570 VN.n28 VN.n21 0.189894
R1571 VN.n24 VN.n21 0.189894
R1572 VN.n6 VN.n3 0.189894
R1573 VN.n10 VN.n3 0.189894
R1574 VN.n11 VN.n10 0.189894
R1575 VN.n12 VN.n11 0.189894
R1576 VN.n12 VN.n1 0.189894
R1577 VN.n16 VN.n1 0.189894
R1578 VDD2.n1 VDD2.t1 77.2875
R1579 VDD2.n2 VDD2.t5 74.8925
R1580 VDD2.n1 VDD2.n0 71.6859
R1581 VDD2 VDD2.n3 71.6831
R1582 VDD2.n2 VDD2.n1 38.6356
R1583 VDD2.n3 VDD2.t0 3.96844
R1584 VDD2.n3 VDD2.t2 3.96844
R1585 VDD2.n0 VDD2.t3 3.96844
R1586 VDD2.n0 VDD2.t4 3.96844
R1587 VDD2 VDD2.n2 2.50912
C0 VDD2 VN 3.16956f
C1 VTAIL VN 4.06428f
C2 VDD1 VN 0.151894f
C3 VN VP 6.463089f
C4 VDD2 VTAIL 5.76414f
C5 VDD2 VDD1 1.74174f
C6 VDD2 VP 0.535032f
C7 VDD1 VTAIL 5.70559f
C8 VTAIL VP 4.07844f
C9 VDD1 VP 3.54624f
C10 VDD2 B 5.400996f
C11 VDD1 B 5.757774f
C12 VTAIL B 5.111527f
C13 VN B 14.761749f
C14 VP B 13.426101f
C15 VDD2.t1 B 0.917402f
C16 VDD2.t3 B 0.087468f
C17 VDD2.t4 B 0.087468f
C18 VDD2.n0 B 0.717147f
C19 VDD2.n1 B 2.50757f
C20 VDD2.t5 B 0.904928f
C21 VDD2.n2 B 2.18416f
C22 VDD2.t0 B 0.087468f
C23 VDD2.t2 B 0.087468f
C24 VDD2.n3 B 0.717118f
C25 VN.t1 B 1.0621f
C26 VN.n0 B 0.496907f
C27 VN.n1 B 0.023522f
C28 VN.n2 B 0.022573f
C29 VN.n3 B 0.023522f
C30 VN.t2 B 1.0621f
C31 VN.n4 B 0.494538f
C32 VN.t4 B 1.34876f
C33 VN.n5 B 0.466997f
C34 VN.n6 B 0.287251f
C35 VN.n7 B 0.043839f
C36 VN.n8 B 0.043839f
C37 VN.n9 B 0.042943f
C38 VN.n10 B 0.023522f
C39 VN.n11 B 0.023522f
C40 VN.n12 B 0.023522f
C41 VN.n13 B 0.047003f
C42 VN.n14 B 0.043839f
C43 VN.n15 B 0.034749f
C44 VN.n16 B 0.037964f
C45 VN.n17 B 0.05895f
C46 VN.t0 B 1.0621f
C47 VN.n18 B 0.496907f
C48 VN.n19 B 0.023522f
C49 VN.n20 B 0.022573f
C50 VN.n21 B 0.023522f
C51 VN.t5 B 1.0621f
C52 VN.n22 B 0.494538f
C53 VN.t3 B 1.34876f
C54 VN.n23 B 0.466997f
C55 VN.n24 B 0.287251f
C56 VN.n25 B 0.043839f
C57 VN.n26 B 0.043839f
C58 VN.n27 B 0.042943f
C59 VN.n28 B 0.023522f
C60 VN.n29 B 0.023522f
C61 VN.n30 B 0.023522f
C62 VN.n31 B 0.047003f
C63 VN.n32 B 0.043839f
C64 VN.n33 B 0.034749f
C65 VN.n34 B 0.037964f
C66 VN.n35 B 1.23127f
C67 VDD1.t4 B 0.930172f
C68 VDD1.t1 B 0.929329f
C69 VDD1.t3 B 0.088605f
C70 VDD1.t2 B 0.088605f
C71 VDD1.n0 B 0.72647f
C72 VDD1.n1 B 2.66531f
C73 VDD1.t0 B 0.088605f
C74 VDD1.t5 B 0.088605f
C75 VDD1.n2 B 0.721367f
C76 VDD1.n3 B 2.23394f
C77 VTAIL.t1 B 0.116205f
C78 VTAIL.t11 B 0.116205f
C79 VTAIL.n0 B 0.875658f
C80 VTAIL.n1 B 0.547806f
C81 VTAIL.t9 B 1.11921f
C82 VTAIL.n2 B 0.848335f
C83 VTAIL.t10 B 0.116205f
C84 VTAIL.t8 B 0.116205f
C85 VTAIL.n3 B 0.875658f
C86 VTAIL.n4 B 2.00451f
C87 VTAIL.t2 B 0.116205f
C88 VTAIL.t0 B 0.116205f
C89 VTAIL.n5 B 0.875663f
C90 VTAIL.n6 B 2.0045f
C91 VTAIL.t4 B 1.11922f
C92 VTAIL.n7 B 0.848328f
C93 VTAIL.t7 B 0.116205f
C94 VTAIL.t5 B 0.116205f
C95 VTAIL.n8 B 0.875663f
C96 VTAIL.n9 B 0.774961f
C97 VTAIL.t6 B 1.11921f
C98 VTAIL.n10 B 1.76763f
C99 VTAIL.t3 B 1.11921f
C100 VTAIL.n11 B 1.68454f
C101 VP.t3 B 1.08779f
C102 VP.n0 B 0.508929f
C103 VP.n1 B 0.024091f
C104 VP.n2 B 0.023119f
C105 VP.n3 B 0.024091f
C106 VP.t2 B 1.08779f
C107 VP.n4 B 0.433453f
C108 VP.n5 B 0.024091f
C109 VP.n6 B 0.023119f
C110 VP.n7 B 0.024091f
C111 VP.t4 B 1.08779f
C112 VP.n8 B 0.508929f
C113 VP.t0 B 1.08779f
C114 VP.n9 B 0.508929f
C115 VP.n10 B 0.024091f
C116 VP.n11 B 0.023119f
C117 VP.n12 B 0.024091f
C118 VP.t5 B 1.08779f
C119 VP.n13 B 0.506503f
C120 VP.t1 B 1.38139f
C121 VP.n14 B 0.478296f
C122 VP.n15 B 0.294201f
C123 VP.n16 B 0.0449f
C124 VP.n17 B 0.0449f
C125 VP.n18 B 0.043982f
C126 VP.n19 B 0.024091f
C127 VP.n20 B 0.024091f
C128 VP.n21 B 0.024091f
C129 VP.n22 B 0.04814f
C130 VP.n23 B 0.0449f
C131 VP.n24 B 0.035589f
C132 VP.n25 B 0.038882f
C133 VP.n26 B 1.25098f
C134 VP.n27 B 1.26946f
C135 VP.n28 B 0.038882f
C136 VP.n29 B 0.035589f
C137 VP.n30 B 0.0449f
C138 VP.n31 B 0.04814f
C139 VP.n32 B 0.024091f
C140 VP.n33 B 0.024091f
C141 VP.n34 B 0.024091f
C142 VP.n35 B 0.043982f
C143 VP.n36 B 0.0449f
C144 VP.n37 B 0.0449f
C145 VP.n38 B 0.024091f
C146 VP.n39 B 0.024091f
C147 VP.n40 B 0.024091f
C148 VP.n41 B 0.0449f
C149 VP.n42 B 0.0449f
C150 VP.n43 B 0.043982f
C151 VP.n44 B 0.024091f
C152 VP.n45 B 0.024091f
C153 VP.n46 B 0.024091f
C154 VP.n47 B 0.04814f
C155 VP.n48 B 0.0449f
C156 VP.n49 B 0.035589f
C157 VP.n50 B 0.038882f
C158 VP.n51 B 0.060376f
.ends

