* NGSPICE file created from diff_pair_sample_0427.ext - technology: sky130A

.subckt diff_pair_sample_0427 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=1.32825 ps=8.38 w=8.05 l=0.31
X1 VDD1.t2 VP.t1 VTAIL.t6 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=1.32825 pd=8.38 as=3.1395 ps=16.88 w=8.05 l=0.31
X2 B.t11 B.t9 B.t10 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=0 ps=0 w=8.05 l=0.31
X3 VDD1.t3 VP.t2 VTAIL.t5 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=1.32825 pd=8.38 as=3.1395 ps=16.88 w=8.05 l=0.31
X4 VTAIL.t0 VN.t0 VDD2.t3 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=1.32825 ps=8.38 w=8.05 l=0.31
X5 B.t8 B.t6 B.t7 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=0 ps=0 w=8.05 l=0.31
X6 B.t5 B.t3 B.t4 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=0 ps=0 w=8.05 l=0.31
X7 VDD2.t2 VN.t1 VTAIL.t3 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=1.32825 pd=8.38 as=3.1395 ps=16.88 w=8.05 l=0.31
X8 VTAIL.t4 VP.t3 VDD1.t0 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=1.32825 ps=8.38 w=8.05 l=0.31
X9 B.t2 B.t0 B.t1 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=0 ps=0 w=8.05 l=0.31
X10 VTAIL.t2 VN.t2 VDD2.t1 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=3.1395 pd=16.88 as=1.32825 ps=8.38 w=8.05 l=0.31
X11 VDD2.t0 VN.t3 VTAIL.t1 w_n1354_n2582# sky130_fd_pr__pfet_01v8 ad=1.32825 pd=8.38 as=3.1395 ps=16.88 w=8.05 l=0.31
R0 VP.n1 VP.t1 774.404
R1 VP.n1 VP.t0 774.404
R2 VP.n0 VP.t3 774.404
R3 VP.n0 VP.t2 774.404
R4 VP.n2 VP.n0 197.633
R5 VP.n2 VP.n1 161.3
R6 VP VP.n2 0.0516364
R7 VDD1 VDD1.n1 113.505
R8 VDD1 VDD1.n0 80.7118
R9 VDD1.n0 VDD1.t0 4.03839
R10 VDD1.n0 VDD1.t3 4.03839
R11 VDD1.n1 VDD1.t1 4.03839
R12 VDD1.n1 VDD1.t2 4.03839
R13 VTAIL.n346 VTAIL.n308 756.745
R14 VTAIL.n38 VTAIL.n0 756.745
R15 VTAIL.n82 VTAIL.n44 756.745
R16 VTAIL.n126 VTAIL.n88 756.745
R17 VTAIL.n302 VTAIL.n264 756.745
R18 VTAIL.n258 VTAIL.n220 756.745
R19 VTAIL.n214 VTAIL.n176 756.745
R20 VTAIL.n170 VTAIL.n132 756.745
R21 VTAIL.n323 VTAIL.n322 585
R22 VTAIL.n320 VTAIL.n319 585
R23 VTAIL.n329 VTAIL.n328 585
R24 VTAIL.n331 VTAIL.n330 585
R25 VTAIL.n316 VTAIL.n315 585
R26 VTAIL.n337 VTAIL.n336 585
R27 VTAIL.n339 VTAIL.n338 585
R28 VTAIL.n312 VTAIL.n311 585
R29 VTAIL.n345 VTAIL.n344 585
R30 VTAIL.n347 VTAIL.n346 585
R31 VTAIL.n15 VTAIL.n14 585
R32 VTAIL.n12 VTAIL.n11 585
R33 VTAIL.n21 VTAIL.n20 585
R34 VTAIL.n23 VTAIL.n22 585
R35 VTAIL.n8 VTAIL.n7 585
R36 VTAIL.n29 VTAIL.n28 585
R37 VTAIL.n31 VTAIL.n30 585
R38 VTAIL.n4 VTAIL.n3 585
R39 VTAIL.n37 VTAIL.n36 585
R40 VTAIL.n39 VTAIL.n38 585
R41 VTAIL.n59 VTAIL.n58 585
R42 VTAIL.n56 VTAIL.n55 585
R43 VTAIL.n65 VTAIL.n64 585
R44 VTAIL.n67 VTAIL.n66 585
R45 VTAIL.n52 VTAIL.n51 585
R46 VTAIL.n73 VTAIL.n72 585
R47 VTAIL.n75 VTAIL.n74 585
R48 VTAIL.n48 VTAIL.n47 585
R49 VTAIL.n81 VTAIL.n80 585
R50 VTAIL.n83 VTAIL.n82 585
R51 VTAIL.n103 VTAIL.n102 585
R52 VTAIL.n100 VTAIL.n99 585
R53 VTAIL.n109 VTAIL.n108 585
R54 VTAIL.n111 VTAIL.n110 585
R55 VTAIL.n96 VTAIL.n95 585
R56 VTAIL.n117 VTAIL.n116 585
R57 VTAIL.n119 VTAIL.n118 585
R58 VTAIL.n92 VTAIL.n91 585
R59 VTAIL.n125 VTAIL.n124 585
R60 VTAIL.n127 VTAIL.n126 585
R61 VTAIL.n303 VTAIL.n302 585
R62 VTAIL.n301 VTAIL.n300 585
R63 VTAIL.n268 VTAIL.n267 585
R64 VTAIL.n295 VTAIL.n294 585
R65 VTAIL.n293 VTAIL.n292 585
R66 VTAIL.n272 VTAIL.n271 585
R67 VTAIL.n287 VTAIL.n286 585
R68 VTAIL.n285 VTAIL.n284 585
R69 VTAIL.n276 VTAIL.n275 585
R70 VTAIL.n279 VTAIL.n278 585
R71 VTAIL.n259 VTAIL.n258 585
R72 VTAIL.n257 VTAIL.n256 585
R73 VTAIL.n224 VTAIL.n223 585
R74 VTAIL.n251 VTAIL.n250 585
R75 VTAIL.n249 VTAIL.n248 585
R76 VTAIL.n228 VTAIL.n227 585
R77 VTAIL.n243 VTAIL.n242 585
R78 VTAIL.n241 VTAIL.n240 585
R79 VTAIL.n232 VTAIL.n231 585
R80 VTAIL.n235 VTAIL.n234 585
R81 VTAIL.n215 VTAIL.n214 585
R82 VTAIL.n213 VTAIL.n212 585
R83 VTAIL.n180 VTAIL.n179 585
R84 VTAIL.n207 VTAIL.n206 585
R85 VTAIL.n205 VTAIL.n204 585
R86 VTAIL.n184 VTAIL.n183 585
R87 VTAIL.n199 VTAIL.n198 585
R88 VTAIL.n197 VTAIL.n196 585
R89 VTAIL.n188 VTAIL.n187 585
R90 VTAIL.n191 VTAIL.n190 585
R91 VTAIL.n171 VTAIL.n170 585
R92 VTAIL.n169 VTAIL.n168 585
R93 VTAIL.n136 VTAIL.n135 585
R94 VTAIL.n163 VTAIL.n162 585
R95 VTAIL.n161 VTAIL.n160 585
R96 VTAIL.n140 VTAIL.n139 585
R97 VTAIL.n155 VTAIL.n154 585
R98 VTAIL.n153 VTAIL.n152 585
R99 VTAIL.n144 VTAIL.n143 585
R100 VTAIL.n147 VTAIL.n146 585
R101 VTAIL.t3 VTAIL.n321 327.473
R102 VTAIL.t2 VTAIL.n13 327.473
R103 VTAIL.t6 VTAIL.n57 327.473
R104 VTAIL.t7 VTAIL.n101 327.473
R105 VTAIL.t5 VTAIL.n277 327.473
R106 VTAIL.t4 VTAIL.n233 327.473
R107 VTAIL.t1 VTAIL.n189 327.473
R108 VTAIL.t0 VTAIL.n145 327.473
R109 VTAIL.n322 VTAIL.n319 171.744
R110 VTAIL.n329 VTAIL.n319 171.744
R111 VTAIL.n330 VTAIL.n329 171.744
R112 VTAIL.n330 VTAIL.n315 171.744
R113 VTAIL.n337 VTAIL.n315 171.744
R114 VTAIL.n338 VTAIL.n337 171.744
R115 VTAIL.n338 VTAIL.n311 171.744
R116 VTAIL.n345 VTAIL.n311 171.744
R117 VTAIL.n346 VTAIL.n345 171.744
R118 VTAIL.n14 VTAIL.n11 171.744
R119 VTAIL.n21 VTAIL.n11 171.744
R120 VTAIL.n22 VTAIL.n21 171.744
R121 VTAIL.n22 VTAIL.n7 171.744
R122 VTAIL.n29 VTAIL.n7 171.744
R123 VTAIL.n30 VTAIL.n29 171.744
R124 VTAIL.n30 VTAIL.n3 171.744
R125 VTAIL.n37 VTAIL.n3 171.744
R126 VTAIL.n38 VTAIL.n37 171.744
R127 VTAIL.n58 VTAIL.n55 171.744
R128 VTAIL.n65 VTAIL.n55 171.744
R129 VTAIL.n66 VTAIL.n65 171.744
R130 VTAIL.n66 VTAIL.n51 171.744
R131 VTAIL.n73 VTAIL.n51 171.744
R132 VTAIL.n74 VTAIL.n73 171.744
R133 VTAIL.n74 VTAIL.n47 171.744
R134 VTAIL.n81 VTAIL.n47 171.744
R135 VTAIL.n82 VTAIL.n81 171.744
R136 VTAIL.n102 VTAIL.n99 171.744
R137 VTAIL.n109 VTAIL.n99 171.744
R138 VTAIL.n110 VTAIL.n109 171.744
R139 VTAIL.n110 VTAIL.n95 171.744
R140 VTAIL.n117 VTAIL.n95 171.744
R141 VTAIL.n118 VTAIL.n117 171.744
R142 VTAIL.n118 VTAIL.n91 171.744
R143 VTAIL.n125 VTAIL.n91 171.744
R144 VTAIL.n126 VTAIL.n125 171.744
R145 VTAIL.n302 VTAIL.n301 171.744
R146 VTAIL.n301 VTAIL.n267 171.744
R147 VTAIL.n294 VTAIL.n267 171.744
R148 VTAIL.n294 VTAIL.n293 171.744
R149 VTAIL.n293 VTAIL.n271 171.744
R150 VTAIL.n286 VTAIL.n271 171.744
R151 VTAIL.n286 VTAIL.n285 171.744
R152 VTAIL.n285 VTAIL.n275 171.744
R153 VTAIL.n278 VTAIL.n275 171.744
R154 VTAIL.n258 VTAIL.n257 171.744
R155 VTAIL.n257 VTAIL.n223 171.744
R156 VTAIL.n250 VTAIL.n223 171.744
R157 VTAIL.n250 VTAIL.n249 171.744
R158 VTAIL.n249 VTAIL.n227 171.744
R159 VTAIL.n242 VTAIL.n227 171.744
R160 VTAIL.n242 VTAIL.n241 171.744
R161 VTAIL.n241 VTAIL.n231 171.744
R162 VTAIL.n234 VTAIL.n231 171.744
R163 VTAIL.n214 VTAIL.n213 171.744
R164 VTAIL.n213 VTAIL.n179 171.744
R165 VTAIL.n206 VTAIL.n179 171.744
R166 VTAIL.n206 VTAIL.n205 171.744
R167 VTAIL.n205 VTAIL.n183 171.744
R168 VTAIL.n198 VTAIL.n183 171.744
R169 VTAIL.n198 VTAIL.n197 171.744
R170 VTAIL.n197 VTAIL.n187 171.744
R171 VTAIL.n190 VTAIL.n187 171.744
R172 VTAIL.n170 VTAIL.n169 171.744
R173 VTAIL.n169 VTAIL.n135 171.744
R174 VTAIL.n162 VTAIL.n135 171.744
R175 VTAIL.n162 VTAIL.n161 171.744
R176 VTAIL.n161 VTAIL.n139 171.744
R177 VTAIL.n154 VTAIL.n139 171.744
R178 VTAIL.n154 VTAIL.n153 171.744
R179 VTAIL.n153 VTAIL.n143 171.744
R180 VTAIL.n146 VTAIL.n143 171.744
R181 VTAIL.n322 VTAIL.t3 85.8723
R182 VTAIL.n14 VTAIL.t2 85.8723
R183 VTAIL.n58 VTAIL.t6 85.8723
R184 VTAIL.n102 VTAIL.t7 85.8723
R185 VTAIL.n278 VTAIL.t5 85.8723
R186 VTAIL.n234 VTAIL.t4 85.8723
R187 VTAIL.n190 VTAIL.t1 85.8723
R188 VTAIL.n146 VTAIL.t0 85.8723
R189 VTAIL.n351 VTAIL.n350 30.052
R190 VTAIL.n43 VTAIL.n42 30.052
R191 VTAIL.n87 VTAIL.n86 30.052
R192 VTAIL.n131 VTAIL.n130 30.052
R193 VTAIL.n307 VTAIL.n306 30.052
R194 VTAIL.n263 VTAIL.n262 30.052
R195 VTAIL.n219 VTAIL.n218 30.052
R196 VTAIL.n175 VTAIL.n174 30.052
R197 VTAIL.n351 VTAIL.n307 19.8755
R198 VTAIL.n175 VTAIL.n131 19.8755
R199 VTAIL.n323 VTAIL.n321 16.3894
R200 VTAIL.n15 VTAIL.n13 16.3894
R201 VTAIL.n59 VTAIL.n57 16.3894
R202 VTAIL.n103 VTAIL.n101 16.3894
R203 VTAIL.n279 VTAIL.n277 16.3894
R204 VTAIL.n235 VTAIL.n233 16.3894
R205 VTAIL.n191 VTAIL.n189 16.3894
R206 VTAIL.n147 VTAIL.n145 16.3894
R207 VTAIL.n324 VTAIL.n320 12.8005
R208 VTAIL.n16 VTAIL.n12 12.8005
R209 VTAIL.n60 VTAIL.n56 12.8005
R210 VTAIL.n104 VTAIL.n100 12.8005
R211 VTAIL.n280 VTAIL.n276 12.8005
R212 VTAIL.n236 VTAIL.n232 12.8005
R213 VTAIL.n192 VTAIL.n188 12.8005
R214 VTAIL.n148 VTAIL.n144 12.8005
R215 VTAIL.n328 VTAIL.n327 12.0247
R216 VTAIL.n20 VTAIL.n19 12.0247
R217 VTAIL.n64 VTAIL.n63 12.0247
R218 VTAIL.n108 VTAIL.n107 12.0247
R219 VTAIL.n284 VTAIL.n283 12.0247
R220 VTAIL.n240 VTAIL.n239 12.0247
R221 VTAIL.n196 VTAIL.n195 12.0247
R222 VTAIL.n152 VTAIL.n151 12.0247
R223 VTAIL.n331 VTAIL.n318 11.249
R224 VTAIL.n23 VTAIL.n10 11.249
R225 VTAIL.n67 VTAIL.n54 11.249
R226 VTAIL.n111 VTAIL.n98 11.249
R227 VTAIL.n287 VTAIL.n274 11.249
R228 VTAIL.n243 VTAIL.n230 11.249
R229 VTAIL.n199 VTAIL.n186 11.249
R230 VTAIL.n155 VTAIL.n142 11.249
R231 VTAIL.n332 VTAIL.n316 10.4732
R232 VTAIL.n24 VTAIL.n8 10.4732
R233 VTAIL.n68 VTAIL.n52 10.4732
R234 VTAIL.n112 VTAIL.n96 10.4732
R235 VTAIL.n288 VTAIL.n272 10.4732
R236 VTAIL.n244 VTAIL.n228 10.4732
R237 VTAIL.n200 VTAIL.n184 10.4732
R238 VTAIL.n156 VTAIL.n140 10.4732
R239 VTAIL.n336 VTAIL.n335 9.69747
R240 VTAIL.n28 VTAIL.n27 9.69747
R241 VTAIL.n72 VTAIL.n71 9.69747
R242 VTAIL.n116 VTAIL.n115 9.69747
R243 VTAIL.n292 VTAIL.n291 9.69747
R244 VTAIL.n248 VTAIL.n247 9.69747
R245 VTAIL.n204 VTAIL.n203 9.69747
R246 VTAIL.n160 VTAIL.n159 9.69747
R247 VTAIL.n350 VTAIL.n349 9.45567
R248 VTAIL.n42 VTAIL.n41 9.45567
R249 VTAIL.n86 VTAIL.n85 9.45567
R250 VTAIL.n130 VTAIL.n129 9.45567
R251 VTAIL.n306 VTAIL.n305 9.45567
R252 VTAIL.n262 VTAIL.n261 9.45567
R253 VTAIL.n218 VTAIL.n217 9.45567
R254 VTAIL.n174 VTAIL.n173 9.45567
R255 VTAIL.n310 VTAIL.n309 9.3005
R256 VTAIL.n349 VTAIL.n348 9.3005
R257 VTAIL.n341 VTAIL.n340 9.3005
R258 VTAIL.n314 VTAIL.n313 9.3005
R259 VTAIL.n335 VTAIL.n334 9.3005
R260 VTAIL.n333 VTAIL.n332 9.3005
R261 VTAIL.n318 VTAIL.n317 9.3005
R262 VTAIL.n327 VTAIL.n326 9.3005
R263 VTAIL.n325 VTAIL.n324 9.3005
R264 VTAIL.n343 VTAIL.n342 9.3005
R265 VTAIL.n2 VTAIL.n1 9.3005
R266 VTAIL.n41 VTAIL.n40 9.3005
R267 VTAIL.n33 VTAIL.n32 9.3005
R268 VTAIL.n6 VTAIL.n5 9.3005
R269 VTAIL.n27 VTAIL.n26 9.3005
R270 VTAIL.n25 VTAIL.n24 9.3005
R271 VTAIL.n10 VTAIL.n9 9.3005
R272 VTAIL.n19 VTAIL.n18 9.3005
R273 VTAIL.n17 VTAIL.n16 9.3005
R274 VTAIL.n35 VTAIL.n34 9.3005
R275 VTAIL.n46 VTAIL.n45 9.3005
R276 VTAIL.n85 VTAIL.n84 9.3005
R277 VTAIL.n77 VTAIL.n76 9.3005
R278 VTAIL.n50 VTAIL.n49 9.3005
R279 VTAIL.n71 VTAIL.n70 9.3005
R280 VTAIL.n69 VTAIL.n68 9.3005
R281 VTAIL.n54 VTAIL.n53 9.3005
R282 VTAIL.n63 VTAIL.n62 9.3005
R283 VTAIL.n61 VTAIL.n60 9.3005
R284 VTAIL.n79 VTAIL.n78 9.3005
R285 VTAIL.n90 VTAIL.n89 9.3005
R286 VTAIL.n129 VTAIL.n128 9.3005
R287 VTAIL.n121 VTAIL.n120 9.3005
R288 VTAIL.n94 VTAIL.n93 9.3005
R289 VTAIL.n115 VTAIL.n114 9.3005
R290 VTAIL.n113 VTAIL.n112 9.3005
R291 VTAIL.n98 VTAIL.n97 9.3005
R292 VTAIL.n107 VTAIL.n106 9.3005
R293 VTAIL.n105 VTAIL.n104 9.3005
R294 VTAIL.n123 VTAIL.n122 9.3005
R295 VTAIL.n266 VTAIL.n265 9.3005
R296 VTAIL.n299 VTAIL.n298 9.3005
R297 VTAIL.n297 VTAIL.n296 9.3005
R298 VTAIL.n270 VTAIL.n269 9.3005
R299 VTAIL.n291 VTAIL.n290 9.3005
R300 VTAIL.n289 VTAIL.n288 9.3005
R301 VTAIL.n274 VTAIL.n273 9.3005
R302 VTAIL.n283 VTAIL.n282 9.3005
R303 VTAIL.n281 VTAIL.n280 9.3005
R304 VTAIL.n305 VTAIL.n304 9.3005
R305 VTAIL.n261 VTAIL.n260 9.3005
R306 VTAIL.n222 VTAIL.n221 9.3005
R307 VTAIL.n255 VTAIL.n254 9.3005
R308 VTAIL.n253 VTAIL.n252 9.3005
R309 VTAIL.n226 VTAIL.n225 9.3005
R310 VTAIL.n247 VTAIL.n246 9.3005
R311 VTAIL.n245 VTAIL.n244 9.3005
R312 VTAIL.n230 VTAIL.n229 9.3005
R313 VTAIL.n239 VTAIL.n238 9.3005
R314 VTAIL.n237 VTAIL.n236 9.3005
R315 VTAIL.n217 VTAIL.n216 9.3005
R316 VTAIL.n178 VTAIL.n177 9.3005
R317 VTAIL.n211 VTAIL.n210 9.3005
R318 VTAIL.n209 VTAIL.n208 9.3005
R319 VTAIL.n182 VTAIL.n181 9.3005
R320 VTAIL.n203 VTAIL.n202 9.3005
R321 VTAIL.n201 VTAIL.n200 9.3005
R322 VTAIL.n186 VTAIL.n185 9.3005
R323 VTAIL.n195 VTAIL.n194 9.3005
R324 VTAIL.n193 VTAIL.n192 9.3005
R325 VTAIL.n173 VTAIL.n172 9.3005
R326 VTAIL.n134 VTAIL.n133 9.3005
R327 VTAIL.n167 VTAIL.n166 9.3005
R328 VTAIL.n165 VTAIL.n164 9.3005
R329 VTAIL.n138 VTAIL.n137 9.3005
R330 VTAIL.n159 VTAIL.n158 9.3005
R331 VTAIL.n157 VTAIL.n156 9.3005
R332 VTAIL.n142 VTAIL.n141 9.3005
R333 VTAIL.n151 VTAIL.n150 9.3005
R334 VTAIL.n149 VTAIL.n148 9.3005
R335 VTAIL.n339 VTAIL.n314 8.92171
R336 VTAIL.n31 VTAIL.n6 8.92171
R337 VTAIL.n75 VTAIL.n50 8.92171
R338 VTAIL.n119 VTAIL.n94 8.92171
R339 VTAIL.n295 VTAIL.n270 8.92171
R340 VTAIL.n251 VTAIL.n226 8.92171
R341 VTAIL.n207 VTAIL.n182 8.92171
R342 VTAIL.n163 VTAIL.n138 8.92171
R343 VTAIL.n340 VTAIL.n312 8.14595
R344 VTAIL.n350 VTAIL.n308 8.14595
R345 VTAIL.n32 VTAIL.n4 8.14595
R346 VTAIL.n42 VTAIL.n0 8.14595
R347 VTAIL.n76 VTAIL.n48 8.14595
R348 VTAIL.n86 VTAIL.n44 8.14595
R349 VTAIL.n120 VTAIL.n92 8.14595
R350 VTAIL.n130 VTAIL.n88 8.14595
R351 VTAIL.n306 VTAIL.n264 8.14595
R352 VTAIL.n296 VTAIL.n268 8.14595
R353 VTAIL.n262 VTAIL.n220 8.14595
R354 VTAIL.n252 VTAIL.n224 8.14595
R355 VTAIL.n218 VTAIL.n176 8.14595
R356 VTAIL.n208 VTAIL.n180 8.14595
R357 VTAIL.n174 VTAIL.n132 8.14595
R358 VTAIL.n164 VTAIL.n136 8.14595
R359 VTAIL.n344 VTAIL.n343 7.3702
R360 VTAIL.n348 VTAIL.n347 7.3702
R361 VTAIL.n36 VTAIL.n35 7.3702
R362 VTAIL.n40 VTAIL.n39 7.3702
R363 VTAIL.n80 VTAIL.n79 7.3702
R364 VTAIL.n84 VTAIL.n83 7.3702
R365 VTAIL.n124 VTAIL.n123 7.3702
R366 VTAIL.n128 VTAIL.n127 7.3702
R367 VTAIL.n304 VTAIL.n303 7.3702
R368 VTAIL.n300 VTAIL.n299 7.3702
R369 VTAIL.n260 VTAIL.n259 7.3702
R370 VTAIL.n256 VTAIL.n255 7.3702
R371 VTAIL.n216 VTAIL.n215 7.3702
R372 VTAIL.n212 VTAIL.n211 7.3702
R373 VTAIL.n172 VTAIL.n171 7.3702
R374 VTAIL.n168 VTAIL.n167 7.3702
R375 VTAIL.n344 VTAIL.n310 6.59444
R376 VTAIL.n347 VTAIL.n310 6.59444
R377 VTAIL.n36 VTAIL.n2 6.59444
R378 VTAIL.n39 VTAIL.n2 6.59444
R379 VTAIL.n80 VTAIL.n46 6.59444
R380 VTAIL.n83 VTAIL.n46 6.59444
R381 VTAIL.n124 VTAIL.n90 6.59444
R382 VTAIL.n127 VTAIL.n90 6.59444
R383 VTAIL.n303 VTAIL.n266 6.59444
R384 VTAIL.n300 VTAIL.n266 6.59444
R385 VTAIL.n259 VTAIL.n222 6.59444
R386 VTAIL.n256 VTAIL.n222 6.59444
R387 VTAIL.n215 VTAIL.n178 6.59444
R388 VTAIL.n212 VTAIL.n178 6.59444
R389 VTAIL.n171 VTAIL.n134 6.59444
R390 VTAIL.n168 VTAIL.n134 6.59444
R391 VTAIL.n343 VTAIL.n312 5.81868
R392 VTAIL.n348 VTAIL.n308 5.81868
R393 VTAIL.n35 VTAIL.n4 5.81868
R394 VTAIL.n40 VTAIL.n0 5.81868
R395 VTAIL.n79 VTAIL.n48 5.81868
R396 VTAIL.n84 VTAIL.n44 5.81868
R397 VTAIL.n123 VTAIL.n92 5.81868
R398 VTAIL.n128 VTAIL.n88 5.81868
R399 VTAIL.n304 VTAIL.n264 5.81868
R400 VTAIL.n299 VTAIL.n268 5.81868
R401 VTAIL.n260 VTAIL.n220 5.81868
R402 VTAIL.n255 VTAIL.n224 5.81868
R403 VTAIL.n216 VTAIL.n176 5.81868
R404 VTAIL.n211 VTAIL.n180 5.81868
R405 VTAIL.n172 VTAIL.n132 5.81868
R406 VTAIL.n167 VTAIL.n136 5.81868
R407 VTAIL.n340 VTAIL.n339 5.04292
R408 VTAIL.n32 VTAIL.n31 5.04292
R409 VTAIL.n76 VTAIL.n75 5.04292
R410 VTAIL.n120 VTAIL.n119 5.04292
R411 VTAIL.n296 VTAIL.n295 5.04292
R412 VTAIL.n252 VTAIL.n251 5.04292
R413 VTAIL.n208 VTAIL.n207 5.04292
R414 VTAIL.n164 VTAIL.n163 5.04292
R415 VTAIL.n336 VTAIL.n314 4.26717
R416 VTAIL.n28 VTAIL.n6 4.26717
R417 VTAIL.n72 VTAIL.n50 4.26717
R418 VTAIL.n116 VTAIL.n94 4.26717
R419 VTAIL.n292 VTAIL.n270 4.26717
R420 VTAIL.n248 VTAIL.n226 4.26717
R421 VTAIL.n204 VTAIL.n182 4.26717
R422 VTAIL.n160 VTAIL.n138 4.26717
R423 VTAIL.n325 VTAIL.n321 3.70995
R424 VTAIL.n17 VTAIL.n13 3.70995
R425 VTAIL.n61 VTAIL.n57 3.70995
R426 VTAIL.n105 VTAIL.n101 3.70995
R427 VTAIL.n237 VTAIL.n233 3.70995
R428 VTAIL.n193 VTAIL.n189 3.70995
R429 VTAIL.n149 VTAIL.n145 3.70995
R430 VTAIL.n281 VTAIL.n277 3.70995
R431 VTAIL.n335 VTAIL.n316 3.49141
R432 VTAIL.n27 VTAIL.n8 3.49141
R433 VTAIL.n71 VTAIL.n52 3.49141
R434 VTAIL.n115 VTAIL.n96 3.49141
R435 VTAIL.n291 VTAIL.n272 3.49141
R436 VTAIL.n247 VTAIL.n228 3.49141
R437 VTAIL.n203 VTAIL.n184 3.49141
R438 VTAIL.n159 VTAIL.n140 3.49141
R439 VTAIL.n332 VTAIL.n331 2.71565
R440 VTAIL.n24 VTAIL.n23 2.71565
R441 VTAIL.n68 VTAIL.n67 2.71565
R442 VTAIL.n112 VTAIL.n111 2.71565
R443 VTAIL.n288 VTAIL.n287 2.71565
R444 VTAIL.n244 VTAIL.n243 2.71565
R445 VTAIL.n200 VTAIL.n199 2.71565
R446 VTAIL.n156 VTAIL.n155 2.71565
R447 VTAIL.n328 VTAIL.n318 1.93989
R448 VTAIL.n20 VTAIL.n10 1.93989
R449 VTAIL.n64 VTAIL.n54 1.93989
R450 VTAIL.n108 VTAIL.n98 1.93989
R451 VTAIL.n284 VTAIL.n274 1.93989
R452 VTAIL.n240 VTAIL.n230 1.93989
R453 VTAIL.n196 VTAIL.n186 1.93989
R454 VTAIL.n152 VTAIL.n142 1.93989
R455 VTAIL.n327 VTAIL.n320 1.16414
R456 VTAIL.n19 VTAIL.n12 1.16414
R457 VTAIL.n63 VTAIL.n56 1.16414
R458 VTAIL.n107 VTAIL.n100 1.16414
R459 VTAIL.n283 VTAIL.n276 1.16414
R460 VTAIL.n239 VTAIL.n232 1.16414
R461 VTAIL.n195 VTAIL.n188 1.16414
R462 VTAIL.n151 VTAIL.n144 1.16414
R463 VTAIL.n219 VTAIL.n175 0.552224
R464 VTAIL.n307 VTAIL.n263 0.552224
R465 VTAIL.n131 VTAIL.n87 0.552224
R466 VTAIL.n263 VTAIL.n219 0.470328
R467 VTAIL.n87 VTAIL.n43 0.470328
R468 VTAIL.n324 VTAIL.n323 0.388379
R469 VTAIL.n16 VTAIL.n15 0.388379
R470 VTAIL.n60 VTAIL.n59 0.388379
R471 VTAIL.n104 VTAIL.n103 0.388379
R472 VTAIL.n280 VTAIL.n279 0.388379
R473 VTAIL.n236 VTAIL.n235 0.388379
R474 VTAIL.n192 VTAIL.n191 0.388379
R475 VTAIL.n148 VTAIL.n147 0.388379
R476 VTAIL VTAIL.n43 0.334552
R477 VTAIL VTAIL.n351 0.218172
R478 VTAIL.n326 VTAIL.n325 0.155672
R479 VTAIL.n326 VTAIL.n317 0.155672
R480 VTAIL.n333 VTAIL.n317 0.155672
R481 VTAIL.n334 VTAIL.n333 0.155672
R482 VTAIL.n334 VTAIL.n313 0.155672
R483 VTAIL.n341 VTAIL.n313 0.155672
R484 VTAIL.n342 VTAIL.n341 0.155672
R485 VTAIL.n342 VTAIL.n309 0.155672
R486 VTAIL.n349 VTAIL.n309 0.155672
R487 VTAIL.n18 VTAIL.n17 0.155672
R488 VTAIL.n18 VTAIL.n9 0.155672
R489 VTAIL.n25 VTAIL.n9 0.155672
R490 VTAIL.n26 VTAIL.n25 0.155672
R491 VTAIL.n26 VTAIL.n5 0.155672
R492 VTAIL.n33 VTAIL.n5 0.155672
R493 VTAIL.n34 VTAIL.n33 0.155672
R494 VTAIL.n34 VTAIL.n1 0.155672
R495 VTAIL.n41 VTAIL.n1 0.155672
R496 VTAIL.n62 VTAIL.n61 0.155672
R497 VTAIL.n62 VTAIL.n53 0.155672
R498 VTAIL.n69 VTAIL.n53 0.155672
R499 VTAIL.n70 VTAIL.n69 0.155672
R500 VTAIL.n70 VTAIL.n49 0.155672
R501 VTAIL.n77 VTAIL.n49 0.155672
R502 VTAIL.n78 VTAIL.n77 0.155672
R503 VTAIL.n78 VTAIL.n45 0.155672
R504 VTAIL.n85 VTAIL.n45 0.155672
R505 VTAIL.n106 VTAIL.n105 0.155672
R506 VTAIL.n106 VTAIL.n97 0.155672
R507 VTAIL.n113 VTAIL.n97 0.155672
R508 VTAIL.n114 VTAIL.n113 0.155672
R509 VTAIL.n114 VTAIL.n93 0.155672
R510 VTAIL.n121 VTAIL.n93 0.155672
R511 VTAIL.n122 VTAIL.n121 0.155672
R512 VTAIL.n122 VTAIL.n89 0.155672
R513 VTAIL.n129 VTAIL.n89 0.155672
R514 VTAIL.n305 VTAIL.n265 0.155672
R515 VTAIL.n298 VTAIL.n265 0.155672
R516 VTAIL.n298 VTAIL.n297 0.155672
R517 VTAIL.n297 VTAIL.n269 0.155672
R518 VTAIL.n290 VTAIL.n269 0.155672
R519 VTAIL.n290 VTAIL.n289 0.155672
R520 VTAIL.n289 VTAIL.n273 0.155672
R521 VTAIL.n282 VTAIL.n273 0.155672
R522 VTAIL.n282 VTAIL.n281 0.155672
R523 VTAIL.n261 VTAIL.n221 0.155672
R524 VTAIL.n254 VTAIL.n221 0.155672
R525 VTAIL.n254 VTAIL.n253 0.155672
R526 VTAIL.n253 VTAIL.n225 0.155672
R527 VTAIL.n246 VTAIL.n225 0.155672
R528 VTAIL.n246 VTAIL.n245 0.155672
R529 VTAIL.n245 VTAIL.n229 0.155672
R530 VTAIL.n238 VTAIL.n229 0.155672
R531 VTAIL.n238 VTAIL.n237 0.155672
R532 VTAIL.n217 VTAIL.n177 0.155672
R533 VTAIL.n210 VTAIL.n177 0.155672
R534 VTAIL.n210 VTAIL.n209 0.155672
R535 VTAIL.n209 VTAIL.n181 0.155672
R536 VTAIL.n202 VTAIL.n181 0.155672
R537 VTAIL.n202 VTAIL.n201 0.155672
R538 VTAIL.n201 VTAIL.n185 0.155672
R539 VTAIL.n194 VTAIL.n185 0.155672
R540 VTAIL.n194 VTAIL.n193 0.155672
R541 VTAIL.n173 VTAIL.n133 0.155672
R542 VTAIL.n166 VTAIL.n133 0.155672
R543 VTAIL.n166 VTAIL.n165 0.155672
R544 VTAIL.n165 VTAIL.n137 0.155672
R545 VTAIL.n158 VTAIL.n137 0.155672
R546 VTAIL.n158 VTAIL.n157 0.155672
R547 VTAIL.n157 VTAIL.n141 0.155672
R548 VTAIL.n150 VTAIL.n141 0.155672
R549 VTAIL.n150 VTAIL.n149 0.155672
R550 B.n83 B.t6 840.794
R551 B.n183 B.t3 840.794
R552 B.n32 B.t9 840.794
R553 B.n24 B.t0 840.794
R554 B.n232 B.n231 585
R555 B.n230 B.n63 585
R556 B.n229 B.n228 585
R557 B.n227 B.n64 585
R558 B.n226 B.n225 585
R559 B.n224 B.n65 585
R560 B.n223 B.n222 585
R561 B.n221 B.n66 585
R562 B.n220 B.n219 585
R563 B.n218 B.n67 585
R564 B.n217 B.n216 585
R565 B.n215 B.n68 585
R566 B.n214 B.n213 585
R567 B.n212 B.n69 585
R568 B.n211 B.n210 585
R569 B.n209 B.n70 585
R570 B.n208 B.n207 585
R571 B.n206 B.n71 585
R572 B.n205 B.n204 585
R573 B.n203 B.n72 585
R574 B.n202 B.n201 585
R575 B.n200 B.n73 585
R576 B.n199 B.n198 585
R577 B.n197 B.n74 585
R578 B.n196 B.n195 585
R579 B.n194 B.n75 585
R580 B.n193 B.n192 585
R581 B.n191 B.n76 585
R582 B.n190 B.n189 585
R583 B.n188 B.n77 585
R584 B.n187 B.n186 585
R585 B.n182 B.n78 585
R586 B.n181 B.n180 585
R587 B.n179 B.n79 585
R588 B.n178 B.n177 585
R589 B.n176 B.n80 585
R590 B.n175 B.n174 585
R591 B.n173 B.n81 585
R592 B.n172 B.n171 585
R593 B.n170 B.n82 585
R594 B.n168 B.n167 585
R595 B.n166 B.n85 585
R596 B.n165 B.n164 585
R597 B.n163 B.n86 585
R598 B.n162 B.n161 585
R599 B.n160 B.n87 585
R600 B.n159 B.n158 585
R601 B.n157 B.n88 585
R602 B.n156 B.n155 585
R603 B.n154 B.n89 585
R604 B.n153 B.n152 585
R605 B.n151 B.n90 585
R606 B.n150 B.n149 585
R607 B.n148 B.n91 585
R608 B.n147 B.n146 585
R609 B.n145 B.n92 585
R610 B.n144 B.n143 585
R611 B.n142 B.n93 585
R612 B.n141 B.n140 585
R613 B.n139 B.n94 585
R614 B.n138 B.n137 585
R615 B.n136 B.n95 585
R616 B.n135 B.n134 585
R617 B.n133 B.n96 585
R618 B.n132 B.n131 585
R619 B.n130 B.n97 585
R620 B.n129 B.n128 585
R621 B.n127 B.n98 585
R622 B.n126 B.n125 585
R623 B.n124 B.n99 585
R624 B.n233 B.n62 585
R625 B.n235 B.n234 585
R626 B.n236 B.n61 585
R627 B.n238 B.n237 585
R628 B.n239 B.n60 585
R629 B.n241 B.n240 585
R630 B.n242 B.n59 585
R631 B.n244 B.n243 585
R632 B.n245 B.n58 585
R633 B.n247 B.n246 585
R634 B.n248 B.n57 585
R635 B.n250 B.n249 585
R636 B.n251 B.n56 585
R637 B.n253 B.n252 585
R638 B.n254 B.n55 585
R639 B.n256 B.n255 585
R640 B.n257 B.n54 585
R641 B.n259 B.n258 585
R642 B.n260 B.n53 585
R643 B.n262 B.n261 585
R644 B.n263 B.n52 585
R645 B.n265 B.n264 585
R646 B.n266 B.n51 585
R647 B.n268 B.n267 585
R648 B.n269 B.n50 585
R649 B.n271 B.n270 585
R650 B.n272 B.n49 585
R651 B.n274 B.n273 585
R652 B.n380 B.n379 585
R653 B.n378 B.n9 585
R654 B.n377 B.n376 585
R655 B.n375 B.n10 585
R656 B.n374 B.n373 585
R657 B.n372 B.n11 585
R658 B.n371 B.n370 585
R659 B.n369 B.n12 585
R660 B.n368 B.n367 585
R661 B.n366 B.n13 585
R662 B.n365 B.n364 585
R663 B.n363 B.n14 585
R664 B.n362 B.n361 585
R665 B.n360 B.n15 585
R666 B.n359 B.n358 585
R667 B.n357 B.n16 585
R668 B.n356 B.n355 585
R669 B.n354 B.n17 585
R670 B.n353 B.n352 585
R671 B.n351 B.n18 585
R672 B.n350 B.n349 585
R673 B.n348 B.n19 585
R674 B.n347 B.n346 585
R675 B.n345 B.n20 585
R676 B.n344 B.n343 585
R677 B.n342 B.n21 585
R678 B.n341 B.n340 585
R679 B.n339 B.n22 585
R680 B.n338 B.n337 585
R681 B.n336 B.n23 585
R682 B.n334 B.n333 585
R683 B.n332 B.n26 585
R684 B.n331 B.n330 585
R685 B.n329 B.n27 585
R686 B.n328 B.n327 585
R687 B.n326 B.n28 585
R688 B.n325 B.n324 585
R689 B.n323 B.n29 585
R690 B.n322 B.n321 585
R691 B.n320 B.n30 585
R692 B.n319 B.n318 585
R693 B.n317 B.n31 585
R694 B.n316 B.n315 585
R695 B.n314 B.n35 585
R696 B.n313 B.n312 585
R697 B.n311 B.n36 585
R698 B.n310 B.n309 585
R699 B.n308 B.n37 585
R700 B.n307 B.n306 585
R701 B.n305 B.n38 585
R702 B.n304 B.n303 585
R703 B.n302 B.n39 585
R704 B.n301 B.n300 585
R705 B.n299 B.n40 585
R706 B.n298 B.n297 585
R707 B.n296 B.n41 585
R708 B.n295 B.n294 585
R709 B.n293 B.n42 585
R710 B.n292 B.n291 585
R711 B.n290 B.n43 585
R712 B.n289 B.n288 585
R713 B.n287 B.n44 585
R714 B.n286 B.n285 585
R715 B.n284 B.n45 585
R716 B.n283 B.n282 585
R717 B.n281 B.n46 585
R718 B.n280 B.n279 585
R719 B.n278 B.n47 585
R720 B.n277 B.n276 585
R721 B.n275 B.n48 585
R722 B.n381 B.n8 585
R723 B.n383 B.n382 585
R724 B.n384 B.n7 585
R725 B.n386 B.n385 585
R726 B.n387 B.n6 585
R727 B.n389 B.n388 585
R728 B.n390 B.n5 585
R729 B.n392 B.n391 585
R730 B.n393 B.n4 585
R731 B.n395 B.n394 585
R732 B.n396 B.n3 585
R733 B.n398 B.n397 585
R734 B.n399 B.n0 585
R735 B.n2 B.n1 585
R736 B.n106 B.n105 585
R737 B.n108 B.n107 585
R738 B.n109 B.n104 585
R739 B.n111 B.n110 585
R740 B.n112 B.n103 585
R741 B.n114 B.n113 585
R742 B.n115 B.n102 585
R743 B.n117 B.n116 585
R744 B.n118 B.n101 585
R745 B.n120 B.n119 585
R746 B.n121 B.n100 585
R747 B.n123 B.n122 585
R748 B.n124 B.n123 516.524
R749 B.n231 B.n62 516.524
R750 B.n273 B.n48 516.524
R751 B.n381 B.n380 516.524
R752 B.n183 B.t4 317.072
R753 B.n32 B.t11 317.072
R754 B.n83 B.t7 317.072
R755 B.n24 B.t2 317.072
R756 B.n184 B.t5 304.659
R757 B.n33 B.t10 304.659
R758 B.n84 B.t8 304.659
R759 B.n25 B.t1 304.659
R760 B.n401 B.n400 256.663
R761 B.n400 B.n399 235.042
R762 B.n400 B.n2 235.042
R763 B.n125 B.n124 163.367
R764 B.n125 B.n98 163.367
R765 B.n129 B.n98 163.367
R766 B.n130 B.n129 163.367
R767 B.n131 B.n130 163.367
R768 B.n131 B.n96 163.367
R769 B.n135 B.n96 163.367
R770 B.n136 B.n135 163.367
R771 B.n137 B.n136 163.367
R772 B.n137 B.n94 163.367
R773 B.n141 B.n94 163.367
R774 B.n142 B.n141 163.367
R775 B.n143 B.n142 163.367
R776 B.n143 B.n92 163.367
R777 B.n147 B.n92 163.367
R778 B.n148 B.n147 163.367
R779 B.n149 B.n148 163.367
R780 B.n149 B.n90 163.367
R781 B.n153 B.n90 163.367
R782 B.n154 B.n153 163.367
R783 B.n155 B.n154 163.367
R784 B.n155 B.n88 163.367
R785 B.n159 B.n88 163.367
R786 B.n160 B.n159 163.367
R787 B.n161 B.n160 163.367
R788 B.n161 B.n86 163.367
R789 B.n165 B.n86 163.367
R790 B.n166 B.n165 163.367
R791 B.n167 B.n166 163.367
R792 B.n167 B.n82 163.367
R793 B.n172 B.n82 163.367
R794 B.n173 B.n172 163.367
R795 B.n174 B.n173 163.367
R796 B.n174 B.n80 163.367
R797 B.n178 B.n80 163.367
R798 B.n179 B.n178 163.367
R799 B.n180 B.n179 163.367
R800 B.n180 B.n78 163.367
R801 B.n187 B.n78 163.367
R802 B.n188 B.n187 163.367
R803 B.n189 B.n188 163.367
R804 B.n189 B.n76 163.367
R805 B.n193 B.n76 163.367
R806 B.n194 B.n193 163.367
R807 B.n195 B.n194 163.367
R808 B.n195 B.n74 163.367
R809 B.n199 B.n74 163.367
R810 B.n200 B.n199 163.367
R811 B.n201 B.n200 163.367
R812 B.n201 B.n72 163.367
R813 B.n205 B.n72 163.367
R814 B.n206 B.n205 163.367
R815 B.n207 B.n206 163.367
R816 B.n207 B.n70 163.367
R817 B.n211 B.n70 163.367
R818 B.n212 B.n211 163.367
R819 B.n213 B.n212 163.367
R820 B.n213 B.n68 163.367
R821 B.n217 B.n68 163.367
R822 B.n218 B.n217 163.367
R823 B.n219 B.n218 163.367
R824 B.n219 B.n66 163.367
R825 B.n223 B.n66 163.367
R826 B.n224 B.n223 163.367
R827 B.n225 B.n224 163.367
R828 B.n225 B.n64 163.367
R829 B.n229 B.n64 163.367
R830 B.n230 B.n229 163.367
R831 B.n231 B.n230 163.367
R832 B.n273 B.n272 163.367
R833 B.n272 B.n271 163.367
R834 B.n271 B.n50 163.367
R835 B.n267 B.n50 163.367
R836 B.n267 B.n266 163.367
R837 B.n266 B.n265 163.367
R838 B.n265 B.n52 163.367
R839 B.n261 B.n52 163.367
R840 B.n261 B.n260 163.367
R841 B.n260 B.n259 163.367
R842 B.n259 B.n54 163.367
R843 B.n255 B.n54 163.367
R844 B.n255 B.n254 163.367
R845 B.n254 B.n253 163.367
R846 B.n253 B.n56 163.367
R847 B.n249 B.n56 163.367
R848 B.n249 B.n248 163.367
R849 B.n248 B.n247 163.367
R850 B.n247 B.n58 163.367
R851 B.n243 B.n58 163.367
R852 B.n243 B.n242 163.367
R853 B.n242 B.n241 163.367
R854 B.n241 B.n60 163.367
R855 B.n237 B.n60 163.367
R856 B.n237 B.n236 163.367
R857 B.n236 B.n235 163.367
R858 B.n235 B.n62 163.367
R859 B.n380 B.n9 163.367
R860 B.n376 B.n9 163.367
R861 B.n376 B.n375 163.367
R862 B.n375 B.n374 163.367
R863 B.n374 B.n11 163.367
R864 B.n370 B.n11 163.367
R865 B.n370 B.n369 163.367
R866 B.n369 B.n368 163.367
R867 B.n368 B.n13 163.367
R868 B.n364 B.n13 163.367
R869 B.n364 B.n363 163.367
R870 B.n363 B.n362 163.367
R871 B.n362 B.n15 163.367
R872 B.n358 B.n15 163.367
R873 B.n358 B.n357 163.367
R874 B.n357 B.n356 163.367
R875 B.n356 B.n17 163.367
R876 B.n352 B.n17 163.367
R877 B.n352 B.n351 163.367
R878 B.n351 B.n350 163.367
R879 B.n350 B.n19 163.367
R880 B.n346 B.n19 163.367
R881 B.n346 B.n345 163.367
R882 B.n345 B.n344 163.367
R883 B.n344 B.n21 163.367
R884 B.n340 B.n21 163.367
R885 B.n340 B.n339 163.367
R886 B.n339 B.n338 163.367
R887 B.n338 B.n23 163.367
R888 B.n333 B.n23 163.367
R889 B.n333 B.n332 163.367
R890 B.n332 B.n331 163.367
R891 B.n331 B.n27 163.367
R892 B.n327 B.n27 163.367
R893 B.n327 B.n326 163.367
R894 B.n326 B.n325 163.367
R895 B.n325 B.n29 163.367
R896 B.n321 B.n29 163.367
R897 B.n321 B.n320 163.367
R898 B.n320 B.n319 163.367
R899 B.n319 B.n31 163.367
R900 B.n315 B.n31 163.367
R901 B.n315 B.n314 163.367
R902 B.n314 B.n313 163.367
R903 B.n313 B.n36 163.367
R904 B.n309 B.n36 163.367
R905 B.n309 B.n308 163.367
R906 B.n308 B.n307 163.367
R907 B.n307 B.n38 163.367
R908 B.n303 B.n38 163.367
R909 B.n303 B.n302 163.367
R910 B.n302 B.n301 163.367
R911 B.n301 B.n40 163.367
R912 B.n297 B.n40 163.367
R913 B.n297 B.n296 163.367
R914 B.n296 B.n295 163.367
R915 B.n295 B.n42 163.367
R916 B.n291 B.n42 163.367
R917 B.n291 B.n290 163.367
R918 B.n290 B.n289 163.367
R919 B.n289 B.n44 163.367
R920 B.n285 B.n44 163.367
R921 B.n285 B.n284 163.367
R922 B.n284 B.n283 163.367
R923 B.n283 B.n46 163.367
R924 B.n279 B.n46 163.367
R925 B.n279 B.n278 163.367
R926 B.n278 B.n277 163.367
R927 B.n277 B.n48 163.367
R928 B.n382 B.n381 163.367
R929 B.n382 B.n7 163.367
R930 B.n386 B.n7 163.367
R931 B.n387 B.n386 163.367
R932 B.n388 B.n387 163.367
R933 B.n388 B.n5 163.367
R934 B.n392 B.n5 163.367
R935 B.n393 B.n392 163.367
R936 B.n394 B.n393 163.367
R937 B.n394 B.n3 163.367
R938 B.n398 B.n3 163.367
R939 B.n399 B.n398 163.367
R940 B.n106 B.n2 163.367
R941 B.n107 B.n106 163.367
R942 B.n107 B.n104 163.367
R943 B.n111 B.n104 163.367
R944 B.n112 B.n111 163.367
R945 B.n113 B.n112 163.367
R946 B.n113 B.n102 163.367
R947 B.n117 B.n102 163.367
R948 B.n118 B.n117 163.367
R949 B.n119 B.n118 163.367
R950 B.n119 B.n100 163.367
R951 B.n123 B.n100 163.367
R952 B.n169 B.n84 59.5399
R953 B.n185 B.n184 59.5399
R954 B.n34 B.n33 59.5399
R955 B.n335 B.n25 59.5399
R956 B.n379 B.n8 33.5615
R957 B.n275 B.n274 33.5615
R958 B.n233 B.n232 33.5615
R959 B.n122 B.n99 33.5615
R960 B B.n401 18.0485
R961 B.n84 B.n83 12.4126
R962 B.n184 B.n183 12.4126
R963 B.n33 B.n32 12.4126
R964 B.n25 B.n24 12.4126
R965 B.n383 B.n8 10.6151
R966 B.n384 B.n383 10.6151
R967 B.n385 B.n384 10.6151
R968 B.n385 B.n6 10.6151
R969 B.n389 B.n6 10.6151
R970 B.n390 B.n389 10.6151
R971 B.n391 B.n390 10.6151
R972 B.n391 B.n4 10.6151
R973 B.n395 B.n4 10.6151
R974 B.n396 B.n395 10.6151
R975 B.n397 B.n396 10.6151
R976 B.n397 B.n0 10.6151
R977 B.n379 B.n378 10.6151
R978 B.n378 B.n377 10.6151
R979 B.n377 B.n10 10.6151
R980 B.n373 B.n10 10.6151
R981 B.n373 B.n372 10.6151
R982 B.n372 B.n371 10.6151
R983 B.n371 B.n12 10.6151
R984 B.n367 B.n12 10.6151
R985 B.n367 B.n366 10.6151
R986 B.n366 B.n365 10.6151
R987 B.n365 B.n14 10.6151
R988 B.n361 B.n14 10.6151
R989 B.n361 B.n360 10.6151
R990 B.n360 B.n359 10.6151
R991 B.n359 B.n16 10.6151
R992 B.n355 B.n16 10.6151
R993 B.n355 B.n354 10.6151
R994 B.n354 B.n353 10.6151
R995 B.n353 B.n18 10.6151
R996 B.n349 B.n18 10.6151
R997 B.n349 B.n348 10.6151
R998 B.n348 B.n347 10.6151
R999 B.n347 B.n20 10.6151
R1000 B.n343 B.n20 10.6151
R1001 B.n343 B.n342 10.6151
R1002 B.n342 B.n341 10.6151
R1003 B.n341 B.n22 10.6151
R1004 B.n337 B.n22 10.6151
R1005 B.n337 B.n336 10.6151
R1006 B.n334 B.n26 10.6151
R1007 B.n330 B.n26 10.6151
R1008 B.n330 B.n329 10.6151
R1009 B.n329 B.n328 10.6151
R1010 B.n328 B.n28 10.6151
R1011 B.n324 B.n28 10.6151
R1012 B.n324 B.n323 10.6151
R1013 B.n323 B.n322 10.6151
R1014 B.n322 B.n30 10.6151
R1015 B.n318 B.n317 10.6151
R1016 B.n317 B.n316 10.6151
R1017 B.n316 B.n35 10.6151
R1018 B.n312 B.n35 10.6151
R1019 B.n312 B.n311 10.6151
R1020 B.n311 B.n310 10.6151
R1021 B.n310 B.n37 10.6151
R1022 B.n306 B.n37 10.6151
R1023 B.n306 B.n305 10.6151
R1024 B.n305 B.n304 10.6151
R1025 B.n304 B.n39 10.6151
R1026 B.n300 B.n39 10.6151
R1027 B.n300 B.n299 10.6151
R1028 B.n299 B.n298 10.6151
R1029 B.n298 B.n41 10.6151
R1030 B.n294 B.n41 10.6151
R1031 B.n294 B.n293 10.6151
R1032 B.n293 B.n292 10.6151
R1033 B.n292 B.n43 10.6151
R1034 B.n288 B.n43 10.6151
R1035 B.n288 B.n287 10.6151
R1036 B.n287 B.n286 10.6151
R1037 B.n286 B.n45 10.6151
R1038 B.n282 B.n45 10.6151
R1039 B.n282 B.n281 10.6151
R1040 B.n281 B.n280 10.6151
R1041 B.n280 B.n47 10.6151
R1042 B.n276 B.n47 10.6151
R1043 B.n276 B.n275 10.6151
R1044 B.n274 B.n49 10.6151
R1045 B.n270 B.n49 10.6151
R1046 B.n270 B.n269 10.6151
R1047 B.n269 B.n268 10.6151
R1048 B.n268 B.n51 10.6151
R1049 B.n264 B.n51 10.6151
R1050 B.n264 B.n263 10.6151
R1051 B.n263 B.n262 10.6151
R1052 B.n262 B.n53 10.6151
R1053 B.n258 B.n53 10.6151
R1054 B.n258 B.n257 10.6151
R1055 B.n257 B.n256 10.6151
R1056 B.n256 B.n55 10.6151
R1057 B.n252 B.n55 10.6151
R1058 B.n252 B.n251 10.6151
R1059 B.n251 B.n250 10.6151
R1060 B.n250 B.n57 10.6151
R1061 B.n246 B.n57 10.6151
R1062 B.n246 B.n245 10.6151
R1063 B.n245 B.n244 10.6151
R1064 B.n244 B.n59 10.6151
R1065 B.n240 B.n59 10.6151
R1066 B.n240 B.n239 10.6151
R1067 B.n239 B.n238 10.6151
R1068 B.n238 B.n61 10.6151
R1069 B.n234 B.n61 10.6151
R1070 B.n234 B.n233 10.6151
R1071 B.n105 B.n1 10.6151
R1072 B.n108 B.n105 10.6151
R1073 B.n109 B.n108 10.6151
R1074 B.n110 B.n109 10.6151
R1075 B.n110 B.n103 10.6151
R1076 B.n114 B.n103 10.6151
R1077 B.n115 B.n114 10.6151
R1078 B.n116 B.n115 10.6151
R1079 B.n116 B.n101 10.6151
R1080 B.n120 B.n101 10.6151
R1081 B.n121 B.n120 10.6151
R1082 B.n122 B.n121 10.6151
R1083 B.n126 B.n99 10.6151
R1084 B.n127 B.n126 10.6151
R1085 B.n128 B.n127 10.6151
R1086 B.n128 B.n97 10.6151
R1087 B.n132 B.n97 10.6151
R1088 B.n133 B.n132 10.6151
R1089 B.n134 B.n133 10.6151
R1090 B.n134 B.n95 10.6151
R1091 B.n138 B.n95 10.6151
R1092 B.n139 B.n138 10.6151
R1093 B.n140 B.n139 10.6151
R1094 B.n140 B.n93 10.6151
R1095 B.n144 B.n93 10.6151
R1096 B.n145 B.n144 10.6151
R1097 B.n146 B.n145 10.6151
R1098 B.n146 B.n91 10.6151
R1099 B.n150 B.n91 10.6151
R1100 B.n151 B.n150 10.6151
R1101 B.n152 B.n151 10.6151
R1102 B.n152 B.n89 10.6151
R1103 B.n156 B.n89 10.6151
R1104 B.n157 B.n156 10.6151
R1105 B.n158 B.n157 10.6151
R1106 B.n158 B.n87 10.6151
R1107 B.n162 B.n87 10.6151
R1108 B.n163 B.n162 10.6151
R1109 B.n164 B.n163 10.6151
R1110 B.n164 B.n85 10.6151
R1111 B.n168 B.n85 10.6151
R1112 B.n171 B.n170 10.6151
R1113 B.n171 B.n81 10.6151
R1114 B.n175 B.n81 10.6151
R1115 B.n176 B.n175 10.6151
R1116 B.n177 B.n176 10.6151
R1117 B.n177 B.n79 10.6151
R1118 B.n181 B.n79 10.6151
R1119 B.n182 B.n181 10.6151
R1120 B.n186 B.n182 10.6151
R1121 B.n190 B.n77 10.6151
R1122 B.n191 B.n190 10.6151
R1123 B.n192 B.n191 10.6151
R1124 B.n192 B.n75 10.6151
R1125 B.n196 B.n75 10.6151
R1126 B.n197 B.n196 10.6151
R1127 B.n198 B.n197 10.6151
R1128 B.n198 B.n73 10.6151
R1129 B.n202 B.n73 10.6151
R1130 B.n203 B.n202 10.6151
R1131 B.n204 B.n203 10.6151
R1132 B.n204 B.n71 10.6151
R1133 B.n208 B.n71 10.6151
R1134 B.n209 B.n208 10.6151
R1135 B.n210 B.n209 10.6151
R1136 B.n210 B.n69 10.6151
R1137 B.n214 B.n69 10.6151
R1138 B.n215 B.n214 10.6151
R1139 B.n216 B.n215 10.6151
R1140 B.n216 B.n67 10.6151
R1141 B.n220 B.n67 10.6151
R1142 B.n221 B.n220 10.6151
R1143 B.n222 B.n221 10.6151
R1144 B.n222 B.n65 10.6151
R1145 B.n226 B.n65 10.6151
R1146 B.n227 B.n226 10.6151
R1147 B.n228 B.n227 10.6151
R1148 B.n228 B.n63 10.6151
R1149 B.n232 B.n63 10.6151
R1150 B.n336 B.n335 8.74196
R1151 B.n318 B.n34 8.74196
R1152 B.n169 B.n168 8.74196
R1153 B.n185 B.n77 8.74196
R1154 B.n401 B.n0 8.11757
R1155 B.n401 B.n1 8.11757
R1156 B.n335 B.n334 1.87367
R1157 B.n34 B.n30 1.87367
R1158 B.n170 B.n169 1.87367
R1159 B.n186 B.n185 1.87367
R1160 VN.n0 VN.t1 774.404
R1161 VN.n0 VN.t2 774.404
R1162 VN.n1 VN.t0 774.404
R1163 VN.n1 VN.t3 774.404
R1164 VN VN.n1 198.014
R1165 VN VN.n0 161.351
R1166 VDD2.n2 VDD2.n0 112.981
R1167 VDD2.n2 VDD2.n1 80.6536
R1168 VDD2.n1 VDD2.t3 4.03839
R1169 VDD2.n1 VDD2.t0 4.03839
R1170 VDD2.n0 VDD2.t1 4.03839
R1171 VDD2.n0 VDD2.t2 4.03839
R1172 VDD2 VDD2.n2 0.0586897
C0 B VDD2 0.766623f
C1 VDD2 w_n1354_n2582# 0.871614f
C2 B VP 0.892054f
C3 VP w_n1354_n2582# 1.96518f
C4 VN VTAIL 1.15919f
C5 VN VDD1 0.14807f
C6 VTAIL VDD1 6.66793f
C7 B w_n1354_n2582# 5.33557f
C8 VN VDD2 1.50648f
C9 VDD2 VTAIL 6.70679f
C10 VDD2 VDD1 0.480601f
C11 VN VP 3.80344f
C12 VP VTAIL 1.1733f
C13 VP VDD1 1.60798f
C14 VN B 0.623475f
C15 VN w_n1354_n2582# 1.79691f
C16 B VTAIL 2.52393f
C17 VP VDD2 0.249729f
C18 VTAIL w_n1354_n2582# 3.20468f
C19 B VDD1 0.750478f
C20 w_n1354_n2582# VDD1 0.86461f
C21 VDD2 VSUBS 0.522196f
C22 VDD1 VSUBS 3.883129f
C23 VTAIL VSUBS 0.597267f
C24 VN VSUBS 3.58283f
C25 VP VSUBS 0.937413f
C26 B VSUBS 1.95409f
C27 w_n1354_n2582# VSUBS 43.3659f
C28 VDD2.t1 VSUBS 0.16716f
C29 VDD2.t2 VSUBS 0.16716f
C30 VDD2.n0 VSUBS 1.61681f
C31 VDD2.t3 VSUBS 0.16716f
C32 VDD2.t0 VSUBS 0.16716f
C33 VDD2.n1 VSUBS 1.18844f
C34 VDD2.n2 VSUBS 3.17374f
C35 VN.t2 VSUBS 0.254653f
C36 VN.t1 VSUBS 0.254653f
C37 VN.n0 VSUBS 0.218642f
C38 VN.t0 VSUBS 0.254653f
C39 VN.t3 VSUBS 0.254653f
C40 VN.n1 VSUBS 0.432435f
C41 B.n0 VSUBS 0.008095f
C42 B.n1 VSUBS 0.008095f
C43 B.n2 VSUBS 0.011973f
C44 B.n3 VSUBS 0.009175f
C45 B.n4 VSUBS 0.009175f
C46 B.n5 VSUBS 0.009175f
C47 B.n6 VSUBS 0.009175f
C48 B.n7 VSUBS 0.009175f
C49 B.n8 VSUBS 0.020995f
C50 B.n9 VSUBS 0.009175f
C51 B.n10 VSUBS 0.009175f
C52 B.n11 VSUBS 0.009175f
C53 B.n12 VSUBS 0.009175f
C54 B.n13 VSUBS 0.009175f
C55 B.n14 VSUBS 0.009175f
C56 B.n15 VSUBS 0.009175f
C57 B.n16 VSUBS 0.009175f
C58 B.n17 VSUBS 0.009175f
C59 B.n18 VSUBS 0.009175f
C60 B.n19 VSUBS 0.009175f
C61 B.n20 VSUBS 0.009175f
C62 B.n21 VSUBS 0.009175f
C63 B.n22 VSUBS 0.009175f
C64 B.n23 VSUBS 0.009175f
C65 B.t1 VSUBS 0.167396f
C66 B.t2 VSUBS 0.176265f
C67 B.t0 VSUBS 0.131114f
C68 B.n24 VSUBS 0.26494f
C69 B.n25 VSUBS 0.239648f
C70 B.n26 VSUBS 0.009175f
C71 B.n27 VSUBS 0.009175f
C72 B.n28 VSUBS 0.009175f
C73 B.n29 VSUBS 0.009175f
C74 B.n30 VSUBS 0.005397f
C75 B.n31 VSUBS 0.009175f
C76 B.t10 VSUBS 0.167399f
C77 B.t11 VSUBS 0.176268f
C78 B.t9 VSUBS 0.131114f
C79 B.n32 VSUBS 0.264937f
C80 B.n33 VSUBS 0.239645f
C81 B.n34 VSUBS 0.021257f
C82 B.n35 VSUBS 0.009175f
C83 B.n36 VSUBS 0.009175f
C84 B.n37 VSUBS 0.009175f
C85 B.n38 VSUBS 0.009175f
C86 B.n39 VSUBS 0.009175f
C87 B.n40 VSUBS 0.009175f
C88 B.n41 VSUBS 0.009175f
C89 B.n42 VSUBS 0.009175f
C90 B.n43 VSUBS 0.009175f
C91 B.n44 VSUBS 0.009175f
C92 B.n45 VSUBS 0.009175f
C93 B.n46 VSUBS 0.009175f
C94 B.n47 VSUBS 0.009175f
C95 B.n48 VSUBS 0.022719f
C96 B.n49 VSUBS 0.009175f
C97 B.n50 VSUBS 0.009175f
C98 B.n51 VSUBS 0.009175f
C99 B.n52 VSUBS 0.009175f
C100 B.n53 VSUBS 0.009175f
C101 B.n54 VSUBS 0.009175f
C102 B.n55 VSUBS 0.009175f
C103 B.n56 VSUBS 0.009175f
C104 B.n57 VSUBS 0.009175f
C105 B.n58 VSUBS 0.009175f
C106 B.n59 VSUBS 0.009175f
C107 B.n60 VSUBS 0.009175f
C108 B.n61 VSUBS 0.009175f
C109 B.n62 VSUBS 0.020995f
C110 B.n63 VSUBS 0.009175f
C111 B.n64 VSUBS 0.009175f
C112 B.n65 VSUBS 0.009175f
C113 B.n66 VSUBS 0.009175f
C114 B.n67 VSUBS 0.009175f
C115 B.n68 VSUBS 0.009175f
C116 B.n69 VSUBS 0.009175f
C117 B.n70 VSUBS 0.009175f
C118 B.n71 VSUBS 0.009175f
C119 B.n72 VSUBS 0.009175f
C120 B.n73 VSUBS 0.009175f
C121 B.n74 VSUBS 0.009175f
C122 B.n75 VSUBS 0.009175f
C123 B.n76 VSUBS 0.009175f
C124 B.n77 VSUBS 0.008365f
C125 B.n78 VSUBS 0.009175f
C126 B.n79 VSUBS 0.009175f
C127 B.n80 VSUBS 0.009175f
C128 B.n81 VSUBS 0.009175f
C129 B.n82 VSUBS 0.009175f
C130 B.t8 VSUBS 0.167396f
C131 B.t7 VSUBS 0.176265f
C132 B.t6 VSUBS 0.131114f
C133 B.n83 VSUBS 0.26494f
C134 B.n84 VSUBS 0.239648f
C135 B.n85 VSUBS 0.009175f
C136 B.n86 VSUBS 0.009175f
C137 B.n87 VSUBS 0.009175f
C138 B.n88 VSUBS 0.009175f
C139 B.n89 VSUBS 0.009175f
C140 B.n90 VSUBS 0.009175f
C141 B.n91 VSUBS 0.009175f
C142 B.n92 VSUBS 0.009175f
C143 B.n93 VSUBS 0.009175f
C144 B.n94 VSUBS 0.009175f
C145 B.n95 VSUBS 0.009175f
C146 B.n96 VSUBS 0.009175f
C147 B.n97 VSUBS 0.009175f
C148 B.n98 VSUBS 0.009175f
C149 B.n99 VSUBS 0.022719f
C150 B.n100 VSUBS 0.009175f
C151 B.n101 VSUBS 0.009175f
C152 B.n102 VSUBS 0.009175f
C153 B.n103 VSUBS 0.009175f
C154 B.n104 VSUBS 0.009175f
C155 B.n105 VSUBS 0.009175f
C156 B.n106 VSUBS 0.009175f
C157 B.n107 VSUBS 0.009175f
C158 B.n108 VSUBS 0.009175f
C159 B.n109 VSUBS 0.009175f
C160 B.n110 VSUBS 0.009175f
C161 B.n111 VSUBS 0.009175f
C162 B.n112 VSUBS 0.009175f
C163 B.n113 VSUBS 0.009175f
C164 B.n114 VSUBS 0.009175f
C165 B.n115 VSUBS 0.009175f
C166 B.n116 VSUBS 0.009175f
C167 B.n117 VSUBS 0.009175f
C168 B.n118 VSUBS 0.009175f
C169 B.n119 VSUBS 0.009175f
C170 B.n120 VSUBS 0.009175f
C171 B.n121 VSUBS 0.009175f
C172 B.n122 VSUBS 0.020995f
C173 B.n123 VSUBS 0.020995f
C174 B.n124 VSUBS 0.022719f
C175 B.n125 VSUBS 0.009175f
C176 B.n126 VSUBS 0.009175f
C177 B.n127 VSUBS 0.009175f
C178 B.n128 VSUBS 0.009175f
C179 B.n129 VSUBS 0.009175f
C180 B.n130 VSUBS 0.009175f
C181 B.n131 VSUBS 0.009175f
C182 B.n132 VSUBS 0.009175f
C183 B.n133 VSUBS 0.009175f
C184 B.n134 VSUBS 0.009175f
C185 B.n135 VSUBS 0.009175f
C186 B.n136 VSUBS 0.009175f
C187 B.n137 VSUBS 0.009175f
C188 B.n138 VSUBS 0.009175f
C189 B.n139 VSUBS 0.009175f
C190 B.n140 VSUBS 0.009175f
C191 B.n141 VSUBS 0.009175f
C192 B.n142 VSUBS 0.009175f
C193 B.n143 VSUBS 0.009175f
C194 B.n144 VSUBS 0.009175f
C195 B.n145 VSUBS 0.009175f
C196 B.n146 VSUBS 0.009175f
C197 B.n147 VSUBS 0.009175f
C198 B.n148 VSUBS 0.009175f
C199 B.n149 VSUBS 0.009175f
C200 B.n150 VSUBS 0.009175f
C201 B.n151 VSUBS 0.009175f
C202 B.n152 VSUBS 0.009175f
C203 B.n153 VSUBS 0.009175f
C204 B.n154 VSUBS 0.009175f
C205 B.n155 VSUBS 0.009175f
C206 B.n156 VSUBS 0.009175f
C207 B.n157 VSUBS 0.009175f
C208 B.n158 VSUBS 0.009175f
C209 B.n159 VSUBS 0.009175f
C210 B.n160 VSUBS 0.009175f
C211 B.n161 VSUBS 0.009175f
C212 B.n162 VSUBS 0.009175f
C213 B.n163 VSUBS 0.009175f
C214 B.n164 VSUBS 0.009175f
C215 B.n165 VSUBS 0.009175f
C216 B.n166 VSUBS 0.009175f
C217 B.n167 VSUBS 0.009175f
C218 B.n168 VSUBS 0.008365f
C219 B.n169 VSUBS 0.021257f
C220 B.n170 VSUBS 0.005397f
C221 B.n171 VSUBS 0.009175f
C222 B.n172 VSUBS 0.009175f
C223 B.n173 VSUBS 0.009175f
C224 B.n174 VSUBS 0.009175f
C225 B.n175 VSUBS 0.009175f
C226 B.n176 VSUBS 0.009175f
C227 B.n177 VSUBS 0.009175f
C228 B.n178 VSUBS 0.009175f
C229 B.n179 VSUBS 0.009175f
C230 B.n180 VSUBS 0.009175f
C231 B.n181 VSUBS 0.009175f
C232 B.n182 VSUBS 0.009175f
C233 B.t5 VSUBS 0.167399f
C234 B.t4 VSUBS 0.176268f
C235 B.t3 VSUBS 0.131114f
C236 B.n183 VSUBS 0.264937f
C237 B.n184 VSUBS 0.239645f
C238 B.n185 VSUBS 0.021257f
C239 B.n186 VSUBS 0.005397f
C240 B.n187 VSUBS 0.009175f
C241 B.n188 VSUBS 0.009175f
C242 B.n189 VSUBS 0.009175f
C243 B.n190 VSUBS 0.009175f
C244 B.n191 VSUBS 0.009175f
C245 B.n192 VSUBS 0.009175f
C246 B.n193 VSUBS 0.009175f
C247 B.n194 VSUBS 0.009175f
C248 B.n195 VSUBS 0.009175f
C249 B.n196 VSUBS 0.009175f
C250 B.n197 VSUBS 0.009175f
C251 B.n198 VSUBS 0.009175f
C252 B.n199 VSUBS 0.009175f
C253 B.n200 VSUBS 0.009175f
C254 B.n201 VSUBS 0.009175f
C255 B.n202 VSUBS 0.009175f
C256 B.n203 VSUBS 0.009175f
C257 B.n204 VSUBS 0.009175f
C258 B.n205 VSUBS 0.009175f
C259 B.n206 VSUBS 0.009175f
C260 B.n207 VSUBS 0.009175f
C261 B.n208 VSUBS 0.009175f
C262 B.n209 VSUBS 0.009175f
C263 B.n210 VSUBS 0.009175f
C264 B.n211 VSUBS 0.009175f
C265 B.n212 VSUBS 0.009175f
C266 B.n213 VSUBS 0.009175f
C267 B.n214 VSUBS 0.009175f
C268 B.n215 VSUBS 0.009175f
C269 B.n216 VSUBS 0.009175f
C270 B.n217 VSUBS 0.009175f
C271 B.n218 VSUBS 0.009175f
C272 B.n219 VSUBS 0.009175f
C273 B.n220 VSUBS 0.009175f
C274 B.n221 VSUBS 0.009175f
C275 B.n222 VSUBS 0.009175f
C276 B.n223 VSUBS 0.009175f
C277 B.n224 VSUBS 0.009175f
C278 B.n225 VSUBS 0.009175f
C279 B.n226 VSUBS 0.009175f
C280 B.n227 VSUBS 0.009175f
C281 B.n228 VSUBS 0.009175f
C282 B.n229 VSUBS 0.009175f
C283 B.n230 VSUBS 0.009175f
C284 B.n231 VSUBS 0.022719f
C285 B.n232 VSUBS 0.021664f
C286 B.n233 VSUBS 0.02205f
C287 B.n234 VSUBS 0.009175f
C288 B.n235 VSUBS 0.009175f
C289 B.n236 VSUBS 0.009175f
C290 B.n237 VSUBS 0.009175f
C291 B.n238 VSUBS 0.009175f
C292 B.n239 VSUBS 0.009175f
C293 B.n240 VSUBS 0.009175f
C294 B.n241 VSUBS 0.009175f
C295 B.n242 VSUBS 0.009175f
C296 B.n243 VSUBS 0.009175f
C297 B.n244 VSUBS 0.009175f
C298 B.n245 VSUBS 0.009175f
C299 B.n246 VSUBS 0.009175f
C300 B.n247 VSUBS 0.009175f
C301 B.n248 VSUBS 0.009175f
C302 B.n249 VSUBS 0.009175f
C303 B.n250 VSUBS 0.009175f
C304 B.n251 VSUBS 0.009175f
C305 B.n252 VSUBS 0.009175f
C306 B.n253 VSUBS 0.009175f
C307 B.n254 VSUBS 0.009175f
C308 B.n255 VSUBS 0.009175f
C309 B.n256 VSUBS 0.009175f
C310 B.n257 VSUBS 0.009175f
C311 B.n258 VSUBS 0.009175f
C312 B.n259 VSUBS 0.009175f
C313 B.n260 VSUBS 0.009175f
C314 B.n261 VSUBS 0.009175f
C315 B.n262 VSUBS 0.009175f
C316 B.n263 VSUBS 0.009175f
C317 B.n264 VSUBS 0.009175f
C318 B.n265 VSUBS 0.009175f
C319 B.n266 VSUBS 0.009175f
C320 B.n267 VSUBS 0.009175f
C321 B.n268 VSUBS 0.009175f
C322 B.n269 VSUBS 0.009175f
C323 B.n270 VSUBS 0.009175f
C324 B.n271 VSUBS 0.009175f
C325 B.n272 VSUBS 0.009175f
C326 B.n273 VSUBS 0.020995f
C327 B.n274 VSUBS 0.020995f
C328 B.n275 VSUBS 0.022719f
C329 B.n276 VSUBS 0.009175f
C330 B.n277 VSUBS 0.009175f
C331 B.n278 VSUBS 0.009175f
C332 B.n279 VSUBS 0.009175f
C333 B.n280 VSUBS 0.009175f
C334 B.n281 VSUBS 0.009175f
C335 B.n282 VSUBS 0.009175f
C336 B.n283 VSUBS 0.009175f
C337 B.n284 VSUBS 0.009175f
C338 B.n285 VSUBS 0.009175f
C339 B.n286 VSUBS 0.009175f
C340 B.n287 VSUBS 0.009175f
C341 B.n288 VSUBS 0.009175f
C342 B.n289 VSUBS 0.009175f
C343 B.n290 VSUBS 0.009175f
C344 B.n291 VSUBS 0.009175f
C345 B.n292 VSUBS 0.009175f
C346 B.n293 VSUBS 0.009175f
C347 B.n294 VSUBS 0.009175f
C348 B.n295 VSUBS 0.009175f
C349 B.n296 VSUBS 0.009175f
C350 B.n297 VSUBS 0.009175f
C351 B.n298 VSUBS 0.009175f
C352 B.n299 VSUBS 0.009175f
C353 B.n300 VSUBS 0.009175f
C354 B.n301 VSUBS 0.009175f
C355 B.n302 VSUBS 0.009175f
C356 B.n303 VSUBS 0.009175f
C357 B.n304 VSUBS 0.009175f
C358 B.n305 VSUBS 0.009175f
C359 B.n306 VSUBS 0.009175f
C360 B.n307 VSUBS 0.009175f
C361 B.n308 VSUBS 0.009175f
C362 B.n309 VSUBS 0.009175f
C363 B.n310 VSUBS 0.009175f
C364 B.n311 VSUBS 0.009175f
C365 B.n312 VSUBS 0.009175f
C366 B.n313 VSUBS 0.009175f
C367 B.n314 VSUBS 0.009175f
C368 B.n315 VSUBS 0.009175f
C369 B.n316 VSUBS 0.009175f
C370 B.n317 VSUBS 0.009175f
C371 B.n318 VSUBS 0.008365f
C372 B.n319 VSUBS 0.009175f
C373 B.n320 VSUBS 0.009175f
C374 B.n321 VSUBS 0.009175f
C375 B.n322 VSUBS 0.009175f
C376 B.n323 VSUBS 0.009175f
C377 B.n324 VSUBS 0.009175f
C378 B.n325 VSUBS 0.009175f
C379 B.n326 VSUBS 0.009175f
C380 B.n327 VSUBS 0.009175f
C381 B.n328 VSUBS 0.009175f
C382 B.n329 VSUBS 0.009175f
C383 B.n330 VSUBS 0.009175f
C384 B.n331 VSUBS 0.009175f
C385 B.n332 VSUBS 0.009175f
C386 B.n333 VSUBS 0.009175f
C387 B.n334 VSUBS 0.005397f
C388 B.n335 VSUBS 0.021257f
C389 B.n336 VSUBS 0.008365f
C390 B.n337 VSUBS 0.009175f
C391 B.n338 VSUBS 0.009175f
C392 B.n339 VSUBS 0.009175f
C393 B.n340 VSUBS 0.009175f
C394 B.n341 VSUBS 0.009175f
C395 B.n342 VSUBS 0.009175f
C396 B.n343 VSUBS 0.009175f
C397 B.n344 VSUBS 0.009175f
C398 B.n345 VSUBS 0.009175f
C399 B.n346 VSUBS 0.009175f
C400 B.n347 VSUBS 0.009175f
C401 B.n348 VSUBS 0.009175f
C402 B.n349 VSUBS 0.009175f
C403 B.n350 VSUBS 0.009175f
C404 B.n351 VSUBS 0.009175f
C405 B.n352 VSUBS 0.009175f
C406 B.n353 VSUBS 0.009175f
C407 B.n354 VSUBS 0.009175f
C408 B.n355 VSUBS 0.009175f
C409 B.n356 VSUBS 0.009175f
C410 B.n357 VSUBS 0.009175f
C411 B.n358 VSUBS 0.009175f
C412 B.n359 VSUBS 0.009175f
C413 B.n360 VSUBS 0.009175f
C414 B.n361 VSUBS 0.009175f
C415 B.n362 VSUBS 0.009175f
C416 B.n363 VSUBS 0.009175f
C417 B.n364 VSUBS 0.009175f
C418 B.n365 VSUBS 0.009175f
C419 B.n366 VSUBS 0.009175f
C420 B.n367 VSUBS 0.009175f
C421 B.n368 VSUBS 0.009175f
C422 B.n369 VSUBS 0.009175f
C423 B.n370 VSUBS 0.009175f
C424 B.n371 VSUBS 0.009175f
C425 B.n372 VSUBS 0.009175f
C426 B.n373 VSUBS 0.009175f
C427 B.n374 VSUBS 0.009175f
C428 B.n375 VSUBS 0.009175f
C429 B.n376 VSUBS 0.009175f
C430 B.n377 VSUBS 0.009175f
C431 B.n378 VSUBS 0.009175f
C432 B.n379 VSUBS 0.022719f
C433 B.n380 VSUBS 0.022719f
C434 B.n381 VSUBS 0.020995f
C435 B.n382 VSUBS 0.009175f
C436 B.n383 VSUBS 0.009175f
C437 B.n384 VSUBS 0.009175f
C438 B.n385 VSUBS 0.009175f
C439 B.n386 VSUBS 0.009175f
C440 B.n387 VSUBS 0.009175f
C441 B.n388 VSUBS 0.009175f
C442 B.n389 VSUBS 0.009175f
C443 B.n390 VSUBS 0.009175f
C444 B.n391 VSUBS 0.009175f
C445 B.n392 VSUBS 0.009175f
C446 B.n393 VSUBS 0.009175f
C447 B.n394 VSUBS 0.009175f
C448 B.n395 VSUBS 0.009175f
C449 B.n396 VSUBS 0.009175f
C450 B.n397 VSUBS 0.009175f
C451 B.n398 VSUBS 0.009175f
C452 B.n399 VSUBS 0.011973f
C453 B.n400 VSUBS 0.012754f
C454 B.n401 VSUBS 0.025362f
C455 VTAIL.n0 VSUBS 0.026108f
C456 VTAIL.n1 VSUBS 0.023759f
C457 VTAIL.n2 VSUBS 0.012767f
C458 VTAIL.n3 VSUBS 0.030177f
C459 VTAIL.n4 VSUBS 0.013518f
C460 VTAIL.n5 VSUBS 0.023759f
C461 VTAIL.n6 VSUBS 0.012767f
C462 VTAIL.n7 VSUBS 0.030177f
C463 VTAIL.n8 VSUBS 0.013518f
C464 VTAIL.n9 VSUBS 0.023759f
C465 VTAIL.n10 VSUBS 0.012767f
C466 VTAIL.n11 VSUBS 0.030177f
C467 VTAIL.n12 VSUBS 0.013518f
C468 VTAIL.n13 VSUBS 0.118919f
C469 VTAIL.t2 VSUBS 0.064337f
C470 VTAIL.n14 VSUBS 0.022633f
C471 VTAIL.n15 VSUBS 0.019197f
C472 VTAIL.n16 VSUBS 0.012767f
C473 VTAIL.n17 VSUBS 0.767156f
C474 VTAIL.n18 VSUBS 0.023759f
C475 VTAIL.n19 VSUBS 0.012767f
C476 VTAIL.n20 VSUBS 0.013518f
C477 VTAIL.n21 VSUBS 0.030177f
C478 VTAIL.n22 VSUBS 0.030177f
C479 VTAIL.n23 VSUBS 0.013518f
C480 VTAIL.n24 VSUBS 0.012767f
C481 VTAIL.n25 VSUBS 0.023759f
C482 VTAIL.n26 VSUBS 0.023759f
C483 VTAIL.n27 VSUBS 0.012767f
C484 VTAIL.n28 VSUBS 0.013518f
C485 VTAIL.n29 VSUBS 0.030177f
C486 VTAIL.n30 VSUBS 0.030177f
C487 VTAIL.n31 VSUBS 0.013518f
C488 VTAIL.n32 VSUBS 0.012767f
C489 VTAIL.n33 VSUBS 0.023759f
C490 VTAIL.n34 VSUBS 0.023759f
C491 VTAIL.n35 VSUBS 0.012767f
C492 VTAIL.n36 VSUBS 0.013518f
C493 VTAIL.n37 VSUBS 0.030177f
C494 VTAIL.n38 VSUBS 0.07306f
C495 VTAIL.n39 VSUBS 0.013518f
C496 VTAIL.n40 VSUBS 0.012767f
C497 VTAIL.n41 VSUBS 0.051348f
C498 VTAIL.n42 VSUBS 0.036628f
C499 VTAIL.n43 VSUBS 0.079823f
C500 VTAIL.n44 VSUBS 0.026108f
C501 VTAIL.n45 VSUBS 0.023759f
C502 VTAIL.n46 VSUBS 0.012767f
C503 VTAIL.n47 VSUBS 0.030177f
C504 VTAIL.n48 VSUBS 0.013518f
C505 VTAIL.n49 VSUBS 0.023759f
C506 VTAIL.n50 VSUBS 0.012767f
C507 VTAIL.n51 VSUBS 0.030177f
C508 VTAIL.n52 VSUBS 0.013518f
C509 VTAIL.n53 VSUBS 0.023759f
C510 VTAIL.n54 VSUBS 0.012767f
C511 VTAIL.n55 VSUBS 0.030177f
C512 VTAIL.n56 VSUBS 0.013518f
C513 VTAIL.n57 VSUBS 0.118919f
C514 VTAIL.t6 VSUBS 0.064337f
C515 VTAIL.n58 VSUBS 0.022633f
C516 VTAIL.n59 VSUBS 0.019197f
C517 VTAIL.n60 VSUBS 0.012767f
C518 VTAIL.n61 VSUBS 0.767156f
C519 VTAIL.n62 VSUBS 0.023759f
C520 VTAIL.n63 VSUBS 0.012767f
C521 VTAIL.n64 VSUBS 0.013518f
C522 VTAIL.n65 VSUBS 0.030177f
C523 VTAIL.n66 VSUBS 0.030177f
C524 VTAIL.n67 VSUBS 0.013518f
C525 VTAIL.n68 VSUBS 0.012767f
C526 VTAIL.n69 VSUBS 0.023759f
C527 VTAIL.n70 VSUBS 0.023759f
C528 VTAIL.n71 VSUBS 0.012767f
C529 VTAIL.n72 VSUBS 0.013518f
C530 VTAIL.n73 VSUBS 0.030177f
C531 VTAIL.n74 VSUBS 0.030177f
C532 VTAIL.n75 VSUBS 0.013518f
C533 VTAIL.n76 VSUBS 0.012767f
C534 VTAIL.n77 VSUBS 0.023759f
C535 VTAIL.n78 VSUBS 0.023759f
C536 VTAIL.n79 VSUBS 0.012767f
C537 VTAIL.n80 VSUBS 0.013518f
C538 VTAIL.n81 VSUBS 0.030177f
C539 VTAIL.n82 VSUBS 0.07306f
C540 VTAIL.n83 VSUBS 0.013518f
C541 VTAIL.n84 VSUBS 0.012767f
C542 VTAIL.n85 VSUBS 0.051348f
C543 VTAIL.n86 VSUBS 0.036628f
C544 VTAIL.n87 VSUBS 0.096488f
C545 VTAIL.n88 VSUBS 0.026108f
C546 VTAIL.n89 VSUBS 0.023759f
C547 VTAIL.n90 VSUBS 0.012767f
C548 VTAIL.n91 VSUBS 0.030177f
C549 VTAIL.n92 VSUBS 0.013518f
C550 VTAIL.n93 VSUBS 0.023759f
C551 VTAIL.n94 VSUBS 0.012767f
C552 VTAIL.n95 VSUBS 0.030177f
C553 VTAIL.n96 VSUBS 0.013518f
C554 VTAIL.n97 VSUBS 0.023759f
C555 VTAIL.n98 VSUBS 0.012767f
C556 VTAIL.n99 VSUBS 0.030177f
C557 VTAIL.n100 VSUBS 0.013518f
C558 VTAIL.n101 VSUBS 0.118919f
C559 VTAIL.t7 VSUBS 0.064337f
C560 VTAIL.n102 VSUBS 0.022633f
C561 VTAIL.n103 VSUBS 0.019197f
C562 VTAIL.n104 VSUBS 0.012767f
C563 VTAIL.n105 VSUBS 0.767156f
C564 VTAIL.n106 VSUBS 0.023759f
C565 VTAIL.n107 VSUBS 0.012767f
C566 VTAIL.n108 VSUBS 0.013518f
C567 VTAIL.n109 VSUBS 0.030177f
C568 VTAIL.n110 VSUBS 0.030177f
C569 VTAIL.n111 VSUBS 0.013518f
C570 VTAIL.n112 VSUBS 0.012767f
C571 VTAIL.n113 VSUBS 0.023759f
C572 VTAIL.n114 VSUBS 0.023759f
C573 VTAIL.n115 VSUBS 0.012767f
C574 VTAIL.n116 VSUBS 0.013518f
C575 VTAIL.n117 VSUBS 0.030177f
C576 VTAIL.n118 VSUBS 0.030177f
C577 VTAIL.n119 VSUBS 0.013518f
C578 VTAIL.n120 VSUBS 0.012767f
C579 VTAIL.n121 VSUBS 0.023759f
C580 VTAIL.n122 VSUBS 0.023759f
C581 VTAIL.n123 VSUBS 0.012767f
C582 VTAIL.n124 VSUBS 0.013518f
C583 VTAIL.n125 VSUBS 0.030177f
C584 VTAIL.n126 VSUBS 0.07306f
C585 VTAIL.n127 VSUBS 0.013518f
C586 VTAIL.n128 VSUBS 0.012767f
C587 VTAIL.n129 VSUBS 0.051348f
C588 VTAIL.n130 VSUBS 0.036628f
C589 VTAIL.n131 VSUBS 0.958099f
C590 VTAIL.n132 VSUBS 0.026108f
C591 VTAIL.n133 VSUBS 0.023759f
C592 VTAIL.n134 VSUBS 0.012767f
C593 VTAIL.n135 VSUBS 0.030177f
C594 VTAIL.n136 VSUBS 0.013518f
C595 VTAIL.n137 VSUBS 0.023759f
C596 VTAIL.n138 VSUBS 0.012767f
C597 VTAIL.n139 VSUBS 0.030177f
C598 VTAIL.n140 VSUBS 0.013518f
C599 VTAIL.n141 VSUBS 0.023759f
C600 VTAIL.n142 VSUBS 0.012767f
C601 VTAIL.n143 VSUBS 0.030177f
C602 VTAIL.n144 VSUBS 0.013518f
C603 VTAIL.n145 VSUBS 0.118919f
C604 VTAIL.t0 VSUBS 0.064337f
C605 VTAIL.n146 VSUBS 0.022633f
C606 VTAIL.n147 VSUBS 0.019197f
C607 VTAIL.n148 VSUBS 0.012767f
C608 VTAIL.n149 VSUBS 0.767156f
C609 VTAIL.n150 VSUBS 0.023759f
C610 VTAIL.n151 VSUBS 0.012767f
C611 VTAIL.n152 VSUBS 0.013518f
C612 VTAIL.n153 VSUBS 0.030177f
C613 VTAIL.n154 VSUBS 0.030177f
C614 VTAIL.n155 VSUBS 0.013518f
C615 VTAIL.n156 VSUBS 0.012767f
C616 VTAIL.n157 VSUBS 0.023759f
C617 VTAIL.n158 VSUBS 0.023759f
C618 VTAIL.n159 VSUBS 0.012767f
C619 VTAIL.n160 VSUBS 0.013518f
C620 VTAIL.n161 VSUBS 0.030177f
C621 VTAIL.n162 VSUBS 0.030177f
C622 VTAIL.n163 VSUBS 0.013518f
C623 VTAIL.n164 VSUBS 0.012767f
C624 VTAIL.n165 VSUBS 0.023759f
C625 VTAIL.n166 VSUBS 0.023759f
C626 VTAIL.n167 VSUBS 0.012767f
C627 VTAIL.n168 VSUBS 0.013518f
C628 VTAIL.n169 VSUBS 0.030177f
C629 VTAIL.n170 VSUBS 0.07306f
C630 VTAIL.n171 VSUBS 0.013518f
C631 VTAIL.n172 VSUBS 0.012767f
C632 VTAIL.n173 VSUBS 0.051348f
C633 VTAIL.n174 VSUBS 0.036628f
C634 VTAIL.n175 VSUBS 0.958099f
C635 VTAIL.n176 VSUBS 0.026108f
C636 VTAIL.n177 VSUBS 0.023759f
C637 VTAIL.n178 VSUBS 0.012767f
C638 VTAIL.n179 VSUBS 0.030177f
C639 VTAIL.n180 VSUBS 0.013518f
C640 VTAIL.n181 VSUBS 0.023759f
C641 VTAIL.n182 VSUBS 0.012767f
C642 VTAIL.n183 VSUBS 0.030177f
C643 VTAIL.n184 VSUBS 0.013518f
C644 VTAIL.n185 VSUBS 0.023759f
C645 VTAIL.n186 VSUBS 0.012767f
C646 VTAIL.n187 VSUBS 0.030177f
C647 VTAIL.n188 VSUBS 0.013518f
C648 VTAIL.n189 VSUBS 0.118919f
C649 VTAIL.t1 VSUBS 0.064337f
C650 VTAIL.n190 VSUBS 0.022633f
C651 VTAIL.n191 VSUBS 0.019197f
C652 VTAIL.n192 VSUBS 0.012767f
C653 VTAIL.n193 VSUBS 0.767156f
C654 VTAIL.n194 VSUBS 0.023759f
C655 VTAIL.n195 VSUBS 0.012767f
C656 VTAIL.n196 VSUBS 0.013518f
C657 VTAIL.n197 VSUBS 0.030177f
C658 VTAIL.n198 VSUBS 0.030177f
C659 VTAIL.n199 VSUBS 0.013518f
C660 VTAIL.n200 VSUBS 0.012767f
C661 VTAIL.n201 VSUBS 0.023759f
C662 VTAIL.n202 VSUBS 0.023759f
C663 VTAIL.n203 VSUBS 0.012767f
C664 VTAIL.n204 VSUBS 0.013518f
C665 VTAIL.n205 VSUBS 0.030177f
C666 VTAIL.n206 VSUBS 0.030177f
C667 VTAIL.n207 VSUBS 0.013518f
C668 VTAIL.n208 VSUBS 0.012767f
C669 VTAIL.n209 VSUBS 0.023759f
C670 VTAIL.n210 VSUBS 0.023759f
C671 VTAIL.n211 VSUBS 0.012767f
C672 VTAIL.n212 VSUBS 0.013518f
C673 VTAIL.n213 VSUBS 0.030177f
C674 VTAIL.n214 VSUBS 0.07306f
C675 VTAIL.n215 VSUBS 0.013518f
C676 VTAIL.n216 VSUBS 0.012767f
C677 VTAIL.n217 VSUBS 0.051348f
C678 VTAIL.n218 VSUBS 0.036628f
C679 VTAIL.n219 VSUBS 0.096488f
C680 VTAIL.n220 VSUBS 0.026108f
C681 VTAIL.n221 VSUBS 0.023759f
C682 VTAIL.n222 VSUBS 0.012767f
C683 VTAIL.n223 VSUBS 0.030177f
C684 VTAIL.n224 VSUBS 0.013518f
C685 VTAIL.n225 VSUBS 0.023759f
C686 VTAIL.n226 VSUBS 0.012767f
C687 VTAIL.n227 VSUBS 0.030177f
C688 VTAIL.n228 VSUBS 0.013518f
C689 VTAIL.n229 VSUBS 0.023759f
C690 VTAIL.n230 VSUBS 0.012767f
C691 VTAIL.n231 VSUBS 0.030177f
C692 VTAIL.n232 VSUBS 0.013518f
C693 VTAIL.n233 VSUBS 0.118919f
C694 VTAIL.t4 VSUBS 0.064337f
C695 VTAIL.n234 VSUBS 0.022633f
C696 VTAIL.n235 VSUBS 0.019197f
C697 VTAIL.n236 VSUBS 0.012767f
C698 VTAIL.n237 VSUBS 0.767156f
C699 VTAIL.n238 VSUBS 0.023759f
C700 VTAIL.n239 VSUBS 0.012767f
C701 VTAIL.n240 VSUBS 0.013518f
C702 VTAIL.n241 VSUBS 0.030177f
C703 VTAIL.n242 VSUBS 0.030177f
C704 VTAIL.n243 VSUBS 0.013518f
C705 VTAIL.n244 VSUBS 0.012767f
C706 VTAIL.n245 VSUBS 0.023759f
C707 VTAIL.n246 VSUBS 0.023759f
C708 VTAIL.n247 VSUBS 0.012767f
C709 VTAIL.n248 VSUBS 0.013518f
C710 VTAIL.n249 VSUBS 0.030177f
C711 VTAIL.n250 VSUBS 0.030177f
C712 VTAIL.n251 VSUBS 0.013518f
C713 VTAIL.n252 VSUBS 0.012767f
C714 VTAIL.n253 VSUBS 0.023759f
C715 VTAIL.n254 VSUBS 0.023759f
C716 VTAIL.n255 VSUBS 0.012767f
C717 VTAIL.n256 VSUBS 0.013518f
C718 VTAIL.n257 VSUBS 0.030177f
C719 VTAIL.n258 VSUBS 0.07306f
C720 VTAIL.n259 VSUBS 0.013518f
C721 VTAIL.n260 VSUBS 0.012767f
C722 VTAIL.n261 VSUBS 0.051348f
C723 VTAIL.n262 VSUBS 0.036628f
C724 VTAIL.n263 VSUBS 0.096488f
C725 VTAIL.n264 VSUBS 0.026108f
C726 VTAIL.n265 VSUBS 0.023759f
C727 VTAIL.n266 VSUBS 0.012767f
C728 VTAIL.n267 VSUBS 0.030177f
C729 VTAIL.n268 VSUBS 0.013518f
C730 VTAIL.n269 VSUBS 0.023759f
C731 VTAIL.n270 VSUBS 0.012767f
C732 VTAIL.n271 VSUBS 0.030177f
C733 VTAIL.n272 VSUBS 0.013518f
C734 VTAIL.n273 VSUBS 0.023759f
C735 VTAIL.n274 VSUBS 0.012767f
C736 VTAIL.n275 VSUBS 0.030177f
C737 VTAIL.n276 VSUBS 0.013518f
C738 VTAIL.n277 VSUBS 0.118919f
C739 VTAIL.t5 VSUBS 0.064337f
C740 VTAIL.n278 VSUBS 0.022633f
C741 VTAIL.n279 VSUBS 0.019197f
C742 VTAIL.n280 VSUBS 0.012767f
C743 VTAIL.n281 VSUBS 0.767156f
C744 VTAIL.n282 VSUBS 0.023759f
C745 VTAIL.n283 VSUBS 0.012767f
C746 VTAIL.n284 VSUBS 0.013518f
C747 VTAIL.n285 VSUBS 0.030177f
C748 VTAIL.n286 VSUBS 0.030177f
C749 VTAIL.n287 VSUBS 0.013518f
C750 VTAIL.n288 VSUBS 0.012767f
C751 VTAIL.n289 VSUBS 0.023759f
C752 VTAIL.n290 VSUBS 0.023759f
C753 VTAIL.n291 VSUBS 0.012767f
C754 VTAIL.n292 VSUBS 0.013518f
C755 VTAIL.n293 VSUBS 0.030177f
C756 VTAIL.n294 VSUBS 0.030177f
C757 VTAIL.n295 VSUBS 0.013518f
C758 VTAIL.n296 VSUBS 0.012767f
C759 VTAIL.n297 VSUBS 0.023759f
C760 VTAIL.n298 VSUBS 0.023759f
C761 VTAIL.n299 VSUBS 0.012767f
C762 VTAIL.n300 VSUBS 0.013518f
C763 VTAIL.n301 VSUBS 0.030177f
C764 VTAIL.n302 VSUBS 0.07306f
C765 VTAIL.n303 VSUBS 0.013518f
C766 VTAIL.n304 VSUBS 0.012767f
C767 VTAIL.n305 VSUBS 0.051348f
C768 VTAIL.n306 VSUBS 0.036628f
C769 VTAIL.n307 VSUBS 0.958099f
C770 VTAIL.n308 VSUBS 0.026108f
C771 VTAIL.n309 VSUBS 0.023759f
C772 VTAIL.n310 VSUBS 0.012767f
C773 VTAIL.n311 VSUBS 0.030177f
C774 VTAIL.n312 VSUBS 0.013518f
C775 VTAIL.n313 VSUBS 0.023759f
C776 VTAIL.n314 VSUBS 0.012767f
C777 VTAIL.n315 VSUBS 0.030177f
C778 VTAIL.n316 VSUBS 0.013518f
C779 VTAIL.n317 VSUBS 0.023759f
C780 VTAIL.n318 VSUBS 0.012767f
C781 VTAIL.n319 VSUBS 0.030177f
C782 VTAIL.n320 VSUBS 0.013518f
C783 VTAIL.n321 VSUBS 0.118919f
C784 VTAIL.t3 VSUBS 0.064337f
C785 VTAIL.n322 VSUBS 0.022633f
C786 VTAIL.n323 VSUBS 0.019197f
C787 VTAIL.n324 VSUBS 0.012767f
C788 VTAIL.n325 VSUBS 0.767156f
C789 VTAIL.n326 VSUBS 0.023759f
C790 VTAIL.n327 VSUBS 0.012767f
C791 VTAIL.n328 VSUBS 0.013518f
C792 VTAIL.n329 VSUBS 0.030177f
C793 VTAIL.n330 VSUBS 0.030177f
C794 VTAIL.n331 VSUBS 0.013518f
C795 VTAIL.n332 VSUBS 0.012767f
C796 VTAIL.n333 VSUBS 0.023759f
C797 VTAIL.n334 VSUBS 0.023759f
C798 VTAIL.n335 VSUBS 0.012767f
C799 VTAIL.n336 VSUBS 0.013518f
C800 VTAIL.n337 VSUBS 0.030177f
C801 VTAIL.n338 VSUBS 0.030177f
C802 VTAIL.n339 VSUBS 0.013518f
C803 VTAIL.n340 VSUBS 0.012767f
C804 VTAIL.n341 VSUBS 0.023759f
C805 VTAIL.n342 VSUBS 0.023759f
C806 VTAIL.n343 VSUBS 0.012767f
C807 VTAIL.n344 VSUBS 0.013518f
C808 VTAIL.n345 VSUBS 0.030177f
C809 VTAIL.n346 VSUBS 0.07306f
C810 VTAIL.n347 VSUBS 0.013518f
C811 VTAIL.n348 VSUBS 0.012767f
C812 VTAIL.n349 VSUBS 0.051348f
C813 VTAIL.n350 VSUBS 0.036628f
C814 VTAIL.n351 VSUBS 0.932525f
C815 VDD1.t0 VSUBS 0.164773f
C816 VDD1.t3 VSUBS 0.164773f
C817 VDD1.n0 VSUBS 1.17185f
C818 VDD1.t1 VSUBS 0.164773f
C819 VDD1.t2 VSUBS 0.164773f
C820 VDD1.n1 VSUBS 1.614f
C821 VP.t3 VSUBS 0.257996f
C822 VP.t2 VSUBS 0.257996f
C823 VP.n0 VSUBS 0.431954f
C824 VP.t0 VSUBS 0.257996f
C825 VP.t1 VSUBS 0.257996f
C826 VP.n1 VSUBS 0.2215f
C827 VP.n2 VSUBS 2.09673f
.ends

