* NGSPICE file created from diff_pair_sample_1572.ext - technology: sky130A

.subckt diff_pair_sample_1572 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.936 ps=5.58 w=2.4 l=2.22
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.936 ps=5.58 w=2.4 l=2.22
X2 B.t11 B.t9 B.t10 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=2.22
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.936 ps=5.58 w=2.4 l=2.22
X4 B.t8 B.t6 B.t7 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=2.22
X5 B.t5 B.t3 B.t4 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=2.22
X6 VDD1.t0 VP.t1 VTAIL.t0 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.936 ps=5.58 w=2.4 l=2.22
X7 B.t2 B.t0 B.t1 w_n1990_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=2.22
R0 VN VN.t1 111.743
R1 VN VN.t0 75.6059
R2 VTAIL.n42 VTAIL.n36 756.745
R3 VTAIL.n6 VTAIL.n0 756.745
R4 VTAIL.n30 VTAIL.n24 756.745
R5 VTAIL.n18 VTAIL.n12 756.745
R6 VTAIL.n41 VTAIL.n40 585
R7 VTAIL.n43 VTAIL.n42 585
R8 VTAIL.n5 VTAIL.n4 585
R9 VTAIL.n7 VTAIL.n6 585
R10 VTAIL.n31 VTAIL.n30 585
R11 VTAIL.n29 VTAIL.n28 585
R12 VTAIL.n19 VTAIL.n18 585
R13 VTAIL.n17 VTAIL.n16 585
R14 VTAIL.n39 VTAIL.t3 355.474
R15 VTAIL.n3 VTAIL.t1 355.474
R16 VTAIL.n27 VTAIL.t0 355.474
R17 VTAIL.n15 VTAIL.t2 355.474
R18 VTAIL.n42 VTAIL.n41 171.744
R19 VTAIL.n6 VTAIL.n5 171.744
R20 VTAIL.n30 VTAIL.n29 171.744
R21 VTAIL.n18 VTAIL.n17 171.744
R22 VTAIL.n41 VTAIL.t3 85.8723
R23 VTAIL.n5 VTAIL.t1 85.8723
R24 VTAIL.n29 VTAIL.t0 85.8723
R25 VTAIL.n17 VTAIL.t2 85.8723
R26 VTAIL.n47 VTAIL.n46 32.1853
R27 VTAIL.n11 VTAIL.n10 32.1853
R28 VTAIL.n35 VTAIL.n34 32.1853
R29 VTAIL.n23 VTAIL.n22 32.1853
R30 VTAIL.n23 VTAIL.n11 18.8324
R31 VTAIL.n47 VTAIL.n35 16.6341
R32 VTAIL.n40 VTAIL.n39 15.8418
R33 VTAIL.n4 VTAIL.n3 15.8418
R34 VTAIL.n28 VTAIL.n27 15.8418
R35 VTAIL.n16 VTAIL.n15 15.8418
R36 VTAIL.n43 VTAIL.n38 12.8005
R37 VTAIL.n7 VTAIL.n2 12.8005
R38 VTAIL.n31 VTAIL.n26 12.8005
R39 VTAIL.n19 VTAIL.n14 12.8005
R40 VTAIL.n44 VTAIL.n36 12.0247
R41 VTAIL.n8 VTAIL.n0 12.0247
R42 VTAIL.n32 VTAIL.n24 12.0247
R43 VTAIL.n20 VTAIL.n12 12.0247
R44 VTAIL.n46 VTAIL.n45 9.45567
R45 VTAIL.n10 VTAIL.n9 9.45567
R46 VTAIL.n34 VTAIL.n33 9.45567
R47 VTAIL.n22 VTAIL.n21 9.45567
R48 VTAIL.n45 VTAIL.n44 9.3005
R49 VTAIL.n38 VTAIL.n37 9.3005
R50 VTAIL.n9 VTAIL.n8 9.3005
R51 VTAIL.n2 VTAIL.n1 9.3005
R52 VTAIL.n33 VTAIL.n32 9.3005
R53 VTAIL.n26 VTAIL.n25 9.3005
R54 VTAIL.n21 VTAIL.n20 9.3005
R55 VTAIL.n14 VTAIL.n13 9.3005
R56 VTAIL.n27 VTAIL.n25 4.29255
R57 VTAIL.n15 VTAIL.n13 4.29255
R58 VTAIL.n39 VTAIL.n37 4.29255
R59 VTAIL.n3 VTAIL.n1 4.29255
R60 VTAIL.n46 VTAIL.n36 1.93989
R61 VTAIL.n10 VTAIL.n0 1.93989
R62 VTAIL.n34 VTAIL.n24 1.93989
R63 VTAIL.n22 VTAIL.n12 1.93989
R64 VTAIL.n35 VTAIL.n23 1.56947
R65 VTAIL.n44 VTAIL.n43 1.16414
R66 VTAIL.n8 VTAIL.n7 1.16414
R67 VTAIL.n32 VTAIL.n31 1.16414
R68 VTAIL.n20 VTAIL.n19 1.16414
R69 VTAIL VTAIL.n11 1.07809
R70 VTAIL VTAIL.n47 0.491879
R71 VTAIL.n40 VTAIL.n38 0.388379
R72 VTAIL.n4 VTAIL.n2 0.388379
R73 VTAIL.n28 VTAIL.n26 0.388379
R74 VTAIL.n16 VTAIL.n14 0.388379
R75 VTAIL.n45 VTAIL.n37 0.155672
R76 VTAIL.n9 VTAIL.n1 0.155672
R77 VTAIL.n33 VTAIL.n25 0.155672
R78 VTAIL.n21 VTAIL.n13 0.155672
R79 VDD2.n17 VDD2.n11 756.745
R80 VDD2.n6 VDD2.n0 756.745
R81 VDD2.n18 VDD2.n17 585
R82 VDD2.n16 VDD2.n15 585
R83 VDD2.n5 VDD2.n4 585
R84 VDD2.n7 VDD2.n6 585
R85 VDD2.n14 VDD2.t0 355.474
R86 VDD2.n3 VDD2.t1 355.474
R87 VDD2.n17 VDD2.n16 171.744
R88 VDD2.n6 VDD2.n5 171.744
R89 VDD2.n16 VDD2.t0 85.8723
R90 VDD2.n5 VDD2.t1 85.8723
R91 VDD2.n22 VDD2.n10 78.9891
R92 VDD2.n22 VDD2.n21 48.8641
R93 VDD2.n15 VDD2.n14 15.8418
R94 VDD2.n4 VDD2.n3 15.8418
R95 VDD2.n18 VDD2.n13 12.8005
R96 VDD2.n7 VDD2.n2 12.8005
R97 VDD2.n19 VDD2.n11 12.0247
R98 VDD2.n8 VDD2.n0 12.0247
R99 VDD2.n21 VDD2.n20 9.45567
R100 VDD2.n10 VDD2.n9 9.45567
R101 VDD2.n20 VDD2.n19 9.3005
R102 VDD2.n13 VDD2.n12 9.3005
R103 VDD2.n9 VDD2.n8 9.3005
R104 VDD2.n2 VDD2.n1 9.3005
R105 VDD2.n14 VDD2.n12 4.29255
R106 VDD2.n3 VDD2.n1 4.29255
R107 VDD2.n21 VDD2.n11 1.93989
R108 VDD2.n10 VDD2.n0 1.93989
R109 VDD2.n19 VDD2.n18 1.16414
R110 VDD2.n8 VDD2.n7 1.16414
R111 VDD2 VDD2.n22 0.608259
R112 VDD2.n15 VDD2.n13 0.388379
R113 VDD2.n4 VDD2.n2 0.388379
R114 VDD2.n20 VDD2.n12 0.155672
R115 VDD2.n9 VDD2.n1 0.155672
R116 VP.n0 VP.t1 111.645
R117 VP.n0 VP.t0 75.2696
R118 VP VP.n0 0.336784
R119 VDD1.n6 VDD1.n0 756.745
R120 VDD1.n17 VDD1.n11 756.745
R121 VDD1.n7 VDD1.n6 585
R122 VDD1.n5 VDD1.n4 585
R123 VDD1.n16 VDD1.n15 585
R124 VDD1.n18 VDD1.n17 585
R125 VDD1.n3 VDD1.t0 355.474
R126 VDD1.n14 VDD1.t1 355.474
R127 VDD1.n6 VDD1.n5 171.744
R128 VDD1.n17 VDD1.n16 171.744
R129 VDD1.n5 VDD1.t0 85.8723
R130 VDD1.n16 VDD1.t1 85.8723
R131 VDD1 VDD1.n21 80.0635
R132 VDD1 VDD1.n10 49.4719
R133 VDD1.n4 VDD1.n3 15.8418
R134 VDD1.n15 VDD1.n14 15.8418
R135 VDD1.n7 VDD1.n2 12.8005
R136 VDD1.n18 VDD1.n13 12.8005
R137 VDD1.n8 VDD1.n0 12.0247
R138 VDD1.n19 VDD1.n11 12.0247
R139 VDD1.n10 VDD1.n9 9.45567
R140 VDD1.n21 VDD1.n20 9.45567
R141 VDD1.n9 VDD1.n8 9.3005
R142 VDD1.n2 VDD1.n1 9.3005
R143 VDD1.n20 VDD1.n19 9.3005
R144 VDD1.n13 VDD1.n12 9.3005
R145 VDD1.n3 VDD1.n1 4.29255
R146 VDD1.n14 VDD1.n12 4.29255
R147 VDD1.n10 VDD1.n0 1.93989
R148 VDD1.n21 VDD1.n11 1.93989
R149 VDD1.n8 VDD1.n7 1.16414
R150 VDD1.n19 VDD1.n18 1.16414
R151 VDD1.n4 VDD1.n2 0.388379
R152 VDD1.n15 VDD1.n13 0.388379
R153 VDD1.n9 VDD1.n1 0.155672
R154 VDD1.n20 VDD1.n12 0.155672
R155 B.n253 B.n252 585
R156 B.n254 B.n35 585
R157 B.n256 B.n255 585
R158 B.n257 B.n34 585
R159 B.n259 B.n258 585
R160 B.n260 B.n33 585
R161 B.n262 B.n261 585
R162 B.n263 B.n32 585
R163 B.n265 B.n264 585
R164 B.n266 B.n31 585
R165 B.n268 B.n267 585
R166 B.n269 B.n30 585
R167 B.n271 B.n270 585
R168 B.n273 B.n27 585
R169 B.n275 B.n274 585
R170 B.n276 B.n26 585
R171 B.n278 B.n277 585
R172 B.n279 B.n25 585
R173 B.n281 B.n280 585
R174 B.n282 B.n24 585
R175 B.n284 B.n283 585
R176 B.n285 B.n23 585
R177 B.n287 B.n286 585
R178 B.n289 B.n288 585
R179 B.n290 B.n19 585
R180 B.n292 B.n291 585
R181 B.n293 B.n18 585
R182 B.n295 B.n294 585
R183 B.n296 B.n17 585
R184 B.n298 B.n297 585
R185 B.n299 B.n16 585
R186 B.n301 B.n300 585
R187 B.n302 B.n15 585
R188 B.n304 B.n303 585
R189 B.n305 B.n14 585
R190 B.n307 B.n306 585
R191 B.n251 B.n36 585
R192 B.n250 B.n249 585
R193 B.n248 B.n37 585
R194 B.n247 B.n246 585
R195 B.n245 B.n38 585
R196 B.n244 B.n243 585
R197 B.n242 B.n39 585
R198 B.n241 B.n240 585
R199 B.n239 B.n40 585
R200 B.n238 B.n237 585
R201 B.n236 B.n41 585
R202 B.n235 B.n234 585
R203 B.n233 B.n42 585
R204 B.n232 B.n231 585
R205 B.n230 B.n43 585
R206 B.n229 B.n228 585
R207 B.n227 B.n44 585
R208 B.n226 B.n225 585
R209 B.n224 B.n45 585
R210 B.n223 B.n222 585
R211 B.n221 B.n46 585
R212 B.n220 B.n219 585
R213 B.n218 B.n47 585
R214 B.n217 B.n216 585
R215 B.n215 B.n48 585
R216 B.n214 B.n213 585
R217 B.n212 B.n49 585
R218 B.n211 B.n210 585
R219 B.n209 B.n50 585
R220 B.n208 B.n207 585
R221 B.n206 B.n51 585
R222 B.n205 B.n204 585
R223 B.n203 B.n52 585
R224 B.n202 B.n201 585
R225 B.n200 B.n53 585
R226 B.n199 B.n198 585
R227 B.n197 B.n54 585
R228 B.n196 B.n195 585
R229 B.n194 B.n55 585
R230 B.n193 B.n192 585
R231 B.n191 B.n56 585
R232 B.n190 B.n189 585
R233 B.n188 B.n57 585
R234 B.n187 B.n186 585
R235 B.n185 B.n58 585
R236 B.n184 B.n183 585
R237 B.n182 B.n59 585
R238 B.n127 B.n126 585
R239 B.n128 B.n81 585
R240 B.n130 B.n129 585
R241 B.n131 B.n80 585
R242 B.n133 B.n132 585
R243 B.n134 B.n79 585
R244 B.n136 B.n135 585
R245 B.n137 B.n78 585
R246 B.n139 B.n138 585
R247 B.n140 B.n77 585
R248 B.n142 B.n141 585
R249 B.n143 B.n76 585
R250 B.n145 B.n144 585
R251 B.n147 B.n73 585
R252 B.n149 B.n148 585
R253 B.n150 B.n72 585
R254 B.n152 B.n151 585
R255 B.n153 B.n71 585
R256 B.n155 B.n154 585
R257 B.n156 B.n70 585
R258 B.n158 B.n157 585
R259 B.n159 B.n69 585
R260 B.n161 B.n160 585
R261 B.n163 B.n162 585
R262 B.n164 B.n65 585
R263 B.n166 B.n165 585
R264 B.n167 B.n64 585
R265 B.n169 B.n168 585
R266 B.n170 B.n63 585
R267 B.n172 B.n171 585
R268 B.n173 B.n62 585
R269 B.n175 B.n174 585
R270 B.n176 B.n61 585
R271 B.n178 B.n177 585
R272 B.n179 B.n60 585
R273 B.n181 B.n180 585
R274 B.n125 B.n82 585
R275 B.n124 B.n123 585
R276 B.n122 B.n83 585
R277 B.n121 B.n120 585
R278 B.n119 B.n84 585
R279 B.n118 B.n117 585
R280 B.n116 B.n85 585
R281 B.n115 B.n114 585
R282 B.n113 B.n86 585
R283 B.n112 B.n111 585
R284 B.n110 B.n87 585
R285 B.n109 B.n108 585
R286 B.n107 B.n88 585
R287 B.n106 B.n105 585
R288 B.n104 B.n89 585
R289 B.n103 B.n102 585
R290 B.n101 B.n90 585
R291 B.n100 B.n99 585
R292 B.n98 B.n91 585
R293 B.n97 B.n96 585
R294 B.n95 B.n92 585
R295 B.n94 B.n93 585
R296 B.n2 B.n0 585
R297 B.n341 B.n1 585
R298 B.n340 B.n339 585
R299 B.n338 B.n3 585
R300 B.n337 B.n336 585
R301 B.n335 B.n4 585
R302 B.n334 B.n333 585
R303 B.n332 B.n5 585
R304 B.n331 B.n330 585
R305 B.n329 B.n6 585
R306 B.n328 B.n327 585
R307 B.n326 B.n7 585
R308 B.n325 B.n324 585
R309 B.n323 B.n8 585
R310 B.n322 B.n321 585
R311 B.n320 B.n9 585
R312 B.n319 B.n318 585
R313 B.n317 B.n10 585
R314 B.n316 B.n315 585
R315 B.n314 B.n11 585
R316 B.n313 B.n312 585
R317 B.n311 B.n12 585
R318 B.n310 B.n309 585
R319 B.n308 B.n13 585
R320 B.n343 B.n342 585
R321 B.n126 B.n125 545.355
R322 B.n306 B.n13 545.355
R323 B.n180 B.n59 545.355
R324 B.n252 B.n251 545.355
R325 B.n66 B.t2 271.767
R326 B.n28 B.t7 271.767
R327 B.n74 B.t11 271.767
R328 B.n20 B.t4 271.767
R329 B.n66 B.t0 233.446
R330 B.n74 B.t9 233.446
R331 B.n20 B.t3 233.446
R332 B.n28 B.t6 233.446
R333 B.n67 B.t1 222.311
R334 B.n29 B.t8 222.311
R335 B.n75 B.t10 222.311
R336 B.n21 B.t5 222.311
R337 B.n125 B.n124 163.367
R338 B.n124 B.n83 163.367
R339 B.n120 B.n83 163.367
R340 B.n120 B.n119 163.367
R341 B.n119 B.n118 163.367
R342 B.n118 B.n85 163.367
R343 B.n114 B.n85 163.367
R344 B.n114 B.n113 163.367
R345 B.n113 B.n112 163.367
R346 B.n112 B.n87 163.367
R347 B.n108 B.n87 163.367
R348 B.n108 B.n107 163.367
R349 B.n107 B.n106 163.367
R350 B.n106 B.n89 163.367
R351 B.n102 B.n89 163.367
R352 B.n102 B.n101 163.367
R353 B.n101 B.n100 163.367
R354 B.n100 B.n91 163.367
R355 B.n96 B.n91 163.367
R356 B.n96 B.n95 163.367
R357 B.n95 B.n94 163.367
R358 B.n94 B.n2 163.367
R359 B.n342 B.n2 163.367
R360 B.n342 B.n341 163.367
R361 B.n341 B.n340 163.367
R362 B.n340 B.n3 163.367
R363 B.n336 B.n3 163.367
R364 B.n336 B.n335 163.367
R365 B.n335 B.n334 163.367
R366 B.n334 B.n5 163.367
R367 B.n330 B.n5 163.367
R368 B.n330 B.n329 163.367
R369 B.n329 B.n328 163.367
R370 B.n328 B.n7 163.367
R371 B.n324 B.n7 163.367
R372 B.n324 B.n323 163.367
R373 B.n323 B.n322 163.367
R374 B.n322 B.n9 163.367
R375 B.n318 B.n9 163.367
R376 B.n318 B.n317 163.367
R377 B.n317 B.n316 163.367
R378 B.n316 B.n11 163.367
R379 B.n312 B.n11 163.367
R380 B.n312 B.n311 163.367
R381 B.n311 B.n310 163.367
R382 B.n310 B.n13 163.367
R383 B.n126 B.n81 163.367
R384 B.n130 B.n81 163.367
R385 B.n131 B.n130 163.367
R386 B.n132 B.n131 163.367
R387 B.n132 B.n79 163.367
R388 B.n136 B.n79 163.367
R389 B.n137 B.n136 163.367
R390 B.n138 B.n137 163.367
R391 B.n138 B.n77 163.367
R392 B.n142 B.n77 163.367
R393 B.n143 B.n142 163.367
R394 B.n144 B.n143 163.367
R395 B.n144 B.n73 163.367
R396 B.n149 B.n73 163.367
R397 B.n150 B.n149 163.367
R398 B.n151 B.n150 163.367
R399 B.n151 B.n71 163.367
R400 B.n155 B.n71 163.367
R401 B.n156 B.n155 163.367
R402 B.n157 B.n156 163.367
R403 B.n157 B.n69 163.367
R404 B.n161 B.n69 163.367
R405 B.n162 B.n161 163.367
R406 B.n162 B.n65 163.367
R407 B.n166 B.n65 163.367
R408 B.n167 B.n166 163.367
R409 B.n168 B.n167 163.367
R410 B.n168 B.n63 163.367
R411 B.n172 B.n63 163.367
R412 B.n173 B.n172 163.367
R413 B.n174 B.n173 163.367
R414 B.n174 B.n61 163.367
R415 B.n178 B.n61 163.367
R416 B.n179 B.n178 163.367
R417 B.n180 B.n179 163.367
R418 B.n184 B.n59 163.367
R419 B.n185 B.n184 163.367
R420 B.n186 B.n185 163.367
R421 B.n186 B.n57 163.367
R422 B.n190 B.n57 163.367
R423 B.n191 B.n190 163.367
R424 B.n192 B.n191 163.367
R425 B.n192 B.n55 163.367
R426 B.n196 B.n55 163.367
R427 B.n197 B.n196 163.367
R428 B.n198 B.n197 163.367
R429 B.n198 B.n53 163.367
R430 B.n202 B.n53 163.367
R431 B.n203 B.n202 163.367
R432 B.n204 B.n203 163.367
R433 B.n204 B.n51 163.367
R434 B.n208 B.n51 163.367
R435 B.n209 B.n208 163.367
R436 B.n210 B.n209 163.367
R437 B.n210 B.n49 163.367
R438 B.n214 B.n49 163.367
R439 B.n215 B.n214 163.367
R440 B.n216 B.n215 163.367
R441 B.n216 B.n47 163.367
R442 B.n220 B.n47 163.367
R443 B.n221 B.n220 163.367
R444 B.n222 B.n221 163.367
R445 B.n222 B.n45 163.367
R446 B.n226 B.n45 163.367
R447 B.n227 B.n226 163.367
R448 B.n228 B.n227 163.367
R449 B.n228 B.n43 163.367
R450 B.n232 B.n43 163.367
R451 B.n233 B.n232 163.367
R452 B.n234 B.n233 163.367
R453 B.n234 B.n41 163.367
R454 B.n238 B.n41 163.367
R455 B.n239 B.n238 163.367
R456 B.n240 B.n239 163.367
R457 B.n240 B.n39 163.367
R458 B.n244 B.n39 163.367
R459 B.n245 B.n244 163.367
R460 B.n246 B.n245 163.367
R461 B.n246 B.n37 163.367
R462 B.n250 B.n37 163.367
R463 B.n251 B.n250 163.367
R464 B.n306 B.n305 163.367
R465 B.n305 B.n304 163.367
R466 B.n304 B.n15 163.367
R467 B.n300 B.n15 163.367
R468 B.n300 B.n299 163.367
R469 B.n299 B.n298 163.367
R470 B.n298 B.n17 163.367
R471 B.n294 B.n17 163.367
R472 B.n294 B.n293 163.367
R473 B.n293 B.n292 163.367
R474 B.n292 B.n19 163.367
R475 B.n288 B.n19 163.367
R476 B.n288 B.n287 163.367
R477 B.n287 B.n23 163.367
R478 B.n283 B.n23 163.367
R479 B.n283 B.n282 163.367
R480 B.n282 B.n281 163.367
R481 B.n281 B.n25 163.367
R482 B.n277 B.n25 163.367
R483 B.n277 B.n276 163.367
R484 B.n276 B.n275 163.367
R485 B.n275 B.n27 163.367
R486 B.n270 B.n27 163.367
R487 B.n270 B.n269 163.367
R488 B.n269 B.n268 163.367
R489 B.n268 B.n31 163.367
R490 B.n264 B.n31 163.367
R491 B.n264 B.n263 163.367
R492 B.n263 B.n262 163.367
R493 B.n262 B.n33 163.367
R494 B.n258 B.n33 163.367
R495 B.n258 B.n257 163.367
R496 B.n257 B.n256 163.367
R497 B.n256 B.n35 163.367
R498 B.n252 B.n35 163.367
R499 B.n68 B.n67 59.5399
R500 B.n146 B.n75 59.5399
R501 B.n22 B.n21 59.5399
R502 B.n272 B.n29 59.5399
R503 B.n67 B.n66 49.455
R504 B.n75 B.n74 49.455
R505 B.n21 B.n20 49.455
R506 B.n29 B.n28 49.455
R507 B.n308 B.n307 35.4346
R508 B.n182 B.n181 35.4346
R509 B.n127 B.n82 35.4346
R510 B.n253 B.n36 35.4346
R511 B B.n343 18.0485
R512 B.n307 B.n14 10.6151
R513 B.n303 B.n14 10.6151
R514 B.n303 B.n302 10.6151
R515 B.n302 B.n301 10.6151
R516 B.n301 B.n16 10.6151
R517 B.n297 B.n16 10.6151
R518 B.n297 B.n296 10.6151
R519 B.n296 B.n295 10.6151
R520 B.n295 B.n18 10.6151
R521 B.n291 B.n18 10.6151
R522 B.n291 B.n290 10.6151
R523 B.n290 B.n289 10.6151
R524 B.n286 B.n285 10.6151
R525 B.n285 B.n284 10.6151
R526 B.n284 B.n24 10.6151
R527 B.n280 B.n24 10.6151
R528 B.n280 B.n279 10.6151
R529 B.n279 B.n278 10.6151
R530 B.n278 B.n26 10.6151
R531 B.n274 B.n26 10.6151
R532 B.n274 B.n273 10.6151
R533 B.n271 B.n30 10.6151
R534 B.n267 B.n30 10.6151
R535 B.n267 B.n266 10.6151
R536 B.n266 B.n265 10.6151
R537 B.n265 B.n32 10.6151
R538 B.n261 B.n32 10.6151
R539 B.n261 B.n260 10.6151
R540 B.n260 B.n259 10.6151
R541 B.n259 B.n34 10.6151
R542 B.n255 B.n34 10.6151
R543 B.n255 B.n254 10.6151
R544 B.n254 B.n253 10.6151
R545 B.n183 B.n182 10.6151
R546 B.n183 B.n58 10.6151
R547 B.n187 B.n58 10.6151
R548 B.n188 B.n187 10.6151
R549 B.n189 B.n188 10.6151
R550 B.n189 B.n56 10.6151
R551 B.n193 B.n56 10.6151
R552 B.n194 B.n193 10.6151
R553 B.n195 B.n194 10.6151
R554 B.n195 B.n54 10.6151
R555 B.n199 B.n54 10.6151
R556 B.n200 B.n199 10.6151
R557 B.n201 B.n200 10.6151
R558 B.n201 B.n52 10.6151
R559 B.n205 B.n52 10.6151
R560 B.n206 B.n205 10.6151
R561 B.n207 B.n206 10.6151
R562 B.n207 B.n50 10.6151
R563 B.n211 B.n50 10.6151
R564 B.n212 B.n211 10.6151
R565 B.n213 B.n212 10.6151
R566 B.n213 B.n48 10.6151
R567 B.n217 B.n48 10.6151
R568 B.n218 B.n217 10.6151
R569 B.n219 B.n218 10.6151
R570 B.n219 B.n46 10.6151
R571 B.n223 B.n46 10.6151
R572 B.n224 B.n223 10.6151
R573 B.n225 B.n224 10.6151
R574 B.n225 B.n44 10.6151
R575 B.n229 B.n44 10.6151
R576 B.n230 B.n229 10.6151
R577 B.n231 B.n230 10.6151
R578 B.n231 B.n42 10.6151
R579 B.n235 B.n42 10.6151
R580 B.n236 B.n235 10.6151
R581 B.n237 B.n236 10.6151
R582 B.n237 B.n40 10.6151
R583 B.n241 B.n40 10.6151
R584 B.n242 B.n241 10.6151
R585 B.n243 B.n242 10.6151
R586 B.n243 B.n38 10.6151
R587 B.n247 B.n38 10.6151
R588 B.n248 B.n247 10.6151
R589 B.n249 B.n248 10.6151
R590 B.n249 B.n36 10.6151
R591 B.n128 B.n127 10.6151
R592 B.n129 B.n128 10.6151
R593 B.n129 B.n80 10.6151
R594 B.n133 B.n80 10.6151
R595 B.n134 B.n133 10.6151
R596 B.n135 B.n134 10.6151
R597 B.n135 B.n78 10.6151
R598 B.n139 B.n78 10.6151
R599 B.n140 B.n139 10.6151
R600 B.n141 B.n140 10.6151
R601 B.n141 B.n76 10.6151
R602 B.n145 B.n76 10.6151
R603 B.n148 B.n147 10.6151
R604 B.n148 B.n72 10.6151
R605 B.n152 B.n72 10.6151
R606 B.n153 B.n152 10.6151
R607 B.n154 B.n153 10.6151
R608 B.n154 B.n70 10.6151
R609 B.n158 B.n70 10.6151
R610 B.n159 B.n158 10.6151
R611 B.n160 B.n159 10.6151
R612 B.n164 B.n163 10.6151
R613 B.n165 B.n164 10.6151
R614 B.n165 B.n64 10.6151
R615 B.n169 B.n64 10.6151
R616 B.n170 B.n169 10.6151
R617 B.n171 B.n170 10.6151
R618 B.n171 B.n62 10.6151
R619 B.n175 B.n62 10.6151
R620 B.n176 B.n175 10.6151
R621 B.n177 B.n176 10.6151
R622 B.n177 B.n60 10.6151
R623 B.n181 B.n60 10.6151
R624 B.n123 B.n82 10.6151
R625 B.n123 B.n122 10.6151
R626 B.n122 B.n121 10.6151
R627 B.n121 B.n84 10.6151
R628 B.n117 B.n84 10.6151
R629 B.n117 B.n116 10.6151
R630 B.n116 B.n115 10.6151
R631 B.n115 B.n86 10.6151
R632 B.n111 B.n86 10.6151
R633 B.n111 B.n110 10.6151
R634 B.n110 B.n109 10.6151
R635 B.n109 B.n88 10.6151
R636 B.n105 B.n88 10.6151
R637 B.n105 B.n104 10.6151
R638 B.n104 B.n103 10.6151
R639 B.n103 B.n90 10.6151
R640 B.n99 B.n90 10.6151
R641 B.n99 B.n98 10.6151
R642 B.n98 B.n97 10.6151
R643 B.n97 B.n92 10.6151
R644 B.n93 B.n92 10.6151
R645 B.n93 B.n0 10.6151
R646 B.n339 B.n1 10.6151
R647 B.n339 B.n338 10.6151
R648 B.n338 B.n337 10.6151
R649 B.n337 B.n4 10.6151
R650 B.n333 B.n4 10.6151
R651 B.n333 B.n332 10.6151
R652 B.n332 B.n331 10.6151
R653 B.n331 B.n6 10.6151
R654 B.n327 B.n6 10.6151
R655 B.n327 B.n326 10.6151
R656 B.n326 B.n325 10.6151
R657 B.n325 B.n8 10.6151
R658 B.n321 B.n8 10.6151
R659 B.n321 B.n320 10.6151
R660 B.n320 B.n319 10.6151
R661 B.n319 B.n10 10.6151
R662 B.n315 B.n10 10.6151
R663 B.n315 B.n314 10.6151
R664 B.n314 B.n313 10.6151
R665 B.n313 B.n12 10.6151
R666 B.n309 B.n12 10.6151
R667 B.n309 B.n308 10.6151
R668 B.n289 B.n22 9.36635
R669 B.n272 B.n271 9.36635
R670 B.n146 B.n145 9.36635
R671 B.n163 B.n68 9.36635
R672 B.n343 B.n0 2.81026
R673 B.n343 B.n1 2.81026
R674 B.n286 B.n22 1.24928
R675 B.n273 B.n272 1.24928
R676 B.n147 B.n146 1.24928
R677 B.n160 B.n68 1.24928
C0 VDD2 VTAIL 2.46338f
C1 VDD1 w_n1990_n1448# 1.06157f
C2 VN VTAIL 0.946183f
C3 VDD1 VP 0.911322f
C4 B w_n1990_n1448# 5.72273f
C5 B VP 1.26522f
C6 VN VDD2 0.743923f
C7 B VDD1 0.901951f
C8 w_n1990_n1448# VTAIL 1.34485f
C9 VTAIL VP 0.960333f
C10 VDD1 VTAIL 2.41319f
C11 VDD2 w_n1990_n1448# 1.08221f
C12 B VTAIL 1.33788f
C13 VDD2 VP 0.323008f
C14 VN w_n1990_n1448# 2.51932f
C15 VDD2 VDD1 0.627957f
C16 VN VP 3.50618f
C17 VN VDD1 0.154052f
C18 B VDD2 0.928929f
C19 VN B 0.851953f
C20 w_n1990_n1448# VP 2.76856f
C21 VDD2 VSUBS 0.527332f
C22 VDD1 VSUBS 2.045151f
C23 VTAIL VSUBS 0.368238f
C24 VN VSUBS 5.16215f
C25 VP VSUBS 1.118931f
C26 B VSUBS 2.669661f
C27 w_n1990_n1448# VSUBS 36.6558f
C28 B.n0 VSUBS 0.005482f
C29 B.n1 VSUBS 0.005482f
C30 B.n2 VSUBS 0.008669f
C31 B.n3 VSUBS 0.008669f
C32 B.n4 VSUBS 0.008669f
C33 B.n5 VSUBS 0.008669f
C34 B.n6 VSUBS 0.008669f
C35 B.n7 VSUBS 0.008669f
C36 B.n8 VSUBS 0.008669f
C37 B.n9 VSUBS 0.008669f
C38 B.n10 VSUBS 0.008669f
C39 B.n11 VSUBS 0.008669f
C40 B.n12 VSUBS 0.008669f
C41 B.n13 VSUBS 0.021016f
C42 B.n14 VSUBS 0.008669f
C43 B.n15 VSUBS 0.008669f
C44 B.n16 VSUBS 0.008669f
C45 B.n17 VSUBS 0.008669f
C46 B.n18 VSUBS 0.008669f
C47 B.n19 VSUBS 0.008669f
C48 B.t5 VSUBS 0.045917f
C49 B.t4 VSUBS 0.061048f
C50 B.t3 VSUBS 0.322118f
C51 B.n20 VSUBS 0.110197f
C52 B.n21 VSUBS 0.095516f
C53 B.n22 VSUBS 0.020086f
C54 B.n23 VSUBS 0.008669f
C55 B.n24 VSUBS 0.008669f
C56 B.n25 VSUBS 0.008669f
C57 B.n26 VSUBS 0.008669f
C58 B.n27 VSUBS 0.008669f
C59 B.t8 VSUBS 0.045917f
C60 B.t7 VSUBS 0.061048f
C61 B.t6 VSUBS 0.322118f
C62 B.n28 VSUBS 0.110197f
C63 B.n29 VSUBS 0.095516f
C64 B.n30 VSUBS 0.008669f
C65 B.n31 VSUBS 0.008669f
C66 B.n32 VSUBS 0.008669f
C67 B.n33 VSUBS 0.008669f
C68 B.n34 VSUBS 0.008669f
C69 B.n35 VSUBS 0.008669f
C70 B.n36 VSUBS 0.02196f
C71 B.n37 VSUBS 0.008669f
C72 B.n38 VSUBS 0.008669f
C73 B.n39 VSUBS 0.008669f
C74 B.n40 VSUBS 0.008669f
C75 B.n41 VSUBS 0.008669f
C76 B.n42 VSUBS 0.008669f
C77 B.n43 VSUBS 0.008669f
C78 B.n44 VSUBS 0.008669f
C79 B.n45 VSUBS 0.008669f
C80 B.n46 VSUBS 0.008669f
C81 B.n47 VSUBS 0.008669f
C82 B.n48 VSUBS 0.008669f
C83 B.n49 VSUBS 0.008669f
C84 B.n50 VSUBS 0.008669f
C85 B.n51 VSUBS 0.008669f
C86 B.n52 VSUBS 0.008669f
C87 B.n53 VSUBS 0.008669f
C88 B.n54 VSUBS 0.008669f
C89 B.n55 VSUBS 0.008669f
C90 B.n56 VSUBS 0.008669f
C91 B.n57 VSUBS 0.008669f
C92 B.n58 VSUBS 0.008669f
C93 B.n59 VSUBS 0.021016f
C94 B.n60 VSUBS 0.008669f
C95 B.n61 VSUBS 0.008669f
C96 B.n62 VSUBS 0.008669f
C97 B.n63 VSUBS 0.008669f
C98 B.n64 VSUBS 0.008669f
C99 B.n65 VSUBS 0.008669f
C100 B.t1 VSUBS 0.045917f
C101 B.t2 VSUBS 0.061048f
C102 B.t0 VSUBS 0.322118f
C103 B.n66 VSUBS 0.110197f
C104 B.n67 VSUBS 0.095516f
C105 B.n68 VSUBS 0.020086f
C106 B.n69 VSUBS 0.008669f
C107 B.n70 VSUBS 0.008669f
C108 B.n71 VSUBS 0.008669f
C109 B.n72 VSUBS 0.008669f
C110 B.n73 VSUBS 0.008669f
C111 B.t10 VSUBS 0.045917f
C112 B.t11 VSUBS 0.061048f
C113 B.t9 VSUBS 0.322118f
C114 B.n74 VSUBS 0.110197f
C115 B.n75 VSUBS 0.095516f
C116 B.n76 VSUBS 0.008669f
C117 B.n77 VSUBS 0.008669f
C118 B.n78 VSUBS 0.008669f
C119 B.n79 VSUBS 0.008669f
C120 B.n80 VSUBS 0.008669f
C121 B.n81 VSUBS 0.008669f
C122 B.n82 VSUBS 0.021016f
C123 B.n83 VSUBS 0.008669f
C124 B.n84 VSUBS 0.008669f
C125 B.n85 VSUBS 0.008669f
C126 B.n86 VSUBS 0.008669f
C127 B.n87 VSUBS 0.008669f
C128 B.n88 VSUBS 0.008669f
C129 B.n89 VSUBS 0.008669f
C130 B.n90 VSUBS 0.008669f
C131 B.n91 VSUBS 0.008669f
C132 B.n92 VSUBS 0.008669f
C133 B.n93 VSUBS 0.008669f
C134 B.n94 VSUBS 0.008669f
C135 B.n95 VSUBS 0.008669f
C136 B.n96 VSUBS 0.008669f
C137 B.n97 VSUBS 0.008669f
C138 B.n98 VSUBS 0.008669f
C139 B.n99 VSUBS 0.008669f
C140 B.n100 VSUBS 0.008669f
C141 B.n101 VSUBS 0.008669f
C142 B.n102 VSUBS 0.008669f
C143 B.n103 VSUBS 0.008669f
C144 B.n104 VSUBS 0.008669f
C145 B.n105 VSUBS 0.008669f
C146 B.n106 VSUBS 0.008669f
C147 B.n107 VSUBS 0.008669f
C148 B.n108 VSUBS 0.008669f
C149 B.n109 VSUBS 0.008669f
C150 B.n110 VSUBS 0.008669f
C151 B.n111 VSUBS 0.008669f
C152 B.n112 VSUBS 0.008669f
C153 B.n113 VSUBS 0.008669f
C154 B.n114 VSUBS 0.008669f
C155 B.n115 VSUBS 0.008669f
C156 B.n116 VSUBS 0.008669f
C157 B.n117 VSUBS 0.008669f
C158 B.n118 VSUBS 0.008669f
C159 B.n119 VSUBS 0.008669f
C160 B.n120 VSUBS 0.008669f
C161 B.n121 VSUBS 0.008669f
C162 B.n122 VSUBS 0.008669f
C163 B.n123 VSUBS 0.008669f
C164 B.n124 VSUBS 0.008669f
C165 B.n125 VSUBS 0.021016f
C166 B.n126 VSUBS 0.021822f
C167 B.n127 VSUBS 0.021822f
C168 B.n128 VSUBS 0.008669f
C169 B.n129 VSUBS 0.008669f
C170 B.n130 VSUBS 0.008669f
C171 B.n131 VSUBS 0.008669f
C172 B.n132 VSUBS 0.008669f
C173 B.n133 VSUBS 0.008669f
C174 B.n134 VSUBS 0.008669f
C175 B.n135 VSUBS 0.008669f
C176 B.n136 VSUBS 0.008669f
C177 B.n137 VSUBS 0.008669f
C178 B.n138 VSUBS 0.008669f
C179 B.n139 VSUBS 0.008669f
C180 B.n140 VSUBS 0.008669f
C181 B.n141 VSUBS 0.008669f
C182 B.n142 VSUBS 0.008669f
C183 B.n143 VSUBS 0.008669f
C184 B.n144 VSUBS 0.008669f
C185 B.n145 VSUBS 0.00816f
C186 B.n146 VSUBS 0.020086f
C187 B.n147 VSUBS 0.004845f
C188 B.n148 VSUBS 0.008669f
C189 B.n149 VSUBS 0.008669f
C190 B.n150 VSUBS 0.008669f
C191 B.n151 VSUBS 0.008669f
C192 B.n152 VSUBS 0.008669f
C193 B.n153 VSUBS 0.008669f
C194 B.n154 VSUBS 0.008669f
C195 B.n155 VSUBS 0.008669f
C196 B.n156 VSUBS 0.008669f
C197 B.n157 VSUBS 0.008669f
C198 B.n158 VSUBS 0.008669f
C199 B.n159 VSUBS 0.008669f
C200 B.n160 VSUBS 0.004845f
C201 B.n161 VSUBS 0.008669f
C202 B.n162 VSUBS 0.008669f
C203 B.n163 VSUBS 0.00816f
C204 B.n164 VSUBS 0.008669f
C205 B.n165 VSUBS 0.008669f
C206 B.n166 VSUBS 0.008669f
C207 B.n167 VSUBS 0.008669f
C208 B.n168 VSUBS 0.008669f
C209 B.n169 VSUBS 0.008669f
C210 B.n170 VSUBS 0.008669f
C211 B.n171 VSUBS 0.008669f
C212 B.n172 VSUBS 0.008669f
C213 B.n173 VSUBS 0.008669f
C214 B.n174 VSUBS 0.008669f
C215 B.n175 VSUBS 0.008669f
C216 B.n176 VSUBS 0.008669f
C217 B.n177 VSUBS 0.008669f
C218 B.n178 VSUBS 0.008669f
C219 B.n179 VSUBS 0.008669f
C220 B.n180 VSUBS 0.021822f
C221 B.n181 VSUBS 0.021822f
C222 B.n182 VSUBS 0.021016f
C223 B.n183 VSUBS 0.008669f
C224 B.n184 VSUBS 0.008669f
C225 B.n185 VSUBS 0.008669f
C226 B.n186 VSUBS 0.008669f
C227 B.n187 VSUBS 0.008669f
C228 B.n188 VSUBS 0.008669f
C229 B.n189 VSUBS 0.008669f
C230 B.n190 VSUBS 0.008669f
C231 B.n191 VSUBS 0.008669f
C232 B.n192 VSUBS 0.008669f
C233 B.n193 VSUBS 0.008669f
C234 B.n194 VSUBS 0.008669f
C235 B.n195 VSUBS 0.008669f
C236 B.n196 VSUBS 0.008669f
C237 B.n197 VSUBS 0.008669f
C238 B.n198 VSUBS 0.008669f
C239 B.n199 VSUBS 0.008669f
C240 B.n200 VSUBS 0.008669f
C241 B.n201 VSUBS 0.008669f
C242 B.n202 VSUBS 0.008669f
C243 B.n203 VSUBS 0.008669f
C244 B.n204 VSUBS 0.008669f
C245 B.n205 VSUBS 0.008669f
C246 B.n206 VSUBS 0.008669f
C247 B.n207 VSUBS 0.008669f
C248 B.n208 VSUBS 0.008669f
C249 B.n209 VSUBS 0.008669f
C250 B.n210 VSUBS 0.008669f
C251 B.n211 VSUBS 0.008669f
C252 B.n212 VSUBS 0.008669f
C253 B.n213 VSUBS 0.008669f
C254 B.n214 VSUBS 0.008669f
C255 B.n215 VSUBS 0.008669f
C256 B.n216 VSUBS 0.008669f
C257 B.n217 VSUBS 0.008669f
C258 B.n218 VSUBS 0.008669f
C259 B.n219 VSUBS 0.008669f
C260 B.n220 VSUBS 0.008669f
C261 B.n221 VSUBS 0.008669f
C262 B.n222 VSUBS 0.008669f
C263 B.n223 VSUBS 0.008669f
C264 B.n224 VSUBS 0.008669f
C265 B.n225 VSUBS 0.008669f
C266 B.n226 VSUBS 0.008669f
C267 B.n227 VSUBS 0.008669f
C268 B.n228 VSUBS 0.008669f
C269 B.n229 VSUBS 0.008669f
C270 B.n230 VSUBS 0.008669f
C271 B.n231 VSUBS 0.008669f
C272 B.n232 VSUBS 0.008669f
C273 B.n233 VSUBS 0.008669f
C274 B.n234 VSUBS 0.008669f
C275 B.n235 VSUBS 0.008669f
C276 B.n236 VSUBS 0.008669f
C277 B.n237 VSUBS 0.008669f
C278 B.n238 VSUBS 0.008669f
C279 B.n239 VSUBS 0.008669f
C280 B.n240 VSUBS 0.008669f
C281 B.n241 VSUBS 0.008669f
C282 B.n242 VSUBS 0.008669f
C283 B.n243 VSUBS 0.008669f
C284 B.n244 VSUBS 0.008669f
C285 B.n245 VSUBS 0.008669f
C286 B.n246 VSUBS 0.008669f
C287 B.n247 VSUBS 0.008669f
C288 B.n248 VSUBS 0.008669f
C289 B.n249 VSUBS 0.008669f
C290 B.n250 VSUBS 0.008669f
C291 B.n251 VSUBS 0.021016f
C292 B.n252 VSUBS 0.021822f
C293 B.n253 VSUBS 0.020878f
C294 B.n254 VSUBS 0.008669f
C295 B.n255 VSUBS 0.008669f
C296 B.n256 VSUBS 0.008669f
C297 B.n257 VSUBS 0.008669f
C298 B.n258 VSUBS 0.008669f
C299 B.n259 VSUBS 0.008669f
C300 B.n260 VSUBS 0.008669f
C301 B.n261 VSUBS 0.008669f
C302 B.n262 VSUBS 0.008669f
C303 B.n263 VSUBS 0.008669f
C304 B.n264 VSUBS 0.008669f
C305 B.n265 VSUBS 0.008669f
C306 B.n266 VSUBS 0.008669f
C307 B.n267 VSUBS 0.008669f
C308 B.n268 VSUBS 0.008669f
C309 B.n269 VSUBS 0.008669f
C310 B.n270 VSUBS 0.008669f
C311 B.n271 VSUBS 0.00816f
C312 B.n272 VSUBS 0.020086f
C313 B.n273 VSUBS 0.004845f
C314 B.n274 VSUBS 0.008669f
C315 B.n275 VSUBS 0.008669f
C316 B.n276 VSUBS 0.008669f
C317 B.n277 VSUBS 0.008669f
C318 B.n278 VSUBS 0.008669f
C319 B.n279 VSUBS 0.008669f
C320 B.n280 VSUBS 0.008669f
C321 B.n281 VSUBS 0.008669f
C322 B.n282 VSUBS 0.008669f
C323 B.n283 VSUBS 0.008669f
C324 B.n284 VSUBS 0.008669f
C325 B.n285 VSUBS 0.008669f
C326 B.n286 VSUBS 0.004845f
C327 B.n287 VSUBS 0.008669f
C328 B.n288 VSUBS 0.008669f
C329 B.n289 VSUBS 0.00816f
C330 B.n290 VSUBS 0.008669f
C331 B.n291 VSUBS 0.008669f
C332 B.n292 VSUBS 0.008669f
C333 B.n293 VSUBS 0.008669f
C334 B.n294 VSUBS 0.008669f
C335 B.n295 VSUBS 0.008669f
C336 B.n296 VSUBS 0.008669f
C337 B.n297 VSUBS 0.008669f
C338 B.n298 VSUBS 0.008669f
C339 B.n299 VSUBS 0.008669f
C340 B.n300 VSUBS 0.008669f
C341 B.n301 VSUBS 0.008669f
C342 B.n302 VSUBS 0.008669f
C343 B.n303 VSUBS 0.008669f
C344 B.n304 VSUBS 0.008669f
C345 B.n305 VSUBS 0.008669f
C346 B.n306 VSUBS 0.021822f
C347 B.n307 VSUBS 0.021822f
C348 B.n308 VSUBS 0.021016f
C349 B.n309 VSUBS 0.008669f
C350 B.n310 VSUBS 0.008669f
C351 B.n311 VSUBS 0.008669f
C352 B.n312 VSUBS 0.008669f
C353 B.n313 VSUBS 0.008669f
C354 B.n314 VSUBS 0.008669f
C355 B.n315 VSUBS 0.008669f
C356 B.n316 VSUBS 0.008669f
C357 B.n317 VSUBS 0.008669f
C358 B.n318 VSUBS 0.008669f
C359 B.n319 VSUBS 0.008669f
C360 B.n320 VSUBS 0.008669f
C361 B.n321 VSUBS 0.008669f
C362 B.n322 VSUBS 0.008669f
C363 B.n323 VSUBS 0.008669f
C364 B.n324 VSUBS 0.008669f
C365 B.n325 VSUBS 0.008669f
C366 B.n326 VSUBS 0.008669f
C367 B.n327 VSUBS 0.008669f
C368 B.n328 VSUBS 0.008669f
C369 B.n329 VSUBS 0.008669f
C370 B.n330 VSUBS 0.008669f
C371 B.n331 VSUBS 0.008669f
C372 B.n332 VSUBS 0.008669f
C373 B.n333 VSUBS 0.008669f
C374 B.n334 VSUBS 0.008669f
C375 B.n335 VSUBS 0.008669f
C376 B.n336 VSUBS 0.008669f
C377 B.n337 VSUBS 0.008669f
C378 B.n338 VSUBS 0.008669f
C379 B.n339 VSUBS 0.008669f
C380 B.n340 VSUBS 0.008669f
C381 B.n341 VSUBS 0.008669f
C382 B.n342 VSUBS 0.008669f
C383 B.n343 VSUBS 0.019631f
C384 VDD1.n0 VSUBS 0.01619f
C385 VDD1.n1 VSUBS 0.108265f
C386 VDD1.n2 VSUBS 0.008615f
C387 VDD1.t0 VSUBS 0.044218f
C388 VDD1.n3 VSUBS 0.051627f
C389 VDD1.n4 VSUBS 0.012007f
C390 VDD1.n5 VSUBS 0.015272f
C391 VDD1.n6 VSUBS 0.044439f
C392 VDD1.n7 VSUBS 0.009122f
C393 VDD1.n8 VSUBS 0.008615f
C394 VDD1.n9 VSUBS 0.037058f
C395 VDD1.n10 VSUBS 0.033967f
C396 VDD1.n11 VSUBS 0.01619f
C397 VDD1.n12 VSUBS 0.108265f
C398 VDD1.n13 VSUBS 0.008615f
C399 VDD1.t1 VSUBS 0.044218f
C400 VDD1.n14 VSUBS 0.051627f
C401 VDD1.n15 VSUBS 0.012007f
C402 VDD1.n16 VSUBS 0.015272f
C403 VDD1.n17 VSUBS 0.044439f
C404 VDD1.n18 VSUBS 0.009122f
C405 VDD1.n19 VSUBS 0.008615f
C406 VDD1.n20 VSUBS 0.037058f
C407 VDD1.n21 VSUBS 0.282942f
C408 VP.t1 VSUBS 1.73559f
C409 VP.t0 VSUBS 1.06441f
C410 VP.n0 VSUBS 3.39412f
C411 VDD2.n0 VSUBS 0.017291f
C412 VDD2.n1 VSUBS 0.115629f
C413 VDD2.n2 VSUBS 0.009201f
C414 VDD2.t1 VSUBS 0.047225f
C415 VDD2.n3 VSUBS 0.055138f
C416 VDD2.n4 VSUBS 0.012823f
C417 VDD2.n5 VSUBS 0.016311f
C418 VDD2.n6 VSUBS 0.047461f
C419 VDD2.n7 VSUBS 0.009742f
C420 VDD2.n8 VSUBS 0.009201f
C421 VDD2.n9 VSUBS 0.039579f
C422 VDD2.n10 VSUBS 0.276981f
C423 VDD2.n11 VSUBS 0.017291f
C424 VDD2.n12 VSUBS 0.115629f
C425 VDD2.n13 VSUBS 0.009201f
C426 VDD2.t0 VSUBS 0.047225f
C427 VDD2.n14 VSUBS 0.055138f
C428 VDD2.n15 VSUBS 0.012823f
C429 VDD2.n16 VSUBS 0.016311f
C430 VDD2.n17 VSUBS 0.047461f
C431 VDD2.n18 VSUBS 0.009742f
C432 VDD2.n19 VSUBS 0.009201f
C433 VDD2.n20 VSUBS 0.039579f
C434 VDD2.n21 VSUBS 0.03546f
C435 VDD2.n22 VSUBS 1.3337f
C436 VTAIL.n0 VSUBS 0.020503f
C437 VTAIL.n1 VSUBS 0.137105f
C438 VTAIL.n2 VSUBS 0.01091f
C439 VTAIL.t1 VSUBS 0.055997f
C440 VTAIL.n3 VSUBS 0.06538f
C441 VTAIL.n4 VSUBS 0.015205f
C442 VTAIL.n5 VSUBS 0.019341f
C443 VTAIL.n6 VSUBS 0.056277f
C444 VTAIL.n7 VSUBS 0.011552f
C445 VTAIL.n8 VSUBS 0.01091f
C446 VTAIL.n9 VSUBS 0.04693f
C447 VTAIL.n10 VSUBS 0.028028f
C448 VTAIL.n11 VSUBS 0.786623f
C449 VTAIL.n12 VSUBS 0.020503f
C450 VTAIL.n13 VSUBS 0.137105f
C451 VTAIL.n14 VSUBS 0.01091f
C452 VTAIL.t2 VSUBS 0.055997f
C453 VTAIL.n15 VSUBS 0.06538f
C454 VTAIL.n16 VSUBS 0.015205f
C455 VTAIL.n17 VSUBS 0.019341f
C456 VTAIL.n18 VSUBS 0.056277f
C457 VTAIL.n19 VSUBS 0.011552f
C458 VTAIL.n20 VSUBS 0.01091f
C459 VTAIL.n21 VSUBS 0.04693f
C460 VTAIL.n22 VSUBS 0.028028f
C461 VTAIL.n23 VSUBS 0.81877f
C462 VTAIL.n24 VSUBS 0.020503f
C463 VTAIL.n25 VSUBS 0.137105f
C464 VTAIL.n26 VSUBS 0.01091f
C465 VTAIL.t0 VSUBS 0.055997f
C466 VTAIL.n27 VSUBS 0.06538f
C467 VTAIL.n28 VSUBS 0.015205f
C468 VTAIL.n29 VSUBS 0.019341f
C469 VTAIL.n30 VSUBS 0.056277f
C470 VTAIL.n31 VSUBS 0.011552f
C471 VTAIL.n32 VSUBS 0.01091f
C472 VTAIL.n33 VSUBS 0.04693f
C473 VTAIL.n34 VSUBS 0.028028f
C474 VTAIL.n35 VSUBS 0.674954f
C475 VTAIL.n36 VSUBS 0.020503f
C476 VTAIL.n37 VSUBS 0.137105f
C477 VTAIL.n38 VSUBS 0.01091f
C478 VTAIL.t3 VSUBS 0.055997f
C479 VTAIL.n39 VSUBS 0.06538f
C480 VTAIL.n40 VSUBS 0.015205f
C481 VTAIL.n41 VSUBS 0.019341f
C482 VTAIL.n42 VSUBS 0.056277f
C483 VTAIL.n43 VSUBS 0.011552f
C484 VTAIL.n44 VSUBS 0.01091f
C485 VTAIL.n45 VSUBS 0.04693f
C486 VTAIL.n46 VSUBS 0.028028f
C487 VTAIL.n47 VSUBS 0.604456f
C488 VN.t0 VSUBS 1.00382f
C489 VN.t1 VSUBS 1.6415f
.ends

