* NGSPICE file created from diff_pair_sample_0786.ext - technology: sky130A

.subckt diff_pair_sample_0786 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t3 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X1 VDD2.t9 VN.t0 VTAIL.t9 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=2.0514 ps=11.3 w=5.26 l=2.26
X2 VTAIL.t18 VP.t1 VDD1.t8 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X3 VTAIL.t4 VN.t1 VDD2.t8 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X4 VDD2.t7 VN.t2 VTAIL.t5 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0.8679 ps=5.59 w=5.26 l=2.26
X5 VDD1.t7 VP.t2 VTAIL.t17 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0.8679 ps=5.59 w=5.26 l=2.26
X6 VDD1.t6 VP.t3 VTAIL.t16 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X7 B.t11 B.t9 B.t10 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0 ps=0 w=5.26 l=2.26
X8 B.t8 B.t6 B.t7 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0 ps=0 w=5.26 l=2.26
X9 VTAIL.t6 VN.t3 VDD2.t6 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X10 VDD2.t5 VN.t4 VTAIL.t8 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=2.0514 ps=11.3 w=5.26 l=2.26
X11 VTAIL.t0 VN.t5 VDD2.t4 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X12 VTAIL.t15 VP.t4 VDD1.t9 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X13 VDD1.t4 VP.t5 VTAIL.t14 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X14 VDD1.t5 VP.t6 VTAIL.t13 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=2.0514 ps=11.3 w=5.26 l=2.26
X15 VDD1.t1 VP.t7 VTAIL.t12 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0.8679 ps=5.59 w=5.26 l=2.26
X16 VDD2.t3 VN.t6 VTAIL.t7 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X17 VDD2.t2 VN.t7 VTAIL.t1 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X18 B.t5 B.t3 B.t4 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0 ps=0 w=5.26 l=2.26
X19 VDD1.t2 VP.t8 VTAIL.t11 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=2.0514 ps=11.3 w=5.26 l=2.26
X20 B.t2 B.t0 B.t1 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0 ps=0 w=5.26 l=2.26
X21 VTAIL.t10 VP.t9 VDD1.t0 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X22 VTAIL.t2 VN.t8 VDD2.t1 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=0.8679 pd=5.59 as=0.8679 ps=5.59 w=5.26 l=2.26
X23 VDD2.t0 VN.t9 VTAIL.t3 w_n4078_n2020# sky130_fd_pr__pfet_01v8 ad=2.0514 pd=11.3 as=0.8679 ps=5.59 w=5.26 l=2.26
R0 VP.n22 VP.n21 161.3
R1 VP.n23 VP.n18 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n17 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n29 VP.n16 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n15 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n14 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n39 VP.n13 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n42 VP.n12 161.3
R14 VP.n44 VP.n43 161.3
R15 VP.n45 VP.n11 161.3
R16 VP.n82 VP.n0 161.3
R17 VP.n81 VP.n80 161.3
R18 VP.n79 VP.n1 161.3
R19 VP.n78 VP.n77 161.3
R20 VP.n76 VP.n2 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n3 161.3
R23 VP.n71 VP.n70 161.3
R24 VP.n69 VP.n4 161.3
R25 VP.n68 VP.n67 161.3
R26 VP.n66 VP.n5 161.3
R27 VP.n65 VP.n64 161.3
R28 VP.n63 VP.n6 161.3
R29 VP.n62 VP.n61 161.3
R30 VP.n60 VP.n7 161.3
R31 VP.n59 VP.n58 161.3
R32 VP.n56 VP.n8 161.3
R33 VP.n55 VP.n54 161.3
R34 VP.n53 VP.n9 161.3
R35 VP.n52 VP.n51 161.3
R36 VP.n50 VP.n10 161.3
R37 VP.n49 VP.n48 102.055
R38 VP.n84 VP.n83 102.055
R39 VP.n47 VP.n46 102.055
R40 VP.n19 VP.t2 86.671
R41 VP.n20 VP.n19 67.8968
R42 VP.n63 VP.n62 56.5617
R43 VP.n70 VP.n69 56.5617
R44 VP.n33 VP.n32 56.5617
R45 VP.n26 VP.n25 56.5617
R46 VP.n5 VP.t3 56.0917
R47 VP.n49 VP.t7 56.0917
R48 VP.n57 VP.t9 56.0917
R49 VP.n75 VP.t4 56.0917
R50 VP.n83 VP.t8 56.0917
R51 VP.n16 VP.t5 56.0917
R52 VP.n46 VP.t6 56.0917
R53 VP.n38 VP.t1 56.0917
R54 VP.n20 VP.t0 56.0917
R55 VP.n55 VP.n9 51.7179
R56 VP.n77 VP.n1 51.7179
R57 VP.n40 VP.n12 51.7179
R58 VP.n48 VP.n47 46.0792
R59 VP.n51 VP.n9 29.4362
R60 VP.n81 VP.n1 29.4362
R61 VP.n44 VP.n12 29.4362
R62 VP.n51 VP.n50 24.5923
R63 VP.n56 VP.n55 24.5923
R64 VP.n58 VP.n7 24.5923
R65 VP.n62 VP.n7 24.5923
R66 VP.n64 VP.n63 24.5923
R67 VP.n64 VP.n5 24.5923
R68 VP.n68 VP.n5 24.5923
R69 VP.n69 VP.n68 24.5923
R70 VP.n70 VP.n3 24.5923
R71 VP.n74 VP.n3 24.5923
R72 VP.n77 VP.n76 24.5923
R73 VP.n82 VP.n81 24.5923
R74 VP.n45 VP.n44 24.5923
R75 VP.n33 VP.n14 24.5923
R76 VP.n37 VP.n14 24.5923
R77 VP.n40 VP.n39 24.5923
R78 VP.n27 VP.n26 24.5923
R79 VP.n27 VP.n16 24.5923
R80 VP.n31 VP.n16 24.5923
R81 VP.n32 VP.n31 24.5923
R82 VP.n21 VP.n18 24.5923
R83 VP.n25 VP.n18 24.5923
R84 VP.n57 VP.n56 20.1658
R85 VP.n76 VP.n75 20.1658
R86 VP.n39 VP.n38 20.1658
R87 VP.n22 VP.n19 10.1113
R88 VP.n50 VP.n49 8.85356
R89 VP.n83 VP.n82 8.85356
R90 VP.n46 VP.n45 8.85356
R91 VP.n58 VP.n57 4.42703
R92 VP.n75 VP.n74 4.42703
R93 VP.n38 VP.n37 4.42703
R94 VP.n21 VP.n20 4.42703
R95 VP.n47 VP.n11 0.278335
R96 VP.n48 VP.n10 0.278335
R97 VP.n84 VP.n0 0.278335
R98 VP.n23 VP.n22 0.189894
R99 VP.n24 VP.n23 0.189894
R100 VP.n24 VP.n17 0.189894
R101 VP.n28 VP.n17 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n30 VP.n29 0.189894
R104 VP.n30 VP.n15 0.189894
R105 VP.n34 VP.n15 0.189894
R106 VP.n35 VP.n34 0.189894
R107 VP.n36 VP.n35 0.189894
R108 VP.n36 VP.n13 0.189894
R109 VP.n41 VP.n13 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n43 VP.n42 0.189894
R112 VP.n43 VP.n11 0.189894
R113 VP.n52 VP.n10 0.189894
R114 VP.n53 VP.n52 0.189894
R115 VP.n54 VP.n53 0.189894
R116 VP.n54 VP.n8 0.189894
R117 VP.n59 VP.n8 0.189894
R118 VP.n60 VP.n59 0.189894
R119 VP.n61 VP.n60 0.189894
R120 VP.n61 VP.n6 0.189894
R121 VP.n65 VP.n6 0.189894
R122 VP.n66 VP.n65 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n67 VP.n4 0.189894
R125 VP.n71 VP.n4 0.189894
R126 VP.n72 VP.n71 0.189894
R127 VP.n73 VP.n72 0.189894
R128 VP.n73 VP.n2 0.189894
R129 VP.n78 VP.n2 0.189894
R130 VP.n79 VP.n78 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n80 VP.n0 0.189894
R133 VP VP.n84 0.153485
R134 VDD1.n22 VDD1.n0 756.745
R135 VDD1.n51 VDD1.n29 756.745
R136 VDD1.n23 VDD1.n22 585
R137 VDD1.n21 VDD1.n20 585
R138 VDD1.n4 VDD1.n3 585
R139 VDD1.n15 VDD1.n14 585
R140 VDD1.n13 VDD1.n12 585
R141 VDD1.n8 VDD1.n7 585
R142 VDD1.n37 VDD1.n36 585
R143 VDD1.n42 VDD1.n41 585
R144 VDD1.n44 VDD1.n43 585
R145 VDD1.n33 VDD1.n32 585
R146 VDD1.n50 VDD1.n49 585
R147 VDD1.n52 VDD1.n51 585
R148 VDD1.n9 VDD1.t7 327.856
R149 VDD1.n38 VDD1.t1 327.856
R150 VDD1.n22 VDD1.n21 171.744
R151 VDD1.n21 VDD1.n3 171.744
R152 VDD1.n14 VDD1.n3 171.744
R153 VDD1.n14 VDD1.n13 171.744
R154 VDD1.n13 VDD1.n7 171.744
R155 VDD1.n42 VDD1.n36 171.744
R156 VDD1.n43 VDD1.n42 171.744
R157 VDD1.n43 VDD1.n32 171.744
R158 VDD1.n50 VDD1.n32 171.744
R159 VDD1.n51 VDD1.n50 171.744
R160 VDD1.n59 VDD1.n58 98.5621
R161 VDD1.n28 VDD1.n27 96.9431
R162 VDD1.n61 VDD1.n60 96.9429
R163 VDD1.n57 VDD1.n56 96.9429
R164 VDD1.t7 VDD1.n7 85.8723
R165 VDD1.t1 VDD1.n36 85.8723
R166 VDD1.n28 VDD1.n26 50.709
R167 VDD1.n57 VDD1.n55 50.709
R168 VDD1.n61 VDD1.n59 40.5548
R169 VDD1.n9 VDD1.n8 16.381
R170 VDD1.n38 VDD1.n37 16.381
R171 VDD1.n12 VDD1.n11 12.8005
R172 VDD1.n41 VDD1.n40 12.8005
R173 VDD1.n15 VDD1.n6 12.0247
R174 VDD1.n44 VDD1.n35 12.0247
R175 VDD1.n16 VDD1.n4 11.249
R176 VDD1.n45 VDD1.n33 11.249
R177 VDD1.n20 VDD1.n19 10.4732
R178 VDD1.n49 VDD1.n48 10.4732
R179 VDD1.n23 VDD1.n2 9.69747
R180 VDD1.n52 VDD1.n31 9.69747
R181 VDD1.n26 VDD1.n25 9.45567
R182 VDD1.n55 VDD1.n54 9.45567
R183 VDD1.n25 VDD1.n24 9.3005
R184 VDD1.n2 VDD1.n1 9.3005
R185 VDD1.n19 VDD1.n18 9.3005
R186 VDD1.n17 VDD1.n16 9.3005
R187 VDD1.n6 VDD1.n5 9.3005
R188 VDD1.n11 VDD1.n10 9.3005
R189 VDD1.n54 VDD1.n53 9.3005
R190 VDD1.n31 VDD1.n30 9.3005
R191 VDD1.n48 VDD1.n47 9.3005
R192 VDD1.n46 VDD1.n45 9.3005
R193 VDD1.n35 VDD1.n34 9.3005
R194 VDD1.n40 VDD1.n39 9.3005
R195 VDD1.n24 VDD1.n0 8.92171
R196 VDD1.n53 VDD1.n29 8.92171
R197 VDD1.n60 VDD1.t8 6.18016
R198 VDD1.n60 VDD1.t5 6.18016
R199 VDD1.n27 VDD1.t3 6.18016
R200 VDD1.n27 VDD1.t4 6.18016
R201 VDD1.n58 VDD1.t9 6.18016
R202 VDD1.n58 VDD1.t2 6.18016
R203 VDD1.n56 VDD1.t0 6.18016
R204 VDD1.n56 VDD1.t6 6.18016
R205 VDD1.n26 VDD1.n0 5.04292
R206 VDD1.n55 VDD1.n29 5.04292
R207 VDD1.n24 VDD1.n23 4.26717
R208 VDD1.n53 VDD1.n52 4.26717
R209 VDD1.n10 VDD1.n9 3.71853
R210 VDD1.n39 VDD1.n38 3.71853
R211 VDD1.n20 VDD1.n2 3.49141
R212 VDD1.n49 VDD1.n31 3.49141
R213 VDD1.n19 VDD1.n4 2.71565
R214 VDD1.n48 VDD1.n33 2.71565
R215 VDD1.n16 VDD1.n15 1.93989
R216 VDD1.n45 VDD1.n44 1.93989
R217 VDD1 VDD1.n61 1.61688
R218 VDD1.n12 VDD1.n6 1.16414
R219 VDD1.n41 VDD1.n35 1.16414
R220 VDD1 VDD1.n28 0.616879
R221 VDD1.n59 VDD1.n57 0.503344
R222 VDD1.n11 VDD1.n8 0.388379
R223 VDD1.n40 VDD1.n37 0.388379
R224 VDD1.n25 VDD1.n1 0.155672
R225 VDD1.n18 VDD1.n1 0.155672
R226 VDD1.n18 VDD1.n17 0.155672
R227 VDD1.n17 VDD1.n5 0.155672
R228 VDD1.n10 VDD1.n5 0.155672
R229 VDD1.n39 VDD1.n34 0.155672
R230 VDD1.n46 VDD1.n34 0.155672
R231 VDD1.n47 VDD1.n46 0.155672
R232 VDD1.n47 VDD1.n30 0.155672
R233 VDD1.n54 VDD1.n30 0.155672
R234 VTAIL.n120 VTAIL.n98 756.745
R235 VTAIL.n24 VTAIL.n2 756.745
R236 VTAIL.n92 VTAIL.n70 756.745
R237 VTAIL.n60 VTAIL.n38 756.745
R238 VTAIL.n106 VTAIL.n105 585
R239 VTAIL.n111 VTAIL.n110 585
R240 VTAIL.n113 VTAIL.n112 585
R241 VTAIL.n102 VTAIL.n101 585
R242 VTAIL.n119 VTAIL.n118 585
R243 VTAIL.n121 VTAIL.n120 585
R244 VTAIL.n10 VTAIL.n9 585
R245 VTAIL.n15 VTAIL.n14 585
R246 VTAIL.n17 VTAIL.n16 585
R247 VTAIL.n6 VTAIL.n5 585
R248 VTAIL.n23 VTAIL.n22 585
R249 VTAIL.n25 VTAIL.n24 585
R250 VTAIL.n93 VTAIL.n92 585
R251 VTAIL.n91 VTAIL.n90 585
R252 VTAIL.n74 VTAIL.n73 585
R253 VTAIL.n85 VTAIL.n84 585
R254 VTAIL.n83 VTAIL.n82 585
R255 VTAIL.n78 VTAIL.n77 585
R256 VTAIL.n61 VTAIL.n60 585
R257 VTAIL.n59 VTAIL.n58 585
R258 VTAIL.n42 VTAIL.n41 585
R259 VTAIL.n53 VTAIL.n52 585
R260 VTAIL.n51 VTAIL.n50 585
R261 VTAIL.n46 VTAIL.n45 585
R262 VTAIL.n107 VTAIL.t9 327.856
R263 VTAIL.n11 VTAIL.t11 327.856
R264 VTAIL.n79 VTAIL.t13 327.856
R265 VTAIL.n47 VTAIL.t8 327.856
R266 VTAIL.n111 VTAIL.n105 171.744
R267 VTAIL.n112 VTAIL.n111 171.744
R268 VTAIL.n112 VTAIL.n101 171.744
R269 VTAIL.n119 VTAIL.n101 171.744
R270 VTAIL.n120 VTAIL.n119 171.744
R271 VTAIL.n15 VTAIL.n9 171.744
R272 VTAIL.n16 VTAIL.n15 171.744
R273 VTAIL.n16 VTAIL.n5 171.744
R274 VTAIL.n23 VTAIL.n5 171.744
R275 VTAIL.n24 VTAIL.n23 171.744
R276 VTAIL.n92 VTAIL.n91 171.744
R277 VTAIL.n91 VTAIL.n73 171.744
R278 VTAIL.n84 VTAIL.n73 171.744
R279 VTAIL.n84 VTAIL.n83 171.744
R280 VTAIL.n83 VTAIL.n77 171.744
R281 VTAIL.n60 VTAIL.n59 171.744
R282 VTAIL.n59 VTAIL.n41 171.744
R283 VTAIL.n52 VTAIL.n41 171.744
R284 VTAIL.n52 VTAIL.n51 171.744
R285 VTAIL.n51 VTAIL.n45 171.744
R286 VTAIL.t9 VTAIL.n105 85.8723
R287 VTAIL.t11 VTAIL.n9 85.8723
R288 VTAIL.t13 VTAIL.n77 85.8723
R289 VTAIL.t8 VTAIL.n45 85.8723
R290 VTAIL.n69 VTAIL.n68 80.2642
R291 VTAIL.n67 VTAIL.n66 80.2642
R292 VTAIL.n37 VTAIL.n36 80.2642
R293 VTAIL.n35 VTAIL.n34 80.2642
R294 VTAIL.n127 VTAIL.n126 80.2641
R295 VTAIL.n1 VTAIL.n0 80.2641
R296 VTAIL.n31 VTAIL.n30 80.2641
R297 VTAIL.n33 VTAIL.n32 80.2641
R298 VTAIL.n125 VTAIL.n124 31.7975
R299 VTAIL.n29 VTAIL.n28 31.7975
R300 VTAIL.n97 VTAIL.n96 31.7975
R301 VTAIL.n65 VTAIL.n64 31.7975
R302 VTAIL.n35 VTAIL.n33 21.3669
R303 VTAIL.n125 VTAIL.n97 19.1341
R304 VTAIL.n107 VTAIL.n106 16.381
R305 VTAIL.n11 VTAIL.n10 16.381
R306 VTAIL.n79 VTAIL.n78 16.381
R307 VTAIL.n47 VTAIL.n46 16.381
R308 VTAIL.n110 VTAIL.n109 12.8005
R309 VTAIL.n14 VTAIL.n13 12.8005
R310 VTAIL.n82 VTAIL.n81 12.8005
R311 VTAIL.n50 VTAIL.n49 12.8005
R312 VTAIL.n113 VTAIL.n104 12.0247
R313 VTAIL.n17 VTAIL.n8 12.0247
R314 VTAIL.n85 VTAIL.n76 12.0247
R315 VTAIL.n53 VTAIL.n44 12.0247
R316 VTAIL.n114 VTAIL.n102 11.249
R317 VTAIL.n18 VTAIL.n6 11.249
R318 VTAIL.n86 VTAIL.n74 11.249
R319 VTAIL.n54 VTAIL.n42 11.249
R320 VTAIL.n118 VTAIL.n117 10.4732
R321 VTAIL.n22 VTAIL.n21 10.4732
R322 VTAIL.n90 VTAIL.n89 10.4732
R323 VTAIL.n58 VTAIL.n57 10.4732
R324 VTAIL.n121 VTAIL.n100 9.69747
R325 VTAIL.n25 VTAIL.n4 9.69747
R326 VTAIL.n93 VTAIL.n72 9.69747
R327 VTAIL.n61 VTAIL.n40 9.69747
R328 VTAIL.n124 VTAIL.n123 9.45567
R329 VTAIL.n28 VTAIL.n27 9.45567
R330 VTAIL.n96 VTAIL.n95 9.45567
R331 VTAIL.n64 VTAIL.n63 9.45567
R332 VTAIL.n123 VTAIL.n122 9.3005
R333 VTAIL.n100 VTAIL.n99 9.3005
R334 VTAIL.n117 VTAIL.n116 9.3005
R335 VTAIL.n115 VTAIL.n114 9.3005
R336 VTAIL.n104 VTAIL.n103 9.3005
R337 VTAIL.n109 VTAIL.n108 9.3005
R338 VTAIL.n27 VTAIL.n26 9.3005
R339 VTAIL.n4 VTAIL.n3 9.3005
R340 VTAIL.n21 VTAIL.n20 9.3005
R341 VTAIL.n19 VTAIL.n18 9.3005
R342 VTAIL.n8 VTAIL.n7 9.3005
R343 VTAIL.n13 VTAIL.n12 9.3005
R344 VTAIL.n95 VTAIL.n94 9.3005
R345 VTAIL.n72 VTAIL.n71 9.3005
R346 VTAIL.n89 VTAIL.n88 9.3005
R347 VTAIL.n87 VTAIL.n86 9.3005
R348 VTAIL.n76 VTAIL.n75 9.3005
R349 VTAIL.n81 VTAIL.n80 9.3005
R350 VTAIL.n63 VTAIL.n62 9.3005
R351 VTAIL.n40 VTAIL.n39 9.3005
R352 VTAIL.n57 VTAIL.n56 9.3005
R353 VTAIL.n55 VTAIL.n54 9.3005
R354 VTAIL.n44 VTAIL.n43 9.3005
R355 VTAIL.n49 VTAIL.n48 9.3005
R356 VTAIL.n122 VTAIL.n98 8.92171
R357 VTAIL.n26 VTAIL.n2 8.92171
R358 VTAIL.n94 VTAIL.n70 8.92171
R359 VTAIL.n62 VTAIL.n38 8.92171
R360 VTAIL.n126 VTAIL.t1 6.18016
R361 VTAIL.n126 VTAIL.t6 6.18016
R362 VTAIL.n0 VTAIL.t3 6.18016
R363 VTAIL.n0 VTAIL.t2 6.18016
R364 VTAIL.n30 VTAIL.t16 6.18016
R365 VTAIL.n30 VTAIL.t15 6.18016
R366 VTAIL.n32 VTAIL.t12 6.18016
R367 VTAIL.n32 VTAIL.t10 6.18016
R368 VTAIL.n68 VTAIL.t14 6.18016
R369 VTAIL.n68 VTAIL.t18 6.18016
R370 VTAIL.n66 VTAIL.t17 6.18016
R371 VTAIL.n66 VTAIL.t19 6.18016
R372 VTAIL.n36 VTAIL.t7 6.18016
R373 VTAIL.n36 VTAIL.t4 6.18016
R374 VTAIL.n34 VTAIL.t5 6.18016
R375 VTAIL.n34 VTAIL.t0 6.18016
R376 VTAIL.n124 VTAIL.n98 5.04292
R377 VTAIL.n28 VTAIL.n2 5.04292
R378 VTAIL.n96 VTAIL.n70 5.04292
R379 VTAIL.n64 VTAIL.n38 5.04292
R380 VTAIL.n122 VTAIL.n121 4.26717
R381 VTAIL.n26 VTAIL.n25 4.26717
R382 VTAIL.n94 VTAIL.n93 4.26717
R383 VTAIL.n62 VTAIL.n61 4.26717
R384 VTAIL.n80 VTAIL.n79 3.71853
R385 VTAIL.n48 VTAIL.n47 3.71853
R386 VTAIL.n108 VTAIL.n107 3.71853
R387 VTAIL.n12 VTAIL.n11 3.71853
R388 VTAIL.n118 VTAIL.n100 3.49141
R389 VTAIL.n22 VTAIL.n4 3.49141
R390 VTAIL.n90 VTAIL.n72 3.49141
R391 VTAIL.n58 VTAIL.n40 3.49141
R392 VTAIL.n117 VTAIL.n102 2.71565
R393 VTAIL.n21 VTAIL.n6 2.71565
R394 VTAIL.n89 VTAIL.n74 2.71565
R395 VTAIL.n57 VTAIL.n42 2.71565
R396 VTAIL.n37 VTAIL.n35 2.23326
R397 VTAIL.n65 VTAIL.n37 2.23326
R398 VTAIL.n69 VTAIL.n67 2.23326
R399 VTAIL.n97 VTAIL.n69 2.23326
R400 VTAIL.n33 VTAIL.n31 2.23326
R401 VTAIL.n31 VTAIL.n29 2.23326
R402 VTAIL.n127 VTAIL.n125 2.23326
R403 VTAIL.n114 VTAIL.n113 1.93989
R404 VTAIL.n18 VTAIL.n17 1.93989
R405 VTAIL.n86 VTAIL.n85 1.93989
R406 VTAIL.n54 VTAIL.n53 1.93989
R407 VTAIL VTAIL.n1 1.73326
R408 VTAIL.n67 VTAIL.n65 1.58671
R409 VTAIL.n29 VTAIL.n1 1.58671
R410 VTAIL.n110 VTAIL.n104 1.16414
R411 VTAIL.n14 VTAIL.n8 1.16414
R412 VTAIL.n82 VTAIL.n76 1.16414
R413 VTAIL.n50 VTAIL.n44 1.16414
R414 VTAIL VTAIL.n127 0.5005
R415 VTAIL.n109 VTAIL.n106 0.388379
R416 VTAIL.n13 VTAIL.n10 0.388379
R417 VTAIL.n81 VTAIL.n78 0.388379
R418 VTAIL.n49 VTAIL.n46 0.388379
R419 VTAIL.n108 VTAIL.n103 0.155672
R420 VTAIL.n115 VTAIL.n103 0.155672
R421 VTAIL.n116 VTAIL.n115 0.155672
R422 VTAIL.n116 VTAIL.n99 0.155672
R423 VTAIL.n123 VTAIL.n99 0.155672
R424 VTAIL.n12 VTAIL.n7 0.155672
R425 VTAIL.n19 VTAIL.n7 0.155672
R426 VTAIL.n20 VTAIL.n19 0.155672
R427 VTAIL.n20 VTAIL.n3 0.155672
R428 VTAIL.n27 VTAIL.n3 0.155672
R429 VTAIL.n95 VTAIL.n71 0.155672
R430 VTAIL.n88 VTAIL.n71 0.155672
R431 VTAIL.n88 VTAIL.n87 0.155672
R432 VTAIL.n87 VTAIL.n75 0.155672
R433 VTAIL.n80 VTAIL.n75 0.155672
R434 VTAIL.n63 VTAIL.n39 0.155672
R435 VTAIL.n56 VTAIL.n39 0.155672
R436 VTAIL.n56 VTAIL.n55 0.155672
R437 VTAIL.n55 VTAIL.n43 0.155672
R438 VTAIL.n48 VTAIL.n43 0.155672
R439 VN.n71 VN.n37 161.3
R440 VN.n70 VN.n69 161.3
R441 VN.n68 VN.n38 161.3
R442 VN.n67 VN.n66 161.3
R443 VN.n65 VN.n39 161.3
R444 VN.n63 VN.n62 161.3
R445 VN.n61 VN.n40 161.3
R446 VN.n60 VN.n59 161.3
R447 VN.n58 VN.n41 161.3
R448 VN.n57 VN.n56 161.3
R449 VN.n55 VN.n42 161.3
R450 VN.n54 VN.n53 161.3
R451 VN.n52 VN.n43 161.3
R452 VN.n51 VN.n50 161.3
R453 VN.n49 VN.n44 161.3
R454 VN.n48 VN.n47 161.3
R455 VN.n34 VN.n0 161.3
R456 VN.n33 VN.n32 161.3
R457 VN.n31 VN.n1 161.3
R458 VN.n30 VN.n29 161.3
R459 VN.n28 VN.n2 161.3
R460 VN.n26 VN.n25 161.3
R461 VN.n24 VN.n3 161.3
R462 VN.n23 VN.n22 161.3
R463 VN.n21 VN.n4 161.3
R464 VN.n20 VN.n19 161.3
R465 VN.n18 VN.n5 161.3
R466 VN.n17 VN.n16 161.3
R467 VN.n15 VN.n6 161.3
R468 VN.n14 VN.n13 161.3
R469 VN.n12 VN.n7 161.3
R470 VN.n11 VN.n10 161.3
R471 VN.n36 VN.n35 102.055
R472 VN.n73 VN.n72 102.055
R473 VN.n8 VN.t9 86.671
R474 VN.n45 VN.t4 86.671
R475 VN.n9 VN.n8 67.8968
R476 VN.n46 VN.n45 67.8968
R477 VN.n15 VN.n14 56.5617
R478 VN.n22 VN.n21 56.5617
R479 VN.n52 VN.n51 56.5617
R480 VN.n59 VN.n58 56.5617
R481 VN.n5 VN.t7 56.0917
R482 VN.n9 VN.t8 56.0917
R483 VN.n27 VN.t3 56.0917
R484 VN.n35 VN.t0 56.0917
R485 VN.n42 VN.t6 56.0917
R486 VN.n46 VN.t1 56.0917
R487 VN.n64 VN.t5 56.0917
R488 VN.n72 VN.t2 56.0917
R489 VN.n29 VN.n1 51.7179
R490 VN.n66 VN.n38 51.7179
R491 VN VN.n73 46.358
R492 VN.n33 VN.n1 29.4362
R493 VN.n70 VN.n38 29.4362
R494 VN.n10 VN.n7 24.5923
R495 VN.n14 VN.n7 24.5923
R496 VN.n16 VN.n15 24.5923
R497 VN.n16 VN.n5 24.5923
R498 VN.n20 VN.n5 24.5923
R499 VN.n21 VN.n20 24.5923
R500 VN.n22 VN.n3 24.5923
R501 VN.n26 VN.n3 24.5923
R502 VN.n29 VN.n28 24.5923
R503 VN.n34 VN.n33 24.5923
R504 VN.n51 VN.n44 24.5923
R505 VN.n47 VN.n44 24.5923
R506 VN.n58 VN.n57 24.5923
R507 VN.n57 VN.n42 24.5923
R508 VN.n53 VN.n42 24.5923
R509 VN.n53 VN.n52 24.5923
R510 VN.n66 VN.n65 24.5923
R511 VN.n63 VN.n40 24.5923
R512 VN.n59 VN.n40 24.5923
R513 VN.n71 VN.n70 24.5923
R514 VN.n28 VN.n27 20.1658
R515 VN.n65 VN.n64 20.1658
R516 VN.n48 VN.n45 10.1113
R517 VN.n11 VN.n8 10.1113
R518 VN.n35 VN.n34 8.85356
R519 VN.n72 VN.n71 8.85356
R520 VN.n10 VN.n9 4.42703
R521 VN.n27 VN.n26 4.42703
R522 VN.n47 VN.n46 4.42703
R523 VN.n64 VN.n63 4.42703
R524 VN.n73 VN.n37 0.278335
R525 VN.n36 VN.n0 0.278335
R526 VN.n69 VN.n37 0.189894
R527 VN.n69 VN.n68 0.189894
R528 VN.n68 VN.n67 0.189894
R529 VN.n67 VN.n39 0.189894
R530 VN.n62 VN.n39 0.189894
R531 VN.n62 VN.n61 0.189894
R532 VN.n61 VN.n60 0.189894
R533 VN.n60 VN.n41 0.189894
R534 VN.n56 VN.n41 0.189894
R535 VN.n56 VN.n55 0.189894
R536 VN.n55 VN.n54 0.189894
R537 VN.n54 VN.n43 0.189894
R538 VN.n50 VN.n43 0.189894
R539 VN.n50 VN.n49 0.189894
R540 VN.n49 VN.n48 0.189894
R541 VN.n12 VN.n11 0.189894
R542 VN.n13 VN.n12 0.189894
R543 VN.n13 VN.n6 0.189894
R544 VN.n17 VN.n6 0.189894
R545 VN.n18 VN.n17 0.189894
R546 VN.n19 VN.n18 0.189894
R547 VN.n19 VN.n4 0.189894
R548 VN.n23 VN.n4 0.189894
R549 VN.n24 VN.n23 0.189894
R550 VN.n25 VN.n24 0.189894
R551 VN.n25 VN.n2 0.189894
R552 VN.n30 VN.n2 0.189894
R553 VN.n31 VN.n30 0.189894
R554 VN.n32 VN.n31 0.189894
R555 VN.n32 VN.n0 0.189894
R556 VN VN.n36 0.153485
R557 VDD2.n53 VDD2.n31 756.745
R558 VDD2.n22 VDD2.n0 756.745
R559 VDD2.n54 VDD2.n53 585
R560 VDD2.n52 VDD2.n51 585
R561 VDD2.n35 VDD2.n34 585
R562 VDD2.n46 VDD2.n45 585
R563 VDD2.n44 VDD2.n43 585
R564 VDD2.n39 VDD2.n38 585
R565 VDD2.n8 VDD2.n7 585
R566 VDD2.n13 VDD2.n12 585
R567 VDD2.n15 VDD2.n14 585
R568 VDD2.n4 VDD2.n3 585
R569 VDD2.n21 VDD2.n20 585
R570 VDD2.n23 VDD2.n22 585
R571 VDD2.n40 VDD2.t7 327.856
R572 VDD2.n9 VDD2.t0 327.856
R573 VDD2.n53 VDD2.n52 171.744
R574 VDD2.n52 VDD2.n34 171.744
R575 VDD2.n45 VDD2.n34 171.744
R576 VDD2.n45 VDD2.n44 171.744
R577 VDD2.n44 VDD2.n38 171.744
R578 VDD2.n13 VDD2.n7 171.744
R579 VDD2.n14 VDD2.n13 171.744
R580 VDD2.n14 VDD2.n3 171.744
R581 VDD2.n21 VDD2.n3 171.744
R582 VDD2.n22 VDD2.n21 171.744
R583 VDD2.n30 VDD2.n29 98.5621
R584 VDD2 VDD2.n61 98.5593
R585 VDD2.n60 VDD2.n59 96.9431
R586 VDD2.n28 VDD2.n27 96.9429
R587 VDD2.t7 VDD2.n38 85.8723
R588 VDD2.t0 VDD2.n7 85.8723
R589 VDD2.n28 VDD2.n26 50.709
R590 VDD2.n58 VDD2.n57 48.4763
R591 VDD2.n58 VDD2.n30 38.8554
R592 VDD2.n40 VDD2.n39 16.381
R593 VDD2.n9 VDD2.n8 16.381
R594 VDD2.n43 VDD2.n42 12.8005
R595 VDD2.n12 VDD2.n11 12.8005
R596 VDD2.n46 VDD2.n37 12.0247
R597 VDD2.n15 VDD2.n6 12.0247
R598 VDD2.n47 VDD2.n35 11.249
R599 VDD2.n16 VDD2.n4 11.249
R600 VDD2.n51 VDD2.n50 10.4732
R601 VDD2.n20 VDD2.n19 10.4732
R602 VDD2.n54 VDD2.n33 9.69747
R603 VDD2.n23 VDD2.n2 9.69747
R604 VDD2.n57 VDD2.n56 9.45567
R605 VDD2.n26 VDD2.n25 9.45567
R606 VDD2.n56 VDD2.n55 9.3005
R607 VDD2.n33 VDD2.n32 9.3005
R608 VDD2.n50 VDD2.n49 9.3005
R609 VDD2.n48 VDD2.n47 9.3005
R610 VDD2.n37 VDD2.n36 9.3005
R611 VDD2.n42 VDD2.n41 9.3005
R612 VDD2.n25 VDD2.n24 9.3005
R613 VDD2.n2 VDD2.n1 9.3005
R614 VDD2.n19 VDD2.n18 9.3005
R615 VDD2.n17 VDD2.n16 9.3005
R616 VDD2.n6 VDD2.n5 9.3005
R617 VDD2.n11 VDD2.n10 9.3005
R618 VDD2.n55 VDD2.n31 8.92171
R619 VDD2.n24 VDD2.n0 8.92171
R620 VDD2.n61 VDD2.t8 6.18016
R621 VDD2.n61 VDD2.t5 6.18016
R622 VDD2.n59 VDD2.t4 6.18016
R623 VDD2.n59 VDD2.t3 6.18016
R624 VDD2.n29 VDD2.t6 6.18016
R625 VDD2.n29 VDD2.t9 6.18016
R626 VDD2.n27 VDD2.t1 6.18016
R627 VDD2.n27 VDD2.t2 6.18016
R628 VDD2.n57 VDD2.n31 5.04292
R629 VDD2.n26 VDD2.n0 5.04292
R630 VDD2.n55 VDD2.n54 4.26717
R631 VDD2.n24 VDD2.n23 4.26717
R632 VDD2.n41 VDD2.n40 3.71853
R633 VDD2.n10 VDD2.n9 3.71853
R634 VDD2.n51 VDD2.n33 3.49141
R635 VDD2.n20 VDD2.n2 3.49141
R636 VDD2.n50 VDD2.n35 2.71565
R637 VDD2.n19 VDD2.n4 2.71565
R638 VDD2.n60 VDD2.n58 2.23326
R639 VDD2.n47 VDD2.n46 1.93989
R640 VDD2.n16 VDD2.n15 1.93989
R641 VDD2.n43 VDD2.n37 1.16414
R642 VDD2.n12 VDD2.n6 1.16414
R643 VDD2 VDD2.n60 0.616879
R644 VDD2.n30 VDD2.n28 0.503344
R645 VDD2.n42 VDD2.n39 0.388379
R646 VDD2.n11 VDD2.n8 0.388379
R647 VDD2.n56 VDD2.n32 0.155672
R648 VDD2.n49 VDD2.n32 0.155672
R649 VDD2.n49 VDD2.n48 0.155672
R650 VDD2.n48 VDD2.n36 0.155672
R651 VDD2.n41 VDD2.n36 0.155672
R652 VDD2.n10 VDD2.n5 0.155672
R653 VDD2.n17 VDD2.n5 0.155672
R654 VDD2.n18 VDD2.n17 0.155672
R655 VDD2.n18 VDD2.n1 0.155672
R656 VDD2.n25 VDD2.n1 0.155672
R657 B.n497 B.n496 585
R658 B.n498 B.n59 585
R659 B.n500 B.n499 585
R660 B.n501 B.n58 585
R661 B.n503 B.n502 585
R662 B.n504 B.n57 585
R663 B.n506 B.n505 585
R664 B.n507 B.n56 585
R665 B.n509 B.n508 585
R666 B.n510 B.n55 585
R667 B.n512 B.n511 585
R668 B.n513 B.n54 585
R669 B.n515 B.n514 585
R670 B.n516 B.n53 585
R671 B.n518 B.n517 585
R672 B.n519 B.n52 585
R673 B.n521 B.n520 585
R674 B.n522 B.n51 585
R675 B.n524 B.n523 585
R676 B.n525 B.n50 585
R677 B.n527 B.n526 585
R678 B.n528 B.n47 585
R679 B.n531 B.n530 585
R680 B.n532 B.n46 585
R681 B.n534 B.n533 585
R682 B.n535 B.n45 585
R683 B.n537 B.n536 585
R684 B.n538 B.n44 585
R685 B.n540 B.n539 585
R686 B.n541 B.n43 585
R687 B.n543 B.n542 585
R688 B.n545 B.n544 585
R689 B.n546 B.n39 585
R690 B.n548 B.n547 585
R691 B.n549 B.n38 585
R692 B.n551 B.n550 585
R693 B.n552 B.n37 585
R694 B.n554 B.n553 585
R695 B.n555 B.n36 585
R696 B.n557 B.n556 585
R697 B.n558 B.n35 585
R698 B.n560 B.n559 585
R699 B.n561 B.n34 585
R700 B.n563 B.n562 585
R701 B.n564 B.n33 585
R702 B.n566 B.n565 585
R703 B.n567 B.n32 585
R704 B.n569 B.n568 585
R705 B.n570 B.n31 585
R706 B.n572 B.n571 585
R707 B.n573 B.n30 585
R708 B.n575 B.n574 585
R709 B.n576 B.n29 585
R710 B.n495 B.n60 585
R711 B.n494 B.n493 585
R712 B.n492 B.n61 585
R713 B.n491 B.n490 585
R714 B.n489 B.n62 585
R715 B.n488 B.n487 585
R716 B.n486 B.n63 585
R717 B.n485 B.n484 585
R718 B.n483 B.n64 585
R719 B.n482 B.n481 585
R720 B.n480 B.n65 585
R721 B.n479 B.n478 585
R722 B.n477 B.n66 585
R723 B.n476 B.n475 585
R724 B.n474 B.n67 585
R725 B.n473 B.n472 585
R726 B.n471 B.n68 585
R727 B.n470 B.n469 585
R728 B.n468 B.n69 585
R729 B.n467 B.n466 585
R730 B.n465 B.n70 585
R731 B.n464 B.n463 585
R732 B.n462 B.n71 585
R733 B.n461 B.n460 585
R734 B.n459 B.n72 585
R735 B.n458 B.n457 585
R736 B.n456 B.n73 585
R737 B.n455 B.n454 585
R738 B.n453 B.n74 585
R739 B.n452 B.n451 585
R740 B.n450 B.n75 585
R741 B.n449 B.n448 585
R742 B.n447 B.n76 585
R743 B.n446 B.n445 585
R744 B.n444 B.n77 585
R745 B.n443 B.n442 585
R746 B.n441 B.n78 585
R747 B.n440 B.n439 585
R748 B.n438 B.n79 585
R749 B.n437 B.n436 585
R750 B.n435 B.n80 585
R751 B.n434 B.n433 585
R752 B.n432 B.n81 585
R753 B.n431 B.n430 585
R754 B.n429 B.n82 585
R755 B.n428 B.n427 585
R756 B.n426 B.n83 585
R757 B.n425 B.n424 585
R758 B.n423 B.n84 585
R759 B.n422 B.n421 585
R760 B.n420 B.n85 585
R761 B.n419 B.n418 585
R762 B.n417 B.n86 585
R763 B.n416 B.n415 585
R764 B.n414 B.n87 585
R765 B.n413 B.n412 585
R766 B.n411 B.n88 585
R767 B.n410 B.n409 585
R768 B.n408 B.n89 585
R769 B.n407 B.n406 585
R770 B.n405 B.n90 585
R771 B.n404 B.n403 585
R772 B.n402 B.n91 585
R773 B.n401 B.n400 585
R774 B.n399 B.n92 585
R775 B.n398 B.n397 585
R776 B.n396 B.n93 585
R777 B.n395 B.n394 585
R778 B.n393 B.n94 585
R779 B.n392 B.n391 585
R780 B.n390 B.n95 585
R781 B.n389 B.n388 585
R782 B.n387 B.n96 585
R783 B.n386 B.n385 585
R784 B.n384 B.n97 585
R785 B.n383 B.n382 585
R786 B.n381 B.n98 585
R787 B.n380 B.n379 585
R788 B.n378 B.n99 585
R789 B.n377 B.n376 585
R790 B.n375 B.n100 585
R791 B.n374 B.n373 585
R792 B.n372 B.n101 585
R793 B.n371 B.n370 585
R794 B.n369 B.n102 585
R795 B.n368 B.n367 585
R796 B.n366 B.n103 585
R797 B.n365 B.n364 585
R798 B.n363 B.n104 585
R799 B.n362 B.n361 585
R800 B.n360 B.n105 585
R801 B.n359 B.n358 585
R802 B.n357 B.n106 585
R803 B.n356 B.n355 585
R804 B.n354 B.n107 585
R805 B.n353 B.n352 585
R806 B.n351 B.n108 585
R807 B.n350 B.n349 585
R808 B.n348 B.n109 585
R809 B.n347 B.n346 585
R810 B.n345 B.n110 585
R811 B.n344 B.n343 585
R812 B.n342 B.n111 585
R813 B.n341 B.n340 585
R814 B.n339 B.n112 585
R815 B.n338 B.n337 585
R816 B.n336 B.n113 585
R817 B.n335 B.n334 585
R818 B.n333 B.n114 585
R819 B.n252 B.n145 585
R820 B.n254 B.n253 585
R821 B.n255 B.n144 585
R822 B.n257 B.n256 585
R823 B.n258 B.n143 585
R824 B.n260 B.n259 585
R825 B.n261 B.n142 585
R826 B.n263 B.n262 585
R827 B.n264 B.n141 585
R828 B.n266 B.n265 585
R829 B.n267 B.n140 585
R830 B.n269 B.n268 585
R831 B.n270 B.n139 585
R832 B.n272 B.n271 585
R833 B.n273 B.n138 585
R834 B.n275 B.n274 585
R835 B.n276 B.n137 585
R836 B.n278 B.n277 585
R837 B.n279 B.n136 585
R838 B.n281 B.n280 585
R839 B.n282 B.n135 585
R840 B.n284 B.n283 585
R841 B.n286 B.n285 585
R842 B.n287 B.n131 585
R843 B.n289 B.n288 585
R844 B.n290 B.n130 585
R845 B.n292 B.n291 585
R846 B.n293 B.n129 585
R847 B.n295 B.n294 585
R848 B.n296 B.n128 585
R849 B.n298 B.n297 585
R850 B.n300 B.n125 585
R851 B.n302 B.n301 585
R852 B.n303 B.n124 585
R853 B.n305 B.n304 585
R854 B.n306 B.n123 585
R855 B.n308 B.n307 585
R856 B.n309 B.n122 585
R857 B.n311 B.n310 585
R858 B.n312 B.n121 585
R859 B.n314 B.n313 585
R860 B.n315 B.n120 585
R861 B.n317 B.n316 585
R862 B.n318 B.n119 585
R863 B.n320 B.n319 585
R864 B.n321 B.n118 585
R865 B.n323 B.n322 585
R866 B.n324 B.n117 585
R867 B.n326 B.n325 585
R868 B.n327 B.n116 585
R869 B.n329 B.n328 585
R870 B.n330 B.n115 585
R871 B.n332 B.n331 585
R872 B.n251 B.n250 585
R873 B.n249 B.n146 585
R874 B.n248 B.n247 585
R875 B.n246 B.n147 585
R876 B.n245 B.n244 585
R877 B.n243 B.n148 585
R878 B.n242 B.n241 585
R879 B.n240 B.n149 585
R880 B.n239 B.n238 585
R881 B.n237 B.n150 585
R882 B.n236 B.n235 585
R883 B.n234 B.n151 585
R884 B.n233 B.n232 585
R885 B.n231 B.n152 585
R886 B.n230 B.n229 585
R887 B.n228 B.n153 585
R888 B.n227 B.n226 585
R889 B.n225 B.n154 585
R890 B.n224 B.n223 585
R891 B.n222 B.n155 585
R892 B.n221 B.n220 585
R893 B.n219 B.n156 585
R894 B.n218 B.n217 585
R895 B.n216 B.n157 585
R896 B.n215 B.n214 585
R897 B.n213 B.n158 585
R898 B.n212 B.n211 585
R899 B.n210 B.n159 585
R900 B.n209 B.n208 585
R901 B.n207 B.n160 585
R902 B.n206 B.n205 585
R903 B.n204 B.n161 585
R904 B.n203 B.n202 585
R905 B.n201 B.n162 585
R906 B.n200 B.n199 585
R907 B.n198 B.n163 585
R908 B.n197 B.n196 585
R909 B.n195 B.n164 585
R910 B.n194 B.n193 585
R911 B.n192 B.n165 585
R912 B.n191 B.n190 585
R913 B.n189 B.n166 585
R914 B.n188 B.n187 585
R915 B.n186 B.n167 585
R916 B.n185 B.n184 585
R917 B.n183 B.n168 585
R918 B.n182 B.n181 585
R919 B.n180 B.n169 585
R920 B.n179 B.n178 585
R921 B.n177 B.n170 585
R922 B.n176 B.n175 585
R923 B.n174 B.n171 585
R924 B.n173 B.n172 585
R925 B.n2 B.n0 585
R926 B.n657 B.n1 585
R927 B.n656 B.n655 585
R928 B.n654 B.n3 585
R929 B.n653 B.n652 585
R930 B.n651 B.n4 585
R931 B.n650 B.n649 585
R932 B.n648 B.n5 585
R933 B.n647 B.n646 585
R934 B.n645 B.n6 585
R935 B.n644 B.n643 585
R936 B.n642 B.n7 585
R937 B.n641 B.n640 585
R938 B.n639 B.n8 585
R939 B.n638 B.n637 585
R940 B.n636 B.n9 585
R941 B.n635 B.n634 585
R942 B.n633 B.n10 585
R943 B.n632 B.n631 585
R944 B.n630 B.n11 585
R945 B.n629 B.n628 585
R946 B.n627 B.n12 585
R947 B.n626 B.n625 585
R948 B.n624 B.n13 585
R949 B.n623 B.n622 585
R950 B.n621 B.n14 585
R951 B.n620 B.n619 585
R952 B.n618 B.n15 585
R953 B.n617 B.n616 585
R954 B.n615 B.n16 585
R955 B.n614 B.n613 585
R956 B.n612 B.n17 585
R957 B.n611 B.n610 585
R958 B.n609 B.n18 585
R959 B.n608 B.n607 585
R960 B.n606 B.n19 585
R961 B.n605 B.n604 585
R962 B.n603 B.n20 585
R963 B.n602 B.n601 585
R964 B.n600 B.n21 585
R965 B.n599 B.n598 585
R966 B.n597 B.n22 585
R967 B.n596 B.n595 585
R968 B.n594 B.n23 585
R969 B.n593 B.n592 585
R970 B.n591 B.n24 585
R971 B.n590 B.n589 585
R972 B.n588 B.n25 585
R973 B.n587 B.n586 585
R974 B.n585 B.n26 585
R975 B.n584 B.n583 585
R976 B.n582 B.n27 585
R977 B.n581 B.n580 585
R978 B.n579 B.n28 585
R979 B.n578 B.n577 585
R980 B.n659 B.n658 585
R981 B.n250 B.n145 482.89
R982 B.n578 B.n29 482.89
R983 B.n333 B.n332 482.89
R984 B.n496 B.n495 482.89
R985 B.n126 B.t8 305.49
R986 B.n48 B.t4 305.49
R987 B.n132 B.t11 305.49
R988 B.n40 B.t1 305.49
R989 B.n126 B.t6 263.56
R990 B.n132 B.t9 263.56
R991 B.n40 B.t0 263.56
R992 B.n48 B.t3 263.56
R993 B.n127 B.t7 255.261
R994 B.n49 B.t5 255.261
R995 B.n133 B.t10 255.261
R996 B.n41 B.t2 255.261
R997 B.n250 B.n249 163.367
R998 B.n249 B.n248 163.367
R999 B.n248 B.n147 163.367
R1000 B.n244 B.n147 163.367
R1001 B.n244 B.n243 163.367
R1002 B.n243 B.n242 163.367
R1003 B.n242 B.n149 163.367
R1004 B.n238 B.n149 163.367
R1005 B.n238 B.n237 163.367
R1006 B.n237 B.n236 163.367
R1007 B.n236 B.n151 163.367
R1008 B.n232 B.n151 163.367
R1009 B.n232 B.n231 163.367
R1010 B.n231 B.n230 163.367
R1011 B.n230 B.n153 163.367
R1012 B.n226 B.n153 163.367
R1013 B.n226 B.n225 163.367
R1014 B.n225 B.n224 163.367
R1015 B.n224 B.n155 163.367
R1016 B.n220 B.n155 163.367
R1017 B.n220 B.n219 163.367
R1018 B.n219 B.n218 163.367
R1019 B.n218 B.n157 163.367
R1020 B.n214 B.n157 163.367
R1021 B.n214 B.n213 163.367
R1022 B.n213 B.n212 163.367
R1023 B.n212 B.n159 163.367
R1024 B.n208 B.n159 163.367
R1025 B.n208 B.n207 163.367
R1026 B.n207 B.n206 163.367
R1027 B.n206 B.n161 163.367
R1028 B.n202 B.n161 163.367
R1029 B.n202 B.n201 163.367
R1030 B.n201 B.n200 163.367
R1031 B.n200 B.n163 163.367
R1032 B.n196 B.n163 163.367
R1033 B.n196 B.n195 163.367
R1034 B.n195 B.n194 163.367
R1035 B.n194 B.n165 163.367
R1036 B.n190 B.n165 163.367
R1037 B.n190 B.n189 163.367
R1038 B.n189 B.n188 163.367
R1039 B.n188 B.n167 163.367
R1040 B.n184 B.n167 163.367
R1041 B.n184 B.n183 163.367
R1042 B.n183 B.n182 163.367
R1043 B.n182 B.n169 163.367
R1044 B.n178 B.n169 163.367
R1045 B.n178 B.n177 163.367
R1046 B.n177 B.n176 163.367
R1047 B.n176 B.n171 163.367
R1048 B.n172 B.n171 163.367
R1049 B.n172 B.n2 163.367
R1050 B.n658 B.n2 163.367
R1051 B.n658 B.n657 163.367
R1052 B.n657 B.n656 163.367
R1053 B.n656 B.n3 163.367
R1054 B.n652 B.n3 163.367
R1055 B.n652 B.n651 163.367
R1056 B.n651 B.n650 163.367
R1057 B.n650 B.n5 163.367
R1058 B.n646 B.n5 163.367
R1059 B.n646 B.n645 163.367
R1060 B.n645 B.n644 163.367
R1061 B.n644 B.n7 163.367
R1062 B.n640 B.n7 163.367
R1063 B.n640 B.n639 163.367
R1064 B.n639 B.n638 163.367
R1065 B.n638 B.n9 163.367
R1066 B.n634 B.n9 163.367
R1067 B.n634 B.n633 163.367
R1068 B.n633 B.n632 163.367
R1069 B.n632 B.n11 163.367
R1070 B.n628 B.n11 163.367
R1071 B.n628 B.n627 163.367
R1072 B.n627 B.n626 163.367
R1073 B.n626 B.n13 163.367
R1074 B.n622 B.n13 163.367
R1075 B.n622 B.n621 163.367
R1076 B.n621 B.n620 163.367
R1077 B.n620 B.n15 163.367
R1078 B.n616 B.n15 163.367
R1079 B.n616 B.n615 163.367
R1080 B.n615 B.n614 163.367
R1081 B.n614 B.n17 163.367
R1082 B.n610 B.n17 163.367
R1083 B.n610 B.n609 163.367
R1084 B.n609 B.n608 163.367
R1085 B.n608 B.n19 163.367
R1086 B.n604 B.n19 163.367
R1087 B.n604 B.n603 163.367
R1088 B.n603 B.n602 163.367
R1089 B.n602 B.n21 163.367
R1090 B.n598 B.n21 163.367
R1091 B.n598 B.n597 163.367
R1092 B.n597 B.n596 163.367
R1093 B.n596 B.n23 163.367
R1094 B.n592 B.n23 163.367
R1095 B.n592 B.n591 163.367
R1096 B.n591 B.n590 163.367
R1097 B.n590 B.n25 163.367
R1098 B.n586 B.n25 163.367
R1099 B.n586 B.n585 163.367
R1100 B.n585 B.n584 163.367
R1101 B.n584 B.n27 163.367
R1102 B.n580 B.n27 163.367
R1103 B.n580 B.n579 163.367
R1104 B.n579 B.n578 163.367
R1105 B.n254 B.n145 163.367
R1106 B.n255 B.n254 163.367
R1107 B.n256 B.n255 163.367
R1108 B.n256 B.n143 163.367
R1109 B.n260 B.n143 163.367
R1110 B.n261 B.n260 163.367
R1111 B.n262 B.n261 163.367
R1112 B.n262 B.n141 163.367
R1113 B.n266 B.n141 163.367
R1114 B.n267 B.n266 163.367
R1115 B.n268 B.n267 163.367
R1116 B.n268 B.n139 163.367
R1117 B.n272 B.n139 163.367
R1118 B.n273 B.n272 163.367
R1119 B.n274 B.n273 163.367
R1120 B.n274 B.n137 163.367
R1121 B.n278 B.n137 163.367
R1122 B.n279 B.n278 163.367
R1123 B.n280 B.n279 163.367
R1124 B.n280 B.n135 163.367
R1125 B.n284 B.n135 163.367
R1126 B.n285 B.n284 163.367
R1127 B.n285 B.n131 163.367
R1128 B.n289 B.n131 163.367
R1129 B.n290 B.n289 163.367
R1130 B.n291 B.n290 163.367
R1131 B.n291 B.n129 163.367
R1132 B.n295 B.n129 163.367
R1133 B.n296 B.n295 163.367
R1134 B.n297 B.n296 163.367
R1135 B.n297 B.n125 163.367
R1136 B.n302 B.n125 163.367
R1137 B.n303 B.n302 163.367
R1138 B.n304 B.n303 163.367
R1139 B.n304 B.n123 163.367
R1140 B.n308 B.n123 163.367
R1141 B.n309 B.n308 163.367
R1142 B.n310 B.n309 163.367
R1143 B.n310 B.n121 163.367
R1144 B.n314 B.n121 163.367
R1145 B.n315 B.n314 163.367
R1146 B.n316 B.n315 163.367
R1147 B.n316 B.n119 163.367
R1148 B.n320 B.n119 163.367
R1149 B.n321 B.n320 163.367
R1150 B.n322 B.n321 163.367
R1151 B.n322 B.n117 163.367
R1152 B.n326 B.n117 163.367
R1153 B.n327 B.n326 163.367
R1154 B.n328 B.n327 163.367
R1155 B.n328 B.n115 163.367
R1156 B.n332 B.n115 163.367
R1157 B.n334 B.n333 163.367
R1158 B.n334 B.n113 163.367
R1159 B.n338 B.n113 163.367
R1160 B.n339 B.n338 163.367
R1161 B.n340 B.n339 163.367
R1162 B.n340 B.n111 163.367
R1163 B.n344 B.n111 163.367
R1164 B.n345 B.n344 163.367
R1165 B.n346 B.n345 163.367
R1166 B.n346 B.n109 163.367
R1167 B.n350 B.n109 163.367
R1168 B.n351 B.n350 163.367
R1169 B.n352 B.n351 163.367
R1170 B.n352 B.n107 163.367
R1171 B.n356 B.n107 163.367
R1172 B.n357 B.n356 163.367
R1173 B.n358 B.n357 163.367
R1174 B.n358 B.n105 163.367
R1175 B.n362 B.n105 163.367
R1176 B.n363 B.n362 163.367
R1177 B.n364 B.n363 163.367
R1178 B.n364 B.n103 163.367
R1179 B.n368 B.n103 163.367
R1180 B.n369 B.n368 163.367
R1181 B.n370 B.n369 163.367
R1182 B.n370 B.n101 163.367
R1183 B.n374 B.n101 163.367
R1184 B.n375 B.n374 163.367
R1185 B.n376 B.n375 163.367
R1186 B.n376 B.n99 163.367
R1187 B.n380 B.n99 163.367
R1188 B.n381 B.n380 163.367
R1189 B.n382 B.n381 163.367
R1190 B.n382 B.n97 163.367
R1191 B.n386 B.n97 163.367
R1192 B.n387 B.n386 163.367
R1193 B.n388 B.n387 163.367
R1194 B.n388 B.n95 163.367
R1195 B.n392 B.n95 163.367
R1196 B.n393 B.n392 163.367
R1197 B.n394 B.n393 163.367
R1198 B.n394 B.n93 163.367
R1199 B.n398 B.n93 163.367
R1200 B.n399 B.n398 163.367
R1201 B.n400 B.n399 163.367
R1202 B.n400 B.n91 163.367
R1203 B.n404 B.n91 163.367
R1204 B.n405 B.n404 163.367
R1205 B.n406 B.n405 163.367
R1206 B.n406 B.n89 163.367
R1207 B.n410 B.n89 163.367
R1208 B.n411 B.n410 163.367
R1209 B.n412 B.n411 163.367
R1210 B.n412 B.n87 163.367
R1211 B.n416 B.n87 163.367
R1212 B.n417 B.n416 163.367
R1213 B.n418 B.n417 163.367
R1214 B.n418 B.n85 163.367
R1215 B.n422 B.n85 163.367
R1216 B.n423 B.n422 163.367
R1217 B.n424 B.n423 163.367
R1218 B.n424 B.n83 163.367
R1219 B.n428 B.n83 163.367
R1220 B.n429 B.n428 163.367
R1221 B.n430 B.n429 163.367
R1222 B.n430 B.n81 163.367
R1223 B.n434 B.n81 163.367
R1224 B.n435 B.n434 163.367
R1225 B.n436 B.n435 163.367
R1226 B.n436 B.n79 163.367
R1227 B.n440 B.n79 163.367
R1228 B.n441 B.n440 163.367
R1229 B.n442 B.n441 163.367
R1230 B.n442 B.n77 163.367
R1231 B.n446 B.n77 163.367
R1232 B.n447 B.n446 163.367
R1233 B.n448 B.n447 163.367
R1234 B.n448 B.n75 163.367
R1235 B.n452 B.n75 163.367
R1236 B.n453 B.n452 163.367
R1237 B.n454 B.n453 163.367
R1238 B.n454 B.n73 163.367
R1239 B.n458 B.n73 163.367
R1240 B.n459 B.n458 163.367
R1241 B.n460 B.n459 163.367
R1242 B.n460 B.n71 163.367
R1243 B.n464 B.n71 163.367
R1244 B.n465 B.n464 163.367
R1245 B.n466 B.n465 163.367
R1246 B.n466 B.n69 163.367
R1247 B.n470 B.n69 163.367
R1248 B.n471 B.n470 163.367
R1249 B.n472 B.n471 163.367
R1250 B.n472 B.n67 163.367
R1251 B.n476 B.n67 163.367
R1252 B.n477 B.n476 163.367
R1253 B.n478 B.n477 163.367
R1254 B.n478 B.n65 163.367
R1255 B.n482 B.n65 163.367
R1256 B.n483 B.n482 163.367
R1257 B.n484 B.n483 163.367
R1258 B.n484 B.n63 163.367
R1259 B.n488 B.n63 163.367
R1260 B.n489 B.n488 163.367
R1261 B.n490 B.n489 163.367
R1262 B.n490 B.n61 163.367
R1263 B.n494 B.n61 163.367
R1264 B.n495 B.n494 163.367
R1265 B.n574 B.n29 163.367
R1266 B.n574 B.n573 163.367
R1267 B.n573 B.n572 163.367
R1268 B.n572 B.n31 163.367
R1269 B.n568 B.n31 163.367
R1270 B.n568 B.n567 163.367
R1271 B.n567 B.n566 163.367
R1272 B.n566 B.n33 163.367
R1273 B.n562 B.n33 163.367
R1274 B.n562 B.n561 163.367
R1275 B.n561 B.n560 163.367
R1276 B.n560 B.n35 163.367
R1277 B.n556 B.n35 163.367
R1278 B.n556 B.n555 163.367
R1279 B.n555 B.n554 163.367
R1280 B.n554 B.n37 163.367
R1281 B.n550 B.n37 163.367
R1282 B.n550 B.n549 163.367
R1283 B.n549 B.n548 163.367
R1284 B.n548 B.n39 163.367
R1285 B.n544 B.n39 163.367
R1286 B.n544 B.n543 163.367
R1287 B.n543 B.n43 163.367
R1288 B.n539 B.n43 163.367
R1289 B.n539 B.n538 163.367
R1290 B.n538 B.n537 163.367
R1291 B.n537 B.n45 163.367
R1292 B.n533 B.n45 163.367
R1293 B.n533 B.n532 163.367
R1294 B.n532 B.n531 163.367
R1295 B.n531 B.n47 163.367
R1296 B.n526 B.n47 163.367
R1297 B.n526 B.n525 163.367
R1298 B.n525 B.n524 163.367
R1299 B.n524 B.n51 163.367
R1300 B.n520 B.n51 163.367
R1301 B.n520 B.n519 163.367
R1302 B.n519 B.n518 163.367
R1303 B.n518 B.n53 163.367
R1304 B.n514 B.n53 163.367
R1305 B.n514 B.n513 163.367
R1306 B.n513 B.n512 163.367
R1307 B.n512 B.n55 163.367
R1308 B.n508 B.n55 163.367
R1309 B.n508 B.n507 163.367
R1310 B.n507 B.n506 163.367
R1311 B.n506 B.n57 163.367
R1312 B.n502 B.n57 163.367
R1313 B.n502 B.n501 163.367
R1314 B.n501 B.n500 163.367
R1315 B.n500 B.n59 163.367
R1316 B.n496 B.n59 163.367
R1317 B.n299 B.n127 59.5399
R1318 B.n134 B.n133 59.5399
R1319 B.n42 B.n41 59.5399
R1320 B.n529 B.n49 59.5399
R1321 B.n127 B.n126 50.2308
R1322 B.n133 B.n132 50.2308
R1323 B.n41 B.n40 50.2308
R1324 B.n49 B.n48 50.2308
R1325 B.n577 B.n576 31.3761
R1326 B.n497 B.n60 31.3761
R1327 B.n331 B.n114 31.3761
R1328 B.n252 B.n251 31.3761
R1329 B B.n659 18.0485
R1330 B.n576 B.n575 10.6151
R1331 B.n575 B.n30 10.6151
R1332 B.n571 B.n30 10.6151
R1333 B.n571 B.n570 10.6151
R1334 B.n570 B.n569 10.6151
R1335 B.n569 B.n32 10.6151
R1336 B.n565 B.n32 10.6151
R1337 B.n565 B.n564 10.6151
R1338 B.n564 B.n563 10.6151
R1339 B.n563 B.n34 10.6151
R1340 B.n559 B.n34 10.6151
R1341 B.n559 B.n558 10.6151
R1342 B.n558 B.n557 10.6151
R1343 B.n557 B.n36 10.6151
R1344 B.n553 B.n36 10.6151
R1345 B.n553 B.n552 10.6151
R1346 B.n552 B.n551 10.6151
R1347 B.n551 B.n38 10.6151
R1348 B.n547 B.n38 10.6151
R1349 B.n547 B.n546 10.6151
R1350 B.n546 B.n545 10.6151
R1351 B.n542 B.n541 10.6151
R1352 B.n541 B.n540 10.6151
R1353 B.n540 B.n44 10.6151
R1354 B.n536 B.n44 10.6151
R1355 B.n536 B.n535 10.6151
R1356 B.n535 B.n534 10.6151
R1357 B.n534 B.n46 10.6151
R1358 B.n530 B.n46 10.6151
R1359 B.n528 B.n527 10.6151
R1360 B.n527 B.n50 10.6151
R1361 B.n523 B.n50 10.6151
R1362 B.n523 B.n522 10.6151
R1363 B.n522 B.n521 10.6151
R1364 B.n521 B.n52 10.6151
R1365 B.n517 B.n52 10.6151
R1366 B.n517 B.n516 10.6151
R1367 B.n516 B.n515 10.6151
R1368 B.n515 B.n54 10.6151
R1369 B.n511 B.n54 10.6151
R1370 B.n511 B.n510 10.6151
R1371 B.n510 B.n509 10.6151
R1372 B.n509 B.n56 10.6151
R1373 B.n505 B.n56 10.6151
R1374 B.n505 B.n504 10.6151
R1375 B.n504 B.n503 10.6151
R1376 B.n503 B.n58 10.6151
R1377 B.n499 B.n58 10.6151
R1378 B.n499 B.n498 10.6151
R1379 B.n498 B.n497 10.6151
R1380 B.n335 B.n114 10.6151
R1381 B.n336 B.n335 10.6151
R1382 B.n337 B.n336 10.6151
R1383 B.n337 B.n112 10.6151
R1384 B.n341 B.n112 10.6151
R1385 B.n342 B.n341 10.6151
R1386 B.n343 B.n342 10.6151
R1387 B.n343 B.n110 10.6151
R1388 B.n347 B.n110 10.6151
R1389 B.n348 B.n347 10.6151
R1390 B.n349 B.n348 10.6151
R1391 B.n349 B.n108 10.6151
R1392 B.n353 B.n108 10.6151
R1393 B.n354 B.n353 10.6151
R1394 B.n355 B.n354 10.6151
R1395 B.n355 B.n106 10.6151
R1396 B.n359 B.n106 10.6151
R1397 B.n360 B.n359 10.6151
R1398 B.n361 B.n360 10.6151
R1399 B.n361 B.n104 10.6151
R1400 B.n365 B.n104 10.6151
R1401 B.n366 B.n365 10.6151
R1402 B.n367 B.n366 10.6151
R1403 B.n367 B.n102 10.6151
R1404 B.n371 B.n102 10.6151
R1405 B.n372 B.n371 10.6151
R1406 B.n373 B.n372 10.6151
R1407 B.n373 B.n100 10.6151
R1408 B.n377 B.n100 10.6151
R1409 B.n378 B.n377 10.6151
R1410 B.n379 B.n378 10.6151
R1411 B.n379 B.n98 10.6151
R1412 B.n383 B.n98 10.6151
R1413 B.n384 B.n383 10.6151
R1414 B.n385 B.n384 10.6151
R1415 B.n385 B.n96 10.6151
R1416 B.n389 B.n96 10.6151
R1417 B.n390 B.n389 10.6151
R1418 B.n391 B.n390 10.6151
R1419 B.n391 B.n94 10.6151
R1420 B.n395 B.n94 10.6151
R1421 B.n396 B.n395 10.6151
R1422 B.n397 B.n396 10.6151
R1423 B.n397 B.n92 10.6151
R1424 B.n401 B.n92 10.6151
R1425 B.n402 B.n401 10.6151
R1426 B.n403 B.n402 10.6151
R1427 B.n403 B.n90 10.6151
R1428 B.n407 B.n90 10.6151
R1429 B.n408 B.n407 10.6151
R1430 B.n409 B.n408 10.6151
R1431 B.n409 B.n88 10.6151
R1432 B.n413 B.n88 10.6151
R1433 B.n414 B.n413 10.6151
R1434 B.n415 B.n414 10.6151
R1435 B.n415 B.n86 10.6151
R1436 B.n419 B.n86 10.6151
R1437 B.n420 B.n419 10.6151
R1438 B.n421 B.n420 10.6151
R1439 B.n421 B.n84 10.6151
R1440 B.n425 B.n84 10.6151
R1441 B.n426 B.n425 10.6151
R1442 B.n427 B.n426 10.6151
R1443 B.n427 B.n82 10.6151
R1444 B.n431 B.n82 10.6151
R1445 B.n432 B.n431 10.6151
R1446 B.n433 B.n432 10.6151
R1447 B.n433 B.n80 10.6151
R1448 B.n437 B.n80 10.6151
R1449 B.n438 B.n437 10.6151
R1450 B.n439 B.n438 10.6151
R1451 B.n439 B.n78 10.6151
R1452 B.n443 B.n78 10.6151
R1453 B.n444 B.n443 10.6151
R1454 B.n445 B.n444 10.6151
R1455 B.n445 B.n76 10.6151
R1456 B.n449 B.n76 10.6151
R1457 B.n450 B.n449 10.6151
R1458 B.n451 B.n450 10.6151
R1459 B.n451 B.n74 10.6151
R1460 B.n455 B.n74 10.6151
R1461 B.n456 B.n455 10.6151
R1462 B.n457 B.n456 10.6151
R1463 B.n457 B.n72 10.6151
R1464 B.n461 B.n72 10.6151
R1465 B.n462 B.n461 10.6151
R1466 B.n463 B.n462 10.6151
R1467 B.n463 B.n70 10.6151
R1468 B.n467 B.n70 10.6151
R1469 B.n468 B.n467 10.6151
R1470 B.n469 B.n468 10.6151
R1471 B.n469 B.n68 10.6151
R1472 B.n473 B.n68 10.6151
R1473 B.n474 B.n473 10.6151
R1474 B.n475 B.n474 10.6151
R1475 B.n475 B.n66 10.6151
R1476 B.n479 B.n66 10.6151
R1477 B.n480 B.n479 10.6151
R1478 B.n481 B.n480 10.6151
R1479 B.n481 B.n64 10.6151
R1480 B.n485 B.n64 10.6151
R1481 B.n486 B.n485 10.6151
R1482 B.n487 B.n486 10.6151
R1483 B.n487 B.n62 10.6151
R1484 B.n491 B.n62 10.6151
R1485 B.n492 B.n491 10.6151
R1486 B.n493 B.n492 10.6151
R1487 B.n493 B.n60 10.6151
R1488 B.n253 B.n252 10.6151
R1489 B.n253 B.n144 10.6151
R1490 B.n257 B.n144 10.6151
R1491 B.n258 B.n257 10.6151
R1492 B.n259 B.n258 10.6151
R1493 B.n259 B.n142 10.6151
R1494 B.n263 B.n142 10.6151
R1495 B.n264 B.n263 10.6151
R1496 B.n265 B.n264 10.6151
R1497 B.n265 B.n140 10.6151
R1498 B.n269 B.n140 10.6151
R1499 B.n270 B.n269 10.6151
R1500 B.n271 B.n270 10.6151
R1501 B.n271 B.n138 10.6151
R1502 B.n275 B.n138 10.6151
R1503 B.n276 B.n275 10.6151
R1504 B.n277 B.n276 10.6151
R1505 B.n277 B.n136 10.6151
R1506 B.n281 B.n136 10.6151
R1507 B.n282 B.n281 10.6151
R1508 B.n283 B.n282 10.6151
R1509 B.n287 B.n286 10.6151
R1510 B.n288 B.n287 10.6151
R1511 B.n288 B.n130 10.6151
R1512 B.n292 B.n130 10.6151
R1513 B.n293 B.n292 10.6151
R1514 B.n294 B.n293 10.6151
R1515 B.n294 B.n128 10.6151
R1516 B.n298 B.n128 10.6151
R1517 B.n301 B.n300 10.6151
R1518 B.n301 B.n124 10.6151
R1519 B.n305 B.n124 10.6151
R1520 B.n306 B.n305 10.6151
R1521 B.n307 B.n306 10.6151
R1522 B.n307 B.n122 10.6151
R1523 B.n311 B.n122 10.6151
R1524 B.n312 B.n311 10.6151
R1525 B.n313 B.n312 10.6151
R1526 B.n313 B.n120 10.6151
R1527 B.n317 B.n120 10.6151
R1528 B.n318 B.n317 10.6151
R1529 B.n319 B.n318 10.6151
R1530 B.n319 B.n118 10.6151
R1531 B.n323 B.n118 10.6151
R1532 B.n324 B.n323 10.6151
R1533 B.n325 B.n324 10.6151
R1534 B.n325 B.n116 10.6151
R1535 B.n329 B.n116 10.6151
R1536 B.n330 B.n329 10.6151
R1537 B.n331 B.n330 10.6151
R1538 B.n251 B.n146 10.6151
R1539 B.n247 B.n146 10.6151
R1540 B.n247 B.n246 10.6151
R1541 B.n246 B.n245 10.6151
R1542 B.n245 B.n148 10.6151
R1543 B.n241 B.n148 10.6151
R1544 B.n241 B.n240 10.6151
R1545 B.n240 B.n239 10.6151
R1546 B.n239 B.n150 10.6151
R1547 B.n235 B.n150 10.6151
R1548 B.n235 B.n234 10.6151
R1549 B.n234 B.n233 10.6151
R1550 B.n233 B.n152 10.6151
R1551 B.n229 B.n152 10.6151
R1552 B.n229 B.n228 10.6151
R1553 B.n228 B.n227 10.6151
R1554 B.n227 B.n154 10.6151
R1555 B.n223 B.n154 10.6151
R1556 B.n223 B.n222 10.6151
R1557 B.n222 B.n221 10.6151
R1558 B.n221 B.n156 10.6151
R1559 B.n217 B.n156 10.6151
R1560 B.n217 B.n216 10.6151
R1561 B.n216 B.n215 10.6151
R1562 B.n215 B.n158 10.6151
R1563 B.n211 B.n158 10.6151
R1564 B.n211 B.n210 10.6151
R1565 B.n210 B.n209 10.6151
R1566 B.n209 B.n160 10.6151
R1567 B.n205 B.n160 10.6151
R1568 B.n205 B.n204 10.6151
R1569 B.n204 B.n203 10.6151
R1570 B.n203 B.n162 10.6151
R1571 B.n199 B.n162 10.6151
R1572 B.n199 B.n198 10.6151
R1573 B.n198 B.n197 10.6151
R1574 B.n197 B.n164 10.6151
R1575 B.n193 B.n164 10.6151
R1576 B.n193 B.n192 10.6151
R1577 B.n192 B.n191 10.6151
R1578 B.n191 B.n166 10.6151
R1579 B.n187 B.n166 10.6151
R1580 B.n187 B.n186 10.6151
R1581 B.n186 B.n185 10.6151
R1582 B.n185 B.n168 10.6151
R1583 B.n181 B.n168 10.6151
R1584 B.n181 B.n180 10.6151
R1585 B.n180 B.n179 10.6151
R1586 B.n179 B.n170 10.6151
R1587 B.n175 B.n170 10.6151
R1588 B.n175 B.n174 10.6151
R1589 B.n174 B.n173 10.6151
R1590 B.n173 B.n0 10.6151
R1591 B.n655 B.n1 10.6151
R1592 B.n655 B.n654 10.6151
R1593 B.n654 B.n653 10.6151
R1594 B.n653 B.n4 10.6151
R1595 B.n649 B.n4 10.6151
R1596 B.n649 B.n648 10.6151
R1597 B.n648 B.n647 10.6151
R1598 B.n647 B.n6 10.6151
R1599 B.n643 B.n6 10.6151
R1600 B.n643 B.n642 10.6151
R1601 B.n642 B.n641 10.6151
R1602 B.n641 B.n8 10.6151
R1603 B.n637 B.n8 10.6151
R1604 B.n637 B.n636 10.6151
R1605 B.n636 B.n635 10.6151
R1606 B.n635 B.n10 10.6151
R1607 B.n631 B.n10 10.6151
R1608 B.n631 B.n630 10.6151
R1609 B.n630 B.n629 10.6151
R1610 B.n629 B.n12 10.6151
R1611 B.n625 B.n12 10.6151
R1612 B.n625 B.n624 10.6151
R1613 B.n624 B.n623 10.6151
R1614 B.n623 B.n14 10.6151
R1615 B.n619 B.n14 10.6151
R1616 B.n619 B.n618 10.6151
R1617 B.n618 B.n617 10.6151
R1618 B.n617 B.n16 10.6151
R1619 B.n613 B.n16 10.6151
R1620 B.n613 B.n612 10.6151
R1621 B.n612 B.n611 10.6151
R1622 B.n611 B.n18 10.6151
R1623 B.n607 B.n18 10.6151
R1624 B.n607 B.n606 10.6151
R1625 B.n606 B.n605 10.6151
R1626 B.n605 B.n20 10.6151
R1627 B.n601 B.n20 10.6151
R1628 B.n601 B.n600 10.6151
R1629 B.n600 B.n599 10.6151
R1630 B.n599 B.n22 10.6151
R1631 B.n595 B.n22 10.6151
R1632 B.n595 B.n594 10.6151
R1633 B.n594 B.n593 10.6151
R1634 B.n593 B.n24 10.6151
R1635 B.n589 B.n24 10.6151
R1636 B.n589 B.n588 10.6151
R1637 B.n588 B.n587 10.6151
R1638 B.n587 B.n26 10.6151
R1639 B.n583 B.n26 10.6151
R1640 B.n583 B.n582 10.6151
R1641 B.n582 B.n581 10.6151
R1642 B.n581 B.n28 10.6151
R1643 B.n577 B.n28 10.6151
R1644 B.n542 B.n42 6.5566
R1645 B.n530 B.n529 6.5566
R1646 B.n286 B.n134 6.5566
R1647 B.n299 B.n298 6.5566
R1648 B.n545 B.n42 4.05904
R1649 B.n529 B.n528 4.05904
R1650 B.n283 B.n134 4.05904
R1651 B.n300 B.n299 4.05904
R1652 B.n659 B.n0 2.81026
R1653 B.n659 B.n1 2.81026
C0 VP VDD1 5.20744f
C1 VDD2 B 1.92431f
C2 VN VDD1 0.152971f
C3 VDD2 w_n4078_n2020# 2.31425f
C4 VP B 2.0502f
C5 VDD1 VTAIL 7.03778f
C6 VN B 1.16105f
C7 VP w_n4078_n2020# 9.03445f
C8 VN w_n4078_n2020# 8.50465f
C9 VTAIL B 2.09693f
C10 VP VDD2 0.544177f
C11 VTAIL w_n4078_n2020# 2.20735f
C12 VDD2 VN 4.82309f
C13 VDD1 B 1.81949f
C14 VDD2 VTAIL 7.08783f
C15 VP VN 6.64776f
C16 VDD1 w_n4078_n2020# 2.18855f
C17 VP VTAIL 5.81819f
C18 VDD2 VDD1 1.95267f
C19 w_n4078_n2020# B 8.09621f
C20 VN VTAIL 5.80399f
C21 VDD2 VSUBS 1.664853f
C22 VDD1 VSUBS 1.598067f
C23 VTAIL VSUBS 0.618251f
C24 VN VSUBS 6.78177f
C25 VP VSUBS 3.29183f
C26 B VSUBS 4.117736f
C27 w_n4078_n2020# VSUBS 0.103108p
C28 B.n0 VSUBS 0.00609f
C29 B.n1 VSUBS 0.00609f
C30 B.n2 VSUBS 0.00963f
C31 B.n3 VSUBS 0.00963f
C32 B.n4 VSUBS 0.00963f
C33 B.n5 VSUBS 0.00963f
C34 B.n6 VSUBS 0.00963f
C35 B.n7 VSUBS 0.00963f
C36 B.n8 VSUBS 0.00963f
C37 B.n9 VSUBS 0.00963f
C38 B.n10 VSUBS 0.00963f
C39 B.n11 VSUBS 0.00963f
C40 B.n12 VSUBS 0.00963f
C41 B.n13 VSUBS 0.00963f
C42 B.n14 VSUBS 0.00963f
C43 B.n15 VSUBS 0.00963f
C44 B.n16 VSUBS 0.00963f
C45 B.n17 VSUBS 0.00963f
C46 B.n18 VSUBS 0.00963f
C47 B.n19 VSUBS 0.00963f
C48 B.n20 VSUBS 0.00963f
C49 B.n21 VSUBS 0.00963f
C50 B.n22 VSUBS 0.00963f
C51 B.n23 VSUBS 0.00963f
C52 B.n24 VSUBS 0.00963f
C53 B.n25 VSUBS 0.00963f
C54 B.n26 VSUBS 0.00963f
C55 B.n27 VSUBS 0.00963f
C56 B.n28 VSUBS 0.00963f
C57 B.n29 VSUBS 0.022255f
C58 B.n30 VSUBS 0.00963f
C59 B.n31 VSUBS 0.00963f
C60 B.n32 VSUBS 0.00963f
C61 B.n33 VSUBS 0.00963f
C62 B.n34 VSUBS 0.00963f
C63 B.n35 VSUBS 0.00963f
C64 B.n36 VSUBS 0.00963f
C65 B.n37 VSUBS 0.00963f
C66 B.n38 VSUBS 0.00963f
C67 B.n39 VSUBS 0.00963f
C68 B.t2 VSUBS 0.105764f
C69 B.t1 VSUBS 0.135377f
C70 B.t0 VSUBS 0.773039f
C71 B.n40 VSUBS 0.23575f
C72 B.n41 VSUBS 0.193834f
C73 B.n42 VSUBS 0.022313f
C74 B.n43 VSUBS 0.00963f
C75 B.n44 VSUBS 0.00963f
C76 B.n45 VSUBS 0.00963f
C77 B.n46 VSUBS 0.00963f
C78 B.n47 VSUBS 0.00963f
C79 B.t5 VSUBS 0.105766f
C80 B.t4 VSUBS 0.135379f
C81 B.t3 VSUBS 0.773039f
C82 B.n48 VSUBS 0.235748f
C83 B.n49 VSUBS 0.193832f
C84 B.n50 VSUBS 0.00963f
C85 B.n51 VSUBS 0.00963f
C86 B.n52 VSUBS 0.00963f
C87 B.n53 VSUBS 0.00963f
C88 B.n54 VSUBS 0.00963f
C89 B.n55 VSUBS 0.00963f
C90 B.n56 VSUBS 0.00963f
C91 B.n57 VSUBS 0.00963f
C92 B.n58 VSUBS 0.00963f
C93 B.n59 VSUBS 0.00963f
C94 B.n60 VSUBS 0.022833f
C95 B.n61 VSUBS 0.00963f
C96 B.n62 VSUBS 0.00963f
C97 B.n63 VSUBS 0.00963f
C98 B.n64 VSUBS 0.00963f
C99 B.n65 VSUBS 0.00963f
C100 B.n66 VSUBS 0.00963f
C101 B.n67 VSUBS 0.00963f
C102 B.n68 VSUBS 0.00963f
C103 B.n69 VSUBS 0.00963f
C104 B.n70 VSUBS 0.00963f
C105 B.n71 VSUBS 0.00963f
C106 B.n72 VSUBS 0.00963f
C107 B.n73 VSUBS 0.00963f
C108 B.n74 VSUBS 0.00963f
C109 B.n75 VSUBS 0.00963f
C110 B.n76 VSUBS 0.00963f
C111 B.n77 VSUBS 0.00963f
C112 B.n78 VSUBS 0.00963f
C113 B.n79 VSUBS 0.00963f
C114 B.n80 VSUBS 0.00963f
C115 B.n81 VSUBS 0.00963f
C116 B.n82 VSUBS 0.00963f
C117 B.n83 VSUBS 0.00963f
C118 B.n84 VSUBS 0.00963f
C119 B.n85 VSUBS 0.00963f
C120 B.n86 VSUBS 0.00963f
C121 B.n87 VSUBS 0.00963f
C122 B.n88 VSUBS 0.00963f
C123 B.n89 VSUBS 0.00963f
C124 B.n90 VSUBS 0.00963f
C125 B.n91 VSUBS 0.00963f
C126 B.n92 VSUBS 0.00963f
C127 B.n93 VSUBS 0.00963f
C128 B.n94 VSUBS 0.00963f
C129 B.n95 VSUBS 0.00963f
C130 B.n96 VSUBS 0.00963f
C131 B.n97 VSUBS 0.00963f
C132 B.n98 VSUBS 0.00963f
C133 B.n99 VSUBS 0.00963f
C134 B.n100 VSUBS 0.00963f
C135 B.n101 VSUBS 0.00963f
C136 B.n102 VSUBS 0.00963f
C137 B.n103 VSUBS 0.00963f
C138 B.n104 VSUBS 0.00963f
C139 B.n105 VSUBS 0.00963f
C140 B.n106 VSUBS 0.00963f
C141 B.n107 VSUBS 0.00963f
C142 B.n108 VSUBS 0.00963f
C143 B.n109 VSUBS 0.00963f
C144 B.n110 VSUBS 0.00963f
C145 B.n111 VSUBS 0.00963f
C146 B.n112 VSUBS 0.00963f
C147 B.n113 VSUBS 0.00963f
C148 B.n114 VSUBS 0.021649f
C149 B.n115 VSUBS 0.00963f
C150 B.n116 VSUBS 0.00963f
C151 B.n117 VSUBS 0.00963f
C152 B.n118 VSUBS 0.00963f
C153 B.n119 VSUBS 0.00963f
C154 B.n120 VSUBS 0.00963f
C155 B.n121 VSUBS 0.00963f
C156 B.n122 VSUBS 0.00963f
C157 B.n123 VSUBS 0.00963f
C158 B.n124 VSUBS 0.00963f
C159 B.n125 VSUBS 0.00963f
C160 B.t7 VSUBS 0.105766f
C161 B.t8 VSUBS 0.135379f
C162 B.t6 VSUBS 0.773039f
C163 B.n126 VSUBS 0.235748f
C164 B.n127 VSUBS 0.193832f
C165 B.n128 VSUBS 0.00963f
C166 B.n129 VSUBS 0.00963f
C167 B.n130 VSUBS 0.00963f
C168 B.n131 VSUBS 0.00963f
C169 B.t10 VSUBS 0.105764f
C170 B.t11 VSUBS 0.135377f
C171 B.t9 VSUBS 0.773039f
C172 B.n132 VSUBS 0.23575f
C173 B.n133 VSUBS 0.193834f
C174 B.n134 VSUBS 0.022313f
C175 B.n135 VSUBS 0.00963f
C176 B.n136 VSUBS 0.00963f
C177 B.n137 VSUBS 0.00963f
C178 B.n138 VSUBS 0.00963f
C179 B.n139 VSUBS 0.00963f
C180 B.n140 VSUBS 0.00963f
C181 B.n141 VSUBS 0.00963f
C182 B.n142 VSUBS 0.00963f
C183 B.n143 VSUBS 0.00963f
C184 B.n144 VSUBS 0.00963f
C185 B.n145 VSUBS 0.022255f
C186 B.n146 VSUBS 0.00963f
C187 B.n147 VSUBS 0.00963f
C188 B.n148 VSUBS 0.00963f
C189 B.n149 VSUBS 0.00963f
C190 B.n150 VSUBS 0.00963f
C191 B.n151 VSUBS 0.00963f
C192 B.n152 VSUBS 0.00963f
C193 B.n153 VSUBS 0.00963f
C194 B.n154 VSUBS 0.00963f
C195 B.n155 VSUBS 0.00963f
C196 B.n156 VSUBS 0.00963f
C197 B.n157 VSUBS 0.00963f
C198 B.n158 VSUBS 0.00963f
C199 B.n159 VSUBS 0.00963f
C200 B.n160 VSUBS 0.00963f
C201 B.n161 VSUBS 0.00963f
C202 B.n162 VSUBS 0.00963f
C203 B.n163 VSUBS 0.00963f
C204 B.n164 VSUBS 0.00963f
C205 B.n165 VSUBS 0.00963f
C206 B.n166 VSUBS 0.00963f
C207 B.n167 VSUBS 0.00963f
C208 B.n168 VSUBS 0.00963f
C209 B.n169 VSUBS 0.00963f
C210 B.n170 VSUBS 0.00963f
C211 B.n171 VSUBS 0.00963f
C212 B.n172 VSUBS 0.00963f
C213 B.n173 VSUBS 0.00963f
C214 B.n174 VSUBS 0.00963f
C215 B.n175 VSUBS 0.00963f
C216 B.n176 VSUBS 0.00963f
C217 B.n177 VSUBS 0.00963f
C218 B.n178 VSUBS 0.00963f
C219 B.n179 VSUBS 0.00963f
C220 B.n180 VSUBS 0.00963f
C221 B.n181 VSUBS 0.00963f
C222 B.n182 VSUBS 0.00963f
C223 B.n183 VSUBS 0.00963f
C224 B.n184 VSUBS 0.00963f
C225 B.n185 VSUBS 0.00963f
C226 B.n186 VSUBS 0.00963f
C227 B.n187 VSUBS 0.00963f
C228 B.n188 VSUBS 0.00963f
C229 B.n189 VSUBS 0.00963f
C230 B.n190 VSUBS 0.00963f
C231 B.n191 VSUBS 0.00963f
C232 B.n192 VSUBS 0.00963f
C233 B.n193 VSUBS 0.00963f
C234 B.n194 VSUBS 0.00963f
C235 B.n195 VSUBS 0.00963f
C236 B.n196 VSUBS 0.00963f
C237 B.n197 VSUBS 0.00963f
C238 B.n198 VSUBS 0.00963f
C239 B.n199 VSUBS 0.00963f
C240 B.n200 VSUBS 0.00963f
C241 B.n201 VSUBS 0.00963f
C242 B.n202 VSUBS 0.00963f
C243 B.n203 VSUBS 0.00963f
C244 B.n204 VSUBS 0.00963f
C245 B.n205 VSUBS 0.00963f
C246 B.n206 VSUBS 0.00963f
C247 B.n207 VSUBS 0.00963f
C248 B.n208 VSUBS 0.00963f
C249 B.n209 VSUBS 0.00963f
C250 B.n210 VSUBS 0.00963f
C251 B.n211 VSUBS 0.00963f
C252 B.n212 VSUBS 0.00963f
C253 B.n213 VSUBS 0.00963f
C254 B.n214 VSUBS 0.00963f
C255 B.n215 VSUBS 0.00963f
C256 B.n216 VSUBS 0.00963f
C257 B.n217 VSUBS 0.00963f
C258 B.n218 VSUBS 0.00963f
C259 B.n219 VSUBS 0.00963f
C260 B.n220 VSUBS 0.00963f
C261 B.n221 VSUBS 0.00963f
C262 B.n222 VSUBS 0.00963f
C263 B.n223 VSUBS 0.00963f
C264 B.n224 VSUBS 0.00963f
C265 B.n225 VSUBS 0.00963f
C266 B.n226 VSUBS 0.00963f
C267 B.n227 VSUBS 0.00963f
C268 B.n228 VSUBS 0.00963f
C269 B.n229 VSUBS 0.00963f
C270 B.n230 VSUBS 0.00963f
C271 B.n231 VSUBS 0.00963f
C272 B.n232 VSUBS 0.00963f
C273 B.n233 VSUBS 0.00963f
C274 B.n234 VSUBS 0.00963f
C275 B.n235 VSUBS 0.00963f
C276 B.n236 VSUBS 0.00963f
C277 B.n237 VSUBS 0.00963f
C278 B.n238 VSUBS 0.00963f
C279 B.n239 VSUBS 0.00963f
C280 B.n240 VSUBS 0.00963f
C281 B.n241 VSUBS 0.00963f
C282 B.n242 VSUBS 0.00963f
C283 B.n243 VSUBS 0.00963f
C284 B.n244 VSUBS 0.00963f
C285 B.n245 VSUBS 0.00963f
C286 B.n246 VSUBS 0.00963f
C287 B.n247 VSUBS 0.00963f
C288 B.n248 VSUBS 0.00963f
C289 B.n249 VSUBS 0.00963f
C290 B.n250 VSUBS 0.021649f
C291 B.n251 VSUBS 0.021649f
C292 B.n252 VSUBS 0.022255f
C293 B.n253 VSUBS 0.00963f
C294 B.n254 VSUBS 0.00963f
C295 B.n255 VSUBS 0.00963f
C296 B.n256 VSUBS 0.00963f
C297 B.n257 VSUBS 0.00963f
C298 B.n258 VSUBS 0.00963f
C299 B.n259 VSUBS 0.00963f
C300 B.n260 VSUBS 0.00963f
C301 B.n261 VSUBS 0.00963f
C302 B.n262 VSUBS 0.00963f
C303 B.n263 VSUBS 0.00963f
C304 B.n264 VSUBS 0.00963f
C305 B.n265 VSUBS 0.00963f
C306 B.n266 VSUBS 0.00963f
C307 B.n267 VSUBS 0.00963f
C308 B.n268 VSUBS 0.00963f
C309 B.n269 VSUBS 0.00963f
C310 B.n270 VSUBS 0.00963f
C311 B.n271 VSUBS 0.00963f
C312 B.n272 VSUBS 0.00963f
C313 B.n273 VSUBS 0.00963f
C314 B.n274 VSUBS 0.00963f
C315 B.n275 VSUBS 0.00963f
C316 B.n276 VSUBS 0.00963f
C317 B.n277 VSUBS 0.00963f
C318 B.n278 VSUBS 0.00963f
C319 B.n279 VSUBS 0.00963f
C320 B.n280 VSUBS 0.00963f
C321 B.n281 VSUBS 0.00963f
C322 B.n282 VSUBS 0.00963f
C323 B.n283 VSUBS 0.006656f
C324 B.n284 VSUBS 0.00963f
C325 B.n285 VSUBS 0.00963f
C326 B.n286 VSUBS 0.007789f
C327 B.n287 VSUBS 0.00963f
C328 B.n288 VSUBS 0.00963f
C329 B.n289 VSUBS 0.00963f
C330 B.n290 VSUBS 0.00963f
C331 B.n291 VSUBS 0.00963f
C332 B.n292 VSUBS 0.00963f
C333 B.n293 VSUBS 0.00963f
C334 B.n294 VSUBS 0.00963f
C335 B.n295 VSUBS 0.00963f
C336 B.n296 VSUBS 0.00963f
C337 B.n297 VSUBS 0.00963f
C338 B.n298 VSUBS 0.007789f
C339 B.n299 VSUBS 0.022313f
C340 B.n300 VSUBS 0.006656f
C341 B.n301 VSUBS 0.00963f
C342 B.n302 VSUBS 0.00963f
C343 B.n303 VSUBS 0.00963f
C344 B.n304 VSUBS 0.00963f
C345 B.n305 VSUBS 0.00963f
C346 B.n306 VSUBS 0.00963f
C347 B.n307 VSUBS 0.00963f
C348 B.n308 VSUBS 0.00963f
C349 B.n309 VSUBS 0.00963f
C350 B.n310 VSUBS 0.00963f
C351 B.n311 VSUBS 0.00963f
C352 B.n312 VSUBS 0.00963f
C353 B.n313 VSUBS 0.00963f
C354 B.n314 VSUBS 0.00963f
C355 B.n315 VSUBS 0.00963f
C356 B.n316 VSUBS 0.00963f
C357 B.n317 VSUBS 0.00963f
C358 B.n318 VSUBS 0.00963f
C359 B.n319 VSUBS 0.00963f
C360 B.n320 VSUBS 0.00963f
C361 B.n321 VSUBS 0.00963f
C362 B.n322 VSUBS 0.00963f
C363 B.n323 VSUBS 0.00963f
C364 B.n324 VSUBS 0.00963f
C365 B.n325 VSUBS 0.00963f
C366 B.n326 VSUBS 0.00963f
C367 B.n327 VSUBS 0.00963f
C368 B.n328 VSUBS 0.00963f
C369 B.n329 VSUBS 0.00963f
C370 B.n330 VSUBS 0.00963f
C371 B.n331 VSUBS 0.022255f
C372 B.n332 VSUBS 0.022255f
C373 B.n333 VSUBS 0.021649f
C374 B.n334 VSUBS 0.00963f
C375 B.n335 VSUBS 0.00963f
C376 B.n336 VSUBS 0.00963f
C377 B.n337 VSUBS 0.00963f
C378 B.n338 VSUBS 0.00963f
C379 B.n339 VSUBS 0.00963f
C380 B.n340 VSUBS 0.00963f
C381 B.n341 VSUBS 0.00963f
C382 B.n342 VSUBS 0.00963f
C383 B.n343 VSUBS 0.00963f
C384 B.n344 VSUBS 0.00963f
C385 B.n345 VSUBS 0.00963f
C386 B.n346 VSUBS 0.00963f
C387 B.n347 VSUBS 0.00963f
C388 B.n348 VSUBS 0.00963f
C389 B.n349 VSUBS 0.00963f
C390 B.n350 VSUBS 0.00963f
C391 B.n351 VSUBS 0.00963f
C392 B.n352 VSUBS 0.00963f
C393 B.n353 VSUBS 0.00963f
C394 B.n354 VSUBS 0.00963f
C395 B.n355 VSUBS 0.00963f
C396 B.n356 VSUBS 0.00963f
C397 B.n357 VSUBS 0.00963f
C398 B.n358 VSUBS 0.00963f
C399 B.n359 VSUBS 0.00963f
C400 B.n360 VSUBS 0.00963f
C401 B.n361 VSUBS 0.00963f
C402 B.n362 VSUBS 0.00963f
C403 B.n363 VSUBS 0.00963f
C404 B.n364 VSUBS 0.00963f
C405 B.n365 VSUBS 0.00963f
C406 B.n366 VSUBS 0.00963f
C407 B.n367 VSUBS 0.00963f
C408 B.n368 VSUBS 0.00963f
C409 B.n369 VSUBS 0.00963f
C410 B.n370 VSUBS 0.00963f
C411 B.n371 VSUBS 0.00963f
C412 B.n372 VSUBS 0.00963f
C413 B.n373 VSUBS 0.00963f
C414 B.n374 VSUBS 0.00963f
C415 B.n375 VSUBS 0.00963f
C416 B.n376 VSUBS 0.00963f
C417 B.n377 VSUBS 0.00963f
C418 B.n378 VSUBS 0.00963f
C419 B.n379 VSUBS 0.00963f
C420 B.n380 VSUBS 0.00963f
C421 B.n381 VSUBS 0.00963f
C422 B.n382 VSUBS 0.00963f
C423 B.n383 VSUBS 0.00963f
C424 B.n384 VSUBS 0.00963f
C425 B.n385 VSUBS 0.00963f
C426 B.n386 VSUBS 0.00963f
C427 B.n387 VSUBS 0.00963f
C428 B.n388 VSUBS 0.00963f
C429 B.n389 VSUBS 0.00963f
C430 B.n390 VSUBS 0.00963f
C431 B.n391 VSUBS 0.00963f
C432 B.n392 VSUBS 0.00963f
C433 B.n393 VSUBS 0.00963f
C434 B.n394 VSUBS 0.00963f
C435 B.n395 VSUBS 0.00963f
C436 B.n396 VSUBS 0.00963f
C437 B.n397 VSUBS 0.00963f
C438 B.n398 VSUBS 0.00963f
C439 B.n399 VSUBS 0.00963f
C440 B.n400 VSUBS 0.00963f
C441 B.n401 VSUBS 0.00963f
C442 B.n402 VSUBS 0.00963f
C443 B.n403 VSUBS 0.00963f
C444 B.n404 VSUBS 0.00963f
C445 B.n405 VSUBS 0.00963f
C446 B.n406 VSUBS 0.00963f
C447 B.n407 VSUBS 0.00963f
C448 B.n408 VSUBS 0.00963f
C449 B.n409 VSUBS 0.00963f
C450 B.n410 VSUBS 0.00963f
C451 B.n411 VSUBS 0.00963f
C452 B.n412 VSUBS 0.00963f
C453 B.n413 VSUBS 0.00963f
C454 B.n414 VSUBS 0.00963f
C455 B.n415 VSUBS 0.00963f
C456 B.n416 VSUBS 0.00963f
C457 B.n417 VSUBS 0.00963f
C458 B.n418 VSUBS 0.00963f
C459 B.n419 VSUBS 0.00963f
C460 B.n420 VSUBS 0.00963f
C461 B.n421 VSUBS 0.00963f
C462 B.n422 VSUBS 0.00963f
C463 B.n423 VSUBS 0.00963f
C464 B.n424 VSUBS 0.00963f
C465 B.n425 VSUBS 0.00963f
C466 B.n426 VSUBS 0.00963f
C467 B.n427 VSUBS 0.00963f
C468 B.n428 VSUBS 0.00963f
C469 B.n429 VSUBS 0.00963f
C470 B.n430 VSUBS 0.00963f
C471 B.n431 VSUBS 0.00963f
C472 B.n432 VSUBS 0.00963f
C473 B.n433 VSUBS 0.00963f
C474 B.n434 VSUBS 0.00963f
C475 B.n435 VSUBS 0.00963f
C476 B.n436 VSUBS 0.00963f
C477 B.n437 VSUBS 0.00963f
C478 B.n438 VSUBS 0.00963f
C479 B.n439 VSUBS 0.00963f
C480 B.n440 VSUBS 0.00963f
C481 B.n441 VSUBS 0.00963f
C482 B.n442 VSUBS 0.00963f
C483 B.n443 VSUBS 0.00963f
C484 B.n444 VSUBS 0.00963f
C485 B.n445 VSUBS 0.00963f
C486 B.n446 VSUBS 0.00963f
C487 B.n447 VSUBS 0.00963f
C488 B.n448 VSUBS 0.00963f
C489 B.n449 VSUBS 0.00963f
C490 B.n450 VSUBS 0.00963f
C491 B.n451 VSUBS 0.00963f
C492 B.n452 VSUBS 0.00963f
C493 B.n453 VSUBS 0.00963f
C494 B.n454 VSUBS 0.00963f
C495 B.n455 VSUBS 0.00963f
C496 B.n456 VSUBS 0.00963f
C497 B.n457 VSUBS 0.00963f
C498 B.n458 VSUBS 0.00963f
C499 B.n459 VSUBS 0.00963f
C500 B.n460 VSUBS 0.00963f
C501 B.n461 VSUBS 0.00963f
C502 B.n462 VSUBS 0.00963f
C503 B.n463 VSUBS 0.00963f
C504 B.n464 VSUBS 0.00963f
C505 B.n465 VSUBS 0.00963f
C506 B.n466 VSUBS 0.00963f
C507 B.n467 VSUBS 0.00963f
C508 B.n468 VSUBS 0.00963f
C509 B.n469 VSUBS 0.00963f
C510 B.n470 VSUBS 0.00963f
C511 B.n471 VSUBS 0.00963f
C512 B.n472 VSUBS 0.00963f
C513 B.n473 VSUBS 0.00963f
C514 B.n474 VSUBS 0.00963f
C515 B.n475 VSUBS 0.00963f
C516 B.n476 VSUBS 0.00963f
C517 B.n477 VSUBS 0.00963f
C518 B.n478 VSUBS 0.00963f
C519 B.n479 VSUBS 0.00963f
C520 B.n480 VSUBS 0.00963f
C521 B.n481 VSUBS 0.00963f
C522 B.n482 VSUBS 0.00963f
C523 B.n483 VSUBS 0.00963f
C524 B.n484 VSUBS 0.00963f
C525 B.n485 VSUBS 0.00963f
C526 B.n486 VSUBS 0.00963f
C527 B.n487 VSUBS 0.00963f
C528 B.n488 VSUBS 0.00963f
C529 B.n489 VSUBS 0.00963f
C530 B.n490 VSUBS 0.00963f
C531 B.n491 VSUBS 0.00963f
C532 B.n492 VSUBS 0.00963f
C533 B.n493 VSUBS 0.00963f
C534 B.n494 VSUBS 0.00963f
C535 B.n495 VSUBS 0.021649f
C536 B.n496 VSUBS 0.022255f
C537 B.n497 VSUBS 0.021071f
C538 B.n498 VSUBS 0.00963f
C539 B.n499 VSUBS 0.00963f
C540 B.n500 VSUBS 0.00963f
C541 B.n501 VSUBS 0.00963f
C542 B.n502 VSUBS 0.00963f
C543 B.n503 VSUBS 0.00963f
C544 B.n504 VSUBS 0.00963f
C545 B.n505 VSUBS 0.00963f
C546 B.n506 VSUBS 0.00963f
C547 B.n507 VSUBS 0.00963f
C548 B.n508 VSUBS 0.00963f
C549 B.n509 VSUBS 0.00963f
C550 B.n510 VSUBS 0.00963f
C551 B.n511 VSUBS 0.00963f
C552 B.n512 VSUBS 0.00963f
C553 B.n513 VSUBS 0.00963f
C554 B.n514 VSUBS 0.00963f
C555 B.n515 VSUBS 0.00963f
C556 B.n516 VSUBS 0.00963f
C557 B.n517 VSUBS 0.00963f
C558 B.n518 VSUBS 0.00963f
C559 B.n519 VSUBS 0.00963f
C560 B.n520 VSUBS 0.00963f
C561 B.n521 VSUBS 0.00963f
C562 B.n522 VSUBS 0.00963f
C563 B.n523 VSUBS 0.00963f
C564 B.n524 VSUBS 0.00963f
C565 B.n525 VSUBS 0.00963f
C566 B.n526 VSUBS 0.00963f
C567 B.n527 VSUBS 0.00963f
C568 B.n528 VSUBS 0.006656f
C569 B.n529 VSUBS 0.022313f
C570 B.n530 VSUBS 0.007789f
C571 B.n531 VSUBS 0.00963f
C572 B.n532 VSUBS 0.00963f
C573 B.n533 VSUBS 0.00963f
C574 B.n534 VSUBS 0.00963f
C575 B.n535 VSUBS 0.00963f
C576 B.n536 VSUBS 0.00963f
C577 B.n537 VSUBS 0.00963f
C578 B.n538 VSUBS 0.00963f
C579 B.n539 VSUBS 0.00963f
C580 B.n540 VSUBS 0.00963f
C581 B.n541 VSUBS 0.00963f
C582 B.n542 VSUBS 0.007789f
C583 B.n543 VSUBS 0.00963f
C584 B.n544 VSUBS 0.00963f
C585 B.n545 VSUBS 0.006656f
C586 B.n546 VSUBS 0.00963f
C587 B.n547 VSUBS 0.00963f
C588 B.n548 VSUBS 0.00963f
C589 B.n549 VSUBS 0.00963f
C590 B.n550 VSUBS 0.00963f
C591 B.n551 VSUBS 0.00963f
C592 B.n552 VSUBS 0.00963f
C593 B.n553 VSUBS 0.00963f
C594 B.n554 VSUBS 0.00963f
C595 B.n555 VSUBS 0.00963f
C596 B.n556 VSUBS 0.00963f
C597 B.n557 VSUBS 0.00963f
C598 B.n558 VSUBS 0.00963f
C599 B.n559 VSUBS 0.00963f
C600 B.n560 VSUBS 0.00963f
C601 B.n561 VSUBS 0.00963f
C602 B.n562 VSUBS 0.00963f
C603 B.n563 VSUBS 0.00963f
C604 B.n564 VSUBS 0.00963f
C605 B.n565 VSUBS 0.00963f
C606 B.n566 VSUBS 0.00963f
C607 B.n567 VSUBS 0.00963f
C608 B.n568 VSUBS 0.00963f
C609 B.n569 VSUBS 0.00963f
C610 B.n570 VSUBS 0.00963f
C611 B.n571 VSUBS 0.00963f
C612 B.n572 VSUBS 0.00963f
C613 B.n573 VSUBS 0.00963f
C614 B.n574 VSUBS 0.00963f
C615 B.n575 VSUBS 0.00963f
C616 B.n576 VSUBS 0.022255f
C617 B.n577 VSUBS 0.021649f
C618 B.n578 VSUBS 0.021649f
C619 B.n579 VSUBS 0.00963f
C620 B.n580 VSUBS 0.00963f
C621 B.n581 VSUBS 0.00963f
C622 B.n582 VSUBS 0.00963f
C623 B.n583 VSUBS 0.00963f
C624 B.n584 VSUBS 0.00963f
C625 B.n585 VSUBS 0.00963f
C626 B.n586 VSUBS 0.00963f
C627 B.n587 VSUBS 0.00963f
C628 B.n588 VSUBS 0.00963f
C629 B.n589 VSUBS 0.00963f
C630 B.n590 VSUBS 0.00963f
C631 B.n591 VSUBS 0.00963f
C632 B.n592 VSUBS 0.00963f
C633 B.n593 VSUBS 0.00963f
C634 B.n594 VSUBS 0.00963f
C635 B.n595 VSUBS 0.00963f
C636 B.n596 VSUBS 0.00963f
C637 B.n597 VSUBS 0.00963f
C638 B.n598 VSUBS 0.00963f
C639 B.n599 VSUBS 0.00963f
C640 B.n600 VSUBS 0.00963f
C641 B.n601 VSUBS 0.00963f
C642 B.n602 VSUBS 0.00963f
C643 B.n603 VSUBS 0.00963f
C644 B.n604 VSUBS 0.00963f
C645 B.n605 VSUBS 0.00963f
C646 B.n606 VSUBS 0.00963f
C647 B.n607 VSUBS 0.00963f
C648 B.n608 VSUBS 0.00963f
C649 B.n609 VSUBS 0.00963f
C650 B.n610 VSUBS 0.00963f
C651 B.n611 VSUBS 0.00963f
C652 B.n612 VSUBS 0.00963f
C653 B.n613 VSUBS 0.00963f
C654 B.n614 VSUBS 0.00963f
C655 B.n615 VSUBS 0.00963f
C656 B.n616 VSUBS 0.00963f
C657 B.n617 VSUBS 0.00963f
C658 B.n618 VSUBS 0.00963f
C659 B.n619 VSUBS 0.00963f
C660 B.n620 VSUBS 0.00963f
C661 B.n621 VSUBS 0.00963f
C662 B.n622 VSUBS 0.00963f
C663 B.n623 VSUBS 0.00963f
C664 B.n624 VSUBS 0.00963f
C665 B.n625 VSUBS 0.00963f
C666 B.n626 VSUBS 0.00963f
C667 B.n627 VSUBS 0.00963f
C668 B.n628 VSUBS 0.00963f
C669 B.n629 VSUBS 0.00963f
C670 B.n630 VSUBS 0.00963f
C671 B.n631 VSUBS 0.00963f
C672 B.n632 VSUBS 0.00963f
C673 B.n633 VSUBS 0.00963f
C674 B.n634 VSUBS 0.00963f
C675 B.n635 VSUBS 0.00963f
C676 B.n636 VSUBS 0.00963f
C677 B.n637 VSUBS 0.00963f
C678 B.n638 VSUBS 0.00963f
C679 B.n639 VSUBS 0.00963f
C680 B.n640 VSUBS 0.00963f
C681 B.n641 VSUBS 0.00963f
C682 B.n642 VSUBS 0.00963f
C683 B.n643 VSUBS 0.00963f
C684 B.n644 VSUBS 0.00963f
C685 B.n645 VSUBS 0.00963f
C686 B.n646 VSUBS 0.00963f
C687 B.n647 VSUBS 0.00963f
C688 B.n648 VSUBS 0.00963f
C689 B.n649 VSUBS 0.00963f
C690 B.n650 VSUBS 0.00963f
C691 B.n651 VSUBS 0.00963f
C692 B.n652 VSUBS 0.00963f
C693 B.n653 VSUBS 0.00963f
C694 B.n654 VSUBS 0.00963f
C695 B.n655 VSUBS 0.00963f
C696 B.n656 VSUBS 0.00963f
C697 B.n657 VSUBS 0.00963f
C698 B.n658 VSUBS 0.00963f
C699 B.n659 VSUBS 0.021807f
C700 VDD2.n0 VSUBS 0.028815f
C701 VDD2.n1 VSUBS 0.026951f
C702 VDD2.n2 VSUBS 0.014482f
C703 VDD2.n3 VSUBS 0.03423f
C704 VDD2.n4 VSUBS 0.015334f
C705 VDD2.n5 VSUBS 0.026951f
C706 VDD2.n6 VSUBS 0.014482f
C707 VDD2.n7 VSUBS 0.025673f
C708 VDD2.n8 VSUBS 0.021743f
C709 VDD2.t0 VSUBS 0.07376f
C710 VDD2.n9 VSUBS 0.113564f
C711 VDD2.n10 VSUBS 0.527065f
C712 VDD2.n11 VSUBS 0.014482f
C713 VDD2.n12 VSUBS 0.015334f
C714 VDD2.n13 VSUBS 0.03423f
C715 VDD2.n14 VSUBS 0.03423f
C716 VDD2.n15 VSUBS 0.015334f
C717 VDD2.n16 VSUBS 0.014482f
C718 VDD2.n17 VSUBS 0.026951f
C719 VDD2.n18 VSUBS 0.026951f
C720 VDD2.n19 VSUBS 0.014482f
C721 VDD2.n20 VSUBS 0.015334f
C722 VDD2.n21 VSUBS 0.03423f
C723 VDD2.n22 VSUBS 0.080149f
C724 VDD2.n23 VSUBS 0.015334f
C725 VDD2.n24 VSUBS 0.014482f
C726 VDD2.n25 VSUBS 0.061559f
C727 VDD2.n26 VSUBS 0.069581f
C728 VDD2.t1 VSUBS 0.112023f
C729 VDD2.t2 VSUBS 0.112023f
C730 VDD2.n27 VSUBS 0.714005f
C731 VDD2.n28 VSUBS 0.893857f
C732 VDD2.t6 VSUBS 0.112023f
C733 VDD2.t9 VSUBS 0.112023f
C734 VDD2.n29 VSUBS 0.726593f
C735 VDD2.n30 VSUBS 2.70087f
C736 VDD2.n31 VSUBS 0.028815f
C737 VDD2.n32 VSUBS 0.026951f
C738 VDD2.n33 VSUBS 0.014482f
C739 VDD2.n34 VSUBS 0.03423f
C740 VDD2.n35 VSUBS 0.015334f
C741 VDD2.n36 VSUBS 0.026951f
C742 VDD2.n37 VSUBS 0.014482f
C743 VDD2.n38 VSUBS 0.025673f
C744 VDD2.n39 VSUBS 0.021743f
C745 VDD2.t7 VSUBS 0.07376f
C746 VDD2.n40 VSUBS 0.113564f
C747 VDD2.n41 VSUBS 0.527065f
C748 VDD2.n42 VSUBS 0.014482f
C749 VDD2.n43 VSUBS 0.015334f
C750 VDD2.n44 VSUBS 0.03423f
C751 VDD2.n45 VSUBS 0.03423f
C752 VDD2.n46 VSUBS 0.015334f
C753 VDD2.n47 VSUBS 0.014482f
C754 VDD2.n48 VSUBS 0.026951f
C755 VDD2.n49 VSUBS 0.026951f
C756 VDD2.n50 VSUBS 0.014482f
C757 VDD2.n51 VSUBS 0.015334f
C758 VDD2.n52 VSUBS 0.03423f
C759 VDD2.n53 VSUBS 0.080149f
C760 VDD2.n54 VSUBS 0.015334f
C761 VDD2.n55 VSUBS 0.014482f
C762 VDD2.n56 VSUBS 0.061559f
C763 VDD2.n57 VSUBS 0.058778f
C764 VDD2.n58 VSUBS 2.40348f
C765 VDD2.t4 VSUBS 0.112023f
C766 VDD2.t3 VSUBS 0.112023f
C767 VDD2.n59 VSUBS 0.714009f
C768 VDD2.n60 VSUBS 0.667906f
C769 VDD2.t8 VSUBS 0.112023f
C770 VDD2.t5 VSUBS 0.112023f
C771 VDD2.n61 VSUBS 0.726561f
C772 VN.n0 VSUBS 0.05166f
C773 VN.t0 VSUBS 1.22273f
C774 VN.n1 VSUBS 0.038794f
C775 VN.n2 VSUBS 0.039186f
C776 VN.t3 VSUBS 1.22273f
C777 VN.n3 VSUBS 0.072666f
C778 VN.n4 VSUBS 0.039186f
C779 VN.t7 VSUBS 1.22273f
C780 VN.n5 VSUBS 0.50782f
C781 VN.n6 VSUBS 0.039186f
C782 VN.n7 VSUBS 0.072666f
C783 VN.t9 VSUBS 1.46183f
C784 VN.n8 VSUBS 0.564296f
C785 VN.t8 VSUBS 1.22273f
C786 VN.n9 VSUBS 0.563609f
C787 VN.n10 VSUBS 0.04325f
C788 VN.n11 VSUBS 0.334973f
C789 VN.n12 VSUBS 0.039186f
C790 VN.n13 VSUBS 0.039186f
C791 VN.n14 VSUBS 0.052084f
C792 VN.n15 VSUBS 0.061841f
C793 VN.n16 VSUBS 0.072666f
C794 VN.n17 VSUBS 0.039186f
C795 VN.n18 VSUBS 0.039186f
C796 VN.n19 VSUBS 0.039186f
C797 VN.n20 VSUBS 0.072666f
C798 VN.n21 VSUBS 0.061841f
C799 VN.n22 VSUBS 0.052084f
C800 VN.n23 VSUBS 0.039186f
C801 VN.n24 VSUBS 0.039186f
C802 VN.n25 VSUBS 0.039186f
C803 VN.n26 VSUBS 0.04325f
C804 VN.n27 VSUBS 0.471027f
C805 VN.n28 VSUBS 0.066209f
C806 VN.n29 VSUBS 0.070409f
C807 VN.n30 VSUBS 0.039186f
C808 VN.n31 VSUBS 0.039186f
C809 VN.n32 VSUBS 0.039186f
C810 VN.n33 VSUBS 0.077389f
C811 VN.n34 VSUBS 0.049707f
C812 VN.n35 VSUBS 0.581212f
C813 VN.n36 VSUBS 0.060548f
C814 VN.n37 VSUBS 0.05166f
C815 VN.t2 VSUBS 1.22273f
C816 VN.n38 VSUBS 0.038794f
C817 VN.n39 VSUBS 0.039186f
C818 VN.t5 VSUBS 1.22273f
C819 VN.n40 VSUBS 0.072666f
C820 VN.n41 VSUBS 0.039186f
C821 VN.t6 VSUBS 1.22273f
C822 VN.n42 VSUBS 0.50782f
C823 VN.n43 VSUBS 0.039186f
C824 VN.n44 VSUBS 0.072666f
C825 VN.t4 VSUBS 1.46183f
C826 VN.n45 VSUBS 0.564296f
C827 VN.t1 VSUBS 1.22273f
C828 VN.n46 VSUBS 0.563609f
C829 VN.n47 VSUBS 0.04325f
C830 VN.n48 VSUBS 0.334973f
C831 VN.n49 VSUBS 0.039186f
C832 VN.n50 VSUBS 0.039186f
C833 VN.n51 VSUBS 0.052084f
C834 VN.n52 VSUBS 0.061841f
C835 VN.n53 VSUBS 0.072666f
C836 VN.n54 VSUBS 0.039186f
C837 VN.n55 VSUBS 0.039186f
C838 VN.n56 VSUBS 0.039186f
C839 VN.n57 VSUBS 0.072666f
C840 VN.n58 VSUBS 0.061841f
C841 VN.n59 VSUBS 0.052084f
C842 VN.n60 VSUBS 0.039186f
C843 VN.n61 VSUBS 0.039186f
C844 VN.n62 VSUBS 0.039186f
C845 VN.n63 VSUBS 0.04325f
C846 VN.n64 VSUBS 0.471027f
C847 VN.n65 VSUBS 0.066209f
C848 VN.n66 VSUBS 0.070409f
C849 VN.n67 VSUBS 0.039186f
C850 VN.n68 VSUBS 0.039186f
C851 VN.n69 VSUBS 0.039186f
C852 VN.n70 VSUBS 0.077389f
C853 VN.n71 VSUBS 0.049707f
C854 VN.n72 VSUBS 0.581212f
C855 VN.n73 VSUBS 1.945f
C856 VTAIL.t3 VSUBS 0.139767f
C857 VTAIL.t2 VSUBS 0.139767f
C858 VTAIL.n0 VSUBS 0.783151f
C859 VTAIL.n1 VSUBS 0.946216f
C860 VTAIL.n2 VSUBS 0.035951f
C861 VTAIL.n3 VSUBS 0.033625f
C862 VTAIL.n4 VSUBS 0.018069f
C863 VTAIL.n5 VSUBS 0.042708f
C864 VTAIL.n6 VSUBS 0.019132f
C865 VTAIL.n7 VSUBS 0.033625f
C866 VTAIL.n8 VSUBS 0.018069f
C867 VTAIL.n9 VSUBS 0.032031f
C868 VTAIL.n10 VSUBS 0.027128f
C869 VTAIL.t11 VSUBS 0.092028f
C870 VTAIL.n11 VSUBS 0.14169f
C871 VTAIL.n12 VSUBS 0.657601f
C872 VTAIL.n13 VSUBS 0.018069f
C873 VTAIL.n14 VSUBS 0.019132f
C874 VTAIL.n15 VSUBS 0.042708f
C875 VTAIL.n16 VSUBS 0.042708f
C876 VTAIL.n17 VSUBS 0.019132f
C877 VTAIL.n18 VSUBS 0.018069f
C878 VTAIL.n19 VSUBS 0.033625f
C879 VTAIL.n20 VSUBS 0.033625f
C880 VTAIL.n21 VSUBS 0.018069f
C881 VTAIL.n22 VSUBS 0.019132f
C882 VTAIL.n23 VSUBS 0.042708f
C883 VTAIL.n24 VSUBS 0.099999f
C884 VTAIL.n25 VSUBS 0.019132f
C885 VTAIL.n26 VSUBS 0.018069f
C886 VTAIL.n27 VSUBS 0.076804f
C887 VTAIL.n28 VSUBS 0.05011f
C888 VTAIL.n29 VSUBS 0.441978f
C889 VTAIL.t16 VSUBS 0.139767f
C890 VTAIL.t15 VSUBS 0.139767f
C891 VTAIL.n30 VSUBS 0.783151f
C892 VTAIL.n31 VSUBS 1.07044f
C893 VTAIL.t12 VSUBS 0.139767f
C894 VTAIL.t10 VSUBS 0.139767f
C895 VTAIL.n32 VSUBS 0.783151f
C896 VTAIL.n33 VSUBS 2.26042f
C897 VTAIL.t5 VSUBS 0.139767f
C898 VTAIL.t0 VSUBS 0.139767f
C899 VTAIL.n34 VSUBS 0.783157f
C900 VTAIL.n35 VSUBS 2.26041f
C901 VTAIL.t7 VSUBS 0.139767f
C902 VTAIL.t4 VSUBS 0.139767f
C903 VTAIL.n36 VSUBS 0.783157f
C904 VTAIL.n37 VSUBS 1.07044f
C905 VTAIL.n38 VSUBS 0.035951f
C906 VTAIL.n39 VSUBS 0.033625f
C907 VTAIL.n40 VSUBS 0.018069f
C908 VTAIL.n41 VSUBS 0.042708f
C909 VTAIL.n42 VSUBS 0.019132f
C910 VTAIL.n43 VSUBS 0.033625f
C911 VTAIL.n44 VSUBS 0.018069f
C912 VTAIL.n45 VSUBS 0.032031f
C913 VTAIL.n46 VSUBS 0.027128f
C914 VTAIL.t8 VSUBS 0.092028f
C915 VTAIL.n47 VSUBS 0.14169f
C916 VTAIL.n48 VSUBS 0.657601f
C917 VTAIL.n49 VSUBS 0.018069f
C918 VTAIL.n50 VSUBS 0.019132f
C919 VTAIL.n51 VSUBS 0.042708f
C920 VTAIL.n52 VSUBS 0.042708f
C921 VTAIL.n53 VSUBS 0.019132f
C922 VTAIL.n54 VSUBS 0.018069f
C923 VTAIL.n55 VSUBS 0.033625f
C924 VTAIL.n56 VSUBS 0.033625f
C925 VTAIL.n57 VSUBS 0.018069f
C926 VTAIL.n58 VSUBS 0.019132f
C927 VTAIL.n59 VSUBS 0.042708f
C928 VTAIL.n60 VSUBS 0.099999f
C929 VTAIL.n61 VSUBS 0.019132f
C930 VTAIL.n62 VSUBS 0.018069f
C931 VTAIL.n63 VSUBS 0.076804f
C932 VTAIL.n64 VSUBS 0.05011f
C933 VTAIL.n65 VSUBS 0.441978f
C934 VTAIL.t17 VSUBS 0.139767f
C935 VTAIL.t19 VSUBS 0.139767f
C936 VTAIL.n66 VSUBS 0.783157f
C937 VTAIL.n67 VSUBS 1.00038f
C938 VTAIL.t14 VSUBS 0.139767f
C939 VTAIL.t18 VSUBS 0.139767f
C940 VTAIL.n68 VSUBS 0.783157f
C941 VTAIL.n69 VSUBS 1.07044f
C942 VTAIL.n70 VSUBS 0.035951f
C943 VTAIL.n71 VSUBS 0.033625f
C944 VTAIL.n72 VSUBS 0.018069f
C945 VTAIL.n73 VSUBS 0.042708f
C946 VTAIL.n74 VSUBS 0.019132f
C947 VTAIL.n75 VSUBS 0.033625f
C948 VTAIL.n76 VSUBS 0.018069f
C949 VTAIL.n77 VSUBS 0.032031f
C950 VTAIL.n78 VSUBS 0.027128f
C951 VTAIL.t13 VSUBS 0.092028f
C952 VTAIL.n79 VSUBS 0.14169f
C953 VTAIL.n80 VSUBS 0.657601f
C954 VTAIL.n81 VSUBS 0.018069f
C955 VTAIL.n82 VSUBS 0.019132f
C956 VTAIL.n83 VSUBS 0.042708f
C957 VTAIL.n84 VSUBS 0.042708f
C958 VTAIL.n85 VSUBS 0.019132f
C959 VTAIL.n86 VSUBS 0.018069f
C960 VTAIL.n87 VSUBS 0.033625f
C961 VTAIL.n88 VSUBS 0.033625f
C962 VTAIL.n89 VSUBS 0.018069f
C963 VTAIL.n90 VSUBS 0.019132f
C964 VTAIL.n91 VSUBS 0.042708f
C965 VTAIL.n92 VSUBS 0.099999f
C966 VTAIL.n93 VSUBS 0.019132f
C967 VTAIL.n94 VSUBS 0.018069f
C968 VTAIL.n95 VSUBS 0.076804f
C969 VTAIL.n96 VSUBS 0.05011f
C970 VTAIL.n97 VSUBS 1.46009f
C971 VTAIL.n98 VSUBS 0.035951f
C972 VTAIL.n99 VSUBS 0.033625f
C973 VTAIL.n100 VSUBS 0.018069f
C974 VTAIL.n101 VSUBS 0.042708f
C975 VTAIL.n102 VSUBS 0.019132f
C976 VTAIL.n103 VSUBS 0.033625f
C977 VTAIL.n104 VSUBS 0.018069f
C978 VTAIL.n105 VSUBS 0.032031f
C979 VTAIL.n106 VSUBS 0.027128f
C980 VTAIL.t9 VSUBS 0.092028f
C981 VTAIL.n107 VSUBS 0.14169f
C982 VTAIL.n108 VSUBS 0.657601f
C983 VTAIL.n109 VSUBS 0.018069f
C984 VTAIL.n110 VSUBS 0.019132f
C985 VTAIL.n111 VSUBS 0.042708f
C986 VTAIL.n112 VSUBS 0.042708f
C987 VTAIL.n113 VSUBS 0.019132f
C988 VTAIL.n114 VSUBS 0.018069f
C989 VTAIL.n115 VSUBS 0.033625f
C990 VTAIL.n116 VSUBS 0.033625f
C991 VTAIL.n117 VSUBS 0.018069f
C992 VTAIL.n118 VSUBS 0.019132f
C993 VTAIL.n119 VSUBS 0.042708f
C994 VTAIL.n120 VSUBS 0.099999f
C995 VTAIL.n121 VSUBS 0.019132f
C996 VTAIL.n122 VSUBS 0.018069f
C997 VTAIL.n123 VSUBS 0.076804f
C998 VTAIL.n124 VSUBS 0.05011f
C999 VTAIL.n125 VSUBS 1.46009f
C1000 VTAIL.t1 VSUBS 0.139767f
C1001 VTAIL.t6 VSUBS 0.139767f
C1002 VTAIL.n126 VSUBS 0.783151f
C1003 VTAIL.n127 VSUBS 0.882701f
C1004 VDD1.n0 VSUBS 0.029017f
C1005 VDD1.n1 VSUBS 0.02714f
C1006 VDD1.n2 VSUBS 0.014584f
C1007 VDD1.n3 VSUBS 0.034471f
C1008 VDD1.n4 VSUBS 0.015442f
C1009 VDD1.n5 VSUBS 0.02714f
C1010 VDD1.n6 VSUBS 0.014584f
C1011 VDD1.n7 VSUBS 0.025853f
C1012 VDD1.n8 VSUBS 0.021896f
C1013 VDD1.t7 VSUBS 0.074279f
C1014 VDD1.n9 VSUBS 0.114362f
C1015 VDD1.n10 VSUBS 0.530768f
C1016 VDD1.n11 VSUBS 0.014584f
C1017 VDD1.n12 VSUBS 0.015442f
C1018 VDD1.n13 VSUBS 0.034471f
C1019 VDD1.n14 VSUBS 0.034471f
C1020 VDD1.n15 VSUBS 0.015442f
C1021 VDD1.n16 VSUBS 0.014584f
C1022 VDD1.n17 VSUBS 0.02714f
C1023 VDD1.n18 VSUBS 0.02714f
C1024 VDD1.n19 VSUBS 0.014584f
C1025 VDD1.n20 VSUBS 0.015442f
C1026 VDD1.n21 VSUBS 0.034471f
C1027 VDD1.n22 VSUBS 0.080712f
C1028 VDD1.n23 VSUBS 0.015442f
C1029 VDD1.n24 VSUBS 0.014584f
C1030 VDD1.n25 VSUBS 0.061991f
C1031 VDD1.n26 VSUBS 0.07007f
C1032 VDD1.t3 VSUBS 0.11281f
C1033 VDD1.t4 VSUBS 0.11281f
C1034 VDD1.n27 VSUBS 0.719025f
C1035 VDD1.n28 VSUBS 0.90881f
C1036 VDD1.n29 VSUBS 0.029017f
C1037 VDD1.n30 VSUBS 0.02714f
C1038 VDD1.n31 VSUBS 0.014584f
C1039 VDD1.n32 VSUBS 0.034471f
C1040 VDD1.n33 VSUBS 0.015442f
C1041 VDD1.n34 VSUBS 0.02714f
C1042 VDD1.n35 VSUBS 0.014584f
C1043 VDD1.n36 VSUBS 0.025853f
C1044 VDD1.n37 VSUBS 0.021896f
C1045 VDD1.t1 VSUBS 0.074279f
C1046 VDD1.n38 VSUBS 0.114362f
C1047 VDD1.n39 VSUBS 0.530768f
C1048 VDD1.n40 VSUBS 0.014584f
C1049 VDD1.n41 VSUBS 0.015442f
C1050 VDD1.n42 VSUBS 0.034471f
C1051 VDD1.n43 VSUBS 0.034471f
C1052 VDD1.n44 VSUBS 0.015442f
C1053 VDD1.n45 VSUBS 0.014584f
C1054 VDD1.n46 VSUBS 0.02714f
C1055 VDD1.n47 VSUBS 0.02714f
C1056 VDD1.n48 VSUBS 0.014584f
C1057 VDD1.n49 VSUBS 0.015442f
C1058 VDD1.n50 VSUBS 0.034471f
C1059 VDD1.n51 VSUBS 0.080712f
C1060 VDD1.n52 VSUBS 0.015442f
C1061 VDD1.n53 VSUBS 0.014584f
C1062 VDD1.n54 VSUBS 0.061991f
C1063 VDD1.n55 VSUBS 0.07007f
C1064 VDD1.t0 VSUBS 0.11281f
C1065 VDD1.t6 VSUBS 0.11281f
C1066 VDD1.n56 VSUBS 0.719021f
C1067 VDD1.n57 VSUBS 0.900136f
C1068 VDD1.t9 VSUBS 0.11281f
C1069 VDD1.t2 VSUBS 0.11281f
C1070 VDD1.n58 VSUBS 0.731698f
C1071 VDD1.n59 VSUBS 2.84006f
C1072 VDD1.t8 VSUBS 0.11281f
C1073 VDD1.t5 VSUBS 0.11281f
C1074 VDD1.n60 VSUBS 0.719021f
C1075 VDD1.n61 VSUBS 2.92428f
C1076 VP.n0 VSUBS 0.057814f
C1077 VP.t8 VSUBS 1.3684f
C1078 VP.n1 VSUBS 0.043416f
C1079 VP.n2 VSUBS 0.043854f
C1080 VP.t4 VSUBS 1.3684f
C1081 VP.n3 VSUBS 0.081323f
C1082 VP.n4 VSUBS 0.043854f
C1083 VP.t3 VSUBS 1.3684f
C1084 VP.n5 VSUBS 0.568317f
C1085 VP.n6 VSUBS 0.043854f
C1086 VP.n7 VSUBS 0.081323f
C1087 VP.n8 VSUBS 0.043854f
C1088 VP.t9 VSUBS 1.3684f
C1089 VP.n9 VSUBS 0.043416f
C1090 VP.n10 VSUBS 0.057814f
C1091 VP.t7 VSUBS 1.3684f
C1092 VP.n11 VSUBS 0.057814f
C1093 VP.t6 VSUBS 1.3684f
C1094 VP.n12 VSUBS 0.043416f
C1095 VP.n13 VSUBS 0.043854f
C1096 VP.t1 VSUBS 1.3684f
C1097 VP.n14 VSUBS 0.081323f
C1098 VP.n15 VSUBS 0.043854f
C1099 VP.t5 VSUBS 1.3684f
C1100 VP.n16 VSUBS 0.568317f
C1101 VP.n17 VSUBS 0.043854f
C1102 VP.n18 VSUBS 0.081323f
C1103 VP.t2 VSUBS 1.63598f
C1104 VP.n19 VSUBS 0.63152f
C1105 VP.t0 VSUBS 1.3684f
C1106 VP.n20 VSUBS 0.630751f
C1107 VP.n21 VSUBS 0.048403f
C1108 VP.n22 VSUBS 0.374879f
C1109 VP.n23 VSUBS 0.043854f
C1110 VP.n24 VSUBS 0.043854f
C1111 VP.n25 VSUBS 0.058289f
C1112 VP.n26 VSUBS 0.069209f
C1113 VP.n27 VSUBS 0.081323f
C1114 VP.n28 VSUBS 0.043854f
C1115 VP.n29 VSUBS 0.043854f
C1116 VP.n30 VSUBS 0.043854f
C1117 VP.n31 VSUBS 0.081323f
C1118 VP.n32 VSUBS 0.069209f
C1119 VP.n33 VSUBS 0.058289f
C1120 VP.n34 VSUBS 0.043854f
C1121 VP.n35 VSUBS 0.043854f
C1122 VP.n36 VSUBS 0.043854f
C1123 VP.n37 VSUBS 0.048403f
C1124 VP.n38 VSUBS 0.527141f
C1125 VP.n39 VSUBS 0.074097f
C1126 VP.n40 VSUBS 0.078796f
C1127 VP.n41 VSUBS 0.043854f
C1128 VP.n42 VSUBS 0.043854f
C1129 VP.n43 VSUBS 0.043854f
C1130 VP.n44 VSUBS 0.086608f
C1131 VP.n45 VSUBS 0.055629f
C1132 VP.n46 VSUBS 0.650452f
C1133 VP.n47 VSUBS 2.15282f
C1134 VP.n48 VSUBS 2.18713f
C1135 VP.n49 VSUBS 0.650452f
C1136 VP.n50 VSUBS 0.055629f
C1137 VP.n51 VSUBS 0.086608f
C1138 VP.n52 VSUBS 0.043854f
C1139 VP.n53 VSUBS 0.043854f
C1140 VP.n54 VSUBS 0.043854f
C1141 VP.n55 VSUBS 0.078796f
C1142 VP.n56 VSUBS 0.074097f
C1143 VP.n57 VSUBS 0.527141f
C1144 VP.n58 VSUBS 0.048403f
C1145 VP.n59 VSUBS 0.043854f
C1146 VP.n60 VSUBS 0.043854f
C1147 VP.n61 VSUBS 0.043854f
C1148 VP.n62 VSUBS 0.058289f
C1149 VP.n63 VSUBS 0.069209f
C1150 VP.n64 VSUBS 0.081323f
C1151 VP.n65 VSUBS 0.043854f
C1152 VP.n66 VSUBS 0.043854f
C1153 VP.n67 VSUBS 0.043854f
C1154 VP.n68 VSUBS 0.081323f
C1155 VP.n69 VSUBS 0.069209f
C1156 VP.n70 VSUBS 0.058289f
C1157 VP.n71 VSUBS 0.043854f
C1158 VP.n72 VSUBS 0.043854f
C1159 VP.n73 VSUBS 0.043854f
C1160 VP.n74 VSUBS 0.048403f
C1161 VP.n75 VSUBS 0.527141f
C1162 VP.n76 VSUBS 0.074097f
C1163 VP.n77 VSUBS 0.078796f
C1164 VP.n78 VSUBS 0.043854f
C1165 VP.n79 VSUBS 0.043854f
C1166 VP.n80 VSUBS 0.043854f
C1167 VP.n81 VSUBS 0.086608f
C1168 VP.n82 VSUBS 0.055629f
C1169 VP.n83 VSUBS 0.650452f
C1170 VP.n84 VSUBS 0.067761f
.ends

