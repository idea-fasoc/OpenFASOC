* NGSPICE file created from diff_pair_sample_1552.ext - technology: sky130A

.subckt diff_pair_sample_1552 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=2.2152 ps=12.14 w=5.68 l=0.78
X1 VDD1.t0 VP.t1 VTAIL.t2 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=2.2152 ps=12.14 w=5.68 l=0.78
X2 B.t11 B.t9 B.t10 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=0.78
X3 B.t8 B.t6 B.t7 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=0.78
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=2.2152 ps=12.14 w=5.68 l=0.78
X5 B.t5 B.t3 B.t4 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=0.78
X6 B.t2 B.t0 B.t1 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=0 ps=0 w=5.68 l=0.78
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1414_n2108# sky130_fd_pr__pfet_01v8 ad=2.2152 pd=12.14 as=2.2152 ps=12.14 w=5.68 l=0.78
R0 VP.n0 VP.t1 422.217
R1 VP.n0 VP.t0 387.161
R2 VP VP.n0 0.0516364
R3 VTAIL.n1 VTAIL.t0 84.4602
R4 VTAIL.n2 VTAIL.t2 84.46
R5 VTAIL.n3 VTAIL.t1 84.4599
R6 VTAIL.n0 VTAIL.t3 84.4599
R7 VTAIL.n1 VTAIL.n0 19.1945
R8 VTAIL.n3 VTAIL.n2 18.2376
R9 VTAIL.n2 VTAIL.n1 0.948776
R10 VTAIL VTAIL.n0 0.767741
R11 VTAIL VTAIL.n3 0.181534
R12 VDD1 VDD1.t1 132.389
R13 VDD1 VDD1.t0 101.436
R14 B.n200 B.n57 585
R15 B.n199 B.n198 585
R16 B.n197 B.n58 585
R17 B.n196 B.n195 585
R18 B.n194 B.n59 585
R19 B.n193 B.n192 585
R20 B.n191 B.n60 585
R21 B.n190 B.n189 585
R22 B.n188 B.n61 585
R23 B.n187 B.n186 585
R24 B.n185 B.n62 585
R25 B.n184 B.n183 585
R26 B.n182 B.n63 585
R27 B.n181 B.n180 585
R28 B.n179 B.n64 585
R29 B.n178 B.n177 585
R30 B.n176 B.n65 585
R31 B.n175 B.n174 585
R32 B.n173 B.n66 585
R33 B.n172 B.n171 585
R34 B.n170 B.n67 585
R35 B.n169 B.n168 585
R36 B.n167 B.n68 585
R37 B.n165 B.n164 585
R38 B.n163 B.n71 585
R39 B.n162 B.n161 585
R40 B.n160 B.n72 585
R41 B.n159 B.n158 585
R42 B.n157 B.n73 585
R43 B.n156 B.n155 585
R44 B.n154 B.n74 585
R45 B.n153 B.n152 585
R46 B.n151 B.n75 585
R47 B.n150 B.n149 585
R48 B.n145 B.n76 585
R49 B.n144 B.n143 585
R50 B.n142 B.n77 585
R51 B.n141 B.n140 585
R52 B.n139 B.n78 585
R53 B.n138 B.n137 585
R54 B.n136 B.n79 585
R55 B.n135 B.n134 585
R56 B.n133 B.n80 585
R57 B.n132 B.n131 585
R58 B.n130 B.n81 585
R59 B.n129 B.n128 585
R60 B.n127 B.n82 585
R61 B.n126 B.n125 585
R62 B.n124 B.n83 585
R63 B.n123 B.n122 585
R64 B.n121 B.n84 585
R65 B.n120 B.n119 585
R66 B.n118 B.n85 585
R67 B.n117 B.n116 585
R68 B.n115 B.n86 585
R69 B.n114 B.n113 585
R70 B.n202 B.n201 585
R71 B.n203 B.n56 585
R72 B.n205 B.n204 585
R73 B.n206 B.n55 585
R74 B.n208 B.n207 585
R75 B.n209 B.n54 585
R76 B.n211 B.n210 585
R77 B.n212 B.n53 585
R78 B.n214 B.n213 585
R79 B.n215 B.n52 585
R80 B.n217 B.n216 585
R81 B.n218 B.n51 585
R82 B.n220 B.n219 585
R83 B.n221 B.n50 585
R84 B.n223 B.n222 585
R85 B.n224 B.n49 585
R86 B.n226 B.n225 585
R87 B.n227 B.n48 585
R88 B.n229 B.n228 585
R89 B.n230 B.n47 585
R90 B.n232 B.n231 585
R91 B.n233 B.n46 585
R92 B.n235 B.n234 585
R93 B.n236 B.n45 585
R94 B.n238 B.n237 585
R95 B.n239 B.n44 585
R96 B.n241 B.n240 585
R97 B.n242 B.n43 585
R98 B.n244 B.n243 585
R99 B.n245 B.n42 585
R100 B.n330 B.n9 585
R101 B.n329 B.n328 585
R102 B.n327 B.n10 585
R103 B.n326 B.n325 585
R104 B.n324 B.n11 585
R105 B.n323 B.n322 585
R106 B.n321 B.n12 585
R107 B.n320 B.n319 585
R108 B.n318 B.n13 585
R109 B.n317 B.n316 585
R110 B.n315 B.n14 585
R111 B.n314 B.n313 585
R112 B.n312 B.n15 585
R113 B.n311 B.n310 585
R114 B.n309 B.n16 585
R115 B.n308 B.n307 585
R116 B.n306 B.n17 585
R117 B.n305 B.n304 585
R118 B.n303 B.n18 585
R119 B.n302 B.n301 585
R120 B.n300 B.n19 585
R121 B.n299 B.n298 585
R122 B.n297 B.n20 585
R123 B.n296 B.n295 585
R124 B.n294 B.n21 585
R125 B.n293 B.n292 585
R126 B.n291 B.n25 585
R127 B.n290 B.n289 585
R128 B.n288 B.n26 585
R129 B.n287 B.n286 585
R130 B.n285 B.n27 585
R131 B.n284 B.n283 585
R132 B.n282 B.n28 585
R133 B.n280 B.n279 585
R134 B.n278 B.n31 585
R135 B.n277 B.n276 585
R136 B.n275 B.n32 585
R137 B.n274 B.n273 585
R138 B.n272 B.n33 585
R139 B.n271 B.n270 585
R140 B.n269 B.n34 585
R141 B.n268 B.n267 585
R142 B.n266 B.n35 585
R143 B.n265 B.n264 585
R144 B.n263 B.n36 585
R145 B.n262 B.n261 585
R146 B.n260 B.n37 585
R147 B.n259 B.n258 585
R148 B.n257 B.n38 585
R149 B.n256 B.n255 585
R150 B.n254 B.n39 585
R151 B.n253 B.n252 585
R152 B.n251 B.n40 585
R153 B.n250 B.n249 585
R154 B.n248 B.n41 585
R155 B.n247 B.n246 585
R156 B.n332 B.n331 585
R157 B.n333 B.n8 585
R158 B.n335 B.n334 585
R159 B.n336 B.n7 585
R160 B.n338 B.n337 585
R161 B.n339 B.n6 585
R162 B.n341 B.n340 585
R163 B.n342 B.n5 585
R164 B.n344 B.n343 585
R165 B.n345 B.n4 585
R166 B.n347 B.n346 585
R167 B.n348 B.n3 585
R168 B.n350 B.n349 585
R169 B.n351 B.n0 585
R170 B.n2 B.n1 585
R171 B.n94 B.n93 585
R172 B.n96 B.n95 585
R173 B.n97 B.n92 585
R174 B.n99 B.n98 585
R175 B.n100 B.n91 585
R176 B.n102 B.n101 585
R177 B.n103 B.n90 585
R178 B.n105 B.n104 585
R179 B.n106 B.n89 585
R180 B.n108 B.n107 585
R181 B.n109 B.n88 585
R182 B.n111 B.n110 585
R183 B.n112 B.n87 585
R184 B.n113 B.n112 502.111
R185 B.n201 B.n200 502.111
R186 B.n247 B.n42 502.111
R187 B.n332 B.n9 502.111
R188 B.n146 B.t9 377.579
R189 B.n69 B.t6 377.579
R190 B.n29 B.t0 377.579
R191 B.n22 B.t3 377.579
R192 B.n353 B.n352 256.663
R193 B.n352 B.n351 235.042
R194 B.n352 B.n2 235.042
R195 B.n113 B.n86 163.367
R196 B.n117 B.n86 163.367
R197 B.n118 B.n117 163.367
R198 B.n119 B.n118 163.367
R199 B.n119 B.n84 163.367
R200 B.n123 B.n84 163.367
R201 B.n124 B.n123 163.367
R202 B.n125 B.n124 163.367
R203 B.n125 B.n82 163.367
R204 B.n129 B.n82 163.367
R205 B.n130 B.n129 163.367
R206 B.n131 B.n130 163.367
R207 B.n131 B.n80 163.367
R208 B.n135 B.n80 163.367
R209 B.n136 B.n135 163.367
R210 B.n137 B.n136 163.367
R211 B.n137 B.n78 163.367
R212 B.n141 B.n78 163.367
R213 B.n142 B.n141 163.367
R214 B.n143 B.n142 163.367
R215 B.n143 B.n76 163.367
R216 B.n150 B.n76 163.367
R217 B.n151 B.n150 163.367
R218 B.n152 B.n151 163.367
R219 B.n152 B.n74 163.367
R220 B.n156 B.n74 163.367
R221 B.n157 B.n156 163.367
R222 B.n158 B.n157 163.367
R223 B.n158 B.n72 163.367
R224 B.n162 B.n72 163.367
R225 B.n163 B.n162 163.367
R226 B.n164 B.n163 163.367
R227 B.n164 B.n68 163.367
R228 B.n169 B.n68 163.367
R229 B.n170 B.n169 163.367
R230 B.n171 B.n170 163.367
R231 B.n171 B.n66 163.367
R232 B.n175 B.n66 163.367
R233 B.n176 B.n175 163.367
R234 B.n177 B.n176 163.367
R235 B.n177 B.n64 163.367
R236 B.n181 B.n64 163.367
R237 B.n182 B.n181 163.367
R238 B.n183 B.n182 163.367
R239 B.n183 B.n62 163.367
R240 B.n187 B.n62 163.367
R241 B.n188 B.n187 163.367
R242 B.n189 B.n188 163.367
R243 B.n189 B.n60 163.367
R244 B.n193 B.n60 163.367
R245 B.n194 B.n193 163.367
R246 B.n195 B.n194 163.367
R247 B.n195 B.n58 163.367
R248 B.n199 B.n58 163.367
R249 B.n200 B.n199 163.367
R250 B.n243 B.n42 163.367
R251 B.n243 B.n242 163.367
R252 B.n242 B.n241 163.367
R253 B.n241 B.n44 163.367
R254 B.n237 B.n44 163.367
R255 B.n237 B.n236 163.367
R256 B.n236 B.n235 163.367
R257 B.n235 B.n46 163.367
R258 B.n231 B.n46 163.367
R259 B.n231 B.n230 163.367
R260 B.n230 B.n229 163.367
R261 B.n229 B.n48 163.367
R262 B.n225 B.n48 163.367
R263 B.n225 B.n224 163.367
R264 B.n224 B.n223 163.367
R265 B.n223 B.n50 163.367
R266 B.n219 B.n50 163.367
R267 B.n219 B.n218 163.367
R268 B.n218 B.n217 163.367
R269 B.n217 B.n52 163.367
R270 B.n213 B.n52 163.367
R271 B.n213 B.n212 163.367
R272 B.n212 B.n211 163.367
R273 B.n211 B.n54 163.367
R274 B.n207 B.n54 163.367
R275 B.n207 B.n206 163.367
R276 B.n206 B.n205 163.367
R277 B.n205 B.n56 163.367
R278 B.n201 B.n56 163.367
R279 B.n328 B.n9 163.367
R280 B.n328 B.n327 163.367
R281 B.n327 B.n326 163.367
R282 B.n326 B.n11 163.367
R283 B.n322 B.n11 163.367
R284 B.n322 B.n321 163.367
R285 B.n321 B.n320 163.367
R286 B.n320 B.n13 163.367
R287 B.n316 B.n13 163.367
R288 B.n316 B.n315 163.367
R289 B.n315 B.n314 163.367
R290 B.n314 B.n15 163.367
R291 B.n310 B.n15 163.367
R292 B.n310 B.n309 163.367
R293 B.n309 B.n308 163.367
R294 B.n308 B.n17 163.367
R295 B.n304 B.n17 163.367
R296 B.n304 B.n303 163.367
R297 B.n303 B.n302 163.367
R298 B.n302 B.n19 163.367
R299 B.n298 B.n19 163.367
R300 B.n298 B.n297 163.367
R301 B.n297 B.n296 163.367
R302 B.n296 B.n21 163.367
R303 B.n292 B.n21 163.367
R304 B.n292 B.n291 163.367
R305 B.n291 B.n290 163.367
R306 B.n290 B.n26 163.367
R307 B.n286 B.n26 163.367
R308 B.n286 B.n285 163.367
R309 B.n285 B.n284 163.367
R310 B.n284 B.n28 163.367
R311 B.n279 B.n28 163.367
R312 B.n279 B.n278 163.367
R313 B.n278 B.n277 163.367
R314 B.n277 B.n32 163.367
R315 B.n273 B.n32 163.367
R316 B.n273 B.n272 163.367
R317 B.n272 B.n271 163.367
R318 B.n271 B.n34 163.367
R319 B.n267 B.n34 163.367
R320 B.n267 B.n266 163.367
R321 B.n266 B.n265 163.367
R322 B.n265 B.n36 163.367
R323 B.n261 B.n36 163.367
R324 B.n261 B.n260 163.367
R325 B.n260 B.n259 163.367
R326 B.n259 B.n38 163.367
R327 B.n255 B.n38 163.367
R328 B.n255 B.n254 163.367
R329 B.n254 B.n253 163.367
R330 B.n253 B.n40 163.367
R331 B.n249 B.n40 163.367
R332 B.n249 B.n248 163.367
R333 B.n248 B.n247 163.367
R334 B.n333 B.n332 163.367
R335 B.n334 B.n333 163.367
R336 B.n334 B.n7 163.367
R337 B.n338 B.n7 163.367
R338 B.n339 B.n338 163.367
R339 B.n340 B.n339 163.367
R340 B.n340 B.n5 163.367
R341 B.n344 B.n5 163.367
R342 B.n345 B.n344 163.367
R343 B.n346 B.n345 163.367
R344 B.n346 B.n3 163.367
R345 B.n350 B.n3 163.367
R346 B.n351 B.n350 163.367
R347 B.n94 B.n2 163.367
R348 B.n95 B.n94 163.367
R349 B.n95 B.n92 163.367
R350 B.n99 B.n92 163.367
R351 B.n100 B.n99 163.367
R352 B.n101 B.n100 163.367
R353 B.n101 B.n90 163.367
R354 B.n105 B.n90 163.367
R355 B.n106 B.n105 163.367
R356 B.n107 B.n106 163.367
R357 B.n107 B.n88 163.367
R358 B.n111 B.n88 163.367
R359 B.n112 B.n111 163.367
R360 B.n69 B.t7 138.263
R361 B.n29 B.t2 138.263
R362 B.n146 B.t10 138.258
R363 B.n22 B.t5 138.258
R364 B.n70 B.t8 116.737
R365 B.n30 B.t1 116.737
R366 B.n147 B.t11 116.731
R367 B.n23 B.t4 116.731
R368 B.n148 B.n147 59.5399
R369 B.n166 B.n70 59.5399
R370 B.n281 B.n30 59.5399
R371 B.n24 B.n23 59.5399
R372 B.n331 B.n330 32.6249
R373 B.n246 B.n245 32.6249
R374 B.n202 B.n57 32.6249
R375 B.n114 B.n87 32.6249
R376 B.n147 B.n146 21.5278
R377 B.n70 B.n69 21.5278
R378 B.n30 B.n29 21.5278
R379 B.n23 B.n22 21.5278
R380 B B.n353 18.0485
R381 B.n331 B.n8 10.6151
R382 B.n335 B.n8 10.6151
R383 B.n336 B.n335 10.6151
R384 B.n337 B.n336 10.6151
R385 B.n337 B.n6 10.6151
R386 B.n341 B.n6 10.6151
R387 B.n342 B.n341 10.6151
R388 B.n343 B.n342 10.6151
R389 B.n343 B.n4 10.6151
R390 B.n347 B.n4 10.6151
R391 B.n348 B.n347 10.6151
R392 B.n349 B.n348 10.6151
R393 B.n349 B.n0 10.6151
R394 B.n330 B.n329 10.6151
R395 B.n329 B.n10 10.6151
R396 B.n325 B.n10 10.6151
R397 B.n325 B.n324 10.6151
R398 B.n324 B.n323 10.6151
R399 B.n323 B.n12 10.6151
R400 B.n319 B.n12 10.6151
R401 B.n319 B.n318 10.6151
R402 B.n318 B.n317 10.6151
R403 B.n317 B.n14 10.6151
R404 B.n313 B.n14 10.6151
R405 B.n313 B.n312 10.6151
R406 B.n312 B.n311 10.6151
R407 B.n311 B.n16 10.6151
R408 B.n307 B.n16 10.6151
R409 B.n307 B.n306 10.6151
R410 B.n306 B.n305 10.6151
R411 B.n305 B.n18 10.6151
R412 B.n301 B.n18 10.6151
R413 B.n301 B.n300 10.6151
R414 B.n300 B.n299 10.6151
R415 B.n299 B.n20 10.6151
R416 B.n295 B.n294 10.6151
R417 B.n294 B.n293 10.6151
R418 B.n293 B.n25 10.6151
R419 B.n289 B.n25 10.6151
R420 B.n289 B.n288 10.6151
R421 B.n288 B.n287 10.6151
R422 B.n287 B.n27 10.6151
R423 B.n283 B.n27 10.6151
R424 B.n283 B.n282 10.6151
R425 B.n280 B.n31 10.6151
R426 B.n276 B.n31 10.6151
R427 B.n276 B.n275 10.6151
R428 B.n275 B.n274 10.6151
R429 B.n274 B.n33 10.6151
R430 B.n270 B.n33 10.6151
R431 B.n270 B.n269 10.6151
R432 B.n269 B.n268 10.6151
R433 B.n268 B.n35 10.6151
R434 B.n264 B.n35 10.6151
R435 B.n264 B.n263 10.6151
R436 B.n263 B.n262 10.6151
R437 B.n262 B.n37 10.6151
R438 B.n258 B.n37 10.6151
R439 B.n258 B.n257 10.6151
R440 B.n257 B.n256 10.6151
R441 B.n256 B.n39 10.6151
R442 B.n252 B.n39 10.6151
R443 B.n252 B.n251 10.6151
R444 B.n251 B.n250 10.6151
R445 B.n250 B.n41 10.6151
R446 B.n246 B.n41 10.6151
R447 B.n245 B.n244 10.6151
R448 B.n244 B.n43 10.6151
R449 B.n240 B.n43 10.6151
R450 B.n240 B.n239 10.6151
R451 B.n239 B.n238 10.6151
R452 B.n238 B.n45 10.6151
R453 B.n234 B.n45 10.6151
R454 B.n234 B.n233 10.6151
R455 B.n233 B.n232 10.6151
R456 B.n232 B.n47 10.6151
R457 B.n228 B.n47 10.6151
R458 B.n228 B.n227 10.6151
R459 B.n227 B.n226 10.6151
R460 B.n226 B.n49 10.6151
R461 B.n222 B.n49 10.6151
R462 B.n222 B.n221 10.6151
R463 B.n221 B.n220 10.6151
R464 B.n220 B.n51 10.6151
R465 B.n216 B.n51 10.6151
R466 B.n216 B.n215 10.6151
R467 B.n215 B.n214 10.6151
R468 B.n214 B.n53 10.6151
R469 B.n210 B.n53 10.6151
R470 B.n210 B.n209 10.6151
R471 B.n209 B.n208 10.6151
R472 B.n208 B.n55 10.6151
R473 B.n204 B.n55 10.6151
R474 B.n204 B.n203 10.6151
R475 B.n203 B.n202 10.6151
R476 B.n93 B.n1 10.6151
R477 B.n96 B.n93 10.6151
R478 B.n97 B.n96 10.6151
R479 B.n98 B.n97 10.6151
R480 B.n98 B.n91 10.6151
R481 B.n102 B.n91 10.6151
R482 B.n103 B.n102 10.6151
R483 B.n104 B.n103 10.6151
R484 B.n104 B.n89 10.6151
R485 B.n108 B.n89 10.6151
R486 B.n109 B.n108 10.6151
R487 B.n110 B.n109 10.6151
R488 B.n110 B.n87 10.6151
R489 B.n115 B.n114 10.6151
R490 B.n116 B.n115 10.6151
R491 B.n116 B.n85 10.6151
R492 B.n120 B.n85 10.6151
R493 B.n121 B.n120 10.6151
R494 B.n122 B.n121 10.6151
R495 B.n122 B.n83 10.6151
R496 B.n126 B.n83 10.6151
R497 B.n127 B.n126 10.6151
R498 B.n128 B.n127 10.6151
R499 B.n128 B.n81 10.6151
R500 B.n132 B.n81 10.6151
R501 B.n133 B.n132 10.6151
R502 B.n134 B.n133 10.6151
R503 B.n134 B.n79 10.6151
R504 B.n138 B.n79 10.6151
R505 B.n139 B.n138 10.6151
R506 B.n140 B.n139 10.6151
R507 B.n140 B.n77 10.6151
R508 B.n144 B.n77 10.6151
R509 B.n145 B.n144 10.6151
R510 B.n149 B.n145 10.6151
R511 B.n153 B.n75 10.6151
R512 B.n154 B.n153 10.6151
R513 B.n155 B.n154 10.6151
R514 B.n155 B.n73 10.6151
R515 B.n159 B.n73 10.6151
R516 B.n160 B.n159 10.6151
R517 B.n161 B.n160 10.6151
R518 B.n161 B.n71 10.6151
R519 B.n165 B.n71 10.6151
R520 B.n168 B.n167 10.6151
R521 B.n168 B.n67 10.6151
R522 B.n172 B.n67 10.6151
R523 B.n173 B.n172 10.6151
R524 B.n174 B.n173 10.6151
R525 B.n174 B.n65 10.6151
R526 B.n178 B.n65 10.6151
R527 B.n179 B.n178 10.6151
R528 B.n180 B.n179 10.6151
R529 B.n180 B.n63 10.6151
R530 B.n184 B.n63 10.6151
R531 B.n185 B.n184 10.6151
R532 B.n186 B.n185 10.6151
R533 B.n186 B.n61 10.6151
R534 B.n190 B.n61 10.6151
R535 B.n191 B.n190 10.6151
R536 B.n192 B.n191 10.6151
R537 B.n192 B.n59 10.6151
R538 B.n196 B.n59 10.6151
R539 B.n197 B.n196 10.6151
R540 B.n198 B.n197 10.6151
R541 B.n198 B.n57 10.6151
R542 B.n24 B.n20 8.74196
R543 B.n281 B.n280 8.74196
R544 B.n149 B.n148 8.74196
R545 B.n167 B.n166 8.74196
R546 B.n353 B.n0 8.11757
R547 B.n353 B.n1 8.11757
R548 B.n295 B.n24 1.87367
R549 B.n282 B.n281 1.87367
R550 B.n148 B.n75 1.87367
R551 B.n166 B.n165 1.87367
R552 VN VN.t1 422.599
R553 VN VN.t0 387.212
R554 VDD2.n0 VDD2.t1 131.625
R555 VDD2.n0 VDD2.t0 101.138
R556 VDD2 VDD2.n0 0.297914
C0 B VP 0.949076f
C1 VP VDD1 1.20895f
C2 w_n1414_n2108# VN 1.67291f
C3 B VN 0.66671f
C4 w_n1414_n2108# B 5.07874f
C5 VDD1 VN 0.148958f
C6 w_n1414_n2108# VDD1 1.11551f
C7 B VDD1 0.967426f
C8 VTAIL VDD2 3.31974f
C9 VP VTAIL 0.94721f
C10 VTAIL VN 0.932879f
C11 w_n1414_n2108# VTAIL 1.85943f
C12 B VTAIL 1.60891f
C13 VDD1 VTAIL 3.28168f
C14 VP VDD2 0.257723f
C15 VN VDD2 1.10228f
C16 w_n1414_n2108# VDD2 1.12088f
C17 VP VN 3.42542f
C18 B VDD2 0.982582f
C19 w_n1414_n2108# VP 1.84911f
C20 VDD1 VDD2 0.468206f
C21 VDD2 VSUBS 0.525457f
C22 VDD1 VSUBS 2.510441f
C23 VTAIL VSUBS 0.426079f
C24 VN VSUBS 3.643759f
C25 VP VSUBS 0.839325f
C26 B VSUBS 1.945086f
C27 w_n1414_n2108# VSUBS 37.2448f
C28 VDD2.t1 VSUBS 0.820221f
C29 VDD2.t0 VSUBS 0.620578f
C30 VDD2.n0 VSUBS 1.81944f
C31 VN.t0 VSUBS 0.520515f
C32 VN.t1 VSUBS 0.617812f
C33 B.n0 VSUBS 0.005894f
C34 B.n1 VSUBS 0.005894f
C35 B.n2 VSUBS 0.008717f
C36 B.n3 VSUBS 0.00668f
C37 B.n4 VSUBS 0.00668f
C38 B.n5 VSUBS 0.00668f
C39 B.n6 VSUBS 0.00668f
C40 B.n7 VSUBS 0.00668f
C41 B.n8 VSUBS 0.00668f
C42 B.n9 VSUBS 0.016168f
C43 B.n10 VSUBS 0.00668f
C44 B.n11 VSUBS 0.00668f
C45 B.n12 VSUBS 0.00668f
C46 B.n13 VSUBS 0.00668f
C47 B.n14 VSUBS 0.00668f
C48 B.n15 VSUBS 0.00668f
C49 B.n16 VSUBS 0.00668f
C50 B.n17 VSUBS 0.00668f
C51 B.n18 VSUBS 0.00668f
C52 B.n19 VSUBS 0.00668f
C53 B.n20 VSUBS 0.00609f
C54 B.n21 VSUBS 0.00668f
C55 B.t4 VSUBS 0.156107f
C56 B.t5 VSUBS 0.164018f
C57 B.t3 VSUBS 0.185277f
C58 B.n22 VSUBS 0.083911f
C59 B.n23 VSUBS 0.060337f
C60 B.n24 VSUBS 0.015476f
C61 B.n25 VSUBS 0.00668f
C62 B.n26 VSUBS 0.00668f
C63 B.n27 VSUBS 0.00668f
C64 B.n28 VSUBS 0.00668f
C65 B.t1 VSUBS 0.156107f
C66 B.t2 VSUBS 0.164018f
C67 B.t0 VSUBS 0.185277f
C68 B.n29 VSUBS 0.083911f
C69 B.n30 VSUBS 0.060337f
C70 B.n31 VSUBS 0.00668f
C71 B.n32 VSUBS 0.00668f
C72 B.n33 VSUBS 0.00668f
C73 B.n34 VSUBS 0.00668f
C74 B.n35 VSUBS 0.00668f
C75 B.n36 VSUBS 0.00668f
C76 B.n37 VSUBS 0.00668f
C77 B.n38 VSUBS 0.00668f
C78 B.n39 VSUBS 0.00668f
C79 B.n40 VSUBS 0.00668f
C80 B.n41 VSUBS 0.00668f
C81 B.n42 VSUBS 0.01507f
C82 B.n43 VSUBS 0.00668f
C83 B.n44 VSUBS 0.00668f
C84 B.n45 VSUBS 0.00668f
C85 B.n46 VSUBS 0.00668f
C86 B.n47 VSUBS 0.00668f
C87 B.n48 VSUBS 0.00668f
C88 B.n49 VSUBS 0.00668f
C89 B.n50 VSUBS 0.00668f
C90 B.n51 VSUBS 0.00668f
C91 B.n52 VSUBS 0.00668f
C92 B.n53 VSUBS 0.00668f
C93 B.n54 VSUBS 0.00668f
C94 B.n55 VSUBS 0.00668f
C95 B.n56 VSUBS 0.00668f
C96 B.n57 VSUBS 0.015378f
C97 B.n58 VSUBS 0.00668f
C98 B.n59 VSUBS 0.00668f
C99 B.n60 VSUBS 0.00668f
C100 B.n61 VSUBS 0.00668f
C101 B.n62 VSUBS 0.00668f
C102 B.n63 VSUBS 0.00668f
C103 B.n64 VSUBS 0.00668f
C104 B.n65 VSUBS 0.00668f
C105 B.n66 VSUBS 0.00668f
C106 B.n67 VSUBS 0.00668f
C107 B.n68 VSUBS 0.00668f
C108 B.t8 VSUBS 0.156107f
C109 B.t7 VSUBS 0.164018f
C110 B.t6 VSUBS 0.185277f
C111 B.n69 VSUBS 0.083911f
C112 B.n70 VSUBS 0.060337f
C113 B.n71 VSUBS 0.00668f
C114 B.n72 VSUBS 0.00668f
C115 B.n73 VSUBS 0.00668f
C116 B.n74 VSUBS 0.00668f
C117 B.n75 VSUBS 0.003929f
C118 B.n76 VSUBS 0.00668f
C119 B.n77 VSUBS 0.00668f
C120 B.n78 VSUBS 0.00668f
C121 B.n79 VSUBS 0.00668f
C122 B.n80 VSUBS 0.00668f
C123 B.n81 VSUBS 0.00668f
C124 B.n82 VSUBS 0.00668f
C125 B.n83 VSUBS 0.00668f
C126 B.n84 VSUBS 0.00668f
C127 B.n85 VSUBS 0.00668f
C128 B.n86 VSUBS 0.00668f
C129 B.n87 VSUBS 0.01507f
C130 B.n88 VSUBS 0.00668f
C131 B.n89 VSUBS 0.00668f
C132 B.n90 VSUBS 0.00668f
C133 B.n91 VSUBS 0.00668f
C134 B.n92 VSUBS 0.00668f
C135 B.n93 VSUBS 0.00668f
C136 B.n94 VSUBS 0.00668f
C137 B.n95 VSUBS 0.00668f
C138 B.n96 VSUBS 0.00668f
C139 B.n97 VSUBS 0.00668f
C140 B.n98 VSUBS 0.00668f
C141 B.n99 VSUBS 0.00668f
C142 B.n100 VSUBS 0.00668f
C143 B.n101 VSUBS 0.00668f
C144 B.n102 VSUBS 0.00668f
C145 B.n103 VSUBS 0.00668f
C146 B.n104 VSUBS 0.00668f
C147 B.n105 VSUBS 0.00668f
C148 B.n106 VSUBS 0.00668f
C149 B.n107 VSUBS 0.00668f
C150 B.n108 VSUBS 0.00668f
C151 B.n109 VSUBS 0.00668f
C152 B.n110 VSUBS 0.00668f
C153 B.n111 VSUBS 0.00668f
C154 B.n112 VSUBS 0.01507f
C155 B.n113 VSUBS 0.016168f
C156 B.n114 VSUBS 0.016168f
C157 B.n115 VSUBS 0.00668f
C158 B.n116 VSUBS 0.00668f
C159 B.n117 VSUBS 0.00668f
C160 B.n118 VSUBS 0.00668f
C161 B.n119 VSUBS 0.00668f
C162 B.n120 VSUBS 0.00668f
C163 B.n121 VSUBS 0.00668f
C164 B.n122 VSUBS 0.00668f
C165 B.n123 VSUBS 0.00668f
C166 B.n124 VSUBS 0.00668f
C167 B.n125 VSUBS 0.00668f
C168 B.n126 VSUBS 0.00668f
C169 B.n127 VSUBS 0.00668f
C170 B.n128 VSUBS 0.00668f
C171 B.n129 VSUBS 0.00668f
C172 B.n130 VSUBS 0.00668f
C173 B.n131 VSUBS 0.00668f
C174 B.n132 VSUBS 0.00668f
C175 B.n133 VSUBS 0.00668f
C176 B.n134 VSUBS 0.00668f
C177 B.n135 VSUBS 0.00668f
C178 B.n136 VSUBS 0.00668f
C179 B.n137 VSUBS 0.00668f
C180 B.n138 VSUBS 0.00668f
C181 B.n139 VSUBS 0.00668f
C182 B.n140 VSUBS 0.00668f
C183 B.n141 VSUBS 0.00668f
C184 B.n142 VSUBS 0.00668f
C185 B.n143 VSUBS 0.00668f
C186 B.n144 VSUBS 0.00668f
C187 B.n145 VSUBS 0.00668f
C188 B.t11 VSUBS 0.156107f
C189 B.t10 VSUBS 0.164018f
C190 B.t9 VSUBS 0.185277f
C191 B.n146 VSUBS 0.083911f
C192 B.n147 VSUBS 0.060337f
C193 B.n148 VSUBS 0.015476f
C194 B.n149 VSUBS 0.00609f
C195 B.n150 VSUBS 0.00668f
C196 B.n151 VSUBS 0.00668f
C197 B.n152 VSUBS 0.00668f
C198 B.n153 VSUBS 0.00668f
C199 B.n154 VSUBS 0.00668f
C200 B.n155 VSUBS 0.00668f
C201 B.n156 VSUBS 0.00668f
C202 B.n157 VSUBS 0.00668f
C203 B.n158 VSUBS 0.00668f
C204 B.n159 VSUBS 0.00668f
C205 B.n160 VSUBS 0.00668f
C206 B.n161 VSUBS 0.00668f
C207 B.n162 VSUBS 0.00668f
C208 B.n163 VSUBS 0.00668f
C209 B.n164 VSUBS 0.00668f
C210 B.n165 VSUBS 0.003929f
C211 B.n166 VSUBS 0.015476f
C212 B.n167 VSUBS 0.00609f
C213 B.n168 VSUBS 0.00668f
C214 B.n169 VSUBS 0.00668f
C215 B.n170 VSUBS 0.00668f
C216 B.n171 VSUBS 0.00668f
C217 B.n172 VSUBS 0.00668f
C218 B.n173 VSUBS 0.00668f
C219 B.n174 VSUBS 0.00668f
C220 B.n175 VSUBS 0.00668f
C221 B.n176 VSUBS 0.00668f
C222 B.n177 VSUBS 0.00668f
C223 B.n178 VSUBS 0.00668f
C224 B.n179 VSUBS 0.00668f
C225 B.n180 VSUBS 0.00668f
C226 B.n181 VSUBS 0.00668f
C227 B.n182 VSUBS 0.00668f
C228 B.n183 VSUBS 0.00668f
C229 B.n184 VSUBS 0.00668f
C230 B.n185 VSUBS 0.00668f
C231 B.n186 VSUBS 0.00668f
C232 B.n187 VSUBS 0.00668f
C233 B.n188 VSUBS 0.00668f
C234 B.n189 VSUBS 0.00668f
C235 B.n190 VSUBS 0.00668f
C236 B.n191 VSUBS 0.00668f
C237 B.n192 VSUBS 0.00668f
C238 B.n193 VSUBS 0.00668f
C239 B.n194 VSUBS 0.00668f
C240 B.n195 VSUBS 0.00668f
C241 B.n196 VSUBS 0.00668f
C242 B.n197 VSUBS 0.00668f
C243 B.n198 VSUBS 0.00668f
C244 B.n199 VSUBS 0.00668f
C245 B.n200 VSUBS 0.016168f
C246 B.n201 VSUBS 0.01507f
C247 B.n202 VSUBS 0.01586f
C248 B.n203 VSUBS 0.00668f
C249 B.n204 VSUBS 0.00668f
C250 B.n205 VSUBS 0.00668f
C251 B.n206 VSUBS 0.00668f
C252 B.n207 VSUBS 0.00668f
C253 B.n208 VSUBS 0.00668f
C254 B.n209 VSUBS 0.00668f
C255 B.n210 VSUBS 0.00668f
C256 B.n211 VSUBS 0.00668f
C257 B.n212 VSUBS 0.00668f
C258 B.n213 VSUBS 0.00668f
C259 B.n214 VSUBS 0.00668f
C260 B.n215 VSUBS 0.00668f
C261 B.n216 VSUBS 0.00668f
C262 B.n217 VSUBS 0.00668f
C263 B.n218 VSUBS 0.00668f
C264 B.n219 VSUBS 0.00668f
C265 B.n220 VSUBS 0.00668f
C266 B.n221 VSUBS 0.00668f
C267 B.n222 VSUBS 0.00668f
C268 B.n223 VSUBS 0.00668f
C269 B.n224 VSUBS 0.00668f
C270 B.n225 VSUBS 0.00668f
C271 B.n226 VSUBS 0.00668f
C272 B.n227 VSUBS 0.00668f
C273 B.n228 VSUBS 0.00668f
C274 B.n229 VSUBS 0.00668f
C275 B.n230 VSUBS 0.00668f
C276 B.n231 VSUBS 0.00668f
C277 B.n232 VSUBS 0.00668f
C278 B.n233 VSUBS 0.00668f
C279 B.n234 VSUBS 0.00668f
C280 B.n235 VSUBS 0.00668f
C281 B.n236 VSUBS 0.00668f
C282 B.n237 VSUBS 0.00668f
C283 B.n238 VSUBS 0.00668f
C284 B.n239 VSUBS 0.00668f
C285 B.n240 VSUBS 0.00668f
C286 B.n241 VSUBS 0.00668f
C287 B.n242 VSUBS 0.00668f
C288 B.n243 VSUBS 0.00668f
C289 B.n244 VSUBS 0.00668f
C290 B.n245 VSUBS 0.01507f
C291 B.n246 VSUBS 0.016168f
C292 B.n247 VSUBS 0.016168f
C293 B.n248 VSUBS 0.00668f
C294 B.n249 VSUBS 0.00668f
C295 B.n250 VSUBS 0.00668f
C296 B.n251 VSUBS 0.00668f
C297 B.n252 VSUBS 0.00668f
C298 B.n253 VSUBS 0.00668f
C299 B.n254 VSUBS 0.00668f
C300 B.n255 VSUBS 0.00668f
C301 B.n256 VSUBS 0.00668f
C302 B.n257 VSUBS 0.00668f
C303 B.n258 VSUBS 0.00668f
C304 B.n259 VSUBS 0.00668f
C305 B.n260 VSUBS 0.00668f
C306 B.n261 VSUBS 0.00668f
C307 B.n262 VSUBS 0.00668f
C308 B.n263 VSUBS 0.00668f
C309 B.n264 VSUBS 0.00668f
C310 B.n265 VSUBS 0.00668f
C311 B.n266 VSUBS 0.00668f
C312 B.n267 VSUBS 0.00668f
C313 B.n268 VSUBS 0.00668f
C314 B.n269 VSUBS 0.00668f
C315 B.n270 VSUBS 0.00668f
C316 B.n271 VSUBS 0.00668f
C317 B.n272 VSUBS 0.00668f
C318 B.n273 VSUBS 0.00668f
C319 B.n274 VSUBS 0.00668f
C320 B.n275 VSUBS 0.00668f
C321 B.n276 VSUBS 0.00668f
C322 B.n277 VSUBS 0.00668f
C323 B.n278 VSUBS 0.00668f
C324 B.n279 VSUBS 0.00668f
C325 B.n280 VSUBS 0.00609f
C326 B.n281 VSUBS 0.015476f
C327 B.n282 VSUBS 0.003929f
C328 B.n283 VSUBS 0.00668f
C329 B.n284 VSUBS 0.00668f
C330 B.n285 VSUBS 0.00668f
C331 B.n286 VSUBS 0.00668f
C332 B.n287 VSUBS 0.00668f
C333 B.n288 VSUBS 0.00668f
C334 B.n289 VSUBS 0.00668f
C335 B.n290 VSUBS 0.00668f
C336 B.n291 VSUBS 0.00668f
C337 B.n292 VSUBS 0.00668f
C338 B.n293 VSUBS 0.00668f
C339 B.n294 VSUBS 0.00668f
C340 B.n295 VSUBS 0.003929f
C341 B.n296 VSUBS 0.00668f
C342 B.n297 VSUBS 0.00668f
C343 B.n298 VSUBS 0.00668f
C344 B.n299 VSUBS 0.00668f
C345 B.n300 VSUBS 0.00668f
C346 B.n301 VSUBS 0.00668f
C347 B.n302 VSUBS 0.00668f
C348 B.n303 VSUBS 0.00668f
C349 B.n304 VSUBS 0.00668f
C350 B.n305 VSUBS 0.00668f
C351 B.n306 VSUBS 0.00668f
C352 B.n307 VSUBS 0.00668f
C353 B.n308 VSUBS 0.00668f
C354 B.n309 VSUBS 0.00668f
C355 B.n310 VSUBS 0.00668f
C356 B.n311 VSUBS 0.00668f
C357 B.n312 VSUBS 0.00668f
C358 B.n313 VSUBS 0.00668f
C359 B.n314 VSUBS 0.00668f
C360 B.n315 VSUBS 0.00668f
C361 B.n316 VSUBS 0.00668f
C362 B.n317 VSUBS 0.00668f
C363 B.n318 VSUBS 0.00668f
C364 B.n319 VSUBS 0.00668f
C365 B.n320 VSUBS 0.00668f
C366 B.n321 VSUBS 0.00668f
C367 B.n322 VSUBS 0.00668f
C368 B.n323 VSUBS 0.00668f
C369 B.n324 VSUBS 0.00668f
C370 B.n325 VSUBS 0.00668f
C371 B.n326 VSUBS 0.00668f
C372 B.n327 VSUBS 0.00668f
C373 B.n328 VSUBS 0.00668f
C374 B.n329 VSUBS 0.00668f
C375 B.n330 VSUBS 0.016168f
C376 B.n331 VSUBS 0.01507f
C377 B.n332 VSUBS 0.01507f
C378 B.n333 VSUBS 0.00668f
C379 B.n334 VSUBS 0.00668f
C380 B.n335 VSUBS 0.00668f
C381 B.n336 VSUBS 0.00668f
C382 B.n337 VSUBS 0.00668f
C383 B.n338 VSUBS 0.00668f
C384 B.n339 VSUBS 0.00668f
C385 B.n340 VSUBS 0.00668f
C386 B.n341 VSUBS 0.00668f
C387 B.n342 VSUBS 0.00668f
C388 B.n343 VSUBS 0.00668f
C389 B.n344 VSUBS 0.00668f
C390 B.n345 VSUBS 0.00668f
C391 B.n346 VSUBS 0.00668f
C392 B.n347 VSUBS 0.00668f
C393 B.n348 VSUBS 0.00668f
C394 B.n349 VSUBS 0.00668f
C395 B.n350 VSUBS 0.00668f
C396 B.n351 VSUBS 0.008717f
C397 B.n352 VSUBS 0.009286f
C398 B.n353 VSUBS 0.018465f
C399 VDD1.t0 VSUBS 0.610721f
C400 VDD1.t1 VSUBS 0.818864f
C401 VTAIL.t3 VSUBS 0.635846f
C402 VTAIL.n0 VSUBS 1.03111f
C403 VTAIL.t0 VSUBS 0.635849f
C404 VTAIL.n1 VSUBS 1.04144f
C405 VTAIL.t2 VSUBS 0.635846f
C406 VTAIL.n2 VSUBS 0.98687f
C407 VTAIL.t1 VSUBS 0.635846f
C408 VTAIL.n3 VSUBS 0.943118f
C409 VP.t1 VSUBS 0.623747f
C410 VP.t0 VSUBS 0.527918f
C411 VP.n0 VSUBS 2.23462f
.ends

