* NGSPICE file created from diff_pair_sample_0964.ext - technology: sky130A

.subckt diff_pair_sample_0964 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t6 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X1 VDD1.t9 VP.t0 VTAIL.t8 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X2 B.t11 B.t9 B.t10 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=2.68
X3 B.t8 B.t6 B.t7 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=2.68
X4 VDD1.t8 VP.t1 VTAIL.t0 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X5 VDD1.t7 VP.t2 VTAIL.t7 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0.65505 ps=4.3 w=3.97 l=2.68
X6 VTAIL.t17 VN.t1 VDD2.t4 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X7 VDD2.t9 VN.t2 VTAIL.t16 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X8 B.t5 B.t3 B.t4 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=2.68
X9 VTAIL.t1 VP.t3 VDD1.t6 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X10 VDD1.t5 VP.t4 VTAIL.t3 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0.65505 ps=4.3 w=3.97 l=2.68
X11 VDD2.t8 VN.t3 VTAIL.t15 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=1.5483 ps=8.72 w=3.97 l=2.68
X12 VTAIL.t4 VP.t5 VDD1.t4 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X13 VDD2.t2 VN.t4 VTAIL.t14 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0.65505 ps=4.3 w=3.97 l=2.68
X14 VDD1.t3 VP.t6 VTAIL.t2 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=1.5483 ps=8.72 w=3.97 l=2.68
X15 VTAIL.t19 VP.t7 VDD1.t2 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X16 VDD2.t3 VN.t5 VTAIL.t13 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X17 VTAIL.t12 VN.t6 VDD2.t1 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X18 VDD1.t1 VP.t8 VTAIL.t5 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=1.5483 ps=8.72 w=3.97 l=2.68
X19 VDD2.t0 VN.t7 VTAIL.t11 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=1.5483 ps=8.72 w=3.97 l=2.68
X20 VDD2.t7 VN.t8 VTAIL.t10 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0.65505 ps=4.3 w=3.97 l=2.68
X21 B.t2 B.t0 B.t1 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=2.68
X22 VTAIL.t6 VP.t9 VDD1.t0 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
X23 VTAIL.t9 VN.t9 VDD2.t5 w_n4582_n1762# sky130_fd_pr__pfet_01v8 ad=0.65505 pd=4.3 as=0.65505 ps=4.3 w=3.97 l=2.68
R0 VN.n83 VN.n43 161.3
R1 VN.n82 VN.n81 161.3
R2 VN.n80 VN.n44 161.3
R3 VN.n79 VN.n78 161.3
R4 VN.n77 VN.n45 161.3
R5 VN.n76 VN.n75 161.3
R6 VN.n74 VN.n73 161.3
R7 VN.n72 VN.n47 161.3
R8 VN.n71 VN.n70 161.3
R9 VN.n69 VN.n48 161.3
R10 VN.n68 VN.n67 161.3
R11 VN.n66 VN.n49 161.3
R12 VN.n65 VN.n64 161.3
R13 VN.n63 VN.n50 161.3
R14 VN.n62 VN.n61 161.3
R15 VN.n60 VN.n51 161.3
R16 VN.n59 VN.n58 161.3
R17 VN.n57 VN.n52 161.3
R18 VN.n56 VN.n55 161.3
R19 VN.n40 VN.n0 161.3
R20 VN.n39 VN.n38 161.3
R21 VN.n37 VN.n1 161.3
R22 VN.n36 VN.n35 161.3
R23 VN.n34 VN.n2 161.3
R24 VN.n33 VN.n32 161.3
R25 VN.n31 VN.n30 161.3
R26 VN.n29 VN.n4 161.3
R27 VN.n28 VN.n27 161.3
R28 VN.n26 VN.n5 161.3
R29 VN.n25 VN.n24 161.3
R30 VN.n23 VN.n6 161.3
R31 VN.n22 VN.n21 161.3
R32 VN.n20 VN.n7 161.3
R33 VN.n19 VN.n18 161.3
R34 VN.n17 VN.n8 161.3
R35 VN.n16 VN.n15 161.3
R36 VN.n14 VN.n9 161.3
R37 VN.n13 VN.n12 161.3
R38 VN.n42 VN.n41 109.778
R39 VN.n85 VN.n84 109.778
R40 VN.n11 VN.n10 72.9374
R41 VN.n54 VN.n53 72.9374
R42 VN.n10 VN.t8 65.9996
R43 VN.n53 VN.t3 65.9996
R44 VN VN.n85 47.6459
R45 VN.n35 VN.n1 41.9503
R46 VN.n78 VN.n44 41.9503
R47 VN.n17 VN.n16 40.979
R48 VN.n28 VN.n5 40.979
R49 VN.n60 VN.n59 40.979
R50 VN.n71 VN.n48 40.979
R51 VN.n18 VN.n17 40.0078
R52 VN.n24 VN.n5 40.0078
R53 VN.n61 VN.n60 40.0078
R54 VN.n67 VN.n48 40.0078
R55 VN.n35 VN.n34 39.0365
R56 VN.n78 VN.n77 39.0365
R57 VN.n22 VN.t2 35.7009
R58 VN.n11 VN.t6 35.7009
R59 VN.n3 VN.t0 35.7009
R60 VN.n41 VN.t7 35.7009
R61 VN.n65 VN.t5 35.7009
R62 VN.n54 VN.t9 35.7009
R63 VN.n46 VN.t1 35.7009
R64 VN.n84 VN.t4 35.7009
R65 VN.n12 VN.n9 24.4675
R66 VN.n16 VN.n9 24.4675
R67 VN.n18 VN.n7 24.4675
R68 VN.n22 VN.n7 24.4675
R69 VN.n23 VN.n22 24.4675
R70 VN.n24 VN.n23 24.4675
R71 VN.n29 VN.n28 24.4675
R72 VN.n30 VN.n29 24.4675
R73 VN.n34 VN.n33 24.4675
R74 VN.n39 VN.n1 24.4675
R75 VN.n40 VN.n39 24.4675
R76 VN.n59 VN.n52 24.4675
R77 VN.n55 VN.n52 24.4675
R78 VN.n67 VN.n66 24.4675
R79 VN.n66 VN.n65 24.4675
R80 VN.n65 VN.n50 24.4675
R81 VN.n61 VN.n50 24.4675
R82 VN.n77 VN.n76 24.4675
R83 VN.n73 VN.n72 24.4675
R84 VN.n72 VN.n71 24.4675
R85 VN.n83 VN.n82 24.4675
R86 VN.n82 VN.n44 24.4675
R87 VN.n33 VN.n3 23.9782
R88 VN.n76 VN.n46 23.9782
R89 VN.n56 VN.n53 7.44194
R90 VN.n13 VN.n10 7.44194
R91 VN.n41 VN.n40 0.97918
R92 VN.n84 VN.n83 0.97918
R93 VN.n12 VN.n11 0.48984
R94 VN.n30 VN.n3 0.48984
R95 VN.n55 VN.n54 0.48984
R96 VN.n73 VN.n46 0.48984
R97 VN.n85 VN.n43 0.278367
R98 VN.n42 VN.n0 0.278367
R99 VN.n81 VN.n43 0.189894
R100 VN.n81 VN.n80 0.189894
R101 VN.n80 VN.n79 0.189894
R102 VN.n79 VN.n45 0.189894
R103 VN.n75 VN.n45 0.189894
R104 VN.n75 VN.n74 0.189894
R105 VN.n74 VN.n47 0.189894
R106 VN.n70 VN.n47 0.189894
R107 VN.n70 VN.n69 0.189894
R108 VN.n69 VN.n68 0.189894
R109 VN.n68 VN.n49 0.189894
R110 VN.n64 VN.n49 0.189894
R111 VN.n64 VN.n63 0.189894
R112 VN.n63 VN.n62 0.189894
R113 VN.n62 VN.n51 0.189894
R114 VN.n58 VN.n51 0.189894
R115 VN.n58 VN.n57 0.189894
R116 VN.n57 VN.n56 0.189894
R117 VN.n14 VN.n13 0.189894
R118 VN.n15 VN.n14 0.189894
R119 VN.n15 VN.n8 0.189894
R120 VN.n19 VN.n8 0.189894
R121 VN.n20 VN.n19 0.189894
R122 VN.n21 VN.n20 0.189894
R123 VN.n21 VN.n6 0.189894
R124 VN.n25 VN.n6 0.189894
R125 VN.n26 VN.n25 0.189894
R126 VN.n27 VN.n26 0.189894
R127 VN.n27 VN.n4 0.189894
R128 VN.n31 VN.n4 0.189894
R129 VN.n32 VN.n31 0.189894
R130 VN.n32 VN.n2 0.189894
R131 VN.n36 VN.n2 0.189894
R132 VN.n37 VN.n36 0.189894
R133 VN.n38 VN.n37 0.189894
R134 VN.n38 VN.n0 0.189894
R135 VN VN.n42 0.153454
R136 VDD2.n37 VDD2.n23 756.745
R137 VDD2.n14 VDD2.n0 756.745
R138 VDD2.n38 VDD2.n37 585
R139 VDD2.n36 VDD2.n35 585
R140 VDD2.n27 VDD2.n26 585
R141 VDD2.n30 VDD2.n29 585
R142 VDD2.n7 VDD2.n6 585
R143 VDD2.n4 VDD2.n3 585
R144 VDD2.n13 VDD2.n12 585
R145 VDD2.n15 VDD2.n14 585
R146 VDD2.t2 VDD2.n28 330.707
R147 VDD2.t7 VDD2.n5 330.707
R148 VDD2.n37 VDD2.n36 171.744
R149 VDD2.n36 VDD2.n26 171.744
R150 VDD2.n29 VDD2.n26 171.744
R151 VDD2.n6 VDD2.n3 171.744
R152 VDD2.n13 VDD2.n3 171.744
R153 VDD2.n14 VDD2.n13 171.744
R154 VDD2.n22 VDD2.n21 117.981
R155 VDD2 VDD2.n45 117.978
R156 VDD2.n44 VDD2.n43 116.09
R157 VDD2.n20 VDD2.n19 116.09
R158 VDD2.n29 VDD2.t2 85.8723
R159 VDD2.n6 VDD2.t7 85.8723
R160 VDD2.n20 VDD2.n18 53.9802
R161 VDD2.n42 VDD2.n41 51.3853
R162 VDD2.n42 VDD2.n22 39.4631
R163 VDD2.n30 VDD2.n28 16.3201
R164 VDD2.n7 VDD2.n5 16.3201
R165 VDD2.n31 VDD2.n27 12.8005
R166 VDD2.n8 VDD2.n4 12.8005
R167 VDD2.n35 VDD2.n34 12.0247
R168 VDD2.n12 VDD2.n11 12.0247
R169 VDD2.n38 VDD2.n25 11.249
R170 VDD2.n15 VDD2.n2 11.249
R171 VDD2.n39 VDD2.n23 10.4732
R172 VDD2.n16 VDD2.n0 10.4732
R173 VDD2.n41 VDD2.n40 9.45567
R174 VDD2.n18 VDD2.n17 9.45567
R175 VDD2.n40 VDD2.n39 9.3005
R176 VDD2.n25 VDD2.n24 9.3005
R177 VDD2.n34 VDD2.n33 9.3005
R178 VDD2.n32 VDD2.n31 9.3005
R179 VDD2.n17 VDD2.n16 9.3005
R180 VDD2.n2 VDD2.n1 9.3005
R181 VDD2.n11 VDD2.n10 9.3005
R182 VDD2.n9 VDD2.n8 9.3005
R183 VDD2.n45 VDD2.t5 8.18816
R184 VDD2.n45 VDD2.t8 8.18816
R185 VDD2.n43 VDD2.t4 8.18816
R186 VDD2.n43 VDD2.t3 8.18816
R187 VDD2.n21 VDD2.t6 8.18816
R188 VDD2.n21 VDD2.t0 8.18816
R189 VDD2.n19 VDD2.t1 8.18816
R190 VDD2.n19 VDD2.t9 8.18816
R191 VDD2.n32 VDD2.n28 3.78097
R192 VDD2.n9 VDD2.n5 3.78097
R193 VDD2.n41 VDD2.n23 3.49141
R194 VDD2.n18 VDD2.n0 3.49141
R195 VDD2.n39 VDD2.n38 2.71565
R196 VDD2.n16 VDD2.n15 2.71565
R197 VDD2.n44 VDD2.n42 2.59533
R198 VDD2.n35 VDD2.n25 1.93989
R199 VDD2.n12 VDD2.n2 1.93989
R200 VDD2.n34 VDD2.n27 1.16414
R201 VDD2.n11 VDD2.n4 1.16414
R202 VDD2 VDD2.n44 0.707397
R203 VDD2.n22 VDD2.n20 0.593861
R204 VDD2.n31 VDD2.n30 0.388379
R205 VDD2.n8 VDD2.n7 0.388379
R206 VDD2.n40 VDD2.n24 0.155672
R207 VDD2.n33 VDD2.n24 0.155672
R208 VDD2.n33 VDD2.n32 0.155672
R209 VDD2.n10 VDD2.n9 0.155672
R210 VDD2.n10 VDD2.n1 0.155672
R211 VDD2.n17 VDD2.n1 0.155672
R212 VTAIL.n88 VTAIL.n74 756.745
R213 VTAIL.n16 VTAIL.n2 756.745
R214 VTAIL.n68 VTAIL.n54 756.745
R215 VTAIL.n44 VTAIL.n30 756.745
R216 VTAIL.n81 VTAIL.n80 585
R217 VTAIL.n78 VTAIL.n77 585
R218 VTAIL.n87 VTAIL.n86 585
R219 VTAIL.n89 VTAIL.n88 585
R220 VTAIL.n9 VTAIL.n8 585
R221 VTAIL.n6 VTAIL.n5 585
R222 VTAIL.n15 VTAIL.n14 585
R223 VTAIL.n17 VTAIL.n16 585
R224 VTAIL.n69 VTAIL.n68 585
R225 VTAIL.n67 VTAIL.n66 585
R226 VTAIL.n58 VTAIL.n57 585
R227 VTAIL.n61 VTAIL.n60 585
R228 VTAIL.n45 VTAIL.n44 585
R229 VTAIL.n43 VTAIL.n42 585
R230 VTAIL.n34 VTAIL.n33 585
R231 VTAIL.n37 VTAIL.n36 585
R232 VTAIL.t11 VTAIL.n79 330.707
R233 VTAIL.t2 VTAIL.n7 330.707
R234 VTAIL.t5 VTAIL.n59 330.707
R235 VTAIL.t15 VTAIL.n35 330.707
R236 VTAIL.n80 VTAIL.n77 171.744
R237 VTAIL.n87 VTAIL.n77 171.744
R238 VTAIL.n88 VTAIL.n87 171.744
R239 VTAIL.n8 VTAIL.n5 171.744
R240 VTAIL.n15 VTAIL.n5 171.744
R241 VTAIL.n16 VTAIL.n15 171.744
R242 VTAIL.n68 VTAIL.n67 171.744
R243 VTAIL.n67 VTAIL.n57 171.744
R244 VTAIL.n60 VTAIL.n57 171.744
R245 VTAIL.n44 VTAIL.n43 171.744
R246 VTAIL.n43 VTAIL.n33 171.744
R247 VTAIL.n36 VTAIL.n33 171.744
R248 VTAIL.n53 VTAIL.n52 99.4107
R249 VTAIL.n51 VTAIL.n50 99.4107
R250 VTAIL.n29 VTAIL.n28 99.4107
R251 VTAIL.n27 VTAIL.n26 99.4107
R252 VTAIL.n95 VTAIL.n94 99.4106
R253 VTAIL.n1 VTAIL.n0 99.4106
R254 VTAIL.n23 VTAIL.n22 99.4106
R255 VTAIL.n25 VTAIL.n24 99.4106
R256 VTAIL.n80 VTAIL.t11 85.8723
R257 VTAIL.n8 VTAIL.t2 85.8723
R258 VTAIL.n60 VTAIL.t5 85.8723
R259 VTAIL.n36 VTAIL.t15 85.8723
R260 VTAIL.n93 VTAIL.n92 34.7066
R261 VTAIL.n21 VTAIL.n20 34.7066
R262 VTAIL.n73 VTAIL.n72 34.7066
R263 VTAIL.n49 VTAIL.n48 34.7066
R264 VTAIL.n27 VTAIL.n25 20.9789
R265 VTAIL.n93 VTAIL.n73 18.3841
R266 VTAIL.n81 VTAIL.n79 16.3201
R267 VTAIL.n9 VTAIL.n7 16.3201
R268 VTAIL.n61 VTAIL.n59 16.3201
R269 VTAIL.n37 VTAIL.n35 16.3201
R270 VTAIL.n82 VTAIL.n78 12.8005
R271 VTAIL.n10 VTAIL.n6 12.8005
R272 VTAIL.n62 VTAIL.n58 12.8005
R273 VTAIL.n38 VTAIL.n34 12.8005
R274 VTAIL.n86 VTAIL.n85 12.0247
R275 VTAIL.n14 VTAIL.n13 12.0247
R276 VTAIL.n66 VTAIL.n65 12.0247
R277 VTAIL.n42 VTAIL.n41 12.0247
R278 VTAIL.n89 VTAIL.n76 11.249
R279 VTAIL.n17 VTAIL.n4 11.249
R280 VTAIL.n69 VTAIL.n56 11.249
R281 VTAIL.n45 VTAIL.n32 11.249
R282 VTAIL.n90 VTAIL.n74 10.4732
R283 VTAIL.n18 VTAIL.n2 10.4732
R284 VTAIL.n70 VTAIL.n54 10.4732
R285 VTAIL.n46 VTAIL.n30 10.4732
R286 VTAIL.n92 VTAIL.n91 9.45567
R287 VTAIL.n20 VTAIL.n19 9.45567
R288 VTAIL.n72 VTAIL.n71 9.45567
R289 VTAIL.n48 VTAIL.n47 9.45567
R290 VTAIL.n91 VTAIL.n90 9.3005
R291 VTAIL.n76 VTAIL.n75 9.3005
R292 VTAIL.n85 VTAIL.n84 9.3005
R293 VTAIL.n83 VTAIL.n82 9.3005
R294 VTAIL.n19 VTAIL.n18 9.3005
R295 VTAIL.n4 VTAIL.n3 9.3005
R296 VTAIL.n13 VTAIL.n12 9.3005
R297 VTAIL.n11 VTAIL.n10 9.3005
R298 VTAIL.n71 VTAIL.n70 9.3005
R299 VTAIL.n56 VTAIL.n55 9.3005
R300 VTAIL.n65 VTAIL.n64 9.3005
R301 VTAIL.n63 VTAIL.n62 9.3005
R302 VTAIL.n47 VTAIL.n46 9.3005
R303 VTAIL.n32 VTAIL.n31 9.3005
R304 VTAIL.n41 VTAIL.n40 9.3005
R305 VTAIL.n39 VTAIL.n38 9.3005
R306 VTAIL.n94 VTAIL.t16 8.18816
R307 VTAIL.n94 VTAIL.t18 8.18816
R308 VTAIL.n0 VTAIL.t10 8.18816
R309 VTAIL.n0 VTAIL.t12 8.18816
R310 VTAIL.n22 VTAIL.t8 8.18816
R311 VTAIL.n22 VTAIL.t1 8.18816
R312 VTAIL.n24 VTAIL.t3 8.18816
R313 VTAIL.n24 VTAIL.t6 8.18816
R314 VTAIL.n52 VTAIL.t0 8.18816
R315 VTAIL.n52 VTAIL.t4 8.18816
R316 VTAIL.n50 VTAIL.t7 8.18816
R317 VTAIL.n50 VTAIL.t19 8.18816
R318 VTAIL.n28 VTAIL.t13 8.18816
R319 VTAIL.n28 VTAIL.t9 8.18816
R320 VTAIL.n26 VTAIL.t14 8.18816
R321 VTAIL.n26 VTAIL.t17 8.18816
R322 VTAIL.n83 VTAIL.n79 3.78097
R323 VTAIL.n11 VTAIL.n7 3.78097
R324 VTAIL.n63 VTAIL.n59 3.78097
R325 VTAIL.n39 VTAIL.n35 3.78097
R326 VTAIL.n92 VTAIL.n74 3.49141
R327 VTAIL.n20 VTAIL.n2 3.49141
R328 VTAIL.n72 VTAIL.n54 3.49141
R329 VTAIL.n48 VTAIL.n30 3.49141
R330 VTAIL.n90 VTAIL.n89 2.71565
R331 VTAIL.n18 VTAIL.n17 2.71565
R332 VTAIL.n70 VTAIL.n69 2.71565
R333 VTAIL.n46 VTAIL.n45 2.71565
R334 VTAIL.n29 VTAIL.n27 2.59533
R335 VTAIL.n49 VTAIL.n29 2.59533
R336 VTAIL.n53 VTAIL.n51 2.59533
R337 VTAIL.n73 VTAIL.n53 2.59533
R338 VTAIL.n25 VTAIL.n23 2.59533
R339 VTAIL.n23 VTAIL.n21 2.59533
R340 VTAIL.n95 VTAIL.n93 2.59533
R341 VTAIL VTAIL.n1 2.00481
R342 VTAIL.n86 VTAIL.n76 1.93989
R343 VTAIL.n14 VTAIL.n4 1.93989
R344 VTAIL.n66 VTAIL.n56 1.93989
R345 VTAIL.n42 VTAIL.n32 1.93989
R346 VTAIL.n51 VTAIL.n49 1.76774
R347 VTAIL.n21 VTAIL.n1 1.76774
R348 VTAIL.n85 VTAIL.n78 1.16414
R349 VTAIL.n13 VTAIL.n6 1.16414
R350 VTAIL.n65 VTAIL.n58 1.16414
R351 VTAIL.n41 VTAIL.n34 1.16414
R352 VTAIL VTAIL.n95 0.591017
R353 VTAIL.n82 VTAIL.n81 0.388379
R354 VTAIL.n10 VTAIL.n9 0.388379
R355 VTAIL.n62 VTAIL.n61 0.388379
R356 VTAIL.n38 VTAIL.n37 0.388379
R357 VTAIL.n84 VTAIL.n83 0.155672
R358 VTAIL.n84 VTAIL.n75 0.155672
R359 VTAIL.n91 VTAIL.n75 0.155672
R360 VTAIL.n12 VTAIL.n11 0.155672
R361 VTAIL.n12 VTAIL.n3 0.155672
R362 VTAIL.n19 VTAIL.n3 0.155672
R363 VTAIL.n71 VTAIL.n55 0.155672
R364 VTAIL.n64 VTAIL.n55 0.155672
R365 VTAIL.n64 VTAIL.n63 0.155672
R366 VTAIL.n47 VTAIL.n31 0.155672
R367 VTAIL.n40 VTAIL.n31 0.155672
R368 VTAIL.n40 VTAIL.n39 0.155672
R369 VP.n27 VP.n26 161.3
R370 VP.n28 VP.n23 161.3
R371 VP.n30 VP.n29 161.3
R372 VP.n31 VP.n22 161.3
R373 VP.n33 VP.n32 161.3
R374 VP.n34 VP.n21 161.3
R375 VP.n36 VP.n35 161.3
R376 VP.n37 VP.n20 161.3
R377 VP.n39 VP.n38 161.3
R378 VP.n40 VP.n19 161.3
R379 VP.n42 VP.n41 161.3
R380 VP.n43 VP.n18 161.3
R381 VP.n45 VP.n44 161.3
R382 VP.n47 VP.n46 161.3
R383 VP.n48 VP.n16 161.3
R384 VP.n50 VP.n49 161.3
R385 VP.n51 VP.n15 161.3
R386 VP.n53 VP.n52 161.3
R387 VP.n54 VP.n14 161.3
R388 VP.n96 VP.n0 161.3
R389 VP.n95 VP.n94 161.3
R390 VP.n93 VP.n1 161.3
R391 VP.n92 VP.n91 161.3
R392 VP.n90 VP.n2 161.3
R393 VP.n89 VP.n88 161.3
R394 VP.n87 VP.n86 161.3
R395 VP.n85 VP.n4 161.3
R396 VP.n84 VP.n83 161.3
R397 VP.n82 VP.n5 161.3
R398 VP.n81 VP.n80 161.3
R399 VP.n79 VP.n6 161.3
R400 VP.n78 VP.n77 161.3
R401 VP.n76 VP.n7 161.3
R402 VP.n75 VP.n74 161.3
R403 VP.n73 VP.n8 161.3
R404 VP.n72 VP.n71 161.3
R405 VP.n70 VP.n9 161.3
R406 VP.n69 VP.n68 161.3
R407 VP.n66 VP.n10 161.3
R408 VP.n65 VP.n64 161.3
R409 VP.n63 VP.n11 161.3
R410 VP.n62 VP.n61 161.3
R411 VP.n60 VP.n12 161.3
R412 VP.n59 VP.n58 161.3
R413 VP.n57 VP.n13 109.778
R414 VP.n98 VP.n97 109.778
R415 VP.n56 VP.n55 109.778
R416 VP.n25 VP.n24 72.9374
R417 VP.n24 VP.t2 65.9996
R418 VP.n57 VP.n56 47.367
R419 VP.n61 VP.n11 41.9503
R420 VP.n91 VP.n1 41.9503
R421 VP.n49 VP.n15 41.9503
R422 VP.n73 VP.n72 40.979
R423 VP.n84 VP.n5 40.979
R424 VP.n42 VP.n19 40.979
R425 VP.n31 VP.n30 40.979
R426 VP.n74 VP.n73 40.0078
R427 VP.n80 VP.n5 40.0078
R428 VP.n38 VP.n19 40.0078
R429 VP.n32 VP.n31 40.0078
R430 VP.n65 VP.n11 39.0365
R431 VP.n91 VP.n90 39.0365
R432 VP.n49 VP.n48 39.0365
R433 VP.n78 VP.t0 35.7009
R434 VP.n13 VP.t4 35.7009
R435 VP.n67 VP.t9 35.7009
R436 VP.n3 VP.t3 35.7009
R437 VP.n97 VP.t6 35.7009
R438 VP.n36 VP.t1 35.7009
R439 VP.n55 VP.t8 35.7009
R440 VP.n17 VP.t5 35.7009
R441 VP.n25 VP.t7 35.7009
R442 VP.n60 VP.n59 24.4675
R443 VP.n61 VP.n60 24.4675
R444 VP.n66 VP.n65 24.4675
R445 VP.n68 VP.n9 24.4675
R446 VP.n72 VP.n9 24.4675
R447 VP.n74 VP.n7 24.4675
R448 VP.n78 VP.n7 24.4675
R449 VP.n79 VP.n78 24.4675
R450 VP.n80 VP.n79 24.4675
R451 VP.n85 VP.n84 24.4675
R452 VP.n86 VP.n85 24.4675
R453 VP.n90 VP.n89 24.4675
R454 VP.n95 VP.n1 24.4675
R455 VP.n96 VP.n95 24.4675
R456 VP.n53 VP.n15 24.4675
R457 VP.n54 VP.n53 24.4675
R458 VP.n43 VP.n42 24.4675
R459 VP.n44 VP.n43 24.4675
R460 VP.n48 VP.n47 24.4675
R461 VP.n32 VP.n21 24.4675
R462 VP.n36 VP.n21 24.4675
R463 VP.n37 VP.n36 24.4675
R464 VP.n38 VP.n37 24.4675
R465 VP.n26 VP.n23 24.4675
R466 VP.n30 VP.n23 24.4675
R467 VP.n67 VP.n66 23.9782
R468 VP.n89 VP.n3 23.9782
R469 VP.n47 VP.n17 23.9782
R470 VP.n27 VP.n24 7.44194
R471 VP.n59 VP.n13 0.97918
R472 VP.n97 VP.n96 0.97918
R473 VP.n55 VP.n54 0.97918
R474 VP.n68 VP.n67 0.48984
R475 VP.n86 VP.n3 0.48984
R476 VP.n44 VP.n17 0.48984
R477 VP.n26 VP.n25 0.48984
R478 VP.n56 VP.n14 0.278367
R479 VP.n58 VP.n57 0.278367
R480 VP.n98 VP.n0 0.278367
R481 VP.n28 VP.n27 0.189894
R482 VP.n29 VP.n28 0.189894
R483 VP.n29 VP.n22 0.189894
R484 VP.n33 VP.n22 0.189894
R485 VP.n34 VP.n33 0.189894
R486 VP.n35 VP.n34 0.189894
R487 VP.n35 VP.n20 0.189894
R488 VP.n39 VP.n20 0.189894
R489 VP.n40 VP.n39 0.189894
R490 VP.n41 VP.n40 0.189894
R491 VP.n41 VP.n18 0.189894
R492 VP.n45 VP.n18 0.189894
R493 VP.n46 VP.n45 0.189894
R494 VP.n46 VP.n16 0.189894
R495 VP.n50 VP.n16 0.189894
R496 VP.n51 VP.n50 0.189894
R497 VP.n52 VP.n51 0.189894
R498 VP.n52 VP.n14 0.189894
R499 VP.n58 VP.n12 0.189894
R500 VP.n62 VP.n12 0.189894
R501 VP.n63 VP.n62 0.189894
R502 VP.n64 VP.n63 0.189894
R503 VP.n64 VP.n10 0.189894
R504 VP.n69 VP.n10 0.189894
R505 VP.n70 VP.n69 0.189894
R506 VP.n71 VP.n70 0.189894
R507 VP.n71 VP.n8 0.189894
R508 VP.n75 VP.n8 0.189894
R509 VP.n76 VP.n75 0.189894
R510 VP.n77 VP.n76 0.189894
R511 VP.n77 VP.n6 0.189894
R512 VP.n81 VP.n6 0.189894
R513 VP.n82 VP.n81 0.189894
R514 VP.n83 VP.n82 0.189894
R515 VP.n83 VP.n4 0.189894
R516 VP.n87 VP.n4 0.189894
R517 VP.n88 VP.n87 0.189894
R518 VP.n88 VP.n2 0.189894
R519 VP.n92 VP.n2 0.189894
R520 VP.n93 VP.n92 0.189894
R521 VP.n94 VP.n93 0.189894
R522 VP.n94 VP.n0 0.189894
R523 VP VP.n98 0.153454
R524 VDD1.n14 VDD1.n0 756.745
R525 VDD1.n35 VDD1.n21 756.745
R526 VDD1.n15 VDD1.n14 585
R527 VDD1.n13 VDD1.n12 585
R528 VDD1.n4 VDD1.n3 585
R529 VDD1.n7 VDD1.n6 585
R530 VDD1.n28 VDD1.n27 585
R531 VDD1.n25 VDD1.n24 585
R532 VDD1.n34 VDD1.n33 585
R533 VDD1.n36 VDD1.n35 585
R534 VDD1.t7 VDD1.n5 330.707
R535 VDD1.t5 VDD1.n26 330.707
R536 VDD1.n14 VDD1.n13 171.744
R537 VDD1.n13 VDD1.n3 171.744
R538 VDD1.n6 VDD1.n3 171.744
R539 VDD1.n27 VDD1.n24 171.744
R540 VDD1.n34 VDD1.n24 171.744
R541 VDD1.n35 VDD1.n34 171.744
R542 VDD1.n43 VDD1.n42 117.981
R543 VDD1.n20 VDD1.n19 116.09
R544 VDD1.n45 VDD1.n44 116.09
R545 VDD1.n41 VDD1.n40 116.09
R546 VDD1.n6 VDD1.t7 85.8723
R547 VDD1.n27 VDD1.t5 85.8723
R548 VDD1.n20 VDD1.n18 53.9802
R549 VDD1.n41 VDD1.n39 53.9802
R550 VDD1.n45 VDD1.n43 41.3436
R551 VDD1.n7 VDD1.n5 16.3201
R552 VDD1.n28 VDD1.n26 16.3201
R553 VDD1.n8 VDD1.n4 12.8005
R554 VDD1.n29 VDD1.n25 12.8005
R555 VDD1.n12 VDD1.n11 12.0247
R556 VDD1.n33 VDD1.n32 12.0247
R557 VDD1.n15 VDD1.n2 11.249
R558 VDD1.n36 VDD1.n23 11.249
R559 VDD1.n16 VDD1.n0 10.4732
R560 VDD1.n37 VDD1.n21 10.4732
R561 VDD1.n18 VDD1.n17 9.45567
R562 VDD1.n39 VDD1.n38 9.45567
R563 VDD1.n17 VDD1.n16 9.3005
R564 VDD1.n2 VDD1.n1 9.3005
R565 VDD1.n11 VDD1.n10 9.3005
R566 VDD1.n9 VDD1.n8 9.3005
R567 VDD1.n38 VDD1.n37 9.3005
R568 VDD1.n23 VDD1.n22 9.3005
R569 VDD1.n32 VDD1.n31 9.3005
R570 VDD1.n30 VDD1.n29 9.3005
R571 VDD1.n44 VDD1.t4 8.18816
R572 VDD1.n44 VDD1.t1 8.18816
R573 VDD1.n19 VDD1.t2 8.18816
R574 VDD1.n19 VDD1.t8 8.18816
R575 VDD1.n42 VDD1.t6 8.18816
R576 VDD1.n42 VDD1.t3 8.18816
R577 VDD1.n40 VDD1.t0 8.18816
R578 VDD1.n40 VDD1.t9 8.18816
R579 VDD1.n9 VDD1.n5 3.78097
R580 VDD1.n30 VDD1.n26 3.78097
R581 VDD1.n18 VDD1.n0 3.49141
R582 VDD1.n39 VDD1.n21 3.49141
R583 VDD1.n16 VDD1.n15 2.71565
R584 VDD1.n37 VDD1.n36 2.71565
R585 VDD1.n12 VDD1.n2 1.93989
R586 VDD1.n33 VDD1.n23 1.93989
R587 VDD1 VDD1.n45 1.88843
R588 VDD1.n11 VDD1.n4 1.16414
R589 VDD1.n32 VDD1.n25 1.16414
R590 VDD1 VDD1.n20 0.707397
R591 VDD1.n43 VDD1.n41 0.593861
R592 VDD1.n8 VDD1.n7 0.388379
R593 VDD1.n29 VDD1.n28 0.388379
R594 VDD1.n17 VDD1.n1 0.155672
R595 VDD1.n10 VDD1.n1 0.155672
R596 VDD1.n10 VDD1.n9 0.155672
R597 VDD1.n31 VDD1.n30 0.155672
R598 VDD1.n31 VDD1.n22 0.155672
R599 VDD1.n38 VDD1.n22 0.155672
R600 B.n525 B.n60 585
R601 B.n527 B.n526 585
R602 B.n528 B.n59 585
R603 B.n530 B.n529 585
R604 B.n531 B.n58 585
R605 B.n533 B.n532 585
R606 B.n534 B.n57 585
R607 B.n536 B.n535 585
R608 B.n537 B.n56 585
R609 B.n539 B.n538 585
R610 B.n540 B.n55 585
R611 B.n542 B.n541 585
R612 B.n543 B.n54 585
R613 B.n545 B.n544 585
R614 B.n546 B.n53 585
R615 B.n548 B.n547 585
R616 B.n549 B.n49 585
R617 B.n551 B.n550 585
R618 B.n552 B.n48 585
R619 B.n554 B.n553 585
R620 B.n555 B.n47 585
R621 B.n557 B.n556 585
R622 B.n558 B.n46 585
R623 B.n560 B.n559 585
R624 B.n561 B.n45 585
R625 B.n563 B.n562 585
R626 B.n564 B.n44 585
R627 B.n566 B.n565 585
R628 B.n568 B.n41 585
R629 B.n570 B.n569 585
R630 B.n571 B.n40 585
R631 B.n573 B.n572 585
R632 B.n574 B.n39 585
R633 B.n576 B.n575 585
R634 B.n577 B.n38 585
R635 B.n579 B.n578 585
R636 B.n580 B.n37 585
R637 B.n582 B.n581 585
R638 B.n583 B.n36 585
R639 B.n585 B.n584 585
R640 B.n586 B.n35 585
R641 B.n588 B.n587 585
R642 B.n589 B.n34 585
R643 B.n591 B.n590 585
R644 B.n592 B.n33 585
R645 B.n594 B.n593 585
R646 B.n524 B.n523 585
R647 B.n522 B.n61 585
R648 B.n521 B.n520 585
R649 B.n519 B.n62 585
R650 B.n518 B.n517 585
R651 B.n516 B.n63 585
R652 B.n515 B.n514 585
R653 B.n513 B.n64 585
R654 B.n512 B.n511 585
R655 B.n510 B.n65 585
R656 B.n509 B.n508 585
R657 B.n507 B.n66 585
R658 B.n506 B.n505 585
R659 B.n504 B.n67 585
R660 B.n503 B.n502 585
R661 B.n501 B.n68 585
R662 B.n500 B.n499 585
R663 B.n498 B.n69 585
R664 B.n497 B.n496 585
R665 B.n495 B.n70 585
R666 B.n494 B.n493 585
R667 B.n492 B.n71 585
R668 B.n491 B.n490 585
R669 B.n489 B.n72 585
R670 B.n488 B.n487 585
R671 B.n486 B.n73 585
R672 B.n485 B.n484 585
R673 B.n483 B.n74 585
R674 B.n482 B.n481 585
R675 B.n480 B.n75 585
R676 B.n479 B.n478 585
R677 B.n477 B.n76 585
R678 B.n476 B.n475 585
R679 B.n474 B.n77 585
R680 B.n473 B.n472 585
R681 B.n471 B.n78 585
R682 B.n470 B.n469 585
R683 B.n468 B.n79 585
R684 B.n467 B.n466 585
R685 B.n465 B.n80 585
R686 B.n464 B.n463 585
R687 B.n462 B.n81 585
R688 B.n461 B.n460 585
R689 B.n459 B.n82 585
R690 B.n458 B.n457 585
R691 B.n456 B.n83 585
R692 B.n455 B.n454 585
R693 B.n453 B.n84 585
R694 B.n452 B.n451 585
R695 B.n450 B.n85 585
R696 B.n449 B.n448 585
R697 B.n447 B.n86 585
R698 B.n446 B.n445 585
R699 B.n444 B.n87 585
R700 B.n443 B.n442 585
R701 B.n441 B.n88 585
R702 B.n440 B.n439 585
R703 B.n438 B.n89 585
R704 B.n437 B.n436 585
R705 B.n435 B.n90 585
R706 B.n434 B.n433 585
R707 B.n432 B.n91 585
R708 B.n431 B.n430 585
R709 B.n429 B.n92 585
R710 B.n428 B.n427 585
R711 B.n426 B.n93 585
R712 B.n425 B.n424 585
R713 B.n423 B.n94 585
R714 B.n422 B.n421 585
R715 B.n420 B.n95 585
R716 B.n419 B.n418 585
R717 B.n417 B.n96 585
R718 B.n416 B.n415 585
R719 B.n414 B.n97 585
R720 B.n413 B.n412 585
R721 B.n411 B.n98 585
R722 B.n410 B.n409 585
R723 B.n408 B.n99 585
R724 B.n407 B.n406 585
R725 B.n405 B.n100 585
R726 B.n404 B.n403 585
R727 B.n402 B.n101 585
R728 B.n401 B.n400 585
R729 B.n399 B.n102 585
R730 B.n398 B.n397 585
R731 B.n396 B.n103 585
R732 B.n395 B.n394 585
R733 B.n393 B.n104 585
R734 B.n392 B.n391 585
R735 B.n390 B.n105 585
R736 B.n389 B.n388 585
R737 B.n387 B.n106 585
R738 B.n386 B.n385 585
R739 B.n384 B.n107 585
R740 B.n383 B.n382 585
R741 B.n381 B.n108 585
R742 B.n380 B.n379 585
R743 B.n378 B.n109 585
R744 B.n377 B.n376 585
R745 B.n375 B.n110 585
R746 B.n374 B.n373 585
R747 B.n372 B.n111 585
R748 B.n371 B.n370 585
R749 B.n369 B.n112 585
R750 B.n368 B.n367 585
R751 B.n366 B.n113 585
R752 B.n365 B.n364 585
R753 B.n363 B.n114 585
R754 B.n362 B.n361 585
R755 B.n360 B.n115 585
R756 B.n359 B.n358 585
R757 B.n357 B.n116 585
R758 B.n356 B.n355 585
R759 B.n354 B.n117 585
R760 B.n353 B.n352 585
R761 B.n351 B.n118 585
R762 B.n350 B.n349 585
R763 B.n348 B.n119 585
R764 B.n347 B.n346 585
R765 B.n345 B.n120 585
R766 B.n344 B.n343 585
R767 B.n342 B.n121 585
R768 B.n341 B.n340 585
R769 B.n270 B.n149 585
R770 B.n272 B.n271 585
R771 B.n273 B.n148 585
R772 B.n275 B.n274 585
R773 B.n276 B.n147 585
R774 B.n278 B.n277 585
R775 B.n279 B.n146 585
R776 B.n281 B.n280 585
R777 B.n282 B.n145 585
R778 B.n284 B.n283 585
R779 B.n285 B.n144 585
R780 B.n287 B.n286 585
R781 B.n288 B.n143 585
R782 B.n290 B.n289 585
R783 B.n291 B.n142 585
R784 B.n293 B.n292 585
R785 B.n294 B.n141 585
R786 B.n296 B.n295 585
R787 B.n298 B.n138 585
R788 B.n300 B.n299 585
R789 B.n301 B.n137 585
R790 B.n303 B.n302 585
R791 B.n304 B.n136 585
R792 B.n306 B.n305 585
R793 B.n307 B.n135 585
R794 B.n309 B.n308 585
R795 B.n310 B.n134 585
R796 B.n312 B.n311 585
R797 B.n314 B.n313 585
R798 B.n315 B.n130 585
R799 B.n317 B.n316 585
R800 B.n318 B.n129 585
R801 B.n320 B.n319 585
R802 B.n321 B.n128 585
R803 B.n323 B.n322 585
R804 B.n324 B.n127 585
R805 B.n326 B.n325 585
R806 B.n327 B.n126 585
R807 B.n329 B.n328 585
R808 B.n330 B.n125 585
R809 B.n332 B.n331 585
R810 B.n333 B.n124 585
R811 B.n335 B.n334 585
R812 B.n336 B.n123 585
R813 B.n338 B.n337 585
R814 B.n339 B.n122 585
R815 B.n269 B.n268 585
R816 B.n267 B.n150 585
R817 B.n266 B.n265 585
R818 B.n264 B.n151 585
R819 B.n263 B.n262 585
R820 B.n261 B.n152 585
R821 B.n260 B.n259 585
R822 B.n258 B.n153 585
R823 B.n257 B.n256 585
R824 B.n255 B.n154 585
R825 B.n254 B.n253 585
R826 B.n252 B.n155 585
R827 B.n251 B.n250 585
R828 B.n249 B.n156 585
R829 B.n248 B.n247 585
R830 B.n246 B.n157 585
R831 B.n245 B.n244 585
R832 B.n243 B.n158 585
R833 B.n242 B.n241 585
R834 B.n240 B.n159 585
R835 B.n239 B.n238 585
R836 B.n237 B.n160 585
R837 B.n236 B.n235 585
R838 B.n234 B.n161 585
R839 B.n233 B.n232 585
R840 B.n231 B.n162 585
R841 B.n230 B.n229 585
R842 B.n228 B.n163 585
R843 B.n227 B.n226 585
R844 B.n225 B.n164 585
R845 B.n224 B.n223 585
R846 B.n222 B.n165 585
R847 B.n221 B.n220 585
R848 B.n219 B.n166 585
R849 B.n218 B.n217 585
R850 B.n216 B.n167 585
R851 B.n215 B.n214 585
R852 B.n213 B.n168 585
R853 B.n212 B.n211 585
R854 B.n210 B.n169 585
R855 B.n209 B.n208 585
R856 B.n207 B.n170 585
R857 B.n206 B.n205 585
R858 B.n204 B.n171 585
R859 B.n203 B.n202 585
R860 B.n201 B.n172 585
R861 B.n200 B.n199 585
R862 B.n198 B.n173 585
R863 B.n197 B.n196 585
R864 B.n195 B.n174 585
R865 B.n194 B.n193 585
R866 B.n192 B.n175 585
R867 B.n191 B.n190 585
R868 B.n189 B.n176 585
R869 B.n188 B.n187 585
R870 B.n186 B.n177 585
R871 B.n185 B.n184 585
R872 B.n183 B.n178 585
R873 B.n182 B.n181 585
R874 B.n180 B.n179 585
R875 B.n2 B.n0 585
R876 B.n685 B.n1 585
R877 B.n684 B.n683 585
R878 B.n682 B.n3 585
R879 B.n681 B.n680 585
R880 B.n679 B.n4 585
R881 B.n678 B.n677 585
R882 B.n676 B.n5 585
R883 B.n675 B.n674 585
R884 B.n673 B.n6 585
R885 B.n672 B.n671 585
R886 B.n670 B.n7 585
R887 B.n669 B.n668 585
R888 B.n667 B.n8 585
R889 B.n666 B.n665 585
R890 B.n664 B.n9 585
R891 B.n663 B.n662 585
R892 B.n661 B.n10 585
R893 B.n660 B.n659 585
R894 B.n658 B.n11 585
R895 B.n657 B.n656 585
R896 B.n655 B.n12 585
R897 B.n654 B.n653 585
R898 B.n652 B.n13 585
R899 B.n651 B.n650 585
R900 B.n649 B.n14 585
R901 B.n648 B.n647 585
R902 B.n646 B.n15 585
R903 B.n645 B.n644 585
R904 B.n643 B.n16 585
R905 B.n642 B.n641 585
R906 B.n640 B.n17 585
R907 B.n639 B.n638 585
R908 B.n637 B.n18 585
R909 B.n636 B.n635 585
R910 B.n634 B.n19 585
R911 B.n633 B.n632 585
R912 B.n631 B.n20 585
R913 B.n630 B.n629 585
R914 B.n628 B.n21 585
R915 B.n627 B.n626 585
R916 B.n625 B.n22 585
R917 B.n624 B.n623 585
R918 B.n622 B.n23 585
R919 B.n621 B.n620 585
R920 B.n619 B.n24 585
R921 B.n618 B.n617 585
R922 B.n616 B.n25 585
R923 B.n615 B.n614 585
R924 B.n613 B.n26 585
R925 B.n612 B.n611 585
R926 B.n610 B.n27 585
R927 B.n609 B.n608 585
R928 B.n607 B.n28 585
R929 B.n606 B.n605 585
R930 B.n604 B.n29 585
R931 B.n603 B.n602 585
R932 B.n601 B.n30 585
R933 B.n600 B.n599 585
R934 B.n598 B.n31 585
R935 B.n597 B.n596 585
R936 B.n595 B.n32 585
R937 B.n687 B.n686 585
R938 B.n270 B.n269 502.111
R939 B.n595 B.n594 502.111
R940 B.n341 B.n122 502.111
R941 B.n523 B.n60 502.111
R942 B.n131 B.t11 293.618
R943 B.n50 B.t1 293.618
R944 B.n139 B.t5 293.618
R945 B.n42 B.t7 293.618
R946 B.n131 B.t9 244.529
R947 B.n50 B.t0 244.529
R948 B.n139 B.t3 244.208
R949 B.n42 B.t6 244.208
R950 B.n132 B.t10 235.242
R951 B.n51 B.t2 235.242
R952 B.n140 B.t4 235.242
R953 B.n43 B.t8 235.242
R954 B.n269 B.n150 163.367
R955 B.n265 B.n150 163.367
R956 B.n265 B.n264 163.367
R957 B.n264 B.n263 163.367
R958 B.n263 B.n152 163.367
R959 B.n259 B.n152 163.367
R960 B.n259 B.n258 163.367
R961 B.n258 B.n257 163.367
R962 B.n257 B.n154 163.367
R963 B.n253 B.n154 163.367
R964 B.n253 B.n252 163.367
R965 B.n252 B.n251 163.367
R966 B.n251 B.n156 163.367
R967 B.n247 B.n156 163.367
R968 B.n247 B.n246 163.367
R969 B.n246 B.n245 163.367
R970 B.n245 B.n158 163.367
R971 B.n241 B.n158 163.367
R972 B.n241 B.n240 163.367
R973 B.n240 B.n239 163.367
R974 B.n239 B.n160 163.367
R975 B.n235 B.n160 163.367
R976 B.n235 B.n234 163.367
R977 B.n234 B.n233 163.367
R978 B.n233 B.n162 163.367
R979 B.n229 B.n162 163.367
R980 B.n229 B.n228 163.367
R981 B.n228 B.n227 163.367
R982 B.n227 B.n164 163.367
R983 B.n223 B.n164 163.367
R984 B.n223 B.n222 163.367
R985 B.n222 B.n221 163.367
R986 B.n221 B.n166 163.367
R987 B.n217 B.n166 163.367
R988 B.n217 B.n216 163.367
R989 B.n216 B.n215 163.367
R990 B.n215 B.n168 163.367
R991 B.n211 B.n168 163.367
R992 B.n211 B.n210 163.367
R993 B.n210 B.n209 163.367
R994 B.n209 B.n170 163.367
R995 B.n205 B.n170 163.367
R996 B.n205 B.n204 163.367
R997 B.n204 B.n203 163.367
R998 B.n203 B.n172 163.367
R999 B.n199 B.n172 163.367
R1000 B.n199 B.n198 163.367
R1001 B.n198 B.n197 163.367
R1002 B.n197 B.n174 163.367
R1003 B.n193 B.n174 163.367
R1004 B.n193 B.n192 163.367
R1005 B.n192 B.n191 163.367
R1006 B.n191 B.n176 163.367
R1007 B.n187 B.n176 163.367
R1008 B.n187 B.n186 163.367
R1009 B.n186 B.n185 163.367
R1010 B.n185 B.n178 163.367
R1011 B.n181 B.n178 163.367
R1012 B.n181 B.n180 163.367
R1013 B.n180 B.n2 163.367
R1014 B.n686 B.n2 163.367
R1015 B.n686 B.n685 163.367
R1016 B.n685 B.n684 163.367
R1017 B.n684 B.n3 163.367
R1018 B.n680 B.n3 163.367
R1019 B.n680 B.n679 163.367
R1020 B.n679 B.n678 163.367
R1021 B.n678 B.n5 163.367
R1022 B.n674 B.n5 163.367
R1023 B.n674 B.n673 163.367
R1024 B.n673 B.n672 163.367
R1025 B.n672 B.n7 163.367
R1026 B.n668 B.n7 163.367
R1027 B.n668 B.n667 163.367
R1028 B.n667 B.n666 163.367
R1029 B.n666 B.n9 163.367
R1030 B.n662 B.n9 163.367
R1031 B.n662 B.n661 163.367
R1032 B.n661 B.n660 163.367
R1033 B.n660 B.n11 163.367
R1034 B.n656 B.n11 163.367
R1035 B.n656 B.n655 163.367
R1036 B.n655 B.n654 163.367
R1037 B.n654 B.n13 163.367
R1038 B.n650 B.n13 163.367
R1039 B.n650 B.n649 163.367
R1040 B.n649 B.n648 163.367
R1041 B.n648 B.n15 163.367
R1042 B.n644 B.n15 163.367
R1043 B.n644 B.n643 163.367
R1044 B.n643 B.n642 163.367
R1045 B.n642 B.n17 163.367
R1046 B.n638 B.n17 163.367
R1047 B.n638 B.n637 163.367
R1048 B.n637 B.n636 163.367
R1049 B.n636 B.n19 163.367
R1050 B.n632 B.n19 163.367
R1051 B.n632 B.n631 163.367
R1052 B.n631 B.n630 163.367
R1053 B.n630 B.n21 163.367
R1054 B.n626 B.n21 163.367
R1055 B.n626 B.n625 163.367
R1056 B.n625 B.n624 163.367
R1057 B.n624 B.n23 163.367
R1058 B.n620 B.n23 163.367
R1059 B.n620 B.n619 163.367
R1060 B.n619 B.n618 163.367
R1061 B.n618 B.n25 163.367
R1062 B.n614 B.n25 163.367
R1063 B.n614 B.n613 163.367
R1064 B.n613 B.n612 163.367
R1065 B.n612 B.n27 163.367
R1066 B.n608 B.n27 163.367
R1067 B.n608 B.n607 163.367
R1068 B.n607 B.n606 163.367
R1069 B.n606 B.n29 163.367
R1070 B.n602 B.n29 163.367
R1071 B.n602 B.n601 163.367
R1072 B.n601 B.n600 163.367
R1073 B.n600 B.n31 163.367
R1074 B.n596 B.n31 163.367
R1075 B.n596 B.n595 163.367
R1076 B.n271 B.n270 163.367
R1077 B.n271 B.n148 163.367
R1078 B.n275 B.n148 163.367
R1079 B.n276 B.n275 163.367
R1080 B.n277 B.n276 163.367
R1081 B.n277 B.n146 163.367
R1082 B.n281 B.n146 163.367
R1083 B.n282 B.n281 163.367
R1084 B.n283 B.n282 163.367
R1085 B.n283 B.n144 163.367
R1086 B.n287 B.n144 163.367
R1087 B.n288 B.n287 163.367
R1088 B.n289 B.n288 163.367
R1089 B.n289 B.n142 163.367
R1090 B.n293 B.n142 163.367
R1091 B.n294 B.n293 163.367
R1092 B.n295 B.n294 163.367
R1093 B.n295 B.n138 163.367
R1094 B.n300 B.n138 163.367
R1095 B.n301 B.n300 163.367
R1096 B.n302 B.n301 163.367
R1097 B.n302 B.n136 163.367
R1098 B.n306 B.n136 163.367
R1099 B.n307 B.n306 163.367
R1100 B.n308 B.n307 163.367
R1101 B.n308 B.n134 163.367
R1102 B.n312 B.n134 163.367
R1103 B.n313 B.n312 163.367
R1104 B.n313 B.n130 163.367
R1105 B.n317 B.n130 163.367
R1106 B.n318 B.n317 163.367
R1107 B.n319 B.n318 163.367
R1108 B.n319 B.n128 163.367
R1109 B.n323 B.n128 163.367
R1110 B.n324 B.n323 163.367
R1111 B.n325 B.n324 163.367
R1112 B.n325 B.n126 163.367
R1113 B.n329 B.n126 163.367
R1114 B.n330 B.n329 163.367
R1115 B.n331 B.n330 163.367
R1116 B.n331 B.n124 163.367
R1117 B.n335 B.n124 163.367
R1118 B.n336 B.n335 163.367
R1119 B.n337 B.n336 163.367
R1120 B.n337 B.n122 163.367
R1121 B.n342 B.n341 163.367
R1122 B.n343 B.n342 163.367
R1123 B.n343 B.n120 163.367
R1124 B.n347 B.n120 163.367
R1125 B.n348 B.n347 163.367
R1126 B.n349 B.n348 163.367
R1127 B.n349 B.n118 163.367
R1128 B.n353 B.n118 163.367
R1129 B.n354 B.n353 163.367
R1130 B.n355 B.n354 163.367
R1131 B.n355 B.n116 163.367
R1132 B.n359 B.n116 163.367
R1133 B.n360 B.n359 163.367
R1134 B.n361 B.n360 163.367
R1135 B.n361 B.n114 163.367
R1136 B.n365 B.n114 163.367
R1137 B.n366 B.n365 163.367
R1138 B.n367 B.n366 163.367
R1139 B.n367 B.n112 163.367
R1140 B.n371 B.n112 163.367
R1141 B.n372 B.n371 163.367
R1142 B.n373 B.n372 163.367
R1143 B.n373 B.n110 163.367
R1144 B.n377 B.n110 163.367
R1145 B.n378 B.n377 163.367
R1146 B.n379 B.n378 163.367
R1147 B.n379 B.n108 163.367
R1148 B.n383 B.n108 163.367
R1149 B.n384 B.n383 163.367
R1150 B.n385 B.n384 163.367
R1151 B.n385 B.n106 163.367
R1152 B.n389 B.n106 163.367
R1153 B.n390 B.n389 163.367
R1154 B.n391 B.n390 163.367
R1155 B.n391 B.n104 163.367
R1156 B.n395 B.n104 163.367
R1157 B.n396 B.n395 163.367
R1158 B.n397 B.n396 163.367
R1159 B.n397 B.n102 163.367
R1160 B.n401 B.n102 163.367
R1161 B.n402 B.n401 163.367
R1162 B.n403 B.n402 163.367
R1163 B.n403 B.n100 163.367
R1164 B.n407 B.n100 163.367
R1165 B.n408 B.n407 163.367
R1166 B.n409 B.n408 163.367
R1167 B.n409 B.n98 163.367
R1168 B.n413 B.n98 163.367
R1169 B.n414 B.n413 163.367
R1170 B.n415 B.n414 163.367
R1171 B.n415 B.n96 163.367
R1172 B.n419 B.n96 163.367
R1173 B.n420 B.n419 163.367
R1174 B.n421 B.n420 163.367
R1175 B.n421 B.n94 163.367
R1176 B.n425 B.n94 163.367
R1177 B.n426 B.n425 163.367
R1178 B.n427 B.n426 163.367
R1179 B.n427 B.n92 163.367
R1180 B.n431 B.n92 163.367
R1181 B.n432 B.n431 163.367
R1182 B.n433 B.n432 163.367
R1183 B.n433 B.n90 163.367
R1184 B.n437 B.n90 163.367
R1185 B.n438 B.n437 163.367
R1186 B.n439 B.n438 163.367
R1187 B.n439 B.n88 163.367
R1188 B.n443 B.n88 163.367
R1189 B.n444 B.n443 163.367
R1190 B.n445 B.n444 163.367
R1191 B.n445 B.n86 163.367
R1192 B.n449 B.n86 163.367
R1193 B.n450 B.n449 163.367
R1194 B.n451 B.n450 163.367
R1195 B.n451 B.n84 163.367
R1196 B.n455 B.n84 163.367
R1197 B.n456 B.n455 163.367
R1198 B.n457 B.n456 163.367
R1199 B.n457 B.n82 163.367
R1200 B.n461 B.n82 163.367
R1201 B.n462 B.n461 163.367
R1202 B.n463 B.n462 163.367
R1203 B.n463 B.n80 163.367
R1204 B.n467 B.n80 163.367
R1205 B.n468 B.n467 163.367
R1206 B.n469 B.n468 163.367
R1207 B.n469 B.n78 163.367
R1208 B.n473 B.n78 163.367
R1209 B.n474 B.n473 163.367
R1210 B.n475 B.n474 163.367
R1211 B.n475 B.n76 163.367
R1212 B.n479 B.n76 163.367
R1213 B.n480 B.n479 163.367
R1214 B.n481 B.n480 163.367
R1215 B.n481 B.n74 163.367
R1216 B.n485 B.n74 163.367
R1217 B.n486 B.n485 163.367
R1218 B.n487 B.n486 163.367
R1219 B.n487 B.n72 163.367
R1220 B.n491 B.n72 163.367
R1221 B.n492 B.n491 163.367
R1222 B.n493 B.n492 163.367
R1223 B.n493 B.n70 163.367
R1224 B.n497 B.n70 163.367
R1225 B.n498 B.n497 163.367
R1226 B.n499 B.n498 163.367
R1227 B.n499 B.n68 163.367
R1228 B.n503 B.n68 163.367
R1229 B.n504 B.n503 163.367
R1230 B.n505 B.n504 163.367
R1231 B.n505 B.n66 163.367
R1232 B.n509 B.n66 163.367
R1233 B.n510 B.n509 163.367
R1234 B.n511 B.n510 163.367
R1235 B.n511 B.n64 163.367
R1236 B.n515 B.n64 163.367
R1237 B.n516 B.n515 163.367
R1238 B.n517 B.n516 163.367
R1239 B.n517 B.n62 163.367
R1240 B.n521 B.n62 163.367
R1241 B.n522 B.n521 163.367
R1242 B.n523 B.n522 163.367
R1243 B.n594 B.n33 163.367
R1244 B.n590 B.n33 163.367
R1245 B.n590 B.n589 163.367
R1246 B.n589 B.n588 163.367
R1247 B.n588 B.n35 163.367
R1248 B.n584 B.n35 163.367
R1249 B.n584 B.n583 163.367
R1250 B.n583 B.n582 163.367
R1251 B.n582 B.n37 163.367
R1252 B.n578 B.n37 163.367
R1253 B.n578 B.n577 163.367
R1254 B.n577 B.n576 163.367
R1255 B.n576 B.n39 163.367
R1256 B.n572 B.n39 163.367
R1257 B.n572 B.n571 163.367
R1258 B.n571 B.n570 163.367
R1259 B.n570 B.n41 163.367
R1260 B.n565 B.n41 163.367
R1261 B.n565 B.n564 163.367
R1262 B.n564 B.n563 163.367
R1263 B.n563 B.n45 163.367
R1264 B.n559 B.n45 163.367
R1265 B.n559 B.n558 163.367
R1266 B.n558 B.n557 163.367
R1267 B.n557 B.n47 163.367
R1268 B.n553 B.n47 163.367
R1269 B.n553 B.n552 163.367
R1270 B.n552 B.n551 163.367
R1271 B.n551 B.n49 163.367
R1272 B.n547 B.n49 163.367
R1273 B.n547 B.n546 163.367
R1274 B.n546 B.n545 163.367
R1275 B.n545 B.n54 163.367
R1276 B.n541 B.n54 163.367
R1277 B.n541 B.n540 163.367
R1278 B.n540 B.n539 163.367
R1279 B.n539 B.n56 163.367
R1280 B.n535 B.n56 163.367
R1281 B.n535 B.n534 163.367
R1282 B.n534 B.n533 163.367
R1283 B.n533 B.n58 163.367
R1284 B.n529 B.n58 163.367
R1285 B.n529 B.n528 163.367
R1286 B.n528 B.n527 163.367
R1287 B.n527 B.n60 163.367
R1288 B.n133 B.n132 59.5399
R1289 B.n297 B.n140 59.5399
R1290 B.n567 B.n43 59.5399
R1291 B.n52 B.n51 59.5399
R1292 B.n132 B.n131 58.3763
R1293 B.n140 B.n139 58.3763
R1294 B.n43 B.n42 58.3763
R1295 B.n51 B.n50 58.3763
R1296 B.n593 B.n32 32.6249
R1297 B.n525 B.n524 32.6249
R1298 B.n340 B.n339 32.6249
R1299 B.n268 B.n149 32.6249
R1300 B B.n687 18.0485
R1301 B.n593 B.n592 10.6151
R1302 B.n592 B.n591 10.6151
R1303 B.n591 B.n34 10.6151
R1304 B.n587 B.n34 10.6151
R1305 B.n587 B.n586 10.6151
R1306 B.n586 B.n585 10.6151
R1307 B.n585 B.n36 10.6151
R1308 B.n581 B.n36 10.6151
R1309 B.n581 B.n580 10.6151
R1310 B.n580 B.n579 10.6151
R1311 B.n579 B.n38 10.6151
R1312 B.n575 B.n38 10.6151
R1313 B.n575 B.n574 10.6151
R1314 B.n574 B.n573 10.6151
R1315 B.n573 B.n40 10.6151
R1316 B.n569 B.n40 10.6151
R1317 B.n569 B.n568 10.6151
R1318 B.n566 B.n44 10.6151
R1319 B.n562 B.n44 10.6151
R1320 B.n562 B.n561 10.6151
R1321 B.n561 B.n560 10.6151
R1322 B.n560 B.n46 10.6151
R1323 B.n556 B.n46 10.6151
R1324 B.n556 B.n555 10.6151
R1325 B.n555 B.n554 10.6151
R1326 B.n554 B.n48 10.6151
R1327 B.n550 B.n549 10.6151
R1328 B.n549 B.n548 10.6151
R1329 B.n548 B.n53 10.6151
R1330 B.n544 B.n53 10.6151
R1331 B.n544 B.n543 10.6151
R1332 B.n543 B.n542 10.6151
R1333 B.n542 B.n55 10.6151
R1334 B.n538 B.n55 10.6151
R1335 B.n538 B.n537 10.6151
R1336 B.n537 B.n536 10.6151
R1337 B.n536 B.n57 10.6151
R1338 B.n532 B.n57 10.6151
R1339 B.n532 B.n531 10.6151
R1340 B.n531 B.n530 10.6151
R1341 B.n530 B.n59 10.6151
R1342 B.n526 B.n59 10.6151
R1343 B.n526 B.n525 10.6151
R1344 B.n340 B.n121 10.6151
R1345 B.n344 B.n121 10.6151
R1346 B.n345 B.n344 10.6151
R1347 B.n346 B.n345 10.6151
R1348 B.n346 B.n119 10.6151
R1349 B.n350 B.n119 10.6151
R1350 B.n351 B.n350 10.6151
R1351 B.n352 B.n351 10.6151
R1352 B.n352 B.n117 10.6151
R1353 B.n356 B.n117 10.6151
R1354 B.n357 B.n356 10.6151
R1355 B.n358 B.n357 10.6151
R1356 B.n358 B.n115 10.6151
R1357 B.n362 B.n115 10.6151
R1358 B.n363 B.n362 10.6151
R1359 B.n364 B.n363 10.6151
R1360 B.n364 B.n113 10.6151
R1361 B.n368 B.n113 10.6151
R1362 B.n369 B.n368 10.6151
R1363 B.n370 B.n369 10.6151
R1364 B.n370 B.n111 10.6151
R1365 B.n374 B.n111 10.6151
R1366 B.n375 B.n374 10.6151
R1367 B.n376 B.n375 10.6151
R1368 B.n376 B.n109 10.6151
R1369 B.n380 B.n109 10.6151
R1370 B.n381 B.n380 10.6151
R1371 B.n382 B.n381 10.6151
R1372 B.n382 B.n107 10.6151
R1373 B.n386 B.n107 10.6151
R1374 B.n387 B.n386 10.6151
R1375 B.n388 B.n387 10.6151
R1376 B.n388 B.n105 10.6151
R1377 B.n392 B.n105 10.6151
R1378 B.n393 B.n392 10.6151
R1379 B.n394 B.n393 10.6151
R1380 B.n394 B.n103 10.6151
R1381 B.n398 B.n103 10.6151
R1382 B.n399 B.n398 10.6151
R1383 B.n400 B.n399 10.6151
R1384 B.n400 B.n101 10.6151
R1385 B.n404 B.n101 10.6151
R1386 B.n405 B.n404 10.6151
R1387 B.n406 B.n405 10.6151
R1388 B.n406 B.n99 10.6151
R1389 B.n410 B.n99 10.6151
R1390 B.n411 B.n410 10.6151
R1391 B.n412 B.n411 10.6151
R1392 B.n412 B.n97 10.6151
R1393 B.n416 B.n97 10.6151
R1394 B.n417 B.n416 10.6151
R1395 B.n418 B.n417 10.6151
R1396 B.n418 B.n95 10.6151
R1397 B.n422 B.n95 10.6151
R1398 B.n423 B.n422 10.6151
R1399 B.n424 B.n423 10.6151
R1400 B.n424 B.n93 10.6151
R1401 B.n428 B.n93 10.6151
R1402 B.n429 B.n428 10.6151
R1403 B.n430 B.n429 10.6151
R1404 B.n430 B.n91 10.6151
R1405 B.n434 B.n91 10.6151
R1406 B.n435 B.n434 10.6151
R1407 B.n436 B.n435 10.6151
R1408 B.n436 B.n89 10.6151
R1409 B.n440 B.n89 10.6151
R1410 B.n441 B.n440 10.6151
R1411 B.n442 B.n441 10.6151
R1412 B.n442 B.n87 10.6151
R1413 B.n446 B.n87 10.6151
R1414 B.n447 B.n446 10.6151
R1415 B.n448 B.n447 10.6151
R1416 B.n448 B.n85 10.6151
R1417 B.n452 B.n85 10.6151
R1418 B.n453 B.n452 10.6151
R1419 B.n454 B.n453 10.6151
R1420 B.n454 B.n83 10.6151
R1421 B.n458 B.n83 10.6151
R1422 B.n459 B.n458 10.6151
R1423 B.n460 B.n459 10.6151
R1424 B.n460 B.n81 10.6151
R1425 B.n464 B.n81 10.6151
R1426 B.n465 B.n464 10.6151
R1427 B.n466 B.n465 10.6151
R1428 B.n466 B.n79 10.6151
R1429 B.n470 B.n79 10.6151
R1430 B.n471 B.n470 10.6151
R1431 B.n472 B.n471 10.6151
R1432 B.n472 B.n77 10.6151
R1433 B.n476 B.n77 10.6151
R1434 B.n477 B.n476 10.6151
R1435 B.n478 B.n477 10.6151
R1436 B.n478 B.n75 10.6151
R1437 B.n482 B.n75 10.6151
R1438 B.n483 B.n482 10.6151
R1439 B.n484 B.n483 10.6151
R1440 B.n484 B.n73 10.6151
R1441 B.n488 B.n73 10.6151
R1442 B.n489 B.n488 10.6151
R1443 B.n490 B.n489 10.6151
R1444 B.n490 B.n71 10.6151
R1445 B.n494 B.n71 10.6151
R1446 B.n495 B.n494 10.6151
R1447 B.n496 B.n495 10.6151
R1448 B.n496 B.n69 10.6151
R1449 B.n500 B.n69 10.6151
R1450 B.n501 B.n500 10.6151
R1451 B.n502 B.n501 10.6151
R1452 B.n502 B.n67 10.6151
R1453 B.n506 B.n67 10.6151
R1454 B.n507 B.n506 10.6151
R1455 B.n508 B.n507 10.6151
R1456 B.n508 B.n65 10.6151
R1457 B.n512 B.n65 10.6151
R1458 B.n513 B.n512 10.6151
R1459 B.n514 B.n513 10.6151
R1460 B.n514 B.n63 10.6151
R1461 B.n518 B.n63 10.6151
R1462 B.n519 B.n518 10.6151
R1463 B.n520 B.n519 10.6151
R1464 B.n520 B.n61 10.6151
R1465 B.n524 B.n61 10.6151
R1466 B.n272 B.n149 10.6151
R1467 B.n273 B.n272 10.6151
R1468 B.n274 B.n273 10.6151
R1469 B.n274 B.n147 10.6151
R1470 B.n278 B.n147 10.6151
R1471 B.n279 B.n278 10.6151
R1472 B.n280 B.n279 10.6151
R1473 B.n280 B.n145 10.6151
R1474 B.n284 B.n145 10.6151
R1475 B.n285 B.n284 10.6151
R1476 B.n286 B.n285 10.6151
R1477 B.n286 B.n143 10.6151
R1478 B.n290 B.n143 10.6151
R1479 B.n291 B.n290 10.6151
R1480 B.n292 B.n291 10.6151
R1481 B.n292 B.n141 10.6151
R1482 B.n296 B.n141 10.6151
R1483 B.n299 B.n298 10.6151
R1484 B.n299 B.n137 10.6151
R1485 B.n303 B.n137 10.6151
R1486 B.n304 B.n303 10.6151
R1487 B.n305 B.n304 10.6151
R1488 B.n305 B.n135 10.6151
R1489 B.n309 B.n135 10.6151
R1490 B.n310 B.n309 10.6151
R1491 B.n311 B.n310 10.6151
R1492 B.n315 B.n314 10.6151
R1493 B.n316 B.n315 10.6151
R1494 B.n316 B.n129 10.6151
R1495 B.n320 B.n129 10.6151
R1496 B.n321 B.n320 10.6151
R1497 B.n322 B.n321 10.6151
R1498 B.n322 B.n127 10.6151
R1499 B.n326 B.n127 10.6151
R1500 B.n327 B.n326 10.6151
R1501 B.n328 B.n327 10.6151
R1502 B.n328 B.n125 10.6151
R1503 B.n332 B.n125 10.6151
R1504 B.n333 B.n332 10.6151
R1505 B.n334 B.n333 10.6151
R1506 B.n334 B.n123 10.6151
R1507 B.n338 B.n123 10.6151
R1508 B.n339 B.n338 10.6151
R1509 B.n268 B.n267 10.6151
R1510 B.n267 B.n266 10.6151
R1511 B.n266 B.n151 10.6151
R1512 B.n262 B.n151 10.6151
R1513 B.n262 B.n261 10.6151
R1514 B.n261 B.n260 10.6151
R1515 B.n260 B.n153 10.6151
R1516 B.n256 B.n153 10.6151
R1517 B.n256 B.n255 10.6151
R1518 B.n255 B.n254 10.6151
R1519 B.n254 B.n155 10.6151
R1520 B.n250 B.n155 10.6151
R1521 B.n250 B.n249 10.6151
R1522 B.n249 B.n248 10.6151
R1523 B.n248 B.n157 10.6151
R1524 B.n244 B.n157 10.6151
R1525 B.n244 B.n243 10.6151
R1526 B.n243 B.n242 10.6151
R1527 B.n242 B.n159 10.6151
R1528 B.n238 B.n159 10.6151
R1529 B.n238 B.n237 10.6151
R1530 B.n237 B.n236 10.6151
R1531 B.n236 B.n161 10.6151
R1532 B.n232 B.n161 10.6151
R1533 B.n232 B.n231 10.6151
R1534 B.n231 B.n230 10.6151
R1535 B.n230 B.n163 10.6151
R1536 B.n226 B.n163 10.6151
R1537 B.n226 B.n225 10.6151
R1538 B.n225 B.n224 10.6151
R1539 B.n224 B.n165 10.6151
R1540 B.n220 B.n165 10.6151
R1541 B.n220 B.n219 10.6151
R1542 B.n219 B.n218 10.6151
R1543 B.n218 B.n167 10.6151
R1544 B.n214 B.n167 10.6151
R1545 B.n214 B.n213 10.6151
R1546 B.n213 B.n212 10.6151
R1547 B.n212 B.n169 10.6151
R1548 B.n208 B.n169 10.6151
R1549 B.n208 B.n207 10.6151
R1550 B.n207 B.n206 10.6151
R1551 B.n206 B.n171 10.6151
R1552 B.n202 B.n171 10.6151
R1553 B.n202 B.n201 10.6151
R1554 B.n201 B.n200 10.6151
R1555 B.n200 B.n173 10.6151
R1556 B.n196 B.n173 10.6151
R1557 B.n196 B.n195 10.6151
R1558 B.n195 B.n194 10.6151
R1559 B.n194 B.n175 10.6151
R1560 B.n190 B.n175 10.6151
R1561 B.n190 B.n189 10.6151
R1562 B.n189 B.n188 10.6151
R1563 B.n188 B.n177 10.6151
R1564 B.n184 B.n177 10.6151
R1565 B.n184 B.n183 10.6151
R1566 B.n183 B.n182 10.6151
R1567 B.n182 B.n179 10.6151
R1568 B.n179 B.n0 10.6151
R1569 B.n683 B.n1 10.6151
R1570 B.n683 B.n682 10.6151
R1571 B.n682 B.n681 10.6151
R1572 B.n681 B.n4 10.6151
R1573 B.n677 B.n4 10.6151
R1574 B.n677 B.n676 10.6151
R1575 B.n676 B.n675 10.6151
R1576 B.n675 B.n6 10.6151
R1577 B.n671 B.n6 10.6151
R1578 B.n671 B.n670 10.6151
R1579 B.n670 B.n669 10.6151
R1580 B.n669 B.n8 10.6151
R1581 B.n665 B.n8 10.6151
R1582 B.n665 B.n664 10.6151
R1583 B.n664 B.n663 10.6151
R1584 B.n663 B.n10 10.6151
R1585 B.n659 B.n10 10.6151
R1586 B.n659 B.n658 10.6151
R1587 B.n658 B.n657 10.6151
R1588 B.n657 B.n12 10.6151
R1589 B.n653 B.n12 10.6151
R1590 B.n653 B.n652 10.6151
R1591 B.n652 B.n651 10.6151
R1592 B.n651 B.n14 10.6151
R1593 B.n647 B.n14 10.6151
R1594 B.n647 B.n646 10.6151
R1595 B.n646 B.n645 10.6151
R1596 B.n645 B.n16 10.6151
R1597 B.n641 B.n16 10.6151
R1598 B.n641 B.n640 10.6151
R1599 B.n640 B.n639 10.6151
R1600 B.n639 B.n18 10.6151
R1601 B.n635 B.n18 10.6151
R1602 B.n635 B.n634 10.6151
R1603 B.n634 B.n633 10.6151
R1604 B.n633 B.n20 10.6151
R1605 B.n629 B.n20 10.6151
R1606 B.n629 B.n628 10.6151
R1607 B.n628 B.n627 10.6151
R1608 B.n627 B.n22 10.6151
R1609 B.n623 B.n22 10.6151
R1610 B.n623 B.n622 10.6151
R1611 B.n622 B.n621 10.6151
R1612 B.n621 B.n24 10.6151
R1613 B.n617 B.n24 10.6151
R1614 B.n617 B.n616 10.6151
R1615 B.n616 B.n615 10.6151
R1616 B.n615 B.n26 10.6151
R1617 B.n611 B.n26 10.6151
R1618 B.n611 B.n610 10.6151
R1619 B.n610 B.n609 10.6151
R1620 B.n609 B.n28 10.6151
R1621 B.n605 B.n28 10.6151
R1622 B.n605 B.n604 10.6151
R1623 B.n604 B.n603 10.6151
R1624 B.n603 B.n30 10.6151
R1625 B.n599 B.n30 10.6151
R1626 B.n599 B.n598 10.6151
R1627 B.n598 B.n597 10.6151
R1628 B.n597 B.n32 10.6151
R1629 B.n568 B.n567 9.52245
R1630 B.n550 B.n52 9.52245
R1631 B.n297 B.n296 9.52245
R1632 B.n314 B.n133 9.52245
R1633 B.n687 B.n0 2.81026
R1634 B.n687 B.n1 2.81026
R1635 B.n567 B.n566 1.09318
R1636 B.n52 B.n48 1.09318
R1637 B.n298 B.n297 1.09318
R1638 B.n311 B.n133 1.09318
C0 B VN 1.24944f
C1 VDD2 VN 3.91286f
C2 VDD2 B 1.99685f
C3 VDD1 w_n4582_n1762# 2.25245f
C4 VDD1 VP 4.34983f
C5 VDD1 VTAIL 6.76217f
C6 w_n4582_n1762# VP 10.3211f
C7 w_n4582_n1762# VTAIL 2.0618f
C8 VP VTAIL 5.21277f
C9 VDD1 VN 0.157504f
C10 B VDD1 1.87566f
C11 w_n4582_n1762# VN 9.72518f
C12 B w_n4582_n1762# 8.46734f
C13 VDD2 VDD1 2.22273f
C14 VP VN 7.03885f
C15 VTAIL VN 5.19861f
C16 B VP 2.25323f
C17 VDD2 w_n4582_n1762# 2.39979f
C18 B VTAIL 1.91957f
C19 VDD2 VP 0.597792f
C20 VDD2 VTAIL 6.81555f
C21 VDD2 VSUBS 1.924528f
C22 VDD1 VSUBS 1.774029f
C23 VTAIL VSUBS 0.61665f
C24 VN VSUBS 7.57042f
C25 VP VSUBS 3.718457f
C26 B VSUBS 4.503272f
C27 w_n4582_n1762# VSUBS 0.101665p
C28 B.n0 VSUBS 0.005593f
C29 B.n1 VSUBS 0.005593f
C30 B.n2 VSUBS 0.008845f
C31 B.n3 VSUBS 0.008845f
C32 B.n4 VSUBS 0.008845f
C33 B.n5 VSUBS 0.008845f
C34 B.n6 VSUBS 0.008845f
C35 B.n7 VSUBS 0.008845f
C36 B.n8 VSUBS 0.008845f
C37 B.n9 VSUBS 0.008845f
C38 B.n10 VSUBS 0.008845f
C39 B.n11 VSUBS 0.008845f
C40 B.n12 VSUBS 0.008845f
C41 B.n13 VSUBS 0.008845f
C42 B.n14 VSUBS 0.008845f
C43 B.n15 VSUBS 0.008845f
C44 B.n16 VSUBS 0.008845f
C45 B.n17 VSUBS 0.008845f
C46 B.n18 VSUBS 0.008845f
C47 B.n19 VSUBS 0.008845f
C48 B.n20 VSUBS 0.008845f
C49 B.n21 VSUBS 0.008845f
C50 B.n22 VSUBS 0.008845f
C51 B.n23 VSUBS 0.008845f
C52 B.n24 VSUBS 0.008845f
C53 B.n25 VSUBS 0.008845f
C54 B.n26 VSUBS 0.008845f
C55 B.n27 VSUBS 0.008845f
C56 B.n28 VSUBS 0.008845f
C57 B.n29 VSUBS 0.008845f
C58 B.n30 VSUBS 0.008845f
C59 B.n31 VSUBS 0.008845f
C60 B.n32 VSUBS 0.0198f
C61 B.n33 VSUBS 0.008845f
C62 B.n34 VSUBS 0.008845f
C63 B.n35 VSUBS 0.008845f
C64 B.n36 VSUBS 0.008845f
C65 B.n37 VSUBS 0.008845f
C66 B.n38 VSUBS 0.008845f
C67 B.n39 VSUBS 0.008845f
C68 B.n40 VSUBS 0.008845f
C69 B.n41 VSUBS 0.008845f
C70 B.t8 VSUBS 0.072823f
C71 B.t7 VSUBS 0.099282f
C72 B.t6 VSUBS 0.647632f
C73 B.n42 VSUBS 0.172462f
C74 B.n43 VSUBS 0.145698f
C75 B.n44 VSUBS 0.008845f
C76 B.n45 VSUBS 0.008845f
C77 B.n46 VSUBS 0.008845f
C78 B.n47 VSUBS 0.008845f
C79 B.n48 VSUBS 0.004877f
C80 B.n49 VSUBS 0.008845f
C81 B.t2 VSUBS 0.072824f
C82 B.t1 VSUBS 0.099283f
C83 B.t0 VSUBS 0.64768f
C84 B.n50 VSUBS 0.172414f
C85 B.n51 VSUBS 0.145697f
C86 B.n52 VSUBS 0.020492f
C87 B.n53 VSUBS 0.008845f
C88 B.n54 VSUBS 0.008845f
C89 B.n55 VSUBS 0.008845f
C90 B.n56 VSUBS 0.008845f
C91 B.n57 VSUBS 0.008845f
C92 B.n58 VSUBS 0.008845f
C93 B.n59 VSUBS 0.008845f
C94 B.n60 VSUBS 0.021561f
C95 B.n61 VSUBS 0.008845f
C96 B.n62 VSUBS 0.008845f
C97 B.n63 VSUBS 0.008845f
C98 B.n64 VSUBS 0.008845f
C99 B.n65 VSUBS 0.008845f
C100 B.n66 VSUBS 0.008845f
C101 B.n67 VSUBS 0.008845f
C102 B.n68 VSUBS 0.008845f
C103 B.n69 VSUBS 0.008845f
C104 B.n70 VSUBS 0.008845f
C105 B.n71 VSUBS 0.008845f
C106 B.n72 VSUBS 0.008845f
C107 B.n73 VSUBS 0.008845f
C108 B.n74 VSUBS 0.008845f
C109 B.n75 VSUBS 0.008845f
C110 B.n76 VSUBS 0.008845f
C111 B.n77 VSUBS 0.008845f
C112 B.n78 VSUBS 0.008845f
C113 B.n79 VSUBS 0.008845f
C114 B.n80 VSUBS 0.008845f
C115 B.n81 VSUBS 0.008845f
C116 B.n82 VSUBS 0.008845f
C117 B.n83 VSUBS 0.008845f
C118 B.n84 VSUBS 0.008845f
C119 B.n85 VSUBS 0.008845f
C120 B.n86 VSUBS 0.008845f
C121 B.n87 VSUBS 0.008845f
C122 B.n88 VSUBS 0.008845f
C123 B.n89 VSUBS 0.008845f
C124 B.n90 VSUBS 0.008845f
C125 B.n91 VSUBS 0.008845f
C126 B.n92 VSUBS 0.008845f
C127 B.n93 VSUBS 0.008845f
C128 B.n94 VSUBS 0.008845f
C129 B.n95 VSUBS 0.008845f
C130 B.n96 VSUBS 0.008845f
C131 B.n97 VSUBS 0.008845f
C132 B.n98 VSUBS 0.008845f
C133 B.n99 VSUBS 0.008845f
C134 B.n100 VSUBS 0.008845f
C135 B.n101 VSUBS 0.008845f
C136 B.n102 VSUBS 0.008845f
C137 B.n103 VSUBS 0.008845f
C138 B.n104 VSUBS 0.008845f
C139 B.n105 VSUBS 0.008845f
C140 B.n106 VSUBS 0.008845f
C141 B.n107 VSUBS 0.008845f
C142 B.n108 VSUBS 0.008845f
C143 B.n109 VSUBS 0.008845f
C144 B.n110 VSUBS 0.008845f
C145 B.n111 VSUBS 0.008845f
C146 B.n112 VSUBS 0.008845f
C147 B.n113 VSUBS 0.008845f
C148 B.n114 VSUBS 0.008845f
C149 B.n115 VSUBS 0.008845f
C150 B.n116 VSUBS 0.008845f
C151 B.n117 VSUBS 0.008845f
C152 B.n118 VSUBS 0.008845f
C153 B.n119 VSUBS 0.008845f
C154 B.n120 VSUBS 0.008845f
C155 B.n121 VSUBS 0.008845f
C156 B.n122 VSUBS 0.021561f
C157 B.n123 VSUBS 0.008845f
C158 B.n124 VSUBS 0.008845f
C159 B.n125 VSUBS 0.008845f
C160 B.n126 VSUBS 0.008845f
C161 B.n127 VSUBS 0.008845f
C162 B.n128 VSUBS 0.008845f
C163 B.n129 VSUBS 0.008845f
C164 B.n130 VSUBS 0.008845f
C165 B.t10 VSUBS 0.072824f
C166 B.t11 VSUBS 0.099283f
C167 B.t9 VSUBS 0.64768f
C168 B.n131 VSUBS 0.172414f
C169 B.n132 VSUBS 0.145697f
C170 B.n133 VSUBS 0.020492f
C171 B.n134 VSUBS 0.008845f
C172 B.n135 VSUBS 0.008845f
C173 B.n136 VSUBS 0.008845f
C174 B.n137 VSUBS 0.008845f
C175 B.n138 VSUBS 0.008845f
C176 B.t4 VSUBS 0.072823f
C177 B.t5 VSUBS 0.099282f
C178 B.t3 VSUBS 0.647632f
C179 B.n139 VSUBS 0.172462f
C180 B.n140 VSUBS 0.145698f
C181 B.n141 VSUBS 0.008845f
C182 B.n142 VSUBS 0.008845f
C183 B.n143 VSUBS 0.008845f
C184 B.n144 VSUBS 0.008845f
C185 B.n145 VSUBS 0.008845f
C186 B.n146 VSUBS 0.008845f
C187 B.n147 VSUBS 0.008845f
C188 B.n148 VSUBS 0.008845f
C189 B.n149 VSUBS 0.021561f
C190 B.n150 VSUBS 0.008845f
C191 B.n151 VSUBS 0.008845f
C192 B.n152 VSUBS 0.008845f
C193 B.n153 VSUBS 0.008845f
C194 B.n154 VSUBS 0.008845f
C195 B.n155 VSUBS 0.008845f
C196 B.n156 VSUBS 0.008845f
C197 B.n157 VSUBS 0.008845f
C198 B.n158 VSUBS 0.008845f
C199 B.n159 VSUBS 0.008845f
C200 B.n160 VSUBS 0.008845f
C201 B.n161 VSUBS 0.008845f
C202 B.n162 VSUBS 0.008845f
C203 B.n163 VSUBS 0.008845f
C204 B.n164 VSUBS 0.008845f
C205 B.n165 VSUBS 0.008845f
C206 B.n166 VSUBS 0.008845f
C207 B.n167 VSUBS 0.008845f
C208 B.n168 VSUBS 0.008845f
C209 B.n169 VSUBS 0.008845f
C210 B.n170 VSUBS 0.008845f
C211 B.n171 VSUBS 0.008845f
C212 B.n172 VSUBS 0.008845f
C213 B.n173 VSUBS 0.008845f
C214 B.n174 VSUBS 0.008845f
C215 B.n175 VSUBS 0.008845f
C216 B.n176 VSUBS 0.008845f
C217 B.n177 VSUBS 0.008845f
C218 B.n178 VSUBS 0.008845f
C219 B.n179 VSUBS 0.008845f
C220 B.n180 VSUBS 0.008845f
C221 B.n181 VSUBS 0.008845f
C222 B.n182 VSUBS 0.008845f
C223 B.n183 VSUBS 0.008845f
C224 B.n184 VSUBS 0.008845f
C225 B.n185 VSUBS 0.008845f
C226 B.n186 VSUBS 0.008845f
C227 B.n187 VSUBS 0.008845f
C228 B.n188 VSUBS 0.008845f
C229 B.n189 VSUBS 0.008845f
C230 B.n190 VSUBS 0.008845f
C231 B.n191 VSUBS 0.008845f
C232 B.n192 VSUBS 0.008845f
C233 B.n193 VSUBS 0.008845f
C234 B.n194 VSUBS 0.008845f
C235 B.n195 VSUBS 0.008845f
C236 B.n196 VSUBS 0.008845f
C237 B.n197 VSUBS 0.008845f
C238 B.n198 VSUBS 0.008845f
C239 B.n199 VSUBS 0.008845f
C240 B.n200 VSUBS 0.008845f
C241 B.n201 VSUBS 0.008845f
C242 B.n202 VSUBS 0.008845f
C243 B.n203 VSUBS 0.008845f
C244 B.n204 VSUBS 0.008845f
C245 B.n205 VSUBS 0.008845f
C246 B.n206 VSUBS 0.008845f
C247 B.n207 VSUBS 0.008845f
C248 B.n208 VSUBS 0.008845f
C249 B.n209 VSUBS 0.008845f
C250 B.n210 VSUBS 0.008845f
C251 B.n211 VSUBS 0.008845f
C252 B.n212 VSUBS 0.008845f
C253 B.n213 VSUBS 0.008845f
C254 B.n214 VSUBS 0.008845f
C255 B.n215 VSUBS 0.008845f
C256 B.n216 VSUBS 0.008845f
C257 B.n217 VSUBS 0.008845f
C258 B.n218 VSUBS 0.008845f
C259 B.n219 VSUBS 0.008845f
C260 B.n220 VSUBS 0.008845f
C261 B.n221 VSUBS 0.008845f
C262 B.n222 VSUBS 0.008845f
C263 B.n223 VSUBS 0.008845f
C264 B.n224 VSUBS 0.008845f
C265 B.n225 VSUBS 0.008845f
C266 B.n226 VSUBS 0.008845f
C267 B.n227 VSUBS 0.008845f
C268 B.n228 VSUBS 0.008845f
C269 B.n229 VSUBS 0.008845f
C270 B.n230 VSUBS 0.008845f
C271 B.n231 VSUBS 0.008845f
C272 B.n232 VSUBS 0.008845f
C273 B.n233 VSUBS 0.008845f
C274 B.n234 VSUBS 0.008845f
C275 B.n235 VSUBS 0.008845f
C276 B.n236 VSUBS 0.008845f
C277 B.n237 VSUBS 0.008845f
C278 B.n238 VSUBS 0.008845f
C279 B.n239 VSUBS 0.008845f
C280 B.n240 VSUBS 0.008845f
C281 B.n241 VSUBS 0.008845f
C282 B.n242 VSUBS 0.008845f
C283 B.n243 VSUBS 0.008845f
C284 B.n244 VSUBS 0.008845f
C285 B.n245 VSUBS 0.008845f
C286 B.n246 VSUBS 0.008845f
C287 B.n247 VSUBS 0.008845f
C288 B.n248 VSUBS 0.008845f
C289 B.n249 VSUBS 0.008845f
C290 B.n250 VSUBS 0.008845f
C291 B.n251 VSUBS 0.008845f
C292 B.n252 VSUBS 0.008845f
C293 B.n253 VSUBS 0.008845f
C294 B.n254 VSUBS 0.008845f
C295 B.n255 VSUBS 0.008845f
C296 B.n256 VSUBS 0.008845f
C297 B.n257 VSUBS 0.008845f
C298 B.n258 VSUBS 0.008845f
C299 B.n259 VSUBS 0.008845f
C300 B.n260 VSUBS 0.008845f
C301 B.n261 VSUBS 0.008845f
C302 B.n262 VSUBS 0.008845f
C303 B.n263 VSUBS 0.008845f
C304 B.n264 VSUBS 0.008845f
C305 B.n265 VSUBS 0.008845f
C306 B.n266 VSUBS 0.008845f
C307 B.n267 VSUBS 0.008845f
C308 B.n268 VSUBS 0.0198f
C309 B.n269 VSUBS 0.0198f
C310 B.n270 VSUBS 0.021561f
C311 B.n271 VSUBS 0.008845f
C312 B.n272 VSUBS 0.008845f
C313 B.n273 VSUBS 0.008845f
C314 B.n274 VSUBS 0.008845f
C315 B.n275 VSUBS 0.008845f
C316 B.n276 VSUBS 0.008845f
C317 B.n277 VSUBS 0.008845f
C318 B.n278 VSUBS 0.008845f
C319 B.n279 VSUBS 0.008845f
C320 B.n280 VSUBS 0.008845f
C321 B.n281 VSUBS 0.008845f
C322 B.n282 VSUBS 0.008845f
C323 B.n283 VSUBS 0.008845f
C324 B.n284 VSUBS 0.008845f
C325 B.n285 VSUBS 0.008845f
C326 B.n286 VSUBS 0.008845f
C327 B.n287 VSUBS 0.008845f
C328 B.n288 VSUBS 0.008845f
C329 B.n289 VSUBS 0.008845f
C330 B.n290 VSUBS 0.008845f
C331 B.n291 VSUBS 0.008845f
C332 B.n292 VSUBS 0.008845f
C333 B.n293 VSUBS 0.008845f
C334 B.n294 VSUBS 0.008845f
C335 B.n295 VSUBS 0.008845f
C336 B.n296 VSUBS 0.008389f
C337 B.n297 VSUBS 0.020492f
C338 B.n298 VSUBS 0.004877f
C339 B.n299 VSUBS 0.008845f
C340 B.n300 VSUBS 0.008845f
C341 B.n301 VSUBS 0.008845f
C342 B.n302 VSUBS 0.008845f
C343 B.n303 VSUBS 0.008845f
C344 B.n304 VSUBS 0.008845f
C345 B.n305 VSUBS 0.008845f
C346 B.n306 VSUBS 0.008845f
C347 B.n307 VSUBS 0.008845f
C348 B.n308 VSUBS 0.008845f
C349 B.n309 VSUBS 0.008845f
C350 B.n310 VSUBS 0.008845f
C351 B.n311 VSUBS 0.004877f
C352 B.n312 VSUBS 0.008845f
C353 B.n313 VSUBS 0.008845f
C354 B.n314 VSUBS 0.008389f
C355 B.n315 VSUBS 0.008845f
C356 B.n316 VSUBS 0.008845f
C357 B.n317 VSUBS 0.008845f
C358 B.n318 VSUBS 0.008845f
C359 B.n319 VSUBS 0.008845f
C360 B.n320 VSUBS 0.008845f
C361 B.n321 VSUBS 0.008845f
C362 B.n322 VSUBS 0.008845f
C363 B.n323 VSUBS 0.008845f
C364 B.n324 VSUBS 0.008845f
C365 B.n325 VSUBS 0.008845f
C366 B.n326 VSUBS 0.008845f
C367 B.n327 VSUBS 0.008845f
C368 B.n328 VSUBS 0.008845f
C369 B.n329 VSUBS 0.008845f
C370 B.n330 VSUBS 0.008845f
C371 B.n331 VSUBS 0.008845f
C372 B.n332 VSUBS 0.008845f
C373 B.n333 VSUBS 0.008845f
C374 B.n334 VSUBS 0.008845f
C375 B.n335 VSUBS 0.008845f
C376 B.n336 VSUBS 0.008845f
C377 B.n337 VSUBS 0.008845f
C378 B.n338 VSUBS 0.008845f
C379 B.n339 VSUBS 0.021561f
C380 B.n340 VSUBS 0.0198f
C381 B.n341 VSUBS 0.0198f
C382 B.n342 VSUBS 0.008845f
C383 B.n343 VSUBS 0.008845f
C384 B.n344 VSUBS 0.008845f
C385 B.n345 VSUBS 0.008845f
C386 B.n346 VSUBS 0.008845f
C387 B.n347 VSUBS 0.008845f
C388 B.n348 VSUBS 0.008845f
C389 B.n349 VSUBS 0.008845f
C390 B.n350 VSUBS 0.008845f
C391 B.n351 VSUBS 0.008845f
C392 B.n352 VSUBS 0.008845f
C393 B.n353 VSUBS 0.008845f
C394 B.n354 VSUBS 0.008845f
C395 B.n355 VSUBS 0.008845f
C396 B.n356 VSUBS 0.008845f
C397 B.n357 VSUBS 0.008845f
C398 B.n358 VSUBS 0.008845f
C399 B.n359 VSUBS 0.008845f
C400 B.n360 VSUBS 0.008845f
C401 B.n361 VSUBS 0.008845f
C402 B.n362 VSUBS 0.008845f
C403 B.n363 VSUBS 0.008845f
C404 B.n364 VSUBS 0.008845f
C405 B.n365 VSUBS 0.008845f
C406 B.n366 VSUBS 0.008845f
C407 B.n367 VSUBS 0.008845f
C408 B.n368 VSUBS 0.008845f
C409 B.n369 VSUBS 0.008845f
C410 B.n370 VSUBS 0.008845f
C411 B.n371 VSUBS 0.008845f
C412 B.n372 VSUBS 0.008845f
C413 B.n373 VSUBS 0.008845f
C414 B.n374 VSUBS 0.008845f
C415 B.n375 VSUBS 0.008845f
C416 B.n376 VSUBS 0.008845f
C417 B.n377 VSUBS 0.008845f
C418 B.n378 VSUBS 0.008845f
C419 B.n379 VSUBS 0.008845f
C420 B.n380 VSUBS 0.008845f
C421 B.n381 VSUBS 0.008845f
C422 B.n382 VSUBS 0.008845f
C423 B.n383 VSUBS 0.008845f
C424 B.n384 VSUBS 0.008845f
C425 B.n385 VSUBS 0.008845f
C426 B.n386 VSUBS 0.008845f
C427 B.n387 VSUBS 0.008845f
C428 B.n388 VSUBS 0.008845f
C429 B.n389 VSUBS 0.008845f
C430 B.n390 VSUBS 0.008845f
C431 B.n391 VSUBS 0.008845f
C432 B.n392 VSUBS 0.008845f
C433 B.n393 VSUBS 0.008845f
C434 B.n394 VSUBS 0.008845f
C435 B.n395 VSUBS 0.008845f
C436 B.n396 VSUBS 0.008845f
C437 B.n397 VSUBS 0.008845f
C438 B.n398 VSUBS 0.008845f
C439 B.n399 VSUBS 0.008845f
C440 B.n400 VSUBS 0.008845f
C441 B.n401 VSUBS 0.008845f
C442 B.n402 VSUBS 0.008845f
C443 B.n403 VSUBS 0.008845f
C444 B.n404 VSUBS 0.008845f
C445 B.n405 VSUBS 0.008845f
C446 B.n406 VSUBS 0.008845f
C447 B.n407 VSUBS 0.008845f
C448 B.n408 VSUBS 0.008845f
C449 B.n409 VSUBS 0.008845f
C450 B.n410 VSUBS 0.008845f
C451 B.n411 VSUBS 0.008845f
C452 B.n412 VSUBS 0.008845f
C453 B.n413 VSUBS 0.008845f
C454 B.n414 VSUBS 0.008845f
C455 B.n415 VSUBS 0.008845f
C456 B.n416 VSUBS 0.008845f
C457 B.n417 VSUBS 0.008845f
C458 B.n418 VSUBS 0.008845f
C459 B.n419 VSUBS 0.008845f
C460 B.n420 VSUBS 0.008845f
C461 B.n421 VSUBS 0.008845f
C462 B.n422 VSUBS 0.008845f
C463 B.n423 VSUBS 0.008845f
C464 B.n424 VSUBS 0.008845f
C465 B.n425 VSUBS 0.008845f
C466 B.n426 VSUBS 0.008845f
C467 B.n427 VSUBS 0.008845f
C468 B.n428 VSUBS 0.008845f
C469 B.n429 VSUBS 0.008845f
C470 B.n430 VSUBS 0.008845f
C471 B.n431 VSUBS 0.008845f
C472 B.n432 VSUBS 0.008845f
C473 B.n433 VSUBS 0.008845f
C474 B.n434 VSUBS 0.008845f
C475 B.n435 VSUBS 0.008845f
C476 B.n436 VSUBS 0.008845f
C477 B.n437 VSUBS 0.008845f
C478 B.n438 VSUBS 0.008845f
C479 B.n439 VSUBS 0.008845f
C480 B.n440 VSUBS 0.008845f
C481 B.n441 VSUBS 0.008845f
C482 B.n442 VSUBS 0.008845f
C483 B.n443 VSUBS 0.008845f
C484 B.n444 VSUBS 0.008845f
C485 B.n445 VSUBS 0.008845f
C486 B.n446 VSUBS 0.008845f
C487 B.n447 VSUBS 0.008845f
C488 B.n448 VSUBS 0.008845f
C489 B.n449 VSUBS 0.008845f
C490 B.n450 VSUBS 0.008845f
C491 B.n451 VSUBS 0.008845f
C492 B.n452 VSUBS 0.008845f
C493 B.n453 VSUBS 0.008845f
C494 B.n454 VSUBS 0.008845f
C495 B.n455 VSUBS 0.008845f
C496 B.n456 VSUBS 0.008845f
C497 B.n457 VSUBS 0.008845f
C498 B.n458 VSUBS 0.008845f
C499 B.n459 VSUBS 0.008845f
C500 B.n460 VSUBS 0.008845f
C501 B.n461 VSUBS 0.008845f
C502 B.n462 VSUBS 0.008845f
C503 B.n463 VSUBS 0.008845f
C504 B.n464 VSUBS 0.008845f
C505 B.n465 VSUBS 0.008845f
C506 B.n466 VSUBS 0.008845f
C507 B.n467 VSUBS 0.008845f
C508 B.n468 VSUBS 0.008845f
C509 B.n469 VSUBS 0.008845f
C510 B.n470 VSUBS 0.008845f
C511 B.n471 VSUBS 0.008845f
C512 B.n472 VSUBS 0.008845f
C513 B.n473 VSUBS 0.008845f
C514 B.n474 VSUBS 0.008845f
C515 B.n475 VSUBS 0.008845f
C516 B.n476 VSUBS 0.008845f
C517 B.n477 VSUBS 0.008845f
C518 B.n478 VSUBS 0.008845f
C519 B.n479 VSUBS 0.008845f
C520 B.n480 VSUBS 0.008845f
C521 B.n481 VSUBS 0.008845f
C522 B.n482 VSUBS 0.008845f
C523 B.n483 VSUBS 0.008845f
C524 B.n484 VSUBS 0.008845f
C525 B.n485 VSUBS 0.008845f
C526 B.n486 VSUBS 0.008845f
C527 B.n487 VSUBS 0.008845f
C528 B.n488 VSUBS 0.008845f
C529 B.n489 VSUBS 0.008845f
C530 B.n490 VSUBS 0.008845f
C531 B.n491 VSUBS 0.008845f
C532 B.n492 VSUBS 0.008845f
C533 B.n493 VSUBS 0.008845f
C534 B.n494 VSUBS 0.008845f
C535 B.n495 VSUBS 0.008845f
C536 B.n496 VSUBS 0.008845f
C537 B.n497 VSUBS 0.008845f
C538 B.n498 VSUBS 0.008845f
C539 B.n499 VSUBS 0.008845f
C540 B.n500 VSUBS 0.008845f
C541 B.n501 VSUBS 0.008845f
C542 B.n502 VSUBS 0.008845f
C543 B.n503 VSUBS 0.008845f
C544 B.n504 VSUBS 0.008845f
C545 B.n505 VSUBS 0.008845f
C546 B.n506 VSUBS 0.008845f
C547 B.n507 VSUBS 0.008845f
C548 B.n508 VSUBS 0.008845f
C549 B.n509 VSUBS 0.008845f
C550 B.n510 VSUBS 0.008845f
C551 B.n511 VSUBS 0.008845f
C552 B.n512 VSUBS 0.008845f
C553 B.n513 VSUBS 0.008845f
C554 B.n514 VSUBS 0.008845f
C555 B.n515 VSUBS 0.008845f
C556 B.n516 VSUBS 0.008845f
C557 B.n517 VSUBS 0.008845f
C558 B.n518 VSUBS 0.008845f
C559 B.n519 VSUBS 0.008845f
C560 B.n520 VSUBS 0.008845f
C561 B.n521 VSUBS 0.008845f
C562 B.n522 VSUBS 0.008845f
C563 B.n523 VSUBS 0.0198f
C564 B.n524 VSUBS 0.020846f
C565 B.n525 VSUBS 0.020515f
C566 B.n526 VSUBS 0.008845f
C567 B.n527 VSUBS 0.008845f
C568 B.n528 VSUBS 0.008845f
C569 B.n529 VSUBS 0.008845f
C570 B.n530 VSUBS 0.008845f
C571 B.n531 VSUBS 0.008845f
C572 B.n532 VSUBS 0.008845f
C573 B.n533 VSUBS 0.008845f
C574 B.n534 VSUBS 0.008845f
C575 B.n535 VSUBS 0.008845f
C576 B.n536 VSUBS 0.008845f
C577 B.n537 VSUBS 0.008845f
C578 B.n538 VSUBS 0.008845f
C579 B.n539 VSUBS 0.008845f
C580 B.n540 VSUBS 0.008845f
C581 B.n541 VSUBS 0.008845f
C582 B.n542 VSUBS 0.008845f
C583 B.n543 VSUBS 0.008845f
C584 B.n544 VSUBS 0.008845f
C585 B.n545 VSUBS 0.008845f
C586 B.n546 VSUBS 0.008845f
C587 B.n547 VSUBS 0.008845f
C588 B.n548 VSUBS 0.008845f
C589 B.n549 VSUBS 0.008845f
C590 B.n550 VSUBS 0.008389f
C591 B.n551 VSUBS 0.008845f
C592 B.n552 VSUBS 0.008845f
C593 B.n553 VSUBS 0.008845f
C594 B.n554 VSUBS 0.008845f
C595 B.n555 VSUBS 0.008845f
C596 B.n556 VSUBS 0.008845f
C597 B.n557 VSUBS 0.008845f
C598 B.n558 VSUBS 0.008845f
C599 B.n559 VSUBS 0.008845f
C600 B.n560 VSUBS 0.008845f
C601 B.n561 VSUBS 0.008845f
C602 B.n562 VSUBS 0.008845f
C603 B.n563 VSUBS 0.008845f
C604 B.n564 VSUBS 0.008845f
C605 B.n565 VSUBS 0.008845f
C606 B.n566 VSUBS 0.004877f
C607 B.n567 VSUBS 0.020492f
C608 B.n568 VSUBS 0.008389f
C609 B.n569 VSUBS 0.008845f
C610 B.n570 VSUBS 0.008845f
C611 B.n571 VSUBS 0.008845f
C612 B.n572 VSUBS 0.008845f
C613 B.n573 VSUBS 0.008845f
C614 B.n574 VSUBS 0.008845f
C615 B.n575 VSUBS 0.008845f
C616 B.n576 VSUBS 0.008845f
C617 B.n577 VSUBS 0.008845f
C618 B.n578 VSUBS 0.008845f
C619 B.n579 VSUBS 0.008845f
C620 B.n580 VSUBS 0.008845f
C621 B.n581 VSUBS 0.008845f
C622 B.n582 VSUBS 0.008845f
C623 B.n583 VSUBS 0.008845f
C624 B.n584 VSUBS 0.008845f
C625 B.n585 VSUBS 0.008845f
C626 B.n586 VSUBS 0.008845f
C627 B.n587 VSUBS 0.008845f
C628 B.n588 VSUBS 0.008845f
C629 B.n589 VSUBS 0.008845f
C630 B.n590 VSUBS 0.008845f
C631 B.n591 VSUBS 0.008845f
C632 B.n592 VSUBS 0.008845f
C633 B.n593 VSUBS 0.021561f
C634 B.n594 VSUBS 0.021561f
C635 B.n595 VSUBS 0.0198f
C636 B.n596 VSUBS 0.008845f
C637 B.n597 VSUBS 0.008845f
C638 B.n598 VSUBS 0.008845f
C639 B.n599 VSUBS 0.008845f
C640 B.n600 VSUBS 0.008845f
C641 B.n601 VSUBS 0.008845f
C642 B.n602 VSUBS 0.008845f
C643 B.n603 VSUBS 0.008845f
C644 B.n604 VSUBS 0.008845f
C645 B.n605 VSUBS 0.008845f
C646 B.n606 VSUBS 0.008845f
C647 B.n607 VSUBS 0.008845f
C648 B.n608 VSUBS 0.008845f
C649 B.n609 VSUBS 0.008845f
C650 B.n610 VSUBS 0.008845f
C651 B.n611 VSUBS 0.008845f
C652 B.n612 VSUBS 0.008845f
C653 B.n613 VSUBS 0.008845f
C654 B.n614 VSUBS 0.008845f
C655 B.n615 VSUBS 0.008845f
C656 B.n616 VSUBS 0.008845f
C657 B.n617 VSUBS 0.008845f
C658 B.n618 VSUBS 0.008845f
C659 B.n619 VSUBS 0.008845f
C660 B.n620 VSUBS 0.008845f
C661 B.n621 VSUBS 0.008845f
C662 B.n622 VSUBS 0.008845f
C663 B.n623 VSUBS 0.008845f
C664 B.n624 VSUBS 0.008845f
C665 B.n625 VSUBS 0.008845f
C666 B.n626 VSUBS 0.008845f
C667 B.n627 VSUBS 0.008845f
C668 B.n628 VSUBS 0.008845f
C669 B.n629 VSUBS 0.008845f
C670 B.n630 VSUBS 0.008845f
C671 B.n631 VSUBS 0.008845f
C672 B.n632 VSUBS 0.008845f
C673 B.n633 VSUBS 0.008845f
C674 B.n634 VSUBS 0.008845f
C675 B.n635 VSUBS 0.008845f
C676 B.n636 VSUBS 0.008845f
C677 B.n637 VSUBS 0.008845f
C678 B.n638 VSUBS 0.008845f
C679 B.n639 VSUBS 0.008845f
C680 B.n640 VSUBS 0.008845f
C681 B.n641 VSUBS 0.008845f
C682 B.n642 VSUBS 0.008845f
C683 B.n643 VSUBS 0.008845f
C684 B.n644 VSUBS 0.008845f
C685 B.n645 VSUBS 0.008845f
C686 B.n646 VSUBS 0.008845f
C687 B.n647 VSUBS 0.008845f
C688 B.n648 VSUBS 0.008845f
C689 B.n649 VSUBS 0.008845f
C690 B.n650 VSUBS 0.008845f
C691 B.n651 VSUBS 0.008845f
C692 B.n652 VSUBS 0.008845f
C693 B.n653 VSUBS 0.008845f
C694 B.n654 VSUBS 0.008845f
C695 B.n655 VSUBS 0.008845f
C696 B.n656 VSUBS 0.008845f
C697 B.n657 VSUBS 0.008845f
C698 B.n658 VSUBS 0.008845f
C699 B.n659 VSUBS 0.008845f
C700 B.n660 VSUBS 0.008845f
C701 B.n661 VSUBS 0.008845f
C702 B.n662 VSUBS 0.008845f
C703 B.n663 VSUBS 0.008845f
C704 B.n664 VSUBS 0.008845f
C705 B.n665 VSUBS 0.008845f
C706 B.n666 VSUBS 0.008845f
C707 B.n667 VSUBS 0.008845f
C708 B.n668 VSUBS 0.008845f
C709 B.n669 VSUBS 0.008845f
C710 B.n670 VSUBS 0.008845f
C711 B.n671 VSUBS 0.008845f
C712 B.n672 VSUBS 0.008845f
C713 B.n673 VSUBS 0.008845f
C714 B.n674 VSUBS 0.008845f
C715 B.n675 VSUBS 0.008845f
C716 B.n676 VSUBS 0.008845f
C717 B.n677 VSUBS 0.008845f
C718 B.n678 VSUBS 0.008845f
C719 B.n679 VSUBS 0.008845f
C720 B.n680 VSUBS 0.008845f
C721 B.n681 VSUBS 0.008845f
C722 B.n682 VSUBS 0.008845f
C723 B.n683 VSUBS 0.008845f
C724 B.n684 VSUBS 0.008845f
C725 B.n685 VSUBS 0.008845f
C726 B.n686 VSUBS 0.008845f
C727 B.n687 VSUBS 0.020027f
C728 VDD1.n0 VSUBS 0.036145f
C729 VDD1.n1 VSUBS 0.032894f
C730 VDD1.n2 VSUBS 0.017676f
C731 VDD1.n3 VSUBS 0.041779f
C732 VDD1.n4 VSUBS 0.018715f
C733 VDD1.n5 VSUBS 0.127945f
C734 VDD1.t7 VSUBS 0.092617f
C735 VDD1.n6 VSUBS 0.031334f
C736 VDD1.n7 VSUBS 0.026278f
C737 VDD1.n8 VSUBS 0.017676f
C738 VDD1.n9 VSUBS 0.446372f
C739 VDD1.n10 VSUBS 0.032894f
C740 VDD1.n11 VSUBS 0.017676f
C741 VDD1.n12 VSUBS 0.018715f
C742 VDD1.n13 VSUBS 0.041779f
C743 VDD1.n14 VSUBS 0.101149f
C744 VDD1.n15 VSUBS 0.018715f
C745 VDD1.n16 VSUBS 0.017676f
C746 VDD1.n17 VSUBS 0.081874f
C747 VDD1.n18 VSUBS 0.090137f
C748 VDD1.t2 VSUBS 0.103195f
C749 VDD1.t8 VSUBS 0.103195f
C750 VDD1.n19 VSUBS 0.601799f
C751 VDD1.n20 VSUBS 1.13906f
C752 VDD1.n21 VSUBS 0.036145f
C753 VDD1.n22 VSUBS 0.032894f
C754 VDD1.n23 VSUBS 0.017676f
C755 VDD1.n24 VSUBS 0.041779f
C756 VDD1.n25 VSUBS 0.018715f
C757 VDD1.n26 VSUBS 0.127945f
C758 VDD1.t5 VSUBS 0.092617f
C759 VDD1.n27 VSUBS 0.031334f
C760 VDD1.n28 VSUBS 0.026278f
C761 VDD1.n29 VSUBS 0.017676f
C762 VDD1.n30 VSUBS 0.446372f
C763 VDD1.n31 VSUBS 0.032894f
C764 VDD1.n32 VSUBS 0.017676f
C765 VDD1.n33 VSUBS 0.018715f
C766 VDD1.n34 VSUBS 0.041779f
C767 VDD1.n35 VSUBS 0.101149f
C768 VDD1.n36 VSUBS 0.018715f
C769 VDD1.n37 VSUBS 0.017676f
C770 VDD1.n38 VSUBS 0.081874f
C771 VDD1.n39 VSUBS 0.090137f
C772 VDD1.t0 VSUBS 0.103195f
C773 VDD1.t9 VSUBS 0.103195f
C774 VDD1.n40 VSUBS 0.601796f
C775 VDD1.n41 VSUBS 1.12831f
C776 VDD1.t6 VSUBS 0.103195f
C777 VDD1.t3 VSUBS 0.103195f
C778 VDD1.n42 VSUBS 0.617067f
C779 VDD1.n43 VSUBS 3.59587f
C780 VDD1.t4 VSUBS 0.103195f
C781 VDD1.t1 VSUBS 0.103195f
C782 VDD1.n44 VSUBS 0.601796f
C783 VDD1.n45 VSUBS 3.59362f
C784 VP.n0 VSUBS 0.060727f
C785 VP.t6 VSUBS 1.25579f
C786 VP.n1 VSUBS 0.090792f
C787 VP.n2 VSUBS 0.046061f
C788 VP.t3 VSUBS 1.25579f
C789 VP.n3 VSUBS 0.500185f
C790 VP.n4 VSUBS 0.046061f
C791 VP.n5 VSUBS 0.037253f
C792 VP.n6 VSUBS 0.046061f
C793 VP.t0 VSUBS 1.25579f
C794 VP.n7 VSUBS 0.085846f
C795 VP.n8 VSUBS 0.046061f
C796 VP.n9 VSUBS 0.085846f
C797 VP.n10 VSUBS 0.046061f
C798 VP.t9 VSUBS 1.25579f
C799 VP.n11 VSUBS 0.037371f
C800 VP.n12 VSUBS 0.046061f
C801 VP.t4 VSUBS 1.25579f
C802 VP.n13 VSUBS 0.63765f
C803 VP.n14 VSUBS 0.060727f
C804 VP.t8 VSUBS 1.25579f
C805 VP.n15 VSUBS 0.090792f
C806 VP.n16 VSUBS 0.046061f
C807 VP.t5 VSUBS 1.25579f
C808 VP.n17 VSUBS 0.500185f
C809 VP.n18 VSUBS 0.046061f
C810 VP.n19 VSUBS 0.037253f
C811 VP.n20 VSUBS 0.046061f
C812 VP.t1 VSUBS 1.25579f
C813 VP.n21 VSUBS 0.085846f
C814 VP.n22 VSUBS 0.046061f
C815 VP.n23 VSUBS 0.085846f
C816 VP.t2 VSUBS 1.61602f
C817 VP.n24 VSUBS 0.618804f
C818 VP.t7 VSUBS 1.25579f
C819 VP.n25 VSUBS 0.61941f
C820 VP.n26 VSUBS 0.044311f
C821 VP.n27 VSUBS 0.447702f
C822 VP.n28 VSUBS 0.046061f
C823 VP.n29 VSUBS 0.046061f
C824 VP.n30 VSUBS 0.091311f
C825 VP.n31 VSUBS 0.037253f
C826 VP.n32 VSUBS 0.091773f
C827 VP.n33 VSUBS 0.046061f
C828 VP.n34 VSUBS 0.046061f
C829 VP.n35 VSUBS 0.046061f
C830 VP.n36 VSUBS 0.543649f
C831 VP.n37 VSUBS 0.085846f
C832 VP.n38 VSUBS 0.091773f
C833 VP.n39 VSUBS 0.046061f
C834 VP.n40 VSUBS 0.046061f
C835 VP.n41 VSUBS 0.046061f
C836 VP.n42 VSUBS 0.091311f
C837 VP.n43 VSUBS 0.085846f
C838 VP.n44 VSUBS 0.044311f
C839 VP.n45 VSUBS 0.046061f
C840 VP.n46 VSUBS 0.046061f
C841 VP.n47 VSUBS 0.084998f
C842 VP.n48 VSUBS 0.092173f
C843 VP.n49 VSUBS 0.037371f
C844 VP.n50 VSUBS 0.046061f
C845 VP.n51 VSUBS 0.046061f
C846 VP.n52 VSUBS 0.046061f
C847 VP.n53 VSUBS 0.085846f
C848 VP.n54 VSUBS 0.045159f
C849 VP.n55 VSUBS 0.63765f
C850 VP.n56 VSUBS 2.37318f
C851 VP.n57 VSUBS 2.40813f
C852 VP.n58 VSUBS 0.060727f
C853 VP.n59 VSUBS 0.045159f
C854 VP.n60 VSUBS 0.085846f
C855 VP.n61 VSUBS 0.090792f
C856 VP.n62 VSUBS 0.046061f
C857 VP.n63 VSUBS 0.046061f
C858 VP.n64 VSUBS 0.046061f
C859 VP.n65 VSUBS 0.092173f
C860 VP.n66 VSUBS 0.084998f
C861 VP.n67 VSUBS 0.500185f
C862 VP.n68 VSUBS 0.044311f
C863 VP.n69 VSUBS 0.046061f
C864 VP.n70 VSUBS 0.046061f
C865 VP.n71 VSUBS 0.046061f
C866 VP.n72 VSUBS 0.091311f
C867 VP.n73 VSUBS 0.037253f
C868 VP.n74 VSUBS 0.091773f
C869 VP.n75 VSUBS 0.046061f
C870 VP.n76 VSUBS 0.046061f
C871 VP.n77 VSUBS 0.046061f
C872 VP.n78 VSUBS 0.543649f
C873 VP.n79 VSUBS 0.085846f
C874 VP.n80 VSUBS 0.091773f
C875 VP.n81 VSUBS 0.046061f
C876 VP.n82 VSUBS 0.046061f
C877 VP.n83 VSUBS 0.046061f
C878 VP.n84 VSUBS 0.091311f
C879 VP.n85 VSUBS 0.085846f
C880 VP.n86 VSUBS 0.044311f
C881 VP.n87 VSUBS 0.046061f
C882 VP.n88 VSUBS 0.046061f
C883 VP.n89 VSUBS 0.084998f
C884 VP.n90 VSUBS 0.092173f
C885 VP.n91 VSUBS 0.037371f
C886 VP.n92 VSUBS 0.046061f
C887 VP.n93 VSUBS 0.046061f
C888 VP.n94 VSUBS 0.046061f
C889 VP.n95 VSUBS 0.085846f
C890 VP.n96 VSUBS 0.045159f
C891 VP.n97 VSUBS 0.63765f
C892 VP.n98 VSUBS 0.085349f
C893 VTAIL.t10 VSUBS 0.107452f
C894 VTAIL.t12 VSUBS 0.107452f
C895 VTAIL.n0 VSUBS 0.546688f
C896 VTAIL.n1 VSUBS 0.932578f
C897 VTAIL.n2 VSUBS 0.037636f
C898 VTAIL.n3 VSUBS 0.034251f
C899 VTAIL.n4 VSUBS 0.018405f
C900 VTAIL.n5 VSUBS 0.043502f
C901 VTAIL.n6 VSUBS 0.019488f
C902 VTAIL.n7 VSUBS 0.133223f
C903 VTAIL.t2 VSUBS 0.096438f
C904 VTAIL.n8 VSUBS 0.032627f
C905 VTAIL.n9 VSUBS 0.027362f
C906 VTAIL.n10 VSUBS 0.018405f
C907 VTAIL.n11 VSUBS 0.464787f
C908 VTAIL.n12 VSUBS 0.034251f
C909 VTAIL.n13 VSUBS 0.018405f
C910 VTAIL.n14 VSUBS 0.019488f
C911 VTAIL.n15 VSUBS 0.043502f
C912 VTAIL.n16 VSUBS 0.105322f
C913 VTAIL.n17 VSUBS 0.019488f
C914 VTAIL.n18 VSUBS 0.018405f
C915 VTAIL.n19 VSUBS 0.085252f
C916 VTAIL.n20 VSUBS 0.053146f
C917 VTAIL.n21 VSUBS 0.514107f
C918 VTAIL.t8 VSUBS 0.107452f
C919 VTAIL.t1 VSUBS 0.107452f
C920 VTAIL.n22 VSUBS 0.546688f
C921 VTAIL.n23 VSUBS 1.08908f
C922 VTAIL.t3 VSUBS 0.107452f
C923 VTAIL.t6 VSUBS 0.107452f
C924 VTAIL.n24 VSUBS 0.546688f
C925 VTAIL.n25 VSUBS 2.21843f
C926 VTAIL.t14 VSUBS 0.107452f
C927 VTAIL.t17 VSUBS 0.107452f
C928 VTAIL.n26 VSUBS 0.546692f
C929 VTAIL.n27 VSUBS 2.21842f
C930 VTAIL.t13 VSUBS 0.107452f
C931 VTAIL.t9 VSUBS 0.107452f
C932 VTAIL.n28 VSUBS 0.546692f
C933 VTAIL.n29 VSUBS 1.08908f
C934 VTAIL.n30 VSUBS 0.037636f
C935 VTAIL.n31 VSUBS 0.034251f
C936 VTAIL.n32 VSUBS 0.018405f
C937 VTAIL.n33 VSUBS 0.043502f
C938 VTAIL.n34 VSUBS 0.019488f
C939 VTAIL.n35 VSUBS 0.133223f
C940 VTAIL.t15 VSUBS 0.096438f
C941 VTAIL.n36 VSUBS 0.032627f
C942 VTAIL.n37 VSUBS 0.027362f
C943 VTAIL.n38 VSUBS 0.018405f
C944 VTAIL.n39 VSUBS 0.464787f
C945 VTAIL.n40 VSUBS 0.034251f
C946 VTAIL.n41 VSUBS 0.018405f
C947 VTAIL.n42 VSUBS 0.019488f
C948 VTAIL.n43 VSUBS 0.043502f
C949 VTAIL.n44 VSUBS 0.105322f
C950 VTAIL.n45 VSUBS 0.019488f
C951 VTAIL.n46 VSUBS 0.018405f
C952 VTAIL.n47 VSUBS 0.085252f
C953 VTAIL.n48 VSUBS 0.053146f
C954 VTAIL.n49 VSUBS 0.514107f
C955 VTAIL.t7 VSUBS 0.107452f
C956 VTAIL.t19 VSUBS 0.107452f
C957 VTAIL.n50 VSUBS 0.546692f
C958 VTAIL.n51 VSUBS 0.997746f
C959 VTAIL.t0 VSUBS 0.107452f
C960 VTAIL.t4 VSUBS 0.107452f
C961 VTAIL.n52 VSUBS 0.546692f
C962 VTAIL.n53 VSUBS 1.08908f
C963 VTAIL.n54 VSUBS 0.037636f
C964 VTAIL.n55 VSUBS 0.034251f
C965 VTAIL.n56 VSUBS 0.018405f
C966 VTAIL.n57 VSUBS 0.043502f
C967 VTAIL.n58 VSUBS 0.019488f
C968 VTAIL.n59 VSUBS 0.133223f
C969 VTAIL.t5 VSUBS 0.096438f
C970 VTAIL.n60 VSUBS 0.032627f
C971 VTAIL.n61 VSUBS 0.027362f
C972 VTAIL.n62 VSUBS 0.018405f
C973 VTAIL.n63 VSUBS 0.464787f
C974 VTAIL.n64 VSUBS 0.034251f
C975 VTAIL.n65 VSUBS 0.018405f
C976 VTAIL.n66 VSUBS 0.019488f
C977 VTAIL.n67 VSUBS 0.043502f
C978 VTAIL.n68 VSUBS 0.105322f
C979 VTAIL.n69 VSUBS 0.019488f
C980 VTAIL.n70 VSUBS 0.018405f
C981 VTAIL.n71 VSUBS 0.085252f
C982 VTAIL.n72 VSUBS 0.053146f
C983 VTAIL.n73 VSUBS 1.44841f
C984 VTAIL.n74 VSUBS 0.037636f
C985 VTAIL.n75 VSUBS 0.034251f
C986 VTAIL.n76 VSUBS 0.018405f
C987 VTAIL.n77 VSUBS 0.043502f
C988 VTAIL.n78 VSUBS 0.019488f
C989 VTAIL.n79 VSUBS 0.133223f
C990 VTAIL.t11 VSUBS 0.096438f
C991 VTAIL.n80 VSUBS 0.032627f
C992 VTAIL.n81 VSUBS 0.027362f
C993 VTAIL.n82 VSUBS 0.018405f
C994 VTAIL.n83 VSUBS 0.464787f
C995 VTAIL.n84 VSUBS 0.034251f
C996 VTAIL.n85 VSUBS 0.018405f
C997 VTAIL.n86 VSUBS 0.019488f
C998 VTAIL.n87 VSUBS 0.043502f
C999 VTAIL.n88 VSUBS 0.105322f
C1000 VTAIL.n89 VSUBS 0.019488f
C1001 VTAIL.n90 VSUBS 0.018405f
C1002 VTAIL.n91 VSUBS 0.085252f
C1003 VTAIL.n92 VSUBS 0.053146f
C1004 VTAIL.n93 VSUBS 1.44841f
C1005 VTAIL.t16 VSUBS 0.107452f
C1006 VTAIL.t18 VSUBS 0.107452f
C1007 VTAIL.n94 VSUBS 0.546688f
C1008 VTAIL.n95 VSUBS 0.867882f
C1009 VDD2.n0 VSUBS 0.035728f
C1010 VDD2.n1 VSUBS 0.032515f
C1011 VDD2.n2 VSUBS 0.017472f
C1012 VDD2.n3 VSUBS 0.041297f
C1013 VDD2.n4 VSUBS 0.0185f
C1014 VDD2.n5 VSUBS 0.126469f
C1015 VDD2.t7 VSUBS 0.091549f
C1016 VDD2.n6 VSUBS 0.030973f
C1017 VDD2.n7 VSUBS 0.025975f
C1018 VDD2.n8 VSUBS 0.017472f
C1019 VDD2.n9 VSUBS 0.441224f
C1020 VDD2.n10 VSUBS 0.032515f
C1021 VDD2.n11 VSUBS 0.017472f
C1022 VDD2.n12 VSUBS 0.0185f
C1023 VDD2.n13 VSUBS 0.041297f
C1024 VDD2.n14 VSUBS 0.099982f
C1025 VDD2.n15 VSUBS 0.0185f
C1026 VDD2.n16 VSUBS 0.017472f
C1027 VDD2.n17 VSUBS 0.08093f
C1028 VDD2.n18 VSUBS 0.089097f
C1029 VDD2.t1 VSUBS 0.102005f
C1030 VDD2.t9 VSUBS 0.102005f
C1031 VDD2.n19 VSUBS 0.594855f
C1032 VDD2.n20 VSUBS 1.1153f
C1033 VDD2.t6 VSUBS 0.102005f
C1034 VDD2.t0 VSUBS 0.102005f
C1035 VDD2.n21 VSUBS 0.609951f
C1036 VDD2.n22 VSUBS 3.39808f
C1037 VDD2.n23 VSUBS 0.035728f
C1038 VDD2.n24 VSUBS 0.032515f
C1039 VDD2.n25 VSUBS 0.017472f
C1040 VDD2.n26 VSUBS 0.041297f
C1041 VDD2.n27 VSUBS 0.0185f
C1042 VDD2.n28 VSUBS 0.126469f
C1043 VDD2.t2 VSUBS 0.091549f
C1044 VDD2.n29 VSUBS 0.030973f
C1045 VDD2.n30 VSUBS 0.025975f
C1046 VDD2.n31 VSUBS 0.017472f
C1047 VDD2.n32 VSUBS 0.441224f
C1048 VDD2.n33 VSUBS 0.032515f
C1049 VDD2.n34 VSUBS 0.017472f
C1050 VDD2.n35 VSUBS 0.0185f
C1051 VDD2.n36 VSUBS 0.041297f
C1052 VDD2.n37 VSUBS 0.099982f
C1053 VDD2.n38 VSUBS 0.0185f
C1054 VDD2.n39 VSUBS 0.017472f
C1055 VDD2.n40 VSUBS 0.08093f
C1056 VDD2.n41 VSUBS 0.072861f
C1057 VDD2.n42 VSUBS 2.98496f
C1058 VDD2.t4 VSUBS 0.102005f
C1059 VDD2.t3 VSUBS 0.102005f
C1060 VDD2.n43 VSUBS 0.594858f
C1061 VDD2.n44 VSUBS 0.804384f
C1062 VDD2.t5 VSUBS 0.102005f
C1063 VDD2.t8 VSUBS 0.102005f
C1064 VDD2.n45 VSUBS 0.609917f
C1065 VN.n0 VSUBS 0.053721f
C1066 VN.t7 VSUBS 1.11091f
C1067 VN.n1 VSUBS 0.080317f
C1068 VN.n2 VSUBS 0.040747f
C1069 VN.t0 VSUBS 1.11091f
C1070 VN.n3 VSUBS 0.442479f
C1071 VN.n4 VSUBS 0.040747f
C1072 VN.n5 VSUBS 0.032955f
C1073 VN.n6 VSUBS 0.040747f
C1074 VN.t2 VSUBS 1.11091f
C1075 VN.n7 VSUBS 0.075942f
C1076 VN.n8 VSUBS 0.040747f
C1077 VN.n9 VSUBS 0.075942f
C1078 VN.t8 VSUBS 1.42958f
C1079 VN.n10 VSUBS 0.547412f
C1080 VN.t6 VSUBS 1.11091f
C1081 VN.n11 VSUBS 0.547948f
C1082 VN.n12 VSUBS 0.039199f
C1083 VN.n13 VSUBS 0.39605f
C1084 VN.n14 VSUBS 0.040747f
C1085 VN.n15 VSUBS 0.040747f
C1086 VN.n16 VSUBS 0.080776f
C1087 VN.n17 VSUBS 0.032955f
C1088 VN.n18 VSUBS 0.081185f
C1089 VN.n19 VSUBS 0.040747f
C1090 VN.n20 VSUBS 0.040747f
C1091 VN.n21 VSUBS 0.040747f
C1092 VN.n22 VSUBS 0.480928f
C1093 VN.n23 VSUBS 0.075942f
C1094 VN.n24 VSUBS 0.081185f
C1095 VN.n25 VSUBS 0.040747f
C1096 VN.n26 VSUBS 0.040747f
C1097 VN.n27 VSUBS 0.040747f
C1098 VN.n28 VSUBS 0.080776f
C1099 VN.n29 VSUBS 0.075942f
C1100 VN.n30 VSUBS 0.039199f
C1101 VN.n31 VSUBS 0.040747f
C1102 VN.n32 VSUBS 0.040747f
C1103 VN.n33 VSUBS 0.075192f
C1104 VN.n34 VSUBS 0.081539f
C1105 VN.n35 VSUBS 0.03306f
C1106 VN.n36 VSUBS 0.040747f
C1107 VN.n37 VSUBS 0.040747f
C1108 VN.n38 VSUBS 0.040747f
C1109 VN.n39 VSUBS 0.075942f
C1110 VN.n40 VSUBS 0.039949f
C1111 VN.n41 VSUBS 0.564084f
C1112 VN.n42 VSUBS 0.075502f
C1113 VN.n43 VSUBS 0.053721f
C1114 VN.t4 VSUBS 1.11091f
C1115 VN.n44 VSUBS 0.080317f
C1116 VN.n45 VSUBS 0.040747f
C1117 VN.t1 VSUBS 1.11091f
C1118 VN.n46 VSUBS 0.442479f
C1119 VN.n47 VSUBS 0.040747f
C1120 VN.n48 VSUBS 0.032955f
C1121 VN.n49 VSUBS 0.040747f
C1122 VN.t5 VSUBS 1.11091f
C1123 VN.n50 VSUBS 0.075942f
C1124 VN.n51 VSUBS 0.040747f
C1125 VN.n52 VSUBS 0.075942f
C1126 VN.t3 VSUBS 1.42958f
C1127 VN.n53 VSUBS 0.547412f
C1128 VN.t9 VSUBS 1.11091f
C1129 VN.n54 VSUBS 0.547948f
C1130 VN.n55 VSUBS 0.039199f
C1131 VN.n56 VSUBS 0.39605f
C1132 VN.n57 VSUBS 0.040747f
C1133 VN.n58 VSUBS 0.040747f
C1134 VN.n59 VSUBS 0.080776f
C1135 VN.n60 VSUBS 0.032955f
C1136 VN.n61 VSUBS 0.081185f
C1137 VN.n62 VSUBS 0.040747f
C1138 VN.n63 VSUBS 0.040747f
C1139 VN.n64 VSUBS 0.040747f
C1140 VN.n65 VSUBS 0.480928f
C1141 VN.n66 VSUBS 0.075942f
C1142 VN.n67 VSUBS 0.081185f
C1143 VN.n68 VSUBS 0.040747f
C1144 VN.n69 VSUBS 0.040747f
C1145 VN.n70 VSUBS 0.040747f
C1146 VN.n71 VSUBS 0.080776f
C1147 VN.n72 VSUBS 0.075942f
C1148 VN.n73 VSUBS 0.039199f
C1149 VN.n74 VSUBS 0.040747f
C1150 VN.n75 VSUBS 0.040747f
C1151 VN.n76 VSUBS 0.075192f
C1152 VN.n77 VSUBS 0.081539f
C1153 VN.n78 VSUBS 0.03306f
C1154 VN.n79 VSUBS 0.040747f
C1155 VN.n80 VSUBS 0.040747f
C1156 VN.n81 VSUBS 0.040747f
C1157 VN.n82 VSUBS 0.075942f
C1158 VN.n83 VSUBS 0.039949f
C1159 VN.n84 VSUBS 0.564084f
C1160 VN.n85 VSUBS 2.12147f
.ends

