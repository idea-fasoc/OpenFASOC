* NGSPICE file created from diff_pair_sample_1638.ext - technology: sky130A

.subckt diff_pair_sample_1638 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=0.89
X1 VDD1.t1 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=0.89
X2 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=0.89
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=0.89
X4 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=0.89
X5 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=0.89
X6 VTAIL.t5 VP.t2 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=0.89
X7 VTAIL.t3 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=0.89
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=0.89
X9 VDD2.t0 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=0.89
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=0.89
X11 VDD1.t3 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=0.89
R0 VP.n1 VP.t0 491.894
R1 VP.n1 VP.t1 491.844
R2 VP.n3 VP.t2 470.899
R3 VP.n5 VP.t3 470.899
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 88.6318
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VDD1 VDD1.n1 102.362
R14 VDD1 VDD1.n0 61.4481
R15 VDD1.n0 VDD1.t2 1.25764
R16 VDD1.n0 VDD1.t1 1.25764
R17 VDD1.n1 VDD1.t0 1.25764
R18 VDD1.n1 VDD1.t3 1.25764
R19 VTAIL.n5 VTAIL.t7 45.9684
R20 VTAIL.n4 VTAIL.t1 45.9684
R21 VTAIL.n3 VTAIL.t3 45.9684
R22 VTAIL.n7 VTAIL.t2 45.9683
R23 VTAIL.n0 VTAIL.t0 45.9683
R24 VTAIL.n1 VTAIL.t4 45.9683
R25 VTAIL.n2 VTAIL.t5 45.9683
R26 VTAIL.n6 VTAIL.t6 45.9683
R27 VTAIL.n7 VTAIL.n6 26.9962
R28 VTAIL.n3 VTAIL.n2 26.9962
R29 VTAIL.n4 VTAIL.n3 1.05222
R30 VTAIL.n6 VTAIL.n5 1.05222
R31 VTAIL.n2 VTAIL.n1 1.05222
R32 VTAIL VTAIL.n0 0.584552
R33 VTAIL.n5 VTAIL.n4 0.470328
R34 VTAIL.n1 VTAIL.n0 0.470328
R35 VTAIL VTAIL.n7 0.468172
R36 B.n424 B.t15 628.606
R37 B.n421 B.t11 628.606
R38 B.n101 B.t4 628.606
R39 B.n98 B.t8 628.606
R40 B.n738 B.n737 585
R41 B.n739 B.n738 585
R42 B.n326 B.n96 585
R43 B.n325 B.n324 585
R44 B.n323 B.n322 585
R45 B.n321 B.n320 585
R46 B.n319 B.n318 585
R47 B.n317 B.n316 585
R48 B.n315 B.n314 585
R49 B.n313 B.n312 585
R50 B.n311 B.n310 585
R51 B.n309 B.n308 585
R52 B.n307 B.n306 585
R53 B.n305 B.n304 585
R54 B.n303 B.n302 585
R55 B.n301 B.n300 585
R56 B.n299 B.n298 585
R57 B.n297 B.n296 585
R58 B.n295 B.n294 585
R59 B.n293 B.n292 585
R60 B.n291 B.n290 585
R61 B.n289 B.n288 585
R62 B.n287 B.n286 585
R63 B.n285 B.n284 585
R64 B.n283 B.n282 585
R65 B.n281 B.n280 585
R66 B.n279 B.n278 585
R67 B.n277 B.n276 585
R68 B.n275 B.n274 585
R69 B.n273 B.n272 585
R70 B.n271 B.n270 585
R71 B.n269 B.n268 585
R72 B.n267 B.n266 585
R73 B.n265 B.n264 585
R74 B.n263 B.n262 585
R75 B.n261 B.n260 585
R76 B.n259 B.n258 585
R77 B.n257 B.n256 585
R78 B.n255 B.n254 585
R79 B.n253 B.n252 585
R80 B.n251 B.n250 585
R81 B.n249 B.n248 585
R82 B.n247 B.n246 585
R83 B.n245 B.n244 585
R84 B.n243 B.n242 585
R85 B.n241 B.n240 585
R86 B.n239 B.n238 585
R87 B.n237 B.n236 585
R88 B.n235 B.n234 585
R89 B.n233 B.n232 585
R90 B.n231 B.n230 585
R91 B.n229 B.n228 585
R92 B.n227 B.n226 585
R93 B.n225 B.n224 585
R94 B.n223 B.n222 585
R95 B.n221 B.n220 585
R96 B.n219 B.n218 585
R97 B.n217 B.n216 585
R98 B.n215 B.n214 585
R99 B.n213 B.n212 585
R100 B.n211 B.n210 585
R101 B.n209 B.n208 585
R102 B.n207 B.n206 585
R103 B.n204 B.n203 585
R104 B.n202 B.n201 585
R105 B.n200 B.n199 585
R106 B.n198 B.n197 585
R107 B.n196 B.n195 585
R108 B.n194 B.n193 585
R109 B.n192 B.n191 585
R110 B.n190 B.n189 585
R111 B.n188 B.n187 585
R112 B.n186 B.n185 585
R113 B.n184 B.n183 585
R114 B.n182 B.n181 585
R115 B.n180 B.n179 585
R116 B.n178 B.n177 585
R117 B.n176 B.n175 585
R118 B.n174 B.n173 585
R119 B.n172 B.n171 585
R120 B.n170 B.n169 585
R121 B.n168 B.n167 585
R122 B.n166 B.n165 585
R123 B.n164 B.n163 585
R124 B.n162 B.n161 585
R125 B.n160 B.n159 585
R126 B.n158 B.n157 585
R127 B.n156 B.n155 585
R128 B.n154 B.n153 585
R129 B.n152 B.n151 585
R130 B.n150 B.n149 585
R131 B.n148 B.n147 585
R132 B.n146 B.n145 585
R133 B.n144 B.n143 585
R134 B.n142 B.n141 585
R135 B.n140 B.n139 585
R136 B.n138 B.n137 585
R137 B.n136 B.n135 585
R138 B.n134 B.n133 585
R139 B.n132 B.n131 585
R140 B.n130 B.n129 585
R141 B.n128 B.n127 585
R142 B.n126 B.n125 585
R143 B.n124 B.n123 585
R144 B.n122 B.n121 585
R145 B.n120 B.n119 585
R146 B.n118 B.n117 585
R147 B.n116 B.n115 585
R148 B.n114 B.n113 585
R149 B.n112 B.n111 585
R150 B.n110 B.n109 585
R151 B.n108 B.n107 585
R152 B.n106 B.n105 585
R153 B.n104 B.n103 585
R154 B.n39 B.n38 585
R155 B.n742 B.n741 585
R156 B.n736 B.n97 585
R157 B.n97 B.n36 585
R158 B.n735 B.n35 585
R159 B.n746 B.n35 585
R160 B.n734 B.n34 585
R161 B.n747 B.n34 585
R162 B.n733 B.n33 585
R163 B.n748 B.n33 585
R164 B.n732 B.n731 585
R165 B.n731 B.n29 585
R166 B.n730 B.n28 585
R167 B.n754 B.n28 585
R168 B.n729 B.n27 585
R169 B.n755 B.n27 585
R170 B.n728 B.n26 585
R171 B.n756 B.n26 585
R172 B.n727 B.n726 585
R173 B.n726 B.n22 585
R174 B.n725 B.n21 585
R175 B.n762 B.n21 585
R176 B.n724 B.n20 585
R177 B.n763 B.n20 585
R178 B.n723 B.n19 585
R179 B.n764 B.n19 585
R180 B.n722 B.n721 585
R181 B.n721 B.n18 585
R182 B.n720 B.n14 585
R183 B.n770 B.n14 585
R184 B.n719 B.n13 585
R185 B.n771 B.n13 585
R186 B.n718 B.n12 585
R187 B.n772 B.n12 585
R188 B.n717 B.n716 585
R189 B.n716 B.n8 585
R190 B.n715 B.n7 585
R191 B.n778 B.n7 585
R192 B.n714 B.n6 585
R193 B.n779 B.n6 585
R194 B.n713 B.n5 585
R195 B.n780 B.n5 585
R196 B.n712 B.n711 585
R197 B.n711 B.n4 585
R198 B.n710 B.n327 585
R199 B.n710 B.n709 585
R200 B.n700 B.n328 585
R201 B.n329 B.n328 585
R202 B.n702 B.n701 585
R203 B.n703 B.n702 585
R204 B.n699 B.n334 585
R205 B.n334 B.n333 585
R206 B.n698 B.n697 585
R207 B.n697 B.n696 585
R208 B.n336 B.n335 585
R209 B.n689 B.n336 585
R210 B.n688 B.n687 585
R211 B.n690 B.n688 585
R212 B.n686 B.n341 585
R213 B.n341 B.n340 585
R214 B.n685 B.n684 585
R215 B.n684 B.n683 585
R216 B.n343 B.n342 585
R217 B.n344 B.n343 585
R218 B.n676 B.n675 585
R219 B.n677 B.n676 585
R220 B.n674 B.n349 585
R221 B.n349 B.n348 585
R222 B.n673 B.n672 585
R223 B.n672 B.n671 585
R224 B.n351 B.n350 585
R225 B.n352 B.n351 585
R226 B.n664 B.n663 585
R227 B.n665 B.n664 585
R228 B.n662 B.n357 585
R229 B.n357 B.n356 585
R230 B.n661 B.n660 585
R231 B.n660 B.n659 585
R232 B.n359 B.n358 585
R233 B.n360 B.n359 585
R234 B.n655 B.n654 585
R235 B.n363 B.n362 585
R236 B.n651 B.n650 585
R237 B.n652 B.n651 585
R238 B.n649 B.n420 585
R239 B.n648 B.n647 585
R240 B.n646 B.n645 585
R241 B.n644 B.n643 585
R242 B.n642 B.n641 585
R243 B.n640 B.n639 585
R244 B.n638 B.n637 585
R245 B.n636 B.n635 585
R246 B.n634 B.n633 585
R247 B.n632 B.n631 585
R248 B.n630 B.n629 585
R249 B.n628 B.n627 585
R250 B.n626 B.n625 585
R251 B.n624 B.n623 585
R252 B.n622 B.n621 585
R253 B.n620 B.n619 585
R254 B.n618 B.n617 585
R255 B.n616 B.n615 585
R256 B.n614 B.n613 585
R257 B.n612 B.n611 585
R258 B.n610 B.n609 585
R259 B.n608 B.n607 585
R260 B.n606 B.n605 585
R261 B.n604 B.n603 585
R262 B.n602 B.n601 585
R263 B.n600 B.n599 585
R264 B.n598 B.n597 585
R265 B.n596 B.n595 585
R266 B.n594 B.n593 585
R267 B.n592 B.n591 585
R268 B.n590 B.n589 585
R269 B.n588 B.n587 585
R270 B.n586 B.n585 585
R271 B.n584 B.n583 585
R272 B.n582 B.n581 585
R273 B.n580 B.n579 585
R274 B.n578 B.n577 585
R275 B.n576 B.n575 585
R276 B.n574 B.n573 585
R277 B.n572 B.n571 585
R278 B.n570 B.n569 585
R279 B.n568 B.n567 585
R280 B.n566 B.n565 585
R281 B.n564 B.n563 585
R282 B.n562 B.n561 585
R283 B.n560 B.n559 585
R284 B.n558 B.n557 585
R285 B.n556 B.n555 585
R286 B.n554 B.n553 585
R287 B.n552 B.n551 585
R288 B.n550 B.n549 585
R289 B.n548 B.n547 585
R290 B.n546 B.n545 585
R291 B.n544 B.n543 585
R292 B.n542 B.n541 585
R293 B.n540 B.n539 585
R294 B.n538 B.n537 585
R295 B.n536 B.n535 585
R296 B.n534 B.n533 585
R297 B.n531 B.n530 585
R298 B.n529 B.n528 585
R299 B.n527 B.n526 585
R300 B.n525 B.n524 585
R301 B.n523 B.n522 585
R302 B.n521 B.n520 585
R303 B.n519 B.n518 585
R304 B.n517 B.n516 585
R305 B.n515 B.n514 585
R306 B.n513 B.n512 585
R307 B.n511 B.n510 585
R308 B.n509 B.n508 585
R309 B.n507 B.n506 585
R310 B.n505 B.n504 585
R311 B.n503 B.n502 585
R312 B.n501 B.n500 585
R313 B.n499 B.n498 585
R314 B.n497 B.n496 585
R315 B.n495 B.n494 585
R316 B.n493 B.n492 585
R317 B.n491 B.n490 585
R318 B.n489 B.n488 585
R319 B.n487 B.n486 585
R320 B.n485 B.n484 585
R321 B.n483 B.n482 585
R322 B.n481 B.n480 585
R323 B.n479 B.n478 585
R324 B.n477 B.n476 585
R325 B.n475 B.n474 585
R326 B.n473 B.n472 585
R327 B.n471 B.n470 585
R328 B.n469 B.n468 585
R329 B.n467 B.n466 585
R330 B.n465 B.n464 585
R331 B.n463 B.n462 585
R332 B.n461 B.n460 585
R333 B.n459 B.n458 585
R334 B.n457 B.n456 585
R335 B.n455 B.n454 585
R336 B.n453 B.n452 585
R337 B.n451 B.n450 585
R338 B.n449 B.n448 585
R339 B.n447 B.n446 585
R340 B.n445 B.n444 585
R341 B.n443 B.n442 585
R342 B.n441 B.n440 585
R343 B.n439 B.n438 585
R344 B.n437 B.n436 585
R345 B.n435 B.n434 585
R346 B.n433 B.n432 585
R347 B.n431 B.n430 585
R348 B.n429 B.n428 585
R349 B.n427 B.n426 585
R350 B.n656 B.n361 585
R351 B.n361 B.n360 585
R352 B.n658 B.n657 585
R353 B.n659 B.n658 585
R354 B.n355 B.n354 585
R355 B.n356 B.n355 585
R356 B.n667 B.n666 585
R357 B.n666 B.n665 585
R358 B.n668 B.n353 585
R359 B.n353 B.n352 585
R360 B.n670 B.n669 585
R361 B.n671 B.n670 585
R362 B.n347 B.n346 585
R363 B.n348 B.n347 585
R364 B.n679 B.n678 585
R365 B.n678 B.n677 585
R366 B.n680 B.n345 585
R367 B.n345 B.n344 585
R368 B.n682 B.n681 585
R369 B.n683 B.n682 585
R370 B.n339 B.n338 585
R371 B.n340 B.n339 585
R372 B.n692 B.n691 585
R373 B.n691 B.n690 585
R374 B.n693 B.n337 585
R375 B.n689 B.n337 585
R376 B.n695 B.n694 585
R377 B.n696 B.n695 585
R378 B.n332 B.n331 585
R379 B.n333 B.n332 585
R380 B.n705 B.n704 585
R381 B.n704 B.n703 585
R382 B.n706 B.n330 585
R383 B.n330 B.n329 585
R384 B.n708 B.n707 585
R385 B.n709 B.n708 585
R386 B.n2 B.n0 585
R387 B.n4 B.n2 585
R388 B.n3 B.n1 585
R389 B.n779 B.n3 585
R390 B.n777 B.n776 585
R391 B.n778 B.n777 585
R392 B.n775 B.n9 585
R393 B.n9 B.n8 585
R394 B.n774 B.n773 585
R395 B.n773 B.n772 585
R396 B.n11 B.n10 585
R397 B.n771 B.n11 585
R398 B.n769 B.n768 585
R399 B.n770 B.n769 585
R400 B.n767 B.n15 585
R401 B.n18 B.n15 585
R402 B.n766 B.n765 585
R403 B.n765 B.n764 585
R404 B.n17 B.n16 585
R405 B.n763 B.n17 585
R406 B.n761 B.n760 585
R407 B.n762 B.n761 585
R408 B.n759 B.n23 585
R409 B.n23 B.n22 585
R410 B.n758 B.n757 585
R411 B.n757 B.n756 585
R412 B.n25 B.n24 585
R413 B.n755 B.n25 585
R414 B.n753 B.n752 585
R415 B.n754 B.n753 585
R416 B.n751 B.n30 585
R417 B.n30 B.n29 585
R418 B.n750 B.n749 585
R419 B.n749 B.n748 585
R420 B.n32 B.n31 585
R421 B.n747 B.n32 585
R422 B.n745 B.n744 585
R423 B.n746 B.n745 585
R424 B.n743 B.n37 585
R425 B.n37 B.n36 585
R426 B.n782 B.n781 585
R427 B.n781 B.n780 585
R428 B.n654 B.n361 468.476
R429 B.n741 B.n37 468.476
R430 B.n426 B.n359 468.476
R431 B.n738 B.n97 468.476
R432 B.n739 B.n95 256.663
R433 B.n739 B.n94 256.663
R434 B.n739 B.n93 256.663
R435 B.n739 B.n92 256.663
R436 B.n739 B.n91 256.663
R437 B.n739 B.n90 256.663
R438 B.n739 B.n89 256.663
R439 B.n739 B.n88 256.663
R440 B.n739 B.n87 256.663
R441 B.n739 B.n86 256.663
R442 B.n739 B.n85 256.663
R443 B.n739 B.n84 256.663
R444 B.n739 B.n83 256.663
R445 B.n739 B.n82 256.663
R446 B.n739 B.n81 256.663
R447 B.n739 B.n80 256.663
R448 B.n739 B.n79 256.663
R449 B.n739 B.n78 256.663
R450 B.n739 B.n77 256.663
R451 B.n739 B.n76 256.663
R452 B.n739 B.n75 256.663
R453 B.n739 B.n74 256.663
R454 B.n739 B.n73 256.663
R455 B.n739 B.n72 256.663
R456 B.n739 B.n71 256.663
R457 B.n739 B.n70 256.663
R458 B.n739 B.n69 256.663
R459 B.n739 B.n68 256.663
R460 B.n739 B.n67 256.663
R461 B.n739 B.n66 256.663
R462 B.n739 B.n65 256.663
R463 B.n739 B.n64 256.663
R464 B.n739 B.n63 256.663
R465 B.n739 B.n62 256.663
R466 B.n739 B.n61 256.663
R467 B.n739 B.n60 256.663
R468 B.n739 B.n59 256.663
R469 B.n739 B.n58 256.663
R470 B.n739 B.n57 256.663
R471 B.n739 B.n56 256.663
R472 B.n739 B.n55 256.663
R473 B.n739 B.n54 256.663
R474 B.n739 B.n53 256.663
R475 B.n739 B.n52 256.663
R476 B.n739 B.n51 256.663
R477 B.n739 B.n50 256.663
R478 B.n739 B.n49 256.663
R479 B.n739 B.n48 256.663
R480 B.n739 B.n47 256.663
R481 B.n739 B.n46 256.663
R482 B.n739 B.n45 256.663
R483 B.n739 B.n44 256.663
R484 B.n739 B.n43 256.663
R485 B.n739 B.n42 256.663
R486 B.n739 B.n41 256.663
R487 B.n739 B.n40 256.663
R488 B.n740 B.n739 256.663
R489 B.n653 B.n652 256.663
R490 B.n652 B.n364 256.663
R491 B.n652 B.n365 256.663
R492 B.n652 B.n366 256.663
R493 B.n652 B.n367 256.663
R494 B.n652 B.n368 256.663
R495 B.n652 B.n369 256.663
R496 B.n652 B.n370 256.663
R497 B.n652 B.n371 256.663
R498 B.n652 B.n372 256.663
R499 B.n652 B.n373 256.663
R500 B.n652 B.n374 256.663
R501 B.n652 B.n375 256.663
R502 B.n652 B.n376 256.663
R503 B.n652 B.n377 256.663
R504 B.n652 B.n378 256.663
R505 B.n652 B.n379 256.663
R506 B.n652 B.n380 256.663
R507 B.n652 B.n381 256.663
R508 B.n652 B.n382 256.663
R509 B.n652 B.n383 256.663
R510 B.n652 B.n384 256.663
R511 B.n652 B.n385 256.663
R512 B.n652 B.n386 256.663
R513 B.n652 B.n387 256.663
R514 B.n652 B.n388 256.663
R515 B.n652 B.n389 256.663
R516 B.n652 B.n390 256.663
R517 B.n652 B.n391 256.663
R518 B.n652 B.n392 256.663
R519 B.n652 B.n393 256.663
R520 B.n652 B.n394 256.663
R521 B.n652 B.n395 256.663
R522 B.n652 B.n396 256.663
R523 B.n652 B.n397 256.663
R524 B.n652 B.n398 256.663
R525 B.n652 B.n399 256.663
R526 B.n652 B.n400 256.663
R527 B.n652 B.n401 256.663
R528 B.n652 B.n402 256.663
R529 B.n652 B.n403 256.663
R530 B.n652 B.n404 256.663
R531 B.n652 B.n405 256.663
R532 B.n652 B.n406 256.663
R533 B.n652 B.n407 256.663
R534 B.n652 B.n408 256.663
R535 B.n652 B.n409 256.663
R536 B.n652 B.n410 256.663
R537 B.n652 B.n411 256.663
R538 B.n652 B.n412 256.663
R539 B.n652 B.n413 256.663
R540 B.n652 B.n414 256.663
R541 B.n652 B.n415 256.663
R542 B.n652 B.n416 256.663
R543 B.n652 B.n417 256.663
R544 B.n652 B.n418 256.663
R545 B.n652 B.n419 256.663
R546 B.n658 B.n361 163.367
R547 B.n658 B.n355 163.367
R548 B.n666 B.n355 163.367
R549 B.n666 B.n353 163.367
R550 B.n670 B.n353 163.367
R551 B.n670 B.n347 163.367
R552 B.n678 B.n347 163.367
R553 B.n678 B.n345 163.367
R554 B.n682 B.n345 163.367
R555 B.n682 B.n339 163.367
R556 B.n691 B.n339 163.367
R557 B.n691 B.n337 163.367
R558 B.n695 B.n337 163.367
R559 B.n695 B.n332 163.367
R560 B.n704 B.n332 163.367
R561 B.n704 B.n330 163.367
R562 B.n708 B.n330 163.367
R563 B.n708 B.n2 163.367
R564 B.n781 B.n2 163.367
R565 B.n781 B.n3 163.367
R566 B.n777 B.n3 163.367
R567 B.n777 B.n9 163.367
R568 B.n773 B.n9 163.367
R569 B.n773 B.n11 163.367
R570 B.n769 B.n11 163.367
R571 B.n769 B.n15 163.367
R572 B.n765 B.n15 163.367
R573 B.n765 B.n17 163.367
R574 B.n761 B.n17 163.367
R575 B.n761 B.n23 163.367
R576 B.n757 B.n23 163.367
R577 B.n757 B.n25 163.367
R578 B.n753 B.n25 163.367
R579 B.n753 B.n30 163.367
R580 B.n749 B.n30 163.367
R581 B.n749 B.n32 163.367
R582 B.n745 B.n32 163.367
R583 B.n745 B.n37 163.367
R584 B.n651 B.n363 163.367
R585 B.n651 B.n420 163.367
R586 B.n647 B.n646 163.367
R587 B.n643 B.n642 163.367
R588 B.n639 B.n638 163.367
R589 B.n635 B.n634 163.367
R590 B.n631 B.n630 163.367
R591 B.n627 B.n626 163.367
R592 B.n623 B.n622 163.367
R593 B.n619 B.n618 163.367
R594 B.n615 B.n614 163.367
R595 B.n611 B.n610 163.367
R596 B.n607 B.n606 163.367
R597 B.n603 B.n602 163.367
R598 B.n599 B.n598 163.367
R599 B.n595 B.n594 163.367
R600 B.n591 B.n590 163.367
R601 B.n587 B.n586 163.367
R602 B.n583 B.n582 163.367
R603 B.n579 B.n578 163.367
R604 B.n575 B.n574 163.367
R605 B.n571 B.n570 163.367
R606 B.n567 B.n566 163.367
R607 B.n563 B.n562 163.367
R608 B.n559 B.n558 163.367
R609 B.n555 B.n554 163.367
R610 B.n551 B.n550 163.367
R611 B.n547 B.n546 163.367
R612 B.n543 B.n542 163.367
R613 B.n539 B.n538 163.367
R614 B.n535 B.n534 163.367
R615 B.n530 B.n529 163.367
R616 B.n526 B.n525 163.367
R617 B.n522 B.n521 163.367
R618 B.n518 B.n517 163.367
R619 B.n514 B.n513 163.367
R620 B.n510 B.n509 163.367
R621 B.n506 B.n505 163.367
R622 B.n502 B.n501 163.367
R623 B.n498 B.n497 163.367
R624 B.n494 B.n493 163.367
R625 B.n490 B.n489 163.367
R626 B.n486 B.n485 163.367
R627 B.n482 B.n481 163.367
R628 B.n478 B.n477 163.367
R629 B.n474 B.n473 163.367
R630 B.n470 B.n469 163.367
R631 B.n466 B.n465 163.367
R632 B.n462 B.n461 163.367
R633 B.n458 B.n457 163.367
R634 B.n454 B.n453 163.367
R635 B.n450 B.n449 163.367
R636 B.n446 B.n445 163.367
R637 B.n442 B.n441 163.367
R638 B.n438 B.n437 163.367
R639 B.n434 B.n433 163.367
R640 B.n430 B.n429 163.367
R641 B.n660 B.n359 163.367
R642 B.n660 B.n357 163.367
R643 B.n664 B.n357 163.367
R644 B.n664 B.n351 163.367
R645 B.n672 B.n351 163.367
R646 B.n672 B.n349 163.367
R647 B.n676 B.n349 163.367
R648 B.n676 B.n343 163.367
R649 B.n684 B.n343 163.367
R650 B.n684 B.n341 163.367
R651 B.n688 B.n341 163.367
R652 B.n688 B.n336 163.367
R653 B.n697 B.n336 163.367
R654 B.n697 B.n334 163.367
R655 B.n702 B.n334 163.367
R656 B.n702 B.n328 163.367
R657 B.n710 B.n328 163.367
R658 B.n711 B.n710 163.367
R659 B.n711 B.n5 163.367
R660 B.n6 B.n5 163.367
R661 B.n7 B.n6 163.367
R662 B.n716 B.n7 163.367
R663 B.n716 B.n12 163.367
R664 B.n13 B.n12 163.367
R665 B.n14 B.n13 163.367
R666 B.n721 B.n14 163.367
R667 B.n721 B.n19 163.367
R668 B.n20 B.n19 163.367
R669 B.n21 B.n20 163.367
R670 B.n726 B.n21 163.367
R671 B.n726 B.n26 163.367
R672 B.n27 B.n26 163.367
R673 B.n28 B.n27 163.367
R674 B.n731 B.n28 163.367
R675 B.n731 B.n33 163.367
R676 B.n34 B.n33 163.367
R677 B.n35 B.n34 163.367
R678 B.n97 B.n35 163.367
R679 B.n103 B.n39 163.367
R680 B.n107 B.n106 163.367
R681 B.n111 B.n110 163.367
R682 B.n115 B.n114 163.367
R683 B.n119 B.n118 163.367
R684 B.n123 B.n122 163.367
R685 B.n127 B.n126 163.367
R686 B.n131 B.n130 163.367
R687 B.n135 B.n134 163.367
R688 B.n139 B.n138 163.367
R689 B.n143 B.n142 163.367
R690 B.n147 B.n146 163.367
R691 B.n151 B.n150 163.367
R692 B.n155 B.n154 163.367
R693 B.n159 B.n158 163.367
R694 B.n163 B.n162 163.367
R695 B.n167 B.n166 163.367
R696 B.n171 B.n170 163.367
R697 B.n175 B.n174 163.367
R698 B.n179 B.n178 163.367
R699 B.n183 B.n182 163.367
R700 B.n187 B.n186 163.367
R701 B.n191 B.n190 163.367
R702 B.n195 B.n194 163.367
R703 B.n199 B.n198 163.367
R704 B.n203 B.n202 163.367
R705 B.n208 B.n207 163.367
R706 B.n212 B.n211 163.367
R707 B.n216 B.n215 163.367
R708 B.n220 B.n219 163.367
R709 B.n224 B.n223 163.367
R710 B.n228 B.n227 163.367
R711 B.n232 B.n231 163.367
R712 B.n236 B.n235 163.367
R713 B.n240 B.n239 163.367
R714 B.n244 B.n243 163.367
R715 B.n248 B.n247 163.367
R716 B.n252 B.n251 163.367
R717 B.n256 B.n255 163.367
R718 B.n260 B.n259 163.367
R719 B.n264 B.n263 163.367
R720 B.n268 B.n267 163.367
R721 B.n272 B.n271 163.367
R722 B.n276 B.n275 163.367
R723 B.n280 B.n279 163.367
R724 B.n284 B.n283 163.367
R725 B.n288 B.n287 163.367
R726 B.n292 B.n291 163.367
R727 B.n296 B.n295 163.367
R728 B.n300 B.n299 163.367
R729 B.n304 B.n303 163.367
R730 B.n308 B.n307 163.367
R731 B.n312 B.n311 163.367
R732 B.n316 B.n315 163.367
R733 B.n320 B.n319 163.367
R734 B.n324 B.n323 163.367
R735 B.n738 B.n96 163.367
R736 B.n424 B.t17 93.1965
R737 B.n98 B.t9 93.1965
R738 B.n421 B.t14 93.1757
R739 B.n101 B.t6 93.1757
R740 B.n654 B.n653 71.676
R741 B.n420 B.n364 71.676
R742 B.n646 B.n365 71.676
R743 B.n642 B.n366 71.676
R744 B.n638 B.n367 71.676
R745 B.n634 B.n368 71.676
R746 B.n630 B.n369 71.676
R747 B.n626 B.n370 71.676
R748 B.n622 B.n371 71.676
R749 B.n618 B.n372 71.676
R750 B.n614 B.n373 71.676
R751 B.n610 B.n374 71.676
R752 B.n606 B.n375 71.676
R753 B.n602 B.n376 71.676
R754 B.n598 B.n377 71.676
R755 B.n594 B.n378 71.676
R756 B.n590 B.n379 71.676
R757 B.n586 B.n380 71.676
R758 B.n582 B.n381 71.676
R759 B.n578 B.n382 71.676
R760 B.n574 B.n383 71.676
R761 B.n570 B.n384 71.676
R762 B.n566 B.n385 71.676
R763 B.n562 B.n386 71.676
R764 B.n558 B.n387 71.676
R765 B.n554 B.n388 71.676
R766 B.n550 B.n389 71.676
R767 B.n546 B.n390 71.676
R768 B.n542 B.n391 71.676
R769 B.n538 B.n392 71.676
R770 B.n534 B.n393 71.676
R771 B.n529 B.n394 71.676
R772 B.n525 B.n395 71.676
R773 B.n521 B.n396 71.676
R774 B.n517 B.n397 71.676
R775 B.n513 B.n398 71.676
R776 B.n509 B.n399 71.676
R777 B.n505 B.n400 71.676
R778 B.n501 B.n401 71.676
R779 B.n497 B.n402 71.676
R780 B.n493 B.n403 71.676
R781 B.n489 B.n404 71.676
R782 B.n485 B.n405 71.676
R783 B.n481 B.n406 71.676
R784 B.n477 B.n407 71.676
R785 B.n473 B.n408 71.676
R786 B.n469 B.n409 71.676
R787 B.n465 B.n410 71.676
R788 B.n461 B.n411 71.676
R789 B.n457 B.n412 71.676
R790 B.n453 B.n413 71.676
R791 B.n449 B.n414 71.676
R792 B.n445 B.n415 71.676
R793 B.n441 B.n416 71.676
R794 B.n437 B.n417 71.676
R795 B.n433 B.n418 71.676
R796 B.n429 B.n419 71.676
R797 B.n741 B.n740 71.676
R798 B.n103 B.n40 71.676
R799 B.n107 B.n41 71.676
R800 B.n111 B.n42 71.676
R801 B.n115 B.n43 71.676
R802 B.n119 B.n44 71.676
R803 B.n123 B.n45 71.676
R804 B.n127 B.n46 71.676
R805 B.n131 B.n47 71.676
R806 B.n135 B.n48 71.676
R807 B.n139 B.n49 71.676
R808 B.n143 B.n50 71.676
R809 B.n147 B.n51 71.676
R810 B.n151 B.n52 71.676
R811 B.n155 B.n53 71.676
R812 B.n159 B.n54 71.676
R813 B.n163 B.n55 71.676
R814 B.n167 B.n56 71.676
R815 B.n171 B.n57 71.676
R816 B.n175 B.n58 71.676
R817 B.n179 B.n59 71.676
R818 B.n183 B.n60 71.676
R819 B.n187 B.n61 71.676
R820 B.n191 B.n62 71.676
R821 B.n195 B.n63 71.676
R822 B.n199 B.n64 71.676
R823 B.n203 B.n65 71.676
R824 B.n208 B.n66 71.676
R825 B.n212 B.n67 71.676
R826 B.n216 B.n68 71.676
R827 B.n220 B.n69 71.676
R828 B.n224 B.n70 71.676
R829 B.n228 B.n71 71.676
R830 B.n232 B.n72 71.676
R831 B.n236 B.n73 71.676
R832 B.n240 B.n74 71.676
R833 B.n244 B.n75 71.676
R834 B.n248 B.n76 71.676
R835 B.n252 B.n77 71.676
R836 B.n256 B.n78 71.676
R837 B.n260 B.n79 71.676
R838 B.n264 B.n80 71.676
R839 B.n268 B.n81 71.676
R840 B.n272 B.n82 71.676
R841 B.n276 B.n83 71.676
R842 B.n280 B.n84 71.676
R843 B.n284 B.n85 71.676
R844 B.n288 B.n86 71.676
R845 B.n292 B.n87 71.676
R846 B.n296 B.n88 71.676
R847 B.n300 B.n89 71.676
R848 B.n304 B.n90 71.676
R849 B.n308 B.n91 71.676
R850 B.n312 B.n92 71.676
R851 B.n316 B.n93 71.676
R852 B.n320 B.n94 71.676
R853 B.n324 B.n95 71.676
R854 B.n96 B.n95 71.676
R855 B.n323 B.n94 71.676
R856 B.n319 B.n93 71.676
R857 B.n315 B.n92 71.676
R858 B.n311 B.n91 71.676
R859 B.n307 B.n90 71.676
R860 B.n303 B.n89 71.676
R861 B.n299 B.n88 71.676
R862 B.n295 B.n87 71.676
R863 B.n291 B.n86 71.676
R864 B.n287 B.n85 71.676
R865 B.n283 B.n84 71.676
R866 B.n279 B.n83 71.676
R867 B.n275 B.n82 71.676
R868 B.n271 B.n81 71.676
R869 B.n267 B.n80 71.676
R870 B.n263 B.n79 71.676
R871 B.n259 B.n78 71.676
R872 B.n255 B.n77 71.676
R873 B.n251 B.n76 71.676
R874 B.n247 B.n75 71.676
R875 B.n243 B.n74 71.676
R876 B.n239 B.n73 71.676
R877 B.n235 B.n72 71.676
R878 B.n231 B.n71 71.676
R879 B.n227 B.n70 71.676
R880 B.n223 B.n69 71.676
R881 B.n219 B.n68 71.676
R882 B.n215 B.n67 71.676
R883 B.n211 B.n66 71.676
R884 B.n207 B.n65 71.676
R885 B.n202 B.n64 71.676
R886 B.n198 B.n63 71.676
R887 B.n194 B.n62 71.676
R888 B.n190 B.n61 71.676
R889 B.n186 B.n60 71.676
R890 B.n182 B.n59 71.676
R891 B.n178 B.n58 71.676
R892 B.n174 B.n57 71.676
R893 B.n170 B.n56 71.676
R894 B.n166 B.n55 71.676
R895 B.n162 B.n54 71.676
R896 B.n158 B.n53 71.676
R897 B.n154 B.n52 71.676
R898 B.n150 B.n51 71.676
R899 B.n146 B.n50 71.676
R900 B.n142 B.n49 71.676
R901 B.n138 B.n48 71.676
R902 B.n134 B.n47 71.676
R903 B.n130 B.n46 71.676
R904 B.n126 B.n45 71.676
R905 B.n122 B.n44 71.676
R906 B.n118 B.n43 71.676
R907 B.n114 B.n42 71.676
R908 B.n110 B.n41 71.676
R909 B.n106 B.n40 71.676
R910 B.n740 B.n39 71.676
R911 B.n653 B.n363 71.676
R912 B.n647 B.n364 71.676
R913 B.n643 B.n365 71.676
R914 B.n639 B.n366 71.676
R915 B.n635 B.n367 71.676
R916 B.n631 B.n368 71.676
R917 B.n627 B.n369 71.676
R918 B.n623 B.n370 71.676
R919 B.n619 B.n371 71.676
R920 B.n615 B.n372 71.676
R921 B.n611 B.n373 71.676
R922 B.n607 B.n374 71.676
R923 B.n603 B.n375 71.676
R924 B.n599 B.n376 71.676
R925 B.n595 B.n377 71.676
R926 B.n591 B.n378 71.676
R927 B.n587 B.n379 71.676
R928 B.n583 B.n380 71.676
R929 B.n579 B.n381 71.676
R930 B.n575 B.n382 71.676
R931 B.n571 B.n383 71.676
R932 B.n567 B.n384 71.676
R933 B.n563 B.n385 71.676
R934 B.n559 B.n386 71.676
R935 B.n555 B.n387 71.676
R936 B.n551 B.n388 71.676
R937 B.n547 B.n389 71.676
R938 B.n543 B.n390 71.676
R939 B.n539 B.n391 71.676
R940 B.n535 B.n392 71.676
R941 B.n530 B.n393 71.676
R942 B.n526 B.n394 71.676
R943 B.n522 B.n395 71.676
R944 B.n518 B.n396 71.676
R945 B.n514 B.n397 71.676
R946 B.n510 B.n398 71.676
R947 B.n506 B.n399 71.676
R948 B.n502 B.n400 71.676
R949 B.n498 B.n401 71.676
R950 B.n494 B.n402 71.676
R951 B.n490 B.n403 71.676
R952 B.n486 B.n404 71.676
R953 B.n482 B.n405 71.676
R954 B.n478 B.n406 71.676
R955 B.n474 B.n407 71.676
R956 B.n470 B.n408 71.676
R957 B.n466 B.n409 71.676
R958 B.n462 B.n410 71.676
R959 B.n458 B.n411 71.676
R960 B.n454 B.n412 71.676
R961 B.n450 B.n413 71.676
R962 B.n446 B.n414 71.676
R963 B.n442 B.n415 71.676
R964 B.n438 B.n416 71.676
R965 B.n434 B.n417 71.676
R966 B.n430 B.n418 71.676
R967 B.n426 B.n419 71.676
R968 B.n425 B.t16 69.5359
R969 B.n99 B.t10 69.5359
R970 B.n422 B.t13 69.5151
R971 B.n102 B.t7 69.5151
R972 B.n652 B.n360 60.167
R973 B.n739 B.n36 60.167
R974 B.n532 B.n425 59.5399
R975 B.n423 B.n422 59.5399
R976 B.n205 B.n102 59.5399
R977 B.n100 B.n99 59.5399
R978 B.n659 B.n360 35.5772
R979 B.n659 B.n356 35.5772
R980 B.n665 B.n356 35.5772
R981 B.n665 B.n352 35.5772
R982 B.n671 B.n352 35.5772
R983 B.n677 B.n348 35.5772
R984 B.n677 B.n344 35.5772
R985 B.n683 B.n344 35.5772
R986 B.n683 B.n340 35.5772
R987 B.n690 B.n340 35.5772
R988 B.n690 B.n689 35.5772
R989 B.n696 B.n333 35.5772
R990 B.n703 B.n333 35.5772
R991 B.n709 B.n329 35.5772
R992 B.n709 B.n4 35.5772
R993 B.n780 B.n4 35.5772
R994 B.n780 B.n779 35.5772
R995 B.n779 B.n778 35.5772
R996 B.n778 B.n8 35.5772
R997 B.n772 B.n771 35.5772
R998 B.n771 B.n770 35.5772
R999 B.n764 B.n18 35.5772
R1000 B.n764 B.n763 35.5772
R1001 B.n763 B.n762 35.5772
R1002 B.n762 B.n22 35.5772
R1003 B.n756 B.n22 35.5772
R1004 B.n756 B.n755 35.5772
R1005 B.n754 B.n29 35.5772
R1006 B.n748 B.n29 35.5772
R1007 B.n748 B.n747 35.5772
R1008 B.n747 B.n746 35.5772
R1009 B.n746 B.n36 35.5772
R1010 B.n696 B.t3 35.054
R1011 B.n770 B.t2 35.054
R1012 B.n743 B.n742 30.4395
R1013 B.n737 B.n736 30.4395
R1014 B.n427 B.n358 30.4395
R1015 B.n656 B.n655 30.4395
R1016 B.t12 B.n348 27.7294
R1017 B.n755 B.t5 27.7294
R1018 B.n425 B.n424 23.6611
R1019 B.n422 B.n421 23.6611
R1020 B.n102 B.n101 23.6611
R1021 B.n99 B.n98 23.6611
R1022 B.n703 B.t1 21.4512
R1023 B.n772 B.t0 21.4512
R1024 B B.n782 18.0485
R1025 B.t1 B.n329 14.1265
R1026 B.t0 B.n8 14.1265
R1027 B.n742 B.n38 10.6151
R1028 B.n104 B.n38 10.6151
R1029 B.n105 B.n104 10.6151
R1030 B.n108 B.n105 10.6151
R1031 B.n109 B.n108 10.6151
R1032 B.n112 B.n109 10.6151
R1033 B.n113 B.n112 10.6151
R1034 B.n116 B.n113 10.6151
R1035 B.n117 B.n116 10.6151
R1036 B.n120 B.n117 10.6151
R1037 B.n121 B.n120 10.6151
R1038 B.n124 B.n121 10.6151
R1039 B.n125 B.n124 10.6151
R1040 B.n128 B.n125 10.6151
R1041 B.n129 B.n128 10.6151
R1042 B.n132 B.n129 10.6151
R1043 B.n133 B.n132 10.6151
R1044 B.n136 B.n133 10.6151
R1045 B.n137 B.n136 10.6151
R1046 B.n140 B.n137 10.6151
R1047 B.n141 B.n140 10.6151
R1048 B.n144 B.n141 10.6151
R1049 B.n145 B.n144 10.6151
R1050 B.n148 B.n145 10.6151
R1051 B.n149 B.n148 10.6151
R1052 B.n152 B.n149 10.6151
R1053 B.n153 B.n152 10.6151
R1054 B.n156 B.n153 10.6151
R1055 B.n157 B.n156 10.6151
R1056 B.n160 B.n157 10.6151
R1057 B.n161 B.n160 10.6151
R1058 B.n164 B.n161 10.6151
R1059 B.n165 B.n164 10.6151
R1060 B.n168 B.n165 10.6151
R1061 B.n169 B.n168 10.6151
R1062 B.n172 B.n169 10.6151
R1063 B.n173 B.n172 10.6151
R1064 B.n176 B.n173 10.6151
R1065 B.n177 B.n176 10.6151
R1066 B.n180 B.n177 10.6151
R1067 B.n181 B.n180 10.6151
R1068 B.n184 B.n181 10.6151
R1069 B.n185 B.n184 10.6151
R1070 B.n188 B.n185 10.6151
R1071 B.n189 B.n188 10.6151
R1072 B.n192 B.n189 10.6151
R1073 B.n193 B.n192 10.6151
R1074 B.n196 B.n193 10.6151
R1075 B.n197 B.n196 10.6151
R1076 B.n200 B.n197 10.6151
R1077 B.n201 B.n200 10.6151
R1078 B.n204 B.n201 10.6151
R1079 B.n209 B.n206 10.6151
R1080 B.n210 B.n209 10.6151
R1081 B.n213 B.n210 10.6151
R1082 B.n214 B.n213 10.6151
R1083 B.n217 B.n214 10.6151
R1084 B.n218 B.n217 10.6151
R1085 B.n221 B.n218 10.6151
R1086 B.n222 B.n221 10.6151
R1087 B.n226 B.n225 10.6151
R1088 B.n229 B.n226 10.6151
R1089 B.n230 B.n229 10.6151
R1090 B.n233 B.n230 10.6151
R1091 B.n234 B.n233 10.6151
R1092 B.n237 B.n234 10.6151
R1093 B.n238 B.n237 10.6151
R1094 B.n241 B.n238 10.6151
R1095 B.n242 B.n241 10.6151
R1096 B.n245 B.n242 10.6151
R1097 B.n246 B.n245 10.6151
R1098 B.n249 B.n246 10.6151
R1099 B.n250 B.n249 10.6151
R1100 B.n253 B.n250 10.6151
R1101 B.n254 B.n253 10.6151
R1102 B.n257 B.n254 10.6151
R1103 B.n258 B.n257 10.6151
R1104 B.n261 B.n258 10.6151
R1105 B.n262 B.n261 10.6151
R1106 B.n265 B.n262 10.6151
R1107 B.n266 B.n265 10.6151
R1108 B.n269 B.n266 10.6151
R1109 B.n270 B.n269 10.6151
R1110 B.n273 B.n270 10.6151
R1111 B.n274 B.n273 10.6151
R1112 B.n277 B.n274 10.6151
R1113 B.n278 B.n277 10.6151
R1114 B.n281 B.n278 10.6151
R1115 B.n282 B.n281 10.6151
R1116 B.n285 B.n282 10.6151
R1117 B.n286 B.n285 10.6151
R1118 B.n289 B.n286 10.6151
R1119 B.n290 B.n289 10.6151
R1120 B.n293 B.n290 10.6151
R1121 B.n294 B.n293 10.6151
R1122 B.n297 B.n294 10.6151
R1123 B.n298 B.n297 10.6151
R1124 B.n301 B.n298 10.6151
R1125 B.n302 B.n301 10.6151
R1126 B.n305 B.n302 10.6151
R1127 B.n306 B.n305 10.6151
R1128 B.n309 B.n306 10.6151
R1129 B.n310 B.n309 10.6151
R1130 B.n313 B.n310 10.6151
R1131 B.n314 B.n313 10.6151
R1132 B.n317 B.n314 10.6151
R1133 B.n318 B.n317 10.6151
R1134 B.n321 B.n318 10.6151
R1135 B.n322 B.n321 10.6151
R1136 B.n325 B.n322 10.6151
R1137 B.n326 B.n325 10.6151
R1138 B.n737 B.n326 10.6151
R1139 B.n661 B.n358 10.6151
R1140 B.n662 B.n661 10.6151
R1141 B.n663 B.n662 10.6151
R1142 B.n663 B.n350 10.6151
R1143 B.n673 B.n350 10.6151
R1144 B.n674 B.n673 10.6151
R1145 B.n675 B.n674 10.6151
R1146 B.n675 B.n342 10.6151
R1147 B.n685 B.n342 10.6151
R1148 B.n686 B.n685 10.6151
R1149 B.n687 B.n686 10.6151
R1150 B.n687 B.n335 10.6151
R1151 B.n698 B.n335 10.6151
R1152 B.n699 B.n698 10.6151
R1153 B.n701 B.n699 10.6151
R1154 B.n701 B.n700 10.6151
R1155 B.n700 B.n327 10.6151
R1156 B.n712 B.n327 10.6151
R1157 B.n713 B.n712 10.6151
R1158 B.n714 B.n713 10.6151
R1159 B.n715 B.n714 10.6151
R1160 B.n717 B.n715 10.6151
R1161 B.n718 B.n717 10.6151
R1162 B.n719 B.n718 10.6151
R1163 B.n720 B.n719 10.6151
R1164 B.n722 B.n720 10.6151
R1165 B.n723 B.n722 10.6151
R1166 B.n724 B.n723 10.6151
R1167 B.n725 B.n724 10.6151
R1168 B.n727 B.n725 10.6151
R1169 B.n728 B.n727 10.6151
R1170 B.n729 B.n728 10.6151
R1171 B.n730 B.n729 10.6151
R1172 B.n732 B.n730 10.6151
R1173 B.n733 B.n732 10.6151
R1174 B.n734 B.n733 10.6151
R1175 B.n735 B.n734 10.6151
R1176 B.n736 B.n735 10.6151
R1177 B.n655 B.n362 10.6151
R1178 B.n650 B.n362 10.6151
R1179 B.n650 B.n649 10.6151
R1180 B.n649 B.n648 10.6151
R1181 B.n648 B.n645 10.6151
R1182 B.n645 B.n644 10.6151
R1183 B.n644 B.n641 10.6151
R1184 B.n641 B.n640 10.6151
R1185 B.n640 B.n637 10.6151
R1186 B.n637 B.n636 10.6151
R1187 B.n636 B.n633 10.6151
R1188 B.n633 B.n632 10.6151
R1189 B.n632 B.n629 10.6151
R1190 B.n629 B.n628 10.6151
R1191 B.n628 B.n625 10.6151
R1192 B.n625 B.n624 10.6151
R1193 B.n624 B.n621 10.6151
R1194 B.n621 B.n620 10.6151
R1195 B.n620 B.n617 10.6151
R1196 B.n617 B.n616 10.6151
R1197 B.n616 B.n613 10.6151
R1198 B.n613 B.n612 10.6151
R1199 B.n612 B.n609 10.6151
R1200 B.n609 B.n608 10.6151
R1201 B.n608 B.n605 10.6151
R1202 B.n605 B.n604 10.6151
R1203 B.n604 B.n601 10.6151
R1204 B.n601 B.n600 10.6151
R1205 B.n600 B.n597 10.6151
R1206 B.n597 B.n596 10.6151
R1207 B.n596 B.n593 10.6151
R1208 B.n593 B.n592 10.6151
R1209 B.n592 B.n589 10.6151
R1210 B.n589 B.n588 10.6151
R1211 B.n588 B.n585 10.6151
R1212 B.n585 B.n584 10.6151
R1213 B.n584 B.n581 10.6151
R1214 B.n581 B.n580 10.6151
R1215 B.n580 B.n577 10.6151
R1216 B.n577 B.n576 10.6151
R1217 B.n576 B.n573 10.6151
R1218 B.n573 B.n572 10.6151
R1219 B.n572 B.n569 10.6151
R1220 B.n569 B.n568 10.6151
R1221 B.n568 B.n565 10.6151
R1222 B.n565 B.n564 10.6151
R1223 B.n564 B.n561 10.6151
R1224 B.n561 B.n560 10.6151
R1225 B.n560 B.n557 10.6151
R1226 B.n557 B.n556 10.6151
R1227 B.n556 B.n553 10.6151
R1228 B.n553 B.n552 10.6151
R1229 B.n549 B.n548 10.6151
R1230 B.n548 B.n545 10.6151
R1231 B.n545 B.n544 10.6151
R1232 B.n544 B.n541 10.6151
R1233 B.n541 B.n540 10.6151
R1234 B.n540 B.n537 10.6151
R1235 B.n537 B.n536 10.6151
R1236 B.n536 B.n533 10.6151
R1237 B.n531 B.n528 10.6151
R1238 B.n528 B.n527 10.6151
R1239 B.n527 B.n524 10.6151
R1240 B.n524 B.n523 10.6151
R1241 B.n523 B.n520 10.6151
R1242 B.n520 B.n519 10.6151
R1243 B.n519 B.n516 10.6151
R1244 B.n516 B.n515 10.6151
R1245 B.n515 B.n512 10.6151
R1246 B.n512 B.n511 10.6151
R1247 B.n511 B.n508 10.6151
R1248 B.n508 B.n507 10.6151
R1249 B.n507 B.n504 10.6151
R1250 B.n504 B.n503 10.6151
R1251 B.n503 B.n500 10.6151
R1252 B.n500 B.n499 10.6151
R1253 B.n499 B.n496 10.6151
R1254 B.n496 B.n495 10.6151
R1255 B.n495 B.n492 10.6151
R1256 B.n492 B.n491 10.6151
R1257 B.n491 B.n488 10.6151
R1258 B.n488 B.n487 10.6151
R1259 B.n487 B.n484 10.6151
R1260 B.n484 B.n483 10.6151
R1261 B.n483 B.n480 10.6151
R1262 B.n480 B.n479 10.6151
R1263 B.n479 B.n476 10.6151
R1264 B.n476 B.n475 10.6151
R1265 B.n475 B.n472 10.6151
R1266 B.n472 B.n471 10.6151
R1267 B.n471 B.n468 10.6151
R1268 B.n468 B.n467 10.6151
R1269 B.n467 B.n464 10.6151
R1270 B.n464 B.n463 10.6151
R1271 B.n463 B.n460 10.6151
R1272 B.n460 B.n459 10.6151
R1273 B.n459 B.n456 10.6151
R1274 B.n456 B.n455 10.6151
R1275 B.n455 B.n452 10.6151
R1276 B.n452 B.n451 10.6151
R1277 B.n451 B.n448 10.6151
R1278 B.n448 B.n447 10.6151
R1279 B.n447 B.n444 10.6151
R1280 B.n444 B.n443 10.6151
R1281 B.n443 B.n440 10.6151
R1282 B.n440 B.n439 10.6151
R1283 B.n439 B.n436 10.6151
R1284 B.n436 B.n435 10.6151
R1285 B.n435 B.n432 10.6151
R1286 B.n432 B.n431 10.6151
R1287 B.n431 B.n428 10.6151
R1288 B.n428 B.n427 10.6151
R1289 B.n657 B.n656 10.6151
R1290 B.n657 B.n354 10.6151
R1291 B.n667 B.n354 10.6151
R1292 B.n668 B.n667 10.6151
R1293 B.n669 B.n668 10.6151
R1294 B.n669 B.n346 10.6151
R1295 B.n679 B.n346 10.6151
R1296 B.n680 B.n679 10.6151
R1297 B.n681 B.n680 10.6151
R1298 B.n681 B.n338 10.6151
R1299 B.n692 B.n338 10.6151
R1300 B.n693 B.n692 10.6151
R1301 B.n694 B.n693 10.6151
R1302 B.n694 B.n331 10.6151
R1303 B.n705 B.n331 10.6151
R1304 B.n706 B.n705 10.6151
R1305 B.n707 B.n706 10.6151
R1306 B.n707 B.n0 10.6151
R1307 B.n776 B.n1 10.6151
R1308 B.n776 B.n775 10.6151
R1309 B.n775 B.n774 10.6151
R1310 B.n774 B.n10 10.6151
R1311 B.n768 B.n10 10.6151
R1312 B.n768 B.n767 10.6151
R1313 B.n767 B.n766 10.6151
R1314 B.n766 B.n16 10.6151
R1315 B.n760 B.n16 10.6151
R1316 B.n760 B.n759 10.6151
R1317 B.n759 B.n758 10.6151
R1318 B.n758 B.n24 10.6151
R1319 B.n752 B.n24 10.6151
R1320 B.n752 B.n751 10.6151
R1321 B.n751 B.n750 10.6151
R1322 B.n750 B.n31 10.6151
R1323 B.n744 B.n31 10.6151
R1324 B.n744 B.n743 10.6151
R1325 B.n671 B.t12 7.8483
R1326 B.t5 B.n754 7.8483
R1327 B.n206 B.n205 6.5566
R1328 B.n222 B.n100 6.5566
R1329 B.n549 B.n423 6.5566
R1330 B.n533 B.n532 6.5566
R1331 B.n205 B.n204 4.05904
R1332 B.n225 B.n100 4.05904
R1333 B.n552 B.n423 4.05904
R1334 B.n532 B.n531 4.05904
R1335 B.n782 B.n0 2.81026
R1336 B.n782 B.n1 2.81026
R1337 B.n689 B.t3 0.523687
R1338 B.n18 B.t2 0.523687
R1339 VN.n0 VN.t0 491.894
R1340 VN.n1 VN.t1 491.894
R1341 VN.n0 VN.t3 491.844
R1342 VN.n1 VN.t2 491.844
R1343 VN VN.n1 89.0125
R1344 VN VN.n0 44.7132
R1345 VDD2.n2 VDD2.n0 101.838
R1346 VDD2.n2 VDD2.n1 61.3899
R1347 VDD2.n1 VDD2.t1 1.25764
R1348 VDD2.n1 VDD2.t2 1.25764
R1349 VDD2.n0 VDD2.t3 1.25764
R1350 VDD2.n0 VDD2.t0 1.25764
R1351 VDD2 VDD2.n2 0.0586897
C0 VDD2 VTAIL 7.77411f
C1 VDD1 VN 0.147263f
C2 VDD2 VDD1 0.610488f
C3 VDD1 VTAIL 7.73137f
C4 VN VP 5.64915f
C5 VDD2 VP 0.285304f
C6 VTAIL VP 4.00779f
C7 VDD2 VN 4.50616f
C8 VTAIL VN 3.99368f
C9 VDD1 VP 4.6439f
C10 VDD2 B 3.099456f
C11 VDD1 B 7.18947f
C12 VTAIL B 11.093533f
C13 VN B 8.849919f
C14 VP B 5.547014f
C15 VDD2.t3 B 0.343377f
C16 VDD2.t0 B 0.343377f
C17 VDD2.n0 B 3.85006f
C18 VDD2.t1 B 0.343377f
C19 VDD2.t2 B 0.343377f
C20 VDD2.n1 B 3.11133f
C21 VDD2.n2 B 3.86567f
C22 VN.t0 B 1.80426f
C23 VN.t3 B 1.80419f
C24 VN.n0 B 1.30222f
C25 VN.t1 B 1.80426f
C26 VN.t2 B 1.80419f
C27 VN.n1 B 2.35791f
C28 VTAIL.t0 B 2.18896f
C29 VTAIL.n0 B 0.26259f
C30 VTAIL.t4 B 2.18896f
C31 VTAIL.n1 B 0.286128f
C32 VTAIL.t5 B 2.18896f
C33 VTAIL.n2 B 1.21096f
C34 VTAIL.t3 B 2.18897f
C35 VTAIL.n3 B 1.21094f
C36 VTAIL.t1 B 2.18897f
C37 VTAIL.n4 B 0.286114f
C38 VTAIL.t7 B 2.18897f
C39 VTAIL.n5 B 0.286114f
C40 VTAIL.t6 B 2.18896f
C41 VTAIL.n6 B 1.21096f
C42 VTAIL.t2 B 2.18896f
C43 VTAIL.n7 B 1.18156f
C44 VDD1.t2 B 0.340556f
C45 VDD1.t1 B 0.340556f
C46 VDD1.n0 B 3.08608f
C47 VDD1.t0 B 0.340556f
C48 VDD1.t3 B 0.340556f
C49 VDD1.n1 B 3.84611f
C50 VP.n0 B 0.045105f
C51 VP.t1 B 1.8251f
C52 VP.t0 B 1.82517f
C53 VP.n1 B 2.36597f
C54 VP.n2 B 3.10951f
C55 VP.t2 B 1.79589f
C56 VP.n3 B 0.682528f
C57 VP.n4 B 0.010235f
C58 VP.t3 B 1.79589f
C59 VP.n5 B 0.682528f
C60 VP.n6 B 0.034955f
.ends

