* NGSPICE file created from diff_pair_sample_1264.ext - technology: sky130A

.subckt diff_pair_sample_1264 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=5.031 ps=26.58 w=12.9 l=2.73
X1 VTAIL.t5 VP.t0 VDD1.t5 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=2.1285 ps=13.23 w=12.9 l=2.73
X2 VDD2.t4 VN.t1 VTAIL.t9 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=2.1285 ps=13.23 w=12.9 l=2.73
X3 B.t11 B.t9 B.t10 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=0 ps=0 w=12.9 l=2.73
X4 B.t8 B.t6 B.t7 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=0 ps=0 w=12.9 l=2.73
X5 VTAIL.t2 VP.t1 VDD1.t4 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=2.1285 ps=13.23 w=12.9 l=2.73
X6 VTAIL.t7 VN.t2 VDD2.t3 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=2.1285 ps=13.23 w=12.9 l=2.73
X7 VDD2.t2 VN.t3 VTAIL.t10 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=5.031 ps=26.58 w=12.9 l=2.73
X8 B.t5 B.t3 B.t4 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=0 ps=0 w=12.9 l=2.73
X9 VDD1.t3 VP.t2 VTAIL.t1 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=5.031 ps=26.58 w=12.9 l=2.73
X10 VDD1.t2 VP.t3 VTAIL.t4 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=5.031 ps=26.58 w=12.9 l=2.73
X11 VDD1.t1 VP.t4 VTAIL.t0 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=2.1285 ps=13.23 w=12.9 l=2.73
X12 VTAIL.t6 VN.t4 VDD2.t1 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=2.1285 pd=13.23 as=2.1285 ps=13.23 w=12.9 l=2.73
X13 B.t2 B.t0 B.t1 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=0 ps=0 w=12.9 l=2.73
X14 VDD2.t0 VN.t5 VTAIL.t8 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=2.1285 ps=13.23 w=12.9 l=2.73
X15 VDD1.t0 VP.t5 VTAIL.t3 w_n3418_n3548# sky130_fd_pr__pfet_01v8 ad=5.031 pd=26.58 as=2.1285 ps=13.23 w=12.9 l=2.73
R0 VN.n29 VN.n16 161.3
R1 VN.n28 VN.n27 161.3
R2 VN.n26 VN.n17 161.3
R3 VN.n25 VN.n24 161.3
R4 VN.n23 VN.n18 161.3
R5 VN.n22 VN.n21 161.3
R6 VN.n13 VN.n0 161.3
R7 VN.n12 VN.n11 161.3
R8 VN.n10 VN.n1 161.3
R9 VN.n9 VN.n8 161.3
R10 VN.n7 VN.n2 161.3
R11 VN.n6 VN.n5 161.3
R12 VN.n4 VN.t5 147.101
R13 VN.n20 VN.t3 147.101
R14 VN.n3 VN.t2 113.879
R15 VN.n14 VN.t0 113.879
R16 VN.n19 VN.t4 113.879
R17 VN.n30 VN.t1 113.879
R18 VN.n15 VN.n14 107.684
R19 VN.n31 VN.n30 107.684
R20 VN VN.n31 50.089
R21 VN.n20 VN.n19 48.82
R22 VN.n4 VN.n3 48.82
R23 VN.n8 VN.n1 43.3318
R24 VN.n24 VN.n17 43.3318
R25 VN.n8 VN.n7 37.4894
R26 VN.n24 VN.n23 37.4894
R27 VN.n6 VN.n3 24.3439
R28 VN.n7 VN.n6 24.3439
R29 VN.n12 VN.n1 24.3439
R30 VN.n13 VN.n12 24.3439
R31 VN.n23 VN.n22 24.3439
R32 VN.n22 VN.n19 24.3439
R33 VN.n29 VN.n28 24.3439
R34 VN.n28 VN.n17 24.3439
R35 VN.n21 VN.n20 5.08087
R36 VN.n5 VN.n4 5.08087
R37 VN.n14 VN.n13 2.92171
R38 VN.n30 VN.n29 2.92171
R39 VN.n31 VN.n16 0.278398
R40 VN.n15 VN.n0 0.278398
R41 VN.n27 VN.n16 0.189894
R42 VN.n27 VN.n26 0.189894
R43 VN.n26 VN.n25 0.189894
R44 VN.n25 VN.n18 0.189894
R45 VN.n21 VN.n18 0.189894
R46 VN.n5 VN.n2 0.189894
R47 VN.n9 VN.n2 0.189894
R48 VN.n10 VN.n9 0.189894
R49 VN.n11 VN.n10 0.189894
R50 VN.n11 VN.n0 0.189894
R51 VN VN.n15 0.153422
R52 VTAIL.n282 VTAIL.n218 756.745
R53 VTAIL.n66 VTAIL.n2 756.745
R54 VTAIL.n212 VTAIL.n148 756.745
R55 VTAIL.n140 VTAIL.n76 756.745
R56 VTAIL.n241 VTAIL.n240 585
R57 VTAIL.n238 VTAIL.n237 585
R58 VTAIL.n247 VTAIL.n246 585
R59 VTAIL.n249 VTAIL.n248 585
R60 VTAIL.n234 VTAIL.n233 585
R61 VTAIL.n255 VTAIL.n254 585
R62 VTAIL.n258 VTAIL.n257 585
R63 VTAIL.n256 VTAIL.n230 585
R64 VTAIL.n263 VTAIL.n229 585
R65 VTAIL.n265 VTAIL.n264 585
R66 VTAIL.n267 VTAIL.n266 585
R67 VTAIL.n226 VTAIL.n225 585
R68 VTAIL.n273 VTAIL.n272 585
R69 VTAIL.n275 VTAIL.n274 585
R70 VTAIL.n222 VTAIL.n221 585
R71 VTAIL.n281 VTAIL.n280 585
R72 VTAIL.n283 VTAIL.n282 585
R73 VTAIL.n25 VTAIL.n24 585
R74 VTAIL.n22 VTAIL.n21 585
R75 VTAIL.n31 VTAIL.n30 585
R76 VTAIL.n33 VTAIL.n32 585
R77 VTAIL.n18 VTAIL.n17 585
R78 VTAIL.n39 VTAIL.n38 585
R79 VTAIL.n42 VTAIL.n41 585
R80 VTAIL.n40 VTAIL.n14 585
R81 VTAIL.n47 VTAIL.n13 585
R82 VTAIL.n49 VTAIL.n48 585
R83 VTAIL.n51 VTAIL.n50 585
R84 VTAIL.n10 VTAIL.n9 585
R85 VTAIL.n57 VTAIL.n56 585
R86 VTAIL.n59 VTAIL.n58 585
R87 VTAIL.n6 VTAIL.n5 585
R88 VTAIL.n65 VTAIL.n64 585
R89 VTAIL.n67 VTAIL.n66 585
R90 VTAIL.n213 VTAIL.n212 585
R91 VTAIL.n211 VTAIL.n210 585
R92 VTAIL.n152 VTAIL.n151 585
R93 VTAIL.n205 VTAIL.n204 585
R94 VTAIL.n203 VTAIL.n202 585
R95 VTAIL.n156 VTAIL.n155 585
R96 VTAIL.n197 VTAIL.n196 585
R97 VTAIL.n195 VTAIL.n194 585
R98 VTAIL.n193 VTAIL.n159 585
R99 VTAIL.n163 VTAIL.n160 585
R100 VTAIL.n188 VTAIL.n187 585
R101 VTAIL.n186 VTAIL.n185 585
R102 VTAIL.n165 VTAIL.n164 585
R103 VTAIL.n180 VTAIL.n179 585
R104 VTAIL.n178 VTAIL.n177 585
R105 VTAIL.n169 VTAIL.n168 585
R106 VTAIL.n172 VTAIL.n171 585
R107 VTAIL.n141 VTAIL.n140 585
R108 VTAIL.n139 VTAIL.n138 585
R109 VTAIL.n80 VTAIL.n79 585
R110 VTAIL.n133 VTAIL.n132 585
R111 VTAIL.n131 VTAIL.n130 585
R112 VTAIL.n84 VTAIL.n83 585
R113 VTAIL.n125 VTAIL.n124 585
R114 VTAIL.n123 VTAIL.n122 585
R115 VTAIL.n121 VTAIL.n87 585
R116 VTAIL.n91 VTAIL.n88 585
R117 VTAIL.n116 VTAIL.n115 585
R118 VTAIL.n114 VTAIL.n113 585
R119 VTAIL.n93 VTAIL.n92 585
R120 VTAIL.n108 VTAIL.n107 585
R121 VTAIL.n106 VTAIL.n105 585
R122 VTAIL.n97 VTAIL.n96 585
R123 VTAIL.n100 VTAIL.n99 585
R124 VTAIL.t11 VTAIL.n239 329.036
R125 VTAIL.t4 VTAIL.n23 329.036
R126 VTAIL.t1 VTAIL.n170 329.036
R127 VTAIL.t10 VTAIL.n98 329.036
R128 VTAIL.n240 VTAIL.n237 171.744
R129 VTAIL.n247 VTAIL.n237 171.744
R130 VTAIL.n248 VTAIL.n247 171.744
R131 VTAIL.n248 VTAIL.n233 171.744
R132 VTAIL.n255 VTAIL.n233 171.744
R133 VTAIL.n257 VTAIL.n255 171.744
R134 VTAIL.n257 VTAIL.n256 171.744
R135 VTAIL.n256 VTAIL.n229 171.744
R136 VTAIL.n265 VTAIL.n229 171.744
R137 VTAIL.n266 VTAIL.n265 171.744
R138 VTAIL.n266 VTAIL.n225 171.744
R139 VTAIL.n273 VTAIL.n225 171.744
R140 VTAIL.n274 VTAIL.n273 171.744
R141 VTAIL.n274 VTAIL.n221 171.744
R142 VTAIL.n281 VTAIL.n221 171.744
R143 VTAIL.n282 VTAIL.n281 171.744
R144 VTAIL.n24 VTAIL.n21 171.744
R145 VTAIL.n31 VTAIL.n21 171.744
R146 VTAIL.n32 VTAIL.n31 171.744
R147 VTAIL.n32 VTAIL.n17 171.744
R148 VTAIL.n39 VTAIL.n17 171.744
R149 VTAIL.n41 VTAIL.n39 171.744
R150 VTAIL.n41 VTAIL.n40 171.744
R151 VTAIL.n40 VTAIL.n13 171.744
R152 VTAIL.n49 VTAIL.n13 171.744
R153 VTAIL.n50 VTAIL.n49 171.744
R154 VTAIL.n50 VTAIL.n9 171.744
R155 VTAIL.n57 VTAIL.n9 171.744
R156 VTAIL.n58 VTAIL.n57 171.744
R157 VTAIL.n58 VTAIL.n5 171.744
R158 VTAIL.n65 VTAIL.n5 171.744
R159 VTAIL.n66 VTAIL.n65 171.744
R160 VTAIL.n212 VTAIL.n211 171.744
R161 VTAIL.n211 VTAIL.n151 171.744
R162 VTAIL.n204 VTAIL.n151 171.744
R163 VTAIL.n204 VTAIL.n203 171.744
R164 VTAIL.n203 VTAIL.n155 171.744
R165 VTAIL.n196 VTAIL.n155 171.744
R166 VTAIL.n196 VTAIL.n195 171.744
R167 VTAIL.n195 VTAIL.n159 171.744
R168 VTAIL.n163 VTAIL.n159 171.744
R169 VTAIL.n187 VTAIL.n163 171.744
R170 VTAIL.n187 VTAIL.n186 171.744
R171 VTAIL.n186 VTAIL.n164 171.744
R172 VTAIL.n179 VTAIL.n164 171.744
R173 VTAIL.n179 VTAIL.n178 171.744
R174 VTAIL.n178 VTAIL.n168 171.744
R175 VTAIL.n171 VTAIL.n168 171.744
R176 VTAIL.n140 VTAIL.n139 171.744
R177 VTAIL.n139 VTAIL.n79 171.744
R178 VTAIL.n132 VTAIL.n79 171.744
R179 VTAIL.n132 VTAIL.n131 171.744
R180 VTAIL.n131 VTAIL.n83 171.744
R181 VTAIL.n124 VTAIL.n83 171.744
R182 VTAIL.n124 VTAIL.n123 171.744
R183 VTAIL.n123 VTAIL.n87 171.744
R184 VTAIL.n91 VTAIL.n87 171.744
R185 VTAIL.n115 VTAIL.n91 171.744
R186 VTAIL.n115 VTAIL.n114 171.744
R187 VTAIL.n114 VTAIL.n92 171.744
R188 VTAIL.n107 VTAIL.n92 171.744
R189 VTAIL.n107 VTAIL.n106 171.744
R190 VTAIL.n106 VTAIL.n96 171.744
R191 VTAIL.n99 VTAIL.n96 171.744
R192 VTAIL.n240 VTAIL.t11 85.8723
R193 VTAIL.n24 VTAIL.t4 85.8723
R194 VTAIL.n171 VTAIL.t1 85.8723
R195 VTAIL.n99 VTAIL.t10 85.8723
R196 VTAIL.n1 VTAIL.n0 57.4962
R197 VTAIL.n73 VTAIL.n72 57.4962
R198 VTAIL.n147 VTAIL.n146 57.4962
R199 VTAIL.n75 VTAIL.n74 57.4962
R200 VTAIL.n287 VTAIL.n286 33.349
R201 VTAIL.n71 VTAIL.n70 33.349
R202 VTAIL.n217 VTAIL.n216 33.349
R203 VTAIL.n145 VTAIL.n144 33.349
R204 VTAIL.n75 VTAIL.n73 28.7634
R205 VTAIL.n287 VTAIL.n217 26.1255
R206 VTAIL.n264 VTAIL.n263 13.1884
R207 VTAIL.n48 VTAIL.n47 13.1884
R208 VTAIL.n194 VTAIL.n193 13.1884
R209 VTAIL.n122 VTAIL.n121 13.1884
R210 VTAIL.n262 VTAIL.n230 12.8005
R211 VTAIL.n267 VTAIL.n228 12.8005
R212 VTAIL.n46 VTAIL.n14 12.8005
R213 VTAIL.n51 VTAIL.n12 12.8005
R214 VTAIL.n197 VTAIL.n158 12.8005
R215 VTAIL.n192 VTAIL.n160 12.8005
R216 VTAIL.n125 VTAIL.n86 12.8005
R217 VTAIL.n120 VTAIL.n88 12.8005
R218 VTAIL.n259 VTAIL.n258 12.0247
R219 VTAIL.n268 VTAIL.n226 12.0247
R220 VTAIL.n43 VTAIL.n42 12.0247
R221 VTAIL.n52 VTAIL.n10 12.0247
R222 VTAIL.n198 VTAIL.n156 12.0247
R223 VTAIL.n189 VTAIL.n188 12.0247
R224 VTAIL.n126 VTAIL.n84 12.0247
R225 VTAIL.n117 VTAIL.n116 12.0247
R226 VTAIL.n254 VTAIL.n232 11.249
R227 VTAIL.n272 VTAIL.n271 11.249
R228 VTAIL.n38 VTAIL.n16 11.249
R229 VTAIL.n56 VTAIL.n55 11.249
R230 VTAIL.n202 VTAIL.n201 11.249
R231 VTAIL.n185 VTAIL.n162 11.249
R232 VTAIL.n130 VTAIL.n129 11.249
R233 VTAIL.n113 VTAIL.n90 11.249
R234 VTAIL.n241 VTAIL.n239 10.7239
R235 VTAIL.n25 VTAIL.n23 10.7239
R236 VTAIL.n172 VTAIL.n170 10.7239
R237 VTAIL.n100 VTAIL.n98 10.7239
R238 VTAIL.n253 VTAIL.n234 10.4732
R239 VTAIL.n275 VTAIL.n224 10.4732
R240 VTAIL.n37 VTAIL.n18 10.4732
R241 VTAIL.n59 VTAIL.n8 10.4732
R242 VTAIL.n205 VTAIL.n154 10.4732
R243 VTAIL.n184 VTAIL.n165 10.4732
R244 VTAIL.n133 VTAIL.n82 10.4732
R245 VTAIL.n112 VTAIL.n93 10.4732
R246 VTAIL.n250 VTAIL.n249 9.69747
R247 VTAIL.n276 VTAIL.n222 9.69747
R248 VTAIL.n34 VTAIL.n33 9.69747
R249 VTAIL.n60 VTAIL.n6 9.69747
R250 VTAIL.n206 VTAIL.n152 9.69747
R251 VTAIL.n181 VTAIL.n180 9.69747
R252 VTAIL.n134 VTAIL.n80 9.69747
R253 VTAIL.n109 VTAIL.n108 9.69747
R254 VTAIL.n286 VTAIL.n285 9.45567
R255 VTAIL.n70 VTAIL.n69 9.45567
R256 VTAIL.n216 VTAIL.n215 9.45567
R257 VTAIL.n144 VTAIL.n143 9.45567
R258 VTAIL.n220 VTAIL.n219 9.3005
R259 VTAIL.n279 VTAIL.n278 9.3005
R260 VTAIL.n277 VTAIL.n276 9.3005
R261 VTAIL.n224 VTAIL.n223 9.3005
R262 VTAIL.n271 VTAIL.n270 9.3005
R263 VTAIL.n269 VTAIL.n268 9.3005
R264 VTAIL.n228 VTAIL.n227 9.3005
R265 VTAIL.n243 VTAIL.n242 9.3005
R266 VTAIL.n245 VTAIL.n244 9.3005
R267 VTAIL.n236 VTAIL.n235 9.3005
R268 VTAIL.n251 VTAIL.n250 9.3005
R269 VTAIL.n253 VTAIL.n252 9.3005
R270 VTAIL.n232 VTAIL.n231 9.3005
R271 VTAIL.n260 VTAIL.n259 9.3005
R272 VTAIL.n262 VTAIL.n261 9.3005
R273 VTAIL.n285 VTAIL.n284 9.3005
R274 VTAIL.n4 VTAIL.n3 9.3005
R275 VTAIL.n63 VTAIL.n62 9.3005
R276 VTAIL.n61 VTAIL.n60 9.3005
R277 VTAIL.n8 VTAIL.n7 9.3005
R278 VTAIL.n55 VTAIL.n54 9.3005
R279 VTAIL.n53 VTAIL.n52 9.3005
R280 VTAIL.n12 VTAIL.n11 9.3005
R281 VTAIL.n27 VTAIL.n26 9.3005
R282 VTAIL.n29 VTAIL.n28 9.3005
R283 VTAIL.n20 VTAIL.n19 9.3005
R284 VTAIL.n35 VTAIL.n34 9.3005
R285 VTAIL.n37 VTAIL.n36 9.3005
R286 VTAIL.n16 VTAIL.n15 9.3005
R287 VTAIL.n44 VTAIL.n43 9.3005
R288 VTAIL.n46 VTAIL.n45 9.3005
R289 VTAIL.n69 VTAIL.n68 9.3005
R290 VTAIL.n174 VTAIL.n173 9.3005
R291 VTAIL.n176 VTAIL.n175 9.3005
R292 VTAIL.n167 VTAIL.n166 9.3005
R293 VTAIL.n182 VTAIL.n181 9.3005
R294 VTAIL.n184 VTAIL.n183 9.3005
R295 VTAIL.n162 VTAIL.n161 9.3005
R296 VTAIL.n190 VTAIL.n189 9.3005
R297 VTAIL.n192 VTAIL.n191 9.3005
R298 VTAIL.n215 VTAIL.n214 9.3005
R299 VTAIL.n150 VTAIL.n149 9.3005
R300 VTAIL.n209 VTAIL.n208 9.3005
R301 VTAIL.n207 VTAIL.n206 9.3005
R302 VTAIL.n154 VTAIL.n153 9.3005
R303 VTAIL.n201 VTAIL.n200 9.3005
R304 VTAIL.n199 VTAIL.n198 9.3005
R305 VTAIL.n158 VTAIL.n157 9.3005
R306 VTAIL.n102 VTAIL.n101 9.3005
R307 VTAIL.n104 VTAIL.n103 9.3005
R308 VTAIL.n95 VTAIL.n94 9.3005
R309 VTAIL.n110 VTAIL.n109 9.3005
R310 VTAIL.n112 VTAIL.n111 9.3005
R311 VTAIL.n90 VTAIL.n89 9.3005
R312 VTAIL.n118 VTAIL.n117 9.3005
R313 VTAIL.n120 VTAIL.n119 9.3005
R314 VTAIL.n143 VTAIL.n142 9.3005
R315 VTAIL.n78 VTAIL.n77 9.3005
R316 VTAIL.n137 VTAIL.n136 9.3005
R317 VTAIL.n135 VTAIL.n134 9.3005
R318 VTAIL.n82 VTAIL.n81 9.3005
R319 VTAIL.n129 VTAIL.n128 9.3005
R320 VTAIL.n127 VTAIL.n126 9.3005
R321 VTAIL.n86 VTAIL.n85 9.3005
R322 VTAIL.n246 VTAIL.n236 8.92171
R323 VTAIL.n280 VTAIL.n279 8.92171
R324 VTAIL.n30 VTAIL.n20 8.92171
R325 VTAIL.n64 VTAIL.n63 8.92171
R326 VTAIL.n210 VTAIL.n209 8.92171
R327 VTAIL.n177 VTAIL.n167 8.92171
R328 VTAIL.n138 VTAIL.n137 8.92171
R329 VTAIL.n105 VTAIL.n95 8.92171
R330 VTAIL.n245 VTAIL.n238 8.14595
R331 VTAIL.n283 VTAIL.n220 8.14595
R332 VTAIL.n29 VTAIL.n22 8.14595
R333 VTAIL.n67 VTAIL.n4 8.14595
R334 VTAIL.n213 VTAIL.n150 8.14595
R335 VTAIL.n176 VTAIL.n169 8.14595
R336 VTAIL.n141 VTAIL.n78 8.14595
R337 VTAIL.n104 VTAIL.n97 8.14595
R338 VTAIL.n242 VTAIL.n241 7.3702
R339 VTAIL.n284 VTAIL.n218 7.3702
R340 VTAIL.n26 VTAIL.n25 7.3702
R341 VTAIL.n68 VTAIL.n2 7.3702
R342 VTAIL.n214 VTAIL.n148 7.3702
R343 VTAIL.n173 VTAIL.n172 7.3702
R344 VTAIL.n142 VTAIL.n76 7.3702
R345 VTAIL.n101 VTAIL.n100 7.3702
R346 VTAIL.n286 VTAIL.n218 6.59444
R347 VTAIL.n70 VTAIL.n2 6.59444
R348 VTAIL.n216 VTAIL.n148 6.59444
R349 VTAIL.n144 VTAIL.n76 6.59444
R350 VTAIL.n242 VTAIL.n238 5.81868
R351 VTAIL.n284 VTAIL.n283 5.81868
R352 VTAIL.n26 VTAIL.n22 5.81868
R353 VTAIL.n68 VTAIL.n67 5.81868
R354 VTAIL.n214 VTAIL.n213 5.81868
R355 VTAIL.n173 VTAIL.n169 5.81868
R356 VTAIL.n142 VTAIL.n141 5.81868
R357 VTAIL.n101 VTAIL.n97 5.81868
R358 VTAIL.n246 VTAIL.n245 5.04292
R359 VTAIL.n280 VTAIL.n220 5.04292
R360 VTAIL.n30 VTAIL.n29 5.04292
R361 VTAIL.n64 VTAIL.n4 5.04292
R362 VTAIL.n210 VTAIL.n150 5.04292
R363 VTAIL.n177 VTAIL.n176 5.04292
R364 VTAIL.n138 VTAIL.n78 5.04292
R365 VTAIL.n105 VTAIL.n104 5.04292
R366 VTAIL.n249 VTAIL.n236 4.26717
R367 VTAIL.n279 VTAIL.n222 4.26717
R368 VTAIL.n33 VTAIL.n20 4.26717
R369 VTAIL.n63 VTAIL.n6 4.26717
R370 VTAIL.n209 VTAIL.n152 4.26717
R371 VTAIL.n180 VTAIL.n167 4.26717
R372 VTAIL.n137 VTAIL.n80 4.26717
R373 VTAIL.n108 VTAIL.n95 4.26717
R374 VTAIL.n250 VTAIL.n234 3.49141
R375 VTAIL.n276 VTAIL.n275 3.49141
R376 VTAIL.n34 VTAIL.n18 3.49141
R377 VTAIL.n60 VTAIL.n59 3.49141
R378 VTAIL.n206 VTAIL.n205 3.49141
R379 VTAIL.n181 VTAIL.n165 3.49141
R380 VTAIL.n134 VTAIL.n133 3.49141
R381 VTAIL.n109 VTAIL.n93 3.49141
R382 VTAIL.n254 VTAIL.n253 2.71565
R383 VTAIL.n272 VTAIL.n224 2.71565
R384 VTAIL.n38 VTAIL.n37 2.71565
R385 VTAIL.n56 VTAIL.n8 2.71565
R386 VTAIL.n202 VTAIL.n154 2.71565
R387 VTAIL.n185 VTAIL.n184 2.71565
R388 VTAIL.n130 VTAIL.n82 2.71565
R389 VTAIL.n113 VTAIL.n112 2.71565
R390 VTAIL.n145 VTAIL.n75 2.63843
R391 VTAIL.n217 VTAIL.n147 2.63843
R392 VTAIL.n73 VTAIL.n71 2.63843
R393 VTAIL.n0 VTAIL.t8 2.52027
R394 VTAIL.n0 VTAIL.t7 2.52027
R395 VTAIL.n72 VTAIL.t0 2.52027
R396 VTAIL.n72 VTAIL.t2 2.52027
R397 VTAIL.n146 VTAIL.t3 2.52027
R398 VTAIL.n146 VTAIL.t5 2.52027
R399 VTAIL.n74 VTAIL.t9 2.52027
R400 VTAIL.n74 VTAIL.t6 2.52027
R401 VTAIL.n243 VTAIL.n239 2.41282
R402 VTAIL.n27 VTAIL.n23 2.41282
R403 VTAIL.n174 VTAIL.n170 2.41282
R404 VTAIL.n102 VTAIL.n98 2.41282
R405 VTAIL.n258 VTAIL.n232 1.93989
R406 VTAIL.n271 VTAIL.n226 1.93989
R407 VTAIL.n42 VTAIL.n16 1.93989
R408 VTAIL.n55 VTAIL.n10 1.93989
R409 VTAIL.n201 VTAIL.n156 1.93989
R410 VTAIL.n188 VTAIL.n162 1.93989
R411 VTAIL.n129 VTAIL.n84 1.93989
R412 VTAIL.n116 VTAIL.n90 1.93989
R413 VTAIL VTAIL.n287 1.92076
R414 VTAIL.n147 VTAIL.n145 1.78929
R415 VTAIL.n71 VTAIL.n1 1.78929
R416 VTAIL.n259 VTAIL.n230 1.16414
R417 VTAIL.n268 VTAIL.n267 1.16414
R418 VTAIL.n43 VTAIL.n14 1.16414
R419 VTAIL.n52 VTAIL.n51 1.16414
R420 VTAIL.n198 VTAIL.n197 1.16414
R421 VTAIL.n189 VTAIL.n160 1.16414
R422 VTAIL.n126 VTAIL.n125 1.16414
R423 VTAIL.n117 VTAIL.n88 1.16414
R424 VTAIL VTAIL.n1 0.718172
R425 VTAIL.n263 VTAIL.n262 0.388379
R426 VTAIL.n264 VTAIL.n228 0.388379
R427 VTAIL.n47 VTAIL.n46 0.388379
R428 VTAIL.n48 VTAIL.n12 0.388379
R429 VTAIL.n194 VTAIL.n158 0.388379
R430 VTAIL.n193 VTAIL.n192 0.388379
R431 VTAIL.n122 VTAIL.n86 0.388379
R432 VTAIL.n121 VTAIL.n120 0.388379
R433 VTAIL.n244 VTAIL.n243 0.155672
R434 VTAIL.n244 VTAIL.n235 0.155672
R435 VTAIL.n251 VTAIL.n235 0.155672
R436 VTAIL.n252 VTAIL.n251 0.155672
R437 VTAIL.n252 VTAIL.n231 0.155672
R438 VTAIL.n260 VTAIL.n231 0.155672
R439 VTAIL.n261 VTAIL.n260 0.155672
R440 VTAIL.n261 VTAIL.n227 0.155672
R441 VTAIL.n269 VTAIL.n227 0.155672
R442 VTAIL.n270 VTAIL.n269 0.155672
R443 VTAIL.n270 VTAIL.n223 0.155672
R444 VTAIL.n277 VTAIL.n223 0.155672
R445 VTAIL.n278 VTAIL.n277 0.155672
R446 VTAIL.n278 VTAIL.n219 0.155672
R447 VTAIL.n285 VTAIL.n219 0.155672
R448 VTAIL.n28 VTAIL.n27 0.155672
R449 VTAIL.n28 VTAIL.n19 0.155672
R450 VTAIL.n35 VTAIL.n19 0.155672
R451 VTAIL.n36 VTAIL.n35 0.155672
R452 VTAIL.n36 VTAIL.n15 0.155672
R453 VTAIL.n44 VTAIL.n15 0.155672
R454 VTAIL.n45 VTAIL.n44 0.155672
R455 VTAIL.n45 VTAIL.n11 0.155672
R456 VTAIL.n53 VTAIL.n11 0.155672
R457 VTAIL.n54 VTAIL.n53 0.155672
R458 VTAIL.n54 VTAIL.n7 0.155672
R459 VTAIL.n61 VTAIL.n7 0.155672
R460 VTAIL.n62 VTAIL.n61 0.155672
R461 VTAIL.n62 VTAIL.n3 0.155672
R462 VTAIL.n69 VTAIL.n3 0.155672
R463 VTAIL.n215 VTAIL.n149 0.155672
R464 VTAIL.n208 VTAIL.n149 0.155672
R465 VTAIL.n208 VTAIL.n207 0.155672
R466 VTAIL.n207 VTAIL.n153 0.155672
R467 VTAIL.n200 VTAIL.n153 0.155672
R468 VTAIL.n200 VTAIL.n199 0.155672
R469 VTAIL.n199 VTAIL.n157 0.155672
R470 VTAIL.n191 VTAIL.n157 0.155672
R471 VTAIL.n191 VTAIL.n190 0.155672
R472 VTAIL.n190 VTAIL.n161 0.155672
R473 VTAIL.n183 VTAIL.n161 0.155672
R474 VTAIL.n183 VTAIL.n182 0.155672
R475 VTAIL.n182 VTAIL.n166 0.155672
R476 VTAIL.n175 VTAIL.n166 0.155672
R477 VTAIL.n175 VTAIL.n174 0.155672
R478 VTAIL.n143 VTAIL.n77 0.155672
R479 VTAIL.n136 VTAIL.n77 0.155672
R480 VTAIL.n136 VTAIL.n135 0.155672
R481 VTAIL.n135 VTAIL.n81 0.155672
R482 VTAIL.n128 VTAIL.n81 0.155672
R483 VTAIL.n128 VTAIL.n127 0.155672
R484 VTAIL.n127 VTAIL.n85 0.155672
R485 VTAIL.n119 VTAIL.n85 0.155672
R486 VTAIL.n119 VTAIL.n118 0.155672
R487 VTAIL.n118 VTAIL.n89 0.155672
R488 VTAIL.n111 VTAIL.n89 0.155672
R489 VTAIL.n111 VTAIL.n110 0.155672
R490 VTAIL.n110 VTAIL.n94 0.155672
R491 VTAIL.n103 VTAIL.n94 0.155672
R492 VTAIL.n103 VTAIL.n102 0.155672
R493 VDD2.n135 VDD2.n71 756.745
R494 VDD2.n64 VDD2.n0 756.745
R495 VDD2.n136 VDD2.n135 585
R496 VDD2.n134 VDD2.n133 585
R497 VDD2.n75 VDD2.n74 585
R498 VDD2.n128 VDD2.n127 585
R499 VDD2.n126 VDD2.n125 585
R500 VDD2.n79 VDD2.n78 585
R501 VDD2.n120 VDD2.n119 585
R502 VDD2.n118 VDD2.n117 585
R503 VDD2.n116 VDD2.n82 585
R504 VDD2.n86 VDD2.n83 585
R505 VDD2.n111 VDD2.n110 585
R506 VDD2.n109 VDD2.n108 585
R507 VDD2.n88 VDD2.n87 585
R508 VDD2.n103 VDD2.n102 585
R509 VDD2.n101 VDD2.n100 585
R510 VDD2.n92 VDD2.n91 585
R511 VDD2.n95 VDD2.n94 585
R512 VDD2.n23 VDD2.n22 585
R513 VDD2.n20 VDD2.n19 585
R514 VDD2.n29 VDD2.n28 585
R515 VDD2.n31 VDD2.n30 585
R516 VDD2.n16 VDD2.n15 585
R517 VDD2.n37 VDD2.n36 585
R518 VDD2.n40 VDD2.n39 585
R519 VDD2.n38 VDD2.n12 585
R520 VDD2.n45 VDD2.n11 585
R521 VDD2.n47 VDD2.n46 585
R522 VDD2.n49 VDD2.n48 585
R523 VDD2.n8 VDD2.n7 585
R524 VDD2.n55 VDD2.n54 585
R525 VDD2.n57 VDD2.n56 585
R526 VDD2.n4 VDD2.n3 585
R527 VDD2.n63 VDD2.n62 585
R528 VDD2.n65 VDD2.n64 585
R529 VDD2.t0 VDD2.n21 329.036
R530 VDD2.t4 VDD2.n93 329.036
R531 VDD2.n135 VDD2.n134 171.744
R532 VDD2.n134 VDD2.n74 171.744
R533 VDD2.n127 VDD2.n74 171.744
R534 VDD2.n127 VDD2.n126 171.744
R535 VDD2.n126 VDD2.n78 171.744
R536 VDD2.n119 VDD2.n78 171.744
R537 VDD2.n119 VDD2.n118 171.744
R538 VDD2.n118 VDD2.n82 171.744
R539 VDD2.n86 VDD2.n82 171.744
R540 VDD2.n110 VDD2.n86 171.744
R541 VDD2.n110 VDD2.n109 171.744
R542 VDD2.n109 VDD2.n87 171.744
R543 VDD2.n102 VDD2.n87 171.744
R544 VDD2.n102 VDD2.n101 171.744
R545 VDD2.n101 VDD2.n91 171.744
R546 VDD2.n94 VDD2.n91 171.744
R547 VDD2.n22 VDD2.n19 171.744
R548 VDD2.n29 VDD2.n19 171.744
R549 VDD2.n30 VDD2.n29 171.744
R550 VDD2.n30 VDD2.n15 171.744
R551 VDD2.n37 VDD2.n15 171.744
R552 VDD2.n39 VDD2.n37 171.744
R553 VDD2.n39 VDD2.n38 171.744
R554 VDD2.n38 VDD2.n11 171.744
R555 VDD2.n47 VDD2.n11 171.744
R556 VDD2.n48 VDD2.n47 171.744
R557 VDD2.n48 VDD2.n7 171.744
R558 VDD2.n55 VDD2.n7 171.744
R559 VDD2.n56 VDD2.n55 171.744
R560 VDD2.n56 VDD2.n3 171.744
R561 VDD2.n63 VDD2.n3 171.744
R562 VDD2.n64 VDD2.n63 171.744
R563 VDD2.n94 VDD2.t4 85.8723
R564 VDD2.n22 VDD2.t0 85.8723
R565 VDD2.n70 VDD2.n69 74.7791
R566 VDD2 VDD2.n141 74.7761
R567 VDD2.n70 VDD2.n68 51.9509
R568 VDD2.n140 VDD2.n139 50.0278
R569 VDD2.n140 VDD2.n70 43.4093
R570 VDD2.n117 VDD2.n116 13.1884
R571 VDD2.n46 VDD2.n45 13.1884
R572 VDD2.n120 VDD2.n81 12.8005
R573 VDD2.n115 VDD2.n83 12.8005
R574 VDD2.n44 VDD2.n12 12.8005
R575 VDD2.n49 VDD2.n10 12.8005
R576 VDD2.n121 VDD2.n79 12.0247
R577 VDD2.n112 VDD2.n111 12.0247
R578 VDD2.n41 VDD2.n40 12.0247
R579 VDD2.n50 VDD2.n8 12.0247
R580 VDD2.n125 VDD2.n124 11.249
R581 VDD2.n108 VDD2.n85 11.249
R582 VDD2.n36 VDD2.n14 11.249
R583 VDD2.n54 VDD2.n53 11.249
R584 VDD2.n95 VDD2.n93 10.7239
R585 VDD2.n23 VDD2.n21 10.7239
R586 VDD2.n128 VDD2.n77 10.4732
R587 VDD2.n107 VDD2.n88 10.4732
R588 VDD2.n35 VDD2.n16 10.4732
R589 VDD2.n57 VDD2.n6 10.4732
R590 VDD2.n129 VDD2.n75 9.69747
R591 VDD2.n104 VDD2.n103 9.69747
R592 VDD2.n32 VDD2.n31 9.69747
R593 VDD2.n58 VDD2.n4 9.69747
R594 VDD2.n139 VDD2.n138 9.45567
R595 VDD2.n68 VDD2.n67 9.45567
R596 VDD2.n97 VDD2.n96 9.3005
R597 VDD2.n99 VDD2.n98 9.3005
R598 VDD2.n90 VDD2.n89 9.3005
R599 VDD2.n105 VDD2.n104 9.3005
R600 VDD2.n107 VDD2.n106 9.3005
R601 VDD2.n85 VDD2.n84 9.3005
R602 VDD2.n113 VDD2.n112 9.3005
R603 VDD2.n115 VDD2.n114 9.3005
R604 VDD2.n138 VDD2.n137 9.3005
R605 VDD2.n73 VDD2.n72 9.3005
R606 VDD2.n132 VDD2.n131 9.3005
R607 VDD2.n130 VDD2.n129 9.3005
R608 VDD2.n77 VDD2.n76 9.3005
R609 VDD2.n124 VDD2.n123 9.3005
R610 VDD2.n122 VDD2.n121 9.3005
R611 VDD2.n81 VDD2.n80 9.3005
R612 VDD2.n2 VDD2.n1 9.3005
R613 VDD2.n61 VDD2.n60 9.3005
R614 VDD2.n59 VDD2.n58 9.3005
R615 VDD2.n6 VDD2.n5 9.3005
R616 VDD2.n53 VDD2.n52 9.3005
R617 VDD2.n51 VDD2.n50 9.3005
R618 VDD2.n10 VDD2.n9 9.3005
R619 VDD2.n25 VDD2.n24 9.3005
R620 VDD2.n27 VDD2.n26 9.3005
R621 VDD2.n18 VDD2.n17 9.3005
R622 VDD2.n33 VDD2.n32 9.3005
R623 VDD2.n35 VDD2.n34 9.3005
R624 VDD2.n14 VDD2.n13 9.3005
R625 VDD2.n42 VDD2.n41 9.3005
R626 VDD2.n44 VDD2.n43 9.3005
R627 VDD2.n67 VDD2.n66 9.3005
R628 VDD2.n133 VDD2.n132 8.92171
R629 VDD2.n100 VDD2.n90 8.92171
R630 VDD2.n28 VDD2.n18 8.92171
R631 VDD2.n62 VDD2.n61 8.92171
R632 VDD2.n136 VDD2.n73 8.14595
R633 VDD2.n99 VDD2.n92 8.14595
R634 VDD2.n27 VDD2.n20 8.14595
R635 VDD2.n65 VDD2.n2 8.14595
R636 VDD2.n137 VDD2.n71 7.3702
R637 VDD2.n96 VDD2.n95 7.3702
R638 VDD2.n24 VDD2.n23 7.3702
R639 VDD2.n66 VDD2.n0 7.3702
R640 VDD2.n139 VDD2.n71 6.59444
R641 VDD2.n68 VDD2.n0 6.59444
R642 VDD2.n137 VDD2.n136 5.81868
R643 VDD2.n96 VDD2.n92 5.81868
R644 VDD2.n24 VDD2.n20 5.81868
R645 VDD2.n66 VDD2.n65 5.81868
R646 VDD2.n133 VDD2.n73 5.04292
R647 VDD2.n100 VDD2.n99 5.04292
R648 VDD2.n28 VDD2.n27 5.04292
R649 VDD2.n62 VDD2.n2 5.04292
R650 VDD2.n132 VDD2.n75 4.26717
R651 VDD2.n103 VDD2.n90 4.26717
R652 VDD2.n31 VDD2.n18 4.26717
R653 VDD2.n61 VDD2.n4 4.26717
R654 VDD2.n129 VDD2.n128 3.49141
R655 VDD2.n104 VDD2.n88 3.49141
R656 VDD2.n32 VDD2.n16 3.49141
R657 VDD2.n58 VDD2.n57 3.49141
R658 VDD2.n125 VDD2.n77 2.71565
R659 VDD2.n108 VDD2.n107 2.71565
R660 VDD2.n36 VDD2.n35 2.71565
R661 VDD2.n54 VDD2.n6 2.71565
R662 VDD2.n141 VDD2.t1 2.52027
R663 VDD2.n141 VDD2.t2 2.52027
R664 VDD2.n69 VDD2.t3 2.52027
R665 VDD2.n69 VDD2.t5 2.52027
R666 VDD2.n97 VDD2.n93 2.41282
R667 VDD2.n25 VDD2.n21 2.41282
R668 VDD2 VDD2.n140 2.03714
R669 VDD2.n124 VDD2.n79 1.93989
R670 VDD2.n111 VDD2.n85 1.93989
R671 VDD2.n40 VDD2.n14 1.93989
R672 VDD2.n53 VDD2.n8 1.93989
R673 VDD2.n121 VDD2.n120 1.16414
R674 VDD2.n112 VDD2.n83 1.16414
R675 VDD2.n41 VDD2.n12 1.16414
R676 VDD2.n50 VDD2.n49 1.16414
R677 VDD2.n117 VDD2.n81 0.388379
R678 VDD2.n116 VDD2.n115 0.388379
R679 VDD2.n45 VDD2.n44 0.388379
R680 VDD2.n46 VDD2.n10 0.388379
R681 VDD2.n138 VDD2.n72 0.155672
R682 VDD2.n131 VDD2.n72 0.155672
R683 VDD2.n131 VDD2.n130 0.155672
R684 VDD2.n130 VDD2.n76 0.155672
R685 VDD2.n123 VDD2.n76 0.155672
R686 VDD2.n123 VDD2.n122 0.155672
R687 VDD2.n122 VDD2.n80 0.155672
R688 VDD2.n114 VDD2.n80 0.155672
R689 VDD2.n114 VDD2.n113 0.155672
R690 VDD2.n113 VDD2.n84 0.155672
R691 VDD2.n106 VDD2.n84 0.155672
R692 VDD2.n106 VDD2.n105 0.155672
R693 VDD2.n105 VDD2.n89 0.155672
R694 VDD2.n98 VDD2.n89 0.155672
R695 VDD2.n98 VDD2.n97 0.155672
R696 VDD2.n26 VDD2.n25 0.155672
R697 VDD2.n26 VDD2.n17 0.155672
R698 VDD2.n33 VDD2.n17 0.155672
R699 VDD2.n34 VDD2.n33 0.155672
R700 VDD2.n34 VDD2.n13 0.155672
R701 VDD2.n42 VDD2.n13 0.155672
R702 VDD2.n43 VDD2.n42 0.155672
R703 VDD2.n43 VDD2.n9 0.155672
R704 VDD2.n51 VDD2.n9 0.155672
R705 VDD2.n52 VDD2.n51 0.155672
R706 VDD2.n52 VDD2.n5 0.155672
R707 VDD2.n59 VDD2.n5 0.155672
R708 VDD2.n60 VDD2.n59 0.155672
R709 VDD2.n60 VDD2.n1 0.155672
R710 VDD2.n67 VDD2.n1 0.155672
R711 VP.n13 VP.n12 161.3
R712 VP.n14 VP.n9 161.3
R713 VP.n16 VP.n15 161.3
R714 VP.n17 VP.n8 161.3
R715 VP.n19 VP.n18 161.3
R716 VP.n20 VP.n7 161.3
R717 VP.n43 VP.n0 161.3
R718 VP.n42 VP.n41 161.3
R719 VP.n40 VP.n1 161.3
R720 VP.n39 VP.n38 161.3
R721 VP.n37 VP.n2 161.3
R722 VP.n36 VP.n35 161.3
R723 VP.n34 VP.n3 161.3
R724 VP.n33 VP.n32 161.3
R725 VP.n31 VP.n4 161.3
R726 VP.n30 VP.n29 161.3
R727 VP.n28 VP.n5 161.3
R728 VP.n27 VP.n26 161.3
R729 VP.n25 VP.n6 161.3
R730 VP.n11 VP.t5 147.101
R731 VP.n3 VP.t1 113.879
R732 VP.n24 VP.t4 113.879
R733 VP.n44 VP.t3 113.879
R734 VP.n10 VP.t0 113.879
R735 VP.n21 VP.t2 113.879
R736 VP.n24 VP.n23 107.684
R737 VP.n45 VP.n44 107.684
R738 VP.n22 VP.n21 107.684
R739 VP.n23 VP.n22 49.8101
R740 VP.n11 VP.n10 48.82
R741 VP.n30 VP.n5 43.3318
R742 VP.n38 VP.n1 43.3318
R743 VP.n15 VP.n8 43.3318
R744 VP.n31 VP.n30 37.4894
R745 VP.n38 VP.n37 37.4894
R746 VP.n15 VP.n14 37.4894
R747 VP.n26 VP.n25 24.3439
R748 VP.n26 VP.n5 24.3439
R749 VP.n32 VP.n31 24.3439
R750 VP.n32 VP.n3 24.3439
R751 VP.n36 VP.n3 24.3439
R752 VP.n37 VP.n36 24.3439
R753 VP.n42 VP.n1 24.3439
R754 VP.n43 VP.n42 24.3439
R755 VP.n19 VP.n8 24.3439
R756 VP.n20 VP.n19 24.3439
R757 VP.n13 VP.n10 24.3439
R758 VP.n14 VP.n13 24.3439
R759 VP.n12 VP.n11 5.08087
R760 VP.n25 VP.n24 2.92171
R761 VP.n44 VP.n43 2.92171
R762 VP.n21 VP.n20 2.92171
R763 VP.n22 VP.n7 0.278398
R764 VP.n23 VP.n6 0.278398
R765 VP.n45 VP.n0 0.278398
R766 VP.n12 VP.n9 0.189894
R767 VP.n16 VP.n9 0.189894
R768 VP.n17 VP.n16 0.189894
R769 VP.n18 VP.n17 0.189894
R770 VP.n18 VP.n7 0.189894
R771 VP.n27 VP.n6 0.189894
R772 VP.n28 VP.n27 0.189894
R773 VP.n29 VP.n28 0.189894
R774 VP.n29 VP.n4 0.189894
R775 VP.n33 VP.n4 0.189894
R776 VP.n34 VP.n33 0.189894
R777 VP.n35 VP.n34 0.189894
R778 VP.n35 VP.n2 0.189894
R779 VP.n39 VP.n2 0.189894
R780 VP.n40 VP.n39 0.189894
R781 VP.n41 VP.n40 0.189894
R782 VP.n41 VP.n0 0.189894
R783 VP VP.n45 0.153422
R784 VDD1.n64 VDD1.n0 756.745
R785 VDD1.n133 VDD1.n69 756.745
R786 VDD1.n65 VDD1.n64 585
R787 VDD1.n63 VDD1.n62 585
R788 VDD1.n4 VDD1.n3 585
R789 VDD1.n57 VDD1.n56 585
R790 VDD1.n55 VDD1.n54 585
R791 VDD1.n8 VDD1.n7 585
R792 VDD1.n49 VDD1.n48 585
R793 VDD1.n47 VDD1.n46 585
R794 VDD1.n45 VDD1.n11 585
R795 VDD1.n15 VDD1.n12 585
R796 VDD1.n40 VDD1.n39 585
R797 VDD1.n38 VDD1.n37 585
R798 VDD1.n17 VDD1.n16 585
R799 VDD1.n32 VDD1.n31 585
R800 VDD1.n30 VDD1.n29 585
R801 VDD1.n21 VDD1.n20 585
R802 VDD1.n24 VDD1.n23 585
R803 VDD1.n92 VDD1.n91 585
R804 VDD1.n89 VDD1.n88 585
R805 VDD1.n98 VDD1.n97 585
R806 VDD1.n100 VDD1.n99 585
R807 VDD1.n85 VDD1.n84 585
R808 VDD1.n106 VDD1.n105 585
R809 VDD1.n109 VDD1.n108 585
R810 VDD1.n107 VDD1.n81 585
R811 VDD1.n114 VDD1.n80 585
R812 VDD1.n116 VDD1.n115 585
R813 VDD1.n118 VDD1.n117 585
R814 VDD1.n77 VDD1.n76 585
R815 VDD1.n124 VDD1.n123 585
R816 VDD1.n126 VDD1.n125 585
R817 VDD1.n73 VDD1.n72 585
R818 VDD1.n132 VDD1.n131 585
R819 VDD1.n134 VDD1.n133 585
R820 VDD1.t1 VDD1.n90 329.036
R821 VDD1.t0 VDD1.n22 329.036
R822 VDD1.n64 VDD1.n63 171.744
R823 VDD1.n63 VDD1.n3 171.744
R824 VDD1.n56 VDD1.n3 171.744
R825 VDD1.n56 VDD1.n55 171.744
R826 VDD1.n55 VDD1.n7 171.744
R827 VDD1.n48 VDD1.n7 171.744
R828 VDD1.n48 VDD1.n47 171.744
R829 VDD1.n47 VDD1.n11 171.744
R830 VDD1.n15 VDD1.n11 171.744
R831 VDD1.n39 VDD1.n15 171.744
R832 VDD1.n39 VDD1.n38 171.744
R833 VDD1.n38 VDD1.n16 171.744
R834 VDD1.n31 VDD1.n16 171.744
R835 VDD1.n31 VDD1.n30 171.744
R836 VDD1.n30 VDD1.n20 171.744
R837 VDD1.n23 VDD1.n20 171.744
R838 VDD1.n91 VDD1.n88 171.744
R839 VDD1.n98 VDD1.n88 171.744
R840 VDD1.n99 VDD1.n98 171.744
R841 VDD1.n99 VDD1.n84 171.744
R842 VDD1.n106 VDD1.n84 171.744
R843 VDD1.n108 VDD1.n106 171.744
R844 VDD1.n108 VDD1.n107 171.744
R845 VDD1.n107 VDD1.n80 171.744
R846 VDD1.n116 VDD1.n80 171.744
R847 VDD1.n117 VDD1.n116 171.744
R848 VDD1.n117 VDD1.n76 171.744
R849 VDD1.n124 VDD1.n76 171.744
R850 VDD1.n125 VDD1.n124 171.744
R851 VDD1.n125 VDD1.n72 171.744
R852 VDD1.n132 VDD1.n72 171.744
R853 VDD1.n133 VDD1.n132 171.744
R854 VDD1.n23 VDD1.t0 85.8723
R855 VDD1.n91 VDD1.t1 85.8723
R856 VDD1.n139 VDD1.n138 74.7791
R857 VDD1.n141 VDD1.n140 74.1748
R858 VDD1 VDD1.n68 52.0644
R859 VDD1.n139 VDD1.n137 51.9509
R860 VDD1.n141 VDD1.n139 45.3112
R861 VDD1.n46 VDD1.n45 13.1884
R862 VDD1.n115 VDD1.n114 13.1884
R863 VDD1.n49 VDD1.n10 12.8005
R864 VDD1.n44 VDD1.n12 12.8005
R865 VDD1.n113 VDD1.n81 12.8005
R866 VDD1.n118 VDD1.n79 12.8005
R867 VDD1.n50 VDD1.n8 12.0247
R868 VDD1.n41 VDD1.n40 12.0247
R869 VDD1.n110 VDD1.n109 12.0247
R870 VDD1.n119 VDD1.n77 12.0247
R871 VDD1.n54 VDD1.n53 11.249
R872 VDD1.n37 VDD1.n14 11.249
R873 VDD1.n105 VDD1.n83 11.249
R874 VDD1.n123 VDD1.n122 11.249
R875 VDD1.n24 VDD1.n22 10.7239
R876 VDD1.n92 VDD1.n90 10.7239
R877 VDD1.n57 VDD1.n6 10.4732
R878 VDD1.n36 VDD1.n17 10.4732
R879 VDD1.n104 VDD1.n85 10.4732
R880 VDD1.n126 VDD1.n75 10.4732
R881 VDD1.n58 VDD1.n4 9.69747
R882 VDD1.n33 VDD1.n32 9.69747
R883 VDD1.n101 VDD1.n100 9.69747
R884 VDD1.n127 VDD1.n73 9.69747
R885 VDD1.n68 VDD1.n67 9.45567
R886 VDD1.n137 VDD1.n136 9.45567
R887 VDD1.n26 VDD1.n25 9.3005
R888 VDD1.n28 VDD1.n27 9.3005
R889 VDD1.n19 VDD1.n18 9.3005
R890 VDD1.n34 VDD1.n33 9.3005
R891 VDD1.n36 VDD1.n35 9.3005
R892 VDD1.n14 VDD1.n13 9.3005
R893 VDD1.n42 VDD1.n41 9.3005
R894 VDD1.n44 VDD1.n43 9.3005
R895 VDD1.n67 VDD1.n66 9.3005
R896 VDD1.n2 VDD1.n1 9.3005
R897 VDD1.n61 VDD1.n60 9.3005
R898 VDD1.n59 VDD1.n58 9.3005
R899 VDD1.n6 VDD1.n5 9.3005
R900 VDD1.n53 VDD1.n52 9.3005
R901 VDD1.n51 VDD1.n50 9.3005
R902 VDD1.n10 VDD1.n9 9.3005
R903 VDD1.n71 VDD1.n70 9.3005
R904 VDD1.n130 VDD1.n129 9.3005
R905 VDD1.n128 VDD1.n127 9.3005
R906 VDD1.n75 VDD1.n74 9.3005
R907 VDD1.n122 VDD1.n121 9.3005
R908 VDD1.n120 VDD1.n119 9.3005
R909 VDD1.n79 VDD1.n78 9.3005
R910 VDD1.n94 VDD1.n93 9.3005
R911 VDD1.n96 VDD1.n95 9.3005
R912 VDD1.n87 VDD1.n86 9.3005
R913 VDD1.n102 VDD1.n101 9.3005
R914 VDD1.n104 VDD1.n103 9.3005
R915 VDD1.n83 VDD1.n82 9.3005
R916 VDD1.n111 VDD1.n110 9.3005
R917 VDD1.n113 VDD1.n112 9.3005
R918 VDD1.n136 VDD1.n135 9.3005
R919 VDD1.n62 VDD1.n61 8.92171
R920 VDD1.n29 VDD1.n19 8.92171
R921 VDD1.n97 VDD1.n87 8.92171
R922 VDD1.n131 VDD1.n130 8.92171
R923 VDD1.n65 VDD1.n2 8.14595
R924 VDD1.n28 VDD1.n21 8.14595
R925 VDD1.n96 VDD1.n89 8.14595
R926 VDD1.n134 VDD1.n71 8.14595
R927 VDD1.n66 VDD1.n0 7.3702
R928 VDD1.n25 VDD1.n24 7.3702
R929 VDD1.n93 VDD1.n92 7.3702
R930 VDD1.n135 VDD1.n69 7.3702
R931 VDD1.n68 VDD1.n0 6.59444
R932 VDD1.n137 VDD1.n69 6.59444
R933 VDD1.n66 VDD1.n65 5.81868
R934 VDD1.n25 VDD1.n21 5.81868
R935 VDD1.n93 VDD1.n89 5.81868
R936 VDD1.n135 VDD1.n134 5.81868
R937 VDD1.n62 VDD1.n2 5.04292
R938 VDD1.n29 VDD1.n28 5.04292
R939 VDD1.n97 VDD1.n96 5.04292
R940 VDD1.n131 VDD1.n71 5.04292
R941 VDD1.n61 VDD1.n4 4.26717
R942 VDD1.n32 VDD1.n19 4.26717
R943 VDD1.n100 VDD1.n87 4.26717
R944 VDD1.n130 VDD1.n73 4.26717
R945 VDD1.n58 VDD1.n57 3.49141
R946 VDD1.n33 VDD1.n17 3.49141
R947 VDD1.n101 VDD1.n85 3.49141
R948 VDD1.n127 VDD1.n126 3.49141
R949 VDD1.n54 VDD1.n6 2.71565
R950 VDD1.n37 VDD1.n36 2.71565
R951 VDD1.n105 VDD1.n104 2.71565
R952 VDD1.n123 VDD1.n75 2.71565
R953 VDD1.n140 VDD1.t5 2.52027
R954 VDD1.n140 VDD1.t3 2.52027
R955 VDD1.n138 VDD1.t4 2.52027
R956 VDD1.n138 VDD1.t2 2.52027
R957 VDD1.n26 VDD1.n22 2.41282
R958 VDD1.n94 VDD1.n90 2.41282
R959 VDD1.n53 VDD1.n8 1.93989
R960 VDD1.n40 VDD1.n14 1.93989
R961 VDD1.n109 VDD1.n83 1.93989
R962 VDD1.n122 VDD1.n77 1.93989
R963 VDD1.n50 VDD1.n49 1.16414
R964 VDD1.n41 VDD1.n12 1.16414
R965 VDD1.n110 VDD1.n81 1.16414
R966 VDD1.n119 VDD1.n118 1.16414
R967 VDD1 VDD1.n141 0.601793
R968 VDD1.n46 VDD1.n10 0.388379
R969 VDD1.n45 VDD1.n44 0.388379
R970 VDD1.n114 VDD1.n113 0.388379
R971 VDD1.n115 VDD1.n79 0.388379
R972 VDD1.n67 VDD1.n1 0.155672
R973 VDD1.n60 VDD1.n1 0.155672
R974 VDD1.n60 VDD1.n59 0.155672
R975 VDD1.n59 VDD1.n5 0.155672
R976 VDD1.n52 VDD1.n5 0.155672
R977 VDD1.n52 VDD1.n51 0.155672
R978 VDD1.n51 VDD1.n9 0.155672
R979 VDD1.n43 VDD1.n9 0.155672
R980 VDD1.n43 VDD1.n42 0.155672
R981 VDD1.n42 VDD1.n13 0.155672
R982 VDD1.n35 VDD1.n13 0.155672
R983 VDD1.n35 VDD1.n34 0.155672
R984 VDD1.n34 VDD1.n18 0.155672
R985 VDD1.n27 VDD1.n18 0.155672
R986 VDD1.n27 VDD1.n26 0.155672
R987 VDD1.n95 VDD1.n94 0.155672
R988 VDD1.n95 VDD1.n86 0.155672
R989 VDD1.n102 VDD1.n86 0.155672
R990 VDD1.n103 VDD1.n102 0.155672
R991 VDD1.n103 VDD1.n82 0.155672
R992 VDD1.n111 VDD1.n82 0.155672
R993 VDD1.n112 VDD1.n111 0.155672
R994 VDD1.n112 VDD1.n78 0.155672
R995 VDD1.n120 VDD1.n78 0.155672
R996 VDD1.n121 VDD1.n120 0.155672
R997 VDD1.n121 VDD1.n74 0.155672
R998 VDD1.n128 VDD1.n74 0.155672
R999 VDD1.n129 VDD1.n128 0.155672
R1000 VDD1.n129 VDD1.n70 0.155672
R1001 VDD1.n136 VDD1.n70 0.155672
R1002 B.n544 B.n77 585
R1003 B.n546 B.n545 585
R1004 B.n547 B.n76 585
R1005 B.n549 B.n548 585
R1006 B.n550 B.n75 585
R1007 B.n552 B.n551 585
R1008 B.n553 B.n74 585
R1009 B.n555 B.n554 585
R1010 B.n556 B.n73 585
R1011 B.n558 B.n557 585
R1012 B.n559 B.n72 585
R1013 B.n561 B.n560 585
R1014 B.n562 B.n71 585
R1015 B.n564 B.n563 585
R1016 B.n565 B.n70 585
R1017 B.n567 B.n566 585
R1018 B.n568 B.n69 585
R1019 B.n570 B.n569 585
R1020 B.n571 B.n68 585
R1021 B.n573 B.n572 585
R1022 B.n574 B.n67 585
R1023 B.n576 B.n575 585
R1024 B.n577 B.n66 585
R1025 B.n579 B.n578 585
R1026 B.n580 B.n65 585
R1027 B.n582 B.n581 585
R1028 B.n583 B.n64 585
R1029 B.n585 B.n584 585
R1030 B.n586 B.n63 585
R1031 B.n588 B.n587 585
R1032 B.n589 B.n62 585
R1033 B.n591 B.n590 585
R1034 B.n592 B.n61 585
R1035 B.n594 B.n593 585
R1036 B.n595 B.n60 585
R1037 B.n597 B.n596 585
R1038 B.n598 B.n59 585
R1039 B.n600 B.n599 585
R1040 B.n601 B.n58 585
R1041 B.n603 B.n602 585
R1042 B.n604 B.n57 585
R1043 B.n606 B.n605 585
R1044 B.n607 B.n56 585
R1045 B.n609 B.n608 585
R1046 B.n611 B.n53 585
R1047 B.n613 B.n612 585
R1048 B.n614 B.n52 585
R1049 B.n616 B.n615 585
R1050 B.n617 B.n51 585
R1051 B.n619 B.n618 585
R1052 B.n620 B.n50 585
R1053 B.n622 B.n621 585
R1054 B.n623 B.n49 585
R1055 B.n625 B.n624 585
R1056 B.n627 B.n626 585
R1057 B.n628 B.n45 585
R1058 B.n630 B.n629 585
R1059 B.n631 B.n44 585
R1060 B.n633 B.n632 585
R1061 B.n634 B.n43 585
R1062 B.n636 B.n635 585
R1063 B.n637 B.n42 585
R1064 B.n639 B.n638 585
R1065 B.n640 B.n41 585
R1066 B.n642 B.n641 585
R1067 B.n643 B.n40 585
R1068 B.n645 B.n644 585
R1069 B.n646 B.n39 585
R1070 B.n648 B.n647 585
R1071 B.n649 B.n38 585
R1072 B.n651 B.n650 585
R1073 B.n652 B.n37 585
R1074 B.n654 B.n653 585
R1075 B.n655 B.n36 585
R1076 B.n657 B.n656 585
R1077 B.n658 B.n35 585
R1078 B.n660 B.n659 585
R1079 B.n661 B.n34 585
R1080 B.n663 B.n662 585
R1081 B.n664 B.n33 585
R1082 B.n666 B.n665 585
R1083 B.n667 B.n32 585
R1084 B.n669 B.n668 585
R1085 B.n670 B.n31 585
R1086 B.n672 B.n671 585
R1087 B.n673 B.n30 585
R1088 B.n675 B.n674 585
R1089 B.n676 B.n29 585
R1090 B.n678 B.n677 585
R1091 B.n679 B.n28 585
R1092 B.n681 B.n680 585
R1093 B.n682 B.n27 585
R1094 B.n684 B.n683 585
R1095 B.n685 B.n26 585
R1096 B.n687 B.n686 585
R1097 B.n688 B.n25 585
R1098 B.n690 B.n689 585
R1099 B.n691 B.n24 585
R1100 B.n543 B.n542 585
R1101 B.n541 B.n78 585
R1102 B.n540 B.n539 585
R1103 B.n538 B.n79 585
R1104 B.n537 B.n536 585
R1105 B.n535 B.n80 585
R1106 B.n534 B.n533 585
R1107 B.n532 B.n81 585
R1108 B.n531 B.n530 585
R1109 B.n529 B.n82 585
R1110 B.n528 B.n527 585
R1111 B.n526 B.n83 585
R1112 B.n525 B.n524 585
R1113 B.n523 B.n84 585
R1114 B.n522 B.n521 585
R1115 B.n520 B.n85 585
R1116 B.n519 B.n518 585
R1117 B.n517 B.n86 585
R1118 B.n516 B.n515 585
R1119 B.n514 B.n87 585
R1120 B.n513 B.n512 585
R1121 B.n511 B.n88 585
R1122 B.n510 B.n509 585
R1123 B.n508 B.n89 585
R1124 B.n507 B.n506 585
R1125 B.n505 B.n90 585
R1126 B.n504 B.n503 585
R1127 B.n502 B.n91 585
R1128 B.n501 B.n500 585
R1129 B.n499 B.n92 585
R1130 B.n498 B.n497 585
R1131 B.n496 B.n93 585
R1132 B.n495 B.n494 585
R1133 B.n493 B.n94 585
R1134 B.n492 B.n491 585
R1135 B.n490 B.n95 585
R1136 B.n489 B.n488 585
R1137 B.n487 B.n96 585
R1138 B.n486 B.n485 585
R1139 B.n484 B.n97 585
R1140 B.n483 B.n482 585
R1141 B.n481 B.n98 585
R1142 B.n480 B.n479 585
R1143 B.n478 B.n99 585
R1144 B.n477 B.n476 585
R1145 B.n475 B.n100 585
R1146 B.n474 B.n473 585
R1147 B.n472 B.n101 585
R1148 B.n471 B.n470 585
R1149 B.n469 B.n102 585
R1150 B.n468 B.n467 585
R1151 B.n466 B.n103 585
R1152 B.n465 B.n464 585
R1153 B.n463 B.n104 585
R1154 B.n462 B.n461 585
R1155 B.n460 B.n105 585
R1156 B.n459 B.n458 585
R1157 B.n457 B.n106 585
R1158 B.n456 B.n455 585
R1159 B.n454 B.n107 585
R1160 B.n453 B.n452 585
R1161 B.n451 B.n108 585
R1162 B.n450 B.n449 585
R1163 B.n448 B.n109 585
R1164 B.n447 B.n446 585
R1165 B.n445 B.n110 585
R1166 B.n444 B.n443 585
R1167 B.n442 B.n111 585
R1168 B.n441 B.n440 585
R1169 B.n439 B.n112 585
R1170 B.n438 B.n437 585
R1171 B.n436 B.n113 585
R1172 B.n435 B.n434 585
R1173 B.n433 B.n114 585
R1174 B.n432 B.n431 585
R1175 B.n430 B.n115 585
R1176 B.n429 B.n428 585
R1177 B.n427 B.n116 585
R1178 B.n426 B.n425 585
R1179 B.n424 B.n117 585
R1180 B.n423 B.n422 585
R1181 B.n421 B.n118 585
R1182 B.n420 B.n419 585
R1183 B.n418 B.n119 585
R1184 B.n417 B.n416 585
R1185 B.n415 B.n120 585
R1186 B.n414 B.n413 585
R1187 B.n412 B.n121 585
R1188 B.n411 B.n410 585
R1189 B.n262 B.n175 585
R1190 B.n264 B.n263 585
R1191 B.n265 B.n174 585
R1192 B.n267 B.n266 585
R1193 B.n268 B.n173 585
R1194 B.n270 B.n269 585
R1195 B.n271 B.n172 585
R1196 B.n273 B.n272 585
R1197 B.n274 B.n171 585
R1198 B.n276 B.n275 585
R1199 B.n277 B.n170 585
R1200 B.n279 B.n278 585
R1201 B.n280 B.n169 585
R1202 B.n282 B.n281 585
R1203 B.n283 B.n168 585
R1204 B.n285 B.n284 585
R1205 B.n286 B.n167 585
R1206 B.n288 B.n287 585
R1207 B.n289 B.n166 585
R1208 B.n291 B.n290 585
R1209 B.n292 B.n165 585
R1210 B.n294 B.n293 585
R1211 B.n295 B.n164 585
R1212 B.n297 B.n296 585
R1213 B.n298 B.n163 585
R1214 B.n300 B.n299 585
R1215 B.n301 B.n162 585
R1216 B.n303 B.n302 585
R1217 B.n304 B.n161 585
R1218 B.n306 B.n305 585
R1219 B.n307 B.n160 585
R1220 B.n309 B.n308 585
R1221 B.n310 B.n159 585
R1222 B.n312 B.n311 585
R1223 B.n313 B.n158 585
R1224 B.n315 B.n314 585
R1225 B.n316 B.n157 585
R1226 B.n318 B.n317 585
R1227 B.n319 B.n156 585
R1228 B.n321 B.n320 585
R1229 B.n322 B.n155 585
R1230 B.n324 B.n323 585
R1231 B.n325 B.n154 585
R1232 B.n327 B.n326 585
R1233 B.n329 B.n151 585
R1234 B.n331 B.n330 585
R1235 B.n332 B.n150 585
R1236 B.n334 B.n333 585
R1237 B.n335 B.n149 585
R1238 B.n337 B.n336 585
R1239 B.n338 B.n148 585
R1240 B.n340 B.n339 585
R1241 B.n341 B.n147 585
R1242 B.n343 B.n342 585
R1243 B.n345 B.n344 585
R1244 B.n346 B.n143 585
R1245 B.n348 B.n347 585
R1246 B.n349 B.n142 585
R1247 B.n351 B.n350 585
R1248 B.n352 B.n141 585
R1249 B.n354 B.n353 585
R1250 B.n355 B.n140 585
R1251 B.n357 B.n356 585
R1252 B.n358 B.n139 585
R1253 B.n360 B.n359 585
R1254 B.n361 B.n138 585
R1255 B.n363 B.n362 585
R1256 B.n364 B.n137 585
R1257 B.n366 B.n365 585
R1258 B.n367 B.n136 585
R1259 B.n369 B.n368 585
R1260 B.n370 B.n135 585
R1261 B.n372 B.n371 585
R1262 B.n373 B.n134 585
R1263 B.n375 B.n374 585
R1264 B.n376 B.n133 585
R1265 B.n378 B.n377 585
R1266 B.n379 B.n132 585
R1267 B.n381 B.n380 585
R1268 B.n382 B.n131 585
R1269 B.n384 B.n383 585
R1270 B.n385 B.n130 585
R1271 B.n387 B.n386 585
R1272 B.n388 B.n129 585
R1273 B.n390 B.n389 585
R1274 B.n391 B.n128 585
R1275 B.n393 B.n392 585
R1276 B.n394 B.n127 585
R1277 B.n396 B.n395 585
R1278 B.n397 B.n126 585
R1279 B.n399 B.n398 585
R1280 B.n400 B.n125 585
R1281 B.n402 B.n401 585
R1282 B.n403 B.n124 585
R1283 B.n405 B.n404 585
R1284 B.n406 B.n123 585
R1285 B.n408 B.n407 585
R1286 B.n409 B.n122 585
R1287 B.n261 B.n260 585
R1288 B.n259 B.n176 585
R1289 B.n258 B.n257 585
R1290 B.n256 B.n177 585
R1291 B.n255 B.n254 585
R1292 B.n253 B.n178 585
R1293 B.n252 B.n251 585
R1294 B.n250 B.n179 585
R1295 B.n249 B.n248 585
R1296 B.n247 B.n180 585
R1297 B.n246 B.n245 585
R1298 B.n244 B.n181 585
R1299 B.n243 B.n242 585
R1300 B.n241 B.n182 585
R1301 B.n240 B.n239 585
R1302 B.n238 B.n183 585
R1303 B.n237 B.n236 585
R1304 B.n235 B.n184 585
R1305 B.n234 B.n233 585
R1306 B.n232 B.n185 585
R1307 B.n231 B.n230 585
R1308 B.n229 B.n186 585
R1309 B.n228 B.n227 585
R1310 B.n226 B.n187 585
R1311 B.n225 B.n224 585
R1312 B.n223 B.n188 585
R1313 B.n222 B.n221 585
R1314 B.n220 B.n189 585
R1315 B.n219 B.n218 585
R1316 B.n217 B.n190 585
R1317 B.n216 B.n215 585
R1318 B.n214 B.n191 585
R1319 B.n213 B.n212 585
R1320 B.n211 B.n192 585
R1321 B.n210 B.n209 585
R1322 B.n208 B.n193 585
R1323 B.n207 B.n206 585
R1324 B.n205 B.n194 585
R1325 B.n204 B.n203 585
R1326 B.n202 B.n195 585
R1327 B.n201 B.n200 585
R1328 B.n199 B.n196 585
R1329 B.n198 B.n197 585
R1330 B.n2 B.n0 585
R1331 B.n757 B.n1 585
R1332 B.n756 B.n755 585
R1333 B.n754 B.n3 585
R1334 B.n753 B.n752 585
R1335 B.n751 B.n4 585
R1336 B.n750 B.n749 585
R1337 B.n748 B.n5 585
R1338 B.n747 B.n746 585
R1339 B.n745 B.n6 585
R1340 B.n744 B.n743 585
R1341 B.n742 B.n7 585
R1342 B.n741 B.n740 585
R1343 B.n739 B.n8 585
R1344 B.n738 B.n737 585
R1345 B.n736 B.n9 585
R1346 B.n735 B.n734 585
R1347 B.n733 B.n10 585
R1348 B.n732 B.n731 585
R1349 B.n730 B.n11 585
R1350 B.n729 B.n728 585
R1351 B.n727 B.n12 585
R1352 B.n726 B.n725 585
R1353 B.n724 B.n13 585
R1354 B.n723 B.n722 585
R1355 B.n721 B.n14 585
R1356 B.n720 B.n719 585
R1357 B.n718 B.n15 585
R1358 B.n717 B.n716 585
R1359 B.n715 B.n16 585
R1360 B.n714 B.n713 585
R1361 B.n712 B.n17 585
R1362 B.n711 B.n710 585
R1363 B.n709 B.n18 585
R1364 B.n708 B.n707 585
R1365 B.n706 B.n19 585
R1366 B.n705 B.n704 585
R1367 B.n703 B.n20 585
R1368 B.n702 B.n701 585
R1369 B.n700 B.n21 585
R1370 B.n699 B.n698 585
R1371 B.n697 B.n22 585
R1372 B.n696 B.n695 585
R1373 B.n694 B.n23 585
R1374 B.n693 B.n692 585
R1375 B.n759 B.n758 585
R1376 B.n260 B.n175 526.135
R1377 B.n692 B.n691 526.135
R1378 B.n410 B.n409 526.135
R1379 B.n542 B.n77 526.135
R1380 B.n144 B.t11 451.389
R1381 B.n54 B.t4 451.389
R1382 B.n152 B.t2 451.389
R1383 B.n46 B.t7 451.389
R1384 B.n145 B.t10 392.043
R1385 B.n55 B.t5 392.043
R1386 B.n153 B.t1 392.043
R1387 B.n47 B.t8 392.043
R1388 B.n144 B.t9 322.115
R1389 B.n152 B.t0 322.115
R1390 B.n46 B.t6 322.115
R1391 B.n54 B.t3 322.115
R1392 B.n260 B.n259 163.367
R1393 B.n259 B.n258 163.367
R1394 B.n258 B.n177 163.367
R1395 B.n254 B.n177 163.367
R1396 B.n254 B.n253 163.367
R1397 B.n253 B.n252 163.367
R1398 B.n252 B.n179 163.367
R1399 B.n248 B.n179 163.367
R1400 B.n248 B.n247 163.367
R1401 B.n247 B.n246 163.367
R1402 B.n246 B.n181 163.367
R1403 B.n242 B.n181 163.367
R1404 B.n242 B.n241 163.367
R1405 B.n241 B.n240 163.367
R1406 B.n240 B.n183 163.367
R1407 B.n236 B.n183 163.367
R1408 B.n236 B.n235 163.367
R1409 B.n235 B.n234 163.367
R1410 B.n234 B.n185 163.367
R1411 B.n230 B.n185 163.367
R1412 B.n230 B.n229 163.367
R1413 B.n229 B.n228 163.367
R1414 B.n228 B.n187 163.367
R1415 B.n224 B.n187 163.367
R1416 B.n224 B.n223 163.367
R1417 B.n223 B.n222 163.367
R1418 B.n222 B.n189 163.367
R1419 B.n218 B.n189 163.367
R1420 B.n218 B.n217 163.367
R1421 B.n217 B.n216 163.367
R1422 B.n216 B.n191 163.367
R1423 B.n212 B.n191 163.367
R1424 B.n212 B.n211 163.367
R1425 B.n211 B.n210 163.367
R1426 B.n210 B.n193 163.367
R1427 B.n206 B.n193 163.367
R1428 B.n206 B.n205 163.367
R1429 B.n205 B.n204 163.367
R1430 B.n204 B.n195 163.367
R1431 B.n200 B.n195 163.367
R1432 B.n200 B.n199 163.367
R1433 B.n199 B.n198 163.367
R1434 B.n198 B.n2 163.367
R1435 B.n758 B.n2 163.367
R1436 B.n758 B.n757 163.367
R1437 B.n757 B.n756 163.367
R1438 B.n756 B.n3 163.367
R1439 B.n752 B.n3 163.367
R1440 B.n752 B.n751 163.367
R1441 B.n751 B.n750 163.367
R1442 B.n750 B.n5 163.367
R1443 B.n746 B.n5 163.367
R1444 B.n746 B.n745 163.367
R1445 B.n745 B.n744 163.367
R1446 B.n744 B.n7 163.367
R1447 B.n740 B.n7 163.367
R1448 B.n740 B.n739 163.367
R1449 B.n739 B.n738 163.367
R1450 B.n738 B.n9 163.367
R1451 B.n734 B.n9 163.367
R1452 B.n734 B.n733 163.367
R1453 B.n733 B.n732 163.367
R1454 B.n732 B.n11 163.367
R1455 B.n728 B.n11 163.367
R1456 B.n728 B.n727 163.367
R1457 B.n727 B.n726 163.367
R1458 B.n726 B.n13 163.367
R1459 B.n722 B.n13 163.367
R1460 B.n722 B.n721 163.367
R1461 B.n721 B.n720 163.367
R1462 B.n720 B.n15 163.367
R1463 B.n716 B.n15 163.367
R1464 B.n716 B.n715 163.367
R1465 B.n715 B.n714 163.367
R1466 B.n714 B.n17 163.367
R1467 B.n710 B.n17 163.367
R1468 B.n710 B.n709 163.367
R1469 B.n709 B.n708 163.367
R1470 B.n708 B.n19 163.367
R1471 B.n704 B.n19 163.367
R1472 B.n704 B.n703 163.367
R1473 B.n703 B.n702 163.367
R1474 B.n702 B.n21 163.367
R1475 B.n698 B.n21 163.367
R1476 B.n698 B.n697 163.367
R1477 B.n697 B.n696 163.367
R1478 B.n696 B.n23 163.367
R1479 B.n692 B.n23 163.367
R1480 B.n264 B.n175 163.367
R1481 B.n265 B.n264 163.367
R1482 B.n266 B.n265 163.367
R1483 B.n266 B.n173 163.367
R1484 B.n270 B.n173 163.367
R1485 B.n271 B.n270 163.367
R1486 B.n272 B.n271 163.367
R1487 B.n272 B.n171 163.367
R1488 B.n276 B.n171 163.367
R1489 B.n277 B.n276 163.367
R1490 B.n278 B.n277 163.367
R1491 B.n278 B.n169 163.367
R1492 B.n282 B.n169 163.367
R1493 B.n283 B.n282 163.367
R1494 B.n284 B.n283 163.367
R1495 B.n284 B.n167 163.367
R1496 B.n288 B.n167 163.367
R1497 B.n289 B.n288 163.367
R1498 B.n290 B.n289 163.367
R1499 B.n290 B.n165 163.367
R1500 B.n294 B.n165 163.367
R1501 B.n295 B.n294 163.367
R1502 B.n296 B.n295 163.367
R1503 B.n296 B.n163 163.367
R1504 B.n300 B.n163 163.367
R1505 B.n301 B.n300 163.367
R1506 B.n302 B.n301 163.367
R1507 B.n302 B.n161 163.367
R1508 B.n306 B.n161 163.367
R1509 B.n307 B.n306 163.367
R1510 B.n308 B.n307 163.367
R1511 B.n308 B.n159 163.367
R1512 B.n312 B.n159 163.367
R1513 B.n313 B.n312 163.367
R1514 B.n314 B.n313 163.367
R1515 B.n314 B.n157 163.367
R1516 B.n318 B.n157 163.367
R1517 B.n319 B.n318 163.367
R1518 B.n320 B.n319 163.367
R1519 B.n320 B.n155 163.367
R1520 B.n324 B.n155 163.367
R1521 B.n325 B.n324 163.367
R1522 B.n326 B.n325 163.367
R1523 B.n326 B.n151 163.367
R1524 B.n331 B.n151 163.367
R1525 B.n332 B.n331 163.367
R1526 B.n333 B.n332 163.367
R1527 B.n333 B.n149 163.367
R1528 B.n337 B.n149 163.367
R1529 B.n338 B.n337 163.367
R1530 B.n339 B.n338 163.367
R1531 B.n339 B.n147 163.367
R1532 B.n343 B.n147 163.367
R1533 B.n344 B.n343 163.367
R1534 B.n344 B.n143 163.367
R1535 B.n348 B.n143 163.367
R1536 B.n349 B.n348 163.367
R1537 B.n350 B.n349 163.367
R1538 B.n350 B.n141 163.367
R1539 B.n354 B.n141 163.367
R1540 B.n355 B.n354 163.367
R1541 B.n356 B.n355 163.367
R1542 B.n356 B.n139 163.367
R1543 B.n360 B.n139 163.367
R1544 B.n361 B.n360 163.367
R1545 B.n362 B.n361 163.367
R1546 B.n362 B.n137 163.367
R1547 B.n366 B.n137 163.367
R1548 B.n367 B.n366 163.367
R1549 B.n368 B.n367 163.367
R1550 B.n368 B.n135 163.367
R1551 B.n372 B.n135 163.367
R1552 B.n373 B.n372 163.367
R1553 B.n374 B.n373 163.367
R1554 B.n374 B.n133 163.367
R1555 B.n378 B.n133 163.367
R1556 B.n379 B.n378 163.367
R1557 B.n380 B.n379 163.367
R1558 B.n380 B.n131 163.367
R1559 B.n384 B.n131 163.367
R1560 B.n385 B.n384 163.367
R1561 B.n386 B.n385 163.367
R1562 B.n386 B.n129 163.367
R1563 B.n390 B.n129 163.367
R1564 B.n391 B.n390 163.367
R1565 B.n392 B.n391 163.367
R1566 B.n392 B.n127 163.367
R1567 B.n396 B.n127 163.367
R1568 B.n397 B.n396 163.367
R1569 B.n398 B.n397 163.367
R1570 B.n398 B.n125 163.367
R1571 B.n402 B.n125 163.367
R1572 B.n403 B.n402 163.367
R1573 B.n404 B.n403 163.367
R1574 B.n404 B.n123 163.367
R1575 B.n408 B.n123 163.367
R1576 B.n409 B.n408 163.367
R1577 B.n410 B.n121 163.367
R1578 B.n414 B.n121 163.367
R1579 B.n415 B.n414 163.367
R1580 B.n416 B.n415 163.367
R1581 B.n416 B.n119 163.367
R1582 B.n420 B.n119 163.367
R1583 B.n421 B.n420 163.367
R1584 B.n422 B.n421 163.367
R1585 B.n422 B.n117 163.367
R1586 B.n426 B.n117 163.367
R1587 B.n427 B.n426 163.367
R1588 B.n428 B.n427 163.367
R1589 B.n428 B.n115 163.367
R1590 B.n432 B.n115 163.367
R1591 B.n433 B.n432 163.367
R1592 B.n434 B.n433 163.367
R1593 B.n434 B.n113 163.367
R1594 B.n438 B.n113 163.367
R1595 B.n439 B.n438 163.367
R1596 B.n440 B.n439 163.367
R1597 B.n440 B.n111 163.367
R1598 B.n444 B.n111 163.367
R1599 B.n445 B.n444 163.367
R1600 B.n446 B.n445 163.367
R1601 B.n446 B.n109 163.367
R1602 B.n450 B.n109 163.367
R1603 B.n451 B.n450 163.367
R1604 B.n452 B.n451 163.367
R1605 B.n452 B.n107 163.367
R1606 B.n456 B.n107 163.367
R1607 B.n457 B.n456 163.367
R1608 B.n458 B.n457 163.367
R1609 B.n458 B.n105 163.367
R1610 B.n462 B.n105 163.367
R1611 B.n463 B.n462 163.367
R1612 B.n464 B.n463 163.367
R1613 B.n464 B.n103 163.367
R1614 B.n468 B.n103 163.367
R1615 B.n469 B.n468 163.367
R1616 B.n470 B.n469 163.367
R1617 B.n470 B.n101 163.367
R1618 B.n474 B.n101 163.367
R1619 B.n475 B.n474 163.367
R1620 B.n476 B.n475 163.367
R1621 B.n476 B.n99 163.367
R1622 B.n480 B.n99 163.367
R1623 B.n481 B.n480 163.367
R1624 B.n482 B.n481 163.367
R1625 B.n482 B.n97 163.367
R1626 B.n486 B.n97 163.367
R1627 B.n487 B.n486 163.367
R1628 B.n488 B.n487 163.367
R1629 B.n488 B.n95 163.367
R1630 B.n492 B.n95 163.367
R1631 B.n493 B.n492 163.367
R1632 B.n494 B.n493 163.367
R1633 B.n494 B.n93 163.367
R1634 B.n498 B.n93 163.367
R1635 B.n499 B.n498 163.367
R1636 B.n500 B.n499 163.367
R1637 B.n500 B.n91 163.367
R1638 B.n504 B.n91 163.367
R1639 B.n505 B.n504 163.367
R1640 B.n506 B.n505 163.367
R1641 B.n506 B.n89 163.367
R1642 B.n510 B.n89 163.367
R1643 B.n511 B.n510 163.367
R1644 B.n512 B.n511 163.367
R1645 B.n512 B.n87 163.367
R1646 B.n516 B.n87 163.367
R1647 B.n517 B.n516 163.367
R1648 B.n518 B.n517 163.367
R1649 B.n518 B.n85 163.367
R1650 B.n522 B.n85 163.367
R1651 B.n523 B.n522 163.367
R1652 B.n524 B.n523 163.367
R1653 B.n524 B.n83 163.367
R1654 B.n528 B.n83 163.367
R1655 B.n529 B.n528 163.367
R1656 B.n530 B.n529 163.367
R1657 B.n530 B.n81 163.367
R1658 B.n534 B.n81 163.367
R1659 B.n535 B.n534 163.367
R1660 B.n536 B.n535 163.367
R1661 B.n536 B.n79 163.367
R1662 B.n540 B.n79 163.367
R1663 B.n541 B.n540 163.367
R1664 B.n542 B.n541 163.367
R1665 B.n691 B.n690 163.367
R1666 B.n690 B.n25 163.367
R1667 B.n686 B.n25 163.367
R1668 B.n686 B.n685 163.367
R1669 B.n685 B.n684 163.367
R1670 B.n684 B.n27 163.367
R1671 B.n680 B.n27 163.367
R1672 B.n680 B.n679 163.367
R1673 B.n679 B.n678 163.367
R1674 B.n678 B.n29 163.367
R1675 B.n674 B.n29 163.367
R1676 B.n674 B.n673 163.367
R1677 B.n673 B.n672 163.367
R1678 B.n672 B.n31 163.367
R1679 B.n668 B.n31 163.367
R1680 B.n668 B.n667 163.367
R1681 B.n667 B.n666 163.367
R1682 B.n666 B.n33 163.367
R1683 B.n662 B.n33 163.367
R1684 B.n662 B.n661 163.367
R1685 B.n661 B.n660 163.367
R1686 B.n660 B.n35 163.367
R1687 B.n656 B.n35 163.367
R1688 B.n656 B.n655 163.367
R1689 B.n655 B.n654 163.367
R1690 B.n654 B.n37 163.367
R1691 B.n650 B.n37 163.367
R1692 B.n650 B.n649 163.367
R1693 B.n649 B.n648 163.367
R1694 B.n648 B.n39 163.367
R1695 B.n644 B.n39 163.367
R1696 B.n644 B.n643 163.367
R1697 B.n643 B.n642 163.367
R1698 B.n642 B.n41 163.367
R1699 B.n638 B.n41 163.367
R1700 B.n638 B.n637 163.367
R1701 B.n637 B.n636 163.367
R1702 B.n636 B.n43 163.367
R1703 B.n632 B.n43 163.367
R1704 B.n632 B.n631 163.367
R1705 B.n631 B.n630 163.367
R1706 B.n630 B.n45 163.367
R1707 B.n626 B.n45 163.367
R1708 B.n626 B.n625 163.367
R1709 B.n625 B.n49 163.367
R1710 B.n621 B.n49 163.367
R1711 B.n621 B.n620 163.367
R1712 B.n620 B.n619 163.367
R1713 B.n619 B.n51 163.367
R1714 B.n615 B.n51 163.367
R1715 B.n615 B.n614 163.367
R1716 B.n614 B.n613 163.367
R1717 B.n613 B.n53 163.367
R1718 B.n608 B.n53 163.367
R1719 B.n608 B.n607 163.367
R1720 B.n607 B.n606 163.367
R1721 B.n606 B.n57 163.367
R1722 B.n602 B.n57 163.367
R1723 B.n602 B.n601 163.367
R1724 B.n601 B.n600 163.367
R1725 B.n600 B.n59 163.367
R1726 B.n596 B.n59 163.367
R1727 B.n596 B.n595 163.367
R1728 B.n595 B.n594 163.367
R1729 B.n594 B.n61 163.367
R1730 B.n590 B.n61 163.367
R1731 B.n590 B.n589 163.367
R1732 B.n589 B.n588 163.367
R1733 B.n588 B.n63 163.367
R1734 B.n584 B.n63 163.367
R1735 B.n584 B.n583 163.367
R1736 B.n583 B.n582 163.367
R1737 B.n582 B.n65 163.367
R1738 B.n578 B.n65 163.367
R1739 B.n578 B.n577 163.367
R1740 B.n577 B.n576 163.367
R1741 B.n576 B.n67 163.367
R1742 B.n572 B.n67 163.367
R1743 B.n572 B.n571 163.367
R1744 B.n571 B.n570 163.367
R1745 B.n570 B.n69 163.367
R1746 B.n566 B.n69 163.367
R1747 B.n566 B.n565 163.367
R1748 B.n565 B.n564 163.367
R1749 B.n564 B.n71 163.367
R1750 B.n560 B.n71 163.367
R1751 B.n560 B.n559 163.367
R1752 B.n559 B.n558 163.367
R1753 B.n558 B.n73 163.367
R1754 B.n554 B.n73 163.367
R1755 B.n554 B.n553 163.367
R1756 B.n553 B.n552 163.367
R1757 B.n552 B.n75 163.367
R1758 B.n548 B.n75 163.367
R1759 B.n548 B.n547 163.367
R1760 B.n547 B.n546 163.367
R1761 B.n546 B.n77 163.367
R1762 B.n146 B.n145 59.5399
R1763 B.n328 B.n153 59.5399
R1764 B.n48 B.n47 59.5399
R1765 B.n610 B.n55 59.5399
R1766 B.n145 B.n144 59.346
R1767 B.n153 B.n152 59.346
R1768 B.n47 B.n46 59.346
R1769 B.n55 B.n54 59.346
R1770 B.n693 B.n24 34.1859
R1771 B.n544 B.n543 34.1859
R1772 B.n411 B.n122 34.1859
R1773 B.n262 B.n261 34.1859
R1774 B B.n759 18.0485
R1775 B.n689 B.n24 10.6151
R1776 B.n689 B.n688 10.6151
R1777 B.n688 B.n687 10.6151
R1778 B.n687 B.n26 10.6151
R1779 B.n683 B.n26 10.6151
R1780 B.n683 B.n682 10.6151
R1781 B.n682 B.n681 10.6151
R1782 B.n681 B.n28 10.6151
R1783 B.n677 B.n28 10.6151
R1784 B.n677 B.n676 10.6151
R1785 B.n676 B.n675 10.6151
R1786 B.n675 B.n30 10.6151
R1787 B.n671 B.n30 10.6151
R1788 B.n671 B.n670 10.6151
R1789 B.n670 B.n669 10.6151
R1790 B.n669 B.n32 10.6151
R1791 B.n665 B.n32 10.6151
R1792 B.n665 B.n664 10.6151
R1793 B.n664 B.n663 10.6151
R1794 B.n663 B.n34 10.6151
R1795 B.n659 B.n34 10.6151
R1796 B.n659 B.n658 10.6151
R1797 B.n658 B.n657 10.6151
R1798 B.n657 B.n36 10.6151
R1799 B.n653 B.n36 10.6151
R1800 B.n653 B.n652 10.6151
R1801 B.n652 B.n651 10.6151
R1802 B.n651 B.n38 10.6151
R1803 B.n647 B.n38 10.6151
R1804 B.n647 B.n646 10.6151
R1805 B.n646 B.n645 10.6151
R1806 B.n645 B.n40 10.6151
R1807 B.n641 B.n40 10.6151
R1808 B.n641 B.n640 10.6151
R1809 B.n640 B.n639 10.6151
R1810 B.n639 B.n42 10.6151
R1811 B.n635 B.n42 10.6151
R1812 B.n635 B.n634 10.6151
R1813 B.n634 B.n633 10.6151
R1814 B.n633 B.n44 10.6151
R1815 B.n629 B.n44 10.6151
R1816 B.n629 B.n628 10.6151
R1817 B.n628 B.n627 10.6151
R1818 B.n624 B.n623 10.6151
R1819 B.n623 B.n622 10.6151
R1820 B.n622 B.n50 10.6151
R1821 B.n618 B.n50 10.6151
R1822 B.n618 B.n617 10.6151
R1823 B.n617 B.n616 10.6151
R1824 B.n616 B.n52 10.6151
R1825 B.n612 B.n52 10.6151
R1826 B.n612 B.n611 10.6151
R1827 B.n609 B.n56 10.6151
R1828 B.n605 B.n56 10.6151
R1829 B.n605 B.n604 10.6151
R1830 B.n604 B.n603 10.6151
R1831 B.n603 B.n58 10.6151
R1832 B.n599 B.n58 10.6151
R1833 B.n599 B.n598 10.6151
R1834 B.n598 B.n597 10.6151
R1835 B.n597 B.n60 10.6151
R1836 B.n593 B.n60 10.6151
R1837 B.n593 B.n592 10.6151
R1838 B.n592 B.n591 10.6151
R1839 B.n591 B.n62 10.6151
R1840 B.n587 B.n62 10.6151
R1841 B.n587 B.n586 10.6151
R1842 B.n586 B.n585 10.6151
R1843 B.n585 B.n64 10.6151
R1844 B.n581 B.n64 10.6151
R1845 B.n581 B.n580 10.6151
R1846 B.n580 B.n579 10.6151
R1847 B.n579 B.n66 10.6151
R1848 B.n575 B.n66 10.6151
R1849 B.n575 B.n574 10.6151
R1850 B.n574 B.n573 10.6151
R1851 B.n573 B.n68 10.6151
R1852 B.n569 B.n68 10.6151
R1853 B.n569 B.n568 10.6151
R1854 B.n568 B.n567 10.6151
R1855 B.n567 B.n70 10.6151
R1856 B.n563 B.n70 10.6151
R1857 B.n563 B.n562 10.6151
R1858 B.n562 B.n561 10.6151
R1859 B.n561 B.n72 10.6151
R1860 B.n557 B.n72 10.6151
R1861 B.n557 B.n556 10.6151
R1862 B.n556 B.n555 10.6151
R1863 B.n555 B.n74 10.6151
R1864 B.n551 B.n74 10.6151
R1865 B.n551 B.n550 10.6151
R1866 B.n550 B.n549 10.6151
R1867 B.n549 B.n76 10.6151
R1868 B.n545 B.n76 10.6151
R1869 B.n545 B.n544 10.6151
R1870 B.n412 B.n411 10.6151
R1871 B.n413 B.n412 10.6151
R1872 B.n413 B.n120 10.6151
R1873 B.n417 B.n120 10.6151
R1874 B.n418 B.n417 10.6151
R1875 B.n419 B.n418 10.6151
R1876 B.n419 B.n118 10.6151
R1877 B.n423 B.n118 10.6151
R1878 B.n424 B.n423 10.6151
R1879 B.n425 B.n424 10.6151
R1880 B.n425 B.n116 10.6151
R1881 B.n429 B.n116 10.6151
R1882 B.n430 B.n429 10.6151
R1883 B.n431 B.n430 10.6151
R1884 B.n431 B.n114 10.6151
R1885 B.n435 B.n114 10.6151
R1886 B.n436 B.n435 10.6151
R1887 B.n437 B.n436 10.6151
R1888 B.n437 B.n112 10.6151
R1889 B.n441 B.n112 10.6151
R1890 B.n442 B.n441 10.6151
R1891 B.n443 B.n442 10.6151
R1892 B.n443 B.n110 10.6151
R1893 B.n447 B.n110 10.6151
R1894 B.n448 B.n447 10.6151
R1895 B.n449 B.n448 10.6151
R1896 B.n449 B.n108 10.6151
R1897 B.n453 B.n108 10.6151
R1898 B.n454 B.n453 10.6151
R1899 B.n455 B.n454 10.6151
R1900 B.n455 B.n106 10.6151
R1901 B.n459 B.n106 10.6151
R1902 B.n460 B.n459 10.6151
R1903 B.n461 B.n460 10.6151
R1904 B.n461 B.n104 10.6151
R1905 B.n465 B.n104 10.6151
R1906 B.n466 B.n465 10.6151
R1907 B.n467 B.n466 10.6151
R1908 B.n467 B.n102 10.6151
R1909 B.n471 B.n102 10.6151
R1910 B.n472 B.n471 10.6151
R1911 B.n473 B.n472 10.6151
R1912 B.n473 B.n100 10.6151
R1913 B.n477 B.n100 10.6151
R1914 B.n478 B.n477 10.6151
R1915 B.n479 B.n478 10.6151
R1916 B.n479 B.n98 10.6151
R1917 B.n483 B.n98 10.6151
R1918 B.n484 B.n483 10.6151
R1919 B.n485 B.n484 10.6151
R1920 B.n485 B.n96 10.6151
R1921 B.n489 B.n96 10.6151
R1922 B.n490 B.n489 10.6151
R1923 B.n491 B.n490 10.6151
R1924 B.n491 B.n94 10.6151
R1925 B.n495 B.n94 10.6151
R1926 B.n496 B.n495 10.6151
R1927 B.n497 B.n496 10.6151
R1928 B.n497 B.n92 10.6151
R1929 B.n501 B.n92 10.6151
R1930 B.n502 B.n501 10.6151
R1931 B.n503 B.n502 10.6151
R1932 B.n503 B.n90 10.6151
R1933 B.n507 B.n90 10.6151
R1934 B.n508 B.n507 10.6151
R1935 B.n509 B.n508 10.6151
R1936 B.n509 B.n88 10.6151
R1937 B.n513 B.n88 10.6151
R1938 B.n514 B.n513 10.6151
R1939 B.n515 B.n514 10.6151
R1940 B.n515 B.n86 10.6151
R1941 B.n519 B.n86 10.6151
R1942 B.n520 B.n519 10.6151
R1943 B.n521 B.n520 10.6151
R1944 B.n521 B.n84 10.6151
R1945 B.n525 B.n84 10.6151
R1946 B.n526 B.n525 10.6151
R1947 B.n527 B.n526 10.6151
R1948 B.n527 B.n82 10.6151
R1949 B.n531 B.n82 10.6151
R1950 B.n532 B.n531 10.6151
R1951 B.n533 B.n532 10.6151
R1952 B.n533 B.n80 10.6151
R1953 B.n537 B.n80 10.6151
R1954 B.n538 B.n537 10.6151
R1955 B.n539 B.n538 10.6151
R1956 B.n539 B.n78 10.6151
R1957 B.n543 B.n78 10.6151
R1958 B.n263 B.n262 10.6151
R1959 B.n263 B.n174 10.6151
R1960 B.n267 B.n174 10.6151
R1961 B.n268 B.n267 10.6151
R1962 B.n269 B.n268 10.6151
R1963 B.n269 B.n172 10.6151
R1964 B.n273 B.n172 10.6151
R1965 B.n274 B.n273 10.6151
R1966 B.n275 B.n274 10.6151
R1967 B.n275 B.n170 10.6151
R1968 B.n279 B.n170 10.6151
R1969 B.n280 B.n279 10.6151
R1970 B.n281 B.n280 10.6151
R1971 B.n281 B.n168 10.6151
R1972 B.n285 B.n168 10.6151
R1973 B.n286 B.n285 10.6151
R1974 B.n287 B.n286 10.6151
R1975 B.n287 B.n166 10.6151
R1976 B.n291 B.n166 10.6151
R1977 B.n292 B.n291 10.6151
R1978 B.n293 B.n292 10.6151
R1979 B.n293 B.n164 10.6151
R1980 B.n297 B.n164 10.6151
R1981 B.n298 B.n297 10.6151
R1982 B.n299 B.n298 10.6151
R1983 B.n299 B.n162 10.6151
R1984 B.n303 B.n162 10.6151
R1985 B.n304 B.n303 10.6151
R1986 B.n305 B.n304 10.6151
R1987 B.n305 B.n160 10.6151
R1988 B.n309 B.n160 10.6151
R1989 B.n310 B.n309 10.6151
R1990 B.n311 B.n310 10.6151
R1991 B.n311 B.n158 10.6151
R1992 B.n315 B.n158 10.6151
R1993 B.n316 B.n315 10.6151
R1994 B.n317 B.n316 10.6151
R1995 B.n317 B.n156 10.6151
R1996 B.n321 B.n156 10.6151
R1997 B.n322 B.n321 10.6151
R1998 B.n323 B.n322 10.6151
R1999 B.n323 B.n154 10.6151
R2000 B.n327 B.n154 10.6151
R2001 B.n330 B.n329 10.6151
R2002 B.n330 B.n150 10.6151
R2003 B.n334 B.n150 10.6151
R2004 B.n335 B.n334 10.6151
R2005 B.n336 B.n335 10.6151
R2006 B.n336 B.n148 10.6151
R2007 B.n340 B.n148 10.6151
R2008 B.n341 B.n340 10.6151
R2009 B.n342 B.n341 10.6151
R2010 B.n346 B.n345 10.6151
R2011 B.n347 B.n346 10.6151
R2012 B.n347 B.n142 10.6151
R2013 B.n351 B.n142 10.6151
R2014 B.n352 B.n351 10.6151
R2015 B.n353 B.n352 10.6151
R2016 B.n353 B.n140 10.6151
R2017 B.n357 B.n140 10.6151
R2018 B.n358 B.n357 10.6151
R2019 B.n359 B.n358 10.6151
R2020 B.n359 B.n138 10.6151
R2021 B.n363 B.n138 10.6151
R2022 B.n364 B.n363 10.6151
R2023 B.n365 B.n364 10.6151
R2024 B.n365 B.n136 10.6151
R2025 B.n369 B.n136 10.6151
R2026 B.n370 B.n369 10.6151
R2027 B.n371 B.n370 10.6151
R2028 B.n371 B.n134 10.6151
R2029 B.n375 B.n134 10.6151
R2030 B.n376 B.n375 10.6151
R2031 B.n377 B.n376 10.6151
R2032 B.n377 B.n132 10.6151
R2033 B.n381 B.n132 10.6151
R2034 B.n382 B.n381 10.6151
R2035 B.n383 B.n382 10.6151
R2036 B.n383 B.n130 10.6151
R2037 B.n387 B.n130 10.6151
R2038 B.n388 B.n387 10.6151
R2039 B.n389 B.n388 10.6151
R2040 B.n389 B.n128 10.6151
R2041 B.n393 B.n128 10.6151
R2042 B.n394 B.n393 10.6151
R2043 B.n395 B.n394 10.6151
R2044 B.n395 B.n126 10.6151
R2045 B.n399 B.n126 10.6151
R2046 B.n400 B.n399 10.6151
R2047 B.n401 B.n400 10.6151
R2048 B.n401 B.n124 10.6151
R2049 B.n405 B.n124 10.6151
R2050 B.n406 B.n405 10.6151
R2051 B.n407 B.n406 10.6151
R2052 B.n407 B.n122 10.6151
R2053 B.n261 B.n176 10.6151
R2054 B.n257 B.n176 10.6151
R2055 B.n257 B.n256 10.6151
R2056 B.n256 B.n255 10.6151
R2057 B.n255 B.n178 10.6151
R2058 B.n251 B.n178 10.6151
R2059 B.n251 B.n250 10.6151
R2060 B.n250 B.n249 10.6151
R2061 B.n249 B.n180 10.6151
R2062 B.n245 B.n180 10.6151
R2063 B.n245 B.n244 10.6151
R2064 B.n244 B.n243 10.6151
R2065 B.n243 B.n182 10.6151
R2066 B.n239 B.n182 10.6151
R2067 B.n239 B.n238 10.6151
R2068 B.n238 B.n237 10.6151
R2069 B.n237 B.n184 10.6151
R2070 B.n233 B.n184 10.6151
R2071 B.n233 B.n232 10.6151
R2072 B.n232 B.n231 10.6151
R2073 B.n231 B.n186 10.6151
R2074 B.n227 B.n186 10.6151
R2075 B.n227 B.n226 10.6151
R2076 B.n226 B.n225 10.6151
R2077 B.n225 B.n188 10.6151
R2078 B.n221 B.n188 10.6151
R2079 B.n221 B.n220 10.6151
R2080 B.n220 B.n219 10.6151
R2081 B.n219 B.n190 10.6151
R2082 B.n215 B.n190 10.6151
R2083 B.n215 B.n214 10.6151
R2084 B.n214 B.n213 10.6151
R2085 B.n213 B.n192 10.6151
R2086 B.n209 B.n192 10.6151
R2087 B.n209 B.n208 10.6151
R2088 B.n208 B.n207 10.6151
R2089 B.n207 B.n194 10.6151
R2090 B.n203 B.n194 10.6151
R2091 B.n203 B.n202 10.6151
R2092 B.n202 B.n201 10.6151
R2093 B.n201 B.n196 10.6151
R2094 B.n197 B.n196 10.6151
R2095 B.n197 B.n0 10.6151
R2096 B.n755 B.n1 10.6151
R2097 B.n755 B.n754 10.6151
R2098 B.n754 B.n753 10.6151
R2099 B.n753 B.n4 10.6151
R2100 B.n749 B.n4 10.6151
R2101 B.n749 B.n748 10.6151
R2102 B.n748 B.n747 10.6151
R2103 B.n747 B.n6 10.6151
R2104 B.n743 B.n6 10.6151
R2105 B.n743 B.n742 10.6151
R2106 B.n742 B.n741 10.6151
R2107 B.n741 B.n8 10.6151
R2108 B.n737 B.n8 10.6151
R2109 B.n737 B.n736 10.6151
R2110 B.n736 B.n735 10.6151
R2111 B.n735 B.n10 10.6151
R2112 B.n731 B.n10 10.6151
R2113 B.n731 B.n730 10.6151
R2114 B.n730 B.n729 10.6151
R2115 B.n729 B.n12 10.6151
R2116 B.n725 B.n12 10.6151
R2117 B.n725 B.n724 10.6151
R2118 B.n724 B.n723 10.6151
R2119 B.n723 B.n14 10.6151
R2120 B.n719 B.n14 10.6151
R2121 B.n719 B.n718 10.6151
R2122 B.n718 B.n717 10.6151
R2123 B.n717 B.n16 10.6151
R2124 B.n713 B.n16 10.6151
R2125 B.n713 B.n712 10.6151
R2126 B.n712 B.n711 10.6151
R2127 B.n711 B.n18 10.6151
R2128 B.n707 B.n18 10.6151
R2129 B.n707 B.n706 10.6151
R2130 B.n706 B.n705 10.6151
R2131 B.n705 B.n20 10.6151
R2132 B.n701 B.n20 10.6151
R2133 B.n701 B.n700 10.6151
R2134 B.n700 B.n699 10.6151
R2135 B.n699 B.n22 10.6151
R2136 B.n695 B.n22 10.6151
R2137 B.n695 B.n694 10.6151
R2138 B.n694 B.n693 10.6151
R2139 B.n627 B.n48 9.36635
R2140 B.n610 B.n609 9.36635
R2141 B.n328 B.n327 9.36635
R2142 B.n345 B.n146 9.36635
R2143 B.n759 B.n0 2.81026
R2144 B.n759 B.n1 2.81026
R2145 B.n624 B.n48 1.24928
R2146 B.n611 B.n610 1.24928
R2147 B.n329 B.n328 1.24928
R2148 B.n342 B.n146 1.24928
C0 w_n3418_n3548# VDD2 2.47186f
C1 VDD1 VTAIL 8.075971f
C2 VDD2 VTAIL 8.12761f
C3 VDD1 VN 0.150419f
C4 VN VDD2 7.26892f
C5 VDD1 VDD2 1.45661f
C6 VP B 1.94028f
C7 VP w_n3418_n3548# 6.98068f
C8 VP VTAIL 7.42885f
C9 VN VP 7.22638f
C10 w_n3418_n3548# B 10.1081f
C11 VDD1 VP 7.58411f
C12 VP VDD2 0.468911f
C13 VTAIL B 3.95012f
C14 VN B 1.20122f
C15 w_n3418_n3548# VTAIL 3.10505f
C16 VN w_n3418_n3548# 6.53842f
C17 VN VTAIL 7.41456f
C18 VDD1 B 2.19839f
C19 VDD2 B 2.2756f
C20 VDD1 w_n3418_n3548# 2.38266f
C21 VDD2 VSUBS 1.975858f
C22 VDD1 VSUBS 1.904109f
C23 VTAIL VSUBS 1.242275f
C24 VN VSUBS 5.969269f
C25 VP VSUBS 3.058545f
C26 B VSUBS 4.843148f
C27 w_n3418_n3548# VSUBS 0.149093p
C28 B.n0 VSUBS 0.004965f
C29 B.n1 VSUBS 0.004965f
C30 B.n2 VSUBS 0.007852f
C31 B.n3 VSUBS 0.007852f
C32 B.n4 VSUBS 0.007852f
C33 B.n5 VSUBS 0.007852f
C34 B.n6 VSUBS 0.007852f
C35 B.n7 VSUBS 0.007852f
C36 B.n8 VSUBS 0.007852f
C37 B.n9 VSUBS 0.007852f
C38 B.n10 VSUBS 0.007852f
C39 B.n11 VSUBS 0.007852f
C40 B.n12 VSUBS 0.007852f
C41 B.n13 VSUBS 0.007852f
C42 B.n14 VSUBS 0.007852f
C43 B.n15 VSUBS 0.007852f
C44 B.n16 VSUBS 0.007852f
C45 B.n17 VSUBS 0.007852f
C46 B.n18 VSUBS 0.007852f
C47 B.n19 VSUBS 0.007852f
C48 B.n20 VSUBS 0.007852f
C49 B.n21 VSUBS 0.007852f
C50 B.n22 VSUBS 0.007852f
C51 B.n23 VSUBS 0.007852f
C52 B.n24 VSUBS 0.019402f
C53 B.n25 VSUBS 0.007852f
C54 B.n26 VSUBS 0.007852f
C55 B.n27 VSUBS 0.007852f
C56 B.n28 VSUBS 0.007852f
C57 B.n29 VSUBS 0.007852f
C58 B.n30 VSUBS 0.007852f
C59 B.n31 VSUBS 0.007852f
C60 B.n32 VSUBS 0.007852f
C61 B.n33 VSUBS 0.007852f
C62 B.n34 VSUBS 0.007852f
C63 B.n35 VSUBS 0.007852f
C64 B.n36 VSUBS 0.007852f
C65 B.n37 VSUBS 0.007852f
C66 B.n38 VSUBS 0.007852f
C67 B.n39 VSUBS 0.007852f
C68 B.n40 VSUBS 0.007852f
C69 B.n41 VSUBS 0.007852f
C70 B.n42 VSUBS 0.007852f
C71 B.n43 VSUBS 0.007852f
C72 B.n44 VSUBS 0.007852f
C73 B.n45 VSUBS 0.007852f
C74 B.t8 VSUBS 0.259635f
C75 B.t7 VSUBS 0.297165f
C76 B.t6 VSUBS 1.79715f
C77 B.n46 VSUBS 0.46898f
C78 B.n47 VSUBS 0.296652f
C79 B.n48 VSUBS 0.018192f
C80 B.n49 VSUBS 0.007852f
C81 B.n50 VSUBS 0.007852f
C82 B.n51 VSUBS 0.007852f
C83 B.n52 VSUBS 0.007852f
C84 B.n53 VSUBS 0.007852f
C85 B.t5 VSUBS 0.259639f
C86 B.t4 VSUBS 0.297168f
C87 B.t3 VSUBS 1.79715f
C88 B.n54 VSUBS 0.468977f
C89 B.n55 VSUBS 0.296649f
C90 B.n56 VSUBS 0.007852f
C91 B.n57 VSUBS 0.007852f
C92 B.n58 VSUBS 0.007852f
C93 B.n59 VSUBS 0.007852f
C94 B.n60 VSUBS 0.007852f
C95 B.n61 VSUBS 0.007852f
C96 B.n62 VSUBS 0.007852f
C97 B.n63 VSUBS 0.007852f
C98 B.n64 VSUBS 0.007852f
C99 B.n65 VSUBS 0.007852f
C100 B.n66 VSUBS 0.007852f
C101 B.n67 VSUBS 0.007852f
C102 B.n68 VSUBS 0.007852f
C103 B.n69 VSUBS 0.007852f
C104 B.n70 VSUBS 0.007852f
C105 B.n71 VSUBS 0.007852f
C106 B.n72 VSUBS 0.007852f
C107 B.n73 VSUBS 0.007852f
C108 B.n74 VSUBS 0.007852f
C109 B.n75 VSUBS 0.007852f
C110 B.n76 VSUBS 0.007852f
C111 B.n77 VSUBS 0.019402f
C112 B.n78 VSUBS 0.007852f
C113 B.n79 VSUBS 0.007852f
C114 B.n80 VSUBS 0.007852f
C115 B.n81 VSUBS 0.007852f
C116 B.n82 VSUBS 0.007852f
C117 B.n83 VSUBS 0.007852f
C118 B.n84 VSUBS 0.007852f
C119 B.n85 VSUBS 0.007852f
C120 B.n86 VSUBS 0.007852f
C121 B.n87 VSUBS 0.007852f
C122 B.n88 VSUBS 0.007852f
C123 B.n89 VSUBS 0.007852f
C124 B.n90 VSUBS 0.007852f
C125 B.n91 VSUBS 0.007852f
C126 B.n92 VSUBS 0.007852f
C127 B.n93 VSUBS 0.007852f
C128 B.n94 VSUBS 0.007852f
C129 B.n95 VSUBS 0.007852f
C130 B.n96 VSUBS 0.007852f
C131 B.n97 VSUBS 0.007852f
C132 B.n98 VSUBS 0.007852f
C133 B.n99 VSUBS 0.007852f
C134 B.n100 VSUBS 0.007852f
C135 B.n101 VSUBS 0.007852f
C136 B.n102 VSUBS 0.007852f
C137 B.n103 VSUBS 0.007852f
C138 B.n104 VSUBS 0.007852f
C139 B.n105 VSUBS 0.007852f
C140 B.n106 VSUBS 0.007852f
C141 B.n107 VSUBS 0.007852f
C142 B.n108 VSUBS 0.007852f
C143 B.n109 VSUBS 0.007852f
C144 B.n110 VSUBS 0.007852f
C145 B.n111 VSUBS 0.007852f
C146 B.n112 VSUBS 0.007852f
C147 B.n113 VSUBS 0.007852f
C148 B.n114 VSUBS 0.007852f
C149 B.n115 VSUBS 0.007852f
C150 B.n116 VSUBS 0.007852f
C151 B.n117 VSUBS 0.007852f
C152 B.n118 VSUBS 0.007852f
C153 B.n119 VSUBS 0.007852f
C154 B.n120 VSUBS 0.007852f
C155 B.n121 VSUBS 0.007852f
C156 B.n122 VSUBS 0.019402f
C157 B.n123 VSUBS 0.007852f
C158 B.n124 VSUBS 0.007852f
C159 B.n125 VSUBS 0.007852f
C160 B.n126 VSUBS 0.007852f
C161 B.n127 VSUBS 0.007852f
C162 B.n128 VSUBS 0.007852f
C163 B.n129 VSUBS 0.007852f
C164 B.n130 VSUBS 0.007852f
C165 B.n131 VSUBS 0.007852f
C166 B.n132 VSUBS 0.007852f
C167 B.n133 VSUBS 0.007852f
C168 B.n134 VSUBS 0.007852f
C169 B.n135 VSUBS 0.007852f
C170 B.n136 VSUBS 0.007852f
C171 B.n137 VSUBS 0.007852f
C172 B.n138 VSUBS 0.007852f
C173 B.n139 VSUBS 0.007852f
C174 B.n140 VSUBS 0.007852f
C175 B.n141 VSUBS 0.007852f
C176 B.n142 VSUBS 0.007852f
C177 B.n143 VSUBS 0.007852f
C178 B.t10 VSUBS 0.259639f
C179 B.t11 VSUBS 0.297168f
C180 B.t9 VSUBS 1.79715f
C181 B.n144 VSUBS 0.468977f
C182 B.n145 VSUBS 0.296649f
C183 B.n146 VSUBS 0.018192f
C184 B.n147 VSUBS 0.007852f
C185 B.n148 VSUBS 0.007852f
C186 B.n149 VSUBS 0.007852f
C187 B.n150 VSUBS 0.007852f
C188 B.n151 VSUBS 0.007852f
C189 B.t1 VSUBS 0.259635f
C190 B.t2 VSUBS 0.297165f
C191 B.t0 VSUBS 1.79715f
C192 B.n152 VSUBS 0.46898f
C193 B.n153 VSUBS 0.296652f
C194 B.n154 VSUBS 0.007852f
C195 B.n155 VSUBS 0.007852f
C196 B.n156 VSUBS 0.007852f
C197 B.n157 VSUBS 0.007852f
C198 B.n158 VSUBS 0.007852f
C199 B.n159 VSUBS 0.007852f
C200 B.n160 VSUBS 0.007852f
C201 B.n161 VSUBS 0.007852f
C202 B.n162 VSUBS 0.007852f
C203 B.n163 VSUBS 0.007852f
C204 B.n164 VSUBS 0.007852f
C205 B.n165 VSUBS 0.007852f
C206 B.n166 VSUBS 0.007852f
C207 B.n167 VSUBS 0.007852f
C208 B.n168 VSUBS 0.007852f
C209 B.n169 VSUBS 0.007852f
C210 B.n170 VSUBS 0.007852f
C211 B.n171 VSUBS 0.007852f
C212 B.n172 VSUBS 0.007852f
C213 B.n173 VSUBS 0.007852f
C214 B.n174 VSUBS 0.007852f
C215 B.n175 VSUBS 0.019402f
C216 B.n176 VSUBS 0.007852f
C217 B.n177 VSUBS 0.007852f
C218 B.n178 VSUBS 0.007852f
C219 B.n179 VSUBS 0.007852f
C220 B.n180 VSUBS 0.007852f
C221 B.n181 VSUBS 0.007852f
C222 B.n182 VSUBS 0.007852f
C223 B.n183 VSUBS 0.007852f
C224 B.n184 VSUBS 0.007852f
C225 B.n185 VSUBS 0.007852f
C226 B.n186 VSUBS 0.007852f
C227 B.n187 VSUBS 0.007852f
C228 B.n188 VSUBS 0.007852f
C229 B.n189 VSUBS 0.007852f
C230 B.n190 VSUBS 0.007852f
C231 B.n191 VSUBS 0.007852f
C232 B.n192 VSUBS 0.007852f
C233 B.n193 VSUBS 0.007852f
C234 B.n194 VSUBS 0.007852f
C235 B.n195 VSUBS 0.007852f
C236 B.n196 VSUBS 0.007852f
C237 B.n197 VSUBS 0.007852f
C238 B.n198 VSUBS 0.007852f
C239 B.n199 VSUBS 0.007852f
C240 B.n200 VSUBS 0.007852f
C241 B.n201 VSUBS 0.007852f
C242 B.n202 VSUBS 0.007852f
C243 B.n203 VSUBS 0.007852f
C244 B.n204 VSUBS 0.007852f
C245 B.n205 VSUBS 0.007852f
C246 B.n206 VSUBS 0.007852f
C247 B.n207 VSUBS 0.007852f
C248 B.n208 VSUBS 0.007852f
C249 B.n209 VSUBS 0.007852f
C250 B.n210 VSUBS 0.007852f
C251 B.n211 VSUBS 0.007852f
C252 B.n212 VSUBS 0.007852f
C253 B.n213 VSUBS 0.007852f
C254 B.n214 VSUBS 0.007852f
C255 B.n215 VSUBS 0.007852f
C256 B.n216 VSUBS 0.007852f
C257 B.n217 VSUBS 0.007852f
C258 B.n218 VSUBS 0.007852f
C259 B.n219 VSUBS 0.007852f
C260 B.n220 VSUBS 0.007852f
C261 B.n221 VSUBS 0.007852f
C262 B.n222 VSUBS 0.007852f
C263 B.n223 VSUBS 0.007852f
C264 B.n224 VSUBS 0.007852f
C265 B.n225 VSUBS 0.007852f
C266 B.n226 VSUBS 0.007852f
C267 B.n227 VSUBS 0.007852f
C268 B.n228 VSUBS 0.007852f
C269 B.n229 VSUBS 0.007852f
C270 B.n230 VSUBS 0.007852f
C271 B.n231 VSUBS 0.007852f
C272 B.n232 VSUBS 0.007852f
C273 B.n233 VSUBS 0.007852f
C274 B.n234 VSUBS 0.007852f
C275 B.n235 VSUBS 0.007852f
C276 B.n236 VSUBS 0.007852f
C277 B.n237 VSUBS 0.007852f
C278 B.n238 VSUBS 0.007852f
C279 B.n239 VSUBS 0.007852f
C280 B.n240 VSUBS 0.007852f
C281 B.n241 VSUBS 0.007852f
C282 B.n242 VSUBS 0.007852f
C283 B.n243 VSUBS 0.007852f
C284 B.n244 VSUBS 0.007852f
C285 B.n245 VSUBS 0.007852f
C286 B.n246 VSUBS 0.007852f
C287 B.n247 VSUBS 0.007852f
C288 B.n248 VSUBS 0.007852f
C289 B.n249 VSUBS 0.007852f
C290 B.n250 VSUBS 0.007852f
C291 B.n251 VSUBS 0.007852f
C292 B.n252 VSUBS 0.007852f
C293 B.n253 VSUBS 0.007852f
C294 B.n254 VSUBS 0.007852f
C295 B.n255 VSUBS 0.007852f
C296 B.n256 VSUBS 0.007852f
C297 B.n257 VSUBS 0.007852f
C298 B.n258 VSUBS 0.007852f
C299 B.n259 VSUBS 0.007852f
C300 B.n260 VSUBS 0.018472f
C301 B.n261 VSUBS 0.018472f
C302 B.n262 VSUBS 0.019402f
C303 B.n263 VSUBS 0.007852f
C304 B.n264 VSUBS 0.007852f
C305 B.n265 VSUBS 0.007852f
C306 B.n266 VSUBS 0.007852f
C307 B.n267 VSUBS 0.007852f
C308 B.n268 VSUBS 0.007852f
C309 B.n269 VSUBS 0.007852f
C310 B.n270 VSUBS 0.007852f
C311 B.n271 VSUBS 0.007852f
C312 B.n272 VSUBS 0.007852f
C313 B.n273 VSUBS 0.007852f
C314 B.n274 VSUBS 0.007852f
C315 B.n275 VSUBS 0.007852f
C316 B.n276 VSUBS 0.007852f
C317 B.n277 VSUBS 0.007852f
C318 B.n278 VSUBS 0.007852f
C319 B.n279 VSUBS 0.007852f
C320 B.n280 VSUBS 0.007852f
C321 B.n281 VSUBS 0.007852f
C322 B.n282 VSUBS 0.007852f
C323 B.n283 VSUBS 0.007852f
C324 B.n284 VSUBS 0.007852f
C325 B.n285 VSUBS 0.007852f
C326 B.n286 VSUBS 0.007852f
C327 B.n287 VSUBS 0.007852f
C328 B.n288 VSUBS 0.007852f
C329 B.n289 VSUBS 0.007852f
C330 B.n290 VSUBS 0.007852f
C331 B.n291 VSUBS 0.007852f
C332 B.n292 VSUBS 0.007852f
C333 B.n293 VSUBS 0.007852f
C334 B.n294 VSUBS 0.007852f
C335 B.n295 VSUBS 0.007852f
C336 B.n296 VSUBS 0.007852f
C337 B.n297 VSUBS 0.007852f
C338 B.n298 VSUBS 0.007852f
C339 B.n299 VSUBS 0.007852f
C340 B.n300 VSUBS 0.007852f
C341 B.n301 VSUBS 0.007852f
C342 B.n302 VSUBS 0.007852f
C343 B.n303 VSUBS 0.007852f
C344 B.n304 VSUBS 0.007852f
C345 B.n305 VSUBS 0.007852f
C346 B.n306 VSUBS 0.007852f
C347 B.n307 VSUBS 0.007852f
C348 B.n308 VSUBS 0.007852f
C349 B.n309 VSUBS 0.007852f
C350 B.n310 VSUBS 0.007852f
C351 B.n311 VSUBS 0.007852f
C352 B.n312 VSUBS 0.007852f
C353 B.n313 VSUBS 0.007852f
C354 B.n314 VSUBS 0.007852f
C355 B.n315 VSUBS 0.007852f
C356 B.n316 VSUBS 0.007852f
C357 B.n317 VSUBS 0.007852f
C358 B.n318 VSUBS 0.007852f
C359 B.n319 VSUBS 0.007852f
C360 B.n320 VSUBS 0.007852f
C361 B.n321 VSUBS 0.007852f
C362 B.n322 VSUBS 0.007852f
C363 B.n323 VSUBS 0.007852f
C364 B.n324 VSUBS 0.007852f
C365 B.n325 VSUBS 0.007852f
C366 B.n326 VSUBS 0.007852f
C367 B.n327 VSUBS 0.00739f
C368 B.n328 VSUBS 0.018192f
C369 B.n329 VSUBS 0.004388f
C370 B.n330 VSUBS 0.007852f
C371 B.n331 VSUBS 0.007852f
C372 B.n332 VSUBS 0.007852f
C373 B.n333 VSUBS 0.007852f
C374 B.n334 VSUBS 0.007852f
C375 B.n335 VSUBS 0.007852f
C376 B.n336 VSUBS 0.007852f
C377 B.n337 VSUBS 0.007852f
C378 B.n338 VSUBS 0.007852f
C379 B.n339 VSUBS 0.007852f
C380 B.n340 VSUBS 0.007852f
C381 B.n341 VSUBS 0.007852f
C382 B.n342 VSUBS 0.004388f
C383 B.n343 VSUBS 0.007852f
C384 B.n344 VSUBS 0.007852f
C385 B.n345 VSUBS 0.00739f
C386 B.n346 VSUBS 0.007852f
C387 B.n347 VSUBS 0.007852f
C388 B.n348 VSUBS 0.007852f
C389 B.n349 VSUBS 0.007852f
C390 B.n350 VSUBS 0.007852f
C391 B.n351 VSUBS 0.007852f
C392 B.n352 VSUBS 0.007852f
C393 B.n353 VSUBS 0.007852f
C394 B.n354 VSUBS 0.007852f
C395 B.n355 VSUBS 0.007852f
C396 B.n356 VSUBS 0.007852f
C397 B.n357 VSUBS 0.007852f
C398 B.n358 VSUBS 0.007852f
C399 B.n359 VSUBS 0.007852f
C400 B.n360 VSUBS 0.007852f
C401 B.n361 VSUBS 0.007852f
C402 B.n362 VSUBS 0.007852f
C403 B.n363 VSUBS 0.007852f
C404 B.n364 VSUBS 0.007852f
C405 B.n365 VSUBS 0.007852f
C406 B.n366 VSUBS 0.007852f
C407 B.n367 VSUBS 0.007852f
C408 B.n368 VSUBS 0.007852f
C409 B.n369 VSUBS 0.007852f
C410 B.n370 VSUBS 0.007852f
C411 B.n371 VSUBS 0.007852f
C412 B.n372 VSUBS 0.007852f
C413 B.n373 VSUBS 0.007852f
C414 B.n374 VSUBS 0.007852f
C415 B.n375 VSUBS 0.007852f
C416 B.n376 VSUBS 0.007852f
C417 B.n377 VSUBS 0.007852f
C418 B.n378 VSUBS 0.007852f
C419 B.n379 VSUBS 0.007852f
C420 B.n380 VSUBS 0.007852f
C421 B.n381 VSUBS 0.007852f
C422 B.n382 VSUBS 0.007852f
C423 B.n383 VSUBS 0.007852f
C424 B.n384 VSUBS 0.007852f
C425 B.n385 VSUBS 0.007852f
C426 B.n386 VSUBS 0.007852f
C427 B.n387 VSUBS 0.007852f
C428 B.n388 VSUBS 0.007852f
C429 B.n389 VSUBS 0.007852f
C430 B.n390 VSUBS 0.007852f
C431 B.n391 VSUBS 0.007852f
C432 B.n392 VSUBS 0.007852f
C433 B.n393 VSUBS 0.007852f
C434 B.n394 VSUBS 0.007852f
C435 B.n395 VSUBS 0.007852f
C436 B.n396 VSUBS 0.007852f
C437 B.n397 VSUBS 0.007852f
C438 B.n398 VSUBS 0.007852f
C439 B.n399 VSUBS 0.007852f
C440 B.n400 VSUBS 0.007852f
C441 B.n401 VSUBS 0.007852f
C442 B.n402 VSUBS 0.007852f
C443 B.n403 VSUBS 0.007852f
C444 B.n404 VSUBS 0.007852f
C445 B.n405 VSUBS 0.007852f
C446 B.n406 VSUBS 0.007852f
C447 B.n407 VSUBS 0.007852f
C448 B.n408 VSUBS 0.007852f
C449 B.n409 VSUBS 0.019402f
C450 B.n410 VSUBS 0.018472f
C451 B.n411 VSUBS 0.018472f
C452 B.n412 VSUBS 0.007852f
C453 B.n413 VSUBS 0.007852f
C454 B.n414 VSUBS 0.007852f
C455 B.n415 VSUBS 0.007852f
C456 B.n416 VSUBS 0.007852f
C457 B.n417 VSUBS 0.007852f
C458 B.n418 VSUBS 0.007852f
C459 B.n419 VSUBS 0.007852f
C460 B.n420 VSUBS 0.007852f
C461 B.n421 VSUBS 0.007852f
C462 B.n422 VSUBS 0.007852f
C463 B.n423 VSUBS 0.007852f
C464 B.n424 VSUBS 0.007852f
C465 B.n425 VSUBS 0.007852f
C466 B.n426 VSUBS 0.007852f
C467 B.n427 VSUBS 0.007852f
C468 B.n428 VSUBS 0.007852f
C469 B.n429 VSUBS 0.007852f
C470 B.n430 VSUBS 0.007852f
C471 B.n431 VSUBS 0.007852f
C472 B.n432 VSUBS 0.007852f
C473 B.n433 VSUBS 0.007852f
C474 B.n434 VSUBS 0.007852f
C475 B.n435 VSUBS 0.007852f
C476 B.n436 VSUBS 0.007852f
C477 B.n437 VSUBS 0.007852f
C478 B.n438 VSUBS 0.007852f
C479 B.n439 VSUBS 0.007852f
C480 B.n440 VSUBS 0.007852f
C481 B.n441 VSUBS 0.007852f
C482 B.n442 VSUBS 0.007852f
C483 B.n443 VSUBS 0.007852f
C484 B.n444 VSUBS 0.007852f
C485 B.n445 VSUBS 0.007852f
C486 B.n446 VSUBS 0.007852f
C487 B.n447 VSUBS 0.007852f
C488 B.n448 VSUBS 0.007852f
C489 B.n449 VSUBS 0.007852f
C490 B.n450 VSUBS 0.007852f
C491 B.n451 VSUBS 0.007852f
C492 B.n452 VSUBS 0.007852f
C493 B.n453 VSUBS 0.007852f
C494 B.n454 VSUBS 0.007852f
C495 B.n455 VSUBS 0.007852f
C496 B.n456 VSUBS 0.007852f
C497 B.n457 VSUBS 0.007852f
C498 B.n458 VSUBS 0.007852f
C499 B.n459 VSUBS 0.007852f
C500 B.n460 VSUBS 0.007852f
C501 B.n461 VSUBS 0.007852f
C502 B.n462 VSUBS 0.007852f
C503 B.n463 VSUBS 0.007852f
C504 B.n464 VSUBS 0.007852f
C505 B.n465 VSUBS 0.007852f
C506 B.n466 VSUBS 0.007852f
C507 B.n467 VSUBS 0.007852f
C508 B.n468 VSUBS 0.007852f
C509 B.n469 VSUBS 0.007852f
C510 B.n470 VSUBS 0.007852f
C511 B.n471 VSUBS 0.007852f
C512 B.n472 VSUBS 0.007852f
C513 B.n473 VSUBS 0.007852f
C514 B.n474 VSUBS 0.007852f
C515 B.n475 VSUBS 0.007852f
C516 B.n476 VSUBS 0.007852f
C517 B.n477 VSUBS 0.007852f
C518 B.n478 VSUBS 0.007852f
C519 B.n479 VSUBS 0.007852f
C520 B.n480 VSUBS 0.007852f
C521 B.n481 VSUBS 0.007852f
C522 B.n482 VSUBS 0.007852f
C523 B.n483 VSUBS 0.007852f
C524 B.n484 VSUBS 0.007852f
C525 B.n485 VSUBS 0.007852f
C526 B.n486 VSUBS 0.007852f
C527 B.n487 VSUBS 0.007852f
C528 B.n488 VSUBS 0.007852f
C529 B.n489 VSUBS 0.007852f
C530 B.n490 VSUBS 0.007852f
C531 B.n491 VSUBS 0.007852f
C532 B.n492 VSUBS 0.007852f
C533 B.n493 VSUBS 0.007852f
C534 B.n494 VSUBS 0.007852f
C535 B.n495 VSUBS 0.007852f
C536 B.n496 VSUBS 0.007852f
C537 B.n497 VSUBS 0.007852f
C538 B.n498 VSUBS 0.007852f
C539 B.n499 VSUBS 0.007852f
C540 B.n500 VSUBS 0.007852f
C541 B.n501 VSUBS 0.007852f
C542 B.n502 VSUBS 0.007852f
C543 B.n503 VSUBS 0.007852f
C544 B.n504 VSUBS 0.007852f
C545 B.n505 VSUBS 0.007852f
C546 B.n506 VSUBS 0.007852f
C547 B.n507 VSUBS 0.007852f
C548 B.n508 VSUBS 0.007852f
C549 B.n509 VSUBS 0.007852f
C550 B.n510 VSUBS 0.007852f
C551 B.n511 VSUBS 0.007852f
C552 B.n512 VSUBS 0.007852f
C553 B.n513 VSUBS 0.007852f
C554 B.n514 VSUBS 0.007852f
C555 B.n515 VSUBS 0.007852f
C556 B.n516 VSUBS 0.007852f
C557 B.n517 VSUBS 0.007852f
C558 B.n518 VSUBS 0.007852f
C559 B.n519 VSUBS 0.007852f
C560 B.n520 VSUBS 0.007852f
C561 B.n521 VSUBS 0.007852f
C562 B.n522 VSUBS 0.007852f
C563 B.n523 VSUBS 0.007852f
C564 B.n524 VSUBS 0.007852f
C565 B.n525 VSUBS 0.007852f
C566 B.n526 VSUBS 0.007852f
C567 B.n527 VSUBS 0.007852f
C568 B.n528 VSUBS 0.007852f
C569 B.n529 VSUBS 0.007852f
C570 B.n530 VSUBS 0.007852f
C571 B.n531 VSUBS 0.007852f
C572 B.n532 VSUBS 0.007852f
C573 B.n533 VSUBS 0.007852f
C574 B.n534 VSUBS 0.007852f
C575 B.n535 VSUBS 0.007852f
C576 B.n536 VSUBS 0.007852f
C577 B.n537 VSUBS 0.007852f
C578 B.n538 VSUBS 0.007852f
C579 B.n539 VSUBS 0.007852f
C580 B.n540 VSUBS 0.007852f
C581 B.n541 VSUBS 0.007852f
C582 B.n542 VSUBS 0.018472f
C583 B.n543 VSUBS 0.019358f
C584 B.n544 VSUBS 0.018515f
C585 B.n545 VSUBS 0.007852f
C586 B.n546 VSUBS 0.007852f
C587 B.n547 VSUBS 0.007852f
C588 B.n548 VSUBS 0.007852f
C589 B.n549 VSUBS 0.007852f
C590 B.n550 VSUBS 0.007852f
C591 B.n551 VSUBS 0.007852f
C592 B.n552 VSUBS 0.007852f
C593 B.n553 VSUBS 0.007852f
C594 B.n554 VSUBS 0.007852f
C595 B.n555 VSUBS 0.007852f
C596 B.n556 VSUBS 0.007852f
C597 B.n557 VSUBS 0.007852f
C598 B.n558 VSUBS 0.007852f
C599 B.n559 VSUBS 0.007852f
C600 B.n560 VSUBS 0.007852f
C601 B.n561 VSUBS 0.007852f
C602 B.n562 VSUBS 0.007852f
C603 B.n563 VSUBS 0.007852f
C604 B.n564 VSUBS 0.007852f
C605 B.n565 VSUBS 0.007852f
C606 B.n566 VSUBS 0.007852f
C607 B.n567 VSUBS 0.007852f
C608 B.n568 VSUBS 0.007852f
C609 B.n569 VSUBS 0.007852f
C610 B.n570 VSUBS 0.007852f
C611 B.n571 VSUBS 0.007852f
C612 B.n572 VSUBS 0.007852f
C613 B.n573 VSUBS 0.007852f
C614 B.n574 VSUBS 0.007852f
C615 B.n575 VSUBS 0.007852f
C616 B.n576 VSUBS 0.007852f
C617 B.n577 VSUBS 0.007852f
C618 B.n578 VSUBS 0.007852f
C619 B.n579 VSUBS 0.007852f
C620 B.n580 VSUBS 0.007852f
C621 B.n581 VSUBS 0.007852f
C622 B.n582 VSUBS 0.007852f
C623 B.n583 VSUBS 0.007852f
C624 B.n584 VSUBS 0.007852f
C625 B.n585 VSUBS 0.007852f
C626 B.n586 VSUBS 0.007852f
C627 B.n587 VSUBS 0.007852f
C628 B.n588 VSUBS 0.007852f
C629 B.n589 VSUBS 0.007852f
C630 B.n590 VSUBS 0.007852f
C631 B.n591 VSUBS 0.007852f
C632 B.n592 VSUBS 0.007852f
C633 B.n593 VSUBS 0.007852f
C634 B.n594 VSUBS 0.007852f
C635 B.n595 VSUBS 0.007852f
C636 B.n596 VSUBS 0.007852f
C637 B.n597 VSUBS 0.007852f
C638 B.n598 VSUBS 0.007852f
C639 B.n599 VSUBS 0.007852f
C640 B.n600 VSUBS 0.007852f
C641 B.n601 VSUBS 0.007852f
C642 B.n602 VSUBS 0.007852f
C643 B.n603 VSUBS 0.007852f
C644 B.n604 VSUBS 0.007852f
C645 B.n605 VSUBS 0.007852f
C646 B.n606 VSUBS 0.007852f
C647 B.n607 VSUBS 0.007852f
C648 B.n608 VSUBS 0.007852f
C649 B.n609 VSUBS 0.00739f
C650 B.n610 VSUBS 0.018192f
C651 B.n611 VSUBS 0.004388f
C652 B.n612 VSUBS 0.007852f
C653 B.n613 VSUBS 0.007852f
C654 B.n614 VSUBS 0.007852f
C655 B.n615 VSUBS 0.007852f
C656 B.n616 VSUBS 0.007852f
C657 B.n617 VSUBS 0.007852f
C658 B.n618 VSUBS 0.007852f
C659 B.n619 VSUBS 0.007852f
C660 B.n620 VSUBS 0.007852f
C661 B.n621 VSUBS 0.007852f
C662 B.n622 VSUBS 0.007852f
C663 B.n623 VSUBS 0.007852f
C664 B.n624 VSUBS 0.004388f
C665 B.n625 VSUBS 0.007852f
C666 B.n626 VSUBS 0.007852f
C667 B.n627 VSUBS 0.00739f
C668 B.n628 VSUBS 0.007852f
C669 B.n629 VSUBS 0.007852f
C670 B.n630 VSUBS 0.007852f
C671 B.n631 VSUBS 0.007852f
C672 B.n632 VSUBS 0.007852f
C673 B.n633 VSUBS 0.007852f
C674 B.n634 VSUBS 0.007852f
C675 B.n635 VSUBS 0.007852f
C676 B.n636 VSUBS 0.007852f
C677 B.n637 VSUBS 0.007852f
C678 B.n638 VSUBS 0.007852f
C679 B.n639 VSUBS 0.007852f
C680 B.n640 VSUBS 0.007852f
C681 B.n641 VSUBS 0.007852f
C682 B.n642 VSUBS 0.007852f
C683 B.n643 VSUBS 0.007852f
C684 B.n644 VSUBS 0.007852f
C685 B.n645 VSUBS 0.007852f
C686 B.n646 VSUBS 0.007852f
C687 B.n647 VSUBS 0.007852f
C688 B.n648 VSUBS 0.007852f
C689 B.n649 VSUBS 0.007852f
C690 B.n650 VSUBS 0.007852f
C691 B.n651 VSUBS 0.007852f
C692 B.n652 VSUBS 0.007852f
C693 B.n653 VSUBS 0.007852f
C694 B.n654 VSUBS 0.007852f
C695 B.n655 VSUBS 0.007852f
C696 B.n656 VSUBS 0.007852f
C697 B.n657 VSUBS 0.007852f
C698 B.n658 VSUBS 0.007852f
C699 B.n659 VSUBS 0.007852f
C700 B.n660 VSUBS 0.007852f
C701 B.n661 VSUBS 0.007852f
C702 B.n662 VSUBS 0.007852f
C703 B.n663 VSUBS 0.007852f
C704 B.n664 VSUBS 0.007852f
C705 B.n665 VSUBS 0.007852f
C706 B.n666 VSUBS 0.007852f
C707 B.n667 VSUBS 0.007852f
C708 B.n668 VSUBS 0.007852f
C709 B.n669 VSUBS 0.007852f
C710 B.n670 VSUBS 0.007852f
C711 B.n671 VSUBS 0.007852f
C712 B.n672 VSUBS 0.007852f
C713 B.n673 VSUBS 0.007852f
C714 B.n674 VSUBS 0.007852f
C715 B.n675 VSUBS 0.007852f
C716 B.n676 VSUBS 0.007852f
C717 B.n677 VSUBS 0.007852f
C718 B.n678 VSUBS 0.007852f
C719 B.n679 VSUBS 0.007852f
C720 B.n680 VSUBS 0.007852f
C721 B.n681 VSUBS 0.007852f
C722 B.n682 VSUBS 0.007852f
C723 B.n683 VSUBS 0.007852f
C724 B.n684 VSUBS 0.007852f
C725 B.n685 VSUBS 0.007852f
C726 B.n686 VSUBS 0.007852f
C727 B.n687 VSUBS 0.007852f
C728 B.n688 VSUBS 0.007852f
C729 B.n689 VSUBS 0.007852f
C730 B.n690 VSUBS 0.007852f
C731 B.n691 VSUBS 0.019402f
C732 B.n692 VSUBS 0.018472f
C733 B.n693 VSUBS 0.018472f
C734 B.n694 VSUBS 0.007852f
C735 B.n695 VSUBS 0.007852f
C736 B.n696 VSUBS 0.007852f
C737 B.n697 VSUBS 0.007852f
C738 B.n698 VSUBS 0.007852f
C739 B.n699 VSUBS 0.007852f
C740 B.n700 VSUBS 0.007852f
C741 B.n701 VSUBS 0.007852f
C742 B.n702 VSUBS 0.007852f
C743 B.n703 VSUBS 0.007852f
C744 B.n704 VSUBS 0.007852f
C745 B.n705 VSUBS 0.007852f
C746 B.n706 VSUBS 0.007852f
C747 B.n707 VSUBS 0.007852f
C748 B.n708 VSUBS 0.007852f
C749 B.n709 VSUBS 0.007852f
C750 B.n710 VSUBS 0.007852f
C751 B.n711 VSUBS 0.007852f
C752 B.n712 VSUBS 0.007852f
C753 B.n713 VSUBS 0.007852f
C754 B.n714 VSUBS 0.007852f
C755 B.n715 VSUBS 0.007852f
C756 B.n716 VSUBS 0.007852f
C757 B.n717 VSUBS 0.007852f
C758 B.n718 VSUBS 0.007852f
C759 B.n719 VSUBS 0.007852f
C760 B.n720 VSUBS 0.007852f
C761 B.n721 VSUBS 0.007852f
C762 B.n722 VSUBS 0.007852f
C763 B.n723 VSUBS 0.007852f
C764 B.n724 VSUBS 0.007852f
C765 B.n725 VSUBS 0.007852f
C766 B.n726 VSUBS 0.007852f
C767 B.n727 VSUBS 0.007852f
C768 B.n728 VSUBS 0.007852f
C769 B.n729 VSUBS 0.007852f
C770 B.n730 VSUBS 0.007852f
C771 B.n731 VSUBS 0.007852f
C772 B.n732 VSUBS 0.007852f
C773 B.n733 VSUBS 0.007852f
C774 B.n734 VSUBS 0.007852f
C775 B.n735 VSUBS 0.007852f
C776 B.n736 VSUBS 0.007852f
C777 B.n737 VSUBS 0.007852f
C778 B.n738 VSUBS 0.007852f
C779 B.n739 VSUBS 0.007852f
C780 B.n740 VSUBS 0.007852f
C781 B.n741 VSUBS 0.007852f
C782 B.n742 VSUBS 0.007852f
C783 B.n743 VSUBS 0.007852f
C784 B.n744 VSUBS 0.007852f
C785 B.n745 VSUBS 0.007852f
C786 B.n746 VSUBS 0.007852f
C787 B.n747 VSUBS 0.007852f
C788 B.n748 VSUBS 0.007852f
C789 B.n749 VSUBS 0.007852f
C790 B.n750 VSUBS 0.007852f
C791 B.n751 VSUBS 0.007852f
C792 B.n752 VSUBS 0.007852f
C793 B.n753 VSUBS 0.007852f
C794 B.n754 VSUBS 0.007852f
C795 B.n755 VSUBS 0.007852f
C796 B.n756 VSUBS 0.007852f
C797 B.n757 VSUBS 0.007852f
C798 B.n758 VSUBS 0.007852f
C799 B.n759 VSUBS 0.017779f
C800 VDD1.n0 VSUBS 0.031834f
C801 VDD1.n1 VSUBS 0.027999f
C802 VDD1.n2 VSUBS 0.015045f
C803 VDD1.n3 VSUBS 0.035562f
C804 VDD1.n4 VSUBS 0.01593f
C805 VDD1.n5 VSUBS 0.027999f
C806 VDD1.n6 VSUBS 0.015045f
C807 VDD1.n7 VSUBS 0.035562f
C808 VDD1.n8 VSUBS 0.01593f
C809 VDD1.n9 VSUBS 0.027999f
C810 VDD1.n10 VSUBS 0.015045f
C811 VDD1.n11 VSUBS 0.035562f
C812 VDD1.n12 VSUBS 0.01593f
C813 VDD1.n13 VSUBS 0.027999f
C814 VDD1.n14 VSUBS 0.015045f
C815 VDD1.n15 VSUBS 0.035562f
C816 VDD1.n16 VSUBS 0.035562f
C817 VDD1.n17 VSUBS 0.01593f
C818 VDD1.n18 VSUBS 0.027999f
C819 VDD1.n19 VSUBS 0.015045f
C820 VDD1.n20 VSUBS 0.035562f
C821 VDD1.n21 VSUBS 0.01593f
C822 VDD1.n22 VSUBS 0.231898f
C823 VDD1.t0 VSUBS 0.076715f
C824 VDD1.n23 VSUBS 0.026671f
C825 VDD1.n24 VSUBS 0.026751f
C826 VDD1.n25 VSUBS 0.015045f
C827 VDD1.n26 VSUBS 1.48608f
C828 VDD1.n27 VSUBS 0.027999f
C829 VDD1.n28 VSUBS 0.015045f
C830 VDD1.n29 VSUBS 0.01593f
C831 VDD1.n30 VSUBS 0.035562f
C832 VDD1.n31 VSUBS 0.035562f
C833 VDD1.n32 VSUBS 0.01593f
C834 VDD1.n33 VSUBS 0.015045f
C835 VDD1.n34 VSUBS 0.027999f
C836 VDD1.n35 VSUBS 0.027999f
C837 VDD1.n36 VSUBS 0.015045f
C838 VDD1.n37 VSUBS 0.01593f
C839 VDD1.n38 VSUBS 0.035562f
C840 VDD1.n39 VSUBS 0.035562f
C841 VDD1.n40 VSUBS 0.01593f
C842 VDD1.n41 VSUBS 0.015045f
C843 VDD1.n42 VSUBS 0.027999f
C844 VDD1.n43 VSUBS 0.027999f
C845 VDD1.n44 VSUBS 0.015045f
C846 VDD1.n45 VSUBS 0.015488f
C847 VDD1.n46 VSUBS 0.015488f
C848 VDD1.n47 VSUBS 0.035562f
C849 VDD1.n48 VSUBS 0.035562f
C850 VDD1.n49 VSUBS 0.01593f
C851 VDD1.n50 VSUBS 0.015045f
C852 VDD1.n51 VSUBS 0.027999f
C853 VDD1.n52 VSUBS 0.027999f
C854 VDD1.n53 VSUBS 0.015045f
C855 VDD1.n54 VSUBS 0.01593f
C856 VDD1.n55 VSUBS 0.035562f
C857 VDD1.n56 VSUBS 0.035562f
C858 VDD1.n57 VSUBS 0.01593f
C859 VDD1.n58 VSUBS 0.015045f
C860 VDD1.n59 VSUBS 0.027999f
C861 VDD1.n60 VSUBS 0.027999f
C862 VDD1.n61 VSUBS 0.015045f
C863 VDD1.n62 VSUBS 0.01593f
C864 VDD1.n63 VSUBS 0.035562f
C865 VDD1.n64 VSUBS 0.089734f
C866 VDD1.n65 VSUBS 0.01593f
C867 VDD1.n66 VSUBS 0.015045f
C868 VDD1.n67 VSUBS 0.067012f
C869 VDD1.n68 VSUBS 0.074021f
C870 VDD1.n69 VSUBS 0.031834f
C871 VDD1.n70 VSUBS 0.027999f
C872 VDD1.n71 VSUBS 0.015045f
C873 VDD1.n72 VSUBS 0.035562f
C874 VDD1.n73 VSUBS 0.01593f
C875 VDD1.n74 VSUBS 0.027999f
C876 VDD1.n75 VSUBS 0.015045f
C877 VDD1.n76 VSUBS 0.035562f
C878 VDD1.n77 VSUBS 0.01593f
C879 VDD1.n78 VSUBS 0.027999f
C880 VDD1.n79 VSUBS 0.015045f
C881 VDD1.n80 VSUBS 0.035562f
C882 VDD1.n81 VSUBS 0.01593f
C883 VDD1.n82 VSUBS 0.027999f
C884 VDD1.n83 VSUBS 0.015045f
C885 VDD1.n84 VSUBS 0.035562f
C886 VDD1.n85 VSUBS 0.01593f
C887 VDD1.n86 VSUBS 0.027999f
C888 VDD1.n87 VSUBS 0.015045f
C889 VDD1.n88 VSUBS 0.035562f
C890 VDD1.n89 VSUBS 0.01593f
C891 VDD1.n90 VSUBS 0.231898f
C892 VDD1.t1 VSUBS 0.076715f
C893 VDD1.n91 VSUBS 0.026671f
C894 VDD1.n92 VSUBS 0.026751f
C895 VDD1.n93 VSUBS 0.015045f
C896 VDD1.n94 VSUBS 1.48607f
C897 VDD1.n95 VSUBS 0.027999f
C898 VDD1.n96 VSUBS 0.015045f
C899 VDD1.n97 VSUBS 0.01593f
C900 VDD1.n98 VSUBS 0.035562f
C901 VDD1.n99 VSUBS 0.035562f
C902 VDD1.n100 VSUBS 0.01593f
C903 VDD1.n101 VSUBS 0.015045f
C904 VDD1.n102 VSUBS 0.027999f
C905 VDD1.n103 VSUBS 0.027999f
C906 VDD1.n104 VSUBS 0.015045f
C907 VDD1.n105 VSUBS 0.01593f
C908 VDD1.n106 VSUBS 0.035562f
C909 VDD1.n107 VSUBS 0.035562f
C910 VDD1.n108 VSUBS 0.035562f
C911 VDD1.n109 VSUBS 0.01593f
C912 VDD1.n110 VSUBS 0.015045f
C913 VDD1.n111 VSUBS 0.027999f
C914 VDD1.n112 VSUBS 0.027999f
C915 VDD1.n113 VSUBS 0.015045f
C916 VDD1.n114 VSUBS 0.015488f
C917 VDD1.n115 VSUBS 0.015488f
C918 VDD1.n116 VSUBS 0.035562f
C919 VDD1.n117 VSUBS 0.035562f
C920 VDD1.n118 VSUBS 0.01593f
C921 VDD1.n119 VSUBS 0.015045f
C922 VDD1.n120 VSUBS 0.027999f
C923 VDD1.n121 VSUBS 0.027999f
C924 VDD1.n122 VSUBS 0.015045f
C925 VDD1.n123 VSUBS 0.01593f
C926 VDD1.n124 VSUBS 0.035562f
C927 VDD1.n125 VSUBS 0.035562f
C928 VDD1.n126 VSUBS 0.01593f
C929 VDD1.n127 VSUBS 0.015045f
C930 VDD1.n128 VSUBS 0.027999f
C931 VDD1.n129 VSUBS 0.027999f
C932 VDD1.n130 VSUBS 0.015045f
C933 VDD1.n131 VSUBS 0.01593f
C934 VDD1.n132 VSUBS 0.035562f
C935 VDD1.n133 VSUBS 0.089734f
C936 VDD1.n134 VSUBS 0.01593f
C937 VDD1.n135 VSUBS 0.015045f
C938 VDD1.n136 VSUBS 0.067012f
C939 VDD1.n137 VSUBS 0.073152f
C940 VDD1.t4 VSUBS 0.285417f
C941 VDD1.t2 VSUBS 0.285417f
C942 VDD1.n138 VSUBS 2.26493f
C943 VDD1.n139 VSUBS 3.56624f
C944 VDD1.t5 VSUBS 0.285417f
C945 VDD1.t3 VSUBS 0.285417f
C946 VDD1.n140 VSUBS 2.25819f
C947 VDD1.n141 VSUBS 3.54055f
C948 VP.n0 VSUBS 0.03937f
C949 VP.t3 VSUBS 2.87093f
C950 VP.n1 VSUBS 0.058594f
C951 VP.n2 VSUBS 0.029861f
C952 VP.t1 VSUBS 2.87093f
C953 VP.n3 VSUBS 1.03829f
C954 VP.n4 VSUBS 0.029861f
C955 VP.n5 VSUBS 0.058594f
C956 VP.n6 VSUBS 0.03937f
C957 VP.t4 VSUBS 2.87093f
C958 VP.n7 VSUBS 0.03937f
C959 VP.t2 VSUBS 2.87093f
C960 VP.n8 VSUBS 0.058594f
C961 VP.n9 VSUBS 0.029861f
C962 VP.t0 VSUBS 2.87093f
C963 VP.n10 VSUBS 1.11645f
C964 VP.t5 VSUBS 3.14358f
C965 VP.n11 VSUBS 1.06776f
C966 VP.n12 VSUBS 0.311319f
C967 VP.n13 VSUBS 0.055932f
C968 VP.n14 VSUBS 0.060386f
C969 VP.n15 VSUBS 0.024513f
C970 VP.n16 VSUBS 0.029861f
C971 VP.n17 VSUBS 0.029861f
C972 VP.n18 VSUBS 0.029861f
C973 VP.n19 VSUBS 0.055932f
C974 VP.n20 VSUBS 0.03163f
C975 VP.n21 VSUBS 1.10451f
C976 VP.n22 VSUBS 1.65799f
C977 VP.n23 VSUBS 1.67948f
C978 VP.n24 VSUBS 1.10451f
C979 VP.n25 VSUBS 0.03163f
C980 VP.n26 VSUBS 0.055932f
C981 VP.n27 VSUBS 0.029861f
C982 VP.n28 VSUBS 0.029861f
C983 VP.n29 VSUBS 0.029861f
C984 VP.n30 VSUBS 0.024513f
C985 VP.n31 VSUBS 0.060386f
C986 VP.n32 VSUBS 0.055932f
C987 VP.n33 VSUBS 0.029861f
C988 VP.n34 VSUBS 0.029861f
C989 VP.n35 VSUBS 0.029861f
C990 VP.n36 VSUBS 0.055932f
C991 VP.n37 VSUBS 0.060386f
C992 VP.n38 VSUBS 0.024513f
C993 VP.n39 VSUBS 0.029861f
C994 VP.n40 VSUBS 0.029861f
C995 VP.n41 VSUBS 0.029861f
C996 VP.n42 VSUBS 0.055932f
C997 VP.n43 VSUBS 0.03163f
C998 VP.n44 VSUBS 1.10451f
C999 VP.n45 VSUBS 0.054866f
C1000 VDD2.n0 VSUBS 0.03184f
C1001 VDD2.n1 VSUBS 0.028003f
C1002 VDD2.n2 VSUBS 0.015048f
C1003 VDD2.n3 VSUBS 0.035568f
C1004 VDD2.n4 VSUBS 0.015933f
C1005 VDD2.n5 VSUBS 0.028003f
C1006 VDD2.n6 VSUBS 0.015048f
C1007 VDD2.n7 VSUBS 0.035568f
C1008 VDD2.n8 VSUBS 0.015933f
C1009 VDD2.n9 VSUBS 0.028003f
C1010 VDD2.n10 VSUBS 0.015048f
C1011 VDD2.n11 VSUBS 0.035568f
C1012 VDD2.n12 VSUBS 0.015933f
C1013 VDD2.n13 VSUBS 0.028003f
C1014 VDD2.n14 VSUBS 0.015048f
C1015 VDD2.n15 VSUBS 0.035568f
C1016 VDD2.n16 VSUBS 0.015933f
C1017 VDD2.n17 VSUBS 0.028003f
C1018 VDD2.n18 VSUBS 0.015048f
C1019 VDD2.n19 VSUBS 0.035568f
C1020 VDD2.n20 VSUBS 0.015933f
C1021 VDD2.n21 VSUBS 0.231938f
C1022 VDD2.t0 VSUBS 0.076728f
C1023 VDD2.n22 VSUBS 0.026676f
C1024 VDD2.n23 VSUBS 0.026756f
C1025 VDD2.n24 VSUBS 0.015048f
C1026 VDD2.n25 VSUBS 1.48633f
C1027 VDD2.n26 VSUBS 0.028003f
C1028 VDD2.n27 VSUBS 0.015048f
C1029 VDD2.n28 VSUBS 0.015933f
C1030 VDD2.n29 VSUBS 0.035568f
C1031 VDD2.n30 VSUBS 0.035568f
C1032 VDD2.n31 VSUBS 0.015933f
C1033 VDD2.n32 VSUBS 0.015048f
C1034 VDD2.n33 VSUBS 0.028003f
C1035 VDD2.n34 VSUBS 0.028003f
C1036 VDD2.n35 VSUBS 0.015048f
C1037 VDD2.n36 VSUBS 0.015933f
C1038 VDD2.n37 VSUBS 0.035568f
C1039 VDD2.n38 VSUBS 0.035568f
C1040 VDD2.n39 VSUBS 0.035568f
C1041 VDD2.n40 VSUBS 0.015933f
C1042 VDD2.n41 VSUBS 0.015048f
C1043 VDD2.n42 VSUBS 0.028003f
C1044 VDD2.n43 VSUBS 0.028003f
C1045 VDD2.n44 VSUBS 0.015048f
C1046 VDD2.n45 VSUBS 0.01549f
C1047 VDD2.n46 VSUBS 0.01549f
C1048 VDD2.n47 VSUBS 0.035568f
C1049 VDD2.n48 VSUBS 0.035568f
C1050 VDD2.n49 VSUBS 0.015933f
C1051 VDD2.n50 VSUBS 0.015048f
C1052 VDD2.n51 VSUBS 0.028003f
C1053 VDD2.n52 VSUBS 0.028003f
C1054 VDD2.n53 VSUBS 0.015048f
C1055 VDD2.n54 VSUBS 0.015933f
C1056 VDD2.n55 VSUBS 0.035568f
C1057 VDD2.n56 VSUBS 0.035568f
C1058 VDD2.n57 VSUBS 0.015933f
C1059 VDD2.n58 VSUBS 0.015048f
C1060 VDD2.n59 VSUBS 0.028003f
C1061 VDD2.n60 VSUBS 0.028003f
C1062 VDD2.n61 VSUBS 0.015048f
C1063 VDD2.n62 VSUBS 0.015933f
C1064 VDD2.n63 VSUBS 0.035568f
C1065 VDD2.n64 VSUBS 0.08975f
C1066 VDD2.n65 VSUBS 0.015933f
C1067 VDD2.n66 VSUBS 0.015048f
C1068 VDD2.n67 VSUBS 0.067024f
C1069 VDD2.n68 VSUBS 0.073164f
C1070 VDD2.t3 VSUBS 0.285465f
C1071 VDD2.t5 VSUBS 0.285465f
C1072 VDD2.n69 VSUBS 2.26531f
C1073 VDD2.n70 VSUBS 3.42323f
C1074 VDD2.n71 VSUBS 0.03184f
C1075 VDD2.n72 VSUBS 0.028003f
C1076 VDD2.n73 VSUBS 0.015048f
C1077 VDD2.n74 VSUBS 0.035568f
C1078 VDD2.n75 VSUBS 0.015933f
C1079 VDD2.n76 VSUBS 0.028003f
C1080 VDD2.n77 VSUBS 0.015048f
C1081 VDD2.n78 VSUBS 0.035568f
C1082 VDD2.n79 VSUBS 0.015933f
C1083 VDD2.n80 VSUBS 0.028003f
C1084 VDD2.n81 VSUBS 0.015048f
C1085 VDD2.n82 VSUBS 0.035568f
C1086 VDD2.n83 VSUBS 0.015933f
C1087 VDD2.n84 VSUBS 0.028003f
C1088 VDD2.n85 VSUBS 0.015048f
C1089 VDD2.n86 VSUBS 0.035568f
C1090 VDD2.n87 VSUBS 0.035568f
C1091 VDD2.n88 VSUBS 0.015933f
C1092 VDD2.n89 VSUBS 0.028003f
C1093 VDD2.n90 VSUBS 0.015048f
C1094 VDD2.n91 VSUBS 0.035568f
C1095 VDD2.n92 VSUBS 0.015933f
C1096 VDD2.n93 VSUBS 0.231938f
C1097 VDD2.t4 VSUBS 0.076728f
C1098 VDD2.n94 VSUBS 0.026676f
C1099 VDD2.n95 VSUBS 0.026756f
C1100 VDD2.n96 VSUBS 0.015048f
C1101 VDD2.n97 VSUBS 1.48633f
C1102 VDD2.n98 VSUBS 0.028003f
C1103 VDD2.n99 VSUBS 0.015048f
C1104 VDD2.n100 VSUBS 0.015933f
C1105 VDD2.n101 VSUBS 0.035568f
C1106 VDD2.n102 VSUBS 0.035568f
C1107 VDD2.n103 VSUBS 0.015933f
C1108 VDD2.n104 VSUBS 0.015048f
C1109 VDD2.n105 VSUBS 0.028003f
C1110 VDD2.n106 VSUBS 0.028003f
C1111 VDD2.n107 VSUBS 0.015048f
C1112 VDD2.n108 VSUBS 0.015933f
C1113 VDD2.n109 VSUBS 0.035568f
C1114 VDD2.n110 VSUBS 0.035568f
C1115 VDD2.n111 VSUBS 0.015933f
C1116 VDD2.n112 VSUBS 0.015048f
C1117 VDD2.n113 VSUBS 0.028003f
C1118 VDD2.n114 VSUBS 0.028003f
C1119 VDD2.n115 VSUBS 0.015048f
C1120 VDD2.n116 VSUBS 0.01549f
C1121 VDD2.n117 VSUBS 0.01549f
C1122 VDD2.n118 VSUBS 0.035568f
C1123 VDD2.n119 VSUBS 0.035568f
C1124 VDD2.n120 VSUBS 0.015933f
C1125 VDD2.n121 VSUBS 0.015048f
C1126 VDD2.n122 VSUBS 0.028003f
C1127 VDD2.n123 VSUBS 0.028003f
C1128 VDD2.n124 VSUBS 0.015048f
C1129 VDD2.n125 VSUBS 0.015933f
C1130 VDD2.n126 VSUBS 0.035568f
C1131 VDD2.n127 VSUBS 0.035568f
C1132 VDD2.n128 VSUBS 0.015933f
C1133 VDD2.n129 VSUBS 0.015048f
C1134 VDD2.n130 VSUBS 0.028003f
C1135 VDD2.n131 VSUBS 0.028003f
C1136 VDD2.n132 VSUBS 0.015048f
C1137 VDD2.n133 VSUBS 0.015933f
C1138 VDD2.n134 VSUBS 0.035568f
C1139 VDD2.n135 VSUBS 0.08975f
C1140 VDD2.n136 VSUBS 0.015933f
C1141 VDD2.n137 VSUBS 0.015048f
C1142 VDD2.n138 VSUBS 0.067024f
C1143 VDD2.n139 VSUBS 0.064684f
C1144 VDD2.n140 VSUBS 2.98786f
C1145 VDD2.t1 VSUBS 0.285465f
C1146 VDD2.t2 VSUBS 0.285465f
C1147 VDD2.n141 VSUBS 2.26527f
C1148 VTAIL.t8 VSUBS 0.294694f
C1149 VTAIL.t7 VSUBS 0.294694f
C1150 VTAIL.n0 VSUBS 2.17479f
C1151 VTAIL.n1 VSUBS 0.897011f
C1152 VTAIL.n2 VSUBS 0.032869f
C1153 VTAIL.n3 VSUBS 0.028909f
C1154 VTAIL.n4 VSUBS 0.015534f
C1155 VTAIL.n5 VSUBS 0.036717f
C1156 VTAIL.n6 VSUBS 0.016448f
C1157 VTAIL.n7 VSUBS 0.028909f
C1158 VTAIL.n8 VSUBS 0.015534f
C1159 VTAIL.n9 VSUBS 0.036717f
C1160 VTAIL.n10 VSUBS 0.016448f
C1161 VTAIL.n11 VSUBS 0.028909f
C1162 VTAIL.n12 VSUBS 0.015534f
C1163 VTAIL.n13 VSUBS 0.036717f
C1164 VTAIL.n14 VSUBS 0.016448f
C1165 VTAIL.n15 VSUBS 0.028909f
C1166 VTAIL.n16 VSUBS 0.015534f
C1167 VTAIL.n17 VSUBS 0.036717f
C1168 VTAIL.n18 VSUBS 0.016448f
C1169 VTAIL.n19 VSUBS 0.028909f
C1170 VTAIL.n20 VSUBS 0.015534f
C1171 VTAIL.n21 VSUBS 0.036717f
C1172 VTAIL.n22 VSUBS 0.016448f
C1173 VTAIL.n23 VSUBS 0.239436f
C1174 VTAIL.t4 VSUBS 0.079209f
C1175 VTAIL.n24 VSUBS 0.027538f
C1176 VTAIL.n25 VSUBS 0.027621f
C1177 VTAIL.n26 VSUBS 0.015534f
C1178 VTAIL.n27 VSUBS 1.53438f
C1179 VTAIL.n28 VSUBS 0.028909f
C1180 VTAIL.n29 VSUBS 0.015534f
C1181 VTAIL.n30 VSUBS 0.016448f
C1182 VTAIL.n31 VSUBS 0.036717f
C1183 VTAIL.n32 VSUBS 0.036717f
C1184 VTAIL.n33 VSUBS 0.016448f
C1185 VTAIL.n34 VSUBS 0.015534f
C1186 VTAIL.n35 VSUBS 0.028909f
C1187 VTAIL.n36 VSUBS 0.028909f
C1188 VTAIL.n37 VSUBS 0.015534f
C1189 VTAIL.n38 VSUBS 0.016448f
C1190 VTAIL.n39 VSUBS 0.036717f
C1191 VTAIL.n40 VSUBS 0.036717f
C1192 VTAIL.n41 VSUBS 0.036717f
C1193 VTAIL.n42 VSUBS 0.016448f
C1194 VTAIL.n43 VSUBS 0.015534f
C1195 VTAIL.n44 VSUBS 0.028909f
C1196 VTAIL.n45 VSUBS 0.028909f
C1197 VTAIL.n46 VSUBS 0.015534f
C1198 VTAIL.n47 VSUBS 0.015991f
C1199 VTAIL.n48 VSUBS 0.015991f
C1200 VTAIL.n49 VSUBS 0.036717f
C1201 VTAIL.n50 VSUBS 0.036717f
C1202 VTAIL.n51 VSUBS 0.016448f
C1203 VTAIL.n52 VSUBS 0.015534f
C1204 VTAIL.n53 VSUBS 0.028909f
C1205 VTAIL.n54 VSUBS 0.028909f
C1206 VTAIL.n55 VSUBS 0.015534f
C1207 VTAIL.n56 VSUBS 0.016448f
C1208 VTAIL.n57 VSUBS 0.036717f
C1209 VTAIL.n58 VSUBS 0.036717f
C1210 VTAIL.n59 VSUBS 0.016448f
C1211 VTAIL.n60 VSUBS 0.015534f
C1212 VTAIL.n61 VSUBS 0.028909f
C1213 VTAIL.n62 VSUBS 0.028909f
C1214 VTAIL.n63 VSUBS 0.015534f
C1215 VTAIL.n64 VSUBS 0.016448f
C1216 VTAIL.n65 VSUBS 0.036717f
C1217 VTAIL.n66 VSUBS 0.092651f
C1218 VTAIL.n67 VSUBS 0.016448f
C1219 VTAIL.n68 VSUBS 0.015534f
C1220 VTAIL.n69 VSUBS 0.069191f
C1221 VTAIL.n70 VSUBS 0.046832f
C1222 VTAIL.n71 VSUBS 0.438379f
C1223 VTAIL.t0 VSUBS 0.294694f
C1224 VTAIL.t2 VSUBS 0.294694f
C1225 VTAIL.n72 VSUBS 2.17479f
C1226 VTAIL.n73 VSUBS 2.82929f
C1227 VTAIL.t9 VSUBS 0.294694f
C1228 VTAIL.t6 VSUBS 0.294694f
C1229 VTAIL.n74 VSUBS 2.1748f
C1230 VTAIL.n75 VSUBS 2.82928f
C1231 VTAIL.n76 VSUBS 0.032869f
C1232 VTAIL.n77 VSUBS 0.028909f
C1233 VTAIL.n78 VSUBS 0.015534f
C1234 VTAIL.n79 VSUBS 0.036717f
C1235 VTAIL.n80 VSUBS 0.016448f
C1236 VTAIL.n81 VSUBS 0.028909f
C1237 VTAIL.n82 VSUBS 0.015534f
C1238 VTAIL.n83 VSUBS 0.036717f
C1239 VTAIL.n84 VSUBS 0.016448f
C1240 VTAIL.n85 VSUBS 0.028909f
C1241 VTAIL.n86 VSUBS 0.015534f
C1242 VTAIL.n87 VSUBS 0.036717f
C1243 VTAIL.n88 VSUBS 0.016448f
C1244 VTAIL.n89 VSUBS 0.028909f
C1245 VTAIL.n90 VSUBS 0.015534f
C1246 VTAIL.n91 VSUBS 0.036717f
C1247 VTAIL.n92 VSUBS 0.036717f
C1248 VTAIL.n93 VSUBS 0.016448f
C1249 VTAIL.n94 VSUBS 0.028909f
C1250 VTAIL.n95 VSUBS 0.015534f
C1251 VTAIL.n96 VSUBS 0.036717f
C1252 VTAIL.n97 VSUBS 0.016448f
C1253 VTAIL.n98 VSUBS 0.239436f
C1254 VTAIL.t10 VSUBS 0.079209f
C1255 VTAIL.n99 VSUBS 0.027538f
C1256 VTAIL.n100 VSUBS 0.027621f
C1257 VTAIL.n101 VSUBS 0.015534f
C1258 VTAIL.n102 VSUBS 1.53438f
C1259 VTAIL.n103 VSUBS 0.028909f
C1260 VTAIL.n104 VSUBS 0.015534f
C1261 VTAIL.n105 VSUBS 0.016448f
C1262 VTAIL.n106 VSUBS 0.036717f
C1263 VTAIL.n107 VSUBS 0.036717f
C1264 VTAIL.n108 VSUBS 0.016448f
C1265 VTAIL.n109 VSUBS 0.015534f
C1266 VTAIL.n110 VSUBS 0.028909f
C1267 VTAIL.n111 VSUBS 0.028909f
C1268 VTAIL.n112 VSUBS 0.015534f
C1269 VTAIL.n113 VSUBS 0.016448f
C1270 VTAIL.n114 VSUBS 0.036717f
C1271 VTAIL.n115 VSUBS 0.036717f
C1272 VTAIL.n116 VSUBS 0.016448f
C1273 VTAIL.n117 VSUBS 0.015534f
C1274 VTAIL.n118 VSUBS 0.028909f
C1275 VTAIL.n119 VSUBS 0.028909f
C1276 VTAIL.n120 VSUBS 0.015534f
C1277 VTAIL.n121 VSUBS 0.015991f
C1278 VTAIL.n122 VSUBS 0.015991f
C1279 VTAIL.n123 VSUBS 0.036717f
C1280 VTAIL.n124 VSUBS 0.036717f
C1281 VTAIL.n125 VSUBS 0.016448f
C1282 VTAIL.n126 VSUBS 0.015534f
C1283 VTAIL.n127 VSUBS 0.028909f
C1284 VTAIL.n128 VSUBS 0.028909f
C1285 VTAIL.n129 VSUBS 0.015534f
C1286 VTAIL.n130 VSUBS 0.016448f
C1287 VTAIL.n131 VSUBS 0.036717f
C1288 VTAIL.n132 VSUBS 0.036717f
C1289 VTAIL.n133 VSUBS 0.016448f
C1290 VTAIL.n134 VSUBS 0.015534f
C1291 VTAIL.n135 VSUBS 0.028909f
C1292 VTAIL.n136 VSUBS 0.028909f
C1293 VTAIL.n137 VSUBS 0.015534f
C1294 VTAIL.n138 VSUBS 0.016448f
C1295 VTAIL.n139 VSUBS 0.036717f
C1296 VTAIL.n140 VSUBS 0.092651f
C1297 VTAIL.n141 VSUBS 0.016448f
C1298 VTAIL.n142 VSUBS 0.015534f
C1299 VTAIL.n143 VSUBS 0.069191f
C1300 VTAIL.n144 VSUBS 0.046832f
C1301 VTAIL.n145 VSUBS 0.438379f
C1302 VTAIL.t3 VSUBS 0.294694f
C1303 VTAIL.t5 VSUBS 0.294694f
C1304 VTAIL.n146 VSUBS 2.1748f
C1305 VTAIL.n147 VSUBS 1.07587f
C1306 VTAIL.n148 VSUBS 0.032869f
C1307 VTAIL.n149 VSUBS 0.028909f
C1308 VTAIL.n150 VSUBS 0.015534f
C1309 VTAIL.n151 VSUBS 0.036717f
C1310 VTAIL.n152 VSUBS 0.016448f
C1311 VTAIL.n153 VSUBS 0.028909f
C1312 VTAIL.n154 VSUBS 0.015534f
C1313 VTAIL.n155 VSUBS 0.036717f
C1314 VTAIL.n156 VSUBS 0.016448f
C1315 VTAIL.n157 VSUBS 0.028909f
C1316 VTAIL.n158 VSUBS 0.015534f
C1317 VTAIL.n159 VSUBS 0.036717f
C1318 VTAIL.n160 VSUBS 0.016448f
C1319 VTAIL.n161 VSUBS 0.028909f
C1320 VTAIL.n162 VSUBS 0.015534f
C1321 VTAIL.n163 VSUBS 0.036717f
C1322 VTAIL.n164 VSUBS 0.036717f
C1323 VTAIL.n165 VSUBS 0.016448f
C1324 VTAIL.n166 VSUBS 0.028909f
C1325 VTAIL.n167 VSUBS 0.015534f
C1326 VTAIL.n168 VSUBS 0.036717f
C1327 VTAIL.n169 VSUBS 0.016448f
C1328 VTAIL.n170 VSUBS 0.239436f
C1329 VTAIL.t1 VSUBS 0.079209f
C1330 VTAIL.n171 VSUBS 0.027538f
C1331 VTAIL.n172 VSUBS 0.027621f
C1332 VTAIL.n173 VSUBS 0.015534f
C1333 VTAIL.n174 VSUBS 1.53438f
C1334 VTAIL.n175 VSUBS 0.028909f
C1335 VTAIL.n176 VSUBS 0.015534f
C1336 VTAIL.n177 VSUBS 0.016448f
C1337 VTAIL.n178 VSUBS 0.036717f
C1338 VTAIL.n179 VSUBS 0.036717f
C1339 VTAIL.n180 VSUBS 0.016448f
C1340 VTAIL.n181 VSUBS 0.015534f
C1341 VTAIL.n182 VSUBS 0.028909f
C1342 VTAIL.n183 VSUBS 0.028909f
C1343 VTAIL.n184 VSUBS 0.015534f
C1344 VTAIL.n185 VSUBS 0.016448f
C1345 VTAIL.n186 VSUBS 0.036717f
C1346 VTAIL.n187 VSUBS 0.036717f
C1347 VTAIL.n188 VSUBS 0.016448f
C1348 VTAIL.n189 VSUBS 0.015534f
C1349 VTAIL.n190 VSUBS 0.028909f
C1350 VTAIL.n191 VSUBS 0.028909f
C1351 VTAIL.n192 VSUBS 0.015534f
C1352 VTAIL.n193 VSUBS 0.015991f
C1353 VTAIL.n194 VSUBS 0.015991f
C1354 VTAIL.n195 VSUBS 0.036717f
C1355 VTAIL.n196 VSUBS 0.036717f
C1356 VTAIL.n197 VSUBS 0.016448f
C1357 VTAIL.n198 VSUBS 0.015534f
C1358 VTAIL.n199 VSUBS 0.028909f
C1359 VTAIL.n200 VSUBS 0.028909f
C1360 VTAIL.n201 VSUBS 0.015534f
C1361 VTAIL.n202 VSUBS 0.016448f
C1362 VTAIL.n203 VSUBS 0.036717f
C1363 VTAIL.n204 VSUBS 0.036717f
C1364 VTAIL.n205 VSUBS 0.016448f
C1365 VTAIL.n206 VSUBS 0.015534f
C1366 VTAIL.n207 VSUBS 0.028909f
C1367 VTAIL.n208 VSUBS 0.028909f
C1368 VTAIL.n209 VSUBS 0.015534f
C1369 VTAIL.n210 VSUBS 0.016448f
C1370 VTAIL.n211 VSUBS 0.036717f
C1371 VTAIL.n212 VSUBS 0.092651f
C1372 VTAIL.n213 VSUBS 0.016448f
C1373 VTAIL.n214 VSUBS 0.015534f
C1374 VTAIL.n215 VSUBS 0.069191f
C1375 VTAIL.n216 VSUBS 0.046832f
C1376 VTAIL.n217 VSUBS 1.94606f
C1377 VTAIL.n218 VSUBS 0.032869f
C1378 VTAIL.n219 VSUBS 0.028909f
C1379 VTAIL.n220 VSUBS 0.015534f
C1380 VTAIL.n221 VSUBS 0.036717f
C1381 VTAIL.n222 VSUBS 0.016448f
C1382 VTAIL.n223 VSUBS 0.028909f
C1383 VTAIL.n224 VSUBS 0.015534f
C1384 VTAIL.n225 VSUBS 0.036717f
C1385 VTAIL.n226 VSUBS 0.016448f
C1386 VTAIL.n227 VSUBS 0.028909f
C1387 VTAIL.n228 VSUBS 0.015534f
C1388 VTAIL.n229 VSUBS 0.036717f
C1389 VTAIL.n230 VSUBS 0.016448f
C1390 VTAIL.n231 VSUBS 0.028909f
C1391 VTAIL.n232 VSUBS 0.015534f
C1392 VTAIL.n233 VSUBS 0.036717f
C1393 VTAIL.n234 VSUBS 0.016448f
C1394 VTAIL.n235 VSUBS 0.028909f
C1395 VTAIL.n236 VSUBS 0.015534f
C1396 VTAIL.n237 VSUBS 0.036717f
C1397 VTAIL.n238 VSUBS 0.016448f
C1398 VTAIL.n239 VSUBS 0.239436f
C1399 VTAIL.t11 VSUBS 0.079209f
C1400 VTAIL.n240 VSUBS 0.027538f
C1401 VTAIL.n241 VSUBS 0.027621f
C1402 VTAIL.n242 VSUBS 0.015534f
C1403 VTAIL.n243 VSUBS 1.53438f
C1404 VTAIL.n244 VSUBS 0.028909f
C1405 VTAIL.n245 VSUBS 0.015534f
C1406 VTAIL.n246 VSUBS 0.016448f
C1407 VTAIL.n247 VSUBS 0.036717f
C1408 VTAIL.n248 VSUBS 0.036717f
C1409 VTAIL.n249 VSUBS 0.016448f
C1410 VTAIL.n250 VSUBS 0.015534f
C1411 VTAIL.n251 VSUBS 0.028909f
C1412 VTAIL.n252 VSUBS 0.028909f
C1413 VTAIL.n253 VSUBS 0.015534f
C1414 VTAIL.n254 VSUBS 0.016448f
C1415 VTAIL.n255 VSUBS 0.036717f
C1416 VTAIL.n256 VSUBS 0.036717f
C1417 VTAIL.n257 VSUBS 0.036717f
C1418 VTAIL.n258 VSUBS 0.016448f
C1419 VTAIL.n259 VSUBS 0.015534f
C1420 VTAIL.n260 VSUBS 0.028909f
C1421 VTAIL.n261 VSUBS 0.028909f
C1422 VTAIL.n262 VSUBS 0.015534f
C1423 VTAIL.n263 VSUBS 0.015991f
C1424 VTAIL.n264 VSUBS 0.015991f
C1425 VTAIL.n265 VSUBS 0.036717f
C1426 VTAIL.n266 VSUBS 0.036717f
C1427 VTAIL.n267 VSUBS 0.016448f
C1428 VTAIL.n268 VSUBS 0.015534f
C1429 VTAIL.n269 VSUBS 0.028909f
C1430 VTAIL.n270 VSUBS 0.028909f
C1431 VTAIL.n271 VSUBS 0.015534f
C1432 VTAIL.n272 VSUBS 0.016448f
C1433 VTAIL.n273 VSUBS 0.036717f
C1434 VTAIL.n274 VSUBS 0.036717f
C1435 VTAIL.n275 VSUBS 0.016448f
C1436 VTAIL.n276 VSUBS 0.015534f
C1437 VTAIL.n277 VSUBS 0.028909f
C1438 VTAIL.n278 VSUBS 0.028909f
C1439 VTAIL.n279 VSUBS 0.015534f
C1440 VTAIL.n280 VSUBS 0.016448f
C1441 VTAIL.n281 VSUBS 0.036717f
C1442 VTAIL.n282 VSUBS 0.092651f
C1443 VTAIL.n283 VSUBS 0.016448f
C1444 VTAIL.n284 VSUBS 0.015534f
C1445 VTAIL.n285 VSUBS 0.069191f
C1446 VTAIL.n286 VSUBS 0.046832f
C1447 VTAIL.n287 VSUBS 1.87921f
C1448 VN.n0 VSUBS 0.038237f
C1449 VN.t0 VSUBS 2.78826f
C1450 VN.n1 VSUBS 0.056907f
C1451 VN.n2 VSUBS 0.029001f
C1452 VN.t2 VSUBS 2.78826f
C1453 VN.n3 VSUBS 1.0843f
C1454 VN.t5 VSUBS 3.05306f
C1455 VN.n4 VSUBS 1.03702f
C1456 VN.n5 VSUBS 0.302355f
C1457 VN.n6 VSUBS 0.054321f
C1458 VN.n7 VSUBS 0.058647f
C1459 VN.n8 VSUBS 0.023807f
C1460 VN.n9 VSUBS 0.029001f
C1461 VN.n10 VSUBS 0.029001f
C1462 VN.n11 VSUBS 0.029001f
C1463 VN.n12 VSUBS 0.054321f
C1464 VN.n13 VSUBS 0.030719f
C1465 VN.n14 VSUBS 1.07271f
C1466 VN.n15 VSUBS 0.053286f
C1467 VN.n16 VSUBS 0.038237f
C1468 VN.t1 VSUBS 2.78826f
C1469 VN.n17 VSUBS 0.056907f
C1470 VN.n18 VSUBS 0.029001f
C1471 VN.t4 VSUBS 2.78826f
C1472 VN.n19 VSUBS 1.0843f
C1473 VN.t3 VSUBS 3.05306f
C1474 VN.n20 VSUBS 1.03702f
C1475 VN.n21 VSUBS 0.302355f
C1476 VN.n22 VSUBS 0.054321f
C1477 VN.n23 VSUBS 0.058647f
C1478 VN.n24 VSUBS 0.023807f
C1479 VN.n25 VSUBS 0.029001f
C1480 VN.n26 VSUBS 0.029001f
C1481 VN.n27 VSUBS 0.029001f
C1482 VN.n28 VSUBS 0.054321f
C1483 VN.n29 VSUBS 0.030719f
C1484 VN.n30 VSUBS 1.07271f
C1485 VN.n31 VSUBS 1.62584f
.ends

