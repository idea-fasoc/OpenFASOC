* NGSPICE file created from diff_pair_sample_0135.ext - technology: sky130A

.subckt diff_pair_sample_0135 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=2.55
X1 B.t8 B.t6 B.t7 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=2.55
X2 VTAIL.t7 VP.t0 VDD1.t2 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=2.55
X3 VTAIL.t0 VN.t0 VDD2.t3 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=2.55
X4 VDD2.t2 VN.t1 VTAIL.t1 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=2.55
X5 VTAIL.t2 VN.t2 VDD2.t1 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=2.55
X6 VDD1.t3 VP.t1 VTAIL.t6 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=2.55
X7 VTAIL.t5 VP.t2 VDD1.t0 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=2.74725 ps=16.98 w=16.65 l=2.55
X8 B.t5 B.t3 B.t4 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=2.55
X9 VDD2.t0 VN.t3 VTAIL.t3 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=2.55
X10 VDD1.t1 VP.t3 VTAIL.t4 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=2.74725 pd=16.98 as=6.4935 ps=34.08 w=16.65 l=2.55
X11 B.t2 B.t0 B.t1 w_n2698_n4298# sky130_fd_pr__pfet_01v8 ad=6.4935 pd=34.08 as=0 ps=0 w=16.65 l=2.55
R0 B.n426 B.n117 585
R1 B.n425 B.n424 585
R2 B.n423 B.n118 585
R3 B.n422 B.n421 585
R4 B.n420 B.n119 585
R5 B.n419 B.n418 585
R6 B.n417 B.n120 585
R7 B.n416 B.n415 585
R8 B.n414 B.n121 585
R9 B.n413 B.n412 585
R10 B.n411 B.n122 585
R11 B.n410 B.n409 585
R12 B.n408 B.n123 585
R13 B.n407 B.n406 585
R14 B.n405 B.n124 585
R15 B.n404 B.n403 585
R16 B.n402 B.n125 585
R17 B.n401 B.n400 585
R18 B.n399 B.n126 585
R19 B.n398 B.n397 585
R20 B.n396 B.n127 585
R21 B.n395 B.n394 585
R22 B.n393 B.n128 585
R23 B.n392 B.n391 585
R24 B.n390 B.n129 585
R25 B.n389 B.n388 585
R26 B.n387 B.n130 585
R27 B.n386 B.n385 585
R28 B.n384 B.n131 585
R29 B.n383 B.n382 585
R30 B.n381 B.n132 585
R31 B.n380 B.n379 585
R32 B.n378 B.n133 585
R33 B.n377 B.n376 585
R34 B.n375 B.n134 585
R35 B.n374 B.n373 585
R36 B.n372 B.n135 585
R37 B.n371 B.n370 585
R38 B.n369 B.n136 585
R39 B.n368 B.n367 585
R40 B.n366 B.n137 585
R41 B.n365 B.n364 585
R42 B.n363 B.n138 585
R43 B.n362 B.n361 585
R44 B.n360 B.n139 585
R45 B.n359 B.n358 585
R46 B.n357 B.n140 585
R47 B.n356 B.n355 585
R48 B.n354 B.n141 585
R49 B.n353 B.n352 585
R50 B.n351 B.n142 585
R51 B.n350 B.n349 585
R52 B.n348 B.n143 585
R53 B.n347 B.n346 585
R54 B.n345 B.n144 585
R55 B.n344 B.n343 585
R56 B.n339 B.n145 585
R57 B.n338 B.n337 585
R58 B.n336 B.n146 585
R59 B.n335 B.n334 585
R60 B.n333 B.n147 585
R61 B.n332 B.n331 585
R62 B.n330 B.n148 585
R63 B.n329 B.n328 585
R64 B.n327 B.n149 585
R65 B.n325 B.n324 585
R66 B.n323 B.n152 585
R67 B.n322 B.n321 585
R68 B.n320 B.n153 585
R69 B.n319 B.n318 585
R70 B.n317 B.n154 585
R71 B.n316 B.n315 585
R72 B.n314 B.n155 585
R73 B.n313 B.n312 585
R74 B.n311 B.n156 585
R75 B.n310 B.n309 585
R76 B.n308 B.n157 585
R77 B.n307 B.n306 585
R78 B.n305 B.n158 585
R79 B.n304 B.n303 585
R80 B.n302 B.n159 585
R81 B.n301 B.n300 585
R82 B.n299 B.n160 585
R83 B.n298 B.n297 585
R84 B.n296 B.n161 585
R85 B.n295 B.n294 585
R86 B.n293 B.n162 585
R87 B.n292 B.n291 585
R88 B.n290 B.n163 585
R89 B.n289 B.n288 585
R90 B.n287 B.n164 585
R91 B.n286 B.n285 585
R92 B.n284 B.n165 585
R93 B.n283 B.n282 585
R94 B.n281 B.n166 585
R95 B.n280 B.n279 585
R96 B.n278 B.n167 585
R97 B.n277 B.n276 585
R98 B.n275 B.n168 585
R99 B.n274 B.n273 585
R100 B.n272 B.n169 585
R101 B.n271 B.n270 585
R102 B.n269 B.n170 585
R103 B.n268 B.n267 585
R104 B.n266 B.n171 585
R105 B.n265 B.n264 585
R106 B.n263 B.n172 585
R107 B.n262 B.n261 585
R108 B.n260 B.n173 585
R109 B.n259 B.n258 585
R110 B.n257 B.n174 585
R111 B.n256 B.n255 585
R112 B.n254 B.n175 585
R113 B.n253 B.n252 585
R114 B.n251 B.n176 585
R115 B.n250 B.n249 585
R116 B.n248 B.n177 585
R117 B.n247 B.n246 585
R118 B.n245 B.n178 585
R119 B.n244 B.n243 585
R120 B.n428 B.n427 585
R121 B.n429 B.n116 585
R122 B.n431 B.n430 585
R123 B.n432 B.n115 585
R124 B.n434 B.n433 585
R125 B.n435 B.n114 585
R126 B.n437 B.n436 585
R127 B.n438 B.n113 585
R128 B.n440 B.n439 585
R129 B.n441 B.n112 585
R130 B.n443 B.n442 585
R131 B.n444 B.n111 585
R132 B.n446 B.n445 585
R133 B.n447 B.n110 585
R134 B.n449 B.n448 585
R135 B.n450 B.n109 585
R136 B.n452 B.n451 585
R137 B.n453 B.n108 585
R138 B.n455 B.n454 585
R139 B.n456 B.n107 585
R140 B.n458 B.n457 585
R141 B.n459 B.n106 585
R142 B.n461 B.n460 585
R143 B.n462 B.n105 585
R144 B.n464 B.n463 585
R145 B.n465 B.n104 585
R146 B.n467 B.n466 585
R147 B.n468 B.n103 585
R148 B.n470 B.n469 585
R149 B.n471 B.n102 585
R150 B.n473 B.n472 585
R151 B.n474 B.n101 585
R152 B.n476 B.n475 585
R153 B.n477 B.n100 585
R154 B.n479 B.n478 585
R155 B.n480 B.n99 585
R156 B.n482 B.n481 585
R157 B.n483 B.n98 585
R158 B.n485 B.n484 585
R159 B.n486 B.n97 585
R160 B.n488 B.n487 585
R161 B.n489 B.n96 585
R162 B.n491 B.n490 585
R163 B.n492 B.n95 585
R164 B.n494 B.n493 585
R165 B.n495 B.n94 585
R166 B.n497 B.n496 585
R167 B.n498 B.n93 585
R168 B.n500 B.n499 585
R169 B.n501 B.n92 585
R170 B.n503 B.n502 585
R171 B.n504 B.n91 585
R172 B.n506 B.n505 585
R173 B.n507 B.n90 585
R174 B.n509 B.n508 585
R175 B.n510 B.n89 585
R176 B.n512 B.n511 585
R177 B.n513 B.n88 585
R178 B.n515 B.n514 585
R179 B.n516 B.n87 585
R180 B.n518 B.n517 585
R181 B.n519 B.n86 585
R182 B.n521 B.n520 585
R183 B.n522 B.n85 585
R184 B.n524 B.n523 585
R185 B.n525 B.n84 585
R186 B.n527 B.n526 585
R187 B.n528 B.n83 585
R188 B.n710 B.n709 585
R189 B.n708 B.n19 585
R190 B.n707 B.n706 585
R191 B.n705 B.n20 585
R192 B.n704 B.n703 585
R193 B.n702 B.n21 585
R194 B.n701 B.n700 585
R195 B.n699 B.n22 585
R196 B.n698 B.n697 585
R197 B.n696 B.n23 585
R198 B.n695 B.n694 585
R199 B.n693 B.n24 585
R200 B.n692 B.n691 585
R201 B.n690 B.n25 585
R202 B.n689 B.n688 585
R203 B.n687 B.n26 585
R204 B.n686 B.n685 585
R205 B.n684 B.n27 585
R206 B.n683 B.n682 585
R207 B.n681 B.n28 585
R208 B.n680 B.n679 585
R209 B.n678 B.n29 585
R210 B.n677 B.n676 585
R211 B.n675 B.n30 585
R212 B.n674 B.n673 585
R213 B.n672 B.n31 585
R214 B.n671 B.n670 585
R215 B.n669 B.n32 585
R216 B.n668 B.n667 585
R217 B.n666 B.n33 585
R218 B.n665 B.n664 585
R219 B.n663 B.n34 585
R220 B.n662 B.n661 585
R221 B.n660 B.n35 585
R222 B.n659 B.n658 585
R223 B.n657 B.n36 585
R224 B.n656 B.n655 585
R225 B.n654 B.n37 585
R226 B.n653 B.n652 585
R227 B.n651 B.n38 585
R228 B.n650 B.n649 585
R229 B.n648 B.n39 585
R230 B.n647 B.n646 585
R231 B.n645 B.n40 585
R232 B.n644 B.n643 585
R233 B.n642 B.n41 585
R234 B.n641 B.n640 585
R235 B.n639 B.n42 585
R236 B.n638 B.n637 585
R237 B.n636 B.n43 585
R238 B.n635 B.n634 585
R239 B.n633 B.n44 585
R240 B.n632 B.n631 585
R241 B.n630 B.n45 585
R242 B.n629 B.n628 585
R243 B.n627 B.n626 585
R244 B.n625 B.n49 585
R245 B.n624 B.n623 585
R246 B.n622 B.n50 585
R247 B.n621 B.n620 585
R248 B.n619 B.n51 585
R249 B.n618 B.n617 585
R250 B.n616 B.n52 585
R251 B.n615 B.n614 585
R252 B.n613 B.n53 585
R253 B.n611 B.n610 585
R254 B.n609 B.n56 585
R255 B.n608 B.n607 585
R256 B.n606 B.n57 585
R257 B.n605 B.n604 585
R258 B.n603 B.n58 585
R259 B.n602 B.n601 585
R260 B.n600 B.n59 585
R261 B.n599 B.n598 585
R262 B.n597 B.n60 585
R263 B.n596 B.n595 585
R264 B.n594 B.n61 585
R265 B.n593 B.n592 585
R266 B.n591 B.n62 585
R267 B.n590 B.n589 585
R268 B.n588 B.n63 585
R269 B.n587 B.n586 585
R270 B.n585 B.n64 585
R271 B.n584 B.n583 585
R272 B.n582 B.n65 585
R273 B.n581 B.n580 585
R274 B.n579 B.n66 585
R275 B.n578 B.n577 585
R276 B.n576 B.n67 585
R277 B.n575 B.n574 585
R278 B.n573 B.n68 585
R279 B.n572 B.n571 585
R280 B.n570 B.n69 585
R281 B.n569 B.n568 585
R282 B.n567 B.n70 585
R283 B.n566 B.n565 585
R284 B.n564 B.n71 585
R285 B.n563 B.n562 585
R286 B.n561 B.n72 585
R287 B.n560 B.n559 585
R288 B.n558 B.n73 585
R289 B.n557 B.n556 585
R290 B.n555 B.n74 585
R291 B.n554 B.n553 585
R292 B.n552 B.n75 585
R293 B.n551 B.n550 585
R294 B.n549 B.n76 585
R295 B.n548 B.n547 585
R296 B.n546 B.n77 585
R297 B.n545 B.n544 585
R298 B.n543 B.n78 585
R299 B.n542 B.n541 585
R300 B.n540 B.n79 585
R301 B.n539 B.n538 585
R302 B.n537 B.n80 585
R303 B.n536 B.n535 585
R304 B.n534 B.n81 585
R305 B.n533 B.n532 585
R306 B.n531 B.n82 585
R307 B.n530 B.n529 585
R308 B.n711 B.n18 585
R309 B.n713 B.n712 585
R310 B.n714 B.n17 585
R311 B.n716 B.n715 585
R312 B.n717 B.n16 585
R313 B.n719 B.n718 585
R314 B.n720 B.n15 585
R315 B.n722 B.n721 585
R316 B.n723 B.n14 585
R317 B.n725 B.n724 585
R318 B.n726 B.n13 585
R319 B.n728 B.n727 585
R320 B.n729 B.n12 585
R321 B.n731 B.n730 585
R322 B.n732 B.n11 585
R323 B.n734 B.n733 585
R324 B.n735 B.n10 585
R325 B.n737 B.n736 585
R326 B.n738 B.n9 585
R327 B.n740 B.n739 585
R328 B.n741 B.n8 585
R329 B.n743 B.n742 585
R330 B.n744 B.n7 585
R331 B.n746 B.n745 585
R332 B.n747 B.n6 585
R333 B.n749 B.n748 585
R334 B.n750 B.n5 585
R335 B.n752 B.n751 585
R336 B.n753 B.n4 585
R337 B.n755 B.n754 585
R338 B.n756 B.n3 585
R339 B.n758 B.n757 585
R340 B.n759 B.n0 585
R341 B.n2 B.n1 585
R342 B.n196 B.n195 585
R343 B.n197 B.n194 585
R344 B.n199 B.n198 585
R345 B.n200 B.n193 585
R346 B.n202 B.n201 585
R347 B.n203 B.n192 585
R348 B.n205 B.n204 585
R349 B.n206 B.n191 585
R350 B.n208 B.n207 585
R351 B.n209 B.n190 585
R352 B.n211 B.n210 585
R353 B.n212 B.n189 585
R354 B.n214 B.n213 585
R355 B.n215 B.n188 585
R356 B.n217 B.n216 585
R357 B.n218 B.n187 585
R358 B.n220 B.n219 585
R359 B.n221 B.n186 585
R360 B.n223 B.n222 585
R361 B.n224 B.n185 585
R362 B.n226 B.n225 585
R363 B.n227 B.n184 585
R364 B.n229 B.n228 585
R365 B.n230 B.n183 585
R366 B.n232 B.n231 585
R367 B.n233 B.n182 585
R368 B.n235 B.n234 585
R369 B.n236 B.n181 585
R370 B.n238 B.n237 585
R371 B.n239 B.n180 585
R372 B.n241 B.n240 585
R373 B.n242 B.n179 585
R374 B.n244 B.n179 516.524
R375 B.n428 B.n117 516.524
R376 B.n530 B.n83 516.524
R377 B.n711 B.n710 516.524
R378 B.n150 B.t0 365.329
R379 B.n340 B.t3 365.329
R380 B.n54 B.t9 365.329
R381 B.n46 B.t6 365.329
R382 B.n761 B.n760 256.663
R383 B.n760 B.n759 235.042
R384 B.n760 B.n2 235.042
R385 B.n340 B.t4 168.602
R386 B.n54 B.t11 168.602
R387 B.n150 B.t1 168.582
R388 B.n46 B.t8 168.582
R389 B.n245 B.n244 163.367
R390 B.n246 B.n245 163.367
R391 B.n246 B.n177 163.367
R392 B.n250 B.n177 163.367
R393 B.n251 B.n250 163.367
R394 B.n252 B.n251 163.367
R395 B.n252 B.n175 163.367
R396 B.n256 B.n175 163.367
R397 B.n257 B.n256 163.367
R398 B.n258 B.n257 163.367
R399 B.n258 B.n173 163.367
R400 B.n262 B.n173 163.367
R401 B.n263 B.n262 163.367
R402 B.n264 B.n263 163.367
R403 B.n264 B.n171 163.367
R404 B.n268 B.n171 163.367
R405 B.n269 B.n268 163.367
R406 B.n270 B.n269 163.367
R407 B.n270 B.n169 163.367
R408 B.n274 B.n169 163.367
R409 B.n275 B.n274 163.367
R410 B.n276 B.n275 163.367
R411 B.n276 B.n167 163.367
R412 B.n280 B.n167 163.367
R413 B.n281 B.n280 163.367
R414 B.n282 B.n281 163.367
R415 B.n282 B.n165 163.367
R416 B.n286 B.n165 163.367
R417 B.n287 B.n286 163.367
R418 B.n288 B.n287 163.367
R419 B.n288 B.n163 163.367
R420 B.n292 B.n163 163.367
R421 B.n293 B.n292 163.367
R422 B.n294 B.n293 163.367
R423 B.n294 B.n161 163.367
R424 B.n298 B.n161 163.367
R425 B.n299 B.n298 163.367
R426 B.n300 B.n299 163.367
R427 B.n300 B.n159 163.367
R428 B.n304 B.n159 163.367
R429 B.n305 B.n304 163.367
R430 B.n306 B.n305 163.367
R431 B.n306 B.n157 163.367
R432 B.n310 B.n157 163.367
R433 B.n311 B.n310 163.367
R434 B.n312 B.n311 163.367
R435 B.n312 B.n155 163.367
R436 B.n316 B.n155 163.367
R437 B.n317 B.n316 163.367
R438 B.n318 B.n317 163.367
R439 B.n318 B.n153 163.367
R440 B.n322 B.n153 163.367
R441 B.n323 B.n322 163.367
R442 B.n324 B.n323 163.367
R443 B.n324 B.n149 163.367
R444 B.n329 B.n149 163.367
R445 B.n330 B.n329 163.367
R446 B.n331 B.n330 163.367
R447 B.n331 B.n147 163.367
R448 B.n335 B.n147 163.367
R449 B.n336 B.n335 163.367
R450 B.n337 B.n336 163.367
R451 B.n337 B.n145 163.367
R452 B.n344 B.n145 163.367
R453 B.n345 B.n344 163.367
R454 B.n346 B.n345 163.367
R455 B.n346 B.n143 163.367
R456 B.n350 B.n143 163.367
R457 B.n351 B.n350 163.367
R458 B.n352 B.n351 163.367
R459 B.n352 B.n141 163.367
R460 B.n356 B.n141 163.367
R461 B.n357 B.n356 163.367
R462 B.n358 B.n357 163.367
R463 B.n358 B.n139 163.367
R464 B.n362 B.n139 163.367
R465 B.n363 B.n362 163.367
R466 B.n364 B.n363 163.367
R467 B.n364 B.n137 163.367
R468 B.n368 B.n137 163.367
R469 B.n369 B.n368 163.367
R470 B.n370 B.n369 163.367
R471 B.n370 B.n135 163.367
R472 B.n374 B.n135 163.367
R473 B.n375 B.n374 163.367
R474 B.n376 B.n375 163.367
R475 B.n376 B.n133 163.367
R476 B.n380 B.n133 163.367
R477 B.n381 B.n380 163.367
R478 B.n382 B.n381 163.367
R479 B.n382 B.n131 163.367
R480 B.n386 B.n131 163.367
R481 B.n387 B.n386 163.367
R482 B.n388 B.n387 163.367
R483 B.n388 B.n129 163.367
R484 B.n392 B.n129 163.367
R485 B.n393 B.n392 163.367
R486 B.n394 B.n393 163.367
R487 B.n394 B.n127 163.367
R488 B.n398 B.n127 163.367
R489 B.n399 B.n398 163.367
R490 B.n400 B.n399 163.367
R491 B.n400 B.n125 163.367
R492 B.n404 B.n125 163.367
R493 B.n405 B.n404 163.367
R494 B.n406 B.n405 163.367
R495 B.n406 B.n123 163.367
R496 B.n410 B.n123 163.367
R497 B.n411 B.n410 163.367
R498 B.n412 B.n411 163.367
R499 B.n412 B.n121 163.367
R500 B.n416 B.n121 163.367
R501 B.n417 B.n416 163.367
R502 B.n418 B.n417 163.367
R503 B.n418 B.n119 163.367
R504 B.n422 B.n119 163.367
R505 B.n423 B.n422 163.367
R506 B.n424 B.n423 163.367
R507 B.n424 B.n117 163.367
R508 B.n526 B.n83 163.367
R509 B.n526 B.n525 163.367
R510 B.n525 B.n524 163.367
R511 B.n524 B.n85 163.367
R512 B.n520 B.n85 163.367
R513 B.n520 B.n519 163.367
R514 B.n519 B.n518 163.367
R515 B.n518 B.n87 163.367
R516 B.n514 B.n87 163.367
R517 B.n514 B.n513 163.367
R518 B.n513 B.n512 163.367
R519 B.n512 B.n89 163.367
R520 B.n508 B.n89 163.367
R521 B.n508 B.n507 163.367
R522 B.n507 B.n506 163.367
R523 B.n506 B.n91 163.367
R524 B.n502 B.n91 163.367
R525 B.n502 B.n501 163.367
R526 B.n501 B.n500 163.367
R527 B.n500 B.n93 163.367
R528 B.n496 B.n93 163.367
R529 B.n496 B.n495 163.367
R530 B.n495 B.n494 163.367
R531 B.n494 B.n95 163.367
R532 B.n490 B.n95 163.367
R533 B.n490 B.n489 163.367
R534 B.n489 B.n488 163.367
R535 B.n488 B.n97 163.367
R536 B.n484 B.n97 163.367
R537 B.n484 B.n483 163.367
R538 B.n483 B.n482 163.367
R539 B.n482 B.n99 163.367
R540 B.n478 B.n99 163.367
R541 B.n478 B.n477 163.367
R542 B.n477 B.n476 163.367
R543 B.n476 B.n101 163.367
R544 B.n472 B.n101 163.367
R545 B.n472 B.n471 163.367
R546 B.n471 B.n470 163.367
R547 B.n470 B.n103 163.367
R548 B.n466 B.n103 163.367
R549 B.n466 B.n465 163.367
R550 B.n465 B.n464 163.367
R551 B.n464 B.n105 163.367
R552 B.n460 B.n105 163.367
R553 B.n460 B.n459 163.367
R554 B.n459 B.n458 163.367
R555 B.n458 B.n107 163.367
R556 B.n454 B.n107 163.367
R557 B.n454 B.n453 163.367
R558 B.n453 B.n452 163.367
R559 B.n452 B.n109 163.367
R560 B.n448 B.n109 163.367
R561 B.n448 B.n447 163.367
R562 B.n447 B.n446 163.367
R563 B.n446 B.n111 163.367
R564 B.n442 B.n111 163.367
R565 B.n442 B.n441 163.367
R566 B.n441 B.n440 163.367
R567 B.n440 B.n113 163.367
R568 B.n436 B.n113 163.367
R569 B.n436 B.n435 163.367
R570 B.n435 B.n434 163.367
R571 B.n434 B.n115 163.367
R572 B.n430 B.n115 163.367
R573 B.n430 B.n429 163.367
R574 B.n429 B.n428 163.367
R575 B.n710 B.n19 163.367
R576 B.n706 B.n19 163.367
R577 B.n706 B.n705 163.367
R578 B.n705 B.n704 163.367
R579 B.n704 B.n21 163.367
R580 B.n700 B.n21 163.367
R581 B.n700 B.n699 163.367
R582 B.n699 B.n698 163.367
R583 B.n698 B.n23 163.367
R584 B.n694 B.n23 163.367
R585 B.n694 B.n693 163.367
R586 B.n693 B.n692 163.367
R587 B.n692 B.n25 163.367
R588 B.n688 B.n25 163.367
R589 B.n688 B.n687 163.367
R590 B.n687 B.n686 163.367
R591 B.n686 B.n27 163.367
R592 B.n682 B.n27 163.367
R593 B.n682 B.n681 163.367
R594 B.n681 B.n680 163.367
R595 B.n680 B.n29 163.367
R596 B.n676 B.n29 163.367
R597 B.n676 B.n675 163.367
R598 B.n675 B.n674 163.367
R599 B.n674 B.n31 163.367
R600 B.n670 B.n31 163.367
R601 B.n670 B.n669 163.367
R602 B.n669 B.n668 163.367
R603 B.n668 B.n33 163.367
R604 B.n664 B.n33 163.367
R605 B.n664 B.n663 163.367
R606 B.n663 B.n662 163.367
R607 B.n662 B.n35 163.367
R608 B.n658 B.n35 163.367
R609 B.n658 B.n657 163.367
R610 B.n657 B.n656 163.367
R611 B.n656 B.n37 163.367
R612 B.n652 B.n37 163.367
R613 B.n652 B.n651 163.367
R614 B.n651 B.n650 163.367
R615 B.n650 B.n39 163.367
R616 B.n646 B.n39 163.367
R617 B.n646 B.n645 163.367
R618 B.n645 B.n644 163.367
R619 B.n644 B.n41 163.367
R620 B.n640 B.n41 163.367
R621 B.n640 B.n639 163.367
R622 B.n639 B.n638 163.367
R623 B.n638 B.n43 163.367
R624 B.n634 B.n43 163.367
R625 B.n634 B.n633 163.367
R626 B.n633 B.n632 163.367
R627 B.n632 B.n45 163.367
R628 B.n628 B.n45 163.367
R629 B.n628 B.n627 163.367
R630 B.n627 B.n49 163.367
R631 B.n623 B.n49 163.367
R632 B.n623 B.n622 163.367
R633 B.n622 B.n621 163.367
R634 B.n621 B.n51 163.367
R635 B.n617 B.n51 163.367
R636 B.n617 B.n616 163.367
R637 B.n616 B.n615 163.367
R638 B.n615 B.n53 163.367
R639 B.n610 B.n53 163.367
R640 B.n610 B.n609 163.367
R641 B.n609 B.n608 163.367
R642 B.n608 B.n57 163.367
R643 B.n604 B.n57 163.367
R644 B.n604 B.n603 163.367
R645 B.n603 B.n602 163.367
R646 B.n602 B.n59 163.367
R647 B.n598 B.n59 163.367
R648 B.n598 B.n597 163.367
R649 B.n597 B.n596 163.367
R650 B.n596 B.n61 163.367
R651 B.n592 B.n61 163.367
R652 B.n592 B.n591 163.367
R653 B.n591 B.n590 163.367
R654 B.n590 B.n63 163.367
R655 B.n586 B.n63 163.367
R656 B.n586 B.n585 163.367
R657 B.n585 B.n584 163.367
R658 B.n584 B.n65 163.367
R659 B.n580 B.n65 163.367
R660 B.n580 B.n579 163.367
R661 B.n579 B.n578 163.367
R662 B.n578 B.n67 163.367
R663 B.n574 B.n67 163.367
R664 B.n574 B.n573 163.367
R665 B.n573 B.n572 163.367
R666 B.n572 B.n69 163.367
R667 B.n568 B.n69 163.367
R668 B.n568 B.n567 163.367
R669 B.n567 B.n566 163.367
R670 B.n566 B.n71 163.367
R671 B.n562 B.n71 163.367
R672 B.n562 B.n561 163.367
R673 B.n561 B.n560 163.367
R674 B.n560 B.n73 163.367
R675 B.n556 B.n73 163.367
R676 B.n556 B.n555 163.367
R677 B.n555 B.n554 163.367
R678 B.n554 B.n75 163.367
R679 B.n550 B.n75 163.367
R680 B.n550 B.n549 163.367
R681 B.n549 B.n548 163.367
R682 B.n548 B.n77 163.367
R683 B.n544 B.n77 163.367
R684 B.n544 B.n543 163.367
R685 B.n543 B.n542 163.367
R686 B.n542 B.n79 163.367
R687 B.n538 B.n79 163.367
R688 B.n538 B.n537 163.367
R689 B.n537 B.n536 163.367
R690 B.n536 B.n81 163.367
R691 B.n532 B.n81 163.367
R692 B.n532 B.n531 163.367
R693 B.n531 B.n530 163.367
R694 B.n712 B.n711 163.367
R695 B.n712 B.n17 163.367
R696 B.n716 B.n17 163.367
R697 B.n717 B.n716 163.367
R698 B.n718 B.n717 163.367
R699 B.n718 B.n15 163.367
R700 B.n722 B.n15 163.367
R701 B.n723 B.n722 163.367
R702 B.n724 B.n723 163.367
R703 B.n724 B.n13 163.367
R704 B.n728 B.n13 163.367
R705 B.n729 B.n728 163.367
R706 B.n730 B.n729 163.367
R707 B.n730 B.n11 163.367
R708 B.n734 B.n11 163.367
R709 B.n735 B.n734 163.367
R710 B.n736 B.n735 163.367
R711 B.n736 B.n9 163.367
R712 B.n740 B.n9 163.367
R713 B.n741 B.n740 163.367
R714 B.n742 B.n741 163.367
R715 B.n742 B.n7 163.367
R716 B.n746 B.n7 163.367
R717 B.n747 B.n746 163.367
R718 B.n748 B.n747 163.367
R719 B.n748 B.n5 163.367
R720 B.n752 B.n5 163.367
R721 B.n753 B.n752 163.367
R722 B.n754 B.n753 163.367
R723 B.n754 B.n3 163.367
R724 B.n758 B.n3 163.367
R725 B.n759 B.n758 163.367
R726 B.n196 B.n2 163.367
R727 B.n197 B.n196 163.367
R728 B.n198 B.n197 163.367
R729 B.n198 B.n193 163.367
R730 B.n202 B.n193 163.367
R731 B.n203 B.n202 163.367
R732 B.n204 B.n203 163.367
R733 B.n204 B.n191 163.367
R734 B.n208 B.n191 163.367
R735 B.n209 B.n208 163.367
R736 B.n210 B.n209 163.367
R737 B.n210 B.n189 163.367
R738 B.n214 B.n189 163.367
R739 B.n215 B.n214 163.367
R740 B.n216 B.n215 163.367
R741 B.n216 B.n187 163.367
R742 B.n220 B.n187 163.367
R743 B.n221 B.n220 163.367
R744 B.n222 B.n221 163.367
R745 B.n222 B.n185 163.367
R746 B.n226 B.n185 163.367
R747 B.n227 B.n226 163.367
R748 B.n228 B.n227 163.367
R749 B.n228 B.n183 163.367
R750 B.n232 B.n183 163.367
R751 B.n233 B.n232 163.367
R752 B.n234 B.n233 163.367
R753 B.n234 B.n181 163.367
R754 B.n238 B.n181 163.367
R755 B.n239 B.n238 163.367
R756 B.n240 B.n239 163.367
R757 B.n240 B.n179 163.367
R758 B.n341 B.t5 112.749
R759 B.n55 B.t10 112.749
R760 B.n151 B.t2 112.728
R761 B.n47 B.t7 112.728
R762 B.n326 B.n151 59.5399
R763 B.n342 B.n341 59.5399
R764 B.n612 B.n55 59.5399
R765 B.n48 B.n47 59.5399
R766 B.n151 B.n150 55.855
R767 B.n341 B.n340 55.855
R768 B.n55 B.n54 55.855
R769 B.n47 B.n46 55.855
R770 B.n709 B.n18 33.5615
R771 B.n529 B.n528 33.5615
R772 B.n427 B.n426 33.5615
R773 B.n243 B.n242 33.5615
R774 B B.n761 18.0485
R775 B.n713 B.n18 10.6151
R776 B.n714 B.n713 10.6151
R777 B.n715 B.n714 10.6151
R778 B.n715 B.n16 10.6151
R779 B.n719 B.n16 10.6151
R780 B.n720 B.n719 10.6151
R781 B.n721 B.n720 10.6151
R782 B.n721 B.n14 10.6151
R783 B.n725 B.n14 10.6151
R784 B.n726 B.n725 10.6151
R785 B.n727 B.n726 10.6151
R786 B.n727 B.n12 10.6151
R787 B.n731 B.n12 10.6151
R788 B.n732 B.n731 10.6151
R789 B.n733 B.n732 10.6151
R790 B.n733 B.n10 10.6151
R791 B.n737 B.n10 10.6151
R792 B.n738 B.n737 10.6151
R793 B.n739 B.n738 10.6151
R794 B.n739 B.n8 10.6151
R795 B.n743 B.n8 10.6151
R796 B.n744 B.n743 10.6151
R797 B.n745 B.n744 10.6151
R798 B.n745 B.n6 10.6151
R799 B.n749 B.n6 10.6151
R800 B.n750 B.n749 10.6151
R801 B.n751 B.n750 10.6151
R802 B.n751 B.n4 10.6151
R803 B.n755 B.n4 10.6151
R804 B.n756 B.n755 10.6151
R805 B.n757 B.n756 10.6151
R806 B.n757 B.n0 10.6151
R807 B.n709 B.n708 10.6151
R808 B.n708 B.n707 10.6151
R809 B.n707 B.n20 10.6151
R810 B.n703 B.n20 10.6151
R811 B.n703 B.n702 10.6151
R812 B.n702 B.n701 10.6151
R813 B.n701 B.n22 10.6151
R814 B.n697 B.n22 10.6151
R815 B.n697 B.n696 10.6151
R816 B.n696 B.n695 10.6151
R817 B.n695 B.n24 10.6151
R818 B.n691 B.n24 10.6151
R819 B.n691 B.n690 10.6151
R820 B.n690 B.n689 10.6151
R821 B.n689 B.n26 10.6151
R822 B.n685 B.n26 10.6151
R823 B.n685 B.n684 10.6151
R824 B.n684 B.n683 10.6151
R825 B.n683 B.n28 10.6151
R826 B.n679 B.n28 10.6151
R827 B.n679 B.n678 10.6151
R828 B.n678 B.n677 10.6151
R829 B.n677 B.n30 10.6151
R830 B.n673 B.n30 10.6151
R831 B.n673 B.n672 10.6151
R832 B.n672 B.n671 10.6151
R833 B.n671 B.n32 10.6151
R834 B.n667 B.n32 10.6151
R835 B.n667 B.n666 10.6151
R836 B.n666 B.n665 10.6151
R837 B.n665 B.n34 10.6151
R838 B.n661 B.n34 10.6151
R839 B.n661 B.n660 10.6151
R840 B.n660 B.n659 10.6151
R841 B.n659 B.n36 10.6151
R842 B.n655 B.n36 10.6151
R843 B.n655 B.n654 10.6151
R844 B.n654 B.n653 10.6151
R845 B.n653 B.n38 10.6151
R846 B.n649 B.n38 10.6151
R847 B.n649 B.n648 10.6151
R848 B.n648 B.n647 10.6151
R849 B.n647 B.n40 10.6151
R850 B.n643 B.n40 10.6151
R851 B.n643 B.n642 10.6151
R852 B.n642 B.n641 10.6151
R853 B.n641 B.n42 10.6151
R854 B.n637 B.n42 10.6151
R855 B.n637 B.n636 10.6151
R856 B.n636 B.n635 10.6151
R857 B.n635 B.n44 10.6151
R858 B.n631 B.n44 10.6151
R859 B.n631 B.n630 10.6151
R860 B.n630 B.n629 10.6151
R861 B.n626 B.n625 10.6151
R862 B.n625 B.n624 10.6151
R863 B.n624 B.n50 10.6151
R864 B.n620 B.n50 10.6151
R865 B.n620 B.n619 10.6151
R866 B.n619 B.n618 10.6151
R867 B.n618 B.n52 10.6151
R868 B.n614 B.n52 10.6151
R869 B.n614 B.n613 10.6151
R870 B.n611 B.n56 10.6151
R871 B.n607 B.n56 10.6151
R872 B.n607 B.n606 10.6151
R873 B.n606 B.n605 10.6151
R874 B.n605 B.n58 10.6151
R875 B.n601 B.n58 10.6151
R876 B.n601 B.n600 10.6151
R877 B.n600 B.n599 10.6151
R878 B.n599 B.n60 10.6151
R879 B.n595 B.n60 10.6151
R880 B.n595 B.n594 10.6151
R881 B.n594 B.n593 10.6151
R882 B.n593 B.n62 10.6151
R883 B.n589 B.n62 10.6151
R884 B.n589 B.n588 10.6151
R885 B.n588 B.n587 10.6151
R886 B.n587 B.n64 10.6151
R887 B.n583 B.n64 10.6151
R888 B.n583 B.n582 10.6151
R889 B.n582 B.n581 10.6151
R890 B.n581 B.n66 10.6151
R891 B.n577 B.n66 10.6151
R892 B.n577 B.n576 10.6151
R893 B.n576 B.n575 10.6151
R894 B.n575 B.n68 10.6151
R895 B.n571 B.n68 10.6151
R896 B.n571 B.n570 10.6151
R897 B.n570 B.n569 10.6151
R898 B.n569 B.n70 10.6151
R899 B.n565 B.n70 10.6151
R900 B.n565 B.n564 10.6151
R901 B.n564 B.n563 10.6151
R902 B.n563 B.n72 10.6151
R903 B.n559 B.n72 10.6151
R904 B.n559 B.n558 10.6151
R905 B.n558 B.n557 10.6151
R906 B.n557 B.n74 10.6151
R907 B.n553 B.n74 10.6151
R908 B.n553 B.n552 10.6151
R909 B.n552 B.n551 10.6151
R910 B.n551 B.n76 10.6151
R911 B.n547 B.n76 10.6151
R912 B.n547 B.n546 10.6151
R913 B.n546 B.n545 10.6151
R914 B.n545 B.n78 10.6151
R915 B.n541 B.n78 10.6151
R916 B.n541 B.n540 10.6151
R917 B.n540 B.n539 10.6151
R918 B.n539 B.n80 10.6151
R919 B.n535 B.n80 10.6151
R920 B.n535 B.n534 10.6151
R921 B.n534 B.n533 10.6151
R922 B.n533 B.n82 10.6151
R923 B.n529 B.n82 10.6151
R924 B.n528 B.n527 10.6151
R925 B.n527 B.n84 10.6151
R926 B.n523 B.n84 10.6151
R927 B.n523 B.n522 10.6151
R928 B.n522 B.n521 10.6151
R929 B.n521 B.n86 10.6151
R930 B.n517 B.n86 10.6151
R931 B.n517 B.n516 10.6151
R932 B.n516 B.n515 10.6151
R933 B.n515 B.n88 10.6151
R934 B.n511 B.n88 10.6151
R935 B.n511 B.n510 10.6151
R936 B.n510 B.n509 10.6151
R937 B.n509 B.n90 10.6151
R938 B.n505 B.n90 10.6151
R939 B.n505 B.n504 10.6151
R940 B.n504 B.n503 10.6151
R941 B.n503 B.n92 10.6151
R942 B.n499 B.n92 10.6151
R943 B.n499 B.n498 10.6151
R944 B.n498 B.n497 10.6151
R945 B.n497 B.n94 10.6151
R946 B.n493 B.n94 10.6151
R947 B.n493 B.n492 10.6151
R948 B.n492 B.n491 10.6151
R949 B.n491 B.n96 10.6151
R950 B.n487 B.n96 10.6151
R951 B.n487 B.n486 10.6151
R952 B.n486 B.n485 10.6151
R953 B.n485 B.n98 10.6151
R954 B.n481 B.n98 10.6151
R955 B.n481 B.n480 10.6151
R956 B.n480 B.n479 10.6151
R957 B.n479 B.n100 10.6151
R958 B.n475 B.n100 10.6151
R959 B.n475 B.n474 10.6151
R960 B.n474 B.n473 10.6151
R961 B.n473 B.n102 10.6151
R962 B.n469 B.n102 10.6151
R963 B.n469 B.n468 10.6151
R964 B.n468 B.n467 10.6151
R965 B.n467 B.n104 10.6151
R966 B.n463 B.n104 10.6151
R967 B.n463 B.n462 10.6151
R968 B.n462 B.n461 10.6151
R969 B.n461 B.n106 10.6151
R970 B.n457 B.n106 10.6151
R971 B.n457 B.n456 10.6151
R972 B.n456 B.n455 10.6151
R973 B.n455 B.n108 10.6151
R974 B.n451 B.n108 10.6151
R975 B.n451 B.n450 10.6151
R976 B.n450 B.n449 10.6151
R977 B.n449 B.n110 10.6151
R978 B.n445 B.n110 10.6151
R979 B.n445 B.n444 10.6151
R980 B.n444 B.n443 10.6151
R981 B.n443 B.n112 10.6151
R982 B.n439 B.n112 10.6151
R983 B.n439 B.n438 10.6151
R984 B.n438 B.n437 10.6151
R985 B.n437 B.n114 10.6151
R986 B.n433 B.n114 10.6151
R987 B.n433 B.n432 10.6151
R988 B.n432 B.n431 10.6151
R989 B.n431 B.n116 10.6151
R990 B.n427 B.n116 10.6151
R991 B.n195 B.n1 10.6151
R992 B.n195 B.n194 10.6151
R993 B.n199 B.n194 10.6151
R994 B.n200 B.n199 10.6151
R995 B.n201 B.n200 10.6151
R996 B.n201 B.n192 10.6151
R997 B.n205 B.n192 10.6151
R998 B.n206 B.n205 10.6151
R999 B.n207 B.n206 10.6151
R1000 B.n207 B.n190 10.6151
R1001 B.n211 B.n190 10.6151
R1002 B.n212 B.n211 10.6151
R1003 B.n213 B.n212 10.6151
R1004 B.n213 B.n188 10.6151
R1005 B.n217 B.n188 10.6151
R1006 B.n218 B.n217 10.6151
R1007 B.n219 B.n218 10.6151
R1008 B.n219 B.n186 10.6151
R1009 B.n223 B.n186 10.6151
R1010 B.n224 B.n223 10.6151
R1011 B.n225 B.n224 10.6151
R1012 B.n225 B.n184 10.6151
R1013 B.n229 B.n184 10.6151
R1014 B.n230 B.n229 10.6151
R1015 B.n231 B.n230 10.6151
R1016 B.n231 B.n182 10.6151
R1017 B.n235 B.n182 10.6151
R1018 B.n236 B.n235 10.6151
R1019 B.n237 B.n236 10.6151
R1020 B.n237 B.n180 10.6151
R1021 B.n241 B.n180 10.6151
R1022 B.n242 B.n241 10.6151
R1023 B.n243 B.n178 10.6151
R1024 B.n247 B.n178 10.6151
R1025 B.n248 B.n247 10.6151
R1026 B.n249 B.n248 10.6151
R1027 B.n249 B.n176 10.6151
R1028 B.n253 B.n176 10.6151
R1029 B.n254 B.n253 10.6151
R1030 B.n255 B.n254 10.6151
R1031 B.n255 B.n174 10.6151
R1032 B.n259 B.n174 10.6151
R1033 B.n260 B.n259 10.6151
R1034 B.n261 B.n260 10.6151
R1035 B.n261 B.n172 10.6151
R1036 B.n265 B.n172 10.6151
R1037 B.n266 B.n265 10.6151
R1038 B.n267 B.n266 10.6151
R1039 B.n267 B.n170 10.6151
R1040 B.n271 B.n170 10.6151
R1041 B.n272 B.n271 10.6151
R1042 B.n273 B.n272 10.6151
R1043 B.n273 B.n168 10.6151
R1044 B.n277 B.n168 10.6151
R1045 B.n278 B.n277 10.6151
R1046 B.n279 B.n278 10.6151
R1047 B.n279 B.n166 10.6151
R1048 B.n283 B.n166 10.6151
R1049 B.n284 B.n283 10.6151
R1050 B.n285 B.n284 10.6151
R1051 B.n285 B.n164 10.6151
R1052 B.n289 B.n164 10.6151
R1053 B.n290 B.n289 10.6151
R1054 B.n291 B.n290 10.6151
R1055 B.n291 B.n162 10.6151
R1056 B.n295 B.n162 10.6151
R1057 B.n296 B.n295 10.6151
R1058 B.n297 B.n296 10.6151
R1059 B.n297 B.n160 10.6151
R1060 B.n301 B.n160 10.6151
R1061 B.n302 B.n301 10.6151
R1062 B.n303 B.n302 10.6151
R1063 B.n303 B.n158 10.6151
R1064 B.n307 B.n158 10.6151
R1065 B.n308 B.n307 10.6151
R1066 B.n309 B.n308 10.6151
R1067 B.n309 B.n156 10.6151
R1068 B.n313 B.n156 10.6151
R1069 B.n314 B.n313 10.6151
R1070 B.n315 B.n314 10.6151
R1071 B.n315 B.n154 10.6151
R1072 B.n319 B.n154 10.6151
R1073 B.n320 B.n319 10.6151
R1074 B.n321 B.n320 10.6151
R1075 B.n321 B.n152 10.6151
R1076 B.n325 B.n152 10.6151
R1077 B.n328 B.n327 10.6151
R1078 B.n328 B.n148 10.6151
R1079 B.n332 B.n148 10.6151
R1080 B.n333 B.n332 10.6151
R1081 B.n334 B.n333 10.6151
R1082 B.n334 B.n146 10.6151
R1083 B.n338 B.n146 10.6151
R1084 B.n339 B.n338 10.6151
R1085 B.n343 B.n339 10.6151
R1086 B.n347 B.n144 10.6151
R1087 B.n348 B.n347 10.6151
R1088 B.n349 B.n348 10.6151
R1089 B.n349 B.n142 10.6151
R1090 B.n353 B.n142 10.6151
R1091 B.n354 B.n353 10.6151
R1092 B.n355 B.n354 10.6151
R1093 B.n355 B.n140 10.6151
R1094 B.n359 B.n140 10.6151
R1095 B.n360 B.n359 10.6151
R1096 B.n361 B.n360 10.6151
R1097 B.n361 B.n138 10.6151
R1098 B.n365 B.n138 10.6151
R1099 B.n366 B.n365 10.6151
R1100 B.n367 B.n366 10.6151
R1101 B.n367 B.n136 10.6151
R1102 B.n371 B.n136 10.6151
R1103 B.n372 B.n371 10.6151
R1104 B.n373 B.n372 10.6151
R1105 B.n373 B.n134 10.6151
R1106 B.n377 B.n134 10.6151
R1107 B.n378 B.n377 10.6151
R1108 B.n379 B.n378 10.6151
R1109 B.n379 B.n132 10.6151
R1110 B.n383 B.n132 10.6151
R1111 B.n384 B.n383 10.6151
R1112 B.n385 B.n384 10.6151
R1113 B.n385 B.n130 10.6151
R1114 B.n389 B.n130 10.6151
R1115 B.n390 B.n389 10.6151
R1116 B.n391 B.n390 10.6151
R1117 B.n391 B.n128 10.6151
R1118 B.n395 B.n128 10.6151
R1119 B.n396 B.n395 10.6151
R1120 B.n397 B.n396 10.6151
R1121 B.n397 B.n126 10.6151
R1122 B.n401 B.n126 10.6151
R1123 B.n402 B.n401 10.6151
R1124 B.n403 B.n402 10.6151
R1125 B.n403 B.n124 10.6151
R1126 B.n407 B.n124 10.6151
R1127 B.n408 B.n407 10.6151
R1128 B.n409 B.n408 10.6151
R1129 B.n409 B.n122 10.6151
R1130 B.n413 B.n122 10.6151
R1131 B.n414 B.n413 10.6151
R1132 B.n415 B.n414 10.6151
R1133 B.n415 B.n120 10.6151
R1134 B.n419 B.n120 10.6151
R1135 B.n420 B.n419 10.6151
R1136 B.n421 B.n420 10.6151
R1137 B.n421 B.n118 10.6151
R1138 B.n425 B.n118 10.6151
R1139 B.n426 B.n425 10.6151
R1140 B.n629 B.n48 9.36635
R1141 B.n612 B.n611 9.36635
R1142 B.n326 B.n325 9.36635
R1143 B.n342 B.n144 9.36635
R1144 B.n761 B.n0 8.11757
R1145 B.n761 B.n1 8.11757
R1146 B.n626 B.n48 1.24928
R1147 B.n613 B.n612 1.24928
R1148 B.n327 B.n326 1.24928
R1149 B.n343 B.n342 1.24928
R1150 VP.n4 VP.t2 193.179
R1151 VP.n4 VP.t1 192.411
R1152 VP.n14 VP.n0 161.3
R1153 VP.n13 VP.n12 161.3
R1154 VP.n11 VP.n1 161.3
R1155 VP.n10 VP.n9 161.3
R1156 VP.n8 VP.n2 161.3
R1157 VP.n7 VP.n6 161.3
R1158 VP.n3 VP.t0 157.359
R1159 VP.n15 VP.t3 157.359
R1160 VP.n5 VP.n3 101.459
R1161 VP.n16 VP.n15 101.459
R1162 VP.n9 VP.n1 56.5193
R1163 VP.n5 VP.n4 54.094
R1164 VP.n8 VP.n7 24.4675
R1165 VP.n9 VP.n8 24.4675
R1166 VP.n13 VP.n1 24.4675
R1167 VP.n14 VP.n13 24.4675
R1168 VP.n7 VP.n3 9.29796
R1169 VP.n15 VP.n14 9.29796
R1170 VP.n6 VP.n5 0.278367
R1171 VP.n16 VP.n0 0.278367
R1172 VP.n6 VP.n2 0.189894
R1173 VP.n10 VP.n2 0.189894
R1174 VP.n11 VP.n10 0.189894
R1175 VP.n12 VP.n11 0.189894
R1176 VP.n12 VP.n0 0.189894
R1177 VP VP.n16 0.153454
R1178 VDD1 VDD1.n1 119.706
R1179 VDD1 VDD1.n0 73.7222
R1180 VDD1.n0 VDD1.t0 1.95275
R1181 VDD1.n0 VDD1.t3 1.95275
R1182 VDD1.n1 VDD1.t2 1.95275
R1183 VDD1.n1 VDD1.t1 1.95275
R1184 VTAIL.n5 VTAIL.t5 58.9377
R1185 VTAIL.n4 VTAIL.t1 58.9377
R1186 VTAIL.n3 VTAIL.t2 58.9377
R1187 VTAIL.n7 VTAIL.t3 58.9374
R1188 VTAIL.n0 VTAIL.t0 58.9374
R1189 VTAIL.n1 VTAIL.t4 58.9374
R1190 VTAIL.n2 VTAIL.t7 58.9374
R1191 VTAIL.n6 VTAIL.t6 58.9374
R1192 VTAIL.n7 VTAIL.n6 29.2031
R1193 VTAIL.n3 VTAIL.n2 29.2031
R1194 VTAIL.n4 VTAIL.n3 2.48326
R1195 VTAIL.n6 VTAIL.n5 2.48326
R1196 VTAIL.n2 VTAIL.n1 2.48326
R1197 VTAIL VTAIL.n0 1.30007
R1198 VTAIL VTAIL.n7 1.18369
R1199 VTAIL.n5 VTAIL.n4 0.470328
R1200 VTAIL.n1 VTAIL.n0 0.470328
R1201 VN.n0 VN.t0 193.179
R1202 VN.n1 VN.t1 193.179
R1203 VN.n0 VN.t3 192.411
R1204 VN.n1 VN.t2 192.411
R1205 VN VN.n1 54.3728
R1206 VN VN.n0 4.42966
R1207 VDD2.n2 VDD2.n0 119.18
R1208 VDD2.n2 VDD2.n1 73.664
R1209 VDD2.n1 VDD2.t1 1.95275
R1210 VDD2.n1 VDD2.t2 1.95275
R1211 VDD2.n0 VDD2.t3 1.95275
R1212 VDD2.n0 VDD2.t0 1.95275
R1213 VDD2 VDD2.n2 0.0586897
C0 VP VDD1 6.68461f
C1 B VP 1.72888f
C2 VTAIL VDD1 6.51405f
C3 VN VDD1 0.149089f
C4 B VTAIL 6.4456f
C5 B VN 1.15376f
C6 w_n2698_n4298# VDD1 1.57122f
C7 VP VDD2 0.391258f
C8 B w_n2698_n4298# 10.488701f
C9 VTAIL VDD2 6.56792f
C10 VN VDD2 6.44317f
C11 B VDD1 1.37716f
C12 w_n2698_n4298# VDD2 1.62625f
C13 VP VTAIL 6.15662f
C14 VP VN 7.01598f
C15 VN VTAIL 6.14251f
C16 VDD1 VDD2 1.0102f
C17 w_n2698_n4298# VP 4.99158f
C18 B VDD2 1.42847f
C19 w_n2698_n4298# VTAIL 5.02102f
C20 w_n2698_n4298# VN 4.64487f
C21 VDD2 VSUBS 1.054986f
C22 VDD1 VSUBS 6.29955f
C23 VTAIL VSUBS 1.428698f
C24 VN VSUBS 5.5927f
C25 VP VSUBS 2.427145f
C26 B VSUBS 4.627097f
C27 w_n2698_n4298# VSUBS 0.141969p
C28 VDD2.t3 VSUBS 0.348884f
C29 VDD2.t0 VSUBS 0.348884f
C30 VDD2.n0 VSUBS 3.74362f
C31 VDD2.t1 VSUBS 0.348884f
C32 VDD2.t2 VSUBS 0.348884f
C33 VDD2.n1 VSUBS 2.88726f
C34 VDD2.n2 VSUBS 4.75574f
C35 VN.t0 VSUBS 3.81304f
C36 VN.t3 VSUBS 3.80748f
C37 VN.n0 VSUBS 2.45604f
C38 VN.t1 VSUBS 3.81304f
C39 VN.t2 VSUBS 3.80748f
C40 VN.n1 VSUBS 4.25866f
C41 VTAIL.t0 VSUBS 3.0331f
C42 VTAIL.n0 VSUBS 0.737018f
C43 VTAIL.t4 VSUBS 3.0331f
C44 VTAIL.n1 VSUBS 0.822593f
C45 VTAIL.t7 VSUBS 3.0331f
C46 VTAIL.n2 VSUBS 2.31121f
C47 VTAIL.t2 VSUBS 3.0331f
C48 VTAIL.n3 VSUBS 2.3112f
C49 VTAIL.t1 VSUBS 3.0331f
C50 VTAIL.n4 VSUBS 0.822589f
C51 VTAIL.t5 VSUBS 3.0331f
C52 VTAIL.n5 VSUBS 0.822589f
C53 VTAIL.t6 VSUBS 3.0331f
C54 VTAIL.n6 VSUBS 2.31121f
C55 VTAIL.t3 VSUBS 3.0331f
C56 VTAIL.n7 VSUBS 2.21721f
C57 VDD1.t0 VSUBS 0.351603f
C58 VDD1.t3 VSUBS 0.351603f
C59 VDD1.n0 VSUBS 2.91033f
C60 VDD1.t2 VSUBS 0.351603f
C61 VDD1.t1 VSUBS 0.351603f
C62 VDD1.n1 VSUBS 3.79919f
C63 VP.n0 VSUBS 0.041522f
C64 VP.t3 VSUBS 3.67238f
C65 VP.n1 VSUBS 0.045976f
C66 VP.n2 VSUBS 0.031494f
C67 VP.t0 VSUBS 3.67238f
C68 VP.n3 VSUBS 1.38042f
C69 VP.t1 VSUBS 3.94086f
C70 VP.t2 VSUBS 3.94662f
C71 VP.n4 VSUBS 4.39143f
C72 VP.n5 VSUBS 1.92534f
C73 VP.n6 VSUBS 0.041522f
C74 VP.n7 VSUBS 0.040731f
C75 VP.n8 VSUBS 0.058698f
C76 VP.n9 VSUBS 0.045976f
C77 VP.n10 VSUBS 0.031494f
C78 VP.n11 VSUBS 0.031494f
C79 VP.n12 VSUBS 0.031494f
C80 VP.n13 VSUBS 0.058698f
C81 VP.n14 VSUBS 0.040731f
C82 VP.n15 VSUBS 1.38042f
C83 VP.n16 VSUBS 0.051294f
C84 B.n0 VSUBS 0.005455f
C85 B.n1 VSUBS 0.005455f
C86 B.n2 VSUBS 0.008068f
C87 B.n3 VSUBS 0.006183f
C88 B.n4 VSUBS 0.006183f
C89 B.n5 VSUBS 0.006183f
C90 B.n6 VSUBS 0.006183f
C91 B.n7 VSUBS 0.006183f
C92 B.n8 VSUBS 0.006183f
C93 B.n9 VSUBS 0.006183f
C94 B.n10 VSUBS 0.006183f
C95 B.n11 VSUBS 0.006183f
C96 B.n12 VSUBS 0.006183f
C97 B.n13 VSUBS 0.006183f
C98 B.n14 VSUBS 0.006183f
C99 B.n15 VSUBS 0.006183f
C100 B.n16 VSUBS 0.006183f
C101 B.n17 VSUBS 0.006183f
C102 B.n18 VSUBS 0.014426f
C103 B.n19 VSUBS 0.006183f
C104 B.n20 VSUBS 0.006183f
C105 B.n21 VSUBS 0.006183f
C106 B.n22 VSUBS 0.006183f
C107 B.n23 VSUBS 0.006183f
C108 B.n24 VSUBS 0.006183f
C109 B.n25 VSUBS 0.006183f
C110 B.n26 VSUBS 0.006183f
C111 B.n27 VSUBS 0.006183f
C112 B.n28 VSUBS 0.006183f
C113 B.n29 VSUBS 0.006183f
C114 B.n30 VSUBS 0.006183f
C115 B.n31 VSUBS 0.006183f
C116 B.n32 VSUBS 0.006183f
C117 B.n33 VSUBS 0.006183f
C118 B.n34 VSUBS 0.006183f
C119 B.n35 VSUBS 0.006183f
C120 B.n36 VSUBS 0.006183f
C121 B.n37 VSUBS 0.006183f
C122 B.n38 VSUBS 0.006183f
C123 B.n39 VSUBS 0.006183f
C124 B.n40 VSUBS 0.006183f
C125 B.n41 VSUBS 0.006183f
C126 B.n42 VSUBS 0.006183f
C127 B.n43 VSUBS 0.006183f
C128 B.n44 VSUBS 0.006183f
C129 B.n45 VSUBS 0.006183f
C130 B.t7 VSUBS 0.493685f
C131 B.t8 VSUBS 0.511784f
C132 B.t6 VSUBS 1.66986f
C133 B.n46 VSUBS 0.275679f
C134 B.n47 VSUBS 0.063445f
C135 B.n48 VSUBS 0.014325f
C136 B.n49 VSUBS 0.006183f
C137 B.n50 VSUBS 0.006183f
C138 B.n51 VSUBS 0.006183f
C139 B.n52 VSUBS 0.006183f
C140 B.n53 VSUBS 0.006183f
C141 B.t10 VSUBS 0.493669f
C142 B.t11 VSUBS 0.511771f
C143 B.t9 VSUBS 1.66986f
C144 B.n54 VSUBS 0.275692f
C145 B.n55 VSUBS 0.06346f
C146 B.n56 VSUBS 0.006183f
C147 B.n57 VSUBS 0.006183f
C148 B.n58 VSUBS 0.006183f
C149 B.n59 VSUBS 0.006183f
C150 B.n60 VSUBS 0.006183f
C151 B.n61 VSUBS 0.006183f
C152 B.n62 VSUBS 0.006183f
C153 B.n63 VSUBS 0.006183f
C154 B.n64 VSUBS 0.006183f
C155 B.n65 VSUBS 0.006183f
C156 B.n66 VSUBS 0.006183f
C157 B.n67 VSUBS 0.006183f
C158 B.n68 VSUBS 0.006183f
C159 B.n69 VSUBS 0.006183f
C160 B.n70 VSUBS 0.006183f
C161 B.n71 VSUBS 0.006183f
C162 B.n72 VSUBS 0.006183f
C163 B.n73 VSUBS 0.006183f
C164 B.n74 VSUBS 0.006183f
C165 B.n75 VSUBS 0.006183f
C166 B.n76 VSUBS 0.006183f
C167 B.n77 VSUBS 0.006183f
C168 B.n78 VSUBS 0.006183f
C169 B.n79 VSUBS 0.006183f
C170 B.n80 VSUBS 0.006183f
C171 B.n81 VSUBS 0.006183f
C172 B.n82 VSUBS 0.006183f
C173 B.n83 VSUBS 0.014426f
C174 B.n84 VSUBS 0.006183f
C175 B.n85 VSUBS 0.006183f
C176 B.n86 VSUBS 0.006183f
C177 B.n87 VSUBS 0.006183f
C178 B.n88 VSUBS 0.006183f
C179 B.n89 VSUBS 0.006183f
C180 B.n90 VSUBS 0.006183f
C181 B.n91 VSUBS 0.006183f
C182 B.n92 VSUBS 0.006183f
C183 B.n93 VSUBS 0.006183f
C184 B.n94 VSUBS 0.006183f
C185 B.n95 VSUBS 0.006183f
C186 B.n96 VSUBS 0.006183f
C187 B.n97 VSUBS 0.006183f
C188 B.n98 VSUBS 0.006183f
C189 B.n99 VSUBS 0.006183f
C190 B.n100 VSUBS 0.006183f
C191 B.n101 VSUBS 0.006183f
C192 B.n102 VSUBS 0.006183f
C193 B.n103 VSUBS 0.006183f
C194 B.n104 VSUBS 0.006183f
C195 B.n105 VSUBS 0.006183f
C196 B.n106 VSUBS 0.006183f
C197 B.n107 VSUBS 0.006183f
C198 B.n108 VSUBS 0.006183f
C199 B.n109 VSUBS 0.006183f
C200 B.n110 VSUBS 0.006183f
C201 B.n111 VSUBS 0.006183f
C202 B.n112 VSUBS 0.006183f
C203 B.n113 VSUBS 0.006183f
C204 B.n114 VSUBS 0.006183f
C205 B.n115 VSUBS 0.006183f
C206 B.n116 VSUBS 0.006183f
C207 B.n117 VSUBS 0.015033f
C208 B.n118 VSUBS 0.006183f
C209 B.n119 VSUBS 0.006183f
C210 B.n120 VSUBS 0.006183f
C211 B.n121 VSUBS 0.006183f
C212 B.n122 VSUBS 0.006183f
C213 B.n123 VSUBS 0.006183f
C214 B.n124 VSUBS 0.006183f
C215 B.n125 VSUBS 0.006183f
C216 B.n126 VSUBS 0.006183f
C217 B.n127 VSUBS 0.006183f
C218 B.n128 VSUBS 0.006183f
C219 B.n129 VSUBS 0.006183f
C220 B.n130 VSUBS 0.006183f
C221 B.n131 VSUBS 0.006183f
C222 B.n132 VSUBS 0.006183f
C223 B.n133 VSUBS 0.006183f
C224 B.n134 VSUBS 0.006183f
C225 B.n135 VSUBS 0.006183f
C226 B.n136 VSUBS 0.006183f
C227 B.n137 VSUBS 0.006183f
C228 B.n138 VSUBS 0.006183f
C229 B.n139 VSUBS 0.006183f
C230 B.n140 VSUBS 0.006183f
C231 B.n141 VSUBS 0.006183f
C232 B.n142 VSUBS 0.006183f
C233 B.n143 VSUBS 0.006183f
C234 B.n144 VSUBS 0.005819f
C235 B.n145 VSUBS 0.006183f
C236 B.n146 VSUBS 0.006183f
C237 B.n147 VSUBS 0.006183f
C238 B.n148 VSUBS 0.006183f
C239 B.n149 VSUBS 0.006183f
C240 B.t2 VSUBS 0.493685f
C241 B.t1 VSUBS 0.511784f
C242 B.t0 VSUBS 1.66986f
C243 B.n150 VSUBS 0.275679f
C244 B.n151 VSUBS 0.063445f
C245 B.n152 VSUBS 0.006183f
C246 B.n153 VSUBS 0.006183f
C247 B.n154 VSUBS 0.006183f
C248 B.n155 VSUBS 0.006183f
C249 B.n156 VSUBS 0.006183f
C250 B.n157 VSUBS 0.006183f
C251 B.n158 VSUBS 0.006183f
C252 B.n159 VSUBS 0.006183f
C253 B.n160 VSUBS 0.006183f
C254 B.n161 VSUBS 0.006183f
C255 B.n162 VSUBS 0.006183f
C256 B.n163 VSUBS 0.006183f
C257 B.n164 VSUBS 0.006183f
C258 B.n165 VSUBS 0.006183f
C259 B.n166 VSUBS 0.006183f
C260 B.n167 VSUBS 0.006183f
C261 B.n168 VSUBS 0.006183f
C262 B.n169 VSUBS 0.006183f
C263 B.n170 VSUBS 0.006183f
C264 B.n171 VSUBS 0.006183f
C265 B.n172 VSUBS 0.006183f
C266 B.n173 VSUBS 0.006183f
C267 B.n174 VSUBS 0.006183f
C268 B.n175 VSUBS 0.006183f
C269 B.n176 VSUBS 0.006183f
C270 B.n177 VSUBS 0.006183f
C271 B.n178 VSUBS 0.006183f
C272 B.n179 VSUBS 0.014426f
C273 B.n180 VSUBS 0.006183f
C274 B.n181 VSUBS 0.006183f
C275 B.n182 VSUBS 0.006183f
C276 B.n183 VSUBS 0.006183f
C277 B.n184 VSUBS 0.006183f
C278 B.n185 VSUBS 0.006183f
C279 B.n186 VSUBS 0.006183f
C280 B.n187 VSUBS 0.006183f
C281 B.n188 VSUBS 0.006183f
C282 B.n189 VSUBS 0.006183f
C283 B.n190 VSUBS 0.006183f
C284 B.n191 VSUBS 0.006183f
C285 B.n192 VSUBS 0.006183f
C286 B.n193 VSUBS 0.006183f
C287 B.n194 VSUBS 0.006183f
C288 B.n195 VSUBS 0.006183f
C289 B.n196 VSUBS 0.006183f
C290 B.n197 VSUBS 0.006183f
C291 B.n198 VSUBS 0.006183f
C292 B.n199 VSUBS 0.006183f
C293 B.n200 VSUBS 0.006183f
C294 B.n201 VSUBS 0.006183f
C295 B.n202 VSUBS 0.006183f
C296 B.n203 VSUBS 0.006183f
C297 B.n204 VSUBS 0.006183f
C298 B.n205 VSUBS 0.006183f
C299 B.n206 VSUBS 0.006183f
C300 B.n207 VSUBS 0.006183f
C301 B.n208 VSUBS 0.006183f
C302 B.n209 VSUBS 0.006183f
C303 B.n210 VSUBS 0.006183f
C304 B.n211 VSUBS 0.006183f
C305 B.n212 VSUBS 0.006183f
C306 B.n213 VSUBS 0.006183f
C307 B.n214 VSUBS 0.006183f
C308 B.n215 VSUBS 0.006183f
C309 B.n216 VSUBS 0.006183f
C310 B.n217 VSUBS 0.006183f
C311 B.n218 VSUBS 0.006183f
C312 B.n219 VSUBS 0.006183f
C313 B.n220 VSUBS 0.006183f
C314 B.n221 VSUBS 0.006183f
C315 B.n222 VSUBS 0.006183f
C316 B.n223 VSUBS 0.006183f
C317 B.n224 VSUBS 0.006183f
C318 B.n225 VSUBS 0.006183f
C319 B.n226 VSUBS 0.006183f
C320 B.n227 VSUBS 0.006183f
C321 B.n228 VSUBS 0.006183f
C322 B.n229 VSUBS 0.006183f
C323 B.n230 VSUBS 0.006183f
C324 B.n231 VSUBS 0.006183f
C325 B.n232 VSUBS 0.006183f
C326 B.n233 VSUBS 0.006183f
C327 B.n234 VSUBS 0.006183f
C328 B.n235 VSUBS 0.006183f
C329 B.n236 VSUBS 0.006183f
C330 B.n237 VSUBS 0.006183f
C331 B.n238 VSUBS 0.006183f
C332 B.n239 VSUBS 0.006183f
C333 B.n240 VSUBS 0.006183f
C334 B.n241 VSUBS 0.006183f
C335 B.n242 VSUBS 0.014426f
C336 B.n243 VSUBS 0.015033f
C337 B.n244 VSUBS 0.015033f
C338 B.n245 VSUBS 0.006183f
C339 B.n246 VSUBS 0.006183f
C340 B.n247 VSUBS 0.006183f
C341 B.n248 VSUBS 0.006183f
C342 B.n249 VSUBS 0.006183f
C343 B.n250 VSUBS 0.006183f
C344 B.n251 VSUBS 0.006183f
C345 B.n252 VSUBS 0.006183f
C346 B.n253 VSUBS 0.006183f
C347 B.n254 VSUBS 0.006183f
C348 B.n255 VSUBS 0.006183f
C349 B.n256 VSUBS 0.006183f
C350 B.n257 VSUBS 0.006183f
C351 B.n258 VSUBS 0.006183f
C352 B.n259 VSUBS 0.006183f
C353 B.n260 VSUBS 0.006183f
C354 B.n261 VSUBS 0.006183f
C355 B.n262 VSUBS 0.006183f
C356 B.n263 VSUBS 0.006183f
C357 B.n264 VSUBS 0.006183f
C358 B.n265 VSUBS 0.006183f
C359 B.n266 VSUBS 0.006183f
C360 B.n267 VSUBS 0.006183f
C361 B.n268 VSUBS 0.006183f
C362 B.n269 VSUBS 0.006183f
C363 B.n270 VSUBS 0.006183f
C364 B.n271 VSUBS 0.006183f
C365 B.n272 VSUBS 0.006183f
C366 B.n273 VSUBS 0.006183f
C367 B.n274 VSUBS 0.006183f
C368 B.n275 VSUBS 0.006183f
C369 B.n276 VSUBS 0.006183f
C370 B.n277 VSUBS 0.006183f
C371 B.n278 VSUBS 0.006183f
C372 B.n279 VSUBS 0.006183f
C373 B.n280 VSUBS 0.006183f
C374 B.n281 VSUBS 0.006183f
C375 B.n282 VSUBS 0.006183f
C376 B.n283 VSUBS 0.006183f
C377 B.n284 VSUBS 0.006183f
C378 B.n285 VSUBS 0.006183f
C379 B.n286 VSUBS 0.006183f
C380 B.n287 VSUBS 0.006183f
C381 B.n288 VSUBS 0.006183f
C382 B.n289 VSUBS 0.006183f
C383 B.n290 VSUBS 0.006183f
C384 B.n291 VSUBS 0.006183f
C385 B.n292 VSUBS 0.006183f
C386 B.n293 VSUBS 0.006183f
C387 B.n294 VSUBS 0.006183f
C388 B.n295 VSUBS 0.006183f
C389 B.n296 VSUBS 0.006183f
C390 B.n297 VSUBS 0.006183f
C391 B.n298 VSUBS 0.006183f
C392 B.n299 VSUBS 0.006183f
C393 B.n300 VSUBS 0.006183f
C394 B.n301 VSUBS 0.006183f
C395 B.n302 VSUBS 0.006183f
C396 B.n303 VSUBS 0.006183f
C397 B.n304 VSUBS 0.006183f
C398 B.n305 VSUBS 0.006183f
C399 B.n306 VSUBS 0.006183f
C400 B.n307 VSUBS 0.006183f
C401 B.n308 VSUBS 0.006183f
C402 B.n309 VSUBS 0.006183f
C403 B.n310 VSUBS 0.006183f
C404 B.n311 VSUBS 0.006183f
C405 B.n312 VSUBS 0.006183f
C406 B.n313 VSUBS 0.006183f
C407 B.n314 VSUBS 0.006183f
C408 B.n315 VSUBS 0.006183f
C409 B.n316 VSUBS 0.006183f
C410 B.n317 VSUBS 0.006183f
C411 B.n318 VSUBS 0.006183f
C412 B.n319 VSUBS 0.006183f
C413 B.n320 VSUBS 0.006183f
C414 B.n321 VSUBS 0.006183f
C415 B.n322 VSUBS 0.006183f
C416 B.n323 VSUBS 0.006183f
C417 B.n324 VSUBS 0.006183f
C418 B.n325 VSUBS 0.005819f
C419 B.n326 VSUBS 0.014325f
C420 B.n327 VSUBS 0.003455f
C421 B.n328 VSUBS 0.006183f
C422 B.n329 VSUBS 0.006183f
C423 B.n330 VSUBS 0.006183f
C424 B.n331 VSUBS 0.006183f
C425 B.n332 VSUBS 0.006183f
C426 B.n333 VSUBS 0.006183f
C427 B.n334 VSUBS 0.006183f
C428 B.n335 VSUBS 0.006183f
C429 B.n336 VSUBS 0.006183f
C430 B.n337 VSUBS 0.006183f
C431 B.n338 VSUBS 0.006183f
C432 B.n339 VSUBS 0.006183f
C433 B.t5 VSUBS 0.493669f
C434 B.t4 VSUBS 0.511771f
C435 B.t3 VSUBS 1.66986f
C436 B.n340 VSUBS 0.275692f
C437 B.n341 VSUBS 0.06346f
C438 B.n342 VSUBS 0.014325f
C439 B.n343 VSUBS 0.003455f
C440 B.n344 VSUBS 0.006183f
C441 B.n345 VSUBS 0.006183f
C442 B.n346 VSUBS 0.006183f
C443 B.n347 VSUBS 0.006183f
C444 B.n348 VSUBS 0.006183f
C445 B.n349 VSUBS 0.006183f
C446 B.n350 VSUBS 0.006183f
C447 B.n351 VSUBS 0.006183f
C448 B.n352 VSUBS 0.006183f
C449 B.n353 VSUBS 0.006183f
C450 B.n354 VSUBS 0.006183f
C451 B.n355 VSUBS 0.006183f
C452 B.n356 VSUBS 0.006183f
C453 B.n357 VSUBS 0.006183f
C454 B.n358 VSUBS 0.006183f
C455 B.n359 VSUBS 0.006183f
C456 B.n360 VSUBS 0.006183f
C457 B.n361 VSUBS 0.006183f
C458 B.n362 VSUBS 0.006183f
C459 B.n363 VSUBS 0.006183f
C460 B.n364 VSUBS 0.006183f
C461 B.n365 VSUBS 0.006183f
C462 B.n366 VSUBS 0.006183f
C463 B.n367 VSUBS 0.006183f
C464 B.n368 VSUBS 0.006183f
C465 B.n369 VSUBS 0.006183f
C466 B.n370 VSUBS 0.006183f
C467 B.n371 VSUBS 0.006183f
C468 B.n372 VSUBS 0.006183f
C469 B.n373 VSUBS 0.006183f
C470 B.n374 VSUBS 0.006183f
C471 B.n375 VSUBS 0.006183f
C472 B.n376 VSUBS 0.006183f
C473 B.n377 VSUBS 0.006183f
C474 B.n378 VSUBS 0.006183f
C475 B.n379 VSUBS 0.006183f
C476 B.n380 VSUBS 0.006183f
C477 B.n381 VSUBS 0.006183f
C478 B.n382 VSUBS 0.006183f
C479 B.n383 VSUBS 0.006183f
C480 B.n384 VSUBS 0.006183f
C481 B.n385 VSUBS 0.006183f
C482 B.n386 VSUBS 0.006183f
C483 B.n387 VSUBS 0.006183f
C484 B.n388 VSUBS 0.006183f
C485 B.n389 VSUBS 0.006183f
C486 B.n390 VSUBS 0.006183f
C487 B.n391 VSUBS 0.006183f
C488 B.n392 VSUBS 0.006183f
C489 B.n393 VSUBS 0.006183f
C490 B.n394 VSUBS 0.006183f
C491 B.n395 VSUBS 0.006183f
C492 B.n396 VSUBS 0.006183f
C493 B.n397 VSUBS 0.006183f
C494 B.n398 VSUBS 0.006183f
C495 B.n399 VSUBS 0.006183f
C496 B.n400 VSUBS 0.006183f
C497 B.n401 VSUBS 0.006183f
C498 B.n402 VSUBS 0.006183f
C499 B.n403 VSUBS 0.006183f
C500 B.n404 VSUBS 0.006183f
C501 B.n405 VSUBS 0.006183f
C502 B.n406 VSUBS 0.006183f
C503 B.n407 VSUBS 0.006183f
C504 B.n408 VSUBS 0.006183f
C505 B.n409 VSUBS 0.006183f
C506 B.n410 VSUBS 0.006183f
C507 B.n411 VSUBS 0.006183f
C508 B.n412 VSUBS 0.006183f
C509 B.n413 VSUBS 0.006183f
C510 B.n414 VSUBS 0.006183f
C511 B.n415 VSUBS 0.006183f
C512 B.n416 VSUBS 0.006183f
C513 B.n417 VSUBS 0.006183f
C514 B.n418 VSUBS 0.006183f
C515 B.n419 VSUBS 0.006183f
C516 B.n420 VSUBS 0.006183f
C517 B.n421 VSUBS 0.006183f
C518 B.n422 VSUBS 0.006183f
C519 B.n423 VSUBS 0.006183f
C520 B.n424 VSUBS 0.006183f
C521 B.n425 VSUBS 0.006183f
C522 B.n426 VSUBS 0.014322f
C523 B.n427 VSUBS 0.015137f
C524 B.n428 VSUBS 0.014426f
C525 B.n429 VSUBS 0.006183f
C526 B.n430 VSUBS 0.006183f
C527 B.n431 VSUBS 0.006183f
C528 B.n432 VSUBS 0.006183f
C529 B.n433 VSUBS 0.006183f
C530 B.n434 VSUBS 0.006183f
C531 B.n435 VSUBS 0.006183f
C532 B.n436 VSUBS 0.006183f
C533 B.n437 VSUBS 0.006183f
C534 B.n438 VSUBS 0.006183f
C535 B.n439 VSUBS 0.006183f
C536 B.n440 VSUBS 0.006183f
C537 B.n441 VSUBS 0.006183f
C538 B.n442 VSUBS 0.006183f
C539 B.n443 VSUBS 0.006183f
C540 B.n444 VSUBS 0.006183f
C541 B.n445 VSUBS 0.006183f
C542 B.n446 VSUBS 0.006183f
C543 B.n447 VSUBS 0.006183f
C544 B.n448 VSUBS 0.006183f
C545 B.n449 VSUBS 0.006183f
C546 B.n450 VSUBS 0.006183f
C547 B.n451 VSUBS 0.006183f
C548 B.n452 VSUBS 0.006183f
C549 B.n453 VSUBS 0.006183f
C550 B.n454 VSUBS 0.006183f
C551 B.n455 VSUBS 0.006183f
C552 B.n456 VSUBS 0.006183f
C553 B.n457 VSUBS 0.006183f
C554 B.n458 VSUBS 0.006183f
C555 B.n459 VSUBS 0.006183f
C556 B.n460 VSUBS 0.006183f
C557 B.n461 VSUBS 0.006183f
C558 B.n462 VSUBS 0.006183f
C559 B.n463 VSUBS 0.006183f
C560 B.n464 VSUBS 0.006183f
C561 B.n465 VSUBS 0.006183f
C562 B.n466 VSUBS 0.006183f
C563 B.n467 VSUBS 0.006183f
C564 B.n468 VSUBS 0.006183f
C565 B.n469 VSUBS 0.006183f
C566 B.n470 VSUBS 0.006183f
C567 B.n471 VSUBS 0.006183f
C568 B.n472 VSUBS 0.006183f
C569 B.n473 VSUBS 0.006183f
C570 B.n474 VSUBS 0.006183f
C571 B.n475 VSUBS 0.006183f
C572 B.n476 VSUBS 0.006183f
C573 B.n477 VSUBS 0.006183f
C574 B.n478 VSUBS 0.006183f
C575 B.n479 VSUBS 0.006183f
C576 B.n480 VSUBS 0.006183f
C577 B.n481 VSUBS 0.006183f
C578 B.n482 VSUBS 0.006183f
C579 B.n483 VSUBS 0.006183f
C580 B.n484 VSUBS 0.006183f
C581 B.n485 VSUBS 0.006183f
C582 B.n486 VSUBS 0.006183f
C583 B.n487 VSUBS 0.006183f
C584 B.n488 VSUBS 0.006183f
C585 B.n489 VSUBS 0.006183f
C586 B.n490 VSUBS 0.006183f
C587 B.n491 VSUBS 0.006183f
C588 B.n492 VSUBS 0.006183f
C589 B.n493 VSUBS 0.006183f
C590 B.n494 VSUBS 0.006183f
C591 B.n495 VSUBS 0.006183f
C592 B.n496 VSUBS 0.006183f
C593 B.n497 VSUBS 0.006183f
C594 B.n498 VSUBS 0.006183f
C595 B.n499 VSUBS 0.006183f
C596 B.n500 VSUBS 0.006183f
C597 B.n501 VSUBS 0.006183f
C598 B.n502 VSUBS 0.006183f
C599 B.n503 VSUBS 0.006183f
C600 B.n504 VSUBS 0.006183f
C601 B.n505 VSUBS 0.006183f
C602 B.n506 VSUBS 0.006183f
C603 B.n507 VSUBS 0.006183f
C604 B.n508 VSUBS 0.006183f
C605 B.n509 VSUBS 0.006183f
C606 B.n510 VSUBS 0.006183f
C607 B.n511 VSUBS 0.006183f
C608 B.n512 VSUBS 0.006183f
C609 B.n513 VSUBS 0.006183f
C610 B.n514 VSUBS 0.006183f
C611 B.n515 VSUBS 0.006183f
C612 B.n516 VSUBS 0.006183f
C613 B.n517 VSUBS 0.006183f
C614 B.n518 VSUBS 0.006183f
C615 B.n519 VSUBS 0.006183f
C616 B.n520 VSUBS 0.006183f
C617 B.n521 VSUBS 0.006183f
C618 B.n522 VSUBS 0.006183f
C619 B.n523 VSUBS 0.006183f
C620 B.n524 VSUBS 0.006183f
C621 B.n525 VSUBS 0.006183f
C622 B.n526 VSUBS 0.006183f
C623 B.n527 VSUBS 0.006183f
C624 B.n528 VSUBS 0.014426f
C625 B.n529 VSUBS 0.015033f
C626 B.n530 VSUBS 0.015033f
C627 B.n531 VSUBS 0.006183f
C628 B.n532 VSUBS 0.006183f
C629 B.n533 VSUBS 0.006183f
C630 B.n534 VSUBS 0.006183f
C631 B.n535 VSUBS 0.006183f
C632 B.n536 VSUBS 0.006183f
C633 B.n537 VSUBS 0.006183f
C634 B.n538 VSUBS 0.006183f
C635 B.n539 VSUBS 0.006183f
C636 B.n540 VSUBS 0.006183f
C637 B.n541 VSUBS 0.006183f
C638 B.n542 VSUBS 0.006183f
C639 B.n543 VSUBS 0.006183f
C640 B.n544 VSUBS 0.006183f
C641 B.n545 VSUBS 0.006183f
C642 B.n546 VSUBS 0.006183f
C643 B.n547 VSUBS 0.006183f
C644 B.n548 VSUBS 0.006183f
C645 B.n549 VSUBS 0.006183f
C646 B.n550 VSUBS 0.006183f
C647 B.n551 VSUBS 0.006183f
C648 B.n552 VSUBS 0.006183f
C649 B.n553 VSUBS 0.006183f
C650 B.n554 VSUBS 0.006183f
C651 B.n555 VSUBS 0.006183f
C652 B.n556 VSUBS 0.006183f
C653 B.n557 VSUBS 0.006183f
C654 B.n558 VSUBS 0.006183f
C655 B.n559 VSUBS 0.006183f
C656 B.n560 VSUBS 0.006183f
C657 B.n561 VSUBS 0.006183f
C658 B.n562 VSUBS 0.006183f
C659 B.n563 VSUBS 0.006183f
C660 B.n564 VSUBS 0.006183f
C661 B.n565 VSUBS 0.006183f
C662 B.n566 VSUBS 0.006183f
C663 B.n567 VSUBS 0.006183f
C664 B.n568 VSUBS 0.006183f
C665 B.n569 VSUBS 0.006183f
C666 B.n570 VSUBS 0.006183f
C667 B.n571 VSUBS 0.006183f
C668 B.n572 VSUBS 0.006183f
C669 B.n573 VSUBS 0.006183f
C670 B.n574 VSUBS 0.006183f
C671 B.n575 VSUBS 0.006183f
C672 B.n576 VSUBS 0.006183f
C673 B.n577 VSUBS 0.006183f
C674 B.n578 VSUBS 0.006183f
C675 B.n579 VSUBS 0.006183f
C676 B.n580 VSUBS 0.006183f
C677 B.n581 VSUBS 0.006183f
C678 B.n582 VSUBS 0.006183f
C679 B.n583 VSUBS 0.006183f
C680 B.n584 VSUBS 0.006183f
C681 B.n585 VSUBS 0.006183f
C682 B.n586 VSUBS 0.006183f
C683 B.n587 VSUBS 0.006183f
C684 B.n588 VSUBS 0.006183f
C685 B.n589 VSUBS 0.006183f
C686 B.n590 VSUBS 0.006183f
C687 B.n591 VSUBS 0.006183f
C688 B.n592 VSUBS 0.006183f
C689 B.n593 VSUBS 0.006183f
C690 B.n594 VSUBS 0.006183f
C691 B.n595 VSUBS 0.006183f
C692 B.n596 VSUBS 0.006183f
C693 B.n597 VSUBS 0.006183f
C694 B.n598 VSUBS 0.006183f
C695 B.n599 VSUBS 0.006183f
C696 B.n600 VSUBS 0.006183f
C697 B.n601 VSUBS 0.006183f
C698 B.n602 VSUBS 0.006183f
C699 B.n603 VSUBS 0.006183f
C700 B.n604 VSUBS 0.006183f
C701 B.n605 VSUBS 0.006183f
C702 B.n606 VSUBS 0.006183f
C703 B.n607 VSUBS 0.006183f
C704 B.n608 VSUBS 0.006183f
C705 B.n609 VSUBS 0.006183f
C706 B.n610 VSUBS 0.006183f
C707 B.n611 VSUBS 0.005819f
C708 B.n612 VSUBS 0.014325f
C709 B.n613 VSUBS 0.003455f
C710 B.n614 VSUBS 0.006183f
C711 B.n615 VSUBS 0.006183f
C712 B.n616 VSUBS 0.006183f
C713 B.n617 VSUBS 0.006183f
C714 B.n618 VSUBS 0.006183f
C715 B.n619 VSUBS 0.006183f
C716 B.n620 VSUBS 0.006183f
C717 B.n621 VSUBS 0.006183f
C718 B.n622 VSUBS 0.006183f
C719 B.n623 VSUBS 0.006183f
C720 B.n624 VSUBS 0.006183f
C721 B.n625 VSUBS 0.006183f
C722 B.n626 VSUBS 0.003455f
C723 B.n627 VSUBS 0.006183f
C724 B.n628 VSUBS 0.006183f
C725 B.n629 VSUBS 0.005819f
C726 B.n630 VSUBS 0.006183f
C727 B.n631 VSUBS 0.006183f
C728 B.n632 VSUBS 0.006183f
C729 B.n633 VSUBS 0.006183f
C730 B.n634 VSUBS 0.006183f
C731 B.n635 VSUBS 0.006183f
C732 B.n636 VSUBS 0.006183f
C733 B.n637 VSUBS 0.006183f
C734 B.n638 VSUBS 0.006183f
C735 B.n639 VSUBS 0.006183f
C736 B.n640 VSUBS 0.006183f
C737 B.n641 VSUBS 0.006183f
C738 B.n642 VSUBS 0.006183f
C739 B.n643 VSUBS 0.006183f
C740 B.n644 VSUBS 0.006183f
C741 B.n645 VSUBS 0.006183f
C742 B.n646 VSUBS 0.006183f
C743 B.n647 VSUBS 0.006183f
C744 B.n648 VSUBS 0.006183f
C745 B.n649 VSUBS 0.006183f
C746 B.n650 VSUBS 0.006183f
C747 B.n651 VSUBS 0.006183f
C748 B.n652 VSUBS 0.006183f
C749 B.n653 VSUBS 0.006183f
C750 B.n654 VSUBS 0.006183f
C751 B.n655 VSUBS 0.006183f
C752 B.n656 VSUBS 0.006183f
C753 B.n657 VSUBS 0.006183f
C754 B.n658 VSUBS 0.006183f
C755 B.n659 VSUBS 0.006183f
C756 B.n660 VSUBS 0.006183f
C757 B.n661 VSUBS 0.006183f
C758 B.n662 VSUBS 0.006183f
C759 B.n663 VSUBS 0.006183f
C760 B.n664 VSUBS 0.006183f
C761 B.n665 VSUBS 0.006183f
C762 B.n666 VSUBS 0.006183f
C763 B.n667 VSUBS 0.006183f
C764 B.n668 VSUBS 0.006183f
C765 B.n669 VSUBS 0.006183f
C766 B.n670 VSUBS 0.006183f
C767 B.n671 VSUBS 0.006183f
C768 B.n672 VSUBS 0.006183f
C769 B.n673 VSUBS 0.006183f
C770 B.n674 VSUBS 0.006183f
C771 B.n675 VSUBS 0.006183f
C772 B.n676 VSUBS 0.006183f
C773 B.n677 VSUBS 0.006183f
C774 B.n678 VSUBS 0.006183f
C775 B.n679 VSUBS 0.006183f
C776 B.n680 VSUBS 0.006183f
C777 B.n681 VSUBS 0.006183f
C778 B.n682 VSUBS 0.006183f
C779 B.n683 VSUBS 0.006183f
C780 B.n684 VSUBS 0.006183f
C781 B.n685 VSUBS 0.006183f
C782 B.n686 VSUBS 0.006183f
C783 B.n687 VSUBS 0.006183f
C784 B.n688 VSUBS 0.006183f
C785 B.n689 VSUBS 0.006183f
C786 B.n690 VSUBS 0.006183f
C787 B.n691 VSUBS 0.006183f
C788 B.n692 VSUBS 0.006183f
C789 B.n693 VSUBS 0.006183f
C790 B.n694 VSUBS 0.006183f
C791 B.n695 VSUBS 0.006183f
C792 B.n696 VSUBS 0.006183f
C793 B.n697 VSUBS 0.006183f
C794 B.n698 VSUBS 0.006183f
C795 B.n699 VSUBS 0.006183f
C796 B.n700 VSUBS 0.006183f
C797 B.n701 VSUBS 0.006183f
C798 B.n702 VSUBS 0.006183f
C799 B.n703 VSUBS 0.006183f
C800 B.n704 VSUBS 0.006183f
C801 B.n705 VSUBS 0.006183f
C802 B.n706 VSUBS 0.006183f
C803 B.n707 VSUBS 0.006183f
C804 B.n708 VSUBS 0.006183f
C805 B.n709 VSUBS 0.015033f
C806 B.n710 VSUBS 0.015033f
C807 B.n711 VSUBS 0.014426f
C808 B.n712 VSUBS 0.006183f
C809 B.n713 VSUBS 0.006183f
C810 B.n714 VSUBS 0.006183f
C811 B.n715 VSUBS 0.006183f
C812 B.n716 VSUBS 0.006183f
C813 B.n717 VSUBS 0.006183f
C814 B.n718 VSUBS 0.006183f
C815 B.n719 VSUBS 0.006183f
C816 B.n720 VSUBS 0.006183f
C817 B.n721 VSUBS 0.006183f
C818 B.n722 VSUBS 0.006183f
C819 B.n723 VSUBS 0.006183f
C820 B.n724 VSUBS 0.006183f
C821 B.n725 VSUBS 0.006183f
C822 B.n726 VSUBS 0.006183f
C823 B.n727 VSUBS 0.006183f
C824 B.n728 VSUBS 0.006183f
C825 B.n729 VSUBS 0.006183f
C826 B.n730 VSUBS 0.006183f
C827 B.n731 VSUBS 0.006183f
C828 B.n732 VSUBS 0.006183f
C829 B.n733 VSUBS 0.006183f
C830 B.n734 VSUBS 0.006183f
C831 B.n735 VSUBS 0.006183f
C832 B.n736 VSUBS 0.006183f
C833 B.n737 VSUBS 0.006183f
C834 B.n738 VSUBS 0.006183f
C835 B.n739 VSUBS 0.006183f
C836 B.n740 VSUBS 0.006183f
C837 B.n741 VSUBS 0.006183f
C838 B.n742 VSUBS 0.006183f
C839 B.n743 VSUBS 0.006183f
C840 B.n744 VSUBS 0.006183f
C841 B.n745 VSUBS 0.006183f
C842 B.n746 VSUBS 0.006183f
C843 B.n747 VSUBS 0.006183f
C844 B.n748 VSUBS 0.006183f
C845 B.n749 VSUBS 0.006183f
C846 B.n750 VSUBS 0.006183f
C847 B.n751 VSUBS 0.006183f
C848 B.n752 VSUBS 0.006183f
C849 B.n753 VSUBS 0.006183f
C850 B.n754 VSUBS 0.006183f
C851 B.n755 VSUBS 0.006183f
C852 B.n756 VSUBS 0.006183f
C853 B.n757 VSUBS 0.006183f
C854 B.n758 VSUBS 0.006183f
C855 B.n759 VSUBS 0.008068f
C856 B.n760 VSUBS 0.008595f
C857 B.n761 VSUBS 0.017091f
.ends

