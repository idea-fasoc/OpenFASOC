* NGSPICE file created from diff_pair_sample_1049.ext - technology: sky130A

.subckt diff_pair_sample_1049 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t19 B.t22 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X1 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=2.96
X2 VTAIL.t6 VN.t0 VDD2.t9 B.t20 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X3 VDD2.t8 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=2.96
X4 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=2.96
X5 VDD1.t8 VP.t1 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=2.96
X6 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=2.96
X7 VTAIL.t17 VP.t2 VDD1.t7 B.t20 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X8 VTAIL.t5 VN.t2 VDD2.t7 B.t19 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X9 VTAIL.t1 VN.t3 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X10 VTAIL.t13 VP.t3 VDD1.t6 B.t19 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X11 VDD1.t5 VP.t4 VTAIL.t16 B.t23 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=2.96
X12 VDD1.t4 VP.t5 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=2.96
X13 VDD2.t5 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X14 VDD1.t3 VP.t6 VTAIL.t12 B.t21 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=2.96
X15 VTAIL.t14 VP.t7 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X16 VDD2.t4 VN.t5 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=2.96
X17 VDD2.t3 VN.t6 VTAIL.t8 B.t22 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X18 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=0 ps=0 w=13.7 l=2.96
X19 VDD1.t1 VP.t8 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X20 VDD2.t2 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.343 pd=28.18 as=2.2605 ps=14.03 w=13.7 l=2.96
X21 VTAIL.t15 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X22 VTAIL.t2 VN.t8 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=2.2605 ps=14.03 w=13.7 l=2.96
X23 VDD2.t0 VN.t9 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=2.2605 pd=14.03 as=5.343 ps=28.18 w=13.7 l=2.96
R0 VP.n27 VP.n24 161.3
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n23 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n22 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n21 161.3
R7 VP.n39 VP.n38 161.3
R8 VP.n40 VP.n20 161.3
R9 VP.n42 VP.n41 161.3
R10 VP.n43 VP.n19 161.3
R11 VP.n45 VP.n44 161.3
R12 VP.n46 VP.n18 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n50 VP.n17 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n16 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n15 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n93 VP.n92 161.3
R27 VP.n91 VP.n4 161.3
R28 VP.n90 VP.n89 161.3
R29 VP.n88 VP.n5 161.3
R30 VP.n87 VP.n86 161.3
R31 VP.n85 VP.n6 161.3
R32 VP.n84 VP.n83 161.3
R33 VP.n81 VP.n7 161.3
R34 VP.n80 VP.n79 161.3
R35 VP.n78 VP.n8 161.3
R36 VP.n77 VP.n76 161.3
R37 VP.n75 VP.n9 161.3
R38 VP.n74 VP.n73 161.3
R39 VP.n72 VP.n10 161.3
R40 VP.n71 VP.n70 161.3
R41 VP.n68 VP.n11 161.3
R42 VP.n67 VP.n66 161.3
R43 VP.n65 VP.n12 161.3
R44 VP.n64 VP.n63 161.3
R45 VP.n62 VP.n13 161.3
R46 VP.n26 VP.t1 143.061
R47 VP.n61 VP.t5 111.544
R48 VP.n69 VP.t9 111.544
R49 VP.n82 VP.t0 111.544
R50 VP.n94 VP.t2 111.544
R51 VP.n0 VP.t4 111.544
R52 VP.n14 VP.t6 111.544
R53 VP.n49 VP.t3 111.544
R54 VP.n37 VP.t8 111.544
R55 VP.n25 VP.t7 111.544
R56 VP.n61 VP.n60 74.0149
R57 VP.n104 VP.n0 74.0149
R58 VP.n59 VP.n14 74.0149
R59 VP.n26 VP.n25 71.6401
R60 VP.n67 VP.n12 56.5617
R61 VP.n100 VP.n2 56.5617
R62 VP.n55 VP.n16 56.5617
R63 VP.n60 VP.n59 56.4124
R64 VP.n76 VP.n8 50.7491
R65 VP.n88 VP.n87 50.7491
R66 VP.n43 VP.n42 50.7491
R67 VP.n31 VP.n22 50.7491
R68 VP.n76 VP.n75 30.405
R69 VP.n89 VP.n88 30.405
R70 VP.n44 VP.n43 30.405
R71 VP.n31 VP.n30 30.405
R72 VP.n63 VP.n62 24.5923
R73 VP.n63 VP.n12 24.5923
R74 VP.n68 VP.n67 24.5923
R75 VP.n70 VP.n68 24.5923
R76 VP.n74 VP.n10 24.5923
R77 VP.n75 VP.n74 24.5923
R78 VP.n80 VP.n8 24.5923
R79 VP.n81 VP.n80 24.5923
R80 VP.n83 VP.n6 24.5923
R81 VP.n87 VP.n6 24.5923
R82 VP.n89 VP.n4 24.5923
R83 VP.n93 VP.n4 24.5923
R84 VP.n96 VP.n95 24.5923
R85 VP.n96 VP.n2 24.5923
R86 VP.n101 VP.n100 24.5923
R87 VP.n102 VP.n101 24.5923
R88 VP.n56 VP.n55 24.5923
R89 VP.n57 VP.n56 24.5923
R90 VP.n44 VP.n18 24.5923
R91 VP.n48 VP.n18 24.5923
R92 VP.n51 VP.n50 24.5923
R93 VP.n51 VP.n16 24.5923
R94 VP.n35 VP.n22 24.5923
R95 VP.n36 VP.n35 24.5923
R96 VP.n38 VP.n20 24.5923
R97 VP.n42 VP.n20 24.5923
R98 VP.n29 VP.n24 24.5923
R99 VP.n30 VP.n29 24.5923
R100 VP.n70 VP.n69 22.625
R101 VP.n95 VP.n94 22.625
R102 VP.n50 VP.n49 22.625
R103 VP.n62 VP.n61 16.2311
R104 VP.n102 VP.n0 16.2311
R105 VP.n57 VP.n14 16.2311
R106 VP.n82 VP.n81 12.2964
R107 VP.n83 VP.n82 12.2964
R108 VP.n37 VP.n36 12.2964
R109 VP.n38 VP.n37 12.2964
R110 VP.n27 VP.n26 5.81313
R111 VP.n69 VP.n10 1.96785
R112 VP.n94 VP.n93 1.96785
R113 VP.n49 VP.n48 1.96785
R114 VP.n25 VP.n24 1.96785
R115 VP.n59 VP.n58 0.354861
R116 VP.n60 VP.n13 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n28 VP.n27 0.189894
R120 VP.n28 VP.n23 0.189894
R121 VP.n32 VP.n23 0.189894
R122 VP.n33 VP.n32 0.189894
R123 VP.n34 VP.n33 0.189894
R124 VP.n34 VP.n21 0.189894
R125 VP.n39 VP.n21 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n19 0.189894
R129 VP.n45 VP.n19 0.189894
R130 VP.n46 VP.n45 0.189894
R131 VP.n47 VP.n46 0.189894
R132 VP.n47 VP.n17 0.189894
R133 VP.n52 VP.n17 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n15 0.189894
R137 VP.n58 VP.n15 0.189894
R138 VP.n64 VP.n13 0.189894
R139 VP.n65 VP.n64 0.189894
R140 VP.n66 VP.n65 0.189894
R141 VP.n66 VP.n11 0.189894
R142 VP.n71 VP.n11 0.189894
R143 VP.n72 VP.n71 0.189894
R144 VP.n73 VP.n72 0.189894
R145 VP.n73 VP.n9 0.189894
R146 VP.n77 VP.n9 0.189894
R147 VP.n78 VP.n77 0.189894
R148 VP.n79 VP.n78 0.189894
R149 VP.n79 VP.n7 0.189894
R150 VP.n84 VP.n7 0.189894
R151 VP.n85 VP.n84 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n86 VP.n5 0.189894
R154 VP.n90 VP.n5 0.189894
R155 VP.n91 VP.n90 0.189894
R156 VP.n92 VP.n91 0.189894
R157 VP.n92 VP.n3 0.189894
R158 VP.n97 VP.n3 0.189894
R159 VP.n98 VP.n97 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n99 VP.n1 0.189894
R162 VP.n103 VP.n1 0.189894
R163 VTAIL.n11 VTAIL.t9 48.5487
R164 VTAIL.n17 VTAIL.t7 48.5485
R165 VTAIL.n2 VTAIL.t16 48.5485
R166 VTAIL.n16 VTAIL.t12 48.5485
R167 VTAIL.n15 VTAIL.n14 47.1035
R168 VTAIL.n13 VTAIL.n12 47.1035
R169 VTAIL.n10 VTAIL.n9 47.1035
R170 VTAIL.n8 VTAIL.n7 47.1035
R171 VTAIL.n19 VTAIL.n18 47.1033
R172 VTAIL.n1 VTAIL.n0 47.1033
R173 VTAIL.n4 VTAIL.n3 47.1033
R174 VTAIL.n6 VTAIL.n5 47.1033
R175 VTAIL.n8 VTAIL.n6 29.8496
R176 VTAIL.n17 VTAIL.n16 27.0134
R177 VTAIL.n10 VTAIL.n8 2.83671
R178 VTAIL.n11 VTAIL.n10 2.83671
R179 VTAIL.n15 VTAIL.n13 2.83671
R180 VTAIL.n16 VTAIL.n15 2.83671
R181 VTAIL.n6 VTAIL.n4 2.83671
R182 VTAIL.n4 VTAIL.n2 2.83671
R183 VTAIL.n19 VTAIL.n17 2.83671
R184 VTAIL VTAIL.n1 2.18584
R185 VTAIL.n13 VTAIL.n11 1.88843
R186 VTAIL.n2 VTAIL.n1 1.88843
R187 VTAIL.n18 VTAIL.t4 1.44576
R188 VTAIL.n18 VTAIL.t5 1.44576
R189 VTAIL.n0 VTAIL.t3 1.44576
R190 VTAIL.n0 VTAIL.t1 1.44576
R191 VTAIL.n3 VTAIL.t19 1.44576
R192 VTAIL.n3 VTAIL.t17 1.44576
R193 VTAIL.n5 VTAIL.t11 1.44576
R194 VTAIL.n5 VTAIL.t15 1.44576
R195 VTAIL.n14 VTAIL.t10 1.44576
R196 VTAIL.n14 VTAIL.t13 1.44576
R197 VTAIL.n12 VTAIL.t18 1.44576
R198 VTAIL.n12 VTAIL.t14 1.44576
R199 VTAIL.n9 VTAIL.t8 1.44576
R200 VTAIL.n9 VTAIL.t6 1.44576
R201 VTAIL.n7 VTAIL.t0 1.44576
R202 VTAIL.n7 VTAIL.t2 1.44576
R203 VTAIL VTAIL.n19 0.651362
R204 VDD1.n1 VDD1.t8 68.0637
R205 VDD1.n3 VDD1.t4 68.0635
R206 VDD1.n5 VDD1.n4 65.8539
R207 VDD1.n1 VDD1.n0 63.7823
R208 VDD1.n7 VDD1.n6 63.7821
R209 VDD1.n3 VDD1.n2 63.7821
R210 VDD1.n7 VDD1.n5 50.9987
R211 VDD1 VDD1.n7 2.06947
R212 VDD1.n6 VDD1.t6 1.44576
R213 VDD1.n6 VDD1.t3 1.44576
R214 VDD1.n0 VDD1.t2 1.44576
R215 VDD1.n0 VDD1.t1 1.44576
R216 VDD1.n4 VDD1.t7 1.44576
R217 VDD1.n4 VDD1.t5 1.44576
R218 VDD1.n2 VDD1.t0 1.44576
R219 VDD1.n2 VDD1.t9 1.44576
R220 VDD1 VDD1.n1 0.767741
R221 VDD1.n5 VDD1.n3 0.654206
R222 B.n852 B.n851 585
R223 B.n852 B.n120 585
R224 B.n855 B.n854 585
R225 B.n856 B.n176 585
R226 B.n858 B.n857 585
R227 B.n860 B.n175 585
R228 B.n863 B.n862 585
R229 B.n864 B.n174 585
R230 B.n866 B.n865 585
R231 B.n868 B.n173 585
R232 B.n871 B.n870 585
R233 B.n872 B.n172 585
R234 B.n874 B.n873 585
R235 B.n876 B.n171 585
R236 B.n879 B.n878 585
R237 B.n880 B.n170 585
R238 B.n882 B.n881 585
R239 B.n884 B.n169 585
R240 B.n887 B.n886 585
R241 B.n888 B.n168 585
R242 B.n890 B.n889 585
R243 B.n892 B.n167 585
R244 B.n895 B.n894 585
R245 B.n896 B.n166 585
R246 B.n898 B.n897 585
R247 B.n900 B.n165 585
R248 B.n903 B.n902 585
R249 B.n904 B.n164 585
R250 B.n906 B.n905 585
R251 B.n908 B.n163 585
R252 B.n911 B.n910 585
R253 B.n912 B.n162 585
R254 B.n914 B.n913 585
R255 B.n916 B.n161 585
R256 B.n919 B.n918 585
R257 B.n920 B.n160 585
R258 B.n922 B.n921 585
R259 B.n924 B.n159 585
R260 B.n927 B.n926 585
R261 B.n928 B.n158 585
R262 B.n930 B.n929 585
R263 B.n932 B.n157 585
R264 B.n935 B.n934 585
R265 B.n936 B.n156 585
R266 B.n938 B.n937 585
R267 B.n940 B.n155 585
R268 B.n943 B.n942 585
R269 B.n944 B.n152 585
R270 B.n947 B.n946 585
R271 B.n949 B.n151 585
R272 B.n952 B.n951 585
R273 B.n953 B.n150 585
R274 B.n955 B.n954 585
R275 B.n957 B.n149 585
R276 B.n960 B.n959 585
R277 B.n961 B.n145 585
R278 B.n963 B.n962 585
R279 B.n965 B.n144 585
R280 B.n968 B.n967 585
R281 B.n969 B.n143 585
R282 B.n971 B.n970 585
R283 B.n973 B.n142 585
R284 B.n976 B.n975 585
R285 B.n977 B.n141 585
R286 B.n979 B.n978 585
R287 B.n981 B.n140 585
R288 B.n984 B.n983 585
R289 B.n985 B.n139 585
R290 B.n987 B.n986 585
R291 B.n989 B.n138 585
R292 B.n992 B.n991 585
R293 B.n993 B.n137 585
R294 B.n995 B.n994 585
R295 B.n997 B.n136 585
R296 B.n1000 B.n999 585
R297 B.n1001 B.n135 585
R298 B.n1003 B.n1002 585
R299 B.n1005 B.n134 585
R300 B.n1008 B.n1007 585
R301 B.n1009 B.n133 585
R302 B.n1011 B.n1010 585
R303 B.n1013 B.n132 585
R304 B.n1016 B.n1015 585
R305 B.n1017 B.n131 585
R306 B.n1019 B.n1018 585
R307 B.n1021 B.n130 585
R308 B.n1024 B.n1023 585
R309 B.n1025 B.n129 585
R310 B.n1027 B.n1026 585
R311 B.n1029 B.n128 585
R312 B.n1032 B.n1031 585
R313 B.n1033 B.n127 585
R314 B.n1035 B.n1034 585
R315 B.n1037 B.n126 585
R316 B.n1040 B.n1039 585
R317 B.n1041 B.n125 585
R318 B.n1043 B.n1042 585
R319 B.n1045 B.n124 585
R320 B.n1048 B.n1047 585
R321 B.n1049 B.n123 585
R322 B.n1051 B.n1050 585
R323 B.n1053 B.n122 585
R324 B.n1056 B.n1055 585
R325 B.n1057 B.n121 585
R326 B.n850 B.n119 585
R327 B.n1060 B.n119 585
R328 B.n849 B.n118 585
R329 B.n1061 B.n118 585
R330 B.n848 B.n117 585
R331 B.n1062 B.n117 585
R332 B.n847 B.n846 585
R333 B.n846 B.n113 585
R334 B.n845 B.n112 585
R335 B.n1068 B.n112 585
R336 B.n844 B.n111 585
R337 B.n1069 B.n111 585
R338 B.n843 B.n110 585
R339 B.n1070 B.n110 585
R340 B.n842 B.n841 585
R341 B.n841 B.n109 585
R342 B.n840 B.n105 585
R343 B.n1076 B.n105 585
R344 B.n839 B.n104 585
R345 B.n1077 B.n104 585
R346 B.n838 B.n103 585
R347 B.n1078 B.n103 585
R348 B.n837 B.n836 585
R349 B.n836 B.n99 585
R350 B.n835 B.n98 585
R351 B.n1084 B.n98 585
R352 B.n834 B.n97 585
R353 B.n1085 B.n97 585
R354 B.n833 B.n96 585
R355 B.n1086 B.n96 585
R356 B.n832 B.n831 585
R357 B.n831 B.n92 585
R358 B.n830 B.n91 585
R359 B.n1092 B.n91 585
R360 B.n829 B.n90 585
R361 B.n1093 B.n90 585
R362 B.n828 B.n89 585
R363 B.n1094 B.n89 585
R364 B.n827 B.n826 585
R365 B.n826 B.n85 585
R366 B.n825 B.n84 585
R367 B.n1100 B.n84 585
R368 B.n824 B.n83 585
R369 B.n1101 B.n83 585
R370 B.n823 B.n82 585
R371 B.n1102 B.n82 585
R372 B.n822 B.n821 585
R373 B.n821 B.n78 585
R374 B.n820 B.n77 585
R375 B.n1108 B.n77 585
R376 B.n819 B.n76 585
R377 B.n1109 B.n76 585
R378 B.n818 B.n75 585
R379 B.n1110 B.n75 585
R380 B.n817 B.n816 585
R381 B.n816 B.n71 585
R382 B.n815 B.n70 585
R383 B.n1116 B.n70 585
R384 B.n814 B.n69 585
R385 B.n1117 B.n69 585
R386 B.n813 B.n68 585
R387 B.n1118 B.n68 585
R388 B.n812 B.n811 585
R389 B.n811 B.n64 585
R390 B.n810 B.n63 585
R391 B.n1124 B.n63 585
R392 B.n809 B.n62 585
R393 B.n1125 B.n62 585
R394 B.n808 B.n61 585
R395 B.n1126 B.n61 585
R396 B.n807 B.n806 585
R397 B.n806 B.n57 585
R398 B.n805 B.n56 585
R399 B.n1132 B.n56 585
R400 B.n804 B.n55 585
R401 B.n1133 B.n55 585
R402 B.n803 B.n54 585
R403 B.n1134 B.n54 585
R404 B.n802 B.n801 585
R405 B.n801 B.n50 585
R406 B.n800 B.n49 585
R407 B.n1140 B.n49 585
R408 B.n799 B.n48 585
R409 B.n1141 B.n48 585
R410 B.n798 B.n47 585
R411 B.n1142 B.n47 585
R412 B.n797 B.n796 585
R413 B.n796 B.n43 585
R414 B.n795 B.n42 585
R415 B.n1148 B.n42 585
R416 B.n794 B.n41 585
R417 B.n1149 B.n41 585
R418 B.n793 B.n40 585
R419 B.n1150 B.n40 585
R420 B.n792 B.n791 585
R421 B.n791 B.n36 585
R422 B.n790 B.n35 585
R423 B.n1156 B.n35 585
R424 B.n789 B.n34 585
R425 B.n1157 B.n34 585
R426 B.n788 B.n33 585
R427 B.n1158 B.n33 585
R428 B.n787 B.n786 585
R429 B.n786 B.n29 585
R430 B.n785 B.n28 585
R431 B.n1164 B.n28 585
R432 B.n784 B.n27 585
R433 B.n1165 B.n27 585
R434 B.n783 B.n26 585
R435 B.n1166 B.n26 585
R436 B.n782 B.n781 585
R437 B.n781 B.n22 585
R438 B.n780 B.n21 585
R439 B.n1172 B.n21 585
R440 B.n779 B.n20 585
R441 B.n1173 B.n20 585
R442 B.n778 B.n19 585
R443 B.n1174 B.n19 585
R444 B.n777 B.n776 585
R445 B.n776 B.n18 585
R446 B.n775 B.n14 585
R447 B.n1180 B.n14 585
R448 B.n774 B.n13 585
R449 B.n1181 B.n13 585
R450 B.n773 B.n12 585
R451 B.n1182 B.n12 585
R452 B.n772 B.n771 585
R453 B.n771 B.n8 585
R454 B.n770 B.n7 585
R455 B.n1188 B.n7 585
R456 B.n769 B.n6 585
R457 B.n1189 B.n6 585
R458 B.n768 B.n5 585
R459 B.n1190 B.n5 585
R460 B.n767 B.n766 585
R461 B.n766 B.n4 585
R462 B.n765 B.n177 585
R463 B.n765 B.n764 585
R464 B.n755 B.n178 585
R465 B.n179 B.n178 585
R466 B.n757 B.n756 585
R467 B.n758 B.n757 585
R468 B.n754 B.n184 585
R469 B.n184 B.n183 585
R470 B.n753 B.n752 585
R471 B.n752 B.n751 585
R472 B.n186 B.n185 585
R473 B.n744 B.n186 585
R474 B.n743 B.n742 585
R475 B.n745 B.n743 585
R476 B.n741 B.n191 585
R477 B.n191 B.n190 585
R478 B.n740 B.n739 585
R479 B.n739 B.n738 585
R480 B.n193 B.n192 585
R481 B.n194 B.n193 585
R482 B.n731 B.n730 585
R483 B.n732 B.n731 585
R484 B.n729 B.n199 585
R485 B.n199 B.n198 585
R486 B.n728 B.n727 585
R487 B.n727 B.n726 585
R488 B.n201 B.n200 585
R489 B.n202 B.n201 585
R490 B.n719 B.n718 585
R491 B.n720 B.n719 585
R492 B.n717 B.n206 585
R493 B.n210 B.n206 585
R494 B.n716 B.n715 585
R495 B.n715 B.n714 585
R496 B.n208 B.n207 585
R497 B.n209 B.n208 585
R498 B.n707 B.n706 585
R499 B.n708 B.n707 585
R500 B.n705 B.n215 585
R501 B.n215 B.n214 585
R502 B.n704 B.n703 585
R503 B.n703 B.n702 585
R504 B.n217 B.n216 585
R505 B.n218 B.n217 585
R506 B.n695 B.n694 585
R507 B.n696 B.n695 585
R508 B.n693 B.n223 585
R509 B.n223 B.n222 585
R510 B.n692 B.n691 585
R511 B.n691 B.n690 585
R512 B.n225 B.n224 585
R513 B.n226 B.n225 585
R514 B.n683 B.n682 585
R515 B.n684 B.n683 585
R516 B.n681 B.n231 585
R517 B.n231 B.n230 585
R518 B.n680 B.n679 585
R519 B.n679 B.n678 585
R520 B.n233 B.n232 585
R521 B.n234 B.n233 585
R522 B.n671 B.n670 585
R523 B.n672 B.n671 585
R524 B.n669 B.n239 585
R525 B.n239 B.n238 585
R526 B.n668 B.n667 585
R527 B.n667 B.n666 585
R528 B.n241 B.n240 585
R529 B.n242 B.n241 585
R530 B.n659 B.n658 585
R531 B.n660 B.n659 585
R532 B.n657 B.n247 585
R533 B.n247 B.n246 585
R534 B.n656 B.n655 585
R535 B.n655 B.n654 585
R536 B.n249 B.n248 585
R537 B.n250 B.n249 585
R538 B.n647 B.n646 585
R539 B.n648 B.n647 585
R540 B.n645 B.n255 585
R541 B.n255 B.n254 585
R542 B.n644 B.n643 585
R543 B.n643 B.n642 585
R544 B.n257 B.n256 585
R545 B.n258 B.n257 585
R546 B.n635 B.n634 585
R547 B.n636 B.n635 585
R548 B.n633 B.n263 585
R549 B.n263 B.n262 585
R550 B.n632 B.n631 585
R551 B.n631 B.n630 585
R552 B.n265 B.n264 585
R553 B.n266 B.n265 585
R554 B.n623 B.n622 585
R555 B.n624 B.n623 585
R556 B.n621 B.n271 585
R557 B.n271 B.n270 585
R558 B.n620 B.n619 585
R559 B.n619 B.n618 585
R560 B.n273 B.n272 585
R561 B.n274 B.n273 585
R562 B.n611 B.n610 585
R563 B.n612 B.n611 585
R564 B.n609 B.n279 585
R565 B.n279 B.n278 585
R566 B.n608 B.n607 585
R567 B.n607 B.n606 585
R568 B.n281 B.n280 585
R569 B.n282 B.n281 585
R570 B.n599 B.n598 585
R571 B.n600 B.n599 585
R572 B.n597 B.n287 585
R573 B.n287 B.n286 585
R574 B.n596 B.n595 585
R575 B.n595 B.n594 585
R576 B.n289 B.n288 585
R577 B.n587 B.n289 585
R578 B.n586 B.n585 585
R579 B.n588 B.n586 585
R580 B.n584 B.n294 585
R581 B.n294 B.n293 585
R582 B.n583 B.n582 585
R583 B.n582 B.n581 585
R584 B.n296 B.n295 585
R585 B.n297 B.n296 585
R586 B.n574 B.n573 585
R587 B.n575 B.n574 585
R588 B.n572 B.n302 585
R589 B.n302 B.n301 585
R590 B.n571 B.n570 585
R591 B.n570 B.n569 585
R592 B.n566 B.n306 585
R593 B.n565 B.n564 585
R594 B.n562 B.n307 585
R595 B.n562 B.n305 585
R596 B.n561 B.n560 585
R597 B.n559 B.n558 585
R598 B.n557 B.n309 585
R599 B.n555 B.n554 585
R600 B.n553 B.n310 585
R601 B.n552 B.n551 585
R602 B.n549 B.n311 585
R603 B.n547 B.n546 585
R604 B.n545 B.n312 585
R605 B.n544 B.n543 585
R606 B.n541 B.n313 585
R607 B.n539 B.n538 585
R608 B.n537 B.n314 585
R609 B.n536 B.n535 585
R610 B.n533 B.n315 585
R611 B.n531 B.n530 585
R612 B.n529 B.n316 585
R613 B.n528 B.n527 585
R614 B.n525 B.n317 585
R615 B.n523 B.n522 585
R616 B.n521 B.n318 585
R617 B.n520 B.n519 585
R618 B.n517 B.n319 585
R619 B.n515 B.n514 585
R620 B.n513 B.n320 585
R621 B.n512 B.n511 585
R622 B.n509 B.n321 585
R623 B.n507 B.n506 585
R624 B.n505 B.n322 585
R625 B.n504 B.n503 585
R626 B.n501 B.n323 585
R627 B.n499 B.n498 585
R628 B.n497 B.n324 585
R629 B.n496 B.n495 585
R630 B.n493 B.n325 585
R631 B.n491 B.n490 585
R632 B.n489 B.n326 585
R633 B.n488 B.n487 585
R634 B.n485 B.n327 585
R635 B.n483 B.n482 585
R636 B.n481 B.n328 585
R637 B.n480 B.n479 585
R638 B.n477 B.n329 585
R639 B.n475 B.n474 585
R640 B.n472 B.n330 585
R641 B.n471 B.n470 585
R642 B.n468 B.n333 585
R643 B.n466 B.n465 585
R644 B.n464 B.n334 585
R645 B.n463 B.n462 585
R646 B.n460 B.n335 585
R647 B.n458 B.n457 585
R648 B.n456 B.n336 585
R649 B.n454 B.n453 585
R650 B.n451 B.n339 585
R651 B.n449 B.n448 585
R652 B.n447 B.n340 585
R653 B.n446 B.n445 585
R654 B.n443 B.n341 585
R655 B.n441 B.n440 585
R656 B.n439 B.n342 585
R657 B.n438 B.n437 585
R658 B.n435 B.n343 585
R659 B.n433 B.n432 585
R660 B.n431 B.n344 585
R661 B.n430 B.n429 585
R662 B.n427 B.n345 585
R663 B.n425 B.n424 585
R664 B.n423 B.n346 585
R665 B.n422 B.n421 585
R666 B.n419 B.n347 585
R667 B.n417 B.n416 585
R668 B.n415 B.n348 585
R669 B.n414 B.n413 585
R670 B.n411 B.n349 585
R671 B.n409 B.n408 585
R672 B.n407 B.n350 585
R673 B.n406 B.n405 585
R674 B.n403 B.n351 585
R675 B.n401 B.n400 585
R676 B.n399 B.n352 585
R677 B.n398 B.n397 585
R678 B.n395 B.n353 585
R679 B.n393 B.n392 585
R680 B.n391 B.n354 585
R681 B.n390 B.n389 585
R682 B.n387 B.n355 585
R683 B.n385 B.n384 585
R684 B.n383 B.n356 585
R685 B.n382 B.n381 585
R686 B.n379 B.n357 585
R687 B.n377 B.n376 585
R688 B.n375 B.n358 585
R689 B.n374 B.n373 585
R690 B.n371 B.n359 585
R691 B.n369 B.n368 585
R692 B.n367 B.n360 585
R693 B.n366 B.n365 585
R694 B.n363 B.n361 585
R695 B.n304 B.n303 585
R696 B.n568 B.n567 585
R697 B.n569 B.n568 585
R698 B.n300 B.n299 585
R699 B.n301 B.n300 585
R700 B.n577 B.n576 585
R701 B.n576 B.n575 585
R702 B.n578 B.n298 585
R703 B.n298 B.n297 585
R704 B.n580 B.n579 585
R705 B.n581 B.n580 585
R706 B.n292 B.n291 585
R707 B.n293 B.n292 585
R708 B.n590 B.n589 585
R709 B.n589 B.n588 585
R710 B.n591 B.n290 585
R711 B.n587 B.n290 585
R712 B.n593 B.n592 585
R713 B.n594 B.n593 585
R714 B.n285 B.n284 585
R715 B.n286 B.n285 585
R716 B.n602 B.n601 585
R717 B.n601 B.n600 585
R718 B.n603 B.n283 585
R719 B.n283 B.n282 585
R720 B.n605 B.n604 585
R721 B.n606 B.n605 585
R722 B.n277 B.n276 585
R723 B.n278 B.n277 585
R724 B.n614 B.n613 585
R725 B.n613 B.n612 585
R726 B.n615 B.n275 585
R727 B.n275 B.n274 585
R728 B.n617 B.n616 585
R729 B.n618 B.n617 585
R730 B.n269 B.n268 585
R731 B.n270 B.n269 585
R732 B.n626 B.n625 585
R733 B.n625 B.n624 585
R734 B.n627 B.n267 585
R735 B.n267 B.n266 585
R736 B.n629 B.n628 585
R737 B.n630 B.n629 585
R738 B.n261 B.n260 585
R739 B.n262 B.n261 585
R740 B.n638 B.n637 585
R741 B.n637 B.n636 585
R742 B.n639 B.n259 585
R743 B.n259 B.n258 585
R744 B.n641 B.n640 585
R745 B.n642 B.n641 585
R746 B.n253 B.n252 585
R747 B.n254 B.n253 585
R748 B.n650 B.n649 585
R749 B.n649 B.n648 585
R750 B.n651 B.n251 585
R751 B.n251 B.n250 585
R752 B.n653 B.n652 585
R753 B.n654 B.n653 585
R754 B.n245 B.n244 585
R755 B.n246 B.n245 585
R756 B.n662 B.n661 585
R757 B.n661 B.n660 585
R758 B.n663 B.n243 585
R759 B.n243 B.n242 585
R760 B.n665 B.n664 585
R761 B.n666 B.n665 585
R762 B.n237 B.n236 585
R763 B.n238 B.n237 585
R764 B.n674 B.n673 585
R765 B.n673 B.n672 585
R766 B.n675 B.n235 585
R767 B.n235 B.n234 585
R768 B.n677 B.n676 585
R769 B.n678 B.n677 585
R770 B.n229 B.n228 585
R771 B.n230 B.n229 585
R772 B.n686 B.n685 585
R773 B.n685 B.n684 585
R774 B.n687 B.n227 585
R775 B.n227 B.n226 585
R776 B.n689 B.n688 585
R777 B.n690 B.n689 585
R778 B.n221 B.n220 585
R779 B.n222 B.n221 585
R780 B.n698 B.n697 585
R781 B.n697 B.n696 585
R782 B.n699 B.n219 585
R783 B.n219 B.n218 585
R784 B.n701 B.n700 585
R785 B.n702 B.n701 585
R786 B.n213 B.n212 585
R787 B.n214 B.n213 585
R788 B.n710 B.n709 585
R789 B.n709 B.n708 585
R790 B.n711 B.n211 585
R791 B.n211 B.n209 585
R792 B.n713 B.n712 585
R793 B.n714 B.n713 585
R794 B.n205 B.n204 585
R795 B.n210 B.n205 585
R796 B.n722 B.n721 585
R797 B.n721 B.n720 585
R798 B.n723 B.n203 585
R799 B.n203 B.n202 585
R800 B.n725 B.n724 585
R801 B.n726 B.n725 585
R802 B.n197 B.n196 585
R803 B.n198 B.n197 585
R804 B.n734 B.n733 585
R805 B.n733 B.n732 585
R806 B.n735 B.n195 585
R807 B.n195 B.n194 585
R808 B.n737 B.n736 585
R809 B.n738 B.n737 585
R810 B.n189 B.n188 585
R811 B.n190 B.n189 585
R812 B.n747 B.n746 585
R813 B.n746 B.n745 585
R814 B.n748 B.n187 585
R815 B.n744 B.n187 585
R816 B.n750 B.n749 585
R817 B.n751 B.n750 585
R818 B.n182 B.n181 585
R819 B.n183 B.n182 585
R820 B.n760 B.n759 585
R821 B.n759 B.n758 585
R822 B.n761 B.n180 585
R823 B.n180 B.n179 585
R824 B.n763 B.n762 585
R825 B.n764 B.n763 585
R826 B.n2 B.n0 585
R827 B.n4 B.n2 585
R828 B.n3 B.n1 585
R829 B.n1189 B.n3 585
R830 B.n1187 B.n1186 585
R831 B.n1188 B.n1187 585
R832 B.n1185 B.n9 585
R833 B.n9 B.n8 585
R834 B.n1184 B.n1183 585
R835 B.n1183 B.n1182 585
R836 B.n11 B.n10 585
R837 B.n1181 B.n11 585
R838 B.n1179 B.n1178 585
R839 B.n1180 B.n1179 585
R840 B.n1177 B.n15 585
R841 B.n18 B.n15 585
R842 B.n1176 B.n1175 585
R843 B.n1175 B.n1174 585
R844 B.n17 B.n16 585
R845 B.n1173 B.n17 585
R846 B.n1171 B.n1170 585
R847 B.n1172 B.n1171 585
R848 B.n1169 B.n23 585
R849 B.n23 B.n22 585
R850 B.n1168 B.n1167 585
R851 B.n1167 B.n1166 585
R852 B.n25 B.n24 585
R853 B.n1165 B.n25 585
R854 B.n1163 B.n1162 585
R855 B.n1164 B.n1163 585
R856 B.n1161 B.n30 585
R857 B.n30 B.n29 585
R858 B.n1160 B.n1159 585
R859 B.n1159 B.n1158 585
R860 B.n32 B.n31 585
R861 B.n1157 B.n32 585
R862 B.n1155 B.n1154 585
R863 B.n1156 B.n1155 585
R864 B.n1153 B.n37 585
R865 B.n37 B.n36 585
R866 B.n1152 B.n1151 585
R867 B.n1151 B.n1150 585
R868 B.n39 B.n38 585
R869 B.n1149 B.n39 585
R870 B.n1147 B.n1146 585
R871 B.n1148 B.n1147 585
R872 B.n1145 B.n44 585
R873 B.n44 B.n43 585
R874 B.n1144 B.n1143 585
R875 B.n1143 B.n1142 585
R876 B.n46 B.n45 585
R877 B.n1141 B.n46 585
R878 B.n1139 B.n1138 585
R879 B.n1140 B.n1139 585
R880 B.n1137 B.n51 585
R881 B.n51 B.n50 585
R882 B.n1136 B.n1135 585
R883 B.n1135 B.n1134 585
R884 B.n53 B.n52 585
R885 B.n1133 B.n53 585
R886 B.n1131 B.n1130 585
R887 B.n1132 B.n1131 585
R888 B.n1129 B.n58 585
R889 B.n58 B.n57 585
R890 B.n1128 B.n1127 585
R891 B.n1127 B.n1126 585
R892 B.n60 B.n59 585
R893 B.n1125 B.n60 585
R894 B.n1123 B.n1122 585
R895 B.n1124 B.n1123 585
R896 B.n1121 B.n65 585
R897 B.n65 B.n64 585
R898 B.n1120 B.n1119 585
R899 B.n1119 B.n1118 585
R900 B.n67 B.n66 585
R901 B.n1117 B.n67 585
R902 B.n1115 B.n1114 585
R903 B.n1116 B.n1115 585
R904 B.n1113 B.n72 585
R905 B.n72 B.n71 585
R906 B.n1112 B.n1111 585
R907 B.n1111 B.n1110 585
R908 B.n74 B.n73 585
R909 B.n1109 B.n74 585
R910 B.n1107 B.n1106 585
R911 B.n1108 B.n1107 585
R912 B.n1105 B.n79 585
R913 B.n79 B.n78 585
R914 B.n1104 B.n1103 585
R915 B.n1103 B.n1102 585
R916 B.n81 B.n80 585
R917 B.n1101 B.n81 585
R918 B.n1099 B.n1098 585
R919 B.n1100 B.n1099 585
R920 B.n1097 B.n86 585
R921 B.n86 B.n85 585
R922 B.n1096 B.n1095 585
R923 B.n1095 B.n1094 585
R924 B.n88 B.n87 585
R925 B.n1093 B.n88 585
R926 B.n1091 B.n1090 585
R927 B.n1092 B.n1091 585
R928 B.n1089 B.n93 585
R929 B.n93 B.n92 585
R930 B.n1088 B.n1087 585
R931 B.n1087 B.n1086 585
R932 B.n95 B.n94 585
R933 B.n1085 B.n95 585
R934 B.n1083 B.n1082 585
R935 B.n1084 B.n1083 585
R936 B.n1081 B.n100 585
R937 B.n100 B.n99 585
R938 B.n1080 B.n1079 585
R939 B.n1079 B.n1078 585
R940 B.n102 B.n101 585
R941 B.n1077 B.n102 585
R942 B.n1075 B.n1074 585
R943 B.n1076 B.n1075 585
R944 B.n1073 B.n106 585
R945 B.n109 B.n106 585
R946 B.n1072 B.n1071 585
R947 B.n1071 B.n1070 585
R948 B.n108 B.n107 585
R949 B.n1069 B.n108 585
R950 B.n1067 B.n1066 585
R951 B.n1068 B.n1067 585
R952 B.n1065 B.n114 585
R953 B.n114 B.n113 585
R954 B.n1064 B.n1063 585
R955 B.n1063 B.n1062 585
R956 B.n116 B.n115 585
R957 B.n1061 B.n116 585
R958 B.n1059 B.n1058 585
R959 B.n1060 B.n1059 585
R960 B.n1192 B.n1191 585
R961 B.n1191 B.n1190 585
R962 B.n568 B.n306 511.721
R963 B.n1059 B.n121 511.721
R964 B.n570 B.n304 511.721
R965 B.n852 B.n119 511.721
R966 B.n337 B.t12 320.077
R967 B.n331 B.t16 320.077
R968 B.n146 B.t9 320.077
R969 B.n153 B.t5 320.077
R970 B.n853 B.n120 256.663
R971 B.n859 B.n120 256.663
R972 B.n861 B.n120 256.663
R973 B.n867 B.n120 256.663
R974 B.n869 B.n120 256.663
R975 B.n875 B.n120 256.663
R976 B.n877 B.n120 256.663
R977 B.n883 B.n120 256.663
R978 B.n885 B.n120 256.663
R979 B.n891 B.n120 256.663
R980 B.n893 B.n120 256.663
R981 B.n899 B.n120 256.663
R982 B.n901 B.n120 256.663
R983 B.n907 B.n120 256.663
R984 B.n909 B.n120 256.663
R985 B.n915 B.n120 256.663
R986 B.n917 B.n120 256.663
R987 B.n923 B.n120 256.663
R988 B.n925 B.n120 256.663
R989 B.n931 B.n120 256.663
R990 B.n933 B.n120 256.663
R991 B.n939 B.n120 256.663
R992 B.n941 B.n120 256.663
R993 B.n948 B.n120 256.663
R994 B.n950 B.n120 256.663
R995 B.n956 B.n120 256.663
R996 B.n958 B.n120 256.663
R997 B.n964 B.n120 256.663
R998 B.n966 B.n120 256.663
R999 B.n972 B.n120 256.663
R1000 B.n974 B.n120 256.663
R1001 B.n980 B.n120 256.663
R1002 B.n982 B.n120 256.663
R1003 B.n988 B.n120 256.663
R1004 B.n990 B.n120 256.663
R1005 B.n996 B.n120 256.663
R1006 B.n998 B.n120 256.663
R1007 B.n1004 B.n120 256.663
R1008 B.n1006 B.n120 256.663
R1009 B.n1012 B.n120 256.663
R1010 B.n1014 B.n120 256.663
R1011 B.n1020 B.n120 256.663
R1012 B.n1022 B.n120 256.663
R1013 B.n1028 B.n120 256.663
R1014 B.n1030 B.n120 256.663
R1015 B.n1036 B.n120 256.663
R1016 B.n1038 B.n120 256.663
R1017 B.n1044 B.n120 256.663
R1018 B.n1046 B.n120 256.663
R1019 B.n1052 B.n120 256.663
R1020 B.n1054 B.n120 256.663
R1021 B.n563 B.n305 256.663
R1022 B.n308 B.n305 256.663
R1023 B.n556 B.n305 256.663
R1024 B.n550 B.n305 256.663
R1025 B.n548 B.n305 256.663
R1026 B.n542 B.n305 256.663
R1027 B.n540 B.n305 256.663
R1028 B.n534 B.n305 256.663
R1029 B.n532 B.n305 256.663
R1030 B.n526 B.n305 256.663
R1031 B.n524 B.n305 256.663
R1032 B.n518 B.n305 256.663
R1033 B.n516 B.n305 256.663
R1034 B.n510 B.n305 256.663
R1035 B.n508 B.n305 256.663
R1036 B.n502 B.n305 256.663
R1037 B.n500 B.n305 256.663
R1038 B.n494 B.n305 256.663
R1039 B.n492 B.n305 256.663
R1040 B.n486 B.n305 256.663
R1041 B.n484 B.n305 256.663
R1042 B.n478 B.n305 256.663
R1043 B.n476 B.n305 256.663
R1044 B.n469 B.n305 256.663
R1045 B.n467 B.n305 256.663
R1046 B.n461 B.n305 256.663
R1047 B.n459 B.n305 256.663
R1048 B.n452 B.n305 256.663
R1049 B.n450 B.n305 256.663
R1050 B.n444 B.n305 256.663
R1051 B.n442 B.n305 256.663
R1052 B.n436 B.n305 256.663
R1053 B.n434 B.n305 256.663
R1054 B.n428 B.n305 256.663
R1055 B.n426 B.n305 256.663
R1056 B.n420 B.n305 256.663
R1057 B.n418 B.n305 256.663
R1058 B.n412 B.n305 256.663
R1059 B.n410 B.n305 256.663
R1060 B.n404 B.n305 256.663
R1061 B.n402 B.n305 256.663
R1062 B.n396 B.n305 256.663
R1063 B.n394 B.n305 256.663
R1064 B.n388 B.n305 256.663
R1065 B.n386 B.n305 256.663
R1066 B.n380 B.n305 256.663
R1067 B.n378 B.n305 256.663
R1068 B.n372 B.n305 256.663
R1069 B.n370 B.n305 256.663
R1070 B.n364 B.n305 256.663
R1071 B.n362 B.n305 256.663
R1072 B.n568 B.n300 163.367
R1073 B.n576 B.n300 163.367
R1074 B.n576 B.n298 163.367
R1075 B.n580 B.n298 163.367
R1076 B.n580 B.n292 163.367
R1077 B.n589 B.n292 163.367
R1078 B.n589 B.n290 163.367
R1079 B.n593 B.n290 163.367
R1080 B.n593 B.n285 163.367
R1081 B.n601 B.n285 163.367
R1082 B.n601 B.n283 163.367
R1083 B.n605 B.n283 163.367
R1084 B.n605 B.n277 163.367
R1085 B.n613 B.n277 163.367
R1086 B.n613 B.n275 163.367
R1087 B.n617 B.n275 163.367
R1088 B.n617 B.n269 163.367
R1089 B.n625 B.n269 163.367
R1090 B.n625 B.n267 163.367
R1091 B.n629 B.n267 163.367
R1092 B.n629 B.n261 163.367
R1093 B.n637 B.n261 163.367
R1094 B.n637 B.n259 163.367
R1095 B.n641 B.n259 163.367
R1096 B.n641 B.n253 163.367
R1097 B.n649 B.n253 163.367
R1098 B.n649 B.n251 163.367
R1099 B.n653 B.n251 163.367
R1100 B.n653 B.n245 163.367
R1101 B.n661 B.n245 163.367
R1102 B.n661 B.n243 163.367
R1103 B.n665 B.n243 163.367
R1104 B.n665 B.n237 163.367
R1105 B.n673 B.n237 163.367
R1106 B.n673 B.n235 163.367
R1107 B.n677 B.n235 163.367
R1108 B.n677 B.n229 163.367
R1109 B.n685 B.n229 163.367
R1110 B.n685 B.n227 163.367
R1111 B.n689 B.n227 163.367
R1112 B.n689 B.n221 163.367
R1113 B.n697 B.n221 163.367
R1114 B.n697 B.n219 163.367
R1115 B.n701 B.n219 163.367
R1116 B.n701 B.n213 163.367
R1117 B.n709 B.n213 163.367
R1118 B.n709 B.n211 163.367
R1119 B.n713 B.n211 163.367
R1120 B.n713 B.n205 163.367
R1121 B.n721 B.n205 163.367
R1122 B.n721 B.n203 163.367
R1123 B.n725 B.n203 163.367
R1124 B.n725 B.n197 163.367
R1125 B.n733 B.n197 163.367
R1126 B.n733 B.n195 163.367
R1127 B.n737 B.n195 163.367
R1128 B.n737 B.n189 163.367
R1129 B.n746 B.n189 163.367
R1130 B.n746 B.n187 163.367
R1131 B.n750 B.n187 163.367
R1132 B.n750 B.n182 163.367
R1133 B.n759 B.n182 163.367
R1134 B.n759 B.n180 163.367
R1135 B.n763 B.n180 163.367
R1136 B.n763 B.n2 163.367
R1137 B.n1191 B.n2 163.367
R1138 B.n1191 B.n3 163.367
R1139 B.n1187 B.n3 163.367
R1140 B.n1187 B.n9 163.367
R1141 B.n1183 B.n9 163.367
R1142 B.n1183 B.n11 163.367
R1143 B.n1179 B.n11 163.367
R1144 B.n1179 B.n15 163.367
R1145 B.n1175 B.n15 163.367
R1146 B.n1175 B.n17 163.367
R1147 B.n1171 B.n17 163.367
R1148 B.n1171 B.n23 163.367
R1149 B.n1167 B.n23 163.367
R1150 B.n1167 B.n25 163.367
R1151 B.n1163 B.n25 163.367
R1152 B.n1163 B.n30 163.367
R1153 B.n1159 B.n30 163.367
R1154 B.n1159 B.n32 163.367
R1155 B.n1155 B.n32 163.367
R1156 B.n1155 B.n37 163.367
R1157 B.n1151 B.n37 163.367
R1158 B.n1151 B.n39 163.367
R1159 B.n1147 B.n39 163.367
R1160 B.n1147 B.n44 163.367
R1161 B.n1143 B.n44 163.367
R1162 B.n1143 B.n46 163.367
R1163 B.n1139 B.n46 163.367
R1164 B.n1139 B.n51 163.367
R1165 B.n1135 B.n51 163.367
R1166 B.n1135 B.n53 163.367
R1167 B.n1131 B.n53 163.367
R1168 B.n1131 B.n58 163.367
R1169 B.n1127 B.n58 163.367
R1170 B.n1127 B.n60 163.367
R1171 B.n1123 B.n60 163.367
R1172 B.n1123 B.n65 163.367
R1173 B.n1119 B.n65 163.367
R1174 B.n1119 B.n67 163.367
R1175 B.n1115 B.n67 163.367
R1176 B.n1115 B.n72 163.367
R1177 B.n1111 B.n72 163.367
R1178 B.n1111 B.n74 163.367
R1179 B.n1107 B.n74 163.367
R1180 B.n1107 B.n79 163.367
R1181 B.n1103 B.n79 163.367
R1182 B.n1103 B.n81 163.367
R1183 B.n1099 B.n81 163.367
R1184 B.n1099 B.n86 163.367
R1185 B.n1095 B.n86 163.367
R1186 B.n1095 B.n88 163.367
R1187 B.n1091 B.n88 163.367
R1188 B.n1091 B.n93 163.367
R1189 B.n1087 B.n93 163.367
R1190 B.n1087 B.n95 163.367
R1191 B.n1083 B.n95 163.367
R1192 B.n1083 B.n100 163.367
R1193 B.n1079 B.n100 163.367
R1194 B.n1079 B.n102 163.367
R1195 B.n1075 B.n102 163.367
R1196 B.n1075 B.n106 163.367
R1197 B.n1071 B.n106 163.367
R1198 B.n1071 B.n108 163.367
R1199 B.n1067 B.n108 163.367
R1200 B.n1067 B.n114 163.367
R1201 B.n1063 B.n114 163.367
R1202 B.n1063 B.n116 163.367
R1203 B.n1059 B.n116 163.367
R1204 B.n564 B.n562 163.367
R1205 B.n562 B.n561 163.367
R1206 B.n558 B.n557 163.367
R1207 B.n555 B.n310 163.367
R1208 B.n551 B.n549 163.367
R1209 B.n547 B.n312 163.367
R1210 B.n543 B.n541 163.367
R1211 B.n539 B.n314 163.367
R1212 B.n535 B.n533 163.367
R1213 B.n531 B.n316 163.367
R1214 B.n527 B.n525 163.367
R1215 B.n523 B.n318 163.367
R1216 B.n519 B.n517 163.367
R1217 B.n515 B.n320 163.367
R1218 B.n511 B.n509 163.367
R1219 B.n507 B.n322 163.367
R1220 B.n503 B.n501 163.367
R1221 B.n499 B.n324 163.367
R1222 B.n495 B.n493 163.367
R1223 B.n491 B.n326 163.367
R1224 B.n487 B.n485 163.367
R1225 B.n483 B.n328 163.367
R1226 B.n479 B.n477 163.367
R1227 B.n475 B.n330 163.367
R1228 B.n470 B.n468 163.367
R1229 B.n466 B.n334 163.367
R1230 B.n462 B.n460 163.367
R1231 B.n458 B.n336 163.367
R1232 B.n453 B.n451 163.367
R1233 B.n449 B.n340 163.367
R1234 B.n445 B.n443 163.367
R1235 B.n441 B.n342 163.367
R1236 B.n437 B.n435 163.367
R1237 B.n433 B.n344 163.367
R1238 B.n429 B.n427 163.367
R1239 B.n425 B.n346 163.367
R1240 B.n421 B.n419 163.367
R1241 B.n417 B.n348 163.367
R1242 B.n413 B.n411 163.367
R1243 B.n409 B.n350 163.367
R1244 B.n405 B.n403 163.367
R1245 B.n401 B.n352 163.367
R1246 B.n397 B.n395 163.367
R1247 B.n393 B.n354 163.367
R1248 B.n389 B.n387 163.367
R1249 B.n385 B.n356 163.367
R1250 B.n381 B.n379 163.367
R1251 B.n377 B.n358 163.367
R1252 B.n373 B.n371 163.367
R1253 B.n369 B.n360 163.367
R1254 B.n365 B.n363 163.367
R1255 B.n570 B.n302 163.367
R1256 B.n574 B.n302 163.367
R1257 B.n574 B.n296 163.367
R1258 B.n582 B.n296 163.367
R1259 B.n582 B.n294 163.367
R1260 B.n586 B.n294 163.367
R1261 B.n586 B.n289 163.367
R1262 B.n595 B.n289 163.367
R1263 B.n595 B.n287 163.367
R1264 B.n599 B.n287 163.367
R1265 B.n599 B.n281 163.367
R1266 B.n607 B.n281 163.367
R1267 B.n607 B.n279 163.367
R1268 B.n611 B.n279 163.367
R1269 B.n611 B.n273 163.367
R1270 B.n619 B.n273 163.367
R1271 B.n619 B.n271 163.367
R1272 B.n623 B.n271 163.367
R1273 B.n623 B.n265 163.367
R1274 B.n631 B.n265 163.367
R1275 B.n631 B.n263 163.367
R1276 B.n635 B.n263 163.367
R1277 B.n635 B.n257 163.367
R1278 B.n643 B.n257 163.367
R1279 B.n643 B.n255 163.367
R1280 B.n647 B.n255 163.367
R1281 B.n647 B.n249 163.367
R1282 B.n655 B.n249 163.367
R1283 B.n655 B.n247 163.367
R1284 B.n659 B.n247 163.367
R1285 B.n659 B.n241 163.367
R1286 B.n667 B.n241 163.367
R1287 B.n667 B.n239 163.367
R1288 B.n671 B.n239 163.367
R1289 B.n671 B.n233 163.367
R1290 B.n679 B.n233 163.367
R1291 B.n679 B.n231 163.367
R1292 B.n683 B.n231 163.367
R1293 B.n683 B.n225 163.367
R1294 B.n691 B.n225 163.367
R1295 B.n691 B.n223 163.367
R1296 B.n695 B.n223 163.367
R1297 B.n695 B.n217 163.367
R1298 B.n703 B.n217 163.367
R1299 B.n703 B.n215 163.367
R1300 B.n707 B.n215 163.367
R1301 B.n707 B.n208 163.367
R1302 B.n715 B.n208 163.367
R1303 B.n715 B.n206 163.367
R1304 B.n719 B.n206 163.367
R1305 B.n719 B.n201 163.367
R1306 B.n727 B.n201 163.367
R1307 B.n727 B.n199 163.367
R1308 B.n731 B.n199 163.367
R1309 B.n731 B.n193 163.367
R1310 B.n739 B.n193 163.367
R1311 B.n739 B.n191 163.367
R1312 B.n743 B.n191 163.367
R1313 B.n743 B.n186 163.367
R1314 B.n752 B.n186 163.367
R1315 B.n752 B.n184 163.367
R1316 B.n757 B.n184 163.367
R1317 B.n757 B.n178 163.367
R1318 B.n765 B.n178 163.367
R1319 B.n766 B.n765 163.367
R1320 B.n766 B.n5 163.367
R1321 B.n6 B.n5 163.367
R1322 B.n7 B.n6 163.367
R1323 B.n771 B.n7 163.367
R1324 B.n771 B.n12 163.367
R1325 B.n13 B.n12 163.367
R1326 B.n14 B.n13 163.367
R1327 B.n776 B.n14 163.367
R1328 B.n776 B.n19 163.367
R1329 B.n20 B.n19 163.367
R1330 B.n21 B.n20 163.367
R1331 B.n781 B.n21 163.367
R1332 B.n781 B.n26 163.367
R1333 B.n27 B.n26 163.367
R1334 B.n28 B.n27 163.367
R1335 B.n786 B.n28 163.367
R1336 B.n786 B.n33 163.367
R1337 B.n34 B.n33 163.367
R1338 B.n35 B.n34 163.367
R1339 B.n791 B.n35 163.367
R1340 B.n791 B.n40 163.367
R1341 B.n41 B.n40 163.367
R1342 B.n42 B.n41 163.367
R1343 B.n796 B.n42 163.367
R1344 B.n796 B.n47 163.367
R1345 B.n48 B.n47 163.367
R1346 B.n49 B.n48 163.367
R1347 B.n801 B.n49 163.367
R1348 B.n801 B.n54 163.367
R1349 B.n55 B.n54 163.367
R1350 B.n56 B.n55 163.367
R1351 B.n806 B.n56 163.367
R1352 B.n806 B.n61 163.367
R1353 B.n62 B.n61 163.367
R1354 B.n63 B.n62 163.367
R1355 B.n811 B.n63 163.367
R1356 B.n811 B.n68 163.367
R1357 B.n69 B.n68 163.367
R1358 B.n70 B.n69 163.367
R1359 B.n816 B.n70 163.367
R1360 B.n816 B.n75 163.367
R1361 B.n76 B.n75 163.367
R1362 B.n77 B.n76 163.367
R1363 B.n821 B.n77 163.367
R1364 B.n821 B.n82 163.367
R1365 B.n83 B.n82 163.367
R1366 B.n84 B.n83 163.367
R1367 B.n826 B.n84 163.367
R1368 B.n826 B.n89 163.367
R1369 B.n90 B.n89 163.367
R1370 B.n91 B.n90 163.367
R1371 B.n831 B.n91 163.367
R1372 B.n831 B.n96 163.367
R1373 B.n97 B.n96 163.367
R1374 B.n98 B.n97 163.367
R1375 B.n836 B.n98 163.367
R1376 B.n836 B.n103 163.367
R1377 B.n104 B.n103 163.367
R1378 B.n105 B.n104 163.367
R1379 B.n841 B.n105 163.367
R1380 B.n841 B.n110 163.367
R1381 B.n111 B.n110 163.367
R1382 B.n112 B.n111 163.367
R1383 B.n846 B.n112 163.367
R1384 B.n846 B.n117 163.367
R1385 B.n118 B.n117 163.367
R1386 B.n119 B.n118 163.367
R1387 B.n1055 B.n1053 163.367
R1388 B.n1051 B.n123 163.367
R1389 B.n1047 B.n1045 163.367
R1390 B.n1043 B.n125 163.367
R1391 B.n1039 B.n1037 163.367
R1392 B.n1035 B.n127 163.367
R1393 B.n1031 B.n1029 163.367
R1394 B.n1027 B.n129 163.367
R1395 B.n1023 B.n1021 163.367
R1396 B.n1019 B.n131 163.367
R1397 B.n1015 B.n1013 163.367
R1398 B.n1011 B.n133 163.367
R1399 B.n1007 B.n1005 163.367
R1400 B.n1003 B.n135 163.367
R1401 B.n999 B.n997 163.367
R1402 B.n995 B.n137 163.367
R1403 B.n991 B.n989 163.367
R1404 B.n987 B.n139 163.367
R1405 B.n983 B.n981 163.367
R1406 B.n979 B.n141 163.367
R1407 B.n975 B.n973 163.367
R1408 B.n971 B.n143 163.367
R1409 B.n967 B.n965 163.367
R1410 B.n963 B.n145 163.367
R1411 B.n959 B.n957 163.367
R1412 B.n955 B.n150 163.367
R1413 B.n951 B.n949 163.367
R1414 B.n947 B.n152 163.367
R1415 B.n942 B.n940 163.367
R1416 B.n938 B.n156 163.367
R1417 B.n934 B.n932 163.367
R1418 B.n930 B.n158 163.367
R1419 B.n926 B.n924 163.367
R1420 B.n922 B.n160 163.367
R1421 B.n918 B.n916 163.367
R1422 B.n914 B.n162 163.367
R1423 B.n910 B.n908 163.367
R1424 B.n906 B.n164 163.367
R1425 B.n902 B.n900 163.367
R1426 B.n898 B.n166 163.367
R1427 B.n894 B.n892 163.367
R1428 B.n890 B.n168 163.367
R1429 B.n886 B.n884 163.367
R1430 B.n882 B.n170 163.367
R1431 B.n878 B.n876 163.367
R1432 B.n874 B.n172 163.367
R1433 B.n870 B.n868 163.367
R1434 B.n866 B.n174 163.367
R1435 B.n862 B.n860 163.367
R1436 B.n858 B.n176 163.367
R1437 B.n854 B.n852 163.367
R1438 B.n337 B.t15 133.333
R1439 B.n153 B.t7 133.333
R1440 B.n331 B.t18 133.315
R1441 B.n146 B.t10 133.315
R1442 B.n569 B.n305 78.2614
R1443 B.n1060 B.n120 78.2614
R1444 B.n563 B.n306 71.676
R1445 B.n561 B.n308 71.676
R1446 B.n557 B.n556 71.676
R1447 B.n550 B.n310 71.676
R1448 B.n549 B.n548 71.676
R1449 B.n542 B.n312 71.676
R1450 B.n541 B.n540 71.676
R1451 B.n534 B.n314 71.676
R1452 B.n533 B.n532 71.676
R1453 B.n526 B.n316 71.676
R1454 B.n525 B.n524 71.676
R1455 B.n518 B.n318 71.676
R1456 B.n517 B.n516 71.676
R1457 B.n510 B.n320 71.676
R1458 B.n509 B.n508 71.676
R1459 B.n502 B.n322 71.676
R1460 B.n501 B.n500 71.676
R1461 B.n494 B.n324 71.676
R1462 B.n493 B.n492 71.676
R1463 B.n486 B.n326 71.676
R1464 B.n485 B.n484 71.676
R1465 B.n478 B.n328 71.676
R1466 B.n477 B.n476 71.676
R1467 B.n469 B.n330 71.676
R1468 B.n468 B.n467 71.676
R1469 B.n461 B.n334 71.676
R1470 B.n460 B.n459 71.676
R1471 B.n452 B.n336 71.676
R1472 B.n451 B.n450 71.676
R1473 B.n444 B.n340 71.676
R1474 B.n443 B.n442 71.676
R1475 B.n436 B.n342 71.676
R1476 B.n435 B.n434 71.676
R1477 B.n428 B.n344 71.676
R1478 B.n427 B.n426 71.676
R1479 B.n420 B.n346 71.676
R1480 B.n419 B.n418 71.676
R1481 B.n412 B.n348 71.676
R1482 B.n411 B.n410 71.676
R1483 B.n404 B.n350 71.676
R1484 B.n403 B.n402 71.676
R1485 B.n396 B.n352 71.676
R1486 B.n395 B.n394 71.676
R1487 B.n388 B.n354 71.676
R1488 B.n387 B.n386 71.676
R1489 B.n380 B.n356 71.676
R1490 B.n379 B.n378 71.676
R1491 B.n372 B.n358 71.676
R1492 B.n371 B.n370 71.676
R1493 B.n364 B.n360 71.676
R1494 B.n363 B.n362 71.676
R1495 B.n1054 B.n121 71.676
R1496 B.n1053 B.n1052 71.676
R1497 B.n1046 B.n123 71.676
R1498 B.n1045 B.n1044 71.676
R1499 B.n1038 B.n125 71.676
R1500 B.n1037 B.n1036 71.676
R1501 B.n1030 B.n127 71.676
R1502 B.n1029 B.n1028 71.676
R1503 B.n1022 B.n129 71.676
R1504 B.n1021 B.n1020 71.676
R1505 B.n1014 B.n131 71.676
R1506 B.n1013 B.n1012 71.676
R1507 B.n1006 B.n133 71.676
R1508 B.n1005 B.n1004 71.676
R1509 B.n998 B.n135 71.676
R1510 B.n997 B.n996 71.676
R1511 B.n990 B.n137 71.676
R1512 B.n989 B.n988 71.676
R1513 B.n982 B.n139 71.676
R1514 B.n981 B.n980 71.676
R1515 B.n974 B.n141 71.676
R1516 B.n973 B.n972 71.676
R1517 B.n966 B.n143 71.676
R1518 B.n965 B.n964 71.676
R1519 B.n958 B.n145 71.676
R1520 B.n957 B.n956 71.676
R1521 B.n950 B.n150 71.676
R1522 B.n949 B.n948 71.676
R1523 B.n941 B.n152 71.676
R1524 B.n940 B.n939 71.676
R1525 B.n933 B.n156 71.676
R1526 B.n932 B.n931 71.676
R1527 B.n925 B.n158 71.676
R1528 B.n924 B.n923 71.676
R1529 B.n917 B.n160 71.676
R1530 B.n916 B.n915 71.676
R1531 B.n909 B.n162 71.676
R1532 B.n908 B.n907 71.676
R1533 B.n901 B.n164 71.676
R1534 B.n900 B.n899 71.676
R1535 B.n893 B.n166 71.676
R1536 B.n892 B.n891 71.676
R1537 B.n885 B.n168 71.676
R1538 B.n884 B.n883 71.676
R1539 B.n877 B.n170 71.676
R1540 B.n876 B.n875 71.676
R1541 B.n869 B.n172 71.676
R1542 B.n868 B.n867 71.676
R1543 B.n861 B.n174 71.676
R1544 B.n860 B.n859 71.676
R1545 B.n853 B.n176 71.676
R1546 B.n854 B.n853 71.676
R1547 B.n859 B.n858 71.676
R1548 B.n862 B.n861 71.676
R1549 B.n867 B.n866 71.676
R1550 B.n870 B.n869 71.676
R1551 B.n875 B.n874 71.676
R1552 B.n878 B.n877 71.676
R1553 B.n883 B.n882 71.676
R1554 B.n886 B.n885 71.676
R1555 B.n891 B.n890 71.676
R1556 B.n894 B.n893 71.676
R1557 B.n899 B.n898 71.676
R1558 B.n902 B.n901 71.676
R1559 B.n907 B.n906 71.676
R1560 B.n910 B.n909 71.676
R1561 B.n915 B.n914 71.676
R1562 B.n918 B.n917 71.676
R1563 B.n923 B.n922 71.676
R1564 B.n926 B.n925 71.676
R1565 B.n931 B.n930 71.676
R1566 B.n934 B.n933 71.676
R1567 B.n939 B.n938 71.676
R1568 B.n942 B.n941 71.676
R1569 B.n948 B.n947 71.676
R1570 B.n951 B.n950 71.676
R1571 B.n956 B.n955 71.676
R1572 B.n959 B.n958 71.676
R1573 B.n964 B.n963 71.676
R1574 B.n967 B.n966 71.676
R1575 B.n972 B.n971 71.676
R1576 B.n975 B.n974 71.676
R1577 B.n980 B.n979 71.676
R1578 B.n983 B.n982 71.676
R1579 B.n988 B.n987 71.676
R1580 B.n991 B.n990 71.676
R1581 B.n996 B.n995 71.676
R1582 B.n999 B.n998 71.676
R1583 B.n1004 B.n1003 71.676
R1584 B.n1007 B.n1006 71.676
R1585 B.n1012 B.n1011 71.676
R1586 B.n1015 B.n1014 71.676
R1587 B.n1020 B.n1019 71.676
R1588 B.n1023 B.n1022 71.676
R1589 B.n1028 B.n1027 71.676
R1590 B.n1031 B.n1030 71.676
R1591 B.n1036 B.n1035 71.676
R1592 B.n1039 B.n1038 71.676
R1593 B.n1044 B.n1043 71.676
R1594 B.n1047 B.n1046 71.676
R1595 B.n1052 B.n1051 71.676
R1596 B.n1055 B.n1054 71.676
R1597 B.n564 B.n563 71.676
R1598 B.n558 B.n308 71.676
R1599 B.n556 B.n555 71.676
R1600 B.n551 B.n550 71.676
R1601 B.n548 B.n547 71.676
R1602 B.n543 B.n542 71.676
R1603 B.n540 B.n539 71.676
R1604 B.n535 B.n534 71.676
R1605 B.n532 B.n531 71.676
R1606 B.n527 B.n526 71.676
R1607 B.n524 B.n523 71.676
R1608 B.n519 B.n518 71.676
R1609 B.n516 B.n515 71.676
R1610 B.n511 B.n510 71.676
R1611 B.n508 B.n507 71.676
R1612 B.n503 B.n502 71.676
R1613 B.n500 B.n499 71.676
R1614 B.n495 B.n494 71.676
R1615 B.n492 B.n491 71.676
R1616 B.n487 B.n486 71.676
R1617 B.n484 B.n483 71.676
R1618 B.n479 B.n478 71.676
R1619 B.n476 B.n475 71.676
R1620 B.n470 B.n469 71.676
R1621 B.n467 B.n466 71.676
R1622 B.n462 B.n461 71.676
R1623 B.n459 B.n458 71.676
R1624 B.n453 B.n452 71.676
R1625 B.n450 B.n449 71.676
R1626 B.n445 B.n444 71.676
R1627 B.n442 B.n441 71.676
R1628 B.n437 B.n436 71.676
R1629 B.n434 B.n433 71.676
R1630 B.n429 B.n428 71.676
R1631 B.n426 B.n425 71.676
R1632 B.n421 B.n420 71.676
R1633 B.n418 B.n417 71.676
R1634 B.n413 B.n412 71.676
R1635 B.n410 B.n409 71.676
R1636 B.n405 B.n404 71.676
R1637 B.n402 B.n401 71.676
R1638 B.n397 B.n396 71.676
R1639 B.n394 B.n393 71.676
R1640 B.n389 B.n388 71.676
R1641 B.n386 B.n385 71.676
R1642 B.n381 B.n380 71.676
R1643 B.n378 B.n377 71.676
R1644 B.n373 B.n372 71.676
R1645 B.n370 B.n369 71.676
R1646 B.n365 B.n364 71.676
R1647 B.n362 B.n304 71.676
R1648 B.n338 B.t14 69.5271
R1649 B.n154 B.t8 69.5271
R1650 B.n332 B.t17 69.5093
R1651 B.n147 B.t11 69.5093
R1652 B.n338 B.n337 63.8066
R1653 B.n332 B.n331 63.8066
R1654 B.n147 B.n146 63.8066
R1655 B.n154 B.n153 63.8066
R1656 B.n455 B.n338 59.5399
R1657 B.n473 B.n332 59.5399
R1658 B.n148 B.n147 59.5399
R1659 B.n945 B.n154 59.5399
R1660 B.n569 B.n301 39.4208
R1661 B.n575 B.n301 39.4208
R1662 B.n575 B.n297 39.4208
R1663 B.n581 B.n297 39.4208
R1664 B.n581 B.n293 39.4208
R1665 B.n588 B.n293 39.4208
R1666 B.n588 B.n587 39.4208
R1667 B.n594 B.n286 39.4208
R1668 B.n600 B.n286 39.4208
R1669 B.n600 B.n282 39.4208
R1670 B.n606 B.n282 39.4208
R1671 B.n606 B.n278 39.4208
R1672 B.n612 B.n278 39.4208
R1673 B.n612 B.n274 39.4208
R1674 B.n618 B.n274 39.4208
R1675 B.n618 B.n270 39.4208
R1676 B.n624 B.n270 39.4208
R1677 B.n624 B.n266 39.4208
R1678 B.n630 B.n266 39.4208
R1679 B.n636 B.n262 39.4208
R1680 B.n636 B.n258 39.4208
R1681 B.n642 B.n258 39.4208
R1682 B.n642 B.n254 39.4208
R1683 B.n648 B.n254 39.4208
R1684 B.n648 B.n250 39.4208
R1685 B.n654 B.n250 39.4208
R1686 B.n654 B.n246 39.4208
R1687 B.n660 B.n246 39.4208
R1688 B.n666 B.n242 39.4208
R1689 B.n666 B.n238 39.4208
R1690 B.n672 B.n238 39.4208
R1691 B.n672 B.n234 39.4208
R1692 B.n678 B.n234 39.4208
R1693 B.n678 B.n230 39.4208
R1694 B.n684 B.n230 39.4208
R1695 B.n684 B.n226 39.4208
R1696 B.n690 B.n226 39.4208
R1697 B.n696 B.n222 39.4208
R1698 B.n696 B.n218 39.4208
R1699 B.n702 B.n218 39.4208
R1700 B.n702 B.n214 39.4208
R1701 B.n708 B.n214 39.4208
R1702 B.n708 B.n209 39.4208
R1703 B.n714 B.n209 39.4208
R1704 B.n714 B.n210 39.4208
R1705 B.n720 B.n202 39.4208
R1706 B.n726 B.n202 39.4208
R1707 B.n726 B.n198 39.4208
R1708 B.n732 B.n198 39.4208
R1709 B.n732 B.n194 39.4208
R1710 B.n738 B.n194 39.4208
R1711 B.n738 B.n190 39.4208
R1712 B.n745 B.n190 39.4208
R1713 B.n745 B.n744 39.4208
R1714 B.n751 B.n183 39.4208
R1715 B.n758 B.n183 39.4208
R1716 B.n758 B.n179 39.4208
R1717 B.n764 B.n179 39.4208
R1718 B.n764 B.n4 39.4208
R1719 B.n1190 B.n4 39.4208
R1720 B.n1190 B.n1189 39.4208
R1721 B.n1189 B.n1188 39.4208
R1722 B.n1188 B.n8 39.4208
R1723 B.n1182 B.n8 39.4208
R1724 B.n1182 B.n1181 39.4208
R1725 B.n1181 B.n1180 39.4208
R1726 B.n1174 B.n18 39.4208
R1727 B.n1174 B.n1173 39.4208
R1728 B.n1173 B.n1172 39.4208
R1729 B.n1172 B.n22 39.4208
R1730 B.n1166 B.n22 39.4208
R1731 B.n1166 B.n1165 39.4208
R1732 B.n1165 B.n1164 39.4208
R1733 B.n1164 B.n29 39.4208
R1734 B.n1158 B.n29 39.4208
R1735 B.n1157 B.n1156 39.4208
R1736 B.n1156 B.n36 39.4208
R1737 B.n1150 B.n36 39.4208
R1738 B.n1150 B.n1149 39.4208
R1739 B.n1149 B.n1148 39.4208
R1740 B.n1148 B.n43 39.4208
R1741 B.n1142 B.n43 39.4208
R1742 B.n1142 B.n1141 39.4208
R1743 B.n1140 B.n50 39.4208
R1744 B.n1134 B.n50 39.4208
R1745 B.n1134 B.n1133 39.4208
R1746 B.n1133 B.n1132 39.4208
R1747 B.n1132 B.n57 39.4208
R1748 B.n1126 B.n57 39.4208
R1749 B.n1126 B.n1125 39.4208
R1750 B.n1125 B.n1124 39.4208
R1751 B.n1124 B.n64 39.4208
R1752 B.n1118 B.n1117 39.4208
R1753 B.n1117 B.n1116 39.4208
R1754 B.n1116 B.n71 39.4208
R1755 B.n1110 B.n71 39.4208
R1756 B.n1110 B.n1109 39.4208
R1757 B.n1109 B.n1108 39.4208
R1758 B.n1108 B.n78 39.4208
R1759 B.n1102 B.n78 39.4208
R1760 B.n1102 B.n1101 39.4208
R1761 B.n1100 B.n85 39.4208
R1762 B.n1094 B.n85 39.4208
R1763 B.n1094 B.n1093 39.4208
R1764 B.n1093 B.n1092 39.4208
R1765 B.n1092 B.n92 39.4208
R1766 B.n1086 B.n92 39.4208
R1767 B.n1086 B.n1085 39.4208
R1768 B.n1085 B.n1084 39.4208
R1769 B.n1084 B.n99 39.4208
R1770 B.n1078 B.n99 39.4208
R1771 B.n1078 B.n1077 39.4208
R1772 B.n1077 B.n1076 39.4208
R1773 B.n1070 B.n109 39.4208
R1774 B.n1070 B.n1069 39.4208
R1775 B.n1069 B.n1068 39.4208
R1776 B.n1068 B.n113 39.4208
R1777 B.n1062 B.n113 39.4208
R1778 B.n1062 B.n1061 39.4208
R1779 B.n1061 B.n1060 39.4208
R1780 B.n587 B.t13 38.2614
R1781 B.n109 B.t6 38.2614
R1782 B.n210 B.t20 34.7831
R1783 B.t1 B.n1157 34.7831
R1784 B.n630 B.t0 33.6237
R1785 B.t21 B.n1100 33.6237
R1786 B.n1058 B.n1057 33.2493
R1787 B.n851 B.n850 33.2493
R1788 B.n571 B.n303 33.2493
R1789 B.n567 B.n566 33.2493
R1790 B.t22 B.n222 31.3048
R1791 B.n1141 B.t4 31.3048
R1792 B.n744 B.t23 22.0295
R1793 B.n18 B.t3 22.0295
R1794 B.n660 B.t2 20.8701
R1795 B.n1118 B.t19 20.8701
R1796 B.t2 B.n242 18.5512
R1797 B.t19 B.n64 18.5512
R1798 B B.n1192 18.0485
R1799 B.n751 B.t23 17.3918
R1800 B.n1180 B.t3 17.3918
R1801 B.n1057 B.n1056 10.6151
R1802 B.n1056 B.n122 10.6151
R1803 B.n1050 B.n122 10.6151
R1804 B.n1050 B.n1049 10.6151
R1805 B.n1049 B.n1048 10.6151
R1806 B.n1048 B.n124 10.6151
R1807 B.n1042 B.n124 10.6151
R1808 B.n1042 B.n1041 10.6151
R1809 B.n1041 B.n1040 10.6151
R1810 B.n1040 B.n126 10.6151
R1811 B.n1034 B.n126 10.6151
R1812 B.n1034 B.n1033 10.6151
R1813 B.n1033 B.n1032 10.6151
R1814 B.n1032 B.n128 10.6151
R1815 B.n1026 B.n128 10.6151
R1816 B.n1026 B.n1025 10.6151
R1817 B.n1025 B.n1024 10.6151
R1818 B.n1024 B.n130 10.6151
R1819 B.n1018 B.n130 10.6151
R1820 B.n1018 B.n1017 10.6151
R1821 B.n1017 B.n1016 10.6151
R1822 B.n1016 B.n132 10.6151
R1823 B.n1010 B.n132 10.6151
R1824 B.n1010 B.n1009 10.6151
R1825 B.n1009 B.n1008 10.6151
R1826 B.n1008 B.n134 10.6151
R1827 B.n1002 B.n134 10.6151
R1828 B.n1002 B.n1001 10.6151
R1829 B.n1001 B.n1000 10.6151
R1830 B.n1000 B.n136 10.6151
R1831 B.n994 B.n136 10.6151
R1832 B.n994 B.n993 10.6151
R1833 B.n993 B.n992 10.6151
R1834 B.n992 B.n138 10.6151
R1835 B.n986 B.n138 10.6151
R1836 B.n986 B.n985 10.6151
R1837 B.n985 B.n984 10.6151
R1838 B.n984 B.n140 10.6151
R1839 B.n978 B.n140 10.6151
R1840 B.n978 B.n977 10.6151
R1841 B.n977 B.n976 10.6151
R1842 B.n976 B.n142 10.6151
R1843 B.n970 B.n142 10.6151
R1844 B.n970 B.n969 10.6151
R1845 B.n969 B.n968 10.6151
R1846 B.n968 B.n144 10.6151
R1847 B.n962 B.n961 10.6151
R1848 B.n961 B.n960 10.6151
R1849 B.n960 B.n149 10.6151
R1850 B.n954 B.n149 10.6151
R1851 B.n954 B.n953 10.6151
R1852 B.n953 B.n952 10.6151
R1853 B.n952 B.n151 10.6151
R1854 B.n946 B.n151 10.6151
R1855 B.n944 B.n943 10.6151
R1856 B.n943 B.n155 10.6151
R1857 B.n937 B.n155 10.6151
R1858 B.n937 B.n936 10.6151
R1859 B.n936 B.n935 10.6151
R1860 B.n935 B.n157 10.6151
R1861 B.n929 B.n157 10.6151
R1862 B.n929 B.n928 10.6151
R1863 B.n928 B.n927 10.6151
R1864 B.n927 B.n159 10.6151
R1865 B.n921 B.n159 10.6151
R1866 B.n921 B.n920 10.6151
R1867 B.n920 B.n919 10.6151
R1868 B.n919 B.n161 10.6151
R1869 B.n913 B.n161 10.6151
R1870 B.n913 B.n912 10.6151
R1871 B.n912 B.n911 10.6151
R1872 B.n911 B.n163 10.6151
R1873 B.n905 B.n163 10.6151
R1874 B.n905 B.n904 10.6151
R1875 B.n904 B.n903 10.6151
R1876 B.n903 B.n165 10.6151
R1877 B.n897 B.n165 10.6151
R1878 B.n897 B.n896 10.6151
R1879 B.n896 B.n895 10.6151
R1880 B.n895 B.n167 10.6151
R1881 B.n889 B.n167 10.6151
R1882 B.n889 B.n888 10.6151
R1883 B.n888 B.n887 10.6151
R1884 B.n887 B.n169 10.6151
R1885 B.n881 B.n169 10.6151
R1886 B.n881 B.n880 10.6151
R1887 B.n880 B.n879 10.6151
R1888 B.n879 B.n171 10.6151
R1889 B.n873 B.n171 10.6151
R1890 B.n873 B.n872 10.6151
R1891 B.n872 B.n871 10.6151
R1892 B.n871 B.n173 10.6151
R1893 B.n865 B.n173 10.6151
R1894 B.n865 B.n864 10.6151
R1895 B.n864 B.n863 10.6151
R1896 B.n863 B.n175 10.6151
R1897 B.n857 B.n175 10.6151
R1898 B.n857 B.n856 10.6151
R1899 B.n856 B.n855 10.6151
R1900 B.n855 B.n851 10.6151
R1901 B.n572 B.n571 10.6151
R1902 B.n573 B.n572 10.6151
R1903 B.n573 B.n295 10.6151
R1904 B.n583 B.n295 10.6151
R1905 B.n584 B.n583 10.6151
R1906 B.n585 B.n584 10.6151
R1907 B.n585 B.n288 10.6151
R1908 B.n596 B.n288 10.6151
R1909 B.n597 B.n596 10.6151
R1910 B.n598 B.n597 10.6151
R1911 B.n598 B.n280 10.6151
R1912 B.n608 B.n280 10.6151
R1913 B.n609 B.n608 10.6151
R1914 B.n610 B.n609 10.6151
R1915 B.n610 B.n272 10.6151
R1916 B.n620 B.n272 10.6151
R1917 B.n621 B.n620 10.6151
R1918 B.n622 B.n621 10.6151
R1919 B.n622 B.n264 10.6151
R1920 B.n632 B.n264 10.6151
R1921 B.n633 B.n632 10.6151
R1922 B.n634 B.n633 10.6151
R1923 B.n634 B.n256 10.6151
R1924 B.n644 B.n256 10.6151
R1925 B.n645 B.n644 10.6151
R1926 B.n646 B.n645 10.6151
R1927 B.n646 B.n248 10.6151
R1928 B.n656 B.n248 10.6151
R1929 B.n657 B.n656 10.6151
R1930 B.n658 B.n657 10.6151
R1931 B.n658 B.n240 10.6151
R1932 B.n668 B.n240 10.6151
R1933 B.n669 B.n668 10.6151
R1934 B.n670 B.n669 10.6151
R1935 B.n670 B.n232 10.6151
R1936 B.n680 B.n232 10.6151
R1937 B.n681 B.n680 10.6151
R1938 B.n682 B.n681 10.6151
R1939 B.n682 B.n224 10.6151
R1940 B.n692 B.n224 10.6151
R1941 B.n693 B.n692 10.6151
R1942 B.n694 B.n693 10.6151
R1943 B.n694 B.n216 10.6151
R1944 B.n704 B.n216 10.6151
R1945 B.n705 B.n704 10.6151
R1946 B.n706 B.n705 10.6151
R1947 B.n706 B.n207 10.6151
R1948 B.n716 B.n207 10.6151
R1949 B.n717 B.n716 10.6151
R1950 B.n718 B.n717 10.6151
R1951 B.n718 B.n200 10.6151
R1952 B.n728 B.n200 10.6151
R1953 B.n729 B.n728 10.6151
R1954 B.n730 B.n729 10.6151
R1955 B.n730 B.n192 10.6151
R1956 B.n740 B.n192 10.6151
R1957 B.n741 B.n740 10.6151
R1958 B.n742 B.n741 10.6151
R1959 B.n742 B.n185 10.6151
R1960 B.n753 B.n185 10.6151
R1961 B.n754 B.n753 10.6151
R1962 B.n756 B.n754 10.6151
R1963 B.n756 B.n755 10.6151
R1964 B.n755 B.n177 10.6151
R1965 B.n767 B.n177 10.6151
R1966 B.n768 B.n767 10.6151
R1967 B.n769 B.n768 10.6151
R1968 B.n770 B.n769 10.6151
R1969 B.n772 B.n770 10.6151
R1970 B.n773 B.n772 10.6151
R1971 B.n774 B.n773 10.6151
R1972 B.n775 B.n774 10.6151
R1973 B.n777 B.n775 10.6151
R1974 B.n778 B.n777 10.6151
R1975 B.n779 B.n778 10.6151
R1976 B.n780 B.n779 10.6151
R1977 B.n782 B.n780 10.6151
R1978 B.n783 B.n782 10.6151
R1979 B.n784 B.n783 10.6151
R1980 B.n785 B.n784 10.6151
R1981 B.n787 B.n785 10.6151
R1982 B.n788 B.n787 10.6151
R1983 B.n789 B.n788 10.6151
R1984 B.n790 B.n789 10.6151
R1985 B.n792 B.n790 10.6151
R1986 B.n793 B.n792 10.6151
R1987 B.n794 B.n793 10.6151
R1988 B.n795 B.n794 10.6151
R1989 B.n797 B.n795 10.6151
R1990 B.n798 B.n797 10.6151
R1991 B.n799 B.n798 10.6151
R1992 B.n800 B.n799 10.6151
R1993 B.n802 B.n800 10.6151
R1994 B.n803 B.n802 10.6151
R1995 B.n804 B.n803 10.6151
R1996 B.n805 B.n804 10.6151
R1997 B.n807 B.n805 10.6151
R1998 B.n808 B.n807 10.6151
R1999 B.n809 B.n808 10.6151
R2000 B.n810 B.n809 10.6151
R2001 B.n812 B.n810 10.6151
R2002 B.n813 B.n812 10.6151
R2003 B.n814 B.n813 10.6151
R2004 B.n815 B.n814 10.6151
R2005 B.n817 B.n815 10.6151
R2006 B.n818 B.n817 10.6151
R2007 B.n819 B.n818 10.6151
R2008 B.n820 B.n819 10.6151
R2009 B.n822 B.n820 10.6151
R2010 B.n823 B.n822 10.6151
R2011 B.n824 B.n823 10.6151
R2012 B.n825 B.n824 10.6151
R2013 B.n827 B.n825 10.6151
R2014 B.n828 B.n827 10.6151
R2015 B.n829 B.n828 10.6151
R2016 B.n830 B.n829 10.6151
R2017 B.n832 B.n830 10.6151
R2018 B.n833 B.n832 10.6151
R2019 B.n834 B.n833 10.6151
R2020 B.n835 B.n834 10.6151
R2021 B.n837 B.n835 10.6151
R2022 B.n838 B.n837 10.6151
R2023 B.n839 B.n838 10.6151
R2024 B.n840 B.n839 10.6151
R2025 B.n842 B.n840 10.6151
R2026 B.n843 B.n842 10.6151
R2027 B.n844 B.n843 10.6151
R2028 B.n845 B.n844 10.6151
R2029 B.n847 B.n845 10.6151
R2030 B.n848 B.n847 10.6151
R2031 B.n849 B.n848 10.6151
R2032 B.n850 B.n849 10.6151
R2033 B.n566 B.n565 10.6151
R2034 B.n565 B.n307 10.6151
R2035 B.n560 B.n307 10.6151
R2036 B.n560 B.n559 10.6151
R2037 B.n559 B.n309 10.6151
R2038 B.n554 B.n309 10.6151
R2039 B.n554 B.n553 10.6151
R2040 B.n553 B.n552 10.6151
R2041 B.n552 B.n311 10.6151
R2042 B.n546 B.n311 10.6151
R2043 B.n546 B.n545 10.6151
R2044 B.n545 B.n544 10.6151
R2045 B.n544 B.n313 10.6151
R2046 B.n538 B.n313 10.6151
R2047 B.n538 B.n537 10.6151
R2048 B.n537 B.n536 10.6151
R2049 B.n536 B.n315 10.6151
R2050 B.n530 B.n315 10.6151
R2051 B.n530 B.n529 10.6151
R2052 B.n529 B.n528 10.6151
R2053 B.n528 B.n317 10.6151
R2054 B.n522 B.n317 10.6151
R2055 B.n522 B.n521 10.6151
R2056 B.n521 B.n520 10.6151
R2057 B.n520 B.n319 10.6151
R2058 B.n514 B.n319 10.6151
R2059 B.n514 B.n513 10.6151
R2060 B.n513 B.n512 10.6151
R2061 B.n512 B.n321 10.6151
R2062 B.n506 B.n321 10.6151
R2063 B.n506 B.n505 10.6151
R2064 B.n505 B.n504 10.6151
R2065 B.n504 B.n323 10.6151
R2066 B.n498 B.n323 10.6151
R2067 B.n498 B.n497 10.6151
R2068 B.n497 B.n496 10.6151
R2069 B.n496 B.n325 10.6151
R2070 B.n490 B.n325 10.6151
R2071 B.n490 B.n489 10.6151
R2072 B.n489 B.n488 10.6151
R2073 B.n488 B.n327 10.6151
R2074 B.n482 B.n327 10.6151
R2075 B.n482 B.n481 10.6151
R2076 B.n481 B.n480 10.6151
R2077 B.n480 B.n329 10.6151
R2078 B.n474 B.n329 10.6151
R2079 B.n472 B.n471 10.6151
R2080 B.n471 B.n333 10.6151
R2081 B.n465 B.n333 10.6151
R2082 B.n465 B.n464 10.6151
R2083 B.n464 B.n463 10.6151
R2084 B.n463 B.n335 10.6151
R2085 B.n457 B.n335 10.6151
R2086 B.n457 B.n456 10.6151
R2087 B.n454 B.n339 10.6151
R2088 B.n448 B.n339 10.6151
R2089 B.n448 B.n447 10.6151
R2090 B.n447 B.n446 10.6151
R2091 B.n446 B.n341 10.6151
R2092 B.n440 B.n341 10.6151
R2093 B.n440 B.n439 10.6151
R2094 B.n439 B.n438 10.6151
R2095 B.n438 B.n343 10.6151
R2096 B.n432 B.n343 10.6151
R2097 B.n432 B.n431 10.6151
R2098 B.n431 B.n430 10.6151
R2099 B.n430 B.n345 10.6151
R2100 B.n424 B.n345 10.6151
R2101 B.n424 B.n423 10.6151
R2102 B.n423 B.n422 10.6151
R2103 B.n422 B.n347 10.6151
R2104 B.n416 B.n347 10.6151
R2105 B.n416 B.n415 10.6151
R2106 B.n415 B.n414 10.6151
R2107 B.n414 B.n349 10.6151
R2108 B.n408 B.n349 10.6151
R2109 B.n408 B.n407 10.6151
R2110 B.n407 B.n406 10.6151
R2111 B.n406 B.n351 10.6151
R2112 B.n400 B.n351 10.6151
R2113 B.n400 B.n399 10.6151
R2114 B.n399 B.n398 10.6151
R2115 B.n398 B.n353 10.6151
R2116 B.n392 B.n353 10.6151
R2117 B.n392 B.n391 10.6151
R2118 B.n391 B.n390 10.6151
R2119 B.n390 B.n355 10.6151
R2120 B.n384 B.n355 10.6151
R2121 B.n384 B.n383 10.6151
R2122 B.n383 B.n382 10.6151
R2123 B.n382 B.n357 10.6151
R2124 B.n376 B.n357 10.6151
R2125 B.n376 B.n375 10.6151
R2126 B.n375 B.n374 10.6151
R2127 B.n374 B.n359 10.6151
R2128 B.n368 B.n359 10.6151
R2129 B.n368 B.n367 10.6151
R2130 B.n367 B.n366 10.6151
R2131 B.n366 B.n361 10.6151
R2132 B.n361 B.n303 10.6151
R2133 B.n567 B.n299 10.6151
R2134 B.n577 B.n299 10.6151
R2135 B.n578 B.n577 10.6151
R2136 B.n579 B.n578 10.6151
R2137 B.n579 B.n291 10.6151
R2138 B.n590 B.n291 10.6151
R2139 B.n591 B.n590 10.6151
R2140 B.n592 B.n591 10.6151
R2141 B.n592 B.n284 10.6151
R2142 B.n602 B.n284 10.6151
R2143 B.n603 B.n602 10.6151
R2144 B.n604 B.n603 10.6151
R2145 B.n604 B.n276 10.6151
R2146 B.n614 B.n276 10.6151
R2147 B.n615 B.n614 10.6151
R2148 B.n616 B.n615 10.6151
R2149 B.n616 B.n268 10.6151
R2150 B.n626 B.n268 10.6151
R2151 B.n627 B.n626 10.6151
R2152 B.n628 B.n627 10.6151
R2153 B.n628 B.n260 10.6151
R2154 B.n638 B.n260 10.6151
R2155 B.n639 B.n638 10.6151
R2156 B.n640 B.n639 10.6151
R2157 B.n640 B.n252 10.6151
R2158 B.n650 B.n252 10.6151
R2159 B.n651 B.n650 10.6151
R2160 B.n652 B.n651 10.6151
R2161 B.n652 B.n244 10.6151
R2162 B.n662 B.n244 10.6151
R2163 B.n663 B.n662 10.6151
R2164 B.n664 B.n663 10.6151
R2165 B.n664 B.n236 10.6151
R2166 B.n674 B.n236 10.6151
R2167 B.n675 B.n674 10.6151
R2168 B.n676 B.n675 10.6151
R2169 B.n676 B.n228 10.6151
R2170 B.n686 B.n228 10.6151
R2171 B.n687 B.n686 10.6151
R2172 B.n688 B.n687 10.6151
R2173 B.n688 B.n220 10.6151
R2174 B.n698 B.n220 10.6151
R2175 B.n699 B.n698 10.6151
R2176 B.n700 B.n699 10.6151
R2177 B.n700 B.n212 10.6151
R2178 B.n710 B.n212 10.6151
R2179 B.n711 B.n710 10.6151
R2180 B.n712 B.n711 10.6151
R2181 B.n712 B.n204 10.6151
R2182 B.n722 B.n204 10.6151
R2183 B.n723 B.n722 10.6151
R2184 B.n724 B.n723 10.6151
R2185 B.n724 B.n196 10.6151
R2186 B.n734 B.n196 10.6151
R2187 B.n735 B.n734 10.6151
R2188 B.n736 B.n735 10.6151
R2189 B.n736 B.n188 10.6151
R2190 B.n747 B.n188 10.6151
R2191 B.n748 B.n747 10.6151
R2192 B.n749 B.n748 10.6151
R2193 B.n749 B.n181 10.6151
R2194 B.n760 B.n181 10.6151
R2195 B.n761 B.n760 10.6151
R2196 B.n762 B.n761 10.6151
R2197 B.n762 B.n0 10.6151
R2198 B.n1186 B.n1 10.6151
R2199 B.n1186 B.n1185 10.6151
R2200 B.n1185 B.n1184 10.6151
R2201 B.n1184 B.n10 10.6151
R2202 B.n1178 B.n10 10.6151
R2203 B.n1178 B.n1177 10.6151
R2204 B.n1177 B.n1176 10.6151
R2205 B.n1176 B.n16 10.6151
R2206 B.n1170 B.n16 10.6151
R2207 B.n1170 B.n1169 10.6151
R2208 B.n1169 B.n1168 10.6151
R2209 B.n1168 B.n24 10.6151
R2210 B.n1162 B.n24 10.6151
R2211 B.n1162 B.n1161 10.6151
R2212 B.n1161 B.n1160 10.6151
R2213 B.n1160 B.n31 10.6151
R2214 B.n1154 B.n31 10.6151
R2215 B.n1154 B.n1153 10.6151
R2216 B.n1153 B.n1152 10.6151
R2217 B.n1152 B.n38 10.6151
R2218 B.n1146 B.n38 10.6151
R2219 B.n1146 B.n1145 10.6151
R2220 B.n1145 B.n1144 10.6151
R2221 B.n1144 B.n45 10.6151
R2222 B.n1138 B.n45 10.6151
R2223 B.n1138 B.n1137 10.6151
R2224 B.n1137 B.n1136 10.6151
R2225 B.n1136 B.n52 10.6151
R2226 B.n1130 B.n52 10.6151
R2227 B.n1130 B.n1129 10.6151
R2228 B.n1129 B.n1128 10.6151
R2229 B.n1128 B.n59 10.6151
R2230 B.n1122 B.n59 10.6151
R2231 B.n1122 B.n1121 10.6151
R2232 B.n1121 B.n1120 10.6151
R2233 B.n1120 B.n66 10.6151
R2234 B.n1114 B.n66 10.6151
R2235 B.n1114 B.n1113 10.6151
R2236 B.n1113 B.n1112 10.6151
R2237 B.n1112 B.n73 10.6151
R2238 B.n1106 B.n73 10.6151
R2239 B.n1106 B.n1105 10.6151
R2240 B.n1105 B.n1104 10.6151
R2241 B.n1104 B.n80 10.6151
R2242 B.n1098 B.n80 10.6151
R2243 B.n1098 B.n1097 10.6151
R2244 B.n1097 B.n1096 10.6151
R2245 B.n1096 B.n87 10.6151
R2246 B.n1090 B.n87 10.6151
R2247 B.n1090 B.n1089 10.6151
R2248 B.n1089 B.n1088 10.6151
R2249 B.n1088 B.n94 10.6151
R2250 B.n1082 B.n94 10.6151
R2251 B.n1082 B.n1081 10.6151
R2252 B.n1081 B.n1080 10.6151
R2253 B.n1080 B.n101 10.6151
R2254 B.n1074 B.n101 10.6151
R2255 B.n1074 B.n1073 10.6151
R2256 B.n1073 B.n1072 10.6151
R2257 B.n1072 B.n107 10.6151
R2258 B.n1066 B.n107 10.6151
R2259 B.n1066 B.n1065 10.6151
R2260 B.n1065 B.n1064 10.6151
R2261 B.n1064 B.n115 10.6151
R2262 B.n1058 B.n115 10.6151
R2263 B.n690 B.t22 8.11644
R2264 B.t4 B.n1140 8.11644
R2265 B.n962 B.n148 6.5566
R2266 B.n946 B.n945 6.5566
R2267 B.n473 B.n472 6.5566
R2268 B.n456 B.n455 6.5566
R2269 B.t0 B.n262 5.7976
R2270 B.n1101 B.t21 5.7976
R2271 B.n720 B.t20 4.63818
R2272 B.n1158 B.t1 4.63818
R2273 B.n148 B.n144 4.05904
R2274 B.n945 B.n944 4.05904
R2275 B.n474 B.n473 4.05904
R2276 B.n455 B.n454 4.05904
R2277 B.n1192 B.n0 2.81026
R2278 B.n1192 B.n1 2.81026
R2279 B.n594 B.t13 1.15992
R2280 B.n1076 B.t6 1.15992
R2281 VN.n90 VN.n89 161.3
R2282 VN.n88 VN.n47 161.3
R2283 VN.n87 VN.n86 161.3
R2284 VN.n85 VN.n48 161.3
R2285 VN.n84 VN.n83 161.3
R2286 VN.n82 VN.n49 161.3
R2287 VN.n80 VN.n79 161.3
R2288 VN.n78 VN.n50 161.3
R2289 VN.n77 VN.n76 161.3
R2290 VN.n75 VN.n51 161.3
R2291 VN.n74 VN.n73 161.3
R2292 VN.n72 VN.n52 161.3
R2293 VN.n71 VN.n70 161.3
R2294 VN.n68 VN.n53 161.3
R2295 VN.n67 VN.n66 161.3
R2296 VN.n65 VN.n54 161.3
R2297 VN.n64 VN.n63 161.3
R2298 VN.n62 VN.n55 161.3
R2299 VN.n61 VN.n60 161.3
R2300 VN.n59 VN.n56 161.3
R2301 VN.n44 VN.n43 161.3
R2302 VN.n42 VN.n1 161.3
R2303 VN.n41 VN.n40 161.3
R2304 VN.n39 VN.n2 161.3
R2305 VN.n38 VN.n37 161.3
R2306 VN.n36 VN.n3 161.3
R2307 VN.n34 VN.n33 161.3
R2308 VN.n32 VN.n4 161.3
R2309 VN.n31 VN.n30 161.3
R2310 VN.n29 VN.n5 161.3
R2311 VN.n28 VN.n27 161.3
R2312 VN.n26 VN.n6 161.3
R2313 VN.n25 VN.n24 161.3
R2314 VN.n22 VN.n7 161.3
R2315 VN.n21 VN.n20 161.3
R2316 VN.n19 VN.n8 161.3
R2317 VN.n18 VN.n17 161.3
R2318 VN.n16 VN.n9 161.3
R2319 VN.n15 VN.n14 161.3
R2320 VN.n13 VN.n10 161.3
R2321 VN.n58 VN.t5 143.061
R2322 VN.n12 VN.t7 143.061
R2323 VN.n11 VN.t3 111.544
R2324 VN.n23 VN.t4 111.544
R2325 VN.n35 VN.t2 111.544
R2326 VN.n0 VN.t9 111.544
R2327 VN.n57 VN.t0 111.544
R2328 VN.n69 VN.t6 111.544
R2329 VN.n81 VN.t8 111.544
R2330 VN.n46 VN.t1 111.544
R2331 VN.n45 VN.n0 74.0149
R2332 VN.n91 VN.n46 74.0149
R2333 VN.n12 VN.n11 71.6401
R2334 VN.n58 VN.n57 71.6401
R2335 VN VN.n91 56.5777
R2336 VN.n41 VN.n2 56.5617
R2337 VN.n87 VN.n48 56.5617
R2338 VN.n17 VN.n8 50.7491
R2339 VN.n29 VN.n28 50.7491
R2340 VN.n63 VN.n54 50.7491
R2341 VN.n75 VN.n74 50.7491
R2342 VN.n17 VN.n16 30.405
R2343 VN.n30 VN.n29 30.405
R2344 VN.n63 VN.n62 30.405
R2345 VN.n76 VN.n75 30.405
R2346 VN.n15 VN.n10 24.5923
R2347 VN.n16 VN.n15 24.5923
R2348 VN.n21 VN.n8 24.5923
R2349 VN.n22 VN.n21 24.5923
R2350 VN.n24 VN.n6 24.5923
R2351 VN.n28 VN.n6 24.5923
R2352 VN.n30 VN.n4 24.5923
R2353 VN.n34 VN.n4 24.5923
R2354 VN.n37 VN.n36 24.5923
R2355 VN.n37 VN.n2 24.5923
R2356 VN.n42 VN.n41 24.5923
R2357 VN.n43 VN.n42 24.5923
R2358 VN.n62 VN.n61 24.5923
R2359 VN.n61 VN.n56 24.5923
R2360 VN.n74 VN.n52 24.5923
R2361 VN.n70 VN.n52 24.5923
R2362 VN.n68 VN.n67 24.5923
R2363 VN.n67 VN.n54 24.5923
R2364 VN.n83 VN.n48 24.5923
R2365 VN.n83 VN.n82 24.5923
R2366 VN.n80 VN.n50 24.5923
R2367 VN.n76 VN.n50 24.5923
R2368 VN.n89 VN.n88 24.5923
R2369 VN.n88 VN.n87 24.5923
R2370 VN.n36 VN.n35 22.625
R2371 VN.n82 VN.n81 22.625
R2372 VN.n43 VN.n0 16.2311
R2373 VN.n89 VN.n46 16.2311
R2374 VN.n23 VN.n22 12.2964
R2375 VN.n24 VN.n23 12.2964
R2376 VN.n70 VN.n69 12.2964
R2377 VN.n69 VN.n68 12.2964
R2378 VN.n59 VN.n58 5.81316
R2379 VN.n13 VN.n12 5.81316
R2380 VN.n11 VN.n10 1.96785
R2381 VN.n35 VN.n34 1.96785
R2382 VN.n57 VN.n56 1.96785
R2383 VN.n81 VN.n80 1.96785
R2384 VN.n91 VN.n90 0.354861
R2385 VN.n45 VN.n44 0.354861
R2386 VN VN.n45 0.267071
R2387 VN.n90 VN.n47 0.189894
R2388 VN.n86 VN.n47 0.189894
R2389 VN.n86 VN.n85 0.189894
R2390 VN.n85 VN.n84 0.189894
R2391 VN.n84 VN.n49 0.189894
R2392 VN.n79 VN.n49 0.189894
R2393 VN.n79 VN.n78 0.189894
R2394 VN.n78 VN.n77 0.189894
R2395 VN.n77 VN.n51 0.189894
R2396 VN.n73 VN.n51 0.189894
R2397 VN.n73 VN.n72 0.189894
R2398 VN.n72 VN.n71 0.189894
R2399 VN.n71 VN.n53 0.189894
R2400 VN.n66 VN.n53 0.189894
R2401 VN.n66 VN.n65 0.189894
R2402 VN.n65 VN.n64 0.189894
R2403 VN.n64 VN.n55 0.189894
R2404 VN.n60 VN.n55 0.189894
R2405 VN.n60 VN.n59 0.189894
R2406 VN.n14 VN.n13 0.189894
R2407 VN.n14 VN.n9 0.189894
R2408 VN.n18 VN.n9 0.189894
R2409 VN.n19 VN.n18 0.189894
R2410 VN.n20 VN.n19 0.189894
R2411 VN.n20 VN.n7 0.189894
R2412 VN.n25 VN.n7 0.189894
R2413 VN.n26 VN.n25 0.189894
R2414 VN.n27 VN.n26 0.189894
R2415 VN.n27 VN.n5 0.189894
R2416 VN.n31 VN.n5 0.189894
R2417 VN.n32 VN.n31 0.189894
R2418 VN.n33 VN.n32 0.189894
R2419 VN.n33 VN.n3 0.189894
R2420 VN.n38 VN.n3 0.189894
R2421 VN.n39 VN.n38 0.189894
R2422 VN.n40 VN.n39 0.189894
R2423 VN.n40 VN.n1 0.189894
R2424 VN.n44 VN.n1 0.189894
R2425 VDD2.n1 VDD2.t2 68.0635
R2426 VDD2.n3 VDD2.n2 65.8539
R2427 VDD2 VDD2.n7 65.8511
R2428 VDD2.n4 VDD2.t8 65.2275
R2429 VDD2.n6 VDD2.n5 63.7823
R2430 VDD2.n1 VDD2.n0 63.7821
R2431 VDD2.n4 VDD2.n3 48.9976
R2432 VDD2.n6 VDD2.n4 2.83671
R2433 VDD2.n7 VDD2.t9 1.44576
R2434 VDD2.n7 VDD2.t4 1.44576
R2435 VDD2.n5 VDD2.t1 1.44576
R2436 VDD2.n5 VDD2.t3 1.44576
R2437 VDD2.n2 VDD2.t7 1.44576
R2438 VDD2.n2 VDD2.t0 1.44576
R2439 VDD2.n0 VDD2.t6 1.44576
R2440 VDD2.n0 VDD2.t5 1.44576
R2441 VDD2 VDD2.n6 0.767741
R2442 VDD2.n3 VDD2.n1 0.654206
C0 VDD1 VDD2 2.40936f
C1 VN VDD1 0.154566f
C2 VN VDD2 12.404599f
C3 VTAIL VDD1 11.243f
C4 VP VDD1 12.8759f
C5 VTAIL VDD2 11.296401f
C6 VN VTAIL 13.1265f
C7 VP VDD2 0.63001f
C8 VP VN 9.24191f
C9 VP VTAIL 13.1407f
C10 VDD2 B 7.926064f
C11 VDD1 B 7.902394f
C12 VTAIL B 9.177164f
C13 VN B 19.991749f
C14 VP B 18.53042f
C15 VDD2.t2 B 3.02272f
C16 VDD2.t6 B 0.2611f
C17 VDD2.t5 B 0.2611f
C18 VDD2.n0 B 2.35252f
C19 VDD2.n1 B 0.930579f
C20 VDD2.t7 B 0.2611f
C21 VDD2.t0 B 0.2611f
C22 VDD2.n2 B 2.37091f
C23 VDD2.n3 B 3.0813f
C24 VDD2.t8 B 3.00249f
C25 VDD2.n4 B 3.2678f
C26 VDD2.t1 B 0.2611f
C27 VDD2.t3 B 0.2611f
C28 VDD2.n5 B 2.35252f
C29 VDD2.n6 B 0.473283f
C30 VDD2.t9 B 0.2611f
C31 VDD2.t4 B 0.2611f
C32 VDD2.n7 B 2.37087f
C33 VN.t9 B 2.14557f
C34 VN.n0 B 0.821014f
C35 VN.n1 B 0.01935f
C36 VN.n2 B 0.024649f
C37 VN.n3 B 0.01935f
C38 VN.t2 B 2.14557f
C39 VN.n4 B 0.035883f
C40 VN.n5 B 0.01935f
C41 VN.n6 B 0.035883f
C42 VN.n7 B 0.01935f
C43 VN.t4 B 2.14557f
C44 VN.n8 B 0.035153f
C45 VN.n9 B 0.01935f
C46 VN.n10 B 0.019586f
C47 VN.t3 B 2.14557f
C48 VN.n11 B 0.804405f
C49 VN.t7 B 2.33841f
C50 VN.n12 B 0.782527f
C51 VN.n13 B 0.209207f
C52 VN.n14 B 0.01935f
C53 VN.n15 B 0.035883f
C54 VN.n16 B 0.038457f
C55 VN.n17 B 0.018531f
C56 VN.n18 B 0.01935f
C57 VN.n19 B 0.01935f
C58 VN.n20 B 0.01935f
C59 VN.n21 B 0.035883f
C60 VN.n22 B 0.027026f
C61 VN.n23 B 0.750741f
C62 VN.n24 B 0.027026f
C63 VN.n25 B 0.01935f
C64 VN.n26 B 0.01935f
C65 VN.n27 B 0.01935f
C66 VN.n28 B 0.035153f
C67 VN.n29 B 0.018531f
C68 VN.n30 B 0.038457f
C69 VN.n31 B 0.01935f
C70 VN.n32 B 0.01935f
C71 VN.n33 B 0.01935f
C72 VN.n34 B 0.019586f
C73 VN.n35 B 0.750741f
C74 VN.n36 B 0.034466f
C75 VN.n37 B 0.035883f
C76 VN.n38 B 0.01935f
C77 VN.n39 B 0.01935f
C78 VN.n40 B 0.01935f
C79 VN.n41 B 0.031609f
C80 VN.n42 B 0.035883f
C81 VN.n43 B 0.02986f
C82 VN.n44 B 0.031226f
C83 VN.n45 B 0.043047f
C84 VN.t1 B 2.14557f
C85 VN.n46 B 0.821014f
C86 VN.n47 B 0.01935f
C87 VN.n48 B 0.024649f
C88 VN.n49 B 0.01935f
C89 VN.t8 B 2.14557f
C90 VN.n50 B 0.035883f
C91 VN.n51 B 0.01935f
C92 VN.n52 B 0.035883f
C93 VN.n53 B 0.01935f
C94 VN.t6 B 2.14557f
C95 VN.n54 B 0.035153f
C96 VN.n55 B 0.01935f
C97 VN.n56 B 0.019586f
C98 VN.t5 B 2.33841f
C99 VN.t0 B 2.14557f
C100 VN.n57 B 0.804405f
C101 VN.n58 B 0.782527f
C102 VN.n59 B 0.209207f
C103 VN.n60 B 0.01935f
C104 VN.n61 B 0.035883f
C105 VN.n62 B 0.038457f
C106 VN.n63 B 0.018531f
C107 VN.n64 B 0.01935f
C108 VN.n65 B 0.01935f
C109 VN.n66 B 0.01935f
C110 VN.n67 B 0.035883f
C111 VN.n68 B 0.027026f
C112 VN.n69 B 0.750741f
C113 VN.n70 B 0.027026f
C114 VN.n71 B 0.01935f
C115 VN.n72 B 0.01935f
C116 VN.n73 B 0.01935f
C117 VN.n74 B 0.035153f
C118 VN.n75 B 0.018531f
C119 VN.n76 B 0.038457f
C120 VN.n77 B 0.01935f
C121 VN.n78 B 0.01935f
C122 VN.n79 B 0.01935f
C123 VN.n80 B 0.019586f
C124 VN.n81 B 0.750741f
C125 VN.n82 B 0.034466f
C126 VN.n83 B 0.035883f
C127 VN.n84 B 0.01935f
C128 VN.n85 B 0.01935f
C129 VN.n86 B 0.01935f
C130 VN.n87 B 0.031609f
C131 VN.n88 B 0.035883f
C132 VN.n89 B 0.02986f
C133 VN.n90 B 0.031226f
C134 VN.n91 B 1.30556f
C135 VDD1.t8 B 3.05861f
C136 VDD1.t2 B 0.264199f
C137 VDD1.t1 B 0.264199f
C138 VDD1.n0 B 2.38045f
C139 VDD1.n1 B 0.949686f
C140 VDD1.t4 B 3.05861f
C141 VDD1.t0 B 0.264199f
C142 VDD1.t9 B 0.264199f
C143 VDD1.n2 B 2.38045f
C144 VDD1.n3 B 0.941627f
C145 VDD1.t7 B 0.264199f
C146 VDD1.t5 B 0.264199f
C147 VDD1.n4 B 2.39906f
C148 VDD1.n5 B 3.25066f
C149 VDD1.t6 B 0.264199f
C150 VDD1.t3 B 0.264199f
C151 VDD1.n6 B 2.38045f
C152 VDD1.n7 B 3.3638f
C153 VTAIL.t3 B 0.267137f
C154 VTAIL.t1 B 0.267137f
C155 VTAIL.n0 B 2.33857f
C156 VTAIL.n1 B 0.556394f
C157 VTAIL.t16 B 2.98377f
C158 VTAIL.n2 B 0.691498f
C159 VTAIL.t19 B 0.267137f
C160 VTAIL.t17 B 0.267137f
C161 VTAIL.n3 B 2.33857f
C162 VTAIL.n4 B 0.68354f
C163 VTAIL.t11 B 0.267137f
C164 VTAIL.t15 B 0.267137f
C165 VTAIL.n5 B 2.33857f
C166 VTAIL.n6 B 2.18326f
C167 VTAIL.t0 B 0.267137f
C168 VTAIL.t2 B 0.267137f
C169 VTAIL.n7 B 2.33857f
C170 VTAIL.n8 B 2.18325f
C171 VTAIL.t8 B 0.267137f
C172 VTAIL.t6 B 0.267137f
C173 VTAIL.n9 B 2.33857f
C174 VTAIL.n10 B 0.683538f
C175 VTAIL.t9 B 2.98377f
C176 VTAIL.n11 B 0.691495f
C177 VTAIL.t18 B 0.267137f
C178 VTAIL.t14 B 0.267137f
C179 VTAIL.n12 B 2.33857f
C180 VTAIL.n13 B 0.608141f
C181 VTAIL.t10 B 0.267137f
C182 VTAIL.t13 B 0.267137f
C183 VTAIL.n14 B 2.33857f
C184 VTAIL.n15 B 0.683538f
C185 VTAIL.t12 B 2.98377f
C186 VTAIL.n16 B 2.04111f
C187 VTAIL.t7 B 2.98377f
C188 VTAIL.n17 B 2.04111f
C189 VTAIL.t4 B 0.267137f
C190 VTAIL.t5 B 0.267137f
C191 VTAIL.n18 B 2.33857f
C192 VTAIL.n19 B 0.509786f
C193 VP.t4 B 2.1782f
C194 VP.n0 B 0.833497f
C195 VP.n1 B 0.019645f
C196 VP.n2 B 0.025024f
C197 VP.n3 B 0.019645f
C198 VP.t2 B 2.1782f
C199 VP.n4 B 0.036429f
C200 VP.n5 B 0.019645f
C201 VP.n6 B 0.036429f
C202 VP.n7 B 0.019645f
C203 VP.t0 B 2.1782f
C204 VP.n8 B 0.035687f
C205 VP.n9 B 0.019645f
C206 VP.n10 B 0.019884f
C207 VP.n11 B 0.019645f
C208 VP.n12 B 0.032089f
C209 VP.n13 B 0.031701f
C210 VP.t5 B 2.1782f
C211 VP.t6 B 2.1782f
C212 VP.n14 B 0.833497f
C213 VP.n15 B 0.019645f
C214 VP.n16 B 0.025024f
C215 VP.n17 B 0.019645f
C216 VP.t3 B 2.1782f
C217 VP.n18 B 0.036429f
C218 VP.n19 B 0.019645f
C219 VP.n20 B 0.036429f
C220 VP.n21 B 0.019645f
C221 VP.t8 B 2.1782f
C222 VP.n22 B 0.035687f
C223 VP.n23 B 0.019645f
C224 VP.n24 B 0.019884f
C225 VP.t1 B 2.37397f
C226 VP.t7 B 2.1782f
C227 VP.n25 B 0.816636f
C228 VP.n26 B 0.794426f
C229 VP.n27 B 0.212389f
C230 VP.n28 B 0.019645f
C231 VP.n29 B 0.036429f
C232 VP.n30 B 0.039042f
C233 VP.n31 B 0.018812f
C234 VP.n32 B 0.019645f
C235 VP.n33 B 0.019645f
C236 VP.n34 B 0.019645f
C237 VP.n35 B 0.036429f
C238 VP.n36 B 0.027437f
C239 VP.n37 B 0.762156f
C240 VP.n38 B 0.027437f
C241 VP.n39 B 0.019645f
C242 VP.n40 B 0.019645f
C243 VP.n41 B 0.019645f
C244 VP.n42 B 0.035687f
C245 VP.n43 B 0.018812f
C246 VP.n44 B 0.039042f
C247 VP.n45 B 0.019645f
C248 VP.n46 B 0.019645f
C249 VP.n47 B 0.019645f
C250 VP.n48 B 0.019884f
C251 VP.n49 B 0.762156f
C252 VP.n50 B 0.03499f
C253 VP.n51 B 0.036429f
C254 VP.n52 B 0.019645f
C255 VP.n53 B 0.019645f
C256 VP.n54 B 0.019645f
C257 VP.n55 B 0.032089f
C258 VP.n56 B 0.036429f
C259 VP.n57 B 0.030314f
C260 VP.n58 B 0.031701f
C261 VP.n59 B 1.31768f
C262 VP.n60 B 1.33023f
C263 VP.n61 B 0.833497f
C264 VP.n62 B 0.030314f
C265 VP.n63 B 0.036429f
C266 VP.n64 B 0.019645f
C267 VP.n65 B 0.019645f
C268 VP.n66 B 0.019645f
C269 VP.n67 B 0.025024f
C270 VP.n68 B 0.036429f
C271 VP.t9 B 2.1782f
C272 VP.n69 B 0.762156f
C273 VP.n70 B 0.03499f
C274 VP.n71 B 0.019645f
C275 VP.n72 B 0.019645f
C276 VP.n73 B 0.019645f
C277 VP.n74 B 0.036429f
C278 VP.n75 B 0.039042f
C279 VP.n76 B 0.018812f
C280 VP.n77 B 0.019645f
C281 VP.n78 B 0.019645f
C282 VP.n79 B 0.019645f
C283 VP.n80 B 0.036429f
C284 VP.n81 B 0.027437f
C285 VP.n82 B 0.762156f
C286 VP.n83 B 0.027437f
C287 VP.n84 B 0.019645f
C288 VP.n85 B 0.019645f
C289 VP.n86 B 0.019645f
C290 VP.n87 B 0.035687f
C291 VP.n88 B 0.018812f
C292 VP.n89 B 0.039042f
C293 VP.n90 B 0.019645f
C294 VP.n91 B 0.019645f
C295 VP.n92 B 0.019645f
C296 VP.n93 B 0.019884f
C297 VP.n94 B 0.762156f
C298 VP.n95 B 0.03499f
C299 VP.n96 B 0.036429f
C300 VP.n97 B 0.019645f
C301 VP.n98 B 0.019645f
C302 VP.n99 B 0.019645f
C303 VP.n100 B 0.032089f
C304 VP.n101 B 0.036429f
C305 VP.n102 B 0.030314f
C306 VP.n103 B 0.031701f
C307 VP.n104 B 0.043701f
.ends

