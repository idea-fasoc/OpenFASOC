* NGSPICE file created from diff_pair_sample_0249.ext - technology: sky130A

.subckt diff_pair_sample_0249 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=0.4488 pd=3.05 as=1.0608 ps=6.22 w=2.72 l=2.5
X1 B.t11 B.t9 B.t10 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0 ps=0 w=2.72 l=2.5
X2 VDD2.t3 VN.t0 VTAIL.t3 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=0.4488 pd=3.05 as=1.0608 ps=6.22 w=2.72 l=2.5
X3 VTAIL.t0 VN.t1 VDD2.t2 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0.4488 ps=3.05 w=2.72 l=2.5
X4 B.t8 B.t6 B.t7 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0 ps=0 w=2.72 l=2.5
X5 VDD1.t2 VP.t1 VTAIL.t7 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=0.4488 pd=3.05 as=1.0608 ps=6.22 w=2.72 l=2.5
X6 VTAIL.t1 VN.t2 VDD2.t1 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0.4488 ps=3.05 w=2.72 l=2.5
X7 VTAIL.t6 VP.t2 VDD1.t1 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0.4488 ps=3.05 w=2.72 l=2.5
X8 VTAIL.t5 VP.t3 VDD1.t0 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0.4488 ps=3.05 w=2.72 l=2.5
X9 VDD2.t0 VN.t3 VTAIL.t2 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=0.4488 pd=3.05 as=1.0608 ps=6.22 w=2.72 l=2.5
X10 B.t5 B.t3 B.t4 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0 ps=0 w=2.72 l=2.5
X11 B.t2 B.t0 B.t1 w_n2668_n1512# sky130_fd_pr__pfet_01v8 ad=1.0608 pd=6.22 as=0 ps=0 w=2.72 l=2.5
R0 VP.n14 VP.n0 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n11 VP.n1 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n8 VP.n2 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n5 VP.n3 102.573
R7 VP.n16 VP.n15 102.573
R8 VP.n4 VP.t3 61.5696
R9 VP.n4 VP.t0 60.8129
R10 VP.n9 VP.n1 56.4773
R11 VP.n5 VP.n4 43.4643
R12 VP.n3 VP.t2 26.2213
R13 VP.n15 VP.t1 26.2213
R14 VP.n8 VP.n7 24.3439
R15 VP.n9 VP.n8 24.3439
R16 VP.n13 VP.n1 24.3439
R17 VP.n14 VP.n13 24.3439
R18 VP.n7 VP.n3 8.03383
R19 VP.n15 VP.n14 8.03383
R20 VP.n6 VP.n5 0.278398
R21 VP.n16 VP.n0 0.278398
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153422
R28 VTAIL.n5 VTAIL.t5 132.566
R29 VTAIL.n4 VTAIL.t3 132.566
R30 VTAIL.n3 VTAIL.t1 132.566
R31 VTAIL.n7 VTAIL.t2 132.565
R32 VTAIL.n0 VTAIL.t0 132.565
R33 VTAIL.n1 VTAIL.t7 132.565
R34 VTAIL.n2 VTAIL.t6 132.565
R35 VTAIL.n6 VTAIL.t4 132.565
R36 VTAIL.n7 VTAIL.n6 17.1514
R37 VTAIL.n3 VTAIL.n2 17.1514
R38 VTAIL.n4 VTAIL.n3 2.44016
R39 VTAIL.n6 VTAIL.n5 2.44016
R40 VTAIL.n2 VTAIL.n1 2.44016
R41 VTAIL VTAIL.n0 1.27852
R42 VTAIL VTAIL.n7 1.16214
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 VDD1 VDD1.n1 171.197
R46 VDD1 VDD1.n0 137.352
R47 VDD1.n0 VDD1.t0 11.9509
R48 VDD1.n0 VDD1.t3 11.9509
R49 VDD1.n1 VDD1.t1 11.9509
R50 VDD1.n1 VDD1.t2 11.9509
R51 B.n323 B.n42 585
R52 B.n325 B.n324 585
R53 B.n326 B.n41 585
R54 B.n328 B.n327 585
R55 B.n329 B.n40 585
R56 B.n331 B.n330 585
R57 B.n332 B.n39 585
R58 B.n334 B.n333 585
R59 B.n335 B.n38 585
R60 B.n337 B.n336 585
R61 B.n338 B.n37 585
R62 B.n340 B.n339 585
R63 B.n341 B.n33 585
R64 B.n343 B.n342 585
R65 B.n344 B.n32 585
R66 B.n346 B.n345 585
R67 B.n347 B.n31 585
R68 B.n349 B.n348 585
R69 B.n350 B.n30 585
R70 B.n352 B.n351 585
R71 B.n353 B.n29 585
R72 B.n355 B.n354 585
R73 B.n356 B.n28 585
R74 B.n358 B.n357 585
R75 B.n360 B.n25 585
R76 B.n362 B.n361 585
R77 B.n363 B.n24 585
R78 B.n365 B.n364 585
R79 B.n366 B.n23 585
R80 B.n368 B.n367 585
R81 B.n369 B.n22 585
R82 B.n371 B.n370 585
R83 B.n372 B.n21 585
R84 B.n374 B.n373 585
R85 B.n375 B.n20 585
R86 B.n377 B.n376 585
R87 B.n378 B.n19 585
R88 B.n380 B.n379 585
R89 B.n322 B.n321 585
R90 B.n320 B.n43 585
R91 B.n319 B.n318 585
R92 B.n317 B.n44 585
R93 B.n316 B.n315 585
R94 B.n314 B.n45 585
R95 B.n313 B.n312 585
R96 B.n311 B.n46 585
R97 B.n310 B.n309 585
R98 B.n308 B.n47 585
R99 B.n307 B.n306 585
R100 B.n305 B.n48 585
R101 B.n304 B.n303 585
R102 B.n302 B.n49 585
R103 B.n301 B.n300 585
R104 B.n299 B.n50 585
R105 B.n298 B.n297 585
R106 B.n296 B.n51 585
R107 B.n295 B.n294 585
R108 B.n293 B.n52 585
R109 B.n292 B.n291 585
R110 B.n290 B.n53 585
R111 B.n289 B.n288 585
R112 B.n287 B.n54 585
R113 B.n286 B.n285 585
R114 B.n284 B.n55 585
R115 B.n283 B.n282 585
R116 B.n281 B.n56 585
R117 B.n280 B.n279 585
R118 B.n278 B.n57 585
R119 B.n277 B.n276 585
R120 B.n275 B.n58 585
R121 B.n274 B.n273 585
R122 B.n272 B.n59 585
R123 B.n271 B.n270 585
R124 B.n269 B.n60 585
R125 B.n268 B.n267 585
R126 B.n266 B.n61 585
R127 B.n265 B.n264 585
R128 B.n263 B.n62 585
R129 B.n262 B.n261 585
R130 B.n260 B.n63 585
R131 B.n259 B.n258 585
R132 B.n257 B.n64 585
R133 B.n256 B.n255 585
R134 B.n254 B.n65 585
R135 B.n253 B.n252 585
R136 B.n251 B.n66 585
R137 B.n250 B.n249 585
R138 B.n248 B.n67 585
R139 B.n247 B.n246 585
R140 B.n245 B.n68 585
R141 B.n244 B.n243 585
R142 B.n242 B.n69 585
R143 B.n241 B.n240 585
R144 B.n239 B.n70 585
R145 B.n238 B.n237 585
R146 B.n236 B.n71 585
R147 B.n235 B.n234 585
R148 B.n233 B.n72 585
R149 B.n232 B.n231 585
R150 B.n230 B.n73 585
R151 B.n229 B.n228 585
R152 B.n227 B.n74 585
R153 B.n226 B.n225 585
R154 B.n224 B.n75 585
R155 B.n223 B.n222 585
R156 B.n164 B.n99 585
R157 B.n166 B.n165 585
R158 B.n167 B.n98 585
R159 B.n169 B.n168 585
R160 B.n170 B.n97 585
R161 B.n172 B.n171 585
R162 B.n173 B.n96 585
R163 B.n175 B.n174 585
R164 B.n176 B.n95 585
R165 B.n178 B.n177 585
R166 B.n179 B.n94 585
R167 B.n181 B.n180 585
R168 B.n182 B.n93 585
R169 B.n184 B.n183 585
R170 B.n186 B.n90 585
R171 B.n188 B.n187 585
R172 B.n189 B.n89 585
R173 B.n191 B.n190 585
R174 B.n192 B.n88 585
R175 B.n194 B.n193 585
R176 B.n195 B.n87 585
R177 B.n197 B.n196 585
R178 B.n198 B.n86 585
R179 B.n200 B.n199 585
R180 B.n202 B.n201 585
R181 B.n203 B.n82 585
R182 B.n205 B.n204 585
R183 B.n206 B.n81 585
R184 B.n208 B.n207 585
R185 B.n209 B.n80 585
R186 B.n211 B.n210 585
R187 B.n212 B.n79 585
R188 B.n214 B.n213 585
R189 B.n215 B.n78 585
R190 B.n217 B.n216 585
R191 B.n218 B.n77 585
R192 B.n220 B.n219 585
R193 B.n221 B.n76 585
R194 B.n163 B.n162 585
R195 B.n161 B.n100 585
R196 B.n160 B.n159 585
R197 B.n158 B.n101 585
R198 B.n157 B.n156 585
R199 B.n155 B.n102 585
R200 B.n154 B.n153 585
R201 B.n152 B.n103 585
R202 B.n151 B.n150 585
R203 B.n149 B.n104 585
R204 B.n148 B.n147 585
R205 B.n146 B.n105 585
R206 B.n145 B.n144 585
R207 B.n143 B.n106 585
R208 B.n142 B.n141 585
R209 B.n140 B.n107 585
R210 B.n139 B.n138 585
R211 B.n137 B.n108 585
R212 B.n136 B.n135 585
R213 B.n134 B.n109 585
R214 B.n133 B.n132 585
R215 B.n131 B.n110 585
R216 B.n130 B.n129 585
R217 B.n128 B.n111 585
R218 B.n127 B.n126 585
R219 B.n125 B.n112 585
R220 B.n124 B.n123 585
R221 B.n122 B.n113 585
R222 B.n121 B.n120 585
R223 B.n119 B.n114 585
R224 B.n118 B.n117 585
R225 B.n116 B.n115 585
R226 B.n2 B.n0 585
R227 B.n429 B.n1 585
R228 B.n428 B.n427 585
R229 B.n426 B.n3 585
R230 B.n425 B.n424 585
R231 B.n423 B.n4 585
R232 B.n422 B.n421 585
R233 B.n420 B.n5 585
R234 B.n419 B.n418 585
R235 B.n417 B.n6 585
R236 B.n416 B.n415 585
R237 B.n414 B.n7 585
R238 B.n413 B.n412 585
R239 B.n411 B.n8 585
R240 B.n410 B.n409 585
R241 B.n408 B.n9 585
R242 B.n407 B.n406 585
R243 B.n405 B.n10 585
R244 B.n404 B.n403 585
R245 B.n402 B.n11 585
R246 B.n401 B.n400 585
R247 B.n399 B.n12 585
R248 B.n398 B.n397 585
R249 B.n396 B.n13 585
R250 B.n395 B.n394 585
R251 B.n393 B.n14 585
R252 B.n392 B.n391 585
R253 B.n390 B.n15 585
R254 B.n389 B.n388 585
R255 B.n387 B.n16 585
R256 B.n386 B.n385 585
R257 B.n384 B.n17 585
R258 B.n383 B.n382 585
R259 B.n381 B.n18 585
R260 B.n431 B.n430 585
R261 B.n164 B.n163 530.939
R262 B.n381 B.n380 530.939
R263 B.n223 B.n76 530.939
R264 B.n321 B.n42 530.939
R265 B.n83 B.t3 234.112
R266 B.n91 B.t9 234.112
R267 B.n26 B.t6 234.112
R268 B.n34 B.t0 234.112
R269 B.n83 B.t5 195.792
R270 B.n34 B.t1 195.792
R271 B.n91 B.t11 195.792
R272 B.n26 B.t7 195.792
R273 B.n163 B.n100 163.367
R274 B.n159 B.n100 163.367
R275 B.n159 B.n158 163.367
R276 B.n158 B.n157 163.367
R277 B.n157 B.n102 163.367
R278 B.n153 B.n102 163.367
R279 B.n153 B.n152 163.367
R280 B.n152 B.n151 163.367
R281 B.n151 B.n104 163.367
R282 B.n147 B.n104 163.367
R283 B.n147 B.n146 163.367
R284 B.n146 B.n145 163.367
R285 B.n145 B.n106 163.367
R286 B.n141 B.n106 163.367
R287 B.n141 B.n140 163.367
R288 B.n140 B.n139 163.367
R289 B.n139 B.n108 163.367
R290 B.n135 B.n108 163.367
R291 B.n135 B.n134 163.367
R292 B.n134 B.n133 163.367
R293 B.n133 B.n110 163.367
R294 B.n129 B.n110 163.367
R295 B.n129 B.n128 163.367
R296 B.n128 B.n127 163.367
R297 B.n127 B.n112 163.367
R298 B.n123 B.n112 163.367
R299 B.n123 B.n122 163.367
R300 B.n122 B.n121 163.367
R301 B.n121 B.n114 163.367
R302 B.n117 B.n114 163.367
R303 B.n117 B.n116 163.367
R304 B.n116 B.n2 163.367
R305 B.n430 B.n2 163.367
R306 B.n430 B.n429 163.367
R307 B.n429 B.n428 163.367
R308 B.n428 B.n3 163.367
R309 B.n424 B.n3 163.367
R310 B.n424 B.n423 163.367
R311 B.n423 B.n422 163.367
R312 B.n422 B.n5 163.367
R313 B.n418 B.n5 163.367
R314 B.n418 B.n417 163.367
R315 B.n417 B.n416 163.367
R316 B.n416 B.n7 163.367
R317 B.n412 B.n7 163.367
R318 B.n412 B.n411 163.367
R319 B.n411 B.n410 163.367
R320 B.n410 B.n9 163.367
R321 B.n406 B.n9 163.367
R322 B.n406 B.n405 163.367
R323 B.n405 B.n404 163.367
R324 B.n404 B.n11 163.367
R325 B.n400 B.n11 163.367
R326 B.n400 B.n399 163.367
R327 B.n399 B.n398 163.367
R328 B.n398 B.n13 163.367
R329 B.n394 B.n13 163.367
R330 B.n394 B.n393 163.367
R331 B.n393 B.n392 163.367
R332 B.n392 B.n15 163.367
R333 B.n388 B.n15 163.367
R334 B.n388 B.n387 163.367
R335 B.n387 B.n386 163.367
R336 B.n386 B.n17 163.367
R337 B.n382 B.n17 163.367
R338 B.n382 B.n381 163.367
R339 B.n165 B.n164 163.367
R340 B.n165 B.n98 163.367
R341 B.n169 B.n98 163.367
R342 B.n170 B.n169 163.367
R343 B.n171 B.n170 163.367
R344 B.n171 B.n96 163.367
R345 B.n175 B.n96 163.367
R346 B.n176 B.n175 163.367
R347 B.n177 B.n176 163.367
R348 B.n177 B.n94 163.367
R349 B.n181 B.n94 163.367
R350 B.n182 B.n181 163.367
R351 B.n183 B.n182 163.367
R352 B.n183 B.n90 163.367
R353 B.n188 B.n90 163.367
R354 B.n189 B.n188 163.367
R355 B.n190 B.n189 163.367
R356 B.n190 B.n88 163.367
R357 B.n194 B.n88 163.367
R358 B.n195 B.n194 163.367
R359 B.n196 B.n195 163.367
R360 B.n196 B.n86 163.367
R361 B.n200 B.n86 163.367
R362 B.n201 B.n200 163.367
R363 B.n201 B.n82 163.367
R364 B.n205 B.n82 163.367
R365 B.n206 B.n205 163.367
R366 B.n207 B.n206 163.367
R367 B.n207 B.n80 163.367
R368 B.n211 B.n80 163.367
R369 B.n212 B.n211 163.367
R370 B.n213 B.n212 163.367
R371 B.n213 B.n78 163.367
R372 B.n217 B.n78 163.367
R373 B.n218 B.n217 163.367
R374 B.n219 B.n218 163.367
R375 B.n219 B.n76 163.367
R376 B.n224 B.n223 163.367
R377 B.n225 B.n224 163.367
R378 B.n225 B.n74 163.367
R379 B.n229 B.n74 163.367
R380 B.n230 B.n229 163.367
R381 B.n231 B.n230 163.367
R382 B.n231 B.n72 163.367
R383 B.n235 B.n72 163.367
R384 B.n236 B.n235 163.367
R385 B.n237 B.n236 163.367
R386 B.n237 B.n70 163.367
R387 B.n241 B.n70 163.367
R388 B.n242 B.n241 163.367
R389 B.n243 B.n242 163.367
R390 B.n243 B.n68 163.367
R391 B.n247 B.n68 163.367
R392 B.n248 B.n247 163.367
R393 B.n249 B.n248 163.367
R394 B.n249 B.n66 163.367
R395 B.n253 B.n66 163.367
R396 B.n254 B.n253 163.367
R397 B.n255 B.n254 163.367
R398 B.n255 B.n64 163.367
R399 B.n259 B.n64 163.367
R400 B.n260 B.n259 163.367
R401 B.n261 B.n260 163.367
R402 B.n261 B.n62 163.367
R403 B.n265 B.n62 163.367
R404 B.n266 B.n265 163.367
R405 B.n267 B.n266 163.367
R406 B.n267 B.n60 163.367
R407 B.n271 B.n60 163.367
R408 B.n272 B.n271 163.367
R409 B.n273 B.n272 163.367
R410 B.n273 B.n58 163.367
R411 B.n277 B.n58 163.367
R412 B.n278 B.n277 163.367
R413 B.n279 B.n278 163.367
R414 B.n279 B.n56 163.367
R415 B.n283 B.n56 163.367
R416 B.n284 B.n283 163.367
R417 B.n285 B.n284 163.367
R418 B.n285 B.n54 163.367
R419 B.n289 B.n54 163.367
R420 B.n290 B.n289 163.367
R421 B.n291 B.n290 163.367
R422 B.n291 B.n52 163.367
R423 B.n295 B.n52 163.367
R424 B.n296 B.n295 163.367
R425 B.n297 B.n296 163.367
R426 B.n297 B.n50 163.367
R427 B.n301 B.n50 163.367
R428 B.n302 B.n301 163.367
R429 B.n303 B.n302 163.367
R430 B.n303 B.n48 163.367
R431 B.n307 B.n48 163.367
R432 B.n308 B.n307 163.367
R433 B.n309 B.n308 163.367
R434 B.n309 B.n46 163.367
R435 B.n313 B.n46 163.367
R436 B.n314 B.n313 163.367
R437 B.n315 B.n314 163.367
R438 B.n315 B.n44 163.367
R439 B.n319 B.n44 163.367
R440 B.n320 B.n319 163.367
R441 B.n321 B.n320 163.367
R442 B.n380 B.n19 163.367
R443 B.n376 B.n19 163.367
R444 B.n376 B.n375 163.367
R445 B.n375 B.n374 163.367
R446 B.n374 B.n21 163.367
R447 B.n370 B.n21 163.367
R448 B.n370 B.n369 163.367
R449 B.n369 B.n368 163.367
R450 B.n368 B.n23 163.367
R451 B.n364 B.n23 163.367
R452 B.n364 B.n363 163.367
R453 B.n363 B.n362 163.367
R454 B.n362 B.n25 163.367
R455 B.n357 B.n25 163.367
R456 B.n357 B.n356 163.367
R457 B.n356 B.n355 163.367
R458 B.n355 B.n29 163.367
R459 B.n351 B.n29 163.367
R460 B.n351 B.n350 163.367
R461 B.n350 B.n349 163.367
R462 B.n349 B.n31 163.367
R463 B.n345 B.n31 163.367
R464 B.n345 B.n344 163.367
R465 B.n344 B.n343 163.367
R466 B.n343 B.n33 163.367
R467 B.n339 B.n33 163.367
R468 B.n339 B.n338 163.367
R469 B.n338 B.n337 163.367
R470 B.n337 B.n38 163.367
R471 B.n333 B.n38 163.367
R472 B.n333 B.n332 163.367
R473 B.n332 B.n331 163.367
R474 B.n331 B.n40 163.367
R475 B.n327 B.n40 163.367
R476 B.n327 B.n326 163.367
R477 B.n326 B.n325 163.367
R478 B.n325 B.n42 163.367
R479 B.n84 B.t4 140.907
R480 B.n35 B.t2 140.907
R481 B.n92 B.t10 140.906
R482 B.n27 B.t8 140.906
R483 B.n85 B.n84 59.5399
R484 B.n185 B.n92 59.5399
R485 B.n359 B.n27 59.5399
R486 B.n36 B.n35 59.5399
R487 B.n84 B.n83 54.8853
R488 B.n92 B.n91 54.8853
R489 B.n27 B.n26 54.8853
R490 B.n35 B.n34 54.8853
R491 B.n379 B.n18 34.4981
R492 B.n323 B.n322 34.4981
R493 B.n222 B.n221 34.4981
R494 B.n162 B.n99 34.4981
R495 B B.n431 18.0485
R496 B.n379 B.n378 10.6151
R497 B.n378 B.n377 10.6151
R498 B.n377 B.n20 10.6151
R499 B.n373 B.n20 10.6151
R500 B.n373 B.n372 10.6151
R501 B.n372 B.n371 10.6151
R502 B.n371 B.n22 10.6151
R503 B.n367 B.n22 10.6151
R504 B.n367 B.n366 10.6151
R505 B.n366 B.n365 10.6151
R506 B.n365 B.n24 10.6151
R507 B.n361 B.n24 10.6151
R508 B.n361 B.n360 10.6151
R509 B.n358 B.n28 10.6151
R510 B.n354 B.n28 10.6151
R511 B.n354 B.n353 10.6151
R512 B.n353 B.n352 10.6151
R513 B.n352 B.n30 10.6151
R514 B.n348 B.n30 10.6151
R515 B.n348 B.n347 10.6151
R516 B.n347 B.n346 10.6151
R517 B.n346 B.n32 10.6151
R518 B.n342 B.n341 10.6151
R519 B.n341 B.n340 10.6151
R520 B.n340 B.n37 10.6151
R521 B.n336 B.n37 10.6151
R522 B.n336 B.n335 10.6151
R523 B.n335 B.n334 10.6151
R524 B.n334 B.n39 10.6151
R525 B.n330 B.n39 10.6151
R526 B.n330 B.n329 10.6151
R527 B.n329 B.n328 10.6151
R528 B.n328 B.n41 10.6151
R529 B.n324 B.n41 10.6151
R530 B.n324 B.n323 10.6151
R531 B.n222 B.n75 10.6151
R532 B.n226 B.n75 10.6151
R533 B.n227 B.n226 10.6151
R534 B.n228 B.n227 10.6151
R535 B.n228 B.n73 10.6151
R536 B.n232 B.n73 10.6151
R537 B.n233 B.n232 10.6151
R538 B.n234 B.n233 10.6151
R539 B.n234 B.n71 10.6151
R540 B.n238 B.n71 10.6151
R541 B.n239 B.n238 10.6151
R542 B.n240 B.n239 10.6151
R543 B.n240 B.n69 10.6151
R544 B.n244 B.n69 10.6151
R545 B.n245 B.n244 10.6151
R546 B.n246 B.n245 10.6151
R547 B.n246 B.n67 10.6151
R548 B.n250 B.n67 10.6151
R549 B.n251 B.n250 10.6151
R550 B.n252 B.n251 10.6151
R551 B.n252 B.n65 10.6151
R552 B.n256 B.n65 10.6151
R553 B.n257 B.n256 10.6151
R554 B.n258 B.n257 10.6151
R555 B.n258 B.n63 10.6151
R556 B.n262 B.n63 10.6151
R557 B.n263 B.n262 10.6151
R558 B.n264 B.n263 10.6151
R559 B.n264 B.n61 10.6151
R560 B.n268 B.n61 10.6151
R561 B.n269 B.n268 10.6151
R562 B.n270 B.n269 10.6151
R563 B.n270 B.n59 10.6151
R564 B.n274 B.n59 10.6151
R565 B.n275 B.n274 10.6151
R566 B.n276 B.n275 10.6151
R567 B.n276 B.n57 10.6151
R568 B.n280 B.n57 10.6151
R569 B.n281 B.n280 10.6151
R570 B.n282 B.n281 10.6151
R571 B.n282 B.n55 10.6151
R572 B.n286 B.n55 10.6151
R573 B.n287 B.n286 10.6151
R574 B.n288 B.n287 10.6151
R575 B.n288 B.n53 10.6151
R576 B.n292 B.n53 10.6151
R577 B.n293 B.n292 10.6151
R578 B.n294 B.n293 10.6151
R579 B.n294 B.n51 10.6151
R580 B.n298 B.n51 10.6151
R581 B.n299 B.n298 10.6151
R582 B.n300 B.n299 10.6151
R583 B.n300 B.n49 10.6151
R584 B.n304 B.n49 10.6151
R585 B.n305 B.n304 10.6151
R586 B.n306 B.n305 10.6151
R587 B.n306 B.n47 10.6151
R588 B.n310 B.n47 10.6151
R589 B.n311 B.n310 10.6151
R590 B.n312 B.n311 10.6151
R591 B.n312 B.n45 10.6151
R592 B.n316 B.n45 10.6151
R593 B.n317 B.n316 10.6151
R594 B.n318 B.n317 10.6151
R595 B.n318 B.n43 10.6151
R596 B.n322 B.n43 10.6151
R597 B.n166 B.n99 10.6151
R598 B.n167 B.n166 10.6151
R599 B.n168 B.n167 10.6151
R600 B.n168 B.n97 10.6151
R601 B.n172 B.n97 10.6151
R602 B.n173 B.n172 10.6151
R603 B.n174 B.n173 10.6151
R604 B.n174 B.n95 10.6151
R605 B.n178 B.n95 10.6151
R606 B.n179 B.n178 10.6151
R607 B.n180 B.n179 10.6151
R608 B.n180 B.n93 10.6151
R609 B.n184 B.n93 10.6151
R610 B.n187 B.n186 10.6151
R611 B.n187 B.n89 10.6151
R612 B.n191 B.n89 10.6151
R613 B.n192 B.n191 10.6151
R614 B.n193 B.n192 10.6151
R615 B.n193 B.n87 10.6151
R616 B.n197 B.n87 10.6151
R617 B.n198 B.n197 10.6151
R618 B.n199 B.n198 10.6151
R619 B.n203 B.n202 10.6151
R620 B.n204 B.n203 10.6151
R621 B.n204 B.n81 10.6151
R622 B.n208 B.n81 10.6151
R623 B.n209 B.n208 10.6151
R624 B.n210 B.n209 10.6151
R625 B.n210 B.n79 10.6151
R626 B.n214 B.n79 10.6151
R627 B.n215 B.n214 10.6151
R628 B.n216 B.n215 10.6151
R629 B.n216 B.n77 10.6151
R630 B.n220 B.n77 10.6151
R631 B.n221 B.n220 10.6151
R632 B.n162 B.n161 10.6151
R633 B.n161 B.n160 10.6151
R634 B.n160 B.n101 10.6151
R635 B.n156 B.n101 10.6151
R636 B.n156 B.n155 10.6151
R637 B.n155 B.n154 10.6151
R638 B.n154 B.n103 10.6151
R639 B.n150 B.n103 10.6151
R640 B.n150 B.n149 10.6151
R641 B.n149 B.n148 10.6151
R642 B.n148 B.n105 10.6151
R643 B.n144 B.n105 10.6151
R644 B.n144 B.n143 10.6151
R645 B.n143 B.n142 10.6151
R646 B.n142 B.n107 10.6151
R647 B.n138 B.n107 10.6151
R648 B.n138 B.n137 10.6151
R649 B.n137 B.n136 10.6151
R650 B.n136 B.n109 10.6151
R651 B.n132 B.n109 10.6151
R652 B.n132 B.n131 10.6151
R653 B.n131 B.n130 10.6151
R654 B.n130 B.n111 10.6151
R655 B.n126 B.n111 10.6151
R656 B.n126 B.n125 10.6151
R657 B.n125 B.n124 10.6151
R658 B.n124 B.n113 10.6151
R659 B.n120 B.n113 10.6151
R660 B.n120 B.n119 10.6151
R661 B.n119 B.n118 10.6151
R662 B.n118 B.n115 10.6151
R663 B.n115 B.n0 10.6151
R664 B.n427 B.n1 10.6151
R665 B.n427 B.n426 10.6151
R666 B.n426 B.n425 10.6151
R667 B.n425 B.n4 10.6151
R668 B.n421 B.n4 10.6151
R669 B.n421 B.n420 10.6151
R670 B.n420 B.n419 10.6151
R671 B.n419 B.n6 10.6151
R672 B.n415 B.n6 10.6151
R673 B.n415 B.n414 10.6151
R674 B.n414 B.n413 10.6151
R675 B.n413 B.n8 10.6151
R676 B.n409 B.n8 10.6151
R677 B.n409 B.n408 10.6151
R678 B.n408 B.n407 10.6151
R679 B.n407 B.n10 10.6151
R680 B.n403 B.n10 10.6151
R681 B.n403 B.n402 10.6151
R682 B.n402 B.n401 10.6151
R683 B.n401 B.n12 10.6151
R684 B.n397 B.n12 10.6151
R685 B.n397 B.n396 10.6151
R686 B.n396 B.n395 10.6151
R687 B.n395 B.n14 10.6151
R688 B.n391 B.n14 10.6151
R689 B.n391 B.n390 10.6151
R690 B.n390 B.n389 10.6151
R691 B.n389 B.n16 10.6151
R692 B.n385 B.n16 10.6151
R693 B.n385 B.n384 10.6151
R694 B.n384 B.n383 10.6151
R695 B.n383 B.n18 10.6151
R696 B.n360 B.n359 9.36635
R697 B.n342 B.n36 9.36635
R698 B.n185 B.n184 9.36635
R699 B.n202 B.n85 9.36635
R700 B.n431 B.n0 2.81026
R701 B.n431 B.n1 2.81026
R702 B.n359 B.n358 1.24928
R703 B.n36 B.n32 1.24928
R704 B.n186 B.n185 1.24928
R705 B.n199 B.n85 1.24928
R706 VN.n0 VN.t1 61.5696
R707 VN.n1 VN.t0 61.5696
R708 VN.n0 VN.t3 60.8129
R709 VN.n1 VN.t2 60.8129
R710 VN VN.n1 43.7432
R711 VN VN.n0 4.54245
R712 VDD2.n2 VDD2.n0 170.673
R713 VDD2.n2 VDD2.n1 137.294
R714 VDD2.n1 VDD2.t1 11.9509
R715 VDD2.n1 VDD2.t3 11.9509
R716 VDD2.n0 VDD2.t2 11.9509
R717 VDD2.n0 VDD2.t0 11.9509
R718 VDD2 VDD2.n2 0.0586897
C0 VN VDD2 1.31487f
C1 VDD2 VDD1 1.00962f
C2 VN VP 4.41255f
C3 VDD2 VTAIL 3.20539f
C4 VDD2 B 1.04295f
C5 VP VDD1 1.55309f
C6 VN VDD1 0.153816f
C7 VP VTAIL 1.80677f
C8 VP B 1.53408f
C9 VN VTAIL 1.79267f
C10 VN B 0.9663f
C11 VTAIL VDD1 3.15185f
C12 B VDD1 0.992244f
C13 B VTAIL 1.80611f
C14 w_n2668_n1512# VDD2 1.23788f
C15 w_n2668_n1512# VP 4.66399f
C16 w_n2668_n1512# VN 4.32406f
C17 w_n2668_n1512# VDD1 1.18452f
C18 w_n2668_n1512# VTAIL 1.84642f
C19 w_n2668_n1512# B 6.54472f
C20 VP VDD2 0.393527f
C21 VDD2 VSUBS 0.637434f
C22 VDD1 VSUBS 3.269874f
C23 VTAIL VSUBS 0.439114f
C24 VN VSUBS 4.77966f
C25 VP VSUBS 1.71824f
C26 B VSUBS 3.218826f
C27 w_n2668_n1512# VSUBS 51.1936f
C28 VDD2.t2 VSUBS 0.04335f
C29 VDD2.t0 VSUBS 0.04335f
C30 VDD2.n0 VSUBS 0.39192f
C31 VDD2.t1 VSUBS 0.04335f
C32 VDD2.t3 VSUBS 0.04335f
C33 VDD2.n1 VSUBS 0.220796f
C34 VDD2.n2 VSUBS 2.251f
C35 VN.t1 VSUBS 0.95379f
C36 VN.t3 VSUBS 0.947357f
C37 VN.n0 VSUBS 0.607477f
C38 VN.t0 VSUBS 0.95379f
C39 VN.t2 VSUBS 0.947357f
C40 VN.n1 VSUBS 2.24172f
C41 B.n0 VSUBS 0.005119f
C42 B.n1 VSUBS 0.005119f
C43 B.n2 VSUBS 0.008096f
C44 B.n3 VSUBS 0.008096f
C45 B.n4 VSUBS 0.008096f
C46 B.n5 VSUBS 0.008096f
C47 B.n6 VSUBS 0.008096f
C48 B.n7 VSUBS 0.008096f
C49 B.n8 VSUBS 0.008096f
C50 B.n9 VSUBS 0.008096f
C51 B.n10 VSUBS 0.008096f
C52 B.n11 VSUBS 0.008096f
C53 B.n12 VSUBS 0.008096f
C54 B.n13 VSUBS 0.008096f
C55 B.n14 VSUBS 0.008096f
C56 B.n15 VSUBS 0.008096f
C57 B.n16 VSUBS 0.008096f
C58 B.n17 VSUBS 0.008096f
C59 B.n18 VSUBS 0.019236f
C60 B.n19 VSUBS 0.008096f
C61 B.n20 VSUBS 0.008096f
C62 B.n21 VSUBS 0.008096f
C63 B.n22 VSUBS 0.008096f
C64 B.n23 VSUBS 0.008096f
C65 B.n24 VSUBS 0.008096f
C66 B.n25 VSUBS 0.008096f
C67 B.t8 VSUBS 0.073925f
C68 B.t7 VSUBS 0.091116f
C69 B.t6 VSUBS 0.383307f
C70 B.n26 VSUBS 0.089187f
C71 B.n27 VSUBS 0.072871f
C72 B.n28 VSUBS 0.008096f
C73 B.n29 VSUBS 0.008096f
C74 B.n30 VSUBS 0.008096f
C75 B.n31 VSUBS 0.008096f
C76 B.n32 VSUBS 0.004524f
C77 B.n33 VSUBS 0.008096f
C78 B.t2 VSUBS 0.073925f
C79 B.t1 VSUBS 0.091116f
C80 B.t0 VSUBS 0.383307f
C81 B.n34 VSUBS 0.089187f
C82 B.n35 VSUBS 0.072871f
C83 B.n36 VSUBS 0.018757f
C84 B.n37 VSUBS 0.008096f
C85 B.n38 VSUBS 0.008096f
C86 B.n39 VSUBS 0.008096f
C87 B.n40 VSUBS 0.008096f
C88 B.n41 VSUBS 0.008096f
C89 B.n42 VSUBS 0.020053f
C90 B.n43 VSUBS 0.008096f
C91 B.n44 VSUBS 0.008096f
C92 B.n45 VSUBS 0.008096f
C93 B.n46 VSUBS 0.008096f
C94 B.n47 VSUBS 0.008096f
C95 B.n48 VSUBS 0.008096f
C96 B.n49 VSUBS 0.008096f
C97 B.n50 VSUBS 0.008096f
C98 B.n51 VSUBS 0.008096f
C99 B.n52 VSUBS 0.008096f
C100 B.n53 VSUBS 0.008096f
C101 B.n54 VSUBS 0.008096f
C102 B.n55 VSUBS 0.008096f
C103 B.n56 VSUBS 0.008096f
C104 B.n57 VSUBS 0.008096f
C105 B.n58 VSUBS 0.008096f
C106 B.n59 VSUBS 0.008096f
C107 B.n60 VSUBS 0.008096f
C108 B.n61 VSUBS 0.008096f
C109 B.n62 VSUBS 0.008096f
C110 B.n63 VSUBS 0.008096f
C111 B.n64 VSUBS 0.008096f
C112 B.n65 VSUBS 0.008096f
C113 B.n66 VSUBS 0.008096f
C114 B.n67 VSUBS 0.008096f
C115 B.n68 VSUBS 0.008096f
C116 B.n69 VSUBS 0.008096f
C117 B.n70 VSUBS 0.008096f
C118 B.n71 VSUBS 0.008096f
C119 B.n72 VSUBS 0.008096f
C120 B.n73 VSUBS 0.008096f
C121 B.n74 VSUBS 0.008096f
C122 B.n75 VSUBS 0.008096f
C123 B.n76 VSUBS 0.020053f
C124 B.n77 VSUBS 0.008096f
C125 B.n78 VSUBS 0.008096f
C126 B.n79 VSUBS 0.008096f
C127 B.n80 VSUBS 0.008096f
C128 B.n81 VSUBS 0.008096f
C129 B.n82 VSUBS 0.008096f
C130 B.t4 VSUBS 0.073925f
C131 B.t5 VSUBS 0.091116f
C132 B.t3 VSUBS 0.383307f
C133 B.n83 VSUBS 0.089187f
C134 B.n84 VSUBS 0.072871f
C135 B.n85 VSUBS 0.018757f
C136 B.n86 VSUBS 0.008096f
C137 B.n87 VSUBS 0.008096f
C138 B.n88 VSUBS 0.008096f
C139 B.n89 VSUBS 0.008096f
C140 B.n90 VSUBS 0.008096f
C141 B.t10 VSUBS 0.073925f
C142 B.t11 VSUBS 0.091116f
C143 B.t9 VSUBS 0.383307f
C144 B.n91 VSUBS 0.089187f
C145 B.n92 VSUBS 0.072871f
C146 B.n93 VSUBS 0.008096f
C147 B.n94 VSUBS 0.008096f
C148 B.n95 VSUBS 0.008096f
C149 B.n96 VSUBS 0.008096f
C150 B.n97 VSUBS 0.008096f
C151 B.n98 VSUBS 0.008096f
C152 B.n99 VSUBS 0.020053f
C153 B.n100 VSUBS 0.008096f
C154 B.n101 VSUBS 0.008096f
C155 B.n102 VSUBS 0.008096f
C156 B.n103 VSUBS 0.008096f
C157 B.n104 VSUBS 0.008096f
C158 B.n105 VSUBS 0.008096f
C159 B.n106 VSUBS 0.008096f
C160 B.n107 VSUBS 0.008096f
C161 B.n108 VSUBS 0.008096f
C162 B.n109 VSUBS 0.008096f
C163 B.n110 VSUBS 0.008096f
C164 B.n111 VSUBS 0.008096f
C165 B.n112 VSUBS 0.008096f
C166 B.n113 VSUBS 0.008096f
C167 B.n114 VSUBS 0.008096f
C168 B.n115 VSUBS 0.008096f
C169 B.n116 VSUBS 0.008096f
C170 B.n117 VSUBS 0.008096f
C171 B.n118 VSUBS 0.008096f
C172 B.n119 VSUBS 0.008096f
C173 B.n120 VSUBS 0.008096f
C174 B.n121 VSUBS 0.008096f
C175 B.n122 VSUBS 0.008096f
C176 B.n123 VSUBS 0.008096f
C177 B.n124 VSUBS 0.008096f
C178 B.n125 VSUBS 0.008096f
C179 B.n126 VSUBS 0.008096f
C180 B.n127 VSUBS 0.008096f
C181 B.n128 VSUBS 0.008096f
C182 B.n129 VSUBS 0.008096f
C183 B.n130 VSUBS 0.008096f
C184 B.n131 VSUBS 0.008096f
C185 B.n132 VSUBS 0.008096f
C186 B.n133 VSUBS 0.008096f
C187 B.n134 VSUBS 0.008096f
C188 B.n135 VSUBS 0.008096f
C189 B.n136 VSUBS 0.008096f
C190 B.n137 VSUBS 0.008096f
C191 B.n138 VSUBS 0.008096f
C192 B.n139 VSUBS 0.008096f
C193 B.n140 VSUBS 0.008096f
C194 B.n141 VSUBS 0.008096f
C195 B.n142 VSUBS 0.008096f
C196 B.n143 VSUBS 0.008096f
C197 B.n144 VSUBS 0.008096f
C198 B.n145 VSUBS 0.008096f
C199 B.n146 VSUBS 0.008096f
C200 B.n147 VSUBS 0.008096f
C201 B.n148 VSUBS 0.008096f
C202 B.n149 VSUBS 0.008096f
C203 B.n150 VSUBS 0.008096f
C204 B.n151 VSUBS 0.008096f
C205 B.n152 VSUBS 0.008096f
C206 B.n153 VSUBS 0.008096f
C207 B.n154 VSUBS 0.008096f
C208 B.n155 VSUBS 0.008096f
C209 B.n156 VSUBS 0.008096f
C210 B.n157 VSUBS 0.008096f
C211 B.n158 VSUBS 0.008096f
C212 B.n159 VSUBS 0.008096f
C213 B.n160 VSUBS 0.008096f
C214 B.n161 VSUBS 0.008096f
C215 B.n162 VSUBS 0.019236f
C216 B.n163 VSUBS 0.019236f
C217 B.n164 VSUBS 0.020053f
C218 B.n165 VSUBS 0.008096f
C219 B.n166 VSUBS 0.008096f
C220 B.n167 VSUBS 0.008096f
C221 B.n168 VSUBS 0.008096f
C222 B.n169 VSUBS 0.008096f
C223 B.n170 VSUBS 0.008096f
C224 B.n171 VSUBS 0.008096f
C225 B.n172 VSUBS 0.008096f
C226 B.n173 VSUBS 0.008096f
C227 B.n174 VSUBS 0.008096f
C228 B.n175 VSUBS 0.008096f
C229 B.n176 VSUBS 0.008096f
C230 B.n177 VSUBS 0.008096f
C231 B.n178 VSUBS 0.008096f
C232 B.n179 VSUBS 0.008096f
C233 B.n180 VSUBS 0.008096f
C234 B.n181 VSUBS 0.008096f
C235 B.n182 VSUBS 0.008096f
C236 B.n183 VSUBS 0.008096f
C237 B.n184 VSUBS 0.00762f
C238 B.n185 VSUBS 0.018757f
C239 B.n186 VSUBS 0.004524f
C240 B.n187 VSUBS 0.008096f
C241 B.n188 VSUBS 0.008096f
C242 B.n189 VSUBS 0.008096f
C243 B.n190 VSUBS 0.008096f
C244 B.n191 VSUBS 0.008096f
C245 B.n192 VSUBS 0.008096f
C246 B.n193 VSUBS 0.008096f
C247 B.n194 VSUBS 0.008096f
C248 B.n195 VSUBS 0.008096f
C249 B.n196 VSUBS 0.008096f
C250 B.n197 VSUBS 0.008096f
C251 B.n198 VSUBS 0.008096f
C252 B.n199 VSUBS 0.004524f
C253 B.n200 VSUBS 0.008096f
C254 B.n201 VSUBS 0.008096f
C255 B.n202 VSUBS 0.00762f
C256 B.n203 VSUBS 0.008096f
C257 B.n204 VSUBS 0.008096f
C258 B.n205 VSUBS 0.008096f
C259 B.n206 VSUBS 0.008096f
C260 B.n207 VSUBS 0.008096f
C261 B.n208 VSUBS 0.008096f
C262 B.n209 VSUBS 0.008096f
C263 B.n210 VSUBS 0.008096f
C264 B.n211 VSUBS 0.008096f
C265 B.n212 VSUBS 0.008096f
C266 B.n213 VSUBS 0.008096f
C267 B.n214 VSUBS 0.008096f
C268 B.n215 VSUBS 0.008096f
C269 B.n216 VSUBS 0.008096f
C270 B.n217 VSUBS 0.008096f
C271 B.n218 VSUBS 0.008096f
C272 B.n219 VSUBS 0.008096f
C273 B.n220 VSUBS 0.008096f
C274 B.n221 VSUBS 0.020053f
C275 B.n222 VSUBS 0.019236f
C276 B.n223 VSUBS 0.019236f
C277 B.n224 VSUBS 0.008096f
C278 B.n225 VSUBS 0.008096f
C279 B.n226 VSUBS 0.008096f
C280 B.n227 VSUBS 0.008096f
C281 B.n228 VSUBS 0.008096f
C282 B.n229 VSUBS 0.008096f
C283 B.n230 VSUBS 0.008096f
C284 B.n231 VSUBS 0.008096f
C285 B.n232 VSUBS 0.008096f
C286 B.n233 VSUBS 0.008096f
C287 B.n234 VSUBS 0.008096f
C288 B.n235 VSUBS 0.008096f
C289 B.n236 VSUBS 0.008096f
C290 B.n237 VSUBS 0.008096f
C291 B.n238 VSUBS 0.008096f
C292 B.n239 VSUBS 0.008096f
C293 B.n240 VSUBS 0.008096f
C294 B.n241 VSUBS 0.008096f
C295 B.n242 VSUBS 0.008096f
C296 B.n243 VSUBS 0.008096f
C297 B.n244 VSUBS 0.008096f
C298 B.n245 VSUBS 0.008096f
C299 B.n246 VSUBS 0.008096f
C300 B.n247 VSUBS 0.008096f
C301 B.n248 VSUBS 0.008096f
C302 B.n249 VSUBS 0.008096f
C303 B.n250 VSUBS 0.008096f
C304 B.n251 VSUBS 0.008096f
C305 B.n252 VSUBS 0.008096f
C306 B.n253 VSUBS 0.008096f
C307 B.n254 VSUBS 0.008096f
C308 B.n255 VSUBS 0.008096f
C309 B.n256 VSUBS 0.008096f
C310 B.n257 VSUBS 0.008096f
C311 B.n258 VSUBS 0.008096f
C312 B.n259 VSUBS 0.008096f
C313 B.n260 VSUBS 0.008096f
C314 B.n261 VSUBS 0.008096f
C315 B.n262 VSUBS 0.008096f
C316 B.n263 VSUBS 0.008096f
C317 B.n264 VSUBS 0.008096f
C318 B.n265 VSUBS 0.008096f
C319 B.n266 VSUBS 0.008096f
C320 B.n267 VSUBS 0.008096f
C321 B.n268 VSUBS 0.008096f
C322 B.n269 VSUBS 0.008096f
C323 B.n270 VSUBS 0.008096f
C324 B.n271 VSUBS 0.008096f
C325 B.n272 VSUBS 0.008096f
C326 B.n273 VSUBS 0.008096f
C327 B.n274 VSUBS 0.008096f
C328 B.n275 VSUBS 0.008096f
C329 B.n276 VSUBS 0.008096f
C330 B.n277 VSUBS 0.008096f
C331 B.n278 VSUBS 0.008096f
C332 B.n279 VSUBS 0.008096f
C333 B.n280 VSUBS 0.008096f
C334 B.n281 VSUBS 0.008096f
C335 B.n282 VSUBS 0.008096f
C336 B.n283 VSUBS 0.008096f
C337 B.n284 VSUBS 0.008096f
C338 B.n285 VSUBS 0.008096f
C339 B.n286 VSUBS 0.008096f
C340 B.n287 VSUBS 0.008096f
C341 B.n288 VSUBS 0.008096f
C342 B.n289 VSUBS 0.008096f
C343 B.n290 VSUBS 0.008096f
C344 B.n291 VSUBS 0.008096f
C345 B.n292 VSUBS 0.008096f
C346 B.n293 VSUBS 0.008096f
C347 B.n294 VSUBS 0.008096f
C348 B.n295 VSUBS 0.008096f
C349 B.n296 VSUBS 0.008096f
C350 B.n297 VSUBS 0.008096f
C351 B.n298 VSUBS 0.008096f
C352 B.n299 VSUBS 0.008096f
C353 B.n300 VSUBS 0.008096f
C354 B.n301 VSUBS 0.008096f
C355 B.n302 VSUBS 0.008096f
C356 B.n303 VSUBS 0.008096f
C357 B.n304 VSUBS 0.008096f
C358 B.n305 VSUBS 0.008096f
C359 B.n306 VSUBS 0.008096f
C360 B.n307 VSUBS 0.008096f
C361 B.n308 VSUBS 0.008096f
C362 B.n309 VSUBS 0.008096f
C363 B.n310 VSUBS 0.008096f
C364 B.n311 VSUBS 0.008096f
C365 B.n312 VSUBS 0.008096f
C366 B.n313 VSUBS 0.008096f
C367 B.n314 VSUBS 0.008096f
C368 B.n315 VSUBS 0.008096f
C369 B.n316 VSUBS 0.008096f
C370 B.n317 VSUBS 0.008096f
C371 B.n318 VSUBS 0.008096f
C372 B.n319 VSUBS 0.008096f
C373 B.n320 VSUBS 0.008096f
C374 B.n321 VSUBS 0.019236f
C375 B.n322 VSUBS 0.020141f
C376 B.n323 VSUBS 0.019147f
C377 B.n324 VSUBS 0.008096f
C378 B.n325 VSUBS 0.008096f
C379 B.n326 VSUBS 0.008096f
C380 B.n327 VSUBS 0.008096f
C381 B.n328 VSUBS 0.008096f
C382 B.n329 VSUBS 0.008096f
C383 B.n330 VSUBS 0.008096f
C384 B.n331 VSUBS 0.008096f
C385 B.n332 VSUBS 0.008096f
C386 B.n333 VSUBS 0.008096f
C387 B.n334 VSUBS 0.008096f
C388 B.n335 VSUBS 0.008096f
C389 B.n336 VSUBS 0.008096f
C390 B.n337 VSUBS 0.008096f
C391 B.n338 VSUBS 0.008096f
C392 B.n339 VSUBS 0.008096f
C393 B.n340 VSUBS 0.008096f
C394 B.n341 VSUBS 0.008096f
C395 B.n342 VSUBS 0.00762f
C396 B.n343 VSUBS 0.008096f
C397 B.n344 VSUBS 0.008096f
C398 B.n345 VSUBS 0.008096f
C399 B.n346 VSUBS 0.008096f
C400 B.n347 VSUBS 0.008096f
C401 B.n348 VSUBS 0.008096f
C402 B.n349 VSUBS 0.008096f
C403 B.n350 VSUBS 0.008096f
C404 B.n351 VSUBS 0.008096f
C405 B.n352 VSUBS 0.008096f
C406 B.n353 VSUBS 0.008096f
C407 B.n354 VSUBS 0.008096f
C408 B.n355 VSUBS 0.008096f
C409 B.n356 VSUBS 0.008096f
C410 B.n357 VSUBS 0.008096f
C411 B.n358 VSUBS 0.004524f
C412 B.n359 VSUBS 0.018757f
C413 B.n360 VSUBS 0.00762f
C414 B.n361 VSUBS 0.008096f
C415 B.n362 VSUBS 0.008096f
C416 B.n363 VSUBS 0.008096f
C417 B.n364 VSUBS 0.008096f
C418 B.n365 VSUBS 0.008096f
C419 B.n366 VSUBS 0.008096f
C420 B.n367 VSUBS 0.008096f
C421 B.n368 VSUBS 0.008096f
C422 B.n369 VSUBS 0.008096f
C423 B.n370 VSUBS 0.008096f
C424 B.n371 VSUBS 0.008096f
C425 B.n372 VSUBS 0.008096f
C426 B.n373 VSUBS 0.008096f
C427 B.n374 VSUBS 0.008096f
C428 B.n375 VSUBS 0.008096f
C429 B.n376 VSUBS 0.008096f
C430 B.n377 VSUBS 0.008096f
C431 B.n378 VSUBS 0.008096f
C432 B.n379 VSUBS 0.020053f
C433 B.n380 VSUBS 0.020053f
C434 B.n381 VSUBS 0.019236f
C435 B.n382 VSUBS 0.008096f
C436 B.n383 VSUBS 0.008096f
C437 B.n384 VSUBS 0.008096f
C438 B.n385 VSUBS 0.008096f
C439 B.n386 VSUBS 0.008096f
C440 B.n387 VSUBS 0.008096f
C441 B.n388 VSUBS 0.008096f
C442 B.n389 VSUBS 0.008096f
C443 B.n390 VSUBS 0.008096f
C444 B.n391 VSUBS 0.008096f
C445 B.n392 VSUBS 0.008096f
C446 B.n393 VSUBS 0.008096f
C447 B.n394 VSUBS 0.008096f
C448 B.n395 VSUBS 0.008096f
C449 B.n396 VSUBS 0.008096f
C450 B.n397 VSUBS 0.008096f
C451 B.n398 VSUBS 0.008096f
C452 B.n399 VSUBS 0.008096f
C453 B.n400 VSUBS 0.008096f
C454 B.n401 VSUBS 0.008096f
C455 B.n402 VSUBS 0.008096f
C456 B.n403 VSUBS 0.008096f
C457 B.n404 VSUBS 0.008096f
C458 B.n405 VSUBS 0.008096f
C459 B.n406 VSUBS 0.008096f
C460 B.n407 VSUBS 0.008096f
C461 B.n408 VSUBS 0.008096f
C462 B.n409 VSUBS 0.008096f
C463 B.n410 VSUBS 0.008096f
C464 B.n411 VSUBS 0.008096f
C465 B.n412 VSUBS 0.008096f
C466 B.n413 VSUBS 0.008096f
C467 B.n414 VSUBS 0.008096f
C468 B.n415 VSUBS 0.008096f
C469 B.n416 VSUBS 0.008096f
C470 B.n417 VSUBS 0.008096f
C471 B.n418 VSUBS 0.008096f
C472 B.n419 VSUBS 0.008096f
C473 B.n420 VSUBS 0.008096f
C474 B.n421 VSUBS 0.008096f
C475 B.n422 VSUBS 0.008096f
C476 B.n423 VSUBS 0.008096f
C477 B.n424 VSUBS 0.008096f
C478 B.n425 VSUBS 0.008096f
C479 B.n426 VSUBS 0.008096f
C480 B.n427 VSUBS 0.008096f
C481 B.n428 VSUBS 0.008096f
C482 B.n429 VSUBS 0.008096f
C483 B.n430 VSUBS 0.008096f
C484 B.n431 VSUBS 0.018332f
C485 VDD1.t0 VSUBS 0.042364f
C486 VDD1.t3 VSUBS 0.042364f
C487 VDD1.n0 VSUBS 0.215944f
C488 VDD1.t1 VSUBS 0.042364f
C489 VDD1.t2 VSUBS 0.042364f
C490 VDD1.n1 VSUBS 0.393024f
C491 VTAIL.t0 VSUBS 0.221205f
C492 VTAIL.n0 VSUBS 0.302428f
C493 VTAIL.t7 VSUBS 0.221205f
C494 VTAIL.n1 VSUBS 0.361586f
C495 VTAIL.t6 VSUBS 0.221205f
C496 VTAIL.n2 VSUBS 0.796003f
C497 VTAIL.t1 VSUBS 0.221206f
C498 VTAIL.n3 VSUBS 0.796003f
C499 VTAIL.t3 VSUBS 0.221206f
C500 VTAIL.n4 VSUBS 0.361585f
C501 VTAIL.t5 VSUBS 0.221206f
C502 VTAIL.n5 VSUBS 0.361585f
C503 VTAIL.t4 VSUBS 0.221205f
C504 VTAIL.n6 VSUBS 0.796003f
C505 VTAIL.t2 VSUBS 0.221205f
C506 VTAIL.n7 VSUBS 0.730919f
C507 VP.n0 VSUBS 0.053996f
C508 VP.t1 VSUBS 0.6848f
C509 VP.n1 VSUBS 0.060045f
C510 VP.n2 VSUBS 0.040954f
C511 VP.t2 VSUBS 0.6848f
C512 VP.n3 VSUBS 0.426341f
C513 VP.t0 VSUBS 0.997183f
C514 VP.t3 VSUBS 1.00395f
C515 VP.n4 VSUBS 2.33771f
C516 VP.n5 VSUBS 1.77609f
C517 VP.n6 VSUBS 0.053996f
C518 VP.n7 VSUBS 0.051334f
C519 VP.n8 VSUBS 0.07671f
C520 VP.n9 VSUBS 0.060045f
C521 VP.n10 VSUBS 0.040954f
C522 VP.n11 VSUBS 0.040954f
C523 VP.n12 VSUBS 0.040954f
C524 VP.n13 VSUBS 0.07671f
C525 VP.n14 VSUBS 0.051334f
C526 VP.n15 VSUBS 0.426341f
C527 VP.n16 VSUBS 0.067245f
.ends

