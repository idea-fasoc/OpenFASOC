* NGSPICE file created from diff_pair_sample_1675.ext - technology: sky130A

.subckt diff_pair_sample_1675 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0 ps=0 w=0.63 l=0.94
X1 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0 ps=0 w=0.63 l=0.94
X2 VDD1.t5 VP.t0 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.2457 ps=2.04 w=0.63 l=0.94
X3 VTAIL.t9 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.10395 ps=0.96 w=0.63 l=0.94
X4 VDD1.t3 VP.t2 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0.10395 ps=0.96 w=0.63 l=0.94
X5 VTAIL.t1 VN.t0 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.10395 ps=0.96 w=0.63 l=0.94
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0 ps=0 w=0.63 l=0.94
X7 VDD2.t4 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0.10395 ps=0.96 w=0.63 l=0.94
X8 VDD2.t3 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.2457 ps=2.04 w=0.63 l=0.94
X9 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0.10395 ps=0.96 w=0.63 l=0.94
X10 VTAIL.t7 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.10395 ps=0.96 w=0.63 l=0.94
X11 VDD2.t1 VN.t4 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.2457 ps=2.04 w=0.63 l=0.94
X12 VDD1.t1 VP.t4 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.2457 ps=2.04 w=0.63 l=0.94
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0 ps=0 w=0.63 l=0.94
X14 VTAIL.t2 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.10395 pd=0.96 as=0.10395 ps=0.96 w=0.63 l=0.94
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2457 pd=2.04 as=0.10395 ps=0.96 w=0.63 l=0.94
R0 B.n324 B.n323 585
R1 B.n110 B.n58 585
R2 B.n109 B.n108 585
R3 B.n107 B.n106 585
R4 B.n105 B.n104 585
R5 B.n103 B.n102 585
R6 B.n101 B.n100 585
R7 B.n99 B.n98 585
R8 B.n97 B.n96 585
R9 B.n95 B.n94 585
R10 B.n93 B.n92 585
R11 B.n91 B.n90 585
R12 B.n89 B.n88 585
R13 B.n87 B.n86 585
R14 B.n85 B.n84 585
R15 B.n83 B.n82 585
R16 B.n81 B.n80 585
R17 B.n79 B.n78 585
R18 B.n77 B.n76 585
R19 B.n75 B.n74 585
R20 B.n73 B.n72 585
R21 B.n71 B.n70 585
R22 B.n69 B.n68 585
R23 B.n67 B.n66 585
R24 B.n46 B.n45 585
R25 B.n329 B.n328 585
R26 B.n322 B.n59 585
R27 B.n59 B.n43 585
R28 B.n321 B.n42 585
R29 B.n333 B.n42 585
R30 B.n320 B.n41 585
R31 B.n334 B.n41 585
R32 B.n319 B.n40 585
R33 B.n335 B.n40 585
R34 B.n318 B.n317 585
R35 B.n317 B.n36 585
R36 B.n316 B.n35 585
R37 B.n341 B.n35 585
R38 B.n315 B.n34 585
R39 B.n342 B.n34 585
R40 B.n314 B.n33 585
R41 B.n343 B.n33 585
R42 B.n313 B.n312 585
R43 B.n312 B.n29 585
R44 B.n311 B.n28 585
R45 B.n349 B.n28 585
R46 B.n310 B.n27 585
R47 B.n350 B.n27 585
R48 B.n309 B.n26 585
R49 B.n351 B.n26 585
R50 B.n308 B.n307 585
R51 B.n307 B.n25 585
R52 B.n306 B.n21 585
R53 B.n357 B.n21 585
R54 B.n305 B.n20 585
R55 B.n358 B.n20 585
R56 B.n304 B.n19 585
R57 B.n359 B.n19 585
R58 B.n303 B.n302 585
R59 B.n302 B.n15 585
R60 B.n301 B.n14 585
R61 B.n365 B.n14 585
R62 B.n300 B.n13 585
R63 B.n366 B.n13 585
R64 B.n299 B.n12 585
R65 B.n367 B.n12 585
R66 B.n298 B.n297 585
R67 B.n297 B.n8 585
R68 B.n296 B.n7 585
R69 B.n373 B.n7 585
R70 B.n295 B.n6 585
R71 B.n374 B.n6 585
R72 B.n294 B.n5 585
R73 B.n375 B.n5 585
R74 B.n293 B.n292 585
R75 B.n292 B.n4 585
R76 B.n291 B.n111 585
R77 B.n291 B.n290 585
R78 B.n281 B.n112 585
R79 B.n113 B.n112 585
R80 B.n283 B.n282 585
R81 B.n284 B.n283 585
R82 B.n280 B.n118 585
R83 B.n118 B.n117 585
R84 B.n279 B.n278 585
R85 B.n278 B.n277 585
R86 B.n120 B.n119 585
R87 B.n121 B.n120 585
R88 B.n270 B.n269 585
R89 B.n271 B.n270 585
R90 B.n268 B.n126 585
R91 B.n126 B.n125 585
R92 B.n267 B.n266 585
R93 B.n266 B.n265 585
R94 B.n128 B.n127 585
R95 B.n258 B.n128 585
R96 B.n257 B.n256 585
R97 B.n259 B.n257 585
R98 B.n255 B.n133 585
R99 B.n133 B.n132 585
R100 B.n254 B.n253 585
R101 B.n253 B.n252 585
R102 B.n135 B.n134 585
R103 B.n136 B.n135 585
R104 B.n245 B.n244 585
R105 B.n246 B.n245 585
R106 B.n243 B.n141 585
R107 B.n141 B.n140 585
R108 B.n242 B.n241 585
R109 B.n241 B.n240 585
R110 B.n143 B.n142 585
R111 B.n144 B.n143 585
R112 B.n233 B.n232 585
R113 B.n234 B.n233 585
R114 B.n231 B.n149 585
R115 B.n149 B.n148 585
R116 B.n230 B.n229 585
R117 B.n229 B.n228 585
R118 B.n151 B.n150 585
R119 B.n152 B.n151 585
R120 B.n224 B.n223 585
R121 B.n155 B.n154 585
R122 B.n220 B.n219 585
R123 B.n221 B.n220 585
R124 B.n218 B.n168 585
R125 B.n217 B.n216 585
R126 B.n215 B.n214 585
R127 B.n213 B.n212 585
R128 B.n211 B.n210 585
R129 B.n208 B.n207 585
R130 B.n206 B.n205 585
R131 B.n204 B.n203 585
R132 B.n202 B.n201 585
R133 B.n200 B.n199 585
R134 B.n198 B.n197 585
R135 B.n196 B.n195 585
R136 B.n194 B.n193 585
R137 B.n192 B.n191 585
R138 B.n190 B.n189 585
R139 B.n187 B.n186 585
R140 B.n185 B.n184 585
R141 B.n183 B.n182 585
R142 B.n181 B.n180 585
R143 B.n179 B.n178 585
R144 B.n177 B.n176 585
R145 B.n175 B.n174 585
R146 B.n173 B.n167 585
R147 B.n221 B.n167 585
R148 B.n225 B.n153 585
R149 B.n153 B.n152 585
R150 B.n227 B.n226 585
R151 B.n228 B.n227 585
R152 B.n147 B.n146 585
R153 B.n148 B.n147 585
R154 B.n236 B.n235 585
R155 B.n235 B.n234 585
R156 B.n237 B.n145 585
R157 B.n145 B.n144 585
R158 B.n239 B.n238 585
R159 B.n240 B.n239 585
R160 B.n139 B.n138 585
R161 B.n140 B.n139 585
R162 B.n248 B.n247 585
R163 B.n247 B.n246 585
R164 B.n249 B.n137 585
R165 B.n137 B.n136 585
R166 B.n251 B.n250 585
R167 B.n252 B.n251 585
R168 B.n131 B.n130 585
R169 B.n132 B.n131 585
R170 B.n261 B.n260 585
R171 B.n260 B.n259 585
R172 B.n262 B.n129 585
R173 B.n258 B.n129 585
R174 B.n264 B.n263 585
R175 B.n265 B.n264 585
R176 B.n124 B.n123 585
R177 B.n125 B.n124 585
R178 B.n273 B.n272 585
R179 B.n272 B.n271 585
R180 B.n274 B.n122 585
R181 B.n122 B.n121 585
R182 B.n276 B.n275 585
R183 B.n277 B.n276 585
R184 B.n116 B.n115 585
R185 B.n117 B.n116 585
R186 B.n286 B.n285 585
R187 B.n285 B.n284 585
R188 B.n287 B.n114 585
R189 B.n114 B.n113 585
R190 B.n289 B.n288 585
R191 B.n290 B.n289 585
R192 B.n2 B.n0 585
R193 B.n4 B.n2 585
R194 B.n3 B.n1 585
R195 B.n374 B.n3 585
R196 B.n372 B.n371 585
R197 B.n373 B.n372 585
R198 B.n370 B.n9 585
R199 B.n9 B.n8 585
R200 B.n369 B.n368 585
R201 B.n368 B.n367 585
R202 B.n11 B.n10 585
R203 B.n366 B.n11 585
R204 B.n364 B.n363 585
R205 B.n365 B.n364 585
R206 B.n362 B.n16 585
R207 B.n16 B.n15 585
R208 B.n361 B.n360 585
R209 B.n360 B.n359 585
R210 B.n18 B.n17 585
R211 B.n358 B.n18 585
R212 B.n356 B.n355 585
R213 B.n357 B.n356 585
R214 B.n354 B.n22 585
R215 B.n25 B.n22 585
R216 B.n353 B.n352 585
R217 B.n352 B.n351 585
R218 B.n24 B.n23 585
R219 B.n350 B.n24 585
R220 B.n348 B.n347 585
R221 B.n349 B.n348 585
R222 B.n346 B.n30 585
R223 B.n30 B.n29 585
R224 B.n345 B.n344 585
R225 B.n344 B.n343 585
R226 B.n32 B.n31 585
R227 B.n342 B.n32 585
R228 B.n340 B.n339 585
R229 B.n341 B.n340 585
R230 B.n338 B.n37 585
R231 B.n37 B.n36 585
R232 B.n337 B.n336 585
R233 B.n336 B.n335 585
R234 B.n39 B.n38 585
R235 B.n334 B.n39 585
R236 B.n332 B.n331 585
R237 B.n333 B.n332 585
R238 B.n330 B.n44 585
R239 B.n44 B.n43 585
R240 B.n377 B.n376 585
R241 B.n376 B.n375 585
R242 B.n223 B.n153 502.111
R243 B.n328 B.n44 502.111
R244 B.n167 B.n151 502.111
R245 B.n324 B.n59 502.111
R246 B.n171 B.t13 262.974
R247 B.n169 B.t19 262.974
R248 B.n63 B.t15 262.974
R249 B.n60 B.t8 262.974
R250 B.n326 B.n325 256.663
R251 B.n326 B.n57 256.663
R252 B.n326 B.n56 256.663
R253 B.n326 B.n55 256.663
R254 B.n326 B.n54 256.663
R255 B.n326 B.n53 256.663
R256 B.n326 B.n52 256.663
R257 B.n326 B.n51 256.663
R258 B.n326 B.n50 256.663
R259 B.n326 B.n49 256.663
R260 B.n326 B.n48 256.663
R261 B.n326 B.n47 256.663
R262 B.n327 B.n326 256.663
R263 B.n222 B.n221 256.663
R264 B.n221 B.n156 256.663
R265 B.n221 B.n157 256.663
R266 B.n221 B.n158 256.663
R267 B.n221 B.n159 256.663
R268 B.n221 B.n160 256.663
R269 B.n221 B.n161 256.663
R270 B.n221 B.n162 256.663
R271 B.n221 B.n163 256.663
R272 B.n221 B.n164 256.663
R273 B.n221 B.n165 256.663
R274 B.n221 B.n166 256.663
R275 B.n172 B.t12 238.345
R276 B.n170 B.t18 238.345
R277 B.n64 B.t16 238.345
R278 B.n61 B.t9 238.345
R279 B.n221 B.n152 236.579
R280 B.n326 B.n43 236.579
R281 B.n171 B.t10 205.225
R282 B.n169 B.t17 205.225
R283 B.n63 B.t14 205.225
R284 B.n60 B.t6 205.225
R285 B.n227 B.n153 163.367
R286 B.n227 B.n147 163.367
R287 B.n235 B.n147 163.367
R288 B.n235 B.n145 163.367
R289 B.n239 B.n145 163.367
R290 B.n239 B.n139 163.367
R291 B.n247 B.n139 163.367
R292 B.n247 B.n137 163.367
R293 B.n251 B.n137 163.367
R294 B.n251 B.n131 163.367
R295 B.n260 B.n131 163.367
R296 B.n260 B.n129 163.367
R297 B.n264 B.n129 163.367
R298 B.n264 B.n124 163.367
R299 B.n272 B.n124 163.367
R300 B.n272 B.n122 163.367
R301 B.n276 B.n122 163.367
R302 B.n276 B.n116 163.367
R303 B.n285 B.n116 163.367
R304 B.n285 B.n114 163.367
R305 B.n289 B.n114 163.367
R306 B.n289 B.n2 163.367
R307 B.n376 B.n2 163.367
R308 B.n376 B.n3 163.367
R309 B.n372 B.n3 163.367
R310 B.n372 B.n9 163.367
R311 B.n368 B.n9 163.367
R312 B.n368 B.n11 163.367
R313 B.n364 B.n11 163.367
R314 B.n364 B.n16 163.367
R315 B.n360 B.n16 163.367
R316 B.n360 B.n18 163.367
R317 B.n356 B.n18 163.367
R318 B.n356 B.n22 163.367
R319 B.n352 B.n22 163.367
R320 B.n352 B.n24 163.367
R321 B.n348 B.n24 163.367
R322 B.n348 B.n30 163.367
R323 B.n344 B.n30 163.367
R324 B.n344 B.n32 163.367
R325 B.n340 B.n32 163.367
R326 B.n340 B.n37 163.367
R327 B.n336 B.n37 163.367
R328 B.n336 B.n39 163.367
R329 B.n332 B.n39 163.367
R330 B.n332 B.n44 163.367
R331 B.n220 B.n155 163.367
R332 B.n220 B.n168 163.367
R333 B.n216 B.n215 163.367
R334 B.n212 B.n211 163.367
R335 B.n207 B.n206 163.367
R336 B.n203 B.n202 163.367
R337 B.n199 B.n198 163.367
R338 B.n195 B.n194 163.367
R339 B.n191 B.n190 163.367
R340 B.n186 B.n185 163.367
R341 B.n182 B.n181 163.367
R342 B.n178 B.n177 163.367
R343 B.n174 B.n167 163.367
R344 B.n229 B.n151 163.367
R345 B.n229 B.n149 163.367
R346 B.n233 B.n149 163.367
R347 B.n233 B.n143 163.367
R348 B.n241 B.n143 163.367
R349 B.n241 B.n141 163.367
R350 B.n245 B.n141 163.367
R351 B.n245 B.n135 163.367
R352 B.n253 B.n135 163.367
R353 B.n253 B.n133 163.367
R354 B.n257 B.n133 163.367
R355 B.n257 B.n128 163.367
R356 B.n266 B.n128 163.367
R357 B.n266 B.n126 163.367
R358 B.n270 B.n126 163.367
R359 B.n270 B.n120 163.367
R360 B.n278 B.n120 163.367
R361 B.n278 B.n118 163.367
R362 B.n283 B.n118 163.367
R363 B.n283 B.n112 163.367
R364 B.n291 B.n112 163.367
R365 B.n292 B.n291 163.367
R366 B.n292 B.n5 163.367
R367 B.n6 B.n5 163.367
R368 B.n7 B.n6 163.367
R369 B.n297 B.n7 163.367
R370 B.n297 B.n12 163.367
R371 B.n13 B.n12 163.367
R372 B.n14 B.n13 163.367
R373 B.n302 B.n14 163.367
R374 B.n302 B.n19 163.367
R375 B.n20 B.n19 163.367
R376 B.n21 B.n20 163.367
R377 B.n307 B.n21 163.367
R378 B.n307 B.n26 163.367
R379 B.n27 B.n26 163.367
R380 B.n28 B.n27 163.367
R381 B.n312 B.n28 163.367
R382 B.n312 B.n33 163.367
R383 B.n34 B.n33 163.367
R384 B.n35 B.n34 163.367
R385 B.n317 B.n35 163.367
R386 B.n317 B.n40 163.367
R387 B.n41 B.n40 163.367
R388 B.n42 B.n41 163.367
R389 B.n59 B.n42 163.367
R390 B.n66 B.n46 163.367
R391 B.n70 B.n69 163.367
R392 B.n74 B.n73 163.367
R393 B.n78 B.n77 163.367
R394 B.n82 B.n81 163.367
R395 B.n86 B.n85 163.367
R396 B.n90 B.n89 163.367
R397 B.n94 B.n93 163.367
R398 B.n98 B.n97 163.367
R399 B.n102 B.n101 163.367
R400 B.n106 B.n105 163.367
R401 B.n108 B.n58 163.367
R402 B.n228 B.n152 126.672
R403 B.n228 B.n148 126.672
R404 B.n234 B.n148 126.672
R405 B.n234 B.n144 126.672
R406 B.n240 B.n144 126.672
R407 B.n246 B.n140 126.672
R408 B.n246 B.n136 126.672
R409 B.n252 B.n136 126.672
R410 B.n252 B.n132 126.672
R411 B.n259 B.n132 126.672
R412 B.n259 B.n258 126.672
R413 B.n265 B.n125 126.672
R414 B.n271 B.n125 126.672
R415 B.n277 B.n121 126.672
R416 B.n277 B.n117 126.672
R417 B.n284 B.n117 126.672
R418 B.n290 B.n113 126.672
R419 B.n290 B.n4 126.672
R420 B.n375 B.n4 126.672
R421 B.n375 B.n374 126.672
R422 B.n374 B.n373 126.672
R423 B.n373 B.n8 126.672
R424 B.n367 B.n366 126.672
R425 B.n366 B.n365 126.672
R426 B.n365 B.n15 126.672
R427 B.n359 B.n358 126.672
R428 B.n358 B.n357 126.672
R429 B.n351 B.n25 126.672
R430 B.n351 B.n350 126.672
R431 B.n350 B.n349 126.672
R432 B.n349 B.n29 126.672
R433 B.n343 B.n29 126.672
R434 B.n343 B.n342 126.672
R435 B.n341 B.n36 126.672
R436 B.n335 B.n36 126.672
R437 B.n335 B.n334 126.672
R438 B.n334 B.n333 126.672
R439 B.n333 B.n43 126.672
R440 B.n265 B.t1 119.222
R441 B.n357 B.t0 119.222
R442 B.t11 B.n140 111.77
R443 B.n342 B.t7 111.77
R444 B.n271 B.t3 100.594
R445 B.n359 B.t5 100.594
R446 B.n223 B.n222 71.676
R447 B.n168 B.n156 71.676
R448 B.n215 B.n157 71.676
R449 B.n211 B.n158 71.676
R450 B.n206 B.n159 71.676
R451 B.n202 B.n160 71.676
R452 B.n198 B.n161 71.676
R453 B.n194 B.n162 71.676
R454 B.n190 B.n163 71.676
R455 B.n185 B.n164 71.676
R456 B.n181 B.n165 71.676
R457 B.n177 B.n166 71.676
R458 B.n328 B.n327 71.676
R459 B.n66 B.n47 71.676
R460 B.n70 B.n48 71.676
R461 B.n74 B.n49 71.676
R462 B.n78 B.n50 71.676
R463 B.n82 B.n51 71.676
R464 B.n86 B.n52 71.676
R465 B.n90 B.n53 71.676
R466 B.n94 B.n54 71.676
R467 B.n98 B.n55 71.676
R468 B.n102 B.n56 71.676
R469 B.n106 B.n57 71.676
R470 B.n325 B.n58 71.676
R471 B.n325 B.n324 71.676
R472 B.n108 B.n57 71.676
R473 B.n105 B.n56 71.676
R474 B.n101 B.n55 71.676
R475 B.n97 B.n54 71.676
R476 B.n93 B.n53 71.676
R477 B.n89 B.n52 71.676
R478 B.n85 B.n51 71.676
R479 B.n81 B.n50 71.676
R480 B.n77 B.n49 71.676
R481 B.n73 B.n48 71.676
R482 B.n69 B.n47 71.676
R483 B.n327 B.n46 71.676
R484 B.n222 B.n155 71.676
R485 B.n216 B.n156 71.676
R486 B.n212 B.n157 71.676
R487 B.n207 B.n158 71.676
R488 B.n203 B.n159 71.676
R489 B.n199 B.n160 71.676
R490 B.n195 B.n161 71.676
R491 B.n191 B.n162 71.676
R492 B.n186 B.n163 71.676
R493 B.n182 B.n164 71.676
R494 B.n178 B.n165 71.676
R495 B.n174 B.n166 71.676
R496 B.n284 B.t2 67.0623
R497 B.n367 B.t4 67.0623
R498 B.t2 B.n113 59.611
R499 B.t4 B.n8 59.611
R500 B.n188 B.n172 59.5399
R501 B.n209 B.n170 59.5399
R502 B.n65 B.n64 59.5399
R503 B.n62 B.n61 59.5399
R504 B.n330 B.n329 32.6249
R505 B.n323 B.n322 32.6249
R506 B.n173 B.n150 32.6249
R507 B.n225 B.n224 32.6249
R508 B.t3 B.n121 26.0801
R509 B.t5 B.n15 26.0801
R510 B.n172 B.n171 24.6308
R511 B.n170 B.n169 24.6308
R512 B.n64 B.n63 24.6308
R513 B.n61 B.n60 24.6308
R514 B B.n377 18.0485
R515 B.n240 B.t11 14.9031
R516 B.t7 B.n341 14.9031
R517 B.n329 B.n45 10.6151
R518 B.n67 B.n45 10.6151
R519 B.n68 B.n67 10.6151
R520 B.n71 B.n68 10.6151
R521 B.n72 B.n71 10.6151
R522 B.n75 B.n72 10.6151
R523 B.n76 B.n75 10.6151
R524 B.n80 B.n79 10.6151
R525 B.n83 B.n80 10.6151
R526 B.n84 B.n83 10.6151
R527 B.n87 B.n84 10.6151
R528 B.n88 B.n87 10.6151
R529 B.n91 B.n88 10.6151
R530 B.n92 B.n91 10.6151
R531 B.n95 B.n92 10.6151
R532 B.n96 B.n95 10.6151
R533 B.n100 B.n99 10.6151
R534 B.n103 B.n100 10.6151
R535 B.n104 B.n103 10.6151
R536 B.n107 B.n104 10.6151
R537 B.n109 B.n107 10.6151
R538 B.n110 B.n109 10.6151
R539 B.n323 B.n110 10.6151
R540 B.n230 B.n150 10.6151
R541 B.n231 B.n230 10.6151
R542 B.n232 B.n231 10.6151
R543 B.n232 B.n142 10.6151
R544 B.n242 B.n142 10.6151
R545 B.n243 B.n242 10.6151
R546 B.n244 B.n243 10.6151
R547 B.n244 B.n134 10.6151
R548 B.n254 B.n134 10.6151
R549 B.n255 B.n254 10.6151
R550 B.n256 B.n255 10.6151
R551 B.n256 B.n127 10.6151
R552 B.n267 B.n127 10.6151
R553 B.n268 B.n267 10.6151
R554 B.n269 B.n268 10.6151
R555 B.n269 B.n119 10.6151
R556 B.n279 B.n119 10.6151
R557 B.n280 B.n279 10.6151
R558 B.n282 B.n280 10.6151
R559 B.n282 B.n281 10.6151
R560 B.n281 B.n111 10.6151
R561 B.n293 B.n111 10.6151
R562 B.n294 B.n293 10.6151
R563 B.n295 B.n294 10.6151
R564 B.n296 B.n295 10.6151
R565 B.n298 B.n296 10.6151
R566 B.n299 B.n298 10.6151
R567 B.n300 B.n299 10.6151
R568 B.n301 B.n300 10.6151
R569 B.n303 B.n301 10.6151
R570 B.n304 B.n303 10.6151
R571 B.n305 B.n304 10.6151
R572 B.n306 B.n305 10.6151
R573 B.n308 B.n306 10.6151
R574 B.n309 B.n308 10.6151
R575 B.n310 B.n309 10.6151
R576 B.n311 B.n310 10.6151
R577 B.n313 B.n311 10.6151
R578 B.n314 B.n313 10.6151
R579 B.n315 B.n314 10.6151
R580 B.n316 B.n315 10.6151
R581 B.n318 B.n316 10.6151
R582 B.n319 B.n318 10.6151
R583 B.n320 B.n319 10.6151
R584 B.n321 B.n320 10.6151
R585 B.n322 B.n321 10.6151
R586 B.n224 B.n154 10.6151
R587 B.n219 B.n154 10.6151
R588 B.n219 B.n218 10.6151
R589 B.n218 B.n217 10.6151
R590 B.n217 B.n214 10.6151
R591 B.n214 B.n213 10.6151
R592 B.n213 B.n210 10.6151
R593 B.n208 B.n205 10.6151
R594 B.n205 B.n204 10.6151
R595 B.n204 B.n201 10.6151
R596 B.n201 B.n200 10.6151
R597 B.n200 B.n197 10.6151
R598 B.n197 B.n196 10.6151
R599 B.n196 B.n193 10.6151
R600 B.n193 B.n192 10.6151
R601 B.n192 B.n189 10.6151
R602 B.n187 B.n184 10.6151
R603 B.n184 B.n183 10.6151
R604 B.n183 B.n180 10.6151
R605 B.n180 B.n179 10.6151
R606 B.n179 B.n176 10.6151
R607 B.n176 B.n175 10.6151
R608 B.n175 B.n173 10.6151
R609 B.n226 B.n225 10.6151
R610 B.n226 B.n146 10.6151
R611 B.n236 B.n146 10.6151
R612 B.n237 B.n236 10.6151
R613 B.n238 B.n237 10.6151
R614 B.n238 B.n138 10.6151
R615 B.n248 B.n138 10.6151
R616 B.n249 B.n248 10.6151
R617 B.n250 B.n249 10.6151
R618 B.n250 B.n130 10.6151
R619 B.n261 B.n130 10.6151
R620 B.n262 B.n261 10.6151
R621 B.n263 B.n262 10.6151
R622 B.n263 B.n123 10.6151
R623 B.n273 B.n123 10.6151
R624 B.n274 B.n273 10.6151
R625 B.n275 B.n274 10.6151
R626 B.n275 B.n115 10.6151
R627 B.n286 B.n115 10.6151
R628 B.n287 B.n286 10.6151
R629 B.n288 B.n287 10.6151
R630 B.n288 B.n0 10.6151
R631 B.n371 B.n1 10.6151
R632 B.n371 B.n370 10.6151
R633 B.n370 B.n369 10.6151
R634 B.n369 B.n10 10.6151
R635 B.n363 B.n10 10.6151
R636 B.n363 B.n362 10.6151
R637 B.n362 B.n361 10.6151
R638 B.n361 B.n17 10.6151
R639 B.n355 B.n17 10.6151
R640 B.n355 B.n354 10.6151
R641 B.n354 B.n353 10.6151
R642 B.n353 B.n23 10.6151
R643 B.n347 B.n23 10.6151
R644 B.n347 B.n346 10.6151
R645 B.n346 B.n345 10.6151
R646 B.n345 B.n31 10.6151
R647 B.n339 B.n31 10.6151
R648 B.n339 B.n338 10.6151
R649 B.n338 B.n337 10.6151
R650 B.n337 B.n38 10.6151
R651 B.n331 B.n38 10.6151
R652 B.n331 B.n330 10.6151
R653 B.n76 B.n65 9.36635
R654 B.n99 B.n62 9.36635
R655 B.n210 B.n209 9.36635
R656 B.n188 B.n187 9.36635
R657 B.n258 B.t1 7.45181
R658 B.n25 B.t0 7.45181
R659 B.n377 B.n0 2.81026
R660 B.n377 B.n1 2.81026
R661 B.n79 B.n65 1.24928
R662 B.n96 B.n62 1.24928
R663 B.n209 B.n208 1.24928
R664 B.n189 B.n188 1.24928
R665 VP.n20 VP.n19 161.3
R666 VP.n7 VP.n6 161.3
R667 VP.n8 VP.n3 161.3
R668 VP.n10 VP.n9 161.3
R669 VP.n18 VP.n0 161.3
R670 VP.n17 VP.n16 161.3
R671 VP.n15 VP.n14 161.3
R672 VP.n13 VP.n2 161.3
R673 VP.n12 VP.n11 161.3
R674 VP.n5 VP.t5 76.5514
R675 VP.n12 VP.t2 58.1994
R676 VP.n19 VP.t0 58.1994
R677 VP.n9 VP.t4 58.1994
R678 VP.n14 VP.n13 51.663
R679 VP.n18 VP.n17 51.663
R680 VP.n8 VP.n7 51.663
R681 VP.n6 VP.n5 43.349
R682 VP.n5 VP.n4 42.3693
R683 VP.n11 VP.n10 33.58
R684 VP.n1 VP.t1 16.1526
R685 VP.n4 VP.t3 16.1526
R686 VP.n14 VP.n1 12.234
R687 VP.n17 VP.n1 12.234
R688 VP.n7 VP.n4 12.234
R689 VP.n13 VP.n12 7.30353
R690 VP.n19 VP.n18 7.30353
R691 VP.n9 VP.n8 7.30353
R692 VP.n6 VP.n3 0.189894
R693 VP.n10 VP.n3 0.189894
R694 VP.n11 VP.n2 0.189894
R695 VP.n15 VP.n2 0.189894
R696 VP.n16 VP.n15 0.189894
R697 VP.n16 VP.n0 0.189894
R698 VP.n20 VP.n0 0.189894
R699 VP VP.n20 0.0516364
R700 VTAIL.n11 VTAIL.t5 249.196
R701 VTAIL.n2 VTAIL.t11 249.196
R702 VTAIL.n10 VTAIL.t10 249.196
R703 VTAIL.n7 VTAIL.t0 249.196
R704 VTAIL.n1 VTAIL.n0 217.768
R705 VTAIL.n4 VTAIL.n3 217.768
R706 VTAIL.n9 VTAIL.n8 217.768
R707 VTAIL.n6 VTAIL.n5 217.768
R708 VTAIL.n0 VTAIL.t4 31.4291
R709 VTAIL.n0 VTAIL.t2 31.4291
R710 VTAIL.n3 VTAIL.t8 31.4291
R711 VTAIL.n3 VTAIL.t9 31.4291
R712 VTAIL.n8 VTAIL.t6 31.4291
R713 VTAIL.n8 VTAIL.t7 31.4291
R714 VTAIL.n5 VTAIL.t3 31.4291
R715 VTAIL.n5 VTAIL.t1 31.4291
R716 VTAIL.n6 VTAIL.n4 15.0996
R717 VTAIL.n11 VTAIL.n10 14.0048
R718 VTAIL.n7 VTAIL.n6 1.09533
R719 VTAIL.n10 VTAIL.n9 1.09533
R720 VTAIL.n4 VTAIL.n2 1.09533
R721 VTAIL.n9 VTAIL.n7 1.01774
R722 VTAIL.n2 VTAIL.n1 1.01774
R723 VTAIL VTAIL.n11 0.763431
R724 VTAIL VTAIL.n1 0.332397
R725 VDD1 VDD1.t0 266.753
R726 VDD1.n1 VDD1.t3 266.64
R727 VDD1.n1 VDD1.n0 234.665
R728 VDD1.n3 VDD1.n2 234.446
R729 VDD1.n2 VDD1.t2 31.4291
R730 VDD1.n2 VDD1.t1 31.4291
R731 VDD1.n0 VDD1.t4 31.4291
R732 VDD1.n0 VDD1.t5 31.4291
R733 VDD1.n3 VDD1.n1 28.947
R734 VDD1 VDD1.n3 0.216017
R735 VN.n7 VN.n6 161.3
R736 VN.n15 VN.n14 161.3
R737 VN.n13 VN.n8 161.3
R738 VN.n12 VN.n11 161.3
R739 VN.n5 VN.n0 161.3
R740 VN.n4 VN.n3 161.3
R741 VN.n2 VN.t3 76.5514
R742 VN.n10 VN.t4 76.5514
R743 VN.n6 VN.t2 58.1994
R744 VN.n14 VN.t1 58.1994
R745 VN.n5 VN.n4 51.663
R746 VN.n13 VN.n12 51.663
R747 VN.n11 VN.n10 43.349
R748 VN.n3 VN.n2 43.349
R749 VN.n2 VN.n1 42.3693
R750 VN.n10 VN.n9 42.3693
R751 VN VN.n15 33.9607
R752 VN.n1 VN.t5 16.1526
R753 VN.n9 VN.t0 16.1526
R754 VN.n4 VN.n1 12.234
R755 VN.n12 VN.n9 12.234
R756 VN.n6 VN.n5 7.30353
R757 VN.n14 VN.n13 7.30353
R758 VN.n15 VN.n8 0.189894
R759 VN.n11 VN.n8 0.189894
R760 VN.n3 VN.n0 0.189894
R761 VN.n7 VN.n0 0.189894
R762 VN VN.n7 0.0516364
R763 VDD2.n1 VDD2.t2 266.64
R764 VDD2.n2 VDD2.t4 265.875
R765 VDD2.n1 VDD2.n0 234.665
R766 VDD2 VDD2.n3 234.661
R767 VDD2.n3 VDD2.t5 31.4291
R768 VDD2.n3 VDD2.t1 31.4291
R769 VDD2.n0 VDD2.t0 31.4291
R770 VDD2.n0 VDD2.t3 31.4291
R771 VDD2.n2 VDD2.n1 27.8166
R772 VDD2 VDD2.n2 0.87981
C0 VN VTAIL 1.01835f
C1 VP VTAIL 1.03248f
C2 VP VN 3.21603f
C3 VDD2 VDD1 0.795333f
C4 VDD1 VTAIL 2.41527f
C5 VDD1 VN 0.156861f
C6 VP VDD1 0.758338f
C7 VDD2 VTAIL 2.45736f
C8 VDD2 VN 0.591333f
C9 VP VDD2 0.32614f
C10 VDD2 B 2.478089f
C11 VDD1 B 2.660571f
C12 VTAIL B 2.028146f
C13 VN B 6.541162f
C14 VP B 5.495349f
C15 VDD2.t2 B 0.051177f
C16 VDD2.t0 B 0.010701f
C17 VDD2.t3 B 0.010701f
C18 VDD2.n0 B 0.027167f
C19 VDD2.n1 B 1.02315f
C20 VDD2.t4 B 0.050826f
C21 VDD2.n2 B 1.04835f
C22 VDD2.t5 B 0.010701f
C23 VDD2.t1 B 0.010701f
C24 VDD2.n3 B 0.027162f
C25 VN.n0 B 0.03243f
C26 VN.t5 B 0.025345f
C27 VN.n1 B 0.079336f
C28 VN.t3 B 0.094552f
C29 VN.n2 B 0.086731f
C30 VN.n3 B 0.138625f
C31 VN.n4 B 0.043637f
C32 VN.n5 B 0.011262f
C33 VN.t2 B 0.072047f
C34 VN.n6 B 0.085199f
C35 VN.n7 B 0.025132f
C36 VN.n8 B 0.03243f
C37 VN.t0 B 0.025345f
C38 VN.n9 B 0.079336f
C39 VN.t4 B 0.094552f
C40 VN.n10 B 0.086731f
C41 VN.n11 B 0.138625f
C42 VN.n12 B 0.043637f
C43 VN.n13 B 0.011262f
C44 VN.t1 B 0.072047f
C45 VN.n14 B 0.085199f
C46 VN.n15 B 0.91231f
C47 VDD1.t0 B 0.047688f
C48 VDD1.t3 B 0.047617f
C49 VDD1.t4 B 0.009957f
C50 VDD1.t5 B 0.009957f
C51 VDD1.n0 B 0.025277f
C52 VDD1.n1 B 1.01226f
C53 VDD1.t2 B 0.009957f
C54 VDD1.t1 B 0.009957f
C55 VDD1.n2 B 0.025142f
C56 VDD1.n3 B 1.01182f
C57 VTAIL.t4 B 0.015983f
C58 VTAIL.t2 B 0.015983f
C59 VTAIL.n0 B 0.03462f
C60 VTAIL.n1 B 0.182713f
C61 VTAIL.t11 B 0.070362f
C62 VTAIL.n2 B 0.269484f
C63 VTAIL.t8 B 0.015983f
C64 VTAIL.t9 B 0.015983f
C65 VTAIL.n3 B 0.03462f
C66 VTAIL.n4 B 0.875197f
C67 VTAIL.t3 B 0.015983f
C68 VTAIL.t1 B 0.015983f
C69 VTAIL.n5 B 0.03462f
C70 VTAIL.n6 B 0.875197f
C71 VTAIL.t0 B 0.070362f
C72 VTAIL.n7 B 0.269484f
C73 VTAIL.t6 B 0.015983f
C74 VTAIL.t7 B 0.015983f
C75 VTAIL.n8 B 0.03462f
C76 VTAIL.n9 B 0.261636f
C77 VTAIL.t10 B 0.070362f
C78 VTAIL.n10 B 0.769788f
C79 VTAIL.t5 B 0.070362f
C80 VTAIL.n11 B 0.735455f
C81 VP.n0 B 0.032899f
C82 VP.t1 B 0.025711f
C83 VP.n1 B 0.048472f
C84 VP.n2 B 0.032899f
C85 VP.n3 B 0.032899f
C86 VP.t4 B 0.073089f
C87 VP.t3 B 0.025711f
C88 VP.n4 B 0.080482f
C89 VP.t5 B 0.095919f
C90 VP.n5 B 0.087984f
C91 VP.n6 B 0.140628f
C92 VP.n7 B 0.044267f
C93 VP.n8 B 0.011425f
C94 VP.n9 B 0.08643f
C95 VP.n10 B 0.903557f
C96 VP.n11 B 0.938775f
C97 VP.t2 B 0.073089f
C98 VP.n12 B 0.08643f
C99 VP.n13 B 0.011425f
C100 VP.n14 B 0.044267f
C101 VP.n15 B 0.032899f
C102 VP.n16 B 0.032899f
C103 VP.n17 B 0.044267f
C104 VP.n18 B 0.011425f
C105 VP.t0 B 0.073089f
C106 VP.n19 B 0.08643f
C107 VP.n20 B 0.025495f
.ends

