* NGSPICE file created from diff_pair_sample_1410.ext - technology: sky130A

.subckt diff_pair_sample_1410 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=3.23895 pd=19.96 as=7.6557 ps=40.04 w=19.63 l=0.44
X1 VTAIL.t6 VP.t1 VDD1.t2 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=3.23895 ps=19.96 w=19.63 l=0.44
X2 VDD2.t3 VN.t0 VTAIL.t1 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=3.23895 pd=19.96 as=7.6557 ps=40.04 w=19.63 l=0.44
X3 VDD2.t2 VN.t1 VTAIL.t2 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=3.23895 pd=19.96 as=7.6557 ps=40.04 w=19.63 l=0.44
X4 B.t11 B.t9 B.t10 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=0 ps=0 w=19.63 l=0.44
X5 VTAIL.t3 VN.t2 VDD2.t1 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=3.23895 ps=19.96 w=19.63 l=0.44
X6 VDD1.t1 VP.t2 VTAIL.t7 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=3.23895 pd=19.96 as=7.6557 ps=40.04 w=19.63 l=0.44
X7 B.t8 B.t6 B.t7 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=0 ps=0 w=19.63 l=0.44
X8 B.t5 B.t3 B.t4 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=0 ps=0 w=19.63 l=0.44
X9 VTAIL.t0 VN.t3 VDD2.t0 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=3.23895 ps=19.96 w=19.63 l=0.44
X10 VTAIL.t5 VP.t3 VDD1.t0 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=3.23895 ps=19.96 w=19.63 l=0.44
X11 B.t2 B.t0 B.t1 w_n1432_n4894# sky130_fd_pr__pfet_01v8 ad=7.6557 pd=40.04 as=0 ps=0 w=19.63 l=0.44
R0 VP.n0 VP.t3 1186
R1 VP.n0 VP.t0 1185.97
R2 VP.n2 VP.t1 1165.02
R3 VP.n3 VP.t2 1165.02
R4 VP.n4 VP.n3 161.3
R5 VP.n2 VP.n1 161.3
R6 VP.n1 VP.n0 115.608
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n874 VTAIL.n770 756.745
R11 VTAIL.n104 VTAIL.n0 756.745
R12 VTAIL.n214 VTAIL.n110 756.745
R13 VTAIL.n324 VTAIL.n220 756.745
R14 VTAIL.n764 VTAIL.n660 756.745
R15 VTAIL.n654 VTAIL.n550 756.745
R16 VTAIL.n544 VTAIL.n440 756.745
R17 VTAIL.n434 VTAIL.n330 756.745
R18 VTAIL.n807 VTAIL.n806 585
R19 VTAIL.n809 VTAIL.n808 585
R20 VTAIL.n802 VTAIL.n801 585
R21 VTAIL.n815 VTAIL.n814 585
R22 VTAIL.n817 VTAIL.n816 585
R23 VTAIL.n798 VTAIL.n797 585
R24 VTAIL.n823 VTAIL.n822 585
R25 VTAIL.n825 VTAIL.n824 585
R26 VTAIL.n794 VTAIL.n793 585
R27 VTAIL.n831 VTAIL.n830 585
R28 VTAIL.n833 VTAIL.n832 585
R29 VTAIL.n790 VTAIL.n789 585
R30 VTAIL.n839 VTAIL.n838 585
R31 VTAIL.n841 VTAIL.n840 585
R32 VTAIL.n786 VTAIL.n785 585
R33 VTAIL.n848 VTAIL.n847 585
R34 VTAIL.n849 VTAIL.n784 585
R35 VTAIL.n851 VTAIL.n850 585
R36 VTAIL.n782 VTAIL.n781 585
R37 VTAIL.n857 VTAIL.n856 585
R38 VTAIL.n859 VTAIL.n858 585
R39 VTAIL.n778 VTAIL.n777 585
R40 VTAIL.n865 VTAIL.n864 585
R41 VTAIL.n867 VTAIL.n866 585
R42 VTAIL.n774 VTAIL.n773 585
R43 VTAIL.n873 VTAIL.n872 585
R44 VTAIL.n875 VTAIL.n874 585
R45 VTAIL.n37 VTAIL.n36 585
R46 VTAIL.n39 VTAIL.n38 585
R47 VTAIL.n32 VTAIL.n31 585
R48 VTAIL.n45 VTAIL.n44 585
R49 VTAIL.n47 VTAIL.n46 585
R50 VTAIL.n28 VTAIL.n27 585
R51 VTAIL.n53 VTAIL.n52 585
R52 VTAIL.n55 VTAIL.n54 585
R53 VTAIL.n24 VTAIL.n23 585
R54 VTAIL.n61 VTAIL.n60 585
R55 VTAIL.n63 VTAIL.n62 585
R56 VTAIL.n20 VTAIL.n19 585
R57 VTAIL.n69 VTAIL.n68 585
R58 VTAIL.n71 VTAIL.n70 585
R59 VTAIL.n16 VTAIL.n15 585
R60 VTAIL.n78 VTAIL.n77 585
R61 VTAIL.n79 VTAIL.n14 585
R62 VTAIL.n81 VTAIL.n80 585
R63 VTAIL.n12 VTAIL.n11 585
R64 VTAIL.n87 VTAIL.n86 585
R65 VTAIL.n89 VTAIL.n88 585
R66 VTAIL.n8 VTAIL.n7 585
R67 VTAIL.n95 VTAIL.n94 585
R68 VTAIL.n97 VTAIL.n96 585
R69 VTAIL.n4 VTAIL.n3 585
R70 VTAIL.n103 VTAIL.n102 585
R71 VTAIL.n105 VTAIL.n104 585
R72 VTAIL.n147 VTAIL.n146 585
R73 VTAIL.n149 VTAIL.n148 585
R74 VTAIL.n142 VTAIL.n141 585
R75 VTAIL.n155 VTAIL.n154 585
R76 VTAIL.n157 VTAIL.n156 585
R77 VTAIL.n138 VTAIL.n137 585
R78 VTAIL.n163 VTAIL.n162 585
R79 VTAIL.n165 VTAIL.n164 585
R80 VTAIL.n134 VTAIL.n133 585
R81 VTAIL.n171 VTAIL.n170 585
R82 VTAIL.n173 VTAIL.n172 585
R83 VTAIL.n130 VTAIL.n129 585
R84 VTAIL.n179 VTAIL.n178 585
R85 VTAIL.n181 VTAIL.n180 585
R86 VTAIL.n126 VTAIL.n125 585
R87 VTAIL.n188 VTAIL.n187 585
R88 VTAIL.n189 VTAIL.n124 585
R89 VTAIL.n191 VTAIL.n190 585
R90 VTAIL.n122 VTAIL.n121 585
R91 VTAIL.n197 VTAIL.n196 585
R92 VTAIL.n199 VTAIL.n198 585
R93 VTAIL.n118 VTAIL.n117 585
R94 VTAIL.n205 VTAIL.n204 585
R95 VTAIL.n207 VTAIL.n206 585
R96 VTAIL.n114 VTAIL.n113 585
R97 VTAIL.n213 VTAIL.n212 585
R98 VTAIL.n215 VTAIL.n214 585
R99 VTAIL.n257 VTAIL.n256 585
R100 VTAIL.n259 VTAIL.n258 585
R101 VTAIL.n252 VTAIL.n251 585
R102 VTAIL.n265 VTAIL.n264 585
R103 VTAIL.n267 VTAIL.n266 585
R104 VTAIL.n248 VTAIL.n247 585
R105 VTAIL.n273 VTAIL.n272 585
R106 VTAIL.n275 VTAIL.n274 585
R107 VTAIL.n244 VTAIL.n243 585
R108 VTAIL.n281 VTAIL.n280 585
R109 VTAIL.n283 VTAIL.n282 585
R110 VTAIL.n240 VTAIL.n239 585
R111 VTAIL.n289 VTAIL.n288 585
R112 VTAIL.n291 VTAIL.n290 585
R113 VTAIL.n236 VTAIL.n235 585
R114 VTAIL.n298 VTAIL.n297 585
R115 VTAIL.n299 VTAIL.n234 585
R116 VTAIL.n301 VTAIL.n300 585
R117 VTAIL.n232 VTAIL.n231 585
R118 VTAIL.n307 VTAIL.n306 585
R119 VTAIL.n309 VTAIL.n308 585
R120 VTAIL.n228 VTAIL.n227 585
R121 VTAIL.n315 VTAIL.n314 585
R122 VTAIL.n317 VTAIL.n316 585
R123 VTAIL.n224 VTAIL.n223 585
R124 VTAIL.n323 VTAIL.n322 585
R125 VTAIL.n325 VTAIL.n324 585
R126 VTAIL.n765 VTAIL.n764 585
R127 VTAIL.n763 VTAIL.n762 585
R128 VTAIL.n664 VTAIL.n663 585
R129 VTAIL.n757 VTAIL.n756 585
R130 VTAIL.n755 VTAIL.n754 585
R131 VTAIL.n668 VTAIL.n667 585
R132 VTAIL.n749 VTAIL.n748 585
R133 VTAIL.n747 VTAIL.n746 585
R134 VTAIL.n672 VTAIL.n671 585
R135 VTAIL.n676 VTAIL.n674 585
R136 VTAIL.n741 VTAIL.n740 585
R137 VTAIL.n739 VTAIL.n738 585
R138 VTAIL.n678 VTAIL.n677 585
R139 VTAIL.n733 VTAIL.n732 585
R140 VTAIL.n731 VTAIL.n730 585
R141 VTAIL.n682 VTAIL.n681 585
R142 VTAIL.n725 VTAIL.n724 585
R143 VTAIL.n723 VTAIL.n722 585
R144 VTAIL.n686 VTAIL.n685 585
R145 VTAIL.n717 VTAIL.n716 585
R146 VTAIL.n715 VTAIL.n714 585
R147 VTAIL.n690 VTAIL.n689 585
R148 VTAIL.n709 VTAIL.n708 585
R149 VTAIL.n707 VTAIL.n706 585
R150 VTAIL.n694 VTAIL.n693 585
R151 VTAIL.n701 VTAIL.n700 585
R152 VTAIL.n699 VTAIL.n698 585
R153 VTAIL.n655 VTAIL.n654 585
R154 VTAIL.n653 VTAIL.n652 585
R155 VTAIL.n554 VTAIL.n553 585
R156 VTAIL.n647 VTAIL.n646 585
R157 VTAIL.n645 VTAIL.n644 585
R158 VTAIL.n558 VTAIL.n557 585
R159 VTAIL.n639 VTAIL.n638 585
R160 VTAIL.n637 VTAIL.n636 585
R161 VTAIL.n562 VTAIL.n561 585
R162 VTAIL.n566 VTAIL.n564 585
R163 VTAIL.n631 VTAIL.n630 585
R164 VTAIL.n629 VTAIL.n628 585
R165 VTAIL.n568 VTAIL.n567 585
R166 VTAIL.n623 VTAIL.n622 585
R167 VTAIL.n621 VTAIL.n620 585
R168 VTAIL.n572 VTAIL.n571 585
R169 VTAIL.n615 VTAIL.n614 585
R170 VTAIL.n613 VTAIL.n612 585
R171 VTAIL.n576 VTAIL.n575 585
R172 VTAIL.n607 VTAIL.n606 585
R173 VTAIL.n605 VTAIL.n604 585
R174 VTAIL.n580 VTAIL.n579 585
R175 VTAIL.n599 VTAIL.n598 585
R176 VTAIL.n597 VTAIL.n596 585
R177 VTAIL.n584 VTAIL.n583 585
R178 VTAIL.n591 VTAIL.n590 585
R179 VTAIL.n589 VTAIL.n588 585
R180 VTAIL.n545 VTAIL.n544 585
R181 VTAIL.n543 VTAIL.n542 585
R182 VTAIL.n444 VTAIL.n443 585
R183 VTAIL.n537 VTAIL.n536 585
R184 VTAIL.n535 VTAIL.n534 585
R185 VTAIL.n448 VTAIL.n447 585
R186 VTAIL.n529 VTAIL.n528 585
R187 VTAIL.n527 VTAIL.n526 585
R188 VTAIL.n452 VTAIL.n451 585
R189 VTAIL.n456 VTAIL.n454 585
R190 VTAIL.n521 VTAIL.n520 585
R191 VTAIL.n519 VTAIL.n518 585
R192 VTAIL.n458 VTAIL.n457 585
R193 VTAIL.n513 VTAIL.n512 585
R194 VTAIL.n511 VTAIL.n510 585
R195 VTAIL.n462 VTAIL.n461 585
R196 VTAIL.n505 VTAIL.n504 585
R197 VTAIL.n503 VTAIL.n502 585
R198 VTAIL.n466 VTAIL.n465 585
R199 VTAIL.n497 VTAIL.n496 585
R200 VTAIL.n495 VTAIL.n494 585
R201 VTAIL.n470 VTAIL.n469 585
R202 VTAIL.n489 VTAIL.n488 585
R203 VTAIL.n487 VTAIL.n486 585
R204 VTAIL.n474 VTAIL.n473 585
R205 VTAIL.n481 VTAIL.n480 585
R206 VTAIL.n479 VTAIL.n478 585
R207 VTAIL.n435 VTAIL.n434 585
R208 VTAIL.n433 VTAIL.n432 585
R209 VTAIL.n334 VTAIL.n333 585
R210 VTAIL.n427 VTAIL.n426 585
R211 VTAIL.n425 VTAIL.n424 585
R212 VTAIL.n338 VTAIL.n337 585
R213 VTAIL.n419 VTAIL.n418 585
R214 VTAIL.n417 VTAIL.n416 585
R215 VTAIL.n342 VTAIL.n341 585
R216 VTAIL.n346 VTAIL.n344 585
R217 VTAIL.n411 VTAIL.n410 585
R218 VTAIL.n409 VTAIL.n408 585
R219 VTAIL.n348 VTAIL.n347 585
R220 VTAIL.n403 VTAIL.n402 585
R221 VTAIL.n401 VTAIL.n400 585
R222 VTAIL.n352 VTAIL.n351 585
R223 VTAIL.n395 VTAIL.n394 585
R224 VTAIL.n393 VTAIL.n392 585
R225 VTAIL.n356 VTAIL.n355 585
R226 VTAIL.n387 VTAIL.n386 585
R227 VTAIL.n385 VTAIL.n384 585
R228 VTAIL.n360 VTAIL.n359 585
R229 VTAIL.n379 VTAIL.n378 585
R230 VTAIL.n377 VTAIL.n376 585
R231 VTAIL.n364 VTAIL.n363 585
R232 VTAIL.n371 VTAIL.n370 585
R233 VTAIL.n369 VTAIL.n368 585
R234 VTAIL.n805 VTAIL.t1 327.466
R235 VTAIL.n35 VTAIL.t0 327.466
R236 VTAIL.n145 VTAIL.t7 327.466
R237 VTAIL.n255 VTAIL.t6 327.466
R238 VTAIL.n697 VTAIL.t4 327.466
R239 VTAIL.n587 VTAIL.t5 327.466
R240 VTAIL.n477 VTAIL.t2 327.466
R241 VTAIL.n367 VTAIL.t3 327.466
R242 VTAIL.n808 VTAIL.n807 171.744
R243 VTAIL.n808 VTAIL.n801 171.744
R244 VTAIL.n815 VTAIL.n801 171.744
R245 VTAIL.n816 VTAIL.n815 171.744
R246 VTAIL.n816 VTAIL.n797 171.744
R247 VTAIL.n823 VTAIL.n797 171.744
R248 VTAIL.n824 VTAIL.n823 171.744
R249 VTAIL.n824 VTAIL.n793 171.744
R250 VTAIL.n831 VTAIL.n793 171.744
R251 VTAIL.n832 VTAIL.n831 171.744
R252 VTAIL.n832 VTAIL.n789 171.744
R253 VTAIL.n839 VTAIL.n789 171.744
R254 VTAIL.n840 VTAIL.n839 171.744
R255 VTAIL.n840 VTAIL.n785 171.744
R256 VTAIL.n848 VTAIL.n785 171.744
R257 VTAIL.n849 VTAIL.n848 171.744
R258 VTAIL.n850 VTAIL.n849 171.744
R259 VTAIL.n850 VTAIL.n781 171.744
R260 VTAIL.n857 VTAIL.n781 171.744
R261 VTAIL.n858 VTAIL.n857 171.744
R262 VTAIL.n858 VTAIL.n777 171.744
R263 VTAIL.n865 VTAIL.n777 171.744
R264 VTAIL.n866 VTAIL.n865 171.744
R265 VTAIL.n866 VTAIL.n773 171.744
R266 VTAIL.n873 VTAIL.n773 171.744
R267 VTAIL.n874 VTAIL.n873 171.744
R268 VTAIL.n38 VTAIL.n37 171.744
R269 VTAIL.n38 VTAIL.n31 171.744
R270 VTAIL.n45 VTAIL.n31 171.744
R271 VTAIL.n46 VTAIL.n45 171.744
R272 VTAIL.n46 VTAIL.n27 171.744
R273 VTAIL.n53 VTAIL.n27 171.744
R274 VTAIL.n54 VTAIL.n53 171.744
R275 VTAIL.n54 VTAIL.n23 171.744
R276 VTAIL.n61 VTAIL.n23 171.744
R277 VTAIL.n62 VTAIL.n61 171.744
R278 VTAIL.n62 VTAIL.n19 171.744
R279 VTAIL.n69 VTAIL.n19 171.744
R280 VTAIL.n70 VTAIL.n69 171.744
R281 VTAIL.n70 VTAIL.n15 171.744
R282 VTAIL.n78 VTAIL.n15 171.744
R283 VTAIL.n79 VTAIL.n78 171.744
R284 VTAIL.n80 VTAIL.n79 171.744
R285 VTAIL.n80 VTAIL.n11 171.744
R286 VTAIL.n87 VTAIL.n11 171.744
R287 VTAIL.n88 VTAIL.n87 171.744
R288 VTAIL.n88 VTAIL.n7 171.744
R289 VTAIL.n95 VTAIL.n7 171.744
R290 VTAIL.n96 VTAIL.n95 171.744
R291 VTAIL.n96 VTAIL.n3 171.744
R292 VTAIL.n103 VTAIL.n3 171.744
R293 VTAIL.n104 VTAIL.n103 171.744
R294 VTAIL.n148 VTAIL.n147 171.744
R295 VTAIL.n148 VTAIL.n141 171.744
R296 VTAIL.n155 VTAIL.n141 171.744
R297 VTAIL.n156 VTAIL.n155 171.744
R298 VTAIL.n156 VTAIL.n137 171.744
R299 VTAIL.n163 VTAIL.n137 171.744
R300 VTAIL.n164 VTAIL.n163 171.744
R301 VTAIL.n164 VTAIL.n133 171.744
R302 VTAIL.n171 VTAIL.n133 171.744
R303 VTAIL.n172 VTAIL.n171 171.744
R304 VTAIL.n172 VTAIL.n129 171.744
R305 VTAIL.n179 VTAIL.n129 171.744
R306 VTAIL.n180 VTAIL.n179 171.744
R307 VTAIL.n180 VTAIL.n125 171.744
R308 VTAIL.n188 VTAIL.n125 171.744
R309 VTAIL.n189 VTAIL.n188 171.744
R310 VTAIL.n190 VTAIL.n189 171.744
R311 VTAIL.n190 VTAIL.n121 171.744
R312 VTAIL.n197 VTAIL.n121 171.744
R313 VTAIL.n198 VTAIL.n197 171.744
R314 VTAIL.n198 VTAIL.n117 171.744
R315 VTAIL.n205 VTAIL.n117 171.744
R316 VTAIL.n206 VTAIL.n205 171.744
R317 VTAIL.n206 VTAIL.n113 171.744
R318 VTAIL.n213 VTAIL.n113 171.744
R319 VTAIL.n214 VTAIL.n213 171.744
R320 VTAIL.n258 VTAIL.n257 171.744
R321 VTAIL.n258 VTAIL.n251 171.744
R322 VTAIL.n265 VTAIL.n251 171.744
R323 VTAIL.n266 VTAIL.n265 171.744
R324 VTAIL.n266 VTAIL.n247 171.744
R325 VTAIL.n273 VTAIL.n247 171.744
R326 VTAIL.n274 VTAIL.n273 171.744
R327 VTAIL.n274 VTAIL.n243 171.744
R328 VTAIL.n281 VTAIL.n243 171.744
R329 VTAIL.n282 VTAIL.n281 171.744
R330 VTAIL.n282 VTAIL.n239 171.744
R331 VTAIL.n289 VTAIL.n239 171.744
R332 VTAIL.n290 VTAIL.n289 171.744
R333 VTAIL.n290 VTAIL.n235 171.744
R334 VTAIL.n298 VTAIL.n235 171.744
R335 VTAIL.n299 VTAIL.n298 171.744
R336 VTAIL.n300 VTAIL.n299 171.744
R337 VTAIL.n300 VTAIL.n231 171.744
R338 VTAIL.n307 VTAIL.n231 171.744
R339 VTAIL.n308 VTAIL.n307 171.744
R340 VTAIL.n308 VTAIL.n227 171.744
R341 VTAIL.n315 VTAIL.n227 171.744
R342 VTAIL.n316 VTAIL.n315 171.744
R343 VTAIL.n316 VTAIL.n223 171.744
R344 VTAIL.n323 VTAIL.n223 171.744
R345 VTAIL.n324 VTAIL.n323 171.744
R346 VTAIL.n764 VTAIL.n763 171.744
R347 VTAIL.n763 VTAIL.n663 171.744
R348 VTAIL.n756 VTAIL.n663 171.744
R349 VTAIL.n756 VTAIL.n755 171.744
R350 VTAIL.n755 VTAIL.n667 171.744
R351 VTAIL.n748 VTAIL.n667 171.744
R352 VTAIL.n748 VTAIL.n747 171.744
R353 VTAIL.n747 VTAIL.n671 171.744
R354 VTAIL.n676 VTAIL.n671 171.744
R355 VTAIL.n740 VTAIL.n676 171.744
R356 VTAIL.n740 VTAIL.n739 171.744
R357 VTAIL.n739 VTAIL.n677 171.744
R358 VTAIL.n732 VTAIL.n677 171.744
R359 VTAIL.n732 VTAIL.n731 171.744
R360 VTAIL.n731 VTAIL.n681 171.744
R361 VTAIL.n724 VTAIL.n681 171.744
R362 VTAIL.n724 VTAIL.n723 171.744
R363 VTAIL.n723 VTAIL.n685 171.744
R364 VTAIL.n716 VTAIL.n685 171.744
R365 VTAIL.n716 VTAIL.n715 171.744
R366 VTAIL.n715 VTAIL.n689 171.744
R367 VTAIL.n708 VTAIL.n689 171.744
R368 VTAIL.n708 VTAIL.n707 171.744
R369 VTAIL.n707 VTAIL.n693 171.744
R370 VTAIL.n700 VTAIL.n693 171.744
R371 VTAIL.n700 VTAIL.n699 171.744
R372 VTAIL.n654 VTAIL.n653 171.744
R373 VTAIL.n653 VTAIL.n553 171.744
R374 VTAIL.n646 VTAIL.n553 171.744
R375 VTAIL.n646 VTAIL.n645 171.744
R376 VTAIL.n645 VTAIL.n557 171.744
R377 VTAIL.n638 VTAIL.n557 171.744
R378 VTAIL.n638 VTAIL.n637 171.744
R379 VTAIL.n637 VTAIL.n561 171.744
R380 VTAIL.n566 VTAIL.n561 171.744
R381 VTAIL.n630 VTAIL.n566 171.744
R382 VTAIL.n630 VTAIL.n629 171.744
R383 VTAIL.n629 VTAIL.n567 171.744
R384 VTAIL.n622 VTAIL.n567 171.744
R385 VTAIL.n622 VTAIL.n621 171.744
R386 VTAIL.n621 VTAIL.n571 171.744
R387 VTAIL.n614 VTAIL.n571 171.744
R388 VTAIL.n614 VTAIL.n613 171.744
R389 VTAIL.n613 VTAIL.n575 171.744
R390 VTAIL.n606 VTAIL.n575 171.744
R391 VTAIL.n606 VTAIL.n605 171.744
R392 VTAIL.n605 VTAIL.n579 171.744
R393 VTAIL.n598 VTAIL.n579 171.744
R394 VTAIL.n598 VTAIL.n597 171.744
R395 VTAIL.n597 VTAIL.n583 171.744
R396 VTAIL.n590 VTAIL.n583 171.744
R397 VTAIL.n590 VTAIL.n589 171.744
R398 VTAIL.n544 VTAIL.n543 171.744
R399 VTAIL.n543 VTAIL.n443 171.744
R400 VTAIL.n536 VTAIL.n443 171.744
R401 VTAIL.n536 VTAIL.n535 171.744
R402 VTAIL.n535 VTAIL.n447 171.744
R403 VTAIL.n528 VTAIL.n447 171.744
R404 VTAIL.n528 VTAIL.n527 171.744
R405 VTAIL.n527 VTAIL.n451 171.744
R406 VTAIL.n456 VTAIL.n451 171.744
R407 VTAIL.n520 VTAIL.n456 171.744
R408 VTAIL.n520 VTAIL.n519 171.744
R409 VTAIL.n519 VTAIL.n457 171.744
R410 VTAIL.n512 VTAIL.n457 171.744
R411 VTAIL.n512 VTAIL.n511 171.744
R412 VTAIL.n511 VTAIL.n461 171.744
R413 VTAIL.n504 VTAIL.n461 171.744
R414 VTAIL.n504 VTAIL.n503 171.744
R415 VTAIL.n503 VTAIL.n465 171.744
R416 VTAIL.n496 VTAIL.n465 171.744
R417 VTAIL.n496 VTAIL.n495 171.744
R418 VTAIL.n495 VTAIL.n469 171.744
R419 VTAIL.n488 VTAIL.n469 171.744
R420 VTAIL.n488 VTAIL.n487 171.744
R421 VTAIL.n487 VTAIL.n473 171.744
R422 VTAIL.n480 VTAIL.n473 171.744
R423 VTAIL.n480 VTAIL.n479 171.744
R424 VTAIL.n434 VTAIL.n433 171.744
R425 VTAIL.n433 VTAIL.n333 171.744
R426 VTAIL.n426 VTAIL.n333 171.744
R427 VTAIL.n426 VTAIL.n425 171.744
R428 VTAIL.n425 VTAIL.n337 171.744
R429 VTAIL.n418 VTAIL.n337 171.744
R430 VTAIL.n418 VTAIL.n417 171.744
R431 VTAIL.n417 VTAIL.n341 171.744
R432 VTAIL.n346 VTAIL.n341 171.744
R433 VTAIL.n410 VTAIL.n346 171.744
R434 VTAIL.n410 VTAIL.n409 171.744
R435 VTAIL.n409 VTAIL.n347 171.744
R436 VTAIL.n402 VTAIL.n347 171.744
R437 VTAIL.n402 VTAIL.n401 171.744
R438 VTAIL.n401 VTAIL.n351 171.744
R439 VTAIL.n394 VTAIL.n351 171.744
R440 VTAIL.n394 VTAIL.n393 171.744
R441 VTAIL.n393 VTAIL.n355 171.744
R442 VTAIL.n386 VTAIL.n355 171.744
R443 VTAIL.n386 VTAIL.n385 171.744
R444 VTAIL.n385 VTAIL.n359 171.744
R445 VTAIL.n378 VTAIL.n359 171.744
R446 VTAIL.n378 VTAIL.n377 171.744
R447 VTAIL.n377 VTAIL.n363 171.744
R448 VTAIL.n370 VTAIL.n363 171.744
R449 VTAIL.n370 VTAIL.n369 171.744
R450 VTAIL.n807 VTAIL.t1 85.8723
R451 VTAIL.n37 VTAIL.t0 85.8723
R452 VTAIL.n147 VTAIL.t7 85.8723
R453 VTAIL.n257 VTAIL.t6 85.8723
R454 VTAIL.n699 VTAIL.t4 85.8723
R455 VTAIL.n589 VTAIL.t5 85.8723
R456 VTAIL.n479 VTAIL.t2 85.8723
R457 VTAIL.n369 VTAIL.t3 85.8723
R458 VTAIL.n879 VTAIL.n878 31.2157
R459 VTAIL.n109 VTAIL.n108 31.2157
R460 VTAIL.n219 VTAIL.n218 31.2157
R461 VTAIL.n329 VTAIL.n328 31.2157
R462 VTAIL.n769 VTAIL.n768 31.2157
R463 VTAIL.n659 VTAIL.n658 31.2157
R464 VTAIL.n549 VTAIL.n548 31.2157
R465 VTAIL.n439 VTAIL.n438 31.2157
R466 VTAIL.n879 VTAIL.n769 29.9531
R467 VTAIL.n439 VTAIL.n329 29.9531
R468 VTAIL.n806 VTAIL.n805 16.3895
R469 VTAIL.n36 VTAIL.n35 16.3895
R470 VTAIL.n146 VTAIL.n145 16.3895
R471 VTAIL.n256 VTAIL.n255 16.3895
R472 VTAIL.n698 VTAIL.n697 16.3895
R473 VTAIL.n588 VTAIL.n587 16.3895
R474 VTAIL.n478 VTAIL.n477 16.3895
R475 VTAIL.n368 VTAIL.n367 16.3895
R476 VTAIL.n851 VTAIL.n782 13.1884
R477 VTAIL.n81 VTAIL.n12 13.1884
R478 VTAIL.n191 VTAIL.n122 13.1884
R479 VTAIL.n301 VTAIL.n232 13.1884
R480 VTAIL.n674 VTAIL.n672 13.1884
R481 VTAIL.n564 VTAIL.n562 13.1884
R482 VTAIL.n454 VTAIL.n452 13.1884
R483 VTAIL.n344 VTAIL.n342 13.1884
R484 VTAIL.n809 VTAIL.n804 12.8005
R485 VTAIL.n852 VTAIL.n784 12.8005
R486 VTAIL.n856 VTAIL.n855 12.8005
R487 VTAIL.n39 VTAIL.n34 12.8005
R488 VTAIL.n82 VTAIL.n14 12.8005
R489 VTAIL.n86 VTAIL.n85 12.8005
R490 VTAIL.n149 VTAIL.n144 12.8005
R491 VTAIL.n192 VTAIL.n124 12.8005
R492 VTAIL.n196 VTAIL.n195 12.8005
R493 VTAIL.n259 VTAIL.n254 12.8005
R494 VTAIL.n302 VTAIL.n234 12.8005
R495 VTAIL.n306 VTAIL.n305 12.8005
R496 VTAIL.n746 VTAIL.n745 12.8005
R497 VTAIL.n742 VTAIL.n741 12.8005
R498 VTAIL.n701 VTAIL.n696 12.8005
R499 VTAIL.n636 VTAIL.n635 12.8005
R500 VTAIL.n632 VTAIL.n631 12.8005
R501 VTAIL.n591 VTAIL.n586 12.8005
R502 VTAIL.n526 VTAIL.n525 12.8005
R503 VTAIL.n522 VTAIL.n521 12.8005
R504 VTAIL.n481 VTAIL.n476 12.8005
R505 VTAIL.n416 VTAIL.n415 12.8005
R506 VTAIL.n412 VTAIL.n411 12.8005
R507 VTAIL.n371 VTAIL.n366 12.8005
R508 VTAIL.n810 VTAIL.n802 12.0247
R509 VTAIL.n847 VTAIL.n846 12.0247
R510 VTAIL.n859 VTAIL.n780 12.0247
R511 VTAIL.n40 VTAIL.n32 12.0247
R512 VTAIL.n77 VTAIL.n76 12.0247
R513 VTAIL.n89 VTAIL.n10 12.0247
R514 VTAIL.n150 VTAIL.n142 12.0247
R515 VTAIL.n187 VTAIL.n186 12.0247
R516 VTAIL.n199 VTAIL.n120 12.0247
R517 VTAIL.n260 VTAIL.n252 12.0247
R518 VTAIL.n297 VTAIL.n296 12.0247
R519 VTAIL.n309 VTAIL.n230 12.0247
R520 VTAIL.n749 VTAIL.n670 12.0247
R521 VTAIL.n738 VTAIL.n675 12.0247
R522 VTAIL.n702 VTAIL.n694 12.0247
R523 VTAIL.n639 VTAIL.n560 12.0247
R524 VTAIL.n628 VTAIL.n565 12.0247
R525 VTAIL.n592 VTAIL.n584 12.0247
R526 VTAIL.n529 VTAIL.n450 12.0247
R527 VTAIL.n518 VTAIL.n455 12.0247
R528 VTAIL.n482 VTAIL.n474 12.0247
R529 VTAIL.n419 VTAIL.n340 12.0247
R530 VTAIL.n408 VTAIL.n345 12.0247
R531 VTAIL.n372 VTAIL.n364 12.0247
R532 VTAIL.n814 VTAIL.n813 11.249
R533 VTAIL.n845 VTAIL.n786 11.249
R534 VTAIL.n860 VTAIL.n778 11.249
R535 VTAIL.n44 VTAIL.n43 11.249
R536 VTAIL.n75 VTAIL.n16 11.249
R537 VTAIL.n90 VTAIL.n8 11.249
R538 VTAIL.n154 VTAIL.n153 11.249
R539 VTAIL.n185 VTAIL.n126 11.249
R540 VTAIL.n200 VTAIL.n118 11.249
R541 VTAIL.n264 VTAIL.n263 11.249
R542 VTAIL.n295 VTAIL.n236 11.249
R543 VTAIL.n310 VTAIL.n228 11.249
R544 VTAIL.n750 VTAIL.n668 11.249
R545 VTAIL.n737 VTAIL.n678 11.249
R546 VTAIL.n706 VTAIL.n705 11.249
R547 VTAIL.n640 VTAIL.n558 11.249
R548 VTAIL.n627 VTAIL.n568 11.249
R549 VTAIL.n596 VTAIL.n595 11.249
R550 VTAIL.n530 VTAIL.n448 11.249
R551 VTAIL.n517 VTAIL.n458 11.249
R552 VTAIL.n486 VTAIL.n485 11.249
R553 VTAIL.n420 VTAIL.n338 11.249
R554 VTAIL.n407 VTAIL.n348 11.249
R555 VTAIL.n376 VTAIL.n375 11.249
R556 VTAIL.n817 VTAIL.n800 10.4732
R557 VTAIL.n842 VTAIL.n841 10.4732
R558 VTAIL.n864 VTAIL.n863 10.4732
R559 VTAIL.n47 VTAIL.n30 10.4732
R560 VTAIL.n72 VTAIL.n71 10.4732
R561 VTAIL.n94 VTAIL.n93 10.4732
R562 VTAIL.n157 VTAIL.n140 10.4732
R563 VTAIL.n182 VTAIL.n181 10.4732
R564 VTAIL.n204 VTAIL.n203 10.4732
R565 VTAIL.n267 VTAIL.n250 10.4732
R566 VTAIL.n292 VTAIL.n291 10.4732
R567 VTAIL.n314 VTAIL.n313 10.4732
R568 VTAIL.n754 VTAIL.n753 10.4732
R569 VTAIL.n734 VTAIL.n733 10.4732
R570 VTAIL.n709 VTAIL.n692 10.4732
R571 VTAIL.n644 VTAIL.n643 10.4732
R572 VTAIL.n624 VTAIL.n623 10.4732
R573 VTAIL.n599 VTAIL.n582 10.4732
R574 VTAIL.n534 VTAIL.n533 10.4732
R575 VTAIL.n514 VTAIL.n513 10.4732
R576 VTAIL.n489 VTAIL.n472 10.4732
R577 VTAIL.n424 VTAIL.n423 10.4732
R578 VTAIL.n404 VTAIL.n403 10.4732
R579 VTAIL.n379 VTAIL.n362 10.4732
R580 VTAIL.n818 VTAIL.n798 9.69747
R581 VTAIL.n838 VTAIL.n788 9.69747
R582 VTAIL.n867 VTAIL.n776 9.69747
R583 VTAIL.n48 VTAIL.n28 9.69747
R584 VTAIL.n68 VTAIL.n18 9.69747
R585 VTAIL.n97 VTAIL.n6 9.69747
R586 VTAIL.n158 VTAIL.n138 9.69747
R587 VTAIL.n178 VTAIL.n128 9.69747
R588 VTAIL.n207 VTAIL.n116 9.69747
R589 VTAIL.n268 VTAIL.n248 9.69747
R590 VTAIL.n288 VTAIL.n238 9.69747
R591 VTAIL.n317 VTAIL.n226 9.69747
R592 VTAIL.n757 VTAIL.n666 9.69747
R593 VTAIL.n730 VTAIL.n680 9.69747
R594 VTAIL.n710 VTAIL.n690 9.69747
R595 VTAIL.n647 VTAIL.n556 9.69747
R596 VTAIL.n620 VTAIL.n570 9.69747
R597 VTAIL.n600 VTAIL.n580 9.69747
R598 VTAIL.n537 VTAIL.n446 9.69747
R599 VTAIL.n510 VTAIL.n460 9.69747
R600 VTAIL.n490 VTAIL.n470 9.69747
R601 VTAIL.n427 VTAIL.n336 9.69747
R602 VTAIL.n400 VTAIL.n350 9.69747
R603 VTAIL.n380 VTAIL.n360 9.69747
R604 VTAIL.n878 VTAIL.n877 9.45567
R605 VTAIL.n108 VTAIL.n107 9.45567
R606 VTAIL.n218 VTAIL.n217 9.45567
R607 VTAIL.n328 VTAIL.n327 9.45567
R608 VTAIL.n768 VTAIL.n767 9.45567
R609 VTAIL.n658 VTAIL.n657 9.45567
R610 VTAIL.n548 VTAIL.n547 9.45567
R611 VTAIL.n438 VTAIL.n437 9.45567
R612 VTAIL.n877 VTAIL.n876 9.3005
R613 VTAIL.n871 VTAIL.n870 9.3005
R614 VTAIL.n869 VTAIL.n868 9.3005
R615 VTAIL.n776 VTAIL.n775 9.3005
R616 VTAIL.n863 VTAIL.n862 9.3005
R617 VTAIL.n861 VTAIL.n860 9.3005
R618 VTAIL.n780 VTAIL.n779 9.3005
R619 VTAIL.n855 VTAIL.n854 9.3005
R620 VTAIL.n827 VTAIL.n826 9.3005
R621 VTAIL.n796 VTAIL.n795 9.3005
R622 VTAIL.n821 VTAIL.n820 9.3005
R623 VTAIL.n819 VTAIL.n818 9.3005
R624 VTAIL.n800 VTAIL.n799 9.3005
R625 VTAIL.n813 VTAIL.n812 9.3005
R626 VTAIL.n811 VTAIL.n810 9.3005
R627 VTAIL.n804 VTAIL.n803 9.3005
R628 VTAIL.n829 VTAIL.n828 9.3005
R629 VTAIL.n792 VTAIL.n791 9.3005
R630 VTAIL.n835 VTAIL.n834 9.3005
R631 VTAIL.n837 VTAIL.n836 9.3005
R632 VTAIL.n788 VTAIL.n787 9.3005
R633 VTAIL.n843 VTAIL.n842 9.3005
R634 VTAIL.n845 VTAIL.n844 9.3005
R635 VTAIL.n846 VTAIL.n783 9.3005
R636 VTAIL.n853 VTAIL.n852 9.3005
R637 VTAIL.n772 VTAIL.n771 9.3005
R638 VTAIL.n107 VTAIL.n106 9.3005
R639 VTAIL.n101 VTAIL.n100 9.3005
R640 VTAIL.n99 VTAIL.n98 9.3005
R641 VTAIL.n6 VTAIL.n5 9.3005
R642 VTAIL.n93 VTAIL.n92 9.3005
R643 VTAIL.n91 VTAIL.n90 9.3005
R644 VTAIL.n10 VTAIL.n9 9.3005
R645 VTAIL.n85 VTAIL.n84 9.3005
R646 VTAIL.n57 VTAIL.n56 9.3005
R647 VTAIL.n26 VTAIL.n25 9.3005
R648 VTAIL.n51 VTAIL.n50 9.3005
R649 VTAIL.n49 VTAIL.n48 9.3005
R650 VTAIL.n30 VTAIL.n29 9.3005
R651 VTAIL.n43 VTAIL.n42 9.3005
R652 VTAIL.n41 VTAIL.n40 9.3005
R653 VTAIL.n34 VTAIL.n33 9.3005
R654 VTAIL.n59 VTAIL.n58 9.3005
R655 VTAIL.n22 VTAIL.n21 9.3005
R656 VTAIL.n65 VTAIL.n64 9.3005
R657 VTAIL.n67 VTAIL.n66 9.3005
R658 VTAIL.n18 VTAIL.n17 9.3005
R659 VTAIL.n73 VTAIL.n72 9.3005
R660 VTAIL.n75 VTAIL.n74 9.3005
R661 VTAIL.n76 VTAIL.n13 9.3005
R662 VTAIL.n83 VTAIL.n82 9.3005
R663 VTAIL.n2 VTAIL.n1 9.3005
R664 VTAIL.n217 VTAIL.n216 9.3005
R665 VTAIL.n211 VTAIL.n210 9.3005
R666 VTAIL.n209 VTAIL.n208 9.3005
R667 VTAIL.n116 VTAIL.n115 9.3005
R668 VTAIL.n203 VTAIL.n202 9.3005
R669 VTAIL.n201 VTAIL.n200 9.3005
R670 VTAIL.n120 VTAIL.n119 9.3005
R671 VTAIL.n195 VTAIL.n194 9.3005
R672 VTAIL.n167 VTAIL.n166 9.3005
R673 VTAIL.n136 VTAIL.n135 9.3005
R674 VTAIL.n161 VTAIL.n160 9.3005
R675 VTAIL.n159 VTAIL.n158 9.3005
R676 VTAIL.n140 VTAIL.n139 9.3005
R677 VTAIL.n153 VTAIL.n152 9.3005
R678 VTAIL.n151 VTAIL.n150 9.3005
R679 VTAIL.n144 VTAIL.n143 9.3005
R680 VTAIL.n169 VTAIL.n168 9.3005
R681 VTAIL.n132 VTAIL.n131 9.3005
R682 VTAIL.n175 VTAIL.n174 9.3005
R683 VTAIL.n177 VTAIL.n176 9.3005
R684 VTAIL.n128 VTAIL.n127 9.3005
R685 VTAIL.n183 VTAIL.n182 9.3005
R686 VTAIL.n185 VTAIL.n184 9.3005
R687 VTAIL.n186 VTAIL.n123 9.3005
R688 VTAIL.n193 VTAIL.n192 9.3005
R689 VTAIL.n112 VTAIL.n111 9.3005
R690 VTAIL.n327 VTAIL.n326 9.3005
R691 VTAIL.n321 VTAIL.n320 9.3005
R692 VTAIL.n319 VTAIL.n318 9.3005
R693 VTAIL.n226 VTAIL.n225 9.3005
R694 VTAIL.n313 VTAIL.n312 9.3005
R695 VTAIL.n311 VTAIL.n310 9.3005
R696 VTAIL.n230 VTAIL.n229 9.3005
R697 VTAIL.n305 VTAIL.n304 9.3005
R698 VTAIL.n277 VTAIL.n276 9.3005
R699 VTAIL.n246 VTAIL.n245 9.3005
R700 VTAIL.n271 VTAIL.n270 9.3005
R701 VTAIL.n269 VTAIL.n268 9.3005
R702 VTAIL.n250 VTAIL.n249 9.3005
R703 VTAIL.n263 VTAIL.n262 9.3005
R704 VTAIL.n261 VTAIL.n260 9.3005
R705 VTAIL.n254 VTAIL.n253 9.3005
R706 VTAIL.n279 VTAIL.n278 9.3005
R707 VTAIL.n242 VTAIL.n241 9.3005
R708 VTAIL.n285 VTAIL.n284 9.3005
R709 VTAIL.n287 VTAIL.n286 9.3005
R710 VTAIL.n238 VTAIL.n237 9.3005
R711 VTAIL.n293 VTAIL.n292 9.3005
R712 VTAIL.n295 VTAIL.n294 9.3005
R713 VTAIL.n296 VTAIL.n233 9.3005
R714 VTAIL.n303 VTAIL.n302 9.3005
R715 VTAIL.n222 VTAIL.n221 9.3005
R716 VTAIL.n684 VTAIL.n683 9.3005
R717 VTAIL.n727 VTAIL.n726 9.3005
R718 VTAIL.n729 VTAIL.n728 9.3005
R719 VTAIL.n680 VTAIL.n679 9.3005
R720 VTAIL.n735 VTAIL.n734 9.3005
R721 VTAIL.n737 VTAIL.n736 9.3005
R722 VTAIL.n675 VTAIL.n673 9.3005
R723 VTAIL.n743 VTAIL.n742 9.3005
R724 VTAIL.n767 VTAIL.n766 9.3005
R725 VTAIL.n662 VTAIL.n661 9.3005
R726 VTAIL.n761 VTAIL.n760 9.3005
R727 VTAIL.n759 VTAIL.n758 9.3005
R728 VTAIL.n666 VTAIL.n665 9.3005
R729 VTAIL.n753 VTAIL.n752 9.3005
R730 VTAIL.n751 VTAIL.n750 9.3005
R731 VTAIL.n670 VTAIL.n669 9.3005
R732 VTAIL.n745 VTAIL.n744 9.3005
R733 VTAIL.n721 VTAIL.n720 9.3005
R734 VTAIL.n719 VTAIL.n718 9.3005
R735 VTAIL.n688 VTAIL.n687 9.3005
R736 VTAIL.n713 VTAIL.n712 9.3005
R737 VTAIL.n711 VTAIL.n710 9.3005
R738 VTAIL.n692 VTAIL.n691 9.3005
R739 VTAIL.n705 VTAIL.n704 9.3005
R740 VTAIL.n703 VTAIL.n702 9.3005
R741 VTAIL.n696 VTAIL.n695 9.3005
R742 VTAIL.n574 VTAIL.n573 9.3005
R743 VTAIL.n617 VTAIL.n616 9.3005
R744 VTAIL.n619 VTAIL.n618 9.3005
R745 VTAIL.n570 VTAIL.n569 9.3005
R746 VTAIL.n625 VTAIL.n624 9.3005
R747 VTAIL.n627 VTAIL.n626 9.3005
R748 VTAIL.n565 VTAIL.n563 9.3005
R749 VTAIL.n633 VTAIL.n632 9.3005
R750 VTAIL.n657 VTAIL.n656 9.3005
R751 VTAIL.n552 VTAIL.n551 9.3005
R752 VTAIL.n651 VTAIL.n650 9.3005
R753 VTAIL.n649 VTAIL.n648 9.3005
R754 VTAIL.n556 VTAIL.n555 9.3005
R755 VTAIL.n643 VTAIL.n642 9.3005
R756 VTAIL.n641 VTAIL.n640 9.3005
R757 VTAIL.n560 VTAIL.n559 9.3005
R758 VTAIL.n635 VTAIL.n634 9.3005
R759 VTAIL.n611 VTAIL.n610 9.3005
R760 VTAIL.n609 VTAIL.n608 9.3005
R761 VTAIL.n578 VTAIL.n577 9.3005
R762 VTAIL.n603 VTAIL.n602 9.3005
R763 VTAIL.n601 VTAIL.n600 9.3005
R764 VTAIL.n582 VTAIL.n581 9.3005
R765 VTAIL.n595 VTAIL.n594 9.3005
R766 VTAIL.n593 VTAIL.n592 9.3005
R767 VTAIL.n586 VTAIL.n585 9.3005
R768 VTAIL.n464 VTAIL.n463 9.3005
R769 VTAIL.n507 VTAIL.n506 9.3005
R770 VTAIL.n509 VTAIL.n508 9.3005
R771 VTAIL.n460 VTAIL.n459 9.3005
R772 VTAIL.n515 VTAIL.n514 9.3005
R773 VTAIL.n517 VTAIL.n516 9.3005
R774 VTAIL.n455 VTAIL.n453 9.3005
R775 VTAIL.n523 VTAIL.n522 9.3005
R776 VTAIL.n547 VTAIL.n546 9.3005
R777 VTAIL.n442 VTAIL.n441 9.3005
R778 VTAIL.n541 VTAIL.n540 9.3005
R779 VTAIL.n539 VTAIL.n538 9.3005
R780 VTAIL.n446 VTAIL.n445 9.3005
R781 VTAIL.n533 VTAIL.n532 9.3005
R782 VTAIL.n531 VTAIL.n530 9.3005
R783 VTAIL.n450 VTAIL.n449 9.3005
R784 VTAIL.n525 VTAIL.n524 9.3005
R785 VTAIL.n501 VTAIL.n500 9.3005
R786 VTAIL.n499 VTAIL.n498 9.3005
R787 VTAIL.n468 VTAIL.n467 9.3005
R788 VTAIL.n493 VTAIL.n492 9.3005
R789 VTAIL.n491 VTAIL.n490 9.3005
R790 VTAIL.n472 VTAIL.n471 9.3005
R791 VTAIL.n485 VTAIL.n484 9.3005
R792 VTAIL.n483 VTAIL.n482 9.3005
R793 VTAIL.n476 VTAIL.n475 9.3005
R794 VTAIL.n354 VTAIL.n353 9.3005
R795 VTAIL.n397 VTAIL.n396 9.3005
R796 VTAIL.n399 VTAIL.n398 9.3005
R797 VTAIL.n350 VTAIL.n349 9.3005
R798 VTAIL.n405 VTAIL.n404 9.3005
R799 VTAIL.n407 VTAIL.n406 9.3005
R800 VTAIL.n345 VTAIL.n343 9.3005
R801 VTAIL.n413 VTAIL.n412 9.3005
R802 VTAIL.n437 VTAIL.n436 9.3005
R803 VTAIL.n332 VTAIL.n331 9.3005
R804 VTAIL.n431 VTAIL.n430 9.3005
R805 VTAIL.n429 VTAIL.n428 9.3005
R806 VTAIL.n336 VTAIL.n335 9.3005
R807 VTAIL.n423 VTAIL.n422 9.3005
R808 VTAIL.n421 VTAIL.n420 9.3005
R809 VTAIL.n340 VTAIL.n339 9.3005
R810 VTAIL.n415 VTAIL.n414 9.3005
R811 VTAIL.n391 VTAIL.n390 9.3005
R812 VTAIL.n389 VTAIL.n388 9.3005
R813 VTAIL.n358 VTAIL.n357 9.3005
R814 VTAIL.n383 VTAIL.n382 9.3005
R815 VTAIL.n381 VTAIL.n380 9.3005
R816 VTAIL.n362 VTAIL.n361 9.3005
R817 VTAIL.n375 VTAIL.n374 9.3005
R818 VTAIL.n373 VTAIL.n372 9.3005
R819 VTAIL.n366 VTAIL.n365 9.3005
R820 VTAIL.n822 VTAIL.n821 8.92171
R821 VTAIL.n837 VTAIL.n790 8.92171
R822 VTAIL.n868 VTAIL.n774 8.92171
R823 VTAIL.n52 VTAIL.n51 8.92171
R824 VTAIL.n67 VTAIL.n20 8.92171
R825 VTAIL.n98 VTAIL.n4 8.92171
R826 VTAIL.n162 VTAIL.n161 8.92171
R827 VTAIL.n177 VTAIL.n130 8.92171
R828 VTAIL.n208 VTAIL.n114 8.92171
R829 VTAIL.n272 VTAIL.n271 8.92171
R830 VTAIL.n287 VTAIL.n240 8.92171
R831 VTAIL.n318 VTAIL.n224 8.92171
R832 VTAIL.n758 VTAIL.n664 8.92171
R833 VTAIL.n729 VTAIL.n682 8.92171
R834 VTAIL.n714 VTAIL.n713 8.92171
R835 VTAIL.n648 VTAIL.n554 8.92171
R836 VTAIL.n619 VTAIL.n572 8.92171
R837 VTAIL.n604 VTAIL.n603 8.92171
R838 VTAIL.n538 VTAIL.n444 8.92171
R839 VTAIL.n509 VTAIL.n462 8.92171
R840 VTAIL.n494 VTAIL.n493 8.92171
R841 VTAIL.n428 VTAIL.n334 8.92171
R842 VTAIL.n399 VTAIL.n352 8.92171
R843 VTAIL.n384 VTAIL.n383 8.92171
R844 VTAIL.n825 VTAIL.n796 8.14595
R845 VTAIL.n834 VTAIL.n833 8.14595
R846 VTAIL.n872 VTAIL.n871 8.14595
R847 VTAIL.n55 VTAIL.n26 8.14595
R848 VTAIL.n64 VTAIL.n63 8.14595
R849 VTAIL.n102 VTAIL.n101 8.14595
R850 VTAIL.n165 VTAIL.n136 8.14595
R851 VTAIL.n174 VTAIL.n173 8.14595
R852 VTAIL.n212 VTAIL.n211 8.14595
R853 VTAIL.n275 VTAIL.n246 8.14595
R854 VTAIL.n284 VTAIL.n283 8.14595
R855 VTAIL.n322 VTAIL.n321 8.14595
R856 VTAIL.n762 VTAIL.n761 8.14595
R857 VTAIL.n726 VTAIL.n725 8.14595
R858 VTAIL.n717 VTAIL.n688 8.14595
R859 VTAIL.n652 VTAIL.n651 8.14595
R860 VTAIL.n616 VTAIL.n615 8.14595
R861 VTAIL.n607 VTAIL.n578 8.14595
R862 VTAIL.n542 VTAIL.n541 8.14595
R863 VTAIL.n506 VTAIL.n505 8.14595
R864 VTAIL.n497 VTAIL.n468 8.14595
R865 VTAIL.n432 VTAIL.n431 8.14595
R866 VTAIL.n396 VTAIL.n395 8.14595
R867 VTAIL.n387 VTAIL.n358 8.14595
R868 VTAIL.n826 VTAIL.n794 7.3702
R869 VTAIL.n830 VTAIL.n792 7.3702
R870 VTAIL.n875 VTAIL.n772 7.3702
R871 VTAIL.n878 VTAIL.n770 7.3702
R872 VTAIL.n56 VTAIL.n24 7.3702
R873 VTAIL.n60 VTAIL.n22 7.3702
R874 VTAIL.n105 VTAIL.n2 7.3702
R875 VTAIL.n108 VTAIL.n0 7.3702
R876 VTAIL.n166 VTAIL.n134 7.3702
R877 VTAIL.n170 VTAIL.n132 7.3702
R878 VTAIL.n215 VTAIL.n112 7.3702
R879 VTAIL.n218 VTAIL.n110 7.3702
R880 VTAIL.n276 VTAIL.n244 7.3702
R881 VTAIL.n280 VTAIL.n242 7.3702
R882 VTAIL.n325 VTAIL.n222 7.3702
R883 VTAIL.n328 VTAIL.n220 7.3702
R884 VTAIL.n768 VTAIL.n660 7.3702
R885 VTAIL.n765 VTAIL.n662 7.3702
R886 VTAIL.n722 VTAIL.n684 7.3702
R887 VTAIL.n718 VTAIL.n686 7.3702
R888 VTAIL.n658 VTAIL.n550 7.3702
R889 VTAIL.n655 VTAIL.n552 7.3702
R890 VTAIL.n612 VTAIL.n574 7.3702
R891 VTAIL.n608 VTAIL.n576 7.3702
R892 VTAIL.n548 VTAIL.n440 7.3702
R893 VTAIL.n545 VTAIL.n442 7.3702
R894 VTAIL.n502 VTAIL.n464 7.3702
R895 VTAIL.n498 VTAIL.n466 7.3702
R896 VTAIL.n438 VTAIL.n330 7.3702
R897 VTAIL.n435 VTAIL.n332 7.3702
R898 VTAIL.n392 VTAIL.n354 7.3702
R899 VTAIL.n388 VTAIL.n356 7.3702
R900 VTAIL.n829 VTAIL.n794 6.59444
R901 VTAIL.n830 VTAIL.n829 6.59444
R902 VTAIL.n876 VTAIL.n875 6.59444
R903 VTAIL.n876 VTAIL.n770 6.59444
R904 VTAIL.n59 VTAIL.n24 6.59444
R905 VTAIL.n60 VTAIL.n59 6.59444
R906 VTAIL.n106 VTAIL.n105 6.59444
R907 VTAIL.n106 VTAIL.n0 6.59444
R908 VTAIL.n169 VTAIL.n134 6.59444
R909 VTAIL.n170 VTAIL.n169 6.59444
R910 VTAIL.n216 VTAIL.n215 6.59444
R911 VTAIL.n216 VTAIL.n110 6.59444
R912 VTAIL.n279 VTAIL.n244 6.59444
R913 VTAIL.n280 VTAIL.n279 6.59444
R914 VTAIL.n326 VTAIL.n325 6.59444
R915 VTAIL.n326 VTAIL.n220 6.59444
R916 VTAIL.n766 VTAIL.n660 6.59444
R917 VTAIL.n766 VTAIL.n765 6.59444
R918 VTAIL.n722 VTAIL.n721 6.59444
R919 VTAIL.n721 VTAIL.n686 6.59444
R920 VTAIL.n656 VTAIL.n550 6.59444
R921 VTAIL.n656 VTAIL.n655 6.59444
R922 VTAIL.n612 VTAIL.n611 6.59444
R923 VTAIL.n611 VTAIL.n576 6.59444
R924 VTAIL.n546 VTAIL.n440 6.59444
R925 VTAIL.n546 VTAIL.n545 6.59444
R926 VTAIL.n502 VTAIL.n501 6.59444
R927 VTAIL.n501 VTAIL.n466 6.59444
R928 VTAIL.n436 VTAIL.n330 6.59444
R929 VTAIL.n436 VTAIL.n435 6.59444
R930 VTAIL.n392 VTAIL.n391 6.59444
R931 VTAIL.n391 VTAIL.n356 6.59444
R932 VTAIL.n826 VTAIL.n825 5.81868
R933 VTAIL.n833 VTAIL.n792 5.81868
R934 VTAIL.n872 VTAIL.n772 5.81868
R935 VTAIL.n56 VTAIL.n55 5.81868
R936 VTAIL.n63 VTAIL.n22 5.81868
R937 VTAIL.n102 VTAIL.n2 5.81868
R938 VTAIL.n166 VTAIL.n165 5.81868
R939 VTAIL.n173 VTAIL.n132 5.81868
R940 VTAIL.n212 VTAIL.n112 5.81868
R941 VTAIL.n276 VTAIL.n275 5.81868
R942 VTAIL.n283 VTAIL.n242 5.81868
R943 VTAIL.n322 VTAIL.n222 5.81868
R944 VTAIL.n762 VTAIL.n662 5.81868
R945 VTAIL.n725 VTAIL.n684 5.81868
R946 VTAIL.n718 VTAIL.n717 5.81868
R947 VTAIL.n652 VTAIL.n552 5.81868
R948 VTAIL.n615 VTAIL.n574 5.81868
R949 VTAIL.n608 VTAIL.n607 5.81868
R950 VTAIL.n542 VTAIL.n442 5.81868
R951 VTAIL.n505 VTAIL.n464 5.81868
R952 VTAIL.n498 VTAIL.n497 5.81868
R953 VTAIL.n432 VTAIL.n332 5.81868
R954 VTAIL.n395 VTAIL.n354 5.81868
R955 VTAIL.n388 VTAIL.n387 5.81868
R956 VTAIL.n822 VTAIL.n796 5.04292
R957 VTAIL.n834 VTAIL.n790 5.04292
R958 VTAIL.n871 VTAIL.n774 5.04292
R959 VTAIL.n52 VTAIL.n26 5.04292
R960 VTAIL.n64 VTAIL.n20 5.04292
R961 VTAIL.n101 VTAIL.n4 5.04292
R962 VTAIL.n162 VTAIL.n136 5.04292
R963 VTAIL.n174 VTAIL.n130 5.04292
R964 VTAIL.n211 VTAIL.n114 5.04292
R965 VTAIL.n272 VTAIL.n246 5.04292
R966 VTAIL.n284 VTAIL.n240 5.04292
R967 VTAIL.n321 VTAIL.n224 5.04292
R968 VTAIL.n761 VTAIL.n664 5.04292
R969 VTAIL.n726 VTAIL.n682 5.04292
R970 VTAIL.n714 VTAIL.n688 5.04292
R971 VTAIL.n651 VTAIL.n554 5.04292
R972 VTAIL.n616 VTAIL.n572 5.04292
R973 VTAIL.n604 VTAIL.n578 5.04292
R974 VTAIL.n541 VTAIL.n444 5.04292
R975 VTAIL.n506 VTAIL.n462 5.04292
R976 VTAIL.n494 VTAIL.n468 5.04292
R977 VTAIL.n431 VTAIL.n334 5.04292
R978 VTAIL.n396 VTAIL.n352 5.04292
R979 VTAIL.n384 VTAIL.n358 5.04292
R980 VTAIL.n821 VTAIL.n798 4.26717
R981 VTAIL.n838 VTAIL.n837 4.26717
R982 VTAIL.n868 VTAIL.n867 4.26717
R983 VTAIL.n51 VTAIL.n28 4.26717
R984 VTAIL.n68 VTAIL.n67 4.26717
R985 VTAIL.n98 VTAIL.n97 4.26717
R986 VTAIL.n161 VTAIL.n138 4.26717
R987 VTAIL.n178 VTAIL.n177 4.26717
R988 VTAIL.n208 VTAIL.n207 4.26717
R989 VTAIL.n271 VTAIL.n248 4.26717
R990 VTAIL.n288 VTAIL.n287 4.26717
R991 VTAIL.n318 VTAIL.n317 4.26717
R992 VTAIL.n758 VTAIL.n757 4.26717
R993 VTAIL.n730 VTAIL.n729 4.26717
R994 VTAIL.n713 VTAIL.n690 4.26717
R995 VTAIL.n648 VTAIL.n647 4.26717
R996 VTAIL.n620 VTAIL.n619 4.26717
R997 VTAIL.n603 VTAIL.n580 4.26717
R998 VTAIL.n538 VTAIL.n537 4.26717
R999 VTAIL.n510 VTAIL.n509 4.26717
R1000 VTAIL.n493 VTAIL.n470 4.26717
R1001 VTAIL.n428 VTAIL.n427 4.26717
R1002 VTAIL.n400 VTAIL.n399 4.26717
R1003 VTAIL.n383 VTAIL.n360 4.26717
R1004 VTAIL.n805 VTAIL.n803 3.70982
R1005 VTAIL.n35 VTAIL.n33 3.70982
R1006 VTAIL.n145 VTAIL.n143 3.70982
R1007 VTAIL.n255 VTAIL.n253 3.70982
R1008 VTAIL.n697 VTAIL.n695 3.70982
R1009 VTAIL.n587 VTAIL.n585 3.70982
R1010 VTAIL.n477 VTAIL.n475 3.70982
R1011 VTAIL.n367 VTAIL.n365 3.70982
R1012 VTAIL.n818 VTAIL.n817 3.49141
R1013 VTAIL.n841 VTAIL.n788 3.49141
R1014 VTAIL.n864 VTAIL.n776 3.49141
R1015 VTAIL.n48 VTAIL.n47 3.49141
R1016 VTAIL.n71 VTAIL.n18 3.49141
R1017 VTAIL.n94 VTAIL.n6 3.49141
R1018 VTAIL.n158 VTAIL.n157 3.49141
R1019 VTAIL.n181 VTAIL.n128 3.49141
R1020 VTAIL.n204 VTAIL.n116 3.49141
R1021 VTAIL.n268 VTAIL.n267 3.49141
R1022 VTAIL.n291 VTAIL.n238 3.49141
R1023 VTAIL.n314 VTAIL.n226 3.49141
R1024 VTAIL.n754 VTAIL.n666 3.49141
R1025 VTAIL.n733 VTAIL.n680 3.49141
R1026 VTAIL.n710 VTAIL.n709 3.49141
R1027 VTAIL.n644 VTAIL.n556 3.49141
R1028 VTAIL.n623 VTAIL.n570 3.49141
R1029 VTAIL.n600 VTAIL.n599 3.49141
R1030 VTAIL.n534 VTAIL.n446 3.49141
R1031 VTAIL.n513 VTAIL.n460 3.49141
R1032 VTAIL.n490 VTAIL.n489 3.49141
R1033 VTAIL.n424 VTAIL.n336 3.49141
R1034 VTAIL.n403 VTAIL.n350 3.49141
R1035 VTAIL.n380 VTAIL.n379 3.49141
R1036 VTAIL.n814 VTAIL.n800 2.71565
R1037 VTAIL.n842 VTAIL.n786 2.71565
R1038 VTAIL.n863 VTAIL.n778 2.71565
R1039 VTAIL.n44 VTAIL.n30 2.71565
R1040 VTAIL.n72 VTAIL.n16 2.71565
R1041 VTAIL.n93 VTAIL.n8 2.71565
R1042 VTAIL.n154 VTAIL.n140 2.71565
R1043 VTAIL.n182 VTAIL.n126 2.71565
R1044 VTAIL.n203 VTAIL.n118 2.71565
R1045 VTAIL.n264 VTAIL.n250 2.71565
R1046 VTAIL.n292 VTAIL.n236 2.71565
R1047 VTAIL.n313 VTAIL.n228 2.71565
R1048 VTAIL.n753 VTAIL.n668 2.71565
R1049 VTAIL.n734 VTAIL.n678 2.71565
R1050 VTAIL.n706 VTAIL.n692 2.71565
R1051 VTAIL.n643 VTAIL.n558 2.71565
R1052 VTAIL.n624 VTAIL.n568 2.71565
R1053 VTAIL.n596 VTAIL.n582 2.71565
R1054 VTAIL.n533 VTAIL.n448 2.71565
R1055 VTAIL.n514 VTAIL.n458 2.71565
R1056 VTAIL.n486 VTAIL.n472 2.71565
R1057 VTAIL.n423 VTAIL.n338 2.71565
R1058 VTAIL.n404 VTAIL.n348 2.71565
R1059 VTAIL.n376 VTAIL.n362 2.71565
R1060 VTAIL.n813 VTAIL.n802 1.93989
R1061 VTAIL.n847 VTAIL.n845 1.93989
R1062 VTAIL.n860 VTAIL.n859 1.93989
R1063 VTAIL.n43 VTAIL.n32 1.93989
R1064 VTAIL.n77 VTAIL.n75 1.93989
R1065 VTAIL.n90 VTAIL.n89 1.93989
R1066 VTAIL.n153 VTAIL.n142 1.93989
R1067 VTAIL.n187 VTAIL.n185 1.93989
R1068 VTAIL.n200 VTAIL.n199 1.93989
R1069 VTAIL.n263 VTAIL.n252 1.93989
R1070 VTAIL.n297 VTAIL.n295 1.93989
R1071 VTAIL.n310 VTAIL.n309 1.93989
R1072 VTAIL.n750 VTAIL.n749 1.93989
R1073 VTAIL.n738 VTAIL.n737 1.93989
R1074 VTAIL.n705 VTAIL.n694 1.93989
R1075 VTAIL.n640 VTAIL.n639 1.93989
R1076 VTAIL.n628 VTAIL.n627 1.93989
R1077 VTAIL.n595 VTAIL.n584 1.93989
R1078 VTAIL.n530 VTAIL.n529 1.93989
R1079 VTAIL.n518 VTAIL.n517 1.93989
R1080 VTAIL.n485 VTAIL.n474 1.93989
R1081 VTAIL.n420 VTAIL.n419 1.93989
R1082 VTAIL.n408 VTAIL.n407 1.93989
R1083 VTAIL.n375 VTAIL.n364 1.93989
R1084 VTAIL.n810 VTAIL.n809 1.16414
R1085 VTAIL.n846 VTAIL.n784 1.16414
R1086 VTAIL.n856 VTAIL.n780 1.16414
R1087 VTAIL.n40 VTAIL.n39 1.16414
R1088 VTAIL.n76 VTAIL.n14 1.16414
R1089 VTAIL.n86 VTAIL.n10 1.16414
R1090 VTAIL.n150 VTAIL.n149 1.16414
R1091 VTAIL.n186 VTAIL.n124 1.16414
R1092 VTAIL.n196 VTAIL.n120 1.16414
R1093 VTAIL.n260 VTAIL.n259 1.16414
R1094 VTAIL.n296 VTAIL.n234 1.16414
R1095 VTAIL.n306 VTAIL.n230 1.16414
R1096 VTAIL.n746 VTAIL.n670 1.16414
R1097 VTAIL.n741 VTAIL.n675 1.16414
R1098 VTAIL.n702 VTAIL.n701 1.16414
R1099 VTAIL.n636 VTAIL.n560 1.16414
R1100 VTAIL.n631 VTAIL.n565 1.16414
R1101 VTAIL.n592 VTAIL.n591 1.16414
R1102 VTAIL.n526 VTAIL.n450 1.16414
R1103 VTAIL.n521 VTAIL.n455 1.16414
R1104 VTAIL.n482 VTAIL.n481 1.16414
R1105 VTAIL.n416 VTAIL.n340 1.16414
R1106 VTAIL.n411 VTAIL.n345 1.16414
R1107 VTAIL.n372 VTAIL.n371 1.16414
R1108 VTAIL.n549 VTAIL.n439 0.664293
R1109 VTAIL.n769 VTAIL.n659 0.664293
R1110 VTAIL.n329 VTAIL.n219 0.664293
R1111 VTAIL.n659 VTAIL.n549 0.470328
R1112 VTAIL.n219 VTAIL.n109 0.470328
R1113 VTAIL VTAIL.n109 0.390586
R1114 VTAIL.n806 VTAIL.n804 0.388379
R1115 VTAIL.n852 VTAIL.n851 0.388379
R1116 VTAIL.n855 VTAIL.n782 0.388379
R1117 VTAIL.n36 VTAIL.n34 0.388379
R1118 VTAIL.n82 VTAIL.n81 0.388379
R1119 VTAIL.n85 VTAIL.n12 0.388379
R1120 VTAIL.n146 VTAIL.n144 0.388379
R1121 VTAIL.n192 VTAIL.n191 0.388379
R1122 VTAIL.n195 VTAIL.n122 0.388379
R1123 VTAIL.n256 VTAIL.n254 0.388379
R1124 VTAIL.n302 VTAIL.n301 0.388379
R1125 VTAIL.n305 VTAIL.n232 0.388379
R1126 VTAIL.n745 VTAIL.n672 0.388379
R1127 VTAIL.n742 VTAIL.n674 0.388379
R1128 VTAIL.n698 VTAIL.n696 0.388379
R1129 VTAIL.n635 VTAIL.n562 0.388379
R1130 VTAIL.n632 VTAIL.n564 0.388379
R1131 VTAIL.n588 VTAIL.n586 0.388379
R1132 VTAIL.n525 VTAIL.n452 0.388379
R1133 VTAIL.n522 VTAIL.n454 0.388379
R1134 VTAIL.n478 VTAIL.n476 0.388379
R1135 VTAIL.n415 VTAIL.n342 0.388379
R1136 VTAIL.n412 VTAIL.n344 0.388379
R1137 VTAIL.n368 VTAIL.n366 0.388379
R1138 VTAIL VTAIL.n879 0.274207
R1139 VTAIL.n811 VTAIL.n803 0.155672
R1140 VTAIL.n812 VTAIL.n811 0.155672
R1141 VTAIL.n812 VTAIL.n799 0.155672
R1142 VTAIL.n819 VTAIL.n799 0.155672
R1143 VTAIL.n820 VTAIL.n819 0.155672
R1144 VTAIL.n820 VTAIL.n795 0.155672
R1145 VTAIL.n827 VTAIL.n795 0.155672
R1146 VTAIL.n828 VTAIL.n827 0.155672
R1147 VTAIL.n828 VTAIL.n791 0.155672
R1148 VTAIL.n835 VTAIL.n791 0.155672
R1149 VTAIL.n836 VTAIL.n835 0.155672
R1150 VTAIL.n836 VTAIL.n787 0.155672
R1151 VTAIL.n843 VTAIL.n787 0.155672
R1152 VTAIL.n844 VTAIL.n843 0.155672
R1153 VTAIL.n844 VTAIL.n783 0.155672
R1154 VTAIL.n853 VTAIL.n783 0.155672
R1155 VTAIL.n854 VTAIL.n853 0.155672
R1156 VTAIL.n854 VTAIL.n779 0.155672
R1157 VTAIL.n861 VTAIL.n779 0.155672
R1158 VTAIL.n862 VTAIL.n861 0.155672
R1159 VTAIL.n862 VTAIL.n775 0.155672
R1160 VTAIL.n869 VTAIL.n775 0.155672
R1161 VTAIL.n870 VTAIL.n869 0.155672
R1162 VTAIL.n870 VTAIL.n771 0.155672
R1163 VTAIL.n877 VTAIL.n771 0.155672
R1164 VTAIL.n41 VTAIL.n33 0.155672
R1165 VTAIL.n42 VTAIL.n41 0.155672
R1166 VTAIL.n42 VTAIL.n29 0.155672
R1167 VTAIL.n49 VTAIL.n29 0.155672
R1168 VTAIL.n50 VTAIL.n49 0.155672
R1169 VTAIL.n50 VTAIL.n25 0.155672
R1170 VTAIL.n57 VTAIL.n25 0.155672
R1171 VTAIL.n58 VTAIL.n57 0.155672
R1172 VTAIL.n58 VTAIL.n21 0.155672
R1173 VTAIL.n65 VTAIL.n21 0.155672
R1174 VTAIL.n66 VTAIL.n65 0.155672
R1175 VTAIL.n66 VTAIL.n17 0.155672
R1176 VTAIL.n73 VTAIL.n17 0.155672
R1177 VTAIL.n74 VTAIL.n73 0.155672
R1178 VTAIL.n74 VTAIL.n13 0.155672
R1179 VTAIL.n83 VTAIL.n13 0.155672
R1180 VTAIL.n84 VTAIL.n83 0.155672
R1181 VTAIL.n84 VTAIL.n9 0.155672
R1182 VTAIL.n91 VTAIL.n9 0.155672
R1183 VTAIL.n92 VTAIL.n91 0.155672
R1184 VTAIL.n92 VTAIL.n5 0.155672
R1185 VTAIL.n99 VTAIL.n5 0.155672
R1186 VTAIL.n100 VTAIL.n99 0.155672
R1187 VTAIL.n100 VTAIL.n1 0.155672
R1188 VTAIL.n107 VTAIL.n1 0.155672
R1189 VTAIL.n151 VTAIL.n143 0.155672
R1190 VTAIL.n152 VTAIL.n151 0.155672
R1191 VTAIL.n152 VTAIL.n139 0.155672
R1192 VTAIL.n159 VTAIL.n139 0.155672
R1193 VTAIL.n160 VTAIL.n159 0.155672
R1194 VTAIL.n160 VTAIL.n135 0.155672
R1195 VTAIL.n167 VTAIL.n135 0.155672
R1196 VTAIL.n168 VTAIL.n167 0.155672
R1197 VTAIL.n168 VTAIL.n131 0.155672
R1198 VTAIL.n175 VTAIL.n131 0.155672
R1199 VTAIL.n176 VTAIL.n175 0.155672
R1200 VTAIL.n176 VTAIL.n127 0.155672
R1201 VTAIL.n183 VTAIL.n127 0.155672
R1202 VTAIL.n184 VTAIL.n183 0.155672
R1203 VTAIL.n184 VTAIL.n123 0.155672
R1204 VTAIL.n193 VTAIL.n123 0.155672
R1205 VTAIL.n194 VTAIL.n193 0.155672
R1206 VTAIL.n194 VTAIL.n119 0.155672
R1207 VTAIL.n201 VTAIL.n119 0.155672
R1208 VTAIL.n202 VTAIL.n201 0.155672
R1209 VTAIL.n202 VTAIL.n115 0.155672
R1210 VTAIL.n209 VTAIL.n115 0.155672
R1211 VTAIL.n210 VTAIL.n209 0.155672
R1212 VTAIL.n210 VTAIL.n111 0.155672
R1213 VTAIL.n217 VTAIL.n111 0.155672
R1214 VTAIL.n261 VTAIL.n253 0.155672
R1215 VTAIL.n262 VTAIL.n261 0.155672
R1216 VTAIL.n262 VTAIL.n249 0.155672
R1217 VTAIL.n269 VTAIL.n249 0.155672
R1218 VTAIL.n270 VTAIL.n269 0.155672
R1219 VTAIL.n270 VTAIL.n245 0.155672
R1220 VTAIL.n277 VTAIL.n245 0.155672
R1221 VTAIL.n278 VTAIL.n277 0.155672
R1222 VTAIL.n278 VTAIL.n241 0.155672
R1223 VTAIL.n285 VTAIL.n241 0.155672
R1224 VTAIL.n286 VTAIL.n285 0.155672
R1225 VTAIL.n286 VTAIL.n237 0.155672
R1226 VTAIL.n293 VTAIL.n237 0.155672
R1227 VTAIL.n294 VTAIL.n293 0.155672
R1228 VTAIL.n294 VTAIL.n233 0.155672
R1229 VTAIL.n303 VTAIL.n233 0.155672
R1230 VTAIL.n304 VTAIL.n303 0.155672
R1231 VTAIL.n304 VTAIL.n229 0.155672
R1232 VTAIL.n311 VTAIL.n229 0.155672
R1233 VTAIL.n312 VTAIL.n311 0.155672
R1234 VTAIL.n312 VTAIL.n225 0.155672
R1235 VTAIL.n319 VTAIL.n225 0.155672
R1236 VTAIL.n320 VTAIL.n319 0.155672
R1237 VTAIL.n320 VTAIL.n221 0.155672
R1238 VTAIL.n327 VTAIL.n221 0.155672
R1239 VTAIL.n767 VTAIL.n661 0.155672
R1240 VTAIL.n760 VTAIL.n661 0.155672
R1241 VTAIL.n760 VTAIL.n759 0.155672
R1242 VTAIL.n759 VTAIL.n665 0.155672
R1243 VTAIL.n752 VTAIL.n665 0.155672
R1244 VTAIL.n752 VTAIL.n751 0.155672
R1245 VTAIL.n751 VTAIL.n669 0.155672
R1246 VTAIL.n744 VTAIL.n669 0.155672
R1247 VTAIL.n744 VTAIL.n743 0.155672
R1248 VTAIL.n743 VTAIL.n673 0.155672
R1249 VTAIL.n736 VTAIL.n673 0.155672
R1250 VTAIL.n736 VTAIL.n735 0.155672
R1251 VTAIL.n735 VTAIL.n679 0.155672
R1252 VTAIL.n728 VTAIL.n679 0.155672
R1253 VTAIL.n728 VTAIL.n727 0.155672
R1254 VTAIL.n727 VTAIL.n683 0.155672
R1255 VTAIL.n720 VTAIL.n683 0.155672
R1256 VTAIL.n720 VTAIL.n719 0.155672
R1257 VTAIL.n719 VTAIL.n687 0.155672
R1258 VTAIL.n712 VTAIL.n687 0.155672
R1259 VTAIL.n712 VTAIL.n711 0.155672
R1260 VTAIL.n711 VTAIL.n691 0.155672
R1261 VTAIL.n704 VTAIL.n691 0.155672
R1262 VTAIL.n704 VTAIL.n703 0.155672
R1263 VTAIL.n703 VTAIL.n695 0.155672
R1264 VTAIL.n657 VTAIL.n551 0.155672
R1265 VTAIL.n650 VTAIL.n551 0.155672
R1266 VTAIL.n650 VTAIL.n649 0.155672
R1267 VTAIL.n649 VTAIL.n555 0.155672
R1268 VTAIL.n642 VTAIL.n555 0.155672
R1269 VTAIL.n642 VTAIL.n641 0.155672
R1270 VTAIL.n641 VTAIL.n559 0.155672
R1271 VTAIL.n634 VTAIL.n559 0.155672
R1272 VTAIL.n634 VTAIL.n633 0.155672
R1273 VTAIL.n633 VTAIL.n563 0.155672
R1274 VTAIL.n626 VTAIL.n563 0.155672
R1275 VTAIL.n626 VTAIL.n625 0.155672
R1276 VTAIL.n625 VTAIL.n569 0.155672
R1277 VTAIL.n618 VTAIL.n569 0.155672
R1278 VTAIL.n618 VTAIL.n617 0.155672
R1279 VTAIL.n617 VTAIL.n573 0.155672
R1280 VTAIL.n610 VTAIL.n573 0.155672
R1281 VTAIL.n610 VTAIL.n609 0.155672
R1282 VTAIL.n609 VTAIL.n577 0.155672
R1283 VTAIL.n602 VTAIL.n577 0.155672
R1284 VTAIL.n602 VTAIL.n601 0.155672
R1285 VTAIL.n601 VTAIL.n581 0.155672
R1286 VTAIL.n594 VTAIL.n581 0.155672
R1287 VTAIL.n594 VTAIL.n593 0.155672
R1288 VTAIL.n593 VTAIL.n585 0.155672
R1289 VTAIL.n547 VTAIL.n441 0.155672
R1290 VTAIL.n540 VTAIL.n441 0.155672
R1291 VTAIL.n540 VTAIL.n539 0.155672
R1292 VTAIL.n539 VTAIL.n445 0.155672
R1293 VTAIL.n532 VTAIL.n445 0.155672
R1294 VTAIL.n532 VTAIL.n531 0.155672
R1295 VTAIL.n531 VTAIL.n449 0.155672
R1296 VTAIL.n524 VTAIL.n449 0.155672
R1297 VTAIL.n524 VTAIL.n523 0.155672
R1298 VTAIL.n523 VTAIL.n453 0.155672
R1299 VTAIL.n516 VTAIL.n453 0.155672
R1300 VTAIL.n516 VTAIL.n515 0.155672
R1301 VTAIL.n515 VTAIL.n459 0.155672
R1302 VTAIL.n508 VTAIL.n459 0.155672
R1303 VTAIL.n508 VTAIL.n507 0.155672
R1304 VTAIL.n507 VTAIL.n463 0.155672
R1305 VTAIL.n500 VTAIL.n463 0.155672
R1306 VTAIL.n500 VTAIL.n499 0.155672
R1307 VTAIL.n499 VTAIL.n467 0.155672
R1308 VTAIL.n492 VTAIL.n467 0.155672
R1309 VTAIL.n492 VTAIL.n491 0.155672
R1310 VTAIL.n491 VTAIL.n471 0.155672
R1311 VTAIL.n484 VTAIL.n471 0.155672
R1312 VTAIL.n484 VTAIL.n483 0.155672
R1313 VTAIL.n483 VTAIL.n475 0.155672
R1314 VTAIL.n437 VTAIL.n331 0.155672
R1315 VTAIL.n430 VTAIL.n331 0.155672
R1316 VTAIL.n430 VTAIL.n429 0.155672
R1317 VTAIL.n429 VTAIL.n335 0.155672
R1318 VTAIL.n422 VTAIL.n335 0.155672
R1319 VTAIL.n422 VTAIL.n421 0.155672
R1320 VTAIL.n421 VTAIL.n339 0.155672
R1321 VTAIL.n414 VTAIL.n339 0.155672
R1322 VTAIL.n414 VTAIL.n413 0.155672
R1323 VTAIL.n413 VTAIL.n343 0.155672
R1324 VTAIL.n406 VTAIL.n343 0.155672
R1325 VTAIL.n406 VTAIL.n405 0.155672
R1326 VTAIL.n405 VTAIL.n349 0.155672
R1327 VTAIL.n398 VTAIL.n349 0.155672
R1328 VTAIL.n398 VTAIL.n397 0.155672
R1329 VTAIL.n397 VTAIL.n353 0.155672
R1330 VTAIL.n390 VTAIL.n353 0.155672
R1331 VTAIL.n390 VTAIL.n389 0.155672
R1332 VTAIL.n389 VTAIL.n357 0.155672
R1333 VTAIL.n382 VTAIL.n357 0.155672
R1334 VTAIL.n382 VTAIL.n381 0.155672
R1335 VTAIL.n381 VTAIL.n361 0.155672
R1336 VTAIL.n374 VTAIL.n361 0.155672
R1337 VTAIL.n374 VTAIL.n373 0.155672
R1338 VTAIL.n373 VTAIL.n365 0.155672
R1339 VDD1 VDD1.n1 110.293
R1340 VDD1 VDD1.n0 67.1981
R1341 VDD1.n0 VDD1.t0 1.65638
R1342 VDD1.n0 VDD1.t3 1.65638
R1343 VDD1.n1 VDD1.t2 1.65638
R1344 VDD1.n1 VDD1.t1 1.65638
R1345 VN.n0 VN.t3 1186
R1346 VN.n1 VN.t1 1186
R1347 VN.n0 VN.t0 1185.97
R1348 VN.n1 VN.t2 1185.97
R1349 VN VN.n1 115.989
R1350 VN VN.n0 70.265
R1351 VDD2.n2 VDD2.n0 109.769
R1352 VDD2.n2 VDD2.n1 67.1399
R1353 VDD2.n1 VDD2.t1 1.65638
R1354 VDD2.n1 VDD2.t2 1.65638
R1355 VDD2.n0 VDD2.t0 1.65638
R1356 VDD2.n0 VDD2.t3 1.65638
R1357 VDD2 VDD2.n2 0.0586897
R1358 B.n131 B.t6 1283.24
R1359 B.n139 B.t9 1283.24
R1360 B.n42 B.t0 1283.24
R1361 B.n50 B.t3 1283.24
R1362 B.n456 B.n83 585
R1363 B.n458 B.n457 585
R1364 B.n459 B.n82 585
R1365 B.n461 B.n460 585
R1366 B.n462 B.n81 585
R1367 B.n464 B.n463 585
R1368 B.n465 B.n80 585
R1369 B.n467 B.n466 585
R1370 B.n468 B.n79 585
R1371 B.n470 B.n469 585
R1372 B.n471 B.n78 585
R1373 B.n473 B.n472 585
R1374 B.n474 B.n77 585
R1375 B.n476 B.n475 585
R1376 B.n477 B.n76 585
R1377 B.n479 B.n478 585
R1378 B.n480 B.n75 585
R1379 B.n482 B.n481 585
R1380 B.n483 B.n74 585
R1381 B.n485 B.n484 585
R1382 B.n486 B.n73 585
R1383 B.n488 B.n487 585
R1384 B.n489 B.n72 585
R1385 B.n491 B.n490 585
R1386 B.n492 B.n71 585
R1387 B.n494 B.n493 585
R1388 B.n495 B.n70 585
R1389 B.n497 B.n496 585
R1390 B.n498 B.n69 585
R1391 B.n500 B.n499 585
R1392 B.n501 B.n68 585
R1393 B.n503 B.n502 585
R1394 B.n504 B.n67 585
R1395 B.n506 B.n505 585
R1396 B.n507 B.n66 585
R1397 B.n509 B.n508 585
R1398 B.n510 B.n65 585
R1399 B.n512 B.n511 585
R1400 B.n513 B.n64 585
R1401 B.n515 B.n514 585
R1402 B.n516 B.n63 585
R1403 B.n518 B.n517 585
R1404 B.n519 B.n62 585
R1405 B.n521 B.n520 585
R1406 B.n522 B.n61 585
R1407 B.n524 B.n523 585
R1408 B.n525 B.n60 585
R1409 B.n527 B.n526 585
R1410 B.n528 B.n59 585
R1411 B.n530 B.n529 585
R1412 B.n531 B.n58 585
R1413 B.n533 B.n532 585
R1414 B.n534 B.n57 585
R1415 B.n536 B.n535 585
R1416 B.n537 B.n56 585
R1417 B.n539 B.n538 585
R1418 B.n540 B.n55 585
R1419 B.n542 B.n541 585
R1420 B.n543 B.n54 585
R1421 B.n545 B.n544 585
R1422 B.n546 B.n53 585
R1423 B.n548 B.n547 585
R1424 B.n549 B.n49 585
R1425 B.n551 B.n550 585
R1426 B.n552 B.n48 585
R1427 B.n554 B.n553 585
R1428 B.n555 B.n47 585
R1429 B.n557 B.n556 585
R1430 B.n558 B.n46 585
R1431 B.n560 B.n559 585
R1432 B.n561 B.n45 585
R1433 B.n563 B.n562 585
R1434 B.n564 B.n44 585
R1435 B.n566 B.n565 585
R1436 B.n568 B.n41 585
R1437 B.n570 B.n569 585
R1438 B.n571 B.n40 585
R1439 B.n573 B.n572 585
R1440 B.n574 B.n39 585
R1441 B.n576 B.n575 585
R1442 B.n577 B.n38 585
R1443 B.n579 B.n578 585
R1444 B.n580 B.n37 585
R1445 B.n582 B.n581 585
R1446 B.n583 B.n36 585
R1447 B.n585 B.n584 585
R1448 B.n586 B.n35 585
R1449 B.n588 B.n587 585
R1450 B.n589 B.n34 585
R1451 B.n591 B.n590 585
R1452 B.n592 B.n33 585
R1453 B.n594 B.n593 585
R1454 B.n595 B.n32 585
R1455 B.n597 B.n596 585
R1456 B.n598 B.n31 585
R1457 B.n600 B.n599 585
R1458 B.n601 B.n30 585
R1459 B.n603 B.n602 585
R1460 B.n604 B.n29 585
R1461 B.n606 B.n605 585
R1462 B.n607 B.n28 585
R1463 B.n609 B.n608 585
R1464 B.n610 B.n27 585
R1465 B.n612 B.n611 585
R1466 B.n613 B.n26 585
R1467 B.n615 B.n614 585
R1468 B.n616 B.n25 585
R1469 B.n618 B.n617 585
R1470 B.n619 B.n24 585
R1471 B.n621 B.n620 585
R1472 B.n622 B.n23 585
R1473 B.n624 B.n623 585
R1474 B.n625 B.n22 585
R1475 B.n627 B.n626 585
R1476 B.n628 B.n21 585
R1477 B.n630 B.n629 585
R1478 B.n631 B.n20 585
R1479 B.n633 B.n632 585
R1480 B.n634 B.n19 585
R1481 B.n636 B.n635 585
R1482 B.n637 B.n18 585
R1483 B.n639 B.n638 585
R1484 B.n640 B.n17 585
R1485 B.n642 B.n641 585
R1486 B.n643 B.n16 585
R1487 B.n645 B.n644 585
R1488 B.n646 B.n15 585
R1489 B.n648 B.n647 585
R1490 B.n649 B.n14 585
R1491 B.n651 B.n650 585
R1492 B.n652 B.n13 585
R1493 B.n654 B.n653 585
R1494 B.n655 B.n12 585
R1495 B.n657 B.n656 585
R1496 B.n658 B.n11 585
R1497 B.n660 B.n659 585
R1498 B.n661 B.n10 585
R1499 B.n663 B.n662 585
R1500 B.n455 B.n454 585
R1501 B.n453 B.n84 585
R1502 B.n452 B.n451 585
R1503 B.n450 B.n85 585
R1504 B.n449 B.n448 585
R1505 B.n447 B.n86 585
R1506 B.n446 B.n445 585
R1507 B.n444 B.n87 585
R1508 B.n443 B.n442 585
R1509 B.n441 B.n88 585
R1510 B.n440 B.n439 585
R1511 B.n438 B.n89 585
R1512 B.n437 B.n436 585
R1513 B.n435 B.n90 585
R1514 B.n434 B.n433 585
R1515 B.n432 B.n91 585
R1516 B.n431 B.n430 585
R1517 B.n429 B.n92 585
R1518 B.n428 B.n427 585
R1519 B.n426 B.n93 585
R1520 B.n425 B.n424 585
R1521 B.n423 B.n94 585
R1522 B.n422 B.n421 585
R1523 B.n420 B.n95 585
R1524 B.n419 B.n418 585
R1525 B.n417 B.n96 585
R1526 B.n416 B.n415 585
R1527 B.n414 B.n97 585
R1528 B.n413 B.n412 585
R1529 B.n411 B.n98 585
R1530 B.n410 B.n409 585
R1531 B.n201 B.n172 585
R1532 B.n203 B.n202 585
R1533 B.n204 B.n171 585
R1534 B.n206 B.n205 585
R1535 B.n207 B.n170 585
R1536 B.n209 B.n208 585
R1537 B.n210 B.n169 585
R1538 B.n212 B.n211 585
R1539 B.n213 B.n168 585
R1540 B.n215 B.n214 585
R1541 B.n216 B.n167 585
R1542 B.n218 B.n217 585
R1543 B.n219 B.n166 585
R1544 B.n221 B.n220 585
R1545 B.n222 B.n165 585
R1546 B.n224 B.n223 585
R1547 B.n225 B.n164 585
R1548 B.n227 B.n226 585
R1549 B.n228 B.n163 585
R1550 B.n230 B.n229 585
R1551 B.n231 B.n162 585
R1552 B.n233 B.n232 585
R1553 B.n234 B.n161 585
R1554 B.n236 B.n235 585
R1555 B.n237 B.n160 585
R1556 B.n239 B.n238 585
R1557 B.n240 B.n159 585
R1558 B.n242 B.n241 585
R1559 B.n243 B.n158 585
R1560 B.n245 B.n244 585
R1561 B.n246 B.n157 585
R1562 B.n248 B.n247 585
R1563 B.n249 B.n156 585
R1564 B.n251 B.n250 585
R1565 B.n252 B.n155 585
R1566 B.n254 B.n253 585
R1567 B.n255 B.n154 585
R1568 B.n257 B.n256 585
R1569 B.n258 B.n153 585
R1570 B.n260 B.n259 585
R1571 B.n261 B.n152 585
R1572 B.n263 B.n262 585
R1573 B.n264 B.n151 585
R1574 B.n266 B.n265 585
R1575 B.n267 B.n150 585
R1576 B.n269 B.n268 585
R1577 B.n270 B.n149 585
R1578 B.n272 B.n271 585
R1579 B.n273 B.n148 585
R1580 B.n275 B.n274 585
R1581 B.n276 B.n147 585
R1582 B.n278 B.n277 585
R1583 B.n279 B.n146 585
R1584 B.n281 B.n280 585
R1585 B.n282 B.n145 585
R1586 B.n284 B.n283 585
R1587 B.n285 B.n144 585
R1588 B.n287 B.n286 585
R1589 B.n288 B.n143 585
R1590 B.n290 B.n289 585
R1591 B.n291 B.n142 585
R1592 B.n293 B.n292 585
R1593 B.n294 B.n141 585
R1594 B.n296 B.n295 585
R1595 B.n298 B.n138 585
R1596 B.n300 B.n299 585
R1597 B.n301 B.n137 585
R1598 B.n303 B.n302 585
R1599 B.n304 B.n136 585
R1600 B.n306 B.n305 585
R1601 B.n307 B.n135 585
R1602 B.n309 B.n308 585
R1603 B.n310 B.n134 585
R1604 B.n312 B.n311 585
R1605 B.n314 B.n313 585
R1606 B.n315 B.n130 585
R1607 B.n317 B.n316 585
R1608 B.n318 B.n129 585
R1609 B.n320 B.n319 585
R1610 B.n321 B.n128 585
R1611 B.n323 B.n322 585
R1612 B.n324 B.n127 585
R1613 B.n326 B.n325 585
R1614 B.n327 B.n126 585
R1615 B.n329 B.n328 585
R1616 B.n330 B.n125 585
R1617 B.n332 B.n331 585
R1618 B.n333 B.n124 585
R1619 B.n335 B.n334 585
R1620 B.n336 B.n123 585
R1621 B.n338 B.n337 585
R1622 B.n339 B.n122 585
R1623 B.n341 B.n340 585
R1624 B.n342 B.n121 585
R1625 B.n344 B.n343 585
R1626 B.n345 B.n120 585
R1627 B.n347 B.n346 585
R1628 B.n348 B.n119 585
R1629 B.n350 B.n349 585
R1630 B.n351 B.n118 585
R1631 B.n353 B.n352 585
R1632 B.n354 B.n117 585
R1633 B.n356 B.n355 585
R1634 B.n357 B.n116 585
R1635 B.n359 B.n358 585
R1636 B.n360 B.n115 585
R1637 B.n362 B.n361 585
R1638 B.n363 B.n114 585
R1639 B.n365 B.n364 585
R1640 B.n366 B.n113 585
R1641 B.n368 B.n367 585
R1642 B.n369 B.n112 585
R1643 B.n371 B.n370 585
R1644 B.n372 B.n111 585
R1645 B.n374 B.n373 585
R1646 B.n375 B.n110 585
R1647 B.n377 B.n376 585
R1648 B.n378 B.n109 585
R1649 B.n380 B.n379 585
R1650 B.n381 B.n108 585
R1651 B.n383 B.n382 585
R1652 B.n384 B.n107 585
R1653 B.n386 B.n385 585
R1654 B.n387 B.n106 585
R1655 B.n389 B.n388 585
R1656 B.n390 B.n105 585
R1657 B.n392 B.n391 585
R1658 B.n393 B.n104 585
R1659 B.n395 B.n394 585
R1660 B.n396 B.n103 585
R1661 B.n398 B.n397 585
R1662 B.n399 B.n102 585
R1663 B.n401 B.n400 585
R1664 B.n402 B.n101 585
R1665 B.n404 B.n403 585
R1666 B.n405 B.n100 585
R1667 B.n407 B.n406 585
R1668 B.n408 B.n99 585
R1669 B.n200 B.n199 585
R1670 B.n198 B.n173 585
R1671 B.n197 B.n196 585
R1672 B.n195 B.n174 585
R1673 B.n194 B.n193 585
R1674 B.n192 B.n175 585
R1675 B.n191 B.n190 585
R1676 B.n189 B.n176 585
R1677 B.n188 B.n187 585
R1678 B.n186 B.n177 585
R1679 B.n185 B.n184 585
R1680 B.n183 B.n178 585
R1681 B.n182 B.n181 585
R1682 B.n180 B.n179 585
R1683 B.n2 B.n0 585
R1684 B.n685 B.n1 585
R1685 B.n684 B.n683 585
R1686 B.n682 B.n3 585
R1687 B.n681 B.n680 585
R1688 B.n679 B.n4 585
R1689 B.n678 B.n677 585
R1690 B.n676 B.n5 585
R1691 B.n675 B.n674 585
R1692 B.n673 B.n6 585
R1693 B.n672 B.n671 585
R1694 B.n670 B.n7 585
R1695 B.n669 B.n668 585
R1696 B.n667 B.n8 585
R1697 B.n666 B.n665 585
R1698 B.n664 B.n9 585
R1699 B.n687 B.n686 585
R1700 B.n131 B.t8 528.101
R1701 B.n50 B.t4 528.101
R1702 B.n139 B.t11 528.101
R1703 B.n42 B.t1 528.101
R1704 B.n132 B.t7 513.168
R1705 B.n51 B.t5 513.168
R1706 B.n140 B.t10 513.168
R1707 B.n43 B.t2 513.168
R1708 B.n199 B.n172 458.866
R1709 B.n662 B.n9 458.866
R1710 B.n409 B.n408 458.866
R1711 B.n456 B.n455 458.866
R1712 B.n199 B.n198 163.367
R1713 B.n198 B.n197 163.367
R1714 B.n197 B.n174 163.367
R1715 B.n193 B.n174 163.367
R1716 B.n193 B.n192 163.367
R1717 B.n192 B.n191 163.367
R1718 B.n191 B.n176 163.367
R1719 B.n187 B.n176 163.367
R1720 B.n187 B.n186 163.367
R1721 B.n186 B.n185 163.367
R1722 B.n185 B.n178 163.367
R1723 B.n181 B.n178 163.367
R1724 B.n181 B.n180 163.367
R1725 B.n180 B.n2 163.367
R1726 B.n686 B.n2 163.367
R1727 B.n686 B.n685 163.367
R1728 B.n685 B.n684 163.367
R1729 B.n684 B.n3 163.367
R1730 B.n680 B.n3 163.367
R1731 B.n680 B.n679 163.367
R1732 B.n679 B.n678 163.367
R1733 B.n678 B.n5 163.367
R1734 B.n674 B.n5 163.367
R1735 B.n674 B.n673 163.367
R1736 B.n673 B.n672 163.367
R1737 B.n672 B.n7 163.367
R1738 B.n668 B.n7 163.367
R1739 B.n668 B.n667 163.367
R1740 B.n667 B.n666 163.367
R1741 B.n666 B.n9 163.367
R1742 B.n203 B.n172 163.367
R1743 B.n204 B.n203 163.367
R1744 B.n205 B.n204 163.367
R1745 B.n205 B.n170 163.367
R1746 B.n209 B.n170 163.367
R1747 B.n210 B.n209 163.367
R1748 B.n211 B.n210 163.367
R1749 B.n211 B.n168 163.367
R1750 B.n215 B.n168 163.367
R1751 B.n216 B.n215 163.367
R1752 B.n217 B.n216 163.367
R1753 B.n217 B.n166 163.367
R1754 B.n221 B.n166 163.367
R1755 B.n222 B.n221 163.367
R1756 B.n223 B.n222 163.367
R1757 B.n223 B.n164 163.367
R1758 B.n227 B.n164 163.367
R1759 B.n228 B.n227 163.367
R1760 B.n229 B.n228 163.367
R1761 B.n229 B.n162 163.367
R1762 B.n233 B.n162 163.367
R1763 B.n234 B.n233 163.367
R1764 B.n235 B.n234 163.367
R1765 B.n235 B.n160 163.367
R1766 B.n239 B.n160 163.367
R1767 B.n240 B.n239 163.367
R1768 B.n241 B.n240 163.367
R1769 B.n241 B.n158 163.367
R1770 B.n245 B.n158 163.367
R1771 B.n246 B.n245 163.367
R1772 B.n247 B.n246 163.367
R1773 B.n247 B.n156 163.367
R1774 B.n251 B.n156 163.367
R1775 B.n252 B.n251 163.367
R1776 B.n253 B.n252 163.367
R1777 B.n253 B.n154 163.367
R1778 B.n257 B.n154 163.367
R1779 B.n258 B.n257 163.367
R1780 B.n259 B.n258 163.367
R1781 B.n259 B.n152 163.367
R1782 B.n263 B.n152 163.367
R1783 B.n264 B.n263 163.367
R1784 B.n265 B.n264 163.367
R1785 B.n265 B.n150 163.367
R1786 B.n269 B.n150 163.367
R1787 B.n270 B.n269 163.367
R1788 B.n271 B.n270 163.367
R1789 B.n271 B.n148 163.367
R1790 B.n275 B.n148 163.367
R1791 B.n276 B.n275 163.367
R1792 B.n277 B.n276 163.367
R1793 B.n277 B.n146 163.367
R1794 B.n281 B.n146 163.367
R1795 B.n282 B.n281 163.367
R1796 B.n283 B.n282 163.367
R1797 B.n283 B.n144 163.367
R1798 B.n287 B.n144 163.367
R1799 B.n288 B.n287 163.367
R1800 B.n289 B.n288 163.367
R1801 B.n289 B.n142 163.367
R1802 B.n293 B.n142 163.367
R1803 B.n294 B.n293 163.367
R1804 B.n295 B.n294 163.367
R1805 B.n295 B.n138 163.367
R1806 B.n300 B.n138 163.367
R1807 B.n301 B.n300 163.367
R1808 B.n302 B.n301 163.367
R1809 B.n302 B.n136 163.367
R1810 B.n306 B.n136 163.367
R1811 B.n307 B.n306 163.367
R1812 B.n308 B.n307 163.367
R1813 B.n308 B.n134 163.367
R1814 B.n312 B.n134 163.367
R1815 B.n313 B.n312 163.367
R1816 B.n313 B.n130 163.367
R1817 B.n317 B.n130 163.367
R1818 B.n318 B.n317 163.367
R1819 B.n319 B.n318 163.367
R1820 B.n319 B.n128 163.367
R1821 B.n323 B.n128 163.367
R1822 B.n324 B.n323 163.367
R1823 B.n325 B.n324 163.367
R1824 B.n325 B.n126 163.367
R1825 B.n329 B.n126 163.367
R1826 B.n330 B.n329 163.367
R1827 B.n331 B.n330 163.367
R1828 B.n331 B.n124 163.367
R1829 B.n335 B.n124 163.367
R1830 B.n336 B.n335 163.367
R1831 B.n337 B.n336 163.367
R1832 B.n337 B.n122 163.367
R1833 B.n341 B.n122 163.367
R1834 B.n342 B.n341 163.367
R1835 B.n343 B.n342 163.367
R1836 B.n343 B.n120 163.367
R1837 B.n347 B.n120 163.367
R1838 B.n348 B.n347 163.367
R1839 B.n349 B.n348 163.367
R1840 B.n349 B.n118 163.367
R1841 B.n353 B.n118 163.367
R1842 B.n354 B.n353 163.367
R1843 B.n355 B.n354 163.367
R1844 B.n355 B.n116 163.367
R1845 B.n359 B.n116 163.367
R1846 B.n360 B.n359 163.367
R1847 B.n361 B.n360 163.367
R1848 B.n361 B.n114 163.367
R1849 B.n365 B.n114 163.367
R1850 B.n366 B.n365 163.367
R1851 B.n367 B.n366 163.367
R1852 B.n367 B.n112 163.367
R1853 B.n371 B.n112 163.367
R1854 B.n372 B.n371 163.367
R1855 B.n373 B.n372 163.367
R1856 B.n373 B.n110 163.367
R1857 B.n377 B.n110 163.367
R1858 B.n378 B.n377 163.367
R1859 B.n379 B.n378 163.367
R1860 B.n379 B.n108 163.367
R1861 B.n383 B.n108 163.367
R1862 B.n384 B.n383 163.367
R1863 B.n385 B.n384 163.367
R1864 B.n385 B.n106 163.367
R1865 B.n389 B.n106 163.367
R1866 B.n390 B.n389 163.367
R1867 B.n391 B.n390 163.367
R1868 B.n391 B.n104 163.367
R1869 B.n395 B.n104 163.367
R1870 B.n396 B.n395 163.367
R1871 B.n397 B.n396 163.367
R1872 B.n397 B.n102 163.367
R1873 B.n401 B.n102 163.367
R1874 B.n402 B.n401 163.367
R1875 B.n403 B.n402 163.367
R1876 B.n403 B.n100 163.367
R1877 B.n407 B.n100 163.367
R1878 B.n408 B.n407 163.367
R1879 B.n409 B.n98 163.367
R1880 B.n413 B.n98 163.367
R1881 B.n414 B.n413 163.367
R1882 B.n415 B.n414 163.367
R1883 B.n415 B.n96 163.367
R1884 B.n419 B.n96 163.367
R1885 B.n420 B.n419 163.367
R1886 B.n421 B.n420 163.367
R1887 B.n421 B.n94 163.367
R1888 B.n425 B.n94 163.367
R1889 B.n426 B.n425 163.367
R1890 B.n427 B.n426 163.367
R1891 B.n427 B.n92 163.367
R1892 B.n431 B.n92 163.367
R1893 B.n432 B.n431 163.367
R1894 B.n433 B.n432 163.367
R1895 B.n433 B.n90 163.367
R1896 B.n437 B.n90 163.367
R1897 B.n438 B.n437 163.367
R1898 B.n439 B.n438 163.367
R1899 B.n439 B.n88 163.367
R1900 B.n443 B.n88 163.367
R1901 B.n444 B.n443 163.367
R1902 B.n445 B.n444 163.367
R1903 B.n445 B.n86 163.367
R1904 B.n449 B.n86 163.367
R1905 B.n450 B.n449 163.367
R1906 B.n451 B.n450 163.367
R1907 B.n451 B.n84 163.367
R1908 B.n455 B.n84 163.367
R1909 B.n662 B.n661 163.367
R1910 B.n661 B.n660 163.367
R1911 B.n660 B.n11 163.367
R1912 B.n656 B.n11 163.367
R1913 B.n656 B.n655 163.367
R1914 B.n655 B.n654 163.367
R1915 B.n654 B.n13 163.367
R1916 B.n650 B.n13 163.367
R1917 B.n650 B.n649 163.367
R1918 B.n649 B.n648 163.367
R1919 B.n648 B.n15 163.367
R1920 B.n644 B.n15 163.367
R1921 B.n644 B.n643 163.367
R1922 B.n643 B.n642 163.367
R1923 B.n642 B.n17 163.367
R1924 B.n638 B.n17 163.367
R1925 B.n638 B.n637 163.367
R1926 B.n637 B.n636 163.367
R1927 B.n636 B.n19 163.367
R1928 B.n632 B.n19 163.367
R1929 B.n632 B.n631 163.367
R1930 B.n631 B.n630 163.367
R1931 B.n630 B.n21 163.367
R1932 B.n626 B.n21 163.367
R1933 B.n626 B.n625 163.367
R1934 B.n625 B.n624 163.367
R1935 B.n624 B.n23 163.367
R1936 B.n620 B.n23 163.367
R1937 B.n620 B.n619 163.367
R1938 B.n619 B.n618 163.367
R1939 B.n618 B.n25 163.367
R1940 B.n614 B.n25 163.367
R1941 B.n614 B.n613 163.367
R1942 B.n613 B.n612 163.367
R1943 B.n612 B.n27 163.367
R1944 B.n608 B.n27 163.367
R1945 B.n608 B.n607 163.367
R1946 B.n607 B.n606 163.367
R1947 B.n606 B.n29 163.367
R1948 B.n602 B.n29 163.367
R1949 B.n602 B.n601 163.367
R1950 B.n601 B.n600 163.367
R1951 B.n600 B.n31 163.367
R1952 B.n596 B.n31 163.367
R1953 B.n596 B.n595 163.367
R1954 B.n595 B.n594 163.367
R1955 B.n594 B.n33 163.367
R1956 B.n590 B.n33 163.367
R1957 B.n590 B.n589 163.367
R1958 B.n589 B.n588 163.367
R1959 B.n588 B.n35 163.367
R1960 B.n584 B.n35 163.367
R1961 B.n584 B.n583 163.367
R1962 B.n583 B.n582 163.367
R1963 B.n582 B.n37 163.367
R1964 B.n578 B.n37 163.367
R1965 B.n578 B.n577 163.367
R1966 B.n577 B.n576 163.367
R1967 B.n576 B.n39 163.367
R1968 B.n572 B.n39 163.367
R1969 B.n572 B.n571 163.367
R1970 B.n571 B.n570 163.367
R1971 B.n570 B.n41 163.367
R1972 B.n565 B.n41 163.367
R1973 B.n565 B.n564 163.367
R1974 B.n564 B.n563 163.367
R1975 B.n563 B.n45 163.367
R1976 B.n559 B.n45 163.367
R1977 B.n559 B.n558 163.367
R1978 B.n558 B.n557 163.367
R1979 B.n557 B.n47 163.367
R1980 B.n553 B.n47 163.367
R1981 B.n553 B.n552 163.367
R1982 B.n552 B.n551 163.367
R1983 B.n551 B.n49 163.367
R1984 B.n547 B.n49 163.367
R1985 B.n547 B.n546 163.367
R1986 B.n546 B.n545 163.367
R1987 B.n545 B.n54 163.367
R1988 B.n541 B.n54 163.367
R1989 B.n541 B.n540 163.367
R1990 B.n540 B.n539 163.367
R1991 B.n539 B.n56 163.367
R1992 B.n535 B.n56 163.367
R1993 B.n535 B.n534 163.367
R1994 B.n534 B.n533 163.367
R1995 B.n533 B.n58 163.367
R1996 B.n529 B.n58 163.367
R1997 B.n529 B.n528 163.367
R1998 B.n528 B.n527 163.367
R1999 B.n527 B.n60 163.367
R2000 B.n523 B.n60 163.367
R2001 B.n523 B.n522 163.367
R2002 B.n522 B.n521 163.367
R2003 B.n521 B.n62 163.367
R2004 B.n517 B.n62 163.367
R2005 B.n517 B.n516 163.367
R2006 B.n516 B.n515 163.367
R2007 B.n515 B.n64 163.367
R2008 B.n511 B.n64 163.367
R2009 B.n511 B.n510 163.367
R2010 B.n510 B.n509 163.367
R2011 B.n509 B.n66 163.367
R2012 B.n505 B.n66 163.367
R2013 B.n505 B.n504 163.367
R2014 B.n504 B.n503 163.367
R2015 B.n503 B.n68 163.367
R2016 B.n499 B.n68 163.367
R2017 B.n499 B.n498 163.367
R2018 B.n498 B.n497 163.367
R2019 B.n497 B.n70 163.367
R2020 B.n493 B.n70 163.367
R2021 B.n493 B.n492 163.367
R2022 B.n492 B.n491 163.367
R2023 B.n491 B.n72 163.367
R2024 B.n487 B.n72 163.367
R2025 B.n487 B.n486 163.367
R2026 B.n486 B.n485 163.367
R2027 B.n485 B.n74 163.367
R2028 B.n481 B.n74 163.367
R2029 B.n481 B.n480 163.367
R2030 B.n480 B.n479 163.367
R2031 B.n479 B.n76 163.367
R2032 B.n475 B.n76 163.367
R2033 B.n475 B.n474 163.367
R2034 B.n474 B.n473 163.367
R2035 B.n473 B.n78 163.367
R2036 B.n469 B.n78 163.367
R2037 B.n469 B.n468 163.367
R2038 B.n468 B.n467 163.367
R2039 B.n467 B.n80 163.367
R2040 B.n463 B.n80 163.367
R2041 B.n463 B.n462 163.367
R2042 B.n462 B.n461 163.367
R2043 B.n461 B.n82 163.367
R2044 B.n457 B.n82 163.367
R2045 B.n457 B.n456 163.367
R2046 B.n133 B.n132 59.5399
R2047 B.n297 B.n140 59.5399
R2048 B.n567 B.n43 59.5399
R2049 B.n52 B.n51 59.5399
R2050 B.n664 B.n663 29.8151
R2051 B.n454 B.n83 29.8151
R2052 B.n410 B.n99 29.8151
R2053 B.n201 B.n200 29.8151
R2054 B B.n687 18.0485
R2055 B.n132 B.n131 14.9338
R2056 B.n140 B.n139 14.9338
R2057 B.n43 B.n42 14.9338
R2058 B.n51 B.n50 14.9338
R2059 B.n663 B.n10 10.6151
R2060 B.n659 B.n10 10.6151
R2061 B.n659 B.n658 10.6151
R2062 B.n658 B.n657 10.6151
R2063 B.n657 B.n12 10.6151
R2064 B.n653 B.n12 10.6151
R2065 B.n653 B.n652 10.6151
R2066 B.n652 B.n651 10.6151
R2067 B.n651 B.n14 10.6151
R2068 B.n647 B.n14 10.6151
R2069 B.n647 B.n646 10.6151
R2070 B.n646 B.n645 10.6151
R2071 B.n645 B.n16 10.6151
R2072 B.n641 B.n16 10.6151
R2073 B.n641 B.n640 10.6151
R2074 B.n640 B.n639 10.6151
R2075 B.n639 B.n18 10.6151
R2076 B.n635 B.n18 10.6151
R2077 B.n635 B.n634 10.6151
R2078 B.n634 B.n633 10.6151
R2079 B.n633 B.n20 10.6151
R2080 B.n629 B.n20 10.6151
R2081 B.n629 B.n628 10.6151
R2082 B.n628 B.n627 10.6151
R2083 B.n627 B.n22 10.6151
R2084 B.n623 B.n22 10.6151
R2085 B.n623 B.n622 10.6151
R2086 B.n622 B.n621 10.6151
R2087 B.n621 B.n24 10.6151
R2088 B.n617 B.n24 10.6151
R2089 B.n617 B.n616 10.6151
R2090 B.n616 B.n615 10.6151
R2091 B.n615 B.n26 10.6151
R2092 B.n611 B.n26 10.6151
R2093 B.n611 B.n610 10.6151
R2094 B.n610 B.n609 10.6151
R2095 B.n609 B.n28 10.6151
R2096 B.n605 B.n28 10.6151
R2097 B.n605 B.n604 10.6151
R2098 B.n604 B.n603 10.6151
R2099 B.n603 B.n30 10.6151
R2100 B.n599 B.n30 10.6151
R2101 B.n599 B.n598 10.6151
R2102 B.n598 B.n597 10.6151
R2103 B.n597 B.n32 10.6151
R2104 B.n593 B.n32 10.6151
R2105 B.n593 B.n592 10.6151
R2106 B.n592 B.n591 10.6151
R2107 B.n591 B.n34 10.6151
R2108 B.n587 B.n34 10.6151
R2109 B.n587 B.n586 10.6151
R2110 B.n586 B.n585 10.6151
R2111 B.n585 B.n36 10.6151
R2112 B.n581 B.n36 10.6151
R2113 B.n581 B.n580 10.6151
R2114 B.n580 B.n579 10.6151
R2115 B.n579 B.n38 10.6151
R2116 B.n575 B.n38 10.6151
R2117 B.n575 B.n574 10.6151
R2118 B.n574 B.n573 10.6151
R2119 B.n573 B.n40 10.6151
R2120 B.n569 B.n40 10.6151
R2121 B.n569 B.n568 10.6151
R2122 B.n566 B.n44 10.6151
R2123 B.n562 B.n44 10.6151
R2124 B.n562 B.n561 10.6151
R2125 B.n561 B.n560 10.6151
R2126 B.n560 B.n46 10.6151
R2127 B.n556 B.n46 10.6151
R2128 B.n556 B.n555 10.6151
R2129 B.n555 B.n554 10.6151
R2130 B.n554 B.n48 10.6151
R2131 B.n550 B.n549 10.6151
R2132 B.n549 B.n548 10.6151
R2133 B.n548 B.n53 10.6151
R2134 B.n544 B.n53 10.6151
R2135 B.n544 B.n543 10.6151
R2136 B.n543 B.n542 10.6151
R2137 B.n542 B.n55 10.6151
R2138 B.n538 B.n55 10.6151
R2139 B.n538 B.n537 10.6151
R2140 B.n537 B.n536 10.6151
R2141 B.n536 B.n57 10.6151
R2142 B.n532 B.n57 10.6151
R2143 B.n532 B.n531 10.6151
R2144 B.n531 B.n530 10.6151
R2145 B.n530 B.n59 10.6151
R2146 B.n526 B.n59 10.6151
R2147 B.n526 B.n525 10.6151
R2148 B.n525 B.n524 10.6151
R2149 B.n524 B.n61 10.6151
R2150 B.n520 B.n61 10.6151
R2151 B.n520 B.n519 10.6151
R2152 B.n519 B.n518 10.6151
R2153 B.n518 B.n63 10.6151
R2154 B.n514 B.n63 10.6151
R2155 B.n514 B.n513 10.6151
R2156 B.n513 B.n512 10.6151
R2157 B.n512 B.n65 10.6151
R2158 B.n508 B.n65 10.6151
R2159 B.n508 B.n507 10.6151
R2160 B.n507 B.n506 10.6151
R2161 B.n506 B.n67 10.6151
R2162 B.n502 B.n67 10.6151
R2163 B.n502 B.n501 10.6151
R2164 B.n501 B.n500 10.6151
R2165 B.n500 B.n69 10.6151
R2166 B.n496 B.n69 10.6151
R2167 B.n496 B.n495 10.6151
R2168 B.n495 B.n494 10.6151
R2169 B.n494 B.n71 10.6151
R2170 B.n490 B.n71 10.6151
R2171 B.n490 B.n489 10.6151
R2172 B.n489 B.n488 10.6151
R2173 B.n488 B.n73 10.6151
R2174 B.n484 B.n73 10.6151
R2175 B.n484 B.n483 10.6151
R2176 B.n483 B.n482 10.6151
R2177 B.n482 B.n75 10.6151
R2178 B.n478 B.n75 10.6151
R2179 B.n478 B.n477 10.6151
R2180 B.n477 B.n476 10.6151
R2181 B.n476 B.n77 10.6151
R2182 B.n472 B.n77 10.6151
R2183 B.n472 B.n471 10.6151
R2184 B.n471 B.n470 10.6151
R2185 B.n470 B.n79 10.6151
R2186 B.n466 B.n79 10.6151
R2187 B.n466 B.n465 10.6151
R2188 B.n465 B.n464 10.6151
R2189 B.n464 B.n81 10.6151
R2190 B.n460 B.n81 10.6151
R2191 B.n460 B.n459 10.6151
R2192 B.n459 B.n458 10.6151
R2193 B.n458 B.n83 10.6151
R2194 B.n411 B.n410 10.6151
R2195 B.n412 B.n411 10.6151
R2196 B.n412 B.n97 10.6151
R2197 B.n416 B.n97 10.6151
R2198 B.n417 B.n416 10.6151
R2199 B.n418 B.n417 10.6151
R2200 B.n418 B.n95 10.6151
R2201 B.n422 B.n95 10.6151
R2202 B.n423 B.n422 10.6151
R2203 B.n424 B.n423 10.6151
R2204 B.n424 B.n93 10.6151
R2205 B.n428 B.n93 10.6151
R2206 B.n429 B.n428 10.6151
R2207 B.n430 B.n429 10.6151
R2208 B.n430 B.n91 10.6151
R2209 B.n434 B.n91 10.6151
R2210 B.n435 B.n434 10.6151
R2211 B.n436 B.n435 10.6151
R2212 B.n436 B.n89 10.6151
R2213 B.n440 B.n89 10.6151
R2214 B.n441 B.n440 10.6151
R2215 B.n442 B.n441 10.6151
R2216 B.n442 B.n87 10.6151
R2217 B.n446 B.n87 10.6151
R2218 B.n447 B.n446 10.6151
R2219 B.n448 B.n447 10.6151
R2220 B.n448 B.n85 10.6151
R2221 B.n452 B.n85 10.6151
R2222 B.n453 B.n452 10.6151
R2223 B.n454 B.n453 10.6151
R2224 B.n202 B.n201 10.6151
R2225 B.n202 B.n171 10.6151
R2226 B.n206 B.n171 10.6151
R2227 B.n207 B.n206 10.6151
R2228 B.n208 B.n207 10.6151
R2229 B.n208 B.n169 10.6151
R2230 B.n212 B.n169 10.6151
R2231 B.n213 B.n212 10.6151
R2232 B.n214 B.n213 10.6151
R2233 B.n214 B.n167 10.6151
R2234 B.n218 B.n167 10.6151
R2235 B.n219 B.n218 10.6151
R2236 B.n220 B.n219 10.6151
R2237 B.n220 B.n165 10.6151
R2238 B.n224 B.n165 10.6151
R2239 B.n225 B.n224 10.6151
R2240 B.n226 B.n225 10.6151
R2241 B.n226 B.n163 10.6151
R2242 B.n230 B.n163 10.6151
R2243 B.n231 B.n230 10.6151
R2244 B.n232 B.n231 10.6151
R2245 B.n232 B.n161 10.6151
R2246 B.n236 B.n161 10.6151
R2247 B.n237 B.n236 10.6151
R2248 B.n238 B.n237 10.6151
R2249 B.n238 B.n159 10.6151
R2250 B.n242 B.n159 10.6151
R2251 B.n243 B.n242 10.6151
R2252 B.n244 B.n243 10.6151
R2253 B.n244 B.n157 10.6151
R2254 B.n248 B.n157 10.6151
R2255 B.n249 B.n248 10.6151
R2256 B.n250 B.n249 10.6151
R2257 B.n250 B.n155 10.6151
R2258 B.n254 B.n155 10.6151
R2259 B.n255 B.n254 10.6151
R2260 B.n256 B.n255 10.6151
R2261 B.n256 B.n153 10.6151
R2262 B.n260 B.n153 10.6151
R2263 B.n261 B.n260 10.6151
R2264 B.n262 B.n261 10.6151
R2265 B.n262 B.n151 10.6151
R2266 B.n266 B.n151 10.6151
R2267 B.n267 B.n266 10.6151
R2268 B.n268 B.n267 10.6151
R2269 B.n268 B.n149 10.6151
R2270 B.n272 B.n149 10.6151
R2271 B.n273 B.n272 10.6151
R2272 B.n274 B.n273 10.6151
R2273 B.n274 B.n147 10.6151
R2274 B.n278 B.n147 10.6151
R2275 B.n279 B.n278 10.6151
R2276 B.n280 B.n279 10.6151
R2277 B.n280 B.n145 10.6151
R2278 B.n284 B.n145 10.6151
R2279 B.n285 B.n284 10.6151
R2280 B.n286 B.n285 10.6151
R2281 B.n286 B.n143 10.6151
R2282 B.n290 B.n143 10.6151
R2283 B.n291 B.n290 10.6151
R2284 B.n292 B.n291 10.6151
R2285 B.n292 B.n141 10.6151
R2286 B.n296 B.n141 10.6151
R2287 B.n299 B.n298 10.6151
R2288 B.n299 B.n137 10.6151
R2289 B.n303 B.n137 10.6151
R2290 B.n304 B.n303 10.6151
R2291 B.n305 B.n304 10.6151
R2292 B.n305 B.n135 10.6151
R2293 B.n309 B.n135 10.6151
R2294 B.n310 B.n309 10.6151
R2295 B.n311 B.n310 10.6151
R2296 B.n315 B.n314 10.6151
R2297 B.n316 B.n315 10.6151
R2298 B.n316 B.n129 10.6151
R2299 B.n320 B.n129 10.6151
R2300 B.n321 B.n320 10.6151
R2301 B.n322 B.n321 10.6151
R2302 B.n322 B.n127 10.6151
R2303 B.n326 B.n127 10.6151
R2304 B.n327 B.n326 10.6151
R2305 B.n328 B.n327 10.6151
R2306 B.n328 B.n125 10.6151
R2307 B.n332 B.n125 10.6151
R2308 B.n333 B.n332 10.6151
R2309 B.n334 B.n333 10.6151
R2310 B.n334 B.n123 10.6151
R2311 B.n338 B.n123 10.6151
R2312 B.n339 B.n338 10.6151
R2313 B.n340 B.n339 10.6151
R2314 B.n340 B.n121 10.6151
R2315 B.n344 B.n121 10.6151
R2316 B.n345 B.n344 10.6151
R2317 B.n346 B.n345 10.6151
R2318 B.n346 B.n119 10.6151
R2319 B.n350 B.n119 10.6151
R2320 B.n351 B.n350 10.6151
R2321 B.n352 B.n351 10.6151
R2322 B.n352 B.n117 10.6151
R2323 B.n356 B.n117 10.6151
R2324 B.n357 B.n356 10.6151
R2325 B.n358 B.n357 10.6151
R2326 B.n358 B.n115 10.6151
R2327 B.n362 B.n115 10.6151
R2328 B.n363 B.n362 10.6151
R2329 B.n364 B.n363 10.6151
R2330 B.n364 B.n113 10.6151
R2331 B.n368 B.n113 10.6151
R2332 B.n369 B.n368 10.6151
R2333 B.n370 B.n369 10.6151
R2334 B.n370 B.n111 10.6151
R2335 B.n374 B.n111 10.6151
R2336 B.n375 B.n374 10.6151
R2337 B.n376 B.n375 10.6151
R2338 B.n376 B.n109 10.6151
R2339 B.n380 B.n109 10.6151
R2340 B.n381 B.n380 10.6151
R2341 B.n382 B.n381 10.6151
R2342 B.n382 B.n107 10.6151
R2343 B.n386 B.n107 10.6151
R2344 B.n387 B.n386 10.6151
R2345 B.n388 B.n387 10.6151
R2346 B.n388 B.n105 10.6151
R2347 B.n392 B.n105 10.6151
R2348 B.n393 B.n392 10.6151
R2349 B.n394 B.n393 10.6151
R2350 B.n394 B.n103 10.6151
R2351 B.n398 B.n103 10.6151
R2352 B.n399 B.n398 10.6151
R2353 B.n400 B.n399 10.6151
R2354 B.n400 B.n101 10.6151
R2355 B.n404 B.n101 10.6151
R2356 B.n405 B.n404 10.6151
R2357 B.n406 B.n405 10.6151
R2358 B.n406 B.n99 10.6151
R2359 B.n200 B.n173 10.6151
R2360 B.n196 B.n173 10.6151
R2361 B.n196 B.n195 10.6151
R2362 B.n195 B.n194 10.6151
R2363 B.n194 B.n175 10.6151
R2364 B.n190 B.n175 10.6151
R2365 B.n190 B.n189 10.6151
R2366 B.n189 B.n188 10.6151
R2367 B.n188 B.n177 10.6151
R2368 B.n184 B.n177 10.6151
R2369 B.n184 B.n183 10.6151
R2370 B.n183 B.n182 10.6151
R2371 B.n182 B.n179 10.6151
R2372 B.n179 B.n0 10.6151
R2373 B.n683 B.n1 10.6151
R2374 B.n683 B.n682 10.6151
R2375 B.n682 B.n681 10.6151
R2376 B.n681 B.n4 10.6151
R2377 B.n677 B.n4 10.6151
R2378 B.n677 B.n676 10.6151
R2379 B.n676 B.n675 10.6151
R2380 B.n675 B.n6 10.6151
R2381 B.n671 B.n6 10.6151
R2382 B.n671 B.n670 10.6151
R2383 B.n670 B.n669 10.6151
R2384 B.n669 B.n8 10.6151
R2385 B.n665 B.n8 10.6151
R2386 B.n665 B.n664 10.6151
R2387 B.n568 B.n567 9.36635
R2388 B.n550 B.n52 9.36635
R2389 B.n297 B.n296 9.36635
R2390 B.n314 B.n133 9.36635
R2391 B.n687 B.n0 2.81026
R2392 B.n687 B.n1 2.81026
R2393 B.n567 B.n566 1.24928
R2394 B.n52 B.n48 1.24928
R2395 B.n298 B.n297 1.24928
R2396 B.n311 B.n133 1.24928
C0 VTAIL VN 3.16044f
C1 w_n1432_n4894# VN 2.17238f
C2 VTAIL w_n1432_n4894# 6.22008f
C3 VP VN 6.04983f
C4 VDD1 VN 0.147151f
C5 VTAIL VP 3.17454f
C6 VTAIL VDD1 12.411599f
C7 VDD2 VN 3.95356f
C8 VTAIL VDD2 12.4513f
C9 w_n1432_n4894# VP 2.351f
C10 VDD1 w_n1432_n4894# 1.21056f
C11 VDD1 VP 4.06318f
C12 B VN 0.784931f
C13 VDD2 w_n1432_n4894# 1.22006f
C14 VTAIL B 5.58655f
C15 VDD2 VP 0.256964f
C16 VDD1 VDD2 0.510386f
C17 w_n1432_n4894# B 8.72723f
C18 B VP 1.0713f
C19 VDD1 B 1.08519f
C20 VDD2 B 1.10308f
C21 VDD2 VSUBS 0.832678f
C22 VDD1 VSUBS 6.422301f
C23 VTAIL VSUBS 1.084035f
C24 VN VSUBS 7.20141f
C25 VP VSUBS 1.443937f
C26 B VSUBS 3.042126f
C27 w_n1432_n4894# VSUBS 85.5935f
C28 B.n0 VSUBS 0.005059f
C29 B.n1 VSUBS 0.005059f
C30 B.n2 VSUBS 0.008001f
C31 B.n3 VSUBS 0.008001f
C32 B.n4 VSUBS 0.008001f
C33 B.n5 VSUBS 0.008001f
C34 B.n6 VSUBS 0.008001f
C35 B.n7 VSUBS 0.008001f
C36 B.n8 VSUBS 0.008001f
C37 B.n9 VSUBS 0.017106f
C38 B.n10 VSUBS 0.008001f
C39 B.n11 VSUBS 0.008001f
C40 B.n12 VSUBS 0.008001f
C41 B.n13 VSUBS 0.008001f
C42 B.n14 VSUBS 0.008001f
C43 B.n15 VSUBS 0.008001f
C44 B.n16 VSUBS 0.008001f
C45 B.n17 VSUBS 0.008001f
C46 B.n18 VSUBS 0.008001f
C47 B.n19 VSUBS 0.008001f
C48 B.n20 VSUBS 0.008001f
C49 B.n21 VSUBS 0.008001f
C50 B.n22 VSUBS 0.008001f
C51 B.n23 VSUBS 0.008001f
C52 B.n24 VSUBS 0.008001f
C53 B.n25 VSUBS 0.008001f
C54 B.n26 VSUBS 0.008001f
C55 B.n27 VSUBS 0.008001f
C56 B.n28 VSUBS 0.008001f
C57 B.n29 VSUBS 0.008001f
C58 B.n30 VSUBS 0.008001f
C59 B.n31 VSUBS 0.008001f
C60 B.n32 VSUBS 0.008001f
C61 B.n33 VSUBS 0.008001f
C62 B.n34 VSUBS 0.008001f
C63 B.n35 VSUBS 0.008001f
C64 B.n36 VSUBS 0.008001f
C65 B.n37 VSUBS 0.008001f
C66 B.n38 VSUBS 0.008001f
C67 B.n39 VSUBS 0.008001f
C68 B.n40 VSUBS 0.008001f
C69 B.n41 VSUBS 0.008001f
C70 B.t2 VSUBS 0.446775f
C71 B.t1 VSUBS 0.457406f
C72 B.t0 VSUBS 0.387309f
C73 B.n42 VSUBS 0.487278f
C74 B.n43 VSUBS 0.387351f
C75 B.n44 VSUBS 0.008001f
C76 B.n45 VSUBS 0.008001f
C77 B.n46 VSUBS 0.008001f
C78 B.n47 VSUBS 0.008001f
C79 B.n48 VSUBS 0.004471f
C80 B.n49 VSUBS 0.008001f
C81 B.t5 VSUBS 0.446779f
C82 B.t4 VSUBS 0.45741f
C83 B.t3 VSUBS 0.387309f
C84 B.n50 VSUBS 0.487274f
C85 B.n51 VSUBS 0.387347f
C86 B.n52 VSUBS 0.018537f
C87 B.n53 VSUBS 0.008001f
C88 B.n54 VSUBS 0.008001f
C89 B.n55 VSUBS 0.008001f
C90 B.n56 VSUBS 0.008001f
C91 B.n57 VSUBS 0.008001f
C92 B.n58 VSUBS 0.008001f
C93 B.n59 VSUBS 0.008001f
C94 B.n60 VSUBS 0.008001f
C95 B.n61 VSUBS 0.008001f
C96 B.n62 VSUBS 0.008001f
C97 B.n63 VSUBS 0.008001f
C98 B.n64 VSUBS 0.008001f
C99 B.n65 VSUBS 0.008001f
C100 B.n66 VSUBS 0.008001f
C101 B.n67 VSUBS 0.008001f
C102 B.n68 VSUBS 0.008001f
C103 B.n69 VSUBS 0.008001f
C104 B.n70 VSUBS 0.008001f
C105 B.n71 VSUBS 0.008001f
C106 B.n72 VSUBS 0.008001f
C107 B.n73 VSUBS 0.008001f
C108 B.n74 VSUBS 0.008001f
C109 B.n75 VSUBS 0.008001f
C110 B.n76 VSUBS 0.008001f
C111 B.n77 VSUBS 0.008001f
C112 B.n78 VSUBS 0.008001f
C113 B.n79 VSUBS 0.008001f
C114 B.n80 VSUBS 0.008001f
C115 B.n81 VSUBS 0.008001f
C116 B.n82 VSUBS 0.008001f
C117 B.n83 VSUBS 0.017157f
C118 B.n84 VSUBS 0.008001f
C119 B.n85 VSUBS 0.008001f
C120 B.n86 VSUBS 0.008001f
C121 B.n87 VSUBS 0.008001f
C122 B.n88 VSUBS 0.008001f
C123 B.n89 VSUBS 0.008001f
C124 B.n90 VSUBS 0.008001f
C125 B.n91 VSUBS 0.008001f
C126 B.n92 VSUBS 0.008001f
C127 B.n93 VSUBS 0.008001f
C128 B.n94 VSUBS 0.008001f
C129 B.n95 VSUBS 0.008001f
C130 B.n96 VSUBS 0.008001f
C131 B.n97 VSUBS 0.008001f
C132 B.n98 VSUBS 0.008001f
C133 B.n99 VSUBS 0.018192f
C134 B.n100 VSUBS 0.008001f
C135 B.n101 VSUBS 0.008001f
C136 B.n102 VSUBS 0.008001f
C137 B.n103 VSUBS 0.008001f
C138 B.n104 VSUBS 0.008001f
C139 B.n105 VSUBS 0.008001f
C140 B.n106 VSUBS 0.008001f
C141 B.n107 VSUBS 0.008001f
C142 B.n108 VSUBS 0.008001f
C143 B.n109 VSUBS 0.008001f
C144 B.n110 VSUBS 0.008001f
C145 B.n111 VSUBS 0.008001f
C146 B.n112 VSUBS 0.008001f
C147 B.n113 VSUBS 0.008001f
C148 B.n114 VSUBS 0.008001f
C149 B.n115 VSUBS 0.008001f
C150 B.n116 VSUBS 0.008001f
C151 B.n117 VSUBS 0.008001f
C152 B.n118 VSUBS 0.008001f
C153 B.n119 VSUBS 0.008001f
C154 B.n120 VSUBS 0.008001f
C155 B.n121 VSUBS 0.008001f
C156 B.n122 VSUBS 0.008001f
C157 B.n123 VSUBS 0.008001f
C158 B.n124 VSUBS 0.008001f
C159 B.n125 VSUBS 0.008001f
C160 B.n126 VSUBS 0.008001f
C161 B.n127 VSUBS 0.008001f
C162 B.n128 VSUBS 0.008001f
C163 B.n129 VSUBS 0.008001f
C164 B.n130 VSUBS 0.008001f
C165 B.t7 VSUBS 0.446779f
C166 B.t8 VSUBS 0.45741f
C167 B.t6 VSUBS 0.387309f
C168 B.n131 VSUBS 0.487274f
C169 B.n132 VSUBS 0.387347f
C170 B.n133 VSUBS 0.018537f
C171 B.n134 VSUBS 0.008001f
C172 B.n135 VSUBS 0.008001f
C173 B.n136 VSUBS 0.008001f
C174 B.n137 VSUBS 0.008001f
C175 B.n138 VSUBS 0.008001f
C176 B.t10 VSUBS 0.446775f
C177 B.t11 VSUBS 0.457406f
C178 B.t9 VSUBS 0.387309f
C179 B.n139 VSUBS 0.487278f
C180 B.n140 VSUBS 0.387351f
C181 B.n141 VSUBS 0.008001f
C182 B.n142 VSUBS 0.008001f
C183 B.n143 VSUBS 0.008001f
C184 B.n144 VSUBS 0.008001f
C185 B.n145 VSUBS 0.008001f
C186 B.n146 VSUBS 0.008001f
C187 B.n147 VSUBS 0.008001f
C188 B.n148 VSUBS 0.008001f
C189 B.n149 VSUBS 0.008001f
C190 B.n150 VSUBS 0.008001f
C191 B.n151 VSUBS 0.008001f
C192 B.n152 VSUBS 0.008001f
C193 B.n153 VSUBS 0.008001f
C194 B.n154 VSUBS 0.008001f
C195 B.n155 VSUBS 0.008001f
C196 B.n156 VSUBS 0.008001f
C197 B.n157 VSUBS 0.008001f
C198 B.n158 VSUBS 0.008001f
C199 B.n159 VSUBS 0.008001f
C200 B.n160 VSUBS 0.008001f
C201 B.n161 VSUBS 0.008001f
C202 B.n162 VSUBS 0.008001f
C203 B.n163 VSUBS 0.008001f
C204 B.n164 VSUBS 0.008001f
C205 B.n165 VSUBS 0.008001f
C206 B.n166 VSUBS 0.008001f
C207 B.n167 VSUBS 0.008001f
C208 B.n168 VSUBS 0.008001f
C209 B.n169 VSUBS 0.008001f
C210 B.n170 VSUBS 0.008001f
C211 B.n171 VSUBS 0.008001f
C212 B.n172 VSUBS 0.018192f
C213 B.n173 VSUBS 0.008001f
C214 B.n174 VSUBS 0.008001f
C215 B.n175 VSUBS 0.008001f
C216 B.n176 VSUBS 0.008001f
C217 B.n177 VSUBS 0.008001f
C218 B.n178 VSUBS 0.008001f
C219 B.n179 VSUBS 0.008001f
C220 B.n180 VSUBS 0.008001f
C221 B.n181 VSUBS 0.008001f
C222 B.n182 VSUBS 0.008001f
C223 B.n183 VSUBS 0.008001f
C224 B.n184 VSUBS 0.008001f
C225 B.n185 VSUBS 0.008001f
C226 B.n186 VSUBS 0.008001f
C227 B.n187 VSUBS 0.008001f
C228 B.n188 VSUBS 0.008001f
C229 B.n189 VSUBS 0.008001f
C230 B.n190 VSUBS 0.008001f
C231 B.n191 VSUBS 0.008001f
C232 B.n192 VSUBS 0.008001f
C233 B.n193 VSUBS 0.008001f
C234 B.n194 VSUBS 0.008001f
C235 B.n195 VSUBS 0.008001f
C236 B.n196 VSUBS 0.008001f
C237 B.n197 VSUBS 0.008001f
C238 B.n198 VSUBS 0.008001f
C239 B.n199 VSUBS 0.017106f
C240 B.n200 VSUBS 0.017106f
C241 B.n201 VSUBS 0.018192f
C242 B.n202 VSUBS 0.008001f
C243 B.n203 VSUBS 0.008001f
C244 B.n204 VSUBS 0.008001f
C245 B.n205 VSUBS 0.008001f
C246 B.n206 VSUBS 0.008001f
C247 B.n207 VSUBS 0.008001f
C248 B.n208 VSUBS 0.008001f
C249 B.n209 VSUBS 0.008001f
C250 B.n210 VSUBS 0.008001f
C251 B.n211 VSUBS 0.008001f
C252 B.n212 VSUBS 0.008001f
C253 B.n213 VSUBS 0.008001f
C254 B.n214 VSUBS 0.008001f
C255 B.n215 VSUBS 0.008001f
C256 B.n216 VSUBS 0.008001f
C257 B.n217 VSUBS 0.008001f
C258 B.n218 VSUBS 0.008001f
C259 B.n219 VSUBS 0.008001f
C260 B.n220 VSUBS 0.008001f
C261 B.n221 VSUBS 0.008001f
C262 B.n222 VSUBS 0.008001f
C263 B.n223 VSUBS 0.008001f
C264 B.n224 VSUBS 0.008001f
C265 B.n225 VSUBS 0.008001f
C266 B.n226 VSUBS 0.008001f
C267 B.n227 VSUBS 0.008001f
C268 B.n228 VSUBS 0.008001f
C269 B.n229 VSUBS 0.008001f
C270 B.n230 VSUBS 0.008001f
C271 B.n231 VSUBS 0.008001f
C272 B.n232 VSUBS 0.008001f
C273 B.n233 VSUBS 0.008001f
C274 B.n234 VSUBS 0.008001f
C275 B.n235 VSUBS 0.008001f
C276 B.n236 VSUBS 0.008001f
C277 B.n237 VSUBS 0.008001f
C278 B.n238 VSUBS 0.008001f
C279 B.n239 VSUBS 0.008001f
C280 B.n240 VSUBS 0.008001f
C281 B.n241 VSUBS 0.008001f
C282 B.n242 VSUBS 0.008001f
C283 B.n243 VSUBS 0.008001f
C284 B.n244 VSUBS 0.008001f
C285 B.n245 VSUBS 0.008001f
C286 B.n246 VSUBS 0.008001f
C287 B.n247 VSUBS 0.008001f
C288 B.n248 VSUBS 0.008001f
C289 B.n249 VSUBS 0.008001f
C290 B.n250 VSUBS 0.008001f
C291 B.n251 VSUBS 0.008001f
C292 B.n252 VSUBS 0.008001f
C293 B.n253 VSUBS 0.008001f
C294 B.n254 VSUBS 0.008001f
C295 B.n255 VSUBS 0.008001f
C296 B.n256 VSUBS 0.008001f
C297 B.n257 VSUBS 0.008001f
C298 B.n258 VSUBS 0.008001f
C299 B.n259 VSUBS 0.008001f
C300 B.n260 VSUBS 0.008001f
C301 B.n261 VSUBS 0.008001f
C302 B.n262 VSUBS 0.008001f
C303 B.n263 VSUBS 0.008001f
C304 B.n264 VSUBS 0.008001f
C305 B.n265 VSUBS 0.008001f
C306 B.n266 VSUBS 0.008001f
C307 B.n267 VSUBS 0.008001f
C308 B.n268 VSUBS 0.008001f
C309 B.n269 VSUBS 0.008001f
C310 B.n270 VSUBS 0.008001f
C311 B.n271 VSUBS 0.008001f
C312 B.n272 VSUBS 0.008001f
C313 B.n273 VSUBS 0.008001f
C314 B.n274 VSUBS 0.008001f
C315 B.n275 VSUBS 0.008001f
C316 B.n276 VSUBS 0.008001f
C317 B.n277 VSUBS 0.008001f
C318 B.n278 VSUBS 0.008001f
C319 B.n279 VSUBS 0.008001f
C320 B.n280 VSUBS 0.008001f
C321 B.n281 VSUBS 0.008001f
C322 B.n282 VSUBS 0.008001f
C323 B.n283 VSUBS 0.008001f
C324 B.n284 VSUBS 0.008001f
C325 B.n285 VSUBS 0.008001f
C326 B.n286 VSUBS 0.008001f
C327 B.n287 VSUBS 0.008001f
C328 B.n288 VSUBS 0.008001f
C329 B.n289 VSUBS 0.008001f
C330 B.n290 VSUBS 0.008001f
C331 B.n291 VSUBS 0.008001f
C332 B.n292 VSUBS 0.008001f
C333 B.n293 VSUBS 0.008001f
C334 B.n294 VSUBS 0.008001f
C335 B.n295 VSUBS 0.008001f
C336 B.n296 VSUBS 0.00753f
C337 B.n297 VSUBS 0.018537f
C338 B.n298 VSUBS 0.004471f
C339 B.n299 VSUBS 0.008001f
C340 B.n300 VSUBS 0.008001f
C341 B.n301 VSUBS 0.008001f
C342 B.n302 VSUBS 0.008001f
C343 B.n303 VSUBS 0.008001f
C344 B.n304 VSUBS 0.008001f
C345 B.n305 VSUBS 0.008001f
C346 B.n306 VSUBS 0.008001f
C347 B.n307 VSUBS 0.008001f
C348 B.n308 VSUBS 0.008001f
C349 B.n309 VSUBS 0.008001f
C350 B.n310 VSUBS 0.008001f
C351 B.n311 VSUBS 0.004471f
C352 B.n312 VSUBS 0.008001f
C353 B.n313 VSUBS 0.008001f
C354 B.n314 VSUBS 0.00753f
C355 B.n315 VSUBS 0.008001f
C356 B.n316 VSUBS 0.008001f
C357 B.n317 VSUBS 0.008001f
C358 B.n318 VSUBS 0.008001f
C359 B.n319 VSUBS 0.008001f
C360 B.n320 VSUBS 0.008001f
C361 B.n321 VSUBS 0.008001f
C362 B.n322 VSUBS 0.008001f
C363 B.n323 VSUBS 0.008001f
C364 B.n324 VSUBS 0.008001f
C365 B.n325 VSUBS 0.008001f
C366 B.n326 VSUBS 0.008001f
C367 B.n327 VSUBS 0.008001f
C368 B.n328 VSUBS 0.008001f
C369 B.n329 VSUBS 0.008001f
C370 B.n330 VSUBS 0.008001f
C371 B.n331 VSUBS 0.008001f
C372 B.n332 VSUBS 0.008001f
C373 B.n333 VSUBS 0.008001f
C374 B.n334 VSUBS 0.008001f
C375 B.n335 VSUBS 0.008001f
C376 B.n336 VSUBS 0.008001f
C377 B.n337 VSUBS 0.008001f
C378 B.n338 VSUBS 0.008001f
C379 B.n339 VSUBS 0.008001f
C380 B.n340 VSUBS 0.008001f
C381 B.n341 VSUBS 0.008001f
C382 B.n342 VSUBS 0.008001f
C383 B.n343 VSUBS 0.008001f
C384 B.n344 VSUBS 0.008001f
C385 B.n345 VSUBS 0.008001f
C386 B.n346 VSUBS 0.008001f
C387 B.n347 VSUBS 0.008001f
C388 B.n348 VSUBS 0.008001f
C389 B.n349 VSUBS 0.008001f
C390 B.n350 VSUBS 0.008001f
C391 B.n351 VSUBS 0.008001f
C392 B.n352 VSUBS 0.008001f
C393 B.n353 VSUBS 0.008001f
C394 B.n354 VSUBS 0.008001f
C395 B.n355 VSUBS 0.008001f
C396 B.n356 VSUBS 0.008001f
C397 B.n357 VSUBS 0.008001f
C398 B.n358 VSUBS 0.008001f
C399 B.n359 VSUBS 0.008001f
C400 B.n360 VSUBS 0.008001f
C401 B.n361 VSUBS 0.008001f
C402 B.n362 VSUBS 0.008001f
C403 B.n363 VSUBS 0.008001f
C404 B.n364 VSUBS 0.008001f
C405 B.n365 VSUBS 0.008001f
C406 B.n366 VSUBS 0.008001f
C407 B.n367 VSUBS 0.008001f
C408 B.n368 VSUBS 0.008001f
C409 B.n369 VSUBS 0.008001f
C410 B.n370 VSUBS 0.008001f
C411 B.n371 VSUBS 0.008001f
C412 B.n372 VSUBS 0.008001f
C413 B.n373 VSUBS 0.008001f
C414 B.n374 VSUBS 0.008001f
C415 B.n375 VSUBS 0.008001f
C416 B.n376 VSUBS 0.008001f
C417 B.n377 VSUBS 0.008001f
C418 B.n378 VSUBS 0.008001f
C419 B.n379 VSUBS 0.008001f
C420 B.n380 VSUBS 0.008001f
C421 B.n381 VSUBS 0.008001f
C422 B.n382 VSUBS 0.008001f
C423 B.n383 VSUBS 0.008001f
C424 B.n384 VSUBS 0.008001f
C425 B.n385 VSUBS 0.008001f
C426 B.n386 VSUBS 0.008001f
C427 B.n387 VSUBS 0.008001f
C428 B.n388 VSUBS 0.008001f
C429 B.n389 VSUBS 0.008001f
C430 B.n390 VSUBS 0.008001f
C431 B.n391 VSUBS 0.008001f
C432 B.n392 VSUBS 0.008001f
C433 B.n393 VSUBS 0.008001f
C434 B.n394 VSUBS 0.008001f
C435 B.n395 VSUBS 0.008001f
C436 B.n396 VSUBS 0.008001f
C437 B.n397 VSUBS 0.008001f
C438 B.n398 VSUBS 0.008001f
C439 B.n399 VSUBS 0.008001f
C440 B.n400 VSUBS 0.008001f
C441 B.n401 VSUBS 0.008001f
C442 B.n402 VSUBS 0.008001f
C443 B.n403 VSUBS 0.008001f
C444 B.n404 VSUBS 0.008001f
C445 B.n405 VSUBS 0.008001f
C446 B.n406 VSUBS 0.008001f
C447 B.n407 VSUBS 0.008001f
C448 B.n408 VSUBS 0.018192f
C449 B.n409 VSUBS 0.017106f
C450 B.n410 VSUBS 0.017106f
C451 B.n411 VSUBS 0.008001f
C452 B.n412 VSUBS 0.008001f
C453 B.n413 VSUBS 0.008001f
C454 B.n414 VSUBS 0.008001f
C455 B.n415 VSUBS 0.008001f
C456 B.n416 VSUBS 0.008001f
C457 B.n417 VSUBS 0.008001f
C458 B.n418 VSUBS 0.008001f
C459 B.n419 VSUBS 0.008001f
C460 B.n420 VSUBS 0.008001f
C461 B.n421 VSUBS 0.008001f
C462 B.n422 VSUBS 0.008001f
C463 B.n423 VSUBS 0.008001f
C464 B.n424 VSUBS 0.008001f
C465 B.n425 VSUBS 0.008001f
C466 B.n426 VSUBS 0.008001f
C467 B.n427 VSUBS 0.008001f
C468 B.n428 VSUBS 0.008001f
C469 B.n429 VSUBS 0.008001f
C470 B.n430 VSUBS 0.008001f
C471 B.n431 VSUBS 0.008001f
C472 B.n432 VSUBS 0.008001f
C473 B.n433 VSUBS 0.008001f
C474 B.n434 VSUBS 0.008001f
C475 B.n435 VSUBS 0.008001f
C476 B.n436 VSUBS 0.008001f
C477 B.n437 VSUBS 0.008001f
C478 B.n438 VSUBS 0.008001f
C479 B.n439 VSUBS 0.008001f
C480 B.n440 VSUBS 0.008001f
C481 B.n441 VSUBS 0.008001f
C482 B.n442 VSUBS 0.008001f
C483 B.n443 VSUBS 0.008001f
C484 B.n444 VSUBS 0.008001f
C485 B.n445 VSUBS 0.008001f
C486 B.n446 VSUBS 0.008001f
C487 B.n447 VSUBS 0.008001f
C488 B.n448 VSUBS 0.008001f
C489 B.n449 VSUBS 0.008001f
C490 B.n450 VSUBS 0.008001f
C491 B.n451 VSUBS 0.008001f
C492 B.n452 VSUBS 0.008001f
C493 B.n453 VSUBS 0.008001f
C494 B.n454 VSUBS 0.018142f
C495 B.n455 VSUBS 0.017106f
C496 B.n456 VSUBS 0.018192f
C497 B.n457 VSUBS 0.008001f
C498 B.n458 VSUBS 0.008001f
C499 B.n459 VSUBS 0.008001f
C500 B.n460 VSUBS 0.008001f
C501 B.n461 VSUBS 0.008001f
C502 B.n462 VSUBS 0.008001f
C503 B.n463 VSUBS 0.008001f
C504 B.n464 VSUBS 0.008001f
C505 B.n465 VSUBS 0.008001f
C506 B.n466 VSUBS 0.008001f
C507 B.n467 VSUBS 0.008001f
C508 B.n468 VSUBS 0.008001f
C509 B.n469 VSUBS 0.008001f
C510 B.n470 VSUBS 0.008001f
C511 B.n471 VSUBS 0.008001f
C512 B.n472 VSUBS 0.008001f
C513 B.n473 VSUBS 0.008001f
C514 B.n474 VSUBS 0.008001f
C515 B.n475 VSUBS 0.008001f
C516 B.n476 VSUBS 0.008001f
C517 B.n477 VSUBS 0.008001f
C518 B.n478 VSUBS 0.008001f
C519 B.n479 VSUBS 0.008001f
C520 B.n480 VSUBS 0.008001f
C521 B.n481 VSUBS 0.008001f
C522 B.n482 VSUBS 0.008001f
C523 B.n483 VSUBS 0.008001f
C524 B.n484 VSUBS 0.008001f
C525 B.n485 VSUBS 0.008001f
C526 B.n486 VSUBS 0.008001f
C527 B.n487 VSUBS 0.008001f
C528 B.n488 VSUBS 0.008001f
C529 B.n489 VSUBS 0.008001f
C530 B.n490 VSUBS 0.008001f
C531 B.n491 VSUBS 0.008001f
C532 B.n492 VSUBS 0.008001f
C533 B.n493 VSUBS 0.008001f
C534 B.n494 VSUBS 0.008001f
C535 B.n495 VSUBS 0.008001f
C536 B.n496 VSUBS 0.008001f
C537 B.n497 VSUBS 0.008001f
C538 B.n498 VSUBS 0.008001f
C539 B.n499 VSUBS 0.008001f
C540 B.n500 VSUBS 0.008001f
C541 B.n501 VSUBS 0.008001f
C542 B.n502 VSUBS 0.008001f
C543 B.n503 VSUBS 0.008001f
C544 B.n504 VSUBS 0.008001f
C545 B.n505 VSUBS 0.008001f
C546 B.n506 VSUBS 0.008001f
C547 B.n507 VSUBS 0.008001f
C548 B.n508 VSUBS 0.008001f
C549 B.n509 VSUBS 0.008001f
C550 B.n510 VSUBS 0.008001f
C551 B.n511 VSUBS 0.008001f
C552 B.n512 VSUBS 0.008001f
C553 B.n513 VSUBS 0.008001f
C554 B.n514 VSUBS 0.008001f
C555 B.n515 VSUBS 0.008001f
C556 B.n516 VSUBS 0.008001f
C557 B.n517 VSUBS 0.008001f
C558 B.n518 VSUBS 0.008001f
C559 B.n519 VSUBS 0.008001f
C560 B.n520 VSUBS 0.008001f
C561 B.n521 VSUBS 0.008001f
C562 B.n522 VSUBS 0.008001f
C563 B.n523 VSUBS 0.008001f
C564 B.n524 VSUBS 0.008001f
C565 B.n525 VSUBS 0.008001f
C566 B.n526 VSUBS 0.008001f
C567 B.n527 VSUBS 0.008001f
C568 B.n528 VSUBS 0.008001f
C569 B.n529 VSUBS 0.008001f
C570 B.n530 VSUBS 0.008001f
C571 B.n531 VSUBS 0.008001f
C572 B.n532 VSUBS 0.008001f
C573 B.n533 VSUBS 0.008001f
C574 B.n534 VSUBS 0.008001f
C575 B.n535 VSUBS 0.008001f
C576 B.n536 VSUBS 0.008001f
C577 B.n537 VSUBS 0.008001f
C578 B.n538 VSUBS 0.008001f
C579 B.n539 VSUBS 0.008001f
C580 B.n540 VSUBS 0.008001f
C581 B.n541 VSUBS 0.008001f
C582 B.n542 VSUBS 0.008001f
C583 B.n543 VSUBS 0.008001f
C584 B.n544 VSUBS 0.008001f
C585 B.n545 VSUBS 0.008001f
C586 B.n546 VSUBS 0.008001f
C587 B.n547 VSUBS 0.008001f
C588 B.n548 VSUBS 0.008001f
C589 B.n549 VSUBS 0.008001f
C590 B.n550 VSUBS 0.00753f
C591 B.n551 VSUBS 0.008001f
C592 B.n552 VSUBS 0.008001f
C593 B.n553 VSUBS 0.008001f
C594 B.n554 VSUBS 0.008001f
C595 B.n555 VSUBS 0.008001f
C596 B.n556 VSUBS 0.008001f
C597 B.n557 VSUBS 0.008001f
C598 B.n558 VSUBS 0.008001f
C599 B.n559 VSUBS 0.008001f
C600 B.n560 VSUBS 0.008001f
C601 B.n561 VSUBS 0.008001f
C602 B.n562 VSUBS 0.008001f
C603 B.n563 VSUBS 0.008001f
C604 B.n564 VSUBS 0.008001f
C605 B.n565 VSUBS 0.008001f
C606 B.n566 VSUBS 0.004471f
C607 B.n567 VSUBS 0.018537f
C608 B.n568 VSUBS 0.00753f
C609 B.n569 VSUBS 0.008001f
C610 B.n570 VSUBS 0.008001f
C611 B.n571 VSUBS 0.008001f
C612 B.n572 VSUBS 0.008001f
C613 B.n573 VSUBS 0.008001f
C614 B.n574 VSUBS 0.008001f
C615 B.n575 VSUBS 0.008001f
C616 B.n576 VSUBS 0.008001f
C617 B.n577 VSUBS 0.008001f
C618 B.n578 VSUBS 0.008001f
C619 B.n579 VSUBS 0.008001f
C620 B.n580 VSUBS 0.008001f
C621 B.n581 VSUBS 0.008001f
C622 B.n582 VSUBS 0.008001f
C623 B.n583 VSUBS 0.008001f
C624 B.n584 VSUBS 0.008001f
C625 B.n585 VSUBS 0.008001f
C626 B.n586 VSUBS 0.008001f
C627 B.n587 VSUBS 0.008001f
C628 B.n588 VSUBS 0.008001f
C629 B.n589 VSUBS 0.008001f
C630 B.n590 VSUBS 0.008001f
C631 B.n591 VSUBS 0.008001f
C632 B.n592 VSUBS 0.008001f
C633 B.n593 VSUBS 0.008001f
C634 B.n594 VSUBS 0.008001f
C635 B.n595 VSUBS 0.008001f
C636 B.n596 VSUBS 0.008001f
C637 B.n597 VSUBS 0.008001f
C638 B.n598 VSUBS 0.008001f
C639 B.n599 VSUBS 0.008001f
C640 B.n600 VSUBS 0.008001f
C641 B.n601 VSUBS 0.008001f
C642 B.n602 VSUBS 0.008001f
C643 B.n603 VSUBS 0.008001f
C644 B.n604 VSUBS 0.008001f
C645 B.n605 VSUBS 0.008001f
C646 B.n606 VSUBS 0.008001f
C647 B.n607 VSUBS 0.008001f
C648 B.n608 VSUBS 0.008001f
C649 B.n609 VSUBS 0.008001f
C650 B.n610 VSUBS 0.008001f
C651 B.n611 VSUBS 0.008001f
C652 B.n612 VSUBS 0.008001f
C653 B.n613 VSUBS 0.008001f
C654 B.n614 VSUBS 0.008001f
C655 B.n615 VSUBS 0.008001f
C656 B.n616 VSUBS 0.008001f
C657 B.n617 VSUBS 0.008001f
C658 B.n618 VSUBS 0.008001f
C659 B.n619 VSUBS 0.008001f
C660 B.n620 VSUBS 0.008001f
C661 B.n621 VSUBS 0.008001f
C662 B.n622 VSUBS 0.008001f
C663 B.n623 VSUBS 0.008001f
C664 B.n624 VSUBS 0.008001f
C665 B.n625 VSUBS 0.008001f
C666 B.n626 VSUBS 0.008001f
C667 B.n627 VSUBS 0.008001f
C668 B.n628 VSUBS 0.008001f
C669 B.n629 VSUBS 0.008001f
C670 B.n630 VSUBS 0.008001f
C671 B.n631 VSUBS 0.008001f
C672 B.n632 VSUBS 0.008001f
C673 B.n633 VSUBS 0.008001f
C674 B.n634 VSUBS 0.008001f
C675 B.n635 VSUBS 0.008001f
C676 B.n636 VSUBS 0.008001f
C677 B.n637 VSUBS 0.008001f
C678 B.n638 VSUBS 0.008001f
C679 B.n639 VSUBS 0.008001f
C680 B.n640 VSUBS 0.008001f
C681 B.n641 VSUBS 0.008001f
C682 B.n642 VSUBS 0.008001f
C683 B.n643 VSUBS 0.008001f
C684 B.n644 VSUBS 0.008001f
C685 B.n645 VSUBS 0.008001f
C686 B.n646 VSUBS 0.008001f
C687 B.n647 VSUBS 0.008001f
C688 B.n648 VSUBS 0.008001f
C689 B.n649 VSUBS 0.008001f
C690 B.n650 VSUBS 0.008001f
C691 B.n651 VSUBS 0.008001f
C692 B.n652 VSUBS 0.008001f
C693 B.n653 VSUBS 0.008001f
C694 B.n654 VSUBS 0.008001f
C695 B.n655 VSUBS 0.008001f
C696 B.n656 VSUBS 0.008001f
C697 B.n657 VSUBS 0.008001f
C698 B.n658 VSUBS 0.008001f
C699 B.n659 VSUBS 0.008001f
C700 B.n660 VSUBS 0.008001f
C701 B.n661 VSUBS 0.008001f
C702 B.n662 VSUBS 0.018192f
C703 B.n663 VSUBS 0.018192f
C704 B.n664 VSUBS 0.017106f
C705 B.n665 VSUBS 0.008001f
C706 B.n666 VSUBS 0.008001f
C707 B.n667 VSUBS 0.008001f
C708 B.n668 VSUBS 0.008001f
C709 B.n669 VSUBS 0.008001f
C710 B.n670 VSUBS 0.008001f
C711 B.n671 VSUBS 0.008001f
C712 B.n672 VSUBS 0.008001f
C713 B.n673 VSUBS 0.008001f
C714 B.n674 VSUBS 0.008001f
C715 B.n675 VSUBS 0.008001f
C716 B.n676 VSUBS 0.008001f
C717 B.n677 VSUBS 0.008001f
C718 B.n678 VSUBS 0.008001f
C719 B.n679 VSUBS 0.008001f
C720 B.n680 VSUBS 0.008001f
C721 B.n681 VSUBS 0.008001f
C722 B.n682 VSUBS 0.008001f
C723 B.n683 VSUBS 0.008001f
C724 B.n684 VSUBS 0.008001f
C725 B.n685 VSUBS 0.008001f
C726 B.n686 VSUBS 0.008001f
C727 B.n687 VSUBS 0.018117f
C728 VDD2.t0 VSUBS 0.481341f
C729 VDD2.t3 VSUBS 0.481341f
C730 VDD2.n0 VSUBS 5.09326f
C731 VDD2.t1 VSUBS 0.481341f
C732 VDD2.t2 VSUBS 0.481341f
C733 VDD2.n1 VSUBS 4.03238f
C734 VDD2.n2 VSUBS 5.37595f
C735 VN.t3 VSUBS 1.62831f
C736 VN.t0 VSUBS 1.62829f
C737 VN.n0 VSUBS 1.2003f
C738 VN.t1 VSUBS 1.62831f
C739 VN.t2 VSUBS 1.62829f
C740 VN.n1 VSUBS 2.46852f
C741 VDD1.t0 VSUBS 0.47802f
C742 VDD1.t3 VSUBS 0.47802f
C743 VDD1.n0 VSUBS 4.00517f
C744 VDD1.t2 VSUBS 0.47802f
C745 VDD1.t1 VSUBS 0.47802f
C746 VDD1.n1 VSUBS 5.09012f
C747 VTAIL.n0 VSUBS 0.026038f
C748 VTAIL.n1 VSUBS 0.023514f
C749 VTAIL.n2 VSUBS 0.012636f
C750 VTAIL.n3 VSUBS 0.029866f
C751 VTAIL.n4 VSUBS 0.013379f
C752 VTAIL.n5 VSUBS 0.023514f
C753 VTAIL.n6 VSUBS 0.012636f
C754 VTAIL.n7 VSUBS 0.029866f
C755 VTAIL.n8 VSUBS 0.013379f
C756 VTAIL.n9 VSUBS 0.023514f
C757 VTAIL.n10 VSUBS 0.012636f
C758 VTAIL.n11 VSUBS 0.029866f
C759 VTAIL.n12 VSUBS 0.013007f
C760 VTAIL.n13 VSUBS 0.023514f
C761 VTAIL.n14 VSUBS 0.013379f
C762 VTAIL.n15 VSUBS 0.029866f
C763 VTAIL.n16 VSUBS 0.013379f
C764 VTAIL.n17 VSUBS 0.023514f
C765 VTAIL.n18 VSUBS 0.012636f
C766 VTAIL.n19 VSUBS 0.029866f
C767 VTAIL.n20 VSUBS 0.013379f
C768 VTAIL.n21 VSUBS 0.023514f
C769 VTAIL.n22 VSUBS 0.012636f
C770 VTAIL.n23 VSUBS 0.029866f
C771 VTAIL.n24 VSUBS 0.013379f
C772 VTAIL.n25 VSUBS 0.023514f
C773 VTAIL.n26 VSUBS 0.012636f
C774 VTAIL.n27 VSUBS 0.029866f
C775 VTAIL.n28 VSUBS 0.013379f
C776 VTAIL.n29 VSUBS 0.023514f
C777 VTAIL.n30 VSUBS 0.012636f
C778 VTAIL.n31 VSUBS 0.029866f
C779 VTAIL.n32 VSUBS 0.013379f
C780 VTAIL.n33 VSUBS 1.9957f
C781 VTAIL.n34 VSUBS 0.012636f
C782 VTAIL.t0 VSUBS 0.064208f
C783 VTAIL.n35 VSUBS 0.19787f
C784 VTAIL.n36 VSUBS 0.019f
C785 VTAIL.n37 VSUBS 0.0224f
C786 VTAIL.n38 VSUBS 0.029866f
C787 VTAIL.n39 VSUBS 0.013379f
C788 VTAIL.n40 VSUBS 0.012636f
C789 VTAIL.n41 VSUBS 0.023514f
C790 VTAIL.n42 VSUBS 0.023514f
C791 VTAIL.n43 VSUBS 0.012636f
C792 VTAIL.n44 VSUBS 0.013379f
C793 VTAIL.n45 VSUBS 0.029866f
C794 VTAIL.n46 VSUBS 0.029866f
C795 VTAIL.n47 VSUBS 0.013379f
C796 VTAIL.n48 VSUBS 0.012636f
C797 VTAIL.n49 VSUBS 0.023514f
C798 VTAIL.n50 VSUBS 0.023514f
C799 VTAIL.n51 VSUBS 0.012636f
C800 VTAIL.n52 VSUBS 0.013379f
C801 VTAIL.n53 VSUBS 0.029866f
C802 VTAIL.n54 VSUBS 0.029866f
C803 VTAIL.n55 VSUBS 0.013379f
C804 VTAIL.n56 VSUBS 0.012636f
C805 VTAIL.n57 VSUBS 0.023514f
C806 VTAIL.n58 VSUBS 0.023514f
C807 VTAIL.n59 VSUBS 0.012636f
C808 VTAIL.n60 VSUBS 0.013379f
C809 VTAIL.n61 VSUBS 0.029866f
C810 VTAIL.n62 VSUBS 0.029866f
C811 VTAIL.n63 VSUBS 0.013379f
C812 VTAIL.n64 VSUBS 0.012636f
C813 VTAIL.n65 VSUBS 0.023514f
C814 VTAIL.n66 VSUBS 0.023514f
C815 VTAIL.n67 VSUBS 0.012636f
C816 VTAIL.n68 VSUBS 0.013379f
C817 VTAIL.n69 VSUBS 0.029866f
C818 VTAIL.n70 VSUBS 0.029866f
C819 VTAIL.n71 VSUBS 0.013379f
C820 VTAIL.n72 VSUBS 0.012636f
C821 VTAIL.n73 VSUBS 0.023514f
C822 VTAIL.n74 VSUBS 0.023514f
C823 VTAIL.n75 VSUBS 0.012636f
C824 VTAIL.n76 VSUBS 0.012636f
C825 VTAIL.n77 VSUBS 0.013379f
C826 VTAIL.n78 VSUBS 0.029866f
C827 VTAIL.n79 VSUBS 0.029866f
C828 VTAIL.n80 VSUBS 0.029866f
C829 VTAIL.n81 VSUBS 0.013007f
C830 VTAIL.n82 VSUBS 0.012636f
C831 VTAIL.n83 VSUBS 0.023514f
C832 VTAIL.n84 VSUBS 0.023514f
C833 VTAIL.n85 VSUBS 0.012636f
C834 VTAIL.n86 VSUBS 0.013379f
C835 VTAIL.n87 VSUBS 0.029866f
C836 VTAIL.n88 VSUBS 0.029866f
C837 VTAIL.n89 VSUBS 0.013379f
C838 VTAIL.n90 VSUBS 0.012636f
C839 VTAIL.n91 VSUBS 0.023514f
C840 VTAIL.n92 VSUBS 0.023514f
C841 VTAIL.n93 VSUBS 0.012636f
C842 VTAIL.n94 VSUBS 0.013379f
C843 VTAIL.n95 VSUBS 0.029866f
C844 VTAIL.n96 VSUBS 0.029866f
C845 VTAIL.n97 VSUBS 0.013379f
C846 VTAIL.n98 VSUBS 0.012636f
C847 VTAIL.n99 VSUBS 0.023514f
C848 VTAIL.n100 VSUBS 0.023514f
C849 VTAIL.n101 VSUBS 0.012636f
C850 VTAIL.n102 VSUBS 0.013379f
C851 VTAIL.n103 VSUBS 0.029866f
C852 VTAIL.n104 VSUBS 0.072987f
C853 VTAIL.n105 VSUBS 0.013379f
C854 VTAIL.n106 VSUBS 0.012636f
C855 VTAIL.n107 VSUBS 0.052747f
C856 VTAIL.n108 VSUBS 0.036685f
C857 VTAIL.n109 VSUBS 0.084332f
C858 VTAIL.n110 VSUBS 0.026038f
C859 VTAIL.n111 VSUBS 0.023514f
C860 VTAIL.n112 VSUBS 0.012636f
C861 VTAIL.n113 VSUBS 0.029866f
C862 VTAIL.n114 VSUBS 0.013379f
C863 VTAIL.n115 VSUBS 0.023514f
C864 VTAIL.n116 VSUBS 0.012636f
C865 VTAIL.n117 VSUBS 0.029866f
C866 VTAIL.n118 VSUBS 0.013379f
C867 VTAIL.n119 VSUBS 0.023514f
C868 VTAIL.n120 VSUBS 0.012636f
C869 VTAIL.n121 VSUBS 0.029866f
C870 VTAIL.n122 VSUBS 0.013007f
C871 VTAIL.n123 VSUBS 0.023514f
C872 VTAIL.n124 VSUBS 0.013379f
C873 VTAIL.n125 VSUBS 0.029866f
C874 VTAIL.n126 VSUBS 0.013379f
C875 VTAIL.n127 VSUBS 0.023514f
C876 VTAIL.n128 VSUBS 0.012636f
C877 VTAIL.n129 VSUBS 0.029866f
C878 VTAIL.n130 VSUBS 0.013379f
C879 VTAIL.n131 VSUBS 0.023514f
C880 VTAIL.n132 VSUBS 0.012636f
C881 VTAIL.n133 VSUBS 0.029866f
C882 VTAIL.n134 VSUBS 0.013379f
C883 VTAIL.n135 VSUBS 0.023514f
C884 VTAIL.n136 VSUBS 0.012636f
C885 VTAIL.n137 VSUBS 0.029866f
C886 VTAIL.n138 VSUBS 0.013379f
C887 VTAIL.n139 VSUBS 0.023514f
C888 VTAIL.n140 VSUBS 0.012636f
C889 VTAIL.n141 VSUBS 0.029866f
C890 VTAIL.n142 VSUBS 0.013379f
C891 VTAIL.n143 VSUBS 1.9957f
C892 VTAIL.n144 VSUBS 0.012636f
C893 VTAIL.t7 VSUBS 0.064208f
C894 VTAIL.n145 VSUBS 0.19787f
C895 VTAIL.n146 VSUBS 0.019f
C896 VTAIL.n147 VSUBS 0.0224f
C897 VTAIL.n148 VSUBS 0.029866f
C898 VTAIL.n149 VSUBS 0.013379f
C899 VTAIL.n150 VSUBS 0.012636f
C900 VTAIL.n151 VSUBS 0.023514f
C901 VTAIL.n152 VSUBS 0.023514f
C902 VTAIL.n153 VSUBS 0.012636f
C903 VTAIL.n154 VSUBS 0.013379f
C904 VTAIL.n155 VSUBS 0.029866f
C905 VTAIL.n156 VSUBS 0.029866f
C906 VTAIL.n157 VSUBS 0.013379f
C907 VTAIL.n158 VSUBS 0.012636f
C908 VTAIL.n159 VSUBS 0.023514f
C909 VTAIL.n160 VSUBS 0.023514f
C910 VTAIL.n161 VSUBS 0.012636f
C911 VTAIL.n162 VSUBS 0.013379f
C912 VTAIL.n163 VSUBS 0.029866f
C913 VTAIL.n164 VSUBS 0.029866f
C914 VTAIL.n165 VSUBS 0.013379f
C915 VTAIL.n166 VSUBS 0.012636f
C916 VTAIL.n167 VSUBS 0.023514f
C917 VTAIL.n168 VSUBS 0.023514f
C918 VTAIL.n169 VSUBS 0.012636f
C919 VTAIL.n170 VSUBS 0.013379f
C920 VTAIL.n171 VSUBS 0.029866f
C921 VTAIL.n172 VSUBS 0.029866f
C922 VTAIL.n173 VSUBS 0.013379f
C923 VTAIL.n174 VSUBS 0.012636f
C924 VTAIL.n175 VSUBS 0.023514f
C925 VTAIL.n176 VSUBS 0.023514f
C926 VTAIL.n177 VSUBS 0.012636f
C927 VTAIL.n178 VSUBS 0.013379f
C928 VTAIL.n179 VSUBS 0.029866f
C929 VTAIL.n180 VSUBS 0.029866f
C930 VTAIL.n181 VSUBS 0.013379f
C931 VTAIL.n182 VSUBS 0.012636f
C932 VTAIL.n183 VSUBS 0.023514f
C933 VTAIL.n184 VSUBS 0.023514f
C934 VTAIL.n185 VSUBS 0.012636f
C935 VTAIL.n186 VSUBS 0.012636f
C936 VTAIL.n187 VSUBS 0.013379f
C937 VTAIL.n188 VSUBS 0.029866f
C938 VTAIL.n189 VSUBS 0.029866f
C939 VTAIL.n190 VSUBS 0.029866f
C940 VTAIL.n191 VSUBS 0.013007f
C941 VTAIL.n192 VSUBS 0.012636f
C942 VTAIL.n193 VSUBS 0.023514f
C943 VTAIL.n194 VSUBS 0.023514f
C944 VTAIL.n195 VSUBS 0.012636f
C945 VTAIL.n196 VSUBS 0.013379f
C946 VTAIL.n197 VSUBS 0.029866f
C947 VTAIL.n198 VSUBS 0.029866f
C948 VTAIL.n199 VSUBS 0.013379f
C949 VTAIL.n200 VSUBS 0.012636f
C950 VTAIL.n201 VSUBS 0.023514f
C951 VTAIL.n202 VSUBS 0.023514f
C952 VTAIL.n203 VSUBS 0.012636f
C953 VTAIL.n204 VSUBS 0.013379f
C954 VTAIL.n205 VSUBS 0.029866f
C955 VTAIL.n206 VSUBS 0.029866f
C956 VTAIL.n207 VSUBS 0.013379f
C957 VTAIL.n208 VSUBS 0.012636f
C958 VTAIL.n209 VSUBS 0.023514f
C959 VTAIL.n210 VSUBS 0.023514f
C960 VTAIL.n211 VSUBS 0.012636f
C961 VTAIL.n212 VSUBS 0.013379f
C962 VTAIL.n213 VSUBS 0.029866f
C963 VTAIL.n214 VSUBS 0.072987f
C964 VTAIL.n215 VSUBS 0.013379f
C965 VTAIL.n216 VSUBS 0.012636f
C966 VTAIL.n217 VSUBS 0.052747f
C967 VTAIL.n218 VSUBS 0.036685f
C968 VTAIL.n219 VSUBS 0.105071f
C969 VTAIL.n220 VSUBS 0.026038f
C970 VTAIL.n221 VSUBS 0.023514f
C971 VTAIL.n222 VSUBS 0.012636f
C972 VTAIL.n223 VSUBS 0.029866f
C973 VTAIL.n224 VSUBS 0.013379f
C974 VTAIL.n225 VSUBS 0.023514f
C975 VTAIL.n226 VSUBS 0.012636f
C976 VTAIL.n227 VSUBS 0.029866f
C977 VTAIL.n228 VSUBS 0.013379f
C978 VTAIL.n229 VSUBS 0.023514f
C979 VTAIL.n230 VSUBS 0.012636f
C980 VTAIL.n231 VSUBS 0.029866f
C981 VTAIL.n232 VSUBS 0.013007f
C982 VTAIL.n233 VSUBS 0.023514f
C983 VTAIL.n234 VSUBS 0.013379f
C984 VTAIL.n235 VSUBS 0.029866f
C985 VTAIL.n236 VSUBS 0.013379f
C986 VTAIL.n237 VSUBS 0.023514f
C987 VTAIL.n238 VSUBS 0.012636f
C988 VTAIL.n239 VSUBS 0.029866f
C989 VTAIL.n240 VSUBS 0.013379f
C990 VTAIL.n241 VSUBS 0.023514f
C991 VTAIL.n242 VSUBS 0.012636f
C992 VTAIL.n243 VSUBS 0.029866f
C993 VTAIL.n244 VSUBS 0.013379f
C994 VTAIL.n245 VSUBS 0.023514f
C995 VTAIL.n246 VSUBS 0.012636f
C996 VTAIL.n247 VSUBS 0.029866f
C997 VTAIL.n248 VSUBS 0.013379f
C998 VTAIL.n249 VSUBS 0.023514f
C999 VTAIL.n250 VSUBS 0.012636f
C1000 VTAIL.n251 VSUBS 0.029866f
C1001 VTAIL.n252 VSUBS 0.013379f
C1002 VTAIL.n253 VSUBS 1.9957f
C1003 VTAIL.n254 VSUBS 0.012636f
C1004 VTAIL.t6 VSUBS 0.064208f
C1005 VTAIL.n255 VSUBS 0.19787f
C1006 VTAIL.n256 VSUBS 0.019f
C1007 VTAIL.n257 VSUBS 0.0224f
C1008 VTAIL.n258 VSUBS 0.029866f
C1009 VTAIL.n259 VSUBS 0.013379f
C1010 VTAIL.n260 VSUBS 0.012636f
C1011 VTAIL.n261 VSUBS 0.023514f
C1012 VTAIL.n262 VSUBS 0.023514f
C1013 VTAIL.n263 VSUBS 0.012636f
C1014 VTAIL.n264 VSUBS 0.013379f
C1015 VTAIL.n265 VSUBS 0.029866f
C1016 VTAIL.n266 VSUBS 0.029866f
C1017 VTAIL.n267 VSUBS 0.013379f
C1018 VTAIL.n268 VSUBS 0.012636f
C1019 VTAIL.n269 VSUBS 0.023514f
C1020 VTAIL.n270 VSUBS 0.023514f
C1021 VTAIL.n271 VSUBS 0.012636f
C1022 VTAIL.n272 VSUBS 0.013379f
C1023 VTAIL.n273 VSUBS 0.029866f
C1024 VTAIL.n274 VSUBS 0.029866f
C1025 VTAIL.n275 VSUBS 0.013379f
C1026 VTAIL.n276 VSUBS 0.012636f
C1027 VTAIL.n277 VSUBS 0.023514f
C1028 VTAIL.n278 VSUBS 0.023514f
C1029 VTAIL.n279 VSUBS 0.012636f
C1030 VTAIL.n280 VSUBS 0.013379f
C1031 VTAIL.n281 VSUBS 0.029866f
C1032 VTAIL.n282 VSUBS 0.029866f
C1033 VTAIL.n283 VSUBS 0.013379f
C1034 VTAIL.n284 VSUBS 0.012636f
C1035 VTAIL.n285 VSUBS 0.023514f
C1036 VTAIL.n286 VSUBS 0.023514f
C1037 VTAIL.n287 VSUBS 0.012636f
C1038 VTAIL.n288 VSUBS 0.013379f
C1039 VTAIL.n289 VSUBS 0.029866f
C1040 VTAIL.n290 VSUBS 0.029866f
C1041 VTAIL.n291 VSUBS 0.013379f
C1042 VTAIL.n292 VSUBS 0.012636f
C1043 VTAIL.n293 VSUBS 0.023514f
C1044 VTAIL.n294 VSUBS 0.023514f
C1045 VTAIL.n295 VSUBS 0.012636f
C1046 VTAIL.n296 VSUBS 0.012636f
C1047 VTAIL.n297 VSUBS 0.013379f
C1048 VTAIL.n298 VSUBS 0.029866f
C1049 VTAIL.n299 VSUBS 0.029866f
C1050 VTAIL.n300 VSUBS 0.029866f
C1051 VTAIL.n301 VSUBS 0.013007f
C1052 VTAIL.n302 VSUBS 0.012636f
C1053 VTAIL.n303 VSUBS 0.023514f
C1054 VTAIL.n304 VSUBS 0.023514f
C1055 VTAIL.n305 VSUBS 0.012636f
C1056 VTAIL.n306 VSUBS 0.013379f
C1057 VTAIL.n307 VSUBS 0.029866f
C1058 VTAIL.n308 VSUBS 0.029866f
C1059 VTAIL.n309 VSUBS 0.013379f
C1060 VTAIL.n310 VSUBS 0.012636f
C1061 VTAIL.n311 VSUBS 0.023514f
C1062 VTAIL.n312 VSUBS 0.023514f
C1063 VTAIL.n313 VSUBS 0.012636f
C1064 VTAIL.n314 VSUBS 0.013379f
C1065 VTAIL.n315 VSUBS 0.029866f
C1066 VTAIL.n316 VSUBS 0.029866f
C1067 VTAIL.n317 VSUBS 0.013379f
C1068 VTAIL.n318 VSUBS 0.012636f
C1069 VTAIL.n319 VSUBS 0.023514f
C1070 VTAIL.n320 VSUBS 0.023514f
C1071 VTAIL.n321 VSUBS 0.012636f
C1072 VTAIL.n322 VSUBS 0.013379f
C1073 VTAIL.n323 VSUBS 0.029866f
C1074 VTAIL.n324 VSUBS 0.072987f
C1075 VTAIL.n325 VSUBS 0.013379f
C1076 VTAIL.n326 VSUBS 0.012636f
C1077 VTAIL.n327 VSUBS 0.052747f
C1078 VTAIL.n328 VSUBS 0.036685f
C1079 VTAIL.n329 VSUBS 1.72138f
C1080 VTAIL.n330 VSUBS 0.026038f
C1081 VTAIL.n331 VSUBS 0.023514f
C1082 VTAIL.n332 VSUBS 0.012636f
C1083 VTAIL.n333 VSUBS 0.029866f
C1084 VTAIL.n334 VSUBS 0.013379f
C1085 VTAIL.n335 VSUBS 0.023514f
C1086 VTAIL.n336 VSUBS 0.012636f
C1087 VTAIL.n337 VSUBS 0.029866f
C1088 VTAIL.n338 VSUBS 0.013379f
C1089 VTAIL.n339 VSUBS 0.023514f
C1090 VTAIL.n340 VSUBS 0.012636f
C1091 VTAIL.n341 VSUBS 0.029866f
C1092 VTAIL.n342 VSUBS 0.013007f
C1093 VTAIL.n343 VSUBS 0.023514f
C1094 VTAIL.n344 VSUBS 0.013007f
C1095 VTAIL.n345 VSUBS 0.012636f
C1096 VTAIL.n346 VSUBS 0.029866f
C1097 VTAIL.n347 VSUBS 0.029866f
C1098 VTAIL.n348 VSUBS 0.013379f
C1099 VTAIL.n349 VSUBS 0.023514f
C1100 VTAIL.n350 VSUBS 0.012636f
C1101 VTAIL.n351 VSUBS 0.029866f
C1102 VTAIL.n352 VSUBS 0.013379f
C1103 VTAIL.n353 VSUBS 0.023514f
C1104 VTAIL.n354 VSUBS 0.012636f
C1105 VTAIL.n355 VSUBS 0.029866f
C1106 VTAIL.n356 VSUBS 0.013379f
C1107 VTAIL.n357 VSUBS 0.023514f
C1108 VTAIL.n358 VSUBS 0.012636f
C1109 VTAIL.n359 VSUBS 0.029866f
C1110 VTAIL.n360 VSUBS 0.013379f
C1111 VTAIL.n361 VSUBS 0.023514f
C1112 VTAIL.n362 VSUBS 0.012636f
C1113 VTAIL.n363 VSUBS 0.029866f
C1114 VTAIL.n364 VSUBS 0.013379f
C1115 VTAIL.n365 VSUBS 1.9957f
C1116 VTAIL.n366 VSUBS 0.012636f
C1117 VTAIL.t3 VSUBS 0.064208f
C1118 VTAIL.n367 VSUBS 0.19787f
C1119 VTAIL.n368 VSUBS 0.019f
C1120 VTAIL.n369 VSUBS 0.0224f
C1121 VTAIL.n370 VSUBS 0.029866f
C1122 VTAIL.n371 VSUBS 0.013379f
C1123 VTAIL.n372 VSUBS 0.012636f
C1124 VTAIL.n373 VSUBS 0.023514f
C1125 VTAIL.n374 VSUBS 0.023514f
C1126 VTAIL.n375 VSUBS 0.012636f
C1127 VTAIL.n376 VSUBS 0.013379f
C1128 VTAIL.n377 VSUBS 0.029866f
C1129 VTAIL.n378 VSUBS 0.029866f
C1130 VTAIL.n379 VSUBS 0.013379f
C1131 VTAIL.n380 VSUBS 0.012636f
C1132 VTAIL.n381 VSUBS 0.023514f
C1133 VTAIL.n382 VSUBS 0.023514f
C1134 VTAIL.n383 VSUBS 0.012636f
C1135 VTAIL.n384 VSUBS 0.013379f
C1136 VTAIL.n385 VSUBS 0.029866f
C1137 VTAIL.n386 VSUBS 0.029866f
C1138 VTAIL.n387 VSUBS 0.013379f
C1139 VTAIL.n388 VSUBS 0.012636f
C1140 VTAIL.n389 VSUBS 0.023514f
C1141 VTAIL.n390 VSUBS 0.023514f
C1142 VTAIL.n391 VSUBS 0.012636f
C1143 VTAIL.n392 VSUBS 0.013379f
C1144 VTAIL.n393 VSUBS 0.029866f
C1145 VTAIL.n394 VSUBS 0.029866f
C1146 VTAIL.n395 VSUBS 0.013379f
C1147 VTAIL.n396 VSUBS 0.012636f
C1148 VTAIL.n397 VSUBS 0.023514f
C1149 VTAIL.n398 VSUBS 0.023514f
C1150 VTAIL.n399 VSUBS 0.012636f
C1151 VTAIL.n400 VSUBS 0.013379f
C1152 VTAIL.n401 VSUBS 0.029866f
C1153 VTAIL.n402 VSUBS 0.029866f
C1154 VTAIL.n403 VSUBS 0.013379f
C1155 VTAIL.n404 VSUBS 0.012636f
C1156 VTAIL.n405 VSUBS 0.023514f
C1157 VTAIL.n406 VSUBS 0.023514f
C1158 VTAIL.n407 VSUBS 0.012636f
C1159 VTAIL.n408 VSUBS 0.013379f
C1160 VTAIL.n409 VSUBS 0.029866f
C1161 VTAIL.n410 VSUBS 0.029866f
C1162 VTAIL.n411 VSUBS 0.013379f
C1163 VTAIL.n412 VSUBS 0.012636f
C1164 VTAIL.n413 VSUBS 0.023514f
C1165 VTAIL.n414 VSUBS 0.023514f
C1166 VTAIL.n415 VSUBS 0.012636f
C1167 VTAIL.n416 VSUBS 0.013379f
C1168 VTAIL.n417 VSUBS 0.029866f
C1169 VTAIL.n418 VSUBS 0.029866f
C1170 VTAIL.n419 VSUBS 0.013379f
C1171 VTAIL.n420 VSUBS 0.012636f
C1172 VTAIL.n421 VSUBS 0.023514f
C1173 VTAIL.n422 VSUBS 0.023514f
C1174 VTAIL.n423 VSUBS 0.012636f
C1175 VTAIL.n424 VSUBS 0.013379f
C1176 VTAIL.n425 VSUBS 0.029866f
C1177 VTAIL.n426 VSUBS 0.029866f
C1178 VTAIL.n427 VSUBS 0.013379f
C1179 VTAIL.n428 VSUBS 0.012636f
C1180 VTAIL.n429 VSUBS 0.023514f
C1181 VTAIL.n430 VSUBS 0.023514f
C1182 VTAIL.n431 VSUBS 0.012636f
C1183 VTAIL.n432 VSUBS 0.013379f
C1184 VTAIL.n433 VSUBS 0.029866f
C1185 VTAIL.n434 VSUBS 0.072987f
C1186 VTAIL.n435 VSUBS 0.013379f
C1187 VTAIL.n436 VSUBS 0.012636f
C1188 VTAIL.n437 VSUBS 0.052747f
C1189 VTAIL.n438 VSUBS 0.036685f
C1190 VTAIL.n439 VSUBS 1.72138f
C1191 VTAIL.n440 VSUBS 0.026038f
C1192 VTAIL.n441 VSUBS 0.023514f
C1193 VTAIL.n442 VSUBS 0.012636f
C1194 VTAIL.n443 VSUBS 0.029866f
C1195 VTAIL.n444 VSUBS 0.013379f
C1196 VTAIL.n445 VSUBS 0.023514f
C1197 VTAIL.n446 VSUBS 0.012636f
C1198 VTAIL.n447 VSUBS 0.029866f
C1199 VTAIL.n448 VSUBS 0.013379f
C1200 VTAIL.n449 VSUBS 0.023514f
C1201 VTAIL.n450 VSUBS 0.012636f
C1202 VTAIL.n451 VSUBS 0.029866f
C1203 VTAIL.n452 VSUBS 0.013007f
C1204 VTAIL.n453 VSUBS 0.023514f
C1205 VTAIL.n454 VSUBS 0.013007f
C1206 VTAIL.n455 VSUBS 0.012636f
C1207 VTAIL.n456 VSUBS 0.029866f
C1208 VTAIL.n457 VSUBS 0.029866f
C1209 VTAIL.n458 VSUBS 0.013379f
C1210 VTAIL.n459 VSUBS 0.023514f
C1211 VTAIL.n460 VSUBS 0.012636f
C1212 VTAIL.n461 VSUBS 0.029866f
C1213 VTAIL.n462 VSUBS 0.013379f
C1214 VTAIL.n463 VSUBS 0.023514f
C1215 VTAIL.n464 VSUBS 0.012636f
C1216 VTAIL.n465 VSUBS 0.029866f
C1217 VTAIL.n466 VSUBS 0.013379f
C1218 VTAIL.n467 VSUBS 0.023514f
C1219 VTAIL.n468 VSUBS 0.012636f
C1220 VTAIL.n469 VSUBS 0.029866f
C1221 VTAIL.n470 VSUBS 0.013379f
C1222 VTAIL.n471 VSUBS 0.023514f
C1223 VTAIL.n472 VSUBS 0.012636f
C1224 VTAIL.n473 VSUBS 0.029866f
C1225 VTAIL.n474 VSUBS 0.013379f
C1226 VTAIL.n475 VSUBS 1.9957f
C1227 VTAIL.n476 VSUBS 0.012636f
C1228 VTAIL.t2 VSUBS 0.064208f
C1229 VTAIL.n477 VSUBS 0.19787f
C1230 VTAIL.n478 VSUBS 0.019f
C1231 VTAIL.n479 VSUBS 0.0224f
C1232 VTAIL.n480 VSUBS 0.029866f
C1233 VTAIL.n481 VSUBS 0.013379f
C1234 VTAIL.n482 VSUBS 0.012636f
C1235 VTAIL.n483 VSUBS 0.023514f
C1236 VTAIL.n484 VSUBS 0.023514f
C1237 VTAIL.n485 VSUBS 0.012636f
C1238 VTAIL.n486 VSUBS 0.013379f
C1239 VTAIL.n487 VSUBS 0.029866f
C1240 VTAIL.n488 VSUBS 0.029866f
C1241 VTAIL.n489 VSUBS 0.013379f
C1242 VTAIL.n490 VSUBS 0.012636f
C1243 VTAIL.n491 VSUBS 0.023514f
C1244 VTAIL.n492 VSUBS 0.023514f
C1245 VTAIL.n493 VSUBS 0.012636f
C1246 VTAIL.n494 VSUBS 0.013379f
C1247 VTAIL.n495 VSUBS 0.029866f
C1248 VTAIL.n496 VSUBS 0.029866f
C1249 VTAIL.n497 VSUBS 0.013379f
C1250 VTAIL.n498 VSUBS 0.012636f
C1251 VTAIL.n499 VSUBS 0.023514f
C1252 VTAIL.n500 VSUBS 0.023514f
C1253 VTAIL.n501 VSUBS 0.012636f
C1254 VTAIL.n502 VSUBS 0.013379f
C1255 VTAIL.n503 VSUBS 0.029866f
C1256 VTAIL.n504 VSUBS 0.029866f
C1257 VTAIL.n505 VSUBS 0.013379f
C1258 VTAIL.n506 VSUBS 0.012636f
C1259 VTAIL.n507 VSUBS 0.023514f
C1260 VTAIL.n508 VSUBS 0.023514f
C1261 VTAIL.n509 VSUBS 0.012636f
C1262 VTAIL.n510 VSUBS 0.013379f
C1263 VTAIL.n511 VSUBS 0.029866f
C1264 VTAIL.n512 VSUBS 0.029866f
C1265 VTAIL.n513 VSUBS 0.013379f
C1266 VTAIL.n514 VSUBS 0.012636f
C1267 VTAIL.n515 VSUBS 0.023514f
C1268 VTAIL.n516 VSUBS 0.023514f
C1269 VTAIL.n517 VSUBS 0.012636f
C1270 VTAIL.n518 VSUBS 0.013379f
C1271 VTAIL.n519 VSUBS 0.029866f
C1272 VTAIL.n520 VSUBS 0.029866f
C1273 VTAIL.n521 VSUBS 0.013379f
C1274 VTAIL.n522 VSUBS 0.012636f
C1275 VTAIL.n523 VSUBS 0.023514f
C1276 VTAIL.n524 VSUBS 0.023514f
C1277 VTAIL.n525 VSUBS 0.012636f
C1278 VTAIL.n526 VSUBS 0.013379f
C1279 VTAIL.n527 VSUBS 0.029866f
C1280 VTAIL.n528 VSUBS 0.029866f
C1281 VTAIL.n529 VSUBS 0.013379f
C1282 VTAIL.n530 VSUBS 0.012636f
C1283 VTAIL.n531 VSUBS 0.023514f
C1284 VTAIL.n532 VSUBS 0.023514f
C1285 VTAIL.n533 VSUBS 0.012636f
C1286 VTAIL.n534 VSUBS 0.013379f
C1287 VTAIL.n535 VSUBS 0.029866f
C1288 VTAIL.n536 VSUBS 0.029866f
C1289 VTAIL.n537 VSUBS 0.013379f
C1290 VTAIL.n538 VSUBS 0.012636f
C1291 VTAIL.n539 VSUBS 0.023514f
C1292 VTAIL.n540 VSUBS 0.023514f
C1293 VTAIL.n541 VSUBS 0.012636f
C1294 VTAIL.n542 VSUBS 0.013379f
C1295 VTAIL.n543 VSUBS 0.029866f
C1296 VTAIL.n544 VSUBS 0.072987f
C1297 VTAIL.n545 VSUBS 0.013379f
C1298 VTAIL.n546 VSUBS 0.012636f
C1299 VTAIL.n547 VSUBS 0.052747f
C1300 VTAIL.n548 VSUBS 0.036685f
C1301 VTAIL.n549 VSUBS 0.105071f
C1302 VTAIL.n550 VSUBS 0.026038f
C1303 VTAIL.n551 VSUBS 0.023514f
C1304 VTAIL.n552 VSUBS 0.012636f
C1305 VTAIL.n553 VSUBS 0.029866f
C1306 VTAIL.n554 VSUBS 0.013379f
C1307 VTAIL.n555 VSUBS 0.023514f
C1308 VTAIL.n556 VSUBS 0.012636f
C1309 VTAIL.n557 VSUBS 0.029866f
C1310 VTAIL.n558 VSUBS 0.013379f
C1311 VTAIL.n559 VSUBS 0.023514f
C1312 VTAIL.n560 VSUBS 0.012636f
C1313 VTAIL.n561 VSUBS 0.029866f
C1314 VTAIL.n562 VSUBS 0.013007f
C1315 VTAIL.n563 VSUBS 0.023514f
C1316 VTAIL.n564 VSUBS 0.013007f
C1317 VTAIL.n565 VSUBS 0.012636f
C1318 VTAIL.n566 VSUBS 0.029866f
C1319 VTAIL.n567 VSUBS 0.029866f
C1320 VTAIL.n568 VSUBS 0.013379f
C1321 VTAIL.n569 VSUBS 0.023514f
C1322 VTAIL.n570 VSUBS 0.012636f
C1323 VTAIL.n571 VSUBS 0.029866f
C1324 VTAIL.n572 VSUBS 0.013379f
C1325 VTAIL.n573 VSUBS 0.023514f
C1326 VTAIL.n574 VSUBS 0.012636f
C1327 VTAIL.n575 VSUBS 0.029866f
C1328 VTAIL.n576 VSUBS 0.013379f
C1329 VTAIL.n577 VSUBS 0.023514f
C1330 VTAIL.n578 VSUBS 0.012636f
C1331 VTAIL.n579 VSUBS 0.029866f
C1332 VTAIL.n580 VSUBS 0.013379f
C1333 VTAIL.n581 VSUBS 0.023514f
C1334 VTAIL.n582 VSUBS 0.012636f
C1335 VTAIL.n583 VSUBS 0.029866f
C1336 VTAIL.n584 VSUBS 0.013379f
C1337 VTAIL.n585 VSUBS 1.9957f
C1338 VTAIL.n586 VSUBS 0.012636f
C1339 VTAIL.t5 VSUBS 0.064208f
C1340 VTAIL.n587 VSUBS 0.19787f
C1341 VTAIL.n588 VSUBS 0.019f
C1342 VTAIL.n589 VSUBS 0.0224f
C1343 VTAIL.n590 VSUBS 0.029866f
C1344 VTAIL.n591 VSUBS 0.013379f
C1345 VTAIL.n592 VSUBS 0.012636f
C1346 VTAIL.n593 VSUBS 0.023514f
C1347 VTAIL.n594 VSUBS 0.023514f
C1348 VTAIL.n595 VSUBS 0.012636f
C1349 VTAIL.n596 VSUBS 0.013379f
C1350 VTAIL.n597 VSUBS 0.029866f
C1351 VTAIL.n598 VSUBS 0.029866f
C1352 VTAIL.n599 VSUBS 0.013379f
C1353 VTAIL.n600 VSUBS 0.012636f
C1354 VTAIL.n601 VSUBS 0.023514f
C1355 VTAIL.n602 VSUBS 0.023514f
C1356 VTAIL.n603 VSUBS 0.012636f
C1357 VTAIL.n604 VSUBS 0.013379f
C1358 VTAIL.n605 VSUBS 0.029866f
C1359 VTAIL.n606 VSUBS 0.029866f
C1360 VTAIL.n607 VSUBS 0.013379f
C1361 VTAIL.n608 VSUBS 0.012636f
C1362 VTAIL.n609 VSUBS 0.023514f
C1363 VTAIL.n610 VSUBS 0.023514f
C1364 VTAIL.n611 VSUBS 0.012636f
C1365 VTAIL.n612 VSUBS 0.013379f
C1366 VTAIL.n613 VSUBS 0.029866f
C1367 VTAIL.n614 VSUBS 0.029866f
C1368 VTAIL.n615 VSUBS 0.013379f
C1369 VTAIL.n616 VSUBS 0.012636f
C1370 VTAIL.n617 VSUBS 0.023514f
C1371 VTAIL.n618 VSUBS 0.023514f
C1372 VTAIL.n619 VSUBS 0.012636f
C1373 VTAIL.n620 VSUBS 0.013379f
C1374 VTAIL.n621 VSUBS 0.029866f
C1375 VTAIL.n622 VSUBS 0.029866f
C1376 VTAIL.n623 VSUBS 0.013379f
C1377 VTAIL.n624 VSUBS 0.012636f
C1378 VTAIL.n625 VSUBS 0.023514f
C1379 VTAIL.n626 VSUBS 0.023514f
C1380 VTAIL.n627 VSUBS 0.012636f
C1381 VTAIL.n628 VSUBS 0.013379f
C1382 VTAIL.n629 VSUBS 0.029866f
C1383 VTAIL.n630 VSUBS 0.029866f
C1384 VTAIL.n631 VSUBS 0.013379f
C1385 VTAIL.n632 VSUBS 0.012636f
C1386 VTAIL.n633 VSUBS 0.023514f
C1387 VTAIL.n634 VSUBS 0.023514f
C1388 VTAIL.n635 VSUBS 0.012636f
C1389 VTAIL.n636 VSUBS 0.013379f
C1390 VTAIL.n637 VSUBS 0.029866f
C1391 VTAIL.n638 VSUBS 0.029866f
C1392 VTAIL.n639 VSUBS 0.013379f
C1393 VTAIL.n640 VSUBS 0.012636f
C1394 VTAIL.n641 VSUBS 0.023514f
C1395 VTAIL.n642 VSUBS 0.023514f
C1396 VTAIL.n643 VSUBS 0.012636f
C1397 VTAIL.n644 VSUBS 0.013379f
C1398 VTAIL.n645 VSUBS 0.029866f
C1399 VTAIL.n646 VSUBS 0.029866f
C1400 VTAIL.n647 VSUBS 0.013379f
C1401 VTAIL.n648 VSUBS 0.012636f
C1402 VTAIL.n649 VSUBS 0.023514f
C1403 VTAIL.n650 VSUBS 0.023514f
C1404 VTAIL.n651 VSUBS 0.012636f
C1405 VTAIL.n652 VSUBS 0.013379f
C1406 VTAIL.n653 VSUBS 0.029866f
C1407 VTAIL.n654 VSUBS 0.072987f
C1408 VTAIL.n655 VSUBS 0.013379f
C1409 VTAIL.n656 VSUBS 0.012636f
C1410 VTAIL.n657 VSUBS 0.052747f
C1411 VTAIL.n658 VSUBS 0.036685f
C1412 VTAIL.n659 VSUBS 0.105071f
C1413 VTAIL.n660 VSUBS 0.026038f
C1414 VTAIL.n661 VSUBS 0.023514f
C1415 VTAIL.n662 VSUBS 0.012636f
C1416 VTAIL.n663 VSUBS 0.029866f
C1417 VTAIL.n664 VSUBS 0.013379f
C1418 VTAIL.n665 VSUBS 0.023514f
C1419 VTAIL.n666 VSUBS 0.012636f
C1420 VTAIL.n667 VSUBS 0.029866f
C1421 VTAIL.n668 VSUBS 0.013379f
C1422 VTAIL.n669 VSUBS 0.023514f
C1423 VTAIL.n670 VSUBS 0.012636f
C1424 VTAIL.n671 VSUBS 0.029866f
C1425 VTAIL.n672 VSUBS 0.013007f
C1426 VTAIL.n673 VSUBS 0.023514f
C1427 VTAIL.n674 VSUBS 0.013007f
C1428 VTAIL.n675 VSUBS 0.012636f
C1429 VTAIL.n676 VSUBS 0.029866f
C1430 VTAIL.n677 VSUBS 0.029866f
C1431 VTAIL.n678 VSUBS 0.013379f
C1432 VTAIL.n679 VSUBS 0.023514f
C1433 VTAIL.n680 VSUBS 0.012636f
C1434 VTAIL.n681 VSUBS 0.029866f
C1435 VTAIL.n682 VSUBS 0.013379f
C1436 VTAIL.n683 VSUBS 0.023514f
C1437 VTAIL.n684 VSUBS 0.012636f
C1438 VTAIL.n685 VSUBS 0.029866f
C1439 VTAIL.n686 VSUBS 0.013379f
C1440 VTAIL.n687 VSUBS 0.023514f
C1441 VTAIL.n688 VSUBS 0.012636f
C1442 VTAIL.n689 VSUBS 0.029866f
C1443 VTAIL.n690 VSUBS 0.013379f
C1444 VTAIL.n691 VSUBS 0.023514f
C1445 VTAIL.n692 VSUBS 0.012636f
C1446 VTAIL.n693 VSUBS 0.029866f
C1447 VTAIL.n694 VSUBS 0.013379f
C1448 VTAIL.n695 VSUBS 1.9957f
C1449 VTAIL.n696 VSUBS 0.012636f
C1450 VTAIL.t4 VSUBS 0.064208f
C1451 VTAIL.n697 VSUBS 0.19787f
C1452 VTAIL.n698 VSUBS 0.019f
C1453 VTAIL.n699 VSUBS 0.0224f
C1454 VTAIL.n700 VSUBS 0.029866f
C1455 VTAIL.n701 VSUBS 0.013379f
C1456 VTAIL.n702 VSUBS 0.012636f
C1457 VTAIL.n703 VSUBS 0.023514f
C1458 VTAIL.n704 VSUBS 0.023514f
C1459 VTAIL.n705 VSUBS 0.012636f
C1460 VTAIL.n706 VSUBS 0.013379f
C1461 VTAIL.n707 VSUBS 0.029866f
C1462 VTAIL.n708 VSUBS 0.029866f
C1463 VTAIL.n709 VSUBS 0.013379f
C1464 VTAIL.n710 VSUBS 0.012636f
C1465 VTAIL.n711 VSUBS 0.023514f
C1466 VTAIL.n712 VSUBS 0.023514f
C1467 VTAIL.n713 VSUBS 0.012636f
C1468 VTAIL.n714 VSUBS 0.013379f
C1469 VTAIL.n715 VSUBS 0.029866f
C1470 VTAIL.n716 VSUBS 0.029866f
C1471 VTAIL.n717 VSUBS 0.013379f
C1472 VTAIL.n718 VSUBS 0.012636f
C1473 VTAIL.n719 VSUBS 0.023514f
C1474 VTAIL.n720 VSUBS 0.023514f
C1475 VTAIL.n721 VSUBS 0.012636f
C1476 VTAIL.n722 VSUBS 0.013379f
C1477 VTAIL.n723 VSUBS 0.029866f
C1478 VTAIL.n724 VSUBS 0.029866f
C1479 VTAIL.n725 VSUBS 0.013379f
C1480 VTAIL.n726 VSUBS 0.012636f
C1481 VTAIL.n727 VSUBS 0.023514f
C1482 VTAIL.n728 VSUBS 0.023514f
C1483 VTAIL.n729 VSUBS 0.012636f
C1484 VTAIL.n730 VSUBS 0.013379f
C1485 VTAIL.n731 VSUBS 0.029866f
C1486 VTAIL.n732 VSUBS 0.029866f
C1487 VTAIL.n733 VSUBS 0.013379f
C1488 VTAIL.n734 VSUBS 0.012636f
C1489 VTAIL.n735 VSUBS 0.023514f
C1490 VTAIL.n736 VSUBS 0.023514f
C1491 VTAIL.n737 VSUBS 0.012636f
C1492 VTAIL.n738 VSUBS 0.013379f
C1493 VTAIL.n739 VSUBS 0.029866f
C1494 VTAIL.n740 VSUBS 0.029866f
C1495 VTAIL.n741 VSUBS 0.013379f
C1496 VTAIL.n742 VSUBS 0.012636f
C1497 VTAIL.n743 VSUBS 0.023514f
C1498 VTAIL.n744 VSUBS 0.023514f
C1499 VTAIL.n745 VSUBS 0.012636f
C1500 VTAIL.n746 VSUBS 0.013379f
C1501 VTAIL.n747 VSUBS 0.029866f
C1502 VTAIL.n748 VSUBS 0.029866f
C1503 VTAIL.n749 VSUBS 0.013379f
C1504 VTAIL.n750 VSUBS 0.012636f
C1505 VTAIL.n751 VSUBS 0.023514f
C1506 VTAIL.n752 VSUBS 0.023514f
C1507 VTAIL.n753 VSUBS 0.012636f
C1508 VTAIL.n754 VSUBS 0.013379f
C1509 VTAIL.n755 VSUBS 0.029866f
C1510 VTAIL.n756 VSUBS 0.029866f
C1511 VTAIL.n757 VSUBS 0.013379f
C1512 VTAIL.n758 VSUBS 0.012636f
C1513 VTAIL.n759 VSUBS 0.023514f
C1514 VTAIL.n760 VSUBS 0.023514f
C1515 VTAIL.n761 VSUBS 0.012636f
C1516 VTAIL.n762 VSUBS 0.013379f
C1517 VTAIL.n763 VSUBS 0.029866f
C1518 VTAIL.n764 VSUBS 0.072987f
C1519 VTAIL.n765 VSUBS 0.013379f
C1520 VTAIL.n766 VSUBS 0.012636f
C1521 VTAIL.n767 VSUBS 0.052747f
C1522 VTAIL.n768 VSUBS 0.036685f
C1523 VTAIL.n769 VSUBS 1.72138f
C1524 VTAIL.n770 VSUBS 0.026038f
C1525 VTAIL.n771 VSUBS 0.023514f
C1526 VTAIL.n772 VSUBS 0.012636f
C1527 VTAIL.n773 VSUBS 0.029866f
C1528 VTAIL.n774 VSUBS 0.013379f
C1529 VTAIL.n775 VSUBS 0.023514f
C1530 VTAIL.n776 VSUBS 0.012636f
C1531 VTAIL.n777 VSUBS 0.029866f
C1532 VTAIL.n778 VSUBS 0.013379f
C1533 VTAIL.n779 VSUBS 0.023514f
C1534 VTAIL.n780 VSUBS 0.012636f
C1535 VTAIL.n781 VSUBS 0.029866f
C1536 VTAIL.n782 VSUBS 0.013007f
C1537 VTAIL.n783 VSUBS 0.023514f
C1538 VTAIL.n784 VSUBS 0.013379f
C1539 VTAIL.n785 VSUBS 0.029866f
C1540 VTAIL.n786 VSUBS 0.013379f
C1541 VTAIL.n787 VSUBS 0.023514f
C1542 VTAIL.n788 VSUBS 0.012636f
C1543 VTAIL.n789 VSUBS 0.029866f
C1544 VTAIL.n790 VSUBS 0.013379f
C1545 VTAIL.n791 VSUBS 0.023514f
C1546 VTAIL.n792 VSUBS 0.012636f
C1547 VTAIL.n793 VSUBS 0.029866f
C1548 VTAIL.n794 VSUBS 0.013379f
C1549 VTAIL.n795 VSUBS 0.023514f
C1550 VTAIL.n796 VSUBS 0.012636f
C1551 VTAIL.n797 VSUBS 0.029866f
C1552 VTAIL.n798 VSUBS 0.013379f
C1553 VTAIL.n799 VSUBS 0.023514f
C1554 VTAIL.n800 VSUBS 0.012636f
C1555 VTAIL.n801 VSUBS 0.029866f
C1556 VTAIL.n802 VSUBS 0.013379f
C1557 VTAIL.n803 VSUBS 1.9957f
C1558 VTAIL.n804 VSUBS 0.012636f
C1559 VTAIL.t1 VSUBS 0.064208f
C1560 VTAIL.n805 VSUBS 0.19787f
C1561 VTAIL.n806 VSUBS 0.019f
C1562 VTAIL.n807 VSUBS 0.0224f
C1563 VTAIL.n808 VSUBS 0.029866f
C1564 VTAIL.n809 VSUBS 0.013379f
C1565 VTAIL.n810 VSUBS 0.012636f
C1566 VTAIL.n811 VSUBS 0.023514f
C1567 VTAIL.n812 VSUBS 0.023514f
C1568 VTAIL.n813 VSUBS 0.012636f
C1569 VTAIL.n814 VSUBS 0.013379f
C1570 VTAIL.n815 VSUBS 0.029866f
C1571 VTAIL.n816 VSUBS 0.029866f
C1572 VTAIL.n817 VSUBS 0.013379f
C1573 VTAIL.n818 VSUBS 0.012636f
C1574 VTAIL.n819 VSUBS 0.023514f
C1575 VTAIL.n820 VSUBS 0.023514f
C1576 VTAIL.n821 VSUBS 0.012636f
C1577 VTAIL.n822 VSUBS 0.013379f
C1578 VTAIL.n823 VSUBS 0.029866f
C1579 VTAIL.n824 VSUBS 0.029866f
C1580 VTAIL.n825 VSUBS 0.013379f
C1581 VTAIL.n826 VSUBS 0.012636f
C1582 VTAIL.n827 VSUBS 0.023514f
C1583 VTAIL.n828 VSUBS 0.023514f
C1584 VTAIL.n829 VSUBS 0.012636f
C1585 VTAIL.n830 VSUBS 0.013379f
C1586 VTAIL.n831 VSUBS 0.029866f
C1587 VTAIL.n832 VSUBS 0.029866f
C1588 VTAIL.n833 VSUBS 0.013379f
C1589 VTAIL.n834 VSUBS 0.012636f
C1590 VTAIL.n835 VSUBS 0.023514f
C1591 VTAIL.n836 VSUBS 0.023514f
C1592 VTAIL.n837 VSUBS 0.012636f
C1593 VTAIL.n838 VSUBS 0.013379f
C1594 VTAIL.n839 VSUBS 0.029866f
C1595 VTAIL.n840 VSUBS 0.029866f
C1596 VTAIL.n841 VSUBS 0.013379f
C1597 VTAIL.n842 VSUBS 0.012636f
C1598 VTAIL.n843 VSUBS 0.023514f
C1599 VTAIL.n844 VSUBS 0.023514f
C1600 VTAIL.n845 VSUBS 0.012636f
C1601 VTAIL.n846 VSUBS 0.012636f
C1602 VTAIL.n847 VSUBS 0.013379f
C1603 VTAIL.n848 VSUBS 0.029866f
C1604 VTAIL.n849 VSUBS 0.029866f
C1605 VTAIL.n850 VSUBS 0.029866f
C1606 VTAIL.n851 VSUBS 0.013007f
C1607 VTAIL.n852 VSUBS 0.012636f
C1608 VTAIL.n853 VSUBS 0.023514f
C1609 VTAIL.n854 VSUBS 0.023514f
C1610 VTAIL.n855 VSUBS 0.012636f
C1611 VTAIL.n856 VSUBS 0.013379f
C1612 VTAIL.n857 VSUBS 0.029866f
C1613 VTAIL.n858 VSUBS 0.029866f
C1614 VTAIL.n859 VSUBS 0.013379f
C1615 VTAIL.n860 VSUBS 0.012636f
C1616 VTAIL.n861 VSUBS 0.023514f
C1617 VTAIL.n862 VSUBS 0.023514f
C1618 VTAIL.n863 VSUBS 0.012636f
C1619 VTAIL.n864 VSUBS 0.013379f
C1620 VTAIL.n865 VSUBS 0.029866f
C1621 VTAIL.n866 VSUBS 0.029866f
C1622 VTAIL.n867 VSUBS 0.013379f
C1623 VTAIL.n868 VSUBS 0.012636f
C1624 VTAIL.n869 VSUBS 0.023514f
C1625 VTAIL.n870 VSUBS 0.023514f
C1626 VTAIL.n871 VSUBS 0.012636f
C1627 VTAIL.n872 VSUBS 0.013379f
C1628 VTAIL.n873 VSUBS 0.029866f
C1629 VTAIL.n874 VSUBS 0.072987f
C1630 VTAIL.n875 VSUBS 0.013379f
C1631 VTAIL.n876 VSUBS 0.012636f
C1632 VTAIL.n877 VSUBS 0.052747f
C1633 VTAIL.n878 VSUBS 0.036685f
C1634 VTAIL.n879 VSUBS 1.69182f
C1635 VP.t0 VSUBS 1.67009f
C1636 VP.t3 VSUBS 1.67011f
C1637 VP.n0 VSUBS 2.50791f
C1638 VP.n1 VSUBS 5.20418f
C1639 VP.t1 VSUBS 1.65902f
C1640 VP.n2 VSUBS 0.626545f
C1641 VP.t2 VSUBS 1.65902f
C1642 VP.n3 VSUBS 0.626545f
C1643 VP.n4 VSUBS 0.052544f
.ends

