* NGSPICE file created from diff_pair_sample_1573.ext - technology: sky130A

.subckt diff_pair_sample_1573 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0.12045 ps=1.06 w=0.73 l=3.27
X1 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0.12045 ps=1.06 w=0.73 l=3.27
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0 ps=0 w=0.73 l=3.27
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0 ps=0 w=0.73 l=3.27
X4 VDD2.t2 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.12045 pd=1.06 as=0.2847 ps=2.24 w=0.73 l=3.27
X5 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0 ps=0 w=0.73 l=3.27
X6 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0.12045 ps=1.06 w=0.73 l=3.27
X7 VDD2.t0 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.12045 pd=1.06 as=0.2847 ps=2.24 w=0.73 l=3.27
X8 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.12045 pd=1.06 as=0.2847 ps=2.24 w=0.73 l=3.27
X9 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.12045 pd=1.06 as=0.2847 ps=2.24 w=0.73 l=3.27
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0 ps=0 w=0.73 l=3.27
X11 VTAIL.t4 VN.t3 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2847 pd=2.24 as=0.12045 ps=1.06 w=0.73 l=3.27
R0 VN VN.n1 42.5683
R1 VN.n0 VN.t3 40.2384
R2 VN.n1 VN.t2 40.2383
R3 VN.n0 VN.t1 39.1264
R4 VN.n1 VN.t0 39.1264
R5 VN VN.n0 2.5266
R6 VDD2.n2 VDD2.n0 270.039
R7 VDD2.n2 VDD2.n1 236.386
R8 VDD2.n1 VDD2.t1 27.1238
R9 VDD2.n1 VDD2.t0 27.1238
R10 VDD2.n0 VDD2.t3 27.1238
R11 VDD2.n0 VDD2.t2 27.1238
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n7 VTAIL.t6 246.829
R14 VTAIL.n0 VTAIL.t4 246.829
R15 VTAIL.n1 VTAIL.t3 246.829
R16 VTAIL.n2 VTAIL.t2 246.829
R17 VTAIL.n6 VTAIL.t0 246.829
R18 VTAIL.n5 VTAIL.t1 246.829
R19 VTAIL.n4 VTAIL.t5 246.829
R20 VTAIL.n3 VTAIL.t7 246.829
R21 VTAIL.n7 VTAIL.n6 16.0996
R22 VTAIL.n3 VTAIL.n2 16.0996
R23 VTAIL.n4 VTAIL.n3 3.10395
R24 VTAIL.n6 VTAIL.n5 3.10395
R25 VTAIL.n2 VTAIL.n1 3.10395
R26 VTAIL VTAIL.n0 1.61041
R27 VTAIL VTAIL.n7 1.49403
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n462 B.n461 585
R31 B.n141 B.n88 585
R32 B.n140 B.n139 585
R33 B.n138 B.n137 585
R34 B.n136 B.n135 585
R35 B.n134 B.n133 585
R36 B.n132 B.n131 585
R37 B.n130 B.n129 585
R38 B.n128 B.n127 585
R39 B.n126 B.n125 585
R40 B.n124 B.n123 585
R41 B.n122 B.n121 585
R42 B.n120 B.n119 585
R43 B.n118 B.n117 585
R44 B.n116 B.n115 585
R45 B.n114 B.n113 585
R46 B.n112 B.n111 585
R47 B.n110 B.n109 585
R48 B.n108 B.n107 585
R49 B.n106 B.n105 585
R50 B.n104 B.n103 585
R51 B.n102 B.n101 585
R52 B.n100 B.n99 585
R53 B.n98 B.n97 585
R54 B.n96 B.n95 585
R55 B.n74 B.n73 585
R56 B.n460 B.n75 585
R57 B.n465 B.n75 585
R58 B.n459 B.n458 585
R59 B.n458 B.n71 585
R60 B.n457 B.n70 585
R61 B.n471 B.n70 585
R62 B.n456 B.n69 585
R63 B.n472 B.n69 585
R64 B.n455 B.n68 585
R65 B.n473 B.n68 585
R66 B.n454 B.n453 585
R67 B.n453 B.n64 585
R68 B.n452 B.n63 585
R69 B.n479 B.n63 585
R70 B.n451 B.n62 585
R71 B.n480 B.n62 585
R72 B.n450 B.n61 585
R73 B.n481 B.n61 585
R74 B.n449 B.n448 585
R75 B.n448 B.n57 585
R76 B.n447 B.n56 585
R77 B.n487 B.n56 585
R78 B.n446 B.n55 585
R79 B.n488 B.n55 585
R80 B.n445 B.n54 585
R81 B.n489 B.n54 585
R82 B.n444 B.n443 585
R83 B.n443 B.n50 585
R84 B.n442 B.n49 585
R85 B.n495 B.n49 585
R86 B.n441 B.n48 585
R87 B.n496 B.n48 585
R88 B.n440 B.n47 585
R89 B.n497 B.n47 585
R90 B.n439 B.n438 585
R91 B.n438 B.n43 585
R92 B.n437 B.n42 585
R93 B.n503 B.n42 585
R94 B.n436 B.n41 585
R95 B.n504 B.n41 585
R96 B.n435 B.n40 585
R97 B.n505 B.n40 585
R98 B.n434 B.n433 585
R99 B.n433 B.n36 585
R100 B.n432 B.n35 585
R101 B.n511 B.n35 585
R102 B.n431 B.n34 585
R103 B.n512 B.n34 585
R104 B.n430 B.n33 585
R105 B.n513 B.n33 585
R106 B.n429 B.n428 585
R107 B.n428 B.n29 585
R108 B.n427 B.n28 585
R109 B.n519 B.n28 585
R110 B.n426 B.n27 585
R111 B.n520 B.n27 585
R112 B.n425 B.n26 585
R113 B.n521 B.n26 585
R114 B.n424 B.n423 585
R115 B.n423 B.n22 585
R116 B.n422 B.n21 585
R117 B.n527 B.n21 585
R118 B.n421 B.n20 585
R119 B.n528 B.n20 585
R120 B.n420 B.n19 585
R121 B.n529 B.n19 585
R122 B.n419 B.n418 585
R123 B.n418 B.n18 585
R124 B.n417 B.n14 585
R125 B.n535 B.n14 585
R126 B.n416 B.n13 585
R127 B.n536 B.n13 585
R128 B.n415 B.n12 585
R129 B.n537 B.n12 585
R130 B.n414 B.n413 585
R131 B.n413 B.n8 585
R132 B.n412 B.n7 585
R133 B.n543 B.n7 585
R134 B.n411 B.n6 585
R135 B.n544 B.n6 585
R136 B.n410 B.n5 585
R137 B.n545 B.n5 585
R138 B.n409 B.n408 585
R139 B.n408 B.n4 585
R140 B.n407 B.n142 585
R141 B.n407 B.n406 585
R142 B.n397 B.n143 585
R143 B.n144 B.n143 585
R144 B.n399 B.n398 585
R145 B.n400 B.n399 585
R146 B.n396 B.n149 585
R147 B.n149 B.n148 585
R148 B.n395 B.n394 585
R149 B.n394 B.n393 585
R150 B.n151 B.n150 585
R151 B.n386 B.n151 585
R152 B.n385 B.n384 585
R153 B.n387 B.n385 585
R154 B.n383 B.n156 585
R155 B.n156 B.n155 585
R156 B.n382 B.n381 585
R157 B.n381 B.n380 585
R158 B.n158 B.n157 585
R159 B.n159 B.n158 585
R160 B.n373 B.n372 585
R161 B.n374 B.n373 585
R162 B.n371 B.n164 585
R163 B.n164 B.n163 585
R164 B.n370 B.n369 585
R165 B.n369 B.n368 585
R166 B.n166 B.n165 585
R167 B.n167 B.n166 585
R168 B.n361 B.n360 585
R169 B.n362 B.n361 585
R170 B.n359 B.n172 585
R171 B.n172 B.n171 585
R172 B.n358 B.n357 585
R173 B.n357 B.n356 585
R174 B.n174 B.n173 585
R175 B.n175 B.n174 585
R176 B.n349 B.n348 585
R177 B.n350 B.n349 585
R178 B.n347 B.n180 585
R179 B.n180 B.n179 585
R180 B.n346 B.n345 585
R181 B.n345 B.n344 585
R182 B.n182 B.n181 585
R183 B.n183 B.n182 585
R184 B.n337 B.n336 585
R185 B.n338 B.n337 585
R186 B.n335 B.n188 585
R187 B.n188 B.n187 585
R188 B.n334 B.n333 585
R189 B.n333 B.n332 585
R190 B.n190 B.n189 585
R191 B.n191 B.n190 585
R192 B.n325 B.n324 585
R193 B.n326 B.n325 585
R194 B.n323 B.n196 585
R195 B.n196 B.n195 585
R196 B.n322 B.n321 585
R197 B.n321 B.n320 585
R198 B.n198 B.n197 585
R199 B.n199 B.n198 585
R200 B.n313 B.n312 585
R201 B.n314 B.n313 585
R202 B.n311 B.n204 585
R203 B.n204 B.n203 585
R204 B.n310 B.n309 585
R205 B.n309 B.n308 585
R206 B.n206 B.n205 585
R207 B.n207 B.n206 585
R208 B.n301 B.n300 585
R209 B.n302 B.n301 585
R210 B.n299 B.n212 585
R211 B.n212 B.n211 585
R212 B.n298 B.n297 585
R213 B.n297 B.n296 585
R214 B.n214 B.n213 585
R215 B.n215 B.n214 585
R216 B.n289 B.n288 585
R217 B.n290 B.n289 585
R218 B.n218 B.n217 585
R219 B.n237 B.n235 585
R220 B.n238 B.n234 585
R221 B.n238 B.n219 585
R222 B.n241 B.n240 585
R223 B.n242 B.n233 585
R224 B.n244 B.n243 585
R225 B.n246 B.n232 585
R226 B.n249 B.n248 585
R227 B.n251 B.n229 585
R228 B.n253 B.n252 585
R229 B.n255 B.n228 585
R230 B.n258 B.n257 585
R231 B.n259 B.n227 585
R232 B.n261 B.n260 585
R233 B.n263 B.n226 585
R234 B.n266 B.n265 585
R235 B.n267 B.n225 585
R236 B.n272 B.n271 585
R237 B.n274 B.n224 585
R238 B.n277 B.n276 585
R239 B.n278 B.n223 585
R240 B.n280 B.n279 585
R241 B.n282 B.n222 585
R242 B.n283 B.n221 585
R243 B.n286 B.n285 585
R244 B.n287 B.n220 585
R245 B.n220 B.n219 585
R246 B.n292 B.n291 585
R247 B.n291 B.n290 585
R248 B.n293 B.n216 585
R249 B.n216 B.n215 585
R250 B.n295 B.n294 585
R251 B.n296 B.n295 585
R252 B.n210 B.n209 585
R253 B.n211 B.n210 585
R254 B.n304 B.n303 585
R255 B.n303 B.n302 585
R256 B.n305 B.n208 585
R257 B.n208 B.n207 585
R258 B.n307 B.n306 585
R259 B.n308 B.n307 585
R260 B.n202 B.n201 585
R261 B.n203 B.n202 585
R262 B.n316 B.n315 585
R263 B.n315 B.n314 585
R264 B.n317 B.n200 585
R265 B.n200 B.n199 585
R266 B.n319 B.n318 585
R267 B.n320 B.n319 585
R268 B.n194 B.n193 585
R269 B.n195 B.n194 585
R270 B.n328 B.n327 585
R271 B.n327 B.n326 585
R272 B.n329 B.n192 585
R273 B.n192 B.n191 585
R274 B.n331 B.n330 585
R275 B.n332 B.n331 585
R276 B.n186 B.n185 585
R277 B.n187 B.n186 585
R278 B.n340 B.n339 585
R279 B.n339 B.n338 585
R280 B.n341 B.n184 585
R281 B.n184 B.n183 585
R282 B.n343 B.n342 585
R283 B.n344 B.n343 585
R284 B.n178 B.n177 585
R285 B.n179 B.n178 585
R286 B.n352 B.n351 585
R287 B.n351 B.n350 585
R288 B.n353 B.n176 585
R289 B.n176 B.n175 585
R290 B.n355 B.n354 585
R291 B.n356 B.n355 585
R292 B.n170 B.n169 585
R293 B.n171 B.n170 585
R294 B.n364 B.n363 585
R295 B.n363 B.n362 585
R296 B.n365 B.n168 585
R297 B.n168 B.n167 585
R298 B.n367 B.n366 585
R299 B.n368 B.n367 585
R300 B.n162 B.n161 585
R301 B.n163 B.n162 585
R302 B.n376 B.n375 585
R303 B.n375 B.n374 585
R304 B.n377 B.n160 585
R305 B.n160 B.n159 585
R306 B.n379 B.n378 585
R307 B.n380 B.n379 585
R308 B.n154 B.n153 585
R309 B.n155 B.n154 585
R310 B.n389 B.n388 585
R311 B.n388 B.n387 585
R312 B.n390 B.n152 585
R313 B.n386 B.n152 585
R314 B.n392 B.n391 585
R315 B.n393 B.n392 585
R316 B.n147 B.n146 585
R317 B.n148 B.n147 585
R318 B.n402 B.n401 585
R319 B.n401 B.n400 585
R320 B.n403 B.n145 585
R321 B.n145 B.n144 585
R322 B.n405 B.n404 585
R323 B.n406 B.n405 585
R324 B.n2 B.n0 585
R325 B.n4 B.n2 585
R326 B.n3 B.n1 585
R327 B.n544 B.n3 585
R328 B.n542 B.n541 585
R329 B.n543 B.n542 585
R330 B.n540 B.n9 585
R331 B.n9 B.n8 585
R332 B.n539 B.n538 585
R333 B.n538 B.n537 585
R334 B.n11 B.n10 585
R335 B.n536 B.n11 585
R336 B.n534 B.n533 585
R337 B.n535 B.n534 585
R338 B.n532 B.n15 585
R339 B.n18 B.n15 585
R340 B.n531 B.n530 585
R341 B.n530 B.n529 585
R342 B.n17 B.n16 585
R343 B.n528 B.n17 585
R344 B.n526 B.n525 585
R345 B.n527 B.n526 585
R346 B.n524 B.n23 585
R347 B.n23 B.n22 585
R348 B.n523 B.n522 585
R349 B.n522 B.n521 585
R350 B.n25 B.n24 585
R351 B.n520 B.n25 585
R352 B.n518 B.n517 585
R353 B.n519 B.n518 585
R354 B.n516 B.n30 585
R355 B.n30 B.n29 585
R356 B.n515 B.n514 585
R357 B.n514 B.n513 585
R358 B.n32 B.n31 585
R359 B.n512 B.n32 585
R360 B.n510 B.n509 585
R361 B.n511 B.n510 585
R362 B.n508 B.n37 585
R363 B.n37 B.n36 585
R364 B.n507 B.n506 585
R365 B.n506 B.n505 585
R366 B.n39 B.n38 585
R367 B.n504 B.n39 585
R368 B.n502 B.n501 585
R369 B.n503 B.n502 585
R370 B.n500 B.n44 585
R371 B.n44 B.n43 585
R372 B.n499 B.n498 585
R373 B.n498 B.n497 585
R374 B.n46 B.n45 585
R375 B.n496 B.n46 585
R376 B.n494 B.n493 585
R377 B.n495 B.n494 585
R378 B.n492 B.n51 585
R379 B.n51 B.n50 585
R380 B.n491 B.n490 585
R381 B.n490 B.n489 585
R382 B.n53 B.n52 585
R383 B.n488 B.n53 585
R384 B.n486 B.n485 585
R385 B.n487 B.n486 585
R386 B.n484 B.n58 585
R387 B.n58 B.n57 585
R388 B.n483 B.n482 585
R389 B.n482 B.n481 585
R390 B.n60 B.n59 585
R391 B.n480 B.n60 585
R392 B.n478 B.n477 585
R393 B.n479 B.n478 585
R394 B.n476 B.n65 585
R395 B.n65 B.n64 585
R396 B.n475 B.n474 585
R397 B.n474 B.n473 585
R398 B.n67 B.n66 585
R399 B.n472 B.n67 585
R400 B.n470 B.n469 585
R401 B.n471 B.n470 585
R402 B.n468 B.n72 585
R403 B.n72 B.n71 585
R404 B.n467 B.n466 585
R405 B.n466 B.n465 585
R406 B.n547 B.n546 585
R407 B.n546 B.n545 585
R408 B.n291 B.n218 521.33
R409 B.n466 B.n74 521.33
R410 B.n289 B.n220 521.33
R411 B.n462 B.n75 521.33
R412 B.n268 B.t17 305.796
R413 B.n230 B.t14 305.796
R414 B.n92 B.t9 305.796
R415 B.n89 B.t6 305.796
R416 B.n464 B.n463 256.663
R417 B.n464 B.n87 256.663
R418 B.n464 B.n86 256.663
R419 B.n464 B.n85 256.663
R420 B.n464 B.n84 256.663
R421 B.n464 B.n83 256.663
R422 B.n464 B.n82 256.663
R423 B.n464 B.n81 256.663
R424 B.n464 B.n80 256.663
R425 B.n464 B.n79 256.663
R426 B.n464 B.n78 256.663
R427 B.n464 B.n77 256.663
R428 B.n464 B.n76 256.663
R429 B.n236 B.n219 256.663
R430 B.n239 B.n219 256.663
R431 B.n245 B.n219 256.663
R432 B.n247 B.n219 256.663
R433 B.n254 B.n219 256.663
R434 B.n256 B.n219 256.663
R435 B.n262 B.n219 256.663
R436 B.n264 B.n219 256.663
R437 B.n273 B.n219 256.663
R438 B.n275 B.n219 256.663
R439 B.n281 B.n219 256.663
R440 B.n284 B.n219 256.663
R441 B.n269 B.t16 235.978
R442 B.n231 B.t13 235.978
R443 B.n93 B.t10 235.978
R444 B.n90 B.t7 235.978
R445 B.n290 B.n219 210.659
R446 B.n465 B.n464 210.659
R447 B.n268 B.t15 209.81
R448 B.n230 B.t11 209.81
R449 B.n92 B.t8 209.81
R450 B.n89 B.t4 209.81
R451 B.n291 B.n216 163.367
R452 B.n295 B.n216 163.367
R453 B.n295 B.n210 163.367
R454 B.n303 B.n210 163.367
R455 B.n303 B.n208 163.367
R456 B.n307 B.n208 163.367
R457 B.n307 B.n202 163.367
R458 B.n315 B.n202 163.367
R459 B.n315 B.n200 163.367
R460 B.n319 B.n200 163.367
R461 B.n319 B.n194 163.367
R462 B.n327 B.n194 163.367
R463 B.n327 B.n192 163.367
R464 B.n331 B.n192 163.367
R465 B.n331 B.n186 163.367
R466 B.n339 B.n186 163.367
R467 B.n339 B.n184 163.367
R468 B.n343 B.n184 163.367
R469 B.n343 B.n178 163.367
R470 B.n351 B.n178 163.367
R471 B.n351 B.n176 163.367
R472 B.n355 B.n176 163.367
R473 B.n355 B.n170 163.367
R474 B.n363 B.n170 163.367
R475 B.n363 B.n168 163.367
R476 B.n367 B.n168 163.367
R477 B.n367 B.n162 163.367
R478 B.n375 B.n162 163.367
R479 B.n375 B.n160 163.367
R480 B.n379 B.n160 163.367
R481 B.n379 B.n154 163.367
R482 B.n388 B.n154 163.367
R483 B.n388 B.n152 163.367
R484 B.n392 B.n152 163.367
R485 B.n392 B.n147 163.367
R486 B.n401 B.n147 163.367
R487 B.n401 B.n145 163.367
R488 B.n405 B.n145 163.367
R489 B.n405 B.n2 163.367
R490 B.n546 B.n2 163.367
R491 B.n546 B.n3 163.367
R492 B.n542 B.n3 163.367
R493 B.n542 B.n9 163.367
R494 B.n538 B.n9 163.367
R495 B.n538 B.n11 163.367
R496 B.n534 B.n11 163.367
R497 B.n534 B.n15 163.367
R498 B.n530 B.n15 163.367
R499 B.n530 B.n17 163.367
R500 B.n526 B.n17 163.367
R501 B.n526 B.n23 163.367
R502 B.n522 B.n23 163.367
R503 B.n522 B.n25 163.367
R504 B.n518 B.n25 163.367
R505 B.n518 B.n30 163.367
R506 B.n514 B.n30 163.367
R507 B.n514 B.n32 163.367
R508 B.n510 B.n32 163.367
R509 B.n510 B.n37 163.367
R510 B.n506 B.n37 163.367
R511 B.n506 B.n39 163.367
R512 B.n502 B.n39 163.367
R513 B.n502 B.n44 163.367
R514 B.n498 B.n44 163.367
R515 B.n498 B.n46 163.367
R516 B.n494 B.n46 163.367
R517 B.n494 B.n51 163.367
R518 B.n490 B.n51 163.367
R519 B.n490 B.n53 163.367
R520 B.n486 B.n53 163.367
R521 B.n486 B.n58 163.367
R522 B.n482 B.n58 163.367
R523 B.n482 B.n60 163.367
R524 B.n478 B.n60 163.367
R525 B.n478 B.n65 163.367
R526 B.n474 B.n65 163.367
R527 B.n474 B.n67 163.367
R528 B.n470 B.n67 163.367
R529 B.n470 B.n72 163.367
R530 B.n466 B.n72 163.367
R531 B.n238 B.n237 163.367
R532 B.n240 B.n238 163.367
R533 B.n244 B.n233 163.367
R534 B.n248 B.n246 163.367
R535 B.n253 B.n229 163.367
R536 B.n257 B.n255 163.367
R537 B.n261 B.n227 163.367
R538 B.n265 B.n263 163.367
R539 B.n272 B.n225 163.367
R540 B.n276 B.n274 163.367
R541 B.n280 B.n223 163.367
R542 B.n283 B.n282 163.367
R543 B.n285 B.n220 163.367
R544 B.n289 B.n214 163.367
R545 B.n297 B.n214 163.367
R546 B.n297 B.n212 163.367
R547 B.n301 B.n212 163.367
R548 B.n301 B.n206 163.367
R549 B.n309 B.n206 163.367
R550 B.n309 B.n204 163.367
R551 B.n313 B.n204 163.367
R552 B.n313 B.n198 163.367
R553 B.n321 B.n198 163.367
R554 B.n321 B.n196 163.367
R555 B.n325 B.n196 163.367
R556 B.n325 B.n190 163.367
R557 B.n333 B.n190 163.367
R558 B.n333 B.n188 163.367
R559 B.n337 B.n188 163.367
R560 B.n337 B.n182 163.367
R561 B.n345 B.n182 163.367
R562 B.n345 B.n180 163.367
R563 B.n349 B.n180 163.367
R564 B.n349 B.n174 163.367
R565 B.n357 B.n174 163.367
R566 B.n357 B.n172 163.367
R567 B.n361 B.n172 163.367
R568 B.n361 B.n166 163.367
R569 B.n369 B.n166 163.367
R570 B.n369 B.n164 163.367
R571 B.n373 B.n164 163.367
R572 B.n373 B.n158 163.367
R573 B.n381 B.n158 163.367
R574 B.n381 B.n156 163.367
R575 B.n385 B.n156 163.367
R576 B.n385 B.n151 163.367
R577 B.n394 B.n151 163.367
R578 B.n394 B.n149 163.367
R579 B.n399 B.n149 163.367
R580 B.n399 B.n143 163.367
R581 B.n407 B.n143 163.367
R582 B.n408 B.n407 163.367
R583 B.n408 B.n5 163.367
R584 B.n6 B.n5 163.367
R585 B.n7 B.n6 163.367
R586 B.n413 B.n7 163.367
R587 B.n413 B.n12 163.367
R588 B.n13 B.n12 163.367
R589 B.n14 B.n13 163.367
R590 B.n418 B.n14 163.367
R591 B.n418 B.n19 163.367
R592 B.n20 B.n19 163.367
R593 B.n21 B.n20 163.367
R594 B.n423 B.n21 163.367
R595 B.n423 B.n26 163.367
R596 B.n27 B.n26 163.367
R597 B.n28 B.n27 163.367
R598 B.n428 B.n28 163.367
R599 B.n428 B.n33 163.367
R600 B.n34 B.n33 163.367
R601 B.n35 B.n34 163.367
R602 B.n433 B.n35 163.367
R603 B.n433 B.n40 163.367
R604 B.n41 B.n40 163.367
R605 B.n42 B.n41 163.367
R606 B.n438 B.n42 163.367
R607 B.n438 B.n47 163.367
R608 B.n48 B.n47 163.367
R609 B.n49 B.n48 163.367
R610 B.n443 B.n49 163.367
R611 B.n443 B.n54 163.367
R612 B.n55 B.n54 163.367
R613 B.n56 B.n55 163.367
R614 B.n448 B.n56 163.367
R615 B.n448 B.n61 163.367
R616 B.n62 B.n61 163.367
R617 B.n63 B.n62 163.367
R618 B.n453 B.n63 163.367
R619 B.n453 B.n68 163.367
R620 B.n69 B.n68 163.367
R621 B.n70 B.n69 163.367
R622 B.n458 B.n70 163.367
R623 B.n458 B.n75 163.367
R624 B.n97 B.n96 163.367
R625 B.n101 B.n100 163.367
R626 B.n105 B.n104 163.367
R627 B.n109 B.n108 163.367
R628 B.n113 B.n112 163.367
R629 B.n117 B.n116 163.367
R630 B.n121 B.n120 163.367
R631 B.n125 B.n124 163.367
R632 B.n129 B.n128 163.367
R633 B.n133 B.n132 163.367
R634 B.n137 B.n136 163.367
R635 B.n139 B.n88 163.367
R636 B.n290 B.n215 124.564
R637 B.n296 B.n215 124.564
R638 B.n296 B.n211 124.564
R639 B.n302 B.n211 124.564
R640 B.n302 B.n207 124.564
R641 B.n308 B.n207 124.564
R642 B.n308 B.n203 124.564
R643 B.n314 B.n203 124.564
R644 B.n320 B.n199 124.564
R645 B.n320 B.n195 124.564
R646 B.n326 B.n195 124.564
R647 B.n326 B.n191 124.564
R648 B.n332 B.n191 124.564
R649 B.n332 B.n187 124.564
R650 B.n338 B.n187 124.564
R651 B.n338 B.n183 124.564
R652 B.n344 B.n183 124.564
R653 B.n344 B.n179 124.564
R654 B.n350 B.n179 124.564
R655 B.n350 B.n175 124.564
R656 B.n356 B.n175 124.564
R657 B.n362 B.n171 124.564
R658 B.n362 B.n167 124.564
R659 B.n368 B.n167 124.564
R660 B.n368 B.n163 124.564
R661 B.n374 B.n163 124.564
R662 B.n374 B.n159 124.564
R663 B.n380 B.n159 124.564
R664 B.n380 B.n155 124.564
R665 B.n387 B.n155 124.564
R666 B.n387 B.n386 124.564
R667 B.n393 B.n148 124.564
R668 B.n400 B.n148 124.564
R669 B.n400 B.n144 124.564
R670 B.n406 B.n144 124.564
R671 B.n406 B.n4 124.564
R672 B.n545 B.n4 124.564
R673 B.n545 B.n544 124.564
R674 B.n544 B.n543 124.564
R675 B.n543 B.n8 124.564
R676 B.n537 B.n8 124.564
R677 B.n537 B.n536 124.564
R678 B.n536 B.n535 124.564
R679 B.n529 B.n18 124.564
R680 B.n529 B.n528 124.564
R681 B.n528 B.n527 124.564
R682 B.n527 B.n22 124.564
R683 B.n521 B.n22 124.564
R684 B.n521 B.n520 124.564
R685 B.n520 B.n519 124.564
R686 B.n519 B.n29 124.564
R687 B.n513 B.n29 124.564
R688 B.n513 B.n512 124.564
R689 B.n511 B.n36 124.564
R690 B.n505 B.n36 124.564
R691 B.n505 B.n504 124.564
R692 B.n504 B.n503 124.564
R693 B.n503 B.n43 124.564
R694 B.n497 B.n43 124.564
R695 B.n497 B.n496 124.564
R696 B.n496 B.n495 124.564
R697 B.n495 B.n50 124.564
R698 B.n489 B.n50 124.564
R699 B.n489 B.n488 124.564
R700 B.n488 B.n487 124.564
R701 B.n487 B.n57 124.564
R702 B.n481 B.n480 124.564
R703 B.n480 B.n479 124.564
R704 B.n479 B.n64 124.564
R705 B.n473 B.n64 124.564
R706 B.n473 B.n472 124.564
R707 B.n472 B.n471 124.564
R708 B.n471 B.n71 124.564
R709 B.n465 B.n71 124.564
R710 B.n393 B.t3 111.74
R711 B.n535 B.t1 111.74
R712 B.n314 B.t12 89.759
R713 B.n481 B.t5 89.759
R714 B.n236 B.n218 71.676
R715 B.n240 B.n239 71.676
R716 B.n245 B.n244 71.676
R717 B.n248 B.n247 71.676
R718 B.n254 B.n253 71.676
R719 B.n257 B.n256 71.676
R720 B.n262 B.n261 71.676
R721 B.n265 B.n264 71.676
R722 B.n273 B.n272 71.676
R723 B.n276 B.n275 71.676
R724 B.n281 B.n280 71.676
R725 B.n284 B.n283 71.676
R726 B.n76 B.n74 71.676
R727 B.n97 B.n77 71.676
R728 B.n101 B.n78 71.676
R729 B.n105 B.n79 71.676
R730 B.n109 B.n80 71.676
R731 B.n113 B.n81 71.676
R732 B.n117 B.n82 71.676
R733 B.n121 B.n83 71.676
R734 B.n125 B.n84 71.676
R735 B.n129 B.n85 71.676
R736 B.n133 B.n86 71.676
R737 B.n137 B.n87 71.676
R738 B.n463 B.n88 71.676
R739 B.n463 B.n462 71.676
R740 B.n139 B.n87 71.676
R741 B.n136 B.n86 71.676
R742 B.n132 B.n85 71.676
R743 B.n128 B.n84 71.676
R744 B.n124 B.n83 71.676
R745 B.n120 B.n82 71.676
R746 B.n116 B.n81 71.676
R747 B.n112 B.n80 71.676
R748 B.n108 B.n79 71.676
R749 B.n104 B.n78 71.676
R750 B.n100 B.n77 71.676
R751 B.n96 B.n76 71.676
R752 B.n237 B.n236 71.676
R753 B.n239 B.n233 71.676
R754 B.n246 B.n245 71.676
R755 B.n247 B.n229 71.676
R756 B.n255 B.n254 71.676
R757 B.n256 B.n227 71.676
R758 B.n263 B.n262 71.676
R759 B.n264 B.n225 71.676
R760 B.n274 B.n273 71.676
R761 B.n275 B.n223 71.676
R762 B.n282 B.n281 71.676
R763 B.n285 B.n284 71.676
R764 B.n269 B.n268 69.8187
R765 B.n231 B.n230 69.8187
R766 B.n93 B.n92 69.8187
R767 B.n90 B.n89 69.8187
R768 B.n356 B.t2 64.1137
R769 B.t0 B.n511 64.1137
R770 B.t2 B.n171 60.4501
R771 B.n512 B.t0 60.4501
R772 B.n270 B.n269 59.5399
R773 B.n250 B.n231 59.5399
R774 B.n94 B.n93 59.5399
R775 B.n91 B.n90 59.5399
R776 B.t12 B.n199 34.8048
R777 B.t5 B.n57 34.8048
R778 B.n467 B.n73 33.8737
R779 B.n461 B.n460 33.8737
R780 B.n288 B.n287 33.8737
R781 B.n292 B.n217 33.8737
R782 B B.n547 18.0485
R783 B.n386 B.t3 12.8231
R784 B.n18 B.t1 12.8231
R785 B.n95 B.n73 10.6151
R786 B.n98 B.n95 10.6151
R787 B.n99 B.n98 10.6151
R788 B.n102 B.n99 10.6151
R789 B.n103 B.n102 10.6151
R790 B.n106 B.n103 10.6151
R791 B.n107 B.n106 10.6151
R792 B.n111 B.n110 10.6151
R793 B.n114 B.n111 10.6151
R794 B.n115 B.n114 10.6151
R795 B.n118 B.n115 10.6151
R796 B.n119 B.n118 10.6151
R797 B.n122 B.n119 10.6151
R798 B.n123 B.n122 10.6151
R799 B.n126 B.n123 10.6151
R800 B.n127 B.n126 10.6151
R801 B.n131 B.n130 10.6151
R802 B.n134 B.n131 10.6151
R803 B.n135 B.n134 10.6151
R804 B.n138 B.n135 10.6151
R805 B.n140 B.n138 10.6151
R806 B.n141 B.n140 10.6151
R807 B.n461 B.n141 10.6151
R808 B.n288 B.n213 10.6151
R809 B.n298 B.n213 10.6151
R810 B.n299 B.n298 10.6151
R811 B.n300 B.n299 10.6151
R812 B.n300 B.n205 10.6151
R813 B.n310 B.n205 10.6151
R814 B.n311 B.n310 10.6151
R815 B.n312 B.n311 10.6151
R816 B.n312 B.n197 10.6151
R817 B.n322 B.n197 10.6151
R818 B.n323 B.n322 10.6151
R819 B.n324 B.n323 10.6151
R820 B.n324 B.n189 10.6151
R821 B.n334 B.n189 10.6151
R822 B.n335 B.n334 10.6151
R823 B.n336 B.n335 10.6151
R824 B.n336 B.n181 10.6151
R825 B.n346 B.n181 10.6151
R826 B.n347 B.n346 10.6151
R827 B.n348 B.n347 10.6151
R828 B.n348 B.n173 10.6151
R829 B.n358 B.n173 10.6151
R830 B.n359 B.n358 10.6151
R831 B.n360 B.n359 10.6151
R832 B.n360 B.n165 10.6151
R833 B.n370 B.n165 10.6151
R834 B.n371 B.n370 10.6151
R835 B.n372 B.n371 10.6151
R836 B.n372 B.n157 10.6151
R837 B.n382 B.n157 10.6151
R838 B.n383 B.n382 10.6151
R839 B.n384 B.n383 10.6151
R840 B.n384 B.n150 10.6151
R841 B.n395 B.n150 10.6151
R842 B.n396 B.n395 10.6151
R843 B.n398 B.n396 10.6151
R844 B.n398 B.n397 10.6151
R845 B.n397 B.n142 10.6151
R846 B.n409 B.n142 10.6151
R847 B.n410 B.n409 10.6151
R848 B.n411 B.n410 10.6151
R849 B.n412 B.n411 10.6151
R850 B.n414 B.n412 10.6151
R851 B.n415 B.n414 10.6151
R852 B.n416 B.n415 10.6151
R853 B.n417 B.n416 10.6151
R854 B.n419 B.n417 10.6151
R855 B.n420 B.n419 10.6151
R856 B.n421 B.n420 10.6151
R857 B.n422 B.n421 10.6151
R858 B.n424 B.n422 10.6151
R859 B.n425 B.n424 10.6151
R860 B.n426 B.n425 10.6151
R861 B.n427 B.n426 10.6151
R862 B.n429 B.n427 10.6151
R863 B.n430 B.n429 10.6151
R864 B.n431 B.n430 10.6151
R865 B.n432 B.n431 10.6151
R866 B.n434 B.n432 10.6151
R867 B.n435 B.n434 10.6151
R868 B.n436 B.n435 10.6151
R869 B.n437 B.n436 10.6151
R870 B.n439 B.n437 10.6151
R871 B.n440 B.n439 10.6151
R872 B.n441 B.n440 10.6151
R873 B.n442 B.n441 10.6151
R874 B.n444 B.n442 10.6151
R875 B.n445 B.n444 10.6151
R876 B.n446 B.n445 10.6151
R877 B.n447 B.n446 10.6151
R878 B.n449 B.n447 10.6151
R879 B.n450 B.n449 10.6151
R880 B.n451 B.n450 10.6151
R881 B.n452 B.n451 10.6151
R882 B.n454 B.n452 10.6151
R883 B.n455 B.n454 10.6151
R884 B.n456 B.n455 10.6151
R885 B.n457 B.n456 10.6151
R886 B.n459 B.n457 10.6151
R887 B.n460 B.n459 10.6151
R888 B.n235 B.n217 10.6151
R889 B.n235 B.n234 10.6151
R890 B.n241 B.n234 10.6151
R891 B.n242 B.n241 10.6151
R892 B.n243 B.n242 10.6151
R893 B.n243 B.n232 10.6151
R894 B.n249 B.n232 10.6151
R895 B.n252 B.n251 10.6151
R896 B.n252 B.n228 10.6151
R897 B.n258 B.n228 10.6151
R898 B.n259 B.n258 10.6151
R899 B.n260 B.n259 10.6151
R900 B.n260 B.n226 10.6151
R901 B.n266 B.n226 10.6151
R902 B.n267 B.n266 10.6151
R903 B.n271 B.n267 10.6151
R904 B.n277 B.n224 10.6151
R905 B.n278 B.n277 10.6151
R906 B.n279 B.n278 10.6151
R907 B.n279 B.n222 10.6151
R908 B.n222 B.n221 10.6151
R909 B.n286 B.n221 10.6151
R910 B.n287 B.n286 10.6151
R911 B.n293 B.n292 10.6151
R912 B.n294 B.n293 10.6151
R913 B.n294 B.n209 10.6151
R914 B.n304 B.n209 10.6151
R915 B.n305 B.n304 10.6151
R916 B.n306 B.n305 10.6151
R917 B.n306 B.n201 10.6151
R918 B.n316 B.n201 10.6151
R919 B.n317 B.n316 10.6151
R920 B.n318 B.n317 10.6151
R921 B.n318 B.n193 10.6151
R922 B.n328 B.n193 10.6151
R923 B.n329 B.n328 10.6151
R924 B.n330 B.n329 10.6151
R925 B.n330 B.n185 10.6151
R926 B.n340 B.n185 10.6151
R927 B.n341 B.n340 10.6151
R928 B.n342 B.n341 10.6151
R929 B.n342 B.n177 10.6151
R930 B.n352 B.n177 10.6151
R931 B.n353 B.n352 10.6151
R932 B.n354 B.n353 10.6151
R933 B.n354 B.n169 10.6151
R934 B.n364 B.n169 10.6151
R935 B.n365 B.n364 10.6151
R936 B.n366 B.n365 10.6151
R937 B.n366 B.n161 10.6151
R938 B.n376 B.n161 10.6151
R939 B.n377 B.n376 10.6151
R940 B.n378 B.n377 10.6151
R941 B.n378 B.n153 10.6151
R942 B.n389 B.n153 10.6151
R943 B.n390 B.n389 10.6151
R944 B.n391 B.n390 10.6151
R945 B.n391 B.n146 10.6151
R946 B.n402 B.n146 10.6151
R947 B.n403 B.n402 10.6151
R948 B.n404 B.n403 10.6151
R949 B.n404 B.n0 10.6151
R950 B.n541 B.n1 10.6151
R951 B.n541 B.n540 10.6151
R952 B.n540 B.n539 10.6151
R953 B.n539 B.n10 10.6151
R954 B.n533 B.n10 10.6151
R955 B.n533 B.n532 10.6151
R956 B.n532 B.n531 10.6151
R957 B.n531 B.n16 10.6151
R958 B.n525 B.n16 10.6151
R959 B.n525 B.n524 10.6151
R960 B.n524 B.n523 10.6151
R961 B.n523 B.n24 10.6151
R962 B.n517 B.n24 10.6151
R963 B.n517 B.n516 10.6151
R964 B.n516 B.n515 10.6151
R965 B.n515 B.n31 10.6151
R966 B.n509 B.n31 10.6151
R967 B.n509 B.n508 10.6151
R968 B.n508 B.n507 10.6151
R969 B.n507 B.n38 10.6151
R970 B.n501 B.n38 10.6151
R971 B.n501 B.n500 10.6151
R972 B.n500 B.n499 10.6151
R973 B.n499 B.n45 10.6151
R974 B.n493 B.n45 10.6151
R975 B.n493 B.n492 10.6151
R976 B.n492 B.n491 10.6151
R977 B.n491 B.n52 10.6151
R978 B.n485 B.n52 10.6151
R979 B.n485 B.n484 10.6151
R980 B.n484 B.n483 10.6151
R981 B.n483 B.n59 10.6151
R982 B.n477 B.n59 10.6151
R983 B.n477 B.n476 10.6151
R984 B.n476 B.n475 10.6151
R985 B.n475 B.n66 10.6151
R986 B.n469 B.n66 10.6151
R987 B.n469 B.n468 10.6151
R988 B.n468 B.n467 10.6151
R989 B.n107 B.n94 9.36635
R990 B.n130 B.n91 9.36635
R991 B.n250 B.n249 9.36635
R992 B.n270 B.n224 9.36635
R993 B.n547 B.n0 2.81026
R994 B.n547 B.n1 2.81026
R995 B.n110 B.n94 1.24928
R996 B.n127 B.n91 1.24928
R997 B.n251 B.n250 1.24928
R998 B.n271 B.n270 1.24928
R999 VP.n17 VP.n16 161.3
R1000 VP.n15 VP.n1 161.3
R1001 VP.n14 VP.n13 161.3
R1002 VP.n12 VP.n2 161.3
R1003 VP.n11 VP.n10 161.3
R1004 VP.n9 VP.n3 161.3
R1005 VP.n8 VP.n7 161.3
R1006 VP.n6 VP.n4 75.3872
R1007 VP.n18 VP.n0 75.3872
R1008 VP.n6 VP.n5 42.4029
R1009 VP.n10 VP.n2 40.4934
R1010 VP.n14 VP.n2 40.4934
R1011 VP.n5 VP.t0 40.2381
R1012 VP.n5 VP.t3 39.1264
R1013 VP.n9 VP.n8 24.4675
R1014 VP.n10 VP.n9 24.4675
R1015 VP.n15 VP.n14 24.4675
R1016 VP.n16 VP.n15 24.4675
R1017 VP.n8 VP.n4 14.6807
R1018 VP.n16 VP.n0 14.6807
R1019 VP.n4 VP.t1 5.38062
R1020 VP.n0 VP.t2 5.38062
R1021 VP.n7 VP.n6 0.354971
R1022 VP.n18 VP.n17 0.354971
R1023 VP VP.n18 0.26696
R1024 VP.n7 VP.n3 0.189894
R1025 VP.n11 VP.n3 0.189894
R1026 VP.n12 VP.n11 0.189894
R1027 VP.n13 VP.n12 0.189894
R1028 VP.n13 VP.n1 0.189894
R1029 VP.n17 VP.n1 0.189894
R1030 VDD1 VDD1.n1 270.565
R1031 VDD1 VDD1.n0 236.444
R1032 VDD1.n0 VDD1.t3 27.1238
R1033 VDD1.n0 VDD1.t0 27.1238
R1034 VDD1.n1 VDD1.t2 27.1238
R1035 VDD1.n1 VDD1.t1 27.1238
C0 VDD1 VTAIL 3.10069f
C1 VDD2 VTAIL 3.15939f
C2 VDD2 VDD1 1.19135f
C3 VP VTAIL 1.55848f
C4 VDD1 VP 0.908805f
C5 VN VTAIL 1.54438f
C6 VDD1 VN 0.15691f
C7 VDD2 VP 0.446008f
C8 VDD2 VN 0.62268f
C9 VP VN 4.59757f
C10 VDD2 B 3.260145f
C11 VDD1 B 6.14133f
C12 VTAIL B 3.088955f
C13 VN B 10.86335f
C14 VP B 9.300426f
C15 VDD1.t3 B 0.015198f
C16 VDD1.t0 B 0.015198f
C17 VDD1.n0 B 0.037351f
C18 VDD1.t2 B 0.015198f
C19 VDD1.t1 B 0.015198f
C20 VDD1.n1 B 0.146786f
C21 VP.t2 B 0.096407f
C22 VP.n0 B 0.187053f
C23 VP.n1 B 0.026521f
C24 VP.n2 B 0.02144f
C25 VP.n3 B 0.026521f
C26 VP.t1 B 0.096407f
C27 VP.n4 B 0.187053f
C28 VP.t0 B 0.340946f
C29 VP.t3 B 0.331841f
C30 VP.n5 B 1.5424f
C31 VP.n6 B 1.1771f
C32 VP.n7 B 0.042805f
C33 VP.n8 B 0.039668f
C34 VP.n9 B 0.049429f
C35 VP.n10 B 0.052711f
C36 VP.n11 B 0.026521f
C37 VP.n12 B 0.026521f
C38 VP.n13 B 0.026521f
C39 VP.n14 B 0.052711f
C40 VP.n15 B 0.049429f
C41 VP.n16 B 0.039668f
C42 VP.n17 B 0.042805f
C43 VP.n18 B 0.06385f
C44 VTAIL.t4 B 0.072708f
C45 VTAIL.n0 B 0.236377f
C46 VTAIL.t3 B 0.072708f
C47 VTAIL.n1 B 0.372924f
C48 VTAIL.t2 B 0.072708f
C49 VTAIL.n2 B 1.05666f
C50 VTAIL.t7 B 0.072708f
C51 VTAIL.n3 B 1.05666f
C52 VTAIL.t5 B 0.072708f
C53 VTAIL.n4 B 0.372924f
C54 VTAIL.t1 B 0.072708f
C55 VTAIL.n5 B 0.372924f
C56 VTAIL.t0 B 0.072708f
C57 VTAIL.n6 B 1.05666f
C58 VTAIL.t6 B 0.072708f
C59 VTAIL.n7 B 0.909472f
C60 VDD2.t3 B 0.016196f
C61 VDD2.t2 B 0.016196f
C62 VDD2.n0 B 0.147802f
C63 VDD2.t1 B 0.016196f
C64 VDD2.t0 B 0.016196f
C65 VDD2.n1 B 0.039715f
C66 VDD2.n2 B 2.66089f
C67 VN.t1 B 0.329173f
C68 VN.t3 B 0.338206f
C69 VN.n0 B 0.281492f
C70 VN.t0 B 0.329173f
C71 VN.t2 B 0.338206f
C72 VN.n1 B 1.54133f
.ends

