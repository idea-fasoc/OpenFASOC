* NGSPICE file created from diff_pair_sample_0279.ext - technology: sky130A

.subckt diff_pair_sample_0279 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0 ps=0 w=4.8 l=2.21
X1 VDD1.t5 VP.t0 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0.792 ps=5.13 w=4.8 l=2.21
X2 VTAIL.t6 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=0.792 ps=5.13 w=4.8 l=2.21
X3 VDD1.t3 VP.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=1.872 ps=10.38 w=4.8 l=2.21
X4 VDD1.t2 VP.t3 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=1.872 ps=10.38 w=4.8 l=2.21
X5 VTAIL.t7 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=0.792 ps=5.13 w=4.8 l=2.21
X6 VTAIL.t1 VN.t0 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=0.792 ps=5.13 w=4.8 l=2.21
X7 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0.792 ps=5.13 w=4.8 l=2.21
X8 VTAIL.t5 VN.t2 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=0.792 ps=5.13 w=4.8 l=2.21
X9 VDD1.t0 VP.t5 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0.792 ps=5.13 w=4.8 l=2.21
X10 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=1.872 ps=10.38 w=4.8 l=2.21
X11 VDD2.t1 VN.t4 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.792 pd=5.13 as=1.872 ps=10.38 w=4.8 l=2.21
X12 VDD2.t0 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0.792 ps=5.13 w=4.8 l=2.21
X13 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0 ps=0 w=4.8 l=2.21
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0 ps=0 w=4.8 l=2.21
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.872 pd=10.38 as=0 ps=0 w=4.8 l=2.21
R0 B.n469 B.n468 585
R1 B.n471 B.n101 585
R2 B.n474 B.n473 585
R3 B.n475 B.n100 585
R4 B.n477 B.n476 585
R5 B.n479 B.n99 585
R6 B.n482 B.n481 585
R7 B.n483 B.n98 585
R8 B.n485 B.n484 585
R9 B.n487 B.n97 585
R10 B.n490 B.n489 585
R11 B.n491 B.n96 585
R12 B.n493 B.n492 585
R13 B.n495 B.n95 585
R14 B.n498 B.n497 585
R15 B.n499 B.n94 585
R16 B.n501 B.n500 585
R17 B.n503 B.n93 585
R18 B.n505 B.n504 585
R19 B.n507 B.n506 585
R20 B.n510 B.n509 585
R21 B.n511 B.n88 585
R22 B.n513 B.n512 585
R23 B.n515 B.n87 585
R24 B.n518 B.n517 585
R25 B.n519 B.n86 585
R26 B.n521 B.n520 585
R27 B.n523 B.n85 585
R28 B.n526 B.n525 585
R29 B.n527 B.n82 585
R30 B.n530 B.n529 585
R31 B.n532 B.n81 585
R32 B.n535 B.n534 585
R33 B.n536 B.n80 585
R34 B.n538 B.n537 585
R35 B.n540 B.n79 585
R36 B.n543 B.n542 585
R37 B.n544 B.n78 585
R38 B.n546 B.n545 585
R39 B.n548 B.n77 585
R40 B.n551 B.n550 585
R41 B.n552 B.n76 585
R42 B.n554 B.n553 585
R43 B.n556 B.n75 585
R44 B.n559 B.n558 585
R45 B.n560 B.n74 585
R46 B.n562 B.n561 585
R47 B.n564 B.n73 585
R48 B.n567 B.n566 585
R49 B.n568 B.n72 585
R50 B.n467 B.n70 585
R51 B.n571 B.n70 585
R52 B.n466 B.n69 585
R53 B.n572 B.n69 585
R54 B.n465 B.n68 585
R55 B.n573 B.n68 585
R56 B.n464 B.n463 585
R57 B.n463 B.n64 585
R58 B.n462 B.n63 585
R59 B.n579 B.n63 585
R60 B.n461 B.n62 585
R61 B.n580 B.n62 585
R62 B.n460 B.n61 585
R63 B.n581 B.n61 585
R64 B.n459 B.n458 585
R65 B.n458 B.n60 585
R66 B.n457 B.n56 585
R67 B.n587 B.n56 585
R68 B.n456 B.n55 585
R69 B.n588 B.n55 585
R70 B.n455 B.n54 585
R71 B.n589 B.n54 585
R72 B.n454 B.n453 585
R73 B.n453 B.n50 585
R74 B.n452 B.n49 585
R75 B.n595 B.n49 585
R76 B.n451 B.n48 585
R77 B.n596 B.n48 585
R78 B.n450 B.n47 585
R79 B.n597 B.n47 585
R80 B.n449 B.n448 585
R81 B.n448 B.n43 585
R82 B.n447 B.n42 585
R83 B.n603 B.n42 585
R84 B.n446 B.n41 585
R85 B.n604 B.n41 585
R86 B.n445 B.n40 585
R87 B.n605 B.n40 585
R88 B.n444 B.n443 585
R89 B.n443 B.n36 585
R90 B.n442 B.n35 585
R91 B.n611 B.n35 585
R92 B.n441 B.n34 585
R93 B.n612 B.n34 585
R94 B.n440 B.n33 585
R95 B.n613 B.n33 585
R96 B.n439 B.n438 585
R97 B.n438 B.n29 585
R98 B.n437 B.n28 585
R99 B.n619 B.n28 585
R100 B.n436 B.n27 585
R101 B.n620 B.n27 585
R102 B.n435 B.n26 585
R103 B.n621 B.n26 585
R104 B.n434 B.n433 585
R105 B.n433 B.n22 585
R106 B.n432 B.n21 585
R107 B.n627 B.n21 585
R108 B.n431 B.n20 585
R109 B.n628 B.n20 585
R110 B.n430 B.n19 585
R111 B.n629 B.n19 585
R112 B.n429 B.n428 585
R113 B.n428 B.n15 585
R114 B.n427 B.n14 585
R115 B.n635 B.n14 585
R116 B.n426 B.n13 585
R117 B.n636 B.n13 585
R118 B.n425 B.n12 585
R119 B.n637 B.n12 585
R120 B.n424 B.n423 585
R121 B.n423 B.n8 585
R122 B.n422 B.n7 585
R123 B.n643 B.n7 585
R124 B.n421 B.n6 585
R125 B.n644 B.n6 585
R126 B.n420 B.n5 585
R127 B.n645 B.n5 585
R128 B.n419 B.n418 585
R129 B.n418 B.n4 585
R130 B.n417 B.n102 585
R131 B.n417 B.n416 585
R132 B.n407 B.n103 585
R133 B.n104 B.n103 585
R134 B.n409 B.n408 585
R135 B.n410 B.n409 585
R136 B.n406 B.n109 585
R137 B.n109 B.n108 585
R138 B.n405 B.n404 585
R139 B.n404 B.n403 585
R140 B.n111 B.n110 585
R141 B.n112 B.n111 585
R142 B.n396 B.n395 585
R143 B.n397 B.n396 585
R144 B.n394 B.n117 585
R145 B.n117 B.n116 585
R146 B.n393 B.n392 585
R147 B.n392 B.n391 585
R148 B.n119 B.n118 585
R149 B.n120 B.n119 585
R150 B.n384 B.n383 585
R151 B.n385 B.n384 585
R152 B.n382 B.n124 585
R153 B.n128 B.n124 585
R154 B.n381 B.n380 585
R155 B.n380 B.n379 585
R156 B.n126 B.n125 585
R157 B.n127 B.n126 585
R158 B.n372 B.n371 585
R159 B.n373 B.n372 585
R160 B.n370 B.n133 585
R161 B.n133 B.n132 585
R162 B.n369 B.n368 585
R163 B.n368 B.n367 585
R164 B.n135 B.n134 585
R165 B.n136 B.n135 585
R166 B.n360 B.n359 585
R167 B.n361 B.n360 585
R168 B.n358 B.n140 585
R169 B.n144 B.n140 585
R170 B.n357 B.n356 585
R171 B.n356 B.n355 585
R172 B.n142 B.n141 585
R173 B.n143 B.n142 585
R174 B.n348 B.n347 585
R175 B.n349 B.n348 585
R176 B.n346 B.n149 585
R177 B.n149 B.n148 585
R178 B.n345 B.n344 585
R179 B.n344 B.n343 585
R180 B.n151 B.n150 585
R181 B.n152 B.n151 585
R182 B.n336 B.n335 585
R183 B.n337 B.n336 585
R184 B.n334 B.n157 585
R185 B.n157 B.n156 585
R186 B.n333 B.n332 585
R187 B.n332 B.n331 585
R188 B.n159 B.n158 585
R189 B.n324 B.n159 585
R190 B.n323 B.n322 585
R191 B.n325 B.n323 585
R192 B.n321 B.n164 585
R193 B.n164 B.n163 585
R194 B.n320 B.n319 585
R195 B.n319 B.n318 585
R196 B.n166 B.n165 585
R197 B.n167 B.n166 585
R198 B.n311 B.n310 585
R199 B.n312 B.n311 585
R200 B.n309 B.n172 585
R201 B.n172 B.n171 585
R202 B.n308 B.n307 585
R203 B.n307 B.n306 585
R204 B.n303 B.n176 585
R205 B.n302 B.n301 585
R206 B.n299 B.n177 585
R207 B.n299 B.n175 585
R208 B.n298 B.n297 585
R209 B.n296 B.n295 585
R210 B.n294 B.n179 585
R211 B.n292 B.n291 585
R212 B.n290 B.n180 585
R213 B.n289 B.n288 585
R214 B.n286 B.n181 585
R215 B.n284 B.n283 585
R216 B.n282 B.n182 585
R217 B.n281 B.n280 585
R218 B.n278 B.n183 585
R219 B.n276 B.n275 585
R220 B.n274 B.n184 585
R221 B.n273 B.n272 585
R222 B.n270 B.n185 585
R223 B.n268 B.n267 585
R224 B.n266 B.n186 585
R225 B.n264 B.n263 585
R226 B.n261 B.n189 585
R227 B.n259 B.n258 585
R228 B.n257 B.n190 585
R229 B.n256 B.n255 585
R230 B.n253 B.n191 585
R231 B.n251 B.n250 585
R232 B.n249 B.n192 585
R233 B.n248 B.n247 585
R234 B.n245 B.n193 585
R235 B.n243 B.n242 585
R236 B.n241 B.n194 585
R237 B.n240 B.n239 585
R238 B.n237 B.n198 585
R239 B.n235 B.n234 585
R240 B.n233 B.n199 585
R241 B.n232 B.n231 585
R242 B.n229 B.n200 585
R243 B.n227 B.n226 585
R244 B.n225 B.n201 585
R245 B.n224 B.n223 585
R246 B.n221 B.n202 585
R247 B.n219 B.n218 585
R248 B.n217 B.n203 585
R249 B.n216 B.n215 585
R250 B.n213 B.n204 585
R251 B.n211 B.n210 585
R252 B.n209 B.n205 585
R253 B.n208 B.n207 585
R254 B.n174 B.n173 585
R255 B.n175 B.n174 585
R256 B.n305 B.n304 585
R257 B.n306 B.n305 585
R258 B.n170 B.n169 585
R259 B.n171 B.n170 585
R260 B.n314 B.n313 585
R261 B.n313 B.n312 585
R262 B.n315 B.n168 585
R263 B.n168 B.n167 585
R264 B.n317 B.n316 585
R265 B.n318 B.n317 585
R266 B.n162 B.n161 585
R267 B.n163 B.n162 585
R268 B.n327 B.n326 585
R269 B.n326 B.n325 585
R270 B.n328 B.n160 585
R271 B.n324 B.n160 585
R272 B.n330 B.n329 585
R273 B.n331 B.n330 585
R274 B.n155 B.n154 585
R275 B.n156 B.n155 585
R276 B.n339 B.n338 585
R277 B.n338 B.n337 585
R278 B.n340 B.n153 585
R279 B.n153 B.n152 585
R280 B.n342 B.n341 585
R281 B.n343 B.n342 585
R282 B.n147 B.n146 585
R283 B.n148 B.n147 585
R284 B.n351 B.n350 585
R285 B.n350 B.n349 585
R286 B.n352 B.n145 585
R287 B.n145 B.n143 585
R288 B.n354 B.n353 585
R289 B.n355 B.n354 585
R290 B.n139 B.n138 585
R291 B.n144 B.n139 585
R292 B.n363 B.n362 585
R293 B.n362 B.n361 585
R294 B.n364 B.n137 585
R295 B.n137 B.n136 585
R296 B.n366 B.n365 585
R297 B.n367 B.n366 585
R298 B.n131 B.n130 585
R299 B.n132 B.n131 585
R300 B.n375 B.n374 585
R301 B.n374 B.n373 585
R302 B.n376 B.n129 585
R303 B.n129 B.n127 585
R304 B.n378 B.n377 585
R305 B.n379 B.n378 585
R306 B.n123 B.n122 585
R307 B.n128 B.n123 585
R308 B.n387 B.n386 585
R309 B.n386 B.n385 585
R310 B.n388 B.n121 585
R311 B.n121 B.n120 585
R312 B.n390 B.n389 585
R313 B.n391 B.n390 585
R314 B.n115 B.n114 585
R315 B.n116 B.n115 585
R316 B.n399 B.n398 585
R317 B.n398 B.n397 585
R318 B.n400 B.n113 585
R319 B.n113 B.n112 585
R320 B.n402 B.n401 585
R321 B.n403 B.n402 585
R322 B.n107 B.n106 585
R323 B.n108 B.n107 585
R324 B.n412 B.n411 585
R325 B.n411 B.n410 585
R326 B.n413 B.n105 585
R327 B.n105 B.n104 585
R328 B.n415 B.n414 585
R329 B.n416 B.n415 585
R330 B.n2 B.n0 585
R331 B.n4 B.n2 585
R332 B.n3 B.n1 585
R333 B.n644 B.n3 585
R334 B.n642 B.n641 585
R335 B.n643 B.n642 585
R336 B.n640 B.n9 585
R337 B.n9 B.n8 585
R338 B.n639 B.n638 585
R339 B.n638 B.n637 585
R340 B.n11 B.n10 585
R341 B.n636 B.n11 585
R342 B.n634 B.n633 585
R343 B.n635 B.n634 585
R344 B.n632 B.n16 585
R345 B.n16 B.n15 585
R346 B.n631 B.n630 585
R347 B.n630 B.n629 585
R348 B.n18 B.n17 585
R349 B.n628 B.n18 585
R350 B.n626 B.n625 585
R351 B.n627 B.n626 585
R352 B.n624 B.n23 585
R353 B.n23 B.n22 585
R354 B.n623 B.n622 585
R355 B.n622 B.n621 585
R356 B.n25 B.n24 585
R357 B.n620 B.n25 585
R358 B.n618 B.n617 585
R359 B.n619 B.n618 585
R360 B.n616 B.n30 585
R361 B.n30 B.n29 585
R362 B.n615 B.n614 585
R363 B.n614 B.n613 585
R364 B.n32 B.n31 585
R365 B.n612 B.n32 585
R366 B.n610 B.n609 585
R367 B.n611 B.n610 585
R368 B.n608 B.n37 585
R369 B.n37 B.n36 585
R370 B.n607 B.n606 585
R371 B.n606 B.n605 585
R372 B.n39 B.n38 585
R373 B.n604 B.n39 585
R374 B.n602 B.n601 585
R375 B.n603 B.n602 585
R376 B.n600 B.n44 585
R377 B.n44 B.n43 585
R378 B.n599 B.n598 585
R379 B.n598 B.n597 585
R380 B.n46 B.n45 585
R381 B.n596 B.n46 585
R382 B.n594 B.n593 585
R383 B.n595 B.n594 585
R384 B.n592 B.n51 585
R385 B.n51 B.n50 585
R386 B.n591 B.n590 585
R387 B.n590 B.n589 585
R388 B.n53 B.n52 585
R389 B.n588 B.n53 585
R390 B.n586 B.n585 585
R391 B.n587 B.n586 585
R392 B.n584 B.n57 585
R393 B.n60 B.n57 585
R394 B.n583 B.n582 585
R395 B.n582 B.n581 585
R396 B.n59 B.n58 585
R397 B.n580 B.n59 585
R398 B.n578 B.n577 585
R399 B.n579 B.n578 585
R400 B.n576 B.n65 585
R401 B.n65 B.n64 585
R402 B.n575 B.n574 585
R403 B.n574 B.n573 585
R404 B.n67 B.n66 585
R405 B.n572 B.n67 585
R406 B.n570 B.n569 585
R407 B.n571 B.n570 585
R408 B.n647 B.n646 585
R409 B.n646 B.n645 585
R410 B.n305 B.n176 535.745
R411 B.n570 B.n72 535.745
R412 B.n307 B.n174 535.745
R413 B.n469 B.n70 535.745
R414 B.n195 B.t17 259.716
R415 B.n187 B.t6 259.716
R416 B.n83 B.t10 259.716
R417 B.n89 B.t14 259.716
R418 B.n470 B.n71 256.663
R419 B.n472 B.n71 256.663
R420 B.n478 B.n71 256.663
R421 B.n480 B.n71 256.663
R422 B.n486 B.n71 256.663
R423 B.n488 B.n71 256.663
R424 B.n494 B.n71 256.663
R425 B.n496 B.n71 256.663
R426 B.n502 B.n71 256.663
R427 B.n92 B.n71 256.663
R428 B.n508 B.n71 256.663
R429 B.n514 B.n71 256.663
R430 B.n516 B.n71 256.663
R431 B.n522 B.n71 256.663
R432 B.n524 B.n71 256.663
R433 B.n531 B.n71 256.663
R434 B.n533 B.n71 256.663
R435 B.n539 B.n71 256.663
R436 B.n541 B.n71 256.663
R437 B.n547 B.n71 256.663
R438 B.n549 B.n71 256.663
R439 B.n555 B.n71 256.663
R440 B.n557 B.n71 256.663
R441 B.n563 B.n71 256.663
R442 B.n565 B.n71 256.663
R443 B.n300 B.n175 256.663
R444 B.n178 B.n175 256.663
R445 B.n293 B.n175 256.663
R446 B.n287 B.n175 256.663
R447 B.n285 B.n175 256.663
R448 B.n279 B.n175 256.663
R449 B.n277 B.n175 256.663
R450 B.n271 B.n175 256.663
R451 B.n269 B.n175 256.663
R452 B.n262 B.n175 256.663
R453 B.n260 B.n175 256.663
R454 B.n254 B.n175 256.663
R455 B.n252 B.n175 256.663
R456 B.n246 B.n175 256.663
R457 B.n244 B.n175 256.663
R458 B.n238 B.n175 256.663
R459 B.n236 B.n175 256.663
R460 B.n230 B.n175 256.663
R461 B.n228 B.n175 256.663
R462 B.n222 B.n175 256.663
R463 B.n220 B.n175 256.663
R464 B.n214 B.n175 256.663
R465 B.n212 B.n175 256.663
R466 B.n206 B.n175 256.663
R467 B.n305 B.n170 163.367
R468 B.n313 B.n170 163.367
R469 B.n313 B.n168 163.367
R470 B.n317 B.n168 163.367
R471 B.n317 B.n162 163.367
R472 B.n326 B.n162 163.367
R473 B.n326 B.n160 163.367
R474 B.n330 B.n160 163.367
R475 B.n330 B.n155 163.367
R476 B.n338 B.n155 163.367
R477 B.n338 B.n153 163.367
R478 B.n342 B.n153 163.367
R479 B.n342 B.n147 163.367
R480 B.n350 B.n147 163.367
R481 B.n350 B.n145 163.367
R482 B.n354 B.n145 163.367
R483 B.n354 B.n139 163.367
R484 B.n362 B.n139 163.367
R485 B.n362 B.n137 163.367
R486 B.n366 B.n137 163.367
R487 B.n366 B.n131 163.367
R488 B.n374 B.n131 163.367
R489 B.n374 B.n129 163.367
R490 B.n378 B.n129 163.367
R491 B.n378 B.n123 163.367
R492 B.n386 B.n123 163.367
R493 B.n386 B.n121 163.367
R494 B.n390 B.n121 163.367
R495 B.n390 B.n115 163.367
R496 B.n398 B.n115 163.367
R497 B.n398 B.n113 163.367
R498 B.n402 B.n113 163.367
R499 B.n402 B.n107 163.367
R500 B.n411 B.n107 163.367
R501 B.n411 B.n105 163.367
R502 B.n415 B.n105 163.367
R503 B.n415 B.n2 163.367
R504 B.n646 B.n2 163.367
R505 B.n646 B.n3 163.367
R506 B.n642 B.n3 163.367
R507 B.n642 B.n9 163.367
R508 B.n638 B.n9 163.367
R509 B.n638 B.n11 163.367
R510 B.n634 B.n11 163.367
R511 B.n634 B.n16 163.367
R512 B.n630 B.n16 163.367
R513 B.n630 B.n18 163.367
R514 B.n626 B.n18 163.367
R515 B.n626 B.n23 163.367
R516 B.n622 B.n23 163.367
R517 B.n622 B.n25 163.367
R518 B.n618 B.n25 163.367
R519 B.n618 B.n30 163.367
R520 B.n614 B.n30 163.367
R521 B.n614 B.n32 163.367
R522 B.n610 B.n32 163.367
R523 B.n610 B.n37 163.367
R524 B.n606 B.n37 163.367
R525 B.n606 B.n39 163.367
R526 B.n602 B.n39 163.367
R527 B.n602 B.n44 163.367
R528 B.n598 B.n44 163.367
R529 B.n598 B.n46 163.367
R530 B.n594 B.n46 163.367
R531 B.n594 B.n51 163.367
R532 B.n590 B.n51 163.367
R533 B.n590 B.n53 163.367
R534 B.n586 B.n53 163.367
R535 B.n586 B.n57 163.367
R536 B.n582 B.n57 163.367
R537 B.n582 B.n59 163.367
R538 B.n578 B.n59 163.367
R539 B.n578 B.n65 163.367
R540 B.n574 B.n65 163.367
R541 B.n574 B.n67 163.367
R542 B.n570 B.n67 163.367
R543 B.n301 B.n299 163.367
R544 B.n299 B.n298 163.367
R545 B.n295 B.n294 163.367
R546 B.n292 B.n180 163.367
R547 B.n288 B.n286 163.367
R548 B.n284 B.n182 163.367
R549 B.n280 B.n278 163.367
R550 B.n276 B.n184 163.367
R551 B.n272 B.n270 163.367
R552 B.n268 B.n186 163.367
R553 B.n263 B.n261 163.367
R554 B.n259 B.n190 163.367
R555 B.n255 B.n253 163.367
R556 B.n251 B.n192 163.367
R557 B.n247 B.n245 163.367
R558 B.n243 B.n194 163.367
R559 B.n239 B.n237 163.367
R560 B.n235 B.n199 163.367
R561 B.n231 B.n229 163.367
R562 B.n227 B.n201 163.367
R563 B.n223 B.n221 163.367
R564 B.n219 B.n203 163.367
R565 B.n215 B.n213 163.367
R566 B.n211 B.n205 163.367
R567 B.n207 B.n174 163.367
R568 B.n307 B.n172 163.367
R569 B.n311 B.n172 163.367
R570 B.n311 B.n166 163.367
R571 B.n319 B.n166 163.367
R572 B.n319 B.n164 163.367
R573 B.n323 B.n164 163.367
R574 B.n323 B.n159 163.367
R575 B.n332 B.n159 163.367
R576 B.n332 B.n157 163.367
R577 B.n336 B.n157 163.367
R578 B.n336 B.n151 163.367
R579 B.n344 B.n151 163.367
R580 B.n344 B.n149 163.367
R581 B.n348 B.n149 163.367
R582 B.n348 B.n142 163.367
R583 B.n356 B.n142 163.367
R584 B.n356 B.n140 163.367
R585 B.n360 B.n140 163.367
R586 B.n360 B.n135 163.367
R587 B.n368 B.n135 163.367
R588 B.n368 B.n133 163.367
R589 B.n372 B.n133 163.367
R590 B.n372 B.n126 163.367
R591 B.n380 B.n126 163.367
R592 B.n380 B.n124 163.367
R593 B.n384 B.n124 163.367
R594 B.n384 B.n119 163.367
R595 B.n392 B.n119 163.367
R596 B.n392 B.n117 163.367
R597 B.n396 B.n117 163.367
R598 B.n396 B.n111 163.367
R599 B.n404 B.n111 163.367
R600 B.n404 B.n109 163.367
R601 B.n409 B.n109 163.367
R602 B.n409 B.n103 163.367
R603 B.n417 B.n103 163.367
R604 B.n418 B.n417 163.367
R605 B.n418 B.n5 163.367
R606 B.n6 B.n5 163.367
R607 B.n7 B.n6 163.367
R608 B.n423 B.n7 163.367
R609 B.n423 B.n12 163.367
R610 B.n13 B.n12 163.367
R611 B.n14 B.n13 163.367
R612 B.n428 B.n14 163.367
R613 B.n428 B.n19 163.367
R614 B.n20 B.n19 163.367
R615 B.n21 B.n20 163.367
R616 B.n433 B.n21 163.367
R617 B.n433 B.n26 163.367
R618 B.n27 B.n26 163.367
R619 B.n28 B.n27 163.367
R620 B.n438 B.n28 163.367
R621 B.n438 B.n33 163.367
R622 B.n34 B.n33 163.367
R623 B.n35 B.n34 163.367
R624 B.n443 B.n35 163.367
R625 B.n443 B.n40 163.367
R626 B.n41 B.n40 163.367
R627 B.n42 B.n41 163.367
R628 B.n448 B.n42 163.367
R629 B.n448 B.n47 163.367
R630 B.n48 B.n47 163.367
R631 B.n49 B.n48 163.367
R632 B.n453 B.n49 163.367
R633 B.n453 B.n54 163.367
R634 B.n55 B.n54 163.367
R635 B.n56 B.n55 163.367
R636 B.n458 B.n56 163.367
R637 B.n458 B.n61 163.367
R638 B.n62 B.n61 163.367
R639 B.n63 B.n62 163.367
R640 B.n463 B.n63 163.367
R641 B.n463 B.n68 163.367
R642 B.n69 B.n68 163.367
R643 B.n70 B.n69 163.367
R644 B.n566 B.n564 163.367
R645 B.n562 B.n74 163.367
R646 B.n558 B.n556 163.367
R647 B.n554 B.n76 163.367
R648 B.n550 B.n548 163.367
R649 B.n546 B.n78 163.367
R650 B.n542 B.n540 163.367
R651 B.n538 B.n80 163.367
R652 B.n534 B.n532 163.367
R653 B.n530 B.n82 163.367
R654 B.n525 B.n523 163.367
R655 B.n521 B.n86 163.367
R656 B.n517 B.n515 163.367
R657 B.n513 B.n88 163.367
R658 B.n509 B.n507 163.367
R659 B.n504 B.n503 163.367
R660 B.n501 B.n94 163.367
R661 B.n497 B.n495 163.367
R662 B.n493 B.n96 163.367
R663 B.n489 B.n487 163.367
R664 B.n485 B.n98 163.367
R665 B.n481 B.n479 163.367
R666 B.n477 B.n100 163.367
R667 B.n473 B.n471 163.367
R668 B.n306 B.n175 134.293
R669 B.n571 B.n71 134.293
R670 B.n195 B.t19 120.389
R671 B.n89 B.t15 120.389
R672 B.n187 B.t9 120.385
R673 B.n83 B.t12 120.385
R674 B.n306 B.n171 74.2437
R675 B.n312 B.n171 74.2437
R676 B.n312 B.n167 74.2437
R677 B.n318 B.n167 74.2437
R678 B.n318 B.n163 74.2437
R679 B.n325 B.n163 74.2437
R680 B.n325 B.n324 74.2437
R681 B.n331 B.n156 74.2437
R682 B.n337 B.n156 74.2437
R683 B.n337 B.n152 74.2437
R684 B.n343 B.n152 74.2437
R685 B.n343 B.n148 74.2437
R686 B.n349 B.n148 74.2437
R687 B.n349 B.n143 74.2437
R688 B.n355 B.n143 74.2437
R689 B.n355 B.n144 74.2437
R690 B.n361 B.n136 74.2437
R691 B.n367 B.n136 74.2437
R692 B.n367 B.n132 74.2437
R693 B.n373 B.n132 74.2437
R694 B.n373 B.n127 74.2437
R695 B.n379 B.n127 74.2437
R696 B.n379 B.n128 74.2437
R697 B.n385 B.n120 74.2437
R698 B.n391 B.n120 74.2437
R699 B.n391 B.n116 74.2437
R700 B.n397 B.n116 74.2437
R701 B.n397 B.n112 74.2437
R702 B.n403 B.n112 74.2437
R703 B.n410 B.n108 74.2437
R704 B.n410 B.n104 74.2437
R705 B.n416 B.n104 74.2437
R706 B.n416 B.n4 74.2437
R707 B.n645 B.n4 74.2437
R708 B.n645 B.n644 74.2437
R709 B.n644 B.n643 74.2437
R710 B.n643 B.n8 74.2437
R711 B.n637 B.n8 74.2437
R712 B.n637 B.n636 74.2437
R713 B.n635 B.n15 74.2437
R714 B.n629 B.n15 74.2437
R715 B.n629 B.n628 74.2437
R716 B.n628 B.n627 74.2437
R717 B.n627 B.n22 74.2437
R718 B.n621 B.n22 74.2437
R719 B.n620 B.n619 74.2437
R720 B.n619 B.n29 74.2437
R721 B.n613 B.n29 74.2437
R722 B.n613 B.n612 74.2437
R723 B.n612 B.n611 74.2437
R724 B.n611 B.n36 74.2437
R725 B.n605 B.n36 74.2437
R726 B.n604 B.n603 74.2437
R727 B.n603 B.n43 74.2437
R728 B.n597 B.n43 74.2437
R729 B.n597 B.n596 74.2437
R730 B.n596 B.n595 74.2437
R731 B.n595 B.n50 74.2437
R732 B.n589 B.n50 74.2437
R733 B.n589 B.n588 74.2437
R734 B.n588 B.n587 74.2437
R735 B.n581 B.n60 74.2437
R736 B.n581 B.n580 74.2437
R737 B.n580 B.n579 74.2437
R738 B.n579 B.n64 74.2437
R739 B.n573 B.n64 74.2437
R740 B.n573 B.n572 74.2437
R741 B.n572 B.n571 74.2437
R742 B.n300 B.n176 71.676
R743 B.n298 B.n178 71.676
R744 B.n294 B.n293 71.676
R745 B.n287 B.n180 71.676
R746 B.n286 B.n285 71.676
R747 B.n279 B.n182 71.676
R748 B.n278 B.n277 71.676
R749 B.n271 B.n184 71.676
R750 B.n270 B.n269 71.676
R751 B.n262 B.n186 71.676
R752 B.n261 B.n260 71.676
R753 B.n254 B.n190 71.676
R754 B.n253 B.n252 71.676
R755 B.n246 B.n192 71.676
R756 B.n245 B.n244 71.676
R757 B.n238 B.n194 71.676
R758 B.n237 B.n236 71.676
R759 B.n230 B.n199 71.676
R760 B.n229 B.n228 71.676
R761 B.n222 B.n201 71.676
R762 B.n221 B.n220 71.676
R763 B.n214 B.n203 71.676
R764 B.n213 B.n212 71.676
R765 B.n206 B.n205 71.676
R766 B.n565 B.n72 71.676
R767 B.n564 B.n563 71.676
R768 B.n557 B.n74 71.676
R769 B.n556 B.n555 71.676
R770 B.n549 B.n76 71.676
R771 B.n548 B.n547 71.676
R772 B.n541 B.n78 71.676
R773 B.n540 B.n539 71.676
R774 B.n533 B.n80 71.676
R775 B.n532 B.n531 71.676
R776 B.n524 B.n82 71.676
R777 B.n523 B.n522 71.676
R778 B.n516 B.n86 71.676
R779 B.n515 B.n514 71.676
R780 B.n508 B.n88 71.676
R781 B.n507 B.n92 71.676
R782 B.n503 B.n502 71.676
R783 B.n496 B.n94 71.676
R784 B.n495 B.n494 71.676
R785 B.n488 B.n96 71.676
R786 B.n487 B.n486 71.676
R787 B.n480 B.n98 71.676
R788 B.n479 B.n478 71.676
R789 B.n472 B.n100 71.676
R790 B.n471 B.n470 71.676
R791 B.n470 B.n469 71.676
R792 B.n473 B.n472 71.676
R793 B.n478 B.n477 71.676
R794 B.n481 B.n480 71.676
R795 B.n486 B.n485 71.676
R796 B.n489 B.n488 71.676
R797 B.n494 B.n493 71.676
R798 B.n497 B.n496 71.676
R799 B.n502 B.n501 71.676
R800 B.n504 B.n92 71.676
R801 B.n509 B.n508 71.676
R802 B.n514 B.n513 71.676
R803 B.n517 B.n516 71.676
R804 B.n522 B.n521 71.676
R805 B.n525 B.n524 71.676
R806 B.n531 B.n530 71.676
R807 B.n534 B.n533 71.676
R808 B.n539 B.n538 71.676
R809 B.n542 B.n541 71.676
R810 B.n547 B.n546 71.676
R811 B.n550 B.n549 71.676
R812 B.n555 B.n554 71.676
R813 B.n558 B.n557 71.676
R814 B.n563 B.n562 71.676
R815 B.n566 B.n565 71.676
R816 B.n301 B.n300 71.676
R817 B.n295 B.n178 71.676
R818 B.n293 B.n292 71.676
R819 B.n288 B.n287 71.676
R820 B.n285 B.n284 71.676
R821 B.n280 B.n279 71.676
R822 B.n277 B.n276 71.676
R823 B.n272 B.n271 71.676
R824 B.n269 B.n268 71.676
R825 B.n263 B.n262 71.676
R826 B.n260 B.n259 71.676
R827 B.n255 B.n254 71.676
R828 B.n252 B.n251 71.676
R829 B.n247 B.n246 71.676
R830 B.n244 B.n243 71.676
R831 B.n239 B.n238 71.676
R832 B.n236 B.n235 71.676
R833 B.n231 B.n230 71.676
R834 B.n228 B.n227 71.676
R835 B.n223 B.n222 71.676
R836 B.n220 B.n219 71.676
R837 B.n215 B.n214 71.676
R838 B.n212 B.n211 71.676
R839 B.n207 B.n206 71.676
R840 B.n196 B.t18 71.1287
R841 B.n90 B.t16 71.1287
R842 B.n188 B.t8 71.1238
R843 B.n84 B.t13 71.1238
R844 B.n331 B.t7 70.9682
R845 B.n587 B.t11 70.9682
R846 B.n385 B.t5 60.0501
R847 B.n621 B.t2 60.0501
R848 B.n197 B.n196 59.5399
R849 B.n265 B.n188 59.5399
R850 B.n528 B.n84 59.5399
R851 B.n91 B.n90 59.5399
R852 B.n144 B.t0 53.4993
R853 B.t1 B.n604 53.4993
R854 B.n196 B.n195 49.2611
R855 B.n188 B.n187 49.2611
R856 B.n84 B.n83 49.2611
R857 B.n90 B.n89 49.2611
R858 B.n403 B.t3 49.132
R859 B.t4 B.n635 49.132
R860 B.n569 B.n568 34.8103
R861 B.n468 B.n467 34.8103
R862 B.n308 B.n173 34.8103
R863 B.n304 B.n303 34.8103
R864 B.t3 B.n108 25.1122
R865 B.n636 B.t4 25.1122
R866 B.n361 B.t0 20.7449
R867 B.n605 B.t1 20.7449
R868 B B.n647 18.0485
R869 B.n128 B.t5 14.194
R870 B.t2 B.n620 14.194
R871 B.n568 B.n567 10.6151
R872 B.n567 B.n73 10.6151
R873 B.n561 B.n73 10.6151
R874 B.n561 B.n560 10.6151
R875 B.n560 B.n559 10.6151
R876 B.n559 B.n75 10.6151
R877 B.n553 B.n75 10.6151
R878 B.n553 B.n552 10.6151
R879 B.n552 B.n551 10.6151
R880 B.n551 B.n77 10.6151
R881 B.n545 B.n77 10.6151
R882 B.n545 B.n544 10.6151
R883 B.n544 B.n543 10.6151
R884 B.n543 B.n79 10.6151
R885 B.n537 B.n79 10.6151
R886 B.n537 B.n536 10.6151
R887 B.n536 B.n535 10.6151
R888 B.n535 B.n81 10.6151
R889 B.n529 B.n81 10.6151
R890 B.n527 B.n526 10.6151
R891 B.n526 B.n85 10.6151
R892 B.n520 B.n85 10.6151
R893 B.n520 B.n519 10.6151
R894 B.n519 B.n518 10.6151
R895 B.n518 B.n87 10.6151
R896 B.n512 B.n87 10.6151
R897 B.n512 B.n511 10.6151
R898 B.n511 B.n510 10.6151
R899 B.n506 B.n505 10.6151
R900 B.n505 B.n93 10.6151
R901 B.n500 B.n93 10.6151
R902 B.n500 B.n499 10.6151
R903 B.n499 B.n498 10.6151
R904 B.n498 B.n95 10.6151
R905 B.n492 B.n95 10.6151
R906 B.n492 B.n491 10.6151
R907 B.n491 B.n490 10.6151
R908 B.n490 B.n97 10.6151
R909 B.n484 B.n97 10.6151
R910 B.n484 B.n483 10.6151
R911 B.n483 B.n482 10.6151
R912 B.n482 B.n99 10.6151
R913 B.n476 B.n99 10.6151
R914 B.n476 B.n475 10.6151
R915 B.n475 B.n474 10.6151
R916 B.n474 B.n101 10.6151
R917 B.n468 B.n101 10.6151
R918 B.n309 B.n308 10.6151
R919 B.n310 B.n309 10.6151
R920 B.n310 B.n165 10.6151
R921 B.n320 B.n165 10.6151
R922 B.n321 B.n320 10.6151
R923 B.n322 B.n321 10.6151
R924 B.n322 B.n158 10.6151
R925 B.n333 B.n158 10.6151
R926 B.n334 B.n333 10.6151
R927 B.n335 B.n334 10.6151
R928 B.n335 B.n150 10.6151
R929 B.n345 B.n150 10.6151
R930 B.n346 B.n345 10.6151
R931 B.n347 B.n346 10.6151
R932 B.n347 B.n141 10.6151
R933 B.n357 B.n141 10.6151
R934 B.n358 B.n357 10.6151
R935 B.n359 B.n358 10.6151
R936 B.n359 B.n134 10.6151
R937 B.n369 B.n134 10.6151
R938 B.n370 B.n369 10.6151
R939 B.n371 B.n370 10.6151
R940 B.n371 B.n125 10.6151
R941 B.n381 B.n125 10.6151
R942 B.n382 B.n381 10.6151
R943 B.n383 B.n382 10.6151
R944 B.n383 B.n118 10.6151
R945 B.n393 B.n118 10.6151
R946 B.n394 B.n393 10.6151
R947 B.n395 B.n394 10.6151
R948 B.n395 B.n110 10.6151
R949 B.n405 B.n110 10.6151
R950 B.n406 B.n405 10.6151
R951 B.n408 B.n406 10.6151
R952 B.n408 B.n407 10.6151
R953 B.n407 B.n102 10.6151
R954 B.n419 B.n102 10.6151
R955 B.n420 B.n419 10.6151
R956 B.n421 B.n420 10.6151
R957 B.n422 B.n421 10.6151
R958 B.n424 B.n422 10.6151
R959 B.n425 B.n424 10.6151
R960 B.n426 B.n425 10.6151
R961 B.n427 B.n426 10.6151
R962 B.n429 B.n427 10.6151
R963 B.n430 B.n429 10.6151
R964 B.n431 B.n430 10.6151
R965 B.n432 B.n431 10.6151
R966 B.n434 B.n432 10.6151
R967 B.n435 B.n434 10.6151
R968 B.n436 B.n435 10.6151
R969 B.n437 B.n436 10.6151
R970 B.n439 B.n437 10.6151
R971 B.n440 B.n439 10.6151
R972 B.n441 B.n440 10.6151
R973 B.n442 B.n441 10.6151
R974 B.n444 B.n442 10.6151
R975 B.n445 B.n444 10.6151
R976 B.n446 B.n445 10.6151
R977 B.n447 B.n446 10.6151
R978 B.n449 B.n447 10.6151
R979 B.n450 B.n449 10.6151
R980 B.n451 B.n450 10.6151
R981 B.n452 B.n451 10.6151
R982 B.n454 B.n452 10.6151
R983 B.n455 B.n454 10.6151
R984 B.n456 B.n455 10.6151
R985 B.n457 B.n456 10.6151
R986 B.n459 B.n457 10.6151
R987 B.n460 B.n459 10.6151
R988 B.n461 B.n460 10.6151
R989 B.n462 B.n461 10.6151
R990 B.n464 B.n462 10.6151
R991 B.n465 B.n464 10.6151
R992 B.n466 B.n465 10.6151
R993 B.n467 B.n466 10.6151
R994 B.n303 B.n302 10.6151
R995 B.n302 B.n177 10.6151
R996 B.n297 B.n177 10.6151
R997 B.n297 B.n296 10.6151
R998 B.n296 B.n179 10.6151
R999 B.n291 B.n179 10.6151
R1000 B.n291 B.n290 10.6151
R1001 B.n290 B.n289 10.6151
R1002 B.n289 B.n181 10.6151
R1003 B.n283 B.n181 10.6151
R1004 B.n283 B.n282 10.6151
R1005 B.n282 B.n281 10.6151
R1006 B.n281 B.n183 10.6151
R1007 B.n275 B.n183 10.6151
R1008 B.n275 B.n274 10.6151
R1009 B.n274 B.n273 10.6151
R1010 B.n273 B.n185 10.6151
R1011 B.n267 B.n185 10.6151
R1012 B.n267 B.n266 10.6151
R1013 B.n264 B.n189 10.6151
R1014 B.n258 B.n189 10.6151
R1015 B.n258 B.n257 10.6151
R1016 B.n257 B.n256 10.6151
R1017 B.n256 B.n191 10.6151
R1018 B.n250 B.n191 10.6151
R1019 B.n250 B.n249 10.6151
R1020 B.n249 B.n248 10.6151
R1021 B.n248 B.n193 10.6151
R1022 B.n242 B.n241 10.6151
R1023 B.n241 B.n240 10.6151
R1024 B.n240 B.n198 10.6151
R1025 B.n234 B.n198 10.6151
R1026 B.n234 B.n233 10.6151
R1027 B.n233 B.n232 10.6151
R1028 B.n232 B.n200 10.6151
R1029 B.n226 B.n200 10.6151
R1030 B.n226 B.n225 10.6151
R1031 B.n225 B.n224 10.6151
R1032 B.n224 B.n202 10.6151
R1033 B.n218 B.n202 10.6151
R1034 B.n218 B.n217 10.6151
R1035 B.n217 B.n216 10.6151
R1036 B.n216 B.n204 10.6151
R1037 B.n210 B.n204 10.6151
R1038 B.n210 B.n209 10.6151
R1039 B.n209 B.n208 10.6151
R1040 B.n208 B.n173 10.6151
R1041 B.n304 B.n169 10.6151
R1042 B.n314 B.n169 10.6151
R1043 B.n315 B.n314 10.6151
R1044 B.n316 B.n315 10.6151
R1045 B.n316 B.n161 10.6151
R1046 B.n327 B.n161 10.6151
R1047 B.n328 B.n327 10.6151
R1048 B.n329 B.n328 10.6151
R1049 B.n329 B.n154 10.6151
R1050 B.n339 B.n154 10.6151
R1051 B.n340 B.n339 10.6151
R1052 B.n341 B.n340 10.6151
R1053 B.n341 B.n146 10.6151
R1054 B.n351 B.n146 10.6151
R1055 B.n352 B.n351 10.6151
R1056 B.n353 B.n352 10.6151
R1057 B.n353 B.n138 10.6151
R1058 B.n363 B.n138 10.6151
R1059 B.n364 B.n363 10.6151
R1060 B.n365 B.n364 10.6151
R1061 B.n365 B.n130 10.6151
R1062 B.n375 B.n130 10.6151
R1063 B.n376 B.n375 10.6151
R1064 B.n377 B.n376 10.6151
R1065 B.n377 B.n122 10.6151
R1066 B.n387 B.n122 10.6151
R1067 B.n388 B.n387 10.6151
R1068 B.n389 B.n388 10.6151
R1069 B.n389 B.n114 10.6151
R1070 B.n399 B.n114 10.6151
R1071 B.n400 B.n399 10.6151
R1072 B.n401 B.n400 10.6151
R1073 B.n401 B.n106 10.6151
R1074 B.n412 B.n106 10.6151
R1075 B.n413 B.n412 10.6151
R1076 B.n414 B.n413 10.6151
R1077 B.n414 B.n0 10.6151
R1078 B.n641 B.n1 10.6151
R1079 B.n641 B.n640 10.6151
R1080 B.n640 B.n639 10.6151
R1081 B.n639 B.n10 10.6151
R1082 B.n633 B.n10 10.6151
R1083 B.n633 B.n632 10.6151
R1084 B.n632 B.n631 10.6151
R1085 B.n631 B.n17 10.6151
R1086 B.n625 B.n17 10.6151
R1087 B.n625 B.n624 10.6151
R1088 B.n624 B.n623 10.6151
R1089 B.n623 B.n24 10.6151
R1090 B.n617 B.n24 10.6151
R1091 B.n617 B.n616 10.6151
R1092 B.n616 B.n615 10.6151
R1093 B.n615 B.n31 10.6151
R1094 B.n609 B.n31 10.6151
R1095 B.n609 B.n608 10.6151
R1096 B.n608 B.n607 10.6151
R1097 B.n607 B.n38 10.6151
R1098 B.n601 B.n38 10.6151
R1099 B.n601 B.n600 10.6151
R1100 B.n600 B.n599 10.6151
R1101 B.n599 B.n45 10.6151
R1102 B.n593 B.n45 10.6151
R1103 B.n593 B.n592 10.6151
R1104 B.n592 B.n591 10.6151
R1105 B.n591 B.n52 10.6151
R1106 B.n585 B.n52 10.6151
R1107 B.n585 B.n584 10.6151
R1108 B.n584 B.n583 10.6151
R1109 B.n583 B.n58 10.6151
R1110 B.n577 B.n58 10.6151
R1111 B.n577 B.n576 10.6151
R1112 B.n576 B.n575 10.6151
R1113 B.n575 B.n66 10.6151
R1114 B.n569 B.n66 10.6151
R1115 B.n529 B.n528 9.36635
R1116 B.n506 B.n91 9.36635
R1117 B.n266 B.n265 9.36635
R1118 B.n242 B.n197 9.36635
R1119 B.n324 B.t7 3.27593
R1120 B.n60 B.t11 3.27593
R1121 B.n647 B.n0 2.81026
R1122 B.n647 B.n1 2.81026
R1123 B.n528 B.n527 1.24928
R1124 B.n510 B.n91 1.24928
R1125 B.n265 B.n264 1.24928
R1126 B.n197 B.n193 1.24928
R1127 VP.n11 VP.n8 161.3
R1128 VP.n13 VP.n12 161.3
R1129 VP.n14 VP.n7 161.3
R1130 VP.n16 VP.n15 161.3
R1131 VP.n17 VP.n6 161.3
R1132 VP.n36 VP.n0 161.3
R1133 VP.n35 VP.n34 161.3
R1134 VP.n33 VP.n1 161.3
R1135 VP.n32 VP.n31 161.3
R1136 VP.n30 VP.n2 161.3
R1137 VP.n28 VP.n27 161.3
R1138 VP.n26 VP.n3 161.3
R1139 VP.n25 VP.n24 161.3
R1140 VP.n23 VP.n4 161.3
R1141 VP.n22 VP.n21 161.3
R1142 VP.n20 VP.n5 96.645
R1143 VP.n38 VP.n37 96.645
R1144 VP.n19 VP.n18 96.645
R1145 VP.n9 VP.t5 84.9908
R1146 VP.n10 VP.n9 59.4181
R1147 VP.n5 VP.t0 52.3444
R1148 VP.n29 VP.t1 52.3444
R1149 VP.n37 VP.t2 52.3444
R1150 VP.n18 VP.t3 52.3444
R1151 VP.n10 VP.t4 52.3444
R1152 VP.n24 VP.n23 42.5146
R1153 VP.n35 VP.n1 42.5146
R1154 VP.n16 VP.n7 42.5146
R1155 VP.n20 VP.n19 41.6815
R1156 VP.n24 VP.n3 38.6395
R1157 VP.n31 VP.n1 38.6395
R1158 VP.n12 VP.n7 38.6395
R1159 VP.n23 VP.n22 24.5923
R1160 VP.n28 VP.n3 24.5923
R1161 VP.n31 VP.n30 24.5923
R1162 VP.n36 VP.n35 24.5923
R1163 VP.n17 VP.n16 24.5923
R1164 VP.n12 VP.n11 24.5923
R1165 VP.n22 VP.n5 14.2638
R1166 VP.n37 VP.n36 14.2638
R1167 VP.n18 VP.n17 14.2638
R1168 VP.n29 VP.n28 12.2964
R1169 VP.n30 VP.n29 12.2964
R1170 VP.n11 VP.n10 12.2964
R1171 VP.n9 VP.n8 9.51334
R1172 VP.n19 VP.n6 0.278335
R1173 VP.n21 VP.n20 0.278335
R1174 VP.n38 VP.n0 0.278335
R1175 VP.n13 VP.n8 0.189894
R1176 VP.n14 VP.n13 0.189894
R1177 VP.n15 VP.n14 0.189894
R1178 VP.n15 VP.n6 0.189894
R1179 VP.n21 VP.n4 0.189894
R1180 VP.n25 VP.n4 0.189894
R1181 VP.n26 VP.n25 0.189894
R1182 VP.n27 VP.n26 0.189894
R1183 VP.n27 VP.n2 0.189894
R1184 VP.n32 VP.n2 0.189894
R1185 VP.n33 VP.n32 0.189894
R1186 VP.n34 VP.n33 0.189894
R1187 VP.n34 VP.n0 0.189894
R1188 VP VP.n38 0.153485
R1189 VTAIL.n7 VTAIL.t3 54.6859
R1190 VTAIL.n11 VTAIL.t2 54.6859
R1191 VTAIL.n2 VTAIL.t11 54.6859
R1192 VTAIL.n10 VTAIL.t8 54.6859
R1193 VTAIL.n9 VTAIL.n8 50.561
R1194 VTAIL.n6 VTAIL.n5 50.561
R1195 VTAIL.n1 VTAIL.n0 50.5608
R1196 VTAIL.n4 VTAIL.n3 50.5608
R1197 VTAIL.n6 VTAIL.n4 20.8841
R1198 VTAIL.n11 VTAIL.n10 18.6945
R1199 VTAIL.n0 VTAIL.t4 4.1255
R1200 VTAIL.n0 VTAIL.t5 4.1255
R1201 VTAIL.n3 VTAIL.t10 4.1255
R1202 VTAIL.n3 VTAIL.t6 4.1255
R1203 VTAIL.n8 VTAIL.t9 4.1255
R1204 VTAIL.n8 VTAIL.t7 4.1255
R1205 VTAIL.n5 VTAIL.t0 4.1255
R1206 VTAIL.n5 VTAIL.t1 4.1255
R1207 VTAIL.n7 VTAIL.n6 2.19016
R1208 VTAIL.n10 VTAIL.n9 2.19016
R1209 VTAIL.n4 VTAIL.n2 2.19016
R1210 VTAIL VTAIL.n11 1.58455
R1211 VTAIL.n9 VTAIL.n7 1.56516
R1212 VTAIL.n2 VTAIL.n1 1.56516
R1213 VTAIL VTAIL.n1 0.606103
R1214 VDD1 VDD1.t0 73.0652
R1215 VDD1.n1 VDD1.t5 72.9515
R1216 VDD1.n1 VDD1.n0 67.7316
R1217 VDD1.n3 VDD1.n2 67.2397
R1218 VDD1.n3 VDD1.n1 36.6474
R1219 VDD1.n2 VDD1.t1 4.1255
R1220 VDD1.n2 VDD1.t2 4.1255
R1221 VDD1.n0 VDD1.t4 4.1255
R1222 VDD1.n0 VDD1.t3 4.1255
R1223 VDD1 VDD1.n3 0.489724
R1224 VN.n25 VN.n14 161.3
R1225 VN.n24 VN.n23 161.3
R1226 VN.n22 VN.n15 161.3
R1227 VN.n21 VN.n20 161.3
R1228 VN.n19 VN.n16 161.3
R1229 VN.n11 VN.n0 161.3
R1230 VN.n10 VN.n9 161.3
R1231 VN.n8 VN.n1 161.3
R1232 VN.n7 VN.n6 161.3
R1233 VN.n5 VN.n2 161.3
R1234 VN.n13 VN.n12 96.645
R1235 VN.n27 VN.n26 96.645
R1236 VN.n3 VN.t5 84.9908
R1237 VN.n17 VN.t3 84.9908
R1238 VN.n4 VN.n3 59.4181
R1239 VN.n18 VN.n17 59.4181
R1240 VN.n4 VN.t2 52.3444
R1241 VN.n12 VN.t4 52.3444
R1242 VN.n18 VN.t0 52.3444
R1243 VN.n26 VN.t1 52.3444
R1244 VN.n10 VN.n1 42.5146
R1245 VN.n24 VN.n15 42.5146
R1246 VN VN.n27 41.9603
R1247 VN.n6 VN.n1 38.6395
R1248 VN.n20 VN.n15 38.6395
R1249 VN.n6 VN.n5 24.5923
R1250 VN.n11 VN.n10 24.5923
R1251 VN.n20 VN.n19 24.5923
R1252 VN.n25 VN.n24 24.5923
R1253 VN.n12 VN.n11 14.2638
R1254 VN.n26 VN.n25 14.2638
R1255 VN.n5 VN.n4 12.2964
R1256 VN.n19 VN.n18 12.2964
R1257 VN.n17 VN.n16 9.51334
R1258 VN.n3 VN.n2 9.51334
R1259 VN.n27 VN.n14 0.278335
R1260 VN.n13 VN.n0 0.278335
R1261 VN.n23 VN.n14 0.189894
R1262 VN.n23 VN.n22 0.189894
R1263 VN.n22 VN.n21 0.189894
R1264 VN.n21 VN.n16 0.189894
R1265 VN.n7 VN.n2 0.189894
R1266 VN.n8 VN.n7 0.189894
R1267 VN.n9 VN.n8 0.189894
R1268 VN.n9 VN.n0 0.189894
R1269 VN VN.n13 0.153485
R1270 VDD2.n1 VDD2.t0 72.9515
R1271 VDD2.n2 VDD2.t4 71.3647
R1272 VDD2.n1 VDD2.n0 67.7316
R1273 VDD2 VDD2.n3 67.7289
R1274 VDD2.n2 VDD2.n1 34.9696
R1275 VDD2.n3 VDD2.t5 4.1255
R1276 VDD2.n3 VDD2.t2 4.1255
R1277 VDD2.n0 VDD2.t3 4.1255
R1278 VDD2.n0 VDD2.t1 4.1255
R1279 VDD2 VDD2.n2 1.70093
C0 VP VDD2 0.429045f
C1 VTAIL VDD1 4.9196f
C2 VN VDD1 0.154205f
C3 VTAIL VP 3.36652f
C4 VP VN 5.21202f
C5 VTAIL VDD2 4.9693f
C6 VP VDD1 3.10662f
C7 VN VDD2 2.83417f
C8 VTAIL VN 3.35232f
C9 VDD2 VDD1 1.25283f
C10 VDD2 B 4.398416f
C11 VDD1 B 4.695908f
C12 VTAIL B 4.409513f
C13 VN B 11.052189f
C14 VP B 9.694203f
C15 VDD2.t0 B 0.863989f
C16 VDD2.t3 B 0.083542f
C17 VDD2.t1 B 0.083542f
C18 VDD2.n0 B 0.678809f
C19 VDD2.n1 B 2.00962f
C20 VDD2.t4 B 0.856508f
C21 VDD2.n2 B 1.85157f
C22 VDD2.t5 B 0.083542f
C23 VDD2.t2 B 0.083542f
C24 VDD2.n3 B 0.678783f
C25 VN.n0 B 0.03896f
C26 VN.t4 B 0.817539f
C27 VN.n1 B 0.02402f
C28 VN.n2 B 0.251855f
C29 VN.t2 B 0.817539f
C30 VN.t5 B 1.00124f
C31 VN.n3 B 0.385101f
C32 VN.n4 B 0.395895f
C33 VN.n5 B 0.041275f
C34 VN.n6 B 0.058933f
C35 VN.n7 B 0.029552f
C36 VN.n8 B 0.029552f
C37 VN.n9 B 0.029552f
C38 VN.n10 B 0.057767f
C39 VN.n11 B 0.043439f
C40 VN.n12 B 0.409466f
C41 VN.n13 B 0.041634f
C42 VN.n14 B 0.03896f
C43 VN.t1 B 0.817539f
C44 VN.n15 B 0.02402f
C45 VN.n16 B 0.251855f
C46 VN.t0 B 0.817539f
C47 VN.t3 B 1.00124f
C48 VN.n17 B 0.385101f
C49 VN.n18 B 0.395895f
C50 VN.n19 B 0.041275f
C51 VN.n20 B 0.058933f
C52 VN.n21 B 0.029552f
C53 VN.n22 B 0.029552f
C54 VN.n23 B 0.029552f
C55 VN.n24 B 0.057767f
C56 VN.n25 B 0.043439f
C57 VN.n26 B 0.409466f
C58 VN.n27 B 1.25115f
C59 VDD1.t0 B 0.877714f
C60 VDD1.t5 B 0.876996f
C61 VDD1.t4 B 0.084799f
C62 VDD1.t3 B 0.084799f
C63 VDD1.n0 B 0.689028f
C64 VDD1.n1 B 2.13615f
C65 VDD1.t1 B 0.084799f
C66 VDD1.t2 B 0.084799f
C67 VDD1.n2 B 0.686261f
C68 VDD1.n3 B 1.8881f
C69 VTAIL.t4 B 0.106184f
C70 VTAIL.t5 B 0.106184f
C71 VTAIL.n0 B 0.78776f
C72 VTAIL.n1 B 0.451546f
C73 VTAIL.t11 B 1.0041f
C74 VTAIL.n2 B 0.66769f
C75 VTAIL.t10 B 0.106184f
C76 VTAIL.t6 B 0.106184f
C77 VTAIL.n3 B 0.78776f
C78 VTAIL.n4 B 1.60184f
C79 VTAIL.t0 B 0.106184f
C80 VTAIL.t1 B 0.106184f
C81 VTAIL.n5 B 0.787764f
C82 VTAIL.n6 B 1.60184f
C83 VTAIL.t3 B 1.0041f
C84 VTAIL.n7 B 0.667684f
C85 VTAIL.t9 B 0.106184f
C86 VTAIL.t7 B 0.106184f
C87 VTAIL.n8 B 0.787764f
C88 VTAIL.n9 B 0.594428f
C89 VTAIL.t8 B 1.0041f
C90 VTAIL.n10 B 1.47759f
C91 VTAIL.t2 B 1.0041f
C92 VTAIL.n11 B 1.42296f
C93 VP.n0 B 0.040131f
C94 VP.t2 B 0.842122f
C95 VP.n1 B 0.024742f
C96 VP.n2 B 0.030441f
C97 VP.t1 B 0.842122f
C98 VP.n3 B 0.060705f
C99 VP.n4 B 0.030441f
C100 VP.t0 B 0.842122f
C101 VP.n5 B 0.421778f
C102 VP.n6 B 0.040131f
C103 VP.t3 B 0.842122f
C104 VP.n7 B 0.024742f
C105 VP.n8 B 0.259428f
C106 VP.t4 B 0.842122f
C107 VP.t5 B 1.03134f
C108 VP.n9 B 0.396681f
C109 VP.n10 B 0.4078f
C110 VP.n11 B 0.042516f
C111 VP.n12 B 0.060705f
C112 VP.n13 B 0.030441f
C113 VP.n14 B 0.030441f
C114 VP.n15 B 0.030441f
C115 VP.n16 B 0.059505f
C116 VP.n17 B 0.044745f
C117 VP.n18 B 0.421778f
C118 VP.n19 B 1.27189f
C119 VP.n20 B 1.29822f
C120 VP.n21 B 0.040131f
C121 VP.n22 B 0.044745f
C122 VP.n23 B 0.059505f
C123 VP.n24 B 0.024742f
C124 VP.n25 B 0.030441f
C125 VP.n26 B 0.030441f
C126 VP.n27 B 0.030441f
C127 VP.n28 B 0.042516f
C128 VP.n29 B 0.329524f
C129 VP.n30 B 0.042516f
C130 VP.n31 B 0.060705f
C131 VP.n32 B 0.030441f
C132 VP.n33 B 0.030441f
C133 VP.n34 B 0.030441f
C134 VP.n35 B 0.059505f
C135 VP.n36 B 0.044745f
C136 VP.n37 B 0.421778f
C137 VP.n38 B 0.042886f
.ends

