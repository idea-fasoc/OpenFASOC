* NGSPICE file created from diff_pair_sample_0325.ext - technology: sky130A

.subckt diff_pair_sample_0325 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t14 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=2.31 ps=14.33 w=14 l=0.6
X1 B.t11 B.t9 B.t10 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=0.6
X2 VDD2.t8 VN.t1 VTAIL.t11 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=2.31 ps=14.33 w=14 l=0.6
X3 VDD1.t9 VP.t0 VTAIL.t2 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X4 VDD1.t8 VP.t1 VTAIL.t1 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=5.46 ps=28.78 w=14 l=0.6
X5 VTAIL.t10 VN.t2 VDD2.t7 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X6 VDD2.t6 VN.t3 VTAIL.t12 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X7 VTAIL.t3 VP.t2 VDD1.t7 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X8 VDD2.t5 VN.t4 VTAIL.t8 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=5.46 ps=28.78 w=14 l=0.6
X9 VTAIL.t15 VN.t5 VDD2.t4 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X10 VDD1.t6 VP.t3 VTAIL.t5 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X11 VTAIL.t7 VP.t4 VDD1.t5 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X12 VTAIL.t16 VN.t6 VDD2.t3 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X13 VDD1.t4 VP.t5 VTAIL.t4 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=5.46 ps=28.78 w=14 l=0.6
X14 VDD1.t3 VP.t6 VTAIL.t18 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=2.31 ps=14.33 w=14 l=0.6
X15 VTAIL.t6 VP.t7 VDD1.t2 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X16 B.t8 B.t6 B.t7 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=0.6
X17 VDD1.t1 VP.t8 VTAIL.t0 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=2.31 ps=14.33 w=14 l=0.6
X18 B.t5 B.t3 B.t4 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=0.6
X19 VDD2.t2 VN.t7 VTAIL.t17 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=5.46 ps=28.78 w=14 l=0.6
X20 VTAIL.t13 VN.t8 VDD2.t1 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X21 B.t2 B.t0 B.t1 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=5.46 pd=28.78 as=0 ps=0 w=14 l=0.6
X22 VDD2.t0 VN.t9 VTAIL.t9 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
X23 VTAIL.t19 VP.t9 VDD1.t0 w_n2086_n3768# sky130_fd_pr__pfet_01v8 ad=2.31 pd=14.33 as=2.31 ps=14.33 w=14 l=0.6
R0 VN.n3 VN.t1 654.006
R1 VN.n13 VN.t4 654.006
R2 VN.n2 VN.t8 627.806
R3 VN.n1 VN.t9 627.806
R4 VN.n6 VN.t6 627.806
R5 VN.n8 VN.t7 627.806
R6 VN.n12 VN.t5 627.806
R7 VN.n11 VN.t3 627.806
R8 VN.n16 VN.t2 627.806
R9 VN.n18 VN.t0 627.806
R10 VN.n9 VN.n8 161.3
R11 VN.n19 VN.n18 161.3
R12 VN.n17 VN.n10 161.3
R13 VN.n16 VN.n15 161.3
R14 VN.n7 VN.n0 161.3
R15 VN.n6 VN.n5 161.3
R16 VN.n14 VN.n11 80.6037
R17 VN.n4 VN.n1 80.6037
R18 VN.n2 VN.n1 48.2005
R19 VN.n6 VN.n1 48.2005
R20 VN.n12 VN.n11 48.2005
R21 VN.n16 VN.n11 48.2005
R22 VN.n8 VN.n7 45.2793
R23 VN.n18 VN.n17 45.2793
R24 VN.n14 VN.n13 45.1669
R25 VN.n4 VN.n3 45.1669
R26 VN VN.n19 44.1501
R27 VN.n3 VN.n2 14.3992
R28 VN.n13 VN.n12 14.3992
R29 VN.n7 VN.n6 2.92171
R30 VN.n17 VN.n16 2.92171
R31 VN.n15 VN.n14 0.285035
R32 VN.n5 VN.n4 0.285035
R33 VN.n19 VN.n10 0.189894
R34 VN.n15 VN.n10 0.189894
R35 VN.n5 VN.n0 0.189894
R36 VN.n9 VN.n0 0.189894
R37 VN VN.n9 0.0516364
R38 VTAIL.n320 VTAIL.n248 756.745
R39 VTAIL.n74 VTAIL.n2 756.745
R40 VTAIL.n242 VTAIL.n170 756.745
R41 VTAIL.n160 VTAIL.n88 756.745
R42 VTAIL.n272 VTAIL.n271 585
R43 VTAIL.n277 VTAIL.n276 585
R44 VTAIL.n279 VTAIL.n278 585
R45 VTAIL.n268 VTAIL.n267 585
R46 VTAIL.n285 VTAIL.n284 585
R47 VTAIL.n287 VTAIL.n286 585
R48 VTAIL.n264 VTAIL.n263 585
R49 VTAIL.n293 VTAIL.n292 585
R50 VTAIL.n295 VTAIL.n294 585
R51 VTAIL.n260 VTAIL.n259 585
R52 VTAIL.n301 VTAIL.n300 585
R53 VTAIL.n303 VTAIL.n302 585
R54 VTAIL.n256 VTAIL.n255 585
R55 VTAIL.n309 VTAIL.n308 585
R56 VTAIL.n311 VTAIL.n310 585
R57 VTAIL.n252 VTAIL.n251 585
R58 VTAIL.n318 VTAIL.n317 585
R59 VTAIL.n319 VTAIL.n250 585
R60 VTAIL.n321 VTAIL.n320 585
R61 VTAIL.n26 VTAIL.n25 585
R62 VTAIL.n31 VTAIL.n30 585
R63 VTAIL.n33 VTAIL.n32 585
R64 VTAIL.n22 VTAIL.n21 585
R65 VTAIL.n39 VTAIL.n38 585
R66 VTAIL.n41 VTAIL.n40 585
R67 VTAIL.n18 VTAIL.n17 585
R68 VTAIL.n47 VTAIL.n46 585
R69 VTAIL.n49 VTAIL.n48 585
R70 VTAIL.n14 VTAIL.n13 585
R71 VTAIL.n55 VTAIL.n54 585
R72 VTAIL.n57 VTAIL.n56 585
R73 VTAIL.n10 VTAIL.n9 585
R74 VTAIL.n63 VTAIL.n62 585
R75 VTAIL.n65 VTAIL.n64 585
R76 VTAIL.n6 VTAIL.n5 585
R77 VTAIL.n72 VTAIL.n71 585
R78 VTAIL.n73 VTAIL.n4 585
R79 VTAIL.n75 VTAIL.n74 585
R80 VTAIL.n243 VTAIL.n242 585
R81 VTAIL.n241 VTAIL.n172 585
R82 VTAIL.n240 VTAIL.n239 585
R83 VTAIL.n175 VTAIL.n173 585
R84 VTAIL.n234 VTAIL.n233 585
R85 VTAIL.n232 VTAIL.n231 585
R86 VTAIL.n179 VTAIL.n178 585
R87 VTAIL.n226 VTAIL.n225 585
R88 VTAIL.n224 VTAIL.n223 585
R89 VTAIL.n183 VTAIL.n182 585
R90 VTAIL.n218 VTAIL.n217 585
R91 VTAIL.n216 VTAIL.n215 585
R92 VTAIL.n187 VTAIL.n186 585
R93 VTAIL.n210 VTAIL.n209 585
R94 VTAIL.n208 VTAIL.n207 585
R95 VTAIL.n191 VTAIL.n190 585
R96 VTAIL.n202 VTAIL.n201 585
R97 VTAIL.n200 VTAIL.n199 585
R98 VTAIL.n195 VTAIL.n194 585
R99 VTAIL.n161 VTAIL.n160 585
R100 VTAIL.n159 VTAIL.n90 585
R101 VTAIL.n158 VTAIL.n157 585
R102 VTAIL.n93 VTAIL.n91 585
R103 VTAIL.n152 VTAIL.n151 585
R104 VTAIL.n150 VTAIL.n149 585
R105 VTAIL.n97 VTAIL.n96 585
R106 VTAIL.n144 VTAIL.n143 585
R107 VTAIL.n142 VTAIL.n141 585
R108 VTAIL.n101 VTAIL.n100 585
R109 VTAIL.n136 VTAIL.n135 585
R110 VTAIL.n134 VTAIL.n133 585
R111 VTAIL.n105 VTAIL.n104 585
R112 VTAIL.n128 VTAIL.n127 585
R113 VTAIL.n126 VTAIL.n125 585
R114 VTAIL.n109 VTAIL.n108 585
R115 VTAIL.n120 VTAIL.n119 585
R116 VTAIL.n118 VTAIL.n117 585
R117 VTAIL.n113 VTAIL.n112 585
R118 VTAIL.n273 VTAIL.t17 327.466
R119 VTAIL.n27 VTAIL.t4 327.466
R120 VTAIL.n196 VTAIL.t1 327.466
R121 VTAIL.n114 VTAIL.t8 327.466
R122 VTAIL.n277 VTAIL.n271 171.744
R123 VTAIL.n278 VTAIL.n277 171.744
R124 VTAIL.n278 VTAIL.n267 171.744
R125 VTAIL.n285 VTAIL.n267 171.744
R126 VTAIL.n286 VTAIL.n285 171.744
R127 VTAIL.n286 VTAIL.n263 171.744
R128 VTAIL.n293 VTAIL.n263 171.744
R129 VTAIL.n294 VTAIL.n293 171.744
R130 VTAIL.n294 VTAIL.n259 171.744
R131 VTAIL.n301 VTAIL.n259 171.744
R132 VTAIL.n302 VTAIL.n301 171.744
R133 VTAIL.n302 VTAIL.n255 171.744
R134 VTAIL.n309 VTAIL.n255 171.744
R135 VTAIL.n310 VTAIL.n309 171.744
R136 VTAIL.n310 VTAIL.n251 171.744
R137 VTAIL.n318 VTAIL.n251 171.744
R138 VTAIL.n319 VTAIL.n318 171.744
R139 VTAIL.n320 VTAIL.n319 171.744
R140 VTAIL.n31 VTAIL.n25 171.744
R141 VTAIL.n32 VTAIL.n31 171.744
R142 VTAIL.n32 VTAIL.n21 171.744
R143 VTAIL.n39 VTAIL.n21 171.744
R144 VTAIL.n40 VTAIL.n39 171.744
R145 VTAIL.n40 VTAIL.n17 171.744
R146 VTAIL.n47 VTAIL.n17 171.744
R147 VTAIL.n48 VTAIL.n47 171.744
R148 VTAIL.n48 VTAIL.n13 171.744
R149 VTAIL.n55 VTAIL.n13 171.744
R150 VTAIL.n56 VTAIL.n55 171.744
R151 VTAIL.n56 VTAIL.n9 171.744
R152 VTAIL.n63 VTAIL.n9 171.744
R153 VTAIL.n64 VTAIL.n63 171.744
R154 VTAIL.n64 VTAIL.n5 171.744
R155 VTAIL.n72 VTAIL.n5 171.744
R156 VTAIL.n73 VTAIL.n72 171.744
R157 VTAIL.n74 VTAIL.n73 171.744
R158 VTAIL.n242 VTAIL.n241 171.744
R159 VTAIL.n241 VTAIL.n240 171.744
R160 VTAIL.n240 VTAIL.n173 171.744
R161 VTAIL.n233 VTAIL.n173 171.744
R162 VTAIL.n233 VTAIL.n232 171.744
R163 VTAIL.n232 VTAIL.n178 171.744
R164 VTAIL.n225 VTAIL.n178 171.744
R165 VTAIL.n225 VTAIL.n224 171.744
R166 VTAIL.n224 VTAIL.n182 171.744
R167 VTAIL.n217 VTAIL.n182 171.744
R168 VTAIL.n217 VTAIL.n216 171.744
R169 VTAIL.n216 VTAIL.n186 171.744
R170 VTAIL.n209 VTAIL.n186 171.744
R171 VTAIL.n209 VTAIL.n208 171.744
R172 VTAIL.n208 VTAIL.n190 171.744
R173 VTAIL.n201 VTAIL.n190 171.744
R174 VTAIL.n201 VTAIL.n200 171.744
R175 VTAIL.n200 VTAIL.n194 171.744
R176 VTAIL.n160 VTAIL.n159 171.744
R177 VTAIL.n159 VTAIL.n158 171.744
R178 VTAIL.n158 VTAIL.n91 171.744
R179 VTAIL.n151 VTAIL.n91 171.744
R180 VTAIL.n151 VTAIL.n150 171.744
R181 VTAIL.n150 VTAIL.n96 171.744
R182 VTAIL.n143 VTAIL.n96 171.744
R183 VTAIL.n143 VTAIL.n142 171.744
R184 VTAIL.n142 VTAIL.n100 171.744
R185 VTAIL.n135 VTAIL.n100 171.744
R186 VTAIL.n135 VTAIL.n134 171.744
R187 VTAIL.n134 VTAIL.n104 171.744
R188 VTAIL.n127 VTAIL.n104 171.744
R189 VTAIL.n127 VTAIL.n126 171.744
R190 VTAIL.n126 VTAIL.n108 171.744
R191 VTAIL.n119 VTAIL.n108 171.744
R192 VTAIL.n119 VTAIL.n118 171.744
R193 VTAIL.n118 VTAIL.n112 171.744
R194 VTAIL.t17 VTAIL.n271 85.8723
R195 VTAIL.t4 VTAIL.n25 85.8723
R196 VTAIL.t1 VTAIL.n194 85.8723
R197 VTAIL.t8 VTAIL.n112 85.8723
R198 VTAIL.n169 VTAIL.n168 56.207
R199 VTAIL.n167 VTAIL.n166 56.207
R200 VTAIL.n87 VTAIL.n86 56.207
R201 VTAIL.n85 VTAIL.n84 56.207
R202 VTAIL.n327 VTAIL.n326 56.2069
R203 VTAIL.n1 VTAIL.n0 56.2069
R204 VTAIL.n81 VTAIL.n80 56.2069
R205 VTAIL.n83 VTAIL.n82 56.2069
R206 VTAIL.n325 VTAIL.n324 33.7369
R207 VTAIL.n79 VTAIL.n78 33.7369
R208 VTAIL.n247 VTAIL.n246 33.7369
R209 VTAIL.n165 VTAIL.n164 33.7369
R210 VTAIL.n85 VTAIL.n83 26.0393
R211 VTAIL.n325 VTAIL.n247 25.2376
R212 VTAIL.n273 VTAIL.n272 16.3895
R213 VTAIL.n27 VTAIL.n26 16.3895
R214 VTAIL.n196 VTAIL.n195 16.3895
R215 VTAIL.n114 VTAIL.n113 16.3895
R216 VTAIL.n321 VTAIL.n250 13.1884
R217 VTAIL.n75 VTAIL.n4 13.1884
R218 VTAIL.n243 VTAIL.n172 13.1884
R219 VTAIL.n161 VTAIL.n90 13.1884
R220 VTAIL.n276 VTAIL.n275 12.8005
R221 VTAIL.n317 VTAIL.n316 12.8005
R222 VTAIL.n322 VTAIL.n248 12.8005
R223 VTAIL.n30 VTAIL.n29 12.8005
R224 VTAIL.n71 VTAIL.n70 12.8005
R225 VTAIL.n76 VTAIL.n2 12.8005
R226 VTAIL.n244 VTAIL.n170 12.8005
R227 VTAIL.n239 VTAIL.n174 12.8005
R228 VTAIL.n199 VTAIL.n198 12.8005
R229 VTAIL.n162 VTAIL.n88 12.8005
R230 VTAIL.n157 VTAIL.n92 12.8005
R231 VTAIL.n117 VTAIL.n116 12.8005
R232 VTAIL.n279 VTAIL.n270 12.0247
R233 VTAIL.n315 VTAIL.n252 12.0247
R234 VTAIL.n33 VTAIL.n24 12.0247
R235 VTAIL.n69 VTAIL.n6 12.0247
R236 VTAIL.n238 VTAIL.n175 12.0247
R237 VTAIL.n202 VTAIL.n193 12.0247
R238 VTAIL.n156 VTAIL.n93 12.0247
R239 VTAIL.n120 VTAIL.n111 12.0247
R240 VTAIL.n280 VTAIL.n268 11.249
R241 VTAIL.n312 VTAIL.n311 11.249
R242 VTAIL.n34 VTAIL.n22 11.249
R243 VTAIL.n66 VTAIL.n65 11.249
R244 VTAIL.n235 VTAIL.n234 11.249
R245 VTAIL.n203 VTAIL.n191 11.249
R246 VTAIL.n153 VTAIL.n152 11.249
R247 VTAIL.n121 VTAIL.n109 11.249
R248 VTAIL.n284 VTAIL.n283 10.4732
R249 VTAIL.n308 VTAIL.n254 10.4732
R250 VTAIL.n38 VTAIL.n37 10.4732
R251 VTAIL.n62 VTAIL.n8 10.4732
R252 VTAIL.n231 VTAIL.n177 10.4732
R253 VTAIL.n207 VTAIL.n206 10.4732
R254 VTAIL.n149 VTAIL.n95 10.4732
R255 VTAIL.n125 VTAIL.n124 10.4732
R256 VTAIL.n287 VTAIL.n266 9.69747
R257 VTAIL.n307 VTAIL.n256 9.69747
R258 VTAIL.n41 VTAIL.n20 9.69747
R259 VTAIL.n61 VTAIL.n10 9.69747
R260 VTAIL.n230 VTAIL.n179 9.69747
R261 VTAIL.n210 VTAIL.n189 9.69747
R262 VTAIL.n148 VTAIL.n97 9.69747
R263 VTAIL.n128 VTAIL.n107 9.69747
R264 VTAIL.n324 VTAIL.n323 9.45567
R265 VTAIL.n78 VTAIL.n77 9.45567
R266 VTAIL.n246 VTAIL.n245 9.45567
R267 VTAIL.n164 VTAIL.n163 9.45567
R268 VTAIL.n323 VTAIL.n322 9.3005
R269 VTAIL.n262 VTAIL.n261 9.3005
R270 VTAIL.n291 VTAIL.n290 9.3005
R271 VTAIL.n289 VTAIL.n288 9.3005
R272 VTAIL.n266 VTAIL.n265 9.3005
R273 VTAIL.n283 VTAIL.n282 9.3005
R274 VTAIL.n281 VTAIL.n280 9.3005
R275 VTAIL.n270 VTAIL.n269 9.3005
R276 VTAIL.n275 VTAIL.n274 9.3005
R277 VTAIL.n297 VTAIL.n296 9.3005
R278 VTAIL.n299 VTAIL.n298 9.3005
R279 VTAIL.n258 VTAIL.n257 9.3005
R280 VTAIL.n305 VTAIL.n304 9.3005
R281 VTAIL.n307 VTAIL.n306 9.3005
R282 VTAIL.n254 VTAIL.n253 9.3005
R283 VTAIL.n313 VTAIL.n312 9.3005
R284 VTAIL.n315 VTAIL.n314 9.3005
R285 VTAIL.n316 VTAIL.n249 9.3005
R286 VTAIL.n77 VTAIL.n76 9.3005
R287 VTAIL.n16 VTAIL.n15 9.3005
R288 VTAIL.n45 VTAIL.n44 9.3005
R289 VTAIL.n43 VTAIL.n42 9.3005
R290 VTAIL.n20 VTAIL.n19 9.3005
R291 VTAIL.n37 VTAIL.n36 9.3005
R292 VTAIL.n35 VTAIL.n34 9.3005
R293 VTAIL.n24 VTAIL.n23 9.3005
R294 VTAIL.n29 VTAIL.n28 9.3005
R295 VTAIL.n51 VTAIL.n50 9.3005
R296 VTAIL.n53 VTAIL.n52 9.3005
R297 VTAIL.n12 VTAIL.n11 9.3005
R298 VTAIL.n59 VTAIL.n58 9.3005
R299 VTAIL.n61 VTAIL.n60 9.3005
R300 VTAIL.n8 VTAIL.n7 9.3005
R301 VTAIL.n67 VTAIL.n66 9.3005
R302 VTAIL.n69 VTAIL.n68 9.3005
R303 VTAIL.n70 VTAIL.n3 9.3005
R304 VTAIL.n222 VTAIL.n221 9.3005
R305 VTAIL.n181 VTAIL.n180 9.3005
R306 VTAIL.n228 VTAIL.n227 9.3005
R307 VTAIL.n230 VTAIL.n229 9.3005
R308 VTAIL.n177 VTAIL.n176 9.3005
R309 VTAIL.n236 VTAIL.n235 9.3005
R310 VTAIL.n238 VTAIL.n237 9.3005
R311 VTAIL.n174 VTAIL.n171 9.3005
R312 VTAIL.n245 VTAIL.n244 9.3005
R313 VTAIL.n220 VTAIL.n219 9.3005
R314 VTAIL.n185 VTAIL.n184 9.3005
R315 VTAIL.n214 VTAIL.n213 9.3005
R316 VTAIL.n212 VTAIL.n211 9.3005
R317 VTAIL.n189 VTAIL.n188 9.3005
R318 VTAIL.n206 VTAIL.n205 9.3005
R319 VTAIL.n204 VTAIL.n203 9.3005
R320 VTAIL.n193 VTAIL.n192 9.3005
R321 VTAIL.n198 VTAIL.n197 9.3005
R322 VTAIL.n140 VTAIL.n139 9.3005
R323 VTAIL.n99 VTAIL.n98 9.3005
R324 VTAIL.n146 VTAIL.n145 9.3005
R325 VTAIL.n148 VTAIL.n147 9.3005
R326 VTAIL.n95 VTAIL.n94 9.3005
R327 VTAIL.n154 VTAIL.n153 9.3005
R328 VTAIL.n156 VTAIL.n155 9.3005
R329 VTAIL.n92 VTAIL.n89 9.3005
R330 VTAIL.n163 VTAIL.n162 9.3005
R331 VTAIL.n138 VTAIL.n137 9.3005
R332 VTAIL.n103 VTAIL.n102 9.3005
R333 VTAIL.n132 VTAIL.n131 9.3005
R334 VTAIL.n130 VTAIL.n129 9.3005
R335 VTAIL.n107 VTAIL.n106 9.3005
R336 VTAIL.n124 VTAIL.n123 9.3005
R337 VTAIL.n122 VTAIL.n121 9.3005
R338 VTAIL.n111 VTAIL.n110 9.3005
R339 VTAIL.n116 VTAIL.n115 9.3005
R340 VTAIL.n288 VTAIL.n264 8.92171
R341 VTAIL.n304 VTAIL.n303 8.92171
R342 VTAIL.n42 VTAIL.n18 8.92171
R343 VTAIL.n58 VTAIL.n57 8.92171
R344 VTAIL.n227 VTAIL.n226 8.92171
R345 VTAIL.n211 VTAIL.n187 8.92171
R346 VTAIL.n145 VTAIL.n144 8.92171
R347 VTAIL.n129 VTAIL.n105 8.92171
R348 VTAIL.n292 VTAIL.n291 8.14595
R349 VTAIL.n300 VTAIL.n258 8.14595
R350 VTAIL.n46 VTAIL.n45 8.14595
R351 VTAIL.n54 VTAIL.n12 8.14595
R352 VTAIL.n223 VTAIL.n181 8.14595
R353 VTAIL.n215 VTAIL.n214 8.14595
R354 VTAIL.n141 VTAIL.n99 8.14595
R355 VTAIL.n133 VTAIL.n132 8.14595
R356 VTAIL.n295 VTAIL.n262 7.3702
R357 VTAIL.n299 VTAIL.n260 7.3702
R358 VTAIL.n49 VTAIL.n16 7.3702
R359 VTAIL.n53 VTAIL.n14 7.3702
R360 VTAIL.n222 VTAIL.n183 7.3702
R361 VTAIL.n218 VTAIL.n185 7.3702
R362 VTAIL.n140 VTAIL.n101 7.3702
R363 VTAIL.n136 VTAIL.n103 7.3702
R364 VTAIL.n296 VTAIL.n295 6.59444
R365 VTAIL.n296 VTAIL.n260 6.59444
R366 VTAIL.n50 VTAIL.n49 6.59444
R367 VTAIL.n50 VTAIL.n14 6.59444
R368 VTAIL.n219 VTAIL.n183 6.59444
R369 VTAIL.n219 VTAIL.n218 6.59444
R370 VTAIL.n137 VTAIL.n101 6.59444
R371 VTAIL.n137 VTAIL.n136 6.59444
R372 VTAIL.n292 VTAIL.n262 5.81868
R373 VTAIL.n300 VTAIL.n299 5.81868
R374 VTAIL.n46 VTAIL.n16 5.81868
R375 VTAIL.n54 VTAIL.n53 5.81868
R376 VTAIL.n223 VTAIL.n222 5.81868
R377 VTAIL.n215 VTAIL.n185 5.81868
R378 VTAIL.n141 VTAIL.n140 5.81868
R379 VTAIL.n133 VTAIL.n103 5.81868
R380 VTAIL.n291 VTAIL.n264 5.04292
R381 VTAIL.n303 VTAIL.n258 5.04292
R382 VTAIL.n45 VTAIL.n18 5.04292
R383 VTAIL.n57 VTAIL.n12 5.04292
R384 VTAIL.n226 VTAIL.n181 5.04292
R385 VTAIL.n214 VTAIL.n187 5.04292
R386 VTAIL.n144 VTAIL.n99 5.04292
R387 VTAIL.n132 VTAIL.n105 5.04292
R388 VTAIL.n288 VTAIL.n287 4.26717
R389 VTAIL.n304 VTAIL.n256 4.26717
R390 VTAIL.n42 VTAIL.n41 4.26717
R391 VTAIL.n58 VTAIL.n10 4.26717
R392 VTAIL.n227 VTAIL.n179 4.26717
R393 VTAIL.n211 VTAIL.n210 4.26717
R394 VTAIL.n145 VTAIL.n97 4.26717
R395 VTAIL.n129 VTAIL.n128 4.26717
R396 VTAIL.n274 VTAIL.n273 3.70982
R397 VTAIL.n28 VTAIL.n27 3.70982
R398 VTAIL.n197 VTAIL.n196 3.70982
R399 VTAIL.n115 VTAIL.n114 3.70982
R400 VTAIL.n284 VTAIL.n266 3.49141
R401 VTAIL.n308 VTAIL.n307 3.49141
R402 VTAIL.n38 VTAIL.n20 3.49141
R403 VTAIL.n62 VTAIL.n61 3.49141
R404 VTAIL.n231 VTAIL.n230 3.49141
R405 VTAIL.n207 VTAIL.n189 3.49141
R406 VTAIL.n149 VTAIL.n148 3.49141
R407 VTAIL.n125 VTAIL.n107 3.49141
R408 VTAIL.n283 VTAIL.n268 2.71565
R409 VTAIL.n311 VTAIL.n254 2.71565
R410 VTAIL.n37 VTAIL.n22 2.71565
R411 VTAIL.n65 VTAIL.n8 2.71565
R412 VTAIL.n234 VTAIL.n177 2.71565
R413 VTAIL.n206 VTAIL.n191 2.71565
R414 VTAIL.n152 VTAIL.n95 2.71565
R415 VTAIL.n124 VTAIL.n109 2.71565
R416 VTAIL.n326 VTAIL.t9 2.32229
R417 VTAIL.n326 VTAIL.t16 2.32229
R418 VTAIL.n0 VTAIL.t11 2.32229
R419 VTAIL.n0 VTAIL.t13 2.32229
R420 VTAIL.n80 VTAIL.t2 2.32229
R421 VTAIL.n80 VTAIL.t19 2.32229
R422 VTAIL.n82 VTAIL.t0 2.32229
R423 VTAIL.n82 VTAIL.t6 2.32229
R424 VTAIL.n168 VTAIL.t5 2.32229
R425 VTAIL.n168 VTAIL.t3 2.32229
R426 VTAIL.n166 VTAIL.t18 2.32229
R427 VTAIL.n166 VTAIL.t7 2.32229
R428 VTAIL.n86 VTAIL.t12 2.32229
R429 VTAIL.n86 VTAIL.t15 2.32229
R430 VTAIL.n84 VTAIL.t14 2.32229
R431 VTAIL.n84 VTAIL.t10 2.32229
R432 VTAIL.n280 VTAIL.n279 1.93989
R433 VTAIL.n312 VTAIL.n252 1.93989
R434 VTAIL.n34 VTAIL.n33 1.93989
R435 VTAIL.n66 VTAIL.n6 1.93989
R436 VTAIL.n235 VTAIL.n175 1.93989
R437 VTAIL.n203 VTAIL.n202 1.93989
R438 VTAIL.n153 VTAIL.n93 1.93989
R439 VTAIL.n121 VTAIL.n120 1.93989
R440 VTAIL.n276 VTAIL.n270 1.16414
R441 VTAIL.n317 VTAIL.n315 1.16414
R442 VTAIL.n324 VTAIL.n248 1.16414
R443 VTAIL.n30 VTAIL.n24 1.16414
R444 VTAIL.n71 VTAIL.n69 1.16414
R445 VTAIL.n78 VTAIL.n2 1.16414
R446 VTAIL.n246 VTAIL.n170 1.16414
R447 VTAIL.n239 VTAIL.n238 1.16414
R448 VTAIL.n199 VTAIL.n193 1.16414
R449 VTAIL.n164 VTAIL.n88 1.16414
R450 VTAIL.n157 VTAIL.n156 1.16414
R451 VTAIL.n117 VTAIL.n111 1.16414
R452 VTAIL.n167 VTAIL.n165 0.87119
R453 VTAIL.n79 VTAIL.n1 0.87119
R454 VTAIL.n87 VTAIL.n85 0.802224
R455 VTAIL.n165 VTAIL.n87 0.802224
R456 VTAIL.n169 VTAIL.n167 0.802224
R457 VTAIL.n247 VTAIL.n169 0.802224
R458 VTAIL.n83 VTAIL.n81 0.802224
R459 VTAIL.n81 VTAIL.n79 0.802224
R460 VTAIL.n327 VTAIL.n325 0.802224
R461 VTAIL VTAIL.n1 0.659983
R462 VTAIL.n275 VTAIL.n272 0.388379
R463 VTAIL.n316 VTAIL.n250 0.388379
R464 VTAIL.n322 VTAIL.n321 0.388379
R465 VTAIL.n29 VTAIL.n26 0.388379
R466 VTAIL.n70 VTAIL.n4 0.388379
R467 VTAIL.n76 VTAIL.n75 0.388379
R468 VTAIL.n244 VTAIL.n243 0.388379
R469 VTAIL.n174 VTAIL.n172 0.388379
R470 VTAIL.n198 VTAIL.n195 0.388379
R471 VTAIL.n162 VTAIL.n161 0.388379
R472 VTAIL.n92 VTAIL.n90 0.388379
R473 VTAIL.n116 VTAIL.n113 0.388379
R474 VTAIL.n274 VTAIL.n269 0.155672
R475 VTAIL.n281 VTAIL.n269 0.155672
R476 VTAIL.n282 VTAIL.n281 0.155672
R477 VTAIL.n282 VTAIL.n265 0.155672
R478 VTAIL.n289 VTAIL.n265 0.155672
R479 VTAIL.n290 VTAIL.n289 0.155672
R480 VTAIL.n290 VTAIL.n261 0.155672
R481 VTAIL.n297 VTAIL.n261 0.155672
R482 VTAIL.n298 VTAIL.n297 0.155672
R483 VTAIL.n298 VTAIL.n257 0.155672
R484 VTAIL.n305 VTAIL.n257 0.155672
R485 VTAIL.n306 VTAIL.n305 0.155672
R486 VTAIL.n306 VTAIL.n253 0.155672
R487 VTAIL.n313 VTAIL.n253 0.155672
R488 VTAIL.n314 VTAIL.n313 0.155672
R489 VTAIL.n314 VTAIL.n249 0.155672
R490 VTAIL.n323 VTAIL.n249 0.155672
R491 VTAIL.n28 VTAIL.n23 0.155672
R492 VTAIL.n35 VTAIL.n23 0.155672
R493 VTAIL.n36 VTAIL.n35 0.155672
R494 VTAIL.n36 VTAIL.n19 0.155672
R495 VTAIL.n43 VTAIL.n19 0.155672
R496 VTAIL.n44 VTAIL.n43 0.155672
R497 VTAIL.n44 VTAIL.n15 0.155672
R498 VTAIL.n51 VTAIL.n15 0.155672
R499 VTAIL.n52 VTAIL.n51 0.155672
R500 VTAIL.n52 VTAIL.n11 0.155672
R501 VTAIL.n59 VTAIL.n11 0.155672
R502 VTAIL.n60 VTAIL.n59 0.155672
R503 VTAIL.n60 VTAIL.n7 0.155672
R504 VTAIL.n67 VTAIL.n7 0.155672
R505 VTAIL.n68 VTAIL.n67 0.155672
R506 VTAIL.n68 VTAIL.n3 0.155672
R507 VTAIL.n77 VTAIL.n3 0.155672
R508 VTAIL.n245 VTAIL.n171 0.155672
R509 VTAIL.n237 VTAIL.n171 0.155672
R510 VTAIL.n237 VTAIL.n236 0.155672
R511 VTAIL.n236 VTAIL.n176 0.155672
R512 VTAIL.n229 VTAIL.n176 0.155672
R513 VTAIL.n229 VTAIL.n228 0.155672
R514 VTAIL.n228 VTAIL.n180 0.155672
R515 VTAIL.n221 VTAIL.n180 0.155672
R516 VTAIL.n221 VTAIL.n220 0.155672
R517 VTAIL.n220 VTAIL.n184 0.155672
R518 VTAIL.n213 VTAIL.n184 0.155672
R519 VTAIL.n213 VTAIL.n212 0.155672
R520 VTAIL.n212 VTAIL.n188 0.155672
R521 VTAIL.n205 VTAIL.n188 0.155672
R522 VTAIL.n205 VTAIL.n204 0.155672
R523 VTAIL.n204 VTAIL.n192 0.155672
R524 VTAIL.n197 VTAIL.n192 0.155672
R525 VTAIL.n163 VTAIL.n89 0.155672
R526 VTAIL.n155 VTAIL.n89 0.155672
R527 VTAIL.n155 VTAIL.n154 0.155672
R528 VTAIL.n154 VTAIL.n94 0.155672
R529 VTAIL.n147 VTAIL.n94 0.155672
R530 VTAIL.n147 VTAIL.n146 0.155672
R531 VTAIL.n146 VTAIL.n98 0.155672
R532 VTAIL.n139 VTAIL.n98 0.155672
R533 VTAIL.n139 VTAIL.n138 0.155672
R534 VTAIL.n138 VTAIL.n102 0.155672
R535 VTAIL.n131 VTAIL.n102 0.155672
R536 VTAIL.n131 VTAIL.n130 0.155672
R537 VTAIL.n130 VTAIL.n106 0.155672
R538 VTAIL.n123 VTAIL.n106 0.155672
R539 VTAIL.n123 VTAIL.n122 0.155672
R540 VTAIL.n122 VTAIL.n110 0.155672
R541 VTAIL.n115 VTAIL.n110 0.155672
R542 VTAIL VTAIL.n327 0.142741
R543 VDD2.n153 VDD2.n81 756.745
R544 VDD2.n72 VDD2.n0 756.745
R545 VDD2.n154 VDD2.n153 585
R546 VDD2.n152 VDD2.n83 585
R547 VDD2.n151 VDD2.n150 585
R548 VDD2.n86 VDD2.n84 585
R549 VDD2.n145 VDD2.n144 585
R550 VDD2.n143 VDD2.n142 585
R551 VDD2.n90 VDD2.n89 585
R552 VDD2.n137 VDD2.n136 585
R553 VDD2.n135 VDD2.n134 585
R554 VDD2.n94 VDD2.n93 585
R555 VDD2.n129 VDD2.n128 585
R556 VDD2.n127 VDD2.n126 585
R557 VDD2.n98 VDD2.n97 585
R558 VDD2.n121 VDD2.n120 585
R559 VDD2.n119 VDD2.n118 585
R560 VDD2.n102 VDD2.n101 585
R561 VDD2.n113 VDD2.n112 585
R562 VDD2.n111 VDD2.n110 585
R563 VDD2.n106 VDD2.n105 585
R564 VDD2.n24 VDD2.n23 585
R565 VDD2.n29 VDD2.n28 585
R566 VDD2.n31 VDD2.n30 585
R567 VDD2.n20 VDD2.n19 585
R568 VDD2.n37 VDD2.n36 585
R569 VDD2.n39 VDD2.n38 585
R570 VDD2.n16 VDD2.n15 585
R571 VDD2.n45 VDD2.n44 585
R572 VDD2.n47 VDD2.n46 585
R573 VDD2.n12 VDD2.n11 585
R574 VDD2.n53 VDD2.n52 585
R575 VDD2.n55 VDD2.n54 585
R576 VDD2.n8 VDD2.n7 585
R577 VDD2.n61 VDD2.n60 585
R578 VDD2.n63 VDD2.n62 585
R579 VDD2.n4 VDD2.n3 585
R580 VDD2.n70 VDD2.n69 585
R581 VDD2.n71 VDD2.n2 585
R582 VDD2.n73 VDD2.n72 585
R583 VDD2.n107 VDD2.t9 327.466
R584 VDD2.n25 VDD2.t8 327.466
R585 VDD2.n153 VDD2.n152 171.744
R586 VDD2.n152 VDD2.n151 171.744
R587 VDD2.n151 VDD2.n84 171.744
R588 VDD2.n144 VDD2.n84 171.744
R589 VDD2.n144 VDD2.n143 171.744
R590 VDD2.n143 VDD2.n89 171.744
R591 VDD2.n136 VDD2.n89 171.744
R592 VDD2.n136 VDD2.n135 171.744
R593 VDD2.n135 VDD2.n93 171.744
R594 VDD2.n128 VDD2.n93 171.744
R595 VDD2.n128 VDD2.n127 171.744
R596 VDD2.n127 VDD2.n97 171.744
R597 VDD2.n120 VDD2.n97 171.744
R598 VDD2.n120 VDD2.n119 171.744
R599 VDD2.n119 VDD2.n101 171.744
R600 VDD2.n112 VDD2.n101 171.744
R601 VDD2.n112 VDD2.n111 171.744
R602 VDD2.n111 VDD2.n105 171.744
R603 VDD2.n29 VDD2.n23 171.744
R604 VDD2.n30 VDD2.n29 171.744
R605 VDD2.n30 VDD2.n19 171.744
R606 VDD2.n37 VDD2.n19 171.744
R607 VDD2.n38 VDD2.n37 171.744
R608 VDD2.n38 VDD2.n15 171.744
R609 VDD2.n45 VDD2.n15 171.744
R610 VDD2.n46 VDD2.n45 171.744
R611 VDD2.n46 VDD2.n11 171.744
R612 VDD2.n53 VDD2.n11 171.744
R613 VDD2.n54 VDD2.n53 171.744
R614 VDD2.n54 VDD2.n7 171.744
R615 VDD2.n61 VDD2.n7 171.744
R616 VDD2.n62 VDD2.n61 171.744
R617 VDD2.n62 VDD2.n3 171.744
R618 VDD2.n70 VDD2.n3 171.744
R619 VDD2.n71 VDD2.n70 171.744
R620 VDD2.n72 VDD2.n71 171.744
R621 VDD2.t9 VDD2.n105 85.8723
R622 VDD2.t8 VDD2.n23 85.8723
R623 VDD2.n80 VDD2.n79 73.4316
R624 VDD2 VDD2.n161 73.4288
R625 VDD2.n160 VDD2.n159 72.8858
R626 VDD2.n78 VDD2.n77 72.8856
R627 VDD2.n78 VDD2.n76 51.2174
R628 VDD2.n158 VDD2.n157 50.4157
R629 VDD2.n158 VDD2.n80 39.5925
R630 VDD2.n107 VDD2.n106 16.3895
R631 VDD2.n25 VDD2.n24 16.3895
R632 VDD2.n154 VDD2.n83 13.1884
R633 VDD2.n73 VDD2.n2 13.1884
R634 VDD2.n155 VDD2.n81 12.8005
R635 VDD2.n150 VDD2.n85 12.8005
R636 VDD2.n110 VDD2.n109 12.8005
R637 VDD2.n28 VDD2.n27 12.8005
R638 VDD2.n69 VDD2.n68 12.8005
R639 VDD2.n74 VDD2.n0 12.8005
R640 VDD2.n149 VDD2.n86 12.0247
R641 VDD2.n113 VDD2.n104 12.0247
R642 VDD2.n31 VDD2.n22 12.0247
R643 VDD2.n67 VDD2.n4 12.0247
R644 VDD2.n146 VDD2.n145 11.249
R645 VDD2.n114 VDD2.n102 11.249
R646 VDD2.n32 VDD2.n20 11.249
R647 VDD2.n64 VDD2.n63 11.249
R648 VDD2.n142 VDD2.n88 10.4732
R649 VDD2.n118 VDD2.n117 10.4732
R650 VDD2.n36 VDD2.n35 10.4732
R651 VDD2.n60 VDD2.n6 10.4732
R652 VDD2.n141 VDD2.n90 9.69747
R653 VDD2.n121 VDD2.n100 9.69747
R654 VDD2.n39 VDD2.n18 9.69747
R655 VDD2.n59 VDD2.n8 9.69747
R656 VDD2.n157 VDD2.n156 9.45567
R657 VDD2.n76 VDD2.n75 9.45567
R658 VDD2.n133 VDD2.n132 9.3005
R659 VDD2.n92 VDD2.n91 9.3005
R660 VDD2.n139 VDD2.n138 9.3005
R661 VDD2.n141 VDD2.n140 9.3005
R662 VDD2.n88 VDD2.n87 9.3005
R663 VDD2.n147 VDD2.n146 9.3005
R664 VDD2.n149 VDD2.n148 9.3005
R665 VDD2.n85 VDD2.n82 9.3005
R666 VDD2.n156 VDD2.n155 9.3005
R667 VDD2.n131 VDD2.n130 9.3005
R668 VDD2.n96 VDD2.n95 9.3005
R669 VDD2.n125 VDD2.n124 9.3005
R670 VDD2.n123 VDD2.n122 9.3005
R671 VDD2.n100 VDD2.n99 9.3005
R672 VDD2.n117 VDD2.n116 9.3005
R673 VDD2.n115 VDD2.n114 9.3005
R674 VDD2.n104 VDD2.n103 9.3005
R675 VDD2.n109 VDD2.n108 9.3005
R676 VDD2.n75 VDD2.n74 9.3005
R677 VDD2.n14 VDD2.n13 9.3005
R678 VDD2.n43 VDD2.n42 9.3005
R679 VDD2.n41 VDD2.n40 9.3005
R680 VDD2.n18 VDD2.n17 9.3005
R681 VDD2.n35 VDD2.n34 9.3005
R682 VDD2.n33 VDD2.n32 9.3005
R683 VDD2.n22 VDD2.n21 9.3005
R684 VDD2.n27 VDD2.n26 9.3005
R685 VDD2.n49 VDD2.n48 9.3005
R686 VDD2.n51 VDD2.n50 9.3005
R687 VDD2.n10 VDD2.n9 9.3005
R688 VDD2.n57 VDD2.n56 9.3005
R689 VDD2.n59 VDD2.n58 9.3005
R690 VDD2.n6 VDD2.n5 9.3005
R691 VDD2.n65 VDD2.n64 9.3005
R692 VDD2.n67 VDD2.n66 9.3005
R693 VDD2.n68 VDD2.n1 9.3005
R694 VDD2.n138 VDD2.n137 8.92171
R695 VDD2.n122 VDD2.n98 8.92171
R696 VDD2.n40 VDD2.n16 8.92171
R697 VDD2.n56 VDD2.n55 8.92171
R698 VDD2.n134 VDD2.n92 8.14595
R699 VDD2.n126 VDD2.n125 8.14595
R700 VDD2.n44 VDD2.n43 8.14595
R701 VDD2.n52 VDD2.n10 8.14595
R702 VDD2.n133 VDD2.n94 7.3702
R703 VDD2.n129 VDD2.n96 7.3702
R704 VDD2.n47 VDD2.n14 7.3702
R705 VDD2.n51 VDD2.n12 7.3702
R706 VDD2.n130 VDD2.n94 6.59444
R707 VDD2.n130 VDD2.n129 6.59444
R708 VDD2.n48 VDD2.n47 6.59444
R709 VDD2.n48 VDD2.n12 6.59444
R710 VDD2.n134 VDD2.n133 5.81868
R711 VDD2.n126 VDD2.n96 5.81868
R712 VDD2.n44 VDD2.n14 5.81868
R713 VDD2.n52 VDD2.n51 5.81868
R714 VDD2.n137 VDD2.n92 5.04292
R715 VDD2.n125 VDD2.n98 5.04292
R716 VDD2.n43 VDD2.n16 5.04292
R717 VDD2.n55 VDD2.n10 5.04292
R718 VDD2.n138 VDD2.n90 4.26717
R719 VDD2.n122 VDD2.n121 4.26717
R720 VDD2.n40 VDD2.n39 4.26717
R721 VDD2.n56 VDD2.n8 4.26717
R722 VDD2.n108 VDD2.n107 3.70982
R723 VDD2.n26 VDD2.n25 3.70982
R724 VDD2.n142 VDD2.n141 3.49141
R725 VDD2.n118 VDD2.n100 3.49141
R726 VDD2.n36 VDD2.n18 3.49141
R727 VDD2.n60 VDD2.n59 3.49141
R728 VDD2.n145 VDD2.n88 2.71565
R729 VDD2.n117 VDD2.n102 2.71565
R730 VDD2.n35 VDD2.n20 2.71565
R731 VDD2.n63 VDD2.n6 2.71565
R732 VDD2.n161 VDD2.t4 2.32229
R733 VDD2.n161 VDD2.t5 2.32229
R734 VDD2.n159 VDD2.t7 2.32229
R735 VDD2.n159 VDD2.t6 2.32229
R736 VDD2.n79 VDD2.t3 2.32229
R737 VDD2.n79 VDD2.t2 2.32229
R738 VDD2.n77 VDD2.t1 2.32229
R739 VDD2.n77 VDD2.t0 2.32229
R740 VDD2.n146 VDD2.n86 1.93989
R741 VDD2.n114 VDD2.n113 1.93989
R742 VDD2.n32 VDD2.n31 1.93989
R743 VDD2.n64 VDD2.n4 1.93989
R744 VDD2.n157 VDD2.n81 1.16414
R745 VDD2.n150 VDD2.n149 1.16414
R746 VDD2.n110 VDD2.n104 1.16414
R747 VDD2.n28 VDD2.n22 1.16414
R748 VDD2.n69 VDD2.n67 1.16414
R749 VDD2.n76 VDD2.n0 1.16414
R750 VDD2.n160 VDD2.n158 0.802224
R751 VDD2.n155 VDD2.n154 0.388379
R752 VDD2.n85 VDD2.n83 0.388379
R753 VDD2.n109 VDD2.n106 0.388379
R754 VDD2.n27 VDD2.n24 0.388379
R755 VDD2.n68 VDD2.n2 0.388379
R756 VDD2.n74 VDD2.n73 0.388379
R757 VDD2 VDD2.n160 0.259121
R758 VDD2.n156 VDD2.n82 0.155672
R759 VDD2.n148 VDD2.n82 0.155672
R760 VDD2.n148 VDD2.n147 0.155672
R761 VDD2.n147 VDD2.n87 0.155672
R762 VDD2.n140 VDD2.n87 0.155672
R763 VDD2.n140 VDD2.n139 0.155672
R764 VDD2.n139 VDD2.n91 0.155672
R765 VDD2.n132 VDD2.n91 0.155672
R766 VDD2.n132 VDD2.n131 0.155672
R767 VDD2.n131 VDD2.n95 0.155672
R768 VDD2.n124 VDD2.n95 0.155672
R769 VDD2.n124 VDD2.n123 0.155672
R770 VDD2.n123 VDD2.n99 0.155672
R771 VDD2.n116 VDD2.n99 0.155672
R772 VDD2.n116 VDD2.n115 0.155672
R773 VDD2.n115 VDD2.n103 0.155672
R774 VDD2.n108 VDD2.n103 0.155672
R775 VDD2.n26 VDD2.n21 0.155672
R776 VDD2.n33 VDD2.n21 0.155672
R777 VDD2.n34 VDD2.n33 0.155672
R778 VDD2.n34 VDD2.n17 0.155672
R779 VDD2.n41 VDD2.n17 0.155672
R780 VDD2.n42 VDD2.n41 0.155672
R781 VDD2.n42 VDD2.n13 0.155672
R782 VDD2.n49 VDD2.n13 0.155672
R783 VDD2.n50 VDD2.n49 0.155672
R784 VDD2.n50 VDD2.n9 0.155672
R785 VDD2.n57 VDD2.n9 0.155672
R786 VDD2.n58 VDD2.n57 0.155672
R787 VDD2.n58 VDD2.n5 0.155672
R788 VDD2.n65 VDD2.n5 0.155672
R789 VDD2.n66 VDD2.n65 0.155672
R790 VDD2.n66 VDD2.n1 0.155672
R791 VDD2.n75 VDD2.n1 0.155672
R792 VDD2.n80 VDD2.n78 0.145585
R793 B.n128 B.t0 766.734
R794 B.n120 B.t9 766.734
R795 B.n46 B.t3 766.734
R796 B.n38 B.t6 766.734
R797 B.n357 B.n96 585
R798 B.n356 B.n355 585
R799 B.n354 B.n97 585
R800 B.n353 B.n352 585
R801 B.n351 B.n98 585
R802 B.n350 B.n349 585
R803 B.n348 B.n99 585
R804 B.n347 B.n346 585
R805 B.n345 B.n100 585
R806 B.n344 B.n343 585
R807 B.n342 B.n101 585
R808 B.n341 B.n340 585
R809 B.n339 B.n102 585
R810 B.n338 B.n337 585
R811 B.n336 B.n103 585
R812 B.n335 B.n334 585
R813 B.n333 B.n104 585
R814 B.n332 B.n331 585
R815 B.n330 B.n105 585
R816 B.n329 B.n328 585
R817 B.n327 B.n106 585
R818 B.n326 B.n325 585
R819 B.n324 B.n107 585
R820 B.n323 B.n322 585
R821 B.n321 B.n108 585
R822 B.n320 B.n319 585
R823 B.n318 B.n109 585
R824 B.n317 B.n316 585
R825 B.n315 B.n110 585
R826 B.n314 B.n313 585
R827 B.n312 B.n111 585
R828 B.n311 B.n310 585
R829 B.n309 B.n112 585
R830 B.n308 B.n307 585
R831 B.n306 B.n113 585
R832 B.n305 B.n304 585
R833 B.n303 B.n114 585
R834 B.n302 B.n301 585
R835 B.n300 B.n115 585
R836 B.n299 B.n298 585
R837 B.n297 B.n116 585
R838 B.n296 B.n295 585
R839 B.n294 B.n117 585
R840 B.n293 B.n292 585
R841 B.n291 B.n118 585
R842 B.n290 B.n289 585
R843 B.n288 B.n119 585
R844 B.n287 B.n286 585
R845 B.n285 B.n284 585
R846 B.n283 B.n123 585
R847 B.n282 B.n281 585
R848 B.n280 B.n124 585
R849 B.n279 B.n278 585
R850 B.n277 B.n125 585
R851 B.n276 B.n275 585
R852 B.n274 B.n126 585
R853 B.n273 B.n272 585
R854 B.n270 B.n127 585
R855 B.n269 B.n268 585
R856 B.n267 B.n130 585
R857 B.n266 B.n265 585
R858 B.n264 B.n131 585
R859 B.n263 B.n262 585
R860 B.n261 B.n132 585
R861 B.n260 B.n259 585
R862 B.n258 B.n133 585
R863 B.n257 B.n256 585
R864 B.n255 B.n134 585
R865 B.n254 B.n253 585
R866 B.n252 B.n135 585
R867 B.n251 B.n250 585
R868 B.n249 B.n136 585
R869 B.n248 B.n247 585
R870 B.n246 B.n137 585
R871 B.n245 B.n244 585
R872 B.n243 B.n138 585
R873 B.n242 B.n241 585
R874 B.n240 B.n139 585
R875 B.n239 B.n238 585
R876 B.n237 B.n140 585
R877 B.n236 B.n235 585
R878 B.n234 B.n141 585
R879 B.n233 B.n232 585
R880 B.n231 B.n142 585
R881 B.n230 B.n229 585
R882 B.n228 B.n143 585
R883 B.n227 B.n226 585
R884 B.n225 B.n144 585
R885 B.n224 B.n223 585
R886 B.n222 B.n145 585
R887 B.n221 B.n220 585
R888 B.n219 B.n146 585
R889 B.n218 B.n217 585
R890 B.n216 B.n147 585
R891 B.n215 B.n214 585
R892 B.n213 B.n148 585
R893 B.n212 B.n211 585
R894 B.n210 B.n149 585
R895 B.n209 B.n208 585
R896 B.n207 B.n150 585
R897 B.n206 B.n205 585
R898 B.n204 B.n151 585
R899 B.n203 B.n202 585
R900 B.n201 B.n152 585
R901 B.n200 B.n199 585
R902 B.n359 B.n358 585
R903 B.n360 B.n95 585
R904 B.n362 B.n361 585
R905 B.n363 B.n94 585
R906 B.n365 B.n364 585
R907 B.n366 B.n93 585
R908 B.n368 B.n367 585
R909 B.n369 B.n92 585
R910 B.n371 B.n370 585
R911 B.n372 B.n91 585
R912 B.n374 B.n373 585
R913 B.n375 B.n90 585
R914 B.n377 B.n376 585
R915 B.n378 B.n89 585
R916 B.n380 B.n379 585
R917 B.n381 B.n88 585
R918 B.n383 B.n382 585
R919 B.n384 B.n87 585
R920 B.n386 B.n385 585
R921 B.n387 B.n86 585
R922 B.n389 B.n388 585
R923 B.n390 B.n85 585
R924 B.n392 B.n391 585
R925 B.n393 B.n84 585
R926 B.n395 B.n394 585
R927 B.n396 B.n83 585
R928 B.n398 B.n397 585
R929 B.n399 B.n82 585
R930 B.n401 B.n400 585
R931 B.n402 B.n81 585
R932 B.n404 B.n403 585
R933 B.n405 B.n80 585
R934 B.n407 B.n406 585
R935 B.n408 B.n79 585
R936 B.n410 B.n409 585
R937 B.n411 B.n78 585
R938 B.n413 B.n412 585
R939 B.n414 B.n77 585
R940 B.n416 B.n415 585
R941 B.n417 B.n76 585
R942 B.n419 B.n418 585
R943 B.n420 B.n75 585
R944 B.n422 B.n421 585
R945 B.n423 B.n74 585
R946 B.n425 B.n424 585
R947 B.n426 B.n73 585
R948 B.n428 B.n427 585
R949 B.n429 B.n72 585
R950 B.n431 B.n430 585
R951 B.n432 B.n71 585
R952 B.n591 B.n14 585
R953 B.n590 B.n589 585
R954 B.n588 B.n15 585
R955 B.n587 B.n586 585
R956 B.n585 B.n16 585
R957 B.n584 B.n583 585
R958 B.n582 B.n17 585
R959 B.n581 B.n580 585
R960 B.n579 B.n18 585
R961 B.n578 B.n577 585
R962 B.n576 B.n19 585
R963 B.n575 B.n574 585
R964 B.n573 B.n20 585
R965 B.n572 B.n571 585
R966 B.n570 B.n21 585
R967 B.n569 B.n568 585
R968 B.n567 B.n22 585
R969 B.n566 B.n565 585
R970 B.n564 B.n23 585
R971 B.n563 B.n562 585
R972 B.n561 B.n24 585
R973 B.n560 B.n559 585
R974 B.n558 B.n25 585
R975 B.n557 B.n556 585
R976 B.n555 B.n26 585
R977 B.n554 B.n553 585
R978 B.n552 B.n27 585
R979 B.n551 B.n550 585
R980 B.n549 B.n28 585
R981 B.n548 B.n547 585
R982 B.n546 B.n29 585
R983 B.n545 B.n544 585
R984 B.n543 B.n30 585
R985 B.n542 B.n541 585
R986 B.n540 B.n31 585
R987 B.n539 B.n538 585
R988 B.n537 B.n32 585
R989 B.n536 B.n535 585
R990 B.n534 B.n33 585
R991 B.n533 B.n532 585
R992 B.n531 B.n34 585
R993 B.n530 B.n529 585
R994 B.n528 B.n35 585
R995 B.n527 B.n526 585
R996 B.n525 B.n36 585
R997 B.n524 B.n523 585
R998 B.n522 B.n37 585
R999 B.n521 B.n520 585
R1000 B.n519 B.n518 585
R1001 B.n517 B.n41 585
R1002 B.n516 B.n515 585
R1003 B.n514 B.n42 585
R1004 B.n513 B.n512 585
R1005 B.n511 B.n43 585
R1006 B.n510 B.n509 585
R1007 B.n508 B.n44 585
R1008 B.n507 B.n506 585
R1009 B.n504 B.n45 585
R1010 B.n503 B.n502 585
R1011 B.n501 B.n48 585
R1012 B.n500 B.n499 585
R1013 B.n498 B.n49 585
R1014 B.n497 B.n496 585
R1015 B.n495 B.n50 585
R1016 B.n494 B.n493 585
R1017 B.n492 B.n51 585
R1018 B.n491 B.n490 585
R1019 B.n489 B.n52 585
R1020 B.n488 B.n487 585
R1021 B.n486 B.n53 585
R1022 B.n485 B.n484 585
R1023 B.n483 B.n54 585
R1024 B.n482 B.n481 585
R1025 B.n480 B.n55 585
R1026 B.n479 B.n478 585
R1027 B.n477 B.n56 585
R1028 B.n476 B.n475 585
R1029 B.n474 B.n57 585
R1030 B.n473 B.n472 585
R1031 B.n471 B.n58 585
R1032 B.n470 B.n469 585
R1033 B.n468 B.n59 585
R1034 B.n467 B.n466 585
R1035 B.n465 B.n60 585
R1036 B.n464 B.n463 585
R1037 B.n462 B.n61 585
R1038 B.n461 B.n460 585
R1039 B.n459 B.n62 585
R1040 B.n458 B.n457 585
R1041 B.n456 B.n63 585
R1042 B.n455 B.n454 585
R1043 B.n453 B.n64 585
R1044 B.n452 B.n451 585
R1045 B.n450 B.n65 585
R1046 B.n449 B.n448 585
R1047 B.n447 B.n66 585
R1048 B.n446 B.n445 585
R1049 B.n444 B.n67 585
R1050 B.n443 B.n442 585
R1051 B.n441 B.n68 585
R1052 B.n440 B.n439 585
R1053 B.n438 B.n69 585
R1054 B.n437 B.n436 585
R1055 B.n435 B.n70 585
R1056 B.n434 B.n433 585
R1057 B.n593 B.n592 585
R1058 B.n594 B.n13 585
R1059 B.n596 B.n595 585
R1060 B.n597 B.n12 585
R1061 B.n599 B.n598 585
R1062 B.n600 B.n11 585
R1063 B.n602 B.n601 585
R1064 B.n603 B.n10 585
R1065 B.n605 B.n604 585
R1066 B.n606 B.n9 585
R1067 B.n608 B.n607 585
R1068 B.n609 B.n8 585
R1069 B.n611 B.n610 585
R1070 B.n612 B.n7 585
R1071 B.n614 B.n613 585
R1072 B.n615 B.n6 585
R1073 B.n617 B.n616 585
R1074 B.n618 B.n5 585
R1075 B.n620 B.n619 585
R1076 B.n621 B.n4 585
R1077 B.n623 B.n622 585
R1078 B.n624 B.n3 585
R1079 B.n626 B.n625 585
R1080 B.n627 B.n0 585
R1081 B.n2 B.n1 585
R1082 B.n165 B.n164 585
R1083 B.n167 B.n166 585
R1084 B.n168 B.n163 585
R1085 B.n170 B.n169 585
R1086 B.n171 B.n162 585
R1087 B.n173 B.n172 585
R1088 B.n174 B.n161 585
R1089 B.n176 B.n175 585
R1090 B.n177 B.n160 585
R1091 B.n179 B.n178 585
R1092 B.n180 B.n159 585
R1093 B.n182 B.n181 585
R1094 B.n183 B.n158 585
R1095 B.n185 B.n184 585
R1096 B.n186 B.n157 585
R1097 B.n188 B.n187 585
R1098 B.n189 B.n156 585
R1099 B.n191 B.n190 585
R1100 B.n192 B.n155 585
R1101 B.n194 B.n193 585
R1102 B.n195 B.n154 585
R1103 B.n197 B.n196 585
R1104 B.n198 B.n153 585
R1105 B.n200 B.n153 468.476
R1106 B.n358 B.n357 468.476
R1107 B.n434 B.n71 468.476
R1108 B.n592 B.n591 468.476
R1109 B.n120 B.t10 429.533
R1110 B.n46 B.t5 429.533
R1111 B.n128 B.t1 429.533
R1112 B.n38 B.t8 429.533
R1113 B.n121 B.t11 411.497
R1114 B.n47 B.t4 411.497
R1115 B.n129 B.t2 411.497
R1116 B.n39 B.t7 411.497
R1117 B.n629 B.n628 256.663
R1118 B.n628 B.n627 235.042
R1119 B.n628 B.n2 235.042
R1120 B.n201 B.n200 163.367
R1121 B.n202 B.n201 163.367
R1122 B.n202 B.n151 163.367
R1123 B.n206 B.n151 163.367
R1124 B.n207 B.n206 163.367
R1125 B.n208 B.n207 163.367
R1126 B.n208 B.n149 163.367
R1127 B.n212 B.n149 163.367
R1128 B.n213 B.n212 163.367
R1129 B.n214 B.n213 163.367
R1130 B.n214 B.n147 163.367
R1131 B.n218 B.n147 163.367
R1132 B.n219 B.n218 163.367
R1133 B.n220 B.n219 163.367
R1134 B.n220 B.n145 163.367
R1135 B.n224 B.n145 163.367
R1136 B.n225 B.n224 163.367
R1137 B.n226 B.n225 163.367
R1138 B.n226 B.n143 163.367
R1139 B.n230 B.n143 163.367
R1140 B.n231 B.n230 163.367
R1141 B.n232 B.n231 163.367
R1142 B.n232 B.n141 163.367
R1143 B.n236 B.n141 163.367
R1144 B.n237 B.n236 163.367
R1145 B.n238 B.n237 163.367
R1146 B.n238 B.n139 163.367
R1147 B.n242 B.n139 163.367
R1148 B.n243 B.n242 163.367
R1149 B.n244 B.n243 163.367
R1150 B.n244 B.n137 163.367
R1151 B.n248 B.n137 163.367
R1152 B.n249 B.n248 163.367
R1153 B.n250 B.n249 163.367
R1154 B.n250 B.n135 163.367
R1155 B.n254 B.n135 163.367
R1156 B.n255 B.n254 163.367
R1157 B.n256 B.n255 163.367
R1158 B.n256 B.n133 163.367
R1159 B.n260 B.n133 163.367
R1160 B.n261 B.n260 163.367
R1161 B.n262 B.n261 163.367
R1162 B.n262 B.n131 163.367
R1163 B.n266 B.n131 163.367
R1164 B.n267 B.n266 163.367
R1165 B.n268 B.n267 163.367
R1166 B.n268 B.n127 163.367
R1167 B.n273 B.n127 163.367
R1168 B.n274 B.n273 163.367
R1169 B.n275 B.n274 163.367
R1170 B.n275 B.n125 163.367
R1171 B.n279 B.n125 163.367
R1172 B.n280 B.n279 163.367
R1173 B.n281 B.n280 163.367
R1174 B.n281 B.n123 163.367
R1175 B.n285 B.n123 163.367
R1176 B.n286 B.n285 163.367
R1177 B.n286 B.n119 163.367
R1178 B.n290 B.n119 163.367
R1179 B.n291 B.n290 163.367
R1180 B.n292 B.n291 163.367
R1181 B.n292 B.n117 163.367
R1182 B.n296 B.n117 163.367
R1183 B.n297 B.n296 163.367
R1184 B.n298 B.n297 163.367
R1185 B.n298 B.n115 163.367
R1186 B.n302 B.n115 163.367
R1187 B.n303 B.n302 163.367
R1188 B.n304 B.n303 163.367
R1189 B.n304 B.n113 163.367
R1190 B.n308 B.n113 163.367
R1191 B.n309 B.n308 163.367
R1192 B.n310 B.n309 163.367
R1193 B.n310 B.n111 163.367
R1194 B.n314 B.n111 163.367
R1195 B.n315 B.n314 163.367
R1196 B.n316 B.n315 163.367
R1197 B.n316 B.n109 163.367
R1198 B.n320 B.n109 163.367
R1199 B.n321 B.n320 163.367
R1200 B.n322 B.n321 163.367
R1201 B.n322 B.n107 163.367
R1202 B.n326 B.n107 163.367
R1203 B.n327 B.n326 163.367
R1204 B.n328 B.n327 163.367
R1205 B.n328 B.n105 163.367
R1206 B.n332 B.n105 163.367
R1207 B.n333 B.n332 163.367
R1208 B.n334 B.n333 163.367
R1209 B.n334 B.n103 163.367
R1210 B.n338 B.n103 163.367
R1211 B.n339 B.n338 163.367
R1212 B.n340 B.n339 163.367
R1213 B.n340 B.n101 163.367
R1214 B.n344 B.n101 163.367
R1215 B.n345 B.n344 163.367
R1216 B.n346 B.n345 163.367
R1217 B.n346 B.n99 163.367
R1218 B.n350 B.n99 163.367
R1219 B.n351 B.n350 163.367
R1220 B.n352 B.n351 163.367
R1221 B.n352 B.n97 163.367
R1222 B.n356 B.n97 163.367
R1223 B.n357 B.n356 163.367
R1224 B.n430 B.n71 163.367
R1225 B.n430 B.n429 163.367
R1226 B.n429 B.n428 163.367
R1227 B.n428 B.n73 163.367
R1228 B.n424 B.n73 163.367
R1229 B.n424 B.n423 163.367
R1230 B.n423 B.n422 163.367
R1231 B.n422 B.n75 163.367
R1232 B.n418 B.n75 163.367
R1233 B.n418 B.n417 163.367
R1234 B.n417 B.n416 163.367
R1235 B.n416 B.n77 163.367
R1236 B.n412 B.n77 163.367
R1237 B.n412 B.n411 163.367
R1238 B.n411 B.n410 163.367
R1239 B.n410 B.n79 163.367
R1240 B.n406 B.n79 163.367
R1241 B.n406 B.n405 163.367
R1242 B.n405 B.n404 163.367
R1243 B.n404 B.n81 163.367
R1244 B.n400 B.n81 163.367
R1245 B.n400 B.n399 163.367
R1246 B.n399 B.n398 163.367
R1247 B.n398 B.n83 163.367
R1248 B.n394 B.n83 163.367
R1249 B.n394 B.n393 163.367
R1250 B.n393 B.n392 163.367
R1251 B.n392 B.n85 163.367
R1252 B.n388 B.n85 163.367
R1253 B.n388 B.n387 163.367
R1254 B.n387 B.n386 163.367
R1255 B.n386 B.n87 163.367
R1256 B.n382 B.n87 163.367
R1257 B.n382 B.n381 163.367
R1258 B.n381 B.n380 163.367
R1259 B.n380 B.n89 163.367
R1260 B.n376 B.n89 163.367
R1261 B.n376 B.n375 163.367
R1262 B.n375 B.n374 163.367
R1263 B.n374 B.n91 163.367
R1264 B.n370 B.n91 163.367
R1265 B.n370 B.n369 163.367
R1266 B.n369 B.n368 163.367
R1267 B.n368 B.n93 163.367
R1268 B.n364 B.n93 163.367
R1269 B.n364 B.n363 163.367
R1270 B.n363 B.n362 163.367
R1271 B.n362 B.n95 163.367
R1272 B.n358 B.n95 163.367
R1273 B.n591 B.n590 163.367
R1274 B.n590 B.n15 163.367
R1275 B.n586 B.n15 163.367
R1276 B.n586 B.n585 163.367
R1277 B.n585 B.n584 163.367
R1278 B.n584 B.n17 163.367
R1279 B.n580 B.n17 163.367
R1280 B.n580 B.n579 163.367
R1281 B.n579 B.n578 163.367
R1282 B.n578 B.n19 163.367
R1283 B.n574 B.n19 163.367
R1284 B.n574 B.n573 163.367
R1285 B.n573 B.n572 163.367
R1286 B.n572 B.n21 163.367
R1287 B.n568 B.n21 163.367
R1288 B.n568 B.n567 163.367
R1289 B.n567 B.n566 163.367
R1290 B.n566 B.n23 163.367
R1291 B.n562 B.n23 163.367
R1292 B.n562 B.n561 163.367
R1293 B.n561 B.n560 163.367
R1294 B.n560 B.n25 163.367
R1295 B.n556 B.n25 163.367
R1296 B.n556 B.n555 163.367
R1297 B.n555 B.n554 163.367
R1298 B.n554 B.n27 163.367
R1299 B.n550 B.n27 163.367
R1300 B.n550 B.n549 163.367
R1301 B.n549 B.n548 163.367
R1302 B.n548 B.n29 163.367
R1303 B.n544 B.n29 163.367
R1304 B.n544 B.n543 163.367
R1305 B.n543 B.n542 163.367
R1306 B.n542 B.n31 163.367
R1307 B.n538 B.n31 163.367
R1308 B.n538 B.n537 163.367
R1309 B.n537 B.n536 163.367
R1310 B.n536 B.n33 163.367
R1311 B.n532 B.n33 163.367
R1312 B.n532 B.n531 163.367
R1313 B.n531 B.n530 163.367
R1314 B.n530 B.n35 163.367
R1315 B.n526 B.n35 163.367
R1316 B.n526 B.n525 163.367
R1317 B.n525 B.n524 163.367
R1318 B.n524 B.n37 163.367
R1319 B.n520 B.n37 163.367
R1320 B.n520 B.n519 163.367
R1321 B.n519 B.n41 163.367
R1322 B.n515 B.n41 163.367
R1323 B.n515 B.n514 163.367
R1324 B.n514 B.n513 163.367
R1325 B.n513 B.n43 163.367
R1326 B.n509 B.n43 163.367
R1327 B.n509 B.n508 163.367
R1328 B.n508 B.n507 163.367
R1329 B.n507 B.n45 163.367
R1330 B.n502 B.n45 163.367
R1331 B.n502 B.n501 163.367
R1332 B.n501 B.n500 163.367
R1333 B.n500 B.n49 163.367
R1334 B.n496 B.n49 163.367
R1335 B.n496 B.n495 163.367
R1336 B.n495 B.n494 163.367
R1337 B.n494 B.n51 163.367
R1338 B.n490 B.n51 163.367
R1339 B.n490 B.n489 163.367
R1340 B.n489 B.n488 163.367
R1341 B.n488 B.n53 163.367
R1342 B.n484 B.n53 163.367
R1343 B.n484 B.n483 163.367
R1344 B.n483 B.n482 163.367
R1345 B.n482 B.n55 163.367
R1346 B.n478 B.n55 163.367
R1347 B.n478 B.n477 163.367
R1348 B.n477 B.n476 163.367
R1349 B.n476 B.n57 163.367
R1350 B.n472 B.n57 163.367
R1351 B.n472 B.n471 163.367
R1352 B.n471 B.n470 163.367
R1353 B.n470 B.n59 163.367
R1354 B.n466 B.n59 163.367
R1355 B.n466 B.n465 163.367
R1356 B.n465 B.n464 163.367
R1357 B.n464 B.n61 163.367
R1358 B.n460 B.n61 163.367
R1359 B.n460 B.n459 163.367
R1360 B.n459 B.n458 163.367
R1361 B.n458 B.n63 163.367
R1362 B.n454 B.n63 163.367
R1363 B.n454 B.n453 163.367
R1364 B.n453 B.n452 163.367
R1365 B.n452 B.n65 163.367
R1366 B.n448 B.n65 163.367
R1367 B.n448 B.n447 163.367
R1368 B.n447 B.n446 163.367
R1369 B.n446 B.n67 163.367
R1370 B.n442 B.n67 163.367
R1371 B.n442 B.n441 163.367
R1372 B.n441 B.n440 163.367
R1373 B.n440 B.n69 163.367
R1374 B.n436 B.n69 163.367
R1375 B.n436 B.n435 163.367
R1376 B.n435 B.n434 163.367
R1377 B.n592 B.n13 163.367
R1378 B.n596 B.n13 163.367
R1379 B.n597 B.n596 163.367
R1380 B.n598 B.n597 163.367
R1381 B.n598 B.n11 163.367
R1382 B.n602 B.n11 163.367
R1383 B.n603 B.n602 163.367
R1384 B.n604 B.n603 163.367
R1385 B.n604 B.n9 163.367
R1386 B.n608 B.n9 163.367
R1387 B.n609 B.n608 163.367
R1388 B.n610 B.n609 163.367
R1389 B.n610 B.n7 163.367
R1390 B.n614 B.n7 163.367
R1391 B.n615 B.n614 163.367
R1392 B.n616 B.n615 163.367
R1393 B.n616 B.n5 163.367
R1394 B.n620 B.n5 163.367
R1395 B.n621 B.n620 163.367
R1396 B.n622 B.n621 163.367
R1397 B.n622 B.n3 163.367
R1398 B.n626 B.n3 163.367
R1399 B.n627 B.n626 163.367
R1400 B.n165 B.n2 163.367
R1401 B.n166 B.n165 163.367
R1402 B.n166 B.n163 163.367
R1403 B.n170 B.n163 163.367
R1404 B.n171 B.n170 163.367
R1405 B.n172 B.n171 163.367
R1406 B.n172 B.n161 163.367
R1407 B.n176 B.n161 163.367
R1408 B.n177 B.n176 163.367
R1409 B.n178 B.n177 163.367
R1410 B.n178 B.n159 163.367
R1411 B.n182 B.n159 163.367
R1412 B.n183 B.n182 163.367
R1413 B.n184 B.n183 163.367
R1414 B.n184 B.n157 163.367
R1415 B.n188 B.n157 163.367
R1416 B.n189 B.n188 163.367
R1417 B.n190 B.n189 163.367
R1418 B.n190 B.n155 163.367
R1419 B.n194 B.n155 163.367
R1420 B.n195 B.n194 163.367
R1421 B.n196 B.n195 163.367
R1422 B.n196 B.n153 163.367
R1423 B.n271 B.n129 59.5399
R1424 B.n122 B.n121 59.5399
R1425 B.n505 B.n47 59.5399
R1426 B.n40 B.n39 59.5399
R1427 B.n359 B.n96 30.4395
R1428 B.n593 B.n14 30.4395
R1429 B.n433 B.n432 30.4395
R1430 B.n199 B.n198 30.4395
R1431 B B.n629 18.0485
R1432 B.n129 B.n128 18.0369
R1433 B.n121 B.n120 18.0369
R1434 B.n47 B.n46 18.0369
R1435 B.n39 B.n38 18.0369
R1436 B.n594 B.n593 10.6151
R1437 B.n595 B.n594 10.6151
R1438 B.n595 B.n12 10.6151
R1439 B.n599 B.n12 10.6151
R1440 B.n600 B.n599 10.6151
R1441 B.n601 B.n600 10.6151
R1442 B.n601 B.n10 10.6151
R1443 B.n605 B.n10 10.6151
R1444 B.n606 B.n605 10.6151
R1445 B.n607 B.n606 10.6151
R1446 B.n607 B.n8 10.6151
R1447 B.n611 B.n8 10.6151
R1448 B.n612 B.n611 10.6151
R1449 B.n613 B.n612 10.6151
R1450 B.n613 B.n6 10.6151
R1451 B.n617 B.n6 10.6151
R1452 B.n618 B.n617 10.6151
R1453 B.n619 B.n618 10.6151
R1454 B.n619 B.n4 10.6151
R1455 B.n623 B.n4 10.6151
R1456 B.n624 B.n623 10.6151
R1457 B.n625 B.n624 10.6151
R1458 B.n625 B.n0 10.6151
R1459 B.n589 B.n14 10.6151
R1460 B.n589 B.n588 10.6151
R1461 B.n588 B.n587 10.6151
R1462 B.n587 B.n16 10.6151
R1463 B.n583 B.n16 10.6151
R1464 B.n583 B.n582 10.6151
R1465 B.n582 B.n581 10.6151
R1466 B.n581 B.n18 10.6151
R1467 B.n577 B.n18 10.6151
R1468 B.n577 B.n576 10.6151
R1469 B.n576 B.n575 10.6151
R1470 B.n575 B.n20 10.6151
R1471 B.n571 B.n20 10.6151
R1472 B.n571 B.n570 10.6151
R1473 B.n570 B.n569 10.6151
R1474 B.n569 B.n22 10.6151
R1475 B.n565 B.n22 10.6151
R1476 B.n565 B.n564 10.6151
R1477 B.n564 B.n563 10.6151
R1478 B.n563 B.n24 10.6151
R1479 B.n559 B.n24 10.6151
R1480 B.n559 B.n558 10.6151
R1481 B.n558 B.n557 10.6151
R1482 B.n557 B.n26 10.6151
R1483 B.n553 B.n26 10.6151
R1484 B.n553 B.n552 10.6151
R1485 B.n552 B.n551 10.6151
R1486 B.n551 B.n28 10.6151
R1487 B.n547 B.n28 10.6151
R1488 B.n547 B.n546 10.6151
R1489 B.n546 B.n545 10.6151
R1490 B.n545 B.n30 10.6151
R1491 B.n541 B.n30 10.6151
R1492 B.n541 B.n540 10.6151
R1493 B.n540 B.n539 10.6151
R1494 B.n539 B.n32 10.6151
R1495 B.n535 B.n32 10.6151
R1496 B.n535 B.n534 10.6151
R1497 B.n534 B.n533 10.6151
R1498 B.n533 B.n34 10.6151
R1499 B.n529 B.n34 10.6151
R1500 B.n529 B.n528 10.6151
R1501 B.n528 B.n527 10.6151
R1502 B.n527 B.n36 10.6151
R1503 B.n523 B.n36 10.6151
R1504 B.n523 B.n522 10.6151
R1505 B.n522 B.n521 10.6151
R1506 B.n518 B.n517 10.6151
R1507 B.n517 B.n516 10.6151
R1508 B.n516 B.n42 10.6151
R1509 B.n512 B.n42 10.6151
R1510 B.n512 B.n511 10.6151
R1511 B.n511 B.n510 10.6151
R1512 B.n510 B.n44 10.6151
R1513 B.n506 B.n44 10.6151
R1514 B.n504 B.n503 10.6151
R1515 B.n503 B.n48 10.6151
R1516 B.n499 B.n48 10.6151
R1517 B.n499 B.n498 10.6151
R1518 B.n498 B.n497 10.6151
R1519 B.n497 B.n50 10.6151
R1520 B.n493 B.n50 10.6151
R1521 B.n493 B.n492 10.6151
R1522 B.n492 B.n491 10.6151
R1523 B.n491 B.n52 10.6151
R1524 B.n487 B.n52 10.6151
R1525 B.n487 B.n486 10.6151
R1526 B.n486 B.n485 10.6151
R1527 B.n485 B.n54 10.6151
R1528 B.n481 B.n54 10.6151
R1529 B.n481 B.n480 10.6151
R1530 B.n480 B.n479 10.6151
R1531 B.n479 B.n56 10.6151
R1532 B.n475 B.n56 10.6151
R1533 B.n475 B.n474 10.6151
R1534 B.n474 B.n473 10.6151
R1535 B.n473 B.n58 10.6151
R1536 B.n469 B.n58 10.6151
R1537 B.n469 B.n468 10.6151
R1538 B.n468 B.n467 10.6151
R1539 B.n467 B.n60 10.6151
R1540 B.n463 B.n60 10.6151
R1541 B.n463 B.n462 10.6151
R1542 B.n462 B.n461 10.6151
R1543 B.n461 B.n62 10.6151
R1544 B.n457 B.n62 10.6151
R1545 B.n457 B.n456 10.6151
R1546 B.n456 B.n455 10.6151
R1547 B.n455 B.n64 10.6151
R1548 B.n451 B.n64 10.6151
R1549 B.n451 B.n450 10.6151
R1550 B.n450 B.n449 10.6151
R1551 B.n449 B.n66 10.6151
R1552 B.n445 B.n66 10.6151
R1553 B.n445 B.n444 10.6151
R1554 B.n444 B.n443 10.6151
R1555 B.n443 B.n68 10.6151
R1556 B.n439 B.n68 10.6151
R1557 B.n439 B.n438 10.6151
R1558 B.n438 B.n437 10.6151
R1559 B.n437 B.n70 10.6151
R1560 B.n433 B.n70 10.6151
R1561 B.n432 B.n431 10.6151
R1562 B.n431 B.n72 10.6151
R1563 B.n427 B.n72 10.6151
R1564 B.n427 B.n426 10.6151
R1565 B.n426 B.n425 10.6151
R1566 B.n425 B.n74 10.6151
R1567 B.n421 B.n74 10.6151
R1568 B.n421 B.n420 10.6151
R1569 B.n420 B.n419 10.6151
R1570 B.n419 B.n76 10.6151
R1571 B.n415 B.n76 10.6151
R1572 B.n415 B.n414 10.6151
R1573 B.n414 B.n413 10.6151
R1574 B.n413 B.n78 10.6151
R1575 B.n409 B.n78 10.6151
R1576 B.n409 B.n408 10.6151
R1577 B.n408 B.n407 10.6151
R1578 B.n407 B.n80 10.6151
R1579 B.n403 B.n80 10.6151
R1580 B.n403 B.n402 10.6151
R1581 B.n402 B.n401 10.6151
R1582 B.n401 B.n82 10.6151
R1583 B.n397 B.n82 10.6151
R1584 B.n397 B.n396 10.6151
R1585 B.n396 B.n395 10.6151
R1586 B.n395 B.n84 10.6151
R1587 B.n391 B.n84 10.6151
R1588 B.n391 B.n390 10.6151
R1589 B.n390 B.n389 10.6151
R1590 B.n389 B.n86 10.6151
R1591 B.n385 B.n86 10.6151
R1592 B.n385 B.n384 10.6151
R1593 B.n384 B.n383 10.6151
R1594 B.n383 B.n88 10.6151
R1595 B.n379 B.n88 10.6151
R1596 B.n379 B.n378 10.6151
R1597 B.n378 B.n377 10.6151
R1598 B.n377 B.n90 10.6151
R1599 B.n373 B.n90 10.6151
R1600 B.n373 B.n372 10.6151
R1601 B.n372 B.n371 10.6151
R1602 B.n371 B.n92 10.6151
R1603 B.n367 B.n92 10.6151
R1604 B.n367 B.n366 10.6151
R1605 B.n366 B.n365 10.6151
R1606 B.n365 B.n94 10.6151
R1607 B.n361 B.n94 10.6151
R1608 B.n361 B.n360 10.6151
R1609 B.n360 B.n359 10.6151
R1610 B.n164 B.n1 10.6151
R1611 B.n167 B.n164 10.6151
R1612 B.n168 B.n167 10.6151
R1613 B.n169 B.n168 10.6151
R1614 B.n169 B.n162 10.6151
R1615 B.n173 B.n162 10.6151
R1616 B.n174 B.n173 10.6151
R1617 B.n175 B.n174 10.6151
R1618 B.n175 B.n160 10.6151
R1619 B.n179 B.n160 10.6151
R1620 B.n180 B.n179 10.6151
R1621 B.n181 B.n180 10.6151
R1622 B.n181 B.n158 10.6151
R1623 B.n185 B.n158 10.6151
R1624 B.n186 B.n185 10.6151
R1625 B.n187 B.n186 10.6151
R1626 B.n187 B.n156 10.6151
R1627 B.n191 B.n156 10.6151
R1628 B.n192 B.n191 10.6151
R1629 B.n193 B.n192 10.6151
R1630 B.n193 B.n154 10.6151
R1631 B.n197 B.n154 10.6151
R1632 B.n198 B.n197 10.6151
R1633 B.n199 B.n152 10.6151
R1634 B.n203 B.n152 10.6151
R1635 B.n204 B.n203 10.6151
R1636 B.n205 B.n204 10.6151
R1637 B.n205 B.n150 10.6151
R1638 B.n209 B.n150 10.6151
R1639 B.n210 B.n209 10.6151
R1640 B.n211 B.n210 10.6151
R1641 B.n211 B.n148 10.6151
R1642 B.n215 B.n148 10.6151
R1643 B.n216 B.n215 10.6151
R1644 B.n217 B.n216 10.6151
R1645 B.n217 B.n146 10.6151
R1646 B.n221 B.n146 10.6151
R1647 B.n222 B.n221 10.6151
R1648 B.n223 B.n222 10.6151
R1649 B.n223 B.n144 10.6151
R1650 B.n227 B.n144 10.6151
R1651 B.n228 B.n227 10.6151
R1652 B.n229 B.n228 10.6151
R1653 B.n229 B.n142 10.6151
R1654 B.n233 B.n142 10.6151
R1655 B.n234 B.n233 10.6151
R1656 B.n235 B.n234 10.6151
R1657 B.n235 B.n140 10.6151
R1658 B.n239 B.n140 10.6151
R1659 B.n240 B.n239 10.6151
R1660 B.n241 B.n240 10.6151
R1661 B.n241 B.n138 10.6151
R1662 B.n245 B.n138 10.6151
R1663 B.n246 B.n245 10.6151
R1664 B.n247 B.n246 10.6151
R1665 B.n247 B.n136 10.6151
R1666 B.n251 B.n136 10.6151
R1667 B.n252 B.n251 10.6151
R1668 B.n253 B.n252 10.6151
R1669 B.n253 B.n134 10.6151
R1670 B.n257 B.n134 10.6151
R1671 B.n258 B.n257 10.6151
R1672 B.n259 B.n258 10.6151
R1673 B.n259 B.n132 10.6151
R1674 B.n263 B.n132 10.6151
R1675 B.n264 B.n263 10.6151
R1676 B.n265 B.n264 10.6151
R1677 B.n265 B.n130 10.6151
R1678 B.n269 B.n130 10.6151
R1679 B.n270 B.n269 10.6151
R1680 B.n272 B.n126 10.6151
R1681 B.n276 B.n126 10.6151
R1682 B.n277 B.n276 10.6151
R1683 B.n278 B.n277 10.6151
R1684 B.n278 B.n124 10.6151
R1685 B.n282 B.n124 10.6151
R1686 B.n283 B.n282 10.6151
R1687 B.n284 B.n283 10.6151
R1688 B.n288 B.n287 10.6151
R1689 B.n289 B.n288 10.6151
R1690 B.n289 B.n118 10.6151
R1691 B.n293 B.n118 10.6151
R1692 B.n294 B.n293 10.6151
R1693 B.n295 B.n294 10.6151
R1694 B.n295 B.n116 10.6151
R1695 B.n299 B.n116 10.6151
R1696 B.n300 B.n299 10.6151
R1697 B.n301 B.n300 10.6151
R1698 B.n301 B.n114 10.6151
R1699 B.n305 B.n114 10.6151
R1700 B.n306 B.n305 10.6151
R1701 B.n307 B.n306 10.6151
R1702 B.n307 B.n112 10.6151
R1703 B.n311 B.n112 10.6151
R1704 B.n312 B.n311 10.6151
R1705 B.n313 B.n312 10.6151
R1706 B.n313 B.n110 10.6151
R1707 B.n317 B.n110 10.6151
R1708 B.n318 B.n317 10.6151
R1709 B.n319 B.n318 10.6151
R1710 B.n319 B.n108 10.6151
R1711 B.n323 B.n108 10.6151
R1712 B.n324 B.n323 10.6151
R1713 B.n325 B.n324 10.6151
R1714 B.n325 B.n106 10.6151
R1715 B.n329 B.n106 10.6151
R1716 B.n330 B.n329 10.6151
R1717 B.n331 B.n330 10.6151
R1718 B.n331 B.n104 10.6151
R1719 B.n335 B.n104 10.6151
R1720 B.n336 B.n335 10.6151
R1721 B.n337 B.n336 10.6151
R1722 B.n337 B.n102 10.6151
R1723 B.n341 B.n102 10.6151
R1724 B.n342 B.n341 10.6151
R1725 B.n343 B.n342 10.6151
R1726 B.n343 B.n100 10.6151
R1727 B.n347 B.n100 10.6151
R1728 B.n348 B.n347 10.6151
R1729 B.n349 B.n348 10.6151
R1730 B.n349 B.n98 10.6151
R1731 B.n353 B.n98 10.6151
R1732 B.n354 B.n353 10.6151
R1733 B.n355 B.n354 10.6151
R1734 B.n355 B.n96 10.6151
R1735 B.n629 B.n0 8.11757
R1736 B.n629 B.n1 8.11757
R1737 B.n518 B.n40 6.5566
R1738 B.n506 B.n505 6.5566
R1739 B.n272 B.n271 6.5566
R1740 B.n284 B.n122 6.5566
R1741 B.n521 B.n40 4.05904
R1742 B.n505 B.n504 4.05904
R1743 B.n271 B.n270 4.05904
R1744 B.n287 B.n122 4.05904
R1745 VP.n6 VP.t6 654.006
R1746 VP.n14 VP.t8 627.806
R1747 VP.n16 VP.t7 627.806
R1748 VP.n1 VP.t0 627.806
R1749 VP.n20 VP.t9 627.806
R1750 VP.n22 VP.t5 627.806
R1751 VP.n11 VP.t1 627.806
R1752 VP.n9 VP.t2 627.806
R1753 VP.n8 VP.t3 627.806
R1754 VP.n7 VP.t4 627.806
R1755 VP.n23 VP.n22 161.3
R1756 VP.n9 VP.n4 161.3
R1757 VP.n10 VP.n3 161.3
R1758 VP.n12 VP.n11 161.3
R1759 VP.n21 VP.n0 161.3
R1760 VP.n20 VP.n19 161.3
R1761 VP.n17 VP.n16 161.3
R1762 VP.n15 VP.n2 161.3
R1763 VP.n14 VP.n13 161.3
R1764 VP.n8 VP.n5 80.6037
R1765 VP.n18 VP.n1 80.6037
R1766 VP.n16 VP.n1 48.2005
R1767 VP.n20 VP.n1 48.2005
R1768 VP.n9 VP.n8 48.2005
R1769 VP.n8 VP.n7 48.2005
R1770 VP.n15 VP.n14 45.2793
R1771 VP.n22 VP.n21 45.2793
R1772 VP.n11 VP.n10 45.2793
R1773 VP.n6 VP.n5 45.1669
R1774 VP.n13 VP.n12 43.7694
R1775 VP.n7 VP.n6 14.3992
R1776 VP.n16 VP.n15 2.92171
R1777 VP.n21 VP.n20 2.92171
R1778 VP.n10 VP.n9 2.92171
R1779 VP.n5 VP.n4 0.285035
R1780 VP.n18 VP.n17 0.285035
R1781 VP.n19 VP.n18 0.285035
R1782 VP.n4 VP.n3 0.189894
R1783 VP.n12 VP.n3 0.189894
R1784 VP.n13 VP.n2 0.189894
R1785 VP.n17 VP.n2 0.189894
R1786 VP.n19 VP.n0 0.189894
R1787 VP.n23 VP.n0 0.189894
R1788 VP VP.n23 0.0516364
R1789 VDD1.n72 VDD1.n0 756.745
R1790 VDD1.n151 VDD1.n79 756.745
R1791 VDD1.n73 VDD1.n72 585
R1792 VDD1.n71 VDD1.n2 585
R1793 VDD1.n70 VDD1.n69 585
R1794 VDD1.n5 VDD1.n3 585
R1795 VDD1.n64 VDD1.n63 585
R1796 VDD1.n62 VDD1.n61 585
R1797 VDD1.n9 VDD1.n8 585
R1798 VDD1.n56 VDD1.n55 585
R1799 VDD1.n54 VDD1.n53 585
R1800 VDD1.n13 VDD1.n12 585
R1801 VDD1.n48 VDD1.n47 585
R1802 VDD1.n46 VDD1.n45 585
R1803 VDD1.n17 VDD1.n16 585
R1804 VDD1.n40 VDD1.n39 585
R1805 VDD1.n38 VDD1.n37 585
R1806 VDD1.n21 VDD1.n20 585
R1807 VDD1.n32 VDD1.n31 585
R1808 VDD1.n30 VDD1.n29 585
R1809 VDD1.n25 VDD1.n24 585
R1810 VDD1.n103 VDD1.n102 585
R1811 VDD1.n108 VDD1.n107 585
R1812 VDD1.n110 VDD1.n109 585
R1813 VDD1.n99 VDD1.n98 585
R1814 VDD1.n116 VDD1.n115 585
R1815 VDD1.n118 VDD1.n117 585
R1816 VDD1.n95 VDD1.n94 585
R1817 VDD1.n124 VDD1.n123 585
R1818 VDD1.n126 VDD1.n125 585
R1819 VDD1.n91 VDD1.n90 585
R1820 VDD1.n132 VDD1.n131 585
R1821 VDD1.n134 VDD1.n133 585
R1822 VDD1.n87 VDD1.n86 585
R1823 VDD1.n140 VDD1.n139 585
R1824 VDD1.n142 VDD1.n141 585
R1825 VDD1.n83 VDD1.n82 585
R1826 VDD1.n149 VDD1.n148 585
R1827 VDD1.n150 VDD1.n81 585
R1828 VDD1.n152 VDD1.n151 585
R1829 VDD1.n26 VDD1.t3 327.466
R1830 VDD1.n104 VDD1.t1 327.466
R1831 VDD1.n72 VDD1.n71 171.744
R1832 VDD1.n71 VDD1.n70 171.744
R1833 VDD1.n70 VDD1.n3 171.744
R1834 VDD1.n63 VDD1.n3 171.744
R1835 VDD1.n63 VDD1.n62 171.744
R1836 VDD1.n62 VDD1.n8 171.744
R1837 VDD1.n55 VDD1.n8 171.744
R1838 VDD1.n55 VDD1.n54 171.744
R1839 VDD1.n54 VDD1.n12 171.744
R1840 VDD1.n47 VDD1.n12 171.744
R1841 VDD1.n47 VDD1.n46 171.744
R1842 VDD1.n46 VDD1.n16 171.744
R1843 VDD1.n39 VDD1.n16 171.744
R1844 VDD1.n39 VDD1.n38 171.744
R1845 VDD1.n38 VDD1.n20 171.744
R1846 VDD1.n31 VDD1.n20 171.744
R1847 VDD1.n31 VDD1.n30 171.744
R1848 VDD1.n30 VDD1.n24 171.744
R1849 VDD1.n108 VDD1.n102 171.744
R1850 VDD1.n109 VDD1.n108 171.744
R1851 VDD1.n109 VDD1.n98 171.744
R1852 VDD1.n116 VDD1.n98 171.744
R1853 VDD1.n117 VDD1.n116 171.744
R1854 VDD1.n117 VDD1.n94 171.744
R1855 VDD1.n124 VDD1.n94 171.744
R1856 VDD1.n125 VDD1.n124 171.744
R1857 VDD1.n125 VDD1.n90 171.744
R1858 VDD1.n132 VDD1.n90 171.744
R1859 VDD1.n133 VDD1.n132 171.744
R1860 VDD1.n133 VDD1.n86 171.744
R1861 VDD1.n140 VDD1.n86 171.744
R1862 VDD1.n141 VDD1.n140 171.744
R1863 VDD1.n141 VDD1.n82 171.744
R1864 VDD1.n149 VDD1.n82 171.744
R1865 VDD1.n150 VDD1.n149 171.744
R1866 VDD1.n151 VDD1.n150 171.744
R1867 VDD1.t3 VDD1.n24 85.8723
R1868 VDD1.t1 VDD1.n102 85.8723
R1869 VDD1.n159 VDD1.n158 73.4316
R1870 VDD1.n78 VDD1.n77 72.8858
R1871 VDD1.n161 VDD1.n160 72.8856
R1872 VDD1.n157 VDD1.n156 72.8856
R1873 VDD1.n78 VDD1.n76 51.2174
R1874 VDD1.n157 VDD1.n155 51.2174
R1875 VDD1.n161 VDD1.n159 40.5763
R1876 VDD1.n26 VDD1.n25 16.3895
R1877 VDD1.n104 VDD1.n103 16.3895
R1878 VDD1.n73 VDD1.n2 13.1884
R1879 VDD1.n152 VDD1.n81 13.1884
R1880 VDD1.n74 VDD1.n0 12.8005
R1881 VDD1.n69 VDD1.n4 12.8005
R1882 VDD1.n29 VDD1.n28 12.8005
R1883 VDD1.n107 VDD1.n106 12.8005
R1884 VDD1.n148 VDD1.n147 12.8005
R1885 VDD1.n153 VDD1.n79 12.8005
R1886 VDD1.n68 VDD1.n5 12.0247
R1887 VDD1.n32 VDD1.n23 12.0247
R1888 VDD1.n110 VDD1.n101 12.0247
R1889 VDD1.n146 VDD1.n83 12.0247
R1890 VDD1.n65 VDD1.n64 11.249
R1891 VDD1.n33 VDD1.n21 11.249
R1892 VDD1.n111 VDD1.n99 11.249
R1893 VDD1.n143 VDD1.n142 11.249
R1894 VDD1.n61 VDD1.n7 10.4732
R1895 VDD1.n37 VDD1.n36 10.4732
R1896 VDD1.n115 VDD1.n114 10.4732
R1897 VDD1.n139 VDD1.n85 10.4732
R1898 VDD1.n60 VDD1.n9 9.69747
R1899 VDD1.n40 VDD1.n19 9.69747
R1900 VDD1.n118 VDD1.n97 9.69747
R1901 VDD1.n138 VDD1.n87 9.69747
R1902 VDD1.n76 VDD1.n75 9.45567
R1903 VDD1.n155 VDD1.n154 9.45567
R1904 VDD1.n52 VDD1.n51 9.3005
R1905 VDD1.n11 VDD1.n10 9.3005
R1906 VDD1.n58 VDD1.n57 9.3005
R1907 VDD1.n60 VDD1.n59 9.3005
R1908 VDD1.n7 VDD1.n6 9.3005
R1909 VDD1.n66 VDD1.n65 9.3005
R1910 VDD1.n68 VDD1.n67 9.3005
R1911 VDD1.n4 VDD1.n1 9.3005
R1912 VDD1.n75 VDD1.n74 9.3005
R1913 VDD1.n50 VDD1.n49 9.3005
R1914 VDD1.n15 VDD1.n14 9.3005
R1915 VDD1.n44 VDD1.n43 9.3005
R1916 VDD1.n42 VDD1.n41 9.3005
R1917 VDD1.n19 VDD1.n18 9.3005
R1918 VDD1.n36 VDD1.n35 9.3005
R1919 VDD1.n34 VDD1.n33 9.3005
R1920 VDD1.n23 VDD1.n22 9.3005
R1921 VDD1.n28 VDD1.n27 9.3005
R1922 VDD1.n154 VDD1.n153 9.3005
R1923 VDD1.n93 VDD1.n92 9.3005
R1924 VDD1.n122 VDD1.n121 9.3005
R1925 VDD1.n120 VDD1.n119 9.3005
R1926 VDD1.n97 VDD1.n96 9.3005
R1927 VDD1.n114 VDD1.n113 9.3005
R1928 VDD1.n112 VDD1.n111 9.3005
R1929 VDD1.n101 VDD1.n100 9.3005
R1930 VDD1.n106 VDD1.n105 9.3005
R1931 VDD1.n128 VDD1.n127 9.3005
R1932 VDD1.n130 VDD1.n129 9.3005
R1933 VDD1.n89 VDD1.n88 9.3005
R1934 VDD1.n136 VDD1.n135 9.3005
R1935 VDD1.n138 VDD1.n137 9.3005
R1936 VDD1.n85 VDD1.n84 9.3005
R1937 VDD1.n144 VDD1.n143 9.3005
R1938 VDD1.n146 VDD1.n145 9.3005
R1939 VDD1.n147 VDD1.n80 9.3005
R1940 VDD1.n57 VDD1.n56 8.92171
R1941 VDD1.n41 VDD1.n17 8.92171
R1942 VDD1.n119 VDD1.n95 8.92171
R1943 VDD1.n135 VDD1.n134 8.92171
R1944 VDD1.n53 VDD1.n11 8.14595
R1945 VDD1.n45 VDD1.n44 8.14595
R1946 VDD1.n123 VDD1.n122 8.14595
R1947 VDD1.n131 VDD1.n89 8.14595
R1948 VDD1.n52 VDD1.n13 7.3702
R1949 VDD1.n48 VDD1.n15 7.3702
R1950 VDD1.n126 VDD1.n93 7.3702
R1951 VDD1.n130 VDD1.n91 7.3702
R1952 VDD1.n49 VDD1.n13 6.59444
R1953 VDD1.n49 VDD1.n48 6.59444
R1954 VDD1.n127 VDD1.n126 6.59444
R1955 VDD1.n127 VDD1.n91 6.59444
R1956 VDD1.n53 VDD1.n52 5.81868
R1957 VDD1.n45 VDD1.n15 5.81868
R1958 VDD1.n123 VDD1.n93 5.81868
R1959 VDD1.n131 VDD1.n130 5.81868
R1960 VDD1.n56 VDD1.n11 5.04292
R1961 VDD1.n44 VDD1.n17 5.04292
R1962 VDD1.n122 VDD1.n95 5.04292
R1963 VDD1.n134 VDD1.n89 5.04292
R1964 VDD1.n57 VDD1.n9 4.26717
R1965 VDD1.n41 VDD1.n40 4.26717
R1966 VDD1.n119 VDD1.n118 4.26717
R1967 VDD1.n135 VDD1.n87 4.26717
R1968 VDD1.n27 VDD1.n26 3.70982
R1969 VDD1.n105 VDD1.n104 3.70982
R1970 VDD1.n61 VDD1.n60 3.49141
R1971 VDD1.n37 VDD1.n19 3.49141
R1972 VDD1.n115 VDD1.n97 3.49141
R1973 VDD1.n139 VDD1.n138 3.49141
R1974 VDD1.n64 VDD1.n7 2.71565
R1975 VDD1.n36 VDD1.n21 2.71565
R1976 VDD1.n114 VDD1.n99 2.71565
R1977 VDD1.n142 VDD1.n85 2.71565
R1978 VDD1.n160 VDD1.t7 2.32229
R1979 VDD1.n160 VDD1.t8 2.32229
R1980 VDD1.n77 VDD1.t5 2.32229
R1981 VDD1.n77 VDD1.t6 2.32229
R1982 VDD1.n158 VDD1.t0 2.32229
R1983 VDD1.n158 VDD1.t4 2.32229
R1984 VDD1.n156 VDD1.t2 2.32229
R1985 VDD1.n156 VDD1.t9 2.32229
R1986 VDD1.n65 VDD1.n5 1.93989
R1987 VDD1.n33 VDD1.n32 1.93989
R1988 VDD1.n111 VDD1.n110 1.93989
R1989 VDD1.n143 VDD1.n83 1.93989
R1990 VDD1.n76 VDD1.n0 1.16414
R1991 VDD1.n69 VDD1.n68 1.16414
R1992 VDD1.n29 VDD1.n23 1.16414
R1993 VDD1.n107 VDD1.n101 1.16414
R1994 VDD1.n148 VDD1.n146 1.16414
R1995 VDD1.n155 VDD1.n79 1.16414
R1996 VDD1 VDD1.n161 0.543603
R1997 VDD1.n74 VDD1.n73 0.388379
R1998 VDD1.n4 VDD1.n2 0.388379
R1999 VDD1.n28 VDD1.n25 0.388379
R2000 VDD1.n106 VDD1.n103 0.388379
R2001 VDD1.n147 VDD1.n81 0.388379
R2002 VDD1.n153 VDD1.n152 0.388379
R2003 VDD1 VDD1.n78 0.259121
R2004 VDD1.n75 VDD1.n1 0.155672
R2005 VDD1.n67 VDD1.n1 0.155672
R2006 VDD1.n67 VDD1.n66 0.155672
R2007 VDD1.n66 VDD1.n6 0.155672
R2008 VDD1.n59 VDD1.n6 0.155672
R2009 VDD1.n59 VDD1.n58 0.155672
R2010 VDD1.n58 VDD1.n10 0.155672
R2011 VDD1.n51 VDD1.n10 0.155672
R2012 VDD1.n51 VDD1.n50 0.155672
R2013 VDD1.n50 VDD1.n14 0.155672
R2014 VDD1.n43 VDD1.n14 0.155672
R2015 VDD1.n43 VDD1.n42 0.155672
R2016 VDD1.n42 VDD1.n18 0.155672
R2017 VDD1.n35 VDD1.n18 0.155672
R2018 VDD1.n35 VDD1.n34 0.155672
R2019 VDD1.n34 VDD1.n22 0.155672
R2020 VDD1.n27 VDD1.n22 0.155672
R2021 VDD1.n105 VDD1.n100 0.155672
R2022 VDD1.n112 VDD1.n100 0.155672
R2023 VDD1.n113 VDD1.n112 0.155672
R2024 VDD1.n113 VDD1.n96 0.155672
R2025 VDD1.n120 VDD1.n96 0.155672
R2026 VDD1.n121 VDD1.n120 0.155672
R2027 VDD1.n121 VDD1.n92 0.155672
R2028 VDD1.n128 VDD1.n92 0.155672
R2029 VDD1.n129 VDD1.n128 0.155672
R2030 VDD1.n129 VDD1.n88 0.155672
R2031 VDD1.n136 VDD1.n88 0.155672
R2032 VDD1.n137 VDD1.n136 0.155672
R2033 VDD1.n137 VDD1.n84 0.155672
R2034 VDD1.n144 VDD1.n84 0.155672
R2035 VDD1.n145 VDD1.n144 0.155672
R2036 VDD1.n145 VDD1.n80 0.155672
R2037 VDD1.n154 VDD1.n80 0.155672
R2038 VDD1.n159 VDD1.n157 0.145585
C0 B VN 0.798132f
C1 VDD1 VN 0.149203f
C2 VP VN 5.81767f
C3 VTAIL VDD2 17.3871f
C4 VDD1 B 1.80389f
C5 VP B 1.23341f
C6 VTAIL w_n2086_n3768# 3.35086f
C7 VDD1 VP 7.27138f
C8 VTAIL VN 6.80012f
C9 w_n2086_n3768# VDD2 2.1861f
C10 VDD2 VN 7.096529f
C11 w_n2086_n3768# VN 3.88317f
C12 VTAIL B 3.01233f
C13 VTAIL VDD1 17.355198f
C14 VTAIL VP 6.81484f
C15 VDD2 B 1.84434f
C16 VDD1 VDD2 0.911342f
C17 VP VDD2 0.329601f
C18 w_n2086_n3768# B 7.74782f
C19 VDD1 w_n2086_n3768# 2.14659f
C20 VP w_n2086_n3768# 4.14858f
C21 VDD2 VSUBS 1.510761f
C22 VDD1 VSUBS 1.189823f
C23 VTAIL VSUBS 0.787623f
C24 VN VSUBS 4.98672f
C25 VP VSUBS 1.771191f
C26 B VSUBS 3.055606f
C27 w_n2086_n3768# VSUBS 96.4984f
C28 VDD1.n0 VSUBS 0.028181f
C29 VDD1.n1 VSUBS 0.027446f
C30 VDD1.n2 VSUBS 0.015182f
C31 VDD1.n3 VSUBS 0.03486f
C32 VDD1.n4 VSUBS 0.014748f
C33 VDD1.n5 VSUBS 0.015616f
C34 VDD1.n6 VSUBS 0.027446f
C35 VDD1.n7 VSUBS 0.014748f
C36 VDD1.n8 VSUBS 0.03486f
C37 VDD1.n9 VSUBS 0.015616f
C38 VDD1.n10 VSUBS 0.027446f
C39 VDD1.n11 VSUBS 0.014748f
C40 VDD1.n12 VSUBS 0.03486f
C41 VDD1.n13 VSUBS 0.015616f
C42 VDD1.n14 VSUBS 0.027446f
C43 VDD1.n15 VSUBS 0.014748f
C44 VDD1.n16 VSUBS 0.03486f
C45 VDD1.n17 VSUBS 0.015616f
C46 VDD1.n18 VSUBS 0.027446f
C47 VDD1.n19 VSUBS 0.014748f
C48 VDD1.n20 VSUBS 0.03486f
C49 VDD1.n21 VSUBS 0.015616f
C50 VDD1.n22 VSUBS 0.027446f
C51 VDD1.n23 VSUBS 0.014748f
C52 VDD1.n24 VSUBS 0.026145f
C53 VDD1.n25 VSUBS 0.022176f
C54 VDD1.t3 VSUBS 0.07456f
C55 VDD1.n26 VSUBS 0.185377f
C56 VDD1.n27 VSUBS 1.6279f
C57 VDD1.n28 VSUBS 0.014748f
C58 VDD1.n29 VSUBS 0.015616f
C59 VDD1.n30 VSUBS 0.03486f
C60 VDD1.n31 VSUBS 0.03486f
C61 VDD1.n32 VSUBS 0.015616f
C62 VDD1.n33 VSUBS 0.014748f
C63 VDD1.n34 VSUBS 0.027446f
C64 VDD1.n35 VSUBS 0.027446f
C65 VDD1.n36 VSUBS 0.014748f
C66 VDD1.n37 VSUBS 0.015616f
C67 VDD1.n38 VSUBS 0.03486f
C68 VDD1.n39 VSUBS 0.03486f
C69 VDD1.n40 VSUBS 0.015616f
C70 VDD1.n41 VSUBS 0.014748f
C71 VDD1.n42 VSUBS 0.027446f
C72 VDD1.n43 VSUBS 0.027446f
C73 VDD1.n44 VSUBS 0.014748f
C74 VDD1.n45 VSUBS 0.015616f
C75 VDD1.n46 VSUBS 0.03486f
C76 VDD1.n47 VSUBS 0.03486f
C77 VDD1.n48 VSUBS 0.015616f
C78 VDD1.n49 VSUBS 0.014748f
C79 VDD1.n50 VSUBS 0.027446f
C80 VDD1.n51 VSUBS 0.027446f
C81 VDD1.n52 VSUBS 0.014748f
C82 VDD1.n53 VSUBS 0.015616f
C83 VDD1.n54 VSUBS 0.03486f
C84 VDD1.n55 VSUBS 0.03486f
C85 VDD1.n56 VSUBS 0.015616f
C86 VDD1.n57 VSUBS 0.014748f
C87 VDD1.n58 VSUBS 0.027446f
C88 VDD1.n59 VSUBS 0.027446f
C89 VDD1.n60 VSUBS 0.014748f
C90 VDD1.n61 VSUBS 0.015616f
C91 VDD1.n62 VSUBS 0.03486f
C92 VDD1.n63 VSUBS 0.03486f
C93 VDD1.n64 VSUBS 0.015616f
C94 VDD1.n65 VSUBS 0.014748f
C95 VDD1.n66 VSUBS 0.027446f
C96 VDD1.n67 VSUBS 0.027446f
C97 VDD1.n68 VSUBS 0.014748f
C98 VDD1.n69 VSUBS 0.015616f
C99 VDD1.n70 VSUBS 0.03486f
C100 VDD1.n71 VSUBS 0.03486f
C101 VDD1.n72 VSUBS 0.07766f
C102 VDD1.n73 VSUBS 0.015182f
C103 VDD1.n74 VSUBS 0.014748f
C104 VDD1.n75 VSUBS 0.06644f
C105 VDD1.n76 VSUBS 0.059739f
C106 VDD1.t5 VSUBS 0.303644f
C107 VDD1.t6 VSUBS 0.303644f
C108 VDD1.n77 VSUBS 2.44568f
C109 VDD1.n78 VSUBS 0.730663f
C110 VDD1.n79 VSUBS 0.028181f
C111 VDD1.n80 VSUBS 0.027446f
C112 VDD1.n81 VSUBS 0.015182f
C113 VDD1.n82 VSUBS 0.03486f
C114 VDD1.n83 VSUBS 0.015616f
C115 VDD1.n84 VSUBS 0.027446f
C116 VDD1.n85 VSUBS 0.014748f
C117 VDD1.n86 VSUBS 0.03486f
C118 VDD1.n87 VSUBS 0.015616f
C119 VDD1.n88 VSUBS 0.027446f
C120 VDD1.n89 VSUBS 0.014748f
C121 VDD1.n90 VSUBS 0.03486f
C122 VDD1.n91 VSUBS 0.015616f
C123 VDD1.n92 VSUBS 0.027446f
C124 VDD1.n93 VSUBS 0.014748f
C125 VDD1.n94 VSUBS 0.03486f
C126 VDD1.n95 VSUBS 0.015616f
C127 VDD1.n96 VSUBS 0.027446f
C128 VDD1.n97 VSUBS 0.014748f
C129 VDD1.n98 VSUBS 0.03486f
C130 VDD1.n99 VSUBS 0.015616f
C131 VDD1.n100 VSUBS 0.027446f
C132 VDD1.n101 VSUBS 0.014748f
C133 VDD1.n102 VSUBS 0.026145f
C134 VDD1.n103 VSUBS 0.022176f
C135 VDD1.t1 VSUBS 0.07456f
C136 VDD1.n104 VSUBS 0.185377f
C137 VDD1.n105 VSUBS 1.6279f
C138 VDD1.n106 VSUBS 0.014748f
C139 VDD1.n107 VSUBS 0.015616f
C140 VDD1.n108 VSUBS 0.03486f
C141 VDD1.n109 VSUBS 0.03486f
C142 VDD1.n110 VSUBS 0.015616f
C143 VDD1.n111 VSUBS 0.014748f
C144 VDD1.n112 VSUBS 0.027446f
C145 VDD1.n113 VSUBS 0.027446f
C146 VDD1.n114 VSUBS 0.014748f
C147 VDD1.n115 VSUBS 0.015616f
C148 VDD1.n116 VSUBS 0.03486f
C149 VDD1.n117 VSUBS 0.03486f
C150 VDD1.n118 VSUBS 0.015616f
C151 VDD1.n119 VSUBS 0.014748f
C152 VDD1.n120 VSUBS 0.027446f
C153 VDD1.n121 VSUBS 0.027446f
C154 VDD1.n122 VSUBS 0.014748f
C155 VDD1.n123 VSUBS 0.015616f
C156 VDD1.n124 VSUBS 0.03486f
C157 VDD1.n125 VSUBS 0.03486f
C158 VDD1.n126 VSUBS 0.015616f
C159 VDD1.n127 VSUBS 0.014748f
C160 VDD1.n128 VSUBS 0.027446f
C161 VDD1.n129 VSUBS 0.027446f
C162 VDD1.n130 VSUBS 0.014748f
C163 VDD1.n131 VSUBS 0.015616f
C164 VDD1.n132 VSUBS 0.03486f
C165 VDD1.n133 VSUBS 0.03486f
C166 VDD1.n134 VSUBS 0.015616f
C167 VDD1.n135 VSUBS 0.014748f
C168 VDD1.n136 VSUBS 0.027446f
C169 VDD1.n137 VSUBS 0.027446f
C170 VDD1.n138 VSUBS 0.014748f
C171 VDD1.n139 VSUBS 0.015616f
C172 VDD1.n140 VSUBS 0.03486f
C173 VDD1.n141 VSUBS 0.03486f
C174 VDD1.n142 VSUBS 0.015616f
C175 VDD1.n143 VSUBS 0.014748f
C176 VDD1.n144 VSUBS 0.027446f
C177 VDD1.n145 VSUBS 0.027446f
C178 VDD1.n146 VSUBS 0.014748f
C179 VDD1.n147 VSUBS 0.014748f
C180 VDD1.n148 VSUBS 0.015616f
C181 VDD1.n149 VSUBS 0.03486f
C182 VDD1.n150 VSUBS 0.03486f
C183 VDD1.n151 VSUBS 0.07766f
C184 VDD1.n152 VSUBS 0.015182f
C185 VDD1.n153 VSUBS 0.014748f
C186 VDD1.n154 VSUBS 0.06644f
C187 VDD1.n155 VSUBS 0.059739f
C188 VDD1.t2 VSUBS 0.303644f
C189 VDD1.t9 VSUBS 0.303644f
C190 VDD1.n156 VSUBS 2.44567f
C191 VDD1.n157 VSUBS 0.725019f
C192 VDD1.t0 VSUBS 0.303644f
C193 VDD1.t4 VSUBS 0.303644f
C194 VDD1.n158 VSUBS 2.45046f
C195 VDD1.n159 VSUBS 2.53319f
C196 VDD1.t7 VSUBS 0.303644f
C197 VDD1.t8 VSUBS 0.303644f
C198 VDD1.n160 VSUBS 2.44567f
C199 VDD1.n161 VSUBS 3.03233f
C200 VP.n0 VSUBS 0.054865f
C201 VP.t0 VSUBS 1.31093f
C202 VP.n1 VSUBS 0.525841f
C203 VP.n2 VSUBS 0.054865f
C204 VP.n3 VSUBS 0.054865f
C205 VP.t1 VSUBS 1.31093f
C206 VP.t2 VSUBS 1.31093f
C207 VP.n4 VSUBS 0.07321f
C208 VP.t3 VSUBS 1.31093f
C209 VP.n5 VSUBS 0.265187f
C210 VP.t4 VSUBS 1.31093f
C211 VP.t6 VSUBS 1.3315f
C212 VP.n6 VSUBS 0.495366f
C213 VP.n7 VSUBS 0.52492f
C214 VP.n8 VSUBS 0.525841f
C215 VP.n9 VSUBS 0.514067f
C216 VP.n10 VSUBS 0.01245f
C217 VP.n11 VSUBS 0.512714f
C218 VP.n12 VSUBS 2.42355f
C219 VP.n13 VSUBS 2.46874f
C220 VP.t8 VSUBS 1.31093f
C221 VP.n14 VSUBS 0.512714f
C222 VP.n15 VSUBS 0.01245f
C223 VP.t7 VSUBS 1.31093f
C224 VP.n16 VSUBS 0.514067f
C225 VP.n17 VSUBS 0.07321f
C226 VP.n18 VSUBS 0.073039f
C227 VP.n19 VSUBS 0.07321f
C228 VP.t9 VSUBS 1.31093f
C229 VP.n20 VSUBS 0.514067f
C230 VP.n21 VSUBS 0.01245f
C231 VP.t5 VSUBS 1.31093f
C232 VP.n22 VSUBS 0.512714f
C233 VP.n23 VSUBS 0.042518f
C234 B.n0 VSUBS 0.00632f
C235 B.n1 VSUBS 0.00632f
C236 B.n2 VSUBS 0.009347f
C237 B.n3 VSUBS 0.007163f
C238 B.n4 VSUBS 0.007163f
C239 B.n5 VSUBS 0.007163f
C240 B.n6 VSUBS 0.007163f
C241 B.n7 VSUBS 0.007163f
C242 B.n8 VSUBS 0.007163f
C243 B.n9 VSUBS 0.007163f
C244 B.n10 VSUBS 0.007163f
C245 B.n11 VSUBS 0.007163f
C246 B.n12 VSUBS 0.007163f
C247 B.n13 VSUBS 0.007163f
C248 B.n14 VSUBS 0.01662f
C249 B.n15 VSUBS 0.007163f
C250 B.n16 VSUBS 0.007163f
C251 B.n17 VSUBS 0.007163f
C252 B.n18 VSUBS 0.007163f
C253 B.n19 VSUBS 0.007163f
C254 B.n20 VSUBS 0.007163f
C255 B.n21 VSUBS 0.007163f
C256 B.n22 VSUBS 0.007163f
C257 B.n23 VSUBS 0.007163f
C258 B.n24 VSUBS 0.007163f
C259 B.n25 VSUBS 0.007163f
C260 B.n26 VSUBS 0.007163f
C261 B.n27 VSUBS 0.007163f
C262 B.n28 VSUBS 0.007163f
C263 B.n29 VSUBS 0.007163f
C264 B.n30 VSUBS 0.007163f
C265 B.n31 VSUBS 0.007163f
C266 B.n32 VSUBS 0.007163f
C267 B.n33 VSUBS 0.007163f
C268 B.n34 VSUBS 0.007163f
C269 B.n35 VSUBS 0.007163f
C270 B.n36 VSUBS 0.007163f
C271 B.n37 VSUBS 0.007163f
C272 B.t7 VSUBS 0.26217f
C273 B.t8 VSUBS 0.273371f
C274 B.t6 VSUBS 0.347877f
C275 B.n38 VSUBS 0.352767f
C276 B.n39 VSUBS 0.276966f
C277 B.n40 VSUBS 0.016595f
C278 B.n41 VSUBS 0.007163f
C279 B.n42 VSUBS 0.007163f
C280 B.n43 VSUBS 0.007163f
C281 B.n44 VSUBS 0.007163f
C282 B.n45 VSUBS 0.007163f
C283 B.t4 VSUBS 0.262173f
C284 B.t5 VSUBS 0.273374f
C285 B.t3 VSUBS 0.347877f
C286 B.n46 VSUBS 0.352763f
C287 B.n47 VSUBS 0.276963f
C288 B.n48 VSUBS 0.007163f
C289 B.n49 VSUBS 0.007163f
C290 B.n50 VSUBS 0.007163f
C291 B.n51 VSUBS 0.007163f
C292 B.n52 VSUBS 0.007163f
C293 B.n53 VSUBS 0.007163f
C294 B.n54 VSUBS 0.007163f
C295 B.n55 VSUBS 0.007163f
C296 B.n56 VSUBS 0.007163f
C297 B.n57 VSUBS 0.007163f
C298 B.n58 VSUBS 0.007163f
C299 B.n59 VSUBS 0.007163f
C300 B.n60 VSUBS 0.007163f
C301 B.n61 VSUBS 0.007163f
C302 B.n62 VSUBS 0.007163f
C303 B.n63 VSUBS 0.007163f
C304 B.n64 VSUBS 0.007163f
C305 B.n65 VSUBS 0.007163f
C306 B.n66 VSUBS 0.007163f
C307 B.n67 VSUBS 0.007163f
C308 B.n68 VSUBS 0.007163f
C309 B.n69 VSUBS 0.007163f
C310 B.n70 VSUBS 0.007163f
C311 B.n71 VSUBS 0.015402f
C312 B.n72 VSUBS 0.007163f
C313 B.n73 VSUBS 0.007163f
C314 B.n74 VSUBS 0.007163f
C315 B.n75 VSUBS 0.007163f
C316 B.n76 VSUBS 0.007163f
C317 B.n77 VSUBS 0.007163f
C318 B.n78 VSUBS 0.007163f
C319 B.n79 VSUBS 0.007163f
C320 B.n80 VSUBS 0.007163f
C321 B.n81 VSUBS 0.007163f
C322 B.n82 VSUBS 0.007163f
C323 B.n83 VSUBS 0.007163f
C324 B.n84 VSUBS 0.007163f
C325 B.n85 VSUBS 0.007163f
C326 B.n86 VSUBS 0.007163f
C327 B.n87 VSUBS 0.007163f
C328 B.n88 VSUBS 0.007163f
C329 B.n89 VSUBS 0.007163f
C330 B.n90 VSUBS 0.007163f
C331 B.n91 VSUBS 0.007163f
C332 B.n92 VSUBS 0.007163f
C333 B.n93 VSUBS 0.007163f
C334 B.n94 VSUBS 0.007163f
C335 B.n95 VSUBS 0.007163f
C336 B.n96 VSUBS 0.015712f
C337 B.n97 VSUBS 0.007163f
C338 B.n98 VSUBS 0.007163f
C339 B.n99 VSUBS 0.007163f
C340 B.n100 VSUBS 0.007163f
C341 B.n101 VSUBS 0.007163f
C342 B.n102 VSUBS 0.007163f
C343 B.n103 VSUBS 0.007163f
C344 B.n104 VSUBS 0.007163f
C345 B.n105 VSUBS 0.007163f
C346 B.n106 VSUBS 0.007163f
C347 B.n107 VSUBS 0.007163f
C348 B.n108 VSUBS 0.007163f
C349 B.n109 VSUBS 0.007163f
C350 B.n110 VSUBS 0.007163f
C351 B.n111 VSUBS 0.007163f
C352 B.n112 VSUBS 0.007163f
C353 B.n113 VSUBS 0.007163f
C354 B.n114 VSUBS 0.007163f
C355 B.n115 VSUBS 0.007163f
C356 B.n116 VSUBS 0.007163f
C357 B.n117 VSUBS 0.007163f
C358 B.n118 VSUBS 0.007163f
C359 B.n119 VSUBS 0.007163f
C360 B.t11 VSUBS 0.262173f
C361 B.t10 VSUBS 0.273374f
C362 B.t9 VSUBS 0.347877f
C363 B.n120 VSUBS 0.352763f
C364 B.n121 VSUBS 0.276963f
C365 B.n122 VSUBS 0.016595f
C366 B.n123 VSUBS 0.007163f
C367 B.n124 VSUBS 0.007163f
C368 B.n125 VSUBS 0.007163f
C369 B.n126 VSUBS 0.007163f
C370 B.n127 VSUBS 0.007163f
C371 B.t2 VSUBS 0.26217f
C372 B.t1 VSUBS 0.273371f
C373 B.t0 VSUBS 0.347877f
C374 B.n128 VSUBS 0.352767f
C375 B.n129 VSUBS 0.276966f
C376 B.n130 VSUBS 0.007163f
C377 B.n131 VSUBS 0.007163f
C378 B.n132 VSUBS 0.007163f
C379 B.n133 VSUBS 0.007163f
C380 B.n134 VSUBS 0.007163f
C381 B.n135 VSUBS 0.007163f
C382 B.n136 VSUBS 0.007163f
C383 B.n137 VSUBS 0.007163f
C384 B.n138 VSUBS 0.007163f
C385 B.n139 VSUBS 0.007163f
C386 B.n140 VSUBS 0.007163f
C387 B.n141 VSUBS 0.007163f
C388 B.n142 VSUBS 0.007163f
C389 B.n143 VSUBS 0.007163f
C390 B.n144 VSUBS 0.007163f
C391 B.n145 VSUBS 0.007163f
C392 B.n146 VSUBS 0.007163f
C393 B.n147 VSUBS 0.007163f
C394 B.n148 VSUBS 0.007163f
C395 B.n149 VSUBS 0.007163f
C396 B.n150 VSUBS 0.007163f
C397 B.n151 VSUBS 0.007163f
C398 B.n152 VSUBS 0.007163f
C399 B.n153 VSUBS 0.015402f
C400 B.n154 VSUBS 0.007163f
C401 B.n155 VSUBS 0.007163f
C402 B.n156 VSUBS 0.007163f
C403 B.n157 VSUBS 0.007163f
C404 B.n158 VSUBS 0.007163f
C405 B.n159 VSUBS 0.007163f
C406 B.n160 VSUBS 0.007163f
C407 B.n161 VSUBS 0.007163f
C408 B.n162 VSUBS 0.007163f
C409 B.n163 VSUBS 0.007163f
C410 B.n164 VSUBS 0.007163f
C411 B.n165 VSUBS 0.007163f
C412 B.n166 VSUBS 0.007163f
C413 B.n167 VSUBS 0.007163f
C414 B.n168 VSUBS 0.007163f
C415 B.n169 VSUBS 0.007163f
C416 B.n170 VSUBS 0.007163f
C417 B.n171 VSUBS 0.007163f
C418 B.n172 VSUBS 0.007163f
C419 B.n173 VSUBS 0.007163f
C420 B.n174 VSUBS 0.007163f
C421 B.n175 VSUBS 0.007163f
C422 B.n176 VSUBS 0.007163f
C423 B.n177 VSUBS 0.007163f
C424 B.n178 VSUBS 0.007163f
C425 B.n179 VSUBS 0.007163f
C426 B.n180 VSUBS 0.007163f
C427 B.n181 VSUBS 0.007163f
C428 B.n182 VSUBS 0.007163f
C429 B.n183 VSUBS 0.007163f
C430 B.n184 VSUBS 0.007163f
C431 B.n185 VSUBS 0.007163f
C432 B.n186 VSUBS 0.007163f
C433 B.n187 VSUBS 0.007163f
C434 B.n188 VSUBS 0.007163f
C435 B.n189 VSUBS 0.007163f
C436 B.n190 VSUBS 0.007163f
C437 B.n191 VSUBS 0.007163f
C438 B.n192 VSUBS 0.007163f
C439 B.n193 VSUBS 0.007163f
C440 B.n194 VSUBS 0.007163f
C441 B.n195 VSUBS 0.007163f
C442 B.n196 VSUBS 0.007163f
C443 B.n197 VSUBS 0.007163f
C444 B.n198 VSUBS 0.015402f
C445 B.n199 VSUBS 0.01662f
C446 B.n200 VSUBS 0.01662f
C447 B.n201 VSUBS 0.007163f
C448 B.n202 VSUBS 0.007163f
C449 B.n203 VSUBS 0.007163f
C450 B.n204 VSUBS 0.007163f
C451 B.n205 VSUBS 0.007163f
C452 B.n206 VSUBS 0.007163f
C453 B.n207 VSUBS 0.007163f
C454 B.n208 VSUBS 0.007163f
C455 B.n209 VSUBS 0.007163f
C456 B.n210 VSUBS 0.007163f
C457 B.n211 VSUBS 0.007163f
C458 B.n212 VSUBS 0.007163f
C459 B.n213 VSUBS 0.007163f
C460 B.n214 VSUBS 0.007163f
C461 B.n215 VSUBS 0.007163f
C462 B.n216 VSUBS 0.007163f
C463 B.n217 VSUBS 0.007163f
C464 B.n218 VSUBS 0.007163f
C465 B.n219 VSUBS 0.007163f
C466 B.n220 VSUBS 0.007163f
C467 B.n221 VSUBS 0.007163f
C468 B.n222 VSUBS 0.007163f
C469 B.n223 VSUBS 0.007163f
C470 B.n224 VSUBS 0.007163f
C471 B.n225 VSUBS 0.007163f
C472 B.n226 VSUBS 0.007163f
C473 B.n227 VSUBS 0.007163f
C474 B.n228 VSUBS 0.007163f
C475 B.n229 VSUBS 0.007163f
C476 B.n230 VSUBS 0.007163f
C477 B.n231 VSUBS 0.007163f
C478 B.n232 VSUBS 0.007163f
C479 B.n233 VSUBS 0.007163f
C480 B.n234 VSUBS 0.007163f
C481 B.n235 VSUBS 0.007163f
C482 B.n236 VSUBS 0.007163f
C483 B.n237 VSUBS 0.007163f
C484 B.n238 VSUBS 0.007163f
C485 B.n239 VSUBS 0.007163f
C486 B.n240 VSUBS 0.007163f
C487 B.n241 VSUBS 0.007163f
C488 B.n242 VSUBS 0.007163f
C489 B.n243 VSUBS 0.007163f
C490 B.n244 VSUBS 0.007163f
C491 B.n245 VSUBS 0.007163f
C492 B.n246 VSUBS 0.007163f
C493 B.n247 VSUBS 0.007163f
C494 B.n248 VSUBS 0.007163f
C495 B.n249 VSUBS 0.007163f
C496 B.n250 VSUBS 0.007163f
C497 B.n251 VSUBS 0.007163f
C498 B.n252 VSUBS 0.007163f
C499 B.n253 VSUBS 0.007163f
C500 B.n254 VSUBS 0.007163f
C501 B.n255 VSUBS 0.007163f
C502 B.n256 VSUBS 0.007163f
C503 B.n257 VSUBS 0.007163f
C504 B.n258 VSUBS 0.007163f
C505 B.n259 VSUBS 0.007163f
C506 B.n260 VSUBS 0.007163f
C507 B.n261 VSUBS 0.007163f
C508 B.n262 VSUBS 0.007163f
C509 B.n263 VSUBS 0.007163f
C510 B.n264 VSUBS 0.007163f
C511 B.n265 VSUBS 0.007163f
C512 B.n266 VSUBS 0.007163f
C513 B.n267 VSUBS 0.007163f
C514 B.n268 VSUBS 0.007163f
C515 B.n269 VSUBS 0.007163f
C516 B.n270 VSUBS 0.004951f
C517 B.n271 VSUBS 0.016595f
C518 B.n272 VSUBS 0.005793f
C519 B.n273 VSUBS 0.007163f
C520 B.n274 VSUBS 0.007163f
C521 B.n275 VSUBS 0.007163f
C522 B.n276 VSUBS 0.007163f
C523 B.n277 VSUBS 0.007163f
C524 B.n278 VSUBS 0.007163f
C525 B.n279 VSUBS 0.007163f
C526 B.n280 VSUBS 0.007163f
C527 B.n281 VSUBS 0.007163f
C528 B.n282 VSUBS 0.007163f
C529 B.n283 VSUBS 0.007163f
C530 B.n284 VSUBS 0.005793f
C531 B.n285 VSUBS 0.007163f
C532 B.n286 VSUBS 0.007163f
C533 B.n287 VSUBS 0.004951f
C534 B.n288 VSUBS 0.007163f
C535 B.n289 VSUBS 0.007163f
C536 B.n290 VSUBS 0.007163f
C537 B.n291 VSUBS 0.007163f
C538 B.n292 VSUBS 0.007163f
C539 B.n293 VSUBS 0.007163f
C540 B.n294 VSUBS 0.007163f
C541 B.n295 VSUBS 0.007163f
C542 B.n296 VSUBS 0.007163f
C543 B.n297 VSUBS 0.007163f
C544 B.n298 VSUBS 0.007163f
C545 B.n299 VSUBS 0.007163f
C546 B.n300 VSUBS 0.007163f
C547 B.n301 VSUBS 0.007163f
C548 B.n302 VSUBS 0.007163f
C549 B.n303 VSUBS 0.007163f
C550 B.n304 VSUBS 0.007163f
C551 B.n305 VSUBS 0.007163f
C552 B.n306 VSUBS 0.007163f
C553 B.n307 VSUBS 0.007163f
C554 B.n308 VSUBS 0.007163f
C555 B.n309 VSUBS 0.007163f
C556 B.n310 VSUBS 0.007163f
C557 B.n311 VSUBS 0.007163f
C558 B.n312 VSUBS 0.007163f
C559 B.n313 VSUBS 0.007163f
C560 B.n314 VSUBS 0.007163f
C561 B.n315 VSUBS 0.007163f
C562 B.n316 VSUBS 0.007163f
C563 B.n317 VSUBS 0.007163f
C564 B.n318 VSUBS 0.007163f
C565 B.n319 VSUBS 0.007163f
C566 B.n320 VSUBS 0.007163f
C567 B.n321 VSUBS 0.007163f
C568 B.n322 VSUBS 0.007163f
C569 B.n323 VSUBS 0.007163f
C570 B.n324 VSUBS 0.007163f
C571 B.n325 VSUBS 0.007163f
C572 B.n326 VSUBS 0.007163f
C573 B.n327 VSUBS 0.007163f
C574 B.n328 VSUBS 0.007163f
C575 B.n329 VSUBS 0.007163f
C576 B.n330 VSUBS 0.007163f
C577 B.n331 VSUBS 0.007163f
C578 B.n332 VSUBS 0.007163f
C579 B.n333 VSUBS 0.007163f
C580 B.n334 VSUBS 0.007163f
C581 B.n335 VSUBS 0.007163f
C582 B.n336 VSUBS 0.007163f
C583 B.n337 VSUBS 0.007163f
C584 B.n338 VSUBS 0.007163f
C585 B.n339 VSUBS 0.007163f
C586 B.n340 VSUBS 0.007163f
C587 B.n341 VSUBS 0.007163f
C588 B.n342 VSUBS 0.007163f
C589 B.n343 VSUBS 0.007163f
C590 B.n344 VSUBS 0.007163f
C591 B.n345 VSUBS 0.007163f
C592 B.n346 VSUBS 0.007163f
C593 B.n347 VSUBS 0.007163f
C594 B.n348 VSUBS 0.007163f
C595 B.n349 VSUBS 0.007163f
C596 B.n350 VSUBS 0.007163f
C597 B.n351 VSUBS 0.007163f
C598 B.n352 VSUBS 0.007163f
C599 B.n353 VSUBS 0.007163f
C600 B.n354 VSUBS 0.007163f
C601 B.n355 VSUBS 0.007163f
C602 B.n356 VSUBS 0.007163f
C603 B.n357 VSUBS 0.01662f
C604 B.n358 VSUBS 0.015402f
C605 B.n359 VSUBS 0.01631f
C606 B.n360 VSUBS 0.007163f
C607 B.n361 VSUBS 0.007163f
C608 B.n362 VSUBS 0.007163f
C609 B.n363 VSUBS 0.007163f
C610 B.n364 VSUBS 0.007163f
C611 B.n365 VSUBS 0.007163f
C612 B.n366 VSUBS 0.007163f
C613 B.n367 VSUBS 0.007163f
C614 B.n368 VSUBS 0.007163f
C615 B.n369 VSUBS 0.007163f
C616 B.n370 VSUBS 0.007163f
C617 B.n371 VSUBS 0.007163f
C618 B.n372 VSUBS 0.007163f
C619 B.n373 VSUBS 0.007163f
C620 B.n374 VSUBS 0.007163f
C621 B.n375 VSUBS 0.007163f
C622 B.n376 VSUBS 0.007163f
C623 B.n377 VSUBS 0.007163f
C624 B.n378 VSUBS 0.007163f
C625 B.n379 VSUBS 0.007163f
C626 B.n380 VSUBS 0.007163f
C627 B.n381 VSUBS 0.007163f
C628 B.n382 VSUBS 0.007163f
C629 B.n383 VSUBS 0.007163f
C630 B.n384 VSUBS 0.007163f
C631 B.n385 VSUBS 0.007163f
C632 B.n386 VSUBS 0.007163f
C633 B.n387 VSUBS 0.007163f
C634 B.n388 VSUBS 0.007163f
C635 B.n389 VSUBS 0.007163f
C636 B.n390 VSUBS 0.007163f
C637 B.n391 VSUBS 0.007163f
C638 B.n392 VSUBS 0.007163f
C639 B.n393 VSUBS 0.007163f
C640 B.n394 VSUBS 0.007163f
C641 B.n395 VSUBS 0.007163f
C642 B.n396 VSUBS 0.007163f
C643 B.n397 VSUBS 0.007163f
C644 B.n398 VSUBS 0.007163f
C645 B.n399 VSUBS 0.007163f
C646 B.n400 VSUBS 0.007163f
C647 B.n401 VSUBS 0.007163f
C648 B.n402 VSUBS 0.007163f
C649 B.n403 VSUBS 0.007163f
C650 B.n404 VSUBS 0.007163f
C651 B.n405 VSUBS 0.007163f
C652 B.n406 VSUBS 0.007163f
C653 B.n407 VSUBS 0.007163f
C654 B.n408 VSUBS 0.007163f
C655 B.n409 VSUBS 0.007163f
C656 B.n410 VSUBS 0.007163f
C657 B.n411 VSUBS 0.007163f
C658 B.n412 VSUBS 0.007163f
C659 B.n413 VSUBS 0.007163f
C660 B.n414 VSUBS 0.007163f
C661 B.n415 VSUBS 0.007163f
C662 B.n416 VSUBS 0.007163f
C663 B.n417 VSUBS 0.007163f
C664 B.n418 VSUBS 0.007163f
C665 B.n419 VSUBS 0.007163f
C666 B.n420 VSUBS 0.007163f
C667 B.n421 VSUBS 0.007163f
C668 B.n422 VSUBS 0.007163f
C669 B.n423 VSUBS 0.007163f
C670 B.n424 VSUBS 0.007163f
C671 B.n425 VSUBS 0.007163f
C672 B.n426 VSUBS 0.007163f
C673 B.n427 VSUBS 0.007163f
C674 B.n428 VSUBS 0.007163f
C675 B.n429 VSUBS 0.007163f
C676 B.n430 VSUBS 0.007163f
C677 B.n431 VSUBS 0.007163f
C678 B.n432 VSUBS 0.015402f
C679 B.n433 VSUBS 0.01662f
C680 B.n434 VSUBS 0.01662f
C681 B.n435 VSUBS 0.007163f
C682 B.n436 VSUBS 0.007163f
C683 B.n437 VSUBS 0.007163f
C684 B.n438 VSUBS 0.007163f
C685 B.n439 VSUBS 0.007163f
C686 B.n440 VSUBS 0.007163f
C687 B.n441 VSUBS 0.007163f
C688 B.n442 VSUBS 0.007163f
C689 B.n443 VSUBS 0.007163f
C690 B.n444 VSUBS 0.007163f
C691 B.n445 VSUBS 0.007163f
C692 B.n446 VSUBS 0.007163f
C693 B.n447 VSUBS 0.007163f
C694 B.n448 VSUBS 0.007163f
C695 B.n449 VSUBS 0.007163f
C696 B.n450 VSUBS 0.007163f
C697 B.n451 VSUBS 0.007163f
C698 B.n452 VSUBS 0.007163f
C699 B.n453 VSUBS 0.007163f
C700 B.n454 VSUBS 0.007163f
C701 B.n455 VSUBS 0.007163f
C702 B.n456 VSUBS 0.007163f
C703 B.n457 VSUBS 0.007163f
C704 B.n458 VSUBS 0.007163f
C705 B.n459 VSUBS 0.007163f
C706 B.n460 VSUBS 0.007163f
C707 B.n461 VSUBS 0.007163f
C708 B.n462 VSUBS 0.007163f
C709 B.n463 VSUBS 0.007163f
C710 B.n464 VSUBS 0.007163f
C711 B.n465 VSUBS 0.007163f
C712 B.n466 VSUBS 0.007163f
C713 B.n467 VSUBS 0.007163f
C714 B.n468 VSUBS 0.007163f
C715 B.n469 VSUBS 0.007163f
C716 B.n470 VSUBS 0.007163f
C717 B.n471 VSUBS 0.007163f
C718 B.n472 VSUBS 0.007163f
C719 B.n473 VSUBS 0.007163f
C720 B.n474 VSUBS 0.007163f
C721 B.n475 VSUBS 0.007163f
C722 B.n476 VSUBS 0.007163f
C723 B.n477 VSUBS 0.007163f
C724 B.n478 VSUBS 0.007163f
C725 B.n479 VSUBS 0.007163f
C726 B.n480 VSUBS 0.007163f
C727 B.n481 VSUBS 0.007163f
C728 B.n482 VSUBS 0.007163f
C729 B.n483 VSUBS 0.007163f
C730 B.n484 VSUBS 0.007163f
C731 B.n485 VSUBS 0.007163f
C732 B.n486 VSUBS 0.007163f
C733 B.n487 VSUBS 0.007163f
C734 B.n488 VSUBS 0.007163f
C735 B.n489 VSUBS 0.007163f
C736 B.n490 VSUBS 0.007163f
C737 B.n491 VSUBS 0.007163f
C738 B.n492 VSUBS 0.007163f
C739 B.n493 VSUBS 0.007163f
C740 B.n494 VSUBS 0.007163f
C741 B.n495 VSUBS 0.007163f
C742 B.n496 VSUBS 0.007163f
C743 B.n497 VSUBS 0.007163f
C744 B.n498 VSUBS 0.007163f
C745 B.n499 VSUBS 0.007163f
C746 B.n500 VSUBS 0.007163f
C747 B.n501 VSUBS 0.007163f
C748 B.n502 VSUBS 0.007163f
C749 B.n503 VSUBS 0.007163f
C750 B.n504 VSUBS 0.004951f
C751 B.n505 VSUBS 0.016595f
C752 B.n506 VSUBS 0.005793f
C753 B.n507 VSUBS 0.007163f
C754 B.n508 VSUBS 0.007163f
C755 B.n509 VSUBS 0.007163f
C756 B.n510 VSUBS 0.007163f
C757 B.n511 VSUBS 0.007163f
C758 B.n512 VSUBS 0.007163f
C759 B.n513 VSUBS 0.007163f
C760 B.n514 VSUBS 0.007163f
C761 B.n515 VSUBS 0.007163f
C762 B.n516 VSUBS 0.007163f
C763 B.n517 VSUBS 0.007163f
C764 B.n518 VSUBS 0.005793f
C765 B.n519 VSUBS 0.007163f
C766 B.n520 VSUBS 0.007163f
C767 B.n521 VSUBS 0.004951f
C768 B.n522 VSUBS 0.007163f
C769 B.n523 VSUBS 0.007163f
C770 B.n524 VSUBS 0.007163f
C771 B.n525 VSUBS 0.007163f
C772 B.n526 VSUBS 0.007163f
C773 B.n527 VSUBS 0.007163f
C774 B.n528 VSUBS 0.007163f
C775 B.n529 VSUBS 0.007163f
C776 B.n530 VSUBS 0.007163f
C777 B.n531 VSUBS 0.007163f
C778 B.n532 VSUBS 0.007163f
C779 B.n533 VSUBS 0.007163f
C780 B.n534 VSUBS 0.007163f
C781 B.n535 VSUBS 0.007163f
C782 B.n536 VSUBS 0.007163f
C783 B.n537 VSUBS 0.007163f
C784 B.n538 VSUBS 0.007163f
C785 B.n539 VSUBS 0.007163f
C786 B.n540 VSUBS 0.007163f
C787 B.n541 VSUBS 0.007163f
C788 B.n542 VSUBS 0.007163f
C789 B.n543 VSUBS 0.007163f
C790 B.n544 VSUBS 0.007163f
C791 B.n545 VSUBS 0.007163f
C792 B.n546 VSUBS 0.007163f
C793 B.n547 VSUBS 0.007163f
C794 B.n548 VSUBS 0.007163f
C795 B.n549 VSUBS 0.007163f
C796 B.n550 VSUBS 0.007163f
C797 B.n551 VSUBS 0.007163f
C798 B.n552 VSUBS 0.007163f
C799 B.n553 VSUBS 0.007163f
C800 B.n554 VSUBS 0.007163f
C801 B.n555 VSUBS 0.007163f
C802 B.n556 VSUBS 0.007163f
C803 B.n557 VSUBS 0.007163f
C804 B.n558 VSUBS 0.007163f
C805 B.n559 VSUBS 0.007163f
C806 B.n560 VSUBS 0.007163f
C807 B.n561 VSUBS 0.007163f
C808 B.n562 VSUBS 0.007163f
C809 B.n563 VSUBS 0.007163f
C810 B.n564 VSUBS 0.007163f
C811 B.n565 VSUBS 0.007163f
C812 B.n566 VSUBS 0.007163f
C813 B.n567 VSUBS 0.007163f
C814 B.n568 VSUBS 0.007163f
C815 B.n569 VSUBS 0.007163f
C816 B.n570 VSUBS 0.007163f
C817 B.n571 VSUBS 0.007163f
C818 B.n572 VSUBS 0.007163f
C819 B.n573 VSUBS 0.007163f
C820 B.n574 VSUBS 0.007163f
C821 B.n575 VSUBS 0.007163f
C822 B.n576 VSUBS 0.007163f
C823 B.n577 VSUBS 0.007163f
C824 B.n578 VSUBS 0.007163f
C825 B.n579 VSUBS 0.007163f
C826 B.n580 VSUBS 0.007163f
C827 B.n581 VSUBS 0.007163f
C828 B.n582 VSUBS 0.007163f
C829 B.n583 VSUBS 0.007163f
C830 B.n584 VSUBS 0.007163f
C831 B.n585 VSUBS 0.007163f
C832 B.n586 VSUBS 0.007163f
C833 B.n587 VSUBS 0.007163f
C834 B.n588 VSUBS 0.007163f
C835 B.n589 VSUBS 0.007163f
C836 B.n590 VSUBS 0.007163f
C837 B.n591 VSUBS 0.01662f
C838 B.n592 VSUBS 0.015402f
C839 B.n593 VSUBS 0.015402f
C840 B.n594 VSUBS 0.007163f
C841 B.n595 VSUBS 0.007163f
C842 B.n596 VSUBS 0.007163f
C843 B.n597 VSUBS 0.007163f
C844 B.n598 VSUBS 0.007163f
C845 B.n599 VSUBS 0.007163f
C846 B.n600 VSUBS 0.007163f
C847 B.n601 VSUBS 0.007163f
C848 B.n602 VSUBS 0.007163f
C849 B.n603 VSUBS 0.007163f
C850 B.n604 VSUBS 0.007163f
C851 B.n605 VSUBS 0.007163f
C852 B.n606 VSUBS 0.007163f
C853 B.n607 VSUBS 0.007163f
C854 B.n608 VSUBS 0.007163f
C855 B.n609 VSUBS 0.007163f
C856 B.n610 VSUBS 0.007163f
C857 B.n611 VSUBS 0.007163f
C858 B.n612 VSUBS 0.007163f
C859 B.n613 VSUBS 0.007163f
C860 B.n614 VSUBS 0.007163f
C861 B.n615 VSUBS 0.007163f
C862 B.n616 VSUBS 0.007163f
C863 B.n617 VSUBS 0.007163f
C864 B.n618 VSUBS 0.007163f
C865 B.n619 VSUBS 0.007163f
C866 B.n620 VSUBS 0.007163f
C867 B.n621 VSUBS 0.007163f
C868 B.n622 VSUBS 0.007163f
C869 B.n623 VSUBS 0.007163f
C870 B.n624 VSUBS 0.007163f
C871 B.n625 VSUBS 0.007163f
C872 B.n626 VSUBS 0.007163f
C873 B.n627 VSUBS 0.009347f
C874 B.n628 VSUBS 0.009957f
C875 B.n629 VSUBS 0.0198f
C876 VDD2.n0 VSUBS 0.028183f
C877 VDD2.n1 VSUBS 0.027448f
C878 VDD2.n2 VSUBS 0.015183f
C879 VDD2.n3 VSUBS 0.034862f
C880 VDD2.n4 VSUBS 0.015617f
C881 VDD2.n5 VSUBS 0.027448f
C882 VDD2.n6 VSUBS 0.014749f
C883 VDD2.n7 VSUBS 0.034862f
C884 VDD2.n8 VSUBS 0.015617f
C885 VDD2.n9 VSUBS 0.027448f
C886 VDD2.n10 VSUBS 0.014749f
C887 VDD2.n11 VSUBS 0.034862f
C888 VDD2.n12 VSUBS 0.015617f
C889 VDD2.n13 VSUBS 0.027448f
C890 VDD2.n14 VSUBS 0.014749f
C891 VDD2.n15 VSUBS 0.034862f
C892 VDD2.n16 VSUBS 0.015617f
C893 VDD2.n17 VSUBS 0.027448f
C894 VDD2.n18 VSUBS 0.014749f
C895 VDD2.n19 VSUBS 0.034862f
C896 VDD2.n20 VSUBS 0.015617f
C897 VDD2.n21 VSUBS 0.027448f
C898 VDD2.n22 VSUBS 0.014749f
C899 VDD2.n23 VSUBS 0.026146f
C900 VDD2.n24 VSUBS 0.022177f
C901 VDD2.t8 VSUBS 0.074564f
C902 VDD2.n25 VSUBS 0.185387f
C903 VDD2.n26 VSUBS 1.62798f
C904 VDD2.n27 VSUBS 0.014749f
C905 VDD2.n28 VSUBS 0.015617f
C906 VDD2.n29 VSUBS 0.034862f
C907 VDD2.n30 VSUBS 0.034862f
C908 VDD2.n31 VSUBS 0.015617f
C909 VDD2.n32 VSUBS 0.014749f
C910 VDD2.n33 VSUBS 0.027448f
C911 VDD2.n34 VSUBS 0.027448f
C912 VDD2.n35 VSUBS 0.014749f
C913 VDD2.n36 VSUBS 0.015617f
C914 VDD2.n37 VSUBS 0.034862f
C915 VDD2.n38 VSUBS 0.034862f
C916 VDD2.n39 VSUBS 0.015617f
C917 VDD2.n40 VSUBS 0.014749f
C918 VDD2.n41 VSUBS 0.027448f
C919 VDD2.n42 VSUBS 0.027448f
C920 VDD2.n43 VSUBS 0.014749f
C921 VDD2.n44 VSUBS 0.015617f
C922 VDD2.n45 VSUBS 0.034862f
C923 VDD2.n46 VSUBS 0.034862f
C924 VDD2.n47 VSUBS 0.015617f
C925 VDD2.n48 VSUBS 0.014749f
C926 VDD2.n49 VSUBS 0.027448f
C927 VDD2.n50 VSUBS 0.027448f
C928 VDD2.n51 VSUBS 0.014749f
C929 VDD2.n52 VSUBS 0.015617f
C930 VDD2.n53 VSUBS 0.034862f
C931 VDD2.n54 VSUBS 0.034862f
C932 VDD2.n55 VSUBS 0.015617f
C933 VDD2.n56 VSUBS 0.014749f
C934 VDD2.n57 VSUBS 0.027448f
C935 VDD2.n58 VSUBS 0.027448f
C936 VDD2.n59 VSUBS 0.014749f
C937 VDD2.n60 VSUBS 0.015617f
C938 VDD2.n61 VSUBS 0.034862f
C939 VDD2.n62 VSUBS 0.034862f
C940 VDD2.n63 VSUBS 0.015617f
C941 VDD2.n64 VSUBS 0.014749f
C942 VDD2.n65 VSUBS 0.027448f
C943 VDD2.n66 VSUBS 0.027448f
C944 VDD2.n67 VSUBS 0.014749f
C945 VDD2.n68 VSUBS 0.014749f
C946 VDD2.n69 VSUBS 0.015617f
C947 VDD2.n70 VSUBS 0.034862f
C948 VDD2.n71 VSUBS 0.034862f
C949 VDD2.n72 VSUBS 0.077664f
C950 VDD2.n73 VSUBS 0.015183f
C951 VDD2.n74 VSUBS 0.014749f
C952 VDD2.n75 VSUBS 0.066444f
C953 VDD2.n76 VSUBS 0.059742f
C954 VDD2.t1 VSUBS 0.30366f
C955 VDD2.t0 VSUBS 0.30366f
C956 VDD2.n77 VSUBS 2.44579f
C957 VDD2.n78 VSUBS 0.725056f
C958 VDD2.t3 VSUBS 0.30366f
C959 VDD2.t2 VSUBS 0.30366f
C960 VDD2.n79 VSUBS 2.45059f
C961 VDD2.n80 VSUBS 2.45077f
C962 VDD2.n81 VSUBS 0.028183f
C963 VDD2.n82 VSUBS 0.027448f
C964 VDD2.n83 VSUBS 0.015183f
C965 VDD2.n84 VSUBS 0.034862f
C966 VDD2.n85 VSUBS 0.014749f
C967 VDD2.n86 VSUBS 0.015617f
C968 VDD2.n87 VSUBS 0.027448f
C969 VDD2.n88 VSUBS 0.014749f
C970 VDD2.n89 VSUBS 0.034862f
C971 VDD2.n90 VSUBS 0.015617f
C972 VDD2.n91 VSUBS 0.027448f
C973 VDD2.n92 VSUBS 0.014749f
C974 VDD2.n93 VSUBS 0.034862f
C975 VDD2.n94 VSUBS 0.015617f
C976 VDD2.n95 VSUBS 0.027448f
C977 VDD2.n96 VSUBS 0.014749f
C978 VDD2.n97 VSUBS 0.034862f
C979 VDD2.n98 VSUBS 0.015617f
C980 VDD2.n99 VSUBS 0.027448f
C981 VDD2.n100 VSUBS 0.014749f
C982 VDD2.n101 VSUBS 0.034862f
C983 VDD2.n102 VSUBS 0.015617f
C984 VDD2.n103 VSUBS 0.027448f
C985 VDD2.n104 VSUBS 0.014749f
C986 VDD2.n105 VSUBS 0.026146f
C987 VDD2.n106 VSUBS 0.022177f
C988 VDD2.t9 VSUBS 0.074564f
C989 VDD2.n107 VSUBS 0.185387f
C990 VDD2.n108 VSUBS 1.62798f
C991 VDD2.n109 VSUBS 0.014749f
C992 VDD2.n110 VSUBS 0.015617f
C993 VDD2.n111 VSUBS 0.034862f
C994 VDD2.n112 VSUBS 0.034862f
C995 VDD2.n113 VSUBS 0.015617f
C996 VDD2.n114 VSUBS 0.014749f
C997 VDD2.n115 VSUBS 0.027448f
C998 VDD2.n116 VSUBS 0.027448f
C999 VDD2.n117 VSUBS 0.014749f
C1000 VDD2.n118 VSUBS 0.015617f
C1001 VDD2.n119 VSUBS 0.034862f
C1002 VDD2.n120 VSUBS 0.034862f
C1003 VDD2.n121 VSUBS 0.015617f
C1004 VDD2.n122 VSUBS 0.014749f
C1005 VDD2.n123 VSUBS 0.027448f
C1006 VDD2.n124 VSUBS 0.027448f
C1007 VDD2.n125 VSUBS 0.014749f
C1008 VDD2.n126 VSUBS 0.015617f
C1009 VDD2.n127 VSUBS 0.034862f
C1010 VDD2.n128 VSUBS 0.034862f
C1011 VDD2.n129 VSUBS 0.015617f
C1012 VDD2.n130 VSUBS 0.014749f
C1013 VDD2.n131 VSUBS 0.027448f
C1014 VDD2.n132 VSUBS 0.027448f
C1015 VDD2.n133 VSUBS 0.014749f
C1016 VDD2.n134 VSUBS 0.015617f
C1017 VDD2.n135 VSUBS 0.034862f
C1018 VDD2.n136 VSUBS 0.034862f
C1019 VDD2.n137 VSUBS 0.015617f
C1020 VDD2.n138 VSUBS 0.014749f
C1021 VDD2.n139 VSUBS 0.027448f
C1022 VDD2.n140 VSUBS 0.027448f
C1023 VDD2.n141 VSUBS 0.014749f
C1024 VDD2.n142 VSUBS 0.015617f
C1025 VDD2.n143 VSUBS 0.034862f
C1026 VDD2.n144 VSUBS 0.034862f
C1027 VDD2.n145 VSUBS 0.015617f
C1028 VDD2.n146 VSUBS 0.014749f
C1029 VDD2.n147 VSUBS 0.027448f
C1030 VDD2.n148 VSUBS 0.027448f
C1031 VDD2.n149 VSUBS 0.014749f
C1032 VDD2.n150 VSUBS 0.015617f
C1033 VDD2.n151 VSUBS 0.034862f
C1034 VDD2.n152 VSUBS 0.034862f
C1035 VDD2.n153 VSUBS 0.077664f
C1036 VDD2.n154 VSUBS 0.015183f
C1037 VDD2.n155 VSUBS 0.014749f
C1038 VDD2.n156 VSUBS 0.066444f
C1039 VDD2.n157 VSUBS 0.057778f
C1040 VDD2.n158 VSUBS 2.49573f
C1041 VDD2.t7 VSUBS 0.30366f
C1042 VDD2.t6 VSUBS 0.30366f
C1043 VDD2.n159 VSUBS 2.4458f
C1044 VDD2.n160 VSUBS 0.607188f
C1045 VDD2.t4 VSUBS 0.30366f
C1046 VDD2.t5 VSUBS 0.30366f
C1047 VDD2.n161 VSUBS 2.45055f
C1048 VTAIL.t11 VSUBS 0.327164f
C1049 VTAIL.t13 VSUBS 0.327164f
C1050 VTAIL.n0 VSUBS 2.47263f
C1051 VTAIL.n1 VSUBS 0.821248f
C1052 VTAIL.n2 VSUBS 0.030364f
C1053 VTAIL.n3 VSUBS 0.029572f
C1054 VTAIL.n4 VSUBS 0.016358f
C1055 VTAIL.n5 VSUBS 0.03756f
C1056 VTAIL.n6 VSUBS 0.016826f
C1057 VTAIL.n7 VSUBS 0.029572f
C1058 VTAIL.n8 VSUBS 0.015891f
C1059 VTAIL.n9 VSUBS 0.03756f
C1060 VTAIL.n10 VSUBS 0.016826f
C1061 VTAIL.n11 VSUBS 0.029572f
C1062 VTAIL.n12 VSUBS 0.015891f
C1063 VTAIL.n13 VSUBS 0.03756f
C1064 VTAIL.n14 VSUBS 0.016826f
C1065 VTAIL.n15 VSUBS 0.029572f
C1066 VTAIL.n16 VSUBS 0.015891f
C1067 VTAIL.n17 VSUBS 0.03756f
C1068 VTAIL.n18 VSUBS 0.016826f
C1069 VTAIL.n19 VSUBS 0.029572f
C1070 VTAIL.n20 VSUBS 0.015891f
C1071 VTAIL.n21 VSUBS 0.03756f
C1072 VTAIL.n22 VSUBS 0.016826f
C1073 VTAIL.n23 VSUBS 0.029572f
C1074 VTAIL.n24 VSUBS 0.015891f
C1075 VTAIL.n25 VSUBS 0.02817f
C1076 VTAIL.n26 VSUBS 0.023894f
C1077 VTAIL.t4 VSUBS 0.080336f
C1078 VTAIL.n27 VSUBS 0.199736f
C1079 VTAIL.n28 VSUBS 1.75399f
C1080 VTAIL.n29 VSUBS 0.015891f
C1081 VTAIL.n30 VSUBS 0.016826f
C1082 VTAIL.n31 VSUBS 0.03756f
C1083 VTAIL.n32 VSUBS 0.03756f
C1084 VTAIL.n33 VSUBS 0.016826f
C1085 VTAIL.n34 VSUBS 0.015891f
C1086 VTAIL.n35 VSUBS 0.029572f
C1087 VTAIL.n36 VSUBS 0.029572f
C1088 VTAIL.n37 VSUBS 0.015891f
C1089 VTAIL.n38 VSUBS 0.016826f
C1090 VTAIL.n39 VSUBS 0.03756f
C1091 VTAIL.n40 VSUBS 0.03756f
C1092 VTAIL.n41 VSUBS 0.016826f
C1093 VTAIL.n42 VSUBS 0.015891f
C1094 VTAIL.n43 VSUBS 0.029572f
C1095 VTAIL.n44 VSUBS 0.029572f
C1096 VTAIL.n45 VSUBS 0.015891f
C1097 VTAIL.n46 VSUBS 0.016826f
C1098 VTAIL.n47 VSUBS 0.03756f
C1099 VTAIL.n48 VSUBS 0.03756f
C1100 VTAIL.n49 VSUBS 0.016826f
C1101 VTAIL.n50 VSUBS 0.015891f
C1102 VTAIL.n51 VSUBS 0.029572f
C1103 VTAIL.n52 VSUBS 0.029572f
C1104 VTAIL.n53 VSUBS 0.015891f
C1105 VTAIL.n54 VSUBS 0.016826f
C1106 VTAIL.n55 VSUBS 0.03756f
C1107 VTAIL.n56 VSUBS 0.03756f
C1108 VTAIL.n57 VSUBS 0.016826f
C1109 VTAIL.n58 VSUBS 0.015891f
C1110 VTAIL.n59 VSUBS 0.029572f
C1111 VTAIL.n60 VSUBS 0.029572f
C1112 VTAIL.n61 VSUBS 0.015891f
C1113 VTAIL.n62 VSUBS 0.016826f
C1114 VTAIL.n63 VSUBS 0.03756f
C1115 VTAIL.n64 VSUBS 0.03756f
C1116 VTAIL.n65 VSUBS 0.016826f
C1117 VTAIL.n66 VSUBS 0.015891f
C1118 VTAIL.n67 VSUBS 0.029572f
C1119 VTAIL.n68 VSUBS 0.029572f
C1120 VTAIL.n69 VSUBS 0.015891f
C1121 VTAIL.n70 VSUBS 0.015891f
C1122 VTAIL.n71 VSUBS 0.016826f
C1123 VTAIL.n72 VSUBS 0.03756f
C1124 VTAIL.n73 VSUBS 0.03756f
C1125 VTAIL.n74 VSUBS 0.083676f
C1126 VTAIL.n75 VSUBS 0.016358f
C1127 VTAIL.n76 VSUBS 0.015891f
C1128 VTAIL.n77 VSUBS 0.071587f
C1129 VTAIL.n78 VSUBS 0.041855f
C1130 VTAIL.n79 VSUBS 0.186444f
C1131 VTAIL.t2 VSUBS 0.327164f
C1132 VTAIL.t19 VSUBS 0.327164f
C1133 VTAIL.n80 VSUBS 2.47263f
C1134 VTAIL.n81 VSUBS 0.82823f
C1135 VTAIL.t0 VSUBS 0.327164f
C1136 VTAIL.t6 VSUBS 0.327164f
C1137 VTAIL.n82 VSUBS 2.47263f
C1138 VTAIL.n83 VSUBS 2.45636f
C1139 VTAIL.t14 VSUBS 0.327164f
C1140 VTAIL.t10 VSUBS 0.327164f
C1141 VTAIL.n84 VSUBS 2.47264f
C1142 VTAIL.n85 VSUBS 2.45634f
C1143 VTAIL.t12 VSUBS 0.327164f
C1144 VTAIL.t15 VSUBS 0.327164f
C1145 VTAIL.n86 VSUBS 2.47264f
C1146 VTAIL.n87 VSUBS 0.828214f
C1147 VTAIL.n88 VSUBS 0.030364f
C1148 VTAIL.n89 VSUBS 0.029572f
C1149 VTAIL.n90 VSUBS 0.016358f
C1150 VTAIL.n91 VSUBS 0.03756f
C1151 VTAIL.n92 VSUBS 0.015891f
C1152 VTAIL.n93 VSUBS 0.016826f
C1153 VTAIL.n94 VSUBS 0.029572f
C1154 VTAIL.n95 VSUBS 0.015891f
C1155 VTAIL.n96 VSUBS 0.03756f
C1156 VTAIL.n97 VSUBS 0.016826f
C1157 VTAIL.n98 VSUBS 0.029572f
C1158 VTAIL.n99 VSUBS 0.015891f
C1159 VTAIL.n100 VSUBS 0.03756f
C1160 VTAIL.n101 VSUBS 0.016826f
C1161 VTAIL.n102 VSUBS 0.029572f
C1162 VTAIL.n103 VSUBS 0.015891f
C1163 VTAIL.n104 VSUBS 0.03756f
C1164 VTAIL.n105 VSUBS 0.016826f
C1165 VTAIL.n106 VSUBS 0.029572f
C1166 VTAIL.n107 VSUBS 0.015891f
C1167 VTAIL.n108 VSUBS 0.03756f
C1168 VTAIL.n109 VSUBS 0.016826f
C1169 VTAIL.n110 VSUBS 0.029572f
C1170 VTAIL.n111 VSUBS 0.015891f
C1171 VTAIL.n112 VSUBS 0.02817f
C1172 VTAIL.n113 VSUBS 0.023894f
C1173 VTAIL.t8 VSUBS 0.080336f
C1174 VTAIL.n114 VSUBS 0.199736f
C1175 VTAIL.n115 VSUBS 1.75399f
C1176 VTAIL.n116 VSUBS 0.015891f
C1177 VTAIL.n117 VSUBS 0.016826f
C1178 VTAIL.n118 VSUBS 0.03756f
C1179 VTAIL.n119 VSUBS 0.03756f
C1180 VTAIL.n120 VSUBS 0.016826f
C1181 VTAIL.n121 VSUBS 0.015891f
C1182 VTAIL.n122 VSUBS 0.029572f
C1183 VTAIL.n123 VSUBS 0.029572f
C1184 VTAIL.n124 VSUBS 0.015891f
C1185 VTAIL.n125 VSUBS 0.016826f
C1186 VTAIL.n126 VSUBS 0.03756f
C1187 VTAIL.n127 VSUBS 0.03756f
C1188 VTAIL.n128 VSUBS 0.016826f
C1189 VTAIL.n129 VSUBS 0.015891f
C1190 VTAIL.n130 VSUBS 0.029572f
C1191 VTAIL.n131 VSUBS 0.029572f
C1192 VTAIL.n132 VSUBS 0.015891f
C1193 VTAIL.n133 VSUBS 0.016826f
C1194 VTAIL.n134 VSUBS 0.03756f
C1195 VTAIL.n135 VSUBS 0.03756f
C1196 VTAIL.n136 VSUBS 0.016826f
C1197 VTAIL.n137 VSUBS 0.015891f
C1198 VTAIL.n138 VSUBS 0.029572f
C1199 VTAIL.n139 VSUBS 0.029572f
C1200 VTAIL.n140 VSUBS 0.015891f
C1201 VTAIL.n141 VSUBS 0.016826f
C1202 VTAIL.n142 VSUBS 0.03756f
C1203 VTAIL.n143 VSUBS 0.03756f
C1204 VTAIL.n144 VSUBS 0.016826f
C1205 VTAIL.n145 VSUBS 0.015891f
C1206 VTAIL.n146 VSUBS 0.029572f
C1207 VTAIL.n147 VSUBS 0.029572f
C1208 VTAIL.n148 VSUBS 0.015891f
C1209 VTAIL.n149 VSUBS 0.016826f
C1210 VTAIL.n150 VSUBS 0.03756f
C1211 VTAIL.n151 VSUBS 0.03756f
C1212 VTAIL.n152 VSUBS 0.016826f
C1213 VTAIL.n153 VSUBS 0.015891f
C1214 VTAIL.n154 VSUBS 0.029572f
C1215 VTAIL.n155 VSUBS 0.029572f
C1216 VTAIL.n156 VSUBS 0.015891f
C1217 VTAIL.n157 VSUBS 0.016826f
C1218 VTAIL.n158 VSUBS 0.03756f
C1219 VTAIL.n159 VSUBS 0.03756f
C1220 VTAIL.n160 VSUBS 0.083676f
C1221 VTAIL.n161 VSUBS 0.016358f
C1222 VTAIL.n162 VSUBS 0.015891f
C1223 VTAIL.n163 VSUBS 0.071587f
C1224 VTAIL.n164 VSUBS 0.041855f
C1225 VTAIL.n165 VSUBS 0.186444f
C1226 VTAIL.t18 VSUBS 0.327164f
C1227 VTAIL.t7 VSUBS 0.327164f
C1228 VTAIL.n166 VSUBS 2.47264f
C1229 VTAIL.n167 VSUBS 0.834786f
C1230 VTAIL.t5 VSUBS 0.327164f
C1231 VTAIL.t3 VSUBS 0.327164f
C1232 VTAIL.n168 VSUBS 2.47264f
C1233 VTAIL.n169 VSUBS 0.828214f
C1234 VTAIL.n170 VSUBS 0.030364f
C1235 VTAIL.n171 VSUBS 0.029572f
C1236 VTAIL.n172 VSUBS 0.016358f
C1237 VTAIL.n173 VSUBS 0.03756f
C1238 VTAIL.n174 VSUBS 0.015891f
C1239 VTAIL.n175 VSUBS 0.016826f
C1240 VTAIL.n176 VSUBS 0.029572f
C1241 VTAIL.n177 VSUBS 0.015891f
C1242 VTAIL.n178 VSUBS 0.03756f
C1243 VTAIL.n179 VSUBS 0.016826f
C1244 VTAIL.n180 VSUBS 0.029572f
C1245 VTAIL.n181 VSUBS 0.015891f
C1246 VTAIL.n182 VSUBS 0.03756f
C1247 VTAIL.n183 VSUBS 0.016826f
C1248 VTAIL.n184 VSUBS 0.029572f
C1249 VTAIL.n185 VSUBS 0.015891f
C1250 VTAIL.n186 VSUBS 0.03756f
C1251 VTAIL.n187 VSUBS 0.016826f
C1252 VTAIL.n188 VSUBS 0.029572f
C1253 VTAIL.n189 VSUBS 0.015891f
C1254 VTAIL.n190 VSUBS 0.03756f
C1255 VTAIL.n191 VSUBS 0.016826f
C1256 VTAIL.n192 VSUBS 0.029572f
C1257 VTAIL.n193 VSUBS 0.015891f
C1258 VTAIL.n194 VSUBS 0.02817f
C1259 VTAIL.n195 VSUBS 0.023894f
C1260 VTAIL.t1 VSUBS 0.080336f
C1261 VTAIL.n196 VSUBS 0.199736f
C1262 VTAIL.n197 VSUBS 1.75399f
C1263 VTAIL.n198 VSUBS 0.015891f
C1264 VTAIL.n199 VSUBS 0.016826f
C1265 VTAIL.n200 VSUBS 0.03756f
C1266 VTAIL.n201 VSUBS 0.03756f
C1267 VTAIL.n202 VSUBS 0.016826f
C1268 VTAIL.n203 VSUBS 0.015891f
C1269 VTAIL.n204 VSUBS 0.029572f
C1270 VTAIL.n205 VSUBS 0.029572f
C1271 VTAIL.n206 VSUBS 0.015891f
C1272 VTAIL.n207 VSUBS 0.016826f
C1273 VTAIL.n208 VSUBS 0.03756f
C1274 VTAIL.n209 VSUBS 0.03756f
C1275 VTAIL.n210 VSUBS 0.016826f
C1276 VTAIL.n211 VSUBS 0.015891f
C1277 VTAIL.n212 VSUBS 0.029572f
C1278 VTAIL.n213 VSUBS 0.029572f
C1279 VTAIL.n214 VSUBS 0.015891f
C1280 VTAIL.n215 VSUBS 0.016826f
C1281 VTAIL.n216 VSUBS 0.03756f
C1282 VTAIL.n217 VSUBS 0.03756f
C1283 VTAIL.n218 VSUBS 0.016826f
C1284 VTAIL.n219 VSUBS 0.015891f
C1285 VTAIL.n220 VSUBS 0.029572f
C1286 VTAIL.n221 VSUBS 0.029572f
C1287 VTAIL.n222 VSUBS 0.015891f
C1288 VTAIL.n223 VSUBS 0.016826f
C1289 VTAIL.n224 VSUBS 0.03756f
C1290 VTAIL.n225 VSUBS 0.03756f
C1291 VTAIL.n226 VSUBS 0.016826f
C1292 VTAIL.n227 VSUBS 0.015891f
C1293 VTAIL.n228 VSUBS 0.029572f
C1294 VTAIL.n229 VSUBS 0.029572f
C1295 VTAIL.n230 VSUBS 0.015891f
C1296 VTAIL.n231 VSUBS 0.016826f
C1297 VTAIL.n232 VSUBS 0.03756f
C1298 VTAIL.n233 VSUBS 0.03756f
C1299 VTAIL.n234 VSUBS 0.016826f
C1300 VTAIL.n235 VSUBS 0.015891f
C1301 VTAIL.n236 VSUBS 0.029572f
C1302 VTAIL.n237 VSUBS 0.029572f
C1303 VTAIL.n238 VSUBS 0.015891f
C1304 VTAIL.n239 VSUBS 0.016826f
C1305 VTAIL.n240 VSUBS 0.03756f
C1306 VTAIL.n241 VSUBS 0.03756f
C1307 VTAIL.n242 VSUBS 0.083676f
C1308 VTAIL.n243 VSUBS 0.016358f
C1309 VTAIL.n244 VSUBS 0.015891f
C1310 VTAIL.n245 VSUBS 0.071587f
C1311 VTAIL.n246 VSUBS 0.041855f
C1312 VTAIL.n247 VSUBS 1.73161f
C1313 VTAIL.n248 VSUBS 0.030364f
C1314 VTAIL.n249 VSUBS 0.029572f
C1315 VTAIL.n250 VSUBS 0.016358f
C1316 VTAIL.n251 VSUBS 0.03756f
C1317 VTAIL.n252 VSUBS 0.016826f
C1318 VTAIL.n253 VSUBS 0.029572f
C1319 VTAIL.n254 VSUBS 0.015891f
C1320 VTAIL.n255 VSUBS 0.03756f
C1321 VTAIL.n256 VSUBS 0.016826f
C1322 VTAIL.n257 VSUBS 0.029572f
C1323 VTAIL.n258 VSUBS 0.015891f
C1324 VTAIL.n259 VSUBS 0.03756f
C1325 VTAIL.n260 VSUBS 0.016826f
C1326 VTAIL.n261 VSUBS 0.029572f
C1327 VTAIL.n262 VSUBS 0.015891f
C1328 VTAIL.n263 VSUBS 0.03756f
C1329 VTAIL.n264 VSUBS 0.016826f
C1330 VTAIL.n265 VSUBS 0.029572f
C1331 VTAIL.n266 VSUBS 0.015891f
C1332 VTAIL.n267 VSUBS 0.03756f
C1333 VTAIL.n268 VSUBS 0.016826f
C1334 VTAIL.n269 VSUBS 0.029572f
C1335 VTAIL.n270 VSUBS 0.015891f
C1336 VTAIL.n271 VSUBS 0.02817f
C1337 VTAIL.n272 VSUBS 0.023894f
C1338 VTAIL.t17 VSUBS 0.080336f
C1339 VTAIL.n273 VSUBS 0.199736f
C1340 VTAIL.n274 VSUBS 1.75399f
C1341 VTAIL.n275 VSUBS 0.015891f
C1342 VTAIL.n276 VSUBS 0.016826f
C1343 VTAIL.n277 VSUBS 0.03756f
C1344 VTAIL.n278 VSUBS 0.03756f
C1345 VTAIL.n279 VSUBS 0.016826f
C1346 VTAIL.n280 VSUBS 0.015891f
C1347 VTAIL.n281 VSUBS 0.029572f
C1348 VTAIL.n282 VSUBS 0.029572f
C1349 VTAIL.n283 VSUBS 0.015891f
C1350 VTAIL.n284 VSUBS 0.016826f
C1351 VTAIL.n285 VSUBS 0.03756f
C1352 VTAIL.n286 VSUBS 0.03756f
C1353 VTAIL.n287 VSUBS 0.016826f
C1354 VTAIL.n288 VSUBS 0.015891f
C1355 VTAIL.n289 VSUBS 0.029572f
C1356 VTAIL.n290 VSUBS 0.029572f
C1357 VTAIL.n291 VSUBS 0.015891f
C1358 VTAIL.n292 VSUBS 0.016826f
C1359 VTAIL.n293 VSUBS 0.03756f
C1360 VTAIL.n294 VSUBS 0.03756f
C1361 VTAIL.n295 VSUBS 0.016826f
C1362 VTAIL.n296 VSUBS 0.015891f
C1363 VTAIL.n297 VSUBS 0.029572f
C1364 VTAIL.n298 VSUBS 0.029572f
C1365 VTAIL.n299 VSUBS 0.015891f
C1366 VTAIL.n300 VSUBS 0.016826f
C1367 VTAIL.n301 VSUBS 0.03756f
C1368 VTAIL.n302 VSUBS 0.03756f
C1369 VTAIL.n303 VSUBS 0.016826f
C1370 VTAIL.n304 VSUBS 0.015891f
C1371 VTAIL.n305 VSUBS 0.029572f
C1372 VTAIL.n306 VSUBS 0.029572f
C1373 VTAIL.n307 VSUBS 0.015891f
C1374 VTAIL.n308 VSUBS 0.016826f
C1375 VTAIL.n309 VSUBS 0.03756f
C1376 VTAIL.n310 VSUBS 0.03756f
C1377 VTAIL.n311 VSUBS 0.016826f
C1378 VTAIL.n312 VSUBS 0.015891f
C1379 VTAIL.n313 VSUBS 0.029572f
C1380 VTAIL.n314 VSUBS 0.029572f
C1381 VTAIL.n315 VSUBS 0.015891f
C1382 VTAIL.n316 VSUBS 0.015891f
C1383 VTAIL.n317 VSUBS 0.016826f
C1384 VTAIL.n318 VSUBS 0.03756f
C1385 VTAIL.n319 VSUBS 0.03756f
C1386 VTAIL.n320 VSUBS 0.083676f
C1387 VTAIL.n321 VSUBS 0.016358f
C1388 VTAIL.n322 VSUBS 0.015891f
C1389 VTAIL.n323 VSUBS 0.071587f
C1390 VTAIL.n324 VSUBS 0.041855f
C1391 VTAIL.n325 VSUBS 1.73161f
C1392 VTAIL.t9 VSUBS 0.327164f
C1393 VTAIL.t16 VSUBS 0.327164f
C1394 VTAIL.n326 VSUBS 2.47263f
C1395 VTAIL.n327 VSUBS 0.765389f
C1396 VN.n0 VSUBS 0.053778f
C1397 VN.t9 VSUBS 1.28496f
C1398 VN.n1 VSUBS 0.515421f
C1399 VN.t1 VSUBS 1.30511f
C1400 VN.t8 VSUBS 1.28496f
C1401 VN.n2 VSUBS 0.514518f
C1402 VN.n3 VSUBS 0.48555f
C1403 VN.n4 VSUBS 0.259932f
C1404 VN.n5 VSUBS 0.07176f
C1405 VN.t6 VSUBS 1.28496f
C1406 VN.n6 VSUBS 0.50388f
C1407 VN.n7 VSUBS 0.012203f
C1408 VN.t7 VSUBS 1.28496f
C1409 VN.n8 VSUBS 0.502554f
C1410 VN.n9 VSUBS 0.041676f
C1411 VN.n10 VSUBS 0.053778f
C1412 VN.t3 VSUBS 1.28496f
C1413 VN.n11 VSUBS 0.515421f
C1414 VN.t2 VSUBS 1.28496f
C1415 VN.t4 VSUBS 1.30511f
C1416 VN.t5 VSUBS 1.28496f
C1417 VN.n12 VSUBS 0.514518f
C1418 VN.n13 VSUBS 0.48555f
C1419 VN.n14 VSUBS 0.259932f
C1420 VN.n15 VSUBS 0.07176f
C1421 VN.n16 VSUBS 0.50388f
C1422 VN.n17 VSUBS 0.012203f
C1423 VN.t0 VSUBS 1.28496f
C1424 VN.n18 VSUBS 0.502554f
C1425 VN.n19 VSUBS 2.41074f
.ends

