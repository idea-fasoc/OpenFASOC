* NGSPICE file created from diff_pair_sample_0489.ext - technology: sky130A

.subckt diff_pair_sample_0489 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=0 ps=0 w=17.14 l=0.22
X1 VDD1.t9 VP.t0 VTAIL.t11 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=2.8281 ps=17.47 w=17.14 l=0.22
X2 VDD1.t8 VP.t1 VTAIL.t18 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=6.6846 ps=35.06 w=17.14 l=0.22
X3 VDD1.t7 VP.t2 VTAIL.t17 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X4 VDD1.t6 VP.t3 VTAIL.t15 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X5 VDD2.t9 VN.t0 VTAIL.t7 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=2.8281 ps=17.47 w=17.14 l=0.22
X6 VTAIL.t4 VN.t1 VDD2.t8 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X7 VDD2.t7 VN.t2 VTAIL.t5 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X8 B.t8 B.t6 B.t7 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=0 ps=0 w=17.14 l=0.22
X9 VDD2.t6 VN.t3 VTAIL.t9 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=6.6846 ps=35.06 w=17.14 l=0.22
X10 VTAIL.t14 VP.t4 VDD1.t5 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X11 B.t5 B.t3 B.t4 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=0 ps=0 w=17.14 l=0.22
X12 VTAIL.t13 VP.t5 VDD1.t4 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X13 VDD1.t3 VP.t6 VTAIL.t12 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=2.8281 ps=17.47 w=17.14 l=0.22
X14 B.t2 B.t0 B.t1 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=0 ps=0 w=17.14 l=0.22
X15 VDD2.t5 VN.t4 VTAIL.t3 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X16 VTAIL.t6 VN.t5 VDD2.t4 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X17 VTAIL.t19 VP.t7 VDD1.t2 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X18 VTAIL.t8 VN.t6 VDD2.t3 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X19 VDD1.t1 VP.t8 VTAIL.t16 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=6.6846 ps=35.06 w=17.14 l=0.22
X20 VTAIL.t10 VP.t9 VDD1.t0 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X21 VTAIL.t0 VN.t7 VDD2.t2 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=2.8281 ps=17.47 w=17.14 l=0.22
X22 VDD2.t1 VN.t8 VTAIL.t1 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=2.8281 pd=17.47 as=6.6846 ps=35.06 w=17.14 l=0.22
X23 VDD2.t0 VN.t9 VTAIL.t2 w_n1630_n4396# sky130_fd_pr__pfet_01v8 ad=6.6846 pd=35.06 as=2.8281 ps=17.47 w=17.14 l=0.22
R0 B.n124 B.t6 2108.48
R1 B.n132 B.t3 2108.48
R2 B.n40 B.t9 2108.48
R3 B.n46 B.t0 2108.48
R4 B.n438 B.n437 585
R5 B.n439 B.n76 585
R6 B.n441 B.n440 585
R7 B.n442 B.n75 585
R8 B.n444 B.n443 585
R9 B.n445 B.n74 585
R10 B.n447 B.n446 585
R11 B.n448 B.n73 585
R12 B.n450 B.n449 585
R13 B.n451 B.n72 585
R14 B.n453 B.n452 585
R15 B.n454 B.n71 585
R16 B.n456 B.n455 585
R17 B.n457 B.n70 585
R18 B.n459 B.n458 585
R19 B.n460 B.n69 585
R20 B.n462 B.n461 585
R21 B.n463 B.n68 585
R22 B.n465 B.n464 585
R23 B.n466 B.n67 585
R24 B.n468 B.n467 585
R25 B.n469 B.n66 585
R26 B.n471 B.n470 585
R27 B.n472 B.n65 585
R28 B.n474 B.n473 585
R29 B.n475 B.n64 585
R30 B.n477 B.n476 585
R31 B.n478 B.n63 585
R32 B.n480 B.n479 585
R33 B.n481 B.n62 585
R34 B.n483 B.n482 585
R35 B.n484 B.n61 585
R36 B.n486 B.n485 585
R37 B.n487 B.n60 585
R38 B.n489 B.n488 585
R39 B.n490 B.n59 585
R40 B.n492 B.n491 585
R41 B.n493 B.n58 585
R42 B.n495 B.n494 585
R43 B.n496 B.n57 585
R44 B.n498 B.n497 585
R45 B.n499 B.n56 585
R46 B.n501 B.n500 585
R47 B.n502 B.n55 585
R48 B.n504 B.n503 585
R49 B.n505 B.n54 585
R50 B.n507 B.n506 585
R51 B.n508 B.n53 585
R52 B.n510 B.n509 585
R53 B.n511 B.n52 585
R54 B.n513 B.n512 585
R55 B.n514 B.n51 585
R56 B.n516 B.n515 585
R57 B.n517 B.n50 585
R58 B.n519 B.n518 585
R59 B.n520 B.n49 585
R60 B.n522 B.n521 585
R61 B.n524 B.n523 585
R62 B.n525 B.n45 585
R63 B.n527 B.n526 585
R64 B.n528 B.n44 585
R65 B.n530 B.n529 585
R66 B.n531 B.n43 585
R67 B.n533 B.n532 585
R68 B.n534 B.n42 585
R69 B.n536 B.n535 585
R70 B.n538 B.n39 585
R71 B.n540 B.n539 585
R72 B.n541 B.n38 585
R73 B.n543 B.n542 585
R74 B.n544 B.n37 585
R75 B.n546 B.n545 585
R76 B.n547 B.n36 585
R77 B.n549 B.n548 585
R78 B.n550 B.n35 585
R79 B.n552 B.n551 585
R80 B.n553 B.n34 585
R81 B.n555 B.n554 585
R82 B.n556 B.n33 585
R83 B.n558 B.n557 585
R84 B.n559 B.n32 585
R85 B.n561 B.n560 585
R86 B.n562 B.n31 585
R87 B.n564 B.n563 585
R88 B.n565 B.n30 585
R89 B.n567 B.n566 585
R90 B.n568 B.n29 585
R91 B.n570 B.n569 585
R92 B.n571 B.n28 585
R93 B.n573 B.n572 585
R94 B.n574 B.n27 585
R95 B.n576 B.n575 585
R96 B.n577 B.n26 585
R97 B.n579 B.n578 585
R98 B.n580 B.n25 585
R99 B.n582 B.n581 585
R100 B.n583 B.n24 585
R101 B.n585 B.n584 585
R102 B.n586 B.n23 585
R103 B.n588 B.n587 585
R104 B.n589 B.n22 585
R105 B.n591 B.n590 585
R106 B.n592 B.n21 585
R107 B.n594 B.n593 585
R108 B.n595 B.n20 585
R109 B.n597 B.n596 585
R110 B.n598 B.n19 585
R111 B.n600 B.n599 585
R112 B.n601 B.n18 585
R113 B.n603 B.n602 585
R114 B.n604 B.n17 585
R115 B.n606 B.n605 585
R116 B.n607 B.n16 585
R117 B.n609 B.n608 585
R118 B.n610 B.n15 585
R119 B.n612 B.n611 585
R120 B.n613 B.n14 585
R121 B.n615 B.n614 585
R122 B.n616 B.n13 585
R123 B.n618 B.n617 585
R124 B.n619 B.n12 585
R125 B.n621 B.n620 585
R126 B.n622 B.n11 585
R127 B.n436 B.n77 585
R128 B.n435 B.n434 585
R129 B.n433 B.n78 585
R130 B.n432 B.n431 585
R131 B.n430 B.n79 585
R132 B.n429 B.n428 585
R133 B.n427 B.n80 585
R134 B.n426 B.n425 585
R135 B.n424 B.n81 585
R136 B.n423 B.n422 585
R137 B.n421 B.n82 585
R138 B.n420 B.n419 585
R139 B.n418 B.n83 585
R140 B.n417 B.n416 585
R141 B.n415 B.n84 585
R142 B.n414 B.n413 585
R143 B.n412 B.n85 585
R144 B.n411 B.n410 585
R145 B.n409 B.n86 585
R146 B.n408 B.n407 585
R147 B.n406 B.n87 585
R148 B.n405 B.n404 585
R149 B.n403 B.n88 585
R150 B.n402 B.n401 585
R151 B.n400 B.n89 585
R152 B.n399 B.n398 585
R153 B.n397 B.n90 585
R154 B.n396 B.n395 585
R155 B.n394 B.n91 585
R156 B.n393 B.n392 585
R157 B.n391 B.n92 585
R158 B.n390 B.n389 585
R159 B.n388 B.n93 585
R160 B.n387 B.n386 585
R161 B.n385 B.n94 585
R162 B.n384 B.n383 585
R163 B.n382 B.n95 585
R164 B.n196 B.n161 585
R165 B.n198 B.n197 585
R166 B.n199 B.n160 585
R167 B.n201 B.n200 585
R168 B.n202 B.n159 585
R169 B.n204 B.n203 585
R170 B.n205 B.n158 585
R171 B.n207 B.n206 585
R172 B.n208 B.n157 585
R173 B.n210 B.n209 585
R174 B.n211 B.n156 585
R175 B.n213 B.n212 585
R176 B.n214 B.n155 585
R177 B.n216 B.n215 585
R178 B.n217 B.n154 585
R179 B.n219 B.n218 585
R180 B.n220 B.n153 585
R181 B.n222 B.n221 585
R182 B.n223 B.n152 585
R183 B.n225 B.n224 585
R184 B.n226 B.n151 585
R185 B.n228 B.n227 585
R186 B.n229 B.n150 585
R187 B.n231 B.n230 585
R188 B.n232 B.n149 585
R189 B.n234 B.n233 585
R190 B.n235 B.n148 585
R191 B.n237 B.n236 585
R192 B.n238 B.n147 585
R193 B.n240 B.n239 585
R194 B.n241 B.n146 585
R195 B.n243 B.n242 585
R196 B.n244 B.n145 585
R197 B.n246 B.n245 585
R198 B.n247 B.n144 585
R199 B.n249 B.n248 585
R200 B.n250 B.n143 585
R201 B.n252 B.n251 585
R202 B.n253 B.n142 585
R203 B.n255 B.n254 585
R204 B.n256 B.n141 585
R205 B.n258 B.n257 585
R206 B.n259 B.n140 585
R207 B.n261 B.n260 585
R208 B.n262 B.n139 585
R209 B.n264 B.n263 585
R210 B.n265 B.n138 585
R211 B.n267 B.n266 585
R212 B.n268 B.n137 585
R213 B.n270 B.n269 585
R214 B.n271 B.n136 585
R215 B.n273 B.n272 585
R216 B.n274 B.n135 585
R217 B.n276 B.n275 585
R218 B.n277 B.n134 585
R219 B.n279 B.n278 585
R220 B.n280 B.n131 585
R221 B.n283 B.n282 585
R222 B.n284 B.n130 585
R223 B.n286 B.n285 585
R224 B.n287 B.n129 585
R225 B.n289 B.n288 585
R226 B.n290 B.n128 585
R227 B.n292 B.n291 585
R228 B.n293 B.n127 585
R229 B.n295 B.n294 585
R230 B.n297 B.n296 585
R231 B.n298 B.n123 585
R232 B.n300 B.n299 585
R233 B.n301 B.n122 585
R234 B.n303 B.n302 585
R235 B.n304 B.n121 585
R236 B.n306 B.n305 585
R237 B.n307 B.n120 585
R238 B.n309 B.n308 585
R239 B.n310 B.n119 585
R240 B.n312 B.n311 585
R241 B.n313 B.n118 585
R242 B.n315 B.n314 585
R243 B.n316 B.n117 585
R244 B.n318 B.n317 585
R245 B.n319 B.n116 585
R246 B.n321 B.n320 585
R247 B.n322 B.n115 585
R248 B.n324 B.n323 585
R249 B.n325 B.n114 585
R250 B.n327 B.n326 585
R251 B.n328 B.n113 585
R252 B.n330 B.n329 585
R253 B.n331 B.n112 585
R254 B.n333 B.n332 585
R255 B.n334 B.n111 585
R256 B.n336 B.n335 585
R257 B.n337 B.n110 585
R258 B.n339 B.n338 585
R259 B.n340 B.n109 585
R260 B.n342 B.n341 585
R261 B.n343 B.n108 585
R262 B.n345 B.n344 585
R263 B.n346 B.n107 585
R264 B.n348 B.n347 585
R265 B.n349 B.n106 585
R266 B.n351 B.n350 585
R267 B.n352 B.n105 585
R268 B.n354 B.n353 585
R269 B.n355 B.n104 585
R270 B.n357 B.n356 585
R271 B.n358 B.n103 585
R272 B.n360 B.n359 585
R273 B.n361 B.n102 585
R274 B.n363 B.n362 585
R275 B.n364 B.n101 585
R276 B.n366 B.n365 585
R277 B.n367 B.n100 585
R278 B.n369 B.n368 585
R279 B.n370 B.n99 585
R280 B.n372 B.n371 585
R281 B.n373 B.n98 585
R282 B.n375 B.n374 585
R283 B.n376 B.n97 585
R284 B.n378 B.n377 585
R285 B.n379 B.n96 585
R286 B.n381 B.n380 585
R287 B.n195 B.n194 585
R288 B.n193 B.n162 585
R289 B.n192 B.n191 585
R290 B.n190 B.n163 585
R291 B.n189 B.n188 585
R292 B.n187 B.n164 585
R293 B.n186 B.n185 585
R294 B.n184 B.n165 585
R295 B.n183 B.n182 585
R296 B.n181 B.n166 585
R297 B.n180 B.n179 585
R298 B.n178 B.n167 585
R299 B.n177 B.n176 585
R300 B.n175 B.n168 585
R301 B.n174 B.n173 585
R302 B.n172 B.n169 585
R303 B.n171 B.n170 585
R304 B.n2 B.n0 585
R305 B.n649 B.n1 585
R306 B.n648 B.n647 585
R307 B.n646 B.n3 585
R308 B.n645 B.n644 585
R309 B.n643 B.n4 585
R310 B.n642 B.n641 585
R311 B.n640 B.n5 585
R312 B.n639 B.n638 585
R313 B.n637 B.n6 585
R314 B.n636 B.n635 585
R315 B.n634 B.n7 585
R316 B.n633 B.n632 585
R317 B.n631 B.n8 585
R318 B.n630 B.n629 585
R319 B.n628 B.n9 585
R320 B.n627 B.n626 585
R321 B.n625 B.n10 585
R322 B.n624 B.n623 585
R323 B.n651 B.n650 585
R324 B.n194 B.n161 473.281
R325 B.n624 B.n11 473.281
R326 B.n380 B.n95 473.281
R327 B.n438 B.n77 473.281
R328 B.n194 B.n193 163.367
R329 B.n193 B.n192 163.367
R330 B.n192 B.n163 163.367
R331 B.n188 B.n163 163.367
R332 B.n188 B.n187 163.367
R333 B.n187 B.n186 163.367
R334 B.n186 B.n165 163.367
R335 B.n182 B.n165 163.367
R336 B.n182 B.n181 163.367
R337 B.n181 B.n180 163.367
R338 B.n180 B.n167 163.367
R339 B.n176 B.n167 163.367
R340 B.n176 B.n175 163.367
R341 B.n175 B.n174 163.367
R342 B.n174 B.n169 163.367
R343 B.n170 B.n169 163.367
R344 B.n170 B.n2 163.367
R345 B.n650 B.n2 163.367
R346 B.n650 B.n649 163.367
R347 B.n649 B.n648 163.367
R348 B.n648 B.n3 163.367
R349 B.n644 B.n3 163.367
R350 B.n644 B.n643 163.367
R351 B.n643 B.n642 163.367
R352 B.n642 B.n5 163.367
R353 B.n638 B.n5 163.367
R354 B.n638 B.n637 163.367
R355 B.n637 B.n636 163.367
R356 B.n636 B.n7 163.367
R357 B.n632 B.n7 163.367
R358 B.n632 B.n631 163.367
R359 B.n631 B.n630 163.367
R360 B.n630 B.n9 163.367
R361 B.n626 B.n9 163.367
R362 B.n626 B.n625 163.367
R363 B.n625 B.n624 163.367
R364 B.n198 B.n161 163.367
R365 B.n199 B.n198 163.367
R366 B.n200 B.n199 163.367
R367 B.n200 B.n159 163.367
R368 B.n204 B.n159 163.367
R369 B.n205 B.n204 163.367
R370 B.n206 B.n205 163.367
R371 B.n206 B.n157 163.367
R372 B.n210 B.n157 163.367
R373 B.n211 B.n210 163.367
R374 B.n212 B.n211 163.367
R375 B.n212 B.n155 163.367
R376 B.n216 B.n155 163.367
R377 B.n217 B.n216 163.367
R378 B.n218 B.n217 163.367
R379 B.n218 B.n153 163.367
R380 B.n222 B.n153 163.367
R381 B.n223 B.n222 163.367
R382 B.n224 B.n223 163.367
R383 B.n224 B.n151 163.367
R384 B.n228 B.n151 163.367
R385 B.n229 B.n228 163.367
R386 B.n230 B.n229 163.367
R387 B.n230 B.n149 163.367
R388 B.n234 B.n149 163.367
R389 B.n235 B.n234 163.367
R390 B.n236 B.n235 163.367
R391 B.n236 B.n147 163.367
R392 B.n240 B.n147 163.367
R393 B.n241 B.n240 163.367
R394 B.n242 B.n241 163.367
R395 B.n242 B.n145 163.367
R396 B.n246 B.n145 163.367
R397 B.n247 B.n246 163.367
R398 B.n248 B.n247 163.367
R399 B.n248 B.n143 163.367
R400 B.n252 B.n143 163.367
R401 B.n253 B.n252 163.367
R402 B.n254 B.n253 163.367
R403 B.n254 B.n141 163.367
R404 B.n258 B.n141 163.367
R405 B.n259 B.n258 163.367
R406 B.n260 B.n259 163.367
R407 B.n260 B.n139 163.367
R408 B.n264 B.n139 163.367
R409 B.n265 B.n264 163.367
R410 B.n266 B.n265 163.367
R411 B.n266 B.n137 163.367
R412 B.n270 B.n137 163.367
R413 B.n271 B.n270 163.367
R414 B.n272 B.n271 163.367
R415 B.n272 B.n135 163.367
R416 B.n276 B.n135 163.367
R417 B.n277 B.n276 163.367
R418 B.n278 B.n277 163.367
R419 B.n278 B.n131 163.367
R420 B.n283 B.n131 163.367
R421 B.n284 B.n283 163.367
R422 B.n285 B.n284 163.367
R423 B.n285 B.n129 163.367
R424 B.n289 B.n129 163.367
R425 B.n290 B.n289 163.367
R426 B.n291 B.n290 163.367
R427 B.n291 B.n127 163.367
R428 B.n295 B.n127 163.367
R429 B.n296 B.n295 163.367
R430 B.n296 B.n123 163.367
R431 B.n300 B.n123 163.367
R432 B.n301 B.n300 163.367
R433 B.n302 B.n301 163.367
R434 B.n302 B.n121 163.367
R435 B.n306 B.n121 163.367
R436 B.n307 B.n306 163.367
R437 B.n308 B.n307 163.367
R438 B.n308 B.n119 163.367
R439 B.n312 B.n119 163.367
R440 B.n313 B.n312 163.367
R441 B.n314 B.n313 163.367
R442 B.n314 B.n117 163.367
R443 B.n318 B.n117 163.367
R444 B.n319 B.n318 163.367
R445 B.n320 B.n319 163.367
R446 B.n320 B.n115 163.367
R447 B.n324 B.n115 163.367
R448 B.n325 B.n324 163.367
R449 B.n326 B.n325 163.367
R450 B.n326 B.n113 163.367
R451 B.n330 B.n113 163.367
R452 B.n331 B.n330 163.367
R453 B.n332 B.n331 163.367
R454 B.n332 B.n111 163.367
R455 B.n336 B.n111 163.367
R456 B.n337 B.n336 163.367
R457 B.n338 B.n337 163.367
R458 B.n338 B.n109 163.367
R459 B.n342 B.n109 163.367
R460 B.n343 B.n342 163.367
R461 B.n344 B.n343 163.367
R462 B.n344 B.n107 163.367
R463 B.n348 B.n107 163.367
R464 B.n349 B.n348 163.367
R465 B.n350 B.n349 163.367
R466 B.n350 B.n105 163.367
R467 B.n354 B.n105 163.367
R468 B.n355 B.n354 163.367
R469 B.n356 B.n355 163.367
R470 B.n356 B.n103 163.367
R471 B.n360 B.n103 163.367
R472 B.n361 B.n360 163.367
R473 B.n362 B.n361 163.367
R474 B.n362 B.n101 163.367
R475 B.n366 B.n101 163.367
R476 B.n367 B.n366 163.367
R477 B.n368 B.n367 163.367
R478 B.n368 B.n99 163.367
R479 B.n372 B.n99 163.367
R480 B.n373 B.n372 163.367
R481 B.n374 B.n373 163.367
R482 B.n374 B.n97 163.367
R483 B.n378 B.n97 163.367
R484 B.n379 B.n378 163.367
R485 B.n380 B.n379 163.367
R486 B.n384 B.n95 163.367
R487 B.n385 B.n384 163.367
R488 B.n386 B.n385 163.367
R489 B.n386 B.n93 163.367
R490 B.n390 B.n93 163.367
R491 B.n391 B.n390 163.367
R492 B.n392 B.n391 163.367
R493 B.n392 B.n91 163.367
R494 B.n396 B.n91 163.367
R495 B.n397 B.n396 163.367
R496 B.n398 B.n397 163.367
R497 B.n398 B.n89 163.367
R498 B.n402 B.n89 163.367
R499 B.n403 B.n402 163.367
R500 B.n404 B.n403 163.367
R501 B.n404 B.n87 163.367
R502 B.n408 B.n87 163.367
R503 B.n409 B.n408 163.367
R504 B.n410 B.n409 163.367
R505 B.n410 B.n85 163.367
R506 B.n414 B.n85 163.367
R507 B.n415 B.n414 163.367
R508 B.n416 B.n415 163.367
R509 B.n416 B.n83 163.367
R510 B.n420 B.n83 163.367
R511 B.n421 B.n420 163.367
R512 B.n422 B.n421 163.367
R513 B.n422 B.n81 163.367
R514 B.n426 B.n81 163.367
R515 B.n427 B.n426 163.367
R516 B.n428 B.n427 163.367
R517 B.n428 B.n79 163.367
R518 B.n432 B.n79 163.367
R519 B.n433 B.n432 163.367
R520 B.n434 B.n433 163.367
R521 B.n434 B.n77 163.367
R522 B.n620 B.n11 163.367
R523 B.n620 B.n619 163.367
R524 B.n619 B.n618 163.367
R525 B.n618 B.n13 163.367
R526 B.n614 B.n13 163.367
R527 B.n614 B.n613 163.367
R528 B.n613 B.n612 163.367
R529 B.n612 B.n15 163.367
R530 B.n608 B.n15 163.367
R531 B.n608 B.n607 163.367
R532 B.n607 B.n606 163.367
R533 B.n606 B.n17 163.367
R534 B.n602 B.n17 163.367
R535 B.n602 B.n601 163.367
R536 B.n601 B.n600 163.367
R537 B.n600 B.n19 163.367
R538 B.n596 B.n19 163.367
R539 B.n596 B.n595 163.367
R540 B.n595 B.n594 163.367
R541 B.n594 B.n21 163.367
R542 B.n590 B.n21 163.367
R543 B.n590 B.n589 163.367
R544 B.n589 B.n588 163.367
R545 B.n588 B.n23 163.367
R546 B.n584 B.n23 163.367
R547 B.n584 B.n583 163.367
R548 B.n583 B.n582 163.367
R549 B.n582 B.n25 163.367
R550 B.n578 B.n25 163.367
R551 B.n578 B.n577 163.367
R552 B.n577 B.n576 163.367
R553 B.n576 B.n27 163.367
R554 B.n572 B.n27 163.367
R555 B.n572 B.n571 163.367
R556 B.n571 B.n570 163.367
R557 B.n570 B.n29 163.367
R558 B.n566 B.n29 163.367
R559 B.n566 B.n565 163.367
R560 B.n565 B.n564 163.367
R561 B.n564 B.n31 163.367
R562 B.n560 B.n31 163.367
R563 B.n560 B.n559 163.367
R564 B.n559 B.n558 163.367
R565 B.n558 B.n33 163.367
R566 B.n554 B.n33 163.367
R567 B.n554 B.n553 163.367
R568 B.n553 B.n552 163.367
R569 B.n552 B.n35 163.367
R570 B.n548 B.n35 163.367
R571 B.n548 B.n547 163.367
R572 B.n547 B.n546 163.367
R573 B.n546 B.n37 163.367
R574 B.n542 B.n37 163.367
R575 B.n542 B.n541 163.367
R576 B.n541 B.n540 163.367
R577 B.n540 B.n39 163.367
R578 B.n535 B.n39 163.367
R579 B.n535 B.n534 163.367
R580 B.n534 B.n533 163.367
R581 B.n533 B.n43 163.367
R582 B.n529 B.n43 163.367
R583 B.n529 B.n528 163.367
R584 B.n528 B.n527 163.367
R585 B.n527 B.n45 163.367
R586 B.n523 B.n45 163.367
R587 B.n523 B.n522 163.367
R588 B.n522 B.n49 163.367
R589 B.n518 B.n49 163.367
R590 B.n518 B.n517 163.367
R591 B.n517 B.n516 163.367
R592 B.n516 B.n51 163.367
R593 B.n512 B.n51 163.367
R594 B.n512 B.n511 163.367
R595 B.n511 B.n510 163.367
R596 B.n510 B.n53 163.367
R597 B.n506 B.n53 163.367
R598 B.n506 B.n505 163.367
R599 B.n505 B.n504 163.367
R600 B.n504 B.n55 163.367
R601 B.n500 B.n55 163.367
R602 B.n500 B.n499 163.367
R603 B.n499 B.n498 163.367
R604 B.n498 B.n57 163.367
R605 B.n494 B.n57 163.367
R606 B.n494 B.n493 163.367
R607 B.n493 B.n492 163.367
R608 B.n492 B.n59 163.367
R609 B.n488 B.n59 163.367
R610 B.n488 B.n487 163.367
R611 B.n487 B.n486 163.367
R612 B.n486 B.n61 163.367
R613 B.n482 B.n61 163.367
R614 B.n482 B.n481 163.367
R615 B.n481 B.n480 163.367
R616 B.n480 B.n63 163.367
R617 B.n476 B.n63 163.367
R618 B.n476 B.n475 163.367
R619 B.n475 B.n474 163.367
R620 B.n474 B.n65 163.367
R621 B.n470 B.n65 163.367
R622 B.n470 B.n469 163.367
R623 B.n469 B.n468 163.367
R624 B.n468 B.n67 163.367
R625 B.n464 B.n67 163.367
R626 B.n464 B.n463 163.367
R627 B.n463 B.n462 163.367
R628 B.n462 B.n69 163.367
R629 B.n458 B.n69 163.367
R630 B.n458 B.n457 163.367
R631 B.n457 B.n456 163.367
R632 B.n456 B.n71 163.367
R633 B.n452 B.n71 163.367
R634 B.n452 B.n451 163.367
R635 B.n451 B.n450 163.367
R636 B.n450 B.n73 163.367
R637 B.n446 B.n73 163.367
R638 B.n446 B.n445 163.367
R639 B.n445 B.n444 163.367
R640 B.n444 B.n75 163.367
R641 B.n440 B.n75 163.367
R642 B.n440 B.n439 163.367
R643 B.n439 B.n438 163.367
R644 B.n124 B.t8 119.675
R645 B.n46 B.t1 119.675
R646 B.n132 B.t5 119.653
R647 B.n40 B.t10 119.653
R648 B.n125 B.t7 109.008
R649 B.n47 B.t2 109.008
R650 B.n133 B.t4 108.987
R651 B.n41 B.t11 108.987
R652 B.n126 B.n125 59.5399
R653 B.n281 B.n133 59.5399
R654 B.n537 B.n41 59.5399
R655 B.n48 B.n47 59.5399
R656 B.n623 B.n622 30.7517
R657 B.n382 B.n381 30.7517
R658 B.n196 B.n195 30.7517
R659 B.n437 B.n436 30.7517
R660 B B.n651 18.0485
R661 B.n125 B.n124 10.6672
R662 B.n133 B.n132 10.6672
R663 B.n41 B.n40 10.6672
R664 B.n47 B.n46 10.6672
R665 B.n622 B.n621 10.6151
R666 B.n621 B.n12 10.6151
R667 B.n617 B.n12 10.6151
R668 B.n617 B.n616 10.6151
R669 B.n616 B.n615 10.6151
R670 B.n615 B.n14 10.6151
R671 B.n611 B.n14 10.6151
R672 B.n611 B.n610 10.6151
R673 B.n610 B.n609 10.6151
R674 B.n609 B.n16 10.6151
R675 B.n605 B.n16 10.6151
R676 B.n605 B.n604 10.6151
R677 B.n604 B.n603 10.6151
R678 B.n603 B.n18 10.6151
R679 B.n599 B.n18 10.6151
R680 B.n599 B.n598 10.6151
R681 B.n598 B.n597 10.6151
R682 B.n597 B.n20 10.6151
R683 B.n593 B.n20 10.6151
R684 B.n593 B.n592 10.6151
R685 B.n592 B.n591 10.6151
R686 B.n591 B.n22 10.6151
R687 B.n587 B.n22 10.6151
R688 B.n587 B.n586 10.6151
R689 B.n586 B.n585 10.6151
R690 B.n585 B.n24 10.6151
R691 B.n581 B.n24 10.6151
R692 B.n581 B.n580 10.6151
R693 B.n580 B.n579 10.6151
R694 B.n579 B.n26 10.6151
R695 B.n575 B.n26 10.6151
R696 B.n575 B.n574 10.6151
R697 B.n574 B.n573 10.6151
R698 B.n573 B.n28 10.6151
R699 B.n569 B.n28 10.6151
R700 B.n569 B.n568 10.6151
R701 B.n568 B.n567 10.6151
R702 B.n567 B.n30 10.6151
R703 B.n563 B.n30 10.6151
R704 B.n563 B.n562 10.6151
R705 B.n562 B.n561 10.6151
R706 B.n561 B.n32 10.6151
R707 B.n557 B.n32 10.6151
R708 B.n557 B.n556 10.6151
R709 B.n556 B.n555 10.6151
R710 B.n555 B.n34 10.6151
R711 B.n551 B.n34 10.6151
R712 B.n551 B.n550 10.6151
R713 B.n550 B.n549 10.6151
R714 B.n549 B.n36 10.6151
R715 B.n545 B.n36 10.6151
R716 B.n545 B.n544 10.6151
R717 B.n544 B.n543 10.6151
R718 B.n543 B.n38 10.6151
R719 B.n539 B.n38 10.6151
R720 B.n539 B.n538 10.6151
R721 B.n536 B.n42 10.6151
R722 B.n532 B.n42 10.6151
R723 B.n532 B.n531 10.6151
R724 B.n531 B.n530 10.6151
R725 B.n530 B.n44 10.6151
R726 B.n526 B.n44 10.6151
R727 B.n526 B.n525 10.6151
R728 B.n525 B.n524 10.6151
R729 B.n521 B.n520 10.6151
R730 B.n520 B.n519 10.6151
R731 B.n519 B.n50 10.6151
R732 B.n515 B.n50 10.6151
R733 B.n515 B.n514 10.6151
R734 B.n514 B.n513 10.6151
R735 B.n513 B.n52 10.6151
R736 B.n509 B.n52 10.6151
R737 B.n509 B.n508 10.6151
R738 B.n508 B.n507 10.6151
R739 B.n507 B.n54 10.6151
R740 B.n503 B.n54 10.6151
R741 B.n503 B.n502 10.6151
R742 B.n502 B.n501 10.6151
R743 B.n501 B.n56 10.6151
R744 B.n497 B.n56 10.6151
R745 B.n497 B.n496 10.6151
R746 B.n496 B.n495 10.6151
R747 B.n495 B.n58 10.6151
R748 B.n491 B.n58 10.6151
R749 B.n491 B.n490 10.6151
R750 B.n490 B.n489 10.6151
R751 B.n489 B.n60 10.6151
R752 B.n485 B.n60 10.6151
R753 B.n485 B.n484 10.6151
R754 B.n484 B.n483 10.6151
R755 B.n483 B.n62 10.6151
R756 B.n479 B.n62 10.6151
R757 B.n479 B.n478 10.6151
R758 B.n478 B.n477 10.6151
R759 B.n477 B.n64 10.6151
R760 B.n473 B.n64 10.6151
R761 B.n473 B.n472 10.6151
R762 B.n472 B.n471 10.6151
R763 B.n471 B.n66 10.6151
R764 B.n467 B.n66 10.6151
R765 B.n467 B.n466 10.6151
R766 B.n466 B.n465 10.6151
R767 B.n465 B.n68 10.6151
R768 B.n461 B.n68 10.6151
R769 B.n461 B.n460 10.6151
R770 B.n460 B.n459 10.6151
R771 B.n459 B.n70 10.6151
R772 B.n455 B.n70 10.6151
R773 B.n455 B.n454 10.6151
R774 B.n454 B.n453 10.6151
R775 B.n453 B.n72 10.6151
R776 B.n449 B.n72 10.6151
R777 B.n449 B.n448 10.6151
R778 B.n448 B.n447 10.6151
R779 B.n447 B.n74 10.6151
R780 B.n443 B.n74 10.6151
R781 B.n443 B.n442 10.6151
R782 B.n442 B.n441 10.6151
R783 B.n441 B.n76 10.6151
R784 B.n437 B.n76 10.6151
R785 B.n383 B.n382 10.6151
R786 B.n383 B.n94 10.6151
R787 B.n387 B.n94 10.6151
R788 B.n388 B.n387 10.6151
R789 B.n389 B.n388 10.6151
R790 B.n389 B.n92 10.6151
R791 B.n393 B.n92 10.6151
R792 B.n394 B.n393 10.6151
R793 B.n395 B.n394 10.6151
R794 B.n395 B.n90 10.6151
R795 B.n399 B.n90 10.6151
R796 B.n400 B.n399 10.6151
R797 B.n401 B.n400 10.6151
R798 B.n401 B.n88 10.6151
R799 B.n405 B.n88 10.6151
R800 B.n406 B.n405 10.6151
R801 B.n407 B.n406 10.6151
R802 B.n407 B.n86 10.6151
R803 B.n411 B.n86 10.6151
R804 B.n412 B.n411 10.6151
R805 B.n413 B.n412 10.6151
R806 B.n413 B.n84 10.6151
R807 B.n417 B.n84 10.6151
R808 B.n418 B.n417 10.6151
R809 B.n419 B.n418 10.6151
R810 B.n419 B.n82 10.6151
R811 B.n423 B.n82 10.6151
R812 B.n424 B.n423 10.6151
R813 B.n425 B.n424 10.6151
R814 B.n425 B.n80 10.6151
R815 B.n429 B.n80 10.6151
R816 B.n430 B.n429 10.6151
R817 B.n431 B.n430 10.6151
R818 B.n431 B.n78 10.6151
R819 B.n435 B.n78 10.6151
R820 B.n436 B.n435 10.6151
R821 B.n197 B.n196 10.6151
R822 B.n197 B.n160 10.6151
R823 B.n201 B.n160 10.6151
R824 B.n202 B.n201 10.6151
R825 B.n203 B.n202 10.6151
R826 B.n203 B.n158 10.6151
R827 B.n207 B.n158 10.6151
R828 B.n208 B.n207 10.6151
R829 B.n209 B.n208 10.6151
R830 B.n209 B.n156 10.6151
R831 B.n213 B.n156 10.6151
R832 B.n214 B.n213 10.6151
R833 B.n215 B.n214 10.6151
R834 B.n215 B.n154 10.6151
R835 B.n219 B.n154 10.6151
R836 B.n220 B.n219 10.6151
R837 B.n221 B.n220 10.6151
R838 B.n221 B.n152 10.6151
R839 B.n225 B.n152 10.6151
R840 B.n226 B.n225 10.6151
R841 B.n227 B.n226 10.6151
R842 B.n227 B.n150 10.6151
R843 B.n231 B.n150 10.6151
R844 B.n232 B.n231 10.6151
R845 B.n233 B.n232 10.6151
R846 B.n233 B.n148 10.6151
R847 B.n237 B.n148 10.6151
R848 B.n238 B.n237 10.6151
R849 B.n239 B.n238 10.6151
R850 B.n239 B.n146 10.6151
R851 B.n243 B.n146 10.6151
R852 B.n244 B.n243 10.6151
R853 B.n245 B.n244 10.6151
R854 B.n245 B.n144 10.6151
R855 B.n249 B.n144 10.6151
R856 B.n250 B.n249 10.6151
R857 B.n251 B.n250 10.6151
R858 B.n251 B.n142 10.6151
R859 B.n255 B.n142 10.6151
R860 B.n256 B.n255 10.6151
R861 B.n257 B.n256 10.6151
R862 B.n257 B.n140 10.6151
R863 B.n261 B.n140 10.6151
R864 B.n262 B.n261 10.6151
R865 B.n263 B.n262 10.6151
R866 B.n263 B.n138 10.6151
R867 B.n267 B.n138 10.6151
R868 B.n268 B.n267 10.6151
R869 B.n269 B.n268 10.6151
R870 B.n269 B.n136 10.6151
R871 B.n273 B.n136 10.6151
R872 B.n274 B.n273 10.6151
R873 B.n275 B.n274 10.6151
R874 B.n275 B.n134 10.6151
R875 B.n279 B.n134 10.6151
R876 B.n280 B.n279 10.6151
R877 B.n282 B.n130 10.6151
R878 B.n286 B.n130 10.6151
R879 B.n287 B.n286 10.6151
R880 B.n288 B.n287 10.6151
R881 B.n288 B.n128 10.6151
R882 B.n292 B.n128 10.6151
R883 B.n293 B.n292 10.6151
R884 B.n294 B.n293 10.6151
R885 B.n298 B.n297 10.6151
R886 B.n299 B.n298 10.6151
R887 B.n299 B.n122 10.6151
R888 B.n303 B.n122 10.6151
R889 B.n304 B.n303 10.6151
R890 B.n305 B.n304 10.6151
R891 B.n305 B.n120 10.6151
R892 B.n309 B.n120 10.6151
R893 B.n310 B.n309 10.6151
R894 B.n311 B.n310 10.6151
R895 B.n311 B.n118 10.6151
R896 B.n315 B.n118 10.6151
R897 B.n316 B.n315 10.6151
R898 B.n317 B.n316 10.6151
R899 B.n317 B.n116 10.6151
R900 B.n321 B.n116 10.6151
R901 B.n322 B.n321 10.6151
R902 B.n323 B.n322 10.6151
R903 B.n323 B.n114 10.6151
R904 B.n327 B.n114 10.6151
R905 B.n328 B.n327 10.6151
R906 B.n329 B.n328 10.6151
R907 B.n329 B.n112 10.6151
R908 B.n333 B.n112 10.6151
R909 B.n334 B.n333 10.6151
R910 B.n335 B.n334 10.6151
R911 B.n335 B.n110 10.6151
R912 B.n339 B.n110 10.6151
R913 B.n340 B.n339 10.6151
R914 B.n341 B.n340 10.6151
R915 B.n341 B.n108 10.6151
R916 B.n345 B.n108 10.6151
R917 B.n346 B.n345 10.6151
R918 B.n347 B.n346 10.6151
R919 B.n347 B.n106 10.6151
R920 B.n351 B.n106 10.6151
R921 B.n352 B.n351 10.6151
R922 B.n353 B.n352 10.6151
R923 B.n353 B.n104 10.6151
R924 B.n357 B.n104 10.6151
R925 B.n358 B.n357 10.6151
R926 B.n359 B.n358 10.6151
R927 B.n359 B.n102 10.6151
R928 B.n363 B.n102 10.6151
R929 B.n364 B.n363 10.6151
R930 B.n365 B.n364 10.6151
R931 B.n365 B.n100 10.6151
R932 B.n369 B.n100 10.6151
R933 B.n370 B.n369 10.6151
R934 B.n371 B.n370 10.6151
R935 B.n371 B.n98 10.6151
R936 B.n375 B.n98 10.6151
R937 B.n376 B.n375 10.6151
R938 B.n377 B.n376 10.6151
R939 B.n377 B.n96 10.6151
R940 B.n381 B.n96 10.6151
R941 B.n195 B.n162 10.6151
R942 B.n191 B.n162 10.6151
R943 B.n191 B.n190 10.6151
R944 B.n190 B.n189 10.6151
R945 B.n189 B.n164 10.6151
R946 B.n185 B.n164 10.6151
R947 B.n185 B.n184 10.6151
R948 B.n184 B.n183 10.6151
R949 B.n183 B.n166 10.6151
R950 B.n179 B.n166 10.6151
R951 B.n179 B.n178 10.6151
R952 B.n178 B.n177 10.6151
R953 B.n177 B.n168 10.6151
R954 B.n173 B.n168 10.6151
R955 B.n173 B.n172 10.6151
R956 B.n172 B.n171 10.6151
R957 B.n171 B.n0 10.6151
R958 B.n647 B.n1 10.6151
R959 B.n647 B.n646 10.6151
R960 B.n646 B.n645 10.6151
R961 B.n645 B.n4 10.6151
R962 B.n641 B.n4 10.6151
R963 B.n641 B.n640 10.6151
R964 B.n640 B.n639 10.6151
R965 B.n639 B.n6 10.6151
R966 B.n635 B.n6 10.6151
R967 B.n635 B.n634 10.6151
R968 B.n634 B.n633 10.6151
R969 B.n633 B.n8 10.6151
R970 B.n629 B.n8 10.6151
R971 B.n629 B.n628 10.6151
R972 B.n628 B.n627 10.6151
R973 B.n627 B.n10 10.6151
R974 B.n623 B.n10 10.6151
R975 B.n537 B.n536 6.5566
R976 B.n524 B.n48 6.5566
R977 B.n282 B.n281 6.5566
R978 B.n294 B.n126 6.5566
R979 B.n538 B.n537 4.05904
R980 B.n521 B.n48 4.05904
R981 B.n281 B.n280 4.05904
R982 B.n297 B.n126 4.05904
R983 B.n651 B.n0 2.81026
R984 B.n651 B.n1 2.81026
R985 VP.n19 VP.t8 2071.14
R986 VP.n12 VP.t6 2071.14
R987 VP.n4 VP.t0 2071.14
R988 VP.n10 VP.t1 2071.14
R989 VP.n18 VP.t5 2020.02
R990 VP.n16 VP.t2 2020.02
R991 VP.n1 VP.t9 2020.02
R992 VP.n3 VP.t4 2020.02
R993 VP.n7 VP.t3 2020.02
R994 VP.n9 VP.t7 2020.02
R995 VP.n5 VP.n4 161.489
R996 VP.n20 VP.n19 161.3
R997 VP.n6 VP.n5 161.3
R998 VP.n8 VP.n2 161.3
R999 VP.n11 VP.n10 161.3
R1000 VP.n17 VP.n0 161.3
R1001 VP.n15 VP.n14 161.3
R1002 VP.n13 VP.n12 161.3
R1003 VP.n13 VP.n11 44.171
R1004 VP.n15 VP.n1 43.8187
R1005 VP.n18 VP.n17 43.8187
R1006 VP.n6 VP.n3 43.8187
R1007 VP.n9 VP.n8 43.8187
R1008 VP.n16 VP.n15 36.5157
R1009 VP.n17 VP.n16 36.5157
R1010 VP.n7 VP.n6 36.5157
R1011 VP.n8 VP.n7 36.5157
R1012 VP.n12 VP.n1 29.2126
R1013 VP.n19 VP.n18 29.2126
R1014 VP.n4 VP.n3 29.2126
R1015 VP.n10 VP.n9 29.2126
R1016 VP.n5 VP.n2 0.189894
R1017 VP.n11 VP.n2 0.189894
R1018 VP.n14 VP.n13 0.189894
R1019 VP.n14 VP.n0 0.189894
R1020 VP.n20 VP.n0 0.189894
R1021 VP VP.n20 0.0516364
R1022 VTAIL.n11 VTAIL.t9 54.0319
R1023 VTAIL.n17 VTAIL.t1 54.0318
R1024 VTAIL.n2 VTAIL.t16 54.0318
R1025 VTAIL.n16 VTAIL.t18 54.0318
R1026 VTAIL.n15 VTAIL.n14 52.1355
R1027 VTAIL.n13 VTAIL.n12 52.1355
R1028 VTAIL.n10 VTAIL.n9 52.1355
R1029 VTAIL.n8 VTAIL.n7 52.1355
R1030 VTAIL.n19 VTAIL.n18 52.1353
R1031 VTAIL.n1 VTAIL.n0 52.1353
R1032 VTAIL.n4 VTAIL.n3 52.1353
R1033 VTAIL.n6 VTAIL.n5 52.1353
R1034 VTAIL.n8 VTAIL.n6 28.091
R1035 VTAIL.n17 VTAIL.n16 27.6169
R1036 VTAIL.n18 VTAIL.t3 1.89694
R1037 VTAIL.n18 VTAIL.t4 1.89694
R1038 VTAIL.n0 VTAIL.t2 1.89694
R1039 VTAIL.n0 VTAIL.t6 1.89694
R1040 VTAIL.n3 VTAIL.t17 1.89694
R1041 VTAIL.n3 VTAIL.t13 1.89694
R1042 VTAIL.n5 VTAIL.t12 1.89694
R1043 VTAIL.n5 VTAIL.t10 1.89694
R1044 VTAIL.n14 VTAIL.t15 1.89694
R1045 VTAIL.n14 VTAIL.t19 1.89694
R1046 VTAIL.n12 VTAIL.t11 1.89694
R1047 VTAIL.n12 VTAIL.t14 1.89694
R1048 VTAIL.n9 VTAIL.t5 1.89694
R1049 VTAIL.n9 VTAIL.t0 1.89694
R1050 VTAIL.n7 VTAIL.t7 1.89694
R1051 VTAIL.n7 VTAIL.t8 1.89694
R1052 VTAIL.n13 VTAIL.n11 0.707397
R1053 VTAIL.n2 VTAIL.n1 0.707397
R1054 VTAIL.n10 VTAIL.n8 0.474638
R1055 VTAIL.n11 VTAIL.n10 0.474638
R1056 VTAIL.n15 VTAIL.n13 0.474638
R1057 VTAIL.n16 VTAIL.n15 0.474638
R1058 VTAIL.n6 VTAIL.n4 0.474638
R1059 VTAIL.n4 VTAIL.n2 0.474638
R1060 VTAIL.n19 VTAIL.n17 0.474638
R1061 VTAIL VTAIL.n1 0.414293
R1062 VTAIL VTAIL.n19 0.0608448
R1063 VDD1.n1 VDD1.t9 71.1848
R1064 VDD1.n3 VDD1.t3 71.1847
R1065 VDD1.n5 VDD1.n4 69.1143
R1066 VDD1.n1 VDD1.n0 68.8143
R1067 VDD1.n7 VDD1.n6 68.8141
R1068 VDD1.n3 VDD1.n2 68.8141
R1069 VDD1.n7 VDD1.n5 41.5634
R1070 VDD1.n6 VDD1.t2 1.89694
R1071 VDD1.n6 VDD1.t8 1.89694
R1072 VDD1.n0 VDD1.t5 1.89694
R1073 VDD1.n0 VDD1.t6 1.89694
R1074 VDD1.n4 VDD1.t4 1.89694
R1075 VDD1.n4 VDD1.t1 1.89694
R1076 VDD1.n2 VDD1.t0 1.89694
R1077 VDD1.n2 VDD1.t7 1.89694
R1078 VDD1 VDD1.n7 0.297914
R1079 VDD1 VDD1.n1 0.177224
R1080 VDD1.n5 VDD1.n3 0.0636885
R1081 VN.n8 VN.t8 2071.14
R1082 VN.n2 VN.t9 2071.14
R1083 VN.n18 VN.t0 2071.14
R1084 VN.n12 VN.t3 2071.14
R1085 VN.n7 VN.t1 2020.02
R1086 VN.n5 VN.t4 2020.02
R1087 VN.n1 VN.t5 2020.02
R1088 VN.n17 VN.t6 2020.02
R1089 VN.n15 VN.t2 2020.02
R1090 VN.n11 VN.t7 2020.02
R1091 VN.n13 VN.n12 161.489
R1092 VN.n3 VN.n2 161.489
R1093 VN.n9 VN.n8 161.3
R1094 VN.n19 VN.n18 161.3
R1095 VN.n16 VN.n10 161.3
R1096 VN.n14 VN.n13 161.3
R1097 VN.n6 VN.n0 161.3
R1098 VN.n4 VN.n3 161.3
R1099 VN VN.n19 44.5516
R1100 VN.n4 VN.n1 43.8187
R1101 VN.n7 VN.n6 43.8187
R1102 VN.n17 VN.n16 43.8187
R1103 VN.n14 VN.n11 43.8187
R1104 VN.n5 VN.n4 36.5157
R1105 VN.n6 VN.n5 36.5157
R1106 VN.n16 VN.n15 36.5157
R1107 VN.n15 VN.n14 36.5157
R1108 VN.n2 VN.n1 29.2126
R1109 VN.n8 VN.n7 29.2126
R1110 VN.n18 VN.n17 29.2126
R1111 VN.n12 VN.n11 29.2126
R1112 VN.n19 VN.n10 0.189894
R1113 VN.n13 VN.n10 0.189894
R1114 VN.n3 VN.n0 0.189894
R1115 VN.n9 VN.n0 0.189894
R1116 VN VN.n9 0.0516364
R1117 VDD2.n1 VDD2.t0 71.1847
R1118 VDD2.n4 VDD2.t9 70.7107
R1119 VDD2.n3 VDD2.n2 69.1143
R1120 VDD2 VDD2.n7 69.1115
R1121 VDD2.n6 VDD2.n5 68.8143
R1122 VDD2.n1 VDD2.n0 68.8141
R1123 VDD2.n4 VDD2.n3 40.7433
R1124 VDD2.n7 VDD2.t2 1.89694
R1125 VDD2.n7 VDD2.t6 1.89694
R1126 VDD2.n5 VDD2.t3 1.89694
R1127 VDD2.n5 VDD2.t7 1.89694
R1128 VDD2.n2 VDD2.t8 1.89694
R1129 VDD2.n2 VDD2.t1 1.89694
R1130 VDD2.n0 VDD2.t4 1.89694
R1131 VDD2.n0 VDD2.t5 1.89694
R1132 VDD2.n6 VDD2.n4 0.474638
R1133 VDD2 VDD2.n6 0.177224
R1134 VDD2.n3 VDD2.n1 0.0636885
C0 VDD2 VN 4.4832f
C1 VDD2 VTAIL 33.2075f
C2 w_n1630_n4396# VDD2 2.22148f
C3 B VDD1 1.8462f
C4 VP VDD1 4.60935f
C5 B VP 1.06662f
C6 VDD1 VN 0.14795f
C7 B VN 0.735245f
C8 VP VN 5.83773f
C9 VTAIL VDD1 33.182697f
C10 B VTAIL 3.2006f
C11 VTAIL VP 3.82931f
C12 w_n1630_n4396# VDD1 2.20148f
C13 VTAIL VN 3.81422f
C14 B w_n1630_n4396# 8.041189f
C15 w_n1630_n4396# VP 3.06159f
C16 w_n1630_n4396# VN 2.85672f
C17 VDD2 VDD1 0.678095f
C18 B VDD2 1.87214f
C19 VDD2 VP 0.281616f
C20 w_n1630_n4396# VTAIL 3.89324f
C21 VDD2 VSUBS 1.705953f
C22 VDD1 VSUBS 1.149996f
C23 VTAIL VSUBS 0.587665f
C24 VN VSUBS 5.14046f
C25 VP VSUBS 1.415082f
C26 B VSUBS 2.843624f
C27 w_n1630_n4396# VSUBS 87.6875f
C28 VDD2.t0 VSUBS 5.06223f
C29 VDD2.t4 VSUBS 0.472126f
C30 VDD2.t5 VSUBS 0.472126f
C31 VDD2.n0 VSUBS 3.89511f
C32 VDD2.n1 VSUBS 1.63281f
C33 VDD2.t8 VSUBS 0.472126f
C34 VDD2.t1 VSUBS 0.472126f
C35 VDD2.n2 VSUBS 3.89854f
C36 VDD2.n3 VSUBS 3.12787f
C37 VDD2.t9 VSUBS 5.05641f
C38 VDD2.n4 VSUBS 4.06086f
C39 VDD2.t3 VSUBS 0.472126f
C40 VDD2.t7 VSUBS 0.472126f
C41 VDD2.n5 VSUBS 3.89511f
C42 VDD2.n6 VSUBS 0.759039f
C43 VDD2.t2 VSUBS 0.472126f
C44 VDD2.t6 VSUBS 0.472126f
C45 VDD2.n7 VSUBS 3.89848f
C46 VN.n0 VSUBS 0.068343f
C47 VN.t1 VSUBS 0.726432f
C48 VN.t4 VSUBS 0.726432f
C49 VN.t5 VSUBS 0.726432f
C50 VN.n1 VSUBS 0.280067f
C51 VN.t9 VSUBS 0.733417f
C52 VN.n2 VSUBS 0.30091f
C53 VN.n3 VSUBS 0.154282f
C54 VN.n4 VSUBS 0.024779f
C55 VN.n5 VSUBS 0.280067f
C56 VN.n6 VSUBS 0.024779f
C57 VN.n7 VSUBS 0.280067f
C58 VN.t8 VSUBS 0.733417f
C59 VN.n8 VSUBS 0.300809f
C60 VN.n9 VSUBS 0.052963f
C61 VN.n10 VSUBS 0.068343f
C62 VN.t0 VSUBS 0.733417f
C63 VN.t6 VSUBS 0.726432f
C64 VN.t2 VSUBS 0.726432f
C65 VN.t7 VSUBS 0.726432f
C66 VN.n11 VSUBS 0.280067f
C67 VN.t3 VSUBS 0.733417f
C68 VN.n12 VSUBS 0.30091f
C69 VN.n13 VSUBS 0.154282f
C70 VN.n14 VSUBS 0.024779f
C71 VN.n15 VSUBS 0.280067f
C72 VN.n16 VSUBS 0.024779f
C73 VN.n17 VSUBS 0.280067f
C74 VN.n18 VSUBS 0.300809f
C75 VN.n19 VSUBS 3.10857f
C76 VDD1.t9 VSUBS 5.05863f
C77 VDD1.t5 VSUBS 0.471787f
C78 VDD1.t6 VSUBS 0.471787f
C79 VDD1.n0 VSUBS 3.89232f
C80 VDD1.n1 VSUBS 1.63157f
C81 VDD1.t3 VSUBS 5.0586f
C82 VDD1.t0 VSUBS 0.471787f
C83 VDD1.t7 VSUBS 0.471787f
C84 VDD1.n2 VSUBS 3.89231f
C85 VDD1.n3 VSUBS 1.63164f
C86 VDD1.t4 VSUBS 0.471787f
C87 VDD1.t1 VSUBS 0.471787f
C88 VDD1.n4 VSUBS 3.89574f
C89 VDD1.n5 VSUBS 3.21852f
C90 VDD1.t2 VSUBS 0.471787f
C91 VDD1.t8 VSUBS 0.471787f
C92 VDD1.n6 VSUBS 3.8923f
C93 VDD1.n7 VSUBS 4.00086f
C94 VTAIL.t2 VSUBS 0.496427f
C95 VTAIL.t6 VSUBS 0.496427f
C96 VTAIL.n0 VSUBS 3.86709f
C97 VTAIL.n1 VSUBS 1.03229f
C98 VTAIL.t16 VSUBS 5.05513f
C99 VTAIL.n2 VSUBS 1.20526f
C100 VTAIL.t17 VSUBS 0.496427f
C101 VTAIL.t13 VSUBS 0.496427f
C102 VTAIL.n3 VSUBS 3.86709f
C103 VTAIL.n4 VSUBS 1.01193f
C104 VTAIL.t12 VSUBS 0.496427f
C105 VTAIL.t10 VSUBS 0.496427f
C106 VTAIL.n5 VSUBS 3.86709f
C107 VTAIL.n6 VSUBS 3.3108f
C108 VTAIL.t7 VSUBS 0.496427f
C109 VTAIL.t8 VSUBS 0.496427f
C110 VTAIL.n7 VSUBS 3.86709f
C111 VTAIL.n8 VSUBS 3.3108f
C112 VTAIL.t5 VSUBS 0.496427f
C113 VTAIL.t0 VSUBS 0.496427f
C114 VTAIL.n9 VSUBS 3.86709f
C115 VTAIL.n10 VSUBS 1.01192f
C116 VTAIL.t9 VSUBS 5.05517f
C117 VTAIL.n11 VSUBS 1.20522f
C118 VTAIL.t11 VSUBS 0.496427f
C119 VTAIL.t14 VSUBS 0.496427f
C120 VTAIL.n12 VSUBS 3.86709f
C121 VTAIL.n13 VSUBS 1.03941f
C122 VTAIL.t15 VSUBS 0.496427f
C123 VTAIL.t19 VSUBS 0.496427f
C124 VTAIL.n14 VSUBS 3.86709f
C125 VTAIL.n15 VSUBS 1.01192f
C126 VTAIL.t18 VSUBS 5.05513f
C127 VTAIL.n16 VSUBS 3.42065f
C128 VTAIL.t1 VSUBS 5.05513f
C129 VTAIL.n17 VSUBS 3.42065f
C130 VTAIL.t3 VSUBS 0.496427f
C131 VTAIL.t4 VSUBS 0.496427f
C132 VTAIL.n18 VSUBS 3.86709f
C133 VTAIL.n19 VSUBS 0.963059f
C134 VP.n0 VSUBS 0.069944f
C135 VP.t5 VSUBS 0.743453f
C136 VP.t2 VSUBS 0.743453f
C137 VP.t9 VSUBS 0.743453f
C138 VP.n1 VSUBS 0.286629f
C139 VP.n2 VSUBS 0.069944f
C140 VP.t7 VSUBS 0.743453f
C141 VP.t3 VSUBS 0.743453f
C142 VP.t4 VSUBS 0.743453f
C143 VP.n3 VSUBS 0.286629f
C144 VP.t0 VSUBS 0.750602f
C145 VP.n4 VSUBS 0.307961f
C146 VP.n5 VSUBS 0.157897f
C147 VP.n6 VSUBS 0.025359f
C148 VP.n7 VSUBS 0.286629f
C149 VP.n8 VSUBS 0.025359f
C150 VP.n9 VSUBS 0.286629f
C151 VP.t1 VSUBS 0.750602f
C152 VP.n10 VSUBS 0.307857f
C153 VP.n11 VSUBS 3.13563f
C154 VP.t6 VSUBS 0.750602f
C155 VP.n12 VSUBS 0.307857f
C156 VP.n13 VSUBS 3.19272f
C157 VP.n14 VSUBS 0.069944f
C158 VP.n15 VSUBS 0.025359f
C159 VP.n16 VSUBS 0.286629f
C160 VP.n17 VSUBS 0.025359f
C161 VP.n18 VSUBS 0.286629f
C162 VP.t8 VSUBS 0.750602f
C163 VP.n19 VSUBS 0.307857f
C164 VP.n20 VSUBS 0.054204f
C165 B.n0 VSUBS 0.004698f
C166 B.n1 VSUBS 0.004698f
C167 B.n2 VSUBS 0.00743f
C168 B.n3 VSUBS 0.00743f
C169 B.n4 VSUBS 0.00743f
C170 B.n5 VSUBS 0.00743f
C171 B.n6 VSUBS 0.00743f
C172 B.n7 VSUBS 0.00743f
C173 B.n8 VSUBS 0.00743f
C174 B.n9 VSUBS 0.00743f
C175 B.n10 VSUBS 0.00743f
C176 B.n11 VSUBS 0.017002f
C177 B.n12 VSUBS 0.00743f
C178 B.n13 VSUBS 0.00743f
C179 B.n14 VSUBS 0.00743f
C180 B.n15 VSUBS 0.00743f
C181 B.n16 VSUBS 0.00743f
C182 B.n17 VSUBS 0.00743f
C183 B.n18 VSUBS 0.00743f
C184 B.n19 VSUBS 0.00743f
C185 B.n20 VSUBS 0.00743f
C186 B.n21 VSUBS 0.00743f
C187 B.n22 VSUBS 0.00743f
C188 B.n23 VSUBS 0.00743f
C189 B.n24 VSUBS 0.00743f
C190 B.n25 VSUBS 0.00743f
C191 B.n26 VSUBS 0.00743f
C192 B.n27 VSUBS 0.00743f
C193 B.n28 VSUBS 0.00743f
C194 B.n29 VSUBS 0.00743f
C195 B.n30 VSUBS 0.00743f
C196 B.n31 VSUBS 0.00743f
C197 B.n32 VSUBS 0.00743f
C198 B.n33 VSUBS 0.00743f
C199 B.n34 VSUBS 0.00743f
C200 B.n35 VSUBS 0.00743f
C201 B.n36 VSUBS 0.00743f
C202 B.n37 VSUBS 0.00743f
C203 B.n38 VSUBS 0.00743f
C204 B.n39 VSUBS 0.00743f
C205 B.t11 VSUBS 0.612045f
C206 B.t10 VSUBS 0.616988f
C207 B.t9 VSUBS 0.154028f
C208 B.n40 VSUBS 0.108101f
C209 B.n41 VSUBS 0.066041f
C210 B.n42 VSUBS 0.00743f
C211 B.n43 VSUBS 0.00743f
C212 B.n44 VSUBS 0.00743f
C213 B.n45 VSUBS 0.00743f
C214 B.t2 VSUBS 0.612024f
C215 B.t1 VSUBS 0.616968f
C216 B.t0 VSUBS 0.154028f
C217 B.n46 VSUBS 0.108121f
C218 B.n47 VSUBS 0.066063f
C219 B.n48 VSUBS 0.017215f
C220 B.n49 VSUBS 0.00743f
C221 B.n50 VSUBS 0.00743f
C222 B.n51 VSUBS 0.00743f
C223 B.n52 VSUBS 0.00743f
C224 B.n53 VSUBS 0.00743f
C225 B.n54 VSUBS 0.00743f
C226 B.n55 VSUBS 0.00743f
C227 B.n56 VSUBS 0.00743f
C228 B.n57 VSUBS 0.00743f
C229 B.n58 VSUBS 0.00743f
C230 B.n59 VSUBS 0.00743f
C231 B.n60 VSUBS 0.00743f
C232 B.n61 VSUBS 0.00743f
C233 B.n62 VSUBS 0.00743f
C234 B.n63 VSUBS 0.00743f
C235 B.n64 VSUBS 0.00743f
C236 B.n65 VSUBS 0.00743f
C237 B.n66 VSUBS 0.00743f
C238 B.n67 VSUBS 0.00743f
C239 B.n68 VSUBS 0.00743f
C240 B.n69 VSUBS 0.00743f
C241 B.n70 VSUBS 0.00743f
C242 B.n71 VSUBS 0.00743f
C243 B.n72 VSUBS 0.00743f
C244 B.n73 VSUBS 0.00743f
C245 B.n74 VSUBS 0.00743f
C246 B.n75 VSUBS 0.00743f
C247 B.n76 VSUBS 0.00743f
C248 B.n77 VSUBS 0.016433f
C249 B.n78 VSUBS 0.00743f
C250 B.n79 VSUBS 0.00743f
C251 B.n80 VSUBS 0.00743f
C252 B.n81 VSUBS 0.00743f
C253 B.n82 VSUBS 0.00743f
C254 B.n83 VSUBS 0.00743f
C255 B.n84 VSUBS 0.00743f
C256 B.n85 VSUBS 0.00743f
C257 B.n86 VSUBS 0.00743f
C258 B.n87 VSUBS 0.00743f
C259 B.n88 VSUBS 0.00743f
C260 B.n89 VSUBS 0.00743f
C261 B.n90 VSUBS 0.00743f
C262 B.n91 VSUBS 0.00743f
C263 B.n92 VSUBS 0.00743f
C264 B.n93 VSUBS 0.00743f
C265 B.n94 VSUBS 0.00743f
C266 B.n95 VSUBS 0.016433f
C267 B.n96 VSUBS 0.00743f
C268 B.n97 VSUBS 0.00743f
C269 B.n98 VSUBS 0.00743f
C270 B.n99 VSUBS 0.00743f
C271 B.n100 VSUBS 0.00743f
C272 B.n101 VSUBS 0.00743f
C273 B.n102 VSUBS 0.00743f
C274 B.n103 VSUBS 0.00743f
C275 B.n104 VSUBS 0.00743f
C276 B.n105 VSUBS 0.00743f
C277 B.n106 VSUBS 0.00743f
C278 B.n107 VSUBS 0.00743f
C279 B.n108 VSUBS 0.00743f
C280 B.n109 VSUBS 0.00743f
C281 B.n110 VSUBS 0.00743f
C282 B.n111 VSUBS 0.00743f
C283 B.n112 VSUBS 0.00743f
C284 B.n113 VSUBS 0.00743f
C285 B.n114 VSUBS 0.00743f
C286 B.n115 VSUBS 0.00743f
C287 B.n116 VSUBS 0.00743f
C288 B.n117 VSUBS 0.00743f
C289 B.n118 VSUBS 0.00743f
C290 B.n119 VSUBS 0.00743f
C291 B.n120 VSUBS 0.00743f
C292 B.n121 VSUBS 0.00743f
C293 B.n122 VSUBS 0.00743f
C294 B.n123 VSUBS 0.00743f
C295 B.t7 VSUBS 0.612024f
C296 B.t8 VSUBS 0.616968f
C297 B.t6 VSUBS 0.154028f
C298 B.n124 VSUBS 0.108121f
C299 B.n125 VSUBS 0.066063f
C300 B.n126 VSUBS 0.017215f
C301 B.n127 VSUBS 0.00743f
C302 B.n128 VSUBS 0.00743f
C303 B.n129 VSUBS 0.00743f
C304 B.n130 VSUBS 0.00743f
C305 B.n131 VSUBS 0.00743f
C306 B.t4 VSUBS 0.612045f
C307 B.t5 VSUBS 0.616988f
C308 B.t3 VSUBS 0.154028f
C309 B.n132 VSUBS 0.108101f
C310 B.n133 VSUBS 0.066041f
C311 B.n134 VSUBS 0.00743f
C312 B.n135 VSUBS 0.00743f
C313 B.n136 VSUBS 0.00743f
C314 B.n137 VSUBS 0.00743f
C315 B.n138 VSUBS 0.00743f
C316 B.n139 VSUBS 0.00743f
C317 B.n140 VSUBS 0.00743f
C318 B.n141 VSUBS 0.00743f
C319 B.n142 VSUBS 0.00743f
C320 B.n143 VSUBS 0.00743f
C321 B.n144 VSUBS 0.00743f
C322 B.n145 VSUBS 0.00743f
C323 B.n146 VSUBS 0.00743f
C324 B.n147 VSUBS 0.00743f
C325 B.n148 VSUBS 0.00743f
C326 B.n149 VSUBS 0.00743f
C327 B.n150 VSUBS 0.00743f
C328 B.n151 VSUBS 0.00743f
C329 B.n152 VSUBS 0.00743f
C330 B.n153 VSUBS 0.00743f
C331 B.n154 VSUBS 0.00743f
C332 B.n155 VSUBS 0.00743f
C333 B.n156 VSUBS 0.00743f
C334 B.n157 VSUBS 0.00743f
C335 B.n158 VSUBS 0.00743f
C336 B.n159 VSUBS 0.00743f
C337 B.n160 VSUBS 0.00743f
C338 B.n161 VSUBS 0.017002f
C339 B.n162 VSUBS 0.00743f
C340 B.n163 VSUBS 0.00743f
C341 B.n164 VSUBS 0.00743f
C342 B.n165 VSUBS 0.00743f
C343 B.n166 VSUBS 0.00743f
C344 B.n167 VSUBS 0.00743f
C345 B.n168 VSUBS 0.00743f
C346 B.n169 VSUBS 0.00743f
C347 B.n170 VSUBS 0.00743f
C348 B.n171 VSUBS 0.00743f
C349 B.n172 VSUBS 0.00743f
C350 B.n173 VSUBS 0.00743f
C351 B.n174 VSUBS 0.00743f
C352 B.n175 VSUBS 0.00743f
C353 B.n176 VSUBS 0.00743f
C354 B.n177 VSUBS 0.00743f
C355 B.n178 VSUBS 0.00743f
C356 B.n179 VSUBS 0.00743f
C357 B.n180 VSUBS 0.00743f
C358 B.n181 VSUBS 0.00743f
C359 B.n182 VSUBS 0.00743f
C360 B.n183 VSUBS 0.00743f
C361 B.n184 VSUBS 0.00743f
C362 B.n185 VSUBS 0.00743f
C363 B.n186 VSUBS 0.00743f
C364 B.n187 VSUBS 0.00743f
C365 B.n188 VSUBS 0.00743f
C366 B.n189 VSUBS 0.00743f
C367 B.n190 VSUBS 0.00743f
C368 B.n191 VSUBS 0.00743f
C369 B.n192 VSUBS 0.00743f
C370 B.n193 VSUBS 0.00743f
C371 B.n194 VSUBS 0.016433f
C372 B.n195 VSUBS 0.016433f
C373 B.n196 VSUBS 0.017002f
C374 B.n197 VSUBS 0.00743f
C375 B.n198 VSUBS 0.00743f
C376 B.n199 VSUBS 0.00743f
C377 B.n200 VSUBS 0.00743f
C378 B.n201 VSUBS 0.00743f
C379 B.n202 VSUBS 0.00743f
C380 B.n203 VSUBS 0.00743f
C381 B.n204 VSUBS 0.00743f
C382 B.n205 VSUBS 0.00743f
C383 B.n206 VSUBS 0.00743f
C384 B.n207 VSUBS 0.00743f
C385 B.n208 VSUBS 0.00743f
C386 B.n209 VSUBS 0.00743f
C387 B.n210 VSUBS 0.00743f
C388 B.n211 VSUBS 0.00743f
C389 B.n212 VSUBS 0.00743f
C390 B.n213 VSUBS 0.00743f
C391 B.n214 VSUBS 0.00743f
C392 B.n215 VSUBS 0.00743f
C393 B.n216 VSUBS 0.00743f
C394 B.n217 VSUBS 0.00743f
C395 B.n218 VSUBS 0.00743f
C396 B.n219 VSUBS 0.00743f
C397 B.n220 VSUBS 0.00743f
C398 B.n221 VSUBS 0.00743f
C399 B.n222 VSUBS 0.00743f
C400 B.n223 VSUBS 0.00743f
C401 B.n224 VSUBS 0.00743f
C402 B.n225 VSUBS 0.00743f
C403 B.n226 VSUBS 0.00743f
C404 B.n227 VSUBS 0.00743f
C405 B.n228 VSUBS 0.00743f
C406 B.n229 VSUBS 0.00743f
C407 B.n230 VSUBS 0.00743f
C408 B.n231 VSUBS 0.00743f
C409 B.n232 VSUBS 0.00743f
C410 B.n233 VSUBS 0.00743f
C411 B.n234 VSUBS 0.00743f
C412 B.n235 VSUBS 0.00743f
C413 B.n236 VSUBS 0.00743f
C414 B.n237 VSUBS 0.00743f
C415 B.n238 VSUBS 0.00743f
C416 B.n239 VSUBS 0.00743f
C417 B.n240 VSUBS 0.00743f
C418 B.n241 VSUBS 0.00743f
C419 B.n242 VSUBS 0.00743f
C420 B.n243 VSUBS 0.00743f
C421 B.n244 VSUBS 0.00743f
C422 B.n245 VSUBS 0.00743f
C423 B.n246 VSUBS 0.00743f
C424 B.n247 VSUBS 0.00743f
C425 B.n248 VSUBS 0.00743f
C426 B.n249 VSUBS 0.00743f
C427 B.n250 VSUBS 0.00743f
C428 B.n251 VSUBS 0.00743f
C429 B.n252 VSUBS 0.00743f
C430 B.n253 VSUBS 0.00743f
C431 B.n254 VSUBS 0.00743f
C432 B.n255 VSUBS 0.00743f
C433 B.n256 VSUBS 0.00743f
C434 B.n257 VSUBS 0.00743f
C435 B.n258 VSUBS 0.00743f
C436 B.n259 VSUBS 0.00743f
C437 B.n260 VSUBS 0.00743f
C438 B.n261 VSUBS 0.00743f
C439 B.n262 VSUBS 0.00743f
C440 B.n263 VSUBS 0.00743f
C441 B.n264 VSUBS 0.00743f
C442 B.n265 VSUBS 0.00743f
C443 B.n266 VSUBS 0.00743f
C444 B.n267 VSUBS 0.00743f
C445 B.n268 VSUBS 0.00743f
C446 B.n269 VSUBS 0.00743f
C447 B.n270 VSUBS 0.00743f
C448 B.n271 VSUBS 0.00743f
C449 B.n272 VSUBS 0.00743f
C450 B.n273 VSUBS 0.00743f
C451 B.n274 VSUBS 0.00743f
C452 B.n275 VSUBS 0.00743f
C453 B.n276 VSUBS 0.00743f
C454 B.n277 VSUBS 0.00743f
C455 B.n278 VSUBS 0.00743f
C456 B.n279 VSUBS 0.00743f
C457 B.n280 VSUBS 0.005136f
C458 B.n281 VSUBS 0.017215f
C459 B.n282 VSUBS 0.00601f
C460 B.n283 VSUBS 0.00743f
C461 B.n284 VSUBS 0.00743f
C462 B.n285 VSUBS 0.00743f
C463 B.n286 VSUBS 0.00743f
C464 B.n287 VSUBS 0.00743f
C465 B.n288 VSUBS 0.00743f
C466 B.n289 VSUBS 0.00743f
C467 B.n290 VSUBS 0.00743f
C468 B.n291 VSUBS 0.00743f
C469 B.n292 VSUBS 0.00743f
C470 B.n293 VSUBS 0.00743f
C471 B.n294 VSUBS 0.00601f
C472 B.n295 VSUBS 0.00743f
C473 B.n296 VSUBS 0.00743f
C474 B.n297 VSUBS 0.005136f
C475 B.n298 VSUBS 0.00743f
C476 B.n299 VSUBS 0.00743f
C477 B.n300 VSUBS 0.00743f
C478 B.n301 VSUBS 0.00743f
C479 B.n302 VSUBS 0.00743f
C480 B.n303 VSUBS 0.00743f
C481 B.n304 VSUBS 0.00743f
C482 B.n305 VSUBS 0.00743f
C483 B.n306 VSUBS 0.00743f
C484 B.n307 VSUBS 0.00743f
C485 B.n308 VSUBS 0.00743f
C486 B.n309 VSUBS 0.00743f
C487 B.n310 VSUBS 0.00743f
C488 B.n311 VSUBS 0.00743f
C489 B.n312 VSUBS 0.00743f
C490 B.n313 VSUBS 0.00743f
C491 B.n314 VSUBS 0.00743f
C492 B.n315 VSUBS 0.00743f
C493 B.n316 VSUBS 0.00743f
C494 B.n317 VSUBS 0.00743f
C495 B.n318 VSUBS 0.00743f
C496 B.n319 VSUBS 0.00743f
C497 B.n320 VSUBS 0.00743f
C498 B.n321 VSUBS 0.00743f
C499 B.n322 VSUBS 0.00743f
C500 B.n323 VSUBS 0.00743f
C501 B.n324 VSUBS 0.00743f
C502 B.n325 VSUBS 0.00743f
C503 B.n326 VSUBS 0.00743f
C504 B.n327 VSUBS 0.00743f
C505 B.n328 VSUBS 0.00743f
C506 B.n329 VSUBS 0.00743f
C507 B.n330 VSUBS 0.00743f
C508 B.n331 VSUBS 0.00743f
C509 B.n332 VSUBS 0.00743f
C510 B.n333 VSUBS 0.00743f
C511 B.n334 VSUBS 0.00743f
C512 B.n335 VSUBS 0.00743f
C513 B.n336 VSUBS 0.00743f
C514 B.n337 VSUBS 0.00743f
C515 B.n338 VSUBS 0.00743f
C516 B.n339 VSUBS 0.00743f
C517 B.n340 VSUBS 0.00743f
C518 B.n341 VSUBS 0.00743f
C519 B.n342 VSUBS 0.00743f
C520 B.n343 VSUBS 0.00743f
C521 B.n344 VSUBS 0.00743f
C522 B.n345 VSUBS 0.00743f
C523 B.n346 VSUBS 0.00743f
C524 B.n347 VSUBS 0.00743f
C525 B.n348 VSUBS 0.00743f
C526 B.n349 VSUBS 0.00743f
C527 B.n350 VSUBS 0.00743f
C528 B.n351 VSUBS 0.00743f
C529 B.n352 VSUBS 0.00743f
C530 B.n353 VSUBS 0.00743f
C531 B.n354 VSUBS 0.00743f
C532 B.n355 VSUBS 0.00743f
C533 B.n356 VSUBS 0.00743f
C534 B.n357 VSUBS 0.00743f
C535 B.n358 VSUBS 0.00743f
C536 B.n359 VSUBS 0.00743f
C537 B.n360 VSUBS 0.00743f
C538 B.n361 VSUBS 0.00743f
C539 B.n362 VSUBS 0.00743f
C540 B.n363 VSUBS 0.00743f
C541 B.n364 VSUBS 0.00743f
C542 B.n365 VSUBS 0.00743f
C543 B.n366 VSUBS 0.00743f
C544 B.n367 VSUBS 0.00743f
C545 B.n368 VSUBS 0.00743f
C546 B.n369 VSUBS 0.00743f
C547 B.n370 VSUBS 0.00743f
C548 B.n371 VSUBS 0.00743f
C549 B.n372 VSUBS 0.00743f
C550 B.n373 VSUBS 0.00743f
C551 B.n374 VSUBS 0.00743f
C552 B.n375 VSUBS 0.00743f
C553 B.n376 VSUBS 0.00743f
C554 B.n377 VSUBS 0.00743f
C555 B.n378 VSUBS 0.00743f
C556 B.n379 VSUBS 0.00743f
C557 B.n380 VSUBS 0.017002f
C558 B.n381 VSUBS 0.017002f
C559 B.n382 VSUBS 0.016433f
C560 B.n383 VSUBS 0.00743f
C561 B.n384 VSUBS 0.00743f
C562 B.n385 VSUBS 0.00743f
C563 B.n386 VSUBS 0.00743f
C564 B.n387 VSUBS 0.00743f
C565 B.n388 VSUBS 0.00743f
C566 B.n389 VSUBS 0.00743f
C567 B.n390 VSUBS 0.00743f
C568 B.n391 VSUBS 0.00743f
C569 B.n392 VSUBS 0.00743f
C570 B.n393 VSUBS 0.00743f
C571 B.n394 VSUBS 0.00743f
C572 B.n395 VSUBS 0.00743f
C573 B.n396 VSUBS 0.00743f
C574 B.n397 VSUBS 0.00743f
C575 B.n398 VSUBS 0.00743f
C576 B.n399 VSUBS 0.00743f
C577 B.n400 VSUBS 0.00743f
C578 B.n401 VSUBS 0.00743f
C579 B.n402 VSUBS 0.00743f
C580 B.n403 VSUBS 0.00743f
C581 B.n404 VSUBS 0.00743f
C582 B.n405 VSUBS 0.00743f
C583 B.n406 VSUBS 0.00743f
C584 B.n407 VSUBS 0.00743f
C585 B.n408 VSUBS 0.00743f
C586 B.n409 VSUBS 0.00743f
C587 B.n410 VSUBS 0.00743f
C588 B.n411 VSUBS 0.00743f
C589 B.n412 VSUBS 0.00743f
C590 B.n413 VSUBS 0.00743f
C591 B.n414 VSUBS 0.00743f
C592 B.n415 VSUBS 0.00743f
C593 B.n416 VSUBS 0.00743f
C594 B.n417 VSUBS 0.00743f
C595 B.n418 VSUBS 0.00743f
C596 B.n419 VSUBS 0.00743f
C597 B.n420 VSUBS 0.00743f
C598 B.n421 VSUBS 0.00743f
C599 B.n422 VSUBS 0.00743f
C600 B.n423 VSUBS 0.00743f
C601 B.n424 VSUBS 0.00743f
C602 B.n425 VSUBS 0.00743f
C603 B.n426 VSUBS 0.00743f
C604 B.n427 VSUBS 0.00743f
C605 B.n428 VSUBS 0.00743f
C606 B.n429 VSUBS 0.00743f
C607 B.n430 VSUBS 0.00743f
C608 B.n431 VSUBS 0.00743f
C609 B.n432 VSUBS 0.00743f
C610 B.n433 VSUBS 0.00743f
C611 B.n434 VSUBS 0.00743f
C612 B.n435 VSUBS 0.00743f
C613 B.n436 VSUBS 0.017366f
C614 B.n437 VSUBS 0.01607f
C615 B.n438 VSUBS 0.017002f
C616 B.n439 VSUBS 0.00743f
C617 B.n440 VSUBS 0.00743f
C618 B.n441 VSUBS 0.00743f
C619 B.n442 VSUBS 0.00743f
C620 B.n443 VSUBS 0.00743f
C621 B.n444 VSUBS 0.00743f
C622 B.n445 VSUBS 0.00743f
C623 B.n446 VSUBS 0.00743f
C624 B.n447 VSUBS 0.00743f
C625 B.n448 VSUBS 0.00743f
C626 B.n449 VSUBS 0.00743f
C627 B.n450 VSUBS 0.00743f
C628 B.n451 VSUBS 0.00743f
C629 B.n452 VSUBS 0.00743f
C630 B.n453 VSUBS 0.00743f
C631 B.n454 VSUBS 0.00743f
C632 B.n455 VSUBS 0.00743f
C633 B.n456 VSUBS 0.00743f
C634 B.n457 VSUBS 0.00743f
C635 B.n458 VSUBS 0.00743f
C636 B.n459 VSUBS 0.00743f
C637 B.n460 VSUBS 0.00743f
C638 B.n461 VSUBS 0.00743f
C639 B.n462 VSUBS 0.00743f
C640 B.n463 VSUBS 0.00743f
C641 B.n464 VSUBS 0.00743f
C642 B.n465 VSUBS 0.00743f
C643 B.n466 VSUBS 0.00743f
C644 B.n467 VSUBS 0.00743f
C645 B.n468 VSUBS 0.00743f
C646 B.n469 VSUBS 0.00743f
C647 B.n470 VSUBS 0.00743f
C648 B.n471 VSUBS 0.00743f
C649 B.n472 VSUBS 0.00743f
C650 B.n473 VSUBS 0.00743f
C651 B.n474 VSUBS 0.00743f
C652 B.n475 VSUBS 0.00743f
C653 B.n476 VSUBS 0.00743f
C654 B.n477 VSUBS 0.00743f
C655 B.n478 VSUBS 0.00743f
C656 B.n479 VSUBS 0.00743f
C657 B.n480 VSUBS 0.00743f
C658 B.n481 VSUBS 0.00743f
C659 B.n482 VSUBS 0.00743f
C660 B.n483 VSUBS 0.00743f
C661 B.n484 VSUBS 0.00743f
C662 B.n485 VSUBS 0.00743f
C663 B.n486 VSUBS 0.00743f
C664 B.n487 VSUBS 0.00743f
C665 B.n488 VSUBS 0.00743f
C666 B.n489 VSUBS 0.00743f
C667 B.n490 VSUBS 0.00743f
C668 B.n491 VSUBS 0.00743f
C669 B.n492 VSUBS 0.00743f
C670 B.n493 VSUBS 0.00743f
C671 B.n494 VSUBS 0.00743f
C672 B.n495 VSUBS 0.00743f
C673 B.n496 VSUBS 0.00743f
C674 B.n497 VSUBS 0.00743f
C675 B.n498 VSUBS 0.00743f
C676 B.n499 VSUBS 0.00743f
C677 B.n500 VSUBS 0.00743f
C678 B.n501 VSUBS 0.00743f
C679 B.n502 VSUBS 0.00743f
C680 B.n503 VSUBS 0.00743f
C681 B.n504 VSUBS 0.00743f
C682 B.n505 VSUBS 0.00743f
C683 B.n506 VSUBS 0.00743f
C684 B.n507 VSUBS 0.00743f
C685 B.n508 VSUBS 0.00743f
C686 B.n509 VSUBS 0.00743f
C687 B.n510 VSUBS 0.00743f
C688 B.n511 VSUBS 0.00743f
C689 B.n512 VSUBS 0.00743f
C690 B.n513 VSUBS 0.00743f
C691 B.n514 VSUBS 0.00743f
C692 B.n515 VSUBS 0.00743f
C693 B.n516 VSUBS 0.00743f
C694 B.n517 VSUBS 0.00743f
C695 B.n518 VSUBS 0.00743f
C696 B.n519 VSUBS 0.00743f
C697 B.n520 VSUBS 0.00743f
C698 B.n521 VSUBS 0.005136f
C699 B.n522 VSUBS 0.00743f
C700 B.n523 VSUBS 0.00743f
C701 B.n524 VSUBS 0.00601f
C702 B.n525 VSUBS 0.00743f
C703 B.n526 VSUBS 0.00743f
C704 B.n527 VSUBS 0.00743f
C705 B.n528 VSUBS 0.00743f
C706 B.n529 VSUBS 0.00743f
C707 B.n530 VSUBS 0.00743f
C708 B.n531 VSUBS 0.00743f
C709 B.n532 VSUBS 0.00743f
C710 B.n533 VSUBS 0.00743f
C711 B.n534 VSUBS 0.00743f
C712 B.n535 VSUBS 0.00743f
C713 B.n536 VSUBS 0.00601f
C714 B.n537 VSUBS 0.017215f
C715 B.n538 VSUBS 0.005136f
C716 B.n539 VSUBS 0.00743f
C717 B.n540 VSUBS 0.00743f
C718 B.n541 VSUBS 0.00743f
C719 B.n542 VSUBS 0.00743f
C720 B.n543 VSUBS 0.00743f
C721 B.n544 VSUBS 0.00743f
C722 B.n545 VSUBS 0.00743f
C723 B.n546 VSUBS 0.00743f
C724 B.n547 VSUBS 0.00743f
C725 B.n548 VSUBS 0.00743f
C726 B.n549 VSUBS 0.00743f
C727 B.n550 VSUBS 0.00743f
C728 B.n551 VSUBS 0.00743f
C729 B.n552 VSUBS 0.00743f
C730 B.n553 VSUBS 0.00743f
C731 B.n554 VSUBS 0.00743f
C732 B.n555 VSUBS 0.00743f
C733 B.n556 VSUBS 0.00743f
C734 B.n557 VSUBS 0.00743f
C735 B.n558 VSUBS 0.00743f
C736 B.n559 VSUBS 0.00743f
C737 B.n560 VSUBS 0.00743f
C738 B.n561 VSUBS 0.00743f
C739 B.n562 VSUBS 0.00743f
C740 B.n563 VSUBS 0.00743f
C741 B.n564 VSUBS 0.00743f
C742 B.n565 VSUBS 0.00743f
C743 B.n566 VSUBS 0.00743f
C744 B.n567 VSUBS 0.00743f
C745 B.n568 VSUBS 0.00743f
C746 B.n569 VSUBS 0.00743f
C747 B.n570 VSUBS 0.00743f
C748 B.n571 VSUBS 0.00743f
C749 B.n572 VSUBS 0.00743f
C750 B.n573 VSUBS 0.00743f
C751 B.n574 VSUBS 0.00743f
C752 B.n575 VSUBS 0.00743f
C753 B.n576 VSUBS 0.00743f
C754 B.n577 VSUBS 0.00743f
C755 B.n578 VSUBS 0.00743f
C756 B.n579 VSUBS 0.00743f
C757 B.n580 VSUBS 0.00743f
C758 B.n581 VSUBS 0.00743f
C759 B.n582 VSUBS 0.00743f
C760 B.n583 VSUBS 0.00743f
C761 B.n584 VSUBS 0.00743f
C762 B.n585 VSUBS 0.00743f
C763 B.n586 VSUBS 0.00743f
C764 B.n587 VSUBS 0.00743f
C765 B.n588 VSUBS 0.00743f
C766 B.n589 VSUBS 0.00743f
C767 B.n590 VSUBS 0.00743f
C768 B.n591 VSUBS 0.00743f
C769 B.n592 VSUBS 0.00743f
C770 B.n593 VSUBS 0.00743f
C771 B.n594 VSUBS 0.00743f
C772 B.n595 VSUBS 0.00743f
C773 B.n596 VSUBS 0.00743f
C774 B.n597 VSUBS 0.00743f
C775 B.n598 VSUBS 0.00743f
C776 B.n599 VSUBS 0.00743f
C777 B.n600 VSUBS 0.00743f
C778 B.n601 VSUBS 0.00743f
C779 B.n602 VSUBS 0.00743f
C780 B.n603 VSUBS 0.00743f
C781 B.n604 VSUBS 0.00743f
C782 B.n605 VSUBS 0.00743f
C783 B.n606 VSUBS 0.00743f
C784 B.n607 VSUBS 0.00743f
C785 B.n608 VSUBS 0.00743f
C786 B.n609 VSUBS 0.00743f
C787 B.n610 VSUBS 0.00743f
C788 B.n611 VSUBS 0.00743f
C789 B.n612 VSUBS 0.00743f
C790 B.n613 VSUBS 0.00743f
C791 B.n614 VSUBS 0.00743f
C792 B.n615 VSUBS 0.00743f
C793 B.n616 VSUBS 0.00743f
C794 B.n617 VSUBS 0.00743f
C795 B.n618 VSUBS 0.00743f
C796 B.n619 VSUBS 0.00743f
C797 B.n620 VSUBS 0.00743f
C798 B.n621 VSUBS 0.00743f
C799 B.n622 VSUBS 0.017002f
C800 B.n623 VSUBS 0.016433f
C801 B.n624 VSUBS 0.016433f
C802 B.n625 VSUBS 0.00743f
C803 B.n626 VSUBS 0.00743f
C804 B.n627 VSUBS 0.00743f
C805 B.n628 VSUBS 0.00743f
C806 B.n629 VSUBS 0.00743f
C807 B.n630 VSUBS 0.00743f
C808 B.n631 VSUBS 0.00743f
C809 B.n632 VSUBS 0.00743f
C810 B.n633 VSUBS 0.00743f
C811 B.n634 VSUBS 0.00743f
C812 B.n635 VSUBS 0.00743f
C813 B.n636 VSUBS 0.00743f
C814 B.n637 VSUBS 0.00743f
C815 B.n638 VSUBS 0.00743f
C816 B.n639 VSUBS 0.00743f
C817 B.n640 VSUBS 0.00743f
C818 B.n641 VSUBS 0.00743f
C819 B.n642 VSUBS 0.00743f
C820 B.n643 VSUBS 0.00743f
C821 B.n644 VSUBS 0.00743f
C822 B.n645 VSUBS 0.00743f
C823 B.n646 VSUBS 0.00743f
C824 B.n647 VSUBS 0.00743f
C825 B.n648 VSUBS 0.00743f
C826 B.n649 VSUBS 0.00743f
C827 B.n650 VSUBS 0.00743f
C828 B.n651 VSUBS 0.016824f
.ends

