* NGSPICE file created from diff_pair_sample_0007.ext - technology: sky130A

.subckt diff_pair_sample_0007 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=0 ps=0 w=18.33 l=0.95
X1 VDD1.t5 VP.t0 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=3.02445 ps=18.66 w=18.33 l=0.95
X2 VDD2.t5 VN.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=3.02445 ps=18.66 w=18.33 l=0.95
X3 VDD1.t4 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=3.02445 ps=18.66 w=18.33 l=0.95
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=0 ps=0 w=18.33 l=0.95
X5 VTAIL.t5 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=3.02445 ps=18.66 w=18.33 l=0.95
X6 VTAIL.t10 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=3.02445 ps=18.66 w=18.33 l=0.95
X7 VDD1.t1 VP.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=7.1487 ps=37.44 w=18.33 l=0.95
X8 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=7.1487 ps=37.44 w=18.33 l=0.95
X9 VDD2.t3 VN.t2 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=7.1487 ps=37.44 w=18.33 l=0.95
X10 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=0 ps=0 w=18.33 l=0.95
X11 VTAIL.t4 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=3.02445 ps=18.66 w=18.33 l=0.95
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=0 ps=0 w=18.33 l=0.95
X13 VDD1.t0 VP.t5 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=7.1487 ps=37.44 w=18.33 l=0.95
X14 VTAIL.t3 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=3.02445 pd=18.66 as=3.02445 ps=18.66 w=18.33 l=0.95
X15 VDD2.t0 VN.t5 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1487 pd=37.44 as=3.02445 ps=18.66 w=18.33 l=0.95
R0 B.n484 B.t17 667.578
R1 B.n482 B.t13 667.578
R2 B.n115 B.t6 667.578
R3 B.n112 B.t10 667.578
R4 B.n844 B.n843 585
R5 B.n370 B.n110 585
R6 B.n369 B.n368 585
R7 B.n367 B.n366 585
R8 B.n365 B.n364 585
R9 B.n363 B.n362 585
R10 B.n361 B.n360 585
R11 B.n359 B.n358 585
R12 B.n357 B.n356 585
R13 B.n355 B.n354 585
R14 B.n353 B.n352 585
R15 B.n351 B.n350 585
R16 B.n349 B.n348 585
R17 B.n347 B.n346 585
R18 B.n345 B.n344 585
R19 B.n343 B.n342 585
R20 B.n341 B.n340 585
R21 B.n339 B.n338 585
R22 B.n337 B.n336 585
R23 B.n335 B.n334 585
R24 B.n333 B.n332 585
R25 B.n331 B.n330 585
R26 B.n329 B.n328 585
R27 B.n327 B.n326 585
R28 B.n325 B.n324 585
R29 B.n323 B.n322 585
R30 B.n321 B.n320 585
R31 B.n319 B.n318 585
R32 B.n317 B.n316 585
R33 B.n315 B.n314 585
R34 B.n313 B.n312 585
R35 B.n311 B.n310 585
R36 B.n309 B.n308 585
R37 B.n307 B.n306 585
R38 B.n305 B.n304 585
R39 B.n303 B.n302 585
R40 B.n301 B.n300 585
R41 B.n299 B.n298 585
R42 B.n297 B.n296 585
R43 B.n295 B.n294 585
R44 B.n293 B.n292 585
R45 B.n291 B.n290 585
R46 B.n289 B.n288 585
R47 B.n287 B.n286 585
R48 B.n285 B.n284 585
R49 B.n283 B.n282 585
R50 B.n281 B.n280 585
R51 B.n279 B.n278 585
R52 B.n277 B.n276 585
R53 B.n275 B.n274 585
R54 B.n273 B.n272 585
R55 B.n271 B.n270 585
R56 B.n269 B.n268 585
R57 B.n267 B.n266 585
R58 B.n265 B.n264 585
R59 B.n263 B.n262 585
R60 B.n261 B.n260 585
R61 B.n259 B.n258 585
R62 B.n257 B.n256 585
R63 B.n255 B.n254 585
R64 B.n253 B.n252 585
R65 B.n251 B.n250 585
R66 B.n249 B.n248 585
R67 B.n247 B.n246 585
R68 B.n245 B.n244 585
R69 B.n243 B.n242 585
R70 B.n241 B.n240 585
R71 B.n239 B.n238 585
R72 B.n237 B.n236 585
R73 B.n235 B.n234 585
R74 B.n233 B.n232 585
R75 B.n231 B.n230 585
R76 B.n229 B.n228 585
R77 B.n227 B.n226 585
R78 B.n225 B.n224 585
R79 B.n223 B.n222 585
R80 B.n221 B.n220 585
R81 B.n219 B.n218 585
R82 B.n217 B.n216 585
R83 B.n215 B.n214 585
R84 B.n213 B.n212 585
R85 B.n211 B.n210 585
R86 B.n209 B.n208 585
R87 B.n207 B.n206 585
R88 B.n205 B.n204 585
R89 B.n203 B.n202 585
R90 B.n201 B.n200 585
R91 B.n199 B.n198 585
R92 B.n197 B.n196 585
R93 B.n195 B.n194 585
R94 B.n193 B.n192 585
R95 B.n191 B.n190 585
R96 B.n189 B.n188 585
R97 B.n187 B.n186 585
R98 B.n185 B.n184 585
R99 B.n183 B.n182 585
R100 B.n181 B.n180 585
R101 B.n179 B.n178 585
R102 B.n177 B.n176 585
R103 B.n175 B.n174 585
R104 B.n173 B.n172 585
R105 B.n171 B.n170 585
R106 B.n169 B.n168 585
R107 B.n167 B.n166 585
R108 B.n165 B.n164 585
R109 B.n163 B.n162 585
R110 B.n161 B.n160 585
R111 B.n159 B.n158 585
R112 B.n157 B.n156 585
R113 B.n155 B.n154 585
R114 B.n153 B.n152 585
R115 B.n151 B.n150 585
R116 B.n149 B.n148 585
R117 B.n147 B.n146 585
R118 B.n145 B.n144 585
R119 B.n143 B.n142 585
R120 B.n141 B.n140 585
R121 B.n139 B.n138 585
R122 B.n137 B.n136 585
R123 B.n135 B.n134 585
R124 B.n133 B.n132 585
R125 B.n131 B.n130 585
R126 B.n129 B.n128 585
R127 B.n127 B.n126 585
R128 B.n125 B.n124 585
R129 B.n123 B.n122 585
R130 B.n121 B.n120 585
R131 B.n119 B.n118 585
R132 B.n46 B.n45 585
R133 B.n849 B.n848 585
R134 B.n842 B.n111 585
R135 B.n111 B.n43 585
R136 B.n841 B.n42 585
R137 B.n853 B.n42 585
R138 B.n840 B.n41 585
R139 B.n854 B.n41 585
R140 B.n839 B.n40 585
R141 B.n855 B.n40 585
R142 B.n838 B.n837 585
R143 B.n837 B.n36 585
R144 B.n836 B.n35 585
R145 B.n861 B.n35 585
R146 B.n835 B.n34 585
R147 B.n862 B.n34 585
R148 B.n834 B.n33 585
R149 B.n863 B.n33 585
R150 B.n833 B.n832 585
R151 B.n832 B.n29 585
R152 B.n831 B.n28 585
R153 B.n869 B.n28 585
R154 B.n830 B.n27 585
R155 B.n870 B.n27 585
R156 B.n829 B.n26 585
R157 B.n871 B.n26 585
R158 B.n828 B.n827 585
R159 B.n827 B.n22 585
R160 B.n826 B.n21 585
R161 B.n877 B.n21 585
R162 B.n825 B.n20 585
R163 B.n878 B.n20 585
R164 B.n824 B.n19 585
R165 B.n879 B.n19 585
R166 B.n823 B.n822 585
R167 B.n822 B.n15 585
R168 B.n821 B.n14 585
R169 B.n885 B.n14 585
R170 B.n820 B.n13 585
R171 B.n886 B.n13 585
R172 B.n819 B.n12 585
R173 B.n887 B.n12 585
R174 B.n818 B.n817 585
R175 B.n817 B.n8 585
R176 B.n816 B.n7 585
R177 B.n893 B.n7 585
R178 B.n815 B.n6 585
R179 B.n894 B.n6 585
R180 B.n814 B.n5 585
R181 B.n895 B.n5 585
R182 B.n813 B.n812 585
R183 B.n812 B.n4 585
R184 B.n811 B.n371 585
R185 B.n811 B.n810 585
R186 B.n801 B.n372 585
R187 B.n373 B.n372 585
R188 B.n803 B.n802 585
R189 B.n804 B.n803 585
R190 B.n800 B.n378 585
R191 B.n378 B.n377 585
R192 B.n799 B.n798 585
R193 B.n798 B.n797 585
R194 B.n380 B.n379 585
R195 B.n381 B.n380 585
R196 B.n790 B.n789 585
R197 B.n791 B.n790 585
R198 B.n788 B.n386 585
R199 B.n386 B.n385 585
R200 B.n787 B.n786 585
R201 B.n786 B.n785 585
R202 B.n388 B.n387 585
R203 B.n389 B.n388 585
R204 B.n778 B.n777 585
R205 B.n779 B.n778 585
R206 B.n776 B.n394 585
R207 B.n394 B.n393 585
R208 B.n775 B.n774 585
R209 B.n774 B.n773 585
R210 B.n396 B.n395 585
R211 B.n397 B.n396 585
R212 B.n766 B.n765 585
R213 B.n767 B.n766 585
R214 B.n764 B.n402 585
R215 B.n402 B.n401 585
R216 B.n763 B.n762 585
R217 B.n762 B.n761 585
R218 B.n404 B.n403 585
R219 B.n405 B.n404 585
R220 B.n754 B.n753 585
R221 B.n755 B.n754 585
R222 B.n752 B.n410 585
R223 B.n410 B.n409 585
R224 B.n751 B.n750 585
R225 B.n750 B.n749 585
R226 B.n412 B.n411 585
R227 B.n413 B.n412 585
R228 B.n745 B.n744 585
R229 B.n416 B.n415 585
R230 B.n741 B.n740 585
R231 B.n742 B.n741 585
R232 B.n739 B.n481 585
R233 B.n738 B.n737 585
R234 B.n736 B.n735 585
R235 B.n734 B.n733 585
R236 B.n732 B.n731 585
R237 B.n730 B.n729 585
R238 B.n728 B.n727 585
R239 B.n726 B.n725 585
R240 B.n724 B.n723 585
R241 B.n722 B.n721 585
R242 B.n720 B.n719 585
R243 B.n718 B.n717 585
R244 B.n716 B.n715 585
R245 B.n714 B.n713 585
R246 B.n712 B.n711 585
R247 B.n710 B.n709 585
R248 B.n708 B.n707 585
R249 B.n706 B.n705 585
R250 B.n704 B.n703 585
R251 B.n702 B.n701 585
R252 B.n700 B.n699 585
R253 B.n698 B.n697 585
R254 B.n696 B.n695 585
R255 B.n694 B.n693 585
R256 B.n692 B.n691 585
R257 B.n690 B.n689 585
R258 B.n688 B.n687 585
R259 B.n686 B.n685 585
R260 B.n684 B.n683 585
R261 B.n682 B.n681 585
R262 B.n680 B.n679 585
R263 B.n678 B.n677 585
R264 B.n676 B.n675 585
R265 B.n674 B.n673 585
R266 B.n672 B.n671 585
R267 B.n670 B.n669 585
R268 B.n668 B.n667 585
R269 B.n666 B.n665 585
R270 B.n664 B.n663 585
R271 B.n662 B.n661 585
R272 B.n660 B.n659 585
R273 B.n658 B.n657 585
R274 B.n656 B.n655 585
R275 B.n654 B.n653 585
R276 B.n652 B.n651 585
R277 B.n650 B.n649 585
R278 B.n648 B.n647 585
R279 B.n646 B.n645 585
R280 B.n644 B.n643 585
R281 B.n642 B.n641 585
R282 B.n640 B.n639 585
R283 B.n638 B.n637 585
R284 B.n636 B.n635 585
R285 B.n634 B.n633 585
R286 B.n632 B.n631 585
R287 B.n630 B.n629 585
R288 B.n628 B.n627 585
R289 B.n625 B.n624 585
R290 B.n623 B.n622 585
R291 B.n621 B.n620 585
R292 B.n619 B.n618 585
R293 B.n617 B.n616 585
R294 B.n615 B.n614 585
R295 B.n613 B.n612 585
R296 B.n611 B.n610 585
R297 B.n609 B.n608 585
R298 B.n607 B.n606 585
R299 B.n604 B.n603 585
R300 B.n602 B.n601 585
R301 B.n600 B.n599 585
R302 B.n598 B.n597 585
R303 B.n596 B.n595 585
R304 B.n594 B.n593 585
R305 B.n592 B.n591 585
R306 B.n590 B.n589 585
R307 B.n588 B.n587 585
R308 B.n586 B.n585 585
R309 B.n584 B.n583 585
R310 B.n582 B.n581 585
R311 B.n580 B.n579 585
R312 B.n578 B.n577 585
R313 B.n576 B.n575 585
R314 B.n574 B.n573 585
R315 B.n572 B.n571 585
R316 B.n570 B.n569 585
R317 B.n568 B.n567 585
R318 B.n566 B.n565 585
R319 B.n564 B.n563 585
R320 B.n562 B.n561 585
R321 B.n560 B.n559 585
R322 B.n558 B.n557 585
R323 B.n556 B.n555 585
R324 B.n554 B.n553 585
R325 B.n552 B.n551 585
R326 B.n550 B.n549 585
R327 B.n548 B.n547 585
R328 B.n546 B.n545 585
R329 B.n544 B.n543 585
R330 B.n542 B.n541 585
R331 B.n540 B.n539 585
R332 B.n538 B.n537 585
R333 B.n536 B.n535 585
R334 B.n534 B.n533 585
R335 B.n532 B.n531 585
R336 B.n530 B.n529 585
R337 B.n528 B.n527 585
R338 B.n526 B.n525 585
R339 B.n524 B.n523 585
R340 B.n522 B.n521 585
R341 B.n520 B.n519 585
R342 B.n518 B.n517 585
R343 B.n516 B.n515 585
R344 B.n514 B.n513 585
R345 B.n512 B.n511 585
R346 B.n510 B.n509 585
R347 B.n508 B.n507 585
R348 B.n506 B.n505 585
R349 B.n504 B.n503 585
R350 B.n502 B.n501 585
R351 B.n500 B.n499 585
R352 B.n498 B.n497 585
R353 B.n496 B.n495 585
R354 B.n494 B.n493 585
R355 B.n492 B.n491 585
R356 B.n490 B.n489 585
R357 B.n488 B.n487 585
R358 B.n486 B.n480 585
R359 B.n742 B.n480 585
R360 B.n746 B.n414 585
R361 B.n414 B.n413 585
R362 B.n748 B.n747 585
R363 B.n749 B.n748 585
R364 B.n408 B.n407 585
R365 B.n409 B.n408 585
R366 B.n757 B.n756 585
R367 B.n756 B.n755 585
R368 B.n758 B.n406 585
R369 B.n406 B.n405 585
R370 B.n760 B.n759 585
R371 B.n761 B.n760 585
R372 B.n400 B.n399 585
R373 B.n401 B.n400 585
R374 B.n769 B.n768 585
R375 B.n768 B.n767 585
R376 B.n770 B.n398 585
R377 B.n398 B.n397 585
R378 B.n772 B.n771 585
R379 B.n773 B.n772 585
R380 B.n392 B.n391 585
R381 B.n393 B.n392 585
R382 B.n781 B.n780 585
R383 B.n780 B.n779 585
R384 B.n782 B.n390 585
R385 B.n390 B.n389 585
R386 B.n784 B.n783 585
R387 B.n785 B.n784 585
R388 B.n384 B.n383 585
R389 B.n385 B.n384 585
R390 B.n793 B.n792 585
R391 B.n792 B.n791 585
R392 B.n794 B.n382 585
R393 B.n382 B.n381 585
R394 B.n796 B.n795 585
R395 B.n797 B.n796 585
R396 B.n376 B.n375 585
R397 B.n377 B.n376 585
R398 B.n806 B.n805 585
R399 B.n805 B.n804 585
R400 B.n807 B.n374 585
R401 B.n374 B.n373 585
R402 B.n809 B.n808 585
R403 B.n810 B.n809 585
R404 B.n2 B.n0 585
R405 B.n4 B.n2 585
R406 B.n3 B.n1 585
R407 B.n894 B.n3 585
R408 B.n892 B.n891 585
R409 B.n893 B.n892 585
R410 B.n890 B.n9 585
R411 B.n9 B.n8 585
R412 B.n889 B.n888 585
R413 B.n888 B.n887 585
R414 B.n11 B.n10 585
R415 B.n886 B.n11 585
R416 B.n884 B.n883 585
R417 B.n885 B.n884 585
R418 B.n882 B.n16 585
R419 B.n16 B.n15 585
R420 B.n881 B.n880 585
R421 B.n880 B.n879 585
R422 B.n18 B.n17 585
R423 B.n878 B.n18 585
R424 B.n876 B.n875 585
R425 B.n877 B.n876 585
R426 B.n874 B.n23 585
R427 B.n23 B.n22 585
R428 B.n873 B.n872 585
R429 B.n872 B.n871 585
R430 B.n25 B.n24 585
R431 B.n870 B.n25 585
R432 B.n868 B.n867 585
R433 B.n869 B.n868 585
R434 B.n866 B.n30 585
R435 B.n30 B.n29 585
R436 B.n865 B.n864 585
R437 B.n864 B.n863 585
R438 B.n32 B.n31 585
R439 B.n862 B.n32 585
R440 B.n860 B.n859 585
R441 B.n861 B.n860 585
R442 B.n858 B.n37 585
R443 B.n37 B.n36 585
R444 B.n857 B.n856 585
R445 B.n856 B.n855 585
R446 B.n39 B.n38 585
R447 B.n854 B.n39 585
R448 B.n852 B.n851 585
R449 B.n853 B.n852 585
R450 B.n850 B.n44 585
R451 B.n44 B.n43 585
R452 B.n897 B.n896 585
R453 B.n896 B.n895 585
R454 B.n744 B.n414 530.939
R455 B.n848 B.n44 530.939
R456 B.n480 B.n412 530.939
R457 B.n844 B.n111 530.939
R458 B.n484 B.t19 416.317
R459 B.n112 B.t11 416.317
R460 B.n482 B.t16 416.317
R461 B.n115 B.t8 416.317
R462 B.n485 B.t18 391.493
R463 B.n113 B.t12 391.493
R464 B.n483 B.t15 391.493
R465 B.n116 B.t9 391.493
R466 B.n846 B.n845 256.663
R467 B.n846 B.n109 256.663
R468 B.n846 B.n108 256.663
R469 B.n846 B.n107 256.663
R470 B.n846 B.n106 256.663
R471 B.n846 B.n105 256.663
R472 B.n846 B.n104 256.663
R473 B.n846 B.n103 256.663
R474 B.n846 B.n102 256.663
R475 B.n846 B.n101 256.663
R476 B.n846 B.n100 256.663
R477 B.n846 B.n99 256.663
R478 B.n846 B.n98 256.663
R479 B.n846 B.n97 256.663
R480 B.n846 B.n96 256.663
R481 B.n846 B.n95 256.663
R482 B.n846 B.n94 256.663
R483 B.n846 B.n93 256.663
R484 B.n846 B.n92 256.663
R485 B.n846 B.n91 256.663
R486 B.n846 B.n90 256.663
R487 B.n846 B.n89 256.663
R488 B.n846 B.n88 256.663
R489 B.n846 B.n87 256.663
R490 B.n846 B.n86 256.663
R491 B.n846 B.n85 256.663
R492 B.n846 B.n84 256.663
R493 B.n846 B.n83 256.663
R494 B.n846 B.n82 256.663
R495 B.n846 B.n81 256.663
R496 B.n846 B.n80 256.663
R497 B.n846 B.n79 256.663
R498 B.n846 B.n78 256.663
R499 B.n846 B.n77 256.663
R500 B.n846 B.n76 256.663
R501 B.n846 B.n75 256.663
R502 B.n846 B.n74 256.663
R503 B.n846 B.n73 256.663
R504 B.n846 B.n72 256.663
R505 B.n846 B.n71 256.663
R506 B.n846 B.n70 256.663
R507 B.n846 B.n69 256.663
R508 B.n846 B.n68 256.663
R509 B.n846 B.n67 256.663
R510 B.n846 B.n66 256.663
R511 B.n846 B.n65 256.663
R512 B.n846 B.n64 256.663
R513 B.n846 B.n63 256.663
R514 B.n846 B.n62 256.663
R515 B.n846 B.n61 256.663
R516 B.n846 B.n60 256.663
R517 B.n846 B.n59 256.663
R518 B.n846 B.n58 256.663
R519 B.n846 B.n57 256.663
R520 B.n846 B.n56 256.663
R521 B.n846 B.n55 256.663
R522 B.n846 B.n54 256.663
R523 B.n846 B.n53 256.663
R524 B.n846 B.n52 256.663
R525 B.n846 B.n51 256.663
R526 B.n846 B.n50 256.663
R527 B.n846 B.n49 256.663
R528 B.n846 B.n48 256.663
R529 B.n846 B.n47 256.663
R530 B.n847 B.n846 256.663
R531 B.n743 B.n742 256.663
R532 B.n742 B.n417 256.663
R533 B.n742 B.n418 256.663
R534 B.n742 B.n419 256.663
R535 B.n742 B.n420 256.663
R536 B.n742 B.n421 256.663
R537 B.n742 B.n422 256.663
R538 B.n742 B.n423 256.663
R539 B.n742 B.n424 256.663
R540 B.n742 B.n425 256.663
R541 B.n742 B.n426 256.663
R542 B.n742 B.n427 256.663
R543 B.n742 B.n428 256.663
R544 B.n742 B.n429 256.663
R545 B.n742 B.n430 256.663
R546 B.n742 B.n431 256.663
R547 B.n742 B.n432 256.663
R548 B.n742 B.n433 256.663
R549 B.n742 B.n434 256.663
R550 B.n742 B.n435 256.663
R551 B.n742 B.n436 256.663
R552 B.n742 B.n437 256.663
R553 B.n742 B.n438 256.663
R554 B.n742 B.n439 256.663
R555 B.n742 B.n440 256.663
R556 B.n742 B.n441 256.663
R557 B.n742 B.n442 256.663
R558 B.n742 B.n443 256.663
R559 B.n742 B.n444 256.663
R560 B.n742 B.n445 256.663
R561 B.n742 B.n446 256.663
R562 B.n742 B.n447 256.663
R563 B.n742 B.n448 256.663
R564 B.n742 B.n449 256.663
R565 B.n742 B.n450 256.663
R566 B.n742 B.n451 256.663
R567 B.n742 B.n452 256.663
R568 B.n742 B.n453 256.663
R569 B.n742 B.n454 256.663
R570 B.n742 B.n455 256.663
R571 B.n742 B.n456 256.663
R572 B.n742 B.n457 256.663
R573 B.n742 B.n458 256.663
R574 B.n742 B.n459 256.663
R575 B.n742 B.n460 256.663
R576 B.n742 B.n461 256.663
R577 B.n742 B.n462 256.663
R578 B.n742 B.n463 256.663
R579 B.n742 B.n464 256.663
R580 B.n742 B.n465 256.663
R581 B.n742 B.n466 256.663
R582 B.n742 B.n467 256.663
R583 B.n742 B.n468 256.663
R584 B.n742 B.n469 256.663
R585 B.n742 B.n470 256.663
R586 B.n742 B.n471 256.663
R587 B.n742 B.n472 256.663
R588 B.n742 B.n473 256.663
R589 B.n742 B.n474 256.663
R590 B.n742 B.n475 256.663
R591 B.n742 B.n476 256.663
R592 B.n742 B.n477 256.663
R593 B.n742 B.n478 256.663
R594 B.n742 B.n479 256.663
R595 B.n748 B.n414 163.367
R596 B.n748 B.n408 163.367
R597 B.n756 B.n408 163.367
R598 B.n756 B.n406 163.367
R599 B.n760 B.n406 163.367
R600 B.n760 B.n400 163.367
R601 B.n768 B.n400 163.367
R602 B.n768 B.n398 163.367
R603 B.n772 B.n398 163.367
R604 B.n772 B.n392 163.367
R605 B.n780 B.n392 163.367
R606 B.n780 B.n390 163.367
R607 B.n784 B.n390 163.367
R608 B.n784 B.n384 163.367
R609 B.n792 B.n384 163.367
R610 B.n792 B.n382 163.367
R611 B.n796 B.n382 163.367
R612 B.n796 B.n376 163.367
R613 B.n805 B.n376 163.367
R614 B.n805 B.n374 163.367
R615 B.n809 B.n374 163.367
R616 B.n809 B.n2 163.367
R617 B.n896 B.n2 163.367
R618 B.n896 B.n3 163.367
R619 B.n892 B.n3 163.367
R620 B.n892 B.n9 163.367
R621 B.n888 B.n9 163.367
R622 B.n888 B.n11 163.367
R623 B.n884 B.n11 163.367
R624 B.n884 B.n16 163.367
R625 B.n880 B.n16 163.367
R626 B.n880 B.n18 163.367
R627 B.n876 B.n18 163.367
R628 B.n876 B.n23 163.367
R629 B.n872 B.n23 163.367
R630 B.n872 B.n25 163.367
R631 B.n868 B.n25 163.367
R632 B.n868 B.n30 163.367
R633 B.n864 B.n30 163.367
R634 B.n864 B.n32 163.367
R635 B.n860 B.n32 163.367
R636 B.n860 B.n37 163.367
R637 B.n856 B.n37 163.367
R638 B.n856 B.n39 163.367
R639 B.n852 B.n39 163.367
R640 B.n852 B.n44 163.367
R641 B.n741 B.n416 163.367
R642 B.n741 B.n481 163.367
R643 B.n737 B.n736 163.367
R644 B.n733 B.n732 163.367
R645 B.n729 B.n728 163.367
R646 B.n725 B.n724 163.367
R647 B.n721 B.n720 163.367
R648 B.n717 B.n716 163.367
R649 B.n713 B.n712 163.367
R650 B.n709 B.n708 163.367
R651 B.n705 B.n704 163.367
R652 B.n701 B.n700 163.367
R653 B.n697 B.n696 163.367
R654 B.n693 B.n692 163.367
R655 B.n689 B.n688 163.367
R656 B.n685 B.n684 163.367
R657 B.n681 B.n680 163.367
R658 B.n677 B.n676 163.367
R659 B.n673 B.n672 163.367
R660 B.n669 B.n668 163.367
R661 B.n665 B.n664 163.367
R662 B.n661 B.n660 163.367
R663 B.n657 B.n656 163.367
R664 B.n653 B.n652 163.367
R665 B.n649 B.n648 163.367
R666 B.n645 B.n644 163.367
R667 B.n641 B.n640 163.367
R668 B.n637 B.n636 163.367
R669 B.n633 B.n632 163.367
R670 B.n629 B.n628 163.367
R671 B.n624 B.n623 163.367
R672 B.n620 B.n619 163.367
R673 B.n616 B.n615 163.367
R674 B.n612 B.n611 163.367
R675 B.n608 B.n607 163.367
R676 B.n603 B.n602 163.367
R677 B.n599 B.n598 163.367
R678 B.n595 B.n594 163.367
R679 B.n591 B.n590 163.367
R680 B.n587 B.n586 163.367
R681 B.n583 B.n582 163.367
R682 B.n579 B.n578 163.367
R683 B.n575 B.n574 163.367
R684 B.n571 B.n570 163.367
R685 B.n567 B.n566 163.367
R686 B.n563 B.n562 163.367
R687 B.n559 B.n558 163.367
R688 B.n555 B.n554 163.367
R689 B.n551 B.n550 163.367
R690 B.n547 B.n546 163.367
R691 B.n543 B.n542 163.367
R692 B.n539 B.n538 163.367
R693 B.n535 B.n534 163.367
R694 B.n531 B.n530 163.367
R695 B.n527 B.n526 163.367
R696 B.n523 B.n522 163.367
R697 B.n519 B.n518 163.367
R698 B.n515 B.n514 163.367
R699 B.n511 B.n510 163.367
R700 B.n507 B.n506 163.367
R701 B.n503 B.n502 163.367
R702 B.n499 B.n498 163.367
R703 B.n495 B.n494 163.367
R704 B.n491 B.n490 163.367
R705 B.n487 B.n480 163.367
R706 B.n750 B.n412 163.367
R707 B.n750 B.n410 163.367
R708 B.n754 B.n410 163.367
R709 B.n754 B.n404 163.367
R710 B.n762 B.n404 163.367
R711 B.n762 B.n402 163.367
R712 B.n766 B.n402 163.367
R713 B.n766 B.n396 163.367
R714 B.n774 B.n396 163.367
R715 B.n774 B.n394 163.367
R716 B.n778 B.n394 163.367
R717 B.n778 B.n388 163.367
R718 B.n786 B.n388 163.367
R719 B.n786 B.n386 163.367
R720 B.n790 B.n386 163.367
R721 B.n790 B.n380 163.367
R722 B.n798 B.n380 163.367
R723 B.n798 B.n378 163.367
R724 B.n803 B.n378 163.367
R725 B.n803 B.n372 163.367
R726 B.n811 B.n372 163.367
R727 B.n812 B.n811 163.367
R728 B.n812 B.n5 163.367
R729 B.n6 B.n5 163.367
R730 B.n7 B.n6 163.367
R731 B.n817 B.n7 163.367
R732 B.n817 B.n12 163.367
R733 B.n13 B.n12 163.367
R734 B.n14 B.n13 163.367
R735 B.n822 B.n14 163.367
R736 B.n822 B.n19 163.367
R737 B.n20 B.n19 163.367
R738 B.n21 B.n20 163.367
R739 B.n827 B.n21 163.367
R740 B.n827 B.n26 163.367
R741 B.n27 B.n26 163.367
R742 B.n28 B.n27 163.367
R743 B.n832 B.n28 163.367
R744 B.n832 B.n33 163.367
R745 B.n34 B.n33 163.367
R746 B.n35 B.n34 163.367
R747 B.n837 B.n35 163.367
R748 B.n837 B.n40 163.367
R749 B.n41 B.n40 163.367
R750 B.n42 B.n41 163.367
R751 B.n111 B.n42 163.367
R752 B.n118 B.n46 163.367
R753 B.n122 B.n121 163.367
R754 B.n126 B.n125 163.367
R755 B.n130 B.n129 163.367
R756 B.n134 B.n133 163.367
R757 B.n138 B.n137 163.367
R758 B.n142 B.n141 163.367
R759 B.n146 B.n145 163.367
R760 B.n150 B.n149 163.367
R761 B.n154 B.n153 163.367
R762 B.n158 B.n157 163.367
R763 B.n162 B.n161 163.367
R764 B.n166 B.n165 163.367
R765 B.n170 B.n169 163.367
R766 B.n174 B.n173 163.367
R767 B.n178 B.n177 163.367
R768 B.n182 B.n181 163.367
R769 B.n186 B.n185 163.367
R770 B.n190 B.n189 163.367
R771 B.n194 B.n193 163.367
R772 B.n198 B.n197 163.367
R773 B.n202 B.n201 163.367
R774 B.n206 B.n205 163.367
R775 B.n210 B.n209 163.367
R776 B.n214 B.n213 163.367
R777 B.n218 B.n217 163.367
R778 B.n222 B.n221 163.367
R779 B.n226 B.n225 163.367
R780 B.n230 B.n229 163.367
R781 B.n234 B.n233 163.367
R782 B.n238 B.n237 163.367
R783 B.n242 B.n241 163.367
R784 B.n246 B.n245 163.367
R785 B.n250 B.n249 163.367
R786 B.n254 B.n253 163.367
R787 B.n258 B.n257 163.367
R788 B.n262 B.n261 163.367
R789 B.n266 B.n265 163.367
R790 B.n270 B.n269 163.367
R791 B.n274 B.n273 163.367
R792 B.n278 B.n277 163.367
R793 B.n282 B.n281 163.367
R794 B.n286 B.n285 163.367
R795 B.n290 B.n289 163.367
R796 B.n294 B.n293 163.367
R797 B.n298 B.n297 163.367
R798 B.n302 B.n301 163.367
R799 B.n306 B.n305 163.367
R800 B.n310 B.n309 163.367
R801 B.n314 B.n313 163.367
R802 B.n318 B.n317 163.367
R803 B.n322 B.n321 163.367
R804 B.n326 B.n325 163.367
R805 B.n330 B.n329 163.367
R806 B.n334 B.n333 163.367
R807 B.n338 B.n337 163.367
R808 B.n342 B.n341 163.367
R809 B.n346 B.n345 163.367
R810 B.n350 B.n349 163.367
R811 B.n354 B.n353 163.367
R812 B.n358 B.n357 163.367
R813 B.n362 B.n361 163.367
R814 B.n366 B.n365 163.367
R815 B.n368 B.n110 163.367
R816 B.n744 B.n743 71.676
R817 B.n481 B.n417 71.676
R818 B.n736 B.n418 71.676
R819 B.n732 B.n419 71.676
R820 B.n728 B.n420 71.676
R821 B.n724 B.n421 71.676
R822 B.n720 B.n422 71.676
R823 B.n716 B.n423 71.676
R824 B.n712 B.n424 71.676
R825 B.n708 B.n425 71.676
R826 B.n704 B.n426 71.676
R827 B.n700 B.n427 71.676
R828 B.n696 B.n428 71.676
R829 B.n692 B.n429 71.676
R830 B.n688 B.n430 71.676
R831 B.n684 B.n431 71.676
R832 B.n680 B.n432 71.676
R833 B.n676 B.n433 71.676
R834 B.n672 B.n434 71.676
R835 B.n668 B.n435 71.676
R836 B.n664 B.n436 71.676
R837 B.n660 B.n437 71.676
R838 B.n656 B.n438 71.676
R839 B.n652 B.n439 71.676
R840 B.n648 B.n440 71.676
R841 B.n644 B.n441 71.676
R842 B.n640 B.n442 71.676
R843 B.n636 B.n443 71.676
R844 B.n632 B.n444 71.676
R845 B.n628 B.n445 71.676
R846 B.n623 B.n446 71.676
R847 B.n619 B.n447 71.676
R848 B.n615 B.n448 71.676
R849 B.n611 B.n449 71.676
R850 B.n607 B.n450 71.676
R851 B.n602 B.n451 71.676
R852 B.n598 B.n452 71.676
R853 B.n594 B.n453 71.676
R854 B.n590 B.n454 71.676
R855 B.n586 B.n455 71.676
R856 B.n582 B.n456 71.676
R857 B.n578 B.n457 71.676
R858 B.n574 B.n458 71.676
R859 B.n570 B.n459 71.676
R860 B.n566 B.n460 71.676
R861 B.n562 B.n461 71.676
R862 B.n558 B.n462 71.676
R863 B.n554 B.n463 71.676
R864 B.n550 B.n464 71.676
R865 B.n546 B.n465 71.676
R866 B.n542 B.n466 71.676
R867 B.n538 B.n467 71.676
R868 B.n534 B.n468 71.676
R869 B.n530 B.n469 71.676
R870 B.n526 B.n470 71.676
R871 B.n522 B.n471 71.676
R872 B.n518 B.n472 71.676
R873 B.n514 B.n473 71.676
R874 B.n510 B.n474 71.676
R875 B.n506 B.n475 71.676
R876 B.n502 B.n476 71.676
R877 B.n498 B.n477 71.676
R878 B.n494 B.n478 71.676
R879 B.n490 B.n479 71.676
R880 B.n848 B.n847 71.676
R881 B.n118 B.n47 71.676
R882 B.n122 B.n48 71.676
R883 B.n126 B.n49 71.676
R884 B.n130 B.n50 71.676
R885 B.n134 B.n51 71.676
R886 B.n138 B.n52 71.676
R887 B.n142 B.n53 71.676
R888 B.n146 B.n54 71.676
R889 B.n150 B.n55 71.676
R890 B.n154 B.n56 71.676
R891 B.n158 B.n57 71.676
R892 B.n162 B.n58 71.676
R893 B.n166 B.n59 71.676
R894 B.n170 B.n60 71.676
R895 B.n174 B.n61 71.676
R896 B.n178 B.n62 71.676
R897 B.n182 B.n63 71.676
R898 B.n186 B.n64 71.676
R899 B.n190 B.n65 71.676
R900 B.n194 B.n66 71.676
R901 B.n198 B.n67 71.676
R902 B.n202 B.n68 71.676
R903 B.n206 B.n69 71.676
R904 B.n210 B.n70 71.676
R905 B.n214 B.n71 71.676
R906 B.n218 B.n72 71.676
R907 B.n222 B.n73 71.676
R908 B.n226 B.n74 71.676
R909 B.n230 B.n75 71.676
R910 B.n234 B.n76 71.676
R911 B.n238 B.n77 71.676
R912 B.n242 B.n78 71.676
R913 B.n246 B.n79 71.676
R914 B.n250 B.n80 71.676
R915 B.n254 B.n81 71.676
R916 B.n258 B.n82 71.676
R917 B.n262 B.n83 71.676
R918 B.n266 B.n84 71.676
R919 B.n270 B.n85 71.676
R920 B.n274 B.n86 71.676
R921 B.n278 B.n87 71.676
R922 B.n282 B.n88 71.676
R923 B.n286 B.n89 71.676
R924 B.n290 B.n90 71.676
R925 B.n294 B.n91 71.676
R926 B.n298 B.n92 71.676
R927 B.n302 B.n93 71.676
R928 B.n306 B.n94 71.676
R929 B.n310 B.n95 71.676
R930 B.n314 B.n96 71.676
R931 B.n318 B.n97 71.676
R932 B.n322 B.n98 71.676
R933 B.n326 B.n99 71.676
R934 B.n330 B.n100 71.676
R935 B.n334 B.n101 71.676
R936 B.n338 B.n102 71.676
R937 B.n342 B.n103 71.676
R938 B.n346 B.n104 71.676
R939 B.n350 B.n105 71.676
R940 B.n354 B.n106 71.676
R941 B.n358 B.n107 71.676
R942 B.n362 B.n108 71.676
R943 B.n366 B.n109 71.676
R944 B.n845 B.n110 71.676
R945 B.n845 B.n844 71.676
R946 B.n368 B.n109 71.676
R947 B.n365 B.n108 71.676
R948 B.n361 B.n107 71.676
R949 B.n357 B.n106 71.676
R950 B.n353 B.n105 71.676
R951 B.n349 B.n104 71.676
R952 B.n345 B.n103 71.676
R953 B.n341 B.n102 71.676
R954 B.n337 B.n101 71.676
R955 B.n333 B.n100 71.676
R956 B.n329 B.n99 71.676
R957 B.n325 B.n98 71.676
R958 B.n321 B.n97 71.676
R959 B.n317 B.n96 71.676
R960 B.n313 B.n95 71.676
R961 B.n309 B.n94 71.676
R962 B.n305 B.n93 71.676
R963 B.n301 B.n92 71.676
R964 B.n297 B.n91 71.676
R965 B.n293 B.n90 71.676
R966 B.n289 B.n89 71.676
R967 B.n285 B.n88 71.676
R968 B.n281 B.n87 71.676
R969 B.n277 B.n86 71.676
R970 B.n273 B.n85 71.676
R971 B.n269 B.n84 71.676
R972 B.n265 B.n83 71.676
R973 B.n261 B.n82 71.676
R974 B.n257 B.n81 71.676
R975 B.n253 B.n80 71.676
R976 B.n249 B.n79 71.676
R977 B.n245 B.n78 71.676
R978 B.n241 B.n77 71.676
R979 B.n237 B.n76 71.676
R980 B.n233 B.n75 71.676
R981 B.n229 B.n74 71.676
R982 B.n225 B.n73 71.676
R983 B.n221 B.n72 71.676
R984 B.n217 B.n71 71.676
R985 B.n213 B.n70 71.676
R986 B.n209 B.n69 71.676
R987 B.n205 B.n68 71.676
R988 B.n201 B.n67 71.676
R989 B.n197 B.n66 71.676
R990 B.n193 B.n65 71.676
R991 B.n189 B.n64 71.676
R992 B.n185 B.n63 71.676
R993 B.n181 B.n62 71.676
R994 B.n177 B.n61 71.676
R995 B.n173 B.n60 71.676
R996 B.n169 B.n59 71.676
R997 B.n165 B.n58 71.676
R998 B.n161 B.n57 71.676
R999 B.n157 B.n56 71.676
R1000 B.n153 B.n55 71.676
R1001 B.n149 B.n54 71.676
R1002 B.n145 B.n53 71.676
R1003 B.n141 B.n52 71.676
R1004 B.n137 B.n51 71.676
R1005 B.n133 B.n50 71.676
R1006 B.n129 B.n49 71.676
R1007 B.n125 B.n48 71.676
R1008 B.n121 B.n47 71.676
R1009 B.n847 B.n46 71.676
R1010 B.n743 B.n416 71.676
R1011 B.n737 B.n417 71.676
R1012 B.n733 B.n418 71.676
R1013 B.n729 B.n419 71.676
R1014 B.n725 B.n420 71.676
R1015 B.n721 B.n421 71.676
R1016 B.n717 B.n422 71.676
R1017 B.n713 B.n423 71.676
R1018 B.n709 B.n424 71.676
R1019 B.n705 B.n425 71.676
R1020 B.n701 B.n426 71.676
R1021 B.n697 B.n427 71.676
R1022 B.n693 B.n428 71.676
R1023 B.n689 B.n429 71.676
R1024 B.n685 B.n430 71.676
R1025 B.n681 B.n431 71.676
R1026 B.n677 B.n432 71.676
R1027 B.n673 B.n433 71.676
R1028 B.n669 B.n434 71.676
R1029 B.n665 B.n435 71.676
R1030 B.n661 B.n436 71.676
R1031 B.n657 B.n437 71.676
R1032 B.n653 B.n438 71.676
R1033 B.n649 B.n439 71.676
R1034 B.n645 B.n440 71.676
R1035 B.n641 B.n441 71.676
R1036 B.n637 B.n442 71.676
R1037 B.n633 B.n443 71.676
R1038 B.n629 B.n444 71.676
R1039 B.n624 B.n445 71.676
R1040 B.n620 B.n446 71.676
R1041 B.n616 B.n447 71.676
R1042 B.n612 B.n448 71.676
R1043 B.n608 B.n449 71.676
R1044 B.n603 B.n450 71.676
R1045 B.n599 B.n451 71.676
R1046 B.n595 B.n452 71.676
R1047 B.n591 B.n453 71.676
R1048 B.n587 B.n454 71.676
R1049 B.n583 B.n455 71.676
R1050 B.n579 B.n456 71.676
R1051 B.n575 B.n457 71.676
R1052 B.n571 B.n458 71.676
R1053 B.n567 B.n459 71.676
R1054 B.n563 B.n460 71.676
R1055 B.n559 B.n461 71.676
R1056 B.n555 B.n462 71.676
R1057 B.n551 B.n463 71.676
R1058 B.n547 B.n464 71.676
R1059 B.n543 B.n465 71.676
R1060 B.n539 B.n466 71.676
R1061 B.n535 B.n467 71.676
R1062 B.n531 B.n468 71.676
R1063 B.n527 B.n469 71.676
R1064 B.n523 B.n470 71.676
R1065 B.n519 B.n471 71.676
R1066 B.n515 B.n472 71.676
R1067 B.n511 B.n473 71.676
R1068 B.n507 B.n474 71.676
R1069 B.n503 B.n475 71.676
R1070 B.n499 B.n476 71.676
R1071 B.n495 B.n477 71.676
R1072 B.n491 B.n478 71.676
R1073 B.n487 B.n479 71.676
R1074 B.n742 B.n413 62.9109
R1075 B.n846 B.n43 62.9109
R1076 B.n605 B.n485 59.5399
R1077 B.n626 B.n483 59.5399
R1078 B.n117 B.n116 59.5399
R1079 B.n114 B.n113 59.5399
R1080 B.n850 B.n849 34.4981
R1081 B.n843 B.n842 34.4981
R1082 B.n486 B.n411 34.4981
R1083 B.n746 B.n745 34.4981
R1084 B.n749 B.n413 31.6887
R1085 B.n749 B.n409 31.6887
R1086 B.n755 B.n409 31.6887
R1087 B.n755 B.n405 31.6887
R1088 B.n761 B.n405 31.6887
R1089 B.n767 B.n401 31.6887
R1090 B.n767 B.n397 31.6887
R1091 B.n773 B.n397 31.6887
R1092 B.n773 B.n393 31.6887
R1093 B.n779 B.n393 31.6887
R1094 B.n785 B.n389 31.6887
R1095 B.n785 B.n385 31.6887
R1096 B.n791 B.n385 31.6887
R1097 B.n797 B.n381 31.6887
R1098 B.n797 B.n377 31.6887
R1099 B.n804 B.n377 31.6887
R1100 B.n810 B.n373 31.6887
R1101 B.n810 B.n4 31.6887
R1102 B.n895 B.n4 31.6887
R1103 B.n895 B.n894 31.6887
R1104 B.n894 B.n893 31.6887
R1105 B.n893 B.n8 31.6887
R1106 B.n887 B.n886 31.6887
R1107 B.n886 B.n885 31.6887
R1108 B.n885 B.n15 31.6887
R1109 B.n879 B.n878 31.6887
R1110 B.n878 B.n877 31.6887
R1111 B.n877 B.n22 31.6887
R1112 B.n871 B.n870 31.6887
R1113 B.n870 B.n869 31.6887
R1114 B.n869 B.n29 31.6887
R1115 B.n863 B.n29 31.6887
R1116 B.n863 B.n862 31.6887
R1117 B.n861 B.n36 31.6887
R1118 B.n855 B.n36 31.6887
R1119 B.n855 B.n854 31.6887
R1120 B.n854 B.n853 31.6887
R1121 B.n853 B.n43 31.6887
R1122 B.t14 B.n401 31.2227
R1123 B.n779 B.t3 31.2227
R1124 B.n871 B.t0 31.2227
R1125 B.n862 B.t7 31.2227
R1126 B.n485 B.n484 24.8247
R1127 B.n483 B.n482 24.8247
R1128 B.n116 B.n115 24.8247
R1129 B.n113 B.n112 24.8247
R1130 B.n791 B.t5 23.7666
R1131 B.n879 B.t4 23.7666
R1132 B B.n897 18.0485
R1133 B.n804 B.t2 16.3106
R1134 B.n887 B.t1 16.3106
R1135 B.t2 B.n373 15.3786
R1136 B.t1 B.n8 15.3786
R1137 B.n849 B.n45 10.6151
R1138 B.n119 B.n45 10.6151
R1139 B.n120 B.n119 10.6151
R1140 B.n123 B.n120 10.6151
R1141 B.n124 B.n123 10.6151
R1142 B.n127 B.n124 10.6151
R1143 B.n128 B.n127 10.6151
R1144 B.n131 B.n128 10.6151
R1145 B.n132 B.n131 10.6151
R1146 B.n135 B.n132 10.6151
R1147 B.n136 B.n135 10.6151
R1148 B.n139 B.n136 10.6151
R1149 B.n140 B.n139 10.6151
R1150 B.n143 B.n140 10.6151
R1151 B.n144 B.n143 10.6151
R1152 B.n147 B.n144 10.6151
R1153 B.n148 B.n147 10.6151
R1154 B.n151 B.n148 10.6151
R1155 B.n152 B.n151 10.6151
R1156 B.n155 B.n152 10.6151
R1157 B.n156 B.n155 10.6151
R1158 B.n159 B.n156 10.6151
R1159 B.n160 B.n159 10.6151
R1160 B.n163 B.n160 10.6151
R1161 B.n164 B.n163 10.6151
R1162 B.n167 B.n164 10.6151
R1163 B.n168 B.n167 10.6151
R1164 B.n171 B.n168 10.6151
R1165 B.n172 B.n171 10.6151
R1166 B.n175 B.n172 10.6151
R1167 B.n176 B.n175 10.6151
R1168 B.n179 B.n176 10.6151
R1169 B.n180 B.n179 10.6151
R1170 B.n183 B.n180 10.6151
R1171 B.n184 B.n183 10.6151
R1172 B.n187 B.n184 10.6151
R1173 B.n188 B.n187 10.6151
R1174 B.n191 B.n188 10.6151
R1175 B.n192 B.n191 10.6151
R1176 B.n195 B.n192 10.6151
R1177 B.n196 B.n195 10.6151
R1178 B.n199 B.n196 10.6151
R1179 B.n200 B.n199 10.6151
R1180 B.n203 B.n200 10.6151
R1181 B.n204 B.n203 10.6151
R1182 B.n207 B.n204 10.6151
R1183 B.n208 B.n207 10.6151
R1184 B.n211 B.n208 10.6151
R1185 B.n212 B.n211 10.6151
R1186 B.n215 B.n212 10.6151
R1187 B.n216 B.n215 10.6151
R1188 B.n219 B.n216 10.6151
R1189 B.n220 B.n219 10.6151
R1190 B.n223 B.n220 10.6151
R1191 B.n224 B.n223 10.6151
R1192 B.n227 B.n224 10.6151
R1193 B.n228 B.n227 10.6151
R1194 B.n231 B.n228 10.6151
R1195 B.n232 B.n231 10.6151
R1196 B.n236 B.n235 10.6151
R1197 B.n239 B.n236 10.6151
R1198 B.n240 B.n239 10.6151
R1199 B.n243 B.n240 10.6151
R1200 B.n244 B.n243 10.6151
R1201 B.n247 B.n244 10.6151
R1202 B.n248 B.n247 10.6151
R1203 B.n251 B.n248 10.6151
R1204 B.n252 B.n251 10.6151
R1205 B.n256 B.n255 10.6151
R1206 B.n259 B.n256 10.6151
R1207 B.n260 B.n259 10.6151
R1208 B.n263 B.n260 10.6151
R1209 B.n264 B.n263 10.6151
R1210 B.n267 B.n264 10.6151
R1211 B.n268 B.n267 10.6151
R1212 B.n271 B.n268 10.6151
R1213 B.n272 B.n271 10.6151
R1214 B.n275 B.n272 10.6151
R1215 B.n276 B.n275 10.6151
R1216 B.n279 B.n276 10.6151
R1217 B.n280 B.n279 10.6151
R1218 B.n283 B.n280 10.6151
R1219 B.n284 B.n283 10.6151
R1220 B.n287 B.n284 10.6151
R1221 B.n288 B.n287 10.6151
R1222 B.n291 B.n288 10.6151
R1223 B.n292 B.n291 10.6151
R1224 B.n295 B.n292 10.6151
R1225 B.n296 B.n295 10.6151
R1226 B.n299 B.n296 10.6151
R1227 B.n300 B.n299 10.6151
R1228 B.n303 B.n300 10.6151
R1229 B.n304 B.n303 10.6151
R1230 B.n307 B.n304 10.6151
R1231 B.n308 B.n307 10.6151
R1232 B.n311 B.n308 10.6151
R1233 B.n312 B.n311 10.6151
R1234 B.n315 B.n312 10.6151
R1235 B.n316 B.n315 10.6151
R1236 B.n319 B.n316 10.6151
R1237 B.n320 B.n319 10.6151
R1238 B.n323 B.n320 10.6151
R1239 B.n324 B.n323 10.6151
R1240 B.n327 B.n324 10.6151
R1241 B.n328 B.n327 10.6151
R1242 B.n331 B.n328 10.6151
R1243 B.n332 B.n331 10.6151
R1244 B.n335 B.n332 10.6151
R1245 B.n336 B.n335 10.6151
R1246 B.n339 B.n336 10.6151
R1247 B.n340 B.n339 10.6151
R1248 B.n343 B.n340 10.6151
R1249 B.n344 B.n343 10.6151
R1250 B.n347 B.n344 10.6151
R1251 B.n348 B.n347 10.6151
R1252 B.n351 B.n348 10.6151
R1253 B.n352 B.n351 10.6151
R1254 B.n355 B.n352 10.6151
R1255 B.n356 B.n355 10.6151
R1256 B.n359 B.n356 10.6151
R1257 B.n360 B.n359 10.6151
R1258 B.n363 B.n360 10.6151
R1259 B.n364 B.n363 10.6151
R1260 B.n367 B.n364 10.6151
R1261 B.n369 B.n367 10.6151
R1262 B.n370 B.n369 10.6151
R1263 B.n843 B.n370 10.6151
R1264 B.n751 B.n411 10.6151
R1265 B.n752 B.n751 10.6151
R1266 B.n753 B.n752 10.6151
R1267 B.n753 B.n403 10.6151
R1268 B.n763 B.n403 10.6151
R1269 B.n764 B.n763 10.6151
R1270 B.n765 B.n764 10.6151
R1271 B.n765 B.n395 10.6151
R1272 B.n775 B.n395 10.6151
R1273 B.n776 B.n775 10.6151
R1274 B.n777 B.n776 10.6151
R1275 B.n777 B.n387 10.6151
R1276 B.n787 B.n387 10.6151
R1277 B.n788 B.n787 10.6151
R1278 B.n789 B.n788 10.6151
R1279 B.n789 B.n379 10.6151
R1280 B.n799 B.n379 10.6151
R1281 B.n800 B.n799 10.6151
R1282 B.n802 B.n800 10.6151
R1283 B.n802 B.n801 10.6151
R1284 B.n801 B.n371 10.6151
R1285 B.n813 B.n371 10.6151
R1286 B.n814 B.n813 10.6151
R1287 B.n815 B.n814 10.6151
R1288 B.n816 B.n815 10.6151
R1289 B.n818 B.n816 10.6151
R1290 B.n819 B.n818 10.6151
R1291 B.n820 B.n819 10.6151
R1292 B.n821 B.n820 10.6151
R1293 B.n823 B.n821 10.6151
R1294 B.n824 B.n823 10.6151
R1295 B.n825 B.n824 10.6151
R1296 B.n826 B.n825 10.6151
R1297 B.n828 B.n826 10.6151
R1298 B.n829 B.n828 10.6151
R1299 B.n830 B.n829 10.6151
R1300 B.n831 B.n830 10.6151
R1301 B.n833 B.n831 10.6151
R1302 B.n834 B.n833 10.6151
R1303 B.n835 B.n834 10.6151
R1304 B.n836 B.n835 10.6151
R1305 B.n838 B.n836 10.6151
R1306 B.n839 B.n838 10.6151
R1307 B.n840 B.n839 10.6151
R1308 B.n841 B.n840 10.6151
R1309 B.n842 B.n841 10.6151
R1310 B.n745 B.n415 10.6151
R1311 B.n740 B.n415 10.6151
R1312 B.n740 B.n739 10.6151
R1313 B.n739 B.n738 10.6151
R1314 B.n738 B.n735 10.6151
R1315 B.n735 B.n734 10.6151
R1316 B.n734 B.n731 10.6151
R1317 B.n731 B.n730 10.6151
R1318 B.n730 B.n727 10.6151
R1319 B.n727 B.n726 10.6151
R1320 B.n726 B.n723 10.6151
R1321 B.n723 B.n722 10.6151
R1322 B.n722 B.n719 10.6151
R1323 B.n719 B.n718 10.6151
R1324 B.n718 B.n715 10.6151
R1325 B.n715 B.n714 10.6151
R1326 B.n714 B.n711 10.6151
R1327 B.n711 B.n710 10.6151
R1328 B.n710 B.n707 10.6151
R1329 B.n707 B.n706 10.6151
R1330 B.n706 B.n703 10.6151
R1331 B.n703 B.n702 10.6151
R1332 B.n702 B.n699 10.6151
R1333 B.n699 B.n698 10.6151
R1334 B.n698 B.n695 10.6151
R1335 B.n695 B.n694 10.6151
R1336 B.n694 B.n691 10.6151
R1337 B.n691 B.n690 10.6151
R1338 B.n690 B.n687 10.6151
R1339 B.n687 B.n686 10.6151
R1340 B.n686 B.n683 10.6151
R1341 B.n683 B.n682 10.6151
R1342 B.n682 B.n679 10.6151
R1343 B.n679 B.n678 10.6151
R1344 B.n678 B.n675 10.6151
R1345 B.n675 B.n674 10.6151
R1346 B.n674 B.n671 10.6151
R1347 B.n671 B.n670 10.6151
R1348 B.n670 B.n667 10.6151
R1349 B.n667 B.n666 10.6151
R1350 B.n666 B.n663 10.6151
R1351 B.n663 B.n662 10.6151
R1352 B.n662 B.n659 10.6151
R1353 B.n659 B.n658 10.6151
R1354 B.n658 B.n655 10.6151
R1355 B.n655 B.n654 10.6151
R1356 B.n654 B.n651 10.6151
R1357 B.n651 B.n650 10.6151
R1358 B.n650 B.n647 10.6151
R1359 B.n647 B.n646 10.6151
R1360 B.n646 B.n643 10.6151
R1361 B.n643 B.n642 10.6151
R1362 B.n642 B.n639 10.6151
R1363 B.n639 B.n638 10.6151
R1364 B.n638 B.n635 10.6151
R1365 B.n635 B.n634 10.6151
R1366 B.n634 B.n631 10.6151
R1367 B.n631 B.n630 10.6151
R1368 B.n630 B.n627 10.6151
R1369 B.n625 B.n622 10.6151
R1370 B.n622 B.n621 10.6151
R1371 B.n621 B.n618 10.6151
R1372 B.n618 B.n617 10.6151
R1373 B.n617 B.n614 10.6151
R1374 B.n614 B.n613 10.6151
R1375 B.n613 B.n610 10.6151
R1376 B.n610 B.n609 10.6151
R1377 B.n609 B.n606 10.6151
R1378 B.n604 B.n601 10.6151
R1379 B.n601 B.n600 10.6151
R1380 B.n600 B.n597 10.6151
R1381 B.n597 B.n596 10.6151
R1382 B.n596 B.n593 10.6151
R1383 B.n593 B.n592 10.6151
R1384 B.n592 B.n589 10.6151
R1385 B.n589 B.n588 10.6151
R1386 B.n588 B.n585 10.6151
R1387 B.n585 B.n584 10.6151
R1388 B.n584 B.n581 10.6151
R1389 B.n581 B.n580 10.6151
R1390 B.n580 B.n577 10.6151
R1391 B.n577 B.n576 10.6151
R1392 B.n576 B.n573 10.6151
R1393 B.n573 B.n572 10.6151
R1394 B.n572 B.n569 10.6151
R1395 B.n569 B.n568 10.6151
R1396 B.n568 B.n565 10.6151
R1397 B.n565 B.n564 10.6151
R1398 B.n564 B.n561 10.6151
R1399 B.n561 B.n560 10.6151
R1400 B.n560 B.n557 10.6151
R1401 B.n557 B.n556 10.6151
R1402 B.n556 B.n553 10.6151
R1403 B.n553 B.n552 10.6151
R1404 B.n552 B.n549 10.6151
R1405 B.n549 B.n548 10.6151
R1406 B.n548 B.n545 10.6151
R1407 B.n545 B.n544 10.6151
R1408 B.n544 B.n541 10.6151
R1409 B.n541 B.n540 10.6151
R1410 B.n540 B.n537 10.6151
R1411 B.n537 B.n536 10.6151
R1412 B.n536 B.n533 10.6151
R1413 B.n533 B.n532 10.6151
R1414 B.n532 B.n529 10.6151
R1415 B.n529 B.n528 10.6151
R1416 B.n528 B.n525 10.6151
R1417 B.n525 B.n524 10.6151
R1418 B.n524 B.n521 10.6151
R1419 B.n521 B.n520 10.6151
R1420 B.n520 B.n517 10.6151
R1421 B.n517 B.n516 10.6151
R1422 B.n516 B.n513 10.6151
R1423 B.n513 B.n512 10.6151
R1424 B.n512 B.n509 10.6151
R1425 B.n509 B.n508 10.6151
R1426 B.n508 B.n505 10.6151
R1427 B.n505 B.n504 10.6151
R1428 B.n504 B.n501 10.6151
R1429 B.n501 B.n500 10.6151
R1430 B.n500 B.n497 10.6151
R1431 B.n497 B.n496 10.6151
R1432 B.n496 B.n493 10.6151
R1433 B.n493 B.n492 10.6151
R1434 B.n492 B.n489 10.6151
R1435 B.n489 B.n488 10.6151
R1436 B.n488 B.n486 10.6151
R1437 B.n747 B.n746 10.6151
R1438 B.n747 B.n407 10.6151
R1439 B.n757 B.n407 10.6151
R1440 B.n758 B.n757 10.6151
R1441 B.n759 B.n758 10.6151
R1442 B.n759 B.n399 10.6151
R1443 B.n769 B.n399 10.6151
R1444 B.n770 B.n769 10.6151
R1445 B.n771 B.n770 10.6151
R1446 B.n771 B.n391 10.6151
R1447 B.n781 B.n391 10.6151
R1448 B.n782 B.n781 10.6151
R1449 B.n783 B.n782 10.6151
R1450 B.n783 B.n383 10.6151
R1451 B.n793 B.n383 10.6151
R1452 B.n794 B.n793 10.6151
R1453 B.n795 B.n794 10.6151
R1454 B.n795 B.n375 10.6151
R1455 B.n806 B.n375 10.6151
R1456 B.n807 B.n806 10.6151
R1457 B.n808 B.n807 10.6151
R1458 B.n808 B.n0 10.6151
R1459 B.n891 B.n1 10.6151
R1460 B.n891 B.n890 10.6151
R1461 B.n890 B.n889 10.6151
R1462 B.n889 B.n10 10.6151
R1463 B.n883 B.n10 10.6151
R1464 B.n883 B.n882 10.6151
R1465 B.n882 B.n881 10.6151
R1466 B.n881 B.n17 10.6151
R1467 B.n875 B.n17 10.6151
R1468 B.n875 B.n874 10.6151
R1469 B.n874 B.n873 10.6151
R1470 B.n873 B.n24 10.6151
R1471 B.n867 B.n24 10.6151
R1472 B.n867 B.n866 10.6151
R1473 B.n866 B.n865 10.6151
R1474 B.n865 B.n31 10.6151
R1475 B.n859 B.n31 10.6151
R1476 B.n859 B.n858 10.6151
R1477 B.n858 B.n857 10.6151
R1478 B.n857 B.n38 10.6151
R1479 B.n851 B.n38 10.6151
R1480 B.n851 B.n850 10.6151
R1481 B.n232 B.n117 9.36635
R1482 B.n255 B.n114 9.36635
R1483 B.n627 B.n626 9.36635
R1484 B.n605 B.n604 9.36635
R1485 B.t5 B.n381 7.92255
R1486 B.t4 B.n15 7.92255
R1487 B.n897 B.n0 2.81026
R1488 B.n897 B.n1 2.81026
R1489 B.n235 B.n117 1.24928
R1490 B.n252 B.n114 1.24928
R1491 B.n626 B.n625 1.24928
R1492 B.n606 B.n605 1.24928
R1493 B.n761 B.t14 0.466503
R1494 B.t3 B.n389 0.466503
R1495 B.t0 B.n22 0.466503
R1496 B.t7 B.n861 0.466503
R1497 VP.n5 VP.t0 525.255
R1498 VP.n12 VP.t1 506.608
R1499 VP.n19 VP.t4 506.608
R1500 VP.n9 VP.t5 506.608
R1501 VP.n1 VP.t2 465.003
R1502 VP.n4 VP.t3 465.003
R1503 VP.n20 VP.n19 161.3
R1504 VP.n7 VP.n6 161.3
R1505 VP.n8 VP.n3 161.3
R1506 VP.n10 VP.n9 161.3
R1507 VP.n18 VP.n0 161.3
R1508 VP.n17 VP.n16 161.3
R1509 VP.n15 VP.n14 161.3
R1510 VP.n13 VP.n2 161.3
R1511 VP.n12 VP.n11 161.3
R1512 VP.n14 VP.n13 51.1773
R1513 VP.n18 VP.n17 51.1773
R1514 VP.n8 VP.n7 51.1773
R1515 VP.n11 VP.n10 47.0384
R1516 VP.n6 VP.n5 43.2994
R1517 VP.n5 VP.n4 42.326
R1518 VP.n14 VP.n1 12.234
R1519 VP.n17 VP.n1 12.234
R1520 VP.n7 VP.n4 12.234
R1521 VP.n13 VP.n12 8.03383
R1522 VP.n19 VP.n18 8.03383
R1523 VP.n9 VP.n8 8.03383
R1524 VP.n6 VP.n3 0.189894
R1525 VP.n10 VP.n3 0.189894
R1526 VP.n11 VP.n2 0.189894
R1527 VP.n15 VP.n2 0.189894
R1528 VP.n16 VP.n15 0.189894
R1529 VP.n16 VP.n0 0.189894
R1530 VP.n20 VP.n0 0.189894
R1531 VP VP.n20 0.0516364
R1532 VTAIL.n410 VTAIL.n314 289.615
R1533 VTAIL.n98 VTAIL.n2 289.615
R1534 VTAIL.n308 VTAIL.n212 289.615
R1535 VTAIL.n204 VTAIL.n108 289.615
R1536 VTAIL.n346 VTAIL.n345 185
R1537 VTAIL.n351 VTAIL.n350 185
R1538 VTAIL.n353 VTAIL.n352 185
R1539 VTAIL.n342 VTAIL.n341 185
R1540 VTAIL.n359 VTAIL.n358 185
R1541 VTAIL.n361 VTAIL.n360 185
R1542 VTAIL.n338 VTAIL.n337 185
R1543 VTAIL.n367 VTAIL.n366 185
R1544 VTAIL.n369 VTAIL.n368 185
R1545 VTAIL.n334 VTAIL.n333 185
R1546 VTAIL.n375 VTAIL.n374 185
R1547 VTAIL.n377 VTAIL.n376 185
R1548 VTAIL.n330 VTAIL.n329 185
R1549 VTAIL.n383 VTAIL.n382 185
R1550 VTAIL.n385 VTAIL.n384 185
R1551 VTAIL.n326 VTAIL.n325 185
R1552 VTAIL.n392 VTAIL.n391 185
R1553 VTAIL.n393 VTAIL.n324 185
R1554 VTAIL.n395 VTAIL.n394 185
R1555 VTAIL.n322 VTAIL.n321 185
R1556 VTAIL.n401 VTAIL.n400 185
R1557 VTAIL.n403 VTAIL.n402 185
R1558 VTAIL.n318 VTAIL.n317 185
R1559 VTAIL.n409 VTAIL.n408 185
R1560 VTAIL.n411 VTAIL.n410 185
R1561 VTAIL.n34 VTAIL.n33 185
R1562 VTAIL.n39 VTAIL.n38 185
R1563 VTAIL.n41 VTAIL.n40 185
R1564 VTAIL.n30 VTAIL.n29 185
R1565 VTAIL.n47 VTAIL.n46 185
R1566 VTAIL.n49 VTAIL.n48 185
R1567 VTAIL.n26 VTAIL.n25 185
R1568 VTAIL.n55 VTAIL.n54 185
R1569 VTAIL.n57 VTAIL.n56 185
R1570 VTAIL.n22 VTAIL.n21 185
R1571 VTAIL.n63 VTAIL.n62 185
R1572 VTAIL.n65 VTAIL.n64 185
R1573 VTAIL.n18 VTAIL.n17 185
R1574 VTAIL.n71 VTAIL.n70 185
R1575 VTAIL.n73 VTAIL.n72 185
R1576 VTAIL.n14 VTAIL.n13 185
R1577 VTAIL.n80 VTAIL.n79 185
R1578 VTAIL.n81 VTAIL.n12 185
R1579 VTAIL.n83 VTAIL.n82 185
R1580 VTAIL.n10 VTAIL.n9 185
R1581 VTAIL.n89 VTAIL.n88 185
R1582 VTAIL.n91 VTAIL.n90 185
R1583 VTAIL.n6 VTAIL.n5 185
R1584 VTAIL.n97 VTAIL.n96 185
R1585 VTAIL.n99 VTAIL.n98 185
R1586 VTAIL.n309 VTAIL.n308 185
R1587 VTAIL.n307 VTAIL.n306 185
R1588 VTAIL.n216 VTAIL.n215 185
R1589 VTAIL.n301 VTAIL.n300 185
R1590 VTAIL.n299 VTAIL.n298 185
R1591 VTAIL.n220 VTAIL.n219 185
R1592 VTAIL.n293 VTAIL.n292 185
R1593 VTAIL.n291 VTAIL.n222 185
R1594 VTAIL.n290 VTAIL.n289 185
R1595 VTAIL.n225 VTAIL.n223 185
R1596 VTAIL.n284 VTAIL.n283 185
R1597 VTAIL.n282 VTAIL.n281 185
R1598 VTAIL.n229 VTAIL.n228 185
R1599 VTAIL.n276 VTAIL.n275 185
R1600 VTAIL.n274 VTAIL.n273 185
R1601 VTAIL.n233 VTAIL.n232 185
R1602 VTAIL.n268 VTAIL.n267 185
R1603 VTAIL.n266 VTAIL.n265 185
R1604 VTAIL.n237 VTAIL.n236 185
R1605 VTAIL.n260 VTAIL.n259 185
R1606 VTAIL.n258 VTAIL.n257 185
R1607 VTAIL.n241 VTAIL.n240 185
R1608 VTAIL.n252 VTAIL.n251 185
R1609 VTAIL.n250 VTAIL.n249 185
R1610 VTAIL.n245 VTAIL.n244 185
R1611 VTAIL.n205 VTAIL.n204 185
R1612 VTAIL.n203 VTAIL.n202 185
R1613 VTAIL.n112 VTAIL.n111 185
R1614 VTAIL.n197 VTAIL.n196 185
R1615 VTAIL.n195 VTAIL.n194 185
R1616 VTAIL.n116 VTAIL.n115 185
R1617 VTAIL.n189 VTAIL.n188 185
R1618 VTAIL.n187 VTAIL.n118 185
R1619 VTAIL.n186 VTAIL.n185 185
R1620 VTAIL.n121 VTAIL.n119 185
R1621 VTAIL.n180 VTAIL.n179 185
R1622 VTAIL.n178 VTAIL.n177 185
R1623 VTAIL.n125 VTAIL.n124 185
R1624 VTAIL.n172 VTAIL.n171 185
R1625 VTAIL.n170 VTAIL.n169 185
R1626 VTAIL.n129 VTAIL.n128 185
R1627 VTAIL.n164 VTAIL.n163 185
R1628 VTAIL.n162 VTAIL.n161 185
R1629 VTAIL.n133 VTAIL.n132 185
R1630 VTAIL.n156 VTAIL.n155 185
R1631 VTAIL.n154 VTAIL.n153 185
R1632 VTAIL.n137 VTAIL.n136 185
R1633 VTAIL.n148 VTAIL.n147 185
R1634 VTAIL.n146 VTAIL.n145 185
R1635 VTAIL.n141 VTAIL.n140 185
R1636 VTAIL.n347 VTAIL.t0 147.659
R1637 VTAIL.n35 VTAIL.t7 147.659
R1638 VTAIL.n246 VTAIL.t8 147.659
R1639 VTAIL.n142 VTAIL.t1 147.659
R1640 VTAIL.n351 VTAIL.n345 104.615
R1641 VTAIL.n352 VTAIL.n351 104.615
R1642 VTAIL.n352 VTAIL.n341 104.615
R1643 VTAIL.n359 VTAIL.n341 104.615
R1644 VTAIL.n360 VTAIL.n359 104.615
R1645 VTAIL.n360 VTAIL.n337 104.615
R1646 VTAIL.n367 VTAIL.n337 104.615
R1647 VTAIL.n368 VTAIL.n367 104.615
R1648 VTAIL.n368 VTAIL.n333 104.615
R1649 VTAIL.n375 VTAIL.n333 104.615
R1650 VTAIL.n376 VTAIL.n375 104.615
R1651 VTAIL.n376 VTAIL.n329 104.615
R1652 VTAIL.n383 VTAIL.n329 104.615
R1653 VTAIL.n384 VTAIL.n383 104.615
R1654 VTAIL.n384 VTAIL.n325 104.615
R1655 VTAIL.n392 VTAIL.n325 104.615
R1656 VTAIL.n393 VTAIL.n392 104.615
R1657 VTAIL.n394 VTAIL.n393 104.615
R1658 VTAIL.n394 VTAIL.n321 104.615
R1659 VTAIL.n401 VTAIL.n321 104.615
R1660 VTAIL.n402 VTAIL.n401 104.615
R1661 VTAIL.n402 VTAIL.n317 104.615
R1662 VTAIL.n409 VTAIL.n317 104.615
R1663 VTAIL.n410 VTAIL.n409 104.615
R1664 VTAIL.n39 VTAIL.n33 104.615
R1665 VTAIL.n40 VTAIL.n39 104.615
R1666 VTAIL.n40 VTAIL.n29 104.615
R1667 VTAIL.n47 VTAIL.n29 104.615
R1668 VTAIL.n48 VTAIL.n47 104.615
R1669 VTAIL.n48 VTAIL.n25 104.615
R1670 VTAIL.n55 VTAIL.n25 104.615
R1671 VTAIL.n56 VTAIL.n55 104.615
R1672 VTAIL.n56 VTAIL.n21 104.615
R1673 VTAIL.n63 VTAIL.n21 104.615
R1674 VTAIL.n64 VTAIL.n63 104.615
R1675 VTAIL.n64 VTAIL.n17 104.615
R1676 VTAIL.n71 VTAIL.n17 104.615
R1677 VTAIL.n72 VTAIL.n71 104.615
R1678 VTAIL.n72 VTAIL.n13 104.615
R1679 VTAIL.n80 VTAIL.n13 104.615
R1680 VTAIL.n81 VTAIL.n80 104.615
R1681 VTAIL.n82 VTAIL.n81 104.615
R1682 VTAIL.n82 VTAIL.n9 104.615
R1683 VTAIL.n89 VTAIL.n9 104.615
R1684 VTAIL.n90 VTAIL.n89 104.615
R1685 VTAIL.n90 VTAIL.n5 104.615
R1686 VTAIL.n97 VTAIL.n5 104.615
R1687 VTAIL.n98 VTAIL.n97 104.615
R1688 VTAIL.n308 VTAIL.n307 104.615
R1689 VTAIL.n307 VTAIL.n215 104.615
R1690 VTAIL.n300 VTAIL.n215 104.615
R1691 VTAIL.n300 VTAIL.n299 104.615
R1692 VTAIL.n299 VTAIL.n219 104.615
R1693 VTAIL.n292 VTAIL.n219 104.615
R1694 VTAIL.n292 VTAIL.n291 104.615
R1695 VTAIL.n291 VTAIL.n290 104.615
R1696 VTAIL.n290 VTAIL.n223 104.615
R1697 VTAIL.n283 VTAIL.n223 104.615
R1698 VTAIL.n283 VTAIL.n282 104.615
R1699 VTAIL.n282 VTAIL.n228 104.615
R1700 VTAIL.n275 VTAIL.n228 104.615
R1701 VTAIL.n275 VTAIL.n274 104.615
R1702 VTAIL.n274 VTAIL.n232 104.615
R1703 VTAIL.n267 VTAIL.n232 104.615
R1704 VTAIL.n267 VTAIL.n266 104.615
R1705 VTAIL.n266 VTAIL.n236 104.615
R1706 VTAIL.n259 VTAIL.n236 104.615
R1707 VTAIL.n259 VTAIL.n258 104.615
R1708 VTAIL.n258 VTAIL.n240 104.615
R1709 VTAIL.n251 VTAIL.n240 104.615
R1710 VTAIL.n251 VTAIL.n250 104.615
R1711 VTAIL.n250 VTAIL.n244 104.615
R1712 VTAIL.n204 VTAIL.n203 104.615
R1713 VTAIL.n203 VTAIL.n111 104.615
R1714 VTAIL.n196 VTAIL.n111 104.615
R1715 VTAIL.n196 VTAIL.n195 104.615
R1716 VTAIL.n195 VTAIL.n115 104.615
R1717 VTAIL.n188 VTAIL.n115 104.615
R1718 VTAIL.n188 VTAIL.n187 104.615
R1719 VTAIL.n187 VTAIL.n186 104.615
R1720 VTAIL.n186 VTAIL.n119 104.615
R1721 VTAIL.n179 VTAIL.n119 104.615
R1722 VTAIL.n179 VTAIL.n178 104.615
R1723 VTAIL.n178 VTAIL.n124 104.615
R1724 VTAIL.n171 VTAIL.n124 104.615
R1725 VTAIL.n171 VTAIL.n170 104.615
R1726 VTAIL.n170 VTAIL.n128 104.615
R1727 VTAIL.n163 VTAIL.n128 104.615
R1728 VTAIL.n163 VTAIL.n162 104.615
R1729 VTAIL.n162 VTAIL.n132 104.615
R1730 VTAIL.n155 VTAIL.n132 104.615
R1731 VTAIL.n155 VTAIL.n154 104.615
R1732 VTAIL.n154 VTAIL.n136 104.615
R1733 VTAIL.n147 VTAIL.n136 104.615
R1734 VTAIL.n147 VTAIL.n146 104.615
R1735 VTAIL.n146 VTAIL.n140 104.615
R1736 VTAIL.t0 VTAIL.n345 52.3082
R1737 VTAIL.t7 VTAIL.n33 52.3082
R1738 VTAIL.t8 VTAIL.n244 52.3082
R1739 VTAIL.t1 VTAIL.n140 52.3082
R1740 VTAIL.n211 VTAIL.n210 45.715
R1741 VTAIL.n107 VTAIL.n106 45.715
R1742 VTAIL.n1 VTAIL.n0 45.7148
R1743 VTAIL.n105 VTAIL.n104 45.7148
R1744 VTAIL.n415 VTAIL.n414 33.9308
R1745 VTAIL.n103 VTAIL.n102 33.9308
R1746 VTAIL.n313 VTAIL.n312 33.9308
R1747 VTAIL.n209 VTAIL.n208 33.9308
R1748 VTAIL.n107 VTAIL.n105 30.3755
R1749 VTAIL.n415 VTAIL.n313 29.2721
R1750 VTAIL.n347 VTAIL.n346 15.6677
R1751 VTAIL.n35 VTAIL.n34 15.6677
R1752 VTAIL.n246 VTAIL.n245 15.6677
R1753 VTAIL.n142 VTAIL.n141 15.6677
R1754 VTAIL.n395 VTAIL.n324 13.1884
R1755 VTAIL.n83 VTAIL.n12 13.1884
R1756 VTAIL.n293 VTAIL.n222 13.1884
R1757 VTAIL.n189 VTAIL.n118 13.1884
R1758 VTAIL.n350 VTAIL.n349 12.8005
R1759 VTAIL.n391 VTAIL.n390 12.8005
R1760 VTAIL.n396 VTAIL.n322 12.8005
R1761 VTAIL.n38 VTAIL.n37 12.8005
R1762 VTAIL.n79 VTAIL.n78 12.8005
R1763 VTAIL.n84 VTAIL.n10 12.8005
R1764 VTAIL.n294 VTAIL.n220 12.8005
R1765 VTAIL.n289 VTAIL.n224 12.8005
R1766 VTAIL.n249 VTAIL.n248 12.8005
R1767 VTAIL.n190 VTAIL.n116 12.8005
R1768 VTAIL.n185 VTAIL.n120 12.8005
R1769 VTAIL.n145 VTAIL.n144 12.8005
R1770 VTAIL.n353 VTAIL.n344 12.0247
R1771 VTAIL.n389 VTAIL.n326 12.0247
R1772 VTAIL.n400 VTAIL.n399 12.0247
R1773 VTAIL.n41 VTAIL.n32 12.0247
R1774 VTAIL.n77 VTAIL.n14 12.0247
R1775 VTAIL.n88 VTAIL.n87 12.0247
R1776 VTAIL.n298 VTAIL.n297 12.0247
R1777 VTAIL.n288 VTAIL.n225 12.0247
R1778 VTAIL.n252 VTAIL.n243 12.0247
R1779 VTAIL.n194 VTAIL.n193 12.0247
R1780 VTAIL.n184 VTAIL.n121 12.0247
R1781 VTAIL.n148 VTAIL.n139 12.0247
R1782 VTAIL.n354 VTAIL.n342 11.249
R1783 VTAIL.n386 VTAIL.n385 11.249
R1784 VTAIL.n403 VTAIL.n320 11.249
R1785 VTAIL.n42 VTAIL.n30 11.249
R1786 VTAIL.n74 VTAIL.n73 11.249
R1787 VTAIL.n91 VTAIL.n8 11.249
R1788 VTAIL.n301 VTAIL.n218 11.249
R1789 VTAIL.n285 VTAIL.n284 11.249
R1790 VTAIL.n253 VTAIL.n241 11.249
R1791 VTAIL.n197 VTAIL.n114 11.249
R1792 VTAIL.n181 VTAIL.n180 11.249
R1793 VTAIL.n149 VTAIL.n137 11.249
R1794 VTAIL.n358 VTAIL.n357 10.4732
R1795 VTAIL.n382 VTAIL.n328 10.4732
R1796 VTAIL.n404 VTAIL.n318 10.4732
R1797 VTAIL.n46 VTAIL.n45 10.4732
R1798 VTAIL.n70 VTAIL.n16 10.4732
R1799 VTAIL.n92 VTAIL.n6 10.4732
R1800 VTAIL.n302 VTAIL.n216 10.4732
R1801 VTAIL.n281 VTAIL.n227 10.4732
R1802 VTAIL.n257 VTAIL.n256 10.4732
R1803 VTAIL.n198 VTAIL.n112 10.4732
R1804 VTAIL.n177 VTAIL.n123 10.4732
R1805 VTAIL.n153 VTAIL.n152 10.4732
R1806 VTAIL.n361 VTAIL.n340 9.69747
R1807 VTAIL.n381 VTAIL.n330 9.69747
R1808 VTAIL.n408 VTAIL.n407 9.69747
R1809 VTAIL.n49 VTAIL.n28 9.69747
R1810 VTAIL.n69 VTAIL.n18 9.69747
R1811 VTAIL.n96 VTAIL.n95 9.69747
R1812 VTAIL.n306 VTAIL.n305 9.69747
R1813 VTAIL.n280 VTAIL.n229 9.69747
R1814 VTAIL.n260 VTAIL.n239 9.69747
R1815 VTAIL.n202 VTAIL.n201 9.69747
R1816 VTAIL.n176 VTAIL.n125 9.69747
R1817 VTAIL.n156 VTAIL.n135 9.69747
R1818 VTAIL.n414 VTAIL.n413 9.45567
R1819 VTAIL.n102 VTAIL.n101 9.45567
R1820 VTAIL.n312 VTAIL.n311 9.45567
R1821 VTAIL.n208 VTAIL.n207 9.45567
R1822 VTAIL.n413 VTAIL.n412 9.3005
R1823 VTAIL.n316 VTAIL.n315 9.3005
R1824 VTAIL.n407 VTAIL.n406 9.3005
R1825 VTAIL.n405 VTAIL.n404 9.3005
R1826 VTAIL.n320 VTAIL.n319 9.3005
R1827 VTAIL.n399 VTAIL.n398 9.3005
R1828 VTAIL.n397 VTAIL.n396 9.3005
R1829 VTAIL.n336 VTAIL.n335 9.3005
R1830 VTAIL.n365 VTAIL.n364 9.3005
R1831 VTAIL.n363 VTAIL.n362 9.3005
R1832 VTAIL.n340 VTAIL.n339 9.3005
R1833 VTAIL.n357 VTAIL.n356 9.3005
R1834 VTAIL.n355 VTAIL.n354 9.3005
R1835 VTAIL.n344 VTAIL.n343 9.3005
R1836 VTAIL.n349 VTAIL.n348 9.3005
R1837 VTAIL.n371 VTAIL.n370 9.3005
R1838 VTAIL.n373 VTAIL.n372 9.3005
R1839 VTAIL.n332 VTAIL.n331 9.3005
R1840 VTAIL.n379 VTAIL.n378 9.3005
R1841 VTAIL.n381 VTAIL.n380 9.3005
R1842 VTAIL.n328 VTAIL.n327 9.3005
R1843 VTAIL.n387 VTAIL.n386 9.3005
R1844 VTAIL.n389 VTAIL.n388 9.3005
R1845 VTAIL.n390 VTAIL.n323 9.3005
R1846 VTAIL.n101 VTAIL.n100 9.3005
R1847 VTAIL.n4 VTAIL.n3 9.3005
R1848 VTAIL.n95 VTAIL.n94 9.3005
R1849 VTAIL.n93 VTAIL.n92 9.3005
R1850 VTAIL.n8 VTAIL.n7 9.3005
R1851 VTAIL.n87 VTAIL.n86 9.3005
R1852 VTAIL.n85 VTAIL.n84 9.3005
R1853 VTAIL.n24 VTAIL.n23 9.3005
R1854 VTAIL.n53 VTAIL.n52 9.3005
R1855 VTAIL.n51 VTAIL.n50 9.3005
R1856 VTAIL.n28 VTAIL.n27 9.3005
R1857 VTAIL.n45 VTAIL.n44 9.3005
R1858 VTAIL.n43 VTAIL.n42 9.3005
R1859 VTAIL.n32 VTAIL.n31 9.3005
R1860 VTAIL.n37 VTAIL.n36 9.3005
R1861 VTAIL.n59 VTAIL.n58 9.3005
R1862 VTAIL.n61 VTAIL.n60 9.3005
R1863 VTAIL.n20 VTAIL.n19 9.3005
R1864 VTAIL.n67 VTAIL.n66 9.3005
R1865 VTAIL.n69 VTAIL.n68 9.3005
R1866 VTAIL.n16 VTAIL.n15 9.3005
R1867 VTAIL.n75 VTAIL.n74 9.3005
R1868 VTAIL.n77 VTAIL.n76 9.3005
R1869 VTAIL.n78 VTAIL.n11 9.3005
R1870 VTAIL.n272 VTAIL.n271 9.3005
R1871 VTAIL.n231 VTAIL.n230 9.3005
R1872 VTAIL.n278 VTAIL.n277 9.3005
R1873 VTAIL.n280 VTAIL.n279 9.3005
R1874 VTAIL.n227 VTAIL.n226 9.3005
R1875 VTAIL.n286 VTAIL.n285 9.3005
R1876 VTAIL.n288 VTAIL.n287 9.3005
R1877 VTAIL.n224 VTAIL.n221 9.3005
R1878 VTAIL.n311 VTAIL.n310 9.3005
R1879 VTAIL.n214 VTAIL.n213 9.3005
R1880 VTAIL.n305 VTAIL.n304 9.3005
R1881 VTAIL.n303 VTAIL.n302 9.3005
R1882 VTAIL.n218 VTAIL.n217 9.3005
R1883 VTAIL.n297 VTAIL.n296 9.3005
R1884 VTAIL.n295 VTAIL.n294 9.3005
R1885 VTAIL.n270 VTAIL.n269 9.3005
R1886 VTAIL.n235 VTAIL.n234 9.3005
R1887 VTAIL.n264 VTAIL.n263 9.3005
R1888 VTAIL.n262 VTAIL.n261 9.3005
R1889 VTAIL.n239 VTAIL.n238 9.3005
R1890 VTAIL.n256 VTAIL.n255 9.3005
R1891 VTAIL.n254 VTAIL.n253 9.3005
R1892 VTAIL.n243 VTAIL.n242 9.3005
R1893 VTAIL.n248 VTAIL.n247 9.3005
R1894 VTAIL.n168 VTAIL.n167 9.3005
R1895 VTAIL.n127 VTAIL.n126 9.3005
R1896 VTAIL.n174 VTAIL.n173 9.3005
R1897 VTAIL.n176 VTAIL.n175 9.3005
R1898 VTAIL.n123 VTAIL.n122 9.3005
R1899 VTAIL.n182 VTAIL.n181 9.3005
R1900 VTAIL.n184 VTAIL.n183 9.3005
R1901 VTAIL.n120 VTAIL.n117 9.3005
R1902 VTAIL.n207 VTAIL.n206 9.3005
R1903 VTAIL.n110 VTAIL.n109 9.3005
R1904 VTAIL.n201 VTAIL.n200 9.3005
R1905 VTAIL.n199 VTAIL.n198 9.3005
R1906 VTAIL.n114 VTAIL.n113 9.3005
R1907 VTAIL.n193 VTAIL.n192 9.3005
R1908 VTAIL.n191 VTAIL.n190 9.3005
R1909 VTAIL.n166 VTAIL.n165 9.3005
R1910 VTAIL.n131 VTAIL.n130 9.3005
R1911 VTAIL.n160 VTAIL.n159 9.3005
R1912 VTAIL.n158 VTAIL.n157 9.3005
R1913 VTAIL.n135 VTAIL.n134 9.3005
R1914 VTAIL.n152 VTAIL.n151 9.3005
R1915 VTAIL.n150 VTAIL.n149 9.3005
R1916 VTAIL.n139 VTAIL.n138 9.3005
R1917 VTAIL.n144 VTAIL.n143 9.3005
R1918 VTAIL.n362 VTAIL.n338 8.92171
R1919 VTAIL.n378 VTAIL.n377 8.92171
R1920 VTAIL.n411 VTAIL.n316 8.92171
R1921 VTAIL.n50 VTAIL.n26 8.92171
R1922 VTAIL.n66 VTAIL.n65 8.92171
R1923 VTAIL.n99 VTAIL.n4 8.92171
R1924 VTAIL.n309 VTAIL.n214 8.92171
R1925 VTAIL.n277 VTAIL.n276 8.92171
R1926 VTAIL.n261 VTAIL.n237 8.92171
R1927 VTAIL.n205 VTAIL.n110 8.92171
R1928 VTAIL.n173 VTAIL.n172 8.92171
R1929 VTAIL.n157 VTAIL.n133 8.92171
R1930 VTAIL.n366 VTAIL.n365 8.14595
R1931 VTAIL.n374 VTAIL.n332 8.14595
R1932 VTAIL.n412 VTAIL.n314 8.14595
R1933 VTAIL.n54 VTAIL.n53 8.14595
R1934 VTAIL.n62 VTAIL.n20 8.14595
R1935 VTAIL.n100 VTAIL.n2 8.14595
R1936 VTAIL.n310 VTAIL.n212 8.14595
R1937 VTAIL.n273 VTAIL.n231 8.14595
R1938 VTAIL.n265 VTAIL.n264 8.14595
R1939 VTAIL.n206 VTAIL.n108 8.14595
R1940 VTAIL.n169 VTAIL.n127 8.14595
R1941 VTAIL.n161 VTAIL.n160 8.14595
R1942 VTAIL.n369 VTAIL.n336 7.3702
R1943 VTAIL.n373 VTAIL.n334 7.3702
R1944 VTAIL.n57 VTAIL.n24 7.3702
R1945 VTAIL.n61 VTAIL.n22 7.3702
R1946 VTAIL.n272 VTAIL.n233 7.3702
R1947 VTAIL.n268 VTAIL.n235 7.3702
R1948 VTAIL.n168 VTAIL.n129 7.3702
R1949 VTAIL.n164 VTAIL.n131 7.3702
R1950 VTAIL.n370 VTAIL.n369 6.59444
R1951 VTAIL.n370 VTAIL.n334 6.59444
R1952 VTAIL.n58 VTAIL.n57 6.59444
R1953 VTAIL.n58 VTAIL.n22 6.59444
R1954 VTAIL.n269 VTAIL.n233 6.59444
R1955 VTAIL.n269 VTAIL.n268 6.59444
R1956 VTAIL.n165 VTAIL.n129 6.59444
R1957 VTAIL.n165 VTAIL.n164 6.59444
R1958 VTAIL.n366 VTAIL.n336 5.81868
R1959 VTAIL.n374 VTAIL.n373 5.81868
R1960 VTAIL.n414 VTAIL.n314 5.81868
R1961 VTAIL.n54 VTAIL.n24 5.81868
R1962 VTAIL.n62 VTAIL.n61 5.81868
R1963 VTAIL.n102 VTAIL.n2 5.81868
R1964 VTAIL.n312 VTAIL.n212 5.81868
R1965 VTAIL.n273 VTAIL.n272 5.81868
R1966 VTAIL.n265 VTAIL.n235 5.81868
R1967 VTAIL.n208 VTAIL.n108 5.81868
R1968 VTAIL.n169 VTAIL.n168 5.81868
R1969 VTAIL.n161 VTAIL.n131 5.81868
R1970 VTAIL.n365 VTAIL.n338 5.04292
R1971 VTAIL.n377 VTAIL.n332 5.04292
R1972 VTAIL.n412 VTAIL.n411 5.04292
R1973 VTAIL.n53 VTAIL.n26 5.04292
R1974 VTAIL.n65 VTAIL.n20 5.04292
R1975 VTAIL.n100 VTAIL.n99 5.04292
R1976 VTAIL.n310 VTAIL.n309 5.04292
R1977 VTAIL.n276 VTAIL.n231 5.04292
R1978 VTAIL.n264 VTAIL.n237 5.04292
R1979 VTAIL.n206 VTAIL.n205 5.04292
R1980 VTAIL.n172 VTAIL.n127 5.04292
R1981 VTAIL.n160 VTAIL.n133 5.04292
R1982 VTAIL.n348 VTAIL.n347 4.38563
R1983 VTAIL.n36 VTAIL.n35 4.38563
R1984 VTAIL.n247 VTAIL.n246 4.38563
R1985 VTAIL.n143 VTAIL.n142 4.38563
R1986 VTAIL.n362 VTAIL.n361 4.26717
R1987 VTAIL.n378 VTAIL.n330 4.26717
R1988 VTAIL.n408 VTAIL.n316 4.26717
R1989 VTAIL.n50 VTAIL.n49 4.26717
R1990 VTAIL.n66 VTAIL.n18 4.26717
R1991 VTAIL.n96 VTAIL.n4 4.26717
R1992 VTAIL.n306 VTAIL.n214 4.26717
R1993 VTAIL.n277 VTAIL.n229 4.26717
R1994 VTAIL.n261 VTAIL.n260 4.26717
R1995 VTAIL.n202 VTAIL.n110 4.26717
R1996 VTAIL.n173 VTAIL.n125 4.26717
R1997 VTAIL.n157 VTAIL.n156 4.26717
R1998 VTAIL.n358 VTAIL.n340 3.49141
R1999 VTAIL.n382 VTAIL.n381 3.49141
R2000 VTAIL.n407 VTAIL.n318 3.49141
R2001 VTAIL.n46 VTAIL.n28 3.49141
R2002 VTAIL.n70 VTAIL.n69 3.49141
R2003 VTAIL.n95 VTAIL.n6 3.49141
R2004 VTAIL.n305 VTAIL.n216 3.49141
R2005 VTAIL.n281 VTAIL.n280 3.49141
R2006 VTAIL.n257 VTAIL.n239 3.49141
R2007 VTAIL.n201 VTAIL.n112 3.49141
R2008 VTAIL.n177 VTAIL.n176 3.49141
R2009 VTAIL.n153 VTAIL.n135 3.49141
R2010 VTAIL.n357 VTAIL.n342 2.71565
R2011 VTAIL.n385 VTAIL.n328 2.71565
R2012 VTAIL.n404 VTAIL.n403 2.71565
R2013 VTAIL.n45 VTAIL.n30 2.71565
R2014 VTAIL.n73 VTAIL.n16 2.71565
R2015 VTAIL.n92 VTAIL.n91 2.71565
R2016 VTAIL.n302 VTAIL.n301 2.71565
R2017 VTAIL.n284 VTAIL.n227 2.71565
R2018 VTAIL.n256 VTAIL.n241 2.71565
R2019 VTAIL.n198 VTAIL.n197 2.71565
R2020 VTAIL.n180 VTAIL.n123 2.71565
R2021 VTAIL.n152 VTAIL.n137 2.71565
R2022 VTAIL.n354 VTAIL.n353 1.93989
R2023 VTAIL.n386 VTAIL.n326 1.93989
R2024 VTAIL.n400 VTAIL.n320 1.93989
R2025 VTAIL.n42 VTAIL.n41 1.93989
R2026 VTAIL.n74 VTAIL.n14 1.93989
R2027 VTAIL.n88 VTAIL.n8 1.93989
R2028 VTAIL.n298 VTAIL.n218 1.93989
R2029 VTAIL.n285 VTAIL.n225 1.93989
R2030 VTAIL.n253 VTAIL.n252 1.93989
R2031 VTAIL.n194 VTAIL.n114 1.93989
R2032 VTAIL.n181 VTAIL.n121 1.93989
R2033 VTAIL.n149 VTAIL.n148 1.93989
R2034 VTAIL.n350 VTAIL.n344 1.16414
R2035 VTAIL.n391 VTAIL.n389 1.16414
R2036 VTAIL.n399 VTAIL.n322 1.16414
R2037 VTAIL.n38 VTAIL.n32 1.16414
R2038 VTAIL.n79 VTAIL.n77 1.16414
R2039 VTAIL.n87 VTAIL.n10 1.16414
R2040 VTAIL.n297 VTAIL.n220 1.16414
R2041 VTAIL.n289 VTAIL.n288 1.16414
R2042 VTAIL.n249 VTAIL.n243 1.16414
R2043 VTAIL.n193 VTAIL.n116 1.16414
R2044 VTAIL.n185 VTAIL.n184 1.16414
R2045 VTAIL.n145 VTAIL.n139 1.16414
R2046 VTAIL.n209 VTAIL.n107 1.10395
R2047 VTAIL.n313 VTAIL.n211 1.10395
R2048 VTAIL.n105 VTAIL.n103 1.10395
R2049 VTAIL.n0 VTAIL.t2 1.0807
R2050 VTAIL.n0 VTAIL.t4 1.0807
R2051 VTAIL.n104 VTAIL.t6 1.0807
R2052 VTAIL.n104 VTAIL.t5 1.0807
R2053 VTAIL.n210 VTAIL.t9 1.0807
R2054 VTAIL.n210 VTAIL.t10 1.0807
R2055 VTAIL.n106 VTAIL.t11 1.0807
R2056 VTAIL.n106 VTAIL.t3 1.0807
R2057 VTAIL.n211 VTAIL.n209 1.02205
R2058 VTAIL.n103 VTAIL.n1 1.02205
R2059 VTAIL VTAIL.n415 0.769897
R2060 VTAIL.n349 VTAIL.n346 0.388379
R2061 VTAIL.n390 VTAIL.n324 0.388379
R2062 VTAIL.n396 VTAIL.n395 0.388379
R2063 VTAIL.n37 VTAIL.n34 0.388379
R2064 VTAIL.n78 VTAIL.n12 0.388379
R2065 VTAIL.n84 VTAIL.n83 0.388379
R2066 VTAIL.n294 VTAIL.n293 0.388379
R2067 VTAIL.n224 VTAIL.n222 0.388379
R2068 VTAIL.n248 VTAIL.n245 0.388379
R2069 VTAIL.n190 VTAIL.n189 0.388379
R2070 VTAIL.n120 VTAIL.n118 0.388379
R2071 VTAIL.n144 VTAIL.n141 0.388379
R2072 VTAIL VTAIL.n1 0.334552
R2073 VTAIL.n348 VTAIL.n343 0.155672
R2074 VTAIL.n355 VTAIL.n343 0.155672
R2075 VTAIL.n356 VTAIL.n355 0.155672
R2076 VTAIL.n356 VTAIL.n339 0.155672
R2077 VTAIL.n363 VTAIL.n339 0.155672
R2078 VTAIL.n364 VTAIL.n363 0.155672
R2079 VTAIL.n364 VTAIL.n335 0.155672
R2080 VTAIL.n371 VTAIL.n335 0.155672
R2081 VTAIL.n372 VTAIL.n371 0.155672
R2082 VTAIL.n372 VTAIL.n331 0.155672
R2083 VTAIL.n379 VTAIL.n331 0.155672
R2084 VTAIL.n380 VTAIL.n379 0.155672
R2085 VTAIL.n380 VTAIL.n327 0.155672
R2086 VTAIL.n387 VTAIL.n327 0.155672
R2087 VTAIL.n388 VTAIL.n387 0.155672
R2088 VTAIL.n388 VTAIL.n323 0.155672
R2089 VTAIL.n397 VTAIL.n323 0.155672
R2090 VTAIL.n398 VTAIL.n397 0.155672
R2091 VTAIL.n398 VTAIL.n319 0.155672
R2092 VTAIL.n405 VTAIL.n319 0.155672
R2093 VTAIL.n406 VTAIL.n405 0.155672
R2094 VTAIL.n406 VTAIL.n315 0.155672
R2095 VTAIL.n413 VTAIL.n315 0.155672
R2096 VTAIL.n36 VTAIL.n31 0.155672
R2097 VTAIL.n43 VTAIL.n31 0.155672
R2098 VTAIL.n44 VTAIL.n43 0.155672
R2099 VTAIL.n44 VTAIL.n27 0.155672
R2100 VTAIL.n51 VTAIL.n27 0.155672
R2101 VTAIL.n52 VTAIL.n51 0.155672
R2102 VTAIL.n52 VTAIL.n23 0.155672
R2103 VTAIL.n59 VTAIL.n23 0.155672
R2104 VTAIL.n60 VTAIL.n59 0.155672
R2105 VTAIL.n60 VTAIL.n19 0.155672
R2106 VTAIL.n67 VTAIL.n19 0.155672
R2107 VTAIL.n68 VTAIL.n67 0.155672
R2108 VTAIL.n68 VTAIL.n15 0.155672
R2109 VTAIL.n75 VTAIL.n15 0.155672
R2110 VTAIL.n76 VTAIL.n75 0.155672
R2111 VTAIL.n76 VTAIL.n11 0.155672
R2112 VTAIL.n85 VTAIL.n11 0.155672
R2113 VTAIL.n86 VTAIL.n85 0.155672
R2114 VTAIL.n86 VTAIL.n7 0.155672
R2115 VTAIL.n93 VTAIL.n7 0.155672
R2116 VTAIL.n94 VTAIL.n93 0.155672
R2117 VTAIL.n94 VTAIL.n3 0.155672
R2118 VTAIL.n101 VTAIL.n3 0.155672
R2119 VTAIL.n311 VTAIL.n213 0.155672
R2120 VTAIL.n304 VTAIL.n213 0.155672
R2121 VTAIL.n304 VTAIL.n303 0.155672
R2122 VTAIL.n303 VTAIL.n217 0.155672
R2123 VTAIL.n296 VTAIL.n217 0.155672
R2124 VTAIL.n296 VTAIL.n295 0.155672
R2125 VTAIL.n295 VTAIL.n221 0.155672
R2126 VTAIL.n287 VTAIL.n221 0.155672
R2127 VTAIL.n287 VTAIL.n286 0.155672
R2128 VTAIL.n286 VTAIL.n226 0.155672
R2129 VTAIL.n279 VTAIL.n226 0.155672
R2130 VTAIL.n279 VTAIL.n278 0.155672
R2131 VTAIL.n278 VTAIL.n230 0.155672
R2132 VTAIL.n271 VTAIL.n230 0.155672
R2133 VTAIL.n271 VTAIL.n270 0.155672
R2134 VTAIL.n270 VTAIL.n234 0.155672
R2135 VTAIL.n263 VTAIL.n234 0.155672
R2136 VTAIL.n263 VTAIL.n262 0.155672
R2137 VTAIL.n262 VTAIL.n238 0.155672
R2138 VTAIL.n255 VTAIL.n238 0.155672
R2139 VTAIL.n255 VTAIL.n254 0.155672
R2140 VTAIL.n254 VTAIL.n242 0.155672
R2141 VTAIL.n247 VTAIL.n242 0.155672
R2142 VTAIL.n207 VTAIL.n109 0.155672
R2143 VTAIL.n200 VTAIL.n109 0.155672
R2144 VTAIL.n200 VTAIL.n199 0.155672
R2145 VTAIL.n199 VTAIL.n113 0.155672
R2146 VTAIL.n192 VTAIL.n113 0.155672
R2147 VTAIL.n192 VTAIL.n191 0.155672
R2148 VTAIL.n191 VTAIL.n117 0.155672
R2149 VTAIL.n183 VTAIL.n117 0.155672
R2150 VTAIL.n183 VTAIL.n182 0.155672
R2151 VTAIL.n182 VTAIL.n122 0.155672
R2152 VTAIL.n175 VTAIL.n122 0.155672
R2153 VTAIL.n175 VTAIL.n174 0.155672
R2154 VTAIL.n174 VTAIL.n126 0.155672
R2155 VTAIL.n167 VTAIL.n126 0.155672
R2156 VTAIL.n167 VTAIL.n166 0.155672
R2157 VTAIL.n166 VTAIL.n130 0.155672
R2158 VTAIL.n159 VTAIL.n130 0.155672
R2159 VTAIL.n159 VTAIL.n158 0.155672
R2160 VTAIL.n158 VTAIL.n134 0.155672
R2161 VTAIL.n151 VTAIL.n134 0.155672
R2162 VTAIL.n151 VTAIL.n150 0.155672
R2163 VTAIL.n150 VTAIL.n138 0.155672
R2164 VTAIL.n143 VTAIL.n138 0.155672
R2165 VDD1.n96 VDD1.n0 289.615
R2166 VDD1.n197 VDD1.n101 289.615
R2167 VDD1.n97 VDD1.n96 185
R2168 VDD1.n95 VDD1.n94 185
R2169 VDD1.n4 VDD1.n3 185
R2170 VDD1.n89 VDD1.n88 185
R2171 VDD1.n87 VDD1.n86 185
R2172 VDD1.n8 VDD1.n7 185
R2173 VDD1.n81 VDD1.n80 185
R2174 VDD1.n79 VDD1.n10 185
R2175 VDD1.n78 VDD1.n77 185
R2176 VDD1.n13 VDD1.n11 185
R2177 VDD1.n72 VDD1.n71 185
R2178 VDD1.n70 VDD1.n69 185
R2179 VDD1.n17 VDD1.n16 185
R2180 VDD1.n64 VDD1.n63 185
R2181 VDD1.n62 VDD1.n61 185
R2182 VDD1.n21 VDD1.n20 185
R2183 VDD1.n56 VDD1.n55 185
R2184 VDD1.n54 VDD1.n53 185
R2185 VDD1.n25 VDD1.n24 185
R2186 VDD1.n48 VDD1.n47 185
R2187 VDD1.n46 VDD1.n45 185
R2188 VDD1.n29 VDD1.n28 185
R2189 VDD1.n40 VDD1.n39 185
R2190 VDD1.n38 VDD1.n37 185
R2191 VDD1.n33 VDD1.n32 185
R2192 VDD1.n133 VDD1.n132 185
R2193 VDD1.n138 VDD1.n137 185
R2194 VDD1.n140 VDD1.n139 185
R2195 VDD1.n129 VDD1.n128 185
R2196 VDD1.n146 VDD1.n145 185
R2197 VDD1.n148 VDD1.n147 185
R2198 VDD1.n125 VDD1.n124 185
R2199 VDD1.n154 VDD1.n153 185
R2200 VDD1.n156 VDD1.n155 185
R2201 VDD1.n121 VDD1.n120 185
R2202 VDD1.n162 VDD1.n161 185
R2203 VDD1.n164 VDD1.n163 185
R2204 VDD1.n117 VDD1.n116 185
R2205 VDD1.n170 VDD1.n169 185
R2206 VDD1.n172 VDD1.n171 185
R2207 VDD1.n113 VDD1.n112 185
R2208 VDD1.n179 VDD1.n178 185
R2209 VDD1.n180 VDD1.n111 185
R2210 VDD1.n182 VDD1.n181 185
R2211 VDD1.n109 VDD1.n108 185
R2212 VDD1.n188 VDD1.n187 185
R2213 VDD1.n190 VDD1.n189 185
R2214 VDD1.n105 VDD1.n104 185
R2215 VDD1.n196 VDD1.n195 185
R2216 VDD1.n198 VDD1.n197 185
R2217 VDD1.n34 VDD1.t5 147.659
R2218 VDD1.n134 VDD1.t4 147.659
R2219 VDD1.n96 VDD1.n95 104.615
R2220 VDD1.n95 VDD1.n3 104.615
R2221 VDD1.n88 VDD1.n3 104.615
R2222 VDD1.n88 VDD1.n87 104.615
R2223 VDD1.n87 VDD1.n7 104.615
R2224 VDD1.n80 VDD1.n7 104.615
R2225 VDD1.n80 VDD1.n79 104.615
R2226 VDD1.n79 VDD1.n78 104.615
R2227 VDD1.n78 VDD1.n11 104.615
R2228 VDD1.n71 VDD1.n11 104.615
R2229 VDD1.n71 VDD1.n70 104.615
R2230 VDD1.n70 VDD1.n16 104.615
R2231 VDD1.n63 VDD1.n16 104.615
R2232 VDD1.n63 VDD1.n62 104.615
R2233 VDD1.n62 VDD1.n20 104.615
R2234 VDD1.n55 VDD1.n20 104.615
R2235 VDD1.n55 VDD1.n54 104.615
R2236 VDD1.n54 VDD1.n24 104.615
R2237 VDD1.n47 VDD1.n24 104.615
R2238 VDD1.n47 VDD1.n46 104.615
R2239 VDD1.n46 VDD1.n28 104.615
R2240 VDD1.n39 VDD1.n28 104.615
R2241 VDD1.n39 VDD1.n38 104.615
R2242 VDD1.n38 VDD1.n32 104.615
R2243 VDD1.n138 VDD1.n132 104.615
R2244 VDD1.n139 VDD1.n138 104.615
R2245 VDD1.n139 VDD1.n128 104.615
R2246 VDD1.n146 VDD1.n128 104.615
R2247 VDD1.n147 VDD1.n146 104.615
R2248 VDD1.n147 VDD1.n124 104.615
R2249 VDD1.n154 VDD1.n124 104.615
R2250 VDD1.n155 VDD1.n154 104.615
R2251 VDD1.n155 VDD1.n120 104.615
R2252 VDD1.n162 VDD1.n120 104.615
R2253 VDD1.n163 VDD1.n162 104.615
R2254 VDD1.n163 VDD1.n116 104.615
R2255 VDD1.n170 VDD1.n116 104.615
R2256 VDD1.n171 VDD1.n170 104.615
R2257 VDD1.n171 VDD1.n112 104.615
R2258 VDD1.n179 VDD1.n112 104.615
R2259 VDD1.n180 VDD1.n179 104.615
R2260 VDD1.n181 VDD1.n180 104.615
R2261 VDD1.n181 VDD1.n108 104.615
R2262 VDD1.n188 VDD1.n108 104.615
R2263 VDD1.n189 VDD1.n188 104.615
R2264 VDD1.n189 VDD1.n104 104.615
R2265 VDD1.n196 VDD1.n104 104.615
R2266 VDD1.n197 VDD1.n196 104.615
R2267 VDD1.n203 VDD1.n202 62.6141
R2268 VDD1.n205 VDD1.n204 62.3936
R2269 VDD1.t5 VDD1.n32 52.3082
R2270 VDD1.t4 VDD1.n132 52.3082
R2271 VDD1 VDD1.n100 51.4954
R2272 VDD1.n203 VDD1.n201 51.3818
R2273 VDD1.n205 VDD1.n203 44.238
R2274 VDD1.n34 VDD1.n33 15.6677
R2275 VDD1.n134 VDD1.n133 15.6677
R2276 VDD1.n81 VDD1.n10 13.1884
R2277 VDD1.n182 VDD1.n111 13.1884
R2278 VDD1.n82 VDD1.n8 12.8005
R2279 VDD1.n77 VDD1.n12 12.8005
R2280 VDD1.n37 VDD1.n36 12.8005
R2281 VDD1.n137 VDD1.n136 12.8005
R2282 VDD1.n178 VDD1.n177 12.8005
R2283 VDD1.n183 VDD1.n109 12.8005
R2284 VDD1.n86 VDD1.n85 12.0247
R2285 VDD1.n76 VDD1.n13 12.0247
R2286 VDD1.n40 VDD1.n31 12.0247
R2287 VDD1.n140 VDD1.n131 12.0247
R2288 VDD1.n176 VDD1.n113 12.0247
R2289 VDD1.n187 VDD1.n186 12.0247
R2290 VDD1.n89 VDD1.n6 11.249
R2291 VDD1.n73 VDD1.n72 11.249
R2292 VDD1.n41 VDD1.n29 11.249
R2293 VDD1.n141 VDD1.n129 11.249
R2294 VDD1.n173 VDD1.n172 11.249
R2295 VDD1.n190 VDD1.n107 11.249
R2296 VDD1.n90 VDD1.n4 10.4732
R2297 VDD1.n69 VDD1.n15 10.4732
R2298 VDD1.n45 VDD1.n44 10.4732
R2299 VDD1.n145 VDD1.n144 10.4732
R2300 VDD1.n169 VDD1.n115 10.4732
R2301 VDD1.n191 VDD1.n105 10.4732
R2302 VDD1.n94 VDD1.n93 9.69747
R2303 VDD1.n68 VDD1.n17 9.69747
R2304 VDD1.n48 VDD1.n27 9.69747
R2305 VDD1.n148 VDD1.n127 9.69747
R2306 VDD1.n168 VDD1.n117 9.69747
R2307 VDD1.n195 VDD1.n194 9.69747
R2308 VDD1.n100 VDD1.n99 9.45567
R2309 VDD1.n201 VDD1.n200 9.45567
R2310 VDD1.n60 VDD1.n59 9.3005
R2311 VDD1.n19 VDD1.n18 9.3005
R2312 VDD1.n66 VDD1.n65 9.3005
R2313 VDD1.n68 VDD1.n67 9.3005
R2314 VDD1.n15 VDD1.n14 9.3005
R2315 VDD1.n74 VDD1.n73 9.3005
R2316 VDD1.n76 VDD1.n75 9.3005
R2317 VDD1.n12 VDD1.n9 9.3005
R2318 VDD1.n99 VDD1.n98 9.3005
R2319 VDD1.n2 VDD1.n1 9.3005
R2320 VDD1.n93 VDD1.n92 9.3005
R2321 VDD1.n91 VDD1.n90 9.3005
R2322 VDD1.n6 VDD1.n5 9.3005
R2323 VDD1.n85 VDD1.n84 9.3005
R2324 VDD1.n83 VDD1.n82 9.3005
R2325 VDD1.n58 VDD1.n57 9.3005
R2326 VDD1.n23 VDD1.n22 9.3005
R2327 VDD1.n52 VDD1.n51 9.3005
R2328 VDD1.n50 VDD1.n49 9.3005
R2329 VDD1.n27 VDD1.n26 9.3005
R2330 VDD1.n44 VDD1.n43 9.3005
R2331 VDD1.n42 VDD1.n41 9.3005
R2332 VDD1.n31 VDD1.n30 9.3005
R2333 VDD1.n36 VDD1.n35 9.3005
R2334 VDD1.n200 VDD1.n199 9.3005
R2335 VDD1.n103 VDD1.n102 9.3005
R2336 VDD1.n194 VDD1.n193 9.3005
R2337 VDD1.n192 VDD1.n191 9.3005
R2338 VDD1.n107 VDD1.n106 9.3005
R2339 VDD1.n186 VDD1.n185 9.3005
R2340 VDD1.n184 VDD1.n183 9.3005
R2341 VDD1.n123 VDD1.n122 9.3005
R2342 VDD1.n152 VDD1.n151 9.3005
R2343 VDD1.n150 VDD1.n149 9.3005
R2344 VDD1.n127 VDD1.n126 9.3005
R2345 VDD1.n144 VDD1.n143 9.3005
R2346 VDD1.n142 VDD1.n141 9.3005
R2347 VDD1.n131 VDD1.n130 9.3005
R2348 VDD1.n136 VDD1.n135 9.3005
R2349 VDD1.n158 VDD1.n157 9.3005
R2350 VDD1.n160 VDD1.n159 9.3005
R2351 VDD1.n119 VDD1.n118 9.3005
R2352 VDD1.n166 VDD1.n165 9.3005
R2353 VDD1.n168 VDD1.n167 9.3005
R2354 VDD1.n115 VDD1.n114 9.3005
R2355 VDD1.n174 VDD1.n173 9.3005
R2356 VDD1.n176 VDD1.n175 9.3005
R2357 VDD1.n177 VDD1.n110 9.3005
R2358 VDD1.n97 VDD1.n2 8.92171
R2359 VDD1.n65 VDD1.n64 8.92171
R2360 VDD1.n49 VDD1.n25 8.92171
R2361 VDD1.n149 VDD1.n125 8.92171
R2362 VDD1.n165 VDD1.n164 8.92171
R2363 VDD1.n198 VDD1.n103 8.92171
R2364 VDD1.n98 VDD1.n0 8.14595
R2365 VDD1.n61 VDD1.n19 8.14595
R2366 VDD1.n53 VDD1.n52 8.14595
R2367 VDD1.n153 VDD1.n152 8.14595
R2368 VDD1.n161 VDD1.n119 8.14595
R2369 VDD1.n199 VDD1.n101 8.14595
R2370 VDD1.n60 VDD1.n21 7.3702
R2371 VDD1.n56 VDD1.n23 7.3702
R2372 VDD1.n156 VDD1.n123 7.3702
R2373 VDD1.n160 VDD1.n121 7.3702
R2374 VDD1.n57 VDD1.n21 6.59444
R2375 VDD1.n57 VDD1.n56 6.59444
R2376 VDD1.n157 VDD1.n156 6.59444
R2377 VDD1.n157 VDD1.n121 6.59444
R2378 VDD1.n100 VDD1.n0 5.81868
R2379 VDD1.n61 VDD1.n60 5.81868
R2380 VDD1.n53 VDD1.n23 5.81868
R2381 VDD1.n153 VDD1.n123 5.81868
R2382 VDD1.n161 VDD1.n160 5.81868
R2383 VDD1.n201 VDD1.n101 5.81868
R2384 VDD1.n98 VDD1.n97 5.04292
R2385 VDD1.n64 VDD1.n19 5.04292
R2386 VDD1.n52 VDD1.n25 5.04292
R2387 VDD1.n152 VDD1.n125 5.04292
R2388 VDD1.n164 VDD1.n119 5.04292
R2389 VDD1.n199 VDD1.n198 5.04292
R2390 VDD1.n35 VDD1.n34 4.38563
R2391 VDD1.n135 VDD1.n134 4.38563
R2392 VDD1.n94 VDD1.n2 4.26717
R2393 VDD1.n65 VDD1.n17 4.26717
R2394 VDD1.n49 VDD1.n48 4.26717
R2395 VDD1.n149 VDD1.n148 4.26717
R2396 VDD1.n165 VDD1.n117 4.26717
R2397 VDD1.n195 VDD1.n103 4.26717
R2398 VDD1.n93 VDD1.n4 3.49141
R2399 VDD1.n69 VDD1.n68 3.49141
R2400 VDD1.n45 VDD1.n27 3.49141
R2401 VDD1.n145 VDD1.n127 3.49141
R2402 VDD1.n169 VDD1.n168 3.49141
R2403 VDD1.n194 VDD1.n105 3.49141
R2404 VDD1.n90 VDD1.n89 2.71565
R2405 VDD1.n72 VDD1.n15 2.71565
R2406 VDD1.n44 VDD1.n29 2.71565
R2407 VDD1.n144 VDD1.n129 2.71565
R2408 VDD1.n172 VDD1.n115 2.71565
R2409 VDD1.n191 VDD1.n190 2.71565
R2410 VDD1.n86 VDD1.n6 1.93989
R2411 VDD1.n73 VDD1.n13 1.93989
R2412 VDD1.n41 VDD1.n40 1.93989
R2413 VDD1.n141 VDD1.n140 1.93989
R2414 VDD1.n173 VDD1.n113 1.93989
R2415 VDD1.n187 VDD1.n107 1.93989
R2416 VDD1.n85 VDD1.n8 1.16414
R2417 VDD1.n77 VDD1.n76 1.16414
R2418 VDD1.n37 VDD1.n31 1.16414
R2419 VDD1.n137 VDD1.n131 1.16414
R2420 VDD1.n178 VDD1.n176 1.16414
R2421 VDD1.n186 VDD1.n109 1.16414
R2422 VDD1.n204 VDD1.t2 1.0807
R2423 VDD1.n204 VDD1.t0 1.0807
R2424 VDD1.n202 VDD1.t3 1.0807
R2425 VDD1.n202 VDD1.t1 1.0807
R2426 VDD1.n82 VDD1.n81 0.388379
R2427 VDD1.n12 VDD1.n10 0.388379
R2428 VDD1.n36 VDD1.n33 0.388379
R2429 VDD1.n136 VDD1.n133 0.388379
R2430 VDD1.n177 VDD1.n111 0.388379
R2431 VDD1.n183 VDD1.n182 0.388379
R2432 VDD1 VDD1.n205 0.218172
R2433 VDD1.n99 VDD1.n1 0.155672
R2434 VDD1.n92 VDD1.n1 0.155672
R2435 VDD1.n92 VDD1.n91 0.155672
R2436 VDD1.n91 VDD1.n5 0.155672
R2437 VDD1.n84 VDD1.n5 0.155672
R2438 VDD1.n84 VDD1.n83 0.155672
R2439 VDD1.n83 VDD1.n9 0.155672
R2440 VDD1.n75 VDD1.n9 0.155672
R2441 VDD1.n75 VDD1.n74 0.155672
R2442 VDD1.n74 VDD1.n14 0.155672
R2443 VDD1.n67 VDD1.n14 0.155672
R2444 VDD1.n67 VDD1.n66 0.155672
R2445 VDD1.n66 VDD1.n18 0.155672
R2446 VDD1.n59 VDD1.n18 0.155672
R2447 VDD1.n59 VDD1.n58 0.155672
R2448 VDD1.n58 VDD1.n22 0.155672
R2449 VDD1.n51 VDD1.n22 0.155672
R2450 VDD1.n51 VDD1.n50 0.155672
R2451 VDD1.n50 VDD1.n26 0.155672
R2452 VDD1.n43 VDD1.n26 0.155672
R2453 VDD1.n43 VDD1.n42 0.155672
R2454 VDD1.n42 VDD1.n30 0.155672
R2455 VDD1.n35 VDD1.n30 0.155672
R2456 VDD1.n135 VDD1.n130 0.155672
R2457 VDD1.n142 VDD1.n130 0.155672
R2458 VDD1.n143 VDD1.n142 0.155672
R2459 VDD1.n143 VDD1.n126 0.155672
R2460 VDD1.n150 VDD1.n126 0.155672
R2461 VDD1.n151 VDD1.n150 0.155672
R2462 VDD1.n151 VDD1.n122 0.155672
R2463 VDD1.n158 VDD1.n122 0.155672
R2464 VDD1.n159 VDD1.n158 0.155672
R2465 VDD1.n159 VDD1.n118 0.155672
R2466 VDD1.n166 VDD1.n118 0.155672
R2467 VDD1.n167 VDD1.n166 0.155672
R2468 VDD1.n167 VDD1.n114 0.155672
R2469 VDD1.n174 VDD1.n114 0.155672
R2470 VDD1.n175 VDD1.n174 0.155672
R2471 VDD1.n175 VDD1.n110 0.155672
R2472 VDD1.n184 VDD1.n110 0.155672
R2473 VDD1.n185 VDD1.n184 0.155672
R2474 VDD1.n185 VDD1.n106 0.155672
R2475 VDD1.n192 VDD1.n106 0.155672
R2476 VDD1.n193 VDD1.n192 0.155672
R2477 VDD1.n193 VDD1.n102 0.155672
R2478 VDD1.n200 VDD1.n102 0.155672
R2479 VN.n2 VN.t5 525.255
R2480 VN.n10 VN.t2 525.255
R2481 VN.n6 VN.t1 506.608
R2482 VN.n14 VN.t0 506.608
R2483 VN.n1 VN.t3 465.003
R2484 VN.n9 VN.t4 465.003
R2485 VN.n7 VN.n6 161.3
R2486 VN.n15 VN.n14 161.3
R2487 VN.n13 VN.n8 161.3
R2488 VN.n12 VN.n11 161.3
R2489 VN.n5 VN.n0 161.3
R2490 VN.n4 VN.n3 161.3
R2491 VN.n5 VN.n4 51.1773
R2492 VN.n13 VN.n12 51.1773
R2493 VN VN.n15 47.4191
R2494 VN.n11 VN.n10 43.2994
R2495 VN.n3 VN.n2 43.2994
R2496 VN.n2 VN.n1 42.326
R2497 VN.n10 VN.n9 42.326
R2498 VN.n4 VN.n1 12.234
R2499 VN.n12 VN.n9 12.234
R2500 VN.n6 VN.n5 8.03383
R2501 VN.n14 VN.n13 8.03383
R2502 VN.n15 VN.n8 0.189894
R2503 VN.n11 VN.n8 0.189894
R2504 VN.n3 VN.n0 0.189894
R2505 VN.n7 VN.n0 0.189894
R2506 VN VN.n7 0.0516364
R2507 VDD2.n199 VDD2.n103 289.615
R2508 VDD2.n96 VDD2.n0 289.615
R2509 VDD2.n200 VDD2.n199 185
R2510 VDD2.n198 VDD2.n197 185
R2511 VDD2.n107 VDD2.n106 185
R2512 VDD2.n192 VDD2.n191 185
R2513 VDD2.n190 VDD2.n189 185
R2514 VDD2.n111 VDD2.n110 185
R2515 VDD2.n184 VDD2.n183 185
R2516 VDD2.n182 VDD2.n113 185
R2517 VDD2.n181 VDD2.n180 185
R2518 VDD2.n116 VDD2.n114 185
R2519 VDD2.n175 VDD2.n174 185
R2520 VDD2.n173 VDD2.n172 185
R2521 VDD2.n120 VDD2.n119 185
R2522 VDD2.n167 VDD2.n166 185
R2523 VDD2.n165 VDD2.n164 185
R2524 VDD2.n124 VDD2.n123 185
R2525 VDD2.n159 VDD2.n158 185
R2526 VDD2.n157 VDD2.n156 185
R2527 VDD2.n128 VDD2.n127 185
R2528 VDD2.n151 VDD2.n150 185
R2529 VDD2.n149 VDD2.n148 185
R2530 VDD2.n132 VDD2.n131 185
R2531 VDD2.n143 VDD2.n142 185
R2532 VDD2.n141 VDD2.n140 185
R2533 VDD2.n136 VDD2.n135 185
R2534 VDD2.n32 VDD2.n31 185
R2535 VDD2.n37 VDD2.n36 185
R2536 VDD2.n39 VDD2.n38 185
R2537 VDD2.n28 VDD2.n27 185
R2538 VDD2.n45 VDD2.n44 185
R2539 VDD2.n47 VDD2.n46 185
R2540 VDD2.n24 VDD2.n23 185
R2541 VDD2.n53 VDD2.n52 185
R2542 VDD2.n55 VDD2.n54 185
R2543 VDD2.n20 VDD2.n19 185
R2544 VDD2.n61 VDD2.n60 185
R2545 VDD2.n63 VDD2.n62 185
R2546 VDD2.n16 VDD2.n15 185
R2547 VDD2.n69 VDD2.n68 185
R2548 VDD2.n71 VDD2.n70 185
R2549 VDD2.n12 VDD2.n11 185
R2550 VDD2.n78 VDD2.n77 185
R2551 VDD2.n79 VDD2.n10 185
R2552 VDD2.n81 VDD2.n80 185
R2553 VDD2.n8 VDD2.n7 185
R2554 VDD2.n87 VDD2.n86 185
R2555 VDD2.n89 VDD2.n88 185
R2556 VDD2.n4 VDD2.n3 185
R2557 VDD2.n95 VDD2.n94 185
R2558 VDD2.n97 VDD2.n96 185
R2559 VDD2.n137 VDD2.t5 147.659
R2560 VDD2.n33 VDD2.t0 147.659
R2561 VDD2.n199 VDD2.n198 104.615
R2562 VDD2.n198 VDD2.n106 104.615
R2563 VDD2.n191 VDD2.n106 104.615
R2564 VDD2.n191 VDD2.n190 104.615
R2565 VDD2.n190 VDD2.n110 104.615
R2566 VDD2.n183 VDD2.n110 104.615
R2567 VDD2.n183 VDD2.n182 104.615
R2568 VDD2.n182 VDD2.n181 104.615
R2569 VDD2.n181 VDD2.n114 104.615
R2570 VDD2.n174 VDD2.n114 104.615
R2571 VDD2.n174 VDD2.n173 104.615
R2572 VDD2.n173 VDD2.n119 104.615
R2573 VDD2.n166 VDD2.n119 104.615
R2574 VDD2.n166 VDD2.n165 104.615
R2575 VDD2.n165 VDD2.n123 104.615
R2576 VDD2.n158 VDD2.n123 104.615
R2577 VDD2.n158 VDD2.n157 104.615
R2578 VDD2.n157 VDD2.n127 104.615
R2579 VDD2.n150 VDD2.n127 104.615
R2580 VDD2.n150 VDD2.n149 104.615
R2581 VDD2.n149 VDD2.n131 104.615
R2582 VDD2.n142 VDD2.n131 104.615
R2583 VDD2.n142 VDD2.n141 104.615
R2584 VDD2.n141 VDD2.n135 104.615
R2585 VDD2.n37 VDD2.n31 104.615
R2586 VDD2.n38 VDD2.n37 104.615
R2587 VDD2.n38 VDD2.n27 104.615
R2588 VDD2.n45 VDD2.n27 104.615
R2589 VDD2.n46 VDD2.n45 104.615
R2590 VDD2.n46 VDD2.n23 104.615
R2591 VDD2.n53 VDD2.n23 104.615
R2592 VDD2.n54 VDD2.n53 104.615
R2593 VDD2.n54 VDD2.n19 104.615
R2594 VDD2.n61 VDD2.n19 104.615
R2595 VDD2.n62 VDD2.n61 104.615
R2596 VDD2.n62 VDD2.n15 104.615
R2597 VDD2.n69 VDD2.n15 104.615
R2598 VDD2.n70 VDD2.n69 104.615
R2599 VDD2.n70 VDD2.n11 104.615
R2600 VDD2.n78 VDD2.n11 104.615
R2601 VDD2.n79 VDD2.n78 104.615
R2602 VDD2.n80 VDD2.n79 104.615
R2603 VDD2.n80 VDD2.n7 104.615
R2604 VDD2.n87 VDD2.n7 104.615
R2605 VDD2.n88 VDD2.n87 104.615
R2606 VDD2.n88 VDD2.n3 104.615
R2607 VDD2.n95 VDD2.n3 104.615
R2608 VDD2.n96 VDD2.n95 104.615
R2609 VDD2.n102 VDD2.n101 62.6141
R2610 VDD2 VDD2.n205 62.6112
R2611 VDD2.t5 VDD2.n135 52.3082
R2612 VDD2.t0 VDD2.n31 52.3082
R2613 VDD2.n102 VDD2.n100 51.3818
R2614 VDD2.n204 VDD2.n203 50.6096
R2615 VDD2.n204 VDD2.n102 43.1032
R2616 VDD2.n137 VDD2.n136 15.6677
R2617 VDD2.n33 VDD2.n32 15.6677
R2618 VDD2.n184 VDD2.n113 13.1884
R2619 VDD2.n81 VDD2.n10 13.1884
R2620 VDD2.n185 VDD2.n111 12.8005
R2621 VDD2.n180 VDD2.n115 12.8005
R2622 VDD2.n140 VDD2.n139 12.8005
R2623 VDD2.n36 VDD2.n35 12.8005
R2624 VDD2.n77 VDD2.n76 12.8005
R2625 VDD2.n82 VDD2.n8 12.8005
R2626 VDD2.n189 VDD2.n188 12.0247
R2627 VDD2.n179 VDD2.n116 12.0247
R2628 VDD2.n143 VDD2.n134 12.0247
R2629 VDD2.n39 VDD2.n30 12.0247
R2630 VDD2.n75 VDD2.n12 12.0247
R2631 VDD2.n86 VDD2.n85 12.0247
R2632 VDD2.n192 VDD2.n109 11.249
R2633 VDD2.n176 VDD2.n175 11.249
R2634 VDD2.n144 VDD2.n132 11.249
R2635 VDD2.n40 VDD2.n28 11.249
R2636 VDD2.n72 VDD2.n71 11.249
R2637 VDD2.n89 VDD2.n6 11.249
R2638 VDD2.n193 VDD2.n107 10.4732
R2639 VDD2.n172 VDD2.n118 10.4732
R2640 VDD2.n148 VDD2.n147 10.4732
R2641 VDD2.n44 VDD2.n43 10.4732
R2642 VDD2.n68 VDD2.n14 10.4732
R2643 VDD2.n90 VDD2.n4 10.4732
R2644 VDD2.n197 VDD2.n196 9.69747
R2645 VDD2.n171 VDD2.n120 9.69747
R2646 VDD2.n151 VDD2.n130 9.69747
R2647 VDD2.n47 VDD2.n26 9.69747
R2648 VDD2.n67 VDD2.n16 9.69747
R2649 VDD2.n94 VDD2.n93 9.69747
R2650 VDD2.n203 VDD2.n202 9.45567
R2651 VDD2.n100 VDD2.n99 9.45567
R2652 VDD2.n163 VDD2.n162 9.3005
R2653 VDD2.n122 VDD2.n121 9.3005
R2654 VDD2.n169 VDD2.n168 9.3005
R2655 VDD2.n171 VDD2.n170 9.3005
R2656 VDD2.n118 VDD2.n117 9.3005
R2657 VDD2.n177 VDD2.n176 9.3005
R2658 VDD2.n179 VDD2.n178 9.3005
R2659 VDD2.n115 VDD2.n112 9.3005
R2660 VDD2.n202 VDD2.n201 9.3005
R2661 VDD2.n105 VDD2.n104 9.3005
R2662 VDD2.n196 VDD2.n195 9.3005
R2663 VDD2.n194 VDD2.n193 9.3005
R2664 VDD2.n109 VDD2.n108 9.3005
R2665 VDD2.n188 VDD2.n187 9.3005
R2666 VDD2.n186 VDD2.n185 9.3005
R2667 VDD2.n161 VDD2.n160 9.3005
R2668 VDD2.n126 VDD2.n125 9.3005
R2669 VDD2.n155 VDD2.n154 9.3005
R2670 VDD2.n153 VDD2.n152 9.3005
R2671 VDD2.n130 VDD2.n129 9.3005
R2672 VDD2.n147 VDD2.n146 9.3005
R2673 VDD2.n145 VDD2.n144 9.3005
R2674 VDD2.n134 VDD2.n133 9.3005
R2675 VDD2.n139 VDD2.n138 9.3005
R2676 VDD2.n99 VDD2.n98 9.3005
R2677 VDD2.n2 VDD2.n1 9.3005
R2678 VDD2.n93 VDD2.n92 9.3005
R2679 VDD2.n91 VDD2.n90 9.3005
R2680 VDD2.n6 VDD2.n5 9.3005
R2681 VDD2.n85 VDD2.n84 9.3005
R2682 VDD2.n83 VDD2.n82 9.3005
R2683 VDD2.n22 VDD2.n21 9.3005
R2684 VDD2.n51 VDD2.n50 9.3005
R2685 VDD2.n49 VDD2.n48 9.3005
R2686 VDD2.n26 VDD2.n25 9.3005
R2687 VDD2.n43 VDD2.n42 9.3005
R2688 VDD2.n41 VDD2.n40 9.3005
R2689 VDD2.n30 VDD2.n29 9.3005
R2690 VDD2.n35 VDD2.n34 9.3005
R2691 VDD2.n57 VDD2.n56 9.3005
R2692 VDD2.n59 VDD2.n58 9.3005
R2693 VDD2.n18 VDD2.n17 9.3005
R2694 VDD2.n65 VDD2.n64 9.3005
R2695 VDD2.n67 VDD2.n66 9.3005
R2696 VDD2.n14 VDD2.n13 9.3005
R2697 VDD2.n73 VDD2.n72 9.3005
R2698 VDD2.n75 VDD2.n74 9.3005
R2699 VDD2.n76 VDD2.n9 9.3005
R2700 VDD2.n200 VDD2.n105 8.92171
R2701 VDD2.n168 VDD2.n167 8.92171
R2702 VDD2.n152 VDD2.n128 8.92171
R2703 VDD2.n48 VDD2.n24 8.92171
R2704 VDD2.n64 VDD2.n63 8.92171
R2705 VDD2.n97 VDD2.n2 8.92171
R2706 VDD2.n201 VDD2.n103 8.14595
R2707 VDD2.n164 VDD2.n122 8.14595
R2708 VDD2.n156 VDD2.n155 8.14595
R2709 VDD2.n52 VDD2.n51 8.14595
R2710 VDD2.n60 VDD2.n18 8.14595
R2711 VDD2.n98 VDD2.n0 8.14595
R2712 VDD2.n163 VDD2.n124 7.3702
R2713 VDD2.n159 VDD2.n126 7.3702
R2714 VDD2.n55 VDD2.n22 7.3702
R2715 VDD2.n59 VDD2.n20 7.3702
R2716 VDD2.n160 VDD2.n124 6.59444
R2717 VDD2.n160 VDD2.n159 6.59444
R2718 VDD2.n56 VDD2.n55 6.59444
R2719 VDD2.n56 VDD2.n20 6.59444
R2720 VDD2.n203 VDD2.n103 5.81868
R2721 VDD2.n164 VDD2.n163 5.81868
R2722 VDD2.n156 VDD2.n126 5.81868
R2723 VDD2.n52 VDD2.n22 5.81868
R2724 VDD2.n60 VDD2.n59 5.81868
R2725 VDD2.n100 VDD2.n0 5.81868
R2726 VDD2.n201 VDD2.n200 5.04292
R2727 VDD2.n167 VDD2.n122 5.04292
R2728 VDD2.n155 VDD2.n128 5.04292
R2729 VDD2.n51 VDD2.n24 5.04292
R2730 VDD2.n63 VDD2.n18 5.04292
R2731 VDD2.n98 VDD2.n97 5.04292
R2732 VDD2.n138 VDD2.n137 4.38563
R2733 VDD2.n34 VDD2.n33 4.38563
R2734 VDD2.n197 VDD2.n105 4.26717
R2735 VDD2.n168 VDD2.n120 4.26717
R2736 VDD2.n152 VDD2.n151 4.26717
R2737 VDD2.n48 VDD2.n47 4.26717
R2738 VDD2.n64 VDD2.n16 4.26717
R2739 VDD2.n94 VDD2.n2 4.26717
R2740 VDD2.n196 VDD2.n107 3.49141
R2741 VDD2.n172 VDD2.n171 3.49141
R2742 VDD2.n148 VDD2.n130 3.49141
R2743 VDD2.n44 VDD2.n26 3.49141
R2744 VDD2.n68 VDD2.n67 3.49141
R2745 VDD2.n93 VDD2.n4 3.49141
R2746 VDD2.n193 VDD2.n192 2.71565
R2747 VDD2.n175 VDD2.n118 2.71565
R2748 VDD2.n147 VDD2.n132 2.71565
R2749 VDD2.n43 VDD2.n28 2.71565
R2750 VDD2.n71 VDD2.n14 2.71565
R2751 VDD2.n90 VDD2.n89 2.71565
R2752 VDD2.n189 VDD2.n109 1.93989
R2753 VDD2.n176 VDD2.n116 1.93989
R2754 VDD2.n144 VDD2.n143 1.93989
R2755 VDD2.n40 VDD2.n39 1.93989
R2756 VDD2.n72 VDD2.n12 1.93989
R2757 VDD2.n86 VDD2.n6 1.93989
R2758 VDD2.n188 VDD2.n111 1.16414
R2759 VDD2.n180 VDD2.n179 1.16414
R2760 VDD2.n140 VDD2.n134 1.16414
R2761 VDD2.n36 VDD2.n30 1.16414
R2762 VDD2.n77 VDD2.n75 1.16414
R2763 VDD2.n85 VDD2.n8 1.16414
R2764 VDD2.n205 VDD2.t1 1.0807
R2765 VDD2.n205 VDD2.t3 1.0807
R2766 VDD2.n101 VDD2.t2 1.0807
R2767 VDD2.n101 VDD2.t4 1.0807
R2768 VDD2 VDD2.n204 0.886276
R2769 VDD2.n185 VDD2.n184 0.388379
R2770 VDD2.n115 VDD2.n113 0.388379
R2771 VDD2.n139 VDD2.n136 0.388379
R2772 VDD2.n35 VDD2.n32 0.388379
R2773 VDD2.n76 VDD2.n10 0.388379
R2774 VDD2.n82 VDD2.n81 0.388379
R2775 VDD2.n202 VDD2.n104 0.155672
R2776 VDD2.n195 VDD2.n104 0.155672
R2777 VDD2.n195 VDD2.n194 0.155672
R2778 VDD2.n194 VDD2.n108 0.155672
R2779 VDD2.n187 VDD2.n108 0.155672
R2780 VDD2.n187 VDD2.n186 0.155672
R2781 VDD2.n186 VDD2.n112 0.155672
R2782 VDD2.n178 VDD2.n112 0.155672
R2783 VDD2.n178 VDD2.n177 0.155672
R2784 VDD2.n177 VDD2.n117 0.155672
R2785 VDD2.n170 VDD2.n117 0.155672
R2786 VDD2.n170 VDD2.n169 0.155672
R2787 VDD2.n169 VDD2.n121 0.155672
R2788 VDD2.n162 VDD2.n121 0.155672
R2789 VDD2.n162 VDD2.n161 0.155672
R2790 VDD2.n161 VDD2.n125 0.155672
R2791 VDD2.n154 VDD2.n125 0.155672
R2792 VDD2.n154 VDD2.n153 0.155672
R2793 VDD2.n153 VDD2.n129 0.155672
R2794 VDD2.n146 VDD2.n129 0.155672
R2795 VDD2.n146 VDD2.n145 0.155672
R2796 VDD2.n145 VDD2.n133 0.155672
R2797 VDD2.n138 VDD2.n133 0.155672
R2798 VDD2.n34 VDD2.n29 0.155672
R2799 VDD2.n41 VDD2.n29 0.155672
R2800 VDD2.n42 VDD2.n41 0.155672
R2801 VDD2.n42 VDD2.n25 0.155672
R2802 VDD2.n49 VDD2.n25 0.155672
R2803 VDD2.n50 VDD2.n49 0.155672
R2804 VDD2.n50 VDD2.n21 0.155672
R2805 VDD2.n57 VDD2.n21 0.155672
R2806 VDD2.n58 VDD2.n57 0.155672
R2807 VDD2.n58 VDD2.n17 0.155672
R2808 VDD2.n65 VDD2.n17 0.155672
R2809 VDD2.n66 VDD2.n65 0.155672
R2810 VDD2.n66 VDD2.n13 0.155672
R2811 VDD2.n73 VDD2.n13 0.155672
R2812 VDD2.n74 VDD2.n73 0.155672
R2813 VDD2.n74 VDD2.n9 0.155672
R2814 VDD2.n83 VDD2.n9 0.155672
R2815 VDD2.n84 VDD2.n83 0.155672
R2816 VDD2.n84 VDD2.n5 0.155672
R2817 VDD2.n91 VDD2.n5 0.155672
R2818 VDD2.n92 VDD2.n91 0.155672
R2819 VDD2.n92 VDD2.n1 0.155672
R2820 VDD2.n99 VDD2.n1 0.155672
C0 VN VDD1 0.148437f
C1 VTAIL VDD2 12.6084f
C2 VP VTAIL 6.94721f
C3 VN VTAIL 6.93245f
C4 VP VDD2 0.319542f
C5 VN VDD2 7.43263f
C6 VP VN 6.4932f
C7 VTAIL VDD1 12.574901f
C8 VDD1 VDD2 0.803199f
C9 VP VDD1 7.59756f
C10 VDD2 B 5.818553f
C11 VDD1 B 5.857514f
C12 VTAIL B 8.980268f
C13 VN B 9.048f
C14 VP B 6.942044f
C15 VDD2.n0 B 0.032818f
C16 VDD2.n1 B 0.022382f
C17 VDD2.n2 B 0.012027f
C18 VDD2.n3 B 0.028427f
C19 VDD2.n4 B 0.012734f
C20 VDD2.n5 B 0.022382f
C21 VDD2.n6 B 0.012027f
C22 VDD2.n7 B 0.028427f
C23 VDD2.n8 B 0.012734f
C24 VDD2.n9 B 0.022382f
C25 VDD2.n10 B 0.012381f
C26 VDD2.n11 B 0.028427f
C27 VDD2.n12 B 0.012734f
C28 VDD2.n13 B 0.022382f
C29 VDD2.n14 B 0.012027f
C30 VDD2.n15 B 0.028427f
C31 VDD2.n16 B 0.012734f
C32 VDD2.n17 B 0.022382f
C33 VDD2.n18 B 0.012027f
C34 VDD2.n19 B 0.028427f
C35 VDD2.n20 B 0.012734f
C36 VDD2.n21 B 0.022382f
C37 VDD2.n22 B 0.012027f
C38 VDD2.n23 B 0.028427f
C39 VDD2.n24 B 0.012734f
C40 VDD2.n25 B 0.022382f
C41 VDD2.n26 B 0.012027f
C42 VDD2.n27 B 0.028427f
C43 VDD2.n28 B 0.012734f
C44 VDD2.n29 B 0.022382f
C45 VDD2.n30 B 0.012027f
C46 VDD2.n31 B 0.02132f
C47 VDD2.n32 B 0.016793f
C48 VDD2.t0 B 0.047129f
C49 VDD2.n33 B 0.164665f
C50 VDD2.n34 B 1.79776f
C51 VDD2.n35 B 0.012027f
C52 VDD2.n36 B 0.012734f
C53 VDD2.n37 B 0.028427f
C54 VDD2.n38 B 0.028427f
C55 VDD2.n39 B 0.012734f
C56 VDD2.n40 B 0.012027f
C57 VDD2.n41 B 0.022382f
C58 VDD2.n42 B 0.022382f
C59 VDD2.n43 B 0.012027f
C60 VDD2.n44 B 0.012734f
C61 VDD2.n45 B 0.028427f
C62 VDD2.n46 B 0.028427f
C63 VDD2.n47 B 0.012734f
C64 VDD2.n48 B 0.012027f
C65 VDD2.n49 B 0.022382f
C66 VDD2.n50 B 0.022382f
C67 VDD2.n51 B 0.012027f
C68 VDD2.n52 B 0.012734f
C69 VDD2.n53 B 0.028427f
C70 VDD2.n54 B 0.028427f
C71 VDD2.n55 B 0.012734f
C72 VDD2.n56 B 0.012027f
C73 VDD2.n57 B 0.022382f
C74 VDD2.n58 B 0.022382f
C75 VDD2.n59 B 0.012027f
C76 VDD2.n60 B 0.012734f
C77 VDD2.n61 B 0.028427f
C78 VDD2.n62 B 0.028427f
C79 VDD2.n63 B 0.012734f
C80 VDD2.n64 B 0.012027f
C81 VDD2.n65 B 0.022382f
C82 VDD2.n66 B 0.022382f
C83 VDD2.n67 B 0.012027f
C84 VDD2.n68 B 0.012734f
C85 VDD2.n69 B 0.028427f
C86 VDD2.n70 B 0.028427f
C87 VDD2.n71 B 0.012734f
C88 VDD2.n72 B 0.012027f
C89 VDD2.n73 B 0.022382f
C90 VDD2.n74 B 0.022382f
C91 VDD2.n75 B 0.012027f
C92 VDD2.n76 B 0.012027f
C93 VDD2.n77 B 0.012734f
C94 VDD2.n78 B 0.028427f
C95 VDD2.n79 B 0.028427f
C96 VDD2.n80 B 0.028427f
C97 VDD2.n81 B 0.012381f
C98 VDD2.n82 B 0.012027f
C99 VDD2.n83 B 0.022382f
C100 VDD2.n84 B 0.022382f
C101 VDD2.n85 B 0.012027f
C102 VDD2.n86 B 0.012734f
C103 VDD2.n87 B 0.028427f
C104 VDD2.n88 B 0.028427f
C105 VDD2.n89 B 0.012734f
C106 VDD2.n90 B 0.012027f
C107 VDD2.n91 B 0.022382f
C108 VDD2.n92 B 0.022382f
C109 VDD2.n93 B 0.012027f
C110 VDD2.n94 B 0.012734f
C111 VDD2.n95 B 0.028427f
C112 VDD2.n96 B 0.063944f
C113 VDD2.n97 B 0.012734f
C114 VDD2.n98 B 0.012027f
C115 VDD2.n99 B 0.054486f
C116 VDD2.n100 B 0.053061f
C117 VDD2.t2 B 0.324197f
C118 VDD2.t4 B 0.324197f
C119 VDD2.n101 B 2.95819f
C120 VDD2.n102 B 2.10922f
C121 VDD2.n103 B 0.032818f
C122 VDD2.n104 B 0.022382f
C123 VDD2.n105 B 0.012027f
C124 VDD2.n106 B 0.028427f
C125 VDD2.n107 B 0.012734f
C126 VDD2.n108 B 0.022382f
C127 VDD2.n109 B 0.012027f
C128 VDD2.n110 B 0.028427f
C129 VDD2.n111 B 0.012734f
C130 VDD2.n112 B 0.022382f
C131 VDD2.n113 B 0.012381f
C132 VDD2.n114 B 0.028427f
C133 VDD2.n115 B 0.012027f
C134 VDD2.n116 B 0.012734f
C135 VDD2.n117 B 0.022382f
C136 VDD2.n118 B 0.012027f
C137 VDD2.n119 B 0.028427f
C138 VDD2.n120 B 0.012734f
C139 VDD2.n121 B 0.022382f
C140 VDD2.n122 B 0.012027f
C141 VDD2.n123 B 0.028427f
C142 VDD2.n124 B 0.012734f
C143 VDD2.n125 B 0.022382f
C144 VDD2.n126 B 0.012027f
C145 VDD2.n127 B 0.028427f
C146 VDD2.n128 B 0.012734f
C147 VDD2.n129 B 0.022382f
C148 VDD2.n130 B 0.012027f
C149 VDD2.n131 B 0.028427f
C150 VDD2.n132 B 0.012734f
C151 VDD2.n133 B 0.022382f
C152 VDD2.n134 B 0.012027f
C153 VDD2.n135 B 0.02132f
C154 VDD2.n136 B 0.016793f
C155 VDD2.t5 B 0.047129f
C156 VDD2.n137 B 0.164665f
C157 VDD2.n138 B 1.79776f
C158 VDD2.n139 B 0.012027f
C159 VDD2.n140 B 0.012734f
C160 VDD2.n141 B 0.028427f
C161 VDD2.n142 B 0.028427f
C162 VDD2.n143 B 0.012734f
C163 VDD2.n144 B 0.012027f
C164 VDD2.n145 B 0.022382f
C165 VDD2.n146 B 0.022382f
C166 VDD2.n147 B 0.012027f
C167 VDD2.n148 B 0.012734f
C168 VDD2.n149 B 0.028427f
C169 VDD2.n150 B 0.028427f
C170 VDD2.n151 B 0.012734f
C171 VDD2.n152 B 0.012027f
C172 VDD2.n153 B 0.022382f
C173 VDD2.n154 B 0.022382f
C174 VDD2.n155 B 0.012027f
C175 VDD2.n156 B 0.012734f
C176 VDD2.n157 B 0.028427f
C177 VDD2.n158 B 0.028427f
C178 VDD2.n159 B 0.012734f
C179 VDD2.n160 B 0.012027f
C180 VDD2.n161 B 0.022382f
C181 VDD2.n162 B 0.022382f
C182 VDD2.n163 B 0.012027f
C183 VDD2.n164 B 0.012734f
C184 VDD2.n165 B 0.028427f
C185 VDD2.n166 B 0.028427f
C186 VDD2.n167 B 0.012734f
C187 VDD2.n168 B 0.012027f
C188 VDD2.n169 B 0.022382f
C189 VDD2.n170 B 0.022382f
C190 VDD2.n171 B 0.012027f
C191 VDD2.n172 B 0.012734f
C192 VDD2.n173 B 0.028427f
C193 VDD2.n174 B 0.028427f
C194 VDD2.n175 B 0.012734f
C195 VDD2.n176 B 0.012027f
C196 VDD2.n177 B 0.022382f
C197 VDD2.n178 B 0.022382f
C198 VDD2.n179 B 0.012027f
C199 VDD2.n180 B 0.012734f
C200 VDD2.n181 B 0.028427f
C201 VDD2.n182 B 0.028427f
C202 VDD2.n183 B 0.028427f
C203 VDD2.n184 B 0.012381f
C204 VDD2.n185 B 0.012027f
C205 VDD2.n186 B 0.022382f
C206 VDD2.n187 B 0.022382f
C207 VDD2.n188 B 0.012027f
C208 VDD2.n189 B 0.012734f
C209 VDD2.n190 B 0.028427f
C210 VDD2.n191 B 0.028427f
C211 VDD2.n192 B 0.012734f
C212 VDD2.n193 B 0.012027f
C213 VDD2.n194 B 0.022382f
C214 VDD2.n195 B 0.022382f
C215 VDD2.n196 B 0.012027f
C216 VDD2.n197 B 0.012734f
C217 VDD2.n198 B 0.028427f
C218 VDD2.n199 B 0.063944f
C219 VDD2.n200 B 0.012734f
C220 VDD2.n201 B 0.012027f
C221 VDD2.n202 B 0.054486f
C222 VDD2.n203 B 0.051542f
C223 VDD2.n204 B 2.32819f
C224 VDD2.t1 B 0.324197f
C225 VDD2.t3 B 0.324197f
C226 VDD2.n205 B 2.95817f
C227 VN.n0 B 0.040014f
C228 VN.t3 B 1.91721f
C229 VN.n1 B 0.727004f
C230 VN.t5 B 2.00191f
C231 VN.n2 B 0.738345f
C232 VN.n3 B 0.171776f
C233 VN.n4 B 0.054242f
C234 VN.n5 B 0.014104f
C235 VN.t1 B 1.97545f
C236 VN.n6 B 0.734878f
C237 VN.n7 B 0.031009f
C238 VN.n8 B 0.040014f
C239 VN.t4 B 1.91721f
C240 VN.n9 B 0.727004f
C241 VN.t2 B 2.00191f
C242 VN.n10 B 0.738345f
C243 VN.n11 B 0.171776f
C244 VN.n12 B 0.054242f
C245 VN.n13 B 0.014104f
C246 VN.t0 B 1.97545f
C247 VN.n14 B 0.734878f
C248 VN.n15 B 2.00774f
C249 VDD1.n0 B 0.03301f
C250 VDD1.n1 B 0.022512f
C251 VDD1.n2 B 0.012097f
C252 VDD1.n3 B 0.028593f
C253 VDD1.n4 B 0.012809f
C254 VDD1.n5 B 0.022512f
C255 VDD1.n6 B 0.012097f
C256 VDD1.n7 B 0.028593f
C257 VDD1.n8 B 0.012809f
C258 VDD1.n9 B 0.022512f
C259 VDD1.n10 B 0.012453f
C260 VDD1.n11 B 0.028593f
C261 VDD1.n12 B 0.012097f
C262 VDD1.n13 B 0.012809f
C263 VDD1.n14 B 0.022512f
C264 VDD1.n15 B 0.012097f
C265 VDD1.n16 B 0.028593f
C266 VDD1.n17 B 0.012809f
C267 VDD1.n18 B 0.022512f
C268 VDD1.n19 B 0.012097f
C269 VDD1.n20 B 0.028593f
C270 VDD1.n21 B 0.012809f
C271 VDD1.n22 B 0.022512f
C272 VDD1.n23 B 0.012097f
C273 VDD1.n24 B 0.028593f
C274 VDD1.n25 B 0.012809f
C275 VDD1.n26 B 0.022512f
C276 VDD1.n27 B 0.012097f
C277 VDD1.n28 B 0.028593f
C278 VDD1.n29 B 0.012809f
C279 VDD1.n30 B 0.022512f
C280 VDD1.n31 B 0.012097f
C281 VDD1.n32 B 0.021445f
C282 VDD1.n33 B 0.016891f
C283 VDD1.t5 B 0.047404f
C284 VDD1.n34 B 0.165627f
C285 VDD1.n35 B 1.80826f
C286 VDD1.n36 B 0.012097f
C287 VDD1.n37 B 0.012809f
C288 VDD1.n38 B 0.028593f
C289 VDD1.n39 B 0.028593f
C290 VDD1.n40 B 0.012809f
C291 VDD1.n41 B 0.012097f
C292 VDD1.n42 B 0.022512f
C293 VDD1.n43 B 0.022512f
C294 VDD1.n44 B 0.012097f
C295 VDD1.n45 B 0.012809f
C296 VDD1.n46 B 0.028593f
C297 VDD1.n47 B 0.028593f
C298 VDD1.n48 B 0.012809f
C299 VDD1.n49 B 0.012097f
C300 VDD1.n50 B 0.022512f
C301 VDD1.n51 B 0.022512f
C302 VDD1.n52 B 0.012097f
C303 VDD1.n53 B 0.012809f
C304 VDD1.n54 B 0.028593f
C305 VDD1.n55 B 0.028593f
C306 VDD1.n56 B 0.012809f
C307 VDD1.n57 B 0.012097f
C308 VDD1.n58 B 0.022512f
C309 VDD1.n59 B 0.022512f
C310 VDD1.n60 B 0.012097f
C311 VDD1.n61 B 0.012809f
C312 VDD1.n62 B 0.028593f
C313 VDD1.n63 B 0.028593f
C314 VDD1.n64 B 0.012809f
C315 VDD1.n65 B 0.012097f
C316 VDD1.n66 B 0.022512f
C317 VDD1.n67 B 0.022512f
C318 VDD1.n68 B 0.012097f
C319 VDD1.n69 B 0.012809f
C320 VDD1.n70 B 0.028593f
C321 VDD1.n71 B 0.028593f
C322 VDD1.n72 B 0.012809f
C323 VDD1.n73 B 0.012097f
C324 VDD1.n74 B 0.022512f
C325 VDD1.n75 B 0.022512f
C326 VDD1.n76 B 0.012097f
C327 VDD1.n77 B 0.012809f
C328 VDD1.n78 B 0.028593f
C329 VDD1.n79 B 0.028593f
C330 VDD1.n80 B 0.028593f
C331 VDD1.n81 B 0.012453f
C332 VDD1.n82 B 0.012097f
C333 VDD1.n83 B 0.022512f
C334 VDD1.n84 B 0.022512f
C335 VDD1.n85 B 0.012097f
C336 VDD1.n86 B 0.012809f
C337 VDD1.n87 B 0.028593f
C338 VDD1.n88 B 0.028593f
C339 VDD1.n89 B 0.012809f
C340 VDD1.n90 B 0.012097f
C341 VDD1.n91 B 0.022512f
C342 VDD1.n92 B 0.022512f
C343 VDD1.n93 B 0.012097f
C344 VDD1.n94 B 0.012809f
C345 VDD1.n95 B 0.028593f
C346 VDD1.n96 B 0.064317f
C347 VDD1.n97 B 0.012809f
C348 VDD1.n98 B 0.012097f
C349 VDD1.n99 B 0.054804f
C350 VDD1.n100 B 0.053721f
C351 VDD1.n101 B 0.03301f
C352 VDD1.n102 B 0.022512f
C353 VDD1.n103 B 0.012097f
C354 VDD1.n104 B 0.028593f
C355 VDD1.n105 B 0.012809f
C356 VDD1.n106 B 0.022512f
C357 VDD1.n107 B 0.012097f
C358 VDD1.n108 B 0.028593f
C359 VDD1.n109 B 0.012809f
C360 VDD1.n110 B 0.022512f
C361 VDD1.n111 B 0.012453f
C362 VDD1.n112 B 0.028593f
C363 VDD1.n113 B 0.012809f
C364 VDD1.n114 B 0.022512f
C365 VDD1.n115 B 0.012097f
C366 VDD1.n116 B 0.028593f
C367 VDD1.n117 B 0.012809f
C368 VDD1.n118 B 0.022512f
C369 VDD1.n119 B 0.012097f
C370 VDD1.n120 B 0.028593f
C371 VDD1.n121 B 0.012809f
C372 VDD1.n122 B 0.022512f
C373 VDD1.n123 B 0.012097f
C374 VDD1.n124 B 0.028593f
C375 VDD1.n125 B 0.012809f
C376 VDD1.n126 B 0.022512f
C377 VDD1.n127 B 0.012097f
C378 VDD1.n128 B 0.028593f
C379 VDD1.n129 B 0.012809f
C380 VDD1.n130 B 0.022512f
C381 VDD1.n131 B 0.012097f
C382 VDD1.n132 B 0.021445f
C383 VDD1.n133 B 0.016891f
C384 VDD1.t4 B 0.047404f
C385 VDD1.n134 B 0.165627f
C386 VDD1.n135 B 1.80826f
C387 VDD1.n136 B 0.012097f
C388 VDD1.n137 B 0.012809f
C389 VDD1.n138 B 0.028593f
C390 VDD1.n139 B 0.028593f
C391 VDD1.n140 B 0.012809f
C392 VDD1.n141 B 0.012097f
C393 VDD1.n142 B 0.022512f
C394 VDD1.n143 B 0.022512f
C395 VDD1.n144 B 0.012097f
C396 VDD1.n145 B 0.012809f
C397 VDD1.n146 B 0.028593f
C398 VDD1.n147 B 0.028593f
C399 VDD1.n148 B 0.012809f
C400 VDD1.n149 B 0.012097f
C401 VDD1.n150 B 0.022512f
C402 VDD1.n151 B 0.022512f
C403 VDD1.n152 B 0.012097f
C404 VDD1.n153 B 0.012809f
C405 VDD1.n154 B 0.028593f
C406 VDD1.n155 B 0.028593f
C407 VDD1.n156 B 0.012809f
C408 VDD1.n157 B 0.012097f
C409 VDD1.n158 B 0.022512f
C410 VDD1.n159 B 0.022512f
C411 VDD1.n160 B 0.012097f
C412 VDD1.n161 B 0.012809f
C413 VDD1.n162 B 0.028593f
C414 VDD1.n163 B 0.028593f
C415 VDD1.n164 B 0.012809f
C416 VDD1.n165 B 0.012097f
C417 VDD1.n166 B 0.022512f
C418 VDD1.n167 B 0.022512f
C419 VDD1.n168 B 0.012097f
C420 VDD1.n169 B 0.012809f
C421 VDD1.n170 B 0.028593f
C422 VDD1.n171 B 0.028593f
C423 VDD1.n172 B 0.012809f
C424 VDD1.n173 B 0.012097f
C425 VDD1.n174 B 0.022512f
C426 VDD1.n175 B 0.022512f
C427 VDD1.n176 B 0.012097f
C428 VDD1.n177 B 0.012097f
C429 VDD1.n178 B 0.012809f
C430 VDD1.n179 B 0.028593f
C431 VDD1.n180 B 0.028593f
C432 VDD1.n181 B 0.028593f
C433 VDD1.n182 B 0.012453f
C434 VDD1.n183 B 0.012097f
C435 VDD1.n184 B 0.022512f
C436 VDD1.n185 B 0.022512f
C437 VDD1.n186 B 0.012097f
C438 VDD1.n187 B 0.012809f
C439 VDD1.n188 B 0.028593f
C440 VDD1.n189 B 0.028593f
C441 VDD1.n190 B 0.012809f
C442 VDD1.n191 B 0.012097f
C443 VDD1.n192 B 0.022512f
C444 VDD1.n193 B 0.022512f
C445 VDD1.n194 B 0.012097f
C446 VDD1.n195 B 0.012809f
C447 VDD1.n196 B 0.028593f
C448 VDD1.n197 B 0.064317f
C449 VDD1.n198 B 0.012809f
C450 VDD1.n199 B 0.012097f
C451 VDD1.n200 B 0.054804f
C452 VDD1.n201 B 0.053371f
C453 VDD1.t3 B 0.326091f
C454 VDD1.t1 B 0.326091f
C455 VDD1.n202 B 2.97548f
C456 VDD1.n203 B 2.19811f
C457 VDD1.t2 B 0.326091f
C458 VDD1.t0 B 0.326091f
C459 VDD1.n204 B 2.97444f
C460 VDD1.n205 B 2.52973f
C461 VTAIL.t2 B 0.330951f
C462 VTAIL.t4 B 0.330951f
C463 VTAIL.n0 B 2.95162f
C464 VTAIL.n1 B 0.324312f
C465 VTAIL.n2 B 0.033502f
C466 VTAIL.n3 B 0.022848f
C467 VTAIL.n4 B 0.012277f
C468 VTAIL.n5 B 0.02902f
C469 VTAIL.n6 B 0.013f
C470 VTAIL.n7 B 0.022848f
C471 VTAIL.n8 B 0.012277f
C472 VTAIL.n9 B 0.02902f
C473 VTAIL.n10 B 0.013f
C474 VTAIL.n11 B 0.022848f
C475 VTAIL.n12 B 0.012639f
C476 VTAIL.n13 B 0.02902f
C477 VTAIL.n14 B 0.013f
C478 VTAIL.n15 B 0.022848f
C479 VTAIL.n16 B 0.012277f
C480 VTAIL.n17 B 0.02902f
C481 VTAIL.n18 B 0.013f
C482 VTAIL.n19 B 0.022848f
C483 VTAIL.n20 B 0.012277f
C484 VTAIL.n21 B 0.02902f
C485 VTAIL.n22 B 0.013f
C486 VTAIL.n23 B 0.022848f
C487 VTAIL.n24 B 0.012277f
C488 VTAIL.n25 B 0.02902f
C489 VTAIL.n26 B 0.013f
C490 VTAIL.n27 B 0.022848f
C491 VTAIL.n28 B 0.012277f
C492 VTAIL.n29 B 0.02902f
C493 VTAIL.n30 B 0.013f
C494 VTAIL.n31 B 0.022848f
C495 VTAIL.n32 B 0.012277f
C496 VTAIL.n33 B 0.021765f
C497 VTAIL.n34 B 0.017143f
C498 VTAIL.t7 B 0.048111f
C499 VTAIL.n35 B 0.168095f
C500 VTAIL.n36 B 1.83521f
C501 VTAIL.n37 B 0.012277f
C502 VTAIL.n38 B 0.013f
C503 VTAIL.n39 B 0.02902f
C504 VTAIL.n40 B 0.02902f
C505 VTAIL.n41 B 0.013f
C506 VTAIL.n42 B 0.012277f
C507 VTAIL.n43 B 0.022848f
C508 VTAIL.n44 B 0.022848f
C509 VTAIL.n45 B 0.012277f
C510 VTAIL.n46 B 0.013f
C511 VTAIL.n47 B 0.02902f
C512 VTAIL.n48 B 0.02902f
C513 VTAIL.n49 B 0.013f
C514 VTAIL.n50 B 0.012277f
C515 VTAIL.n51 B 0.022848f
C516 VTAIL.n52 B 0.022848f
C517 VTAIL.n53 B 0.012277f
C518 VTAIL.n54 B 0.013f
C519 VTAIL.n55 B 0.02902f
C520 VTAIL.n56 B 0.02902f
C521 VTAIL.n57 B 0.013f
C522 VTAIL.n58 B 0.012277f
C523 VTAIL.n59 B 0.022848f
C524 VTAIL.n60 B 0.022848f
C525 VTAIL.n61 B 0.012277f
C526 VTAIL.n62 B 0.013f
C527 VTAIL.n63 B 0.02902f
C528 VTAIL.n64 B 0.02902f
C529 VTAIL.n65 B 0.013f
C530 VTAIL.n66 B 0.012277f
C531 VTAIL.n67 B 0.022848f
C532 VTAIL.n68 B 0.022848f
C533 VTAIL.n69 B 0.012277f
C534 VTAIL.n70 B 0.013f
C535 VTAIL.n71 B 0.02902f
C536 VTAIL.n72 B 0.02902f
C537 VTAIL.n73 B 0.013f
C538 VTAIL.n74 B 0.012277f
C539 VTAIL.n75 B 0.022848f
C540 VTAIL.n76 B 0.022848f
C541 VTAIL.n77 B 0.012277f
C542 VTAIL.n78 B 0.012277f
C543 VTAIL.n79 B 0.013f
C544 VTAIL.n80 B 0.02902f
C545 VTAIL.n81 B 0.02902f
C546 VTAIL.n82 B 0.02902f
C547 VTAIL.n83 B 0.012639f
C548 VTAIL.n84 B 0.012277f
C549 VTAIL.n85 B 0.022848f
C550 VTAIL.n86 B 0.022848f
C551 VTAIL.n87 B 0.012277f
C552 VTAIL.n88 B 0.013f
C553 VTAIL.n89 B 0.02902f
C554 VTAIL.n90 B 0.02902f
C555 VTAIL.n91 B 0.013f
C556 VTAIL.n92 B 0.012277f
C557 VTAIL.n93 B 0.022848f
C558 VTAIL.n94 B 0.022848f
C559 VTAIL.n95 B 0.012277f
C560 VTAIL.n96 B 0.013f
C561 VTAIL.n97 B 0.02902f
C562 VTAIL.n98 B 0.065276f
C563 VTAIL.n99 B 0.013f
C564 VTAIL.n100 B 0.012277f
C565 VTAIL.n101 B 0.055621f
C566 VTAIL.n102 B 0.036861f
C567 VTAIL.n103 B 0.177546f
C568 VTAIL.t6 B 0.330951f
C569 VTAIL.t5 B 0.330951f
C570 VTAIL.n104 B 2.95162f
C571 VTAIL.n105 B 1.94193f
C572 VTAIL.t11 B 0.330951f
C573 VTAIL.t3 B 0.330951f
C574 VTAIL.n106 B 2.95163f
C575 VTAIL.n107 B 1.94191f
C576 VTAIL.n108 B 0.033502f
C577 VTAIL.n109 B 0.022848f
C578 VTAIL.n110 B 0.012277f
C579 VTAIL.n111 B 0.02902f
C580 VTAIL.n112 B 0.013f
C581 VTAIL.n113 B 0.022848f
C582 VTAIL.n114 B 0.012277f
C583 VTAIL.n115 B 0.02902f
C584 VTAIL.n116 B 0.013f
C585 VTAIL.n117 B 0.022848f
C586 VTAIL.n118 B 0.012639f
C587 VTAIL.n119 B 0.02902f
C588 VTAIL.n120 B 0.012277f
C589 VTAIL.n121 B 0.013f
C590 VTAIL.n122 B 0.022848f
C591 VTAIL.n123 B 0.012277f
C592 VTAIL.n124 B 0.02902f
C593 VTAIL.n125 B 0.013f
C594 VTAIL.n126 B 0.022848f
C595 VTAIL.n127 B 0.012277f
C596 VTAIL.n128 B 0.02902f
C597 VTAIL.n129 B 0.013f
C598 VTAIL.n130 B 0.022848f
C599 VTAIL.n131 B 0.012277f
C600 VTAIL.n132 B 0.02902f
C601 VTAIL.n133 B 0.013f
C602 VTAIL.n134 B 0.022848f
C603 VTAIL.n135 B 0.012277f
C604 VTAIL.n136 B 0.02902f
C605 VTAIL.n137 B 0.013f
C606 VTAIL.n138 B 0.022848f
C607 VTAIL.n139 B 0.012277f
C608 VTAIL.n140 B 0.021765f
C609 VTAIL.n141 B 0.017143f
C610 VTAIL.t1 B 0.048111f
C611 VTAIL.n142 B 0.168095f
C612 VTAIL.n143 B 1.83521f
C613 VTAIL.n144 B 0.012277f
C614 VTAIL.n145 B 0.013f
C615 VTAIL.n146 B 0.02902f
C616 VTAIL.n147 B 0.02902f
C617 VTAIL.n148 B 0.013f
C618 VTAIL.n149 B 0.012277f
C619 VTAIL.n150 B 0.022848f
C620 VTAIL.n151 B 0.022848f
C621 VTAIL.n152 B 0.012277f
C622 VTAIL.n153 B 0.013f
C623 VTAIL.n154 B 0.02902f
C624 VTAIL.n155 B 0.02902f
C625 VTAIL.n156 B 0.013f
C626 VTAIL.n157 B 0.012277f
C627 VTAIL.n158 B 0.022848f
C628 VTAIL.n159 B 0.022848f
C629 VTAIL.n160 B 0.012277f
C630 VTAIL.n161 B 0.013f
C631 VTAIL.n162 B 0.02902f
C632 VTAIL.n163 B 0.02902f
C633 VTAIL.n164 B 0.013f
C634 VTAIL.n165 B 0.012277f
C635 VTAIL.n166 B 0.022848f
C636 VTAIL.n167 B 0.022848f
C637 VTAIL.n168 B 0.012277f
C638 VTAIL.n169 B 0.013f
C639 VTAIL.n170 B 0.02902f
C640 VTAIL.n171 B 0.02902f
C641 VTAIL.n172 B 0.013f
C642 VTAIL.n173 B 0.012277f
C643 VTAIL.n174 B 0.022848f
C644 VTAIL.n175 B 0.022848f
C645 VTAIL.n176 B 0.012277f
C646 VTAIL.n177 B 0.013f
C647 VTAIL.n178 B 0.02902f
C648 VTAIL.n179 B 0.02902f
C649 VTAIL.n180 B 0.013f
C650 VTAIL.n181 B 0.012277f
C651 VTAIL.n182 B 0.022848f
C652 VTAIL.n183 B 0.022848f
C653 VTAIL.n184 B 0.012277f
C654 VTAIL.n185 B 0.013f
C655 VTAIL.n186 B 0.02902f
C656 VTAIL.n187 B 0.02902f
C657 VTAIL.n188 B 0.02902f
C658 VTAIL.n189 B 0.012639f
C659 VTAIL.n190 B 0.012277f
C660 VTAIL.n191 B 0.022848f
C661 VTAIL.n192 B 0.022848f
C662 VTAIL.n193 B 0.012277f
C663 VTAIL.n194 B 0.013f
C664 VTAIL.n195 B 0.02902f
C665 VTAIL.n196 B 0.02902f
C666 VTAIL.n197 B 0.013f
C667 VTAIL.n198 B 0.012277f
C668 VTAIL.n199 B 0.022848f
C669 VTAIL.n200 B 0.022848f
C670 VTAIL.n201 B 0.012277f
C671 VTAIL.n202 B 0.013f
C672 VTAIL.n203 B 0.02902f
C673 VTAIL.n204 B 0.065276f
C674 VTAIL.n205 B 0.013f
C675 VTAIL.n206 B 0.012277f
C676 VTAIL.n207 B 0.055621f
C677 VTAIL.n208 B 0.036861f
C678 VTAIL.n209 B 0.177546f
C679 VTAIL.t9 B 0.330951f
C680 VTAIL.t10 B 0.330951f
C681 VTAIL.n210 B 2.95163f
C682 VTAIL.n211 B 0.380943f
C683 VTAIL.n212 B 0.033502f
C684 VTAIL.n213 B 0.022848f
C685 VTAIL.n214 B 0.012277f
C686 VTAIL.n215 B 0.02902f
C687 VTAIL.n216 B 0.013f
C688 VTAIL.n217 B 0.022848f
C689 VTAIL.n218 B 0.012277f
C690 VTAIL.n219 B 0.02902f
C691 VTAIL.n220 B 0.013f
C692 VTAIL.n221 B 0.022848f
C693 VTAIL.n222 B 0.012639f
C694 VTAIL.n223 B 0.02902f
C695 VTAIL.n224 B 0.012277f
C696 VTAIL.n225 B 0.013f
C697 VTAIL.n226 B 0.022848f
C698 VTAIL.n227 B 0.012277f
C699 VTAIL.n228 B 0.02902f
C700 VTAIL.n229 B 0.013f
C701 VTAIL.n230 B 0.022848f
C702 VTAIL.n231 B 0.012277f
C703 VTAIL.n232 B 0.02902f
C704 VTAIL.n233 B 0.013f
C705 VTAIL.n234 B 0.022848f
C706 VTAIL.n235 B 0.012277f
C707 VTAIL.n236 B 0.02902f
C708 VTAIL.n237 B 0.013f
C709 VTAIL.n238 B 0.022848f
C710 VTAIL.n239 B 0.012277f
C711 VTAIL.n240 B 0.02902f
C712 VTAIL.n241 B 0.013f
C713 VTAIL.n242 B 0.022848f
C714 VTAIL.n243 B 0.012277f
C715 VTAIL.n244 B 0.021765f
C716 VTAIL.n245 B 0.017143f
C717 VTAIL.t8 B 0.048111f
C718 VTAIL.n246 B 0.168095f
C719 VTAIL.n247 B 1.83521f
C720 VTAIL.n248 B 0.012277f
C721 VTAIL.n249 B 0.013f
C722 VTAIL.n250 B 0.02902f
C723 VTAIL.n251 B 0.02902f
C724 VTAIL.n252 B 0.013f
C725 VTAIL.n253 B 0.012277f
C726 VTAIL.n254 B 0.022848f
C727 VTAIL.n255 B 0.022848f
C728 VTAIL.n256 B 0.012277f
C729 VTAIL.n257 B 0.013f
C730 VTAIL.n258 B 0.02902f
C731 VTAIL.n259 B 0.02902f
C732 VTAIL.n260 B 0.013f
C733 VTAIL.n261 B 0.012277f
C734 VTAIL.n262 B 0.022848f
C735 VTAIL.n263 B 0.022848f
C736 VTAIL.n264 B 0.012277f
C737 VTAIL.n265 B 0.013f
C738 VTAIL.n266 B 0.02902f
C739 VTAIL.n267 B 0.02902f
C740 VTAIL.n268 B 0.013f
C741 VTAIL.n269 B 0.012277f
C742 VTAIL.n270 B 0.022848f
C743 VTAIL.n271 B 0.022848f
C744 VTAIL.n272 B 0.012277f
C745 VTAIL.n273 B 0.013f
C746 VTAIL.n274 B 0.02902f
C747 VTAIL.n275 B 0.02902f
C748 VTAIL.n276 B 0.013f
C749 VTAIL.n277 B 0.012277f
C750 VTAIL.n278 B 0.022848f
C751 VTAIL.n279 B 0.022848f
C752 VTAIL.n280 B 0.012277f
C753 VTAIL.n281 B 0.013f
C754 VTAIL.n282 B 0.02902f
C755 VTAIL.n283 B 0.02902f
C756 VTAIL.n284 B 0.013f
C757 VTAIL.n285 B 0.012277f
C758 VTAIL.n286 B 0.022848f
C759 VTAIL.n287 B 0.022848f
C760 VTAIL.n288 B 0.012277f
C761 VTAIL.n289 B 0.013f
C762 VTAIL.n290 B 0.02902f
C763 VTAIL.n291 B 0.02902f
C764 VTAIL.n292 B 0.02902f
C765 VTAIL.n293 B 0.012639f
C766 VTAIL.n294 B 0.012277f
C767 VTAIL.n295 B 0.022848f
C768 VTAIL.n296 B 0.022848f
C769 VTAIL.n297 B 0.012277f
C770 VTAIL.n298 B 0.013f
C771 VTAIL.n299 B 0.02902f
C772 VTAIL.n300 B 0.02902f
C773 VTAIL.n301 B 0.013f
C774 VTAIL.n302 B 0.012277f
C775 VTAIL.n303 B 0.022848f
C776 VTAIL.n304 B 0.022848f
C777 VTAIL.n305 B 0.012277f
C778 VTAIL.n306 B 0.013f
C779 VTAIL.n307 B 0.02902f
C780 VTAIL.n308 B 0.065276f
C781 VTAIL.n309 B 0.013f
C782 VTAIL.n310 B 0.012277f
C783 VTAIL.n311 B 0.055621f
C784 VTAIL.n312 B 0.036861f
C785 VTAIL.n313 B 1.65728f
C786 VTAIL.n314 B 0.033502f
C787 VTAIL.n315 B 0.022848f
C788 VTAIL.n316 B 0.012277f
C789 VTAIL.n317 B 0.02902f
C790 VTAIL.n318 B 0.013f
C791 VTAIL.n319 B 0.022848f
C792 VTAIL.n320 B 0.012277f
C793 VTAIL.n321 B 0.02902f
C794 VTAIL.n322 B 0.013f
C795 VTAIL.n323 B 0.022848f
C796 VTAIL.n324 B 0.012639f
C797 VTAIL.n325 B 0.02902f
C798 VTAIL.n326 B 0.013f
C799 VTAIL.n327 B 0.022848f
C800 VTAIL.n328 B 0.012277f
C801 VTAIL.n329 B 0.02902f
C802 VTAIL.n330 B 0.013f
C803 VTAIL.n331 B 0.022848f
C804 VTAIL.n332 B 0.012277f
C805 VTAIL.n333 B 0.02902f
C806 VTAIL.n334 B 0.013f
C807 VTAIL.n335 B 0.022848f
C808 VTAIL.n336 B 0.012277f
C809 VTAIL.n337 B 0.02902f
C810 VTAIL.n338 B 0.013f
C811 VTAIL.n339 B 0.022848f
C812 VTAIL.n340 B 0.012277f
C813 VTAIL.n341 B 0.02902f
C814 VTAIL.n342 B 0.013f
C815 VTAIL.n343 B 0.022848f
C816 VTAIL.n344 B 0.012277f
C817 VTAIL.n345 B 0.021765f
C818 VTAIL.n346 B 0.017143f
C819 VTAIL.t0 B 0.048111f
C820 VTAIL.n347 B 0.168095f
C821 VTAIL.n348 B 1.83521f
C822 VTAIL.n349 B 0.012277f
C823 VTAIL.n350 B 0.013f
C824 VTAIL.n351 B 0.02902f
C825 VTAIL.n352 B 0.02902f
C826 VTAIL.n353 B 0.013f
C827 VTAIL.n354 B 0.012277f
C828 VTAIL.n355 B 0.022848f
C829 VTAIL.n356 B 0.022848f
C830 VTAIL.n357 B 0.012277f
C831 VTAIL.n358 B 0.013f
C832 VTAIL.n359 B 0.02902f
C833 VTAIL.n360 B 0.02902f
C834 VTAIL.n361 B 0.013f
C835 VTAIL.n362 B 0.012277f
C836 VTAIL.n363 B 0.022848f
C837 VTAIL.n364 B 0.022848f
C838 VTAIL.n365 B 0.012277f
C839 VTAIL.n366 B 0.013f
C840 VTAIL.n367 B 0.02902f
C841 VTAIL.n368 B 0.02902f
C842 VTAIL.n369 B 0.013f
C843 VTAIL.n370 B 0.012277f
C844 VTAIL.n371 B 0.022848f
C845 VTAIL.n372 B 0.022848f
C846 VTAIL.n373 B 0.012277f
C847 VTAIL.n374 B 0.013f
C848 VTAIL.n375 B 0.02902f
C849 VTAIL.n376 B 0.02902f
C850 VTAIL.n377 B 0.013f
C851 VTAIL.n378 B 0.012277f
C852 VTAIL.n379 B 0.022848f
C853 VTAIL.n380 B 0.022848f
C854 VTAIL.n381 B 0.012277f
C855 VTAIL.n382 B 0.013f
C856 VTAIL.n383 B 0.02902f
C857 VTAIL.n384 B 0.02902f
C858 VTAIL.n385 B 0.013f
C859 VTAIL.n386 B 0.012277f
C860 VTAIL.n387 B 0.022848f
C861 VTAIL.n388 B 0.022848f
C862 VTAIL.n389 B 0.012277f
C863 VTAIL.n390 B 0.012277f
C864 VTAIL.n391 B 0.013f
C865 VTAIL.n392 B 0.02902f
C866 VTAIL.n393 B 0.02902f
C867 VTAIL.n394 B 0.02902f
C868 VTAIL.n395 B 0.012639f
C869 VTAIL.n396 B 0.012277f
C870 VTAIL.n397 B 0.022848f
C871 VTAIL.n398 B 0.022848f
C872 VTAIL.n399 B 0.012277f
C873 VTAIL.n400 B 0.013f
C874 VTAIL.n401 B 0.02902f
C875 VTAIL.n402 B 0.02902f
C876 VTAIL.n403 B 0.013f
C877 VTAIL.n404 B 0.012277f
C878 VTAIL.n405 B 0.022848f
C879 VTAIL.n406 B 0.022848f
C880 VTAIL.n407 B 0.012277f
C881 VTAIL.n408 B 0.013f
C882 VTAIL.n409 B 0.02902f
C883 VTAIL.n410 B 0.065276f
C884 VTAIL.n411 B 0.013f
C885 VTAIL.n412 B 0.012277f
C886 VTAIL.n413 B 0.055621f
C887 VTAIL.n414 B 0.036861f
C888 VTAIL.n415 B 1.63269f
C889 VP.n0 B 0.040509f
C890 VP.t2 B 1.9409f
C891 VP.n1 B 0.696222f
C892 VP.n2 B 0.040509f
C893 VP.n3 B 0.040509f
C894 VP.t5 B 1.99985f
C895 VP.t3 B 1.9409f
C896 VP.n4 B 0.735984f
C897 VP.t0 B 2.02664f
C898 VP.n5 B 0.747465f
C899 VP.n6 B 0.173898f
C900 VP.n7 B 0.054912f
C901 VP.n8 B 0.014278f
C902 VP.n9 B 0.743956f
C903 VP.n10 B 2.00613f
C904 VP.n11 B 2.03708f
C905 VP.t1 B 1.99985f
C906 VP.n12 B 0.743956f
C907 VP.n13 B 0.014278f
C908 VP.n14 B 0.054912f
C909 VP.n15 B 0.040509f
C910 VP.n16 B 0.040509f
C911 VP.n17 B 0.054912f
C912 VP.n18 B 0.014278f
C913 VP.t4 B 1.99985f
C914 VP.n19 B 0.743956f
C915 VP.n20 B 0.031392f
.ends

