* NGSPICE file created from diff_pair_sample_0223.ext - technology: sky130A

.subckt diff_pair_sample_0223 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=2.937 ps=18.13 w=17.8 l=0.18
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=0 ps=0 w=17.8 l=0.18
X2 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=2.937 ps=18.13 w=17.8 l=0.18
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=0 ps=0 w=17.8 l=0.18
X4 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=0 ps=0 w=17.8 l=0.18
X5 VDD1.t4 VP.t1 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=6.942 ps=36.38 w=17.8 l=0.18
X6 VTAIL.t2 VN.t1 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=2.937 ps=18.13 w=17.8 l=0.18
X7 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=6.942 ps=36.38 w=17.8 l=0.18
X8 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=6.942 ps=36.38 w=17.8 l=0.18
X9 VTAIL.t11 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=2.937 ps=18.13 w=17.8 l=0.18
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=0 ps=0 w=17.8 l=0.18
X11 VDD2.t0 VN.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=2.937 ps=18.13 w=17.8 l=0.18
X12 VTAIL.t8 VP.t2 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=2.937 ps=18.13 w=17.8 l=0.18
X13 VDD1.t2 VP.t3 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=6.942 pd=36.38 as=2.937 ps=18.13 w=17.8 l=0.18
X14 VDD1.t1 VP.t4 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=6.942 ps=36.38 w=17.8 l=0.18
X15 VTAIL.t5 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.937 pd=18.13 as=2.937 ps=18.13 w=17.8 l=0.18
R0 VP.n7 VP.t1 2595.25
R1 VP.n5 VP.t0 2595.25
R2 VP.n0 VP.t3 2595.25
R3 VP.n2 VP.t4 2595.25
R4 VP.n6 VP.t2 2557.28
R5 VP.n1 VP.t5 2557.28
R6 VP.n3 VP.n0 161.489
R7 VP.n8 VP.n7 161.3
R8 VP.n3 VP.n2 161.3
R9 VP.n5 VP.n4 161.3
R10 VP.n4 VP.n3 43.6028
R11 VP.n6 VP.n5 36.5157
R12 VP.n7 VP.n6 36.5157
R13 VP.n1 VP.n0 36.5157
R14 VP.n2 VP.n1 36.5157
R15 VP.n8 VP.n4 0.189894
R16 VP VP.n8 0.0516364
R17 VTAIL.n7 VTAIL.t3 43.546
R18 VTAIL.n11 VTAIL.t1 43.5458
R19 VTAIL.n2 VTAIL.t4 43.5458
R20 VTAIL.n10 VTAIL.t6 43.5458
R21 VTAIL.n9 VTAIL.n8 42.4337
R22 VTAIL.n6 VTAIL.n5 42.4337
R23 VTAIL.n1 VTAIL.n0 42.4335
R24 VTAIL.n4 VTAIL.n3 42.4335
R25 VTAIL.n6 VTAIL.n4 28.591
R26 VTAIL.n11 VTAIL.n10 28.1514
R27 VTAIL.n0 VTAIL.t0 1.11286
R28 VTAIL.n0 VTAIL.t2 1.11286
R29 VTAIL.n3 VTAIL.t7 1.11286
R30 VTAIL.n3 VTAIL.t8 1.11286
R31 VTAIL.n8 VTAIL.t9 1.11286
R32 VTAIL.n8 VTAIL.t5 1.11286
R33 VTAIL.n5 VTAIL.t10 1.11286
R34 VTAIL.n5 VTAIL.t11 1.11286
R35 VTAIL.n9 VTAIL.n7 0.690155
R36 VTAIL.n2 VTAIL.n1 0.690155
R37 VTAIL.n7 VTAIL.n6 0.440155
R38 VTAIL.n10 VTAIL.n9 0.440155
R39 VTAIL.n4 VTAIL.n2 0.440155
R40 VTAIL VTAIL.n11 0.272052
R41 VTAIL VTAIL.n1 0.168603
R42 VDD1 VDD1.t2 60.6128
R43 VDD1.n1 VDD1.t5 60.499
R44 VDD1.n1 VDD1.n0 59.1668
R45 VDD1.n3 VDD1.n2 59.1123
R46 VDD1.n3 VDD1.n1 41.2918
R47 VDD1.n2 VDD1.t0 1.11286
R48 VDD1.n2 VDD1.t1 1.11286
R49 VDD1.n0 VDD1.t3 1.11286
R50 VDD1.n0 VDD1.t4 1.11286
R51 VDD1 VDD1.n3 0.0522241
R52 B.n159 B.t14 2626.27
R53 B.n153 B.t10 2626.27
R54 B.n60 B.t6 2626.27
R55 B.n67 B.t17 2626.27
R56 B.n508 B.n507 585
R57 B.n508 B.n28 585
R58 B.n511 B.n510 585
R59 B.n512 B.n96 585
R60 B.n514 B.n513 585
R61 B.n516 B.n95 585
R62 B.n519 B.n518 585
R63 B.n520 B.n94 585
R64 B.n522 B.n521 585
R65 B.n524 B.n93 585
R66 B.n527 B.n526 585
R67 B.n528 B.n92 585
R68 B.n530 B.n529 585
R69 B.n532 B.n91 585
R70 B.n535 B.n534 585
R71 B.n536 B.n90 585
R72 B.n538 B.n537 585
R73 B.n540 B.n89 585
R74 B.n543 B.n542 585
R75 B.n544 B.n88 585
R76 B.n546 B.n545 585
R77 B.n548 B.n87 585
R78 B.n551 B.n550 585
R79 B.n552 B.n86 585
R80 B.n554 B.n553 585
R81 B.n556 B.n85 585
R82 B.n559 B.n558 585
R83 B.n560 B.n84 585
R84 B.n562 B.n561 585
R85 B.n564 B.n83 585
R86 B.n567 B.n566 585
R87 B.n568 B.n82 585
R88 B.n570 B.n569 585
R89 B.n572 B.n81 585
R90 B.n575 B.n574 585
R91 B.n576 B.n80 585
R92 B.n578 B.n577 585
R93 B.n580 B.n79 585
R94 B.n583 B.n582 585
R95 B.n584 B.n78 585
R96 B.n586 B.n585 585
R97 B.n588 B.n77 585
R98 B.n591 B.n590 585
R99 B.n592 B.n76 585
R100 B.n594 B.n593 585
R101 B.n596 B.n75 585
R102 B.n599 B.n598 585
R103 B.n600 B.n74 585
R104 B.n602 B.n601 585
R105 B.n604 B.n73 585
R106 B.n607 B.n606 585
R107 B.n608 B.n72 585
R108 B.n610 B.n609 585
R109 B.n612 B.n71 585
R110 B.n615 B.n614 585
R111 B.n616 B.n70 585
R112 B.n618 B.n617 585
R113 B.n620 B.n69 585
R114 B.n623 B.n622 585
R115 B.n624 B.n66 585
R116 B.n627 B.n626 585
R117 B.n629 B.n65 585
R118 B.n632 B.n631 585
R119 B.n633 B.n64 585
R120 B.n635 B.n634 585
R121 B.n637 B.n63 585
R122 B.n640 B.n639 585
R123 B.n641 B.n59 585
R124 B.n643 B.n642 585
R125 B.n645 B.n58 585
R126 B.n648 B.n647 585
R127 B.n649 B.n57 585
R128 B.n651 B.n650 585
R129 B.n653 B.n56 585
R130 B.n656 B.n655 585
R131 B.n657 B.n55 585
R132 B.n659 B.n658 585
R133 B.n661 B.n54 585
R134 B.n664 B.n663 585
R135 B.n665 B.n53 585
R136 B.n667 B.n666 585
R137 B.n669 B.n52 585
R138 B.n672 B.n671 585
R139 B.n673 B.n51 585
R140 B.n675 B.n674 585
R141 B.n677 B.n50 585
R142 B.n680 B.n679 585
R143 B.n681 B.n49 585
R144 B.n683 B.n682 585
R145 B.n685 B.n48 585
R146 B.n688 B.n687 585
R147 B.n689 B.n47 585
R148 B.n691 B.n690 585
R149 B.n693 B.n46 585
R150 B.n696 B.n695 585
R151 B.n697 B.n45 585
R152 B.n699 B.n698 585
R153 B.n701 B.n44 585
R154 B.n704 B.n703 585
R155 B.n705 B.n43 585
R156 B.n707 B.n706 585
R157 B.n709 B.n42 585
R158 B.n712 B.n711 585
R159 B.n713 B.n41 585
R160 B.n715 B.n714 585
R161 B.n717 B.n40 585
R162 B.n720 B.n719 585
R163 B.n721 B.n39 585
R164 B.n723 B.n722 585
R165 B.n725 B.n38 585
R166 B.n728 B.n727 585
R167 B.n729 B.n37 585
R168 B.n731 B.n730 585
R169 B.n733 B.n36 585
R170 B.n736 B.n735 585
R171 B.n737 B.n35 585
R172 B.n739 B.n738 585
R173 B.n741 B.n34 585
R174 B.n744 B.n743 585
R175 B.n745 B.n33 585
R176 B.n747 B.n746 585
R177 B.n749 B.n32 585
R178 B.n752 B.n751 585
R179 B.n753 B.n31 585
R180 B.n755 B.n754 585
R181 B.n757 B.n30 585
R182 B.n760 B.n759 585
R183 B.n761 B.n29 585
R184 B.n506 B.n27 585
R185 B.n764 B.n27 585
R186 B.n505 B.n26 585
R187 B.n765 B.n26 585
R188 B.n504 B.n25 585
R189 B.n766 B.n25 585
R190 B.n503 B.n502 585
R191 B.n502 B.n24 585
R192 B.n501 B.n20 585
R193 B.n772 B.n20 585
R194 B.n500 B.n19 585
R195 B.n773 B.n19 585
R196 B.n499 B.n18 585
R197 B.n774 B.n18 585
R198 B.n498 B.n497 585
R199 B.n497 B.n14 585
R200 B.n496 B.n13 585
R201 B.n780 B.n13 585
R202 B.n495 B.n12 585
R203 B.n781 B.n12 585
R204 B.n494 B.n11 585
R205 B.n782 B.n11 585
R206 B.n493 B.n492 585
R207 B.n492 B.n491 585
R208 B.n490 B.n7 585
R209 B.n788 B.n7 585
R210 B.n489 B.n6 585
R211 B.n789 B.n6 585
R212 B.n488 B.n5 585
R213 B.n790 B.n5 585
R214 B.n487 B.n486 585
R215 B.n486 B.n4 585
R216 B.n485 B.n97 585
R217 B.n485 B.n484 585
R218 B.n474 B.n98 585
R219 B.n477 B.n98 585
R220 B.n476 B.n475 585
R221 B.n478 B.n476 585
R222 B.n473 B.n103 585
R223 B.n103 B.n102 585
R224 B.n472 B.n471 585
R225 B.n471 B.n470 585
R226 B.n105 B.n104 585
R227 B.n106 B.n105 585
R228 B.n463 B.n462 585
R229 B.n464 B.n463 585
R230 B.n461 B.n111 585
R231 B.n111 B.n110 585
R232 B.n460 B.n459 585
R233 B.n459 B.n458 585
R234 B.n113 B.n112 585
R235 B.n451 B.n113 585
R236 B.n450 B.n449 585
R237 B.n452 B.n450 585
R238 B.n448 B.n118 585
R239 B.n118 B.n117 585
R240 B.n447 B.n446 585
R241 B.n446 B.n445 585
R242 B.n442 B.n122 585
R243 B.n441 B.n440 585
R244 B.n438 B.n123 585
R245 B.n438 B.n121 585
R246 B.n437 B.n436 585
R247 B.n435 B.n434 585
R248 B.n433 B.n125 585
R249 B.n431 B.n430 585
R250 B.n429 B.n126 585
R251 B.n428 B.n427 585
R252 B.n425 B.n127 585
R253 B.n423 B.n422 585
R254 B.n421 B.n128 585
R255 B.n420 B.n419 585
R256 B.n417 B.n129 585
R257 B.n415 B.n414 585
R258 B.n413 B.n130 585
R259 B.n412 B.n411 585
R260 B.n409 B.n131 585
R261 B.n407 B.n406 585
R262 B.n405 B.n132 585
R263 B.n404 B.n403 585
R264 B.n401 B.n133 585
R265 B.n399 B.n398 585
R266 B.n397 B.n134 585
R267 B.n396 B.n395 585
R268 B.n393 B.n135 585
R269 B.n391 B.n390 585
R270 B.n389 B.n136 585
R271 B.n388 B.n387 585
R272 B.n385 B.n137 585
R273 B.n383 B.n382 585
R274 B.n381 B.n138 585
R275 B.n380 B.n379 585
R276 B.n377 B.n139 585
R277 B.n375 B.n374 585
R278 B.n373 B.n140 585
R279 B.n372 B.n371 585
R280 B.n369 B.n141 585
R281 B.n367 B.n366 585
R282 B.n365 B.n142 585
R283 B.n364 B.n363 585
R284 B.n361 B.n143 585
R285 B.n359 B.n358 585
R286 B.n357 B.n144 585
R287 B.n356 B.n355 585
R288 B.n353 B.n145 585
R289 B.n351 B.n350 585
R290 B.n349 B.n146 585
R291 B.n348 B.n347 585
R292 B.n345 B.n147 585
R293 B.n343 B.n342 585
R294 B.n341 B.n148 585
R295 B.n340 B.n339 585
R296 B.n337 B.n149 585
R297 B.n335 B.n334 585
R298 B.n333 B.n150 585
R299 B.n332 B.n331 585
R300 B.n329 B.n151 585
R301 B.n327 B.n326 585
R302 B.n324 B.n152 585
R303 B.n323 B.n322 585
R304 B.n320 B.n155 585
R305 B.n318 B.n317 585
R306 B.n316 B.n156 585
R307 B.n315 B.n314 585
R308 B.n312 B.n157 585
R309 B.n310 B.n309 585
R310 B.n308 B.n158 585
R311 B.n306 B.n305 585
R312 B.n303 B.n161 585
R313 B.n301 B.n300 585
R314 B.n299 B.n162 585
R315 B.n298 B.n297 585
R316 B.n295 B.n163 585
R317 B.n293 B.n292 585
R318 B.n291 B.n164 585
R319 B.n290 B.n289 585
R320 B.n287 B.n165 585
R321 B.n285 B.n284 585
R322 B.n283 B.n166 585
R323 B.n282 B.n281 585
R324 B.n279 B.n167 585
R325 B.n277 B.n276 585
R326 B.n275 B.n168 585
R327 B.n274 B.n273 585
R328 B.n271 B.n169 585
R329 B.n269 B.n268 585
R330 B.n267 B.n170 585
R331 B.n266 B.n265 585
R332 B.n263 B.n171 585
R333 B.n261 B.n260 585
R334 B.n259 B.n172 585
R335 B.n258 B.n257 585
R336 B.n255 B.n173 585
R337 B.n253 B.n252 585
R338 B.n251 B.n174 585
R339 B.n250 B.n249 585
R340 B.n247 B.n175 585
R341 B.n245 B.n244 585
R342 B.n243 B.n176 585
R343 B.n242 B.n241 585
R344 B.n239 B.n177 585
R345 B.n237 B.n236 585
R346 B.n235 B.n178 585
R347 B.n234 B.n233 585
R348 B.n231 B.n179 585
R349 B.n229 B.n228 585
R350 B.n227 B.n180 585
R351 B.n226 B.n225 585
R352 B.n223 B.n181 585
R353 B.n221 B.n220 585
R354 B.n219 B.n182 585
R355 B.n218 B.n217 585
R356 B.n215 B.n183 585
R357 B.n213 B.n212 585
R358 B.n211 B.n184 585
R359 B.n210 B.n209 585
R360 B.n207 B.n185 585
R361 B.n205 B.n204 585
R362 B.n203 B.n186 585
R363 B.n202 B.n201 585
R364 B.n199 B.n187 585
R365 B.n197 B.n196 585
R366 B.n195 B.n188 585
R367 B.n194 B.n193 585
R368 B.n191 B.n189 585
R369 B.n120 B.n119 585
R370 B.n444 B.n443 585
R371 B.n445 B.n444 585
R372 B.n116 B.n115 585
R373 B.n117 B.n116 585
R374 B.n454 B.n453 585
R375 B.n453 B.n452 585
R376 B.n455 B.n114 585
R377 B.n451 B.n114 585
R378 B.n457 B.n456 585
R379 B.n458 B.n457 585
R380 B.n109 B.n108 585
R381 B.n110 B.n109 585
R382 B.n466 B.n465 585
R383 B.n465 B.n464 585
R384 B.n467 B.n107 585
R385 B.n107 B.n106 585
R386 B.n469 B.n468 585
R387 B.n470 B.n469 585
R388 B.n101 B.n100 585
R389 B.n102 B.n101 585
R390 B.n480 B.n479 585
R391 B.n479 B.n478 585
R392 B.n481 B.n99 585
R393 B.n477 B.n99 585
R394 B.n483 B.n482 585
R395 B.n484 B.n483 585
R396 B.n2 B.n0 585
R397 B.n4 B.n2 585
R398 B.n3 B.n1 585
R399 B.n789 B.n3 585
R400 B.n787 B.n786 585
R401 B.n788 B.n787 585
R402 B.n785 B.n8 585
R403 B.n491 B.n8 585
R404 B.n784 B.n783 585
R405 B.n783 B.n782 585
R406 B.n10 B.n9 585
R407 B.n781 B.n10 585
R408 B.n779 B.n778 585
R409 B.n780 B.n779 585
R410 B.n777 B.n15 585
R411 B.n15 B.n14 585
R412 B.n776 B.n775 585
R413 B.n775 B.n774 585
R414 B.n17 B.n16 585
R415 B.n773 B.n17 585
R416 B.n771 B.n770 585
R417 B.n772 B.n771 585
R418 B.n769 B.n21 585
R419 B.n24 B.n21 585
R420 B.n768 B.n767 585
R421 B.n767 B.n766 585
R422 B.n23 B.n22 585
R423 B.n765 B.n23 585
R424 B.n763 B.n762 585
R425 B.n764 B.n763 585
R426 B.n792 B.n791 585
R427 B.n791 B.n790 585
R428 B.n444 B.n122 511.721
R429 B.n763 B.n29 511.721
R430 B.n446 B.n120 511.721
R431 B.n508 B.n27 511.721
R432 B.n509 B.n28 256.663
R433 B.n515 B.n28 256.663
R434 B.n517 B.n28 256.663
R435 B.n523 B.n28 256.663
R436 B.n525 B.n28 256.663
R437 B.n531 B.n28 256.663
R438 B.n533 B.n28 256.663
R439 B.n539 B.n28 256.663
R440 B.n541 B.n28 256.663
R441 B.n547 B.n28 256.663
R442 B.n549 B.n28 256.663
R443 B.n555 B.n28 256.663
R444 B.n557 B.n28 256.663
R445 B.n563 B.n28 256.663
R446 B.n565 B.n28 256.663
R447 B.n571 B.n28 256.663
R448 B.n573 B.n28 256.663
R449 B.n579 B.n28 256.663
R450 B.n581 B.n28 256.663
R451 B.n587 B.n28 256.663
R452 B.n589 B.n28 256.663
R453 B.n595 B.n28 256.663
R454 B.n597 B.n28 256.663
R455 B.n603 B.n28 256.663
R456 B.n605 B.n28 256.663
R457 B.n611 B.n28 256.663
R458 B.n613 B.n28 256.663
R459 B.n619 B.n28 256.663
R460 B.n621 B.n28 256.663
R461 B.n628 B.n28 256.663
R462 B.n630 B.n28 256.663
R463 B.n636 B.n28 256.663
R464 B.n638 B.n28 256.663
R465 B.n644 B.n28 256.663
R466 B.n646 B.n28 256.663
R467 B.n652 B.n28 256.663
R468 B.n654 B.n28 256.663
R469 B.n660 B.n28 256.663
R470 B.n662 B.n28 256.663
R471 B.n668 B.n28 256.663
R472 B.n670 B.n28 256.663
R473 B.n676 B.n28 256.663
R474 B.n678 B.n28 256.663
R475 B.n684 B.n28 256.663
R476 B.n686 B.n28 256.663
R477 B.n692 B.n28 256.663
R478 B.n694 B.n28 256.663
R479 B.n700 B.n28 256.663
R480 B.n702 B.n28 256.663
R481 B.n708 B.n28 256.663
R482 B.n710 B.n28 256.663
R483 B.n716 B.n28 256.663
R484 B.n718 B.n28 256.663
R485 B.n724 B.n28 256.663
R486 B.n726 B.n28 256.663
R487 B.n732 B.n28 256.663
R488 B.n734 B.n28 256.663
R489 B.n740 B.n28 256.663
R490 B.n742 B.n28 256.663
R491 B.n748 B.n28 256.663
R492 B.n750 B.n28 256.663
R493 B.n756 B.n28 256.663
R494 B.n758 B.n28 256.663
R495 B.n439 B.n121 256.663
R496 B.n124 B.n121 256.663
R497 B.n432 B.n121 256.663
R498 B.n426 B.n121 256.663
R499 B.n424 B.n121 256.663
R500 B.n418 B.n121 256.663
R501 B.n416 B.n121 256.663
R502 B.n410 B.n121 256.663
R503 B.n408 B.n121 256.663
R504 B.n402 B.n121 256.663
R505 B.n400 B.n121 256.663
R506 B.n394 B.n121 256.663
R507 B.n392 B.n121 256.663
R508 B.n386 B.n121 256.663
R509 B.n384 B.n121 256.663
R510 B.n378 B.n121 256.663
R511 B.n376 B.n121 256.663
R512 B.n370 B.n121 256.663
R513 B.n368 B.n121 256.663
R514 B.n362 B.n121 256.663
R515 B.n360 B.n121 256.663
R516 B.n354 B.n121 256.663
R517 B.n352 B.n121 256.663
R518 B.n346 B.n121 256.663
R519 B.n344 B.n121 256.663
R520 B.n338 B.n121 256.663
R521 B.n336 B.n121 256.663
R522 B.n330 B.n121 256.663
R523 B.n328 B.n121 256.663
R524 B.n321 B.n121 256.663
R525 B.n319 B.n121 256.663
R526 B.n313 B.n121 256.663
R527 B.n311 B.n121 256.663
R528 B.n304 B.n121 256.663
R529 B.n302 B.n121 256.663
R530 B.n296 B.n121 256.663
R531 B.n294 B.n121 256.663
R532 B.n288 B.n121 256.663
R533 B.n286 B.n121 256.663
R534 B.n280 B.n121 256.663
R535 B.n278 B.n121 256.663
R536 B.n272 B.n121 256.663
R537 B.n270 B.n121 256.663
R538 B.n264 B.n121 256.663
R539 B.n262 B.n121 256.663
R540 B.n256 B.n121 256.663
R541 B.n254 B.n121 256.663
R542 B.n248 B.n121 256.663
R543 B.n246 B.n121 256.663
R544 B.n240 B.n121 256.663
R545 B.n238 B.n121 256.663
R546 B.n232 B.n121 256.663
R547 B.n230 B.n121 256.663
R548 B.n224 B.n121 256.663
R549 B.n222 B.n121 256.663
R550 B.n216 B.n121 256.663
R551 B.n214 B.n121 256.663
R552 B.n208 B.n121 256.663
R553 B.n206 B.n121 256.663
R554 B.n200 B.n121 256.663
R555 B.n198 B.n121 256.663
R556 B.n192 B.n121 256.663
R557 B.n190 B.n121 256.663
R558 B.n444 B.n116 163.367
R559 B.n453 B.n116 163.367
R560 B.n453 B.n114 163.367
R561 B.n457 B.n114 163.367
R562 B.n457 B.n109 163.367
R563 B.n465 B.n109 163.367
R564 B.n465 B.n107 163.367
R565 B.n469 B.n107 163.367
R566 B.n469 B.n101 163.367
R567 B.n479 B.n101 163.367
R568 B.n479 B.n99 163.367
R569 B.n483 B.n99 163.367
R570 B.n483 B.n2 163.367
R571 B.n791 B.n2 163.367
R572 B.n791 B.n3 163.367
R573 B.n787 B.n3 163.367
R574 B.n787 B.n8 163.367
R575 B.n783 B.n8 163.367
R576 B.n783 B.n10 163.367
R577 B.n779 B.n10 163.367
R578 B.n779 B.n15 163.367
R579 B.n775 B.n15 163.367
R580 B.n775 B.n17 163.367
R581 B.n771 B.n17 163.367
R582 B.n771 B.n21 163.367
R583 B.n767 B.n21 163.367
R584 B.n767 B.n23 163.367
R585 B.n763 B.n23 163.367
R586 B.n440 B.n438 163.367
R587 B.n438 B.n437 163.367
R588 B.n434 B.n433 163.367
R589 B.n431 B.n126 163.367
R590 B.n427 B.n425 163.367
R591 B.n423 B.n128 163.367
R592 B.n419 B.n417 163.367
R593 B.n415 B.n130 163.367
R594 B.n411 B.n409 163.367
R595 B.n407 B.n132 163.367
R596 B.n403 B.n401 163.367
R597 B.n399 B.n134 163.367
R598 B.n395 B.n393 163.367
R599 B.n391 B.n136 163.367
R600 B.n387 B.n385 163.367
R601 B.n383 B.n138 163.367
R602 B.n379 B.n377 163.367
R603 B.n375 B.n140 163.367
R604 B.n371 B.n369 163.367
R605 B.n367 B.n142 163.367
R606 B.n363 B.n361 163.367
R607 B.n359 B.n144 163.367
R608 B.n355 B.n353 163.367
R609 B.n351 B.n146 163.367
R610 B.n347 B.n345 163.367
R611 B.n343 B.n148 163.367
R612 B.n339 B.n337 163.367
R613 B.n335 B.n150 163.367
R614 B.n331 B.n329 163.367
R615 B.n327 B.n152 163.367
R616 B.n322 B.n320 163.367
R617 B.n318 B.n156 163.367
R618 B.n314 B.n312 163.367
R619 B.n310 B.n158 163.367
R620 B.n305 B.n303 163.367
R621 B.n301 B.n162 163.367
R622 B.n297 B.n295 163.367
R623 B.n293 B.n164 163.367
R624 B.n289 B.n287 163.367
R625 B.n285 B.n166 163.367
R626 B.n281 B.n279 163.367
R627 B.n277 B.n168 163.367
R628 B.n273 B.n271 163.367
R629 B.n269 B.n170 163.367
R630 B.n265 B.n263 163.367
R631 B.n261 B.n172 163.367
R632 B.n257 B.n255 163.367
R633 B.n253 B.n174 163.367
R634 B.n249 B.n247 163.367
R635 B.n245 B.n176 163.367
R636 B.n241 B.n239 163.367
R637 B.n237 B.n178 163.367
R638 B.n233 B.n231 163.367
R639 B.n229 B.n180 163.367
R640 B.n225 B.n223 163.367
R641 B.n221 B.n182 163.367
R642 B.n217 B.n215 163.367
R643 B.n213 B.n184 163.367
R644 B.n209 B.n207 163.367
R645 B.n205 B.n186 163.367
R646 B.n201 B.n199 163.367
R647 B.n197 B.n188 163.367
R648 B.n193 B.n191 163.367
R649 B.n446 B.n118 163.367
R650 B.n450 B.n118 163.367
R651 B.n450 B.n113 163.367
R652 B.n459 B.n113 163.367
R653 B.n459 B.n111 163.367
R654 B.n463 B.n111 163.367
R655 B.n463 B.n105 163.367
R656 B.n471 B.n105 163.367
R657 B.n471 B.n103 163.367
R658 B.n476 B.n103 163.367
R659 B.n476 B.n98 163.367
R660 B.n485 B.n98 163.367
R661 B.n486 B.n485 163.367
R662 B.n486 B.n5 163.367
R663 B.n6 B.n5 163.367
R664 B.n7 B.n6 163.367
R665 B.n492 B.n7 163.367
R666 B.n492 B.n11 163.367
R667 B.n12 B.n11 163.367
R668 B.n13 B.n12 163.367
R669 B.n497 B.n13 163.367
R670 B.n497 B.n18 163.367
R671 B.n19 B.n18 163.367
R672 B.n20 B.n19 163.367
R673 B.n502 B.n20 163.367
R674 B.n502 B.n25 163.367
R675 B.n26 B.n25 163.367
R676 B.n27 B.n26 163.367
R677 B.n759 B.n757 163.367
R678 B.n755 B.n31 163.367
R679 B.n751 B.n749 163.367
R680 B.n747 B.n33 163.367
R681 B.n743 B.n741 163.367
R682 B.n739 B.n35 163.367
R683 B.n735 B.n733 163.367
R684 B.n731 B.n37 163.367
R685 B.n727 B.n725 163.367
R686 B.n723 B.n39 163.367
R687 B.n719 B.n717 163.367
R688 B.n715 B.n41 163.367
R689 B.n711 B.n709 163.367
R690 B.n707 B.n43 163.367
R691 B.n703 B.n701 163.367
R692 B.n699 B.n45 163.367
R693 B.n695 B.n693 163.367
R694 B.n691 B.n47 163.367
R695 B.n687 B.n685 163.367
R696 B.n683 B.n49 163.367
R697 B.n679 B.n677 163.367
R698 B.n675 B.n51 163.367
R699 B.n671 B.n669 163.367
R700 B.n667 B.n53 163.367
R701 B.n663 B.n661 163.367
R702 B.n659 B.n55 163.367
R703 B.n655 B.n653 163.367
R704 B.n651 B.n57 163.367
R705 B.n647 B.n645 163.367
R706 B.n643 B.n59 163.367
R707 B.n639 B.n637 163.367
R708 B.n635 B.n64 163.367
R709 B.n631 B.n629 163.367
R710 B.n627 B.n66 163.367
R711 B.n622 B.n620 163.367
R712 B.n618 B.n70 163.367
R713 B.n614 B.n612 163.367
R714 B.n610 B.n72 163.367
R715 B.n606 B.n604 163.367
R716 B.n602 B.n74 163.367
R717 B.n598 B.n596 163.367
R718 B.n594 B.n76 163.367
R719 B.n590 B.n588 163.367
R720 B.n586 B.n78 163.367
R721 B.n582 B.n580 163.367
R722 B.n578 B.n80 163.367
R723 B.n574 B.n572 163.367
R724 B.n570 B.n82 163.367
R725 B.n566 B.n564 163.367
R726 B.n562 B.n84 163.367
R727 B.n558 B.n556 163.367
R728 B.n554 B.n86 163.367
R729 B.n550 B.n548 163.367
R730 B.n546 B.n88 163.367
R731 B.n542 B.n540 163.367
R732 B.n538 B.n90 163.367
R733 B.n534 B.n532 163.367
R734 B.n530 B.n92 163.367
R735 B.n526 B.n524 163.367
R736 B.n522 B.n94 163.367
R737 B.n518 B.n516 163.367
R738 B.n514 B.n96 163.367
R739 B.n510 B.n508 163.367
R740 B.n159 B.t16 79.4789
R741 B.n67 B.t18 79.4789
R742 B.n153 B.t13 79.4552
R743 B.n60 B.t8 79.4552
R744 B.n439 B.n122 71.676
R745 B.n437 B.n124 71.676
R746 B.n433 B.n432 71.676
R747 B.n426 B.n126 71.676
R748 B.n425 B.n424 71.676
R749 B.n418 B.n128 71.676
R750 B.n417 B.n416 71.676
R751 B.n410 B.n130 71.676
R752 B.n409 B.n408 71.676
R753 B.n402 B.n132 71.676
R754 B.n401 B.n400 71.676
R755 B.n394 B.n134 71.676
R756 B.n393 B.n392 71.676
R757 B.n386 B.n136 71.676
R758 B.n385 B.n384 71.676
R759 B.n378 B.n138 71.676
R760 B.n377 B.n376 71.676
R761 B.n370 B.n140 71.676
R762 B.n369 B.n368 71.676
R763 B.n362 B.n142 71.676
R764 B.n361 B.n360 71.676
R765 B.n354 B.n144 71.676
R766 B.n353 B.n352 71.676
R767 B.n346 B.n146 71.676
R768 B.n345 B.n344 71.676
R769 B.n338 B.n148 71.676
R770 B.n337 B.n336 71.676
R771 B.n330 B.n150 71.676
R772 B.n329 B.n328 71.676
R773 B.n321 B.n152 71.676
R774 B.n320 B.n319 71.676
R775 B.n313 B.n156 71.676
R776 B.n312 B.n311 71.676
R777 B.n304 B.n158 71.676
R778 B.n303 B.n302 71.676
R779 B.n296 B.n162 71.676
R780 B.n295 B.n294 71.676
R781 B.n288 B.n164 71.676
R782 B.n287 B.n286 71.676
R783 B.n280 B.n166 71.676
R784 B.n279 B.n278 71.676
R785 B.n272 B.n168 71.676
R786 B.n271 B.n270 71.676
R787 B.n264 B.n170 71.676
R788 B.n263 B.n262 71.676
R789 B.n256 B.n172 71.676
R790 B.n255 B.n254 71.676
R791 B.n248 B.n174 71.676
R792 B.n247 B.n246 71.676
R793 B.n240 B.n176 71.676
R794 B.n239 B.n238 71.676
R795 B.n232 B.n178 71.676
R796 B.n231 B.n230 71.676
R797 B.n224 B.n180 71.676
R798 B.n223 B.n222 71.676
R799 B.n216 B.n182 71.676
R800 B.n215 B.n214 71.676
R801 B.n208 B.n184 71.676
R802 B.n207 B.n206 71.676
R803 B.n200 B.n186 71.676
R804 B.n199 B.n198 71.676
R805 B.n192 B.n188 71.676
R806 B.n191 B.n190 71.676
R807 B.n758 B.n29 71.676
R808 B.n757 B.n756 71.676
R809 B.n750 B.n31 71.676
R810 B.n749 B.n748 71.676
R811 B.n742 B.n33 71.676
R812 B.n741 B.n740 71.676
R813 B.n734 B.n35 71.676
R814 B.n733 B.n732 71.676
R815 B.n726 B.n37 71.676
R816 B.n725 B.n724 71.676
R817 B.n718 B.n39 71.676
R818 B.n717 B.n716 71.676
R819 B.n710 B.n41 71.676
R820 B.n709 B.n708 71.676
R821 B.n702 B.n43 71.676
R822 B.n701 B.n700 71.676
R823 B.n694 B.n45 71.676
R824 B.n693 B.n692 71.676
R825 B.n686 B.n47 71.676
R826 B.n685 B.n684 71.676
R827 B.n678 B.n49 71.676
R828 B.n677 B.n676 71.676
R829 B.n670 B.n51 71.676
R830 B.n669 B.n668 71.676
R831 B.n662 B.n53 71.676
R832 B.n661 B.n660 71.676
R833 B.n654 B.n55 71.676
R834 B.n653 B.n652 71.676
R835 B.n646 B.n57 71.676
R836 B.n645 B.n644 71.676
R837 B.n638 B.n59 71.676
R838 B.n637 B.n636 71.676
R839 B.n630 B.n64 71.676
R840 B.n629 B.n628 71.676
R841 B.n621 B.n66 71.676
R842 B.n620 B.n619 71.676
R843 B.n613 B.n70 71.676
R844 B.n612 B.n611 71.676
R845 B.n605 B.n72 71.676
R846 B.n604 B.n603 71.676
R847 B.n597 B.n74 71.676
R848 B.n596 B.n595 71.676
R849 B.n589 B.n76 71.676
R850 B.n588 B.n587 71.676
R851 B.n581 B.n78 71.676
R852 B.n580 B.n579 71.676
R853 B.n573 B.n80 71.676
R854 B.n572 B.n571 71.676
R855 B.n565 B.n82 71.676
R856 B.n564 B.n563 71.676
R857 B.n557 B.n84 71.676
R858 B.n556 B.n555 71.676
R859 B.n549 B.n86 71.676
R860 B.n548 B.n547 71.676
R861 B.n541 B.n88 71.676
R862 B.n540 B.n539 71.676
R863 B.n533 B.n90 71.676
R864 B.n532 B.n531 71.676
R865 B.n525 B.n92 71.676
R866 B.n524 B.n523 71.676
R867 B.n517 B.n94 71.676
R868 B.n516 B.n515 71.676
R869 B.n509 B.n96 71.676
R870 B.n510 B.n509 71.676
R871 B.n515 B.n514 71.676
R872 B.n518 B.n517 71.676
R873 B.n523 B.n522 71.676
R874 B.n526 B.n525 71.676
R875 B.n531 B.n530 71.676
R876 B.n534 B.n533 71.676
R877 B.n539 B.n538 71.676
R878 B.n542 B.n541 71.676
R879 B.n547 B.n546 71.676
R880 B.n550 B.n549 71.676
R881 B.n555 B.n554 71.676
R882 B.n558 B.n557 71.676
R883 B.n563 B.n562 71.676
R884 B.n566 B.n565 71.676
R885 B.n571 B.n570 71.676
R886 B.n574 B.n573 71.676
R887 B.n579 B.n578 71.676
R888 B.n582 B.n581 71.676
R889 B.n587 B.n586 71.676
R890 B.n590 B.n589 71.676
R891 B.n595 B.n594 71.676
R892 B.n598 B.n597 71.676
R893 B.n603 B.n602 71.676
R894 B.n606 B.n605 71.676
R895 B.n611 B.n610 71.676
R896 B.n614 B.n613 71.676
R897 B.n619 B.n618 71.676
R898 B.n622 B.n621 71.676
R899 B.n628 B.n627 71.676
R900 B.n631 B.n630 71.676
R901 B.n636 B.n635 71.676
R902 B.n639 B.n638 71.676
R903 B.n644 B.n643 71.676
R904 B.n647 B.n646 71.676
R905 B.n652 B.n651 71.676
R906 B.n655 B.n654 71.676
R907 B.n660 B.n659 71.676
R908 B.n663 B.n662 71.676
R909 B.n668 B.n667 71.676
R910 B.n671 B.n670 71.676
R911 B.n676 B.n675 71.676
R912 B.n679 B.n678 71.676
R913 B.n684 B.n683 71.676
R914 B.n687 B.n686 71.676
R915 B.n692 B.n691 71.676
R916 B.n695 B.n694 71.676
R917 B.n700 B.n699 71.676
R918 B.n703 B.n702 71.676
R919 B.n708 B.n707 71.676
R920 B.n711 B.n710 71.676
R921 B.n716 B.n715 71.676
R922 B.n719 B.n718 71.676
R923 B.n724 B.n723 71.676
R924 B.n727 B.n726 71.676
R925 B.n732 B.n731 71.676
R926 B.n735 B.n734 71.676
R927 B.n740 B.n739 71.676
R928 B.n743 B.n742 71.676
R929 B.n748 B.n747 71.676
R930 B.n751 B.n750 71.676
R931 B.n756 B.n755 71.676
R932 B.n759 B.n758 71.676
R933 B.n440 B.n439 71.676
R934 B.n434 B.n124 71.676
R935 B.n432 B.n431 71.676
R936 B.n427 B.n426 71.676
R937 B.n424 B.n423 71.676
R938 B.n419 B.n418 71.676
R939 B.n416 B.n415 71.676
R940 B.n411 B.n410 71.676
R941 B.n408 B.n407 71.676
R942 B.n403 B.n402 71.676
R943 B.n400 B.n399 71.676
R944 B.n395 B.n394 71.676
R945 B.n392 B.n391 71.676
R946 B.n387 B.n386 71.676
R947 B.n384 B.n383 71.676
R948 B.n379 B.n378 71.676
R949 B.n376 B.n375 71.676
R950 B.n371 B.n370 71.676
R951 B.n368 B.n367 71.676
R952 B.n363 B.n362 71.676
R953 B.n360 B.n359 71.676
R954 B.n355 B.n354 71.676
R955 B.n352 B.n351 71.676
R956 B.n347 B.n346 71.676
R957 B.n344 B.n343 71.676
R958 B.n339 B.n338 71.676
R959 B.n336 B.n335 71.676
R960 B.n331 B.n330 71.676
R961 B.n328 B.n327 71.676
R962 B.n322 B.n321 71.676
R963 B.n319 B.n318 71.676
R964 B.n314 B.n313 71.676
R965 B.n311 B.n310 71.676
R966 B.n305 B.n304 71.676
R967 B.n302 B.n301 71.676
R968 B.n297 B.n296 71.676
R969 B.n294 B.n293 71.676
R970 B.n289 B.n288 71.676
R971 B.n286 B.n285 71.676
R972 B.n281 B.n280 71.676
R973 B.n278 B.n277 71.676
R974 B.n273 B.n272 71.676
R975 B.n270 B.n269 71.676
R976 B.n265 B.n264 71.676
R977 B.n262 B.n261 71.676
R978 B.n257 B.n256 71.676
R979 B.n254 B.n253 71.676
R980 B.n249 B.n248 71.676
R981 B.n246 B.n245 71.676
R982 B.n241 B.n240 71.676
R983 B.n238 B.n237 71.676
R984 B.n233 B.n232 71.676
R985 B.n230 B.n229 71.676
R986 B.n225 B.n224 71.676
R987 B.n222 B.n221 71.676
R988 B.n217 B.n216 71.676
R989 B.n214 B.n213 71.676
R990 B.n209 B.n208 71.676
R991 B.n206 B.n205 71.676
R992 B.n201 B.n200 71.676
R993 B.n198 B.n197 71.676
R994 B.n193 B.n192 71.676
R995 B.n190 B.n120 71.676
R996 B.n160 B.t15 69.588
R997 B.n68 B.t19 69.588
R998 B.n154 B.t12 69.5643
R999 B.n61 B.t9 69.5643
R1000 B.n445 B.n121 62.449
R1001 B.n764 B.n28 62.449
R1002 B.n307 B.n160 59.5399
R1003 B.n325 B.n154 59.5399
R1004 B.n62 B.n61 59.5399
R1005 B.n625 B.n68 59.5399
R1006 B.n762 B.n761 33.2493
R1007 B.n507 B.n506 33.2493
R1008 B.n447 B.n119 33.2493
R1009 B.n443 B.n442 33.2493
R1010 B.n445 B.n117 32.4165
R1011 B.n452 B.n117 32.4165
R1012 B.n452 B.n451 32.4165
R1013 B.n458 B.n110 32.4165
R1014 B.n464 B.n110 32.4165
R1015 B.n464 B.n106 32.4165
R1016 B.n470 B.n106 32.4165
R1017 B.n478 B.n102 32.4165
R1018 B.n484 B.n4 32.4165
R1019 B.n790 B.n4 32.4165
R1020 B.n790 B.n789 32.4165
R1021 B.n789 B.n788 32.4165
R1022 B.n782 B.n781 32.4165
R1023 B.n780 B.n14 32.4165
R1024 B.n774 B.n14 32.4165
R1025 B.n774 B.n773 32.4165
R1026 B.n773 B.n772 32.4165
R1027 B.n766 B.n24 32.4165
R1028 B.n766 B.n765 32.4165
R1029 B.n765 B.n764 32.4165
R1030 B.n451 B.t11 30.5097
R1031 B.n24 B.t7 30.5097
R1032 B.t4 B.n477 27.6495
R1033 B.n491 B.t2 27.6495
R1034 B.n470 B.t5 20.9756
R1035 B.n477 B.t3 20.9756
R1036 B.n491 B.t0 20.9756
R1037 B.t1 B.n780 20.9756
R1038 B B.n792 18.0485
R1039 B.t5 B.n102 11.4415
R1040 B.n484 B.t3 11.4415
R1041 B.n788 B.t0 11.4415
R1042 B.n781 B.t1 11.4415
R1043 B.n761 B.n760 10.6151
R1044 B.n760 B.n30 10.6151
R1045 B.n754 B.n30 10.6151
R1046 B.n754 B.n753 10.6151
R1047 B.n753 B.n752 10.6151
R1048 B.n752 B.n32 10.6151
R1049 B.n746 B.n32 10.6151
R1050 B.n746 B.n745 10.6151
R1051 B.n745 B.n744 10.6151
R1052 B.n744 B.n34 10.6151
R1053 B.n738 B.n34 10.6151
R1054 B.n738 B.n737 10.6151
R1055 B.n737 B.n736 10.6151
R1056 B.n736 B.n36 10.6151
R1057 B.n730 B.n36 10.6151
R1058 B.n730 B.n729 10.6151
R1059 B.n729 B.n728 10.6151
R1060 B.n728 B.n38 10.6151
R1061 B.n722 B.n38 10.6151
R1062 B.n722 B.n721 10.6151
R1063 B.n721 B.n720 10.6151
R1064 B.n720 B.n40 10.6151
R1065 B.n714 B.n40 10.6151
R1066 B.n714 B.n713 10.6151
R1067 B.n713 B.n712 10.6151
R1068 B.n712 B.n42 10.6151
R1069 B.n706 B.n42 10.6151
R1070 B.n706 B.n705 10.6151
R1071 B.n705 B.n704 10.6151
R1072 B.n704 B.n44 10.6151
R1073 B.n698 B.n44 10.6151
R1074 B.n698 B.n697 10.6151
R1075 B.n697 B.n696 10.6151
R1076 B.n696 B.n46 10.6151
R1077 B.n690 B.n46 10.6151
R1078 B.n690 B.n689 10.6151
R1079 B.n689 B.n688 10.6151
R1080 B.n688 B.n48 10.6151
R1081 B.n682 B.n48 10.6151
R1082 B.n682 B.n681 10.6151
R1083 B.n681 B.n680 10.6151
R1084 B.n680 B.n50 10.6151
R1085 B.n674 B.n50 10.6151
R1086 B.n674 B.n673 10.6151
R1087 B.n673 B.n672 10.6151
R1088 B.n672 B.n52 10.6151
R1089 B.n666 B.n52 10.6151
R1090 B.n666 B.n665 10.6151
R1091 B.n665 B.n664 10.6151
R1092 B.n664 B.n54 10.6151
R1093 B.n658 B.n54 10.6151
R1094 B.n658 B.n657 10.6151
R1095 B.n657 B.n656 10.6151
R1096 B.n656 B.n56 10.6151
R1097 B.n650 B.n56 10.6151
R1098 B.n650 B.n649 10.6151
R1099 B.n649 B.n648 10.6151
R1100 B.n648 B.n58 10.6151
R1101 B.n642 B.n641 10.6151
R1102 B.n641 B.n640 10.6151
R1103 B.n640 B.n63 10.6151
R1104 B.n634 B.n63 10.6151
R1105 B.n634 B.n633 10.6151
R1106 B.n633 B.n632 10.6151
R1107 B.n632 B.n65 10.6151
R1108 B.n626 B.n65 10.6151
R1109 B.n624 B.n623 10.6151
R1110 B.n623 B.n69 10.6151
R1111 B.n617 B.n69 10.6151
R1112 B.n617 B.n616 10.6151
R1113 B.n616 B.n615 10.6151
R1114 B.n615 B.n71 10.6151
R1115 B.n609 B.n71 10.6151
R1116 B.n609 B.n608 10.6151
R1117 B.n608 B.n607 10.6151
R1118 B.n607 B.n73 10.6151
R1119 B.n601 B.n73 10.6151
R1120 B.n601 B.n600 10.6151
R1121 B.n600 B.n599 10.6151
R1122 B.n599 B.n75 10.6151
R1123 B.n593 B.n75 10.6151
R1124 B.n593 B.n592 10.6151
R1125 B.n592 B.n591 10.6151
R1126 B.n591 B.n77 10.6151
R1127 B.n585 B.n77 10.6151
R1128 B.n585 B.n584 10.6151
R1129 B.n584 B.n583 10.6151
R1130 B.n583 B.n79 10.6151
R1131 B.n577 B.n79 10.6151
R1132 B.n577 B.n576 10.6151
R1133 B.n576 B.n575 10.6151
R1134 B.n575 B.n81 10.6151
R1135 B.n569 B.n81 10.6151
R1136 B.n569 B.n568 10.6151
R1137 B.n568 B.n567 10.6151
R1138 B.n567 B.n83 10.6151
R1139 B.n561 B.n83 10.6151
R1140 B.n561 B.n560 10.6151
R1141 B.n560 B.n559 10.6151
R1142 B.n559 B.n85 10.6151
R1143 B.n553 B.n85 10.6151
R1144 B.n553 B.n552 10.6151
R1145 B.n552 B.n551 10.6151
R1146 B.n551 B.n87 10.6151
R1147 B.n545 B.n87 10.6151
R1148 B.n545 B.n544 10.6151
R1149 B.n544 B.n543 10.6151
R1150 B.n543 B.n89 10.6151
R1151 B.n537 B.n89 10.6151
R1152 B.n537 B.n536 10.6151
R1153 B.n536 B.n535 10.6151
R1154 B.n535 B.n91 10.6151
R1155 B.n529 B.n91 10.6151
R1156 B.n529 B.n528 10.6151
R1157 B.n528 B.n527 10.6151
R1158 B.n527 B.n93 10.6151
R1159 B.n521 B.n93 10.6151
R1160 B.n521 B.n520 10.6151
R1161 B.n520 B.n519 10.6151
R1162 B.n519 B.n95 10.6151
R1163 B.n513 B.n95 10.6151
R1164 B.n513 B.n512 10.6151
R1165 B.n512 B.n511 10.6151
R1166 B.n511 B.n507 10.6151
R1167 B.n448 B.n447 10.6151
R1168 B.n449 B.n448 10.6151
R1169 B.n449 B.n112 10.6151
R1170 B.n460 B.n112 10.6151
R1171 B.n461 B.n460 10.6151
R1172 B.n462 B.n461 10.6151
R1173 B.n462 B.n104 10.6151
R1174 B.n472 B.n104 10.6151
R1175 B.n473 B.n472 10.6151
R1176 B.n475 B.n473 10.6151
R1177 B.n475 B.n474 10.6151
R1178 B.n474 B.n97 10.6151
R1179 B.n487 B.n97 10.6151
R1180 B.n488 B.n487 10.6151
R1181 B.n489 B.n488 10.6151
R1182 B.n490 B.n489 10.6151
R1183 B.n493 B.n490 10.6151
R1184 B.n494 B.n493 10.6151
R1185 B.n495 B.n494 10.6151
R1186 B.n496 B.n495 10.6151
R1187 B.n498 B.n496 10.6151
R1188 B.n499 B.n498 10.6151
R1189 B.n500 B.n499 10.6151
R1190 B.n501 B.n500 10.6151
R1191 B.n503 B.n501 10.6151
R1192 B.n504 B.n503 10.6151
R1193 B.n505 B.n504 10.6151
R1194 B.n506 B.n505 10.6151
R1195 B.n442 B.n441 10.6151
R1196 B.n441 B.n123 10.6151
R1197 B.n436 B.n123 10.6151
R1198 B.n436 B.n435 10.6151
R1199 B.n435 B.n125 10.6151
R1200 B.n430 B.n125 10.6151
R1201 B.n430 B.n429 10.6151
R1202 B.n429 B.n428 10.6151
R1203 B.n428 B.n127 10.6151
R1204 B.n422 B.n127 10.6151
R1205 B.n422 B.n421 10.6151
R1206 B.n421 B.n420 10.6151
R1207 B.n420 B.n129 10.6151
R1208 B.n414 B.n129 10.6151
R1209 B.n414 B.n413 10.6151
R1210 B.n413 B.n412 10.6151
R1211 B.n412 B.n131 10.6151
R1212 B.n406 B.n131 10.6151
R1213 B.n406 B.n405 10.6151
R1214 B.n405 B.n404 10.6151
R1215 B.n404 B.n133 10.6151
R1216 B.n398 B.n133 10.6151
R1217 B.n398 B.n397 10.6151
R1218 B.n397 B.n396 10.6151
R1219 B.n396 B.n135 10.6151
R1220 B.n390 B.n135 10.6151
R1221 B.n390 B.n389 10.6151
R1222 B.n389 B.n388 10.6151
R1223 B.n388 B.n137 10.6151
R1224 B.n382 B.n137 10.6151
R1225 B.n382 B.n381 10.6151
R1226 B.n381 B.n380 10.6151
R1227 B.n380 B.n139 10.6151
R1228 B.n374 B.n139 10.6151
R1229 B.n374 B.n373 10.6151
R1230 B.n373 B.n372 10.6151
R1231 B.n372 B.n141 10.6151
R1232 B.n366 B.n141 10.6151
R1233 B.n366 B.n365 10.6151
R1234 B.n365 B.n364 10.6151
R1235 B.n364 B.n143 10.6151
R1236 B.n358 B.n143 10.6151
R1237 B.n358 B.n357 10.6151
R1238 B.n357 B.n356 10.6151
R1239 B.n356 B.n145 10.6151
R1240 B.n350 B.n145 10.6151
R1241 B.n350 B.n349 10.6151
R1242 B.n349 B.n348 10.6151
R1243 B.n348 B.n147 10.6151
R1244 B.n342 B.n147 10.6151
R1245 B.n342 B.n341 10.6151
R1246 B.n341 B.n340 10.6151
R1247 B.n340 B.n149 10.6151
R1248 B.n334 B.n149 10.6151
R1249 B.n334 B.n333 10.6151
R1250 B.n333 B.n332 10.6151
R1251 B.n332 B.n151 10.6151
R1252 B.n326 B.n151 10.6151
R1253 B.n324 B.n323 10.6151
R1254 B.n323 B.n155 10.6151
R1255 B.n317 B.n155 10.6151
R1256 B.n317 B.n316 10.6151
R1257 B.n316 B.n315 10.6151
R1258 B.n315 B.n157 10.6151
R1259 B.n309 B.n157 10.6151
R1260 B.n309 B.n308 10.6151
R1261 B.n306 B.n161 10.6151
R1262 B.n300 B.n161 10.6151
R1263 B.n300 B.n299 10.6151
R1264 B.n299 B.n298 10.6151
R1265 B.n298 B.n163 10.6151
R1266 B.n292 B.n163 10.6151
R1267 B.n292 B.n291 10.6151
R1268 B.n291 B.n290 10.6151
R1269 B.n290 B.n165 10.6151
R1270 B.n284 B.n165 10.6151
R1271 B.n284 B.n283 10.6151
R1272 B.n283 B.n282 10.6151
R1273 B.n282 B.n167 10.6151
R1274 B.n276 B.n167 10.6151
R1275 B.n276 B.n275 10.6151
R1276 B.n275 B.n274 10.6151
R1277 B.n274 B.n169 10.6151
R1278 B.n268 B.n169 10.6151
R1279 B.n268 B.n267 10.6151
R1280 B.n267 B.n266 10.6151
R1281 B.n266 B.n171 10.6151
R1282 B.n260 B.n171 10.6151
R1283 B.n260 B.n259 10.6151
R1284 B.n259 B.n258 10.6151
R1285 B.n258 B.n173 10.6151
R1286 B.n252 B.n173 10.6151
R1287 B.n252 B.n251 10.6151
R1288 B.n251 B.n250 10.6151
R1289 B.n250 B.n175 10.6151
R1290 B.n244 B.n175 10.6151
R1291 B.n244 B.n243 10.6151
R1292 B.n243 B.n242 10.6151
R1293 B.n242 B.n177 10.6151
R1294 B.n236 B.n177 10.6151
R1295 B.n236 B.n235 10.6151
R1296 B.n235 B.n234 10.6151
R1297 B.n234 B.n179 10.6151
R1298 B.n228 B.n179 10.6151
R1299 B.n228 B.n227 10.6151
R1300 B.n227 B.n226 10.6151
R1301 B.n226 B.n181 10.6151
R1302 B.n220 B.n181 10.6151
R1303 B.n220 B.n219 10.6151
R1304 B.n219 B.n218 10.6151
R1305 B.n218 B.n183 10.6151
R1306 B.n212 B.n183 10.6151
R1307 B.n212 B.n211 10.6151
R1308 B.n211 B.n210 10.6151
R1309 B.n210 B.n185 10.6151
R1310 B.n204 B.n185 10.6151
R1311 B.n204 B.n203 10.6151
R1312 B.n203 B.n202 10.6151
R1313 B.n202 B.n187 10.6151
R1314 B.n196 B.n187 10.6151
R1315 B.n196 B.n195 10.6151
R1316 B.n195 B.n194 10.6151
R1317 B.n194 B.n189 10.6151
R1318 B.n189 B.n119 10.6151
R1319 B.n443 B.n115 10.6151
R1320 B.n454 B.n115 10.6151
R1321 B.n455 B.n454 10.6151
R1322 B.n456 B.n455 10.6151
R1323 B.n456 B.n108 10.6151
R1324 B.n466 B.n108 10.6151
R1325 B.n467 B.n466 10.6151
R1326 B.n468 B.n467 10.6151
R1327 B.n468 B.n100 10.6151
R1328 B.n480 B.n100 10.6151
R1329 B.n481 B.n480 10.6151
R1330 B.n482 B.n481 10.6151
R1331 B.n482 B.n0 10.6151
R1332 B.n786 B.n1 10.6151
R1333 B.n786 B.n785 10.6151
R1334 B.n785 B.n784 10.6151
R1335 B.n784 B.n9 10.6151
R1336 B.n778 B.n9 10.6151
R1337 B.n778 B.n777 10.6151
R1338 B.n777 B.n776 10.6151
R1339 B.n776 B.n16 10.6151
R1340 B.n770 B.n16 10.6151
R1341 B.n770 B.n769 10.6151
R1342 B.n769 B.n768 10.6151
R1343 B.n768 B.n22 10.6151
R1344 B.n762 B.n22 10.6151
R1345 B.n160 B.n159 9.89141
R1346 B.n154 B.n153 9.89141
R1347 B.n61 B.n60 9.89141
R1348 B.n68 B.n67 9.89141
R1349 B.n642 B.n62 6.5566
R1350 B.n626 B.n625 6.5566
R1351 B.n325 B.n324 6.5566
R1352 B.n308 B.n307 6.5566
R1353 B.n478 B.t4 4.76756
R1354 B.n782 B.t2 4.76756
R1355 B.n62 B.n58 4.05904
R1356 B.n625 B.n624 4.05904
R1357 B.n326 B.n325 4.05904
R1358 B.n307 B.n306 4.05904
R1359 B.n792 B.n0 2.81026
R1360 B.n792 B.n1 2.81026
R1361 B.n458 B.t11 1.90733
R1362 B.n772 B.t7 1.90733
R1363 VN.n2 VN.t2 2595.25
R1364 VN.n0 VN.t0 2595.25
R1365 VN.n6 VN.t5 2595.25
R1366 VN.n4 VN.t3 2595.25
R1367 VN.n1 VN.t1 2557.28
R1368 VN.n5 VN.t4 2557.28
R1369 VN.n7 VN.n4 161.489
R1370 VN.n3 VN.n0 161.489
R1371 VN.n3 VN.n2 161.3
R1372 VN.n7 VN.n6 161.3
R1373 VN VN.n7 43.9835
R1374 VN.n1 VN.n0 36.5157
R1375 VN.n2 VN.n1 36.5157
R1376 VN.n6 VN.n5 36.5157
R1377 VN.n5 VN.n4 36.5157
R1378 VN VN.n3 0.0516364
R1379 VDD2.n1 VDD2.t5 60.499
R1380 VDD2.n2 VDD2.t0 60.2248
R1381 VDD2.n1 VDD2.n0 59.1668
R1382 VDD2 VDD2.n3 59.164
R1383 VDD2.n2 VDD2.n1 40.489
R1384 VDD2.n3 VDD2.t1 1.11286
R1385 VDD2.n3 VDD2.t2 1.11286
R1386 VDD2.n0 VDD2.t4 1.11286
R1387 VDD2.n0 VDD2.t3 1.11286
R1388 VDD2 VDD2.n2 0.388431
C0 VDD1 VP 2.98254f
C1 VDD2 VP 0.255051f
C2 VDD2 VDD1 0.53124f
C3 VN VTAIL 2.08425f
C4 VP VN 5.64926f
C5 VP VTAIL 2.09941f
C6 VDD1 VN 0.147524f
C7 VDD2 VN 2.88288f
C8 VDD1 VTAIL 24.2706f
C9 VDD2 VTAIL 24.2941f
C10 VDD2 B 5.181761f
C11 VDD1 B 5.400463f
C12 VTAIL B 7.955803f
C13 VN B 7.47441f
C14 VP B 4.59224f
C15 VDD2.t5 B 5.27223f
C16 VDD2.t4 B 0.453311f
C17 VDD2.t3 B 0.453311f
C18 VDD2.n0 B 4.12506f
C19 VDD2.n1 B 2.87095f
C20 VDD2.t0 B 5.27039f
C21 VDD2.n2 B 3.34314f
C22 VDD2.t1 B 0.453311f
C23 VDD2.t2 B 0.453311f
C24 VDD2.n3 B 4.12502f
C25 VN.t0 B 0.57029f
C26 VN.n0 B 0.236843f
C27 VN.t1 B 0.567089f
C28 VN.n1 B 0.221063f
C29 VN.t2 B 0.57029f
C30 VN.n2 B 0.23676f
C31 VN.n3 B 0.119136f
C32 VN.t3 B 0.57029f
C33 VN.n4 B 0.236843f
C34 VN.t5 B 0.57029f
C35 VN.t4 B 0.567089f
C36 VN.n5 B 0.221063f
C37 VN.n6 B 0.23676f
C38 VN.n7 B 2.8687f
C39 VDD1.t2 B 5.26937f
C40 VDD1.t5 B 5.26856f
C41 VDD1.t3 B 0.452995f
C42 VDD1.t4 B 0.452995f
C43 VDD1.n0 B 4.12218f
C44 VDD1.n1 B 2.95387f
C45 VDD1.t0 B 0.452995f
C46 VDD1.t1 B 0.452995f
C47 VDD1.n2 B 4.12185f
C48 VDD1.n3 B 3.29501f
C49 VTAIL.t0 B 0.456471f
C50 VTAIL.t2 B 0.456471f
C51 VTAIL.n0 B 4.04882f
C52 VTAIL.n1 B 0.422735f
C53 VTAIL.t4 B 5.17018f
C54 VTAIL.n2 B 0.574698f
C55 VTAIL.t7 B 0.456471f
C56 VTAIL.t8 B 0.456471f
C57 VTAIL.n3 B 4.04882f
C58 VTAIL.n4 B 2.51635f
C59 VTAIL.t10 B 0.456471f
C60 VTAIL.t11 B 0.456471f
C61 VTAIL.n5 B 4.04883f
C62 VTAIL.n6 B 2.51634f
C63 VTAIL.t3 B 5.17018f
C64 VTAIL.n7 B 0.574692f
C65 VTAIL.t9 B 0.456471f
C66 VTAIL.t5 B 0.456471f
C67 VTAIL.n8 B 4.04883f
C68 VTAIL.n9 B 0.451125f
C69 VTAIL.t6 B 5.17018f
C70 VTAIL.n10 B 2.59394f
C71 VTAIL.t1 B 5.17018f
C72 VTAIL.n11 B 2.57637f
C73 VP.t3 B 0.580505f
C74 VP.n0 B 0.241085f
C75 VP.t5 B 0.577247f
C76 VP.n1 B 0.225022f
C77 VP.t4 B 0.580505f
C78 VP.n2 B 0.241001f
C79 VP.n3 B 2.87821f
C80 VP.n4 B 2.85934f
C81 VP.t2 B 0.577247f
C82 VP.t0 B 0.580505f
C83 VP.n5 B 0.241001f
C84 VP.n6 B 0.225022f
C85 VP.t1 B 0.580505f
C86 VP.n7 B 0.241001f
C87 VP.n8 B 0.049542f
.ends

