* NGSPICE file created from diff_pair_sample_1176.ext - technology: sky130A

.subckt diff_pair_sample_1176 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X1 VTAIL.t13 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.79
X3 VTAIL.t11 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X4 VTAIL.t6 VP.t1 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X5 VTAIL.t5 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.79
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.79
X7 VDD1.t1 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.79
X8 VDD1.t6 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.79
X9 VDD2.t5 VN.t2 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X10 VDD1.t3 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X11 VTAIL.t1 VP.t6 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.79
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.79
X13 VDD2.t4 VN.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X14 VDD2.t3 VN.t4 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.79
X15 VTAIL.t14 VN.t5 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.79
X16 VDD2.t1 VN.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=1.4508 ps=8.22 w=3.72 l=2.79
X17 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6138 pd=4.05 as=0.6138 ps=4.05 w=3.72 l=2.79
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0 ps=0 w=3.72 l=2.79
X19 VTAIL.t8 VN.t7 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4508 pd=8.22 as=0.6138 ps=4.05 w=3.72 l=2.79
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n27 VP.n26 161.3
R6 VP.n29 VP.n13 161.3
R7 VP.n31 VP.n30 161.3
R8 VP.n32 VP.n12 161.3
R9 VP.n34 VP.n33 161.3
R10 VP.n35 VP.n11 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n69 VP.n68 161.3
R13 VP.n67 VP.n1 161.3
R14 VP.n66 VP.n65 161.3
R15 VP.n64 VP.n2 161.3
R16 VP.n63 VP.n62 161.3
R17 VP.n61 VP.n3 161.3
R18 VP.n59 VP.n58 161.3
R19 VP.n57 VP.n4 161.3
R20 VP.n56 VP.n55 161.3
R21 VP.n54 VP.n5 161.3
R22 VP.n53 VP.n52 161.3
R23 VP.n51 VP.n6 161.3
R24 VP.n50 VP.n49 161.3
R25 VP.n47 VP.n7 161.3
R26 VP.n46 VP.n45 161.3
R27 VP.n44 VP.n8 161.3
R28 VP.n43 VP.n42 161.3
R29 VP.n41 VP.n9 161.3
R30 VP.n40 VP.n39 68.9556
R31 VP.n70 VP.n0 68.9556
R32 VP.n38 VP.n10 68.9556
R33 VP.n18 VP.t2 63.8957
R34 VP.n18 VP.n17 58.3046
R35 VP.n55 VP.n54 56.4773
R36 VP.n23 VP.n22 56.4773
R37 VP.n46 VP.n8 53.0692
R38 VP.n66 VP.n2 53.0692
R39 VP.n34 VP.n12 53.0692
R40 VP.n39 VP.n38 45.5976
R41 VP.n40 VP.t6 32.1338
R42 VP.n48 VP.t5 32.1338
R43 VP.n60 VP.t0 32.1338
R44 VP.n0 VP.t4 32.1338
R45 VP.n10 VP.t3 32.1338
R46 VP.n28 VP.t1 32.1338
R47 VP.n17 VP.t7 32.1338
R48 VP.n42 VP.n8 27.752
R49 VP.n67 VP.n66 27.752
R50 VP.n35 VP.n34 27.752
R51 VP.n42 VP.n41 24.3439
R52 VP.n47 VP.n46 24.3439
R53 VP.n49 VP.n47 24.3439
R54 VP.n53 VP.n6 24.3439
R55 VP.n54 VP.n53 24.3439
R56 VP.n55 VP.n4 24.3439
R57 VP.n59 VP.n4 24.3439
R58 VP.n62 VP.n61 24.3439
R59 VP.n62 VP.n2 24.3439
R60 VP.n68 VP.n67 24.3439
R61 VP.n36 VP.n35 24.3439
R62 VP.n23 VP.n14 24.3439
R63 VP.n27 VP.n14 24.3439
R64 VP.n30 VP.n29 24.3439
R65 VP.n30 VP.n12 24.3439
R66 VP.n21 VP.n16 24.3439
R67 VP.n22 VP.n21 24.3439
R68 VP.n41 VP.n40 20.9359
R69 VP.n68 VP.n0 20.9359
R70 VP.n36 VP.n10 20.9359
R71 VP.n48 VP.n6 15.0934
R72 VP.n60 VP.n59 15.0934
R73 VP.n28 VP.n27 15.0934
R74 VP.n17 VP.n16 15.0934
R75 VP.n49 VP.n48 9.251
R76 VP.n61 VP.n60 9.251
R77 VP.n29 VP.n28 9.251
R78 VP.n19 VP.n18 5.48081
R79 VP.n38 VP.n37 0.355081
R80 VP.n39 VP.n9 0.355081
R81 VP.n70 VP.n69 0.355081
R82 VP VP.n70 0.26685
R83 VP.n20 VP.n19 0.189894
R84 VP.n20 VP.n15 0.189894
R85 VP.n24 VP.n15 0.189894
R86 VP.n25 VP.n24 0.189894
R87 VP.n26 VP.n25 0.189894
R88 VP.n26 VP.n13 0.189894
R89 VP.n31 VP.n13 0.189894
R90 VP.n32 VP.n31 0.189894
R91 VP.n33 VP.n32 0.189894
R92 VP.n33 VP.n11 0.189894
R93 VP.n37 VP.n11 0.189894
R94 VP.n43 VP.n9 0.189894
R95 VP.n44 VP.n43 0.189894
R96 VP.n45 VP.n44 0.189894
R97 VP.n45 VP.n7 0.189894
R98 VP.n50 VP.n7 0.189894
R99 VP.n51 VP.n50 0.189894
R100 VP.n52 VP.n51 0.189894
R101 VP.n52 VP.n5 0.189894
R102 VP.n56 VP.n5 0.189894
R103 VP.n57 VP.n56 0.189894
R104 VP.n58 VP.n57 0.189894
R105 VP.n58 VP.n3 0.189894
R106 VP.n63 VP.n3 0.189894
R107 VP.n64 VP.n63 0.189894
R108 VP.n65 VP.n64 0.189894
R109 VP.n65 VP.n1 0.189894
R110 VP.n69 VP.n1 0.189894
R111 VDD1 VDD1.n0 75.4436
R112 VDD1.n3 VDD1.n2 75.33
R113 VDD1.n3 VDD1.n1 75.33
R114 VDD1.n5 VDD1.n4 74.0406
R115 VDD1.n5 VDD1.n3 39.6087
R116 VDD1.n4 VDD1.t0 5.32308
R117 VDD1.n4 VDD1.t1 5.32308
R118 VDD1.n0 VDD1.t7 5.32308
R119 VDD1.n0 VDD1.t2 5.32308
R120 VDD1.n2 VDD1.t5 5.32308
R121 VDD1.n2 VDD1.t6 5.32308
R122 VDD1.n1 VDD1.t4 5.32308
R123 VDD1.n1 VDD1.t3 5.32308
R124 VDD1 VDD1.n5 1.28714
R125 VTAIL.n14 VTAIL.t4 62.6844
R126 VTAIL.n11 VTAIL.t5 62.6844
R127 VTAIL.n10 VTAIL.t9 62.6844
R128 VTAIL.n7 VTAIL.t8 62.6844
R129 VTAIL.n15 VTAIL.t15 62.6843
R130 VTAIL.n2 VTAIL.t14 62.6843
R131 VTAIL.n3 VTAIL.t3 62.6843
R132 VTAIL.n6 VTAIL.t1 62.6843
R133 VTAIL.n13 VTAIL.n12 57.3618
R134 VTAIL.n9 VTAIL.n8 57.3618
R135 VTAIL.n1 VTAIL.n0 57.3617
R136 VTAIL.n5 VTAIL.n4 57.3617
R137 VTAIL.n15 VTAIL.n14 18.2634
R138 VTAIL.n7 VTAIL.n6 18.2634
R139 VTAIL.n0 VTAIL.t10 5.32308
R140 VTAIL.n0 VTAIL.t11 5.32308
R141 VTAIL.n4 VTAIL.t2 5.32308
R142 VTAIL.n4 VTAIL.t7 5.32308
R143 VTAIL.n12 VTAIL.t0 5.32308
R144 VTAIL.n12 VTAIL.t6 5.32308
R145 VTAIL.n8 VTAIL.t12 5.32308
R146 VTAIL.n8 VTAIL.t13 5.32308
R147 VTAIL.n9 VTAIL.n7 2.69016
R148 VTAIL.n10 VTAIL.n9 2.69016
R149 VTAIL.n13 VTAIL.n11 2.69016
R150 VTAIL.n14 VTAIL.n13 2.69016
R151 VTAIL.n6 VTAIL.n5 2.69016
R152 VTAIL.n5 VTAIL.n3 2.69016
R153 VTAIL.n2 VTAIL.n1 2.69016
R154 VTAIL VTAIL.n15 2.63197
R155 VTAIL.n11 VTAIL.n10 0.470328
R156 VTAIL.n3 VTAIL.n2 0.470328
R157 VTAIL VTAIL.n1 0.0586897
R158 B.n579 B.n578 585
R159 B.n581 B.n126 585
R160 B.n584 B.n583 585
R161 B.n585 B.n125 585
R162 B.n587 B.n586 585
R163 B.n589 B.n124 585
R164 B.n592 B.n591 585
R165 B.n593 B.n123 585
R166 B.n595 B.n594 585
R167 B.n597 B.n122 585
R168 B.n600 B.n599 585
R169 B.n601 B.n121 585
R170 B.n603 B.n602 585
R171 B.n605 B.n120 585
R172 B.n608 B.n607 585
R173 B.n609 B.n116 585
R174 B.n611 B.n610 585
R175 B.n613 B.n115 585
R176 B.n616 B.n615 585
R177 B.n617 B.n114 585
R178 B.n619 B.n618 585
R179 B.n621 B.n113 585
R180 B.n624 B.n623 585
R181 B.n625 B.n112 585
R182 B.n627 B.n626 585
R183 B.n629 B.n111 585
R184 B.n632 B.n631 585
R185 B.n634 B.n108 585
R186 B.n636 B.n635 585
R187 B.n638 B.n107 585
R188 B.n641 B.n640 585
R189 B.n642 B.n106 585
R190 B.n644 B.n643 585
R191 B.n646 B.n105 585
R192 B.n649 B.n648 585
R193 B.n650 B.n104 585
R194 B.n652 B.n651 585
R195 B.n654 B.n103 585
R196 B.n657 B.n656 585
R197 B.n658 B.n102 585
R198 B.n660 B.n659 585
R199 B.n662 B.n101 585
R200 B.n665 B.n664 585
R201 B.n666 B.n100 585
R202 B.n577 B.n98 585
R203 B.n669 B.n98 585
R204 B.n576 B.n97 585
R205 B.n670 B.n97 585
R206 B.n575 B.n96 585
R207 B.n671 B.n96 585
R208 B.n574 B.n573 585
R209 B.n573 B.n92 585
R210 B.n572 B.n91 585
R211 B.n677 B.n91 585
R212 B.n571 B.n90 585
R213 B.n678 B.n90 585
R214 B.n570 B.n89 585
R215 B.n679 B.n89 585
R216 B.n569 B.n568 585
R217 B.n568 B.n88 585
R218 B.n567 B.n84 585
R219 B.n685 B.n84 585
R220 B.n566 B.n83 585
R221 B.n686 B.n83 585
R222 B.n565 B.n82 585
R223 B.n687 B.n82 585
R224 B.n564 B.n563 585
R225 B.n563 B.n78 585
R226 B.n562 B.n77 585
R227 B.n693 B.n77 585
R228 B.n561 B.n76 585
R229 B.n694 B.n76 585
R230 B.n560 B.n75 585
R231 B.n695 B.n75 585
R232 B.n559 B.n558 585
R233 B.n558 B.n71 585
R234 B.n557 B.n70 585
R235 B.n701 B.n70 585
R236 B.n556 B.n69 585
R237 B.n702 B.n69 585
R238 B.n555 B.n68 585
R239 B.n703 B.n68 585
R240 B.n554 B.n553 585
R241 B.n553 B.n64 585
R242 B.n552 B.n63 585
R243 B.n709 B.n63 585
R244 B.n551 B.n62 585
R245 B.n710 B.n62 585
R246 B.n550 B.n61 585
R247 B.n711 B.n61 585
R248 B.n549 B.n548 585
R249 B.n548 B.n57 585
R250 B.n547 B.n56 585
R251 B.n717 B.n56 585
R252 B.n546 B.n55 585
R253 B.n718 B.n55 585
R254 B.n545 B.n54 585
R255 B.n719 B.n54 585
R256 B.n544 B.n543 585
R257 B.n543 B.n50 585
R258 B.n542 B.n49 585
R259 B.n725 B.n49 585
R260 B.n541 B.n48 585
R261 B.n726 B.n48 585
R262 B.n540 B.n47 585
R263 B.n727 B.n47 585
R264 B.n539 B.n538 585
R265 B.n538 B.n43 585
R266 B.n537 B.n42 585
R267 B.n733 B.n42 585
R268 B.n536 B.n41 585
R269 B.n734 B.n41 585
R270 B.n535 B.n40 585
R271 B.n735 B.n40 585
R272 B.n534 B.n533 585
R273 B.n533 B.n36 585
R274 B.n532 B.n35 585
R275 B.n741 B.n35 585
R276 B.n531 B.n34 585
R277 B.n742 B.n34 585
R278 B.n530 B.n33 585
R279 B.n743 B.n33 585
R280 B.n529 B.n528 585
R281 B.n528 B.n29 585
R282 B.n527 B.n28 585
R283 B.n749 B.n28 585
R284 B.n526 B.n27 585
R285 B.n750 B.n27 585
R286 B.n525 B.n26 585
R287 B.n751 B.n26 585
R288 B.n524 B.n523 585
R289 B.n523 B.n22 585
R290 B.n522 B.n21 585
R291 B.n757 B.n21 585
R292 B.n521 B.n20 585
R293 B.n758 B.n20 585
R294 B.n520 B.n19 585
R295 B.n759 B.n19 585
R296 B.n519 B.n518 585
R297 B.n518 B.n18 585
R298 B.n517 B.n14 585
R299 B.n765 B.n14 585
R300 B.n516 B.n13 585
R301 B.n766 B.n13 585
R302 B.n515 B.n12 585
R303 B.n767 B.n12 585
R304 B.n514 B.n513 585
R305 B.n513 B.n8 585
R306 B.n512 B.n7 585
R307 B.n773 B.n7 585
R308 B.n511 B.n6 585
R309 B.n774 B.n6 585
R310 B.n510 B.n5 585
R311 B.n775 B.n5 585
R312 B.n509 B.n508 585
R313 B.n508 B.n4 585
R314 B.n507 B.n127 585
R315 B.n507 B.n506 585
R316 B.n497 B.n128 585
R317 B.n129 B.n128 585
R318 B.n499 B.n498 585
R319 B.n500 B.n499 585
R320 B.n496 B.n134 585
R321 B.n134 B.n133 585
R322 B.n495 B.n494 585
R323 B.n494 B.n493 585
R324 B.n136 B.n135 585
R325 B.n486 B.n136 585
R326 B.n485 B.n484 585
R327 B.n487 B.n485 585
R328 B.n483 B.n141 585
R329 B.n141 B.n140 585
R330 B.n482 B.n481 585
R331 B.n481 B.n480 585
R332 B.n143 B.n142 585
R333 B.n144 B.n143 585
R334 B.n473 B.n472 585
R335 B.n474 B.n473 585
R336 B.n471 B.n149 585
R337 B.n149 B.n148 585
R338 B.n470 B.n469 585
R339 B.n469 B.n468 585
R340 B.n151 B.n150 585
R341 B.n152 B.n151 585
R342 B.n461 B.n460 585
R343 B.n462 B.n461 585
R344 B.n459 B.n157 585
R345 B.n157 B.n156 585
R346 B.n458 B.n457 585
R347 B.n457 B.n456 585
R348 B.n159 B.n158 585
R349 B.n160 B.n159 585
R350 B.n449 B.n448 585
R351 B.n450 B.n449 585
R352 B.n447 B.n165 585
R353 B.n165 B.n164 585
R354 B.n446 B.n445 585
R355 B.n445 B.n444 585
R356 B.n167 B.n166 585
R357 B.n168 B.n167 585
R358 B.n437 B.n436 585
R359 B.n438 B.n437 585
R360 B.n435 B.n172 585
R361 B.n176 B.n172 585
R362 B.n434 B.n433 585
R363 B.n433 B.n432 585
R364 B.n174 B.n173 585
R365 B.n175 B.n174 585
R366 B.n425 B.n424 585
R367 B.n426 B.n425 585
R368 B.n423 B.n181 585
R369 B.n181 B.n180 585
R370 B.n422 B.n421 585
R371 B.n421 B.n420 585
R372 B.n183 B.n182 585
R373 B.n184 B.n183 585
R374 B.n413 B.n412 585
R375 B.n414 B.n413 585
R376 B.n411 B.n189 585
R377 B.n189 B.n188 585
R378 B.n410 B.n409 585
R379 B.n409 B.n408 585
R380 B.n191 B.n190 585
R381 B.n192 B.n191 585
R382 B.n401 B.n400 585
R383 B.n402 B.n401 585
R384 B.n399 B.n197 585
R385 B.n197 B.n196 585
R386 B.n398 B.n397 585
R387 B.n397 B.n396 585
R388 B.n199 B.n198 585
R389 B.n200 B.n199 585
R390 B.n389 B.n388 585
R391 B.n390 B.n389 585
R392 B.n387 B.n205 585
R393 B.n205 B.n204 585
R394 B.n386 B.n385 585
R395 B.n385 B.n384 585
R396 B.n207 B.n206 585
R397 B.n208 B.n207 585
R398 B.n377 B.n376 585
R399 B.n378 B.n377 585
R400 B.n375 B.n213 585
R401 B.n213 B.n212 585
R402 B.n374 B.n373 585
R403 B.n373 B.n372 585
R404 B.n215 B.n214 585
R405 B.n365 B.n215 585
R406 B.n364 B.n363 585
R407 B.n366 B.n364 585
R408 B.n362 B.n220 585
R409 B.n220 B.n219 585
R410 B.n361 B.n360 585
R411 B.n360 B.n359 585
R412 B.n222 B.n221 585
R413 B.n223 B.n222 585
R414 B.n352 B.n351 585
R415 B.n353 B.n352 585
R416 B.n350 B.n228 585
R417 B.n228 B.n227 585
R418 B.n349 B.n348 585
R419 B.n348 B.n347 585
R420 B.n344 B.n232 585
R421 B.n343 B.n342 585
R422 B.n340 B.n233 585
R423 B.n340 B.n231 585
R424 B.n339 B.n338 585
R425 B.n337 B.n336 585
R426 B.n335 B.n235 585
R427 B.n333 B.n332 585
R428 B.n331 B.n236 585
R429 B.n330 B.n329 585
R430 B.n327 B.n237 585
R431 B.n325 B.n324 585
R432 B.n323 B.n238 585
R433 B.n322 B.n321 585
R434 B.n319 B.n239 585
R435 B.n317 B.n316 585
R436 B.n315 B.n240 585
R437 B.n314 B.n313 585
R438 B.n311 B.n310 585
R439 B.n309 B.n308 585
R440 B.n307 B.n245 585
R441 B.n305 B.n304 585
R442 B.n303 B.n246 585
R443 B.n302 B.n301 585
R444 B.n299 B.n247 585
R445 B.n297 B.n296 585
R446 B.n295 B.n248 585
R447 B.n294 B.n293 585
R448 B.n291 B.n290 585
R449 B.n289 B.n288 585
R450 B.n287 B.n253 585
R451 B.n285 B.n284 585
R452 B.n283 B.n254 585
R453 B.n282 B.n281 585
R454 B.n279 B.n255 585
R455 B.n277 B.n276 585
R456 B.n275 B.n256 585
R457 B.n274 B.n273 585
R458 B.n271 B.n257 585
R459 B.n269 B.n268 585
R460 B.n267 B.n258 585
R461 B.n266 B.n265 585
R462 B.n263 B.n259 585
R463 B.n261 B.n260 585
R464 B.n230 B.n229 585
R465 B.n231 B.n230 585
R466 B.n346 B.n345 585
R467 B.n347 B.n346 585
R468 B.n226 B.n225 585
R469 B.n227 B.n226 585
R470 B.n355 B.n354 585
R471 B.n354 B.n353 585
R472 B.n356 B.n224 585
R473 B.n224 B.n223 585
R474 B.n358 B.n357 585
R475 B.n359 B.n358 585
R476 B.n218 B.n217 585
R477 B.n219 B.n218 585
R478 B.n368 B.n367 585
R479 B.n367 B.n366 585
R480 B.n369 B.n216 585
R481 B.n365 B.n216 585
R482 B.n371 B.n370 585
R483 B.n372 B.n371 585
R484 B.n211 B.n210 585
R485 B.n212 B.n211 585
R486 B.n380 B.n379 585
R487 B.n379 B.n378 585
R488 B.n381 B.n209 585
R489 B.n209 B.n208 585
R490 B.n383 B.n382 585
R491 B.n384 B.n383 585
R492 B.n203 B.n202 585
R493 B.n204 B.n203 585
R494 B.n392 B.n391 585
R495 B.n391 B.n390 585
R496 B.n393 B.n201 585
R497 B.n201 B.n200 585
R498 B.n395 B.n394 585
R499 B.n396 B.n395 585
R500 B.n195 B.n194 585
R501 B.n196 B.n195 585
R502 B.n404 B.n403 585
R503 B.n403 B.n402 585
R504 B.n405 B.n193 585
R505 B.n193 B.n192 585
R506 B.n407 B.n406 585
R507 B.n408 B.n407 585
R508 B.n187 B.n186 585
R509 B.n188 B.n187 585
R510 B.n416 B.n415 585
R511 B.n415 B.n414 585
R512 B.n417 B.n185 585
R513 B.n185 B.n184 585
R514 B.n419 B.n418 585
R515 B.n420 B.n419 585
R516 B.n179 B.n178 585
R517 B.n180 B.n179 585
R518 B.n428 B.n427 585
R519 B.n427 B.n426 585
R520 B.n429 B.n177 585
R521 B.n177 B.n175 585
R522 B.n431 B.n430 585
R523 B.n432 B.n431 585
R524 B.n171 B.n170 585
R525 B.n176 B.n171 585
R526 B.n440 B.n439 585
R527 B.n439 B.n438 585
R528 B.n441 B.n169 585
R529 B.n169 B.n168 585
R530 B.n443 B.n442 585
R531 B.n444 B.n443 585
R532 B.n163 B.n162 585
R533 B.n164 B.n163 585
R534 B.n452 B.n451 585
R535 B.n451 B.n450 585
R536 B.n453 B.n161 585
R537 B.n161 B.n160 585
R538 B.n455 B.n454 585
R539 B.n456 B.n455 585
R540 B.n155 B.n154 585
R541 B.n156 B.n155 585
R542 B.n464 B.n463 585
R543 B.n463 B.n462 585
R544 B.n465 B.n153 585
R545 B.n153 B.n152 585
R546 B.n467 B.n466 585
R547 B.n468 B.n467 585
R548 B.n147 B.n146 585
R549 B.n148 B.n147 585
R550 B.n476 B.n475 585
R551 B.n475 B.n474 585
R552 B.n477 B.n145 585
R553 B.n145 B.n144 585
R554 B.n479 B.n478 585
R555 B.n480 B.n479 585
R556 B.n139 B.n138 585
R557 B.n140 B.n139 585
R558 B.n489 B.n488 585
R559 B.n488 B.n487 585
R560 B.n490 B.n137 585
R561 B.n486 B.n137 585
R562 B.n492 B.n491 585
R563 B.n493 B.n492 585
R564 B.n132 B.n131 585
R565 B.n133 B.n132 585
R566 B.n502 B.n501 585
R567 B.n501 B.n500 585
R568 B.n503 B.n130 585
R569 B.n130 B.n129 585
R570 B.n505 B.n504 585
R571 B.n506 B.n505 585
R572 B.n2 B.n0 585
R573 B.n4 B.n2 585
R574 B.n3 B.n1 585
R575 B.n774 B.n3 585
R576 B.n772 B.n771 585
R577 B.n773 B.n772 585
R578 B.n770 B.n9 585
R579 B.n9 B.n8 585
R580 B.n769 B.n768 585
R581 B.n768 B.n767 585
R582 B.n11 B.n10 585
R583 B.n766 B.n11 585
R584 B.n764 B.n763 585
R585 B.n765 B.n764 585
R586 B.n762 B.n15 585
R587 B.n18 B.n15 585
R588 B.n761 B.n760 585
R589 B.n760 B.n759 585
R590 B.n17 B.n16 585
R591 B.n758 B.n17 585
R592 B.n756 B.n755 585
R593 B.n757 B.n756 585
R594 B.n754 B.n23 585
R595 B.n23 B.n22 585
R596 B.n753 B.n752 585
R597 B.n752 B.n751 585
R598 B.n25 B.n24 585
R599 B.n750 B.n25 585
R600 B.n748 B.n747 585
R601 B.n749 B.n748 585
R602 B.n746 B.n30 585
R603 B.n30 B.n29 585
R604 B.n745 B.n744 585
R605 B.n744 B.n743 585
R606 B.n32 B.n31 585
R607 B.n742 B.n32 585
R608 B.n740 B.n739 585
R609 B.n741 B.n740 585
R610 B.n738 B.n37 585
R611 B.n37 B.n36 585
R612 B.n737 B.n736 585
R613 B.n736 B.n735 585
R614 B.n39 B.n38 585
R615 B.n734 B.n39 585
R616 B.n732 B.n731 585
R617 B.n733 B.n732 585
R618 B.n730 B.n44 585
R619 B.n44 B.n43 585
R620 B.n729 B.n728 585
R621 B.n728 B.n727 585
R622 B.n46 B.n45 585
R623 B.n726 B.n46 585
R624 B.n724 B.n723 585
R625 B.n725 B.n724 585
R626 B.n722 B.n51 585
R627 B.n51 B.n50 585
R628 B.n721 B.n720 585
R629 B.n720 B.n719 585
R630 B.n53 B.n52 585
R631 B.n718 B.n53 585
R632 B.n716 B.n715 585
R633 B.n717 B.n716 585
R634 B.n714 B.n58 585
R635 B.n58 B.n57 585
R636 B.n713 B.n712 585
R637 B.n712 B.n711 585
R638 B.n60 B.n59 585
R639 B.n710 B.n60 585
R640 B.n708 B.n707 585
R641 B.n709 B.n708 585
R642 B.n706 B.n65 585
R643 B.n65 B.n64 585
R644 B.n705 B.n704 585
R645 B.n704 B.n703 585
R646 B.n67 B.n66 585
R647 B.n702 B.n67 585
R648 B.n700 B.n699 585
R649 B.n701 B.n700 585
R650 B.n698 B.n72 585
R651 B.n72 B.n71 585
R652 B.n697 B.n696 585
R653 B.n696 B.n695 585
R654 B.n74 B.n73 585
R655 B.n694 B.n74 585
R656 B.n692 B.n691 585
R657 B.n693 B.n692 585
R658 B.n690 B.n79 585
R659 B.n79 B.n78 585
R660 B.n689 B.n688 585
R661 B.n688 B.n687 585
R662 B.n81 B.n80 585
R663 B.n686 B.n81 585
R664 B.n684 B.n683 585
R665 B.n685 B.n684 585
R666 B.n682 B.n85 585
R667 B.n88 B.n85 585
R668 B.n681 B.n680 585
R669 B.n680 B.n679 585
R670 B.n87 B.n86 585
R671 B.n678 B.n87 585
R672 B.n676 B.n675 585
R673 B.n677 B.n676 585
R674 B.n674 B.n93 585
R675 B.n93 B.n92 585
R676 B.n673 B.n672 585
R677 B.n672 B.n671 585
R678 B.n95 B.n94 585
R679 B.n670 B.n95 585
R680 B.n668 B.n667 585
R681 B.n669 B.n668 585
R682 B.n777 B.n776 585
R683 B.n776 B.n775 585
R684 B.n346 B.n232 506.916
R685 B.n668 B.n100 506.916
R686 B.n348 B.n230 506.916
R687 B.n579 B.n98 506.916
R688 B.n580 B.n99 256.663
R689 B.n582 B.n99 256.663
R690 B.n588 B.n99 256.663
R691 B.n590 B.n99 256.663
R692 B.n596 B.n99 256.663
R693 B.n598 B.n99 256.663
R694 B.n604 B.n99 256.663
R695 B.n606 B.n99 256.663
R696 B.n612 B.n99 256.663
R697 B.n614 B.n99 256.663
R698 B.n620 B.n99 256.663
R699 B.n622 B.n99 256.663
R700 B.n628 B.n99 256.663
R701 B.n630 B.n99 256.663
R702 B.n637 B.n99 256.663
R703 B.n639 B.n99 256.663
R704 B.n645 B.n99 256.663
R705 B.n647 B.n99 256.663
R706 B.n653 B.n99 256.663
R707 B.n655 B.n99 256.663
R708 B.n661 B.n99 256.663
R709 B.n663 B.n99 256.663
R710 B.n341 B.n231 256.663
R711 B.n234 B.n231 256.663
R712 B.n334 B.n231 256.663
R713 B.n328 B.n231 256.663
R714 B.n326 B.n231 256.663
R715 B.n320 B.n231 256.663
R716 B.n318 B.n231 256.663
R717 B.n312 B.n231 256.663
R718 B.n244 B.n231 256.663
R719 B.n306 B.n231 256.663
R720 B.n300 B.n231 256.663
R721 B.n298 B.n231 256.663
R722 B.n292 B.n231 256.663
R723 B.n252 B.n231 256.663
R724 B.n286 B.n231 256.663
R725 B.n280 B.n231 256.663
R726 B.n278 B.n231 256.663
R727 B.n272 B.n231 256.663
R728 B.n270 B.n231 256.663
R729 B.n264 B.n231 256.663
R730 B.n262 B.n231 256.663
R731 B.n249 B.t19 241.115
R732 B.n117 B.t12 241.115
R733 B.n241 B.t8 240.804
R734 B.n109 B.t16 240.804
R735 B.n346 B.n226 163.367
R736 B.n354 B.n226 163.367
R737 B.n354 B.n224 163.367
R738 B.n358 B.n224 163.367
R739 B.n358 B.n218 163.367
R740 B.n367 B.n218 163.367
R741 B.n367 B.n216 163.367
R742 B.n371 B.n216 163.367
R743 B.n371 B.n211 163.367
R744 B.n379 B.n211 163.367
R745 B.n379 B.n209 163.367
R746 B.n383 B.n209 163.367
R747 B.n383 B.n203 163.367
R748 B.n391 B.n203 163.367
R749 B.n391 B.n201 163.367
R750 B.n395 B.n201 163.367
R751 B.n395 B.n195 163.367
R752 B.n403 B.n195 163.367
R753 B.n403 B.n193 163.367
R754 B.n407 B.n193 163.367
R755 B.n407 B.n187 163.367
R756 B.n415 B.n187 163.367
R757 B.n415 B.n185 163.367
R758 B.n419 B.n185 163.367
R759 B.n419 B.n179 163.367
R760 B.n427 B.n179 163.367
R761 B.n427 B.n177 163.367
R762 B.n431 B.n177 163.367
R763 B.n431 B.n171 163.367
R764 B.n439 B.n171 163.367
R765 B.n439 B.n169 163.367
R766 B.n443 B.n169 163.367
R767 B.n443 B.n163 163.367
R768 B.n451 B.n163 163.367
R769 B.n451 B.n161 163.367
R770 B.n455 B.n161 163.367
R771 B.n455 B.n155 163.367
R772 B.n463 B.n155 163.367
R773 B.n463 B.n153 163.367
R774 B.n467 B.n153 163.367
R775 B.n467 B.n147 163.367
R776 B.n475 B.n147 163.367
R777 B.n475 B.n145 163.367
R778 B.n479 B.n145 163.367
R779 B.n479 B.n139 163.367
R780 B.n488 B.n139 163.367
R781 B.n488 B.n137 163.367
R782 B.n492 B.n137 163.367
R783 B.n492 B.n132 163.367
R784 B.n501 B.n132 163.367
R785 B.n501 B.n130 163.367
R786 B.n505 B.n130 163.367
R787 B.n505 B.n2 163.367
R788 B.n776 B.n2 163.367
R789 B.n776 B.n3 163.367
R790 B.n772 B.n3 163.367
R791 B.n772 B.n9 163.367
R792 B.n768 B.n9 163.367
R793 B.n768 B.n11 163.367
R794 B.n764 B.n11 163.367
R795 B.n764 B.n15 163.367
R796 B.n760 B.n15 163.367
R797 B.n760 B.n17 163.367
R798 B.n756 B.n17 163.367
R799 B.n756 B.n23 163.367
R800 B.n752 B.n23 163.367
R801 B.n752 B.n25 163.367
R802 B.n748 B.n25 163.367
R803 B.n748 B.n30 163.367
R804 B.n744 B.n30 163.367
R805 B.n744 B.n32 163.367
R806 B.n740 B.n32 163.367
R807 B.n740 B.n37 163.367
R808 B.n736 B.n37 163.367
R809 B.n736 B.n39 163.367
R810 B.n732 B.n39 163.367
R811 B.n732 B.n44 163.367
R812 B.n728 B.n44 163.367
R813 B.n728 B.n46 163.367
R814 B.n724 B.n46 163.367
R815 B.n724 B.n51 163.367
R816 B.n720 B.n51 163.367
R817 B.n720 B.n53 163.367
R818 B.n716 B.n53 163.367
R819 B.n716 B.n58 163.367
R820 B.n712 B.n58 163.367
R821 B.n712 B.n60 163.367
R822 B.n708 B.n60 163.367
R823 B.n708 B.n65 163.367
R824 B.n704 B.n65 163.367
R825 B.n704 B.n67 163.367
R826 B.n700 B.n67 163.367
R827 B.n700 B.n72 163.367
R828 B.n696 B.n72 163.367
R829 B.n696 B.n74 163.367
R830 B.n692 B.n74 163.367
R831 B.n692 B.n79 163.367
R832 B.n688 B.n79 163.367
R833 B.n688 B.n81 163.367
R834 B.n684 B.n81 163.367
R835 B.n684 B.n85 163.367
R836 B.n680 B.n85 163.367
R837 B.n680 B.n87 163.367
R838 B.n676 B.n87 163.367
R839 B.n676 B.n93 163.367
R840 B.n672 B.n93 163.367
R841 B.n672 B.n95 163.367
R842 B.n668 B.n95 163.367
R843 B.n342 B.n340 163.367
R844 B.n340 B.n339 163.367
R845 B.n336 B.n335 163.367
R846 B.n333 B.n236 163.367
R847 B.n329 B.n327 163.367
R848 B.n325 B.n238 163.367
R849 B.n321 B.n319 163.367
R850 B.n317 B.n240 163.367
R851 B.n313 B.n311 163.367
R852 B.n308 B.n307 163.367
R853 B.n305 B.n246 163.367
R854 B.n301 B.n299 163.367
R855 B.n297 B.n248 163.367
R856 B.n293 B.n291 163.367
R857 B.n288 B.n287 163.367
R858 B.n285 B.n254 163.367
R859 B.n281 B.n279 163.367
R860 B.n277 B.n256 163.367
R861 B.n273 B.n271 163.367
R862 B.n269 B.n258 163.367
R863 B.n265 B.n263 163.367
R864 B.n261 B.n230 163.367
R865 B.n348 B.n228 163.367
R866 B.n352 B.n228 163.367
R867 B.n352 B.n222 163.367
R868 B.n360 B.n222 163.367
R869 B.n360 B.n220 163.367
R870 B.n364 B.n220 163.367
R871 B.n364 B.n215 163.367
R872 B.n373 B.n215 163.367
R873 B.n373 B.n213 163.367
R874 B.n377 B.n213 163.367
R875 B.n377 B.n207 163.367
R876 B.n385 B.n207 163.367
R877 B.n385 B.n205 163.367
R878 B.n389 B.n205 163.367
R879 B.n389 B.n199 163.367
R880 B.n397 B.n199 163.367
R881 B.n397 B.n197 163.367
R882 B.n401 B.n197 163.367
R883 B.n401 B.n191 163.367
R884 B.n409 B.n191 163.367
R885 B.n409 B.n189 163.367
R886 B.n413 B.n189 163.367
R887 B.n413 B.n183 163.367
R888 B.n421 B.n183 163.367
R889 B.n421 B.n181 163.367
R890 B.n425 B.n181 163.367
R891 B.n425 B.n174 163.367
R892 B.n433 B.n174 163.367
R893 B.n433 B.n172 163.367
R894 B.n437 B.n172 163.367
R895 B.n437 B.n167 163.367
R896 B.n445 B.n167 163.367
R897 B.n445 B.n165 163.367
R898 B.n449 B.n165 163.367
R899 B.n449 B.n159 163.367
R900 B.n457 B.n159 163.367
R901 B.n457 B.n157 163.367
R902 B.n461 B.n157 163.367
R903 B.n461 B.n151 163.367
R904 B.n469 B.n151 163.367
R905 B.n469 B.n149 163.367
R906 B.n473 B.n149 163.367
R907 B.n473 B.n143 163.367
R908 B.n481 B.n143 163.367
R909 B.n481 B.n141 163.367
R910 B.n485 B.n141 163.367
R911 B.n485 B.n136 163.367
R912 B.n494 B.n136 163.367
R913 B.n494 B.n134 163.367
R914 B.n499 B.n134 163.367
R915 B.n499 B.n128 163.367
R916 B.n507 B.n128 163.367
R917 B.n508 B.n507 163.367
R918 B.n508 B.n5 163.367
R919 B.n6 B.n5 163.367
R920 B.n7 B.n6 163.367
R921 B.n513 B.n7 163.367
R922 B.n513 B.n12 163.367
R923 B.n13 B.n12 163.367
R924 B.n14 B.n13 163.367
R925 B.n518 B.n14 163.367
R926 B.n518 B.n19 163.367
R927 B.n20 B.n19 163.367
R928 B.n21 B.n20 163.367
R929 B.n523 B.n21 163.367
R930 B.n523 B.n26 163.367
R931 B.n27 B.n26 163.367
R932 B.n28 B.n27 163.367
R933 B.n528 B.n28 163.367
R934 B.n528 B.n33 163.367
R935 B.n34 B.n33 163.367
R936 B.n35 B.n34 163.367
R937 B.n533 B.n35 163.367
R938 B.n533 B.n40 163.367
R939 B.n41 B.n40 163.367
R940 B.n42 B.n41 163.367
R941 B.n538 B.n42 163.367
R942 B.n538 B.n47 163.367
R943 B.n48 B.n47 163.367
R944 B.n49 B.n48 163.367
R945 B.n543 B.n49 163.367
R946 B.n543 B.n54 163.367
R947 B.n55 B.n54 163.367
R948 B.n56 B.n55 163.367
R949 B.n548 B.n56 163.367
R950 B.n548 B.n61 163.367
R951 B.n62 B.n61 163.367
R952 B.n63 B.n62 163.367
R953 B.n553 B.n63 163.367
R954 B.n553 B.n68 163.367
R955 B.n69 B.n68 163.367
R956 B.n70 B.n69 163.367
R957 B.n558 B.n70 163.367
R958 B.n558 B.n75 163.367
R959 B.n76 B.n75 163.367
R960 B.n77 B.n76 163.367
R961 B.n563 B.n77 163.367
R962 B.n563 B.n82 163.367
R963 B.n83 B.n82 163.367
R964 B.n84 B.n83 163.367
R965 B.n568 B.n84 163.367
R966 B.n568 B.n89 163.367
R967 B.n90 B.n89 163.367
R968 B.n91 B.n90 163.367
R969 B.n573 B.n91 163.367
R970 B.n573 B.n96 163.367
R971 B.n97 B.n96 163.367
R972 B.n98 B.n97 163.367
R973 B.n664 B.n662 163.367
R974 B.n660 B.n102 163.367
R975 B.n656 B.n654 163.367
R976 B.n652 B.n104 163.367
R977 B.n648 B.n646 163.367
R978 B.n644 B.n106 163.367
R979 B.n640 B.n638 163.367
R980 B.n636 B.n108 163.367
R981 B.n631 B.n629 163.367
R982 B.n627 B.n112 163.367
R983 B.n623 B.n621 163.367
R984 B.n619 B.n114 163.367
R985 B.n615 B.n613 163.367
R986 B.n611 B.n116 163.367
R987 B.n607 B.n605 163.367
R988 B.n603 B.n121 163.367
R989 B.n599 B.n597 163.367
R990 B.n595 B.n123 163.367
R991 B.n591 B.n589 163.367
R992 B.n587 B.n125 163.367
R993 B.n583 B.n581 163.367
R994 B.n347 B.n231 150.417
R995 B.n669 B.n99 150.417
R996 B.n249 B.t21 139.194
R997 B.n117 B.t14 139.194
R998 B.n241 B.t11 139.19
R999 B.n109 B.t17 139.19
R1000 B.n347 B.n227 83.1578
R1001 B.n353 B.n227 83.1578
R1002 B.n353 B.n223 83.1578
R1003 B.n359 B.n223 83.1578
R1004 B.n359 B.n219 83.1578
R1005 B.n366 B.n219 83.1578
R1006 B.n366 B.n365 83.1578
R1007 B.n372 B.n212 83.1578
R1008 B.n378 B.n212 83.1578
R1009 B.n378 B.n208 83.1578
R1010 B.n384 B.n208 83.1578
R1011 B.n384 B.n204 83.1578
R1012 B.n390 B.n204 83.1578
R1013 B.n390 B.n200 83.1578
R1014 B.n396 B.n200 83.1578
R1015 B.n396 B.n196 83.1578
R1016 B.n402 B.n196 83.1578
R1017 B.n402 B.n192 83.1578
R1018 B.n408 B.n192 83.1578
R1019 B.n414 B.n188 83.1578
R1020 B.n414 B.n184 83.1578
R1021 B.n420 B.n184 83.1578
R1022 B.n420 B.n180 83.1578
R1023 B.n426 B.n180 83.1578
R1024 B.n426 B.n175 83.1578
R1025 B.n432 B.n175 83.1578
R1026 B.n432 B.n176 83.1578
R1027 B.n438 B.n168 83.1578
R1028 B.n444 B.n168 83.1578
R1029 B.n444 B.n164 83.1578
R1030 B.n450 B.n164 83.1578
R1031 B.n450 B.n160 83.1578
R1032 B.n456 B.n160 83.1578
R1033 B.n456 B.n156 83.1578
R1034 B.n462 B.n156 83.1578
R1035 B.n468 B.n152 83.1578
R1036 B.n468 B.n148 83.1578
R1037 B.n474 B.n148 83.1578
R1038 B.n474 B.n144 83.1578
R1039 B.n480 B.n144 83.1578
R1040 B.n480 B.n140 83.1578
R1041 B.n487 B.n140 83.1578
R1042 B.n487 B.n486 83.1578
R1043 B.n493 B.n133 83.1578
R1044 B.n500 B.n133 83.1578
R1045 B.n500 B.n129 83.1578
R1046 B.n506 B.n129 83.1578
R1047 B.n506 B.n4 83.1578
R1048 B.n775 B.n4 83.1578
R1049 B.n775 B.n774 83.1578
R1050 B.n774 B.n773 83.1578
R1051 B.n773 B.n8 83.1578
R1052 B.n767 B.n8 83.1578
R1053 B.n767 B.n766 83.1578
R1054 B.n766 B.n765 83.1578
R1055 B.n759 B.n18 83.1578
R1056 B.n759 B.n758 83.1578
R1057 B.n758 B.n757 83.1578
R1058 B.n757 B.n22 83.1578
R1059 B.n751 B.n22 83.1578
R1060 B.n751 B.n750 83.1578
R1061 B.n750 B.n749 83.1578
R1062 B.n749 B.n29 83.1578
R1063 B.n743 B.n742 83.1578
R1064 B.n742 B.n741 83.1578
R1065 B.n741 B.n36 83.1578
R1066 B.n735 B.n36 83.1578
R1067 B.n735 B.n734 83.1578
R1068 B.n734 B.n733 83.1578
R1069 B.n733 B.n43 83.1578
R1070 B.n727 B.n43 83.1578
R1071 B.n726 B.n725 83.1578
R1072 B.n725 B.n50 83.1578
R1073 B.n719 B.n50 83.1578
R1074 B.n719 B.n718 83.1578
R1075 B.n718 B.n717 83.1578
R1076 B.n717 B.n57 83.1578
R1077 B.n711 B.n57 83.1578
R1078 B.n711 B.n710 83.1578
R1079 B.n709 B.n64 83.1578
R1080 B.n703 B.n64 83.1578
R1081 B.n703 B.n702 83.1578
R1082 B.n702 B.n701 83.1578
R1083 B.n701 B.n71 83.1578
R1084 B.n695 B.n71 83.1578
R1085 B.n695 B.n694 83.1578
R1086 B.n694 B.n693 83.1578
R1087 B.n693 B.n78 83.1578
R1088 B.n687 B.n78 83.1578
R1089 B.n687 B.n686 83.1578
R1090 B.n686 B.n685 83.1578
R1091 B.n679 B.n88 83.1578
R1092 B.n679 B.n678 83.1578
R1093 B.n678 B.n677 83.1578
R1094 B.n677 B.n92 83.1578
R1095 B.n671 B.n92 83.1578
R1096 B.n671 B.n670 83.1578
R1097 B.n670 B.n669 83.1578
R1098 B.n250 B.t20 78.6841
R1099 B.n118 B.t15 78.6841
R1100 B.n242 B.t10 78.6812
R1101 B.n110 B.t18 78.6812
R1102 B.n365 B.t9 74.5975
R1103 B.n88 B.t13 74.5975
R1104 B.n341 B.n232 71.676
R1105 B.n339 B.n234 71.676
R1106 B.n335 B.n334 71.676
R1107 B.n328 B.n236 71.676
R1108 B.n327 B.n326 71.676
R1109 B.n320 B.n238 71.676
R1110 B.n319 B.n318 71.676
R1111 B.n312 B.n240 71.676
R1112 B.n311 B.n244 71.676
R1113 B.n307 B.n306 71.676
R1114 B.n300 B.n246 71.676
R1115 B.n299 B.n298 71.676
R1116 B.n292 B.n248 71.676
R1117 B.n291 B.n252 71.676
R1118 B.n287 B.n286 71.676
R1119 B.n280 B.n254 71.676
R1120 B.n279 B.n278 71.676
R1121 B.n272 B.n256 71.676
R1122 B.n271 B.n270 71.676
R1123 B.n264 B.n258 71.676
R1124 B.n263 B.n262 71.676
R1125 B.n663 B.n100 71.676
R1126 B.n662 B.n661 71.676
R1127 B.n655 B.n102 71.676
R1128 B.n654 B.n653 71.676
R1129 B.n647 B.n104 71.676
R1130 B.n646 B.n645 71.676
R1131 B.n639 B.n106 71.676
R1132 B.n638 B.n637 71.676
R1133 B.n630 B.n108 71.676
R1134 B.n629 B.n628 71.676
R1135 B.n622 B.n112 71.676
R1136 B.n621 B.n620 71.676
R1137 B.n614 B.n114 71.676
R1138 B.n613 B.n612 71.676
R1139 B.n606 B.n116 71.676
R1140 B.n605 B.n604 71.676
R1141 B.n598 B.n121 71.676
R1142 B.n597 B.n596 71.676
R1143 B.n590 B.n123 71.676
R1144 B.n589 B.n588 71.676
R1145 B.n582 B.n125 71.676
R1146 B.n581 B.n580 71.676
R1147 B.n580 B.n579 71.676
R1148 B.n583 B.n582 71.676
R1149 B.n588 B.n587 71.676
R1150 B.n591 B.n590 71.676
R1151 B.n596 B.n595 71.676
R1152 B.n599 B.n598 71.676
R1153 B.n604 B.n603 71.676
R1154 B.n607 B.n606 71.676
R1155 B.n612 B.n611 71.676
R1156 B.n615 B.n614 71.676
R1157 B.n620 B.n619 71.676
R1158 B.n623 B.n622 71.676
R1159 B.n628 B.n627 71.676
R1160 B.n631 B.n630 71.676
R1161 B.n637 B.n636 71.676
R1162 B.n640 B.n639 71.676
R1163 B.n645 B.n644 71.676
R1164 B.n648 B.n647 71.676
R1165 B.n653 B.n652 71.676
R1166 B.n656 B.n655 71.676
R1167 B.n661 B.n660 71.676
R1168 B.n664 B.n663 71.676
R1169 B.n342 B.n341 71.676
R1170 B.n336 B.n234 71.676
R1171 B.n334 B.n333 71.676
R1172 B.n329 B.n328 71.676
R1173 B.n326 B.n325 71.676
R1174 B.n321 B.n320 71.676
R1175 B.n318 B.n317 71.676
R1176 B.n313 B.n312 71.676
R1177 B.n308 B.n244 71.676
R1178 B.n306 B.n305 71.676
R1179 B.n301 B.n300 71.676
R1180 B.n298 B.n297 71.676
R1181 B.n293 B.n292 71.676
R1182 B.n288 B.n252 71.676
R1183 B.n286 B.n285 71.676
R1184 B.n281 B.n280 71.676
R1185 B.n278 B.n277 71.676
R1186 B.n273 B.n272 71.676
R1187 B.n270 B.n269 71.676
R1188 B.n265 B.n264 71.676
R1189 B.n262 B.n261 71.676
R1190 B.n486 B.t3 67.2601
R1191 B.n18 B.t5 67.2601
R1192 B.n250 B.n249 60.5096
R1193 B.n242 B.n241 60.5096
R1194 B.n110 B.n109 60.5096
R1195 B.n118 B.n117 60.5096
R1196 B.t1 B.n188 59.9227
R1197 B.n710 B.t4 59.9227
R1198 B.n251 B.n250 59.5399
R1199 B.n243 B.n242 59.5399
R1200 B.n633 B.n110 59.5399
R1201 B.n119 B.n118 59.5399
R1202 B.n462 B.t7 52.5853
R1203 B.n743 B.t0 52.5853
R1204 B.n438 B.t2 45.2479
R1205 B.n727 B.t6 45.2479
R1206 B.n176 B.t2 37.9105
R1207 B.t6 B.n726 37.9105
R1208 B.n667 B.n666 32.9371
R1209 B.n578 B.n577 32.9371
R1210 B.n349 B.n229 32.9371
R1211 B.n345 B.n344 32.9371
R1212 B.t7 B.n152 30.573
R1213 B.t0 B.n29 30.573
R1214 B.n408 B.t1 23.2356
R1215 B.t4 B.n709 23.2356
R1216 B B.n777 18.0485
R1217 B.n493 B.t3 15.8982
R1218 B.n765 B.t5 15.8982
R1219 B.n666 B.n665 10.6151
R1220 B.n665 B.n101 10.6151
R1221 B.n659 B.n101 10.6151
R1222 B.n659 B.n658 10.6151
R1223 B.n658 B.n657 10.6151
R1224 B.n657 B.n103 10.6151
R1225 B.n651 B.n103 10.6151
R1226 B.n651 B.n650 10.6151
R1227 B.n650 B.n649 10.6151
R1228 B.n649 B.n105 10.6151
R1229 B.n643 B.n105 10.6151
R1230 B.n643 B.n642 10.6151
R1231 B.n642 B.n641 10.6151
R1232 B.n641 B.n107 10.6151
R1233 B.n635 B.n107 10.6151
R1234 B.n635 B.n634 10.6151
R1235 B.n632 B.n111 10.6151
R1236 B.n626 B.n111 10.6151
R1237 B.n626 B.n625 10.6151
R1238 B.n625 B.n624 10.6151
R1239 B.n624 B.n113 10.6151
R1240 B.n618 B.n113 10.6151
R1241 B.n618 B.n617 10.6151
R1242 B.n617 B.n616 10.6151
R1243 B.n616 B.n115 10.6151
R1244 B.n610 B.n609 10.6151
R1245 B.n609 B.n608 10.6151
R1246 B.n608 B.n120 10.6151
R1247 B.n602 B.n120 10.6151
R1248 B.n602 B.n601 10.6151
R1249 B.n601 B.n600 10.6151
R1250 B.n600 B.n122 10.6151
R1251 B.n594 B.n122 10.6151
R1252 B.n594 B.n593 10.6151
R1253 B.n593 B.n592 10.6151
R1254 B.n592 B.n124 10.6151
R1255 B.n586 B.n124 10.6151
R1256 B.n586 B.n585 10.6151
R1257 B.n585 B.n584 10.6151
R1258 B.n584 B.n126 10.6151
R1259 B.n578 B.n126 10.6151
R1260 B.n350 B.n349 10.6151
R1261 B.n351 B.n350 10.6151
R1262 B.n351 B.n221 10.6151
R1263 B.n361 B.n221 10.6151
R1264 B.n362 B.n361 10.6151
R1265 B.n363 B.n362 10.6151
R1266 B.n363 B.n214 10.6151
R1267 B.n374 B.n214 10.6151
R1268 B.n375 B.n374 10.6151
R1269 B.n376 B.n375 10.6151
R1270 B.n376 B.n206 10.6151
R1271 B.n386 B.n206 10.6151
R1272 B.n387 B.n386 10.6151
R1273 B.n388 B.n387 10.6151
R1274 B.n388 B.n198 10.6151
R1275 B.n398 B.n198 10.6151
R1276 B.n399 B.n398 10.6151
R1277 B.n400 B.n399 10.6151
R1278 B.n400 B.n190 10.6151
R1279 B.n410 B.n190 10.6151
R1280 B.n411 B.n410 10.6151
R1281 B.n412 B.n411 10.6151
R1282 B.n412 B.n182 10.6151
R1283 B.n422 B.n182 10.6151
R1284 B.n423 B.n422 10.6151
R1285 B.n424 B.n423 10.6151
R1286 B.n424 B.n173 10.6151
R1287 B.n434 B.n173 10.6151
R1288 B.n435 B.n434 10.6151
R1289 B.n436 B.n435 10.6151
R1290 B.n436 B.n166 10.6151
R1291 B.n446 B.n166 10.6151
R1292 B.n447 B.n446 10.6151
R1293 B.n448 B.n447 10.6151
R1294 B.n448 B.n158 10.6151
R1295 B.n458 B.n158 10.6151
R1296 B.n459 B.n458 10.6151
R1297 B.n460 B.n459 10.6151
R1298 B.n460 B.n150 10.6151
R1299 B.n470 B.n150 10.6151
R1300 B.n471 B.n470 10.6151
R1301 B.n472 B.n471 10.6151
R1302 B.n472 B.n142 10.6151
R1303 B.n482 B.n142 10.6151
R1304 B.n483 B.n482 10.6151
R1305 B.n484 B.n483 10.6151
R1306 B.n484 B.n135 10.6151
R1307 B.n495 B.n135 10.6151
R1308 B.n496 B.n495 10.6151
R1309 B.n498 B.n496 10.6151
R1310 B.n498 B.n497 10.6151
R1311 B.n497 B.n127 10.6151
R1312 B.n509 B.n127 10.6151
R1313 B.n510 B.n509 10.6151
R1314 B.n511 B.n510 10.6151
R1315 B.n512 B.n511 10.6151
R1316 B.n514 B.n512 10.6151
R1317 B.n515 B.n514 10.6151
R1318 B.n516 B.n515 10.6151
R1319 B.n517 B.n516 10.6151
R1320 B.n519 B.n517 10.6151
R1321 B.n520 B.n519 10.6151
R1322 B.n521 B.n520 10.6151
R1323 B.n522 B.n521 10.6151
R1324 B.n524 B.n522 10.6151
R1325 B.n525 B.n524 10.6151
R1326 B.n526 B.n525 10.6151
R1327 B.n527 B.n526 10.6151
R1328 B.n529 B.n527 10.6151
R1329 B.n530 B.n529 10.6151
R1330 B.n531 B.n530 10.6151
R1331 B.n532 B.n531 10.6151
R1332 B.n534 B.n532 10.6151
R1333 B.n535 B.n534 10.6151
R1334 B.n536 B.n535 10.6151
R1335 B.n537 B.n536 10.6151
R1336 B.n539 B.n537 10.6151
R1337 B.n540 B.n539 10.6151
R1338 B.n541 B.n540 10.6151
R1339 B.n542 B.n541 10.6151
R1340 B.n544 B.n542 10.6151
R1341 B.n545 B.n544 10.6151
R1342 B.n546 B.n545 10.6151
R1343 B.n547 B.n546 10.6151
R1344 B.n549 B.n547 10.6151
R1345 B.n550 B.n549 10.6151
R1346 B.n551 B.n550 10.6151
R1347 B.n552 B.n551 10.6151
R1348 B.n554 B.n552 10.6151
R1349 B.n555 B.n554 10.6151
R1350 B.n556 B.n555 10.6151
R1351 B.n557 B.n556 10.6151
R1352 B.n559 B.n557 10.6151
R1353 B.n560 B.n559 10.6151
R1354 B.n561 B.n560 10.6151
R1355 B.n562 B.n561 10.6151
R1356 B.n564 B.n562 10.6151
R1357 B.n565 B.n564 10.6151
R1358 B.n566 B.n565 10.6151
R1359 B.n567 B.n566 10.6151
R1360 B.n569 B.n567 10.6151
R1361 B.n570 B.n569 10.6151
R1362 B.n571 B.n570 10.6151
R1363 B.n572 B.n571 10.6151
R1364 B.n574 B.n572 10.6151
R1365 B.n575 B.n574 10.6151
R1366 B.n576 B.n575 10.6151
R1367 B.n577 B.n576 10.6151
R1368 B.n344 B.n343 10.6151
R1369 B.n343 B.n233 10.6151
R1370 B.n338 B.n233 10.6151
R1371 B.n338 B.n337 10.6151
R1372 B.n337 B.n235 10.6151
R1373 B.n332 B.n235 10.6151
R1374 B.n332 B.n331 10.6151
R1375 B.n331 B.n330 10.6151
R1376 B.n330 B.n237 10.6151
R1377 B.n324 B.n237 10.6151
R1378 B.n324 B.n323 10.6151
R1379 B.n323 B.n322 10.6151
R1380 B.n322 B.n239 10.6151
R1381 B.n316 B.n239 10.6151
R1382 B.n316 B.n315 10.6151
R1383 B.n315 B.n314 10.6151
R1384 B.n310 B.n309 10.6151
R1385 B.n309 B.n245 10.6151
R1386 B.n304 B.n245 10.6151
R1387 B.n304 B.n303 10.6151
R1388 B.n303 B.n302 10.6151
R1389 B.n302 B.n247 10.6151
R1390 B.n296 B.n247 10.6151
R1391 B.n296 B.n295 10.6151
R1392 B.n295 B.n294 10.6151
R1393 B.n290 B.n289 10.6151
R1394 B.n289 B.n253 10.6151
R1395 B.n284 B.n253 10.6151
R1396 B.n284 B.n283 10.6151
R1397 B.n283 B.n282 10.6151
R1398 B.n282 B.n255 10.6151
R1399 B.n276 B.n255 10.6151
R1400 B.n276 B.n275 10.6151
R1401 B.n275 B.n274 10.6151
R1402 B.n274 B.n257 10.6151
R1403 B.n268 B.n257 10.6151
R1404 B.n268 B.n267 10.6151
R1405 B.n267 B.n266 10.6151
R1406 B.n266 B.n259 10.6151
R1407 B.n260 B.n259 10.6151
R1408 B.n260 B.n229 10.6151
R1409 B.n345 B.n225 10.6151
R1410 B.n355 B.n225 10.6151
R1411 B.n356 B.n355 10.6151
R1412 B.n357 B.n356 10.6151
R1413 B.n357 B.n217 10.6151
R1414 B.n368 B.n217 10.6151
R1415 B.n369 B.n368 10.6151
R1416 B.n370 B.n369 10.6151
R1417 B.n370 B.n210 10.6151
R1418 B.n380 B.n210 10.6151
R1419 B.n381 B.n380 10.6151
R1420 B.n382 B.n381 10.6151
R1421 B.n382 B.n202 10.6151
R1422 B.n392 B.n202 10.6151
R1423 B.n393 B.n392 10.6151
R1424 B.n394 B.n393 10.6151
R1425 B.n394 B.n194 10.6151
R1426 B.n404 B.n194 10.6151
R1427 B.n405 B.n404 10.6151
R1428 B.n406 B.n405 10.6151
R1429 B.n406 B.n186 10.6151
R1430 B.n416 B.n186 10.6151
R1431 B.n417 B.n416 10.6151
R1432 B.n418 B.n417 10.6151
R1433 B.n418 B.n178 10.6151
R1434 B.n428 B.n178 10.6151
R1435 B.n429 B.n428 10.6151
R1436 B.n430 B.n429 10.6151
R1437 B.n430 B.n170 10.6151
R1438 B.n440 B.n170 10.6151
R1439 B.n441 B.n440 10.6151
R1440 B.n442 B.n441 10.6151
R1441 B.n442 B.n162 10.6151
R1442 B.n452 B.n162 10.6151
R1443 B.n453 B.n452 10.6151
R1444 B.n454 B.n453 10.6151
R1445 B.n454 B.n154 10.6151
R1446 B.n464 B.n154 10.6151
R1447 B.n465 B.n464 10.6151
R1448 B.n466 B.n465 10.6151
R1449 B.n466 B.n146 10.6151
R1450 B.n476 B.n146 10.6151
R1451 B.n477 B.n476 10.6151
R1452 B.n478 B.n477 10.6151
R1453 B.n478 B.n138 10.6151
R1454 B.n489 B.n138 10.6151
R1455 B.n490 B.n489 10.6151
R1456 B.n491 B.n490 10.6151
R1457 B.n491 B.n131 10.6151
R1458 B.n502 B.n131 10.6151
R1459 B.n503 B.n502 10.6151
R1460 B.n504 B.n503 10.6151
R1461 B.n504 B.n0 10.6151
R1462 B.n771 B.n1 10.6151
R1463 B.n771 B.n770 10.6151
R1464 B.n770 B.n769 10.6151
R1465 B.n769 B.n10 10.6151
R1466 B.n763 B.n10 10.6151
R1467 B.n763 B.n762 10.6151
R1468 B.n762 B.n761 10.6151
R1469 B.n761 B.n16 10.6151
R1470 B.n755 B.n16 10.6151
R1471 B.n755 B.n754 10.6151
R1472 B.n754 B.n753 10.6151
R1473 B.n753 B.n24 10.6151
R1474 B.n747 B.n24 10.6151
R1475 B.n747 B.n746 10.6151
R1476 B.n746 B.n745 10.6151
R1477 B.n745 B.n31 10.6151
R1478 B.n739 B.n31 10.6151
R1479 B.n739 B.n738 10.6151
R1480 B.n738 B.n737 10.6151
R1481 B.n737 B.n38 10.6151
R1482 B.n731 B.n38 10.6151
R1483 B.n731 B.n730 10.6151
R1484 B.n730 B.n729 10.6151
R1485 B.n729 B.n45 10.6151
R1486 B.n723 B.n45 10.6151
R1487 B.n723 B.n722 10.6151
R1488 B.n722 B.n721 10.6151
R1489 B.n721 B.n52 10.6151
R1490 B.n715 B.n52 10.6151
R1491 B.n715 B.n714 10.6151
R1492 B.n714 B.n713 10.6151
R1493 B.n713 B.n59 10.6151
R1494 B.n707 B.n59 10.6151
R1495 B.n707 B.n706 10.6151
R1496 B.n706 B.n705 10.6151
R1497 B.n705 B.n66 10.6151
R1498 B.n699 B.n66 10.6151
R1499 B.n699 B.n698 10.6151
R1500 B.n698 B.n697 10.6151
R1501 B.n697 B.n73 10.6151
R1502 B.n691 B.n73 10.6151
R1503 B.n691 B.n690 10.6151
R1504 B.n690 B.n689 10.6151
R1505 B.n689 B.n80 10.6151
R1506 B.n683 B.n80 10.6151
R1507 B.n683 B.n682 10.6151
R1508 B.n682 B.n681 10.6151
R1509 B.n681 B.n86 10.6151
R1510 B.n675 B.n86 10.6151
R1511 B.n675 B.n674 10.6151
R1512 B.n674 B.n673 10.6151
R1513 B.n673 B.n94 10.6151
R1514 B.n667 B.n94 10.6151
R1515 B.n634 B.n633 9.52245
R1516 B.n610 B.n119 9.52245
R1517 B.n314 B.n243 9.52245
R1518 B.n290 B.n251 9.52245
R1519 B.n372 B.t9 8.56081
R1520 B.n685 B.t13 8.56081
R1521 B.n777 B.n0 2.81026
R1522 B.n777 B.n1 2.81026
R1523 B.n633 B.n632 1.09318
R1524 B.n119 B.n115 1.09318
R1525 B.n310 B.n243 1.09318
R1526 B.n294 B.n251 1.09318
R1527 VN.n56 VN.n55 161.3
R1528 VN.n54 VN.n30 161.3
R1529 VN.n53 VN.n52 161.3
R1530 VN.n51 VN.n31 161.3
R1531 VN.n50 VN.n49 161.3
R1532 VN.n48 VN.n32 161.3
R1533 VN.n46 VN.n45 161.3
R1534 VN.n44 VN.n33 161.3
R1535 VN.n43 VN.n42 161.3
R1536 VN.n41 VN.n34 161.3
R1537 VN.n40 VN.n39 161.3
R1538 VN.n38 VN.n35 161.3
R1539 VN.n27 VN.n26 161.3
R1540 VN.n25 VN.n1 161.3
R1541 VN.n24 VN.n23 161.3
R1542 VN.n22 VN.n2 161.3
R1543 VN.n21 VN.n20 161.3
R1544 VN.n19 VN.n3 161.3
R1545 VN.n17 VN.n16 161.3
R1546 VN.n15 VN.n4 161.3
R1547 VN.n14 VN.n13 161.3
R1548 VN.n12 VN.n5 161.3
R1549 VN.n11 VN.n10 161.3
R1550 VN.n9 VN.n6 161.3
R1551 VN.n28 VN.n0 68.9556
R1552 VN.n57 VN.n29 68.9556
R1553 VN.n37 VN.t6 63.896
R1554 VN.n8 VN.t5 63.896
R1555 VN.n8 VN.n7 58.3046
R1556 VN.n37 VN.n36 58.3046
R1557 VN.n13 VN.n12 56.4773
R1558 VN.n42 VN.n41 56.4773
R1559 VN.n24 VN.n2 53.0692
R1560 VN.n53 VN.n31 53.0692
R1561 VN VN.n57 45.7631
R1562 VN.n7 VN.t2 32.1338
R1563 VN.n18 VN.t1 32.1338
R1564 VN.n0 VN.t4 32.1338
R1565 VN.n36 VN.t0 32.1338
R1566 VN.n47 VN.t3 32.1338
R1567 VN.n29 VN.t7 32.1338
R1568 VN.n25 VN.n24 27.752
R1569 VN.n54 VN.n53 27.752
R1570 VN.n11 VN.n6 24.3439
R1571 VN.n12 VN.n11 24.3439
R1572 VN.n13 VN.n4 24.3439
R1573 VN.n17 VN.n4 24.3439
R1574 VN.n20 VN.n19 24.3439
R1575 VN.n20 VN.n2 24.3439
R1576 VN.n26 VN.n25 24.3439
R1577 VN.n41 VN.n40 24.3439
R1578 VN.n40 VN.n35 24.3439
R1579 VN.n49 VN.n31 24.3439
R1580 VN.n49 VN.n48 24.3439
R1581 VN.n46 VN.n33 24.3439
R1582 VN.n42 VN.n33 24.3439
R1583 VN.n55 VN.n54 24.3439
R1584 VN.n26 VN.n0 20.9359
R1585 VN.n55 VN.n29 20.9359
R1586 VN.n7 VN.n6 15.0934
R1587 VN.n18 VN.n17 15.0934
R1588 VN.n36 VN.n35 15.0934
R1589 VN.n47 VN.n46 15.0934
R1590 VN.n19 VN.n18 9.251
R1591 VN.n48 VN.n47 9.251
R1592 VN.n38 VN.n37 5.48085
R1593 VN.n9 VN.n8 5.48085
R1594 VN.n57 VN.n56 0.355081
R1595 VN.n28 VN.n27 0.355081
R1596 VN VN.n28 0.26685
R1597 VN.n56 VN.n30 0.189894
R1598 VN.n52 VN.n30 0.189894
R1599 VN.n52 VN.n51 0.189894
R1600 VN.n51 VN.n50 0.189894
R1601 VN.n50 VN.n32 0.189894
R1602 VN.n45 VN.n32 0.189894
R1603 VN.n45 VN.n44 0.189894
R1604 VN.n44 VN.n43 0.189894
R1605 VN.n43 VN.n34 0.189894
R1606 VN.n39 VN.n34 0.189894
R1607 VN.n39 VN.n38 0.189894
R1608 VN.n10 VN.n9 0.189894
R1609 VN.n10 VN.n5 0.189894
R1610 VN.n14 VN.n5 0.189894
R1611 VN.n15 VN.n14 0.189894
R1612 VN.n16 VN.n15 0.189894
R1613 VN.n16 VN.n3 0.189894
R1614 VN.n21 VN.n3 0.189894
R1615 VN.n22 VN.n21 0.189894
R1616 VN.n23 VN.n22 0.189894
R1617 VN.n23 VN.n1 0.189894
R1618 VN.n27 VN.n1 0.189894
R1619 VDD2.n2 VDD2.n1 75.33
R1620 VDD2.n2 VDD2.n0 75.33
R1621 VDD2 VDD2.n5 75.3272
R1622 VDD2.n4 VDD2.n3 74.0406
R1623 VDD2.n4 VDD2.n2 39.0256
R1624 VDD2.n5 VDD2.t7 5.32308
R1625 VDD2.n5 VDD2.t1 5.32308
R1626 VDD2.n3 VDD2.t0 5.32308
R1627 VDD2.n3 VDD2.t4 5.32308
R1628 VDD2.n1 VDD2.t6 5.32308
R1629 VDD2.n1 VDD2.t3 5.32308
R1630 VDD2.n0 VDD2.t2 5.32308
R1631 VDD2.n0 VDD2.t5 5.32308
R1632 VDD2 VDD2.n4 1.40352
C0 VTAIL VN 4.10838f
C1 VDD1 VDD2 1.87613f
C2 VDD2 VP 0.544701f
C3 VDD1 VTAIL 5.4411f
C4 VTAIL VP 4.12249f
C5 VDD1 VN 0.156201f
C6 VN VP 6.37875f
C7 VTAIL VDD2 5.49679f
C8 VDD1 VP 3.43519f
C9 VN VDD2 3.04903f
C10 VDD2 B 4.871132f
C11 VDD1 B 5.33688f
C12 VTAIL B 5.223108f
C13 VN B 15.50414f
C14 VP B 14.076917f
C15 VDD2.t2 B 0.070626f
C16 VDD2.t5 B 0.070626f
C17 VDD2.n0 B 0.544669f
C18 VDD2.t6 B 0.070626f
C19 VDD2.t3 B 0.070626f
C20 VDD2.n1 B 0.544669f
C21 VDD2.n2 B 2.76969f
C22 VDD2.t0 B 0.070626f
C23 VDD2.t4 B 0.070626f
C24 VDD2.n3 B 0.535848f
C25 VDD2.n4 B 2.28124f
C26 VDD2.t7 B 0.070626f
C27 VDD2.t1 B 0.070626f
C28 VDD2.n5 B 0.544641f
C29 VN.t4 B 0.690848f
C30 VN.n0 B 0.376916f
C31 VN.n1 B 0.026141f
C32 VN.n2 B 0.046609f
C33 VN.n3 B 0.026141f
C34 VN.t1 B 0.690848f
C35 VN.n4 B 0.048964f
C36 VN.n5 B 0.026141f
C37 VN.n6 B 0.039778f
C38 VN.t2 B 0.690848f
C39 VN.n7 B 0.360976f
C40 VN.t5 B 0.912968f
C41 VN.n8 B 0.347535f
C42 VN.n9 B 0.275934f
C43 VN.n10 B 0.026141f
C44 VN.n11 B 0.048964f
C45 VN.n12 B 0.038327f
C46 VN.n13 B 0.038327f
C47 VN.n14 B 0.026141f
C48 VN.n15 B 0.026141f
C49 VN.n16 B 0.026141f
C50 VN.n17 B 0.039778f
C51 VN.n18 B 0.277623f
C52 VN.n19 B 0.033975f
C53 VN.n20 B 0.048964f
C54 VN.n21 B 0.026141f
C55 VN.n22 B 0.026141f
C56 VN.n23 B 0.026141f
C57 VN.n24 B 0.027492f
C58 VN.n25 B 0.051518f
C59 VN.n26 B 0.04558f
C60 VN.n27 B 0.042197f
C61 VN.n28 B 0.051465f
C62 VN.t7 B 0.690848f
C63 VN.n29 B 0.376916f
C64 VN.n30 B 0.026141f
C65 VN.n31 B 0.046609f
C66 VN.n32 B 0.026141f
C67 VN.t3 B 0.690848f
C68 VN.n33 B 0.048964f
C69 VN.n34 B 0.026141f
C70 VN.n35 B 0.039778f
C71 VN.t6 B 0.912968f
C72 VN.t0 B 0.690848f
C73 VN.n36 B 0.360976f
C74 VN.n37 B 0.347535f
C75 VN.n38 B 0.275934f
C76 VN.n39 B 0.026141f
C77 VN.n40 B 0.048964f
C78 VN.n41 B 0.038327f
C79 VN.n42 B 0.038327f
C80 VN.n43 B 0.026141f
C81 VN.n44 B 0.026141f
C82 VN.n45 B 0.026141f
C83 VN.n46 B 0.039778f
C84 VN.n47 B 0.277623f
C85 VN.n48 B 0.033975f
C86 VN.n49 B 0.048964f
C87 VN.n50 B 0.026141f
C88 VN.n51 B 0.026141f
C89 VN.n52 B 0.026141f
C90 VN.n53 B 0.027492f
C91 VN.n54 B 0.051518f
C92 VN.n55 B 0.04558f
C93 VN.n56 B 0.042197f
C94 VN.n57 B 1.29604f
C95 VTAIL.t10 B 0.078793f
C96 VTAIL.t11 B 0.078793f
C97 VTAIL.n0 B 0.535288f
C98 VTAIL.n1 B 0.483536f
C99 VTAIL.t14 B 0.69317f
C100 VTAIL.n2 B 0.576096f
C101 VTAIL.t3 B 0.69317f
C102 VTAIL.n3 B 0.576096f
C103 VTAIL.t2 B 0.078793f
C104 VTAIL.t7 B 0.078793f
C105 VTAIL.n4 B 0.535288f
C106 VTAIL.n5 B 0.710808f
C107 VTAIL.t1 B 0.69317f
C108 VTAIL.n6 B 1.40888f
C109 VTAIL.t8 B 0.693174f
C110 VTAIL.n7 B 1.40888f
C111 VTAIL.t12 B 0.078793f
C112 VTAIL.t13 B 0.078793f
C113 VTAIL.n8 B 0.535292f
C114 VTAIL.n9 B 0.710804f
C115 VTAIL.t9 B 0.693174f
C116 VTAIL.n10 B 0.576093f
C117 VTAIL.t5 B 0.693174f
C118 VTAIL.n11 B 0.576093f
C119 VTAIL.t0 B 0.078793f
C120 VTAIL.t6 B 0.078793f
C121 VTAIL.n12 B 0.535292f
C122 VTAIL.n13 B 0.710804f
C123 VTAIL.t4 B 0.693174f
C124 VTAIL.n14 B 1.40888f
C125 VTAIL.t15 B 0.69317f
C126 VTAIL.n15 B 1.40386f
C127 VDD1.t7 B 0.072364f
C128 VDD1.t2 B 0.072364f
C129 VDD1.n0 B 0.55901f
C130 VDD1.t4 B 0.072364f
C131 VDD1.t3 B 0.072364f
C132 VDD1.n1 B 0.558067f
C133 VDD1.t5 B 0.072364f
C134 VDD1.t6 B 0.072364f
C135 VDD1.n2 B 0.558067f
C136 VDD1.n3 B 2.88919f
C137 VDD1.t0 B 0.072364f
C138 VDD1.t1 B 0.072364f
C139 VDD1.n4 B 0.549029f
C140 VDD1.n5 B 2.36767f
C141 VP.t4 B 0.713259f
C142 VP.n0 B 0.389143f
C143 VP.n1 B 0.026989f
C144 VP.n2 B 0.048121f
C145 VP.n3 B 0.026989f
C146 VP.t0 B 0.713259f
C147 VP.n4 B 0.050553f
C148 VP.n5 B 0.026989f
C149 VP.n6 B 0.041068f
C150 VP.n7 B 0.026989f
C151 VP.n8 B 0.028384f
C152 VP.n9 B 0.043566f
C153 VP.t6 B 0.713259f
C154 VP.t3 B 0.713259f
C155 VP.n10 B 0.389143f
C156 VP.n11 B 0.026989f
C157 VP.n12 B 0.048121f
C158 VP.n13 B 0.026989f
C159 VP.t1 B 0.713259f
C160 VP.n14 B 0.050553f
C161 VP.n15 B 0.026989f
C162 VP.n16 B 0.041068f
C163 VP.t2 B 0.942583f
C164 VP.t7 B 0.713259f
C165 VP.n17 B 0.372686f
C166 VP.n18 B 0.35881f
C167 VP.n19 B 0.284886f
C168 VP.n20 B 0.026989f
C169 VP.n21 B 0.050553f
C170 VP.n22 B 0.03957f
C171 VP.n23 B 0.03957f
C172 VP.n24 B 0.026989f
C173 VP.n25 B 0.026989f
C174 VP.n26 B 0.026989f
C175 VP.n27 B 0.041068f
C176 VP.n28 B 0.286629f
C177 VP.n29 B 0.035078f
C178 VP.n30 B 0.050553f
C179 VP.n31 B 0.026989f
C180 VP.n32 B 0.026989f
C181 VP.n33 B 0.026989f
C182 VP.n34 B 0.028384f
C183 VP.n35 B 0.053189f
C184 VP.n36 B 0.047058f
C185 VP.n37 B 0.043566f
C186 VP.n38 B 1.32666f
C187 VP.n39 B 1.34787f
C188 VP.n40 B 0.389143f
C189 VP.n41 B 0.047058f
C190 VP.n42 B 0.053189f
C191 VP.n43 B 0.026989f
C192 VP.n44 B 0.026989f
C193 VP.n45 B 0.026989f
C194 VP.n46 B 0.048121f
C195 VP.n47 B 0.050553f
C196 VP.t5 B 0.713259f
C197 VP.n48 B 0.286629f
C198 VP.n49 B 0.035078f
C199 VP.n50 B 0.026989f
C200 VP.n51 B 0.026989f
C201 VP.n52 B 0.026989f
C202 VP.n53 B 0.050553f
C203 VP.n54 B 0.03957f
C204 VP.n55 B 0.03957f
C205 VP.n56 B 0.026989f
C206 VP.n57 B 0.026989f
C207 VP.n58 B 0.026989f
C208 VP.n59 B 0.041068f
C209 VP.n60 B 0.286629f
C210 VP.n61 B 0.035078f
C211 VP.n62 B 0.050553f
C212 VP.n63 B 0.026989f
C213 VP.n64 B 0.026989f
C214 VP.n65 B 0.026989f
C215 VP.n66 B 0.028384f
C216 VP.n67 B 0.053189f
C217 VP.n68 B 0.047058f
C218 VP.n69 B 0.043566f
C219 VP.n70 B 0.053135f
.ends

