* NGSPICE file created from diff_pair_sample_0982.ext - technology: sky130A

.subckt diff_pair_sample_0982 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VP.t0 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X1 VDD2.t9 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0.10725 ps=0.98 w=0.65 l=2.23
X2 VDD1.t2 VP.t1 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0.10725 ps=0.98 w=0.65 l=2.23
X3 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0 ps=0 w=0.65 l=2.23
X4 VDD2.t8 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X5 VTAIL.t19 VN.t2 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X6 VTAIL.t2 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0 ps=0 w=0.65 l=2.23
X8 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0 ps=0 w=0.65 l=2.23
X9 VDD1.t8 VP.t2 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0.10725 ps=0.98 w=0.65 l=2.23
X10 VDD2.t5 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.2535 ps=2.08 w=0.65 l=2.23
X11 VTAIL.t0 VN.t5 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X12 VTAIL.t18 VN.t6 VDD2.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0 ps=0 w=0.65 l=2.23
X14 VTAIL.t13 VP.t3 VDD1.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X15 VDD1.t3 VP.t4 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X16 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.2535 ps=2.08 w=0.65 l=2.23
X17 VDD1.t4 VP.t5 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.2535 ps=2.08 w=0.65 l=2.23
X18 VDD1.t6 VP.t6 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.2535 ps=2.08 w=0.65 l=2.23
X19 VTAIL.t9 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X20 VDD1.t9 VP.t8 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X21 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0.10725 ps=0.98 w=0.65 l=2.23
X22 VTAIL.t7 VP.t9 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
X23 VDD2.t0 VN.t9 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=2.23
R0 VP.n22 VP.n21 161.3
R1 VP.n23 VP.n18 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n17 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n31 VP.n15 161.3
R7 VP.n33 VP.n32 161.3
R8 VP.n34 VP.n14 161.3
R9 VP.n36 VP.n35 161.3
R10 VP.n38 VP.n13 161.3
R11 VP.n40 VP.n39 161.3
R12 VP.n41 VP.n12 161.3
R13 VP.n43 VP.n42 161.3
R14 VP.n44 VP.n11 161.3
R15 VP.n80 VP.n0 161.3
R16 VP.n79 VP.n78 161.3
R17 VP.n77 VP.n1 161.3
R18 VP.n76 VP.n75 161.3
R19 VP.n74 VP.n2 161.3
R20 VP.n72 VP.n71 161.3
R21 VP.n70 VP.n3 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n67 VP.n4 161.3
R24 VP.n66 VP.n65 161.3
R25 VP.n64 VP.n63 161.3
R26 VP.n62 VP.n6 161.3
R27 VP.n61 VP.n60 161.3
R28 VP.n59 VP.n7 161.3
R29 VP.n58 VP.n57 161.3
R30 VP.n55 VP.n8 161.3
R31 VP.n54 VP.n53 161.3
R32 VP.n52 VP.n9 161.3
R33 VP.n51 VP.n50 161.3
R34 VP.n49 VP.n10 161.3
R35 VP.n48 VP.n47 92.6509
R36 VP.n82 VP.n81 92.6509
R37 VP.n46 VP.n45 92.6509
R38 VP.n20 VP.n19 56.0043
R39 VP.n50 VP.n9 49.2348
R40 VP.n79 VP.n1 49.2348
R41 VP.n43 VP.n12 49.2348
R42 VP.n61 VP.n7 43.4072
R43 VP.n68 VP.n3 43.4072
R44 VP.n32 VP.n14 43.4072
R45 VP.n25 VP.n18 43.4072
R46 VP.n47 VP.n46 42.5602
R47 VP.n19 VP.t2 40.6547
R48 VP.n62 VP.n61 37.5796
R49 VP.n68 VP.n67 37.5796
R50 VP.n32 VP.n31 37.5796
R51 VP.n26 VP.n25 37.5796
R52 VP.n54 VP.n9 31.752
R53 VP.n75 VP.n1 31.752
R54 VP.n39 VP.n12 31.752
R55 VP.n50 VP.n49 24.4675
R56 VP.n55 VP.n54 24.4675
R57 VP.n57 VP.n7 24.4675
R58 VP.n63 VP.n62 24.4675
R59 VP.n67 VP.n66 24.4675
R60 VP.n72 VP.n3 24.4675
R61 VP.n75 VP.n74 24.4675
R62 VP.n80 VP.n79 24.4675
R63 VP.n44 VP.n43 24.4675
R64 VP.n36 VP.n14 24.4675
R65 VP.n39 VP.n38 24.4675
R66 VP.n27 VP.n26 24.4675
R67 VP.n31 VP.n30 24.4675
R68 VP.n21 VP.n18 24.4675
R69 VP.n49 VP.n48 18.1061
R70 VP.n81 VP.n80 18.1061
R71 VP.n45 VP.n44 18.1061
R72 VP.n57 VP.n56 15.17
R73 VP.n73 VP.n72 15.17
R74 VP.n37 VP.n36 15.17
R75 VP.n21 VP.n20 15.17
R76 VP.n63 VP.n5 12.234
R77 VP.n66 VP.n5 12.234
R78 VP.n27 VP.n16 12.234
R79 VP.n30 VP.n16 12.234
R80 VP.n56 VP.n55 9.29796
R81 VP.n74 VP.n73 9.29796
R82 VP.n38 VP.n37 9.29796
R83 VP.n22 VP.n19 9.14908
R84 VP.n48 VP.t1 7.02516
R85 VP.n56 VP.t3 7.02516
R86 VP.n5 VP.t4 7.02516
R87 VP.n73 VP.t7 7.02516
R88 VP.n81 VP.t6 7.02516
R89 VP.n45 VP.t5 7.02516
R90 VP.n37 VP.t0 7.02516
R91 VP.n16 VP.t8 7.02516
R92 VP.n20 VP.t9 7.02516
R93 VP.n46 VP.n11 0.278367
R94 VP.n47 VP.n10 0.278367
R95 VP.n82 VP.n0 0.278367
R96 VP.n23 VP.n22 0.189894
R97 VP.n24 VP.n23 0.189894
R98 VP.n24 VP.n17 0.189894
R99 VP.n28 VP.n17 0.189894
R100 VP.n29 VP.n28 0.189894
R101 VP.n29 VP.n15 0.189894
R102 VP.n33 VP.n15 0.189894
R103 VP.n34 VP.n33 0.189894
R104 VP.n35 VP.n34 0.189894
R105 VP.n35 VP.n13 0.189894
R106 VP.n40 VP.n13 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n11 0.189894
R110 VP.n51 VP.n10 0.189894
R111 VP.n52 VP.n51 0.189894
R112 VP.n53 VP.n52 0.189894
R113 VP.n53 VP.n8 0.189894
R114 VP.n58 VP.n8 0.189894
R115 VP.n59 VP.n58 0.189894
R116 VP.n60 VP.n59 0.189894
R117 VP.n60 VP.n6 0.189894
R118 VP.n64 VP.n6 0.189894
R119 VP.n65 VP.n64 0.189894
R120 VP.n65 VP.n4 0.189894
R121 VP.n69 VP.n4 0.189894
R122 VP.n70 VP.n69 0.189894
R123 VP.n71 VP.n70 0.189894
R124 VP.n71 VP.n2 0.189894
R125 VP.n76 VP.n2 0.189894
R126 VP.n77 VP.n76 0.189894
R127 VP.n78 VP.n77 0.189894
R128 VP.n78 VP.n0 0.189894
R129 VP VP.n82 0.153454
R130 VDD1.n1 VDD1.t8 267.502
R131 VDD1.n3 VDD1.t2 267.502
R132 VDD1.n5 VDD1.n4 236.434
R133 VDD1.n7 VDD1.n6 234.833
R134 VDD1.n1 VDD1.n0 234.833
R135 VDD1.n3 VDD1.n2 234.833
R136 VDD1.n7 VDD1.n5 36.4449
R137 VDD1.n6 VDD1.t7 30.462
R138 VDD1.n6 VDD1.t4 30.462
R139 VDD1.n0 VDD1.t5 30.462
R140 VDD1.n0 VDD1.t9 30.462
R141 VDD1.n4 VDD1.t0 30.462
R142 VDD1.n4 VDD1.t6 30.462
R143 VDD1.n2 VDD1.t1 30.462
R144 VDD1.n2 VDD1.t3 30.462
R145 VDD1 VDD1.n7 1.59748
R146 VDD1 VDD1.n1 0.610414
R147 VDD1.n5 VDD1.n3 0.496878
R148 VTAIL.n17 VTAIL.t1 248.617
R149 VTAIL.n2 VTAIL.t10 248.617
R150 VTAIL.n16 VTAIL.t11 248.617
R151 VTAIL.n11 VTAIL.t6 248.617
R152 VTAIL.n19 VTAIL.n18 218.155
R153 VTAIL.n1 VTAIL.n0 218.155
R154 VTAIL.n4 VTAIL.n3 218.155
R155 VTAIL.n6 VTAIL.n5 218.155
R156 VTAIL.n15 VTAIL.n14 218.155
R157 VTAIL.n13 VTAIL.n12 218.155
R158 VTAIL.n10 VTAIL.n9 218.155
R159 VTAIL.n8 VTAIL.n7 218.155
R160 VTAIL.n18 VTAIL.t3 30.462
R161 VTAIL.n18 VTAIL.t0 30.462
R162 VTAIL.n0 VTAIL.t4 30.462
R163 VTAIL.n0 VTAIL.t19 30.462
R164 VTAIL.n3 VTAIL.t12 30.462
R165 VTAIL.n3 VTAIL.t9 30.462
R166 VTAIL.n5 VTAIL.t15 30.462
R167 VTAIL.n5 VTAIL.t13 30.462
R168 VTAIL.n14 VTAIL.t8 30.462
R169 VTAIL.n14 VTAIL.t16 30.462
R170 VTAIL.n12 VTAIL.t14 30.462
R171 VTAIL.n12 VTAIL.t7 30.462
R172 VTAIL.n9 VTAIL.t17 30.462
R173 VTAIL.n9 VTAIL.t2 30.462
R174 VTAIL.n7 VTAIL.t5 30.462
R175 VTAIL.n7 VTAIL.t18 30.462
R176 VTAIL.n8 VTAIL.n6 17.341
R177 VTAIL.n17 VTAIL.n16 15.1341
R178 VTAIL.n10 VTAIL.n8 2.2074
R179 VTAIL.n11 VTAIL.n10 2.2074
R180 VTAIL.n15 VTAIL.n13 2.2074
R181 VTAIL.n16 VTAIL.n15 2.2074
R182 VTAIL.n6 VTAIL.n4 2.2074
R183 VTAIL.n4 VTAIL.n2 2.2074
R184 VTAIL.n19 VTAIL.n17 2.2074
R185 VTAIL VTAIL.n1 1.71386
R186 VTAIL.n13 VTAIL.n11 1.57378
R187 VTAIL.n2 VTAIL.n1 1.57378
R188 VTAIL VTAIL.n19 0.494034
R189 B.n570 B.n569 585
R190 B.n166 B.n111 585
R191 B.n165 B.n164 585
R192 B.n163 B.n162 585
R193 B.n161 B.n160 585
R194 B.n159 B.n158 585
R195 B.n157 B.n156 585
R196 B.n155 B.n154 585
R197 B.n153 B.n152 585
R198 B.n151 B.n150 585
R199 B.n149 B.n148 585
R200 B.n147 B.n146 585
R201 B.n145 B.n144 585
R202 B.n143 B.n142 585
R203 B.n141 B.n140 585
R204 B.n139 B.n138 585
R205 B.n137 B.n136 585
R206 B.n135 B.n134 585
R207 B.n133 B.n132 585
R208 B.n131 B.n130 585
R209 B.n129 B.n128 585
R210 B.n127 B.n126 585
R211 B.n125 B.n124 585
R212 B.n123 B.n122 585
R213 B.n121 B.n120 585
R214 B.n119 B.n118 585
R215 B.n568 B.n98 585
R216 B.n573 B.n98 585
R217 B.n567 B.n97 585
R218 B.n574 B.n97 585
R219 B.n566 B.n565 585
R220 B.n565 B.n93 585
R221 B.n564 B.n92 585
R222 B.n580 B.n92 585
R223 B.n563 B.n91 585
R224 B.n581 B.n91 585
R225 B.n562 B.n90 585
R226 B.n582 B.n90 585
R227 B.n561 B.n560 585
R228 B.n560 B.n86 585
R229 B.n559 B.n85 585
R230 B.n588 B.n85 585
R231 B.n558 B.n84 585
R232 B.n589 B.n84 585
R233 B.n557 B.n83 585
R234 B.n590 B.n83 585
R235 B.n556 B.n555 585
R236 B.n555 B.n79 585
R237 B.n554 B.n78 585
R238 B.n596 B.n78 585
R239 B.n553 B.n77 585
R240 B.n597 B.n77 585
R241 B.n552 B.n76 585
R242 B.n598 B.n76 585
R243 B.n551 B.n550 585
R244 B.n550 B.n72 585
R245 B.n549 B.n71 585
R246 B.n604 B.n71 585
R247 B.n548 B.n70 585
R248 B.n605 B.n70 585
R249 B.n547 B.n69 585
R250 B.n606 B.n69 585
R251 B.n546 B.n545 585
R252 B.n545 B.n68 585
R253 B.n544 B.n64 585
R254 B.n612 B.n64 585
R255 B.n543 B.n63 585
R256 B.n613 B.n63 585
R257 B.n542 B.n62 585
R258 B.n614 B.n62 585
R259 B.n541 B.n540 585
R260 B.n540 B.n58 585
R261 B.n539 B.n57 585
R262 B.n620 B.n57 585
R263 B.n538 B.n56 585
R264 B.n621 B.n56 585
R265 B.n537 B.n55 585
R266 B.n622 B.n55 585
R267 B.n536 B.n535 585
R268 B.n535 B.n51 585
R269 B.n534 B.n50 585
R270 B.n628 B.n50 585
R271 B.n533 B.n49 585
R272 B.n629 B.n49 585
R273 B.n532 B.n48 585
R274 B.n630 B.n48 585
R275 B.n531 B.n530 585
R276 B.n530 B.n44 585
R277 B.n529 B.n43 585
R278 B.n636 B.n43 585
R279 B.n528 B.n42 585
R280 B.n637 B.n42 585
R281 B.n527 B.n41 585
R282 B.n638 B.n41 585
R283 B.n526 B.n525 585
R284 B.n525 B.n37 585
R285 B.n524 B.n36 585
R286 B.n644 B.n36 585
R287 B.n523 B.n35 585
R288 B.n645 B.n35 585
R289 B.n522 B.n34 585
R290 B.n646 B.n34 585
R291 B.n521 B.n520 585
R292 B.n520 B.n30 585
R293 B.n519 B.n29 585
R294 B.n652 B.n29 585
R295 B.n518 B.n28 585
R296 B.n653 B.n28 585
R297 B.n517 B.n27 585
R298 B.n654 B.n27 585
R299 B.n516 B.n515 585
R300 B.n515 B.n23 585
R301 B.n514 B.n22 585
R302 B.n660 B.n22 585
R303 B.n513 B.n21 585
R304 B.n661 B.n21 585
R305 B.n512 B.n20 585
R306 B.n662 B.n20 585
R307 B.n511 B.n510 585
R308 B.n510 B.n16 585
R309 B.n509 B.n15 585
R310 B.n668 B.n15 585
R311 B.n508 B.n14 585
R312 B.n669 B.n14 585
R313 B.n507 B.n13 585
R314 B.n670 B.n13 585
R315 B.n506 B.n505 585
R316 B.n505 B.n12 585
R317 B.n504 B.n503 585
R318 B.n504 B.n8 585
R319 B.n502 B.n7 585
R320 B.n677 B.n7 585
R321 B.n501 B.n6 585
R322 B.n678 B.n6 585
R323 B.n500 B.n5 585
R324 B.n679 B.n5 585
R325 B.n499 B.n498 585
R326 B.n498 B.n4 585
R327 B.n497 B.n167 585
R328 B.n497 B.n496 585
R329 B.n487 B.n168 585
R330 B.n169 B.n168 585
R331 B.n489 B.n488 585
R332 B.n490 B.n489 585
R333 B.n486 B.n173 585
R334 B.n177 B.n173 585
R335 B.n485 B.n484 585
R336 B.n484 B.n483 585
R337 B.n175 B.n174 585
R338 B.n176 B.n175 585
R339 B.n476 B.n475 585
R340 B.n477 B.n476 585
R341 B.n474 B.n182 585
R342 B.n182 B.n181 585
R343 B.n473 B.n472 585
R344 B.n472 B.n471 585
R345 B.n184 B.n183 585
R346 B.n185 B.n184 585
R347 B.n464 B.n463 585
R348 B.n465 B.n464 585
R349 B.n462 B.n189 585
R350 B.n193 B.n189 585
R351 B.n461 B.n460 585
R352 B.n460 B.n459 585
R353 B.n191 B.n190 585
R354 B.n192 B.n191 585
R355 B.n452 B.n451 585
R356 B.n453 B.n452 585
R357 B.n450 B.n198 585
R358 B.n198 B.n197 585
R359 B.n449 B.n448 585
R360 B.n448 B.n447 585
R361 B.n200 B.n199 585
R362 B.n201 B.n200 585
R363 B.n440 B.n439 585
R364 B.n441 B.n440 585
R365 B.n438 B.n206 585
R366 B.n206 B.n205 585
R367 B.n437 B.n436 585
R368 B.n436 B.n435 585
R369 B.n208 B.n207 585
R370 B.n209 B.n208 585
R371 B.n428 B.n427 585
R372 B.n429 B.n428 585
R373 B.n426 B.n214 585
R374 B.n214 B.n213 585
R375 B.n425 B.n424 585
R376 B.n424 B.n423 585
R377 B.n216 B.n215 585
R378 B.n217 B.n216 585
R379 B.n416 B.n415 585
R380 B.n417 B.n416 585
R381 B.n414 B.n222 585
R382 B.n222 B.n221 585
R383 B.n413 B.n412 585
R384 B.n412 B.n411 585
R385 B.n224 B.n223 585
R386 B.n225 B.n224 585
R387 B.n404 B.n403 585
R388 B.n405 B.n404 585
R389 B.n402 B.n230 585
R390 B.n230 B.n229 585
R391 B.n401 B.n400 585
R392 B.n400 B.n399 585
R393 B.n232 B.n231 585
R394 B.n392 B.n232 585
R395 B.n391 B.n390 585
R396 B.n393 B.n391 585
R397 B.n389 B.n237 585
R398 B.n237 B.n236 585
R399 B.n388 B.n387 585
R400 B.n387 B.n386 585
R401 B.n239 B.n238 585
R402 B.n240 B.n239 585
R403 B.n379 B.n378 585
R404 B.n380 B.n379 585
R405 B.n377 B.n245 585
R406 B.n245 B.n244 585
R407 B.n376 B.n375 585
R408 B.n375 B.n374 585
R409 B.n247 B.n246 585
R410 B.n248 B.n247 585
R411 B.n367 B.n366 585
R412 B.n368 B.n367 585
R413 B.n365 B.n253 585
R414 B.n253 B.n252 585
R415 B.n364 B.n363 585
R416 B.n363 B.n362 585
R417 B.n255 B.n254 585
R418 B.n256 B.n255 585
R419 B.n355 B.n354 585
R420 B.n356 B.n355 585
R421 B.n353 B.n261 585
R422 B.n261 B.n260 585
R423 B.n352 B.n351 585
R424 B.n351 B.n350 585
R425 B.n263 B.n262 585
R426 B.n264 B.n263 585
R427 B.n343 B.n342 585
R428 B.n344 B.n343 585
R429 B.n341 B.n269 585
R430 B.n269 B.n268 585
R431 B.n336 B.n335 585
R432 B.n334 B.n284 585
R433 B.n333 B.n283 585
R434 B.n338 B.n283 585
R435 B.n332 B.n331 585
R436 B.n330 B.n329 585
R437 B.n328 B.n327 585
R438 B.n326 B.n325 585
R439 B.n324 B.n323 585
R440 B.n321 B.n320 585
R441 B.n319 B.n318 585
R442 B.n317 B.n316 585
R443 B.n315 B.n314 585
R444 B.n313 B.n312 585
R445 B.n311 B.n310 585
R446 B.n309 B.n308 585
R447 B.n307 B.n306 585
R448 B.n305 B.n304 585
R449 B.n303 B.n302 585
R450 B.n300 B.n299 585
R451 B.n298 B.n297 585
R452 B.n296 B.n295 585
R453 B.n294 B.n293 585
R454 B.n292 B.n291 585
R455 B.n290 B.n289 585
R456 B.n271 B.n270 585
R457 B.n340 B.n339 585
R458 B.n339 B.n338 585
R459 B.n267 B.n266 585
R460 B.n268 B.n267 585
R461 B.n346 B.n345 585
R462 B.n345 B.n344 585
R463 B.n347 B.n265 585
R464 B.n265 B.n264 585
R465 B.n349 B.n348 585
R466 B.n350 B.n349 585
R467 B.n259 B.n258 585
R468 B.n260 B.n259 585
R469 B.n358 B.n357 585
R470 B.n357 B.n356 585
R471 B.n359 B.n257 585
R472 B.n257 B.n256 585
R473 B.n361 B.n360 585
R474 B.n362 B.n361 585
R475 B.n251 B.n250 585
R476 B.n252 B.n251 585
R477 B.n370 B.n369 585
R478 B.n369 B.n368 585
R479 B.n371 B.n249 585
R480 B.n249 B.n248 585
R481 B.n373 B.n372 585
R482 B.n374 B.n373 585
R483 B.n243 B.n242 585
R484 B.n244 B.n243 585
R485 B.n382 B.n381 585
R486 B.n381 B.n380 585
R487 B.n383 B.n241 585
R488 B.n241 B.n240 585
R489 B.n385 B.n384 585
R490 B.n386 B.n385 585
R491 B.n235 B.n234 585
R492 B.n236 B.n235 585
R493 B.n395 B.n394 585
R494 B.n394 B.n393 585
R495 B.n396 B.n233 585
R496 B.n392 B.n233 585
R497 B.n398 B.n397 585
R498 B.n399 B.n398 585
R499 B.n228 B.n227 585
R500 B.n229 B.n228 585
R501 B.n407 B.n406 585
R502 B.n406 B.n405 585
R503 B.n408 B.n226 585
R504 B.n226 B.n225 585
R505 B.n410 B.n409 585
R506 B.n411 B.n410 585
R507 B.n220 B.n219 585
R508 B.n221 B.n220 585
R509 B.n419 B.n418 585
R510 B.n418 B.n417 585
R511 B.n420 B.n218 585
R512 B.n218 B.n217 585
R513 B.n422 B.n421 585
R514 B.n423 B.n422 585
R515 B.n212 B.n211 585
R516 B.n213 B.n212 585
R517 B.n431 B.n430 585
R518 B.n430 B.n429 585
R519 B.n432 B.n210 585
R520 B.n210 B.n209 585
R521 B.n434 B.n433 585
R522 B.n435 B.n434 585
R523 B.n204 B.n203 585
R524 B.n205 B.n204 585
R525 B.n443 B.n442 585
R526 B.n442 B.n441 585
R527 B.n444 B.n202 585
R528 B.n202 B.n201 585
R529 B.n446 B.n445 585
R530 B.n447 B.n446 585
R531 B.n196 B.n195 585
R532 B.n197 B.n196 585
R533 B.n455 B.n454 585
R534 B.n454 B.n453 585
R535 B.n456 B.n194 585
R536 B.n194 B.n192 585
R537 B.n458 B.n457 585
R538 B.n459 B.n458 585
R539 B.n188 B.n187 585
R540 B.n193 B.n188 585
R541 B.n467 B.n466 585
R542 B.n466 B.n465 585
R543 B.n468 B.n186 585
R544 B.n186 B.n185 585
R545 B.n470 B.n469 585
R546 B.n471 B.n470 585
R547 B.n180 B.n179 585
R548 B.n181 B.n180 585
R549 B.n479 B.n478 585
R550 B.n478 B.n477 585
R551 B.n480 B.n178 585
R552 B.n178 B.n176 585
R553 B.n482 B.n481 585
R554 B.n483 B.n482 585
R555 B.n172 B.n171 585
R556 B.n177 B.n172 585
R557 B.n492 B.n491 585
R558 B.n491 B.n490 585
R559 B.n493 B.n170 585
R560 B.n170 B.n169 585
R561 B.n495 B.n494 585
R562 B.n496 B.n495 585
R563 B.n3 B.n0 585
R564 B.n4 B.n3 585
R565 B.n676 B.n1 585
R566 B.n677 B.n676 585
R567 B.n675 B.n674 585
R568 B.n675 B.n8 585
R569 B.n673 B.n9 585
R570 B.n12 B.n9 585
R571 B.n672 B.n671 585
R572 B.n671 B.n670 585
R573 B.n11 B.n10 585
R574 B.n669 B.n11 585
R575 B.n667 B.n666 585
R576 B.n668 B.n667 585
R577 B.n665 B.n17 585
R578 B.n17 B.n16 585
R579 B.n664 B.n663 585
R580 B.n663 B.n662 585
R581 B.n19 B.n18 585
R582 B.n661 B.n19 585
R583 B.n659 B.n658 585
R584 B.n660 B.n659 585
R585 B.n657 B.n24 585
R586 B.n24 B.n23 585
R587 B.n656 B.n655 585
R588 B.n655 B.n654 585
R589 B.n26 B.n25 585
R590 B.n653 B.n26 585
R591 B.n651 B.n650 585
R592 B.n652 B.n651 585
R593 B.n649 B.n31 585
R594 B.n31 B.n30 585
R595 B.n648 B.n647 585
R596 B.n647 B.n646 585
R597 B.n33 B.n32 585
R598 B.n645 B.n33 585
R599 B.n643 B.n642 585
R600 B.n644 B.n643 585
R601 B.n641 B.n38 585
R602 B.n38 B.n37 585
R603 B.n640 B.n639 585
R604 B.n639 B.n638 585
R605 B.n40 B.n39 585
R606 B.n637 B.n40 585
R607 B.n635 B.n634 585
R608 B.n636 B.n635 585
R609 B.n633 B.n45 585
R610 B.n45 B.n44 585
R611 B.n632 B.n631 585
R612 B.n631 B.n630 585
R613 B.n47 B.n46 585
R614 B.n629 B.n47 585
R615 B.n627 B.n626 585
R616 B.n628 B.n627 585
R617 B.n625 B.n52 585
R618 B.n52 B.n51 585
R619 B.n624 B.n623 585
R620 B.n623 B.n622 585
R621 B.n54 B.n53 585
R622 B.n621 B.n54 585
R623 B.n619 B.n618 585
R624 B.n620 B.n619 585
R625 B.n617 B.n59 585
R626 B.n59 B.n58 585
R627 B.n616 B.n615 585
R628 B.n615 B.n614 585
R629 B.n61 B.n60 585
R630 B.n613 B.n61 585
R631 B.n611 B.n610 585
R632 B.n612 B.n611 585
R633 B.n609 B.n65 585
R634 B.n68 B.n65 585
R635 B.n608 B.n607 585
R636 B.n607 B.n606 585
R637 B.n67 B.n66 585
R638 B.n605 B.n67 585
R639 B.n603 B.n602 585
R640 B.n604 B.n603 585
R641 B.n601 B.n73 585
R642 B.n73 B.n72 585
R643 B.n600 B.n599 585
R644 B.n599 B.n598 585
R645 B.n75 B.n74 585
R646 B.n597 B.n75 585
R647 B.n595 B.n594 585
R648 B.n596 B.n595 585
R649 B.n593 B.n80 585
R650 B.n80 B.n79 585
R651 B.n592 B.n591 585
R652 B.n591 B.n590 585
R653 B.n82 B.n81 585
R654 B.n589 B.n82 585
R655 B.n587 B.n586 585
R656 B.n588 B.n587 585
R657 B.n585 B.n87 585
R658 B.n87 B.n86 585
R659 B.n584 B.n583 585
R660 B.n583 B.n582 585
R661 B.n89 B.n88 585
R662 B.n581 B.n89 585
R663 B.n579 B.n578 585
R664 B.n580 B.n579 585
R665 B.n577 B.n94 585
R666 B.n94 B.n93 585
R667 B.n576 B.n575 585
R668 B.n575 B.n574 585
R669 B.n96 B.n95 585
R670 B.n573 B.n96 585
R671 B.n680 B.n679 585
R672 B.n678 B.n2 585
R673 B.n118 B.n96 468.476
R674 B.n570 B.n98 468.476
R675 B.n339 B.n269 468.476
R676 B.n336 B.n267 468.476
R677 B.n115 B.t12 287.413
R678 B.n112 B.t22 287.413
R679 B.n287 B.t17 287.413
R680 B.n285 B.t20 287.413
R681 B.n572 B.n571 256.663
R682 B.n572 B.n110 256.663
R683 B.n572 B.n109 256.663
R684 B.n572 B.n108 256.663
R685 B.n572 B.n107 256.663
R686 B.n572 B.n106 256.663
R687 B.n572 B.n105 256.663
R688 B.n572 B.n104 256.663
R689 B.n572 B.n103 256.663
R690 B.n572 B.n102 256.663
R691 B.n572 B.n101 256.663
R692 B.n572 B.n100 256.663
R693 B.n572 B.n99 256.663
R694 B.n338 B.n337 256.663
R695 B.n338 B.n272 256.663
R696 B.n338 B.n273 256.663
R697 B.n338 B.n274 256.663
R698 B.n338 B.n275 256.663
R699 B.n338 B.n276 256.663
R700 B.n338 B.n277 256.663
R701 B.n338 B.n278 256.663
R702 B.n338 B.n279 256.663
R703 B.n338 B.n280 256.663
R704 B.n338 B.n281 256.663
R705 B.n338 B.n282 256.663
R706 B.n682 B.n681 256.663
R707 B.n116 B.t13 237.766
R708 B.n113 B.t23 237.766
R709 B.n288 B.t16 237.766
R710 B.n286 B.t19 237.766
R711 B.n115 B.t10 208.819
R712 B.n112 B.t21 208.819
R713 B.n287 B.t14 208.819
R714 B.n285 B.t18 208.819
R715 B.n338 B.n268 202.363
R716 B.n573 B.n572 202.363
R717 B.n122 B.n121 163.367
R718 B.n126 B.n125 163.367
R719 B.n130 B.n129 163.367
R720 B.n134 B.n133 163.367
R721 B.n138 B.n137 163.367
R722 B.n142 B.n141 163.367
R723 B.n146 B.n145 163.367
R724 B.n150 B.n149 163.367
R725 B.n154 B.n153 163.367
R726 B.n158 B.n157 163.367
R727 B.n162 B.n161 163.367
R728 B.n164 B.n111 163.367
R729 B.n343 B.n269 163.367
R730 B.n343 B.n263 163.367
R731 B.n351 B.n263 163.367
R732 B.n351 B.n261 163.367
R733 B.n355 B.n261 163.367
R734 B.n355 B.n255 163.367
R735 B.n363 B.n255 163.367
R736 B.n363 B.n253 163.367
R737 B.n367 B.n253 163.367
R738 B.n367 B.n247 163.367
R739 B.n375 B.n247 163.367
R740 B.n375 B.n245 163.367
R741 B.n379 B.n245 163.367
R742 B.n379 B.n239 163.367
R743 B.n387 B.n239 163.367
R744 B.n387 B.n237 163.367
R745 B.n391 B.n237 163.367
R746 B.n391 B.n232 163.367
R747 B.n400 B.n232 163.367
R748 B.n400 B.n230 163.367
R749 B.n404 B.n230 163.367
R750 B.n404 B.n224 163.367
R751 B.n412 B.n224 163.367
R752 B.n412 B.n222 163.367
R753 B.n416 B.n222 163.367
R754 B.n416 B.n216 163.367
R755 B.n424 B.n216 163.367
R756 B.n424 B.n214 163.367
R757 B.n428 B.n214 163.367
R758 B.n428 B.n208 163.367
R759 B.n436 B.n208 163.367
R760 B.n436 B.n206 163.367
R761 B.n440 B.n206 163.367
R762 B.n440 B.n200 163.367
R763 B.n448 B.n200 163.367
R764 B.n448 B.n198 163.367
R765 B.n452 B.n198 163.367
R766 B.n452 B.n191 163.367
R767 B.n460 B.n191 163.367
R768 B.n460 B.n189 163.367
R769 B.n464 B.n189 163.367
R770 B.n464 B.n184 163.367
R771 B.n472 B.n184 163.367
R772 B.n472 B.n182 163.367
R773 B.n476 B.n182 163.367
R774 B.n476 B.n175 163.367
R775 B.n484 B.n175 163.367
R776 B.n484 B.n173 163.367
R777 B.n489 B.n173 163.367
R778 B.n489 B.n168 163.367
R779 B.n497 B.n168 163.367
R780 B.n498 B.n497 163.367
R781 B.n498 B.n5 163.367
R782 B.n6 B.n5 163.367
R783 B.n7 B.n6 163.367
R784 B.n504 B.n7 163.367
R785 B.n505 B.n504 163.367
R786 B.n505 B.n13 163.367
R787 B.n14 B.n13 163.367
R788 B.n15 B.n14 163.367
R789 B.n510 B.n15 163.367
R790 B.n510 B.n20 163.367
R791 B.n21 B.n20 163.367
R792 B.n22 B.n21 163.367
R793 B.n515 B.n22 163.367
R794 B.n515 B.n27 163.367
R795 B.n28 B.n27 163.367
R796 B.n29 B.n28 163.367
R797 B.n520 B.n29 163.367
R798 B.n520 B.n34 163.367
R799 B.n35 B.n34 163.367
R800 B.n36 B.n35 163.367
R801 B.n525 B.n36 163.367
R802 B.n525 B.n41 163.367
R803 B.n42 B.n41 163.367
R804 B.n43 B.n42 163.367
R805 B.n530 B.n43 163.367
R806 B.n530 B.n48 163.367
R807 B.n49 B.n48 163.367
R808 B.n50 B.n49 163.367
R809 B.n535 B.n50 163.367
R810 B.n535 B.n55 163.367
R811 B.n56 B.n55 163.367
R812 B.n57 B.n56 163.367
R813 B.n540 B.n57 163.367
R814 B.n540 B.n62 163.367
R815 B.n63 B.n62 163.367
R816 B.n64 B.n63 163.367
R817 B.n545 B.n64 163.367
R818 B.n545 B.n69 163.367
R819 B.n70 B.n69 163.367
R820 B.n71 B.n70 163.367
R821 B.n550 B.n71 163.367
R822 B.n550 B.n76 163.367
R823 B.n77 B.n76 163.367
R824 B.n78 B.n77 163.367
R825 B.n555 B.n78 163.367
R826 B.n555 B.n83 163.367
R827 B.n84 B.n83 163.367
R828 B.n85 B.n84 163.367
R829 B.n560 B.n85 163.367
R830 B.n560 B.n90 163.367
R831 B.n91 B.n90 163.367
R832 B.n92 B.n91 163.367
R833 B.n565 B.n92 163.367
R834 B.n565 B.n97 163.367
R835 B.n98 B.n97 163.367
R836 B.n284 B.n283 163.367
R837 B.n331 B.n283 163.367
R838 B.n329 B.n328 163.367
R839 B.n325 B.n324 163.367
R840 B.n320 B.n319 163.367
R841 B.n316 B.n315 163.367
R842 B.n312 B.n311 163.367
R843 B.n308 B.n307 163.367
R844 B.n304 B.n303 163.367
R845 B.n299 B.n298 163.367
R846 B.n295 B.n294 163.367
R847 B.n291 B.n290 163.367
R848 B.n339 B.n271 163.367
R849 B.n345 B.n267 163.367
R850 B.n345 B.n265 163.367
R851 B.n349 B.n265 163.367
R852 B.n349 B.n259 163.367
R853 B.n357 B.n259 163.367
R854 B.n357 B.n257 163.367
R855 B.n361 B.n257 163.367
R856 B.n361 B.n251 163.367
R857 B.n369 B.n251 163.367
R858 B.n369 B.n249 163.367
R859 B.n373 B.n249 163.367
R860 B.n373 B.n243 163.367
R861 B.n381 B.n243 163.367
R862 B.n381 B.n241 163.367
R863 B.n385 B.n241 163.367
R864 B.n385 B.n235 163.367
R865 B.n394 B.n235 163.367
R866 B.n394 B.n233 163.367
R867 B.n398 B.n233 163.367
R868 B.n398 B.n228 163.367
R869 B.n406 B.n228 163.367
R870 B.n406 B.n226 163.367
R871 B.n410 B.n226 163.367
R872 B.n410 B.n220 163.367
R873 B.n418 B.n220 163.367
R874 B.n418 B.n218 163.367
R875 B.n422 B.n218 163.367
R876 B.n422 B.n212 163.367
R877 B.n430 B.n212 163.367
R878 B.n430 B.n210 163.367
R879 B.n434 B.n210 163.367
R880 B.n434 B.n204 163.367
R881 B.n442 B.n204 163.367
R882 B.n442 B.n202 163.367
R883 B.n446 B.n202 163.367
R884 B.n446 B.n196 163.367
R885 B.n454 B.n196 163.367
R886 B.n454 B.n194 163.367
R887 B.n458 B.n194 163.367
R888 B.n458 B.n188 163.367
R889 B.n466 B.n188 163.367
R890 B.n466 B.n186 163.367
R891 B.n470 B.n186 163.367
R892 B.n470 B.n180 163.367
R893 B.n478 B.n180 163.367
R894 B.n478 B.n178 163.367
R895 B.n482 B.n178 163.367
R896 B.n482 B.n172 163.367
R897 B.n491 B.n172 163.367
R898 B.n491 B.n170 163.367
R899 B.n495 B.n170 163.367
R900 B.n495 B.n3 163.367
R901 B.n680 B.n3 163.367
R902 B.n676 B.n2 163.367
R903 B.n676 B.n675 163.367
R904 B.n675 B.n9 163.367
R905 B.n671 B.n9 163.367
R906 B.n671 B.n11 163.367
R907 B.n667 B.n11 163.367
R908 B.n667 B.n17 163.367
R909 B.n663 B.n17 163.367
R910 B.n663 B.n19 163.367
R911 B.n659 B.n19 163.367
R912 B.n659 B.n24 163.367
R913 B.n655 B.n24 163.367
R914 B.n655 B.n26 163.367
R915 B.n651 B.n26 163.367
R916 B.n651 B.n31 163.367
R917 B.n647 B.n31 163.367
R918 B.n647 B.n33 163.367
R919 B.n643 B.n33 163.367
R920 B.n643 B.n38 163.367
R921 B.n639 B.n38 163.367
R922 B.n639 B.n40 163.367
R923 B.n635 B.n40 163.367
R924 B.n635 B.n45 163.367
R925 B.n631 B.n45 163.367
R926 B.n631 B.n47 163.367
R927 B.n627 B.n47 163.367
R928 B.n627 B.n52 163.367
R929 B.n623 B.n52 163.367
R930 B.n623 B.n54 163.367
R931 B.n619 B.n54 163.367
R932 B.n619 B.n59 163.367
R933 B.n615 B.n59 163.367
R934 B.n615 B.n61 163.367
R935 B.n611 B.n61 163.367
R936 B.n611 B.n65 163.367
R937 B.n607 B.n65 163.367
R938 B.n607 B.n67 163.367
R939 B.n603 B.n67 163.367
R940 B.n603 B.n73 163.367
R941 B.n599 B.n73 163.367
R942 B.n599 B.n75 163.367
R943 B.n595 B.n75 163.367
R944 B.n595 B.n80 163.367
R945 B.n591 B.n80 163.367
R946 B.n591 B.n82 163.367
R947 B.n587 B.n82 163.367
R948 B.n587 B.n87 163.367
R949 B.n583 B.n87 163.367
R950 B.n583 B.n89 163.367
R951 B.n579 B.n89 163.367
R952 B.n579 B.n94 163.367
R953 B.n575 B.n94 163.367
R954 B.n575 B.n96 163.367
R955 B.n344 B.n268 126.246
R956 B.n344 B.n264 126.246
R957 B.n350 B.n264 126.246
R958 B.n350 B.n260 126.246
R959 B.n356 B.n260 126.246
R960 B.n356 B.n256 126.246
R961 B.n362 B.n256 126.246
R962 B.n368 B.n252 126.246
R963 B.n368 B.n248 126.246
R964 B.n374 B.n248 126.246
R965 B.n374 B.n244 126.246
R966 B.n380 B.n244 126.246
R967 B.n380 B.n240 126.246
R968 B.n386 B.n240 126.246
R969 B.n386 B.n236 126.246
R970 B.n393 B.n236 126.246
R971 B.n393 B.n392 126.246
R972 B.n399 B.n229 126.246
R973 B.n405 B.n229 126.246
R974 B.n405 B.n225 126.246
R975 B.n411 B.n225 126.246
R976 B.n411 B.n221 126.246
R977 B.n417 B.n221 126.246
R978 B.n423 B.n217 126.246
R979 B.n423 B.n213 126.246
R980 B.n429 B.n213 126.246
R981 B.n429 B.n209 126.246
R982 B.n435 B.n209 126.246
R983 B.n435 B.n205 126.246
R984 B.n441 B.n205 126.246
R985 B.n447 B.n201 126.246
R986 B.n447 B.n197 126.246
R987 B.n453 B.n197 126.246
R988 B.n453 B.n192 126.246
R989 B.n459 B.n192 126.246
R990 B.n459 B.n193 126.246
R991 B.n465 B.n185 126.246
R992 B.n471 B.n185 126.246
R993 B.n471 B.n181 126.246
R994 B.n477 B.n181 126.246
R995 B.n477 B.n176 126.246
R996 B.n483 B.n176 126.246
R997 B.n483 B.n177 126.246
R998 B.n490 B.n169 126.246
R999 B.n496 B.n169 126.246
R1000 B.n496 B.n4 126.246
R1001 B.n679 B.n4 126.246
R1002 B.n679 B.n678 126.246
R1003 B.n678 B.n677 126.246
R1004 B.n677 B.n8 126.246
R1005 B.n12 B.n8 126.246
R1006 B.n670 B.n12 126.246
R1007 B.n669 B.n668 126.246
R1008 B.n668 B.n16 126.246
R1009 B.n662 B.n16 126.246
R1010 B.n662 B.n661 126.246
R1011 B.n661 B.n660 126.246
R1012 B.n660 B.n23 126.246
R1013 B.n654 B.n23 126.246
R1014 B.n653 B.n652 126.246
R1015 B.n652 B.n30 126.246
R1016 B.n646 B.n30 126.246
R1017 B.n646 B.n645 126.246
R1018 B.n645 B.n644 126.246
R1019 B.n644 B.n37 126.246
R1020 B.n638 B.n637 126.246
R1021 B.n637 B.n636 126.246
R1022 B.n636 B.n44 126.246
R1023 B.n630 B.n44 126.246
R1024 B.n630 B.n629 126.246
R1025 B.n629 B.n628 126.246
R1026 B.n628 B.n51 126.246
R1027 B.n622 B.n621 126.246
R1028 B.n621 B.n620 126.246
R1029 B.n620 B.n58 126.246
R1030 B.n614 B.n58 126.246
R1031 B.n614 B.n613 126.246
R1032 B.n613 B.n612 126.246
R1033 B.n606 B.n68 126.246
R1034 B.n606 B.n605 126.246
R1035 B.n605 B.n604 126.246
R1036 B.n604 B.n72 126.246
R1037 B.n598 B.n72 126.246
R1038 B.n598 B.n597 126.246
R1039 B.n597 B.n596 126.246
R1040 B.n596 B.n79 126.246
R1041 B.n590 B.n79 126.246
R1042 B.n590 B.n589 126.246
R1043 B.n588 B.n86 126.246
R1044 B.n582 B.n86 126.246
R1045 B.n582 B.n581 126.246
R1046 B.n581 B.n580 126.246
R1047 B.n580 B.n93 126.246
R1048 B.n574 B.n93 126.246
R1049 B.n574 B.n573 126.246
R1050 B.n399 B.t5 124.388
R1051 B.n612 B.t1 124.388
R1052 B.t8 B.n201 116.963
R1053 B.t3 B.n37 116.963
R1054 B.n490 B.t6 109.537
R1055 B.n670 B.t4 109.537
R1056 B.t15 B.n252 90.971
R1057 B.n589 B.t11 90.971
R1058 B.n193 B.t2 76.1186
R1059 B.t7 B.n653 76.1186
R1060 B.n118 B.n99 71.676
R1061 B.n122 B.n100 71.676
R1062 B.n126 B.n101 71.676
R1063 B.n130 B.n102 71.676
R1064 B.n134 B.n103 71.676
R1065 B.n138 B.n104 71.676
R1066 B.n142 B.n105 71.676
R1067 B.n146 B.n106 71.676
R1068 B.n150 B.n107 71.676
R1069 B.n154 B.n108 71.676
R1070 B.n158 B.n109 71.676
R1071 B.n162 B.n110 71.676
R1072 B.n571 B.n111 71.676
R1073 B.n571 B.n570 71.676
R1074 B.n164 B.n110 71.676
R1075 B.n161 B.n109 71.676
R1076 B.n157 B.n108 71.676
R1077 B.n153 B.n107 71.676
R1078 B.n149 B.n106 71.676
R1079 B.n145 B.n105 71.676
R1080 B.n141 B.n104 71.676
R1081 B.n137 B.n103 71.676
R1082 B.n133 B.n102 71.676
R1083 B.n129 B.n101 71.676
R1084 B.n125 B.n100 71.676
R1085 B.n121 B.n99 71.676
R1086 B.n337 B.n336 71.676
R1087 B.n331 B.n272 71.676
R1088 B.n328 B.n273 71.676
R1089 B.n324 B.n274 71.676
R1090 B.n319 B.n275 71.676
R1091 B.n315 B.n276 71.676
R1092 B.n311 B.n277 71.676
R1093 B.n307 B.n278 71.676
R1094 B.n303 B.n279 71.676
R1095 B.n298 B.n280 71.676
R1096 B.n294 B.n281 71.676
R1097 B.n290 B.n282 71.676
R1098 B.n337 B.n284 71.676
R1099 B.n329 B.n272 71.676
R1100 B.n325 B.n273 71.676
R1101 B.n320 B.n274 71.676
R1102 B.n316 B.n275 71.676
R1103 B.n312 B.n276 71.676
R1104 B.n308 B.n277 71.676
R1105 B.n304 B.n278 71.676
R1106 B.n299 B.n279 71.676
R1107 B.n295 B.n280 71.676
R1108 B.n291 B.n281 71.676
R1109 B.n282 B.n271 71.676
R1110 B.n681 B.n680 71.676
R1111 B.n681 B.n2 71.676
R1112 B.n417 B.t9 68.6925
R1113 B.n622 B.t0 68.6925
R1114 B.n117 B.n116 59.5399
R1115 B.n114 B.n113 59.5399
R1116 B.n301 B.n288 59.5399
R1117 B.n322 B.n286 59.5399
R1118 B.t9 B.n217 57.5532
R1119 B.t0 B.n51 57.5532
R1120 B.n465 B.t2 50.1271
R1121 B.n654 B.t7 50.1271
R1122 B.n116 B.n115 49.649
R1123 B.n113 B.n112 49.649
R1124 B.n288 B.n287 49.649
R1125 B.n286 B.n285 49.649
R1126 B.n362 B.t15 35.2748
R1127 B.t11 B.n588 35.2748
R1128 B.n335 B.n266 30.4395
R1129 B.n341 B.n340 30.4395
R1130 B.n119 B.n95 30.4395
R1131 B.n569 B.n568 30.4395
R1132 B B.n682 18.0485
R1133 B.n177 B.t6 16.7094
R1134 B.t4 B.n669 16.7094
R1135 B.n346 B.n266 10.6151
R1136 B.n347 B.n346 10.6151
R1137 B.n348 B.n347 10.6151
R1138 B.n348 B.n258 10.6151
R1139 B.n358 B.n258 10.6151
R1140 B.n359 B.n358 10.6151
R1141 B.n360 B.n359 10.6151
R1142 B.n360 B.n250 10.6151
R1143 B.n370 B.n250 10.6151
R1144 B.n371 B.n370 10.6151
R1145 B.n372 B.n371 10.6151
R1146 B.n372 B.n242 10.6151
R1147 B.n382 B.n242 10.6151
R1148 B.n383 B.n382 10.6151
R1149 B.n384 B.n383 10.6151
R1150 B.n384 B.n234 10.6151
R1151 B.n395 B.n234 10.6151
R1152 B.n396 B.n395 10.6151
R1153 B.n397 B.n396 10.6151
R1154 B.n397 B.n227 10.6151
R1155 B.n407 B.n227 10.6151
R1156 B.n408 B.n407 10.6151
R1157 B.n409 B.n408 10.6151
R1158 B.n409 B.n219 10.6151
R1159 B.n419 B.n219 10.6151
R1160 B.n420 B.n419 10.6151
R1161 B.n421 B.n420 10.6151
R1162 B.n421 B.n211 10.6151
R1163 B.n431 B.n211 10.6151
R1164 B.n432 B.n431 10.6151
R1165 B.n433 B.n432 10.6151
R1166 B.n433 B.n203 10.6151
R1167 B.n443 B.n203 10.6151
R1168 B.n444 B.n443 10.6151
R1169 B.n445 B.n444 10.6151
R1170 B.n445 B.n195 10.6151
R1171 B.n455 B.n195 10.6151
R1172 B.n456 B.n455 10.6151
R1173 B.n457 B.n456 10.6151
R1174 B.n457 B.n187 10.6151
R1175 B.n467 B.n187 10.6151
R1176 B.n468 B.n467 10.6151
R1177 B.n469 B.n468 10.6151
R1178 B.n469 B.n179 10.6151
R1179 B.n479 B.n179 10.6151
R1180 B.n480 B.n479 10.6151
R1181 B.n481 B.n480 10.6151
R1182 B.n481 B.n171 10.6151
R1183 B.n492 B.n171 10.6151
R1184 B.n493 B.n492 10.6151
R1185 B.n494 B.n493 10.6151
R1186 B.n494 B.n0 10.6151
R1187 B.n335 B.n334 10.6151
R1188 B.n334 B.n333 10.6151
R1189 B.n333 B.n332 10.6151
R1190 B.n332 B.n330 10.6151
R1191 B.n330 B.n327 10.6151
R1192 B.n327 B.n326 10.6151
R1193 B.n326 B.n323 10.6151
R1194 B.n321 B.n318 10.6151
R1195 B.n318 B.n317 10.6151
R1196 B.n317 B.n314 10.6151
R1197 B.n314 B.n313 10.6151
R1198 B.n313 B.n310 10.6151
R1199 B.n310 B.n309 10.6151
R1200 B.n309 B.n306 10.6151
R1201 B.n306 B.n305 10.6151
R1202 B.n305 B.n302 10.6151
R1203 B.n300 B.n297 10.6151
R1204 B.n297 B.n296 10.6151
R1205 B.n296 B.n293 10.6151
R1206 B.n293 B.n292 10.6151
R1207 B.n292 B.n289 10.6151
R1208 B.n289 B.n270 10.6151
R1209 B.n340 B.n270 10.6151
R1210 B.n342 B.n341 10.6151
R1211 B.n342 B.n262 10.6151
R1212 B.n352 B.n262 10.6151
R1213 B.n353 B.n352 10.6151
R1214 B.n354 B.n353 10.6151
R1215 B.n354 B.n254 10.6151
R1216 B.n364 B.n254 10.6151
R1217 B.n365 B.n364 10.6151
R1218 B.n366 B.n365 10.6151
R1219 B.n366 B.n246 10.6151
R1220 B.n376 B.n246 10.6151
R1221 B.n377 B.n376 10.6151
R1222 B.n378 B.n377 10.6151
R1223 B.n378 B.n238 10.6151
R1224 B.n388 B.n238 10.6151
R1225 B.n389 B.n388 10.6151
R1226 B.n390 B.n389 10.6151
R1227 B.n390 B.n231 10.6151
R1228 B.n401 B.n231 10.6151
R1229 B.n402 B.n401 10.6151
R1230 B.n403 B.n402 10.6151
R1231 B.n403 B.n223 10.6151
R1232 B.n413 B.n223 10.6151
R1233 B.n414 B.n413 10.6151
R1234 B.n415 B.n414 10.6151
R1235 B.n415 B.n215 10.6151
R1236 B.n425 B.n215 10.6151
R1237 B.n426 B.n425 10.6151
R1238 B.n427 B.n426 10.6151
R1239 B.n427 B.n207 10.6151
R1240 B.n437 B.n207 10.6151
R1241 B.n438 B.n437 10.6151
R1242 B.n439 B.n438 10.6151
R1243 B.n439 B.n199 10.6151
R1244 B.n449 B.n199 10.6151
R1245 B.n450 B.n449 10.6151
R1246 B.n451 B.n450 10.6151
R1247 B.n451 B.n190 10.6151
R1248 B.n461 B.n190 10.6151
R1249 B.n462 B.n461 10.6151
R1250 B.n463 B.n462 10.6151
R1251 B.n463 B.n183 10.6151
R1252 B.n473 B.n183 10.6151
R1253 B.n474 B.n473 10.6151
R1254 B.n475 B.n474 10.6151
R1255 B.n475 B.n174 10.6151
R1256 B.n485 B.n174 10.6151
R1257 B.n486 B.n485 10.6151
R1258 B.n488 B.n486 10.6151
R1259 B.n488 B.n487 10.6151
R1260 B.n487 B.n167 10.6151
R1261 B.n499 B.n167 10.6151
R1262 B.n500 B.n499 10.6151
R1263 B.n501 B.n500 10.6151
R1264 B.n502 B.n501 10.6151
R1265 B.n503 B.n502 10.6151
R1266 B.n506 B.n503 10.6151
R1267 B.n507 B.n506 10.6151
R1268 B.n508 B.n507 10.6151
R1269 B.n509 B.n508 10.6151
R1270 B.n511 B.n509 10.6151
R1271 B.n512 B.n511 10.6151
R1272 B.n513 B.n512 10.6151
R1273 B.n514 B.n513 10.6151
R1274 B.n516 B.n514 10.6151
R1275 B.n517 B.n516 10.6151
R1276 B.n518 B.n517 10.6151
R1277 B.n519 B.n518 10.6151
R1278 B.n521 B.n519 10.6151
R1279 B.n522 B.n521 10.6151
R1280 B.n523 B.n522 10.6151
R1281 B.n524 B.n523 10.6151
R1282 B.n526 B.n524 10.6151
R1283 B.n527 B.n526 10.6151
R1284 B.n528 B.n527 10.6151
R1285 B.n529 B.n528 10.6151
R1286 B.n531 B.n529 10.6151
R1287 B.n532 B.n531 10.6151
R1288 B.n533 B.n532 10.6151
R1289 B.n534 B.n533 10.6151
R1290 B.n536 B.n534 10.6151
R1291 B.n537 B.n536 10.6151
R1292 B.n538 B.n537 10.6151
R1293 B.n539 B.n538 10.6151
R1294 B.n541 B.n539 10.6151
R1295 B.n542 B.n541 10.6151
R1296 B.n543 B.n542 10.6151
R1297 B.n544 B.n543 10.6151
R1298 B.n546 B.n544 10.6151
R1299 B.n547 B.n546 10.6151
R1300 B.n548 B.n547 10.6151
R1301 B.n549 B.n548 10.6151
R1302 B.n551 B.n549 10.6151
R1303 B.n552 B.n551 10.6151
R1304 B.n553 B.n552 10.6151
R1305 B.n554 B.n553 10.6151
R1306 B.n556 B.n554 10.6151
R1307 B.n557 B.n556 10.6151
R1308 B.n558 B.n557 10.6151
R1309 B.n559 B.n558 10.6151
R1310 B.n561 B.n559 10.6151
R1311 B.n562 B.n561 10.6151
R1312 B.n563 B.n562 10.6151
R1313 B.n564 B.n563 10.6151
R1314 B.n566 B.n564 10.6151
R1315 B.n567 B.n566 10.6151
R1316 B.n568 B.n567 10.6151
R1317 B.n674 B.n1 10.6151
R1318 B.n674 B.n673 10.6151
R1319 B.n673 B.n672 10.6151
R1320 B.n672 B.n10 10.6151
R1321 B.n666 B.n10 10.6151
R1322 B.n666 B.n665 10.6151
R1323 B.n665 B.n664 10.6151
R1324 B.n664 B.n18 10.6151
R1325 B.n658 B.n18 10.6151
R1326 B.n658 B.n657 10.6151
R1327 B.n657 B.n656 10.6151
R1328 B.n656 B.n25 10.6151
R1329 B.n650 B.n25 10.6151
R1330 B.n650 B.n649 10.6151
R1331 B.n649 B.n648 10.6151
R1332 B.n648 B.n32 10.6151
R1333 B.n642 B.n32 10.6151
R1334 B.n642 B.n641 10.6151
R1335 B.n641 B.n640 10.6151
R1336 B.n640 B.n39 10.6151
R1337 B.n634 B.n39 10.6151
R1338 B.n634 B.n633 10.6151
R1339 B.n633 B.n632 10.6151
R1340 B.n632 B.n46 10.6151
R1341 B.n626 B.n46 10.6151
R1342 B.n626 B.n625 10.6151
R1343 B.n625 B.n624 10.6151
R1344 B.n624 B.n53 10.6151
R1345 B.n618 B.n53 10.6151
R1346 B.n618 B.n617 10.6151
R1347 B.n617 B.n616 10.6151
R1348 B.n616 B.n60 10.6151
R1349 B.n610 B.n60 10.6151
R1350 B.n610 B.n609 10.6151
R1351 B.n609 B.n608 10.6151
R1352 B.n608 B.n66 10.6151
R1353 B.n602 B.n66 10.6151
R1354 B.n602 B.n601 10.6151
R1355 B.n601 B.n600 10.6151
R1356 B.n600 B.n74 10.6151
R1357 B.n594 B.n74 10.6151
R1358 B.n594 B.n593 10.6151
R1359 B.n593 B.n592 10.6151
R1360 B.n592 B.n81 10.6151
R1361 B.n586 B.n81 10.6151
R1362 B.n586 B.n585 10.6151
R1363 B.n585 B.n584 10.6151
R1364 B.n584 B.n88 10.6151
R1365 B.n578 B.n88 10.6151
R1366 B.n578 B.n577 10.6151
R1367 B.n577 B.n576 10.6151
R1368 B.n576 B.n95 10.6151
R1369 B.n120 B.n119 10.6151
R1370 B.n123 B.n120 10.6151
R1371 B.n124 B.n123 10.6151
R1372 B.n127 B.n124 10.6151
R1373 B.n128 B.n127 10.6151
R1374 B.n131 B.n128 10.6151
R1375 B.n132 B.n131 10.6151
R1376 B.n136 B.n135 10.6151
R1377 B.n139 B.n136 10.6151
R1378 B.n140 B.n139 10.6151
R1379 B.n143 B.n140 10.6151
R1380 B.n144 B.n143 10.6151
R1381 B.n147 B.n144 10.6151
R1382 B.n148 B.n147 10.6151
R1383 B.n151 B.n148 10.6151
R1384 B.n152 B.n151 10.6151
R1385 B.n156 B.n155 10.6151
R1386 B.n159 B.n156 10.6151
R1387 B.n160 B.n159 10.6151
R1388 B.n163 B.n160 10.6151
R1389 B.n165 B.n163 10.6151
R1390 B.n166 B.n165 10.6151
R1391 B.n569 B.n166 10.6151
R1392 B.n323 B.n322 9.36635
R1393 B.n301 B.n300 9.36635
R1394 B.n132 B.n117 9.36635
R1395 B.n155 B.n114 9.36635
R1396 B.n441 B.t8 9.2832
R1397 B.n638 B.t3 9.2832
R1398 B.n682 B.n0 8.11757
R1399 B.n682 B.n1 8.11757
R1400 B.n392 B.t5 1.85704
R1401 B.n68 B.t1 1.85704
R1402 B.n322 B.n321 1.24928
R1403 B.n302 B.n301 1.24928
R1404 B.n135 B.n117 1.24928
R1405 B.n152 B.n114 1.24928
R1406 VN.n69 VN.n36 161.3
R1407 VN.n68 VN.n67 161.3
R1408 VN.n66 VN.n37 161.3
R1409 VN.n65 VN.n64 161.3
R1410 VN.n63 VN.n38 161.3
R1411 VN.n61 VN.n60 161.3
R1412 VN.n59 VN.n39 161.3
R1413 VN.n58 VN.n57 161.3
R1414 VN.n56 VN.n40 161.3
R1415 VN.n55 VN.n54 161.3
R1416 VN.n53 VN.n52 161.3
R1417 VN.n51 VN.n42 161.3
R1418 VN.n50 VN.n49 161.3
R1419 VN.n48 VN.n43 161.3
R1420 VN.n47 VN.n46 161.3
R1421 VN.n33 VN.n0 161.3
R1422 VN.n32 VN.n31 161.3
R1423 VN.n30 VN.n1 161.3
R1424 VN.n29 VN.n28 161.3
R1425 VN.n27 VN.n2 161.3
R1426 VN.n25 VN.n24 161.3
R1427 VN.n23 VN.n3 161.3
R1428 VN.n22 VN.n21 161.3
R1429 VN.n20 VN.n4 161.3
R1430 VN.n19 VN.n18 161.3
R1431 VN.n17 VN.n16 161.3
R1432 VN.n15 VN.n6 161.3
R1433 VN.n14 VN.n13 161.3
R1434 VN.n12 VN.n7 161.3
R1435 VN.n11 VN.n10 161.3
R1436 VN.n35 VN.n34 92.6509
R1437 VN.n71 VN.n70 92.6509
R1438 VN.n9 VN.n8 56.0043
R1439 VN.n45 VN.n44 56.0043
R1440 VN.n32 VN.n1 49.2348
R1441 VN.n68 VN.n37 49.2348
R1442 VN.n14 VN.n7 43.4072
R1443 VN.n21 VN.n3 43.4072
R1444 VN.n50 VN.n43 43.4072
R1445 VN.n57 VN.n39 43.4072
R1446 VN VN.n71 42.8391
R1447 VN.n8 VN.t0 40.6547
R1448 VN.n44 VN.t7 40.6547
R1449 VN.n15 VN.n14 37.5796
R1450 VN.n21 VN.n20 37.5796
R1451 VN.n51 VN.n50 37.5796
R1452 VN.n57 VN.n56 37.5796
R1453 VN.n28 VN.n1 31.752
R1454 VN.n64 VN.n37 31.752
R1455 VN.n10 VN.n7 24.4675
R1456 VN.n16 VN.n15 24.4675
R1457 VN.n20 VN.n19 24.4675
R1458 VN.n25 VN.n3 24.4675
R1459 VN.n28 VN.n27 24.4675
R1460 VN.n33 VN.n32 24.4675
R1461 VN.n46 VN.n43 24.4675
R1462 VN.n56 VN.n55 24.4675
R1463 VN.n52 VN.n51 24.4675
R1464 VN.n64 VN.n63 24.4675
R1465 VN.n61 VN.n39 24.4675
R1466 VN.n69 VN.n68 24.4675
R1467 VN.n34 VN.n33 18.1061
R1468 VN.n70 VN.n69 18.1061
R1469 VN.n10 VN.n9 15.17
R1470 VN.n26 VN.n25 15.17
R1471 VN.n46 VN.n45 15.17
R1472 VN.n62 VN.n61 15.17
R1473 VN.n16 VN.n5 12.234
R1474 VN.n19 VN.n5 12.234
R1475 VN.n55 VN.n41 12.234
R1476 VN.n52 VN.n41 12.234
R1477 VN.n27 VN.n26 9.29796
R1478 VN.n63 VN.n62 9.29796
R1479 VN.n47 VN.n44 9.14908
R1480 VN.n11 VN.n8 9.14908
R1481 VN.n9 VN.t2 7.02516
R1482 VN.n5 VN.t1 7.02516
R1483 VN.n26 VN.t5 7.02516
R1484 VN.n34 VN.t4 7.02516
R1485 VN.n45 VN.t3 7.02516
R1486 VN.n41 VN.t9 7.02516
R1487 VN.n62 VN.t6 7.02516
R1488 VN.n70 VN.t8 7.02516
R1489 VN.n71 VN.n36 0.278367
R1490 VN.n35 VN.n0 0.278367
R1491 VN.n67 VN.n36 0.189894
R1492 VN.n67 VN.n66 0.189894
R1493 VN.n66 VN.n65 0.189894
R1494 VN.n65 VN.n38 0.189894
R1495 VN.n60 VN.n38 0.189894
R1496 VN.n60 VN.n59 0.189894
R1497 VN.n59 VN.n58 0.189894
R1498 VN.n58 VN.n40 0.189894
R1499 VN.n54 VN.n40 0.189894
R1500 VN.n54 VN.n53 0.189894
R1501 VN.n53 VN.n42 0.189894
R1502 VN.n49 VN.n42 0.189894
R1503 VN.n49 VN.n48 0.189894
R1504 VN.n48 VN.n47 0.189894
R1505 VN.n12 VN.n11 0.189894
R1506 VN.n13 VN.n12 0.189894
R1507 VN.n13 VN.n6 0.189894
R1508 VN.n17 VN.n6 0.189894
R1509 VN.n18 VN.n17 0.189894
R1510 VN.n18 VN.n4 0.189894
R1511 VN.n22 VN.n4 0.189894
R1512 VN.n23 VN.n22 0.189894
R1513 VN.n24 VN.n23 0.189894
R1514 VN.n24 VN.n2 0.189894
R1515 VN.n29 VN.n2 0.189894
R1516 VN.n30 VN.n29 0.189894
R1517 VN.n31 VN.n30 0.189894
R1518 VN.n31 VN.n0 0.189894
R1519 VN VN.n35 0.153454
R1520 VDD2.n1 VDD2.t9 267.502
R1521 VDD2.n4 VDD2.t1 265.296
R1522 VDD2.n3 VDD2.n2 236.434
R1523 VDD2 VDD2.n7 236.43
R1524 VDD2.n6 VDD2.n5 234.833
R1525 VDD2.n1 VDD2.n0 234.833
R1526 VDD2.n4 VDD2.n3 34.7584
R1527 VDD2.n7 VDD2.t6 30.462
R1528 VDD2.n7 VDD2.t2 30.462
R1529 VDD2.n5 VDD2.t3 30.462
R1530 VDD2.n5 VDD2.t0 30.462
R1531 VDD2.n2 VDD2.t4 30.462
R1532 VDD2.n2 VDD2.t5 30.462
R1533 VDD2.n0 VDD2.t7 30.462
R1534 VDD2.n0 VDD2.t8 30.462
R1535 VDD2.n6 VDD2.n4 2.2074
R1536 VDD2 VDD2.n6 0.610414
R1537 VDD2.n3 VDD2.n1 0.496878
C0 VTAIL VN 2.49459f
C1 VDD1 VP 1.43202f
C2 VTAIL VDD2 4.76504f
C3 VDD2 VN 1.0514f
C4 VTAIL VDD1 4.71397f
C5 VTAIL VP 2.50871f
C6 VDD1 VN 0.160796f
C7 VN VP 5.76038f
C8 VDD1 VDD2 1.93054f
C9 VDD2 VP 0.546006f
C10 VDD2 B 4.571026f
C11 VDD1 B 4.68656f
C12 VTAIL B 2.958557f
C13 VN B 15.435739f
C14 VP B 13.841603f
C15 VDD2.t9 B 0.054835f
C16 VDD2.t7 B 0.011157f
C17 VDD2.t8 B 0.011157f
C18 VDD2.n0 B 0.02799f
C19 VDD2.n1 B 0.466993f
C20 VDD2.t4 B 0.011157f
C21 VDD2.t5 B 0.011157f
C22 VDD2.n2 B 0.030226f
C23 VDD2.n3 B 1.65466f
C24 VDD2.t1 B 0.05299f
C25 VDD2.n4 B 1.63051f
C26 VDD2.t3 B 0.011157f
C27 VDD2.t0 B 0.011157f
C28 VDD2.n5 B 0.02799f
C29 VDD2.n6 B 0.25214f
C30 VDD2.t6 B 0.011157f
C31 VDD2.t2 B 0.011157f
C32 VDD2.n7 B 0.030219f
C33 VN.n0 B 0.043364f
C34 VN.t4 B 0.065093f
C35 VN.n1 B 0.030179f
C36 VN.n2 B 0.032892f
C37 VN.t5 B 0.065093f
C38 VN.n3 B 0.064205f
C39 VN.n4 B 0.032892f
C40 VN.t1 B 0.065093f
C41 VN.n5 B 0.074802f
C42 VN.n6 B 0.032892f
C43 VN.n7 B 0.064205f
C44 VN.t0 B 0.278502f
C45 VN.n8 B 0.146183f
C46 VN.t2 B 0.065093f
C47 VN.n9 B 0.163704f
C48 VN.n10 B 0.049801f
C49 VN.n11 B 0.280936f
C50 VN.n12 B 0.032892f
C51 VN.n13 B 0.032892f
C52 VN.n14 B 0.026972f
C53 VN.n15 B 0.066157f
C54 VN.n16 B 0.046169f
C55 VN.n17 B 0.032892f
C56 VN.n18 B 0.032892f
C57 VN.n19 B 0.046169f
C58 VN.n20 B 0.066157f
C59 VN.n21 B 0.026972f
C60 VN.n22 B 0.032892f
C61 VN.n23 B 0.032892f
C62 VN.n24 B 0.032892f
C63 VN.n25 B 0.049801f
C64 VN.n26 B 0.074802f
C65 VN.n27 B 0.042537f
C66 VN.n28 B 0.06616f
C67 VN.n29 B 0.032892f
C68 VN.n30 B 0.032892f
C69 VN.n31 B 0.032892f
C70 VN.n32 B 0.060995f
C71 VN.n33 B 0.053433f
C72 VN.n34 B 0.183616f
C73 VN.n35 B 0.042915f
C74 VN.n36 B 0.043364f
C75 VN.t8 B 0.065093f
C76 VN.n37 B 0.030179f
C77 VN.n38 B 0.032892f
C78 VN.t6 B 0.065093f
C79 VN.n39 B 0.064205f
C80 VN.n40 B 0.032892f
C81 VN.t9 B 0.065093f
C82 VN.n41 B 0.074802f
C83 VN.n42 B 0.032892f
C84 VN.n43 B 0.064205f
C85 VN.t7 B 0.278502f
C86 VN.n44 B 0.146183f
C87 VN.t3 B 0.065093f
C88 VN.n45 B 0.163704f
C89 VN.n46 B 0.049801f
C90 VN.n47 B 0.280936f
C91 VN.n48 B 0.032892f
C92 VN.n49 B 0.032892f
C93 VN.n50 B 0.026972f
C94 VN.n51 B 0.066157f
C95 VN.n52 B 0.046169f
C96 VN.n53 B 0.032892f
C97 VN.n54 B 0.032892f
C98 VN.n55 B 0.046169f
C99 VN.n56 B 0.066157f
C100 VN.n57 B 0.026972f
C101 VN.n58 B 0.032892f
C102 VN.n59 B 0.032892f
C103 VN.n60 B 0.032892f
C104 VN.n61 B 0.049801f
C105 VN.n62 B 0.074802f
C106 VN.n63 B 0.042537f
C107 VN.n64 B 0.06616f
C108 VN.n65 B 0.032892f
C109 VN.n66 B 0.032892f
C110 VN.n67 B 0.032892f
C111 VN.n68 B 0.060995f
C112 VN.n69 B 0.053433f
C113 VN.n70 B 0.183616f
C114 VN.n71 B 1.43737f
C115 VTAIL.t4 B 0.026445f
C116 VTAIL.t19 B 0.026445f
C117 VTAIL.n0 B 0.057128f
C118 VTAIL.n1 B 0.614837f
C119 VTAIL.t10 B 0.116654f
C120 VTAIL.n2 B 0.709307f
C121 VTAIL.t12 B 0.026445f
C122 VTAIL.t9 B 0.026445f
C123 VTAIL.n3 B 0.057128f
C124 VTAIL.n4 B 0.801824f
C125 VTAIL.t15 B 0.026445f
C126 VTAIL.t13 B 0.026445f
C127 VTAIL.n5 B 0.057128f
C128 VTAIL.n6 B 1.96023f
C129 VTAIL.t5 B 0.026445f
C130 VTAIL.t18 B 0.026445f
C131 VTAIL.n7 B 0.057128f
C132 VTAIL.n8 B 1.96023f
C133 VTAIL.t17 B 0.026445f
C134 VTAIL.t2 B 0.026445f
C135 VTAIL.n9 B 0.057128f
C136 VTAIL.n10 B 0.801824f
C137 VTAIL.t6 B 0.116654f
C138 VTAIL.n11 B 0.709307f
C139 VTAIL.t14 B 0.026445f
C140 VTAIL.t7 B 0.026445f
C141 VTAIL.n12 B 0.057128f
C142 VTAIL.n13 B 0.696711f
C143 VTAIL.t8 B 0.026445f
C144 VTAIL.t16 B 0.026445f
C145 VTAIL.n14 B 0.057128f
C146 VTAIL.n15 B 0.801824f
C147 VTAIL.t11 B 0.116654f
C148 VTAIL.n16 B 1.60672f
C149 VTAIL.t1 B 0.116654f
C150 VTAIL.n17 B 1.60672f
C151 VTAIL.t3 B 0.026445f
C152 VTAIL.t0 B 0.026445f
C153 VTAIL.n18 B 0.057128f
C154 VTAIL.n19 B 0.51759f
C155 VDD1.t8 B 0.05281f
C156 VDD1.t5 B 0.010744f
C157 VDD1.t9 B 0.010744f
C158 VDD1.n0 B 0.026956f
C159 VDD1.n1 B 0.456422f
C160 VDD1.t2 B 0.05281f
C161 VDD1.t1 B 0.010744f
C162 VDD1.t3 B 0.010744f
C163 VDD1.n2 B 0.026956f
C164 VDD1.n3 B 0.449747f
C165 VDD1.t0 B 0.010744f
C166 VDD1.t6 B 0.010744f
C167 VDD1.n4 B 0.02911f
C168 VDD1.n5 B 1.68132f
C169 VDD1.t7 B 0.010744f
C170 VDD1.t4 B 0.010744f
C171 VDD1.n6 B 0.026956f
C172 VDD1.n7 B 1.66221f
C173 VP.n0 B 0.043607f
C174 VP.t6 B 0.065458f
C175 VP.n1 B 0.030348f
C176 VP.n2 B 0.033076f
C177 VP.t7 B 0.065458f
C178 VP.n3 B 0.064564f
C179 VP.n4 B 0.033076f
C180 VP.t4 B 0.065458f
C181 VP.n5 B 0.075221f
C182 VP.n6 B 0.033076f
C183 VP.n7 B 0.064564f
C184 VP.n8 B 0.033076f
C185 VP.t3 B 0.065458f
C186 VP.n9 B 0.030348f
C187 VP.n10 B 0.043607f
C188 VP.t1 B 0.065458f
C189 VP.n11 B 0.043607f
C190 VP.t5 B 0.065458f
C191 VP.n12 B 0.030348f
C192 VP.n13 B 0.033076f
C193 VP.t0 B 0.065458f
C194 VP.n14 B 0.064564f
C195 VP.n15 B 0.033076f
C196 VP.t8 B 0.065458f
C197 VP.n16 B 0.075221f
C198 VP.n17 B 0.033076f
C199 VP.n18 B 0.064564f
C200 VP.t2 B 0.280062f
C201 VP.n19 B 0.147002f
C202 VP.t9 B 0.065458f
C203 VP.n20 B 0.164621f
C204 VP.n21 B 0.05008f
C205 VP.n22 B 0.28251f
C206 VP.n23 B 0.033076f
C207 VP.n24 B 0.033076f
C208 VP.n25 B 0.027123f
C209 VP.n26 B 0.066528f
C210 VP.n27 B 0.046428f
C211 VP.n28 B 0.033076f
C212 VP.n29 B 0.033076f
C213 VP.n30 B 0.046428f
C214 VP.n31 B 0.066528f
C215 VP.n32 B 0.027123f
C216 VP.n33 B 0.033076f
C217 VP.n34 B 0.033076f
C218 VP.n35 B 0.033076f
C219 VP.n36 B 0.05008f
C220 VP.n37 B 0.075221f
C221 VP.n38 B 0.042776f
C222 VP.n39 B 0.066531f
C223 VP.n40 B 0.033076f
C224 VP.n41 B 0.033076f
C225 VP.n42 B 0.033076f
C226 VP.n43 B 0.061336f
C227 VP.n44 B 0.053732f
C228 VP.n45 B 0.184645f
C229 VP.n46 B 1.42715f
C230 VP.n47 B 1.45509f
C231 VP.n48 B 0.184645f
C232 VP.n49 B 0.053732f
C233 VP.n50 B 0.061336f
C234 VP.n51 B 0.033076f
C235 VP.n52 B 0.033076f
C236 VP.n53 B 0.033076f
C237 VP.n54 B 0.066531f
C238 VP.n55 B 0.042776f
C239 VP.n56 B 0.075221f
C240 VP.n57 B 0.05008f
C241 VP.n58 B 0.033076f
C242 VP.n59 B 0.033076f
C243 VP.n60 B 0.033076f
C244 VP.n61 B 0.027123f
C245 VP.n62 B 0.066528f
C246 VP.n63 B 0.046428f
C247 VP.n64 B 0.033076f
C248 VP.n65 B 0.033076f
C249 VP.n66 B 0.046428f
C250 VP.n67 B 0.066528f
C251 VP.n68 B 0.027123f
C252 VP.n69 B 0.033076f
C253 VP.n70 B 0.033076f
C254 VP.n71 B 0.033076f
C255 VP.n72 B 0.05008f
C256 VP.n73 B 0.075221f
C257 VP.n74 B 0.042776f
C258 VP.n75 B 0.066531f
C259 VP.n76 B 0.033076f
C260 VP.n77 B 0.033076f
C261 VP.n78 B 0.033076f
C262 VP.n79 B 0.061336f
C263 VP.n80 B 0.053732f
C264 VP.n81 B 0.184645f
C265 VP.n82 B 0.043155f
.ends

