* NGSPICE file created from diff_pair_sample_0015.ext - technology: sky130A

.subckt diff_pair_sample_0015 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=2.71095 ps=16.76 w=16.43 l=1.51
X1 VDD1.t2 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.71095 pd=16.76 as=6.4077 ps=33.64 w=16.43 l=1.51
X2 VDD1.t3 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.71095 pd=16.76 as=6.4077 ps=33.64 w=16.43 l=1.51
X3 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=0 ps=0 w=16.43 l=1.51
X4 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=0 ps=0 w=16.43 l=1.51
X5 VDD2.t3 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.71095 pd=16.76 as=6.4077 ps=33.64 w=16.43 l=1.51
X6 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=2.71095 ps=16.76 w=16.43 l=1.51
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=0 ps=0 w=16.43 l=1.51
X8 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.71095 pd=16.76 as=6.4077 ps=33.64 w=16.43 l=1.51
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=0 ps=0 w=16.43 l=1.51
X10 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=2.71095 ps=16.76 w=16.43 l=1.51
X11 VTAIL.t4 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4077 pd=33.64 as=2.71095 ps=16.76 w=16.43 l=1.51
R0 VP.n2 VP.t3 298.733
R1 VP.n2 VP.t2 298.416
R2 VP.n4 VP.t0 262.228
R3 VP.n11 VP.t1 262.228
R4 VP.n4 VP.n3 177.448
R5 VP.n12 VP.n11 177.448
R6 VP.n10 VP.n0 161.3
R7 VP.n9 VP.n8 161.3
R8 VP.n7 VP.n1 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n3 VP.n2 59.2431
R11 VP.n9 VP.n1 56.5193
R12 VP.n5 VP.n1 24.4675
R13 VP.n10 VP.n9 24.4675
R14 VP.n5 VP.n4 8.31928
R15 VP.n11 VP.n10 8.31928
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VDD1 VDD1.n1 103.718
R23 VDD1 VDD1.n0 60.6137
R24 VDD1.n0 VDD1.t0 1.20561
R25 VDD1.n0 VDD1.t3 1.20561
R26 VDD1.n1 VDD1.t1 1.20561
R27 VDD1.n1 VDD1.t2 1.20561
R28 VTAIL.n5 VTAIL.t4 45.082
R29 VTAIL.n4 VTAIL.t3 45.082
R30 VTAIL.n3 VTAIL.t0 45.082
R31 VTAIL.n7 VTAIL.t1 45.0818
R32 VTAIL.n0 VTAIL.t2 45.0818
R33 VTAIL.n1 VTAIL.t6 45.0818
R34 VTAIL.n2 VTAIL.t7 45.0818
R35 VTAIL.n6 VTAIL.t5 45.0818
R36 VTAIL.n7 VTAIL.n6 28.1169
R37 VTAIL.n3 VTAIL.n2 28.1169
R38 VTAIL.n4 VTAIL.n3 1.58671
R39 VTAIL.n6 VTAIL.n5 1.58671
R40 VTAIL.n2 VTAIL.n1 1.58671
R41 VTAIL VTAIL.n0 0.851793
R42 VTAIL VTAIL.n7 0.735414
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 B.n803 B.n802 585
R46 B.n804 B.n803 585
R47 B.n346 B.n107 585
R48 B.n345 B.n344 585
R49 B.n343 B.n342 585
R50 B.n341 B.n340 585
R51 B.n339 B.n338 585
R52 B.n337 B.n336 585
R53 B.n335 B.n334 585
R54 B.n333 B.n332 585
R55 B.n331 B.n330 585
R56 B.n329 B.n328 585
R57 B.n327 B.n326 585
R58 B.n325 B.n324 585
R59 B.n323 B.n322 585
R60 B.n321 B.n320 585
R61 B.n319 B.n318 585
R62 B.n317 B.n316 585
R63 B.n315 B.n314 585
R64 B.n313 B.n312 585
R65 B.n311 B.n310 585
R66 B.n309 B.n308 585
R67 B.n307 B.n306 585
R68 B.n305 B.n304 585
R69 B.n303 B.n302 585
R70 B.n301 B.n300 585
R71 B.n299 B.n298 585
R72 B.n297 B.n296 585
R73 B.n295 B.n294 585
R74 B.n293 B.n292 585
R75 B.n291 B.n290 585
R76 B.n289 B.n288 585
R77 B.n287 B.n286 585
R78 B.n285 B.n284 585
R79 B.n283 B.n282 585
R80 B.n281 B.n280 585
R81 B.n279 B.n278 585
R82 B.n277 B.n276 585
R83 B.n275 B.n274 585
R84 B.n273 B.n272 585
R85 B.n271 B.n270 585
R86 B.n269 B.n268 585
R87 B.n267 B.n266 585
R88 B.n265 B.n264 585
R89 B.n263 B.n262 585
R90 B.n261 B.n260 585
R91 B.n259 B.n258 585
R92 B.n257 B.n256 585
R93 B.n255 B.n254 585
R94 B.n253 B.n252 585
R95 B.n251 B.n250 585
R96 B.n249 B.n248 585
R97 B.n247 B.n246 585
R98 B.n245 B.n244 585
R99 B.n243 B.n242 585
R100 B.n241 B.n240 585
R101 B.n239 B.n238 585
R102 B.n237 B.n236 585
R103 B.n235 B.n234 585
R104 B.n233 B.n232 585
R105 B.n231 B.n230 585
R106 B.n229 B.n228 585
R107 B.n227 B.n226 585
R108 B.n225 B.n224 585
R109 B.n223 B.n222 585
R110 B.n220 B.n219 585
R111 B.n218 B.n217 585
R112 B.n216 B.n215 585
R113 B.n214 B.n213 585
R114 B.n212 B.n211 585
R115 B.n210 B.n209 585
R116 B.n208 B.n207 585
R117 B.n206 B.n205 585
R118 B.n204 B.n203 585
R119 B.n202 B.n201 585
R120 B.n200 B.n199 585
R121 B.n198 B.n197 585
R122 B.n196 B.n195 585
R123 B.n194 B.n193 585
R124 B.n192 B.n191 585
R125 B.n190 B.n189 585
R126 B.n188 B.n187 585
R127 B.n186 B.n185 585
R128 B.n184 B.n183 585
R129 B.n182 B.n181 585
R130 B.n180 B.n179 585
R131 B.n178 B.n177 585
R132 B.n176 B.n175 585
R133 B.n174 B.n173 585
R134 B.n172 B.n171 585
R135 B.n170 B.n169 585
R136 B.n168 B.n167 585
R137 B.n166 B.n165 585
R138 B.n164 B.n163 585
R139 B.n162 B.n161 585
R140 B.n160 B.n159 585
R141 B.n158 B.n157 585
R142 B.n156 B.n155 585
R143 B.n154 B.n153 585
R144 B.n152 B.n151 585
R145 B.n150 B.n149 585
R146 B.n148 B.n147 585
R147 B.n146 B.n145 585
R148 B.n144 B.n143 585
R149 B.n142 B.n141 585
R150 B.n140 B.n139 585
R151 B.n138 B.n137 585
R152 B.n136 B.n135 585
R153 B.n134 B.n133 585
R154 B.n132 B.n131 585
R155 B.n130 B.n129 585
R156 B.n128 B.n127 585
R157 B.n126 B.n125 585
R158 B.n124 B.n123 585
R159 B.n122 B.n121 585
R160 B.n120 B.n119 585
R161 B.n118 B.n117 585
R162 B.n116 B.n115 585
R163 B.n114 B.n113 585
R164 B.n46 B.n45 585
R165 B.n801 B.n47 585
R166 B.n805 B.n47 585
R167 B.n800 B.n799 585
R168 B.n799 B.n43 585
R169 B.n798 B.n42 585
R170 B.n811 B.n42 585
R171 B.n797 B.n41 585
R172 B.n812 B.n41 585
R173 B.n796 B.n40 585
R174 B.n813 B.n40 585
R175 B.n795 B.n794 585
R176 B.n794 B.n36 585
R177 B.n793 B.n35 585
R178 B.n819 B.n35 585
R179 B.n792 B.n34 585
R180 B.n820 B.n34 585
R181 B.n791 B.n33 585
R182 B.n821 B.n33 585
R183 B.n790 B.n789 585
R184 B.n789 B.n29 585
R185 B.n788 B.n28 585
R186 B.n827 B.n28 585
R187 B.n787 B.n27 585
R188 B.n828 B.n27 585
R189 B.n786 B.n26 585
R190 B.n829 B.n26 585
R191 B.n785 B.n784 585
R192 B.n784 B.n22 585
R193 B.n783 B.n21 585
R194 B.n835 B.n21 585
R195 B.n782 B.n20 585
R196 B.n836 B.n20 585
R197 B.n781 B.n19 585
R198 B.n837 B.n19 585
R199 B.n780 B.n779 585
R200 B.n779 B.n15 585
R201 B.n778 B.n14 585
R202 B.n843 B.n14 585
R203 B.n777 B.n13 585
R204 B.n844 B.n13 585
R205 B.n776 B.n12 585
R206 B.n845 B.n12 585
R207 B.n775 B.n774 585
R208 B.n774 B.n773 585
R209 B.n772 B.n771 585
R210 B.n772 B.n8 585
R211 B.n770 B.n7 585
R212 B.n852 B.n7 585
R213 B.n769 B.n6 585
R214 B.n853 B.n6 585
R215 B.n768 B.n5 585
R216 B.n854 B.n5 585
R217 B.n767 B.n766 585
R218 B.n766 B.n4 585
R219 B.n765 B.n347 585
R220 B.n765 B.n764 585
R221 B.n755 B.n348 585
R222 B.n349 B.n348 585
R223 B.n757 B.n756 585
R224 B.n758 B.n757 585
R225 B.n754 B.n354 585
R226 B.n354 B.n353 585
R227 B.n753 B.n752 585
R228 B.n752 B.n751 585
R229 B.n356 B.n355 585
R230 B.n357 B.n356 585
R231 B.n744 B.n743 585
R232 B.n745 B.n744 585
R233 B.n742 B.n362 585
R234 B.n362 B.n361 585
R235 B.n741 B.n740 585
R236 B.n740 B.n739 585
R237 B.n364 B.n363 585
R238 B.n365 B.n364 585
R239 B.n732 B.n731 585
R240 B.n733 B.n732 585
R241 B.n730 B.n370 585
R242 B.n370 B.n369 585
R243 B.n729 B.n728 585
R244 B.n728 B.n727 585
R245 B.n372 B.n371 585
R246 B.n373 B.n372 585
R247 B.n720 B.n719 585
R248 B.n721 B.n720 585
R249 B.n718 B.n378 585
R250 B.n378 B.n377 585
R251 B.n717 B.n716 585
R252 B.n716 B.n715 585
R253 B.n380 B.n379 585
R254 B.n381 B.n380 585
R255 B.n708 B.n707 585
R256 B.n709 B.n708 585
R257 B.n706 B.n386 585
R258 B.n386 B.n385 585
R259 B.n705 B.n704 585
R260 B.n704 B.n703 585
R261 B.n388 B.n387 585
R262 B.n389 B.n388 585
R263 B.n696 B.n695 585
R264 B.n697 B.n696 585
R265 B.n392 B.n391 585
R266 B.n457 B.n456 585
R267 B.n458 B.n454 585
R268 B.n454 B.n393 585
R269 B.n460 B.n459 585
R270 B.n462 B.n453 585
R271 B.n465 B.n464 585
R272 B.n466 B.n452 585
R273 B.n468 B.n467 585
R274 B.n470 B.n451 585
R275 B.n473 B.n472 585
R276 B.n474 B.n450 585
R277 B.n476 B.n475 585
R278 B.n478 B.n449 585
R279 B.n481 B.n480 585
R280 B.n482 B.n448 585
R281 B.n484 B.n483 585
R282 B.n486 B.n447 585
R283 B.n489 B.n488 585
R284 B.n490 B.n446 585
R285 B.n492 B.n491 585
R286 B.n494 B.n445 585
R287 B.n497 B.n496 585
R288 B.n498 B.n444 585
R289 B.n500 B.n499 585
R290 B.n502 B.n443 585
R291 B.n505 B.n504 585
R292 B.n506 B.n442 585
R293 B.n508 B.n507 585
R294 B.n510 B.n441 585
R295 B.n513 B.n512 585
R296 B.n514 B.n440 585
R297 B.n516 B.n515 585
R298 B.n518 B.n439 585
R299 B.n521 B.n520 585
R300 B.n522 B.n438 585
R301 B.n524 B.n523 585
R302 B.n526 B.n437 585
R303 B.n529 B.n528 585
R304 B.n530 B.n436 585
R305 B.n532 B.n531 585
R306 B.n534 B.n435 585
R307 B.n537 B.n536 585
R308 B.n538 B.n434 585
R309 B.n540 B.n539 585
R310 B.n542 B.n433 585
R311 B.n545 B.n544 585
R312 B.n546 B.n432 585
R313 B.n548 B.n547 585
R314 B.n550 B.n431 585
R315 B.n553 B.n552 585
R316 B.n554 B.n430 585
R317 B.n556 B.n555 585
R318 B.n558 B.n429 585
R319 B.n561 B.n560 585
R320 B.n562 B.n426 585
R321 B.n565 B.n564 585
R322 B.n567 B.n425 585
R323 B.n570 B.n569 585
R324 B.n571 B.n424 585
R325 B.n573 B.n572 585
R326 B.n575 B.n423 585
R327 B.n578 B.n577 585
R328 B.n579 B.n422 585
R329 B.n584 B.n583 585
R330 B.n586 B.n421 585
R331 B.n589 B.n588 585
R332 B.n590 B.n420 585
R333 B.n592 B.n591 585
R334 B.n594 B.n419 585
R335 B.n597 B.n596 585
R336 B.n598 B.n418 585
R337 B.n600 B.n599 585
R338 B.n602 B.n417 585
R339 B.n605 B.n604 585
R340 B.n606 B.n416 585
R341 B.n608 B.n607 585
R342 B.n610 B.n415 585
R343 B.n613 B.n612 585
R344 B.n614 B.n414 585
R345 B.n616 B.n615 585
R346 B.n618 B.n413 585
R347 B.n621 B.n620 585
R348 B.n622 B.n412 585
R349 B.n624 B.n623 585
R350 B.n626 B.n411 585
R351 B.n629 B.n628 585
R352 B.n630 B.n410 585
R353 B.n632 B.n631 585
R354 B.n634 B.n409 585
R355 B.n637 B.n636 585
R356 B.n638 B.n408 585
R357 B.n640 B.n639 585
R358 B.n642 B.n407 585
R359 B.n645 B.n644 585
R360 B.n646 B.n406 585
R361 B.n648 B.n647 585
R362 B.n650 B.n405 585
R363 B.n653 B.n652 585
R364 B.n654 B.n404 585
R365 B.n656 B.n655 585
R366 B.n658 B.n403 585
R367 B.n661 B.n660 585
R368 B.n662 B.n402 585
R369 B.n664 B.n663 585
R370 B.n666 B.n401 585
R371 B.n669 B.n668 585
R372 B.n670 B.n400 585
R373 B.n672 B.n671 585
R374 B.n674 B.n399 585
R375 B.n677 B.n676 585
R376 B.n678 B.n398 585
R377 B.n680 B.n679 585
R378 B.n682 B.n397 585
R379 B.n685 B.n684 585
R380 B.n686 B.n396 585
R381 B.n688 B.n687 585
R382 B.n690 B.n395 585
R383 B.n693 B.n692 585
R384 B.n694 B.n394 585
R385 B.n699 B.n698 585
R386 B.n698 B.n697 585
R387 B.n700 B.n390 585
R388 B.n390 B.n389 585
R389 B.n702 B.n701 585
R390 B.n703 B.n702 585
R391 B.n384 B.n383 585
R392 B.n385 B.n384 585
R393 B.n711 B.n710 585
R394 B.n710 B.n709 585
R395 B.n712 B.n382 585
R396 B.n382 B.n381 585
R397 B.n714 B.n713 585
R398 B.n715 B.n714 585
R399 B.n376 B.n375 585
R400 B.n377 B.n376 585
R401 B.n723 B.n722 585
R402 B.n722 B.n721 585
R403 B.n724 B.n374 585
R404 B.n374 B.n373 585
R405 B.n726 B.n725 585
R406 B.n727 B.n726 585
R407 B.n368 B.n367 585
R408 B.n369 B.n368 585
R409 B.n735 B.n734 585
R410 B.n734 B.n733 585
R411 B.n736 B.n366 585
R412 B.n366 B.n365 585
R413 B.n738 B.n737 585
R414 B.n739 B.n738 585
R415 B.n360 B.n359 585
R416 B.n361 B.n360 585
R417 B.n747 B.n746 585
R418 B.n746 B.n745 585
R419 B.n748 B.n358 585
R420 B.n358 B.n357 585
R421 B.n750 B.n749 585
R422 B.n751 B.n750 585
R423 B.n352 B.n351 585
R424 B.n353 B.n352 585
R425 B.n760 B.n759 585
R426 B.n759 B.n758 585
R427 B.n761 B.n350 585
R428 B.n350 B.n349 585
R429 B.n763 B.n762 585
R430 B.n764 B.n763 585
R431 B.n3 B.n0 585
R432 B.n4 B.n3 585
R433 B.n851 B.n1 585
R434 B.n852 B.n851 585
R435 B.n850 B.n849 585
R436 B.n850 B.n8 585
R437 B.n848 B.n9 585
R438 B.n773 B.n9 585
R439 B.n847 B.n846 585
R440 B.n846 B.n845 585
R441 B.n11 B.n10 585
R442 B.n844 B.n11 585
R443 B.n842 B.n841 585
R444 B.n843 B.n842 585
R445 B.n840 B.n16 585
R446 B.n16 B.n15 585
R447 B.n839 B.n838 585
R448 B.n838 B.n837 585
R449 B.n18 B.n17 585
R450 B.n836 B.n18 585
R451 B.n834 B.n833 585
R452 B.n835 B.n834 585
R453 B.n832 B.n23 585
R454 B.n23 B.n22 585
R455 B.n831 B.n830 585
R456 B.n830 B.n829 585
R457 B.n25 B.n24 585
R458 B.n828 B.n25 585
R459 B.n826 B.n825 585
R460 B.n827 B.n826 585
R461 B.n824 B.n30 585
R462 B.n30 B.n29 585
R463 B.n823 B.n822 585
R464 B.n822 B.n821 585
R465 B.n32 B.n31 585
R466 B.n820 B.n32 585
R467 B.n818 B.n817 585
R468 B.n819 B.n818 585
R469 B.n816 B.n37 585
R470 B.n37 B.n36 585
R471 B.n815 B.n814 585
R472 B.n814 B.n813 585
R473 B.n39 B.n38 585
R474 B.n812 B.n39 585
R475 B.n810 B.n809 585
R476 B.n811 B.n810 585
R477 B.n808 B.n44 585
R478 B.n44 B.n43 585
R479 B.n807 B.n806 585
R480 B.n806 B.n805 585
R481 B.n855 B.n854 585
R482 B.n853 B.n2 585
R483 B.n111 B.t8 467.704
R484 B.n108 B.t15 467.704
R485 B.n580 B.t4 467.704
R486 B.n427 B.t12 467.704
R487 B.n806 B.n46 463.671
R488 B.n803 B.n47 463.671
R489 B.n696 B.n394 463.671
R490 B.n698 B.n392 463.671
R491 B.n804 B.n106 256.663
R492 B.n804 B.n105 256.663
R493 B.n804 B.n104 256.663
R494 B.n804 B.n103 256.663
R495 B.n804 B.n102 256.663
R496 B.n804 B.n101 256.663
R497 B.n804 B.n100 256.663
R498 B.n804 B.n99 256.663
R499 B.n804 B.n98 256.663
R500 B.n804 B.n97 256.663
R501 B.n804 B.n96 256.663
R502 B.n804 B.n95 256.663
R503 B.n804 B.n94 256.663
R504 B.n804 B.n93 256.663
R505 B.n804 B.n92 256.663
R506 B.n804 B.n91 256.663
R507 B.n804 B.n90 256.663
R508 B.n804 B.n89 256.663
R509 B.n804 B.n88 256.663
R510 B.n804 B.n87 256.663
R511 B.n804 B.n86 256.663
R512 B.n804 B.n85 256.663
R513 B.n804 B.n84 256.663
R514 B.n804 B.n83 256.663
R515 B.n804 B.n82 256.663
R516 B.n804 B.n81 256.663
R517 B.n804 B.n80 256.663
R518 B.n804 B.n79 256.663
R519 B.n804 B.n78 256.663
R520 B.n804 B.n77 256.663
R521 B.n804 B.n76 256.663
R522 B.n804 B.n75 256.663
R523 B.n804 B.n74 256.663
R524 B.n804 B.n73 256.663
R525 B.n804 B.n72 256.663
R526 B.n804 B.n71 256.663
R527 B.n804 B.n70 256.663
R528 B.n804 B.n69 256.663
R529 B.n804 B.n68 256.663
R530 B.n804 B.n67 256.663
R531 B.n804 B.n66 256.663
R532 B.n804 B.n65 256.663
R533 B.n804 B.n64 256.663
R534 B.n804 B.n63 256.663
R535 B.n804 B.n62 256.663
R536 B.n804 B.n61 256.663
R537 B.n804 B.n60 256.663
R538 B.n804 B.n59 256.663
R539 B.n804 B.n58 256.663
R540 B.n804 B.n57 256.663
R541 B.n804 B.n56 256.663
R542 B.n804 B.n55 256.663
R543 B.n804 B.n54 256.663
R544 B.n804 B.n53 256.663
R545 B.n804 B.n52 256.663
R546 B.n804 B.n51 256.663
R547 B.n804 B.n50 256.663
R548 B.n804 B.n49 256.663
R549 B.n804 B.n48 256.663
R550 B.n455 B.n393 256.663
R551 B.n461 B.n393 256.663
R552 B.n463 B.n393 256.663
R553 B.n469 B.n393 256.663
R554 B.n471 B.n393 256.663
R555 B.n477 B.n393 256.663
R556 B.n479 B.n393 256.663
R557 B.n485 B.n393 256.663
R558 B.n487 B.n393 256.663
R559 B.n493 B.n393 256.663
R560 B.n495 B.n393 256.663
R561 B.n501 B.n393 256.663
R562 B.n503 B.n393 256.663
R563 B.n509 B.n393 256.663
R564 B.n511 B.n393 256.663
R565 B.n517 B.n393 256.663
R566 B.n519 B.n393 256.663
R567 B.n525 B.n393 256.663
R568 B.n527 B.n393 256.663
R569 B.n533 B.n393 256.663
R570 B.n535 B.n393 256.663
R571 B.n541 B.n393 256.663
R572 B.n543 B.n393 256.663
R573 B.n549 B.n393 256.663
R574 B.n551 B.n393 256.663
R575 B.n557 B.n393 256.663
R576 B.n559 B.n393 256.663
R577 B.n566 B.n393 256.663
R578 B.n568 B.n393 256.663
R579 B.n574 B.n393 256.663
R580 B.n576 B.n393 256.663
R581 B.n585 B.n393 256.663
R582 B.n587 B.n393 256.663
R583 B.n593 B.n393 256.663
R584 B.n595 B.n393 256.663
R585 B.n601 B.n393 256.663
R586 B.n603 B.n393 256.663
R587 B.n609 B.n393 256.663
R588 B.n611 B.n393 256.663
R589 B.n617 B.n393 256.663
R590 B.n619 B.n393 256.663
R591 B.n625 B.n393 256.663
R592 B.n627 B.n393 256.663
R593 B.n633 B.n393 256.663
R594 B.n635 B.n393 256.663
R595 B.n641 B.n393 256.663
R596 B.n643 B.n393 256.663
R597 B.n649 B.n393 256.663
R598 B.n651 B.n393 256.663
R599 B.n657 B.n393 256.663
R600 B.n659 B.n393 256.663
R601 B.n665 B.n393 256.663
R602 B.n667 B.n393 256.663
R603 B.n673 B.n393 256.663
R604 B.n675 B.n393 256.663
R605 B.n681 B.n393 256.663
R606 B.n683 B.n393 256.663
R607 B.n689 B.n393 256.663
R608 B.n691 B.n393 256.663
R609 B.n857 B.n856 256.663
R610 B.n115 B.n114 163.367
R611 B.n119 B.n118 163.367
R612 B.n123 B.n122 163.367
R613 B.n127 B.n126 163.367
R614 B.n131 B.n130 163.367
R615 B.n135 B.n134 163.367
R616 B.n139 B.n138 163.367
R617 B.n143 B.n142 163.367
R618 B.n147 B.n146 163.367
R619 B.n151 B.n150 163.367
R620 B.n155 B.n154 163.367
R621 B.n159 B.n158 163.367
R622 B.n163 B.n162 163.367
R623 B.n167 B.n166 163.367
R624 B.n171 B.n170 163.367
R625 B.n175 B.n174 163.367
R626 B.n179 B.n178 163.367
R627 B.n183 B.n182 163.367
R628 B.n187 B.n186 163.367
R629 B.n191 B.n190 163.367
R630 B.n195 B.n194 163.367
R631 B.n199 B.n198 163.367
R632 B.n203 B.n202 163.367
R633 B.n207 B.n206 163.367
R634 B.n211 B.n210 163.367
R635 B.n215 B.n214 163.367
R636 B.n219 B.n218 163.367
R637 B.n224 B.n223 163.367
R638 B.n228 B.n227 163.367
R639 B.n232 B.n231 163.367
R640 B.n236 B.n235 163.367
R641 B.n240 B.n239 163.367
R642 B.n244 B.n243 163.367
R643 B.n248 B.n247 163.367
R644 B.n252 B.n251 163.367
R645 B.n256 B.n255 163.367
R646 B.n260 B.n259 163.367
R647 B.n264 B.n263 163.367
R648 B.n268 B.n267 163.367
R649 B.n272 B.n271 163.367
R650 B.n276 B.n275 163.367
R651 B.n280 B.n279 163.367
R652 B.n284 B.n283 163.367
R653 B.n288 B.n287 163.367
R654 B.n292 B.n291 163.367
R655 B.n296 B.n295 163.367
R656 B.n300 B.n299 163.367
R657 B.n304 B.n303 163.367
R658 B.n308 B.n307 163.367
R659 B.n312 B.n311 163.367
R660 B.n316 B.n315 163.367
R661 B.n320 B.n319 163.367
R662 B.n324 B.n323 163.367
R663 B.n328 B.n327 163.367
R664 B.n332 B.n331 163.367
R665 B.n336 B.n335 163.367
R666 B.n340 B.n339 163.367
R667 B.n344 B.n343 163.367
R668 B.n803 B.n107 163.367
R669 B.n696 B.n388 163.367
R670 B.n704 B.n388 163.367
R671 B.n704 B.n386 163.367
R672 B.n708 B.n386 163.367
R673 B.n708 B.n380 163.367
R674 B.n716 B.n380 163.367
R675 B.n716 B.n378 163.367
R676 B.n720 B.n378 163.367
R677 B.n720 B.n372 163.367
R678 B.n728 B.n372 163.367
R679 B.n728 B.n370 163.367
R680 B.n732 B.n370 163.367
R681 B.n732 B.n364 163.367
R682 B.n740 B.n364 163.367
R683 B.n740 B.n362 163.367
R684 B.n744 B.n362 163.367
R685 B.n744 B.n356 163.367
R686 B.n752 B.n356 163.367
R687 B.n752 B.n354 163.367
R688 B.n757 B.n354 163.367
R689 B.n757 B.n348 163.367
R690 B.n765 B.n348 163.367
R691 B.n766 B.n765 163.367
R692 B.n766 B.n5 163.367
R693 B.n6 B.n5 163.367
R694 B.n7 B.n6 163.367
R695 B.n772 B.n7 163.367
R696 B.n774 B.n772 163.367
R697 B.n774 B.n12 163.367
R698 B.n13 B.n12 163.367
R699 B.n14 B.n13 163.367
R700 B.n779 B.n14 163.367
R701 B.n779 B.n19 163.367
R702 B.n20 B.n19 163.367
R703 B.n21 B.n20 163.367
R704 B.n784 B.n21 163.367
R705 B.n784 B.n26 163.367
R706 B.n27 B.n26 163.367
R707 B.n28 B.n27 163.367
R708 B.n789 B.n28 163.367
R709 B.n789 B.n33 163.367
R710 B.n34 B.n33 163.367
R711 B.n35 B.n34 163.367
R712 B.n794 B.n35 163.367
R713 B.n794 B.n40 163.367
R714 B.n41 B.n40 163.367
R715 B.n42 B.n41 163.367
R716 B.n799 B.n42 163.367
R717 B.n799 B.n47 163.367
R718 B.n456 B.n454 163.367
R719 B.n460 B.n454 163.367
R720 B.n464 B.n462 163.367
R721 B.n468 B.n452 163.367
R722 B.n472 B.n470 163.367
R723 B.n476 B.n450 163.367
R724 B.n480 B.n478 163.367
R725 B.n484 B.n448 163.367
R726 B.n488 B.n486 163.367
R727 B.n492 B.n446 163.367
R728 B.n496 B.n494 163.367
R729 B.n500 B.n444 163.367
R730 B.n504 B.n502 163.367
R731 B.n508 B.n442 163.367
R732 B.n512 B.n510 163.367
R733 B.n516 B.n440 163.367
R734 B.n520 B.n518 163.367
R735 B.n524 B.n438 163.367
R736 B.n528 B.n526 163.367
R737 B.n532 B.n436 163.367
R738 B.n536 B.n534 163.367
R739 B.n540 B.n434 163.367
R740 B.n544 B.n542 163.367
R741 B.n548 B.n432 163.367
R742 B.n552 B.n550 163.367
R743 B.n556 B.n430 163.367
R744 B.n560 B.n558 163.367
R745 B.n565 B.n426 163.367
R746 B.n569 B.n567 163.367
R747 B.n573 B.n424 163.367
R748 B.n577 B.n575 163.367
R749 B.n584 B.n422 163.367
R750 B.n588 B.n586 163.367
R751 B.n592 B.n420 163.367
R752 B.n596 B.n594 163.367
R753 B.n600 B.n418 163.367
R754 B.n604 B.n602 163.367
R755 B.n608 B.n416 163.367
R756 B.n612 B.n610 163.367
R757 B.n616 B.n414 163.367
R758 B.n620 B.n618 163.367
R759 B.n624 B.n412 163.367
R760 B.n628 B.n626 163.367
R761 B.n632 B.n410 163.367
R762 B.n636 B.n634 163.367
R763 B.n640 B.n408 163.367
R764 B.n644 B.n642 163.367
R765 B.n648 B.n406 163.367
R766 B.n652 B.n650 163.367
R767 B.n656 B.n404 163.367
R768 B.n660 B.n658 163.367
R769 B.n664 B.n402 163.367
R770 B.n668 B.n666 163.367
R771 B.n672 B.n400 163.367
R772 B.n676 B.n674 163.367
R773 B.n680 B.n398 163.367
R774 B.n684 B.n682 163.367
R775 B.n688 B.n396 163.367
R776 B.n692 B.n690 163.367
R777 B.n698 B.n390 163.367
R778 B.n702 B.n390 163.367
R779 B.n702 B.n384 163.367
R780 B.n710 B.n384 163.367
R781 B.n710 B.n382 163.367
R782 B.n714 B.n382 163.367
R783 B.n714 B.n376 163.367
R784 B.n722 B.n376 163.367
R785 B.n722 B.n374 163.367
R786 B.n726 B.n374 163.367
R787 B.n726 B.n368 163.367
R788 B.n734 B.n368 163.367
R789 B.n734 B.n366 163.367
R790 B.n738 B.n366 163.367
R791 B.n738 B.n360 163.367
R792 B.n746 B.n360 163.367
R793 B.n746 B.n358 163.367
R794 B.n750 B.n358 163.367
R795 B.n750 B.n352 163.367
R796 B.n759 B.n352 163.367
R797 B.n759 B.n350 163.367
R798 B.n763 B.n350 163.367
R799 B.n763 B.n3 163.367
R800 B.n855 B.n3 163.367
R801 B.n851 B.n2 163.367
R802 B.n851 B.n850 163.367
R803 B.n850 B.n9 163.367
R804 B.n846 B.n9 163.367
R805 B.n846 B.n11 163.367
R806 B.n842 B.n11 163.367
R807 B.n842 B.n16 163.367
R808 B.n838 B.n16 163.367
R809 B.n838 B.n18 163.367
R810 B.n834 B.n18 163.367
R811 B.n834 B.n23 163.367
R812 B.n830 B.n23 163.367
R813 B.n830 B.n25 163.367
R814 B.n826 B.n25 163.367
R815 B.n826 B.n30 163.367
R816 B.n822 B.n30 163.367
R817 B.n822 B.n32 163.367
R818 B.n818 B.n32 163.367
R819 B.n818 B.n37 163.367
R820 B.n814 B.n37 163.367
R821 B.n814 B.n39 163.367
R822 B.n810 B.n39 163.367
R823 B.n810 B.n44 163.367
R824 B.n806 B.n44 163.367
R825 B.n108 B.t16 105.169
R826 B.n580 B.t7 105.169
R827 B.n111 B.t10 105.147
R828 B.n427 B.t14 105.147
R829 B.n48 B.n46 71.676
R830 B.n115 B.n49 71.676
R831 B.n119 B.n50 71.676
R832 B.n123 B.n51 71.676
R833 B.n127 B.n52 71.676
R834 B.n131 B.n53 71.676
R835 B.n135 B.n54 71.676
R836 B.n139 B.n55 71.676
R837 B.n143 B.n56 71.676
R838 B.n147 B.n57 71.676
R839 B.n151 B.n58 71.676
R840 B.n155 B.n59 71.676
R841 B.n159 B.n60 71.676
R842 B.n163 B.n61 71.676
R843 B.n167 B.n62 71.676
R844 B.n171 B.n63 71.676
R845 B.n175 B.n64 71.676
R846 B.n179 B.n65 71.676
R847 B.n183 B.n66 71.676
R848 B.n187 B.n67 71.676
R849 B.n191 B.n68 71.676
R850 B.n195 B.n69 71.676
R851 B.n199 B.n70 71.676
R852 B.n203 B.n71 71.676
R853 B.n207 B.n72 71.676
R854 B.n211 B.n73 71.676
R855 B.n215 B.n74 71.676
R856 B.n219 B.n75 71.676
R857 B.n224 B.n76 71.676
R858 B.n228 B.n77 71.676
R859 B.n232 B.n78 71.676
R860 B.n236 B.n79 71.676
R861 B.n240 B.n80 71.676
R862 B.n244 B.n81 71.676
R863 B.n248 B.n82 71.676
R864 B.n252 B.n83 71.676
R865 B.n256 B.n84 71.676
R866 B.n260 B.n85 71.676
R867 B.n264 B.n86 71.676
R868 B.n268 B.n87 71.676
R869 B.n272 B.n88 71.676
R870 B.n276 B.n89 71.676
R871 B.n280 B.n90 71.676
R872 B.n284 B.n91 71.676
R873 B.n288 B.n92 71.676
R874 B.n292 B.n93 71.676
R875 B.n296 B.n94 71.676
R876 B.n300 B.n95 71.676
R877 B.n304 B.n96 71.676
R878 B.n308 B.n97 71.676
R879 B.n312 B.n98 71.676
R880 B.n316 B.n99 71.676
R881 B.n320 B.n100 71.676
R882 B.n324 B.n101 71.676
R883 B.n328 B.n102 71.676
R884 B.n332 B.n103 71.676
R885 B.n336 B.n104 71.676
R886 B.n340 B.n105 71.676
R887 B.n344 B.n106 71.676
R888 B.n107 B.n106 71.676
R889 B.n343 B.n105 71.676
R890 B.n339 B.n104 71.676
R891 B.n335 B.n103 71.676
R892 B.n331 B.n102 71.676
R893 B.n327 B.n101 71.676
R894 B.n323 B.n100 71.676
R895 B.n319 B.n99 71.676
R896 B.n315 B.n98 71.676
R897 B.n311 B.n97 71.676
R898 B.n307 B.n96 71.676
R899 B.n303 B.n95 71.676
R900 B.n299 B.n94 71.676
R901 B.n295 B.n93 71.676
R902 B.n291 B.n92 71.676
R903 B.n287 B.n91 71.676
R904 B.n283 B.n90 71.676
R905 B.n279 B.n89 71.676
R906 B.n275 B.n88 71.676
R907 B.n271 B.n87 71.676
R908 B.n267 B.n86 71.676
R909 B.n263 B.n85 71.676
R910 B.n259 B.n84 71.676
R911 B.n255 B.n83 71.676
R912 B.n251 B.n82 71.676
R913 B.n247 B.n81 71.676
R914 B.n243 B.n80 71.676
R915 B.n239 B.n79 71.676
R916 B.n235 B.n78 71.676
R917 B.n231 B.n77 71.676
R918 B.n227 B.n76 71.676
R919 B.n223 B.n75 71.676
R920 B.n218 B.n74 71.676
R921 B.n214 B.n73 71.676
R922 B.n210 B.n72 71.676
R923 B.n206 B.n71 71.676
R924 B.n202 B.n70 71.676
R925 B.n198 B.n69 71.676
R926 B.n194 B.n68 71.676
R927 B.n190 B.n67 71.676
R928 B.n186 B.n66 71.676
R929 B.n182 B.n65 71.676
R930 B.n178 B.n64 71.676
R931 B.n174 B.n63 71.676
R932 B.n170 B.n62 71.676
R933 B.n166 B.n61 71.676
R934 B.n162 B.n60 71.676
R935 B.n158 B.n59 71.676
R936 B.n154 B.n58 71.676
R937 B.n150 B.n57 71.676
R938 B.n146 B.n56 71.676
R939 B.n142 B.n55 71.676
R940 B.n138 B.n54 71.676
R941 B.n134 B.n53 71.676
R942 B.n130 B.n52 71.676
R943 B.n126 B.n51 71.676
R944 B.n122 B.n50 71.676
R945 B.n118 B.n49 71.676
R946 B.n114 B.n48 71.676
R947 B.n455 B.n392 71.676
R948 B.n461 B.n460 71.676
R949 B.n464 B.n463 71.676
R950 B.n469 B.n468 71.676
R951 B.n472 B.n471 71.676
R952 B.n477 B.n476 71.676
R953 B.n480 B.n479 71.676
R954 B.n485 B.n484 71.676
R955 B.n488 B.n487 71.676
R956 B.n493 B.n492 71.676
R957 B.n496 B.n495 71.676
R958 B.n501 B.n500 71.676
R959 B.n504 B.n503 71.676
R960 B.n509 B.n508 71.676
R961 B.n512 B.n511 71.676
R962 B.n517 B.n516 71.676
R963 B.n520 B.n519 71.676
R964 B.n525 B.n524 71.676
R965 B.n528 B.n527 71.676
R966 B.n533 B.n532 71.676
R967 B.n536 B.n535 71.676
R968 B.n541 B.n540 71.676
R969 B.n544 B.n543 71.676
R970 B.n549 B.n548 71.676
R971 B.n552 B.n551 71.676
R972 B.n557 B.n556 71.676
R973 B.n560 B.n559 71.676
R974 B.n566 B.n565 71.676
R975 B.n569 B.n568 71.676
R976 B.n574 B.n573 71.676
R977 B.n577 B.n576 71.676
R978 B.n585 B.n584 71.676
R979 B.n588 B.n587 71.676
R980 B.n593 B.n592 71.676
R981 B.n596 B.n595 71.676
R982 B.n601 B.n600 71.676
R983 B.n604 B.n603 71.676
R984 B.n609 B.n608 71.676
R985 B.n612 B.n611 71.676
R986 B.n617 B.n616 71.676
R987 B.n620 B.n619 71.676
R988 B.n625 B.n624 71.676
R989 B.n628 B.n627 71.676
R990 B.n633 B.n632 71.676
R991 B.n636 B.n635 71.676
R992 B.n641 B.n640 71.676
R993 B.n644 B.n643 71.676
R994 B.n649 B.n648 71.676
R995 B.n652 B.n651 71.676
R996 B.n657 B.n656 71.676
R997 B.n660 B.n659 71.676
R998 B.n665 B.n664 71.676
R999 B.n668 B.n667 71.676
R1000 B.n673 B.n672 71.676
R1001 B.n676 B.n675 71.676
R1002 B.n681 B.n680 71.676
R1003 B.n684 B.n683 71.676
R1004 B.n689 B.n688 71.676
R1005 B.n692 B.n691 71.676
R1006 B.n456 B.n455 71.676
R1007 B.n462 B.n461 71.676
R1008 B.n463 B.n452 71.676
R1009 B.n470 B.n469 71.676
R1010 B.n471 B.n450 71.676
R1011 B.n478 B.n477 71.676
R1012 B.n479 B.n448 71.676
R1013 B.n486 B.n485 71.676
R1014 B.n487 B.n446 71.676
R1015 B.n494 B.n493 71.676
R1016 B.n495 B.n444 71.676
R1017 B.n502 B.n501 71.676
R1018 B.n503 B.n442 71.676
R1019 B.n510 B.n509 71.676
R1020 B.n511 B.n440 71.676
R1021 B.n518 B.n517 71.676
R1022 B.n519 B.n438 71.676
R1023 B.n526 B.n525 71.676
R1024 B.n527 B.n436 71.676
R1025 B.n534 B.n533 71.676
R1026 B.n535 B.n434 71.676
R1027 B.n542 B.n541 71.676
R1028 B.n543 B.n432 71.676
R1029 B.n550 B.n549 71.676
R1030 B.n551 B.n430 71.676
R1031 B.n558 B.n557 71.676
R1032 B.n559 B.n426 71.676
R1033 B.n567 B.n566 71.676
R1034 B.n568 B.n424 71.676
R1035 B.n575 B.n574 71.676
R1036 B.n576 B.n422 71.676
R1037 B.n586 B.n585 71.676
R1038 B.n587 B.n420 71.676
R1039 B.n594 B.n593 71.676
R1040 B.n595 B.n418 71.676
R1041 B.n602 B.n601 71.676
R1042 B.n603 B.n416 71.676
R1043 B.n610 B.n609 71.676
R1044 B.n611 B.n414 71.676
R1045 B.n618 B.n617 71.676
R1046 B.n619 B.n412 71.676
R1047 B.n626 B.n625 71.676
R1048 B.n627 B.n410 71.676
R1049 B.n634 B.n633 71.676
R1050 B.n635 B.n408 71.676
R1051 B.n642 B.n641 71.676
R1052 B.n643 B.n406 71.676
R1053 B.n650 B.n649 71.676
R1054 B.n651 B.n404 71.676
R1055 B.n658 B.n657 71.676
R1056 B.n659 B.n402 71.676
R1057 B.n666 B.n665 71.676
R1058 B.n667 B.n400 71.676
R1059 B.n674 B.n673 71.676
R1060 B.n675 B.n398 71.676
R1061 B.n682 B.n681 71.676
R1062 B.n683 B.n396 71.676
R1063 B.n690 B.n689 71.676
R1064 B.n691 B.n394 71.676
R1065 B.n856 B.n855 71.676
R1066 B.n856 B.n2 71.676
R1067 B.n109 B.t17 69.4848
R1068 B.n581 B.t6 69.4848
R1069 B.n112 B.t11 69.4631
R1070 B.n428 B.t13 69.4631
R1071 B.n221 B.n112 59.5399
R1072 B.n110 B.n109 59.5399
R1073 B.n582 B.n581 59.5399
R1074 B.n563 B.n428 59.5399
R1075 B.n697 B.n393 57.2684
R1076 B.n805 B.n804 57.2684
R1077 B.n112 B.n111 35.6853
R1078 B.n109 B.n108 35.6853
R1079 B.n581 B.n580 35.6853
R1080 B.n428 B.n427 35.6853
R1081 B.n697 B.n389 34.4626
R1082 B.n703 B.n389 34.4626
R1083 B.n703 B.n385 34.4626
R1084 B.n709 B.n385 34.4626
R1085 B.n709 B.n381 34.4626
R1086 B.n715 B.n381 34.4626
R1087 B.n721 B.n377 34.4626
R1088 B.n721 B.n373 34.4626
R1089 B.n727 B.n373 34.4626
R1090 B.n727 B.n369 34.4626
R1091 B.n733 B.n369 34.4626
R1092 B.n733 B.n365 34.4626
R1093 B.n739 B.n365 34.4626
R1094 B.n745 B.n361 34.4626
R1095 B.n745 B.n357 34.4626
R1096 B.n751 B.n357 34.4626
R1097 B.n751 B.n353 34.4626
R1098 B.n758 B.n353 34.4626
R1099 B.n764 B.n349 34.4626
R1100 B.n764 B.n4 34.4626
R1101 B.n854 B.n4 34.4626
R1102 B.n854 B.n853 34.4626
R1103 B.n853 B.n852 34.4626
R1104 B.n852 B.n8 34.4626
R1105 B.n773 B.n8 34.4626
R1106 B.n845 B.n844 34.4626
R1107 B.n844 B.n843 34.4626
R1108 B.n843 B.n15 34.4626
R1109 B.n837 B.n15 34.4626
R1110 B.n837 B.n836 34.4626
R1111 B.n835 B.n22 34.4626
R1112 B.n829 B.n22 34.4626
R1113 B.n829 B.n828 34.4626
R1114 B.n828 B.n827 34.4626
R1115 B.n827 B.n29 34.4626
R1116 B.n821 B.n29 34.4626
R1117 B.n821 B.n820 34.4626
R1118 B.n819 B.n36 34.4626
R1119 B.n813 B.n36 34.4626
R1120 B.n813 B.n812 34.4626
R1121 B.n812 B.n811 34.4626
R1122 B.n811 B.n43 34.4626
R1123 B.n805 B.n43 34.4626
R1124 B.n699 B.n391 30.1273
R1125 B.n695 B.n694 30.1273
R1126 B.n802 B.n801 30.1273
R1127 B.n807 B.n45 30.1273
R1128 B.t5 B.n377 28.8879
R1129 B.n820 B.t9 28.8879
R1130 B.t3 B.n349 27.8743
R1131 B.n773 B.t2 27.8743
R1132 B.n739 B.t0 26.8607
R1133 B.t1 B.n835 26.8607
R1134 B B.n857 18.0485
R1135 B.n700 B.n699 10.6151
R1136 B.n701 B.n700 10.6151
R1137 B.n701 B.n383 10.6151
R1138 B.n711 B.n383 10.6151
R1139 B.n712 B.n711 10.6151
R1140 B.n713 B.n712 10.6151
R1141 B.n713 B.n375 10.6151
R1142 B.n723 B.n375 10.6151
R1143 B.n724 B.n723 10.6151
R1144 B.n725 B.n724 10.6151
R1145 B.n725 B.n367 10.6151
R1146 B.n735 B.n367 10.6151
R1147 B.n736 B.n735 10.6151
R1148 B.n737 B.n736 10.6151
R1149 B.n737 B.n359 10.6151
R1150 B.n747 B.n359 10.6151
R1151 B.n748 B.n747 10.6151
R1152 B.n749 B.n748 10.6151
R1153 B.n749 B.n351 10.6151
R1154 B.n760 B.n351 10.6151
R1155 B.n761 B.n760 10.6151
R1156 B.n762 B.n761 10.6151
R1157 B.n762 B.n0 10.6151
R1158 B.n457 B.n391 10.6151
R1159 B.n458 B.n457 10.6151
R1160 B.n459 B.n458 10.6151
R1161 B.n459 B.n453 10.6151
R1162 B.n465 B.n453 10.6151
R1163 B.n466 B.n465 10.6151
R1164 B.n467 B.n466 10.6151
R1165 B.n467 B.n451 10.6151
R1166 B.n473 B.n451 10.6151
R1167 B.n474 B.n473 10.6151
R1168 B.n475 B.n474 10.6151
R1169 B.n475 B.n449 10.6151
R1170 B.n481 B.n449 10.6151
R1171 B.n482 B.n481 10.6151
R1172 B.n483 B.n482 10.6151
R1173 B.n483 B.n447 10.6151
R1174 B.n489 B.n447 10.6151
R1175 B.n490 B.n489 10.6151
R1176 B.n491 B.n490 10.6151
R1177 B.n491 B.n445 10.6151
R1178 B.n497 B.n445 10.6151
R1179 B.n498 B.n497 10.6151
R1180 B.n499 B.n498 10.6151
R1181 B.n499 B.n443 10.6151
R1182 B.n505 B.n443 10.6151
R1183 B.n506 B.n505 10.6151
R1184 B.n507 B.n506 10.6151
R1185 B.n507 B.n441 10.6151
R1186 B.n513 B.n441 10.6151
R1187 B.n514 B.n513 10.6151
R1188 B.n515 B.n514 10.6151
R1189 B.n515 B.n439 10.6151
R1190 B.n521 B.n439 10.6151
R1191 B.n522 B.n521 10.6151
R1192 B.n523 B.n522 10.6151
R1193 B.n523 B.n437 10.6151
R1194 B.n529 B.n437 10.6151
R1195 B.n530 B.n529 10.6151
R1196 B.n531 B.n530 10.6151
R1197 B.n531 B.n435 10.6151
R1198 B.n537 B.n435 10.6151
R1199 B.n538 B.n537 10.6151
R1200 B.n539 B.n538 10.6151
R1201 B.n539 B.n433 10.6151
R1202 B.n545 B.n433 10.6151
R1203 B.n546 B.n545 10.6151
R1204 B.n547 B.n546 10.6151
R1205 B.n547 B.n431 10.6151
R1206 B.n553 B.n431 10.6151
R1207 B.n554 B.n553 10.6151
R1208 B.n555 B.n554 10.6151
R1209 B.n555 B.n429 10.6151
R1210 B.n561 B.n429 10.6151
R1211 B.n562 B.n561 10.6151
R1212 B.n564 B.n425 10.6151
R1213 B.n570 B.n425 10.6151
R1214 B.n571 B.n570 10.6151
R1215 B.n572 B.n571 10.6151
R1216 B.n572 B.n423 10.6151
R1217 B.n578 B.n423 10.6151
R1218 B.n579 B.n578 10.6151
R1219 B.n583 B.n579 10.6151
R1220 B.n589 B.n421 10.6151
R1221 B.n590 B.n589 10.6151
R1222 B.n591 B.n590 10.6151
R1223 B.n591 B.n419 10.6151
R1224 B.n597 B.n419 10.6151
R1225 B.n598 B.n597 10.6151
R1226 B.n599 B.n598 10.6151
R1227 B.n599 B.n417 10.6151
R1228 B.n605 B.n417 10.6151
R1229 B.n606 B.n605 10.6151
R1230 B.n607 B.n606 10.6151
R1231 B.n607 B.n415 10.6151
R1232 B.n613 B.n415 10.6151
R1233 B.n614 B.n613 10.6151
R1234 B.n615 B.n614 10.6151
R1235 B.n615 B.n413 10.6151
R1236 B.n621 B.n413 10.6151
R1237 B.n622 B.n621 10.6151
R1238 B.n623 B.n622 10.6151
R1239 B.n623 B.n411 10.6151
R1240 B.n629 B.n411 10.6151
R1241 B.n630 B.n629 10.6151
R1242 B.n631 B.n630 10.6151
R1243 B.n631 B.n409 10.6151
R1244 B.n637 B.n409 10.6151
R1245 B.n638 B.n637 10.6151
R1246 B.n639 B.n638 10.6151
R1247 B.n639 B.n407 10.6151
R1248 B.n645 B.n407 10.6151
R1249 B.n646 B.n645 10.6151
R1250 B.n647 B.n646 10.6151
R1251 B.n647 B.n405 10.6151
R1252 B.n653 B.n405 10.6151
R1253 B.n654 B.n653 10.6151
R1254 B.n655 B.n654 10.6151
R1255 B.n655 B.n403 10.6151
R1256 B.n661 B.n403 10.6151
R1257 B.n662 B.n661 10.6151
R1258 B.n663 B.n662 10.6151
R1259 B.n663 B.n401 10.6151
R1260 B.n669 B.n401 10.6151
R1261 B.n670 B.n669 10.6151
R1262 B.n671 B.n670 10.6151
R1263 B.n671 B.n399 10.6151
R1264 B.n677 B.n399 10.6151
R1265 B.n678 B.n677 10.6151
R1266 B.n679 B.n678 10.6151
R1267 B.n679 B.n397 10.6151
R1268 B.n685 B.n397 10.6151
R1269 B.n686 B.n685 10.6151
R1270 B.n687 B.n686 10.6151
R1271 B.n687 B.n395 10.6151
R1272 B.n693 B.n395 10.6151
R1273 B.n694 B.n693 10.6151
R1274 B.n695 B.n387 10.6151
R1275 B.n705 B.n387 10.6151
R1276 B.n706 B.n705 10.6151
R1277 B.n707 B.n706 10.6151
R1278 B.n707 B.n379 10.6151
R1279 B.n717 B.n379 10.6151
R1280 B.n718 B.n717 10.6151
R1281 B.n719 B.n718 10.6151
R1282 B.n719 B.n371 10.6151
R1283 B.n729 B.n371 10.6151
R1284 B.n730 B.n729 10.6151
R1285 B.n731 B.n730 10.6151
R1286 B.n731 B.n363 10.6151
R1287 B.n741 B.n363 10.6151
R1288 B.n742 B.n741 10.6151
R1289 B.n743 B.n742 10.6151
R1290 B.n743 B.n355 10.6151
R1291 B.n753 B.n355 10.6151
R1292 B.n754 B.n753 10.6151
R1293 B.n756 B.n754 10.6151
R1294 B.n756 B.n755 10.6151
R1295 B.n755 B.n347 10.6151
R1296 B.n767 B.n347 10.6151
R1297 B.n768 B.n767 10.6151
R1298 B.n769 B.n768 10.6151
R1299 B.n770 B.n769 10.6151
R1300 B.n771 B.n770 10.6151
R1301 B.n775 B.n771 10.6151
R1302 B.n776 B.n775 10.6151
R1303 B.n777 B.n776 10.6151
R1304 B.n778 B.n777 10.6151
R1305 B.n780 B.n778 10.6151
R1306 B.n781 B.n780 10.6151
R1307 B.n782 B.n781 10.6151
R1308 B.n783 B.n782 10.6151
R1309 B.n785 B.n783 10.6151
R1310 B.n786 B.n785 10.6151
R1311 B.n787 B.n786 10.6151
R1312 B.n788 B.n787 10.6151
R1313 B.n790 B.n788 10.6151
R1314 B.n791 B.n790 10.6151
R1315 B.n792 B.n791 10.6151
R1316 B.n793 B.n792 10.6151
R1317 B.n795 B.n793 10.6151
R1318 B.n796 B.n795 10.6151
R1319 B.n797 B.n796 10.6151
R1320 B.n798 B.n797 10.6151
R1321 B.n800 B.n798 10.6151
R1322 B.n801 B.n800 10.6151
R1323 B.n849 B.n1 10.6151
R1324 B.n849 B.n848 10.6151
R1325 B.n848 B.n847 10.6151
R1326 B.n847 B.n10 10.6151
R1327 B.n841 B.n10 10.6151
R1328 B.n841 B.n840 10.6151
R1329 B.n840 B.n839 10.6151
R1330 B.n839 B.n17 10.6151
R1331 B.n833 B.n17 10.6151
R1332 B.n833 B.n832 10.6151
R1333 B.n832 B.n831 10.6151
R1334 B.n831 B.n24 10.6151
R1335 B.n825 B.n24 10.6151
R1336 B.n825 B.n824 10.6151
R1337 B.n824 B.n823 10.6151
R1338 B.n823 B.n31 10.6151
R1339 B.n817 B.n31 10.6151
R1340 B.n817 B.n816 10.6151
R1341 B.n816 B.n815 10.6151
R1342 B.n815 B.n38 10.6151
R1343 B.n809 B.n38 10.6151
R1344 B.n809 B.n808 10.6151
R1345 B.n808 B.n807 10.6151
R1346 B.n113 B.n45 10.6151
R1347 B.n116 B.n113 10.6151
R1348 B.n117 B.n116 10.6151
R1349 B.n120 B.n117 10.6151
R1350 B.n121 B.n120 10.6151
R1351 B.n124 B.n121 10.6151
R1352 B.n125 B.n124 10.6151
R1353 B.n128 B.n125 10.6151
R1354 B.n129 B.n128 10.6151
R1355 B.n132 B.n129 10.6151
R1356 B.n133 B.n132 10.6151
R1357 B.n136 B.n133 10.6151
R1358 B.n137 B.n136 10.6151
R1359 B.n140 B.n137 10.6151
R1360 B.n141 B.n140 10.6151
R1361 B.n144 B.n141 10.6151
R1362 B.n145 B.n144 10.6151
R1363 B.n148 B.n145 10.6151
R1364 B.n149 B.n148 10.6151
R1365 B.n152 B.n149 10.6151
R1366 B.n153 B.n152 10.6151
R1367 B.n156 B.n153 10.6151
R1368 B.n157 B.n156 10.6151
R1369 B.n160 B.n157 10.6151
R1370 B.n161 B.n160 10.6151
R1371 B.n164 B.n161 10.6151
R1372 B.n165 B.n164 10.6151
R1373 B.n168 B.n165 10.6151
R1374 B.n169 B.n168 10.6151
R1375 B.n172 B.n169 10.6151
R1376 B.n173 B.n172 10.6151
R1377 B.n176 B.n173 10.6151
R1378 B.n177 B.n176 10.6151
R1379 B.n180 B.n177 10.6151
R1380 B.n181 B.n180 10.6151
R1381 B.n184 B.n181 10.6151
R1382 B.n185 B.n184 10.6151
R1383 B.n188 B.n185 10.6151
R1384 B.n189 B.n188 10.6151
R1385 B.n192 B.n189 10.6151
R1386 B.n193 B.n192 10.6151
R1387 B.n196 B.n193 10.6151
R1388 B.n197 B.n196 10.6151
R1389 B.n200 B.n197 10.6151
R1390 B.n201 B.n200 10.6151
R1391 B.n204 B.n201 10.6151
R1392 B.n205 B.n204 10.6151
R1393 B.n208 B.n205 10.6151
R1394 B.n209 B.n208 10.6151
R1395 B.n212 B.n209 10.6151
R1396 B.n213 B.n212 10.6151
R1397 B.n216 B.n213 10.6151
R1398 B.n217 B.n216 10.6151
R1399 B.n220 B.n217 10.6151
R1400 B.n225 B.n222 10.6151
R1401 B.n226 B.n225 10.6151
R1402 B.n229 B.n226 10.6151
R1403 B.n230 B.n229 10.6151
R1404 B.n233 B.n230 10.6151
R1405 B.n234 B.n233 10.6151
R1406 B.n237 B.n234 10.6151
R1407 B.n238 B.n237 10.6151
R1408 B.n242 B.n241 10.6151
R1409 B.n245 B.n242 10.6151
R1410 B.n246 B.n245 10.6151
R1411 B.n249 B.n246 10.6151
R1412 B.n250 B.n249 10.6151
R1413 B.n253 B.n250 10.6151
R1414 B.n254 B.n253 10.6151
R1415 B.n257 B.n254 10.6151
R1416 B.n258 B.n257 10.6151
R1417 B.n261 B.n258 10.6151
R1418 B.n262 B.n261 10.6151
R1419 B.n265 B.n262 10.6151
R1420 B.n266 B.n265 10.6151
R1421 B.n269 B.n266 10.6151
R1422 B.n270 B.n269 10.6151
R1423 B.n273 B.n270 10.6151
R1424 B.n274 B.n273 10.6151
R1425 B.n277 B.n274 10.6151
R1426 B.n278 B.n277 10.6151
R1427 B.n281 B.n278 10.6151
R1428 B.n282 B.n281 10.6151
R1429 B.n285 B.n282 10.6151
R1430 B.n286 B.n285 10.6151
R1431 B.n289 B.n286 10.6151
R1432 B.n290 B.n289 10.6151
R1433 B.n293 B.n290 10.6151
R1434 B.n294 B.n293 10.6151
R1435 B.n297 B.n294 10.6151
R1436 B.n298 B.n297 10.6151
R1437 B.n301 B.n298 10.6151
R1438 B.n302 B.n301 10.6151
R1439 B.n305 B.n302 10.6151
R1440 B.n306 B.n305 10.6151
R1441 B.n309 B.n306 10.6151
R1442 B.n310 B.n309 10.6151
R1443 B.n313 B.n310 10.6151
R1444 B.n314 B.n313 10.6151
R1445 B.n317 B.n314 10.6151
R1446 B.n318 B.n317 10.6151
R1447 B.n321 B.n318 10.6151
R1448 B.n322 B.n321 10.6151
R1449 B.n325 B.n322 10.6151
R1450 B.n326 B.n325 10.6151
R1451 B.n329 B.n326 10.6151
R1452 B.n330 B.n329 10.6151
R1453 B.n333 B.n330 10.6151
R1454 B.n334 B.n333 10.6151
R1455 B.n337 B.n334 10.6151
R1456 B.n338 B.n337 10.6151
R1457 B.n341 B.n338 10.6151
R1458 B.n342 B.n341 10.6151
R1459 B.n345 B.n342 10.6151
R1460 B.n346 B.n345 10.6151
R1461 B.n802 B.n346 10.6151
R1462 B.n857 B.n0 8.11757
R1463 B.n857 B.n1 8.11757
R1464 B.t0 B.n361 7.60243
R1465 B.n836 B.t1 7.60243
R1466 B.n758 B.t3 6.58884
R1467 B.n845 B.t2 6.58884
R1468 B.n564 B.n563 6.5566
R1469 B.n583 B.n582 6.5566
R1470 B.n222 B.n221 6.5566
R1471 B.n238 B.n110 6.5566
R1472 B.n715 B.t5 5.57525
R1473 B.t9 B.n819 5.57525
R1474 B.n563 B.n562 4.05904
R1475 B.n582 B.n421 4.05904
R1476 B.n221 B.n220 4.05904
R1477 B.n241 B.n110 4.05904
R1478 VN.n0 VN.t1 298.733
R1479 VN.n1 VN.t2 298.733
R1480 VN.n0 VN.t0 298.416
R1481 VN.n1 VN.t3 298.416
R1482 VN VN.n1 59.6237
R1483 VN VN.n0 13.029
R1484 VDD2.n2 VDD2.n0 103.192
R1485 VDD2.n2 VDD2.n1 60.5555
R1486 VDD2.n1 VDD2.t0 1.20561
R1487 VDD2.n1 VDD2.t1 1.20561
R1488 VDD2.n0 VDD2.t2 1.20561
R1489 VDD2.n0 VDD2.t3 1.20561
R1490 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 5.80471f
C1 VDD1 VTAIL 6.85795f
C2 VP VN 6.22654f
C3 VN VTAIL 5.19593f
C4 VP VTAIL 5.21003f
C5 VDD2 VDD1 0.76218f
C6 VDD2 VN 5.62825f
C7 VDD1 VN 0.148133f
C8 VDD2 VP 0.325065f
C9 VDD2 VTAIL 6.90485f
C10 VDD2 B 3.501921f
C11 VDD1 B 7.76584f
C12 VTAIL B 12.01322f
C13 VN B 9.30397f
C14 VP B 6.90754f
C15 VDD2.t2 B 0.34487f
C16 VDD2.t3 B 0.34487f
C17 VDD2.n0 B 3.90611f
C18 VDD2.t0 B 0.34487f
C19 VDD2.t1 B 0.34487f
C20 VDD2.n1 B 3.12954f
C21 VDD2.n2 B 3.94339f
C22 VN.t1 B 2.44447f
C23 VN.t0 B 2.44342f
C24 VN.n0 B 1.73883f
C25 VN.t2 B 2.44447f
C26 VN.t3 B 2.44342f
C27 VN.n1 B 3.19247f
C28 VTAIL.t2 B 2.23617f
C29 VTAIL.n0 B 0.27322f
C30 VTAIL.t6 B 2.23617f
C31 VTAIL.n1 B 0.309368f
C32 VTAIL.t7 B 2.23617f
C33 VTAIL.n2 B 1.2683f
C34 VTAIL.t0 B 2.23617f
C35 VTAIL.n3 B 1.26829f
C36 VTAIL.t3 B 2.23617f
C37 VTAIL.n4 B 0.309365f
C38 VTAIL.t4 B 2.23617f
C39 VTAIL.n5 B 0.309365f
C40 VTAIL.t5 B 2.23617f
C41 VTAIL.n6 B 1.2683f
C42 VTAIL.t1 B 2.23617f
C43 VTAIL.n7 B 1.22642f
C44 VDD1.t0 B 0.34766f
C45 VDD1.t3 B 0.34766f
C46 VDD1.n0 B 3.15521f
C47 VDD1.t1 B 0.34766f
C48 VDD1.t2 B 0.34766f
C49 VDD1.n1 B 3.96552f
C50 VP.n0 B 0.034662f
C51 VP.t1 B 2.36105f
C52 VP.n1 B 0.0506f
C53 VP.t3 B 2.48023f
C54 VP.t2 B 2.47917f
C55 VP.n2 B 3.21887f
C56 VP.n3 B 2.11487f
C57 VP.t0 B 2.36105f
C58 VP.n4 B 0.904367f
C59 VP.n5 B 0.043551f
C60 VP.n6 B 0.034662f
C61 VP.n7 B 0.034662f
C62 VP.n8 B 0.034662f
C63 VP.n9 B 0.0506f
C64 VP.n10 B 0.043551f
C65 VP.n11 B 0.904367f
C66 VP.n12 B 0.033785f
.ends

