* NGSPICE file created from diff_pair_sample_0809.ext - technology: sky130A

.subckt diff_pair_sample_0809 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=5.9826 ps=31.46 w=15.34 l=3.01
X1 B.t11 B.t9 B.t10 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.01
X2 B.t8 B.t6 B.t7 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.01
X3 B.t5 B.t3 B.t4 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.01
X4 B.t2 B.t0 B.t1 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.01
X5 VDD1.t1 VP.t0 VTAIL.t0 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=5.9826 ps=31.46 w=15.34 l=3.01
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=5.9826 ps=31.46 w=15.34 l=3.01
X7 VDD2.t0 VN.t1 VTAIL.t3 w_n2306_n4036# sky130_fd_pr__pfet_01v8 ad=5.9826 pd=31.46 as=5.9826 ps=31.46 w=15.34 l=3.01
R0 VN VN.t0 212.237
R1 VN VN.t1 164.392
R2 VTAIL.n338 VTAIL.n258 756.745
R3 VTAIL.n80 VTAIL.n0 756.745
R4 VTAIL.n252 VTAIL.n172 756.745
R5 VTAIL.n166 VTAIL.n86 756.745
R6 VTAIL.n287 VTAIL.n286 585
R7 VTAIL.n289 VTAIL.n288 585
R8 VTAIL.n282 VTAIL.n281 585
R9 VTAIL.n295 VTAIL.n294 585
R10 VTAIL.n297 VTAIL.n296 585
R11 VTAIL.n278 VTAIL.n277 585
R12 VTAIL.n303 VTAIL.n302 585
R13 VTAIL.n305 VTAIL.n304 585
R14 VTAIL.n274 VTAIL.n273 585
R15 VTAIL.n311 VTAIL.n310 585
R16 VTAIL.n313 VTAIL.n312 585
R17 VTAIL.n270 VTAIL.n269 585
R18 VTAIL.n319 VTAIL.n318 585
R19 VTAIL.n321 VTAIL.n320 585
R20 VTAIL.n266 VTAIL.n265 585
R21 VTAIL.n328 VTAIL.n327 585
R22 VTAIL.n329 VTAIL.n264 585
R23 VTAIL.n331 VTAIL.n330 585
R24 VTAIL.n262 VTAIL.n261 585
R25 VTAIL.n337 VTAIL.n336 585
R26 VTAIL.n339 VTAIL.n338 585
R27 VTAIL.n29 VTAIL.n28 585
R28 VTAIL.n31 VTAIL.n30 585
R29 VTAIL.n24 VTAIL.n23 585
R30 VTAIL.n37 VTAIL.n36 585
R31 VTAIL.n39 VTAIL.n38 585
R32 VTAIL.n20 VTAIL.n19 585
R33 VTAIL.n45 VTAIL.n44 585
R34 VTAIL.n47 VTAIL.n46 585
R35 VTAIL.n16 VTAIL.n15 585
R36 VTAIL.n53 VTAIL.n52 585
R37 VTAIL.n55 VTAIL.n54 585
R38 VTAIL.n12 VTAIL.n11 585
R39 VTAIL.n61 VTAIL.n60 585
R40 VTAIL.n63 VTAIL.n62 585
R41 VTAIL.n8 VTAIL.n7 585
R42 VTAIL.n70 VTAIL.n69 585
R43 VTAIL.n71 VTAIL.n6 585
R44 VTAIL.n73 VTAIL.n72 585
R45 VTAIL.n4 VTAIL.n3 585
R46 VTAIL.n79 VTAIL.n78 585
R47 VTAIL.n81 VTAIL.n80 585
R48 VTAIL.n253 VTAIL.n252 585
R49 VTAIL.n251 VTAIL.n250 585
R50 VTAIL.n176 VTAIL.n175 585
R51 VTAIL.n180 VTAIL.n178 585
R52 VTAIL.n245 VTAIL.n244 585
R53 VTAIL.n243 VTAIL.n242 585
R54 VTAIL.n182 VTAIL.n181 585
R55 VTAIL.n237 VTAIL.n236 585
R56 VTAIL.n235 VTAIL.n234 585
R57 VTAIL.n186 VTAIL.n185 585
R58 VTAIL.n229 VTAIL.n228 585
R59 VTAIL.n227 VTAIL.n226 585
R60 VTAIL.n190 VTAIL.n189 585
R61 VTAIL.n221 VTAIL.n220 585
R62 VTAIL.n219 VTAIL.n218 585
R63 VTAIL.n194 VTAIL.n193 585
R64 VTAIL.n213 VTAIL.n212 585
R65 VTAIL.n211 VTAIL.n210 585
R66 VTAIL.n198 VTAIL.n197 585
R67 VTAIL.n205 VTAIL.n204 585
R68 VTAIL.n203 VTAIL.n202 585
R69 VTAIL.n167 VTAIL.n166 585
R70 VTAIL.n165 VTAIL.n164 585
R71 VTAIL.n90 VTAIL.n89 585
R72 VTAIL.n94 VTAIL.n92 585
R73 VTAIL.n159 VTAIL.n158 585
R74 VTAIL.n157 VTAIL.n156 585
R75 VTAIL.n96 VTAIL.n95 585
R76 VTAIL.n151 VTAIL.n150 585
R77 VTAIL.n149 VTAIL.n148 585
R78 VTAIL.n100 VTAIL.n99 585
R79 VTAIL.n143 VTAIL.n142 585
R80 VTAIL.n141 VTAIL.n140 585
R81 VTAIL.n104 VTAIL.n103 585
R82 VTAIL.n135 VTAIL.n134 585
R83 VTAIL.n133 VTAIL.n132 585
R84 VTAIL.n108 VTAIL.n107 585
R85 VTAIL.n127 VTAIL.n126 585
R86 VTAIL.n125 VTAIL.n124 585
R87 VTAIL.n112 VTAIL.n111 585
R88 VTAIL.n119 VTAIL.n118 585
R89 VTAIL.n117 VTAIL.n116 585
R90 VTAIL.n285 VTAIL.t3 327.466
R91 VTAIL.n27 VTAIL.t0 327.466
R92 VTAIL.n201 VTAIL.t1 327.466
R93 VTAIL.n115 VTAIL.t2 327.466
R94 VTAIL.n288 VTAIL.n287 171.744
R95 VTAIL.n288 VTAIL.n281 171.744
R96 VTAIL.n295 VTAIL.n281 171.744
R97 VTAIL.n296 VTAIL.n295 171.744
R98 VTAIL.n296 VTAIL.n277 171.744
R99 VTAIL.n303 VTAIL.n277 171.744
R100 VTAIL.n304 VTAIL.n303 171.744
R101 VTAIL.n304 VTAIL.n273 171.744
R102 VTAIL.n311 VTAIL.n273 171.744
R103 VTAIL.n312 VTAIL.n311 171.744
R104 VTAIL.n312 VTAIL.n269 171.744
R105 VTAIL.n319 VTAIL.n269 171.744
R106 VTAIL.n320 VTAIL.n319 171.744
R107 VTAIL.n320 VTAIL.n265 171.744
R108 VTAIL.n328 VTAIL.n265 171.744
R109 VTAIL.n329 VTAIL.n328 171.744
R110 VTAIL.n330 VTAIL.n329 171.744
R111 VTAIL.n330 VTAIL.n261 171.744
R112 VTAIL.n337 VTAIL.n261 171.744
R113 VTAIL.n338 VTAIL.n337 171.744
R114 VTAIL.n30 VTAIL.n29 171.744
R115 VTAIL.n30 VTAIL.n23 171.744
R116 VTAIL.n37 VTAIL.n23 171.744
R117 VTAIL.n38 VTAIL.n37 171.744
R118 VTAIL.n38 VTAIL.n19 171.744
R119 VTAIL.n45 VTAIL.n19 171.744
R120 VTAIL.n46 VTAIL.n45 171.744
R121 VTAIL.n46 VTAIL.n15 171.744
R122 VTAIL.n53 VTAIL.n15 171.744
R123 VTAIL.n54 VTAIL.n53 171.744
R124 VTAIL.n54 VTAIL.n11 171.744
R125 VTAIL.n61 VTAIL.n11 171.744
R126 VTAIL.n62 VTAIL.n61 171.744
R127 VTAIL.n62 VTAIL.n7 171.744
R128 VTAIL.n70 VTAIL.n7 171.744
R129 VTAIL.n71 VTAIL.n70 171.744
R130 VTAIL.n72 VTAIL.n71 171.744
R131 VTAIL.n72 VTAIL.n3 171.744
R132 VTAIL.n79 VTAIL.n3 171.744
R133 VTAIL.n80 VTAIL.n79 171.744
R134 VTAIL.n252 VTAIL.n251 171.744
R135 VTAIL.n251 VTAIL.n175 171.744
R136 VTAIL.n180 VTAIL.n175 171.744
R137 VTAIL.n244 VTAIL.n180 171.744
R138 VTAIL.n244 VTAIL.n243 171.744
R139 VTAIL.n243 VTAIL.n181 171.744
R140 VTAIL.n236 VTAIL.n181 171.744
R141 VTAIL.n236 VTAIL.n235 171.744
R142 VTAIL.n235 VTAIL.n185 171.744
R143 VTAIL.n228 VTAIL.n185 171.744
R144 VTAIL.n228 VTAIL.n227 171.744
R145 VTAIL.n227 VTAIL.n189 171.744
R146 VTAIL.n220 VTAIL.n189 171.744
R147 VTAIL.n220 VTAIL.n219 171.744
R148 VTAIL.n219 VTAIL.n193 171.744
R149 VTAIL.n212 VTAIL.n193 171.744
R150 VTAIL.n212 VTAIL.n211 171.744
R151 VTAIL.n211 VTAIL.n197 171.744
R152 VTAIL.n204 VTAIL.n197 171.744
R153 VTAIL.n204 VTAIL.n203 171.744
R154 VTAIL.n166 VTAIL.n165 171.744
R155 VTAIL.n165 VTAIL.n89 171.744
R156 VTAIL.n94 VTAIL.n89 171.744
R157 VTAIL.n158 VTAIL.n94 171.744
R158 VTAIL.n158 VTAIL.n157 171.744
R159 VTAIL.n157 VTAIL.n95 171.744
R160 VTAIL.n150 VTAIL.n95 171.744
R161 VTAIL.n150 VTAIL.n149 171.744
R162 VTAIL.n149 VTAIL.n99 171.744
R163 VTAIL.n142 VTAIL.n99 171.744
R164 VTAIL.n142 VTAIL.n141 171.744
R165 VTAIL.n141 VTAIL.n103 171.744
R166 VTAIL.n134 VTAIL.n103 171.744
R167 VTAIL.n134 VTAIL.n133 171.744
R168 VTAIL.n133 VTAIL.n107 171.744
R169 VTAIL.n126 VTAIL.n107 171.744
R170 VTAIL.n126 VTAIL.n125 171.744
R171 VTAIL.n125 VTAIL.n111 171.744
R172 VTAIL.n118 VTAIL.n111 171.744
R173 VTAIL.n118 VTAIL.n117 171.744
R174 VTAIL.n287 VTAIL.t3 85.8723
R175 VTAIL.n29 VTAIL.t0 85.8723
R176 VTAIL.n203 VTAIL.t1 85.8723
R177 VTAIL.n117 VTAIL.t2 85.8723
R178 VTAIL.n343 VTAIL.n342 31.7975
R179 VTAIL.n85 VTAIL.n84 31.7975
R180 VTAIL.n257 VTAIL.n256 31.7975
R181 VTAIL.n171 VTAIL.n170 31.7975
R182 VTAIL.n171 VTAIL.n85 31.3496
R183 VTAIL.n343 VTAIL.n257 28.4703
R184 VTAIL.n286 VTAIL.n285 16.3895
R185 VTAIL.n28 VTAIL.n27 16.3895
R186 VTAIL.n202 VTAIL.n201 16.3895
R187 VTAIL.n116 VTAIL.n115 16.3895
R188 VTAIL.n331 VTAIL.n262 13.1884
R189 VTAIL.n73 VTAIL.n4 13.1884
R190 VTAIL.n178 VTAIL.n176 13.1884
R191 VTAIL.n92 VTAIL.n90 13.1884
R192 VTAIL.n289 VTAIL.n284 12.8005
R193 VTAIL.n332 VTAIL.n264 12.8005
R194 VTAIL.n336 VTAIL.n335 12.8005
R195 VTAIL.n31 VTAIL.n26 12.8005
R196 VTAIL.n74 VTAIL.n6 12.8005
R197 VTAIL.n78 VTAIL.n77 12.8005
R198 VTAIL.n250 VTAIL.n249 12.8005
R199 VTAIL.n246 VTAIL.n245 12.8005
R200 VTAIL.n205 VTAIL.n200 12.8005
R201 VTAIL.n164 VTAIL.n163 12.8005
R202 VTAIL.n160 VTAIL.n159 12.8005
R203 VTAIL.n119 VTAIL.n114 12.8005
R204 VTAIL.n290 VTAIL.n282 12.0247
R205 VTAIL.n327 VTAIL.n326 12.0247
R206 VTAIL.n339 VTAIL.n260 12.0247
R207 VTAIL.n32 VTAIL.n24 12.0247
R208 VTAIL.n69 VTAIL.n68 12.0247
R209 VTAIL.n81 VTAIL.n2 12.0247
R210 VTAIL.n253 VTAIL.n174 12.0247
R211 VTAIL.n242 VTAIL.n179 12.0247
R212 VTAIL.n206 VTAIL.n198 12.0247
R213 VTAIL.n167 VTAIL.n88 12.0247
R214 VTAIL.n156 VTAIL.n93 12.0247
R215 VTAIL.n120 VTAIL.n112 12.0247
R216 VTAIL.n294 VTAIL.n293 11.249
R217 VTAIL.n325 VTAIL.n266 11.249
R218 VTAIL.n340 VTAIL.n258 11.249
R219 VTAIL.n36 VTAIL.n35 11.249
R220 VTAIL.n67 VTAIL.n8 11.249
R221 VTAIL.n82 VTAIL.n0 11.249
R222 VTAIL.n254 VTAIL.n172 11.249
R223 VTAIL.n241 VTAIL.n182 11.249
R224 VTAIL.n210 VTAIL.n209 11.249
R225 VTAIL.n168 VTAIL.n86 11.249
R226 VTAIL.n155 VTAIL.n96 11.249
R227 VTAIL.n124 VTAIL.n123 11.249
R228 VTAIL.n297 VTAIL.n280 10.4732
R229 VTAIL.n322 VTAIL.n321 10.4732
R230 VTAIL.n39 VTAIL.n22 10.4732
R231 VTAIL.n64 VTAIL.n63 10.4732
R232 VTAIL.n238 VTAIL.n237 10.4732
R233 VTAIL.n213 VTAIL.n196 10.4732
R234 VTAIL.n152 VTAIL.n151 10.4732
R235 VTAIL.n127 VTAIL.n110 10.4732
R236 VTAIL.n298 VTAIL.n278 9.69747
R237 VTAIL.n318 VTAIL.n268 9.69747
R238 VTAIL.n40 VTAIL.n20 9.69747
R239 VTAIL.n60 VTAIL.n10 9.69747
R240 VTAIL.n234 VTAIL.n184 9.69747
R241 VTAIL.n214 VTAIL.n194 9.69747
R242 VTAIL.n148 VTAIL.n98 9.69747
R243 VTAIL.n128 VTAIL.n108 9.69747
R244 VTAIL.n342 VTAIL.n341 9.45567
R245 VTAIL.n84 VTAIL.n83 9.45567
R246 VTAIL.n256 VTAIL.n255 9.45567
R247 VTAIL.n170 VTAIL.n169 9.45567
R248 VTAIL.n341 VTAIL.n340 9.3005
R249 VTAIL.n260 VTAIL.n259 9.3005
R250 VTAIL.n335 VTAIL.n334 9.3005
R251 VTAIL.n307 VTAIL.n306 9.3005
R252 VTAIL.n276 VTAIL.n275 9.3005
R253 VTAIL.n301 VTAIL.n300 9.3005
R254 VTAIL.n299 VTAIL.n298 9.3005
R255 VTAIL.n280 VTAIL.n279 9.3005
R256 VTAIL.n293 VTAIL.n292 9.3005
R257 VTAIL.n291 VTAIL.n290 9.3005
R258 VTAIL.n284 VTAIL.n283 9.3005
R259 VTAIL.n309 VTAIL.n308 9.3005
R260 VTAIL.n272 VTAIL.n271 9.3005
R261 VTAIL.n315 VTAIL.n314 9.3005
R262 VTAIL.n317 VTAIL.n316 9.3005
R263 VTAIL.n268 VTAIL.n267 9.3005
R264 VTAIL.n323 VTAIL.n322 9.3005
R265 VTAIL.n325 VTAIL.n324 9.3005
R266 VTAIL.n326 VTAIL.n263 9.3005
R267 VTAIL.n333 VTAIL.n332 9.3005
R268 VTAIL.n83 VTAIL.n82 9.3005
R269 VTAIL.n2 VTAIL.n1 9.3005
R270 VTAIL.n77 VTAIL.n76 9.3005
R271 VTAIL.n49 VTAIL.n48 9.3005
R272 VTAIL.n18 VTAIL.n17 9.3005
R273 VTAIL.n43 VTAIL.n42 9.3005
R274 VTAIL.n41 VTAIL.n40 9.3005
R275 VTAIL.n22 VTAIL.n21 9.3005
R276 VTAIL.n35 VTAIL.n34 9.3005
R277 VTAIL.n33 VTAIL.n32 9.3005
R278 VTAIL.n26 VTAIL.n25 9.3005
R279 VTAIL.n51 VTAIL.n50 9.3005
R280 VTAIL.n14 VTAIL.n13 9.3005
R281 VTAIL.n57 VTAIL.n56 9.3005
R282 VTAIL.n59 VTAIL.n58 9.3005
R283 VTAIL.n10 VTAIL.n9 9.3005
R284 VTAIL.n65 VTAIL.n64 9.3005
R285 VTAIL.n67 VTAIL.n66 9.3005
R286 VTAIL.n68 VTAIL.n5 9.3005
R287 VTAIL.n75 VTAIL.n74 9.3005
R288 VTAIL.n188 VTAIL.n187 9.3005
R289 VTAIL.n231 VTAIL.n230 9.3005
R290 VTAIL.n233 VTAIL.n232 9.3005
R291 VTAIL.n184 VTAIL.n183 9.3005
R292 VTAIL.n239 VTAIL.n238 9.3005
R293 VTAIL.n241 VTAIL.n240 9.3005
R294 VTAIL.n179 VTAIL.n177 9.3005
R295 VTAIL.n247 VTAIL.n246 9.3005
R296 VTAIL.n255 VTAIL.n254 9.3005
R297 VTAIL.n174 VTAIL.n173 9.3005
R298 VTAIL.n249 VTAIL.n248 9.3005
R299 VTAIL.n225 VTAIL.n224 9.3005
R300 VTAIL.n223 VTAIL.n222 9.3005
R301 VTAIL.n192 VTAIL.n191 9.3005
R302 VTAIL.n217 VTAIL.n216 9.3005
R303 VTAIL.n215 VTAIL.n214 9.3005
R304 VTAIL.n196 VTAIL.n195 9.3005
R305 VTAIL.n209 VTAIL.n208 9.3005
R306 VTAIL.n207 VTAIL.n206 9.3005
R307 VTAIL.n200 VTAIL.n199 9.3005
R308 VTAIL.n102 VTAIL.n101 9.3005
R309 VTAIL.n145 VTAIL.n144 9.3005
R310 VTAIL.n147 VTAIL.n146 9.3005
R311 VTAIL.n98 VTAIL.n97 9.3005
R312 VTAIL.n153 VTAIL.n152 9.3005
R313 VTAIL.n155 VTAIL.n154 9.3005
R314 VTAIL.n93 VTAIL.n91 9.3005
R315 VTAIL.n161 VTAIL.n160 9.3005
R316 VTAIL.n169 VTAIL.n168 9.3005
R317 VTAIL.n88 VTAIL.n87 9.3005
R318 VTAIL.n163 VTAIL.n162 9.3005
R319 VTAIL.n139 VTAIL.n138 9.3005
R320 VTAIL.n137 VTAIL.n136 9.3005
R321 VTAIL.n106 VTAIL.n105 9.3005
R322 VTAIL.n131 VTAIL.n130 9.3005
R323 VTAIL.n129 VTAIL.n128 9.3005
R324 VTAIL.n110 VTAIL.n109 9.3005
R325 VTAIL.n123 VTAIL.n122 9.3005
R326 VTAIL.n121 VTAIL.n120 9.3005
R327 VTAIL.n114 VTAIL.n113 9.3005
R328 VTAIL.n302 VTAIL.n301 8.92171
R329 VTAIL.n317 VTAIL.n270 8.92171
R330 VTAIL.n44 VTAIL.n43 8.92171
R331 VTAIL.n59 VTAIL.n12 8.92171
R332 VTAIL.n233 VTAIL.n186 8.92171
R333 VTAIL.n218 VTAIL.n217 8.92171
R334 VTAIL.n147 VTAIL.n100 8.92171
R335 VTAIL.n132 VTAIL.n131 8.92171
R336 VTAIL.n305 VTAIL.n276 8.14595
R337 VTAIL.n314 VTAIL.n313 8.14595
R338 VTAIL.n47 VTAIL.n18 8.14595
R339 VTAIL.n56 VTAIL.n55 8.14595
R340 VTAIL.n230 VTAIL.n229 8.14595
R341 VTAIL.n221 VTAIL.n192 8.14595
R342 VTAIL.n144 VTAIL.n143 8.14595
R343 VTAIL.n135 VTAIL.n106 8.14595
R344 VTAIL.n306 VTAIL.n274 7.3702
R345 VTAIL.n310 VTAIL.n272 7.3702
R346 VTAIL.n48 VTAIL.n16 7.3702
R347 VTAIL.n52 VTAIL.n14 7.3702
R348 VTAIL.n226 VTAIL.n188 7.3702
R349 VTAIL.n222 VTAIL.n190 7.3702
R350 VTAIL.n140 VTAIL.n102 7.3702
R351 VTAIL.n136 VTAIL.n104 7.3702
R352 VTAIL.n309 VTAIL.n274 6.59444
R353 VTAIL.n310 VTAIL.n309 6.59444
R354 VTAIL.n51 VTAIL.n16 6.59444
R355 VTAIL.n52 VTAIL.n51 6.59444
R356 VTAIL.n226 VTAIL.n225 6.59444
R357 VTAIL.n225 VTAIL.n190 6.59444
R358 VTAIL.n140 VTAIL.n139 6.59444
R359 VTAIL.n139 VTAIL.n104 6.59444
R360 VTAIL.n306 VTAIL.n305 5.81868
R361 VTAIL.n313 VTAIL.n272 5.81868
R362 VTAIL.n48 VTAIL.n47 5.81868
R363 VTAIL.n55 VTAIL.n14 5.81868
R364 VTAIL.n229 VTAIL.n188 5.81868
R365 VTAIL.n222 VTAIL.n221 5.81868
R366 VTAIL.n143 VTAIL.n102 5.81868
R367 VTAIL.n136 VTAIL.n135 5.81868
R368 VTAIL.n302 VTAIL.n276 5.04292
R369 VTAIL.n314 VTAIL.n270 5.04292
R370 VTAIL.n44 VTAIL.n18 5.04292
R371 VTAIL.n56 VTAIL.n12 5.04292
R372 VTAIL.n230 VTAIL.n186 5.04292
R373 VTAIL.n218 VTAIL.n192 5.04292
R374 VTAIL.n144 VTAIL.n100 5.04292
R375 VTAIL.n132 VTAIL.n106 5.04292
R376 VTAIL.n301 VTAIL.n278 4.26717
R377 VTAIL.n318 VTAIL.n317 4.26717
R378 VTAIL.n43 VTAIL.n20 4.26717
R379 VTAIL.n60 VTAIL.n59 4.26717
R380 VTAIL.n234 VTAIL.n233 4.26717
R381 VTAIL.n217 VTAIL.n194 4.26717
R382 VTAIL.n148 VTAIL.n147 4.26717
R383 VTAIL.n131 VTAIL.n108 4.26717
R384 VTAIL.n285 VTAIL.n283 3.70982
R385 VTAIL.n27 VTAIL.n25 3.70982
R386 VTAIL.n201 VTAIL.n199 3.70982
R387 VTAIL.n115 VTAIL.n113 3.70982
R388 VTAIL.n298 VTAIL.n297 3.49141
R389 VTAIL.n321 VTAIL.n268 3.49141
R390 VTAIL.n40 VTAIL.n39 3.49141
R391 VTAIL.n63 VTAIL.n10 3.49141
R392 VTAIL.n237 VTAIL.n184 3.49141
R393 VTAIL.n214 VTAIL.n213 3.49141
R394 VTAIL.n151 VTAIL.n98 3.49141
R395 VTAIL.n128 VTAIL.n127 3.49141
R396 VTAIL.n294 VTAIL.n280 2.71565
R397 VTAIL.n322 VTAIL.n266 2.71565
R398 VTAIL.n342 VTAIL.n258 2.71565
R399 VTAIL.n36 VTAIL.n22 2.71565
R400 VTAIL.n64 VTAIL.n8 2.71565
R401 VTAIL.n84 VTAIL.n0 2.71565
R402 VTAIL.n256 VTAIL.n172 2.71565
R403 VTAIL.n238 VTAIL.n182 2.71565
R404 VTAIL.n210 VTAIL.n196 2.71565
R405 VTAIL.n170 VTAIL.n86 2.71565
R406 VTAIL.n152 VTAIL.n96 2.71565
R407 VTAIL.n124 VTAIL.n110 2.71565
R408 VTAIL.n293 VTAIL.n282 1.93989
R409 VTAIL.n327 VTAIL.n325 1.93989
R410 VTAIL.n340 VTAIL.n339 1.93989
R411 VTAIL.n35 VTAIL.n24 1.93989
R412 VTAIL.n69 VTAIL.n67 1.93989
R413 VTAIL.n82 VTAIL.n81 1.93989
R414 VTAIL.n254 VTAIL.n253 1.93989
R415 VTAIL.n242 VTAIL.n241 1.93989
R416 VTAIL.n209 VTAIL.n198 1.93989
R417 VTAIL.n168 VTAIL.n167 1.93989
R418 VTAIL.n156 VTAIL.n155 1.93989
R419 VTAIL.n123 VTAIL.n112 1.93989
R420 VTAIL.n257 VTAIL.n171 1.90998
R421 VTAIL VTAIL.n85 1.24834
R422 VTAIL.n290 VTAIL.n289 1.16414
R423 VTAIL.n326 VTAIL.n264 1.16414
R424 VTAIL.n336 VTAIL.n260 1.16414
R425 VTAIL.n32 VTAIL.n31 1.16414
R426 VTAIL.n68 VTAIL.n6 1.16414
R427 VTAIL.n78 VTAIL.n2 1.16414
R428 VTAIL.n250 VTAIL.n174 1.16414
R429 VTAIL.n245 VTAIL.n179 1.16414
R430 VTAIL.n206 VTAIL.n205 1.16414
R431 VTAIL.n164 VTAIL.n88 1.16414
R432 VTAIL.n159 VTAIL.n93 1.16414
R433 VTAIL.n120 VTAIL.n119 1.16414
R434 VTAIL VTAIL.n343 0.662138
R435 VTAIL.n286 VTAIL.n284 0.388379
R436 VTAIL.n332 VTAIL.n331 0.388379
R437 VTAIL.n335 VTAIL.n262 0.388379
R438 VTAIL.n28 VTAIL.n26 0.388379
R439 VTAIL.n74 VTAIL.n73 0.388379
R440 VTAIL.n77 VTAIL.n4 0.388379
R441 VTAIL.n249 VTAIL.n176 0.388379
R442 VTAIL.n246 VTAIL.n178 0.388379
R443 VTAIL.n202 VTAIL.n200 0.388379
R444 VTAIL.n163 VTAIL.n90 0.388379
R445 VTAIL.n160 VTAIL.n92 0.388379
R446 VTAIL.n116 VTAIL.n114 0.388379
R447 VTAIL.n291 VTAIL.n283 0.155672
R448 VTAIL.n292 VTAIL.n291 0.155672
R449 VTAIL.n292 VTAIL.n279 0.155672
R450 VTAIL.n299 VTAIL.n279 0.155672
R451 VTAIL.n300 VTAIL.n299 0.155672
R452 VTAIL.n300 VTAIL.n275 0.155672
R453 VTAIL.n307 VTAIL.n275 0.155672
R454 VTAIL.n308 VTAIL.n307 0.155672
R455 VTAIL.n308 VTAIL.n271 0.155672
R456 VTAIL.n315 VTAIL.n271 0.155672
R457 VTAIL.n316 VTAIL.n315 0.155672
R458 VTAIL.n316 VTAIL.n267 0.155672
R459 VTAIL.n323 VTAIL.n267 0.155672
R460 VTAIL.n324 VTAIL.n323 0.155672
R461 VTAIL.n324 VTAIL.n263 0.155672
R462 VTAIL.n333 VTAIL.n263 0.155672
R463 VTAIL.n334 VTAIL.n333 0.155672
R464 VTAIL.n334 VTAIL.n259 0.155672
R465 VTAIL.n341 VTAIL.n259 0.155672
R466 VTAIL.n33 VTAIL.n25 0.155672
R467 VTAIL.n34 VTAIL.n33 0.155672
R468 VTAIL.n34 VTAIL.n21 0.155672
R469 VTAIL.n41 VTAIL.n21 0.155672
R470 VTAIL.n42 VTAIL.n41 0.155672
R471 VTAIL.n42 VTAIL.n17 0.155672
R472 VTAIL.n49 VTAIL.n17 0.155672
R473 VTAIL.n50 VTAIL.n49 0.155672
R474 VTAIL.n50 VTAIL.n13 0.155672
R475 VTAIL.n57 VTAIL.n13 0.155672
R476 VTAIL.n58 VTAIL.n57 0.155672
R477 VTAIL.n58 VTAIL.n9 0.155672
R478 VTAIL.n65 VTAIL.n9 0.155672
R479 VTAIL.n66 VTAIL.n65 0.155672
R480 VTAIL.n66 VTAIL.n5 0.155672
R481 VTAIL.n75 VTAIL.n5 0.155672
R482 VTAIL.n76 VTAIL.n75 0.155672
R483 VTAIL.n76 VTAIL.n1 0.155672
R484 VTAIL.n83 VTAIL.n1 0.155672
R485 VTAIL.n255 VTAIL.n173 0.155672
R486 VTAIL.n248 VTAIL.n173 0.155672
R487 VTAIL.n248 VTAIL.n247 0.155672
R488 VTAIL.n247 VTAIL.n177 0.155672
R489 VTAIL.n240 VTAIL.n177 0.155672
R490 VTAIL.n240 VTAIL.n239 0.155672
R491 VTAIL.n239 VTAIL.n183 0.155672
R492 VTAIL.n232 VTAIL.n183 0.155672
R493 VTAIL.n232 VTAIL.n231 0.155672
R494 VTAIL.n231 VTAIL.n187 0.155672
R495 VTAIL.n224 VTAIL.n187 0.155672
R496 VTAIL.n224 VTAIL.n223 0.155672
R497 VTAIL.n223 VTAIL.n191 0.155672
R498 VTAIL.n216 VTAIL.n191 0.155672
R499 VTAIL.n216 VTAIL.n215 0.155672
R500 VTAIL.n215 VTAIL.n195 0.155672
R501 VTAIL.n208 VTAIL.n195 0.155672
R502 VTAIL.n208 VTAIL.n207 0.155672
R503 VTAIL.n207 VTAIL.n199 0.155672
R504 VTAIL.n169 VTAIL.n87 0.155672
R505 VTAIL.n162 VTAIL.n87 0.155672
R506 VTAIL.n162 VTAIL.n161 0.155672
R507 VTAIL.n161 VTAIL.n91 0.155672
R508 VTAIL.n154 VTAIL.n91 0.155672
R509 VTAIL.n154 VTAIL.n153 0.155672
R510 VTAIL.n153 VTAIL.n97 0.155672
R511 VTAIL.n146 VTAIL.n97 0.155672
R512 VTAIL.n146 VTAIL.n145 0.155672
R513 VTAIL.n145 VTAIL.n101 0.155672
R514 VTAIL.n138 VTAIL.n101 0.155672
R515 VTAIL.n138 VTAIL.n137 0.155672
R516 VTAIL.n137 VTAIL.n105 0.155672
R517 VTAIL.n130 VTAIL.n105 0.155672
R518 VTAIL.n130 VTAIL.n129 0.155672
R519 VTAIL.n129 VTAIL.n109 0.155672
R520 VTAIL.n122 VTAIL.n109 0.155672
R521 VTAIL.n122 VTAIL.n121 0.155672
R522 VTAIL.n121 VTAIL.n113 0.155672
R523 VDD2.n165 VDD2.n85 756.745
R524 VDD2.n80 VDD2.n0 756.745
R525 VDD2.n166 VDD2.n165 585
R526 VDD2.n164 VDD2.n163 585
R527 VDD2.n89 VDD2.n88 585
R528 VDD2.n93 VDD2.n91 585
R529 VDD2.n158 VDD2.n157 585
R530 VDD2.n156 VDD2.n155 585
R531 VDD2.n95 VDD2.n94 585
R532 VDD2.n150 VDD2.n149 585
R533 VDD2.n148 VDD2.n147 585
R534 VDD2.n99 VDD2.n98 585
R535 VDD2.n142 VDD2.n141 585
R536 VDD2.n140 VDD2.n139 585
R537 VDD2.n103 VDD2.n102 585
R538 VDD2.n134 VDD2.n133 585
R539 VDD2.n132 VDD2.n131 585
R540 VDD2.n107 VDD2.n106 585
R541 VDD2.n126 VDD2.n125 585
R542 VDD2.n124 VDD2.n123 585
R543 VDD2.n111 VDD2.n110 585
R544 VDD2.n118 VDD2.n117 585
R545 VDD2.n116 VDD2.n115 585
R546 VDD2.n29 VDD2.n28 585
R547 VDD2.n31 VDD2.n30 585
R548 VDD2.n24 VDD2.n23 585
R549 VDD2.n37 VDD2.n36 585
R550 VDD2.n39 VDD2.n38 585
R551 VDD2.n20 VDD2.n19 585
R552 VDD2.n45 VDD2.n44 585
R553 VDD2.n47 VDD2.n46 585
R554 VDD2.n16 VDD2.n15 585
R555 VDD2.n53 VDD2.n52 585
R556 VDD2.n55 VDD2.n54 585
R557 VDD2.n12 VDD2.n11 585
R558 VDD2.n61 VDD2.n60 585
R559 VDD2.n63 VDD2.n62 585
R560 VDD2.n8 VDD2.n7 585
R561 VDD2.n70 VDD2.n69 585
R562 VDD2.n71 VDD2.n6 585
R563 VDD2.n73 VDD2.n72 585
R564 VDD2.n4 VDD2.n3 585
R565 VDD2.n79 VDD2.n78 585
R566 VDD2.n81 VDD2.n80 585
R567 VDD2.n114 VDD2.t1 327.466
R568 VDD2.n27 VDD2.t0 327.466
R569 VDD2.n165 VDD2.n164 171.744
R570 VDD2.n164 VDD2.n88 171.744
R571 VDD2.n93 VDD2.n88 171.744
R572 VDD2.n157 VDD2.n93 171.744
R573 VDD2.n157 VDD2.n156 171.744
R574 VDD2.n156 VDD2.n94 171.744
R575 VDD2.n149 VDD2.n94 171.744
R576 VDD2.n149 VDD2.n148 171.744
R577 VDD2.n148 VDD2.n98 171.744
R578 VDD2.n141 VDD2.n98 171.744
R579 VDD2.n141 VDD2.n140 171.744
R580 VDD2.n140 VDD2.n102 171.744
R581 VDD2.n133 VDD2.n102 171.744
R582 VDD2.n133 VDD2.n132 171.744
R583 VDD2.n132 VDD2.n106 171.744
R584 VDD2.n125 VDD2.n106 171.744
R585 VDD2.n125 VDD2.n124 171.744
R586 VDD2.n124 VDD2.n110 171.744
R587 VDD2.n117 VDD2.n110 171.744
R588 VDD2.n117 VDD2.n116 171.744
R589 VDD2.n30 VDD2.n29 171.744
R590 VDD2.n30 VDD2.n23 171.744
R591 VDD2.n37 VDD2.n23 171.744
R592 VDD2.n38 VDD2.n37 171.744
R593 VDD2.n38 VDD2.n19 171.744
R594 VDD2.n45 VDD2.n19 171.744
R595 VDD2.n46 VDD2.n45 171.744
R596 VDD2.n46 VDD2.n15 171.744
R597 VDD2.n53 VDD2.n15 171.744
R598 VDD2.n54 VDD2.n53 171.744
R599 VDD2.n54 VDD2.n11 171.744
R600 VDD2.n61 VDD2.n11 171.744
R601 VDD2.n62 VDD2.n61 171.744
R602 VDD2.n62 VDD2.n7 171.744
R603 VDD2.n70 VDD2.n7 171.744
R604 VDD2.n71 VDD2.n70 171.744
R605 VDD2.n72 VDD2.n71 171.744
R606 VDD2.n72 VDD2.n3 171.744
R607 VDD2.n79 VDD2.n3 171.744
R608 VDD2.n80 VDD2.n79 171.744
R609 VDD2.n170 VDD2.n84 91.1185
R610 VDD2.n116 VDD2.t1 85.8723
R611 VDD2.n29 VDD2.t0 85.8723
R612 VDD2.n170 VDD2.n169 48.4763
R613 VDD2.n115 VDD2.n114 16.3895
R614 VDD2.n28 VDD2.n27 16.3895
R615 VDD2.n91 VDD2.n89 13.1884
R616 VDD2.n73 VDD2.n4 13.1884
R617 VDD2.n163 VDD2.n162 12.8005
R618 VDD2.n159 VDD2.n158 12.8005
R619 VDD2.n118 VDD2.n113 12.8005
R620 VDD2.n31 VDD2.n26 12.8005
R621 VDD2.n74 VDD2.n6 12.8005
R622 VDD2.n78 VDD2.n77 12.8005
R623 VDD2.n166 VDD2.n87 12.0247
R624 VDD2.n155 VDD2.n92 12.0247
R625 VDD2.n119 VDD2.n111 12.0247
R626 VDD2.n32 VDD2.n24 12.0247
R627 VDD2.n69 VDD2.n68 12.0247
R628 VDD2.n81 VDD2.n2 12.0247
R629 VDD2.n167 VDD2.n85 11.249
R630 VDD2.n154 VDD2.n95 11.249
R631 VDD2.n123 VDD2.n122 11.249
R632 VDD2.n36 VDD2.n35 11.249
R633 VDD2.n67 VDD2.n8 11.249
R634 VDD2.n82 VDD2.n0 11.249
R635 VDD2.n151 VDD2.n150 10.4732
R636 VDD2.n126 VDD2.n109 10.4732
R637 VDD2.n39 VDD2.n22 10.4732
R638 VDD2.n64 VDD2.n63 10.4732
R639 VDD2.n147 VDD2.n97 9.69747
R640 VDD2.n127 VDD2.n107 9.69747
R641 VDD2.n40 VDD2.n20 9.69747
R642 VDD2.n60 VDD2.n10 9.69747
R643 VDD2.n169 VDD2.n168 9.45567
R644 VDD2.n84 VDD2.n83 9.45567
R645 VDD2.n101 VDD2.n100 9.3005
R646 VDD2.n144 VDD2.n143 9.3005
R647 VDD2.n146 VDD2.n145 9.3005
R648 VDD2.n97 VDD2.n96 9.3005
R649 VDD2.n152 VDD2.n151 9.3005
R650 VDD2.n154 VDD2.n153 9.3005
R651 VDD2.n92 VDD2.n90 9.3005
R652 VDD2.n160 VDD2.n159 9.3005
R653 VDD2.n168 VDD2.n167 9.3005
R654 VDD2.n87 VDD2.n86 9.3005
R655 VDD2.n162 VDD2.n161 9.3005
R656 VDD2.n138 VDD2.n137 9.3005
R657 VDD2.n136 VDD2.n135 9.3005
R658 VDD2.n105 VDD2.n104 9.3005
R659 VDD2.n130 VDD2.n129 9.3005
R660 VDD2.n128 VDD2.n127 9.3005
R661 VDD2.n109 VDD2.n108 9.3005
R662 VDD2.n122 VDD2.n121 9.3005
R663 VDD2.n120 VDD2.n119 9.3005
R664 VDD2.n113 VDD2.n112 9.3005
R665 VDD2.n83 VDD2.n82 9.3005
R666 VDD2.n2 VDD2.n1 9.3005
R667 VDD2.n77 VDD2.n76 9.3005
R668 VDD2.n49 VDD2.n48 9.3005
R669 VDD2.n18 VDD2.n17 9.3005
R670 VDD2.n43 VDD2.n42 9.3005
R671 VDD2.n41 VDD2.n40 9.3005
R672 VDD2.n22 VDD2.n21 9.3005
R673 VDD2.n35 VDD2.n34 9.3005
R674 VDD2.n33 VDD2.n32 9.3005
R675 VDD2.n26 VDD2.n25 9.3005
R676 VDD2.n51 VDD2.n50 9.3005
R677 VDD2.n14 VDD2.n13 9.3005
R678 VDD2.n57 VDD2.n56 9.3005
R679 VDD2.n59 VDD2.n58 9.3005
R680 VDD2.n10 VDD2.n9 9.3005
R681 VDD2.n65 VDD2.n64 9.3005
R682 VDD2.n67 VDD2.n66 9.3005
R683 VDD2.n68 VDD2.n5 9.3005
R684 VDD2.n75 VDD2.n74 9.3005
R685 VDD2.n146 VDD2.n99 8.92171
R686 VDD2.n131 VDD2.n130 8.92171
R687 VDD2.n44 VDD2.n43 8.92171
R688 VDD2.n59 VDD2.n12 8.92171
R689 VDD2.n143 VDD2.n142 8.14595
R690 VDD2.n134 VDD2.n105 8.14595
R691 VDD2.n47 VDD2.n18 8.14595
R692 VDD2.n56 VDD2.n55 8.14595
R693 VDD2.n139 VDD2.n101 7.3702
R694 VDD2.n135 VDD2.n103 7.3702
R695 VDD2.n48 VDD2.n16 7.3702
R696 VDD2.n52 VDD2.n14 7.3702
R697 VDD2.n139 VDD2.n138 6.59444
R698 VDD2.n138 VDD2.n103 6.59444
R699 VDD2.n51 VDD2.n16 6.59444
R700 VDD2.n52 VDD2.n51 6.59444
R701 VDD2.n142 VDD2.n101 5.81868
R702 VDD2.n135 VDD2.n134 5.81868
R703 VDD2.n48 VDD2.n47 5.81868
R704 VDD2.n55 VDD2.n14 5.81868
R705 VDD2.n143 VDD2.n99 5.04292
R706 VDD2.n131 VDD2.n105 5.04292
R707 VDD2.n44 VDD2.n18 5.04292
R708 VDD2.n56 VDD2.n12 5.04292
R709 VDD2.n147 VDD2.n146 4.26717
R710 VDD2.n130 VDD2.n107 4.26717
R711 VDD2.n43 VDD2.n20 4.26717
R712 VDD2.n60 VDD2.n59 4.26717
R713 VDD2.n114 VDD2.n112 3.70982
R714 VDD2.n27 VDD2.n25 3.70982
R715 VDD2.n150 VDD2.n97 3.49141
R716 VDD2.n127 VDD2.n126 3.49141
R717 VDD2.n40 VDD2.n39 3.49141
R718 VDD2.n63 VDD2.n10 3.49141
R719 VDD2.n169 VDD2.n85 2.71565
R720 VDD2.n151 VDD2.n95 2.71565
R721 VDD2.n123 VDD2.n109 2.71565
R722 VDD2.n36 VDD2.n22 2.71565
R723 VDD2.n64 VDD2.n8 2.71565
R724 VDD2.n84 VDD2.n0 2.71565
R725 VDD2.n167 VDD2.n166 1.93989
R726 VDD2.n155 VDD2.n154 1.93989
R727 VDD2.n122 VDD2.n111 1.93989
R728 VDD2.n35 VDD2.n24 1.93989
R729 VDD2.n69 VDD2.n67 1.93989
R730 VDD2.n82 VDD2.n81 1.93989
R731 VDD2.n163 VDD2.n87 1.16414
R732 VDD2.n158 VDD2.n92 1.16414
R733 VDD2.n119 VDD2.n118 1.16414
R734 VDD2.n32 VDD2.n31 1.16414
R735 VDD2.n68 VDD2.n6 1.16414
R736 VDD2.n78 VDD2.n2 1.16414
R737 VDD2 VDD2.n170 0.778517
R738 VDD2.n162 VDD2.n89 0.388379
R739 VDD2.n159 VDD2.n91 0.388379
R740 VDD2.n115 VDD2.n113 0.388379
R741 VDD2.n28 VDD2.n26 0.388379
R742 VDD2.n74 VDD2.n73 0.388379
R743 VDD2.n77 VDD2.n4 0.388379
R744 VDD2.n168 VDD2.n86 0.155672
R745 VDD2.n161 VDD2.n86 0.155672
R746 VDD2.n161 VDD2.n160 0.155672
R747 VDD2.n160 VDD2.n90 0.155672
R748 VDD2.n153 VDD2.n90 0.155672
R749 VDD2.n153 VDD2.n152 0.155672
R750 VDD2.n152 VDD2.n96 0.155672
R751 VDD2.n145 VDD2.n96 0.155672
R752 VDD2.n145 VDD2.n144 0.155672
R753 VDD2.n144 VDD2.n100 0.155672
R754 VDD2.n137 VDD2.n100 0.155672
R755 VDD2.n137 VDD2.n136 0.155672
R756 VDD2.n136 VDD2.n104 0.155672
R757 VDD2.n129 VDD2.n104 0.155672
R758 VDD2.n129 VDD2.n128 0.155672
R759 VDD2.n128 VDD2.n108 0.155672
R760 VDD2.n121 VDD2.n108 0.155672
R761 VDD2.n121 VDD2.n120 0.155672
R762 VDD2.n120 VDD2.n112 0.155672
R763 VDD2.n33 VDD2.n25 0.155672
R764 VDD2.n34 VDD2.n33 0.155672
R765 VDD2.n34 VDD2.n21 0.155672
R766 VDD2.n41 VDD2.n21 0.155672
R767 VDD2.n42 VDD2.n41 0.155672
R768 VDD2.n42 VDD2.n17 0.155672
R769 VDD2.n49 VDD2.n17 0.155672
R770 VDD2.n50 VDD2.n49 0.155672
R771 VDD2.n50 VDD2.n13 0.155672
R772 VDD2.n57 VDD2.n13 0.155672
R773 VDD2.n58 VDD2.n57 0.155672
R774 VDD2.n58 VDD2.n9 0.155672
R775 VDD2.n65 VDD2.n9 0.155672
R776 VDD2.n66 VDD2.n65 0.155672
R777 VDD2.n66 VDD2.n5 0.155672
R778 VDD2.n75 VDD2.n5 0.155672
R779 VDD2.n76 VDD2.n75 0.155672
R780 VDD2.n76 VDD2.n1 0.155672
R781 VDD2.n83 VDD2.n1 0.155672
R782 B.n385 B.n104 585
R783 B.n384 B.n383 585
R784 B.n382 B.n105 585
R785 B.n381 B.n380 585
R786 B.n379 B.n106 585
R787 B.n378 B.n377 585
R788 B.n376 B.n107 585
R789 B.n375 B.n374 585
R790 B.n373 B.n108 585
R791 B.n372 B.n371 585
R792 B.n370 B.n109 585
R793 B.n369 B.n368 585
R794 B.n367 B.n110 585
R795 B.n366 B.n365 585
R796 B.n364 B.n111 585
R797 B.n363 B.n362 585
R798 B.n361 B.n112 585
R799 B.n360 B.n359 585
R800 B.n358 B.n113 585
R801 B.n357 B.n356 585
R802 B.n355 B.n114 585
R803 B.n354 B.n353 585
R804 B.n352 B.n115 585
R805 B.n351 B.n350 585
R806 B.n349 B.n116 585
R807 B.n348 B.n347 585
R808 B.n346 B.n117 585
R809 B.n345 B.n344 585
R810 B.n343 B.n118 585
R811 B.n342 B.n341 585
R812 B.n340 B.n119 585
R813 B.n339 B.n338 585
R814 B.n337 B.n120 585
R815 B.n336 B.n335 585
R816 B.n334 B.n121 585
R817 B.n333 B.n332 585
R818 B.n331 B.n122 585
R819 B.n330 B.n329 585
R820 B.n328 B.n123 585
R821 B.n327 B.n326 585
R822 B.n325 B.n124 585
R823 B.n324 B.n323 585
R824 B.n322 B.n125 585
R825 B.n321 B.n320 585
R826 B.n319 B.n126 585
R827 B.n318 B.n317 585
R828 B.n316 B.n127 585
R829 B.n315 B.n314 585
R830 B.n313 B.n128 585
R831 B.n312 B.n311 585
R832 B.n310 B.n129 585
R833 B.n308 B.n307 585
R834 B.n306 B.n132 585
R835 B.n305 B.n304 585
R836 B.n303 B.n133 585
R837 B.n302 B.n301 585
R838 B.n300 B.n134 585
R839 B.n299 B.n298 585
R840 B.n297 B.n135 585
R841 B.n296 B.n295 585
R842 B.n294 B.n136 585
R843 B.n293 B.n292 585
R844 B.n288 B.n137 585
R845 B.n287 B.n286 585
R846 B.n285 B.n138 585
R847 B.n284 B.n283 585
R848 B.n282 B.n139 585
R849 B.n281 B.n280 585
R850 B.n279 B.n140 585
R851 B.n278 B.n277 585
R852 B.n276 B.n141 585
R853 B.n275 B.n274 585
R854 B.n273 B.n142 585
R855 B.n272 B.n271 585
R856 B.n270 B.n143 585
R857 B.n269 B.n268 585
R858 B.n267 B.n144 585
R859 B.n266 B.n265 585
R860 B.n264 B.n145 585
R861 B.n263 B.n262 585
R862 B.n261 B.n146 585
R863 B.n260 B.n259 585
R864 B.n258 B.n147 585
R865 B.n257 B.n256 585
R866 B.n255 B.n148 585
R867 B.n254 B.n253 585
R868 B.n252 B.n149 585
R869 B.n251 B.n250 585
R870 B.n249 B.n150 585
R871 B.n248 B.n247 585
R872 B.n246 B.n151 585
R873 B.n245 B.n244 585
R874 B.n243 B.n152 585
R875 B.n242 B.n241 585
R876 B.n240 B.n153 585
R877 B.n239 B.n238 585
R878 B.n237 B.n154 585
R879 B.n236 B.n235 585
R880 B.n234 B.n155 585
R881 B.n233 B.n232 585
R882 B.n231 B.n156 585
R883 B.n230 B.n229 585
R884 B.n228 B.n157 585
R885 B.n227 B.n226 585
R886 B.n225 B.n158 585
R887 B.n224 B.n223 585
R888 B.n222 B.n159 585
R889 B.n221 B.n220 585
R890 B.n219 B.n160 585
R891 B.n218 B.n217 585
R892 B.n216 B.n161 585
R893 B.n215 B.n214 585
R894 B.n387 B.n386 585
R895 B.n388 B.n103 585
R896 B.n390 B.n389 585
R897 B.n391 B.n102 585
R898 B.n393 B.n392 585
R899 B.n394 B.n101 585
R900 B.n396 B.n395 585
R901 B.n397 B.n100 585
R902 B.n399 B.n398 585
R903 B.n400 B.n99 585
R904 B.n402 B.n401 585
R905 B.n403 B.n98 585
R906 B.n405 B.n404 585
R907 B.n406 B.n97 585
R908 B.n408 B.n407 585
R909 B.n409 B.n96 585
R910 B.n411 B.n410 585
R911 B.n412 B.n95 585
R912 B.n414 B.n413 585
R913 B.n415 B.n94 585
R914 B.n417 B.n416 585
R915 B.n418 B.n93 585
R916 B.n420 B.n419 585
R917 B.n421 B.n92 585
R918 B.n423 B.n422 585
R919 B.n424 B.n91 585
R920 B.n426 B.n425 585
R921 B.n427 B.n90 585
R922 B.n429 B.n428 585
R923 B.n430 B.n89 585
R924 B.n432 B.n431 585
R925 B.n433 B.n88 585
R926 B.n435 B.n434 585
R927 B.n436 B.n87 585
R928 B.n438 B.n437 585
R929 B.n439 B.n86 585
R930 B.n441 B.n440 585
R931 B.n442 B.n85 585
R932 B.n444 B.n443 585
R933 B.n445 B.n84 585
R934 B.n447 B.n446 585
R935 B.n448 B.n83 585
R936 B.n450 B.n449 585
R937 B.n451 B.n82 585
R938 B.n453 B.n452 585
R939 B.n454 B.n81 585
R940 B.n456 B.n455 585
R941 B.n457 B.n80 585
R942 B.n459 B.n458 585
R943 B.n460 B.n79 585
R944 B.n462 B.n461 585
R945 B.n463 B.n78 585
R946 B.n465 B.n464 585
R947 B.n466 B.n77 585
R948 B.n468 B.n467 585
R949 B.n469 B.n76 585
R950 B.n639 B.n638 585
R951 B.n637 B.n16 585
R952 B.n636 B.n635 585
R953 B.n634 B.n17 585
R954 B.n633 B.n632 585
R955 B.n631 B.n18 585
R956 B.n630 B.n629 585
R957 B.n628 B.n19 585
R958 B.n627 B.n626 585
R959 B.n625 B.n20 585
R960 B.n624 B.n623 585
R961 B.n622 B.n21 585
R962 B.n621 B.n620 585
R963 B.n619 B.n22 585
R964 B.n618 B.n617 585
R965 B.n616 B.n23 585
R966 B.n615 B.n614 585
R967 B.n613 B.n24 585
R968 B.n612 B.n611 585
R969 B.n610 B.n25 585
R970 B.n609 B.n608 585
R971 B.n607 B.n26 585
R972 B.n606 B.n605 585
R973 B.n604 B.n27 585
R974 B.n603 B.n602 585
R975 B.n601 B.n28 585
R976 B.n600 B.n599 585
R977 B.n598 B.n29 585
R978 B.n597 B.n596 585
R979 B.n595 B.n30 585
R980 B.n594 B.n593 585
R981 B.n592 B.n31 585
R982 B.n591 B.n590 585
R983 B.n589 B.n32 585
R984 B.n588 B.n587 585
R985 B.n586 B.n33 585
R986 B.n585 B.n584 585
R987 B.n583 B.n34 585
R988 B.n582 B.n581 585
R989 B.n580 B.n35 585
R990 B.n579 B.n578 585
R991 B.n577 B.n36 585
R992 B.n576 B.n575 585
R993 B.n574 B.n37 585
R994 B.n573 B.n572 585
R995 B.n571 B.n38 585
R996 B.n570 B.n569 585
R997 B.n568 B.n39 585
R998 B.n567 B.n566 585
R999 B.n565 B.n40 585
R1000 B.n564 B.n563 585
R1001 B.n561 B.n41 585
R1002 B.n560 B.n559 585
R1003 B.n558 B.n44 585
R1004 B.n557 B.n556 585
R1005 B.n555 B.n45 585
R1006 B.n554 B.n553 585
R1007 B.n552 B.n46 585
R1008 B.n551 B.n550 585
R1009 B.n549 B.n47 585
R1010 B.n548 B.n547 585
R1011 B.n546 B.n545 585
R1012 B.n544 B.n51 585
R1013 B.n543 B.n542 585
R1014 B.n541 B.n52 585
R1015 B.n540 B.n539 585
R1016 B.n538 B.n53 585
R1017 B.n537 B.n536 585
R1018 B.n535 B.n54 585
R1019 B.n534 B.n533 585
R1020 B.n532 B.n55 585
R1021 B.n531 B.n530 585
R1022 B.n529 B.n56 585
R1023 B.n528 B.n527 585
R1024 B.n526 B.n57 585
R1025 B.n525 B.n524 585
R1026 B.n523 B.n58 585
R1027 B.n522 B.n521 585
R1028 B.n520 B.n59 585
R1029 B.n519 B.n518 585
R1030 B.n517 B.n60 585
R1031 B.n516 B.n515 585
R1032 B.n514 B.n61 585
R1033 B.n513 B.n512 585
R1034 B.n511 B.n62 585
R1035 B.n510 B.n509 585
R1036 B.n508 B.n63 585
R1037 B.n507 B.n506 585
R1038 B.n505 B.n64 585
R1039 B.n504 B.n503 585
R1040 B.n502 B.n65 585
R1041 B.n501 B.n500 585
R1042 B.n499 B.n66 585
R1043 B.n498 B.n497 585
R1044 B.n496 B.n67 585
R1045 B.n495 B.n494 585
R1046 B.n493 B.n68 585
R1047 B.n492 B.n491 585
R1048 B.n490 B.n69 585
R1049 B.n489 B.n488 585
R1050 B.n487 B.n70 585
R1051 B.n486 B.n485 585
R1052 B.n484 B.n71 585
R1053 B.n483 B.n482 585
R1054 B.n481 B.n72 585
R1055 B.n480 B.n479 585
R1056 B.n478 B.n73 585
R1057 B.n477 B.n476 585
R1058 B.n475 B.n74 585
R1059 B.n474 B.n473 585
R1060 B.n472 B.n75 585
R1061 B.n471 B.n470 585
R1062 B.n640 B.n15 585
R1063 B.n642 B.n641 585
R1064 B.n643 B.n14 585
R1065 B.n645 B.n644 585
R1066 B.n646 B.n13 585
R1067 B.n648 B.n647 585
R1068 B.n649 B.n12 585
R1069 B.n651 B.n650 585
R1070 B.n652 B.n11 585
R1071 B.n654 B.n653 585
R1072 B.n655 B.n10 585
R1073 B.n657 B.n656 585
R1074 B.n658 B.n9 585
R1075 B.n660 B.n659 585
R1076 B.n661 B.n8 585
R1077 B.n663 B.n662 585
R1078 B.n664 B.n7 585
R1079 B.n666 B.n665 585
R1080 B.n667 B.n6 585
R1081 B.n669 B.n668 585
R1082 B.n670 B.n5 585
R1083 B.n672 B.n671 585
R1084 B.n673 B.n4 585
R1085 B.n675 B.n674 585
R1086 B.n676 B.n3 585
R1087 B.n678 B.n677 585
R1088 B.n679 B.n0 585
R1089 B.n2 B.n1 585
R1090 B.n176 B.n175 585
R1091 B.n177 B.n174 585
R1092 B.n179 B.n178 585
R1093 B.n180 B.n173 585
R1094 B.n182 B.n181 585
R1095 B.n183 B.n172 585
R1096 B.n185 B.n184 585
R1097 B.n186 B.n171 585
R1098 B.n188 B.n187 585
R1099 B.n189 B.n170 585
R1100 B.n191 B.n190 585
R1101 B.n192 B.n169 585
R1102 B.n194 B.n193 585
R1103 B.n195 B.n168 585
R1104 B.n197 B.n196 585
R1105 B.n198 B.n167 585
R1106 B.n200 B.n199 585
R1107 B.n201 B.n166 585
R1108 B.n203 B.n202 585
R1109 B.n204 B.n165 585
R1110 B.n206 B.n205 585
R1111 B.n207 B.n164 585
R1112 B.n209 B.n208 585
R1113 B.n210 B.n163 585
R1114 B.n212 B.n211 585
R1115 B.n213 B.n162 585
R1116 B.n214 B.n213 578.989
R1117 B.n386 B.n385 578.989
R1118 B.n470 B.n469 578.989
R1119 B.n638 B.n15 578.989
R1120 B.n130 B.t1 500.38
R1121 B.n48 B.t8 500.38
R1122 B.n289 B.t4 500.38
R1123 B.n42 B.t11 500.38
R1124 B.n131 B.t2 435.604
R1125 B.n49 B.t7 435.604
R1126 B.n290 B.t5 435.604
R1127 B.n43 B.t10 435.604
R1128 B.n289 B.t3 331.413
R1129 B.n130 B.t0 331.413
R1130 B.n48 B.t6 331.413
R1131 B.n42 B.t9 331.413
R1132 B.n681 B.n680 256.663
R1133 B.n680 B.n679 235.042
R1134 B.n680 B.n2 235.042
R1135 B.n214 B.n161 163.367
R1136 B.n218 B.n161 163.367
R1137 B.n219 B.n218 163.367
R1138 B.n220 B.n219 163.367
R1139 B.n220 B.n159 163.367
R1140 B.n224 B.n159 163.367
R1141 B.n225 B.n224 163.367
R1142 B.n226 B.n225 163.367
R1143 B.n226 B.n157 163.367
R1144 B.n230 B.n157 163.367
R1145 B.n231 B.n230 163.367
R1146 B.n232 B.n231 163.367
R1147 B.n232 B.n155 163.367
R1148 B.n236 B.n155 163.367
R1149 B.n237 B.n236 163.367
R1150 B.n238 B.n237 163.367
R1151 B.n238 B.n153 163.367
R1152 B.n242 B.n153 163.367
R1153 B.n243 B.n242 163.367
R1154 B.n244 B.n243 163.367
R1155 B.n244 B.n151 163.367
R1156 B.n248 B.n151 163.367
R1157 B.n249 B.n248 163.367
R1158 B.n250 B.n249 163.367
R1159 B.n250 B.n149 163.367
R1160 B.n254 B.n149 163.367
R1161 B.n255 B.n254 163.367
R1162 B.n256 B.n255 163.367
R1163 B.n256 B.n147 163.367
R1164 B.n260 B.n147 163.367
R1165 B.n261 B.n260 163.367
R1166 B.n262 B.n261 163.367
R1167 B.n262 B.n145 163.367
R1168 B.n266 B.n145 163.367
R1169 B.n267 B.n266 163.367
R1170 B.n268 B.n267 163.367
R1171 B.n268 B.n143 163.367
R1172 B.n272 B.n143 163.367
R1173 B.n273 B.n272 163.367
R1174 B.n274 B.n273 163.367
R1175 B.n274 B.n141 163.367
R1176 B.n278 B.n141 163.367
R1177 B.n279 B.n278 163.367
R1178 B.n280 B.n279 163.367
R1179 B.n280 B.n139 163.367
R1180 B.n284 B.n139 163.367
R1181 B.n285 B.n284 163.367
R1182 B.n286 B.n285 163.367
R1183 B.n286 B.n137 163.367
R1184 B.n293 B.n137 163.367
R1185 B.n294 B.n293 163.367
R1186 B.n295 B.n294 163.367
R1187 B.n295 B.n135 163.367
R1188 B.n299 B.n135 163.367
R1189 B.n300 B.n299 163.367
R1190 B.n301 B.n300 163.367
R1191 B.n301 B.n133 163.367
R1192 B.n305 B.n133 163.367
R1193 B.n306 B.n305 163.367
R1194 B.n307 B.n306 163.367
R1195 B.n307 B.n129 163.367
R1196 B.n312 B.n129 163.367
R1197 B.n313 B.n312 163.367
R1198 B.n314 B.n313 163.367
R1199 B.n314 B.n127 163.367
R1200 B.n318 B.n127 163.367
R1201 B.n319 B.n318 163.367
R1202 B.n320 B.n319 163.367
R1203 B.n320 B.n125 163.367
R1204 B.n324 B.n125 163.367
R1205 B.n325 B.n324 163.367
R1206 B.n326 B.n325 163.367
R1207 B.n326 B.n123 163.367
R1208 B.n330 B.n123 163.367
R1209 B.n331 B.n330 163.367
R1210 B.n332 B.n331 163.367
R1211 B.n332 B.n121 163.367
R1212 B.n336 B.n121 163.367
R1213 B.n337 B.n336 163.367
R1214 B.n338 B.n337 163.367
R1215 B.n338 B.n119 163.367
R1216 B.n342 B.n119 163.367
R1217 B.n343 B.n342 163.367
R1218 B.n344 B.n343 163.367
R1219 B.n344 B.n117 163.367
R1220 B.n348 B.n117 163.367
R1221 B.n349 B.n348 163.367
R1222 B.n350 B.n349 163.367
R1223 B.n350 B.n115 163.367
R1224 B.n354 B.n115 163.367
R1225 B.n355 B.n354 163.367
R1226 B.n356 B.n355 163.367
R1227 B.n356 B.n113 163.367
R1228 B.n360 B.n113 163.367
R1229 B.n361 B.n360 163.367
R1230 B.n362 B.n361 163.367
R1231 B.n362 B.n111 163.367
R1232 B.n366 B.n111 163.367
R1233 B.n367 B.n366 163.367
R1234 B.n368 B.n367 163.367
R1235 B.n368 B.n109 163.367
R1236 B.n372 B.n109 163.367
R1237 B.n373 B.n372 163.367
R1238 B.n374 B.n373 163.367
R1239 B.n374 B.n107 163.367
R1240 B.n378 B.n107 163.367
R1241 B.n379 B.n378 163.367
R1242 B.n380 B.n379 163.367
R1243 B.n380 B.n105 163.367
R1244 B.n384 B.n105 163.367
R1245 B.n385 B.n384 163.367
R1246 B.n469 B.n468 163.367
R1247 B.n468 B.n77 163.367
R1248 B.n464 B.n77 163.367
R1249 B.n464 B.n463 163.367
R1250 B.n463 B.n462 163.367
R1251 B.n462 B.n79 163.367
R1252 B.n458 B.n79 163.367
R1253 B.n458 B.n457 163.367
R1254 B.n457 B.n456 163.367
R1255 B.n456 B.n81 163.367
R1256 B.n452 B.n81 163.367
R1257 B.n452 B.n451 163.367
R1258 B.n451 B.n450 163.367
R1259 B.n450 B.n83 163.367
R1260 B.n446 B.n83 163.367
R1261 B.n446 B.n445 163.367
R1262 B.n445 B.n444 163.367
R1263 B.n444 B.n85 163.367
R1264 B.n440 B.n85 163.367
R1265 B.n440 B.n439 163.367
R1266 B.n439 B.n438 163.367
R1267 B.n438 B.n87 163.367
R1268 B.n434 B.n87 163.367
R1269 B.n434 B.n433 163.367
R1270 B.n433 B.n432 163.367
R1271 B.n432 B.n89 163.367
R1272 B.n428 B.n89 163.367
R1273 B.n428 B.n427 163.367
R1274 B.n427 B.n426 163.367
R1275 B.n426 B.n91 163.367
R1276 B.n422 B.n91 163.367
R1277 B.n422 B.n421 163.367
R1278 B.n421 B.n420 163.367
R1279 B.n420 B.n93 163.367
R1280 B.n416 B.n93 163.367
R1281 B.n416 B.n415 163.367
R1282 B.n415 B.n414 163.367
R1283 B.n414 B.n95 163.367
R1284 B.n410 B.n95 163.367
R1285 B.n410 B.n409 163.367
R1286 B.n409 B.n408 163.367
R1287 B.n408 B.n97 163.367
R1288 B.n404 B.n97 163.367
R1289 B.n404 B.n403 163.367
R1290 B.n403 B.n402 163.367
R1291 B.n402 B.n99 163.367
R1292 B.n398 B.n99 163.367
R1293 B.n398 B.n397 163.367
R1294 B.n397 B.n396 163.367
R1295 B.n396 B.n101 163.367
R1296 B.n392 B.n101 163.367
R1297 B.n392 B.n391 163.367
R1298 B.n391 B.n390 163.367
R1299 B.n390 B.n103 163.367
R1300 B.n386 B.n103 163.367
R1301 B.n638 B.n637 163.367
R1302 B.n637 B.n636 163.367
R1303 B.n636 B.n17 163.367
R1304 B.n632 B.n17 163.367
R1305 B.n632 B.n631 163.367
R1306 B.n631 B.n630 163.367
R1307 B.n630 B.n19 163.367
R1308 B.n626 B.n19 163.367
R1309 B.n626 B.n625 163.367
R1310 B.n625 B.n624 163.367
R1311 B.n624 B.n21 163.367
R1312 B.n620 B.n21 163.367
R1313 B.n620 B.n619 163.367
R1314 B.n619 B.n618 163.367
R1315 B.n618 B.n23 163.367
R1316 B.n614 B.n23 163.367
R1317 B.n614 B.n613 163.367
R1318 B.n613 B.n612 163.367
R1319 B.n612 B.n25 163.367
R1320 B.n608 B.n25 163.367
R1321 B.n608 B.n607 163.367
R1322 B.n607 B.n606 163.367
R1323 B.n606 B.n27 163.367
R1324 B.n602 B.n27 163.367
R1325 B.n602 B.n601 163.367
R1326 B.n601 B.n600 163.367
R1327 B.n600 B.n29 163.367
R1328 B.n596 B.n29 163.367
R1329 B.n596 B.n595 163.367
R1330 B.n595 B.n594 163.367
R1331 B.n594 B.n31 163.367
R1332 B.n590 B.n31 163.367
R1333 B.n590 B.n589 163.367
R1334 B.n589 B.n588 163.367
R1335 B.n588 B.n33 163.367
R1336 B.n584 B.n33 163.367
R1337 B.n584 B.n583 163.367
R1338 B.n583 B.n582 163.367
R1339 B.n582 B.n35 163.367
R1340 B.n578 B.n35 163.367
R1341 B.n578 B.n577 163.367
R1342 B.n577 B.n576 163.367
R1343 B.n576 B.n37 163.367
R1344 B.n572 B.n37 163.367
R1345 B.n572 B.n571 163.367
R1346 B.n571 B.n570 163.367
R1347 B.n570 B.n39 163.367
R1348 B.n566 B.n39 163.367
R1349 B.n566 B.n565 163.367
R1350 B.n565 B.n564 163.367
R1351 B.n564 B.n41 163.367
R1352 B.n559 B.n41 163.367
R1353 B.n559 B.n558 163.367
R1354 B.n558 B.n557 163.367
R1355 B.n557 B.n45 163.367
R1356 B.n553 B.n45 163.367
R1357 B.n553 B.n552 163.367
R1358 B.n552 B.n551 163.367
R1359 B.n551 B.n47 163.367
R1360 B.n547 B.n47 163.367
R1361 B.n547 B.n546 163.367
R1362 B.n546 B.n51 163.367
R1363 B.n542 B.n51 163.367
R1364 B.n542 B.n541 163.367
R1365 B.n541 B.n540 163.367
R1366 B.n540 B.n53 163.367
R1367 B.n536 B.n53 163.367
R1368 B.n536 B.n535 163.367
R1369 B.n535 B.n534 163.367
R1370 B.n534 B.n55 163.367
R1371 B.n530 B.n55 163.367
R1372 B.n530 B.n529 163.367
R1373 B.n529 B.n528 163.367
R1374 B.n528 B.n57 163.367
R1375 B.n524 B.n57 163.367
R1376 B.n524 B.n523 163.367
R1377 B.n523 B.n522 163.367
R1378 B.n522 B.n59 163.367
R1379 B.n518 B.n59 163.367
R1380 B.n518 B.n517 163.367
R1381 B.n517 B.n516 163.367
R1382 B.n516 B.n61 163.367
R1383 B.n512 B.n61 163.367
R1384 B.n512 B.n511 163.367
R1385 B.n511 B.n510 163.367
R1386 B.n510 B.n63 163.367
R1387 B.n506 B.n63 163.367
R1388 B.n506 B.n505 163.367
R1389 B.n505 B.n504 163.367
R1390 B.n504 B.n65 163.367
R1391 B.n500 B.n65 163.367
R1392 B.n500 B.n499 163.367
R1393 B.n499 B.n498 163.367
R1394 B.n498 B.n67 163.367
R1395 B.n494 B.n67 163.367
R1396 B.n494 B.n493 163.367
R1397 B.n493 B.n492 163.367
R1398 B.n492 B.n69 163.367
R1399 B.n488 B.n69 163.367
R1400 B.n488 B.n487 163.367
R1401 B.n487 B.n486 163.367
R1402 B.n486 B.n71 163.367
R1403 B.n482 B.n71 163.367
R1404 B.n482 B.n481 163.367
R1405 B.n481 B.n480 163.367
R1406 B.n480 B.n73 163.367
R1407 B.n476 B.n73 163.367
R1408 B.n476 B.n475 163.367
R1409 B.n475 B.n474 163.367
R1410 B.n474 B.n75 163.367
R1411 B.n470 B.n75 163.367
R1412 B.n642 B.n15 163.367
R1413 B.n643 B.n642 163.367
R1414 B.n644 B.n643 163.367
R1415 B.n644 B.n13 163.367
R1416 B.n648 B.n13 163.367
R1417 B.n649 B.n648 163.367
R1418 B.n650 B.n649 163.367
R1419 B.n650 B.n11 163.367
R1420 B.n654 B.n11 163.367
R1421 B.n655 B.n654 163.367
R1422 B.n656 B.n655 163.367
R1423 B.n656 B.n9 163.367
R1424 B.n660 B.n9 163.367
R1425 B.n661 B.n660 163.367
R1426 B.n662 B.n661 163.367
R1427 B.n662 B.n7 163.367
R1428 B.n666 B.n7 163.367
R1429 B.n667 B.n666 163.367
R1430 B.n668 B.n667 163.367
R1431 B.n668 B.n5 163.367
R1432 B.n672 B.n5 163.367
R1433 B.n673 B.n672 163.367
R1434 B.n674 B.n673 163.367
R1435 B.n674 B.n3 163.367
R1436 B.n678 B.n3 163.367
R1437 B.n679 B.n678 163.367
R1438 B.n176 B.n2 163.367
R1439 B.n177 B.n176 163.367
R1440 B.n178 B.n177 163.367
R1441 B.n178 B.n173 163.367
R1442 B.n182 B.n173 163.367
R1443 B.n183 B.n182 163.367
R1444 B.n184 B.n183 163.367
R1445 B.n184 B.n171 163.367
R1446 B.n188 B.n171 163.367
R1447 B.n189 B.n188 163.367
R1448 B.n190 B.n189 163.367
R1449 B.n190 B.n169 163.367
R1450 B.n194 B.n169 163.367
R1451 B.n195 B.n194 163.367
R1452 B.n196 B.n195 163.367
R1453 B.n196 B.n167 163.367
R1454 B.n200 B.n167 163.367
R1455 B.n201 B.n200 163.367
R1456 B.n202 B.n201 163.367
R1457 B.n202 B.n165 163.367
R1458 B.n206 B.n165 163.367
R1459 B.n207 B.n206 163.367
R1460 B.n208 B.n207 163.367
R1461 B.n208 B.n163 163.367
R1462 B.n212 B.n163 163.367
R1463 B.n213 B.n212 163.367
R1464 B.n290 B.n289 64.7763
R1465 B.n131 B.n130 64.7763
R1466 B.n49 B.n48 64.7763
R1467 B.n43 B.n42 64.7763
R1468 B.n291 B.n290 59.5399
R1469 B.n309 B.n131 59.5399
R1470 B.n50 B.n49 59.5399
R1471 B.n562 B.n43 59.5399
R1472 B.n640 B.n639 37.62
R1473 B.n471 B.n76 37.62
R1474 B.n387 B.n104 37.62
R1475 B.n215 B.n162 37.62
R1476 B B.n681 18.0485
R1477 B.n641 B.n640 10.6151
R1478 B.n641 B.n14 10.6151
R1479 B.n645 B.n14 10.6151
R1480 B.n646 B.n645 10.6151
R1481 B.n647 B.n646 10.6151
R1482 B.n647 B.n12 10.6151
R1483 B.n651 B.n12 10.6151
R1484 B.n652 B.n651 10.6151
R1485 B.n653 B.n652 10.6151
R1486 B.n653 B.n10 10.6151
R1487 B.n657 B.n10 10.6151
R1488 B.n658 B.n657 10.6151
R1489 B.n659 B.n658 10.6151
R1490 B.n659 B.n8 10.6151
R1491 B.n663 B.n8 10.6151
R1492 B.n664 B.n663 10.6151
R1493 B.n665 B.n664 10.6151
R1494 B.n665 B.n6 10.6151
R1495 B.n669 B.n6 10.6151
R1496 B.n670 B.n669 10.6151
R1497 B.n671 B.n670 10.6151
R1498 B.n671 B.n4 10.6151
R1499 B.n675 B.n4 10.6151
R1500 B.n676 B.n675 10.6151
R1501 B.n677 B.n676 10.6151
R1502 B.n677 B.n0 10.6151
R1503 B.n639 B.n16 10.6151
R1504 B.n635 B.n16 10.6151
R1505 B.n635 B.n634 10.6151
R1506 B.n634 B.n633 10.6151
R1507 B.n633 B.n18 10.6151
R1508 B.n629 B.n18 10.6151
R1509 B.n629 B.n628 10.6151
R1510 B.n628 B.n627 10.6151
R1511 B.n627 B.n20 10.6151
R1512 B.n623 B.n20 10.6151
R1513 B.n623 B.n622 10.6151
R1514 B.n622 B.n621 10.6151
R1515 B.n621 B.n22 10.6151
R1516 B.n617 B.n22 10.6151
R1517 B.n617 B.n616 10.6151
R1518 B.n616 B.n615 10.6151
R1519 B.n615 B.n24 10.6151
R1520 B.n611 B.n24 10.6151
R1521 B.n611 B.n610 10.6151
R1522 B.n610 B.n609 10.6151
R1523 B.n609 B.n26 10.6151
R1524 B.n605 B.n26 10.6151
R1525 B.n605 B.n604 10.6151
R1526 B.n604 B.n603 10.6151
R1527 B.n603 B.n28 10.6151
R1528 B.n599 B.n28 10.6151
R1529 B.n599 B.n598 10.6151
R1530 B.n598 B.n597 10.6151
R1531 B.n597 B.n30 10.6151
R1532 B.n593 B.n30 10.6151
R1533 B.n593 B.n592 10.6151
R1534 B.n592 B.n591 10.6151
R1535 B.n591 B.n32 10.6151
R1536 B.n587 B.n32 10.6151
R1537 B.n587 B.n586 10.6151
R1538 B.n586 B.n585 10.6151
R1539 B.n585 B.n34 10.6151
R1540 B.n581 B.n34 10.6151
R1541 B.n581 B.n580 10.6151
R1542 B.n580 B.n579 10.6151
R1543 B.n579 B.n36 10.6151
R1544 B.n575 B.n36 10.6151
R1545 B.n575 B.n574 10.6151
R1546 B.n574 B.n573 10.6151
R1547 B.n573 B.n38 10.6151
R1548 B.n569 B.n38 10.6151
R1549 B.n569 B.n568 10.6151
R1550 B.n568 B.n567 10.6151
R1551 B.n567 B.n40 10.6151
R1552 B.n563 B.n40 10.6151
R1553 B.n561 B.n560 10.6151
R1554 B.n560 B.n44 10.6151
R1555 B.n556 B.n44 10.6151
R1556 B.n556 B.n555 10.6151
R1557 B.n555 B.n554 10.6151
R1558 B.n554 B.n46 10.6151
R1559 B.n550 B.n46 10.6151
R1560 B.n550 B.n549 10.6151
R1561 B.n549 B.n548 10.6151
R1562 B.n545 B.n544 10.6151
R1563 B.n544 B.n543 10.6151
R1564 B.n543 B.n52 10.6151
R1565 B.n539 B.n52 10.6151
R1566 B.n539 B.n538 10.6151
R1567 B.n538 B.n537 10.6151
R1568 B.n537 B.n54 10.6151
R1569 B.n533 B.n54 10.6151
R1570 B.n533 B.n532 10.6151
R1571 B.n532 B.n531 10.6151
R1572 B.n531 B.n56 10.6151
R1573 B.n527 B.n56 10.6151
R1574 B.n527 B.n526 10.6151
R1575 B.n526 B.n525 10.6151
R1576 B.n525 B.n58 10.6151
R1577 B.n521 B.n58 10.6151
R1578 B.n521 B.n520 10.6151
R1579 B.n520 B.n519 10.6151
R1580 B.n519 B.n60 10.6151
R1581 B.n515 B.n60 10.6151
R1582 B.n515 B.n514 10.6151
R1583 B.n514 B.n513 10.6151
R1584 B.n513 B.n62 10.6151
R1585 B.n509 B.n62 10.6151
R1586 B.n509 B.n508 10.6151
R1587 B.n508 B.n507 10.6151
R1588 B.n507 B.n64 10.6151
R1589 B.n503 B.n64 10.6151
R1590 B.n503 B.n502 10.6151
R1591 B.n502 B.n501 10.6151
R1592 B.n501 B.n66 10.6151
R1593 B.n497 B.n66 10.6151
R1594 B.n497 B.n496 10.6151
R1595 B.n496 B.n495 10.6151
R1596 B.n495 B.n68 10.6151
R1597 B.n491 B.n68 10.6151
R1598 B.n491 B.n490 10.6151
R1599 B.n490 B.n489 10.6151
R1600 B.n489 B.n70 10.6151
R1601 B.n485 B.n70 10.6151
R1602 B.n485 B.n484 10.6151
R1603 B.n484 B.n483 10.6151
R1604 B.n483 B.n72 10.6151
R1605 B.n479 B.n72 10.6151
R1606 B.n479 B.n478 10.6151
R1607 B.n478 B.n477 10.6151
R1608 B.n477 B.n74 10.6151
R1609 B.n473 B.n74 10.6151
R1610 B.n473 B.n472 10.6151
R1611 B.n472 B.n471 10.6151
R1612 B.n467 B.n76 10.6151
R1613 B.n467 B.n466 10.6151
R1614 B.n466 B.n465 10.6151
R1615 B.n465 B.n78 10.6151
R1616 B.n461 B.n78 10.6151
R1617 B.n461 B.n460 10.6151
R1618 B.n460 B.n459 10.6151
R1619 B.n459 B.n80 10.6151
R1620 B.n455 B.n80 10.6151
R1621 B.n455 B.n454 10.6151
R1622 B.n454 B.n453 10.6151
R1623 B.n453 B.n82 10.6151
R1624 B.n449 B.n82 10.6151
R1625 B.n449 B.n448 10.6151
R1626 B.n448 B.n447 10.6151
R1627 B.n447 B.n84 10.6151
R1628 B.n443 B.n84 10.6151
R1629 B.n443 B.n442 10.6151
R1630 B.n442 B.n441 10.6151
R1631 B.n441 B.n86 10.6151
R1632 B.n437 B.n86 10.6151
R1633 B.n437 B.n436 10.6151
R1634 B.n436 B.n435 10.6151
R1635 B.n435 B.n88 10.6151
R1636 B.n431 B.n88 10.6151
R1637 B.n431 B.n430 10.6151
R1638 B.n430 B.n429 10.6151
R1639 B.n429 B.n90 10.6151
R1640 B.n425 B.n90 10.6151
R1641 B.n425 B.n424 10.6151
R1642 B.n424 B.n423 10.6151
R1643 B.n423 B.n92 10.6151
R1644 B.n419 B.n92 10.6151
R1645 B.n419 B.n418 10.6151
R1646 B.n418 B.n417 10.6151
R1647 B.n417 B.n94 10.6151
R1648 B.n413 B.n94 10.6151
R1649 B.n413 B.n412 10.6151
R1650 B.n412 B.n411 10.6151
R1651 B.n411 B.n96 10.6151
R1652 B.n407 B.n96 10.6151
R1653 B.n407 B.n406 10.6151
R1654 B.n406 B.n405 10.6151
R1655 B.n405 B.n98 10.6151
R1656 B.n401 B.n98 10.6151
R1657 B.n401 B.n400 10.6151
R1658 B.n400 B.n399 10.6151
R1659 B.n399 B.n100 10.6151
R1660 B.n395 B.n100 10.6151
R1661 B.n395 B.n394 10.6151
R1662 B.n394 B.n393 10.6151
R1663 B.n393 B.n102 10.6151
R1664 B.n389 B.n102 10.6151
R1665 B.n389 B.n388 10.6151
R1666 B.n388 B.n387 10.6151
R1667 B.n175 B.n1 10.6151
R1668 B.n175 B.n174 10.6151
R1669 B.n179 B.n174 10.6151
R1670 B.n180 B.n179 10.6151
R1671 B.n181 B.n180 10.6151
R1672 B.n181 B.n172 10.6151
R1673 B.n185 B.n172 10.6151
R1674 B.n186 B.n185 10.6151
R1675 B.n187 B.n186 10.6151
R1676 B.n187 B.n170 10.6151
R1677 B.n191 B.n170 10.6151
R1678 B.n192 B.n191 10.6151
R1679 B.n193 B.n192 10.6151
R1680 B.n193 B.n168 10.6151
R1681 B.n197 B.n168 10.6151
R1682 B.n198 B.n197 10.6151
R1683 B.n199 B.n198 10.6151
R1684 B.n199 B.n166 10.6151
R1685 B.n203 B.n166 10.6151
R1686 B.n204 B.n203 10.6151
R1687 B.n205 B.n204 10.6151
R1688 B.n205 B.n164 10.6151
R1689 B.n209 B.n164 10.6151
R1690 B.n210 B.n209 10.6151
R1691 B.n211 B.n210 10.6151
R1692 B.n211 B.n162 10.6151
R1693 B.n216 B.n215 10.6151
R1694 B.n217 B.n216 10.6151
R1695 B.n217 B.n160 10.6151
R1696 B.n221 B.n160 10.6151
R1697 B.n222 B.n221 10.6151
R1698 B.n223 B.n222 10.6151
R1699 B.n223 B.n158 10.6151
R1700 B.n227 B.n158 10.6151
R1701 B.n228 B.n227 10.6151
R1702 B.n229 B.n228 10.6151
R1703 B.n229 B.n156 10.6151
R1704 B.n233 B.n156 10.6151
R1705 B.n234 B.n233 10.6151
R1706 B.n235 B.n234 10.6151
R1707 B.n235 B.n154 10.6151
R1708 B.n239 B.n154 10.6151
R1709 B.n240 B.n239 10.6151
R1710 B.n241 B.n240 10.6151
R1711 B.n241 B.n152 10.6151
R1712 B.n245 B.n152 10.6151
R1713 B.n246 B.n245 10.6151
R1714 B.n247 B.n246 10.6151
R1715 B.n247 B.n150 10.6151
R1716 B.n251 B.n150 10.6151
R1717 B.n252 B.n251 10.6151
R1718 B.n253 B.n252 10.6151
R1719 B.n253 B.n148 10.6151
R1720 B.n257 B.n148 10.6151
R1721 B.n258 B.n257 10.6151
R1722 B.n259 B.n258 10.6151
R1723 B.n259 B.n146 10.6151
R1724 B.n263 B.n146 10.6151
R1725 B.n264 B.n263 10.6151
R1726 B.n265 B.n264 10.6151
R1727 B.n265 B.n144 10.6151
R1728 B.n269 B.n144 10.6151
R1729 B.n270 B.n269 10.6151
R1730 B.n271 B.n270 10.6151
R1731 B.n271 B.n142 10.6151
R1732 B.n275 B.n142 10.6151
R1733 B.n276 B.n275 10.6151
R1734 B.n277 B.n276 10.6151
R1735 B.n277 B.n140 10.6151
R1736 B.n281 B.n140 10.6151
R1737 B.n282 B.n281 10.6151
R1738 B.n283 B.n282 10.6151
R1739 B.n283 B.n138 10.6151
R1740 B.n287 B.n138 10.6151
R1741 B.n288 B.n287 10.6151
R1742 B.n292 B.n288 10.6151
R1743 B.n296 B.n136 10.6151
R1744 B.n297 B.n296 10.6151
R1745 B.n298 B.n297 10.6151
R1746 B.n298 B.n134 10.6151
R1747 B.n302 B.n134 10.6151
R1748 B.n303 B.n302 10.6151
R1749 B.n304 B.n303 10.6151
R1750 B.n304 B.n132 10.6151
R1751 B.n308 B.n132 10.6151
R1752 B.n311 B.n310 10.6151
R1753 B.n311 B.n128 10.6151
R1754 B.n315 B.n128 10.6151
R1755 B.n316 B.n315 10.6151
R1756 B.n317 B.n316 10.6151
R1757 B.n317 B.n126 10.6151
R1758 B.n321 B.n126 10.6151
R1759 B.n322 B.n321 10.6151
R1760 B.n323 B.n322 10.6151
R1761 B.n323 B.n124 10.6151
R1762 B.n327 B.n124 10.6151
R1763 B.n328 B.n327 10.6151
R1764 B.n329 B.n328 10.6151
R1765 B.n329 B.n122 10.6151
R1766 B.n333 B.n122 10.6151
R1767 B.n334 B.n333 10.6151
R1768 B.n335 B.n334 10.6151
R1769 B.n335 B.n120 10.6151
R1770 B.n339 B.n120 10.6151
R1771 B.n340 B.n339 10.6151
R1772 B.n341 B.n340 10.6151
R1773 B.n341 B.n118 10.6151
R1774 B.n345 B.n118 10.6151
R1775 B.n346 B.n345 10.6151
R1776 B.n347 B.n346 10.6151
R1777 B.n347 B.n116 10.6151
R1778 B.n351 B.n116 10.6151
R1779 B.n352 B.n351 10.6151
R1780 B.n353 B.n352 10.6151
R1781 B.n353 B.n114 10.6151
R1782 B.n357 B.n114 10.6151
R1783 B.n358 B.n357 10.6151
R1784 B.n359 B.n358 10.6151
R1785 B.n359 B.n112 10.6151
R1786 B.n363 B.n112 10.6151
R1787 B.n364 B.n363 10.6151
R1788 B.n365 B.n364 10.6151
R1789 B.n365 B.n110 10.6151
R1790 B.n369 B.n110 10.6151
R1791 B.n370 B.n369 10.6151
R1792 B.n371 B.n370 10.6151
R1793 B.n371 B.n108 10.6151
R1794 B.n375 B.n108 10.6151
R1795 B.n376 B.n375 10.6151
R1796 B.n377 B.n376 10.6151
R1797 B.n377 B.n106 10.6151
R1798 B.n381 B.n106 10.6151
R1799 B.n382 B.n381 10.6151
R1800 B.n383 B.n382 10.6151
R1801 B.n383 B.n104 10.6151
R1802 B.n563 B.n562 9.36635
R1803 B.n545 B.n50 9.36635
R1804 B.n292 B.n291 9.36635
R1805 B.n310 B.n309 9.36635
R1806 B.n681 B.n0 8.11757
R1807 B.n681 B.n1 8.11757
R1808 B.n562 B.n561 1.24928
R1809 B.n548 B.n50 1.24928
R1810 B.n291 B.n136 1.24928
R1811 B.n309 B.n308 1.24928
R1812 VP.n0 VP.t1 212.234
R1813 VP.n0 VP.t0 163.96
R1814 VP VP.n0 0.431812
R1815 VDD1.n80 VDD1.n0 756.745
R1816 VDD1.n165 VDD1.n85 756.745
R1817 VDD1.n81 VDD1.n80 585
R1818 VDD1.n79 VDD1.n78 585
R1819 VDD1.n4 VDD1.n3 585
R1820 VDD1.n8 VDD1.n6 585
R1821 VDD1.n73 VDD1.n72 585
R1822 VDD1.n71 VDD1.n70 585
R1823 VDD1.n10 VDD1.n9 585
R1824 VDD1.n65 VDD1.n64 585
R1825 VDD1.n63 VDD1.n62 585
R1826 VDD1.n14 VDD1.n13 585
R1827 VDD1.n57 VDD1.n56 585
R1828 VDD1.n55 VDD1.n54 585
R1829 VDD1.n18 VDD1.n17 585
R1830 VDD1.n49 VDD1.n48 585
R1831 VDD1.n47 VDD1.n46 585
R1832 VDD1.n22 VDD1.n21 585
R1833 VDD1.n41 VDD1.n40 585
R1834 VDD1.n39 VDD1.n38 585
R1835 VDD1.n26 VDD1.n25 585
R1836 VDD1.n33 VDD1.n32 585
R1837 VDD1.n31 VDD1.n30 585
R1838 VDD1.n114 VDD1.n113 585
R1839 VDD1.n116 VDD1.n115 585
R1840 VDD1.n109 VDD1.n108 585
R1841 VDD1.n122 VDD1.n121 585
R1842 VDD1.n124 VDD1.n123 585
R1843 VDD1.n105 VDD1.n104 585
R1844 VDD1.n130 VDD1.n129 585
R1845 VDD1.n132 VDD1.n131 585
R1846 VDD1.n101 VDD1.n100 585
R1847 VDD1.n138 VDD1.n137 585
R1848 VDD1.n140 VDD1.n139 585
R1849 VDD1.n97 VDD1.n96 585
R1850 VDD1.n146 VDD1.n145 585
R1851 VDD1.n148 VDD1.n147 585
R1852 VDD1.n93 VDD1.n92 585
R1853 VDD1.n155 VDD1.n154 585
R1854 VDD1.n156 VDD1.n91 585
R1855 VDD1.n158 VDD1.n157 585
R1856 VDD1.n89 VDD1.n88 585
R1857 VDD1.n164 VDD1.n163 585
R1858 VDD1.n166 VDD1.n165 585
R1859 VDD1.n29 VDD1.t0 327.466
R1860 VDD1.n112 VDD1.t1 327.466
R1861 VDD1.n80 VDD1.n79 171.744
R1862 VDD1.n79 VDD1.n3 171.744
R1863 VDD1.n8 VDD1.n3 171.744
R1864 VDD1.n72 VDD1.n8 171.744
R1865 VDD1.n72 VDD1.n71 171.744
R1866 VDD1.n71 VDD1.n9 171.744
R1867 VDD1.n64 VDD1.n9 171.744
R1868 VDD1.n64 VDD1.n63 171.744
R1869 VDD1.n63 VDD1.n13 171.744
R1870 VDD1.n56 VDD1.n13 171.744
R1871 VDD1.n56 VDD1.n55 171.744
R1872 VDD1.n55 VDD1.n17 171.744
R1873 VDD1.n48 VDD1.n17 171.744
R1874 VDD1.n48 VDD1.n47 171.744
R1875 VDD1.n47 VDD1.n21 171.744
R1876 VDD1.n40 VDD1.n21 171.744
R1877 VDD1.n40 VDD1.n39 171.744
R1878 VDD1.n39 VDD1.n25 171.744
R1879 VDD1.n32 VDD1.n25 171.744
R1880 VDD1.n32 VDD1.n31 171.744
R1881 VDD1.n115 VDD1.n114 171.744
R1882 VDD1.n115 VDD1.n108 171.744
R1883 VDD1.n122 VDD1.n108 171.744
R1884 VDD1.n123 VDD1.n122 171.744
R1885 VDD1.n123 VDD1.n104 171.744
R1886 VDD1.n130 VDD1.n104 171.744
R1887 VDD1.n131 VDD1.n130 171.744
R1888 VDD1.n131 VDD1.n100 171.744
R1889 VDD1.n138 VDD1.n100 171.744
R1890 VDD1.n139 VDD1.n138 171.744
R1891 VDD1.n139 VDD1.n96 171.744
R1892 VDD1.n146 VDD1.n96 171.744
R1893 VDD1.n147 VDD1.n146 171.744
R1894 VDD1.n147 VDD1.n92 171.744
R1895 VDD1.n155 VDD1.n92 171.744
R1896 VDD1.n156 VDD1.n155 171.744
R1897 VDD1.n157 VDD1.n156 171.744
R1898 VDD1.n157 VDD1.n88 171.744
R1899 VDD1.n164 VDD1.n88 171.744
R1900 VDD1.n165 VDD1.n164 171.744
R1901 VDD1 VDD1.n169 92.3631
R1902 VDD1.n31 VDD1.t0 85.8723
R1903 VDD1.n114 VDD1.t1 85.8723
R1904 VDD1 VDD1.n84 49.2543
R1905 VDD1.n30 VDD1.n29 16.3895
R1906 VDD1.n113 VDD1.n112 16.3895
R1907 VDD1.n6 VDD1.n4 13.1884
R1908 VDD1.n158 VDD1.n89 13.1884
R1909 VDD1.n78 VDD1.n77 12.8005
R1910 VDD1.n74 VDD1.n73 12.8005
R1911 VDD1.n33 VDD1.n28 12.8005
R1912 VDD1.n116 VDD1.n111 12.8005
R1913 VDD1.n159 VDD1.n91 12.8005
R1914 VDD1.n163 VDD1.n162 12.8005
R1915 VDD1.n81 VDD1.n2 12.0247
R1916 VDD1.n70 VDD1.n7 12.0247
R1917 VDD1.n34 VDD1.n26 12.0247
R1918 VDD1.n117 VDD1.n109 12.0247
R1919 VDD1.n154 VDD1.n153 12.0247
R1920 VDD1.n166 VDD1.n87 12.0247
R1921 VDD1.n82 VDD1.n0 11.249
R1922 VDD1.n69 VDD1.n10 11.249
R1923 VDD1.n38 VDD1.n37 11.249
R1924 VDD1.n121 VDD1.n120 11.249
R1925 VDD1.n152 VDD1.n93 11.249
R1926 VDD1.n167 VDD1.n85 11.249
R1927 VDD1.n66 VDD1.n65 10.4732
R1928 VDD1.n41 VDD1.n24 10.4732
R1929 VDD1.n124 VDD1.n107 10.4732
R1930 VDD1.n149 VDD1.n148 10.4732
R1931 VDD1.n62 VDD1.n12 9.69747
R1932 VDD1.n42 VDD1.n22 9.69747
R1933 VDD1.n125 VDD1.n105 9.69747
R1934 VDD1.n145 VDD1.n95 9.69747
R1935 VDD1.n84 VDD1.n83 9.45567
R1936 VDD1.n169 VDD1.n168 9.45567
R1937 VDD1.n16 VDD1.n15 9.3005
R1938 VDD1.n59 VDD1.n58 9.3005
R1939 VDD1.n61 VDD1.n60 9.3005
R1940 VDD1.n12 VDD1.n11 9.3005
R1941 VDD1.n67 VDD1.n66 9.3005
R1942 VDD1.n69 VDD1.n68 9.3005
R1943 VDD1.n7 VDD1.n5 9.3005
R1944 VDD1.n75 VDD1.n74 9.3005
R1945 VDD1.n83 VDD1.n82 9.3005
R1946 VDD1.n2 VDD1.n1 9.3005
R1947 VDD1.n77 VDD1.n76 9.3005
R1948 VDD1.n53 VDD1.n52 9.3005
R1949 VDD1.n51 VDD1.n50 9.3005
R1950 VDD1.n20 VDD1.n19 9.3005
R1951 VDD1.n45 VDD1.n44 9.3005
R1952 VDD1.n43 VDD1.n42 9.3005
R1953 VDD1.n24 VDD1.n23 9.3005
R1954 VDD1.n37 VDD1.n36 9.3005
R1955 VDD1.n35 VDD1.n34 9.3005
R1956 VDD1.n28 VDD1.n27 9.3005
R1957 VDD1.n168 VDD1.n167 9.3005
R1958 VDD1.n87 VDD1.n86 9.3005
R1959 VDD1.n162 VDD1.n161 9.3005
R1960 VDD1.n134 VDD1.n133 9.3005
R1961 VDD1.n103 VDD1.n102 9.3005
R1962 VDD1.n128 VDD1.n127 9.3005
R1963 VDD1.n126 VDD1.n125 9.3005
R1964 VDD1.n107 VDD1.n106 9.3005
R1965 VDD1.n120 VDD1.n119 9.3005
R1966 VDD1.n118 VDD1.n117 9.3005
R1967 VDD1.n111 VDD1.n110 9.3005
R1968 VDD1.n136 VDD1.n135 9.3005
R1969 VDD1.n99 VDD1.n98 9.3005
R1970 VDD1.n142 VDD1.n141 9.3005
R1971 VDD1.n144 VDD1.n143 9.3005
R1972 VDD1.n95 VDD1.n94 9.3005
R1973 VDD1.n150 VDD1.n149 9.3005
R1974 VDD1.n152 VDD1.n151 9.3005
R1975 VDD1.n153 VDD1.n90 9.3005
R1976 VDD1.n160 VDD1.n159 9.3005
R1977 VDD1.n61 VDD1.n14 8.92171
R1978 VDD1.n46 VDD1.n45 8.92171
R1979 VDD1.n129 VDD1.n128 8.92171
R1980 VDD1.n144 VDD1.n97 8.92171
R1981 VDD1.n58 VDD1.n57 8.14595
R1982 VDD1.n49 VDD1.n20 8.14595
R1983 VDD1.n132 VDD1.n103 8.14595
R1984 VDD1.n141 VDD1.n140 8.14595
R1985 VDD1.n54 VDD1.n16 7.3702
R1986 VDD1.n50 VDD1.n18 7.3702
R1987 VDD1.n133 VDD1.n101 7.3702
R1988 VDD1.n137 VDD1.n99 7.3702
R1989 VDD1.n54 VDD1.n53 6.59444
R1990 VDD1.n53 VDD1.n18 6.59444
R1991 VDD1.n136 VDD1.n101 6.59444
R1992 VDD1.n137 VDD1.n136 6.59444
R1993 VDD1.n57 VDD1.n16 5.81868
R1994 VDD1.n50 VDD1.n49 5.81868
R1995 VDD1.n133 VDD1.n132 5.81868
R1996 VDD1.n140 VDD1.n99 5.81868
R1997 VDD1.n58 VDD1.n14 5.04292
R1998 VDD1.n46 VDD1.n20 5.04292
R1999 VDD1.n129 VDD1.n103 5.04292
R2000 VDD1.n141 VDD1.n97 5.04292
R2001 VDD1.n62 VDD1.n61 4.26717
R2002 VDD1.n45 VDD1.n22 4.26717
R2003 VDD1.n128 VDD1.n105 4.26717
R2004 VDD1.n145 VDD1.n144 4.26717
R2005 VDD1.n29 VDD1.n27 3.70982
R2006 VDD1.n112 VDD1.n110 3.70982
R2007 VDD1.n65 VDD1.n12 3.49141
R2008 VDD1.n42 VDD1.n41 3.49141
R2009 VDD1.n125 VDD1.n124 3.49141
R2010 VDD1.n148 VDD1.n95 3.49141
R2011 VDD1.n84 VDD1.n0 2.71565
R2012 VDD1.n66 VDD1.n10 2.71565
R2013 VDD1.n38 VDD1.n24 2.71565
R2014 VDD1.n121 VDD1.n107 2.71565
R2015 VDD1.n149 VDD1.n93 2.71565
R2016 VDD1.n169 VDD1.n85 2.71565
R2017 VDD1.n82 VDD1.n81 1.93989
R2018 VDD1.n70 VDD1.n69 1.93989
R2019 VDD1.n37 VDD1.n26 1.93989
R2020 VDD1.n120 VDD1.n109 1.93989
R2021 VDD1.n154 VDD1.n152 1.93989
R2022 VDD1.n167 VDD1.n166 1.93989
R2023 VDD1.n78 VDD1.n2 1.16414
R2024 VDD1.n73 VDD1.n7 1.16414
R2025 VDD1.n34 VDD1.n33 1.16414
R2026 VDD1.n117 VDD1.n116 1.16414
R2027 VDD1.n153 VDD1.n91 1.16414
R2028 VDD1.n163 VDD1.n87 1.16414
R2029 VDD1.n77 VDD1.n4 0.388379
R2030 VDD1.n74 VDD1.n6 0.388379
R2031 VDD1.n30 VDD1.n28 0.388379
R2032 VDD1.n113 VDD1.n111 0.388379
R2033 VDD1.n159 VDD1.n158 0.388379
R2034 VDD1.n162 VDD1.n89 0.388379
R2035 VDD1.n83 VDD1.n1 0.155672
R2036 VDD1.n76 VDD1.n1 0.155672
R2037 VDD1.n76 VDD1.n75 0.155672
R2038 VDD1.n75 VDD1.n5 0.155672
R2039 VDD1.n68 VDD1.n5 0.155672
R2040 VDD1.n68 VDD1.n67 0.155672
R2041 VDD1.n67 VDD1.n11 0.155672
R2042 VDD1.n60 VDD1.n11 0.155672
R2043 VDD1.n60 VDD1.n59 0.155672
R2044 VDD1.n59 VDD1.n15 0.155672
R2045 VDD1.n52 VDD1.n15 0.155672
R2046 VDD1.n52 VDD1.n51 0.155672
R2047 VDD1.n51 VDD1.n19 0.155672
R2048 VDD1.n44 VDD1.n19 0.155672
R2049 VDD1.n44 VDD1.n43 0.155672
R2050 VDD1.n43 VDD1.n23 0.155672
R2051 VDD1.n36 VDD1.n23 0.155672
R2052 VDD1.n36 VDD1.n35 0.155672
R2053 VDD1.n35 VDD1.n27 0.155672
R2054 VDD1.n118 VDD1.n110 0.155672
R2055 VDD1.n119 VDD1.n118 0.155672
R2056 VDD1.n119 VDD1.n106 0.155672
R2057 VDD1.n126 VDD1.n106 0.155672
R2058 VDD1.n127 VDD1.n126 0.155672
R2059 VDD1.n127 VDD1.n102 0.155672
R2060 VDD1.n134 VDD1.n102 0.155672
R2061 VDD1.n135 VDD1.n134 0.155672
R2062 VDD1.n135 VDD1.n98 0.155672
R2063 VDD1.n142 VDD1.n98 0.155672
R2064 VDD1.n143 VDD1.n142 0.155672
R2065 VDD1.n143 VDD1.n94 0.155672
R2066 VDD1.n150 VDD1.n94 0.155672
R2067 VDD1.n151 VDD1.n150 0.155672
R2068 VDD1.n151 VDD1.n90 0.155672
R2069 VDD1.n160 VDD1.n90 0.155672
R2070 VDD1.n161 VDD1.n160 0.155672
R2071 VDD1.n161 VDD1.n86 0.155672
R2072 VDD1.n168 VDD1.n86 0.155672
C0 B VTAIL 4.58362f
C1 w_n2306_n4036# VTAIL 3.20872f
C2 VTAIL VN 3.10535f
C3 w_n2306_n4036# B 10.1881f
C4 B VN 1.16222f
C5 w_n2306_n4036# VN 3.28121f
C6 VP VTAIL 3.11965f
C7 VDD1 VTAIL 5.99528f
C8 B VP 1.64824f
C9 w_n2306_n4036# VP 3.57583f
C10 B VDD1 2.02698f
C11 w_n2306_n4036# VDD1 2.05751f
C12 VP VN 6.26164f
C13 VDD1 VN 0.148644f
C14 VDD1 VP 3.75874f
C15 VDD2 VTAIL 6.04836f
C16 B VDD2 2.06071f
C17 w_n2306_n4036# VDD2 2.08845f
C18 VDD2 VN 3.5594f
C19 VP VDD2 0.350856f
C20 VDD1 VDD2 0.724697f
C21 VDD2 VSUBS 1.085454f
C22 VDD1 VSUBS 5.40788f
C23 VTAIL VSUBS 1.185055f
C24 VN VSUBS 8.65303f
C25 VP VSUBS 1.925865f
C26 B VSUBS 4.493237f
C27 w_n2306_n4036# VSUBS 0.114092p
C28 VDD1.n0 VSUBS 0.029376f
C29 VDD1.n1 VSUBS 0.028848f
C30 VDD1.n2 VSUBS 0.015502f
C31 VDD1.n3 VSUBS 0.036641f
C32 VDD1.n4 VSUBS 0.015958f
C33 VDD1.n5 VSUBS 0.028848f
C34 VDD1.n6 VSUBS 0.015958f
C35 VDD1.n7 VSUBS 0.015502f
C36 VDD1.n8 VSUBS 0.036641f
C37 VDD1.n9 VSUBS 0.036641f
C38 VDD1.n10 VSUBS 0.016414f
C39 VDD1.n11 VSUBS 0.028848f
C40 VDD1.n12 VSUBS 0.015502f
C41 VDD1.n13 VSUBS 0.036641f
C42 VDD1.n14 VSUBS 0.016414f
C43 VDD1.n15 VSUBS 0.028848f
C44 VDD1.n16 VSUBS 0.015502f
C45 VDD1.n17 VSUBS 0.036641f
C46 VDD1.n18 VSUBS 0.016414f
C47 VDD1.n19 VSUBS 0.028848f
C48 VDD1.n20 VSUBS 0.015502f
C49 VDD1.n21 VSUBS 0.036641f
C50 VDD1.n22 VSUBS 0.016414f
C51 VDD1.n23 VSUBS 0.028848f
C52 VDD1.n24 VSUBS 0.015502f
C53 VDD1.n25 VSUBS 0.036641f
C54 VDD1.n26 VSUBS 0.016414f
C55 VDD1.n27 VSUBS 1.88655f
C56 VDD1.n28 VSUBS 0.015502f
C57 VDD1.t0 VSUBS 0.078465f
C58 VDD1.n29 VSUBS 0.206248f
C59 VDD1.n30 VSUBS 0.023309f
C60 VDD1.n31 VSUBS 0.02748f
C61 VDD1.n32 VSUBS 0.036641f
C62 VDD1.n33 VSUBS 0.016414f
C63 VDD1.n34 VSUBS 0.015502f
C64 VDD1.n35 VSUBS 0.028848f
C65 VDD1.n36 VSUBS 0.028848f
C66 VDD1.n37 VSUBS 0.015502f
C67 VDD1.n38 VSUBS 0.016414f
C68 VDD1.n39 VSUBS 0.036641f
C69 VDD1.n40 VSUBS 0.036641f
C70 VDD1.n41 VSUBS 0.016414f
C71 VDD1.n42 VSUBS 0.015502f
C72 VDD1.n43 VSUBS 0.028848f
C73 VDD1.n44 VSUBS 0.028848f
C74 VDD1.n45 VSUBS 0.015502f
C75 VDD1.n46 VSUBS 0.016414f
C76 VDD1.n47 VSUBS 0.036641f
C77 VDD1.n48 VSUBS 0.036641f
C78 VDD1.n49 VSUBS 0.016414f
C79 VDD1.n50 VSUBS 0.015502f
C80 VDD1.n51 VSUBS 0.028848f
C81 VDD1.n52 VSUBS 0.028848f
C82 VDD1.n53 VSUBS 0.015502f
C83 VDD1.n54 VSUBS 0.016414f
C84 VDD1.n55 VSUBS 0.036641f
C85 VDD1.n56 VSUBS 0.036641f
C86 VDD1.n57 VSUBS 0.016414f
C87 VDD1.n58 VSUBS 0.015502f
C88 VDD1.n59 VSUBS 0.028848f
C89 VDD1.n60 VSUBS 0.028848f
C90 VDD1.n61 VSUBS 0.015502f
C91 VDD1.n62 VSUBS 0.016414f
C92 VDD1.n63 VSUBS 0.036641f
C93 VDD1.n64 VSUBS 0.036641f
C94 VDD1.n65 VSUBS 0.016414f
C95 VDD1.n66 VSUBS 0.015502f
C96 VDD1.n67 VSUBS 0.028848f
C97 VDD1.n68 VSUBS 0.028848f
C98 VDD1.n69 VSUBS 0.015502f
C99 VDD1.n70 VSUBS 0.016414f
C100 VDD1.n71 VSUBS 0.036641f
C101 VDD1.n72 VSUBS 0.036641f
C102 VDD1.n73 VSUBS 0.016414f
C103 VDD1.n74 VSUBS 0.015502f
C104 VDD1.n75 VSUBS 0.028848f
C105 VDD1.n76 VSUBS 0.028848f
C106 VDD1.n77 VSUBS 0.015502f
C107 VDD1.n78 VSUBS 0.016414f
C108 VDD1.n79 VSUBS 0.036641f
C109 VDD1.n80 VSUBS 0.080794f
C110 VDD1.n81 VSUBS 0.016414f
C111 VDD1.n82 VSUBS 0.015502f
C112 VDD1.n83 VSUBS 0.065893f
C113 VDD1.n84 VSUBS 0.062193f
C114 VDD1.n85 VSUBS 0.029376f
C115 VDD1.n86 VSUBS 0.028848f
C116 VDD1.n87 VSUBS 0.015502f
C117 VDD1.n88 VSUBS 0.036641f
C118 VDD1.n89 VSUBS 0.015958f
C119 VDD1.n90 VSUBS 0.028848f
C120 VDD1.n91 VSUBS 0.016414f
C121 VDD1.n92 VSUBS 0.036641f
C122 VDD1.n93 VSUBS 0.016414f
C123 VDD1.n94 VSUBS 0.028848f
C124 VDD1.n95 VSUBS 0.015502f
C125 VDD1.n96 VSUBS 0.036641f
C126 VDD1.n97 VSUBS 0.016414f
C127 VDD1.n98 VSUBS 0.028848f
C128 VDD1.n99 VSUBS 0.015502f
C129 VDD1.n100 VSUBS 0.036641f
C130 VDD1.n101 VSUBS 0.016414f
C131 VDD1.n102 VSUBS 0.028848f
C132 VDD1.n103 VSUBS 0.015502f
C133 VDD1.n104 VSUBS 0.036641f
C134 VDD1.n105 VSUBS 0.016414f
C135 VDD1.n106 VSUBS 0.028848f
C136 VDD1.n107 VSUBS 0.015502f
C137 VDD1.n108 VSUBS 0.036641f
C138 VDD1.n109 VSUBS 0.016414f
C139 VDD1.n110 VSUBS 1.88655f
C140 VDD1.n111 VSUBS 0.015502f
C141 VDD1.t1 VSUBS 0.078465f
C142 VDD1.n112 VSUBS 0.206248f
C143 VDD1.n113 VSUBS 0.023309f
C144 VDD1.n114 VSUBS 0.02748f
C145 VDD1.n115 VSUBS 0.036641f
C146 VDD1.n116 VSUBS 0.016414f
C147 VDD1.n117 VSUBS 0.015502f
C148 VDD1.n118 VSUBS 0.028848f
C149 VDD1.n119 VSUBS 0.028848f
C150 VDD1.n120 VSUBS 0.015502f
C151 VDD1.n121 VSUBS 0.016414f
C152 VDD1.n122 VSUBS 0.036641f
C153 VDD1.n123 VSUBS 0.036641f
C154 VDD1.n124 VSUBS 0.016414f
C155 VDD1.n125 VSUBS 0.015502f
C156 VDD1.n126 VSUBS 0.028848f
C157 VDD1.n127 VSUBS 0.028848f
C158 VDD1.n128 VSUBS 0.015502f
C159 VDD1.n129 VSUBS 0.016414f
C160 VDD1.n130 VSUBS 0.036641f
C161 VDD1.n131 VSUBS 0.036641f
C162 VDD1.n132 VSUBS 0.016414f
C163 VDD1.n133 VSUBS 0.015502f
C164 VDD1.n134 VSUBS 0.028848f
C165 VDD1.n135 VSUBS 0.028848f
C166 VDD1.n136 VSUBS 0.015502f
C167 VDD1.n137 VSUBS 0.016414f
C168 VDD1.n138 VSUBS 0.036641f
C169 VDD1.n139 VSUBS 0.036641f
C170 VDD1.n140 VSUBS 0.016414f
C171 VDD1.n141 VSUBS 0.015502f
C172 VDD1.n142 VSUBS 0.028848f
C173 VDD1.n143 VSUBS 0.028848f
C174 VDD1.n144 VSUBS 0.015502f
C175 VDD1.n145 VSUBS 0.016414f
C176 VDD1.n146 VSUBS 0.036641f
C177 VDD1.n147 VSUBS 0.036641f
C178 VDD1.n148 VSUBS 0.016414f
C179 VDD1.n149 VSUBS 0.015502f
C180 VDD1.n150 VSUBS 0.028848f
C181 VDD1.n151 VSUBS 0.028848f
C182 VDD1.n152 VSUBS 0.015502f
C183 VDD1.n153 VSUBS 0.015502f
C184 VDD1.n154 VSUBS 0.016414f
C185 VDD1.n155 VSUBS 0.036641f
C186 VDD1.n156 VSUBS 0.036641f
C187 VDD1.n157 VSUBS 0.036641f
C188 VDD1.n158 VSUBS 0.015958f
C189 VDD1.n159 VSUBS 0.015502f
C190 VDD1.n160 VSUBS 0.028848f
C191 VDD1.n161 VSUBS 0.028848f
C192 VDD1.n162 VSUBS 0.015502f
C193 VDD1.n163 VSUBS 0.016414f
C194 VDD1.n164 VSUBS 0.036641f
C195 VDD1.n165 VSUBS 0.080794f
C196 VDD1.n166 VSUBS 0.016414f
C197 VDD1.n167 VSUBS 0.015502f
C198 VDD1.n168 VSUBS 0.065893f
C199 VDD1.n169 VSUBS 1.08583f
C200 VP.t0 VSUBS 4.96983f
C201 VP.t1 VSUBS 5.74703f
C202 VP.n0 VSUBS 5.97661f
C203 B.n0 VSUBS 0.006146f
C204 B.n1 VSUBS 0.006146f
C205 B.n2 VSUBS 0.00909f
C206 B.n3 VSUBS 0.006966f
C207 B.n4 VSUBS 0.006966f
C208 B.n5 VSUBS 0.006966f
C209 B.n6 VSUBS 0.006966f
C210 B.n7 VSUBS 0.006966f
C211 B.n8 VSUBS 0.006966f
C212 B.n9 VSUBS 0.006966f
C213 B.n10 VSUBS 0.006966f
C214 B.n11 VSUBS 0.006966f
C215 B.n12 VSUBS 0.006966f
C216 B.n13 VSUBS 0.006966f
C217 B.n14 VSUBS 0.006966f
C218 B.n15 VSUBS 0.017569f
C219 B.n16 VSUBS 0.006966f
C220 B.n17 VSUBS 0.006966f
C221 B.n18 VSUBS 0.006966f
C222 B.n19 VSUBS 0.006966f
C223 B.n20 VSUBS 0.006966f
C224 B.n21 VSUBS 0.006966f
C225 B.n22 VSUBS 0.006966f
C226 B.n23 VSUBS 0.006966f
C227 B.n24 VSUBS 0.006966f
C228 B.n25 VSUBS 0.006966f
C229 B.n26 VSUBS 0.006966f
C230 B.n27 VSUBS 0.006966f
C231 B.n28 VSUBS 0.006966f
C232 B.n29 VSUBS 0.006966f
C233 B.n30 VSUBS 0.006966f
C234 B.n31 VSUBS 0.006966f
C235 B.n32 VSUBS 0.006966f
C236 B.n33 VSUBS 0.006966f
C237 B.n34 VSUBS 0.006966f
C238 B.n35 VSUBS 0.006966f
C239 B.n36 VSUBS 0.006966f
C240 B.n37 VSUBS 0.006966f
C241 B.n38 VSUBS 0.006966f
C242 B.n39 VSUBS 0.006966f
C243 B.n40 VSUBS 0.006966f
C244 B.n41 VSUBS 0.006966f
C245 B.t10 VSUBS 0.285988f
C246 B.t11 VSUBS 0.323079f
C247 B.t9 VSUBS 2.08157f
C248 B.n42 VSUBS 0.508061f
C249 B.n43 VSUBS 0.296453f
C250 B.n44 VSUBS 0.006966f
C251 B.n45 VSUBS 0.006966f
C252 B.n46 VSUBS 0.006966f
C253 B.n47 VSUBS 0.006966f
C254 B.t7 VSUBS 0.285992f
C255 B.t8 VSUBS 0.323082f
C256 B.t6 VSUBS 2.08157f
C257 B.n48 VSUBS 0.508058f
C258 B.n49 VSUBS 0.29645f
C259 B.n50 VSUBS 0.016139f
C260 B.n51 VSUBS 0.006966f
C261 B.n52 VSUBS 0.006966f
C262 B.n53 VSUBS 0.006966f
C263 B.n54 VSUBS 0.006966f
C264 B.n55 VSUBS 0.006966f
C265 B.n56 VSUBS 0.006966f
C266 B.n57 VSUBS 0.006966f
C267 B.n58 VSUBS 0.006966f
C268 B.n59 VSUBS 0.006966f
C269 B.n60 VSUBS 0.006966f
C270 B.n61 VSUBS 0.006966f
C271 B.n62 VSUBS 0.006966f
C272 B.n63 VSUBS 0.006966f
C273 B.n64 VSUBS 0.006966f
C274 B.n65 VSUBS 0.006966f
C275 B.n66 VSUBS 0.006966f
C276 B.n67 VSUBS 0.006966f
C277 B.n68 VSUBS 0.006966f
C278 B.n69 VSUBS 0.006966f
C279 B.n70 VSUBS 0.006966f
C280 B.n71 VSUBS 0.006966f
C281 B.n72 VSUBS 0.006966f
C282 B.n73 VSUBS 0.006966f
C283 B.n74 VSUBS 0.006966f
C284 B.n75 VSUBS 0.006966f
C285 B.n76 VSUBS 0.017569f
C286 B.n77 VSUBS 0.006966f
C287 B.n78 VSUBS 0.006966f
C288 B.n79 VSUBS 0.006966f
C289 B.n80 VSUBS 0.006966f
C290 B.n81 VSUBS 0.006966f
C291 B.n82 VSUBS 0.006966f
C292 B.n83 VSUBS 0.006966f
C293 B.n84 VSUBS 0.006966f
C294 B.n85 VSUBS 0.006966f
C295 B.n86 VSUBS 0.006966f
C296 B.n87 VSUBS 0.006966f
C297 B.n88 VSUBS 0.006966f
C298 B.n89 VSUBS 0.006966f
C299 B.n90 VSUBS 0.006966f
C300 B.n91 VSUBS 0.006966f
C301 B.n92 VSUBS 0.006966f
C302 B.n93 VSUBS 0.006966f
C303 B.n94 VSUBS 0.006966f
C304 B.n95 VSUBS 0.006966f
C305 B.n96 VSUBS 0.006966f
C306 B.n97 VSUBS 0.006966f
C307 B.n98 VSUBS 0.006966f
C308 B.n99 VSUBS 0.006966f
C309 B.n100 VSUBS 0.006966f
C310 B.n101 VSUBS 0.006966f
C311 B.n102 VSUBS 0.006966f
C312 B.n103 VSUBS 0.006966f
C313 B.n104 VSUBS 0.017569f
C314 B.n105 VSUBS 0.006966f
C315 B.n106 VSUBS 0.006966f
C316 B.n107 VSUBS 0.006966f
C317 B.n108 VSUBS 0.006966f
C318 B.n109 VSUBS 0.006966f
C319 B.n110 VSUBS 0.006966f
C320 B.n111 VSUBS 0.006966f
C321 B.n112 VSUBS 0.006966f
C322 B.n113 VSUBS 0.006966f
C323 B.n114 VSUBS 0.006966f
C324 B.n115 VSUBS 0.006966f
C325 B.n116 VSUBS 0.006966f
C326 B.n117 VSUBS 0.006966f
C327 B.n118 VSUBS 0.006966f
C328 B.n119 VSUBS 0.006966f
C329 B.n120 VSUBS 0.006966f
C330 B.n121 VSUBS 0.006966f
C331 B.n122 VSUBS 0.006966f
C332 B.n123 VSUBS 0.006966f
C333 B.n124 VSUBS 0.006966f
C334 B.n125 VSUBS 0.006966f
C335 B.n126 VSUBS 0.006966f
C336 B.n127 VSUBS 0.006966f
C337 B.n128 VSUBS 0.006966f
C338 B.n129 VSUBS 0.006966f
C339 B.t2 VSUBS 0.285992f
C340 B.t1 VSUBS 0.323082f
C341 B.t0 VSUBS 2.08157f
C342 B.n130 VSUBS 0.508058f
C343 B.n131 VSUBS 0.29645f
C344 B.n132 VSUBS 0.006966f
C345 B.n133 VSUBS 0.006966f
C346 B.n134 VSUBS 0.006966f
C347 B.n135 VSUBS 0.006966f
C348 B.n136 VSUBS 0.003893f
C349 B.n137 VSUBS 0.006966f
C350 B.n138 VSUBS 0.006966f
C351 B.n139 VSUBS 0.006966f
C352 B.n140 VSUBS 0.006966f
C353 B.n141 VSUBS 0.006966f
C354 B.n142 VSUBS 0.006966f
C355 B.n143 VSUBS 0.006966f
C356 B.n144 VSUBS 0.006966f
C357 B.n145 VSUBS 0.006966f
C358 B.n146 VSUBS 0.006966f
C359 B.n147 VSUBS 0.006966f
C360 B.n148 VSUBS 0.006966f
C361 B.n149 VSUBS 0.006966f
C362 B.n150 VSUBS 0.006966f
C363 B.n151 VSUBS 0.006966f
C364 B.n152 VSUBS 0.006966f
C365 B.n153 VSUBS 0.006966f
C366 B.n154 VSUBS 0.006966f
C367 B.n155 VSUBS 0.006966f
C368 B.n156 VSUBS 0.006966f
C369 B.n157 VSUBS 0.006966f
C370 B.n158 VSUBS 0.006966f
C371 B.n159 VSUBS 0.006966f
C372 B.n160 VSUBS 0.006966f
C373 B.n161 VSUBS 0.006966f
C374 B.n162 VSUBS 0.017569f
C375 B.n163 VSUBS 0.006966f
C376 B.n164 VSUBS 0.006966f
C377 B.n165 VSUBS 0.006966f
C378 B.n166 VSUBS 0.006966f
C379 B.n167 VSUBS 0.006966f
C380 B.n168 VSUBS 0.006966f
C381 B.n169 VSUBS 0.006966f
C382 B.n170 VSUBS 0.006966f
C383 B.n171 VSUBS 0.006966f
C384 B.n172 VSUBS 0.006966f
C385 B.n173 VSUBS 0.006966f
C386 B.n174 VSUBS 0.006966f
C387 B.n175 VSUBS 0.006966f
C388 B.n176 VSUBS 0.006966f
C389 B.n177 VSUBS 0.006966f
C390 B.n178 VSUBS 0.006966f
C391 B.n179 VSUBS 0.006966f
C392 B.n180 VSUBS 0.006966f
C393 B.n181 VSUBS 0.006966f
C394 B.n182 VSUBS 0.006966f
C395 B.n183 VSUBS 0.006966f
C396 B.n184 VSUBS 0.006966f
C397 B.n185 VSUBS 0.006966f
C398 B.n186 VSUBS 0.006966f
C399 B.n187 VSUBS 0.006966f
C400 B.n188 VSUBS 0.006966f
C401 B.n189 VSUBS 0.006966f
C402 B.n190 VSUBS 0.006966f
C403 B.n191 VSUBS 0.006966f
C404 B.n192 VSUBS 0.006966f
C405 B.n193 VSUBS 0.006966f
C406 B.n194 VSUBS 0.006966f
C407 B.n195 VSUBS 0.006966f
C408 B.n196 VSUBS 0.006966f
C409 B.n197 VSUBS 0.006966f
C410 B.n198 VSUBS 0.006966f
C411 B.n199 VSUBS 0.006966f
C412 B.n200 VSUBS 0.006966f
C413 B.n201 VSUBS 0.006966f
C414 B.n202 VSUBS 0.006966f
C415 B.n203 VSUBS 0.006966f
C416 B.n204 VSUBS 0.006966f
C417 B.n205 VSUBS 0.006966f
C418 B.n206 VSUBS 0.006966f
C419 B.n207 VSUBS 0.006966f
C420 B.n208 VSUBS 0.006966f
C421 B.n209 VSUBS 0.006966f
C422 B.n210 VSUBS 0.006966f
C423 B.n211 VSUBS 0.006966f
C424 B.n212 VSUBS 0.006966f
C425 B.n213 VSUBS 0.017569f
C426 B.n214 VSUBS 0.018284f
C427 B.n215 VSUBS 0.018284f
C428 B.n216 VSUBS 0.006966f
C429 B.n217 VSUBS 0.006966f
C430 B.n218 VSUBS 0.006966f
C431 B.n219 VSUBS 0.006966f
C432 B.n220 VSUBS 0.006966f
C433 B.n221 VSUBS 0.006966f
C434 B.n222 VSUBS 0.006966f
C435 B.n223 VSUBS 0.006966f
C436 B.n224 VSUBS 0.006966f
C437 B.n225 VSUBS 0.006966f
C438 B.n226 VSUBS 0.006966f
C439 B.n227 VSUBS 0.006966f
C440 B.n228 VSUBS 0.006966f
C441 B.n229 VSUBS 0.006966f
C442 B.n230 VSUBS 0.006966f
C443 B.n231 VSUBS 0.006966f
C444 B.n232 VSUBS 0.006966f
C445 B.n233 VSUBS 0.006966f
C446 B.n234 VSUBS 0.006966f
C447 B.n235 VSUBS 0.006966f
C448 B.n236 VSUBS 0.006966f
C449 B.n237 VSUBS 0.006966f
C450 B.n238 VSUBS 0.006966f
C451 B.n239 VSUBS 0.006966f
C452 B.n240 VSUBS 0.006966f
C453 B.n241 VSUBS 0.006966f
C454 B.n242 VSUBS 0.006966f
C455 B.n243 VSUBS 0.006966f
C456 B.n244 VSUBS 0.006966f
C457 B.n245 VSUBS 0.006966f
C458 B.n246 VSUBS 0.006966f
C459 B.n247 VSUBS 0.006966f
C460 B.n248 VSUBS 0.006966f
C461 B.n249 VSUBS 0.006966f
C462 B.n250 VSUBS 0.006966f
C463 B.n251 VSUBS 0.006966f
C464 B.n252 VSUBS 0.006966f
C465 B.n253 VSUBS 0.006966f
C466 B.n254 VSUBS 0.006966f
C467 B.n255 VSUBS 0.006966f
C468 B.n256 VSUBS 0.006966f
C469 B.n257 VSUBS 0.006966f
C470 B.n258 VSUBS 0.006966f
C471 B.n259 VSUBS 0.006966f
C472 B.n260 VSUBS 0.006966f
C473 B.n261 VSUBS 0.006966f
C474 B.n262 VSUBS 0.006966f
C475 B.n263 VSUBS 0.006966f
C476 B.n264 VSUBS 0.006966f
C477 B.n265 VSUBS 0.006966f
C478 B.n266 VSUBS 0.006966f
C479 B.n267 VSUBS 0.006966f
C480 B.n268 VSUBS 0.006966f
C481 B.n269 VSUBS 0.006966f
C482 B.n270 VSUBS 0.006966f
C483 B.n271 VSUBS 0.006966f
C484 B.n272 VSUBS 0.006966f
C485 B.n273 VSUBS 0.006966f
C486 B.n274 VSUBS 0.006966f
C487 B.n275 VSUBS 0.006966f
C488 B.n276 VSUBS 0.006966f
C489 B.n277 VSUBS 0.006966f
C490 B.n278 VSUBS 0.006966f
C491 B.n279 VSUBS 0.006966f
C492 B.n280 VSUBS 0.006966f
C493 B.n281 VSUBS 0.006966f
C494 B.n282 VSUBS 0.006966f
C495 B.n283 VSUBS 0.006966f
C496 B.n284 VSUBS 0.006966f
C497 B.n285 VSUBS 0.006966f
C498 B.n286 VSUBS 0.006966f
C499 B.n287 VSUBS 0.006966f
C500 B.n288 VSUBS 0.006966f
C501 B.t5 VSUBS 0.285988f
C502 B.t4 VSUBS 0.323079f
C503 B.t3 VSUBS 2.08157f
C504 B.n289 VSUBS 0.508061f
C505 B.n290 VSUBS 0.296453f
C506 B.n291 VSUBS 0.016139f
C507 B.n292 VSUBS 0.006556f
C508 B.n293 VSUBS 0.006966f
C509 B.n294 VSUBS 0.006966f
C510 B.n295 VSUBS 0.006966f
C511 B.n296 VSUBS 0.006966f
C512 B.n297 VSUBS 0.006966f
C513 B.n298 VSUBS 0.006966f
C514 B.n299 VSUBS 0.006966f
C515 B.n300 VSUBS 0.006966f
C516 B.n301 VSUBS 0.006966f
C517 B.n302 VSUBS 0.006966f
C518 B.n303 VSUBS 0.006966f
C519 B.n304 VSUBS 0.006966f
C520 B.n305 VSUBS 0.006966f
C521 B.n306 VSUBS 0.006966f
C522 B.n307 VSUBS 0.006966f
C523 B.n308 VSUBS 0.003893f
C524 B.n309 VSUBS 0.016139f
C525 B.n310 VSUBS 0.006556f
C526 B.n311 VSUBS 0.006966f
C527 B.n312 VSUBS 0.006966f
C528 B.n313 VSUBS 0.006966f
C529 B.n314 VSUBS 0.006966f
C530 B.n315 VSUBS 0.006966f
C531 B.n316 VSUBS 0.006966f
C532 B.n317 VSUBS 0.006966f
C533 B.n318 VSUBS 0.006966f
C534 B.n319 VSUBS 0.006966f
C535 B.n320 VSUBS 0.006966f
C536 B.n321 VSUBS 0.006966f
C537 B.n322 VSUBS 0.006966f
C538 B.n323 VSUBS 0.006966f
C539 B.n324 VSUBS 0.006966f
C540 B.n325 VSUBS 0.006966f
C541 B.n326 VSUBS 0.006966f
C542 B.n327 VSUBS 0.006966f
C543 B.n328 VSUBS 0.006966f
C544 B.n329 VSUBS 0.006966f
C545 B.n330 VSUBS 0.006966f
C546 B.n331 VSUBS 0.006966f
C547 B.n332 VSUBS 0.006966f
C548 B.n333 VSUBS 0.006966f
C549 B.n334 VSUBS 0.006966f
C550 B.n335 VSUBS 0.006966f
C551 B.n336 VSUBS 0.006966f
C552 B.n337 VSUBS 0.006966f
C553 B.n338 VSUBS 0.006966f
C554 B.n339 VSUBS 0.006966f
C555 B.n340 VSUBS 0.006966f
C556 B.n341 VSUBS 0.006966f
C557 B.n342 VSUBS 0.006966f
C558 B.n343 VSUBS 0.006966f
C559 B.n344 VSUBS 0.006966f
C560 B.n345 VSUBS 0.006966f
C561 B.n346 VSUBS 0.006966f
C562 B.n347 VSUBS 0.006966f
C563 B.n348 VSUBS 0.006966f
C564 B.n349 VSUBS 0.006966f
C565 B.n350 VSUBS 0.006966f
C566 B.n351 VSUBS 0.006966f
C567 B.n352 VSUBS 0.006966f
C568 B.n353 VSUBS 0.006966f
C569 B.n354 VSUBS 0.006966f
C570 B.n355 VSUBS 0.006966f
C571 B.n356 VSUBS 0.006966f
C572 B.n357 VSUBS 0.006966f
C573 B.n358 VSUBS 0.006966f
C574 B.n359 VSUBS 0.006966f
C575 B.n360 VSUBS 0.006966f
C576 B.n361 VSUBS 0.006966f
C577 B.n362 VSUBS 0.006966f
C578 B.n363 VSUBS 0.006966f
C579 B.n364 VSUBS 0.006966f
C580 B.n365 VSUBS 0.006966f
C581 B.n366 VSUBS 0.006966f
C582 B.n367 VSUBS 0.006966f
C583 B.n368 VSUBS 0.006966f
C584 B.n369 VSUBS 0.006966f
C585 B.n370 VSUBS 0.006966f
C586 B.n371 VSUBS 0.006966f
C587 B.n372 VSUBS 0.006966f
C588 B.n373 VSUBS 0.006966f
C589 B.n374 VSUBS 0.006966f
C590 B.n375 VSUBS 0.006966f
C591 B.n376 VSUBS 0.006966f
C592 B.n377 VSUBS 0.006966f
C593 B.n378 VSUBS 0.006966f
C594 B.n379 VSUBS 0.006966f
C595 B.n380 VSUBS 0.006966f
C596 B.n381 VSUBS 0.006966f
C597 B.n382 VSUBS 0.006966f
C598 B.n383 VSUBS 0.006966f
C599 B.n384 VSUBS 0.006966f
C600 B.n385 VSUBS 0.018284f
C601 B.n386 VSUBS 0.017569f
C602 B.n387 VSUBS 0.018284f
C603 B.n388 VSUBS 0.006966f
C604 B.n389 VSUBS 0.006966f
C605 B.n390 VSUBS 0.006966f
C606 B.n391 VSUBS 0.006966f
C607 B.n392 VSUBS 0.006966f
C608 B.n393 VSUBS 0.006966f
C609 B.n394 VSUBS 0.006966f
C610 B.n395 VSUBS 0.006966f
C611 B.n396 VSUBS 0.006966f
C612 B.n397 VSUBS 0.006966f
C613 B.n398 VSUBS 0.006966f
C614 B.n399 VSUBS 0.006966f
C615 B.n400 VSUBS 0.006966f
C616 B.n401 VSUBS 0.006966f
C617 B.n402 VSUBS 0.006966f
C618 B.n403 VSUBS 0.006966f
C619 B.n404 VSUBS 0.006966f
C620 B.n405 VSUBS 0.006966f
C621 B.n406 VSUBS 0.006966f
C622 B.n407 VSUBS 0.006966f
C623 B.n408 VSUBS 0.006966f
C624 B.n409 VSUBS 0.006966f
C625 B.n410 VSUBS 0.006966f
C626 B.n411 VSUBS 0.006966f
C627 B.n412 VSUBS 0.006966f
C628 B.n413 VSUBS 0.006966f
C629 B.n414 VSUBS 0.006966f
C630 B.n415 VSUBS 0.006966f
C631 B.n416 VSUBS 0.006966f
C632 B.n417 VSUBS 0.006966f
C633 B.n418 VSUBS 0.006966f
C634 B.n419 VSUBS 0.006966f
C635 B.n420 VSUBS 0.006966f
C636 B.n421 VSUBS 0.006966f
C637 B.n422 VSUBS 0.006966f
C638 B.n423 VSUBS 0.006966f
C639 B.n424 VSUBS 0.006966f
C640 B.n425 VSUBS 0.006966f
C641 B.n426 VSUBS 0.006966f
C642 B.n427 VSUBS 0.006966f
C643 B.n428 VSUBS 0.006966f
C644 B.n429 VSUBS 0.006966f
C645 B.n430 VSUBS 0.006966f
C646 B.n431 VSUBS 0.006966f
C647 B.n432 VSUBS 0.006966f
C648 B.n433 VSUBS 0.006966f
C649 B.n434 VSUBS 0.006966f
C650 B.n435 VSUBS 0.006966f
C651 B.n436 VSUBS 0.006966f
C652 B.n437 VSUBS 0.006966f
C653 B.n438 VSUBS 0.006966f
C654 B.n439 VSUBS 0.006966f
C655 B.n440 VSUBS 0.006966f
C656 B.n441 VSUBS 0.006966f
C657 B.n442 VSUBS 0.006966f
C658 B.n443 VSUBS 0.006966f
C659 B.n444 VSUBS 0.006966f
C660 B.n445 VSUBS 0.006966f
C661 B.n446 VSUBS 0.006966f
C662 B.n447 VSUBS 0.006966f
C663 B.n448 VSUBS 0.006966f
C664 B.n449 VSUBS 0.006966f
C665 B.n450 VSUBS 0.006966f
C666 B.n451 VSUBS 0.006966f
C667 B.n452 VSUBS 0.006966f
C668 B.n453 VSUBS 0.006966f
C669 B.n454 VSUBS 0.006966f
C670 B.n455 VSUBS 0.006966f
C671 B.n456 VSUBS 0.006966f
C672 B.n457 VSUBS 0.006966f
C673 B.n458 VSUBS 0.006966f
C674 B.n459 VSUBS 0.006966f
C675 B.n460 VSUBS 0.006966f
C676 B.n461 VSUBS 0.006966f
C677 B.n462 VSUBS 0.006966f
C678 B.n463 VSUBS 0.006966f
C679 B.n464 VSUBS 0.006966f
C680 B.n465 VSUBS 0.006966f
C681 B.n466 VSUBS 0.006966f
C682 B.n467 VSUBS 0.006966f
C683 B.n468 VSUBS 0.006966f
C684 B.n469 VSUBS 0.017569f
C685 B.n470 VSUBS 0.018284f
C686 B.n471 VSUBS 0.018284f
C687 B.n472 VSUBS 0.006966f
C688 B.n473 VSUBS 0.006966f
C689 B.n474 VSUBS 0.006966f
C690 B.n475 VSUBS 0.006966f
C691 B.n476 VSUBS 0.006966f
C692 B.n477 VSUBS 0.006966f
C693 B.n478 VSUBS 0.006966f
C694 B.n479 VSUBS 0.006966f
C695 B.n480 VSUBS 0.006966f
C696 B.n481 VSUBS 0.006966f
C697 B.n482 VSUBS 0.006966f
C698 B.n483 VSUBS 0.006966f
C699 B.n484 VSUBS 0.006966f
C700 B.n485 VSUBS 0.006966f
C701 B.n486 VSUBS 0.006966f
C702 B.n487 VSUBS 0.006966f
C703 B.n488 VSUBS 0.006966f
C704 B.n489 VSUBS 0.006966f
C705 B.n490 VSUBS 0.006966f
C706 B.n491 VSUBS 0.006966f
C707 B.n492 VSUBS 0.006966f
C708 B.n493 VSUBS 0.006966f
C709 B.n494 VSUBS 0.006966f
C710 B.n495 VSUBS 0.006966f
C711 B.n496 VSUBS 0.006966f
C712 B.n497 VSUBS 0.006966f
C713 B.n498 VSUBS 0.006966f
C714 B.n499 VSUBS 0.006966f
C715 B.n500 VSUBS 0.006966f
C716 B.n501 VSUBS 0.006966f
C717 B.n502 VSUBS 0.006966f
C718 B.n503 VSUBS 0.006966f
C719 B.n504 VSUBS 0.006966f
C720 B.n505 VSUBS 0.006966f
C721 B.n506 VSUBS 0.006966f
C722 B.n507 VSUBS 0.006966f
C723 B.n508 VSUBS 0.006966f
C724 B.n509 VSUBS 0.006966f
C725 B.n510 VSUBS 0.006966f
C726 B.n511 VSUBS 0.006966f
C727 B.n512 VSUBS 0.006966f
C728 B.n513 VSUBS 0.006966f
C729 B.n514 VSUBS 0.006966f
C730 B.n515 VSUBS 0.006966f
C731 B.n516 VSUBS 0.006966f
C732 B.n517 VSUBS 0.006966f
C733 B.n518 VSUBS 0.006966f
C734 B.n519 VSUBS 0.006966f
C735 B.n520 VSUBS 0.006966f
C736 B.n521 VSUBS 0.006966f
C737 B.n522 VSUBS 0.006966f
C738 B.n523 VSUBS 0.006966f
C739 B.n524 VSUBS 0.006966f
C740 B.n525 VSUBS 0.006966f
C741 B.n526 VSUBS 0.006966f
C742 B.n527 VSUBS 0.006966f
C743 B.n528 VSUBS 0.006966f
C744 B.n529 VSUBS 0.006966f
C745 B.n530 VSUBS 0.006966f
C746 B.n531 VSUBS 0.006966f
C747 B.n532 VSUBS 0.006966f
C748 B.n533 VSUBS 0.006966f
C749 B.n534 VSUBS 0.006966f
C750 B.n535 VSUBS 0.006966f
C751 B.n536 VSUBS 0.006966f
C752 B.n537 VSUBS 0.006966f
C753 B.n538 VSUBS 0.006966f
C754 B.n539 VSUBS 0.006966f
C755 B.n540 VSUBS 0.006966f
C756 B.n541 VSUBS 0.006966f
C757 B.n542 VSUBS 0.006966f
C758 B.n543 VSUBS 0.006966f
C759 B.n544 VSUBS 0.006966f
C760 B.n545 VSUBS 0.006556f
C761 B.n546 VSUBS 0.006966f
C762 B.n547 VSUBS 0.006966f
C763 B.n548 VSUBS 0.003893f
C764 B.n549 VSUBS 0.006966f
C765 B.n550 VSUBS 0.006966f
C766 B.n551 VSUBS 0.006966f
C767 B.n552 VSUBS 0.006966f
C768 B.n553 VSUBS 0.006966f
C769 B.n554 VSUBS 0.006966f
C770 B.n555 VSUBS 0.006966f
C771 B.n556 VSUBS 0.006966f
C772 B.n557 VSUBS 0.006966f
C773 B.n558 VSUBS 0.006966f
C774 B.n559 VSUBS 0.006966f
C775 B.n560 VSUBS 0.006966f
C776 B.n561 VSUBS 0.003893f
C777 B.n562 VSUBS 0.016139f
C778 B.n563 VSUBS 0.006556f
C779 B.n564 VSUBS 0.006966f
C780 B.n565 VSUBS 0.006966f
C781 B.n566 VSUBS 0.006966f
C782 B.n567 VSUBS 0.006966f
C783 B.n568 VSUBS 0.006966f
C784 B.n569 VSUBS 0.006966f
C785 B.n570 VSUBS 0.006966f
C786 B.n571 VSUBS 0.006966f
C787 B.n572 VSUBS 0.006966f
C788 B.n573 VSUBS 0.006966f
C789 B.n574 VSUBS 0.006966f
C790 B.n575 VSUBS 0.006966f
C791 B.n576 VSUBS 0.006966f
C792 B.n577 VSUBS 0.006966f
C793 B.n578 VSUBS 0.006966f
C794 B.n579 VSUBS 0.006966f
C795 B.n580 VSUBS 0.006966f
C796 B.n581 VSUBS 0.006966f
C797 B.n582 VSUBS 0.006966f
C798 B.n583 VSUBS 0.006966f
C799 B.n584 VSUBS 0.006966f
C800 B.n585 VSUBS 0.006966f
C801 B.n586 VSUBS 0.006966f
C802 B.n587 VSUBS 0.006966f
C803 B.n588 VSUBS 0.006966f
C804 B.n589 VSUBS 0.006966f
C805 B.n590 VSUBS 0.006966f
C806 B.n591 VSUBS 0.006966f
C807 B.n592 VSUBS 0.006966f
C808 B.n593 VSUBS 0.006966f
C809 B.n594 VSUBS 0.006966f
C810 B.n595 VSUBS 0.006966f
C811 B.n596 VSUBS 0.006966f
C812 B.n597 VSUBS 0.006966f
C813 B.n598 VSUBS 0.006966f
C814 B.n599 VSUBS 0.006966f
C815 B.n600 VSUBS 0.006966f
C816 B.n601 VSUBS 0.006966f
C817 B.n602 VSUBS 0.006966f
C818 B.n603 VSUBS 0.006966f
C819 B.n604 VSUBS 0.006966f
C820 B.n605 VSUBS 0.006966f
C821 B.n606 VSUBS 0.006966f
C822 B.n607 VSUBS 0.006966f
C823 B.n608 VSUBS 0.006966f
C824 B.n609 VSUBS 0.006966f
C825 B.n610 VSUBS 0.006966f
C826 B.n611 VSUBS 0.006966f
C827 B.n612 VSUBS 0.006966f
C828 B.n613 VSUBS 0.006966f
C829 B.n614 VSUBS 0.006966f
C830 B.n615 VSUBS 0.006966f
C831 B.n616 VSUBS 0.006966f
C832 B.n617 VSUBS 0.006966f
C833 B.n618 VSUBS 0.006966f
C834 B.n619 VSUBS 0.006966f
C835 B.n620 VSUBS 0.006966f
C836 B.n621 VSUBS 0.006966f
C837 B.n622 VSUBS 0.006966f
C838 B.n623 VSUBS 0.006966f
C839 B.n624 VSUBS 0.006966f
C840 B.n625 VSUBS 0.006966f
C841 B.n626 VSUBS 0.006966f
C842 B.n627 VSUBS 0.006966f
C843 B.n628 VSUBS 0.006966f
C844 B.n629 VSUBS 0.006966f
C845 B.n630 VSUBS 0.006966f
C846 B.n631 VSUBS 0.006966f
C847 B.n632 VSUBS 0.006966f
C848 B.n633 VSUBS 0.006966f
C849 B.n634 VSUBS 0.006966f
C850 B.n635 VSUBS 0.006966f
C851 B.n636 VSUBS 0.006966f
C852 B.n637 VSUBS 0.006966f
C853 B.n638 VSUBS 0.018284f
C854 B.n639 VSUBS 0.018284f
C855 B.n640 VSUBS 0.017569f
C856 B.n641 VSUBS 0.006966f
C857 B.n642 VSUBS 0.006966f
C858 B.n643 VSUBS 0.006966f
C859 B.n644 VSUBS 0.006966f
C860 B.n645 VSUBS 0.006966f
C861 B.n646 VSUBS 0.006966f
C862 B.n647 VSUBS 0.006966f
C863 B.n648 VSUBS 0.006966f
C864 B.n649 VSUBS 0.006966f
C865 B.n650 VSUBS 0.006966f
C866 B.n651 VSUBS 0.006966f
C867 B.n652 VSUBS 0.006966f
C868 B.n653 VSUBS 0.006966f
C869 B.n654 VSUBS 0.006966f
C870 B.n655 VSUBS 0.006966f
C871 B.n656 VSUBS 0.006966f
C872 B.n657 VSUBS 0.006966f
C873 B.n658 VSUBS 0.006966f
C874 B.n659 VSUBS 0.006966f
C875 B.n660 VSUBS 0.006966f
C876 B.n661 VSUBS 0.006966f
C877 B.n662 VSUBS 0.006966f
C878 B.n663 VSUBS 0.006966f
C879 B.n664 VSUBS 0.006966f
C880 B.n665 VSUBS 0.006966f
C881 B.n666 VSUBS 0.006966f
C882 B.n667 VSUBS 0.006966f
C883 B.n668 VSUBS 0.006966f
C884 B.n669 VSUBS 0.006966f
C885 B.n670 VSUBS 0.006966f
C886 B.n671 VSUBS 0.006966f
C887 B.n672 VSUBS 0.006966f
C888 B.n673 VSUBS 0.006966f
C889 B.n674 VSUBS 0.006966f
C890 B.n675 VSUBS 0.006966f
C891 B.n676 VSUBS 0.006966f
C892 B.n677 VSUBS 0.006966f
C893 B.n678 VSUBS 0.006966f
C894 B.n679 VSUBS 0.00909f
C895 B.n680 VSUBS 0.009683f
C896 B.n681 VSUBS 0.019255f
C897 VDD2.n0 VSUBS 0.02939f
C898 VDD2.n1 VSUBS 0.028862f
C899 VDD2.n2 VSUBS 0.015509f
C900 VDD2.n3 VSUBS 0.036658f
C901 VDD2.n4 VSUBS 0.015965f
C902 VDD2.n5 VSUBS 0.028862f
C903 VDD2.n6 VSUBS 0.016421f
C904 VDD2.n7 VSUBS 0.036658f
C905 VDD2.n8 VSUBS 0.016421f
C906 VDD2.n9 VSUBS 0.028862f
C907 VDD2.n10 VSUBS 0.015509f
C908 VDD2.n11 VSUBS 0.036658f
C909 VDD2.n12 VSUBS 0.016421f
C910 VDD2.n13 VSUBS 0.028862f
C911 VDD2.n14 VSUBS 0.015509f
C912 VDD2.n15 VSUBS 0.036658f
C913 VDD2.n16 VSUBS 0.016421f
C914 VDD2.n17 VSUBS 0.028862f
C915 VDD2.n18 VSUBS 0.015509f
C916 VDD2.n19 VSUBS 0.036658f
C917 VDD2.n20 VSUBS 0.016421f
C918 VDD2.n21 VSUBS 0.028862f
C919 VDD2.n22 VSUBS 0.015509f
C920 VDD2.n23 VSUBS 0.036658f
C921 VDD2.n24 VSUBS 0.016421f
C922 VDD2.n25 VSUBS 1.88744f
C923 VDD2.n26 VSUBS 0.015509f
C924 VDD2.t0 VSUBS 0.078502f
C925 VDD2.n27 VSUBS 0.206346f
C926 VDD2.n28 VSUBS 0.02332f
C927 VDD2.n29 VSUBS 0.027493f
C928 VDD2.n30 VSUBS 0.036658f
C929 VDD2.n31 VSUBS 0.016421f
C930 VDD2.n32 VSUBS 0.015509f
C931 VDD2.n33 VSUBS 0.028862f
C932 VDD2.n34 VSUBS 0.028862f
C933 VDD2.n35 VSUBS 0.015509f
C934 VDD2.n36 VSUBS 0.016421f
C935 VDD2.n37 VSUBS 0.036658f
C936 VDD2.n38 VSUBS 0.036658f
C937 VDD2.n39 VSUBS 0.016421f
C938 VDD2.n40 VSUBS 0.015509f
C939 VDD2.n41 VSUBS 0.028862f
C940 VDD2.n42 VSUBS 0.028862f
C941 VDD2.n43 VSUBS 0.015509f
C942 VDD2.n44 VSUBS 0.016421f
C943 VDD2.n45 VSUBS 0.036658f
C944 VDD2.n46 VSUBS 0.036658f
C945 VDD2.n47 VSUBS 0.016421f
C946 VDD2.n48 VSUBS 0.015509f
C947 VDD2.n49 VSUBS 0.028862f
C948 VDD2.n50 VSUBS 0.028862f
C949 VDD2.n51 VSUBS 0.015509f
C950 VDD2.n52 VSUBS 0.016421f
C951 VDD2.n53 VSUBS 0.036658f
C952 VDD2.n54 VSUBS 0.036658f
C953 VDD2.n55 VSUBS 0.016421f
C954 VDD2.n56 VSUBS 0.015509f
C955 VDD2.n57 VSUBS 0.028862f
C956 VDD2.n58 VSUBS 0.028862f
C957 VDD2.n59 VSUBS 0.015509f
C958 VDD2.n60 VSUBS 0.016421f
C959 VDD2.n61 VSUBS 0.036658f
C960 VDD2.n62 VSUBS 0.036658f
C961 VDD2.n63 VSUBS 0.016421f
C962 VDD2.n64 VSUBS 0.015509f
C963 VDD2.n65 VSUBS 0.028862f
C964 VDD2.n66 VSUBS 0.028862f
C965 VDD2.n67 VSUBS 0.015509f
C966 VDD2.n68 VSUBS 0.015509f
C967 VDD2.n69 VSUBS 0.016421f
C968 VDD2.n70 VSUBS 0.036658f
C969 VDD2.n71 VSUBS 0.036658f
C970 VDD2.n72 VSUBS 0.036658f
C971 VDD2.n73 VSUBS 0.015965f
C972 VDD2.n74 VSUBS 0.015509f
C973 VDD2.n75 VSUBS 0.028862f
C974 VDD2.n76 VSUBS 0.028862f
C975 VDD2.n77 VSUBS 0.015509f
C976 VDD2.n78 VSUBS 0.016421f
C977 VDD2.n79 VSUBS 0.036658f
C978 VDD2.n80 VSUBS 0.080833f
C979 VDD2.n81 VSUBS 0.016421f
C980 VDD2.n82 VSUBS 0.015509f
C981 VDD2.n83 VSUBS 0.065925f
C982 VDD2.n84 VSUBS 1.02194f
C983 VDD2.n85 VSUBS 0.02939f
C984 VDD2.n86 VSUBS 0.028862f
C985 VDD2.n87 VSUBS 0.015509f
C986 VDD2.n88 VSUBS 0.036658f
C987 VDD2.n89 VSUBS 0.015965f
C988 VDD2.n90 VSUBS 0.028862f
C989 VDD2.n91 VSUBS 0.015965f
C990 VDD2.n92 VSUBS 0.015509f
C991 VDD2.n93 VSUBS 0.036658f
C992 VDD2.n94 VSUBS 0.036658f
C993 VDD2.n95 VSUBS 0.016421f
C994 VDD2.n96 VSUBS 0.028862f
C995 VDD2.n97 VSUBS 0.015509f
C996 VDD2.n98 VSUBS 0.036658f
C997 VDD2.n99 VSUBS 0.016421f
C998 VDD2.n100 VSUBS 0.028862f
C999 VDD2.n101 VSUBS 0.015509f
C1000 VDD2.n102 VSUBS 0.036658f
C1001 VDD2.n103 VSUBS 0.016421f
C1002 VDD2.n104 VSUBS 0.028862f
C1003 VDD2.n105 VSUBS 0.015509f
C1004 VDD2.n106 VSUBS 0.036658f
C1005 VDD2.n107 VSUBS 0.016421f
C1006 VDD2.n108 VSUBS 0.028862f
C1007 VDD2.n109 VSUBS 0.015509f
C1008 VDD2.n110 VSUBS 0.036658f
C1009 VDD2.n111 VSUBS 0.016421f
C1010 VDD2.n112 VSUBS 1.88744f
C1011 VDD2.n113 VSUBS 0.015509f
C1012 VDD2.t1 VSUBS 0.078502f
C1013 VDD2.n114 VSUBS 0.206346f
C1014 VDD2.n115 VSUBS 0.02332f
C1015 VDD2.n116 VSUBS 0.027493f
C1016 VDD2.n117 VSUBS 0.036658f
C1017 VDD2.n118 VSUBS 0.016421f
C1018 VDD2.n119 VSUBS 0.015509f
C1019 VDD2.n120 VSUBS 0.028862f
C1020 VDD2.n121 VSUBS 0.028862f
C1021 VDD2.n122 VSUBS 0.015509f
C1022 VDD2.n123 VSUBS 0.016421f
C1023 VDD2.n124 VSUBS 0.036658f
C1024 VDD2.n125 VSUBS 0.036658f
C1025 VDD2.n126 VSUBS 0.016421f
C1026 VDD2.n127 VSUBS 0.015509f
C1027 VDD2.n128 VSUBS 0.028862f
C1028 VDD2.n129 VSUBS 0.028862f
C1029 VDD2.n130 VSUBS 0.015509f
C1030 VDD2.n131 VSUBS 0.016421f
C1031 VDD2.n132 VSUBS 0.036658f
C1032 VDD2.n133 VSUBS 0.036658f
C1033 VDD2.n134 VSUBS 0.016421f
C1034 VDD2.n135 VSUBS 0.015509f
C1035 VDD2.n136 VSUBS 0.028862f
C1036 VDD2.n137 VSUBS 0.028862f
C1037 VDD2.n138 VSUBS 0.015509f
C1038 VDD2.n139 VSUBS 0.016421f
C1039 VDD2.n140 VSUBS 0.036658f
C1040 VDD2.n141 VSUBS 0.036658f
C1041 VDD2.n142 VSUBS 0.016421f
C1042 VDD2.n143 VSUBS 0.015509f
C1043 VDD2.n144 VSUBS 0.028862f
C1044 VDD2.n145 VSUBS 0.028862f
C1045 VDD2.n146 VSUBS 0.015509f
C1046 VDD2.n147 VSUBS 0.016421f
C1047 VDD2.n148 VSUBS 0.036658f
C1048 VDD2.n149 VSUBS 0.036658f
C1049 VDD2.n150 VSUBS 0.016421f
C1050 VDD2.n151 VSUBS 0.015509f
C1051 VDD2.n152 VSUBS 0.028862f
C1052 VDD2.n153 VSUBS 0.028862f
C1053 VDD2.n154 VSUBS 0.015509f
C1054 VDD2.n155 VSUBS 0.016421f
C1055 VDD2.n156 VSUBS 0.036658f
C1056 VDD2.n157 VSUBS 0.036658f
C1057 VDD2.n158 VSUBS 0.016421f
C1058 VDD2.n159 VSUBS 0.015509f
C1059 VDD2.n160 VSUBS 0.028862f
C1060 VDD2.n161 VSUBS 0.028862f
C1061 VDD2.n162 VSUBS 0.015509f
C1062 VDD2.n163 VSUBS 0.016421f
C1063 VDD2.n164 VSUBS 0.036658f
C1064 VDD2.n165 VSUBS 0.080833f
C1065 VDD2.n166 VSUBS 0.016421f
C1066 VDD2.n167 VSUBS 0.015509f
C1067 VDD2.n168 VSUBS 0.065925f
C1068 VDD2.n169 VSUBS 0.060209f
C1069 VDD2.n170 VSUBS 4.00487f
C1070 VTAIL.n0 VSUBS 0.029306f
C1071 VTAIL.n1 VSUBS 0.02878f
C1072 VTAIL.n2 VSUBS 0.015465f
C1073 VTAIL.n3 VSUBS 0.036554f
C1074 VTAIL.n4 VSUBS 0.01592f
C1075 VTAIL.n5 VSUBS 0.02878f
C1076 VTAIL.n6 VSUBS 0.016375f
C1077 VTAIL.n7 VSUBS 0.036554f
C1078 VTAIL.n8 VSUBS 0.016375f
C1079 VTAIL.n9 VSUBS 0.02878f
C1080 VTAIL.n10 VSUBS 0.015465f
C1081 VTAIL.n11 VSUBS 0.036554f
C1082 VTAIL.n12 VSUBS 0.016375f
C1083 VTAIL.n13 VSUBS 0.02878f
C1084 VTAIL.n14 VSUBS 0.015465f
C1085 VTAIL.n15 VSUBS 0.036554f
C1086 VTAIL.n16 VSUBS 0.016375f
C1087 VTAIL.n17 VSUBS 0.02878f
C1088 VTAIL.n18 VSUBS 0.015465f
C1089 VTAIL.n19 VSUBS 0.036554f
C1090 VTAIL.n20 VSUBS 0.016375f
C1091 VTAIL.n21 VSUBS 0.02878f
C1092 VTAIL.n22 VSUBS 0.015465f
C1093 VTAIL.n23 VSUBS 0.036554f
C1094 VTAIL.n24 VSUBS 0.016375f
C1095 VTAIL.n25 VSUBS 1.88206f
C1096 VTAIL.n26 VSUBS 0.015465f
C1097 VTAIL.t0 VSUBS 0.078278f
C1098 VTAIL.n27 VSUBS 0.205758f
C1099 VTAIL.n28 VSUBS 0.023254f
C1100 VTAIL.n29 VSUBS 0.027415f
C1101 VTAIL.n30 VSUBS 0.036554f
C1102 VTAIL.n31 VSUBS 0.016375f
C1103 VTAIL.n32 VSUBS 0.015465f
C1104 VTAIL.n33 VSUBS 0.02878f
C1105 VTAIL.n34 VSUBS 0.02878f
C1106 VTAIL.n35 VSUBS 0.015465f
C1107 VTAIL.n36 VSUBS 0.016375f
C1108 VTAIL.n37 VSUBS 0.036554f
C1109 VTAIL.n38 VSUBS 0.036554f
C1110 VTAIL.n39 VSUBS 0.016375f
C1111 VTAIL.n40 VSUBS 0.015465f
C1112 VTAIL.n41 VSUBS 0.02878f
C1113 VTAIL.n42 VSUBS 0.02878f
C1114 VTAIL.n43 VSUBS 0.015465f
C1115 VTAIL.n44 VSUBS 0.016375f
C1116 VTAIL.n45 VSUBS 0.036554f
C1117 VTAIL.n46 VSUBS 0.036554f
C1118 VTAIL.n47 VSUBS 0.016375f
C1119 VTAIL.n48 VSUBS 0.015465f
C1120 VTAIL.n49 VSUBS 0.02878f
C1121 VTAIL.n50 VSUBS 0.02878f
C1122 VTAIL.n51 VSUBS 0.015465f
C1123 VTAIL.n52 VSUBS 0.016375f
C1124 VTAIL.n53 VSUBS 0.036554f
C1125 VTAIL.n54 VSUBS 0.036554f
C1126 VTAIL.n55 VSUBS 0.016375f
C1127 VTAIL.n56 VSUBS 0.015465f
C1128 VTAIL.n57 VSUBS 0.02878f
C1129 VTAIL.n58 VSUBS 0.02878f
C1130 VTAIL.n59 VSUBS 0.015465f
C1131 VTAIL.n60 VSUBS 0.016375f
C1132 VTAIL.n61 VSUBS 0.036554f
C1133 VTAIL.n62 VSUBS 0.036554f
C1134 VTAIL.n63 VSUBS 0.016375f
C1135 VTAIL.n64 VSUBS 0.015465f
C1136 VTAIL.n65 VSUBS 0.02878f
C1137 VTAIL.n66 VSUBS 0.02878f
C1138 VTAIL.n67 VSUBS 0.015465f
C1139 VTAIL.n68 VSUBS 0.015465f
C1140 VTAIL.n69 VSUBS 0.016375f
C1141 VTAIL.n70 VSUBS 0.036554f
C1142 VTAIL.n71 VSUBS 0.036554f
C1143 VTAIL.n72 VSUBS 0.036554f
C1144 VTAIL.n73 VSUBS 0.01592f
C1145 VTAIL.n74 VSUBS 0.015465f
C1146 VTAIL.n75 VSUBS 0.02878f
C1147 VTAIL.n76 VSUBS 0.02878f
C1148 VTAIL.n77 VSUBS 0.015465f
C1149 VTAIL.n78 VSUBS 0.016375f
C1150 VTAIL.n79 VSUBS 0.036554f
C1151 VTAIL.n80 VSUBS 0.080602f
C1152 VTAIL.n81 VSUBS 0.016375f
C1153 VTAIL.n82 VSUBS 0.015465f
C1154 VTAIL.n83 VSUBS 0.065737f
C1155 VTAIL.n84 VSUBS 0.04016f
C1156 VTAIL.n85 VSUBS 2.29115f
C1157 VTAIL.n86 VSUBS 0.029306f
C1158 VTAIL.n87 VSUBS 0.02878f
C1159 VTAIL.n88 VSUBS 0.015465f
C1160 VTAIL.n89 VSUBS 0.036554f
C1161 VTAIL.n90 VSUBS 0.01592f
C1162 VTAIL.n91 VSUBS 0.02878f
C1163 VTAIL.n92 VSUBS 0.01592f
C1164 VTAIL.n93 VSUBS 0.015465f
C1165 VTAIL.n94 VSUBS 0.036554f
C1166 VTAIL.n95 VSUBS 0.036554f
C1167 VTAIL.n96 VSUBS 0.016375f
C1168 VTAIL.n97 VSUBS 0.02878f
C1169 VTAIL.n98 VSUBS 0.015465f
C1170 VTAIL.n99 VSUBS 0.036554f
C1171 VTAIL.n100 VSUBS 0.016375f
C1172 VTAIL.n101 VSUBS 0.02878f
C1173 VTAIL.n102 VSUBS 0.015465f
C1174 VTAIL.n103 VSUBS 0.036554f
C1175 VTAIL.n104 VSUBS 0.016375f
C1176 VTAIL.n105 VSUBS 0.02878f
C1177 VTAIL.n106 VSUBS 0.015465f
C1178 VTAIL.n107 VSUBS 0.036554f
C1179 VTAIL.n108 VSUBS 0.016375f
C1180 VTAIL.n109 VSUBS 0.02878f
C1181 VTAIL.n110 VSUBS 0.015465f
C1182 VTAIL.n111 VSUBS 0.036554f
C1183 VTAIL.n112 VSUBS 0.016375f
C1184 VTAIL.n113 VSUBS 1.88206f
C1185 VTAIL.n114 VSUBS 0.015465f
C1186 VTAIL.t2 VSUBS 0.078278f
C1187 VTAIL.n115 VSUBS 0.205758f
C1188 VTAIL.n116 VSUBS 0.023254f
C1189 VTAIL.n117 VSUBS 0.027415f
C1190 VTAIL.n118 VSUBS 0.036554f
C1191 VTAIL.n119 VSUBS 0.016375f
C1192 VTAIL.n120 VSUBS 0.015465f
C1193 VTAIL.n121 VSUBS 0.02878f
C1194 VTAIL.n122 VSUBS 0.02878f
C1195 VTAIL.n123 VSUBS 0.015465f
C1196 VTAIL.n124 VSUBS 0.016375f
C1197 VTAIL.n125 VSUBS 0.036554f
C1198 VTAIL.n126 VSUBS 0.036554f
C1199 VTAIL.n127 VSUBS 0.016375f
C1200 VTAIL.n128 VSUBS 0.015465f
C1201 VTAIL.n129 VSUBS 0.02878f
C1202 VTAIL.n130 VSUBS 0.02878f
C1203 VTAIL.n131 VSUBS 0.015465f
C1204 VTAIL.n132 VSUBS 0.016375f
C1205 VTAIL.n133 VSUBS 0.036554f
C1206 VTAIL.n134 VSUBS 0.036554f
C1207 VTAIL.n135 VSUBS 0.016375f
C1208 VTAIL.n136 VSUBS 0.015465f
C1209 VTAIL.n137 VSUBS 0.02878f
C1210 VTAIL.n138 VSUBS 0.02878f
C1211 VTAIL.n139 VSUBS 0.015465f
C1212 VTAIL.n140 VSUBS 0.016375f
C1213 VTAIL.n141 VSUBS 0.036554f
C1214 VTAIL.n142 VSUBS 0.036554f
C1215 VTAIL.n143 VSUBS 0.016375f
C1216 VTAIL.n144 VSUBS 0.015465f
C1217 VTAIL.n145 VSUBS 0.02878f
C1218 VTAIL.n146 VSUBS 0.02878f
C1219 VTAIL.n147 VSUBS 0.015465f
C1220 VTAIL.n148 VSUBS 0.016375f
C1221 VTAIL.n149 VSUBS 0.036554f
C1222 VTAIL.n150 VSUBS 0.036554f
C1223 VTAIL.n151 VSUBS 0.016375f
C1224 VTAIL.n152 VSUBS 0.015465f
C1225 VTAIL.n153 VSUBS 0.02878f
C1226 VTAIL.n154 VSUBS 0.02878f
C1227 VTAIL.n155 VSUBS 0.015465f
C1228 VTAIL.n156 VSUBS 0.016375f
C1229 VTAIL.n157 VSUBS 0.036554f
C1230 VTAIL.n158 VSUBS 0.036554f
C1231 VTAIL.n159 VSUBS 0.016375f
C1232 VTAIL.n160 VSUBS 0.015465f
C1233 VTAIL.n161 VSUBS 0.02878f
C1234 VTAIL.n162 VSUBS 0.02878f
C1235 VTAIL.n163 VSUBS 0.015465f
C1236 VTAIL.n164 VSUBS 0.016375f
C1237 VTAIL.n165 VSUBS 0.036554f
C1238 VTAIL.n166 VSUBS 0.080602f
C1239 VTAIL.n167 VSUBS 0.016375f
C1240 VTAIL.n168 VSUBS 0.015465f
C1241 VTAIL.n169 VSUBS 0.065737f
C1242 VTAIL.n170 VSUBS 0.04016f
C1243 VTAIL.n171 VSUBS 2.3525f
C1244 VTAIL.n172 VSUBS 0.029306f
C1245 VTAIL.n173 VSUBS 0.02878f
C1246 VTAIL.n174 VSUBS 0.015465f
C1247 VTAIL.n175 VSUBS 0.036554f
C1248 VTAIL.n176 VSUBS 0.01592f
C1249 VTAIL.n177 VSUBS 0.02878f
C1250 VTAIL.n178 VSUBS 0.01592f
C1251 VTAIL.n179 VSUBS 0.015465f
C1252 VTAIL.n180 VSUBS 0.036554f
C1253 VTAIL.n181 VSUBS 0.036554f
C1254 VTAIL.n182 VSUBS 0.016375f
C1255 VTAIL.n183 VSUBS 0.02878f
C1256 VTAIL.n184 VSUBS 0.015465f
C1257 VTAIL.n185 VSUBS 0.036554f
C1258 VTAIL.n186 VSUBS 0.016375f
C1259 VTAIL.n187 VSUBS 0.02878f
C1260 VTAIL.n188 VSUBS 0.015465f
C1261 VTAIL.n189 VSUBS 0.036554f
C1262 VTAIL.n190 VSUBS 0.016375f
C1263 VTAIL.n191 VSUBS 0.02878f
C1264 VTAIL.n192 VSUBS 0.015465f
C1265 VTAIL.n193 VSUBS 0.036554f
C1266 VTAIL.n194 VSUBS 0.016375f
C1267 VTAIL.n195 VSUBS 0.02878f
C1268 VTAIL.n196 VSUBS 0.015465f
C1269 VTAIL.n197 VSUBS 0.036554f
C1270 VTAIL.n198 VSUBS 0.016375f
C1271 VTAIL.n199 VSUBS 1.88206f
C1272 VTAIL.n200 VSUBS 0.015465f
C1273 VTAIL.t1 VSUBS 0.078278f
C1274 VTAIL.n201 VSUBS 0.205758f
C1275 VTAIL.n202 VSUBS 0.023254f
C1276 VTAIL.n203 VSUBS 0.027415f
C1277 VTAIL.n204 VSUBS 0.036554f
C1278 VTAIL.n205 VSUBS 0.016375f
C1279 VTAIL.n206 VSUBS 0.015465f
C1280 VTAIL.n207 VSUBS 0.02878f
C1281 VTAIL.n208 VSUBS 0.02878f
C1282 VTAIL.n209 VSUBS 0.015465f
C1283 VTAIL.n210 VSUBS 0.016375f
C1284 VTAIL.n211 VSUBS 0.036554f
C1285 VTAIL.n212 VSUBS 0.036554f
C1286 VTAIL.n213 VSUBS 0.016375f
C1287 VTAIL.n214 VSUBS 0.015465f
C1288 VTAIL.n215 VSUBS 0.02878f
C1289 VTAIL.n216 VSUBS 0.02878f
C1290 VTAIL.n217 VSUBS 0.015465f
C1291 VTAIL.n218 VSUBS 0.016375f
C1292 VTAIL.n219 VSUBS 0.036554f
C1293 VTAIL.n220 VSUBS 0.036554f
C1294 VTAIL.n221 VSUBS 0.016375f
C1295 VTAIL.n222 VSUBS 0.015465f
C1296 VTAIL.n223 VSUBS 0.02878f
C1297 VTAIL.n224 VSUBS 0.02878f
C1298 VTAIL.n225 VSUBS 0.015465f
C1299 VTAIL.n226 VSUBS 0.016375f
C1300 VTAIL.n227 VSUBS 0.036554f
C1301 VTAIL.n228 VSUBS 0.036554f
C1302 VTAIL.n229 VSUBS 0.016375f
C1303 VTAIL.n230 VSUBS 0.015465f
C1304 VTAIL.n231 VSUBS 0.02878f
C1305 VTAIL.n232 VSUBS 0.02878f
C1306 VTAIL.n233 VSUBS 0.015465f
C1307 VTAIL.n234 VSUBS 0.016375f
C1308 VTAIL.n235 VSUBS 0.036554f
C1309 VTAIL.n236 VSUBS 0.036554f
C1310 VTAIL.n237 VSUBS 0.016375f
C1311 VTAIL.n238 VSUBS 0.015465f
C1312 VTAIL.n239 VSUBS 0.02878f
C1313 VTAIL.n240 VSUBS 0.02878f
C1314 VTAIL.n241 VSUBS 0.015465f
C1315 VTAIL.n242 VSUBS 0.016375f
C1316 VTAIL.n243 VSUBS 0.036554f
C1317 VTAIL.n244 VSUBS 0.036554f
C1318 VTAIL.n245 VSUBS 0.016375f
C1319 VTAIL.n246 VSUBS 0.015465f
C1320 VTAIL.n247 VSUBS 0.02878f
C1321 VTAIL.n248 VSUBS 0.02878f
C1322 VTAIL.n249 VSUBS 0.015465f
C1323 VTAIL.n250 VSUBS 0.016375f
C1324 VTAIL.n251 VSUBS 0.036554f
C1325 VTAIL.n252 VSUBS 0.080602f
C1326 VTAIL.n253 VSUBS 0.016375f
C1327 VTAIL.n254 VSUBS 0.015465f
C1328 VTAIL.n255 VSUBS 0.065737f
C1329 VTAIL.n256 VSUBS 0.04016f
C1330 VTAIL.n257 VSUBS 2.08549f
C1331 VTAIL.n258 VSUBS 0.029306f
C1332 VTAIL.n259 VSUBS 0.02878f
C1333 VTAIL.n260 VSUBS 0.015465f
C1334 VTAIL.n261 VSUBS 0.036554f
C1335 VTAIL.n262 VSUBS 0.01592f
C1336 VTAIL.n263 VSUBS 0.02878f
C1337 VTAIL.n264 VSUBS 0.016375f
C1338 VTAIL.n265 VSUBS 0.036554f
C1339 VTAIL.n266 VSUBS 0.016375f
C1340 VTAIL.n267 VSUBS 0.02878f
C1341 VTAIL.n268 VSUBS 0.015465f
C1342 VTAIL.n269 VSUBS 0.036554f
C1343 VTAIL.n270 VSUBS 0.016375f
C1344 VTAIL.n271 VSUBS 0.02878f
C1345 VTAIL.n272 VSUBS 0.015465f
C1346 VTAIL.n273 VSUBS 0.036554f
C1347 VTAIL.n274 VSUBS 0.016375f
C1348 VTAIL.n275 VSUBS 0.02878f
C1349 VTAIL.n276 VSUBS 0.015465f
C1350 VTAIL.n277 VSUBS 0.036554f
C1351 VTAIL.n278 VSUBS 0.016375f
C1352 VTAIL.n279 VSUBS 0.02878f
C1353 VTAIL.n280 VSUBS 0.015465f
C1354 VTAIL.n281 VSUBS 0.036554f
C1355 VTAIL.n282 VSUBS 0.016375f
C1356 VTAIL.n283 VSUBS 1.88206f
C1357 VTAIL.n284 VSUBS 0.015465f
C1358 VTAIL.t3 VSUBS 0.078278f
C1359 VTAIL.n285 VSUBS 0.205758f
C1360 VTAIL.n286 VSUBS 0.023254f
C1361 VTAIL.n287 VSUBS 0.027415f
C1362 VTAIL.n288 VSUBS 0.036554f
C1363 VTAIL.n289 VSUBS 0.016375f
C1364 VTAIL.n290 VSUBS 0.015465f
C1365 VTAIL.n291 VSUBS 0.02878f
C1366 VTAIL.n292 VSUBS 0.02878f
C1367 VTAIL.n293 VSUBS 0.015465f
C1368 VTAIL.n294 VSUBS 0.016375f
C1369 VTAIL.n295 VSUBS 0.036554f
C1370 VTAIL.n296 VSUBS 0.036554f
C1371 VTAIL.n297 VSUBS 0.016375f
C1372 VTAIL.n298 VSUBS 0.015465f
C1373 VTAIL.n299 VSUBS 0.02878f
C1374 VTAIL.n300 VSUBS 0.02878f
C1375 VTAIL.n301 VSUBS 0.015465f
C1376 VTAIL.n302 VSUBS 0.016375f
C1377 VTAIL.n303 VSUBS 0.036554f
C1378 VTAIL.n304 VSUBS 0.036554f
C1379 VTAIL.n305 VSUBS 0.016375f
C1380 VTAIL.n306 VSUBS 0.015465f
C1381 VTAIL.n307 VSUBS 0.02878f
C1382 VTAIL.n308 VSUBS 0.02878f
C1383 VTAIL.n309 VSUBS 0.015465f
C1384 VTAIL.n310 VSUBS 0.016375f
C1385 VTAIL.n311 VSUBS 0.036554f
C1386 VTAIL.n312 VSUBS 0.036554f
C1387 VTAIL.n313 VSUBS 0.016375f
C1388 VTAIL.n314 VSUBS 0.015465f
C1389 VTAIL.n315 VSUBS 0.02878f
C1390 VTAIL.n316 VSUBS 0.02878f
C1391 VTAIL.n317 VSUBS 0.015465f
C1392 VTAIL.n318 VSUBS 0.016375f
C1393 VTAIL.n319 VSUBS 0.036554f
C1394 VTAIL.n320 VSUBS 0.036554f
C1395 VTAIL.n321 VSUBS 0.016375f
C1396 VTAIL.n322 VSUBS 0.015465f
C1397 VTAIL.n323 VSUBS 0.02878f
C1398 VTAIL.n324 VSUBS 0.02878f
C1399 VTAIL.n325 VSUBS 0.015465f
C1400 VTAIL.n326 VSUBS 0.015465f
C1401 VTAIL.n327 VSUBS 0.016375f
C1402 VTAIL.n328 VSUBS 0.036554f
C1403 VTAIL.n329 VSUBS 0.036554f
C1404 VTAIL.n330 VSUBS 0.036554f
C1405 VTAIL.n331 VSUBS 0.01592f
C1406 VTAIL.n332 VSUBS 0.015465f
C1407 VTAIL.n333 VSUBS 0.02878f
C1408 VTAIL.n334 VSUBS 0.02878f
C1409 VTAIL.n335 VSUBS 0.015465f
C1410 VTAIL.n336 VSUBS 0.016375f
C1411 VTAIL.n337 VSUBS 0.036554f
C1412 VTAIL.n338 VSUBS 0.080602f
C1413 VTAIL.n339 VSUBS 0.016375f
C1414 VTAIL.n340 VSUBS 0.015465f
C1415 VTAIL.n341 VSUBS 0.065737f
C1416 VTAIL.n342 VSUBS 0.04016f
C1417 VTAIL.n343 VSUBS 1.96978f
C1418 VN.t1 VSUBS 4.81156f
C1419 VN.t0 VSUBS 5.56123f
.ends

