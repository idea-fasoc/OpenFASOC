* NGSPICE file created from diff_pair_sample_0227.ext - technology: sky130A

.subckt diff_pair_sample_0227 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=0 ps=0 w=10.55 l=2.49
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=0 ps=0 w=10.55 l=2.49
X2 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=4.1145 ps=21.88 w=10.55 l=2.49
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=0 ps=0 w=10.55 l=2.49
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=4.1145 ps=21.88 w=10.55 l=2.49
X5 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=4.1145 ps=21.88 w=10.55 l=2.49
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=0 ps=0 w=10.55 l=2.49
X7 VDD2.t0 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1145 pd=21.88 as=4.1145 ps=21.88 w=10.55 l=2.49
R0 B.n627 B.n626 585
R1 B.n259 B.n90 585
R2 B.n258 B.n257 585
R3 B.n256 B.n255 585
R4 B.n254 B.n253 585
R5 B.n252 B.n251 585
R6 B.n250 B.n249 585
R7 B.n248 B.n247 585
R8 B.n246 B.n245 585
R9 B.n244 B.n243 585
R10 B.n242 B.n241 585
R11 B.n240 B.n239 585
R12 B.n238 B.n237 585
R13 B.n236 B.n235 585
R14 B.n234 B.n233 585
R15 B.n232 B.n231 585
R16 B.n230 B.n229 585
R17 B.n228 B.n227 585
R18 B.n226 B.n225 585
R19 B.n224 B.n223 585
R20 B.n222 B.n221 585
R21 B.n220 B.n219 585
R22 B.n218 B.n217 585
R23 B.n216 B.n215 585
R24 B.n214 B.n213 585
R25 B.n212 B.n211 585
R26 B.n210 B.n209 585
R27 B.n208 B.n207 585
R28 B.n206 B.n205 585
R29 B.n204 B.n203 585
R30 B.n202 B.n201 585
R31 B.n200 B.n199 585
R32 B.n198 B.n197 585
R33 B.n196 B.n195 585
R34 B.n194 B.n193 585
R35 B.n192 B.n191 585
R36 B.n190 B.n189 585
R37 B.n187 B.n186 585
R38 B.n185 B.n184 585
R39 B.n183 B.n182 585
R40 B.n181 B.n180 585
R41 B.n179 B.n178 585
R42 B.n177 B.n176 585
R43 B.n175 B.n174 585
R44 B.n173 B.n172 585
R45 B.n171 B.n170 585
R46 B.n169 B.n168 585
R47 B.n166 B.n165 585
R48 B.n164 B.n163 585
R49 B.n162 B.n161 585
R50 B.n160 B.n159 585
R51 B.n158 B.n157 585
R52 B.n156 B.n155 585
R53 B.n154 B.n153 585
R54 B.n152 B.n151 585
R55 B.n150 B.n149 585
R56 B.n148 B.n147 585
R57 B.n146 B.n145 585
R58 B.n144 B.n143 585
R59 B.n142 B.n141 585
R60 B.n140 B.n139 585
R61 B.n138 B.n137 585
R62 B.n136 B.n135 585
R63 B.n134 B.n133 585
R64 B.n132 B.n131 585
R65 B.n130 B.n129 585
R66 B.n128 B.n127 585
R67 B.n126 B.n125 585
R68 B.n124 B.n123 585
R69 B.n122 B.n121 585
R70 B.n120 B.n119 585
R71 B.n118 B.n117 585
R72 B.n116 B.n115 585
R73 B.n114 B.n113 585
R74 B.n112 B.n111 585
R75 B.n110 B.n109 585
R76 B.n108 B.n107 585
R77 B.n106 B.n105 585
R78 B.n104 B.n103 585
R79 B.n102 B.n101 585
R80 B.n100 B.n99 585
R81 B.n98 B.n97 585
R82 B.n96 B.n95 585
R83 B.n47 B.n46 585
R84 B.n625 B.n48 585
R85 B.n630 B.n48 585
R86 B.n624 B.n623 585
R87 B.n623 B.n44 585
R88 B.n622 B.n43 585
R89 B.n636 B.n43 585
R90 B.n621 B.n42 585
R91 B.n637 B.n42 585
R92 B.n620 B.n41 585
R93 B.n638 B.n41 585
R94 B.n619 B.n618 585
R95 B.n618 B.n37 585
R96 B.n617 B.n36 585
R97 B.n644 B.n36 585
R98 B.n616 B.n35 585
R99 B.n645 B.n35 585
R100 B.n615 B.n34 585
R101 B.n646 B.n34 585
R102 B.n614 B.n613 585
R103 B.n613 B.n30 585
R104 B.n612 B.n29 585
R105 B.n652 B.n29 585
R106 B.n611 B.n28 585
R107 B.n653 B.n28 585
R108 B.n610 B.n27 585
R109 B.n654 B.n27 585
R110 B.n609 B.n608 585
R111 B.n608 B.n23 585
R112 B.n607 B.n22 585
R113 B.n660 B.n22 585
R114 B.n606 B.n21 585
R115 B.n661 B.n21 585
R116 B.n605 B.n20 585
R117 B.n662 B.n20 585
R118 B.n604 B.n603 585
R119 B.n603 B.n16 585
R120 B.n602 B.n15 585
R121 B.n668 B.n15 585
R122 B.n601 B.n14 585
R123 B.n669 B.n14 585
R124 B.n600 B.n13 585
R125 B.n670 B.n13 585
R126 B.n599 B.n598 585
R127 B.n598 B.n12 585
R128 B.n597 B.n596 585
R129 B.n597 B.n8 585
R130 B.n595 B.n7 585
R131 B.n677 B.n7 585
R132 B.n594 B.n6 585
R133 B.n678 B.n6 585
R134 B.n593 B.n5 585
R135 B.n679 B.n5 585
R136 B.n592 B.n591 585
R137 B.n591 B.n4 585
R138 B.n590 B.n260 585
R139 B.n590 B.n589 585
R140 B.n580 B.n261 585
R141 B.n262 B.n261 585
R142 B.n582 B.n581 585
R143 B.n583 B.n582 585
R144 B.n579 B.n267 585
R145 B.n267 B.n266 585
R146 B.n578 B.n577 585
R147 B.n577 B.n576 585
R148 B.n269 B.n268 585
R149 B.n270 B.n269 585
R150 B.n569 B.n568 585
R151 B.n570 B.n569 585
R152 B.n567 B.n275 585
R153 B.n275 B.n274 585
R154 B.n566 B.n565 585
R155 B.n565 B.n564 585
R156 B.n277 B.n276 585
R157 B.n278 B.n277 585
R158 B.n557 B.n556 585
R159 B.n558 B.n557 585
R160 B.n555 B.n283 585
R161 B.n283 B.n282 585
R162 B.n554 B.n553 585
R163 B.n553 B.n552 585
R164 B.n285 B.n284 585
R165 B.n286 B.n285 585
R166 B.n545 B.n544 585
R167 B.n546 B.n545 585
R168 B.n543 B.n290 585
R169 B.n294 B.n290 585
R170 B.n542 B.n541 585
R171 B.n541 B.n540 585
R172 B.n292 B.n291 585
R173 B.n293 B.n292 585
R174 B.n533 B.n532 585
R175 B.n534 B.n533 585
R176 B.n531 B.n299 585
R177 B.n299 B.n298 585
R178 B.n530 B.n529 585
R179 B.n529 B.n528 585
R180 B.n301 B.n300 585
R181 B.n302 B.n301 585
R182 B.n521 B.n520 585
R183 B.n522 B.n521 585
R184 B.n305 B.n304 585
R185 B.n356 B.n355 585
R186 B.n357 B.n353 585
R187 B.n353 B.n306 585
R188 B.n359 B.n358 585
R189 B.n361 B.n352 585
R190 B.n364 B.n363 585
R191 B.n365 B.n351 585
R192 B.n367 B.n366 585
R193 B.n369 B.n350 585
R194 B.n372 B.n371 585
R195 B.n373 B.n349 585
R196 B.n375 B.n374 585
R197 B.n377 B.n348 585
R198 B.n380 B.n379 585
R199 B.n381 B.n347 585
R200 B.n383 B.n382 585
R201 B.n385 B.n346 585
R202 B.n388 B.n387 585
R203 B.n389 B.n345 585
R204 B.n391 B.n390 585
R205 B.n393 B.n344 585
R206 B.n396 B.n395 585
R207 B.n397 B.n343 585
R208 B.n399 B.n398 585
R209 B.n401 B.n342 585
R210 B.n404 B.n403 585
R211 B.n405 B.n341 585
R212 B.n407 B.n406 585
R213 B.n409 B.n340 585
R214 B.n412 B.n411 585
R215 B.n413 B.n339 585
R216 B.n415 B.n414 585
R217 B.n417 B.n338 585
R218 B.n420 B.n419 585
R219 B.n421 B.n337 585
R220 B.n423 B.n422 585
R221 B.n425 B.n336 585
R222 B.n428 B.n427 585
R223 B.n429 B.n332 585
R224 B.n431 B.n430 585
R225 B.n433 B.n331 585
R226 B.n436 B.n435 585
R227 B.n437 B.n330 585
R228 B.n439 B.n438 585
R229 B.n441 B.n329 585
R230 B.n444 B.n443 585
R231 B.n445 B.n326 585
R232 B.n448 B.n447 585
R233 B.n450 B.n325 585
R234 B.n453 B.n452 585
R235 B.n454 B.n324 585
R236 B.n456 B.n455 585
R237 B.n458 B.n323 585
R238 B.n461 B.n460 585
R239 B.n462 B.n322 585
R240 B.n464 B.n463 585
R241 B.n466 B.n321 585
R242 B.n469 B.n468 585
R243 B.n470 B.n320 585
R244 B.n472 B.n471 585
R245 B.n474 B.n319 585
R246 B.n477 B.n476 585
R247 B.n478 B.n318 585
R248 B.n480 B.n479 585
R249 B.n482 B.n317 585
R250 B.n485 B.n484 585
R251 B.n486 B.n316 585
R252 B.n488 B.n487 585
R253 B.n490 B.n315 585
R254 B.n493 B.n492 585
R255 B.n494 B.n314 585
R256 B.n496 B.n495 585
R257 B.n498 B.n313 585
R258 B.n501 B.n500 585
R259 B.n502 B.n312 585
R260 B.n504 B.n503 585
R261 B.n506 B.n311 585
R262 B.n509 B.n508 585
R263 B.n510 B.n310 585
R264 B.n512 B.n511 585
R265 B.n514 B.n309 585
R266 B.n515 B.n308 585
R267 B.n518 B.n517 585
R268 B.n519 B.n307 585
R269 B.n307 B.n306 585
R270 B.n524 B.n523 585
R271 B.n523 B.n522 585
R272 B.n525 B.n303 585
R273 B.n303 B.n302 585
R274 B.n527 B.n526 585
R275 B.n528 B.n527 585
R276 B.n297 B.n296 585
R277 B.n298 B.n297 585
R278 B.n536 B.n535 585
R279 B.n535 B.n534 585
R280 B.n537 B.n295 585
R281 B.n295 B.n293 585
R282 B.n539 B.n538 585
R283 B.n540 B.n539 585
R284 B.n289 B.n288 585
R285 B.n294 B.n289 585
R286 B.n548 B.n547 585
R287 B.n547 B.n546 585
R288 B.n549 B.n287 585
R289 B.n287 B.n286 585
R290 B.n551 B.n550 585
R291 B.n552 B.n551 585
R292 B.n281 B.n280 585
R293 B.n282 B.n281 585
R294 B.n560 B.n559 585
R295 B.n559 B.n558 585
R296 B.n561 B.n279 585
R297 B.n279 B.n278 585
R298 B.n563 B.n562 585
R299 B.n564 B.n563 585
R300 B.n273 B.n272 585
R301 B.n274 B.n273 585
R302 B.n572 B.n571 585
R303 B.n571 B.n570 585
R304 B.n573 B.n271 585
R305 B.n271 B.n270 585
R306 B.n575 B.n574 585
R307 B.n576 B.n575 585
R308 B.n265 B.n264 585
R309 B.n266 B.n265 585
R310 B.n585 B.n584 585
R311 B.n584 B.n583 585
R312 B.n586 B.n263 585
R313 B.n263 B.n262 585
R314 B.n588 B.n587 585
R315 B.n589 B.n588 585
R316 B.n3 B.n0 585
R317 B.n4 B.n3 585
R318 B.n676 B.n1 585
R319 B.n677 B.n676 585
R320 B.n675 B.n674 585
R321 B.n675 B.n8 585
R322 B.n673 B.n9 585
R323 B.n12 B.n9 585
R324 B.n672 B.n671 585
R325 B.n671 B.n670 585
R326 B.n11 B.n10 585
R327 B.n669 B.n11 585
R328 B.n667 B.n666 585
R329 B.n668 B.n667 585
R330 B.n665 B.n17 585
R331 B.n17 B.n16 585
R332 B.n664 B.n663 585
R333 B.n663 B.n662 585
R334 B.n19 B.n18 585
R335 B.n661 B.n19 585
R336 B.n659 B.n658 585
R337 B.n660 B.n659 585
R338 B.n657 B.n24 585
R339 B.n24 B.n23 585
R340 B.n656 B.n655 585
R341 B.n655 B.n654 585
R342 B.n26 B.n25 585
R343 B.n653 B.n26 585
R344 B.n651 B.n650 585
R345 B.n652 B.n651 585
R346 B.n649 B.n31 585
R347 B.n31 B.n30 585
R348 B.n648 B.n647 585
R349 B.n647 B.n646 585
R350 B.n33 B.n32 585
R351 B.n645 B.n33 585
R352 B.n643 B.n642 585
R353 B.n644 B.n643 585
R354 B.n641 B.n38 585
R355 B.n38 B.n37 585
R356 B.n640 B.n639 585
R357 B.n639 B.n638 585
R358 B.n40 B.n39 585
R359 B.n637 B.n40 585
R360 B.n635 B.n634 585
R361 B.n636 B.n635 585
R362 B.n633 B.n45 585
R363 B.n45 B.n44 585
R364 B.n632 B.n631 585
R365 B.n631 B.n630 585
R366 B.n680 B.n679 585
R367 B.n678 B.n2 585
R368 B.n631 B.n47 554.963
R369 B.n627 B.n48 554.963
R370 B.n521 B.n307 554.963
R371 B.n523 B.n305 554.963
R372 B.n91 B.t4 311.529
R373 B.n327 B.t9 311.529
R374 B.n93 B.t14 311.529
R375 B.n333 B.t12 311.529
R376 B.n93 B.t13 309.986
R377 B.n91 B.t2 309.986
R378 B.n327 B.t6 309.986
R379 B.n333 B.t10 309.986
R380 B.n92 B.t5 256.839
R381 B.n328 B.t8 256.839
R382 B.n94 B.t15 256.837
R383 B.n334 B.t11 256.837
R384 B.n629 B.n628 256.663
R385 B.n629 B.n89 256.663
R386 B.n629 B.n88 256.663
R387 B.n629 B.n87 256.663
R388 B.n629 B.n86 256.663
R389 B.n629 B.n85 256.663
R390 B.n629 B.n84 256.663
R391 B.n629 B.n83 256.663
R392 B.n629 B.n82 256.663
R393 B.n629 B.n81 256.663
R394 B.n629 B.n80 256.663
R395 B.n629 B.n79 256.663
R396 B.n629 B.n78 256.663
R397 B.n629 B.n77 256.663
R398 B.n629 B.n76 256.663
R399 B.n629 B.n75 256.663
R400 B.n629 B.n74 256.663
R401 B.n629 B.n73 256.663
R402 B.n629 B.n72 256.663
R403 B.n629 B.n71 256.663
R404 B.n629 B.n70 256.663
R405 B.n629 B.n69 256.663
R406 B.n629 B.n68 256.663
R407 B.n629 B.n67 256.663
R408 B.n629 B.n66 256.663
R409 B.n629 B.n65 256.663
R410 B.n629 B.n64 256.663
R411 B.n629 B.n63 256.663
R412 B.n629 B.n62 256.663
R413 B.n629 B.n61 256.663
R414 B.n629 B.n60 256.663
R415 B.n629 B.n59 256.663
R416 B.n629 B.n58 256.663
R417 B.n629 B.n57 256.663
R418 B.n629 B.n56 256.663
R419 B.n629 B.n55 256.663
R420 B.n629 B.n54 256.663
R421 B.n629 B.n53 256.663
R422 B.n629 B.n52 256.663
R423 B.n629 B.n51 256.663
R424 B.n629 B.n50 256.663
R425 B.n629 B.n49 256.663
R426 B.n354 B.n306 256.663
R427 B.n360 B.n306 256.663
R428 B.n362 B.n306 256.663
R429 B.n368 B.n306 256.663
R430 B.n370 B.n306 256.663
R431 B.n376 B.n306 256.663
R432 B.n378 B.n306 256.663
R433 B.n384 B.n306 256.663
R434 B.n386 B.n306 256.663
R435 B.n392 B.n306 256.663
R436 B.n394 B.n306 256.663
R437 B.n400 B.n306 256.663
R438 B.n402 B.n306 256.663
R439 B.n408 B.n306 256.663
R440 B.n410 B.n306 256.663
R441 B.n416 B.n306 256.663
R442 B.n418 B.n306 256.663
R443 B.n424 B.n306 256.663
R444 B.n426 B.n306 256.663
R445 B.n432 B.n306 256.663
R446 B.n434 B.n306 256.663
R447 B.n440 B.n306 256.663
R448 B.n442 B.n306 256.663
R449 B.n449 B.n306 256.663
R450 B.n451 B.n306 256.663
R451 B.n457 B.n306 256.663
R452 B.n459 B.n306 256.663
R453 B.n465 B.n306 256.663
R454 B.n467 B.n306 256.663
R455 B.n473 B.n306 256.663
R456 B.n475 B.n306 256.663
R457 B.n481 B.n306 256.663
R458 B.n483 B.n306 256.663
R459 B.n489 B.n306 256.663
R460 B.n491 B.n306 256.663
R461 B.n497 B.n306 256.663
R462 B.n499 B.n306 256.663
R463 B.n505 B.n306 256.663
R464 B.n507 B.n306 256.663
R465 B.n513 B.n306 256.663
R466 B.n516 B.n306 256.663
R467 B.n682 B.n681 256.663
R468 B.n97 B.n96 163.367
R469 B.n101 B.n100 163.367
R470 B.n105 B.n104 163.367
R471 B.n109 B.n108 163.367
R472 B.n113 B.n112 163.367
R473 B.n117 B.n116 163.367
R474 B.n121 B.n120 163.367
R475 B.n125 B.n124 163.367
R476 B.n129 B.n128 163.367
R477 B.n133 B.n132 163.367
R478 B.n137 B.n136 163.367
R479 B.n141 B.n140 163.367
R480 B.n145 B.n144 163.367
R481 B.n149 B.n148 163.367
R482 B.n153 B.n152 163.367
R483 B.n157 B.n156 163.367
R484 B.n161 B.n160 163.367
R485 B.n165 B.n164 163.367
R486 B.n170 B.n169 163.367
R487 B.n174 B.n173 163.367
R488 B.n178 B.n177 163.367
R489 B.n182 B.n181 163.367
R490 B.n186 B.n185 163.367
R491 B.n191 B.n190 163.367
R492 B.n195 B.n194 163.367
R493 B.n199 B.n198 163.367
R494 B.n203 B.n202 163.367
R495 B.n207 B.n206 163.367
R496 B.n211 B.n210 163.367
R497 B.n215 B.n214 163.367
R498 B.n219 B.n218 163.367
R499 B.n223 B.n222 163.367
R500 B.n227 B.n226 163.367
R501 B.n231 B.n230 163.367
R502 B.n235 B.n234 163.367
R503 B.n239 B.n238 163.367
R504 B.n243 B.n242 163.367
R505 B.n247 B.n246 163.367
R506 B.n251 B.n250 163.367
R507 B.n255 B.n254 163.367
R508 B.n257 B.n90 163.367
R509 B.n521 B.n301 163.367
R510 B.n529 B.n301 163.367
R511 B.n529 B.n299 163.367
R512 B.n533 B.n299 163.367
R513 B.n533 B.n292 163.367
R514 B.n541 B.n292 163.367
R515 B.n541 B.n290 163.367
R516 B.n545 B.n290 163.367
R517 B.n545 B.n285 163.367
R518 B.n553 B.n285 163.367
R519 B.n553 B.n283 163.367
R520 B.n557 B.n283 163.367
R521 B.n557 B.n277 163.367
R522 B.n565 B.n277 163.367
R523 B.n565 B.n275 163.367
R524 B.n569 B.n275 163.367
R525 B.n569 B.n269 163.367
R526 B.n577 B.n269 163.367
R527 B.n577 B.n267 163.367
R528 B.n582 B.n267 163.367
R529 B.n582 B.n261 163.367
R530 B.n590 B.n261 163.367
R531 B.n591 B.n590 163.367
R532 B.n591 B.n5 163.367
R533 B.n6 B.n5 163.367
R534 B.n7 B.n6 163.367
R535 B.n597 B.n7 163.367
R536 B.n598 B.n597 163.367
R537 B.n598 B.n13 163.367
R538 B.n14 B.n13 163.367
R539 B.n15 B.n14 163.367
R540 B.n603 B.n15 163.367
R541 B.n603 B.n20 163.367
R542 B.n21 B.n20 163.367
R543 B.n22 B.n21 163.367
R544 B.n608 B.n22 163.367
R545 B.n608 B.n27 163.367
R546 B.n28 B.n27 163.367
R547 B.n29 B.n28 163.367
R548 B.n613 B.n29 163.367
R549 B.n613 B.n34 163.367
R550 B.n35 B.n34 163.367
R551 B.n36 B.n35 163.367
R552 B.n618 B.n36 163.367
R553 B.n618 B.n41 163.367
R554 B.n42 B.n41 163.367
R555 B.n43 B.n42 163.367
R556 B.n623 B.n43 163.367
R557 B.n623 B.n48 163.367
R558 B.n355 B.n353 163.367
R559 B.n359 B.n353 163.367
R560 B.n363 B.n361 163.367
R561 B.n367 B.n351 163.367
R562 B.n371 B.n369 163.367
R563 B.n375 B.n349 163.367
R564 B.n379 B.n377 163.367
R565 B.n383 B.n347 163.367
R566 B.n387 B.n385 163.367
R567 B.n391 B.n345 163.367
R568 B.n395 B.n393 163.367
R569 B.n399 B.n343 163.367
R570 B.n403 B.n401 163.367
R571 B.n407 B.n341 163.367
R572 B.n411 B.n409 163.367
R573 B.n415 B.n339 163.367
R574 B.n419 B.n417 163.367
R575 B.n423 B.n337 163.367
R576 B.n427 B.n425 163.367
R577 B.n431 B.n332 163.367
R578 B.n435 B.n433 163.367
R579 B.n439 B.n330 163.367
R580 B.n443 B.n441 163.367
R581 B.n448 B.n326 163.367
R582 B.n452 B.n450 163.367
R583 B.n456 B.n324 163.367
R584 B.n460 B.n458 163.367
R585 B.n464 B.n322 163.367
R586 B.n468 B.n466 163.367
R587 B.n472 B.n320 163.367
R588 B.n476 B.n474 163.367
R589 B.n480 B.n318 163.367
R590 B.n484 B.n482 163.367
R591 B.n488 B.n316 163.367
R592 B.n492 B.n490 163.367
R593 B.n496 B.n314 163.367
R594 B.n500 B.n498 163.367
R595 B.n504 B.n312 163.367
R596 B.n508 B.n506 163.367
R597 B.n512 B.n310 163.367
R598 B.n515 B.n514 163.367
R599 B.n517 B.n307 163.367
R600 B.n523 B.n303 163.367
R601 B.n527 B.n303 163.367
R602 B.n527 B.n297 163.367
R603 B.n535 B.n297 163.367
R604 B.n535 B.n295 163.367
R605 B.n539 B.n295 163.367
R606 B.n539 B.n289 163.367
R607 B.n547 B.n289 163.367
R608 B.n547 B.n287 163.367
R609 B.n551 B.n287 163.367
R610 B.n551 B.n281 163.367
R611 B.n559 B.n281 163.367
R612 B.n559 B.n279 163.367
R613 B.n563 B.n279 163.367
R614 B.n563 B.n273 163.367
R615 B.n571 B.n273 163.367
R616 B.n571 B.n271 163.367
R617 B.n575 B.n271 163.367
R618 B.n575 B.n265 163.367
R619 B.n584 B.n265 163.367
R620 B.n584 B.n263 163.367
R621 B.n588 B.n263 163.367
R622 B.n588 B.n3 163.367
R623 B.n680 B.n3 163.367
R624 B.n676 B.n2 163.367
R625 B.n676 B.n675 163.367
R626 B.n675 B.n9 163.367
R627 B.n671 B.n9 163.367
R628 B.n671 B.n11 163.367
R629 B.n667 B.n11 163.367
R630 B.n667 B.n17 163.367
R631 B.n663 B.n17 163.367
R632 B.n663 B.n19 163.367
R633 B.n659 B.n19 163.367
R634 B.n659 B.n24 163.367
R635 B.n655 B.n24 163.367
R636 B.n655 B.n26 163.367
R637 B.n651 B.n26 163.367
R638 B.n651 B.n31 163.367
R639 B.n647 B.n31 163.367
R640 B.n647 B.n33 163.367
R641 B.n643 B.n33 163.367
R642 B.n643 B.n38 163.367
R643 B.n639 B.n38 163.367
R644 B.n639 B.n40 163.367
R645 B.n635 B.n40 163.367
R646 B.n635 B.n45 163.367
R647 B.n631 B.n45 163.367
R648 B.n522 B.n306 95.2296
R649 B.n630 B.n629 95.2296
R650 B.n49 B.n47 71.676
R651 B.n97 B.n50 71.676
R652 B.n101 B.n51 71.676
R653 B.n105 B.n52 71.676
R654 B.n109 B.n53 71.676
R655 B.n113 B.n54 71.676
R656 B.n117 B.n55 71.676
R657 B.n121 B.n56 71.676
R658 B.n125 B.n57 71.676
R659 B.n129 B.n58 71.676
R660 B.n133 B.n59 71.676
R661 B.n137 B.n60 71.676
R662 B.n141 B.n61 71.676
R663 B.n145 B.n62 71.676
R664 B.n149 B.n63 71.676
R665 B.n153 B.n64 71.676
R666 B.n157 B.n65 71.676
R667 B.n161 B.n66 71.676
R668 B.n165 B.n67 71.676
R669 B.n170 B.n68 71.676
R670 B.n174 B.n69 71.676
R671 B.n178 B.n70 71.676
R672 B.n182 B.n71 71.676
R673 B.n186 B.n72 71.676
R674 B.n191 B.n73 71.676
R675 B.n195 B.n74 71.676
R676 B.n199 B.n75 71.676
R677 B.n203 B.n76 71.676
R678 B.n207 B.n77 71.676
R679 B.n211 B.n78 71.676
R680 B.n215 B.n79 71.676
R681 B.n219 B.n80 71.676
R682 B.n223 B.n81 71.676
R683 B.n227 B.n82 71.676
R684 B.n231 B.n83 71.676
R685 B.n235 B.n84 71.676
R686 B.n239 B.n85 71.676
R687 B.n243 B.n86 71.676
R688 B.n247 B.n87 71.676
R689 B.n251 B.n88 71.676
R690 B.n255 B.n89 71.676
R691 B.n628 B.n90 71.676
R692 B.n628 B.n627 71.676
R693 B.n257 B.n89 71.676
R694 B.n254 B.n88 71.676
R695 B.n250 B.n87 71.676
R696 B.n246 B.n86 71.676
R697 B.n242 B.n85 71.676
R698 B.n238 B.n84 71.676
R699 B.n234 B.n83 71.676
R700 B.n230 B.n82 71.676
R701 B.n226 B.n81 71.676
R702 B.n222 B.n80 71.676
R703 B.n218 B.n79 71.676
R704 B.n214 B.n78 71.676
R705 B.n210 B.n77 71.676
R706 B.n206 B.n76 71.676
R707 B.n202 B.n75 71.676
R708 B.n198 B.n74 71.676
R709 B.n194 B.n73 71.676
R710 B.n190 B.n72 71.676
R711 B.n185 B.n71 71.676
R712 B.n181 B.n70 71.676
R713 B.n177 B.n69 71.676
R714 B.n173 B.n68 71.676
R715 B.n169 B.n67 71.676
R716 B.n164 B.n66 71.676
R717 B.n160 B.n65 71.676
R718 B.n156 B.n64 71.676
R719 B.n152 B.n63 71.676
R720 B.n148 B.n62 71.676
R721 B.n144 B.n61 71.676
R722 B.n140 B.n60 71.676
R723 B.n136 B.n59 71.676
R724 B.n132 B.n58 71.676
R725 B.n128 B.n57 71.676
R726 B.n124 B.n56 71.676
R727 B.n120 B.n55 71.676
R728 B.n116 B.n54 71.676
R729 B.n112 B.n53 71.676
R730 B.n108 B.n52 71.676
R731 B.n104 B.n51 71.676
R732 B.n100 B.n50 71.676
R733 B.n96 B.n49 71.676
R734 B.n354 B.n305 71.676
R735 B.n360 B.n359 71.676
R736 B.n363 B.n362 71.676
R737 B.n368 B.n367 71.676
R738 B.n371 B.n370 71.676
R739 B.n376 B.n375 71.676
R740 B.n379 B.n378 71.676
R741 B.n384 B.n383 71.676
R742 B.n387 B.n386 71.676
R743 B.n392 B.n391 71.676
R744 B.n395 B.n394 71.676
R745 B.n400 B.n399 71.676
R746 B.n403 B.n402 71.676
R747 B.n408 B.n407 71.676
R748 B.n411 B.n410 71.676
R749 B.n416 B.n415 71.676
R750 B.n419 B.n418 71.676
R751 B.n424 B.n423 71.676
R752 B.n427 B.n426 71.676
R753 B.n432 B.n431 71.676
R754 B.n435 B.n434 71.676
R755 B.n440 B.n439 71.676
R756 B.n443 B.n442 71.676
R757 B.n449 B.n448 71.676
R758 B.n452 B.n451 71.676
R759 B.n457 B.n456 71.676
R760 B.n460 B.n459 71.676
R761 B.n465 B.n464 71.676
R762 B.n468 B.n467 71.676
R763 B.n473 B.n472 71.676
R764 B.n476 B.n475 71.676
R765 B.n481 B.n480 71.676
R766 B.n484 B.n483 71.676
R767 B.n489 B.n488 71.676
R768 B.n492 B.n491 71.676
R769 B.n497 B.n496 71.676
R770 B.n500 B.n499 71.676
R771 B.n505 B.n504 71.676
R772 B.n508 B.n507 71.676
R773 B.n513 B.n512 71.676
R774 B.n516 B.n515 71.676
R775 B.n355 B.n354 71.676
R776 B.n361 B.n360 71.676
R777 B.n362 B.n351 71.676
R778 B.n369 B.n368 71.676
R779 B.n370 B.n349 71.676
R780 B.n377 B.n376 71.676
R781 B.n378 B.n347 71.676
R782 B.n385 B.n384 71.676
R783 B.n386 B.n345 71.676
R784 B.n393 B.n392 71.676
R785 B.n394 B.n343 71.676
R786 B.n401 B.n400 71.676
R787 B.n402 B.n341 71.676
R788 B.n409 B.n408 71.676
R789 B.n410 B.n339 71.676
R790 B.n417 B.n416 71.676
R791 B.n418 B.n337 71.676
R792 B.n425 B.n424 71.676
R793 B.n426 B.n332 71.676
R794 B.n433 B.n432 71.676
R795 B.n434 B.n330 71.676
R796 B.n441 B.n440 71.676
R797 B.n442 B.n326 71.676
R798 B.n450 B.n449 71.676
R799 B.n451 B.n324 71.676
R800 B.n458 B.n457 71.676
R801 B.n459 B.n322 71.676
R802 B.n466 B.n465 71.676
R803 B.n467 B.n320 71.676
R804 B.n474 B.n473 71.676
R805 B.n475 B.n318 71.676
R806 B.n482 B.n481 71.676
R807 B.n483 B.n316 71.676
R808 B.n490 B.n489 71.676
R809 B.n491 B.n314 71.676
R810 B.n498 B.n497 71.676
R811 B.n499 B.n312 71.676
R812 B.n506 B.n505 71.676
R813 B.n507 B.n310 71.676
R814 B.n514 B.n513 71.676
R815 B.n517 B.n516 71.676
R816 B.n681 B.n680 71.676
R817 B.n681 B.n2 71.676
R818 B.n167 B.n94 59.5399
R819 B.n188 B.n92 59.5399
R820 B.n446 B.n328 59.5399
R821 B.n335 B.n334 59.5399
R822 B.n94 B.n93 54.6914
R823 B.n92 B.n91 54.6914
R824 B.n328 B.n327 54.6914
R825 B.n334 B.n333 54.6914
R826 B.n522 B.n302 47.2675
R827 B.n528 B.n302 47.2675
R828 B.n528 B.n298 47.2675
R829 B.n534 B.n298 47.2675
R830 B.n534 B.n293 47.2675
R831 B.n540 B.n293 47.2675
R832 B.n540 B.n294 47.2675
R833 B.n546 B.n286 47.2675
R834 B.n552 B.n286 47.2675
R835 B.n552 B.n282 47.2675
R836 B.n558 B.n282 47.2675
R837 B.n558 B.n278 47.2675
R838 B.n564 B.n278 47.2675
R839 B.n564 B.n274 47.2675
R840 B.n570 B.n274 47.2675
R841 B.n570 B.n270 47.2675
R842 B.n576 B.n270 47.2675
R843 B.n583 B.n266 47.2675
R844 B.n583 B.n262 47.2675
R845 B.n589 B.n262 47.2675
R846 B.n589 B.n4 47.2675
R847 B.n679 B.n4 47.2675
R848 B.n679 B.n678 47.2675
R849 B.n678 B.n677 47.2675
R850 B.n677 B.n8 47.2675
R851 B.n12 B.n8 47.2675
R852 B.n670 B.n12 47.2675
R853 B.n670 B.n669 47.2675
R854 B.n668 B.n16 47.2675
R855 B.n662 B.n16 47.2675
R856 B.n662 B.n661 47.2675
R857 B.n661 B.n660 47.2675
R858 B.n660 B.n23 47.2675
R859 B.n654 B.n23 47.2675
R860 B.n654 B.n653 47.2675
R861 B.n653 B.n652 47.2675
R862 B.n652 B.n30 47.2675
R863 B.n646 B.n30 47.2675
R864 B.n645 B.n644 47.2675
R865 B.n644 B.n37 47.2675
R866 B.n638 B.n37 47.2675
R867 B.n638 B.n637 47.2675
R868 B.n637 B.n636 47.2675
R869 B.n636 B.n44 47.2675
R870 B.n630 B.n44 47.2675
R871 B.n524 B.n304 36.059
R872 B.n520 B.n519 36.059
R873 B.n626 B.n625 36.059
R874 B.n632 B.n46 36.059
R875 B.n546 B.t7 35.4507
R876 B.n576 B.t1 35.4507
R877 B.t0 B.n668 35.4507
R878 B.n646 B.t3 35.4507
R879 B B.n682 18.0485
R880 B.n294 B.t7 11.8172
R881 B.t1 B.n266 11.8172
R882 B.n669 B.t0 11.8172
R883 B.t3 B.n645 11.8172
R884 B.n525 B.n524 10.6151
R885 B.n526 B.n525 10.6151
R886 B.n526 B.n296 10.6151
R887 B.n536 B.n296 10.6151
R888 B.n537 B.n536 10.6151
R889 B.n538 B.n537 10.6151
R890 B.n538 B.n288 10.6151
R891 B.n548 B.n288 10.6151
R892 B.n549 B.n548 10.6151
R893 B.n550 B.n549 10.6151
R894 B.n550 B.n280 10.6151
R895 B.n560 B.n280 10.6151
R896 B.n561 B.n560 10.6151
R897 B.n562 B.n561 10.6151
R898 B.n562 B.n272 10.6151
R899 B.n572 B.n272 10.6151
R900 B.n573 B.n572 10.6151
R901 B.n574 B.n573 10.6151
R902 B.n574 B.n264 10.6151
R903 B.n585 B.n264 10.6151
R904 B.n586 B.n585 10.6151
R905 B.n587 B.n586 10.6151
R906 B.n587 B.n0 10.6151
R907 B.n356 B.n304 10.6151
R908 B.n357 B.n356 10.6151
R909 B.n358 B.n357 10.6151
R910 B.n358 B.n352 10.6151
R911 B.n364 B.n352 10.6151
R912 B.n365 B.n364 10.6151
R913 B.n366 B.n365 10.6151
R914 B.n366 B.n350 10.6151
R915 B.n372 B.n350 10.6151
R916 B.n373 B.n372 10.6151
R917 B.n374 B.n373 10.6151
R918 B.n374 B.n348 10.6151
R919 B.n380 B.n348 10.6151
R920 B.n381 B.n380 10.6151
R921 B.n382 B.n381 10.6151
R922 B.n382 B.n346 10.6151
R923 B.n388 B.n346 10.6151
R924 B.n389 B.n388 10.6151
R925 B.n390 B.n389 10.6151
R926 B.n390 B.n344 10.6151
R927 B.n396 B.n344 10.6151
R928 B.n397 B.n396 10.6151
R929 B.n398 B.n397 10.6151
R930 B.n398 B.n342 10.6151
R931 B.n404 B.n342 10.6151
R932 B.n405 B.n404 10.6151
R933 B.n406 B.n405 10.6151
R934 B.n406 B.n340 10.6151
R935 B.n412 B.n340 10.6151
R936 B.n413 B.n412 10.6151
R937 B.n414 B.n413 10.6151
R938 B.n414 B.n338 10.6151
R939 B.n420 B.n338 10.6151
R940 B.n421 B.n420 10.6151
R941 B.n422 B.n421 10.6151
R942 B.n422 B.n336 10.6151
R943 B.n429 B.n428 10.6151
R944 B.n430 B.n429 10.6151
R945 B.n430 B.n331 10.6151
R946 B.n436 B.n331 10.6151
R947 B.n437 B.n436 10.6151
R948 B.n438 B.n437 10.6151
R949 B.n438 B.n329 10.6151
R950 B.n444 B.n329 10.6151
R951 B.n445 B.n444 10.6151
R952 B.n447 B.n325 10.6151
R953 B.n453 B.n325 10.6151
R954 B.n454 B.n453 10.6151
R955 B.n455 B.n454 10.6151
R956 B.n455 B.n323 10.6151
R957 B.n461 B.n323 10.6151
R958 B.n462 B.n461 10.6151
R959 B.n463 B.n462 10.6151
R960 B.n463 B.n321 10.6151
R961 B.n469 B.n321 10.6151
R962 B.n470 B.n469 10.6151
R963 B.n471 B.n470 10.6151
R964 B.n471 B.n319 10.6151
R965 B.n477 B.n319 10.6151
R966 B.n478 B.n477 10.6151
R967 B.n479 B.n478 10.6151
R968 B.n479 B.n317 10.6151
R969 B.n485 B.n317 10.6151
R970 B.n486 B.n485 10.6151
R971 B.n487 B.n486 10.6151
R972 B.n487 B.n315 10.6151
R973 B.n493 B.n315 10.6151
R974 B.n494 B.n493 10.6151
R975 B.n495 B.n494 10.6151
R976 B.n495 B.n313 10.6151
R977 B.n501 B.n313 10.6151
R978 B.n502 B.n501 10.6151
R979 B.n503 B.n502 10.6151
R980 B.n503 B.n311 10.6151
R981 B.n509 B.n311 10.6151
R982 B.n510 B.n509 10.6151
R983 B.n511 B.n510 10.6151
R984 B.n511 B.n309 10.6151
R985 B.n309 B.n308 10.6151
R986 B.n518 B.n308 10.6151
R987 B.n519 B.n518 10.6151
R988 B.n520 B.n300 10.6151
R989 B.n530 B.n300 10.6151
R990 B.n531 B.n530 10.6151
R991 B.n532 B.n531 10.6151
R992 B.n532 B.n291 10.6151
R993 B.n542 B.n291 10.6151
R994 B.n543 B.n542 10.6151
R995 B.n544 B.n543 10.6151
R996 B.n544 B.n284 10.6151
R997 B.n554 B.n284 10.6151
R998 B.n555 B.n554 10.6151
R999 B.n556 B.n555 10.6151
R1000 B.n556 B.n276 10.6151
R1001 B.n566 B.n276 10.6151
R1002 B.n567 B.n566 10.6151
R1003 B.n568 B.n567 10.6151
R1004 B.n568 B.n268 10.6151
R1005 B.n578 B.n268 10.6151
R1006 B.n579 B.n578 10.6151
R1007 B.n581 B.n579 10.6151
R1008 B.n581 B.n580 10.6151
R1009 B.n580 B.n260 10.6151
R1010 B.n592 B.n260 10.6151
R1011 B.n593 B.n592 10.6151
R1012 B.n594 B.n593 10.6151
R1013 B.n595 B.n594 10.6151
R1014 B.n596 B.n595 10.6151
R1015 B.n599 B.n596 10.6151
R1016 B.n600 B.n599 10.6151
R1017 B.n601 B.n600 10.6151
R1018 B.n602 B.n601 10.6151
R1019 B.n604 B.n602 10.6151
R1020 B.n605 B.n604 10.6151
R1021 B.n606 B.n605 10.6151
R1022 B.n607 B.n606 10.6151
R1023 B.n609 B.n607 10.6151
R1024 B.n610 B.n609 10.6151
R1025 B.n611 B.n610 10.6151
R1026 B.n612 B.n611 10.6151
R1027 B.n614 B.n612 10.6151
R1028 B.n615 B.n614 10.6151
R1029 B.n616 B.n615 10.6151
R1030 B.n617 B.n616 10.6151
R1031 B.n619 B.n617 10.6151
R1032 B.n620 B.n619 10.6151
R1033 B.n621 B.n620 10.6151
R1034 B.n622 B.n621 10.6151
R1035 B.n624 B.n622 10.6151
R1036 B.n625 B.n624 10.6151
R1037 B.n674 B.n1 10.6151
R1038 B.n674 B.n673 10.6151
R1039 B.n673 B.n672 10.6151
R1040 B.n672 B.n10 10.6151
R1041 B.n666 B.n10 10.6151
R1042 B.n666 B.n665 10.6151
R1043 B.n665 B.n664 10.6151
R1044 B.n664 B.n18 10.6151
R1045 B.n658 B.n18 10.6151
R1046 B.n658 B.n657 10.6151
R1047 B.n657 B.n656 10.6151
R1048 B.n656 B.n25 10.6151
R1049 B.n650 B.n25 10.6151
R1050 B.n650 B.n649 10.6151
R1051 B.n649 B.n648 10.6151
R1052 B.n648 B.n32 10.6151
R1053 B.n642 B.n32 10.6151
R1054 B.n642 B.n641 10.6151
R1055 B.n641 B.n640 10.6151
R1056 B.n640 B.n39 10.6151
R1057 B.n634 B.n39 10.6151
R1058 B.n634 B.n633 10.6151
R1059 B.n633 B.n632 10.6151
R1060 B.n95 B.n46 10.6151
R1061 B.n98 B.n95 10.6151
R1062 B.n99 B.n98 10.6151
R1063 B.n102 B.n99 10.6151
R1064 B.n103 B.n102 10.6151
R1065 B.n106 B.n103 10.6151
R1066 B.n107 B.n106 10.6151
R1067 B.n110 B.n107 10.6151
R1068 B.n111 B.n110 10.6151
R1069 B.n114 B.n111 10.6151
R1070 B.n115 B.n114 10.6151
R1071 B.n118 B.n115 10.6151
R1072 B.n119 B.n118 10.6151
R1073 B.n122 B.n119 10.6151
R1074 B.n123 B.n122 10.6151
R1075 B.n126 B.n123 10.6151
R1076 B.n127 B.n126 10.6151
R1077 B.n130 B.n127 10.6151
R1078 B.n131 B.n130 10.6151
R1079 B.n134 B.n131 10.6151
R1080 B.n135 B.n134 10.6151
R1081 B.n138 B.n135 10.6151
R1082 B.n139 B.n138 10.6151
R1083 B.n142 B.n139 10.6151
R1084 B.n143 B.n142 10.6151
R1085 B.n146 B.n143 10.6151
R1086 B.n147 B.n146 10.6151
R1087 B.n150 B.n147 10.6151
R1088 B.n151 B.n150 10.6151
R1089 B.n154 B.n151 10.6151
R1090 B.n155 B.n154 10.6151
R1091 B.n158 B.n155 10.6151
R1092 B.n159 B.n158 10.6151
R1093 B.n162 B.n159 10.6151
R1094 B.n163 B.n162 10.6151
R1095 B.n166 B.n163 10.6151
R1096 B.n171 B.n168 10.6151
R1097 B.n172 B.n171 10.6151
R1098 B.n175 B.n172 10.6151
R1099 B.n176 B.n175 10.6151
R1100 B.n179 B.n176 10.6151
R1101 B.n180 B.n179 10.6151
R1102 B.n183 B.n180 10.6151
R1103 B.n184 B.n183 10.6151
R1104 B.n187 B.n184 10.6151
R1105 B.n192 B.n189 10.6151
R1106 B.n193 B.n192 10.6151
R1107 B.n196 B.n193 10.6151
R1108 B.n197 B.n196 10.6151
R1109 B.n200 B.n197 10.6151
R1110 B.n201 B.n200 10.6151
R1111 B.n204 B.n201 10.6151
R1112 B.n205 B.n204 10.6151
R1113 B.n208 B.n205 10.6151
R1114 B.n209 B.n208 10.6151
R1115 B.n212 B.n209 10.6151
R1116 B.n213 B.n212 10.6151
R1117 B.n216 B.n213 10.6151
R1118 B.n217 B.n216 10.6151
R1119 B.n220 B.n217 10.6151
R1120 B.n221 B.n220 10.6151
R1121 B.n224 B.n221 10.6151
R1122 B.n225 B.n224 10.6151
R1123 B.n228 B.n225 10.6151
R1124 B.n229 B.n228 10.6151
R1125 B.n232 B.n229 10.6151
R1126 B.n233 B.n232 10.6151
R1127 B.n236 B.n233 10.6151
R1128 B.n237 B.n236 10.6151
R1129 B.n240 B.n237 10.6151
R1130 B.n241 B.n240 10.6151
R1131 B.n244 B.n241 10.6151
R1132 B.n245 B.n244 10.6151
R1133 B.n248 B.n245 10.6151
R1134 B.n249 B.n248 10.6151
R1135 B.n252 B.n249 10.6151
R1136 B.n253 B.n252 10.6151
R1137 B.n256 B.n253 10.6151
R1138 B.n258 B.n256 10.6151
R1139 B.n259 B.n258 10.6151
R1140 B.n626 B.n259 10.6151
R1141 B.n336 B.n335 9.36635
R1142 B.n447 B.n446 9.36635
R1143 B.n167 B.n166 9.36635
R1144 B.n189 B.n188 9.36635
R1145 B.n682 B.n0 8.11757
R1146 B.n682 B.n1 8.11757
R1147 B.n428 B.n335 1.24928
R1148 B.n446 B.n445 1.24928
R1149 B.n168 B.n167 1.24928
R1150 B.n188 B.n187 1.24928
R1151 VP.n0 VP.t1 194.548
R1152 VP.n0 VP.t0 151.281
R1153 VP VP.n0 0.336784
R1154 VTAIL.n230 VTAIL.n229 289.615
R1155 VTAIL.n56 VTAIL.n55 289.615
R1156 VTAIL.n172 VTAIL.n171 289.615
R1157 VTAIL.n114 VTAIL.n113 289.615
R1158 VTAIL.n192 VTAIL.n191 185
R1159 VTAIL.n197 VTAIL.n196 185
R1160 VTAIL.n199 VTAIL.n198 185
R1161 VTAIL.n188 VTAIL.n187 185
R1162 VTAIL.n205 VTAIL.n204 185
R1163 VTAIL.n207 VTAIL.n206 185
R1164 VTAIL.n184 VTAIL.n183 185
R1165 VTAIL.n213 VTAIL.n212 185
R1166 VTAIL.n215 VTAIL.n214 185
R1167 VTAIL.n180 VTAIL.n179 185
R1168 VTAIL.n221 VTAIL.n220 185
R1169 VTAIL.n223 VTAIL.n222 185
R1170 VTAIL.n176 VTAIL.n175 185
R1171 VTAIL.n229 VTAIL.n228 185
R1172 VTAIL.n18 VTAIL.n17 185
R1173 VTAIL.n23 VTAIL.n22 185
R1174 VTAIL.n25 VTAIL.n24 185
R1175 VTAIL.n14 VTAIL.n13 185
R1176 VTAIL.n31 VTAIL.n30 185
R1177 VTAIL.n33 VTAIL.n32 185
R1178 VTAIL.n10 VTAIL.n9 185
R1179 VTAIL.n39 VTAIL.n38 185
R1180 VTAIL.n41 VTAIL.n40 185
R1181 VTAIL.n6 VTAIL.n5 185
R1182 VTAIL.n47 VTAIL.n46 185
R1183 VTAIL.n49 VTAIL.n48 185
R1184 VTAIL.n2 VTAIL.n1 185
R1185 VTAIL.n55 VTAIL.n54 185
R1186 VTAIL.n171 VTAIL.n170 185
R1187 VTAIL.n118 VTAIL.n117 185
R1188 VTAIL.n165 VTAIL.n164 185
R1189 VTAIL.n163 VTAIL.n162 185
R1190 VTAIL.n122 VTAIL.n121 185
R1191 VTAIL.n157 VTAIL.n156 185
R1192 VTAIL.n155 VTAIL.n154 185
R1193 VTAIL.n126 VTAIL.n125 185
R1194 VTAIL.n149 VTAIL.n148 185
R1195 VTAIL.n147 VTAIL.n146 185
R1196 VTAIL.n130 VTAIL.n129 185
R1197 VTAIL.n141 VTAIL.n140 185
R1198 VTAIL.n139 VTAIL.n138 185
R1199 VTAIL.n134 VTAIL.n133 185
R1200 VTAIL.n113 VTAIL.n112 185
R1201 VTAIL.n60 VTAIL.n59 185
R1202 VTAIL.n107 VTAIL.n106 185
R1203 VTAIL.n105 VTAIL.n104 185
R1204 VTAIL.n64 VTAIL.n63 185
R1205 VTAIL.n99 VTAIL.n98 185
R1206 VTAIL.n97 VTAIL.n96 185
R1207 VTAIL.n68 VTAIL.n67 185
R1208 VTAIL.n91 VTAIL.n90 185
R1209 VTAIL.n89 VTAIL.n88 185
R1210 VTAIL.n72 VTAIL.n71 185
R1211 VTAIL.n83 VTAIL.n82 185
R1212 VTAIL.n81 VTAIL.n80 185
R1213 VTAIL.n76 VTAIL.n75 185
R1214 VTAIL.n193 VTAIL.t1 147.659
R1215 VTAIL.n19 VTAIL.t2 147.659
R1216 VTAIL.n135 VTAIL.t3 147.659
R1217 VTAIL.n77 VTAIL.t0 147.659
R1218 VTAIL.n197 VTAIL.n191 104.615
R1219 VTAIL.n198 VTAIL.n197 104.615
R1220 VTAIL.n198 VTAIL.n187 104.615
R1221 VTAIL.n205 VTAIL.n187 104.615
R1222 VTAIL.n206 VTAIL.n205 104.615
R1223 VTAIL.n206 VTAIL.n183 104.615
R1224 VTAIL.n213 VTAIL.n183 104.615
R1225 VTAIL.n214 VTAIL.n213 104.615
R1226 VTAIL.n214 VTAIL.n179 104.615
R1227 VTAIL.n221 VTAIL.n179 104.615
R1228 VTAIL.n222 VTAIL.n221 104.615
R1229 VTAIL.n222 VTAIL.n175 104.615
R1230 VTAIL.n229 VTAIL.n175 104.615
R1231 VTAIL.n23 VTAIL.n17 104.615
R1232 VTAIL.n24 VTAIL.n23 104.615
R1233 VTAIL.n24 VTAIL.n13 104.615
R1234 VTAIL.n31 VTAIL.n13 104.615
R1235 VTAIL.n32 VTAIL.n31 104.615
R1236 VTAIL.n32 VTAIL.n9 104.615
R1237 VTAIL.n39 VTAIL.n9 104.615
R1238 VTAIL.n40 VTAIL.n39 104.615
R1239 VTAIL.n40 VTAIL.n5 104.615
R1240 VTAIL.n47 VTAIL.n5 104.615
R1241 VTAIL.n48 VTAIL.n47 104.615
R1242 VTAIL.n48 VTAIL.n1 104.615
R1243 VTAIL.n55 VTAIL.n1 104.615
R1244 VTAIL.n171 VTAIL.n117 104.615
R1245 VTAIL.n164 VTAIL.n117 104.615
R1246 VTAIL.n164 VTAIL.n163 104.615
R1247 VTAIL.n163 VTAIL.n121 104.615
R1248 VTAIL.n156 VTAIL.n121 104.615
R1249 VTAIL.n156 VTAIL.n155 104.615
R1250 VTAIL.n155 VTAIL.n125 104.615
R1251 VTAIL.n148 VTAIL.n125 104.615
R1252 VTAIL.n148 VTAIL.n147 104.615
R1253 VTAIL.n147 VTAIL.n129 104.615
R1254 VTAIL.n140 VTAIL.n129 104.615
R1255 VTAIL.n140 VTAIL.n139 104.615
R1256 VTAIL.n139 VTAIL.n133 104.615
R1257 VTAIL.n113 VTAIL.n59 104.615
R1258 VTAIL.n106 VTAIL.n59 104.615
R1259 VTAIL.n106 VTAIL.n105 104.615
R1260 VTAIL.n105 VTAIL.n63 104.615
R1261 VTAIL.n98 VTAIL.n63 104.615
R1262 VTAIL.n98 VTAIL.n97 104.615
R1263 VTAIL.n97 VTAIL.n67 104.615
R1264 VTAIL.n90 VTAIL.n67 104.615
R1265 VTAIL.n90 VTAIL.n89 104.615
R1266 VTAIL.n89 VTAIL.n71 104.615
R1267 VTAIL.n82 VTAIL.n71 104.615
R1268 VTAIL.n82 VTAIL.n81 104.615
R1269 VTAIL.n81 VTAIL.n75 104.615
R1270 VTAIL.t1 VTAIL.n191 52.3082
R1271 VTAIL.t2 VTAIL.n17 52.3082
R1272 VTAIL.t3 VTAIL.n133 52.3082
R1273 VTAIL.t0 VTAIL.n75 52.3082
R1274 VTAIL.n231 VTAIL.n230 33.9308
R1275 VTAIL.n57 VTAIL.n56 33.9308
R1276 VTAIL.n173 VTAIL.n172 33.9308
R1277 VTAIL.n115 VTAIL.n114 33.9308
R1278 VTAIL.n115 VTAIL.n57 26.3238
R1279 VTAIL.n231 VTAIL.n173 23.8927
R1280 VTAIL.n193 VTAIL.n192 15.6677
R1281 VTAIL.n19 VTAIL.n18 15.6677
R1282 VTAIL.n135 VTAIL.n134 15.6677
R1283 VTAIL.n77 VTAIL.n76 15.6677
R1284 VTAIL.n196 VTAIL.n195 12.8005
R1285 VTAIL.n22 VTAIL.n21 12.8005
R1286 VTAIL.n138 VTAIL.n137 12.8005
R1287 VTAIL.n80 VTAIL.n79 12.8005
R1288 VTAIL.n199 VTAIL.n190 12.0247
R1289 VTAIL.n25 VTAIL.n16 12.0247
R1290 VTAIL.n141 VTAIL.n132 12.0247
R1291 VTAIL.n83 VTAIL.n74 12.0247
R1292 VTAIL.n200 VTAIL.n188 11.249
R1293 VTAIL.n26 VTAIL.n14 11.249
R1294 VTAIL.n142 VTAIL.n130 11.249
R1295 VTAIL.n84 VTAIL.n72 11.249
R1296 VTAIL.n204 VTAIL.n203 10.4732
R1297 VTAIL.n228 VTAIL.n174 10.4732
R1298 VTAIL.n30 VTAIL.n29 10.4732
R1299 VTAIL.n54 VTAIL.n0 10.4732
R1300 VTAIL.n170 VTAIL.n116 10.4732
R1301 VTAIL.n146 VTAIL.n145 10.4732
R1302 VTAIL.n112 VTAIL.n58 10.4732
R1303 VTAIL.n88 VTAIL.n87 10.4732
R1304 VTAIL.n207 VTAIL.n186 9.69747
R1305 VTAIL.n227 VTAIL.n176 9.69747
R1306 VTAIL.n33 VTAIL.n12 9.69747
R1307 VTAIL.n53 VTAIL.n2 9.69747
R1308 VTAIL.n169 VTAIL.n118 9.69747
R1309 VTAIL.n149 VTAIL.n128 9.69747
R1310 VTAIL.n111 VTAIL.n60 9.69747
R1311 VTAIL.n91 VTAIL.n70 9.69747
R1312 VTAIL.n226 VTAIL.n174 9.45567
R1313 VTAIL.n52 VTAIL.n0 9.45567
R1314 VTAIL.n168 VTAIL.n116 9.45567
R1315 VTAIL.n110 VTAIL.n58 9.45567
R1316 VTAIL.n217 VTAIL.n216 9.3005
R1317 VTAIL.n219 VTAIL.n218 9.3005
R1318 VTAIL.n178 VTAIL.n177 9.3005
R1319 VTAIL.n225 VTAIL.n224 9.3005
R1320 VTAIL.n227 VTAIL.n226 9.3005
R1321 VTAIL.n211 VTAIL.n210 9.3005
R1322 VTAIL.n209 VTAIL.n208 9.3005
R1323 VTAIL.n186 VTAIL.n185 9.3005
R1324 VTAIL.n203 VTAIL.n202 9.3005
R1325 VTAIL.n201 VTAIL.n200 9.3005
R1326 VTAIL.n190 VTAIL.n189 9.3005
R1327 VTAIL.n195 VTAIL.n194 9.3005
R1328 VTAIL.n182 VTAIL.n181 9.3005
R1329 VTAIL.n43 VTAIL.n42 9.3005
R1330 VTAIL.n45 VTAIL.n44 9.3005
R1331 VTAIL.n4 VTAIL.n3 9.3005
R1332 VTAIL.n51 VTAIL.n50 9.3005
R1333 VTAIL.n53 VTAIL.n52 9.3005
R1334 VTAIL.n37 VTAIL.n36 9.3005
R1335 VTAIL.n35 VTAIL.n34 9.3005
R1336 VTAIL.n12 VTAIL.n11 9.3005
R1337 VTAIL.n29 VTAIL.n28 9.3005
R1338 VTAIL.n27 VTAIL.n26 9.3005
R1339 VTAIL.n16 VTAIL.n15 9.3005
R1340 VTAIL.n21 VTAIL.n20 9.3005
R1341 VTAIL.n8 VTAIL.n7 9.3005
R1342 VTAIL.n169 VTAIL.n168 9.3005
R1343 VTAIL.n167 VTAIL.n166 9.3005
R1344 VTAIL.n120 VTAIL.n119 9.3005
R1345 VTAIL.n161 VTAIL.n160 9.3005
R1346 VTAIL.n159 VTAIL.n158 9.3005
R1347 VTAIL.n124 VTAIL.n123 9.3005
R1348 VTAIL.n153 VTAIL.n152 9.3005
R1349 VTAIL.n151 VTAIL.n150 9.3005
R1350 VTAIL.n128 VTAIL.n127 9.3005
R1351 VTAIL.n145 VTAIL.n144 9.3005
R1352 VTAIL.n143 VTAIL.n142 9.3005
R1353 VTAIL.n132 VTAIL.n131 9.3005
R1354 VTAIL.n137 VTAIL.n136 9.3005
R1355 VTAIL.n103 VTAIL.n102 9.3005
R1356 VTAIL.n62 VTAIL.n61 9.3005
R1357 VTAIL.n109 VTAIL.n108 9.3005
R1358 VTAIL.n111 VTAIL.n110 9.3005
R1359 VTAIL.n101 VTAIL.n100 9.3005
R1360 VTAIL.n66 VTAIL.n65 9.3005
R1361 VTAIL.n95 VTAIL.n94 9.3005
R1362 VTAIL.n93 VTAIL.n92 9.3005
R1363 VTAIL.n70 VTAIL.n69 9.3005
R1364 VTAIL.n87 VTAIL.n86 9.3005
R1365 VTAIL.n85 VTAIL.n84 9.3005
R1366 VTAIL.n74 VTAIL.n73 9.3005
R1367 VTAIL.n79 VTAIL.n78 9.3005
R1368 VTAIL.n208 VTAIL.n184 8.92171
R1369 VTAIL.n224 VTAIL.n223 8.92171
R1370 VTAIL.n34 VTAIL.n10 8.92171
R1371 VTAIL.n50 VTAIL.n49 8.92171
R1372 VTAIL.n166 VTAIL.n165 8.92171
R1373 VTAIL.n150 VTAIL.n126 8.92171
R1374 VTAIL.n108 VTAIL.n107 8.92171
R1375 VTAIL.n92 VTAIL.n68 8.92171
R1376 VTAIL.n212 VTAIL.n211 8.14595
R1377 VTAIL.n220 VTAIL.n178 8.14595
R1378 VTAIL.n38 VTAIL.n37 8.14595
R1379 VTAIL.n46 VTAIL.n4 8.14595
R1380 VTAIL.n162 VTAIL.n120 8.14595
R1381 VTAIL.n154 VTAIL.n153 8.14595
R1382 VTAIL.n104 VTAIL.n62 8.14595
R1383 VTAIL.n96 VTAIL.n95 8.14595
R1384 VTAIL.n215 VTAIL.n182 7.3702
R1385 VTAIL.n219 VTAIL.n180 7.3702
R1386 VTAIL.n41 VTAIL.n8 7.3702
R1387 VTAIL.n45 VTAIL.n6 7.3702
R1388 VTAIL.n161 VTAIL.n122 7.3702
R1389 VTAIL.n157 VTAIL.n124 7.3702
R1390 VTAIL.n103 VTAIL.n64 7.3702
R1391 VTAIL.n99 VTAIL.n66 7.3702
R1392 VTAIL.n216 VTAIL.n215 6.59444
R1393 VTAIL.n216 VTAIL.n180 6.59444
R1394 VTAIL.n42 VTAIL.n41 6.59444
R1395 VTAIL.n42 VTAIL.n6 6.59444
R1396 VTAIL.n158 VTAIL.n122 6.59444
R1397 VTAIL.n158 VTAIL.n157 6.59444
R1398 VTAIL.n100 VTAIL.n64 6.59444
R1399 VTAIL.n100 VTAIL.n99 6.59444
R1400 VTAIL.n212 VTAIL.n182 5.81868
R1401 VTAIL.n220 VTAIL.n219 5.81868
R1402 VTAIL.n38 VTAIL.n8 5.81868
R1403 VTAIL.n46 VTAIL.n45 5.81868
R1404 VTAIL.n162 VTAIL.n161 5.81868
R1405 VTAIL.n154 VTAIL.n124 5.81868
R1406 VTAIL.n104 VTAIL.n103 5.81868
R1407 VTAIL.n96 VTAIL.n66 5.81868
R1408 VTAIL.n211 VTAIL.n184 5.04292
R1409 VTAIL.n223 VTAIL.n178 5.04292
R1410 VTAIL.n37 VTAIL.n10 5.04292
R1411 VTAIL.n49 VTAIL.n4 5.04292
R1412 VTAIL.n165 VTAIL.n120 5.04292
R1413 VTAIL.n153 VTAIL.n126 5.04292
R1414 VTAIL.n107 VTAIL.n62 5.04292
R1415 VTAIL.n95 VTAIL.n68 5.04292
R1416 VTAIL.n194 VTAIL.n193 4.38563
R1417 VTAIL.n20 VTAIL.n19 4.38563
R1418 VTAIL.n136 VTAIL.n135 4.38563
R1419 VTAIL.n78 VTAIL.n77 4.38563
R1420 VTAIL.n208 VTAIL.n207 4.26717
R1421 VTAIL.n224 VTAIL.n176 4.26717
R1422 VTAIL.n34 VTAIL.n33 4.26717
R1423 VTAIL.n50 VTAIL.n2 4.26717
R1424 VTAIL.n166 VTAIL.n118 4.26717
R1425 VTAIL.n150 VTAIL.n149 4.26717
R1426 VTAIL.n108 VTAIL.n60 4.26717
R1427 VTAIL.n92 VTAIL.n91 4.26717
R1428 VTAIL.n204 VTAIL.n186 3.49141
R1429 VTAIL.n228 VTAIL.n227 3.49141
R1430 VTAIL.n30 VTAIL.n12 3.49141
R1431 VTAIL.n54 VTAIL.n53 3.49141
R1432 VTAIL.n170 VTAIL.n169 3.49141
R1433 VTAIL.n146 VTAIL.n128 3.49141
R1434 VTAIL.n112 VTAIL.n111 3.49141
R1435 VTAIL.n88 VTAIL.n70 3.49141
R1436 VTAIL.n203 VTAIL.n188 2.71565
R1437 VTAIL.n230 VTAIL.n174 2.71565
R1438 VTAIL.n29 VTAIL.n14 2.71565
R1439 VTAIL.n56 VTAIL.n0 2.71565
R1440 VTAIL.n172 VTAIL.n116 2.71565
R1441 VTAIL.n145 VTAIL.n130 2.71565
R1442 VTAIL.n114 VTAIL.n58 2.71565
R1443 VTAIL.n87 VTAIL.n72 2.71565
R1444 VTAIL.n200 VTAIL.n199 1.93989
R1445 VTAIL.n26 VTAIL.n25 1.93989
R1446 VTAIL.n142 VTAIL.n141 1.93989
R1447 VTAIL.n84 VTAIL.n83 1.93989
R1448 VTAIL.n173 VTAIL.n115 1.68584
R1449 VTAIL.n196 VTAIL.n190 1.16414
R1450 VTAIL.n22 VTAIL.n16 1.16414
R1451 VTAIL.n138 VTAIL.n132 1.16414
R1452 VTAIL.n80 VTAIL.n74 1.16414
R1453 VTAIL VTAIL.n57 1.13628
R1454 VTAIL VTAIL.n231 0.550069
R1455 VTAIL.n195 VTAIL.n192 0.388379
R1456 VTAIL.n21 VTAIL.n18 0.388379
R1457 VTAIL.n137 VTAIL.n134 0.388379
R1458 VTAIL.n79 VTAIL.n76 0.388379
R1459 VTAIL.n194 VTAIL.n189 0.155672
R1460 VTAIL.n201 VTAIL.n189 0.155672
R1461 VTAIL.n202 VTAIL.n201 0.155672
R1462 VTAIL.n202 VTAIL.n185 0.155672
R1463 VTAIL.n209 VTAIL.n185 0.155672
R1464 VTAIL.n210 VTAIL.n209 0.155672
R1465 VTAIL.n210 VTAIL.n181 0.155672
R1466 VTAIL.n217 VTAIL.n181 0.155672
R1467 VTAIL.n218 VTAIL.n217 0.155672
R1468 VTAIL.n218 VTAIL.n177 0.155672
R1469 VTAIL.n225 VTAIL.n177 0.155672
R1470 VTAIL.n226 VTAIL.n225 0.155672
R1471 VTAIL.n20 VTAIL.n15 0.155672
R1472 VTAIL.n27 VTAIL.n15 0.155672
R1473 VTAIL.n28 VTAIL.n27 0.155672
R1474 VTAIL.n28 VTAIL.n11 0.155672
R1475 VTAIL.n35 VTAIL.n11 0.155672
R1476 VTAIL.n36 VTAIL.n35 0.155672
R1477 VTAIL.n36 VTAIL.n7 0.155672
R1478 VTAIL.n43 VTAIL.n7 0.155672
R1479 VTAIL.n44 VTAIL.n43 0.155672
R1480 VTAIL.n44 VTAIL.n3 0.155672
R1481 VTAIL.n51 VTAIL.n3 0.155672
R1482 VTAIL.n52 VTAIL.n51 0.155672
R1483 VTAIL.n168 VTAIL.n167 0.155672
R1484 VTAIL.n167 VTAIL.n119 0.155672
R1485 VTAIL.n160 VTAIL.n119 0.155672
R1486 VTAIL.n160 VTAIL.n159 0.155672
R1487 VTAIL.n159 VTAIL.n123 0.155672
R1488 VTAIL.n152 VTAIL.n123 0.155672
R1489 VTAIL.n152 VTAIL.n151 0.155672
R1490 VTAIL.n151 VTAIL.n127 0.155672
R1491 VTAIL.n144 VTAIL.n127 0.155672
R1492 VTAIL.n144 VTAIL.n143 0.155672
R1493 VTAIL.n143 VTAIL.n131 0.155672
R1494 VTAIL.n136 VTAIL.n131 0.155672
R1495 VTAIL.n110 VTAIL.n109 0.155672
R1496 VTAIL.n109 VTAIL.n61 0.155672
R1497 VTAIL.n102 VTAIL.n61 0.155672
R1498 VTAIL.n102 VTAIL.n101 0.155672
R1499 VTAIL.n101 VTAIL.n65 0.155672
R1500 VTAIL.n94 VTAIL.n65 0.155672
R1501 VTAIL.n94 VTAIL.n93 0.155672
R1502 VTAIL.n93 VTAIL.n69 0.155672
R1503 VTAIL.n86 VTAIL.n69 0.155672
R1504 VTAIL.n86 VTAIL.n85 0.155672
R1505 VTAIL.n85 VTAIL.n73 0.155672
R1506 VTAIL.n78 VTAIL.n73 0.155672
R1507 VDD1.n56 VDD1.n55 289.615
R1508 VDD1.n113 VDD1.n112 289.615
R1509 VDD1.n55 VDD1.n54 185
R1510 VDD1.n2 VDD1.n1 185
R1511 VDD1.n49 VDD1.n48 185
R1512 VDD1.n47 VDD1.n46 185
R1513 VDD1.n6 VDD1.n5 185
R1514 VDD1.n41 VDD1.n40 185
R1515 VDD1.n39 VDD1.n38 185
R1516 VDD1.n10 VDD1.n9 185
R1517 VDD1.n33 VDD1.n32 185
R1518 VDD1.n31 VDD1.n30 185
R1519 VDD1.n14 VDD1.n13 185
R1520 VDD1.n25 VDD1.n24 185
R1521 VDD1.n23 VDD1.n22 185
R1522 VDD1.n18 VDD1.n17 185
R1523 VDD1.n75 VDD1.n74 185
R1524 VDD1.n80 VDD1.n79 185
R1525 VDD1.n82 VDD1.n81 185
R1526 VDD1.n71 VDD1.n70 185
R1527 VDD1.n88 VDD1.n87 185
R1528 VDD1.n90 VDD1.n89 185
R1529 VDD1.n67 VDD1.n66 185
R1530 VDD1.n96 VDD1.n95 185
R1531 VDD1.n98 VDD1.n97 185
R1532 VDD1.n63 VDD1.n62 185
R1533 VDD1.n104 VDD1.n103 185
R1534 VDD1.n106 VDD1.n105 185
R1535 VDD1.n59 VDD1.n58 185
R1536 VDD1.n112 VDD1.n111 185
R1537 VDD1.n76 VDD1.t1 147.659
R1538 VDD1.n19 VDD1.t0 147.659
R1539 VDD1.n55 VDD1.n1 104.615
R1540 VDD1.n48 VDD1.n1 104.615
R1541 VDD1.n48 VDD1.n47 104.615
R1542 VDD1.n47 VDD1.n5 104.615
R1543 VDD1.n40 VDD1.n5 104.615
R1544 VDD1.n40 VDD1.n39 104.615
R1545 VDD1.n39 VDD1.n9 104.615
R1546 VDD1.n32 VDD1.n9 104.615
R1547 VDD1.n32 VDD1.n31 104.615
R1548 VDD1.n31 VDD1.n13 104.615
R1549 VDD1.n24 VDD1.n13 104.615
R1550 VDD1.n24 VDD1.n23 104.615
R1551 VDD1.n23 VDD1.n17 104.615
R1552 VDD1.n80 VDD1.n74 104.615
R1553 VDD1.n81 VDD1.n80 104.615
R1554 VDD1.n81 VDD1.n70 104.615
R1555 VDD1.n88 VDD1.n70 104.615
R1556 VDD1.n89 VDD1.n88 104.615
R1557 VDD1.n89 VDD1.n66 104.615
R1558 VDD1.n96 VDD1.n66 104.615
R1559 VDD1.n97 VDD1.n96 104.615
R1560 VDD1.n97 VDD1.n62 104.615
R1561 VDD1.n104 VDD1.n62 104.615
R1562 VDD1.n105 VDD1.n104 104.615
R1563 VDD1.n105 VDD1.n58 104.615
R1564 VDD1.n112 VDD1.n58 104.615
R1565 VDD1 VDD1.n113 89.3585
R1566 VDD1.t0 VDD1.n17 52.3082
R1567 VDD1.t1 VDD1.n74 52.3082
R1568 VDD1 VDD1.n56 51.2755
R1569 VDD1.n19 VDD1.n18 15.6677
R1570 VDD1.n76 VDD1.n75 15.6677
R1571 VDD1.n22 VDD1.n21 12.8005
R1572 VDD1.n79 VDD1.n78 12.8005
R1573 VDD1.n25 VDD1.n16 12.0247
R1574 VDD1.n82 VDD1.n73 12.0247
R1575 VDD1.n26 VDD1.n14 11.249
R1576 VDD1.n83 VDD1.n71 11.249
R1577 VDD1.n54 VDD1.n0 10.4732
R1578 VDD1.n30 VDD1.n29 10.4732
R1579 VDD1.n87 VDD1.n86 10.4732
R1580 VDD1.n111 VDD1.n57 10.4732
R1581 VDD1.n53 VDD1.n2 9.69747
R1582 VDD1.n33 VDD1.n12 9.69747
R1583 VDD1.n90 VDD1.n69 9.69747
R1584 VDD1.n110 VDD1.n59 9.69747
R1585 VDD1.n52 VDD1.n0 9.45567
R1586 VDD1.n109 VDD1.n57 9.45567
R1587 VDD1.n53 VDD1.n52 9.3005
R1588 VDD1.n51 VDD1.n50 9.3005
R1589 VDD1.n4 VDD1.n3 9.3005
R1590 VDD1.n45 VDD1.n44 9.3005
R1591 VDD1.n43 VDD1.n42 9.3005
R1592 VDD1.n8 VDD1.n7 9.3005
R1593 VDD1.n37 VDD1.n36 9.3005
R1594 VDD1.n35 VDD1.n34 9.3005
R1595 VDD1.n12 VDD1.n11 9.3005
R1596 VDD1.n29 VDD1.n28 9.3005
R1597 VDD1.n27 VDD1.n26 9.3005
R1598 VDD1.n16 VDD1.n15 9.3005
R1599 VDD1.n21 VDD1.n20 9.3005
R1600 VDD1.n100 VDD1.n99 9.3005
R1601 VDD1.n102 VDD1.n101 9.3005
R1602 VDD1.n61 VDD1.n60 9.3005
R1603 VDD1.n108 VDD1.n107 9.3005
R1604 VDD1.n110 VDD1.n109 9.3005
R1605 VDD1.n94 VDD1.n93 9.3005
R1606 VDD1.n92 VDD1.n91 9.3005
R1607 VDD1.n69 VDD1.n68 9.3005
R1608 VDD1.n86 VDD1.n85 9.3005
R1609 VDD1.n84 VDD1.n83 9.3005
R1610 VDD1.n73 VDD1.n72 9.3005
R1611 VDD1.n78 VDD1.n77 9.3005
R1612 VDD1.n65 VDD1.n64 9.3005
R1613 VDD1.n50 VDD1.n49 8.92171
R1614 VDD1.n34 VDD1.n10 8.92171
R1615 VDD1.n91 VDD1.n67 8.92171
R1616 VDD1.n107 VDD1.n106 8.92171
R1617 VDD1.n46 VDD1.n4 8.14595
R1618 VDD1.n38 VDD1.n37 8.14595
R1619 VDD1.n95 VDD1.n94 8.14595
R1620 VDD1.n103 VDD1.n61 8.14595
R1621 VDD1.n45 VDD1.n6 7.3702
R1622 VDD1.n41 VDD1.n8 7.3702
R1623 VDD1.n98 VDD1.n65 7.3702
R1624 VDD1.n102 VDD1.n63 7.3702
R1625 VDD1.n42 VDD1.n6 6.59444
R1626 VDD1.n42 VDD1.n41 6.59444
R1627 VDD1.n99 VDD1.n98 6.59444
R1628 VDD1.n99 VDD1.n63 6.59444
R1629 VDD1.n46 VDD1.n45 5.81868
R1630 VDD1.n38 VDD1.n8 5.81868
R1631 VDD1.n95 VDD1.n65 5.81868
R1632 VDD1.n103 VDD1.n102 5.81868
R1633 VDD1.n49 VDD1.n4 5.04292
R1634 VDD1.n37 VDD1.n10 5.04292
R1635 VDD1.n94 VDD1.n67 5.04292
R1636 VDD1.n106 VDD1.n61 5.04292
R1637 VDD1.n77 VDD1.n76 4.38563
R1638 VDD1.n20 VDD1.n19 4.38563
R1639 VDD1.n50 VDD1.n2 4.26717
R1640 VDD1.n34 VDD1.n33 4.26717
R1641 VDD1.n91 VDD1.n90 4.26717
R1642 VDD1.n107 VDD1.n59 4.26717
R1643 VDD1.n54 VDD1.n53 3.49141
R1644 VDD1.n30 VDD1.n12 3.49141
R1645 VDD1.n87 VDD1.n69 3.49141
R1646 VDD1.n111 VDD1.n110 3.49141
R1647 VDD1.n56 VDD1.n0 2.71565
R1648 VDD1.n29 VDD1.n14 2.71565
R1649 VDD1.n86 VDD1.n71 2.71565
R1650 VDD1.n113 VDD1.n57 2.71565
R1651 VDD1.n26 VDD1.n25 1.93989
R1652 VDD1.n83 VDD1.n82 1.93989
R1653 VDD1.n22 VDD1.n16 1.16414
R1654 VDD1.n79 VDD1.n73 1.16414
R1655 VDD1.n21 VDD1.n18 0.388379
R1656 VDD1.n78 VDD1.n75 0.388379
R1657 VDD1.n52 VDD1.n51 0.155672
R1658 VDD1.n51 VDD1.n3 0.155672
R1659 VDD1.n44 VDD1.n3 0.155672
R1660 VDD1.n44 VDD1.n43 0.155672
R1661 VDD1.n43 VDD1.n7 0.155672
R1662 VDD1.n36 VDD1.n7 0.155672
R1663 VDD1.n36 VDD1.n35 0.155672
R1664 VDD1.n35 VDD1.n11 0.155672
R1665 VDD1.n28 VDD1.n11 0.155672
R1666 VDD1.n28 VDD1.n27 0.155672
R1667 VDD1.n27 VDD1.n15 0.155672
R1668 VDD1.n20 VDD1.n15 0.155672
R1669 VDD1.n77 VDD1.n72 0.155672
R1670 VDD1.n84 VDD1.n72 0.155672
R1671 VDD1.n85 VDD1.n84 0.155672
R1672 VDD1.n85 VDD1.n68 0.155672
R1673 VDD1.n92 VDD1.n68 0.155672
R1674 VDD1.n93 VDD1.n92 0.155672
R1675 VDD1.n93 VDD1.n64 0.155672
R1676 VDD1.n100 VDD1.n64 0.155672
R1677 VDD1.n101 VDD1.n100 0.155672
R1678 VDD1.n101 VDD1.n60 0.155672
R1679 VDD1.n108 VDD1.n60 0.155672
R1680 VDD1.n109 VDD1.n108 0.155672
R1681 VN VN.t0 194.644
R1682 VN VN.t1 151.618
R1683 VDD2.n113 VDD2.n112 289.615
R1684 VDD2.n56 VDD2.n55 289.615
R1685 VDD2.n112 VDD2.n111 185
R1686 VDD2.n59 VDD2.n58 185
R1687 VDD2.n106 VDD2.n105 185
R1688 VDD2.n104 VDD2.n103 185
R1689 VDD2.n63 VDD2.n62 185
R1690 VDD2.n98 VDD2.n97 185
R1691 VDD2.n96 VDD2.n95 185
R1692 VDD2.n67 VDD2.n66 185
R1693 VDD2.n90 VDD2.n89 185
R1694 VDD2.n88 VDD2.n87 185
R1695 VDD2.n71 VDD2.n70 185
R1696 VDD2.n82 VDD2.n81 185
R1697 VDD2.n80 VDD2.n79 185
R1698 VDD2.n75 VDD2.n74 185
R1699 VDD2.n18 VDD2.n17 185
R1700 VDD2.n23 VDD2.n22 185
R1701 VDD2.n25 VDD2.n24 185
R1702 VDD2.n14 VDD2.n13 185
R1703 VDD2.n31 VDD2.n30 185
R1704 VDD2.n33 VDD2.n32 185
R1705 VDD2.n10 VDD2.n9 185
R1706 VDD2.n39 VDD2.n38 185
R1707 VDD2.n41 VDD2.n40 185
R1708 VDD2.n6 VDD2.n5 185
R1709 VDD2.n47 VDD2.n46 185
R1710 VDD2.n49 VDD2.n48 185
R1711 VDD2.n2 VDD2.n1 185
R1712 VDD2.n55 VDD2.n54 185
R1713 VDD2.n19 VDD2.t0 147.659
R1714 VDD2.n76 VDD2.t1 147.659
R1715 VDD2.n112 VDD2.n58 104.615
R1716 VDD2.n105 VDD2.n58 104.615
R1717 VDD2.n105 VDD2.n104 104.615
R1718 VDD2.n104 VDD2.n62 104.615
R1719 VDD2.n97 VDD2.n62 104.615
R1720 VDD2.n97 VDD2.n96 104.615
R1721 VDD2.n96 VDD2.n66 104.615
R1722 VDD2.n89 VDD2.n66 104.615
R1723 VDD2.n89 VDD2.n88 104.615
R1724 VDD2.n88 VDD2.n70 104.615
R1725 VDD2.n81 VDD2.n70 104.615
R1726 VDD2.n81 VDD2.n80 104.615
R1727 VDD2.n80 VDD2.n74 104.615
R1728 VDD2.n23 VDD2.n17 104.615
R1729 VDD2.n24 VDD2.n23 104.615
R1730 VDD2.n24 VDD2.n13 104.615
R1731 VDD2.n31 VDD2.n13 104.615
R1732 VDD2.n32 VDD2.n31 104.615
R1733 VDD2.n32 VDD2.n9 104.615
R1734 VDD2.n39 VDD2.n9 104.615
R1735 VDD2.n40 VDD2.n39 104.615
R1736 VDD2.n40 VDD2.n5 104.615
R1737 VDD2.n47 VDD2.n5 104.615
R1738 VDD2.n48 VDD2.n47 104.615
R1739 VDD2.n48 VDD2.n1 104.615
R1740 VDD2.n55 VDD2.n1 104.615
R1741 VDD2.n114 VDD2.n56 88.2259
R1742 VDD2.t1 VDD2.n74 52.3082
R1743 VDD2.t0 VDD2.n17 52.3082
R1744 VDD2.n114 VDD2.n113 50.6096
R1745 VDD2.n76 VDD2.n75 15.6677
R1746 VDD2.n19 VDD2.n18 15.6677
R1747 VDD2.n79 VDD2.n78 12.8005
R1748 VDD2.n22 VDD2.n21 12.8005
R1749 VDD2.n82 VDD2.n73 12.0247
R1750 VDD2.n25 VDD2.n16 12.0247
R1751 VDD2.n83 VDD2.n71 11.249
R1752 VDD2.n26 VDD2.n14 11.249
R1753 VDD2.n111 VDD2.n57 10.4732
R1754 VDD2.n87 VDD2.n86 10.4732
R1755 VDD2.n30 VDD2.n29 10.4732
R1756 VDD2.n54 VDD2.n0 10.4732
R1757 VDD2.n110 VDD2.n59 9.69747
R1758 VDD2.n90 VDD2.n69 9.69747
R1759 VDD2.n33 VDD2.n12 9.69747
R1760 VDD2.n53 VDD2.n2 9.69747
R1761 VDD2.n109 VDD2.n57 9.45567
R1762 VDD2.n52 VDD2.n0 9.45567
R1763 VDD2.n110 VDD2.n109 9.3005
R1764 VDD2.n108 VDD2.n107 9.3005
R1765 VDD2.n61 VDD2.n60 9.3005
R1766 VDD2.n102 VDD2.n101 9.3005
R1767 VDD2.n100 VDD2.n99 9.3005
R1768 VDD2.n65 VDD2.n64 9.3005
R1769 VDD2.n94 VDD2.n93 9.3005
R1770 VDD2.n92 VDD2.n91 9.3005
R1771 VDD2.n69 VDD2.n68 9.3005
R1772 VDD2.n86 VDD2.n85 9.3005
R1773 VDD2.n84 VDD2.n83 9.3005
R1774 VDD2.n73 VDD2.n72 9.3005
R1775 VDD2.n78 VDD2.n77 9.3005
R1776 VDD2.n43 VDD2.n42 9.3005
R1777 VDD2.n45 VDD2.n44 9.3005
R1778 VDD2.n4 VDD2.n3 9.3005
R1779 VDD2.n51 VDD2.n50 9.3005
R1780 VDD2.n53 VDD2.n52 9.3005
R1781 VDD2.n37 VDD2.n36 9.3005
R1782 VDD2.n35 VDD2.n34 9.3005
R1783 VDD2.n12 VDD2.n11 9.3005
R1784 VDD2.n29 VDD2.n28 9.3005
R1785 VDD2.n27 VDD2.n26 9.3005
R1786 VDD2.n16 VDD2.n15 9.3005
R1787 VDD2.n21 VDD2.n20 9.3005
R1788 VDD2.n8 VDD2.n7 9.3005
R1789 VDD2.n107 VDD2.n106 8.92171
R1790 VDD2.n91 VDD2.n67 8.92171
R1791 VDD2.n34 VDD2.n10 8.92171
R1792 VDD2.n50 VDD2.n49 8.92171
R1793 VDD2.n103 VDD2.n61 8.14595
R1794 VDD2.n95 VDD2.n94 8.14595
R1795 VDD2.n38 VDD2.n37 8.14595
R1796 VDD2.n46 VDD2.n4 8.14595
R1797 VDD2.n102 VDD2.n63 7.3702
R1798 VDD2.n98 VDD2.n65 7.3702
R1799 VDD2.n41 VDD2.n8 7.3702
R1800 VDD2.n45 VDD2.n6 7.3702
R1801 VDD2.n99 VDD2.n63 6.59444
R1802 VDD2.n99 VDD2.n98 6.59444
R1803 VDD2.n42 VDD2.n41 6.59444
R1804 VDD2.n42 VDD2.n6 6.59444
R1805 VDD2.n103 VDD2.n102 5.81868
R1806 VDD2.n95 VDD2.n65 5.81868
R1807 VDD2.n38 VDD2.n8 5.81868
R1808 VDD2.n46 VDD2.n45 5.81868
R1809 VDD2.n106 VDD2.n61 5.04292
R1810 VDD2.n94 VDD2.n67 5.04292
R1811 VDD2.n37 VDD2.n10 5.04292
R1812 VDD2.n49 VDD2.n4 5.04292
R1813 VDD2.n20 VDD2.n19 4.38563
R1814 VDD2.n77 VDD2.n76 4.38563
R1815 VDD2.n107 VDD2.n59 4.26717
R1816 VDD2.n91 VDD2.n90 4.26717
R1817 VDD2.n34 VDD2.n33 4.26717
R1818 VDD2.n50 VDD2.n2 4.26717
R1819 VDD2.n111 VDD2.n110 3.49141
R1820 VDD2.n87 VDD2.n69 3.49141
R1821 VDD2.n30 VDD2.n12 3.49141
R1822 VDD2.n54 VDD2.n53 3.49141
R1823 VDD2.n113 VDD2.n57 2.71565
R1824 VDD2.n86 VDD2.n71 2.71565
R1825 VDD2.n29 VDD2.n14 2.71565
R1826 VDD2.n56 VDD2.n0 2.71565
R1827 VDD2.n83 VDD2.n82 1.93989
R1828 VDD2.n26 VDD2.n25 1.93989
R1829 VDD2.n79 VDD2.n73 1.16414
R1830 VDD2.n22 VDD2.n16 1.16414
R1831 VDD2 VDD2.n114 0.666448
R1832 VDD2.n78 VDD2.n75 0.388379
R1833 VDD2.n21 VDD2.n18 0.388379
R1834 VDD2.n109 VDD2.n108 0.155672
R1835 VDD2.n108 VDD2.n60 0.155672
R1836 VDD2.n101 VDD2.n60 0.155672
R1837 VDD2.n101 VDD2.n100 0.155672
R1838 VDD2.n100 VDD2.n64 0.155672
R1839 VDD2.n93 VDD2.n64 0.155672
R1840 VDD2.n93 VDD2.n92 0.155672
R1841 VDD2.n92 VDD2.n68 0.155672
R1842 VDD2.n85 VDD2.n68 0.155672
R1843 VDD2.n85 VDD2.n84 0.155672
R1844 VDD2.n84 VDD2.n72 0.155672
R1845 VDD2.n77 VDD2.n72 0.155672
R1846 VDD2.n20 VDD2.n15 0.155672
R1847 VDD2.n27 VDD2.n15 0.155672
R1848 VDD2.n28 VDD2.n27 0.155672
R1849 VDD2.n28 VDD2.n11 0.155672
R1850 VDD2.n35 VDD2.n11 0.155672
R1851 VDD2.n36 VDD2.n35 0.155672
R1852 VDD2.n36 VDD2.n7 0.155672
R1853 VDD2.n43 VDD2.n7 0.155672
R1854 VDD2.n44 VDD2.n43 0.155672
R1855 VDD2.n44 VDD2.n3 0.155672
R1856 VDD2.n51 VDD2.n3 0.155672
R1857 VDD2.n52 VDD2.n51 0.155672
C0 VTAIL VN 2.17867f
C1 VTAIL VDD2 4.71636f
C2 VDD1 VN 0.148071f
C3 VP VN 5.13382f
C4 VDD1 VDD2 0.661241f
C5 VP VDD2 0.328331f
C6 VTAIL VDD1 4.66625f
C7 VTAIL VP 2.19295f
C8 VP VDD1 2.63538f
C9 VDD2 VN 2.45745f
C10 VDD2 B 4.133081f
C11 VDD1 B 6.74504f
C12 VTAIL B 6.734996f
C13 VN B 10.230969f
C14 VP B 6.159474f
C15 VDD2.n0 B 0.011535f
C16 VDD2.n1 B 0.025954f
C17 VDD2.n2 B 0.011626f
C18 VDD2.n3 B 0.020434f
C19 VDD2.n4 B 0.010981f
C20 VDD2.n5 B 0.025954f
C21 VDD2.n6 B 0.011626f
C22 VDD2.n7 B 0.020434f
C23 VDD2.n8 B 0.010981f
C24 VDD2.n9 B 0.025954f
C25 VDD2.n10 B 0.011626f
C26 VDD2.n11 B 0.020434f
C27 VDD2.n12 B 0.010981f
C28 VDD2.n13 B 0.025954f
C29 VDD2.n14 B 0.011626f
C30 VDD2.n15 B 0.020434f
C31 VDD2.n16 B 0.010981f
C32 VDD2.n17 B 0.019466f
C33 VDD2.n18 B 0.015332f
C34 VDD2.t0 B 0.042484f
C35 VDD2.n19 B 0.11048f
C36 VDD2.n20 B 0.912742f
C37 VDD2.n21 B 0.010981f
C38 VDD2.n22 B 0.011626f
C39 VDD2.n23 B 0.025954f
C40 VDD2.n24 B 0.025954f
C41 VDD2.n25 B 0.011626f
C42 VDD2.n26 B 0.010981f
C43 VDD2.n27 B 0.020434f
C44 VDD2.n28 B 0.020434f
C45 VDD2.n29 B 0.010981f
C46 VDD2.n30 B 0.011626f
C47 VDD2.n31 B 0.025954f
C48 VDD2.n32 B 0.025954f
C49 VDD2.n33 B 0.011626f
C50 VDD2.n34 B 0.010981f
C51 VDD2.n35 B 0.020434f
C52 VDD2.n36 B 0.020434f
C53 VDD2.n37 B 0.010981f
C54 VDD2.n38 B 0.011626f
C55 VDD2.n39 B 0.025954f
C56 VDD2.n40 B 0.025954f
C57 VDD2.n41 B 0.011626f
C58 VDD2.n42 B 0.010981f
C59 VDD2.n43 B 0.020434f
C60 VDD2.n44 B 0.020434f
C61 VDD2.n45 B 0.010981f
C62 VDD2.n46 B 0.011626f
C63 VDD2.n47 B 0.025954f
C64 VDD2.n48 B 0.025954f
C65 VDD2.n49 B 0.011626f
C66 VDD2.n50 B 0.010981f
C67 VDD2.n51 B 0.020434f
C68 VDD2.n52 B 0.053654f
C69 VDD2.n53 B 0.010981f
C70 VDD2.n54 B 0.011626f
C71 VDD2.n55 B 0.051066f
C72 VDD2.n56 B 0.556825f
C73 VDD2.n57 B 0.011535f
C74 VDD2.n58 B 0.025954f
C75 VDD2.n59 B 0.011626f
C76 VDD2.n60 B 0.020434f
C77 VDD2.n61 B 0.010981f
C78 VDD2.n62 B 0.025954f
C79 VDD2.n63 B 0.011626f
C80 VDD2.n64 B 0.020434f
C81 VDD2.n65 B 0.010981f
C82 VDD2.n66 B 0.025954f
C83 VDD2.n67 B 0.011626f
C84 VDD2.n68 B 0.020434f
C85 VDD2.n69 B 0.010981f
C86 VDD2.n70 B 0.025954f
C87 VDD2.n71 B 0.011626f
C88 VDD2.n72 B 0.020434f
C89 VDD2.n73 B 0.010981f
C90 VDD2.n74 B 0.019466f
C91 VDD2.n75 B 0.015332f
C92 VDD2.t1 B 0.042484f
C93 VDD2.n76 B 0.11048f
C94 VDD2.n77 B 0.912742f
C95 VDD2.n78 B 0.010981f
C96 VDD2.n79 B 0.011626f
C97 VDD2.n80 B 0.025954f
C98 VDD2.n81 B 0.025954f
C99 VDD2.n82 B 0.011626f
C100 VDD2.n83 B 0.010981f
C101 VDD2.n84 B 0.020434f
C102 VDD2.n85 B 0.020434f
C103 VDD2.n86 B 0.010981f
C104 VDD2.n87 B 0.011626f
C105 VDD2.n88 B 0.025954f
C106 VDD2.n89 B 0.025954f
C107 VDD2.n90 B 0.011626f
C108 VDD2.n91 B 0.010981f
C109 VDD2.n92 B 0.020434f
C110 VDD2.n93 B 0.020434f
C111 VDD2.n94 B 0.010981f
C112 VDD2.n95 B 0.011626f
C113 VDD2.n96 B 0.025954f
C114 VDD2.n97 B 0.025954f
C115 VDD2.n98 B 0.011626f
C116 VDD2.n99 B 0.010981f
C117 VDD2.n100 B 0.020434f
C118 VDD2.n101 B 0.020434f
C119 VDD2.n102 B 0.010981f
C120 VDD2.n103 B 0.011626f
C121 VDD2.n104 B 0.025954f
C122 VDD2.n105 B 0.025954f
C123 VDD2.n106 B 0.011626f
C124 VDD2.n107 B 0.010981f
C125 VDD2.n108 B 0.020434f
C126 VDD2.n109 B 0.053654f
C127 VDD2.n110 B 0.010981f
C128 VDD2.n111 B 0.011626f
C129 VDD2.n112 B 0.051066f
C130 VDD2.n113 B 0.058186f
C131 VDD2.n114 B 2.36678f
C132 VN.t1 B 2.63781f
C133 VN.t0 B 3.13489f
C134 VDD1.n0 B 0.011574f
C135 VDD1.n1 B 0.026042f
C136 VDD1.n2 B 0.011666f
C137 VDD1.n3 B 0.020503f
C138 VDD1.n4 B 0.011018f
C139 VDD1.n5 B 0.026042f
C140 VDD1.n6 B 0.011666f
C141 VDD1.n7 B 0.020503f
C142 VDD1.n8 B 0.011018f
C143 VDD1.n9 B 0.026042f
C144 VDD1.n10 B 0.011666f
C145 VDD1.n11 B 0.020503f
C146 VDD1.n12 B 0.011018f
C147 VDD1.n13 B 0.026042f
C148 VDD1.n14 B 0.011666f
C149 VDD1.n15 B 0.020503f
C150 VDD1.n16 B 0.011018f
C151 VDD1.n17 B 0.019531f
C152 VDD1.n18 B 0.015383f
C153 VDD1.t0 B 0.042627f
C154 VDD1.n19 B 0.110852f
C155 VDD1.n20 B 0.915818f
C156 VDD1.n21 B 0.011018f
C157 VDD1.n22 B 0.011666f
C158 VDD1.n23 B 0.026042f
C159 VDD1.n24 B 0.026042f
C160 VDD1.n25 B 0.011666f
C161 VDD1.n26 B 0.011018f
C162 VDD1.n27 B 0.020503f
C163 VDD1.n28 B 0.020503f
C164 VDD1.n29 B 0.011018f
C165 VDD1.n30 B 0.011666f
C166 VDD1.n31 B 0.026042f
C167 VDD1.n32 B 0.026042f
C168 VDD1.n33 B 0.011666f
C169 VDD1.n34 B 0.011018f
C170 VDD1.n35 B 0.020503f
C171 VDD1.n36 B 0.020503f
C172 VDD1.n37 B 0.011018f
C173 VDD1.n38 B 0.011666f
C174 VDD1.n39 B 0.026042f
C175 VDD1.n40 B 0.026042f
C176 VDD1.n41 B 0.011666f
C177 VDD1.n42 B 0.011018f
C178 VDD1.n43 B 0.020503f
C179 VDD1.n44 B 0.020503f
C180 VDD1.n45 B 0.011018f
C181 VDD1.n46 B 0.011666f
C182 VDD1.n47 B 0.026042f
C183 VDD1.n48 B 0.026042f
C184 VDD1.n49 B 0.011666f
C185 VDD1.n50 B 0.011018f
C186 VDD1.n51 B 0.020503f
C187 VDD1.n52 B 0.053834f
C188 VDD1.n53 B 0.011018f
C189 VDD1.n54 B 0.011666f
C190 VDD1.n55 B 0.051238f
C191 VDD1.n56 B 0.059485f
C192 VDD1.n57 B 0.011574f
C193 VDD1.n58 B 0.026042f
C194 VDD1.n59 B 0.011666f
C195 VDD1.n60 B 0.020503f
C196 VDD1.n61 B 0.011018f
C197 VDD1.n62 B 0.026042f
C198 VDD1.n63 B 0.011666f
C199 VDD1.n64 B 0.020503f
C200 VDD1.n65 B 0.011018f
C201 VDD1.n66 B 0.026042f
C202 VDD1.n67 B 0.011666f
C203 VDD1.n68 B 0.020503f
C204 VDD1.n69 B 0.011018f
C205 VDD1.n70 B 0.026042f
C206 VDD1.n71 B 0.011666f
C207 VDD1.n72 B 0.020503f
C208 VDD1.n73 B 0.011018f
C209 VDD1.n74 B 0.019531f
C210 VDD1.n75 B 0.015383f
C211 VDD1.t1 B 0.042627f
C212 VDD1.n76 B 0.110852f
C213 VDD1.n77 B 0.915818f
C214 VDD1.n78 B 0.011018f
C215 VDD1.n79 B 0.011666f
C216 VDD1.n80 B 0.026042f
C217 VDD1.n81 B 0.026042f
C218 VDD1.n82 B 0.011666f
C219 VDD1.n83 B 0.011018f
C220 VDD1.n84 B 0.020503f
C221 VDD1.n85 B 0.020503f
C222 VDD1.n86 B 0.011018f
C223 VDD1.n87 B 0.011666f
C224 VDD1.n88 B 0.026042f
C225 VDD1.n89 B 0.026042f
C226 VDD1.n90 B 0.011666f
C227 VDD1.n91 B 0.011018f
C228 VDD1.n92 B 0.020503f
C229 VDD1.n93 B 0.020503f
C230 VDD1.n94 B 0.011018f
C231 VDD1.n95 B 0.011666f
C232 VDD1.n96 B 0.026042f
C233 VDD1.n97 B 0.026042f
C234 VDD1.n98 B 0.011666f
C235 VDD1.n99 B 0.011018f
C236 VDD1.n100 B 0.020503f
C237 VDD1.n101 B 0.020503f
C238 VDD1.n102 B 0.011018f
C239 VDD1.n103 B 0.011666f
C240 VDD1.n104 B 0.026042f
C241 VDD1.n105 B 0.026042f
C242 VDD1.n106 B 0.011666f
C243 VDD1.n107 B 0.011018f
C244 VDD1.n108 B 0.020503f
C245 VDD1.n109 B 0.053834f
C246 VDD1.n110 B 0.011018f
C247 VDD1.n111 B 0.011666f
C248 VDD1.n112 B 0.051238f
C249 VDD1.n113 B 0.596514f
C250 VTAIL.n0 B 0.011924f
C251 VTAIL.n1 B 0.02683f
C252 VTAIL.n2 B 0.012019f
C253 VTAIL.n3 B 0.021124f
C254 VTAIL.n4 B 0.011351f
C255 VTAIL.n5 B 0.02683f
C256 VTAIL.n6 B 0.012019f
C257 VTAIL.n7 B 0.021124f
C258 VTAIL.n8 B 0.011351f
C259 VTAIL.n9 B 0.02683f
C260 VTAIL.n10 B 0.012019f
C261 VTAIL.n11 B 0.021124f
C262 VTAIL.n12 B 0.011351f
C263 VTAIL.n13 B 0.02683f
C264 VTAIL.n14 B 0.012019f
C265 VTAIL.n15 B 0.021124f
C266 VTAIL.n16 B 0.011351f
C267 VTAIL.n17 B 0.020123f
C268 VTAIL.n18 B 0.015849f
C269 VTAIL.t2 B 0.043918f
C270 VTAIL.n19 B 0.11421f
C271 VTAIL.n20 B 0.943554f
C272 VTAIL.n21 B 0.011351f
C273 VTAIL.n22 B 0.012019f
C274 VTAIL.n23 B 0.02683f
C275 VTAIL.n24 B 0.02683f
C276 VTAIL.n25 B 0.012019f
C277 VTAIL.n26 B 0.011351f
C278 VTAIL.n27 B 0.021124f
C279 VTAIL.n28 B 0.021124f
C280 VTAIL.n29 B 0.011351f
C281 VTAIL.n30 B 0.012019f
C282 VTAIL.n31 B 0.02683f
C283 VTAIL.n32 B 0.02683f
C284 VTAIL.n33 B 0.012019f
C285 VTAIL.n34 B 0.011351f
C286 VTAIL.n35 B 0.021124f
C287 VTAIL.n36 B 0.021124f
C288 VTAIL.n37 B 0.011351f
C289 VTAIL.n38 B 0.012019f
C290 VTAIL.n39 B 0.02683f
C291 VTAIL.n40 B 0.02683f
C292 VTAIL.n41 B 0.012019f
C293 VTAIL.n42 B 0.011351f
C294 VTAIL.n43 B 0.021124f
C295 VTAIL.n44 B 0.021124f
C296 VTAIL.n45 B 0.011351f
C297 VTAIL.n46 B 0.012019f
C298 VTAIL.n47 B 0.02683f
C299 VTAIL.n48 B 0.02683f
C300 VTAIL.n49 B 0.012019f
C301 VTAIL.n50 B 0.011351f
C302 VTAIL.n51 B 0.021124f
C303 VTAIL.n52 B 0.055465f
C304 VTAIL.n53 B 0.011351f
C305 VTAIL.n54 B 0.012019f
C306 VTAIL.n55 B 0.05279f
C307 VTAIL.n56 B 0.045584f
C308 VTAIL.n57 B 1.33377f
C309 VTAIL.n58 B 0.011924f
C310 VTAIL.n59 B 0.02683f
C311 VTAIL.n60 B 0.012019f
C312 VTAIL.n61 B 0.021124f
C313 VTAIL.n62 B 0.011351f
C314 VTAIL.n63 B 0.02683f
C315 VTAIL.n64 B 0.012019f
C316 VTAIL.n65 B 0.021124f
C317 VTAIL.n66 B 0.011351f
C318 VTAIL.n67 B 0.02683f
C319 VTAIL.n68 B 0.012019f
C320 VTAIL.n69 B 0.021124f
C321 VTAIL.n70 B 0.011351f
C322 VTAIL.n71 B 0.02683f
C323 VTAIL.n72 B 0.012019f
C324 VTAIL.n73 B 0.021124f
C325 VTAIL.n74 B 0.011351f
C326 VTAIL.n75 B 0.020123f
C327 VTAIL.n76 B 0.015849f
C328 VTAIL.t0 B 0.043918f
C329 VTAIL.n77 B 0.11421f
C330 VTAIL.n78 B 0.943554f
C331 VTAIL.n79 B 0.011351f
C332 VTAIL.n80 B 0.012019f
C333 VTAIL.n81 B 0.02683f
C334 VTAIL.n82 B 0.02683f
C335 VTAIL.n83 B 0.012019f
C336 VTAIL.n84 B 0.011351f
C337 VTAIL.n85 B 0.021124f
C338 VTAIL.n86 B 0.021124f
C339 VTAIL.n87 B 0.011351f
C340 VTAIL.n88 B 0.012019f
C341 VTAIL.n89 B 0.02683f
C342 VTAIL.n90 B 0.02683f
C343 VTAIL.n91 B 0.012019f
C344 VTAIL.n92 B 0.011351f
C345 VTAIL.n93 B 0.021124f
C346 VTAIL.n94 B 0.021124f
C347 VTAIL.n95 B 0.011351f
C348 VTAIL.n96 B 0.012019f
C349 VTAIL.n97 B 0.02683f
C350 VTAIL.n98 B 0.02683f
C351 VTAIL.n99 B 0.012019f
C352 VTAIL.n100 B 0.011351f
C353 VTAIL.n101 B 0.021124f
C354 VTAIL.n102 B 0.021124f
C355 VTAIL.n103 B 0.011351f
C356 VTAIL.n104 B 0.012019f
C357 VTAIL.n105 B 0.02683f
C358 VTAIL.n106 B 0.02683f
C359 VTAIL.n107 B 0.012019f
C360 VTAIL.n108 B 0.011351f
C361 VTAIL.n109 B 0.021124f
C362 VTAIL.n110 B 0.055465f
C363 VTAIL.n111 B 0.011351f
C364 VTAIL.n112 B 0.012019f
C365 VTAIL.n113 B 0.05279f
C366 VTAIL.n114 B 0.045584f
C367 VTAIL.n115 B 1.37118f
C368 VTAIL.n116 B 0.011924f
C369 VTAIL.n117 B 0.02683f
C370 VTAIL.n118 B 0.012019f
C371 VTAIL.n119 B 0.021124f
C372 VTAIL.n120 B 0.011351f
C373 VTAIL.n121 B 0.02683f
C374 VTAIL.n122 B 0.012019f
C375 VTAIL.n123 B 0.021124f
C376 VTAIL.n124 B 0.011351f
C377 VTAIL.n125 B 0.02683f
C378 VTAIL.n126 B 0.012019f
C379 VTAIL.n127 B 0.021124f
C380 VTAIL.n128 B 0.011351f
C381 VTAIL.n129 B 0.02683f
C382 VTAIL.n130 B 0.012019f
C383 VTAIL.n131 B 0.021124f
C384 VTAIL.n132 B 0.011351f
C385 VTAIL.n133 B 0.020123f
C386 VTAIL.n134 B 0.015849f
C387 VTAIL.t3 B 0.043918f
C388 VTAIL.n135 B 0.11421f
C389 VTAIL.n136 B 0.943554f
C390 VTAIL.n137 B 0.011351f
C391 VTAIL.n138 B 0.012019f
C392 VTAIL.n139 B 0.02683f
C393 VTAIL.n140 B 0.02683f
C394 VTAIL.n141 B 0.012019f
C395 VTAIL.n142 B 0.011351f
C396 VTAIL.n143 B 0.021124f
C397 VTAIL.n144 B 0.021124f
C398 VTAIL.n145 B 0.011351f
C399 VTAIL.n146 B 0.012019f
C400 VTAIL.n147 B 0.02683f
C401 VTAIL.n148 B 0.02683f
C402 VTAIL.n149 B 0.012019f
C403 VTAIL.n150 B 0.011351f
C404 VTAIL.n151 B 0.021124f
C405 VTAIL.n152 B 0.021124f
C406 VTAIL.n153 B 0.011351f
C407 VTAIL.n154 B 0.012019f
C408 VTAIL.n155 B 0.02683f
C409 VTAIL.n156 B 0.02683f
C410 VTAIL.n157 B 0.012019f
C411 VTAIL.n158 B 0.011351f
C412 VTAIL.n159 B 0.021124f
C413 VTAIL.n160 B 0.021124f
C414 VTAIL.n161 B 0.011351f
C415 VTAIL.n162 B 0.012019f
C416 VTAIL.n163 B 0.02683f
C417 VTAIL.n164 B 0.02683f
C418 VTAIL.n165 B 0.012019f
C419 VTAIL.n166 B 0.011351f
C420 VTAIL.n167 B 0.021124f
C421 VTAIL.n168 B 0.055465f
C422 VTAIL.n169 B 0.011351f
C423 VTAIL.n170 B 0.012019f
C424 VTAIL.n171 B 0.05279f
C425 VTAIL.n172 B 0.045584f
C426 VTAIL.n173 B 1.2057f
C427 VTAIL.n174 B 0.011924f
C428 VTAIL.n175 B 0.02683f
C429 VTAIL.n176 B 0.012019f
C430 VTAIL.n177 B 0.021124f
C431 VTAIL.n178 B 0.011351f
C432 VTAIL.n179 B 0.02683f
C433 VTAIL.n180 B 0.012019f
C434 VTAIL.n181 B 0.021124f
C435 VTAIL.n182 B 0.011351f
C436 VTAIL.n183 B 0.02683f
C437 VTAIL.n184 B 0.012019f
C438 VTAIL.n185 B 0.021124f
C439 VTAIL.n186 B 0.011351f
C440 VTAIL.n187 B 0.02683f
C441 VTAIL.n188 B 0.012019f
C442 VTAIL.n189 B 0.021124f
C443 VTAIL.n190 B 0.011351f
C444 VTAIL.n191 B 0.020123f
C445 VTAIL.n192 B 0.015849f
C446 VTAIL.t1 B 0.043918f
C447 VTAIL.n193 B 0.11421f
C448 VTAIL.n194 B 0.943554f
C449 VTAIL.n195 B 0.011351f
C450 VTAIL.n196 B 0.012019f
C451 VTAIL.n197 B 0.02683f
C452 VTAIL.n198 B 0.02683f
C453 VTAIL.n199 B 0.012019f
C454 VTAIL.n200 B 0.011351f
C455 VTAIL.n201 B 0.021124f
C456 VTAIL.n202 B 0.021124f
C457 VTAIL.n203 B 0.011351f
C458 VTAIL.n204 B 0.012019f
C459 VTAIL.n205 B 0.02683f
C460 VTAIL.n206 B 0.02683f
C461 VTAIL.n207 B 0.012019f
C462 VTAIL.n208 B 0.011351f
C463 VTAIL.n209 B 0.021124f
C464 VTAIL.n210 B 0.021124f
C465 VTAIL.n211 B 0.011351f
C466 VTAIL.n212 B 0.012019f
C467 VTAIL.n213 B 0.02683f
C468 VTAIL.n214 B 0.02683f
C469 VTAIL.n215 B 0.012019f
C470 VTAIL.n216 B 0.011351f
C471 VTAIL.n217 B 0.021124f
C472 VTAIL.n218 B 0.021124f
C473 VTAIL.n219 B 0.011351f
C474 VTAIL.n220 B 0.012019f
C475 VTAIL.n221 B 0.02683f
C476 VTAIL.n222 B 0.02683f
C477 VTAIL.n223 B 0.012019f
C478 VTAIL.n224 B 0.011351f
C479 VTAIL.n225 B 0.021124f
C480 VTAIL.n226 B 0.055465f
C481 VTAIL.n227 B 0.011351f
C482 VTAIL.n228 B 0.012019f
C483 VTAIL.n229 B 0.05279f
C484 VTAIL.n230 B 0.045584f
C485 VTAIL.n231 B 1.1284f
C486 VP.t1 B 3.17812f
C487 VP.t0 B 2.67524f
C488 VP.n0 B 3.97149f
.ends

