**** sch_path: /home/chandru/MPW4_workdir/xschem_mpw4/LC_Cell
.subckt LC_Cell_3 Ibias outn outp ind_sub VDD GND
** Higher current mirrorring ratio 1:4, increased by 2, increasing Cap W by 4X
*.ipin Ibias
*.opin outn
*.opin outp
XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5 
XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5
XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=12
XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=12
XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC2 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC3 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC4 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
*XC5 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.3 W=2.4 nf=2
.ends

**
***Sw C1 
**XC1 outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
**XC2 net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
**XM6 net3 sw<0> net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1
***Sw C2
**XC3 outp net3 sky130_fd_pr__cap_mim_m3_1 W=32 L=5 MF=1 m=1
**XC4 net4 outn sky130_fd_pr__cap_mim_m3_1 W=32 L=5 MF=1 m=1
**XM7 net3 sw<1> net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=5
**.ends
