* NGSPICE file created from diff_pair_sample_0075.ext - technology: sky130A

.subckt diff_pair_sample_0075 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=0 ps=0 w=6.11 l=2.13
X1 VDD1.t3 VP.t0 VTAIL.t6 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=1.00815 pd=6.44 as=2.3829 ps=13 w=6.11 l=2.13
X2 B.t8 B.t6 B.t7 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=0 ps=0 w=6.11 l=2.13
X3 B.t5 B.t3 B.t4 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=0 ps=0 w=6.11 l=2.13
X4 VTAIL.t4 VP.t1 VDD1.t2 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=1.00815 ps=6.44 w=6.11 l=2.13
X5 B.t2 B.t0 B.t1 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=0 ps=0 w=6.11 l=2.13
X6 VDD2.t3 VN.t0 VTAIL.t0 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=1.00815 pd=6.44 as=2.3829 ps=13 w=6.11 l=2.13
X7 VTAIL.t1 VN.t1 VDD2.t2 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=1.00815 ps=6.44 w=6.11 l=2.13
X8 VTAIL.t7 VP.t2 VDD1.t1 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=1.00815 ps=6.44 w=6.11 l=2.13
X9 VDD1.t0 VP.t3 VTAIL.t5 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=1.00815 pd=6.44 as=2.3829 ps=13 w=6.11 l=2.13
X10 VTAIL.t3 VN.t2 VDD2.t1 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=2.3829 pd=13 as=1.00815 ps=6.44 w=6.11 l=2.13
X11 VDD2.t0 VN.t3 VTAIL.t2 w_n2446_n2190# sky130_fd_pr__pfet_01v8 ad=1.00815 pd=6.44 as=2.3829 ps=13 w=6.11 l=2.13
R0 B.n353 B.n50 585
R1 B.n355 B.n354 585
R2 B.n356 B.n49 585
R3 B.n358 B.n357 585
R4 B.n359 B.n48 585
R5 B.n361 B.n360 585
R6 B.n362 B.n47 585
R7 B.n364 B.n363 585
R8 B.n365 B.n46 585
R9 B.n367 B.n366 585
R10 B.n368 B.n45 585
R11 B.n370 B.n369 585
R12 B.n371 B.n44 585
R13 B.n373 B.n372 585
R14 B.n374 B.n43 585
R15 B.n376 B.n375 585
R16 B.n377 B.n42 585
R17 B.n379 B.n378 585
R18 B.n380 B.n41 585
R19 B.n382 B.n381 585
R20 B.n383 B.n40 585
R21 B.n385 B.n384 585
R22 B.n386 B.n39 585
R23 B.n388 B.n387 585
R24 B.n390 B.n389 585
R25 B.n391 B.n35 585
R26 B.n393 B.n392 585
R27 B.n394 B.n34 585
R28 B.n396 B.n395 585
R29 B.n397 B.n33 585
R30 B.n399 B.n398 585
R31 B.n400 B.n32 585
R32 B.n402 B.n401 585
R33 B.n403 B.n29 585
R34 B.n406 B.n405 585
R35 B.n407 B.n28 585
R36 B.n409 B.n408 585
R37 B.n410 B.n27 585
R38 B.n412 B.n411 585
R39 B.n413 B.n26 585
R40 B.n415 B.n414 585
R41 B.n416 B.n25 585
R42 B.n418 B.n417 585
R43 B.n419 B.n24 585
R44 B.n421 B.n420 585
R45 B.n422 B.n23 585
R46 B.n424 B.n423 585
R47 B.n425 B.n22 585
R48 B.n427 B.n426 585
R49 B.n428 B.n21 585
R50 B.n430 B.n429 585
R51 B.n431 B.n20 585
R52 B.n433 B.n432 585
R53 B.n434 B.n19 585
R54 B.n436 B.n435 585
R55 B.n437 B.n18 585
R56 B.n439 B.n438 585
R57 B.n440 B.n17 585
R58 B.n352 B.n351 585
R59 B.n350 B.n51 585
R60 B.n349 B.n348 585
R61 B.n347 B.n52 585
R62 B.n346 B.n345 585
R63 B.n344 B.n53 585
R64 B.n343 B.n342 585
R65 B.n341 B.n54 585
R66 B.n340 B.n339 585
R67 B.n338 B.n55 585
R68 B.n337 B.n336 585
R69 B.n335 B.n56 585
R70 B.n334 B.n333 585
R71 B.n332 B.n57 585
R72 B.n331 B.n330 585
R73 B.n329 B.n58 585
R74 B.n328 B.n327 585
R75 B.n326 B.n59 585
R76 B.n325 B.n324 585
R77 B.n323 B.n60 585
R78 B.n322 B.n321 585
R79 B.n320 B.n61 585
R80 B.n319 B.n318 585
R81 B.n317 B.n62 585
R82 B.n316 B.n315 585
R83 B.n314 B.n63 585
R84 B.n313 B.n312 585
R85 B.n311 B.n64 585
R86 B.n310 B.n309 585
R87 B.n308 B.n65 585
R88 B.n307 B.n306 585
R89 B.n305 B.n66 585
R90 B.n304 B.n303 585
R91 B.n302 B.n67 585
R92 B.n301 B.n300 585
R93 B.n299 B.n68 585
R94 B.n298 B.n297 585
R95 B.n296 B.n69 585
R96 B.n295 B.n294 585
R97 B.n293 B.n70 585
R98 B.n292 B.n291 585
R99 B.n290 B.n71 585
R100 B.n289 B.n288 585
R101 B.n287 B.n72 585
R102 B.n286 B.n285 585
R103 B.n284 B.n73 585
R104 B.n283 B.n282 585
R105 B.n281 B.n74 585
R106 B.n280 B.n279 585
R107 B.n278 B.n75 585
R108 B.n277 B.n276 585
R109 B.n275 B.n76 585
R110 B.n274 B.n273 585
R111 B.n272 B.n77 585
R112 B.n271 B.n270 585
R113 B.n269 B.n78 585
R114 B.n268 B.n267 585
R115 B.n266 B.n79 585
R116 B.n265 B.n264 585
R117 B.n263 B.n80 585
R118 B.n262 B.n261 585
R119 B.n173 B.n114 585
R120 B.n175 B.n174 585
R121 B.n176 B.n113 585
R122 B.n178 B.n177 585
R123 B.n179 B.n112 585
R124 B.n181 B.n180 585
R125 B.n182 B.n111 585
R126 B.n184 B.n183 585
R127 B.n185 B.n110 585
R128 B.n187 B.n186 585
R129 B.n188 B.n109 585
R130 B.n190 B.n189 585
R131 B.n191 B.n108 585
R132 B.n193 B.n192 585
R133 B.n194 B.n107 585
R134 B.n196 B.n195 585
R135 B.n197 B.n106 585
R136 B.n199 B.n198 585
R137 B.n200 B.n105 585
R138 B.n202 B.n201 585
R139 B.n203 B.n104 585
R140 B.n205 B.n204 585
R141 B.n206 B.n103 585
R142 B.n208 B.n207 585
R143 B.n210 B.n209 585
R144 B.n211 B.n99 585
R145 B.n213 B.n212 585
R146 B.n214 B.n98 585
R147 B.n216 B.n215 585
R148 B.n217 B.n97 585
R149 B.n219 B.n218 585
R150 B.n220 B.n96 585
R151 B.n222 B.n221 585
R152 B.n223 B.n93 585
R153 B.n226 B.n225 585
R154 B.n227 B.n92 585
R155 B.n229 B.n228 585
R156 B.n230 B.n91 585
R157 B.n232 B.n231 585
R158 B.n233 B.n90 585
R159 B.n235 B.n234 585
R160 B.n236 B.n89 585
R161 B.n238 B.n237 585
R162 B.n239 B.n88 585
R163 B.n241 B.n240 585
R164 B.n242 B.n87 585
R165 B.n244 B.n243 585
R166 B.n245 B.n86 585
R167 B.n247 B.n246 585
R168 B.n248 B.n85 585
R169 B.n250 B.n249 585
R170 B.n251 B.n84 585
R171 B.n253 B.n252 585
R172 B.n254 B.n83 585
R173 B.n256 B.n255 585
R174 B.n257 B.n82 585
R175 B.n259 B.n258 585
R176 B.n260 B.n81 585
R177 B.n172 B.n171 585
R178 B.n170 B.n115 585
R179 B.n169 B.n168 585
R180 B.n167 B.n116 585
R181 B.n166 B.n165 585
R182 B.n164 B.n117 585
R183 B.n163 B.n162 585
R184 B.n161 B.n118 585
R185 B.n160 B.n159 585
R186 B.n158 B.n119 585
R187 B.n157 B.n156 585
R188 B.n155 B.n120 585
R189 B.n154 B.n153 585
R190 B.n152 B.n121 585
R191 B.n151 B.n150 585
R192 B.n149 B.n122 585
R193 B.n148 B.n147 585
R194 B.n146 B.n123 585
R195 B.n145 B.n144 585
R196 B.n143 B.n124 585
R197 B.n142 B.n141 585
R198 B.n140 B.n125 585
R199 B.n139 B.n138 585
R200 B.n137 B.n126 585
R201 B.n136 B.n135 585
R202 B.n134 B.n127 585
R203 B.n133 B.n132 585
R204 B.n131 B.n128 585
R205 B.n130 B.n129 585
R206 B.n2 B.n0 585
R207 B.n485 B.n1 585
R208 B.n484 B.n483 585
R209 B.n482 B.n3 585
R210 B.n481 B.n480 585
R211 B.n479 B.n4 585
R212 B.n478 B.n477 585
R213 B.n476 B.n5 585
R214 B.n475 B.n474 585
R215 B.n473 B.n6 585
R216 B.n472 B.n471 585
R217 B.n470 B.n7 585
R218 B.n469 B.n468 585
R219 B.n467 B.n8 585
R220 B.n466 B.n465 585
R221 B.n464 B.n9 585
R222 B.n463 B.n462 585
R223 B.n461 B.n10 585
R224 B.n460 B.n459 585
R225 B.n458 B.n11 585
R226 B.n457 B.n456 585
R227 B.n455 B.n12 585
R228 B.n454 B.n453 585
R229 B.n452 B.n13 585
R230 B.n451 B.n450 585
R231 B.n449 B.n14 585
R232 B.n448 B.n447 585
R233 B.n446 B.n15 585
R234 B.n445 B.n444 585
R235 B.n443 B.n16 585
R236 B.n442 B.n441 585
R237 B.n487 B.n486 585
R238 B.n173 B.n172 482.89
R239 B.n442 B.n17 482.89
R240 B.n262 B.n81 482.89
R241 B.n353 B.n352 482.89
R242 B.n94 B.t8 318.036
R243 B.n36 B.t10 318.036
R244 B.n100 B.t5 318.036
R245 B.n30 B.t1 318.036
R246 B.n94 B.t6 276.339
R247 B.n100 B.t3 276.339
R248 B.n30 B.t0 276.339
R249 B.n36 B.t9 276.339
R250 B.n95 B.t7 270.327
R251 B.n37 B.t11 270.327
R252 B.n101 B.t4 270.327
R253 B.n31 B.t2 270.327
R254 B.n172 B.n115 163.367
R255 B.n168 B.n115 163.367
R256 B.n168 B.n167 163.367
R257 B.n167 B.n166 163.367
R258 B.n166 B.n117 163.367
R259 B.n162 B.n117 163.367
R260 B.n162 B.n161 163.367
R261 B.n161 B.n160 163.367
R262 B.n160 B.n119 163.367
R263 B.n156 B.n119 163.367
R264 B.n156 B.n155 163.367
R265 B.n155 B.n154 163.367
R266 B.n154 B.n121 163.367
R267 B.n150 B.n121 163.367
R268 B.n150 B.n149 163.367
R269 B.n149 B.n148 163.367
R270 B.n148 B.n123 163.367
R271 B.n144 B.n123 163.367
R272 B.n144 B.n143 163.367
R273 B.n143 B.n142 163.367
R274 B.n142 B.n125 163.367
R275 B.n138 B.n125 163.367
R276 B.n138 B.n137 163.367
R277 B.n137 B.n136 163.367
R278 B.n136 B.n127 163.367
R279 B.n132 B.n127 163.367
R280 B.n132 B.n131 163.367
R281 B.n131 B.n130 163.367
R282 B.n130 B.n2 163.367
R283 B.n486 B.n2 163.367
R284 B.n486 B.n485 163.367
R285 B.n485 B.n484 163.367
R286 B.n484 B.n3 163.367
R287 B.n480 B.n3 163.367
R288 B.n480 B.n479 163.367
R289 B.n479 B.n478 163.367
R290 B.n478 B.n5 163.367
R291 B.n474 B.n5 163.367
R292 B.n474 B.n473 163.367
R293 B.n473 B.n472 163.367
R294 B.n472 B.n7 163.367
R295 B.n468 B.n7 163.367
R296 B.n468 B.n467 163.367
R297 B.n467 B.n466 163.367
R298 B.n466 B.n9 163.367
R299 B.n462 B.n9 163.367
R300 B.n462 B.n461 163.367
R301 B.n461 B.n460 163.367
R302 B.n460 B.n11 163.367
R303 B.n456 B.n11 163.367
R304 B.n456 B.n455 163.367
R305 B.n455 B.n454 163.367
R306 B.n454 B.n13 163.367
R307 B.n450 B.n13 163.367
R308 B.n450 B.n449 163.367
R309 B.n449 B.n448 163.367
R310 B.n448 B.n15 163.367
R311 B.n444 B.n15 163.367
R312 B.n444 B.n443 163.367
R313 B.n443 B.n442 163.367
R314 B.n174 B.n173 163.367
R315 B.n174 B.n113 163.367
R316 B.n178 B.n113 163.367
R317 B.n179 B.n178 163.367
R318 B.n180 B.n179 163.367
R319 B.n180 B.n111 163.367
R320 B.n184 B.n111 163.367
R321 B.n185 B.n184 163.367
R322 B.n186 B.n185 163.367
R323 B.n186 B.n109 163.367
R324 B.n190 B.n109 163.367
R325 B.n191 B.n190 163.367
R326 B.n192 B.n191 163.367
R327 B.n192 B.n107 163.367
R328 B.n196 B.n107 163.367
R329 B.n197 B.n196 163.367
R330 B.n198 B.n197 163.367
R331 B.n198 B.n105 163.367
R332 B.n202 B.n105 163.367
R333 B.n203 B.n202 163.367
R334 B.n204 B.n203 163.367
R335 B.n204 B.n103 163.367
R336 B.n208 B.n103 163.367
R337 B.n209 B.n208 163.367
R338 B.n209 B.n99 163.367
R339 B.n213 B.n99 163.367
R340 B.n214 B.n213 163.367
R341 B.n215 B.n214 163.367
R342 B.n215 B.n97 163.367
R343 B.n219 B.n97 163.367
R344 B.n220 B.n219 163.367
R345 B.n221 B.n220 163.367
R346 B.n221 B.n93 163.367
R347 B.n226 B.n93 163.367
R348 B.n227 B.n226 163.367
R349 B.n228 B.n227 163.367
R350 B.n228 B.n91 163.367
R351 B.n232 B.n91 163.367
R352 B.n233 B.n232 163.367
R353 B.n234 B.n233 163.367
R354 B.n234 B.n89 163.367
R355 B.n238 B.n89 163.367
R356 B.n239 B.n238 163.367
R357 B.n240 B.n239 163.367
R358 B.n240 B.n87 163.367
R359 B.n244 B.n87 163.367
R360 B.n245 B.n244 163.367
R361 B.n246 B.n245 163.367
R362 B.n246 B.n85 163.367
R363 B.n250 B.n85 163.367
R364 B.n251 B.n250 163.367
R365 B.n252 B.n251 163.367
R366 B.n252 B.n83 163.367
R367 B.n256 B.n83 163.367
R368 B.n257 B.n256 163.367
R369 B.n258 B.n257 163.367
R370 B.n258 B.n81 163.367
R371 B.n263 B.n262 163.367
R372 B.n264 B.n263 163.367
R373 B.n264 B.n79 163.367
R374 B.n268 B.n79 163.367
R375 B.n269 B.n268 163.367
R376 B.n270 B.n269 163.367
R377 B.n270 B.n77 163.367
R378 B.n274 B.n77 163.367
R379 B.n275 B.n274 163.367
R380 B.n276 B.n275 163.367
R381 B.n276 B.n75 163.367
R382 B.n280 B.n75 163.367
R383 B.n281 B.n280 163.367
R384 B.n282 B.n281 163.367
R385 B.n282 B.n73 163.367
R386 B.n286 B.n73 163.367
R387 B.n287 B.n286 163.367
R388 B.n288 B.n287 163.367
R389 B.n288 B.n71 163.367
R390 B.n292 B.n71 163.367
R391 B.n293 B.n292 163.367
R392 B.n294 B.n293 163.367
R393 B.n294 B.n69 163.367
R394 B.n298 B.n69 163.367
R395 B.n299 B.n298 163.367
R396 B.n300 B.n299 163.367
R397 B.n300 B.n67 163.367
R398 B.n304 B.n67 163.367
R399 B.n305 B.n304 163.367
R400 B.n306 B.n305 163.367
R401 B.n306 B.n65 163.367
R402 B.n310 B.n65 163.367
R403 B.n311 B.n310 163.367
R404 B.n312 B.n311 163.367
R405 B.n312 B.n63 163.367
R406 B.n316 B.n63 163.367
R407 B.n317 B.n316 163.367
R408 B.n318 B.n317 163.367
R409 B.n318 B.n61 163.367
R410 B.n322 B.n61 163.367
R411 B.n323 B.n322 163.367
R412 B.n324 B.n323 163.367
R413 B.n324 B.n59 163.367
R414 B.n328 B.n59 163.367
R415 B.n329 B.n328 163.367
R416 B.n330 B.n329 163.367
R417 B.n330 B.n57 163.367
R418 B.n334 B.n57 163.367
R419 B.n335 B.n334 163.367
R420 B.n336 B.n335 163.367
R421 B.n336 B.n55 163.367
R422 B.n340 B.n55 163.367
R423 B.n341 B.n340 163.367
R424 B.n342 B.n341 163.367
R425 B.n342 B.n53 163.367
R426 B.n346 B.n53 163.367
R427 B.n347 B.n346 163.367
R428 B.n348 B.n347 163.367
R429 B.n348 B.n51 163.367
R430 B.n352 B.n51 163.367
R431 B.n438 B.n17 163.367
R432 B.n438 B.n437 163.367
R433 B.n437 B.n436 163.367
R434 B.n436 B.n19 163.367
R435 B.n432 B.n19 163.367
R436 B.n432 B.n431 163.367
R437 B.n431 B.n430 163.367
R438 B.n430 B.n21 163.367
R439 B.n426 B.n21 163.367
R440 B.n426 B.n425 163.367
R441 B.n425 B.n424 163.367
R442 B.n424 B.n23 163.367
R443 B.n420 B.n23 163.367
R444 B.n420 B.n419 163.367
R445 B.n419 B.n418 163.367
R446 B.n418 B.n25 163.367
R447 B.n414 B.n25 163.367
R448 B.n414 B.n413 163.367
R449 B.n413 B.n412 163.367
R450 B.n412 B.n27 163.367
R451 B.n408 B.n27 163.367
R452 B.n408 B.n407 163.367
R453 B.n407 B.n406 163.367
R454 B.n406 B.n29 163.367
R455 B.n401 B.n29 163.367
R456 B.n401 B.n400 163.367
R457 B.n400 B.n399 163.367
R458 B.n399 B.n33 163.367
R459 B.n395 B.n33 163.367
R460 B.n395 B.n394 163.367
R461 B.n394 B.n393 163.367
R462 B.n393 B.n35 163.367
R463 B.n389 B.n35 163.367
R464 B.n389 B.n388 163.367
R465 B.n388 B.n39 163.367
R466 B.n384 B.n39 163.367
R467 B.n384 B.n383 163.367
R468 B.n383 B.n382 163.367
R469 B.n382 B.n41 163.367
R470 B.n378 B.n41 163.367
R471 B.n378 B.n377 163.367
R472 B.n377 B.n376 163.367
R473 B.n376 B.n43 163.367
R474 B.n372 B.n43 163.367
R475 B.n372 B.n371 163.367
R476 B.n371 B.n370 163.367
R477 B.n370 B.n45 163.367
R478 B.n366 B.n45 163.367
R479 B.n366 B.n365 163.367
R480 B.n365 B.n364 163.367
R481 B.n364 B.n47 163.367
R482 B.n360 B.n47 163.367
R483 B.n360 B.n359 163.367
R484 B.n359 B.n358 163.367
R485 B.n358 B.n49 163.367
R486 B.n354 B.n49 163.367
R487 B.n354 B.n353 163.367
R488 B.n224 B.n95 59.5399
R489 B.n102 B.n101 59.5399
R490 B.n404 B.n31 59.5399
R491 B.n38 B.n37 59.5399
R492 B.n95 B.n94 47.7096
R493 B.n101 B.n100 47.7096
R494 B.n31 B.n30 47.7096
R495 B.n37 B.n36 47.7096
R496 B.n441 B.n440 31.3761
R497 B.n351 B.n50 31.3761
R498 B.n261 B.n260 31.3761
R499 B.n171 B.n114 31.3761
R500 B B.n487 18.0485
R501 B.n440 B.n439 10.6151
R502 B.n439 B.n18 10.6151
R503 B.n435 B.n18 10.6151
R504 B.n435 B.n434 10.6151
R505 B.n434 B.n433 10.6151
R506 B.n433 B.n20 10.6151
R507 B.n429 B.n20 10.6151
R508 B.n429 B.n428 10.6151
R509 B.n428 B.n427 10.6151
R510 B.n427 B.n22 10.6151
R511 B.n423 B.n22 10.6151
R512 B.n423 B.n422 10.6151
R513 B.n422 B.n421 10.6151
R514 B.n421 B.n24 10.6151
R515 B.n417 B.n24 10.6151
R516 B.n417 B.n416 10.6151
R517 B.n416 B.n415 10.6151
R518 B.n415 B.n26 10.6151
R519 B.n411 B.n26 10.6151
R520 B.n411 B.n410 10.6151
R521 B.n410 B.n409 10.6151
R522 B.n409 B.n28 10.6151
R523 B.n405 B.n28 10.6151
R524 B.n403 B.n402 10.6151
R525 B.n402 B.n32 10.6151
R526 B.n398 B.n32 10.6151
R527 B.n398 B.n397 10.6151
R528 B.n397 B.n396 10.6151
R529 B.n396 B.n34 10.6151
R530 B.n392 B.n34 10.6151
R531 B.n392 B.n391 10.6151
R532 B.n391 B.n390 10.6151
R533 B.n387 B.n386 10.6151
R534 B.n386 B.n385 10.6151
R535 B.n385 B.n40 10.6151
R536 B.n381 B.n40 10.6151
R537 B.n381 B.n380 10.6151
R538 B.n380 B.n379 10.6151
R539 B.n379 B.n42 10.6151
R540 B.n375 B.n42 10.6151
R541 B.n375 B.n374 10.6151
R542 B.n374 B.n373 10.6151
R543 B.n373 B.n44 10.6151
R544 B.n369 B.n44 10.6151
R545 B.n369 B.n368 10.6151
R546 B.n368 B.n367 10.6151
R547 B.n367 B.n46 10.6151
R548 B.n363 B.n46 10.6151
R549 B.n363 B.n362 10.6151
R550 B.n362 B.n361 10.6151
R551 B.n361 B.n48 10.6151
R552 B.n357 B.n48 10.6151
R553 B.n357 B.n356 10.6151
R554 B.n356 B.n355 10.6151
R555 B.n355 B.n50 10.6151
R556 B.n261 B.n80 10.6151
R557 B.n265 B.n80 10.6151
R558 B.n266 B.n265 10.6151
R559 B.n267 B.n266 10.6151
R560 B.n267 B.n78 10.6151
R561 B.n271 B.n78 10.6151
R562 B.n272 B.n271 10.6151
R563 B.n273 B.n272 10.6151
R564 B.n273 B.n76 10.6151
R565 B.n277 B.n76 10.6151
R566 B.n278 B.n277 10.6151
R567 B.n279 B.n278 10.6151
R568 B.n279 B.n74 10.6151
R569 B.n283 B.n74 10.6151
R570 B.n284 B.n283 10.6151
R571 B.n285 B.n284 10.6151
R572 B.n285 B.n72 10.6151
R573 B.n289 B.n72 10.6151
R574 B.n290 B.n289 10.6151
R575 B.n291 B.n290 10.6151
R576 B.n291 B.n70 10.6151
R577 B.n295 B.n70 10.6151
R578 B.n296 B.n295 10.6151
R579 B.n297 B.n296 10.6151
R580 B.n297 B.n68 10.6151
R581 B.n301 B.n68 10.6151
R582 B.n302 B.n301 10.6151
R583 B.n303 B.n302 10.6151
R584 B.n303 B.n66 10.6151
R585 B.n307 B.n66 10.6151
R586 B.n308 B.n307 10.6151
R587 B.n309 B.n308 10.6151
R588 B.n309 B.n64 10.6151
R589 B.n313 B.n64 10.6151
R590 B.n314 B.n313 10.6151
R591 B.n315 B.n314 10.6151
R592 B.n315 B.n62 10.6151
R593 B.n319 B.n62 10.6151
R594 B.n320 B.n319 10.6151
R595 B.n321 B.n320 10.6151
R596 B.n321 B.n60 10.6151
R597 B.n325 B.n60 10.6151
R598 B.n326 B.n325 10.6151
R599 B.n327 B.n326 10.6151
R600 B.n327 B.n58 10.6151
R601 B.n331 B.n58 10.6151
R602 B.n332 B.n331 10.6151
R603 B.n333 B.n332 10.6151
R604 B.n333 B.n56 10.6151
R605 B.n337 B.n56 10.6151
R606 B.n338 B.n337 10.6151
R607 B.n339 B.n338 10.6151
R608 B.n339 B.n54 10.6151
R609 B.n343 B.n54 10.6151
R610 B.n344 B.n343 10.6151
R611 B.n345 B.n344 10.6151
R612 B.n345 B.n52 10.6151
R613 B.n349 B.n52 10.6151
R614 B.n350 B.n349 10.6151
R615 B.n351 B.n350 10.6151
R616 B.n175 B.n114 10.6151
R617 B.n176 B.n175 10.6151
R618 B.n177 B.n176 10.6151
R619 B.n177 B.n112 10.6151
R620 B.n181 B.n112 10.6151
R621 B.n182 B.n181 10.6151
R622 B.n183 B.n182 10.6151
R623 B.n183 B.n110 10.6151
R624 B.n187 B.n110 10.6151
R625 B.n188 B.n187 10.6151
R626 B.n189 B.n188 10.6151
R627 B.n189 B.n108 10.6151
R628 B.n193 B.n108 10.6151
R629 B.n194 B.n193 10.6151
R630 B.n195 B.n194 10.6151
R631 B.n195 B.n106 10.6151
R632 B.n199 B.n106 10.6151
R633 B.n200 B.n199 10.6151
R634 B.n201 B.n200 10.6151
R635 B.n201 B.n104 10.6151
R636 B.n205 B.n104 10.6151
R637 B.n206 B.n205 10.6151
R638 B.n207 B.n206 10.6151
R639 B.n211 B.n210 10.6151
R640 B.n212 B.n211 10.6151
R641 B.n212 B.n98 10.6151
R642 B.n216 B.n98 10.6151
R643 B.n217 B.n216 10.6151
R644 B.n218 B.n217 10.6151
R645 B.n218 B.n96 10.6151
R646 B.n222 B.n96 10.6151
R647 B.n223 B.n222 10.6151
R648 B.n225 B.n92 10.6151
R649 B.n229 B.n92 10.6151
R650 B.n230 B.n229 10.6151
R651 B.n231 B.n230 10.6151
R652 B.n231 B.n90 10.6151
R653 B.n235 B.n90 10.6151
R654 B.n236 B.n235 10.6151
R655 B.n237 B.n236 10.6151
R656 B.n237 B.n88 10.6151
R657 B.n241 B.n88 10.6151
R658 B.n242 B.n241 10.6151
R659 B.n243 B.n242 10.6151
R660 B.n243 B.n86 10.6151
R661 B.n247 B.n86 10.6151
R662 B.n248 B.n247 10.6151
R663 B.n249 B.n248 10.6151
R664 B.n249 B.n84 10.6151
R665 B.n253 B.n84 10.6151
R666 B.n254 B.n253 10.6151
R667 B.n255 B.n254 10.6151
R668 B.n255 B.n82 10.6151
R669 B.n259 B.n82 10.6151
R670 B.n260 B.n259 10.6151
R671 B.n171 B.n170 10.6151
R672 B.n170 B.n169 10.6151
R673 B.n169 B.n116 10.6151
R674 B.n165 B.n116 10.6151
R675 B.n165 B.n164 10.6151
R676 B.n164 B.n163 10.6151
R677 B.n163 B.n118 10.6151
R678 B.n159 B.n118 10.6151
R679 B.n159 B.n158 10.6151
R680 B.n158 B.n157 10.6151
R681 B.n157 B.n120 10.6151
R682 B.n153 B.n120 10.6151
R683 B.n153 B.n152 10.6151
R684 B.n152 B.n151 10.6151
R685 B.n151 B.n122 10.6151
R686 B.n147 B.n122 10.6151
R687 B.n147 B.n146 10.6151
R688 B.n146 B.n145 10.6151
R689 B.n145 B.n124 10.6151
R690 B.n141 B.n124 10.6151
R691 B.n141 B.n140 10.6151
R692 B.n140 B.n139 10.6151
R693 B.n139 B.n126 10.6151
R694 B.n135 B.n126 10.6151
R695 B.n135 B.n134 10.6151
R696 B.n134 B.n133 10.6151
R697 B.n133 B.n128 10.6151
R698 B.n129 B.n128 10.6151
R699 B.n129 B.n0 10.6151
R700 B.n483 B.n1 10.6151
R701 B.n483 B.n482 10.6151
R702 B.n482 B.n481 10.6151
R703 B.n481 B.n4 10.6151
R704 B.n477 B.n4 10.6151
R705 B.n477 B.n476 10.6151
R706 B.n476 B.n475 10.6151
R707 B.n475 B.n6 10.6151
R708 B.n471 B.n6 10.6151
R709 B.n471 B.n470 10.6151
R710 B.n470 B.n469 10.6151
R711 B.n469 B.n8 10.6151
R712 B.n465 B.n8 10.6151
R713 B.n465 B.n464 10.6151
R714 B.n464 B.n463 10.6151
R715 B.n463 B.n10 10.6151
R716 B.n459 B.n10 10.6151
R717 B.n459 B.n458 10.6151
R718 B.n458 B.n457 10.6151
R719 B.n457 B.n12 10.6151
R720 B.n453 B.n12 10.6151
R721 B.n453 B.n452 10.6151
R722 B.n452 B.n451 10.6151
R723 B.n451 B.n14 10.6151
R724 B.n447 B.n14 10.6151
R725 B.n447 B.n446 10.6151
R726 B.n446 B.n445 10.6151
R727 B.n445 B.n16 10.6151
R728 B.n441 B.n16 10.6151
R729 B.n405 B.n404 9.36635
R730 B.n387 B.n38 9.36635
R731 B.n207 B.n102 9.36635
R732 B.n225 B.n224 9.36635
R733 B.n487 B.n0 2.81026
R734 B.n487 B.n1 2.81026
R735 B.n404 B.n403 1.24928
R736 B.n390 B.n38 1.24928
R737 B.n210 B.n102 1.24928
R738 B.n224 B.n223 1.24928
R739 VP.n10 VP.n0 161.3
R740 VP.n9 VP.n8 161.3
R741 VP.n7 VP.n1 161.3
R742 VP.n6 VP.n5 161.3
R743 VP.n2 VP.t2 105.379
R744 VP.n2 VP.t3 104.826
R745 VP.n4 VP.n3 87.2681
R746 VP.n12 VP.n11 87.2681
R747 VP.n4 VP.t1 69.1324
R748 VP.n11 VP.t0 69.1324
R749 VP.n9 VP.n1 56.5193
R750 VP.n3 VP.n2 47.2629
R751 VP.n5 VP.n1 24.4675
R752 VP.n10 VP.n9 24.4675
R753 VP.n5 VP.n4 23.4888
R754 VP.n11 VP.n10 23.4888
R755 VP.n6 VP.n3 0.278367
R756 VP.n12 VP.n0 0.278367
R757 VP.n7 VP.n6 0.189894
R758 VP.n8 VP.n7 0.189894
R759 VP.n8 VP.n0 0.189894
R760 VP VP.n12 0.153454
R761 VTAIL.n250 VTAIL.n224 756.745
R762 VTAIL.n26 VTAIL.n0 756.745
R763 VTAIL.n58 VTAIL.n32 756.745
R764 VTAIL.n90 VTAIL.n64 756.745
R765 VTAIL.n218 VTAIL.n192 756.745
R766 VTAIL.n186 VTAIL.n160 756.745
R767 VTAIL.n154 VTAIL.n128 756.745
R768 VTAIL.n122 VTAIL.n96 756.745
R769 VTAIL.n235 VTAIL.n234 585
R770 VTAIL.n232 VTAIL.n231 585
R771 VTAIL.n241 VTAIL.n240 585
R772 VTAIL.n243 VTAIL.n242 585
R773 VTAIL.n228 VTAIL.n227 585
R774 VTAIL.n249 VTAIL.n248 585
R775 VTAIL.n251 VTAIL.n250 585
R776 VTAIL.n11 VTAIL.n10 585
R777 VTAIL.n8 VTAIL.n7 585
R778 VTAIL.n17 VTAIL.n16 585
R779 VTAIL.n19 VTAIL.n18 585
R780 VTAIL.n4 VTAIL.n3 585
R781 VTAIL.n25 VTAIL.n24 585
R782 VTAIL.n27 VTAIL.n26 585
R783 VTAIL.n43 VTAIL.n42 585
R784 VTAIL.n40 VTAIL.n39 585
R785 VTAIL.n49 VTAIL.n48 585
R786 VTAIL.n51 VTAIL.n50 585
R787 VTAIL.n36 VTAIL.n35 585
R788 VTAIL.n57 VTAIL.n56 585
R789 VTAIL.n59 VTAIL.n58 585
R790 VTAIL.n75 VTAIL.n74 585
R791 VTAIL.n72 VTAIL.n71 585
R792 VTAIL.n81 VTAIL.n80 585
R793 VTAIL.n83 VTAIL.n82 585
R794 VTAIL.n68 VTAIL.n67 585
R795 VTAIL.n89 VTAIL.n88 585
R796 VTAIL.n91 VTAIL.n90 585
R797 VTAIL.n219 VTAIL.n218 585
R798 VTAIL.n217 VTAIL.n216 585
R799 VTAIL.n196 VTAIL.n195 585
R800 VTAIL.n211 VTAIL.n210 585
R801 VTAIL.n209 VTAIL.n208 585
R802 VTAIL.n200 VTAIL.n199 585
R803 VTAIL.n203 VTAIL.n202 585
R804 VTAIL.n187 VTAIL.n186 585
R805 VTAIL.n185 VTAIL.n184 585
R806 VTAIL.n164 VTAIL.n163 585
R807 VTAIL.n179 VTAIL.n178 585
R808 VTAIL.n177 VTAIL.n176 585
R809 VTAIL.n168 VTAIL.n167 585
R810 VTAIL.n171 VTAIL.n170 585
R811 VTAIL.n155 VTAIL.n154 585
R812 VTAIL.n153 VTAIL.n152 585
R813 VTAIL.n132 VTAIL.n131 585
R814 VTAIL.n147 VTAIL.n146 585
R815 VTAIL.n145 VTAIL.n144 585
R816 VTAIL.n136 VTAIL.n135 585
R817 VTAIL.n139 VTAIL.n138 585
R818 VTAIL.n123 VTAIL.n122 585
R819 VTAIL.n121 VTAIL.n120 585
R820 VTAIL.n100 VTAIL.n99 585
R821 VTAIL.n115 VTAIL.n114 585
R822 VTAIL.n113 VTAIL.n112 585
R823 VTAIL.n104 VTAIL.n103 585
R824 VTAIL.n107 VTAIL.n106 585
R825 VTAIL.t2 VTAIL.n233 327.601
R826 VTAIL.t3 VTAIL.n9 327.601
R827 VTAIL.t6 VTAIL.n41 327.601
R828 VTAIL.t4 VTAIL.n73 327.601
R829 VTAIL.t5 VTAIL.n201 327.601
R830 VTAIL.t7 VTAIL.n169 327.601
R831 VTAIL.t0 VTAIL.n137 327.601
R832 VTAIL.t1 VTAIL.n105 327.601
R833 VTAIL.n234 VTAIL.n231 171.744
R834 VTAIL.n241 VTAIL.n231 171.744
R835 VTAIL.n242 VTAIL.n241 171.744
R836 VTAIL.n242 VTAIL.n227 171.744
R837 VTAIL.n249 VTAIL.n227 171.744
R838 VTAIL.n250 VTAIL.n249 171.744
R839 VTAIL.n10 VTAIL.n7 171.744
R840 VTAIL.n17 VTAIL.n7 171.744
R841 VTAIL.n18 VTAIL.n17 171.744
R842 VTAIL.n18 VTAIL.n3 171.744
R843 VTAIL.n25 VTAIL.n3 171.744
R844 VTAIL.n26 VTAIL.n25 171.744
R845 VTAIL.n42 VTAIL.n39 171.744
R846 VTAIL.n49 VTAIL.n39 171.744
R847 VTAIL.n50 VTAIL.n49 171.744
R848 VTAIL.n50 VTAIL.n35 171.744
R849 VTAIL.n57 VTAIL.n35 171.744
R850 VTAIL.n58 VTAIL.n57 171.744
R851 VTAIL.n74 VTAIL.n71 171.744
R852 VTAIL.n81 VTAIL.n71 171.744
R853 VTAIL.n82 VTAIL.n81 171.744
R854 VTAIL.n82 VTAIL.n67 171.744
R855 VTAIL.n89 VTAIL.n67 171.744
R856 VTAIL.n90 VTAIL.n89 171.744
R857 VTAIL.n218 VTAIL.n217 171.744
R858 VTAIL.n217 VTAIL.n195 171.744
R859 VTAIL.n210 VTAIL.n195 171.744
R860 VTAIL.n210 VTAIL.n209 171.744
R861 VTAIL.n209 VTAIL.n199 171.744
R862 VTAIL.n202 VTAIL.n199 171.744
R863 VTAIL.n186 VTAIL.n185 171.744
R864 VTAIL.n185 VTAIL.n163 171.744
R865 VTAIL.n178 VTAIL.n163 171.744
R866 VTAIL.n178 VTAIL.n177 171.744
R867 VTAIL.n177 VTAIL.n167 171.744
R868 VTAIL.n170 VTAIL.n167 171.744
R869 VTAIL.n154 VTAIL.n153 171.744
R870 VTAIL.n153 VTAIL.n131 171.744
R871 VTAIL.n146 VTAIL.n131 171.744
R872 VTAIL.n146 VTAIL.n145 171.744
R873 VTAIL.n145 VTAIL.n135 171.744
R874 VTAIL.n138 VTAIL.n135 171.744
R875 VTAIL.n122 VTAIL.n121 171.744
R876 VTAIL.n121 VTAIL.n99 171.744
R877 VTAIL.n114 VTAIL.n99 171.744
R878 VTAIL.n114 VTAIL.n113 171.744
R879 VTAIL.n113 VTAIL.n103 171.744
R880 VTAIL.n106 VTAIL.n103 171.744
R881 VTAIL.n234 VTAIL.t2 85.8723
R882 VTAIL.n10 VTAIL.t3 85.8723
R883 VTAIL.n42 VTAIL.t6 85.8723
R884 VTAIL.n74 VTAIL.t4 85.8723
R885 VTAIL.n202 VTAIL.t5 85.8723
R886 VTAIL.n170 VTAIL.t7 85.8723
R887 VTAIL.n138 VTAIL.t0 85.8723
R888 VTAIL.n106 VTAIL.t1 85.8723
R889 VTAIL.n255 VTAIL.n254 34.3187
R890 VTAIL.n31 VTAIL.n30 34.3187
R891 VTAIL.n63 VTAIL.n62 34.3187
R892 VTAIL.n95 VTAIL.n94 34.3187
R893 VTAIL.n223 VTAIL.n222 34.3187
R894 VTAIL.n191 VTAIL.n190 34.3187
R895 VTAIL.n159 VTAIL.n158 34.3187
R896 VTAIL.n127 VTAIL.n126 34.3187
R897 VTAIL.n255 VTAIL.n223 19.7548
R898 VTAIL.n127 VTAIL.n95 19.7548
R899 VTAIL.n235 VTAIL.n233 16.3865
R900 VTAIL.n11 VTAIL.n9 16.3865
R901 VTAIL.n43 VTAIL.n41 16.3865
R902 VTAIL.n75 VTAIL.n73 16.3865
R903 VTAIL.n203 VTAIL.n201 16.3865
R904 VTAIL.n171 VTAIL.n169 16.3865
R905 VTAIL.n139 VTAIL.n137 16.3865
R906 VTAIL.n107 VTAIL.n105 16.3865
R907 VTAIL.n236 VTAIL.n232 12.8005
R908 VTAIL.n12 VTAIL.n8 12.8005
R909 VTAIL.n44 VTAIL.n40 12.8005
R910 VTAIL.n76 VTAIL.n72 12.8005
R911 VTAIL.n204 VTAIL.n200 12.8005
R912 VTAIL.n172 VTAIL.n168 12.8005
R913 VTAIL.n140 VTAIL.n136 12.8005
R914 VTAIL.n108 VTAIL.n104 12.8005
R915 VTAIL.n240 VTAIL.n239 12.0247
R916 VTAIL.n16 VTAIL.n15 12.0247
R917 VTAIL.n48 VTAIL.n47 12.0247
R918 VTAIL.n80 VTAIL.n79 12.0247
R919 VTAIL.n208 VTAIL.n207 12.0247
R920 VTAIL.n176 VTAIL.n175 12.0247
R921 VTAIL.n144 VTAIL.n143 12.0247
R922 VTAIL.n112 VTAIL.n111 12.0247
R923 VTAIL.n243 VTAIL.n230 11.249
R924 VTAIL.n19 VTAIL.n6 11.249
R925 VTAIL.n51 VTAIL.n38 11.249
R926 VTAIL.n83 VTAIL.n70 11.249
R927 VTAIL.n211 VTAIL.n198 11.249
R928 VTAIL.n179 VTAIL.n166 11.249
R929 VTAIL.n147 VTAIL.n134 11.249
R930 VTAIL.n115 VTAIL.n102 11.249
R931 VTAIL.n244 VTAIL.n228 10.4732
R932 VTAIL.n20 VTAIL.n4 10.4732
R933 VTAIL.n52 VTAIL.n36 10.4732
R934 VTAIL.n84 VTAIL.n68 10.4732
R935 VTAIL.n212 VTAIL.n196 10.4732
R936 VTAIL.n180 VTAIL.n164 10.4732
R937 VTAIL.n148 VTAIL.n132 10.4732
R938 VTAIL.n116 VTAIL.n100 10.4732
R939 VTAIL.n248 VTAIL.n247 9.69747
R940 VTAIL.n24 VTAIL.n23 9.69747
R941 VTAIL.n56 VTAIL.n55 9.69747
R942 VTAIL.n88 VTAIL.n87 9.69747
R943 VTAIL.n216 VTAIL.n215 9.69747
R944 VTAIL.n184 VTAIL.n183 9.69747
R945 VTAIL.n152 VTAIL.n151 9.69747
R946 VTAIL.n120 VTAIL.n119 9.69747
R947 VTAIL.n254 VTAIL.n253 9.45567
R948 VTAIL.n30 VTAIL.n29 9.45567
R949 VTAIL.n62 VTAIL.n61 9.45567
R950 VTAIL.n94 VTAIL.n93 9.45567
R951 VTAIL.n222 VTAIL.n221 9.45567
R952 VTAIL.n190 VTAIL.n189 9.45567
R953 VTAIL.n158 VTAIL.n157 9.45567
R954 VTAIL.n126 VTAIL.n125 9.45567
R955 VTAIL.n253 VTAIL.n252 9.3005
R956 VTAIL.n226 VTAIL.n225 9.3005
R957 VTAIL.n247 VTAIL.n246 9.3005
R958 VTAIL.n245 VTAIL.n244 9.3005
R959 VTAIL.n230 VTAIL.n229 9.3005
R960 VTAIL.n239 VTAIL.n238 9.3005
R961 VTAIL.n237 VTAIL.n236 9.3005
R962 VTAIL.n29 VTAIL.n28 9.3005
R963 VTAIL.n2 VTAIL.n1 9.3005
R964 VTAIL.n23 VTAIL.n22 9.3005
R965 VTAIL.n21 VTAIL.n20 9.3005
R966 VTAIL.n6 VTAIL.n5 9.3005
R967 VTAIL.n15 VTAIL.n14 9.3005
R968 VTAIL.n13 VTAIL.n12 9.3005
R969 VTAIL.n61 VTAIL.n60 9.3005
R970 VTAIL.n34 VTAIL.n33 9.3005
R971 VTAIL.n55 VTAIL.n54 9.3005
R972 VTAIL.n53 VTAIL.n52 9.3005
R973 VTAIL.n38 VTAIL.n37 9.3005
R974 VTAIL.n47 VTAIL.n46 9.3005
R975 VTAIL.n45 VTAIL.n44 9.3005
R976 VTAIL.n93 VTAIL.n92 9.3005
R977 VTAIL.n66 VTAIL.n65 9.3005
R978 VTAIL.n87 VTAIL.n86 9.3005
R979 VTAIL.n85 VTAIL.n84 9.3005
R980 VTAIL.n70 VTAIL.n69 9.3005
R981 VTAIL.n79 VTAIL.n78 9.3005
R982 VTAIL.n77 VTAIL.n76 9.3005
R983 VTAIL.n221 VTAIL.n220 9.3005
R984 VTAIL.n194 VTAIL.n193 9.3005
R985 VTAIL.n215 VTAIL.n214 9.3005
R986 VTAIL.n213 VTAIL.n212 9.3005
R987 VTAIL.n198 VTAIL.n197 9.3005
R988 VTAIL.n207 VTAIL.n206 9.3005
R989 VTAIL.n205 VTAIL.n204 9.3005
R990 VTAIL.n189 VTAIL.n188 9.3005
R991 VTAIL.n162 VTAIL.n161 9.3005
R992 VTAIL.n183 VTAIL.n182 9.3005
R993 VTAIL.n181 VTAIL.n180 9.3005
R994 VTAIL.n166 VTAIL.n165 9.3005
R995 VTAIL.n175 VTAIL.n174 9.3005
R996 VTAIL.n173 VTAIL.n172 9.3005
R997 VTAIL.n157 VTAIL.n156 9.3005
R998 VTAIL.n130 VTAIL.n129 9.3005
R999 VTAIL.n151 VTAIL.n150 9.3005
R1000 VTAIL.n149 VTAIL.n148 9.3005
R1001 VTAIL.n134 VTAIL.n133 9.3005
R1002 VTAIL.n143 VTAIL.n142 9.3005
R1003 VTAIL.n141 VTAIL.n140 9.3005
R1004 VTAIL.n125 VTAIL.n124 9.3005
R1005 VTAIL.n98 VTAIL.n97 9.3005
R1006 VTAIL.n119 VTAIL.n118 9.3005
R1007 VTAIL.n117 VTAIL.n116 9.3005
R1008 VTAIL.n102 VTAIL.n101 9.3005
R1009 VTAIL.n111 VTAIL.n110 9.3005
R1010 VTAIL.n109 VTAIL.n108 9.3005
R1011 VTAIL.n251 VTAIL.n226 8.92171
R1012 VTAIL.n27 VTAIL.n2 8.92171
R1013 VTAIL.n59 VTAIL.n34 8.92171
R1014 VTAIL.n91 VTAIL.n66 8.92171
R1015 VTAIL.n219 VTAIL.n194 8.92171
R1016 VTAIL.n187 VTAIL.n162 8.92171
R1017 VTAIL.n155 VTAIL.n130 8.92171
R1018 VTAIL.n123 VTAIL.n98 8.92171
R1019 VTAIL.n252 VTAIL.n224 8.14595
R1020 VTAIL.n28 VTAIL.n0 8.14595
R1021 VTAIL.n60 VTAIL.n32 8.14595
R1022 VTAIL.n92 VTAIL.n64 8.14595
R1023 VTAIL.n220 VTAIL.n192 8.14595
R1024 VTAIL.n188 VTAIL.n160 8.14595
R1025 VTAIL.n156 VTAIL.n128 8.14595
R1026 VTAIL.n124 VTAIL.n96 8.14595
R1027 VTAIL.n254 VTAIL.n224 5.81868
R1028 VTAIL.n30 VTAIL.n0 5.81868
R1029 VTAIL.n62 VTAIL.n32 5.81868
R1030 VTAIL.n94 VTAIL.n64 5.81868
R1031 VTAIL.n222 VTAIL.n192 5.81868
R1032 VTAIL.n190 VTAIL.n160 5.81868
R1033 VTAIL.n158 VTAIL.n128 5.81868
R1034 VTAIL.n126 VTAIL.n96 5.81868
R1035 VTAIL.n252 VTAIL.n251 5.04292
R1036 VTAIL.n28 VTAIL.n27 5.04292
R1037 VTAIL.n60 VTAIL.n59 5.04292
R1038 VTAIL.n92 VTAIL.n91 5.04292
R1039 VTAIL.n220 VTAIL.n219 5.04292
R1040 VTAIL.n188 VTAIL.n187 5.04292
R1041 VTAIL.n156 VTAIL.n155 5.04292
R1042 VTAIL.n124 VTAIL.n123 5.04292
R1043 VTAIL.n248 VTAIL.n226 4.26717
R1044 VTAIL.n24 VTAIL.n2 4.26717
R1045 VTAIL.n56 VTAIL.n34 4.26717
R1046 VTAIL.n88 VTAIL.n66 4.26717
R1047 VTAIL.n216 VTAIL.n194 4.26717
R1048 VTAIL.n184 VTAIL.n162 4.26717
R1049 VTAIL.n152 VTAIL.n130 4.26717
R1050 VTAIL.n120 VTAIL.n98 4.26717
R1051 VTAIL.n205 VTAIL.n201 3.71286
R1052 VTAIL.n173 VTAIL.n169 3.71286
R1053 VTAIL.n141 VTAIL.n137 3.71286
R1054 VTAIL.n109 VTAIL.n105 3.71286
R1055 VTAIL.n237 VTAIL.n233 3.71286
R1056 VTAIL.n13 VTAIL.n9 3.71286
R1057 VTAIL.n45 VTAIL.n41 3.71286
R1058 VTAIL.n77 VTAIL.n73 3.71286
R1059 VTAIL.n247 VTAIL.n228 3.49141
R1060 VTAIL.n23 VTAIL.n4 3.49141
R1061 VTAIL.n55 VTAIL.n36 3.49141
R1062 VTAIL.n87 VTAIL.n68 3.49141
R1063 VTAIL.n215 VTAIL.n196 3.49141
R1064 VTAIL.n183 VTAIL.n164 3.49141
R1065 VTAIL.n151 VTAIL.n132 3.49141
R1066 VTAIL.n119 VTAIL.n100 3.49141
R1067 VTAIL.n244 VTAIL.n243 2.71565
R1068 VTAIL.n20 VTAIL.n19 2.71565
R1069 VTAIL.n52 VTAIL.n51 2.71565
R1070 VTAIL.n84 VTAIL.n83 2.71565
R1071 VTAIL.n212 VTAIL.n211 2.71565
R1072 VTAIL.n180 VTAIL.n179 2.71565
R1073 VTAIL.n148 VTAIL.n147 2.71565
R1074 VTAIL.n116 VTAIL.n115 2.71565
R1075 VTAIL.n159 VTAIL.n127 2.12119
R1076 VTAIL.n223 VTAIL.n191 2.12119
R1077 VTAIL.n95 VTAIL.n63 2.12119
R1078 VTAIL.n240 VTAIL.n230 1.93989
R1079 VTAIL.n16 VTAIL.n6 1.93989
R1080 VTAIL.n48 VTAIL.n38 1.93989
R1081 VTAIL.n80 VTAIL.n70 1.93989
R1082 VTAIL.n208 VTAIL.n198 1.93989
R1083 VTAIL.n176 VTAIL.n166 1.93989
R1084 VTAIL.n144 VTAIL.n134 1.93989
R1085 VTAIL.n112 VTAIL.n102 1.93989
R1086 VTAIL.n239 VTAIL.n232 1.16414
R1087 VTAIL.n15 VTAIL.n8 1.16414
R1088 VTAIL.n47 VTAIL.n40 1.16414
R1089 VTAIL.n79 VTAIL.n72 1.16414
R1090 VTAIL.n207 VTAIL.n200 1.16414
R1091 VTAIL.n175 VTAIL.n168 1.16414
R1092 VTAIL.n143 VTAIL.n136 1.16414
R1093 VTAIL.n111 VTAIL.n104 1.16414
R1094 VTAIL VTAIL.n31 1.11903
R1095 VTAIL VTAIL.n255 1.00266
R1096 VTAIL.n191 VTAIL.n159 0.470328
R1097 VTAIL.n63 VTAIL.n31 0.470328
R1098 VTAIL.n236 VTAIL.n235 0.388379
R1099 VTAIL.n12 VTAIL.n11 0.388379
R1100 VTAIL.n44 VTAIL.n43 0.388379
R1101 VTAIL.n76 VTAIL.n75 0.388379
R1102 VTAIL.n204 VTAIL.n203 0.388379
R1103 VTAIL.n172 VTAIL.n171 0.388379
R1104 VTAIL.n140 VTAIL.n139 0.388379
R1105 VTAIL.n108 VTAIL.n107 0.388379
R1106 VTAIL.n238 VTAIL.n237 0.155672
R1107 VTAIL.n238 VTAIL.n229 0.155672
R1108 VTAIL.n245 VTAIL.n229 0.155672
R1109 VTAIL.n246 VTAIL.n245 0.155672
R1110 VTAIL.n246 VTAIL.n225 0.155672
R1111 VTAIL.n253 VTAIL.n225 0.155672
R1112 VTAIL.n14 VTAIL.n13 0.155672
R1113 VTAIL.n14 VTAIL.n5 0.155672
R1114 VTAIL.n21 VTAIL.n5 0.155672
R1115 VTAIL.n22 VTAIL.n21 0.155672
R1116 VTAIL.n22 VTAIL.n1 0.155672
R1117 VTAIL.n29 VTAIL.n1 0.155672
R1118 VTAIL.n46 VTAIL.n45 0.155672
R1119 VTAIL.n46 VTAIL.n37 0.155672
R1120 VTAIL.n53 VTAIL.n37 0.155672
R1121 VTAIL.n54 VTAIL.n53 0.155672
R1122 VTAIL.n54 VTAIL.n33 0.155672
R1123 VTAIL.n61 VTAIL.n33 0.155672
R1124 VTAIL.n78 VTAIL.n77 0.155672
R1125 VTAIL.n78 VTAIL.n69 0.155672
R1126 VTAIL.n85 VTAIL.n69 0.155672
R1127 VTAIL.n86 VTAIL.n85 0.155672
R1128 VTAIL.n86 VTAIL.n65 0.155672
R1129 VTAIL.n93 VTAIL.n65 0.155672
R1130 VTAIL.n221 VTAIL.n193 0.155672
R1131 VTAIL.n214 VTAIL.n193 0.155672
R1132 VTAIL.n214 VTAIL.n213 0.155672
R1133 VTAIL.n213 VTAIL.n197 0.155672
R1134 VTAIL.n206 VTAIL.n197 0.155672
R1135 VTAIL.n206 VTAIL.n205 0.155672
R1136 VTAIL.n189 VTAIL.n161 0.155672
R1137 VTAIL.n182 VTAIL.n161 0.155672
R1138 VTAIL.n182 VTAIL.n181 0.155672
R1139 VTAIL.n181 VTAIL.n165 0.155672
R1140 VTAIL.n174 VTAIL.n165 0.155672
R1141 VTAIL.n174 VTAIL.n173 0.155672
R1142 VTAIL.n157 VTAIL.n129 0.155672
R1143 VTAIL.n150 VTAIL.n129 0.155672
R1144 VTAIL.n150 VTAIL.n149 0.155672
R1145 VTAIL.n149 VTAIL.n133 0.155672
R1146 VTAIL.n142 VTAIL.n133 0.155672
R1147 VTAIL.n142 VTAIL.n141 0.155672
R1148 VTAIL.n125 VTAIL.n97 0.155672
R1149 VTAIL.n118 VTAIL.n97 0.155672
R1150 VTAIL.n118 VTAIL.n117 0.155672
R1151 VTAIL.n117 VTAIL.n101 0.155672
R1152 VTAIL.n110 VTAIL.n101 0.155672
R1153 VTAIL.n110 VTAIL.n109 0.155672
R1154 VDD1 VDD1.n1 130.297
R1155 VDD1 VDD1.n0 94.4856
R1156 VDD1.n0 VDD1.t1 5.32047
R1157 VDD1.n0 VDD1.t0 5.32047
R1158 VDD1.n1 VDD1.t2 5.32047
R1159 VDD1.n1 VDD1.t3 5.32047
R1160 VN.n0 VN.t2 105.379
R1161 VN.n1 VN.t0 105.379
R1162 VN.n0 VN.t3 104.826
R1163 VN.n1 VN.t1 104.826
R1164 VN VN.n1 47.5418
R1165 VN VN.n0 6.79559
R1166 VDD2.n2 VDD2.n0 129.772
R1167 VDD2.n2 VDD2.n1 94.4274
R1168 VDD2.n1 VDD2.t2 5.32047
R1169 VDD2.n1 VDD2.t3 5.32047
R1170 VDD2.n0 VDD2.t1 5.32047
R1171 VDD2.n0 VDD2.t0 5.32047
R1172 VDD2 VDD2.n2 0.0586897
C0 B VDD2 1.06593f
C1 VDD2 w_n2446_n2190# 1.25154f
C2 B VP 1.46455f
C3 VP w_n2446_n2190# 4.24993f
C4 VN VTAIL 2.67439f
C5 VN VDD1 0.148703f
C6 VTAIL VDD1 3.85533f
C7 B w_n2446_n2190# 7.02436f
C8 VN VDD2 2.47761f
C9 VDD2 VTAIL 3.90639f
C10 VDD2 VDD1 0.916374f
C11 VN VP 4.75855f
C12 VP VTAIL 2.6885f
C13 VP VDD1 2.69282f
C14 VN B 0.946909f
C15 VN w_n2446_n2190# 3.93667f
C16 B VTAIL 2.84102f
C17 VP VDD2 0.364526f
C18 VTAIL w_n2446_n2190# 2.62009f
C19 B VDD1 1.02149f
C20 w_n2446_n2190# VDD1 1.20594f
C21 VDD2 VSUBS 0.722942f
C22 VDD1 VSUBS 4.708567f
C23 VTAIL VSUBS 0.669378f
C24 VN VSUBS 5.05861f
C25 VP VSUBS 1.730252f
C26 B VSUBS 3.369387f
C27 w_n2446_n2190# VSUBS 66.834496f
C28 VDD2.t1 VSUBS 0.132025f
C29 VDD2.t0 VSUBS 0.132025f
C30 VDD2.n0 VSUBS 1.28994f
C31 VDD2.t2 VSUBS 0.132025f
C32 VDD2.t3 VSUBS 0.132025f
C33 VDD2.n1 VSUBS 0.881932f
C34 VDD2.n2 VSUBS 3.50729f
C35 VN.t2 VSUBS 1.81553f
C36 VN.t3 VSUBS 1.81129f
C37 VN.n0 VSUBS 1.21187f
C38 VN.t0 VSUBS 1.81553f
C39 VN.t1 VSUBS 1.81129f
C40 VN.n1 VSUBS 3.00465f
C41 VDD1.t1 VSUBS 0.134036f
C42 VDD1.t0 VSUBS 0.134036f
C43 VDD1.n0 VSUBS 0.895768f
C44 VDD1.t2 VSUBS 0.134036f
C45 VDD1.t3 VSUBS 0.134036f
C46 VDD1.n1 VSUBS 1.3295f
C47 VTAIL.n0 VSUBS 0.030646f
C48 VTAIL.n1 VSUBS 0.026854f
C49 VTAIL.n2 VSUBS 0.01443f
C50 VTAIL.n3 VSUBS 0.034107f
C51 VTAIL.n4 VSUBS 0.015279f
C52 VTAIL.n5 VSUBS 0.026854f
C53 VTAIL.n6 VSUBS 0.01443f
C54 VTAIL.n7 VSUBS 0.034107f
C55 VTAIL.n8 VSUBS 0.015279f
C56 VTAIL.n9 VSUBS 0.119764f
C57 VTAIL.t3 VSUBS 0.073352f
C58 VTAIL.n10 VSUBS 0.02558f
C59 VTAIL.n11 VSUBS 0.021686f
C60 VTAIL.n12 VSUBS 0.01443f
C61 VTAIL.n13 VSUBS 0.629095f
C62 VTAIL.n14 VSUBS 0.026854f
C63 VTAIL.n15 VSUBS 0.01443f
C64 VTAIL.n16 VSUBS 0.015279f
C65 VTAIL.n17 VSUBS 0.034107f
C66 VTAIL.n18 VSUBS 0.034107f
C67 VTAIL.n19 VSUBS 0.015279f
C68 VTAIL.n20 VSUBS 0.01443f
C69 VTAIL.n21 VSUBS 0.026854f
C70 VTAIL.n22 VSUBS 0.026854f
C71 VTAIL.n23 VSUBS 0.01443f
C72 VTAIL.n24 VSUBS 0.015279f
C73 VTAIL.n25 VSUBS 0.034107f
C74 VTAIL.n26 VSUBS 0.086452f
C75 VTAIL.n27 VSUBS 0.015279f
C76 VTAIL.n28 VSUBS 0.01443f
C77 VTAIL.n29 VSUBS 0.066106f
C78 VTAIL.n30 VSUBS 0.043769f
C79 VTAIL.n31 VSUBS 0.162654f
C80 VTAIL.n32 VSUBS 0.030646f
C81 VTAIL.n33 VSUBS 0.026854f
C82 VTAIL.n34 VSUBS 0.01443f
C83 VTAIL.n35 VSUBS 0.034107f
C84 VTAIL.n36 VSUBS 0.015279f
C85 VTAIL.n37 VSUBS 0.026854f
C86 VTAIL.n38 VSUBS 0.01443f
C87 VTAIL.n39 VSUBS 0.034107f
C88 VTAIL.n40 VSUBS 0.015279f
C89 VTAIL.n41 VSUBS 0.119764f
C90 VTAIL.t6 VSUBS 0.073352f
C91 VTAIL.n42 VSUBS 0.02558f
C92 VTAIL.n43 VSUBS 0.021686f
C93 VTAIL.n44 VSUBS 0.01443f
C94 VTAIL.n45 VSUBS 0.629095f
C95 VTAIL.n46 VSUBS 0.026854f
C96 VTAIL.n47 VSUBS 0.01443f
C97 VTAIL.n48 VSUBS 0.015279f
C98 VTAIL.n49 VSUBS 0.034107f
C99 VTAIL.n50 VSUBS 0.034107f
C100 VTAIL.n51 VSUBS 0.015279f
C101 VTAIL.n52 VSUBS 0.01443f
C102 VTAIL.n53 VSUBS 0.026854f
C103 VTAIL.n54 VSUBS 0.026854f
C104 VTAIL.n55 VSUBS 0.01443f
C105 VTAIL.n56 VSUBS 0.015279f
C106 VTAIL.n57 VSUBS 0.034107f
C107 VTAIL.n58 VSUBS 0.086452f
C108 VTAIL.n59 VSUBS 0.015279f
C109 VTAIL.n60 VSUBS 0.01443f
C110 VTAIL.n61 VSUBS 0.066106f
C111 VTAIL.n62 VSUBS 0.043769f
C112 VTAIL.n63 VSUBS 0.249369f
C113 VTAIL.n64 VSUBS 0.030646f
C114 VTAIL.n65 VSUBS 0.026854f
C115 VTAIL.n66 VSUBS 0.01443f
C116 VTAIL.n67 VSUBS 0.034107f
C117 VTAIL.n68 VSUBS 0.015279f
C118 VTAIL.n69 VSUBS 0.026854f
C119 VTAIL.n70 VSUBS 0.01443f
C120 VTAIL.n71 VSUBS 0.034107f
C121 VTAIL.n72 VSUBS 0.015279f
C122 VTAIL.n73 VSUBS 0.119764f
C123 VTAIL.t4 VSUBS 0.073352f
C124 VTAIL.n74 VSUBS 0.02558f
C125 VTAIL.n75 VSUBS 0.021686f
C126 VTAIL.n76 VSUBS 0.01443f
C127 VTAIL.n77 VSUBS 0.629095f
C128 VTAIL.n78 VSUBS 0.026854f
C129 VTAIL.n79 VSUBS 0.01443f
C130 VTAIL.n80 VSUBS 0.015279f
C131 VTAIL.n81 VSUBS 0.034107f
C132 VTAIL.n82 VSUBS 0.034107f
C133 VTAIL.n83 VSUBS 0.015279f
C134 VTAIL.n84 VSUBS 0.01443f
C135 VTAIL.n85 VSUBS 0.026854f
C136 VTAIL.n86 VSUBS 0.026854f
C137 VTAIL.n87 VSUBS 0.01443f
C138 VTAIL.n88 VSUBS 0.015279f
C139 VTAIL.n89 VSUBS 0.034107f
C140 VTAIL.n90 VSUBS 0.086452f
C141 VTAIL.n91 VSUBS 0.015279f
C142 VTAIL.n92 VSUBS 0.01443f
C143 VTAIL.n93 VSUBS 0.066106f
C144 VTAIL.n94 VSUBS 0.043769f
C145 VTAIL.n95 VSUBS 1.21276f
C146 VTAIL.n96 VSUBS 0.030646f
C147 VTAIL.n97 VSUBS 0.026854f
C148 VTAIL.n98 VSUBS 0.01443f
C149 VTAIL.n99 VSUBS 0.034107f
C150 VTAIL.n100 VSUBS 0.015279f
C151 VTAIL.n101 VSUBS 0.026854f
C152 VTAIL.n102 VSUBS 0.01443f
C153 VTAIL.n103 VSUBS 0.034107f
C154 VTAIL.n104 VSUBS 0.015279f
C155 VTAIL.n105 VSUBS 0.119764f
C156 VTAIL.t1 VSUBS 0.073352f
C157 VTAIL.n106 VSUBS 0.02558f
C158 VTAIL.n107 VSUBS 0.021686f
C159 VTAIL.n108 VSUBS 0.01443f
C160 VTAIL.n109 VSUBS 0.629095f
C161 VTAIL.n110 VSUBS 0.026854f
C162 VTAIL.n111 VSUBS 0.01443f
C163 VTAIL.n112 VSUBS 0.015279f
C164 VTAIL.n113 VSUBS 0.034107f
C165 VTAIL.n114 VSUBS 0.034107f
C166 VTAIL.n115 VSUBS 0.015279f
C167 VTAIL.n116 VSUBS 0.01443f
C168 VTAIL.n117 VSUBS 0.026854f
C169 VTAIL.n118 VSUBS 0.026854f
C170 VTAIL.n119 VSUBS 0.01443f
C171 VTAIL.n120 VSUBS 0.015279f
C172 VTAIL.n121 VSUBS 0.034107f
C173 VTAIL.n122 VSUBS 0.086452f
C174 VTAIL.n123 VSUBS 0.015279f
C175 VTAIL.n124 VSUBS 0.01443f
C176 VTAIL.n125 VSUBS 0.066106f
C177 VTAIL.n126 VSUBS 0.043769f
C178 VTAIL.n127 VSUBS 1.21276f
C179 VTAIL.n128 VSUBS 0.030646f
C180 VTAIL.n129 VSUBS 0.026854f
C181 VTAIL.n130 VSUBS 0.01443f
C182 VTAIL.n131 VSUBS 0.034107f
C183 VTAIL.n132 VSUBS 0.015279f
C184 VTAIL.n133 VSUBS 0.026854f
C185 VTAIL.n134 VSUBS 0.01443f
C186 VTAIL.n135 VSUBS 0.034107f
C187 VTAIL.n136 VSUBS 0.015279f
C188 VTAIL.n137 VSUBS 0.119764f
C189 VTAIL.t0 VSUBS 0.073352f
C190 VTAIL.n138 VSUBS 0.02558f
C191 VTAIL.n139 VSUBS 0.021686f
C192 VTAIL.n140 VSUBS 0.01443f
C193 VTAIL.n141 VSUBS 0.629095f
C194 VTAIL.n142 VSUBS 0.026854f
C195 VTAIL.n143 VSUBS 0.01443f
C196 VTAIL.n144 VSUBS 0.015279f
C197 VTAIL.n145 VSUBS 0.034107f
C198 VTAIL.n146 VSUBS 0.034107f
C199 VTAIL.n147 VSUBS 0.015279f
C200 VTAIL.n148 VSUBS 0.01443f
C201 VTAIL.n149 VSUBS 0.026854f
C202 VTAIL.n150 VSUBS 0.026854f
C203 VTAIL.n151 VSUBS 0.01443f
C204 VTAIL.n152 VSUBS 0.015279f
C205 VTAIL.n153 VSUBS 0.034107f
C206 VTAIL.n154 VSUBS 0.086452f
C207 VTAIL.n155 VSUBS 0.015279f
C208 VTAIL.n156 VSUBS 0.01443f
C209 VTAIL.n157 VSUBS 0.066106f
C210 VTAIL.n158 VSUBS 0.043769f
C211 VTAIL.n159 VSUBS 0.249369f
C212 VTAIL.n160 VSUBS 0.030646f
C213 VTAIL.n161 VSUBS 0.026854f
C214 VTAIL.n162 VSUBS 0.01443f
C215 VTAIL.n163 VSUBS 0.034107f
C216 VTAIL.n164 VSUBS 0.015279f
C217 VTAIL.n165 VSUBS 0.026854f
C218 VTAIL.n166 VSUBS 0.01443f
C219 VTAIL.n167 VSUBS 0.034107f
C220 VTAIL.n168 VSUBS 0.015279f
C221 VTAIL.n169 VSUBS 0.119764f
C222 VTAIL.t7 VSUBS 0.073352f
C223 VTAIL.n170 VSUBS 0.02558f
C224 VTAIL.n171 VSUBS 0.021686f
C225 VTAIL.n172 VSUBS 0.01443f
C226 VTAIL.n173 VSUBS 0.629095f
C227 VTAIL.n174 VSUBS 0.026854f
C228 VTAIL.n175 VSUBS 0.01443f
C229 VTAIL.n176 VSUBS 0.015279f
C230 VTAIL.n177 VSUBS 0.034107f
C231 VTAIL.n178 VSUBS 0.034107f
C232 VTAIL.n179 VSUBS 0.015279f
C233 VTAIL.n180 VSUBS 0.01443f
C234 VTAIL.n181 VSUBS 0.026854f
C235 VTAIL.n182 VSUBS 0.026854f
C236 VTAIL.n183 VSUBS 0.01443f
C237 VTAIL.n184 VSUBS 0.015279f
C238 VTAIL.n185 VSUBS 0.034107f
C239 VTAIL.n186 VSUBS 0.086452f
C240 VTAIL.n187 VSUBS 0.015279f
C241 VTAIL.n188 VSUBS 0.01443f
C242 VTAIL.n189 VSUBS 0.066106f
C243 VTAIL.n190 VSUBS 0.043769f
C244 VTAIL.n191 VSUBS 0.249369f
C245 VTAIL.n192 VSUBS 0.030646f
C246 VTAIL.n193 VSUBS 0.026854f
C247 VTAIL.n194 VSUBS 0.01443f
C248 VTAIL.n195 VSUBS 0.034107f
C249 VTAIL.n196 VSUBS 0.015279f
C250 VTAIL.n197 VSUBS 0.026854f
C251 VTAIL.n198 VSUBS 0.01443f
C252 VTAIL.n199 VSUBS 0.034107f
C253 VTAIL.n200 VSUBS 0.015279f
C254 VTAIL.n201 VSUBS 0.119764f
C255 VTAIL.t5 VSUBS 0.073352f
C256 VTAIL.n202 VSUBS 0.02558f
C257 VTAIL.n203 VSUBS 0.021686f
C258 VTAIL.n204 VSUBS 0.01443f
C259 VTAIL.n205 VSUBS 0.629095f
C260 VTAIL.n206 VSUBS 0.026854f
C261 VTAIL.n207 VSUBS 0.01443f
C262 VTAIL.n208 VSUBS 0.015279f
C263 VTAIL.n209 VSUBS 0.034107f
C264 VTAIL.n210 VSUBS 0.034107f
C265 VTAIL.n211 VSUBS 0.015279f
C266 VTAIL.n212 VSUBS 0.01443f
C267 VTAIL.n213 VSUBS 0.026854f
C268 VTAIL.n214 VSUBS 0.026854f
C269 VTAIL.n215 VSUBS 0.01443f
C270 VTAIL.n216 VSUBS 0.015279f
C271 VTAIL.n217 VSUBS 0.034107f
C272 VTAIL.n218 VSUBS 0.086452f
C273 VTAIL.n219 VSUBS 0.015279f
C274 VTAIL.n220 VSUBS 0.01443f
C275 VTAIL.n221 VSUBS 0.066106f
C276 VTAIL.n222 VSUBS 0.043769f
C277 VTAIL.n223 VSUBS 1.21276f
C278 VTAIL.n224 VSUBS 0.030646f
C279 VTAIL.n225 VSUBS 0.026854f
C280 VTAIL.n226 VSUBS 0.01443f
C281 VTAIL.n227 VSUBS 0.034107f
C282 VTAIL.n228 VSUBS 0.015279f
C283 VTAIL.n229 VSUBS 0.026854f
C284 VTAIL.n230 VSUBS 0.01443f
C285 VTAIL.n231 VSUBS 0.034107f
C286 VTAIL.n232 VSUBS 0.015279f
C287 VTAIL.n233 VSUBS 0.119764f
C288 VTAIL.t2 VSUBS 0.073352f
C289 VTAIL.n234 VSUBS 0.02558f
C290 VTAIL.n235 VSUBS 0.021686f
C291 VTAIL.n236 VSUBS 0.01443f
C292 VTAIL.n237 VSUBS 0.629095f
C293 VTAIL.n238 VSUBS 0.026854f
C294 VTAIL.n239 VSUBS 0.01443f
C295 VTAIL.n240 VSUBS 0.015279f
C296 VTAIL.n241 VSUBS 0.034107f
C297 VTAIL.n242 VSUBS 0.034107f
C298 VTAIL.n243 VSUBS 0.015279f
C299 VTAIL.n244 VSUBS 0.01443f
C300 VTAIL.n245 VSUBS 0.026854f
C301 VTAIL.n246 VSUBS 0.026854f
C302 VTAIL.n247 VSUBS 0.01443f
C303 VTAIL.n248 VSUBS 0.015279f
C304 VTAIL.n249 VSUBS 0.034107f
C305 VTAIL.n250 VSUBS 0.086452f
C306 VTAIL.n251 VSUBS 0.015279f
C307 VTAIL.n252 VSUBS 0.01443f
C308 VTAIL.n253 VSUBS 0.066106f
C309 VTAIL.n254 VSUBS 0.043769f
C310 VTAIL.n255 VSUBS 1.11597f
C311 VP.n0 VSUBS 0.060832f
C312 VP.t0 VSUBS 1.59103f
C313 VP.n1 VSUBS 0.067357f
C314 VP.t3 VSUBS 1.88489f
C315 VP.t2 VSUBS 1.88931f
C316 VP.n2 VSUBS 3.10287f
C317 VP.n3 VSUBS 2.17954f
C318 VP.t1 VSUBS 1.59103f
C319 VP.n4 VSUBS 0.764974f
C320 VP.n5 VSUBS 0.084296f
C321 VP.n6 VSUBS 0.060832f
C322 VP.n7 VSUBS 0.04614f
C323 VP.n8 VSUBS 0.04614f
C324 VP.n9 VSUBS 0.067357f
C325 VP.n10 VSUBS 0.084296f
C326 VP.n11 VSUBS 0.764974f
C327 VP.n12 VSUBS 0.051229f
C328 B.n0 VSUBS 0.00529f
C329 B.n1 VSUBS 0.00529f
C330 B.n2 VSUBS 0.008366f
C331 B.n3 VSUBS 0.008366f
C332 B.n4 VSUBS 0.008366f
C333 B.n5 VSUBS 0.008366f
C334 B.n6 VSUBS 0.008366f
C335 B.n7 VSUBS 0.008366f
C336 B.n8 VSUBS 0.008366f
C337 B.n9 VSUBS 0.008366f
C338 B.n10 VSUBS 0.008366f
C339 B.n11 VSUBS 0.008366f
C340 B.n12 VSUBS 0.008366f
C341 B.n13 VSUBS 0.008366f
C342 B.n14 VSUBS 0.008366f
C343 B.n15 VSUBS 0.008366f
C344 B.n16 VSUBS 0.008366f
C345 B.n17 VSUBS 0.019333f
C346 B.n18 VSUBS 0.008366f
C347 B.n19 VSUBS 0.008366f
C348 B.n20 VSUBS 0.008366f
C349 B.n21 VSUBS 0.008366f
C350 B.n22 VSUBS 0.008366f
C351 B.n23 VSUBS 0.008366f
C352 B.n24 VSUBS 0.008366f
C353 B.n25 VSUBS 0.008366f
C354 B.n26 VSUBS 0.008366f
C355 B.n27 VSUBS 0.008366f
C356 B.n28 VSUBS 0.008366f
C357 B.n29 VSUBS 0.008366f
C358 B.t2 VSUBS 0.109543f
C359 B.t1 VSUBS 0.135775f
C360 B.t0 VSUBS 0.727364f
C361 B.n30 VSUBS 0.233205f
C362 B.n31 VSUBS 0.186801f
C363 B.n32 VSUBS 0.008366f
C364 B.n33 VSUBS 0.008366f
C365 B.n34 VSUBS 0.008366f
C366 B.n35 VSUBS 0.008366f
C367 B.t11 VSUBS 0.109545f
C368 B.t10 VSUBS 0.135777f
C369 B.t9 VSUBS 0.727364f
C370 B.n36 VSUBS 0.233204f
C371 B.n37 VSUBS 0.186799f
C372 B.n38 VSUBS 0.019383f
C373 B.n39 VSUBS 0.008366f
C374 B.n40 VSUBS 0.008366f
C375 B.n41 VSUBS 0.008366f
C376 B.n42 VSUBS 0.008366f
C377 B.n43 VSUBS 0.008366f
C378 B.n44 VSUBS 0.008366f
C379 B.n45 VSUBS 0.008366f
C380 B.n46 VSUBS 0.008366f
C381 B.n47 VSUBS 0.008366f
C382 B.n48 VSUBS 0.008366f
C383 B.n49 VSUBS 0.008366f
C384 B.n50 VSUBS 0.018304f
C385 B.n51 VSUBS 0.008366f
C386 B.n52 VSUBS 0.008366f
C387 B.n53 VSUBS 0.008366f
C388 B.n54 VSUBS 0.008366f
C389 B.n55 VSUBS 0.008366f
C390 B.n56 VSUBS 0.008366f
C391 B.n57 VSUBS 0.008366f
C392 B.n58 VSUBS 0.008366f
C393 B.n59 VSUBS 0.008366f
C394 B.n60 VSUBS 0.008366f
C395 B.n61 VSUBS 0.008366f
C396 B.n62 VSUBS 0.008366f
C397 B.n63 VSUBS 0.008366f
C398 B.n64 VSUBS 0.008366f
C399 B.n65 VSUBS 0.008366f
C400 B.n66 VSUBS 0.008366f
C401 B.n67 VSUBS 0.008366f
C402 B.n68 VSUBS 0.008366f
C403 B.n69 VSUBS 0.008366f
C404 B.n70 VSUBS 0.008366f
C405 B.n71 VSUBS 0.008366f
C406 B.n72 VSUBS 0.008366f
C407 B.n73 VSUBS 0.008366f
C408 B.n74 VSUBS 0.008366f
C409 B.n75 VSUBS 0.008366f
C410 B.n76 VSUBS 0.008366f
C411 B.n77 VSUBS 0.008366f
C412 B.n78 VSUBS 0.008366f
C413 B.n79 VSUBS 0.008366f
C414 B.n80 VSUBS 0.008366f
C415 B.n81 VSUBS 0.019333f
C416 B.n82 VSUBS 0.008366f
C417 B.n83 VSUBS 0.008366f
C418 B.n84 VSUBS 0.008366f
C419 B.n85 VSUBS 0.008366f
C420 B.n86 VSUBS 0.008366f
C421 B.n87 VSUBS 0.008366f
C422 B.n88 VSUBS 0.008366f
C423 B.n89 VSUBS 0.008366f
C424 B.n90 VSUBS 0.008366f
C425 B.n91 VSUBS 0.008366f
C426 B.n92 VSUBS 0.008366f
C427 B.n93 VSUBS 0.008366f
C428 B.t7 VSUBS 0.109545f
C429 B.t8 VSUBS 0.135777f
C430 B.t6 VSUBS 0.727364f
C431 B.n94 VSUBS 0.233204f
C432 B.n95 VSUBS 0.186799f
C433 B.n96 VSUBS 0.008366f
C434 B.n97 VSUBS 0.008366f
C435 B.n98 VSUBS 0.008366f
C436 B.n99 VSUBS 0.008366f
C437 B.t4 VSUBS 0.109543f
C438 B.t5 VSUBS 0.135775f
C439 B.t3 VSUBS 0.727364f
C440 B.n100 VSUBS 0.233205f
C441 B.n101 VSUBS 0.186801f
C442 B.n102 VSUBS 0.019383f
C443 B.n103 VSUBS 0.008366f
C444 B.n104 VSUBS 0.008366f
C445 B.n105 VSUBS 0.008366f
C446 B.n106 VSUBS 0.008366f
C447 B.n107 VSUBS 0.008366f
C448 B.n108 VSUBS 0.008366f
C449 B.n109 VSUBS 0.008366f
C450 B.n110 VSUBS 0.008366f
C451 B.n111 VSUBS 0.008366f
C452 B.n112 VSUBS 0.008366f
C453 B.n113 VSUBS 0.008366f
C454 B.n114 VSUBS 0.019333f
C455 B.n115 VSUBS 0.008366f
C456 B.n116 VSUBS 0.008366f
C457 B.n117 VSUBS 0.008366f
C458 B.n118 VSUBS 0.008366f
C459 B.n119 VSUBS 0.008366f
C460 B.n120 VSUBS 0.008366f
C461 B.n121 VSUBS 0.008366f
C462 B.n122 VSUBS 0.008366f
C463 B.n123 VSUBS 0.008366f
C464 B.n124 VSUBS 0.008366f
C465 B.n125 VSUBS 0.008366f
C466 B.n126 VSUBS 0.008366f
C467 B.n127 VSUBS 0.008366f
C468 B.n128 VSUBS 0.008366f
C469 B.n129 VSUBS 0.008366f
C470 B.n130 VSUBS 0.008366f
C471 B.n131 VSUBS 0.008366f
C472 B.n132 VSUBS 0.008366f
C473 B.n133 VSUBS 0.008366f
C474 B.n134 VSUBS 0.008366f
C475 B.n135 VSUBS 0.008366f
C476 B.n136 VSUBS 0.008366f
C477 B.n137 VSUBS 0.008366f
C478 B.n138 VSUBS 0.008366f
C479 B.n139 VSUBS 0.008366f
C480 B.n140 VSUBS 0.008366f
C481 B.n141 VSUBS 0.008366f
C482 B.n142 VSUBS 0.008366f
C483 B.n143 VSUBS 0.008366f
C484 B.n144 VSUBS 0.008366f
C485 B.n145 VSUBS 0.008366f
C486 B.n146 VSUBS 0.008366f
C487 B.n147 VSUBS 0.008366f
C488 B.n148 VSUBS 0.008366f
C489 B.n149 VSUBS 0.008366f
C490 B.n150 VSUBS 0.008366f
C491 B.n151 VSUBS 0.008366f
C492 B.n152 VSUBS 0.008366f
C493 B.n153 VSUBS 0.008366f
C494 B.n154 VSUBS 0.008366f
C495 B.n155 VSUBS 0.008366f
C496 B.n156 VSUBS 0.008366f
C497 B.n157 VSUBS 0.008366f
C498 B.n158 VSUBS 0.008366f
C499 B.n159 VSUBS 0.008366f
C500 B.n160 VSUBS 0.008366f
C501 B.n161 VSUBS 0.008366f
C502 B.n162 VSUBS 0.008366f
C503 B.n163 VSUBS 0.008366f
C504 B.n164 VSUBS 0.008366f
C505 B.n165 VSUBS 0.008366f
C506 B.n166 VSUBS 0.008366f
C507 B.n167 VSUBS 0.008366f
C508 B.n168 VSUBS 0.008366f
C509 B.n169 VSUBS 0.008366f
C510 B.n170 VSUBS 0.008366f
C511 B.n171 VSUBS 0.018806f
C512 B.n172 VSUBS 0.018806f
C513 B.n173 VSUBS 0.019333f
C514 B.n174 VSUBS 0.008366f
C515 B.n175 VSUBS 0.008366f
C516 B.n176 VSUBS 0.008366f
C517 B.n177 VSUBS 0.008366f
C518 B.n178 VSUBS 0.008366f
C519 B.n179 VSUBS 0.008366f
C520 B.n180 VSUBS 0.008366f
C521 B.n181 VSUBS 0.008366f
C522 B.n182 VSUBS 0.008366f
C523 B.n183 VSUBS 0.008366f
C524 B.n184 VSUBS 0.008366f
C525 B.n185 VSUBS 0.008366f
C526 B.n186 VSUBS 0.008366f
C527 B.n187 VSUBS 0.008366f
C528 B.n188 VSUBS 0.008366f
C529 B.n189 VSUBS 0.008366f
C530 B.n190 VSUBS 0.008366f
C531 B.n191 VSUBS 0.008366f
C532 B.n192 VSUBS 0.008366f
C533 B.n193 VSUBS 0.008366f
C534 B.n194 VSUBS 0.008366f
C535 B.n195 VSUBS 0.008366f
C536 B.n196 VSUBS 0.008366f
C537 B.n197 VSUBS 0.008366f
C538 B.n198 VSUBS 0.008366f
C539 B.n199 VSUBS 0.008366f
C540 B.n200 VSUBS 0.008366f
C541 B.n201 VSUBS 0.008366f
C542 B.n202 VSUBS 0.008366f
C543 B.n203 VSUBS 0.008366f
C544 B.n204 VSUBS 0.008366f
C545 B.n205 VSUBS 0.008366f
C546 B.n206 VSUBS 0.008366f
C547 B.n207 VSUBS 0.007874f
C548 B.n208 VSUBS 0.008366f
C549 B.n209 VSUBS 0.008366f
C550 B.n210 VSUBS 0.004675f
C551 B.n211 VSUBS 0.008366f
C552 B.n212 VSUBS 0.008366f
C553 B.n213 VSUBS 0.008366f
C554 B.n214 VSUBS 0.008366f
C555 B.n215 VSUBS 0.008366f
C556 B.n216 VSUBS 0.008366f
C557 B.n217 VSUBS 0.008366f
C558 B.n218 VSUBS 0.008366f
C559 B.n219 VSUBS 0.008366f
C560 B.n220 VSUBS 0.008366f
C561 B.n221 VSUBS 0.008366f
C562 B.n222 VSUBS 0.008366f
C563 B.n223 VSUBS 0.004675f
C564 B.n224 VSUBS 0.019383f
C565 B.n225 VSUBS 0.007874f
C566 B.n226 VSUBS 0.008366f
C567 B.n227 VSUBS 0.008366f
C568 B.n228 VSUBS 0.008366f
C569 B.n229 VSUBS 0.008366f
C570 B.n230 VSUBS 0.008366f
C571 B.n231 VSUBS 0.008366f
C572 B.n232 VSUBS 0.008366f
C573 B.n233 VSUBS 0.008366f
C574 B.n234 VSUBS 0.008366f
C575 B.n235 VSUBS 0.008366f
C576 B.n236 VSUBS 0.008366f
C577 B.n237 VSUBS 0.008366f
C578 B.n238 VSUBS 0.008366f
C579 B.n239 VSUBS 0.008366f
C580 B.n240 VSUBS 0.008366f
C581 B.n241 VSUBS 0.008366f
C582 B.n242 VSUBS 0.008366f
C583 B.n243 VSUBS 0.008366f
C584 B.n244 VSUBS 0.008366f
C585 B.n245 VSUBS 0.008366f
C586 B.n246 VSUBS 0.008366f
C587 B.n247 VSUBS 0.008366f
C588 B.n248 VSUBS 0.008366f
C589 B.n249 VSUBS 0.008366f
C590 B.n250 VSUBS 0.008366f
C591 B.n251 VSUBS 0.008366f
C592 B.n252 VSUBS 0.008366f
C593 B.n253 VSUBS 0.008366f
C594 B.n254 VSUBS 0.008366f
C595 B.n255 VSUBS 0.008366f
C596 B.n256 VSUBS 0.008366f
C597 B.n257 VSUBS 0.008366f
C598 B.n258 VSUBS 0.008366f
C599 B.n259 VSUBS 0.008366f
C600 B.n260 VSUBS 0.019333f
C601 B.n261 VSUBS 0.018806f
C602 B.n262 VSUBS 0.018806f
C603 B.n263 VSUBS 0.008366f
C604 B.n264 VSUBS 0.008366f
C605 B.n265 VSUBS 0.008366f
C606 B.n266 VSUBS 0.008366f
C607 B.n267 VSUBS 0.008366f
C608 B.n268 VSUBS 0.008366f
C609 B.n269 VSUBS 0.008366f
C610 B.n270 VSUBS 0.008366f
C611 B.n271 VSUBS 0.008366f
C612 B.n272 VSUBS 0.008366f
C613 B.n273 VSUBS 0.008366f
C614 B.n274 VSUBS 0.008366f
C615 B.n275 VSUBS 0.008366f
C616 B.n276 VSUBS 0.008366f
C617 B.n277 VSUBS 0.008366f
C618 B.n278 VSUBS 0.008366f
C619 B.n279 VSUBS 0.008366f
C620 B.n280 VSUBS 0.008366f
C621 B.n281 VSUBS 0.008366f
C622 B.n282 VSUBS 0.008366f
C623 B.n283 VSUBS 0.008366f
C624 B.n284 VSUBS 0.008366f
C625 B.n285 VSUBS 0.008366f
C626 B.n286 VSUBS 0.008366f
C627 B.n287 VSUBS 0.008366f
C628 B.n288 VSUBS 0.008366f
C629 B.n289 VSUBS 0.008366f
C630 B.n290 VSUBS 0.008366f
C631 B.n291 VSUBS 0.008366f
C632 B.n292 VSUBS 0.008366f
C633 B.n293 VSUBS 0.008366f
C634 B.n294 VSUBS 0.008366f
C635 B.n295 VSUBS 0.008366f
C636 B.n296 VSUBS 0.008366f
C637 B.n297 VSUBS 0.008366f
C638 B.n298 VSUBS 0.008366f
C639 B.n299 VSUBS 0.008366f
C640 B.n300 VSUBS 0.008366f
C641 B.n301 VSUBS 0.008366f
C642 B.n302 VSUBS 0.008366f
C643 B.n303 VSUBS 0.008366f
C644 B.n304 VSUBS 0.008366f
C645 B.n305 VSUBS 0.008366f
C646 B.n306 VSUBS 0.008366f
C647 B.n307 VSUBS 0.008366f
C648 B.n308 VSUBS 0.008366f
C649 B.n309 VSUBS 0.008366f
C650 B.n310 VSUBS 0.008366f
C651 B.n311 VSUBS 0.008366f
C652 B.n312 VSUBS 0.008366f
C653 B.n313 VSUBS 0.008366f
C654 B.n314 VSUBS 0.008366f
C655 B.n315 VSUBS 0.008366f
C656 B.n316 VSUBS 0.008366f
C657 B.n317 VSUBS 0.008366f
C658 B.n318 VSUBS 0.008366f
C659 B.n319 VSUBS 0.008366f
C660 B.n320 VSUBS 0.008366f
C661 B.n321 VSUBS 0.008366f
C662 B.n322 VSUBS 0.008366f
C663 B.n323 VSUBS 0.008366f
C664 B.n324 VSUBS 0.008366f
C665 B.n325 VSUBS 0.008366f
C666 B.n326 VSUBS 0.008366f
C667 B.n327 VSUBS 0.008366f
C668 B.n328 VSUBS 0.008366f
C669 B.n329 VSUBS 0.008366f
C670 B.n330 VSUBS 0.008366f
C671 B.n331 VSUBS 0.008366f
C672 B.n332 VSUBS 0.008366f
C673 B.n333 VSUBS 0.008366f
C674 B.n334 VSUBS 0.008366f
C675 B.n335 VSUBS 0.008366f
C676 B.n336 VSUBS 0.008366f
C677 B.n337 VSUBS 0.008366f
C678 B.n338 VSUBS 0.008366f
C679 B.n339 VSUBS 0.008366f
C680 B.n340 VSUBS 0.008366f
C681 B.n341 VSUBS 0.008366f
C682 B.n342 VSUBS 0.008366f
C683 B.n343 VSUBS 0.008366f
C684 B.n344 VSUBS 0.008366f
C685 B.n345 VSUBS 0.008366f
C686 B.n346 VSUBS 0.008366f
C687 B.n347 VSUBS 0.008366f
C688 B.n348 VSUBS 0.008366f
C689 B.n349 VSUBS 0.008366f
C690 B.n350 VSUBS 0.008366f
C691 B.n351 VSUBS 0.019835f
C692 B.n352 VSUBS 0.018806f
C693 B.n353 VSUBS 0.019333f
C694 B.n354 VSUBS 0.008366f
C695 B.n355 VSUBS 0.008366f
C696 B.n356 VSUBS 0.008366f
C697 B.n357 VSUBS 0.008366f
C698 B.n358 VSUBS 0.008366f
C699 B.n359 VSUBS 0.008366f
C700 B.n360 VSUBS 0.008366f
C701 B.n361 VSUBS 0.008366f
C702 B.n362 VSUBS 0.008366f
C703 B.n363 VSUBS 0.008366f
C704 B.n364 VSUBS 0.008366f
C705 B.n365 VSUBS 0.008366f
C706 B.n366 VSUBS 0.008366f
C707 B.n367 VSUBS 0.008366f
C708 B.n368 VSUBS 0.008366f
C709 B.n369 VSUBS 0.008366f
C710 B.n370 VSUBS 0.008366f
C711 B.n371 VSUBS 0.008366f
C712 B.n372 VSUBS 0.008366f
C713 B.n373 VSUBS 0.008366f
C714 B.n374 VSUBS 0.008366f
C715 B.n375 VSUBS 0.008366f
C716 B.n376 VSUBS 0.008366f
C717 B.n377 VSUBS 0.008366f
C718 B.n378 VSUBS 0.008366f
C719 B.n379 VSUBS 0.008366f
C720 B.n380 VSUBS 0.008366f
C721 B.n381 VSUBS 0.008366f
C722 B.n382 VSUBS 0.008366f
C723 B.n383 VSUBS 0.008366f
C724 B.n384 VSUBS 0.008366f
C725 B.n385 VSUBS 0.008366f
C726 B.n386 VSUBS 0.008366f
C727 B.n387 VSUBS 0.007874f
C728 B.n388 VSUBS 0.008366f
C729 B.n389 VSUBS 0.008366f
C730 B.n390 VSUBS 0.004675f
C731 B.n391 VSUBS 0.008366f
C732 B.n392 VSUBS 0.008366f
C733 B.n393 VSUBS 0.008366f
C734 B.n394 VSUBS 0.008366f
C735 B.n395 VSUBS 0.008366f
C736 B.n396 VSUBS 0.008366f
C737 B.n397 VSUBS 0.008366f
C738 B.n398 VSUBS 0.008366f
C739 B.n399 VSUBS 0.008366f
C740 B.n400 VSUBS 0.008366f
C741 B.n401 VSUBS 0.008366f
C742 B.n402 VSUBS 0.008366f
C743 B.n403 VSUBS 0.004675f
C744 B.n404 VSUBS 0.019383f
C745 B.n405 VSUBS 0.007874f
C746 B.n406 VSUBS 0.008366f
C747 B.n407 VSUBS 0.008366f
C748 B.n408 VSUBS 0.008366f
C749 B.n409 VSUBS 0.008366f
C750 B.n410 VSUBS 0.008366f
C751 B.n411 VSUBS 0.008366f
C752 B.n412 VSUBS 0.008366f
C753 B.n413 VSUBS 0.008366f
C754 B.n414 VSUBS 0.008366f
C755 B.n415 VSUBS 0.008366f
C756 B.n416 VSUBS 0.008366f
C757 B.n417 VSUBS 0.008366f
C758 B.n418 VSUBS 0.008366f
C759 B.n419 VSUBS 0.008366f
C760 B.n420 VSUBS 0.008366f
C761 B.n421 VSUBS 0.008366f
C762 B.n422 VSUBS 0.008366f
C763 B.n423 VSUBS 0.008366f
C764 B.n424 VSUBS 0.008366f
C765 B.n425 VSUBS 0.008366f
C766 B.n426 VSUBS 0.008366f
C767 B.n427 VSUBS 0.008366f
C768 B.n428 VSUBS 0.008366f
C769 B.n429 VSUBS 0.008366f
C770 B.n430 VSUBS 0.008366f
C771 B.n431 VSUBS 0.008366f
C772 B.n432 VSUBS 0.008366f
C773 B.n433 VSUBS 0.008366f
C774 B.n434 VSUBS 0.008366f
C775 B.n435 VSUBS 0.008366f
C776 B.n436 VSUBS 0.008366f
C777 B.n437 VSUBS 0.008366f
C778 B.n438 VSUBS 0.008366f
C779 B.n439 VSUBS 0.008366f
C780 B.n440 VSUBS 0.019333f
C781 B.n441 VSUBS 0.018806f
C782 B.n442 VSUBS 0.018806f
C783 B.n443 VSUBS 0.008366f
C784 B.n444 VSUBS 0.008366f
C785 B.n445 VSUBS 0.008366f
C786 B.n446 VSUBS 0.008366f
C787 B.n447 VSUBS 0.008366f
C788 B.n448 VSUBS 0.008366f
C789 B.n449 VSUBS 0.008366f
C790 B.n450 VSUBS 0.008366f
C791 B.n451 VSUBS 0.008366f
C792 B.n452 VSUBS 0.008366f
C793 B.n453 VSUBS 0.008366f
C794 B.n454 VSUBS 0.008366f
C795 B.n455 VSUBS 0.008366f
C796 B.n456 VSUBS 0.008366f
C797 B.n457 VSUBS 0.008366f
C798 B.n458 VSUBS 0.008366f
C799 B.n459 VSUBS 0.008366f
C800 B.n460 VSUBS 0.008366f
C801 B.n461 VSUBS 0.008366f
C802 B.n462 VSUBS 0.008366f
C803 B.n463 VSUBS 0.008366f
C804 B.n464 VSUBS 0.008366f
C805 B.n465 VSUBS 0.008366f
C806 B.n466 VSUBS 0.008366f
C807 B.n467 VSUBS 0.008366f
C808 B.n468 VSUBS 0.008366f
C809 B.n469 VSUBS 0.008366f
C810 B.n470 VSUBS 0.008366f
C811 B.n471 VSUBS 0.008366f
C812 B.n472 VSUBS 0.008366f
C813 B.n473 VSUBS 0.008366f
C814 B.n474 VSUBS 0.008366f
C815 B.n475 VSUBS 0.008366f
C816 B.n476 VSUBS 0.008366f
C817 B.n477 VSUBS 0.008366f
C818 B.n478 VSUBS 0.008366f
C819 B.n479 VSUBS 0.008366f
C820 B.n480 VSUBS 0.008366f
C821 B.n481 VSUBS 0.008366f
C822 B.n482 VSUBS 0.008366f
C823 B.n483 VSUBS 0.008366f
C824 B.n484 VSUBS 0.008366f
C825 B.n485 VSUBS 0.008366f
C826 B.n486 VSUBS 0.008366f
C827 B.n487 VSUBS 0.018943f
.ends

