* NGSPICE file created from diff_pair_sample_0319.ext - technology: sky130A

.subckt diff_pair_sample_0319 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=0 ps=0 w=4.19 l=3.34
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=0 ps=0 w=4.19 l=3.34
X2 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=1.6341 ps=9.16 w=4.19 l=3.34
X3 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=1.6341 ps=9.16 w=4.19 l=3.34
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=0 ps=0 w=4.19 l=3.34
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=1.6341 ps=9.16 w=4.19 l=3.34
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=1.6341 ps=9.16 w=4.19 l=3.34
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6341 pd=9.16 as=0 ps=0 w=4.19 l=3.34
R0 B.n484 B.n483 585
R1 B.n485 B.n484 585
R2 B.n177 B.n80 585
R3 B.n176 B.n175 585
R4 B.n174 B.n173 585
R5 B.n172 B.n171 585
R6 B.n170 B.n169 585
R7 B.n168 B.n167 585
R8 B.n166 B.n165 585
R9 B.n164 B.n163 585
R10 B.n162 B.n161 585
R11 B.n160 B.n159 585
R12 B.n158 B.n157 585
R13 B.n156 B.n155 585
R14 B.n154 B.n153 585
R15 B.n152 B.n151 585
R16 B.n150 B.n149 585
R17 B.n148 B.n147 585
R18 B.n146 B.n145 585
R19 B.n144 B.n143 585
R20 B.n142 B.n141 585
R21 B.n140 B.n139 585
R22 B.n138 B.n137 585
R23 B.n136 B.n135 585
R24 B.n134 B.n133 585
R25 B.n132 B.n131 585
R26 B.n130 B.n129 585
R27 B.n128 B.n127 585
R28 B.n126 B.n125 585
R29 B.n123 B.n122 585
R30 B.n121 B.n120 585
R31 B.n119 B.n118 585
R32 B.n117 B.n116 585
R33 B.n115 B.n114 585
R34 B.n113 B.n112 585
R35 B.n111 B.n110 585
R36 B.n109 B.n108 585
R37 B.n107 B.n106 585
R38 B.n105 B.n104 585
R39 B.n103 B.n102 585
R40 B.n101 B.n100 585
R41 B.n99 B.n98 585
R42 B.n97 B.n96 585
R43 B.n95 B.n94 585
R44 B.n93 B.n92 585
R45 B.n91 B.n90 585
R46 B.n89 B.n88 585
R47 B.n87 B.n86 585
R48 B.n482 B.n56 585
R49 B.n486 B.n56 585
R50 B.n481 B.n55 585
R51 B.n487 B.n55 585
R52 B.n480 B.n479 585
R53 B.n479 B.n51 585
R54 B.n478 B.n50 585
R55 B.n493 B.n50 585
R56 B.n477 B.n49 585
R57 B.n494 B.n49 585
R58 B.n476 B.n48 585
R59 B.n495 B.n48 585
R60 B.n475 B.n474 585
R61 B.n474 B.n44 585
R62 B.n473 B.n43 585
R63 B.n501 B.n43 585
R64 B.n472 B.n42 585
R65 B.n502 B.n42 585
R66 B.n471 B.n41 585
R67 B.n503 B.n41 585
R68 B.n470 B.n469 585
R69 B.n469 B.n37 585
R70 B.n468 B.n36 585
R71 B.n509 B.n36 585
R72 B.n467 B.n35 585
R73 B.n510 B.n35 585
R74 B.n466 B.n34 585
R75 B.n511 B.n34 585
R76 B.n465 B.n464 585
R77 B.n464 B.n30 585
R78 B.n463 B.n29 585
R79 B.n517 B.n29 585
R80 B.n462 B.n28 585
R81 B.n518 B.n28 585
R82 B.n461 B.n27 585
R83 B.n519 B.n27 585
R84 B.n460 B.n459 585
R85 B.n459 B.n23 585
R86 B.n458 B.n22 585
R87 B.n525 B.n22 585
R88 B.n457 B.n21 585
R89 B.n526 B.n21 585
R90 B.n456 B.n20 585
R91 B.n527 B.n20 585
R92 B.n455 B.n454 585
R93 B.n454 B.n19 585
R94 B.n453 B.n15 585
R95 B.n533 B.n15 585
R96 B.n452 B.n14 585
R97 B.n534 B.n14 585
R98 B.n451 B.n13 585
R99 B.n535 B.n13 585
R100 B.n450 B.n449 585
R101 B.n449 B.n12 585
R102 B.n448 B.n447 585
R103 B.n448 B.n8 585
R104 B.n446 B.n7 585
R105 B.n542 B.n7 585
R106 B.n445 B.n6 585
R107 B.n543 B.n6 585
R108 B.n444 B.n5 585
R109 B.n544 B.n5 585
R110 B.n443 B.n442 585
R111 B.n442 B.n4 585
R112 B.n441 B.n178 585
R113 B.n441 B.n440 585
R114 B.n431 B.n179 585
R115 B.n180 B.n179 585
R116 B.n433 B.n432 585
R117 B.n434 B.n433 585
R118 B.n430 B.n185 585
R119 B.n185 B.n184 585
R120 B.n429 B.n428 585
R121 B.n428 B.n427 585
R122 B.n187 B.n186 585
R123 B.n420 B.n187 585
R124 B.n419 B.n418 585
R125 B.n421 B.n419 585
R126 B.n417 B.n192 585
R127 B.n192 B.n191 585
R128 B.n416 B.n415 585
R129 B.n415 B.n414 585
R130 B.n194 B.n193 585
R131 B.n195 B.n194 585
R132 B.n407 B.n406 585
R133 B.n408 B.n407 585
R134 B.n405 B.n200 585
R135 B.n200 B.n199 585
R136 B.n404 B.n403 585
R137 B.n403 B.n402 585
R138 B.n202 B.n201 585
R139 B.n203 B.n202 585
R140 B.n395 B.n394 585
R141 B.n396 B.n395 585
R142 B.n393 B.n208 585
R143 B.n208 B.n207 585
R144 B.n392 B.n391 585
R145 B.n391 B.n390 585
R146 B.n210 B.n209 585
R147 B.n211 B.n210 585
R148 B.n383 B.n382 585
R149 B.n384 B.n383 585
R150 B.n381 B.n215 585
R151 B.n219 B.n215 585
R152 B.n380 B.n379 585
R153 B.n379 B.n378 585
R154 B.n217 B.n216 585
R155 B.n218 B.n217 585
R156 B.n371 B.n370 585
R157 B.n372 B.n371 585
R158 B.n369 B.n224 585
R159 B.n224 B.n223 585
R160 B.n368 B.n367 585
R161 B.n367 B.n366 585
R162 B.n226 B.n225 585
R163 B.n227 B.n226 585
R164 B.n359 B.n358 585
R165 B.n360 B.n359 585
R166 B.n357 B.n232 585
R167 B.n232 B.n231 585
R168 B.n351 B.n350 585
R169 B.n349 B.n257 585
R170 B.n348 B.n256 585
R171 B.n353 B.n256 585
R172 B.n347 B.n346 585
R173 B.n345 B.n344 585
R174 B.n343 B.n342 585
R175 B.n341 B.n340 585
R176 B.n339 B.n338 585
R177 B.n337 B.n336 585
R178 B.n335 B.n334 585
R179 B.n333 B.n332 585
R180 B.n331 B.n330 585
R181 B.n329 B.n328 585
R182 B.n327 B.n326 585
R183 B.n325 B.n324 585
R184 B.n323 B.n322 585
R185 B.n321 B.n320 585
R186 B.n319 B.n318 585
R187 B.n317 B.n316 585
R188 B.n315 B.n314 585
R189 B.n313 B.n312 585
R190 B.n311 B.n310 585
R191 B.n309 B.n308 585
R192 B.n307 B.n306 585
R193 B.n305 B.n304 585
R194 B.n303 B.n302 585
R195 B.n301 B.n300 585
R196 B.n299 B.n298 585
R197 B.n296 B.n295 585
R198 B.n294 B.n293 585
R199 B.n292 B.n291 585
R200 B.n290 B.n289 585
R201 B.n288 B.n287 585
R202 B.n286 B.n285 585
R203 B.n284 B.n283 585
R204 B.n282 B.n281 585
R205 B.n280 B.n279 585
R206 B.n278 B.n277 585
R207 B.n276 B.n275 585
R208 B.n274 B.n273 585
R209 B.n272 B.n271 585
R210 B.n270 B.n269 585
R211 B.n268 B.n267 585
R212 B.n266 B.n265 585
R213 B.n264 B.n263 585
R214 B.n234 B.n233 585
R215 B.n356 B.n355 585
R216 B.n230 B.n229 585
R217 B.n231 B.n230 585
R218 B.n362 B.n361 585
R219 B.n361 B.n360 585
R220 B.n363 B.n228 585
R221 B.n228 B.n227 585
R222 B.n365 B.n364 585
R223 B.n366 B.n365 585
R224 B.n222 B.n221 585
R225 B.n223 B.n222 585
R226 B.n374 B.n373 585
R227 B.n373 B.n372 585
R228 B.n375 B.n220 585
R229 B.n220 B.n218 585
R230 B.n377 B.n376 585
R231 B.n378 B.n377 585
R232 B.n214 B.n213 585
R233 B.n219 B.n214 585
R234 B.n386 B.n385 585
R235 B.n385 B.n384 585
R236 B.n387 B.n212 585
R237 B.n212 B.n211 585
R238 B.n389 B.n388 585
R239 B.n390 B.n389 585
R240 B.n206 B.n205 585
R241 B.n207 B.n206 585
R242 B.n398 B.n397 585
R243 B.n397 B.n396 585
R244 B.n399 B.n204 585
R245 B.n204 B.n203 585
R246 B.n401 B.n400 585
R247 B.n402 B.n401 585
R248 B.n198 B.n197 585
R249 B.n199 B.n198 585
R250 B.n410 B.n409 585
R251 B.n409 B.n408 585
R252 B.n411 B.n196 585
R253 B.n196 B.n195 585
R254 B.n413 B.n412 585
R255 B.n414 B.n413 585
R256 B.n190 B.n189 585
R257 B.n191 B.n190 585
R258 B.n423 B.n422 585
R259 B.n422 B.n421 585
R260 B.n424 B.n188 585
R261 B.n420 B.n188 585
R262 B.n426 B.n425 585
R263 B.n427 B.n426 585
R264 B.n183 B.n182 585
R265 B.n184 B.n183 585
R266 B.n436 B.n435 585
R267 B.n435 B.n434 585
R268 B.n437 B.n181 585
R269 B.n181 B.n180 585
R270 B.n439 B.n438 585
R271 B.n440 B.n439 585
R272 B.n3 B.n0 585
R273 B.n4 B.n3 585
R274 B.n541 B.n1 585
R275 B.n542 B.n541 585
R276 B.n540 B.n539 585
R277 B.n540 B.n8 585
R278 B.n538 B.n9 585
R279 B.n12 B.n9 585
R280 B.n537 B.n536 585
R281 B.n536 B.n535 585
R282 B.n11 B.n10 585
R283 B.n534 B.n11 585
R284 B.n532 B.n531 585
R285 B.n533 B.n532 585
R286 B.n530 B.n16 585
R287 B.n19 B.n16 585
R288 B.n529 B.n528 585
R289 B.n528 B.n527 585
R290 B.n18 B.n17 585
R291 B.n526 B.n18 585
R292 B.n524 B.n523 585
R293 B.n525 B.n524 585
R294 B.n522 B.n24 585
R295 B.n24 B.n23 585
R296 B.n521 B.n520 585
R297 B.n520 B.n519 585
R298 B.n26 B.n25 585
R299 B.n518 B.n26 585
R300 B.n516 B.n515 585
R301 B.n517 B.n516 585
R302 B.n514 B.n31 585
R303 B.n31 B.n30 585
R304 B.n513 B.n512 585
R305 B.n512 B.n511 585
R306 B.n33 B.n32 585
R307 B.n510 B.n33 585
R308 B.n508 B.n507 585
R309 B.n509 B.n508 585
R310 B.n506 B.n38 585
R311 B.n38 B.n37 585
R312 B.n505 B.n504 585
R313 B.n504 B.n503 585
R314 B.n40 B.n39 585
R315 B.n502 B.n40 585
R316 B.n500 B.n499 585
R317 B.n501 B.n500 585
R318 B.n498 B.n45 585
R319 B.n45 B.n44 585
R320 B.n497 B.n496 585
R321 B.n496 B.n495 585
R322 B.n47 B.n46 585
R323 B.n494 B.n47 585
R324 B.n492 B.n491 585
R325 B.n493 B.n492 585
R326 B.n490 B.n52 585
R327 B.n52 B.n51 585
R328 B.n489 B.n488 585
R329 B.n488 B.n487 585
R330 B.n54 B.n53 585
R331 B.n486 B.n54 585
R332 B.n545 B.n544 585
R333 B.n543 B.n2 585
R334 B.n86 B.n54 521.33
R335 B.n484 B.n56 521.33
R336 B.n355 B.n232 521.33
R337 B.n351 B.n230 521.33
R338 B.n485 B.n79 256.663
R339 B.n485 B.n78 256.663
R340 B.n485 B.n77 256.663
R341 B.n485 B.n76 256.663
R342 B.n485 B.n75 256.663
R343 B.n485 B.n74 256.663
R344 B.n485 B.n73 256.663
R345 B.n485 B.n72 256.663
R346 B.n485 B.n71 256.663
R347 B.n485 B.n70 256.663
R348 B.n485 B.n69 256.663
R349 B.n485 B.n68 256.663
R350 B.n485 B.n67 256.663
R351 B.n485 B.n66 256.663
R352 B.n485 B.n65 256.663
R353 B.n485 B.n64 256.663
R354 B.n485 B.n63 256.663
R355 B.n485 B.n62 256.663
R356 B.n485 B.n61 256.663
R357 B.n485 B.n60 256.663
R358 B.n485 B.n59 256.663
R359 B.n485 B.n58 256.663
R360 B.n485 B.n57 256.663
R361 B.n353 B.n352 256.663
R362 B.n353 B.n235 256.663
R363 B.n353 B.n236 256.663
R364 B.n353 B.n237 256.663
R365 B.n353 B.n238 256.663
R366 B.n353 B.n239 256.663
R367 B.n353 B.n240 256.663
R368 B.n353 B.n241 256.663
R369 B.n353 B.n242 256.663
R370 B.n353 B.n243 256.663
R371 B.n353 B.n244 256.663
R372 B.n353 B.n245 256.663
R373 B.n353 B.n246 256.663
R374 B.n353 B.n247 256.663
R375 B.n353 B.n248 256.663
R376 B.n353 B.n249 256.663
R377 B.n353 B.n250 256.663
R378 B.n353 B.n251 256.663
R379 B.n353 B.n252 256.663
R380 B.n353 B.n253 256.663
R381 B.n353 B.n254 256.663
R382 B.n353 B.n255 256.663
R383 B.n354 B.n353 256.663
R384 B.n547 B.n546 256.663
R385 B.n84 B.t10 239.178
R386 B.n81 B.t2 239.178
R387 B.n261 B.t6 239.178
R388 B.n258 B.t13 239.178
R389 B.n90 B.n89 163.367
R390 B.n94 B.n93 163.367
R391 B.n98 B.n97 163.367
R392 B.n102 B.n101 163.367
R393 B.n106 B.n105 163.367
R394 B.n110 B.n109 163.367
R395 B.n114 B.n113 163.367
R396 B.n118 B.n117 163.367
R397 B.n122 B.n121 163.367
R398 B.n127 B.n126 163.367
R399 B.n131 B.n130 163.367
R400 B.n135 B.n134 163.367
R401 B.n139 B.n138 163.367
R402 B.n143 B.n142 163.367
R403 B.n147 B.n146 163.367
R404 B.n151 B.n150 163.367
R405 B.n155 B.n154 163.367
R406 B.n159 B.n158 163.367
R407 B.n163 B.n162 163.367
R408 B.n167 B.n166 163.367
R409 B.n171 B.n170 163.367
R410 B.n175 B.n174 163.367
R411 B.n484 B.n80 163.367
R412 B.n359 B.n232 163.367
R413 B.n359 B.n226 163.367
R414 B.n367 B.n226 163.367
R415 B.n367 B.n224 163.367
R416 B.n371 B.n224 163.367
R417 B.n371 B.n217 163.367
R418 B.n379 B.n217 163.367
R419 B.n379 B.n215 163.367
R420 B.n383 B.n215 163.367
R421 B.n383 B.n210 163.367
R422 B.n391 B.n210 163.367
R423 B.n391 B.n208 163.367
R424 B.n395 B.n208 163.367
R425 B.n395 B.n202 163.367
R426 B.n403 B.n202 163.367
R427 B.n403 B.n200 163.367
R428 B.n407 B.n200 163.367
R429 B.n407 B.n194 163.367
R430 B.n415 B.n194 163.367
R431 B.n415 B.n192 163.367
R432 B.n419 B.n192 163.367
R433 B.n419 B.n187 163.367
R434 B.n428 B.n187 163.367
R435 B.n428 B.n185 163.367
R436 B.n433 B.n185 163.367
R437 B.n433 B.n179 163.367
R438 B.n441 B.n179 163.367
R439 B.n442 B.n441 163.367
R440 B.n442 B.n5 163.367
R441 B.n6 B.n5 163.367
R442 B.n7 B.n6 163.367
R443 B.n448 B.n7 163.367
R444 B.n449 B.n448 163.367
R445 B.n449 B.n13 163.367
R446 B.n14 B.n13 163.367
R447 B.n15 B.n14 163.367
R448 B.n454 B.n15 163.367
R449 B.n454 B.n20 163.367
R450 B.n21 B.n20 163.367
R451 B.n22 B.n21 163.367
R452 B.n459 B.n22 163.367
R453 B.n459 B.n27 163.367
R454 B.n28 B.n27 163.367
R455 B.n29 B.n28 163.367
R456 B.n464 B.n29 163.367
R457 B.n464 B.n34 163.367
R458 B.n35 B.n34 163.367
R459 B.n36 B.n35 163.367
R460 B.n469 B.n36 163.367
R461 B.n469 B.n41 163.367
R462 B.n42 B.n41 163.367
R463 B.n43 B.n42 163.367
R464 B.n474 B.n43 163.367
R465 B.n474 B.n48 163.367
R466 B.n49 B.n48 163.367
R467 B.n50 B.n49 163.367
R468 B.n479 B.n50 163.367
R469 B.n479 B.n55 163.367
R470 B.n56 B.n55 163.367
R471 B.n257 B.n256 163.367
R472 B.n346 B.n256 163.367
R473 B.n344 B.n343 163.367
R474 B.n340 B.n339 163.367
R475 B.n336 B.n335 163.367
R476 B.n332 B.n331 163.367
R477 B.n328 B.n327 163.367
R478 B.n324 B.n323 163.367
R479 B.n320 B.n319 163.367
R480 B.n316 B.n315 163.367
R481 B.n312 B.n311 163.367
R482 B.n308 B.n307 163.367
R483 B.n304 B.n303 163.367
R484 B.n300 B.n299 163.367
R485 B.n295 B.n294 163.367
R486 B.n291 B.n290 163.367
R487 B.n287 B.n286 163.367
R488 B.n283 B.n282 163.367
R489 B.n279 B.n278 163.367
R490 B.n275 B.n274 163.367
R491 B.n271 B.n270 163.367
R492 B.n267 B.n266 163.367
R493 B.n263 B.n234 163.367
R494 B.n361 B.n230 163.367
R495 B.n361 B.n228 163.367
R496 B.n365 B.n228 163.367
R497 B.n365 B.n222 163.367
R498 B.n373 B.n222 163.367
R499 B.n373 B.n220 163.367
R500 B.n377 B.n220 163.367
R501 B.n377 B.n214 163.367
R502 B.n385 B.n214 163.367
R503 B.n385 B.n212 163.367
R504 B.n389 B.n212 163.367
R505 B.n389 B.n206 163.367
R506 B.n397 B.n206 163.367
R507 B.n397 B.n204 163.367
R508 B.n401 B.n204 163.367
R509 B.n401 B.n198 163.367
R510 B.n409 B.n198 163.367
R511 B.n409 B.n196 163.367
R512 B.n413 B.n196 163.367
R513 B.n413 B.n190 163.367
R514 B.n422 B.n190 163.367
R515 B.n422 B.n188 163.367
R516 B.n426 B.n188 163.367
R517 B.n426 B.n183 163.367
R518 B.n435 B.n183 163.367
R519 B.n435 B.n181 163.367
R520 B.n439 B.n181 163.367
R521 B.n439 B.n3 163.367
R522 B.n545 B.n3 163.367
R523 B.n541 B.n2 163.367
R524 B.n541 B.n540 163.367
R525 B.n540 B.n9 163.367
R526 B.n536 B.n9 163.367
R527 B.n536 B.n11 163.367
R528 B.n532 B.n11 163.367
R529 B.n532 B.n16 163.367
R530 B.n528 B.n16 163.367
R531 B.n528 B.n18 163.367
R532 B.n524 B.n18 163.367
R533 B.n524 B.n24 163.367
R534 B.n520 B.n24 163.367
R535 B.n520 B.n26 163.367
R536 B.n516 B.n26 163.367
R537 B.n516 B.n31 163.367
R538 B.n512 B.n31 163.367
R539 B.n512 B.n33 163.367
R540 B.n508 B.n33 163.367
R541 B.n508 B.n38 163.367
R542 B.n504 B.n38 163.367
R543 B.n504 B.n40 163.367
R544 B.n500 B.n40 163.367
R545 B.n500 B.n45 163.367
R546 B.n496 B.n45 163.367
R547 B.n496 B.n47 163.367
R548 B.n492 B.n47 163.367
R549 B.n492 B.n52 163.367
R550 B.n488 B.n52 163.367
R551 B.n488 B.n54 163.367
R552 B.n353 B.n231 159.219
R553 B.n486 B.n485 159.219
R554 B.n81 B.t4 144.45
R555 B.n261 B.t9 144.45
R556 B.n84 B.t11 144.446
R557 B.n258 B.t15 144.446
R558 B.n360 B.n231 79.0285
R559 B.n360 B.n227 79.0285
R560 B.n366 B.n227 79.0285
R561 B.n366 B.n223 79.0285
R562 B.n372 B.n223 79.0285
R563 B.n372 B.n218 79.0285
R564 B.n378 B.n218 79.0285
R565 B.n378 B.n219 79.0285
R566 B.n384 B.n211 79.0285
R567 B.n390 B.n211 79.0285
R568 B.n390 B.n207 79.0285
R569 B.n396 B.n207 79.0285
R570 B.n396 B.n203 79.0285
R571 B.n402 B.n203 79.0285
R572 B.n402 B.n199 79.0285
R573 B.n408 B.n199 79.0285
R574 B.n408 B.n195 79.0285
R575 B.n414 B.n195 79.0285
R576 B.n414 B.n191 79.0285
R577 B.n421 B.n191 79.0285
R578 B.n421 B.n420 79.0285
R579 B.n427 B.n184 79.0285
R580 B.n434 B.n184 79.0285
R581 B.n434 B.n180 79.0285
R582 B.n440 B.n180 79.0285
R583 B.n440 B.n4 79.0285
R584 B.n544 B.n4 79.0285
R585 B.n544 B.n543 79.0285
R586 B.n543 B.n542 79.0285
R587 B.n542 B.n8 79.0285
R588 B.n12 B.n8 79.0285
R589 B.n535 B.n12 79.0285
R590 B.n535 B.n534 79.0285
R591 B.n534 B.n533 79.0285
R592 B.n527 B.n19 79.0285
R593 B.n527 B.n526 79.0285
R594 B.n526 B.n525 79.0285
R595 B.n525 B.n23 79.0285
R596 B.n519 B.n23 79.0285
R597 B.n519 B.n518 79.0285
R598 B.n518 B.n517 79.0285
R599 B.n517 B.n30 79.0285
R600 B.n511 B.n30 79.0285
R601 B.n511 B.n510 79.0285
R602 B.n510 B.n509 79.0285
R603 B.n509 B.n37 79.0285
R604 B.n503 B.n37 79.0285
R605 B.n502 B.n501 79.0285
R606 B.n501 B.n44 79.0285
R607 B.n495 B.n44 79.0285
R608 B.n495 B.n494 79.0285
R609 B.n494 B.n493 79.0285
R610 B.n493 B.n51 79.0285
R611 B.n487 B.n51 79.0285
R612 B.n487 B.n486 79.0285
R613 B.n82 B.t5 73.2734
R614 B.n262 B.t8 73.2734
R615 B.n85 B.t12 73.2695
R616 B.n259 B.t14 73.2695
R617 B.n86 B.n57 71.676
R618 B.n90 B.n58 71.676
R619 B.n94 B.n59 71.676
R620 B.n98 B.n60 71.676
R621 B.n102 B.n61 71.676
R622 B.n106 B.n62 71.676
R623 B.n110 B.n63 71.676
R624 B.n114 B.n64 71.676
R625 B.n118 B.n65 71.676
R626 B.n122 B.n66 71.676
R627 B.n127 B.n67 71.676
R628 B.n131 B.n68 71.676
R629 B.n135 B.n69 71.676
R630 B.n139 B.n70 71.676
R631 B.n143 B.n71 71.676
R632 B.n147 B.n72 71.676
R633 B.n151 B.n73 71.676
R634 B.n155 B.n74 71.676
R635 B.n159 B.n75 71.676
R636 B.n163 B.n76 71.676
R637 B.n167 B.n77 71.676
R638 B.n171 B.n78 71.676
R639 B.n175 B.n79 71.676
R640 B.n80 B.n79 71.676
R641 B.n174 B.n78 71.676
R642 B.n170 B.n77 71.676
R643 B.n166 B.n76 71.676
R644 B.n162 B.n75 71.676
R645 B.n158 B.n74 71.676
R646 B.n154 B.n73 71.676
R647 B.n150 B.n72 71.676
R648 B.n146 B.n71 71.676
R649 B.n142 B.n70 71.676
R650 B.n138 B.n69 71.676
R651 B.n134 B.n68 71.676
R652 B.n130 B.n67 71.676
R653 B.n126 B.n66 71.676
R654 B.n121 B.n65 71.676
R655 B.n117 B.n64 71.676
R656 B.n113 B.n63 71.676
R657 B.n109 B.n62 71.676
R658 B.n105 B.n61 71.676
R659 B.n101 B.n60 71.676
R660 B.n97 B.n59 71.676
R661 B.n93 B.n58 71.676
R662 B.n89 B.n57 71.676
R663 B.n352 B.n351 71.676
R664 B.n346 B.n235 71.676
R665 B.n343 B.n236 71.676
R666 B.n339 B.n237 71.676
R667 B.n335 B.n238 71.676
R668 B.n331 B.n239 71.676
R669 B.n327 B.n240 71.676
R670 B.n323 B.n241 71.676
R671 B.n319 B.n242 71.676
R672 B.n315 B.n243 71.676
R673 B.n311 B.n244 71.676
R674 B.n307 B.n245 71.676
R675 B.n303 B.n246 71.676
R676 B.n299 B.n247 71.676
R677 B.n294 B.n248 71.676
R678 B.n290 B.n249 71.676
R679 B.n286 B.n250 71.676
R680 B.n282 B.n251 71.676
R681 B.n278 B.n252 71.676
R682 B.n274 B.n253 71.676
R683 B.n270 B.n254 71.676
R684 B.n266 B.n255 71.676
R685 B.n354 B.n234 71.676
R686 B.n352 B.n257 71.676
R687 B.n344 B.n235 71.676
R688 B.n340 B.n236 71.676
R689 B.n336 B.n237 71.676
R690 B.n332 B.n238 71.676
R691 B.n328 B.n239 71.676
R692 B.n324 B.n240 71.676
R693 B.n320 B.n241 71.676
R694 B.n316 B.n242 71.676
R695 B.n312 B.n243 71.676
R696 B.n308 B.n244 71.676
R697 B.n304 B.n245 71.676
R698 B.n300 B.n246 71.676
R699 B.n295 B.n247 71.676
R700 B.n291 B.n248 71.676
R701 B.n287 B.n249 71.676
R702 B.n283 B.n250 71.676
R703 B.n279 B.n251 71.676
R704 B.n275 B.n252 71.676
R705 B.n271 B.n253 71.676
R706 B.n267 B.n254 71.676
R707 B.n263 B.n255 71.676
R708 B.n355 B.n354 71.676
R709 B.n546 B.n545 71.676
R710 B.n546 B.n2 71.676
R711 B.n85 B.n84 71.1763
R712 B.n82 B.n81 71.1763
R713 B.n262 B.n261 71.1763
R714 B.n259 B.n258 71.1763
R715 B.n124 B.n85 59.5399
R716 B.n83 B.n82 59.5399
R717 B.n297 B.n262 59.5399
R718 B.n260 B.n259 59.5399
R719 B.n219 B.t7 39.5145
R720 B.n384 B.t7 39.5145
R721 B.n420 B.t0 39.5145
R722 B.n427 B.t0 39.5145
R723 B.n533 B.t1 39.5145
R724 B.n19 B.t1 39.5145
R725 B.n503 B.t3 39.5145
R726 B.t3 B.n502 39.5145
R727 B.n350 B.n229 33.8737
R728 B.n357 B.n356 33.8737
R729 B.n483 B.n482 33.8737
R730 B.n87 B.n53 33.8737
R731 B B.n547 18.0485
R732 B.n362 B.n229 10.6151
R733 B.n363 B.n362 10.6151
R734 B.n364 B.n363 10.6151
R735 B.n364 B.n221 10.6151
R736 B.n374 B.n221 10.6151
R737 B.n375 B.n374 10.6151
R738 B.n376 B.n375 10.6151
R739 B.n376 B.n213 10.6151
R740 B.n386 B.n213 10.6151
R741 B.n387 B.n386 10.6151
R742 B.n388 B.n387 10.6151
R743 B.n388 B.n205 10.6151
R744 B.n398 B.n205 10.6151
R745 B.n399 B.n398 10.6151
R746 B.n400 B.n399 10.6151
R747 B.n400 B.n197 10.6151
R748 B.n410 B.n197 10.6151
R749 B.n411 B.n410 10.6151
R750 B.n412 B.n411 10.6151
R751 B.n412 B.n189 10.6151
R752 B.n423 B.n189 10.6151
R753 B.n424 B.n423 10.6151
R754 B.n425 B.n424 10.6151
R755 B.n425 B.n182 10.6151
R756 B.n436 B.n182 10.6151
R757 B.n437 B.n436 10.6151
R758 B.n438 B.n437 10.6151
R759 B.n438 B.n0 10.6151
R760 B.n350 B.n349 10.6151
R761 B.n349 B.n348 10.6151
R762 B.n348 B.n347 10.6151
R763 B.n347 B.n345 10.6151
R764 B.n345 B.n342 10.6151
R765 B.n342 B.n341 10.6151
R766 B.n341 B.n338 10.6151
R767 B.n338 B.n337 10.6151
R768 B.n337 B.n334 10.6151
R769 B.n334 B.n333 10.6151
R770 B.n333 B.n330 10.6151
R771 B.n330 B.n329 10.6151
R772 B.n329 B.n326 10.6151
R773 B.n326 B.n325 10.6151
R774 B.n325 B.n322 10.6151
R775 B.n322 B.n321 10.6151
R776 B.n321 B.n318 10.6151
R777 B.n318 B.n317 10.6151
R778 B.n314 B.n313 10.6151
R779 B.n313 B.n310 10.6151
R780 B.n310 B.n309 10.6151
R781 B.n309 B.n306 10.6151
R782 B.n306 B.n305 10.6151
R783 B.n305 B.n302 10.6151
R784 B.n302 B.n301 10.6151
R785 B.n301 B.n298 10.6151
R786 B.n296 B.n293 10.6151
R787 B.n293 B.n292 10.6151
R788 B.n292 B.n289 10.6151
R789 B.n289 B.n288 10.6151
R790 B.n288 B.n285 10.6151
R791 B.n285 B.n284 10.6151
R792 B.n284 B.n281 10.6151
R793 B.n281 B.n280 10.6151
R794 B.n280 B.n277 10.6151
R795 B.n277 B.n276 10.6151
R796 B.n276 B.n273 10.6151
R797 B.n273 B.n272 10.6151
R798 B.n272 B.n269 10.6151
R799 B.n269 B.n268 10.6151
R800 B.n268 B.n265 10.6151
R801 B.n265 B.n264 10.6151
R802 B.n264 B.n233 10.6151
R803 B.n356 B.n233 10.6151
R804 B.n358 B.n357 10.6151
R805 B.n358 B.n225 10.6151
R806 B.n368 B.n225 10.6151
R807 B.n369 B.n368 10.6151
R808 B.n370 B.n369 10.6151
R809 B.n370 B.n216 10.6151
R810 B.n380 B.n216 10.6151
R811 B.n381 B.n380 10.6151
R812 B.n382 B.n381 10.6151
R813 B.n382 B.n209 10.6151
R814 B.n392 B.n209 10.6151
R815 B.n393 B.n392 10.6151
R816 B.n394 B.n393 10.6151
R817 B.n394 B.n201 10.6151
R818 B.n404 B.n201 10.6151
R819 B.n405 B.n404 10.6151
R820 B.n406 B.n405 10.6151
R821 B.n406 B.n193 10.6151
R822 B.n416 B.n193 10.6151
R823 B.n417 B.n416 10.6151
R824 B.n418 B.n417 10.6151
R825 B.n418 B.n186 10.6151
R826 B.n429 B.n186 10.6151
R827 B.n430 B.n429 10.6151
R828 B.n432 B.n430 10.6151
R829 B.n432 B.n431 10.6151
R830 B.n431 B.n178 10.6151
R831 B.n443 B.n178 10.6151
R832 B.n444 B.n443 10.6151
R833 B.n445 B.n444 10.6151
R834 B.n446 B.n445 10.6151
R835 B.n447 B.n446 10.6151
R836 B.n450 B.n447 10.6151
R837 B.n451 B.n450 10.6151
R838 B.n452 B.n451 10.6151
R839 B.n453 B.n452 10.6151
R840 B.n455 B.n453 10.6151
R841 B.n456 B.n455 10.6151
R842 B.n457 B.n456 10.6151
R843 B.n458 B.n457 10.6151
R844 B.n460 B.n458 10.6151
R845 B.n461 B.n460 10.6151
R846 B.n462 B.n461 10.6151
R847 B.n463 B.n462 10.6151
R848 B.n465 B.n463 10.6151
R849 B.n466 B.n465 10.6151
R850 B.n467 B.n466 10.6151
R851 B.n468 B.n467 10.6151
R852 B.n470 B.n468 10.6151
R853 B.n471 B.n470 10.6151
R854 B.n472 B.n471 10.6151
R855 B.n473 B.n472 10.6151
R856 B.n475 B.n473 10.6151
R857 B.n476 B.n475 10.6151
R858 B.n477 B.n476 10.6151
R859 B.n478 B.n477 10.6151
R860 B.n480 B.n478 10.6151
R861 B.n481 B.n480 10.6151
R862 B.n482 B.n481 10.6151
R863 B.n539 B.n1 10.6151
R864 B.n539 B.n538 10.6151
R865 B.n538 B.n537 10.6151
R866 B.n537 B.n10 10.6151
R867 B.n531 B.n10 10.6151
R868 B.n531 B.n530 10.6151
R869 B.n530 B.n529 10.6151
R870 B.n529 B.n17 10.6151
R871 B.n523 B.n17 10.6151
R872 B.n523 B.n522 10.6151
R873 B.n522 B.n521 10.6151
R874 B.n521 B.n25 10.6151
R875 B.n515 B.n25 10.6151
R876 B.n515 B.n514 10.6151
R877 B.n514 B.n513 10.6151
R878 B.n513 B.n32 10.6151
R879 B.n507 B.n32 10.6151
R880 B.n507 B.n506 10.6151
R881 B.n506 B.n505 10.6151
R882 B.n505 B.n39 10.6151
R883 B.n499 B.n39 10.6151
R884 B.n499 B.n498 10.6151
R885 B.n498 B.n497 10.6151
R886 B.n497 B.n46 10.6151
R887 B.n491 B.n46 10.6151
R888 B.n491 B.n490 10.6151
R889 B.n490 B.n489 10.6151
R890 B.n489 B.n53 10.6151
R891 B.n88 B.n87 10.6151
R892 B.n91 B.n88 10.6151
R893 B.n92 B.n91 10.6151
R894 B.n95 B.n92 10.6151
R895 B.n96 B.n95 10.6151
R896 B.n99 B.n96 10.6151
R897 B.n100 B.n99 10.6151
R898 B.n103 B.n100 10.6151
R899 B.n104 B.n103 10.6151
R900 B.n107 B.n104 10.6151
R901 B.n108 B.n107 10.6151
R902 B.n111 B.n108 10.6151
R903 B.n112 B.n111 10.6151
R904 B.n115 B.n112 10.6151
R905 B.n116 B.n115 10.6151
R906 B.n119 B.n116 10.6151
R907 B.n120 B.n119 10.6151
R908 B.n123 B.n120 10.6151
R909 B.n128 B.n125 10.6151
R910 B.n129 B.n128 10.6151
R911 B.n132 B.n129 10.6151
R912 B.n133 B.n132 10.6151
R913 B.n136 B.n133 10.6151
R914 B.n137 B.n136 10.6151
R915 B.n140 B.n137 10.6151
R916 B.n141 B.n140 10.6151
R917 B.n145 B.n144 10.6151
R918 B.n148 B.n145 10.6151
R919 B.n149 B.n148 10.6151
R920 B.n152 B.n149 10.6151
R921 B.n153 B.n152 10.6151
R922 B.n156 B.n153 10.6151
R923 B.n157 B.n156 10.6151
R924 B.n160 B.n157 10.6151
R925 B.n161 B.n160 10.6151
R926 B.n164 B.n161 10.6151
R927 B.n165 B.n164 10.6151
R928 B.n168 B.n165 10.6151
R929 B.n169 B.n168 10.6151
R930 B.n172 B.n169 10.6151
R931 B.n173 B.n172 10.6151
R932 B.n176 B.n173 10.6151
R933 B.n177 B.n176 10.6151
R934 B.n483 B.n177 10.6151
R935 B.n547 B.n0 8.11757
R936 B.n547 B.n1 8.11757
R937 B.n314 B.n260 6.5566
R938 B.n298 B.n297 6.5566
R939 B.n125 B.n124 6.5566
R940 B.n141 B.n83 6.5566
R941 B.n317 B.n260 4.05904
R942 B.n297 B.n296 4.05904
R943 B.n124 B.n123 4.05904
R944 B.n144 B.n83 4.05904
R945 VP.n0 VP.t1 109.724
R946 VP.n0 VP.t0 69.0215
R947 VP VP.n0 0.52637
R948 VTAIL.n1 VTAIL.t0 59.7712
R949 VTAIL.n2 VTAIL.t2 59.771
R950 VTAIL.n3 VTAIL.t1 59.771
R951 VTAIL.n0 VTAIL.t3 59.771
R952 VTAIL.n1 VTAIL.n0 22.3065
R953 VTAIL.n3 VTAIL.n2 19.1427
R954 VTAIL.n2 VTAIL.n1 2.05222
R955 VTAIL VTAIL.n0 1.31947
R956 VTAIL VTAIL.n3 0.733259
R957 VDD1 VDD1.t1 111.365
R958 VDD1 VDD1.t0 77.299
R959 VN VN.t0 109.63
R960 VN VN.t1 69.5473
R961 VDD2.n0 VDD2.t0 110.049
R962 VDD2.n0 VDD2.t1 76.4498
R963 VDD2 VDD2.n0 0.849638
C0 VN VP 4.36341f
C1 VTAIL VDD1 3.22247f
C2 VDD2 VP 0.368164f
C3 VDD1 VN 0.152597f
C4 VTAIL VN 1.38195f
C5 VDD2 VDD1 0.764169f
C6 VDD2 VTAIL 3.28011f
C7 VDD2 VN 1.17372f
C8 VDD1 VP 1.38774f
C9 VTAIL VP 1.39611f
C10 VDD2 B 3.242504f
C11 VDD1 B 5.23695f
C12 VTAIL B 4.209258f
C13 VN B 8.625521f
C14 VP B 6.604544f
C15 VDD2.t0 B 0.803443f
C16 VDD2.t1 B 0.537155f
C17 VDD2.n0 B 1.8326f
C18 VN.t1 B 1.00835f
C19 VN.t0 B 1.44063f
C20 VDD1.t0 B 0.513821f
C21 VDD1.t1 B 0.789089f
C22 VTAIL.t3 B 0.560127f
C23 VTAIL.n0 B 1.11492f
C24 VTAIL.t0 B 0.560129f
C25 VTAIL.n1 B 1.1581f
C26 VTAIL.t2 B 0.560127f
C27 VTAIL.n2 B 0.971645f
C28 VTAIL.t1 B 0.560127f
C29 VTAIL.n3 B 0.893912f
C30 VP.t1 B 1.4496f
C31 VP.t0 B 1.01253f
C32 VP.n0 B 1.86346f
.ends

