* NGSPICE file created from diff_pair_sample_1175.ext - technology: sky130A

.subckt diff_pair_sample_1175 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=2.51295 ps=15.56 w=15.23 l=0.69
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=0 ps=0 w=15.23 l=0.69
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=0 ps=0 w=15.23 l=0.69
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=0 ps=0 w=15.23 l=0.69
X4 VDD2.t3 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.51295 pd=15.56 as=5.9397 ps=31.24 w=15.23 l=0.69
X5 VTAIL.t0 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=2.51295 ps=15.56 w=15.23 l=0.69
X6 VDD2.t2 VN.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.51295 pd=15.56 as=5.9397 ps=31.24 w=15.23 l=0.69
X7 VTAIL.t4 VN.t3 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=2.51295 ps=15.56 w=15.23 l=0.69
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=0 ps=0 w=15.23 l=0.69
X9 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=5.9397 pd=31.24 as=2.51295 ps=15.56 w=15.23 l=0.69
X10 VDD1.t1 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.51295 pd=15.56 as=5.9397 ps=31.24 w=15.23 l=0.69
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.51295 pd=15.56 as=5.9397 ps=31.24 w=15.23 l=0.69
R0 VN.n0 VN.t0 610.225
R1 VN.n1 VN.t2 610.225
R2 VN.n0 VN.t1 610.174
R3 VN.n1 VN.t3 610.174
R4 VN VN.n1 87.861
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 104.823
R7 VDD2.n2 VDD2.n1 65.3402
R8 VDD2.n1 VDD2.t1 1.30057
R9 VDD2.n1 VDD2.t2 1.30057
R10 VDD2.n0 VDD2.t0 1.30057
R11 VDD2.n0 VDD2.t3 1.30057
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t3 49.9617
R14 VTAIL.n4 VTAIL.t5 49.9617
R15 VTAIL.n3 VTAIL.t4 49.9617
R16 VTAIL.n7 VTAIL.t6 49.9614
R17 VTAIL.n0 VTAIL.t7 49.9614
R18 VTAIL.n1 VTAIL.t2 49.9614
R19 VTAIL.n2 VTAIL.t0 49.9614
R20 VTAIL.n6 VTAIL.t1 49.9614
R21 VTAIL.n7 VTAIL.n6 26.3755
R22 VTAIL.n3 VTAIL.n2 26.3755
R23 VTAIL.n4 VTAIL.n3 0.87981
R24 VTAIL.n6 VTAIL.n5 0.87981
R25 VTAIL.n2 VTAIL.n1 0.87981
R26 VTAIL VTAIL.n0 0.498345
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.381966
R30 B.n410 B.t15 735.037
R31 B.n407 B.t8 735.037
R32 B.n93 B.t4 735.037
R33 B.n91 B.t12 735.037
R34 B.n709 B.n708 585
R35 B.n317 B.n90 585
R36 B.n316 B.n315 585
R37 B.n314 B.n313 585
R38 B.n312 B.n311 585
R39 B.n310 B.n309 585
R40 B.n308 B.n307 585
R41 B.n306 B.n305 585
R42 B.n304 B.n303 585
R43 B.n302 B.n301 585
R44 B.n300 B.n299 585
R45 B.n298 B.n297 585
R46 B.n296 B.n295 585
R47 B.n294 B.n293 585
R48 B.n292 B.n291 585
R49 B.n290 B.n289 585
R50 B.n288 B.n287 585
R51 B.n286 B.n285 585
R52 B.n284 B.n283 585
R53 B.n282 B.n281 585
R54 B.n280 B.n279 585
R55 B.n278 B.n277 585
R56 B.n276 B.n275 585
R57 B.n274 B.n273 585
R58 B.n272 B.n271 585
R59 B.n270 B.n269 585
R60 B.n268 B.n267 585
R61 B.n266 B.n265 585
R62 B.n264 B.n263 585
R63 B.n262 B.n261 585
R64 B.n260 B.n259 585
R65 B.n258 B.n257 585
R66 B.n256 B.n255 585
R67 B.n254 B.n253 585
R68 B.n252 B.n251 585
R69 B.n250 B.n249 585
R70 B.n248 B.n247 585
R71 B.n246 B.n245 585
R72 B.n244 B.n243 585
R73 B.n242 B.n241 585
R74 B.n240 B.n239 585
R75 B.n238 B.n237 585
R76 B.n236 B.n235 585
R77 B.n234 B.n233 585
R78 B.n232 B.n231 585
R79 B.n230 B.n229 585
R80 B.n228 B.n227 585
R81 B.n226 B.n225 585
R82 B.n224 B.n223 585
R83 B.n222 B.n221 585
R84 B.n220 B.n219 585
R85 B.n217 B.n216 585
R86 B.n215 B.n214 585
R87 B.n213 B.n212 585
R88 B.n211 B.n210 585
R89 B.n209 B.n208 585
R90 B.n207 B.n206 585
R91 B.n205 B.n204 585
R92 B.n203 B.n202 585
R93 B.n201 B.n200 585
R94 B.n199 B.n198 585
R95 B.n196 B.n195 585
R96 B.n194 B.n193 585
R97 B.n192 B.n191 585
R98 B.n190 B.n189 585
R99 B.n188 B.n187 585
R100 B.n186 B.n185 585
R101 B.n184 B.n183 585
R102 B.n182 B.n181 585
R103 B.n180 B.n179 585
R104 B.n178 B.n177 585
R105 B.n176 B.n175 585
R106 B.n174 B.n173 585
R107 B.n172 B.n171 585
R108 B.n170 B.n169 585
R109 B.n168 B.n167 585
R110 B.n166 B.n165 585
R111 B.n164 B.n163 585
R112 B.n162 B.n161 585
R113 B.n160 B.n159 585
R114 B.n158 B.n157 585
R115 B.n156 B.n155 585
R116 B.n154 B.n153 585
R117 B.n152 B.n151 585
R118 B.n150 B.n149 585
R119 B.n148 B.n147 585
R120 B.n146 B.n145 585
R121 B.n144 B.n143 585
R122 B.n142 B.n141 585
R123 B.n140 B.n139 585
R124 B.n138 B.n137 585
R125 B.n136 B.n135 585
R126 B.n134 B.n133 585
R127 B.n132 B.n131 585
R128 B.n130 B.n129 585
R129 B.n128 B.n127 585
R130 B.n126 B.n125 585
R131 B.n124 B.n123 585
R132 B.n122 B.n121 585
R133 B.n120 B.n119 585
R134 B.n118 B.n117 585
R135 B.n116 B.n115 585
R136 B.n114 B.n113 585
R137 B.n112 B.n111 585
R138 B.n110 B.n109 585
R139 B.n108 B.n107 585
R140 B.n106 B.n105 585
R141 B.n104 B.n103 585
R142 B.n102 B.n101 585
R143 B.n100 B.n99 585
R144 B.n98 B.n97 585
R145 B.n96 B.n95 585
R146 B.n707 B.n34 585
R147 B.n712 B.n34 585
R148 B.n706 B.n33 585
R149 B.n713 B.n33 585
R150 B.n705 B.n704 585
R151 B.n704 B.n29 585
R152 B.n703 B.n28 585
R153 B.n719 B.n28 585
R154 B.n702 B.n27 585
R155 B.n720 B.n27 585
R156 B.n701 B.n26 585
R157 B.n721 B.n26 585
R158 B.n700 B.n699 585
R159 B.n699 B.n22 585
R160 B.n698 B.n21 585
R161 B.n727 B.n21 585
R162 B.n697 B.n20 585
R163 B.n728 B.n20 585
R164 B.n696 B.n19 585
R165 B.n729 B.n19 585
R166 B.n695 B.n694 585
R167 B.n694 B.n18 585
R168 B.n693 B.n14 585
R169 B.n735 B.n14 585
R170 B.n692 B.n13 585
R171 B.n736 B.n13 585
R172 B.n691 B.n12 585
R173 B.n737 B.n12 585
R174 B.n690 B.n689 585
R175 B.n689 B.n8 585
R176 B.n688 B.n7 585
R177 B.n743 B.n7 585
R178 B.n687 B.n6 585
R179 B.n744 B.n6 585
R180 B.n686 B.n5 585
R181 B.n745 B.n5 585
R182 B.n685 B.n684 585
R183 B.n684 B.n4 585
R184 B.n683 B.n318 585
R185 B.n683 B.n682 585
R186 B.n673 B.n319 585
R187 B.n320 B.n319 585
R188 B.n675 B.n674 585
R189 B.n676 B.n675 585
R190 B.n672 B.n325 585
R191 B.n325 B.n324 585
R192 B.n671 B.n670 585
R193 B.n670 B.n669 585
R194 B.n327 B.n326 585
R195 B.n662 B.n327 585
R196 B.n661 B.n660 585
R197 B.n663 B.n661 585
R198 B.n659 B.n332 585
R199 B.n332 B.n331 585
R200 B.n658 B.n657 585
R201 B.n657 B.n656 585
R202 B.n334 B.n333 585
R203 B.n335 B.n334 585
R204 B.n649 B.n648 585
R205 B.n650 B.n649 585
R206 B.n647 B.n339 585
R207 B.n343 B.n339 585
R208 B.n646 B.n645 585
R209 B.n645 B.n644 585
R210 B.n341 B.n340 585
R211 B.n342 B.n341 585
R212 B.n637 B.n636 585
R213 B.n638 B.n637 585
R214 B.n635 B.n348 585
R215 B.n348 B.n347 585
R216 B.n630 B.n629 585
R217 B.n628 B.n406 585
R218 B.n627 B.n405 585
R219 B.n632 B.n405 585
R220 B.n626 B.n625 585
R221 B.n624 B.n623 585
R222 B.n622 B.n621 585
R223 B.n620 B.n619 585
R224 B.n618 B.n617 585
R225 B.n616 B.n615 585
R226 B.n614 B.n613 585
R227 B.n612 B.n611 585
R228 B.n610 B.n609 585
R229 B.n608 B.n607 585
R230 B.n606 B.n605 585
R231 B.n604 B.n603 585
R232 B.n602 B.n601 585
R233 B.n600 B.n599 585
R234 B.n598 B.n597 585
R235 B.n596 B.n595 585
R236 B.n594 B.n593 585
R237 B.n592 B.n591 585
R238 B.n590 B.n589 585
R239 B.n588 B.n587 585
R240 B.n586 B.n585 585
R241 B.n584 B.n583 585
R242 B.n582 B.n581 585
R243 B.n580 B.n579 585
R244 B.n578 B.n577 585
R245 B.n576 B.n575 585
R246 B.n574 B.n573 585
R247 B.n572 B.n571 585
R248 B.n570 B.n569 585
R249 B.n568 B.n567 585
R250 B.n566 B.n565 585
R251 B.n564 B.n563 585
R252 B.n562 B.n561 585
R253 B.n560 B.n559 585
R254 B.n558 B.n557 585
R255 B.n556 B.n555 585
R256 B.n554 B.n553 585
R257 B.n552 B.n551 585
R258 B.n550 B.n549 585
R259 B.n548 B.n547 585
R260 B.n546 B.n545 585
R261 B.n544 B.n543 585
R262 B.n542 B.n541 585
R263 B.n540 B.n539 585
R264 B.n538 B.n537 585
R265 B.n536 B.n535 585
R266 B.n534 B.n533 585
R267 B.n532 B.n531 585
R268 B.n530 B.n529 585
R269 B.n528 B.n527 585
R270 B.n526 B.n525 585
R271 B.n524 B.n523 585
R272 B.n522 B.n521 585
R273 B.n520 B.n519 585
R274 B.n518 B.n517 585
R275 B.n516 B.n515 585
R276 B.n514 B.n513 585
R277 B.n512 B.n511 585
R278 B.n510 B.n509 585
R279 B.n508 B.n507 585
R280 B.n506 B.n505 585
R281 B.n504 B.n503 585
R282 B.n502 B.n501 585
R283 B.n500 B.n499 585
R284 B.n498 B.n497 585
R285 B.n496 B.n495 585
R286 B.n494 B.n493 585
R287 B.n492 B.n491 585
R288 B.n490 B.n489 585
R289 B.n488 B.n487 585
R290 B.n486 B.n485 585
R291 B.n484 B.n483 585
R292 B.n482 B.n481 585
R293 B.n480 B.n479 585
R294 B.n478 B.n477 585
R295 B.n476 B.n475 585
R296 B.n474 B.n473 585
R297 B.n472 B.n471 585
R298 B.n470 B.n469 585
R299 B.n468 B.n467 585
R300 B.n466 B.n465 585
R301 B.n464 B.n463 585
R302 B.n462 B.n461 585
R303 B.n460 B.n459 585
R304 B.n458 B.n457 585
R305 B.n456 B.n455 585
R306 B.n454 B.n453 585
R307 B.n452 B.n451 585
R308 B.n450 B.n449 585
R309 B.n448 B.n447 585
R310 B.n446 B.n445 585
R311 B.n444 B.n443 585
R312 B.n442 B.n441 585
R313 B.n440 B.n439 585
R314 B.n438 B.n437 585
R315 B.n436 B.n435 585
R316 B.n434 B.n433 585
R317 B.n432 B.n431 585
R318 B.n430 B.n429 585
R319 B.n428 B.n427 585
R320 B.n426 B.n425 585
R321 B.n424 B.n423 585
R322 B.n422 B.n421 585
R323 B.n420 B.n419 585
R324 B.n418 B.n417 585
R325 B.n416 B.n415 585
R326 B.n414 B.n413 585
R327 B.n350 B.n349 585
R328 B.n634 B.n633 585
R329 B.n633 B.n632 585
R330 B.n346 B.n345 585
R331 B.n347 B.n346 585
R332 B.n640 B.n639 585
R333 B.n639 B.n638 585
R334 B.n641 B.n344 585
R335 B.n344 B.n342 585
R336 B.n643 B.n642 585
R337 B.n644 B.n643 585
R338 B.n338 B.n337 585
R339 B.n343 B.n338 585
R340 B.n652 B.n651 585
R341 B.n651 B.n650 585
R342 B.n653 B.n336 585
R343 B.n336 B.n335 585
R344 B.n655 B.n654 585
R345 B.n656 B.n655 585
R346 B.n330 B.n329 585
R347 B.n331 B.n330 585
R348 B.n665 B.n664 585
R349 B.n664 B.n663 585
R350 B.n666 B.n328 585
R351 B.n662 B.n328 585
R352 B.n668 B.n667 585
R353 B.n669 B.n668 585
R354 B.n323 B.n322 585
R355 B.n324 B.n323 585
R356 B.n678 B.n677 585
R357 B.n677 B.n676 585
R358 B.n679 B.n321 585
R359 B.n321 B.n320 585
R360 B.n681 B.n680 585
R361 B.n682 B.n681 585
R362 B.n2 B.n0 585
R363 B.n4 B.n2 585
R364 B.n3 B.n1 585
R365 B.n744 B.n3 585
R366 B.n742 B.n741 585
R367 B.n743 B.n742 585
R368 B.n740 B.n9 585
R369 B.n9 B.n8 585
R370 B.n739 B.n738 585
R371 B.n738 B.n737 585
R372 B.n11 B.n10 585
R373 B.n736 B.n11 585
R374 B.n734 B.n733 585
R375 B.n735 B.n734 585
R376 B.n732 B.n15 585
R377 B.n18 B.n15 585
R378 B.n731 B.n730 585
R379 B.n730 B.n729 585
R380 B.n17 B.n16 585
R381 B.n728 B.n17 585
R382 B.n726 B.n725 585
R383 B.n727 B.n726 585
R384 B.n724 B.n23 585
R385 B.n23 B.n22 585
R386 B.n723 B.n722 585
R387 B.n722 B.n721 585
R388 B.n25 B.n24 585
R389 B.n720 B.n25 585
R390 B.n718 B.n717 585
R391 B.n719 B.n718 585
R392 B.n716 B.n30 585
R393 B.n30 B.n29 585
R394 B.n715 B.n714 585
R395 B.n714 B.n713 585
R396 B.n32 B.n31 585
R397 B.n712 B.n32 585
R398 B.n747 B.n746 585
R399 B.n746 B.n745 585
R400 B.n630 B.n346 502.111
R401 B.n95 B.n32 502.111
R402 B.n633 B.n348 502.111
R403 B.n709 B.n34 502.111
R404 B.n711 B.n710 256.663
R405 B.n711 B.n89 256.663
R406 B.n711 B.n88 256.663
R407 B.n711 B.n87 256.663
R408 B.n711 B.n86 256.663
R409 B.n711 B.n85 256.663
R410 B.n711 B.n84 256.663
R411 B.n711 B.n83 256.663
R412 B.n711 B.n82 256.663
R413 B.n711 B.n81 256.663
R414 B.n711 B.n80 256.663
R415 B.n711 B.n79 256.663
R416 B.n711 B.n78 256.663
R417 B.n711 B.n77 256.663
R418 B.n711 B.n76 256.663
R419 B.n711 B.n75 256.663
R420 B.n711 B.n74 256.663
R421 B.n711 B.n73 256.663
R422 B.n711 B.n72 256.663
R423 B.n711 B.n71 256.663
R424 B.n711 B.n70 256.663
R425 B.n711 B.n69 256.663
R426 B.n711 B.n68 256.663
R427 B.n711 B.n67 256.663
R428 B.n711 B.n66 256.663
R429 B.n711 B.n65 256.663
R430 B.n711 B.n64 256.663
R431 B.n711 B.n63 256.663
R432 B.n711 B.n62 256.663
R433 B.n711 B.n61 256.663
R434 B.n711 B.n60 256.663
R435 B.n711 B.n59 256.663
R436 B.n711 B.n58 256.663
R437 B.n711 B.n57 256.663
R438 B.n711 B.n56 256.663
R439 B.n711 B.n55 256.663
R440 B.n711 B.n54 256.663
R441 B.n711 B.n53 256.663
R442 B.n711 B.n52 256.663
R443 B.n711 B.n51 256.663
R444 B.n711 B.n50 256.663
R445 B.n711 B.n49 256.663
R446 B.n711 B.n48 256.663
R447 B.n711 B.n47 256.663
R448 B.n711 B.n46 256.663
R449 B.n711 B.n45 256.663
R450 B.n711 B.n44 256.663
R451 B.n711 B.n43 256.663
R452 B.n711 B.n42 256.663
R453 B.n711 B.n41 256.663
R454 B.n711 B.n40 256.663
R455 B.n711 B.n39 256.663
R456 B.n711 B.n38 256.663
R457 B.n711 B.n37 256.663
R458 B.n711 B.n36 256.663
R459 B.n711 B.n35 256.663
R460 B.n632 B.n631 256.663
R461 B.n632 B.n351 256.663
R462 B.n632 B.n352 256.663
R463 B.n632 B.n353 256.663
R464 B.n632 B.n354 256.663
R465 B.n632 B.n355 256.663
R466 B.n632 B.n356 256.663
R467 B.n632 B.n357 256.663
R468 B.n632 B.n358 256.663
R469 B.n632 B.n359 256.663
R470 B.n632 B.n360 256.663
R471 B.n632 B.n361 256.663
R472 B.n632 B.n362 256.663
R473 B.n632 B.n363 256.663
R474 B.n632 B.n364 256.663
R475 B.n632 B.n365 256.663
R476 B.n632 B.n366 256.663
R477 B.n632 B.n367 256.663
R478 B.n632 B.n368 256.663
R479 B.n632 B.n369 256.663
R480 B.n632 B.n370 256.663
R481 B.n632 B.n371 256.663
R482 B.n632 B.n372 256.663
R483 B.n632 B.n373 256.663
R484 B.n632 B.n374 256.663
R485 B.n632 B.n375 256.663
R486 B.n632 B.n376 256.663
R487 B.n632 B.n377 256.663
R488 B.n632 B.n378 256.663
R489 B.n632 B.n379 256.663
R490 B.n632 B.n380 256.663
R491 B.n632 B.n381 256.663
R492 B.n632 B.n382 256.663
R493 B.n632 B.n383 256.663
R494 B.n632 B.n384 256.663
R495 B.n632 B.n385 256.663
R496 B.n632 B.n386 256.663
R497 B.n632 B.n387 256.663
R498 B.n632 B.n388 256.663
R499 B.n632 B.n389 256.663
R500 B.n632 B.n390 256.663
R501 B.n632 B.n391 256.663
R502 B.n632 B.n392 256.663
R503 B.n632 B.n393 256.663
R504 B.n632 B.n394 256.663
R505 B.n632 B.n395 256.663
R506 B.n632 B.n396 256.663
R507 B.n632 B.n397 256.663
R508 B.n632 B.n398 256.663
R509 B.n632 B.n399 256.663
R510 B.n632 B.n400 256.663
R511 B.n632 B.n401 256.663
R512 B.n632 B.n402 256.663
R513 B.n632 B.n403 256.663
R514 B.n632 B.n404 256.663
R515 B.n639 B.n346 163.367
R516 B.n639 B.n344 163.367
R517 B.n643 B.n344 163.367
R518 B.n643 B.n338 163.367
R519 B.n651 B.n338 163.367
R520 B.n651 B.n336 163.367
R521 B.n655 B.n336 163.367
R522 B.n655 B.n330 163.367
R523 B.n664 B.n330 163.367
R524 B.n664 B.n328 163.367
R525 B.n668 B.n328 163.367
R526 B.n668 B.n323 163.367
R527 B.n677 B.n323 163.367
R528 B.n677 B.n321 163.367
R529 B.n681 B.n321 163.367
R530 B.n681 B.n2 163.367
R531 B.n746 B.n2 163.367
R532 B.n746 B.n3 163.367
R533 B.n742 B.n3 163.367
R534 B.n742 B.n9 163.367
R535 B.n738 B.n9 163.367
R536 B.n738 B.n11 163.367
R537 B.n734 B.n11 163.367
R538 B.n734 B.n15 163.367
R539 B.n730 B.n15 163.367
R540 B.n730 B.n17 163.367
R541 B.n726 B.n17 163.367
R542 B.n726 B.n23 163.367
R543 B.n722 B.n23 163.367
R544 B.n722 B.n25 163.367
R545 B.n718 B.n25 163.367
R546 B.n718 B.n30 163.367
R547 B.n714 B.n30 163.367
R548 B.n714 B.n32 163.367
R549 B.n406 B.n405 163.367
R550 B.n625 B.n405 163.367
R551 B.n623 B.n622 163.367
R552 B.n619 B.n618 163.367
R553 B.n615 B.n614 163.367
R554 B.n611 B.n610 163.367
R555 B.n607 B.n606 163.367
R556 B.n603 B.n602 163.367
R557 B.n599 B.n598 163.367
R558 B.n595 B.n594 163.367
R559 B.n591 B.n590 163.367
R560 B.n587 B.n586 163.367
R561 B.n583 B.n582 163.367
R562 B.n579 B.n578 163.367
R563 B.n575 B.n574 163.367
R564 B.n571 B.n570 163.367
R565 B.n567 B.n566 163.367
R566 B.n563 B.n562 163.367
R567 B.n559 B.n558 163.367
R568 B.n555 B.n554 163.367
R569 B.n551 B.n550 163.367
R570 B.n547 B.n546 163.367
R571 B.n543 B.n542 163.367
R572 B.n539 B.n538 163.367
R573 B.n535 B.n534 163.367
R574 B.n531 B.n530 163.367
R575 B.n527 B.n526 163.367
R576 B.n523 B.n522 163.367
R577 B.n519 B.n518 163.367
R578 B.n515 B.n514 163.367
R579 B.n511 B.n510 163.367
R580 B.n507 B.n506 163.367
R581 B.n503 B.n502 163.367
R582 B.n499 B.n498 163.367
R583 B.n495 B.n494 163.367
R584 B.n491 B.n490 163.367
R585 B.n487 B.n486 163.367
R586 B.n483 B.n482 163.367
R587 B.n479 B.n478 163.367
R588 B.n475 B.n474 163.367
R589 B.n471 B.n470 163.367
R590 B.n467 B.n466 163.367
R591 B.n463 B.n462 163.367
R592 B.n459 B.n458 163.367
R593 B.n455 B.n454 163.367
R594 B.n451 B.n450 163.367
R595 B.n447 B.n446 163.367
R596 B.n443 B.n442 163.367
R597 B.n439 B.n438 163.367
R598 B.n435 B.n434 163.367
R599 B.n431 B.n430 163.367
R600 B.n427 B.n426 163.367
R601 B.n423 B.n422 163.367
R602 B.n419 B.n418 163.367
R603 B.n415 B.n414 163.367
R604 B.n633 B.n350 163.367
R605 B.n637 B.n348 163.367
R606 B.n637 B.n341 163.367
R607 B.n645 B.n341 163.367
R608 B.n645 B.n339 163.367
R609 B.n649 B.n339 163.367
R610 B.n649 B.n334 163.367
R611 B.n657 B.n334 163.367
R612 B.n657 B.n332 163.367
R613 B.n661 B.n332 163.367
R614 B.n661 B.n327 163.367
R615 B.n670 B.n327 163.367
R616 B.n670 B.n325 163.367
R617 B.n675 B.n325 163.367
R618 B.n675 B.n319 163.367
R619 B.n683 B.n319 163.367
R620 B.n684 B.n683 163.367
R621 B.n684 B.n5 163.367
R622 B.n6 B.n5 163.367
R623 B.n7 B.n6 163.367
R624 B.n689 B.n7 163.367
R625 B.n689 B.n12 163.367
R626 B.n13 B.n12 163.367
R627 B.n14 B.n13 163.367
R628 B.n694 B.n14 163.367
R629 B.n694 B.n19 163.367
R630 B.n20 B.n19 163.367
R631 B.n21 B.n20 163.367
R632 B.n699 B.n21 163.367
R633 B.n699 B.n26 163.367
R634 B.n27 B.n26 163.367
R635 B.n28 B.n27 163.367
R636 B.n704 B.n28 163.367
R637 B.n704 B.n33 163.367
R638 B.n34 B.n33 163.367
R639 B.n99 B.n98 163.367
R640 B.n103 B.n102 163.367
R641 B.n107 B.n106 163.367
R642 B.n111 B.n110 163.367
R643 B.n115 B.n114 163.367
R644 B.n119 B.n118 163.367
R645 B.n123 B.n122 163.367
R646 B.n127 B.n126 163.367
R647 B.n131 B.n130 163.367
R648 B.n135 B.n134 163.367
R649 B.n139 B.n138 163.367
R650 B.n143 B.n142 163.367
R651 B.n147 B.n146 163.367
R652 B.n151 B.n150 163.367
R653 B.n155 B.n154 163.367
R654 B.n159 B.n158 163.367
R655 B.n163 B.n162 163.367
R656 B.n167 B.n166 163.367
R657 B.n171 B.n170 163.367
R658 B.n175 B.n174 163.367
R659 B.n179 B.n178 163.367
R660 B.n183 B.n182 163.367
R661 B.n187 B.n186 163.367
R662 B.n191 B.n190 163.367
R663 B.n195 B.n194 163.367
R664 B.n200 B.n199 163.367
R665 B.n204 B.n203 163.367
R666 B.n208 B.n207 163.367
R667 B.n212 B.n211 163.367
R668 B.n216 B.n215 163.367
R669 B.n221 B.n220 163.367
R670 B.n225 B.n224 163.367
R671 B.n229 B.n228 163.367
R672 B.n233 B.n232 163.367
R673 B.n237 B.n236 163.367
R674 B.n241 B.n240 163.367
R675 B.n245 B.n244 163.367
R676 B.n249 B.n248 163.367
R677 B.n253 B.n252 163.367
R678 B.n257 B.n256 163.367
R679 B.n261 B.n260 163.367
R680 B.n265 B.n264 163.367
R681 B.n269 B.n268 163.367
R682 B.n273 B.n272 163.367
R683 B.n277 B.n276 163.367
R684 B.n281 B.n280 163.367
R685 B.n285 B.n284 163.367
R686 B.n289 B.n288 163.367
R687 B.n293 B.n292 163.367
R688 B.n297 B.n296 163.367
R689 B.n301 B.n300 163.367
R690 B.n305 B.n304 163.367
R691 B.n309 B.n308 163.367
R692 B.n313 B.n312 163.367
R693 B.n315 B.n90 163.367
R694 B.n410 B.t17 92.4627
R695 B.n91 B.t13 92.4627
R696 B.n407 B.t11 92.4429
R697 B.n93 B.t6 92.4429
R698 B.n411 B.t16 72.6808
R699 B.n92 B.t14 72.6808
R700 B.n408 B.t10 72.6611
R701 B.n94 B.t7 72.6611
R702 B.n631 B.n630 71.676
R703 B.n625 B.n351 71.676
R704 B.n622 B.n352 71.676
R705 B.n618 B.n353 71.676
R706 B.n614 B.n354 71.676
R707 B.n610 B.n355 71.676
R708 B.n606 B.n356 71.676
R709 B.n602 B.n357 71.676
R710 B.n598 B.n358 71.676
R711 B.n594 B.n359 71.676
R712 B.n590 B.n360 71.676
R713 B.n586 B.n361 71.676
R714 B.n582 B.n362 71.676
R715 B.n578 B.n363 71.676
R716 B.n574 B.n364 71.676
R717 B.n570 B.n365 71.676
R718 B.n566 B.n366 71.676
R719 B.n562 B.n367 71.676
R720 B.n558 B.n368 71.676
R721 B.n554 B.n369 71.676
R722 B.n550 B.n370 71.676
R723 B.n546 B.n371 71.676
R724 B.n542 B.n372 71.676
R725 B.n538 B.n373 71.676
R726 B.n534 B.n374 71.676
R727 B.n530 B.n375 71.676
R728 B.n526 B.n376 71.676
R729 B.n522 B.n377 71.676
R730 B.n518 B.n378 71.676
R731 B.n514 B.n379 71.676
R732 B.n510 B.n380 71.676
R733 B.n506 B.n381 71.676
R734 B.n502 B.n382 71.676
R735 B.n498 B.n383 71.676
R736 B.n494 B.n384 71.676
R737 B.n490 B.n385 71.676
R738 B.n486 B.n386 71.676
R739 B.n482 B.n387 71.676
R740 B.n478 B.n388 71.676
R741 B.n474 B.n389 71.676
R742 B.n470 B.n390 71.676
R743 B.n466 B.n391 71.676
R744 B.n462 B.n392 71.676
R745 B.n458 B.n393 71.676
R746 B.n454 B.n394 71.676
R747 B.n450 B.n395 71.676
R748 B.n446 B.n396 71.676
R749 B.n442 B.n397 71.676
R750 B.n438 B.n398 71.676
R751 B.n434 B.n399 71.676
R752 B.n430 B.n400 71.676
R753 B.n426 B.n401 71.676
R754 B.n422 B.n402 71.676
R755 B.n418 B.n403 71.676
R756 B.n414 B.n404 71.676
R757 B.n95 B.n35 71.676
R758 B.n99 B.n36 71.676
R759 B.n103 B.n37 71.676
R760 B.n107 B.n38 71.676
R761 B.n111 B.n39 71.676
R762 B.n115 B.n40 71.676
R763 B.n119 B.n41 71.676
R764 B.n123 B.n42 71.676
R765 B.n127 B.n43 71.676
R766 B.n131 B.n44 71.676
R767 B.n135 B.n45 71.676
R768 B.n139 B.n46 71.676
R769 B.n143 B.n47 71.676
R770 B.n147 B.n48 71.676
R771 B.n151 B.n49 71.676
R772 B.n155 B.n50 71.676
R773 B.n159 B.n51 71.676
R774 B.n163 B.n52 71.676
R775 B.n167 B.n53 71.676
R776 B.n171 B.n54 71.676
R777 B.n175 B.n55 71.676
R778 B.n179 B.n56 71.676
R779 B.n183 B.n57 71.676
R780 B.n187 B.n58 71.676
R781 B.n191 B.n59 71.676
R782 B.n195 B.n60 71.676
R783 B.n200 B.n61 71.676
R784 B.n204 B.n62 71.676
R785 B.n208 B.n63 71.676
R786 B.n212 B.n64 71.676
R787 B.n216 B.n65 71.676
R788 B.n221 B.n66 71.676
R789 B.n225 B.n67 71.676
R790 B.n229 B.n68 71.676
R791 B.n233 B.n69 71.676
R792 B.n237 B.n70 71.676
R793 B.n241 B.n71 71.676
R794 B.n245 B.n72 71.676
R795 B.n249 B.n73 71.676
R796 B.n253 B.n74 71.676
R797 B.n257 B.n75 71.676
R798 B.n261 B.n76 71.676
R799 B.n265 B.n77 71.676
R800 B.n269 B.n78 71.676
R801 B.n273 B.n79 71.676
R802 B.n277 B.n80 71.676
R803 B.n281 B.n81 71.676
R804 B.n285 B.n82 71.676
R805 B.n289 B.n83 71.676
R806 B.n293 B.n84 71.676
R807 B.n297 B.n85 71.676
R808 B.n301 B.n86 71.676
R809 B.n305 B.n87 71.676
R810 B.n309 B.n88 71.676
R811 B.n313 B.n89 71.676
R812 B.n710 B.n90 71.676
R813 B.n710 B.n709 71.676
R814 B.n315 B.n89 71.676
R815 B.n312 B.n88 71.676
R816 B.n308 B.n87 71.676
R817 B.n304 B.n86 71.676
R818 B.n300 B.n85 71.676
R819 B.n296 B.n84 71.676
R820 B.n292 B.n83 71.676
R821 B.n288 B.n82 71.676
R822 B.n284 B.n81 71.676
R823 B.n280 B.n80 71.676
R824 B.n276 B.n79 71.676
R825 B.n272 B.n78 71.676
R826 B.n268 B.n77 71.676
R827 B.n264 B.n76 71.676
R828 B.n260 B.n75 71.676
R829 B.n256 B.n74 71.676
R830 B.n252 B.n73 71.676
R831 B.n248 B.n72 71.676
R832 B.n244 B.n71 71.676
R833 B.n240 B.n70 71.676
R834 B.n236 B.n69 71.676
R835 B.n232 B.n68 71.676
R836 B.n228 B.n67 71.676
R837 B.n224 B.n66 71.676
R838 B.n220 B.n65 71.676
R839 B.n215 B.n64 71.676
R840 B.n211 B.n63 71.676
R841 B.n207 B.n62 71.676
R842 B.n203 B.n61 71.676
R843 B.n199 B.n60 71.676
R844 B.n194 B.n59 71.676
R845 B.n190 B.n58 71.676
R846 B.n186 B.n57 71.676
R847 B.n182 B.n56 71.676
R848 B.n178 B.n55 71.676
R849 B.n174 B.n54 71.676
R850 B.n170 B.n53 71.676
R851 B.n166 B.n52 71.676
R852 B.n162 B.n51 71.676
R853 B.n158 B.n50 71.676
R854 B.n154 B.n49 71.676
R855 B.n150 B.n48 71.676
R856 B.n146 B.n47 71.676
R857 B.n142 B.n46 71.676
R858 B.n138 B.n45 71.676
R859 B.n134 B.n44 71.676
R860 B.n130 B.n43 71.676
R861 B.n126 B.n42 71.676
R862 B.n122 B.n41 71.676
R863 B.n118 B.n40 71.676
R864 B.n114 B.n39 71.676
R865 B.n110 B.n38 71.676
R866 B.n106 B.n37 71.676
R867 B.n102 B.n36 71.676
R868 B.n98 B.n35 71.676
R869 B.n631 B.n406 71.676
R870 B.n623 B.n351 71.676
R871 B.n619 B.n352 71.676
R872 B.n615 B.n353 71.676
R873 B.n611 B.n354 71.676
R874 B.n607 B.n355 71.676
R875 B.n603 B.n356 71.676
R876 B.n599 B.n357 71.676
R877 B.n595 B.n358 71.676
R878 B.n591 B.n359 71.676
R879 B.n587 B.n360 71.676
R880 B.n583 B.n361 71.676
R881 B.n579 B.n362 71.676
R882 B.n575 B.n363 71.676
R883 B.n571 B.n364 71.676
R884 B.n567 B.n365 71.676
R885 B.n563 B.n366 71.676
R886 B.n559 B.n367 71.676
R887 B.n555 B.n368 71.676
R888 B.n551 B.n369 71.676
R889 B.n547 B.n370 71.676
R890 B.n543 B.n371 71.676
R891 B.n539 B.n372 71.676
R892 B.n535 B.n373 71.676
R893 B.n531 B.n374 71.676
R894 B.n527 B.n375 71.676
R895 B.n523 B.n376 71.676
R896 B.n519 B.n377 71.676
R897 B.n515 B.n378 71.676
R898 B.n511 B.n379 71.676
R899 B.n507 B.n380 71.676
R900 B.n503 B.n381 71.676
R901 B.n499 B.n382 71.676
R902 B.n495 B.n383 71.676
R903 B.n491 B.n384 71.676
R904 B.n487 B.n385 71.676
R905 B.n483 B.n386 71.676
R906 B.n479 B.n387 71.676
R907 B.n475 B.n388 71.676
R908 B.n471 B.n389 71.676
R909 B.n467 B.n390 71.676
R910 B.n463 B.n391 71.676
R911 B.n459 B.n392 71.676
R912 B.n455 B.n393 71.676
R913 B.n451 B.n394 71.676
R914 B.n447 B.n395 71.676
R915 B.n443 B.n396 71.676
R916 B.n439 B.n397 71.676
R917 B.n435 B.n398 71.676
R918 B.n431 B.n399 71.676
R919 B.n427 B.n400 71.676
R920 B.n423 B.n401 71.676
R921 B.n419 B.n402 71.676
R922 B.n415 B.n403 71.676
R923 B.n404 B.n350 71.676
R924 B.n632 B.n347 70.276
R925 B.n712 B.n711 70.276
R926 B.n412 B.n411 59.5399
R927 B.n409 B.n408 59.5399
R928 B.n197 B.n94 59.5399
R929 B.n218 B.n92 59.5399
R930 B.n638 B.n347 36.4794
R931 B.n638 B.n342 36.4794
R932 B.n644 B.n342 36.4794
R933 B.n644 B.n343 36.4794
R934 B.n650 B.n335 36.4794
R935 B.n656 B.n335 36.4794
R936 B.n656 B.n331 36.4794
R937 B.n663 B.n331 36.4794
R938 B.n663 B.n662 36.4794
R939 B.n669 B.n324 36.4794
R940 B.n676 B.n324 36.4794
R941 B.n682 B.n320 36.4794
R942 B.n682 B.n4 36.4794
R943 B.n745 B.n4 36.4794
R944 B.n745 B.n744 36.4794
R945 B.n744 B.n743 36.4794
R946 B.n743 B.n8 36.4794
R947 B.n737 B.n736 36.4794
R948 B.n736 B.n735 36.4794
R949 B.n729 B.n18 36.4794
R950 B.n729 B.n728 36.4794
R951 B.n728 B.n727 36.4794
R952 B.n727 B.n22 36.4794
R953 B.n721 B.n22 36.4794
R954 B.n720 B.n719 36.4794
R955 B.n719 B.n29 36.4794
R956 B.n713 B.n29 36.4794
R957 B.n713 B.n712 36.4794
R958 B.n662 B.t0 32.7242
R959 B.n676 B.t2 32.7242
R960 B.n737 B.t3 32.7242
R961 B.n18 B.t1 32.7242
R962 B.n96 B.n31 32.6249
R963 B.n708 B.n707 32.6249
R964 B.n635 B.n634 32.6249
R965 B.n629 B.n345 32.6249
R966 B.n343 B.t9 25.2139
R967 B.t5 B.n720 25.2139
R968 B.n411 B.n410 19.7823
R969 B.n408 B.n407 19.7823
R970 B.n94 B.n93 19.7823
R971 B.n92 B.n91 19.7823
R972 B B.n747 18.0485
R973 B.n650 B.t9 11.266
R974 B.n721 B.t5 11.266
R975 B.n97 B.n96 10.6151
R976 B.n100 B.n97 10.6151
R977 B.n101 B.n100 10.6151
R978 B.n104 B.n101 10.6151
R979 B.n105 B.n104 10.6151
R980 B.n108 B.n105 10.6151
R981 B.n109 B.n108 10.6151
R982 B.n112 B.n109 10.6151
R983 B.n113 B.n112 10.6151
R984 B.n116 B.n113 10.6151
R985 B.n117 B.n116 10.6151
R986 B.n120 B.n117 10.6151
R987 B.n121 B.n120 10.6151
R988 B.n124 B.n121 10.6151
R989 B.n125 B.n124 10.6151
R990 B.n128 B.n125 10.6151
R991 B.n129 B.n128 10.6151
R992 B.n132 B.n129 10.6151
R993 B.n133 B.n132 10.6151
R994 B.n136 B.n133 10.6151
R995 B.n137 B.n136 10.6151
R996 B.n140 B.n137 10.6151
R997 B.n141 B.n140 10.6151
R998 B.n144 B.n141 10.6151
R999 B.n145 B.n144 10.6151
R1000 B.n148 B.n145 10.6151
R1001 B.n149 B.n148 10.6151
R1002 B.n152 B.n149 10.6151
R1003 B.n153 B.n152 10.6151
R1004 B.n156 B.n153 10.6151
R1005 B.n157 B.n156 10.6151
R1006 B.n160 B.n157 10.6151
R1007 B.n161 B.n160 10.6151
R1008 B.n164 B.n161 10.6151
R1009 B.n165 B.n164 10.6151
R1010 B.n168 B.n165 10.6151
R1011 B.n169 B.n168 10.6151
R1012 B.n172 B.n169 10.6151
R1013 B.n173 B.n172 10.6151
R1014 B.n176 B.n173 10.6151
R1015 B.n177 B.n176 10.6151
R1016 B.n180 B.n177 10.6151
R1017 B.n181 B.n180 10.6151
R1018 B.n184 B.n181 10.6151
R1019 B.n185 B.n184 10.6151
R1020 B.n188 B.n185 10.6151
R1021 B.n189 B.n188 10.6151
R1022 B.n192 B.n189 10.6151
R1023 B.n193 B.n192 10.6151
R1024 B.n196 B.n193 10.6151
R1025 B.n201 B.n198 10.6151
R1026 B.n202 B.n201 10.6151
R1027 B.n205 B.n202 10.6151
R1028 B.n206 B.n205 10.6151
R1029 B.n209 B.n206 10.6151
R1030 B.n210 B.n209 10.6151
R1031 B.n213 B.n210 10.6151
R1032 B.n214 B.n213 10.6151
R1033 B.n217 B.n214 10.6151
R1034 B.n222 B.n219 10.6151
R1035 B.n223 B.n222 10.6151
R1036 B.n226 B.n223 10.6151
R1037 B.n227 B.n226 10.6151
R1038 B.n230 B.n227 10.6151
R1039 B.n231 B.n230 10.6151
R1040 B.n234 B.n231 10.6151
R1041 B.n235 B.n234 10.6151
R1042 B.n238 B.n235 10.6151
R1043 B.n239 B.n238 10.6151
R1044 B.n242 B.n239 10.6151
R1045 B.n243 B.n242 10.6151
R1046 B.n246 B.n243 10.6151
R1047 B.n247 B.n246 10.6151
R1048 B.n250 B.n247 10.6151
R1049 B.n251 B.n250 10.6151
R1050 B.n254 B.n251 10.6151
R1051 B.n255 B.n254 10.6151
R1052 B.n258 B.n255 10.6151
R1053 B.n259 B.n258 10.6151
R1054 B.n262 B.n259 10.6151
R1055 B.n263 B.n262 10.6151
R1056 B.n266 B.n263 10.6151
R1057 B.n267 B.n266 10.6151
R1058 B.n270 B.n267 10.6151
R1059 B.n271 B.n270 10.6151
R1060 B.n274 B.n271 10.6151
R1061 B.n275 B.n274 10.6151
R1062 B.n278 B.n275 10.6151
R1063 B.n279 B.n278 10.6151
R1064 B.n282 B.n279 10.6151
R1065 B.n283 B.n282 10.6151
R1066 B.n286 B.n283 10.6151
R1067 B.n287 B.n286 10.6151
R1068 B.n290 B.n287 10.6151
R1069 B.n291 B.n290 10.6151
R1070 B.n294 B.n291 10.6151
R1071 B.n295 B.n294 10.6151
R1072 B.n298 B.n295 10.6151
R1073 B.n299 B.n298 10.6151
R1074 B.n302 B.n299 10.6151
R1075 B.n303 B.n302 10.6151
R1076 B.n306 B.n303 10.6151
R1077 B.n307 B.n306 10.6151
R1078 B.n310 B.n307 10.6151
R1079 B.n311 B.n310 10.6151
R1080 B.n314 B.n311 10.6151
R1081 B.n316 B.n314 10.6151
R1082 B.n317 B.n316 10.6151
R1083 B.n708 B.n317 10.6151
R1084 B.n636 B.n635 10.6151
R1085 B.n636 B.n340 10.6151
R1086 B.n646 B.n340 10.6151
R1087 B.n647 B.n646 10.6151
R1088 B.n648 B.n647 10.6151
R1089 B.n648 B.n333 10.6151
R1090 B.n658 B.n333 10.6151
R1091 B.n659 B.n658 10.6151
R1092 B.n660 B.n659 10.6151
R1093 B.n660 B.n326 10.6151
R1094 B.n671 B.n326 10.6151
R1095 B.n672 B.n671 10.6151
R1096 B.n674 B.n672 10.6151
R1097 B.n674 B.n673 10.6151
R1098 B.n673 B.n318 10.6151
R1099 B.n685 B.n318 10.6151
R1100 B.n686 B.n685 10.6151
R1101 B.n687 B.n686 10.6151
R1102 B.n688 B.n687 10.6151
R1103 B.n690 B.n688 10.6151
R1104 B.n691 B.n690 10.6151
R1105 B.n692 B.n691 10.6151
R1106 B.n693 B.n692 10.6151
R1107 B.n695 B.n693 10.6151
R1108 B.n696 B.n695 10.6151
R1109 B.n697 B.n696 10.6151
R1110 B.n698 B.n697 10.6151
R1111 B.n700 B.n698 10.6151
R1112 B.n701 B.n700 10.6151
R1113 B.n702 B.n701 10.6151
R1114 B.n703 B.n702 10.6151
R1115 B.n705 B.n703 10.6151
R1116 B.n706 B.n705 10.6151
R1117 B.n707 B.n706 10.6151
R1118 B.n629 B.n628 10.6151
R1119 B.n628 B.n627 10.6151
R1120 B.n627 B.n626 10.6151
R1121 B.n626 B.n624 10.6151
R1122 B.n624 B.n621 10.6151
R1123 B.n621 B.n620 10.6151
R1124 B.n620 B.n617 10.6151
R1125 B.n617 B.n616 10.6151
R1126 B.n616 B.n613 10.6151
R1127 B.n613 B.n612 10.6151
R1128 B.n612 B.n609 10.6151
R1129 B.n609 B.n608 10.6151
R1130 B.n608 B.n605 10.6151
R1131 B.n605 B.n604 10.6151
R1132 B.n604 B.n601 10.6151
R1133 B.n601 B.n600 10.6151
R1134 B.n600 B.n597 10.6151
R1135 B.n597 B.n596 10.6151
R1136 B.n596 B.n593 10.6151
R1137 B.n593 B.n592 10.6151
R1138 B.n592 B.n589 10.6151
R1139 B.n589 B.n588 10.6151
R1140 B.n588 B.n585 10.6151
R1141 B.n585 B.n584 10.6151
R1142 B.n584 B.n581 10.6151
R1143 B.n581 B.n580 10.6151
R1144 B.n580 B.n577 10.6151
R1145 B.n577 B.n576 10.6151
R1146 B.n576 B.n573 10.6151
R1147 B.n573 B.n572 10.6151
R1148 B.n572 B.n569 10.6151
R1149 B.n569 B.n568 10.6151
R1150 B.n568 B.n565 10.6151
R1151 B.n565 B.n564 10.6151
R1152 B.n564 B.n561 10.6151
R1153 B.n561 B.n560 10.6151
R1154 B.n560 B.n557 10.6151
R1155 B.n557 B.n556 10.6151
R1156 B.n556 B.n553 10.6151
R1157 B.n553 B.n552 10.6151
R1158 B.n552 B.n549 10.6151
R1159 B.n549 B.n548 10.6151
R1160 B.n548 B.n545 10.6151
R1161 B.n545 B.n544 10.6151
R1162 B.n544 B.n541 10.6151
R1163 B.n541 B.n540 10.6151
R1164 B.n540 B.n537 10.6151
R1165 B.n537 B.n536 10.6151
R1166 B.n536 B.n533 10.6151
R1167 B.n533 B.n532 10.6151
R1168 B.n529 B.n528 10.6151
R1169 B.n528 B.n525 10.6151
R1170 B.n525 B.n524 10.6151
R1171 B.n524 B.n521 10.6151
R1172 B.n521 B.n520 10.6151
R1173 B.n520 B.n517 10.6151
R1174 B.n517 B.n516 10.6151
R1175 B.n516 B.n513 10.6151
R1176 B.n513 B.n512 10.6151
R1177 B.n509 B.n508 10.6151
R1178 B.n508 B.n505 10.6151
R1179 B.n505 B.n504 10.6151
R1180 B.n504 B.n501 10.6151
R1181 B.n501 B.n500 10.6151
R1182 B.n500 B.n497 10.6151
R1183 B.n497 B.n496 10.6151
R1184 B.n496 B.n493 10.6151
R1185 B.n493 B.n492 10.6151
R1186 B.n492 B.n489 10.6151
R1187 B.n489 B.n488 10.6151
R1188 B.n488 B.n485 10.6151
R1189 B.n485 B.n484 10.6151
R1190 B.n484 B.n481 10.6151
R1191 B.n481 B.n480 10.6151
R1192 B.n480 B.n477 10.6151
R1193 B.n477 B.n476 10.6151
R1194 B.n476 B.n473 10.6151
R1195 B.n473 B.n472 10.6151
R1196 B.n472 B.n469 10.6151
R1197 B.n469 B.n468 10.6151
R1198 B.n468 B.n465 10.6151
R1199 B.n465 B.n464 10.6151
R1200 B.n464 B.n461 10.6151
R1201 B.n461 B.n460 10.6151
R1202 B.n460 B.n457 10.6151
R1203 B.n457 B.n456 10.6151
R1204 B.n456 B.n453 10.6151
R1205 B.n453 B.n452 10.6151
R1206 B.n452 B.n449 10.6151
R1207 B.n449 B.n448 10.6151
R1208 B.n448 B.n445 10.6151
R1209 B.n445 B.n444 10.6151
R1210 B.n444 B.n441 10.6151
R1211 B.n441 B.n440 10.6151
R1212 B.n440 B.n437 10.6151
R1213 B.n437 B.n436 10.6151
R1214 B.n436 B.n433 10.6151
R1215 B.n433 B.n432 10.6151
R1216 B.n432 B.n429 10.6151
R1217 B.n429 B.n428 10.6151
R1218 B.n428 B.n425 10.6151
R1219 B.n425 B.n424 10.6151
R1220 B.n424 B.n421 10.6151
R1221 B.n421 B.n420 10.6151
R1222 B.n420 B.n417 10.6151
R1223 B.n417 B.n416 10.6151
R1224 B.n416 B.n413 10.6151
R1225 B.n413 B.n349 10.6151
R1226 B.n634 B.n349 10.6151
R1227 B.n640 B.n345 10.6151
R1228 B.n641 B.n640 10.6151
R1229 B.n642 B.n641 10.6151
R1230 B.n642 B.n337 10.6151
R1231 B.n652 B.n337 10.6151
R1232 B.n653 B.n652 10.6151
R1233 B.n654 B.n653 10.6151
R1234 B.n654 B.n329 10.6151
R1235 B.n665 B.n329 10.6151
R1236 B.n666 B.n665 10.6151
R1237 B.n667 B.n666 10.6151
R1238 B.n667 B.n322 10.6151
R1239 B.n678 B.n322 10.6151
R1240 B.n679 B.n678 10.6151
R1241 B.n680 B.n679 10.6151
R1242 B.n680 B.n0 10.6151
R1243 B.n741 B.n1 10.6151
R1244 B.n741 B.n740 10.6151
R1245 B.n740 B.n739 10.6151
R1246 B.n739 B.n10 10.6151
R1247 B.n733 B.n10 10.6151
R1248 B.n733 B.n732 10.6151
R1249 B.n732 B.n731 10.6151
R1250 B.n731 B.n16 10.6151
R1251 B.n725 B.n16 10.6151
R1252 B.n725 B.n724 10.6151
R1253 B.n724 B.n723 10.6151
R1254 B.n723 B.n24 10.6151
R1255 B.n717 B.n24 10.6151
R1256 B.n717 B.n716 10.6151
R1257 B.n716 B.n715 10.6151
R1258 B.n715 B.n31 10.6151
R1259 B.n197 B.n196 9.36635
R1260 B.n219 B.n218 9.36635
R1261 B.n532 B.n409 9.36635
R1262 B.n509 B.n412 9.36635
R1263 B.n669 B.t0 3.75568
R1264 B.t2 B.n320 3.75568
R1265 B.t3 B.n8 3.75568
R1266 B.n735 B.t1 3.75568
R1267 B.n747 B.n0 2.81026
R1268 B.n747 B.n1 2.81026
R1269 B.n198 B.n197 1.24928
R1270 B.n218 B.n217 1.24928
R1271 B.n529 B.n409 1.24928
R1272 B.n512 B.n412 1.24928
R1273 VP.n1 VP.t1 610.225
R1274 VP.n1 VP.t3 610.174
R1275 VP.n3 VP.t0 589.229
R1276 VP.n5 VP.t2 589.229
R1277 VP.n6 VP.n5 161.3
R1278 VP.n4 VP.n0 161.3
R1279 VP.n3 VP.n2 161.3
R1280 VP.n2 VP.n1 87.4803
R1281 VP.n4 VP.n3 24.1005
R1282 VP.n5 VP.n4 24.1005
R1283 VP.n2 VP.n0 0.189894
R1284 VP.n6 VP.n0 0.189894
R1285 VP VP.n6 0.0516364
R1286 VDD1 VDD1.n1 105.347
R1287 VDD1 VDD1.n0 65.3984
R1288 VDD1.n0 VDD1.t2 1.30057
R1289 VDD1.n0 VDD1.t0 1.30057
R1290 VDD1.n1 VDD1.t3 1.30057
R1291 VDD1.n1 VDD1.t1 1.30057
C0 VDD1 VDD2 0.564133f
C1 VTAIL VDD1 8.267079f
C2 VP VDD1 4.03628f
C3 VN VDD2 3.91104f
C4 VTAIL VN 3.38163f
C5 VP VN 5.41525f
C6 VTAIL VDD2 8.30848f
C7 VP VDD2 0.272575f
C8 VN VDD1 0.14708f
C9 VP VTAIL 3.39573f
C10 VDD2 B 2.946175f
C11 VDD1 B 7.05272f
C12 VTAIL B 10.589967f
C13 VN B 8.60707f
C14 VP B 5.09647f
C15 VDD1.t2 B 0.340782f
C16 VDD1.t0 B 0.340782f
C17 VDD1.n0 B 3.08797f
C18 VDD1.t3 B 0.340782f
C19 VDD1.t1 B 0.340782f
C20 VDD1.n1 B 3.81298f
C21 VP.n0 B 0.050012f
C22 VP.t3 B 1.51325f
C23 VP.t1 B 1.5133f
C24 VP.n1 B 2.2101f
C25 VP.n2 B 3.31576f
C26 VP.t0 B 1.49351f
C27 VP.n3 B 0.571364f
C28 VP.n4 B 0.011349f
C29 VP.t2 B 1.49351f
C30 VP.n5 B 0.571364f
C31 VP.n6 B 0.038758f
C32 VTAIL.t7 B 2.19006f
C33 VTAIL.n0 B 0.254093f
C34 VTAIL.t2 B 2.19006f
C35 VTAIL.n1 B 0.273905f
C36 VTAIL.t0 B 2.19006f
C37 VTAIL.n2 B 1.19598f
C38 VTAIL.t4 B 2.19006f
C39 VTAIL.n3 B 1.19598f
C40 VTAIL.t5 B 2.19006f
C41 VTAIL.n4 B 0.273903f
C42 VTAIL.t3 B 2.19006f
C43 VTAIL.n5 B 0.273903f
C44 VTAIL.t1 B 2.19006f
C45 VTAIL.n6 B 1.19598f
C46 VTAIL.t6 B 2.19006f
C47 VTAIL.n7 B 1.17013f
C48 VDD2.t0 B 0.34091f
C49 VDD2.t3 B 0.34091f
C50 VDD2.n0 B 3.787f
C51 VDD2.t1 B 0.34091f
C52 VDD2.t2 B 0.34091f
C53 VDD2.n1 B 3.08884f
C54 VDD2.n2 B 3.87416f
C55 VN.t0 B 1.49328f
C56 VN.t1 B 1.49322f
C57 VN.n0 B 1.10029f
C58 VN.t2 B 1.49328f
C59 VN.t3 B 1.49322f
C60 VN.n1 B 2.20165f
.ends

