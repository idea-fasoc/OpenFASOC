* NGSPICE file created from diff_pair_sample_1298.ext - technology: sky130A

.subckt diff_pair_sample_1298 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.04425 pd=18.78 as=7.1955 ps=37.68 w=18.45 l=1.78
X1 VTAIL.t5 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=3.04425 ps=18.78 w=18.45 l=1.78
X2 VTAIL.t4 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=3.04425 ps=18.78 w=18.45 l=1.78
X3 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.04425 pd=18.78 as=7.1955 ps=37.68 w=18.45 l=1.78
X4 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.04425 pd=18.78 as=7.1955 ps=37.68 w=18.45 l=1.78
X5 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=0 ps=0 w=18.45 l=1.78
X6 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=3.04425 ps=18.78 w=18.45 l=1.78
X7 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=0 ps=0 w=18.45 l=1.78
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=0 ps=0 w=18.45 l=1.78
X9 VDD2.t0 VN.t3 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.04425 pd=18.78 as=7.1955 ps=37.68 w=18.45 l=1.78
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=0 ps=0 w=18.45 l=1.78
X11 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1955 pd=37.68 as=3.04425 ps=18.78 w=18.45 l=1.78
R0 VN.n0 VN.t2 286.048
R1 VN.n1 VN.t3 286.048
R2 VN.n0 VN.t0 285.618
R3 VN.n1 VN.t1 285.618
R4 VN VN.n1 58.3248
R5 VN VN.n0 9.36643
R6 VTAIL.n5 VTAIL.t3 48.6049
R7 VTAIL.n4 VTAIL.t6 48.6049
R8 VTAIL.n3 VTAIL.t5 48.6049
R9 VTAIL.n7 VTAIL.t7 48.6039
R10 VTAIL.n0 VTAIL.t4 48.6039
R11 VTAIL.n1 VTAIL.t0 48.6039
R12 VTAIL.n2 VTAIL.t1 48.6039
R13 VTAIL.n6 VTAIL.t2 48.6038
R14 VTAIL.n7 VTAIL.n6 30.091
R15 VTAIL.n3 VTAIL.n2 30.091
R16 VTAIL.n4 VTAIL.n3 1.81947
R17 VTAIL.n6 VTAIL.n5 1.81947
R18 VTAIL.n2 VTAIL.n1 1.81947
R19 VTAIL VTAIL.n0 0.968172
R20 VTAIL VTAIL.n7 0.851793
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 109.287
R24 VDD2.n2 VDD2.n1 64.2095
R25 VDD2.n1 VDD2.t2 1.07367
R26 VDD2.n1 VDD2.t0 1.07367
R27 VDD2.n0 VDD2.t1 1.07367
R28 VDD2.n0 VDD2.t3 1.07367
R29 VDD2 VDD2.n2 0.0586897
R30 B.n619 B.n122 585
R31 B.n122 B.n51 585
R32 B.n621 B.n620 585
R33 B.n623 B.n121 585
R34 B.n626 B.n625 585
R35 B.n627 B.n120 585
R36 B.n629 B.n628 585
R37 B.n631 B.n119 585
R38 B.n634 B.n633 585
R39 B.n635 B.n118 585
R40 B.n637 B.n636 585
R41 B.n639 B.n117 585
R42 B.n642 B.n641 585
R43 B.n643 B.n116 585
R44 B.n645 B.n644 585
R45 B.n647 B.n115 585
R46 B.n650 B.n649 585
R47 B.n651 B.n114 585
R48 B.n653 B.n652 585
R49 B.n655 B.n113 585
R50 B.n658 B.n657 585
R51 B.n659 B.n112 585
R52 B.n661 B.n660 585
R53 B.n663 B.n111 585
R54 B.n666 B.n665 585
R55 B.n667 B.n110 585
R56 B.n669 B.n668 585
R57 B.n671 B.n109 585
R58 B.n674 B.n673 585
R59 B.n675 B.n108 585
R60 B.n677 B.n676 585
R61 B.n679 B.n107 585
R62 B.n682 B.n681 585
R63 B.n683 B.n106 585
R64 B.n685 B.n684 585
R65 B.n687 B.n105 585
R66 B.n690 B.n689 585
R67 B.n691 B.n104 585
R68 B.n693 B.n692 585
R69 B.n695 B.n103 585
R70 B.n698 B.n697 585
R71 B.n699 B.n102 585
R72 B.n701 B.n700 585
R73 B.n703 B.n101 585
R74 B.n706 B.n705 585
R75 B.n707 B.n100 585
R76 B.n709 B.n708 585
R77 B.n711 B.n99 585
R78 B.n714 B.n713 585
R79 B.n715 B.n98 585
R80 B.n717 B.n716 585
R81 B.n719 B.n97 585
R82 B.n722 B.n721 585
R83 B.n723 B.n96 585
R84 B.n725 B.n724 585
R85 B.n727 B.n95 585
R86 B.n730 B.n729 585
R87 B.n731 B.n94 585
R88 B.n733 B.n732 585
R89 B.n735 B.n93 585
R90 B.n737 B.n736 585
R91 B.n739 B.n738 585
R92 B.n742 B.n741 585
R93 B.n743 B.n88 585
R94 B.n745 B.n744 585
R95 B.n747 B.n87 585
R96 B.n750 B.n749 585
R97 B.n751 B.n86 585
R98 B.n753 B.n752 585
R99 B.n755 B.n85 585
R100 B.n758 B.n757 585
R101 B.n760 B.n82 585
R102 B.n762 B.n761 585
R103 B.n764 B.n81 585
R104 B.n767 B.n766 585
R105 B.n768 B.n80 585
R106 B.n770 B.n769 585
R107 B.n772 B.n79 585
R108 B.n775 B.n774 585
R109 B.n776 B.n78 585
R110 B.n778 B.n777 585
R111 B.n780 B.n77 585
R112 B.n783 B.n782 585
R113 B.n784 B.n76 585
R114 B.n786 B.n785 585
R115 B.n788 B.n75 585
R116 B.n791 B.n790 585
R117 B.n792 B.n74 585
R118 B.n794 B.n793 585
R119 B.n796 B.n73 585
R120 B.n799 B.n798 585
R121 B.n800 B.n72 585
R122 B.n802 B.n801 585
R123 B.n804 B.n71 585
R124 B.n807 B.n806 585
R125 B.n808 B.n70 585
R126 B.n810 B.n809 585
R127 B.n812 B.n69 585
R128 B.n815 B.n814 585
R129 B.n816 B.n68 585
R130 B.n818 B.n817 585
R131 B.n820 B.n67 585
R132 B.n823 B.n822 585
R133 B.n824 B.n66 585
R134 B.n826 B.n825 585
R135 B.n828 B.n65 585
R136 B.n831 B.n830 585
R137 B.n832 B.n64 585
R138 B.n834 B.n833 585
R139 B.n836 B.n63 585
R140 B.n839 B.n838 585
R141 B.n840 B.n62 585
R142 B.n842 B.n841 585
R143 B.n844 B.n61 585
R144 B.n847 B.n846 585
R145 B.n848 B.n60 585
R146 B.n850 B.n849 585
R147 B.n852 B.n59 585
R148 B.n855 B.n854 585
R149 B.n856 B.n58 585
R150 B.n858 B.n857 585
R151 B.n860 B.n57 585
R152 B.n863 B.n862 585
R153 B.n864 B.n56 585
R154 B.n866 B.n865 585
R155 B.n868 B.n55 585
R156 B.n871 B.n870 585
R157 B.n872 B.n54 585
R158 B.n874 B.n873 585
R159 B.n876 B.n53 585
R160 B.n879 B.n878 585
R161 B.n880 B.n52 585
R162 B.n618 B.n50 585
R163 B.n883 B.n50 585
R164 B.n617 B.n49 585
R165 B.n884 B.n49 585
R166 B.n616 B.n48 585
R167 B.n885 B.n48 585
R168 B.n615 B.n614 585
R169 B.n614 B.n44 585
R170 B.n613 B.n43 585
R171 B.n891 B.n43 585
R172 B.n612 B.n42 585
R173 B.n892 B.n42 585
R174 B.n611 B.n41 585
R175 B.n893 B.n41 585
R176 B.n610 B.n609 585
R177 B.n609 B.n37 585
R178 B.n608 B.n36 585
R179 B.n899 B.n36 585
R180 B.n607 B.n35 585
R181 B.n900 B.n35 585
R182 B.n606 B.n34 585
R183 B.n901 B.n34 585
R184 B.n605 B.n604 585
R185 B.n604 B.n30 585
R186 B.n603 B.n29 585
R187 B.n907 B.n29 585
R188 B.n602 B.n28 585
R189 B.n908 B.n28 585
R190 B.n601 B.n27 585
R191 B.n909 B.n27 585
R192 B.n600 B.n599 585
R193 B.n599 B.n26 585
R194 B.n598 B.n22 585
R195 B.n915 B.n22 585
R196 B.n597 B.n21 585
R197 B.n916 B.n21 585
R198 B.n596 B.n20 585
R199 B.n917 B.n20 585
R200 B.n595 B.n594 585
R201 B.n594 B.n16 585
R202 B.n593 B.n15 585
R203 B.n923 B.n15 585
R204 B.n592 B.n14 585
R205 B.n924 B.n14 585
R206 B.n591 B.n13 585
R207 B.n925 B.n13 585
R208 B.n590 B.n589 585
R209 B.n589 B.n12 585
R210 B.n588 B.n587 585
R211 B.n588 B.n8 585
R212 B.n586 B.n7 585
R213 B.n932 B.n7 585
R214 B.n585 B.n6 585
R215 B.n933 B.n6 585
R216 B.n584 B.n5 585
R217 B.n934 B.n5 585
R218 B.n583 B.n582 585
R219 B.n582 B.n4 585
R220 B.n581 B.n123 585
R221 B.n581 B.n580 585
R222 B.n571 B.n124 585
R223 B.n125 B.n124 585
R224 B.n573 B.n572 585
R225 B.n574 B.n573 585
R226 B.n570 B.n129 585
R227 B.n133 B.n129 585
R228 B.n569 B.n568 585
R229 B.n568 B.n567 585
R230 B.n131 B.n130 585
R231 B.n132 B.n131 585
R232 B.n560 B.n559 585
R233 B.n561 B.n560 585
R234 B.n558 B.n138 585
R235 B.n138 B.n137 585
R236 B.n557 B.n556 585
R237 B.n556 B.n555 585
R238 B.n140 B.n139 585
R239 B.n548 B.n140 585
R240 B.n547 B.n546 585
R241 B.n549 B.n547 585
R242 B.n545 B.n145 585
R243 B.n145 B.n144 585
R244 B.n544 B.n543 585
R245 B.n543 B.n542 585
R246 B.n147 B.n146 585
R247 B.n148 B.n147 585
R248 B.n535 B.n534 585
R249 B.n536 B.n535 585
R250 B.n533 B.n153 585
R251 B.n153 B.n152 585
R252 B.n532 B.n531 585
R253 B.n531 B.n530 585
R254 B.n155 B.n154 585
R255 B.n156 B.n155 585
R256 B.n523 B.n522 585
R257 B.n524 B.n523 585
R258 B.n521 B.n161 585
R259 B.n161 B.n160 585
R260 B.n520 B.n519 585
R261 B.n519 B.n518 585
R262 B.n163 B.n162 585
R263 B.n164 B.n163 585
R264 B.n511 B.n510 585
R265 B.n512 B.n511 585
R266 B.n509 B.n169 585
R267 B.n169 B.n168 585
R268 B.n508 B.n507 585
R269 B.n507 B.n506 585
R270 B.n503 B.n173 585
R271 B.n502 B.n501 585
R272 B.n499 B.n174 585
R273 B.n499 B.n172 585
R274 B.n498 B.n497 585
R275 B.n496 B.n495 585
R276 B.n494 B.n176 585
R277 B.n492 B.n491 585
R278 B.n490 B.n177 585
R279 B.n489 B.n488 585
R280 B.n486 B.n178 585
R281 B.n484 B.n483 585
R282 B.n482 B.n179 585
R283 B.n481 B.n480 585
R284 B.n478 B.n180 585
R285 B.n476 B.n475 585
R286 B.n474 B.n181 585
R287 B.n473 B.n472 585
R288 B.n470 B.n182 585
R289 B.n468 B.n467 585
R290 B.n466 B.n183 585
R291 B.n465 B.n464 585
R292 B.n462 B.n184 585
R293 B.n460 B.n459 585
R294 B.n458 B.n185 585
R295 B.n457 B.n456 585
R296 B.n454 B.n186 585
R297 B.n452 B.n451 585
R298 B.n450 B.n187 585
R299 B.n449 B.n448 585
R300 B.n446 B.n188 585
R301 B.n444 B.n443 585
R302 B.n442 B.n189 585
R303 B.n441 B.n440 585
R304 B.n438 B.n190 585
R305 B.n436 B.n435 585
R306 B.n434 B.n191 585
R307 B.n433 B.n432 585
R308 B.n430 B.n192 585
R309 B.n428 B.n427 585
R310 B.n426 B.n193 585
R311 B.n425 B.n424 585
R312 B.n422 B.n194 585
R313 B.n420 B.n419 585
R314 B.n418 B.n195 585
R315 B.n417 B.n416 585
R316 B.n414 B.n196 585
R317 B.n412 B.n411 585
R318 B.n410 B.n197 585
R319 B.n409 B.n408 585
R320 B.n406 B.n198 585
R321 B.n404 B.n403 585
R322 B.n402 B.n199 585
R323 B.n401 B.n400 585
R324 B.n398 B.n200 585
R325 B.n396 B.n395 585
R326 B.n394 B.n201 585
R327 B.n393 B.n392 585
R328 B.n390 B.n202 585
R329 B.n388 B.n387 585
R330 B.n386 B.n203 585
R331 B.n385 B.n384 585
R332 B.n382 B.n381 585
R333 B.n380 B.n379 585
R334 B.n378 B.n208 585
R335 B.n376 B.n375 585
R336 B.n374 B.n209 585
R337 B.n373 B.n372 585
R338 B.n370 B.n210 585
R339 B.n368 B.n367 585
R340 B.n366 B.n211 585
R341 B.n364 B.n363 585
R342 B.n361 B.n214 585
R343 B.n359 B.n358 585
R344 B.n357 B.n215 585
R345 B.n356 B.n355 585
R346 B.n353 B.n216 585
R347 B.n351 B.n350 585
R348 B.n349 B.n217 585
R349 B.n348 B.n347 585
R350 B.n345 B.n218 585
R351 B.n343 B.n342 585
R352 B.n341 B.n219 585
R353 B.n340 B.n339 585
R354 B.n337 B.n220 585
R355 B.n335 B.n334 585
R356 B.n333 B.n221 585
R357 B.n332 B.n331 585
R358 B.n329 B.n222 585
R359 B.n327 B.n326 585
R360 B.n325 B.n223 585
R361 B.n324 B.n323 585
R362 B.n321 B.n224 585
R363 B.n319 B.n318 585
R364 B.n317 B.n225 585
R365 B.n316 B.n315 585
R366 B.n313 B.n226 585
R367 B.n311 B.n310 585
R368 B.n309 B.n227 585
R369 B.n308 B.n307 585
R370 B.n305 B.n228 585
R371 B.n303 B.n302 585
R372 B.n301 B.n229 585
R373 B.n300 B.n299 585
R374 B.n297 B.n230 585
R375 B.n295 B.n294 585
R376 B.n293 B.n231 585
R377 B.n292 B.n291 585
R378 B.n289 B.n232 585
R379 B.n287 B.n286 585
R380 B.n285 B.n233 585
R381 B.n284 B.n283 585
R382 B.n281 B.n234 585
R383 B.n279 B.n278 585
R384 B.n277 B.n235 585
R385 B.n276 B.n275 585
R386 B.n273 B.n236 585
R387 B.n271 B.n270 585
R388 B.n269 B.n237 585
R389 B.n268 B.n267 585
R390 B.n265 B.n238 585
R391 B.n263 B.n262 585
R392 B.n261 B.n239 585
R393 B.n260 B.n259 585
R394 B.n257 B.n240 585
R395 B.n255 B.n254 585
R396 B.n253 B.n241 585
R397 B.n252 B.n251 585
R398 B.n249 B.n242 585
R399 B.n247 B.n246 585
R400 B.n245 B.n244 585
R401 B.n171 B.n170 585
R402 B.n505 B.n504 585
R403 B.n506 B.n505 585
R404 B.n167 B.n166 585
R405 B.n168 B.n167 585
R406 B.n514 B.n513 585
R407 B.n513 B.n512 585
R408 B.n515 B.n165 585
R409 B.n165 B.n164 585
R410 B.n517 B.n516 585
R411 B.n518 B.n517 585
R412 B.n159 B.n158 585
R413 B.n160 B.n159 585
R414 B.n526 B.n525 585
R415 B.n525 B.n524 585
R416 B.n527 B.n157 585
R417 B.n157 B.n156 585
R418 B.n529 B.n528 585
R419 B.n530 B.n529 585
R420 B.n151 B.n150 585
R421 B.n152 B.n151 585
R422 B.n538 B.n537 585
R423 B.n537 B.n536 585
R424 B.n539 B.n149 585
R425 B.n149 B.n148 585
R426 B.n541 B.n540 585
R427 B.n542 B.n541 585
R428 B.n143 B.n142 585
R429 B.n144 B.n143 585
R430 B.n551 B.n550 585
R431 B.n550 B.n549 585
R432 B.n552 B.n141 585
R433 B.n548 B.n141 585
R434 B.n554 B.n553 585
R435 B.n555 B.n554 585
R436 B.n136 B.n135 585
R437 B.n137 B.n136 585
R438 B.n563 B.n562 585
R439 B.n562 B.n561 585
R440 B.n564 B.n134 585
R441 B.n134 B.n132 585
R442 B.n566 B.n565 585
R443 B.n567 B.n566 585
R444 B.n128 B.n127 585
R445 B.n133 B.n128 585
R446 B.n576 B.n575 585
R447 B.n575 B.n574 585
R448 B.n577 B.n126 585
R449 B.n126 B.n125 585
R450 B.n579 B.n578 585
R451 B.n580 B.n579 585
R452 B.n3 B.n0 585
R453 B.n4 B.n3 585
R454 B.n931 B.n1 585
R455 B.n932 B.n931 585
R456 B.n930 B.n929 585
R457 B.n930 B.n8 585
R458 B.n928 B.n9 585
R459 B.n12 B.n9 585
R460 B.n927 B.n926 585
R461 B.n926 B.n925 585
R462 B.n11 B.n10 585
R463 B.n924 B.n11 585
R464 B.n922 B.n921 585
R465 B.n923 B.n922 585
R466 B.n920 B.n17 585
R467 B.n17 B.n16 585
R468 B.n919 B.n918 585
R469 B.n918 B.n917 585
R470 B.n19 B.n18 585
R471 B.n916 B.n19 585
R472 B.n914 B.n913 585
R473 B.n915 B.n914 585
R474 B.n912 B.n23 585
R475 B.n26 B.n23 585
R476 B.n911 B.n910 585
R477 B.n910 B.n909 585
R478 B.n25 B.n24 585
R479 B.n908 B.n25 585
R480 B.n906 B.n905 585
R481 B.n907 B.n906 585
R482 B.n904 B.n31 585
R483 B.n31 B.n30 585
R484 B.n903 B.n902 585
R485 B.n902 B.n901 585
R486 B.n33 B.n32 585
R487 B.n900 B.n33 585
R488 B.n898 B.n897 585
R489 B.n899 B.n898 585
R490 B.n896 B.n38 585
R491 B.n38 B.n37 585
R492 B.n895 B.n894 585
R493 B.n894 B.n893 585
R494 B.n40 B.n39 585
R495 B.n892 B.n40 585
R496 B.n890 B.n889 585
R497 B.n891 B.n890 585
R498 B.n888 B.n45 585
R499 B.n45 B.n44 585
R500 B.n887 B.n886 585
R501 B.n886 B.n885 585
R502 B.n47 B.n46 585
R503 B.n884 B.n47 585
R504 B.n882 B.n881 585
R505 B.n883 B.n882 585
R506 B.n935 B.n934 585
R507 B.n933 B.n2 585
R508 B.n882 B.n52 516.524
R509 B.n122 B.n50 516.524
R510 B.n507 B.n171 516.524
R511 B.n505 B.n173 516.524
R512 B.n83 B.t15 456.151
R513 B.n89 B.t8 456.151
R514 B.n212 B.t12 456.151
R515 B.n204 B.t4 456.151
R516 B.n622 B.n51 256.663
R517 B.n624 B.n51 256.663
R518 B.n630 B.n51 256.663
R519 B.n632 B.n51 256.663
R520 B.n638 B.n51 256.663
R521 B.n640 B.n51 256.663
R522 B.n646 B.n51 256.663
R523 B.n648 B.n51 256.663
R524 B.n654 B.n51 256.663
R525 B.n656 B.n51 256.663
R526 B.n662 B.n51 256.663
R527 B.n664 B.n51 256.663
R528 B.n670 B.n51 256.663
R529 B.n672 B.n51 256.663
R530 B.n678 B.n51 256.663
R531 B.n680 B.n51 256.663
R532 B.n686 B.n51 256.663
R533 B.n688 B.n51 256.663
R534 B.n694 B.n51 256.663
R535 B.n696 B.n51 256.663
R536 B.n702 B.n51 256.663
R537 B.n704 B.n51 256.663
R538 B.n710 B.n51 256.663
R539 B.n712 B.n51 256.663
R540 B.n718 B.n51 256.663
R541 B.n720 B.n51 256.663
R542 B.n726 B.n51 256.663
R543 B.n728 B.n51 256.663
R544 B.n734 B.n51 256.663
R545 B.n92 B.n51 256.663
R546 B.n740 B.n51 256.663
R547 B.n746 B.n51 256.663
R548 B.n748 B.n51 256.663
R549 B.n754 B.n51 256.663
R550 B.n756 B.n51 256.663
R551 B.n763 B.n51 256.663
R552 B.n765 B.n51 256.663
R553 B.n771 B.n51 256.663
R554 B.n773 B.n51 256.663
R555 B.n779 B.n51 256.663
R556 B.n781 B.n51 256.663
R557 B.n787 B.n51 256.663
R558 B.n789 B.n51 256.663
R559 B.n795 B.n51 256.663
R560 B.n797 B.n51 256.663
R561 B.n803 B.n51 256.663
R562 B.n805 B.n51 256.663
R563 B.n811 B.n51 256.663
R564 B.n813 B.n51 256.663
R565 B.n819 B.n51 256.663
R566 B.n821 B.n51 256.663
R567 B.n827 B.n51 256.663
R568 B.n829 B.n51 256.663
R569 B.n835 B.n51 256.663
R570 B.n837 B.n51 256.663
R571 B.n843 B.n51 256.663
R572 B.n845 B.n51 256.663
R573 B.n851 B.n51 256.663
R574 B.n853 B.n51 256.663
R575 B.n859 B.n51 256.663
R576 B.n861 B.n51 256.663
R577 B.n867 B.n51 256.663
R578 B.n869 B.n51 256.663
R579 B.n875 B.n51 256.663
R580 B.n877 B.n51 256.663
R581 B.n500 B.n172 256.663
R582 B.n175 B.n172 256.663
R583 B.n493 B.n172 256.663
R584 B.n487 B.n172 256.663
R585 B.n485 B.n172 256.663
R586 B.n479 B.n172 256.663
R587 B.n477 B.n172 256.663
R588 B.n471 B.n172 256.663
R589 B.n469 B.n172 256.663
R590 B.n463 B.n172 256.663
R591 B.n461 B.n172 256.663
R592 B.n455 B.n172 256.663
R593 B.n453 B.n172 256.663
R594 B.n447 B.n172 256.663
R595 B.n445 B.n172 256.663
R596 B.n439 B.n172 256.663
R597 B.n437 B.n172 256.663
R598 B.n431 B.n172 256.663
R599 B.n429 B.n172 256.663
R600 B.n423 B.n172 256.663
R601 B.n421 B.n172 256.663
R602 B.n415 B.n172 256.663
R603 B.n413 B.n172 256.663
R604 B.n407 B.n172 256.663
R605 B.n405 B.n172 256.663
R606 B.n399 B.n172 256.663
R607 B.n397 B.n172 256.663
R608 B.n391 B.n172 256.663
R609 B.n389 B.n172 256.663
R610 B.n383 B.n172 256.663
R611 B.n207 B.n172 256.663
R612 B.n377 B.n172 256.663
R613 B.n371 B.n172 256.663
R614 B.n369 B.n172 256.663
R615 B.n362 B.n172 256.663
R616 B.n360 B.n172 256.663
R617 B.n354 B.n172 256.663
R618 B.n352 B.n172 256.663
R619 B.n346 B.n172 256.663
R620 B.n344 B.n172 256.663
R621 B.n338 B.n172 256.663
R622 B.n336 B.n172 256.663
R623 B.n330 B.n172 256.663
R624 B.n328 B.n172 256.663
R625 B.n322 B.n172 256.663
R626 B.n320 B.n172 256.663
R627 B.n314 B.n172 256.663
R628 B.n312 B.n172 256.663
R629 B.n306 B.n172 256.663
R630 B.n304 B.n172 256.663
R631 B.n298 B.n172 256.663
R632 B.n296 B.n172 256.663
R633 B.n290 B.n172 256.663
R634 B.n288 B.n172 256.663
R635 B.n282 B.n172 256.663
R636 B.n280 B.n172 256.663
R637 B.n274 B.n172 256.663
R638 B.n272 B.n172 256.663
R639 B.n266 B.n172 256.663
R640 B.n264 B.n172 256.663
R641 B.n258 B.n172 256.663
R642 B.n256 B.n172 256.663
R643 B.n250 B.n172 256.663
R644 B.n248 B.n172 256.663
R645 B.n243 B.n172 256.663
R646 B.n937 B.n936 256.663
R647 B.n878 B.n876 163.367
R648 B.n874 B.n54 163.367
R649 B.n870 B.n868 163.367
R650 B.n866 B.n56 163.367
R651 B.n862 B.n860 163.367
R652 B.n858 B.n58 163.367
R653 B.n854 B.n852 163.367
R654 B.n850 B.n60 163.367
R655 B.n846 B.n844 163.367
R656 B.n842 B.n62 163.367
R657 B.n838 B.n836 163.367
R658 B.n834 B.n64 163.367
R659 B.n830 B.n828 163.367
R660 B.n826 B.n66 163.367
R661 B.n822 B.n820 163.367
R662 B.n818 B.n68 163.367
R663 B.n814 B.n812 163.367
R664 B.n810 B.n70 163.367
R665 B.n806 B.n804 163.367
R666 B.n802 B.n72 163.367
R667 B.n798 B.n796 163.367
R668 B.n794 B.n74 163.367
R669 B.n790 B.n788 163.367
R670 B.n786 B.n76 163.367
R671 B.n782 B.n780 163.367
R672 B.n778 B.n78 163.367
R673 B.n774 B.n772 163.367
R674 B.n770 B.n80 163.367
R675 B.n766 B.n764 163.367
R676 B.n762 B.n82 163.367
R677 B.n757 B.n755 163.367
R678 B.n753 B.n86 163.367
R679 B.n749 B.n747 163.367
R680 B.n745 B.n88 163.367
R681 B.n741 B.n739 163.367
R682 B.n736 B.n735 163.367
R683 B.n733 B.n94 163.367
R684 B.n729 B.n727 163.367
R685 B.n725 B.n96 163.367
R686 B.n721 B.n719 163.367
R687 B.n717 B.n98 163.367
R688 B.n713 B.n711 163.367
R689 B.n709 B.n100 163.367
R690 B.n705 B.n703 163.367
R691 B.n701 B.n102 163.367
R692 B.n697 B.n695 163.367
R693 B.n693 B.n104 163.367
R694 B.n689 B.n687 163.367
R695 B.n685 B.n106 163.367
R696 B.n681 B.n679 163.367
R697 B.n677 B.n108 163.367
R698 B.n673 B.n671 163.367
R699 B.n669 B.n110 163.367
R700 B.n665 B.n663 163.367
R701 B.n661 B.n112 163.367
R702 B.n657 B.n655 163.367
R703 B.n653 B.n114 163.367
R704 B.n649 B.n647 163.367
R705 B.n645 B.n116 163.367
R706 B.n641 B.n639 163.367
R707 B.n637 B.n118 163.367
R708 B.n633 B.n631 163.367
R709 B.n629 B.n120 163.367
R710 B.n625 B.n623 163.367
R711 B.n621 B.n122 163.367
R712 B.n507 B.n169 163.367
R713 B.n511 B.n169 163.367
R714 B.n511 B.n163 163.367
R715 B.n519 B.n163 163.367
R716 B.n519 B.n161 163.367
R717 B.n523 B.n161 163.367
R718 B.n523 B.n155 163.367
R719 B.n531 B.n155 163.367
R720 B.n531 B.n153 163.367
R721 B.n535 B.n153 163.367
R722 B.n535 B.n147 163.367
R723 B.n543 B.n147 163.367
R724 B.n543 B.n145 163.367
R725 B.n547 B.n145 163.367
R726 B.n547 B.n140 163.367
R727 B.n556 B.n140 163.367
R728 B.n556 B.n138 163.367
R729 B.n560 B.n138 163.367
R730 B.n560 B.n131 163.367
R731 B.n568 B.n131 163.367
R732 B.n568 B.n129 163.367
R733 B.n573 B.n129 163.367
R734 B.n573 B.n124 163.367
R735 B.n581 B.n124 163.367
R736 B.n582 B.n581 163.367
R737 B.n582 B.n5 163.367
R738 B.n6 B.n5 163.367
R739 B.n7 B.n6 163.367
R740 B.n588 B.n7 163.367
R741 B.n589 B.n588 163.367
R742 B.n589 B.n13 163.367
R743 B.n14 B.n13 163.367
R744 B.n15 B.n14 163.367
R745 B.n594 B.n15 163.367
R746 B.n594 B.n20 163.367
R747 B.n21 B.n20 163.367
R748 B.n22 B.n21 163.367
R749 B.n599 B.n22 163.367
R750 B.n599 B.n27 163.367
R751 B.n28 B.n27 163.367
R752 B.n29 B.n28 163.367
R753 B.n604 B.n29 163.367
R754 B.n604 B.n34 163.367
R755 B.n35 B.n34 163.367
R756 B.n36 B.n35 163.367
R757 B.n609 B.n36 163.367
R758 B.n609 B.n41 163.367
R759 B.n42 B.n41 163.367
R760 B.n43 B.n42 163.367
R761 B.n614 B.n43 163.367
R762 B.n614 B.n48 163.367
R763 B.n49 B.n48 163.367
R764 B.n50 B.n49 163.367
R765 B.n501 B.n499 163.367
R766 B.n499 B.n498 163.367
R767 B.n495 B.n494 163.367
R768 B.n492 B.n177 163.367
R769 B.n488 B.n486 163.367
R770 B.n484 B.n179 163.367
R771 B.n480 B.n478 163.367
R772 B.n476 B.n181 163.367
R773 B.n472 B.n470 163.367
R774 B.n468 B.n183 163.367
R775 B.n464 B.n462 163.367
R776 B.n460 B.n185 163.367
R777 B.n456 B.n454 163.367
R778 B.n452 B.n187 163.367
R779 B.n448 B.n446 163.367
R780 B.n444 B.n189 163.367
R781 B.n440 B.n438 163.367
R782 B.n436 B.n191 163.367
R783 B.n432 B.n430 163.367
R784 B.n428 B.n193 163.367
R785 B.n424 B.n422 163.367
R786 B.n420 B.n195 163.367
R787 B.n416 B.n414 163.367
R788 B.n412 B.n197 163.367
R789 B.n408 B.n406 163.367
R790 B.n404 B.n199 163.367
R791 B.n400 B.n398 163.367
R792 B.n396 B.n201 163.367
R793 B.n392 B.n390 163.367
R794 B.n388 B.n203 163.367
R795 B.n384 B.n382 163.367
R796 B.n379 B.n378 163.367
R797 B.n376 B.n209 163.367
R798 B.n372 B.n370 163.367
R799 B.n368 B.n211 163.367
R800 B.n363 B.n361 163.367
R801 B.n359 B.n215 163.367
R802 B.n355 B.n353 163.367
R803 B.n351 B.n217 163.367
R804 B.n347 B.n345 163.367
R805 B.n343 B.n219 163.367
R806 B.n339 B.n337 163.367
R807 B.n335 B.n221 163.367
R808 B.n331 B.n329 163.367
R809 B.n327 B.n223 163.367
R810 B.n323 B.n321 163.367
R811 B.n319 B.n225 163.367
R812 B.n315 B.n313 163.367
R813 B.n311 B.n227 163.367
R814 B.n307 B.n305 163.367
R815 B.n303 B.n229 163.367
R816 B.n299 B.n297 163.367
R817 B.n295 B.n231 163.367
R818 B.n291 B.n289 163.367
R819 B.n287 B.n233 163.367
R820 B.n283 B.n281 163.367
R821 B.n279 B.n235 163.367
R822 B.n275 B.n273 163.367
R823 B.n271 B.n237 163.367
R824 B.n267 B.n265 163.367
R825 B.n263 B.n239 163.367
R826 B.n259 B.n257 163.367
R827 B.n255 B.n241 163.367
R828 B.n251 B.n249 163.367
R829 B.n247 B.n244 163.367
R830 B.n505 B.n167 163.367
R831 B.n513 B.n167 163.367
R832 B.n513 B.n165 163.367
R833 B.n517 B.n165 163.367
R834 B.n517 B.n159 163.367
R835 B.n525 B.n159 163.367
R836 B.n525 B.n157 163.367
R837 B.n529 B.n157 163.367
R838 B.n529 B.n151 163.367
R839 B.n537 B.n151 163.367
R840 B.n537 B.n149 163.367
R841 B.n541 B.n149 163.367
R842 B.n541 B.n143 163.367
R843 B.n550 B.n143 163.367
R844 B.n550 B.n141 163.367
R845 B.n554 B.n141 163.367
R846 B.n554 B.n136 163.367
R847 B.n562 B.n136 163.367
R848 B.n562 B.n134 163.367
R849 B.n566 B.n134 163.367
R850 B.n566 B.n128 163.367
R851 B.n575 B.n128 163.367
R852 B.n575 B.n126 163.367
R853 B.n579 B.n126 163.367
R854 B.n579 B.n3 163.367
R855 B.n935 B.n3 163.367
R856 B.n931 B.n2 163.367
R857 B.n931 B.n930 163.367
R858 B.n930 B.n9 163.367
R859 B.n926 B.n9 163.367
R860 B.n926 B.n11 163.367
R861 B.n922 B.n11 163.367
R862 B.n922 B.n17 163.367
R863 B.n918 B.n17 163.367
R864 B.n918 B.n19 163.367
R865 B.n914 B.n19 163.367
R866 B.n914 B.n23 163.367
R867 B.n910 B.n23 163.367
R868 B.n910 B.n25 163.367
R869 B.n906 B.n25 163.367
R870 B.n906 B.n31 163.367
R871 B.n902 B.n31 163.367
R872 B.n902 B.n33 163.367
R873 B.n898 B.n33 163.367
R874 B.n898 B.n38 163.367
R875 B.n894 B.n38 163.367
R876 B.n894 B.n40 163.367
R877 B.n890 B.n40 163.367
R878 B.n890 B.n45 163.367
R879 B.n886 B.n45 163.367
R880 B.n886 B.n47 163.367
R881 B.n882 B.n47 163.367
R882 B.n89 B.t10 109.889
R883 B.n212 B.t14 109.889
R884 B.n83 B.t16 109.865
R885 B.n204 B.t7 109.865
R886 B.n877 B.n52 71.676
R887 B.n876 B.n875 71.676
R888 B.n869 B.n54 71.676
R889 B.n868 B.n867 71.676
R890 B.n861 B.n56 71.676
R891 B.n860 B.n859 71.676
R892 B.n853 B.n58 71.676
R893 B.n852 B.n851 71.676
R894 B.n845 B.n60 71.676
R895 B.n844 B.n843 71.676
R896 B.n837 B.n62 71.676
R897 B.n836 B.n835 71.676
R898 B.n829 B.n64 71.676
R899 B.n828 B.n827 71.676
R900 B.n821 B.n66 71.676
R901 B.n820 B.n819 71.676
R902 B.n813 B.n68 71.676
R903 B.n812 B.n811 71.676
R904 B.n805 B.n70 71.676
R905 B.n804 B.n803 71.676
R906 B.n797 B.n72 71.676
R907 B.n796 B.n795 71.676
R908 B.n789 B.n74 71.676
R909 B.n788 B.n787 71.676
R910 B.n781 B.n76 71.676
R911 B.n780 B.n779 71.676
R912 B.n773 B.n78 71.676
R913 B.n772 B.n771 71.676
R914 B.n765 B.n80 71.676
R915 B.n764 B.n763 71.676
R916 B.n756 B.n82 71.676
R917 B.n755 B.n754 71.676
R918 B.n748 B.n86 71.676
R919 B.n747 B.n746 71.676
R920 B.n740 B.n88 71.676
R921 B.n739 B.n92 71.676
R922 B.n735 B.n734 71.676
R923 B.n728 B.n94 71.676
R924 B.n727 B.n726 71.676
R925 B.n720 B.n96 71.676
R926 B.n719 B.n718 71.676
R927 B.n712 B.n98 71.676
R928 B.n711 B.n710 71.676
R929 B.n704 B.n100 71.676
R930 B.n703 B.n702 71.676
R931 B.n696 B.n102 71.676
R932 B.n695 B.n694 71.676
R933 B.n688 B.n104 71.676
R934 B.n687 B.n686 71.676
R935 B.n680 B.n106 71.676
R936 B.n679 B.n678 71.676
R937 B.n672 B.n108 71.676
R938 B.n671 B.n670 71.676
R939 B.n664 B.n110 71.676
R940 B.n663 B.n662 71.676
R941 B.n656 B.n112 71.676
R942 B.n655 B.n654 71.676
R943 B.n648 B.n114 71.676
R944 B.n647 B.n646 71.676
R945 B.n640 B.n116 71.676
R946 B.n639 B.n638 71.676
R947 B.n632 B.n118 71.676
R948 B.n631 B.n630 71.676
R949 B.n624 B.n120 71.676
R950 B.n623 B.n622 71.676
R951 B.n622 B.n621 71.676
R952 B.n625 B.n624 71.676
R953 B.n630 B.n629 71.676
R954 B.n633 B.n632 71.676
R955 B.n638 B.n637 71.676
R956 B.n641 B.n640 71.676
R957 B.n646 B.n645 71.676
R958 B.n649 B.n648 71.676
R959 B.n654 B.n653 71.676
R960 B.n657 B.n656 71.676
R961 B.n662 B.n661 71.676
R962 B.n665 B.n664 71.676
R963 B.n670 B.n669 71.676
R964 B.n673 B.n672 71.676
R965 B.n678 B.n677 71.676
R966 B.n681 B.n680 71.676
R967 B.n686 B.n685 71.676
R968 B.n689 B.n688 71.676
R969 B.n694 B.n693 71.676
R970 B.n697 B.n696 71.676
R971 B.n702 B.n701 71.676
R972 B.n705 B.n704 71.676
R973 B.n710 B.n709 71.676
R974 B.n713 B.n712 71.676
R975 B.n718 B.n717 71.676
R976 B.n721 B.n720 71.676
R977 B.n726 B.n725 71.676
R978 B.n729 B.n728 71.676
R979 B.n734 B.n733 71.676
R980 B.n736 B.n92 71.676
R981 B.n741 B.n740 71.676
R982 B.n746 B.n745 71.676
R983 B.n749 B.n748 71.676
R984 B.n754 B.n753 71.676
R985 B.n757 B.n756 71.676
R986 B.n763 B.n762 71.676
R987 B.n766 B.n765 71.676
R988 B.n771 B.n770 71.676
R989 B.n774 B.n773 71.676
R990 B.n779 B.n778 71.676
R991 B.n782 B.n781 71.676
R992 B.n787 B.n786 71.676
R993 B.n790 B.n789 71.676
R994 B.n795 B.n794 71.676
R995 B.n798 B.n797 71.676
R996 B.n803 B.n802 71.676
R997 B.n806 B.n805 71.676
R998 B.n811 B.n810 71.676
R999 B.n814 B.n813 71.676
R1000 B.n819 B.n818 71.676
R1001 B.n822 B.n821 71.676
R1002 B.n827 B.n826 71.676
R1003 B.n830 B.n829 71.676
R1004 B.n835 B.n834 71.676
R1005 B.n838 B.n837 71.676
R1006 B.n843 B.n842 71.676
R1007 B.n846 B.n845 71.676
R1008 B.n851 B.n850 71.676
R1009 B.n854 B.n853 71.676
R1010 B.n859 B.n858 71.676
R1011 B.n862 B.n861 71.676
R1012 B.n867 B.n866 71.676
R1013 B.n870 B.n869 71.676
R1014 B.n875 B.n874 71.676
R1015 B.n878 B.n877 71.676
R1016 B.n500 B.n173 71.676
R1017 B.n498 B.n175 71.676
R1018 B.n494 B.n493 71.676
R1019 B.n487 B.n177 71.676
R1020 B.n486 B.n485 71.676
R1021 B.n479 B.n179 71.676
R1022 B.n478 B.n477 71.676
R1023 B.n471 B.n181 71.676
R1024 B.n470 B.n469 71.676
R1025 B.n463 B.n183 71.676
R1026 B.n462 B.n461 71.676
R1027 B.n455 B.n185 71.676
R1028 B.n454 B.n453 71.676
R1029 B.n447 B.n187 71.676
R1030 B.n446 B.n445 71.676
R1031 B.n439 B.n189 71.676
R1032 B.n438 B.n437 71.676
R1033 B.n431 B.n191 71.676
R1034 B.n430 B.n429 71.676
R1035 B.n423 B.n193 71.676
R1036 B.n422 B.n421 71.676
R1037 B.n415 B.n195 71.676
R1038 B.n414 B.n413 71.676
R1039 B.n407 B.n197 71.676
R1040 B.n406 B.n405 71.676
R1041 B.n399 B.n199 71.676
R1042 B.n398 B.n397 71.676
R1043 B.n391 B.n201 71.676
R1044 B.n390 B.n389 71.676
R1045 B.n383 B.n203 71.676
R1046 B.n382 B.n207 71.676
R1047 B.n378 B.n377 71.676
R1048 B.n371 B.n209 71.676
R1049 B.n370 B.n369 71.676
R1050 B.n362 B.n211 71.676
R1051 B.n361 B.n360 71.676
R1052 B.n354 B.n215 71.676
R1053 B.n353 B.n352 71.676
R1054 B.n346 B.n217 71.676
R1055 B.n345 B.n344 71.676
R1056 B.n338 B.n219 71.676
R1057 B.n337 B.n336 71.676
R1058 B.n330 B.n221 71.676
R1059 B.n329 B.n328 71.676
R1060 B.n322 B.n223 71.676
R1061 B.n321 B.n320 71.676
R1062 B.n314 B.n225 71.676
R1063 B.n313 B.n312 71.676
R1064 B.n306 B.n227 71.676
R1065 B.n305 B.n304 71.676
R1066 B.n298 B.n229 71.676
R1067 B.n297 B.n296 71.676
R1068 B.n290 B.n231 71.676
R1069 B.n289 B.n288 71.676
R1070 B.n282 B.n233 71.676
R1071 B.n281 B.n280 71.676
R1072 B.n274 B.n235 71.676
R1073 B.n273 B.n272 71.676
R1074 B.n266 B.n237 71.676
R1075 B.n265 B.n264 71.676
R1076 B.n258 B.n239 71.676
R1077 B.n257 B.n256 71.676
R1078 B.n250 B.n241 71.676
R1079 B.n249 B.n248 71.676
R1080 B.n244 B.n243 71.676
R1081 B.n501 B.n500 71.676
R1082 B.n495 B.n175 71.676
R1083 B.n493 B.n492 71.676
R1084 B.n488 B.n487 71.676
R1085 B.n485 B.n484 71.676
R1086 B.n480 B.n479 71.676
R1087 B.n477 B.n476 71.676
R1088 B.n472 B.n471 71.676
R1089 B.n469 B.n468 71.676
R1090 B.n464 B.n463 71.676
R1091 B.n461 B.n460 71.676
R1092 B.n456 B.n455 71.676
R1093 B.n453 B.n452 71.676
R1094 B.n448 B.n447 71.676
R1095 B.n445 B.n444 71.676
R1096 B.n440 B.n439 71.676
R1097 B.n437 B.n436 71.676
R1098 B.n432 B.n431 71.676
R1099 B.n429 B.n428 71.676
R1100 B.n424 B.n423 71.676
R1101 B.n421 B.n420 71.676
R1102 B.n416 B.n415 71.676
R1103 B.n413 B.n412 71.676
R1104 B.n408 B.n407 71.676
R1105 B.n405 B.n404 71.676
R1106 B.n400 B.n399 71.676
R1107 B.n397 B.n396 71.676
R1108 B.n392 B.n391 71.676
R1109 B.n389 B.n388 71.676
R1110 B.n384 B.n383 71.676
R1111 B.n379 B.n207 71.676
R1112 B.n377 B.n376 71.676
R1113 B.n372 B.n371 71.676
R1114 B.n369 B.n368 71.676
R1115 B.n363 B.n362 71.676
R1116 B.n360 B.n359 71.676
R1117 B.n355 B.n354 71.676
R1118 B.n352 B.n351 71.676
R1119 B.n347 B.n346 71.676
R1120 B.n344 B.n343 71.676
R1121 B.n339 B.n338 71.676
R1122 B.n336 B.n335 71.676
R1123 B.n331 B.n330 71.676
R1124 B.n328 B.n327 71.676
R1125 B.n323 B.n322 71.676
R1126 B.n320 B.n319 71.676
R1127 B.n315 B.n314 71.676
R1128 B.n312 B.n311 71.676
R1129 B.n307 B.n306 71.676
R1130 B.n304 B.n303 71.676
R1131 B.n299 B.n298 71.676
R1132 B.n296 B.n295 71.676
R1133 B.n291 B.n290 71.676
R1134 B.n288 B.n287 71.676
R1135 B.n283 B.n282 71.676
R1136 B.n280 B.n279 71.676
R1137 B.n275 B.n274 71.676
R1138 B.n272 B.n271 71.676
R1139 B.n267 B.n266 71.676
R1140 B.n264 B.n263 71.676
R1141 B.n259 B.n258 71.676
R1142 B.n256 B.n255 71.676
R1143 B.n251 B.n250 71.676
R1144 B.n248 B.n247 71.676
R1145 B.n243 B.n171 71.676
R1146 B.n936 B.n935 71.676
R1147 B.n936 B.n2 71.676
R1148 B.n90 B.t11 68.968
R1149 B.n213 B.t13 68.968
R1150 B.n84 B.t17 68.9433
R1151 B.n205 B.t6 68.9433
R1152 B.n506 B.n172 64.4473
R1153 B.n883 B.n51 64.4473
R1154 B.n759 B.n84 59.5399
R1155 B.n91 B.n90 59.5399
R1156 B.n365 B.n213 59.5399
R1157 B.n206 B.n205 59.5399
R1158 B.n84 B.n83 40.9217
R1159 B.n90 B.n89 40.9217
R1160 B.n213 B.n212 40.9217
R1161 B.n205 B.n204 40.9217
R1162 B.n504 B.n503 33.5615
R1163 B.n508 B.n170 33.5615
R1164 B.n619 B.n618 33.5615
R1165 B.n881 B.n880 33.5615
R1166 B.n506 B.n168 31.5284
R1167 B.n512 B.n168 31.5284
R1168 B.n512 B.n164 31.5284
R1169 B.n518 B.n164 31.5284
R1170 B.n518 B.n160 31.5284
R1171 B.n524 B.n160 31.5284
R1172 B.n530 B.n156 31.5284
R1173 B.n530 B.n152 31.5284
R1174 B.n536 B.n152 31.5284
R1175 B.n536 B.n148 31.5284
R1176 B.n542 B.n148 31.5284
R1177 B.n542 B.n144 31.5284
R1178 B.n549 B.n144 31.5284
R1179 B.n549 B.n548 31.5284
R1180 B.n555 B.n137 31.5284
R1181 B.n561 B.n137 31.5284
R1182 B.n561 B.n132 31.5284
R1183 B.n567 B.n132 31.5284
R1184 B.n567 B.n133 31.5284
R1185 B.n574 B.n125 31.5284
R1186 B.n580 B.n125 31.5284
R1187 B.n580 B.n4 31.5284
R1188 B.n934 B.n4 31.5284
R1189 B.n934 B.n933 31.5284
R1190 B.n933 B.n932 31.5284
R1191 B.n932 B.n8 31.5284
R1192 B.n12 B.n8 31.5284
R1193 B.n925 B.n12 31.5284
R1194 B.n924 B.n923 31.5284
R1195 B.n923 B.n16 31.5284
R1196 B.n917 B.n16 31.5284
R1197 B.n917 B.n916 31.5284
R1198 B.n916 B.n915 31.5284
R1199 B.n909 B.n26 31.5284
R1200 B.n909 B.n908 31.5284
R1201 B.n908 B.n907 31.5284
R1202 B.n907 B.n30 31.5284
R1203 B.n901 B.n30 31.5284
R1204 B.n901 B.n900 31.5284
R1205 B.n900 B.n899 31.5284
R1206 B.n899 B.n37 31.5284
R1207 B.n893 B.n892 31.5284
R1208 B.n892 B.n891 31.5284
R1209 B.n891 B.n44 31.5284
R1210 B.n885 B.n44 31.5284
R1211 B.n885 B.n884 31.5284
R1212 B.n884 B.n883 31.5284
R1213 B.t5 B.n156 25.9647
R1214 B.t9 B.n37 25.9647
R1215 B.n133 B.t0 25.0374
R1216 B.t3 B.n924 25.0374
R1217 B.n548 B.t1 18.5463
R1218 B.n26 B.t2 18.5463
R1219 B B.n937 18.0485
R1220 B.n555 B.t1 12.9826
R1221 B.n915 B.t2 12.9826
R1222 B.n504 B.n166 10.6151
R1223 B.n514 B.n166 10.6151
R1224 B.n515 B.n514 10.6151
R1225 B.n516 B.n515 10.6151
R1226 B.n516 B.n158 10.6151
R1227 B.n526 B.n158 10.6151
R1228 B.n527 B.n526 10.6151
R1229 B.n528 B.n527 10.6151
R1230 B.n528 B.n150 10.6151
R1231 B.n538 B.n150 10.6151
R1232 B.n539 B.n538 10.6151
R1233 B.n540 B.n539 10.6151
R1234 B.n540 B.n142 10.6151
R1235 B.n551 B.n142 10.6151
R1236 B.n552 B.n551 10.6151
R1237 B.n553 B.n552 10.6151
R1238 B.n553 B.n135 10.6151
R1239 B.n563 B.n135 10.6151
R1240 B.n564 B.n563 10.6151
R1241 B.n565 B.n564 10.6151
R1242 B.n565 B.n127 10.6151
R1243 B.n576 B.n127 10.6151
R1244 B.n577 B.n576 10.6151
R1245 B.n578 B.n577 10.6151
R1246 B.n578 B.n0 10.6151
R1247 B.n503 B.n502 10.6151
R1248 B.n502 B.n174 10.6151
R1249 B.n497 B.n174 10.6151
R1250 B.n497 B.n496 10.6151
R1251 B.n496 B.n176 10.6151
R1252 B.n491 B.n176 10.6151
R1253 B.n491 B.n490 10.6151
R1254 B.n490 B.n489 10.6151
R1255 B.n489 B.n178 10.6151
R1256 B.n483 B.n178 10.6151
R1257 B.n483 B.n482 10.6151
R1258 B.n482 B.n481 10.6151
R1259 B.n481 B.n180 10.6151
R1260 B.n475 B.n180 10.6151
R1261 B.n475 B.n474 10.6151
R1262 B.n474 B.n473 10.6151
R1263 B.n473 B.n182 10.6151
R1264 B.n467 B.n182 10.6151
R1265 B.n467 B.n466 10.6151
R1266 B.n466 B.n465 10.6151
R1267 B.n465 B.n184 10.6151
R1268 B.n459 B.n184 10.6151
R1269 B.n459 B.n458 10.6151
R1270 B.n458 B.n457 10.6151
R1271 B.n457 B.n186 10.6151
R1272 B.n451 B.n186 10.6151
R1273 B.n451 B.n450 10.6151
R1274 B.n450 B.n449 10.6151
R1275 B.n449 B.n188 10.6151
R1276 B.n443 B.n188 10.6151
R1277 B.n443 B.n442 10.6151
R1278 B.n442 B.n441 10.6151
R1279 B.n441 B.n190 10.6151
R1280 B.n435 B.n190 10.6151
R1281 B.n435 B.n434 10.6151
R1282 B.n434 B.n433 10.6151
R1283 B.n433 B.n192 10.6151
R1284 B.n427 B.n192 10.6151
R1285 B.n427 B.n426 10.6151
R1286 B.n426 B.n425 10.6151
R1287 B.n425 B.n194 10.6151
R1288 B.n419 B.n194 10.6151
R1289 B.n419 B.n418 10.6151
R1290 B.n418 B.n417 10.6151
R1291 B.n417 B.n196 10.6151
R1292 B.n411 B.n196 10.6151
R1293 B.n411 B.n410 10.6151
R1294 B.n410 B.n409 10.6151
R1295 B.n409 B.n198 10.6151
R1296 B.n403 B.n198 10.6151
R1297 B.n403 B.n402 10.6151
R1298 B.n402 B.n401 10.6151
R1299 B.n401 B.n200 10.6151
R1300 B.n395 B.n200 10.6151
R1301 B.n395 B.n394 10.6151
R1302 B.n394 B.n393 10.6151
R1303 B.n393 B.n202 10.6151
R1304 B.n387 B.n202 10.6151
R1305 B.n387 B.n386 10.6151
R1306 B.n386 B.n385 10.6151
R1307 B.n381 B.n380 10.6151
R1308 B.n380 B.n208 10.6151
R1309 B.n375 B.n208 10.6151
R1310 B.n375 B.n374 10.6151
R1311 B.n374 B.n373 10.6151
R1312 B.n373 B.n210 10.6151
R1313 B.n367 B.n210 10.6151
R1314 B.n367 B.n366 10.6151
R1315 B.n364 B.n214 10.6151
R1316 B.n358 B.n214 10.6151
R1317 B.n358 B.n357 10.6151
R1318 B.n357 B.n356 10.6151
R1319 B.n356 B.n216 10.6151
R1320 B.n350 B.n216 10.6151
R1321 B.n350 B.n349 10.6151
R1322 B.n349 B.n348 10.6151
R1323 B.n348 B.n218 10.6151
R1324 B.n342 B.n218 10.6151
R1325 B.n342 B.n341 10.6151
R1326 B.n341 B.n340 10.6151
R1327 B.n340 B.n220 10.6151
R1328 B.n334 B.n220 10.6151
R1329 B.n334 B.n333 10.6151
R1330 B.n333 B.n332 10.6151
R1331 B.n332 B.n222 10.6151
R1332 B.n326 B.n222 10.6151
R1333 B.n326 B.n325 10.6151
R1334 B.n325 B.n324 10.6151
R1335 B.n324 B.n224 10.6151
R1336 B.n318 B.n224 10.6151
R1337 B.n318 B.n317 10.6151
R1338 B.n317 B.n316 10.6151
R1339 B.n316 B.n226 10.6151
R1340 B.n310 B.n226 10.6151
R1341 B.n310 B.n309 10.6151
R1342 B.n309 B.n308 10.6151
R1343 B.n308 B.n228 10.6151
R1344 B.n302 B.n228 10.6151
R1345 B.n302 B.n301 10.6151
R1346 B.n301 B.n300 10.6151
R1347 B.n300 B.n230 10.6151
R1348 B.n294 B.n230 10.6151
R1349 B.n294 B.n293 10.6151
R1350 B.n293 B.n292 10.6151
R1351 B.n292 B.n232 10.6151
R1352 B.n286 B.n232 10.6151
R1353 B.n286 B.n285 10.6151
R1354 B.n285 B.n284 10.6151
R1355 B.n284 B.n234 10.6151
R1356 B.n278 B.n234 10.6151
R1357 B.n278 B.n277 10.6151
R1358 B.n277 B.n276 10.6151
R1359 B.n276 B.n236 10.6151
R1360 B.n270 B.n236 10.6151
R1361 B.n270 B.n269 10.6151
R1362 B.n269 B.n268 10.6151
R1363 B.n268 B.n238 10.6151
R1364 B.n262 B.n238 10.6151
R1365 B.n262 B.n261 10.6151
R1366 B.n261 B.n260 10.6151
R1367 B.n260 B.n240 10.6151
R1368 B.n254 B.n240 10.6151
R1369 B.n254 B.n253 10.6151
R1370 B.n253 B.n252 10.6151
R1371 B.n252 B.n242 10.6151
R1372 B.n246 B.n242 10.6151
R1373 B.n246 B.n245 10.6151
R1374 B.n245 B.n170 10.6151
R1375 B.n509 B.n508 10.6151
R1376 B.n510 B.n509 10.6151
R1377 B.n510 B.n162 10.6151
R1378 B.n520 B.n162 10.6151
R1379 B.n521 B.n520 10.6151
R1380 B.n522 B.n521 10.6151
R1381 B.n522 B.n154 10.6151
R1382 B.n532 B.n154 10.6151
R1383 B.n533 B.n532 10.6151
R1384 B.n534 B.n533 10.6151
R1385 B.n534 B.n146 10.6151
R1386 B.n544 B.n146 10.6151
R1387 B.n545 B.n544 10.6151
R1388 B.n546 B.n545 10.6151
R1389 B.n546 B.n139 10.6151
R1390 B.n557 B.n139 10.6151
R1391 B.n558 B.n557 10.6151
R1392 B.n559 B.n558 10.6151
R1393 B.n559 B.n130 10.6151
R1394 B.n569 B.n130 10.6151
R1395 B.n570 B.n569 10.6151
R1396 B.n572 B.n570 10.6151
R1397 B.n572 B.n571 10.6151
R1398 B.n571 B.n123 10.6151
R1399 B.n583 B.n123 10.6151
R1400 B.n584 B.n583 10.6151
R1401 B.n585 B.n584 10.6151
R1402 B.n586 B.n585 10.6151
R1403 B.n587 B.n586 10.6151
R1404 B.n590 B.n587 10.6151
R1405 B.n591 B.n590 10.6151
R1406 B.n592 B.n591 10.6151
R1407 B.n593 B.n592 10.6151
R1408 B.n595 B.n593 10.6151
R1409 B.n596 B.n595 10.6151
R1410 B.n597 B.n596 10.6151
R1411 B.n598 B.n597 10.6151
R1412 B.n600 B.n598 10.6151
R1413 B.n601 B.n600 10.6151
R1414 B.n602 B.n601 10.6151
R1415 B.n603 B.n602 10.6151
R1416 B.n605 B.n603 10.6151
R1417 B.n606 B.n605 10.6151
R1418 B.n607 B.n606 10.6151
R1419 B.n608 B.n607 10.6151
R1420 B.n610 B.n608 10.6151
R1421 B.n611 B.n610 10.6151
R1422 B.n612 B.n611 10.6151
R1423 B.n613 B.n612 10.6151
R1424 B.n615 B.n613 10.6151
R1425 B.n616 B.n615 10.6151
R1426 B.n617 B.n616 10.6151
R1427 B.n618 B.n617 10.6151
R1428 B.n929 B.n1 10.6151
R1429 B.n929 B.n928 10.6151
R1430 B.n928 B.n927 10.6151
R1431 B.n927 B.n10 10.6151
R1432 B.n921 B.n10 10.6151
R1433 B.n921 B.n920 10.6151
R1434 B.n920 B.n919 10.6151
R1435 B.n919 B.n18 10.6151
R1436 B.n913 B.n18 10.6151
R1437 B.n913 B.n912 10.6151
R1438 B.n912 B.n911 10.6151
R1439 B.n911 B.n24 10.6151
R1440 B.n905 B.n24 10.6151
R1441 B.n905 B.n904 10.6151
R1442 B.n904 B.n903 10.6151
R1443 B.n903 B.n32 10.6151
R1444 B.n897 B.n32 10.6151
R1445 B.n897 B.n896 10.6151
R1446 B.n896 B.n895 10.6151
R1447 B.n895 B.n39 10.6151
R1448 B.n889 B.n39 10.6151
R1449 B.n889 B.n888 10.6151
R1450 B.n888 B.n887 10.6151
R1451 B.n887 B.n46 10.6151
R1452 B.n881 B.n46 10.6151
R1453 B.n880 B.n879 10.6151
R1454 B.n879 B.n53 10.6151
R1455 B.n873 B.n53 10.6151
R1456 B.n873 B.n872 10.6151
R1457 B.n872 B.n871 10.6151
R1458 B.n871 B.n55 10.6151
R1459 B.n865 B.n55 10.6151
R1460 B.n865 B.n864 10.6151
R1461 B.n864 B.n863 10.6151
R1462 B.n863 B.n57 10.6151
R1463 B.n857 B.n57 10.6151
R1464 B.n857 B.n856 10.6151
R1465 B.n856 B.n855 10.6151
R1466 B.n855 B.n59 10.6151
R1467 B.n849 B.n59 10.6151
R1468 B.n849 B.n848 10.6151
R1469 B.n848 B.n847 10.6151
R1470 B.n847 B.n61 10.6151
R1471 B.n841 B.n61 10.6151
R1472 B.n841 B.n840 10.6151
R1473 B.n840 B.n839 10.6151
R1474 B.n839 B.n63 10.6151
R1475 B.n833 B.n63 10.6151
R1476 B.n833 B.n832 10.6151
R1477 B.n832 B.n831 10.6151
R1478 B.n831 B.n65 10.6151
R1479 B.n825 B.n65 10.6151
R1480 B.n825 B.n824 10.6151
R1481 B.n824 B.n823 10.6151
R1482 B.n823 B.n67 10.6151
R1483 B.n817 B.n67 10.6151
R1484 B.n817 B.n816 10.6151
R1485 B.n816 B.n815 10.6151
R1486 B.n815 B.n69 10.6151
R1487 B.n809 B.n69 10.6151
R1488 B.n809 B.n808 10.6151
R1489 B.n808 B.n807 10.6151
R1490 B.n807 B.n71 10.6151
R1491 B.n801 B.n71 10.6151
R1492 B.n801 B.n800 10.6151
R1493 B.n800 B.n799 10.6151
R1494 B.n799 B.n73 10.6151
R1495 B.n793 B.n73 10.6151
R1496 B.n793 B.n792 10.6151
R1497 B.n792 B.n791 10.6151
R1498 B.n791 B.n75 10.6151
R1499 B.n785 B.n75 10.6151
R1500 B.n785 B.n784 10.6151
R1501 B.n784 B.n783 10.6151
R1502 B.n783 B.n77 10.6151
R1503 B.n777 B.n77 10.6151
R1504 B.n777 B.n776 10.6151
R1505 B.n776 B.n775 10.6151
R1506 B.n775 B.n79 10.6151
R1507 B.n769 B.n79 10.6151
R1508 B.n769 B.n768 10.6151
R1509 B.n768 B.n767 10.6151
R1510 B.n767 B.n81 10.6151
R1511 B.n761 B.n81 10.6151
R1512 B.n761 B.n760 10.6151
R1513 B.n758 B.n85 10.6151
R1514 B.n752 B.n85 10.6151
R1515 B.n752 B.n751 10.6151
R1516 B.n751 B.n750 10.6151
R1517 B.n750 B.n87 10.6151
R1518 B.n744 B.n87 10.6151
R1519 B.n744 B.n743 10.6151
R1520 B.n743 B.n742 10.6151
R1521 B.n738 B.n737 10.6151
R1522 B.n737 B.n93 10.6151
R1523 B.n732 B.n93 10.6151
R1524 B.n732 B.n731 10.6151
R1525 B.n731 B.n730 10.6151
R1526 B.n730 B.n95 10.6151
R1527 B.n724 B.n95 10.6151
R1528 B.n724 B.n723 10.6151
R1529 B.n723 B.n722 10.6151
R1530 B.n722 B.n97 10.6151
R1531 B.n716 B.n97 10.6151
R1532 B.n716 B.n715 10.6151
R1533 B.n715 B.n714 10.6151
R1534 B.n714 B.n99 10.6151
R1535 B.n708 B.n99 10.6151
R1536 B.n708 B.n707 10.6151
R1537 B.n707 B.n706 10.6151
R1538 B.n706 B.n101 10.6151
R1539 B.n700 B.n101 10.6151
R1540 B.n700 B.n699 10.6151
R1541 B.n699 B.n698 10.6151
R1542 B.n698 B.n103 10.6151
R1543 B.n692 B.n103 10.6151
R1544 B.n692 B.n691 10.6151
R1545 B.n691 B.n690 10.6151
R1546 B.n690 B.n105 10.6151
R1547 B.n684 B.n105 10.6151
R1548 B.n684 B.n683 10.6151
R1549 B.n683 B.n682 10.6151
R1550 B.n682 B.n107 10.6151
R1551 B.n676 B.n107 10.6151
R1552 B.n676 B.n675 10.6151
R1553 B.n675 B.n674 10.6151
R1554 B.n674 B.n109 10.6151
R1555 B.n668 B.n109 10.6151
R1556 B.n668 B.n667 10.6151
R1557 B.n667 B.n666 10.6151
R1558 B.n666 B.n111 10.6151
R1559 B.n660 B.n111 10.6151
R1560 B.n660 B.n659 10.6151
R1561 B.n659 B.n658 10.6151
R1562 B.n658 B.n113 10.6151
R1563 B.n652 B.n113 10.6151
R1564 B.n652 B.n651 10.6151
R1565 B.n651 B.n650 10.6151
R1566 B.n650 B.n115 10.6151
R1567 B.n644 B.n115 10.6151
R1568 B.n644 B.n643 10.6151
R1569 B.n643 B.n642 10.6151
R1570 B.n642 B.n117 10.6151
R1571 B.n636 B.n117 10.6151
R1572 B.n636 B.n635 10.6151
R1573 B.n635 B.n634 10.6151
R1574 B.n634 B.n119 10.6151
R1575 B.n628 B.n119 10.6151
R1576 B.n628 B.n627 10.6151
R1577 B.n627 B.n626 10.6151
R1578 B.n626 B.n121 10.6151
R1579 B.n620 B.n121 10.6151
R1580 B.n620 B.n619 10.6151
R1581 B.n937 B.n0 8.11757
R1582 B.n937 B.n1 8.11757
R1583 B.n381 B.n206 6.5566
R1584 B.n366 B.n365 6.5566
R1585 B.n759 B.n758 6.5566
R1586 B.n742 B.n91 6.5566
R1587 B.n574 B.t0 6.49154
R1588 B.n925 B.t3 6.49154
R1589 B.n524 B.t5 5.56425
R1590 B.n893 B.t9 5.56425
R1591 B.n385 B.n206 4.05904
R1592 B.n365 B.n364 4.05904
R1593 B.n760 B.n759 4.05904
R1594 B.n738 B.n91 4.05904
R1595 VP.n3 VP.t2 286.048
R1596 VP.n3 VP.t1 285.618
R1597 VP.n5 VP.t3 249.802
R1598 VP.n13 VP.t0 249.802
R1599 VP.n5 VP.n4 183.077
R1600 VP.n14 VP.n13 183.077
R1601 VP.n12 VP.n0 161.3
R1602 VP.n11 VP.n10 161.3
R1603 VP.n9 VP.n1 161.3
R1604 VP.n8 VP.n7 161.3
R1605 VP.n6 VP.n2 161.3
R1606 VP.n4 VP.n3 57.9441
R1607 VP.n7 VP.n1 40.4934
R1608 VP.n11 VP.n1 40.4934
R1609 VP.n7 VP.n6 24.4675
R1610 VP.n12 VP.n11 24.4675
R1611 VP.n6 VP.n5 2.69187
R1612 VP.n13 VP.n12 2.69187
R1613 VP.n4 VP.n2 0.189894
R1614 VP.n8 VP.n2 0.189894
R1615 VP.n9 VP.n8 0.189894
R1616 VP.n10 VP.n9 0.189894
R1617 VP.n10 VP.n0 0.189894
R1618 VP.n14 VP.n0 0.189894
R1619 VP VP.n14 0.0516364
R1620 VDD1 VDD1.n1 109.812
R1621 VDD1 VDD1.n0 64.2677
R1622 VDD1.n0 VDD1.t1 1.07367
R1623 VDD1.n0 VDD1.t2 1.07367
R1624 VDD1.n1 VDD1.t0 1.07367
R1625 VDD1.n1 VDD1.t3 1.07367
C0 VTAIL VDD1 7.21697f
C1 VP VN 6.79467f
C2 VP VTAIL 6.12099f
C3 VDD1 VDD2 0.826815f
C4 VN VTAIL 6.10689f
C5 VP VDD2 0.341949f
C6 VN VDD2 6.5783f
C7 VTAIL VDD2 7.26568f
C8 VP VDD1 6.77164f
C9 VN VDD1 0.14808f
C10 VDD2 B 3.804843f
C11 VDD1 B 8.359241f
C12 VTAIL B 13.386457f
C13 VN B 9.88209f
C14 VP B 7.617009f
C15 VDD1.t1 B 0.388038f
C16 VDD1.t2 B 0.388038f
C17 VDD1.n0 B 3.54941f
C18 VDD1.t0 B 0.388038f
C19 VDD1.t3 B 0.388038f
C20 VDD1.n1 B 4.41345f
C21 VP.n0 B 0.031318f
C22 VP.t0 B 2.83033f
C23 VP.n1 B 0.025318f
C24 VP.n2 B 0.031318f
C25 VP.t3 B 2.83033f
C26 VP.t2 B 2.97486f
C27 VP.t1 B 2.97314f
C28 VP.n3 B 3.59462f
C29 VP.n4 B 1.96068f
C30 VP.n5 B 1.05805f
C31 VP.n6 B 0.032721f
C32 VP.n7 B 0.062245f
C33 VP.n8 B 0.031318f
C34 VP.n9 B 0.031318f
C35 VP.n10 B 0.031318f
C36 VP.n11 B 0.062245f
C37 VP.n12 B 0.032721f
C38 VP.n13 B 1.05805f
C39 VP.n14 B 0.03351f
C40 VDD2.t1 B 0.387991f
C41 VDD2.t3 B 0.387991f
C42 VDD2.n0 B 4.38535f
C43 VDD2.t2 B 0.387991f
C44 VDD2.t0 B 0.387991f
C45 VDD2.n1 B 3.54863f
C46 VDD2.n2 B 4.25236f
C47 VTAIL.t4 B 2.51406f
C48 VTAIL.n0 B 0.261266f
C49 VTAIL.t0 B 2.51406f
C50 VTAIL.n1 B 0.302571f
C51 VTAIL.t1 B 2.51406f
C52 VTAIL.n2 B 1.3443f
C53 VTAIL.t5 B 2.51406f
C54 VTAIL.n3 B 1.34431f
C55 VTAIL.t6 B 2.51406f
C56 VTAIL.n4 B 0.302578f
C57 VTAIL.t3 B 2.51406f
C58 VTAIL.n5 B 0.302578f
C59 VTAIL.t2 B 2.51406f
C60 VTAIL.n6 B 1.34431f
C61 VTAIL.t7 B 2.51406f
C62 VTAIL.n7 B 1.29735f
C63 VN.t2 B 2.93809f
C64 VN.t0 B 2.93639f
C65 VN.n0 B 2.02626f
C66 VN.t3 B 2.93809f
C67 VN.t1 B 2.93639f
C68 VN.n1 B 3.56902f
.ends

