* NGSPICE file created from diff_pair_sample_0817.ext - technology: sky130A

.subckt diff_pair_sample_0817 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t8 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0.3729 ps=2.59 w=2.26 l=3.83
X1 VDD2.t9 VN.t0 VTAIL.t18 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0.3729 ps=2.59 w=2.26 l=3.83
X2 VDD1.t8 VP.t1 VTAIL.t16 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X3 B.t11 B.t9 B.t10 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0 ps=0 w=2.26 l=3.83
X4 VTAIL.t1 VN.t1 VDD2.t8 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X5 VTAIL.t11 VP.t2 VDD1.t7 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X6 VDD2.t7 VN.t2 VTAIL.t19 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X7 VDD2.t6 VN.t3 VTAIL.t3 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.8814 ps=5.3 w=2.26 l=3.83
X8 VDD1.t6 VP.t3 VTAIL.t7 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.8814 ps=5.3 w=2.26 l=3.83
X9 VTAIL.t4 VN.t4 VDD2.t5 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X10 VTAIL.t6 VN.t5 VDD2.t4 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X11 VTAIL.t15 VP.t4 VDD1.t5 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X12 VTAIL.t13 VP.t5 VDD1.t4 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X13 VDD2.t3 VN.t6 VTAIL.t2 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.8814 ps=5.3 w=2.26 l=3.83
X14 VDD2.t2 VN.t7 VTAIL.t17 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X15 VDD2.t1 VN.t8 VTAIL.t5 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0.3729 ps=2.59 w=2.26 l=3.83
X16 B.t8 B.t6 B.t7 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0 ps=0 w=2.26 l=3.83
X17 VTAIL.t0 VN.t9 VDD2.t0 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X18 VDD1.t3 VP.t6 VTAIL.t12 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.8814 ps=5.3 w=2.26 l=3.83
X19 VDD1.t2 VP.t7 VTAIL.t10 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X20 VTAIL.t9 VP.t8 VDD1.t1 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.3729 pd=2.59 as=0.3729 ps=2.59 w=2.26 l=3.83
X21 B.t5 B.t3 B.t4 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0 ps=0 w=2.26 l=3.83
X22 B.t2 B.t0 B.t1 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0 ps=0 w=2.26 l=3.83
X23 VDD1.t0 VP.t9 VTAIL.t14 w_n5962_n1420# sky130_fd_pr__pfet_01v8 ad=0.8814 pd=5.3 as=0.3729 ps=2.59 w=2.26 l=3.83
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n75 VP.n74 86.8027
R60 VP.n130 VP.n0 86.8027
R61 VP.n73 VP.n18 86.8027
R62 VP.n96 VP.n95 56.5617
R63 VP.n109 VP.n108 56.5617
R64 VP.n52 VP.n51 56.5617
R65 VP.n39 VP.n38 56.5617
R66 VP.n32 VP.n31 55.106
R67 VP.n74 VP.n73 52.492
R68 VP.n31 VP.t0 47.3096
R69 VP.n83 VP.n82 41.5458
R70 VP.n122 VP.n121 41.5458
R71 VP.n65 VP.n64 41.5458
R72 VP.n82 VP.n81 39.6083
R73 VP.n122 VP.n2 39.6083
R74 VP.n65 VP.n20 39.6083
R75 VP.n77 VP.n76 24.5923
R76 VP.n77 VP.n16 24.5923
R77 VP.n81 VP.n16 24.5923
R78 VP.n83 VP.n14 24.5923
R79 VP.n87 VP.n14 24.5923
R80 VP.n88 VP.n87 24.5923
R81 VP.n90 VP.n12 24.5923
R82 VP.n94 VP.n12 24.5923
R83 VP.n95 VP.n94 24.5923
R84 VP.n96 VP.n10 24.5923
R85 VP.n100 VP.n10 24.5923
R86 VP.n101 VP.n100 24.5923
R87 VP.n103 VP.n8 24.5923
R88 VP.n107 VP.n8 24.5923
R89 VP.n108 VP.n107 24.5923
R90 VP.n109 VP.n6 24.5923
R91 VP.n113 VP.n6 24.5923
R92 VP.n114 VP.n113 24.5923
R93 VP.n116 VP.n4 24.5923
R94 VP.n120 VP.n4 24.5923
R95 VP.n121 VP.n120 24.5923
R96 VP.n126 VP.n2 24.5923
R97 VP.n127 VP.n126 24.5923
R98 VP.n128 VP.n127 24.5923
R99 VP.n69 VP.n20 24.5923
R100 VP.n70 VP.n69 24.5923
R101 VP.n71 VP.n70 24.5923
R102 VP.n52 VP.n24 24.5923
R103 VP.n56 VP.n24 24.5923
R104 VP.n57 VP.n56 24.5923
R105 VP.n59 VP.n22 24.5923
R106 VP.n63 VP.n22 24.5923
R107 VP.n64 VP.n63 24.5923
R108 VP.n39 VP.n28 24.5923
R109 VP.n43 VP.n28 24.5923
R110 VP.n44 VP.n43 24.5923
R111 VP.n46 VP.n26 24.5923
R112 VP.n50 VP.n26 24.5923
R113 VP.n51 VP.n50 24.5923
R114 VP.n33 VP.n30 24.5923
R115 VP.n37 VP.n30 24.5923
R116 VP.n38 VP.n37 24.5923
R117 VP.n90 VP.n89 20.1658
R118 VP.n115 VP.n114 20.1658
R119 VP.n58 VP.n57 20.1658
R120 VP.n33 VP.n32 20.1658
R121 VP.n75 VP.t9 14.2214
R122 VP.n89 VP.t8 14.2214
R123 VP.n102 VP.t7 14.2214
R124 VP.n115 VP.t5 14.2214
R125 VP.n0 VP.t6 14.2214
R126 VP.n18 VP.t3 14.2214
R127 VP.n58 VP.t4 14.2214
R128 VP.n45 VP.t1 14.2214
R129 VP.n32 VP.t2 14.2214
R130 VP.n102 VP.n101 12.2964
R131 VP.n103 VP.n102 12.2964
R132 VP.n45 VP.n44 12.2964
R133 VP.n46 VP.n45 12.2964
R134 VP.n89 VP.n88 4.42703
R135 VP.n116 VP.n115 4.42703
R136 VP.n59 VP.n58 4.42703
R137 VP.n76 VP.n75 3.44336
R138 VP.n128 VP.n0 3.44336
R139 VP.n71 VP.n18 3.44336
R140 VP.n34 VP.n31 2.44068
R141 VP.n73 VP.n72 0.354861
R142 VP.n74 VP.n17 0.354861
R143 VP.n130 VP.n129 0.354861
R144 VP VP.n130 0.267071
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VTAIL.n17 VTAIL.t3 172.81
R203 VTAIL.n2 VTAIL.t12 172.81
R204 VTAIL.n16 VTAIL.t7 172.81
R205 VTAIL.n11 VTAIL.t2 172.81
R206 VTAIL.n15 VTAIL.n14 158.428
R207 VTAIL.n13 VTAIL.n12 158.428
R208 VTAIL.n10 VTAIL.n9 158.428
R209 VTAIL.n8 VTAIL.n7 158.428
R210 VTAIL.n19 VTAIL.n18 158.427
R211 VTAIL.n1 VTAIL.n0 158.427
R212 VTAIL.n4 VTAIL.n3 158.427
R213 VTAIL.n6 VTAIL.n5 158.427
R214 VTAIL.n8 VTAIL.n6 21.4876
R215 VTAIL.n17 VTAIL.n16 17.9014
R216 VTAIL.n18 VTAIL.t17 14.3832
R217 VTAIL.n18 VTAIL.t4 14.3832
R218 VTAIL.n0 VTAIL.t5 14.3832
R219 VTAIL.n0 VTAIL.t6 14.3832
R220 VTAIL.n3 VTAIL.t10 14.3832
R221 VTAIL.n3 VTAIL.t13 14.3832
R222 VTAIL.n5 VTAIL.t14 14.3832
R223 VTAIL.n5 VTAIL.t9 14.3832
R224 VTAIL.n14 VTAIL.t16 14.3832
R225 VTAIL.n14 VTAIL.t15 14.3832
R226 VTAIL.n12 VTAIL.t8 14.3832
R227 VTAIL.n12 VTAIL.t11 14.3832
R228 VTAIL.n9 VTAIL.t19 14.3832
R229 VTAIL.n9 VTAIL.t0 14.3832
R230 VTAIL.n7 VTAIL.t18 14.3832
R231 VTAIL.n7 VTAIL.t1 14.3832
R232 VTAIL.n10 VTAIL.n8 3.58671
R233 VTAIL.n11 VTAIL.n10 3.58671
R234 VTAIL.n15 VTAIL.n13 3.58671
R235 VTAIL.n16 VTAIL.n15 3.58671
R236 VTAIL.n6 VTAIL.n4 3.58671
R237 VTAIL.n4 VTAIL.n2 3.58671
R238 VTAIL.n19 VTAIL.n17 3.58671
R239 VTAIL VTAIL.n1 2.74834
R240 VTAIL.n13 VTAIL.n11 2.26343
R241 VTAIL.n2 VTAIL.n1 2.26343
R242 VTAIL VTAIL.n19 0.838862
R243 VDD1.n3 VDD1.t0 193.075
R244 VDD1.n1 VDD1.t9 193.075
R245 VDD1.n5 VDD1.n4 177.74
R246 VDD1.n1 VDD1.n0 175.107
R247 VDD1.n7 VDD1.n6 175.106
R248 VDD1.n3 VDD1.n2 175.106
R249 VDD1.n7 VDD1.n5 45.0742
R250 VDD1.n6 VDD1.t5 14.3832
R251 VDD1.n6 VDD1.t6 14.3832
R252 VDD1.n0 VDD1.t7 14.3832
R253 VDD1.n0 VDD1.t8 14.3832
R254 VDD1.n4 VDD1.t4 14.3832
R255 VDD1.n4 VDD1.t3 14.3832
R256 VDD1.n2 VDD1.t1 14.3832
R257 VDD1.n2 VDD1.t2 14.3832
R258 VDD1 VDD1.n7 2.63197
R259 VDD1 VDD1.n1 0.955241
R260 VDD1.n5 VDD1.n3 0.841706
R261 VN.n110 VN.n109 161.3
R262 VN.n108 VN.n57 161.3
R263 VN.n107 VN.n106 161.3
R264 VN.n105 VN.n58 161.3
R265 VN.n104 VN.n103 161.3
R266 VN.n102 VN.n59 161.3
R267 VN.n101 VN.n100 161.3
R268 VN.n99 VN.n60 161.3
R269 VN.n98 VN.n97 161.3
R270 VN.n95 VN.n61 161.3
R271 VN.n94 VN.n93 161.3
R272 VN.n92 VN.n62 161.3
R273 VN.n91 VN.n90 161.3
R274 VN.n89 VN.n63 161.3
R275 VN.n88 VN.n87 161.3
R276 VN.n86 VN.n64 161.3
R277 VN.n85 VN.n84 161.3
R278 VN.n82 VN.n65 161.3
R279 VN.n81 VN.n80 161.3
R280 VN.n79 VN.n66 161.3
R281 VN.n78 VN.n77 161.3
R282 VN.n76 VN.n67 161.3
R283 VN.n75 VN.n74 161.3
R284 VN.n73 VN.n68 161.3
R285 VN.n72 VN.n71 161.3
R286 VN.n54 VN.n53 161.3
R287 VN.n52 VN.n1 161.3
R288 VN.n51 VN.n50 161.3
R289 VN.n49 VN.n2 161.3
R290 VN.n48 VN.n47 161.3
R291 VN.n46 VN.n3 161.3
R292 VN.n45 VN.n44 161.3
R293 VN.n43 VN.n4 161.3
R294 VN.n42 VN.n41 161.3
R295 VN.n39 VN.n5 161.3
R296 VN.n38 VN.n37 161.3
R297 VN.n36 VN.n6 161.3
R298 VN.n35 VN.n34 161.3
R299 VN.n33 VN.n7 161.3
R300 VN.n32 VN.n31 161.3
R301 VN.n30 VN.n8 161.3
R302 VN.n29 VN.n28 161.3
R303 VN.n26 VN.n9 161.3
R304 VN.n25 VN.n24 161.3
R305 VN.n23 VN.n10 161.3
R306 VN.n22 VN.n21 161.3
R307 VN.n20 VN.n11 161.3
R308 VN.n19 VN.n18 161.3
R309 VN.n17 VN.n12 161.3
R310 VN.n16 VN.n15 161.3
R311 VN.n55 VN.n0 86.8027
R312 VN.n111 VN.n56 86.8027
R313 VN.n21 VN.n20 56.5617
R314 VN.n34 VN.n33 56.5617
R315 VN.n77 VN.n76 56.5617
R316 VN.n90 VN.n89 56.5617
R317 VN.n14 VN.n13 55.106
R318 VN.n70 VN.n69 55.106
R319 VN VN.n111 52.6572
R320 VN.n69 VN.t6 47.3097
R321 VN.n13 VN.t8 47.3097
R322 VN.n47 VN.n46 41.5458
R323 VN.n103 VN.n102 41.5458
R324 VN.n47 VN.n2 39.6083
R325 VN.n103 VN.n58 39.6083
R326 VN.n15 VN.n12 24.5923
R327 VN.n19 VN.n12 24.5923
R328 VN.n20 VN.n19 24.5923
R329 VN.n21 VN.n10 24.5923
R330 VN.n25 VN.n10 24.5923
R331 VN.n26 VN.n25 24.5923
R332 VN.n28 VN.n8 24.5923
R333 VN.n32 VN.n8 24.5923
R334 VN.n33 VN.n32 24.5923
R335 VN.n34 VN.n6 24.5923
R336 VN.n38 VN.n6 24.5923
R337 VN.n39 VN.n38 24.5923
R338 VN.n41 VN.n4 24.5923
R339 VN.n45 VN.n4 24.5923
R340 VN.n46 VN.n45 24.5923
R341 VN.n51 VN.n2 24.5923
R342 VN.n52 VN.n51 24.5923
R343 VN.n53 VN.n52 24.5923
R344 VN.n76 VN.n75 24.5923
R345 VN.n75 VN.n68 24.5923
R346 VN.n71 VN.n68 24.5923
R347 VN.n89 VN.n88 24.5923
R348 VN.n88 VN.n64 24.5923
R349 VN.n84 VN.n64 24.5923
R350 VN.n82 VN.n81 24.5923
R351 VN.n81 VN.n66 24.5923
R352 VN.n77 VN.n66 24.5923
R353 VN.n102 VN.n101 24.5923
R354 VN.n101 VN.n60 24.5923
R355 VN.n97 VN.n60 24.5923
R356 VN.n95 VN.n94 24.5923
R357 VN.n94 VN.n62 24.5923
R358 VN.n90 VN.n62 24.5923
R359 VN.n109 VN.n108 24.5923
R360 VN.n108 VN.n107 24.5923
R361 VN.n107 VN.n58 24.5923
R362 VN.n15 VN.n14 20.1658
R363 VN.n40 VN.n39 20.1658
R364 VN.n71 VN.n70 20.1658
R365 VN.n96 VN.n95 20.1658
R366 VN.n14 VN.t5 14.2214
R367 VN.n27 VN.t7 14.2214
R368 VN.n40 VN.t4 14.2214
R369 VN.n0 VN.t3 14.2214
R370 VN.n70 VN.t9 14.2214
R371 VN.n83 VN.t2 14.2214
R372 VN.n96 VN.t1 14.2214
R373 VN.n56 VN.t0 14.2214
R374 VN.n27 VN.n26 12.2964
R375 VN.n28 VN.n27 12.2964
R376 VN.n84 VN.n83 12.2964
R377 VN.n83 VN.n82 12.2964
R378 VN.n41 VN.n40 4.42703
R379 VN.n97 VN.n96 4.42703
R380 VN.n53 VN.n0 3.44336
R381 VN.n109 VN.n56 3.44336
R382 VN.n16 VN.n13 2.44069
R383 VN.n72 VN.n69 2.44069
R384 VN.n111 VN.n110 0.354861
R385 VN.n55 VN.n54 0.354861
R386 VN VN.n55 0.267071
R387 VN.n110 VN.n57 0.189894
R388 VN.n106 VN.n57 0.189894
R389 VN.n106 VN.n105 0.189894
R390 VN.n105 VN.n104 0.189894
R391 VN.n104 VN.n59 0.189894
R392 VN.n100 VN.n59 0.189894
R393 VN.n100 VN.n99 0.189894
R394 VN.n99 VN.n98 0.189894
R395 VN.n98 VN.n61 0.189894
R396 VN.n93 VN.n61 0.189894
R397 VN.n93 VN.n92 0.189894
R398 VN.n92 VN.n91 0.189894
R399 VN.n91 VN.n63 0.189894
R400 VN.n87 VN.n63 0.189894
R401 VN.n87 VN.n86 0.189894
R402 VN.n86 VN.n85 0.189894
R403 VN.n85 VN.n65 0.189894
R404 VN.n80 VN.n65 0.189894
R405 VN.n80 VN.n79 0.189894
R406 VN.n79 VN.n78 0.189894
R407 VN.n78 VN.n67 0.189894
R408 VN.n74 VN.n67 0.189894
R409 VN.n74 VN.n73 0.189894
R410 VN.n73 VN.n72 0.189894
R411 VN.n17 VN.n16 0.189894
R412 VN.n18 VN.n17 0.189894
R413 VN.n18 VN.n11 0.189894
R414 VN.n22 VN.n11 0.189894
R415 VN.n23 VN.n22 0.189894
R416 VN.n24 VN.n23 0.189894
R417 VN.n24 VN.n9 0.189894
R418 VN.n29 VN.n9 0.189894
R419 VN.n30 VN.n29 0.189894
R420 VN.n31 VN.n30 0.189894
R421 VN.n31 VN.n7 0.189894
R422 VN.n35 VN.n7 0.189894
R423 VN.n36 VN.n35 0.189894
R424 VN.n37 VN.n36 0.189894
R425 VN.n37 VN.n5 0.189894
R426 VN.n42 VN.n5 0.189894
R427 VN.n43 VN.n42 0.189894
R428 VN.n44 VN.n43 0.189894
R429 VN.n44 VN.n3 0.189894
R430 VN.n48 VN.n3 0.189894
R431 VN.n49 VN.n48 0.189894
R432 VN.n50 VN.n49 0.189894
R433 VN.n50 VN.n1 0.189894
R434 VN.n54 VN.n1 0.189894
R435 VDD2.n1 VDD2.t1 193.075
R436 VDD2.n4 VDD2.t9 189.488
R437 VDD2.n3 VDD2.n2 177.74
R438 VDD2 VDD2.n7 177.738
R439 VDD2.n6 VDD2.n5 175.107
R440 VDD2.n1 VDD2.n0 175.106
R441 VDD2.n4 VDD2.n3 42.6981
R442 VDD2.n7 VDD2.t0 14.3832
R443 VDD2.n7 VDD2.t3 14.3832
R444 VDD2.n5 VDD2.t8 14.3832
R445 VDD2.n5 VDD2.t7 14.3832
R446 VDD2.n2 VDD2.t5 14.3832
R447 VDD2.n2 VDD2.t6 14.3832
R448 VDD2.n0 VDD2.t4 14.3832
R449 VDD2.n0 VDD2.t2 14.3832
R450 VDD2.n6 VDD2.n4 3.58671
R451 VDD2 VDD2.n6 0.955241
R452 VDD2.n3 VDD2.n1 0.841706
R453 B.n384 B.n147 585
R454 B.n383 B.n382 585
R455 B.n381 B.n148 585
R456 B.n380 B.n379 585
R457 B.n378 B.n149 585
R458 B.n377 B.n376 585
R459 B.n375 B.n150 585
R460 B.n374 B.n373 585
R461 B.n372 B.n151 585
R462 B.n371 B.n370 585
R463 B.n369 B.n152 585
R464 B.n368 B.n367 585
R465 B.n366 B.n153 585
R466 B.n364 B.n363 585
R467 B.n362 B.n156 585
R468 B.n361 B.n360 585
R469 B.n359 B.n157 585
R470 B.n358 B.n357 585
R471 B.n356 B.n158 585
R472 B.n355 B.n354 585
R473 B.n353 B.n159 585
R474 B.n352 B.n351 585
R475 B.n350 B.n160 585
R476 B.n349 B.n348 585
R477 B.n344 B.n161 585
R478 B.n343 B.n342 585
R479 B.n341 B.n162 585
R480 B.n340 B.n339 585
R481 B.n338 B.n163 585
R482 B.n337 B.n336 585
R483 B.n335 B.n164 585
R484 B.n334 B.n333 585
R485 B.n332 B.n165 585
R486 B.n331 B.n330 585
R487 B.n329 B.n166 585
R488 B.n328 B.n327 585
R489 B.n386 B.n385 585
R490 B.n387 B.n146 585
R491 B.n389 B.n388 585
R492 B.n390 B.n145 585
R493 B.n392 B.n391 585
R494 B.n393 B.n144 585
R495 B.n395 B.n394 585
R496 B.n396 B.n143 585
R497 B.n398 B.n397 585
R498 B.n399 B.n142 585
R499 B.n401 B.n400 585
R500 B.n402 B.n141 585
R501 B.n404 B.n403 585
R502 B.n405 B.n140 585
R503 B.n407 B.n406 585
R504 B.n408 B.n139 585
R505 B.n410 B.n409 585
R506 B.n411 B.n138 585
R507 B.n413 B.n412 585
R508 B.n414 B.n137 585
R509 B.n416 B.n415 585
R510 B.n417 B.n136 585
R511 B.n419 B.n418 585
R512 B.n420 B.n135 585
R513 B.n422 B.n421 585
R514 B.n423 B.n134 585
R515 B.n425 B.n424 585
R516 B.n426 B.n133 585
R517 B.n428 B.n427 585
R518 B.n429 B.n132 585
R519 B.n431 B.n430 585
R520 B.n432 B.n131 585
R521 B.n434 B.n433 585
R522 B.n435 B.n130 585
R523 B.n437 B.n436 585
R524 B.n438 B.n129 585
R525 B.n440 B.n439 585
R526 B.n441 B.n128 585
R527 B.n443 B.n442 585
R528 B.n444 B.n127 585
R529 B.n446 B.n445 585
R530 B.n447 B.n126 585
R531 B.n449 B.n448 585
R532 B.n450 B.n125 585
R533 B.n452 B.n451 585
R534 B.n453 B.n124 585
R535 B.n455 B.n454 585
R536 B.n456 B.n123 585
R537 B.n458 B.n457 585
R538 B.n459 B.n122 585
R539 B.n461 B.n460 585
R540 B.n462 B.n121 585
R541 B.n464 B.n463 585
R542 B.n465 B.n120 585
R543 B.n467 B.n466 585
R544 B.n468 B.n119 585
R545 B.n470 B.n469 585
R546 B.n471 B.n118 585
R547 B.n473 B.n472 585
R548 B.n474 B.n117 585
R549 B.n476 B.n475 585
R550 B.n477 B.n116 585
R551 B.n479 B.n478 585
R552 B.n480 B.n115 585
R553 B.n482 B.n481 585
R554 B.n483 B.n114 585
R555 B.n485 B.n484 585
R556 B.n486 B.n113 585
R557 B.n488 B.n487 585
R558 B.n489 B.n112 585
R559 B.n491 B.n490 585
R560 B.n492 B.n111 585
R561 B.n494 B.n493 585
R562 B.n495 B.n110 585
R563 B.n497 B.n496 585
R564 B.n498 B.n109 585
R565 B.n500 B.n499 585
R566 B.n501 B.n108 585
R567 B.n503 B.n502 585
R568 B.n504 B.n107 585
R569 B.n506 B.n505 585
R570 B.n507 B.n106 585
R571 B.n509 B.n508 585
R572 B.n510 B.n105 585
R573 B.n512 B.n511 585
R574 B.n513 B.n104 585
R575 B.n515 B.n514 585
R576 B.n516 B.n103 585
R577 B.n518 B.n517 585
R578 B.n519 B.n102 585
R579 B.n521 B.n520 585
R580 B.n522 B.n101 585
R581 B.n524 B.n523 585
R582 B.n525 B.n100 585
R583 B.n527 B.n526 585
R584 B.n528 B.n99 585
R585 B.n530 B.n529 585
R586 B.n531 B.n98 585
R587 B.n533 B.n532 585
R588 B.n534 B.n97 585
R589 B.n536 B.n535 585
R590 B.n537 B.n96 585
R591 B.n539 B.n538 585
R592 B.n540 B.n95 585
R593 B.n542 B.n541 585
R594 B.n543 B.n94 585
R595 B.n545 B.n544 585
R596 B.n546 B.n93 585
R597 B.n548 B.n547 585
R598 B.n549 B.n92 585
R599 B.n551 B.n550 585
R600 B.n552 B.n91 585
R601 B.n554 B.n553 585
R602 B.n555 B.n90 585
R603 B.n557 B.n556 585
R604 B.n558 B.n89 585
R605 B.n560 B.n559 585
R606 B.n561 B.n88 585
R607 B.n563 B.n562 585
R608 B.n564 B.n87 585
R609 B.n566 B.n565 585
R610 B.n567 B.n86 585
R611 B.n569 B.n568 585
R612 B.n570 B.n85 585
R613 B.n572 B.n571 585
R614 B.n573 B.n84 585
R615 B.n575 B.n574 585
R616 B.n576 B.n83 585
R617 B.n578 B.n577 585
R618 B.n579 B.n82 585
R619 B.n581 B.n580 585
R620 B.n582 B.n81 585
R621 B.n584 B.n583 585
R622 B.n585 B.n80 585
R623 B.n587 B.n586 585
R624 B.n588 B.n79 585
R625 B.n590 B.n589 585
R626 B.n591 B.n78 585
R627 B.n593 B.n592 585
R628 B.n594 B.n77 585
R629 B.n596 B.n595 585
R630 B.n597 B.n76 585
R631 B.n599 B.n598 585
R632 B.n600 B.n75 585
R633 B.n602 B.n601 585
R634 B.n603 B.n74 585
R635 B.n605 B.n604 585
R636 B.n606 B.n73 585
R637 B.n608 B.n607 585
R638 B.n609 B.n72 585
R639 B.n611 B.n610 585
R640 B.n612 B.n71 585
R641 B.n614 B.n613 585
R642 B.n615 B.n70 585
R643 B.n617 B.n616 585
R644 B.n618 B.n69 585
R645 B.n620 B.n619 585
R646 B.n621 B.n68 585
R647 B.n623 B.n622 585
R648 B.n624 B.n67 585
R649 B.n626 B.n625 585
R650 B.n627 B.n66 585
R651 B.n629 B.n628 585
R652 B.n630 B.n65 585
R653 B.n686 B.n685 585
R654 B.n684 B.n43 585
R655 B.n683 B.n682 585
R656 B.n681 B.n44 585
R657 B.n680 B.n679 585
R658 B.n678 B.n45 585
R659 B.n677 B.n676 585
R660 B.n675 B.n46 585
R661 B.n674 B.n673 585
R662 B.n672 B.n47 585
R663 B.n671 B.n670 585
R664 B.n669 B.n48 585
R665 B.n668 B.n667 585
R666 B.n665 B.n49 585
R667 B.n664 B.n663 585
R668 B.n662 B.n52 585
R669 B.n661 B.n660 585
R670 B.n659 B.n53 585
R671 B.n658 B.n657 585
R672 B.n656 B.n54 585
R673 B.n655 B.n654 585
R674 B.n653 B.n55 585
R675 B.n652 B.n651 585
R676 B.n650 B.n649 585
R677 B.n648 B.n59 585
R678 B.n647 B.n646 585
R679 B.n645 B.n60 585
R680 B.n644 B.n643 585
R681 B.n642 B.n61 585
R682 B.n641 B.n640 585
R683 B.n639 B.n62 585
R684 B.n638 B.n637 585
R685 B.n636 B.n63 585
R686 B.n635 B.n634 585
R687 B.n633 B.n64 585
R688 B.n632 B.n631 585
R689 B.n687 B.n42 585
R690 B.n689 B.n688 585
R691 B.n690 B.n41 585
R692 B.n692 B.n691 585
R693 B.n693 B.n40 585
R694 B.n695 B.n694 585
R695 B.n696 B.n39 585
R696 B.n698 B.n697 585
R697 B.n699 B.n38 585
R698 B.n701 B.n700 585
R699 B.n702 B.n37 585
R700 B.n704 B.n703 585
R701 B.n705 B.n36 585
R702 B.n707 B.n706 585
R703 B.n708 B.n35 585
R704 B.n710 B.n709 585
R705 B.n711 B.n34 585
R706 B.n713 B.n712 585
R707 B.n714 B.n33 585
R708 B.n716 B.n715 585
R709 B.n717 B.n32 585
R710 B.n719 B.n718 585
R711 B.n720 B.n31 585
R712 B.n722 B.n721 585
R713 B.n723 B.n30 585
R714 B.n725 B.n724 585
R715 B.n726 B.n29 585
R716 B.n728 B.n727 585
R717 B.n729 B.n28 585
R718 B.n731 B.n730 585
R719 B.n732 B.n27 585
R720 B.n734 B.n733 585
R721 B.n735 B.n26 585
R722 B.n737 B.n736 585
R723 B.n738 B.n25 585
R724 B.n740 B.n739 585
R725 B.n741 B.n24 585
R726 B.n743 B.n742 585
R727 B.n744 B.n23 585
R728 B.n746 B.n745 585
R729 B.n747 B.n22 585
R730 B.n749 B.n748 585
R731 B.n750 B.n21 585
R732 B.n752 B.n751 585
R733 B.n753 B.n20 585
R734 B.n755 B.n754 585
R735 B.n756 B.n19 585
R736 B.n758 B.n757 585
R737 B.n759 B.n18 585
R738 B.n761 B.n760 585
R739 B.n762 B.n17 585
R740 B.n764 B.n763 585
R741 B.n765 B.n16 585
R742 B.n767 B.n766 585
R743 B.n768 B.n15 585
R744 B.n770 B.n769 585
R745 B.n771 B.n14 585
R746 B.n773 B.n772 585
R747 B.n774 B.n13 585
R748 B.n776 B.n775 585
R749 B.n777 B.n12 585
R750 B.n779 B.n778 585
R751 B.n780 B.n11 585
R752 B.n782 B.n781 585
R753 B.n783 B.n10 585
R754 B.n785 B.n784 585
R755 B.n786 B.n9 585
R756 B.n788 B.n787 585
R757 B.n789 B.n8 585
R758 B.n791 B.n790 585
R759 B.n792 B.n7 585
R760 B.n794 B.n793 585
R761 B.n795 B.n6 585
R762 B.n797 B.n796 585
R763 B.n798 B.n5 585
R764 B.n800 B.n799 585
R765 B.n801 B.n4 585
R766 B.n803 B.n802 585
R767 B.n804 B.n3 585
R768 B.n806 B.n805 585
R769 B.n807 B.n0 585
R770 B.n2 B.n1 585
R771 B.n208 B.n207 585
R772 B.n209 B.n206 585
R773 B.n211 B.n210 585
R774 B.n212 B.n205 585
R775 B.n214 B.n213 585
R776 B.n215 B.n204 585
R777 B.n217 B.n216 585
R778 B.n218 B.n203 585
R779 B.n220 B.n219 585
R780 B.n221 B.n202 585
R781 B.n223 B.n222 585
R782 B.n224 B.n201 585
R783 B.n226 B.n225 585
R784 B.n227 B.n200 585
R785 B.n229 B.n228 585
R786 B.n230 B.n199 585
R787 B.n232 B.n231 585
R788 B.n233 B.n198 585
R789 B.n235 B.n234 585
R790 B.n236 B.n197 585
R791 B.n238 B.n237 585
R792 B.n239 B.n196 585
R793 B.n241 B.n240 585
R794 B.n242 B.n195 585
R795 B.n244 B.n243 585
R796 B.n245 B.n194 585
R797 B.n247 B.n246 585
R798 B.n248 B.n193 585
R799 B.n250 B.n249 585
R800 B.n251 B.n192 585
R801 B.n253 B.n252 585
R802 B.n254 B.n191 585
R803 B.n256 B.n255 585
R804 B.n257 B.n190 585
R805 B.n259 B.n258 585
R806 B.n260 B.n189 585
R807 B.n262 B.n261 585
R808 B.n263 B.n188 585
R809 B.n265 B.n264 585
R810 B.n266 B.n187 585
R811 B.n268 B.n267 585
R812 B.n269 B.n186 585
R813 B.n271 B.n270 585
R814 B.n272 B.n185 585
R815 B.n274 B.n273 585
R816 B.n275 B.n184 585
R817 B.n277 B.n276 585
R818 B.n278 B.n183 585
R819 B.n280 B.n279 585
R820 B.n281 B.n182 585
R821 B.n283 B.n282 585
R822 B.n284 B.n181 585
R823 B.n286 B.n285 585
R824 B.n287 B.n180 585
R825 B.n289 B.n288 585
R826 B.n290 B.n179 585
R827 B.n292 B.n291 585
R828 B.n293 B.n178 585
R829 B.n295 B.n294 585
R830 B.n296 B.n177 585
R831 B.n298 B.n297 585
R832 B.n299 B.n176 585
R833 B.n301 B.n300 585
R834 B.n302 B.n175 585
R835 B.n304 B.n303 585
R836 B.n305 B.n174 585
R837 B.n307 B.n306 585
R838 B.n308 B.n173 585
R839 B.n310 B.n309 585
R840 B.n311 B.n172 585
R841 B.n313 B.n312 585
R842 B.n314 B.n171 585
R843 B.n316 B.n315 585
R844 B.n317 B.n170 585
R845 B.n319 B.n318 585
R846 B.n320 B.n169 585
R847 B.n322 B.n321 585
R848 B.n323 B.n168 585
R849 B.n325 B.n324 585
R850 B.n326 B.n167 585
R851 B.n328 B.n167 463.671
R852 B.n386 B.n147 463.671
R853 B.n632 B.n65 463.671
R854 B.n687 B.n686 463.671
R855 B.n809 B.n808 256.663
R856 B.n154 B.t7 254.298
R857 B.n56 B.t11 254.298
R858 B.n345 B.t4 254.298
R859 B.n50 B.t2 254.298
R860 B.n808 B.n807 235.042
R861 B.n808 B.n2 235.042
R862 B.n345 B.t3 223.588
R863 B.n154 B.t6 223.588
R864 B.n56 B.t9 223.588
R865 B.n50 B.t0 223.588
R866 B.n155 B.t8 173.619
R867 B.n57 B.t10 173.619
R868 B.n346 B.t5 173.619
R869 B.n51 B.t1 173.619
R870 B.n329 B.n328 163.367
R871 B.n330 B.n329 163.367
R872 B.n330 B.n165 163.367
R873 B.n334 B.n165 163.367
R874 B.n335 B.n334 163.367
R875 B.n336 B.n335 163.367
R876 B.n336 B.n163 163.367
R877 B.n340 B.n163 163.367
R878 B.n341 B.n340 163.367
R879 B.n342 B.n341 163.367
R880 B.n342 B.n161 163.367
R881 B.n349 B.n161 163.367
R882 B.n350 B.n349 163.367
R883 B.n351 B.n350 163.367
R884 B.n351 B.n159 163.367
R885 B.n355 B.n159 163.367
R886 B.n356 B.n355 163.367
R887 B.n357 B.n356 163.367
R888 B.n357 B.n157 163.367
R889 B.n361 B.n157 163.367
R890 B.n362 B.n361 163.367
R891 B.n363 B.n362 163.367
R892 B.n363 B.n153 163.367
R893 B.n368 B.n153 163.367
R894 B.n369 B.n368 163.367
R895 B.n370 B.n369 163.367
R896 B.n370 B.n151 163.367
R897 B.n374 B.n151 163.367
R898 B.n375 B.n374 163.367
R899 B.n376 B.n375 163.367
R900 B.n376 B.n149 163.367
R901 B.n380 B.n149 163.367
R902 B.n381 B.n380 163.367
R903 B.n382 B.n381 163.367
R904 B.n382 B.n147 163.367
R905 B.n628 B.n65 163.367
R906 B.n628 B.n627 163.367
R907 B.n627 B.n626 163.367
R908 B.n626 B.n67 163.367
R909 B.n622 B.n67 163.367
R910 B.n622 B.n621 163.367
R911 B.n621 B.n620 163.367
R912 B.n620 B.n69 163.367
R913 B.n616 B.n69 163.367
R914 B.n616 B.n615 163.367
R915 B.n615 B.n614 163.367
R916 B.n614 B.n71 163.367
R917 B.n610 B.n71 163.367
R918 B.n610 B.n609 163.367
R919 B.n609 B.n608 163.367
R920 B.n608 B.n73 163.367
R921 B.n604 B.n73 163.367
R922 B.n604 B.n603 163.367
R923 B.n603 B.n602 163.367
R924 B.n602 B.n75 163.367
R925 B.n598 B.n75 163.367
R926 B.n598 B.n597 163.367
R927 B.n597 B.n596 163.367
R928 B.n596 B.n77 163.367
R929 B.n592 B.n77 163.367
R930 B.n592 B.n591 163.367
R931 B.n591 B.n590 163.367
R932 B.n590 B.n79 163.367
R933 B.n586 B.n79 163.367
R934 B.n586 B.n585 163.367
R935 B.n585 B.n584 163.367
R936 B.n584 B.n81 163.367
R937 B.n580 B.n81 163.367
R938 B.n580 B.n579 163.367
R939 B.n579 B.n578 163.367
R940 B.n578 B.n83 163.367
R941 B.n574 B.n83 163.367
R942 B.n574 B.n573 163.367
R943 B.n573 B.n572 163.367
R944 B.n572 B.n85 163.367
R945 B.n568 B.n85 163.367
R946 B.n568 B.n567 163.367
R947 B.n567 B.n566 163.367
R948 B.n566 B.n87 163.367
R949 B.n562 B.n87 163.367
R950 B.n562 B.n561 163.367
R951 B.n561 B.n560 163.367
R952 B.n560 B.n89 163.367
R953 B.n556 B.n89 163.367
R954 B.n556 B.n555 163.367
R955 B.n555 B.n554 163.367
R956 B.n554 B.n91 163.367
R957 B.n550 B.n91 163.367
R958 B.n550 B.n549 163.367
R959 B.n549 B.n548 163.367
R960 B.n548 B.n93 163.367
R961 B.n544 B.n93 163.367
R962 B.n544 B.n543 163.367
R963 B.n543 B.n542 163.367
R964 B.n542 B.n95 163.367
R965 B.n538 B.n95 163.367
R966 B.n538 B.n537 163.367
R967 B.n537 B.n536 163.367
R968 B.n536 B.n97 163.367
R969 B.n532 B.n97 163.367
R970 B.n532 B.n531 163.367
R971 B.n531 B.n530 163.367
R972 B.n530 B.n99 163.367
R973 B.n526 B.n99 163.367
R974 B.n526 B.n525 163.367
R975 B.n525 B.n524 163.367
R976 B.n524 B.n101 163.367
R977 B.n520 B.n101 163.367
R978 B.n520 B.n519 163.367
R979 B.n519 B.n518 163.367
R980 B.n518 B.n103 163.367
R981 B.n514 B.n103 163.367
R982 B.n514 B.n513 163.367
R983 B.n513 B.n512 163.367
R984 B.n512 B.n105 163.367
R985 B.n508 B.n105 163.367
R986 B.n508 B.n507 163.367
R987 B.n507 B.n506 163.367
R988 B.n506 B.n107 163.367
R989 B.n502 B.n107 163.367
R990 B.n502 B.n501 163.367
R991 B.n501 B.n500 163.367
R992 B.n500 B.n109 163.367
R993 B.n496 B.n109 163.367
R994 B.n496 B.n495 163.367
R995 B.n495 B.n494 163.367
R996 B.n494 B.n111 163.367
R997 B.n490 B.n111 163.367
R998 B.n490 B.n489 163.367
R999 B.n489 B.n488 163.367
R1000 B.n488 B.n113 163.367
R1001 B.n484 B.n113 163.367
R1002 B.n484 B.n483 163.367
R1003 B.n483 B.n482 163.367
R1004 B.n482 B.n115 163.367
R1005 B.n478 B.n115 163.367
R1006 B.n478 B.n477 163.367
R1007 B.n477 B.n476 163.367
R1008 B.n476 B.n117 163.367
R1009 B.n472 B.n117 163.367
R1010 B.n472 B.n471 163.367
R1011 B.n471 B.n470 163.367
R1012 B.n470 B.n119 163.367
R1013 B.n466 B.n119 163.367
R1014 B.n466 B.n465 163.367
R1015 B.n465 B.n464 163.367
R1016 B.n464 B.n121 163.367
R1017 B.n460 B.n121 163.367
R1018 B.n460 B.n459 163.367
R1019 B.n459 B.n458 163.367
R1020 B.n458 B.n123 163.367
R1021 B.n454 B.n123 163.367
R1022 B.n454 B.n453 163.367
R1023 B.n453 B.n452 163.367
R1024 B.n452 B.n125 163.367
R1025 B.n448 B.n125 163.367
R1026 B.n448 B.n447 163.367
R1027 B.n447 B.n446 163.367
R1028 B.n446 B.n127 163.367
R1029 B.n442 B.n127 163.367
R1030 B.n442 B.n441 163.367
R1031 B.n441 B.n440 163.367
R1032 B.n440 B.n129 163.367
R1033 B.n436 B.n129 163.367
R1034 B.n436 B.n435 163.367
R1035 B.n435 B.n434 163.367
R1036 B.n434 B.n131 163.367
R1037 B.n430 B.n131 163.367
R1038 B.n430 B.n429 163.367
R1039 B.n429 B.n428 163.367
R1040 B.n428 B.n133 163.367
R1041 B.n424 B.n133 163.367
R1042 B.n424 B.n423 163.367
R1043 B.n423 B.n422 163.367
R1044 B.n422 B.n135 163.367
R1045 B.n418 B.n135 163.367
R1046 B.n418 B.n417 163.367
R1047 B.n417 B.n416 163.367
R1048 B.n416 B.n137 163.367
R1049 B.n412 B.n137 163.367
R1050 B.n412 B.n411 163.367
R1051 B.n411 B.n410 163.367
R1052 B.n410 B.n139 163.367
R1053 B.n406 B.n139 163.367
R1054 B.n406 B.n405 163.367
R1055 B.n405 B.n404 163.367
R1056 B.n404 B.n141 163.367
R1057 B.n400 B.n141 163.367
R1058 B.n400 B.n399 163.367
R1059 B.n399 B.n398 163.367
R1060 B.n398 B.n143 163.367
R1061 B.n394 B.n143 163.367
R1062 B.n394 B.n393 163.367
R1063 B.n393 B.n392 163.367
R1064 B.n392 B.n145 163.367
R1065 B.n388 B.n145 163.367
R1066 B.n388 B.n387 163.367
R1067 B.n387 B.n386 163.367
R1068 B.n686 B.n43 163.367
R1069 B.n682 B.n43 163.367
R1070 B.n682 B.n681 163.367
R1071 B.n681 B.n680 163.367
R1072 B.n680 B.n45 163.367
R1073 B.n676 B.n45 163.367
R1074 B.n676 B.n675 163.367
R1075 B.n675 B.n674 163.367
R1076 B.n674 B.n47 163.367
R1077 B.n670 B.n47 163.367
R1078 B.n670 B.n669 163.367
R1079 B.n669 B.n668 163.367
R1080 B.n668 B.n49 163.367
R1081 B.n663 B.n49 163.367
R1082 B.n663 B.n662 163.367
R1083 B.n662 B.n661 163.367
R1084 B.n661 B.n53 163.367
R1085 B.n657 B.n53 163.367
R1086 B.n657 B.n656 163.367
R1087 B.n656 B.n655 163.367
R1088 B.n655 B.n55 163.367
R1089 B.n651 B.n55 163.367
R1090 B.n651 B.n650 163.367
R1091 B.n650 B.n59 163.367
R1092 B.n646 B.n59 163.367
R1093 B.n646 B.n645 163.367
R1094 B.n645 B.n644 163.367
R1095 B.n644 B.n61 163.367
R1096 B.n640 B.n61 163.367
R1097 B.n640 B.n639 163.367
R1098 B.n639 B.n638 163.367
R1099 B.n638 B.n63 163.367
R1100 B.n634 B.n63 163.367
R1101 B.n634 B.n633 163.367
R1102 B.n633 B.n632 163.367
R1103 B.n688 B.n687 163.367
R1104 B.n688 B.n41 163.367
R1105 B.n692 B.n41 163.367
R1106 B.n693 B.n692 163.367
R1107 B.n694 B.n693 163.367
R1108 B.n694 B.n39 163.367
R1109 B.n698 B.n39 163.367
R1110 B.n699 B.n698 163.367
R1111 B.n700 B.n699 163.367
R1112 B.n700 B.n37 163.367
R1113 B.n704 B.n37 163.367
R1114 B.n705 B.n704 163.367
R1115 B.n706 B.n705 163.367
R1116 B.n706 B.n35 163.367
R1117 B.n710 B.n35 163.367
R1118 B.n711 B.n710 163.367
R1119 B.n712 B.n711 163.367
R1120 B.n712 B.n33 163.367
R1121 B.n716 B.n33 163.367
R1122 B.n717 B.n716 163.367
R1123 B.n718 B.n717 163.367
R1124 B.n718 B.n31 163.367
R1125 B.n722 B.n31 163.367
R1126 B.n723 B.n722 163.367
R1127 B.n724 B.n723 163.367
R1128 B.n724 B.n29 163.367
R1129 B.n728 B.n29 163.367
R1130 B.n729 B.n728 163.367
R1131 B.n730 B.n729 163.367
R1132 B.n730 B.n27 163.367
R1133 B.n734 B.n27 163.367
R1134 B.n735 B.n734 163.367
R1135 B.n736 B.n735 163.367
R1136 B.n736 B.n25 163.367
R1137 B.n740 B.n25 163.367
R1138 B.n741 B.n740 163.367
R1139 B.n742 B.n741 163.367
R1140 B.n742 B.n23 163.367
R1141 B.n746 B.n23 163.367
R1142 B.n747 B.n746 163.367
R1143 B.n748 B.n747 163.367
R1144 B.n748 B.n21 163.367
R1145 B.n752 B.n21 163.367
R1146 B.n753 B.n752 163.367
R1147 B.n754 B.n753 163.367
R1148 B.n754 B.n19 163.367
R1149 B.n758 B.n19 163.367
R1150 B.n759 B.n758 163.367
R1151 B.n760 B.n759 163.367
R1152 B.n760 B.n17 163.367
R1153 B.n764 B.n17 163.367
R1154 B.n765 B.n764 163.367
R1155 B.n766 B.n765 163.367
R1156 B.n766 B.n15 163.367
R1157 B.n770 B.n15 163.367
R1158 B.n771 B.n770 163.367
R1159 B.n772 B.n771 163.367
R1160 B.n772 B.n13 163.367
R1161 B.n776 B.n13 163.367
R1162 B.n777 B.n776 163.367
R1163 B.n778 B.n777 163.367
R1164 B.n778 B.n11 163.367
R1165 B.n782 B.n11 163.367
R1166 B.n783 B.n782 163.367
R1167 B.n784 B.n783 163.367
R1168 B.n784 B.n9 163.367
R1169 B.n788 B.n9 163.367
R1170 B.n789 B.n788 163.367
R1171 B.n790 B.n789 163.367
R1172 B.n790 B.n7 163.367
R1173 B.n794 B.n7 163.367
R1174 B.n795 B.n794 163.367
R1175 B.n796 B.n795 163.367
R1176 B.n796 B.n5 163.367
R1177 B.n800 B.n5 163.367
R1178 B.n801 B.n800 163.367
R1179 B.n802 B.n801 163.367
R1180 B.n802 B.n3 163.367
R1181 B.n806 B.n3 163.367
R1182 B.n807 B.n806 163.367
R1183 B.n208 B.n2 163.367
R1184 B.n209 B.n208 163.367
R1185 B.n210 B.n209 163.367
R1186 B.n210 B.n205 163.367
R1187 B.n214 B.n205 163.367
R1188 B.n215 B.n214 163.367
R1189 B.n216 B.n215 163.367
R1190 B.n216 B.n203 163.367
R1191 B.n220 B.n203 163.367
R1192 B.n221 B.n220 163.367
R1193 B.n222 B.n221 163.367
R1194 B.n222 B.n201 163.367
R1195 B.n226 B.n201 163.367
R1196 B.n227 B.n226 163.367
R1197 B.n228 B.n227 163.367
R1198 B.n228 B.n199 163.367
R1199 B.n232 B.n199 163.367
R1200 B.n233 B.n232 163.367
R1201 B.n234 B.n233 163.367
R1202 B.n234 B.n197 163.367
R1203 B.n238 B.n197 163.367
R1204 B.n239 B.n238 163.367
R1205 B.n240 B.n239 163.367
R1206 B.n240 B.n195 163.367
R1207 B.n244 B.n195 163.367
R1208 B.n245 B.n244 163.367
R1209 B.n246 B.n245 163.367
R1210 B.n246 B.n193 163.367
R1211 B.n250 B.n193 163.367
R1212 B.n251 B.n250 163.367
R1213 B.n252 B.n251 163.367
R1214 B.n252 B.n191 163.367
R1215 B.n256 B.n191 163.367
R1216 B.n257 B.n256 163.367
R1217 B.n258 B.n257 163.367
R1218 B.n258 B.n189 163.367
R1219 B.n262 B.n189 163.367
R1220 B.n263 B.n262 163.367
R1221 B.n264 B.n263 163.367
R1222 B.n264 B.n187 163.367
R1223 B.n268 B.n187 163.367
R1224 B.n269 B.n268 163.367
R1225 B.n270 B.n269 163.367
R1226 B.n270 B.n185 163.367
R1227 B.n274 B.n185 163.367
R1228 B.n275 B.n274 163.367
R1229 B.n276 B.n275 163.367
R1230 B.n276 B.n183 163.367
R1231 B.n280 B.n183 163.367
R1232 B.n281 B.n280 163.367
R1233 B.n282 B.n281 163.367
R1234 B.n282 B.n181 163.367
R1235 B.n286 B.n181 163.367
R1236 B.n287 B.n286 163.367
R1237 B.n288 B.n287 163.367
R1238 B.n288 B.n179 163.367
R1239 B.n292 B.n179 163.367
R1240 B.n293 B.n292 163.367
R1241 B.n294 B.n293 163.367
R1242 B.n294 B.n177 163.367
R1243 B.n298 B.n177 163.367
R1244 B.n299 B.n298 163.367
R1245 B.n300 B.n299 163.367
R1246 B.n300 B.n175 163.367
R1247 B.n304 B.n175 163.367
R1248 B.n305 B.n304 163.367
R1249 B.n306 B.n305 163.367
R1250 B.n306 B.n173 163.367
R1251 B.n310 B.n173 163.367
R1252 B.n311 B.n310 163.367
R1253 B.n312 B.n311 163.367
R1254 B.n312 B.n171 163.367
R1255 B.n316 B.n171 163.367
R1256 B.n317 B.n316 163.367
R1257 B.n318 B.n317 163.367
R1258 B.n318 B.n169 163.367
R1259 B.n322 B.n169 163.367
R1260 B.n323 B.n322 163.367
R1261 B.n324 B.n323 163.367
R1262 B.n324 B.n167 163.367
R1263 B.n346 B.n345 80.6793
R1264 B.n155 B.n154 80.6793
R1265 B.n57 B.n56 80.6793
R1266 B.n51 B.n50 80.6793
R1267 B.n347 B.n346 59.5399
R1268 B.n365 B.n155 59.5399
R1269 B.n58 B.n57 59.5399
R1270 B.n666 B.n51 59.5399
R1271 B.n385 B.n384 30.1273
R1272 B.n685 B.n42 30.1273
R1273 B.n631 B.n630 30.1273
R1274 B.n327 B.n326 30.1273
R1275 B B.n809 18.0485
R1276 B.n689 B.n42 10.6151
R1277 B.n690 B.n689 10.6151
R1278 B.n691 B.n690 10.6151
R1279 B.n691 B.n40 10.6151
R1280 B.n695 B.n40 10.6151
R1281 B.n696 B.n695 10.6151
R1282 B.n697 B.n696 10.6151
R1283 B.n697 B.n38 10.6151
R1284 B.n701 B.n38 10.6151
R1285 B.n702 B.n701 10.6151
R1286 B.n703 B.n702 10.6151
R1287 B.n703 B.n36 10.6151
R1288 B.n707 B.n36 10.6151
R1289 B.n708 B.n707 10.6151
R1290 B.n709 B.n708 10.6151
R1291 B.n709 B.n34 10.6151
R1292 B.n713 B.n34 10.6151
R1293 B.n714 B.n713 10.6151
R1294 B.n715 B.n714 10.6151
R1295 B.n715 B.n32 10.6151
R1296 B.n719 B.n32 10.6151
R1297 B.n720 B.n719 10.6151
R1298 B.n721 B.n720 10.6151
R1299 B.n721 B.n30 10.6151
R1300 B.n725 B.n30 10.6151
R1301 B.n726 B.n725 10.6151
R1302 B.n727 B.n726 10.6151
R1303 B.n727 B.n28 10.6151
R1304 B.n731 B.n28 10.6151
R1305 B.n732 B.n731 10.6151
R1306 B.n733 B.n732 10.6151
R1307 B.n733 B.n26 10.6151
R1308 B.n737 B.n26 10.6151
R1309 B.n738 B.n737 10.6151
R1310 B.n739 B.n738 10.6151
R1311 B.n739 B.n24 10.6151
R1312 B.n743 B.n24 10.6151
R1313 B.n744 B.n743 10.6151
R1314 B.n745 B.n744 10.6151
R1315 B.n745 B.n22 10.6151
R1316 B.n749 B.n22 10.6151
R1317 B.n750 B.n749 10.6151
R1318 B.n751 B.n750 10.6151
R1319 B.n751 B.n20 10.6151
R1320 B.n755 B.n20 10.6151
R1321 B.n756 B.n755 10.6151
R1322 B.n757 B.n756 10.6151
R1323 B.n757 B.n18 10.6151
R1324 B.n761 B.n18 10.6151
R1325 B.n762 B.n761 10.6151
R1326 B.n763 B.n762 10.6151
R1327 B.n763 B.n16 10.6151
R1328 B.n767 B.n16 10.6151
R1329 B.n768 B.n767 10.6151
R1330 B.n769 B.n768 10.6151
R1331 B.n769 B.n14 10.6151
R1332 B.n773 B.n14 10.6151
R1333 B.n774 B.n773 10.6151
R1334 B.n775 B.n774 10.6151
R1335 B.n775 B.n12 10.6151
R1336 B.n779 B.n12 10.6151
R1337 B.n780 B.n779 10.6151
R1338 B.n781 B.n780 10.6151
R1339 B.n781 B.n10 10.6151
R1340 B.n785 B.n10 10.6151
R1341 B.n786 B.n785 10.6151
R1342 B.n787 B.n786 10.6151
R1343 B.n787 B.n8 10.6151
R1344 B.n791 B.n8 10.6151
R1345 B.n792 B.n791 10.6151
R1346 B.n793 B.n792 10.6151
R1347 B.n793 B.n6 10.6151
R1348 B.n797 B.n6 10.6151
R1349 B.n798 B.n797 10.6151
R1350 B.n799 B.n798 10.6151
R1351 B.n799 B.n4 10.6151
R1352 B.n803 B.n4 10.6151
R1353 B.n804 B.n803 10.6151
R1354 B.n805 B.n804 10.6151
R1355 B.n805 B.n0 10.6151
R1356 B.n685 B.n684 10.6151
R1357 B.n684 B.n683 10.6151
R1358 B.n683 B.n44 10.6151
R1359 B.n679 B.n44 10.6151
R1360 B.n679 B.n678 10.6151
R1361 B.n678 B.n677 10.6151
R1362 B.n677 B.n46 10.6151
R1363 B.n673 B.n46 10.6151
R1364 B.n673 B.n672 10.6151
R1365 B.n672 B.n671 10.6151
R1366 B.n671 B.n48 10.6151
R1367 B.n667 B.n48 10.6151
R1368 B.n665 B.n664 10.6151
R1369 B.n664 B.n52 10.6151
R1370 B.n660 B.n52 10.6151
R1371 B.n660 B.n659 10.6151
R1372 B.n659 B.n658 10.6151
R1373 B.n658 B.n54 10.6151
R1374 B.n654 B.n54 10.6151
R1375 B.n654 B.n653 10.6151
R1376 B.n653 B.n652 10.6151
R1377 B.n649 B.n648 10.6151
R1378 B.n648 B.n647 10.6151
R1379 B.n647 B.n60 10.6151
R1380 B.n643 B.n60 10.6151
R1381 B.n643 B.n642 10.6151
R1382 B.n642 B.n641 10.6151
R1383 B.n641 B.n62 10.6151
R1384 B.n637 B.n62 10.6151
R1385 B.n637 B.n636 10.6151
R1386 B.n636 B.n635 10.6151
R1387 B.n635 B.n64 10.6151
R1388 B.n631 B.n64 10.6151
R1389 B.n630 B.n629 10.6151
R1390 B.n629 B.n66 10.6151
R1391 B.n625 B.n66 10.6151
R1392 B.n625 B.n624 10.6151
R1393 B.n624 B.n623 10.6151
R1394 B.n623 B.n68 10.6151
R1395 B.n619 B.n68 10.6151
R1396 B.n619 B.n618 10.6151
R1397 B.n618 B.n617 10.6151
R1398 B.n617 B.n70 10.6151
R1399 B.n613 B.n70 10.6151
R1400 B.n613 B.n612 10.6151
R1401 B.n612 B.n611 10.6151
R1402 B.n611 B.n72 10.6151
R1403 B.n607 B.n72 10.6151
R1404 B.n607 B.n606 10.6151
R1405 B.n606 B.n605 10.6151
R1406 B.n605 B.n74 10.6151
R1407 B.n601 B.n74 10.6151
R1408 B.n601 B.n600 10.6151
R1409 B.n600 B.n599 10.6151
R1410 B.n599 B.n76 10.6151
R1411 B.n595 B.n76 10.6151
R1412 B.n595 B.n594 10.6151
R1413 B.n594 B.n593 10.6151
R1414 B.n593 B.n78 10.6151
R1415 B.n589 B.n78 10.6151
R1416 B.n589 B.n588 10.6151
R1417 B.n588 B.n587 10.6151
R1418 B.n587 B.n80 10.6151
R1419 B.n583 B.n80 10.6151
R1420 B.n583 B.n582 10.6151
R1421 B.n582 B.n581 10.6151
R1422 B.n581 B.n82 10.6151
R1423 B.n577 B.n82 10.6151
R1424 B.n577 B.n576 10.6151
R1425 B.n576 B.n575 10.6151
R1426 B.n575 B.n84 10.6151
R1427 B.n571 B.n84 10.6151
R1428 B.n571 B.n570 10.6151
R1429 B.n570 B.n569 10.6151
R1430 B.n569 B.n86 10.6151
R1431 B.n565 B.n86 10.6151
R1432 B.n565 B.n564 10.6151
R1433 B.n564 B.n563 10.6151
R1434 B.n563 B.n88 10.6151
R1435 B.n559 B.n88 10.6151
R1436 B.n559 B.n558 10.6151
R1437 B.n558 B.n557 10.6151
R1438 B.n557 B.n90 10.6151
R1439 B.n553 B.n90 10.6151
R1440 B.n553 B.n552 10.6151
R1441 B.n552 B.n551 10.6151
R1442 B.n551 B.n92 10.6151
R1443 B.n547 B.n92 10.6151
R1444 B.n547 B.n546 10.6151
R1445 B.n546 B.n545 10.6151
R1446 B.n545 B.n94 10.6151
R1447 B.n541 B.n94 10.6151
R1448 B.n541 B.n540 10.6151
R1449 B.n540 B.n539 10.6151
R1450 B.n539 B.n96 10.6151
R1451 B.n535 B.n96 10.6151
R1452 B.n535 B.n534 10.6151
R1453 B.n534 B.n533 10.6151
R1454 B.n533 B.n98 10.6151
R1455 B.n529 B.n98 10.6151
R1456 B.n529 B.n528 10.6151
R1457 B.n528 B.n527 10.6151
R1458 B.n527 B.n100 10.6151
R1459 B.n523 B.n100 10.6151
R1460 B.n523 B.n522 10.6151
R1461 B.n522 B.n521 10.6151
R1462 B.n521 B.n102 10.6151
R1463 B.n517 B.n102 10.6151
R1464 B.n517 B.n516 10.6151
R1465 B.n516 B.n515 10.6151
R1466 B.n515 B.n104 10.6151
R1467 B.n511 B.n104 10.6151
R1468 B.n511 B.n510 10.6151
R1469 B.n510 B.n509 10.6151
R1470 B.n509 B.n106 10.6151
R1471 B.n505 B.n106 10.6151
R1472 B.n505 B.n504 10.6151
R1473 B.n504 B.n503 10.6151
R1474 B.n503 B.n108 10.6151
R1475 B.n499 B.n108 10.6151
R1476 B.n499 B.n498 10.6151
R1477 B.n498 B.n497 10.6151
R1478 B.n497 B.n110 10.6151
R1479 B.n493 B.n110 10.6151
R1480 B.n493 B.n492 10.6151
R1481 B.n492 B.n491 10.6151
R1482 B.n491 B.n112 10.6151
R1483 B.n487 B.n112 10.6151
R1484 B.n487 B.n486 10.6151
R1485 B.n486 B.n485 10.6151
R1486 B.n485 B.n114 10.6151
R1487 B.n481 B.n114 10.6151
R1488 B.n481 B.n480 10.6151
R1489 B.n480 B.n479 10.6151
R1490 B.n479 B.n116 10.6151
R1491 B.n475 B.n116 10.6151
R1492 B.n475 B.n474 10.6151
R1493 B.n474 B.n473 10.6151
R1494 B.n473 B.n118 10.6151
R1495 B.n469 B.n118 10.6151
R1496 B.n469 B.n468 10.6151
R1497 B.n468 B.n467 10.6151
R1498 B.n467 B.n120 10.6151
R1499 B.n463 B.n120 10.6151
R1500 B.n463 B.n462 10.6151
R1501 B.n462 B.n461 10.6151
R1502 B.n461 B.n122 10.6151
R1503 B.n457 B.n122 10.6151
R1504 B.n457 B.n456 10.6151
R1505 B.n456 B.n455 10.6151
R1506 B.n455 B.n124 10.6151
R1507 B.n451 B.n124 10.6151
R1508 B.n451 B.n450 10.6151
R1509 B.n450 B.n449 10.6151
R1510 B.n449 B.n126 10.6151
R1511 B.n445 B.n126 10.6151
R1512 B.n445 B.n444 10.6151
R1513 B.n444 B.n443 10.6151
R1514 B.n443 B.n128 10.6151
R1515 B.n439 B.n128 10.6151
R1516 B.n439 B.n438 10.6151
R1517 B.n438 B.n437 10.6151
R1518 B.n437 B.n130 10.6151
R1519 B.n433 B.n130 10.6151
R1520 B.n433 B.n432 10.6151
R1521 B.n432 B.n431 10.6151
R1522 B.n431 B.n132 10.6151
R1523 B.n427 B.n132 10.6151
R1524 B.n427 B.n426 10.6151
R1525 B.n426 B.n425 10.6151
R1526 B.n425 B.n134 10.6151
R1527 B.n421 B.n134 10.6151
R1528 B.n421 B.n420 10.6151
R1529 B.n420 B.n419 10.6151
R1530 B.n419 B.n136 10.6151
R1531 B.n415 B.n136 10.6151
R1532 B.n415 B.n414 10.6151
R1533 B.n414 B.n413 10.6151
R1534 B.n413 B.n138 10.6151
R1535 B.n409 B.n138 10.6151
R1536 B.n409 B.n408 10.6151
R1537 B.n408 B.n407 10.6151
R1538 B.n407 B.n140 10.6151
R1539 B.n403 B.n140 10.6151
R1540 B.n403 B.n402 10.6151
R1541 B.n402 B.n401 10.6151
R1542 B.n401 B.n142 10.6151
R1543 B.n397 B.n142 10.6151
R1544 B.n397 B.n396 10.6151
R1545 B.n396 B.n395 10.6151
R1546 B.n395 B.n144 10.6151
R1547 B.n391 B.n144 10.6151
R1548 B.n391 B.n390 10.6151
R1549 B.n390 B.n389 10.6151
R1550 B.n389 B.n146 10.6151
R1551 B.n385 B.n146 10.6151
R1552 B.n207 B.n1 10.6151
R1553 B.n207 B.n206 10.6151
R1554 B.n211 B.n206 10.6151
R1555 B.n212 B.n211 10.6151
R1556 B.n213 B.n212 10.6151
R1557 B.n213 B.n204 10.6151
R1558 B.n217 B.n204 10.6151
R1559 B.n218 B.n217 10.6151
R1560 B.n219 B.n218 10.6151
R1561 B.n219 B.n202 10.6151
R1562 B.n223 B.n202 10.6151
R1563 B.n224 B.n223 10.6151
R1564 B.n225 B.n224 10.6151
R1565 B.n225 B.n200 10.6151
R1566 B.n229 B.n200 10.6151
R1567 B.n230 B.n229 10.6151
R1568 B.n231 B.n230 10.6151
R1569 B.n231 B.n198 10.6151
R1570 B.n235 B.n198 10.6151
R1571 B.n236 B.n235 10.6151
R1572 B.n237 B.n236 10.6151
R1573 B.n237 B.n196 10.6151
R1574 B.n241 B.n196 10.6151
R1575 B.n242 B.n241 10.6151
R1576 B.n243 B.n242 10.6151
R1577 B.n243 B.n194 10.6151
R1578 B.n247 B.n194 10.6151
R1579 B.n248 B.n247 10.6151
R1580 B.n249 B.n248 10.6151
R1581 B.n249 B.n192 10.6151
R1582 B.n253 B.n192 10.6151
R1583 B.n254 B.n253 10.6151
R1584 B.n255 B.n254 10.6151
R1585 B.n255 B.n190 10.6151
R1586 B.n259 B.n190 10.6151
R1587 B.n260 B.n259 10.6151
R1588 B.n261 B.n260 10.6151
R1589 B.n261 B.n188 10.6151
R1590 B.n265 B.n188 10.6151
R1591 B.n266 B.n265 10.6151
R1592 B.n267 B.n266 10.6151
R1593 B.n267 B.n186 10.6151
R1594 B.n271 B.n186 10.6151
R1595 B.n272 B.n271 10.6151
R1596 B.n273 B.n272 10.6151
R1597 B.n273 B.n184 10.6151
R1598 B.n277 B.n184 10.6151
R1599 B.n278 B.n277 10.6151
R1600 B.n279 B.n278 10.6151
R1601 B.n279 B.n182 10.6151
R1602 B.n283 B.n182 10.6151
R1603 B.n284 B.n283 10.6151
R1604 B.n285 B.n284 10.6151
R1605 B.n285 B.n180 10.6151
R1606 B.n289 B.n180 10.6151
R1607 B.n290 B.n289 10.6151
R1608 B.n291 B.n290 10.6151
R1609 B.n291 B.n178 10.6151
R1610 B.n295 B.n178 10.6151
R1611 B.n296 B.n295 10.6151
R1612 B.n297 B.n296 10.6151
R1613 B.n297 B.n176 10.6151
R1614 B.n301 B.n176 10.6151
R1615 B.n302 B.n301 10.6151
R1616 B.n303 B.n302 10.6151
R1617 B.n303 B.n174 10.6151
R1618 B.n307 B.n174 10.6151
R1619 B.n308 B.n307 10.6151
R1620 B.n309 B.n308 10.6151
R1621 B.n309 B.n172 10.6151
R1622 B.n313 B.n172 10.6151
R1623 B.n314 B.n313 10.6151
R1624 B.n315 B.n314 10.6151
R1625 B.n315 B.n170 10.6151
R1626 B.n319 B.n170 10.6151
R1627 B.n320 B.n319 10.6151
R1628 B.n321 B.n320 10.6151
R1629 B.n321 B.n168 10.6151
R1630 B.n325 B.n168 10.6151
R1631 B.n326 B.n325 10.6151
R1632 B.n327 B.n166 10.6151
R1633 B.n331 B.n166 10.6151
R1634 B.n332 B.n331 10.6151
R1635 B.n333 B.n332 10.6151
R1636 B.n333 B.n164 10.6151
R1637 B.n337 B.n164 10.6151
R1638 B.n338 B.n337 10.6151
R1639 B.n339 B.n338 10.6151
R1640 B.n339 B.n162 10.6151
R1641 B.n343 B.n162 10.6151
R1642 B.n344 B.n343 10.6151
R1643 B.n348 B.n344 10.6151
R1644 B.n352 B.n160 10.6151
R1645 B.n353 B.n352 10.6151
R1646 B.n354 B.n353 10.6151
R1647 B.n354 B.n158 10.6151
R1648 B.n358 B.n158 10.6151
R1649 B.n359 B.n358 10.6151
R1650 B.n360 B.n359 10.6151
R1651 B.n360 B.n156 10.6151
R1652 B.n364 B.n156 10.6151
R1653 B.n367 B.n366 10.6151
R1654 B.n367 B.n152 10.6151
R1655 B.n371 B.n152 10.6151
R1656 B.n372 B.n371 10.6151
R1657 B.n373 B.n372 10.6151
R1658 B.n373 B.n150 10.6151
R1659 B.n377 B.n150 10.6151
R1660 B.n378 B.n377 10.6151
R1661 B.n379 B.n378 10.6151
R1662 B.n379 B.n148 10.6151
R1663 B.n383 B.n148 10.6151
R1664 B.n384 B.n383 10.6151
R1665 B.n667 B.n666 9.36635
R1666 B.n649 B.n58 9.36635
R1667 B.n348 B.n347 9.36635
R1668 B.n366 B.n365 9.36635
R1669 B.n809 B.n0 8.11757
R1670 B.n809 B.n1 8.11757
R1671 B.n666 B.n665 1.24928
R1672 B.n652 B.n58 1.24928
R1673 B.n347 B.n160 1.24928
R1674 B.n365 B.n364 1.24928
C0 w_n5962_n1420# B 9.96926f
C1 VP VN 8.4066f
C2 VTAIL VP 4.68204f
C3 VN VDD2 2.60131f
C4 VTAIL VDD2 7.3339f
C5 w_n5962_n1420# VP 13.754701f
C6 VTAIL VN 4.6678f
C7 w_n5962_n1420# VDD2 2.79011f
C8 w_n5962_n1420# VN 12.9784f
C9 w_n5962_n1420# VTAIL 2.03483f
C10 VDD1 B 2.16943f
C11 VDD1 VP 3.18183f
C12 VDD1 VDD2 2.97434f
C13 VDD1 VN 0.162481f
C14 VDD1 VTAIL 7.27224f
C15 w_n5962_n1420# VDD1 2.58331f
C16 VP B 2.82905f
C17 B VDD2 2.33568f
C18 B VN 1.51127f
C19 VTAIL B 1.74268f
C20 VP VDD2 0.747684f
C21 VDD2 VSUBS 2.602129f
C22 VDD1 VSUBS 2.315657f
C23 VTAIL VSUBS 0.750726f
C24 VN VSUBS 10.04651f
C25 VP VSUBS 5.047292f
C26 B VSUBS 5.680255f
C27 w_n5962_n1420# VSUBS 0.107817p
C28 B.n0 VSUBS 0.012446f
C29 B.n1 VSUBS 0.012446f
C30 B.n2 VSUBS 0.018408f
C31 B.n3 VSUBS 0.014106f
C32 B.n4 VSUBS 0.014106f
C33 B.n5 VSUBS 0.014106f
C34 B.n6 VSUBS 0.014106f
C35 B.n7 VSUBS 0.014106f
C36 B.n8 VSUBS 0.014106f
C37 B.n9 VSUBS 0.014106f
C38 B.n10 VSUBS 0.014106f
C39 B.n11 VSUBS 0.014106f
C40 B.n12 VSUBS 0.014106f
C41 B.n13 VSUBS 0.014106f
C42 B.n14 VSUBS 0.014106f
C43 B.n15 VSUBS 0.014106f
C44 B.n16 VSUBS 0.014106f
C45 B.n17 VSUBS 0.014106f
C46 B.n18 VSUBS 0.014106f
C47 B.n19 VSUBS 0.014106f
C48 B.n20 VSUBS 0.014106f
C49 B.n21 VSUBS 0.014106f
C50 B.n22 VSUBS 0.014106f
C51 B.n23 VSUBS 0.014106f
C52 B.n24 VSUBS 0.014106f
C53 B.n25 VSUBS 0.014106f
C54 B.n26 VSUBS 0.014106f
C55 B.n27 VSUBS 0.014106f
C56 B.n28 VSUBS 0.014106f
C57 B.n29 VSUBS 0.014106f
C58 B.n30 VSUBS 0.014106f
C59 B.n31 VSUBS 0.014106f
C60 B.n32 VSUBS 0.014106f
C61 B.n33 VSUBS 0.014106f
C62 B.n34 VSUBS 0.014106f
C63 B.n35 VSUBS 0.014106f
C64 B.n36 VSUBS 0.014106f
C65 B.n37 VSUBS 0.014106f
C66 B.n38 VSUBS 0.014106f
C67 B.n39 VSUBS 0.014106f
C68 B.n40 VSUBS 0.014106f
C69 B.n41 VSUBS 0.014106f
C70 B.n42 VSUBS 0.030068f
C71 B.n43 VSUBS 0.014106f
C72 B.n44 VSUBS 0.014106f
C73 B.n45 VSUBS 0.014106f
C74 B.n46 VSUBS 0.014106f
C75 B.n47 VSUBS 0.014106f
C76 B.n48 VSUBS 0.014106f
C77 B.n49 VSUBS 0.014106f
C78 B.t1 VSUBS 0.100921f
C79 B.t2 VSUBS 0.136557f
C80 B.t0 VSUBS 0.86151f
C81 B.n50 VSUBS 0.171543f
C82 B.n51 VSUBS 0.132443f
C83 B.n52 VSUBS 0.014106f
C84 B.n53 VSUBS 0.014106f
C85 B.n54 VSUBS 0.014106f
C86 B.n55 VSUBS 0.014106f
C87 B.t10 VSUBS 0.100921f
C88 B.t11 VSUBS 0.136557f
C89 B.t9 VSUBS 0.86151f
C90 B.n56 VSUBS 0.171543f
C91 B.n57 VSUBS 0.132443f
C92 B.n58 VSUBS 0.032682f
C93 B.n59 VSUBS 0.014106f
C94 B.n60 VSUBS 0.014106f
C95 B.n61 VSUBS 0.014106f
C96 B.n62 VSUBS 0.014106f
C97 B.n63 VSUBS 0.014106f
C98 B.n64 VSUBS 0.014106f
C99 B.n65 VSUBS 0.030068f
C100 B.n66 VSUBS 0.014106f
C101 B.n67 VSUBS 0.014106f
C102 B.n68 VSUBS 0.014106f
C103 B.n69 VSUBS 0.014106f
C104 B.n70 VSUBS 0.014106f
C105 B.n71 VSUBS 0.014106f
C106 B.n72 VSUBS 0.014106f
C107 B.n73 VSUBS 0.014106f
C108 B.n74 VSUBS 0.014106f
C109 B.n75 VSUBS 0.014106f
C110 B.n76 VSUBS 0.014106f
C111 B.n77 VSUBS 0.014106f
C112 B.n78 VSUBS 0.014106f
C113 B.n79 VSUBS 0.014106f
C114 B.n80 VSUBS 0.014106f
C115 B.n81 VSUBS 0.014106f
C116 B.n82 VSUBS 0.014106f
C117 B.n83 VSUBS 0.014106f
C118 B.n84 VSUBS 0.014106f
C119 B.n85 VSUBS 0.014106f
C120 B.n86 VSUBS 0.014106f
C121 B.n87 VSUBS 0.014106f
C122 B.n88 VSUBS 0.014106f
C123 B.n89 VSUBS 0.014106f
C124 B.n90 VSUBS 0.014106f
C125 B.n91 VSUBS 0.014106f
C126 B.n92 VSUBS 0.014106f
C127 B.n93 VSUBS 0.014106f
C128 B.n94 VSUBS 0.014106f
C129 B.n95 VSUBS 0.014106f
C130 B.n96 VSUBS 0.014106f
C131 B.n97 VSUBS 0.014106f
C132 B.n98 VSUBS 0.014106f
C133 B.n99 VSUBS 0.014106f
C134 B.n100 VSUBS 0.014106f
C135 B.n101 VSUBS 0.014106f
C136 B.n102 VSUBS 0.014106f
C137 B.n103 VSUBS 0.014106f
C138 B.n104 VSUBS 0.014106f
C139 B.n105 VSUBS 0.014106f
C140 B.n106 VSUBS 0.014106f
C141 B.n107 VSUBS 0.014106f
C142 B.n108 VSUBS 0.014106f
C143 B.n109 VSUBS 0.014106f
C144 B.n110 VSUBS 0.014106f
C145 B.n111 VSUBS 0.014106f
C146 B.n112 VSUBS 0.014106f
C147 B.n113 VSUBS 0.014106f
C148 B.n114 VSUBS 0.014106f
C149 B.n115 VSUBS 0.014106f
C150 B.n116 VSUBS 0.014106f
C151 B.n117 VSUBS 0.014106f
C152 B.n118 VSUBS 0.014106f
C153 B.n119 VSUBS 0.014106f
C154 B.n120 VSUBS 0.014106f
C155 B.n121 VSUBS 0.014106f
C156 B.n122 VSUBS 0.014106f
C157 B.n123 VSUBS 0.014106f
C158 B.n124 VSUBS 0.014106f
C159 B.n125 VSUBS 0.014106f
C160 B.n126 VSUBS 0.014106f
C161 B.n127 VSUBS 0.014106f
C162 B.n128 VSUBS 0.014106f
C163 B.n129 VSUBS 0.014106f
C164 B.n130 VSUBS 0.014106f
C165 B.n131 VSUBS 0.014106f
C166 B.n132 VSUBS 0.014106f
C167 B.n133 VSUBS 0.014106f
C168 B.n134 VSUBS 0.014106f
C169 B.n135 VSUBS 0.014106f
C170 B.n136 VSUBS 0.014106f
C171 B.n137 VSUBS 0.014106f
C172 B.n138 VSUBS 0.014106f
C173 B.n139 VSUBS 0.014106f
C174 B.n140 VSUBS 0.014106f
C175 B.n141 VSUBS 0.014106f
C176 B.n142 VSUBS 0.014106f
C177 B.n143 VSUBS 0.014106f
C178 B.n144 VSUBS 0.014106f
C179 B.n145 VSUBS 0.014106f
C180 B.n146 VSUBS 0.014106f
C181 B.n147 VSUBS 0.03258f
C182 B.n148 VSUBS 0.014106f
C183 B.n149 VSUBS 0.014106f
C184 B.n150 VSUBS 0.014106f
C185 B.n151 VSUBS 0.014106f
C186 B.n152 VSUBS 0.014106f
C187 B.n153 VSUBS 0.014106f
C188 B.t8 VSUBS 0.100921f
C189 B.t7 VSUBS 0.136557f
C190 B.t6 VSUBS 0.86151f
C191 B.n154 VSUBS 0.171543f
C192 B.n155 VSUBS 0.132443f
C193 B.n156 VSUBS 0.014106f
C194 B.n157 VSUBS 0.014106f
C195 B.n158 VSUBS 0.014106f
C196 B.n159 VSUBS 0.014106f
C197 B.n160 VSUBS 0.007883f
C198 B.n161 VSUBS 0.014106f
C199 B.n162 VSUBS 0.014106f
C200 B.n163 VSUBS 0.014106f
C201 B.n164 VSUBS 0.014106f
C202 B.n165 VSUBS 0.014106f
C203 B.n166 VSUBS 0.014106f
C204 B.n167 VSUBS 0.030068f
C205 B.n168 VSUBS 0.014106f
C206 B.n169 VSUBS 0.014106f
C207 B.n170 VSUBS 0.014106f
C208 B.n171 VSUBS 0.014106f
C209 B.n172 VSUBS 0.014106f
C210 B.n173 VSUBS 0.014106f
C211 B.n174 VSUBS 0.014106f
C212 B.n175 VSUBS 0.014106f
C213 B.n176 VSUBS 0.014106f
C214 B.n177 VSUBS 0.014106f
C215 B.n178 VSUBS 0.014106f
C216 B.n179 VSUBS 0.014106f
C217 B.n180 VSUBS 0.014106f
C218 B.n181 VSUBS 0.014106f
C219 B.n182 VSUBS 0.014106f
C220 B.n183 VSUBS 0.014106f
C221 B.n184 VSUBS 0.014106f
C222 B.n185 VSUBS 0.014106f
C223 B.n186 VSUBS 0.014106f
C224 B.n187 VSUBS 0.014106f
C225 B.n188 VSUBS 0.014106f
C226 B.n189 VSUBS 0.014106f
C227 B.n190 VSUBS 0.014106f
C228 B.n191 VSUBS 0.014106f
C229 B.n192 VSUBS 0.014106f
C230 B.n193 VSUBS 0.014106f
C231 B.n194 VSUBS 0.014106f
C232 B.n195 VSUBS 0.014106f
C233 B.n196 VSUBS 0.014106f
C234 B.n197 VSUBS 0.014106f
C235 B.n198 VSUBS 0.014106f
C236 B.n199 VSUBS 0.014106f
C237 B.n200 VSUBS 0.014106f
C238 B.n201 VSUBS 0.014106f
C239 B.n202 VSUBS 0.014106f
C240 B.n203 VSUBS 0.014106f
C241 B.n204 VSUBS 0.014106f
C242 B.n205 VSUBS 0.014106f
C243 B.n206 VSUBS 0.014106f
C244 B.n207 VSUBS 0.014106f
C245 B.n208 VSUBS 0.014106f
C246 B.n209 VSUBS 0.014106f
C247 B.n210 VSUBS 0.014106f
C248 B.n211 VSUBS 0.014106f
C249 B.n212 VSUBS 0.014106f
C250 B.n213 VSUBS 0.014106f
C251 B.n214 VSUBS 0.014106f
C252 B.n215 VSUBS 0.014106f
C253 B.n216 VSUBS 0.014106f
C254 B.n217 VSUBS 0.014106f
C255 B.n218 VSUBS 0.014106f
C256 B.n219 VSUBS 0.014106f
C257 B.n220 VSUBS 0.014106f
C258 B.n221 VSUBS 0.014106f
C259 B.n222 VSUBS 0.014106f
C260 B.n223 VSUBS 0.014106f
C261 B.n224 VSUBS 0.014106f
C262 B.n225 VSUBS 0.014106f
C263 B.n226 VSUBS 0.014106f
C264 B.n227 VSUBS 0.014106f
C265 B.n228 VSUBS 0.014106f
C266 B.n229 VSUBS 0.014106f
C267 B.n230 VSUBS 0.014106f
C268 B.n231 VSUBS 0.014106f
C269 B.n232 VSUBS 0.014106f
C270 B.n233 VSUBS 0.014106f
C271 B.n234 VSUBS 0.014106f
C272 B.n235 VSUBS 0.014106f
C273 B.n236 VSUBS 0.014106f
C274 B.n237 VSUBS 0.014106f
C275 B.n238 VSUBS 0.014106f
C276 B.n239 VSUBS 0.014106f
C277 B.n240 VSUBS 0.014106f
C278 B.n241 VSUBS 0.014106f
C279 B.n242 VSUBS 0.014106f
C280 B.n243 VSUBS 0.014106f
C281 B.n244 VSUBS 0.014106f
C282 B.n245 VSUBS 0.014106f
C283 B.n246 VSUBS 0.014106f
C284 B.n247 VSUBS 0.014106f
C285 B.n248 VSUBS 0.014106f
C286 B.n249 VSUBS 0.014106f
C287 B.n250 VSUBS 0.014106f
C288 B.n251 VSUBS 0.014106f
C289 B.n252 VSUBS 0.014106f
C290 B.n253 VSUBS 0.014106f
C291 B.n254 VSUBS 0.014106f
C292 B.n255 VSUBS 0.014106f
C293 B.n256 VSUBS 0.014106f
C294 B.n257 VSUBS 0.014106f
C295 B.n258 VSUBS 0.014106f
C296 B.n259 VSUBS 0.014106f
C297 B.n260 VSUBS 0.014106f
C298 B.n261 VSUBS 0.014106f
C299 B.n262 VSUBS 0.014106f
C300 B.n263 VSUBS 0.014106f
C301 B.n264 VSUBS 0.014106f
C302 B.n265 VSUBS 0.014106f
C303 B.n266 VSUBS 0.014106f
C304 B.n267 VSUBS 0.014106f
C305 B.n268 VSUBS 0.014106f
C306 B.n269 VSUBS 0.014106f
C307 B.n270 VSUBS 0.014106f
C308 B.n271 VSUBS 0.014106f
C309 B.n272 VSUBS 0.014106f
C310 B.n273 VSUBS 0.014106f
C311 B.n274 VSUBS 0.014106f
C312 B.n275 VSUBS 0.014106f
C313 B.n276 VSUBS 0.014106f
C314 B.n277 VSUBS 0.014106f
C315 B.n278 VSUBS 0.014106f
C316 B.n279 VSUBS 0.014106f
C317 B.n280 VSUBS 0.014106f
C318 B.n281 VSUBS 0.014106f
C319 B.n282 VSUBS 0.014106f
C320 B.n283 VSUBS 0.014106f
C321 B.n284 VSUBS 0.014106f
C322 B.n285 VSUBS 0.014106f
C323 B.n286 VSUBS 0.014106f
C324 B.n287 VSUBS 0.014106f
C325 B.n288 VSUBS 0.014106f
C326 B.n289 VSUBS 0.014106f
C327 B.n290 VSUBS 0.014106f
C328 B.n291 VSUBS 0.014106f
C329 B.n292 VSUBS 0.014106f
C330 B.n293 VSUBS 0.014106f
C331 B.n294 VSUBS 0.014106f
C332 B.n295 VSUBS 0.014106f
C333 B.n296 VSUBS 0.014106f
C334 B.n297 VSUBS 0.014106f
C335 B.n298 VSUBS 0.014106f
C336 B.n299 VSUBS 0.014106f
C337 B.n300 VSUBS 0.014106f
C338 B.n301 VSUBS 0.014106f
C339 B.n302 VSUBS 0.014106f
C340 B.n303 VSUBS 0.014106f
C341 B.n304 VSUBS 0.014106f
C342 B.n305 VSUBS 0.014106f
C343 B.n306 VSUBS 0.014106f
C344 B.n307 VSUBS 0.014106f
C345 B.n308 VSUBS 0.014106f
C346 B.n309 VSUBS 0.014106f
C347 B.n310 VSUBS 0.014106f
C348 B.n311 VSUBS 0.014106f
C349 B.n312 VSUBS 0.014106f
C350 B.n313 VSUBS 0.014106f
C351 B.n314 VSUBS 0.014106f
C352 B.n315 VSUBS 0.014106f
C353 B.n316 VSUBS 0.014106f
C354 B.n317 VSUBS 0.014106f
C355 B.n318 VSUBS 0.014106f
C356 B.n319 VSUBS 0.014106f
C357 B.n320 VSUBS 0.014106f
C358 B.n321 VSUBS 0.014106f
C359 B.n322 VSUBS 0.014106f
C360 B.n323 VSUBS 0.014106f
C361 B.n324 VSUBS 0.014106f
C362 B.n325 VSUBS 0.014106f
C363 B.n326 VSUBS 0.030068f
C364 B.n327 VSUBS 0.03258f
C365 B.n328 VSUBS 0.03258f
C366 B.n329 VSUBS 0.014106f
C367 B.n330 VSUBS 0.014106f
C368 B.n331 VSUBS 0.014106f
C369 B.n332 VSUBS 0.014106f
C370 B.n333 VSUBS 0.014106f
C371 B.n334 VSUBS 0.014106f
C372 B.n335 VSUBS 0.014106f
C373 B.n336 VSUBS 0.014106f
C374 B.n337 VSUBS 0.014106f
C375 B.n338 VSUBS 0.014106f
C376 B.n339 VSUBS 0.014106f
C377 B.n340 VSUBS 0.014106f
C378 B.n341 VSUBS 0.014106f
C379 B.n342 VSUBS 0.014106f
C380 B.n343 VSUBS 0.014106f
C381 B.n344 VSUBS 0.014106f
C382 B.t5 VSUBS 0.100921f
C383 B.t4 VSUBS 0.136557f
C384 B.t3 VSUBS 0.86151f
C385 B.n345 VSUBS 0.171543f
C386 B.n346 VSUBS 0.132443f
C387 B.n347 VSUBS 0.032682f
C388 B.n348 VSUBS 0.013276f
C389 B.n349 VSUBS 0.014106f
C390 B.n350 VSUBS 0.014106f
C391 B.n351 VSUBS 0.014106f
C392 B.n352 VSUBS 0.014106f
C393 B.n353 VSUBS 0.014106f
C394 B.n354 VSUBS 0.014106f
C395 B.n355 VSUBS 0.014106f
C396 B.n356 VSUBS 0.014106f
C397 B.n357 VSUBS 0.014106f
C398 B.n358 VSUBS 0.014106f
C399 B.n359 VSUBS 0.014106f
C400 B.n360 VSUBS 0.014106f
C401 B.n361 VSUBS 0.014106f
C402 B.n362 VSUBS 0.014106f
C403 B.n363 VSUBS 0.014106f
C404 B.n364 VSUBS 0.007883f
C405 B.n365 VSUBS 0.032682f
C406 B.n366 VSUBS 0.013276f
C407 B.n367 VSUBS 0.014106f
C408 B.n368 VSUBS 0.014106f
C409 B.n369 VSUBS 0.014106f
C410 B.n370 VSUBS 0.014106f
C411 B.n371 VSUBS 0.014106f
C412 B.n372 VSUBS 0.014106f
C413 B.n373 VSUBS 0.014106f
C414 B.n374 VSUBS 0.014106f
C415 B.n375 VSUBS 0.014106f
C416 B.n376 VSUBS 0.014106f
C417 B.n377 VSUBS 0.014106f
C418 B.n378 VSUBS 0.014106f
C419 B.n379 VSUBS 0.014106f
C420 B.n380 VSUBS 0.014106f
C421 B.n381 VSUBS 0.014106f
C422 B.n382 VSUBS 0.014106f
C423 B.n383 VSUBS 0.014106f
C424 B.n384 VSUBS 0.030773f
C425 B.n385 VSUBS 0.031875f
C426 B.n386 VSUBS 0.030068f
C427 B.n387 VSUBS 0.014106f
C428 B.n388 VSUBS 0.014106f
C429 B.n389 VSUBS 0.014106f
C430 B.n390 VSUBS 0.014106f
C431 B.n391 VSUBS 0.014106f
C432 B.n392 VSUBS 0.014106f
C433 B.n393 VSUBS 0.014106f
C434 B.n394 VSUBS 0.014106f
C435 B.n395 VSUBS 0.014106f
C436 B.n396 VSUBS 0.014106f
C437 B.n397 VSUBS 0.014106f
C438 B.n398 VSUBS 0.014106f
C439 B.n399 VSUBS 0.014106f
C440 B.n400 VSUBS 0.014106f
C441 B.n401 VSUBS 0.014106f
C442 B.n402 VSUBS 0.014106f
C443 B.n403 VSUBS 0.014106f
C444 B.n404 VSUBS 0.014106f
C445 B.n405 VSUBS 0.014106f
C446 B.n406 VSUBS 0.014106f
C447 B.n407 VSUBS 0.014106f
C448 B.n408 VSUBS 0.014106f
C449 B.n409 VSUBS 0.014106f
C450 B.n410 VSUBS 0.014106f
C451 B.n411 VSUBS 0.014106f
C452 B.n412 VSUBS 0.014106f
C453 B.n413 VSUBS 0.014106f
C454 B.n414 VSUBS 0.014106f
C455 B.n415 VSUBS 0.014106f
C456 B.n416 VSUBS 0.014106f
C457 B.n417 VSUBS 0.014106f
C458 B.n418 VSUBS 0.014106f
C459 B.n419 VSUBS 0.014106f
C460 B.n420 VSUBS 0.014106f
C461 B.n421 VSUBS 0.014106f
C462 B.n422 VSUBS 0.014106f
C463 B.n423 VSUBS 0.014106f
C464 B.n424 VSUBS 0.014106f
C465 B.n425 VSUBS 0.014106f
C466 B.n426 VSUBS 0.014106f
C467 B.n427 VSUBS 0.014106f
C468 B.n428 VSUBS 0.014106f
C469 B.n429 VSUBS 0.014106f
C470 B.n430 VSUBS 0.014106f
C471 B.n431 VSUBS 0.014106f
C472 B.n432 VSUBS 0.014106f
C473 B.n433 VSUBS 0.014106f
C474 B.n434 VSUBS 0.014106f
C475 B.n435 VSUBS 0.014106f
C476 B.n436 VSUBS 0.014106f
C477 B.n437 VSUBS 0.014106f
C478 B.n438 VSUBS 0.014106f
C479 B.n439 VSUBS 0.014106f
C480 B.n440 VSUBS 0.014106f
C481 B.n441 VSUBS 0.014106f
C482 B.n442 VSUBS 0.014106f
C483 B.n443 VSUBS 0.014106f
C484 B.n444 VSUBS 0.014106f
C485 B.n445 VSUBS 0.014106f
C486 B.n446 VSUBS 0.014106f
C487 B.n447 VSUBS 0.014106f
C488 B.n448 VSUBS 0.014106f
C489 B.n449 VSUBS 0.014106f
C490 B.n450 VSUBS 0.014106f
C491 B.n451 VSUBS 0.014106f
C492 B.n452 VSUBS 0.014106f
C493 B.n453 VSUBS 0.014106f
C494 B.n454 VSUBS 0.014106f
C495 B.n455 VSUBS 0.014106f
C496 B.n456 VSUBS 0.014106f
C497 B.n457 VSUBS 0.014106f
C498 B.n458 VSUBS 0.014106f
C499 B.n459 VSUBS 0.014106f
C500 B.n460 VSUBS 0.014106f
C501 B.n461 VSUBS 0.014106f
C502 B.n462 VSUBS 0.014106f
C503 B.n463 VSUBS 0.014106f
C504 B.n464 VSUBS 0.014106f
C505 B.n465 VSUBS 0.014106f
C506 B.n466 VSUBS 0.014106f
C507 B.n467 VSUBS 0.014106f
C508 B.n468 VSUBS 0.014106f
C509 B.n469 VSUBS 0.014106f
C510 B.n470 VSUBS 0.014106f
C511 B.n471 VSUBS 0.014106f
C512 B.n472 VSUBS 0.014106f
C513 B.n473 VSUBS 0.014106f
C514 B.n474 VSUBS 0.014106f
C515 B.n475 VSUBS 0.014106f
C516 B.n476 VSUBS 0.014106f
C517 B.n477 VSUBS 0.014106f
C518 B.n478 VSUBS 0.014106f
C519 B.n479 VSUBS 0.014106f
C520 B.n480 VSUBS 0.014106f
C521 B.n481 VSUBS 0.014106f
C522 B.n482 VSUBS 0.014106f
C523 B.n483 VSUBS 0.014106f
C524 B.n484 VSUBS 0.014106f
C525 B.n485 VSUBS 0.014106f
C526 B.n486 VSUBS 0.014106f
C527 B.n487 VSUBS 0.014106f
C528 B.n488 VSUBS 0.014106f
C529 B.n489 VSUBS 0.014106f
C530 B.n490 VSUBS 0.014106f
C531 B.n491 VSUBS 0.014106f
C532 B.n492 VSUBS 0.014106f
C533 B.n493 VSUBS 0.014106f
C534 B.n494 VSUBS 0.014106f
C535 B.n495 VSUBS 0.014106f
C536 B.n496 VSUBS 0.014106f
C537 B.n497 VSUBS 0.014106f
C538 B.n498 VSUBS 0.014106f
C539 B.n499 VSUBS 0.014106f
C540 B.n500 VSUBS 0.014106f
C541 B.n501 VSUBS 0.014106f
C542 B.n502 VSUBS 0.014106f
C543 B.n503 VSUBS 0.014106f
C544 B.n504 VSUBS 0.014106f
C545 B.n505 VSUBS 0.014106f
C546 B.n506 VSUBS 0.014106f
C547 B.n507 VSUBS 0.014106f
C548 B.n508 VSUBS 0.014106f
C549 B.n509 VSUBS 0.014106f
C550 B.n510 VSUBS 0.014106f
C551 B.n511 VSUBS 0.014106f
C552 B.n512 VSUBS 0.014106f
C553 B.n513 VSUBS 0.014106f
C554 B.n514 VSUBS 0.014106f
C555 B.n515 VSUBS 0.014106f
C556 B.n516 VSUBS 0.014106f
C557 B.n517 VSUBS 0.014106f
C558 B.n518 VSUBS 0.014106f
C559 B.n519 VSUBS 0.014106f
C560 B.n520 VSUBS 0.014106f
C561 B.n521 VSUBS 0.014106f
C562 B.n522 VSUBS 0.014106f
C563 B.n523 VSUBS 0.014106f
C564 B.n524 VSUBS 0.014106f
C565 B.n525 VSUBS 0.014106f
C566 B.n526 VSUBS 0.014106f
C567 B.n527 VSUBS 0.014106f
C568 B.n528 VSUBS 0.014106f
C569 B.n529 VSUBS 0.014106f
C570 B.n530 VSUBS 0.014106f
C571 B.n531 VSUBS 0.014106f
C572 B.n532 VSUBS 0.014106f
C573 B.n533 VSUBS 0.014106f
C574 B.n534 VSUBS 0.014106f
C575 B.n535 VSUBS 0.014106f
C576 B.n536 VSUBS 0.014106f
C577 B.n537 VSUBS 0.014106f
C578 B.n538 VSUBS 0.014106f
C579 B.n539 VSUBS 0.014106f
C580 B.n540 VSUBS 0.014106f
C581 B.n541 VSUBS 0.014106f
C582 B.n542 VSUBS 0.014106f
C583 B.n543 VSUBS 0.014106f
C584 B.n544 VSUBS 0.014106f
C585 B.n545 VSUBS 0.014106f
C586 B.n546 VSUBS 0.014106f
C587 B.n547 VSUBS 0.014106f
C588 B.n548 VSUBS 0.014106f
C589 B.n549 VSUBS 0.014106f
C590 B.n550 VSUBS 0.014106f
C591 B.n551 VSUBS 0.014106f
C592 B.n552 VSUBS 0.014106f
C593 B.n553 VSUBS 0.014106f
C594 B.n554 VSUBS 0.014106f
C595 B.n555 VSUBS 0.014106f
C596 B.n556 VSUBS 0.014106f
C597 B.n557 VSUBS 0.014106f
C598 B.n558 VSUBS 0.014106f
C599 B.n559 VSUBS 0.014106f
C600 B.n560 VSUBS 0.014106f
C601 B.n561 VSUBS 0.014106f
C602 B.n562 VSUBS 0.014106f
C603 B.n563 VSUBS 0.014106f
C604 B.n564 VSUBS 0.014106f
C605 B.n565 VSUBS 0.014106f
C606 B.n566 VSUBS 0.014106f
C607 B.n567 VSUBS 0.014106f
C608 B.n568 VSUBS 0.014106f
C609 B.n569 VSUBS 0.014106f
C610 B.n570 VSUBS 0.014106f
C611 B.n571 VSUBS 0.014106f
C612 B.n572 VSUBS 0.014106f
C613 B.n573 VSUBS 0.014106f
C614 B.n574 VSUBS 0.014106f
C615 B.n575 VSUBS 0.014106f
C616 B.n576 VSUBS 0.014106f
C617 B.n577 VSUBS 0.014106f
C618 B.n578 VSUBS 0.014106f
C619 B.n579 VSUBS 0.014106f
C620 B.n580 VSUBS 0.014106f
C621 B.n581 VSUBS 0.014106f
C622 B.n582 VSUBS 0.014106f
C623 B.n583 VSUBS 0.014106f
C624 B.n584 VSUBS 0.014106f
C625 B.n585 VSUBS 0.014106f
C626 B.n586 VSUBS 0.014106f
C627 B.n587 VSUBS 0.014106f
C628 B.n588 VSUBS 0.014106f
C629 B.n589 VSUBS 0.014106f
C630 B.n590 VSUBS 0.014106f
C631 B.n591 VSUBS 0.014106f
C632 B.n592 VSUBS 0.014106f
C633 B.n593 VSUBS 0.014106f
C634 B.n594 VSUBS 0.014106f
C635 B.n595 VSUBS 0.014106f
C636 B.n596 VSUBS 0.014106f
C637 B.n597 VSUBS 0.014106f
C638 B.n598 VSUBS 0.014106f
C639 B.n599 VSUBS 0.014106f
C640 B.n600 VSUBS 0.014106f
C641 B.n601 VSUBS 0.014106f
C642 B.n602 VSUBS 0.014106f
C643 B.n603 VSUBS 0.014106f
C644 B.n604 VSUBS 0.014106f
C645 B.n605 VSUBS 0.014106f
C646 B.n606 VSUBS 0.014106f
C647 B.n607 VSUBS 0.014106f
C648 B.n608 VSUBS 0.014106f
C649 B.n609 VSUBS 0.014106f
C650 B.n610 VSUBS 0.014106f
C651 B.n611 VSUBS 0.014106f
C652 B.n612 VSUBS 0.014106f
C653 B.n613 VSUBS 0.014106f
C654 B.n614 VSUBS 0.014106f
C655 B.n615 VSUBS 0.014106f
C656 B.n616 VSUBS 0.014106f
C657 B.n617 VSUBS 0.014106f
C658 B.n618 VSUBS 0.014106f
C659 B.n619 VSUBS 0.014106f
C660 B.n620 VSUBS 0.014106f
C661 B.n621 VSUBS 0.014106f
C662 B.n622 VSUBS 0.014106f
C663 B.n623 VSUBS 0.014106f
C664 B.n624 VSUBS 0.014106f
C665 B.n625 VSUBS 0.014106f
C666 B.n626 VSUBS 0.014106f
C667 B.n627 VSUBS 0.014106f
C668 B.n628 VSUBS 0.014106f
C669 B.n629 VSUBS 0.014106f
C670 B.n630 VSUBS 0.030068f
C671 B.n631 VSUBS 0.03258f
C672 B.n632 VSUBS 0.03258f
C673 B.n633 VSUBS 0.014106f
C674 B.n634 VSUBS 0.014106f
C675 B.n635 VSUBS 0.014106f
C676 B.n636 VSUBS 0.014106f
C677 B.n637 VSUBS 0.014106f
C678 B.n638 VSUBS 0.014106f
C679 B.n639 VSUBS 0.014106f
C680 B.n640 VSUBS 0.014106f
C681 B.n641 VSUBS 0.014106f
C682 B.n642 VSUBS 0.014106f
C683 B.n643 VSUBS 0.014106f
C684 B.n644 VSUBS 0.014106f
C685 B.n645 VSUBS 0.014106f
C686 B.n646 VSUBS 0.014106f
C687 B.n647 VSUBS 0.014106f
C688 B.n648 VSUBS 0.014106f
C689 B.n649 VSUBS 0.013276f
C690 B.n650 VSUBS 0.014106f
C691 B.n651 VSUBS 0.014106f
C692 B.n652 VSUBS 0.007883f
C693 B.n653 VSUBS 0.014106f
C694 B.n654 VSUBS 0.014106f
C695 B.n655 VSUBS 0.014106f
C696 B.n656 VSUBS 0.014106f
C697 B.n657 VSUBS 0.014106f
C698 B.n658 VSUBS 0.014106f
C699 B.n659 VSUBS 0.014106f
C700 B.n660 VSUBS 0.014106f
C701 B.n661 VSUBS 0.014106f
C702 B.n662 VSUBS 0.014106f
C703 B.n663 VSUBS 0.014106f
C704 B.n664 VSUBS 0.014106f
C705 B.n665 VSUBS 0.007883f
C706 B.n666 VSUBS 0.032682f
C707 B.n667 VSUBS 0.013276f
C708 B.n668 VSUBS 0.014106f
C709 B.n669 VSUBS 0.014106f
C710 B.n670 VSUBS 0.014106f
C711 B.n671 VSUBS 0.014106f
C712 B.n672 VSUBS 0.014106f
C713 B.n673 VSUBS 0.014106f
C714 B.n674 VSUBS 0.014106f
C715 B.n675 VSUBS 0.014106f
C716 B.n676 VSUBS 0.014106f
C717 B.n677 VSUBS 0.014106f
C718 B.n678 VSUBS 0.014106f
C719 B.n679 VSUBS 0.014106f
C720 B.n680 VSUBS 0.014106f
C721 B.n681 VSUBS 0.014106f
C722 B.n682 VSUBS 0.014106f
C723 B.n683 VSUBS 0.014106f
C724 B.n684 VSUBS 0.014106f
C725 B.n685 VSUBS 0.03258f
C726 B.n686 VSUBS 0.03258f
C727 B.n687 VSUBS 0.030068f
C728 B.n688 VSUBS 0.014106f
C729 B.n689 VSUBS 0.014106f
C730 B.n690 VSUBS 0.014106f
C731 B.n691 VSUBS 0.014106f
C732 B.n692 VSUBS 0.014106f
C733 B.n693 VSUBS 0.014106f
C734 B.n694 VSUBS 0.014106f
C735 B.n695 VSUBS 0.014106f
C736 B.n696 VSUBS 0.014106f
C737 B.n697 VSUBS 0.014106f
C738 B.n698 VSUBS 0.014106f
C739 B.n699 VSUBS 0.014106f
C740 B.n700 VSUBS 0.014106f
C741 B.n701 VSUBS 0.014106f
C742 B.n702 VSUBS 0.014106f
C743 B.n703 VSUBS 0.014106f
C744 B.n704 VSUBS 0.014106f
C745 B.n705 VSUBS 0.014106f
C746 B.n706 VSUBS 0.014106f
C747 B.n707 VSUBS 0.014106f
C748 B.n708 VSUBS 0.014106f
C749 B.n709 VSUBS 0.014106f
C750 B.n710 VSUBS 0.014106f
C751 B.n711 VSUBS 0.014106f
C752 B.n712 VSUBS 0.014106f
C753 B.n713 VSUBS 0.014106f
C754 B.n714 VSUBS 0.014106f
C755 B.n715 VSUBS 0.014106f
C756 B.n716 VSUBS 0.014106f
C757 B.n717 VSUBS 0.014106f
C758 B.n718 VSUBS 0.014106f
C759 B.n719 VSUBS 0.014106f
C760 B.n720 VSUBS 0.014106f
C761 B.n721 VSUBS 0.014106f
C762 B.n722 VSUBS 0.014106f
C763 B.n723 VSUBS 0.014106f
C764 B.n724 VSUBS 0.014106f
C765 B.n725 VSUBS 0.014106f
C766 B.n726 VSUBS 0.014106f
C767 B.n727 VSUBS 0.014106f
C768 B.n728 VSUBS 0.014106f
C769 B.n729 VSUBS 0.014106f
C770 B.n730 VSUBS 0.014106f
C771 B.n731 VSUBS 0.014106f
C772 B.n732 VSUBS 0.014106f
C773 B.n733 VSUBS 0.014106f
C774 B.n734 VSUBS 0.014106f
C775 B.n735 VSUBS 0.014106f
C776 B.n736 VSUBS 0.014106f
C777 B.n737 VSUBS 0.014106f
C778 B.n738 VSUBS 0.014106f
C779 B.n739 VSUBS 0.014106f
C780 B.n740 VSUBS 0.014106f
C781 B.n741 VSUBS 0.014106f
C782 B.n742 VSUBS 0.014106f
C783 B.n743 VSUBS 0.014106f
C784 B.n744 VSUBS 0.014106f
C785 B.n745 VSUBS 0.014106f
C786 B.n746 VSUBS 0.014106f
C787 B.n747 VSUBS 0.014106f
C788 B.n748 VSUBS 0.014106f
C789 B.n749 VSUBS 0.014106f
C790 B.n750 VSUBS 0.014106f
C791 B.n751 VSUBS 0.014106f
C792 B.n752 VSUBS 0.014106f
C793 B.n753 VSUBS 0.014106f
C794 B.n754 VSUBS 0.014106f
C795 B.n755 VSUBS 0.014106f
C796 B.n756 VSUBS 0.014106f
C797 B.n757 VSUBS 0.014106f
C798 B.n758 VSUBS 0.014106f
C799 B.n759 VSUBS 0.014106f
C800 B.n760 VSUBS 0.014106f
C801 B.n761 VSUBS 0.014106f
C802 B.n762 VSUBS 0.014106f
C803 B.n763 VSUBS 0.014106f
C804 B.n764 VSUBS 0.014106f
C805 B.n765 VSUBS 0.014106f
C806 B.n766 VSUBS 0.014106f
C807 B.n767 VSUBS 0.014106f
C808 B.n768 VSUBS 0.014106f
C809 B.n769 VSUBS 0.014106f
C810 B.n770 VSUBS 0.014106f
C811 B.n771 VSUBS 0.014106f
C812 B.n772 VSUBS 0.014106f
C813 B.n773 VSUBS 0.014106f
C814 B.n774 VSUBS 0.014106f
C815 B.n775 VSUBS 0.014106f
C816 B.n776 VSUBS 0.014106f
C817 B.n777 VSUBS 0.014106f
C818 B.n778 VSUBS 0.014106f
C819 B.n779 VSUBS 0.014106f
C820 B.n780 VSUBS 0.014106f
C821 B.n781 VSUBS 0.014106f
C822 B.n782 VSUBS 0.014106f
C823 B.n783 VSUBS 0.014106f
C824 B.n784 VSUBS 0.014106f
C825 B.n785 VSUBS 0.014106f
C826 B.n786 VSUBS 0.014106f
C827 B.n787 VSUBS 0.014106f
C828 B.n788 VSUBS 0.014106f
C829 B.n789 VSUBS 0.014106f
C830 B.n790 VSUBS 0.014106f
C831 B.n791 VSUBS 0.014106f
C832 B.n792 VSUBS 0.014106f
C833 B.n793 VSUBS 0.014106f
C834 B.n794 VSUBS 0.014106f
C835 B.n795 VSUBS 0.014106f
C836 B.n796 VSUBS 0.014106f
C837 B.n797 VSUBS 0.014106f
C838 B.n798 VSUBS 0.014106f
C839 B.n799 VSUBS 0.014106f
C840 B.n800 VSUBS 0.014106f
C841 B.n801 VSUBS 0.014106f
C842 B.n802 VSUBS 0.014106f
C843 B.n803 VSUBS 0.014106f
C844 B.n804 VSUBS 0.014106f
C845 B.n805 VSUBS 0.014106f
C846 B.n806 VSUBS 0.014106f
C847 B.n807 VSUBS 0.018408f
C848 B.n808 VSUBS 0.019609f
C849 B.n809 VSUBS 0.038994f
C850 VDD2.t1 VSUBS 0.534489f
C851 VDD2.t4 VSUBS 0.075105f
C852 VDD2.t2 VSUBS 0.075105f
C853 VDD2.n0 VSUBS 0.347016f
C854 VDD2.n1 VSUBS 2.0706f
C855 VDD2.t5 VSUBS 0.075105f
C856 VDD2.t6 VSUBS 0.075105f
C857 VDD2.n2 VSUBS 0.3668f
C858 VDD2.n3 VSUBS 5.12007f
C859 VDD2.t9 VSUBS 0.515662f
C860 VDD2.n4 VSUBS 4.8405f
C861 VDD2.t8 VSUBS 0.075105f
C862 VDD2.t7 VSUBS 0.075105f
C863 VDD2.n5 VSUBS 0.347017f
C864 VDD2.n6 VSUBS 1.08995f
C865 VDD2.t0 VSUBS 0.075105f
C866 VDD2.t3 VSUBS 0.075105f
C867 VDD2.n7 VSUBS 0.366768f
C868 VN.t3 VSUBS 0.943298f
C869 VN.n0 VSUBS 0.583195f
C870 VN.n1 VSUBS 0.045614f
C871 VN.n2 VSUBS 0.090604f
C872 VN.n3 VSUBS 0.045614f
C873 VN.n4 VSUBS 0.084588f
C874 VN.n5 VSUBS 0.045614f
C875 VN.t4 VSUBS 0.943298f
C876 VN.n6 VSUBS 0.084588f
C877 VN.n7 VSUBS 0.045614f
C878 VN.n8 VSUBS 0.084588f
C879 VN.n9 VSUBS 0.045614f
C880 VN.t7 VSUBS 0.943298f
C881 VN.n10 VSUBS 0.084588f
C882 VN.n11 VSUBS 0.045614f
C883 VN.n12 VSUBS 0.084588f
C884 VN.t8 VSUBS 1.48456f
C885 VN.n13 VSUBS 0.652769f
C886 VN.t5 VSUBS 0.943298f
C887 VN.n14 VSUBS 0.588177f
C888 VN.n15 VSUBS 0.077071f
C889 VN.n16 VSUBS 0.58693f
C890 VN.n17 VSUBS 0.045614f
C891 VN.n18 VSUBS 0.045614f
C892 VN.n19 VSUBS 0.084588f
C893 VN.n20 VSUBS 0.056211f
C894 VN.n21 VSUBS 0.076404f
C895 VN.n22 VSUBS 0.045614f
C896 VN.n23 VSUBS 0.045614f
C897 VN.n24 VSUBS 0.045614f
C898 VN.n25 VSUBS 0.084588f
C899 VN.n26 VSUBS 0.063708f
C900 VN.n27 VSUBS 0.410591f
C901 VN.n28 VSUBS 0.063708f
C902 VN.n29 VSUBS 0.045614f
C903 VN.n30 VSUBS 0.045614f
C904 VN.n31 VSUBS 0.045614f
C905 VN.n32 VSUBS 0.084588f
C906 VN.n33 VSUBS 0.076404f
C907 VN.n34 VSUBS 0.056211f
C908 VN.n35 VSUBS 0.045614f
C909 VN.n36 VSUBS 0.045614f
C910 VN.n37 VSUBS 0.045614f
C911 VN.n38 VSUBS 0.084588f
C912 VN.n39 VSUBS 0.077071f
C913 VN.n40 VSUBS 0.410591f
C914 VN.n41 VSUBS 0.050346f
C915 VN.n42 VSUBS 0.045614f
C916 VN.n43 VSUBS 0.045614f
C917 VN.n44 VSUBS 0.045614f
C918 VN.n45 VSUBS 0.084588f
C919 VN.n46 VSUBS 0.0897f
C920 VN.n47 VSUBS 0.036899f
C921 VN.n48 VSUBS 0.045614f
C922 VN.n49 VSUBS 0.045614f
C923 VN.n50 VSUBS 0.045614f
C924 VN.n51 VSUBS 0.084588f
C925 VN.n52 VSUBS 0.084588f
C926 VN.n53 VSUBS 0.048675f
C927 VN.n54 VSUBS 0.073609f
C928 VN.n55 VSUBS 0.139948f
C929 VN.t0 VSUBS 0.943298f
C930 VN.n56 VSUBS 0.583195f
C931 VN.n57 VSUBS 0.045614f
C932 VN.n58 VSUBS 0.090604f
C933 VN.n59 VSUBS 0.045614f
C934 VN.n60 VSUBS 0.084588f
C935 VN.n61 VSUBS 0.045614f
C936 VN.t1 VSUBS 0.943298f
C937 VN.n62 VSUBS 0.084588f
C938 VN.n63 VSUBS 0.045614f
C939 VN.n64 VSUBS 0.084588f
C940 VN.n65 VSUBS 0.045614f
C941 VN.t2 VSUBS 0.943298f
C942 VN.n66 VSUBS 0.084588f
C943 VN.n67 VSUBS 0.045614f
C944 VN.n68 VSUBS 0.084588f
C945 VN.t6 VSUBS 1.48456f
C946 VN.n69 VSUBS 0.652769f
C947 VN.t9 VSUBS 0.943298f
C948 VN.n70 VSUBS 0.588177f
C949 VN.n71 VSUBS 0.077071f
C950 VN.n72 VSUBS 0.58693f
C951 VN.n73 VSUBS 0.045614f
C952 VN.n74 VSUBS 0.045614f
C953 VN.n75 VSUBS 0.084588f
C954 VN.n76 VSUBS 0.056211f
C955 VN.n77 VSUBS 0.076404f
C956 VN.n78 VSUBS 0.045614f
C957 VN.n79 VSUBS 0.045614f
C958 VN.n80 VSUBS 0.045614f
C959 VN.n81 VSUBS 0.084588f
C960 VN.n82 VSUBS 0.063708f
C961 VN.n83 VSUBS 0.410591f
C962 VN.n84 VSUBS 0.063708f
C963 VN.n85 VSUBS 0.045614f
C964 VN.n86 VSUBS 0.045614f
C965 VN.n87 VSUBS 0.045614f
C966 VN.n88 VSUBS 0.084588f
C967 VN.n89 VSUBS 0.076404f
C968 VN.n90 VSUBS 0.056211f
C969 VN.n91 VSUBS 0.045614f
C970 VN.n92 VSUBS 0.045614f
C971 VN.n93 VSUBS 0.045614f
C972 VN.n94 VSUBS 0.084588f
C973 VN.n95 VSUBS 0.077071f
C974 VN.n96 VSUBS 0.410591f
C975 VN.n97 VSUBS 0.050346f
C976 VN.n98 VSUBS 0.045614f
C977 VN.n99 VSUBS 0.045614f
C978 VN.n100 VSUBS 0.045614f
C979 VN.n101 VSUBS 0.084588f
C980 VN.n102 VSUBS 0.0897f
C981 VN.n103 VSUBS 0.036899f
C982 VN.n104 VSUBS 0.045614f
C983 VN.n105 VSUBS 0.045614f
C984 VN.n106 VSUBS 0.045614f
C985 VN.n107 VSUBS 0.084588f
C986 VN.n108 VSUBS 0.084588f
C987 VN.n109 VSUBS 0.048675f
C988 VN.n110 VSUBS 0.073609f
C989 VN.n111 VSUBS 2.82982f
C990 VDD1.t9 VSUBS 0.53875f
C991 VDD1.t7 VSUBS 0.075703f
C992 VDD1.t8 VSUBS 0.075703f
C993 VDD1.n0 VSUBS 0.349783f
C994 VDD1.n1 VSUBS 2.10143f
C995 VDD1.t0 VSUBS 0.538748f
C996 VDD1.t1 VSUBS 0.075703f
C997 VDD1.t2 VSUBS 0.075703f
C998 VDD1.n2 VSUBS 0.349782f
C999 VDD1.n3 VSUBS 2.0871f
C1000 VDD1.t4 VSUBS 0.075703f
C1001 VDD1.t3 VSUBS 0.075703f
C1002 VDD1.n4 VSUBS 0.369723f
C1003 VDD1.n5 VSUBS 5.41352f
C1004 VDD1.t5 VSUBS 0.075703f
C1005 VDD1.t6 VSUBS 0.075703f
C1006 VDD1.n6 VSUBS 0.349781f
C1007 VDD1.n7 VSUBS 5.10593f
C1008 VTAIL.t5 VSUBS 0.073817f
C1009 VTAIL.t6 VSUBS 0.073817f
C1010 VTAIL.n0 VSUBS 0.292787f
C1011 VTAIL.n1 VSUBS 1.12595f
C1012 VTAIL.t12 VSUBS 0.459127f
C1013 VTAIL.n2 VSUBS 1.27259f
C1014 VTAIL.t10 VSUBS 0.073817f
C1015 VTAIL.t13 VSUBS 0.073817f
C1016 VTAIL.n3 VSUBS 0.292787f
C1017 VTAIL.n4 VSUBS 1.41384f
C1018 VTAIL.t14 VSUBS 0.073817f
C1019 VTAIL.t9 VSUBS 0.073817f
C1020 VTAIL.n5 VSUBS 0.292787f
C1021 VTAIL.n6 VSUBS 2.71241f
C1022 VTAIL.t18 VSUBS 0.073817f
C1023 VTAIL.t1 VSUBS 0.073817f
C1024 VTAIL.n7 VSUBS 0.292788f
C1025 VTAIL.n8 VSUBS 2.71241f
C1026 VTAIL.t19 VSUBS 0.073817f
C1027 VTAIL.t0 VSUBS 0.073817f
C1028 VTAIL.n9 VSUBS 0.292788f
C1029 VTAIL.n10 VSUBS 1.41384f
C1030 VTAIL.t2 VSUBS 0.459129f
C1031 VTAIL.n11 VSUBS 1.27258f
C1032 VTAIL.t8 VSUBS 0.073817f
C1033 VTAIL.t11 VSUBS 0.073817f
C1034 VTAIL.n12 VSUBS 0.292788f
C1035 VTAIL.n13 VSUBS 1.2376f
C1036 VTAIL.t16 VSUBS 0.073817f
C1037 VTAIL.t15 VSUBS 0.073817f
C1038 VTAIL.n14 VSUBS 0.292788f
C1039 VTAIL.n15 VSUBS 1.41384f
C1040 VTAIL.t7 VSUBS 0.459127f
C1041 VTAIL.n16 VSUBS 2.26977f
C1042 VTAIL.t3 VSUBS 0.459127f
C1043 VTAIL.n17 VSUBS 2.26977f
C1044 VTAIL.t17 VSUBS 0.073817f
C1045 VTAIL.t4 VSUBS 0.073817f
C1046 VTAIL.n18 VSUBS 0.292787f
C1047 VTAIL.n19 VSUBS 1.04787f
C1048 VP.t6 VSUBS 1.08376f
C1049 VP.n0 VSUBS 0.670037f
C1050 VP.n1 VSUBS 0.052407f
C1051 VP.n2 VSUBS 0.104095f
C1052 VP.n3 VSUBS 0.052407f
C1053 VP.n4 VSUBS 0.097184f
C1054 VP.n5 VSUBS 0.052407f
C1055 VP.t5 VSUBS 1.08376f
C1056 VP.n6 VSUBS 0.097184f
C1057 VP.n7 VSUBS 0.052407f
C1058 VP.n8 VSUBS 0.097184f
C1059 VP.n9 VSUBS 0.052407f
C1060 VP.t7 VSUBS 1.08376f
C1061 VP.n10 VSUBS 0.097184f
C1062 VP.n11 VSUBS 0.052407f
C1063 VP.n12 VSUBS 0.097184f
C1064 VP.n13 VSUBS 0.052407f
C1065 VP.t8 VSUBS 1.08376f
C1066 VP.n14 VSUBS 0.097184f
C1067 VP.n15 VSUBS 0.052407f
C1068 VP.n16 VSUBS 0.097184f
C1069 VP.n17 VSUBS 0.08457f
C1070 VP.t9 VSUBS 1.08376f
C1071 VP.t3 VSUBS 1.08376f
C1072 VP.n18 VSUBS 0.670037f
C1073 VP.n19 VSUBS 0.052407f
C1074 VP.n20 VSUBS 0.104095f
C1075 VP.n21 VSUBS 0.052407f
C1076 VP.n22 VSUBS 0.097184f
C1077 VP.n23 VSUBS 0.052407f
C1078 VP.t4 VSUBS 1.08376f
C1079 VP.n24 VSUBS 0.097184f
C1080 VP.n25 VSUBS 0.052407f
C1081 VP.n26 VSUBS 0.097184f
C1082 VP.n27 VSUBS 0.052407f
C1083 VP.t1 VSUBS 1.08376f
C1084 VP.n28 VSUBS 0.097184f
C1085 VP.n29 VSUBS 0.052407f
C1086 VP.n30 VSUBS 0.097184f
C1087 VP.t0 VSUBS 1.70562f
C1088 VP.n31 VSUBS 0.749973f
C1089 VP.t2 VSUBS 1.08376f
C1090 VP.n32 VSUBS 0.675761f
C1091 VP.n33 VSUBS 0.088548f
C1092 VP.n34 VSUBS 0.674329f
C1093 VP.n35 VSUBS 0.052407f
C1094 VP.n36 VSUBS 0.052407f
C1095 VP.n37 VSUBS 0.097184f
C1096 VP.n38 VSUBS 0.064582f
C1097 VP.n39 VSUBS 0.087781f
C1098 VP.n40 VSUBS 0.052407f
C1099 VP.n41 VSUBS 0.052407f
C1100 VP.n42 VSUBS 0.052407f
C1101 VP.n43 VSUBS 0.097184f
C1102 VP.n44 VSUBS 0.073195f
C1103 VP.n45 VSUBS 0.471732f
C1104 VP.n46 VSUBS 0.073195f
C1105 VP.n47 VSUBS 0.052407f
C1106 VP.n48 VSUBS 0.052407f
C1107 VP.n49 VSUBS 0.052407f
C1108 VP.n50 VSUBS 0.097184f
C1109 VP.n51 VSUBS 0.087781f
C1110 VP.n52 VSUBS 0.064582f
C1111 VP.n53 VSUBS 0.052407f
C1112 VP.n54 VSUBS 0.052407f
C1113 VP.n55 VSUBS 0.052407f
C1114 VP.n56 VSUBS 0.097184f
C1115 VP.n57 VSUBS 0.088548f
C1116 VP.n58 VSUBS 0.471732f
C1117 VP.n59 VSUBS 0.057842f
C1118 VP.n60 VSUBS 0.052407f
C1119 VP.n61 VSUBS 0.052407f
C1120 VP.n62 VSUBS 0.052407f
C1121 VP.n63 VSUBS 0.097184f
C1122 VP.n64 VSUBS 0.103057f
C1123 VP.n65 VSUBS 0.042394f
C1124 VP.n66 VSUBS 0.052407f
C1125 VP.n67 VSUBS 0.052407f
C1126 VP.n68 VSUBS 0.052407f
C1127 VP.n69 VSUBS 0.097184f
C1128 VP.n70 VSUBS 0.097184f
C1129 VP.n71 VSUBS 0.055923f
C1130 VP.n72 VSUBS 0.08457f
C1131 VP.n73 VSUBS 3.23012f
C1132 VP.n74 VSUBS 3.26612f
C1133 VP.n75 VSUBS 0.670037f
C1134 VP.n76 VSUBS 0.055923f
C1135 VP.n77 VSUBS 0.097184f
C1136 VP.n78 VSUBS 0.052407f
C1137 VP.n79 VSUBS 0.052407f
C1138 VP.n80 VSUBS 0.052407f
C1139 VP.n81 VSUBS 0.104095f
C1140 VP.n82 VSUBS 0.042394f
C1141 VP.n83 VSUBS 0.103057f
C1142 VP.n84 VSUBS 0.052407f
C1143 VP.n85 VSUBS 0.052407f
C1144 VP.n86 VSUBS 0.052407f
C1145 VP.n87 VSUBS 0.097184f
C1146 VP.n88 VSUBS 0.057842f
C1147 VP.n89 VSUBS 0.471732f
C1148 VP.n90 VSUBS 0.088548f
C1149 VP.n91 VSUBS 0.052407f
C1150 VP.n92 VSUBS 0.052407f
C1151 VP.n93 VSUBS 0.052407f
C1152 VP.n94 VSUBS 0.097184f
C1153 VP.n95 VSUBS 0.064582f
C1154 VP.n96 VSUBS 0.087781f
C1155 VP.n97 VSUBS 0.052407f
C1156 VP.n98 VSUBS 0.052407f
C1157 VP.n99 VSUBS 0.052407f
C1158 VP.n100 VSUBS 0.097184f
C1159 VP.n101 VSUBS 0.073195f
C1160 VP.n102 VSUBS 0.471732f
C1161 VP.n103 VSUBS 0.073195f
C1162 VP.n104 VSUBS 0.052407f
C1163 VP.n105 VSUBS 0.052407f
C1164 VP.n106 VSUBS 0.052407f
C1165 VP.n107 VSUBS 0.097184f
C1166 VP.n108 VSUBS 0.087781f
C1167 VP.n109 VSUBS 0.064582f
C1168 VP.n110 VSUBS 0.052407f
C1169 VP.n111 VSUBS 0.052407f
C1170 VP.n112 VSUBS 0.052407f
C1171 VP.n113 VSUBS 0.097184f
C1172 VP.n114 VSUBS 0.088548f
C1173 VP.n115 VSUBS 0.471732f
C1174 VP.n116 VSUBS 0.057842f
C1175 VP.n117 VSUBS 0.052407f
C1176 VP.n118 VSUBS 0.052407f
C1177 VP.n119 VSUBS 0.052407f
C1178 VP.n120 VSUBS 0.097184f
C1179 VP.n121 VSUBS 0.103057f
C1180 VP.n122 VSUBS 0.042394f
C1181 VP.n123 VSUBS 0.052407f
C1182 VP.n124 VSUBS 0.052407f
C1183 VP.n125 VSUBS 0.052407f
C1184 VP.n126 VSUBS 0.097184f
C1185 VP.n127 VSUBS 0.097184f
C1186 VP.n128 VSUBS 0.055923f
C1187 VP.n129 VSUBS 0.08457f
C1188 VP.n130 VSUBS 0.160788f
.ends

