* NGSPICE file created from diff_pair_sample_0900.ext - technology: sky130A

.subckt diff_pair_sample_0900 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=0.92565 ps=5.94 w=5.61 l=0.35
X1 VDD2.t5 VN.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=2.1879 ps=12 w=5.61 l=0.35
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0 ps=0 w=5.61 l=0.35
X3 VDD1.t3 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0.92565 ps=5.94 w=5.61 l=0.35
X4 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0.92565 ps=5.94 w=5.61 l=0.35
X5 VDD2.t3 VN.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=2.1879 ps=12 w=5.61 l=0.35
X6 VTAIL.t9 VN.t3 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=0.92565 ps=5.94 w=5.61 l=0.35
X7 VDD1.t0 VP.t2 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=2.1879 ps=12 w=5.61 l=0.35
X8 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0 ps=0 w=5.61 l=0.35
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0 ps=0 w=5.61 l=0.35
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0 ps=0 w=5.61 l=0.35
X11 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0.92565 ps=5.94 w=5.61 l=0.35
X12 VDD1.t1 VP.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=2.1879 ps=12 w=5.61 l=0.35
X13 VTAIL.t8 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=0.92565 ps=5.94 w=5.61 l=0.35
X14 VTAIL.t3 VP.t4 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.92565 pd=5.94 as=0.92565 ps=5.94 w=5.61 l=0.35
X15 VDD1.t5 VP.t5 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1879 pd=12 as=0.92565 ps=5.94 w=5.61 l=0.35
R0 VP.n1 VP.t5 520.649
R1 VP.n8 VP.t2 499.945
R2 VP.n6 VP.t1 499.945
R3 VP.n3 VP.t3 499.945
R4 VP.n7 VP.t0 499.214
R5 VP.n2 VP.t4 499.214
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n7 VP.n0 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n4 VP.n1 70.5418
R11 VP.n7 VP.n6 47.4702
R12 VP.n8 VP.n7 47.4702
R13 VP.n3 VP.n2 47.4702
R14 VP.n5 VP.n4 35.0157
R15 VP.n2 VP.n1 20.6807
R16 VP.n5 VP.n0 0.189894
R17 VP.n9 VP.n0 0.189894
R18 VP VP.n9 0.0516364
R19 VDD1 VDD1.t5 71.3155
R20 VDD1.n1 VDD1.t3 71.2017
R21 VDD1.n1 VDD1.n0 67.3792
R22 VDD1.n3 VDD1.n2 67.288
R23 VDD1.n3 VDD1.n1 31.3328
R24 VDD1.n2 VDD1.t4 3.52991
R25 VDD1.n2 VDD1.t1 3.52991
R26 VDD1.n0 VDD1.t2 3.52991
R27 VDD1.n0 VDD1.t0 3.52991
R28 VDD1 VDD1.n3 0.0888621
R29 VTAIL.n7 VTAIL.t10 54.1388
R30 VTAIL.n11 VTAIL.t11 54.1386
R31 VTAIL.n2 VTAIL.t5 54.1386
R32 VTAIL.n10 VTAIL.t4 54.1386
R33 VTAIL.n9 VTAIL.n8 50.6094
R34 VTAIL.n6 VTAIL.n5 50.6094
R35 VTAIL.n1 VTAIL.n0 50.6092
R36 VTAIL.n4 VTAIL.n3 50.6092
R37 VTAIL.n6 VTAIL.n4 18.3755
R38 VTAIL.n11 VTAIL.n10 17.7893
R39 VTAIL.n0 VTAIL.t0 3.52991
R40 VTAIL.n0 VTAIL.t8 3.52991
R41 VTAIL.n3 VTAIL.t6 3.52991
R42 VTAIL.n3 VTAIL.t7 3.52991
R43 VTAIL.n8 VTAIL.t2 3.52991
R44 VTAIL.n8 VTAIL.t3 3.52991
R45 VTAIL.n5 VTAIL.t1 3.52991
R46 VTAIL.n5 VTAIL.t9 3.52991
R47 VTAIL.n9 VTAIL.n7 0.763431
R48 VTAIL.n2 VTAIL.n1 0.763431
R49 VTAIL.n7 VTAIL.n6 0.586707
R50 VTAIL.n10 VTAIL.n9 0.586707
R51 VTAIL.n4 VTAIL.n2 0.586707
R52 VTAIL VTAIL.n11 0.381966
R53 VTAIL VTAIL.n1 0.205241
R54 B.n292 B.t6 597.861
R55 B.n219 B.t17 597.861
R56 B.n65 B.t14 597.861
R57 B.n62 B.t10 597.861
R58 B.n416 B.n415 585
R59 B.n417 B.n416 585
R60 B.n172 B.n61 585
R61 B.n171 B.n170 585
R62 B.n169 B.n168 585
R63 B.n167 B.n166 585
R64 B.n165 B.n164 585
R65 B.n163 B.n162 585
R66 B.n161 B.n160 585
R67 B.n159 B.n158 585
R68 B.n157 B.n156 585
R69 B.n155 B.n154 585
R70 B.n153 B.n152 585
R71 B.n151 B.n150 585
R72 B.n149 B.n148 585
R73 B.n147 B.n146 585
R74 B.n145 B.n144 585
R75 B.n143 B.n142 585
R76 B.n141 B.n140 585
R77 B.n139 B.n138 585
R78 B.n137 B.n136 585
R79 B.n135 B.n134 585
R80 B.n133 B.n132 585
R81 B.n131 B.n130 585
R82 B.n129 B.n128 585
R83 B.n127 B.n126 585
R84 B.n125 B.n124 585
R85 B.n123 B.n122 585
R86 B.n121 B.n120 585
R87 B.n119 B.n118 585
R88 B.n117 B.n116 585
R89 B.n115 B.n114 585
R90 B.n113 B.n112 585
R91 B.n110 B.n109 585
R92 B.n108 B.n107 585
R93 B.n106 B.n105 585
R94 B.n104 B.n103 585
R95 B.n102 B.n101 585
R96 B.n100 B.n99 585
R97 B.n98 B.n97 585
R98 B.n96 B.n95 585
R99 B.n94 B.n93 585
R100 B.n92 B.n91 585
R101 B.n90 B.n89 585
R102 B.n88 B.n87 585
R103 B.n86 B.n85 585
R104 B.n84 B.n83 585
R105 B.n82 B.n81 585
R106 B.n80 B.n79 585
R107 B.n78 B.n77 585
R108 B.n76 B.n75 585
R109 B.n74 B.n73 585
R110 B.n72 B.n71 585
R111 B.n70 B.n69 585
R112 B.n68 B.n67 585
R113 B.n32 B.n31 585
R114 B.n414 B.n33 585
R115 B.n418 B.n33 585
R116 B.n413 B.n412 585
R117 B.n412 B.n29 585
R118 B.n411 B.n28 585
R119 B.n424 B.n28 585
R120 B.n410 B.n27 585
R121 B.n425 B.n27 585
R122 B.n409 B.n26 585
R123 B.n426 B.n26 585
R124 B.n408 B.n407 585
R125 B.n407 B.n22 585
R126 B.n406 B.n21 585
R127 B.n432 B.n21 585
R128 B.n405 B.n20 585
R129 B.n433 B.n20 585
R130 B.n404 B.n19 585
R131 B.n434 B.n19 585
R132 B.n403 B.n402 585
R133 B.n402 B.n18 585
R134 B.n401 B.n14 585
R135 B.n440 B.n14 585
R136 B.n400 B.n13 585
R137 B.n441 B.n13 585
R138 B.n399 B.n12 585
R139 B.n442 B.n12 585
R140 B.n398 B.n397 585
R141 B.n397 B.n11 585
R142 B.n396 B.n7 585
R143 B.n448 B.n7 585
R144 B.n395 B.n6 585
R145 B.n449 B.n6 585
R146 B.n394 B.n5 585
R147 B.n450 B.n5 585
R148 B.n393 B.n392 585
R149 B.n392 B.n4 585
R150 B.n391 B.n173 585
R151 B.n391 B.n390 585
R152 B.n380 B.n174 585
R153 B.n383 B.n174 585
R154 B.n382 B.n381 585
R155 B.n384 B.n382 585
R156 B.n379 B.n178 585
R157 B.n181 B.n178 585
R158 B.n378 B.n377 585
R159 B.n377 B.n376 585
R160 B.n180 B.n179 585
R161 B.n369 B.n180 585
R162 B.n368 B.n367 585
R163 B.n370 B.n368 585
R164 B.n366 B.n186 585
R165 B.n186 B.n185 585
R166 B.n365 B.n364 585
R167 B.n364 B.n363 585
R168 B.n188 B.n187 585
R169 B.n189 B.n188 585
R170 B.n356 B.n355 585
R171 B.n357 B.n356 585
R172 B.n354 B.n194 585
R173 B.n194 B.n193 585
R174 B.n353 B.n352 585
R175 B.n352 B.n351 585
R176 B.n196 B.n195 585
R177 B.n197 B.n196 585
R178 B.n344 B.n343 585
R179 B.n345 B.n344 585
R180 B.n200 B.n199 585
R181 B.n233 B.n232 585
R182 B.n234 B.n230 585
R183 B.n230 B.n201 585
R184 B.n236 B.n235 585
R185 B.n238 B.n229 585
R186 B.n241 B.n240 585
R187 B.n242 B.n228 585
R188 B.n244 B.n243 585
R189 B.n246 B.n227 585
R190 B.n249 B.n248 585
R191 B.n250 B.n226 585
R192 B.n252 B.n251 585
R193 B.n254 B.n225 585
R194 B.n257 B.n256 585
R195 B.n258 B.n224 585
R196 B.n260 B.n259 585
R197 B.n262 B.n223 585
R198 B.n265 B.n264 585
R199 B.n266 B.n222 585
R200 B.n268 B.n267 585
R201 B.n270 B.n221 585
R202 B.n273 B.n272 585
R203 B.n274 B.n218 585
R204 B.n277 B.n276 585
R205 B.n279 B.n217 585
R206 B.n282 B.n281 585
R207 B.n283 B.n216 585
R208 B.n285 B.n284 585
R209 B.n287 B.n215 585
R210 B.n290 B.n289 585
R211 B.n291 B.n214 585
R212 B.n296 B.n295 585
R213 B.n298 B.n213 585
R214 B.n301 B.n300 585
R215 B.n302 B.n212 585
R216 B.n304 B.n303 585
R217 B.n306 B.n211 585
R218 B.n309 B.n308 585
R219 B.n310 B.n210 585
R220 B.n312 B.n311 585
R221 B.n314 B.n209 585
R222 B.n317 B.n316 585
R223 B.n318 B.n208 585
R224 B.n320 B.n319 585
R225 B.n322 B.n207 585
R226 B.n325 B.n324 585
R227 B.n326 B.n206 585
R228 B.n328 B.n327 585
R229 B.n330 B.n205 585
R230 B.n333 B.n332 585
R231 B.n334 B.n204 585
R232 B.n336 B.n335 585
R233 B.n338 B.n203 585
R234 B.n341 B.n340 585
R235 B.n342 B.n202 585
R236 B.n347 B.n346 585
R237 B.n346 B.n345 585
R238 B.n348 B.n198 585
R239 B.n198 B.n197 585
R240 B.n350 B.n349 585
R241 B.n351 B.n350 585
R242 B.n192 B.n191 585
R243 B.n193 B.n192 585
R244 B.n359 B.n358 585
R245 B.n358 B.n357 585
R246 B.n360 B.n190 585
R247 B.n190 B.n189 585
R248 B.n362 B.n361 585
R249 B.n363 B.n362 585
R250 B.n184 B.n183 585
R251 B.n185 B.n184 585
R252 B.n372 B.n371 585
R253 B.n371 B.n370 585
R254 B.n373 B.n182 585
R255 B.n369 B.n182 585
R256 B.n375 B.n374 585
R257 B.n376 B.n375 585
R258 B.n177 B.n176 585
R259 B.n181 B.n177 585
R260 B.n386 B.n385 585
R261 B.n385 B.n384 585
R262 B.n387 B.n175 585
R263 B.n383 B.n175 585
R264 B.n389 B.n388 585
R265 B.n390 B.n389 585
R266 B.n2 B.n0 585
R267 B.n4 B.n2 585
R268 B.n3 B.n1 585
R269 B.n449 B.n3 585
R270 B.n447 B.n446 585
R271 B.n448 B.n447 585
R272 B.n445 B.n8 585
R273 B.n11 B.n8 585
R274 B.n444 B.n443 585
R275 B.n443 B.n442 585
R276 B.n10 B.n9 585
R277 B.n441 B.n10 585
R278 B.n439 B.n438 585
R279 B.n440 B.n439 585
R280 B.n437 B.n15 585
R281 B.n18 B.n15 585
R282 B.n436 B.n435 585
R283 B.n435 B.n434 585
R284 B.n17 B.n16 585
R285 B.n433 B.n17 585
R286 B.n431 B.n430 585
R287 B.n432 B.n431 585
R288 B.n429 B.n23 585
R289 B.n23 B.n22 585
R290 B.n428 B.n427 585
R291 B.n427 B.n426 585
R292 B.n25 B.n24 585
R293 B.n425 B.n25 585
R294 B.n423 B.n422 585
R295 B.n424 B.n423 585
R296 B.n421 B.n30 585
R297 B.n30 B.n29 585
R298 B.n420 B.n419 585
R299 B.n419 B.n418 585
R300 B.n452 B.n451 585
R301 B.n451 B.n450 585
R302 B.n346 B.n200 535.745
R303 B.n419 B.n32 535.745
R304 B.n344 B.n202 535.745
R305 B.n416 B.n33 535.745
R306 B.n417 B.n60 256.663
R307 B.n417 B.n59 256.663
R308 B.n417 B.n58 256.663
R309 B.n417 B.n57 256.663
R310 B.n417 B.n56 256.663
R311 B.n417 B.n55 256.663
R312 B.n417 B.n54 256.663
R313 B.n417 B.n53 256.663
R314 B.n417 B.n52 256.663
R315 B.n417 B.n51 256.663
R316 B.n417 B.n50 256.663
R317 B.n417 B.n49 256.663
R318 B.n417 B.n48 256.663
R319 B.n417 B.n47 256.663
R320 B.n417 B.n46 256.663
R321 B.n417 B.n45 256.663
R322 B.n417 B.n44 256.663
R323 B.n417 B.n43 256.663
R324 B.n417 B.n42 256.663
R325 B.n417 B.n41 256.663
R326 B.n417 B.n40 256.663
R327 B.n417 B.n39 256.663
R328 B.n417 B.n38 256.663
R329 B.n417 B.n37 256.663
R330 B.n417 B.n36 256.663
R331 B.n417 B.n35 256.663
R332 B.n417 B.n34 256.663
R333 B.n231 B.n201 256.663
R334 B.n237 B.n201 256.663
R335 B.n239 B.n201 256.663
R336 B.n245 B.n201 256.663
R337 B.n247 B.n201 256.663
R338 B.n253 B.n201 256.663
R339 B.n255 B.n201 256.663
R340 B.n261 B.n201 256.663
R341 B.n263 B.n201 256.663
R342 B.n269 B.n201 256.663
R343 B.n271 B.n201 256.663
R344 B.n278 B.n201 256.663
R345 B.n280 B.n201 256.663
R346 B.n286 B.n201 256.663
R347 B.n288 B.n201 256.663
R348 B.n297 B.n201 256.663
R349 B.n299 B.n201 256.663
R350 B.n305 B.n201 256.663
R351 B.n307 B.n201 256.663
R352 B.n313 B.n201 256.663
R353 B.n315 B.n201 256.663
R354 B.n321 B.n201 256.663
R355 B.n323 B.n201 256.663
R356 B.n329 B.n201 256.663
R357 B.n331 B.n201 256.663
R358 B.n337 B.n201 256.663
R359 B.n339 B.n201 256.663
R360 B.n346 B.n198 163.367
R361 B.n350 B.n198 163.367
R362 B.n350 B.n192 163.367
R363 B.n358 B.n192 163.367
R364 B.n358 B.n190 163.367
R365 B.n362 B.n190 163.367
R366 B.n362 B.n184 163.367
R367 B.n371 B.n184 163.367
R368 B.n371 B.n182 163.367
R369 B.n375 B.n182 163.367
R370 B.n375 B.n177 163.367
R371 B.n385 B.n177 163.367
R372 B.n385 B.n175 163.367
R373 B.n389 B.n175 163.367
R374 B.n389 B.n2 163.367
R375 B.n451 B.n2 163.367
R376 B.n451 B.n3 163.367
R377 B.n447 B.n3 163.367
R378 B.n447 B.n8 163.367
R379 B.n443 B.n8 163.367
R380 B.n443 B.n10 163.367
R381 B.n439 B.n10 163.367
R382 B.n439 B.n15 163.367
R383 B.n435 B.n15 163.367
R384 B.n435 B.n17 163.367
R385 B.n431 B.n17 163.367
R386 B.n431 B.n23 163.367
R387 B.n427 B.n23 163.367
R388 B.n427 B.n25 163.367
R389 B.n423 B.n25 163.367
R390 B.n423 B.n30 163.367
R391 B.n419 B.n30 163.367
R392 B.n232 B.n230 163.367
R393 B.n236 B.n230 163.367
R394 B.n240 B.n238 163.367
R395 B.n244 B.n228 163.367
R396 B.n248 B.n246 163.367
R397 B.n252 B.n226 163.367
R398 B.n256 B.n254 163.367
R399 B.n260 B.n224 163.367
R400 B.n264 B.n262 163.367
R401 B.n268 B.n222 163.367
R402 B.n272 B.n270 163.367
R403 B.n277 B.n218 163.367
R404 B.n281 B.n279 163.367
R405 B.n285 B.n216 163.367
R406 B.n289 B.n287 163.367
R407 B.n296 B.n214 163.367
R408 B.n300 B.n298 163.367
R409 B.n304 B.n212 163.367
R410 B.n308 B.n306 163.367
R411 B.n312 B.n210 163.367
R412 B.n316 B.n314 163.367
R413 B.n320 B.n208 163.367
R414 B.n324 B.n322 163.367
R415 B.n328 B.n206 163.367
R416 B.n332 B.n330 163.367
R417 B.n336 B.n204 163.367
R418 B.n340 B.n338 163.367
R419 B.n344 B.n196 163.367
R420 B.n352 B.n196 163.367
R421 B.n352 B.n194 163.367
R422 B.n356 B.n194 163.367
R423 B.n356 B.n188 163.367
R424 B.n364 B.n188 163.367
R425 B.n364 B.n186 163.367
R426 B.n368 B.n186 163.367
R427 B.n368 B.n180 163.367
R428 B.n377 B.n180 163.367
R429 B.n377 B.n178 163.367
R430 B.n382 B.n178 163.367
R431 B.n382 B.n174 163.367
R432 B.n391 B.n174 163.367
R433 B.n392 B.n391 163.367
R434 B.n392 B.n5 163.367
R435 B.n6 B.n5 163.367
R436 B.n7 B.n6 163.367
R437 B.n397 B.n7 163.367
R438 B.n397 B.n12 163.367
R439 B.n13 B.n12 163.367
R440 B.n14 B.n13 163.367
R441 B.n402 B.n14 163.367
R442 B.n402 B.n19 163.367
R443 B.n20 B.n19 163.367
R444 B.n21 B.n20 163.367
R445 B.n407 B.n21 163.367
R446 B.n407 B.n26 163.367
R447 B.n27 B.n26 163.367
R448 B.n28 B.n27 163.367
R449 B.n412 B.n28 163.367
R450 B.n412 B.n33 163.367
R451 B.n69 B.n68 163.367
R452 B.n73 B.n72 163.367
R453 B.n77 B.n76 163.367
R454 B.n81 B.n80 163.367
R455 B.n85 B.n84 163.367
R456 B.n89 B.n88 163.367
R457 B.n93 B.n92 163.367
R458 B.n97 B.n96 163.367
R459 B.n101 B.n100 163.367
R460 B.n105 B.n104 163.367
R461 B.n109 B.n108 163.367
R462 B.n114 B.n113 163.367
R463 B.n118 B.n117 163.367
R464 B.n122 B.n121 163.367
R465 B.n126 B.n125 163.367
R466 B.n130 B.n129 163.367
R467 B.n134 B.n133 163.367
R468 B.n138 B.n137 163.367
R469 B.n142 B.n141 163.367
R470 B.n146 B.n145 163.367
R471 B.n150 B.n149 163.367
R472 B.n154 B.n153 163.367
R473 B.n158 B.n157 163.367
R474 B.n162 B.n161 163.367
R475 B.n166 B.n165 163.367
R476 B.n170 B.n169 163.367
R477 B.n416 B.n61 163.367
R478 B.n345 B.n201 132.385
R479 B.n418 B.n417 132.385
R480 B.n292 B.t9 86.1786
R481 B.n62 B.t12 86.1786
R482 B.n219 B.t19 86.1728
R483 B.n65 B.t15 86.1728
R484 B.n293 B.t8 72.9907
R485 B.n63 B.t13 72.9907
R486 B.n220 B.t18 72.985
R487 B.n66 B.t16 72.985
R488 B.n231 B.n200 71.676
R489 B.n237 B.n236 71.676
R490 B.n240 B.n239 71.676
R491 B.n245 B.n244 71.676
R492 B.n248 B.n247 71.676
R493 B.n253 B.n252 71.676
R494 B.n256 B.n255 71.676
R495 B.n261 B.n260 71.676
R496 B.n264 B.n263 71.676
R497 B.n269 B.n268 71.676
R498 B.n272 B.n271 71.676
R499 B.n278 B.n277 71.676
R500 B.n281 B.n280 71.676
R501 B.n286 B.n285 71.676
R502 B.n289 B.n288 71.676
R503 B.n297 B.n296 71.676
R504 B.n300 B.n299 71.676
R505 B.n305 B.n304 71.676
R506 B.n308 B.n307 71.676
R507 B.n313 B.n312 71.676
R508 B.n316 B.n315 71.676
R509 B.n321 B.n320 71.676
R510 B.n324 B.n323 71.676
R511 B.n329 B.n328 71.676
R512 B.n332 B.n331 71.676
R513 B.n337 B.n336 71.676
R514 B.n340 B.n339 71.676
R515 B.n34 B.n32 71.676
R516 B.n69 B.n35 71.676
R517 B.n73 B.n36 71.676
R518 B.n77 B.n37 71.676
R519 B.n81 B.n38 71.676
R520 B.n85 B.n39 71.676
R521 B.n89 B.n40 71.676
R522 B.n93 B.n41 71.676
R523 B.n97 B.n42 71.676
R524 B.n101 B.n43 71.676
R525 B.n105 B.n44 71.676
R526 B.n109 B.n45 71.676
R527 B.n114 B.n46 71.676
R528 B.n118 B.n47 71.676
R529 B.n122 B.n48 71.676
R530 B.n126 B.n49 71.676
R531 B.n130 B.n50 71.676
R532 B.n134 B.n51 71.676
R533 B.n138 B.n52 71.676
R534 B.n142 B.n53 71.676
R535 B.n146 B.n54 71.676
R536 B.n150 B.n55 71.676
R537 B.n154 B.n56 71.676
R538 B.n158 B.n57 71.676
R539 B.n162 B.n58 71.676
R540 B.n166 B.n59 71.676
R541 B.n170 B.n60 71.676
R542 B.n61 B.n60 71.676
R543 B.n169 B.n59 71.676
R544 B.n165 B.n58 71.676
R545 B.n161 B.n57 71.676
R546 B.n157 B.n56 71.676
R547 B.n153 B.n55 71.676
R548 B.n149 B.n54 71.676
R549 B.n145 B.n53 71.676
R550 B.n141 B.n52 71.676
R551 B.n137 B.n51 71.676
R552 B.n133 B.n50 71.676
R553 B.n129 B.n49 71.676
R554 B.n125 B.n48 71.676
R555 B.n121 B.n47 71.676
R556 B.n117 B.n46 71.676
R557 B.n113 B.n45 71.676
R558 B.n108 B.n44 71.676
R559 B.n104 B.n43 71.676
R560 B.n100 B.n42 71.676
R561 B.n96 B.n41 71.676
R562 B.n92 B.n40 71.676
R563 B.n88 B.n39 71.676
R564 B.n84 B.n38 71.676
R565 B.n80 B.n37 71.676
R566 B.n76 B.n36 71.676
R567 B.n72 B.n35 71.676
R568 B.n68 B.n34 71.676
R569 B.n232 B.n231 71.676
R570 B.n238 B.n237 71.676
R571 B.n239 B.n228 71.676
R572 B.n246 B.n245 71.676
R573 B.n247 B.n226 71.676
R574 B.n254 B.n253 71.676
R575 B.n255 B.n224 71.676
R576 B.n262 B.n261 71.676
R577 B.n263 B.n222 71.676
R578 B.n270 B.n269 71.676
R579 B.n271 B.n218 71.676
R580 B.n279 B.n278 71.676
R581 B.n280 B.n216 71.676
R582 B.n287 B.n286 71.676
R583 B.n288 B.n214 71.676
R584 B.n298 B.n297 71.676
R585 B.n299 B.n212 71.676
R586 B.n306 B.n305 71.676
R587 B.n307 B.n210 71.676
R588 B.n314 B.n313 71.676
R589 B.n315 B.n208 71.676
R590 B.n322 B.n321 71.676
R591 B.n323 B.n206 71.676
R592 B.n330 B.n329 71.676
R593 B.n331 B.n204 71.676
R594 B.n338 B.n337 71.676
R595 B.n339 B.n202 71.676
R596 B.n345 B.n197 68.7189
R597 B.n351 B.n197 68.7189
R598 B.n351 B.n193 68.7189
R599 B.n357 B.n193 68.7189
R600 B.n363 B.n189 68.7189
R601 B.n363 B.n185 68.7189
R602 B.n370 B.n185 68.7189
R603 B.n370 B.n369 68.7189
R604 B.n376 B.n181 68.7189
R605 B.n384 B.n383 68.7189
R606 B.n390 B.n4 68.7189
R607 B.n450 B.n4 68.7189
R608 B.n450 B.n449 68.7189
R609 B.n449 B.n448 68.7189
R610 B.n442 B.n11 68.7189
R611 B.n441 B.n440 68.7189
R612 B.n434 B.n18 68.7189
R613 B.n434 B.n433 68.7189
R614 B.n433 B.n432 68.7189
R615 B.n432 B.n22 68.7189
R616 B.n426 B.n425 68.7189
R617 B.n425 B.n424 68.7189
R618 B.n424 B.n29 68.7189
R619 B.n418 B.n29 68.7189
R620 B.n294 B.n293 59.5399
R621 B.n275 B.n220 59.5399
R622 B.n111 B.n66 59.5399
R623 B.n64 B.n63 59.5399
R624 B.t7 B.n189 55.5816
R625 B.t11 B.n22 55.5816
R626 B.n376 B.t1 41.4337
R627 B.n384 B.t5 41.4337
R628 B.n390 B.t4 41.4337
R629 B.n448 B.t0 41.4337
R630 B.n442 B.t2 41.4337
R631 B.n440 B.t3 41.4337
R632 B.n420 B.n31 34.8103
R633 B.n415 B.n414 34.8103
R634 B.n343 B.n342 34.8103
R635 B.n347 B.n199 34.8103
R636 B.n369 B.t1 27.2858
R637 B.n181 B.t5 27.2858
R638 B.n383 B.t4 27.2858
R639 B.n11 B.t0 27.2858
R640 B.t2 B.n441 27.2858
R641 B.n18 B.t3 27.2858
R642 B B.n452 18.0485
R643 B.n293 B.n292 13.1884
R644 B.n220 B.n219 13.1884
R645 B.n66 B.n65 13.1884
R646 B.n63 B.n62 13.1884
R647 B.n357 B.t7 13.1378
R648 B.n426 B.t11 13.1378
R649 B.n67 B.n31 10.6151
R650 B.n70 B.n67 10.6151
R651 B.n71 B.n70 10.6151
R652 B.n74 B.n71 10.6151
R653 B.n75 B.n74 10.6151
R654 B.n78 B.n75 10.6151
R655 B.n79 B.n78 10.6151
R656 B.n82 B.n79 10.6151
R657 B.n83 B.n82 10.6151
R658 B.n86 B.n83 10.6151
R659 B.n87 B.n86 10.6151
R660 B.n90 B.n87 10.6151
R661 B.n91 B.n90 10.6151
R662 B.n94 B.n91 10.6151
R663 B.n95 B.n94 10.6151
R664 B.n98 B.n95 10.6151
R665 B.n99 B.n98 10.6151
R666 B.n102 B.n99 10.6151
R667 B.n103 B.n102 10.6151
R668 B.n106 B.n103 10.6151
R669 B.n107 B.n106 10.6151
R670 B.n110 B.n107 10.6151
R671 B.n115 B.n112 10.6151
R672 B.n116 B.n115 10.6151
R673 B.n119 B.n116 10.6151
R674 B.n120 B.n119 10.6151
R675 B.n123 B.n120 10.6151
R676 B.n124 B.n123 10.6151
R677 B.n127 B.n124 10.6151
R678 B.n128 B.n127 10.6151
R679 B.n132 B.n131 10.6151
R680 B.n135 B.n132 10.6151
R681 B.n136 B.n135 10.6151
R682 B.n139 B.n136 10.6151
R683 B.n140 B.n139 10.6151
R684 B.n143 B.n140 10.6151
R685 B.n144 B.n143 10.6151
R686 B.n147 B.n144 10.6151
R687 B.n148 B.n147 10.6151
R688 B.n151 B.n148 10.6151
R689 B.n152 B.n151 10.6151
R690 B.n155 B.n152 10.6151
R691 B.n156 B.n155 10.6151
R692 B.n159 B.n156 10.6151
R693 B.n160 B.n159 10.6151
R694 B.n163 B.n160 10.6151
R695 B.n164 B.n163 10.6151
R696 B.n167 B.n164 10.6151
R697 B.n168 B.n167 10.6151
R698 B.n171 B.n168 10.6151
R699 B.n172 B.n171 10.6151
R700 B.n415 B.n172 10.6151
R701 B.n343 B.n195 10.6151
R702 B.n353 B.n195 10.6151
R703 B.n354 B.n353 10.6151
R704 B.n355 B.n354 10.6151
R705 B.n355 B.n187 10.6151
R706 B.n365 B.n187 10.6151
R707 B.n366 B.n365 10.6151
R708 B.n367 B.n366 10.6151
R709 B.n367 B.n179 10.6151
R710 B.n378 B.n179 10.6151
R711 B.n379 B.n378 10.6151
R712 B.n381 B.n379 10.6151
R713 B.n381 B.n380 10.6151
R714 B.n380 B.n173 10.6151
R715 B.n393 B.n173 10.6151
R716 B.n394 B.n393 10.6151
R717 B.n395 B.n394 10.6151
R718 B.n396 B.n395 10.6151
R719 B.n398 B.n396 10.6151
R720 B.n399 B.n398 10.6151
R721 B.n400 B.n399 10.6151
R722 B.n401 B.n400 10.6151
R723 B.n403 B.n401 10.6151
R724 B.n404 B.n403 10.6151
R725 B.n405 B.n404 10.6151
R726 B.n406 B.n405 10.6151
R727 B.n408 B.n406 10.6151
R728 B.n409 B.n408 10.6151
R729 B.n410 B.n409 10.6151
R730 B.n411 B.n410 10.6151
R731 B.n413 B.n411 10.6151
R732 B.n414 B.n413 10.6151
R733 B.n233 B.n199 10.6151
R734 B.n234 B.n233 10.6151
R735 B.n235 B.n234 10.6151
R736 B.n235 B.n229 10.6151
R737 B.n241 B.n229 10.6151
R738 B.n242 B.n241 10.6151
R739 B.n243 B.n242 10.6151
R740 B.n243 B.n227 10.6151
R741 B.n249 B.n227 10.6151
R742 B.n250 B.n249 10.6151
R743 B.n251 B.n250 10.6151
R744 B.n251 B.n225 10.6151
R745 B.n257 B.n225 10.6151
R746 B.n258 B.n257 10.6151
R747 B.n259 B.n258 10.6151
R748 B.n259 B.n223 10.6151
R749 B.n265 B.n223 10.6151
R750 B.n266 B.n265 10.6151
R751 B.n267 B.n266 10.6151
R752 B.n267 B.n221 10.6151
R753 B.n273 B.n221 10.6151
R754 B.n274 B.n273 10.6151
R755 B.n276 B.n217 10.6151
R756 B.n282 B.n217 10.6151
R757 B.n283 B.n282 10.6151
R758 B.n284 B.n283 10.6151
R759 B.n284 B.n215 10.6151
R760 B.n290 B.n215 10.6151
R761 B.n291 B.n290 10.6151
R762 B.n295 B.n291 10.6151
R763 B.n301 B.n213 10.6151
R764 B.n302 B.n301 10.6151
R765 B.n303 B.n302 10.6151
R766 B.n303 B.n211 10.6151
R767 B.n309 B.n211 10.6151
R768 B.n310 B.n309 10.6151
R769 B.n311 B.n310 10.6151
R770 B.n311 B.n209 10.6151
R771 B.n317 B.n209 10.6151
R772 B.n318 B.n317 10.6151
R773 B.n319 B.n318 10.6151
R774 B.n319 B.n207 10.6151
R775 B.n325 B.n207 10.6151
R776 B.n326 B.n325 10.6151
R777 B.n327 B.n326 10.6151
R778 B.n327 B.n205 10.6151
R779 B.n333 B.n205 10.6151
R780 B.n334 B.n333 10.6151
R781 B.n335 B.n334 10.6151
R782 B.n335 B.n203 10.6151
R783 B.n341 B.n203 10.6151
R784 B.n342 B.n341 10.6151
R785 B.n348 B.n347 10.6151
R786 B.n349 B.n348 10.6151
R787 B.n349 B.n191 10.6151
R788 B.n359 B.n191 10.6151
R789 B.n360 B.n359 10.6151
R790 B.n361 B.n360 10.6151
R791 B.n361 B.n183 10.6151
R792 B.n372 B.n183 10.6151
R793 B.n373 B.n372 10.6151
R794 B.n374 B.n373 10.6151
R795 B.n374 B.n176 10.6151
R796 B.n386 B.n176 10.6151
R797 B.n387 B.n386 10.6151
R798 B.n388 B.n387 10.6151
R799 B.n388 B.n0 10.6151
R800 B.n446 B.n1 10.6151
R801 B.n446 B.n445 10.6151
R802 B.n445 B.n444 10.6151
R803 B.n444 B.n9 10.6151
R804 B.n438 B.n9 10.6151
R805 B.n438 B.n437 10.6151
R806 B.n437 B.n436 10.6151
R807 B.n436 B.n16 10.6151
R808 B.n430 B.n16 10.6151
R809 B.n430 B.n429 10.6151
R810 B.n429 B.n428 10.6151
R811 B.n428 B.n24 10.6151
R812 B.n422 B.n24 10.6151
R813 B.n422 B.n421 10.6151
R814 B.n421 B.n420 10.6151
R815 B.n112 B.n111 6.5566
R816 B.n128 B.n64 6.5566
R817 B.n276 B.n275 6.5566
R818 B.n295 B.n294 6.5566
R819 B.n111 B.n110 4.05904
R820 B.n131 B.n64 4.05904
R821 B.n275 B.n274 4.05904
R822 B.n294 B.n213 4.05904
R823 B.n452 B.n0 2.81026
R824 B.n452 B.n1 2.81026
R825 VN.n0 VN.t1 520.649
R826 VN.n4 VN.t2 520.649
R827 VN.n2 VN.t0 499.945
R828 VN.n6 VN.t4 499.945
R829 VN.n1 VN.t5 499.214
R830 VN.n5 VN.t3 499.214
R831 VN.n3 VN.n2 161.3
R832 VN.n7 VN.n6 161.3
R833 VN.n7 VN.n4 70.5418
R834 VN.n3 VN.n0 70.5418
R835 VN.n2 VN.n1 47.4702
R836 VN.n6 VN.n5 47.4702
R837 VN VN.n7 35.3963
R838 VN.n5 VN.n4 20.6807
R839 VN.n1 VN.n0 20.6807
R840 VN VN.n3 0.0516364
R841 VDD2.n1 VDD2.t4 71.2017
R842 VDD2.n2 VDD2.t1 70.8176
R843 VDD2.n1 VDD2.n0 67.3792
R844 VDD2 VDD2.n3 67.3764
R845 VDD2.n2 VDD2.n1 30.4567
R846 VDD2.n3 VDD2.t2 3.52991
R847 VDD2.n3 VDD2.t3 3.52991
R848 VDD2.n0 VDD2.t0 3.52991
R849 VDD2.n0 VDD2.t5 3.52991
R850 VDD2 VDD2.n2 0.498345
C0 VTAIL VP 1.43906f
C1 VDD1 VP 1.6701f
C2 VDD1 VTAIL 6.98929f
C3 VP VDD2 0.267063f
C4 VN VP 3.55917f
C5 VTAIL VDD2 7.02385f
C6 VDD1 VDD2 0.585596f
C7 VN VTAIL 1.42466f
C8 VDD1 VN 0.147699f
C9 VN VDD2 1.55317f
C10 VDD2 B 3.020224f
C11 VDD1 B 3.206603f
C12 VTAIL B 3.676684f
C13 VN B 5.241317f
C14 VP B 4.210046f
C15 VDD2.t4 B 1.0054f
C16 VDD2.t0 B 0.095637f
C17 VDD2.t5 B 0.095637f
C18 VDD2.n0 B 0.791142f
C19 VDD2.n1 B 1.32555f
C20 VDD2.t1 B 1.00401f
C21 VDD2.n2 B 1.43012f
C22 VDD2.t2 B 0.095637f
C23 VDD2.t3 B 0.095637f
C24 VDD2.n3 B 0.791124f
C25 VN.t1 B 0.177949f
C26 VN.n0 B 0.082678f
C27 VN.t5 B 0.174417f
C28 VN.n1 B 0.091925f
C29 VN.t0 B 0.174532f
C30 VN.n2 B 0.085879f
C31 VN.n3 B 0.088474f
C32 VN.t2 B 0.177949f
C33 VN.n4 B 0.082678f
C34 VN.t4 B 0.174532f
C35 VN.t3 B 0.174417f
C36 VN.n5 B 0.091925f
C37 VN.n6 B 0.085879f
C38 VN.n7 B 0.99578f
C39 VTAIL.t0 B 0.106327f
C40 VTAIL.t8 B 0.106327f
C41 VTAIL.n0 B 0.816937f
C42 VTAIL.n1 B 0.297991f
C43 VTAIL.t5 B 1.04169f
C44 VTAIL.n2 B 0.392703f
C45 VTAIL.t6 B 0.106327f
C46 VTAIL.t7 B 0.106327f
C47 VTAIL.n3 B 0.816937f
C48 VTAIL.n4 B 1.05867f
C49 VTAIL.t1 B 0.106327f
C50 VTAIL.t9 B 0.106327f
C51 VTAIL.n5 B 0.816942f
C52 VTAIL.n6 B 1.05867f
C53 VTAIL.t10 B 1.04169f
C54 VTAIL.n7 B 0.392699f
C55 VTAIL.t2 B 0.106327f
C56 VTAIL.t3 B 0.106327f
C57 VTAIL.n8 B 0.816942f
C58 VTAIL.n9 B 0.327467f
C59 VTAIL.t4 B 1.04169f
C60 VTAIL.n10 B 1.0786f
C61 VTAIL.t11 B 1.04169f
C62 VTAIL.n11 B 1.06277f
C63 VDD1.t5 B 0.994539f
C64 VDD1.t3 B 0.994086f
C65 VDD1.t2 B 0.094561f
C66 VDD1.t0 B 0.094561f
C67 VDD1.n0 B 0.782238f
C68 VDD1.n1 B 1.36802f
C69 VDD1.t4 B 0.094561f
C70 VDD1.t1 B 0.094561f
C71 VDD1.n2 B 0.781922f
C72 VDD1.n3 B 1.40046f
C73 VP.n0 B 0.030904f
C74 VP.t1 B 0.176638f
C75 VP.t5 B 0.180096f
C76 VP.n1 B 0.083675f
C77 VP.t4 B 0.176521f
C78 VP.n2 B 0.093035f
C79 VP.t3 B 0.176638f
C80 VP.n3 B 0.086916f
C81 VP.n4 B 0.987256f
C82 VP.n5 B 0.95339f
C83 VP.n6 B 0.086916f
C84 VP.t0 B 0.176521f
C85 VP.n7 B 0.093035f
C86 VP.t2 B 0.176638f
C87 VP.n8 B 0.086916f
C88 VP.n9 B 0.023949f
.ends

