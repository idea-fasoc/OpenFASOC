* NGSPICE file created from diff_pair_sample_0438.ext - technology: sky130A

.subckt diff_pair_sample_0438 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=4.4343 ps=23.52 w=11.37 l=2.03
X1 VTAIL.t3 VN.t0 VDD2.t5 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=1.87605 ps=11.7 w=11.37 l=2.03
X2 VDD1.t4 VP.t1 VTAIL.t7 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=1.87605 ps=11.7 w=11.37 l=2.03
X3 VTAIL.t9 VP.t2 VDD1.t3 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=1.87605 ps=11.7 w=11.37 l=2.03
X4 VTAIL.t5 VN.t1 VDD2.t4 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=1.87605 ps=11.7 w=11.37 l=2.03
X5 VDD1.t2 VP.t3 VTAIL.t6 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=1.87605 ps=11.7 w=11.37 l=2.03
X6 VDD2.t3 VN.t2 VTAIL.t1 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=4.4343 ps=23.52 w=11.37 l=2.03
X7 VDD2.t2 VN.t3 VTAIL.t2 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=4.4343 ps=23.52 w=11.37 l=2.03
X8 VDD2.t1 VN.t4 VTAIL.t4 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=1.87605 ps=11.7 w=11.37 l=2.03
X9 VDD1.t1 VP.t4 VTAIL.t8 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=4.4343 ps=23.52 w=11.37 l=2.03
X10 B.t11 B.t9 B.t10 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=2.03
X11 VDD2.t0 VN.t5 VTAIL.t0 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=1.87605 ps=11.7 w=11.37 l=2.03
X12 VTAIL.t10 VP.t5 VDD1.t0 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=1.87605 pd=11.7 as=1.87605 ps=11.7 w=11.37 l=2.03
X13 B.t8 B.t6 B.t7 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=2.03
X14 B.t5 B.t3 B.t4 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=2.03
X15 B.t2 B.t0 B.t1 w_n2858_n3242# sky130_fd_pr__pfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=2.03
R0 VP.n7 VP.t1 168.714
R1 VP.n10 VP.n9 161.3
R2 VP.n11 VP.n6 161.3
R3 VP.n13 VP.n12 161.3
R4 VP.n14 VP.n5 161.3
R5 VP.n31 VP.n0 161.3
R6 VP.n30 VP.n29 161.3
R7 VP.n28 VP.n1 161.3
R8 VP.n27 VP.n26 161.3
R9 VP.n25 VP.n2 161.3
R10 VP.n24 VP.n23 161.3
R11 VP.n22 VP.n3 161.3
R12 VP.n21 VP.n20 161.3
R13 VP.n19 VP.n4 161.3
R14 VP.n25 VP.t2 134.984
R15 VP.n18 VP.t3 134.984
R16 VP.n32 VP.t4 134.984
R17 VP.n8 VP.t5 134.984
R18 VP.n15 VP.t0 134.984
R19 VP.n18 VP.n17 93.1402
R20 VP.n33 VP.n32 93.1402
R21 VP.n16 VP.n15 93.1402
R22 VP.n30 VP.n1 56.5193
R23 VP.n20 VP.n3 56.5193
R24 VP.n13 VP.n6 56.5193
R25 VP.n17 VP.n16 45.9617
R26 VP.n8 VP.n7 45.8473
R27 VP.n20 VP.n19 24.4675
R28 VP.n24 VP.n3 24.4675
R29 VP.n25 VP.n24 24.4675
R30 VP.n26 VP.n25 24.4675
R31 VP.n26 VP.n1 24.4675
R32 VP.n31 VP.n30 24.4675
R33 VP.n14 VP.n13 24.4675
R34 VP.n9 VP.n8 24.4675
R35 VP.n9 VP.n6 24.4675
R36 VP.n19 VP.n18 17.6167
R37 VP.n32 VP.n31 17.6167
R38 VP.n15 VP.n14 17.6167
R39 VP.n10 VP.n7 9.19303
R40 VP.n16 VP.n5 0.278367
R41 VP.n17 VP.n4 0.278367
R42 VP.n33 VP.n0 0.278367
R43 VP.n11 VP.n10 0.189894
R44 VP.n12 VP.n11 0.189894
R45 VP.n12 VP.n5 0.189894
R46 VP.n21 VP.n4 0.189894
R47 VP.n22 VP.n21 0.189894
R48 VP.n23 VP.n22 0.189894
R49 VP.n23 VP.n2 0.189894
R50 VP.n27 VP.n2 0.189894
R51 VP.n28 VP.n27 0.189894
R52 VP.n29 VP.n28 0.189894
R53 VP.n29 VP.n0 0.189894
R54 VP VP.n33 0.153454
R55 VTAIL.n250 VTAIL.n194 756.745
R56 VTAIL.n58 VTAIL.n2 756.745
R57 VTAIL.n188 VTAIL.n132 756.745
R58 VTAIL.n124 VTAIL.n68 756.745
R59 VTAIL.n215 VTAIL.n214 585
R60 VTAIL.n217 VTAIL.n216 585
R61 VTAIL.n210 VTAIL.n209 585
R62 VTAIL.n223 VTAIL.n222 585
R63 VTAIL.n225 VTAIL.n224 585
R64 VTAIL.n206 VTAIL.n205 585
R65 VTAIL.n232 VTAIL.n231 585
R66 VTAIL.n233 VTAIL.n204 585
R67 VTAIL.n235 VTAIL.n234 585
R68 VTAIL.n202 VTAIL.n201 585
R69 VTAIL.n241 VTAIL.n240 585
R70 VTAIL.n243 VTAIL.n242 585
R71 VTAIL.n198 VTAIL.n197 585
R72 VTAIL.n249 VTAIL.n248 585
R73 VTAIL.n251 VTAIL.n250 585
R74 VTAIL.n23 VTAIL.n22 585
R75 VTAIL.n25 VTAIL.n24 585
R76 VTAIL.n18 VTAIL.n17 585
R77 VTAIL.n31 VTAIL.n30 585
R78 VTAIL.n33 VTAIL.n32 585
R79 VTAIL.n14 VTAIL.n13 585
R80 VTAIL.n40 VTAIL.n39 585
R81 VTAIL.n41 VTAIL.n12 585
R82 VTAIL.n43 VTAIL.n42 585
R83 VTAIL.n10 VTAIL.n9 585
R84 VTAIL.n49 VTAIL.n48 585
R85 VTAIL.n51 VTAIL.n50 585
R86 VTAIL.n6 VTAIL.n5 585
R87 VTAIL.n57 VTAIL.n56 585
R88 VTAIL.n59 VTAIL.n58 585
R89 VTAIL.n189 VTAIL.n188 585
R90 VTAIL.n187 VTAIL.n186 585
R91 VTAIL.n136 VTAIL.n135 585
R92 VTAIL.n181 VTAIL.n180 585
R93 VTAIL.n179 VTAIL.n178 585
R94 VTAIL.n140 VTAIL.n139 585
R95 VTAIL.n144 VTAIL.n142 585
R96 VTAIL.n173 VTAIL.n172 585
R97 VTAIL.n171 VTAIL.n170 585
R98 VTAIL.n146 VTAIL.n145 585
R99 VTAIL.n165 VTAIL.n164 585
R100 VTAIL.n163 VTAIL.n162 585
R101 VTAIL.n150 VTAIL.n149 585
R102 VTAIL.n157 VTAIL.n156 585
R103 VTAIL.n155 VTAIL.n154 585
R104 VTAIL.n125 VTAIL.n124 585
R105 VTAIL.n123 VTAIL.n122 585
R106 VTAIL.n72 VTAIL.n71 585
R107 VTAIL.n117 VTAIL.n116 585
R108 VTAIL.n115 VTAIL.n114 585
R109 VTAIL.n76 VTAIL.n75 585
R110 VTAIL.n80 VTAIL.n78 585
R111 VTAIL.n109 VTAIL.n108 585
R112 VTAIL.n107 VTAIL.n106 585
R113 VTAIL.n82 VTAIL.n81 585
R114 VTAIL.n101 VTAIL.n100 585
R115 VTAIL.n99 VTAIL.n98 585
R116 VTAIL.n86 VTAIL.n85 585
R117 VTAIL.n93 VTAIL.n92 585
R118 VTAIL.n91 VTAIL.n90 585
R119 VTAIL.n213 VTAIL.t2 329.036
R120 VTAIL.n21 VTAIL.t8 329.036
R121 VTAIL.n153 VTAIL.t11 329.036
R122 VTAIL.n89 VTAIL.t1 329.036
R123 VTAIL.n216 VTAIL.n215 171.744
R124 VTAIL.n216 VTAIL.n209 171.744
R125 VTAIL.n223 VTAIL.n209 171.744
R126 VTAIL.n224 VTAIL.n223 171.744
R127 VTAIL.n224 VTAIL.n205 171.744
R128 VTAIL.n232 VTAIL.n205 171.744
R129 VTAIL.n233 VTAIL.n232 171.744
R130 VTAIL.n234 VTAIL.n233 171.744
R131 VTAIL.n234 VTAIL.n201 171.744
R132 VTAIL.n241 VTAIL.n201 171.744
R133 VTAIL.n242 VTAIL.n241 171.744
R134 VTAIL.n242 VTAIL.n197 171.744
R135 VTAIL.n249 VTAIL.n197 171.744
R136 VTAIL.n250 VTAIL.n249 171.744
R137 VTAIL.n24 VTAIL.n23 171.744
R138 VTAIL.n24 VTAIL.n17 171.744
R139 VTAIL.n31 VTAIL.n17 171.744
R140 VTAIL.n32 VTAIL.n31 171.744
R141 VTAIL.n32 VTAIL.n13 171.744
R142 VTAIL.n40 VTAIL.n13 171.744
R143 VTAIL.n41 VTAIL.n40 171.744
R144 VTAIL.n42 VTAIL.n41 171.744
R145 VTAIL.n42 VTAIL.n9 171.744
R146 VTAIL.n49 VTAIL.n9 171.744
R147 VTAIL.n50 VTAIL.n49 171.744
R148 VTAIL.n50 VTAIL.n5 171.744
R149 VTAIL.n57 VTAIL.n5 171.744
R150 VTAIL.n58 VTAIL.n57 171.744
R151 VTAIL.n188 VTAIL.n187 171.744
R152 VTAIL.n187 VTAIL.n135 171.744
R153 VTAIL.n180 VTAIL.n135 171.744
R154 VTAIL.n180 VTAIL.n179 171.744
R155 VTAIL.n179 VTAIL.n139 171.744
R156 VTAIL.n144 VTAIL.n139 171.744
R157 VTAIL.n172 VTAIL.n144 171.744
R158 VTAIL.n172 VTAIL.n171 171.744
R159 VTAIL.n171 VTAIL.n145 171.744
R160 VTAIL.n164 VTAIL.n145 171.744
R161 VTAIL.n164 VTAIL.n163 171.744
R162 VTAIL.n163 VTAIL.n149 171.744
R163 VTAIL.n156 VTAIL.n149 171.744
R164 VTAIL.n156 VTAIL.n155 171.744
R165 VTAIL.n124 VTAIL.n123 171.744
R166 VTAIL.n123 VTAIL.n71 171.744
R167 VTAIL.n116 VTAIL.n71 171.744
R168 VTAIL.n116 VTAIL.n115 171.744
R169 VTAIL.n115 VTAIL.n75 171.744
R170 VTAIL.n80 VTAIL.n75 171.744
R171 VTAIL.n108 VTAIL.n80 171.744
R172 VTAIL.n108 VTAIL.n107 171.744
R173 VTAIL.n107 VTAIL.n81 171.744
R174 VTAIL.n100 VTAIL.n81 171.744
R175 VTAIL.n100 VTAIL.n99 171.744
R176 VTAIL.n99 VTAIL.n85 171.744
R177 VTAIL.n92 VTAIL.n85 171.744
R178 VTAIL.n92 VTAIL.n91 171.744
R179 VTAIL.n215 VTAIL.t2 85.8723
R180 VTAIL.n23 VTAIL.t8 85.8723
R181 VTAIL.n155 VTAIL.t11 85.8723
R182 VTAIL.n91 VTAIL.t1 85.8723
R183 VTAIL.n131 VTAIL.n130 57.5224
R184 VTAIL.n67 VTAIL.n66 57.5224
R185 VTAIL.n1 VTAIL.n0 57.5222
R186 VTAIL.n65 VTAIL.n64 57.5222
R187 VTAIL.n255 VTAIL.n254 31.6035
R188 VTAIL.n63 VTAIL.n62 31.6035
R189 VTAIL.n193 VTAIL.n192 31.6035
R190 VTAIL.n129 VTAIL.n128 31.6035
R191 VTAIL.n67 VTAIL.n65 26.2376
R192 VTAIL.n255 VTAIL.n193 24.2031
R193 VTAIL.n235 VTAIL.n202 13.1884
R194 VTAIL.n43 VTAIL.n10 13.1884
R195 VTAIL.n142 VTAIL.n140 13.1884
R196 VTAIL.n78 VTAIL.n76 13.1884
R197 VTAIL.n236 VTAIL.n204 12.8005
R198 VTAIL.n240 VTAIL.n239 12.8005
R199 VTAIL.n44 VTAIL.n12 12.8005
R200 VTAIL.n48 VTAIL.n47 12.8005
R201 VTAIL.n178 VTAIL.n177 12.8005
R202 VTAIL.n174 VTAIL.n173 12.8005
R203 VTAIL.n114 VTAIL.n113 12.8005
R204 VTAIL.n110 VTAIL.n109 12.8005
R205 VTAIL.n231 VTAIL.n230 12.0247
R206 VTAIL.n243 VTAIL.n200 12.0247
R207 VTAIL.n39 VTAIL.n38 12.0247
R208 VTAIL.n51 VTAIL.n8 12.0247
R209 VTAIL.n181 VTAIL.n138 12.0247
R210 VTAIL.n170 VTAIL.n143 12.0247
R211 VTAIL.n117 VTAIL.n74 12.0247
R212 VTAIL.n106 VTAIL.n79 12.0247
R213 VTAIL.n229 VTAIL.n206 11.249
R214 VTAIL.n244 VTAIL.n198 11.249
R215 VTAIL.n37 VTAIL.n14 11.249
R216 VTAIL.n52 VTAIL.n6 11.249
R217 VTAIL.n182 VTAIL.n136 11.249
R218 VTAIL.n169 VTAIL.n146 11.249
R219 VTAIL.n118 VTAIL.n72 11.249
R220 VTAIL.n105 VTAIL.n82 11.249
R221 VTAIL.n214 VTAIL.n213 10.7239
R222 VTAIL.n22 VTAIL.n21 10.7239
R223 VTAIL.n154 VTAIL.n153 10.7239
R224 VTAIL.n90 VTAIL.n89 10.7239
R225 VTAIL.n226 VTAIL.n225 10.4732
R226 VTAIL.n248 VTAIL.n247 10.4732
R227 VTAIL.n34 VTAIL.n33 10.4732
R228 VTAIL.n56 VTAIL.n55 10.4732
R229 VTAIL.n186 VTAIL.n185 10.4732
R230 VTAIL.n166 VTAIL.n165 10.4732
R231 VTAIL.n122 VTAIL.n121 10.4732
R232 VTAIL.n102 VTAIL.n101 10.4732
R233 VTAIL.n222 VTAIL.n208 9.69747
R234 VTAIL.n251 VTAIL.n196 9.69747
R235 VTAIL.n30 VTAIL.n16 9.69747
R236 VTAIL.n59 VTAIL.n4 9.69747
R237 VTAIL.n189 VTAIL.n134 9.69747
R238 VTAIL.n162 VTAIL.n148 9.69747
R239 VTAIL.n125 VTAIL.n70 9.69747
R240 VTAIL.n98 VTAIL.n84 9.69747
R241 VTAIL.n254 VTAIL.n253 9.45567
R242 VTAIL.n62 VTAIL.n61 9.45567
R243 VTAIL.n192 VTAIL.n191 9.45567
R244 VTAIL.n128 VTAIL.n127 9.45567
R245 VTAIL.n253 VTAIL.n252 9.3005
R246 VTAIL.n196 VTAIL.n195 9.3005
R247 VTAIL.n247 VTAIL.n246 9.3005
R248 VTAIL.n245 VTAIL.n244 9.3005
R249 VTAIL.n200 VTAIL.n199 9.3005
R250 VTAIL.n239 VTAIL.n238 9.3005
R251 VTAIL.n212 VTAIL.n211 9.3005
R252 VTAIL.n219 VTAIL.n218 9.3005
R253 VTAIL.n221 VTAIL.n220 9.3005
R254 VTAIL.n208 VTAIL.n207 9.3005
R255 VTAIL.n227 VTAIL.n226 9.3005
R256 VTAIL.n229 VTAIL.n228 9.3005
R257 VTAIL.n230 VTAIL.n203 9.3005
R258 VTAIL.n237 VTAIL.n236 9.3005
R259 VTAIL.n61 VTAIL.n60 9.3005
R260 VTAIL.n4 VTAIL.n3 9.3005
R261 VTAIL.n55 VTAIL.n54 9.3005
R262 VTAIL.n53 VTAIL.n52 9.3005
R263 VTAIL.n8 VTAIL.n7 9.3005
R264 VTAIL.n47 VTAIL.n46 9.3005
R265 VTAIL.n20 VTAIL.n19 9.3005
R266 VTAIL.n27 VTAIL.n26 9.3005
R267 VTAIL.n29 VTAIL.n28 9.3005
R268 VTAIL.n16 VTAIL.n15 9.3005
R269 VTAIL.n35 VTAIL.n34 9.3005
R270 VTAIL.n37 VTAIL.n36 9.3005
R271 VTAIL.n38 VTAIL.n11 9.3005
R272 VTAIL.n45 VTAIL.n44 9.3005
R273 VTAIL.n152 VTAIL.n151 9.3005
R274 VTAIL.n159 VTAIL.n158 9.3005
R275 VTAIL.n161 VTAIL.n160 9.3005
R276 VTAIL.n148 VTAIL.n147 9.3005
R277 VTAIL.n167 VTAIL.n166 9.3005
R278 VTAIL.n169 VTAIL.n168 9.3005
R279 VTAIL.n143 VTAIL.n141 9.3005
R280 VTAIL.n175 VTAIL.n174 9.3005
R281 VTAIL.n191 VTAIL.n190 9.3005
R282 VTAIL.n134 VTAIL.n133 9.3005
R283 VTAIL.n185 VTAIL.n184 9.3005
R284 VTAIL.n183 VTAIL.n182 9.3005
R285 VTAIL.n138 VTAIL.n137 9.3005
R286 VTAIL.n177 VTAIL.n176 9.3005
R287 VTAIL.n88 VTAIL.n87 9.3005
R288 VTAIL.n95 VTAIL.n94 9.3005
R289 VTAIL.n97 VTAIL.n96 9.3005
R290 VTAIL.n84 VTAIL.n83 9.3005
R291 VTAIL.n103 VTAIL.n102 9.3005
R292 VTAIL.n105 VTAIL.n104 9.3005
R293 VTAIL.n79 VTAIL.n77 9.3005
R294 VTAIL.n111 VTAIL.n110 9.3005
R295 VTAIL.n127 VTAIL.n126 9.3005
R296 VTAIL.n70 VTAIL.n69 9.3005
R297 VTAIL.n121 VTAIL.n120 9.3005
R298 VTAIL.n119 VTAIL.n118 9.3005
R299 VTAIL.n74 VTAIL.n73 9.3005
R300 VTAIL.n113 VTAIL.n112 9.3005
R301 VTAIL.n221 VTAIL.n210 8.92171
R302 VTAIL.n252 VTAIL.n194 8.92171
R303 VTAIL.n29 VTAIL.n18 8.92171
R304 VTAIL.n60 VTAIL.n2 8.92171
R305 VTAIL.n190 VTAIL.n132 8.92171
R306 VTAIL.n161 VTAIL.n150 8.92171
R307 VTAIL.n126 VTAIL.n68 8.92171
R308 VTAIL.n97 VTAIL.n86 8.92171
R309 VTAIL.n218 VTAIL.n217 8.14595
R310 VTAIL.n26 VTAIL.n25 8.14595
R311 VTAIL.n158 VTAIL.n157 8.14595
R312 VTAIL.n94 VTAIL.n93 8.14595
R313 VTAIL.n214 VTAIL.n212 7.3702
R314 VTAIL.n22 VTAIL.n20 7.3702
R315 VTAIL.n154 VTAIL.n152 7.3702
R316 VTAIL.n90 VTAIL.n88 7.3702
R317 VTAIL.n217 VTAIL.n212 5.81868
R318 VTAIL.n25 VTAIL.n20 5.81868
R319 VTAIL.n157 VTAIL.n152 5.81868
R320 VTAIL.n93 VTAIL.n88 5.81868
R321 VTAIL.n218 VTAIL.n210 5.04292
R322 VTAIL.n254 VTAIL.n194 5.04292
R323 VTAIL.n26 VTAIL.n18 5.04292
R324 VTAIL.n62 VTAIL.n2 5.04292
R325 VTAIL.n192 VTAIL.n132 5.04292
R326 VTAIL.n158 VTAIL.n150 5.04292
R327 VTAIL.n128 VTAIL.n68 5.04292
R328 VTAIL.n94 VTAIL.n86 5.04292
R329 VTAIL.n222 VTAIL.n221 4.26717
R330 VTAIL.n252 VTAIL.n251 4.26717
R331 VTAIL.n30 VTAIL.n29 4.26717
R332 VTAIL.n60 VTAIL.n59 4.26717
R333 VTAIL.n190 VTAIL.n189 4.26717
R334 VTAIL.n162 VTAIL.n161 4.26717
R335 VTAIL.n126 VTAIL.n125 4.26717
R336 VTAIL.n98 VTAIL.n97 4.26717
R337 VTAIL.n225 VTAIL.n208 3.49141
R338 VTAIL.n248 VTAIL.n196 3.49141
R339 VTAIL.n33 VTAIL.n16 3.49141
R340 VTAIL.n56 VTAIL.n4 3.49141
R341 VTAIL.n186 VTAIL.n134 3.49141
R342 VTAIL.n165 VTAIL.n148 3.49141
R343 VTAIL.n122 VTAIL.n70 3.49141
R344 VTAIL.n101 VTAIL.n84 3.49141
R345 VTAIL.n0 VTAIL.t0 2.85934
R346 VTAIL.n0 VTAIL.t5 2.85934
R347 VTAIL.n64 VTAIL.t6 2.85934
R348 VTAIL.n64 VTAIL.t9 2.85934
R349 VTAIL.n130 VTAIL.t7 2.85934
R350 VTAIL.n130 VTAIL.t10 2.85934
R351 VTAIL.n66 VTAIL.t4 2.85934
R352 VTAIL.n66 VTAIL.t3 2.85934
R353 VTAIL.n226 VTAIL.n206 2.71565
R354 VTAIL.n247 VTAIL.n198 2.71565
R355 VTAIL.n34 VTAIL.n14 2.71565
R356 VTAIL.n55 VTAIL.n6 2.71565
R357 VTAIL.n185 VTAIL.n136 2.71565
R358 VTAIL.n166 VTAIL.n146 2.71565
R359 VTAIL.n121 VTAIL.n72 2.71565
R360 VTAIL.n102 VTAIL.n82 2.71565
R361 VTAIL.n213 VTAIL.n211 2.41282
R362 VTAIL.n21 VTAIL.n19 2.41282
R363 VTAIL.n153 VTAIL.n151 2.41282
R364 VTAIL.n89 VTAIL.n87 2.41282
R365 VTAIL.n129 VTAIL.n67 2.03498
R366 VTAIL.n193 VTAIL.n131 2.03498
R367 VTAIL.n65 VTAIL.n63 2.03498
R368 VTAIL.n231 VTAIL.n229 1.93989
R369 VTAIL.n244 VTAIL.n243 1.93989
R370 VTAIL.n39 VTAIL.n37 1.93989
R371 VTAIL.n52 VTAIL.n51 1.93989
R372 VTAIL.n182 VTAIL.n181 1.93989
R373 VTAIL.n170 VTAIL.n169 1.93989
R374 VTAIL.n118 VTAIL.n117 1.93989
R375 VTAIL.n106 VTAIL.n105 1.93989
R376 VTAIL.n131 VTAIL.n129 1.48757
R377 VTAIL.n63 VTAIL.n1 1.48757
R378 VTAIL VTAIL.n255 1.46817
R379 VTAIL.n230 VTAIL.n204 1.16414
R380 VTAIL.n240 VTAIL.n200 1.16414
R381 VTAIL.n38 VTAIL.n12 1.16414
R382 VTAIL.n48 VTAIL.n8 1.16414
R383 VTAIL.n178 VTAIL.n138 1.16414
R384 VTAIL.n173 VTAIL.n143 1.16414
R385 VTAIL.n114 VTAIL.n74 1.16414
R386 VTAIL.n109 VTAIL.n79 1.16414
R387 VTAIL VTAIL.n1 0.56731
R388 VTAIL.n236 VTAIL.n235 0.388379
R389 VTAIL.n239 VTAIL.n202 0.388379
R390 VTAIL.n44 VTAIL.n43 0.388379
R391 VTAIL.n47 VTAIL.n10 0.388379
R392 VTAIL.n177 VTAIL.n140 0.388379
R393 VTAIL.n174 VTAIL.n142 0.388379
R394 VTAIL.n113 VTAIL.n76 0.388379
R395 VTAIL.n110 VTAIL.n78 0.388379
R396 VTAIL.n219 VTAIL.n211 0.155672
R397 VTAIL.n220 VTAIL.n219 0.155672
R398 VTAIL.n220 VTAIL.n207 0.155672
R399 VTAIL.n227 VTAIL.n207 0.155672
R400 VTAIL.n228 VTAIL.n227 0.155672
R401 VTAIL.n228 VTAIL.n203 0.155672
R402 VTAIL.n237 VTAIL.n203 0.155672
R403 VTAIL.n238 VTAIL.n237 0.155672
R404 VTAIL.n238 VTAIL.n199 0.155672
R405 VTAIL.n245 VTAIL.n199 0.155672
R406 VTAIL.n246 VTAIL.n245 0.155672
R407 VTAIL.n246 VTAIL.n195 0.155672
R408 VTAIL.n253 VTAIL.n195 0.155672
R409 VTAIL.n27 VTAIL.n19 0.155672
R410 VTAIL.n28 VTAIL.n27 0.155672
R411 VTAIL.n28 VTAIL.n15 0.155672
R412 VTAIL.n35 VTAIL.n15 0.155672
R413 VTAIL.n36 VTAIL.n35 0.155672
R414 VTAIL.n36 VTAIL.n11 0.155672
R415 VTAIL.n45 VTAIL.n11 0.155672
R416 VTAIL.n46 VTAIL.n45 0.155672
R417 VTAIL.n46 VTAIL.n7 0.155672
R418 VTAIL.n53 VTAIL.n7 0.155672
R419 VTAIL.n54 VTAIL.n53 0.155672
R420 VTAIL.n54 VTAIL.n3 0.155672
R421 VTAIL.n61 VTAIL.n3 0.155672
R422 VTAIL.n191 VTAIL.n133 0.155672
R423 VTAIL.n184 VTAIL.n133 0.155672
R424 VTAIL.n184 VTAIL.n183 0.155672
R425 VTAIL.n183 VTAIL.n137 0.155672
R426 VTAIL.n176 VTAIL.n137 0.155672
R427 VTAIL.n176 VTAIL.n175 0.155672
R428 VTAIL.n175 VTAIL.n141 0.155672
R429 VTAIL.n168 VTAIL.n141 0.155672
R430 VTAIL.n168 VTAIL.n167 0.155672
R431 VTAIL.n167 VTAIL.n147 0.155672
R432 VTAIL.n160 VTAIL.n147 0.155672
R433 VTAIL.n160 VTAIL.n159 0.155672
R434 VTAIL.n159 VTAIL.n151 0.155672
R435 VTAIL.n127 VTAIL.n69 0.155672
R436 VTAIL.n120 VTAIL.n69 0.155672
R437 VTAIL.n120 VTAIL.n119 0.155672
R438 VTAIL.n119 VTAIL.n73 0.155672
R439 VTAIL.n112 VTAIL.n73 0.155672
R440 VTAIL.n112 VTAIL.n111 0.155672
R441 VTAIL.n111 VTAIL.n77 0.155672
R442 VTAIL.n104 VTAIL.n77 0.155672
R443 VTAIL.n104 VTAIL.n103 0.155672
R444 VTAIL.n103 VTAIL.n83 0.155672
R445 VTAIL.n96 VTAIL.n83 0.155672
R446 VTAIL.n96 VTAIL.n95 0.155672
R447 VTAIL.n95 VTAIL.n87 0.155672
R448 VDD1.n56 VDD1.n0 756.745
R449 VDD1.n117 VDD1.n61 756.745
R450 VDD1.n57 VDD1.n56 585
R451 VDD1.n55 VDD1.n54 585
R452 VDD1.n4 VDD1.n3 585
R453 VDD1.n49 VDD1.n48 585
R454 VDD1.n47 VDD1.n46 585
R455 VDD1.n8 VDD1.n7 585
R456 VDD1.n12 VDD1.n10 585
R457 VDD1.n41 VDD1.n40 585
R458 VDD1.n39 VDD1.n38 585
R459 VDD1.n14 VDD1.n13 585
R460 VDD1.n33 VDD1.n32 585
R461 VDD1.n31 VDD1.n30 585
R462 VDD1.n18 VDD1.n17 585
R463 VDD1.n25 VDD1.n24 585
R464 VDD1.n23 VDD1.n22 585
R465 VDD1.n82 VDD1.n81 585
R466 VDD1.n84 VDD1.n83 585
R467 VDD1.n77 VDD1.n76 585
R468 VDD1.n90 VDD1.n89 585
R469 VDD1.n92 VDD1.n91 585
R470 VDD1.n73 VDD1.n72 585
R471 VDD1.n99 VDD1.n98 585
R472 VDD1.n100 VDD1.n71 585
R473 VDD1.n102 VDD1.n101 585
R474 VDD1.n69 VDD1.n68 585
R475 VDD1.n108 VDD1.n107 585
R476 VDD1.n110 VDD1.n109 585
R477 VDD1.n65 VDD1.n64 585
R478 VDD1.n116 VDD1.n115 585
R479 VDD1.n118 VDD1.n117 585
R480 VDD1.n21 VDD1.t4 329.036
R481 VDD1.n80 VDD1.t2 329.036
R482 VDD1.n56 VDD1.n55 171.744
R483 VDD1.n55 VDD1.n3 171.744
R484 VDD1.n48 VDD1.n3 171.744
R485 VDD1.n48 VDD1.n47 171.744
R486 VDD1.n47 VDD1.n7 171.744
R487 VDD1.n12 VDD1.n7 171.744
R488 VDD1.n40 VDD1.n12 171.744
R489 VDD1.n40 VDD1.n39 171.744
R490 VDD1.n39 VDD1.n13 171.744
R491 VDD1.n32 VDD1.n13 171.744
R492 VDD1.n32 VDD1.n31 171.744
R493 VDD1.n31 VDD1.n17 171.744
R494 VDD1.n24 VDD1.n17 171.744
R495 VDD1.n24 VDD1.n23 171.744
R496 VDD1.n83 VDD1.n82 171.744
R497 VDD1.n83 VDD1.n76 171.744
R498 VDD1.n90 VDD1.n76 171.744
R499 VDD1.n91 VDD1.n90 171.744
R500 VDD1.n91 VDD1.n72 171.744
R501 VDD1.n99 VDD1.n72 171.744
R502 VDD1.n100 VDD1.n99 171.744
R503 VDD1.n101 VDD1.n100 171.744
R504 VDD1.n101 VDD1.n68 171.744
R505 VDD1.n108 VDD1.n68 171.744
R506 VDD1.n109 VDD1.n108 171.744
R507 VDD1.n109 VDD1.n64 171.744
R508 VDD1.n116 VDD1.n64 171.744
R509 VDD1.n117 VDD1.n116 171.744
R510 VDD1.n23 VDD1.t4 85.8723
R511 VDD1.n82 VDD1.t2 85.8723
R512 VDD1.n123 VDD1.n122 74.6542
R513 VDD1.n125 VDD1.n124 74.201
R514 VDD1 VDD1.n60 49.8664
R515 VDD1.n123 VDD1.n121 49.7528
R516 VDD1.n125 VDD1.n123 41.7293
R517 VDD1.n10 VDD1.n8 13.1884
R518 VDD1.n102 VDD1.n69 13.1884
R519 VDD1.n46 VDD1.n45 12.8005
R520 VDD1.n42 VDD1.n41 12.8005
R521 VDD1.n103 VDD1.n71 12.8005
R522 VDD1.n107 VDD1.n106 12.8005
R523 VDD1.n49 VDD1.n6 12.0247
R524 VDD1.n38 VDD1.n11 12.0247
R525 VDD1.n98 VDD1.n97 12.0247
R526 VDD1.n110 VDD1.n67 12.0247
R527 VDD1.n50 VDD1.n4 11.249
R528 VDD1.n37 VDD1.n14 11.249
R529 VDD1.n96 VDD1.n73 11.249
R530 VDD1.n111 VDD1.n65 11.249
R531 VDD1.n22 VDD1.n21 10.7239
R532 VDD1.n81 VDD1.n80 10.7239
R533 VDD1.n54 VDD1.n53 10.4732
R534 VDD1.n34 VDD1.n33 10.4732
R535 VDD1.n93 VDD1.n92 10.4732
R536 VDD1.n115 VDD1.n114 10.4732
R537 VDD1.n57 VDD1.n2 9.69747
R538 VDD1.n30 VDD1.n16 9.69747
R539 VDD1.n89 VDD1.n75 9.69747
R540 VDD1.n118 VDD1.n63 9.69747
R541 VDD1.n60 VDD1.n59 9.45567
R542 VDD1.n121 VDD1.n120 9.45567
R543 VDD1.n20 VDD1.n19 9.3005
R544 VDD1.n27 VDD1.n26 9.3005
R545 VDD1.n29 VDD1.n28 9.3005
R546 VDD1.n16 VDD1.n15 9.3005
R547 VDD1.n35 VDD1.n34 9.3005
R548 VDD1.n37 VDD1.n36 9.3005
R549 VDD1.n11 VDD1.n9 9.3005
R550 VDD1.n43 VDD1.n42 9.3005
R551 VDD1.n59 VDD1.n58 9.3005
R552 VDD1.n2 VDD1.n1 9.3005
R553 VDD1.n53 VDD1.n52 9.3005
R554 VDD1.n51 VDD1.n50 9.3005
R555 VDD1.n6 VDD1.n5 9.3005
R556 VDD1.n45 VDD1.n44 9.3005
R557 VDD1.n120 VDD1.n119 9.3005
R558 VDD1.n63 VDD1.n62 9.3005
R559 VDD1.n114 VDD1.n113 9.3005
R560 VDD1.n112 VDD1.n111 9.3005
R561 VDD1.n67 VDD1.n66 9.3005
R562 VDD1.n106 VDD1.n105 9.3005
R563 VDD1.n79 VDD1.n78 9.3005
R564 VDD1.n86 VDD1.n85 9.3005
R565 VDD1.n88 VDD1.n87 9.3005
R566 VDD1.n75 VDD1.n74 9.3005
R567 VDD1.n94 VDD1.n93 9.3005
R568 VDD1.n96 VDD1.n95 9.3005
R569 VDD1.n97 VDD1.n70 9.3005
R570 VDD1.n104 VDD1.n103 9.3005
R571 VDD1.n58 VDD1.n0 8.92171
R572 VDD1.n29 VDD1.n18 8.92171
R573 VDD1.n88 VDD1.n77 8.92171
R574 VDD1.n119 VDD1.n61 8.92171
R575 VDD1.n26 VDD1.n25 8.14595
R576 VDD1.n85 VDD1.n84 8.14595
R577 VDD1.n22 VDD1.n20 7.3702
R578 VDD1.n81 VDD1.n79 7.3702
R579 VDD1.n25 VDD1.n20 5.81868
R580 VDD1.n84 VDD1.n79 5.81868
R581 VDD1.n60 VDD1.n0 5.04292
R582 VDD1.n26 VDD1.n18 5.04292
R583 VDD1.n85 VDD1.n77 5.04292
R584 VDD1.n121 VDD1.n61 5.04292
R585 VDD1.n58 VDD1.n57 4.26717
R586 VDD1.n30 VDD1.n29 4.26717
R587 VDD1.n89 VDD1.n88 4.26717
R588 VDD1.n119 VDD1.n118 4.26717
R589 VDD1.n54 VDD1.n2 3.49141
R590 VDD1.n33 VDD1.n16 3.49141
R591 VDD1.n92 VDD1.n75 3.49141
R592 VDD1.n115 VDD1.n63 3.49141
R593 VDD1.n124 VDD1.t0 2.85934
R594 VDD1.n124 VDD1.t5 2.85934
R595 VDD1.n122 VDD1.t3 2.85934
R596 VDD1.n122 VDD1.t1 2.85934
R597 VDD1.n53 VDD1.n4 2.71565
R598 VDD1.n34 VDD1.n14 2.71565
R599 VDD1.n93 VDD1.n73 2.71565
R600 VDD1.n114 VDD1.n65 2.71565
R601 VDD1.n21 VDD1.n19 2.41282
R602 VDD1.n80 VDD1.n78 2.41282
R603 VDD1.n50 VDD1.n49 1.93989
R604 VDD1.n38 VDD1.n37 1.93989
R605 VDD1.n98 VDD1.n96 1.93989
R606 VDD1.n111 VDD1.n110 1.93989
R607 VDD1.n46 VDD1.n6 1.16414
R608 VDD1.n41 VDD1.n11 1.16414
R609 VDD1.n97 VDD1.n71 1.16414
R610 VDD1.n107 VDD1.n67 1.16414
R611 VDD1 VDD1.n125 0.450931
R612 VDD1.n45 VDD1.n8 0.388379
R613 VDD1.n42 VDD1.n10 0.388379
R614 VDD1.n103 VDD1.n102 0.388379
R615 VDD1.n106 VDD1.n69 0.388379
R616 VDD1.n59 VDD1.n1 0.155672
R617 VDD1.n52 VDD1.n1 0.155672
R618 VDD1.n52 VDD1.n51 0.155672
R619 VDD1.n51 VDD1.n5 0.155672
R620 VDD1.n44 VDD1.n5 0.155672
R621 VDD1.n44 VDD1.n43 0.155672
R622 VDD1.n43 VDD1.n9 0.155672
R623 VDD1.n36 VDD1.n9 0.155672
R624 VDD1.n36 VDD1.n35 0.155672
R625 VDD1.n35 VDD1.n15 0.155672
R626 VDD1.n28 VDD1.n15 0.155672
R627 VDD1.n28 VDD1.n27 0.155672
R628 VDD1.n27 VDD1.n19 0.155672
R629 VDD1.n86 VDD1.n78 0.155672
R630 VDD1.n87 VDD1.n86 0.155672
R631 VDD1.n87 VDD1.n74 0.155672
R632 VDD1.n94 VDD1.n74 0.155672
R633 VDD1.n95 VDD1.n94 0.155672
R634 VDD1.n95 VDD1.n70 0.155672
R635 VDD1.n104 VDD1.n70 0.155672
R636 VDD1.n105 VDD1.n104 0.155672
R637 VDD1.n105 VDD1.n66 0.155672
R638 VDD1.n112 VDD1.n66 0.155672
R639 VDD1.n113 VDD1.n112 0.155672
R640 VDD1.n113 VDD1.n62 0.155672
R641 VDD1.n120 VDD1.n62 0.155672
R642 VN.n2 VN.t5 168.714
R643 VN.n14 VN.t2 168.714
R644 VN.n21 VN.n12 161.3
R645 VN.n20 VN.n19 161.3
R646 VN.n18 VN.n13 161.3
R647 VN.n17 VN.n16 161.3
R648 VN.n9 VN.n0 161.3
R649 VN.n8 VN.n7 161.3
R650 VN.n6 VN.n1 161.3
R651 VN.n5 VN.n4 161.3
R652 VN.n3 VN.t1 134.984
R653 VN.n10 VN.t3 134.984
R654 VN.n15 VN.t0 134.984
R655 VN.n22 VN.t4 134.984
R656 VN.n11 VN.n10 93.1402
R657 VN.n23 VN.n22 93.1402
R658 VN.n8 VN.n1 56.5193
R659 VN.n20 VN.n13 56.5193
R660 VN VN.n23 46.2406
R661 VN.n15 VN.n14 45.8473
R662 VN.n3 VN.n2 45.8473
R663 VN.n4 VN.n3 24.4675
R664 VN.n4 VN.n1 24.4675
R665 VN.n9 VN.n8 24.4675
R666 VN.n16 VN.n13 24.4675
R667 VN.n16 VN.n15 24.4675
R668 VN.n21 VN.n20 24.4675
R669 VN.n10 VN.n9 17.6167
R670 VN.n22 VN.n21 17.6167
R671 VN.n17 VN.n14 9.19303
R672 VN.n5 VN.n2 9.19303
R673 VN.n23 VN.n12 0.278367
R674 VN.n11 VN.n0 0.278367
R675 VN.n19 VN.n12 0.189894
R676 VN.n19 VN.n18 0.189894
R677 VN.n18 VN.n17 0.189894
R678 VN.n6 VN.n5 0.189894
R679 VN.n7 VN.n6 0.189894
R680 VN.n7 VN.n0 0.189894
R681 VN VN.n11 0.153454
R682 VDD2.n119 VDD2.n63 756.745
R683 VDD2.n56 VDD2.n0 756.745
R684 VDD2.n120 VDD2.n119 585
R685 VDD2.n118 VDD2.n117 585
R686 VDD2.n67 VDD2.n66 585
R687 VDD2.n112 VDD2.n111 585
R688 VDD2.n110 VDD2.n109 585
R689 VDD2.n71 VDD2.n70 585
R690 VDD2.n75 VDD2.n73 585
R691 VDD2.n104 VDD2.n103 585
R692 VDD2.n102 VDD2.n101 585
R693 VDD2.n77 VDD2.n76 585
R694 VDD2.n96 VDD2.n95 585
R695 VDD2.n94 VDD2.n93 585
R696 VDD2.n81 VDD2.n80 585
R697 VDD2.n88 VDD2.n87 585
R698 VDD2.n86 VDD2.n85 585
R699 VDD2.n21 VDD2.n20 585
R700 VDD2.n23 VDD2.n22 585
R701 VDD2.n16 VDD2.n15 585
R702 VDD2.n29 VDD2.n28 585
R703 VDD2.n31 VDD2.n30 585
R704 VDD2.n12 VDD2.n11 585
R705 VDD2.n38 VDD2.n37 585
R706 VDD2.n39 VDD2.n10 585
R707 VDD2.n41 VDD2.n40 585
R708 VDD2.n8 VDD2.n7 585
R709 VDD2.n47 VDD2.n46 585
R710 VDD2.n49 VDD2.n48 585
R711 VDD2.n4 VDD2.n3 585
R712 VDD2.n55 VDD2.n54 585
R713 VDD2.n57 VDD2.n56 585
R714 VDD2.n84 VDD2.t1 329.036
R715 VDD2.n19 VDD2.t0 329.036
R716 VDD2.n119 VDD2.n118 171.744
R717 VDD2.n118 VDD2.n66 171.744
R718 VDD2.n111 VDD2.n66 171.744
R719 VDD2.n111 VDD2.n110 171.744
R720 VDD2.n110 VDD2.n70 171.744
R721 VDD2.n75 VDD2.n70 171.744
R722 VDD2.n103 VDD2.n75 171.744
R723 VDD2.n103 VDD2.n102 171.744
R724 VDD2.n102 VDD2.n76 171.744
R725 VDD2.n95 VDD2.n76 171.744
R726 VDD2.n95 VDD2.n94 171.744
R727 VDD2.n94 VDD2.n80 171.744
R728 VDD2.n87 VDD2.n80 171.744
R729 VDD2.n87 VDD2.n86 171.744
R730 VDD2.n22 VDD2.n21 171.744
R731 VDD2.n22 VDD2.n15 171.744
R732 VDD2.n29 VDD2.n15 171.744
R733 VDD2.n30 VDD2.n29 171.744
R734 VDD2.n30 VDD2.n11 171.744
R735 VDD2.n38 VDD2.n11 171.744
R736 VDD2.n39 VDD2.n38 171.744
R737 VDD2.n40 VDD2.n39 171.744
R738 VDD2.n40 VDD2.n7 171.744
R739 VDD2.n47 VDD2.n7 171.744
R740 VDD2.n48 VDD2.n47 171.744
R741 VDD2.n48 VDD2.n3 171.744
R742 VDD2.n55 VDD2.n3 171.744
R743 VDD2.n56 VDD2.n55 171.744
R744 VDD2.n86 VDD2.t1 85.8723
R745 VDD2.n21 VDD2.t0 85.8723
R746 VDD2.n62 VDD2.n61 74.6542
R747 VDD2 VDD2.n125 74.6514
R748 VDD2.n62 VDD2.n60 49.7528
R749 VDD2.n124 VDD2.n123 48.2823
R750 VDD2.n124 VDD2.n62 40.1291
R751 VDD2.n73 VDD2.n71 13.1884
R752 VDD2.n41 VDD2.n8 13.1884
R753 VDD2.n109 VDD2.n108 12.8005
R754 VDD2.n105 VDD2.n104 12.8005
R755 VDD2.n42 VDD2.n10 12.8005
R756 VDD2.n46 VDD2.n45 12.8005
R757 VDD2.n112 VDD2.n69 12.0247
R758 VDD2.n101 VDD2.n74 12.0247
R759 VDD2.n37 VDD2.n36 12.0247
R760 VDD2.n49 VDD2.n6 12.0247
R761 VDD2.n113 VDD2.n67 11.249
R762 VDD2.n100 VDD2.n77 11.249
R763 VDD2.n35 VDD2.n12 11.249
R764 VDD2.n50 VDD2.n4 11.249
R765 VDD2.n85 VDD2.n84 10.7239
R766 VDD2.n20 VDD2.n19 10.7239
R767 VDD2.n117 VDD2.n116 10.4732
R768 VDD2.n97 VDD2.n96 10.4732
R769 VDD2.n32 VDD2.n31 10.4732
R770 VDD2.n54 VDD2.n53 10.4732
R771 VDD2.n120 VDD2.n65 9.69747
R772 VDD2.n93 VDD2.n79 9.69747
R773 VDD2.n28 VDD2.n14 9.69747
R774 VDD2.n57 VDD2.n2 9.69747
R775 VDD2.n123 VDD2.n122 9.45567
R776 VDD2.n60 VDD2.n59 9.45567
R777 VDD2.n83 VDD2.n82 9.3005
R778 VDD2.n90 VDD2.n89 9.3005
R779 VDD2.n92 VDD2.n91 9.3005
R780 VDD2.n79 VDD2.n78 9.3005
R781 VDD2.n98 VDD2.n97 9.3005
R782 VDD2.n100 VDD2.n99 9.3005
R783 VDD2.n74 VDD2.n72 9.3005
R784 VDD2.n106 VDD2.n105 9.3005
R785 VDD2.n122 VDD2.n121 9.3005
R786 VDD2.n65 VDD2.n64 9.3005
R787 VDD2.n116 VDD2.n115 9.3005
R788 VDD2.n114 VDD2.n113 9.3005
R789 VDD2.n69 VDD2.n68 9.3005
R790 VDD2.n108 VDD2.n107 9.3005
R791 VDD2.n59 VDD2.n58 9.3005
R792 VDD2.n2 VDD2.n1 9.3005
R793 VDD2.n53 VDD2.n52 9.3005
R794 VDD2.n51 VDD2.n50 9.3005
R795 VDD2.n6 VDD2.n5 9.3005
R796 VDD2.n45 VDD2.n44 9.3005
R797 VDD2.n18 VDD2.n17 9.3005
R798 VDD2.n25 VDD2.n24 9.3005
R799 VDD2.n27 VDD2.n26 9.3005
R800 VDD2.n14 VDD2.n13 9.3005
R801 VDD2.n33 VDD2.n32 9.3005
R802 VDD2.n35 VDD2.n34 9.3005
R803 VDD2.n36 VDD2.n9 9.3005
R804 VDD2.n43 VDD2.n42 9.3005
R805 VDD2.n121 VDD2.n63 8.92171
R806 VDD2.n92 VDD2.n81 8.92171
R807 VDD2.n27 VDD2.n16 8.92171
R808 VDD2.n58 VDD2.n0 8.92171
R809 VDD2.n89 VDD2.n88 8.14595
R810 VDD2.n24 VDD2.n23 8.14595
R811 VDD2.n85 VDD2.n83 7.3702
R812 VDD2.n20 VDD2.n18 7.3702
R813 VDD2.n88 VDD2.n83 5.81868
R814 VDD2.n23 VDD2.n18 5.81868
R815 VDD2.n123 VDD2.n63 5.04292
R816 VDD2.n89 VDD2.n81 5.04292
R817 VDD2.n24 VDD2.n16 5.04292
R818 VDD2.n60 VDD2.n0 5.04292
R819 VDD2.n121 VDD2.n120 4.26717
R820 VDD2.n93 VDD2.n92 4.26717
R821 VDD2.n28 VDD2.n27 4.26717
R822 VDD2.n58 VDD2.n57 4.26717
R823 VDD2.n117 VDD2.n65 3.49141
R824 VDD2.n96 VDD2.n79 3.49141
R825 VDD2.n31 VDD2.n14 3.49141
R826 VDD2.n54 VDD2.n2 3.49141
R827 VDD2.n125 VDD2.t5 2.85934
R828 VDD2.n125 VDD2.t3 2.85934
R829 VDD2.n61 VDD2.t4 2.85934
R830 VDD2.n61 VDD2.t2 2.85934
R831 VDD2.n116 VDD2.n67 2.71565
R832 VDD2.n97 VDD2.n77 2.71565
R833 VDD2.n32 VDD2.n12 2.71565
R834 VDD2.n53 VDD2.n4 2.71565
R835 VDD2.n84 VDD2.n82 2.41282
R836 VDD2.n19 VDD2.n17 2.41282
R837 VDD2.n113 VDD2.n112 1.93989
R838 VDD2.n101 VDD2.n100 1.93989
R839 VDD2.n37 VDD2.n35 1.93989
R840 VDD2.n50 VDD2.n49 1.93989
R841 VDD2 VDD2.n124 1.58455
R842 VDD2.n109 VDD2.n69 1.16414
R843 VDD2.n104 VDD2.n74 1.16414
R844 VDD2.n36 VDD2.n10 1.16414
R845 VDD2.n46 VDD2.n6 1.16414
R846 VDD2.n108 VDD2.n71 0.388379
R847 VDD2.n105 VDD2.n73 0.388379
R848 VDD2.n42 VDD2.n41 0.388379
R849 VDD2.n45 VDD2.n8 0.388379
R850 VDD2.n122 VDD2.n64 0.155672
R851 VDD2.n115 VDD2.n64 0.155672
R852 VDD2.n115 VDD2.n114 0.155672
R853 VDD2.n114 VDD2.n68 0.155672
R854 VDD2.n107 VDD2.n68 0.155672
R855 VDD2.n107 VDD2.n106 0.155672
R856 VDD2.n106 VDD2.n72 0.155672
R857 VDD2.n99 VDD2.n72 0.155672
R858 VDD2.n99 VDD2.n98 0.155672
R859 VDD2.n98 VDD2.n78 0.155672
R860 VDD2.n91 VDD2.n78 0.155672
R861 VDD2.n91 VDD2.n90 0.155672
R862 VDD2.n90 VDD2.n82 0.155672
R863 VDD2.n25 VDD2.n17 0.155672
R864 VDD2.n26 VDD2.n25 0.155672
R865 VDD2.n26 VDD2.n13 0.155672
R866 VDD2.n33 VDD2.n13 0.155672
R867 VDD2.n34 VDD2.n33 0.155672
R868 VDD2.n34 VDD2.n9 0.155672
R869 VDD2.n43 VDD2.n9 0.155672
R870 VDD2.n44 VDD2.n43 0.155672
R871 VDD2.n44 VDD2.n5 0.155672
R872 VDD2.n51 VDD2.n5 0.155672
R873 VDD2.n52 VDD2.n51 0.155672
R874 VDD2.n52 VDD2.n1 0.155672
R875 VDD2.n59 VDD2.n1 0.155672
R876 B.n470 B.n469 585
R877 B.n471 B.n68 585
R878 B.n473 B.n472 585
R879 B.n474 B.n67 585
R880 B.n476 B.n475 585
R881 B.n477 B.n66 585
R882 B.n479 B.n478 585
R883 B.n480 B.n65 585
R884 B.n482 B.n481 585
R885 B.n483 B.n64 585
R886 B.n485 B.n484 585
R887 B.n486 B.n63 585
R888 B.n488 B.n487 585
R889 B.n489 B.n62 585
R890 B.n491 B.n490 585
R891 B.n492 B.n61 585
R892 B.n494 B.n493 585
R893 B.n495 B.n60 585
R894 B.n497 B.n496 585
R895 B.n498 B.n59 585
R896 B.n500 B.n499 585
R897 B.n501 B.n58 585
R898 B.n503 B.n502 585
R899 B.n504 B.n57 585
R900 B.n506 B.n505 585
R901 B.n507 B.n56 585
R902 B.n509 B.n508 585
R903 B.n510 B.n55 585
R904 B.n512 B.n511 585
R905 B.n513 B.n54 585
R906 B.n515 B.n514 585
R907 B.n516 B.n53 585
R908 B.n518 B.n517 585
R909 B.n519 B.n52 585
R910 B.n521 B.n520 585
R911 B.n522 B.n51 585
R912 B.n524 B.n523 585
R913 B.n525 B.n50 585
R914 B.n527 B.n526 585
R915 B.n528 B.n47 585
R916 B.n531 B.n530 585
R917 B.n532 B.n46 585
R918 B.n534 B.n533 585
R919 B.n535 B.n45 585
R920 B.n537 B.n536 585
R921 B.n538 B.n44 585
R922 B.n540 B.n539 585
R923 B.n541 B.n43 585
R924 B.n543 B.n542 585
R925 B.n545 B.n544 585
R926 B.n546 B.n39 585
R927 B.n548 B.n547 585
R928 B.n549 B.n38 585
R929 B.n551 B.n550 585
R930 B.n552 B.n37 585
R931 B.n554 B.n553 585
R932 B.n555 B.n36 585
R933 B.n557 B.n556 585
R934 B.n558 B.n35 585
R935 B.n560 B.n559 585
R936 B.n561 B.n34 585
R937 B.n563 B.n562 585
R938 B.n564 B.n33 585
R939 B.n566 B.n565 585
R940 B.n567 B.n32 585
R941 B.n569 B.n568 585
R942 B.n570 B.n31 585
R943 B.n572 B.n571 585
R944 B.n573 B.n30 585
R945 B.n575 B.n574 585
R946 B.n576 B.n29 585
R947 B.n578 B.n577 585
R948 B.n579 B.n28 585
R949 B.n581 B.n580 585
R950 B.n582 B.n27 585
R951 B.n584 B.n583 585
R952 B.n585 B.n26 585
R953 B.n587 B.n586 585
R954 B.n588 B.n25 585
R955 B.n590 B.n589 585
R956 B.n591 B.n24 585
R957 B.n593 B.n592 585
R958 B.n594 B.n23 585
R959 B.n596 B.n595 585
R960 B.n597 B.n22 585
R961 B.n599 B.n598 585
R962 B.n600 B.n21 585
R963 B.n602 B.n601 585
R964 B.n603 B.n20 585
R965 B.n468 B.n69 585
R966 B.n467 B.n466 585
R967 B.n465 B.n70 585
R968 B.n464 B.n463 585
R969 B.n462 B.n71 585
R970 B.n461 B.n460 585
R971 B.n459 B.n72 585
R972 B.n458 B.n457 585
R973 B.n456 B.n73 585
R974 B.n455 B.n454 585
R975 B.n453 B.n74 585
R976 B.n452 B.n451 585
R977 B.n450 B.n75 585
R978 B.n449 B.n448 585
R979 B.n447 B.n76 585
R980 B.n446 B.n445 585
R981 B.n444 B.n77 585
R982 B.n443 B.n442 585
R983 B.n441 B.n78 585
R984 B.n440 B.n439 585
R985 B.n438 B.n79 585
R986 B.n437 B.n436 585
R987 B.n435 B.n80 585
R988 B.n434 B.n433 585
R989 B.n432 B.n81 585
R990 B.n431 B.n430 585
R991 B.n429 B.n82 585
R992 B.n428 B.n427 585
R993 B.n426 B.n83 585
R994 B.n425 B.n424 585
R995 B.n423 B.n84 585
R996 B.n422 B.n421 585
R997 B.n420 B.n85 585
R998 B.n419 B.n418 585
R999 B.n417 B.n86 585
R1000 B.n416 B.n415 585
R1001 B.n414 B.n87 585
R1002 B.n413 B.n412 585
R1003 B.n411 B.n88 585
R1004 B.n410 B.n409 585
R1005 B.n408 B.n89 585
R1006 B.n407 B.n406 585
R1007 B.n405 B.n90 585
R1008 B.n404 B.n403 585
R1009 B.n402 B.n91 585
R1010 B.n401 B.n400 585
R1011 B.n399 B.n92 585
R1012 B.n398 B.n397 585
R1013 B.n396 B.n93 585
R1014 B.n395 B.n394 585
R1015 B.n393 B.n94 585
R1016 B.n392 B.n391 585
R1017 B.n390 B.n95 585
R1018 B.n389 B.n388 585
R1019 B.n387 B.n96 585
R1020 B.n386 B.n385 585
R1021 B.n384 B.n97 585
R1022 B.n383 B.n382 585
R1023 B.n381 B.n98 585
R1024 B.n380 B.n379 585
R1025 B.n378 B.n99 585
R1026 B.n377 B.n376 585
R1027 B.n375 B.n100 585
R1028 B.n374 B.n373 585
R1029 B.n372 B.n101 585
R1030 B.n371 B.n370 585
R1031 B.n369 B.n102 585
R1032 B.n368 B.n367 585
R1033 B.n366 B.n103 585
R1034 B.n365 B.n364 585
R1035 B.n363 B.n104 585
R1036 B.n362 B.n361 585
R1037 B.n360 B.n105 585
R1038 B.n225 B.n154 585
R1039 B.n227 B.n226 585
R1040 B.n228 B.n153 585
R1041 B.n230 B.n229 585
R1042 B.n231 B.n152 585
R1043 B.n233 B.n232 585
R1044 B.n234 B.n151 585
R1045 B.n236 B.n235 585
R1046 B.n237 B.n150 585
R1047 B.n239 B.n238 585
R1048 B.n240 B.n149 585
R1049 B.n242 B.n241 585
R1050 B.n243 B.n148 585
R1051 B.n245 B.n244 585
R1052 B.n246 B.n147 585
R1053 B.n248 B.n247 585
R1054 B.n249 B.n146 585
R1055 B.n251 B.n250 585
R1056 B.n252 B.n145 585
R1057 B.n254 B.n253 585
R1058 B.n255 B.n144 585
R1059 B.n257 B.n256 585
R1060 B.n258 B.n143 585
R1061 B.n260 B.n259 585
R1062 B.n261 B.n142 585
R1063 B.n263 B.n262 585
R1064 B.n264 B.n141 585
R1065 B.n266 B.n265 585
R1066 B.n267 B.n140 585
R1067 B.n269 B.n268 585
R1068 B.n270 B.n139 585
R1069 B.n272 B.n271 585
R1070 B.n273 B.n138 585
R1071 B.n275 B.n274 585
R1072 B.n276 B.n137 585
R1073 B.n278 B.n277 585
R1074 B.n279 B.n136 585
R1075 B.n281 B.n280 585
R1076 B.n282 B.n135 585
R1077 B.n284 B.n283 585
R1078 B.n286 B.n285 585
R1079 B.n287 B.n131 585
R1080 B.n289 B.n288 585
R1081 B.n290 B.n130 585
R1082 B.n292 B.n291 585
R1083 B.n293 B.n129 585
R1084 B.n295 B.n294 585
R1085 B.n296 B.n128 585
R1086 B.n298 B.n297 585
R1087 B.n300 B.n125 585
R1088 B.n302 B.n301 585
R1089 B.n303 B.n124 585
R1090 B.n305 B.n304 585
R1091 B.n306 B.n123 585
R1092 B.n308 B.n307 585
R1093 B.n309 B.n122 585
R1094 B.n311 B.n310 585
R1095 B.n312 B.n121 585
R1096 B.n314 B.n313 585
R1097 B.n315 B.n120 585
R1098 B.n317 B.n316 585
R1099 B.n318 B.n119 585
R1100 B.n320 B.n319 585
R1101 B.n321 B.n118 585
R1102 B.n323 B.n322 585
R1103 B.n324 B.n117 585
R1104 B.n326 B.n325 585
R1105 B.n327 B.n116 585
R1106 B.n329 B.n328 585
R1107 B.n330 B.n115 585
R1108 B.n332 B.n331 585
R1109 B.n333 B.n114 585
R1110 B.n335 B.n334 585
R1111 B.n336 B.n113 585
R1112 B.n338 B.n337 585
R1113 B.n339 B.n112 585
R1114 B.n341 B.n340 585
R1115 B.n342 B.n111 585
R1116 B.n344 B.n343 585
R1117 B.n345 B.n110 585
R1118 B.n347 B.n346 585
R1119 B.n348 B.n109 585
R1120 B.n350 B.n349 585
R1121 B.n351 B.n108 585
R1122 B.n353 B.n352 585
R1123 B.n354 B.n107 585
R1124 B.n356 B.n355 585
R1125 B.n357 B.n106 585
R1126 B.n359 B.n358 585
R1127 B.n224 B.n223 585
R1128 B.n222 B.n155 585
R1129 B.n221 B.n220 585
R1130 B.n219 B.n156 585
R1131 B.n218 B.n217 585
R1132 B.n216 B.n157 585
R1133 B.n215 B.n214 585
R1134 B.n213 B.n158 585
R1135 B.n212 B.n211 585
R1136 B.n210 B.n159 585
R1137 B.n209 B.n208 585
R1138 B.n207 B.n160 585
R1139 B.n206 B.n205 585
R1140 B.n204 B.n161 585
R1141 B.n203 B.n202 585
R1142 B.n201 B.n162 585
R1143 B.n200 B.n199 585
R1144 B.n198 B.n163 585
R1145 B.n197 B.n196 585
R1146 B.n195 B.n164 585
R1147 B.n194 B.n193 585
R1148 B.n192 B.n165 585
R1149 B.n191 B.n190 585
R1150 B.n189 B.n166 585
R1151 B.n188 B.n187 585
R1152 B.n186 B.n167 585
R1153 B.n185 B.n184 585
R1154 B.n183 B.n168 585
R1155 B.n182 B.n181 585
R1156 B.n180 B.n169 585
R1157 B.n179 B.n178 585
R1158 B.n177 B.n170 585
R1159 B.n176 B.n175 585
R1160 B.n174 B.n171 585
R1161 B.n173 B.n172 585
R1162 B.n2 B.n0 585
R1163 B.n657 B.n1 585
R1164 B.n656 B.n655 585
R1165 B.n654 B.n3 585
R1166 B.n653 B.n652 585
R1167 B.n651 B.n4 585
R1168 B.n650 B.n649 585
R1169 B.n648 B.n5 585
R1170 B.n647 B.n646 585
R1171 B.n645 B.n6 585
R1172 B.n644 B.n643 585
R1173 B.n642 B.n7 585
R1174 B.n641 B.n640 585
R1175 B.n639 B.n8 585
R1176 B.n638 B.n637 585
R1177 B.n636 B.n9 585
R1178 B.n635 B.n634 585
R1179 B.n633 B.n10 585
R1180 B.n632 B.n631 585
R1181 B.n630 B.n11 585
R1182 B.n629 B.n628 585
R1183 B.n627 B.n12 585
R1184 B.n626 B.n625 585
R1185 B.n624 B.n13 585
R1186 B.n623 B.n622 585
R1187 B.n621 B.n14 585
R1188 B.n620 B.n619 585
R1189 B.n618 B.n15 585
R1190 B.n617 B.n616 585
R1191 B.n615 B.n16 585
R1192 B.n614 B.n613 585
R1193 B.n612 B.n17 585
R1194 B.n611 B.n610 585
R1195 B.n609 B.n18 585
R1196 B.n608 B.n607 585
R1197 B.n606 B.n19 585
R1198 B.n605 B.n604 585
R1199 B.n659 B.n658 585
R1200 B.n225 B.n224 487.695
R1201 B.n604 B.n603 487.695
R1202 B.n358 B.n105 487.695
R1203 B.n470 B.n69 487.695
R1204 B.n126 B.t2 410.024
R1205 B.n48 B.t7 410.024
R1206 B.n132 B.t11 410.024
R1207 B.n40 B.t4 410.024
R1208 B.n127 B.t1 364.255
R1209 B.n49 B.t8 364.255
R1210 B.n133 B.t10 364.255
R1211 B.n41 B.t5 364.255
R1212 B.n126 B.t0 341.971
R1213 B.n132 B.t9 341.971
R1214 B.n40 B.t3 341.971
R1215 B.n48 B.t6 341.971
R1216 B.n224 B.n155 163.367
R1217 B.n220 B.n155 163.367
R1218 B.n220 B.n219 163.367
R1219 B.n219 B.n218 163.367
R1220 B.n218 B.n157 163.367
R1221 B.n214 B.n157 163.367
R1222 B.n214 B.n213 163.367
R1223 B.n213 B.n212 163.367
R1224 B.n212 B.n159 163.367
R1225 B.n208 B.n159 163.367
R1226 B.n208 B.n207 163.367
R1227 B.n207 B.n206 163.367
R1228 B.n206 B.n161 163.367
R1229 B.n202 B.n161 163.367
R1230 B.n202 B.n201 163.367
R1231 B.n201 B.n200 163.367
R1232 B.n200 B.n163 163.367
R1233 B.n196 B.n163 163.367
R1234 B.n196 B.n195 163.367
R1235 B.n195 B.n194 163.367
R1236 B.n194 B.n165 163.367
R1237 B.n190 B.n165 163.367
R1238 B.n190 B.n189 163.367
R1239 B.n189 B.n188 163.367
R1240 B.n188 B.n167 163.367
R1241 B.n184 B.n167 163.367
R1242 B.n184 B.n183 163.367
R1243 B.n183 B.n182 163.367
R1244 B.n182 B.n169 163.367
R1245 B.n178 B.n169 163.367
R1246 B.n178 B.n177 163.367
R1247 B.n177 B.n176 163.367
R1248 B.n176 B.n171 163.367
R1249 B.n172 B.n171 163.367
R1250 B.n172 B.n2 163.367
R1251 B.n658 B.n2 163.367
R1252 B.n658 B.n657 163.367
R1253 B.n657 B.n656 163.367
R1254 B.n656 B.n3 163.367
R1255 B.n652 B.n3 163.367
R1256 B.n652 B.n651 163.367
R1257 B.n651 B.n650 163.367
R1258 B.n650 B.n5 163.367
R1259 B.n646 B.n5 163.367
R1260 B.n646 B.n645 163.367
R1261 B.n645 B.n644 163.367
R1262 B.n644 B.n7 163.367
R1263 B.n640 B.n7 163.367
R1264 B.n640 B.n639 163.367
R1265 B.n639 B.n638 163.367
R1266 B.n638 B.n9 163.367
R1267 B.n634 B.n9 163.367
R1268 B.n634 B.n633 163.367
R1269 B.n633 B.n632 163.367
R1270 B.n632 B.n11 163.367
R1271 B.n628 B.n11 163.367
R1272 B.n628 B.n627 163.367
R1273 B.n627 B.n626 163.367
R1274 B.n626 B.n13 163.367
R1275 B.n622 B.n13 163.367
R1276 B.n622 B.n621 163.367
R1277 B.n621 B.n620 163.367
R1278 B.n620 B.n15 163.367
R1279 B.n616 B.n15 163.367
R1280 B.n616 B.n615 163.367
R1281 B.n615 B.n614 163.367
R1282 B.n614 B.n17 163.367
R1283 B.n610 B.n17 163.367
R1284 B.n610 B.n609 163.367
R1285 B.n609 B.n608 163.367
R1286 B.n608 B.n19 163.367
R1287 B.n604 B.n19 163.367
R1288 B.n226 B.n225 163.367
R1289 B.n226 B.n153 163.367
R1290 B.n230 B.n153 163.367
R1291 B.n231 B.n230 163.367
R1292 B.n232 B.n231 163.367
R1293 B.n232 B.n151 163.367
R1294 B.n236 B.n151 163.367
R1295 B.n237 B.n236 163.367
R1296 B.n238 B.n237 163.367
R1297 B.n238 B.n149 163.367
R1298 B.n242 B.n149 163.367
R1299 B.n243 B.n242 163.367
R1300 B.n244 B.n243 163.367
R1301 B.n244 B.n147 163.367
R1302 B.n248 B.n147 163.367
R1303 B.n249 B.n248 163.367
R1304 B.n250 B.n249 163.367
R1305 B.n250 B.n145 163.367
R1306 B.n254 B.n145 163.367
R1307 B.n255 B.n254 163.367
R1308 B.n256 B.n255 163.367
R1309 B.n256 B.n143 163.367
R1310 B.n260 B.n143 163.367
R1311 B.n261 B.n260 163.367
R1312 B.n262 B.n261 163.367
R1313 B.n262 B.n141 163.367
R1314 B.n266 B.n141 163.367
R1315 B.n267 B.n266 163.367
R1316 B.n268 B.n267 163.367
R1317 B.n268 B.n139 163.367
R1318 B.n272 B.n139 163.367
R1319 B.n273 B.n272 163.367
R1320 B.n274 B.n273 163.367
R1321 B.n274 B.n137 163.367
R1322 B.n278 B.n137 163.367
R1323 B.n279 B.n278 163.367
R1324 B.n280 B.n279 163.367
R1325 B.n280 B.n135 163.367
R1326 B.n284 B.n135 163.367
R1327 B.n285 B.n284 163.367
R1328 B.n285 B.n131 163.367
R1329 B.n289 B.n131 163.367
R1330 B.n290 B.n289 163.367
R1331 B.n291 B.n290 163.367
R1332 B.n291 B.n129 163.367
R1333 B.n295 B.n129 163.367
R1334 B.n296 B.n295 163.367
R1335 B.n297 B.n296 163.367
R1336 B.n297 B.n125 163.367
R1337 B.n302 B.n125 163.367
R1338 B.n303 B.n302 163.367
R1339 B.n304 B.n303 163.367
R1340 B.n304 B.n123 163.367
R1341 B.n308 B.n123 163.367
R1342 B.n309 B.n308 163.367
R1343 B.n310 B.n309 163.367
R1344 B.n310 B.n121 163.367
R1345 B.n314 B.n121 163.367
R1346 B.n315 B.n314 163.367
R1347 B.n316 B.n315 163.367
R1348 B.n316 B.n119 163.367
R1349 B.n320 B.n119 163.367
R1350 B.n321 B.n320 163.367
R1351 B.n322 B.n321 163.367
R1352 B.n322 B.n117 163.367
R1353 B.n326 B.n117 163.367
R1354 B.n327 B.n326 163.367
R1355 B.n328 B.n327 163.367
R1356 B.n328 B.n115 163.367
R1357 B.n332 B.n115 163.367
R1358 B.n333 B.n332 163.367
R1359 B.n334 B.n333 163.367
R1360 B.n334 B.n113 163.367
R1361 B.n338 B.n113 163.367
R1362 B.n339 B.n338 163.367
R1363 B.n340 B.n339 163.367
R1364 B.n340 B.n111 163.367
R1365 B.n344 B.n111 163.367
R1366 B.n345 B.n344 163.367
R1367 B.n346 B.n345 163.367
R1368 B.n346 B.n109 163.367
R1369 B.n350 B.n109 163.367
R1370 B.n351 B.n350 163.367
R1371 B.n352 B.n351 163.367
R1372 B.n352 B.n107 163.367
R1373 B.n356 B.n107 163.367
R1374 B.n357 B.n356 163.367
R1375 B.n358 B.n357 163.367
R1376 B.n362 B.n105 163.367
R1377 B.n363 B.n362 163.367
R1378 B.n364 B.n363 163.367
R1379 B.n364 B.n103 163.367
R1380 B.n368 B.n103 163.367
R1381 B.n369 B.n368 163.367
R1382 B.n370 B.n369 163.367
R1383 B.n370 B.n101 163.367
R1384 B.n374 B.n101 163.367
R1385 B.n375 B.n374 163.367
R1386 B.n376 B.n375 163.367
R1387 B.n376 B.n99 163.367
R1388 B.n380 B.n99 163.367
R1389 B.n381 B.n380 163.367
R1390 B.n382 B.n381 163.367
R1391 B.n382 B.n97 163.367
R1392 B.n386 B.n97 163.367
R1393 B.n387 B.n386 163.367
R1394 B.n388 B.n387 163.367
R1395 B.n388 B.n95 163.367
R1396 B.n392 B.n95 163.367
R1397 B.n393 B.n392 163.367
R1398 B.n394 B.n393 163.367
R1399 B.n394 B.n93 163.367
R1400 B.n398 B.n93 163.367
R1401 B.n399 B.n398 163.367
R1402 B.n400 B.n399 163.367
R1403 B.n400 B.n91 163.367
R1404 B.n404 B.n91 163.367
R1405 B.n405 B.n404 163.367
R1406 B.n406 B.n405 163.367
R1407 B.n406 B.n89 163.367
R1408 B.n410 B.n89 163.367
R1409 B.n411 B.n410 163.367
R1410 B.n412 B.n411 163.367
R1411 B.n412 B.n87 163.367
R1412 B.n416 B.n87 163.367
R1413 B.n417 B.n416 163.367
R1414 B.n418 B.n417 163.367
R1415 B.n418 B.n85 163.367
R1416 B.n422 B.n85 163.367
R1417 B.n423 B.n422 163.367
R1418 B.n424 B.n423 163.367
R1419 B.n424 B.n83 163.367
R1420 B.n428 B.n83 163.367
R1421 B.n429 B.n428 163.367
R1422 B.n430 B.n429 163.367
R1423 B.n430 B.n81 163.367
R1424 B.n434 B.n81 163.367
R1425 B.n435 B.n434 163.367
R1426 B.n436 B.n435 163.367
R1427 B.n436 B.n79 163.367
R1428 B.n440 B.n79 163.367
R1429 B.n441 B.n440 163.367
R1430 B.n442 B.n441 163.367
R1431 B.n442 B.n77 163.367
R1432 B.n446 B.n77 163.367
R1433 B.n447 B.n446 163.367
R1434 B.n448 B.n447 163.367
R1435 B.n448 B.n75 163.367
R1436 B.n452 B.n75 163.367
R1437 B.n453 B.n452 163.367
R1438 B.n454 B.n453 163.367
R1439 B.n454 B.n73 163.367
R1440 B.n458 B.n73 163.367
R1441 B.n459 B.n458 163.367
R1442 B.n460 B.n459 163.367
R1443 B.n460 B.n71 163.367
R1444 B.n464 B.n71 163.367
R1445 B.n465 B.n464 163.367
R1446 B.n466 B.n465 163.367
R1447 B.n466 B.n69 163.367
R1448 B.n603 B.n602 163.367
R1449 B.n602 B.n21 163.367
R1450 B.n598 B.n21 163.367
R1451 B.n598 B.n597 163.367
R1452 B.n597 B.n596 163.367
R1453 B.n596 B.n23 163.367
R1454 B.n592 B.n23 163.367
R1455 B.n592 B.n591 163.367
R1456 B.n591 B.n590 163.367
R1457 B.n590 B.n25 163.367
R1458 B.n586 B.n25 163.367
R1459 B.n586 B.n585 163.367
R1460 B.n585 B.n584 163.367
R1461 B.n584 B.n27 163.367
R1462 B.n580 B.n27 163.367
R1463 B.n580 B.n579 163.367
R1464 B.n579 B.n578 163.367
R1465 B.n578 B.n29 163.367
R1466 B.n574 B.n29 163.367
R1467 B.n574 B.n573 163.367
R1468 B.n573 B.n572 163.367
R1469 B.n572 B.n31 163.367
R1470 B.n568 B.n31 163.367
R1471 B.n568 B.n567 163.367
R1472 B.n567 B.n566 163.367
R1473 B.n566 B.n33 163.367
R1474 B.n562 B.n33 163.367
R1475 B.n562 B.n561 163.367
R1476 B.n561 B.n560 163.367
R1477 B.n560 B.n35 163.367
R1478 B.n556 B.n35 163.367
R1479 B.n556 B.n555 163.367
R1480 B.n555 B.n554 163.367
R1481 B.n554 B.n37 163.367
R1482 B.n550 B.n37 163.367
R1483 B.n550 B.n549 163.367
R1484 B.n549 B.n548 163.367
R1485 B.n548 B.n39 163.367
R1486 B.n544 B.n39 163.367
R1487 B.n544 B.n543 163.367
R1488 B.n543 B.n43 163.367
R1489 B.n539 B.n43 163.367
R1490 B.n539 B.n538 163.367
R1491 B.n538 B.n537 163.367
R1492 B.n537 B.n45 163.367
R1493 B.n533 B.n45 163.367
R1494 B.n533 B.n532 163.367
R1495 B.n532 B.n531 163.367
R1496 B.n531 B.n47 163.367
R1497 B.n526 B.n47 163.367
R1498 B.n526 B.n525 163.367
R1499 B.n525 B.n524 163.367
R1500 B.n524 B.n51 163.367
R1501 B.n520 B.n51 163.367
R1502 B.n520 B.n519 163.367
R1503 B.n519 B.n518 163.367
R1504 B.n518 B.n53 163.367
R1505 B.n514 B.n53 163.367
R1506 B.n514 B.n513 163.367
R1507 B.n513 B.n512 163.367
R1508 B.n512 B.n55 163.367
R1509 B.n508 B.n55 163.367
R1510 B.n508 B.n507 163.367
R1511 B.n507 B.n506 163.367
R1512 B.n506 B.n57 163.367
R1513 B.n502 B.n57 163.367
R1514 B.n502 B.n501 163.367
R1515 B.n501 B.n500 163.367
R1516 B.n500 B.n59 163.367
R1517 B.n496 B.n59 163.367
R1518 B.n496 B.n495 163.367
R1519 B.n495 B.n494 163.367
R1520 B.n494 B.n61 163.367
R1521 B.n490 B.n61 163.367
R1522 B.n490 B.n489 163.367
R1523 B.n489 B.n488 163.367
R1524 B.n488 B.n63 163.367
R1525 B.n484 B.n63 163.367
R1526 B.n484 B.n483 163.367
R1527 B.n483 B.n482 163.367
R1528 B.n482 B.n65 163.367
R1529 B.n478 B.n65 163.367
R1530 B.n478 B.n477 163.367
R1531 B.n477 B.n476 163.367
R1532 B.n476 B.n67 163.367
R1533 B.n472 B.n67 163.367
R1534 B.n472 B.n471 163.367
R1535 B.n471 B.n470 163.367
R1536 B.n299 B.n127 59.5399
R1537 B.n134 B.n133 59.5399
R1538 B.n42 B.n41 59.5399
R1539 B.n529 B.n49 59.5399
R1540 B.n127 B.n126 45.7702
R1541 B.n133 B.n132 45.7702
R1542 B.n41 B.n40 45.7702
R1543 B.n49 B.n48 45.7702
R1544 B.n605 B.n20 31.6883
R1545 B.n469 B.n468 31.6883
R1546 B.n360 B.n359 31.6883
R1547 B.n223 B.n154 31.6883
R1548 B B.n659 18.0485
R1549 B.n601 B.n20 10.6151
R1550 B.n601 B.n600 10.6151
R1551 B.n600 B.n599 10.6151
R1552 B.n599 B.n22 10.6151
R1553 B.n595 B.n22 10.6151
R1554 B.n595 B.n594 10.6151
R1555 B.n594 B.n593 10.6151
R1556 B.n593 B.n24 10.6151
R1557 B.n589 B.n24 10.6151
R1558 B.n589 B.n588 10.6151
R1559 B.n588 B.n587 10.6151
R1560 B.n587 B.n26 10.6151
R1561 B.n583 B.n26 10.6151
R1562 B.n583 B.n582 10.6151
R1563 B.n582 B.n581 10.6151
R1564 B.n581 B.n28 10.6151
R1565 B.n577 B.n28 10.6151
R1566 B.n577 B.n576 10.6151
R1567 B.n576 B.n575 10.6151
R1568 B.n575 B.n30 10.6151
R1569 B.n571 B.n30 10.6151
R1570 B.n571 B.n570 10.6151
R1571 B.n570 B.n569 10.6151
R1572 B.n569 B.n32 10.6151
R1573 B.n565 B.n32 10.6151
R1574 B.n565 B.n564 10.6151
R1575 B.n564 B.n563 10.6151
R1576 B.n563 B.n34 10.6151
R1577 B.n559 B.n34 10.6151
R1578 B.n559 B.n558 10.6151
R1579 B.n558 B.n557 10.6151
R1580 B.n557 B.n36 10.6151
R1581 B.n553 B.n36 10.6151
R1582 B.n553 B.n552 10.6151
R1583 B.n552 B.n551 10.6151
R1584 B.n551 B.n38 10.6151
R1585 B.n547 B.n38 10.6151
R1586 B.n547 B.n546 10.6151
R1587 B.n546 B.n545 10.6151
R1588 B.n542 B.n541 10.6151
R1589 B.n541 B.n540 10.6151
R1590 B.n540 B.n44 10.6151
R1591 B.n536 B.n44 10.6151
R1592 B.n536 B.n535 10.6151
R1593 B.n535 B.n534 10.6151
R1594 B.n534 B.n46 10.6151
R1595 B.n530 B.n46 10.6151
R1596 B.n528 B.n527 10.6151
R1597 B.n527 B.n50 10.6151
R1598 B.n523 B.n50 10.6151
R1599 B.n523 B.n522 10.6151
R1600 B.n522 B.n521 10.6151
R1601 B.n521 B.n52 10.6151
R1602 B.n517 B.n52 10.6151
R1603 B.n517 B.n516 10.6151
R1604 B.n516 B.n515 10.6151
R1605 B.n515 B.n54 10.6151
R1606 B.n511 B.n54 10.6151
R1607 B.n511 B.n510 10.6151
R1608 B.n510 B.n509 10.6151
R1609 B.n509 B.n56 10.6151
R1610 B.n505 B.n56 10.6151
R1611 B.n505 B.n504 10.6151
R1612 B.n504 B.n503 10.6151
R1613 B.n503 B.n58 10.6151
R1614 B.n499 B.n58 10.6151
R1615 B.n499 B.n498 10.6151
R1616 B.n498 B.n497 10.6151
R1617 B.n497 B.n60 10.6151
R1618 B.n493 B.n60 10.6151
R1619 B.n493 B.n492 10.6151
R1620 B.n492 B.n491 10.6151
R1621 B.n491 B.n62 10.6151
R1622 B.n487 B.n62 10.6151
R1623 B.n487 B.n486 10.6151
R1624 B.n486 B.n485 10.6151
R1625 B.n485 B.n64 10.6151
R1626 B.n481 B.n64 10.6151
R1627 B.n481 B.n480 10.6151
R1628 B.n480 B.n479 10.6151
R1629 B.n479 B.n66 10.6151
R1630 B.n475 B.n66 10.6151
R1631 B.n475 B.n474 10.6151
R1632 B.n474 B.n473 10.6151
R1633 B.n473 B.n68 10.6151
R1634 B.n469 B.n68 10.6151
R1635 B.n361 B.n360 10.6151
R1636 B.n361 B.n104 10.6151
R1637 B.n365 B.n104 10.6151
R1638 B.n366 B.n365 10.6151
R1639 B.n367 B.n366 10.6151
R1640 B.n367 B.n102 10.6151
R1641 B.n371 B.n102 10.6151
R1642 B.n372 B.n371 10.6151
R1643 B.n373 B.n372 10.6151
R1644 B.n373 B.n100 10.6151
R1645 B.n377 B.n100 10.6151
R1646 B.n378 B.n377 10.6151
R1647 B.n379 B.n378 10.6151
R1648 B.n379 B.n98 10.6151
R1649 B.n383 B.n98 10.6151
R1650 B.n384 B.n383 10.6151
R1651 B.n385 B.n384 10.6151
R1652 B.n385 B.n96 10.6151
R1653 B.n389 B.n96 10.6151
R1654 B.n390 B.n389 10.6151
R1655 B.n391 B.n390 10.6151
R1656 B.n391 B.n94 10.6151
R1657 B.n395 B.n94 10.6151
R1658 B.n396 B.n395 10.6151
R1659 B.n397 B.n396 10.6151
R1660 B.n397 B.n92 10.6151
R1661 B.n401 B.n92 10.6151
R1662 B.n402 B.n401 10.6151
R1663 B.n403 B.n402 10.6151
R1664 B.n403 B.n90 10.6151
R1665 B.n407 B.n90 10.6151
R1666 B.n408 B.n407 10.6151
R1667 B.n409 B.n408 10.6151
R1668 B.n409 B.n88 10.6151
R1669 B.n413 B.n88 10.6151
R1670 B.n414 B.n413 10.6151
R1671 B.n415 B.n414 10.6151
R1672 B.n415 B.n86 10.6151
R1673 B.n419 B.n86 10.6151
R1674 B.n420 B.n419 10.6151
R1675 B.n421 B.n420 10.6151
R1676 B.n421 B.n84 10.6151
R1677 B.n425 B.n84 10.6151
R1678 B.n426 B.n425 10.6151
R1679 B.n427 B.n426 10.6151
R1680 B.n427 B.n82 10.6151
R1681 B.n431 B.n82 10.6151
R1682 B.n432 B.n431 10.6151
R1683 B.n433 B.n432 10.6151
R1684 B.n433 B.n80 10.6151
R1685 B.n437 B.n80 10.6151
R1686 B.n438 B.n437 10.6151
R1687 B.n439 B.n438 10.6151
R1688 B.n439 B.n78 10.6151
R1689 B.n443 B.n78 10.6151
R1690 B.n444 B.n443 10.6151
R1691 B.n445 B.n444 10.6151
R1692 B.n445 B.n76 10.6151
R1693 B.n449 B.n76 10.6151
R1694 B.n450 B.n449 10.6151
R1695 B.n451 B.n450 10.6151
R1696 B.n451 B.n74 10.6151
R1697 B.n455 B.n74 10.6151
R1698 B.n456 B.n455 10.6151
R1699 B.n457 B.n456 10.6151
R1700 B.n457 B.n72 10.6151
R1701 B.n461 B.n72 10.6151
R1702 B.n462 B.n461 10.6151
R1703 B.n463 B.n462 10.6151
R1704 B.n463 B.n70 10.6151
R1705 B.n467 B.n70 10.6151
R1706 B.n468 B.n467 10.6151
R1707 B.n227 B.n154 10.6151
R1708 B.n228 B.n227 10.6151
R1709 B.n229 B.n228 10.6151
R1710 B.n229 B.n152 10.6151
R1711 B.n233 B.n152 10.6151
R1712 B.n234 B.n233 10.6151
R1713 B.n235 B.n234 10.6151
R1714 B.n235 B.n150 10.6151
R1715 B.n239 B.n150 10.6151
R1716 B.n240 B.n239 10.6151
R1717 B.n241 B.n240 10.6151
R1718 B.n241 B.n148 10.6151
R1719 B.n245 B.n148 10.6151
R1720 B.n246 B.n245 10.6151
R1721 B.n247 B.n246 10.6151
R1722 B.n247 B.n146 10.6151
R1723 B.n251 B.n146 10.6151
R1724 B.n252 B.n251 10.6151
R1725 B.n253 B.n252 10.6151
R1726 B.n253 B.n144 10.6151
R1727 B.n257 B.n144 10.6151
R1728 B.n258 B.n257 10.6151
R1729 B.n259 B.n258 10.6151
R1730 B.n259 B.n142 10.6151
R1731 B.n263 B.n142 10.6151
R1732 B.n264 B.n263 10.6151
R1733 B.n265 B.n264 10.6151
R1734 B.n265 B.n140 10.6151
R1735 B.n269 B.n140 10.6151
R1736 B.n270 B.n269 10.6151
R1737 B.n271 B.n270 10.6151
R1738 B.n271 B.n138 10.6151
R1739 B.n275 B.n138 10.6151
R1740 B.n276 B.n275 10.6151
R1741 B.n277 B.n276 10.6151
R1742 B.n277 B.n136 10.6151
R1743 B.n281 B.n136 10.6151
R1744 B.n282 B.n281 10.6151
R1745 B.n283 B.n282 10.6151
R1746 B.n287 B.n286 10.6151
R1747 B.n288 B.n287 10.6151
R1748 B.n288 B.n130 10.6151
R1749 B.n292 B.n130 10.6151
R1750 B.n293 B.n292 10.6151
R1751 B.n294 B.n293 10.6151
R1752 B.n294 B.n128 10.6151
R1753 B.n298 B.n128 10.6151
R1754 B.n301 B.n300 10.6151
R1755 B.n301 B.n124 10.6151
R1756 B.n305 B.n124 10.6151
R1757 B.n306 B.n305 10.6151
R1758 B.n307 B.n306 10.6151
R1759 B.n307 B.n122 10.6151
R1760 B.n311 B.n122 10.6151
R1761 B.n312 B.n311 10.6151
R1762 B.n313 B.n312 10.6151
R1763 B.n313 B.n120 10.6151
R1764 B.n317 B.n120 10.6151
R1765 B.n318 B.n317 10.6151
R1766 B.n319 B.n318 10.6151
R1767 B.n319 B.n118 10.6151
R1768 B.n323 B.n118 10.6151
R1769 B.n324 B.n323 10.6151
R1770 B.n325 B.n324 10.6151
R1771 B.n325 B.n116 10.6151
R1772 B.n329 B.n116 10.6151
R1773 B.n330 B.n329 10.6151
R1774 B.n331 B.n330 10.6151
R1775 B.n331 B.n114 10.6151
R1776 B.n335 B.n114 10.6151
R1777 B.n336 B.n335 10.6151
R1778 B.n337 B.n336 10.6151
R1779 B.n337 B.n112 10.6151
R1780 B.n341 B.n112 10.6151
R1781 B.n342 B.n341 10.6151
R1782 B.n343 B.n342 10.6151
R1783 B.n343 B.n110 10.6151
R1784 B.n347 B.n110 10.6151
R1785 B.n348 B.n347 10.6151
R1786 B.n349 B.n348 10.6151
R1787 B.n349 B.n108 10.6151
R1788 B.n353 B.n108 10.6151
R1789 B.n354 B.n353 10.6151
R1790 B.n355 B.n354 10.6151
R1791 B.n355 B.n106 10.6151
R1792 B.n359 B.n106 10.6151
R1793 B.n223 B.n222 10.6151
R1794 B.n222 B.n221 10.6151
R1795 B.n221 B.n156 10.6151
R1796 B.n217 B.n156 10.6151
R1797 B.n217 B.n216 10.6151
R1798 B.n216 B.n215 10.6151
R1799 B.n215 B.n158 10.6151
R1800 B.n211 B.n158 10.6151
R1801 B.n211 B.n210 10.6151
R1802 B.n210 B.n209 10.6151
R1803 B.n209 B.n160 10.6151
R1804 B.n205 B.n160 10.6151
R1805 B.n205 B.n204 10.6151
R1806 B.n204 B.n203 10.6151
R1807 B.n203 B.n162 10.6151
R1808 B.n199 B.n162 10.6151
R1809 B.n199 B.n198 10.6151
R1810 B.n198 B.n197 10.6151
R1811 B.n197 B.n164 10.6151
R1812 B.n193 B.n164 10.6151
R1813 B.n193 B.n192 10.6151
R1814 B.n192 B.n191 10.6151
R1815 B.n191 B.n166 10.6151
R1816 B.n187 B.n166 10.6151
R1817 B.n187 B.n186 10.6151
R1818 B.n186 B.n185 10.6151
R1819 B.n185 B.n168 10.6151
R1820 B.n181 B.n168 10.6151
R1821 B.n181 B.n180 10.6151
R1822 B.n180 B.n179 10.6151
R1823 B.n179 B.n170 10.6151
R1824 B.n175 B.n170 10.6151
R1825 B.n175 B.n174 10.6151
R1826 B.n174 B.n173 10.6151
R1827 B.n173 B.n0 10.6151
R1828 B.n655 B.n1 10.6151
R1829 B.n655 B.n654 10.6151
R1830 B.n654 B.n653 10.6151
R1831 B.n653 B.n4 10.6151
R1832 B.n649 B.n4 10.6151
R1833 B.n649 B.n648 10.6151
R1834 B.n648 B.n647 10.6151
R1835 B.n647 B.n6 10.6151
R1836 B.n643 B.n6 10.6151
R1837 B.n643 B.n642 10.6151
R1838 B.n642 B.n641 10.6151
R1839 B.n641 B.n8 10.6151
R1840 B.n637 B.n8 10.6151
R1841 B.n637 B.n636 10.6151
R1842 B.n636 B.n635 10.6151
R1843 B.n635 B.n10 10.6151
R1844 B.n631 B.n10 10.6151
R1845 B.n631 B.n630 10.6151
R1846 B.n630 B.n629 10.6151
R1847 B.n629 B.n12 10.6151
R1848 B.n625 B.n12 10.6151
R1849 B.n625 B.n624 10.6151
R1850 B.n624 B.n623 10.6151
R1851 B.n623 B.n14 10.6151
R1852 B.n619 B.n14 10.6151
R1853 B.n619 B.n618 10.6151
R1854 B.n618 B.n617 10.6151
R1855 B.n617 B.n16 10.6151
R1856 B.n613 B.n16 10.6151
R1857 B.n613 B.n612 10.6151
R1858 B.n612 B.n611 10.6151
R1859 B.n611 B.n18 10.6151
R1860 B.n607 B.n18 10.6151
R1861 B.n607 B.n606 10.6151
R1862 B.n606 B.n605 10.6151
R1863 B.n542 B.n42 6.5566
R1864 B.n530 B.n529 6.5566
R1865 B.n286 B.n134 6.5566
R1866 B.n299 B.n298 6.5566
R1867 B.n545 B.n42 4.05904
R1868 B.n529 B.n528 4.05904
R1869 B.n283 B.n134 4.05904
R1870 B.n300 B.n299 4.05904
R1871 B.n659 B.n0 2.81026
R1872 B.n659 B.n1 2.81026
C0 VDD2 w_n2858_n3242# 2.17733f
C1 VTAIL VDD2 7.51902f
C2 VDD2 VN 6.06048f
C3 B w_n2858_n3242# 8.71166f
C4 VP w_n2858_n3242# 5.63674f
C5 VTAIL B 3.31217f
C6 B VN 1.03942f
C7 VTAIL VP 6.12824f
C8 VP VN 6.25883f
C9 VDD1 VDD2 1.1943f
C10 VTAIL w_n2858_n3242# 2.84722f
C11 VN w_n2858_n3242# 5.26883f
C12 VDD1 B 1.89236f
C13 VDD1 VP 6.31723f
C14 VTAIL VN 6.11391f
C15 B VDD2 1.95278f
C16 VP VDD2 0.410047f
C17 VDD1 w_n2858_n3242# 2.11043f
C18 VDD1 VTAIL 7.47255f
C19 VDD1 VN 0.150033f
C20 B VP 1.65082f
C21 VDD2 VSUBS 1.6437f
C22 VDD1 VSUBS 1.570322f
C23 VTAIL VSUBS 1.060162f
C24 VN VSUBS 5.28843f
C25 VP VSUBS 2.475417f
C26 B VSUBS 4.018236f
C27 w_n2858_n3242# VSUBS 0.114171p
C28 B.n0 VSUBS 0.004104f
C29 B.n1 VSUBS 0.004104f
C30 B.n2 VSUBS 0.00649f
C31 B.n3 VSUBS 0.00649f
C32 B.n4 VSUBS 0.00649f
C33 B.n5 VSUBS 0.00649f
C34 B.n6 VSUBS 0.00649f
C35 B.n7 VSUBS 0.00649f
C36 B.n8 VSUBS 0.00649f
C37 B.n9 VSUBS 0.00649f
C38 B.n10 VSUBS 0.00649f
C39 B.n11 VSUBS 0.00649f
C40 B.n12 VSUBS 0.00649f
C41 B.n13 VSUBS 0.00649f
C42 B.n14 VSUBS 0.00649f
C43 B.n15 VSUBS 0.00649f
C44 B.n16 VSUBS 0.00649f
C45 B.n17 VSUBS 0.00649f
C46 B.n18 VSUBS 0.00649f
C47 B.n19 VSUBS 0.00649f
C48 B.n20 VSUBS 0.01515f
C49 B.n21 VSUBS 0.00649f
C50 B.n22 VSUBS 0.00649f
C51 B.n23 VSUBS 0.00649f
C52 B.n24 VSUBS 0.00649f
C53 B.n25 VSUBS 0.00649f
C54 B.n26 VSUBS 0.00649f
C55 B.n27 VSUBS 0.00649f
C56 B.n28 VSUBS 0.00649f
C57 B.n29 VSUBS 0.00649f
C58 B.n30 VSUBS 0.00649f
C59 B.n31 VSUBS 0.00649f
C60 B.n32 VSUBS 0.00649f
C61 B.n33 VSUBS 0.00649f
C62 B.n34 VSUBS 0.00649f
C63 B.n35 VSUBS 0.00649f
C64 B.n36 VSUBS 0.00649f
C65 B.n37 VSUBS 0.00649f
C66 B.n38 VSUBS 0.00649f
C67 B.n39 VSUBS 0.00649f
C68 B.t5 VSUBS 0.182709f
C69 B.t4 VSUBS 0.206584f
C70 B.t3 VSUBS 0.961261f
C71 B.n40 VSUBS 0.326577f
C72 B.n41 VSUBS 0.223139f
C73 B.n42 VSUBS 0.015037f
C74 B.n43 VSUBS 0.00649f
C75 B.n44 VSUBS 0.00649f
C76 B.n45 VSUBS 0.00649f
C77 B.n46 VSUBS 0.00649f
C78 B.n47 VSUBS 0.00649f
C79 B.t8 VSUBS 0.182712f
C80 B.t7 VSUBS 0.206587f
C81 B.t6 VSUBS 0.961261f
C82 B.n48 VSUBS 0.326574f
C83 B.n49 VSUBS 0.223136f
C84 B.n50 VSUBS 0.00649f
C85 B.n51 VSUBS 0.00649f
C86 B.n52 VSUBS 0.00649f
C87 B.n53 VSUBS 0.00649f
C88 B.n54 VSUBS 0.00649f
C89 B.n55 VSUBS 0.00649f
C90 B.n56 VSUBS 0.00649f
C91 B.n57 VSUBS 0.00649f
C92 B.n58 VSUBS 0.00649f
C93 B.n59 VSUBS 0.00649f
C94 B.n60 VSUBS 0.00649f
C95 B.n61 VSUBS 0.00649f
C96 B.n62 VSUBS 0.00649f
C97 B.n63 VSUBS 0.00649f
C98 B.n64 VSUBS 0.00649f
C99 B.n65 VSUBS 0.00649f
C100 B.n66 VSUBS 0.00649f
C101 B.n67 VSUBS 0.00649f
C102 B.n68 VSUBS 0.00649f
C103 B.n69 VSUBS 0.014629f
C104 B.n70 VSUBS 0.00649f
C105 B.n71 VSUBS 0.00649f
C106 B.n72 VSUBS 0.00649f
C107 B.n73 VSUBS 0.00649f
C108 B.n74 VSUBS 0.00649f
C109 B.n75 VSUBS 0.00649f
C110 B.n76 VSUBS 0.00649f
C111 B.n77 VSUBS 0.00649f
C112 B.n78 VSUBS 0.00649f
C113 B.n79 VSUBS 0.00649f
C114 B.n80 VSUBS 0.00649f
C115 B.n81 VSUBS 0.00649f
C116 B.n82 VSUBS 0.00649f
C117 B.n83 VSUBS 0.00649f
C118 B.n84 VSUBS 0.00649f
C119 B.n85 VSUBS 0.00649f
C120 B.n86 VSUBS 0.00649f
C121 B.n87 VSUBS 0.00649f
C122 B.n88 VSUBS 0.00649f
C123 B.n89 VSUBS 0.00649f
C124 B.n90 VSUBS 0.00649f
C125 B.n91 VSUBS 0.00649f
C126 B.n92 VSUBS 0.00649f
C127 B.n93 VSUBS 0.00649f
C128 B.n94 VSUBS 0.00649f
C129 B.n95 VSUBS 0.00649f
C130 B.n96 VSUBS 0.00649f
C131 B.n97 VSUBS 0.00649f
C132 B.n98 VSUBS 0.00649f
C133 B.n99 VSUBS 0.00649f
C134 B.n100 VSUBS 0.00649f
C135 B.n101 VSUBS 0.00649f
C136 B.n102 VSUBS 0.00649f
C137 B.n103 VSUBS 0.00649f
C138 B.n104 VSUBS 0.00649f
C139 B.n105 VSUBS 0.014629f
C140 B.n106 VSUBS 0.00649f
C141 B.n107 VSUBS 0.00649f
C142 B.n108 VSUBS 0.00649f
C143 B.n109 VSUBS 0.00649f
C144 B.n110 VSUBS 0.00649f
C145 B.n111 VSUBS 0.00649f
C146 B.n112 VSUBS 0.00649f
C147 B.n113 VSUBS 0.00649f
C148 B.n114 VSUBS 0.00649f
C149 B.n115 VSUBS 0.00649f
C150 B.n116 VSUBS 0.00649f
C151 B.n117 VSUBS 0.00649f
C152 B.n118 VSUBS 0.00649f
C153 B.n119 VSUBS 0.00649f
C154 B.n120 VSUBS 0.00649f
C155 B.n121 VSUBS 0.00649f
C156 B.n122 VSUBS 0.00649f
C157 B.n123 VSUBS 0.00649f
C158 B.n124 VSUBS 0.00649f
C159 B.n125 VSUBS 0.00649f
C160 B.t1 VSUBS 0.182712f
C161 B.t2 VSUBS 0.206587f
C162 B.t0 VSUBS 0.961261f
C163 B.n126 VSUBS 0.326574f
C164 B.n127 VSUBS 0.223136f
C165 B.n128 VSUBS 0.00649f
C166 B.n129 VSUBS 0.00649f
C167 B.n130 VSUBS 0.00649f
C168 B.n131 VSUBS 0.00649f
C169 B.t10 VSUBS 0.182709f
C170 B.t11 VSUBS 0.206584f
C171 B.t9 VSUBS 0.961261f
C172 B.n132 VSUBS 0.326577f
C173 B.n133 VSUBS 0.223139f
C174 B.n134 VSUBS 0.015037f
C175 B.n135 VSUBS 0.00649f
C176 B.n136 VSUBS 0.00649f
C177 B.n137 VSUBS 0.00649f
C178 B.n138 VSUBS 0.00649f
C179 B.n139 VSUBS 0.00649f
C180 B.n140 VSUBS 0.00649f
C181 B.n141 VSUBS 0.00649f
C182 B.n142 VSUBS 0.00649f
C183 B.n143 VSUBS 0.00649f
C184 B.n144 VSUBS 0.00649f
C185 B.n145 VSUBS 0.00649f
C186 B.n146 VSUBS 0.00649f
C187 B.n147 VSUBS 0.00649f
C188 B.n148 VSUBS 0.00649f
C189 B.n149 VSUBS 0.00649f
C190 B.n150 VSUBS 0.00649f
C191 B.n151 VSUBS 0.00649f
C192 B.n152 VSUBS 0.00649f
C193 B.n153 VSUBS 0.00649f
C194 B.n154 VSUBS 0.01515f
C195 B.n155 VSUBS 0.00649f
C196 B.n156 VSUBS 0.00649f
C197 B.n157 VSUBS 0.00649f
C198 B.n158 VSUBS 0.00649f
C199 B.n159 VSUBS 0.00649f
C200 B.n160 VSUBS 0.00649f
C201 B.n161 VSUBS 0.00649f
C202 B.n162 VSUBS 0.00649f
C203 B.n163 VSUBS 0.00649f
C204 B.n164 VSUBS 0.00649f
C205 B.n165 VSUBS 0.00649f
C206 B.n166 VSUBS 0.00649f
C207 B.n167 VSUBS 0.00649f
C208 B.n168 VSUBS 0.00649f
C209 B.n169 VSUBS 0.00649f
C210 B.n170 VSUBS 0.00649f
C211 B.n171 VSUBS 0.00649f
C212 B.n172 VSUBS 0.00649f
C213 B.n173 VSUBS 0.00649f
C214 B.n174 VSUBS 0.00649f
C215 B.n175 VSUBS 0.00649f
C216 B.n176 VSUBS 0.00649f
C217 B.n177 VSUBS 0.00649f
C218 B.n178 VSUBS 0.00649f
C219 B.n179 VSUBS 0.00649f
C220 B.n180 VSUBS 0.00649f
C221 B.n181 VSUBS 0.00649f
C222 B.n182 VSUBS 0.00649f
C223 B.n183 VSUBS 0.00649f
C224 B.n184 VSUBS 0.00649f
C225 B.n185 VSUBS 0.00649f
C226 B.n186 VSUBS 0.00649f
C227 B.n187 VSUBS 0.00649f
C228 B.n188 VSUBS 0.00649f
C229 B.n189 VSUBS 0.00649f
C230 B.n190 VSUBS 0.00649f
C231 B.n191 VSUBS 0.00649f
C232 B.n192 VSUBS 0.00649f
C233 B.n193 VSUBS 0.00649f
C234 B.n194 VSUBS 0.00649f
C235 B.n195 VSUBS 0.00649f
C236 B.n196 VSUBS 0.00649f
C237 B.n197 VSUBS 0.00649f
C238 B.n198 VSUBS 0.00649f
C239 B.n199 VSUBS 0.00649f
C240 B.n200 VSUBS 0.00649f
C241 B.n201 VSUBS 0.00649f
C242 B.n202 VSUBS 0.00649f
C243 B.n203 VSUBS 0.00649f
C244 B.n204 VSUBS 0.00649f
C245 B.n205 VSUBS 0.00649f
C246 B.n206 VSUBS 0.00649f
C247 B.n207 VSUBS 0.00649f
C248 B.n208 VSUBS 0.00649f
C249 B.n209 VSUBS 0.00649f
C250 B.n210 VSUBS 0.00649f
C251 B.n211 VSUBS 0.00649f
C252 B.n212 VSUBS 0.00649f
C253 B.n213 VSUBS 0.00649f
C254 B.n214 VSUBS 0.00649f
C255 B.n215 VSUBS 0.00649f
C256 B.n216 VSUBS 0.00649f
C257 B.n217 VSUBS 0.00649f
C258 B.n218 VSUBS 0.00649f
C259 B.n219 VSUBS 0.00649f
C260 B.n220 VSUBS 0.00649f
C261 B.n221 VSUBS 0.00649f
C262 B.n222 VSUBS 0.00649f
C263 B.n223 VSUBS 0.014629f
C264 B.n224 VSUBS 0.014629f
C265 B.n225 VSUBS 0.01515f
C266 B.n226 VSUBS 0.00649f
C267 B.n227 VSUBS 0.00649f
C268 B.n228 VSUBS 0.00649f
C269 B.n229 VSUBS 0.00649f
C270 B.n230 VSUBS 0.00649f
C271 B.n231 VSUBS 0.00649f
C272 B.n232 VSUBS 0.00649f
C273 B.n233 VSUBS 0.00649f
C274 B.n234 VSUBS 0.00649f
C275 B.n235 VSUBS 0.00649f
C276 B.n236 VSUBS 0.00649f
C277 B.n237 VSUBS 0.00649f
C278 B.n238 VSUBS 0.00649f
C279 B.n239 VSUBS 0.00649f
C280 B.n240 VSUBS 0.00649f
C281 B.n241 VSUBS 0.00649f
C282 B.n242 VSUBS 0.00649f
C283 B.n243 VSUBS 0.00649f
C284 B.n244 VSUBS 0.00649f
C285 B.n245 VSUBS 0.00649f
C286 B.n246 VSUBS 0.00649f
C287 B.n247 VSUBS 0.00649f
C288 B.n248 VSUBS 0.00649f
C289 B.n249 VSUBS 0.00649f
C290 B.n250 VSUBS 0.00649f
C291 B.n251 VSUBS 0.00649f
C292 B.n252 VSUBS 0.00649f
C293 B.n253 VSUBS 0.00649f
C294 B.n254 VSUBS 0.00649f
C295 B.n255 VSUBS 0.00649f
C296 B.n256 VSUBS 0.00649f
C297 B.n257 VSUBS 0.00649f
C298 B.n258 VSUBS 0.00649f
C299 B.n259 VSUBS 0.00649f
C300 B.n260 VSUBS 0.00649f
C301 B.n261 VSUBS 0.00649f
C302 B.n262 VSUBS 0.00649f
C303 B.n263 VSUBS 0.00649f
C304 B.n264 VSUBS 0.00649f
C305 B.n265 VSUBS 0.00649f
C306 B.n266 VSUBS 0.00649f
C307 B.n267 VSUBS 0.00649f
C308 B.n268 VSUBS 0.00649f
C309 B.n269 VSUBS 0.00649f
C310 B.n270 VSUBS 0.00649f
C311 B.n271 VSUBS 0.00649f
C312 B.n272 VSUBS 0.00649f
C313 B.n273 VSUBS 0.00649f
C314 B.n274 VSUBS 0.00649f
C315 B.n275 VSUBS 0.00649f
C316 B.n276 VSUBS 0.00649f
C317 B.n277 VSUBS 0.00649f
C318 B.n278 VSUBS 0.00649f
C319 B.n279 VSUBS 0.00649f
C320 B.n280 VSUBS 0.00649f
C321 B.n281 VSUBS 0.00649f
C322 B.n282 VSUBS 0.00649f
C323 B.n283 VSUBS 0.004486f
C324 B.n284 VSUBS 0.00649f
C325 B.n285 VSUBS 0.00649f
C326 B.n286 VSUBS 0.00525f
C327 B.n287 VSUBS 0.00649f
C328 B.n288 VSUBS 0.00649f
C329 B.n289 VSUBS 0.00649f
C330 B.n290 VSUBS 0.00649f
C331 B.n291 VSUBS 0.00649f
C332 B.n292 VSUBS 0.00649f
C333 B.n293 VSUBS 0.00649f
C334 B.n294 VSUBS 0.00649f
C335 B.n295 VSUBS 0.00649f
C336 B.n296 VSUBS 0.00649f
C337 B.n297 VSUBS 0.00649f
C338 B.n298 VSUBS 0.00525f
C339 B.n299 VSUBS 0.015037f
C340 B.n300 VSUBS 0.004486f
C341 B.n301 VSUBS 0.00649f
C342 B.n302 VSUBS 0.00649f
C343 B.n303 VSUBS 0.00649f
C344 B.n304 VSUBS 0.00649f
C345 B.n305 VSUBS 0.00649f
C346 B.n306 VSUBS 0.00649f
C347 B.n307 VSUBS 0.00649f
C348 B.n308 VSUBS 0.00649f
C349 B.n309 VSUBS 0.00649f
C350 B.n310 VSUBS 0.00649f
C351 B.n311 VSUBS 0.00649f
C352 B.n312 VSUBS 0.00649f
C353 B.n313 VSUBS 0.00649f
C354 B.n314 VSUBS 0.00649f
C355 B.n315 VSUBS 0.00649f
C356 B.n316 VSUBS 0.00649f
C357 B.n317 VSUBS 0.00649f
C358 B.n318 VSUBS 0.00649f
C359 B.n319 VSUBS 0.00649f
C360 B.n320 VSUBS 0.00649f
C361 B.n321 VSUBS 0.00649f
C362 B.n322 VSUBS 0.00649f
C363 B.n323 VSUBS 0.00649f
C364 B.n324 VSUBS 0.00649f
C365 B.n325 VSUBS 0.00649f
C366 B.n326 VSUBS 0.00649f
C367 B.n327 VSUBS 0.00649f
C368 B.n328 VSUBS 0.00649f
C369 B.n329 VSUBS 0.00649f
C370 B.n330 VSUBS 0.00649f
C371 B.n331 VSUBS 0.00649f
C372 B.n332 VSUBS 0.00649f
C373 B.n333 VSUBS 0.00649f
C374 B.n334 VSUBS 0.00649f
C375 B.n335 VSUBS 0.00649f
C376 B.n336 VSUBS 0.00649f
C377 B.n337 VSUBS 0.00649f
C378 B.n338 VSUBS 0.00649f
C379 B.n339 VSUBS 0.00649f
C380 B.n340 VSUBS 0.00649f
C381 B.n341 VSUBS 0.00649f
C382 B.n342 VSUBS 0.00649f
C383 B.n343 VSUBS 0.00649f
C384 B.n344 VSUBS 0.00649f
C385 B.n345 VSUBS 0.00649f
C386 B.n346 VSUBS 0.00649f
C387 B.n347 VSUBS 0.00649f
C388 B.n348 VSUBS 0.00649f
C389 B.n349 VSUBS 0.00649f
C390 B.n350 VSUBS 0.00649f
C391 B.n351 VSUBS 0.00649f
C392 B.n352 VSUBS 0.00649f
C393 B.n353 VSUBS 0.00649f
C394 B.n354 VSUBS 0.00649f
C395 B.n355 VSUBS 0.00649f
C396 B.n356 VSUBS 0.00649f
C397 B.n357 VSUBS 0.00649f
C398 B.n358 VSUBS 0.01515f
C399 B.n359 VSUBS 0.01515f
C400 B.n360 VSUBS 0.014629f
C401 B.n361 VSUBS 0.00649f
C402 B.n362 VSUBS 0.00649f
C403 B.n363 VSUBS 0.00649f
C404 B.n364 VSUBS 0.00649f
C405 B.n365 VSUBS 0.00649f
C406 B.n366 VSUBS 0.00649f
C407 B.n367 VSUBS 0.00649f
C408 B.n368 VSUBS 0.00649f
C409 B.n369 VSUBS 0.00649f
C410 B.n370 VSUBS 0.00649f
C411 B.n371 VSUBS 0.00649f
C412 B.n372 VSUBS 0.00649f
C413 B.n373 VSUBS 0.00649f
C414 B.n374 VSUBS 0.00649f
C415 B.n375 VSUBS 0.00649f
C416 B.n376 VSUBS 0.00649f
C417 B.n377 VSUBS 0.00649f
C418 B.n378 VSUBS 0.00649f
C419 B.n379 VSUBS 0.00649f
C420 B.n380 VSUBS 0.00649f
C421 B.n381 VSUBS 0.00649f
C422 B.n382 VSUBS 0.00649f
C423 B.n383 VSUBS 0.00649f
C424 B.n384 VSUBS 0.00649f
C425 B.n385 VSUBS 0.00649f
C426 B.n386 VSUBS 0.00649f
C427 B.n387 VSUBS 0.00649f
C428 B.n388 VSUBS 0.00649f
C429 B.n389 VSUBS 0.00649f
C430 B.n390 VSUBS 0.00649f
C431 B.n391 VSUBS 0.00649f
C432 B.n392 VSUBS 0.00649f
C433 B.n393 VSUBS 0.00649f
C434 B.n394 VSUBS 0.00649f
C435 B.n395 VSUBS 0.00649f
C436 B.n396 VSUBS 0.00649f
C437 B.n397 VSUBS 0.00649f
C438 B.n398 VSUBS 0.00649f
C439 B.n399 VSUBS 0.00649f
C440 B.n400 VSUBS 0.00649f
C441 B.n401 VSUBS 0.00649f
C442 B.n402 VSUBS 0.00649f
C443 B.n403 VSUBS 0.00649f
C444 B.n404 VSUBS 0.00649f
C445 B.n405 VSUBS 0.00649f
C446 B.n406 VSUBS 0.00649f
C447 B.n407 VSUBS 0.00649f
C448 B.n408 VSUBS 0.00649f
C449 B.n409 VSUBS 0.00649f
C450 B.n410 VSUBS 0.00649f
C451 B.n411 VSUBS 0.00649f
C452 B.n412 VSUBS 0.00649f
C453 B.n413 VSUBS 0.00649f
C454 B.n414 VSUBS 0.00649f
C455 B.n415 VSUBS 0.00649f
C456 B.n416 VSUBS 0.00649f
C457 B.n417 VSUBS 0.00649f
C458 B.n418 VSUBS 0.00649f
C459 B.n419 VSUBS 0.00649f
C460 B.n420 VSUBS 0.00649f
C461 B.n421 VSUBS 0.00649f
C462 B.n422 VSUBS 0.00649f
C463 B.n423 VSUBS 0.00649f
C464 B.n424 VSUBS 0.00649f
C465 B.n425 VSUBS 0.00649f
C466 B.n426 VSUBS 0.00649f
C467 B.n427 VSUBS 0.00649f
C468 B.n428 VSUBS 0.00649f
C469 B.n429 VSUBS 0.00649f
C470 B.n430 VSUBS 0.00649f
C471 B.n431 VSUBS 0.00649f
C472 B.n432 VSUBS 0.00649f
C473 B.n433 VSUBS 0.00649f
C474 B.n434 VSUBS 0.00649f
C475 B.n435 VSUBS 0.00649f
C476 B.n436 VSUBS 0.00649f
C477 B.n437 VSUBS 0.00649f
C478 B.n438 VSUBS 0.00649f
C479 B.n439 VSUBS 0.00649f
C480 B.n440 VSUBS 0.00649f
C481 B.n441 VSUBS 0.00649f
C482 B.n442 VSUBS 0.00649f
C483 B.n443 VSUBS 0.00649f
C484 B.n444 VSUBS 0.00649f
C485 B.n445 VSUBS 0.00649f
C486 B.n446 VSUBS 0.00649f
C487 B.n447 VSUBS 0.00649f
C488 B.n448 VSUBS 0.00649f
C489 B.n449 VSUBS 0.00649f
C490 B.n450 VSUBS 0.00649f
C491 B.n451 VSUBS 0.00649f
C492 B.n452 VSUBS 0.00649f
C493 B.n453 VSUBS 0.00649f
C494 B.n454 VSUBS 0.00649f
C495 B.n455 VSUBS 0.00649f
C496 B.n456 VSUBS 0.00649f
C497 B.n457 VSUBS 0.00649f
C498 B.n458 VSUBS 0.00649f
C499 B.n459 VSUBS 0.00649f
C500 B.n460 VSUBS 0.00649f
C501 B.n461 VSUBS 0.00649f
C502 B.n462 VSUBS 0.00649f
C503 B.n463 VSUBS 0.00649f
C504 B.n464 VSUBS 0.00649f
C505 B.n465 VSUBS 0.00649f
C506 B.n466 VSUBS 0.00649f
C507 B.n467 VSUBS 0.00649f
C508 B.n468 VSUBS 0.01542f
C509 B.n469 VSUBS 0.014359f
C510 B.n470 VSUBS 0.01515f
C511 B.n471 VSUBS 0.00649f
C512 B.n472 VSUBS 0.00649f
C513 B.n473 VSUBS 0.00649f
C514 B.n474 VSUBS 0.00649f
C515 B.n475 VSUBS 0.00649f
C516 B.n476 VSUBS 0.00649f
C517 B.n477 VSUBS 0.00649f
C518 B.n478 VSUBS 0.00649f
C519 B.n479 VSUBS 0.00649f
C520 B.n480 VSUBS 0.00649f
C521 B.n481 VSUBS 0.00649f
C522 B.n482 VSUBS 0.00649f
C523 B.n483 VSUBS 0.00649f
C524 B.n484 VSUBS 0.00649f
C525 B.n485 VSUBS 0.00649f
C526 B.n486 VSUBS 0.00649f
C527 B.n487 VSUBS 0.00649f
C528 B.n488 VSUBS 0.00649f
C529 B.n489 VSUBS 0.00649f
C530 B.n490 VSUBS 0.00649f
C531 B.n491 VSUBS 0.00649f
C532 B.n492 VSUBS 0.00649f
C533 B.n493 VSUBS 0.00649f
C534 B.n494 VSUBS 0.00649f
C535 B.n495 VSUBS 0.00649f
C536 B.n496 VSUBS 0.00649f
C537 B.n497 VSUBS 0.00649f
C538 B.n498 VSUBS 0.00649f
C539 B.n499 VSUBS 0.00649f
C540 B.n500 VSUBS 0.00649f
C541 B.n501 VSUBS 0.00649f
C542 B.n502 VSUBS 0.00649f
C543 B.n503 VSUBS 0.00649f
C544 B.n504 VSUBS 0.00649f
C545 B.n505 VSUBS 0.00649f
C546 B.n506 VSUBS 0.00649f
C547 B.n507 VSUBS 0.00649f
C548 B.n508 VSUBS 0.00649f
C549 B.n509 VSUBS 0.00649f
C550 B.n510 VSUBS 0.00649f
C551 B.n511 VSUBS 0.00649f
C552 B.n512 VSUBS 0.00649f
C553 B.n513 VSUBS 0.00649f
C554 B.n514 VSUBS 0.00649f
C555 B.n515 VSUBS 0.00649f
C556 B.n516 VSUBS 0.00649f
C557 B.n517 VSUBS 0.00649f
C558 B.n518 VSUBS 0.00649f
C559 B.n519 VSUBS 0.00649f
C560 B.n520 VSUBS 0.00649f
C561 B.n521 VSUBS 0.00649f
C562 B.n522 VSUBS 0.00649f
C563 B.n523 VSUBS 0.00649f
C564 B.n524 VSUBS 0.00649f
C565 B.n525 VSUBS 0.00649f
C566 B.n526 VSUBS 0.00649f
C567 B.n527 VSUBS 0.00649f
C568 B.n528 VSUBS 0.004486f
C569 B.n529 VSUBS 0.015037f
C570 B.n530 VSUBS 0.00525f
C571 B.n531 VSUBS 0.00649f
C572 B.n532 VSUBS 0.00649f
C573 B.n533 VSUBS 0.00649f
C574 B.n534 VSUBS 0.00649f
C575 B.n535 VSUBS 0.00649f
C576 B.n536 VSUBS 0.00649f
C577 B.n537 VSUBS 0.00649f
C578 B.n538 VSUBS 0.00649f
C579 B.n539 VSUBS 0.00649f
C580 B.n540 VSUBS 0.00649f
C581 B.n541 VSUBS 0.00649f
C582 B.n542 VSUBS 0.00525f
C583 B.n543 VSUBS 0.00649f
C584 B.n544 VSUBS 0.00649f
C585 B.n545 VSUBS 0.004486f
C586 B.n546 VSUBS 0.00649f
C587 B.n547 VSUBS 0.00649f
C588 B.n548 VSUBS 0.00649f
C589 B.n549 VSUBS 0.00649f
C590 B.n550 VSUBS 0.00649f
C591 B.n551 VSUBS 0.00649f
C592 B.n552 VSUBS 0.00649f
C593 B.n553 VSUBS 0.00649f
C594 B.n554 VSUBS 0.00649f
C595 B.n555 VSUBS 0.00649f
C596 B.n556 VSUBS 0.00649f
C597 B.n557 VSUBS 0.00649f
C598 B.n558 VSUBS 0.00649f
C599 B.n559 VSUBS 0.00649f
C600 B.n560 VSUBS 0.00649f
C601 B.n561 VSUBS 0.00649f
C602 B.n562 VSUBS 0.00649f
C603 B.n563 VSUBS 0.00649f
C604 B.n564 VSUBS 0.00649f
C605 B.n565 VSUBS 0.00649f
C606 B.n566 VSUBS 0.00649f
C607 B.n567 VSUBS 0.00649f
C608 B.n568 VSUBS 0.00649f
C609 B.n569 VSUBS 0.00649f
C610 B.n570 VSUBS 0.00649f
C611 B.n571 VSUBS 0.00649f
C612 B.n572 VSUBS 0.00649f
C613 B.n573 VSUBS 0.00649f
C614 B.n574 VSUBS 0.00649f
C615 B.n575 VSUBS 0.00649f
C616 B.n576 VSUBS 0.00649f
C617 B.n577 VSUBS 0.00649f
C618 B.n578 VSUBS 0.00649f
C619 B.n579 VSUBS 0.00649f
C620 B.n580 VSUBS 0.00649f
C621 B.n581 VSUBS 0.00649f
C622 B.n582 VSUBS 0.00649f
C623 B.n583 VSUBS 0.00649f
C624 B.n584 VSUBS 0.00649f
C625 B.n585 VSUBS 0.00649f
C626 B.n586 VSUBS 0.00649f
C627 B.n587 VSUBS 0.00649f
C628 B.n588 VSUBS 0.00649f
C629 B.n589 VSUBS 0.00649f
C630 B.n590 VSUBS 0.00649f
C631 B.n591 VSUBS 0.00649f
C632 B.n592 VSUBS 0.00649f
C633 B.n593 VSUBS 0.00649f
C634 B.n594 VSUBS 0.00649f
C635 B.n595 VSUBS 0.00649f
C636 B.n596 VSUBS 0.00649f
C637 B.n597 VSUBS 0.00649f
C638 B.n598 VSUBS 0.00649f
C639 B.n599 VSUBS 0.00649f
C640 B.n600 VSUBS 0.00649f
C641 B.n601 VSUBS 0.00649f
C642 B.n602 VSUBS 0.00649f
C643 B.n603 VSUBS 0.01515f
C644 B.n604 VSUBS 0.014629f
C645 B.n605 VSUBS 0.014629f
C646 B.n606 VSUBS 0.00649f
C647 B.n607 VSUBS 0.00649f
C648 B.n608 VSUBS 0.00649f
C649 B.n609 VSUBS 0.00649f
C650 B.n610 VSUBS 0.00649f
C651 B.n611 VSUBS 0.00649f
C652 B.n612 VSUBS 0.00649f
C653 B.n613 VSUBS 0.00649f
C654 B.n614 VSUBS 0.00649f
C655 B.n615 VSUBS 0.00649f
C656 B.n616 VSUBS 0.00649f
C657 B.n617 VSUBS 0.00649f
C658 B.n618 VSUBS 0.00649f
C659 B.n619 VSUBS 0.00649f
C660 B.n620 VSUBS 0.00649f
C661 B.n621 VSUBS 0.00649f
C662 B.n622 VSUBS 0.00649f
C663 B.n623 VSUBS 0.00649f
C664 B.n624 VSUBS 0.00649f
C665 B.n625 VSUBS 0.00649f
C666 B.n626 VSUBS 0.00649f
C667 B.n627 VSUBS 0.00649f
C668 B.n628 VSUBS 0.00649f
C669 B.n629 VSUBS 0.00649f
C670 B.n630 VSUBS 0.00649f
C671 B.n631 VSUBS 0.00649f
C672 B.n632 VSUBS 0.00649f
C673 B.n633 VSUBS 0.00649f
C674 B.n634 VSUBS 0.00649f
C675 B.n635 VSUBS 0.00649f
C676 B.n636 VSUBS 0.00649f
C677 B.n637 VSUBS 0.00649f
C678 B.n638 VSUBS 0.00649f
C679 B.n639 VSUBS 0.00649f
C680 B.n640 VSUBS 0.00649f
C681 B.n641 VSUBS 0.00649f
C682 B.n642 VSUBS 0.00649f
C683 B.n643 VSUBS 0.00649f
C684 B.n644 VSUBS 0.00649f
C685 B.n645 VSUBS 0.00649f
C686 B.n646 VSUBS 0.00649f
C687 B.n647 VSUBS 0.00649f
C688 B.n648 VSUBS 0.00649f
C689 B.n649 VSUBS 0.00649f
C690 B.n650 VSUBS 0.00649f
C691 B.n651 VSUBS 0.00649f
C692 B.n652 VSUBS 0.00649f
C693 B.n653 VSUBS 0.00649f
C694 B.n654 VSUBS 0.00649f
C695 B.n655 VSUBS 0.00649f
C696 B.n656 VSUBS 0.00649f
C697 B.n657 VSUBS 0.00649f
C698 B.n658 VSUBS 0.00649f
C699 B.n659 VSUBS 0.014696f
C700 VDD2.n0 VSUBS 0.026662f
C701 VDD2.n1 VSUBS 0.025036f
C702 VDD2.n2 VSUBS 0.013453f
C703 VDD2.n3 VSUBS 0.031799f
C704 VDD2.n4 VSUBS 0.014245f
C705 VDD2.n5 VSUBS 0.025036f
C706 VDD2.n6 VSUBS 0.013453f
C707 VDD2.n7 VSUBS 0.031799f
C708 VDD2.n8 VSUBS 0.013849f
C709 VDD2.n9 VSUBS 0.025036f
C710 VDD2.n10 VSUBS 0.014245f
C711 VDD2.n11 VSUBS 0.031799f
C712 VDD2.n12 VSUBS 0.014245f
C713 VDD2.n13 VSUBS 0.025036f
C714 VDD2.n14 VSUBS 0.013453f
C715 VDD2.n15 VSUBS 0.031799f
C716 VDD2.n16 VSUBS 0.014245f
C717 VDD2.n17 VSUBS 1.16099f
C718 VDD2.n18 VSUBS 0.013453f
C719 VDD2.t0 VSUBS 0.068472f
C720 VDD2.n19 VSUBS 0.190045f
C721 VDD2.n20 VSUBS 0.023921f
C722 VDD2.n21 VSUBS 0.023849f
C723 VDD2.n22 VSUBS 0.031799f
C724 VDD2.n23 VSUBS 0.014245f
C725 VDD2.n24 VSUBS 0.013453f
C726 VDD2.n25 VSUBS 0.025036f
C727 VDD2.n26 VSUBS 0.025036f
C728 VDD2.n27 VSUBS 0.013453f
C729 VDD2.n28 VSUBS 0.014245f
C730 VDD2.n29 VSUBS 0.031799f
C731 VDD2.n30 VSUBS 0.031799f
C732 VDD2.n31 VSUBS 0.014245f
C733 VDD2.n32 VSUBS 0.013453f
C734 VDD2.n33 VSUBS 0.025036f
C735 VDD2.n34 VSUBS 0.025036f
C736 VDD2.n35 VSUBS 0.013453f
C737 VDD2.n36 VSUBS 0.013453f
C738 VDD2.n37 VSUBS 0.014245f
C739 VDD2.n38 VSUBS 0.031799f
C740 VDD2.n39 VSUBS 0.031799f
C741 VDD2.n40 VSUBS 0.031799f
C742 VDD2.n41 VSUBS 0.013849f
C743 VDD2.n42 VSUBS 0.013453f
C744 VDD2.n43 VSUBS 0.025036f
C745 VDD2.n44 VSUBS 0.025036f
C746 VDD2.n45 VSUBS 0.013453f
C747 VDD2.n46 VSUBS 0.014245f
C748 VDD2.n47 VSUBS 0.031799f
C749 VDD2.n48 VSUBS 0.031799f
C750 VDD2.n49 VSUBS 0.014245f
C751 VDD2.n50 VSUBS 0.013453f
C752 VDD2.n51 VSUBS 0.025036f
C753 VDD2.n52 VSUBS 0.025036f
C754 VDD2.n53 VSUBS 0.013453f
C755 VDD2.n54 VSUBS 0.014245f
C756 VDD2.n55 VSUBS 0.031799f
C757 VDD2.n56 VSUBS 0.074094f
C758 VDD2.n57 VSUBS 0.014245f
C759 VDD2.n58 VSUBS 0.013453f
C760 VDD2.n59 VSUBS 0.056844f
C761 VDD2.n60 VSUBS 0.059322f
C762 VDD2.t4 VSUBS 0.224947f
C763 VDD2.t2 VSUBS 0.224947f
C764 VDD2.n61 VSUBS 1.7408f
C765 VDD2.n62 VSUBS 2.65573f
C766 VDD2.n63 VSUBS 0.026662f
C767 VDD2.n64 VSUBS 0.025036f
C768 VDD2.n65 VSUBS 0.013453f
C769 VDD2.n66 VSUBS 0.031799f
C770 VDD2.n67 VSUBS 0.014245f
C771 VDD2.n68 VSUBS 0.025036f
C772 VDD2.n69 VSUBS 0.013453f
C773 VDD2.n70 VSUBS 0.031799f
C774 VDD2.n71 VSUBS 0.013849f
C775 VDD2.n72 VSUBS 0.025036f
C776 VDD2.n73 VSUBS 0.013849f
C777 VDD2.n74 VSUBS 0.013453f
C778 VDD2.n75 VSUBS 0.031799f
C779 VDD2.n76 VSUBS 0.031799f
C780 VDD2.n77 VSUBS 0.014245f
C781 VDD2.n78 VSUBS 0.025036f
C782 VDD2.n79 VSUBS 0.013453f
C783 VDD2.n80 VSUBS 0.031799f
C784 VDD2.n81 VSUBS 0.014245f
C785 VDD2.n82 VSUBS 1.16099f
C786 VDD2.n83 VSUBS 0.013453f
C787 VDD2.t1 VSUBS 0.068472f
C788 VDD2.n84 VSUBS 0.190045f
C789 VDD2.n85 VSUBS 0.023921f
C790 VDD2.n86 VSUBS 0.023849f
C791 VDD2.n87 VSUBS 0.031799f
C792 VDD2.n88 VSUBS 0.014245f
C793 VDD2.n89 VSUBS 0.013453f
C794 VDD2.n90 VSUBS 0.025036f
C795 VDD2.n91 VSUBS 0.025036f
C796 VDD2.n92 VSUBS 0.013453f
C797 VDD2.n93 VSUBS 0.014245f
C798 VDD2.n94 VSUBS 0.031799f
C799 VDD2.n95 VSUBS 0.031799f
C800 VDD2.n96 VSUBS 0.014245f
C801 VDD2.n97 VSUBS 0.013453f
C802 VDD2.n98 VSUBS 0.025036f
C803 VDD2.n99 VSUBS 0.025036f
C804 VDD2.n100 VSUBS 0.013453f
C805 VDD2.n101 VSUBS 0.014245f
C806 VDD2.n102 VSUBS 0.031799f
C807 VDD2.n103 VSUBS 0.031799f
C808 VDD2.n104 VSUBS 0.014245f
C809 VDD2.n105 VSUBS 0.013453f
C810 VDD2.n106 VSUBS 0.025036f
C811 VDD2.n107 VSUBS 0.025036f
C812 VDD2.n108 VSUBS 0.013453f
C813 VDD2.n109 VSUBS 0.014245f
C814 VDD2.n110 VSUBS 0.031799f
C815 VDD2.n111 VSUBS 0.031799f
C816 VDD2.n112 VSUBS 0.014245f
C817 VDD2.n113 VSUBS 0.013453f
C818 VDD2.n114 VSUBS 0.025036f
C819 VDD2.n115 VSUBS 0.025036f
C820 VDD2.n116 VSUBS 0.013453f
C821 VDD2.n117 VSUBS 0.014245f
C822 VDD2.n118 VSUBS 0.031799f
C823 VDD2.n119 VSUBS 0.074094f
C824 VDD2.n120 VSUBS 0.014245f
C825 VDD2.n121 VSUBS 0.013453f
C826 VDD2.n122 VSUBS 0.056844f
C827 VDD2.n123 VSUBS 0.054396f
C828 VDD2.n124 VSUBS 2.35983f
C829 VDD2.t5 VSUBS 0.224947f
C830 VDD2.t3 VSUBS 0.224947f
C831 VDD2.n125 VSUBS 1.74076f
C832 VN.n0 VSUBS 0.046519f
C833 VN.t3 VSUBS 2.21543f
C834 VN.n1 VSUBS 0.044626f
C835 VN.t5 VSUBS 2.41058f
C836 VN.n2 VSUBS 0.870297f
C837 VN.t1 VSUBS 2.21543f
C838 VN.n3 VSUBS 0.897068f
C839 VN.n4 VSUBS 0.065761f
C840 VN.n5 VSUBS 0.294816f
C841 VN.n6 VSUBS 0.035284f
C842 VN.n7 VSUBS 0.035284f
C843 VN.n8 VSUBS 0.058392f
C844 VN.n9 VSUBS 0.056671f
C845 VN.n10 VSUBS 0.898473f
C846 VN.n11 VSUBS 0.045156f
C847 VN.n12 VSUBS 0.046519f
C848 VN.t4 VSUBS 2.21543f
C849 VN.n13 VSUBS 0.044626f
C850 VN.t2 VSUBS 2.41058f
C851 VN.n14 VSUBS 0.870297f
C852 VN.t0 VSUBS 2.21543f
C853 VN.n15 VSUBS 0.897068f
C854 VN.n16 VSUBS 0.065761f
C855 VN.n17 VSUBS 0.294816f
C856 VN.n18 VSUBS 0.035284f
C857 VN.n19 VSUBS 0.035284f
C858 VN.n20 VSUBS 0.058392f
C859 VN.n21 VSUBS 0.056671f
C860 VN.n22 VSUBS 0.898473f
C861 VN.n23 VSUBS 1.736f
C862 VDD1.n0 VSUBS 0.026674f
C863 VDD1.n1 VSUBS 0.025048f
C864 VDD1.n2 VSUBS 0.01346f
C865 VDD1.n3 VSUBS 0.031814f
C866 VDD1.n4 VSUBS 0.014251f
C867 VDD1.n5 VSUBS 0.025048f
C868 VDD1.n6 VSUBS 0.01346f
C869 VDD1.n7 VSUBS 0.031814f
C870 VDD1.n8 VSUBS 0.013856f
C871 VDD1.n9 VSUBS 0.025048f
C872 VDD1.n10 VSUBS 0.013856f
C873 VDD1.n11 VSUBS 0.01346f
C874 VDD1.n12 VSUBS 0.031814f
C875 VDD1.n13 VSUBS 0.031814f
C876 VDD1.n14 VSUBS 0.014251f
C877 VDD1.n15 VSUBS 0.025048f
C878 VDD1.n16 VSUBS 0.01346f
C879 VDD1.n17 VSUBS 0.031814f
C880 VDD1.n18 VSUBS 0.014251f
C881 VDD1.n19 VSUBS 1.16154f
C882 VDD1.n20 VSUBS 0.01346f
C883 VDD1.t4 VSUBS 0.068505f
C884 VDD1.n21 VSUBS 0.190135f
C885 VDD1.n22 VSUBS 0.023932f
C886 VDD1.n23 VSUBS 0.02386f
C887 VDD1.n24 VSUBS 0.031814f
C888 VDD1.n25 VSUBS 0.014251f
C889 VDD1.n26 VSUBS 0.01346f
C890 VDD1.n27 VSUBS 0.025048f
C891 VDD1.n28 VSUBS 0.025048f
C892 VDD1.n29 VSUBS 0.01346f
C893 VDD1.n30 VSUBS 0.014251f
C894 VDD1.n31 VSUBS 0.031814f
C895 VDD1.n32 VSUBS 0.031814f
C896 VDD1.n33 VSUBS 0.014251f
C897 VDD1.n34 VSUBS 0.01346f
C898 VDD1.n35 VSUBS 0.025048f
C899 VDD1.n36 VSUBS 0.025048f
C900 VDD1.n37 VSUBS 0.01346f
C901 VDD1.n38 VSUBS 0.014251f
C902 VDD1.n39 VSUBS 0.031814f
C903 VDD1.n40 VSUBS 0.031814f
C904 VDD1.n41 VSUBS 0.014251f
C905 VDD1.n42 VSUBS 0.01346f
C906 VDD1.n43 VSUBS 0.025048f
C907 VDD1.n44 VSUBS 0.025048f
C908 VDD1.n45 VSUBS 0.01346f
C909 VDD1.n46 VSUBS 0.014251f
C910 VDD1.n47 VSUBS 0.031814f
C911 VDD1.n48 VSUBS 0.031814f
C912 VDD1.n49 VSUBS 0.014251f
C913 VDD1.n50 VSUBS 0.01346f
C914 VDD1.n51 VSUBS 0.025048f
C915 VDD1.n52 VSUBS 0.025048f
C916 VDD1.n53 VSUBS 0.01346f
C917 VDD1.n54 VSUBS 0.014251f
C918 VDD1.n55 VSUBS 0.031814f
C919 VDD1.n56 VSUBS 0.074129f
C920 VDD1.n57 VSUBS 0.014251f
C921 VDD1.n58 VSUBS 0.01346f
C922 VDD1.n59 VSUBS 0.056871f
C923 VDD1.n60 VSUBS 0.059997f
C924 VDD1.n61 VSUBS 0.026674f
C925 VDD1.n62 VSUBS 0.025048f
C926 VDD1.n63 VSUBS 0.01346f
C927 VDD1.n64 VSUBS 0.031814f
C928 VDD1.n65 VSUBS 0.014251f
C929 VDD1.n66 VSUBS 0.025048f
C930 VDD1.n67 VSUBS 0.01346f
C931 VDD1.n68 VSUBS 0.031814f
C932 VDD1.n69 VSUBS 0.013856f
C933 VDD1.n70 VSUBS 0.025048f
C934 VDD1.n71 VSUBS 0.014251f
C935 VDD1.n72 VSUBS 0.031814f
C936 VDD1.n73 VSUBS 0.014251f
C937 VDD1.n74 VSUBS 0.025048f
C938 VDD1.n75 VSUBS 0.01346f
C939 VDD1.n76 VSUBS 0.031814f
C940 VDD1.n77 VSUBS 0.014251f
C941 VDD1.n78 VSUBS 1.16154f
C942 VDD1.n79 VSUBS 0.01346f
C943 VDD1.t2 VSUBS 0.068505f
C944 VDD1.n80 VSUBS 0.190135f
C945 VDD1.n81 VSUBS 0.023932f
C946 VDD1.n82 VSUBS 0.02386f
C947 VDD1.n83 VSUBS 0.031814f
C948 VDD1.n84 VSUBS 0.014251f
C949 VDD1.n85 VSUBS 0.01346f
C950 VDD1.n86 VSUBS 0.025048f
C951 VDD1.n87 VSUBS 0.025048f
C952 VDD1.n88 VSUBS 0.01346f
C953 VDD1.n89 VSUBS 0.014251f
C954 VDD1.n90 VSUBS 0.031814f
C955 VDD1.n91 VSUBS 0.031814f
C956 VDD1.n92 VSUBS 0.014251f
C957 VDD1.n93 VSUBS 0.01346f
C958 VDD1.n94 VSUBS 0.025048f
C959 VDD1.n95 VSUBS 0.025048f
C960 VDD1.n96 VSUBS 0.01346f
C961 VDD1.n97 VSUBS 0.01346f
C962 VDD1.n98 VSUBS 0.014251f
C963 VDD1.n99 VSUBS 0.031814f
C964 VDD1.n100 VSUBS 0.031814f
C965 VDD1.n101 VSUBS 0.031814f
C966 VDD1.n102 VSUBS 0.013856f
C967 VDD1.n103 VSUBS 0.01346f
C968 VDD1.n104 VSUBS 0.025048f
C969 VDD1.n105 VSUBS 0.025048f
C970 VDD1.n106 VSUBS 0.01346f
C971 VDD1.n107 VSUBS 0.014251f
C972 VDD1.n108 VSUBS 0.031814f
C973 VDD1.n109 VSUBS 0.031814f
C974 VDD1.n110 VSUBS 0.014251f
C975 VDD1.n111 VSUBS 0.01346f
C976 VDD1.n112 VSUBS 0.025048f
C977 VDD1.n113 VSUBS 0.025048f
C978 VDD1.n114 VSUBS 0.01346f
C979 VDD1.n115 VSUBS 0.014251f
C980 VDD1.n116 VSUBS 0.031814f
C981 VDD1.n117 VSUBS 0.074129f
C982 VDD1.n118 VSUBS 0.014251f
C983 VDD1.n119 VSUBS 0.01346f
C984 VDD1.n120 VSUBS 0.056871f
C985 VDD1.n121 VSUBS 0.05935f
C986 VDD1.t3 VSUBS 0.225054f
C987 VDD1.t1 VSUBS 0.225054f
C988 VDD1.n122 VSUBS 1.74162f
C989 VDD1.n123 VSUBS 2.76624f
C990 VDD1.t0 VSUBS 0.225054f
C991 VDD1.t5 VSUBS 0.225054f
C992 VDD1.n124 VSUBS 1.73749f
C993 VDD1.n125 VSUBS 2.84702f
C994 VTAIL.t0 VSUBS 0.25906f
C995 VTAIL.t5 VSUBS 0.25906f
C996 VTAIL.n0 VSUBS 1.84553f
C997 VTAIL.n1 VSUBS 0.844456f
C998 VTAIL.n2 VSUBS 0.030705f
C999 VTAIL.n3 VSUBS 0.028833f
C1000 VTAIL.n4 VSUBS 0.015494f
C1001 VTAIL.n5 VSUBS 0.036621f
C1002 VTAIL.n6 VSUBS 0.016405f
C1003 VTAIL.n7 VSUBS 0.028833f
C1004 VTAIL.n8 VSUBS 0.015494f
C1005 VTAIL.n9 VSUBS 0.036621f
C1006 VTAIL.n10 VSUBS 0.015949f
C1007 VTAIL.n11 VSUBS 0.028833f
C1008 VTAIL.n12 VSUBS 0.016405f
C1009 VTAIL.n13 VSUBS 0.036621f
C1010 VTAIL.n14 VSUBS 0.016405f
C1011 VTAIL.n15 VSUBS 0.028833f
C1012 VTAIL.n16 VSUBS 0.015494f
C1013 VTAIL.n17 VSUBS 0.036621f
C1014 VTAIL.n18 VSUBS 0.016405f
C1015 VTAIL.n19 VSUBS 1.33705f
C1016 VTAIL.n20 VSUBS 0.015494f
C1017 VTAIL.t8 VSUBS 0.078856f
C1018 VTAIL.n21 VSUBS 0.218864f
C1019 VTAIL.n22 VSUBS 0.027548f
C1020 VTAIL.n23 VSUBS 0.027466f
C1021 VTAIL.n24 VSUBS 0.036621f
C1022 VTAIL.n25 VSUBS 0.016405f
C1023 VTAIL.n26 VSUBS 0.015494f
C1024 VTAIL.n27 VSUBS 0.028833f
C1025 VTAIL.n28 VSUBS 0.028833f
C1026 VTAIL.n29 VSUBS 0.015494f
C1027 VTAIL.n30 VSUBS 0.016405f
C1028 VTAIL.n31 VSUBS 0.036621f
C1029 VTAIL.n32 VSUBS 0.036621f
C1030 VTAIL.n33 VSUBS 0.016405f
C1031 VTAIL.n34 VSUBS 0.015494f
C1032 VTAIL.n35 VSUBS 0.028833f
C1033 VTAIL.n36 VSUBS 0.028833f
C1034 VTAIL.n37 VSUBS 0.015494f
C1035 VTAIL.n38 VSUBS 0.015494f
C1036 VTAIL.n39 VSUBS 0.016405f
C1037 VTAIL.n40 VSUBS 0.036621f
C1038 VTAIL.n41 VSUBS 0.036621f
C1039 VTAIL.n42 VSUBS 0.036621f
C1040 VTAIL.n43 VSUBS 0.015949f
C1041 VTAIL.n44 VSUBS 0.015494f
C1042 VTAIL.n45 VSUBS 0.028833f
C1043 VTAIL.n46 VSUBS 0.028833f
C1044 VTAIL.n47 VSUBS 0.015494f
C1045 VTAIL.n48 VSUBS 0.016405f
C1046 VTAIL.n49 VSUBS 0.036621f
C1047 VTAIL.n50 VSUBS 0.036621f
C1048 VTAIL.n51 VSUBS 0.016405f
C1049 VTAIL.n52 VSUBS 0.015494f
C1050 VTAIL.n53 VSUBS 0.028833f
C1051 VTAIL.n54 VSUBS 0.028833f
C1052 VTAIL.n55 VSUBS 0.015494f
C1053 VTAIL.n56 VSUBS 0.016405f
C1054 VTAIL.n57 VSUBS 0.036621f
C1055 VTAIL.n58 VSUBS 0.08533f
C1056 VTAIL.n59 VSUBS 0.016405f
C1057 VTAIL.n60 VSUBS 0.015494f
C1058 VTAIL.n61 VSUBS 0.065464f
C1059 VTAIL.n62 VSUBS 0.042728f
C1060 VTAIL.n63 VSUBS 0.351131f
C1061 VTAIL.t6 VSUBS 0.25906f
C1062 VTAIL.t9 VSUBS 0.25906f
C1063 VTAIL.n64 VSUBS 1.84553f
C1064 VTAIL.n65 VSUBS 2.52298f
C1065 VTAIL.t4 VSUBS 0.25906f
C1066 VTAIL.t3 VSUBS 0.25906f
C1067 VTAIL.n66 VSUBS 1.84555f
C1068 VTAIL.n67 VSUBS 2.52297f
C1069 VTAIL.n68 VSUBS 0.030705f
C1070 VTAIL.n69 VSUBS 0.028833f
C1071 VTAIL.n70 VSUBS 0.015494f
C1072 VTAIL.n71 VSUBS 0.036621f
C1073 VTAIL.n72 VSUBS 0.016405f
C1074 VTAIL.n73 VSUBS 0.028833f
C1075 VTAIL.n74 VSUBS 0.015494f
C1076 VTAIL.n75 VSUBS 0.036621f
C1077 VTAIL.n76 VSUBS 0.015949f
C1078 VTAIL.n77 VSUBS 0.028833f
C1079 VTAIL.n78 VSUBS 0.015949f
C1080 VTAIL.n79 VSUBS 0.015494f
C1081 VTAIL.n80 VSUBS 0.036621f
C1082 VTAIL.n81 VSUBS 0.036621f
C1083 VTAIL.n82 VSUBS 0.016405f
C1084 VTAIL.n83 VSUBS 0.028833f
C1085 VTAIL.n84 VSUBS 0.015494f
C1086 VTAIL.n85 VSUBS 0.036621f
C1087 VTAIL.n86 VSUBS 0.016405f
C1088 VTAIL.n87 VSUBS 1.33705f
C1089 VTAIL.n88 VSUBS 0.015494f
C1090 VTAIL.t1 VSUBS 0.078856f
C1091 VTAIL.n89 VSUBS 0.218864f
C1092 VTAIL.n90 VSUBS 0.027548f
C1093 VTAIL.n91 VSUBS 0.027466f
C1094 VTAIL.n92 VSUBS 0.036621f
C1095 VTAIL.n93 VSUBS 0.016405f
C1096 VTAIL.n94 VSUBS 0.015494f
C1097 VTAIL.n95 VSUBS 0.028833f
C1098 VTAIL.n96 VSUBS 0.028833f
C1099 VTAIL.n97 VSUBS 0.015494f
C1100 VTAIL.n98 VSUBS 0.016405f
C1101 VTAIL.n99 VSUBS 0.036621f
C1102 VTAIL.n100 VSUBS 0.036621f
C1103 VTAIL.n101 VSUBS 0.016405f
C1104 VTAIL.n102 VSUBS 0.015494f
C1105 VTAIL.n103 VSUBS 0.028833f
C1106 VTAIL.n104 VSUBS 0.028833f
C1107 VTAIL.n105 VSUBS 0.015494f
C1108 VTAIL.n106 VSUBS 0.016405f
C1109 VTAIL.n107 VSUBS 0.036621f
C1110 VTAIL.n108 VSUBS 0.036621f
C1111 VTAIL.n109 VSUBS 0.016405f
C1112 VTAIL.n110 VSUBS 0.015494f
C1113 VTAIL.n111 VSUBS 0.028833f
C1114 VTAIL.n112 VSUBS 0.028833f
C1115 VTAIL.n113 VSUBS 0.015494f
C1116 VTAIL.n114 VSUBS 0.016405f
C1117 VTAIL.n115 VSUBS 0.036621f
C1118 VTAIL.n116 VSUBS 0.036621f
C1119 VTAIL.n117 VSUBS 0.016405f
C1120 VTAIL.n118 VSUBS 0.015494f
C1121 VTAIL.n119 VSUBS 0.028833f
C1122 VTAIL.n120 VSUBS 0.028833f
C1123 VTAIL.n121 VSUBS 0.015494f
C1124 VTAIL.n122 VSUBS 0.016405f
C1125 VTAIL.n123 VSUBS 0.036621f
C1126 VTAIL.n124 VSUBS 0.08533f
C1127 VTAIL.n125 VSUBS 0.016405f
C1128 VTAIL.n126 VSUBS 0.015494f
C1129 VTAIL.n127 VSUBS 0.065464f
C1130 VTAIL.n128 VSUBS 0.042728f
C1131 VTAIL.n129 VSUBS 0.351131f
C1132 VTAIL.t7 VSUBS 0.25906f
C1133 VTAIL.t10 VSUBS 0.25906f
C1134 VTAIL.n130 VSUBS 1.84555f
C1135 VTAIL.n131 VSUBS 0.980798f
C1136 VTAIL.n132 VSUBS 0.030705f
C1137 VTAIL.n133 VSUBS 0.028833f
C1138 VTAIL.n134 VSUBS 0.015494f
C1139 VTAIL.n135 VSUBS 0.036621f
C1140 VTAIL.n136 VSUBS 0.016405f
C1141 VTAIL.n137 VSUBS 0.028833f
C1142 VTAIL.n138 VSUBS 0.015494f
C1143 VTAIL.n139 VSUBS 0.036621f
C1144 VTAIL.n140 VSUBS 0.015949f
C1145 VTAIL.n141 VSUBS 0.028833f
C1146 VTAIL.n142 VSUBS 0.015949f
C1147 VTAIL.n143 VSUBS 0.015494f
C1148 VTAIL.n144 VSUBS 0.036621f
C1149 VTAIL.n145 VSUBS 0.036621f
C1150 VTAIL.n146 VSUBS 0.016405f
C1151 VTAIL.n147 VSUBS 0.028833f
C1152 VTAIL.n148 VSUBS 0.015494f
C1153 VTAIL.n149 VSUBS 0.036621f
C1154 VTAIL.n150 VSUBS 0.016405f
C1155 VTAIL.n151 VSUBS 1.33705f
C1156 VTAIL.n152 VSUBS 0.015494f
C1157 VTAIL.t11 VSUBS 0.078856f
C1158 VTAIL.n153 VSUBS 0.218864f
C1159 VTAIL.n154 VSUBS 0.027548f
C1160 VTAIL.n155 VSUBS 0.027466f
C1161 VTAIL.n156 VSUBS 0.036621f
C1162 VTAIL.n157 VSUBS 0.016405f
C1163 VTAIL.n158 VSUBS 0.015494f
C1164 VTAIL.n159 VSUBS 0.028833f
C1165 VTAIL.n160 VSUBS 0.028833f
C1166 VTAIL.n161 VSUBS 0.015494f
C1167 VTAIL.n162 VSUBS 0.016405f
C1168 VTAIL.n163 VSUBS 0.036621f
C1169 VTAIL.n164 VSUBS 0.036621f
C1170 VTAIL.n165 VSUBS 0.016405f
C1171 VTAIL.n166 VSUBS 0.015494f
C1172 VTAIL.n167 VSUBS 0.028833f
C1173 VTAIL.n168 VSUBS 0.028833f
C1174 VTAIL.n169 VSUBS 0.015494f
C1175 VTAIL.n170 VSUBS 0.016405f
C1176 VTAIL.n171 VSUBS 0.036621f
C1177 VTAIL.n172 VSUBS 0.036621f
C1178 VTAIL.n173 VSUBS 0.016405f
C1179 VTAIL.n174 VSUBS 0.015494f
C1180 VTAIL.n175 VSUBS 0.028833f
C1181 VTAIL.n176 VSUBS 0.028833f
C1182 VTAIL.n177 VSUBS 0.015494f
C1183 VTAIL.n178 VSUBS 0.016405f
C1184 VTAIL.n179 VSUBS 0.036621f
C1185 VTAIL.n180 VSUBS 0.036621f
C1186 VTAIL.n181 VSUBS 0.016405f
C1187 VTAIL.n182 VSUBS 0.015494f
C1188 VTAIL.n183 VSUBS 0.028833f
C1189 VTAIL.n184 VSUBS 0.028833f
C1190 VTAIL.n185 VSUBS 0.015494f
C1191 VTAIL.n186 VSUBS 0.016405f
C1192 VTAIL.n187 VSUBS 0.036621f
C1193 VTAIL.n188 VSUBS 0.08533f
C1194 VTAIL.n189 VSUBS 0.016405f
C1195 VTAIL.n190 VSUBS 0.015494f
C1196 VTAIL.n191 VSUBS 0.065464f
C1197 VTAIL.n192 VSUBS 0.042728f
C1198 VTAIL.n193 VSUBS 1.70428f
C1199 VTAIL.n194 VSUBS 0.030705f
C1200 VTAIL.n195 VSUBS 0.028833f
C1201 VTAIL.n196 VSUBS 0.015494f
C1202 VTAIL.n197 VSUBS 0.036621f
C1203 VTAIL.n198 VSUBS 0.016405f
C1204 VTAIL.n199 VSUBS 0.028833f
C1205 VTAIL.n200 VSUBS 0.015494f
C1206 VTAIL.n201 VSUBS 0.036621f
C1207 VTAIL.n202 VSUBS 0.015949f
C1208 VTAIL.n203 VSUBS 0.028833f
C1209 VTAIL.n204 VSUBS 0.016405f
C1210 VTAIL.n205 VSUBS 0.036621f
C1211 VTAIL.n206 VSUBS 0.016405f
C1212 VTAIL.n207 VSUBS 0.028833f
C1213 VTAIL.n208 VSUBS 0.015494f
C1214 VTAIL.n209 VSUBS 0.036621f
C1215 VTAIL.n210 VSUBS 0.016405f
C1216 VTAIL.n211 VSUBS 1.33705f
C1217 VTAIL.n212 VSUBS 0.015494f
C1218 VTAIL.t2 VSUBS 0.078856f
C1219 VTAIL.n213 VSUBS 0.218864f
C1220 VTAIL.n214 VSUBS 0.027548f
C1221 VTAIL.n215 VSUBS 0.027466f
C1222 VTAIL.n216 VSUBS 0.036621f
C1223 VTAIL.n217 VSUBS 0.016405f
C1224 VTAIL.n218 VSUBS 0.015494f
C1225 VTAIL.n219 VSUBS 0.028833f
C1226 VTAIL.n220 VSUBS 0.028833f
C1227 VTAIL.n221 VSUBS 0.015494f
C1228 VTAIL.n222 VSUBS 0.016405f
C1229 VTAIL.n223 VSUBS 0.036621f
C1230 VTAIL.n224 VSUBS 0.036621f
C1231 VTAIL.n225 VSUBS 0.016405f
C1232 VTAIL.n226 VSUBS 0.015494f
C1233 VTAIL.n227 VSUBS 0.028833f
C1234 VTAIL.n228 VSUBS 0.028833f
C1235 VTAIL.n229 VSUBS 0.015494f
C1236 VTAIL.n230 VSUBS 0.015494f
C1237 VTAIL.n231 VSUBS 0.016405f
C1238 VTAIL.n232 VSUBS 0.036621f
C1239 VTAIL.n233 VSUBS 0.036621f
C1240 VTAIL.n234 VSUBS 0.036621f
C1241 VTAIL.n235 VSUBS 0.015949f
C1242 VTAIL.n236 VSUBS 0.015494f
C1243 VTAIL.n237 VSUBS 0.028833f
C1244 VTAIL.n238 VSUBS 0.028833f
C1245 VTAIL.n239 VSUBS 0.015494f
C1246 VTAIL.n240 VSUBS 0.016405f
C1247 VTAIL.n241 VSUBS 0.036621f
C1248 VTAIL.n242 VSUBS 0.036621f
C1249 VTAIL.n243 VSUBS 0.016405f
C1250 VTAIL.n244 VSUBS 0.015494f
C1251 VTAIL.n245 VSUBS 0.028833f
C1252 VTAIL.n246 VSUBS 0.028833f
C1253 VTAIL.n247 VSUBS 0.015494f
C1254 VTAIL.n248 VSUBS 0.016405f
C1255 VTAIL.n249 VSUBS 0.036621f
C1256 VTAIL.n250 VSUBS 0.08533f
C1257 VTAIL.n251 VSUBS 0.016405f
C1258 VTAIL.n252 VSUBS 0.015494f
C1259 VTAIL.n253 VSUBS 0.065464f
C1260 VTAIL.n254 VSUBS 0.042728f
C1261 VTAIL.n255 VSUBS 1.65162f
C1262 VP.n0 VSUBS 0.047596f
C1263 VP.t4 VSUBS 2.2667f
C1264 VP.n1 VSUBS 0.045659f
C1265 VP.n2 VSUBS 0.036101f
C1266 VP.t2 VSUBS 2.2667f
C1267 VP.n3 VSUBS 0.045659f
C1268 VP.n4 VSUBS 0.047596f
C1269 VP.t3 VSUBS 2.2667f
C1270 VP.n5 VSUBS 0.047596f
C1271 VP.t0 VSUBS 2.2667f
C1272 VP.n6 VSUBS 0.045659f
C1273 VP.t1 VSUBS 2.46636f
C1274 VP.n7 VSUBS 0.890436f
C1275 VP.t5 VSUBS 2.2667f
C1276 VP.n8 VSUBS 0.917827f
C1277 VP.n9 VSUBS 0.067283f
C1278 VP.n10 VSUBS 0.301638f
C1279 VP.n11 VSUBS 0.036101f
C1280 VP.n12 VSUBS 0.036101f
C1281 VP.n13 VSUBS 0.059743f
C1282 VP.n14 VSUBS 0.057982f
C1283 VP.n15 VSUBS 0.919265f
C1284 VP.n16 VSUBS 1.7565f
C1285 VP.n17 VSUBS 1.78473f
C1286 VP.n18 VSUBS 0.919265f
C1287 VP.n19 VSUBS 0.057982f
C1288 VP.n20 VSUBS 0.059743f
C1289 VP.n21 VSUBS 0.036101f
C1290 VP.n22 VSUBS 0.036101f
C1291 VP.n23 VSUBS 0.036101f
C1292 VP.n24 VSUBS 0.067283f
C1293 VP.n25 VSUBS 0.845668f
C1294 VP.n26 VSUBS 0.067283f
C1295 VP.n27 VSUBS 0.036101f
C1296 VP.n28 VSUBS 0.036101f
C1297 VP.n29 VSUBS 0.036101f
C1298 VP.n30 VSUBS 0.059743f
C1299 VP.n31 VSUBS 0.057982f
C1300 VP.n32 VSUBS 0.919265f
C1301 VP.n33 VSUBS 0.046201f
.ends

