* NGSPICE file created from diff_pair_sample_0312.ext - technology: sky130A

.subckt diff_pair_sample_0312 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=0 ps=0 w=17.32 l=0.76
X1 VTAIL.t7 VP.t0 VDD1.t1 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=2.8578 ps=17.65 w=17.32 l=0.76
X2 VTAIL.t6 VP.t1 VDD1.t0 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=2.8578 ps=17.65 w=17.32 l=0.76
X3 VDD1.t2 VP.t2 VTAIL.t5 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=2.8578 pd=17.65 as=6.7548 ps=35.42 w=17.32 l=0.76
X4 B.t8 B.t6 B.t7 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=0 ps=0 w=17.32 l=0.76
X5 VDD2.t3 VN.t0 VTAIL.t3 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=2.8578 pd=17.65 as=6.7548 ps=35.42 w=17.32 l=0.76
X6 VTAIL.t0 VN.t1 VDD2.t2 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=2.8578 ps=17.65 w=17.32 l=0.76
X7 VDD2.t1 VN.t2 VTAIL.t1 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=2.8578 pd=17.65 as=6.7548 ps=35.42 w=17.32 l=0.76
X8 VDD1.t3 VP.t3 VTAIL.t4 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=2.8578 pd=17.65 as=6.7548 ps=35.42 w=17.32 l=0.76
X9 B.t5 B.t3 B.t4 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=0 ps=0 w=17.32 l=0.76
X10 VTAIL.t2 VN.t3 VDD2.t0 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=2.8578 ps=17.65 w=17.32 l=0.76
X11 B.t2 B.t0 B.t1 w_n1624_n4432# sky130_fd_pr__pfet_01v8 ad=6.7548 pd=35.42 as=0 ps=0 w=17.32 l=0.76
R0 B.n275 B.t3 751.511
R1 B.n124 B.t0 751.511
R2 B.n46 B.t6 751.511
R3 B.n40 B.t9 751.511
R4 B.n380 B.n95 585
R5 B.n379 B.n378 585
R6 B.n377 B.n96 585
R7 B.n376 B.n375 585
R8 B.n374 B.n97 585
R9 B.n373 B.n372 585
R10 B.n371 B.n98 585
R11 B.n370 B.n369 585
R12 B.n368 B.n99 585
R13 B.n367 B.n366 585
R14 B.n365 B.n100 585
R15 B.n364 B.n363 585
R16 B.n362 B.n101 585
R17 B.n361 B.n360 585
R18 B.n359 B.n102 585
R19 B.n358 B.n357 585
R20 B.n356 B.n103 585
R21 B.n355 B.n354 585
R22 B.n353 B.n104 585
R23 B.n352 B.n351 585
R24 B.n350 B.n105 585
R25 B.n349 B.n348 585
R26 B.n347 B.n106 585
R27 B.n346 B.n345 585
R28 B.n344 B.n107 585
R29 B.n343 B.n342 585
R30 B.n341 B.n108 585
R31 B.n340 B.n339 585
R32 B.n338 B.n109 585
R33 B.n337 B.n336 585
R34 B.n335 B.n110 585
R35 B.n334 B.n333 585
R36 B.n332 B.n111 585
R37 B.n331 B.n330 585
R38 B.n329 B.n112 585
R39 B.n328 B.n327 585
R40 B.n326 B.n113 585
R41 B.n325 B.n324 585
R42 B.n323 B.n114 585
R43 B.n322 B.n321 585
R44 B.n320 B.n115 585
R45 B.n319 B.n318 585
R46 B.n317 B.n116 585
R47 B.n316 B.n315 585
R48 B.n314 B.n117 585
R49 B.n313 B.n312 585
R50 B.n311 B.n118 585
R51 B.n310 B.n309 585
R52 B.n308 B.n119 585
R53 B.n307 B.n306 585
R54 B.n305 B.n120 585
R55 B.n304 B.n303 585
R56 B.n302 B.n121 585
R57 B.n301 B.n300 585
R58 B.n299 B.n122 585
R59 B.n298 B.n297 585
R60 B.n296 B.n123 585
R61 B.n294 B.n293 585
R62 B.n292 B.n126 585
R63 B.n291 B.n290 585
R64 B.n289 B.n127 585
R65 B.n288 B.n287 585
R66 B.n286 B.n128 585
R67 B.n285 B.n284 585
R68 B.n283 B.n129 585
R69 B.n282 B.n281 585
R70 B.n280 B.n130 585
R71 B.n279 B.n278 585
R72 B.n274 B.n131 585
R73 B.n273 B.n272 585
R74 B.n271 B.n132 585
R75 B.n270 B.n269 585
R76 B.n268 B.n133 585
R77 B.n267 B.n266 585
R78 B.n265 B.n134 585
R79 B.n264 B.n263 585
R80 B.n262 B.n135 585
R81 B.n261 B.n260 585
R82 B.n259 B.n136 585
R83 B.n258 B.n257 585
R84 B.n256 B.n137 585
R85 B.n255 B.n254 585
R86 B.n253 B.n138 585
R87 B.n252 B.n251 585
R88 B.n250 B.n139 585
R89 B.n249 B.n248 585
R90 B.n247 B.n140 585
R91 B.n246 B.n245 585
R92 B.n244 B.n141 585
R93 B.n243 B.n242 585
R94 B.n241 B.n142 585
R95 B.n240 B.n239 585
R96 B.n238 B.n143 585
R97 B.n237 B.n236 585
R98 B.n235 B.n144 585
R99 B.n234 B.n233 585
R100 B.n232 B.n145 585
R101 B.n231 B.n230 585
R102 B.n229 B.n146 585
R103 B.n228 B.n227 585
R104 B.n226 B.n147 585
R105 B.n225 B.n224 585
R106 B.n223 B.n148 585
R107 B.n222 B.n221 585
R108 B.n220 B.n149 585
R109 B.n219 B.n218 585
R110 B.n217 B.n150 585
R111 B.n216 B.n215 585
R112 B.n214 B.n151 585
R113 B.n213 B.n212 585
R114 B.n211 B.n152 585
R115 B.n210 B.n209 585
R116 B.n208 B.n153 585
R117 B.n207 B.n206 585
R118 B.n205 B.n154 585
R119 B.n204 B.n203 585
R120 B.n202 B.n155 585
R121 B.n201 B.n200 585
R122 B.n199 B.n156 585
R123 B.n198 B.n197 585
R124 B.n196 B.n157 585
R125 B.n195 B.n194 585
R126 B.n193 B.n158 585
R127 B.n192 B.n191 585
R128 B.n382 B.n381 585
R129 B.n383 B.n94 585
R130 B.n385 B.n384 585
R131 B.n386 B.n93 585
R132 B.n388 B.n387 585
R133 B.n389 B.n92 585
R134 B.n391 B.n390 585
R135 B.n392 B.n91 585
R136 B.n394 B.n393 585
R137 B.n395 B.n90 585
R138 B.n397 B.n396 585
R139 B.n398 B.n89 585
R140 B.n400 B.n399 585
R141 B.n401 B.n88 585
R142 B.n403 B.n402 585
R143 B.n404 B.n87 585
R144 B.n406 B.n405 585
R145 B.n407 B.n86 585
R146 B.n409 B.n408 585
R147 B.n410 B.n85 585
R148 B.n412 B.n411 585
R149 B.n413 B.n84 585
R150 B.n415 B.n414 585
R151 B.n416 B.n83 585
R152 B.n418 B.n417 585
R153 B.n419 B.n82 585
R154 B.n421 B.n420 585
R155 B.n422 B.n81 585
R156 B.n424 B.n423 585
R157 B.n425 B.n80 585
R158 B.n427 B.n426 585
R159 B.n428 B.n79 585
R160 B.n430 B.n429 585
R161 B.n431 B.n78 585
R162 B.n433 B.n432 585
R163 B.n434 B.n77 585
R164 B.n622 B.n621 585
R165 B.n620 B.n11 585
R166 B.n619 B.n618 585
R167 B.n617 B.n12 585
R168 B.n616 B.n615 585
R169 B.n614 B.n13 585
R170 B.n613 B.n612 585
R171 B.n611 B.n14 585
R172 B.n610 B.n609 585
R173 B.n608 B.n15 585
R174 B.n607 B.n606 585
R175 B.n605 B.n16 585
R176 B.n604 B.n603 585
R177 B.n602 B.n17 585
R178 B.n601 B.n600 585
R179 B.n599 B.n18 585
R180 B.n598 B.n597 585
R181 B.n596 B.n19 585
R182 B.n595 B.n594 585
R183 B.n593 B.n20 585
R184 B.n592 B.n591 585
R185 B.n590 B.n21 585
R186 B.n589 B.n588 585
R187 B.n587 B.n22 585
R188 B.n586 B.n585 585
R189 B.n584 B.n23 585
R190 B.n583 B.n582 585
R191 B.n581 B.n24 585
R192 B.n580 B.n579 585
R193 B.n578 B.n25 585
R194 B.n577 B.n576 585
R195 B.n575 B.n26 585
R196 B.n574 B.n573 585
R197 B.n572 B.n27 585
R198 B.n571 B.n570 585
R199 B.n569 B.n28 585
R200 B.n568 B.n567 585
R201 B.n566 B.n29 585
R202 B.n565 B.n564 585
R203 B.n563 B.n30 585
R204 B.n562 B.n561 585
R205 B.n560 B.n31 585
R206 B.n559 B.n558 585
R207 B.n557 B.n32 585
R208 B.n556 B.n555 585
R209 B.n554 B.n33 585
R210 B.n553 B.n552 585
R211 B.n551 B.n34 585
R212 B.n550 B.n549 585
R213 B.n548 B.n35 585
R214 B.n547 B.n546 585
R215 B.n545 B.n36 585
R216 B.n544 B.n543 585
R217 B.n542 B.n37 585
R218 B.n541 B.n540 585
R219 B.n539 B.n38 585
R220 B.n538 B.n537 585
R221 B.n535 B.n39 585
R222 B.n534 B.n533 585
R223 B.n532 B.n42 585
R224 B.n531 B.n530 585
R225 B.n529 B.n43 585
R226 B.n528 B.n527 585
R227 B.n526 B.n44 585
R228 B.n525 B.n524 585
R229 B.n523 B.n45 585
R230 B.n522 B.n521 585
R231 B.n520 B.n519 585
R232 B.n518 B.n49 585
R233 B.n517 B.n516 585
R234 B.n515 B.n50 585
R235 B.n514 B.n513 585
R236 B.n512 B.n51 585
R237 B.n511 B.n510 585
R238 B.n509 B.n52 585
R239 B.n508 B.n507 585
R240 B.n506 B.n53 585
R241 B.n505 B.n504 585
R242 B.n503 B.n54 585
R243 B.n502 B.n501 585
R244 B.n500 B.n55 585
R245 B.n499 B.n498 585
R246 B.n497 B.n56 585
R247 B.n496 B.n495 585
R248 B.n494 B.n57 585
R249 B.n493 B.n492 585
R250 B.n491 B.n58 585
R251 B.n490 B.n489 585
R252 B.n488 B.n59 585
R253 B.n487 B.n486 585
R254 B.n485 B.n60 585
R255 B.n484 B.n483 585
R256 B.n482 B.n61 585
R257 B.n481 B.n480 585
R258 B.n479 B.n62 585
R259 B.n478 B.n477 585
R260 B.n476 B.n63 585
R261 B.n475 B.n474 585
R262 B.n473 B.n64 585
R263 B.n472 B.n471 585
R264 B.n470 B.n65 585
R265 B.n469 B.n468 585
R266 B.n467 B.n66 585
R267 B.n466 B.n465 585
R268 B.n464 B.n67 585
R269 B.n463 B.n462 585
R270 B.n461 B.n68 585
R271 B.n460 B.n459 585
R272 B.n458 B.n69 585
R273 B.n457 B.n456 585
R274 B.n455 B.n70 585
R275 B.n454 B.n453 585
R276 B.n452 B.n71 585
R277 B.n451 B.n450 585
R278 B.n449 B.n72 585
R279 B.n448 B.n447 585
R280 B.n446 B.n73 585
R281 B.n445 B.n444 585
R282 B.n443 B.n74 585
R283 B.n442 B.n441 585
R284 B.n440 B.n75 585
R285 B.n439 B.n438 585
R286 B.n437 B.n76 585
R287 B.n436 B.n435 585
R288 B.n623 B.n10 585
R289 B.n625 B.n624 585
R290 B.n626 B.n9 585
R291 B.n628 B.n627 585
R292 B.n629 B.n8 585
R293 B.n631 B.n630 585
R294 B.n632 B.n7 585
R295 B.n634 B.n633 585
R296 B.n635 B.n6 585
R297 B.n637 B.n636 585
R298 B.n638 B.n5 585
R299 B.n640 B.n639 585
R300 B.n641 B.n4 585
R301 B.n643 B.n642 585
R302 B.n644 B.n3 585
R303 B.n646 B.n645 585
R304 B.n647 B.n0 585
R305 B.n2 B.n1 585
R306 B.n168 B.n167 585
R307 B.n169 B.n166 585
R308 B.n171 B.n170 585
R309 B.n172 B.n165 585
R310 B.n174 B.n173 585
R311 B.n175 B.n164 585
R312 B.n177 B.n176 585
R313 B.n178 B.n163 585
R314 B.n180 B.n179 585
R315 B.n181 B.n162 585
R316 B.n183 B.n182 585
R317 B.n184 B.n161 585
R318 B.n186 B.n185 585
R319 B.n187 B.n160 585
R320 B.n189 B.n188 585
R321 B.n190 B.n159 585
R322 B.n192 B.n159 545.355
R323 B.n382 B.n95 545.355
R324 B.n436 B.n77 545.355
R325 B.n623 B.n622 545.355
R326 B.n649 B.n648 256.663
R327 B.n648 B.n647 235.042
R328 B.n648 B.n2 235.042
R329 B.n193 B.n192 163.367
R330 B.n194 B.n193 163.367
R331 B.n194 B.n157 163.367
R332 B.n198 B.n157 163.367
R333 B.n199 B.n198 163.367
R334 B.n200 B.n199 163.367
R335 B.n200 B.n155 163.367
R336 B.n204 B.n155 163.367
R337 B.n205 B.n204 163.367
R338 B.n206 B.n205 163.367
R339 B.n206 B.n153 163.367
R340 B.n210 B.n153 163.367
R341 B.n211 B.n210 163.367
R342 B.n212 B.n211 163.367
R343 B.n212 B.n151 163.367
R344 B.n216 B.n151 163.367
R345 B.n217 B.n216 163.367
R346 B.n218 B.n217 163.367
R347 B.n218 B.n149 163.367
R348 B.n222 B.n149 163.367
R349 B.n223 B.n222 163.367
R350 B.n224 B.n223 163.367
R351 B.n224 B.n147 163.367
R352 B.n228 B.n147 163.367
R353 B.n229 B.n228 163.367
R354 B.n230 B.n229 163.367
R355 B.n230 B.n145 163.367
R356 B.n234 B.n145 163.367
R357 B.n235 B.n234 163.367
R358 B.n236 B.n235 163.367
R359 B.n236 B.n143 163.367
R360 B.n240 B.n143 163.367
R361 B.n241 B.n240 163.367
R362 B.n242 B.n241 163.367
R363 B.n242 B.n141 163.367
R364 B.n246 B.n141 163.367
R365 B.n247 B.n246 163.367
R366 B.n248 B.n247 163.367
R367 B.n248 B.n139 163.367
R368 B.n252 B.n139 163.367
R369 B.n253 B.n252 163.367
R370 B.n254 B.n253 163.367
R371 B.n254 B.n137 163.367
R372 B.n258 B.n137 163.367
R373 B.n259 B.n258 163.367
R374 B.n260 B.n259 163.367
R375 B.n260 B.n135 163.367
R376 B.n264 B.n135 163.367
R377 B.n265 B.n264 163.367
R378 B.n266 B.n265 163.367
R379 B.n266 B.n133 163.367
R380 B.n270 B.n133 163.367
R381 B.n271 B.n270 163.367
R382 B.n272 B.n271 163.367
R383 B.n272 B.n131 163.367
R384 B.n279 B.n131 163.367
R385 B.n280 B.n279 163.367
R386 B.n281 B.n280 163.367
R387 B.n281 B.n129 163.367
R388 B.n285 B.n129 163.367
R389 B.n286 B.n285 163.367
R390 B.n287 B.n286 163.367
R391 B.n287 B.n127 163.367
R392 B.n291 B.n127 163.367
R393 B.n292 B.n291 163.367
R394 B.n293 B.n292 163.367
R395 B.n293 B.n123 163.367
R396 B.n298 B.n123 163.367
R397 B.n299 B.n298 163.367
R398 B.n300 B.n299 163.367
R399 B.n300 B.n121 163.367
R400 B.n304 B.n121 163.367
R401 B.n305 B.n304 163.367
R402 B.n306 B.n305 163.367
R403 B.n306 B.n119 163.367
R404 B.n310 B.n119 163.367
R405 B.n311 B.n310 163.367
R406 B.n312 B.n311 163.367
R407 B.n312 B.n117 163.367
R408 B.n316 B.n117 163.367
R409 B.n317 B.n316 163.367
R410 B.n318 B.n317 163.367
R411 B.n318 B.n115 163.367
R412 B.n322 B.n115 163.367
R413 B.n323 B.n322 163.367
R414 B.n324 B.n323 163.367
R415 B.n324 B.n113 163.367
R416 B.n328 B.n113 163.367
R417 B.n329 B.n328 163.367
R418 B.n330 B.n329 163.367
R419 B.n330 B.n111 163.367
R420 B.n334 B.n111 163.367
R421 B.n335 B.n334 163.367
R422 B.n336 B.n335 163.367
R423 B.n336 B.n109 163.367
R424 B.n340 B.n109 163.367
R425 B.n341 B.n340 163.367
R426 B.n342 B.n341 163.367
R427 B.n342 B.n107 163.367
R428 B.n346 B.n107 163.367
R429 B.n347 B.n346 163.367
R430 B.n348 B.n347 163.367
R431 B.n348 B.n105 163.367
R432 B.n352 B.n105 163.367
R433 B.n353 B.n352 163.367
R434 B.n354 B.n353 163.367
R435 B.n354 B.n103 163.367
R436 B.n358 B.n103 163.367
R437 B.n359 B.n358 163.367
R438 B.n360 B.n359 163.367
R439 B.n360 B.n101 163.367
R440 B.n364 B.n101 163.367
R441 B.n365 B.n364 163.367
R442 B.n366 B.n365 163.367
R443 B.n366 B.n99 163.367
R444 B.n370 B.n99 163.367
R445 B.n371 B.n370 163.367
R446 B.n372 B.n371 163.367
R447 B.n372 B.n97 163.367
R448 B.n376 B.n97 163.367
R449 B.n377 B.n376 163.367
R450 B.n378 B.n377 163.367
R451 B.n378 B.n95 163.367
R452 B.n432 B.n77 163.367
R453 B.n432 B.n431 163.367
R454 B.n431 B.n430 163.367
R455 B.n430 B.n79 163.367
R456 B.n426 B.n79 163.367
R457 B.n426 B.n425 163.367
R458 B.n425 B.n424 163.367
R459 B.n424 B.n81 163.367
R460 B.n420 B.n81 163.367
R461 B.n420 B.n419 163.367
R462 B.n419 B.n418 163.367
R463 B.n418 B.n83 163.367
R464 B.n414 B.n83 163.367
R465 B.n414 B.n413 163.367
R466 B.n413 B.n412 163.367
R467 B.n412 B.n85 163.367
R468 B.n408 B.n85 163.367
R469 B.n408 B.n407 163.367
R470 B.n407 B.n406 163.367
R471 B.n406 B.n87 163.367
R472 B.n402 B.n87 163.367
R473 B.n402 B.n401 163.367
R474 B.n401 B.n400 163.367
R475 B.n400 B.n89 163.367
R476 B.n396 B.n89 163.367
R477 B.n396 B.n395 163.367
R478 B.n395 B.n394 163.367
R479 B.n394 B.n91 163.367
R480 B.n390 B.n91 163.367
R481 B.n390 B.n389 163.367
R482 B.n389 B.n388 163.367
R483 B.n388 B.n93 163.367
R484 B.n384 B.n93 163.367
R485 B.n384 B.n383 163.367
R486 B.n383 B.n382 163.367
R487 B.n622 B.n11 163.367
R488 B.n618 B.n11 163.367
R489 B.n618 B.n617 163.367
R490 B.n617 B.n616 163.367
R491 B.n616 B.n13 163.367
R492 B.n612 B.n13 163.367
R493 B.n612 B.n611 163.367
R494 B.n611 B.n610 163.367
R495 B.n610 B.n15 163.367
R496 B.n606 B.n15 163.367
R497 B.n606 B.n605 163.367
R498 B.n605 B.n604 163.367
R499 B.n604 B.n17 163.367
R500 B.n600 B.n17 163.367
R501 B.n600 B.n599 163.367
R502 B.n599 B.n598 163.367
R503 B.n598 B.n19 163.367
R504 B.n594 B.n19 163.367
R505 B.n594 B.n593 163.367
R506 B.n593 B.n592 163.367
R507 B.n592 B.n21 163.367
R508 B.n588 B.n21 163.367
R509 B.n588 B.n587 163.367
R510 B.n587 B.n586 163.367
R511 B.n586 B.n23 163.367
R512 B.n582 B.n23 163.367
R513 B.n582 B.n581 163.367
R514 B.n581 B.n580 163.367
R515 B.n580 B.n25 163.367
R516 B.n576 B.n25 163.367
R517 B.n576 B.n575 163.367
R518 B.n575 B.n574 163.367
R519 B.n574 B.n27 163.367
R520 B.n570 B.n27 163.367
R521 B.n570 B.n569 163.367
R522 B.n569 B.n568 163.367
R523 B.n568 B.n29 163.367
R524 B.n564 B.n29 163.367
R525 B.n564 B.n563 163.367
R526 B.n563 B.n562 163.367
R527 B.n562 B.n31 163.367
R528 B.n558 B.n31 163.367
R529 B.n558 B.n557 163.367
R530 B.n557 B.n556 163.367
R531 B.n556 B.n33 163.367
R532 B.n552 B.n33 163.367
R533 B.n552 B.n551 163.367
R534 B.n551 B.n550 163.367
R535 B.n550 B.n35 163.367
R536 B.n546 B.n35 163.367
R537 B.n546 B.n545 163.367
R538 B.n545 B.n544 163.367
R539 B.n544 B.n37 163.367
R540 B.n540 B.n37 163.367
R541 B.n540 B.n539 163.367
R542 B.n539 B.n538 163.367
R543 B.n538 B.n39 163.367
R544 B.n533 B.n39 163.367
R545 B.n533 B.n532 163.367
R546 B.n532 B.n531 163.367
R547 B.n531 B.n43 163.367
R548 B.n527 B.n43 163.367
R549 B.n527 B.n526 163.367
R550 B.n526 B.n525 163.367
R551 B.n525 B.n45 163.367
R552 B.n521 B.n45 163.367
R553 B.n521 B.n520 163.367
R554 B.n520 B.n49 163.367
R555 B.n516 B.n49 163.367
R556 B.n516 B.n515 163.367
R557 B.n515 B.n514 163.367
R558 B.n514 B.n51 163.367
R559 B.n510 B.n51 163.367
R560 B.n510 B.n509 163.367
R561 B.n509 B.n508 163.367
R562 B.n508 B.n53 163.367
R563 B.n504 B.n53 163.367
R564 B.n504 B.n503 163.367
R565 B.n503 B.n502 163.367
R566 B.n502 B.n55 163.367
R567 B.n498 B.n55 163.367
R568 B.n498 B.n497 163.367
R569 B.n497 B.n496 163.367
R570 B.n496 B.n57 163.367
R571 B.n492 B.n57 163.367
R572 B.n492 B.n491 163.367
R573 B.n491 B.n490 163.367
R574 B.n490 B.n59 163.367
R575 B.n486 B.n59 163.367
R576 B.n486 B.n485 163.367
R577 B.n485 B.n484 163.367
R578 B.n484 B.n61 163.367
R579 B.n480 B.n61 163.367
R580 B.n480 B.n479 163.367
R581 B.n479 B.n478 163.367
R582 B.n478 B.n63 163.367
R583 B.n474 B.n63 163.367
R584 B.n474 B.n473 163.367
R585 B.n473 B.n472 163.367
R586 B.n472 B.n65 163.367
R587 B.n468 B.n65 163.367
R588 B.n468 B.n467 163.367
R589 B.n467 B.n466 163.367
R590 B.n466 B.n67 163.367
R591 B.n462 B.n67 163.367
R592 B.n462 B.n461 163.367
R593 B.n461 B.n460 163.367
R594 B.n460 B.n69 163.367
R595 B.n456 B.n69 163.367
R596 B.n456 B.n455 163.367
R597 B.n455 B.n454 163.367
R598 B.n454 B.n71 163.367
R599 B.n450 B.n71 163.367
R600 B.n450 B.n449 163.367
R601 B.n449 B.n448 163.367
R602 B.n448 B.n73 163.367
R603 B.n444 B.n73 163.367
R604 B.n444 B.n443 163.367
R605 B.n443 B.n442 163.367
R606 B.n442 B.n75 163.367
R607 B.n438 B.n75 163.367
R608 B.n438 B.n437 163.367
R609 B.n437 B.n436 163.367
R610 B.n624 B.n623 163.367
R611 B.n624 B.n9 163.367
R612 B.n628 B.n9 163.367
R613 B.n629 B.n628 163.367
R614 B.n630 B.n629 163.367
R615 B.n630 B.n7 163.367
R616 B.n634 B.n7 163.367
R617 B.n635 B.n634 163.367
R618 B.n636 B.n635 163.367
R619 B.n636 B.n5 163.367
R620 B.n640 B.n5 163.367
R621 B.n641 B.n640 163.367
R622 B.n642 B.n641 163.367
R623 B.n642 B.n3 163.367
R624 B.n646 B.n3 163.367
R625 B.n647 B.n646 163.367
R626 B.n168 B.n2 163.367
R627 B.n169 B.n168 163.367
R628 B.n170 B.n169 163.367
R629 B.n170 B.n165 163.367
R630 B.n174 B.n165 163.367
R631 B.n175 B.n174 163.367
R632 B.n176 B.n175 163.367
R633 B.n176 B.n163 163.367
R634 B.n180 B.n163 163.367
R635 B.n181 B.n180 163.367
R636 B.n182 B.n181 163.367
R637 B.n182 B.n161 163.367
R638 B.n186 B.n161 163.367
R639 B.n187 B.n186 163.367
R640 B.n188 B.n187 163.367
R641 B.n188 B.n159 163.367
R642 B.n124 B.t1 133.619
R643 B.n46 B.t8 133.619
R644 B.n275 B.t4 133.597
R645 B.n40 B.t11 133.597
R646 B.n125 B.t2 112.48
R647 B.n47 B.t7 112.48
R648 B.n276 B.t5 112.457
R649 B.n41 B.t10 112.457
R650 B.n277 B.n276 59.5399
R651 B.n295 B.n125 59.5399
R652 B.n48 B.n47 59.5399
R653 B.n536 B.n41 59.5399
R654 B.n381 B.n380 35.4346
R655 B.n621 B.n10 35.4346
R656 B.n435 B.n434 35.4346
R657 B.n191 B.n190 35.4346
R658 B.n276 B.n275 21.1399
R659 B.n125 B.n124 21.1399
R660 B.n47 B.n46 21.1399
R661 B.n41 B.n40 21.1399
R662 B B.n649 18.0485
R663 B.n625 B.n10 10.6151
R664 B.n626 B.n625 10.6151
R665 B.n627 B.n626 10.6151
R666 B.n627 B.n8 10.6151
R667 B.n631 B.n8 10.6151
R668 B.n632 B.n631 10.6151
R669 B.n633 B.n632 10.6151
R670 B.n633 B.n6 10.6151
R671 B.n637 B.n6 10.6151
R672 B.n638 B.n637 10.6151
R673 B.n639 B.n638 10.6151
R674 B.n639 B.n4 10.6151
R675 B.n643 B.n4 10.6151
R676 B.n644 B.n643 10.6151
R677 B.n645 B.n644 10.6151
R678 B.n645 B.n0 10.6151
R679 B.n621 B.n620 10.6151
R680 B.n620 B.n619 10.6151
R681 B.n619 B.n12 10.6151
R682 B.n615 B.n12 10.6151
R683 B.n615 B.n614 10.6151
R684 B.n614 B.n613 10.6151
R685 B.n613 B.n14 10.6151
R686 B.n609 B.n14 10.6151
R687 B.n609 B.n608 10.6151
R688 B.n608 B.n607 10.6151
R689 B.n607 B.n16 10.6151
R690 B.n603 B.n16 10.6151
R691 B.n603 B.n602 10.6151
R692 B.n602 B.n601 10.6151
R693 B.n601 B.n18 10.6151
R694 B.n597 B.n18 10.6151
R695 B.n597 B.n596 10.6151
R696 B.n596 B.n595 10.6151
R697 B.n595 B.n20 10.6151
R698 B.n591 B.n20 10.6151
R699 B.n591 B.n590 10.6151
R700 B.n590 B.n589 10.6151
R701 B.n589 B.n22 10.6151
R702 B.n585 B.n22 10.6151
R703 B.n585 B.n584 10.6151
R704 B.n584 B.n583 10.6151
R705 B.n583 B.n24 10.6151
R706 B.n579 B.n24 10.6151
R707 B.n579 B.n578 10.6151
R708 B.n578 B.n577 10.6151
R709 B.n577 B.n26 10.6151
R710 B.n573 B.n26 10.6151
R711 B.n573 B.n572 10.6151
R712 B.n572 B.n571 10.6151
R713 B.n571 B.n28 10.6151
R714 B.n567 B.n28 10.6151
R715 B.n567 B.n566 10.6151
R716 B.n566 B.n565 10.6151
R717 B.n565 B.n30 10.6151
R718 B.n561 B.n30 10.6151
R719 B.n561 B.n560 10.6151
R720 B.n560 B.n559 10.6151
R721 B.n559 B.n32 10.6151
R722 B.n555 B.n32 10.6151
R723 B.n555 B.n554 10.6151
R724 B.n554 B.n553 10.6151
R725 B.n553 B.n34 10.6151
R726 B.n549 B.n34 10.6151
R727 B.n549 B.n548 10.6151
R728 B.n548 B.n547 10.6151
R729 B.n547 B.n36 10.6151
R730 B.n543 B.n36 10.6151
R731 B.n543 B.n542 10.6151
R732 B.n542 B.n541 10.6151
R733 B.n541 B.n38 10.6151
R734 B.n537 B.n38 10.6151
R735 B.n535 B.n534 10.6151
R736 B.n534 B.n42 10.6151
R737 B.n530 B.n42 10.6151
R738 B.n530 B.n529 10.6151
R739 B.n529 B.n528 10.6151
R740 B.n528 B.n44 10.6151
R741 B.n524 B.n44 10.6151
R742 B.n524 B.n523 10.6151
R743 B.n523 B.n522 10.6151
R744 B.n519 B.n518 10.6151
R745 B.n518 B.n517 10.6151
R746 B.n517 B.n50 10.6151
R747 B.n513 B.n50 10.6151
R748 B.n513 B.n512 10.6151
R749 B.n512 B.n511 10.6151
R750 B.n511 B.n52 10.6151
R751 B.n507 B.n52 10.6151
R752 B.n507 B.n506 10.6151
R753 B.n506 B.n505 10.6151
R754 B.n505 B.n54 10.6151
R755 B.n501 B.n54 10.6151
R756 B.n501 B.n500 10.6151
R757 B.n500 B.n499 10.6151
R758 B.n499 B.n56 10.6151
R759 B.n495 B.n56 10.6151
R760 B.n495 B.n494 10.6151
R761 B.n494 B.n493 10.6151
R762 B.n493 B.n58 10.6151
R763 B.n489 B.n58 10.6151
R764 B.n489 B.n488 10.6151
R765 B.n488 B.n487 10.6151
R766 B.n487 B.n60 10.6151
R767 B.n483 B.n60 10.6151
R768 B.n483 B.n482 10.6151
R769 B.n482 B.n481 10.6151
R770 B.n481 B.n62 10.6151
R771 B.n477 B.n62 10.6151
R772 B.n477 B.n476 10.6151
R773 B.n476 B.n475 10.6151
R774 B.n475 B.n64 10.6151
R775 B.n471 B.n64 10.6151
R776 B.n471 B.n470 10.6151
R777 B.n470 B.n469 10.6151
R778 B.n469 B.n66 10.6151
R779 B.n465 B.n66 10.6151
R780 B.n465 B.n464 10.6151
R781 B.n464 B.n463 10.6151
R782 B.n463 B.n68 10.6151
R783 B.n459 B.n68 10.6151
R784 B.n459 B.n458 10.6151
R785 B.n458 B.n457 10.6151
R786 B.n457 B.n70 10.6151
R787 B.n453 B.n70 10.6151
R788 B.n453 B.n452 10.6151
R789 B.n452 B.n451 10.6151
R790 B.n451 B.n72 10.6151
R791 B.n447 B.n72 10.6151
R792 B.n447 B.n446 10.6151
R793 B.n446 B.n445 10.6151
R794 B.n445 B.n74 10.6151
R795 B.n441 B.n74 10.6151
R796 B.n441 B.n440 10.6151
R797 B.n440 B.n439 10.6151
R798 B.n439 B.n76 10.6151
R799 B.n435 B.n76 10.6151
R800 B.n434 B.n433 10.6151
R801 B.n433 B.n78 10.6151
R802 B.n429 B.n78 10.6151
R803 B.n429 B.n428 10.6151
R804 B.n428 B.n427 10.6151
R805 B.n427 B.n80 10.6151
R806 B.n423 B.n80 10.6151
R807 B.n423 B.n422 10.6151
R808 B.n422 B.n421 10.6151
R809 B.n421 B.n82 10.6151
R810 B.n417 B.n82 10.6151
R811 B.n417 B.n416 10.6151
R812 B.n416 B.n415 10.6151
R813 B.n415 B.n84 10.6151
R814 B.n411 B.n84 10.6151
R815 B.n411 B.n410 10.6151
R816 B.n410 B.n409 10.6151
R817 B.n409 B.n86 10.6151
R818 B.n405 B.n86 10.6151
R819 B.n405 B.n404 10.6151
R820 B.n404 B.n403 10.6151
R821 B.n403 B.n88 10.6151
R822 B.n399 B.n88 10.6151
R823 B.n399 B.n398 10.6151
R824 B.n398 B.n397 10.6151
R825 B.n397 B.n90 10.6151
R826 B.n393 B.n90 10.6151
R827 B.n393 B.n392 10.6151
R828 B.n392 B.n391 10.6151
R829 B.n391 B.n92 10.6151
R830 B.n387 B.n92 10.6151
R831 B.n387 B.n386 10.6151
R832 B.n386 B.n385 10.6151
R833 B.n385 B.n94 10.6151
R834 B.n381 B.n94 10.6151
R835 B.n167 B.n1 10.6151
R836 B.n167 B.n166 10.6151
R837 B.n171 B.n166 10.6151
R838 B.n172 B.n171 10.6151
R839 B.n173 B.n172 10.6151
R840 B.n173 B.n164 10.6151
R841 B.n177 B.n164 10.6151
R842 B.n178 B.n177 10.6151
R843 B.n179 B.n178 10.6151
R844 B.n179 B.n162 10.6151
R845 B.n183 B.n162 10.6151
R846 B.n184 B.n183 10.6151
R847 B.n185 B.n184 10.6151
R848 B.n185 B.n160 10.6151
R849 B.n189 B.n160 10.6151
R850 B.n190 B.n189 10.6151
R851 B.n191 B.n158 10.6151
R852 B.n195 B.n158 10.6151
R853 B.n196 B.n195 10.6151
R854 B.n197 B.n196 10.6151
R855 B.n197 B.n156 10.6151
R856 B.n201 B.n156 10.6151
R857 B.n202 B.n201 10.6151
R858 B.n203 B.n202 10.6151
R859 B.n203 B.n154 10.6151
R860 B.n207 B.n154 10.6151
R861 B.n208 B.n207 10.6151
R862 B.n209 B.n208 10.6151
R863 B.n209 B.n152 10.6151
R864 B.n213 B.n152 10.6151
R865 B.n214 B.n213 10.6151
R866 B.n215 B.n214 10.6151
R867 B.n215 B.n150 10.6151
R868 B.n219 B.n150 10.6151
R869 B.n220 B.n219 10.6151
R870 B.n221 B.n220 10.6151
R871 B.n221 B.n148 10.6151
R872 B.n225 B.n148 10.6151
R873 B.n226 B.n225 10.6151
R874 B.n227 B.n226 10.6151
R875 B.n227 B.n146 10.6151
R876 B.n231 B.n146 10.6151
R877 B.n232 B.n231 10.6151
R878 B.n233 B.n232 10.6151
R879 B.n233 B.n144 10.6151
R880 B.n237 B.n144 10.6151
R881 B.n238 B.n237 10.6151
R882 B.n239 B.n238 10.6151
R883 B.n239 B.n142 10.6151
R884 B.n243 B.n142 10.6151
R885 B.n244 B.n243 10.6151
R886 B.n245 B.n244 10.6151
R887 B.n245 B.n140 10.6151
R888 B.n249 B.n140 10.6151
R889 B.n250 B.n249 10.6151
R890 B.n251 B.n250 10.6151
R891 B.n251 B.n138 10.6151
R892 B.n255 B.n138 10.6151
R893 B.n256 B.n255 10.6151
R894 B.n257 B.n256 10.6151
R895 B.n257 B.n136 10.6151
R896 B.n261 B.n136 10.6151
R897 B.n262 B.n261 10.6151
R898 B.n263 B.n262 10.6151
R899 B.n263 B.n134 10.6151
R900 B.n267 B.n134 10.6151
R901 B.n268 B.n267 10.6151
R902 B.n269 B.n268 10.6151
R903 B.n269 B.n132 10.6151
R904 B.n273 B.n132 10.6151
R905 B.n274 B.n273 10.6151
R906 B.n278 B.n274 10.6151
R907 B.n282 B.n130 10.6151
R908 B.n283 B.n282 10.6151
R909 B.n284 B.n283 10.6151
R910 B.n284 B.n128 10.6151
R911 B.n288 B.n128 10.6151
R912 B.n289 B.n288 10.6151
R913 B.n290 B.n289 10.6151
R914 B.n290 B.n126 10.6151
R915 B.n294 B.n126 10.6151
R916 B.n297 B.n296 10.6151
R917 B.n297 B.n122 10.6151
R918 B.n301 B.n122 10.6151
R919 B.n302 B.n301 10.6151
R920 B.n303 B.n302 10.6151
R921 B.n303 B.n120 10.6151
R922 B.n307 B.n120 10.6151
R923 B.n308 B.n307 10.6151
R924 B.n309 B.n308 10.6151
R925 B.n309 B.n118 10.6151
R926 B.n313 B.n118 10.6151
R927 B.n314 B.n313 10.6151
R928 B.n315 B.n314 10.6151
R929 B.n315 B.n116 10.6151
R930 B.n319 B.n116 10.6151
R931 B.n320 B.n319 10.6151
R932 B.n321 B.n320 10.6151
R933 B.n321 B.n114 10.6151
R934 B.n325 B.n114 10.6151
R935 B.n326 B.n325 10.6151
R936 B.n327 B.n326 10.6151
R937 B.n327 B.n112 10.6151
R938 B.n331 B.n112 10.6151
R939 B.n332 B.n331 10.6151
R940 B.n333 B.n332 10.6151
R941 B.n333 B.n110 10.6151
R942 B.n337 B.n110 10.6151
R943 B.n338 B.n337 10.6151
R944 B.n339 B.n338 10.6151
R945 B.n339 B.n108 10.6151
R946 B.n343 B.n108 10.6151
R947 B.n344 B.n343 10.6151
R948 B.n345 B.n344 10.6151
R949 B.n345 B.n106 10.6151
R950 B.n349 B.n106 10.6151
R951 B.n350 B.n349 10.6151
R952 B.n351 B.n350 10.6151
R953 B.n351 B.n104 10.6151
R954 B.n355 B.n104 10.6151
R955 B.n356 B.n355 10.6151
R956 B.n357 B.n356 10.6151
R957 B.n357 B.n102 10.6151
R958 B.n361 B.n102 10.6151
R959 B.n362 B.n361 10.6151
R960 B.n363 B.n362 10.6151
R961 B.n363 B.n100 10.6151
R962 B.n367 B.n100 10.6151
R963 B.n368 B.n367 10.6151
R964 B.n369 B.n368 10.6151
R965 B.n369 B.n98 10.6151
R966 B.n373 B.n98 10.6151
R967 B.n374 B.n373 10.6151
R968 B.n375 B.n374 10.6151
R969 B.n375 B.n96 10.6151
R970 B.n379 B.n96 10.6151
R971 B.n380 B.n379 10.6151
R972 B.n537 B.n536 9.36635
R973 B.n519 B.n48 9.36635
R974 B.n278 B.n277 9.36635
R975 B.n296 B.n295 9.36635
R976 B.n649 B.n0 8.11757
R977 B.n649 B.n1 8.11757
R978 B.n536 B.n535 1.24928
R979 B.n522 B.n48 1.24928
R980 B.n277 B.n130 1.24928
R981 B.n295 B.n294 1.24928
R982 VP.n1 VP.t0 621.912
R983 VP.n1 VP.t3 621.861
R984 VP.n3 VP.t1 600.914
R985 VP.n5 VP.t2 600.914
R986 VP.n6 VP.n5 161.3
R987 VP.n4 VP.n0 161.3
R988 VP.n3 VP.n2 161.3
R989 VP.n2 VP.n1 89.3287
R990 VP.n4 VP.n3 24.1005
R991 VP.n5 VP.n4 24.1005
R992 VP.n2 VP.n0 0.189894
R993 VP.n6 VP.n0 0.189894
R994 VP VP.n6 0.0516364
R995 VDD1 VDD1.n1 114.294
R996 VDD1 VDD1.n0 72.3632
R997 VDD1.n0 VDD1.t1 1.87723
R998 VDD1.n0 VDD1.t3 1.87723
R999 VDD1.n1 VDD1.t0 1.87723
R1000 VDD1.n1 VDD1.t2 1.87723
R1001 VTAIL.n5 VTAIL.t7 57.5031
R1002 VTAIL.n4 VTAIL.t3 57.5031
R1003 VTAIL.n3 VTAIL.t2 57.5031
R1004 VTAIL.n7 VTAIL.t1 57.503
R1005 VTAIL.n0 VTAIL.t0 57.503
R1006 VTAIL.n1 VTAIL.t5 57.503
R1007 VTAIL.n2 VTAIL.t6 57.503
R1008 VTAIL.n6 VTAIL.t4 57.503
R1009 VTAIL.n7 VTAIL.n6 28.2376
R1010 VTAIL.n3 VTAIL.n2 28.2376
R1011 VTAIL.n4 VTAIL.n3 0.940155
R1012 VTAIL.n6 VTAIL.n5 0.940155
R1013 VTAIL.n2 VTAIL.n1 0.940155
R1014 VTAIL VTAIL.n0 0.528517
R1015 VTAIL.n5 VTAIL.n4 0.470328
R1016 VTAIL.n1 VTAIL.n0 0.470328
R1017 VTAIL VTAIL.n7 0.412138
R1018 VN.n0 VN.t1 621.912
R1019 VN.n1 VN.t0 621.912
R1020 VN.n0 VN.t2 621.861
R1021 VN.n1 VN.t3 621.861
R1022 VN VN.n1 89.7094
R1023 VN VN.n0 44.7132
R1024 VDD2.n2 VDD2.n0 113.769
R1025 VDD2.n2 VDD2.n1 72.305
R1026 VDD2.n1 VDD2.t0 1.87723
R1027 VDD2.n1 VDD2.t3 1.87723
R1028 VDD2.n0 VDD2.t2 1.87723
R1029 VDD2.n0 VDD2.t1 1.87723
R1030 VDD2 VDD2.n2 0.0586897
C0 VDD2 VP 0.277364f
C1 w_n1624_n4432# VP 2.71429f
C2 VP VDD1 4.73546f
C3 VTAIL VN 4.01121f
C4 VDD2 VTAIL 8.89782f
C5 VTAIL w_n1624_n4432# 5.44989f
C6 VTAIL VDD1 8.85595f
C7 B VP 1.15288f
C8 VDD2 VN 4.60585f
C9 w_n1624_n4432# VN 2.51017f
C10 VN VDD1 0.147478f
C11 VTAIL B 5.31423f
C12 VDD2 w_n1624_n4432# 1.23285f
C13 VDD2 VDD1 0.580232f
C14 w_n1624_n4432# VDD1 1.21712f
C15 VTAIL VP 4.02532f
C16 B VN 0.822723f
C17 VDD2 B 1.10246f
C18 B w_n1624_n4432# 8.473001f
C19 B VDD1 1.08008f
C20 VN VP 5.84798f
C21 VDD2 VSUBS 0.813453f
C22 VDD1 VSUBS 5.746703f
C23 VTAIL VSUBS 1.128602f
C24 VN VSUBS 6.22444f
C25 VP VSUBS 1.520454f
C26 B VSUBS 3.121181f
C27 w_n1624_n4432# VSUBS 88.0663f
C28 VDD2.t2 VSUBS 0.383887f
C29 VDD2.t1 VSUBS 0.383887f
C30 VDD2.n0 VSUBS 4.02569f
C31 VDD2.t0 VSUBS 0.383887f
C32 VDD2.t3 VSUBS 0.383887f
C33 VDD2.n1 VSUBS 3.18804f
C34 VDD2.n2 VSUBS 4.65976f
C35 VN.t1 VSUBS 2.10269f
C36 VN.t2 VSUBS 2.10262f
C37 VN.n0 VSUBS 1.5225f
C38 VN.t0 VSUBS 2.10269f
C39 VN.t3 VSUBS 2.10262f
C40 VN.n1 VSUBS 2.87673f
C41 VTAIL.t0 VSUBS 3.14027f
C42 VTAIL.n0 VSUBS 0.68893f
C43 VTAIL.t5 VSUBS 3.14027f
C44 VTAIL.n1 VSUBS 0.718466f
C45 VTAIL.t6 VSUBS 3.14027f
C46 VTAIL.n2 VSUBS 2.126f
C47 VTAIL.t2 VSUBS 3.14029f
C48 VTAIL.n3 VSUBS 2.12598f
C49 VTAIL.t3 VSUBS 3.14029f
C50 VTAIL.n4 VSUBS 0.718444f
C51 VTAIL.t7 VSUBS 3.14029f
C52 VTAIL.n5 VSUBS 0.718444f
C53 VTAIL.t4 VSUBS 3.14027f
C54 VTAIL.n6 VSUBS 2.126f
C55 VTAIL.t1 VSUBS 3.14027f
C56 VTAIL.n7 VSUBS 2.08811f
C57 VDD1.t1 VSUBS 0.383785f
C58 VDD1.t3 VSUBS 0.383785f
C59 VDD1.n0 VSUBS 3.18771f
C60 VDD1.t0 VSUBS 0.383785f
C61 VDD1.t2 VSUBS 0.383785f
C62 VDD1.n1 VSUBS 4.05196f
C63 VP.n0 VSUBS 0.056857f
C64 VP.t3 VSUBS 2.14989f
C65 VP.t0 VSUBS 2.14996f
C66 VP.n1 VSUBS 2.91695f
C67 VP.n2 VSUBS 4.00124f
C68 VP.t1 VSUBS 2.12285f
C69 VP.n3 VSUBS 0.798695f
C70 VP.n4 VSUBS 0.012902f
C71 VP.t2 VSUBS 2.12285f
C72 VP.n5 VSUBS 0.798695f
C73 VP.n6 VSUBS 0.044062f
C74 B.n0 VSUBS 0.006791f
C75 B.n1 VSUBS 0.006791f
C76 B.n2 VSUBS 0.010044f
C77 B.n3 VSUBS 0.007697f
C78 B.n4 VSUBS 0.007697f
C79 B.n5 VSUBS 0.007697f
C80 B.n6 VSUBS 0.007697f
C81 B.n7 VSUBS 0.007697f
C82 B.n8 VSUBS 0.007697f
C83 B.n9 VSUBS 0.007697f
C84 B.n10 VSUBS 0.018494f
C85 B.n11 VSUBS 0.007697f
C86 B.n12 VSUBS 0.007697f
C87 B.n13 VSUBS 0.007697f
C88 B.n14 VSUBS 0.007697f
C89 B.n15 VSUBS 0.007697f
C90 B.n16 VSUBS 0.007697f
C91 B.n17 VSUBS 0.007697f
C92 B.n18 VSUBS 0.007697f
C93 B.n19 VSUBS 0.007697f
C94 B.n20 VSUBS 0.007697f
C95 B.n21 VSUBS 0.007697f
C96 B.n22 VSUBS 0.007697f
C97 B.n23 VSUBS 0.007697f
C98 B.n24 VSUBS 0.007697f
C99 B.n25 VSUBS 0.007697f
C100 B.n26 VSUBS 0.007697f
C101 B.n27 VSUBS 0.007697f
C102 B.n28 VSUBS 0.007697f
C103 B.n29 VSUBS 0.007697f
C104 B.n30 VSUBS 0.007697f
C105 B.n31 VSUBS 0.007697f
C106 B.n32 VSUBS 0.007697f
C107 B.n33 VSUBS 0.007697f
C108 B.n34 VSUBS 0.007697f
C109 B.n35 VSUBS 0.007697f
C110 B.n36 VSUBS 0.007697f
C111 B.n37 VSUBS 0.007697f
C112 B.n38 VSUBS 0.007697f
C113 B.n39 VSUBS 0.007697f
C114 B.t10 VSUBS 0.641179f
C115 B.t11 VSUBS 0.650654f
C116 B.t9 VSUBS 0.58748f
C117 B.n40 VSUBS 0.205646f
C118 B.n41 VSUBS 0.070856f
C119 B.n42 VSUBS 0.007697f
C120 B.n43 VSUBS 0.007697f
C121 B.n44 VSUBS 0.007697f
C122 B.n45 VSUBS 0.007697f
C123 B.t7 VSUBS 0.641157f
C124 B.t8 VSUBS 0.650634f
C125 B.t6 VSUBS 0.58748f
C126 B.n46 VSUBS 0.205666f
C127 B.n47 VSUBS 0.070878f
C128 B.n48 VSUBS 0.017833f
C129 B.n49 VSUBS 0.007697f
C130 B.n50 VSUBS 0.007697f
C131 B.n51 VSUBS 0.007697f
C132 B.n52 VSUBS 0.007697f
C133 B.n53 VSUBS 0.007697f
C134 B.n54 VSUBS 0.007697f
C135 B.n55 VSUBS 0.007697f
C136 B.n56 VSUBS 0.007697f
C137 B.n57 VSUBS 0.007697f
C138 B.n58 VSUBS 0.007697f
C139 B.n59 VSUBS 0.007697f
C140 B.n60 VSUBS 0.007697f
C141 B.n61 VSUBS 0.007697f
C142 B.n62 VSUBS 0.007697f
C143 B.n63 VSUBS 0.007697f
C144 B.n64 VSUBS 0.007697f
C145 B.n65 VSUBS 0.007697f
C146 B.n66 VSUBS 0.007697f
C147 B.n67 VSUBS 0.007697f
C148 B.n68 VSUBS 0.007697f
C149 B.n69 VSUBS 0.007697f
C150 B.n70 VSUBS 0.007697f
C151 B.n71 VSUBS 0.007697f
C152 B.n72 VSUBS 0.007697f
C153 B.n73 VSUBS 0.007697f
C154 B.n74 VSUBS 0.007697f
C155 B.n75 VSUBS 0.007697f
C156 B.n76 VSUBS 0.007697f
C157 B.n77 VSUBS 0.018494f
C158 B.n78 VSUBS 0.007697f
C159 B.n79 VSUBS 0.007697f
C160 B.n80 VSUBS 0.007697f
C161 B.n81 VSUBS 0.007697f
C162 B.n82 VSUBS 0.007697f
C163 B.n83 VSUBS 0.007697f
C164 B.n84 VSUBS 0.007697f
C165 B.n85 VSUBS 0.007697f
C166 B.n86 VSUBS 0.007697f
C167 B.n87 VSUBS 0.007697f
C168 B.n88 VSUBS 0.007697f
C169 B.n89 VSUBS 0.007697f
C170 B.n90 VSUBS 0.007697f
C171 B.n91 VSUBS 0.007697f
C172 B.n92 VSUBS 0.007697f
C173 B.n93 VSUBS 0.007697f
C174 B.n94 VSUBS 0.007697f
C175 B.n95 VSUBS 0.019537f
C176 B.n96 VSUBS 0.007697f
C177 B.n97 VSUBS 0.007697f
C178 B.n98 VSUBS 0.007697f
C179 B.n99 VSUBS 0.007697f
C180 B.n100 VSUBS 0.007697f
C181 B.n101 VSUBS 0.007697f
C182 B.n102 VSUBS 0.007697f
C183 B.n103 VSUBS 0.007697f
C184 B.n104 VSUBS 0.007697f
C185 B.n105 VSUBS 0.007697f
C186 B.n106 VSUBS 0.007697f
C187 B.n107 VSUBS 0.007697f
C188 B.n108 VSUBS 0.007697f
C189 B.n109 VSUBS 0.007697f
C190 B.n110 VSUBS 0.007697f
C191 B.n111 VSUBS 0.007697f
C192 B.n112 VSUBS 0.007697f
C193 B.n113 VSUBS 0.007697f
C194 B.n114 VSUBS 0.007697f
C195 B.n115 VSUBS 0.007697f
C196 B.n116 VSUBS 0.007697f
C197 B.n117 VSUBS 0.007697f
C198 B.n118 VSUBS 0.007697f
C199 B.n119 VSUBS 0.007697f
C200 B.n120 VSUBS 0.007697f
C201 B.n121 VSUBS 0.007697f
C202 B.n122 VSUBS 0.007697f
C203 B.n123 VSUBS 0.007697f
C204 B.t2 VSUBS 0.641157f
C205 B.t1 VSUBS 0.650634f
C206 B.t0 VSUBS 0.58748f
C207 B.n124 VSUBS 0.205666f
C208 B.n125 VSUBS 0.070878f
C209 B.n126 VSUBS 0.007697f
C210 B.n127 VSUBS 0.007697f
C211 B.n128 VSUBS 0.007697f
C212 B.n129 VSUBS 0.007697f
C213 B.n130 VSUBS 0.004301f
C214 B.n131 VSUBS 0.007697f
C215 B.n132 VSUBS 0.007697f
C216 B.n133 VSUBS 0.007697f
C217 B.n134 VSUBS 0.007697f
C218 B.n135 VSUBS 0.007697f
C219 B.n136 VSUBS 0.007697f
C220 B.n137 VSUBS 0.007697f
C221 B.n138 VSUBS 0.007697f
C222 B.n139 VSUBS 0.007697f
C223 B.n140 VSUBS 0.007697f
C224 B.n141 VSUBS 0.007697f
C225 B.n142 VSUBS 0.007697f
C226 B.n143 VSUBS 0.007697f
C227 B.n144 VSUBS 0.007697f
C228 B.n145 VSUBS 0.007697f
C229 B.n146 VSUBS 0.007697f
C230 B.n147 VSUBS 0.007697f
C231 B.n148 VSUBS 0.007697f
C232 B.n149 VSUBS 0.007697f
C233 B.n150 VSUBS 0.007697f
C234 B.n151 VSUBS 0.007697f
C235 B.n152 VSUBS 0.007697f
C236 B.n153 VSUBS 0.007697f
C237 B.n154 VSUBS 0.007697f
C238 B.n155 VSUBS 0.007697f
C239 B.n156 VSUBS 0.007697f
C240 B.n157 VSUBS 0.007697f
C241 B.n158 VSUBS 0.007697f
C242 B.n159 VSUBS 0.018494f
C243 B.n160 VSUBS 0.007697f
C244 B.n161 VSUBS 0.007697f
C245 B.n162 VSUBS 0.007697f
C246 B.n163 VSUBS 0.007697f
C247 B.n164 VSUBS 0.007697f
C248 B.n165 VSUBS 0.007697f
C249 B.n166 VSUBS 0.007697f
C250 B.n167 VSUBS 0.007697f
C251 B.n168 VSUBS 0.007697f
C252 B.n169 VSUBS 0.007697f
C253 B.n170 VSUBS 0.007697f
C254 B.n171 VSUBS 0.007697f
C255 B.n172 VSUBS 0.007697f
C256 B.n173 VSUBS 0.007697f
C257 B.n174 VSUBS 0.007697f
C258 B.n175 VSUBS 0.007697f
C259 B.n176 VSUBS 0.007697f
C260 B.n177 VSUBS 0.007697f
C261 B.n178 VSUBS 0.007697f
C262 B.n179 VSUBS 0.007697f
C263 B.n180 VSUBS 0.007697f
C264 B.n181 VSUBS 0.007697f
C265 B.n182 VSUBS 0.007697f
C266 B.n183 VSUBS 0.007697f
C267 B.n184 VSUBS 0.007697f
C268 B.n185 VSUBS 0.007697f
C269 B.n186 VSUBS 0.007697f
C270 B.n187 VSUBS 0.007697f
C271 B.n188 VSUBS 0.007697f
C272 B.n189 VSUBS 0.007697f
C273 B.n190 VSUBS 0.018494f
C274 B.n191 VSUBS 0.019537f
C275 B.n192 VSUBS 0.019537f
C276 B.n193 VSUBS 0.007697f
C277 B.n194 VSUBS 0.007697f
C278 B.n195 VSUBS 0.007697f
C279 B.n196 VSUBS 0.007697f
C280 B.n197 VSUBS 0.007697f
C281 B.n198 VSUBS 0.007697f
C282 B.n199 VSUBS 0.007697f
C283 B.n200 VSUBS 0.007697f
C284 B.n201 VSUBS 0.007697f
C285 B.n202 VSUBS 0.007697f
C286 B.n203 VSUBS 0.007697f
C287 B.n204 VSUBS 0.007697f
C288 B.n205 VSUBS 0.007697f
C289 B.n206 VSUBS 0.007697f
C290 B.n207 VSUBS 0.007697f
C291 B.n208 VSUBS 0.007697f
C292 B.n209 VSUBS 0.007697f
C293 B.n210 VSUBS 0.007697f
C294 B.n211 VSUBS 0.007697f
C295 B.n212 VSUBS 0.007697f
C296 B.n213 VSUBS 0.007697f
C297 B.n214 VSUBS 0.007697f
C298 B.n215 VSUBS 0.007697f
C299 B.n216 VSUBS 0.007697f
C300 B.n217 VSUBS 0.007697f
C301 B.n218 VSUBS 0.007697f
C302 B.n219 VSUBS 0.007697f
C303 B.n220 VSUBS 0.007697f
C304 B.n221 VSUBS 0.007697f
C305 B.n222 VSUBS 0.007697f
C306 B.n223 VSUBS 0.007697f
C307 B.n224 VSUBS 0.007697f
C308 B.n225 VSUBS 0.007697f
C309 B.n226 VSUBS 0.007697f
C310 B.n227 VSUBS 0.007697f
C311 B.n228 VSUBS 0.007697f
C312 B.n229 VSUBS 0.007697f
C313 B.n230 VSUBS 0.007697f
C314 B.n231 VSUBS 0.007697f
C315 B.n232 VSUBS 0.007697f
C316 B.n233 VSUBS 0.007697f
C317 B.n234 VSUBS 0.007697f
C318 B.n235 VSUBS 0.007697f
C319 B.n236 VSUBS 0.007697f
C320 B.n237 VSUBS 0.007697f
C321 B.n238 VSUBS 0.007697f
C322 B.n239 VSUBS 0.007697f
C323 B.n240 VSUBS 0.007697f
C324 B.n241 VSUBS 0.007697f
C325 B.n242 VSUBS 0.007697f
C326 B.n243 VSUBS 0.007697f
C327 B.n244 VSUBS 0.007697f
C328 B.n245 VSUBS 0.007697f
C329 B.n246 VSUBS 0.007697f
C330 B.n247 VSUBS 0.007697f
C331 B.n248 VSUBS 0.007697f
C332 B.n249 VSUBS 0.007697f
C333 B.n250 VSUBS 0.007697f
C334 B.n251 VSUBS 0.007697f
C335 B.n252 VSUBS 0.007697f
C336 B.n253 VSUBS 0.007697f
C337 B.n254 VSUBS 0.007697f
C338 B.n255 VSUBS 0.007697f
C339 B.n256 VSUBS 0.007697f
C340 B.n257 VSUBS 0.007697f
C341 B.n258 VSUBS 0.007697f
C342 B.n259 VSUBS 0.007697f
C343 B.n260 VSUBS 0.007697f
C344 B.n261 VSUBS 0.007697f
C345 B.n262 VSUBS 0.007697f
C346 B.n263 VSUBS 0.007697f
C347 B.n264 VSUBS 0.007697f
C348 B.n265 VSUBS 0.007697f
C349 B.n266 VSUBS 0.007697f
C350 B.n267 VSUBS 0.007697f
C351 B.n268 VSUBS 0.007697f
C352 B.n269 VSUBS 0.007697f
C353 B.n270 VSUBS 0.007697f
C354 B.n271 VSUBS 0.007697f
C355 B.n272 VSUBS 0.007697f
C356 B.n273 VSUBS 0.007697f
C357 B.n274 VSUBS 0.007697f
C358 B.t5 VSUBS 0.641179f
C359 B.t4 VSUBS 0.650654f
C360 B.t3 VSUBS 0.58748f
C361 B.n275 VSUBS 0.205646f
C362 B.n276 VSUBS 0.070856f
C363 B.n277 VSUBS 0.017833f
C364 B.n278 VSUBS 0.007244f
C365 B.n279 VSUBS 0.007697f
C366 B.n280 VSUBS 0.007697f
C367 B.n281 VSUBS 0.007697f
C368 B.n282 VSUBS 0.007697f
C369 B.n283 VSUBS 0.007697f
C370 B.n284 VSUBS 0.007697f
C371 B.n285 VSUBS 0.007697f
C372 B.n286 VSUBS 0.007697f
C373 B.n287 VSUBS 0.007697f
C374 B.n288 VSUBS 0.007697f
C375 B.n289 VSUBS 0.007697f
C376 B.n290 VSUBS 0.007697f
C377 B.n291 VSUBS 0.007697f
C378 B.n292 VSUBS 0.007697f
C379 B.n293 VSUBS 0.007697f
C380 B.n294 VSUBS 0.004301f
C381 B.n295 VSUBS 0.017833f
C382 B.n296 VSUBS 0.007244f
C383 B.n297 VSUBS 0.007697f
C384 B.n298 VSUBS 0.007697f
C385 B.n299 VSUBS 0.007697f
C386 B.n300 VSUBS 0.007697f
C387 B.n301 VSUBS 0.007697f
C388 B.n302 VSUBS 0.007697f
C389 B.n303 VSUBS 0.007697f
C390 B.n304 VSUBS 0.007697f
C391 B.n305 VSUBS 0.007697f
C392 B.n306 VSUBS 0.007697f
C393 B.n307 VSUBS 0.007697f
C394 B.n308 VSUBS 0.007697f
C395 B.n309 VSUBS 0.007697f
C396 B.n310 VSUBS 0.007697f
C397 B.n311 VSUBS 0.007697f
C398 B.n312 VSUBS 0.007697f
C399 B.n313 VSUBS 0.007697f
C400 B.n314 VSUBS 0.007697f
C401 B.n315 VSUBS 0.007697f
C402 B.n316 VSUBS 0.007697f
C403 B.n317 VSUBS 0.007697f
C404 B.n318 VSUBS 0.007697f
C405 B.n319 VSUBS 0.007697f
C406 B.n320 VSUBS 0.007697f
C407 B.n321 VSUBS 0.007697f
C408 B.n322 VSUBS 0.007697f
C409 B.n323 VSUBS 0.007697f
C410 B.n324 VSUBS 0.007697f
C411 B.n325 VSUBS 0.007697f
C412 B.n326 VSUBS 0.007697f
C413 B.n327 VSUBS 0.007697f
C414 B.n328 VSUBS 0.007697f
C415 B.n329 VSUBS 0.007697f
C416 B.n330 VSUBS 0.007697f
C417 B.n331 VSUBS 0.007697f
C418 B.n332 VSUBS 0.007697f
C419 B.n333 VSUBS 0.007697f
C420 B.n334 VSUBS 0.007697f
C421 B.n335 VSUBS 0.007697f
C422 B.n336 VSUBS 0.007697f
C423 B.n337 VSUBS 0.007697f
C424 B.n338 VSUBS 0.007697f
C425 B.n339 VSUBS 0.007697f
C426 B.n340 VSUBS 0.007697f
C427 B.n341 VSUBS 0.007697f
C428 B.n342 VSUBS 0.007697f
C429 B.n343 VSUBS 0.007697f
C430 B.n344 VSUBS 0.007697f
C431 B.n345 VSUBS 0.007697f
C432 B.n346 VSUBS 0.007697f
C433 B.n347 VSUBS 0.007697f
C434 B.n348 VSUBS 0.007697f
C435 B.n349 VSUBS 0.007697f
C436 B.n350 VSUBS 0.007697f
C437 B.n351 VSUBS 0.007697f
C438 B.n352 VSUBS 0.007697f
C439 B.n353 VSUBS 0.007697f
C440 B.n354 VSUBS 0.007697f
C441 B.n355 VSUBS 0.007697f
C442 B.n356 VSUBS 0.007697f
C443 B.n357 VSUBS 0.007697f
C444 B.n358 VSUBS 0.007697f
C445 B.n359 VSUBS 0.007697f
C446 B.n360 VSUBS 0.007697f
C447 B.n361 VSUBS 0.007697f
C448 B.n362 VSUBS 0.007697f
C449 B.n363 VSUBS 0.007697f
C450 B.n364 VSUBS 0.007697f
C451 B.n365 VSUBS 0.007697f
C452 B.n366 VSUBS 0.007697f
C453 B.n367 VSUBS 0.007697f
C454 B.n368 VSUBS 0.007697f
C455 B.n369 VSUBS 0.007697f
C456 B.n370 VSUBS 0.007697f
C457 B.n371 VSUBS 0.007697f
C458 B.n372 VSUBS 0.007697f
C459 B.n373 VSUBS 0.007697f
C460 B.n374 VSUBS 0.007697f
C461 B.n375 VSUBS 0.007697f
C462 B.n376 VSUBS 0.007697f
C463 B.n377 VSUBS 0.007697f
C464 B.n378 VSUBS 0.007697f
C465 B.n379 VSUBS 0.007697f
C466 B.n380 VSUBS 0.018699f
C467 B.n381 VSUBS 0.019332f
C468 B.n382 VSUBS 0.018494f
C469 B.n383 VSUBS 0.007697f
C470 B.n384 VSUBS 0.007697f
C471 B.n385 VSUBS 0.007697f
C472 B.n386 VSUBS 0.007697f
C473 B.n387 VSUBS 0.007697f
C474 B.n388 VSUBS 0.007697f
C475 B.n389 VSUBS 0.007697f
C476 B.n390 VSUBS 0.007697f
C477 B.n391 VSUBS 0.007697f
C478 B.n392 VSUBS 0.007697f
C479 B.n393 VSUBS 0.007697f
C480 B.n394 VSUBS 0.007697f
C481 B.n395 VSUBS 0.007697f
C482 B.n396 VSUBS 0.007697f
C483 B.n397 VSUBS 0.007697f
C484 B.n398 VSUBS 0.007697f
C485 B.n399 VSUBS 0.007697f
C486 B.n400 VSUBS 0.007697f
C487 B.n401 VSUBS 0.007697f
C488 B.n402 VSUBS 0.007697f
C489 B.n403 VSUBS 0.007697f
C490 B.n404 VSUBS 0.007697f
C491 B.n405 VSUBS 0.007697f
C492 B.n406 VSUBS 0.007697f
C493 B.n407 VSUBS 0.007697f
C494 B.n408 VSUBS 0.007697f
C495 B.n409 VSUBS 0.007697f
C496 B.n410 VSUBS 0.007697f
C497 B.n411 VSUBS 0.007697f
C498 B.n412 VSUBS 0.007697f
C499 B.n413 VSUBS 0.007697f
C500 B.n414 VSUBS 0.007697f
C501 B.n415 VSUBS 0.007697f
C502 B.n416 VSUBS 0.007697f
C503 B.n417 VSUBS 0.007697f
C504 B.n418 VSUBS 0.007697f
C505 B.n419 VSUBS 0.007697f
C506 B.n420 VSUBS 0.007697f
C507 B.n421 VSUBS 0.007697f
C508 B.n422 VSUBS 0.007697f
C509 B.n423 VSUBS 0.007697f
C510 B.n424 VSUBS 0.007697f
C511 B.n425 VSUBS 0.007697f
C512 B.n426 VSUBS 0.007697f
C513 B.n427 VSUBS 0.007697f
C514 B.n428 VSUBS 0.007697f
C515 B.n429 VSUBS 0.007697f
C516 B.n430 VSUBS 0.007697f
C517 B.n431 VSUBS 0.007697f
C518 B.n432 VSUBS 0.007697f
C519 B.n433 VSUBS 0.007697f
C520 B.n434 VSUBS 0.018494f
C521 B.n435 VSUBS 0.019537f
C522 B.n436 VSUBS 0.019537f
C523 B.n437 VSUBS 0.007697f
C524 B.n438 VSUBS 0.007697f
C525 B.n439 VSUBS 0.007697f
C526 B.n440 VSUBS 0.007697f
C527 B.n441 VSUBS 0.007697f
C528 B.n442 VSUBS 0.007697f
C529 B.n443 VSUBS 0.007697f
C530 B.n444 VSUBS 0.007697f
C531 B.n445 VSUBS 0.007697f
C532 B.n446 VSUBS 0.007697f
C533 B.n447 VSUBS 0.007697f
C534 B.n448 VSUBS 0.007697f
C535 B.n449 VSUBS 0.007697f
C536 B.n450 VSUBS 0.007697f
C537 B.n451 VSUBS 0.007697f
C538 B.n452 VSUBS 0.007697f
C539 B.n453 VSUBS 0.007697f
C540 B.n454 VSUBS 0.007697f
C541 B.n455 VSUBS 0.007697f
C542 B.n456 VSUBS 0.007697f
C543 B.n457 VSUBS 0.007697f
C544 B.n458 VSUBS 0.007697f
C545 B.n459 VSUBS 0.007697f
C546 B.n460 VSUBS 0.007697f
C547 B.n461 VSUBS 0.007697f
C548 B.n462 VSUBS 0.007697f
C549 B.n463 VSUBS 0.007697f
C550 B.n464 VSUBS 0.007697f
C551 B.n465 VSUBS 0.007697f
C552 B.n466 VSUBS 0.007697f
C553 B.n467 VSUBS 0.007697f
C554 B.n468 VSUBS 0.007697f
C555 B.n469 VSUBS 0.007697f
C556 B.n470 VSUBS 0.007697f
C557 B.n471 VSUBS 0.007697f
C558 B.n472 VSUBS 0.007697f
C559 B.n473 VSUBS 0.007697f
C560 B.n474 VSUBS 0.007697f
C561 B.n475 VSUBS 0.007697f
C562 B.n476 VSUBS 0.007697f
C563 B.n477 VSUBS 0.007697f
C564 B.n478 VSUBS 0.007697f
C565 B.n479 VSUBS 0.007697f
C566 B.n480 VSUBS 0.007697f
C567 B.n481 VSUBS 0.007697f
C568 B.n482 VSUBS 0.007697f
C569 B.n483 VSUBS 0.007697f
C570 B.n484 VSUBS 0.007697f
C571 B.n485 VSUBS 0.007697f
C572 B.n486 VSUBS 0.007697f
C573 B.n487 VSUBS 0.007697f
C574 B.n488 VSUBS 0.007697f
C575 B.n489 VSUBS 0.007697f
C576 B.n490 VSUBS 0.007697f
C577 B.n491 VSUBS 0.007697f
C578 B.n492 VSUBS 0.007697f
C579 B.n493 VSUBS 0.007697f
C580 B.n494 VSUBS 0.007697f
C581 B.n495 VSUBS 0.007697f
C582 B.n496 VSUBS 0.007697f
C583 B.n497 VSUBS 0.007697f
C584 B.n498 VSUBS 0.007697f
C585 B.n499 VSUBS 0.007697f
C586 B.n500 VSUBS 0.007697f
C587 B.n501 VSUBS 0.007697f
C588 B.n502 VSUBS 0.007697f
C589 B.n503 VSUBS 0.007697f
C590 B.n504 VSUBS 0.007697f
C591 B.n505 VSUBS 0.007697f
C592 B.n506 VSUBS 0.007697f
C593 B.n507 VSUBS 0.007697f
C594 B.n508 VSUBS 0.007697f
C595 B.n509 VSUBS 0.007697f
C596 B.n510 VSUBS 0.007697f
C597 B.n511 VSUBS 0.007697f
C598 B.n512 VSUBS 0.007697f
C599 B.n513 VSUBS 0.007697f
C600 B.n514 VSUBS 0.007697f
C601 B.n515 VSUBS 0.007697f
C602 B.n516 VSUBS 0.007697f
C603 B.n517 VSUBS 0.007697f
C604 B.n518 VSUBS 0.007697f
C605 B.n519 VSUBS 0.007244f
C606 B.n520 VSUBS 0.007697f
C607 B.n521 VSUBS 0.007697f
C608 B.n522 VSUBS 0.004301f
C609 B.n523 VSUBS 0.007697f
C610 B.n524 VSUBS 0.007697f
C611 B.n525 VSUBS 0.007697f
C612 B.n526 VSUBS 0.007697f
C613 B.n527 VSUBS 0.007697f
C614 B.n528 VSUBS 0.007697f
C615 B.n529 VSUBS 0.007697f
C616 B.n530 VSUBS 0.007697f
C617 B.n531 VSUBS 0.007697f
C618 B.n532 VSUBS 0.007697f
C619 B.n533 VSUBS 0.007697f
C620 B.n534 VSUBS 0.007697f
C621 B.n535 VSUBS 0.004301f
C622 B.n536 VSUBS 0.017833f
C623 B.n537 VSUBS 0.007244f
C624 B.n538 VSUBS 0.007697f
C625 B.n539 VSUBS 0.007697f
C626 B.n540 VSUBS 0.007697f
C627 B.n541 VSUBS 0.007697f
C628 B.n542 VSUBS 0.007697f
C629 B.n543 VSUBS 0.007697f
C630 B.n544 VSUBS 0.007697f
C631 B.n545 VSUBS 0.007697f
C632 B.n546 VSUBS 0.007697f
C633 B.n547 VSUBS 0.007697f
C634 B.n548 VSUBS 0.007697f
C635 B.n549 VSUBS 0.007697f
C636 B.n550 VSUBS 0.007697f
C637 B.n551 VSUBS 0.007697f
C638 B.n552 VSUBS 0.007697f
C639 B.n553 VSUBS 0.007697f
C640 B.n554 VSUBS 0.007697f
C641 B.n555 VSUBS 0.007697f
C642 B.n556 VSUBS 0.007697f
C643 B.n557 VSUBS 0.007697f
C644 B.n558 VSUBS 0.007697f
C645 B.n559 VSUBS 0.007697f
C646 B.n560 VSUBS 0.007697f
C647 B.n561 VSUBS 0.007697f
C648 B.n562 VSUBS 0.007697f
C649 B.n563 VSUBS 0.007697f
C650 B.n564 VSUBS 0.007697f
C651 B.n565 VSUBS 0.007697f
C652 B.n566 VSUBS 0.007697f
C653 B.n567 VSUBS 0.007697f
C654 B.n568 VSUBS 0.007697f
C655 B.n569 VSUBS 0.007697f
C656 B.n570 VSUBS 0.007697f
C657 B.n571 VSUBS 0.007697f
C658 B.n572 VSUBS 0.007697f
C659 B.n573 VSUBS 0.007697f
C660 B.n574 VSUBS 0.007697f
C661 B.n575 VSUBS 0.007697f
C662 B.n576 VSUBS 0.007697f
C663 B.n577 VSUBS 0.007697f
C664 B.n578 VSUBS 0.007697f
C665 B.n579 VSUBS 0.007697f
C666 B.n580 VSUBS 0.007697f
C667 B.n581 VSUBS 0.007697f
C668 B.n582 VSUBS 0.007697f
C669 B.n583 VSUBS 0.007697f
C670 B.n584 VSUBS 0.007697f
C671 B.n585 VSUBS 0.007697f
C672 B.n586 VSUBS 0.007697f
C673 B.n587 VSUBS 0.007697f
C674 B.n588 VSUBS 0.007697f
C675 B.n589 VSUBS 0.007697f
C676 B.n590 VSUBS 0.007697f
C677 B.n591 VSUBS 0.007697f
C678 B.n592 VSUBS 0.007697f
C679 B.n593 VSUBS 0.007697f
C680 B.n594 VSUBS 0.007697f
C681 B.n595 VSUBS 0.007697f
C682 B.n596 VSUBS 0.007697f
C683 B.n597 VSUBS 0.007697f
C684 B.n598 VSUBS 0.007697f
C685 B.n599 VSUBS 0.007697f
C686 B.n600 VSUBS 0.007697f
C687 B.n601 VSUBS 0.007697f
C688 B.n602 VSUBS 0.007697f
C689 B.n603 VSUBS 0.007697f
C690 B.n604 VSUBS 0.007697f
C691 B.n605 VSUBS 0.007697f
C692 B.n606 VSUBS 0.007697f
C693 B.n607 VSUBS 0.007697f
C694 B.n608 VSUBS 0.007697f
C695 B.n609 VSUBS 0.007697f
C696 B.n610 VSUBS 0.007697f
C697 B.n611 VSUBS 0.007697f
C698 B.n612 VSUBS 0.007697f
C699 B.n613 VSUBS 0.007697f
C700 B.n614 VSUBS 0.007697f
C701 B.n615 VSUBS 0.007697f
C702 B.n616 VSUBS 0.007697f
C703 B.n617 VSUBS 0.007697f
C704 B.n618 VSUBS 0.007697f
C705 B.n619 VSUBS 0.007697f
C706 B.n620 VSUBS 0.007697f
C707 B.n621 VSUBS 0.019537f
C708 B.n622 VSUBS 0.019537f
C709 B.n623 VSUBS 0.018494f
C710 B.n624 VSUBS 0.007697f
C711 B.n625 VSUBS 0.007697f
C712 B.n626 VSUBS 0.007697f
C713 B.n627 VSUBS 0.007697f
C714 B.n628 VSUBS 0.007697f
C715 B.n629 VSUBS 0.007697f
C716 B.n630 VSUBS 0.007697f
C717 B.n631 VSUBS 0.007697f
C718 B.n632 VSUBS 0.007697f
C719 B.n633 VSUBS 0.007697f
C720 B.n634 VSUBS 0.007697f
C721 B.n635 VSUBS 0.007697f
C722 B.n636 VSUBS 0.007697f
C723 B.n637 VSUBS 0.007697f
C724 B.n638 VSUBS 0.007697f
C725 B.n639 VSUBS 0.007697f
C726 B.n640 VSUBS 0.007697f
C727 B.n641 VSUBS 0.007697f
C728 B.n642 VSUBS 0.007697f
C729 B.n643 VSUBS 0.007697f
C730 B.n644 VSUBS 0.007697f
C731 B.n645 VSUBS 0.007697f
C732 B.n646 VSUBS 0.007697f
C733 B.n647 VSUBS 0.010044f
C734 B.n648 VSUBS 0.010699f
C735 B.n649 VSUBS 0.021276f
.ends

