* NGSPICE file created from diff_pair_sample_1546.ext - technology: sky130A

.subckt diff_pair_sample_1546 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0.5577 ps=3.71 w=3.38 l=3.64
X1 VDD1.t9 VP.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X2 VTAIL.t14 VN.t1 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X3 VTAIL.t11 VN.t2 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X4 VTAIL.t19 VN.t3 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X5 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0 ps=0 w=3.38 l=3.64
X6 VTAIL.t13 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X7 VDD1.t8 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0.5577 ps=3.71 w=3.38 l=3.64
X8 VDD2.t4 VN.t5 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X9 VDD1.t7 VP.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=1.3182 ps=7.54 w=3.38 l=3.64
X10 VTAIL.t7 VP.t3 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X11 VDD2.t3 VN.t6 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0.5577 ps=3.71 w=3.38 l=3.64
X12 VDD2.t2 VN.t7 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=1.3182 ps=7.54 w=3.38 l=3.64
X13 VDD1.t5 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X14 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0 ps=0 w=3.38 l=3.64
X15 VDD2.t1 VN.t8 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=1.3182 ps=7.54 w=3.38 l=3.64
X16 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0 ps=0 w=3.38 l=3.64
X17 VTAIL.t6 VP.t5 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X18 VDD1.t3 VP.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=1.3182 ps=7.54 w=3.38 l=3.64
X19 VTAIL.t0 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X20 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0 ps=0 w=3.38 l=3.64
X22 VDD2.t0 VN.t9 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5577 pd=3.71 as=0.5577 ps=3.71 w=3.38 l=3.64
X23 VDD1.t0 VP.t9 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3182 pd=7.54 as=0.5577 ps=3.71 w=3.38 l=3.64
R0 VN.n106 VN.n105 161.3
R1 VN.n104 VN.n55 161.3
R2 VN.n103 VN.n102 161.3
R3 VN.n101 VN.n56 161.3
R4 VN.n100 VN.n99 161.3
R5 VN.n98 VN.n57 161.3
R6 VN.n97 VN.n96 161.3
R7 VN.n95 VN.n58 161.3
R8 VN.n94 VN.n93 161.3
R9 VN.n92 VN.n59 161.3
R10 VN.n91 VN.n90 161.3
R11 VN.n89 VN.n61 161.3
R12 VN.n88 VN.n87 161.3
R13 VN.n86 VN.n62 161.3
R14 VN.n85 VN.n84 161.3
R15 VN.n83 VN.n63 161.3
R16 VN.n82 VN.n81 161.3
R17 VN.n80 VN.n64 161.3
R18 VN.n79 VN.n78 161.3
R19 VN.n77 VN.n66 161.3
R20 VN.n76 VN.n75 161.3
R21 VN.n74 VN.n67 161.3
R22 VN.n73 VN.n72 161.3
R23 VN.n71 VN.n68 161.3
R24 VN.n52 VN.n51 161.3
R25 VN.n50 VN.n1 161.3
R26 VN.n49 VN.n48 161.3
R27 VN.n47 VN.n2 161.3
R28 VN.n46 VN.n45 161.3
R29 VN.n44 VN.n3 161.3
R30 VN.n43 VN.n42 161.3
R31 VN.n41 VN.n4 161.3
R32 VN.n40 VN.n39 161.3
R33 VN.n37 VN.n5 161.3
R34 VN.n36 VN.n35 161.3
R35 VN.n34 VN.n6 161.3
R36 VN.n33 VN.n32 161.3
R37 VN.n31 VN.n7 161.3
R38 VN.n30 VN.n29 161.3
R39 VN.n28 VN.n8 161.3
R40 VN.n27 VN.n26 161.3
R41 VN.n24 VN.n9 161.3
R42 VN.n23 VN.n22 161.3
R43 VN.n21 VN.n10 161.3
R44 VN.n20 VN.n19 161.3
R45 VN.n18 VN.n11 161.3
R46 VN.n17 VN.n16 161.3
R47 VN.n15 VN.n12 161.3
R48 VN.n53 VN.n0 80.9007
R49 VN.n107 VN.n54 80.9007
R50 VN.n14 VN.n13 63.9939
R51 VN.n70 VN.n69 63.9939
R52 VN.n45 VN.n2 56.5617
R53 VN.n99 VN.n56 56.5617
R54 VN.n19 VN.n10 56.5617
R55 VN.n32 VN.n6 56.5617
R56 VN.n75 VN.n66 56.5617
R57 VN.n87 VN.n61 56.5617
R58 VN.n70 VN.t8 55.7439
R59 VN.n14 VN.t0 55.7439
R60 VN VN.n107 52.5171
R61 VN.n17 VN.n12 24.5923
R62 VN.n18 VN.n17 24.5923
R63 VN.n19 VN.n18 24.5923
R64 VN.n23 VN.n10 24.5923
R65 VN.n24 VN.n23 24.5923
R66 VN.n26 VN.n24 24.5923
R67 VN.n30 VN.n8 24.5923
R68 VN.n31 VN.n30 24.5923
R69 VN.n32 VN.n31 24.5923
R70 VN.n36 VN.n6 24.5923
R71 VN.n37 VN.n36 24.5923
R72 VN.n39 VN.n37 24.5923
R73 VN.n43 VN.n4 24.5923
R74 VN.n44 VN.n43 24.5923
R75 VN.n45 VN.n44 24.5923
R76 VN.n49 VN.n2 24.5923
R77 VN.n50 VN.n49 24.5923
R78 VN.n51 VN.n50 24.5923
R79 VN.n75 VN.n74 24.5923
R80 VN.n74 VN.n73 24.5923
R81 VN.n73 VN.n68 24.5923
R82 VN.n87 VN.n86 24.5923
R83 VN.n86 VN.n85 24.5923
R84 VN.n85 VN.n63 24.5923
R85 VN.n81 VN.n80 24.5923
R86 VN.n80 VN.n79 24.5923
R87 VN.n79 VN.n66 24.5923
R88 VN.n99 VN.n98 24.5923
R89 VN.n98 VN.n97 24.5923
R90 VN.n97 VN.n58 24.5923
R91 VN.n93 VN.n92 24.5923
R92 VN.n92 VN.n91 24.5923
R93 VN.n91 VN.n61 24.5923
R94 VN.n105 VN.n104 24.5923
R95 VN.n104 VN.n103 24.5923
R96 VN.n103 VN.n56 24.5923
R97 VN.n13 VN.t2 22.3791
R98 VN.n25 VN.t5 22.3791
R99 VN.n38 VN.t4 22.3791
R100 VN.n0 VN.t7 22.3791
R101 VN.n69 VN.t3 22.3791
R102 VN.n65 VN.t9 22.3791
R103 VN.n60 VN.t1 22.3791
R104 VN.n54 VN.t6 22.3791
R105 VN.n38 VN.n4 13.7719
R106 VN.n60 VN.n58 13.7719
R107 VN.n26 VN.n25 12.2964
R108 VN.n25 VN.n8 12.2964
R109 VN.n65 VN.n63 12.2964
R110 VN.n81 VN.n65 12.2964
R111 VN.n13 VN.n12 10.8209
R112 VN.n39 VN.n38 10.8209
R113 VN.n69 VN.n68 10.8209
R114 VN.n93 VN.n60 10.8209
R115 VN.n51 VN.n0 9.3454
R116 VN.n105 VN.n54 9.3454
R117 VN.n71 VN.n70 3.16706
R118 VN.n15 VN.n14 3.16706
R119 VN.n107 VN.n106 0.354861
R120 VN.n53 VN.n52 0.354861
R121 VN VN.n53 0.267071
R122 VN.n106 VN.n55 0.189894
R123 VN.n102 VN.n55 0.189894
R124 VN.n102 VN.n101 0.189894
R125 VN.n101 VN.n100 0.189894
R126 VN.n100 VN.n57 0.189894
R127 VN.n96 VN.n57 0.189894
R128 VN.n96 VN.n95 0.189894
R129 VN.n95 VN.n94 0.189894
R130 VN.n94 VN.n59 0.189894
R131 VN.n90 VN.n59 0.189894
R132 VN.n90 VN.n89 0.189894
R133 VN.n89 VN.n88 0.189894
R134 VN.n88 VN.n62 0.189894
R135 VN.n84 VN.n62 0.189894
R136 VN.n84 VN.n83 0.189894
R137 VN.n83 VN.n82 0.189894
R138 VN.n82 VN.n64 0.189894
R139 VN.n78 VN.n64 0.189894
R140 VN.n78 VN.n77 0.189894
R141 VN.n77 VN.n76 0.189894
R142 VN.n76 VN.n67 0.189894
R143 VN.n72 VN.n67 0.189894
R144 VN.n72 VN.n71 0.189894
R145 VN.n16 VN.n15 0.189894
R146 VN.n16 VN.n11 0.189894
R147 VN.n20 VN.n11 0.189894
R148 VN.n21 VN.n20 0.189894
R149 VN.n22 VN.n21 0.189894
R150 VN.n22 VN.n9 0.189894
R151 VN.n27 VN.n9 0.189894
R152 VN.n28 VN.n27 0.189894
R153 VN.n29 VN.n28 0.189894
R154 VN.n29 VN.n7 0.189894
R155 VN.n33 VN.n7 0.189894
R156 VN.n34 VN.n33 0.189894
R157 VN.n35 VN.n34 0.189894
R158 VN.n35 VN.n5 0.189894
R159 VN.n40 VN.n5 0.189894
R160 VN.n41 VN.n40 0.189894
R161 VN.n42 VN.n41 0.189894
R162 VN.n42 VN.n3 0.189894
R163 VN.n46 VN.n3 0.189894
R164 VN.n47 VN.n46 0.189894
R165 VN.n48 VN.n47 0.189894
R166 VN.n48 VN.n1 0.189894
R167 VN.n52 VN.n1 0.189894
R168 VTAIL.n72 VTAIL.n62 289.615
R169 VTAIL.n12 VTAIL.n2 289.615
R170 VTAIL.n56 VTAIL.n46 289.615
R171 VTAIL.n36 VTAIL.n26 289.615
R172 VTAIL.n66 VTAIL.n65 185
R173 VTAIL.n71 VTAIL.n70 185
R174 VTAIL.n73 VTAIL.n72 185
R175 VTAIL.n6 VTAIL.n5 185
R176 VTAIL.n11 VTAIL.n10 185
R177 VTAIL.n13 VTAIL.n12 185
R178 VTAIL.n57 VTAIL.n56 185
R179 VTAIL.n55 VTAIL.n54 185
R180 VTAIL.n50 VTAIL.n49 185
R181 VTAIL.n37 VTAIL.n36 185
R182 VTAIL.n35 VTAIL.n34 185
R183 VTAIL.n30 VTAIL.n29 185
R184 VTAIL.n67 VTAIL.t15 150.499
R185 VTAIL.n7 VTAIL.t8 150.499
R186 VTAIL.n31 VTAIL.t10 150.499
R187 VTAIL.n51 VTAIL.t3 150.499
R188 VTAIL.n71 VTAIL.n65 104.615
R189 VTAIL.n72 VTAIL.n71 104.615
R190 VTAIL.n11 VTAIL.n5 104.615
R191 VTAIL.n12 VTAIL.n11 104.615
R192 VTAIL.n56 VTAIL.n55 104.615
R193 VTAIL.n55 VTAIL.n49 104.615
R194 VTAIL.n36 VTAIL.n35 104.615
R195 VTAIL.n35 VTAIL.n29 104.615
R196 VTAIL.n45 VTAIL.n44 60.2527
R197 VTAIL.n43 VTAIL.n42 60.2527
R198 VTAIL.n25 VTAIL.n24 60.2527
R199 VTAIL.n23 VTAIL.n22 60.2527
R200 VTAIL.n79 VTAIL.n78 60.2527
R201 VTAIL.n1 VTAIL.n0 60.2527
R202 VTAIL.n19 VTAIL.n18 60.2527
R203 VTAIL.n21 VTAIL.n20 60.2527
R204 VTAIL.t15 VTAIL.n65 52.3082
R205 VTAIL.t8 VTAIL.n5 52.3082
R206 VTAIL.t3 VTAIL.n49 52.3082
R207 VTAIL.t10 VTAIL.n29 52.3082
R208 VTAIL.n77 VTAIL.n76 30.246
R209 VTAIL.n17 VTAIL.n16 30.246
R210 VTAIL.n61 VTAIL.n60 30.246
R211 VTAIL.n41 VTAIL.n40 30.246
R212 VTAIL.n23 VTAIL.n21 22.1255
R213 VTAIL.n77 VTAIL.n61 18.7031
R214 VTAIL.n67 VTAIL.n66 10.2326
R215 VTAIL.n7 VTAIL.n6 10.2326
R216 VTAIL.n51 VTAIL.n50 10.2326
R217 VTAIL.n31 VTAIL.n30 10.2326
R218 VTAIL.n76 VTAIL.n62 9.69747
R219 VTAIL.n16 VTAIL.n2 9.69747
R220 VTAIL.n60 VTAIL.n46 9.69747
R221 VTAIL.n40 VTAIL.n26 9.69747
R222 VTAIL.n76 VTAIL.n75 9.45567
R223 VTAIL.n16 VTAIL.n15 9.45567
R224 VTAIL.n60 VTAIL.n59 9.45567
R225 VTAIL.n40 VTAIL.n39 9.45567
R226 VTAIL.n69 VTAIL.n68 9.3005
R227 VTAIL.n64 VTAIL.n63 9.3005
R228 VTAIL.n75 VTAIL.n74 9.3005
R229 VTAIL.n9 VTAIL.n8 9.3005
R230 VTAIL.n4 VTAIL.n3 9.3005
R231 VTAIL.n15 VTAIL.n14 9.3005
R232 VTAIL.n48 VTAIL.n47 9.3005
R233 VTAIL.n53 VTAIL.n52 9.3005
R234 VTAIL.n59 VTAIL.n58 9.3005
R235 VTAIL.n28 VTAIL.n27 9.3005
R236 VTAIL.n39 VTAIL.n38 9.3005
R237 VTAIL.n33 VTAIL.n32 9.3005
R238 VTAIL.n74 VTAIL.n73 8.92171
R239 VTAIL.n14 VTAIL.n13 8.92171
R240 VTAIL.n58 VTAIL.n57 8.92171
R241 VTAIL.n38 VTAIL.n37 8.92171
R242 VTAIL.n70 VTAIL.n64 8.14595
R243 VTAIL.n10 VTAIL.n4 8.14595
R244 VTAIL.n54 VTAIL.n48 8.14595
R245 VTAIL.n34 VTAIL.n28 8.14595
R246 VTAIL.n69 VTAIL.n66 7.3702
R247 VTAIL.n9 VTAIL.n6 7.3702
R248 VTAIL.n53 VTAIL.n50 7.3702
R249 VTAIL.n33 VTAIL.n30 7.3702
R250 VTAIL.n78 VTAIL.t12 5.85849
R251 VTAIL.n78 VTAIL.t13 5.85849
R252 VTAIL.n0 VTAIL.t16 5.85849
R253 VTAIL.n0 VTAIL.t11 5.85849
R254 VTAIL.n18 VTAIL.t4 5.85849
R255 VTAIL.n18 VTAIL.t6 5.85849
R256 VTAIL.n20 VTAIL.t5 5.85849
R257 VTAIL.n20 VTAIL.t0 5.85849
R258 VTAIL.n44 VTAIL.t9 5.85849
R259 VTAIL.n44 VTAIL.t7 5.85849
R260 VTAIL.n42 VTAIL.t2 5.85849
R261 VTAIL.n42 VTAIL.t1 5.85849
R262 VTAIL.n24 VTAIL.t18 5.85849
R263 VTAIL.n24 VTAIL.t19 5.85849
R264 VTAIL.n22 VTAIL.t17 5.85849
R265 VTAIL.n22 VTAIL.t14 5.85849
R266 VTAIL.n70 VTAIL.n69 5.81868
R267 VTAIL.n10 VTAIL.n9 5.81868
R268 VTAIL.n54 VTAIL.n53 5.81868
R269 VTAIL.n34 VTAIL.n33 5.81868
R270 VTAIL.n73 VTAIL.n64 5.04292
R271 VTAIL.n13 VTAIL.n4 5.04292
R272 VTAIL.n57 VTAIL.n48 5.04292
R273 VTAIL.n37 VTAIL.n28 5.04292
R274 VTAIL.n74 VTAIL.n62 4.26717
R275 VTAIL.n14 VTAIL.n2 4.26717
R276 VTAIL.n58 VTAIL.n46 4.26717
R277 VTAIL.n38 VTAIL.n26 4.26717
R278 VTAIL.n25 VTAIL.n23 3.42291
R279 VTAIL.n41 VTAIL.n25 3.42291
R280 VTAIL.n45 VTAIL.n43 3.42291
R281 VTAIL.n61 VTAIL.n45 3.42291
R282 VTAIL.n21 VTAIL.n19 3.42291
R283 VTAIL.n19 VTAIL.n17 3.42291
R284 VTAIL.n79 VTAIL.n77 3.42291
R285 VTAIL.n68 VTAIL.n67 2.88718
R286 VTAIL.n8 VTAIL.n7 2.88718
R287 VTAIL.n52 VTAIL.n51 2.88718
R288 VTAIL.n32 VTAIL.n31 2.88718
R289 VTAIL VTAIL.n1 2.6255
R290 VTAIL.n43 VTAIL.n41 2.18153
R291 VTAIL.n17 VTAIL.n1 2.18153
R292 VTAIL VTAIL.n79 0.797914
R293 VTAIL.n68 VTAIL.n63 0.155672
R294 VTAIL.n75 VTAIL.n63 0.155672
R295 VTAIL.n8 VTAIL.n3 0.155672
R296 VTAIL.n15 VTAIL.n3 0.155672
R297 VTAIL.n59 VTAIL.n47 0.155672
R298 VTAIL.n52 VTAIL.n47 0.155672
R299 VTAIL.n39 VTAIL.n27 0.155672
R300 VTAIL.n32 VTAIL.n27 0.155672
R301 VDD2.n29 VDD2.n19 289.615
R302 VDD2.n10 VDD2.n0 289.615
R303 VDD2.n30 VDD2.n29 185
R304 VDD2.n28 VDD2.n27 185
R305 VDD2.n23 VDD2.n22 185
R306 VDD2.n4 VDD2.n3 185
R307 VDD2.n9 VDD2.n8 185
R308 VDD2.n11 VDD2.n10 185
R309 VDD2.n24 VDD2.t3 150.499
R310 VDD2.n5 VDD2.t9 150.499
R311 VDD2.n29 VDD2.n28 104.615
R312 VDD2.n28 VDD2.n22 104.615
R313 VDD2.n9 VDD2.n3 104.615
R314 VDD2.n10 VDD2.n9 104.615
R315 VDD2.n18 VDD2.n17 79.443
R316 VDD2 VDD2.n37 79.4401
R317 VDD2.n36 VDD2.n35 76.9315
R318 VDD2.n16 VDD2.n15 76.9315
R319 VDD2.t3 VDD2.n22 52.3082
R320 VDD2.t9 VDD2.n3 52.3082
R321 VDD2.n16 VDD2.n14 50.3472
R322 VDD2.n34 VDD2.n33 46.9247
R323 VDD2.n34 VDD2.n18 42.8856
R324 VDD2.n24 VDD2.n23 10.2326
R325 VDD2.n5 VDD2.n4 10.2326
R326 VDD2.n33 VDD2.n19 9.69747
R327 VDD2.n14 VDD2.n0 9.69747
R328 VDD2.n33 VDD2.n32 9.45567
R329 VDD2.n14 VDD2.n13 9.45567
R330 VDD2.n21 VDD2.n20 9.3005
R331 VDD2.n32 VDD2.n31 9.3005
R332 VDD2.n26 VDD2.n25 9.3005
R333 VDD2.n7 VDD2.n6 9.3005
R334 VDD2.n2 VDD2.n1 9.3005
R335 VDD2.n13 VDD2.n12 9.3005
R336 VDD2.n31 VDD2.n30 8.92171
R337 VDD2.n12 VDD2.n11 8.92171
R338 VDD2.n27 VDD2.n21 8.14595
R339 VDD2.n8 VDD2.n2 8.14595
R340 VDD2.n26 VDD2.n23 7.3702
R341 VDD2.n7 VDD2.n4 7.3702
R342 VDD2.n37 VDD2.t6 5.85849
R343 VDD2.n37 VDD2.t1 5.85849
R344 VDD2.n35 VDD2.t8 5.85849
R345 VDD2.n35 VDD2.t0 5.85849
R346 VDD2.n17 VDD2.t5 5.85849
R347 VDD2.n17 VDD2.t2 5.85849
R348 VDD2.n15 VDD2.t7 5.85849
R349 VDD2.n15 VDD2.t4 5.85849
R350 VDD2.n27 VDD2.n26 5.81868
R351 VDD2.n8 VDD2.n7 5.81868
R352 VDD2.n30 VDD2.n21 5.04292
R353 VDD2.n11 VDD2.n2 5.04292
R354 VDD2.n31 VDD2.n19 4.26717
R355 VDD2.n12 VDD2.n0 4.26717
R356 VDD2.n36 VDD2.n34 3.42291
R357 VDD2.n25 VDD2.n24 2.88718
R358 VDD2.n6 VDD2.n5 2.88718
R359 VDD2 VDD2.n36 0.914293
R360 VDD2.n18 VDD2.n16 0.800757
R361 VDD2.n32 VDD2.n20 0.155672
R362 VDD2.n25 VDD2.n20 0.155672
R363 VDD2.n6 VDD2.n1 0.155672
R364 VDD2.n13 VDD2.n1 0.155672
R365 B.n765 B.n764 585
R366 B.n767 B.n167 585
R367 B.n770 B.n769 585
R368 B.n771 B.n166 585
R369 B.n773 B.n772 585
R370 B.n775 B.n165 585
R371 B.n778 B.n777 585
R372 B.n779 B.n164 585
R373 B.n781 B.n780 585
R374 B.n783 B.n163 585
R375 B.n786 B.n785 585
R376 B.n787 B.n162 585
R377 B.n789 B.n788 585
R378 B.n791 B.n161 585
R379 B.n793 B.n792 585
R380 B.n795 B.n794 585
R381 B.n798 B.n797 585
R382 B.n799 B.n156 585
R383 B.n801 B.n800 585
R384 B.n803 B.n155 585
R385 B.n806 B.n805 585
R386 B.n807 B.n154 585
R387 B.n809 B.n808 585
R388 B.n811 B.n153 585
R389 B.n814 B.n813 585
R390 B.n815 B.n150 585
R391 B.n818 B.n817 585
R392 B.n820 B.n149 585
R393 B.n823 B.n822 585
R394 B.n824 B.n148 585
R395 B.n826 B.n825 585
R396 B.n828 B.n147 585
R397 B.n831 B.n830 585
R398 B.n832 B.n146 585
R399 B.n834 B.n833 585
R400 B.n836 B.n145 585
R401 B.n839 B.n838 585
R402 B.n840 B.n144 585
R403 B.n842 B.n841 585
R404 B.n844 B.n143 585
R405 B.n847 B.n846 585
R406 B.n848 B.n142 585
R407 B.n763 B.n140 585
R408 B.n851 B.n140 585
R409 B.n762 B.n139 585
R410 B.n852 B.n139 585
R411 B.n761 B.n138 585
R412 B.n853 B.n138 585
R413 B.n760 B.n759 585
R414 B.n759 B.n134 585
R415 B.n758 B.n133 585
R416 B.n859 B.n133 585
R417 B.n757 B.n132 585
R418 B.n860 B.n132 585
R419 B.n756 B.n131 585
R420 B.n861 B.n131 585
R421 B.n755 B.n754 585
R422 B.n754 B.n127 585
R423 B.n753 B.n126 585
R424 B.n867 B.n126 585
R425 B.n752 B.n125 585
R426 B.n868 B.n125 585
R427 B.n751 B.n124 585
R428 B.n869 B.n124 585
R429 B.n750 B.n749 585
R430 B.n749 B.n120 585
R431 B.n748 B.n119 585
R432 B.n875 B.n119 585
R433 B.n747 B.n118 585
R434 B.n876 B.n118 585
R435 B.n746 B.n117 585
R436 B.n877 B.n117 585
R437 B.n745 B.n744 585
R438 B.n744 B.n113 585
R439 B.n743 B.n112 585
R440 B.n883 B.n112 585
R441 B.n742 B.n111 585
R442 B.n884 B.n111 585
R443 B.n741 B.n110 585
R444 B.n885 B.n110 585
R445 B.n740 B.n739 585
R446 B.n739 B.n106 585
R447 B.n738 B.n105 585
R448 B.n891 B.n105 585
R449 B.n737 B.n104 585
R450 B.n892 B.n104 585
R451 B.n736 B.n103 585
R452 B.n893 B.n103 585
R453 B.n735 B.n734 585
R454 B.n734 B.n102 585
R455 B.n733 B.n98 585
R456 B.n899 B.n98 585
R457 B.n732 B.n97 585
R458 B.n900 B.n97 585
R459 B.n731 B.n96 585
R460 B.n901 B.n96 585
R461 B.n730 B.n729 585
R462 B.n729 B.n92 585
R463 B.n728 B.n91 585
R464 B.n907 B.n91 585
R465 B.n727 B.n90 585
R466 B.n908 B.n90 585
R467 B.n726 B.n89 585
R468 B.n909 B.n89 585
R469 B.n725 B.n724 585
R470 B.n724 B.n85 585
R471 B.n723 B.n84 585
R472 B.n915 B.n84 585
R473 B.n722 B.n83 585
R474 B.n916 B.n83 585
R475 B.n721 B.n82 585
R476 B.n917 B.n82 585
R477 B.n720 B.n719 585
R478 B.n719 B.n81 585
R479 B.n718 B.n77 585
R480 B.n923 B.n77 585
R481 B.n717 B.n76 585
R482 B.n924 B.n76 585
R483 B.n716 B.n75 585
R484 B.n925 B.n75 585
R485 B.n715 B.n714 585
R486 B.n714 B.n71 585
R487 B.n713 B.n70 585
R488 B.n931 B.n70 585
R489 B.n712 B.n69 585
R490 B.n932 B.n69 585
R491 B.n711 B.n68 585
R492 B.n933 B.n68 585
R493 B.n710 B.n709 585
R494 B.n709 B.n64 585
R495 B.n708 B.n63 585
R496 B.n939 B.n63 585
R497 B.n707 B.n62 585
R498 B.n940 B.n62 585
R499 B.n706 B.n61 585
R500 B.n941 B.n61 585
R501 B.n705 B.n704 585
R502 B.n704 B.n60 585
R503 B.n703 B.n56 585
R504 B.n947 B.n56 585
R505 B.n702 B.n55 585
R506 B.n948 B.n55 585
R507 B.n701 B.n54 585
R508 B.n949 B.n54 585
R509 B.n700 B.n699 585
R510 B.n699 B.n50 585
R511 B.n698 B.n49 585
R512 B.n955 B.n49 585
R513 B.n697 B.n48 585
R514 B.n956 B.n48 585
R515 B.n696 B.n47 585
R516 B.n957 B.n47 585
R517 B.n695 B.n694 585
R518 B.n694 B.n43 585
R519 B.n693 B.n42 585
R520 B.n963 B.n42 585
R521 B.n692 B.n41 585
R522 B.n964 B.n41 585
R523 B.n691 B.n40 585
R524 B.n965 B.n40 585
R525 B.n690 B.n689 585
R526 B.n689 B.n36 585
R527 B.n688 B.n35 585
R528 B.n971 B.n35 585
R529 B.n687 B.n34 585
R530 B.n972 B.n34 585
R531 B.n686 B.n33 585
R532 B.n973 B.n33 585
R533 B.n685 B.n684 585
R534 B.n684 B.n29 585
R535 B.n683 B.n28 585
R536 B.n979 B.n28 585
R537 B.n682 B.n27 585
R538 B.n980 B.n27 585
R539 B.n681 B.n26 585
R540 B.n981 B.n26 585
R541 B.n680 B.n679 585
R542 B.n679 B.n22 585
R543 B.n678 B.n21 585
R544 B.n987 B.n21 585
R545 B.n677 B.n20 585
R546 B.n988 B.n20 585
R547 B.n676 B.n19 585
R548 B.n989 B.n19 585
R549 B.n675 B.n674 585
R550 B.n674 B.n15 585
R551 B.n673 B.n14 585
R552 B.n995 B.n14 585
R553 B.n672 B.n13 585
R554 B.n996 B.n13 585
R555 B.n671 B.n12 585
R556 B.n997 B.n12 585
R557 B.n670 B.n669 585
R558 B.n669 B.n8 585
R559 B.n668 B.n7 585
R560 B.n1003 B.n7 585
R561 B.n667 B.n6 585
R562 B.n1004 B.n6 585
R563 B.n666 B.n5 585
R564 B.n1005 B.n5 585
R565 B.n665 B.n664 585
R566 B.n664 B.n4 585
R567 B.n663 B.n168 585
R568 B.n663 B.n662 585
R569 B.n653 B.n169 585
R570 B.n170 B.n169 585
R571 B.n655 B.n654 585
R572 B.n656 B.n655 585
R573 B.n652 B.n175 585
R574 B.n175 B.n174 585
R575 B.n651 B.n650 585
R576 B.n650 B.n649 585
R577 B.n177 B.n176 585
R578 B.n178 B.n177 585
R579 B.n642 B.n641 585
R580 B.n643 B.n642 585
R581 B.n640 B.n183 585
R582 B.n183 B.n182 585
R583 B.n639 B.n638 585
R584 B.n638 B.n637 585
R585 B.n185 B.n184 585
R586 B.n186 B.n185 585
R587 B.n630 B.n629 585
R588 B.n631 B.n630 585
R589 B.n628 B.n191 585
R590 B.n191 B.n190 585
R591 B.n627 B.n626 585
R592 B.n626 B.n625 585
R593 B.n193 B.n192 585
R594 B.n194 B.n193 585
R595 B.n618 B.n617 585
R596 B.n619 B.n618 585
R597 B.n616 B.n199 585
R598 B.n199 B.n198 585
R599 B.n615 B.n614 585
R600 B.n614 B.n613 585
R601 B.n201 B.n200 585
R602 B.n202 B.n201 585
R603 B.n606 B.n605 585
R604 B.n607 B.n606 585
R605 B.n604 B.n207 585
R606 B.n207 B.n206 585
R607 B.n603 B.n602 585
R608 B.n602 B.n601 585
R609 B.n209 B.n208 585
R610 B.n210 B.n209 585
R611 B.n594 B.n593 585
R612 B.n595 B.n594 585
R613 B.n592 B.n215 585
R614 B.n215 B.n214 585
R615 B.n591 B.n590 585
R616 B.n590 B.n589 585
R617 B.n217 B.n216 585
R618 B.n218 B.n217 585
R619 B.n582 B.n581 585
R620 B.n583 B.n582 585
R621 B.n580 B.n223 585
R622 B.n223 B.n222 585
R623 B.n579 B.n578 585
R624 B.n578 B.n577 585
R625 B.n225 B.n224 585
R626 B.n570 B.n225 585
R627 B.n569 B.n568 585
R628 B.n571 B.n569 585
R629 B.n567 B.n230 585
R630 B.n230 B.n229 585
R631 B.n566 B.n565 585
R632 B.n565 B.n564 585
R633 B.n232 B.n231 585
R634 B.n233 B.n232 585
R635 B.n557 B.n556 585
R636 B.n558 B.n557 585
R637 B.n555 B.n238 585
R638 B.n238 B.n237 585
R639 B.n554 B.n553 585
R640 B.n553 B.n552 585
R641 B.n240 B.n239 585
R642 B.n241 B.n240 585
R643 B.n545 B.n544 585
R644 B.n546 B.n545 585
R645 B.n543 B.n246 585
R646 B.n246 B.n245 585
R647 B.n542 B.n541 585
R648 B.n541 B.n540 585
R649 B.n248 B.n247 585
R650 B.n533 B.n248 585
R651 B.n532 B.n531 585
R652 B.n534 B.n532 585
R653 B.n530 B.n253 585
R654 B.n253 B.n252 585
R655 B.n529 B.n528 585
R656 B.n528 B.n527 585
R657 B.n255 B.n254 585
R658 B.n256 B.n255 585
R659 B.n520 B.n519 585
R660 B.n521 B.n520 585
R661 B.n518 B.n261 585
R662 B.n261 B.n260 585
R663 B.n517 B.n516 585
R664 B.n516 B.n515 585
R665 B.n263 B.n262 585
R666 B.n264 B.n263 585
R667 B.n508 B.n507 585
R668 B.n509 B.n508 585
R669 B.n506 B.n269 585
R670 B.n269 B.n268 585
R671 B.n505 B.n504 585
R672 B.n504 B.n503 585
R673 B.n271 B.n270 585
R674 B.n496 B.n271 585
R675 B.n495 B.n494 585
R676 B.n497 B.n495 585
R677 B.n493 B.n276 585
R678 B.n276 B.n275 585
R679 B.n492 B.n491 585
R680 B.n491 B.n490 585
R681 B.n278 B.n277 585
R682 B.n279 B.n278 585
R683 B.n483 B.n482 585
R684 B.n484 B.n483 585
R685 B.n481 B.n284 585
R686 B.n284 B.n283 585
R687 B.n480 B.n479 585
R688 B.n479 B.n478 585
R689 B.n286 B.n285 585
R690 B.n287 B.n286 585
R691 B.n471 B.n470 585
R692 B.n472 B.n471 585
R693 B.n469 B.n292 585
R694 B.n292 B.n291 585
R695 B.n468 B.n467 585
R696 B.n467 B.n466 585
R697 B.n294 B.n293 585
R698 B.n295 B.n294 585
R699 B.n459 B.n458 585
R700 B.n460 B.n459 585
R701 B.n457 B.n300 585
R702 B.n300 B.n299 585
R703 B.n456 B.n455 585
R704 B.n455 B.n454 585
R705 B.n302 B.n301 585
R706 B.n303 B.n302 585
R707 B.n447 B.n446 585
R708 B.n448 B.n447 585
R709 B.n445 B.n308 585
R710 B.n308 B.n307 585
R711 B.n444 B.n443 585
R712 B.n443 B.n442 585
R713 B.n310 B.n309 585
R714 B.n311 B.n310 585
R715 B.n435 B.n434 585
R716 B.n436 B.n435 585
R717 B.n433 B.n316 585
R718 B.n316 B.n315 585
R719 B.n432 B.n431 585
R720 B.n431 B.n430 585
R721 B.n427 B.n320 585
R722 B.n426 B.n425 585
R723 B.n423 B.n321 585
R724 B.n423 B.n319 585
R725 B.n422 B.n421 585
R726 B.n420 B.n419 585
R727 B.n418 B.n323 585
R728 B.n416 B.n415 585
R729 B.n414 B.n324 585
R730 B.n413 B.n412 585
R731 B.n410 B.n325 585
R732 B.n408 B.n407 585
R733 B.n406 B.n326 585
R734 B.n405 B.n404 585
R735 B.n402 B.n327 585
R736 B.n400 B.n399 585
R737 B.n398 B.n328 585
R738 B.n396 B.n395 585
R739 B.n393 B.n331 585
R740 B.n391 B.n390 585
R741 B.n389 B.n332 585
R742 B.n388 B.n387 585
R743 B.n385 B.n333 585
R744 B.n383 B.n382 585
R745 B.n381 B.n334 585
R746 B.n380 B.n379 585
R747 B.n377 B.n335 585
R748 B.n375 B.n374 585
R749 B.n373 B.n336 585
R750 B.n372 B.n371 585
R751 B.n369 B.n340 585
R752 B.n367 B.n366 585
R753 B.n365 B.n341 585
R754 B.n364 B.n363 585
R755 B.n361 B.n342 585
R756 B.n359 B.n358 585
R757 B.n357 B.n343 585
R758 B.n356 B.n355 585
R759 B.n353 B.n344 585
R760 B.n351 B.n350 585
R761 B.n349 B.n345 585
R762 B.n348 B.n347 585
R763 B.n318 B.n317 585
R764 B.n319 B.n318 585
R765 B.n429 B.n428 585
R766 B.n430 B.n429 585
R767 B.n314 B.n313 585
R768 B.n315 B.n314 585
R769 B.n438 B.n437 585
R770 B.n437 B.n436 585
R771 B.n439 B.n312 585
R772 B.n312 B.n311 585
R773 B.n441 B.n440 585
R774 B.n442 B.n441 585
R775 B.n306 B.n305 585
R776 B.n307 B.n306 585
R777 B.n450 B.n449 585
R778 B.n449 B.n448 585
R779 B.n451 B.n304 585
R780 B.n304 B.n303 585
R781 B.n453 B.n452 585
R782 B.n454 B.n453 585
R783 B.n298 B.n297 585
R784 B.n299 B.n298 585
R785 B.n462 B.n461 585
R786 B.n461 B.n460 585
R787 B.n463 B.n296 585
R788 B.n296 B.n295 585
R789 B.n465 B.n464 585
R790 B.n466 B.n465 585
R791 B.n290 B.n289 585
R792 B.n291 B.n290 585
R793 B.n474 B.n473 585
R794 B.n473 B.n472 585
R795 B.n475 B.n288 585
R796 B.n288 B.n287 585
R797 B.n477 B.n476 585
R798 B.n478 B.n477 585
R799 B.n282 B.n281 585
R800 B.n283 B.n282 585
R801 B.n486 B.n485 585
R802 B.n485 B.n484 585
R803 B.n487 B.n280 585
R804 B.n280 B.n279 585
R805 B.n489 B.n488 585
R806 B.n490 B.n489 585
R807 B.n274 B.n273 585
R808 B.n275 B.n274 585
R809 B.n499 B.n498 585
R810 B.n498 B.n497 585
R811 B.n500 B.n272 585
R812 B.n496 B.n272 585
R813 B.n502 B.n501 585
R814 B.n503 B.n502 585
R815 B.n267 B.n266 585
R816 B.n268 B.n267 585
R817 B.n511 B.n510 585
R818 B.n510 B.n509 585
R819 B.n512 B.n265 585
R820 B.n265 B.n264 585
R821 B.n514 B.n513 585
R822 B.n515 B.n514 585
R823 B.n259 B.n258 585
R824 B.n260 B.n259 585
R825 B.n523 B.n522 585
R826 B.n522 B.n521 585
R827 B.n524 B.n257 585
R828 B.n257 B.n256 585
R829 B.n526 B.n525 585
R830 B.n527 B.n526 585
R831 B.n251 B.n250 585
R832 B.n252 B.n251 585
R833 B.n536 B.n535 585
R834 B.n535 B.n534 585
R835 B.n537 B.n249 585
R836 B.n533 B.n249 585
R837 B.n539 B.n538 585
R838 B.n540 B.n539 585
R839 B.n244 B.n243 585
R840 B.n245 B.n244 585
R841 B.n548 B.n547 585
R842 B.n547 B.n546 585
R843 B.n549 B.n242 585
R844 B.n242 B.n241 585
R845 B.n551 B.n550 585
R846 B.n552 B.n551 585
R847 B.n236 B.n235 585
R848 B.n237 B.n236 585
R849 B.n560 B.n559 585
R850 B.n559 B.n558 585
R851 B.n561 B.n234 585
R852 B.n234 B.n233 585
R853 B.n563 B.n562 585
R854 B.n564 B.n563 585
R855 B.n228 B.n227 585
R856 B.n229 B.n228 585
R857 B.n573 B.n572 585
R858 B.n572 B.n571 585
R859 B.n574 B.n226 585
R860 B.n570 B.n226 585
R861 B.n576 B.n575 585
R862 B.n577 B.n576 585
R863 B.n221 B.n220 585
R864 B.n222 B.n221 585
R865 B.n585 B.n584 585
R866 B.n584 B.n583 585
R867 B.n586 B.n219 585
R868 B.n219 B.n218 585
R869 B.n588 B.n587 585
R870 B.n589 B.n588 585
R871 B.n213 B.n212 585
R872 B.n214 B.n213 585
R873 B.n597 B.n596 585
R874 B.n596 B.n595 585
R875 B.n598 B.n211 585
R876 B.n211 B.n210 585
R877 B.n600 B.n599 585
R878 B.n601 B.n600 585
R879 B.n205 B.n204 585
R880 B.n206 B.n205 585
R881 B.n609 B.n608 585
R882 B.n608 B.n607 585
R883 B.n610 B.n203 585
R884 B.n203 B.n202 585
R885 B.n612 B.n611 585
R886 B.n613 B.n612 585
R887 B.n197 B.n196 585
R888 B.n198 B.n197 585
R889 B.n621 B.n620 585
R890 B.n620 B.n619 585
R891 B.n622 B.n195 585
R892 B.n195 B.n194 585
R893 B.n624 B.n623 585
R894 B.n625 B.n624 585
R895 B.n189 B.n188 585
R896 B.n190 B.n189 585
R897 B.n633 B.n632 585
R898 B.n632 B.n631 585
R899 B.n634 B.n187 585
R900 B.n187 B.n186 585
R901 B.n636 B.n635 585
R902 B.n637 B.n636 585
R903 B.n181 B.n180 585
R904 B.n182 B.n181 585
R905 B.n645 B.n644 585
R906 B.n644 B.n643 585
R907 B.n646 B.n179 585
R908 B.n179 B.n178 585
R909 B.n648 B.n647 585
R910 B.n649 B.n648 585
R911 B.n173 B.n172 585
R912 B.n174 B.n173 585
R913 B.n658 B.n657 585
R914 B.n657 B.n656 585
R915 B.n659 B.n171 585
R916 B.n171 B.n170 585
R917 B.n661 B.n660 585
R918 B.n662 B.n661 585
R919 B.n2 B.n0 585
R920 B.n4 B.n2 585
R921 B.n3 B.n1 585
R922 B.n1004 B.n3 585
R923 B.n1002 B.n1001 585
R924 B.n1003 B.n1002 585
R925 B.n1000 B.n9 585
R926 B.n9 B.n8 585
R927 B.n999 B.n998 585
R928 B.n998 B.n997 585
R929 B.n11 B.n10 585
R930 B.n996 B.n11 585
R931 B.n994 B.n993 585
R932 B.n995 B.n994 585
R933 B.n992 B.n16 585
R934 B.n16 B.n15 585
R935 B.n991 B.n990 585
R936 B.n990 B.n989 585
R937 B.n18 B.n17 585
R938 B.n988 B.n18 585
R939 B.n986 B.n985 585
R940 B.n987 B.n986 585
R941 B.n984 B.n23 585
R942 B.n23 B.n22 585
R943 B.n983 B.n982 585
R944 B.n982 B.n981 585
R945 B.n25 B.n24 585
R946 B.n980 B.n25 585
R947 B.n978 B.n977 585
R948 B.n979 B.n978 585
R949 B.n976 B.n30 585
R950 B.n30 B.n29 585
R951 B.n975 B.n974 585
R952 B.n974 B.n973 585
R953 B.n32 B.n31 585
R954 B.n972 B.n32 585
R955 B.n970 B.n969 585
R956 B.n971 B.n970 585
R957 B.n968 B.n37 585
R958 B.n37 B.n36 585
R959 B.n967 B.n966 585
R960 B.n966 B.n965 585
R961 B.n39 B.n38 585
R962 B.n964 B.n39 585
R963 B.n962 B.n961 585
R964 B.n963 B.n962 585
R965 B.n960 B.n44 585
R966 B.n44 B.n43 585
R967 B.n959 B.n958 585
R968 B.n958 B.n957 585
R969 B.n46 B.n45 585
R970 B.n956 B.n46 585
R971 B.n954 B.n953 585
R972 B.n955 B.n954 585
R973 B.n952 B.n51 585
R974 B.n51 B.n50 585
R975 B.n951 B.n950 585
R976 B.n950 B.n949 585
R977 B.n53 B.n52 585
R978 B.n948 B.n53 585
R979 B.n946 B.n945 585
R980 B.n947 B.n946 585
R981 B.n944 B.n57 585
R982 B.n60 B.n57 585
R983 B.n943 B.n942 585
R984 B.n942 B.n941 585
R985 B.n59 B.n58 585
R986 B.n940 B.n59 585
R987 B.n938 B.n937 585
R988 B.n939 B.n938 585
R989 B.n936 B.n65 585
R990 B.n65 B.n64 585
R991 B.n935 B.n934 585
R992 B.n934 B.n933 585
R993 B.n67 B.n66 585
R994 B.n932 B.n67 585
R995 B.n930 B.n929 585
R996 B.n931 B.n930 585
R997 B.n928 B.n72 585
R998 B.n72 B.n71 585
R999 B.n927 B.n926 585
R1000 B.n926 B.n925 585
R1001 B.n74 B.n73 585
R1002 B.n924 B.n74 585
R1003 B.n922 B.n921 585
R1004 B.n923 B.n922 585
R1005 B.n920 B.n78 585
R1006 B.n81 B.n78 585
R1007 B.n919 B.n918 585
R1008 B.n918 B.n917 585
R1009 B.n80 B.n79 585
R1010 B.n916 B.n80 585
R1011 B.n914 B.n913 585
R1012 B.n915 B.n914 585
R1013 B.n912 B.n86 585
R1014 B.n86 B.n85 585
R1015 B.n911 B.n910 585
R1016 B.n910 B.n909 585
R1017 B.n88 B.n87 585
R1018 B.n908 B.n88 585
R1019 B.n906 B.n905 585
R1020 B.n907 B.n906 585
R1021 B.n904 B.n93 585
R1022 B.n93 B.n92 585
R1023 B.n903 B.n902 585
R1024 B.n902 B.n901 585
R1025 B.n95 B.n94 585
R1026 B.n900 B.n95 585
R1027 B.n898 B.n897 585
R1028 B.n899 B.n898 585
R1029 B.n896 B.n99 585
R1030 B.n102 B.n99 585
R1031 B.n895 B.n894 585
R1032 B.n894 B.n893 585
R1033 B.n101 B.n100 585
R1034 B.n892 B.n101 585
R1035 B.n890 B.n889 585
R1036 B.n891 B.n890 585
R1037 B.n888 B.n107 585
R1038 B.n107 B.n106 585
R1039 B.n887 B.n886 585
R1040 B.n886 B.n885 585
R1041 B.n109 B.n108 585
R1042 B.n884 B.n109 585
R1043 B.n882 B.n881 585
R1044 B.n883 B.n882 585
R1045 B.n880 B.n114 585
R1046 B.n114 B.n113 585
R1047 B.n879 B.n878 585
R1048 B.n878 B.n877 585
R1049 B.n116 B.n115 585
R1050 B.n876 B.n116 585
R1051 B.n874 B.n873 585
R1052 B.n875 B.n874 585
R1053 B.n872 B.n121 585
R1054 B.n121 B.n120 585
R1055 B.n871 B.n870 585
R1056 B.n870 B.n869 585
R1057 B.n123 B.n122 585
R1058 B.n868 B.n123 585
R1059 B.n866 B.n865 585
R1060 B.n867 B.n866 585
R1061 B.n864 B.n128 585
R1062 B.n128 B.n127 585
R1063 B.n863 B.n862 585
R1064 B.n862 B.n861 585
R1065 B.n130 B.n129 585
R1066 B.n860 B.n130 585
R1067 B.n858 B.n857 585
R1068 B.n859 B.n858 585
R1069 B.n856 B.n135 585
R1070 B.n135 B.n134 585
R1071 B.n855 B.n854 585
R1072 B.n854 B.n853 585
R1073 B.n137 B.n136 585
R1074 B.n852 B.n137 585
R1075 B.n850 B.n849 585
R1076 B.n851 B.n850 585
R1077 B.n1007 B.n1006 585
R1078 B.n1006 B.n1005 585
R1079 B.n429 B.n320 535.745
R1080 B.n850 B.n142 535.745
R1081 B.n431 B.n318 535.745
R1082 B.n765 B.n140 535.745
R1083 B.n766 B.n141 256.663
R1084 B.n768 B.n141 256.663
R1085 B.n774 B.n141 256.663
R1086 B.n776 B.n141 256.663
R1087 B.n782 B.n141 256.663
R1088 B.n784 B.n141 256.663
R1089 B.n790 B.n141 256.663
R1090 B.n160 B.n141 256.663
R1091 B.n796 B.n141 256.663
R1092 B.n802 B.n141 256.663
R1093 B.n804 B.n141 256.663
R1094 B.n810 B.n141 256.663
R1095 B.n812 B.n141 256.663
R1096 B.n819 B.n141 256.663
R1097 B.n821 B.n141 256.663
R1098 B.n827 B.n141 256.663
R1099 B.n829 B.n141 256.663
R1100 B.n835 B.n141 256.663
R1101 B.n837 B.n141 256.663
R1102 B.n843 B.n141 256.663
R1103 B.n845 B.n141 256.663
R1104 B.n424 B.n319 256.663
R1105 B.n322 B.n319 256.663
R1106 B.n417 B.n319 256.663
R1107 B.n411 B.n319 256.663
R1108 B.n409 B.n319 256.663
R1109 B.n403 B.n319 256.663
R1110 B.n401 B.n319 256.663
R1111 B.n394 B.n319 256.663
R1112 B.n392 B.n319 256.663
R1113 B.n386 B.n319 256.663
R1114 B.n384 B.n319 256.663
R1115 B.n378 B.n319 256.663
R1116 B.n376 B.n319 256.663
R1117 B.n370 B.n319 256.663
R1118 B.n368 B.n319 256.663
R1119 B.n362 B.n319 256.663
R1120 B.n360 B.n319 256.663
R1121 B.n354 B.n319 256.663
R1122 B.n352 B.n319 256.663
R1123 B.n346 B.n319 256.663
R1124 B.n337 B.t10 231.594
R1125 B.n329 B.t21 231.594
R1126 B.n151 B.t18 231.594
R1127 B.n157 B.t14 231.594
R1128 B.n337 B.t13 212.665
R1129 B.n157 B.t16 212.665
R1130 B.n329 B.t23 212.665
R1131 B.n151 B.t19 212.665
R1132 B.n430 B.n319 171.577
R1133 B.n851 B.n141 171.577
R1134 B.n429 B.n314 163.367
R1135 B.n437 B.n314 163.367
R1136 B.n437 B.n312 163.367
R1137 B.n441 B.n312 163.367
R1138 B.n441 B.n306 163.367
R1139 B.n449 B.n306 163.367
R1140 B.n449 B.n304 163.367
R1141 B.n453 B.n304 163.367
R1142 B.n453 B.n298 163.367
R1143 B.n461 B.n298 163.367
R1144 B.n461 B.n296 163.367
R1145 B.n465 B.n296 163.367
R1146 B.n465 B.n290 163.367
R1147 B.n473 B.n290 163.367
R1148 B.n473 B.n288 163.367
R1149 B.n477 B.n288 163.367
R1150 B.n477 B.n282 163.367
R1151 B.n485 B.n282 163.367
R1152 B.n485 B.n280 163.367
R1153 B.n489 B.n280 163.367
R1154 B.n489 B.n274 163.367
R1155 B.n498 B.n274 163.367
R1156 B.n498 B.n272 163.367
R1157 B.n502 B.n272 163.367
R1158 B.n502 B.n267 163.367
R1159 B.n510 B.n267 163.367
R1160 B.n510 B.n265 163.367
R1161 B.n514 B.n265 163.367
R1162 B.n514 B.n259 163.367
R1163 B.n522 B.n259 163.367
R1164 B.n522 B.n257 163.367
R1165 B.n526 B.n257 163.367
R1166 B.n526 B.n251 163.367
R1167 B.n535 B.n251 163.367
R1168 B.n535 B.n249 163.367
R1169 B.n539 B.n249 163.367
R1170 B.n539 B.n244 163.367
R1171 B.n547 B.n244 163.367
R1172 B.n547 B.n242 163.367
R1173 B.n551 B.n242 163.367
R1174 B.n551 B.n236 163.367
R1175 B.n559 B.n236 163.367
R1176 B.n559 B.n234 163.367
R1177 B.n563 B.n234 163.367
R1178 B.n563 B.n228 163.367
R1179 B.n572 B.n228 163.367
R1180 B.n572 B.n226 163.367
R1181 B.n576 B.n226 163.367
R1182 B.n576 B.n221 163.367
R1183 B.n584 B.n221 163.367
R1184 B.n584 B.n219 163.367
R1185 B.n588 B.n219 163.367
R1186 B.n588 B.n213 163.367
R1187 B.n596 B.n213 163.367
R1188 B.n596 B.n211 163.367
R1189 B.n600 B.n211 163.367
R1190 B.n600 B.n205 163.367
R1191 B.n608 B.n205 163.367
R1192 B.n608 B.n203 163.367
R1193 B.n612 B.n203 163.367
R1194 B.n612 B.n197 163.367
R1195 B.n620 B.n197 163.367
R1196 B.n620 B.n195 163.367
R1197 B.n624 B.n195 163.367
R1198 B.n624 B.n189 163.367
R1199 B.n632 B.n189 163.367
R1200 B.n632 B.n187 163.367
R1201 B.n636 B.n187 163.367
R1202 B.n636 B.n181 163.367
R1203 B.n644 B.n181 163.367
R1204 B.n644 B.n179 163.367
R1205 B.n648 B.n179 163.367
R1206 B.n648 B.n173 163.367
R1207 B.n657 B.n173 163.367
R1208 B.n657 B.n171 163.367
R1209 B.n661 B.n171 163.367
R1210 B.n661 B.n2 163.367
R1211 B.n1006 B.n2 163.367
R1212 B.n1006 B.n3 163.367
R1213 B.n1002 B.n3 163.367
R1214 B.n1002 B.n9 163.367
R1215 B.n998 B.n9 163.367
R1216 B.n998 B.n11 163.367
R1217 B.n994 B.n11 163.367
R1218 B.n994 B.n16 163.367
R1219 B.n990 B.n16 163.367
R1220 B.n990 B.n18 163.367
R1221 B.n986 B.n18 163.367
R1222 B.n986 B.n23 163.367
R1223 B.n982 B.n23 163.367
R1224 B.n982 B.n25 163.367
R1225 B.n978 B.n25 163.367
R1226 B.n978 B.n30 163.367
R1227 B.n974 B.n30 163.367
R1228 B.n974 B.n32 163.367
R1229 B.n970 B.n32 163.367
R1230 B.n970 B.n37 163.367
R1231 B.n966 B.n37 163.367
R1232 B.n966 B.n39 163.367
R1233 B.n962 B.n39 163.367
R1234 B.n962 B.n44 163.367
R1235 B.n958 B.n44 163.367
R1236 B.n958 B.n46 163.367
R1237 B.n954 B.n46 163.367
R1238 B.n954 B.n51 163.367
R1239 B.n950 B.n51 163.367
R1240 B.n950 B.n53 163.367
R1241 B.n946 B.n53 163.367
R1242 B.n946 B.n57 163.367
R1243 B.n942 B.n57 163.367
R1244 B.n942 B.n59 163.367
R1245 B.n938 B.n59 163.367
R1246 B.n938 B.n65 163.367
R1247 B.n934 B.n65 163.367
R1248 B.n934 B.n67 163.367
R1249 B.n930 B.n67 163.367
R1250 B.n930 B.n72 163.367
R1251 B.n926 B.n72 163.367
R1252 B.n926 B.n74 163.367
R1253 B.n922 B.n74 163.367
R1254 B.n922 B.n78 163.367
R1255 B.n918 B.n78 163.367
R1256 B.n918 B.n80 163.367
R1257 B.n914 B.n80 163.367
R1258 B.n914 B.n86 163.367
R1259 B.n910 B.n86 163.367
R1260 B.n910 B.n88 163.367
R1261 B.n906 B.n88 163.367
R1262 B.n906 B.n93 163.367
R1263 B.n902 B.n93 163.367
R1264 B.n902 B.n95 163.367
R1265 B.n898 B.n95 163.367
R1266 B.n898 B.n99 163.367
R1267 B.n894 B.n99 163.367
R1268 B.n894 B.n101 163.367
R1269 B.n890 B.n101 163.367
R1270 B.n890 B.n107 163.367
R1271 B.n886 B.n107 163.367
R1272 B.n886 B.n109 163.367
R1273 B.n882 B.n109 163.367
R1274 B.n882 B.n114 163.367
R1275 B.n878 B.n114 163.367
R1276 B.n878 B.n116 163.367
R1277 B.n874 B.n116 163.367
R1278 B.n874 B.n121 163.367
R1279 B.n870 B.n121 163.367
R1280 B.n870 B.n123 163.367
R1281 B.n866 B.n123 163.367
R1282 B.n866 B.n128 163.367
R1283 B.n862 B.n128 163.367
R1284 B.n862 B.n130 163.367
R1285 B.n858 B.n130 163.367
R1286 B.n858 B.n135 163.367
R1287 B.n854 B.n135 163.367
R1288 B.n854 B.n137 163.367
R1289 B.n850 B.n137 163.367
R1290 B.n425 B.n423 163.367
R1291 B.n423 B.n422 163.367
R1292 B.n419 B.n418 163.367
R1293 B.n416 B.n324 163.367
R1294 B.n412 B.n410 163.367
R1295 B.n408 B.n326 163.367
R1296 B.n404 B.n402 163.367
R1297 B.n400 B.n328 163.367
R1298 B.n395 B.n393 163.367
R1299 B.n391 B.n332 163.367
R1300 B.n387 B.n385 163.367
R1301 B.n383 B.n334 163.367
R1302 B.n379 B.n377 163.367
R1303 B.n375 B.n336 163.367
R1304 B.n371 B.n369 163.367
R1305 B.n367 B.n341 163.367
R1306 B.n363 B.n361 163.367
R1307 B.n359 B.n343 163.367
R1308 B.n355 B.n353 163.367
R1309 B.n351 B.n345 163.367
R1310 B.n347 B.n318 163.367
R1311 B.n431 B.n316 163.367
R1312 B.n435 B.n316 163.367
R1313 B.n435 B.n310 163.367
R1314 B.n443 B.n310 163.367
R1315 B.n443 B.n308 163.367
R1316 B.n447 B.n308 163.367
R1317 B.n447 B.n302 163.367
R1318 B.n455 B.n302 163.367
R1319 B.n455 B.n300 163.367
R1320 B.n459 B.n300 163.367
R1321 B.n459 B.n294 163.367
R1322 B.n467 B.n294 163.367
R1323 B.n467 B.n292 163.367
R1324 B.n471 B.n292 163.367
R1325 B.n471 B.n286 163.367
R1326 B.n479 B.n286 163.367
R1327 B.n479 B.n284 163.367
R1328 B.n483 B.n284 163.367
R1329 B.n483 B.n278 163.367
R1330 B.n491 B.n278 163.367
R1331 B.n491 B.n276 163.367
R1332 B.n495 B.n276 163.367
R1333 B.n495 B.n271 163.367
R1334 B.n504 B.n271 163.367
R1335 B.n504 B.n269 163.367
R1336 B.n508 B.n269 163.367
R1337 B.n508 B.n263 163.367
R1338 B.n516 B.n263 163.367
R1339 B.n516 B.n261 163.367
R1340 B.n520 B.n261 163.367
R1341 B.n520 B.n255 163.367
R1342 B.n528 B.n255 163.367
R1343 B.n528 B.n253 163.367
R1344 B.n532 B.n253 163.367
R1345 B.n532 B.n248 163.367
R1346 B.n541 B.n248 163.367
R1347 B.n541 B.n246 163.367
R1348 B.n545 B.n246 163.367
R1349 B.n545 B.n240 163.367
R1350 B.n553 B.n240 163.367
R1351 B.n553 B.n238 163.367
R1352 B.n557 B.n238 163.367
R1353 B.n557 B.n232 163.367
R1354 B.n565 B.n232 163.367
R1355 B.n565 B.n230 163.367
R1356 B.n569 B.n230 163.367
R1357 B.n569 B.n225 163.367
R1358 B.n578 B.n225 163.367
R1359 B.n578 B.n223 163.367
R1360 B.n582 B.n223 163.367
R1361 B.n582 B.n217 163.367
R1362 B.n590 B.n217 163.367
R1363 B.n590 B.n215 163.367
R1364 B.n594 B.n215 163.367
R1365 B.n594 B.n209 163.367
R1366 B.n602 B.n209 163.367
R1367 B.n602 B.n207 163.367
R1368 B.n606 B.n207 163.367
R1369 B.n606 B.n201 163.367
R1370 B.n614 B.n201 163.367
R1371 B.n614 B.n199 163.367
R1372 B.n618 B.n199 163.367
R1373 B.n618 B.n193 163.367
R1374 B.n626 B.n193 163.367
R1375 B.n626 B.n191 163.367
R1376 B.n630 B.n191 163.367
R1377 B.n630 B.n185 163.367
R1378 B.n638 B.n185 163.367
R1379 B.n638 B.n183 163.367
R1380 B.n642 B.n183 163.367
R1381 B.n642 B.n177 163.367
R1382 B.n650 B.n177 163.367
R1383 B.n650 B.n175 163.367
R1384 B.n655 B.n175 163.367
R1385 B.n655 B.n169 163.367
R1386 B.n663 B.n169 163.367
R1387 B.n664 B.n663 163.367
R1388 B.n664 B.n5 163.367
R1389 B.n6 B.n5 163.367
R1390 B.n7 B.n6 163.367
R1391 B.n669 B.n7 163.367
R1392 B.n669 B.n12 163.367
R1393 B.n13 B.n12 163.367
R1394 B.n14 B.n13 163.367
R1395 B.n674 B.n14 163.367
R1396 B.n674 B.n19 163.367
R1397 B.n20 B.n19 163.367
R1398 B.n21 B.n20 163.367
R1399 B.n679 B.n21 163.367
R1400 B.n679 B.n26 163.367
R1401 B.n27 B.n26 163.367
R1402 B.n28 B.n27 163.367
R1403 B.n684 B.n28 163.367
R1404 B.n684 B.n33 163.367
R1405 B.n34 B.n33 163.367
R1406 B.n35 B.n34 163.367
R1407 B.n689 B.n35 163.367
R1408 B.n689 B.n40 163.367
R1409 B.n41 B.n40 163.367
R1410 B.n42 B.n41 163.367
R1411 B.n694 B.n42 163.367
R1412 B.n694 B.n47 163.367
R1413 B.n48 B.n47 163.367
R1414 B.n49 B.n48 163.367
R1415 B.n699 B.n49 163.367
R1416 B.n699 B.n54 163.367
R1417 B.n55 B.n54 163.367
R1418 B.n56 B.n55 163.367
R1419 B.n704 B.n56 163.367
R1420 B.n704 B.n61 163.367
R1421 B.n62 B.n61 163.367
R1422 B.n63 B.n62 163.367
R1423 B.n709 B.n63 163.367
R1424 B.n709 B.n68 163.367
R1425 B.n69 B.n68 163.367
R1426 B.n70 B.n69 163.367
R1427 B.n714 B.n70 163.367
R1428 B.n714 B.n75 163.367
R1429 B.n76 B.n75 163.367
R1430 B.n77 B.n76 163.367
R1431 B.n719 B.n77 163.367
R1432 B.n719 B.n82 163.367
R1433 B.n83 B.n82 163.367
R1434 B.n84 B.n83 163.367
R1435 B.n724 B.n84 163.367
R1436 B.n724 B.n89 163.367
R1437 B.n90 B.n89 163.367
R1438 B.n91 B.n90 163.367
R1439 B.n729 B.n91 163.367
R1440 B.n729 B.n96 163.367
R1441 B.n97 B.n96 163.367
R1442 B.n98 B.n97 163.367
R1443 B.n734 B.n98 163.367
R1444 B.n734 B.n103 163.367
R1445 B.n104 B.n103 163.367
R1446 B.n105 B.n104 163.367
R1447 B.n739 B.n105 163.367
R1448 B.n739 B.n110 163.367
R1449 B.n111 B.n110 163.367
R1450 B.n112 B.n111 163.367
R1451 B.n744 B.n112 163.367
R1452 B.n744 B.n117 163.367
R1453 B.n118 B.n117 163.367
R1454 B.n119 B.n118 163.367
R1455 B.n749 B.n119 163.367
R1456 B.n749 B.n124 163.367
R1457 B.n125 B.n124 163.367
R1458 B.n126 B.n125 163.367
R1459 B.n754 B.n126 163.367
R1460 B.n754 B.n131 163.367
R1461 B.n132 B.n131 163.367
R1462 B.n133 B.n132 163.367
R1463 B.n759 B.n133 163.367
R1464 B.n759 B.n138 163.367
R1465 B.n139 B.n138 163.367
R1466 B.n140 B.n139 163.367
R1467 B.n846 B.n844 163.367
R1468 B.n842 B.n144 163.367
R1469 B.n838 B.n836 163.367
R1470 B.n834 B.n146 163.367
R1471 B.n830 B.n828 163.367
R1472 B.n826 B.n148 163.367
R1473 B.n822 B.n820 163.367
R1474 B.n818 B.n150 163.367
R1475 B.n813 B.n811 163.367
R1476 B.n809 B.n154 163.367
R1477 B.n805 B.n803 163.367
R1478 B.n801 B.n156 163.367
R1479 B.n797 B.n795 163.367
R1480 B.n792 B.n791 163.367
R1481 B.n789 B.n162 163.367
R1482 B.n785 B.n783 163.367
R1483 B.n781 B.n164 163.367
R1484 B.n777 B.n775 163.367
R1485 B.n773 B.n166 163.367
R1486 B.n769 B.n767 163.367
R1487 B.n338 B.t12 135.671
R1488 B.n158 B.t17 135.671
R1489 B.n330 B.t22 135.671
R1490 B.n152 B.t20 135.671
R1491 B.n430 B.n315 86.4245
R1492 B.n436 B.n315 86.4245
R1493 B.n436 B.n311 86.4245
R1494 B.n442 B.n311 86.4245
R1495 B.n442 B.n307 86.4245
R1496 B.n448 B.n307 86.4245
R1497 B.n448 B.n303 86.4245
R1498 B.n454 B.n303 86.4245
R1499 B.n460 B.n299 86.4245
R1500 B.n460 B.n295 86.4245
R1501 B.n466 B.n295 86.4245
R1502 B.n466 B.n291 86.4245
R1503 B.n472 B.n291 86.4245
R1504 B.n472 B.n287 86.4245
R1505 B.n478 B.n287 86.4245
R1506 B.n478 B.n283 86.4245
R1507 B.n484 B.n283 86.4245
R1508 B.n484 B.n279 86.4245
R1509 B.n490 B.n279 86.4245
R1510 B.n490 B.n275 86.4245
R1511 B.n497 B.n275 86.4245
R1512 B.n497 B.n496 86.4245
R1513 B.n503 B.n268 86.4245
R1514 B.n509 B.n268 86.4245
R1515 B.n509 B.n264 86.4245
R1516 B.n515 B.n264 86.4245
R1517 B.n515 B.n260 86.4245
R1518 B.n521 B.n260 86.4245
R1519 B.n521 B.n256 86.4245
R1520 B.n527 B.n256 86.4245
R1521 B.n527 B.n252 86.4245
R1522 B.n534 B.n252 86.4245
R1523 B.n534 B.n533 86.4245
R1524 B.n540 B.n245 86.4245
R1525 B.n546 B.n245 86.4245
R1526 B.n546 B.n241 86.4245
R1527 B.n552 B.n241 86.4245
R1528 B.n552 B.n237 86.4245
R1529 B.n558 B.n237 86.4245
R1530 B.n558 B.n233 86.4245
R1531 B.n564 B.n233 86.4245
R1532 B.n564 B.n229 86.4245
R1533 B.n571 B.n229 86.4245
R1534 B.n571 B.n570 86.4245
R1535 B.n577 B.n222 86.4245
R1536 B.n583 B.n222 86.4245
R1537 B.n583 B.n218 86.4245
R1538 B.n589 B.n218 86.4245
R1539 B.n589 B.n214 86.4245
R1540 B.n595 B.n214 86.4245
R1541 B.n595 B.n210 86.4245
R1542 B.n601 B.n210 86.4245
R1543 B.n601 B.n206 86.4245
R1544 B.n607 B.n206 86.4245
R1545 B.n613 B.n202 86.4245
R1546 B.n613 B.n198 86.4245
R1547 B.n619 B.n198 86.4245
R1548 B.n619 B.n194 86.4245
R1549 B.n625 B.n194 86.4245
R1550 B.n625 B.n190 86.4245
R1551 B.n631 B.n190 86.4245
R1552 B.n631 B.n186 86.4245
R1553 B.n637 B.n186 86.4245
R1554 B.n637 B.n182 86.4245
R1555 B.n643 B.n182 86.4245
R1556 B.n649 B.n178 86.4245
R1557 B.n649 B.n174 86.4245
R1558 B.n656 B.n174 86.4245
R1559 B.n656 B.n170 86.4245
R1560 B.n662 B.n170 86.4245
R1561 B.n662 B.n4 86.4245
R1562 B.n1005 B.n4 86.4245
R1563 B.n1005 B.n1004 86.4245
R1564 B.n1004 B.n1003 86.4245
R1565 B.n1003 B.n8 86.4245
R1566 B.n997 B.n8 86.4245
R1567 B.n997 B.n996 86.4245
R1568 B.n996 B.n995 86.4245
R1569 B.n995 B.n15 86.4245
R1570 B.n989 B.n988 86.4245
R1571 B.n988 B.n987 86.4245
R1572 B.n987 B.n22 86.4245
R1573 B.n981 B.n22 86.4245
R1574 B.n981 B.n980 86.4245
R1575 B.n980 B.n979 86.4245
R1576 B.n979 B.n29 86.4245
R1577 B.n973 B.n29 86.4245
R1578 B.n973 B.n972 86.4245
R1579 B.n972 B.n971 86.4245
R1580 B.n971 B.n36 86.4245
R1581 B.n965 B.n964 86.4245
R1582 B.n964 B.n963 86.4245
R1583 B.n963 B.n43 86.4245
R1584 B.n957 B.n43 86.4245
R1585 B.n957 B.n956 86.4245
R1586 B.n956 B.n955 86.4245
R1587 B.n955 B.n50 86.4245
R1588 B.n949 B.n50 86.4245
R1589 B.n949 B.n948 86.4245
R1590 B.n948 B.n947 86.4245
R1591 B.n941 B.n60 86.4245
R1592 B.n941 B.n940 86.4245
R1593 B.n940 B.n939 86.4245
R1594 B.n939 B.n64 86.4245
R1595 B.n933 B.n64 86.4245
R1596 B.n933 B.n932 86.4245
R1597 B.n932 B.n931 86.4245
R1598 B.n931 B.n71 86.4245
R1599 B.n925 B.n71 86.4245
R1600 B.n925 B.n924 86.4245
R1601 B.n924 B.n923 86.4245
R1602 B.n917 B.n81 86.4245
R1603 B.n917 B.n916 86.4245
R1604 B.n916 B.n915 86.4245
R1605 B.n915 B.n85 86.4245
R1606 B.n909 B.n85 86.4245
R1607 B.n909 B.n908 86.4245
R1608 B.n908 B.n907 86.4245
R1609 B.n907 B.n92 86.4245
R1610 B.n901 B.n92 86.4245
R1611 B.n901 B.n900 86.4245
R1612 B.n900 B.n899 86.4245
R1613 B.n893 B.n102 86.4245
R1614 B.n893 B.n892 86.4245
R1615 B.n892 B.n891 86.4245
R1616 B.n891 B.n106 86.4245
R1617 B.n885 B.n106 86.4245
R1618 B.n885 B.n884 86.4245
R1619 B.n884 B.n883 86.4245
R1620 B.n883 B.n113 86.4245
R1621 B.n877 B.n113 86.4245
R1622 B.n877 B.n876 86.4245
R1623 B.n876 B.n875 86.4245
R1624 B.n875 B.n120 86.4245
R1625 B.n869 B.n120 86.4245
R1626 B.n869 B.n868 86.4245
R1627 B.n867 B.n127 86.4245
R1628 B.n861 B.n127 86.4245
R1629 B.n861 B.n860 86.4245
R1630 B.n860 B.n859 86.4245
R1631 B.n859 B.n134 86.4245
R1632 B.n853 B.n134 86.4245
R1633 B.n853 B.n852 86.4245
R1634 B.n852 B.n851 86.4245
R1635 B.n454 B.t11 83.8826
R1636 B.t15 B.n867 83.8826
R1637 B.n338 B.n337 76.9944
R1638 B.n330 B.n329 76.9944
R1639 B.n152 B.n151 76.9944
R1640 B.n158 B.n157 76.9944
R1641 B.n607 B.t6 76.257
R1642 B.n965 B.t1 76.257
R1643 B.n496 B.t5 73.7151
R1644 B.n102 B.t3 73.7151
R1645 B.n424 B.n320 71.676
R1646 B.n422 B.n322 71.676
R1647 B.n418 B.n417 71.676
R1648 B.n411 B.n324 71.676
R1649 B.n410 B.n409 71.676
R1650 B.n403 B.n326 71.676
R1651 B.n402 B.n401 71.676
R1652 B.n394 B.n328 71.676
R1653 B.n393 B.n392 71.676
R1654 B.n386 B.n332 71.676
R1655 B.n385 B.n384 71.676
R1656 B.n378 B.n334 71.676
R1657 B.n377 B.n376 71.676
R1658 B.n370 B.n336 71.676
R1659 B.n369 B.n368 71.676
R1660 B.n362 B.n341 71.676
R1661 B.n361 B.n360 71.676
R1662 B.n354 B.n343 71.676
R1663 B.n353 B.n352 71.676
R1664 B.n346 B.n345 71.676
R1665 B.n845 B.n142 71.676
R1666 B.n844 B.n843 71.676
R1667 B.n837 B.n144 71.676
R1668 B.n836 B.n835 71.676
R1669 B.n829 B.n146 71.676
R1670 B.n828 B.n827 71.676
R1671 B.n821 B.n148 71.676
R1672 B.n820 B.n819 71.676
R1673 B.n812 B.n150 71.676
R1674 B.n811 B.n810 71.676
R1675 B.n804 B.n154 71.676
R1676 B.n803 B.n802 71.676
R1677 B.n796 B.n156 71.676
R1678 B.n795 B.n160 71.676
R1679 B.n791 B.n790 71.676
R1680 B.n784 B.n162 71.676
R1681 B.n783 B.n782 71.676
R1682 B.n776 B.n164 71.676
R1683 B.n775 B.n774 71.676
R1684 B.n768 B.n166 71.676
R1685 B.n767 B.n766 71.676
R1686 B.n766 B.n765 71.676
R1687 B.n769 B.n768 71.676
R1688 B.n774 B.n773 71.676
R1689 B.n777 B.n776 71.676
R1690 B.n782 B.n781 71.676
R1691 B.n785 B.n784 71.676
R1692 B.n790 B.n789 71.676
R1693 B.n792 B.n160 71.676
R1694 B.n797 B.n796 71.676
R1695 B.n802 B.n801 71.676
R1696 B.n805 B.n804 71.676
R1697 B.n810 B.n809 71.676
R1698 B.n813 B.n812 71.676
R1699 B.n819 B.n818 71.676
R1700 B.n822 B.n821 71.676
R1701 B.n827 B.n826 71.676
R1702 B.n830 B.n829 71.676
R1703 B.n835 B.n834 71.676
R1704 B.n838 B.n837 71.676
R1705 B.n843 B.n842 71.676
R1706 B.n846 B.n845 71.676
R1707 B.n425 B.n424 71.676
R1708 B.n419 B.n322 71.676
R1709 B.n417 B.n416 71.676
R1710 B.n412 B.n411 71.676
R1711 B.n409 B.n408 71.676
R1712 B.n404 B.n403 71.676
R1713 B.n401 B.n400 71.676
R1714 B.n395 B.n394 71.676
R1715 B.n392 B.n391 71.676
R1716 B.n387 B.n386 71.676
R1717 B.n384 B.n383 71.676
R1718 B.n379 B.n378 71.676
R1719 B.n376 B.n375 71.676
R1720 B.n371 B.n370 71.676
R1721 B.n368 B.n367 71.676
R1722 B.n363 B.n362 71.676
R1723 B.n360 B.n359 71.676
R1724 B.n355 B.n354 71.676
R1725 B.n352 B.n351 71.676
R1726 B.n347 B.n346 71.676
R1727 B.n577 B.t4 68.6314
R1728 B.n947 B.t9 68.6314
R1729 B.n339 B.n338 59.5399
R1730 B.n397 B.n330 59.5399
R1731 B.n816 B.n152 59.5399
R1732 B.n159 B.n158 59.5399
R1733 B.n643 B.t8 48.2963
R1734 B.n989 B.t2 48.2963
R1735 B.n533 B.t0 45.7544
R1736 B.n81 B.t7 45.7544
R1737 B.n540 B.t0 40.6706
R1738 B.n923 B.t7 40.6706
R1739 B.t8 B.n178 38.1288
R1740 B.t2 B.n15 38.1288
R1741 B.n764 B.n763 34.8103
R1742 B.n849 B.n848 34.8103
R1743 B.n432 B.n317 34.8103
R1744 B.n428 B.n427 34.8103
R1745 B B.n1007 18.0485
R1746 B.n570 B.t4 17.7937
R1747 B.n60 B.t9 17.7937
R1748 B.n503 B.t5 12.7099
R1749 B.n899 B.t3 12.7099
R1750 B.n848 B.n847 10.6151
R1751 B.n847 B.n143 10.6151
R1752 B.n841 B.n143 10.6151
R1753 B.n841 B.n840 10.6151
R1754 B.n840 B.n839 10.6151
R1755 B.n839 B.n145 10.6151
R1756 B.n833 B.n145 10.6151
R1757 B.n833 B.n832 10.6151
R1758 B.n832 B.n831 10.6151
R1759 B.n831 B.n147 10.6151
R1760 B.n825 B.n147 10.6151
R1761 B.n825 B.n824 10.6151
R1762 B.n824 B.n823 10.6151
R1763 B.n823 B.n149 10.6151
R1764 B.n817 B.n149 10.6151
R1765 B.n815 B.n814 10.6151
R1766 B.n814 B.n153 10.6151
R1767 B.n808 B.n153 10.6151
R1768 B.n808 B.n807 10.6151
R1769 B.n807 B.n806 10.6151
R1770 B.n806 B.n155 10.6151
R1771 B.n800 B.n155 10.6151
R1772 B.n800 B.n799 10.6151
R1773 B.n799 B.n798 10.6151
R1774 B.n794 B.n793 10.6151
R1775 B.n793 B.n161 10.6151
R1776 B.n788 B.n161 10.6151
R1777 B.n788 B.n787 10.6151
R1778 B.n787 B.n786 10.6151
R1779 B.n786 B.n163 10.6151
R1780 B.n780 B.n163 10.6151
R1781 B.n780 B.n779 10.6151
R1782 B.n779 B.n778 10.6151
R1783 B.n778 B.n165 10.6151
R1784 B.n772 B.n165 10.6151
R1785 B.n772 B.n771 10.6151
R1786 B.n771 B.n770 10.6151
R1787 B.n770 B.n167 10.6151
R1788 B.n764 B.n167 10.6151
R1789 B.n433 B.n432 10.6151
R1790 B.n434 B.n433 10.6151
R1791 B.n434 B.n309 10.6151
R1792 B.n444 B.n309 10.6151
R1793 B.n445 B.n444 10.6151
R1794 B.n446 B.n445 10.6151
R1795 B.n446 B.n301 10.6151
R1796 B.n456 B.n301 10.6151
R1797 B.n457 B.n456 10.6151
R1798 B.n458 B.n457 10.6151
R1799 B.n458 B.n293 10.6151
R1800 B.n468 B.n293 10.6151
R1801 B.n469 B.n468 10.6151
R1802 B.n470 B.n469 10.6151
R1803 B.n470 B.n285 10.6151
R1804 B.n480 B.n285 10.6151
R1805 B.n481 B.n480 10.6151
R1806 B.n482 B.n481 10.6151
R1807 B.n482 B.n277 10.6151
R1808 B.n492 B.n277 10.6151
R1809 B.n493 B.n492 10.6151
R1810 B.n494 B.n493 10.6151
R1811 B.n494 B.n270 10.6151
R1812 B.n505 B.n270 10.6151
R1813 B.n506 B.n505 10.6151
R1814 B.n507 B.n506 10.6151
R1815 B.n507 B.n262 10.6151
R1816 B.n517 B.n262 10.6151
R1817 B.n518 B.n517 10.6151
R1818 B.n519 B.n518 10.6151
R1819 B.n519 B.n254 10.6151
R1820 B.n529 B.n254 10.6151
R1821 B.n530 B.n529 10.6151
R1822 B.n531 B.n530 10.6151
R1823 B.n531 B.n247 10.6151
R1824 B.n542 B.n247 10.6151
R1825 B.n543 B.n542 10.6151
R1826 B.n544 B.n543 10.6151
R1827 B.n544 B.n239 10.6151
R1828 B.n554 B.n239 10.6151
R1829 B.n555 B.n554 10.6151
R1830 B.n556 B.n555 10.6151
R1831 B.n556 B.n231 10.6151
R1832 B.n566 B.n231 10.6151
R1833 B.n567 B.n566 10.6151
R1834 B.n568 B.n567 10.6151
R1835 B.n568 B.n224 10.6151
R1836 B.n579 B.n224 10.6151
R1837 B.n580 B.n579 10.6151
R1838 B.n581 B.n580 10.6151
R1839 B.n581 B.n216 10.6151
R1840 B.n591 B.n216 10.6151
R1841 B.n592 B.n591 10.6151
R1842 B.n593 B.n592 10.6151
R1843 B.n593 B.n208 10.6151
R1844 B.n603 B.n208 10.6151
R1845 B.n604 B.n603 10.6151
R1846 B.n605 B.n604 10.6151
R1847 B.n605 B.n200 10.6151
R1848 B.n615 B.n200 10.6151
R1849 B.n616 B.n615 10.6151
R1850 B.n617 B.n616 10.6151
R1851 B.n617 B.n192 10.6151
R1852 B.n627 B.n192 10.6151
R1853 B.n628 B.n627 10.6151
R1854 B.n629 B.n628 10.6151
R1855 B.n629 B.n184 10.6151
R1856 B.n639 B.n184 10.6151
R1857 B.n640 B.n639 10.6151
R1858 B.n641 B.n640 10.6151
R1859 B.n641 B.n176 10.6151
R1860 B.n651 B.n176 10.6151
R1861 B.n652 B.n651 10.6151
R1862 B.n654 B.n652 10.6151
R1863 B.n654 B.n653 10.6151
R1864 B.n653 B.n168 10.6151
R1865 B.n665 B.n168 10.6151
R1866 B.n666 B.n665 10.6151
R1867 B.n667 B.n666 10.6151
R1868 B.n668 B.n667 10.6151
R1869 B.n670 B.n668 10.6151
R1870 B.n671 B.n670 10.6151
R1871 B.n672 B.n671 10.6151
R1872 B.n673 B.n672 10.6151
R1873 B.n675 B.n673 10.6151
R1874 B.n676 B.n675 10.6151
R1875 B.n677 B.n676 10.6151
R1876 B.n678 B.n677 10.6151
R1877 B.n680 B.n678 10.6151
R1878 B.n681 B.n680 10.6151
R1879 B.n682 B.n681 10.6151
R1880 B.n683 B.n682 10.6151
R1881 B.n685 B.n683 10.6151
R1882 B.n686 B.n685 10.6151
R1883 B.n687 B.n686 10.6151
R1884 B.n688 B.n687 10.6151
R1885 B.n690 B.n688 10.6151
R1886 B.n691 B.n690 10.6151
R1887 B.n692 B.n691 10.6151
R1888 B.n693 B.n692 10.6151
R1889 B.n695 B.n693 10.6151
R1890 B.n696 B.n695 10.6151
R1891 B.n697 B.n696 10.6151
R1892 B.n698 B.n697 10.6151
R1893 B.n700 B.n698 10.6151
R1894 B.n701 B.n700 10.6151
R1895 B.n702 B.n701 10.6151
R1896 B.n703 B.n702 10.6151
R1897 B.n705 B.n703 10.6151
R1898 B.n706 B.n705 10.6151
R1899 B.n707 B.n706 10.6151
R1900 B.n708 B.n707 10.6151
R1901 B.n710 B.n708 10.6151
R1902 B.n711 B.n710 10.6151
R1903 B.n712 B.n711 10.6151
R1904 B.n713 B.n712 10.6151
R1905 B.n715 B.n713 10.6151
R1906 B.n716 B.n715 10.6151
R1907 B.n717 B.n716 10.6151
R1908 B.n718 B.n717 10.6151
R1909 B.n720 B.n718 10.6151
R1910 B.n721 B.n720 10.6151
R1911 B.n722 B.n721 10.6151
R1912 B.n723 B.n722 10.6151
R1913 B.n725 B.n723 10.6151
R1914 B.n726 B.n725 10.6151
R1915 B.n727 B.n726 10.6151
R1916 B.n728 B.n727 10.6151
R1917 B.n730 B.n728 10.6151
R1918 B.n731 B.n730 10.6151
R1919 B.n732 B.n731 10.6151
R1920 B.n733 B.n732 10.6151
R1921 B.n735 B.n733 10.6151
R1922 B.n736 B.n735 10.6151
R1923 B.n737 B.n736 10.6151
R1924 B.n738 B.n737 10.6151
R1925 B.n740 B.n738 10.6151
R1926 B.n741 B.n740 10.6151
R1927 B.n742 B.n741 10.6151
R1928 B.n743 B.n742 10.6151
R1929 B.n745 B.n743 10.6151
R1930 B.n746 B.n745 10.6151
R1931 B.n747 B.n746 10.6151
R1932 B.n748 B.n747 10.6151
R1933 B.n750 B.n748 10.6151
R1934 B.n751 B.n750 10.6151
R1935 B.n752 B.n751 10.6151
R1936 B.n753 B.n752 10.6151
R1937 B.n755 B.n753 10.6151
R1938 B.n756 B.n755 10.6151
R1939 B.n757 B.n756 10.6151
R1940 B.n758 B.n757 10.6151
R1941 B.n760 B.n758 10.6151
R1942 B.n761 B.n760 10.6151
R1943 B.n762 B.n761 10.6151
R1944 B.n763 B.n762 10.6151
R1945 B.n427 B.n426 10.6151
R1946 B.n426 B.n321 10.6151
R1947 B.n421 B.n321 10.6151
R1948 B.n421 B.n420 10.6151
R1949 B.n420 B.n323 10.6151
R1950 B.n415 B.n323 10.6151
R1951 B.n415 B.n414 10.6151
R1952 B.n414 B.n413 10.6151
R1953 B.n413 B.n325 10.6151
R1954 B.n407 B.n325 10.6151
R1955 B.n407 B.n406 10.6151
R1956 B.n406 B.n405 10.6151
R1957 B.n405 B.n327 10.6151
R1958 B.n399 B.n327 10.6151
R1959 B.n399 B.n398 10.6151
R1960 B.n396 B.n331 10.6151
R1961 B.n390 B.n331 10.6151
R1962 B.n390 B.n389 10.6151
R1963 B.n389 B.n388 10.6151
R1964 B.n388 B.n333 10.6151
R1965 B.n382 B.n333 10.6151
R1966 B.n382 B.n381 10.6151
R1967 B.n381 B.n380 10.6151
R1968 B.n380 B.n335 10.6151
R1969 B.n374 B.n373 10.6151
R1970 B.n373 B.n372 10.6151
R1971 B.n372 B.n340 10.6151
R1972 B.n366 B.n340 10.6151
R1973 B.n366 B.n365 10.6151
R1974 B.n365 B.n364 10.6151
R1975 B.n364 B.n342 10.6151
R1976 B.n358 B.n342 10.6151
R1977 B.n358 B.n357 10.6151
R1978 B.n357 B.n356 10.6151
R1979 B.n356 B.n344 10.6151
R1980 B.n350 B.n344 10.6151
R1981 B.n350 B.n349 10.6151
R1982 B.n349 B.n348 10.6151
R1983 B.n348 B.n317 10.6151
R1984 B.n428 B.n313 10.6151
R1985 B.n438 B.n313 10.6151
R1986 B.n439 B.n438 10.6151
R1987 B.n440 B.n439 10.6151
R1988 B.n440 B.n305 10.6151
R1989 B.n450 B.n305 10.6151
R1990 B.n451 B.n450 10.6151
R1991 B.n452 B.n451 10.6151
R1992 B.n452 B.n297 10.6151
R1993 B.n462 B.n297 10.6151
R1994 B.n463 B.n462 10.6151
R1995 B.n464 B.n463 10.6151
R1996 B.n464 B.n289 10.6151
R1997 B.n474 B.n289 10.6151
R1998 B.n475 B.n474 10.6151
R1999 B.n476 B.n475 10.6151
R2000 B.n476 B.n281 10.6151
R2001 B.n486 B.n281 10.6151
R2002 B.n487 B.n486 10.6151
R2003 B.n488 B.n487 10.6151
R2004 B.n488 B.n273 10.6151
R2005 B.n499 B.n273 10.6151
R2006 B.n500 B.n499 10.6151
R2007 B.n501 B.n500 10.6151
R2008 B.n501 B.n266 10.6151
R2009 B.n511 B.n266 10.6151
R2010 B.n512 B.n511 10.6151
R2011 B.n513 B.n512 10.6151
R2012 B.n513 B.n258 10.6151
R2013 B.n523 B.n258 10.6151
R2014 B.n524 B.n523 10.6151
R2015 B.n525 B.n524 10.6151
R2016 B.n525 B.n250 10.6151
R2017 B.n536 B.n250 10.6151
R2018 B.n537 B.n536 10.6151
R2019 B.n538 B.n537 10.6151
R2020 B.n538 B.n243 10.6151
R2021 B.n548 B.n243 10.6151
R2022 B.n549 B.n548 10.6151
R2023 B.n550 B.n549 10.6151
R2024 B.n550 B.n235 10.6151
R2025 B.n560 B.n235 10.6151
R2026 B.n561 B.n560 10.6151
R2027 B.n562 B.n561 10.6151
R2028 B.n562 B.n227 10.6151
R2029 B.n573 B.n227 10.6151
R2030 B.n574 B.n573 10.6151
R2031 B.n575 B.n574 10.6151
R2032 B.n575 B.n220 10.6151
R2033 B.n585 B.n220 10.6151
R2034 B.n586 B.n585 10.6151
R2035 B.n587 B.n586 10.6151
R2036 B.n587 B.n212 10.6151
R2037 B.n597 B.n212 10.6151
R2038 B.n598 B.n597 10.6151
R2039 B.n599 B.n598 10.6151
R2040 B.n599 B.n204 10.6151
R2041 B.n609 B.n204 10.6151
R2042 B.n610 B.n609 10.6151
R2043 B.n611 B.n610 10.6151
R2044 B.n611 B.n196 10.6151
R2045 B.n621 B.n196 10.6151
R2046 B.n622 B.n621 10.6151
R2047 B.n623 B.n622 10.6151
R2048 B.n623 B.n188 10.6151
R2049 B.n633 B.n188 10.6151
R2050 B.n634 B.n633 10.6151
R2051 B.n635 B.n634 10.6151
R2052 B.n635 B.n180 10.6151
R2053 B.n645 B.n180 10.6151
R2054 B.n646 B.n645 10.6151
R2055 B.n647 B.n646 10.6151
R2056 B.n647 B.n172 10.6151
R2057 B.n658 B.n172 10.6151
R2058 B.n659 B.n658 10.6151
R2059 B.n660 B.n659 10.6151
R2060 B.n660 B.n0 10.6151
R2061 B.n1001 B.n1 10.6151
R2062 B.n1001 B.n1000 10.6151
R2063 B.n1000 B.n999 10.6151
R2064 B.n999 B.n10 10.6151
R2065 B.n993 B.n10 10.6151
R2066 B.n993 B.n992 10.6151
R2067 B.n992 B.n991 10.6151
R2068 B.n991 B.n17 10.6151
R2069 B.n985 B.n17 10.6151
R2070 B.n985 B.n984 10.6151
R2071 B.n984 B.n983 10.6151
R2072 B.n983 B.n24 10.6151
R2073 B.n977 B.n24 10.6151
R2074 B.n977 B.n976 10.6151
R2075 B.n976 B.n975 10.6151
R2076 B.n975 B.n31 10.6151
R2077 B.n969 B.n31 10.6151
R2078 B.n969 B.n968 10.6151
R2079 B.n968 B.n967 10.6151
R2080 B.n967 B.n38 10.6151
R2081 B.n961 B.n38 10.6151
R2082 B.n961 B.n960 10.6151
R2083 B.n960 B.n959 10.6151
R2084 B.n959 B.n45 10.6151
R2085 B.n953 B.n45 10.6151
R2086 B.n953 B.n952 10.6151
R2087 B.n952 B.n951 10.6151
R2088 B.n951 B.n52 10.6151
R2089 B.n945 B.n52 10.6151
R2090 B.n945 B.n944 10.6151
R2091 B.n944 B.n943 10.6151
R2092 B.n943 B.n58 10.6151
R2093 B.n937 B.n58 10.6151
R2094 B.n937 B.n936 10.6151
R2095 B.n936 B.n935 10.6151
R2096 B.n935 B.n66 10.6151
R2097 B.n929 B.n66 10.6151
R2098 B.n929 B.n928 10.6151
R2099 B.n928 B.n927 10.6151
R2100 B.n927 B.n73 10.6151
R2101 B.n921 B.n73 10.6151
R2102 B.n921 B.n920 10.6151
R2103 B.n920 B.n919 10.6151
R2104 B.n919 B.n79 10.6151
R2105 B.n913 B.n79 10.6151
R2106 B.n913 B.n912 10.6151
R2107 B.n912 B.n911 10.6151
R2108 B.n911 B.n87 10.6151
R2109 B.n905 B.n87 10.6151
R2110 B.n905 B.n904 10.6151
R2111 B.n904 B.n903 10.6151
R2112 B.n903 B.n94 10.6151
R2113 B.n897 B.n94 10.6151
R2114 B.n897 B.n896 10.6151
R2115 B.n896 B.n895 10.6151
R2116 B.n895 B.n100 10.6151
R2117 B.n889 B.n100 10.6151
R2118 B.n889 B.n888 10.6151
R2119 B.n888 B.n887 10.6151
R2120 B.n887 B.n108 10.6151
R2121 B.n881 B.n108 10.6151
R2122 B.n881 B.n880 10.6151
R2123 B.n880 B.n879 10.6151
R2124 B.n879 B.n115 10.6151
R2125 B.n873 B.n115 10.6151
R2126 B.n873 B.n872 10.6151
R2127 B.n872 B.n871 10.6151
R2128 B.n871 B.n122 10.6151
R2129 B.n865 B.n122 10.6151
R2130 B.n865 B.n864 10.6151
R2131 B.n864 B.n863 10.6151
R2132 B.n863 B.n129 10.6151
R2133 B.n857 B.n129 10.6151
R2134 B.n857 B.n856 10.6151
R2135 B.n856 B.n855 10.6151
R2136 B.n855 B.n136 10.6151
R2137 B.n849 B.n136 10.6151
R2138 B.t6 B.n202 10.168
R2139 B.t1 B.n36 10.168
R2140 B.n817 B.n816 9.36635
R2141 B.n794 B.n159 9.36635
R2142 B.n398 B.n397 9.36635
R2143 B.n374 B.n339 9.36635
R2144 B.n1007 B.n0 2.81026
R2145 B.n1007 B.n1 2.81026
R2146 B.t11 B.n299 2.54238
R2147 B.n868 B.t15 2.54238
R2148 B.n816 B.n815 1.24928
R2149 B.n798 B.n159 1.24928
R2150 B.n397 B.n396 1.24928
R2151 B.n339 B.n335 1.24928
R2152 VP.n32 VP.n29 161.3
R2153 VP.n34 VP.n33 161.3
R2154 VP.n35 VP.n28 161.3
R2155 VP.n37 VP.n36 161.3
R2156 VP.n38 VP.n27 161.3
R2157 VP.n40 VP.n39 161.3
R2158 VP.n41 VP.n26 161.3
R2159 VP.n44 VP.n43 161.3
R2160 VP.n45 VP.n25 161.3
R2161 VP.n47 VP.n46 161.3
R2162 VP.n48 VP.n24 161.3
R2163 VP.n50 VP.n49 161.3
R2164 VP.n51 VP.n23 161.3
R2165 VP.n53 VP.n52 161.3
R2166 VP.n54 VP.n22 161.3
R2167 VP.n57 VP.n56 161.3
R2168 VP.n58 VP.n21 161.3
R2169 VP.n60 VP.n59 161.3
R2170 VP.n61 VP.n20 161.3
R2171 VP.n63 VP.n62 161.3
R2172 VP.n64 VP.n19 161.3
R2173 VP.n66 VP.n65 161.3
R2174 VP.n67 VP.n18 161.3
R2175 VP.n69 VP.n68 161.3
R2176 VP.n123 VP.n122 161.3
R2177 VP.n121 VP.n1 161.3
R2178 VP.n120 VP.n119 161.3
R2179 VP.n118 VP.n2 161.3
R2180 VP.n117 VP.n116 161.3
R2181 VP.n115 VP.n3 161.3
R2182 VP.n114 VP.n113 161.3
R2183 VP.n112 VP.n4 161.3
R2184 VP.n111 VP.n110 161.3
R2185 VP.n108 VP.n5 161.3
R2186 VP.n107 VP.n106 161.3
R2187 VP.n105 VP.n6 161.3
R2188 VP.n104 VP.n103 161.3
R2189 VP.n102 VP.n7 161.3
R2190 VP.n101 VP.n100 161.3
R2191 VP.n99 VP.n8 161.3
R2192 VP.n98 VP.n97 161.3
R2193 VP.n95 VP.n9 161.3
R2194 VP.n94 VP.n93 161.3
R2195 VP.n92 VP.n10 161.3
R2196 VP.n91 VP.n90 161.3
R2197 VP.n89 VP.n11 161.3
R2198 VP.n88 VP.n87 161.3
R2199 VP.n86 VP.n12 161.3
R2200 VP.n85 VP.n84 161.3
R2201 VP.n82 VP.n13 161.3
R2202 VP.n81 VP.n80 161.3
R2203 VP.n79 VP.n14 161.3
R2204 VP.n78 VP.n77 161.3
R2205 VP.n76 VP.n15 161.3
R2206 VP.n75 VP.n74 161.3
R2207 VP.n73 VP.n16 161.3
R2208 VP.n72 VP.n71 80.9007
R2209 VP.n124 VP.n0 80.9007
R2210 VP.n70 VP.n17 80.9007
R2211 VP.n31 VP.n30 63.9939
R2212 VP.n77 VP.n14 56.5617
R2213 VP.n116 VP.n2 56.5617
R2214 VP.n62 VP.n19 56.5617
R2215 VP.n90 VP.n10 56.5617
R2216 VP.n103 VP.n6 56.5617
R2217 VP.n49 VP.n23 56.5617
R2218 VP.n36 VP.n27 56.5617
R2219 VP.n31 VP.t1 55.7437
R2220 VP.n72 VP.n70 52.3518
R2221 VP.n75 VP.n16 24.5923
R2222 VP.n76 VP.n75 24.5923
R2223 VP.n77 VP.n76 24.5923
R2224 VP.n81 VP.n14 24.5923
R2225 VP.n82 VP.n81 24.5923
R2226 VP.n84 VP.n82 24.5923
R2227 VP.n88 VP.n12 24.5923
R2228 VP.n89 VP.n88 24.5923
R2229 VP.n90 VP.n89 24.5923
R2230 VP.n94 VP.n10 24.5923
R2231 VP.n95 VP.n94 24.5923
R2232 VP.n97 VP.n95 24.5923
R2233 VP.n101 VP.n8 24.5923
R2234 VP.n102 VP.n101 24.5923
R2235 VP.n103 VP.n102 24.5923
R2236 VP.n107 VP.n6 24.5923
R2237 VP.n108 VP.n107 24.5923
R2238 VP.n110 VP.n108 24.5923
R2239 VP.n114 VP.n4 24.5923
R2240 VP.n115 VP.n114 24.5923
R2241 VP.n116 VP.n115 24.5923
R2242 VP.n120 VP.n2 24.5923
R2243 VP.n121 VP.n120 24.5923
R2244 VP.n122 VP.n121 24.5923
R2245 VP.n66 VP.n19 24.5923
R2246 VP.n67 VP.n66 24.5923
R2247 VP.n68 VP.n67 24.5923
R2248 VP.n53 VP.n23 24.5923
R2249 VP.n54 VP.n53 24.5923
R2250 VP.n56 VP.n54 24.5923
R2251 VP.n60 VP.n21 24.5923
R2252 VP.n61 VP.n60 24.5923
R2253 VP.n62 VP.n61 24.5923
R2254 VP.n40 VP.n27 24.5923
R2255 VP.n41 VP.n40 24.5923
R2256 VP.n43 VP.n41 24.5923
R2257 VP.n47 VP.n25 24.5923
R2258 VP.n48 VP.n47 24.5923
R2259 VP.n49 VP.n48 24.5923
R2260 VP.n34 VP.n29 24.5923
R2261 VP.n35 VP.n34 24.5923
R2262 VP.n36 VP.n35 24.5923
R2263 VP.n71 VP.t9 22.3791
R2264 VP.n83 VP.t7 22.3791
R2265 VP.n96 VP.t4 22.3791
R2266 VP.n109 VP.t5 22.3791
R2267 VP.n0 VP.t2 22.3791
R2268 VP.n17 VP.t6 22.3791
R2269 VP.n55 VP.t3 22.3791
R2270 VP.n42 VP.t0 22.3791
R2271 VP.n30 VP.t8 22.3791
R2272 VP.n84 VP.n83 13.7719
R2273 VP.n109 VP.n4 13.7719
R2274 VP.n55 VP.n21 13.7719
R2275 VP.n97 VP.n96 12.2964
R2276 VP.n96 VP.n8 12.2964
R2277 VP.n43 VP.n42 12.2964
R2278 VP.n42 VP.n25 12.2964
R2279 VP.n83 VP.n12 10.8209
R2280 VP.n110 VP.n109 10.8209
R2281 VP.n56 VP.n55 10.8209
R2282 VP.n30 VP.n29 10.8209
R2283 VP.n71 VP.n16 9.3454
R2284 VP.n122 VP.n0 9.3454
R2285 VP.n68 VP.n17 9.3454
R2286 VP.n32 VP.n31 3.16704
R2287 VP.n70 VP.n69 0.354861
R2288 VP.n73 VP.n72 0.354861
R2289 VP.n124 VP.n123 0.354861
R2290 VP VP.n124 0.267071
R2291 VP.n33 VP.n32 0.189894
R2292 VP.n33 VP.n28 0.189894
R2293 VP.n37 VP.n28 0.189894
R2294 VP.n38 VP.n37 0.189894
R2295 VP.n39 VP.n38 0.189894
R2296 VP.n39 VP.n26 0.189894
R2297 VP.n44 VP.n26 0.189894
R2298 VP.n45 VP.n44 0.189894
R2299 VP.n46 VP.n45 0.189894
R2300 VP.n46 VP.n24 0.189894
R2301 VP.n50 VP.n24 0.189894
R2302 VP.n51 VP.n50 0.189894
R2303 VP.n52 VP.n51 0.189894
R2304 VP.n52 VP.n22 0.189894
R2305 VP.n57 VP.n22 0.189894
R2306 VP.n58 VP.n57 0.189894
R2307 VP.n59 VP.n58 0.189894
R2308 VP.n59 VP.n20 0.189894
R2309 VP.n63 VP.n20 0.189894
R2310 VP.n64 VP.n63 0.189894
R2311 VP.n65 VP.n64 0.189894
R2312 VP.n65 VP.n18 0.189894
R2313 VP.n69 VP.n18 0.189894
R2314 VP.n74 VP.n73 0.189894
R2315 VP.n74 VP.n15 0.189894
R2316 VP.n78 VP.n15 0.189894
R2317 VP.n79 VP.n78 0.189894
R2318 VP.n80 VP.n79 0.189894
R2319 VP.n80 VP.n13 0.189894
R2320 VP.n85 VP.n13 0.189894
R2321 VP.n86 VP.n85 0.189894
R2322 VP.n87 VP.n86 0.189894
R2323 VP.n87 VP.n11 0.189894
R2324 VP.n91 VP.n11 0.189894
R2325 VP.n92 VP.n91 0.189894
R2326 VP.n93 VP.n92 0.189894
R2327 VP.n93 VP.n9 0.189894
R2328 VP.n98 VP.n9 0.189894
R2329 VP.n99 VP.n98 0.189894
R2330 VP.n100 VP.n99 0.189894
R2331 VP.n100 VP.n7 0.189894
R2332 VP.n104 VP.n7 0.189894
R2333 VP.n105 VP.n104 0.189894
R2334 VP.n106 VP.n105 0.189894
R2335 VP.n106 VP.n5 0.189894
R2336 VP.n111 VP.n5 0.189894
R2337 VP.n112 VP.n111 0.189894
R2338 VP.n113 VP.n112 0.189894
R2339 VP.n113 VP.n3 0.189894
R2340 VP.n117 VP.n3 0.189894
R2341 VP.n118 VP.n117 0.189894
R2342 VP.n119 VP.n118 0.189894
R2343 VP.n119 VP.n1 0.189894
R2344 VP.n123 VP.n1 0.189894
R2345 VDD1.n10 VDD1.n0 289.615
R2346 VDD1.n27 VDD1.n17 289.615
R2347 VDD1.n11 VDD1.n10 185
R2348 VDD1.n9 VDD1.n8 185
R2349 VDD1.n4 VDD1.n3 185
R2350 VDD1.n21 VDD1.n20 185
R2351 VDD1.n26 VDD1.n25 185
R2352 VDD1.n28 VDD1.n27 185
R2353 VDD1.n5 VDD1.t8 150.499
R2354 VDD1.n22 VDD1.t0 150.499
R2355 VDD1.n10 VDD1.n9 104.615
R2356 VDD1.n9 VDD1.n3 104.615
R2357 VDD1.n26 VDD1.n20 104.615
R2358 VDD1.n27 VDD1.n26 104.615
R2359 VDD1.n35 VDD1.n34 79.443
R2360 VDD1.n37 VDD1.n36 76.9315
R2361 VDD1.n16 VDD1.n15 76.9315
R2362 VDD1.n33 VDD1.n32 76.9315
R2363 VDD1.t8 VDD1.n3 52.3082
R2364 VDD1.t0 VDD1.n20 52.3082
R2365 VDD1.n16 VDD1.n14 50.3472
R2366 VDD1.n33 VDD1.n31 50.3472
R2367 VDD1.n37 VDD1.n35 45.1798
R2368 VDD1.n5 VDD1.n4 10.2326
R2369 VDD1.n22 VDD1.n21 10.2326
R2370 VDD1.n14 VDD1.n0 9.69747
R2371 VDD1.n31 VDD1.n17 9.69747
R2372 VDD1.n14 VDD1.n13 9.45567
R2373 VDD1.n31 VDD1.n30 9.45567
R2374 VDD1.n2 VDD1.n1 9.3005
R2375 VDD1.n13 VDD1.n12 9.3005
R2376 VDD1.n7 VDD1.n6 9.3005
R2377 VDD1.n24 VDD1.n23 9.3005
R2378 VDD1.n19 VDD1.n18 9.3005
R2379 VDD1.n30 VDD1.n29 9.3005
R2380 VDD1.n12 VDD1.n11 8.92171
R2381 VDD1.n29 VDD1.n28 8.92171
R2382 VDD1.n8 VDD1.n2 8.14595
R2383 VDD1.n25 VDD1.n19 8.14595
R2384 VDD1.n7 VDD1.n4 7.3702
R2385 VDD1.n24 VDD1.n21 7.3702
R2386 VDD1.n36 VDD1.t6 5.85849
R2387 VDD1.n36 VDD1.t3 5.85849
R2388 VDD1.n15 VDD1.t1 5.85849
R2389 VDD1.n15 VDD1.t9 5.85849
R2390 VDD1.n34 VDD1.t4 5.85849
R2391 VDD1.n34 VDD1.t7 5.85849
R2392 VDD1.n32 VDD1.t2 5.85849
R2393 VDD1.n32 VDD1.t5 5.85849
R2394 VDD1.n8 VDD1.n7 5.81868
R2395 VDD1.n25 VDD1.n24 5.81868
R2396 VDD1.n11 VDD1.n2 5.04292
R2397 VDD1.n28 VDD1.n19 5.04292
R2398 VDD1.n12 VDD1.n0 4.26717
R2399 VDD1.n29 VDD1.n17 4.26717
R2400 VDD1.n6 VDD1.n5 2.88718
R2401 VDD1.n23 VDD1.n22 2.88718
R2402 VDD1 VDD1.n37 2.50912
R2403 VDD1 VDD1.n16 0.914293
R2404 VDD1.n35 VDD1.n33 0.800757
R2405 VDD1.n13 VDD1.n1 0.155672
R2406 VDD1.n6 VDD1.n1 0.155672
R2407 VDD1.n23 VDD1.n18 0.155672
R2408 VDD1.n30 VDD1.n18 0.155672
C0 VP VDD2 0.722029f
C1 VN VDD2 3.57624f
C2 VTAIL VDD2 7.55563f
C3 VDD1 VP 4.13311f
C4 VN VDD1 0.161065f
C5 VDD1 VTAIL 7.49544f
C6 VDD1 VDD2 2.85248f
C7 VN VP 8.332139f
C8 VTAIL VP 5.43259f
C9 VN VTAIL 5.4184f
C10 VDD2 B 7.04736f
C11 VDD1 B 6.904426f
C12 VTAIL B 4.882223f
C13 VN B 22.32426f
C14 VP B 20.751549f
C15 VDD1.n0 B 0.043583f
C16 VDD1.n1 B 0.029587f
C17 VDD1.n2 B 0.015899f
C18 VDD1.n3 B 0.028184f
C19 VDD1.n4 B 0.026311f
C20 VDD1.t8 B 0.065769f
C21 VDD1.n5 B 0.119372f
C22 VDD1.n6 B 0.350837f
C23 VDD1.n7 B 0.015899f
C24 VDD1.n8 B 0.016834f
C25 VDD1.n9 B 0.037578f
C26 VDD1.n10 B 0.084881f
C27 VDD1.n11 B 0.016834f
C28 VDD1.n12 B 0.015899f
C29 VDD1.n13 B 0.064346f
C30 VDD1.n14 B 0.094088f
C31 VDD1.t1 B 0.079025f
C32 VDD1.t9 B 0.079025f
C33 VDD1.n15 B 0.586606f
C34 VDD1.n16 B 1.00905f
C35 VDD1.n17 B 0.043583f
C36 VDD1.n18 B 0.029587f
C37 VDD1.n19 B 0.015899f
C38 VDD1.n20 B 0.028184f
C39 VDD1.n21 B 0.026311f
C40 VDD1.t0 B 0.065769f
C41 VDD1.n22 B 0.119372f
C42 VDD1.n23 B 0.350837f
C43 VDD1.n24 B 0.015899f
C44 VDD1.n25 B 0.016834f
C45 VDD1.n26 B 0.037578f
C46 VDD1.n27 B 0.084881f
C47 VDD1.n28 B 0.016834f
C48 VDD1.n29 B 0.015899f
C49 VDD1.n30 B 0.064346f
C50 VDD1.n31 B 0.094088f
C51 VDD1.t2 B 0.079025f
C52 VDD1.t5 B 0.079025f
C53 VDD1.n32 B 0.586604f
C54 VDD1.n33 B 0.999085f
C55 VDD1.t4 B 0.079025f
C56 VDD1.t7 B 0.079025f
C57 VDD1.n34 B 0.612481f
C58 VDD1.n35 B 3.62995f
C59 VDD1.t6 B 0.079025f
C60 VDD1.t3 B 0.079025f
C61 VDD1.n36 B 0.586606f
C62 VDD1.n37 B 3.47933f
C63 VP.t2 B 0.733307f
C64 VP.n0 B 0.385552f
C65 VP.n1 B 0.023595f
C66 VP.n2 B 0.037237f
C67 VP.n3 B 0.023595f
C68 VP.n4 B 0.03425f
C69 VP.n5 B 0.023595f
C70 VP.n6 B 0.035278f
C71 VP.n7 B 0.023595f
C72 VP.n8 B 0.032954f
C73 VP.n9 B 0.023595f
C74 VP.n10 B 0.03332f
C75 VP.n11 B 0.023595f
C76 VP.n12 B 0.031658f
C77 VP.n13 B 0.023595f
C78 VP.n14 B 0.031361f
C79 VP.n15 B 0.023595f
C80 VP.n16 B 0.030362f
C81 VP.t6 B 0.733307f
C82 VP.n17 B 0.385552f
C83 VP.n18 B 0.023595f
C84 VP.n19 B 0.037237f
C85 VP.n20 B 0.023595f
C86 VP.n21 B 0.03425f
C87 VP.n22 B 0.023595f
C88 VP.n23 B 0.035278f
C89 VP.n24 B 0.023595f
C90 VP.n25 B 0.032954f
C91 VP.n26 B 0.023595f
C92 VP.n27 B 0.03332f
C93 VP.n28 B 0.023595f
C94 VP.n29 B 0.031658f
C95 VP.t1 B 1.01598f
C96 VP.t8 B 0.733307f
C97 VP.n30 B 0.373286f
C98 VP.n31 B 0.378466f
C99 VP.n32 B 0.295591f
C100 VP.n33 B 0.023595f
C101 VP.n34 B 0.043755f
C102 VP.n35 B 0.043755f
C103 VP.n36 B 0.035278f
C104 VP.n37 B 0.023595f
C105 VP.n38 B 0.023595f
C106 VP.n39 B 0.023595f
C107 VP.n40 B 0.043755f
C108 VP.n41 B 0.043755f
C109 VP.t0 B 0.733307f
C110 VP.n42 B 0.29278f
C111 VP.n43 B 0.032954f
C112 VP.n44 B 0.023595f
C113 VP.n45 B 0.023595f
C114 VP.n46 B 0.023595f
C115 VP.n47 B 0.043755f
C116 VP.n48 B 0.043755f
C117 VP.n49 B 0.03332f
C118 VP.n50 B 0.023595f
C119 VP.n51 B 0.023595f
C120 VP.n52 B 0.023595f
C121 VP.n53 B 0.043755f
C122 VP.n54 B 0.043755f
C123 VP.t3 B 0.733307f
C124 VP.n55 B 0.29278f
C125 VP.n56 B 0.031658f
C126 VP.n57 B 0.023595f
C127 VP.n58 B 0.023595f
C128 VP.n59 B 0.023595f
C129 VP.n60 B 0.043755f
C130 VP.n61 B 0.043755f
C131 VP.n62 B 0.031361f
C132 VP.n63 B 0.023595f
C133 VP.n64 B 0.023595f
C134 VP.n65 B 0.023595f
C135 VP.n66 B 0.043755f
C136 VP.n67 B 0.043755f
C137 VP.n68 B 0.030362f
C138 VP.n69 B 0.038076f
C139 VP.n70 B 1.44237f
C140 VP.t9 B 0.733307f
C141 VP.n71 B 0.385552f
C142 VP.n72 B 1.45862f
C143 VP.n73 B 0.038076f
C144 VP.n74 B 0.023595f
C145 VP.n75 B 0.043755f
C146 VP.n76 B 0.043755f
C147 VP.n77 B 0.037237f
C148 VP.n78 B 0.023595f
C149 VP.n79 B 0.023595f
C150 VP.n80 B 0.023595f
C151 VP.n81 B 0.043755f
C152 VP.n82 B 0.043755f
C153 VP.t7 B 0.733307f
C154 VP.n83 B 0.29278f
C155 VP.n84 B 0.03425f
C156 VP.n85 B 0.023595f
C157 VP.n86 B 0.023595f
C158 VP.n87 B 0.023595f
C159 VP.n88 B 0.043755f
C160 VP.n89 B 0.043755f
C161 VP.n90 B 0.035278f
C162 VP.n91 B 0.023595f
C163 VP.n92 B 0.023595f
C164 VP.n93 B 0.023595f
C165 VP.n94 B 0.043755f
C166 VP.n95 B 0.043755f
C167 VP.t4 B 0.733307f
C168 VP.n96 B 0.29278f
C169 VP.n97 B 0.032954f
C170 VP.n98 B 0.023595f
C171 VP.n99 B 0.023595f
C172 VP.n100 B 0.023595f
C173 VP.n101 B 0.043755f
C174 VP.n102 B 0.043755f
C175 VP.n103 B 0.03332f
C176 VP.n104 B 0.023595f
C177 VP.n105 B 0.023595f
C178 VP.n106 B 0.023595f
C179 VP.n107 B 0.043755f
C180 VP.n108 B 0.043755f
C181 VP.t5 B 0.733307f
C182 VP.n109 B 0.29278f
C183 VP.n110 B 0.031658f
C184 VP.n111 B 0.023595f
C185 VP.n112 B 0.023595f
C186 VP.n113 B 0.023595f
C187 VP.n114 B 0.043755f
C188 VP.n115 B 0.043755f
C189 VP.n116 B 0.031361f
C190 VP.n117 B 0.023595f
C191 VP.n118 B 0.023595f
C192 VP.n119 B 0.023595f
C193 VP.n120 B 0.043755f
C194 VP.n121 B 0.043755f
C195 VP.n122 B 0.030362f
C196 VP.n123 B 0.038076f
C197 VP.n124 B 0.065468f
C198 VDD2.n0 B 0.042702f
C199 VDD2.n1 B 0.028989f
C200 VDD2.n2 B 0.015577f
C201 VDD2.n3 B 0.027615f
C202 VDD2.n4 B 0.025779f
C203 VDD2.t9 B 0.06444f
C204 VDD2.n5 B 0.116961f
C205 VDD2.n6 B 0.343749f
C206 VDD2.n7 B 0.015577f
C207 VDD2.n8 B 0.016494f
C208 VDD2.n9 B 0.036819f
C209 VDD2.n10 B 0.083167f
C210 VDD2.n11 B 0.016494f
C211 VDD2.n12 B 0.015577f
C212 VDD2.n13 B 0.063047f
C213 VDD2.n14 B 0.092187f
C214 VDD2.t7 B 0.077429f
C215 VDD2.t4 B 0.077429f
C216 VDD2.n15 B 0.574754f
C217 VDD2.n16 B 0.978901f
C218 VDD2.t5 B 0.077429f
C219 VDD2.t2 B 0.077429f
C220 VDD2.n17 B 0.600107f
C221 VDD2.n18 B 3.38827f
C222 VDD2.n19 B 0.042702f
C223 VDD2.n20 B 0.028989f
C224 VDD2.n21 B 0.015577f
C225 VDD2.n22 B 0.027615f
C226 VDD2.n23 B 0.025779f
C227 VDD2.t3 B 0.06444f
C228 VDD2.n24 B 0.116961f
C229 VDD2.n25 B 0.343749f
C230 VDD2.n26 B 0.015577f
C231 VDD2.n27 B 0.016494f
C232 VDD2.n28 B 0.036819f
C233 VDD2.n29 B 0.083167f
C234 VDD2.n30 B 0.016494f
C235 VDD2.n31 B 0.015577f
C236 VDD2.n32 B 0.063047f
C237 VDD2.n33 B 0.066815f
C238 VDD2.n34 B 3.04212f
C239 VDD2.t8 B 0.077429f
C240 VDD2.t0 B 0.077429f
C241 VDD2.n35 B 0.574756f
C242 VDD2.n36 B 0.640797f
C243 VDD2.t6 B 0.077429f
C244 VDD2.t1 B 0.077429f
C245 VDD2.n37 B 0.600065f
C246 VTAIL.t16 B 0.091786f
C247 VTAIL.t11 B 0.091786f
C248 VTAIL.n0 B 0.605777f
C249 VTAIL.n1 B 0.840489f
C250 VTAIL.n2 B 0.050621f
C251 VTAIL.n3 B 0.034364f
C252 VTAIL.n4 B 0.018466f
C253 VTAIL.n5 B 0.032735f
C254 VTAIL.n6 B 0.03056f
C255 VTAIL.t8 B 0.07639f
C256 VTAIL.n7 B 0.138648f
C257 VTAIL.n8 B 0.40749f
C258 VTAIL.n9 B 0.018466f
C259 VTAIL.n10 B 0.019552f
C260 VTAIL.n11 B 0.043647f
C261 VTAIL.n12 B 0.098588f
C262 VTAIL.n13 B 0.019552f
C263 VTAIL.n14 B 0.018466f
C264 VTAIL.n15 B 0.074737f
C265 VTAIL.n16 B 0.055437f
C266 VTAIL.n17 B 0.647172f
C267 VTAIL.t4 B 0.091786f
C268 VTAIL.t6 B 0.091786f
C269 VTAIL.n18 B 0.605777f
C270 VTAIL.n19 B 1.06624f
C271 VTAIL.t5 B 0.091786f
C272 VTAIL.t0 B 0.091786f
C273 VTAIL.n20 B 0.605777f
C274 VTAIL.n21 B 2.23465f
C275 VTAIL.t17 B 0.091786f
C276 VTAIL.t14 B 0.091786f
C277 VTAIL.n22 B 0.60578f
C278 VTAIL.n23 B 2.23464f
C279 VTAIL.t18 B 0.091786f
C280 VTAIL.t19 B 0.091786f
C281 VTAIL.n24 B 0.60578f
C282 VTAIL.n25 B 1.06624f
C283 VTAIL.n26 B 0.050621f
C284 VTAIL.n27 B 0.034364f
C285 VTAIL.n28 B 0.018466f
C286 VTAIL.n29 B 0.032735f
C287 VTAIL.n30 B 0.03056f
C288 VTAIL.t10 B 0.07639f
C289 VTAIL.n31 B 0.138648f
C290 VTAIL.n32 B 0.40749f
C291 VTAIL.n33 B 0.018466f
C292 VTAIL.n34 B 0.019552f
C293 VTAIL.n35 B 0.043647f
C294 VTAIL.n36 B 0.098588f
C295 VTAIL.n37 B 0.019552f
C296 VTAIL.n38 B 0.018466f
C297 VTAIL.n39 B 0.074737f
C298 VTAIL.n40 B 0.055437f
C299 VTAIL.n41 B 0.647172f
C300 VTAIL.t2 B 0.091786f
C301 VTAIL.t1 B 0.091786f
C302 VTAIL.n42 B 0.60578f
C303 VTAIL.n43 B 0.928783f
C304 VTAIL.t9 B 0.091786f
C305 VTAIL.t7 B 0.091786f
C306 VTAIL.n44 B 0.60578f
C307 VTAIL.n45 B 1.06624f
C308 VTAIL.n46 B 0.050621f
C309 VTAIL.n47 B 0.034364f
C310 VTAIL.n48 B 0.018466f
C311 VTAIL.n49 B 0.032735f
C312 VTAIL.n50 B 0.03056f
C313 VTAIL.t3 B 0.07639f
C314 VTAIL.n51 B 0.138648f
C315 VTAIL.n52 B 0.40749f
C316 VTAIL.n53 B 0.018466f
C317 VTAIL.n54 B 0.019552f
C318 VTAIL.n55 B 0.043647f
C319 VTAIL.n56 B 0.098588f
C320 VTAIL.n57 B 0.019552f
C321 VTAIL.n58 B 0.018466f
C322 VTAIL.n59 B 0.074737f
C323 VTAIL.n60 B 0.055437f
C324 VTAIL.n61 B 1.57407f
C325 VTAIL.n62 B 0.050621f
C326 VTAIL.n63 B 0.034364f
C327 VTAIL.n64 B 0.018466f
C328 VTAIL.n65 B 0.032735f
C329 VTAIL.n66 B 0.03056f
C330 VTAIL.t15 B 0.07639f
C331 VTAIL.n67 B 0.138648f
C332 VTAIL.n68 B 0.40749f
C333 VTAIL.n69 B 0.018466f
C334 VTAIL.n70 B 0.019552f
C335 VTAIL.n71 B 0.043647f
C336 VTAIL.n72 B 0.098588f
C337 VTAIL.n73 B 0.019552f
C338 VTAIL.n74 B 0.018466f
C339 VTAIL.n75 B 0.074737f
C340 VTAIL.n76 B 0.055437f
C341 VTAIL.n77 B 1.57407f
C342 VTAIL.t12 B 0.091786f
C343 VTAIL.t13 B 0.091786f
C344 VTAIL.n78 B 0.605777f
C345 VTAIL.n79 B 0.775578f
C346 VN.t7 B 0.711383f
C347 VN.n0 B 0.374025f
C348 VN.n1 B 0.02289f
C349 VN.n2 B 0.036123f
C350 VN.n3 B 0.02289f
C351 VN.n4 B 0.033226f
C352 VN.n5 B 0.02289f
C353 VN.n6 B 0.034223f
C354 VN.n7 B 0.02289f
C355 VN.n8 B 0.031969f
C356 VN.n9 B 0.02289f
C357 VN.n10 B 0.032324f
C358 VN.n11 B 0.02289f
C359 VN.n12 B 0.030712f
C360 VN.t2 B 0.711383f
C361 VN.n13 B 0.362125f
C362 VN.t0 B 0.985602f
C363 VN.n14 B 0.36715f
C364 VN.n15 B 0.286753f
C365 VN.n16 B 0.02289f
C366 VN.n17 B 0.042446f
C367 VN.n18 B 0.042446f
C368 VN.n19 B 0.034223f
C369 VN.n20 B 0.02289f
C370 VN.n21 B 0.02289f
C371 VN.n22 B 0.02289f
C372 VN.n23 B 0.042446f
C373 VN.n24 B 0.042446f
C374 VN.t5 B 0.711383f
C375 VN.n25 B 0.284026f
C376 VN.n26 B 0.031969f
C377 VN.n27 B 0.02289f
C378 VN.n28 B 0.02289f
C379 VN.n29 B 0.02289f
C380 VN.n30 B 0.042446f
C381 VN.n31 B 0.042446f
C382 VN.n32 B 0.032324f
C383 VN.n33 B 0.02289f
C384 VN.n34 B 0.02289f
C385 VN.n35 B 0.02289f
C386 VN.n36 B 0.042446f
C387 VN.n37 B 0.042446f
C388 VN.t4 B 0.711383f
C389 VN.n38 B 0.284026f
C390 VN.n39 B 0.030712f
C391 VN.n40 B 0.02289f
C392 VN.n41 B 0.02289f
C393 VN.n42 B 0.02289f
C394 VN.n43 B 0.042446f
C395 VN.n44 B 0.042446f
C396 VN.n45 B 0.030424f
C397 VN.n46 B 0.02289f
C398 VN.n47 B 0.02289f
C399 VN.n48 B 0.02289f
C400 VN.n49 B 0.042446f
C401 VN.n50 B 0.042446f
C402 VN.n51 B 0.029454f
C403 VN.n52 B 0.036937f
C404 VN.n53 B 0.063511f
C405 VN.t6 B 0.711383f
C406 VN.n54 B 0.374025f
C407 VN.n55 B 0.02289f
C408 VN.n56 B 0.036123f
C409 VN.n57 B 0.02289f
C410 VN.n58 B 0.033226f
C411 VN.n59 B 0.02289f
C412 VN.t1 B 0.711383f
C413 VN.n60 B 0.284026f
C414 VN.n61 B 0.034223f
C415 VN.n62 B 0.02289f
C416 VN.n63 B 0.031969f
C417 VN.n64 B 0.02289f
C418 VN.t9 B 0.711383f
C419 VN.n65 B 0.284026f
C420 VN.n66 B 0.032324f
C421 VN.n67 B 0.02289f
C422 VN.n68 B 0.030712f
C423 VN.t8 B 0.985602f
C424 VN.t3 B 0.711383f
C425 VN.n69 B 0.362125f
C426 VN.n70 B 0.36715f
C427 VN.n71 B 0.286753f
C428 VN.n72 B 0.02289f
C429 VN.n73 B 0.042446f
C430 VN.n74 B 0.042446f
C431 VN.n75 B 0.034223f
C432 VN.n76 B 0.02289f
C433 VN.n77 B 0.02289f
C434 VN.n78 B 0.02289f
C435 VN.n79 B 0.042446f
C436 VN.n80 B 0.042446f
C437 VN.n81 B 0.031969f
C438 VN.n82 B 0.02289f
C439 VN.n83 B 0.02289f
C440 VN.n84 B 0.02289f
C441 VN.n85 B 0.042446f
C442 VN.n86 B 0.042446f
C443 VN.n87 B 0.032324f
C444 VN.n88 B 0.02289f
C445 VN.n89 B 0.02289f
C446 VN.n90 B 0.02289f
C447 VN.n91 B 0.042446f
C448 VN.n92 B 0.042446f
C449 VN.n93 B 0.030712f
C450 VN.n94 B 0.02289f
C451 VN.n95 B 0.02289f
C452 VN.n96 B 0.02289f
C453 VN.n97 B 0.042446f
C454 VN.n98 B 0.042446f
C455 VN.n99 B 0.030424f
C456 VN.n100 B 0.02289f
C457 VN.n101 B 0.02289f
C458 VN.n102 B 0.02289f
C459 VN.n103 B 0.042446f
C460 VN.n104 B 0.042446f
C461 VN.n105 B 0.029454f
C462 VN.n106 B 0.036937f
C463 VN.n107 B 1.40846f
.ends

