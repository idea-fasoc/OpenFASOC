* NGSPICE file created from diff_pair_sample_1716.ext - technology: sky130A

.subckt diff_pair_sample_1716 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.78
X1 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.78
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.78
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.78
X4 VTAIL.t6 VP.t1 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.78
X5 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.78
X6 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.78
X7 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.78
X8 VDD1.t1 VP.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.78
X9 VDD1.t0 VP.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.78
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.78
X11 VDD2.t0 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.78
R0 VP.n21 VP.n20 161.3
R1 VP.n19 VP.n1 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n16 VP.n2 161.3
R4 VP.n15 VP.n14 161.3
R5 VP.n13 VP.n3 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n4 161.3
R8 VP.n9 VP.n8 161.3
R9 VP.n5 VP.t1 159.225
R10 VP.n5 VP.t3 157.88
R11 VP.n7 VP.t0 125.409
R12 VP.n0 VP.t2 125.409
R13 VP.n7 VP.n6 87.376
R14 VP.n22 VP.n0 87.376
R15 VP.n6 VP.n5 57.6509
R16 VP.n14 VP.n13 40.4934
R17 VP.n14 VP.n2 40.4934
R18 VP.n8 VP.n4 24.4675
R19 VP.n12 VP.n4 24.4675
R20 VP.n13 VP.n12 24.4675
R21 VP.n18 VP.n2 24.4675
R22 VP.n19 VP.n18 24.4675
R23 VP.n20 VP.n19 24.4675
R24 VP.n8 VP.n7 2.69187
R25 VP.n20 VP.n0 2.69187
R26 VP.n9 VP.n6 0.354971
R27 VP.n22 VP.n21 0.354971
R28 VP VP.n22 0.26696
R29 VP.n10 VP.n9 0.189894
R30 VP.n11 VP.n10 0.189894
R31 VP.n11 VP.n3 0.189894
R32 VP.n15 VP.n3 0.189894
R33 VP.n16 VP.n15 0.189894
R34 VP.n17 VP.n16 0.189894
R35 VP.n17 VP.n1 0.189894
R36 VP.n21 VP.n1 0.189894
R37 VDD1 VDD1.n1 112.234
R38 VDD1 VDD1.n0 60.4662
R39 VDD1.n0 VDD1.t3 1.00711
R40 VDD1.n0 VDD1.t0 1.00711
R41 VDD1.n1 VDD1.t2 1.00711
R42 VDD1.n1 VDD1.t1 1.00711
R43 VTAIL.n874 VTAIL.n770 289.615
R44 VTAIL.n104 VTAIL.n0 289.615
R45 VTAIL.n214 VTAIL.n110 289.615
R46 VTAIL.n324 VTAIL.n220 289.615
R47 VTAIL.n764 VTAIL.n660 289.615
R48 VTAIL.n654 VTAIL.n550 289.615
R49 VTAIL.n544 VTAIL.n440 289.615
R50 VTAIL.n434 VTAIL.n330 289.615
R51 VTAIL.n807 VTAIL.n806 185
R52 VTAIL.n809 VTAIL.n808 185
R53 VTAIL.n802 VTAIL.n801 185
R54 VTAIL.n815 VTAIL.n814 185
R55 VTAIL.n817 VTAIL.n816 185
R56 VTAIL.n798 VTAIL.n797 185
R57 VTAIL.n823 VTAIL.n822 185
R58 VTAIL.n825 VTAIL.n824 185
R59 VTAIL.n794 VTAIL.n793 185
R60 VTAIL.n831 VTAIL.n830 185
R61 VTAIL.n833 VTAIL.n832 185
R62 VTAIL.n790 VTAIL.n789 185
R63 VTAIL.n839 VTAIL.n838 185
R64 VTAIL.n841 VTAIL.n840 185
R65 VTAIL.n786 VTAIL.n785 185
R66 VTAIL.n848 VTAIL.n847 185
R67 VTAIL.n849 VTAIL.n784 185
R68 VTAIL.n851 VTAIL.n850 185
R69 VTAIL.n782 VTAIL.n781 185
R70 VTAIL.n857 VTAIL.n856 185
R71 VTAIL.n859 VTAIL.n858 185
R72 VTAIL.n778 VTAIL.n777 185
R73 VTAIL.n865 VTAIL.n864 185
R74 VTAIL.n867 VTAIL.n866 185
R75 VTAIL.n774 VTAIL.n773 185
R76 VTAIL.n873 VTAIL.n872 185
R77 VTAIL.n875 VTAIL.n874 185
R78 VTAIL.n37 VTAIL.n36 185
R79 VTAIL.n39 VTAIL.n38 185
R80 VTAIL.n32 VTAIL.n31 185
R81 VTAIL.n45 VTAIL.n44 185
R82 VTAIL.n47 VTAIL.n46 185
R83 VTAIL.n28 VTAIL.n27 185
R84 VTAIL.n53 VTAIL.n52 185
R85 VTAIL.n55 VTAIL.n54 185
R86 VTAIL.n24 VTAIL.n23 185
R87 VTAIL.n61 VTAIL.n60 185
R88 VTAIL.n63 VTAIL.n62 185
R89 VTAIL.n20 VTAIL.n19 185
R90 VTAIL.n69 VTAIL.n68 185
R91 VTAIL.n71 VTAIL.n70 185
R92 VTAIL.n16 VTAIL.n15 185
R93 VTAIL.n78 VTAIL.n77 185
R94 VTAIL.n79 VTAIL.n14 185
R95 VTAIL.n81 VTAIL.n80 185
R96 VTAIL.n12 VTAIL.n11 185
R97 VTAIL.n87 VTAIL.n86 185
R98 VTAIL.n89 VTAIL.n88 185
R99 VTAIL.n8 VTAIL.n7 185
R100 VTAIL.n95 VTAIL.n94 185
R101 VTAIL.n97 VTAIL.n96 185
R102 VTAIL.n4 VTAIL.n3 185
R103 VTAIL.n103 VTAIL.n102 185
R104 VTAIL.n105 VTAIL.n104 185
R105 VTAIL.n147 VTAIL.n146 185
R106 VTAIL.n149 VTAIL.n148 185
R107 VTAIL.n142 VTAIL.n141 185
R108 VTAIL.n155 VTAIL.n154 185
R109 VTAIL.n157 VTAIL.n156 185
R110 VTAIL.n138 VTAIL.n137 185
R111 VTAIL.n163 VTAIL.n162 185
R112 VTAIL.n165 VTAIL.n164 185
R113 VTAIL.n134 VTAIL.n133 185
R114 VTAIL.n171 VTAIL.n170 185
R115 VTAIL.n173 VTAIL.n172 185
R116 VTAIL.n130 VTAIL.n129 185
R117 VTAIL.n179 VTAIL.n178 185
R118 VTAIL.n181 VTAIL.n180 185
R119 VTAIL.n126 VTAIL.n125 185
R120 VTAIL.n188 VTAIL.n187 185
R121 VTAIL.n189 VTAIL.n124 185
R122 VTAIL.n191 VTAIL.n190 185
R123 VTAIL.n122 VTAIL.n121 185
R124 VTAIL.n197 VTAIL.n196 185
R125 VTAIL.n199 VTAIL.n198 185
R126 VTAIL.n118 VTAIL.n117 185
R127 VTAIL.n205 VTAIL.n204 185
R128 VTAIL.n207 VTAIL.n206 185
R129 VTAIL.n114 VTAIL.n113 185
R130 VTAIL.n213 VTAIL.n212 185
R131 VTAIL.n215 VTAIL.n214 185
R132 VTAIL.n257 VTAIL.n256 185
R133 VTAIL.n259 VTAIL.n258 185
R134 VTAIL.n252 VTAIL.n251 185
R135 VTAIL.n265 VTAIL.n264 185
R136 VTAIL.n267 VTAIL.n266 185
R137 VTAIL.n248 VTAIL.n247 185
R138 VTAIL.n273 VTAIL.n272 185
R139 VTAIL.n275 VTAIL.n274 185
R140 VTAIL.n244 VTAIL.n243 185
R141 VTAIL.n281 VTAIL.n280 185
R142 VTAIL.n283 VTAIL.n282 185
R143 VTAIL.n240 VTAIL.n239 185
R144 VTAIL.n289 VTAIL.n288 185
R145 VTAIL.n291 VTAIL.n290 185
R146 VTAIL.n236 VTAIL.n235 185
R147 VTAIL.n298 VTAIL.n297 185
R148 VTAIL.n299 VTAIL.n234 185
R149 VTAIL.n301 VTAIL.n300 185
R150 VTAIL.n232 VTAIL.n231 185
R151 VTAIL.n307 VTAIL.n306 185
R152 VTAIL.n309 VTAIL.n308 185
R153 VTAIL.n228 VTAIL.n227 185
R154 VTAIL.n315 VTAIL.n314 185
R155 VTAIL.n317 VTAIL.n316 185
R156 VTAIL.n224 VTAIL.n223 185
R157 VTAIL.n323 VTAIL.n322 185
R158 VTAIL.n325 VTAIL.n324 185
R159 VTAIL.n765 VTAIL.n764 185
R160 VTAIL.n763 VTAIL.n762 185
R161 VTAIL.n664 VTAIL.n663 185
R162 VTAIL.n757 VTAIL.n756 185
R163 VTAIL.n755 VTAIL.n754 185
R164 VTAIL.n668 VTAIL.n667 185
R165 VTAIL.n749 VTAIL.n748 185
R166 VTAIL.n747 VTAIL.n746 185
R167 VTAIL.n672 VTAIL.n671 185
R168 VTAIL.n676 VTAIL.n674 185
R169 VTAIL.n741 VTAIL.n740 185
R170 VTAIL.n739 VTAIL.n738 185
R171 VTAIL.n678 VTAIL.n677 185
R172 VTAIL.n733 VTAIL.n732 185
R173 VTAIL.n731 VTAIL.n730 185
R174 VTAIL.n682 VTAIL.n681 185
R175 VTAIL.n725 VTAIL.n724 185
R176 VTAIL.n723 VTAIL.n722 185
R177 VTAIL.n686 VTAIL.n685 185
R178 VTAIL.n717 VTAIL.n716 185
R179 VTAIL.n715 VTAIL.n714 185
R180 VTAIL.n690 VTAIL.n689 185
R181 VTAIL.n709 VTAIL.n708 185
R182 VTAIL.n707 VTAIL.n706 185
R183 VTAIL.n694 VTAIL.n693 185
R184 VTAIL.n701 VTAIL.n700 185
R185 VTAIL.n699 VTAIL.n698 185
R186 VTAIL.n655 VTAIL.n654 185
R187 VTAIL.n653 VTAIL.n652 185
R188 VTAIL.n554 VTAIL.n553 185
R189 VTAIL.n647 VTAIL.n646 185
R190 VTAIL.n645 VTAIL.n644 185
R191 VTAIL.n558 VTAIL.n557 185
R192 VTAIL.n639 VTAIL.n638 185
R193 VTAIL.n637 VTAIL.n636 185
R194 VTAIL.n562 VTAIL.n561 185
R195 VTAIL.n566 VTAIL.n564 185
R196 VTAIL.n631 VTAIL.n630 185
R197 VTAIL.n629 VTAIL.n628 185
R198 VTAIL.n568 VTAIL.n567 185
R199 VTAIL.n623 VTAIL.n622 185
R200 VTAIL.n621 VTAIL.n620 185
R201 VTAIL.n572 VTAIL.n571 185
R202 VTAIL.n615 VTAIL.n614 185
R203 VTAIL.n613 VTAIL.n612 185
R204 VTAIL.n576 VTAIL.n575 185
R205 VTAIL.n607 VTAIL.n606 185
R206 VTAIL.n605 VTAIL.n604 185
R207 VTAIL.n580 VTAIL.n579 185
R208 VTAIL.n599 VTAIL.n598 185
R209 VTAIL.n597 VTAIL.n596 185
R210 VTAIL.n584 VTAIL.n583 185
R211 VTAIL.n591 VTAIL.n590 185
R212 VTAIL.n589 VTAIL.n588 185
R213 VTAIL.n545 VTAIL.n544 185
R214 VTAIL.n543 VTAIL.n542 185
R215 VTAIL.n444 VTAIL.n443 185
R216 VTAIL.n537 VTAIL.n536 185
R217 VTAIL.n535 VTAIL.n534 185
R218 VTAIL.n448 VTAIL.n447 185
R219 VTAIL.n529 VTAIL.n528 185
R220 VTAIL.n527 VTAIL.n526 185
R221 VTAIL.n452 VTAIL.n451 185
R222 VTAIL.n456 VTAIL.n454 185
R223 VTAIL.n521 VTAIL.n520 185
R224 VTAIL.n519 VTAIL.n518 185
R225 VTAIL.n458 VTAIL.n457 185
R226 VTAIL.n513 VTAIL.n512 185
R227 VTAIL.n511 VTAIL.n510 185
R228 VTAIL.n462 VTAIL.n461 185
R229 VTAIL.n505 VTAIL.n504 185
R230 VTAIL.n503 VTAIL.n502 185
R231 VTAIL.n466 VTAIL.n465 185
R232 VTAIL.n497 VTAIL.n496 185
R233 VTAIL.n495 VTAIL.n494 185
R234 VTAIL.n470 VTAIL.n469 185
R235 VTAIL.n489 VTAIL.n488 185
R236 VTAIL.n487 VTAIL.n486 185
R237 VTAIL.n474 VTAIL.n473 185
R238 VTAIL.n481 VTAIL.n480 185
R239 VTAIL.n479 VTAIL.n478 185
R240 VTAIL.n435 VTAIL.n434 185
R241 VTAIL.n433 VTAIL.n432 185
R242 VTAIL.n334 VTAIL.n333 185
R243 VTAIL.n427 VTAIL.n426 185
R244 VTAIL.n425 VTAIL.n424 185
R245 VTAIL.n338 VTAIL.n337 185
R246 VTAIL.n419 VTAIL.n418 185
R247 VTAIL.n417 VTAIL.n416 185
R248 VTAIL.n342 VTAIL.n341 185
R249 VTAIL.n346 VTAIL.n344 185
R250 VTAIL.n411 VTAIL.n410 185
R251 VTAIL.n409 VTAIL.n408 185
R252 VTAIL.n348 VTAIL.n347 185
R253 VTAIL.n403 VTAIL.n402 185
R254 VTAIL.n401 VTAIL.n400 185
R255 VTAIL.n352 VTAIL.n351 185
R256 VTAIL.n395 VTAIL.n394 185
R257 VTAIL.n393 VTAIL.n392 185
R258 VTAIL.n356 VTAIL.n355 185
R259 VTAIL.n387 VTAIL.n386 185
R260 VTAIL.n385 VTAIL.n384 185
R261 VTAIL.n360 VTAIL.n359 185
R262 VTAIL.n379 VTAIL.n378 185
R263 VTAIL.n377 VTAIL.n376 185
R264 VTAIL.n364 VTAIL.n363 185
R265 VTAIL.n371 VTAIL.n370 185
R266 VTAIL.n369 VTAIL.n368 185
R267 VTAIL.n805 VTAIL.t0 147.659
R268 VTAIL.n35 VTAIL.t2 147.659
R269 VTAIL.n145 VTAIL.t5 147.659
R270 VTAIL.n255 VTAIL.t7 147.659
R271 VTAIL.n697 VTAIL.t4 147.659
R272 VTAIL.n587 VTAIL.t6 147.659
R273 VTAIL.n477 VTAIL.t3 147.659
R274 VTAIL.n367 VTAIL.t1 147.659
R275 VTAIL.n808 VTAIL.n807 104.615
R276 VTAIL.n808 VTAIL.n801 104.615
R277 VTAIL.n815 VTAIL.n801 104.615
R278 VTAIL.n816 VTAIL.n815 104.615
R279 VTAIL.n816 VTAIL.n797 104.615
R280 VTAIL.n823 VTAIL.n797 104.615
R281 VTAIL.n824 VTAIL.n823 104.615
R282 VTAIL.n824 VTAIL.n793 104.615
R283 VTAIL.n831 VTAIL.n793 104.615
R284 VTAIL.n832 VTAIL.n831 104.615
R285 VTAIL.n832 VTAIL.n789 104.615
R286 VTAIL.n839 VTAIL.n789 104.615
R287 VTAIL.n840 VTAIL.n839 104.615
R288 VTAIL.n840 VTAIL.n785 104.615
R289 VTAIL.n848 VTAIL.n785 104.615
R290 VTAIL.n849 VTAIL.n848 104.615
R291 VTAIL.n850 VTAIL.n849 104.615
R292 VTAIL.n850 VTAIL.n781 104.615
R293 VTAIL.n857 VTAIL.n781 104.615
R294 VTAIL.n858 VTAIL.n857 104.615
R295 VTAIL.n858 VTAIL.n777 104.615
R296 VTAIL.n865 VTAIL.n777 104.615
R297 VTAIL.n866 VTAIL.n865 104.615
R298 VTAIL.n866 VTAIL.n773 104.615
R299 VTAIL.n873 VTAIL.n773 104.615
R300 VTAIL.n874 VTAIL.n873 104.615
R301 VTAIL.n38 VTAIL.n37 104.615
R302 VTAIL.n38 VTAIL.n31 104.615
R303 VTAIL.n45 VTAIL.n31 104.615
R304 VTAIL.n46 VTAIL.n45 104.615
R305 VTAIL.n46 VTAIL.n27 104.615
R306 VTAIL.n53 VTAIL.n27 104.615
R307 VTAIL.n54 VTAIL.n53 104.615
R308 VTAIL.n54 VTAIL.n23 104.615
R309 VTAIL.n61 VTAIL.n23 104.615
R310 VTAIL.n62 VTAIL.n61 104.615
R311 VTAIL.n62 VTAIL.n19 104.615
R312 VTAIL.n69 VTAIL.n19 104.615
R313 VTAIL.n70 VTAIL.n69 104.615
R314 VTAIL.n70 VTAIL.n15 104.615
R315 VTAIL.n78 VTAIL.n15 104.615
R316 VTAIL.n79 VTAIL.n78 104.615
R317 VTAIL.n80 VTAIL.n79 104.615
R318 VTAIL.n80 VTAIL.n11 104.615
R319 VTAIL.n87 VTAIL.n11 104.615
R320 VTAIL.n88 VTAIL.n87 104.615
R321 VTAIL.n88 VTAIL.n7 104.615
R322 VTAIL.n95 VTAIL.n7 104.615
R323 VTAIL.n96 VTAIL.n95 104.615
R324 VTAIL.n96 VTAIL.n3 104.615
R325 VTAIL.n103 VTAIL.n3 104.615
R326 VTAIL.n104 VTAIL.n103 104.615
R327 VTAIL.n148 VTAIL.n147 104.615
R328 VTAIL.n148 VTAIL.n141 104.615
R329 VTAIL.n155 VTAIL.n141 104.615
R330 VTAIL.n156 VTAIL.n155 104.615
R331 VTAIL.n156 VTAIL.n137 104.615
R332 VTAIL.n163 VTAIL.n137 104.615
R333 VTAIL.n164 VTAIL.n163 104.615
R334 VTAIL.n164 VTAIL.n133 104.615
R335 VTAIL.n171 VTAIL.n133 104.615
R336 VTAIL.n172 VTAIL.n171 104.615
R337 VTAIL.n172 VTAIL.n129 104.615
R338 VTAIL.n179 VTAIL.n129 104.615
R339 VTAIL.n180 VTAIL.n179 104.615
R340 VTAIL.n180 VTAIL.n125 104.615
R341 VTAIL.n188 VTAIL.n125 104.615
R342 VTAIL.n189 VTAIL.n188 104.615
R343 VTAIL.n190 VTAIL.n189 104.615
R344 VTAIL.n190 VTAIL.n121 104.615
R345 VTAIL.n197 VTAIL.n121 104.615
R346 VTAIL.n198 VTAIL.n197 104.615
R347 VTAIL.n198 VTAIL.n117 104.615
R348 VTAIL.n205 VTAIL.n117 104.615
R349 VTAIL.n206 VTAIL.n205 104.615
R350 VTAIL.n206 VTAIL.n113 104.615
R351 VTAIL.n213 VTAIL.n113 104.615
R352 VTAIL.n214 VTAIL.n213 104.615
R353 VTAIL.n258 VTAIL.n257 104.615
R354 VTAIL.n258 VTAIL.n251 104.615
R355 VTAIL.n265 VTAIL.n251 104.615
R356 VTAIL.n266 VTAIL.n265 104.615
R357 VTAIL.n266 VTAIL.n247 104.615
R358 VTAIL.n273 VTAIL.n247 104.615
R359 VTAIL.n274 VTAIL.n273 104.615
R360 VTAIL.n274 VTAIL.n243 104.615
R361 VTAIL.n281 VTAIL.n243 104.615
R362 VTAIL.n282 VTAIL.n281 104.615
R363 VTAIL.n282 VTAIL.n239 104.615
R364 VTAIL.n289 VTAIL.n239 104.615
R365 VTAIL.n290 VTAIL.n289 104.615
R366 VTAIL.n290 VTAIL.n235 104.615
R367 VTAIL.n298 VTAIL.n235 104.615
R368 VTAIL.n299 VTAIL.n298 104.615
R369 VTAIL.n300 VTAIL.n299 104.615
R370 VTAIL.n300 VTAIL.n231 104.615
R371 VTAIL.n307 VTAIL.n231 104.615
R372 VTAIL.n308 VTAIL.n307 104.615
R373 VTAIL.n308 VTAIL.n227 104.615
R374 VTAIL.n315 VTAIL.n227 104.615
R375 VTAIL.n316 VTAIL.n315 104.615
R376 VTAIL.n316 VTAIL.n223 104.615
R377 VTAIL.n323 VTAIL.n223 104.615
R378 VTAIL.n324 VTAIL.n323 104.615
R379 VTAIL.n764 VTAIL.n763 104.615
R380 VTAIL.n763 VTAIL.n663 104.615
R381 VTAIL.n756 VTAIL.n663 104.615
R382 VTAIL.n756 VTAIL.n755 104.615
R383 VTAIL.n755 VTAIL.n667 104.615
R384 VTAIL.n748 VTAIL.n667 104.615
R385 VTAIL.n748 VTAIL.n747 104.615
R386 VTAIL.n747 VTAIL.n671 104.615
R387 VTAIL.n676 VTAIL.n671 104.615
R388 VTAIL.n740 VTAIL.n676 104.615
R389 VTAIL.n740 VTAIL.n739 104.615
R390 VTAIL.n739 VTAIL.n677 104.615
R391 VTAIL.n732 VTAIL.n677 104.615
R392 VTAIL.n732 VTAIL.n731 104.615
R393 VTAIL.n731 VTAIL.n681 104.615
R394 VTAIL.n724 VTAIL.n681 104.615
R395 VTAIL.n724 VTAIL.n723 104.615
R396 VTAIL.n723 VTAIL.n685 104.615
R397 VTAIL.n716 VTAIL.n685 104.615
R398 VTAIL.n716 VTAIL.n715 104.615
R399 VTAIL.n715 VTAIL.n689 104.615
R400 VTAIL.n708 VTAIL.n689 104.615
R401 VTAIL.n708 VTAIL.n707 104.615
R402 VTAIL.n707 VTAIL.n693 104.615
R403 VTAIL.n700 VTAIL.n693 104.615
R404 VTAIL.n700 VTAIL.n699 104.615
R405 VTAIL.n654 VTAIL.n653 104.615
R406 VTAIL.n653 VTAIL.n553 104.615
R407 VTAIL.n646 VTAIL.n553 104.615
R408 VTAIL.n646 VTAIL.n645 104.615
R409 VTAIL.n645 VTAIL.n557 104.615
R410 VTAIL.n638 VTAIL.n557 104.615
R411 VTAIL.n638 VTAIL.n637 104.615
R412 VTAIL.n637 VTAIL.n561 104.615
R413 VTAIL.n566 VTAIL.n561 104.615
R414 VTAIL.n630 VTAIL.n566 104.615
R415 VTAIL.n630 VTAIL.n629 104.615
R416 VTAIL.n629 VTAIL.n567 104.615
R417 VTAIL.n622 VTAIL.n567 104.615
R418 VTAIL.n622 VTAIL.n621 104.615
R419 VTAIL.n621 VTAIL.n571 104.615
R420 VTAIL.n614 VTAIL.n571 104.615
R421 VTAIL.n614 VTAIL.n613 104.615
R422 VTAIL.n613 VTAIL.n575 104.615
R423 VTAIL.n606 VTAIL.n575 104.615
R424 VTAIL.n606 VTAIL.n605 104.615
R425 VTAIL.n605 VTAIL.n579 104.615
R426 VTAIL.n598 VTAIL.n579 104.615
R427 VTAIL.n598 VTAIL.n597 104.615
R428 VTAIL.n597 VTAIL.n583 104.615
R429 VTAIL.n590 VTAIL.n583 104.615
R430 VTAIL.n590 VTAIL.n589 104.615
R431 VTAIL.n544 VTAIL.n543 104.615
R432 VTAIL.n543 VTAIL.n443 104.615
R433 VTAIL.n536 VTAIL.n443 104.615
R434 VTAIL.n536 VTAIL.n535 104.615
R435 VTAIL.n535 VTAIL.n447 104.615
R436 VTAIL.n528 VTAIL.n447 104.615
R437 VTAIL.n528 VTAIL.n527 104.615
R438 VTAIL.n527 VTAIL.n451 104.615
R439 VTAIL.n456 VTAIL.n451 104.615
R440 VTAIL.n520 VTAIL.n456 104.615
R441 VTAIL.n520 VTAIL.n519 104.615
R442 VTAIL.n519 VTAIL.n457 104.615
R443 VTAIL.n512 VTAIL.n457 104.615
R444 VTAIL.n512 VTAIL.n511 104.615
R445 VTAIL.n511 VTAIL.n461 104.615
R446 VTAIL.n504 VTAIL.n461 104.615
R447 VTAIL.n504 VTAIL.n503 104.615
R448 VTAIL.n503 VTAIL.n465 104.615
R449 VTAIL.n496 VTAIL.n465 104.615
R450 VTAIL.n496 VTAIL.n495 104.615
R451 VTAIL.n495 VTAIL.n469 104.615
R452 VTAIL.n488 VTAIL.n469 104.615
R453 VTAIL.n488 VTAIL.n487 104.615
R454 VTAIL.n487 VTAIL.n473 104.615
R455 VTAIL.n480 VTAIL.n473 104.615
R456 VTAIL.n480 VTAIL.n479 104.615
R457 VTAIL.n434 VTAIL.n433 104.615
R458 VTAIL.n433 VTAIL.n333 104.615
R459 VTAIL.n426 VTAIL.n333 104.615
R460 VTAIL.n426 VTAIL.n425 104.615
R461 VTAIL.n425 VTAIL.n337 104.615
R462 VTAIL.n418 VTAIL.n337 104.615
R463 VTAIL.n418 VTAIL.n417 104.615
R464 VTAIL.n417 VTAIL.n341 104.615
R465 VTAIL.n346 VTAIL.n341 104.615
R466 VTAIL.n410 VTAIL.n346 104.615
R467 VTAIL.n410 VTAIL.n409 104.615
R468 VTAIL.n409 VTAIL.n347 104.615
R469 VTAIL.n402 VTAIL.n347 104.615
R470 VTAIL.n402 VTAIL.n401 104.615
R471 VTAIL.n401 VTAIL.n351 104.615
R472 VTAIL.n394 VTAIL.n351 104.615
R473 VTAIL.n394 VTAIL.n393 104.615
R474 VTAIL.n393 VTAIL.n355 104.615
R475 VTAIL.n386 VTAIL.n355 104.615
R476 VTAIL.n386 VTAIL.n385 104.615
R477 VTAIL.n385 VTAIL.n359 104.615
R478 VTAIL.n378 VTAIL.n359 104.615
R479 VTAIL.n378 VTAIL.n377 104.615
R480 VTAIL.n377 VTAIL.n363 104.615
R481 VTAIL.n370 VTAIL.n363 104.615
R482 VTAIL.n370 VTAIL.n369 104.615
R483 VTAIL.n807 VTAIL.t0 52.3082
R484 VTAIL.n37 VTAIL.t2 52.3082
R485 VTAIL.n147 VTAIL.t5 52.3082
R486 VTAIL.n257 VTAIL.t7 52.3082
R487 VTAIL.n699 VTAIL.t4 52.3082
R488 VTAIL.n589 VTAIL.t6 52.3082
R489 VTAIL.n479 VTAIL.t3 52.3082
R490 VTAIL.n369 VTAIL.t1 52.3082
R491 VTAIL.n879 VTAIL.n769 32.8669
R492 VTAIL.n439 VTAIL.n329 32.8669
R493 VTAIL.n879 VTAIL.n878 31.9914
R494 VTAIL.n109 VTAIL.n108 31.9914
R495 VTAIL.n219 VTAIL.n218 31.9914
R496 VTAIL.n329 VTAIL.n328 31.9914
R497 VTAIL.n769 VTAIL.n768 31.9914
R498 VTAIL.n659 VTAIL.n658 31.9914
R499 VTAIL.n549 VTAIL.n548 31.9914
R500 VTAIL.n439 VTAIL.n438 31.9914
R501 VTAIL.n806 VTAIL.n805 15.6677
R502 VTAIL.n36 VTAIL.n35 15.6677
R503 VTAIL.n146 VTAIL.n145 15.6677
R504 VTAIL.n256 VTAIL.n255 15.6677
R505 VTAIL.n698 VTAIL.n697 15.6677
R506 VTAIL.n588 VTAIL.n587 15.6677
R507 VTAIL.n478 VTAIL.n477 15.6677
R508 VTAIL.n368 VTAIL.n367 15.6677
R509 VTAIL.n851 VTAIL.n782 13.1884
R510 VTAIL.n81 VTAIL.n12 13.1884
R511 VTAIL.n191 VTAIL.n122 13.1884
R512 VTAIL.n301 VTAIL.n232 13.1884
R513 VTAIL.n674 VTAIL.n672 13.1884
R514 VTAIL.n564 VTAIL.n562 13.1884
R515 VTAIL.n454 VTAIL.n452 13.1884
R516 VTAIL.n344 VTAIL.n342 13.1884
R517 VTAIL.n809 VTAIL.n804 12.8005
R518 VTAIL.n852 VTAIL.n784 12.8005
R519 VTAIL.n856 VTAIL.n855 12.8005
R520 VTAIL.n39 VTAIL.n34 12.8005
R521 VTAIL.n82 VTAIL.n14 12.8005
R522 VTAIL.n86 VTAIL.n85 12.8005
R523 VTAIL.n149 VTAIL.n144 12.8005
R524 VTAIL.n192 VTAIL.n124 12.8005
R525 VTAIL.n196 VTAIL.n195 12.8005
R526 VTAIL.n259 VTAIL.n254 12.8005
R527 VTAIL.n302 VTAIL.n234 12.8005
R528 VTAIL.n306 VTAIL.n305 12.8005
R529 VTAIL.n746 VTAIL.n745 12.8005
R530 VTAIL.n742 VTAIL.n741 12.8005
R531 VTAIL.n701 VTAIL.n696 12.8005
R532 VTAIL.n636 VTAIL.n635 12.8005
R533 VTAIL.n632 VTAIL.n631 12.8005
R534 VTAIL.n591 VTAIL.n586 12.8005
R535 VTAIL.n526 VTAIL.n525 12.8005
R536 VTAIL.n522 VTAIL.n521 12.8005
R537 VTAIL.n481 VTAIL.n476 12.8005
R538 VTAIL.n416 VTAIL.n415 12.8005
R539 VTAIL.n412 VTAIL.n411 12.8005
R540 VTAIL.n371 VTAIL.n366 12.8005
R541 VTAIL.n810 VTAIL.n802 12.0247
R542 VTAIL.n847 VTAIL.n846 12.0247
R543 VTAIL.n859 VTAIL.n780 12.0247
R544 VTAIL.n40 VTAIL.n32 12.0247
R545 VTAIL.n77 VTAIL.n76 12.0247
R546 VTAIL.n89 VTAIL.n10 12.0247
R547 VTAIL.n150 VTAIL.n142 12.0247
R548 VTAIL.n187 VTAIL.n186 12.0247
R549 VTAIL.n199 VTAIL.n120 12.0247
R550 VTAIL.n260 VTAIL.n252 12.0247
R551 VTAIL.n297 VTAIL.n296 12.0247
R552 VTAIL.n309 VTAIL.n230 12.0247
R553 VTAIL.n749 VTAIL.n670 12.0247
R554 VTAIL.n738 VTAIL.n675 12.0247
R555 VTAIL.n702 VTAIL.n694 12.0247
R556 VTAIL.n639 VTAIL.n560 12.0247
R557 VTAIL.n628 VTAIL.n565 12.0247
R558 VTAIL.n592 VTAIL.n584 12.0247
R559 VTAIL.n529 VTAIL.n450 12.0247
R560 VTAIL.n518 VTAIL.n455 12.0247
R561 VTAIL.n482 VTAIL.n474 12.0247
R562 VTAIL.n419 VTAIL.n340 12.0247
R563 VTAIL.n408 VTAIL.n345 12.0247
R564 VTAIL.n372 VTAIL.n364 12.0247
R565 VTAIL.n814 VTAIL.n813 11.249
R566 VTAIL.n845 VTAIL.n786 11.249
R567 VTAIL.n860 VTAIL.n778 11.249
R568 VTAIL.n44 VTAIL.n43 11.249
R569 VTAIL.n75 VTAIL.n16 11.249
R570 VTAIL.n90 VTAIL.n8 11.249
R571 VTAIL.n154 VTAIL.n153 11.249
R572 VTAIL.n185 VTAIL.n126 11.249
R573 VTAIL.n200 VTAIL.n118 11.249
R574 VTAIL.n264 VTAIL.n263 11.249
R575 VTAIL.n295 VTAIL.n236 11.249
R576 VTAIL.n310 VTAIL.n228 11.249
R577 VTAIL.n750 VTAIL.n668 11.249
R578 VTAIL.n737 VTAIL.n678 11.249
R579 VTAIL.n706 VTAIL.n705 11.249
R580 VTAIL.n640 VTAIL.n558 11.249
R581 VTAIL.n627 VTAIL.n568 11.249
R582 VTAIL.n596 VTAIL.n595 11.249
R583 VTAIL.n530 VTAIL.n448 11.249
R584 VTAIL.n517 VTAIL.n458 11.249
R585 VTAIL.n486 VTAIL.n485 11.249
R586 VTAIL.n420 VTAIL.n338 11.249
R587 VTAIL.n407 VTAIL.n348 11.249
R588 VTAIL.n376 VTAIL.n375 11.249
R589 VTAIL.n817 VTAIL.n800 10.4732
R590 VTAIL.n842 VTAIL.n841 10.4732
R591 VTAIL.n864 VTAIL.n863 10.4732
R592 VTAIL.n47 VTAIL.n30 10.4732
R593 VTAIL.n72 VTAIL.n71 10.4732
R594 VTAIL.n94 VTAIL.n93 10.4732
R595 VTAIL.n157 VTAIL.n140 10.4732
R596 VTAIL.n182 VTAIL.n181 10.4732
R597 VTAIL.n204 VTAIL.n203 10.4732
R598 VTAIL.n267 VTAIL.n250 10.4732
R599 VTAIL.n292 VTAIL.n291 10.4732
R600 VTAIL.n314 VTAIL.n313 10.4732
R601 VTAIL.n754 VTAIL.n753 10.4732
R602 VTAIL.n734 VTAIL.n733 10.4732
R603 VTAIL.n709 VTAIL.n692 10.4732
R604 VTAIL.n644 VTAIL.n643 10.4732
R605 VTAIL.n624 VTAIL.n623 10.4732
R606 VTAIL.n599 VTAIL.n582 10.4732
R607 VTAIL.n534 VTAIL.n533 10.4732
R608 VTAIL.n514 VTAIL.n513 10.4732
R609 VTAIL.n489 VTAIL.n472 10.4732
R610 VTAIL.n424 VTAIL.n423 10.4732
R611 VTAIL.n404 VTAIL.n403 10.4732
R612 VTAIL.n379 VTAIL.n362 10.4732
R613 VTAIL.n818 VTAIL.n798 9.69747
R614 VTAIL.n838 VTAIL.n788 9.69747
R615 VTAIL.n867 VTAIL.n776 9.69747
R616 VTAIL.n48 VTAIL.n28 9.69747
R617 VTAIL.n68 VTAIL.n18 9.69747
R618 VTAIL.n97 VTAIL.n6 9.69747
R619 VTAIL.n158 VTAIL.n138 9.69747
R620 VTAIL.n178 VTAIL.n128 9.69747
R621 VTAIL.n207 VTAIL.n116 9.69747
R622 VTAIL.n268 VTAIL.n248 9.69747
R623 VTAIL.n288 VTAIL.n238 9.69747
R624 VTAIL.n317 VTAIL.n226 9.69747
R625 VTAIL.n757 VTAIL.n666 9.69747
R626 VTAIL.n730 VTAIL.n680 9.69747
R627 VTAIL.n710 VTAIL.n690 9.69747
R628 VTAIL.n647 VTAIL.n556 9.69747
R629 VTAIL.n620 VTAIL.n570 9.69747
R630 VTAIL.n600 VTAIL.n580 9.69747
R631 VTAIL.n537 VTAIL.n446 9.69747
R632 VTAIL.n510 VTAIL.n460 9.69747
R633 VTAIL.n490 VTAIL.n470 9.69747
R634 VTAIL.n427 VTAIL.n336 9.69747
R635 VTAIL.n400 VTAIL.n350 9.69747
R636 VTAIL.n380 VTAIL.n360 9.69747
R637 VTAIL.n878 VTAIL.n877 9.45567
R638 VTAIL.n108 VTAIL.n107 9.45567
R639 VTAIL.n218 VTAIL.n217 9.45567
R640 VTAIL.n328 VTAIL.n327 9.45567
R641 VTAIL.n768 VTAIL.n767 9.45567
R642 VTAIL.n658 VTAIL.n657 9.45567
R643 VTAIL.n548 VTAIL.n547 9.45567
R644 VTAIL.n438 VTAIL.n437 9.45567
R645 VTAIL.n877 VTAIL.n876 9.3005
R646 VTAIL.n871 VTAIL.n870 9.3005
R647 VTAIL.n869 VTAIL.n868 9.3005
R648 VTAIL.n776 VTAIL.n775 9.3005
R649 VTAIL.n863 VTAIL.n862 9.3005
R650 VTAIL.n861 VTAIL.n860 9.3005
R651 VTAIL.n780 VTAIL.n779 9.3005
R652 VTAIL.n855 VTAIL.n854 9.3005
R653 VTAIL.n827 VTAIL.n826 9.3005
R654 VTAIL.n796 VTAIL.n795 9.3005
R655 VTAIL.n821 VTAIL.n820 9.3005
R656 VTAIL.n819 VTAIL.n818 9.3005
R657 VTAIL.n800 VTAIL.n799 9.3005
R658 VTAIL.n813 VTAIL.n812 9.3005
R659 VTAIL.n811 VTAIL.n810 9.3005
R660 VTAIL.n804 VTAIL.n803 9.3005
R661 VTAIL.n829 VTAIL.n828 9.3005
R662 VTAIL.n792 VTAIL.n791 9.3005
R663 VTAIL.n835 VTAIL.n834 9.3005
R664 VTAIL.n837 VTAIL.n836 9.3005
R665 VTAIL.n788 VTAIL.n787 9.3005
R666 VTAIL.n843 VTAIL.n842 9.3005
R667 VTAIL.n845 VTAIL.n844 9.3005
R668 VTAIL.n846 VTAIL.n783 9.3005
R669 VTAIL.n853 VTAIL.n852 9.3005
R670 VTAIL.n772 VTAIL.n771 9.3005
R671 VTAIL.n107 VTAIL.n106 9.3005
R672 VTAIL.n101 VTAIL.n100 9.3005
R673 VTAIL.n99 VTAIL.n98 9.3005
R674 VTAIL.n6 VTAIL.n5 9.3005
R675 VTAIL.n93 VTAIL.n92 9.3005
R676 VTAIL.n91 VTAIL.n90 9.3005
R677 VTAIL.n10 VTAIL.n9 9.3005
R678 VTAIL.n85 VTAIL.n84 9.3005
R679 VTAIL.n57 VTAIL.n56 9.3005
R680 VTAIL.n26 VTAIL.n25 9.3005
R681 VTAIL.n51 VTAIL.n50 9.3005
R682 VTAIL.n49 VTAIL.n48 9.3005
R683 VTAIL.n30 VTAIL.n29 9.3005
R684 VTAIL.n43 VTAIL.n42 9.3005
R685 VTAIL.n41 VTAIL.n40 9.3005
R686 VTAIL.n34 VTAIL.n33 9.3005
R687 VTAIL.n59 VTAIL.n58 9.3005
R688 VTAIL.n22 VTAIL.n21 9.3005
R689 VTAIL.n65 VTAIL.n64 9.3005
R690 VTAIL.n67 VTAIL.n66 9.3005
R691 VTAIL.n18 VTAIL.n17 9.3005
R692 VTAIL.n73 VTAIL.n72 9.3005
R693 VTAIL.n75 VTAIL.n74 9.3005
R694 VTAIL.n76 VTAIL.n13 9.3005
R695 VTAIL.n83 VTAIL.n82 9.3005
R696 VTAIL.n2 VTAIL.n1 9.3005
R697 VTAIL.n217 VTAIL.n216 9.3005
R698 VTAIL.n211 VTAIL.n210 9.3005
R699 VTAIL.n209 VTAIL.n208 9.3005
R700 VTAIL.n116 VTAIL.n115 9.3005
R701 VTAIL.n203 VTAIL.n202 9.3005
R702 VTAIL.n201 VTAIL.n200 9.3005
R703 VTAIL.n120 VTAIL.n119 9.3005
R704 VTAIL.n195 VTAIL.n194 9.3005
R705 VTAIL.n167 VTAIL.n166 9.3005
R706 VTAIL.n136 VTAIL.n135 9.3005
R707 VTAIL.n161 VTAIL.n160 9.3005
R708 VTAIL.n159 VTAIL.n158 9.3005
R709 VTAIL.n140 VTAIL.n139 9.3005
R710 VTAIL.n153 VTAIL.n152 9.3005
R711 VTAIL.n151 VTAIL.n150 9.3005
R712 VTAIL.n144 VTAIL.n143 9.3005
R713 VTAIL.n169 VTAIL.n168 9.3005
R714 VTAIL.n132 VTAIL.n131 9.3005
R715 VTAIL.n175 VTAIL.n174 9.3005
R716 VTAIL.n177 VTAIL.n176 9.3005
R717 VTAIL.n128 VTAIL.n127 9.3005
R718 VTAIL.n183 VTAIL.n182 9.3005
R719 VTAIL.n185 VTAIL.n184 9.3005
R720 VTAIL.n186 VTAIL.n123 9.3005
R721 VTAIL.n193 VTAIL.n192 9.3005
R722 VTAIL.n112 VTAIL.n111 9.3005
R723 VTAIL.n327 VTAIL.n326 9.3005
R724 VTAIL.n321 VTAIL.n320 9.3005
R725 VTAIL.n319 VTAIL.n318 9.3005
R726 VTAIL.n226 VTAIL.n225 9.3005
R727 VTAIL.n313 VTAIL.n312 9.3005
R728 VTAIL.n311 VTAIL.n310 9.3005
R729 VTAIL.n230 VTAIL.n229 9.3005
R730 VTAIL.n305 VTAIL.n304 9.3005
R731 VTAIL.n277 VTAIL.n276 9.3005
R732 VTAIL.n246 VTAIL.n245 9.3005
R733 VTAIL.n271 VTAIL.n270 9.3005
R734 VTAIL.n269 VTAIL.n268 9.3005
R735 VTAIL.n250 VTAIL.n249 9.3005
R736 VTAIL.n263 VTAIL.n262 9.3005
R737 VTAIL.n261 VTAIL.n260 9.3005
R738 VTAIL.n254 VTAIL.n253 9.3005
R739 VTAIL.n279 VTAIL.n278 9.3005
R740 VTAIL.n242 VTAIL.n241 9.3005
R741 VTAIL.n285 VTAIL.n284 9.3005
R742 VTAIL.n287 VTAIL.n286 9.3005
R743 VTAIL.n238 VTAIL.n237 9.3005
R744 VTAIL.n293 VTAIL.n292 9.3005
R745 VTAIL.n295 VTAIL.n294 9.3005
R746 VTAIL.n296 VTAIL.n233 9.3005
R747 VTAIL.n303 VTAIL.n302 9.3005
R748 VTAIL.n222 VTAIL.n221 9.3005
R749 VTAIL.n684 VTAIL.n683 9.3005
R750 VTAIL.n727 VTAIL.n726 9.3005
R751 VTAIL.n729 VTAIL.n728 9.3005
R752 VTAIL.n680 VTAIL.n679 9.3005
R753 VTAIL.n735 VTAIL.n734 9.3005
R754 VTAIL.n737 VTAIL.n736 9.3005
R755 VTAIL.n675 VTAIL.n673 9.3005
R756 VTAIL.n743 VTAIL.n742 9.3005
R757 VTAIL.n767 VTAIL.n766 9.3005
R758 VTAIL.n662 VTAIL.n661 9.3005
R759 VTAIL.n761 VTAIL.n760 9.3005
R760 VTAIL.n759 VTAIL.n758 9.3005
R761 VTAIL.n666 VTAIL.n665 9.3005
R762 VTAIL.n753 VTAIL.n752 9.3005
R763 VTAIL.n751 VTAIL.n750 9.3005
R764 VTAIL.n670 VTAIL.n669 9.3005
R765 VTAIL.n745 VTAIL.n744 9.3005
R766 VTAIL.n721 VTAIL.n720 9.3005
R767 VTAIL.n719 VTAIL.n718 9.3005
R768 VTAIL.n688 VTAIL.n687 9.3005
R769 VTAIL.n713 VTAIL.n712 9.3005
R770 VTAIL.n711 VTAIL.n710 9.3005
R771 VTAIL.n692 VTAIL.n691 9.3005
R772 VTAIL.n705 VTAIL.n704 9.3005
R773 VTAIL.n703 VTAIL.n702 9.3005
R774 VTAIL.n696 VTAIL.n695 9.3005
R775 VTAIL.n574 VTAIL.n573 9.3005
R776 VTAIL.n617 VTAIL.n616 9.3005
R777 VTAIL.n619 VTAIL.n618 9.3005
R778 VTAIL.n570 VTAIL.n569 9.3005
R779 VTAIL.n625 VTAIL.n624 9.3005
R780 VTAIL.n627 VTAIL.n626 9.3005
R781 VTAIL.n565 VTAIL.n563 9.3005
R782 VTAIL.n633 VTAIL.n632 9.3005
R783 VTAIL.n657 VTAIL.n656 9.3005
R784 VTAIL.n552 VTAIL.n551 9.3005
R785 VTAIL.n651 VTAIL.n650 9.3005
R786 VTAIL.n649 VTAIL.n648 9.3005
R787 VTAIL.n556 VTAIL.n555 9.3005
R788 VTAIL.n643 VTAIL.n642 9.3005
R789 VTAIL.n641 VTAIL.n640 9.3005
R790 VTAIL.n560 VTAIL.n559 9.3005
R791 VTAIL.n635 VTAIL.n634 9.3005
R792 VTAIL.n611 VTAIL.n610 9.3005
R793 VTAIL.n609 VTAIL.n608 9.3005
R794 VTAIL.n578 VTAIL.n577 9.3005
R795 VTAIL.n603 VTAIL.n602 9.3005
R796 VTAIL.n601 VTAIL.n600 9.3005
R797 VTAIL.n582 VTAIL.n581 9.3005
R798 VTAIL.n595 VTAIL.n594 9.3005
R799 VTAIL.n593 VTAIL.n592 9.3005
R800 VTAIL.n586 VTAIL.n585 9.3005
R801 VTAIL.n464 VTAIL.n463 9.3005
R802 VTAIL.n507 VTAIL.n506 9.3005
R803 VTAIL.n509 VTAIL.n508 9.3005
R804 VTAIL.n460 VTAIL.n459 9.3005
R805 VTAIL.n515 VTAIL.n514 9.3005
R806 VTAIL.n517 VTAIL.n516 9.3005
R807 VTAIL.n455 VTAIL.n453 9.3005
R808 VTAIL.n523 VTAIL.n522 9.3005
R809 VTAIL.n547 VTAIL.n546 9.3005
R810 VTAIL.n442 VTAIL.n441 9.3005
R811 VTAIL.n541 VTAIL.n540 9.3005
R812 VTAIL.n539 VTAIL.n538 9.3005
R813 VTAIL.n446 VTAIL.n445 9.3005
R814 VTAIL.n533 VTAIL.n532 9.3005
R815 VTAIL.n531 VTAIL.n530 9.3005
R816 VTAIL.n450 VTAIL.n449 9.3005
R817 VTAIL.n525 VTAIL.n524 9.3005
R818 VTAIL.n501 VTAIL.n500 9.3005
R819 VTAIL.n499 VTAIL.n498 9.3005
R820 VTAIL.n468 VTAIL.n467 9.3005
R821 VTAIL.n493 VTAIL.n492 9.3005
R822 VTAIL.n491 VTAIL.n490 9.3005
R823 VTAIL.n472 VTAIL.n471 9.3005
R824 VTAIL.n485 VTAIL.n484 9.3005
R825 VTAIL.n483 VTAIL.n482 9.3005
R826 VTAIL.n476 VTAIL.n475 9.3005
R827 VTAIL.n354 VTAIL.n353 9.3005
R828 VTAIL.n397 VTAIL.n396 9.3005
R829 VTAIL.n399 VTAIL.n398 9.3005
R830 VTAIL.n350 VTAIL.n349 9.3005
R831 VTAIL.n405 VTAIL.n404 9.3005
R832 VTAIL.n407 VTAIL.n406 9.3005
R833 VTAIL.n345 VTAIL.n343 9.3005
R834 VTAIL.n413 VTAIL.n412 9.3005
R835 VTAIL.n437 VTAIL.n436 9.3005
R836 VTAIL.n332 VTAIL.n331 9.3005
R837 VTAIL.n431 VTAIL.n430 9.3005
R838 VTAIL.n429 VTAIL.n428 9.3005
R839 VTAIL.n336 VTAIL.n335 9.3005
R840 VTAIL.n423 VTAIL.n422 9.3005
R841 VTAIL.n421 VTAIL.n420 9.3005
R842 VTAIL.n340 VTAIL.n339 9.3005
R843 VTAIL.n415 VTAIL.n414 9.3005
R844 VTAIL.n391 VTAIL.n390 9.3005
R845 VTAIL.n389 VTAIL.n388 9.3005
R846 VTAIL.n358 VTAIL.n357 9.3005
R847 VTAIL.n383 VTAIL.n382 9.3005
R848 VTAIL.n381 VTAIL.n380 9.3005
R849 VTAIL.n362 VTAIL.n361 9.3005
R850 VTAIL.n375 VTAIL.n374 9.3005
R851 VTAIL.n373 VTAIL.n372 9.3005
R852 VTAIL.n366 VTAIL.n365 9.3005
R853 VTAIL.n822 VTAIL.n821 8.92171
R854 VTAIL.n837 VTAIL.n790 8.92171
R855 VTAIL.n868 VTAIL.n774 8.92171
R856 VTAIL.n52 VTAIL.n51 8.92171
R857 VTAIL.n67 VTAIL.n20 8.92171
R858 VTAIL.n98 VTAIL.n4 8.92171
R859 VTAIL.n162 VTAIL.n161 8.92171
R860 VTAIL.n177 VTAIL.n130 8.92171
R861 VTAIL.n208 VTAIL.n114 8.92171
R862 VTAIL.n272 VTAIL.n271 8.92171
R863 VTAIL.n287 VTAIL.n240 8.92171
R864 VTAIL.n318 VTAIL.n224 8.92171
R865 VTAIL.n758 VTAIL.n664 8.92171
R866 VTAIL.n729 VTAIL.n682 8.92171
R867 VTAIL.n714 VTAIL.n713 8.92171
R868 VTAIL.n648 VTAIL.n554 8.92171
R869 VTAIL.n619 VTAIL.n572 8.92171
R870 VTAIL.n604 VTAIL.n603 8.92171
R871 VTAIL.n538 VTAIL.n444 8.92171
R872 VTAIL.n509 VTAIL.n462 8.92171
R873 VTAIL.n494 VTAIL.n493 8.92171
R874 VTAIL.n428 VTAIL.n334 8.92171
R875 VTAIL.n399 VTAIL.n352 8.92171
R876 VTAIL.n384 VTAIL.n383 8.92171
R877 VTAIL.n825 VTAIL.n796 8.14595
R878 VTAIL.n834 VTAIL.n833 8.14595
R879 VTAIL.n872 VTAIL.n871 8.14595
R880 VTAIL.n55 VTAIL.n26 8.14595
R881 VTAIL.n64 VTAIL.n63 8.14595
R882 VTAIL.n102 VTAIL.n101 8.14595
R883 VTAIL.n165 VTAIL.n136 8.14595
R884 VTAIL.n174 VTAIL.n173 8.14595
R885 VTAIL.n212 VTAIL.n211 8.14595
R886 VTAIL.n275 VTAIL.n246 8.14595
R887 VTAIL.n284 VTAIL.n283 8.14595
R888 VTAIL.n322 VTAIL.n321 8.14595
R889 VTAIL.n762 VTAIL.n761 8.14595
R890 VTAIL.n726 VTAIL.n725 8.14595
R891 VTAIL.n717 VTAIL.n688 8.14595
R892 VTAIL.n652 VTAIL.n651 8.14595
R893 VTAIL.n616 VTAIL.n615 8.14595
R894 VTAIL.n607 VTAIL.n578 8.14595
R895 VTAIL.n542 VTAIL.n541 8.14595
R896 VTAIL.n506 VTAIL.n505 8.14595
R897 VTAIL.n497 VTAIL.n468 8.14595
R898 VTAIL.n432 VTAIL.n431 8.14595
R899 VTAIL.n396 VTAIL.n395 8.14595
R900 VTAIL.n387 VTAIL.n358 8.14595
R901 VTAIL.n826 VTAIL.n794 7.3702
R902 VTAIL.n830 VTAIL.n792 7.3702
R903 VTAIL.n875 VTAIL.n772 7.3702
R904 VTAIL.n878 VTAIL.n770 7.3702
R905 VTAIL.n56 VTAIL.n24 7.3702
R906 VTAIL.n60 VTAIL.n22 7.3702
R907 VTAIL.n105 VTAIL.n2 7.3702
R908 VTAIL.n108 VTAIL.n0 7.3702
R909 VTAIL.n166 VTAIL.n134 7.3702
R910 VTAIL.n170 VTAIL.n132 7.3702
R911 VTAIL.n215 VTAIL.n112 7.3702
R912 VTAIL.n218 VTAIL.n110 7.3702
R913 VTAIL.n276 VTAIL.n244 7.3702
R914 VTAIL.n280 VTAIL.n242 7.3702
R915 VTAIL.n325 VTAIL.n222 7.3702
R916 VTAIL.n328 VTAIL.n220 7.3702
R917 VTAIL.n768 VTAIL.n660 7.3702
R918 VTAIL.n765 VTAIL.n662 7.3702
R919 VTAIL.n722 VTAIL.n684 7.3702
R920 VTAIL.n718 VTAIL.n686 7.3702
R921 VTAIL.n658 VTAIL.n550 7.3702
R922 VTAIL.n655 VTAIL.n552 7.3702
R923 VTAIL.n612 VTAIL.n574 7.3702
R924 VTAIL.n608 VTAIL.n576 7.3702
R925 VTAIL.n548 VTAIL.n440 7.3702
R926 VTAIL.n545 VTAIL.n442 7.3702
R927 VTAIL.n502 VTAIL.n464 7.3702
R928 VTAIL.n498 VTAIL.n466 7.3702
R929 VTAIL.n438 VTAIL.n330 7.3702
R930 VTAIL.n435 VTAIL.n332 7.3702
R931 VTAIL.n392 VTAIL.n354 7.3702
R932 VTAIL.n388 VTAIL.n356 7.3702
R933 VTAIL.n829 VTAIL.n794 6.59444
R934 VTAIL.n830 VTAIL.n829 6.59444
R935 VTAIL.n876 VTAIL.n875 6.59444
R936 VTAIL.n876 VTAIL.n770 6.59444
R937 VTAIL.n59 VTAIL.n24 6.59444
R938 VTAIL.n60 VTAIL.n59 6.59444
R939 VTAIL.n106 VTAIL.n105 6.59444
R940 VTAIL.n106 VTAIL.n0 6.59444
R941 VTAIL.n169 VTAIL.n134 6.59444
R942 VTAIL.n170 VTAIL.n169 6.59444
R943 VTAIL.n216 VTAIL.n215 6.59444
R944 VTAIL.n216 VTAIL.n110 6.59444
R945 VTAIL.n279 VTAIL.n244 6.59444
R946 VTAIL.n280 VTAIL.n279 6.59444
R947 VTAIL.n326 VTAIL.n325 6.59444
R948 VTAIL.n326 VTAIL.n220 6.59444
R949 VTAIL.n766 VTAIL.n660 6.59444
R950 VTAIL.n766 VTAIL.n765 6.59444
R951 VTAIL.n722 VTAIL.n721 6.59444
R952 VTAIL.n721 VTAIL.n686 6.59444
R953 VTAIL.n656 VTAIL.n550 6.59444
R954 VTAIL.n656 VTAIL.n655 6.59444
R955 VTAIL.n612 VTAIL.n611 6.59444
R956 VTAIL.n611 VTAIL.n576 6.59444
R957 VTAIL.n546 VTAIL.n440 6.59444
R958 VTAIL.n546 VTAIL.n545 6.59444
R959 VTAIL.n502 VTAIL.n501 6.59444
R960 VTAIL.n501 VTAIL.n466 6.59444
R961 VTAIL.n436 VTAIL.n330 6.59444
R962 VTAIL.n436 VTAIL.n435 6.59444
R963 VTAIL.n392 VTAIL.n391 6.59444
R964 VTAIL.n391 VTAIL.n356 6.59444
R965 VTAIL.n826 VTAIL.n825 5.81868
R966 VTAIL.n833 VTAIL.n792 5.81868
R967 VTAIL.n872 VTAIL.n772 5.81868
R968 VTAIL.n56 VTAIL.n55 5.81868
R969 VTAIL.n63 VTAIL.n22 5.81868
R970 VTAIL.n102 VTAIL.n2 5.81868
R971 VTAIL.n166 VTAIL.n165 5.81868
R972 VTAIL.n173 VTAIL.n132 5.81868
R973 VTAIL.n212 VTAIL.n112 5.81868
R974 VTAIL.n276 VTAIL.n275 5.81868
R975 VTAIL.n283 VTAIL.n242 5.81868
R976 VTAIL.n322 VTAIL.n222 5.81868
R977 VTAIL.n762 VTAIL.n662 5.81868
R978 VTAIL.n725 VTAIL.n684 5.81868
R979 VTAIL.n718 VTAIL.n717 5.81868
R980 VTAIL.n652 VTAIL.n552 5.81868
R981 VTAIL.n615 VTAIL.n574 5.81868
R982 VTAIL.n608 VTAIL.n607 5.81868
R983 VTAIL.n542 VTAIL.n442 5.81868
R984 VTAIL.n505 VTAIL.n464 5.81868
R985 VTAIL.n498 VTAIL.n497 5.81868
R986 VTAIL.n432 VTAIL.n332 5.81868
R987 VTAIL.n395 VTAIL.n354 5.81868
R988 VTAIL.n388 VTAIL.n387 5.81868
R989 VTAIL.n822 VTAIL.n796 5.04292
R990 VTAIL.n834 VTAIL.n790 5.04292
R991 VTAIL.n871 VTAIL.n774 5.04292
R992 VTAIL.n52 VTAIL.n26 5.04292
R993 VTAIL.n64 VTAIL.n20 5.04292
R994 VTAIL.n101 VTAIL.n4 5.04292
R995 VTAIL.n162 VTAIL.n136 5.04292
R996 VTAIL.n174 VTAIL.n130 5.04292
R997 VTAIL.n211 VTAIL.n114 5.04292
R998 VTAIL.n272 VTAIL.n246 5.04292
R999 VTAIL.n284 VTAIL.n240 5.04292
R1000 VTAIL.n321 VTAIL.n224 5.04292
R1001 VTAIL.n761 VTAIL.n664 5.04292
R1002 VTAIL.n726 VTAIL.n682 5.04292
R1003 VTAIL.n714 VTAIL.n688 5.04292
R1004 VTAIL.n651 VTAIL.n554 5.04292
R1005 VTAIL.n616 VTAIL.n572 5.04292
R1006 VTAIL.n604 VTAIL.n578 5.04292
R1007 VTAIL.n541 VTAIL.n444 5.04292
R1008 VTAIL.n506 VTAIL.n462 5.04292
R1009 VTAIL.n494 VTAIL.n468 5.04292
R1010 VTAIL.n431 VTAIL.n334 5.04292
R1011 VTAIL.n396 VTAIL.n352 5.04292
R1012 VTAIL.n384 VTAIL.n358 5.04292
R1013 VTAIL.n805 VTAIL.n803 4.38563
R1014 VTAIL.n35 VTAIL.n33 4.38563
R1015 VTAIL.n145 VTAIL.n143 4.38563
R1016 VTAIL.n255 VTAIL.n253 4.38563
R1017 VTAIL.n697 VTAIL.n695 4.38563
R1018 VTAIL.n587 VTAIL.n585 4.38563
R1019 VTAIL.n477 VTAIL.n475 4.38563
R1020 VTAIL.n367 VTAIL.n365 4.38563
R1021 VTAIL.n821 VTAIL.n798 4.26717
R1022 VTAIL.n838 VTAIL.n837 4.26717
R1023 VTAIL.n868 VTAIL.n867 4.26717
R1024 VTAIL.n51 VTAIL.n28 4.26717
R1025 VTAIL.n68 VTAIL.n67 4.26717
R1026 VTAIL.n98 VTAIL.n97 4.26717
R1027 VTAIL.n161 VTAIL.n138 4.26717
R1028 VTAIL.n178 VTAIL.n177 4.26717
R1029 VTAIL.n208 VTAIL.n207 4.26717
R1030 VTAIL.n271 VTAIL.n248 4.26717
R1031 VTAIL.n288 VTAIL.n287 4.26717
R1032 VTAIL.n318 VTAIL.n317 4.26717
R1033 VTAIL.n758 VTAIL.n757 4.26717
R1034 VTAIL.n730 VTAIL.n729 4.26717
R1035 VTAIL.n713 VTAIL.n690 4.26717
R1036 VTAIL.n648 VTAIL.n647 4.26717
R1037 VTAIL.n620 VTAIL.n619 4.26717
R1038 VTAIL.n603 VTAIL.n580 4.26717
R1039 VTAIL.n538 VTAIL.n537 4.26717
R1040 VTAIL.n510 VTAIL.n509 4.26717
R1041 VTAIL.n493 VTAIL.n470 4.26717
R1042 VTAIL.n428 VTAIL.n427 4.26717
R1043 VTAIL.n400 VTAIL.n399 4.26717
R1044 VTAIL.n383 VTAIL.n360 4.26717
R1045 VTAIL.n549 VTAIL.n439 3.5436
R1046 VTAIL.n769 VTAIL.n659 3.5436
R1047 VTAIL.n329 VTAIL.n219 3.5436
R1048 VTAIL.n818 VTAIL.n817 3.49141
R1049 VTAIL.n841 VTAIL.n788 3.49141
R1050 VTAIL.n864 VTAIL.n776 3.49141
R1051 VTAIL.n48 VTAIL.n47 3.49141
R1052 VTAIL.n71 VTAIL.n18 3.49141
R1053 VTAIL.n94 VTAIL.n6 3.49141
R1054 VTAIL.n158 VTAIL.n157 3.49141
R1055 VTAIL.n181 VTAIL.n128 3.49141
R1056 VTAIL.n204 VTAIL.n116 3.49141
R1057 VTAIL.n268 VTAIL.n267 3.49141
R1058 VTAIL.n291 VTAIL.n238 3.49141
R1059 VTAIL.n314 VTAIL.n226 3.49141
R1060 VTAIL.n754 VTAIL.n666 3.49141
R1061 VTAIL.n733 VTAIL.n680 3.49141
R1062 VTAIL.n710 VTAIL.n709 3.49141
R1063 VTAIL.n644 VTAIL.n556 3.49141
R1064 VTAIL.n623 VTAIL.n570 3.49141
R1065 VTAIL.n600 VTAIL.n599 3.49141
R1066 VTAIL.n534 VTAIL.n446 3.49141
R1067 VTAIL.n513 VTAIL.n460 3.49141
R1068 VTAIL.n490 VTAIL.n489 3.49141
R1069 VTAIL.n424 VTAIL.n336 3.49141
R1070 VTAIL.n403 VTAIL.n350 3.49141
R1071 VTAIL.n380 VTAIL.n379 3.49141
R1072 VTAIL.n814 VTAIL.n800 2.71565
R1073 VTAIL.n842 VTAIL.n786 2.71565
R1074 VTAIL.n863 VTAIL.n778 2.71565
R1075 VTAIL.n44 VTAIL.n30 2.71565
R1076 VTAIL.n72 VTAIL.n16 2.71565
R1077 VTAIL.n93 VTAIL.n8 2.71565
R1078 VTAIL.n154 VTAIL.n140 2.71565
R1079 VTAIL.n182 VTAIL.n126 2.71565
R1080 VTAIL.n203 VTAIL.n118 2.71565
R1081 VTAIL.n264 VTAIL.n250 2.71565
R1082 VTAIL.n292 VTAIL.n236 2.71565
R1083 VTAIL.n313 VTAIL.n228 2.71565
R1084 VTAIL.n753 VTAIL.n668 2.71565
R1085 VTAIL.n734 VTAIL.n678 2.71565
R1086 VTAIL.n706 VTAIL.n692 2.71565
R1087 VTAIL.n643 VTAIL.n558 2.71565
R1088 VTAIL.n624 VTAIL.n568 2.71565
R1089 VTAIL.n596 VTAIL.n582 2.71565
R1090 VTAIL.n533 VTAIL.n448 2.71565
R1091 VTAIL.n514 VTAIL.n458 2.71565
R1092 VTAIL.n486 VTAIL.n472 2.71565
R1093 VTAIL.n423 VTAIL.n338 2.71565
R1094 VTAIL.n404 VTAIL.n348 2.71565
R1095 VTAIL.n376 VTAIL.n362 2.71565
R1096 VTAIL.n813 VTAIL.n802 1.93989
R1097 VTAIL.n847 VTAIL.n845 1.93989
R1098 VTAIL.n860 VTAIL.n859 1.93989
R1099 VTAIL.n43 VTAIL.n32 1.93989
R1100 VTAIL.n77 VTAIL.n75 1.93989
R1101 VTAIL.n90 VTAIL.n89 1.93989
R1102 VTAIL.n153 VTAIL.n142 1.93989
R1103 VTAIL.n187 VTAIL.n185 1.93989
R1104 VTAIL.n200 VTAIL.n199 1.93989
R1105 VTAIL.n263 VTAIL.n252 1.93989
R1106 VTAIL.n297 VTAIL.n295 1.93989
R1107 VTAIL.n310 VTAIL.n309 1.93989
R1108 VTAIL.n750 VTAIL.n749 1.93989
R1109 VTAIL.n738 VTAIL.n737 1.93989
R1110 VTAIL.n705 VTAIL.n694 1.93989
R1111 VTAIL.n640 VTAIL.n639 1.93989
R1112 VTAIL.n628 VTAIL.n627 1.93989
R1113 VTAIL.n595 VTAIL.n584 1.93989
R1114 VTAIL.n530 VTAIL.n529 1.93989
R1115 VTAIL.n518 VTAIL.n517 1.93989
R1116 VTAIL.n485 VTAIL.n474 1.93989
R1117 VTAIL.n420 VTAIL.n419 1.93989
R1118 VTAIL.n408 VTAIL.n407 1.93989
R1119 VTAIL.n375 VTAIL.n364 1.93989
R1120 VTAIL VTAIL.n109 1.83024
R1121 VTAIL VTAIL.n879 1.71386
R1122 VTAIL.n810 VTAIL.n809 1.16414
R1123 VTAIL.n846 VTAIL.n784 1.16414
R1124 VTAIL.n856 VTAIL.n780 1.16414
R1125 VTAIL.n40 VTAIL.n39 1.16414
R1126 VTAIL.n76 VTAIL.n14 1.16414
R1127 VTAIL.n86 VTAIL.n10 1.16414
R1128 VTAIL.n150 VTAIL.n149 1.16414
R1129 VTAIL.n186 VTAIL.n124 1.16414
R1130 VTAIL.n196 VTAIL.n120 1.16414
R1131 VTAIL.n260 VTAIL.n259 1.16414
R1132 VTAIL.n296 VTAIL.n234 1.16414
R1133 VTAIL.n306 VTAIL.n230 1.16414
R1134 VTAIL.n746 VTAIL.n670 1.16414
R1135 VTAIL.n741 VTAIL.n675 1.16414
R1136 VTAIL.n702 VTAIL.n701 1.16414
R1137 VTAIL.n636 VTAIL.n560 1.16414
R1138 VTAIL.n631 VTAIL.n565 1.16414
R1139 VTAIL.n592 VTAIL.n591 1.16414
R1140 VTAIL.n526 VTAIL.n450 1.16414
R1141 VTAIL.n521 VTAIL.n455 1.16414
R1142 VTAIL.n482 VTAIL.n481 1.16414
R1143 VTAIL.n416 VTAIL.n340 1.16414
R1144 VTAIL.n411 VTAIL.n345 1.16414
R1145 VTAIL.n372 VTAIL.n371 1.16414
R1146 VTAIL.n659 VTAIL.n549 0.470328
R1147 VTAIL.n219 VTAIL.n109 0.470328
R1148 VTAIL.n806 VTAIL.n804 0.388379
R1149 VTAIL.n852 VTAIL.n851 0.388379
R1150 VTAIL.n855 VTAIL.n782 0.388379
R1151 VTAIL.n36 VTAIL.n34 0.388379
R1152 VTAIL.n82 VTAIL.n81 0.388379
R1153 VTAIL.n85 VTAIL.n12 0.388379
R1154 VTAIL.n146 VTAIL.n144 0.388379
R1155 VTAIL.n192 VTAIL.n191 0.388379
R1156 VTAIL.n195 VTAIL.n122 0.388379
R1157 VTAIL.n256 VTAIL.n254 0.388379
R1158 VTAIL.n302 VTAIL.n301 0.388379
R1159 VTAIL.n305 VTAIL.n232 0.388379
R1160 VTAIL.n745 VTAIL.n672 0.388379
R1161 VTAIL.n742 VTAIL.n674 0.388379
R1162 VTAIL.n698 VTAIL.n696 0.388379
R1163 VTAIL.n635 VTAIL.n562 0.388379
R1164 VTAIL.n632 VTAIL.n564 0.388379
R1165 VTAIL.n588 VTAIL.n586 0.388379
R1166 VTAIL.n525 VTAIL.n452 0.388379
R1167 VTAIL.n522 VTAIL.n454 0.388379
R1168 VTAIL.n478 VTAIL.n476 0.388379
R1169 VTAIL.n415 VTAIL.n342 0.388379
R1170 VTAIL.n412 VTAIL.n344 0.388379
R1171 VTAIL.n368 VTAIL.n366 0.388379
R1172 VTAIL.n811 VTAIL.n803 0.155672
R1173 VTAIL.n812 VTAIL.n811 0.155672
R1174 VTAIL.n812 VTAIL.n799 0.155672
R1175 VTAIL.n819 VTAIL.n799 0.155672
R1176 VTAIL.n820 VTAIL.n819 0.155672
R1177 VTAIL.n820 VTAIL.n795 0.155672
R1178 VTAIL.n827 VTAIL.n795 0.155672
R1179 VTAIL.n828 VTAIL.n827 0.155672
R1180 VTAIL.n828 VTAIL.n791 0.155672
R1181 VTAIL.n835 VTAIL.n791 0.155672
R1182 VTAIL.n836 VTAIL.n835 0.155672
R1183 VTAIL.n836 VTAIL.n787 0.155672
R1184 VTAIL.n843 VTAIL.n787 0.155672
R1185 VTAIL.n844 VTAIL.n843 0.155672
R1186 VTAIL.n844 VTAIL.n783 0.155672
R1187 VTAIL.n853 VTAIL.n783 0.155672
R1188 VTAIL.n854 VTAIL.n853 0.155672
R1189 VTAIL.n854 VTAIL.n779 0.155672
R1190 VTAIL.n861 VTAIL.n779 0.155672
R1191 VTAIL.n862 VTAIL.n861 0.155672
R1192 VTAIL.n862 VTAIL.n775 0.155672
R1193 VTAIL.n869 VTAIL.n775 0.155672
R1194 VTAIL.n870 VTAIL.n869 0.155672
R1195 VTAIL.n870 VTAIL.n771 0.155672
R1196 VTAIL.n877 VTAIL.n771 0.155672
R1197 VTAIL.n41 VTAIL.n33 0.155672
R1198 VTAIL.n42 VTAIL.n41 0.155672
R1199 VTAIL.n42 VTAIL.n29 0.155672
R1200 VTAIL.n49 VTAIL.n29 0.155672
R1201 VTAIL.n50 VTAIL.n49 0.155672
R1202 VTAIL.n50 VTAIL.n25 0.155672
R1203 VTAIL.n57 VTAIL.n25 0.155672
R1204 VTAIL.n58 VTAIL.n57 0.155672
R1205 VTAIL.n58 VTAIL.n21 0.155672
R1206 VTAIL.n65 VTAIL.n21 0.155672
R1207 VTAIL.n66 VTAIL.n65 0.155672
R1208 VTAIL.n66 VTAIL.n17 0.155672
R1209 VTAIL.n73 VTAIL.n17 0.155672
R1210 VTAIL.n74 VTAIL.n73 0.155672
R1211 VTAIL.n74 VTAIL.n13 0.155672
R1212 VTAIL.n83 VTAIL.n13 0.155672
R1213 VTAIL.n84 VTAIL.n83 0.155672
R1214 VTAIL.n84 VTAIL.n9 0.155672
R1215 VTAIL.n91 VTAIL.n9 0.155672
R1216 VTAIL.n92 VTAIL.n91 0.155672
R1217 VTAIL.n92 VTAIL.n5 0.155672
R1218 VTAIL.n99 VTAIL.n5 0.155672
R1219 VTAIL.n100 VTAIL.n99 0.155672
R1220 VTAIL.n100 VTAIL.n1 0.155672
R1221 VTAIL.n107 VTAIL.n1 0.155672
R1222 VTAIL.n151 VTAIL.n143 0.155672
R1223 VTAIL.n152 VTAIL.n151 0.155672
R1224 VTAIL.n152 VTAIL.n139 0.155672
R1225 VTAIL.n159 VTAIL.n139 0.155672
R1226 VTAIL.n160 VTAIL.n159 0.155672
R1227 VTAIL.n160 VTAIL.n135 0.155672
R1228 VTAIL.n167 VTAIL.n135 0.155672
R1229 VTAIL.n168 VTAIL.n167 0.155672
R1230 VTAIL.n168 VTAIL.n131 0.155672
R1231 VTAIL.n175 VTAIL.n131 0.155672
R1232 VTAIL.n176 VTAIL.n175 0.155672
R1233 VTAIL.n176 VTAIL.n127 0.155672
R1234 VTAIL.n183 VTAIL.n127 0.155672
R1235 VTAIL.n184 VTAIL.n183 0.155672
R1236 VTAIL.n184 VTAIL.n123 0.155672
R1237 VTAIL.n193 VTAIL.n123 0.155672
R1238 VTAIL.n194 VTAIL.n193 0.155672
R1239 VTAIL.n194 VTAIL.n119 0.155672
R1240 VTAIL.n201 VTAIL.n119 0.155672
R1241 VTAIL.n202 VTAIL.n201 0.155672
R1242 VTAIL.n202 VTAIL.n115 0.155672
R1243 VTAIL.n209 VTAIL.n115 0.155672
R1244 VTAIL.n210 VTAIL.n209 0.155672
R1245 VTAIL.n210 VTAIL.n111 0.155672
R1246 VTAIL.n217 VTAIL.n111 0.155672
R1247 VTAIL.n261 VTAIL.n253 0.155672
R1248 VTAIL.n262 VTAIL.n261 0.155672
R1249 VTAIL.n262 VTAIL.n249 0.155672
R1250 VTAIL.n269 VTAIL.n249 0.155672
R1251 VTAIL.n270 VTAIL.n269 0.155672
R1252 VTAIL.n270 VTAIL.n245 0.155672
R1253 VTAIL.n277 VTAIL.n245 0.155672
R1254 VTAIL.n278 VTAIL.n277 0.155672
R1255 VTAIL.n278 VTAIL.n241 0.155672
R1256 VTAIL.n285 VTAIL.n241 0.155672
R1257 VTAIL.n286 VTAIL.n285 0.155672
R1258 VTAIL.n286 VTAIL.n237 0.155672
R1259 VTAIL.n293 VTAIL.n237 0.155672
R1260 VTAIL.n294 VTAIL.n293 0.155672
R1261 VTAIL.n294 VTAIL.n233 0.155672
R1262 VTAIL.n303 VTAIL.n233 0.155672
R1263 VTAIL.n304 VTAIL.n303 0.155672
R1264 VTAIL.n304 VTAIL.n229 0.155672
R1265 VTAIL.n311 VTAIL.n229 0.155672
R1266 VTAIL.n312 VTAIL.n311 0.155672
R1267 VTAIL.n312 VTAIL.n225 0.155672
R1268 VTAIL.n319 VTAIL.n225 0.155672
R1269 VTAIL.n320 VTAIL.n319 0.155672
R1270 VTAIL.n320 VTAIL.n221 0.155672
R1271 VTAIL.n327 VTAIL.n221 0.155672
R1272 VTAIL.n767 VTAIL.n661 0.155672
R1273 VTAIL.n760 VTAIL.n661 0.155672
R1274 VTAIL.n760 VTAIL.n759 0.155672
R1275 VTAIL.n759 VTAIL.n665 0.155672
R1276 VTAIL.n752 VTAIL.n665 0.155672
R1277 VTAIL.n752 VTAIL.n751 0.155672
R1278 VTAIL.n751 VTAIL.n669 0.155672
R1279 VTAIL.n744 VTAIL.n669 0.155672
R1280 VTAIL.n744 VTAIL.n743 0.155672
R1281 VTAIL.n743 VTAIL.n673 0.155672
R1282 VTAIL.n736 VTAIL.n673 0.155672
R1283 VTAIL.n736 VTAIL.n735 0.155672
R1284 VTAIL.n735 VTAIL.n679 0.155672
R1285 VTAIL.n728 VTAIL.n679 0.155672
R1286 VTAIL.n728 VTAIL.n727 0.155672
R1287 VTAIL.n727 VTAIL.n683 0.155672
R1288 VTAIL.n720 VTAIL.n683 0.155672
R1289 VTAIL.n720 VTAIL.n719 0.155672
R1290 VTAIL.n719 VTAIL.n687 0.155672
R1291 VTAIL.n712 VTAIL.n687 0.155672
R1292 VTAIL.n712 VTAIL.n711 0.155672
R1293 VTAIL.n711 VTAIL.n691 0.155672
R1294 VTAIL.n704 VTAIL.n691 0.155672
R1295 VTAIL.n704 VTAIL.n703 0.155672
R1296 VTAIL.n703 VTAIL.n695 0.155672
R1297 VTAIL.n657 VTAIL.n551 0.155672
R1298 VTAIL.n650 VTAIL.n551 0.155672
R1299 VTAIL.n650 VTAIL.n649 0.155672
R1300 VTAIL.n649 VTAIL.n555 0.155672
R1301 VTAIL.n642 VTAIL.n555 0.155672
R1302 VTAIL.n642 VTAIL.n641 0.155672
R1303 VTAIL.n641 VTAIL.n559 0.155672
R1304 VTAIL.n634 VTAIL.n559 0.155672
R1305 VTAIL.n634 VTAIL.n633 0.155672
R1306 VTAIL.n633 VTAIL.n563 0.155672
R1307 VTAIL.n626 VTAIL.n563 0.155672
R1308 VTAIL.n626 VTAIL.n625 0.155672
R1309 VTAIL.n625 VTAIL.n569 0.155672
R1310 VTAIL.n618 VTAIL.n569 0.155672
R1311 VTAIL.n618 VTAIL.n617 0.155672
R1312 VTAIL.n617 VTAIL.n573 0.155672
R1313 VTAIL.n610 VTAIL.n573 0.155672
R1314 VTAIL.n610 VTAIL.n609 0.155672
R1315 VTAIL.n609 VTAIL.n577 0.155672
R1316 VTAIL.n602 VTAIL.n577 0.155672
R1317 VTAIL.n602 VTAIL.n601 0.155672
R1318 VTAIL.n601 VTAIL.n581 0.155672
R1319 VTAIL.n594 VTAIL.n581 0.155672
R1320 VTAIL.n594 VTAIL.n593 0.155672
R1321 VTAIL.n593 VTAIL.n585 0.155672
R1322 VTAIL.n547 VTAIL.n441 0.155672
R1323 VTAIL.n540 VTAIL.n441 0.155672
R1324 VTAIL.n540 VTAIL.n539 0.155672
R1325 VTAIL.n539 VTAIL.n445 0.155672
R1326 VTAIL.n532 VTAIL.n445 0.155672
R1327 VTAIL.n532 VTAIL.n531 0.155672
R1328 VTAIL.n531 VTAIL.n449 0.155672
R1329 VTAIL.n524 VTAIL.n449 0.155672
R1330 VTAIL.n524 VTAIL.n523 0.155672
R1331 VTAIL.n523 VTAIL.n453 0.155672
R1332 VTAIL.n516 VTAIL.n453 0.155672
R1333 VTAIL.n516 VTAIL.n515 0.155672
R1334 VTAIL.n515 VTAIL.n459 0.155672
R1335 VTAIL.n508 VTAIL.n459 0.155672
R1336 VTAIL.n508 VTAIL.n507 0.155672
R1337 VTAIL.n507 VTAIL.n463 0.155672
R1338 VTAIL.n500 VTAIL.n463 0.155672
R1339 VTAIL.n500 VTAIL.n499 0.155672
R1340 VTAIL.n499 VTAIL.n467 0.155672
R1341 VTAIL.n492 VTAIL.n467 0.155672
R1342 VTAIL.n492 VTAIL.n491 0.155672
R1343 VTAIL.n491 VTAIL.n471 0.155672
R1344 VTAIL.n484 VTAIL.n471 0.155672
R1345 VTAIL.n484 VTAIL.n483 0.155672
R1346 VTAIL.n483 VTAIL.n475 0.155672
R1347 VTAIL.n437 VTAIL.n331 0.155672
R1348 VTAIL.n430 VTAIL.n331 0.155672
R1349 VTAIL.n430 VTAIL.n429 0.155672
R1350 VTAIL.n429 VTAIL.n335 0.155672
R1351 VTAIL.n422 VTAIL.n335 0.155672
R1352 VTAIL.n422 VTAIL.n421 0.155672
R1353 VTAIL.n421 VTAIL.n339 0.155672
R1354 VTAIL.n414 VTAIL.n339 0.155672
R1355 VTAIL.n414 VTAIL.n413 0.155672
R1356 VTAIL.n413 VTAIL.n343 0.155672
R1357 VTAIL.n406 VTAIL.n343 0.155672
R1358 VTAIL.n406 VTAIL.n405 0.155672
R1359 VTAIL.n405 VTAIL.n349 0.155672
R1360 VTAIL.n398 VTAIL.n349 0.155672
R1361 VTAIL.n398 VTAIL.n397 0.155672
R1362 VTAIL.n397 VTAIL.n353 0.155672
R1363 VTAIL.n390 VTAIL.n353 0.155672
R1364 VTAIL.n390 VTAIL.n389 0.155672
R1365 VTAIL.n389 VTAIL.n357 0.155672
R1366 VTAIL.n382 VTAIL.n357 0.155672
R1367 VTAIL.n382 VTAIL.n381 0.155672
R1368 VTAIL.n381 VTAIL.n361 0.155672
R1369 VTAIL.n374 VTAIL.n361 0.155672
R1370 VTAIL.n374 VTAIL.n373 0.155672
R1371 VTAIL.n373 VTAIL.n365 0.155672
R1372 B.n1057 B.n1056 585
R1373 B.n429 B.n152 585
R1374 B.n428 B.n427 585
R1375 B.n426 B.n425 585
R1376 B.n424 B.n423 585
R1377 B.n422 B.n421 585
R1378 B.n420 B.n419 585
R1379 B.n418 B.n417 585
R1380 B.n416 B.n415 585
R1381 B.n414 B.n413 585
R1382 B.n412 B.n411 585
R1383 B.n410 B.n409 585
R1384 B.n408 B.n407 585
R1385 B.n406 B.n405 585
R1386 B.n404 B.n403 585
R1387 B.n402 B.n401 585
R1388 B.n400 B.n399 585
R1389 B.n398 B.n397 585
R1390 B.n396 B.n395 585
R1391 B.n394 B.n393 585
R1392 B.n392 B.n391 585
R1393 B.n390 B.n389 585
R1394 B.n388 B.n387 585
R1395 B.n386 B.n385 585
R1396 B.n384 B.n383 585
R1397 B.n382 B.n381 585
R1398 B.n380 B.n379 585
R1399 B.n378 B.n377 585
R1400 B.n376 B.n375 585
R1401 B.n374 B.n373 585
R1402 B.n372 B.n371 585
R1403 B.n370 B.n369 585
R1404 B.n368 B.n367 585
R1405 B.n366 B.n365 585
R1406 B.n364 B.n363 585
R1407 B.n362 B.n361 585
R1408 B.n360 B.n359 585
R1409 B.n358 B.n357 585
R1410 B.n356 B.n355 585
R1411 B.n354 B.n353 585
R1412 B.n352 B.n351 585
R1413 B.n350 B.n349 585
R1414 B.n348 B.n347 585
R1415 B.n346 B.n345 585
R1416 B.n344 B.n343 585
R1417 B.n342 B.n341 585
R1418 B.n340 B.n339 585
R1419 B.n338 B.n337 585
R1420 B.n336 B.n335 585
R1421 B.n334 B.n333 585
R1422 B.n332 B.n331 585
R1423 B.n330 B.n329 585
R1424 B.n328 B.n327 585
R1425 B.n326 B.n325 585
R1426 B.n324 B.n323 585
R1427 B.n322 B.n321 585
R1428 B.n320 B.n319 585
R1429 B.n318 B.n317 585
R1430 B.n316 B.n315 585
R1431 B.n314 B.n313 585
R1432 B.n312 B.n311 585
R1433 B.n310 B.n309 585
R1434 B.n308 B.n307 585
R1435 B.n306 B.n305 585
R1436 B.n304 B.n303 585
R1437 B.n302 B.n301 585
R1438 B.n300 B.n299 585
R1439 B.n298 B.n297 585
R1440 B.n296 B.n295 585
R1441 B.n294 B.n293 585
R1442 B.n292 B.n291 585
R1443 B.n290 B.n289 585
R1444 B.n288 B.n287 585
R1445 B.n286 B.n285 585
R1446 B.n284 B.n283 585
R1447 B.n282 B.n281 585
R1448 B.n280 B.n279 585
R1449 B.n278 B.n277 585
R1450 B.n276 B.n275 585
R1451 B.n274 B.n273 585
R1452 B.n272 B.n271 585
R1453 B.n270 B.n269 585
R1454 B.n268 B.n267 585
R1455 B.n266 B.n265 585
R1456 B.n264 B.n263 585
R1457 B.n262 B.n261 585
R1458 B.n260 B.n259 585
R1459 B.n258 B.n257 585
R1460 B.n256 B.n255 585
R1461 B.n254 B.n253 585
R1462 B.n252 B.n251 585
R1463 B.n250 B.n249 585
R1464 B.n248 B.n247 585
R1465 B.n246 B.n245 585
R1466 B.n244 B.n243 585
R1467 B.n242 B.n241 585
R1468 B.n240 B.n239 585
R1469 B.n238 B.n237 585
R1470 B.n236 B.n235 585
R1471 B.n234 B.n233 585
R1472 B.n232 B.n231 585
R1473 B.n230 B.n229 585
R1474 B.n228 B.n227 585
R1475 B.n226 B.n225 585
R1476 B.n224 B.n223 585
R1477 B.n222 B.n221 585
R1478 B.n220 B.n219 585
R1479 B.n218 B.n217 585
R1480 B.n216 B.n215 585
R1481 B.n214 B.n213 585
R1482 B.n212 B.n211 585
R1483 B.n210 B.n209 585
R1484 B.n208 B.n207 585
R1485 B.n206 B.n205 585
R1486 B.n204 B.n203 585
R1487 B.n202 B.n201 585
R1488 B.n200 B.n199 585
R1489 B.n198 B.n197 585
R1490 B.n196 B.n195 585
R1491 B.n194 B.n193 585
R1492 B.n192 B.n191 585
R1493 B.n190 B.n189 585
R1494 B.n188 B.n187 585
R1495 B.n186 B.n185 585
R1496 B.n184 B.n183 585
R1497 B.n182 B.n181 585
R1498 B.n180 B.n179 585
R1499 B.n178 B.n177 585
R1500 B.n176 B.n175 585
R1501 B.n174 B.n173 585
R1502 B.n172 B.n171 585
R1503 B.n170 B.n169 585
R1504 B.n168 B.n167 585
R1505 B.n166 B.n165 585
R1506 B.n164 B.n163 585
R1507 B.n162 B.n161 585
R1508 B.n160 B.n159 585
R1509 B.n82 B.n81 585
R1510 B.n1055 B.n83 585
R1511 B.n1060 B.n83 585
R1512 B.n1054 B.n1053 585
R1513 B.n1053 B.n79 585
R1514 B.n1052 B.n78 585
R1515 B.n1066 B.n78 585
R1516 B.n1051 B.n77 585
R1517 B.n1067 B.n77 585
R1518 B.n1050 B.n76 585
R1519 B.n1068 B.n76 585
R1520 B.n1049 B.n1048 585
R1521 B.n1048 B.n72 585
R1522 B.n1047 B.n71 585
R1523 B.n1074 B.n71 585
R1524 B.n1046 B.n70 585
R1525 B.n1075 B.n70 585
R1526 B.n1045 B.n69 585
R1527 B.n1076 B.n69 585
R1528 B.n1044 B.n1043 585
R1529 B.n1043 B.n68 585
R1530 B.n1042 B.n64 585
R1531 B.n1082 B.n64 585
R1532 B.n1041 B.n63 585
R1533 B.n1083 B.n63 585
R1534 B.n1040 B.n62 585
R1535 B.n1084 B.n62 585
R1536 B.n1039 B.n1038 585
R1537 B.n1038 B.n58 585
R1538 B.n1037 B.n57 585
R1539 B.n1090 B.n57 585
R1540 B.n1036 B.n56 585
R1541 B.n1091 B.n56 585
R1542 B.n1035 B.n55 585
R1543 B.n1092 B.n55 585
R1544 B.n1034 B.n1033 585
R1545 B.n1033 B.n51 585
R1546 B.n1032 B.n50 585
R1547 B.n1098 B.n50 585
R1548 B.n1031 B.n49 585
R1549 B.n1099 B.n49 585
R1550 B.n1030 B.n48 585
R1551 B.n1100 B.n48 585
R1552 B.n1029 B.n1028 585
R1553 B.n1028 B.n44 585
R1554 B.n1027 B.n43 585
R1555 B.n1106 B.n43 585
R1556 B.n1026 B.n42 585
R1557 B.n1107 B.n42 585
R1558 B.n1025 B.n41 585
R1559 B.n1108 B.n41 585
R1560 B.n1024 B.n1023 585
R1561 B.n1023 B.n37 585
R1562 B.n1022 B.n36 585
R1563 B.n1114 B.n36 585
R1564 B.n1021 B.n35 585
R1565 B.n1115 B.n35 585
R1566 B.n1020 B.n34 585
R1567 B.n1116 B.n34 585
R1568 B.n1019 B.n1018 585
R1569 B.n1018 B.n30 585
R1570 B.n1017 B.n29 585
R1571 B.n1122 B.n29 585
R1572 B.n1016 B.n28 585
R1573 B.n1123 B.n28 585
R1574 B.n1015 B.n27 585
R1575 B.n1124 B.n27 585
R1576 B.n1014 B.n1013 585
R1577 B.n1013 B.n23 585
R1578 B.n1012 B.n22 585
R1579 B.n1130 B.n22 585
R1580 B.n1011 B.n21 585
R1581 B.n1131 B.n21 585
R1582 B.n1010 B.n20 585
R1583 B.n1132 B.n20 585
R1584 B.n1009 B.n1008 585
R1585 B.n1008 B.n16 585
R1586 B.n1007 B.n15 585
R1587 B.n1138 B.n15 585
R1588 B.n1006 B.n14 585
R1589 B.n1139 B.n14 585
R1590 B.n1005 B.n13 585
R1591 B.n1140 B.n13 585
R1592 B.n1004 B.n1003 585
R1593 B.n1003 B.n12 585
R1594 B.n1002 B.n1001 585
R1595 B.n1002 B.n8 585
R1596 B.n1000 B.n7 585
R1597 B.n1147 B.n7 585
R1598 B.n999 B.n6 585
R1599 B.n1148 B.n6 585
R1600 B.n998 B.n5 585
R1601 B.n1149 B.n5 585
R1602 B.n997 B.n996 585
R1603 B.n996 B.n4 585
R1604 B.n995 B.n430 585
R1605 B.n995 B.n994 585
R1606 B.n985 B.n431 585
R1607 B.n432 B.n431 585
R1608 B.n987 B.n986 585
R1609 B.n988 B.n987 585
R1610 B.n984 B.n437 585
R1611 B.n437 B.n436 585
R1612 B.n983 B.n982 585
R1613 B.n982 B.n981 585
R1614 B.n439 B.n438 585
R1615 B.n440 B.n439 585
R1616 B.n974 B.n973 585
R1617 B.n975 B.n974 585
R1618 B.n972 B.n445 585
R1619 B.n445 B.n444 585
R1620 B.n971 B.n970 585
R1621 B.n970 B.n969 585
R1622 B.n447 B.n446 585
R1623 B.n448 B.n447 585
R1624 B.n962 B.n961 585
R1625 B.n963 B.n962 585
R1626 B.n960 B.n453 585
R1627 B.n453 B.n452 585
R1628 B.n959 B.n958 585
R1629 B.n958 B.n957 585
R1630 B.n455 B.n454 585
R1631 B.n456 B.n455 585
R1632 B.n950 B.n949 585
R1633 B.n951 B.n950 585
R1634 B.n948 B.n461 585
R1635 B.n461 B.n460 585
R1636 B.n947 B.n946 585
R1637 B.n946 B.n945 585
R1638 B.n463 B.n462 585
R1639 B.n464 B.n463 585
R1640 B.n938 B.n937 585
R1641 B.n939 B.n938 585
R1642 B.n936 B.n469 585
R1643 B.n469 B.n468 585
R1644 B.n935 B.n934 585
R1645 B.n934 B.n933 585
R1646 B.n471 B.n470 585
R1647 B.n472 B.n471 585
R1648 B.n926 B.n925 585
R1649 B.n927 B.n926 585
R1650 B.n924 B.n477 585
R1651 B.n477 B.n476 585
R1652 B.n923 B.n922 585
R1653 B.n922 B.n921 585
R1654 B.n479 B.n478 585
R1655 B.n480 B.n479 585
R1656 B.n914 B.n913 585
R1657 B.n915 B.n914 585
R1658 B.n912 B.n485 585
R1659 B.n485 B.n484 585
R1660 B.n911 B.n910 585
R1661 B.n910 B.n909 585
R1662 B.n487 B.n486 585
R1663 B.n488 B.n487 585
R1664 B.n902 B.n901 585
R1665 B.n903 B.n902 585
R1666 B.n900 B.n493 585
R1667 B.n493 B.n492 585
R1668 B.n899 B.n898 585
R1669 B.n898 B.n897 585
R1670 B.n495 B.n494 585
R1671 B.n890 B.n495 585
R1672 B.n889 B.n888 585
R1673 B.n891 B.n889 585
R1674 B.n887 B.n500 585
R1675 B.n500 B.n499 585
R1676 B.n886 B.n885 585
R1677 B.n885 B.n884 585
R1678 B.n502 B.n501 585
R1679 B.n503 B.n502 585
R1680 B.n877 B.n876 585
R1681 B.n878 B.n877 585
R1682 B.n875 B.n508 585
R1683 B.n508 B.n507 585
R1684 B.n874 B.n873 585
R1685 B.n873 B.n872 585
R1686 B.n510 B.n509 585
R1687 B.n511 B.n510 585
R1688 B.n865 B.n864 585
R1689 B.n866 B.n865 585
R1690 B.n514 B.n513 585
R1691 B.n589 B.n587 585
R1692 B.n590 B.n586 585
R1693 B.n590 B.n515 585
R1694 B.n593 B.n592 585
R1695 B.n594 B.n585 585
R1696 B.n596 B.n595 585
R1697 B.n598 B.n584 585
R1698 B.n601 B.n600 585
R1699 B.n602 B.n583 585
R1700 B.n604 B.n603 585
R1701 B.n606 B.n582 585
R1702 B.n609 B.n608 585
R1703 B.n610 B.n581 585
R1704 B.n612 B.n611 585
R1705 B.n614 B.n580 585
R1706 B.n617 B.n616 585
R1707 B.n618 B.n579 585
R1708 B.n620 B.n619 585
R1709 B.n622 B.n578 585
R1710 B.n625 B.n624 585
R1711 B.n626 B.n577 585
R1712 B.n628 B.n627 585
R1713 B.n630 B.n576 585
R1714 B.n633 B.n632 585
R1715 B.n634 B.n575 585
R1716 B.n636 B.n635 585
R1717 B.n638 B.n574 585
R1718 B.n641 B.n640 585
R1719 B.n642 B.n573 585
R1720 B.n644 B.n643 585
R1721 B.n646 B.n572 585
R1722 B.n649 B.n648 585
R1723 B.n650 B.n571 585
R1724 B.n652 B.n651 585
R1725 B.n654 B.n570 585
R1726 B.n657 B.n656 585
R1727 B.n658 B.n569 585
R1728 B.n660 B.n659 585
R1729 B.n662 B.n568 585
R1730 B.n665 B.n664 585
R1731 B.n666 B.n567 585
R1732 B.n668 B.n667 585
R1733 B.n670 B.n566 585
R1734 B.n673 B.n672 585
R1735 B.n674 B.n565 585
R1736 B.n676 B.n675 585
R1737 B.n678 B.n564 585
R1738 B.n681 B.n680 585
R1739 B.n682 B.n563 585
R1740 B.n684 B.n683 585
R1741 B.n686 B.n562 585
R1742 B.n689 B.n688 585
R1743 B.n690 B.n561 585
R1744 B.n692 B.n691 585
R1745 B.n694 B.n560 585
R1746 B.n697 B.n696 585
R1747 B.n698 B.n559 585
R1748 B.n700 B.n699 585
R1749 B.n702 B.n558 585
R1750 B.n705 B.n704 585
R1751 B.n706 B.n557 585
R1752 B.n708 B.n707 585
R1753 B.n710 B.n556 585
R1754 B.n713 B.n712 585
R1755 B.n715 B.n553 585
R1756 B.n717 B.n716 585
R1757 B.n719 B.n552 585
R1758 B.n722 B.n721 585
R1759 B.n723 B.n551 585
R1760 B.n725 B.n724 585
R1761 B.n727 B.n550 585
R1762 B.n730 B.n729 585
R1763 B.n731 B.n549 585
R1764 B.n736 B.n735 585
R1765 B.n738 B.n548 585
R1766 B.n741 B.n740 585
R1767 B.n742 B.n547 585
R1768 B.n744 B.n743 585
R1769 B.n746 B.n546 585
R1770 B.n749 B.n748 585
R1771 B.n750 B.n545 585
R1772 B.n752 B.n751 585
R1773 B.n754 B.n544 585
R1774 B.n757 B.n756 585
R1775 B.n758 B.n543 585
R1776 B.n760 B.n759 585
R1777 B.n762 B.n542 585
R1778 B.n765 B.n764 585
R1779 B.n766 B.n541 585
R1780 B.n768 B.n767 585
R1781 B.n770 B.n540 585
R1782 B.n773 B.n772 585
R1783 B.n774 B.n539 585
R1784 B.n776 B.n775 585
R1785 B.n778 B.n538 585
R1786 B.n781 B.n780 585
R1787 B.n782 B.n537 585
R1788 B.n784 B.n783 585
R1789 B.n786 B.n536 585
R1790 B.n789 B.n788 585
R1791 B.n790 B.n535 585
R1792 B.n792 B.n791 585
R1793 B.n794 B.n534 585
R1794 B.n797 B.n796 585
R1795 B.n798 B.n533 585
R1796 B.n800 B.n799 585
R1797 B.n802 B.n532 585
R1798 B.n805 B.n804 585
R1799 B.n806 B.n531 585
R1800 B.n808 B.n807 585
R1801 B.n810 B.n530 585
R1802 B.n813 B.n812 585
R1803 B.n814 B.n529 585
R1804 B.n816 B.n815 585
R1805 B.n818 B.n528 585
R1806 B.n821 B.n820 585
R1807 B.n822 B.n527 585
R1808 B.n824 B.n823 585
R1809 B.n826 B.n526 585
R1810 B.n829 B.n828 585
R1811 B.n830 B.n525 585
R1812 B.n832 B.n831 585
R1813 B.n834 B.n524 585
R1814 B.n837 B.n836 585
R1815 B.n838 B.n523 585
R1816 B.n840 B.n839 585
R1817 B.n842 B.n522 585
R1818 B.n845 B.n844 585
R1819 B.n846 B.n521 585
R1820 B.n848 B.n847 585
R1821 B.n850 B.n520 585
R1822 B.n853 B.n852 585
R1823 B.n854 B.n519 585
R1824 B.n856 B.n855 585
R1825 B.n858 B.n518 585
R1826 B.n859 B.n517 585
R1827 B.n862 B.n861 585
R1828 B.n863 B.n516 585
R1829 B.n516 B.n515 585
R1830 B.n868 B.n867 585
R1831 B.n867 B.n866 585
R1832 B.n869 B.n512 585
R1833 B.n512 B.n511 585
R1834 B.n871 B.n870 585
R1835 B.n872 B.n871 585
R1836 B.n506 B.n505 585
R1837 B.n507 B.n506 585
R1838 B.n880 B.n879 585
R1839 B.n879 B.n878 585
R1840 B.n881 B.n504 585
R1841 B.n504 B.n503 585
R1842 B.n883 B.n882 585
R1843 B.n884 B.n883 585
R1844 B.n498 B.n497 585
R1845 B.n499 B.n498 585
R1846 B.n893 B.n892 585
R1847 B.n892 B.n891 585
R1848 B.n894 B.n496 585
R1849 B.n890 B.n496 585
R1850 B.n896 B.n895 585
R1851 B.n897 B.n896 585
R1852 B.n491 B.n490 585
R1853 B.n492 B.n491 585
R1854 B.n905 B.n904 585
R1855 B.n904 B.n903 585
R1856 B.n906 B.n489 585
R1857 B.n489 B.n488 585
R1858 B.n908 B.n907 585
R1859 B.n909 B.n908 585
R1860 B.n483 B.n482 585
R1861 B.n484 B.n483 585
R1862 B.n917 B.n916 585
R1863 B.n916 B.n915 585
R1864 B.n918 B.n481 585
R1865 B.n481 B.n480 585
R1866 B.n920 B.n919 585
R1867 B.n921 B.n920 585
R1868 B.n475 B.n474 585
R1869 B.n476 B.n475 585
R1870 B.n929 B.n928 585
R1871 B.n928 B.n927 585
R1872 B.n930 B.n473 585
R1873 B.n473 B.n472 585
R1874 B.n932 B.n931 585
R1875 B.n933 B.n932 585
R1876 B.n467 B.n466 585
R1877 B.n468 B.n467 585
R1878 B.n941 B.n940 585
R1879 B.n940 B.n939 585
R1880 B.n942 B.n465 585
R1881 B.n465 B.n464 585
R1882 B.n944 B.n943 585
R1883 B.n945 B.n944 585
R1884 B.n459 B.n458 585
R1885 B.n460 B.n459 585
R1886 B.n953 B.n952 585
R1887 B.n952 B.n951 585
R1888 B.n954 B.n457 585
R1889 B.n457 B.n456 585
R1890 B.n956 B.n955 585
R1891 B.n957 B.n956 585
R1892 B.n451 B.n450 585
R1893 B.n452 B.n451 585
R1894 B.n965 B.n964 585
R1895 B.n964 B.n963 585
R1896 B.n966 B.n449 585
R1897 B.n449 B.n448 585
R1898 B.n968 B.n967 585
R1899 B.n969 B.n968 585
R1900 B.n443 B.n442 585
R1901 B.n444 B.n443 585
R1902 B.n977 B.n976 585
R1903 B.n976 B.n975 585
R1904 B.n978 B.n441 585
R1905 B.n441 B.n440 585
R1906 B.n980 B.n979 585
R1907 B.n981 B.n980 585
R1908 B.n435 B.n434 585
R1909 B.n436 B.n435 585
R1910 B.n990 B.n989 585
R1911 B.n989 B.n988 585
R1912 B.n991 B.n433 585
R1913 B.n433 B.n432 585
R1914 B.n993 B.n992 585
R1915 B.n994 B.n993 585
R1916 B.n3 B.n0 585
R1917 B.n4 B.n3 585
R1918 B.n1146 B.n1 585
R1919 B.n1147 B.n1146 585
R1920 B.n1145 B.n1144 585
R1921 B.n1145 B.n8 585
R1922 B.n1143 B.n9 585
R1923 B.n12 B.n9 585
R1924 B.n1142 B.n1141 585
R1925 B.n1141 B.n1140 585
R1926 B.n11 B.n10 585
R1927 B.n1139 B.n11 585
R1928 B.n1137 B.n1136 585
R1929 B.n1138 B.n1137 585
R1930 B.n1135 B.n17 585
R1931 B.n17 B.n16 585
R1932 B.n1134 B.n1133 585
R1933 B.n1133 B.n1132 585
R1934 B.n19 B.n18 585
R1935 B.n1131 B.n19 585
R1936 B.n1129 B.n1128 585
R1937 B.n1130 B.n1129 585
R1938 B.n1127 B.n24 585
R1939 B.n24 B.n23 585
R1940 B.n1126 B.n1125 585
R1941 B.n1125 B.n1124 585
R1942 B.n26 B.n25 585
R1943 B.n1123 B.n26 585
R1944 B.n1121 B.n1120 585
R1945 B.n1122 B.n1121 585
R1946 B.n1119 B.n31 585
R1947 B.n31 B.n30 585
R1948 B.n1118 B.n1117 585
R1949 B.n1117 B.n1116 585
R1950 B.n33 B.n32 585
R1951 B.n1115 B.n33 585
R1952 B.n1113 B.n1112 585
R1953 B.n1114 B.n1113 585
R1954 B.n1111 B.n38 585
R1955 B.n38 B.n37 585
R1956 B.n1110 B.n1109 585
R1957 B.n1109 B.n1108 585
R1958 B.n40 B.n39 585
R1959 B.n1107 B.n40 585
R1960 B.n1105 B.n1104 585
R1961 B.n1106 B.n1105 585
R1962 B.n1103 B.n45 585
R1963 B.n45 B.n44 585
R1964 B.n1102 B.n1101 585
R1965 B.n1101 B.n1100 585
R1966 B.n47 B.n46 585
R1967 B.n1099 B.n47 585
R1968 B.n1097 B.n1096 585
R1969 B.n1098 B.n1097 585
R1970 B.n1095 B.n52 585
R1971 B.n52 B.n51 585
R1972 B.n1094 B.n1093 585
R1973 B.n1093 B.n1092 585
R1974 B.n54 B.n53 585
R1975 B.n1091 B.n54 585
R1976 B.n1089 B.n1088 585
R1977 B.n1090 B.n1089 585
R1978 B.n1087 B.n59 585
R1979 B.n59 B.n58 585
R1980 B.n1086 B.n1085 585
R1981 B.n1085 B.n1084 585
R1982 B.n61 B.n60 585
R1983 B.n1083 B.n61 585
R1984 B.n1081 B.n1080 585
R1985 B.n1082 B.n1081 585
R1986 B.n1079 B.n65 585
R1987 B.n68 B.n65 585
R1988 B.n1078 B.n1077 585
R1989 B.n1077 B.n1076 585
R1990 B.n67 B.n66 585
R1991 B.n1075 B.n67 585
R1992 B.n1073 B.n1072 585
R1993 B.n1074 B.n1073 585
R1994 B.n1071 B.n73 585
R1995 B.n73 B.n72 585
R1996 B.n1070 B.n1069 585
R1997 B.n1069 B.n1068 585
R1998 B.n75 B.n74 585
R1999 B.n1067 B.n75 585
R2000 B.n1065 B.n1064 585
R2001 B.n1066 B.n1065 585
R2002 B.n1063 B.n80 585
R2003 B.n80 B.n79 585
R2004 B.n1062 B.n1061 585
R2005 B.n1061 B.n1060 585
R2006 B.n1150 B.n1149 585
R2007 B.n1148 B.n2 585
R2008 B.n153 B.t6 494.238
R2009 B.n732 B.t14 494.238
R2010 B.n156 B.t9 494.238
R2011 B.n554 B.t17 494.238
R2012 B.n1061 B.n82 473.281
R2013 B.n1057 B.n83 473.281
R2014 B.n865 B.n516 473.281
R2015 B.n867 B.n514 473.281
R2016 B.n154 B.t7 414.529
R2017 B.n733 B.t13 414.529
R2018 B.n157 B.t10 414.529
R2019 B.n555 B.t16 414.529
R2020 B.n156 B.t8 334.738
R2021 B.n153 B.t4 334.738
R2022 B.n732 B.t11 334.738
R2023 B.n554 B.t15 334.738
R2024 B.n1059 B.n1058 256.663
R2025 B.n1059 B.n151 256.663
R2026 B.n1059 B.n150 256.663
R2027 B.n1059 B.n149 256.663
R2028 B.n1059 B.n148 256.663
R2029 B.n1059 B.n147 256.663
R2030 B.n1059 B.n146 256.663
R2031 B.n1059 B.n145 256.663
R2032 B.n1059 B.n144 256.663
R2033 B.n1059 B.n143 256.663
R2034 B.n1059 B.n142 256.663
R2035 B.n1059 B.n141 256.663
R2036 B.n1059 B.n140 256.663
R2037 B.n1059 B.n139 256.663
R2038 B.n1059 B.n138 256.663
R2039 B.n1059 B.n137 256.663
R2040 B.n1059 B.n136 256.663
R2041 B.n1059 B.n135 256.663
R2042 B.n1059 B.n134 256.663
R2043 B.n1059 B.n133 256.663
R2044 B.n1059 B.n132 256.663
R2045 B.n1059 B.n131 256.663
R2046 B.n1059 B.n130 256.663
R2047 B.n1059 B.n129 256.663
R2048 B.n1059 B.n128 256.663
R2049 B.n1059 B.n127 256.663
R2050 B.n1059 B.n126 256.663
R2051 B.n1059 B.n125 256.663
R2052 B.n1059 B.n124 256.663
R2053 B.n1059 B.n123 256.663
R2054 B.n1059 B.n122 256.663
R2055 B.n1059 B.n121 256.663
R2056 B.n1059 B.n120 256.663
R2057 B.n1059 B.n119 256.663
R2058 B.n1059 B.n118 256.663
R2059 B.n1059 B.n117 256.663
R2060 B.n1059 B.n116 256.663
R2061 B.n1059 B.n115 256.663
R2062 B.n1059 B.n114 256.663
R2063 B.n1059 B.n113 256.663
R2064 B.n1059 B.n112 256.663
R2065 B.n1059 B.n111 256.663
R2066 B.n1059 B.n110 256.663
R2067 B.n1059 B.n109 256.663
R2068 B.n1059 B.n108 256.663
R2069 B.n1059 B.n107 256.663
R2070 B.n1059 B.n106 256.663
R2071 B.n1059 B.n105 256.663
R2072 B.n1059 B.n104 256.663
R2073 B.n1059 B.n103 256.663
R2074 B.n1059 B.n102 256.663
R2075 B.n1059 B.n101 256.663
R2076 B.n1059 B.n100 256.663
R2077 B.n1059 B.n99 256.663
R2078 B.n1059 B.n98 256.663
R2079 B.n1059 B.n97 256.663
R2080 B.n1059 B.n96 256.663
R2081 B.n1059 B.n95 256.663
R2082 B.n1059 B.n94 256.663
R2083 B.n1059 B.n93 256.663
R2084 B.n1059 B.n92 256.663
R2085 B.n1059 B.n91 256.663
R2086 B.n1059 B.n90 256.663
R2087 B.n1059 B.n89 256.663
R2088 B.n1059 B.n88 256.663
R2089 B.n1059 B.n87 256.663
R2090 B.n1059 B.n86 256.663
R2091 B.n1059 B.n85 256.663
R2092 B.n1059 B.n84 256.663
R2093 B.n588 B.n515 256.663
R2094 B.n591 B.n515 256.663
R2095 B.n597 B.n515 256.663
R2096 B.n599 B.n515 256.663
R2097 B.n605 B.n515 256.663
R2098 B.n607 B.n515 256.663
R2099 B.n613 B.n515 256.663
R2100 B.n615 B.n515 256.663
R2101 B.n621 B.n515 256.663
R2102 B.n623 B.n515 256.663
R2103 B.n629 B.n515 256.663
R2104 B.n631 B.n515 256.663
R2105 B.n637 B.n515 256.663
R2106 B.n639 B.n515 256.663
R2107 B.n645 B.n515 256.663
R2108 B.n647 B.n515 256.663
R2109 B.n653 B.n515 256.663
R2110 B.n655 B.n515 256.663
R2111 B.n661 B.n515 256.663
R2112 B.n663 B.n515 256.663
R2113 B.n669 B.n515 256.663
R2114 B.n671 B.n515 256.663
R2115 B.n677 B.n515 256.663
R2116 B.n679 B.n515 256.663
R2117 B.n685 B.n515 256.663
R2118 B.n687 B.n515 256.663
R2119 B.n693 B.n515 256.663
R2120 B.n695 B.n515 256.663
R2121 B.n701 B.n515 256.663
R2122 B.n703 B.n515 256.663
R2123 B.n709 B.n515 256.663
R2124 B.n711 B.n515 256.663
R2125 B.n718 B.n515 256.663
R2126 B.n720 B.n515 256.663
R2127 B.n726 B.n515 256.663
R2128 B.n728 B.n515 256.663
R2129 B.n737 B.n515 256.663
R2130 B.n739 B.n515 256.663
R2131 B.n745 B.n515 256.663
R2132 B.n747 B.n515 256.663
R2133 B.n753 B.n515 256.663
R2134 B.n755 B.n515 256.663
R2135 B.n761 B.n515 256.663
R2136 B.n763 B.n515 256.663
R2137 B.n769 B.n515 256.663
R2138 B.n771 B.n515 256.663
R2139 B.n777 B.n515 256.663
R2140 B.n779 B.n515 256.663
R2141 B.n785 B.n515 256.663
R2142 B.n787 B.n515 256.663
R2143 B.n793 B.n515 256.663
R2144 B.n795 B.n515 256.663
R2145 B.n801 B.n515 256.663
R2146 B.n803 B.n515 256.663
R2147 B.n809 B.n515 256.663
R2148 B.n811 B.n515 256.663
R2149 B.n817 B.n515 256.663
R2150 B.n819 B.n515 256.663
R2151 B.n825 B.n515 256.663
R2152 B.n827 B.n515 256.663
R2153 B.n833 B.n515 256.663
R2154 B.n835 B.n515 256.663
R2155 B.n841 B.n515 256.663
R2156 B.n843 B.n515 256.663
R2157 B.n849 B.n515 256.663
R2158 B.n851 B.n515 256.663
R2159 B.n857 B.n515 256.663
R2160 B.n860 B.n515 256.663
R2161 B.n1152 B.n1151 256.663
R2162 B.n161 B.n160 163.367
R2163 B.n165 B.n164 163.367
R2164 B.n169 B.n168 163.367
R2165 B.n173 B.n172 163.367
R2166 B.n177 B.n176 163.367
R2167 B.n181 B.n180 163.367
R2168 B.n185 B.n184 163.367
R2169 B.n189 B.n188 163.367
R2170 B.n193 B.n192 163.367
R2171 B.n197 B.n196 163.367
R2172 B.n201 B.n200 163.367
R2173 B.n205 B.n204 163.367
R2174 B.n209 B.n208 163.367
R2175 B.n213 B.n212 163.367
R2176 B.n217 B.n216 163.367
R2177 B.n221 B.n220 163.367
R2178 B.n225 B.n224 163.367
R2179 B.n229 B.n228 163.367
R2180 B.n233 B.n232 163.367
R2181 B.n237 B.n236 163.367
R2182 B.n241 B.n240 163.367
R2183 B.n245 B.n244 163.367
R2184 B.n249 B.n248 163.367
R2185 B.n253 B.n252 163.367
R2186 B.n257 B.n256 163.367
R2187 B.n261 B.n260 163.367
R2188 B.n265 B.n264 163.367
R2189 B.n269 B.n268 163.367
R2190 B.n273 B.n272 163.367
R2191 B.n277 B.n276 163.367
R2192 B.n281 B.n280 163.367
R2193 B.n285 B.n284 163.367
R2194 B.n289 B.n288 163.367
R2195 B.n293 B.n292 163.367
R2196 B.n297 B.n296 163.367
R2197 B.n301 B.n300 163.367
R2198 B.n305 B.n304 163.367
R2199 B.n309 B.n308 163.367
R2200 B.n313 B.n312 163.367
R2201 B.n317 B.n316 163.367
R2202 B.n321 B.n320 163.367
R2203 B.n325 B.n324 163.367
R2204 B.n329 B.n328 163.367
R2205 B.n333 B.n332 163.367
R2206 B.n337 B.n336 163.367
R2207 B.n341 B.n340 163.367
R2208 B.n345 B.n344 163.367
R2209 B.n349 B.n348 163.367
R2210 B.n353 B.n352 163.367
R2211 B.n357 B.n356 163.367
R2212 B.n361 B.n360 163.367
R2213 B.n365 B.n364 163.367
R2214 B.n369 B.n368 163.367
R2215 B.n373 B.n372 163.367
R2216 B.n377 B.n376 163.367
R2217 B.n381 B.n380 163.367
R2218 B.n385 B.n384 163.367
R2219 B.n389 B.n388 163.367
R2220 B.n393 B.n392 163.367
R2221 B.n397 B.n396 163.367
R2222 B.n401 B.n400 163.367
R2223 B.n405 B.n404 163.367
R2224 B.n409 B.n408 163.367
R2225 B.n413 B.n412 163.367
R2226 B.n417 B.n416 163.367
R2227 B.n421 B.n420 163.367
R2228 B.n425 B.n424 163.367
R2229 B.n427 B.n152 163.367
R2230 B.n865 B.n510 163.367
R2231 B.n873 B.n510 163.367
R2232 B.n873 B.n508 163.367
R2233 B.n877 B.n508 163.367
R2234 B.n877 B.n502 163.367
R2235 B.n885 B.n502 163.367
R2236 B.n885 B.n500 163.367
R2237 B.n889 B.n500 163.367
R2238 B.n889 B.n495 163.367
R2239 B.n898 B.n495 163.367
R2240 B.n898 B.n493 163.367
R2241 B.n902 B.n493 163.367
R2242 B.n902 B.n487 163.367
R2243 B.n910 B.n487 163.367
R2244 B.n910 B.n485 163.367
R2245 B.n914 B.n485 163.367
R2246 B.n914 B.n479 163.367
R2247 B.n922 B.n479 163.367
R2248 B.n922 B.n477 163.367
R2249 B.n926 B.n477 163.367
R2250 B.n926 B.n471 163.367
R2251 B.n934 B.n471 163.367
R2252 B.n934 B.n469 163.367
R2253 B.n938 B.n469 163.367
R2254 B.n938 B.n463 163.367
R2255 B.n946 B.n463 163.367
R2256 B.n946 B.n461 163.367
R2257 B.n950 B.n461 163.367
R2258 B.n950 B.n455 163.367
R2259 B.n958 B.n455 163.367
R2260 B.n958 B.n453 163.367
R2261 B.n962 B.n453 163.367
R2262 B.n962 B.n447 163.367
R2263 B.n970 B.n447 163.367
R2264 B.n970 B.n445 163.367
R2265 B.n974 B.n445 163.367
R2266 B.n974 B.n439 163.367
R2267 B.n982 B.n439 163.367
R2268 B.n982 B.n437 163.367
R2269 B.n987 B.n437 163.367
R2270 B.n987 B.n431 163.367
R2271 B.n995 B.n431 163.367
R2272 B.n996 B.n995 163.367
R2273 B.n996 B.n5 163.367
R2274 B.n6 B.n5 163.367
R2275 B.n7 B.n6 163.367
R2276 B.n1002 B.n7 163.367
R2277 B.n1003 B.n1002 163.367
R2278 B.n1003 B.n13 163.367
R2279 B.n14 B.n13 163.367
R2280 B.n15 B.n14 163.367
R2281 B.n1008 B.n15 163.367
R2282 B.n1008 B.n20 163.367
R2283 B.n21 B.n20 163.367
R2284 B.n22 B.n21 163.367
R2285 B.n1013 B.n22 163.367
R2286 B.n1013 B.n27 163.367
R2287 B.n28 B.n27 163.367
R2288 B.n29 B.n28 163.367
R2289 B.n1018 B.n29 163.367
R2290 B.n1018 B.n34 163.367
R2291 B.n35 B.n34 163.367
R2292 B.n36 B.n35 163.367
R2293 B.n1023 B.n36 163.367
R2294 B.n1023 B.n41 163.367
R2295 B.n42 B.n41 163.367
R2296 B.n43 B.n42 163.367
R2297 B.n1028 B.n43 163.367
R2298 B.n1028 B.n48 163.367
R2299 B.n49 B.n48 163.367
R2300 B.n50 B.n49 163.367
R2301 B.n1033 B.n50 163.367
R2302 B.n1033 B.n55 163.367
R2303 B.n56 B.n55 163.367
R2304 B.n57 B.n56 163.367
R2305 B.n1038 B.n57 163.367
R2306 B.n1038 B.n62 163.367
R2307 B.n63 B.n62 163.367
R2308 B.n64 B.n63 163.367
R2309 B.n1043 B.n64 163.367
R2310 B.n1043 B.n69 163.367
R2311 B.n70 B.n69 163.367
R2312 B.n71 B.n70 163.367
R2313 B.n1048 B.n71 163.367
R2314 B.n1048 B.n76 163.367
R2315 B.n77 B.n76 163.367
R2316 B.n78 B.n77 163.367
R2317 B.n1053 B.n78 163.367
R2318 B.n1053 B.n83 163.367
R2319 B.n590 B.n589 163.367
R2320 B.n592 B.n590 163.367
R2321 B.n596 B.n585 163.367
R2322 B.n600 B.n598 163.367
R2323 B.n604 B.n583 163.367
R2324 B.n608 B.n606 163.367
R2325 B.n612 B.n581 163.367
R2326 B.n616 B.n614 163.367
R2327 B.n620 B.n579 163.367
R2328 B.n624 B.n622 163.367
R2329 B.n628 B.n577 163.367
R2330 B.n632 B.n630 163.367
R2331 B.n636 B.n575 163.367
R2332 B.n640 B.n638 163.367
R2333 B.n644 B.n573 163.367
R2334 B.n648 B.n646 163.367
R2335 B.n652 B.n571 163.367
R2336 B.n656 B.n654 163.367
R2337 B.n660 B.n569 163.367
R2338 B.n664 B.n662 163.367
R2339 B.n668 B.n567 163.367
R2340 B.n672 B.n670 163.367
R2341 B.n676 B.n565 163.367
R2342 B.n680 B.n678 163.367
R2343 B.n684 B.n563 163.367
R2344 B.n688 B.n686 163.367
R2345 B.n692 B.n561 163.367
R2346 B.n696 B.n694 163.367
R2347 B.n700 B.n559 163.367
R2348 B.n704 B.n702 163.367
R2349 B.n708 B.n557 163.367
R2350 B.n712 B.n710 163.367
R2351 B.n717 B.n553 163.367
R2352 B.n721 B.n719 163.367
R2353 B.n725 B.n551 163.367
R2354 B.n729 B.n727 163.367
R2355 B.n736 B.n549 163.367
R2356 B.n740 B.n738 163.367
R2357 B.n744 B.n547 163.367
R2358 B.n748 B.n746 163.367
R2359 B.n752 B.n545 163.367
R2360 B.n756 B.n754 163.367
R2361 B.n760 B.n543 163.367
R2362 B.n764 B.n762 163.367
R2363 B.n768 B.n541 163.367
R2364 B.n772 B.n770 163.367
R2365 B.n776 B.n539 163.367
R2366 B.n780 B.n778 163.367
R2367 B.n784 B.n537 163.367
R2368 B.n788 B.n786 163.367
R2369 B.n792 B.n535 163.367
R2370 B.n796 B.n794 163.367
R2371 B.n800 B.n533 163.367
R2372 B.n804 B.n802 163.367
R2373 B.n808 B.n531 163.367
R2374 B.n812 B.n810 163.367
R2375 B.n816 B.n529 163.367
R2376 B.n820 B.n818 163.367
R2377 B.n824 B.n527 163.367
R2378 B.n828 B.n826 163.367
R2379 B.n832 B.n525 163.367
R2380 B.n836 B.n834 163.367
R2381 B.n840 B.n523 163.367
R2382 B.n844 B.n842 163.367
R2383 B.n848 B.n521 163.367
R2384 B.n852 B.n850 163.367
R2385 B.n856 B.n519 163.367
R2386 B.n859 B.n858 163.367
R2387 B.n861 B.n516 163.367
R2388 B.n867 B.n512 163.367
R2389 B.n871 B.n512 163.367
R2390 B.n871 B.n506 163.367
R2391 B.n879 B.n506 163.367
R2392 B.n879 B.n504 163.367
R2393 B.n883 B.n504 163.367
R2394 B.n883 B.n498 163.367
R2395 B.n892 B.n498 163.367
R2396 B.n892 B.n496 163.367
R2397 B.n896 B.n496 163.367
R2398 B.n896 B.n491 163.367
R2399 B.n904 B.n491 163.367
R2400 B.n904 B.n489 163.367
R2401 B.n908 B.n489 163.367
R2402 B.n908 B.n483 163.367
R2403 B.n916 B.n483 163.367
R2404 B.n916 B.n481 163.367
R2405 B.n920 B.n481 163.367
R2406 B.n920 B.n475 163.367
R2407 B.n928 B.n475 163.367
R2408 B.n928 B.n473 163.367
R2409 B.n932 B.n473 163.367
R2410 B.n932 B.n467 163.367
R2411 B.n940 B.n467 163.367
R2412 B.n940 B.n465 163.367
R2413 B.n944 B.n465 163.367
R2414 B.n944 B.n459 163.367
R2415 B.n952 B.n459 163.367
R2416 B.n952 B.n457 163.367
R2417 B.n956 B.n457 163.367
R2418 B.n956 B.n451 163.367
R2419 B.n964 B.n451 163.367
R2420 B.n964 B.n449 163.367
R2421 B.n968 B.n449 163.367
R2422 B.n968 B.n443 163.367
R2423 B.n976 B.n443 163.367
R2424 B.n976 B.n441 163.367
R2425 B.n980 B.n441 163.367
R2426 B.n980 B.n435 163.367
R2427 B.n989 B.n435 163.367
R2428 B.n989 B.n433 163.367
R2429 B.n993 B.n433 163.367
R2430 B.n993 B.n3 163.367
R2431 B.n1150 B.n3 163.367
R2432 B.n1146 B.n2 163.367
R2433 B.n1146 B.n1145 163.367
R2434 B.n1145 B.n9 163.367
R2435 B.n1141 B.n9 163.367
R2436 B.n1141 B.n11 163.367
R2437 B.n1137 B.n11 163.367
R2438 B.n1137 B.n17 163.367
R2439 B.n1133 B.n17 163.367
R2440 B.n1133 B.n19 163.367
R2441 B.n1129 B.n19 163.367
R2442 B.n1129 B.n24 163.367
R2443 B.n1125 B.n24 163.367
R2444 B.n1125 B.n26 163.367
R2445 B.n1121 B.n26 163.367
R2446 B.n1121 B.n31 163.367
R2447 B.n1117 B.n31 163.367
R2448 B.n1117 B.n33 163.367
R2449 B.n1113 B.n33 163.367
R2450 B.n1113 B.n38 163.367
R2451 B.n1109 B.n38 163.367
R2452 B.n1109 B.n40 163.367
R2453 B.n1105 B.n40 163.367
R2454 B.n1105 B.n45 163.367
R2455 B.n1101 B.n45 163.367
R2456 B.n1101 B.n47 163.367
R2457 B.n1097 B.n47 163.367
R2458 B.n1097 B.n52 163.367
R2459 B.n1093 B.n52 163.367
R2460 B.n1093 B.n54 163.367
R2461 B.n1089 B.n54 163.367
R2462 B.n1089 B.n59 163.367
R2463 B.n1085 B.n59 163.367
R2464 B.n1085 B.n61 163.367
R2465 B.n1081 B.n61 163.367
R2466 B.n1081 B.n65 163.367
R2467 B.n1077 B.n65 163.367
R2468 B.n1077 B.n67 163.367
R2469 B.n1073 B.n67 163.367
R2470 B.n1073 B.n73 163.367
R2471 B.n1069 B.n73 163.367
R2472 B.n1069 B.n75 163.367
R2473 B.n1065 B.n75 163.367
R2474 B.n1065 B.n80 163.367
R2475 B.n1061 B.n80 163.367
R2476 B.n157 B.n156 79.7096
R2477 B.n154 B.n153 79.7096
R2478 B.n733 B.n732 79.7096
R2479 B.n555 B.n554 79.7096
R2480 B.n84 B.n82 71.676
R2481 B.n161 B.n85 71.676
R2482 B.n165 B.n86 71.676
R2483 B.n169 B.n87 71.676
R2484 B.n173 B.n88 71.676
R2485 B.n177 B.n89 71.676
R2486 B.n181 B.n90 71.676
R2487 B.n185 B.n91 71.676
R2488 B.n189 B.n92 71.676
R2489 B.n193 B.n93 71.676
R2490 B.n197 B.n94 71.676
R2491 B.n201 B.n95 71.676
R2492 B.n205 B.n96 71.676
R2493 B.n209 B.n97 71.676
R2494 B.n213 B.n98 71.676
R2495 B.n217 B.n99 71.676
R2496 B.n221 B.n100 71.676
R2497 B.n225 B.n101 71.676
R2498 B.n229 B.n102 71.676
R2499 B.n233 B.n103 71.676
R2500 B.n237 B.n104 71.676
R2501 B.n241 B.n105 71.676
R2502 B.n245 B.n106 71.676
R2503 B.n249 B.n107 71.676
R2504 B.n253 B.n108 71.676
R2505 B.n257 B.n109 71.676
R2506 B.n261 B.n110 71.676
R2507 B.n265 B.n111 71.676
R2508 B.n269 B.n112 71.676
R2509 B.n273 B.n113 71.676
R2510 B.n277 B.n114 71.676
R2511 B.n281 B.n115 71.676
R2512 B.n285 B.n116 71.676
R2513 B.n289 B.n117 71.676
R2514 B.n293 B.n118 71.676
R2515 B.n297 B.n119 71.676
R2516 B.n301 B.n120 71.676
R2517 B.n305 B.n121 71.676
R2518 B.n309 B.n122 71.676
R2519 B.n313 B.n123 71.676
R2520 B.n317 B.n124 71.676
R2521 B.n321 B.n125 71.676
R2522 B.n325 B.n126 71.676
R2523 B.n329 B.n127 71.676
R2524 B.n333 B.n128 71.676
R2525 B.n337 B.n129 71.676
R2526 B.n341 B.n130 71.676
R2527 B.n345 B.n131 71.676
R2528 B.n349 B.n132 71.676
R2529 B.n353 B.n133 71.676
R2530 B.n357 B.n134 71.676
R2531 B.n361 B.n135 71.676
R2532 B.n365 B.n136 71.676
R2533 B.n369 B.n137 71.676
R2534 B.n373 B.n138 71.676
R2535 B.n377 B.n139 71.676
R2536 B.n381 B.n140 71.676
R2537 B.n385 B.n141 71.676
R2538 B.n389 B.n142 71.676
R2539 B.n393 B.n143 71.676
R2540 B.n397 B.n144 71.676
R2541 B.n401 B.n145 71.676
R2542 B.n405 B.n146 71.676
R2543 B.n409 B.n147 71.676
R2544 B.n413 B.n148 71.676
R2545 B.n417 B.n149 71.676
R2546 B.n421 B.n150 71.676
R2547 B.n425 B.n151 71.676
R2548 B.n1058 B.n152 71.676
R2549 B.n1058 B.n1057 71.676
R2550 B.n427 B.n151 71.676
R2551 B.n424 B.n150 71.676
R2552 B.n420 B.n149 71.676
R2553 B.n416 B.n148 71.676
R2554 B.n412 B.n147 71.676
R2555 B.n408 B.n146 71.676
R2556 B.n404 B.n145 71.676
R2557 B.n400 B.n144 71.676
R2558 B.n396 B.n143 71.676
R2559 B.n392 B.n142 71.676
R2560 B.n388 B.n141 71.676
R2561 B.n384 B.n140 71.676
R2562 B.n380 B.n139 71.676
R2563 B.n376 B.n138 71.676
R2564 B.n372 B.n137 71.676
R2565 B.n368 B.n136 71.676
R2566 B.n364 B.n135 71.676
R2567 B.n360 B.n134 71.676
R2568 B.n356 B.n133 71.676
R2569 B.n352 B.n132 71.676
R2570 B.n348 B.n131 71.676
R2571 B.n344 B.n130 71.676
R2572 B.n340 B.n129 71.676
R2573 B.n336 B.n128 71.676
R2574 B.n332 B.n127 71.676
R2575 B.n328 B.n126 71.676
R2576 B.n324 B.n125 71.676
R2577 B.n320 B.n124 71.676
R2578 B.n316 B.n123 71.676
R2579 B.n312 B.n122 71.676
R2580 B.n308 B.n121 71.676
R2581 B.n304 B.n120 71.676
R2582 B.n300 B.n119 71.676
R2583 B.n296 B.n118 71.676
R2584 B.n292 B.n117 71.676
R2585 B.n288 B.n116 71.676
R2586 B.n284 B.n115 71.676
R2587 B.n280 B.n114 71.676
R2588 B.n276 B.n113 71.676
R2589 B.n272 B.n112 71.676
R2590 B.n268 B.n111 71.676
R2591 B.n264 B.n110 71.676
R2592 B.n260 B.n109 71.676
R2593 B.n256 B.n108 71.676
R2594 B.n252 B.n107 71.676
R2595 B.n248 B.n106 71.676
R2596 B.n244 B.n105 71.676
R2597 B.n240 B.n104 71.676
R2598 B.n236 B.n103 71.676
R2599 B.n232 B.n102 71.676
R2600 B.n228 B.n101 71.676
R2601 B.n224 B.n100 71.676
R2602 B.n220 B.n99 71.676
R2603 B.n216 B.n98 71.676
R2604 B.n212 B.n97 71.676
R2605 B.n208 B.n96 71.676
R2606 B.n204 B.n95 71.676
R2607 B.n200 B.n94 71.676
R2608 B.n196 B.n93 71.676
R2609 B.n192 B.n92 71.676
R2610 B.n188 B.n91 71.676
R2611 B.n184 B.n90 71.676
R2612 B.n180 B.n89 71.676
R2613 B.n176 B.n88 71.676
R2614 B.n172 B.n87 71.676
R2615 B.n168 B.n86 71.676
R2616 B.n164 B.n85 71.676
R2617 B.n160 B.n84 71.676
R2618 B.n588 B.n514 71.676
R2619 B.n592 B.n591 71.676
R2620 B.n597 B.n596 71.676
R2621 B.n600 B.n599 71.676
R2622 B.n605 B.n604 71.676
R2623 B.n608 B.n607 71.676
R2624 B.n613 B.n612 71.676
R2625 B.n616 B.n615 71.676
R2626 B.n621 B.n620 71.676
R2627 B.n624 B.n623 71.676
R2628 B.n629 B.n628 71.676
R2629 B.n632 B.n631 71.676
R2630 B.n637 B.n636 71.676
R2631 B.n640 B.n639 71.676
R2632 B.n645 B.n644 71.676
R2633 B.n648 B.n647 71.676
R2634 B.n653 B.n652 71.676
R2635 B.n656 B.n655 71.676
R2636 B.n661 B.n660 71.676
R2637 B.n664 B.n663 71.676
R2638 B.n669 B.n668 71.676
R2639 B.n672 B.n671 71.676
R2640 B.n677 B.n676 71.676
R2641 B.n680 B.n679 71.676
R2642 B.n685 B.n684 71.676
R2643 B.n688 B.n687 71.676
R2644 B.n693 B.n692 71.676
R2645 B.n696 B.n695 71.676
R2646 B.n701 B.n700 71.676
R2647 B.n704 B.n703 71.676
R2648 B.n709 B.n708 71.676
R2649 B.n712 B.n711 71.676
R2650 B.n718 B.n717 71.676
R2651 B.n721 B.n720 71.676
R2652 B.n726 B.n725 71.676
R2653 B.n729 B.n728 71.676
R2654 B.n737 B.n736 71.676
R2655 B.n740 B.n739 71.676
R2656 B.n745 B.n744 71.676
R2657 B.n748 B.n747 71.676
R2658 B.n753 B.n752 71.676
R2659 B.n756 B.n755 71.676
R2660 B.n761 B.n760 71.676
R2661 B.n764 B.n763 71.676
R2662 B.n769 B.n768 71.676
R2663 B.n772 B.n771 71.676
R2664 B.n777 B.n776 71.676
R2665 B.n780 B.n779 71.676
R2666 B.n785 B.n784 71.676
R2667 B.n788 B.n787 71.676
R2668 B.n793 B.n792 71.676
R2669 B.n796 B.n795 71.676
R2670 B.n801 B.n800 71.676
R2671 B.n804 B.n803 71.676
R2672 B.n809 B.n808 71.676
R2673 B.n812 B.n811 71.676
R2674 B.n817 B.n816 71.676
R2675 B.n820 B.n819 71.676
R2676 B.n825 B.n824 71.676
R2677 B.n828 B.n827 71.676
R2678 B.n833 B.n832 71.676
R2679 B.n836 B.n835 71.676
R2680 B.n841 B.n840 71.676
R2681 B.n844 B.n843 71.676
R2682 B.n849 B.n848 71.676
R2683 B.n852 B.n851 71.676
R2684 B.n857 B.n856 71.676
R2685 B.n860 B.n859 71.676
R2686 B.n589 B.n588 71.676
R2687 B.n591 B.n585 71.676
R2688 B.n598 B.n597 71.676
R2689 B.n599 B.n583 71.676
R2690 B.n606 B.n605 71.676
R2691 B.n607 B.n581 71.676
R2692 B.n614 B.n613 71.676
R2693 B.n615 B.n579 71.676
R2694 B.n622 B.n621 71.676
R2695 B.n623 B.n577 71.676
R2696 B.n630 B.n629 71.676
R2697 B.n631 B.n575 71.676
R2698 B.n638 B.n637 71.676
R2699 B.n639 B.n573 71.676
R2700 B.n646 B.n645 71.676
R2701 B.n647 B.n571 71.676
R2702 B.n654 B.n653 71.676
R2703 B.n655 B.n569 71.676
R2704 B.n662 B.n661 71.676
R2705 B.n663 B.n567 71.676
R2706 B.n670 B.n669 71.676
R2707 B.n671 B.n565 71.676
R2708 B.n678 B.n677 71.676
R2709 B.n679 B.n563 71.676
R2710 B.n686 B.n685 71.676
R2711 B.n687 B.n561 71.676
R2712 B.n694 B.n693 71.676
R2713 B.n695 B.n559 71.676
R2714 B.n702 B.n701 71.676
R2715 B.n703 B.n557 71.676
R2716 B.n710 B.n709 71.676
R2717 B.n711 B.n553 71.676
R2718 B.n719 B.n718 71.676
R2719 B.n720 B.n551 71.676
R2720 B.n727 B.n726 71.676
R2721 B.n728 B.n549 71.676
R2722 B.n738 B.n737 71.676
R2723 B.n739 B.n547 71.676
R2724 B.n746 B.n745 71.676
R2725 B.n747 B.n545 71.676
R2726 B.n754 B.n753 71.676
R2727 B.n755 B.n543 71.676
R2728 B.n762 B.n761 71.676
R2729 B.n763 B.n541 71.676
R2730 B.n770 B.n769 71.676
R2731 B.n771 B.n539 71.676
R2732 B.n778 B.n777 71.676
R2733 B.n779 B.n537 71.676
R2734 B.n786 B.n785 71.676
R2735 B.n787 B.n535 71.676
R2736 B.n794 B.n793 71.676
R2737 B.n795 B.n533 71.676
R2738 B.n802 B.n801 71.676
R2739 B.n803 B.n531 71.676
R2740 B.n810 B.n809 71.676
R2741 B.n811 B.n529 71.676
R2742 B.n818 B.n817 71.676
R2743 B.n819 B.n527 71.676
R2744 B.n826 B.n825 71.676
R2745 B.n827 B.n525 71.676
R2746 B.n834 B.n833 71.676
R2747 B.n835 B.n523 71.676
R2748 B.n842 B.n841 71.676
R2749 B.n843 B.n521 71.676
R2750 B.n850 B.n849 71.676
R2751 B.n851 B.n519 71.676
R2752 B.n858 B.n857 71.676
R2753 B.n861 B.n860 71.676
R2754 B.n1151 B.n1150 71.676
R2755 B.n1151 B.n2 71.676
R2756 B.n158 B.n157 59.5399
R2757 B.n155 B.n154 59.5399
R2758 B.n734 B.n733 59.5399
R2759 B.n714 B.n555 59.5399
R2760 B.n866 B.n515 50.7121
R2761 B.n1060 B.n1059 50.7121
R2762 B.n868 B.n513 30.7517
R2763 B.n864 B.n863 30.7517
R2764 B.n1056 B.n1055 30.7517
R2765 B.n1062 B.n81 30.7517
R2766 B.n866 B.n511 29.9865
R2767 B.n872 B.n511 29.9865
R2768 B.n872 B.n507 29.9865
R2769 B.n878 B.n507 29.9865
R2770 B.n878 B.n503 29.9865
R2771 B.n884 B.n503 29.9865
R2772 B.n884 B.n499 29.9865
R2773 B.n891 B.n499 29.9865
R2774 B.n891 B.n890 29.9865
R2775 B.n897 B.n492 29.9865
R2776 B.n903 B.n492 29.9865
R2777 B.n903 B.n488 29.9865
R2778 B.n909 B.n488 29.9865
R2779 B.n909 B.n484 29.9865
R2780 B.n915 B.n484 29.9865
R2781 B.n915 B.n480 29.9865
R2782 B.n921 B.n480 29.9865
R2783 B.n921 B.n476 29.9865
R2784 B.n927 B.n476 29.9865
R2785 B.n927 B.n472 29.9865
R2786 B.n933 B.n472 29.9865
R2787 B.n933 B.n468 29.9865
R2788 B.n939 B.n468 29.9865
R2789 B.n945 B.n464 29.9865
R2790 B.n945 B.n460 29.9865
R2791 B.n951 B.n460 29.9865
R2792 B.n951 B.n456 29.9865
R2793 B.n957 B.n456 29.9865
R2794 B.n957 B.n452 29.9865
R2795 B.n963 B.n452 29.9865
R2796 B.n963 B.n448 29.9865
R2797 B.n969 B.n448 29.9865
R2798 B.n969 B.n444 29.9865
R2799 B.n975 B.n444 29.9865
R2800 B.n981 B.n440 29.9865
R2801 B.n981 B.n436 29.9865
R2802 B.n988 B.n436 29.9865
R2803 B.n988 B.n432 29.9865
R2804 B.n994 B.n432 29.9865
R2805 B.n994 B.n4 29.9865
R2806 B.n1149 B.n4 29.9865
R2807 B.n1149 B.n1148 29.9865
R2808 B.n1148 B.n1147 29.9865
R2809 B.n1147 B.n8 29.9865
R2810 B.n12 B.n8 29.9865
R2811 B.n1140 B.n12 29.9865
R2812 B.n1140 B.n1139 29.9865
R2813 B.n1139 B.n1138 29.9865
R2814 B.n1138 B.n16 29.9865
R2815 B.n1132 B.n1131 29.9865
R2816 B.n1131 B.n1130 29.9865
R2817 B.n1130 B.n23 29.9865
R2818 B.n1124 B.n23 29.9865
R2819 B.n1124 B.n1123 29.9865
R2820 B.n1123 B.n1122 29.9865
R2821 B.n1122 B.n30 29.9865
R2822 B.n1116 B.n30 29.9865
R2823 B.n1116 B.n1115 29.9865
R2824 B.n1115 B.n1114 29.9865
R2825 B.n1114 B.n37 29.9865
R2826 B.n1108 B.n1107 29.9865
R2827 B.n1107 B.n1106 29.9865
R2828 B.n1106 B.n44 29.9865
R2829 B.n1100 B.n44 29.9865
R2830 B.n1100 B.n1099 29.9865
R2831 B.n1099 B.n1098 29.9865
R2832 B.n1098 B.n51 29.9865
R2833 B.n1092 B.n51 29.9865
R2834 B.n1092 B.n1091 29.9865
R2835 B.n1091 B.n1090 29.9865
R2836 B.n1090 B.n58 29.9865
R2837 B.n1084 B.n58 29.9865
R2838 B.n1084 B.n1083 29.9865
R2839 B.n1083 B.n1082 29.9865
R2840 B.n1076 B.n68 29.9865
R2841 B.n1076 B.n1075 29.9865
R2842 B.n1075 B.n1074 29.9865
R2843 B.n1074 B.n72 29.9865
R2844 B.n1068 B.n72 29.9865
R2845 B.n1068 B.n1067 29.9865
R2846 B.n1067 B.n1066 29.9865
R2847 B.n1066 B.n79 29.9865
R2848 B.n1060 B.n79 29.9865
R2849 B.n975 B.t3 25.5768
R2850 B.n1132 B.t2 25.5768
R2851 B.n939 B.t1 22.9309
R2852 B.n1108 B.t0 22.9309
R2853 B B.n1152 18.0485
R2854 B.n897 B.t12 15.8754
R2855 B.n1082 B.t5 15.8754
R2856 B.n890 B.t12 14.1115
R2857 B.n68 B.t5 14.1115
R2858 B.n869 B.n868 10.6151
R2859 B.n870 B.n869 10.6151
R2860 B.n870 B.n505 10.6151
R2861 B.n880 B.n505 10.6151
R2862 B.n881 B.n880 10.6151
R2863 B.n882 B.n881 10.6151
R2864 B.n882 B.n497 10.6151
R2865 B.n893 B.n497 10.6151
R2866 B.n894 B.n893 10.6151
R2867 B.n895 B.n894 10.6151
R2868 B.n895 B.n490 10.6151
R2869 B.n905 B.n490 10.6151
R2870 B.n906 B.n905 10.6151
R2871 B.n907 B.n906 10.6151
R2872 B.n907 B.n482 10.6151
R2873 B.n917 B.n482 10.6151
R2874 B.n918 B.n917 10.6151
R2875 B.n919 B.n918 10.6151
R2876 B.n919 B.n474 10.6151
R2877 B.n929 B.n474 10.6151
R2878 B.n930 B.n929 10.6151
R2879 B.n931 B.n930 10.6151
R2880 B.n931 B.n466 10.6151
R2881 B.n941 B.n466 10.6151
R2882 B.n942 B.n941 10.6151
R2883 B.n943 B.n942 10.6151
R2884 B.n943 B.n458 10.6151
R2885 B.n953 B.n458 10.6151
R2886 B.n954 B.n953 10.6151
R2887 B.n955 B.n954 10.6151
R2888 B.n955 B.n450 10.6151
R2889 B.n965 B.n450 10.6151
R2890 B.n966 B.n965 10.6151
R2891 B.n967 B.n966 10.6151
R2892 B.n967 B.n442 10.6151
R2893 B.n977 B.n442 10.6151
R2894 B.n978 B.n977 10.6151
R2895 B.n979 B.n978 10.6151
R2896 B.n979 B.n434 10.6151
R2897 B.n990 B.n434 10.6151
R2898 B.n991 B.n990 10.6151
R2899 B.n992 B.n991 10.6151
R2900 B.n992 B.n0 10.6151
R2901 B.n587 B.n513 10.6151
R2902 B.n587 B.n586 10.6151
R2903 B.n593 B.n586 10.6151
R2904 B.n594 B.n593 10.6151
R2905 B.n595 B.n594 10.6151
R2906 B.n595 B.n584 10.6151
R2907 B.n601 B.n584 10.6151
R2908 B.n602 B.n601 10.6151
R2909 B.n603 B.n602 10.6151
R2910 B.n603 B.n582 10.6151
R2911 B.n609 B.n582 10.6151
R2912 B.n610 B.n609 10.6151
R2913 B.n611 B.n610 10.6151
R2914 B.n611 B.n580 10.6151
R2915 B.n617 B.n580 10.6151
R2916 B.n618 B.n617 10.6151
R2917 B.n619 B.n618 10.6151
R2918 B.n619 B.n578 10.6151
R2919 B.n625 B.n578 10.6151
R2920 B.n626 B.n625 10.6151
R2921 B.n627 B.n626 10.6151
R2922 B.n627 B.n576 10.6151
R2923 B.n633 B.n576 10.6151
R2924 B.n634 B.n633 10.6151
R2925 B.n635 B.n634 10.6151
R2926 B.n635 B.n574 10.6151
R2927 B.n641 B.n574 10.6151
R2928 B.n642 B.n641 10.6151
R2929 B.n643 B.n642 10.6151
R2930 B.n643 B.n572 10.6151
R2931 B.n649 B.n572 10.6151
R2932 B.n650 B.n649 10.6151
R2933 B.n651 B.n650 10.6151
R2934 B.n651 B.n570 10.6151
R2935 B.n657 B.n570 10.6151
R2936 B.n658 B.n657 10.6151
R2937 B.n659 B.n658 10.6151
R2938 B.n659 B.n568 10.6151
R2939 B.n665 B.n568 10.6151
R2940 B.n666 B.n665 10.6151
R2941 B.n667 B.n666 10.6151
R2942 B.n667 B.n566 10.6151
R2943 B.n673 B.n566 10.6151
R2944 B.n674 B.n673 10.6151
R2945 B.n675 B.n674 10.6151
R2946 B.n675 B.n564 10.6151
R2947 B.n681 B.n564 10.6151
R2948 B.n682 B.n681 10.6151
R2949 B.n683 B.n682 10.6151
R2950 B.n683 B.n562 10.6151
R2951 B.n689 B.n562 10.6151
R2952 B.n690 B.n689 10.6151
R2953 B.n691 B.n690 10.6151
R2954 B.n691 B.n560 10.6151
R2955 B.n697 B.n560 10.6151
R2956 B.n698 B.n697 10.6151
R2957 B.n699 B.n698 10.6151
R2958 B.n699 B.n558 10.6151
R2959 B.n705 B.n558 10.6151
R2960 B.n706 B.n705 10.6151
R2961 B.n707 B.n706 10.6151
R2962 B.n707 B.n556 10.6151
R2963 B.n713 B.n556 10.6151
R2964 B.n716 B.n715 10.6151
R2965 B.n716 B.n552 10.6151
R2966 B.n722 B.n552 10.6151
R2967 B.n723 B.n722 10.6151
R2968 B.n724 B.n723 10.6151
R2969 B.n724 B.n550 10.6151
R2970 B.n730 B.n550 10.6151
R2971 B.n731 B.n730 10.6151
R2972 B.n735 B.n731 10.6151
R2973 B.n741 B.n548 10.6151
R2974 B.n742 B.n741 10.6151
R2975 B.n743 B.n742 10.6151
R2976 B.n743 B.n546 10.6151
R2977 B.n749 B.n546 10.6151
R2978 B.n750 B.n749 10.6151
R2979 B.n751 B.n750 10.6151
R2980 B.n751 B.n544 10.6151
R2981 B.n757 B.n544 10.6151
R2982 B.n758 B.n757 10.6151
R2983 B.n759 B.n758 10.6151
R2984 B.n759 B.n542 10.6151
R2985 B.n765 B.n542 10.6151
R2986 B.n766 B.n765 10.6151
R2987 B.n767 B.n766 10.6151
R2988 B.n767 B.n540 10.6151
R2989 B.n773 B.n540 10.6151
R2990 B.n774 B.n773 10.6151
R2991 B.n775 B.n774 10.6151
R2992 B.n775 B.n538 10.6151
R2993 B.n781 B.n538 10.6151
R2994 B.n782 B.n781 10.6151
R2995 B.n783 B.n782 10.6151
R2996 B.n783 B.n536 10.6151
R2997 B.n789 B.n536 10.6151
R2998 B.n790 B.n789 10.6151
R2999 B.n791 B.n790 10.6151
R3000 B.n791 B.n534 10.6151
R3001 B.n797 B.n534 10.6151
R3002 B.n798 B.n797 10.6151
R3003 B.n799 B.n798 10.6151
R3004 B.n799 B.n532 10.6151
R3005 B.n805 B.n532 10.6151
R3006 B.n806 B.n805 10.6151
R3007 B.n807 B.n806 10.6151
R3008 B.n807 B.n530 10.6151
R3009 B.n813 B.n530 10.6151
R3010 B.n814 B.n813 10.6151
R3011 B.n815 B.n814 10.6151
R3012 B.n815 B.n528 10.6151
R3013 B.n821 B.n528 10.6151
R3014 B.n822 B.n821 10.6151
R3015 B.n823 B.n822 10.6151
R3016 B.n823 B.n526 10.6151
R3017 B.n829 B.n526 10.6151
R3018 B.n830 B.n829 10.6151
R3019 B.n831 B.n830 10.6151
R3020 B.n831 B.n524 10.6151
R3021 B.n837 B.n524 10.6151
R3022 B.n838 B.n837 10.6151
R3023 B.n839 B.n838 10.6151
R3024 B.n839 B.n522 10.6151
R3025 B.n845 B.n522 10.6151
R3026 B.n846 B.n845 10.6151
R3027 B.n847 B.n846 10.6151
R3028 B.n847 B.n520 10.6151
R3029 B.n853 B.n520 10.6151
R3030 B.n854 B.n853 10.6151
R3031 B.n855 B.n854 10.6151
R3032 B.n855 B.n518 10.6151
R3033 B.n518 B.n517 10.6151
R3034 B.n862 B.n517 10.6151
R3035 B.n863 B.n862 10.6151
R3036 B.n864 B.n509 10.6151
R3037 B.n874 B.n509 10.6151
R3038 B.n875 B.n874 10.6151
R3039 B.n876 B.n875 10.6151
R3040 B.n876 B.n501 10.6151
R3041 B.n886 B.n501 10.6151
R3042 B.n887 B.n886 10.6151
R3043 B.n888 B.n887 10.6151
R3044 B.n888 B.n494 10.6151
R3045 B.n899 B.n494 10.6151
R3046 B.n900 B.n899 10.6151
R3047 B.n901 B.n900 10.6151
R3048 B.n901 B.n486 10.6151
R3049 B.n911 B.n486 10.6151
R3050 B.n912 B.n911 10.6151
R3051 B.n913 B.n912 10.6151
R3052 B.n913 B.n478 10.6151
R3053 B.n923 B.n478 10.6151
R3054 B.n924 B.n923 10.6151
R3055 B.n925 B.n924 10.6151
R3056 B.n925 B.n470 10.6151
R3057 B.n935 B.n470 10.6151
R3058 B.n936 B.n935 10.6151
R3059 B.n937 B.n936 10.6151
R3060 B.n937 B.n462 10.6151
R3061 B.n947 B.n462 10.6151
R3062 B.n948 B.n947 10.6151
R3063 B.n949 B.n948 10.6151
R3064 B.n949 B.n454 10.6151
R3065 B.n959 B.n454 10.6151
R3066 B.n960 B.n959 10.6151
R3067 B.n961 B.n960 10.6151
R3068 B.n961 B.n446 10.6151
R3069 B.n971 B.n446 10.6151
R3070 B.n972 B.n971 10.6151
R3071 B.n973 B.n972 10.6151
R3072 B.n973 B.n438 10.6151
R3073 B.n983 B.n438 10.6151
R3074 B.n984 B.n983 10.6151
R3075 B.n986 B.n984 10.6151
R3076 B.n986 B.n985 10.6151
R3077 B.n985 B.n430 10.6151
R3078 B.n997 B.n430 10.6151
R3079 B.n998 B.n997 10.6151
R3080 B.n999 B.n998 10.6151
R3081 B.n1000 B.n999 10.6151
R3082 B.n1001 B.n1000 10.6151
R3083 B.n1004 B.n1001 10.6151
R3084 B.n1005 B.n1004 10.6151
R3085 B.n1006 B.n1005 10.6151
R3086 B.n1007 B.n1006 10.6151
R3087 B.n1009 B.n1007 10.6151
R3088 B.n1010 B.n1009 10.6151
R3089 B.n1011 B.n1010 10.6151
R3090 B.n1012 B.n1011 10.6151
R3091 B.n1014 B.n1012 10.6151
R3092 B.n1015 B.n1014 10.6151
R3093 B.n1016 B.n1015 10.6151
R3094 B.n1017 B.n1016 10.6151
R3095 B.n1019 B.n1017 10.6151
R3096 B.n1020 B.n1019 10.6151
R3097 B.n1021 B.n1020 10.6151
R3098 B.n1022 B.n1021 10.6151
R3099 B.n1024 B.n1022 10.6151
R3100 B.n1025 B.n1024 10.6151
R3101 B.n1026 B.n1025 10.6151
R3102 B.n1027 B.n1026 10.6151
R3103 B.n1029 B.n1027 10.6151
R3104 B.n1030 B.n1029 10.6151
R3105 B.n1031 B.n1030 10.6151
R3106 B.n1032 B.n1031 10.6151
R3107 B.n1034 B.n1032 10.6151
R3108 B.n1035 B.n1034 10.6151
R3109 B.n1036 B.n1035 10.6151
R3110 B.n1037 B.n1036 10.6151
R3111 B.n1039 B.n1037 10.6151
R3112 B.n1040 B.n1039 10.6151
R3113 B.n1041 B.n1040 10.6151
R3114 B.n1042 B.n1041 10.6151
R3115 B.n1044 B.n1042 10.6151
R3116 B.n1045 B.n1044 10.6151
R3117 B.n1046 B.n1045 10.6151
R3118 B.n1047 B.n1046 10.6151
R3119 B.n1049 B.n1047 10.6151
R3120 B.n1050 B.n1049 10.6151
R3121 B.n1051 B.n1050 10.6151
R3122 B.n1052 B.n1051 10.6151
R3123 B.n1054 B.n1052 10.6151
R3124 B.n1055 B.n1054 10.6151
R3125 B.n1144 B.n1 10.6151
R3126 B.n1144 B.n1143 10.6151
R3127 B.n1143 B.n1142 10.6151
R3128 B.n1142 B.n10 10.6151
R3129 B.n1136 B.n10 10.6151
R3130 B.n1136 B.n1135 10.6151
R3131 B.n1135 B.n1134 10.6151
R3132 B.n1134 B.n18 10.6151
R3133 B.n1128 B.n18 10.6151
R3134 B.n1128 B.n1127 10.6151
R3135 B.n1127 B.n1126 10.6151
R3136 B.n1126 B.n25 10.6151
R3137 B.n1120 B.n25 10.6151
R3138 B.n1120 B.n1119 10.6151
R3139 B.n1119 B.n1118 10.6151
R3140 B.n1118 B.n32 10.6151
R3141 B.n1112 B.n32 10.6151
R3142 B.n1112 B.n1111 10.6151
R3143 B.n1111 B.n1110 10.6151
R3144 B.n1110 B.n39 10.6151
R3145 B.n1104 B.n39 10.6151
R3146 B.n1104 B.n1103 10.6151
R3147 B.n1103 B.n1102 10.6151
R3148 B.n1102 B.n46 10.6151
R3149 B.n1096 B.n46 10.6151
R3150 B.n1096 B.n1095 10.6151
R3151 B.n1095 B.n1094 10.6151
R3152 B.n1094 B.n53 10.6151
R3153 B.n1088 B.n53 10.6151
R3154 B.n1088 B.n1087 10.6151
R3155 B.n1087 B.n1086 10.6151
R3156 B.n1086 B.n60 10.6151
R3157 B.n1080 B.n60 10.6151
R3158 B.n1080 B.n1079 10.6151
R3159 B.n1079 B.n1078 10.6151
R3160 B.n1078 B.n66 10.6151
R3161 B.n1072 B.n66 10.6151
R3162 B.n1072 B.n1071 10.6151
R3163 B.n1071 B.n1070 10.6151
R3164 B.n1070 B.n74 10.6151
R3165 B.n1064 B.n74 10.6151
R3166 B.n1064 B.n1063 10.6151
R3167 B.n1063 B.n1062 10.6151
R3168 B.n159 B.n81 10.6151
R3169 B.n162 B.n159 10.6151
R3170 B.n163 B.n162 10.6151
R3171 B.n166 B.n163 10.6151
R3172 B.n167 B.n166 10.6151
R3173 B.n170 B.n167 10.6151
R3174 B.n171 B.n170 10.6151
R3175 B.n174 B.n171 10.6151
R3176 B.n175 B.n174 10.6151
R3177 B.n178 B.n175 10.6151
R3178 B.n179 B.n178 10.6151
R3179 B.n182 B.n179 10.6151
R3180 B.n183 B.n182 10.6151
R3181 B.n186 B.n183 10.6151
R3182 B.n187 B.n186 10.6151
R3183 B.n190 B.n187 10.6151
R3184 B.n191 B.n190 10.6151
R3185 B.n194 B.n191 10.6151
R3186 B.n195 B.n194 10.6151
R3187 B.n198 B.n195 10.6151
R3188 B.n199 B.n198 10.6151
R3189 B.n202 B.n199 10.6151
R3190 B.n203 B.n202 10.6151
R3191 B.n206 B.n203 10.6151
R3192 B.n207 B.n206 10.6151
R3193 B.n210 B.n207 10.6151
R3194 B.n211 B.n210 10.6151
R3195 B.n214 B.n211 10.6151
R3196 B.n215 B.n214 10.6151
R3197 B.n218 B.n215 10.6151
R3198 B.n219 B.n218 10.6151
R3199 B.n222 B.n219 10.6151
R3200 B.n223 B.n222 10.6151
R3201 B.n226 B.n223 10.6151
R3202 B.n227 B.n226 10.6151
R3203 B.n230 B.n227 10.6151
R3204 B.n231 B.n230 10.6151
R3205 B.n234 B.n231 10.6151
R3206 B.n235 B.n234 10.6151
R3207 B.n238 B.n235 10.6151
R3208 B.n239 B.n238 10.6151
R3209 B.n242 B.n239 10.6151
R3210 B.n243 B.n242 10.6151
R3211 B.n246 B.n243 10.6151
R3212 B.n247 B.n246 10.6151
R3213 B.n250 B.n247 10.6151
R3214 B.n251 B.n250 10.6151
R3215 B.n254 B.n251 10.6151
R3216 B.n255 B.n254 10.6151
R3217 B.n258 B.n255 10.6151
R3218 B.n259 B.n258 10.6151
R3219 B.n262 B.n259 10.6151
R3220 B.n263 B.n262 10.6151
R3221 B.n266 B.n263 10.6151
R3222 B.n267 B.n266 10.6151
R3223 B.n270 B.n267 10.6151
R3224 B.n271 B.n270 10.6151
R3225 B.n274 B.n271 10.6151
R3226 B.n275 B.n274 10.6151
R3227 B.n278 B.n275 10.6151
R3228 B.n279 B.n278 10.6151
R3229 B.n282 B.n279 10.6151
R3230 B.n283 B.n282 10.6151
R3231 B.n287 B.n286 10.6151
R3232 B.n290 B.n287 10.6151
R3233 B.n291 B.n290 10.6151
R3234 B.n294 B.n291 10.6151
R3235 B.n295 B.n294 10.6151
R3236 B.n298 B.n295 10.6151
R3237 B.n299 B.n298 10.6151
R3238 B.n302 B.n299 10.6151
R3239 B.n303 B.n302 10.6151
R3240 B.n307 B.n306 10.6151
R3241 B.n310 B.n307 10.6151
R3242 B.n311 B.n310 10.6151
R3243 B.n314 B.n311 10.6151
R3244 B.n315 B.n314 10.6151
R3245 B.n318 B.n315 10.6151
R3246 B.n319 B.n318 10.6151
R3247 B.n322 B.n319 10.6151
R3248 B.n323 B.n322 10.6151
R3249 B.n326 B.n323 10.6151
R3250 B.n327 B.n326 10.6151
R3251 B.n330 B.n327 10.6151
R3252 B.n331 B.n330 10.6151
R3253 B.n334 B.n331 10.6151
R3254 B.n335 B.n334 10.6151
R3255 B.n338 B.n335 10.6151
R3256 B.n339 B.n338 10.6151
R3257 B.n342 B.n339 10.6151
R3258 B.n343 B.n342 10.6151
R3259 B.n346 B.n343 10.6151
R3260 B.n347 B.n346 10.6151
R3261 B.n350 B.n347 10.6151
R3262 B.n351 B.n350 10.6151
R3263 B.n354 B.n351 10.6151
R3264 B.n355 B.n354 10.6151
R3265 B.n358 B.n355 10.6151
R3266 B.n359 B.n358 10.6151
R3267 B.n362 B.n359 10.6151
R3268 B.n363 B.n362 10.6151
R3269 B.n366 B.n363 10.6151
R3270 B.n367 B.n366 10.6151
R3271 B.n370 B.n367 10.6151
R3272 B.n371 B.n370 10.6151
R3273 B.n374 B.n371 10.6151
R3274 B.n375 B.n374 10.6151
R3275 B.n378 B.n375 10.6151
R3276 B.n379 B.n378 10.6151
R3277 B.n382 B.n379 10.6151
R3278 B.n383 B.n382 10.6151
R3279 B.n386 B.n383 10.6151
R3280 B.n387 B.n386 10.6151
R3281 B.n390 B.n387 10.6151
R3282 B.n391 B.n390 10.6151
R3283 B.n394 B.n391 10.6151
R3284 B.n395 B.n394 10.6151
R3285 B.n398 B.n395 10.6151
R3286 B.n399 B.n398 10.6151
R3287 B.n402 B.n399 10.6151
R3288 B.n403 B.n402 10.6151
R3289 B.n406 B.n403 10.6151
R3290 B.n407 B.n406 10.6151
R3291 B.n410 B.n407 10.6151
R3292 B.n411 B.n410 10.6151
R3293 B.n414 B.n411 10.6151
R3294 B.n415 B.n414 10.6151
R3295 B.n418 B.n415 10.6151
R3296 B.n419 B.n418 10.6151
R3297 B.n422 B.n419 10.6151
R3298 B.n423 B.n422 10.6151
R3299 B.n426 B.n423 10.6151
R3300 B.n428 B.n426 10.6151
R3301 B.n429 B.n428 10.6151
R3302 B.n1056 B.n429 10.6151
R3303 B.n714 B.n713 9.36635
R3304 B.n734 B.n548 9.36635
R3305 B.n283 B.n158 9.36635
R3306 B.n306 B.n155 9.36635
R3307 B.n1152 B.n0 8.11757
R3308 B.n1152 B.n1 8.11757
R3309 B.t1 B.n464 7.05602
R3310 B.t0 B.n37 7.05602
R3311 B.t3 B.n440 4.4102
R3312 B.t2 B.n16 4.4102
R3313 B.n715 B.n714 1.24928
R3314 B.n735 B.n734 1.24928
R3315 B.n286 B.n158 1.24928
R3316 B.n303 B.n155 1.24928
R3317 VN.n1 VN.t2 159.226
R3318 VN.n0 VN.t1 159.226
R3319 VN.n0 VN.t3 157.88
R3320 VN.n1 VN.t0 157.88
R3321 VN VN.n1 57.8163
R3322 VN VN.n0 1.87307
R3323 VDD2.n2 VDD2.n0 111.71
R3324 VDD2.n2 VDD2.n1 60.408
R3325 VDD2.n1 VDD2.t3 1.00711
R3326 VDD2.n1 VDD2.t1 1.00711
R3327 VDD2.n0 VDD2.t2 1.00711
R3328 VDD2.n0 VDD2.t0 1.00711
R3329 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 8.35676f
C1 VTAIL VN 7.7528f
C2 VDD1 VN 0.149921f
C3 VTAIL VDD1 7.33986f
C4 VDD2 VP 0.469245f
C5 VDD2 VN 8.03847f
C6 VDD2 VTAIL 7.40198f
C7 VDD2 VDD1 1.31245f
C8 VP VN 8.462911f
C9 VTAIL VP 7.76691f
C10 VDD2 B 5.023706f
C11 VDD1 B 10.340321f
C12 VTAIL B 15.3922f
C13 VN B 13.58346f
C14 VP B 11.963607f
C15 VDD2.t2 B 0.413367f
C16 VDD2.t0 B 0.413367f
C17 VDD2.n0 B 4.81649f
C18 VDD2.t3 B 0.413367f
C19 VDD2.t1 B 0.413367f
C20 VDD2.n1 B 3.77767f
C21 VDD2.n2 B 4.84304f
C22 VN.t3 B 4.09144f
C23 VN.t1 B 4.10323f
C24 VN.n0 B 2.5112f
C25 VN.t0 B 4.09144f
C26 VN.t2 B 4.10323f
C27 VN.n1 B 3.90279f
C28 VTAIL.n0 B 0.0226f
C29 VTAIL.n1 B 0.015556f
C30 VTAIL.n2 B 0.008359f
C31 VTAIL.n3 B 0.019758f
C32 VTAIL.n4 B 0.008851f
C33 VTAIL.n5 B 0.015556f
C34 VTAIL.n6 B 0.008359f
C35 VTAIL.n7 B 0.019758f
C36 VTAIL.n8 B 0.008851f
C37 VTAIL.n9 B 0.015556f
C38 VTAIL.n10 B 0.008359f
C39 VTAIL.n11 B 0.019758f
C40 VTAIL.n12 B 0.008605f
C41 VTAIL.n13 B 0.015556f
C42 VTAIL.n14 B 0.008851f
C43 VTAIL.n15 B 0.019758f
C44 VTAIL.n16 B 0.008851f
C45 VTAIL.n17 B 0.015556f
C46 VTAIL.n18 B 0.008359f
C47 VTAIL.n19 B 0.019758f
C48 VTAIL.n20 B 0.008851f
C49 VTAIL.n21 B 0.015556f
C50 VTAIL.n22 B 0.008359f
C51 VTAIL.n23 B 0.019758f
C52 VTAIL.n24 B 0.008851f
C53 VTAIL.n25 B 0.015556f
C54 VTAIL.n26 B 0.008359f
C55 VTAIL.n27 B 0.019758f
C56 VTAIL.n28 B 0.008851f
C57 VTAIL.n29 B 0.015556f
C58 VTAIL.n30 B 0.008359f
C59 VTAIL.n31 B 0.019758f
C60 VTAIL.n32 B 0.008851f
C61 VTAIL.n33 B 1.34505f
C62 VTAIL.n34 B 0.008359f
C63 VTAIL.t2 B 0.032828f
C64 VTAIL.n35 B 0.119675f
C65 VTAIL.n36 B 0.011672f
C66 VTAIL.n37 B 0.014819f
C67 VTAIL.n38 B 0.019758f
C68 VTAIL.n39 B 0.008851f
C69 VTAIL.n40 B 0.008359f
C70 VTAIL.n41 B 0.015556f
C71 VTAIL.n42 B 0.015556f
C72 VTAIL.n43 B 0.008359f
C73 VTAIL.n44 B 0.008851f
C74 VTAIL.n45 B 0.019758f
C75 VTAIL.n46 B 0.019758f
C76 VTAIL.n47 B 0.008851f
C77 VTAIL.n48 B 0.008359f
C78 VTAIL.n49 B 0.015556f
C79 VTAIL.n50 B 0.015556f
C80 VTAIL.n51 B 0.008359f
C81 VTAIL.n52 B 0.008851f
C82 VTAIL.n53 B 0.019758f
C83 VTAIL.n54 B 0.019758f
C84 VTAIL.n55 B 0.008851f
C85 VTAIL.n56 B 0.008359f
C86 VTAIL.n57 B 0.015556f
C87 VTAIL.n58 B 0.015556f
C88 VTAIL.n59 B 0.008359f
C89 VTAIL.n60 B 0.008851f
C90 VTAIL.n61 B 0.019758f
C91 VTAIL.n62 B 0.019758f
C92 VTAIL.n63 B 0.008851f
C93 VTAIL.n64 B 0.008359f
C94 VTAIL.n65 B 0.015556f
C95 VTAIL.n66 B 0.015556f
C96 VTAIL.n67 B 0.008359f
C97 VTAIL.n68 B 0.008851f
C98 VTAIL.n69 B 0.019758f
C99 VTAIL.n70 B 0.019758f
C100 VTAIL.n71 B 0.008851f
C101 VTAIL.n72 B 0.008359f
C102 VTAIL.n73 B 0.015556f
C103 VTAIL.n74 B 0.015556f
C104 VTAIL.n75 B 0.008359f
C105 VTAIL.n76 B 0.008359f
C106 VTAIL.n77 B 0.008851f
C107 VTAIL.n78 B 0.019758f
C108 VTAIL.n79 B 0.019758f
C109 VTAIL.n80 B 0.019758f
C110 VTAIL.n81 B 0.008605f
C111 VTAIL.n82 B 0.008359f
C112 VTAIL.n83 B 0.015556f
C113 VTAIL.n84 B 0.015556f
C114 VTAIL.n85 B 0.008359f
C115 VTAIL.n86 B 0.008851f
C116 VTAIL.n87 B 0.019758f
C117 VTAIL.n88 B 0.019758f
C118 VTAIL.n89 B 0.008851f
C119 VTAIL.n90 B 0.008359f
C120 VTAIL.n91 B 0.015556f
C121 VTAIL.n92 B 0.015556f
C122 VTAIL.n93 B 0.008359f
C123 VTAIL.n94 B 0.008851f
C124 VTAIL.n95 B 0.019758f
C125 VTAIL.n96 B 0.019758f
C126 VTAIL.n97 B 0.008851f
C127 VTAIL.n98 B 0.008359f
C128 VTAIL.n99 B 0.015556f
C129 VTAIL.n100 B 0.015556f
C130 VTAIL.n101 B 0.008359f
C131 VTAIL.n102 B 0.008851f
C132 VTAIL.n103 B 0.019758f
C133 VTAIL.n104 B 0.044072f
C134 VTAIL.n105 B 0.008851f
C135 VTAIL.n106 B 0.008359f
C136 VTAIL.n107 B 0.035745f
C137 VTAIL.n108 B 0.024787f
C138 VTAIL.n109 B 0.128433f
C139 VTAIL.n110 B 0.0226f
C140 VTAIL.n111 B 0.015556f
C141 VTAIL.n112 B 0.008359f
C142 VTAIL.n113 B 0.019758f
C143 VTAIL.n114 B 0.008851f
C144 VTAIL.n115 B 0.015556f
C145 VTAIL.n116 B 0.008359f
C146 VTAIL.n117 B 0.019758f
C147 VTAIL.n118 B 0.008851f
C148 VTAIL.n119 B 0.015556f
C149 VTAIL.n120 B 0.008359f
C150 VTAIL.n121 B 0.019758f
C151 VTAIL.n122 B 0.008605f
C152 VTAIL.n123 B 0.015556f
C153 VTAIL.n124 B 0.008851f
C154 VTAIL.n125 B 0.019758f
C155 VTAIL.n126 B 0.008851f
C156 VTAIL.n127 B 0.015556f
C157 VTAIL.n128 B 0.008359f
C158 VTAIL.n129 B 0.019758f
C159 VTAIL.n130 B 0.008851f
C160 VTAIL.n131 B 0.015556f
C161 VTAIL.n132 B 0.008359f
C162 VTAIL.n133 B 0.019758f
C163 VTAIL.n134 B 0.008851f
C164 VTAIL.n135 B 0.015556f
C165 VTAIL.n136 B 0.008359f
C166 VTAIL.n137 B 0.019758f
C167 VTAIL.n138 B 0.008851f
C168 VTAIL.n139 B 0.015556f
C169 VTAIL.n140 B 0.008359f
C170 VTAIL.n141 B 0.019758f
C171 VTAIL.n142 B 0.008851f
C172 VTAIL.n143 B 1.34505f
C173 VTAIL.n144 B 0.008359f
C174 VTAIL.t5 B 0.032828f
C175 VTAIL.n145 B 0.119675f
C176 VTAIL.n146 B 0.011672f
C177 VTAIL.n147 B 0.014819f
C178 VTAIL.n148 B 0.019758f
C179 VTAIL.n149 B 0.008851f
C180 VTAIL.n150 B 0.008359f
C181 VTAIL.n151 B 0.015556f
C182 VTAIL.n152 B 0.015556f
C183 VTAIL.n153 B 0.008359f
C184 VTAIL.n154 B 0.008851f
C185 VTAIL.n155 B 0.019758f
C186 VTAIL.n156 B 0.019758f
C187 VTAIL.n157 B 0.008851f
C188 VTAIL.n158 B 0.008359f
C189 VTAIL.n159 B 0.015556f
C190 VTAIL.n160 B 0.015556f
C191 VTAIL.n161 B 0.008359f
C192 VTAIL.n162 B 0.008851f
C193 VTAIL.n163 B 0.019758f
C194 VTAIL.n164 B 0.019758f
C195 VTAIL.n165 B 0.008851f
C196 VTAIL.n166 B 0.008359f
C197 VTAIL.n167 B 0.015556f
C198 VTAIL.n168 B 0.015556f
C199 VTAIL.n169 B 0.008359f
C200 VTAIL.n170 B 0.008851f
C201 VTAIL.n171 B 0.019758f
C202 VTAIL.n172 B 0.019758f
C203 VTAIL.n173 B 0.008851f
C204 VTAIL.n174 B 0.008359f
C205 VTAIL.n175 B 0.015556f
C206 VTAIL.n176 B 0.015556f
C207 VTAIL.n177 B 0.008359f
C208 VTAIL.n178 B 0.008851f
C209 VTAIL.n179 B 0.019758f
C210 VTAIL.n180 B 0.019758f
C211 VTAIL.n181 B 0.008851f
C212 VTAIL.n182 B 0.008359f
C213 VTAIL.n183 B 0.015556f
C214 VTAIL.n184 B 0.015556f
C215 VTAIL.n185 B 0.008359f
C216 VTAIL.n186 B 0.008359f
C217 VTAIL.n187 B 0.008851f
C218 VTAIL.n188 B 0.019758f
C219 VTAIL.n189 B 0.019758f
C220 VTAIL.n190 B 0.019758f
C221 VTAIL.n191 B 0.008605f
C222 VTAIL.n192 B 0.008359f
C223 VTAIL.n193 B 0.015556f
C224 VTAIL.n194 B 0.015556f
C225 VTAIL.n195 B 0.008359f
C226 VTAIL.n196 B 0.008851f
C227 VTAIL.n197 B 0.019758f
C228 VTAIL.n198 B 0.019758f
C229 VTAIL.n199 B 0.008851f
C230 VTAIL.n200 B 0.008359f
C231 VTAIL.n201 B 0.015556f
C232 VTAIL.n202 B 0.015556f
C233 VTAIL.n203 B 0.008359f
C234 VTAIL.n204 B 0.008851f
C235 VTAIL.n205 B 0.019758f
C236 VTAIL.n206 B 0.019758f
C237 VTAIL.n207 B 0.008851f
C238 VTAIL.n208 B 0.008359f
C239 VTAIL.n209 B 0.015556f
C240 VTAIL.n210 B 0.015556f
C241 VTAIL.n211 B 0.008359f
C242 VTAIL.n212 B 0.008851f
C243 VTAIL.n213 B 0.019758f
C244 VTAIL.n214 B 0.044072f
C245 VTAIL.n215 B 0.008851f
C246 VTAIL.n216 B 0.008359f
C247 VTAIL.n217 B 0.035745f
C248 VTAIL.n218 B 0.024787f
C249 VTAIL.n219 B 0.214316f
C250 VTAIL.n220 B 0.0226f
C251 VTAIL.n221 B 0.015556f
C252 VTAIL.n222 B 0.008359f
C253 VTAIL.n223 B 0.019758f
C254 VTAIL.n224 B 0.008851f
C255 VTAIL.n225 B 0.015556f
C256 VTAIL.n226 B 0.008359f
C257 VTAIL.n227 B 0.019758f
C258 VTAIL.n228 B 0.008851f
C259 VTAIL.n229 B 0.015556f
C260 VTAIL.n230 B 0.008359f
C261 VTAIL.n231 B 0.019758f
C262 VTAIL.n232 B 0.008605f
C263 VTAIL.n233 B 0.015556f
C264 VTAIL.n234 B 0.008851f
C265 VTAIL.n235 B 0.019758f
C266 VTAIL.n236 B 0.008851f
C267 VTAIL.n237 B 0.015556f
C268 VTAIL.n238 B 0.008359f
C269 VTAIL.n239 B 0.019758f
C270 VTAIL.n240 B 0.008851f
C271 VTAIL.n241 B 0.015556f
C272 VTAIL.n242 B 0.008359f
C273 VTAIL.n243 B 0.019758f
C274 VTAIL.n244 B 0.008851f
C275 VTAIL.n245 B 0.015556f
C276 VTAIL.n246 B 0.008359f
C277 VTAIL.n247 B 0.019758f
C278 VTAIL.n248 B 0.008851f
C279 VTAIL.n249 B 0.015556f
C280 VTAIL.n250 B 0.008359f
C281 VTAIL.n251 B 0.019758f
C282 VTAIL.n252 B 0.008851f
C283 VTAIL.n253 B 1.34505f
C284 VTAIL.n254 B 0.008359f
C285 VTAIL.t7 B 0.032828f
C286 VTAIL.n255 B 0.119675f
C287 VTAIL.n256 B 0.011672f
C288 VTAIL.n257 B 0.014819f
C289 VTAIL.n258 B 0.019758f
C290 VTAIL.n259 B 0.008851f
C291 VTAIL.n260 B 0.008359f
C292 VTAIL.n261 B 0.015556f
C293 VTAIL.n262 B 0.015556f
C294 VTAIL.n263 B 0.008359f
C295 VTAIL.n264 B 0.008851f
C296 VTAIL.n265 B 0.019758f
C297 VTAIL.n266 B 0.019758f
C298 VTAIL.n267 B 0.008851f
C299 VTAIL.n268 B 0.008359f
C300 VTAIL.n269 B 0.015556f
C301 VTAIL.n270 B 0.015556f
C302 VTAIL.n271 B 0.008359f
C303 VTAIL.n272 B 0.008851f
C304 VTAIL.n273 B 0.019758f
C305 VTAIL.n274 B 0.019758f
C306 VTAIL.n275 B 0.008851f
C307 VTAIL.n276 B 0.008359f
C308 VTAIL.n277 B 0.015556f
C309 VTAIL.n278 B 0.015556f
C310 VTAIL.n279 B 0.008359f
C311 VTAIL.n280 B 0.008851f
C312 VTAIL.n281 B 0.019758f
C313 VTAIL.n282 B 0.019758f
C314 VTAIL.n283 B 0.008851f
C315 VTAIL.n284 B 0.008359f
C316 VTAIL.n285 B 0.015556f
C317 VTAIL.n286 B 0.015556f
C318 VTAIL.n287 B 0.008359f
C319 VTAIL.n288 B 0.008851f
C320 VTAIL.n289 B 0.019758f
C321 VTAIL.n290 B 0.019758f
C322 VTAIL.n291 B 0.008851f
C323 VTAIL.n292 B 0.008359f
C324 VTAIL.n293 B 0.015556f
C325 VTAIL.n294 B 0.015556f
C326 VTAIL.n295 B 0.008359f
C327 VTAIL.n296 B 0.008359f
C328 VTAIL.n297 B 0.008851f
C329 VTAIL.n298 B 0.019758f
C330 VTAIL.n299 B 0.019758f
C331 VTAIL.n300 B 0.019758f
C332 VTAIL.n301 B 0.008605f
C333 VTAIL.n302 B 0.008359f
C334 VTAIL.n303 B 0.015556f
C335 VTAIL.n304 B 0.015556f
C336 VTAIL.n305 B 0.008359f
C337 VTAIL.n306 B 0.008851f
C338 VTAIL.n307 B 0.019758f
C339 VTAIL.n308 B 0.019758f
C340 VTAIL.n309 B 0.008851f
C341 VTAIL.n310 B 0.008359f
C342 VTAIL.n311 B 0.015556f
C343 VTAIL.n312 B 0.015556f
C344 VTAIL.n313 B 0.008359f
C345 VTAIL.n314 B 0.008851f
C346 VTAIL.n315 B 0.019758f
C347 VTAIL.n316 B 0.019758f
C348 VTAIL.n317 B 0.008851f
C349 VTAIL.n318 B 0.008359f
C350 VTAIL.n319 B 0.015556f
C351 VTAIL.n320 B 0.015556f
C352 VTAIL.n321 B 0.008359f
C353 VTAIL.n322 B 0.008851f
C354 VTAIL.n323 B 0.019758f
C355 VTAIL.n324 B 0.044072f
C356 VTAIL.n325 B 0.008851f
C357 VTAIL.n326 B 0.008359f
C358 VTAIL.n327 B 0.035745f
C359 VTAIL.n328 B 0.024787f
C360 VTAIL.n329 B 1.42965f
C361 VTAIL.n330 B 0.0226f
C362 VTAIL.n331 B 0.015556f
C363 VTAIL.n332 B 0.008359f
C364 VTAIL.n333 B 0.019758f
C365 VTAIL.n334 B 0.008851f
C366 VTAIL.n335 B 0.015556f
C367 VTAIL.n336 B 0.008359f
C368 VTAIL.n337 B 0.019758f
C369 VTAIL.n338 B 0.008851f
C370 VTAIL.n339 B 0.015556f
C371 VTAIL.n340 B 0.008359f
C372 VTAIL.n341 B 0.019758f
C373 VTAIL.n342 B 0.008605f
C374 VTAIL.n343 B 0.015556f
C375 VTAIL.n344 B 0.008605f
C376 VTAIL.n345 B 0.008359f
C377 VTAIL.n346 B 0.019758f
C378 VTAIL.n347 B 0.019758f
C379 VTAIL.n348 B 0.008851f
C380 VTAIL.n349 B 0.015556f
C381 VTAIL.n350 B 0.008359f
C382 VTAIL.n351 B 0.019758f
C383 VTAIL.n352 B 0.008851f
C384 VTAIL.n353 B 0.015556f
C385 VTAIL.n354 B 0.008359f
C386 VTAIL.n355 B 0.019758f
C387 VTAIL.n356 B 0.008851f
C388 VTAIL.n357 B 0.015556f
C389 VTAIL.n358 B 0.008359f
C390 VTAIL.n359 B 0.019758f
C391 VTAIL.n360 B 0.008851f
C392 VTAIL.n361 B 0.015556f
C393 VTAIL.n362 B 0.008359f
C394 VTAIL.n363 B 0.019758f
C395 VTAIL.n364 B 0.008851f
C396 VTAIL.n365 B 1.34505f
C397 VTAIL.n366 B 0.008359f
C398 VTAIL.t1 B 0.032828f
C399 VTAIL.n367 B 0.119675f
C400 VTAIL.n368 B 0.011672f
C401 VTAIL.n369 B 0.014819f
C402 VTAIL.n370 B 0.019758f
C403 VTAIL.n371 B 0.008851f
C404 VTAIL.n372 B 0.008359f
C405 VTAIL.n373 B 0.015556f
C406 VTAIL.n374 B 0.015556f
C407 VTAIL.n375 B 0.008359f
C408 VTAIL.n376 B 0.008851f
C409 VTAIL.n377 B 0.019758f
C410 VTAIL.n378 B 0.019758f
C411 VTAIL.n379 B 0.008851f
C412 VTAIL.n380 B 0.008359f
C413 VTAIL.n381 B 0.015556f
C414 VTAIL.n382 B 0.015556f
C415 VTAIL.n383 B 0.008359f
C416 VTAIL.n384 B 0.008851f
C417 VTAIL.n385 B 0.019758f
C418 VTAIL.n386 B 0.019758f
C419 VTAIL.n387 B 0.008851f
C420 VTAIL.n388 B 0.008359f
C421 VTAIL.n389 B 0.015556f
C422 VTAIL.n390 B 0.015556f
C423 VTAIL.n391 B 0.008359f
C424 VTAIL.n392 B 0.008851f
C425 VTAIL.n393 B 0.019758f
C426 VTAIL.n394 B 0.019758f
C427 VTAIL.n395 B 0.008851f
C428 VTAIL.n396 B 0.008359f
C429 VTAIL.n397 B 0.015556f
C430 VTAIL.n398 B 0.015556f
C431 VTAIL.n399 B 0.008359f
C432 VTAIL.n400 B 0.008851f
C433 VTAIL.n401 B 0.019758f
C434 VTAIL.n402 B 0.019758f
C435 VTAIL.n403 B 0.008851f
C436 VTAIL.n404 B 0.008359f
C437 VTAIL.n405 B 0.015556f
C438 VTAIL.n406 B 0.015556f
C439 VTAIL.n407 B 0.008359f
C440 VTAIL.n408 B 0.008851f
C441 VTAIL.n409 B 0.019758f
C442 VTAIL.n410 B 0.019758f
C443 VTAIL.n411 B 0.008851f
C444 VTAIL.n412 B 0.008359f
C445 VTAIL.n413 B 0.015556f
C446 VTAIL.n414 B 0.015556f
C447 VTAIL.n415 B 0.008359f
C448 VTAIL.n416 B 0.008851f
C449 VTAIL.n417 B 0.019758f
C450 VTAIL.n418 B 0.019758f
C451 VTAIL.n419 B 0.008851f
C452 VTAIL.n420 B 0.008359f
C453 VTAIL.n421 B 0.015556f
C454 VTAIL.n422 B 0.015556f
C455 VTAIL.n423 B 0.008359f
C456 VTAIL.n424 B 0.008851f
C457 VTAIL.n425 B 0.019758f
C458 VTAIL.n426 B 0.019758f
C459 VTAIL.n427 B 0.008851f
C460 VTAIL.n428 B 0.008359f
C461 VTAIL.n429 B 0.015556f
C462 VTAIL.n430 B 0.015556f
C463 VTAIL.n431 B 0.008359f
C464 VTAIL.n432 B 0.008851f
C465 VTAIL.n433 B 0.019758f
C466 VTAIL.n434 B 0.044072f
C467 VTAIL.n435 B 0.008851f
C468 VTAIL.n436 B 0.008359f
C469 VTAIL.n437 B 0.035745f
C470 VTAIL.n438 B 0.024787f
C471 VTAIL.n439 B 1.42965f
C472 VTAIL.n440 B 0.0226f
C473 VTAIL.n441 B 0.015556f
C474 VTAIL.n442 B 0.008359f
C475 VTAIL.n443 B 0.019758f
C476 VTAIL.n444 B 0.008851f
C477 VTAIL.n445 B 0.015556f
C478 VTAIL.n446 B 0.008359f
C479 VTAIL.n447 B 0.019758f
C480 VTAIL.n448 B 0.008851f
C481 VTAIL.n449 B 0.015556f
C482 VTAIL.n450 B 0.008359f
C483 VTAIL.n451 B 0.019758f
C484 VTAIL.n452 B 0.008605f
C485 VTAIL.n453 B 0.015556f
C486 VTAIL.n454 B 0.008605f
C487 VTAIL.n455 B 0.008359f
C488 VTAIL.n456 B 0.019758f
C489 VTAIL.n457 B 0.019758f
C490 VTAIL.n458 B 0.008851f
C491 VTAIL.n459 B 0.015556f
C492 VTAIL.n460 B 0.008359f
C493 VTAIL.n461 B 0.019758f
C494 VTAIL.n462 B 0.008851f
C495 VTAIL.n463 B 0.015556f
C496 VTAIL.n464 B 0.008359f
C497 VTAIL.n465 B 0.019758f
C498 VTAIL.n466 B 0.008851f
C499 VTAIL.n467 B 0.015556f
C500 VTAIL.n468 B 0.008359f
C501 VTAIL.n469 B 0.019758f
C502 VTAIL.n470 B 0.008851f
C503 VTAIL.n471 B 0.015556f
C504 VTAIL.n472 B 0.008359f
C505 VTAIL.n473 B 0.019758f
C506 VTAIL.n474 B 0.008851f
C507 VTAIL.n475 B 1.34505f
C508 VTAIL.n476 B 0.008359f
C509 VTAIL.t3 B 0.032828f
C510 VTAIL.n477 B 0.119675f
C511 VTAIL.n478 B 0.011672f
C512 VTAIL.n479 B 0.014819f
C513 VTAIL.n480 B 0.019758f
C514 VTAIL.n481 B 0.008851f
C515 VTAIL.n482 B 0.008359f
C516 VTAIL.n483 B 0.015556f
C517 VTAIL.n484 B 0.015556f
C518 VTAIL.n485 B 0.008359f
C519 VTAIL.n486 B 0.008851f
C520 VTAIL.n487 B 0.019758f
C521 VTAIL.n488 B 0.019758f
C522 VTAIL.n489 B 0.008851f
C523 VTAIL.n490 B 0.008359f
C524 VTAIL.n491 B 0.015556f
C525 VTAIL.n492 B 0.015556f
C526 VTAIL.n493 B 0.008359f
C527 VTAIL.n494 B 0.008851f
C528 VTAIL.n495 B 0.019758f
C529 VTAIL.n496 B 0.019758f
C530 VTAIL.n497 B 0.008851f
C531 VTAIL.n498 B 0.008359f
C532 VTAIL.n499 B 0.015556f
C533 VTAIL.n500 B 0.015556f
C534 VTAIL.n501 B 0.008359f
C535 VTAIL.n502 B 0.008851f
C536 VTAIL.n503 B 0.019758f
C537 VTAIL.n504 B 0.019758f
C538 VTAIL.n505 B 0.008851f
C539 VTAIL.n506 B 0.008359f
C540 VTAIL.n507 B 0.015556f
C541 VTAIL.n508 B 0.015556f
C542 VTAIL.n509 B 0.008359f
C543 VTAIL.n510 B 0.008851f
C544 VTAIL.n511 B 0.019758f
C545 VTAIL.n512 B 0.019758f
C546 VTAIL.n513 B 0.008851f
C547 VTAIL.n514 B 0.008359f
C548 VTAIL.n515 B 0.015556f
C549 VTAIL.n516 B 0.015556f
C550 VTAIL.n517 B 0.008359f
C551 VTAIL.n518 B 0.008851f
C552 VTAIL.n519 B 0.019758f
C553 VTAIL.n520 B 0.019758f
C554 VTAIL.n521 B 0.008851f
C555 VTAIL.n522 B 0.008359f
C556 VTAIL.n523 B 0.015556f
C557 VTAIL.n524 B 0.015556f
C558 VTAIL.n525 B 0.008359f
C559 VTAIL.n526 B 0.008851f
C560 VTAIL.n527 B 0.019758f
C561 VTAIL.n528 B 0.019758f
C562 VTAIL.n529 B 0.008851f
C563 VTAIL.n530 B 0.008359f
C564 VTAIL.n531 B 0.015556f
C565 VTAIL.n532 B 0.015556f
C566 VTAIL.n533 B 0.008359f
C567 VTAIL.n534 B 0.008851f
C568 VTAIL.n535 B 0.019758f
C569 VTAIL.n536 B 0.019758f
C570 VTAIL.n537 B 0.008851f
C571 VTAIL.n538 B 0.008359f
C572 VTAIL.n539 B 0.015556f
C573 VTAIL.n540 B 0.015556f
C574 VTAIL.n541 B 0.008359f
C575 VTAIL.n542 B 0.008851f
C576 VTAIL.n543 B 0.019758f
C577 VTAIL.n544 B 0.044072f
C578 VTAIL.n545 B 0.008851f
C579 VTAIL.n546 B 0.008359f
C580 VTAIL.n547 B 0.035745f
C581 VTAIL.n548 B 0.024787f
C582 VTAIL.n549 B 0.214316f
C583 VTAIL.n550 B 0.0226f
C584 VTAIL.n551 B 0.015556f
C585 VTAIL.n552 B 0.008359f
C586 VTAIL.n553 B 0.019758f
C587 VTAIL.n554 B 0.008851f
C588 VTAIL.n555 B 0.015556f
C589 VTAIL.n556 B 0.008359f
C590 VTAIL.n557 B 0.019758f
C591 VTAIL.n558 B 0.008851f
C592 VTAIL.n559 B 0.015556f
C593 VTAIL.n560 B 0.008359f
C594 VTAIL.n561 B 0.019758f
C595 VTAIL.n562 B 0.008605f
C596 VTAIL.n563 B 0.015556f
C597 VTAIL.n564 B 0.008605f
C598 VTAIL.n565 B 0.008359f
C599 VTAIL.n566 B 0.019758f
C600 VTAIL.n567 B 0.019758f
C601 VTAIL.n568 B 0.008851f
C602 VTAIL.n569 B 0.015556f
C603 VTAIL.n570 B 0.008359f
C604 VTAIL.n571 B 0.019758f
C605 VTAIL.n572 B 0.008851f
C606 VTAIL.n573 B 0.015556f
C607 VTAIL.n574 B 0.008359f
C608 VTAIL.n575 B 0.019758f
C609 VTAIL.n576 B 0.008851f
C610 VTAIL.n577 B 0.015556f
C611 VTAIL.n578 B 0.008359f
C612 VTAIL.n579 B 0.019758f
C613 VTAIL.n580 B 0.008851f
C614 VTAIL.n581 B 0.015556f
C615 VTAIL.n582 B 0.008359f
C616 VTAIL.n583 B 0.019758f
C617 VTAIL.n584 B 0.008851f
C618 VTAIL.n585 B 1.34505f
C619 VTAIL.n586 B 0.008359f
C620 VTAIL.t6 B 0.032828f
C621 VTAIL.n587 B 0.119675f
C622 VTAIL.n588 B 0.011672f
C623 VTAIL.n589 B 0.014819f
C624 VTAIL.n590 B 0.019758f
C625 VTAIL.n591 B 0.008851f
C626 VTAIL.n592 B 0.008359f
C627 VTAIL.n593 B 0.015556f
C628 VTAIL.n594 B 0.015556f
C629 VTAIL.n595 B 0.008359f
C630 VTAIL.n596 B 0.008851f
C631 VTAIL.n597 B 0.019758f
C632 VTAIL.n598 B 0.019758f
C633 VTAIL.n599 B 0.008851f
C634 VTAIL.n600 B 0.008359f
C635 VTAIL.n601 B 0.015556f
C636 VTAIL.n602 B 0.015556f
C637 VTAIL.n603 B 0.008359f
C638 VTAIL.n604 B 0.008851f
C639 VTAIL.n605 B 0.019758f
C640 VTAIL.n606 B 0.019758f
C641 VTAIL.n607 B 0.008851f
C642 VTAIL.n608 B 0.008359f
C643 VTAIL.n609 B 0.015556f
C644 VTAIL.n610 B 0.015556f
C645 VTAIL.n611 B 0.008359f
C646 VTAIL.n612 B 0.008851f
C647 VTAIL.n613 B 0.019758f
C648 VTAIL.n614 B 0.019758f
C649 VTAIL.n615 B 0.008851f
C650 VTAIL.n616 B 0.008359f
C651 VTAIL.n617 B 0.015556f
C652 VTAIL.n618 B 0.015556f
C653 VTAIL.n619 B 0.008359f
C654 VTAIL.n620 B 0.008851f
C655 VTAIL.n621 B 0.019758f
C656 VTAIL.n622 B 0.019758f
C657 VTAIL.n623 B 0.008851f
C658 VTAIL.n624 B 0.008359f
C659 VTAIL.n625 B 0.015556f
C660 VTAIL.n626 B 0.015556f
C661 VTAIL.n627 B 0.008359f
C662 VTAIL.n628 B 0.008851f
C663 VTAIL.n629 B 0.019758f
C664 VTAIL.n630 B 0.019758f
C665 VTAIL.n631 B 0.008851f
C666 VTAIL.n632 B 0.008359f
C667 VTAIL.n633 B 0.015556f
C668 VTAIL.n634 B 0.015556f
C669 VTAIL.n635 B 0.008359f
C670 VTAIL.n636 B 0.008851f
C671 VTAIL.n637 B 0.019758f
C672 VTAIL.n638 B 0.019758f
C673 VTAIL.n639 B 0.008851f
C674 VTAIL.n640 B 0.008359f
C675 VTAIL.n641 B 0.015556f
C676 VTAIL.n642 B 0.015556f
C677 VTAIL.n643 B 0.008359f
C678 VTAIL.n644 B 0.008851f
C679 VTAIL.n645 B 0.019758f
C680 VTAIL.n646 B 0.019758f
C681 VTAIL.n647 B 0.008851f
C682 VTAIL.n648 B 0.008359f
C683 VTAIL.n649 B 0.015556f
C684 VTAIL.n650 B 0.015556f
C685 VTAIL.n651 B 0.008359f
C686 VTAIL.n652 B 0.008851f
C687 VTAIL.n653 B 0.019758f
C688 VTAIL.n654 B 0.044072f
C689 VTAIL.n655 B 0.008851f
C690 VTAIL.n656 B 0.008359f
C691 VTAIL.n657 B 0.035745f
C692 VTAIL.n658 B 0.024787f
C693 VTAIL.n659 B 0.214316f
C694 VTAIL.n660 B 0.0226f
C695 VTAIL.n661 B 0.015556f
C696 VTAIL.n662 B 0.008359f
C697 VTAIL.n663 B 0.019758f
C698 VTAIL.n664 B 0.008851f
C699 VTAIL.n665 B 0.015556f
C700 VTAIL.n666 B 0.008359f
C701 VTAIL.n667 B 0.019758f
C702 VTAIL.n668 B 0.008851f
C703 VTAIL.n669 B 0.015556f
C704 VTAIL.n670 B 0.008359f
C705 VTAIL.n671 B 0.019758f
C706 VTAIL.n672 B 0.008605f
C707 VTAIL.n673 B 0.015556f
C708 VTAIL.n674 B 0.008605f
C709 VTAIL.n675 B 0.008359f
C710 VTAIL.n676 B 0.019758f
C711 VTAIL.n677 B 0.019758f
C712 VTAIL.n678 B 0.008851f
C713 VTAIL.n679 B 0.015556f
C714 VTAIL.n680 B 0.008359f
C715 VTAIL.n681 B 0.019758f
C716 VTAIL.n682 B 0.008851f
C717 VTAIL.n683 B 0.015556f
C718 VTAIL.n684 B 0.008359f
C719 VTAIL.n685 B 0.019758f
C720 VTAIL.n686 B 0.008851f
C721 VTAIL.n687 B 0.015556f
C722 VTAIL.n688 B 0.008359f
C723 VTAIL.n689 B 0.019758f
C724 VTAIL.n690 B 0.008851f
C725 VTAIL.n691 B 0.015556f
C726 VTAIL.n692 B 0.008359f
C727 VTAIL.n693 B 0.019758f
C728 VTAIL.n694 B 0.008851f
C729 VTAIL.n695 B 1.34505f
C730 VTAIL.n696 B 0.008359f
C731 VTAIL.t4 B 0.032828f
C732 VTAIL.n697 B 0.119675f
C733 VTAIL.n698 B 0.011672f
C734 VTAIL.n699 B 0.014819f
C735 VTAIL.n700 B 0.019758f
C736 VTAIL.n701 B 0.008851f
C737 VTAIL.n702 B 0.008359f
C738 VTAIL.n703 B 0.015556f
C739 VTAIL.n704 B 0.015556f
C740 VTAIL.n705 B 0.008359f
C741 VTAIL.n706 B 0.008851f
C742 VTAIL.n707 B 0.019758f
C743 VTAIL.n708 B 0.019758f
C744 VTAIL.n709 B 0.008851f
C745 VTAIL.n710 B 0.008359f
C746 VTAIL.n711 B 0.015556f
C747 VTAIL.n712 B 0.015556f
C748 VTAIL.n713 B 0.008359f
C749 VTAIL.n714 B 0.008851f
C750 VTAIL.n715 B 0.019758f
C751 VTAIL.n716 B 0.019758f
C752 VTAIL.n717 B 0.008851f
C753 VTAIL.n718 B 0.008359f
C754 VTAIL.n719 B 0.015556f
C755 VTAIL.n720 B 0.015556f
C756 VTAIL.n721 B 0.008359f
C757 VTAIL.n722 B 0.008851f
C758 VTAIL.n723 B 0.019758f
C759 VTAIL.n724 B 0.019758f
C760 VTAIL.n725 B 0.008851f
C761 VTAIL.n726 B 0.008359f
C762 VTAIL.n727 B 0.015556f
C763 VTAIL.n728 B 0.015556f
C764 VTAIL.n729 B 0.008359f
C765 VTAIL.n730 B 0.008851f
C766 VTAIL.n731 B 0.019758f
C767 VTAIL.n732 B 0.019758f
C768 VTAIL.n733 B 0.008851f
C769 VTAIL.n734 B 0.008359f
C770 VTAIL.n735 B 0.015556f
C771 VTAIL.n736 B 0.015556f
C772 VTAIL.n737 B 0.008359f
C773 VTAIL.n738 B 0.008851f
C774 VTAIL.n739 B 0.019758f
C775 VTAIL.n740 B 0.019758f
C776 VTAIL.n741 B 0.008851f
C777 VTAIL.n742 B 0.008359f
C778 VTAIL.n743 B 0.015556f
C779 VTAIL.n744 B 0.015556f
C780 VTAIL.n745 B 0.008359f
C781 VTAIL.n746 B 0.008851f
C782 VTAIL.n747 B 0.019758f
C783 VTAIL.n748 B 0.019758f
C784 VTAIL.n749 B 0.008851f
C785 VTAIL.n750 B 0.008359f
C786 VTAIL.n751 B 0.015556f
C787 VTAIL.n752 B 0.015556f
C788 VTAIL.n753 B 0.008359f
C789 VTAIL.n754 B 0.008851f
C790 VTAIL.n755 B 0.019758f
C791 VTAIL.n756 B 0.019758f
C792 VTAIL.n757 B 0.008851f
C793 VTAIL.n758 B 0.008359f
C794 VTAIL.n759 B 0.015556f
C795 VTAIL.n760 B 0.015556f
C796 VTAIL.n761 B 0.008359f
C797 VTAIL.n762 B 0.008851f
C798 VTAIL.n763 B 0.019758f
C799 VTAIL.n764 B 0.044072f
C800 VTAIL.n765 B 0.008851f
C801 VTAIL.n766 B 0.008359f
C802 VTAIL.n767 B 0.035745f
C803 VTAIL.n768 B 0.024787f
C804 VTAIL.n769 B 1.42965f
C805 VTAIL.n770 B 0.0226f
C806 VTAIL.n771 B 0.015556f
C807 VTAIL.n772 B 0.008359f
C808 VTAIL.n773 B 0.019758f
C809 VTAIL.n774 B 0.008851f
C810 VTAIL.n775 B 0.015556f
C811 VTAIL.n776 B 0.008359f
C812 VTAIL.n777 B 0.019758f
C813 VTAIL.n778 B 0.008851f
C814 VTAIL.n779 B 0.015556f
C815 VTAIL.n780 B 0.008359f
C816 VTAIL.n781 B 0.019758f
C817 VTAIL.n782 B 0.008605f
C818 VTAIL.n783 B 0.015556f
C819 VTAIL.n784 B 0.008851f
C820 VTAIL.n785 B 0.019758f
C821 VTAIL.n786 B 0.008851f
C822 VTAIL.n787 B 0.015556f
C823 VTAIL.n788 B 0.008359f
C824 VTAIL.n789 B 0.019758f
C825 VTAIL.n790 B 0.008851f
C826 VTAIL.n791 B 0.015556f
C827 VTAIL.n792 B 0.008359f
C828 VTAIL.n793 B 0.019758f
C829 VTAIL.n794 B 0.008851f
C830 VTAIL.n795 B 0.015556f
C831 VTAIL.n796 B 0.008359f
C832 VTAIL.n797 B 0.019758f
C833 VTAIL.n798 B 0.008851f
C834 VTAIL.n799 B 0.015556f
C835 VTAIL.n800 B 0.008359f
C836 VTAIL.n801 B 0.019758f
C837 VTAIL.n802 B 0.008851f
C838 VTAIL.n803 B 1.34505f
C839 VTAIL.n804 B 0.008359f
C840 VTAIL.t0 B 0.032828f
C841 VTAIL.n805 B 0.119675f
C842 VTAIL.n806 B 0.011672f
C843 VTAIL.n807 B 0.014819f
C844 VTAIL.n808 B 0.019758f
C845 VTAIL.n809 B 0.008851f
C846 VTAIL.n810 B 0.008359f
C847 VTAIL.n811 B 0.015556f
C848 VTAIL.n812 B 0.015556f
C849 VTAIL.n813 B 0.008359f
C850 VTAIL.n814 B 0.008851f
C851 VTAIL.n815 B 0.019758f
C852 VTAIL.n816 B 0.019758f
C853 VTAIL.n817 B 0.008851f
C854 VTAIL.n818 B 0.008359f
C855 VTAIL.n819 B 0.015556f
C856 VTAIL.n820 B 0.015556f
C857 VTAIL.n821 B 0.008359f
C858 VTAIL.n822 B 0.008851f
C859 VTAIL.n823 B 0.019758f
C860 VTAIL.n824 B 0.019758f
C861 VTAIL.n825 B 0.008851f
C862 VTAIL.n826 B 0.008359f
C863 VTAIL.n827 B 0.015556f
C864 VTAIL.n828 B 0.015556f
C865 VTAIL.n829 B 0.008359f
C866 VTAIL.n830 B 0.008851f
C867 VTAIL.n831 B 0.019758f
C868 VTAIL.n832 B 0.019758f
C869 VTAIL.n833 B 0.008851f
C870 VTAIL.n834 B 0.008359f
C871 VTAIL.n835 B 0.015556f
C872 VTAIL.n836 B 0.015556f
C873 VTAIL.n837 B 0.008359f
C874 VTAIL.n838 B 0.008851f
C875 VTAIL.n839 B 0.019758f
C876 VTAIL.n840 B 0.019758f
C877 VTAIL.n841 B 0.008851f
C878 VTAIL.n842 B 0.008359f
C879 VTAIL.n843 B 0.015556f
C880 VTAIL.n844 B 0.015556f
C881 VTAIL.n845 B 0.008359f
C882 VTAIL.n846 B 0.008359f
C883 VTAIL.n847 B 0.008851f
C884 VTAIL.n848 B 0.019758f
C885 VTAIL.n849 B 0.019758f
C886 VTAIL.n850 B 0.019758f
C887 VTAIL.n851 B 0.008605f
C888 VTAIL.n852 B 0.008359f
C889 VTAIL.n853 B 0.015556f
C890 VTAIL.n854 B 0.015556f
C891 VTAIL.n855 B 0.008359f
C892 VTAIL.n856 B 0.008851f
C893 VTAIL.n857 B 0.019758f
C894 VTAIL.n858 B 0.019758f
C895 VTAIL.n859 B 0.008851f
C896 VTAIL.n860 B 0.008359f
C897 VTAIL.n861 B 0.015556f
C898 VTAIL.n862 B 0.015556f
C899 VTAIL.n863 B 0.008359f
C900 VTAIL.n864 B 0.008851f
C901 VTAIL.n865 B 0.019758f
C902 VTAIL.n866 B 0.019758f
C903 VTAIL.n867 B 0.008851f
C904 VTAIL.n868 B 0.008359f
C905 VTAIL.n869 B 0.015556f
C906 VTAIL.n870 B 0.015556f
C907 VTAIL.n871 B 0.008359f
C908 VTAIL.n872 B 0.008851f
C909 VTAIL.n873 B 0.019758f
C910 VTAIL.n874 B 0.044072f
C911 VTAIL.n875 B 0.008851f
C912 VTAIL.n876 B 0.008359f
C913 VTAIL.n877 B 0.035745f
C914 VTAIL.n878 B 0.024787f
C915 VTAIL.n879 B 1.33793f
C916 VDD1.t3 B 0.418748f
C917 VDD1.t0 B 0.418748f
C918 VDD1.n0 B 3.82738f
C919 VDD1.t2 B 0.418748f
C920 VDD1.t1 B 0.418748f
C921 VDD1.n1 B 4.90915f
C922 VP.t2 B 3.86059f
C923 VP.n0 B 1.39658f
C924 VP.n1 B 0.018847f
C925 VP.n2 B 0.037458f
C926 VP.n3 B 0.018847f
C927 VP.n4 B 0.035126f
C928 VP.t1 B 4.17525f
C929 VP.t3 B 4.16325f
C930 VP.n5 B 3.96396f
C931 VP.n6 B 1.32411f
C932 VP.t0 B 3.86059f
C933 VP.n7 B 1.39658f
C934 VP.n8 B 0.019691f
C935 VP.n9 B 0.030419f
C936 VP.n10 B 0.018847f
C937 VP.n11 B 0.018847f
C938 VP.n12 B 0.035126f
C939 VP.n13 B 0.037458f
C940 VP.n14 B 0.015236f
C941 VP.n15 B 0.018847f
C942 VP.n16 B 0.018847f
C943 VP.n17 B 0.018847f
C944 VP.n18 B 0.035126f
C945 VP.n19 B 0.035126f
C946 VP.n20 B 0.019691f
C947 VP.n21 B 0.030419f
C948 VP.n22 B 0.057795f
.ends

