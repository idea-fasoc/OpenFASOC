* NGSPICE file created from diff_pair_sample_1524.ext - technology: sky130A

.subckt diff_pair_sample_1524 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X1 VTAIL.t18 VP.t1 VDD1.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X2 VTAIL.t19 VN.t0 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X3 VDD2.t8 VN.t1 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X4 VDD1.t7 VP.t2 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.29
X5 VDD1.t6 VP.t3 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.29
X6 VDD2.t7 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X7 VTAIL.t10 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X8 VTAIL.t6 VN.t3 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X9 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.29
X10 VTAIL.t5 VN.t4 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X11 VDD1.t4 VP.t5 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.29
X12 VDD1.t3 VP.t6 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X13 VTAIL.t9 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X14 VDD1.t1 VP.t8 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.29
X15 VDD2.t4 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.29
X16 VDD2.t3 VN.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.29
X17 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.29
X18 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.29
X19 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.29
X20 VTAIL.t13 VP.t9 VDD1.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X21 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.29
X22 VTAIL.t0 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.29
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.29
R0 VP.n19 VP.t8 233.322
R1 VP.n5 VP.t6 201.745
R2 VP.n49 VP.t5 201.745
R3 VP.n57 VP.t9 201.745
R4 VP.n75 VP.t1 201.745
R5 VP.n83 VP.t3 201.745
R6 VP.n16 VP.t0 201.745
R7 VP.n46 VP.t2 201.745
R8 VP.n38 VP.t7 201.745
R9 VP.n20 VP.t4 201.745
R10 VP.n22 VP.n21 161.3
R11 VP.n23 VP.n18 161.3
R12 VP.n25 VP.n24 161.3
R13 VP.n26 VP.n17 161.3
R14 VP.n28 VP.n27 161.3
R15 VP.n29 VP.n16 161.3
R16 VP.n31 VP.n30 161.3
R17 VP.n32 VP.n15 161.3
R18 VP.n34 VP.n33 161.3
R19 VP.n35 VP.n14 161.3
R20 VP.n37 VP.n36 161.3
R21 VP.n39 VP.n13 161.3
R22 VP.n41 VP.n40 161.3
R23 VP.n42 VP.n12 161.3
R24 VP.n44 VP.n43 161.3
R25 VP.n45 VP.n11 161.3
R26 VP.n82 VP.n0 161.3
R27 VP.n81 VP.n80 161.3
R28 VP.n79 VP.n1 161.3
R29 VP.n78 VP.n77 161.3
R30 VP.n76 VP.n2 161.3
R31 VP.n74 VP.n73 161.3
R32 VP.n72 VP.n3 161.3
R33 VP.n71 VP.n70 161.3
R34 VP.n69 VP.n4 161.3
R35 VP.n68 VP.n67 161.3
R36 VP.n66 VP.n5 161.3
R37 VP.n65 VP.n64 161.3
R38 VP.n63 VP.n6 161.3
R39 VP.n62 VP.n61 161.3
R40 VP.n60 VP.n7 161.3
R41 VP.n59 VP.n58 161.3
R42 VP.n56 VP.n8 161.3
R43 VP.n55 VP.n54 161.3
R44 VP.n53 VP.n9 161.3
R45 VP.n52 VP.n51 161.3
R46 VP.n50 VP.n10 161.3
R47 VP.n49 VP.n48 99.0123
R48 VP.n84 VP.n83 99.0123
R49 VP.n47 VP.n46 99.0123
R50 VP.n20 VP.n19 66.166
R51 VP.n48 VP.n47 56.8329
R52 VP.n63 VP.n62 56.5193
R53 VP.n70 VP.n69 56.5193
R54 VP.n33 VP.n32 56.5193
R55 VP.n26 VP.n25 56.5193
R56 VP.n55 VP.n9 47.2923
R57 VP.n77 VP.n1 47.2923
R58 VP.n40 VP.n12 47.2923
R59 VP.n51 VP.n9 33.6945
R60 VP.n81 VP.n1 33.6945
R61 VP.n44 VP.n12 33.6945
R62 VP.n51 VP.n50 24.4675
R63 VP.n56 VP.n55 24.4675
R64 VP.n58 VP.n7 24.4675
R65 VP.n62 VP.n7 24.4675
R66 VP.n64 VP.n63 24.4675
R67 VP.n64 VP.n5 24.4675
R68 VP.n68 VP.n5 24.4675
R69 VP.n69 VP.n68 24.4675
R70 VP.n70 VP.n3 24.4675
R71 VP.n74 VP.n3 24.4675
R72 VP.n77 VP.n76 24.4675
R73 VP.n82 VP.n81 24.4675
R74 VP.n45 VP.n44 24.4675
R75 VP.n33 VP.n14 24.4675
R76 VP.n37 VP.n14 24.4675
R77 VP.n40 VP.n39 24.4675
R78 VP.n27 VP.n26 24.4675
R79 VP.n27 VP.n16 24.4675
R80 VP.n31 VP.n16 24.4675
R81 VP.n32 VP.n31 24.4675
R82 VP.n21 VP.n18 24.4675
R83 VP.n25 VP.n18 24.4675
R84 VP.n57 VP.n56 18.5954
R85 VP.n76 VP.n75 18.5954
R86 VP.n39 VP.n38 18.5954
R87 VP.n50 VP.n49 11.7447
R88 VP.n83 VP.n82 11.7447
R89 VP.n46 VP.n45 11.7447
R90 VP.n22 VP.n19 9.81663
R91 VP.n58 VP.n57 5.87258
R92 VP.n75 VP.n74 5.87258
R93 VP.n38 VP.n37 5.87258
R94 VP.n21 VP.n20 5.87258
R95 VP.n47 VP.n11 0.278367
R96 VP.n48 VP.n10 0.278367
R97 VP.n84 VP.n0 0.278367
R98 VP.n23 VP.n22 0.189894
R99 VP.n24 VP.n23 0.189894
R100 VP.n24 VP.n17 0.189894
R101 VP.n28 VP.n17 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n30 VP.n29 0.189894
R104 VP.n30 VP.n15 0.189894
R105 VP.n34 VP.n15 0.189894
R106 VP.n35 VP.n34 0.189894
R107 VP.n36 VP.n35 0.189894
R108 VP.n36 VP.n13 0.189894
R109 VP.n41 VP.n13 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n43 VP.n42 0.189894
R112 VP.n43 VP.n11 0.189894
R113 VP.n52 VP.n10 0.189894
R114 VP.n53 VP.n52 0.189894
R115 VP.n54 VP.n53 0.189894
R116 VP.n54 VP.n8 0.189894
R117 VP.n59 VP.n8 0.189894
R118 VP.n60 VP.n59 0.189894
R119 VP.n61 VP.n60 0.189894
R120 VP.n61 VP.n6 0.189894
R121 VP.n65 VP.n6 0.189894
R122 VP.n66 VP.n65 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n67 VP.n4 0.189894
R125 VP.n71 VP.n4 0.189894
R126 VP.n72 VP.n71 0.189894
R127 VP.n73 VP.n72 0.189894
R128 VP.n73 VP.n2 0.189894
R129 VP.n78 VP.n2 0.189894
R130 VP.n79 VP.n78 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n80 VP.n0 0.189894
R133 VP VP.n84 0.153454
R134 VTAIL.n11 VTAIL.t1 48.6263
R135 VTAIL.n17 VTAIL.t2 48.6262
R136 VTAIL.n2 VTAIL.t15 48.6262
R137 VTAIL.n16 VTAIL.t17 48.6262
R138 VTAIL.n15 VTAIL.n14 47.5935
R139 VTAIL.n13 VTAIL.n12 47.5935
R140 VTAIL.n10 VTAIL.n9 47.5935
R141 VTAIL.n8 VTAIL.n7 47.5935
R142 VTAIL.n19 VTAIL.n18 47.5923
R143 VTAIL.n1 VTAIL.n0 47.5923
R144 VTAIL.n4 VTAIL.n3 47.5923
R145 VTAIL.n6 VTAIL.n5 47.5923
R146 VTAIL.n8 VTAIL.n6 33.41
R147 VTAIL.n17 VTAIL.n16 31.1514
R148 VTAIL.n10 VTAIL.n8 2.25912
R149 VTAIL.n11 VTAIL.n10 2.25912
R150 VTAIL.n15 VTAIL.n13 2.25912
R151 VTAIL.n16 VTAIL.n15 2.25912
R152 VTAIL.n6 VTAIL.n4 2.25912
R153 VTAIL.n4 VTAIL.n2 2.25912
R154 VTAIL.n19 VTAIL.n17 2.25912
R155 VTAIL VTAIL.n1 1.75266
R156 VTAIL.n13 VTAIL.n11 1.59964
R157 VTAIL.n2 VTAIL.n1 1.59964
R158 VTAIL.n18 VTAIL.t7 1.03336
R159 VTAIL.n18 VTAIL.t0 1.03336
R160 VTAIL.n0 VTAIL.t4 1.03336
R161 VTAIL.n0 VTAIL.t5 1.03336
R162 VTAIL.n3 VTAIL.t14 1.03336
R163 VTAIL.n3 VTAIL.t18 1.03336
R164 VTAIL.n5 VTAIL.t12 1.03336
R165 VTAIL.n5 VTAIL.t13 1.03336
R166 VTAIL.n14 VTAIL.t11 1.03336
R167 VTAIL.n14 VTAIL.t9 1.03336
R168 VTAIL.n12 VTAIL.t16 1.03336
R169 VTAIL.n12 VTAIL.t10 1.03336
R170 VTAIL.n9 VTAIL.t8 1.03336
R171 VTAIL.n9 VTAIL.t6 1.03336
R172 VTAIL.n7 VTAIL.t3 1.03336
R173 VTAIL.n7 VTAIL.t19 1.03336
R174 VTAIL VTAIL.n19 0.506965
R175 VDD1.n1 VDD1.t1 67.5637
R176 VDD1.n3 VDD1.t4 67.5636
R177 VDD1.n5 VDD1.n4 65.9097
R178 VDD1.n1 VDD1.n0 64.2723
R179 VDD1.n7 VDD1.n6 64.2721
R180 VDD1.n3 VDD1.n2 64.2711
R181 VDD1.n7 VDD1.n5 52.6819
R182 VDD1 VDD1.n7 1.63628
R183 VDD1.n6 VDD1.t2 1.03336
R184 VDD1.n6 VDD1.t7 1.03336
R185 VDD1.n0 VDD1.t5 1.03336
R186 VDD1.n0 VDD1.t9 1.03336
R187 VDD1.n4 VDD1.t8 1.03336
R188 VDD1.n4 VDD1.t6 1.03336
R189 VDD1.n2 VDD1.t0 1.03336
R190 VDD1.n2 VDD1.t3 1.03336
R191 VDD1 VDD1.n1 0.623345
R192 VDD1.n5 VDD1.n3 0.509809
R193 B.n855 B.n854 585
R194 B.n855 B.n100 585
R195 B.n858 B.n857 585
R196 B.n859 B.n172 585
R197 B.n861 B.n860 585
R198 B.n863 B.n171 585
R199 B.n866 B.n865 585
R200 B.n867 B.n170 585
R201 B.n869 B.n868 585
R202 B.n871 B.n169 585
R203 B.n874 B.n873 585
R204 B.n875 B.n168 585
R205 B.n877 B.n876 585
R206 B.n879 B.n167 585
R207 B.n882 B.n881 585
R208 B.n883 B.n166 585
R209 B.n885 B.n884 585
R210 B.n887 B.n165 585
R211 B.n890 B.n889 585
R212 B.n891 B.n164 585
R213 B.n893 B.n892 585
R214 B.n895 B.n163 585
R215 B.n898 B.n897 585
R216 B.n899 B.n162 585
R217 B.n901 B.n900 585
R218 B.n903 B.n161 585
R219 B.n906 B.n905 585
R220 B.n907 B.n160 585
R221 B.n909 B.n908 585
R222 B.n911 B.n159 585
R223 B.n914 B.n913 585
R224 B.n915 B.n158 585
R225 B.n917 B.n916 585
R226 B.n919 B.n157 585
R227 B.n922 B.n921 585
R228 B.n923 B.n156 585
R229 B.n925 B.n924 585
R230 B.n927 B.n155 585
R231 B.n930 B.n929 585
R232 B.n931 B.n154 585
R233 B.n933 B.n932 585
R234 B.n935 B.n153 585
R235 B.n938 B.n937 585
R236 B.n939 B.n152 585
R237 B.n941 B.n940 585
R238 B.n943 B.n151 585
R239 B.n946 B.n945 585
R240 B.n947 B.n150 585
R241 B.n949 B.n948 585
R242 B.n951 B.n149 585
R243 B.n954 B.n953 585
R244 B.n955 B.n148 585
R245 B.n957 B.n956 585
R246 B.n959 B.n147 585
R247 B.n962 B.n961 585
R248 B.n963 B.n146 585
R249 B.n965 B.n964 585
R250 B.n967 B.n145 585
R251 B.n970 B.n969 585
R252 B.n971 B.n144 585
R253 B.n973 B.n972 585
R254 B.n975 B.n143 585
R255 B.n978 B.n977 585
R256 B.n979 B.n140 585
R257 B.n982 B.n981 585
R258 B.n984 B.n139 585
R259 B.n987 B.n986 585
R260 B.n988 B.n138 585
R261 B.n990 B.n989 585
R262 B.n992 B.n137 585
R263 B.n995 B.n994 585
R264 B.n996 B.n133 585
R265 B.n998 B.n997 585
R266 B.n1000 B.n132 585
R267 B.n1003 B.n1002 585
R268 B.n1004 B.n131 585
R269 B.n1006 B.n1005 585
R270 B.n1008 B.n130 585
R271 B.n1011 B.n1010 585
R272 B.n1012 B.n129 585
R273 B.n1014 B.n1013 585
R274 B.n1016 B.n128 585
R275 B.n1019 B.n1018 585
R276 B.n1020 B.n127 585
R277 B.n1022 B.n1021 585
R278 B.n1024 B.n126 585
R279 B.n1027 B.n1026 585
R280 B.n1028 B.n125 585
R281 B.n1030 B.n1029 585
R282 B.n1032 B.n124 585
R283 B.n1035 B.n1034 585
R284 B.n1036 B.n123 585
R285 B.n1038 B.n1037 585
R286 B.n1040 B.n122 585
R287 B.n1043 B.n1042 585
R288 B.n1044 B.n121 585
R289 B.n1046 B.n1045 585
R290 B.n1048 B.n120 585
R291 B.n1051 B.n1050 585
R292 B.n1052 B.n119 585
R293 B.n1054 B.n1053 585
R294 B.n1056 B.n118 585
R295 B.n1059 B.n1058 585
R296 B.n1060 B.n117 585
R297 B.n1062 B.n1061 585
R298 B.n1064 B.n116 585
R299 B.n1067 B.n1066 585
R300 B.n1068 B.n115 585
R301 B.n1070 B.n1069 585
R302 B.n1072 B.n114 585
R303 B.n1075 B.n1074 585
R304 B.n1076 B.n113 585
R305 B.n1078 B.n1077 585
R306 B.n1080 B.n112 585
R307 B.n1083 B.n1082 585
R308 B.n1084 B.n111 585
R309 B.n1086 B.n1085 585
R310 B.n1088 B.n110 585
R311 B.n1091 B.n1090 585
R312 B.n1092 B.n109 585
R313 B.n1094 B.n1093 585
R314 B.n1096 B.n108 585
R315 B.n1099 B.n1098 585
R316 B.n1100 B.n107 585
R317 B.n1102 B.n1101 585
R318 B.n1104 B.n106 585
R319 B.n1107 B.n1106 585
R320 B.n1108 B.n105 585
R321 B.n1110 B.n1109 585
R322 B.n1112 B.n104 585
R323 B.n1115 B.n1114 585
R324 B.n1116 B.n103 585
R325 B.n1118 B.n1117 585
R326 B.n1120 B.n102 585
R327 B.n1123 B.n1122 585
R328 B.n1124 B.n101 585
R329 B.n853 B.n99 585
R330 B.n1127 B.n99 585
R331 B.n852 B.n98 585
R332 B.n1128 B.n98 585
R333 B.n851 B.n97 585
R334 B.n1129 B.n97 585
R335 B.n850 B.n849 585
R336 B.n849 B.n93 585
R337 B.n848 B.n92 585
R338 B.n1135 B.n92 585
R339 B.n847 B.n91 585
R340 B.n1136 B.n91 585
R341 B.n846 B.n90 585
R342 B.n1137 B.n90 585
R343 B.n845 B.n844 585
R344 B.n844 B.n89 585
R345 B.n843 B.n85 585
R346 B.n1143 B.n85 585
R347 B.n842 B.n84 585
R348 B.n1144 B.n84 585
R349 B.n841 B.n83 585
R350 B.n1145 B.n83 585
R351 B.n840 B.n839 585
R352 B.n839 B.n79 585
R353 B.n838 B.n78 585
R354 B.n1151 B.n78 585
R355 B.n837 B.n77 585
R356 B.n1152 B.n77 585
R357 B.n836 B.n76 585
R358 B.n1153 B.n76 585
R359 B.n835 B.n834 585
R360 B.n834 B.n72 585
R361 B.n833 B.n71 585
R362 B.n1159 B.n71 585
R363 B.n832 B.n70 585
R364 B.n1160 B.n70 585
R365 B.n831 B.n69 585
R366 B.n1161 B.n69 585
R367 B.n830 B.n829 585
R368 B.n829 B.n65 585
R369 B.n828 B.n64 585
R370 B.n1167 B.n64 585
R371 B.n827 B.n63 585
R372 B.n1168 B.n63 585
R373 B.n826 B.n62 585
R374 B.n1169 B.n62 585
R375 B.n825 B.n824 585
R376 B.n824 B.n58 585
R377 B.n823 B.n57 585
R378 B.n1175 B.n57 585
R379 B.n822 B.n56 585
R380 B.n1176 B.n56 585
R381 B.n821 B.n55 585
R382 B.n1177 B.n55 585
R383 B.n820 B.n819 585
R384 B.n819 B.n51 585
R385 B.n818 B.n50 585
R386 B.n1183 B.n50 585
R387 B.n817 B.n49 585
R388 B.n1184 B.n49 585
R389 B.n816 B.n48 585
R390 B.n1185 B.n48 585
R391 B.n815 B.n814 585
R392 B.n814 B.n44 585
R393 B.n813 B.n43 585
R394 B.n1191 B.n43 585
R395 B.n812 B.n42 585
R396 B.n1192 B.n42 585
R397 B.n811 B.n41 585
R398 B.n1193 B.n41 585
R399 B.n810 B.n809 585
R400 B.n809 B.n37 585
R401 B.n808 B.n36 585
R402 B.n1199 B.n36 585
R403 B.n807 B.n35 585
R404 B.n1200 B.n35 585
R405 B.n806 B.n34 585
R406 B.n1201 B.n34 585
R407 B.n805 B.n804 585
R408 B.n804 B.n30 585
R409 B.n803 B.n29 585
R410 B.n1207 B.n29 585
R411 B.n802 B.n28 585
R412 B.n1208 B.n28 585
R413 B.n801 B.n27 585
R414 B.n1209 B.n27 585
R415 B.n800 B.n799 585
R416 B.n799 B.n23 585
R417 B.n798 B.n22 585
R418 B.n1215 B.n22 585
R419 B.n797 B.n21 585
R420 B.n1216 B.n21 585
R421 B.n796 B.n20 585
R422 B.n1217 B.n20 585
R423 B.n795 B.n794 585
R424 B.n794 B.n16 585
R425 B.n793 B.n15 585
R426 B.n1223 B.n15 585
R427 B.n792 B.n14 585
R428 B.n1224 B.n14 585
R429 B.n791 B.n13 585
R430 B.n1225 B.n13 585
R431 B.n790 B.n789 585
R432 B.n789 B.n12 585
R433 B.n788 B.n787 585
R434 B.n788 B.n8 585
R435 B.n786 B.n7 585
R436 B.n1232 B.n7 585
R437 B.n785 B.n6 585
R438 B.n1233 B.n6 585
R439 B.n784 B.n5 585
R440 B.n1234 B.n5 585
R441 B.n783 B.n782 585
R442 B.n782 B.n4 585
R443 B.n781 B.n173 585
R444 B.n781 B.n780 585
R445 B.n771 B.n174 585
R446 B.n175 B.n174 585
R447 B.n773 B.n772 585
R448 B.n774 B.n773 585
R449 B.n770 B.n179 585
R450 B.n183 B.n179 585
R451 B.n769 B.n768 585
R452 B.n768 B.n767 585
R453 B.n181 B.n180 585
R454 B.n182 B.n181 585
R455 B.n760 B.n759 585
R456 B.n761 B.n760 585
R457 B.n758 B.n188 585
R458 B.n188 B.n187 585
R459 B.n757 B.n756 585
R460 B.n756 B.n755 585
R461 B.n190 B.n189 585
R462 B.n191 B.n190 585
R463 B.n748 B.n747 585
R464 B.n749 B.n748 585
R465 B.n746 B.n195 585
R466 B.n199 B.n195 585
R467 B.n745 B.n744 585
R468 B.n744 B.n743 585
R469 B.n197 B.n196 585
R470 B.n198 B.n197 585
R471 B.n736 B.n735 585
R472 B.n737 B.n736 585
R473 B.n734 B.n204 585
R474 B.n204 B.n203 585
R475 B.n733 B.n732 585
R476 B.n732 B.n731 585
R477 B.n206 B.n205 585
R478 B.n207 B.n206 585
R479 B.n724 B.n723 585
R480 B.n725 B.n724 585
R481 B.n722 B.n211 585
R482 B.n215 B.n211 585
R483 B.n721 B.n720 585
R484 B.n720 B.n719 585
R485 B.n213 B.n212 585
R486 B.n214 B.n213 585
R487 B.n712 B.n711 585
R488 B.n713 B.n712 585
R489 B.n710 B.n220 585
R490 B.n220 B.n219 585
R491 B.n709 B.n708 585
R492 B.n708 B.n707 585
R493 B.n222 B.n221 585
R494 B.n223 B.n222 585
R495 B.n700 B.n699 585
R496 B.n701 B.n700 585
R497 B.n698 B.n227 585
R498 B.n231 B.n227 585
R499 B.n697 B.n696 585
R500 B.n696 B.n695 585
R501 B.n229 B.n228 585
R502 B.n230 B.n229 585
R503 B.n688 B.n687 585
R504 B.n689 B.n688 585
R505 B.n686 B.n236 585
R506 B.n236 B.n235 585
R507 B.n685 B.n684 585
R508 B.n684 B.n683 585
R509 B.n238 B.n237 585
R510 B.n239 B.n238 585
R511 B.n676 B.n675 585
R512 B.n677 B.n676 585
R513 B.n674 B.n244 585
R514 B.n244 B.n243 585
R515 B.n673 B.n672 585
R516 B.n672 B.n671 585
R517 B.n246 B.n245 585
R518 B.n247 B.n246 585
R519 B.n664 B.n663 585
R520 B.n665 B.n664 585
R521 B.n662 B.n252 585
R522 B.n252 B.n251 585
R523 B.n661 B.n660 585
R524 B.n660 B.n659 585
R525 B.n254 B.n253 585
R526 B.n255 B.n254 585
R527 B.n652 B.n651 585
R528 B.n653 B.n652 585
R529 B.n650 B.n260 585
R530 B.n260 B.n259 585
R531 B.n649 B.n648 585
R532 B.n648 B.n647 585
R533 B.n262 B.n261 585
R534 B.n640 B.n262 585
R535 B.n639 B.n638 585
R536 B.n641 B.n639 585
R537 B.n637 B.n267 585
R538 B.n267 B.n266 585
R539 B.n636 B.n635 585
R540 B.n635 B.n634 585
R541 B.n269 B.n268 585
R542 B.n270 B.n269 585
R543 B.n627 B.n626 585
R544 B.n628 B.n627 585
R545 B.n625 B.n275 585
R546 B.n275 B.n274 585
R547 B.n624 B.n623 585
R548 B.n623 B.n622 585
R549 B.n619 B.n279 585
R550 B.n618 B.n617 585
R551 B.n615 B.n280 585
R552 B.n615 B.n278 585
R553 B.n614 B.n613 585
R554 B.n612 B.n611 585
R555 B.n610 B.n282 585
R556 B.n608 B.n607 585
R557 B.n606 B.n283 585
R558 B.n605 B.n604 585
R559 B.n602 B.n284 585
R560 B.n600 B.n599 585
R561 B.n598 B.n285 585
R562 B.n597 B.n596 585
R563 B.n594 B.n286 585
R564 B.n592 B.n591 585
R565 B.n590 B.n287 585
R566 B.n589 B.n588 585
R567 B.n586 B.n288 585
R568 B.n584 B.n583 585
R569 B.n582 B.n289 585
R570 B.n581 B.n580 585
R571 B.n578 B.n290 585
R572 B.n576 B.n575 585
R573 B.n574 B.n291 585
R574 B.n573 B.n572 585
R575 B.n570 B.n292 585
R576 B.n568 B.n567 585
R577 B.n566 B.n293 585
R578 B.n565 B.n564 585
R579 B.n562 B.n294 585
R580 B.n560 B.n559 585
R581 B.n558 B.n295 585
R582 B.n557 B.n556 585
R583 B.n554 B.n296 585
R584 B.n552 B.n551 585
R585 B.n550 B.n297 585
R586 B.n549 B.n548 585
R587 B.n546 B.n298 585
R588 B.n544 B.n543 585
R589 B.n542 B.n299 585
R590 B.n541 B.n540 585
R591 B.n538 B.n300 585
R592 B.n536 B.n535 585
R593 B.n534 B.n301 585
R594 B.n533 B.n532 585
R595 B.n530 B.n302 585
R596 B.n528 B.n527 585
R597 B.n526 B.n303 585
R598 B.n525 B.n524 585
R599 B.n522 B.n304 585
R600 B.n520 B.n519 585
R601 B.n518 B.n305 585
R602 B.n517 B.n516 585
R603 B.n514 B.n306 585
R604 B.n512 B.n511 585
R605 B.n510 B.n307 585
R606 B.n509 B.n508 585
R607 B.n506 B.n308 585
R608 B.n504 B.n503 585
R609 B.n502 B.n309 585
R610 B.n501 B.n500 585
R611 B.n498 B.n310 585
R612 B.n496 B.n495 585
R613 B.n493 B.n311 585
R614 B.n492 B.n491 585
R615 B.n489 B.n314 585
R616 B.n487 B.n486 585
R617 B.n485 B.n315 585
R618 B.n484 B.n483 585
R619 B.n481 B.n316 585
R620 B.n479 B.n478 585
R621 B.n477 B.n317 585
R622 B.n475 B.n474 585
R623 B.n472 B.n320 585
R624 B.n470 B.n469 585
R625 B.n468 B.n321 585
R626 B.n467 B.n466 585
R627 B.n464 B.n322 585
R628 B.n462 B.n461 585
R629 B.n460 B.n323 585
R630 B.n459 B.n458 585
R631 B.n456 B.n324 585
R632 B.n454 B.n453 585
R633 B.n452 B.n325 585
R634 B.n451 B.n450 585
R635 B.n448 B.n326 585
R636 B.n446 B.n445 585
R637 B.n444 B.n327 585
R638 B.n443 B.n442 585
R639 B.n440 B.n328 585
R640 B.n438 B.n437 585
R641 B.n436 B.n329 585
R642 B.n435 B.n434 585
R643 B.n432 B.n330 585
R644 B.n430 B.n429 585
R645 B.n428 B.n331 585
R646 B.n427 B.n426 585
R647 B.n424 B.n332 585
R648 B.n422 B.n421 585
R649 B.n420 B.n333 585
R650 B.n419 B.n418 585
R651 B.n416 B.n334 585
R652 B.n414 B.n413 585
R653 B.n412 B.n335 585
R654 B.n411 B.n410 585
R655 B.n408 B.n336 585
R656 B.n406 B.n405 585
R657 B.n404 B.n337 585
R658 B.n403 B.n402 585
R659 B.n400 B.n338 585
R660 B.n398 B.n397 585
R661 B.n396 B.n339 585
R662 B.n395 B.n394 585
R663 B.n392 B.n340 585
R664 B.n390 B.n389 585
R665 B.n388 B.n341 585
R666 B.n387 B.n386 585
R667 B.n384 B.n342 585
R668 B.n382 B.n381 585
R669 B.n380 B.n343 585
R670 B.n379 B.n378 585
R671 B.n376 B.n344 585
R672 B.n374 B.n373 585
R673 B.n372 B.n345 585
R674 B.n371 B.n370 585
R675 B.n368 B.n346 585
R676 B.n366 B.n365 585
R677 B.n364 B.n347 585
R678 B.n363 B.n362 585
R679 B.n360 B.n348 585
R680 B.n358 B.n357 585
R681 B.n356 B.n349 585
R682 B.n355 B.n354 585
R683 B.n352 B.n350 585
R684 B.n277 B.n276 585
R685 B.n621 B.n620 585
R686 B.n622 B.n621 585
R687 B.n273 B.n272 585
R688 B.n274 B.n273 585
R689 B.n630 B.n629 585
R690 B.n629 B.n628 585
R691 B.n631 B.n271 585
R692 B.n271 B.n270 585
R693 B.n633 B.n632 585
R694 B.n634 B.n633 585
R695 B.n265 B.n264 585
R696 B.n266 B.n265 585
R697 B.n643 B.n642 585
R698 B.n642 B.n641 585
R699 B.n644 B.n263 585
R700 B.n640 B.n263 585
R701 B.n646 B.n645 585
R702 B.n647 B.n646 585
R703 B.n258 B.n257 585
R704 B.n259 B.n258 585
R705 B.n655 B.n654 585
R706 B.n654 B.n653 585
R707 B.n656 B.n256 585
R708 B.n256 B.n255 585
R709 B.n658 B.n657 585
R710 B.n659 B.n658 585
R711 B.n250 B.n249 585
R712 B.n251 B.n250 585
R713 B.n667 B.n666 585
R714 B.n666 B.n665 585
R715 B.n668 B.n248 585
R716 B.n248 B.n247 585
R717 B.n670 B.n669 585
R718 B.n671 B.n670 585
R719 B.n242 B.n241 585
R720 B.n243 B.n242 585
R721 B.n679 B.n678 585
R722 B.n678 B.n677 585
R723 B.n680 B.n240 585
R724 B.n240 B.n239 585
R725 B.n682 B.n681 585
R726 B.n683 B.n682 585
R727 B.n234 B.n233 585
R728 B.n235 B.n234 585
R729 B.n691 B.n690 585
R730 B.n690 B.n689 585
R731 B.n692 B.n232 585
R732 B.n232 B.n230 585
R733 B.n694 B.n693 585
R734 B.n695 B.n694 585
R735 B.n226 B.n225 585
R736 B.n231 B.n226 585
R737 B.n703 B.n702 585
R738 B.n702 B.n701 585
R739 B.n704 B.n224 585
R740 B.n224 B.n223 585
R741 B.n706 B.n705 585
R742 B.n707 B.n706 585
R743 B.n218 B.n217 585
R744 B.n219 B.n218 585
R745 B.n715 B.n714 585
R746 B.n714 B.n713 585
R747 B.n716 B.n216 585
R748 B.n216 B.n214 585
R749 B.n718 B.n717 585
R750 B.n719 B.n718 585
R751 B.n210 B.n209 585
R752 B.n215 B.n210 585
R753 B.n727 B.n726 585
R754 B.n726 B.n725 585
R755 B.n728 B.n208 585
R756 B.n208 B.n207 585
R757 B.n730 B.n729 585
R758 B.n731 B.n730 585
R759 B.n202 B.n201 585
R760 B.n203 B.n202 585
R761 B.n739 B.n738 585
R762 B.n738 B.n737 585
R763 B.n740 B.n200 585
R764 B.n200 B.n198 585
R765 B.n742 B.n741 585
R766 B.n743 B.n742 585
R767 B.n194 B.n193 585
R768 B.n199 B.n194 585
R769 B.n751 B.n750 585
R770 B.n750 B.n749 585
R771 B.n752 B.n192 585
R772 B.n192 B.n191 585
R773 B.n754 B.n753 585
R774 B.n755 B.n754 585
R775 B.n186 B.n185 585
R776 B.n187 B.n186 585
R777 B.n763 B.n762 585
R778 B.n762 B.n761 585
R779 B.n764 B.n184 585
R780 B.n184 B.n182 585
R781 B.n766 B.n765 585
R782 B.n767 B.n766 585
R783 B.n178 B.n177 585
R784 B.n183 B.n178 585
R785 B.n776 B.n775 585
R786 B.n775 B.n774 585
R787 B.n777 B.n176 585
R788 B.n176 B.n175 585
R789 B.n779 B.n778 585
R790 B.n780 B.n779 585
R791 B.n3 B.n0 585
R792 B.n4 B.n3 585
R793 B.n1231 B.n1 585
R794 B.n1232 B.n1231 585
R795 B.n1230 B.n1229 585
R796 B.n1230 B.n8 585
R797 B.n1228 B.n9 585
R798 B.n12 B.n9 585
R799 B.n1227 B.n1226 585
R800 B.n1226 B.n1225 585
R801 B.n11 B.n10 585
R802 B.n1224 B.n11 585
R803 B.n1222 B.n1221 585
R804 B.n1223 B.n1222 585
R805 B.n1220 B.n17 585
R806 B.n17 B.n16 585
R807 B.n1219 B.n1218 585
R808 B.n1218 B.n1217 585
R809 B.n19 B.n18 585
R810 B.n1216 B.n19 585
R811 B.n1214 B.n1213 585
R812 B.n1215 B.n1214 585
R813 B.n1212 B.n24 585
R814 B.n24 B.n23 585
R815 B.n1211 B.n1210 585
R816 B.n1210 B.n1209 585
R817 B.n26 B.n25 585
R818 B.n1208 B.n26 585
R819 B.n1206 B.n1205 585
R820 B.n1207 B.n1206 585
R821 B.n1204 B.n31 585
R822 B.n31 B.n30 585
R823 B.n1203 B.n1202 585
R824 B.n1202 B.n1201 585
R825 B.n33 B.n32 585
R826 B.n1200 B.n33 585
R827 B.n1198 B.n1197 585
R828 B.n1199 B.n1198 585
R829 B.n1196 B.n38 585
R830 B.n38 B.n37 585
R831 B.n1195 B.n1194 585
R832 B.n1194 B.n1193 585
R833 B.n40 B.n39 585
R834 B.n1192 B.n40 585
R835 B.n1190 B.n1189 585
R836 B.n1191 B.n1190 585
R837 B.n1188 B.n45 585
R838 B.n45 B.n44 585
R839 B.n1187 B.n1186 585
R840 B.n1186 B.n1185 585
R841 B.n47 B.n46 585
R842 B.n1184 B.n47 585
R843 B.n1182 B.n1181 585
R844 B.n1183 B.n1182 585
R845 B.n1180 B.n52 585
R846 B.n52 B.n51 585
R847 B.n1179 B.n1178 585
R848 B.n1178 B.n1177 585
R849 B.n54 B.n53 585
R850 B.n1176 B.n54 585
R851 B.n1174 B.n1173 585
R852 B.n1175 B.n1174 585
R853 B.n1172 B.n59 585
R854 B.n59 B.n58 585
R855 B.n1171 B.n1170 585
R856 B.n1170 B.n1169 585
R857 B.n61 B.n60 585
R858 B.n1168 B.n61 585
R859 B.n1166 B.n1165 585
R860 B.n1167 B.n1166 585
R861 B.n1164 B.n66 585
R862 B.n66 B.n65 585
R863 B.n1163 B.n1162 585
R864 B.n1162 B.n1161 585
R865 B.n68 B.n67 585
R866 B.n1160 B.n68 585
R867 B.n1158 B.n1157 585
R868 B.n1159 B.n1158 585
R869 B.n1156 B.n73 585
R870 B.n73 B.n72 585
R871 B.n1155 B.n1154 585
R872 B.n1154 B.n1153 585
R873 B.n75 B.n74 585
R874 B.n1152 B.n75 585
R875 B.n1150 B.n1149 585
R876 B.n1151 B.n1150 585
R877 B.n1148 B.n80 585
R878 B.n80 B.n79 585
R879 B.n1147 B.n1146 585
R880 B.n1146 B.n1145 585
R881 B.n82 B.n81 585
R882 B.n1144 B.n82 585
R883 B.n1142 B.n1141 585
R884 B.n1143 B.n1142 585
R885 B.n1140 B.n86 585
R886 B.n89 B.n86 585
R887 B.n1139 B.n1138 585
R888 B.n1138 B.n1137 585
R889 B.n88 B.n87 585
R890 B.n1136 B.n88 585
R891 B.n1134 B.n1133 585
R892 B.n1135 B.n1134 585
R893 B.n1132 B.n94 585
R894 B.n94 B.n93 585
R895 B.n1131 B.n1130 585
R896 B.n1130 B.n1129 585
R897 B.n96 B.n95 585
R898 B.n1128 B.n96 585
R899 B.n1126 B.n1125 585
R900 B.n1127 B.n1126 585
R901 B.n1235 B.n1234 585
R902 B.n1233 B.n2 585
R903 B.n1126 B.n101 473.281
R904 B.n855 B.n99 473.281
R905 B.n623 B.n277 473.281
R906 B.n621 B.n279 473.281
R907 B.n134 B.t21 409.272
R908 B.n141 B.t17 409.272
R909 B.n318 B.t10 409.272
R910 B.n312 B.t14 409.272
R911 B.n856 B.n100 256.663
R912 B.n862 B.n100 256.663
R913 B.n864 B.n100 256.663
R914 B.n870 B.n100 256.663
R915 B.n872 B.n100 256.663
R916 B.n878 B.n100 256.663
R917 B.n880 B.n100 256.663
R918 B.n886 B.n100 256.663
R919 B.n888 B.n100 256.663
R920 B.n894 B.n100 256.663
R921 B.n896 B.n100 256.663
R922 B.n902 B.n100 256.663
R923 B.n904 B.n100 256.663
R924 B.n910 B.n100 256.663
R925 B.n912 B.n100 256.663
R926 B.n918 B.n100 256.663
R927 B.n920 B.n100 256.663
R928 B.n926 B.n100 256.663
R929 B.n928 B.n100 256.663
R930 B.n934 B.n100 256.663
R931 B.n936 B.n100 256.663
R932 B.n942 B.n100 256.663
R933 B.n944 B.n100 256.663
R934 B.n950 B.n100 256.663
R935 B.n952 B.n100 256.663
R936 B.n958 B.n100 256.663
R937 B.n960 B.n100 256.663
R938 B.n966 B.n100 256.663
R939 B.n968 B.n100 256.663
R940 B.n974 B.n100 256.663
R941 B.n976 B.n100 256.663
R942 B.n983 B.n100 256.663
R943 B.n985 B.n100 256.663
R944 B.n991 B.n100 256.663
R945 B.n993 B.n100 256.663
R946 B.n999 B.n100 256.663
R947 B.n1001 B.n100 256.663
R948 B.n1007 B.n100 256.663
R949 B.n1009 B.n100 256.663
R950 B.n1015 B.n100 256.663
R951 B.n1017 B.n100 256.663
R952 B.n1023 B.n100 256.663
R953 B.n1025 B.n100 256.663
R954 B.n1031 B.n100 256.663
R955 B.n1033 B.n100 256.663
R956 B.n1039 B.n100 256.663
R957 B.n1041 B.n100 256.663
R958 B.n1047 B.n100 256.663
R959 B.n1049 B.n100 256.663
R960 B.n1055 B.n100 256.663
R961 B.n1057 B.n100 256.663
R962 B.n1063 B.n100 256.663
R963 B.n1065 B.n100 256.663
R964 B.n1071 B.n100 256.663
R965 B.n1073 B.n100 256.663
R966 B.n1079 B.n100 256.663
R967 B.n1081 B.n100 256.663
R968 B.n1087 B.n100 256.663
R969 B.n1089 B.n100 256.663
R970 B.n1095 B.n100 256.663
R971 B.n1097 B.n100 256.663
R972 B.n1103 B.n100 256.663
R973 B.n1105 B.n100 256.663
R974 B.n1111 B.n100 256.663
R975 B.n1113 B.n100 256.663
R976 B.n1119 B.n100 256.663
R977 B.n1121 B.n100 256.663
R978 B.n616 B.n278 256.663
R979 B.n281 B.n278 256.663
R980 B.n609 B.n278 256.663
R981 B.n603 B.n278 256.663
R982 B.n601 B.n278 256.663
R983 B.n595 B.n278 256.663
R984 B.n593 B.n278 256.663
R985 B.n587 B.n278 256.663
R986 B.n585 B.n278 256.663
R987 B.n579 B.n278 256.663
R988 B.n577 B.n278 256.663
R989 B.n571 B.n278 256.663
R990 B.n569 B.n278 256.663
R991 B.n563 B.n278 256.663
R992 B.n561 B.n278 256.663
R993 B.n555 B.n278 256.663
R994 B.n553 B.n278 256.663
R995 B.n547 B.n278 256.663
R996 B.n545 B.n278 256.663
R997 B.n539 B.n278 256.663
R998 B.n537 B.n278 256.663
R999 B.n531 B.n278 256.663
R1000 B.n529 B.n278 256.663
R1001 B.n523 B.n278 256.663
R1002 B.n521 B.n278 256.663
R1003 B.n515 B.n278 256.663
R1004 B.n513 B.n278 256.663
R1005 B.n507 B.n278 256.663
R1006 B.n505 B.n278 256.663
R1007 B.n499 B.n278 256.663
R1008 B.n497 B.n278 256.663
R1009 B.n490 B.n278 256.663
R1010 B.n488 B.n278 256.663
R1011 B.n482 B.n278 256.663
R1012 B.n480 B.n278 256.663
R1013 B.n473 B.n278 256.663
R1014 B.n471 B.n278 256.663
R1015 B.n465 B.n278 256.663
R1016 B.n463 B.n278 256.663
R1017 B.n457 B.n278 256.663
R1018 B.n455 B.n278 256.663
R1019 B.n449 B.n278 256.663
R1020 B.n447 B.n278 256.663
R1021 B.n441 B.n278 256.663
R1022 B.n439 B.n278 256.663
R1023 B.n433 B.n278 256.663
R1024 B.n431 B.n278 256.663
R1025 B.n425 B.n278 256.663
R1026 B.n423 B.n278 256.663
R1027 B.n417 B.n278 256.663
R1028 B.n415 B.n278 256.663
R1029 B.n409 B.n278 256.663
R1030 B.n407 B.n278 256.663
R1031 B.n401 B.n278 256.663
R1032 B.n399 B.n278 256.663
R1033 B.n393 B.n278 256.663
R1034 B.n391 B.n278 256.663
R1035 B.n385 B.n278 256.663
R1036 B.n383 B.n278 256.663
R1037 B.n377 B.n278 256.663
R1038 B.n375 B.n278 256.663
R1039 B.n369 B.n278 256.663
R1040 B.n367 B.n278 256.663
R1041 B.n361 B.n278 256.663
R1042 B.n359 B.n278 256.663
R1043 B.n353 B.n278 256.663
R1044 B.n351 B.n278 256.663
R1045 B.n1237 B.n1236 256.663
R1046 B.n1122 B.n1120 163.367
R1047 B.n1118 B.n103 163.367
R1048 B.n1114 B.n1112 163.367
R1049 B.n1110 B.n105 163.367
R1050 B.n1106 B.n1104 163.367
R1051 B.n1102 B.n107 163.367
R1052 B.n1098 B.n1096 163.367
R1053 B.n1094 B.n109 163.367
R1054 B.n1090 B.n1088 163.367
R1055 B.n1086 B.n111 163.367
R1056 B.n1082 B.n1080 163.367
R1057 B.n1078 B.n113 163.367
R1058 B.n1074 B.n1072 163.367
R1059 B.n1070 B.n115 163.367
R1060 B.n1066 B.n1064 163.367
R1061 B.n1062 B.n117 163.367
R1062 B.n1058 B.n1056 163.367
R1063 B.n1054 B.n119 163.367
R1064 B.n1050 B.n1048 163.367
R1065 B.n1046 B.n121 163.367
R1066 B.n1042 B.n1040 163.367
R1067 B.n1038 B.n123 163.367
R1068 B.n1034 B.n1032 163.367
R1069 B.n1030 B.n125 163.367
R1070 B.n1026 B.n1024 163.367
R1071 B.n1022 B.n127 163.367
R1072 B.n1018 B.n1016 163.367
R1073 B.n1014 B.n129 163.367
R1074 B.n1010 B.n1008 163.367
R1075 B.n1006 B.n131 163.367
R1076 B.n1002 B.n1000 163.367
R1077 B.n998 B.n133 163.367
R1078 B.n994 B.n992 163.367
R1079 B.n990 B.n138 163.367
R1080 B.n986 B.n984 163.367
R1081 B.n982 B.n140 163.367
R1082 B.n977 B.n975 163.367
R1083 B.n973 B.n144 163.367
R1084 B.n969 B.n967 163.367
R1085 B.n965 B.n146 163.367
R1086 B.n961 B.n959 163.367
R1087 B.n957 B.n148 163.367
R1088 B.n953 B.n951 163.367
R1089 B.n949 B.n150 163.367
R1090 B.n945 B.n943 163.367
R1091 B.n941 B.n152 163.367
R1092 B.n937 B.n935 163.367
R1093 B.n933 B.n154 163.367
R1094 B.n929 B.n927 163.367
R1095 B.n925 B.n156 163.367
R1096 B.n921 B.n919 163.367
R1097 B.n917 B.n158 163.367
R1098 B.n913 B.n911 163.367
R1099 B.n909 B.n160 163.367
R1100 B.n905 B.n903 163.367
R1101 B.n901 B.n162 163.367
R1102 B.n897 B.n895 163.367
R1103 B.n893 B.n164 163.367
R1104 B.n889 B.n887 163.367
R1105 B.n885 B.n166 163.367
R1106 B.n881 B.n879 163.367
R1107 B.n877 B.n168 163.367
R1108 B.n873 B.n871 163.367
R1109 B.n869 B.n170 163.367
R1110 B.n865 B.n863 163.367
R1111 B.n861 B.n172 163.367
R1112 B.n857 B.n855 163.367
R1113 B.n623 B.n275 163.367
R1114 B.n627 B.n275 163.367
R1115 B.n627 B.n269 163.367
R1116 B.n635 B.n269 163.367
R1117 B.n635 B.n267 163.367
R1118 B.n639 B.n267 163.367
R1119 B.n639 B.n262 163.367
R1120 B.n648 B.n262 163.367
R1121 B.n648 B.n260 163.367
R1122 B.n652 B.n260 163.367
R1123 B.n652 B.n254 163.367
R1124 B.n660 B.n254 163.367
R1125 B.n660 B.n252 163.367
R1126 B.n664 B.n252 163.367
R1127 B.n664 B.n246 163.367
R1128 B.n672 B.n246 163.367
R1129 B.n672 B.n244 163.367
R1130 B.n676 B.n244 163.367
R1131 B.n676 B.n238 163.367
R1132 B.n684 B.n238 163.367
R1133 B.n684 B.n236 163.367
R1134 B.n688 B.n236 163.367
R1135 B.n688 B.n229 163.367
R1136 B.n696 B.n229 163.367
R1137 B.n696 B.n227 163.367
R1138 B.n700 B.n227 163.367
R1139 B.n700 B.n222 163.367
R1140 B.n708 B.n222 163.367
R1141 B.n708 B.n220 163.367
R1142 B.n712 B.n220 163.367
R1143 B.n712 B.n213 163.367
R1144 B.n720 B.n213 163.367
R1145 B.n720 B.n211 163.367
R1146 B.n724 B.n211 163.367
R1147 B.n724 B.n206 163.367
R1148 B.n732 B.n206 163.367
R1149 B.n732 B.n204 163.367
R1150 B.n736 B.n204 163.367
R1151 B.n736 B.n197 163.367
R1152 B.n744 B.n197 163.367
R1153 B.n744 B.n195 163.367
R1154 B.n748 B.n195 163.367
R1155 B.n748 B.n190 163.367
R1156 B.n756 B.n190 163.367
R1157 B.n756 B.n188 163.367
R1158 B.n760 B.n188 163.367
R1159 B.n760 B.n181 163.367
R1160 B.n768 B.n181 163.367
R1161 B.n768 B.n179 163.367
R1162 B.n773 B.n179 163.367
R1163 B.n773 B.n174 163.367
R1164 B.n781 B.n174 163.367
R1165 B.n782 B.n781 163.367
R1166 B.n782 B.n5 163.367
R1167 B.n6 B.n5 163.367
R1168 B.n7 B.n6 163.367
R1169 B.n788 B.n7 163.367
R1170 B.n789 B.n788 163.367
R1171 B.n789 B.n13 163.367
R1172 B.n14 B.n13 163.367
R1173 B.n15 B.n14 163.367
R1174 B.n794 B.n15 163.367
R1175 B.n794 B.n20 163.367
R1176 B.n21 B.n20 163.367
R1177 B.n22 B.n21 163.367
R1178 B.n799 B.n22 163.367
R1179 B.n799 B.n27 163.367
R1180 B.n28 B.n27 163.367
R1181 B.n29 B.n28 163.367
R1182 B.n804 B.n29 163.367
R1183 B.n804 B.n34 163.367
R1184 B.n35 B.n34 163.367
R1185 B.n36 B.n35 163.367
R1186 B.n809 B.n36 163.367
R1187 B.n809 B.n41 163.367
R1188 B.n42 B.n41 163.367
R1189 B.n43 B.n42 163.367
R1190 B.n814 B.n43 163.367
R1191 B.n814 B.n48 163.367
R1192 B.n49 B.n48 163.367
R1193 B.n50 B.n49 163.367
R1194 B.n819 B.n50 163.367
R1195 B.n819 B.n55 163.367
R1196 B.n56 B.n55 163.367
R1197 B.n57 B.n56 163.367
R1198 B.n824 B.n57 163.367
R1199 B.n824 B.n62 163.367
R1200 B.n63 B.n62 163.367
R1201 B.n64 B.n63 163.367
R1202 B.n829 B.n64 163.367
R1203 B.n829 B.n69 163.367
R1204 B.n70 B.n69 163.367
R1205 B.n71 B.n70 163.367
R1206 B.n834 B.n71 163.367
R1207 B.n834 B.n76 163.367
R1208 B.n77 B.n76 163.367
R1209 B.n78 B.n77 163.367
R1210 B.n839 B.n78 163.367
R1211 B.n839 B.n83 163.367
R1212 B.n84 B.n83 163.367
R1213 B.n85 B.n84 163.367
R1214 B.n844 B.n85 163.367
R1215 B.n844 B.n90 163.367
R1216 B.n91 B.n90 163.367
R1217 B.n92 B.n91 163.367
R1218 B.n849 B.n92 163.367
R1219 B.n849 B.n97 163.367
R1220 B.n98 B.n97 163.367
R1221 B.n99 B.n98 163.367
R1222 B.n617 B.n615 163.367
R1223 B.n615 B.n614 163.367
R1224 B.n611 B.n610 163.367
R1225 B.n608 B.n283 163.367
R1226 B.n604 B.n602 163.367
R1227 B.n600 B.n285 163.367
R1228 B.n596 B.n594 163.367
R1229 B.n592 B.n287 163.367
R1230 B.n588 B.n586 163.367
R1231 B.n584 B.n289 163.367
R1232 B.n580 B.n578 163.367
R1233 B.n576 B.n291 163.367
R1234 B.n572 B.n570 163.367
R1235 B.n568 B.n293 163.367
R1236 B.n564 B.n562 163.367
R1237 B.n560 B.n295 163.367
R1238 B.n556 B.n554 163.367
R1239 B.n552 B.n297 163.367
R1240 B.n548 B.n546 163.367
R1241 B.n544 B.n299 163.367
R1242 B.n540 B.n538 163.367
R1243 B.n536 B.n301 163.367
R1244 B.n532 B.n530 163.367
R1245 B.n528 B.n303 163.367
R1246 B.n524 B.n522 163.367
R1247 B.n520 B.n305 163.367
R1248 B.n516 B.n514 163.367
R1249 B.n512 B.n307 163.367
R1250 B.n508 B.n506 163.367
R1251 B.n504 B.n309 163.367
R1252 B.n500 B.n498 163.367
R1253 B.n496 B.n311 163.367
R1254 B.n491 B.n489 163.367
R1255 B.n487 B.n315 163.367
R1256 B.n483 B.n481 163.367
R1257 B.n479 B.n317 163.367
R1258 B.n474 B.n472 163.367
R1259 B.n470 B.n321 163.367
R1260 B.n466 B.n464 163.367
R1261 B.n462 B.n323 163.367
R1262 B.n458 B.n456 163.367
R1263 B.n454 B.n325 163.367
R1264 B.n450 B.n448 163.367
R1265 B.n446 B.n327 163.367
R1266 B.n442 B.n440 163.367
R1267 B.n438 B.n329 163.367
R1268 B.n434 B.n432 163.367
R1269 B.n430 B.n331 163.367
R1270 B.n426 B.n424 163.367
R1271 B.n422 B.n333 163.367
R1272 B.n418 B.n416 163.367
R1273 B.n414 B.n335 163.367
R1274 B.n410 B.n408 163.367
R1275 B.n406 B.n337 163.367
R1276 B.n402 B.n400 163.367
R1277 B.n398 B.n339 163.367
R1278 B.n394 B.n392 163.367
R1279 B.n390 B.n341 163.367
R1280 B.n386 B.n384 163.367
R1281 B.n382 B.n343 163.367
R1282 B.n378 B.n376 163.367
R1283 B.n374 B.n345 163.367
R1284 B.n370 B.n368 163.367
R1285 B.n366 B.n347 163.367
R1286 B.n362 B.n360 163.367
R1287 B.n358 B.n349 163.367
R1288 B.n354 B.n352 163.367
R1289 B.n621 B.n273 163.367
R1290 B.n629 B.n273 163.367
R1291 B.n629 B.n271 163.367
R1292 B.n633 B.n271 163.367
R1293 B.n633 B.n265 163.367
R1294 B.n642 B.n265 163.367
R1295 B.n642 B.n263 163.367
R1296 B.n646 B.n263 163.367
R1297 B.n646 B.n258 163.367
R1298 B.n654 B.n258 163.367
R1299 B.n654 B.n256 163.367
R1300 B.n658 B.n256 163.367
R1301 B.n658 B.n250 163.367
R1302 B.n666 B.n250 163.367
R1303 B.n666 B.n248 163.367
R1304 B.n670 B.n248 163.367
R1305 B.n670 B.n242 163.367
R1306 B.n678 B.n242 163.367
R1307 B.n678 B.n240 163.367
R1308 B.n682 B.n240 163.367
R1309 B.n682 B.n234 163.367
R1310 B.n690 B.n234 163.367
R1311 B.n690 B.n232 163.367
R1312 B.n694 B.n232 163.367
R1313 B.n694 B.n226 163.367
R1314 B.n702 B.n226 163.367
R1315 B.n702 B.n224 163.367
R1316 B.n706 B.n224 163.367
R1317 B.n706 B.n218 163.367
R1318 B.n714 B.n218 163.367
R1319 B.n714 B.n216 163.367
R1320 B.n718 B.n216 163.367
R1321 B.n718 B.n210 163.367
R1322 B.n726 B.n210 163.367
R1323 B.n726 B.n208 163.367
R1324 B.n730 B.n208 163.367
R1325 B.n730 B.n202 163.367
R1326 B.n738 B.n202 163.367
R1327 B.n738 B.n200 163.367
R1328 B.n742 B.n200 163.367
R1329 B.n742 B.n194 163.367
R1330 B.n750 B.n194 163.367
R1331 B.n750 B.n192 163.367
R1332 B.n754 B.n192 163.367
R1333 B.n754 B.n186 163.367
R1334 B.n762 B.n186 163.367
R1335 B.n762 B.n184 163.367
R1336 B.n766 B.n184 163.367
R1337 B.n766 B.n178 163.367
R1338 B.n775 B.n178 163.367
R1339 B.n775 B.n176 163.367
R1340 B.n779 B.n176 163.367
R1341 B.n779 B.n3 163.367
R1342 B.n1235 B.n3 163.367
R1343 B.n1231 B.n2 163.367
R1344 B.n1231 B.n1230 163.367
R1345 B.n1230 B.n9 163.367
R1346 B.n1226 B.n9 163.367
R1347 B.n1226 B.n11 163.367
R1348 B.n1222 B.n11 163.367
R1349 B.n1222 B.n17 163.367
R1350 B.n1218 B.n17 163.367
R1351 B.n1218 B.n19 163.367
R1352 B.n1214 B.n19 163.367
R1353 B.n1214 B.n24 163.367
R1354 B.n1210 B.n24 163.367
R1355 B.n1210 B.n26 163.367
R1356 B.n1206 B.n26 163.367
R1357 B.n1206 B.n31 163.367
R1358 B.n1202 B.n31 163.367
R1359 B.n1202 B.n33 163.367
R1360 B.n1198 B.n33 163.367
R1361 B.n1198 B.n38 163.367
R1362 B.n1194 B.n38 163.367
R1363 B.n1194 B.n40 163.367
R1364 B.n1190 B.n40 163.367
R1365 B.n1190 B.n45 163.367
R1366 B.n1186 B.n45 163.367
R1367 B.n1186 B.n47 163.367
R1368 B.n1182 B.n47 163.367
R1369 B.n1182 B.n52 163.367
R1370 B.n1178 B.n52 163.367
R1371 B.n1178 B.n54 163.367
R1372 B.n1174 B.n54 163.367
R1373 B.n1174 B.n59 163.367
R1374 B.n1170 B.n59 163.367
R1375 B.n1170 B.n61 163.367
R1376 B.n1166 B.n61 163.367
R1377 B.n1166 B.n66 163.367
R1378 B.n1162 B.n66 163.367
R1379 B.n1162 B.n68 163.367
R1380 B.n1158 B.n68 163.367
R1381 B.n1158 B.n73 163.367
R1382 B.n1154 B.n73 163.367
R1383 B.n1154 B.n75 163.367
R1384 B.n1150 B.n75 163.367
R1385 B.n1150 B.n80 163.367
R1386 B.n1146 B.n80 163.367
R1387 B.n1146 B.n82 163.367
R1388 B.n1142 B.n82 163.367
R1389 B.n1142 B.n86 163.367
R1390 B.n1138 B.n86 163.367
R1391 B.n1138 B.n88 163.367
R1392 B.n1134 B.n88 163.367
R1393 B.n1134 B.n94 163.367
R1394 B.n1130 B.n94 163.367
R1395 B.n1130 B.n96 163.367
R1396 B.n1126 B.n96 163.367
R1397 B.n141 B.t19 120.516
R1398 B.n318 B.t13 120.516
R1399 B.n134 B.t22 120.49
R1400 B.n312 B.t16 120.49
R1401 B.n1121 B.n101 71.676
R1402 B.n1120 B.n1119 71.676
R1403 B.n1113 B.n103 71.676
R1404 B.n1112 B.n1111 71.676
R1405 B.n1105 B.n105 71.676
R1406 B.n1104 B.n1103 71.676
R1407 B.n1097 B.n107 71.676
R1408 B.n1096 B.n1095 71.676
R1409 B.n1089 B.n109 71.676
R1410 B.n1088 B.n1087 71.676
R1411 B.n1081 B.n111 71.676
R1412 B.n1080 B.n1079 71.676
R1413 B.n1073 B.n113 71.676
R1414 B.n1072 B.n1071 71.676
R1415 B.n1065 B.n115 71.676
R1416 B.n1064 B.n1063 71.676
R1417 B.n1057 B.n117 71.676
R1418 B.n1056 B.n1055 71.676
R1419 B.n1049 B.n119 71.676
R1420 B.n1048 B.n1047 71.676
R1421 B.n1041 B.n121 71.676
R1422 B.n1040 B.n1039 71.676
R1423 B.n1033 B.n123 71.676
R1424 B.n1032 B.n1031 71.676
R1425 B.n1025 B.n125 71.676
R1426 B.n1024 B.n1023 71.676
R1427 B.n1017 B.n127 71.676
R1428 B.n1016 B.n1015 71.676
R1429 B.n1009 B.n129 71.676
R1430 B.n1008 B.n1007 71.676
R1431 B.n1001 B.n131 71.676
R1432 B.n1000 B.n999 71.676
R1433 B.n993 B.n133 71.676
R1434 B.n992 B.n991 71.676
R1435 B.n985 B.n138 71.676
R1436 B.n984 B.n983 71.676
R1437 B.n976 B.n140 71.676
R1438 B.n975 B.n974 71.676
R1439 B.n968 B.n144 71.676
R1440 B.n967 B.n966 71.676
R1441 B.n960 B.n146 71.676
R1442 B.n959 B.n958 71.676
R1443 B.n952 B.n148 71.676
R1444 B.n951 B.n950 71.676
R1445 B.n944 B.n150 71.676
R1446 B.n943 B.n942 71.676
R1447 B.n936 B.n152 71.676
R1448 B.n935 B.n934 71.676
R1449 B.n928 B.n154 71.676
R1450 B.n927 B.n926 71.676
R1451 B.n920 B.n156 71.676
R1452 B.n919 B.n918 71.676
R1453 B.n912 B.n158 71.676
R1454 B.n911 B.n910 71.676
R1455 B.n904 B.n160 71.676
R1456 B.n903 B.n902 71.676
R1457 B.n896 B.n162 71.676
R1458 B.n895 B.n894 71.676
R1459 B.n888 B.n164 71.676
R1460 B.n887 B.n886 71.676
R1461 B.n880 B.n166 71.676
R1462 B.n879 B.n878 71.676
R1463 B.n872 B.n168 71.676
R1464 B.n871 B.n870 71.676
R1465 B.n864 B.n170 71.676
R1466 B.n863 B.n862 71.676
R1467 B.n856 B.n172 71.676
R1468 B.n857 B.n856 71.676
R1469 B.n862 B.n861 71.676
R1470 B.n865 B.n864 71.676
R1471 B.n870 B.n869 71.676
R1472 B.n873 B.n872 71.676
R1473 B.n878 B.n877 71.676
R1474 B.n881 B.n880 71.676
R1475 B.n886 B.n885 71.676
R1476 B.n889 B.n888 71.676
R1477 B.n894 B.n893 71.676
R1478 B.n897 B.n896 71.676
R1479 B.n902 B.n901 71.676
R1480 B.n905 B.n904 71.676
R1481 B.n910 B.n909 71.676
R1482 B.n913 B.n912 71.676
R1483 B.n918 B.n917 71.676
R1484 B.n921 B.n920 71.676
R1485 B.n926 B.n925 71.676
R1486 B.n929 B.n928 71.676
R1487 B.n934 B.n933 71.676
R1488 B.n937 B.n936 71.676
R1489 B.n942 B.n941 71.676
R1490 B.n945 B.n944 71.676
R1491 B.n950 B.n949 71.676
R1492 B.n953 B.n952 71.676
R1493 B.n958 B.n957 71.676
R1494 B.n961 B.n960 71.676
R1495 B.n966 B.n965 71.676
R1496 B.n969 B.n968 71.676
R1497 B.n974 B.n973 71.676
R1498 B.n977 B.n976 71.676
R1499 B.n983 B.n982 71.676
R1500 B.n986 B.n985 71.676
R1501 B.n991 B.n990 71.676
R1502 B.n994 B.n993 71.676
R1503 B.n999 B.n998 71.676
R1504 B.n1002 B.n1001 71.676
R1505 B.n1007 B.n1006 71.676
R1506 B.n1010 B.n1009 71.676
R1507 B.n1015 B.n1014 71.676
R1508 B.n1018 B.n1017 71.676
R1509 B.n1023 B.n1022 71.676
R1510 B.n1026 B.n1025 71.676
R1511 B.n1031 B.n1030 71.676
R1512 B.n1034 B.n1033 71.676
R1513 B.n1039 B.n1038 71.676
R1514 B.n1042 B.n1041 71.676
R1515 B.n1047 B.n1046 71.676
R1516 B.n1050 B.n1049 71.676
R1517 B.n1055 B.n1054 71.676
R1518 B.n1058 B.n1057 71.676
R1519 B.n1063 B.n1062 71.676
R1520 B.n1066 B.n1065 71.676
R1521 B.n1071 B.n1070 71.676
R1522 B.n1074 B.n1073 71.676
R1523 B.n1079 B.n1078 71.676
R1524 B.n1082 B.n1081 71.676
R1525 B.n1087 B.n1086 71.676
R1526 B.n1090 B.n1089 71.676
R1527 B.n1095 B.n1094 71.676
R1528 B.n1098 B.n1097 71.676
R1529 B.n1103 B.n1102 71.676
R1530 B.n1106 B.n1105 71.676
R1531 B.n1111 B.n1110 71.676
R1532 B.n1114 B.n1113 71.676
R1533 B.n1119 B.n1118 71.676
R1534 B.n1122 B.n1121 71.676
R1535 B.n616 B.n279 71.676
R1536 B.n614 B.n281 71.676
R1537 B.n610 B.n609 71.676
R1538 B.n603 B.n283 71.676
R1539 B.n602 B.n601 71.676
R1540 B.n595 B.n285 71.676
R1541 B.n594 B.n593 71.676
R1542 B.n587 B.n287 71.676
R1543 B.n586 B.n585 71.676
R1544 B.n579 B.n289 71.676
R1545 B.n578 B.n577 71.676
R1546 B.n571 B.n291 71.676
R1547 B.n570 B.n569 71.676
R1548 B.n563 B.n293 71.676
R1549 B.n562 B.n561 71.676
R1550 B.n555 B.n295 71.676
R1551 B.n554 B.n553 71.676
R1552 B.n547 B.n297 71.676
R1553 B.n546 B.n545 71.676
R1554 B.n539 B.n299 71.676
R1555 B.n538 B.n537 71.676
R1556 B.n531 B.n301 71.676
R1557 B.n530 B.n529 71.676
R1558 B.n523 B.n303 71.676
R1559 B.n522 B.n521 71.676
R1560 B.n515 B.n305 71.676
R1561 B.n514 B.n513 71.676
R1562 B.n507 B.n307 71.676
R1563 B.n506 B.n505 71.676
R1564 B.n499 B.n309 71.676
R1565 B.n498 B.n497 71.676
R1566 B.n490 B.n311 71.676
R1567 B.n489 B.n488 71.676
R1568 B.n482 B.n315 71.676
R1569 B.n481 B.n480 71.676
R1570 B.n473 B.n317 71.676
R1571 B.n472 B.n471 71.676
R1572 B.n465 B.n321 71.676
R1573 B.n464 B.n463 71.676
R1574 B.n457 B.n323 71.676
R1575 B.n456 B.n455 71.676
R1576 B.n449 B.n325 71.676
R1577 B.n448 B.n447 71.676
R1578 B.n441 B.n327 71.676
R1579 B.n440 B.n439 71.676
R1580 B.n433 B.n329 71.676
R1581 B.n432 B.n431 71.676
R1582 B.n425 B.n331 71.676
R1583 B.n424 B.n423 71.676
R1584 B.n417 B.n333 71.676
R1585 B.n416 B.n415 71.676
R1586 B.n409 B.n335 71.676
R1587 B.n408 B.n407 71.676
R1588 B.n401 B.n337 71.676
R1589 B.n400 B.n399 71.676
R1590 B.n393 B.n339 71.676
R1591 B.n392 B.n391 71.676
R1592 B.n385 B.n341 71.676
R1593 B.n384 B.n383 71.676
R1594 B.n377 B.n343 71.676
R1595 B.n376 B.n375 71.676
R1596 B.n369 B.n345 71.676
R1597 B.n368 B.n367 71.676
R1598 B.n361 B.n347 71.676
R1599 B.n360 B.n359 71.676
R1600 B.n353 B.n349 71.676
R1601 B.n352 B.n351 71.676
R1602 B.n617 B.n616 71.676
R1603 B.n611 B.n281 71.676
R1604 B.n609 B.n608 71.676
R1605 B.n604 B.n603 71.676
R1606 B.n601 B.n600 71.676
R1607 B.n596 B.n595 71.676
R1608 B.n593 B.n592 71.676
R1609 B.n588 B.n587 71.676
R1610 B.n585 B.n584 71.676
R1611 B.n580 B.n579 71.676
R1612 B.n577 B.n576 71.676
R1613 B.n572 B.n571 71.676
R1614 B.n569 B.n568 71.676
R1615 B.n564 B.n563 71.676
R1616 B.n561 B.n560 71.676
R1617 B.n556 B.n555 71.676
R1618 B.n553 B.n552 71.676
R1619 B.n548 B.n547 71.676
R1620 B.n545 B.n544 71.676
R1621 B.n540 B.n539 71.676
R1622 B.n537 B.n536 71.676
R1623 B.n532 B.n531 71.676
R1624 B.n529 B.n528 71.676
R1625 B.n524 B.n523 71.676
R1626 B.n521 B.n520 71.676
R1627 B.n516 B.n515 71.676
R1628 B.n513 B.n512 71.676
R1629 B.n508 B.n507 71.676
R1630 B.n505 B.n504 71.676
R1631 B.n500 B.n499 71.676
R1632 B.n497 B.n496 71.676
R1633 B.n491 B.n490 71.676
R1634 B.n488 B.n487 71.676
R1635 B.n483 B.n482 71.676
R1636 B.n480 B.n479 71.676
R1637 B.n474 B.n473 71.676
R1638 B.n471 B.n470 71.676
R1639 B.n466 B.n465 71.676
R1640 B.n463 B.n462 71.676
R1641 B.n458 B.n457 71.676
R1642 B.n455 B.n454 71.676
R1643 B.n450 B.n449 71.676
R1644 B.n447 B.n446 71.676
R1645 B.n442 B.n441 71.676
R1646 B.n439 B.n438 71.676
R1647 B.n434 B.n433 71.676
R1648 B.n431 B.n430 71.676
R1649 B.n426 B.n425 71.676
R1650 B.n423 B.n422 71.676
R1651 B.n418 B.n417 71.676
R1652 B.n415 B.n414 71.676
R1653 B.n410 B.n409 71.676
R1654 B.n407 B.n406 71.676
R1655 B.n402 B.n401 71.676
R1656 B.n399 B.n398 71.676
R1657 B.n394 B.n393 71.676
R1658 B.n391 B.n390 71.676
R1659 B.n386 B.n385 71.676
R1660 B.n383 B.n382 71.676
R1661 B.n378 B.n377 71.676
R1662 B.n375 B.n374 71.676
R1663 B.n370 B.n369 71.676
R1664 B.n367 B.n366 71.676
R1665 B.n362 B.n361 71.676
R1666 B.n359 B.n358 71.676
R1667 B.n354 B.n353 71.676
R1668 B.n351 B.n277 71.676
R1669 B.n1236 B.n1235 71.676
R1670 B.n1236 B.n2 71.676
R1671 B.n142 B.t20 69.7045
R1672 B.n319 B.t12 69.7045
R1673 B.n135 B.t23 69.6787
R1674 B.n313 B.t15 69.6787
R1675 B.n136 B.n135 59.5399
R1676 B.n980 B.n142 59.5399
R1677 B.n476 B.n319 59.5399
R1678 B.n494 B.n313 59.5399
R1679 B.n622 B.n278 50.8493
R1680 B.n1127 B.n100 50.8493
R1681 B.n135 B.n134 50.8126
R1682 B.n142 B.n141 50.8126
R1683 B.n319 B.n318 50.8126
R1684 B.n313 B.n312 50.8126
R1685 B.n620 B.n619 30.7517
R1686 B.n624 B.n276 30.7517
R1687 B.n854 B.n853 30.7517
R1688 B.n1125 B.n1124 30.7517
R1689 B.n622 B.n274 30.5998
R1690 B.n628 B.n274 30.5998
R1691 B.n628 B.n270 30.5998
R1692 B.n634 B.n270 30.5998
R1693 B.n634 B.n266 30.5998
R1694 B.n641 B.n266 30.5998
R1695 B.n641 B.n640 30.5998
R1696 B.n647 B.n259 30.5998
R1697 B.n653 B.n259 30.5998
R1698 B.n653 B.n255 30.5998
R1699 B.n659 B.n255 30.5998
R1700 B.n659 B.n251 30.5998
R1701 B.n665 B.n251 30.5998
R1702 B.n665 B.n247 30.5998
R1703 B.n671 B.n247 30.5998
R1704 B.n671 B.n243 30.5998
R1705 B.n677 B.n243 30.5998
R1706 B.n683 B.n239 30.5998
R1707 B.n683 B.n235 30.5998
R1708 B.n689 B.n235 30.5998
R1709 B.n689 B.n230 30.5998
R1710 B.n695 B.n230 30.5998
R1711 B.n695 B.n231 30.5998
R1712 B.n701 B.n223 30.5998
R1713 B.n707 B.n223 30.5998
R1714 B.n707 B.n219 30.5998
R1715 B.n713 B.n219 30.5998
R1716 B.n713 B.n214 30.5998
R1717 B.n719 B.n214 30.5998
R1718 B.n719 B.n215 30.5998
R1719 B.n725 B.n207 30.5998
R1720 B.n731 B.n207 30.5998
R1721 B.n731 B.n203 30.5998
R1722 B.n737 B.n203 30.5998
R1723 B.n737 B.n198 30.5998
R1724 B.n743 B.n198 30.5998
R1725 B.n743 B.n199 30.5998
R1726 B.n749 B.n191 30.5998
R1727 B.n755 B.n191 30.5998
R1728 B.n755 B.n187 30.5998
R1729 B.n761 B.n187 30.5998
R1730 B.n761 B.n182 30.5998
R1731 B.n767 B.n182 30.5998
R1732 B.n767 B.n183 30.5998
R1733 B.n774 B.n175 30.5998
R1734 B.n780 B.n175 30.5998
R1735 B.n780 B.n4 30.5998
R1736 B.n1234 B.n4 30.5998
R1737 B.n1234 B.n1233 30.5998
R1738 B.n1233 B.n1232 30.5998
R1739 B.n1232 B.n8 30.5998
R1740 B.n12 B.n8 30.5998
R1741 B.n1225 B.n12 30.5998
R1742 B.n1224 B.n1223 30.5998
R1743 B.n1223 B.n16 30.5998
R1744 B.n1217 B.n16 30.5998
R1745 B.n1217 B.n1216 30.5998
R1746 B.n1216 B.n1215 30.5998
R1747 B.n1215 B.n23 30.5998
R1748 B.n1209 B.n23 30.5998
R1749 B.n1208 B.n1207 30.5998
R1750 B.n1207 B.n30 30.5998
R1751 B.n1201 B.n30 30.5998
R1752 B.n1201 B.n1200 30.5998
R1753 B.n1200 B.n1199 30.5998
R1754 B.n1199 B.n37 30.5998
R1755 B.n1193 B.n37 30.5998
R1756 B.n1192 B.n1191 30.5998
R1757 B.n1191 B.n44 30.5998
R1758 B.n1185 B.n44 30.5998
R1759 B.n1185 B.n1184 30.5998
R1760 B.n1184 B.n1183 30.5998
R1761 B.n1183 B.n51 30.5998
R1762 B.n1177 B.n51 30.5998
R1763 B.n1176 B.n1175 30.5998
R1764 B.n1175 B.n58 30.5998
R1765 B.n1169 B.n58 30.5998
R1766 B.n1169 B.n1168 30.5998
R1767 B.n1168 B.n1167 30.5998
R1768 B.n1167 B.n65 30.5998
R1769 B.n1161 B.n1160 30.5998
R1770 B.n1160 B.n1159 30.5998
R1771 B.n1159 B.n72 30.5998
R1772 B.n1153 B.n72 30.5998
R1773 B.n1153 B.n1152 30.5998
R1774 B.n1152 B.n1151 30.5998
R1775 B.n1151 B.n79 30.5998
R1776 B.n1145 B.n79 30.5998
R1777 B.n1145 B.n1144 30.5998
R1778 B.n1144 B.n1143 30.5998
R1779 B.n1137 B.n89 30.5998
R1780 B.n1137 B.n1136 30.5998
R1781 B.n1136 B.n1135 30.5998
R1782 B.n1135 B.n93 30.5998
R1783 B.n1129 B.n93 30.5998
R1784 B.n1129 B.n1128 30.5998
R1785 B.n1128 B.n1127 30.5998
R1786 B.n774 B.t1 29.2498
R1787 B.n1225 B.t4 29.2498
R1788 B.n231 B.t9 28.3499
R1789 B.t0 B.n1176 28.3499
R1790 B.t3 B.n239 23.85
R1791 B.t2 B.n65 23.85
R1792 B.n647 B.t11 21.15
R1793 B.n1143 B.t18 21.15
R1794 B.n749 B.t6 20.25
R1795 B.n1209 B.t5 20.25
R1796 B.n215 B.t8 19.3501
R1797 B.t7 B.n1192 19.3501
R1798 B B.n1237 18.0485
R1799 B.n725 B.t8 11.2502
R1800 B.n1193 B.t7 11.2502
R1801 B.n620 B.n272 10.6151
R1802 B.n630 B.n272 10.6151
R1803 B.n631 B.n630 10.6151
R1804 B.n632 B.n631 10.6151
R1805 B.n632 B.n264 10.6151
R1806 B.n643 B.n264 10.6151
R1807 B.n644 B.n643 10.6151
R1808 B.n645 B.n644 10.6151
R1809 B.n645 B.n257 10.6151
R1810 B.n655 B.n257 10.6151
R1811 B.n656 B.n655 10.6151
R1812 B.n657 B.n656 10.6151
R1813 B.n657 B.n249 10.6151
R1814 B.n667 B.n249 10.6151
R1815 B.n668 B.n667 10.6151
R1816 B.n669 B.n668 10.6151
R1817 B.n669 B.n241 10.6151
R1818 B.n679 B.n241 10.6151
R1819 B.n680 B.n679 10.6151
R1820 B.n681 B.n680 10.6151
R1821 B.n681 B.n233 10.6151
R1822 B.n691 B.n233 10.6151
R1823 B.n692 B.n691 10.6151
R1824 B.n693 B.n692 10.6151
R1825 B.n693 B.n225 10.6151
R1826 B.n703 B.n225 10.6151
R1827 B.n704 B.n703 10.6151
R1828 B.n705 B.n704 10.6151
R1829 B.n705 B.n217 10.6151
R1830 B.n715 B.n217 10.6151
R1831 B.n716 B.n715 10.6151
R1832 B.n717 B.n716 10.6151
R1833 B.n717 B.n209 10.6151
R1834 B.n727 B.n209 10.6151
R1835 B.n728 B.n727 10.6151
R1836 B.n729 B.n728 10.6151
R1837 B.n729 B.n201 10.6151
R1838 B.n739 B.n201 10.6151
R1839 B.n740 B.n739 10.6151
R1840 B.n741 B.n740 10.6151
R1841 B.n741 B.n193 10.6151
R1842 B.n751 B.n193 10.6151
R1843 B.n752 B.n751 10.6151
R1844 B.n753 B.n752 10.6151
R1845 B.n753 B.n185 10.6151
R1846 B.n763 B.n185 10.6151
R1847 B.n764 B.n763 10.6151
R1848 B.n765 B.n764 10.6151
R1849 B.n765 B.n177 10.6151
R1850 B.n776 B.n177 10.6151
R1851 B.n777 B.n776 10.6151
R1852 B.n778 B.n777 10.6151
R1853 B.n778 B.n0 10.6151
R1854 B.n619 B.n618 10.6151
R1855 B.n618 B.n280 10.6151
R1856 B.n613 B.n280 10.6151
R1857 B.n613 B.n612 10.6151
R1858 B.n612 B.n282 10.6151
R1859 B.n607 B.n282 10.6151
R1860 B.n607 B.n606 10.6151
R1861 B.n606 B.n605 10.6151
R1862 B.n605 B.n284 10.6151
R1863 B.n599 B.n284 10.6151
R1864 B.n599 B.n598 10.6151
R1865 B.n598 B.n597 10.6151
R1866 B.n597 B.n286 10.6151
R1867 B.n591 B.n286 10.6151
R1868 B.n591 B.n590 10.6151
R1869 B.n590 B.n589 10.6151
R1870 B.n589 B.n288 10.6151
R1871 B.n583 B.n288 10.6151
R1872 B.n583 B.n582 10.6151
R1873 B.n582 B.n581 10.6151
R1874 B.n581 B.n290 10.6151
R1875 B.n575 B.n290 10.6151
R1876 B.n575 B.n574 10.6151
R1877 B.n574 B.n573 10.6151
R1878 B.n573 B.n292 10.6151
R1879 B.n567 B.n292 10.6151
R1880 B.n567 B.n566 10.6151
R1881 B.n566 B.n565 10.6151
R1882 B.n565 B.n294 10.6151
R1883 B.n559 B.n294 10.6151
R1884 B.n559 B.n558 10.6151
R1885 B.n558 B.n557 10.6151
R1886 B.n557 B.n296 10.6151
R1887 B.n551 B.n296 10.6151
R1888 B.n551 B.n550 10.6151
R1889 B.n550 B.n549 10.6151
R1890 B.n549 B.n298 10.6151
R1891 B.n543 B.n298 10.6151
R1892 B.n543 B.n542 10.6151
R1893 B.n542 B.n541 10.6151
R1894 B.n541 B.n300 10.6151
R1895 B.n535 B.n300 10.6151
R1896 B.n535 B.n534 10.6151
R1897 B.n534 B.n533 10.6151
R1898 B.n533 B.n302 10.6151
R1899 B.n527 B.n302 10.6151
R1900 B.n527 B.n526 10.6151
R1901 B.n526 B.n525 10.6151
R1902 B.n525 B.n304 10.6151
R1903 B.n519 B.n304 10.6151
R1904 B.n519 B.n518 10.6151
R1905 B.n518 B.n517 10.6151
R1906 B.n517 B.n306 10.6151
R1907 B.n511 B.n306 10.6151
R1908 B.n511 B.n510 10.6151
R1909 B.n510 B.n509 10.6151
R1910 B.n509 B.n308 10.6151
R1911 B.n503 B.n308 10.6151
R1912 B.n503 B.n502 10.6151
R1913 B.n502 B.n501 10.6151
R1914 B.n501 B.n310 10.6151
R1915 B.n495 B.n310 10.6151
R1916 B.n493 B.n492 10.6151
R1917 B.n492 B.n314 10.6151
R1918 B.n486 B.n314 10.6151
R1919 B.n486 B.n485 10.6151
R1920 B.n485 B.n484 10.6151
R1921 B.n484 B.n316 10.6151
R1922 B.n478 B.n316 10.6151
R1923 B.n478 B.n477 10.6151
R1924 B.n475 B.n320 10.6151
R1925 B.n469 B.n320 10.6151
R1926 B.n469 B.n468 10.6151
R1927 B.n468 B.n467 10.6151
R1928 B.n467 B.n322 10.6151
R1929 B.n461 B.n322 10.6151
R1930 B.n461 B.n460 10.6151
R1931 B.n460 B.n459 10.6151
R1932 B.n459 B.n324 10.6151
R1933 B.n453 B.n324 10.6151
R1934 B.n453 B.n452 10.6151
R1935 B.n452 B.n451 10.6151
R1936 B.n451 B.n326 10.6151
R1937 B.n445 B.n326 10.6151
R1938 B.n445 B.n444 10.6151
R1939 B.n444 B.n443 10.6151
R1940 B.n443 B.n328 10.6151
R1941 B.n437 B.n328 10.6151
R1942 B.n437 B.n436 10.6151
R1943 B.n436 B.n435 10.6151
R1944 B.n435 B.n330 10.6151
R1945 B.n429 B.n330 10.6151
R1946 B.n429 B.n428 10.6151
R1947 B.n428 B.n427 10.6151
R1948 B.n427 B.n332 10.6151
R1949 B.n421 B.n332 10.6151
R1950 B.n421 B.n420 10.6151
R1951 B.n420 B.n419 10.6151
R1952 B.n419 B.n334 10.6151
R1953 B.n413 B.n334 10.6151
R1954 B.n413 B.n412 10.6151
R1955 B.n412 B.n411 10.6151
R1956 B.n411 B.n336 10.6151
R1957 B.n405 B.n336 10.6151
R1958 B.n405 B.n404 10.6151
R1959 B.n404 B.n403 10.6151
R1960 B.n403 B.n338 10.6151
R1961 B.n397 B.n338 10.6151
R1962 B.n397 B.n396 10.6151
R1963 B.n396 B.n395 10.6151
R1964 B.n395 B.n340 10.6151
R1965 B.n389 B.n340 10.6151
R1966 B.n389 B.n388 10.6151
R1967 B.n388 B.n387 10.6151
R1968 B.n387 B.n342 10.6151
R1969 B.n381 B.n342 10.6151
R1970 B.n381 B.n380 10.6151
R1971 B.n380 B.n379 10.6151
R1972 B.n379 B.n344 10.6151
R1973 B.n373 B.n344 10.6151
R1974 B.n373 B.n372 10.6151
R1975 B.n372 B.n371 10.6151
R1976 B.n371 B.n346 10.6151
R1977 B.n365 B.n346 10.6151
R1978 B.n365 B.n364 10.6151
R1979 B.n364 B.n363 10.6151
R1980 B.n363 B.n348 10.6151
R1981 B.n357 B.n348 10.6151
R1982 B.n357 B.n356 10.6151
R1983 B.n356 B.n355 10.6151
R1984 B.n355 B.n350 10.6151
R1985 B.n350 B.n276 10.6151
R1986 B.n625 B.n624 10.6151
R1987 B.n626 B.n625 10.6151
R1988 B.n626 B.n268 10.6151
R1989 B.n636 B.n268 10.6151
R1990 B.n637 B.n636 10.6151
R1991 B.n638 B.n637 10.6151
R1992 B.n638 B.n261 10.6151
R1993 B.n649 B.n261 10.6151
R1994 B.n650 B.n649 10.6151
R1995 B.n651 B.n650 10.6151
R1996 B.n651 B.n253 10.6151
R1997 B.n661 B.n253 10.6151
R1998 B.n662 B.n661 10.6151
R1999 B.n663 B.n662 10.6151
R2000 B.n663 B.n245 10.6151
R2001 B.n673 B.n245 10.6151
R2002 B.n674 B.n673 10.6151
R2003 B.n675 B.n674 10.6151
R2004 B.n675 B.n237 10.6151
R2005 B.n685 B.n237 10.6151
R2006 B.n686 B.n685 10.6151
R2007 B.n687 B.n686 10.6151
R2008 B.n687 B.n228 10.6151
R2009 B.n697 B.n228 10.6151
R2010 B.n698 B.n697 10.6151
R2011 B.n699 B.n698 10.6151
R2012 B.n699 B.n221 10.6151
R2013 B.n709 B.n221 10.6151
R2014 B.n710 B.n709 10.6151
R2015 B.n711 B.n710 10.6151
R2016 B.n711 B.n212 10.6151
R2017 B.n721 B.n212 10.6151
R2018 B.n722 B.n721 10.6151
R2019 B.n723 B.n722 10.6151
R2020 B.n723 B.n205 10.6151
R2021 B.n733 B.n205 10.6151
R2022 B.n734 B.n733 10.6151
R2023 B.n735 B.n734 10.6151
R2024 B.n735 B.n196 10.6151
R2025 B.n745 B.n196 10.6151
R2026 B.n746 B.n745 10.6151
R2027 B.n747 B.n746 10.6151
R2028 B.n747 B.n189 10.6151
R2029 B.n757 B.n189 10.6151
R2030 B.n758 B.n757 10.6151
R2031 B.n759 B.n758 10.6151
R2032 B.n759 B.n180 10.6151
R2033 B.n769 B.n180 10.6151
R2034 B.n770 B.n769 10.6151
R2035 B.n772 B.n770 10.6151
R2036 B.n772 B.n771 10.6151
R2037 B.n771 B.n173 10.6151
R2038 B.n783 B.n173 10.6151
R2039 B.n784 B.n783 10.6151
R2040 B.n785 B.n784 10.6151
R2041 B.n786 B.n785 10.6151
R2042 B.n787 B.n786 10.6151
R2043 B.n790 B.n787 10.6151
R2044 B.n791 B.n790 10.6151
R2045 B.n792 B.n791 10.6151
R2046 B.n793 B.n792 10.6151
R2047 B.n795 B.n793 10.6151
R2048 B.n796 B.n795 10.6151
R2049 B.n797 B.n796 10.6151
R2050 B.n798 B.n797 10.6151
R2051 B.n800 B.n798 10.6151
R2052 B.n801 B.n800 10.6151
R2053 B.n802 B.n801 10.6151
R2054 B.n803 B.n802 10.6151
R2055 B.n805 B.n803 10.6151
R2056 B.n806 B.n805 10.6151
R2057 B.n807 B.n806 10.6151
R2058 B.n808 B.n807 10.6151
R2059 B.n810 B.n808 10.6151
R2060 B.n811 B.n810 10.6151
R2061 B.n812 B.n811 10.6151
R2062 B.n813 B.n812 10.6151
R2063 B.n815 B.n813 10.6151
R2064 B.n816 B.n815 10.6151
R2065 B.n817 B.n816 10.6151
R2066 B.n818 B.n817 10.6151
R2067 B.n820 B.n818 10.6151
R2068 B.n821 B.n820 10.6151
R2069 B.n822 B.n821 10.6151
R2070 B.n823 B.n822 10.6151
R2071 B.n825 B.n823 10.6151
R2072 B.n826 B.n825 10.6151
R2073 B.n827 B.n826 10.6151
R2074 B.n828 B.n827 10.6151
R2075 B.n830 B.n828 10.6151
R2076 B.n831 B.n830 10.6151
R2077 B.n832 B.n831 10.6151
R2078 B.n833 B.n832 10.6151
R2079 B.n835 B.n833 10.6151
R2080 B.n836 B.n835 10.6151
R2081 B.n837 B.n836 10.6151
R2082 B.n838 B.n837 10.6151
R2083 B.n840 B.n838 10.6151
R2084 B.n841 B.n840 10.6151
R2085 B.n842 B.n841 10.6151
R2086 B.n843 B.n842 10.6151
R2087 B.n845 B.n843 10.6151
R2088 B.n846 B.n845 10.6151
R2089 B.n847 B.n846 10.6151
R2090 B.n848 B.n847 10.6151
R2091 B.n850 B.n848 10.6151
R2092 B.n851 B.n850 10.6151
R2093 B.n852 B.n851 10.6151
R2094 B.n853 B.n852 10.6151
R2095 B.n1229 B.n1 10.6151
R2096 B.n1229 B.n1228 10.6151
R2097 B.n1228 B.n1227 10.6151
R2098 B.n1227 B.n10 10.6151
R2099 B.n1221 B.n10 10.6151
R2100 B.n1221 B.n1220 10.6151
R2101 B.n1220 B.n1219 10.6151
R2102 B.n1219 B.n18 10.6151
R2103 B.n1213 B.n18 10.6151
R2104 B.n1213 B.n1212 10.6151
R2105 B.n1212 B.n1211 10.6151
R2106 B.n1211 B.n25 10.6151
R2107 B.n1205 B.n25 10.6151
R2108 B.n1205 B.n1204 10.6151
R2109 B.n1204 B.n1203 10.6151
R2110 B.n1203 B.n32 10.6151
R2111 B.n1197 B.n32 10.6151
R2112 B.n1197 B.n1196 10.6151
R2113 B.n1196 B.n1195 10.6151
R2114 B.n1195 B.n39 10.6151
R2115 B.n1189 B.n39 10.6151
R2116 B.n1189 B.n1188 10.6151
R2117 B.n1188 B.n1187 10.6151
R2118 B.n1187 B.n46 10.6151
R2119 B.n1181 B.n46 10.6151
R2120 B.n1181 B.n1180 10.6151
R2121 B.n1180 B.n1179 10.6151
R2122 B.n1179 B.n53 10.6151
R2123 B.n1173 B.n53 10.6151
R2124 B.n1173 B.n1172 10.6151
R2125 B.n1172 B.n1171 10.6151
R2126 B.n1171 B.n60 10.6151
R2127 B.n1165 B.n60 10.6151
R2128 B.n1165 B.n1164 10.6151
R2129 B.n1164 B.n1163 10.6151
R2130 B.n1163 B.n67 10.6151
R2131 B.n1157 B.n67 10.6151
R2132 B.n1157 B.n1156 10.6151
R2133 B.n1156 B.n1155 10.6151
R2134 B.n1155 B.n74 10.6151
R2135 B.n1149 B.n74 10.6151
R2136 B.n1149 B.n1148 10.6151
R2137 B.n1148 B.n1147 10.6151
R2138 B.n1147 B.n81 10.6151
R2139 B.n1141 B.n81 10.6151
R2140 B.n1141 B.n1140 10.6151
R2141 B.n1140 B.n1139 10.6151
R2142 B.n1139 B.n87 10.6151
R2143 B.n1133 B.n87 10.6151
R2144 B.n1133 B.n1132 10.6151
R2145 B.n1132 B.n1131 10.6151
R2146 B.n1131 B.n95 10.6151
R2147 B.n1125 B.n95 10.6151
R2148 B.n1124 B.n1123 10.6151
R2149 B.n1123 B.n102 10.6151
R2150 B.n1117 B.n102 10.6151
R2151 B.n1117 B.n1116 10.6151
R2152 B.n1116 B.n1115 10.6151
R2153 B.n1115 B.n104 10.6151
R2154 B.n1109 B.n104 10.6151
R2155 B.n1109 B.n1108 10.6151
R2156 B.n1108 B.n1107 10.6151
R2157 B.n1107 B.n106 10.6151
R2158 B.n1101 B.n106 10.6151
R2159 B.n1101 B.n1100 10.6151
R2160 B.n1100 B.n1099 10.6151
R2161 B.n1099 B.n108 10.6151
R2162 B.n1093 B.n108 10.6151
R2163 B.n1093 B.n1092 10.6151
R2164 B.n1092 B.n1091 10.6151
R2165 B.n1091 B.n110 10.6151
R2166 B.n1085 B.n110 10.6151
R2167 B.n1085 B.n1084 10.6151
R2168 B.n1084 B.n1083 10.6151
R2169 B.n1083 B.n112 10.6151
R2170 B.n1077 B.n112 10.6151
R2171 B.n1077 B.n1076 10.6151
R2172 B.n1076 B.n1075 10.6151
R2173 B.n1075 B.n114 10.6151
R2174 B.n1069 B.n114 10.6151
R2175 B.n1069 B.n1068 10.6151
R2176 B.n1068 B.n1067 10.6151
R2177 B.n1067 B.n116 10.6151
R2178 B.n1061 B.n116 10.6151
R2179 B.n1061 B.n1060 10.6151
R2180 B.n1060 B.n1059 10.6151
R2181 B.n1059 B.n118 10.6151
R2182 B.n1053 B.n118 10.6151
R2183 B.n1053 B.n1052 10.6151
R2184 B.n1052 B.n1051 10.6151
R2185 B.n1051 B.n120 10.6151
R2186 B.n1045 B.n120 10.6151
R2187 B.n1045 B.n1044 10.6151
R2188 B.n1044 B.n1043 10.6151
R2189 B.n1043 B.n122 10.6151
R2190 B.n1037 B.n122 10.6151
R2191 B.n1037 B.n1036 10.6151
R2192 B.n1036 B.n1035 10.6151
R2193 B.n1035 B.n124 10.6151
R2194 B.n1029 B.n124 10.6151
R2195 B.n1029 B.n1028 10.6151
R2196 B.n1028 B.n1027 10.6151
R2197 B.n1027 B.n126 10.6151
R2198 B.n1021 B.n126 10.6151
R2199 B.n1021 B.n1020 10.6151
R2200 B.n1020 B.n1019 10.6151
R2201 B.n1019 B.n128 10.6151
R2202 B.n1013 B.n128 10.6151
R2203 B.n1013 B.n1012 10.6151
R2204 B.n1012 B.n1011 10.6151
R2205 B.n1011 B.n130 10.6151
R2206 B.n1005 B.n130 10.6151
R2207 B.n1005 B.n1004 10.6151
R2208 B.n1004 B.n1003 10.6151
R2209 B.n1003 B.n132 10.6151
R2210 B.n997 B.n996 10.6151
R2211 B.n996 B.n995 10.6151
R2212 B.n995 B.n137 10.6151
R2213 B.n989 B.n137 10.6151
R2214 B.n989 B.n988 10.6151
R2215 B.n988 B.n987 10.6151
R2216 B.n987 B.n139 10.6151
R2217 B.n981 B.n139 10.6151
R2218 B.n979 B.n978 10.6151
R2219 B.n978 B.n143 10.6151
R2220 B.n972 B.n143 10.6151
R2221 B.n972 B.n971 10.6151
R2222 B.n971 B.n970 10.6151
R2223 B.n970 B.n145 10.6151
R2224 B.n964 B.n145 10.6151
R2225 B.n964 B.n963 10.6151
R2226 B.n963 B.n962 10.6151
R2227 B.n962 B.n147 10.6151
R2228 B.n956 B.n147 10.6151
R2229 B.n956 B.n955 10.6151
R2230 B.n955 B.n954 10.6151
R2231 B.n954 B.n149 10.6151
R2232 B.n948 B.n149 10.6151
R2233 B.n948 B.n947 10.6151
R2234 B.n947 B.n946 10.6151
R2235 B.n946 B.n151 10.6151
R2236 B.n940 B.n151 10.6151
R2237 B.n940 B.n939 10.6151
R2238 B.n939 B.n938 10.6151
R2239 B.n938 B.n153 10.6151
R2240 B.n932 B.n153 10.6151
R2241 B.n932 B.n931 10.6151
R2242 B.n931 B.n930 10.6151
R2243 B.n930 B.n155 10.6151
R2244 B.n924 B.n155 10.6151
R2245 B.n924 B.n923 10.6151
R2246 B.n923 B.n922 10.6151
R2247 B.n922 B.n157 10.6151
R2248 B.n916 B.n157 10.6151
R2249 B.n916 B.n915 10.6151
R2250 B.n915 B.n914 10.6151
R2251 B.n914 B.n159 10.6151
R2252 B.n908 B.n159 10.6151
R2253 B.n908 B.n907 10.6151
R2254 B.n907 B.n906 10.6151
R2255 B.n906 B.n161 10.6151
R2256 B.n900 B.n161 10.6151
R2257 B.n900 B.n899 10.6151
R2258 B.n899 B.n898 10.6151
R2259 B.n898 B.n163 10.6151
R2260 B.n892 B.n163 10.6151
R2261 B.n892 B.n891 10.6151
R2262 B.n891 B.n890 10.6151
R2263 B.n890 B.n165 10.6151
R2264 B.n884 B.n165 10.6151
R2265 B.n884 B.n883 10.6151
R2266 B.n883 B.n882 10.6151
R2267 B.n882 B.n167 10.6151
R2268 B.n876 B.n167 10.6151
R2269 B.n876 B.n875 10.6151
R2270 B.n875 B.n874 10.6151
R2271 B.n874 B.n169 10.6151
R2272 B.n868 B.n169 10.6151
R2273 B.n868 B.n867 10.6151
R2274 B.n867 B.n866 10.6151
R2275 B.n866 B.n171 10.6151
R2276 B.n860 B.n171 10.6151
R2277 B.n860 B.n859 10.6151
R2278 B.n859 B.n858 10.6151
R2279 B.n858 B.n854 10.6151
R2280 B.n199 B.t6 10.3503
R2281 B.t5 B.n1208 10.3503
R2282 B.n640 B.t11 9.45029
R2283 B.n89 B.t18 9.45029
R2284 B.n1237 B.n0 8.11757
R2285 B.n1237 B.n1 8.11757
R2286 B.n677 B.t3 6.75035
R2287 B.n1161 B.t2 6.75035
R2288 B.n494 B.n493 6.5566
R2289 B.n477 B.n476 6.5566
R2290 B.n997 B.n136 6.5566
R2291 B.n981 B.n980 6.5566
R2292 B.n495 B.n494 4.05904
R2293 B.n476 B.n475 4.05904
R2294 B.n136 B.n132 4.05904
R2295 B.n980 B.n979 4.05904
R2296 B.n701 B.t9 2.25045
R2297 B.n1177 B.t0 2.25045
R2298 B.n183 B.t1 1.35047
R2299 B.t4 B.n1224 1.35047
R2300 VN.n8 VN.t5 233.322
R2301 VN.n45 VN.t8 233.322
R2302 VN.n5 VN.t2 201.745
R2303 VN.n9 VN.t4 201.745
R2304 VN.n27 VN.t9 201.745
R2305 VN.n35 VN.t7 201.745
R2306 VN.n42 VN.t1 201.745
R2307 VN.n46 VN.t3 201.745
R2308 VN.n64 VN.t0 201.745
R2309 VN.n72 VN.t6 201.745
R2310 VN.n71 VN.n37 161.3
R2311 VN.n70 VN.n69 161.3
R2312 VN.n68 VN.n38 161.3
R2313 VN.n67 VN.n66 161.3
R2314 VN.n65 VN.n39 161.3
R2315 VN.n63 VN.n62 161.3
R2316 VN.n61 VN.n40 161.3
R2317 VN.n60 VN.n59 161.3
R2318 VN.n58 VN.n41 161.3
R2319 VN.n57 VN.n56 161.3
R2320 VN.n55 VN.n42 161.3
R2321 VN.n54 VN.n53 161.3
R2322 VN.n52 VN.n43 161.3
R2323 VN.n51 VN.n50 161.3
R2324 VN.n49 VN.n44 161.3
R2325 VN.n48 VN.n47 161.3
R2326 VN.n34 VN.n0 161.3
R2327 VN.n33 VN.n32 161.3
R2328 VN.n31 VN.n1 161.3
R2329 VN.n30 VN.n29 161.3
R2330 VN.n28 VN.n2 161.3
R2331 VN.n26 VN.n25 161.3
R2332 VN.n24 VN.n3 161.3
R2333 VN.n23 VN.n22 161.3
R2334 VN.n21 VN.n4 161.3
R2335 VN.n20 VN.n19 161.3
R2336 VN.n18 VN.n5 161.3
R2337 VN.n17 VN.n16 161.3
R2338 VN.n15 VN.n6 161.3
R2339 VN.n14 VN.n13 161.3
R2340 VN.n12 VN.n7 161.3
R2341 VN.n11 VN.n10 161.3
R2342 VN.n36 VN.n35 99.0123
R2343 VN.n73 VN.n72 99.0123
R2344 VN.n9 VN.n8 66.166
R2345 VN.n46 VN.n45 66.166
R2346 VN VN.n73 57.1118
R2347 VN.n15 VN.n14 56.5193
R2348 VN.n22 VN.n21 56.5193
R2349 VN.n52 VN.n51 56.5193
R2350 VN.n59 VN.n58 56.5193
R2351 VN.n29 VN.n1 47.2923
R2352 VN.n66 VN.n38 47.2923
R2353 VN.n33 VN.n1 33.6945
R2354 VN.n70 VN.n38 33.6945
R2355 VN.n10 VN.n7 24.4675
R2356 VN.n14 VN.n7 24.4675
R2357 VN.n16 VN.n15 24.4675
R2358 VN.n16 VN.n5 24.4675
R2359 VN.n20 VN.n5 24.4675
R2360 VN.n21 VN.n20 24.4675
R2361 VN.n22 VN.n3 24.4675
R2362 VN.n26 VN.n3 24.4675
R2363 VN.n29 VN.n28 24.4675
R2364 VN.n34 VN.n33 24.4675
R2365 VN.n51 VN.n44 24.4675
R2366 VN.n47 VN.n44 24.4675
R2367 VN.n58 VN.n57 24.4675
R2368 VN.n57 VN.n42 24.4675
R2369 VN.n53 VN.n42 24.4675
R2370 VN.n53 VN.n52 24.4675
R2371 VN.n66 VN.n65 24.4675
R2372 VN.n63 VN.n40 24.4675
R2373 VN.n59 VN.n40 24.4675
R2374 VN.n71 VN.n70 24.4675
R2375 VN.n28 VN.n27 18.5954
R2376 VN.n65 VN.n64 18.5954
R2377 VN.n35 VN.n34 11.7447
R2378 VN.n72 VN.n71 11.7447
R2379 VN.n48 VN.n45 9.81663
R2380 VN.n11 VN.n8 9.81663
R2381 VN.n10 VN.n9 5.87258
R2382 VN.n27 VN.n26 5.87258
R2383 VN.n47 VN.n46 5.87258
R2384 VN.n64 VN.n63 5.87258
R2385 VN.n73 VN.n37 0.278367
R2386 VN.n36 VN.n0 0.278367
R2387 VN.n69 VN.n37 0.189894
R2388 VN.n69 VN.n68 0.189894
R2389 VN.n68 VN.n67 0.189894
R2390 VN.n67 VN.n39 0.189894
R2391 VN.n62 VN.n39 0.189894
R2392 VN.n62 VN.n61 0.189894
R2393 VN.n61 VN.n60 0.189894
R2394 VN.n60 VN.n41 0.189894
R2395 VN.n56 VN.n41 0.189894
R2396 VN.n56 VN.n55 0.189894
R2397 VN.n55 VN.n54 0.189894
R2398 VN.n54 VN.n43 0.189894
R2399 VN.n50 VN.n43 0.189894
R2400 VN.n50 VN.n49 0.189894
R2401 VN.n49 VN.n48 0.189894
R2402 VN.n12 VN.n11 0.189894
R2403 VN.n13 VN.n12 0.189894
R2404 VN.n13 VN.n6 0.189894
R2405 VN.n17 VN.n6 0.189894
R2406 VN.n18 VN.n17 0.189894
R2407 VN.n19 VN.n18 0.189894
R2408 VN.n19 VN.n4 0.189894
R2409 VN.n23 VN.n4 0.189894
R2410 VN.n24 VN.n23 0.189894
R2411 VN.n25 VN.n24 0.189894
R2412 VN.n25 VN.n2 0.189894
R2413 VN.n30 VN.n2 0.189894
R2414 VN.n31 VN.n30 0.189894
R2415 VN.n32 VN.n31 0.189894
R2416 VN.n32 VN.n0 0.189894
R2417 VN VN.n36 0.153454
R2418 VDD2.n1 VDD2.t4 67.5636
R2419 VDD2.n3 VDD2.n2 65.9097
R2420 VDD2 VDD2.n7 65.9079
R2421 VDD2.n4 VDD2.t3 65.3051
R2422 VDD2.n6 VDD2.n5 64.2723
R2423 VDD2.n1 VDD2.n0 64.2711
R2424 VDD2.n4 VDD2.n3 50.9696
R2425 VDD2.n6 VDD2.n4 2.25912
R2426 VDD2.n7 VDD2.t6 1.03336
R2427 VDD2.n7 VDD2.t1 1.03336
R2428 VDD2.n5 VDD2.t9 1.03336
R2429 VDD2.n5 VDD2.t8 1.03336
R2430 VDD2.n2 VDD2.t0 1.03336
R2431 VDD2.n2 VDD2.t2 1.03336
R2432 VDD2.n0 VDD2.t5 1.03336
R2433 VDD2.n0 VDD2.t7 1.03336
R2434 VDD2 VDD2.n6 0.623345
R2435 VDD2.n3 VDD2.n1 0.509809
C0 VP VN 9.271791f
C1 VTAIL VP 16.5031f
C2 VDD2 VP 0.54465f
C3 VTAIL VN 16.488699f
C4 VDD2 VN 16.2883f
C5 VDD1 VP 16.675098f
C6 VDD2 VTAIL 13.944099f
C7 VDD1 VN 0.152628f
C8 VTAIL VDD1 13.8975f
C9 VDD2 VDD1 1.97347f
C10 VDD2 B 8.070951f
C11 VDD1 B 8.080392f
C12 VTAIL B 10.796312f
C13 VN B 17.30907f
C14 VP B 15.664197f
C15 VDD2.t4 B 3.89274f
C16 VDD2.t5 B 0.331219f
C17 VDD2.t7 B 0.331219f
C18 VDD2.n0 B 3.0331f
C19 VDD2.n1 B 0.75588f
C20 VDD2.t0 B 0.331219f
C21 VDD2.t2 B 0.331219f
C22 VDD2.n2 B 3.04448f
C23 VDD2.n3 B 2.78667f
C24 VDD2.t3 B 3.87941f
C25 VDD2.n4 B 3.0982f
C26 VDD2.t9 B 0.331219f
C27 VDD2.t8 B 0.331219f
C28 VDD2.n5 B 3.03311f
C29 VDD2.n6 B 0.377129f
C30 VDD2.t6 B 0.331219f
C31 VDD2.t1 B 0.331219f
C32 VDD2.n7 B 3.04444f
C33 VN.n0 B 0.029392f
C34 VN.t7 B 2.695f
C35 VN.n1 B 0.019466f
C36 VN.n2 B 0.022294f
C37 VN.t9 B 2.695f
C38 VN.n3 B 0.04155f
C39 VN.n4 B 0.022294f
C40 VN.t2 B 2.695f
C41 VN.n5 B 0.955779f
C42 VN.n6 B 0.022294f
C43 VN.n7 B 0.04155f
C44 VN.t5 B 2.83792f
C45 VN.n8 B 0.986274f
C46 VN.t4 B 2.695f
C47 VN.n9 B 0.989164f
C48 VN.n10 B 0.025959f
C49 VN.n11 B 0.191664f
C50 VN.n12 B 0.022294f
C51 VN.n13 B 0.022294f
C52 VN.n14 B 0.028817f
C53 VN.n15 B 0.036272f
C54 VN.n16 B 0.04155f
C55 VN.n17 B 0.022294f
C56 VN.n18 B 0.022294f
C57 VN.n19 B 0.022294f
C58 VN.n20 B 0.04155f
C59 VN.n21 B 0.036272f
C60 VN.n22 B 0.028817f
C61 VN.n23 B 0.022294f
C62 VN.n24 B 0.022294f
C63 VN.n25 B 0.022294f
C64 VN.n26 B 0.025959f
C65 VN.n27 B 0.934742f
C66 VN.n28 B 0.036626f
C67 VN.n29 B 0.042142f
C68 VN.n30 B 0.022294f
C69 VN.n31 B 0.022294f
C70 VN.n32 B 0.022294f
C71 VN.n33 B 0.045031f
C72 VN.n34 B 0.030883f
C73 VN.n35 B 1.0022f
C74 VN.n36 B 0.033234f
C75 VN.n37 B 0.029392f
C76 VN.t6 B 2.695f
C77 VN.n38 B 0.019466f
C78 VN.n39 B 0.022294f
C79 VN.t0 B 2.695f
C80 VN.n40 B 0.04155f
C81 VN.n41 B 0.022294f
C82 VN.t1 B 2.695f
C83 VN.n42 B 0.955779f
C84 VN.n43 B 0.022294f
C85 VN.n44 B 0.04155f
C86 VN.t8 B 2.83792f
C87 VN.n45 B 0.986274f
C88 VN.t3 B 2.695f
C89 VN.n46 B 0.989164f
C90 VN.n47 B 0.025959f
C91 VN.n48 B 0.191664f
C92 VN.n49 B 0.022294f
C93 VN.n50 B 0.022294f
C94 VN.n51 B 0.028817f
C95 VN.n52 B 0.036272f
C96 VN.n53 B 0.04155f
C97 VN.n54 B 0.022294f
C98 VN.n55 B 0.022294f
C99 VN.n56 B 0.022294f
C100 VN.n57 B 0.04155f
C101 VN.n58 B 0.036272f
C102 VN.n59 B 0.028817f
C103 VN.n60 B 0.022294f
C104 VN.n61 B 0.022294f
C105 VN.n62 B 0.022294f
C106 VN.n63 B 0.025959f
C107 VN.n64 B 0.934742f
C108 VN.n65 B 0.036626f
C109 VN.n66 B 0.042142f
C110 VN.n67 B 0.022294f
C111 VN.n68 B 0.022294f
C112 VN.n69 B 0.022294f
C113 VN.n70 B 0.045031f
C114 VN.n71 B 0.030883f
C115 VN.n72 B 1.0022f
C116 VN.n73 B 1.49737f
C117 VDD1.t1 B 3.9338f
C118 VDD1.t5 B 0.334711f
C119 VDD1.t9 B 0.334711f
C120 VDD1.n0 B 3.06508f
C121 VDD1.n1 B 0.770902f
C122 VDD1.t4 B 3.93378f
C123 VDD1.t0 B 0.334711f
C124 VDD1.t3 B 0.334711f
C125 VDD1.n2 B 3.06508f
C126 VDD1.n3 B 0.763849f
C127 VDD1.t8 B 0.334711f
C128 VDD1.t6 B 0.334711f
C129 VDD1.n4 B 3.07658f
C130 VDD1.n5 B 2.92271f
C131 VDD1.t2 B 0.334711f
C132 VDD1.t7 B 0.334711f
C133 VDD1.n6 B 3.06507f
C134 VDD1.n7 B 3.16467f
C135 VTAIL.t4 B 0.354298f
C136 VTAIL.t5 B 0.354298f
C137 VTAIL.n0 B 3.18073f
C138 VTAIL.n1 B 0.470746f
C139 VTAIL.t15 B 4.06642f
C140 VTAIL.n2 B 0.58949f
C141 VTAIL.t14 B 0.354298f
C142 VTAIL.t18 B 0.354298f
C143 VTAIL.n3 B 3.18073f
C144 VTAIL.n4 B 0.558613f
C145 VTAIL.t12 B 0.354298f
C146 VTAIL.t13 B 0.354298f
C147 VTAIL.n5 B 3.18073f
C148 VTAIL.n6 B 2.29193f
C149 VTAIL.t3 B 0.354298f
C150 VTAIL.t19 B 0.354298f
C151 VTAIL.n7 B 3.18074f
C152 VTAIL.n8 B 2.29192f
C153 VTAIL.t8 B 0.354298f
C154 VTAIL.t6 B 0.354298f
C155 VTAIL.n9 B 3.18074f
C156 VTAIL.n10 B 0.558604f
C157 VTAIL.t1 B 4.06645f
C158 VTAIL.n11 B 0.589461f
C159 VTAIL.t16 B 0.354298f
C160 VTAIL.t10 B 0.354298f
C161 VTAIL.n12 B 3.18074f
C162 VTAIL.n13 B 0.508905f
C163 VTAIL.t11 B 0.354298f
C164 VTAIL.t9 B 0.354298f
C165 VTAIL.n14 B 3.18074f
C166 VTAIL.n15 B 0.558604f
C167 VTAIL.t17 B 4.06642f
C168 VTAIL.n16 B 2.2023f
C169 VTAIL.t2 B 4.06642f
C170 VTAIL.n17 B 2.2023f
C171 VTAIL.t7 B 0.354298f
C172 VTAIL.t0 B 0.354298f
C173 VTAIL.n18 B 3.18073f
C174 VTAIL.n19 B 0.426568f
C175 VP.n0 B 0.029693f
C176 VP.t3 B 2.72263f
C177 VP.n1 B 0.019666f
C178 VP.n2 B 0.022522f
C179 VP.t1 B 2.72263f
C180 VP.n3 B 0.041975f
C181 VP.n4 B 0.022522f
C182 VP.t6 B 2.72263f
C183 VP.n5 B 0.965578f
C184 VP.n6 B 0.022522f
C185 VP.n7 B 0.041975f
C186 VP.n8 B 0.022522f
C187 VP.t9 B 2.72263f
C188 VP.n9 B 0.019666f
C189 VP.n10 B 0.029693f
C190 VP.t5 B 2.72263f
C191 VP.n11 B 0.029693f
C192 VP.t2 B 2.72263f
C193 VP.n12 B 0.019666f
C194 VP.n13 B 0.022522f
C195 VP.t7 B 2.72263f
C196 VP.n14 B 0.041975f
C197 VP.n15 B 0.022522f
C198 VP.t0 B 2.72263f
C199 VP.n16 B 0.965578f
C200 VP.n17 B 0.022522f
C201 VP.n18 B 0.041975f
C202 VP.t8 B 2.86701f
C203 VP.n19 B 0.996386f
C204 VP.t4 B 2.72263f
C205 VP.n20 B 0.999306f
C206 VP.n21 B 0.026226f
C207 VP.n22 B 0.19363f
C208 VP.n23 B 0.022522f
C209 VP.n24 B 0.022522f
C210 VP.n25 B 0.029112f
C211 VP.n26 B 0.036644f
C212 VP.n27 B 0.041975f
C213 VP.n28 B 0.022522f
C214 VP.n29 B 0.022522f
C215 VP.n30 B 0.022522f
C216 VP.n31 B 0.041975f
C217 VP.n32 B 0.036644f
C218 VP.n33 B 0.029112f
C219 VP.n34 B 0.022522f
C220 VP.n35 B 0.022522f
C221 VP.n36 B 0.022522f
C222 VP.n37 B 0.026226f
C223 VP.n38 B 0.944326f
C224 VP.n39 B 0.037002f
C225 VP.n40 B 0.042574f
C226 VP.n41 B 0.022522f
C227 VP.n42 B 0.022522f
C228 VP.n43 B 0.022522f
C229 VP.n44 B 0.045493f
C230 VP.n45 B 0.031199f
C231 VP.n46 B 1.01247f
C232 VP.n47 B 1.50085f
C233 VP.n48 B 1.51509f
C234 VP.n49 B 1.01247f
C235 VP.n50 B 0.031199f
C236 VP.n51 B 0.045493f
C237 VP.n52 B 0.022522f
C238 VP.n53 B 0.022522f
C239 VP.n54 B 0.022522f
C240 VP.n55 B 0.042574f
C241 VP.n56 B 0.037002f
C242 VP.n57 B 0.944326f
C243 VP.n58 B 0.026226f
C244 VP.n59 B 0.022522f
C245 VP.n60 B 0.022522f
C246 VP.n61 B 0.022522f
C247 VP.n62 B 0.029112f
C248 VP.n63 B 0.036644f
C249 VP.n64 B 0.041975f
C250 VP.n65 B 0.022522f
C251 VP.n66 B 0.022522f
C252 VP.n67 B 0.022522f
C253 VP.n68 B 0.041975f
C254 VP.n69 B 0.036644f
C255 VP.n70 B 0.029112f
C256 VP.n71 B 0.022522f
C257 VP.n72 B 0.022522f
C258 VP.n73 B 0.022522f
C259 VP.n74 B 0.026226f
C260 VP.n75 B 0.944326f
C261 VP.n76 B 0.037002f
C262 VP.n77 B 0.042574f
C263 VP.n78 B 0.022522f
C264 VP.n79 B 0.022522f
C265 VP.n80 B 0.022522f
C266 VP.n81 B 0.045493f
C267 VP.n82 B 0.031199f
C268 VP.n83 B 1.01247f
C269 VP.n84 B 0.033575f
.ends

