* NGSPICE file created from diff_pair_sample_0527.ext - technology: sky130A

.subckt diff_pair_sample_0527 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=1.21935 pd=7.72 as=2.8821 ps=15.56 w=7.39 l=1.75
X1 B.t11 B.t9 B.t10 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=0 ps=0 w=7.39 l=1.75
X2 B.t8 B.t6 B.t7 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=0 ps=0 w=7.39 l=1.75
X3 VTAIL.t0 VN.t0 VDD2.t3 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=1.21935 ps=7.72 w=7.39 l=1.75
X4 VDD2.t2 VN.t1 VTAIL.t2 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=1.21935 pd=7.72 as=2.8821 ps=15.56 w=7.39 l=1.75
X5 VTAIL.t5 VP.t1 VDD1.t2 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=1.21935 ps=7.72 w=7.39 l=1.75
X6 VTAIL.t1 VN.t2 VDD2.t1 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=1.21935 ps=7.72 w=7.39 l=1.75
X7 B.t5 B.t3 B.t4 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=0 ps=0 w=7.39 l=1.75
X8 B.t2 B.t0 B.t1 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=0 ps=0 w=7.39 l=1.75
X9 VDD1.t1 VP.t2 VTAIL.t6 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=1.21935 pd=7.72 as=2.8821 ps=15.56 w=7.39 l=1.75
X10 VDD2.t0 VN.t3 VTAIL.t3 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=1.21935 pd=7.72 as=2.8821 ps=15.56 w=7.39 l=1.75
X11 VTAIL.t7 VP.t3 VDD1.t0 w_n2218_n2446# sky130_fd_pr__pfet_01v8 ad=2.8821 pd=15.56 as=1.21935 ps=7.72 w=7.39 l=1.75
R0 VP.n5 VP.n4 183.81
R1 VP.n14 VP.n13 183.81
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n3 VP.t1 137.567
R8 VP.n3 VP.t0 137.142
R9 VP.n5 VP.t3 101.772
R10 VP.n13 VP.t2 101.772
R11 VP.n4 VP.n3 49.5251
R12 VP.n7 VP.n1 40.4934
R13 VP.n11 VP.n1 40.4934
R14 VP.n7 VP.n6 24.4675
R15 VP.n12 VP.n11 24.4675
R16 VP.n6 VP.n5 1.95786
R17 VP.n13 VP.n12 1.95786
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VTAIL.n314 VTAIL.n280 756.745
R26 VTAIL.n34 VTAIL.n0 756.745
R27 VTAIL.n74 VTAIL.n40 756.745
R28 VTAIL.n114 VTAIL.n80 756.745
R29 VTAIL.n274 VTAIL.n240 756.745
R30 VTAIL.n234 VTAIL.n200 756.745
R31 VTAIL.n194 VTAIL.n160 756.745
R32 VTAIL.n154 VTAIL.n120 756.745
R33 VTAIL.n292 VTAIL.n291 585
R34 VTAIL.n297 VTAIL.n296 585
R35 VTAIL.n299 VTAIL.n298 585
R36 VTAIL.n288 VTAIL.n287 585
R37 VTAIL.n305 VTAIL.n304 585
R38 VTAIL.n307 VTAIL.n306 585
R39 VTAIL.n284 VTAIL.n283 585
R40 VTAIL.n313 VTAIL.n312 585
R41 VTAIL.n315 VTAIL.n314 585
R42 VTAIL.n12 VTAIL.n11 585
R43 VTAIL.n17 VTAIL.n16 585
R44 VTAIL.n19 VTAIL.n18 585
R45 VTAIL.n8 VTAIL.n7 585
R46 VTAIL.n25 VTAIL.n24 585
R47 VTAIL.n27 VTAIL.n26 585
R48 VTAIL.n4 VTAIL.n3 585
R49 VTAIL.n33 VTAIL.n32 585
R50 VTAIL.n35 VTAIL.n34 585
R51 VTAIL.n52 VTAIL.n51 585
R52 VTAIL.n57 VTAIL.n56 585
R53 VTAIL.n59 VTAIL.n58 585
R54 VTAIL.n48 VTAIL.n47 585
R55 VTAIL.n65 VTAIL.n64 585
R56 VTAIL.n67 VTAIL.n66 585
R57 VTAIL.n44 VTAIL.n43 585
R58 VTAIL.n73 VTAIL.n72 585
R59 VTAIL.n75 VTAIL.n74 585
R60 VTAIL.n92 VTAIL.n91 585
R61 VTAIL.n97 VTAIL.n96 585
R62 VTAIL.n99 VTAIL.n98 585
R63 VTAIL.n88 VTAIL.n87 585
R64 VTAIL.n105 VTAIL.n104 585
R65 VTAIL.n107 VTAIL.n106 585
R66 VTAIL.n84 VTAIL.n83 585
R67 VTAIL.n113 VTAIL.n112 585
R68 VTAIL.n115 VTAIL.n114 585
R69 VTAIL.n275 VTAIL.n274 585
R70 VTAIL.n273 VTAIL.n272 585
R71 VTAIL.n244 VTAIL.n243 585
R72 VTAIL.n267 VTAIL.n266 585
R73 VTAIL.n265 VTAIL.n264 585
R74 VTAIL.n248 VTAIL.n247 585
R75 VTAIL.n259 VTAIL.n258 585
R76 VTAIL.n257 VTAIL.n256 585
R77 VTAIL.n252 VTAIL.n251 585
R78 VTAIL.n235 VTAIL.n234 585
R79 VTAIL.n233 VTAIL.n232 585
R80 VTAIL.n204 VTAIL.n203 585
R81 VTAIL.n227 VTAIL.n226 585
R82 VTAIL.n225 VTAIL.n224 585
R83 VTAIL.n208 VTAIL.n207 585
R84 VTAIL.n219 VTAIL.n218 585
R85 VTAIL.n217 VTAIL.n216 585
R86 VTAIL.n212 VTAIL.n211 585
R87 VTAIL.n195 VTAIL.n194 585
R88 VTAIL.n193 VTAIL.n192 585
R89 VTAIL.n164 VTAIL.n163 585
R90 VTAIL.n187 VTAIL.n186 585
R91 VTAIL.n185 VTAIL.n184 585
R92 VTAIL.n168 VTAIL.n167 585
R93 VTAIL.n179 VTAIL.n178 585
R94 VTAIL.n177 VTAIL.n176 585
R95 VTAIL.n172 VTAIL.n171 585
R96 VTAIL.n155 VTAIL.n154 585
R97 VTAIL.n153 VTAIL.n152 585
R98 VTAIL.n124 VTAIL.n123 585
R99 VTAIL.n147 VTAIL.n146 585
R100 VTAIL.n145 VTAIL.n144 585
R101 VTAIL.n128 VTAIL.n127 585
R102 VTAIL.n139 VTAIL.n138 585
R103 VTAIL.n137 VTAIL.n136 585
R104 VTAIL.n132 VTAIL.n131 585
R105 VTAIL.n293 VTAIL.t2 327.483
R106 VTAIL.n13 VTAIL.t1 327.483
R107 VTAIL.n53 VTAIL.t6 327.483
R108 VTAIL.n93 VTAIL.t7 327.483
R109 VTAIL.n253 VTAIL.t4 327.483
R110 VTAIL.n213 VTAIL.t5 327.483
R111 VTAIL.n173 VTAIL.t3 327.483
R112 VTAIL.n133 VTAIL.t0 327.483
R113 VTAIL.n297 VTAIL.n291 171.744
R114 VTAIL.n298 VTAIL.n297 171.744
R115 VTAIL.n298 VTAIL.n287 171.744
R116 VTAIL.n305 VTAIL.n287 171.744
R117 VTAIL.n306 VTAIL.n305 171.744
R118 VTAIL.n306 VTAIL.n283 171.744
R119 VTAIL.n313 VTAIL.n283 171.744
R120 VTAIL.n314 VTAIL.n313 171.744
R121 VTAIL.n17 VTAIL.n11 171.744
R122 VTAIL.n18 VTAIL.n17 171.744
R123 VTAIL.n18 VTAIL.n7 171.744
R124 VTAIL.n25 VTAIL.n7 171.744
R125 VTAIL.n26 VTAIL.n25 171.744
R126 VTAIL.n26 VTAIL.n3 171.744
R127 VTAIL.n33 VTAIL.n3 171.744
R128 VTAIL.n34 VTAIL.n33 171.744
R129 VTAIL.n57 VTAIL.n51 171.744
R130 VTAIL.n58 VTAIL.n57 171.744
R131 VTAIL.n58 VTAIL.n47 171.744
R132 VTAIL.n65 VTAIL.n47 171.744
R133 VTAIL.n66 VTAIL.n65 171.744
R134 VTAIL.n66 VTAIL.n43 171.744
R135 VTAIL.n73 VTAIL.n43 171.744
R136 VTAIL.n74 VTAIL.n73 171.744
R137 VTAIL.n97 VTAIL.n91 171.744
R138 VTAIL.n98 VTAIL.n97 171.744
R139 VTAIL.n98 VTAIL.n87 171.744
R140 VTAIL.n105 VTAIL.n87 171.744
R141 VTAIL.n106 VTAIL.n105 171.744
R142 VTAIL.n106 VTAIL.n83 171.744
R143 VTAIL.n113 VTAIL.n83 171.744
R144 VTAIL.n114 VTAIL.n113 171.744
R145 VTAIL.n274 VTAIL.n273 171.744
R146 VTAIL.n273 VTAIL.n243 171.744
R147 VTAIL.n266 VTAIL.n243 171.744
R148 VTAIL.n266 VTAIL.n265 171.744
R149 VTAIL.n265 VTAIL.n247 171.744
R150 VTAIL.n258 VTAIL.n247 171.744
R151 VTAIL.n258 VTAIL.n257 171.744
R152 VTAIL.n257 VTAIL.n251 171.744
R153 VTAIL.n234 VTAIL.n233 171.744
R154 VTAIL.n233 VTAIL.n203 171.744
R155 VTAIL.n226 VTAIL.n203 171.744
R156 VTAIL.n226 VTAIL.n225 171.744
R157 VTAIL.n225 VTAIL.n207 171.744
R158 VTAIL.n218 VTAIL.n207 171.744
R159 VTAIL.n218 VTAIL.n217 171.744
R160 VTAIL.n217 VTAIL.n211 171.744
R161 VTAIL.n194 VTAIL.n193 171.744
R162 VTAIL.n193 VTAIL.n163 171.744
R163 VTAIL.n186 VTAIL.n163 171.744
R164 VTAIL.n186 VTAIL.n185 171.744
R165 VTAIL.n185 VTAIL.n167 171.744
R166 VTAIL.n178 VTAIL.n167 171.744
R167 VTAIL.n178 VTAIL.n177 171.744
R168 VTAIL.n177 VTAIL.n171 171.744
R169 VTAIL.n154 VTAIL.n153 171.744
R170 VTAIL.n153 VTAIL.n123 171.744
R171 VTAIL.n146 VTAIL.n123 171.744
R172 VTAIL.n146 VTAIL.n145 171.744
R173 VTAIL.n145 VTAIL.n127 171.744
R174 VTAIL.n138 VTAIL.n127 171.744
R175 VTAIL.n138 VTAIL.n137 171.744
R176 VTAIL.n137 VTAIL.n131 171.744
R177 VTAIL.t2 VTAIL.n291 85.8723
R178 VTAIL.t1 VTAIL.n11 85.8723
R179 VTAIL.t6 VTAIL.n51 85.8723
R180 VTAIL.t7 VTAIL.n91 85.8723
R181 VTAIL.t4 VTAIL.n251 85.8723
R182 VTAIL.t5 VTAIL.n211 85.8723
R183 VTAIL.t3 VTAIL.n171 85.8723
R184 VTAIL.t0 VTAIL.n131 85.8723
R185 VTAIL.n319 VTAIL.n318 31.2157
R186 VTAIL.n39 VTAIL.n38 31.2157
R187 VTAIL.n79 VTAIL.n78 31.2157
R188 VTAIL.n119 VTAIL.n118 31.2157
R189 VTAIL.n279 VTAIL.n278 31.2157
R190 VTAIL.n239 VTAIL.n238 31.2157
R191 VTAIL.n199 VTAIL.n198 31.2157
R192 VTAIL.n159 VTAIL.n158 31.2157
R193 VTAIL.n319 VTAIL.n279 20.5307
R194 VTAIL.n159 VTAIL.n119 20.5307
R195 VTAIL.n293 VTAIL.n292 16.3891
R196 VTAIL.n13 VTAIL.n12 16.3891
R197 VTAIL.n53 VTAIL.n52 16.3891
R198 VTAIL.n93 VTAIL.n92 16.3891
R199 VTAIL.n253 VTAIL.n252 16.3891
R200 VTAIL.n213 VTAIL.n212 16.3891
R201 VTAIL.n173 VTAIL.n172 16.3891
R202 VTAIL.n133 VTAIL.n132 16.3891
R203 VTAIL.n296 VTAIL.n295 12.8005
R204 VTAIL.n16 VTAIL.n15 12.8005
R205 VTAIL.n56 VTAIL.n55 12.8005
R206 VTAIL.n96 VTAIL.n95 12.8005
R207 VTAIL.n256 VTAIL.n255 12.8005
R208 VTAIL.n216 VTAIL.n215 12.8005
R209 VTAIL.n176 VTAIL.n175 12.8005
R210 VTAIL.n136 VTAIL.n135 12.8005
R211 VTAIL.n299 VTAIL.n290 12.0247
R212 VTAIL.n19 VTAIL.n10 12.0247
R213 VTAIL.n59 VTAIL.n50 12.0247
R214 VTAIL.n99 VTAIL.n90 12.0247
R215 VTAIL.n259 VTAIL.n250 12.0247
R216 VTAIL.n219 VTAIL.n210 12.0247
R217 VTAIL.n179 VTAIL.n170 12.0247
R218 VTAIL.n139 VTAIL.n130 12.0247
R219 VTAIL.n300 VTAIL.n288 11.249
R220 VTAIL.n20 VTAIL.n8 11.249
R221 VTAIL.n60 VTAIL.n48 11.249
R222 VTAIL.n100 VTAIL.n88 11.249
R223 VTAIL.n260 VTAIL.n248 11.249
R224 VTAIL.n220 VTAIL.n208 11.249
R225 VTAIL.n180 VTAIL.n168 11.249
R226 VTAIL.n140 VTAIL.n128 11.249
R227 VTAIL.n304 VTAIL.n303 10.4732
R228 VTAIL.n24 VTAIL.n23 10.4732
R229 VTAIL.n64 VTAIL.n63 10.4732
R230 VTAIL.n104 VTAIL.n103 10.4732
R231 VTAIL.n264 VTAIL.n263 10.4732
R232 VTAIL.n224 VTAIL.n223 10.4732
R233 VTAIL.n184 VTAIL.n183 10.4732
R234 VTAIL.n144 VTAIL.n143 10.4732
R235 VTAIL.n307 VTAIL.n286 9.69747
R236 VTAIL.n27 VTAIL.n6 9.69747
R237 VTAIL.n67 VTAIL.n46 9.69747
R238 VTAIL.n107 VTAIL.n86 9.69747
R239 VTAIL.n267 VTAIL.n246 9.69747
R240 VTAIL.n227 VTAIL.n206 9.69747
R241 VTAIL.n187 VTAIL.n166 9.69747
R242 VTAIL.n147 VTAIL.n126 9.69747
R243 VTAIL.n318 VTAIL.n317 9.45567
R244 VTAIL.n38 VTAIL.n37 9.45567
R245 VTAIL.n78 VTAIL.n77 9.45567
R246 VTAIL.n118 VTAIL.n117 9.45567
R247 VTAIL.n278 VTAIL.n277 9.45567
R248 VTAIL.n238 VTAIL.n237 9.45567
R249 VTAIL.n198 VTAIL.n197 9.45567
R250 VTAIL.n158 VTAIL.n157 9.45567
R251 VTAIL.n317 VTAIL.n316 9.3005
R252 VTAIL.n311 VTAIL.n310 9.3005
R253 VTAIL.n309 VTAIL.n308 9.3005
R254 VTAIL.n286 VTAIL.n285 9.3005
R255 VTAIL.n303 VTAIL.n302 9.3005
R256 VTAIL.n301 VTAIL.n300 9.3005
R257 VTAIL.n290 VTAIL.n289 9.3005
R258 VTAIL.n295 VTAIL.n294 9.3005
R259 VTAIL.n282 VTAIL.n281 9.3005
R260 VTAIL.n37 VTAIL.n36 9.3005
R261 VTAIL.n31 VTAIL.n30 9.3005
R262 VTAIL.n29 VTAIL.n28 9.3005
R263 VTAIL.n6 VTAIL.n5 9.3005
R264 VTAIL.n23 VTAIL.n22 9.3005
R265 VTAIL.n21 VTAIL.n20 9.3005
R266 VTAIL.n10 VTAIL.n9 9.3005
R267 VTAIL.n15 VTAIL.n14 9.3005
R268 VTAIL.n2 VTAIL.n1 9.3005
R269 VTAIL.n77 VTAIL.n76 9.3005
R270 VTAIL.n71 VTAIL.n70 9.3005
R271 VTAIL.n69 VTAIL.n68 9.3005
R272 VTAIL.n46 VTAIL.n45 9.3005
R273 VTAIL.n63 VTAIL.n62 9.3005
R274 VTAIL.n61 VTAIL.n60 9.3005
R275 VTAIL.n50 VTAIL.n49 9.3005
R276 VTAIL.n55 VTAIL.n54 9.3005
R277 VTAIL.n42 VTAIL.n41 9.3005
R278 VTAIL.n117 VTAIL.n116 9.3005
R279 VTAIL.n111 VTAIL.n110 9.3005
R280 VTAIL.n109 VTAIL.n108 9.3005
R281 VTAIL.n86 VTAIL.n85 9.3005
R282 VTAIL.n103 VTAIL.n102 9.3005
R283 VTAIL.n101 VTAIL.n100 9.3005
R284 VTAIL.n90 VTAIL.n89 9.3005
R285 VTAIL.n95 VTAIL.n94 9.3005
R286 VTAIL.n82 VTAIL.n81 9.3005
R287 VTAIL.n277 VTAIL.n276 9.3005
R288 VTAIL.n242 VTAIL.n241 9.3005
R289 VTAIL.n271 VTAIL.n270 9.3005
R290 VTAIL.n269 VTAIL.n268 9.3005
R291 VTAIL.n246 VTAIL.n245 9.3005
R292 VTAIL.n263 VTAIL.n262 9.3005
R293 VTAIL.n261 VTAIL.n260 9.3005
R294 VTAIL.n250 VTAIL.n249 9.3005
R295 VTAIL.n255 VTAIL.n254 9.3005
R296 VTAIL.n237 VTAIL.n236 9.3005
R297 VTAIL.n202 VTAIL.n201 9.3005
R298 VTAIL.n231 VTAIL.n230 9.3005
R299 VTAIL.n229 VTAIL.n228 9.3005
R300 VTAIL.n206 VTAIL.n205 9.3005
R301 VTAIL.n223 VTAIL.n222 9.3005
R302 VTAIL.n221 VTAIL.n220 9.3005
R303 VTAIL.n210 VTAIL.n209 9.3005
R304 VTAIL.n215 VTAIL.n214 9.3005
R305 VTAIL.n197 VTAIL.n196 9.3005
R306 VTAIL.n162 VTAIL.n161 9.3005
R307 VTAIL.n191 VTAIL.n190 9.3005
R308 VTAIL.n189 VTAIL.n188 9.3005
R309 VTAIL.n166 VTAIL.n165 9.3005
R310 VTAIL.n183 VTAIL.n182 9.3005
R311 VTAIL.n181 VTAIL.n180 9.3005
R312 VTAIL.n170 VTAIL.n169 9.3005
R313 VTAIL.n175 VTAIL.n174 9.3005
R314 VTAIL.n157 VTAIL.n156 9.3005
R315 VTAIL.n122 VTAIL.n121 9.3005
R316 VTAIL.n151 VTAIL.n150 9.3005
R317 VTAIL.n149 VTAIL.n148 9.3005
R318 VTAIL.n126 VTAIL.n125 9.3005
R319 VTAIL.n143 VTAIL.n142 9.3005
R320 VTAIL.n141 VTAIL.n140 9.3005
R321 VTAIL.n130 VTAIL.n129 9.3005
R322 VTAIL.n135 VTAIL.n134 9.3005
R323 VTAIL.n308 VTAIL.n284 8.92171
R324 VTAIL.n28 VTAIL.n4 8.92171
R325 VTAIL.n68 VTAIL.n44 8.92171
R326 VTAIL.n108 VTAIL.n84 8.92171
R327 VTAIL.n268 VTAIL.n244 8.92171
R328 VTAIL.n228 VTAIL.n204 8.92171
R329 VTAIL.n188 VTAIL.n164 8.92171
R330 VTAIL.n148 VTAIL.n124 8.92171
R331 VTAIL.n312 VTAIL.n311 8.14595
R332 VTAIL.n32 VTAIL.n31 8.14595
R333 VTAIL.n72 VTAIL.n71 8.14595
R334 VTAIL.n112 VTAIL.n111 8.14595
R335 VTAIL.n272 VTAIL.n271 8.14595
R336 VTAIL.n232 VTAIL.n231 8.14595
R337 VTAIL.n192 VTAIL.n191 8.14595
R338 VTAIL.n152 VTAIL.n151 8.14595
R339 VTAIL.n315 VTAIL.n282 7.3702
R340 VTAIL.n318 VTAIL.n280 7.3702
R341 VTAIL.n35 VTAIL.n2 7.3702
R342 VTAIL.n38 VTAIL.n0 7.3702
R343 VTAIL.n75 VTAIL.n42 7.3702
R344 VTAIL.n78 VTAIL.n40 7.3702
R345 VTAIL.n115 VTAIL.n82 7.3702
R346 VTAIL.n118 VTAIL.n80 7.3702
R347 VTAIL.n278 VTAIL.n240 7.3702
R348 VTAIL.n275 VTAIL.n242 7.3702
R349 VTAIL.n238 VTAIL.n200 7.3702
R350 VTAIL.n235 VTAIL.n202 7.3702
R351 VTAIL.n198 VTAIL.n160 7.3702
R352 VTAIL.n195 VTAIL.n162 7.3702
R353 VTAIL.n158 VTAIL.n120 7.3702
R354 VTAIL.n155 VTAIL.n122 7.3702
R355 VTAIL.n316 VTAIL.n315 6.59444
R356 VTAIL.n316 VTAIL.n280 6.59444
R357 VTAIL.n36 VTAIL.n35 6.59444
R358 VTAIL.n36 VTAIL.n0 6.59444
R359 VTAIL.n76 VTAIL.n75 6.59444
R360 VTAIL.n76 VTAIL.n40 6.59444
R361 VTAIL.n116 VTAIL.n115 6.59444
R362 VTAIL.n116 VTAIL.n80 6.59444
R363 VTAIL.n276 VTAIL.n240 6.59444
R364 VTAIL.n276 VTAIL.n275 6.59444
R365 VTAIL.n236 VTAIL.n200 6.59444
R366 VTAIL.n236 VTAIL.n235 6.59444
R367 VTAIL.n196 VTAIL.n160 6.59444
R368 VTAIL.n196 VTAIL.n195 6.59444
R369 VTAIL.n156 VTAIL.n120 6.59444
R370 VTAIL.n156 VTAIL.n155 6.59444
R371 VTAIL.n312 VTAIL.n282 5.81868
R372 VTAIL.n32 VTAIL.n2 5.81868
R373 VTAIL.n72 VTAIL.n42 5.81868
R374 VTAIL.n112 VTAIL.n82 5.81868
R375 VTAIL.n272 VTAIL.n242 5.81868
R376 VTAIL.n232 VTAIL.n202 5.81868
R377 VTAIL.n192 VTAIL.n162 5.81868
R378 VTAIL.n152 VTAIL.n122 5.81868
R379 VTAIL.n311 VTAIL.n284 5.04292
R380 VTAIL.n31 VTAIL.n4 5.04292
R381 VTAIL.n71 VTAIL.n44 5.04292
R382 VTAIL.n111 VTAIL.n84 5.04292
R383 VTAIL.n271 VTAIL.n244 5.04292
R384 VTAIL.n231 VTAIL.n204 5.04292
R385 VTAIL.n191 VTAIL.n164 5.04292
R386 VTAIL.n151 VTAIL.n124 5.04292
R387 VTAIL.n308 VTAIL.n307 4.26717
R388 VTAIL.n28 VTAIL.n27 4.26717
R389 VTAIL.n68 VTAIL.n67 4.26717
R390 VTAIL.n108 VTAIL.n107 4.26717
R391 VTAIL.n268 VTAIL.n267 4.26717
R392 VTAIL.n228 VTAIL.n227 4.26717
R393 VTAIL.n188 VTAIL.n187 4.26717
R394 VTAIL.n148 VTAIL.n147 4.26717
R395 VTAIL.n294 VTAIL.n293 3.71019
R396 VTAIL.n14 VTAIL.n13 3.71019
R397 VTAIL.n54 VTAIL.n53 3.71019
R398 VTAIL.n94 VTAIL.n93 3.71019
R399 VTAIL.n254 VTAIL.n253 3.71019
R400 VTAIL.n214 VTAIL.n213 3.71019
R401 VTAIL.n174 VTAIL.n173 3.71019
R402 VTAIL.n134 VTAIL.n133 3.71019
R403 VTAIL.n304 VTAIL.n286 3.49141
R404 VTAIL.n24 VTAIL.n6 3.49141
R405 VTAIL.n64 VTAIL.n46 3.49141
R406 VTAIL.n104 VTAIL.n86 3.49141
R407 VTAIL.n264 VTAIL.n246 3.49141
R408 VTAIL.n224 VTAIL.n206 3.49141
R409 VTAIL.n184 VTAIL.n166 3.49141
R410 VTAIL.n144 VTAIL.n126 3.49141
R411 VTAIL.n303 VTAIL.n288 2.71565
R412 VTAIL.n23 VTAIL.n8 2.71565
R413 VTAIL.n63 VTAIL.n48 2.71565
R414 VTAIL.n103 VTAIL.n88 2.71565
R415 VTAIL.n263 VTAIL.n248 2.71565
R416 VTAIL.n223 VTAIL.n208 2.71565
R417 VTAIL.n183 VTAIL.n168 2.71565
R418 VTAIL.n143 VTAIL.n128 2.71565
R419 VTAIL.n300 VTAIL.n299 1.93989
R420 VTAIL.n20 VTAIL.n19 1.93989
R421 VTAIL.n60 VTAIL.n59 1.93989
R422 VTAIL.n100 VTAIL.n99 1.93989
R423 VTAIL.n260 VTAIL.n259 1.93989
R424 VTAIL.n220 VTAIL.n219 1.93989
R425 VTAIL.n180 VTAIL.n179 1.93989
R426 VTAIL.n140 VTAIL.n139 1.93989
R427 VTAIL.n199 VTAIL.n159 1.7936
R428 VTAIL.n279 VTAIL.n239 1.7936
R429 VTAIL.n119 VTAIL.n79 1.7936
R430 VTAIL.n296 VTAIL.n290 1.16414
R431 VTAIL.n16 VTAIL.n10 1.16414
R432 VTAIL.n56 VTAIL.n50 1.16414
R433 VTAIL.n96 VTAIL.n90 1.16414
R434 VTAIL.n256 VTAIL.n250 1.16414
R435 VTAIL.n216 VTAIL.n210 1.16414
R436 VTAIL.n176 VTAIL.n170 1.16414
R437 VTAIL.n136 VTAIL.n130 1.16414
R438 VTAIL VTAIL.n39 0.955241
R439 VTAIL VTAIL.n319 0.838862
R440 VTAIL.n239 VTAIL.n199 0.470328
R441 VTAIL.n79 VTAIL.n39 0.470328
R442 VTAIL.n295 VTAIL.n292 0.388379
R443 VTAIL.n15 VTAIL.n12 0.388379
R444 VTAIL.n55 VTAIL.n52 0.388379
R445 VTAIL.n95 VTAIL.n92 0.388379
R446 VTAIL.n255 VTAIL.n252 0.388379
R447 VTAIL.n215 VTAIL.n212 0.388379
R448 VTAIL.n175 VTAIL.n172 0.388379
R449 VTAIL.n135 VTAIL.n132 0.388379
R450 VTAIL.n294 VTAIL.n289 0.155672
R451 VTAIL.n301 VTAIL.n289 0.155672
R452 VTAIL.n302 VTAIL.n301 0.155672
R453 VTAIL.n302 VTAIL.n285 0.155672
R454 VTAIL.n309 VTAIL.n285 0.155672
R455 VTAIL.n310 VTAIL.n309 0.155672
R456 VTAIL.n310 VTAIL.n281 0.155672
R457 VTAIL.n317 VTAIL.n281 0.155672
R458 VTAIL.n14 VTAIL.n9 0.155672
R459 VTAIL.n21 VTAIL.n9 0.155672
R460 VTAIL.n22 VTAIL.n21 0.155672
R461 VTAIL.n22 VTAIL.n5 0.155672
R462 VTAIL.n29 VTAIL.n5 0.155672
R463 VTAIL.n30 VTAIL.n29 0.155672
R464 VTAIL.n30 VTAIL.n1 0.155672
R465 VTAIL.n37 VTAIL.n1 0.155672
R466 VTAIL.n54 VTAIL.n49 0.155672
R467 VTAIL.n61 VTAIL.n49 0.155672
R468 VTAIL.n62 VTAIL.n61 0.155672
R469 VTAIL.n62 VTAIL.n45 0.155672
R470 VTAIL.n69 VTAIL.n45 0.155672
R471 VTAIL.n70 VTAIL.n69 0.155672
R472 VTAIL.n70 VTAIL.n41 0.155672
R473 VTAIL.n77 VTAIL.n41 0.155672
R474 VTAIL.n94 VTAIL.n89 0.155672
R475 VTAIL.n101 VTAIL.n89 0.155672
R476 VTAIL.n102 VTAIL.n101 0.155672
R477 VTAIL.n102 VTAIL.n85 0.155672
R478 VTAIL.n109 VTAIL.n85 0.155672
R479 VTAIL.n110 VTAIL.n109 0.155672
R480 VTAIL.n110 VTAIL.n81 0.155672
R481 VTAIL.n117 VTAIL.n81 0.155672
R482 VTAIL.n277 VTAIL.n241 0.155672
R483 VTAIL.n270 VTAIL.n241 0.155672
R484 VTAIL.n270 VTAIL.n269 0.155672
R485 VTAIL.n269 VTAIL.n245 0.155672
R486 VTAIL.n262 VTAIL.n245 0.155672
R487 VTAIL.n262 VTAIL.n261 0.155672
R488 VTAIL.n261 VTAIL.n249 0.155672
R489 VTAIL.n254 VTAIL.n249 0.155672
R490 VTAIL.n237 VTAIL.n201 0.155672
R491 VTAIL.n230 VTAIL.n201 0.155672
R492 VTAIL.n230 VTAIL.n229 0.155672
R493 VTAIL.n229 VTAIL.n205 0.155672
R494 VTAIL.n222 VTAIL.n205 0.155672
R495 VTAIL.n222 VTAIL.n221 0.155672
R496 VTAIL.n221 VTAIL.n209 0.155672
R497 VTAIL.n214 VTAIL.n209 0.155672
R498 VTAIL.n197 VTAIL.n161 0.155672
R499 VTAIL.n190 VTAIL.n161 0.155672
R500 VTAIL.n190 VTAIL.n189 0.155672
R501 VTAIL.n189 VTAIL.n165 0.155672
R502 VTAIL.n182 VTAIL.n165 0.155672
R503 VTAIL.n182 VTAIL.n181 0.155672
R504 VTAIL.n181 VTAIL.n169 0.155672
R505 VTAIL.n174 VTAIL.n169 0.155672
R506 VTAIL.n157 VTAIL.n121 0.155672
R507 VTAIL.n150 VTAIL.n121 0.155672
R508 VTAIL.n150 VTAIL.n149 0.155672
R509 VTAIL.n149 VTAIL.n125 0.155672
R510 VTAIL.n142 VTAIL.n125 0.155672
R511 VTAIL.n142 VTAIL.n141 0.155672
R512 VTAIL.n141 VTAIL.n129 0.155672
R513 VTAIL.n134 VTAIL.n129 0.155672
R514 VDD1 VDD1.n1 120.323
R515 VDD1 VDD1.n0 84.3909
R516 VDD1.n0 VDD1.t2 4.39901
R517 VDD1.n0 VDD1.t3 4.39901
R518 VDD1.n1 VDD1.t0 4.39901
R519 VDD1.n1 VDD1.t1 4.39901
R520 B.n267 B.n266 585
R521 B.n265 B.n80 585
R522 B.n264 B.n263 585
R523 B.n262 B.n81 585
R524 B.n261 B.n260 585
R525 B.n259 B.n82 585
R526 B.n258 B.n257 585
R527 B.n256 B.n83 585
R528 B.n255 B.n254 585
R529 B.n253 B.n84 585
R530 B.n252 B.n251 585
R531 B.n250 B.n85 585
R532 B.n249 B.n248 585
R533 B.n247 B.n86 585
R534 B.n246 B.n245 585
R535 B.n244 B.n87 585
R536 B.n243 B.n242 585
R537 B.n241 B.n88 585
R538 B.n240 B.n239 585
R539 B.n238 B.n89 585
R540 B.n237 B.n236 585
R541 B.n235 B.n90 585
R542 B.n234 B.n233 585
R543 B.n232 B.n91 585
R544 B.n231 B.n230 585
R545 B.n229 B.n92 585
R546 B.n228 B.n227 585
R547 B.n226 B.n93 585
R548 B.n224 B.n223 585
R549 B.n222 B.n96 585
R550 B.n221 B.n220 585
R551 B.n219 B.n97 585
R552 B.n218 B.n217 585
R553 B.n216 B.n98 585
R554 B.n215 B.n214 585
R555 B.n213 B.n99 585
R556 B.n212 B.n211 585
R557 B.n210 B.n100 585
R558 B.n209 B.n208 585
R559 B.n204 B.n101 585
R560 B.n203 B.n202 585
R561 B.n201 B.n102 585
R562 B.n200 B.n199 585
R563 B.n198 B.n103 585
R564 B.n197 B.n196 585
R565 B.n195 B.n104 585
R566 B.n194 B.n193 585
R567 B.n192 B.n105 585
R568 B.n191 B.n190 585
R569 B.n189 B.n106 585
R570 B.n188 B.n187 585
R571 B.n186 B.n107 585
R572 B.n185 B.n184 585
R573 B.n183 B.n108 585
R574 B.n182 B.n181 585
R575 B.n180 B.n109 585
R576 B.n179 B.n178 585
R577 B.n177 B.n110 585
R578 B.n176 B.n175 585
R579 B.n174 B.n111 585
R580 B.n173 B.n172 585
R581 B.n171 B.n112 585
R582 B.n170 B.n169 585
R583 B.n168 B.n113 585
R584 B.n167 B.n166 585
R585 B.n165 B.n114 585
R586 B.n268 B.n79 585
R587 B.n270 B.n269 585
R588 B.n271 B.n78 585
R589 B.n273 B.n272 585
R590 B.n274 B.n77 585
R591 B.n276 B.n275 585
R592 B.n277 B.n76 585
R593 B.n279 B.n278 585
R594 B.n280 B.n75 585
R595 B.n282 B.n281 585
R596 B.n283 B.n74 585
R597 B.n285 B.n284 585
R598 B.n286 B.n73 585
R599 B.n288 B.n287 585
R600 B.n289 B.n72 585
R601 B.n291 B.n290 585
R602 B.n292 B.n71 585
R603 B.n294 B.n293 585
R604 B.n295 B.n70 585
R605 B.n297 B.n296 585
R606 B.n298 B.n69 585
R607 B.n300 B.n299 585
R608 B.n301 B.n68 585
R609 B.n303 B.n302 585
R610 B.n304 B.n67 585
R611 B.n306 B.n305 585
R612 B.n307 B.n66 585
R613 B.n309 B.n308 585
R614 B.n310 B.n65 585
R615 B.n312 B.n311 585
R616 B.n313 B.n64 585
R617 B.n315 B.n314 585
R618 B.n316 B.n63 585
R619 B.n318 B.n317 585
R620 B.n319 B.n62 585
R621 B.n321 B.n320 585
R622 B.n322 B.n61 585
R623 B.n324 B.n323 585
R624 B.n325 B.n60 585
R625 B.n327 B.n326 585
R626 B.n328 B.n59 585
R627 B.n330 B.n329 585
R628 B.n331 B.n58 585
R629 B.n333 B.n332 585
R630 B.n334 B.n57 585
R631 B.n336 B.n335 585
R632 B.n337 B.n56 585
R633 B.n339 B.n338 585
R634 B.n340 B.n55 585
R635 B.n342 B.n341 585
R636 B.n343 B.n54 585
R637 B.n345 B.n344 585
R638 B.n346 B.n53 585
R639 B.n348 B.n347 585
R640 B.n448 B.n15 585
R641 B.n447 B.n446 585
R642 B.n445 B.n16 585
R643 B.n444 B.n443 585
R644 B.n442 B.n17 585
R645 B.n441 B.n440 585
R646 B.n439 B.n18 585
R647 B.n438 B.n437 585
R648 B.n436 B.n19 585
R649 B.n435 B.n434 585
R650 B.n433 B.n20 585
R651 B.n432 B.n431 585
R652 B.n430 B.n21 585
R653 B.n429 B.n428 585
R654 B.n427 B.n22 585
R655 B.n426 B.n425 585
R656 B.n424 B.n23 585
R657 B.n423 B.n422 585
R658 B.n421 B.n24 585
R659 B.n420 B.n419 585
R660 B.n418 B.n25 585
R661 B.n417 B.n416 585
R662 B.n415 B.n26 585
R663 B.n414 B.n413 585
R664 B.n412 B.n27 585
R665 B.n411 B.n410 585
R666 B.n409 B.n28 585
R667 B.n408 B.n407 585
R668 B.n405 B.n29 585
R669 B.n404 B.n403 585
R670 B.n402 B.n32 585
R671 B.n401 B.n400 585
R672 B.n399 B.n33 585
R673 B.n398 B.n397 585
R674 B.n396 B.n34 585
R675 B.n395 B.n394 585
R676 B.n393 B.n35 585
R677 B.n392 B.n391 585
R678 B.n390 B.n389 585
R679 B.n388 B.n39 585
R680 B.n387 B.n386 585
R681 B.n385 B.n40 585
R682 B.n384 B.n383 585
R683 B.n382 B.n41 585
R684 B.n381 B.n380 585
R685 B.n379 B.n42 585
R686 B.n378 B.n377 585
R687 B.n376 B.n43 585
R688 B.n375 B.n374 585
R689 B.n373 B.n44 585
R690 B.n372 B.n371 585
R691 B.n370 B.n45 585
R692 B.n369 B.n368 585
R693 B.n367 B.n46 585
R694 B.n366 B.n365 585
R695 B.n364 B.n47 585
R696 B.n363 B.n362 585
R697 B.n361 B.n48 585
R698 B.n360 B.n359 585
R699 B.n358 B.n49 585
R700 B.n357 B.n356 585
R701 B.n355 B.n50 585
R702 B.n354 B.n353 585
R703 B.n352 B.n51 585
R704 B.n351 B.n350 585
R705 B.n349 B.n52 585
R706 B.n450 B.n449 585
R707 B.n451 B.n14 585
R708 B.n453 B.n452 585
R709 B.n454 B.n13 585
R710 B.n456 B.n455 585
R711 B.n457 B.n12 585
R712 B.n459 B.n458 585
R713 B.n460 B.n11 585
R714 B.n462 B.n461 585
R715 B.n463 B.n10 585
R716 B.n465 B.n464 585
R717 B.n466 B.n9 585
R718 B.n468 B.n467 585
R719 B.n469 B.n8 585
R720 B.n471 B.n470 585
R721 B.n472 B.n7 585
R722 B.n474 B.n473 585
R723 B.n475 B.n6 585
R724 B.n477 B.n476 585
R725 B.n478 B.n5 585
R726 B.n480 B.n479 585
R727 B.n481 B.n4 585
R728 B.n483 B.n482 585
R729 B.n484 B.n3 585
R730 B.n486 B.n485 585
R731 B.n487 B.n0 585
R732 B.n2 B.n1 585
R733 B.n128 B.n127 585
R734 B.n129 B.n126 585
R735 B.n131 B.n130 585
R736 B.n132 B.n125 585
R737 B.n134 B.n133 585
R738 B.n135 B.n124 585
R739 B.n137 B.n136 585
R740 B.n138 B.n123 585
R741 B.n140 B.n139 585
R742 B.n141 B.n122 585
R743 B.n143 B.n142 585
R744 B.n144 B.n121 585
R745 B.n146 B.n145 585
R746 B.n147 B.n120 585
R747 B.n149 B.n148 585
R748 B.n150 B.n119 585
R749 B.n152 B.n151 585
R750 B.n153 B.n118 585
R751 B.n155 B.n154 585
R752 B.n156 B.n117 585
R753 B.n158 B.n157 585
R754 B.n159 B.n116 585
R755 B.n161 B.n160 585
R756 B.n162 B.n115 585
R757 B.n164 B.n163 585
R758 B.n165 B.n164 468.476
R759 B.n266 B.n79 468.476
R760 B.n349 B.n348 468.476
R761 B.n450 B.n15 468.476
R762 B.n94 B.t1 333.216
R763 B.n36 B.t11 333.216
R764 B.n205 B.t7 333.216
R765 B.n30 B.t5 333.216
R766 B.n205 B.t6 308.034
R767 B.n94 B.t0 308.034
R768 B.n36 B.t9 308.034
R769 B.n30 B.t3 308.034
R770 B.n95 B.t2 292.877
R771 B.n37 B.t10 292.877
R772 B.n206 B.t8 292.877
R773 B.n31 B.t4 292.877
R774 B.n489 B.n488 256.663
R775 B.n488 B.n487 235.042
R776 B.n488 B.n2 235.042
R777 B.n166 B.n165 163.367
R778 B.n166 B.n113 163.367
R779 B.n170 B.n113 163.367
R780 B.n171 B.n170 163.367
R781 B.n172 B.n171 163.367
R782 B.n172 B.n111 163.367
R783 B.n176 B.n111 163.367
R784 B.n177 B.n176 163.367
R785 B.n178 B.n177 163.367
R786 B.n178 B.n109 163.367
R787 B.n182 B.n109 163.367
R788 B.n183 B.n182 163.367
R789 B.n184 B.n183 163.367
R790 B.n184 B.n107 163.367
R791 B.n188 B.n107 163.367
R792 B.n189 B.n188 163.367
R793 B.n190 B.n189 163.367
R794 B.n190 B.n105 163.367
R795 B.n194 B.n105 163.367
R796 B.n195 B.n194 163.367
R797 B.n196 B.n195 163.367
R798 B.n196 B.n103 163.367
R799 B.n200 B.n103 163.367
R800 B.n201 B.n200 163.367
R801 B.n202 B.n201 163.367
R802 B.n202 B.n101 163.367
R803 B.n209 B.n101 163.367
R804 B.n210 B.n209 163.367
R805 B.n211 B.n210 163.367
R806 B.n211 B.n99 163.367
R807 B.n215 B.n99 163.367
R808 B.n216 B.n215 163.367
R809 B.n217 B.n216 163.367
R810 B.n217 B.n97 163.367
R811 B.n221 B.n97 163.367
R812 B.n222 B.n221 163.367
R813 B.n223 B.n222 163.367
R814 B.n223 B.n93 163.367
R815 B.n228 B.n93 163.367
R816 B.n229 B.n228 163.367
R817 B.n230 B.n229 163.367
R818 B.n230 B.n91 163.367
R819 B.n234 B.n91 163.367
R820 B.n235 B.n234 163.367
R821 B.n236 B.n235 163.367
R822 B.n236 B.n89 163.367
R823 B.n240 B.n89 163.367
R824 B.n241 B.n240 163.367
R825 B.n242 B.n241 163.367
R826 B.n242 B.n87 163.367
R827 B.n246 B.n87 163.367
R828 B.n247 B.n246 163.367
R829 B.n248 B.n247 163.367
R830 B.n248 B.n85 163.367
R831 B.n252 B.n85 163.367
R832 B.n253 B.n252 163.367
R833 B.n254 B.n253 163.367
R834 B.n254 B.n83 163.367
R835 B.n258 B.n83 163.367
R836 B.n259 B.n258 163.367
R837 B.n260 B.n259 163.367
R838 B.n260 B.n81 163.367
R839 B.n264 B.n81 163.367
R840 B.n265 B.n264 163.367
R841 B.n266 B.n265 163.367
R842 B.n348 B.n53 163.367
R843 B.n344 B.n53 163.367
R844 B.n344 B.n343 163.367
R845 B.n343 B.n342 163.367
R846 B.n342 B.n55 163.367
R847 B.n338 B.n55 163.367
R848 B.n338 B.n337 163.367
R849 B.n337 B.n336 163.367
R850 B.n336 B.n57 163.367
R851 B.n332 B.n57 163.367
R852 B.n332 B.n331 163.367
R853 B.n331 B.n330 163.367
R854 B.n330 B.n59 163.367
R855 B.n326 B.n59 163.367
R856 B.n326 B.n325 163.367
R857 B.n325 B.n324 163.367
R858 B.n324 B.n61 163.367
R859 B.n320 B.n61 163.367
R860 B.n320 B.n319 163.367
R861 B.n319 B.n318 163.367
R862 B.n318 B.n63 163.367
R863 B.n314 B.n63 163.367
R864 B.n314 B.n313 163.367
R865 B.n313 B.n312 163.367
R866 B.n312 B.n65 163.367
R867 B.n308 B.n65 163.367
R868 B.n308 B.n307 163.367
R869 B.n307 B.n306 163.367
R870 B.n306 B.n67 163.367
R871 B.n302 B.n67 163.367
R872 B.n302 B.n301 163.367
R873 B.n301 B.n300 163.367
R874 B.n300 B.n69 163.367
R875 B.n296 B.n69 163.367
R876 B.n296 B.n295 163.367
R877 B.n295 B.n294 163.367
R878 B.n294 B.n71 163.367
R879 B.n290 B.n71 163.367
R880 B.n290 B.n289 163.367
R881 B.n289 B.n288 163.367
R882 B.n288 B.n73 163.367
R883 B.n284 B.n73 163.367
R884 B.n284 B.n283 163.367
R885 B.n283 B.n282 163.367
R886 B.n282 B.n75 163.367
R887 B.n278 B.n75 163.367
R888 B.n278 B.n277 163.367
R889 B.n277 B.n276 163.367
R890 B.n276 B.n77 163.367
R891 B.n272 B.n77 163.367
R892 B.n272 B.n271 163.367
R893 B.n271 B.n270 163.367
R894 B.n270 B.n79 163.367
R895 B.n446 B.n15 163.367
R896 B.n446 B.n445 163.367
R897 B.n445 B.n444 163.367
R898 B.n444 B.n17 163.367
R899 B.n440 B.n17 163.367
R900 B.n440 B.n439 163.367
R901 B.n439 B.n438 163.367
R902 B.n438 B.n19 163.367
R903 B.n434 B.n19 163.367
R904 B.n434 B.n433 163.367
R905 B.n433 B.n432 163.367
R906 B.n432 B.n21 163.367
R907 B.n428 B.n21 163.367
R908 B.n428 B.n427 163.367
R909 B.n427 B.n426 163.367
R910 B.n426 B.n23 163.367
R911 B.n422 B.n23 163.367
R912 B.n422 B.n421 163.367
R913 B.n421 B.n420 163.367
R914 B.n420 B.n25 163.367
R915 B.n416 B.n25 163.367
R916 B.n416 B.n415 163.367
R917 B.n415 B.n414 163.367
R918 B.n414 B.n27 163.367
R919 B.n410 B.n27 163.367
R920 B.n410 B.n409 163.367
R921 B.n409 B.n408 163.367
R922 B.n408 B.n29 163.367
R923 B.n403 B.n29 163.367
R924 B.n403 B.n402 163.367
R925 B.n402 B.n401 163.367
R926 B.n401 B.n33 163.367
R927 B.n397 B.n33 163.367
R928 B.n397 B.n396 163.367
R929 B.n396 B.n395 163.367
R930 B.n395 B.n35 163.367
R931 B.n391 B.n35 163.367
R932 B.n391 B.n390 163.367
R933 B.n390 B.n39 163.367
R934 B.n386 B.n39 163.367
R935 B.n386 B.n385 163.367
R936 B.n385 B.n384 163.367
R937 B.n384 B.n41 163.367
R938 B.n380 B.n41 163.367
R939 B.n380 B.n379 163.367
R940 B.n379 B.n378 163.367
R941 B.n378 B.n43 163.367
R942 B.n374 B.n43 163.367
R943 B.n374 B.n373 163.367
R944 B.n373 B.n372 163.367
R945 B.n372 B.n45 163.367
R946 B.n368 B.n45 163.367
R947 B.n368 B.n367 163.367
R948 B.n367 B.n366 163.367
R949 B.n366 B.n47 163.367
R950 B.n362 B.n47 163.367
R951 B.n362 B.n361 163.367
R952 B.n361 B.n360 163.367
R953 B.n360 B.n49 163.367
R954 B.n356 B.n49 163.367
R955 B.n356 B.n355 163.367
R956 B.n355 B.n354 163.367
R957 B.n354 B.n51 163.367
R958 B.n350 B.n51 163.367
R959 B.n350 B.n349 163.367
R960 B.n451 B.n450 163.367
R961 B.n452 B.n451 163.367
R962 B.n452 B.n13 163.367
R963 B.n456 B.n13 163.367
R964 B.n457 B.n456 163.367
R965 B.n458 B.n457 163.367
R966 B.n458 B.n11 163.367
R967 B.n462 B.n11 163.367
R968 B.n463 B.n462 163.367
R969 B.n464 B.n463 163.367
R970 B.n464 B.n9 163.367
R971 B.n468 B.n9 163.367
R972 B.n469 B.n468 163.367
R973 B.n470 B.n469 163.367
R974 B.n470 B.n7 163.367
R975 B.n474 B.n7 163.367
R976 B.n475 B.n474 163.367
R977 B.n476 B.n475 163.367
R978 B.n476 B.n5 163.367
R979 B.n480 B.n5 163.367
R980 B.n481 B.n480 163.367
R981 B.n482 B.n481 163.367
R982 B.n482 B.n3 163.367
R983 B.n486 B.n3 163.367
R984 B.n487 B.n486 163.367
R985 B.n128 B.n2 163.367
R986 B.n129 B.n128 163.367
R987 B.n130 B.n129 163.367
R988 B.n130 B.n125 163.367
R989 B.n134 B.n125 163.367
R990 B.n135 B.n134 163.367
R991 B.n136 B.n135 163.367
R992 B.n136 B.n123 163.367
R993 B.n140 B.n123 163.367
R994 B.n141 B.n140 163.367
R995 B.n142 B.n141 163.367
R996 B.n142 B.n121 163.367
R997 B.n146 B.n121 163.367
R998 B.n147 B.n146 163.367
R999 B.n148 B.n147 163.367
R1000 B.n148 B.n119 163.367
R1001 B.n152 B.n119 163.367
R1002 B.n153 B.n152 163.367
R1003 B.n154 B.n153 163.367
R1004 B.n154 B.n117 163.367
R1005 B.n158 B.n117 163.367
R1006 B.n159 B.n158 163.367
R1007 B.n160 B.n159 163.367
R1008 B.n160 B.n115 163.367
R1009 B.n164 B.n115 163.367
R1010 B.n207 B.n206 59.5399
R1011 B.n225 B.n95 59.5399
R1012 B.n38 B.n37 59.5399
R1013 B.n406 B.n31 59.5399
R1014 B.n206 B.n205 40.3399
R1015 B.n95 B.n94 40.3399
R1016 B.n37 B.n36 40.3399
R1017 B.n31 B.n30 40.3399
R1018 B.n449 B.n448 30.4395
R1019 B.n347 B.n52 30.4395
R1020 B.n268 B.n267 30.4395
R1021 B.n163 B.n114 30.4395
R1022 B B.n489 18.0485
R1023 B.n449 B.n14 10.6151
R1024 B.n453 B.n14 10.6151
R1025 B.n454 B.n453 10.6151
R1026 B.n455 B.n454 10.6151
R1027 B.n455 B.n12 10.6151
R1028 B.n459 B.n12 10.6151
R1029 B.n460 B.n459 10.6151
R1030 B.n461 B.n460 10.6151
R1031 B.n461 B.n10 10.6151
R1032 B.n465 B.n10 10.6151
R1033 B.n466 B.n465 10.6151
R1034 B.n467 B.n466 10.6151
R1035 B.n467 B.n8 10.6151
R1036 B.n471 B.n8 10.6151
R1037 B.n472 B.n471 10.6151
R1038 B.n473 B.n472 10.6151
R1039 B.n473 B.n6 10.6151
R1040 B.n477 B.n6 10.6151
R1041 B.n478 B.n477 10.6151
R1042 B.n479 B.n478 10.6151
R1043 B.n479 B.n4 10.6151
R1044 B.n483 B.n4 10.6151
R1045 B.n484 B.n483 10.6151
R1046 B.n485 B.n484 10.6151
R1047 B.n485 B.n0 10.6151
R1048 B.n448 B.n447 10.6151
R1049 B.n447 B.n16 10.6151
R1050 B.n443 B.n16 10.6151
R1051 B.n443 B.n442 10.6151
R1052 B.n442 B.n441 10.6151
R1053 B.n441 B.n18 10.6151
R1054 B.n437 B.n18 10.6151
R1055 B.n437 B.n436 10.6151
R1056 B.n436 B.n435 10.6151
R1057 B.n435 B.n20 10.6151
R1058 B.n431 B.n20 10.6151
R1059 B.n431 B.n430 10.6151
R1060 B.n430 B.n429 10.6151
R1061 B.n429 B.n22 10.6151
R1062 B.n425 B.n22 10.6151
R1063 B.n425 B.n424 10.6151
R1064 B.n424 B.n423 10.6151
R1065 B.n423 B.n24 10.6151
R1066 B.n419 B.n24 10.6151
R1067 B.n419 B.n418 10.6151
R1068 B.n418 B.n417 10.6151
R1069 B.n417 B.n26 10.6151
R1070 B.n413 B.n26 10.6151
R1071 B.n413 B.n412 10.6151
R1072 B.n412 B.n411 10.6151
R1073 B.n411 B.n28 10.6151
R1074 B.n407 B.n28 10.6151
R1075 B.n405 B.n404 10.6151
R1076 B.n404 B.n32 10.6151
R1077 B.n400 B.n32 10.6151
R1078 B.n400 B.n399 10.6151
R1079 B.n399 B.n398 10.6151
R1080 B.n398 B.n34 10.6151
R1081 B.n394 B.n34 10.6151
R1082 B.n394 B.n393 10.6151
R1083 B.n393 B.n392 10.6151
R1084 B.n389 B.n388 10.6151
R1085 B.n388 B.n387 10.6151
R1086 B.n387 B.n40 10.6151
R1087 B.n383 B.n40 10.6151
R1088 B.n383 B.n382 10.6151
R1089 B.n382 B.n381 10.6151
R1090 B.n381 B.n42 10.6151
R1091 B.n377 B.n42 10.6151
R1092 B.n377 B.n376 10.6151
R1093 B.n376 B.n375 10.6151
R1094 B.n375 B.n44 10.6151
R1095 B.n371 B.n44 10.6151
R1096 B.n371 B.n370 10.6151
R1097 B.n370 B.n369 10.6151
R1098 B.n369 B.n46 10.6151
R1099 B.n365 B.n46 10.6151
R1100 B.n365 B.n364 10.6151
R1101 B.n364 B.n363 10.6151
R1102 B.n363 B.n48 10.6151
R1103 B.n359 B.n48 10.6151
R1104 B.n359 B.n358 10.6151
R1105 B.n358 B.n357 10.6151
R1106 B.n357 B.n50 10.6151
R1107 B.n353 B.n50 10.6151
R1108 B.n353 B.n352 10.6151
R1109 B.n352 B.n351 10.6151
R1110 B.n351 B.n52 10.6151
R1111 B.n347 B.n346 10.6151
R1112 B.n346 B.n345 10.6151
R1113 B.n345 B.n54 10.6151
R1114 B.n341 B.n54 10.6151
R1115 B.n341 B.n340 10.6151
R1116 B.n340 B.n339 10.6151
R1117 B.n339 B.n56 10.6151
R1118 B.n335 B.n56 10.6151
R1119 B.n335 B.n334 10.6151
R1120 B.n334 B.n333 10.6151
R1121 B.n333 B.n58 10.6151
R1122 B.n329 B.n58 10.6151
R1123 B.n329 B.n328 10.6151
R1124 B.n328 B.n327 10.6151
R1125 B.n327 B.n60 10.6151
R1126 B.n323 B.n60 10.6151
R1127 B.n323 B.n322 10.6151
R1128 B.n322 B.n321 10.6151
R1129 B.n321 B.n62 10.6151
R1130 B.n317 B.n62 10.6151
R1131 B.n317 B.n316 10.6151
R1132 B.n316 B.n315 10.6151
R1133 B.n315 B.n64 10.6151
R1134 B.n311 B.n64 10.6151
R1135 B.n311 B.n310 10.6151
R1136 B.n310 B.n309 10.6151
R1137 B.n309 B.n66 10.6151
R1138 B.n305 B.n66 10.6151
R1139 B.n305 B.n304 10.6151
R1140 B.n304 B.n303 10.6151
R1141 B.n303 B.n68 10.6151
R1142 B.n299 B.n68 10.6151
R1143 B.n299 B.n298 10.6151
R1144 B.n298 B.n297 10.6151
R1145 B.n297 B.n70 10.6151
R1146 B.n293 B.n70 10.6151
R1147 B.n293 B.n292 10.6151
R1148 B.n292 B.n291 10.6151
R1149 B.n291 B.n72 10.6151
R1150 B.n287 B.n72 10.6151
R1151 B.n287 B.n286 10.6151
R1152 B.n286 B.n285 10.6151
R1153 B.n285 B.n74 10.6151
R1154 B.n281 B.n74 10.6151
R1155 B.n281 B.n280 10.6151
R1156 B.n280 B.n279 10.6151
R1157 B.n279 B.n76 10.6151
R1158 B.n275 B.n76 10.6151
R1159 B.n275 B.n274 10.6151
R1160 B.n274 B.n273 10.6151
R1161 B.n273 B.n78 10.6151
R1162 B.n269 B.n78 10.6151
R1163 B.n269 B.n268 10.6151
R1164 B.n127 B.n1 10.6151
R1165 B.n127 B.n126 10.6151
R1166 B.n131 B.n126 10.6151
R1167 B.n132 B.n131 10.6151
R1168 B.n133 B.n132 10.6151
R1169 B.n133 B.n124 10.6151
R1170 B.n137 B.n124 10.6151
R1171 B.n138 B.n137 10.6151
R1172 B.n139 B.n138 10.6151
R1173 B.n139 B.n122 10.6151
R1174 B.n143 B.n122 10.6151
R1175 B.n144 B.n143 10.6151
R1176 B.n145 B.n144 10.6151
R1177 B.n145 B.n120 10.6151
R1178 B.n149 B.n120 10.6151
R1179 B.n150 B.n149 10.6151
R1180 B.n151 B.n150 10.6151
R1181 B.n151 B.n118 10.6151
R1182 B.n155 B.n118 10.6151
R1183 B.n156 B.n155 10.6151
R1184 B.n157 B.n156 10.6151
R1185 B.n157 B.n116 10.6151
R1186 B.n161 B.n116 10.6151
R1187 B.n162 B.n161 10.6151
R1188 B.n163 B.n162 10.6151
R1189 B.n167 B.n114 10.6151
R1190 B.n168 B.n167 10.6151
R1191 B.n169 B.n168 10.6151
R1192 B.n169 B.n112 10.6151
R1193 B.n173 B.n112 10.6151
R1194 B.n174 B.n173 10.6151
R1195 B.n175 B.n174 10.6151
R1196 B.n175 B.n110 10.6151
R1197 B.n179 B.n110 10.6151
R1198 B.n180 B.n179 10.6151
R1199 B.n181 B.n180 10.6151
R1200 B.n181 B.n108 10.6151
R1201 B.n185 B.n108 10.6151
R1202 B.n186 B.n185 10.6151
R1203 B.n187 B.n186 10.6151
R1204 B.n187 B.n106 10.6151
R1205 B.n191 B.n106 10.6151
R1206 B.n192 B.n191 10.6151
R1207 B.n193 B.n192 10.6151
R1208 B.n193 B.n104 10.6151
R1209 B.n197 B.n104 10.6151
R1210 B.n198 B.n197 10.6151
R1211 B.n199 B.n198 10.6151
R1212 B.n199 B.n102 10.6151
R1213 B.n203 B.n102 10.6151
R1214 B.n204 B.n203 10.6151
R1215 B.n208 B.n204 10.6151
R1216 B.n212 B.n100 10.6151
R1217 B.n213 B.n212 10.6151
R1218 B.n214 B.n213 10.6151
R1219 B.n214 B.n98 10.6151
R1220 B.n218 B.n98 10.6151
R1221 B.n219 B.n218 10.6151
R1222 B.n220 B.n219 10.6151
R1223 B.n220 B.n96 10.6151
R1224 B.n224 B.n96 10.6151
R1225 B.n227 B.n226 10.6151
R1226 B.n227 B.n92 10.6151
R1227 B.n231 B.n92 10.6151
R1228 B.n232 B.n231 10.6151
R1229 B.n233 B.n232 10.6151
R1230 B.n233 B.n90 10.6151
R1231 B.n237 B.n90 10.6151
R1232 B.n238 B.n237 10.6151
R1233 B.n239 B.n238 10.6151
R1234 B.n239 B.n88 10.6151
R1235 B.n243 B.n88 10.6151
R1236 B.n244 B.n243 10.6151
R1237 B.n245 B.n244 10.6151
R1238 B.n245 B.n86 10.6151
R1239 B.n249 B.n86 10.6151
R1240 B.n250 B.n249 10.6151
R1241 B.n251 B.n250 10.6151
R1242 B.n251 B.n84 10.6151
R1243 B.n255 B.n84 10.6151
R1244 B.n256 B.n255 10.6151
R1245 B.n257 B.n256 10.6151
R1246 B.n257 B.n82 10.6151
R1247 B.n261 B.n82 10.6151
R1248 B.n262 B.n261 10.6151
R1249 B.n263 B.n262 10.6151
R1250 B.n263 B.n80 10.6151
R1251 B.n267 B.n80 10.6151
R1252 B.n407 B.n406 9.36635
R1253 B.n389 B.n38 9.36635
R1254 B.n208 B.n207 9.36635
R1255 B.n226 B.n225 9.36635
R1256 B.n489 B.n0 8.11757
R1257 B.n489 B.n1 8.11757
R1258 B.n406 B.n405 1.24928
R1259 B.n392 B.n38 1.24928
R1260 B.n207 B.n100 1.24928
R1261 B.n225 B.n224 1.24928
R1262 VN.n0 VN.t2 137.567
R1263 VN.n1 VN.t3 137.567
R1264 VN.n0 VN.t1 137.142
R1265 VN.n1 VN.t0 137.142
R1266 VN VN.n1 49.9058
R1267 VN VN.n0 9.43984
R1268 VDD2.n2 VDD2.n0 119.797
R1269 VDD2.n2 VDD2.n1 84.3327
R1270 VDD2.n1 VDD2.t3 4.39901
R1271 VDD2.n1 VDD2.t0 4.39901
R1272 VDD2.n0 VDD2.t1 4.39901
R1273 VDD2.n0 VDD2.t2 4.39901
R1274 VDD2 VDD2.n2 0.0586897
C0 VN w_n2218_n2446# 3.51868f
C1 VP w_n2218_n2446# 3.80166f
C2 VDD2 B 1.02653f
C3 VDD1 VDD2 0.819364f
C4 VDD1 B 0.988279f
C5 VTAIL VDD2 4.18398f
C6 VTAIL B 3.09892f
C7 VTAIL VDD1 4.13547f
C8 VN VDD2 2.80709f
C9 VN B 0.893319f
C10 VN VDD1 0.148053f
C11 VP VDD2 0.340039f
C12 VP B 1.35896f
C13 VTAIL VN 2.78542f
C14 VP VDD1 2.99855f
C15 VDD2 w_n2218_n2446# 1.19698f
C16 VTAIL VP 2.79952f
C17 B w_n2218_n2446# 6.90769f
C18 VDD1 w_n2218_n2446# 1.15987f
C19 VN VP 4.72588f
C20 VTAIL w_n2218_n2446# 2.90535f
C21 VDD2 VSUBS 0.703122f
C22 VDD1 VSUBS 4.626422f
C23 VTAIL VSUBS 0.873432f
C24 VN VSUBS 4.99239f
C25 VP VSUBS 1.651835f
C26 B VSUBS 3.15089f
C27 w_n2218_n2446# VSUBS 67.4183f
C28 VDD2.t1 VSUBS 0.157721f
C29 VDD2.t2 VSUBS 0.157721f
C30 VDD2.n0 VSUBS 1.56578f
C31 VDD2.t3 VSUBS 0.157721f
C32 VDD2.t0 VSUBS 0.157721f
C33 VDD2.n1 VSUBS 1.10132f
C34 VDD2.n2 VSUBS 3.54016f
C35 VN.t2 VSUBS 1.77589f
C36 VN.t1 VSUBS 1.77338f
C37 VN.n0 VSUBS 1.27154f
C38 VN.t3 VSUBS 1.77589f
C39 VN.t0 VSUBS 1.77338f
C40 VN.n1 VSUBS 2.94116f
C41 B.n0 VSUBS 0.007223f
C42 B.n1 VSUBS 0.007223f
C43 B.n2 VSUBS 0.010682f
C44 B.n3 VSUBS 0.008186f
C45 B.n4 VSUBS 0.008186f
C46 B.n5 VSUBS 0.008186f
C47 B.n6 VSUBS 0.008186f
C48 B.n7 VSUBS 0.008186f
C49 B.n8 VSUBS 0.008186f
C50 B.n9 VSUBS 0.008186f
C51 B.n10 VSUBS 0.008186f
C52 B.n11 VSUBS 0.008186f
C53 B.n12 VSUBS 0.008186f
C54 B.n13 VSUBS 0.008186f
C55 B.n14 VSUBS 0.008186f
C56 B.n15 VSUBS 0.018892f
C57 B.n16 VSUBS 0.008186f
C58 B.n17 VSUBS 0.008186f
C59 B.n18 VSUBS 0.008186f
C60 B.n19 VSUBS 0.008186f
C61 B.n20 VSUBS 0.008186f
C62 B.n21 VSUBS 0.008186f
C63 B.n22 VSUBS 0.008186f
C64 B.n23 VSUBS 0.008186f
C65 B.n24 VSUBS 0.008186f
C66 B.n25 VSUBS 0.008186f
C67 B.n26 VSUBS 0.008186f
C68 B.n27 VSUBS 0.008186f
C69 B.n28 VSUBS 0.008186f
C70 B.n29 VSUBS 0.008186f
C71 B.t4 VSUBS 0.134431f
C72 B.t5 VSUBS 0.158174f
C73 B.t3 VSUBS 0.691056f
C74 B.n30 VSUBS 0.267275f
C75 B.n31 VSUBS 0.207801f
C76 B.n32 VSUBS 0.008186f
C77 B.n33 VSUBS 0.008186f
C78 B.n34 VSUBS 0.008186f
C79 B.n35 VSUBS 0.008186f
C80 B.t10 VSUBS 0.134434f
C81 B.t11 VSUBS 0.158177f
C82 B.t9 VSUBS 0.691056f
C83 B.n36 VSUBS 0.267273f
C84 B.n37 VSUBS 0.207799f
C85 B.n38 VSUBS 0.018965f
C86 B.n39 VSUBS 0.008186f
C87 B.n40 VSUBS 0.008186f
C88 B.n41 VSUBS 0.008186f
C89 B.n42 VSUBS 0.008186f
C90 B.n43 VSUBS 0.008186f
C91 B.n44 VSUBS 0.008186f
C92 B.n45 VSUBS 0.008186f
C93 B.n46 VSUBS 0.008186f
C94 B.n47 VSUBS 0.008186f
C95 B.n48 VSUBS 0.008186f
C96 B.n49 VSUBS 0.008186f
C97 B.n50 VSUBS 0.008186f
C98 B.n51 VSUBS 0.008186f
C99 B.n52 VSUBS 0.018892f
C100 B.n53 VSUBS 0.008186f
C101 B.n54 VSUBS 0.008186f
C102 B.n55 VSUBS 0.008186f
C103 B.n56 VSUBS 0.008186f
C104 B.n57 VSUBS 0.008186f
C105 B.n58 VSUBS 0.008186f
C106 B.n59 VSUBS 0.008186f
C107 B.n60 VSUBS 0.008186f
C108 B.n61 VSUBS 0.008186f
C109 B.n62 VSUBS 0.008186f
C110 B.n63 VSUBS 0.008186f
C111 B.n64 VSUBS 0.008186f
C112 B.n65 VSUBS 0.008186f
C113 B.n66 VSUBS 0.008186f
C114 B.n67 VSUBS 0.008186f
C115 B.n68 VSUBS 0.008186f
C116 B.n69 VSUBS 0.008186f
C117 B.n70 VSUBS 0.008186f
C118 B.n71 VSUBS 0.008186f
C119 B.n72 VSUBS 0.008186f
C120 B.n73 VSUBS 0.008186f
C121 B.n74 VSUBS 0.008186f
C122 B.n75 VSUBS 0.008186f
C123 B.n76 VSUBS 0.008186f
C124 B.n77 VSUBS 0.008186f
C125 B.n78 VSUBS 0.008186f
C126 B.n79 VSUBS 0.017702f
C127 B.n80 VSUBS 0.008186f
C128 B.n81 VSUBS 0.008186f
C129 B.n82 VSUBS 0.008186f
C130 B.n83 VSUBS 0.008186f
C131 B.n84 VSUBS 0.008186f
C132 B.n85 VSUBS 0.008186f
C133 B.n86 VSUBS 0.008186f
C134 B.n87 VSUBS 0.008186f
C135 B.n88 VSUBS 0.008186f
C136 B.n89 VSUBS 0.008186f
C137 B.n90 VSUBS 0.008186f
C138 B.n91 VSUBS 0.008186f
C139 B.n92 VSUBS 0.008186f
C140 B.n93 VSUBS 0.008186f
C141 B.t2 VSUBS 0.134434f
C142 B.t1 VSUBS 0.158177f
C143 B.t0 VSUBS 0.691056f
C144 B.n94 VSUBS 0.267273f
C145 B.n95 VSUBS 0.207799f
C146 B.n96 VSUBS 0.008186f
C147 B.n97 VSUBS 0.008186f
C148 B.n98 VSUBS 0.008186f
C149 B.n99 VSUBS 0.008186f
C150 B.n100 VSUBS 0.004574f
C151 B.n101 VSUBS 0.008186f
C152 B.n102 VSUBS 0.008186f
C153 B.n103 VSUBS 0.008186f
C154 B.n104 VSUBS 0.008186f
C155 B.n105 VSUBS 0.008186f
C156 B.n106 VSUBS 0.008186f
C157 B.n107 VSUBS 0.008186f
C158 B.n108 VSUBS 0.008186f
C159 B.n109 VSUBS 0.008186f
C160 B.n110 VSUBS 0.008186f
C161 B.n111 VSUBS 0.008186f
C162 B.n112 VSUBS 0.008186f
C163 B.n113 VSUBS 0.008186f
C164 B.n114 VSUBS 0.018892f
C165 B.n115 VSUBS 0.008186f
C166 B.n116 VSUBS 0.008186f
C167 B.n117 VSUBS 0.008186f
C168 B.n118 VSUBS 0.008186f
C169 B.n119 VSUBS 0.008186f
C170 B.n120 VSUBS 0.008186f
C171 B.n121 VSUBS 0.008186f
C172 B.n122 VSUBS 0.008186f
C173 B.n123 VSUBS 0.008186f
C174 B.n124 VSUBS 0.008186f
C175 B.n125 VSUBS 0.008186f
C176 B.n126 VSUBS 0.008186f
C177 B.n127 VSUBS 0.008186f
C178 B.n128 VSUBS 0.008186f
C179 B.n129 VSUBS 0.008186f
C180 B.n130 VSUBS 0.008186f
C181 B.n131 VSUBS 0.008186f
C182 B.n132 VSUBS 0.008186f
C183 B.n133 VSUBS 0.008186f
C184 B.n134 VSUBS 0.008186f
C185 B.n135 VSUBS 0.008186f
C186 B.n136 VSUBS 0.008186f
C187 B.n137 VSUBS 0.008186f
C188 B.n138 VSUBS 0.008186f
C189 B.n139 VSUBS 0.008186f
C190 B.n140 VSUBS 0.008186f
C191 B.n141 VSUBS 0.008186f
C192 B.n142 VSUBS 0.008186f
C193 B.n143 VSUBS 0.008186f
C194 B.n144 VSUBS 0.008186f
C195 B.n145 VSUBS 0.008186f
C196 B.n146 VSUBS 0.008186f
C197 B.n147 VSUBS 0.008186f
C198 B.n148 VSUBS 0.008186f
C199 B.n149 VSUBS 0.008186f
C200 B.n150 VSUBS 0.008186f
C201 B.n151 VSUBS 0.008186f
C202 B.n152 VSUBS 0.008186f
C203 B.n153 VSUBS 0.008186f
C204 B.n154 VSUBS 0.008186f
C205 B.n155 VSUBS 0.008186f
C206 B.n156 VSUBS 0.008186f
C207 B.n157 VSUBS 0.008186f
C208 B.n158 VSUBS 0.008186f
C209 B.n159 VSUBS 0.008186f
C210 B.n160 VSUBS 0.008186f
C211 B.n161 VSUBS 0.008186f
C212 B.n162 VSUBS 0.008186f
C213 B.n163 VSUBS 0.017702f
C214 B.n164 VSUBS 0.017702f
C215 B.n165 VSUBS 0.018892f
C216 B.n166 VSUBS 0.008186f
C217 B.n167 VSUBS 0.008186f
C218 B.n168 VSUBS 0.008186f
C219 B.n169 VSUBS 0.008186f
C220 B.n170 VSUBS 0.008186f
C221 B.n171 VSUBS 0.008186f
C222 B.n172 VSUBS 0.008186f
C223 B.n173 VSUBS 0.008186f
C224 B.n174 VSUBS 0.008186f
C225 B.n175 VSUBS 0.008186f
C226 B.n176 VSUBS 0.008186f
C227 B.n177 VSUBS 0.008186f
C228 B.n178 VSUBS 0.008186f
C229 B.n179 VSUBS 0.008186f
C230 B.n180 VSUBS 0.008186f
C231 B.n181 VSUBS 0.008186f
C232 B.n182 VSUBS 0.008186f
C233 B.n183 VSUBS 0.008186f
C234 B.n184 VSUBS 0.008186f
C235 B.n185 VSUBS 0.008186f
C236 B.n186 VSUBS 0.008186f
C237 B.n187 VSUBS 0.008186f
C238 B.n188 VSUBS 0.008186f
C239 B.n189 VSUBS 0.008186f
C240 B.n190 VSUBS 0.008186f
C241 B.n191 VSUBS 0.008186f
C242 B.n192 VSUBS 0.008186f
C243 B.n193 VSUBS 0.008186f
C244 B.n194 VSUBS 0.008186f
C245 B.n195 VSUBS 0.008186f
C246 B.n196 VSUBS 0.008186f
C247 B.n197 VSUBS 0.008186f
C248 B.n198 VSUBS 0.008186f
C249 B.n199 VSUBS 0.008186f
C250 B.n200 VSUBS 0.008186f
C251 B.n201 VSUBS 0.008186f
C252 B.n202 VSUBS 0.008186f
C253 B.n203 VSUBS 0.008186f
C254 B.n204 VSUBS 0.008186f
C255 B.t8 VSUBS 0.134431f
C256 B.t7 VSUBS 0.158174f
C257 B.t6 VSUBS 0.691056f
C258 B.n205 VSUBS 0.267275f
C259 B.n206 VSUBS 0.207801f
C260 B.n207 VSUBS 0.018965f
C261 B.n208 VSUBS 0.007704f
C262 B.n209 VSUBS 0.008186f
C263 B.n210 VSUBS 0.008186f
C264 B.n211 VSUBS 0.008186f
C265 B.n212 VSUBS 0.008186f
C266 B.n213 VSUBS 0.008186f
C267 B.n214 VSUBS 0.008186f
C268 B.n215 VSUBS 0.008186f
C269 B.n216 VSUBS 0.008186f
C270 B.n217 VSUBS 0.008186f
C271 B.n218 VSUBS 0.008186f
C272 B.n219 VSUBS 0.008186f
C273 B.n220 VSUBS 0.008186f
C274 B.n221 VSUBS 0.008186f
C275 B.n222 VSUBS 0.008186f
C276 B.n223 VSUBS 0.008186f
C277 B.n224 VSUBS 0.004574f
C278 B.n225 VSUBS 0.018965f
C279 B.n226 VSUBS 0.007704f
C280 B.n227 VSUBS 0.008186f
C281 B.n228 VSUBS 0.008186f
C282 B.n229 VSUBS 0.008186f
C283 B.n230 VSUBS 0.008186f
C284 B.n231 VSUBS 0.008186f
C285 B.n232 VSUBS 0.008186f
C286 B.n233 VSUBS 0.008186f
C287 B.n234 VSUBS 0.008186f
C288 B.n235 VSUBS 0.008186f
C289 B.n236 VSUBS 0.008186f
C290 B.n237 VSUBS 0.008186f
C291 B.n238 VSUBS 0.008186f
C292 B.n239 VSUBS 0.008186f
C293 B.n240 VSUBS 0.008186f
C294 B.n241 VSUBS 0.008186f
C295 B.n242 VSUBS 0.008186f
C296 B.n243 VSUBS 0.008186f
C297 B.n244 VSUBS 0.008186f
C298 B.n245 VSUBS 0.008186f
C299 B.n246 VSUBS 0.008186f
C300 B.n247 VSUBS 0.008186f
C301 B.n248 VSUBS 0.008186f
C302 B.n249 VSUBS 0.008186f
C303 B.n250 VSUBS 0.008186f
C304 B.n251 VSUBS 0.008186f
C305 B.n252 VSUBS 0.008186f
C306 B.n253 VSUBS 0.008186f
C307 B.n254 VSUBS 0.008186f
C308 B.n255 VSUBS 0.008186f
C309 B.n256 VSUBS 0.008186f
C310 B.n257 VSUBS 0.008186f
C311 B.n258 VSUBS 0.008186f
C312 B.n259 VSUBS 0.008186f
C313 B.n260 VSUBS 0.008186f
C314 B.n261 VSUBS 0.008186f
C315 B.n262 VSUBS 0.008186f
C316 B.n263 VSUBS 0.008186f
C317 B.n264 VSUBS 0.008186f
C318 B.n265 VSUBS 0.008186f
C319 B.n266 VSUBS 0.018892f
C320 B.n267 VSUBS 0.017854f
C321 B.n268 VSUBS 0.01874f
C322 B.n269 VSUBS 0.008186f
C323 B.n270 VSUBS 0.008186f
C324 B.n271 VSUBS 0.008186f
C325 B.n272 VSUBS 0.008186f
C326 B.n273 VSUBS 0.008186f
C327 B.n274 VSUBS 0.008186f
C328 B.n275 VSUBS 0.008186f
C329 B.n276 VSUBS 0.008186f
C330 B.n277 VSUBS 0.008186f
C331 B.n278 VSUBS 0.008186f
C332 B.n279 VSUBS 0.008186f
C333 B.n280 VSUBS 0.008186f
C334 B.n281 VSUBS 0.008186f
C335 B.n282 VSUBS 0.008186f
C336 B.n283 VSUBS 0.008186f
C337 B.n284 VSUBS 0.008186f
C338 B.n285 VSUBS 0.008186f
C339 B.n286 VSUBS 0.008186f
C340 B.n287 VSUBS 0.008186f
C341 B.n288 VSUBS 0.008186f
C342 B.n289 VSUBS 0.008186f
C343 B.n290 VSUBS 0.008186f
C344 B.n291 VSUBS 0.008186f
C345 B.n292 VSUBS 0.008186f
C346 B.n293 VSUBS 0.008186f
C347 B.n294 VSUBS 0.008186f
C348 B.n295 VSUBS 0.008186f
C349 B.n296 VSUBS 0.008186f
C350 B.n297 VSUBS 0.008186f
C351 B.n298 VSUBS 0.008186f
C352 B.n299 VSUBS 0.008186f
C353 B.n300 VSUBS 0.008186f
C354 B.n301 VSUBS 0.008186f
C355 B.n302 VSUBS 0.008186f
C356 B.n303 VSUBS 0.008186f
C357 B.n304 VSUBS 0.008186f
C358 B.n305 VSUBS 0.008186f
C359 B.n306 VSUBS 0.008186f
C360 B.n307 VSUBS 0.008186f
C361 B.n308 VSUBS 0.008186f
C362 B.n309 VSUBS 0.008186f
C363 B.n310 VSUBS 0.008186f
C364 B.n311 VSUBS 0.008186f
C365 B.n312 VSUBS 0.008186f
C366 B.n313 VSUBS 0.008186f
C367 B.n314 VSUBS 0.008186f
C368 B.n315 VSUBS 0.008186f
C369 B.n316 VSUBS 0.008186f
C370 B.n317 VSUBS 0.008186f
C371 B.n318 VSUBS 0.008186f
C372 B.n319 VSUBS 0.008186f
C373 B.n320 VSUBS 0.008186f
C374 B.n321 VSUBS 0.008186f
C375 B.n322 VSUBS 0.008186f
C376 B.n323 VSUBS 0.008186f
C377 B.n324 VSUBS 0.008186f
C378 B.n325 VSUBS 0.008186f
C379 B.n326 VSUBS 0.008186f
C380 B.n327 VSUBS 0.008186f
C381 B.n328 VSUBS 0.008186f
C382 B.n329 VSUBS 0.008186f
C383 B.n330 VSUBS 0.008186f
C384 B.n331 VSUBS 0.008186f
C385 B.n332 VSUBS 0.008186f
C386 B.n333 VSUBS 0.008186f
C387 B.n334 VSUBS 0.008186f
C388 B.n335 VSUBS 0.008186f
C389 B.n336 VSUBS 0.008186f
C390 B.n337 VSUBS 0.008186f
C391 B.n338 VSUBS 0.008186f
C392 B.n339 VSUBS 0.008186f
C393 B.n340 VSUBS 0.008186f
C394 B.n341 VSUBS 0.008186f
C395 B.n342 VSUBS 0.008186f
C396 B.n343 VSUBS 0.008186f
C397 B.n344 VSUBS 0.008186f
C398 B.n345 VSUBS 0.008186f
C399 B.n346 VSUBS 0.008186f
C400 B.n347 VSUBS 0.017702f
C401 B.n348 VSUBS 0.017702f
C402 B.n349 VSUBS 0.018892f
C403 B.n350 VSUBS 0.008186f
C404 B.n351 VSUBS 0.008186f
C405 B.n352 VSUBS 0.008186f
C406 B.n353 VSUBS 0.008186f
C407 B.n354 VSUBS 0.008186f
C408 B.n355 VSUBS 0.008186f
C409 B.n356 VSUBS 0.008186f
C410 B.n357 VSUBS 0.008186f
C411 B.n358 VSUBS 0.008186f
C412 B.n359 VSUBS 0.008186f
C413 B.n360 VSUBS 0.008186f
C414 B.n361 VSUBS 0.008186f
C415 B.n362 VSUBS 0.008186f
C416 B.n363 VSUBS 0.008186f
C417 B.n364 VSUBS 0.008186f
C418 B.n365 VSUBS 0.008186f
C419 B.n366 VSUBS 0.008186f
C420 B.n367 VSUBS 0.008186f
C421 B.n368 VSUBS 0.008186f
C422 B.n369 VSUBS 0.008186f
C423 B.n370 VSUBS 0.008186f
C424 B.n371 VSUBS 0.008186f
C425 B.n372 VSUBS 0.008186f
C426 B.n373 VSUBS 0.008186f
C427 B.n374 VSUBS 0.008186f
C428 B.n375 VSUBS 0.008186f
C429 B.n376 VSUBS 0.008186f
C430 B.n377 VSUBS 0.008186f
C431 B.n378 VSUBS 0.008186f
C432 B.n379 VSUBS 0.008186f
C433 B.n380 VSUBS 0.008186f
C434 B.n381 VSUBS 0.008186f
C435 B.n382 VSUBS 0.008186f
C436 B.n383 VSUBS 0.008186f
C437 B.n384 VSUBS 0.008186f
C438 B.n385 VSUBS 0.008186f
C439 B.n386 VSUBS 0.008186f
C440 B.n387 VSUBS 0.008186f
C441 B.n388 VSUBS 0.008186f
C442 B.n389 VSUBS 0.007704f
C443 B.n390 VSUBS 0.008186f
C444 B.n391 VSUBS 0.008186f
C445 B.n392 VSUBS 0.004574f
C446 B.n393 VSUBS 0.008186f
C447 B.n394 VSUBS 0.008186f
C448 B.n395 VSUBS 0.008186f
C449 B.n396 VSUBS 0.008186f
C450 B.n397 VSUBS 0.008186f
C451 B.n398 VSUBS 0.008186f
C452 B.n399 VSUBS 0.008186f
C453 B.n400 VSUBS 0.008186f
C454 B.n401 VSUBS 0.008186f
C455 B.n402 VSUBS 0.008186f
C456 B.n403 VSUBS 0.008186f
C457 B.n404 VSUBS 0.008186f
C458 B.n405 VSUBS 0.004574f
C459 B.n406 VSUBS 0.018965f
C460 B.n407 VSUBS 0.007704f
C461 B.n408 VSUBS 0.008186f
C462 B.n409 VSUBS 0.008186f
C463 B.n410 VSUBS 0.008186f
C464 B.n411 VSUBS 0.008186f
C465 B.n412 VSUBS 0.008186f
C466 B.n413 VSUBS 0.008186f
C467 B.n414 VSUBS 0.008186f
C468 B.n415 VSUBS 0.008186f
C469 B.n416 VSUBS 0.008186f
C470 B.n417 VSUBS 0.008186f
C471 B.n418 VSUBS 0.008186f
C472 B.n419 VSUBS 0.008186f
C473 B.n420 VSUBS 0.008186f
C474 B.n421 VSUBS 0.008186f
C475 B.n422 VSUBS 0.008186f
C476 B.n423 VSUBS 0.008186f
C477 B.n424 VSUBS 0.008186f
C478 B.n425 VSUBS 0.008186f
C479 B.n426 VSUBS 0.008186f
C480 B.n427 VSUBS 0.008186f
C481 B.n428 VSUBS 0.008186f
C482 B.n429 VSUBS 0.008186f
C483 B.n430 VSUBS 0.008186f
C484 B.n431 VSUBS 0.008186f
C485 B.n432 VSUBS 0.008186f
C486 B.n433 VSUBS 0.008186f
C487 B.n434 VSUBS 0.008186f
C488 B.n435 VSUBS 0.008186f
C489 B.n436 VSUBS 0.008186f
C490 B.n437 VSUBS 0.008186f
C491 B.n438 VSUBS 0.008186f
C492 B.n439 VSUBS 0.008186f
C493 B.n440 VSUBS 0.008186f
C494 B.n441 VSUBS 0.008186f
C495 B.n442 VSUBS 0.008186f
C496 B.n443 VSUBS 0.008186f
C497 B.n444 VSUBS 0.008186f
C498 B.n445 VSUBS 0.008186f
C499 B.n446 VSUBS 0.008186f
C500 B.n447 VSUBS 0.008186f
C501 B.n448 VSUBS 0.018892f
C502 B.n449 VSUBS 0.017702f
C503 B.n450 VSUBS 0.017702f
C504 B.n451 VSUBS 0.008186f
C505 B.n452 VSUBS 0.008186f
C506 B.n453 VSUBS 0.008186f
C507 B.n454 VSUBS 0.008186f
C508 B.n455 VSUBS 0.008186f
C509 B.n456 VSUBS 0.008186f
C510 B.n457 VSUBS 0.008186f
C511 B.n458 VSUBS 0.008186f
C512 B.n459 VSUBS 0.008186f
C513 B.n460 VSUBS 0.008186f
C514 B.n461 VSUBS 0.008186f
C515 B.n462 VSUBS 0.008186f
C516 B.n463 VSUBS 0.008186f
C517 B.n464 VSUBS 0.008186f
C518 B.n465 VSUBS 0.008186f
C519 B.n466 VSUBS 0.008186f
C520 B.n467 VSUBS 0.008186f
C521 B.n468 VSUBS 0.008186f
C522 B.n469 VSUBS 0.008186f
C523 B.n470 VSUBS 0.008186f
C524 B.n471 VSUBS 0.008186f
C525 B.n472 VSUBS 0.008186f
C526 B.n473 VSUBS 0.008186f
C527 B.n474 VSUBS 0.008186f
C528 B.n475 VSUBS 0.008186f
C529 B.n476 VSUBS 0.008186f
C530 B.n477 VSUBS 0.008186f
C531 B.n478 VSUBS 0.008186f
C532 B.n479 VSUBS 0.008186f
C533 B.n480 VSUBS 0.008186f
C534 B.n481 VSUBS 0.008186f
C535 B.n482 VSUBS 0.008186f
C536 B.n483 VSUBS 0.008186f
C537 B.n484 VSUBS 0.008186f
C538 B.n485 VSUBS 0.008186f
C539 B.n486 VSUBS 0.008186f
C540 B.n487 VSUBS 0.010682f
C541 B.n488 VSUBS 0.011379f
C542 B.n489 VSUBS 0.022628f
C543 VDD1.t2 VSUBS 0.157726f
C544 VDD1.t3 VSUBS 0.157726f
C545 VDD1.n0 VSUBS 1.1018f
C546 VDD1.t0 VSUBS 0.157726f
C547 VDD1.t1 VSUBS 0.157726f
C548 VDD1.n1 VSUBS 1.58701f
C549 VTAIL.n0 VSUBS 0.027778f
C550 VTAIL.n1 VSUBS 0.025086f
C551 VTAIL.n2 VSUBS 0.01348f
C552 VTAIL.n3 VSUBS 0.031862f
C553 VTAIL.n4 VSUBS 0.014273f
C554 VTAIL.n5 VSUBS 0.025086f
C555 VTAIL.n6 VSUBS 0.01348f
C556 VTAIL.n7 VSUBS 0.031862f
C557 VTAIL.n8 VSUBS 0.014273f
C558 VTAIL.n9 VSUBS 0.025086f
C559 VTAIL.n10 VSUBS 0.01348f
C560 VTAIL.n11 VSUBS 0.023897f
C561 VTAIL.n12 VSUBS 0.020268f
C562 VTAIL.t1 VSUBS 0.068005f
C563 VTAIL.n13 VSUBS 0.12079f
C564 VTAIL.n14 VSUBS 0.734614f
C565 VTAIL.n15 VSUBS 0.01348f
C566 VTAIL.n16 VSUBS 0.014273f
C567 VTAIL.n17 VSUBS 0.031862f
C568 VTAIL.n18 VSUBS 0.031862f
C569 VTAIL.n19 VSUBS 0.014273f
C570 VTAIL.n20 VSUBS 0.01348f
C571 VTAIL.n21 VSUBS 0.025086f
C572 VTAIL.n22 VSUBS 0.025086f
C573 VTAIL.n23 VSUBS 0.01348f
C574 VTAIL.n24 VSUBS 0.014273f
C575 VTAIL.n25 VSUBS 0.031862f
C576 VTAIL.n26 VSUBS 0.031862f
C577 VTAIL.n27 VSUBS 0.014273f
C578 VTAIL.n28 VSUBS 0.01348f
C579 VTAIL.n29 VSUBS 0.025086f
C580 VTAIL.n30 VSUBS 0.025086f
C581 VTAIL.n31 VSUBS 0.01348f
C582 VTAIL.n32 VSUBS 0.014273f
C583 VTAIL.n33 VSUBS 0.031862f
C584 VTAIL.n34 VSUBS 0.077865f
C585 VTAIL.n35 VSUBS 0.014273f
C586 VTAIL.n36 VSUBS 0.01348f
C587 VTAIL.n37 VSUBS 0.056272f
C588 VTAIL.n38 VSUBS 0.039136f
C589 VTAIL.n39 VSUBS 0.135612f
C590 VTAIL.n40 VSUBS 0.027778f
C591 VTAIL.n41 VSUBS 0.025086f
C592 VTAIL.n42 VSUBS 0.01348f
C593 VTAIL.n43 VSUBS 0.031862f
C594 VTAIL.n44 VSUBS 0.014273f
C595 VTAIL.n45 VSUBS 0.025086f
C596 VTAIL.n46 VSUBS 0.01348f
C597 VTAIL.n47 VSUBS 0.031862f
C598 VTAIL.n48 VSUBS 0.014273f
C599 VTAIL.n49 VSUBS 0.025086f
C600 VTAIL.n50 VSUBS 0.01348f
C601 VTAIL.n51 VSUBS 0.023897f
C602 VTAIL.n52 VSUBS 0.020268f
C603 VTAIL.t6 VSUBS 0.068005f
C604 VTAIL.n53 VSUBS 0.12079f
C605 VTAIL.n54 VSUBS 0.734614f
C606 VTAIL.n55 VSUBS 0.01348f
C607 VTAIL.n56 VSUBS 0.014273f
C608 VTAIL.n57 VSUBS 0.031862f
C609 VTAIL.n58 VSUBS 0.031862f
C610 VTAIL.n59 VSUBS 0.014273f
C611 VTAIL.n60 VSUBS 0.01348f
C612 VTAIL.n61 VSUBS 0.025086f
C613 VTAIL.n62 VSUBS 0.025086f
C614 VTAIL.n63 VSUBS 0.01348f
C615 VTAIL.n64 VSUBS 0.014273f
C616 VTAIL.n65 VSUBS 0.031862f
C617 VTAIL.n66 VSUBS 0.031862f
C618 VTAIL.n67 VSUBS 0.014273f
C619 VTAIL.n68 VSUBS 0.01348f
C620 VTAIL.n69 VSUBS 0.025086f
C621 VTAIL.n70 VSUBS 0.025086f
C622 VTAIL.n71 VSUBS 0.01348f
C623 VTAIL.n72 VSUBS 0.014273f
C624 VTAIL.n73 VSUBS 0.031862f
C625 VTAIL.n74 VSUBS 0.077865f
C626 VTAIL.n75 VSUBS 0.014273f
C627 VTAIL.n76 VSUBS 0.01348f
C628 VTAIL.n77 VSUBS 0.056272f
C629 VTAIL.n78 VSUBS 0.039136f
C630 VTAIL.n79 VSUBS 0.203379f
C631 VTAIL.n80 VSUBS 0.027778f
C632 VTAIL.n81 VSUBS 0.025086f
C633 VTAIL.n82 VSUBS 0.01348f
C634 VTAIL.n83 VSUBS 0.031862f
C635 VTAIL.n84 VSUBS 0.014273f
C636 VTAIL.n85 VSUBS 0.025086f
C637 VTAIL.n86 VSUBS 0.01348f
C638 VTAIL.n87 VSUBS 0.031862f
C639 VTAIL.n88 VSUBS 0.014273f
C640 VTAIL.n89 VSUBS 0.025086f
C641 VTAIL.n90 VSUBS 0.01348f
C642 VTAIL.n91 VSUBS 0.023897f
C643 VTAIL.n92 VSUBS 0.020268f
C644 VTAIL.t7 VSUBS 0.068005f
C645 VTAIL.n93 VSUBS 0.12079f
C646 VTAIL.n94 VSUBS 0.734614f
C647 VTAIL.n95 VSUBS 0.01348f
C648 VTAIL.n96 VSUBS 0.014273f
C649 VTAIL.n97 VSUBS 0.031862f
C650 VTAIL.n98 VSUBS 0.031862f
C651 VTAIL.n99 VSUBS 0.014273f
C652 VTAIL.n100 VSUBS 0.01348f
C653 VTAIL.n101 VSUBS 0.025086f
C654 VTAIL.n102 VSUBS 0.025086f
C655 VTAIL.n103 VSUBS 0.01348f
C656 VTAIL.n104 VSUBS 0.014273f
C657 VTAIL.n105 VSUBS 0.031862f
C658 VTAIL.n106 VSUBS 0.031862f
C659 VTAIL.n107 VSUBS 0.014273f
C660 VTAIL.n108 VSUBS 0.01348f
C661 VTAIL.n109 VSUBS 0.025086f
C662 VTAIL.n110 VSUBS 0.025086f
C663 VTAIL.n111 VSUBS 0.01348f
C664 VTAIL.n112 VSUBS 0.014273f
C665 VTAIL.n113 VSUBS 0.031862f
C666 VTAIL.n114 VSUBS 0.077865f
C667 VTAIL.n115 VSUBS 0.014273f
C668 VTAIL.n116 VSUBS 0.01348f
C669 VTAIL.n117 VSUBS 0.056272f
C670 VTAIL.n118 VSUBS 0.039136f
C671 VTAIL.n119 VSUBS 1.16607f
C672 VTAIL.n120 VSUBS 0.027778f
C673 VTAIL.n121 VSUBS 0.025086f
C674 VTAIL.n122 VSUBS 0.01348f
C675 VTAIL.n123 VSUBS 0.031862f
C676 VTAIL.n124 VSUBS 0.014273f
C677 VTAIL.n125 VSUBS 0.025086f
C678 VTAIL.n126 VSUBS 0.01348f
C679 VTAIL.n127 VSUBS 0.031862f
C680 VTAIL.n128 VSUBS 0.014273f
C681 VTAIL.n129 VSUBS 0.025086f
C682 VTAIL.n130 VSUBS 0.01348f
C683 VTAIL.n131 VSUBS 0.023897f
C684 VTAIL.n132 VSUBS 0.020268f
C685 VTAIL.t0 VSUBS 0.068005f
C686 VTAIL.n133 VSUBS 0.12079f
C687 VTAIL.n134 VSUBS 0.734614f
C688 VTAIL.n135 VSUBS 0.01348f
C689 VTAIL.n136 VSUBS 0.014273f
C690 VTAIL.n137 VSUBS 0.031862f
C691 VTAIL.n138 VSUBS 0.031862f
C692 VTAIL.n139 VSUBS 0.014273f
C693 VTAIL.n140 VSUBS 0.01348f
C694 VTAIL.n141 VSUBS 0.025086f
C695 VTAIL.n142 VSUBS 0.025086f
C696 VTAIL.n143 VSUBS 0.01348f
C697 VTAIL.n144 VSUBS 0.014273f
C698 VTAIL.n145 VSUBS 0.031862f
C699 VTAIL.n146 VSUBS 0.031862f
C700 VTAIL.n147 VSUBS 0.014273f
C701 VTAIL.n148 VSUBS 0.01348f
C702 VTAIL.n149 VSUBS 0.025086f
C703 VTAIL.n150 VSUBS 0.025086f
C704 VTAIL.n151 VSUBS 0.01348f
C705 VTAIL.n152 VSUBS 0.014273f
C706 VTAIL.n153 VSUBS 0.031862f
C707 VTAIL.n154 VSUBS 0.077865f
C708 VTAIL.n155 VSUBS 0.014273f
C709 VTAIL.n156 VSUBS 0.01348f
C710 VTAIL.n157 VSUBS 0.056272f
C711 VTAIL.n158 VSUBS 0.039136f
C712 VTAIL.n159 VSUBS 1.16607f
C713 VTAIL.n160 VSUBS 0.027778f
C714 VTAIL.n161 VSUBS 0.025086f
C715 VTAIL.n162 VSUBS 0.01348f
C716 VTAIL.n163 VSUBS 0.031862f
C717 VTAIL.n164 VSUBS 0.014273f
C718 VTAIL.n165 VSUBS 0.025086f
C719 VTAIL.n166 VSUBS 0.01348f
C720 VTAIL.n167 VSUBS 0.031862f
C721 VTAIL.n168 VSUBS 0.014273f
C722 VTAIL.n169 VSUBS 0.025086f
C723 VTAIL.n170 VSUBS 0.01348f
C724 VTAIL.n171 VSUBS 0.023897f
C725 VTAIL.n172 VSUBS 0.020268f
C726 VTAIL.t3 VSUBS 0.068005f
C727 VTAIL.n173 VSUBS 0.12079f
C728 VTAIL.n174 VSUBS 0.734614f
C729 VTAIL.n175 VSUBS 0.01348f
C730 VTAIL.n176 VSUBS 0.014273f
C731 VTAIL.n177 VSUBS 0.031862f
C732 VTAIL.n178 VSUBS 0.031862f
C733 VTAIL.n179 VSUBS 0.014273f
C734 VTAIL.n180 VSUBS 0.01348f
C735 VTAIL.n181 VSUBS 0.025086f
C736 VTAIL.n182 VSUBS 0.025086f
C737 VTAIL.n183 VSUBS 0.01348f
C738 VTAIL.n184 VSUBS 0.014273f
C739 VTAIL.n185 VSUBS 0.031862f
C740 VTAIL.n186 VSUBS 0.031862f
C741 VTAIL.n187 VSUBS 0.014273f
C742 VTAIL.n188 VSUBS 0.01348f
C743 VTAIL.n189 VSUBS 0.025086f
C744 VTAIL.n190 VSUBS 0.025086f
C745 VTAIL.n191 VSUBS 0.01348f
C746 VTAIL.n192 VSUBS 0.014273f
C747 VTAIL.n193 VSUBS 0.031862f
C748 VTAIL.n194 VSUBS 0.077865f
C749 VTAIL.n195 VSUBS 0.014273f
C750 VTAIL.n196 VSUBS 0.01348f
C751 VTAIL.n197 VSUBS 0.056272f
C752 VTAIL.n198 VSUBS 0.039136f
C753 VTAIL.n199 VSUBS 0.203379f
C754 VTAIL.n200 VSUBS 0.027778f
C755 VTAIL.n201 VSUBS 0.025086f
C756 VTAIL.n202 VSUBS 0.01348f
C757 VTAIL.n203 VSUBS 0.031862f
C758 VTAIL.n204 VSUBS 0.014273f
C759 VTAIL.n205 VSUBS 0.025086f
C760 VTAIL.n206 VSUBS 0.01348f
C761 VTAIL.n207 VSUBS 0.031862f
C762 VTAIL.n208 VSUBS 0.014273f
C763 VTAIL.n209 VSUBS 0.025086f
C764 VTAIL.n210 VSUBS 0.01348f
C765 VTAIL.n211 VSUBS 0.023897f
C766 VTAIL.n212 VSUBS 0.020268f
C767 VTAIL.t5 VSUBS 0.068005f
C768 VTAIL.n213 VSUBS 0.12079f
C769 VTAIL.n214 VSUBS 0.734614f
C770 VTAIL.n215 VSUBS 0.01348f
C771 VTAIL.n216 VSUBS 0.014273f
C772 VTAIL.n217 VSUBS 0.031862f
C773 VTAIL.n218 VSUBS 0.031862f
C774 VTAIL.n219 VSUBS 0.014273f
C775 VTAIL.n220 VSUBS 0.01348f
C776 VTAIL.n221 VSUBS 0.025086f
C777 VTAIL.n222 VSUBS 0.025086f
C778 VTAIL.n223 VSUBS 0.01348f
C779 VTAIL.n224 VSUBS 0.014273f
C780 VTAIL.n225 VSUBS 0.031862f
C781 VTAIL.n226 VSUBS 0.031862f
C782 VTAIL.n227 VSUBS 0.014273f
C783 VTAIL.n228 VSUBS 0.01348f
C784 VTAIL.n229 VSUBS 0.025086f
C785 VTAIL.n230 VSUBS 0.025086f
C786 VTAIL.n231 VSUBS 0.01348f
C787 VTAIL.n232 VSUBS 0.014273f
C788 VTAIL.n233 VSUBS 0.031862f
C789 VTAIL.n234 VSUBS 0.077865f
C790 VTAIL.n235 VSUBS 0.014273f
C791 VTAIL.n236 VSUBS 0.01348f
C792 VTAIL.n237 VSUBS 0.056272f
C793 VTAIL.n238 VSUBS 0.039136f
C794 VTAIL.n239 VSUBS 0.203379f
C795 VTAIL.n240 VSUBS 0.027778f
C796 VTAIL.n241 VSUBS 0.025086f
C797 VTAIL.n242 VSUBS 0.01348f
C798 VTAIL.n243 VSUBS 0.031862f
C799 VTAIL.n244 VSUBS 0.014273f
C800 VTAIL.n245 VSUBS 0.025086f
C801 VTAIL.n246 VSUBS 0.01348f
C802 VTAIL.n247 VSUBS 0.031862f
C803 VTAIL.n248 VSUBS 0.014273f
C804 VTAIL.n249 VSUBS 0.025086f
C805 VTAIL.n250 VSUBS 0.01348f
C806 VTAIL.n251 VSUBS 0.023897f
C807 VTAIL.n252 VSUBS 0.020268f
C808 VTAIL.t4 VSUBS 0.068005f
C809 VTAIL.n253 VSUBS 0.12079f
C810 VTAIL.n254 VSUBS 0.734614f
C811 VTAIL.n255 VSUBS 0.01348f
C812 VTAIL.n256 VSUBS 0.014273f
C813 VTAIL.n257 VSUBS 0.031862f
C814 VTAIL.n258 VSUBS 0.031862f
C815 VTAIL.n259 VSUBS 0.014273f
C816 VTAIL.n260 VSUBS 0.01348f
C817 VTAIL.n261 VSUBS 0.025086f
C818 VTAIL.n262 VSUBS 0.025086f
C819 VTAIL.n263 VSUBS 0.01348f
C820 VTAIL.n264 VSUBS 0.014273f
C821 VTAIL.n265 VSUBS 0.031862f
C822 VTAIL.n266 VSUBS 0.031862f
C823 VTAIL.n267 VSUBS 0.014273f
C824 VTAIL.n268 VSUBS 0.01348f
C825 VTAIL.n269 VSUBS 0.025086f
C826 VTAIL.n270 VSUBS 0.025086f
C827 VTAIL.n271 VSUBS 0.01348f
C828 VTAIL.n272 VSUBS 0.014273f
C829 VTAIL.n273 VSUBS 0.031862f
C830 VTAIL.n274 VSUBS 0.077865f
C831 VTAIL.n275 VSUBS 0.014273f
C832 VTAIL.n276 VSUBS 0.01348f
C833 VTAIL.n277 VSUBS 0.056272f
C834 VTAIL.n278 VSUBS 0.039136f
C835 VTAIL.n279 VSUBS 1.16607f
C836 VTAIL.n280 VSUBS 0.027778f
C837 VTAIL.n281 VSUBS 0.025086f
C838 VTAIL.n282 VSUBS 0.01348f
C839 VTAIL.n283 VSUBS 0.031862f
C840 VTAIL.n284 VSUBS 0.014273f
C841 VTAIL.n285 VSUBS 0.025086f
C842 VTAIL.n286 VSUBS 0.01348f
C843 VTAIL.n287 VSUBS 0.031862f
C844 VTAIL.n288 VSUBS 0.014273f
C845 VTAIL.n289 VSUBS 0.025086f
C846 VTAIL.n290 VSUBS 0.01348f
C847 VTAIL.n291 VSUBS 0.023897f
C848 VTAIL.n292 VSUBS 0.020268f
C849 VTAIL.t2 VSUBS 0.068005f
C850 VTAIL.n293 VSUBS 0.12079f
C851 VTAIL.n294 VSUBS 0.734614f
C852 VTAIL.n295 VSUBS 0.01348f
C853 VTAIL.n296 VSUBS 0.014273f
C854 VTAIL.n297 VSUBS 0.031862f
C855 VTAIL.n298 VSUBS 0.031862f
C856 VTAIL.n299 VSUBS 0.014273f
C857 VTAIL.n300 VSUBS 0.01348f
C858 VTAIL.n301 VSUBS 0.025086f
C859 VTAIL.n302 VSUBS 0.025086f
C860 VTAIL.n303 VSUBS 0.01348f
C861 VTAIL.n304 VSUBS 0.014273f
C862 VTAIL.n305 VSUBS 0.031862f
C863 VTAIL.n306 VSUBS 0.031862f
C864 VTAIL.n307 VSUBS 0.014273f
C865 VTAIL.n308 VSUBS 0.01348f
C866 VTAIL.n309 VSUBS 0.025086f
C867 VTAIL.n310 VSUBS 0.025086f
C868 VTAIL.n311 VSUBS 0.01348f
C869 VTAIL.n312 VSUBS 0.014273f
C870 VTAIL.n313 VSUBS 0.031862f
C871 VTAIL.n314 VSUBS 0.077865f
C872 VTAIL.n315 VSUBS 0.014273f
C873 VTAIL.n316 VSUBS 0.01348f
C874 VTAIL.n317 VSUBS 0.056272f
C875 VTAIL.n318 VSUBS 0.039136f
C876 VTAIL.n319 VSUBS 1.0889f
C877 VP.n0 VSUBS 0.04713f
C878 VP.t2 VSUBS 1.63109f
C879 VP.n1 VSUBS 0.0381f
C880 VP.n2 VSUBS 0.04713f
C881 VP.t3 VSUBS 1.63109f
C882 VP.t1 VSUBS 1.84876f
C883 VP.t0 VSUBS 1.84614f
C884 VP.n3 VSUBS 3.0336f
C885 VP.n4 VSUBS 2.25798f
C886 VP.n5 VSUBS 0.711902f
C887 VP.n6 VSUBS 0.047942f
C888 VP.n7 VSUBS 0.093671f
C889 VP.n8 VSUBS 0.04713f
C890 VP.n9 VSUBS 0.04713f
C891 VP.n10 VSUBS 0.04713f
C892 VP.n11 VSUBS 0.093671f
C893 VP.n12 VSUBS 0.047942f
C894 VP.n13 VSUBS 0.711902f
C895 VP.n14 VSUBS 0.050361f
.ends

