* NGSPICE file created from diff_pair_sample_0762.ext - technology: sky130A

.subckt diff_pair_sample_0762 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=1.0197 ps=6.51 w=6.18 l=3
X1 VTAIL.t3 VN.t0 VDD2.t3 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=1.0197 ps=6.51 w=6.18 l=3
X2 B.t11 B.t9 B.t10 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=0 ps=0 w=6.18 l=3
X3 VDD2.t2 VN.t1 VTAIL.t1 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=1.0197 pd=6.51 as=2.4102 ps=13.14 w=6.18 l=3
X4 VTAIL.t2 VN.t2 VDD2.t1 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=1.0197 ps=6.51 w=6.18 l=3
X5 VDD1.t3 VP.t1 VTAIL.t6 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=1.0197 pd=6.51 as=2.4102 ps=13.14 w=6.18 l=3
X6 VDD1.t1 VP.t2 VTAIL.t5 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=1.0197 pd=6.51 as=2.4102 ps=13.14 w=6.18 l=3
X7 VTAIL.t4 VP.t3 VDD1.t0 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=1.0197 ps=6.51 w=6.18 l=3
X8 B.t8 B.t6 B.t7 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=0 ps=0 w=6.18 l=3
X9 B.t5 B.t3 B.t4 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=0 ps=0 w=6.18 l=3
X10 B.t2 B.t0 B.t1 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=2.4102 pd=13.14 as=0 ps=0 w=6.18 l=3
X11 VDD2.t0 VN.t3 VTAIL.t0 w_n2968_n2204# sky130_fd_pr__pfet_01v8 ad=1.0197 pd=6.51 as=2.4102 ps=13.14 w=6.18 l=3
R0 VP.n15 VP.n14 161.3
R1 VP.n13 VP.n1 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n10 VP.n2 161.3
R4 VP.n9 VP.n8 161.3
R5 VP.n7 VP.n3 161.3
R6 VP.n4 VP.t3 84.1648
R7 VP.n4 VP.t1 83.1726
R8 VP.n6 VP.n5 69.8343
R9 VP.n16 VP.n0 69.8343
R10 VP.n12 VP.n2 56.5617
R11 VP.n6 VP.t0 49.6465
R12 VP.n0 VP.t2 49.6465
R13 VP.n5 VP.n4 46.1699
R14 VP.n8 VP.n7 24.5923
R15 VP.n8 VP.n2 24.5923
R16 VP.n13 VP.n12 24.5923
R17 VP.n14 VP.n13 24.5923
R18 VP.n7 VP.n6 20.4117
R19 VP.n14 VP.n0 20.4117
R20 VP.n5 VP.n3 0.354861
R21 VP.n16 VP.n15 0.354861
R22 VP VP.n16 0.267071
R23 VP.n9 VP.n3 0.189894
R24 VP.n10 VP.n9 0.189894
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n1 0.189894
R27 VP.n15 VP.n1 0.189894
R28 VDD1 VDD1.n1 131.294
R29 VDD1 VDD1.n0 93.1729
R30 VDD1.n0 VDD1.t0 5.26021
R31 VDD1.n0 VDD1.t3 5.26021
R32 VDD1.n1 VDD1.t2 5.26021
R33 VDD1.n1 VDD1.t1 5.26021
R34 VTAIL.n5 VTAIL.t4 81.6967
R35 VTAIL.n4 VTAIL.t1 81.6967
R36 VTAIL.n3 VTAIL.t2 81.6967
R37 VTAIL.n7 VTAIL.t0 81.6957
R38 VTAIL.n0 VTAIL.t3 81.6957
R39 VTAIL.n1 VTAIL.t5 81.6957
R40 VTAIL.n2 VTAIL.t7 81.6957
R41 VTAIL.n6 VTAIL.t6 81.6956
R42 VTAIL.n7 VTAIL.n6 20.5652
R43 VTAIL.n3 VTAIL.n2 20.5652
R44 VTAIL.n4 VTAIL.n3 2.87119
R45 VTAIL.n6 VTAIL.n5 2.87119
R46 VTAIL.n2 VTAIL.n1 2.87119
R47 VTAIL VTAIL.n0 1.49403
R48 VTAIL VTAIL.n7 1.37766
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 VN.n1 VN.t1 84.1651
R52 VN.n0 VN.t0 84.1651
R53 VN.n0 VN.t3 83.1725
R54 VN.n1 VN.t2 83.1725
R55 VN VN.n1 46.3352
R56 VN VN.n0 2.99808
R57 VDD2.n2 VDD2.n0 130.77
R58 VDD2.n2 VDD2.n1 93.1147
R59 VDD2.n1 VDD2.t1 5.26021
R60 VDD2.n1 VDD2.t2 5.26021
R61 VDD2.n0 VDD2.t3 5.26021
R62 VDD2.n0 VDD2.t0 5.26021
R63 VDD2 VDD2.n2 0.0586897
R64 B.n287 B.n92 585
R65 B.n286 B.n285 585
R66 B.n284 B.n93 585
R67 B.n283 B.n282 585
R68 B.n281 B.n94 585
R69 B.n280 B.n279 585
R70 B.n278 B.n95 585
R71 B.n277 B.n276 585
R72 B.n275 B.n96 585
R73 B.n274 B.n273 585
R74 B.n272 B.n97 585
R75 B.n271 B.n270 585
R76 B.n269 B.n98 585
R77 B.n268 B.n267 585
R78 B.n266 B.n99 585
R79 B.n265 B.n264 585
R80 B.n263 B.n100 585
R81 B.n262 B.n261 585
R82 B.n260 B.n101 585
R83 B.n259 B.n258 585
R84 B.n257 B.n102 585
R85 B.n256 B.n255 585
R86 B.n254 B.n103 585
R87 B.n253 B.n252 585
R88 B.n251 B.n104 585
R89 B.n250 B.n249 585
R90 B.n245 B.n105 585
R91 B.n244 B.n243 585
R92 B.n242 B.n106 585
R93 B.n241 B.n240 585
R94 B.n239 B.n107 585
R95 B.n238 B.n237 585
R96 B.n236 B.n108 585
R97 B.n235 B.n234 585
R98 B.n232 B.n109 585
R99 B.n231 B.n230 585
R100 B.n229 B.n112 585
R101 B.n228 B.n227 585
R102 B.n226 B.n113 585
R103 B.n225 B.n224 585
R104 B.n223 B.n114 585
R105 B.n222 B.n221 585
R106 B.n220 B.n115 585
R107 B.n219 B.n218 585
R108 B.n217 B.n116 585
R109 B.n216 B.n215 585
R110 B.n214 B.n117 585
R111 B.n213 B.n212 585
R112 B.n211 B.n118 585
R113 B.n210 B.n209 585
R114 B.n208 B.n119 585
R115 B.n207 B.n206 585
R116 B.n205 B.n120 585
R117 B.n204 B.n203 585
R118 B.n202 B.n121 585
R119 B.n201 B.n200 585
R120 B.n199 B.n122 585
R121 B.n198 B.n197 585
R122 B.n196 B.n123 585
R123 B.n289 B.n288 585
R124 B.n290 B.n91 585
R125 B.n292 B.n291 585
R126 B.n293 B.n90 585
R127 B.n295 B.n294 585
R128 B.n296 B.n89 585
R129 B.n298 B.n297 585
R130 B.n299 B.n88 585
R131 B.n301 B.n300 585
R132 B.n302 B.n87 585
R133 B.n304 B.n303 585
R134 B.n305 B.n86 585
R135 B.n307 B.n306 585
R136 B.n308 B.n85 585
R137 B.n310 B.n309 585
R138 B.n311 B.n84 585
R139 B.n313 B.n312 585
R140 B.n314 B.n83 585
R141 B.n316 B.n315 585
R142 B.n317 B.n82 585
R143 B.n319 B.n318 585
R144 B.n320 B.n81 585
R145 B.n322 B.n321 585
R146 B.n323 B.n80 585
R147 B.n325 B.n324 585
R148 B.n326 B.n79 585
R149 B.n328 B.n327 585
R150 B.n329 B.n78 585
R151 B.n331 B.n330 585
R152 B.n332 B.n77 585
R153 B.n334 B.n333 585
R154 B.n335 B.n76 585
R155 B.n337 B.n336 585
R156 B.n338 B.n75 585
R157 B.n340 B.n339 585
R158 B.n341 B.n74 585
R159 B.n343 B.n342 585
R160 B.n344 B.n73 585
R161 B.n346 B.n345 585
R162 B.n347 B.n72 585
R163 B.n349 B.n348 585
R164 B.n350 B.n71 585
R165 B.n352 B.n351 585
R166 B.n353 B.n70 585
R167 B.n355 B.n354 585
R168 B.n356 B.n69 585
R169 B.n358 B.n357 585
R170 B.n359 B.n68 585
R171 B.n361 B.n360 585
R172 B.n362 B.n67 585
R173 B.n364 B.n363 585
R174 B.n365 B.n66 585
R175 B.n367 B.n366 585
R176 B.n368 B.n65 585
R177 B.n370 B.n369 585
R178 B.n371 B.n64 585
R179 B.n373 B.n372 585
R180 B.n374 B.n63 585
R181 B.n376 B.n375 585
R182 B.n377 B.n62 585
R183 B.n379 B.n378 585
R184 B.n380 B.n61 585
R185 B.n382 B.n381 585
R186 B.n383 B.n60 585
R187 B.n385 B.n384 585
R188 B.n386 B.n59 585
R189 B.n388 B.n387 585
R190 B.n389 B.n58 585
R191 B.n391 B.n390 585
R192 B.n392 B.n57 585
R193 B.n394 B.n393 585
R194 B.n395 B.n56 585
R195 B.n397 B.n396 585
R196 B.n398 B.n55 585
R197 B.n400 B.n399 585
R198 B.n401 B.n54 585
R199 B.n492 B.n491 585
R200 B.n490 B.n21 585
R201 B.n489 B.n488 585
R202 B.n487 B.n22 585
R203 B.n486 B.n485 585
R204 B.n484 B.n23 585
R205 B.n483 B.n482 585
R206 B.n481 B.n24 585
R207 B.n480 B.n479 585
R208 B.n478 B.n25 585
R209 B.n477 B.n476 585
R210 B.n475 B.n26 585
R211 B.n474 B.n473 585
R212 B.n472 B.n27 585
R213 B.n471 B.n470 585
R214 B.n469 B.n28 585
R215 B.n468 B.n467 585
R216 B.n466 B.n29 585
R217 B.n465 B.n464 585
R218 B.n463 B.n30 585
R219 B.n462 B.n461 585
R220 B.n460 B.n31 585
R221 B.n459 B.n458 585
R222 B.n457 B.n32 585
R223 B.n456 B.n455 585
R224 B.n453 B.n33 585
R225 B.n452 B.n451 585
R226 B.n450 B.n36 585
R227 B.n449 B.n448 585
R228 B.n447 B.n37 585
R229 B.n446 B.n445 585
R230 B.n444 B.n38 585
R231 B.n443 B.n442 585
R232 B.n441 B.n39 585
R233 B.n439 B.n438 585
R234 B.n437 B.n42 585
R235 B.n436 B.n435 585
R236 B.n434 B.n43 585
R237 B.n433 B.n432 585
R238 B.n431 B.n44 585
R239 B.n430 B.n429 585
R240 B.n428 B.n45 585
R241 B.n427 B.n426 585
R242 B.n425 B.n46 585
R243 B.n424 B.n423 585
R244 B.n422 B.n47 585
R245 B.n421 B.n420 585
R246 B.n419 B.n48 585
R247 B.n418 B.n417 585
R248 B.n416 B.n49 585
R249 B.n415 B.n414 585
R250 B.n413 B.n50 585
R251 B.n412 B.n411 585
R252 B.n410 B.n51 585
R253 B.n409 B.n408 585
R254 B.n407 B.n52 585
R255 B.n406 B.n405 585
R256 B.n404 B.n53 585
R257 B.n403 B.n402 585
R258 B.n493 B.n20 585
R259 B.n495 B.n494 585
R260 B.n496 B.n19 585
R261 B.n498 B.n497 585
R262 B.n499 B.n18 585
R263 B.n501 B.n500 585
R264 B.n502 B.n17 585
R265 B.n504 B.n503 585
R266 B.n505 B.n16 585
R267 B.n507 B.n506 585
R268 B.n508 B.n15 585
R269 B.n510 B.n509 585
R270 B.n511 B.n14 585
R271 B.n513 B.n512 585
R272 B.n514 B.n13 585
R273 B.n516 B.n515 585
R274 B.n517 B.n12 585
R275 B.n519 B.n518 585
R276 B.n520 B.n11 585
R277 B.n522 B.n521 585
R278 B.n523 B.n10 585
R279 B.n525 B.n524 585
R280 B.n526 B.n9 585
R281 B.n528 B.n527 585
R282 B.n529 B.n8 585
R283 B.n531 B.n530 585
R284 B.n532 B.n7 585
R285 B.n534 B.n533 585
R286 B.n535 B.n6 585
R287 B.n537 B.n536 585
R288 B.n538 B.n5 585
R289 B.n540 B.n539 585
R290 B.n541 B.n4 585
R291 B.n543 B.n542 585
R292 B.n544 B.n3 585
R293 B.n546 B.n545 585
R294 B.n547 B.n0 585
R295 B.n2 B.n1 585
R296 B.n142 B.n141 585
R297 B.n144 B.n143 585
R298 B.n145 B.n140 585
R299 B.n147 B.n146 585
R300 B.n148 B.n139 585
R301 B.n150 B.n149 585
R302 B.n151 B.n138 585
R303 B.n153 B.n152 585
R304 B.n154 B.n137 585
R305 B.n156 B.n155 585
R306 B.n157 B.n136 585
R307 B.n159 B.n158 585
R308 B.n160 B.n135 585
R309 B.n162 B.n161 585
R310 B.n163 B.n134 585
R311 B.n165 B.n164 585
R312 B.n166 B.n133 585
R313 B.n168 B.n167 585
R314 B.n169 B.n132 585
R315 B.n171 B.n170 585
R316 B.n172 B.n131 585
R317 B.n174 B.n173 585
R318 B.n175 B.n130 585
R319 B.n177 B.n176 585
R320 B.n178 B.n129 585
R321 B.n180 B.n179 585
R322 B.n181 B.n128 585
R323 B.n183 B.n182 585
R324 B.n184 B.n127 585
R325 B.n186 B.n185 585
R326 B.n187 B.n126 585
R327 B.n189 B.n188 585
R328 B.n190 B.n125 585
R329 B.n192 B.n191 585
R330 B.n193 B.n124 585
R331 B.n195 B.n194 585
R332 B.n194 B.n123 463.671
R333 B.n288 B.n287 463.671
R334 B.n402 B.n401 463.671
R335 B.n493 B.n492 463.671
R336 B.n110 B.t9 258.226
R337 B.n246 B.t6 258.226
R338 B.n40 B.t3 258.226
R339 B.n34 B.t0 258.226
R340 B.n549 B.n548 256.663
R341 B.n548 B.n547 235.042
R342 B.n548 B.n2 235.042
R343 B.n246 B.t7 176.466
R344 B.n40 B.t5 176.466
R345 B.n110 B.t10 176.46
R346 B.n34 B.t2 176.46
R347 B.n198 B.n123 163.367
R348 B.n199 B.n198 163.367
R349 B.n200 B.n199 163.367
R350 B.n200 B.n121 163.367
R351 B.n204 B.n121 163.367
R352 B.n205 B.n204 163.367
R353 B.n206 B.n205 163.367
R354 B.n206 B.n119 163.367
R355 B.n210 B.n119 163.367
R356 B.n211 B.n210 163.367
R357 B.n212 B.n211 163.367
R358 B.n212 B.n117 163.367
R359 B.n216 B.n117 163.367
R360 B.n217 B.n216 163.367
R361 B.n218 B.n217 163.367
R362 B.n218 B.n115 163.367
R363 B.n222 B.n115 163.367
R364 B.n223 B.n222 163.367
R365 B.n224 B.n223 163.367
R366 B.n224 B.n113 163.367
R367 B.n228 B.n113 163.367
R368 B.n229 B.n228 163.367
R369 B.n230 B.n229 163.367
R370 B.n230 B.n109 163.367
R371 B.n235 B.n109 163.367
R372 B.n236 B.n235 163.367
R373 B.n237 B.n236 163.367
R374 B.n237 B.n107 163.367
R375 B.n241 B.n107 163.367
R376 B.n242 B.n241 163.367
R377 B.n243 B.n242 163.367
R378 B.n243 B.n105 163.367
R379 B.n250 B.n105 163.367
R380 B.n251 B.n250 163.367
R381 B.n252 B.n251 163.367
R382 B.n252 B.n103 163.367
R383 B.n256 B.n103 163.367
R384 B.n257 B.n256 163.367
R385 B.n258 B.n257 163.367
R386 B.n258 B.n101 163.367
R387 B.n262 B.n101 163.367
R388 B.n263 B.n262 163.367
R389 B.n264 B.n263 163.367
R390 B.n264 B.n99 163.367
R391 B.n268 B.n99 163.367
R392 B.n269 B.n268 163.367
R393 B.n270 B.n269 163.367
R394 B.n270 B.n97 163.367
R395 B.n274 B.n97 163.367
R396 B.n275 B.n274 163.367
R397 B.n276 B.n275 163.367
R398 B.n276 B.n95 163.367
R399 B.n280 B.n95 163.367
R400 B.n281 B.n280 163.367
R401 B.n282 B.n281 163.367
R402 B.n282 B.n93 163.367
R403 B.n286 B.n93 163.367
R404 B.n287 B.n286 163.367
R405 B.n401 B.n400 163.367
R406 B.n400 B.n55 163.367
R407 B.n396 B.n55 163.367
R408 B.n396 B.n395 163.367
R409 B.n395 B.n394 163.367
R410 B.n394 B.n57 163.367
R411 B.n390 B.n57 163.367
R412 B.n390 B.n389 163.367
R413 B.n389 B.n388 163.367
R414 B.n388 B.n59 163.367
R415 B.n384 B.n59 163.367
R416 B.n384 B.n383 163.367
R417 B.n383 B.n382 163.367
R418 B.n382 B.n61 163.367
R419 B.n378 B.n61 163.367
R420 B.n378 B.n377 163.367
R421 B.n377 B.n376 163.367
R422 B.n376 B.n63 163.367
R423 B.n372 B.n63 163.367
R424 B.n372 B.n371 163.367
R425 B.n371 B.n370 163.367
R426 B.n370 B.n65 163.367
R427 B.n366 B.n65 163.367
R428 B.n366 B.n365 163.367
R429 B.n365 B.n364 163.367
R430 B.n364 B.n67 163.367
R431 B.n360 B.n67 163.367
R432 B.n360 B.n359 163.367
R433 B.n359 B.n358 163.367
R434 B.n358 B.n69 163.367
R435 B.n354 B.n69 163.367
R436 B.n354 B.n353 163.367
R437 B.n353 B.n352 163.367
R438 B.n352 B.n71 163.367
R439 B.n348 B.n71 163.367
R440 B.n348 B.n347 163.367
R441 B.n347 B.n346 163.367
R442 B.n346 B.n73 163.367
R443 B.n342 B.n73 163.367
R444 B.n342 B.n341 163.367
R445 B.n341 B.n340 163.367
R446 B.n340 B.n75 163.367
R447 B.n336 B.n75 163.367
R448 B.n336 B.n335 163.367
R449 B.n335 B.n334 163.367
R450 B.n334 B.n77 163.367
R451 B.n330 B.n77 163.367
R452 B.n330 B.n329 163.367
R453 B.n329 B.n328 163.367
R454 B.n328 B.n79 163.367
R455 B.n324 B.n79 163.367
R456 B.n324 B.n323 163.367
R457 B.n323 B.n322 163.367
R458 B.n322 B.n81 163.367
R459 B.n318 B.n81 163.367
R460 B.n318 B.n317 163.367
R461 B.n317 B.n316 163.367
R462 B.n316 B.n83 163.367
R463 B.n312 B.n83 163.367
R464 B.n312 B.n311 163.367
R465 B.n311 B.n310 163.367
R466 B.n310 B.n85 163.367
R467 B.n306 B.n85 163.367
R468 B.n306 B.n305 163.367
R469 B.n305 B.n304 163.367
R470 B.n304 B.n87 163.367
R471 B.n300 B.n87 163.367
R472 B.n300 B.n299 163.367
R473 B.n299 B.n298 163.367
R474 B.n298 B.n89 163.367
R475 B.n294 B.n89 163.367
R476 B.n294 B.n293 163.367
R477 B.n293 B.n292 163.367
R478 B.n292 B.n91 163.367
R479 B.n288 B.n91 163.367
R480 B.n492 B.n21 163.367
R481 B.n488 B.n21 163.367
R482 B.n488 B.n487 163.367
R483 B.n487 B.n486 163.367
R484 B.n486 B.n23 163.367
R485 B.n482 B.n23 163.367
R486 B.n482 B.n481 163.367
R487 B.n481 B.n480 163.367
R488 B.n480 B.n25 163.367
R489 B.n476 B.n25 163.367
R490 B.n476 B.n475 163.367
R491 B.n475 B.n474 163.367
R492 B.n474 B.n27 163.367
R493 B.n470 B.n27 163.367
R494 B.n470 B.n469 163.367
R495 B.n469 B.n468 163.367
R496 B.n468 B.n29 163.367
R497 B.n464 B.n29 163.367
R498 B.n464 B.n463 163.367
R499 B.n463 B.n462 163.367
R500 B.n462 B.n31 163.367
R501 B.n458 B.n31 163.367
R502 B.n458 B.n457 163.367
R503 B.n457 B.n456 163.367
R504 B.n456 B.n33 163.367
R505 B.n451 B.n33 163.367
R506 B.n451 B.n450 163.367
R507 B.n450 B.n449 163.367
R508 B.n449 B.n37 163.367
R509 B.n445 B.n37 163.367
R510 B.n445 B.n444 163.367
R511 B.n444 B.n443 163.367
R512 B.n443 B.n39 163.367
R513 B.n438 B.n39 163.367
R514 B.n438 B.n437 163.367
R515 B.n437 B.n436 163.367
R516 B.n436 B.n43 163.367
R517 B.n432 B.n43 163.367
R518 B.n432 B.n431 163.367
R519 B.n431 B.n430 163.367
R520 B.n430 B.n45 163.367
R521 B.n426 B.n45 163.367
R522 B.n426 B.n425 163.367
R523 B.n425 B.n424 163.367
R524 B.n424 B.n47 163.367
R525 B.n420 B.n47 163.367
R526 B.n420 B.n419 163.367
R527 B.n419 B.n418 163.367
R528 B.n418 B.n49 163.367
R529 B.n414 B.n49 163.367
R530 B.n414 B.n413 163.367
R531 B.n413 B.n412 163.367
R532 B.n412 B.n51 163.367
R533 B.n408 B.n51 163.367
R534 B.n408 B.n407 163.367
R535 B.n407 B.n406 163.367
R536 B.n406 B.n53 163.367
R537 B.n402 B.n53 163.367
R538 B.n494 B.n493 163.367
R539 B.n494 B.n19 163.367
R540 B.n498 B.n19 163.367
R541 B.n499 B.n498 163.367
R542 B.n500 B.n499 163.367
R543 B.n500 B.n17 163.367
R544 B.n504 B.n17 163.367
R545 B.n505 B.n504 163.367
R546 B.n506 B.n505 163.367
R547 B.n506 B.n15 163.367
R548 B.n510 B.n15 163.367
R549 B.n511 B.n510 163.367
R550 B.n512 B.n511 163.367
R551 B.n512 B.n13 163.367
R552 B.n516 B.n13 163.367
R553 B.n517 B.n516 163.367
R554 B.n518 B.n517 163.367
R555 B.n518 B.n11 163.367
R556 B.n522 B.n11 163.367
R557 B.n523 B.n522 163.367
R558 B.n524 B.n523 163.367
R559 B.n524 B.n9 163.367
R560 B.n528 B.n9 163.367
R561 B.n529 B.n528 163.367
R562 B.n530 B.n529 163.367
R563 B.n530 B.n7 163.367
R564 B.n534 B.n7 163.367
R565 B.n535 B.n534 163.367
R566 B.n536 B.n535 163.367
R567 B.n536 B.n5 163.367
R568 B.n540 B.n5 163.367
R569 B.n541 B.n540 163.367
R570 B.n542 B.n541 163.367
R571 B.n542 B.n3 163.367
R572 B.n546 B.n3 163.367
R573 B.n547 B.n546 163.367
R574 B.n141 B.n2 163.367
R575 B.n144 B.n141 163.367
R576 B.n145 B.n144 163.367
R577 B.n146 B.n145 163.367
R578 B.n146 B.n139 163.367
R579 B.n150 B.n139 163.367
R580 B.n151 B.n150 163.367
R581 B.n152 B.n151 163.367
R582 B.n152 B.n137 163.367
R583 B.n156 B.n137 163.367
R584 B.n157 B.n156 163.367
R585 B.n158 B.n157 163.367
R586 B.n158 B.n135 163.367
R587 B.n162 B.n135 163.367
R588 B.n163 B.n162 163.367
R589 B.n164 B.n163 163.367
R590 B.n164 B.n133 163.367
R591 B.n168 B.n133 163.367
R592 B.n169 B.n168 163.367
R593 B.n170 B.n169 163.367
R594 B.n170 B.n131 163.367
R595 B.n174 B.n131 163.367
R596 B.n175 B.n174 163.367
R597 B.n176 B.n175 163.367
R598 B.n176 B.n129 163.367
R599 B.n180 B.n129 163.367
R600 B.n181 B.n180 163.367
R601 B.n182 B.n181 163.367
R602 B.n182 B.n127 163.367
R603 B.n186 B.n127 163.367
R604 B.n187 B.n186 163.367
R605 B.n188 B.n187 163.367
R606 B.n188 B.n125 163.367
R607 B.n192 B.n125 163.367
R608 B.n193 B.n192 163.367
R609 B.n194 B.n193 163.367
R610 B.n247 B.t8 111.885
R611 B.n41 B.t4 111.885
R612 B.n111 B.t11 111.879
R613 B.n35 B.t1 111.879
R614 B.n111 B.n110 64.5823
R615 B.n247 B.n246 64.5823
R616 B.n41 B.n40 64.5823
R617 B.n35 B.n34 64.5823
R618 B.n233 B.n111 59.5399
R619 B.n248 B.n247 59.5399
R620 B.n440 B.n41 59.5399
R621 B.n454 B.n35 59.5399
R622 B.n289 B.n92 30.1273
R623 B.n491 B.n20 30.1273
R624 B.n403 B.n54 30.1273
R625 B.n196 B.n195 30.1273
R626 B B.n549 18.0485
R627 B.n495 B.n20 10.6151
R628 B.n496 B.n495 10.6151
R629 B.n497 B.n496 10.6151
R630 B.n497 B.n18 10.6151
R631 B.n501 B.n18 10.6151
R632 B.n502 B.n501 10.6151
R633 B.n503 B.n502 10.6151
R634 B.n503 B.n16 10.6151
R635 B.n507 B.n16 10.6151
R636 B.n508 B.n507 10.6151
R637 B.n509 B.n508 10.6151
R638 B.n509 B.n14 10.6151
R639 B.n513 B.n14 10.6151
R640 B.n514 B.n513 10.6151
R641 B.n515 B.n514 10.6151
R642 B.n515 B.n12 10.6151
R643 B.n519 B.n12 10.6151
R644 B.n520 B.n519 10.6151
R645 B.n521 B.n520 10.6151
R646 B.n521 B.n10 10.6151
R647 B.n525 B.n10 10.6151
R648 B.n526 B.n525 10.6151
R649 B.n527 B.n526 10.6151
R650 B.n527 B.n8 10.6151
R651 B.n531 B.n8 10.6151
R652 B.n532 B.n531 10.6151
R653 B.n533 B.n532 10.6151
R654 B.n533 B.n6 10.6151
R655 B.n537 B.n6 10.6151
R656 B.n538 B.n537 10.6151
R657 B.n539 B.n538 10.6151
R658 B.n539 B.n4 10.6151
R659 B.n543 B.n4 10.6151
R660 B.n544 B.n543 10.6151
R661 B.n545 B.n544 10.6151
R662 B.n545 B.n0 10.6151
R663 B.n491 B.n490 10.6151
R664 B.n490 B.n489 10.6151
R665 B.n489 B.n22 10.6151
R666 B.n485 B.n22 10.6151
R667 B.n485 B.n484 10.6151
R668 B.n484 B.n483 10.6151
R669 B.n483 B.n24 10.6151
R670 B.n479 B.n24 10.6151
R671 B.n479 B.n478 10.6151
R672 B.n478 B.n477 10.6151
R673 B.n477 B.n26 10.6151
R674 B.n473 B.n26 10.6151
R675 B.n473 B.n472 10.6151
R676 B.n472 B.n471 10.6151
R677 B.n471 B.n28 10.6151
R678 B.n467 B.n28 10.6151
R679 B.n467 B.n466 10.6151
R680 B.n466 B.n465 10.6151
R681 B.n465 B.n30 10.6151
R682 B.n461 B.n30 10.6151
R683 B.n461 B.n460 10.6151
R684 B.n460 B.n459 10.6151
R685 B.n459 B.n32 10.6151
R686 B.n455 B.n32 10.6151
R687 B.n453 B.n452 10.6151
R688 B.n452 B.n36 10.6151
R689 B.n448 B.n36 10.6151
R690 B.n448 B.n447 10.6151
R691 B.n447 B.n446 10.6151
R692 B.n446 B.n38 10.6151
R693 B.n442 B.n38 10.6151
R694 B.n442 B.n441 10.6151
R695 B.n439 B.n42 10.6151
R696 B.n435 B.n42 10.6151
R697 B.n435 B.n434 10.6151
R698 B.n434 B.n433 10.6151
R699 B.n433 B.n44 10.6151
R700 B.n429 B.n44 10.6151
R701 B.n429 B.n428 10.6151
R702 B.n428 B.n427 10.6151
R703 B.n427 B.n46 10.6151
R704 B.n423 B.n46 10.6151
R705 B.n423 B.n422 10.6151
R706 B.n422 B.n421 10.6151
R707 B.n421 B.n48 10.6151
R708 B.n417 B.n48 10.6151
R709 B.n417 B.n416 10.6151
R710 B.n416 B.n415 10.6151
R711 B.n415 B.n50 10.6151
R712 B.n411 B.n50 10.6151
R713 B.n411 B.n410 10.6151
R714 B.n410 B.n409 10.6151
R715 B.n409 B.n52 10.6151
R716 B.n405 B.n52 10.6151
R717 B.n405 B.n404 10.6151
R718 B.n404 B.n403 10.6151
R719 B.n399 B.n54 10.6151
R720 B.n399 B.n398 10.6151
R721 B.n398 B.n397 10.6151
R722 B.n397 B.n56 10.6151
R723 B.n393 B.n56 10.6151
R724 B.n393 B.n392 10.6151
R725 B.n392 B.n391 10.6151
R726 B.n391 B.n58 10.6151
R727 B.n387 B.n58 10.6151
R728 B.n387 B.n386 10.6151
R729 B.n386 B.n385 10.6151
R730 B.n385 B.n60 10.6151
R731 B.n381 B.n60 10.6151
R732 B.n381 B.n380 10.6151
R733 B.n380 B.n379 10.6151
R734 B.n379 B.n62 10.6151
R735 B.n375 B.n62 10.6151
R736 B.n375 B.n374 10.6151
R737 B.n374 B.n373 10.6151
R738 B.n373 B.n64 10.6151
R739 B.n369 B.n64 10.6151
R740 B.n369 B.n368 10.6151
R741 B.n368 B.n367 10.6151
R742 B.n367 B.n66 10.6151
R743 B.n363 B.n66 10.6151
R744 B.n363 B.n362 10.6151
R745 B.n362 B.n361 10.6151
R746 B.n361 B.n68 10.6151
R747 B.n357 B.n68 10.6151
R748 B.n357 B.n356 10.6151
R749 B.n356 B.n355 10.6151
R750 B.n355 B.n70 10.6151
R751 B.n351 B.n70 10.6151
R752 B.n351 B.n350 10.6151
R753 B.n350 B.n349 10.6151
R754 B.n349 B.n72 10.6151
R755 B.n345 B.n72 10.6151
R756 B.n345 B.n344 10.6151
R757 B.n344 B.n343 10.6151
R758 B.n343 B.n74 10.6151
R759 B.n339 B.n74 10.6151
R760 B.n339 B.n338 10.6151
R761 B.n338 B.n337 10.6151
R762 B.n337 B.n76 10.6151
R763 B.n333 B.n76 10.6151
R764 B.n333 B.n332 10.6151
R765 B.n332 B.n331 10.6151
R766 B.n331 B.n78 10.6151
R767 B.n327 B.n78 10.6151
R768 B.n327 B.n326 10.6151
R769 B.n326 B.n325 10.6151
R770 B.n325 B.n80 10.6151
R771 B.n321 B.n80 10.6151
R772 B.n321 B.n320 10.6151
R773 B.n320 B.n319 10.6151
R774 B.n319 B.n82 10.6151
R775 B.n315 B.n82 10.6151
R776 B.n315 B.n314 10.6151
R777 B.n314 B.n313 10.6151
R778 B.n313 B.n84 10.6151
R779 B.n309 B.n84 10.6151
R780 B.n309 B.n308 10.6151
R781 B.n308 B.n307 10.6151
R782 B.n307 B.n86 10.6151
R783 B.n303 B.n86 10.6151
R784 B.n303 B.n302 10.6151
R785 B.n302 B.n301 10.6151
R786 B.n301 B.n88 10.6151
R787 B.n297 B.n88 10.6151
R788 B.n297 B.n296 10.6151
R789 B.n296 B.n295 10.6151
R790 B.n295 B.n90 10.6151
R791 B.n291 B.n90 10.6151
R792 B.n291 B.n290 10.6151
R793 B.n290 B.n289 10.6151
R794 B.n142 B.n1 10.6151
R795 B.n143 B.n142 10.6151
R796 B.n143 B.n140 10.6151
R797 B.n147 B.n140 10.6151
R798 B.n148 B.n147 10.6151
R799 B.n149 B.n148 10.6151
R800 B.n149 B.n138 10.6151
R801 B.n153 B.n138 10.6151
R802 B.n154 B.n153 10.6151
R803 B.n155 B.n154 10.6151
R804 B.n155 B.n136 10.6151
R805 B.n159 B.n136 10.6151
R806 B.n160 B.n159 10.6151
R807 B.n161 B.n160 10.6151
R808 B.n161 B.n134 10.6151
R809 B.n165 B.n134 10.6151
R810 B.n166 B.n165 10.6151
R811 B.n167 B.n166 10.6151
R812 B.n167 B.n132 10.6151
R813 B.n171 B.n132 10.6151
R814 B.n172 B.n171 10.6151
R815 B.n173 B.n172 10.6151
R816 B.n173 B.n130 10.6151
R817 B.n177 B.n130 10.6151
R818 B.n178 B.n177 10.6151
R819 B.n179 B.n178 10.6151
R820 B.n179 B.n128 10.6151
R821 B.n183 B.n128 10.6151
R822 B.n184 B.n183 10.6151
R823 B.n185 B.n184 10.6151
R824 B.n185 B.n126 10.6151
R825 B.n189 B.n126 10.6151
R826 B.n190 B.n189 10.6151
R827 B.n191 B.n190 10.6151
R828 B.n191 B.n124 10.6151
R829 B.n195 B.n124 10.6151
R830 B.n197 B.n196 10.6151
R831 B.n197 B.n122 10.6151
R832 B.n201 B.n122 10.6151
R833 B.n202 B.n201 10.6151
R834 B.n203 B.n202 10.6151
R835 B.n203 B.n120 10.6151
R836 B.n207 B.n120 10.6151
R837 B.n208 B.n207 10.6151
R838 B.n209 B.n208 10.6151
R839 B.n209 B.n118 10.6151
R840 B.n213 B.n118 10.6151
R841 B.n214 B.n213 10.6151
R842 B.n215 B.n214 10.6151
R843 B.n215 B.n116 10.6151
R844 B.n219 B.n116 10.6151
R845 B.n220 B.n219 10.6151
R846 B.n221 B.n220 10.6151
R847 B.n221 B.n114 10.6151
R848 B.n225 B.n114 10.6151
R849 B.n226 B.n225 10.6151
R850 B.n227 B.n226 10.6151
R851 B.n227 B.n112 10.6151
R852 B.n231 B.n112 10.6151
R853 B.n232 B.n231 10.6151
R854 B.n234 B.n108 10.6151
R855 B.n238 B.n108 10.6151
R856 B.n239 B.n238 10.6151
R857 B.n240 B.n239 10.6151
R858 B.n240 B.n106 10.6151
R859 B.n244 B.n106 10.6151
R860 B.n245 B.n244 10.6151
R861 B.n249 B.n245 10.6151
R862 B.n253 B.n104 10.6151
R863 B.n254 B.n253 10.6151
R864 B.n255 B.n254 10.6151
R865 B.n255 B.n102 10.6151
R866 B.n259 B.n102 10.6151
R867 B.n260 B.n259 10.6151
R868 B.n261 B.n260 10.6151
R869 B.n261 B.n100 10.6151
R870 B.n265 B.n100 10.6151
R871 B.n266 B.n265 10.6151
R872 B.n267 B.n266 10.6151
R873 B.n267 B.n98 10.6151
R874 B.n271 B.n98 10.6151
R875 B.n272 B.n271 10.6151
R876 B.n273 B.n272 10.6151
R877 B.n273 B.n96 10.6151
R878 B.n277 B.n96 10.6151
R879 B.n278 B.n277 10.6151
R880 B.n279 B.n278 10.6151
R881 B.n279 B.n94 10.6151
R882 B.n283 B.n94 10.6151
R883 B.n284 B.n283 10.6151
R884 B.n285 B.n284 10.6151
R885 B.n285 B.n92 10.6151
R886 B.n549 B.n0 8.11757
R887 B.n549 B.n1 8.11757
R888 B.n454 B.n453 6.5566
R889 B.n441 B.n440 6.5566
R890 B.n234 B.n233 6.5566
R891 B.n249 B.n248 6.5566
R892 B.n455 B.n454 4.05904
R893 B.n440 B.n439 4.05904
R894 B.n233 B.n232 4.05904
R895 B.n248 B.n104 4.05904
C0 w_n2968_n2204# B 8.11621f
C1 VTAIL B 3.15797f
C2 VDD1 B 1.17539f
C3 VDD2 B 1.23418f
C4 VP B 1.75287f
C5 VTAIL w_n2968_n2204# 2.68982f
C6 VDD1 w_n2968_n2204# 1.37509f
C7 VN B 1.11617f
C8 VDD2 w_n2968_n2204# 1.44007f
C9 VP w_n2968_n2204# 5.37265f
C10 VN w_n2968_n2204# 4.99009f
C11 VDD1 VTAIL 4.17802f
C12 VDD2 VTAIL 4.23491f
C13 VDD2 VDD1 1.12335f
C14 VP VTAIL 3.0411f
C15 VDD1 VP 2.93122f
C16 VN VTAIL 3.02699f
C17 VDD1 VN 0.149837f
C18 VDD2 VP 0.420233f
C19 VDD2 VN 2.66167f
C20 VP VN 5.39893f
C21 VDD2 VSUBS 0.873567f
C22 VDD1 VSUBS 5.21576f
C23 VTAIL VSUBS 0.737297f
C24 VN VSUBS 5.53897f
C25 VP VSUBS 2.164113f
C26 B VSUBS 4.130165f
C27 w_n2968_n2204# VSUBS 81.5963f
C28 B.n0 VSUBS 0.007101f
C29 B.n1 VSUBS 0.007101f
C30 B.n2 VSUBS 0.010502f
C31 B.n3 VSUBS 0.008047f
C32 B.n4 VSUBS 0.008047f
C33 B.n5 VSUBS 0.008047f
C34 B.n6 VSUBS 0.008047f
C35 B.n7 VSUBS 0.008047f
C36 B.n8 VSUBS 0.008047f
C37 B.n9 VSUBS 0.008047f
C38 B.n10 VSUBS 0.008047f
C39 B.n11 VSUBS 0.008047f
C40 B.n12 VSUBS 0.008047f
C41 B.n13 VSUBS 0.008047f
C42 B.n14 VSUBS 0.008047f
C43 B.n15 VSUBS 0.008047f
C44 B.n16 VSUBS 0.008047f
C45 B.n17 VSUBS 0.008047f
C46 B.n18 VSUBS 0.008047f
C47 B.n19 VSUBS 0.008047f
C48 B.n20 VSUBS 0.017204f
C49 B.n21 VSUBS 0.008047f
C50 B.n22 VSUBS 0.008047f
C51 B.n23 VSUBS 0.008047f
C52 B.n24 VSUBS 0.008047f
C53 B.n25 VSUBS 0.008047f
C54 B.n26 VSUBS 0.008047f
C55 B.n27 VSUBS 0.008047f
C56 B.n28 VSUBS 0.008047f
C57 B.n29 VSUBS 0.008047f
C58 B.n30 VSUBS 0.008047f
C59 B.n31 VSUBS 0.008047f
C60 B.n32 VSUBS 0.008047f
C61 B.n33 VSUBS 0.008047f
C62 B.t1 VSUBS 0.208783f
C63 B.t2 VSUBS 0.235081f
C64 B.t0 VSUBS 1.01357f
C65 B.n34 VSUBS 0.140296f
C66 B.n35 VSUBS 0.083335f
C67 B.n36 VSUBS 0.008047f
C68 B.n37 VSUBS 0.008047f
C69 B.n38 VSUBS 0.008047f
C70 B.n39 VSUBS 0.008047f
C71 B.t4 VSUBS 0.208782f
C72 B.t5 VSUBS 0.23508f
C73 B.t3 VSUBS 1.01357f
C74 B.n40 VSUBS 0.140298f
C75 B.n41 VSUBS 0.083335f
C76 B.n42 VSUBS 0.008047f
C77 B.n43 VSUBS 0.008047f
C78 B.n44 VSUBS 0.008047f
C79 B.n45 VSUBS 0.008047f
C80 B.n46 VSUBS 0.008047f
C81 B.n47 VSUBS 0.008047f
C82 B.n48 VSUBS 0.008047f
C83 B.n49 VSUBS 0.008047f
C84 B.n50 VSUBS 0.008047f
C85 B.n51 VSUBS 0.008047f
C86 B.n52 VSUBS 0.008047f
C87 B.n53 VSUBS 0.008047f
C88 B.n54 VSUBS 0.017204f
C89 B.n55 VSUBS 0.008047f
C90 B.n56 VSUBS 0.008047f
C91 B.n57 VSUBS 0.008047f
C92 B.n58 VSUBS 0.008047f
C93 B.n59 VSUBS 0.008047f
C94 B.n60 VSUBS 0.008047f
C95 B.n61 VSUBS 0.008047f
C96 B.n62 VSUBS 0.008047f
C97 B.n63 VSUBS 0.008047f
C98 B.n64 VSUBS 0.008047f
C99 B.n65 VSUBS 0.008047f
C100 B.n66 VSUBS 0.008047f
C101 B.n67 VSUBS 0.008047f
C102 B.n68 VSUBS 0.008047f
C103 B.n69 VSUBS 0.008047f
C104 B.n70 VSUBS 0.008047f
C105 B.n71 VSUBS 0.008047f
C106 B.n72 VSUBS 0.008047f
C107 B.n73 VSUBS 0.008047f
C108 B.n74 VSUBS 0.008047f
C109 B.n75 VSUBS 0.008047f
C110 B.n76 VSUBS 0.008047f
C111 B.n77 VSUBS 0.008047f
C112 B.n78 VSUBS 0.008047f
C113 B.n79 VSUBS 0.008047f
C114 B.n80 VSUBS 0.008047f
C115 B.n81 VSUBS 0.008047f
C116 B.n82 VSUBS 0.008047f
C117 B.n83 VSUBS 0.008047f
C118 B.n84 VSUBS 0.008047f
C119 B.n85 VSUBS 0.008047f
C120 B.n86 VSUBS 0.008047f
C121 B.n87 VSUBS 0.008047f
C122 B.n88 VSUBS 0.008047f
C123 B.n89 VSUBS 0.008047f
C124 B.n90 VSUBS 0.008047f
C125 B.n91 VSUBS 0.008047f
C126 B.n92 VSUBS 0.017506f
C127 B.n93 VSUBS 0.008047f
C128 B.n94 VSUBS 0.008047f
C129 B.n95 VSUBS 0.008047f
C130 B.n96 VSUBS 0.008047f
C131 B.n97 VSUBS 0.008047f
C132 B.n98 VSUBS 0.008047f
C133 B.n99 VSUBS 0.008047f
C134 B.n100 VSUBS 0.008047f
C135 B.n101 VSUBS 0.008047f
C136 B.n102 VSUBS 0.008047f
C137 B.n103 VSUBS 0.008047f
C138 B.n104 VSUBS 0.005562f
C139 B.n105 VSUBS 0.008047f
C140 B.n106 VSUBS 0.008047f
C141 B.n107 VSUBS 0.008047f
C142 B.n108 VSUBS 0.008047f
C143 B.n109 VSUBS 0.008047f
C144 B.t11 VSUBS 0.208783f
C145 B.t10 VSUBS 0.235081f
C146 B.t9 VSUBS 1.01357f
C147 B.n110 VSUBS 0.140296f
C148 B.n111 VSUBS 0.083335f
C149 B.n112 VSUBS 0.008047f
C150 B.n113 VSUBS 0.008047f
C151 B.n114 VSUBS 0.008047f
C152 B.n115 VSUBS 0.008047f
C153 B.n116 VSUBS 0.008047f
C154 B.n117 VSUBS 0.008047f
C155 B.n118 VSUBS 0.008047f
C156 B.n119 VSUBS 0.008047f
C157 B.n120 VSUBS 0.008047f
C158 B.n121 VSUBS 0.008047f
C159 B.n122 VSUBS 0.008047f
C160 B.n123 VSUBS 0.018536f
C161 B.n124 VSUBS 0.008047f
C162 B.n125 VSUBS 0.008047f
C163 B.n126 VSUBS 0.008047f
C164 B.n127 VSUBS 0.008047f
C165 B.n128 VSUBS 0.008047f
C166 B.n129 VSUBS 0.008047f
C167 B.n130 VSUBS 0.008047f
C168 B.n131 VSUBS 0.008047f
C169 B.n132 VSUBS 0.008047f
C170 B.n133 VSUBS 0.008047f
C171 B.n134 VSUBS 0.008047f
C172 B.n135 VSUBS 0.008047f
C173 B.n136 VSUBS 0.008047f
C174 B.n137 VSUBS 0.008047f
C175 B.n138 VSUBS 0.008047f
C176 B.n139 VSUBS 0.008047f
C177 B.n140 VSUBS 0.008047f
C178 B.n141 VSUBS 0.008047f
C179 B.n142 VSUBS 0.008047f
C180 B.n143 VSUBS 0.008047f
C181 B.n144 VSUBS 0.008047f
C182 B.n145 VSUBS 0.008047f
C183 B.n146 VSUBS 0.008047f
C184 B.n147 VSUBS 0.008047f
C185 B.n148 VSUBS 0.008047f
C186 B.n149 VSUBS 0.008047f
C187 B.n150 VSUBS 0.008047f
C188 B.n151 VSUBS 0.008047f
C189 B.n152 VSUBS 0.008047f
C190 B.n153 VSUBS 0.008047f
C191 B.n154 VSUBS 0.008047f
C192 B.n155 VSUBS 0.008047f
C193 B.n156 VSUBS 0.008047f
C194 B.n157 VSUBS 0.008047f
C195 B.n158 VSUBS 0.008047f
C196 B.n159 VSUBS 0.008047f
C197 B.n160 VSUBS 0.008047f
C198 B.n161 VSUBS 0.008047f
C199 B.n162 VSUBS 0.008047f
C200 B.n163 VSUBS 0.008047f
C201 B.n164 VSUBS 0.008047f
C202 B.n165 VSUBS 0.008047f
C203 B.n166 VSUBS 0.008047f
C204 B.n167 VSUBS 0.008047f
C205 B.n168 VSUBS 0.008047f
C206 B.n169 VSUBS 0.008047f
C207 B.n170 VSUBS 0.008047f
C208 B.n171 VSUBS 0.008047f
C209 B.n172 VSUBS 0.008047f
C210 B.n173 VSUBS 0.008047f
C211 B.n174 VSUBS 0.008047f
C212 B.n175 VSUBS 0.008047f
C213 B.n176 VSUBS 0.008047f
C214 B.n177 VSUBS 0.008047f
C215 B.n178 VSUBS 0.008047f
C216 B.n179 VSUBS 0.008047f
C217 B.n180 VSUBS 0.008047f
C218 B.n181 VSUBS 0.008047f
C219 B.n182 VSUBS 0.008047f
C220 B.n183 VSUBS 0.008047f
C221 B.n184 VSUBS 0.008047f
C222 B.n185 VSUBS 0.008047f
C223 B.n186 VSUBS 0.008047f
C224 B.n187 VSUBS 0.008047f
C225 B.n188 VSUBS 0.008047f
C226 B.n189 VSUBS 0.008047f
C227 B.n190 VSUBS 0.008047f
C228 B.n191 VSUBS 0.008047f
C229 B.n192 VSUBS 0.008047f
C230 B.n193 VSUBS 0.008047f
C231 B.n194 VSUBS 0.017204f
C232 B.n195 VSUBS 0.017204f
C233 B.n196 VSUBS 0.018536f
C234 B.n197 VSUBS 0.008047f
C235 B.n198 VSUBS 0.008047f
C236 B.n199 VSUBS 0.008047f
C237 B.n200 VSUBS 0.008047f
C238 B.n201 VSUBS 0.008047f
C239 B.n202 VSUBS 0.008047f
C240 B.n203 VSUBS 0.008047f
C241 B.n204 VSUBS 0.008047f
C242 B.n205 VSUBS 0.008047f
C243 B.n206 VSUBS 0.008047f
C244 B.n207 VSUBS 0.008047f
C245 B.n208 VSUBS 0.008047f
C246 B.n209 VSUBS 0.008047f
C247 B.n210 VSUBS 0.008047f
C248 B.n211 VSUBS 0.008047f
C249 B.n212 VSUBS 0.008047f
C250 B.n213 VSUBS 0.008047f
C251 B.n214 VSUBS 0.008047f
C252 B.n215 VSUBS 0.008047f
C253 B.n216 VSUBS 0.008047f
C254 B.n217 VSUBS 0.008047f
C255 B.n218 VSUBS 0.008047f
C256 B.n219 VSUBS 0.008047f
C257 B.n220 VSUBS 0.008047f
C258 B.n221 VSUBS 0.008047f
C259 B.n222 VSUBS 0.008047f
C260 B.n223 VSUBS 0.008047f
C261 B.n224 VSUBS 0.008047f
C262 B.n225 VSUBS 0.008047f
C263 B.n226 VSUBS 0.008047f
C264 B.n227 VSUBS 0.008047f
C265 B.n228 VSUBS 0.008047f
C266 B.n229 VSUBS 0.008047f
C267 B.n230 VSUBS 0.008047f
C268 B.n231 VSUBS 0.008047f
C269 B.n232 VSUBS 0.005562f
C270 B.n233 VSUBS 0.018645f
C271 B.n234 VSUBS 0.006509f
C272 B.n235 VSUBS 0.008047f
C273 B.n236 VSUBS 0.008047f
C274 B.n237 VSUBS 0.008047f
C275 B.n238 VSUBS 0.008047f
C276 B.n239 VSUBS 0.008047f
C277 B.n240 VSUBS 0.008047f
C278 B.n241 VSUBS 0.008047f
C279 B.n242 VSUBS 0.008047f
C280 B.n243 VSUBS 0.008047f
C281 B.n244 VSUBS 0.008047f
C282 B.n245 VSUBS 0.008047f
C283 B.t8 VSUBS 0.208782f
C284 B.t7 VSUBS 0.23508f
C285 B.t6 VSUBS 1.01357f
C286 B.n246 VSUBS 0.140298f
C287 B.n247 VSUBS 0.083335f
C288 B.n248 VSUBS 0.018645f
C289 B.n249 VSUBS 0.006509f
C290 B.n250 VSUBS 0.008047f
C291 B.n251 VSUBS 0.008047f
C292 B.n252 VSUBS 0.008047f
C293 B.n253 VSUBS 0.008047f
C294 B.n254 VSUBS 0.008047f
C295 B.n255 VSUBS 0.008047f
C296 B.n256 VSUBS 0.008047f
C297 B.n257 VSUBS 0.008047f
C298 B.n258 VSUBS 0.008047f
C299 B.n259 VSUBS 0.008047f
C300 B.n260 VSUBS 0.008047f
C301 B.n261 VSUBS 0.008047f
C302 B.n262 VSUBS 0.008047f
C303 B.n263 VSUBS 0.008047f
C304 B.n264 VSUBS 0.008047f
C305 B.n265 VSUBS 0.008047f
C306 B.n266 VSUBS 0.008047f
C307 B.n267 VSUBS 0.008047f
C308 B.n268 VSUBS 0.008047f
C309 B.n269 VSUBS 0.008047f
C310 B.n270 VSUBS 0.008047f
C311 B.n271 VSUBS 0.008047f
C312 B.n272 VSUBS 0.008047f
C313 B.n273 VSUBS 0.008047f
C314 B.n274 VSUBS 0.008047f
C315 B.n275 VSUBS 0.008047f
C316 B.n276 VSUBS 0.008047f
C317 B.n277 VSUBS 0.008047f
C318 B.n278 VSUBS 0.008047f
C319 B.n279 VSUBS 0.008047f
C320 B.n280 VSUBS 0.008047f
C321 B.n281 VSUBS 0.008047f
C322 B.n282 VSUBS 0.008047f
C323 B.n283 VSUBS 0.008047f
C324 B.n284 VSUBS 0.008047f
C325 B.n285 VSUBS 0.008047f
C326 B.n286 VSUBS 0.008047f
C327 B.n287 VSUBS 0.018536f
C328 B.n288 VSUBS 0.017204f
C329 B.n289 VSUBS 0.018235f
C330 B.n290 VSUBS 0.008047f
C331 B.n291 VSUBS 0.008047f
C332 B.n292 VSUBS 0.008047f
C333 B.n293 VSUBS 0.008047f
C334 B.n294 VSUBS 0.008047f
C335 B.n295 VSUBS 0.008047f
C336 B.n296 VSUBS 0.008047f
C337 B.n297 VSUBS 0.008047f
C338 B.n298 VSUBS 0.008047f
C339 B.n299 VSUBS 0.008047f
C340 B.n300 VSUBS 0.008047f
C341 B.n301 VSUBS 0.008047f
C342 B.n302 VSUBS 0.008047f
C343 B.n303 VSUBS 0.008047f
C344 B.n304 VSUBS 0.008047f
C345 B.n305 VSUBS 0.008047f
C346 B.n306 VSUBS 0.008047f
C347 B.n307 VSUBS 0.008047f
C348 B.n308 VSUBS 0.008047f
C349 B.n309 VSUBS 0.008047f
C350 B.n310 VSUBS 0.008047f
C351 B.n311 VSUBS 0.008047f
C352 B.n312 VSUBS 0.008047f
C353 B.n313 VSUBS 0.008047f
C354 B.n314 VSUBS 0.008047f
C355 B.n315 VSUBS 0.008047f
C356 B.n316 VSUBS 0.008047f
C357 B.n317 VSUBS 0.008047f
C358 B.n318 VSUBS 0.008047f
C359 B.n319 VSUBS 0.008047f
C360 B.n320 VSUBS 0.008047f
C361 B.n321 VSUBS 0.008047f
C362 B.n322 VSUBS 0.008047f
C363 B.n323 VSUBS 0.008047f
C364 B.n324 VSUBS 0.008047f
C365 B.n325 VSUBS 0.008047f
C366 B.n326 VSUBS 0.008047f
C367 B.n327 VSUBS 0.008047f
C368 B.n328 VSUBS 0.008047f
C369 B.n329 VSUBS 0.008047f
C370 B.n330 VSUBS 0.008047f
C371 B.n331 VSUBS 0.008047f
C372 B.n332 VSUBS 0.008047f
C373 B.n333 VSUBS 0.008047f
C374 B.n334 VSUBS 0.008047f
C375 B.n335 VSUBS 0.008047f
C376 B.n336 VSUBS 0.008047f
C377 B.n337 VSUBS 0.008047f
C378 B.n338 VSUBS 0.008047f
C379 B.n339 VSUBS 0.008047f
C380 B.n340 VSUBS 0.008047f
C381 B.n341 VSUBS 0.008047f
C382 B.n342 VSUBS 0.008047f
C383 B.n343 VSUBS 0.008047f
C384 B.n344 VSUBS 0.008047f
C385 B.n345 VSUBS 0.008047f
C386 B.n346 VSUBS 0.008047f
C387 B.n347 VSUBS 0.008047f
C388 B.n348 VSUBS 0.008047f
C389 B.n349 VSUBS 0.008047f
C390 B.n350 VSUBS 0.008047f
C391 B.n351 VSUBS 0.008047f
C392 B.n352 VSUBS 0.008047f
C393 B.n353 VSUBS 0.008047f
C394 B.n354 VSUBS 0.008047f
C395 B.n355 VSUBS 0.008047f
C396 B.n356 VSUBS 0.008047f
C397 B.n357 VSUBS 0.008047f
C398 B.n358 VSUBS 0.008047f
C399 B.n359 VSUBS 0.008047f
C400 B.n360 VSUBS 0.008047f
C401 B.n361 VSUBS 0.008047f
C402 B.n362 VSUBS 0.008047f
C403 B.n363 VSUBS 0.008047f
C404 B.n364 VSUBS 0.008047f
C405 B.n365 VSUBS 0.008047f
C406 B.n366 VSUBS 0.008047f
C407 B.n367 VSUBS 0.008047f
C408 B.n368 VSUBS 0.008047f
C409 B.n369 VSUBS 0.008047f
C410 B.n370 VSUBS 0.008047f
C411 B.n371 VSUBS 0.008047f
C412 B.n372 VSUBS 0.008047f
C413 B.n373 VSUBS 0.008047f
C414 B.n374 VSUBS 0.008047f
C415 B.n375 VSUBS 0.008047f
C416 B.n376 VSUBS 0.008047f
C417 B.n377 VSUBS 0.008047f
C418 B.n378 VSUBS 0.008047f
C419 B.n379 VSUBS 0.008047f
C420 B.n380 VSUBS 0.008047f
C421 B.n381 VSUBS 0.008047f
C422 B.n382 VSUBS 0.008047f
C423 B.n383 VSUBS 0.008047f
C424 B.n384 VSUBS 0.008047f
C425 B.n385 VSUBS 0.008047f
C426 B.n386 VSUBS 0.008047f
C427 B.n387 VSUBS 0.008047f
C428 B.n388 VSUBS 0.008047f
C429 B.n389 VSUBS 0.008047f
C430 B.n390 VSUBS 0.008047f
C431 B.n391 VSUBS 0.008047f
C432 B.n392 VSUBS 0.008047f
C433 B.n393 VSUBS 0.008047f
C434 B.n394 VSUBS 0.008047f
C435 B.n395 VSUBS 0.008047f
C436 B.n396 VSUBS 0.008047f
C437 B.n397 VSUBS 0.008047f
C438 B.n398 VSUBS 0.008047f
C439 B.n399 VSUBS 0.008047f
C440 B.n400 VSUBS 0.008047f
C441 B.n401 VSUBS 0.017204f
C442 B.n402 VSUBS 0.018536f
C443 B.n403 VSUBS 0.018536f
C444 B.n404 VSUBS 0.008047f
C445 B.n405 VSUBS 0.008047f
C446 B.n406 VSUBS 0.008047f
C447 B.n407 VSUBS 0.008047f
C448 B.n408 VSUBS 0.008047f
C449 B.n409 VSUBS 0.008047f
C450 B.n410 VSUBS 0.008047f
C451 B.n411 VSUBS 0.008047f
C452 B.n412 VSUBS 0.008047f
C453 B.n413 VSUBS 0.008047f
C454 B.n414 VSUBS 0.008047f
C455 B.n415 VSUBS 0.008047f
C456 B.n416 VSUBS 0.008047f
C457 B.n417 VSUBS 0.008047f
C458 B.n418 VSUBS 0.008047f
C459 B.n419 VSUBS 0.008047f
C460 B.n420 VSUBS 0.008047f
C461 B.n421 VSUBS 0.008047f
C462 B.n422 VSUBS 0.008047f
C463 B.n423 VSUBS 0.008047f
C464 B.n424 VSUBS 0.008047f
C465 B.n425 VSUBS 0.008047f
C466 B.n426 VSUBS 0.008047f
C467 B.n427 VSUBS 0.008047f
C468 B.n428 VSUBS 0.008047f
C469 B.n429 VSUBS 0.008047f
C470 B.n430 VSUBS 0.008047f
C471 B.n431 VSUBS 0.008047f
C472 B.n432 VSUBS 0.008047f
C473 B.n433 VSUBS 0.008047f
C474 B.n434 VSUBS 0.008047f
C475 B.n435 VSUBS 0.008047f
C476 B.n436 VSUBS 0.008047f
C477 B.n437 VSUBS 0.008047f
C478 B.n438 VSUBS 0.008047f
C479 B.n439 VSUBS 0.005562f
C480 B.n440 VSUBS 0.018645f
C481 B.n441 VSUBS 0.006509f
C482 B.n442 VSUBS 0.008047f
C483 B.n443 VSUBS 0.008047f
C484 B.n444 VSUBS 0.008047f
C485 B.n445 VSUBS 0.008047f
C486 B.n446 VSUBS 0.008047f
C487 B.n447 VSUBS 0.008047f
C488 B.n448 VSUBS 0.008047f
C489 B.n449 VSUBS 0.008047f
C490 B.n450 VSUBS 0.008047f
C491 B.n451 VSUBS 0.008047f
C492 B.n452 VSUBS 0.008047f
C493 B.n453 VSUBS 0.006509f
C494 B.n454 VSUBS 0.018645f
C495 B.n455 VSUBS 0.005562f
C496 B.n456 VSUBS 0.008047f
C497 B.n457 VSUBS 0.008047f
C498 B.n458 VSUBS 0.008047f
C499 B.n459 VSUBS 0.008047f
C500 B.n460 VSUBS 0.008047f
C501 B.n461 VSUBS 0.008047f
C502 B.n462 VSUBS 0.008047f
C503 B.n463 VSUBS 0.008047f
C504 B.n464 VSUBS 0.008047f
C505 B.n465 VSUBS 0.008047f
C506 B.n466 VSUBS 0.008047f
C507 B.n467 VSUBS 0.008047f
C508 B.n468 VSUBS 0.008047f
C509 B.n469 VSUBS 0.008047f
C510 B.n470 VSUBS 0.008047f
C511 B.n471 VSUBS 0.008047f
C512 B.n472 VSUBS 0.008047f
C513 B.n473 VSUBS 0.008047f
C514 B.n474 VSUBS 0.008047f
C515 B.n475 VSUBS 0.008047f
C516 B.n476 VSUBS 0.008047f
C517 B.n477 VSUBS 0.008047f
C518 B.n478 VSUBS 0.008047f
C519 B.n479 VSUBS 0.008047f
C520 B.n480 VSUBS 0.008047f
C521 B.n481 VSUBS 0.008047f
C522 B.n482 VSUBS 0.008047f
C523 B.n483 VSUBS 0.008047f
C524 B.n484 VSUBS 0.008047f
C525 B.n485 VSUBS 0.008047f
C526 B.n486 VSUBS 0.008047f
C527 B.n487 VSUBS 0.008047f
C528 B.n488 VSUBS 0.008047f
C529 B.n489 VSUBS 0.008047f
C530 B.n490 VSUBS 0.008047f
C531 B.n491 VSUBS 0.018536f
C532 B.n492 VSUBS 0.018536f
C533 B.n493 VSUBS 0.017204f
C534 B.n494 VSUBS 0.008047f
C535 B.n495 VSUBS 0.008047f
C536 B.n496 VSUBS 0.008047f
C537 B.n497 VSUBS 0.008047f
C538 B.n498 VSUBS 0.008047f
C539 B.n499 VSUBS 0.008047f
C540 B.n500 VSUBS 0.008047f
C541 B.n501 VSUBS 0.008047f
C542 B.n502 VSUBS 0.008047f
C543 B.n503 VSUBS 0.008047f
C544 B.n504 VSUBS 0.008047f
C545 B.n505 VSUBS 0.008047f
C546 B.n506 VSUBS 0.008047f
C547 B.n507 VSUBS 0.008047f
C548 B.n508 VSUBS 0.008047f
C549 B.n509 VSUBS 0.008047f
C550 B.n510 VSUBS 0.008047f
C551 B.n511 VSUBS 0.008047f
C552 B.n512 VSUBS 0.008047f
C553 B.n513 VSUBS 0.008047f
C554 B.n514 VSUBS 0.008047f
C555 B.n515 VSUBS 0.008047f
C556 B.n516 VSUBS 0.008047f
C557 B.n517 VSUBS 0.008047f
C558 B.n518 VSUBS 0.008047f
C559 B.n519 VSUBS 0.008047f
C560 B.n520 VSUBS 0.008047f
C561 B.n521 VSUBS 0.008047f
C562 B.n522 VSUBS 0.008047f
C563 B.n523 VSUBS 0.008047f
C564 B.n524 VSUBS 0.008047f
C565 B.n525 VSUBS 0.008047f
C566 B.n526 VSUBS 0.008047f
C567 B.n527 VSUBS 0.008047f
C568 B.n528 VSUBS 0.008047f
C569 B.n529 VSUBS 0.008047f
C570 B.n530 VSUBS 0.008047f
C571 B.n531 VSUBS 0.008047f
C572 B.n532 VSUBS 0.008047f
C573 B.n533 VSUBS 0.008047f
C574 B.n534 VSUBS 0.008047f
C575 B.n535 VSUBS 0.008047f
C576 B.n536 VSUBS 0.008047f
C577 B.n537 VSUBS 0.008047f
C578 B.n538 VSUBS 0.008047f
C579 B.n539 VSUBS 0.008047f
C580 B.n540 VSUBS 0.008047f
C581 B.n541 VSUBS 0.008047f
C582 B.n542 VSUBS 0.008047f
C583 B.n543 VSUBS 0.008047f
C584 B.n544 VSUBS 0.008047f
C585 B.n545 VSUBS 0.008047f
C586 B.n546 VSUBS 0.008047f
C587 B.n547 VSUBS 0.010502f
C588 B.n548 VSUBS 0.011187f
C589 B.n549 VSUBS 0.022246f
C590 VDD2.t3 VSUBS 0.135984f
C591 VDD2.t0 VSUBS 0.135984f
C592 VDD2.n0 VSUBS 1.38058f
C593 VDD2.t1 VSUBS 0.135984f
C594 VDD2.t2 VSUBS 0.135984f
C595 VDD2.n1 VSUBS 0.928383f
C596 VDD2.n2 VSUBS 3.78354f
C597 VN.t3 VSUBS 2.26216f
C598 VN.t0 VSUBS 2.27329f
C599 VN.n0 VSUBS 1.38003f
C600 VN.t1 VSUBS 2.27329f
C601 VN.t2 VSUBS 2.26216f
C602 VN.n1 VSUBS 3.3616f
C603 VTAIL.t3 VSUBS 1.13822f
C604 VTAIL.n0 VSUBS 0.738803f
C605 VTAIL.t5 VSUBS 1.13822f
C606 VTAIL.n1 VSUBS 0.862568f
C607 VTAIL.t7 VSUBS 1.13822f
C608 VTAIL.n2 VSUBS 1.93599f
C609 VTAIL.t2 VSUBS 1.13823f
C610 VTAIL.n3 VSUBS 1.93598f
C611 VTAIL.t1 VSUBS 1.13823f
C612 VTAIL.n4 VSUBS 0.862564f
C613 VTAIL.t4 VSUBS 1.13823f
C614 VTAIL.n5 VSUBS 0.862564f
C615 VTAIL.t6 VSUBS 1.13822f
C616 VTAIL.n6 VSUBS 1.93599f
C617 VTAIL.t0 VSUBS 1.13822f
C618 VTAIL.n7 VSUBS 1.80177f
C619 VDD1.t0 VSUBS 0.137871f
C620 VDD1.t3 VSUBS 0.137871f
C621 VDD1.n0 VSUBS 0.941713f
C622 VDD1.t2 VSUBS 0.137871f
C623 VDD1.t1 VSUBS 0.137871f
C624 VDD1.n1 VSUBS 1.42072f
C625 VP.t2 VSUBS 1.95304f
C626 VP.n0 VSUBS 0.881316f
C627 VP.n1 VSUBS 0.039732f
C628 VP.n2 VSUBS 0.057757f
C629 VP.n3 VSUBS 0.064117f
C630 VP.t0 VSUBS 1.95304f
C631 VP.t3 VSUBS 2.36589f
C632 VP.t1 VSUBS 2.35432f
C633 VP.n4 VSUBS 3.48199f
C634 VP.n5 VSUBS 1.98314f
C635 VP.n6 VSUBS 0.881316f
C636 VP.n7 VSUBS 0.067496f
C637 VP.n8 VSUBS 0.073679f
C638 VP.n9 VSUBS 0.039732f
C639 VP.n10 VSUBS 0.039732f
C640 VP.n11 VSUBS 0.039732f
C641 VP.n12 VSUBS 0.057757f
C642 VP.n13 VSUBS 0.073679f
C643 VP.n14 VSUBS 0.067496f
C644 VP.n15 VSUBS 0.064117f
C645 VP.n16 VSUBS 0.082072f
.ends

